`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
sWumofZYST6mcnnY+SwyRTvh77swIBrhjt/XKPTEp5kzCOV6F9FKQgFe4oGFWYqfN2TJmqipIKDr
R0JoZRTteE1al1+8iorfqNN5u85DMU9vxwr3iVjrtAb1hSgtkkk+rhEMP6C2sthttnexF78MuEBa
cl4heg5wmxvY1vVpWI2mQ4WJMTtgaWSeh8hQlT7MaqIfS8L0KxVgj63tO6ivIsnAilzak/TWvVbR
0vl1ukC7LMgyxTkixTuiNQyJVv9XJLyKN8CPgPAA6fYAiJMP8KHDu1T4LRLuLrv8+4oYod+Bg7EG
g1+5G+Rnh8KvNRALo2EfDoUq5/L4MIuWANLPiw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="VxNWF8gxYv9utWUJQAsXldcuC6C1Qjy/t171FHbtcSA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18368)
`protect data_block
gCtg/3wX+DuoyCjZcOi5uP81HeRv+/sX79418JDbrCnbymoKwk54RmYqotoYEK0hz7n1LknsoapC
rT7oK3PchXgiGHoWDg7dUDJSt4itJy8MGnCySlH4Cu9QZ66NQsSvfdzBMNb5tyF2LURDv3wEu9Ww
Y+rOh4aFww6cYcoHQzyZGo/QuavMS4Ih/yi2IRv5DeuZT01MhNVc+8n5PRGdAfyxNiiclUt4uDdL
PI29gVxO7KTjf3jUBOLV1kWnVcVPGJg8b/EvlBXiZl9uKV5ekHEXcuVUNo0g5PhLHCVom51qQOqv
ZTpOx5QDB12x116uyAmvLcIE9aZ5V95v5UrRtekrURjhTXo3E9nEnNzexs/gfj6VRFlekq9p73xl
70udWJrZJSt7Gj9a3VwCkfY81//YnCVhD+/Yrz7W7dO9XTHv3CLOIEuzcUThb3Dfkv63+F+J3o9j
ai30VPa2KqzOh97ivITGvMbsGIEBC0wH7uC5y7PqlRPXGzkwCqvkLFKSXqbgECC0kzm/HR6Ob88z
lZZG6o/GamhcWWN+tl7xNyQQ/lDZbbhvdmWGC/QFKe9Zm4sCFbythJMFlpmxtyUu8JRwMjaLaJHQ
A+wYOJ2bNfCLWFvKmrpnZqAf5P2cAkOnwh5zLsLI4u8xDQWpe93L6iG+TXu/GQt5SQeah/goFo7A
LUHKn37KdYXdNj6GNDHJLteph4LDqRegqqD4K/jrG918ZRREFFNc3YrcNwXWZ7iwWqMgYVqCtklp
HW4u3Kq1wBF5hkqFCN4enjco1by5cbPSA/BnZf1dIVtgnZXNHwTkbMpmQpRlIUkP2F6UrerdpZUW
Tx9vcL94kk9Olg+I6Xlj3qrc1M/qGFmQ1JnBU045tB5HtuWhGbChw+JLKXJ+eOv7e+cBtinM8TGD
ijP+ZCF4cHvbw93RSiex9LZ9mWQS5Fow41wKOdpiqDKAiBSifh2Kq5p+wqfYMZzyaan7TSPNlqMS
gftSFa6Hd56b4NEkS5NntDXw9yDpyp3yrEDhmlYjuOpJXcbvRqnT2gQ522+/u1AYgHwpOavL+IIA
cBZGf1lgb4r3EJIxl3y5FpyVoK2iWRq71MqY1gMR1SexSr5tzEFRMbxe+teBmK6Z00bBNSBaaWAo
YGr3RJgDkhnnZkRFGvWQX4d9WJeRHSRdjxHgxeX/7RqDWNLSo8f1Zrd7xQkrQgbn4H3yCXGCARhP
e3o0VJ08Wck7TdzhFZ5h7qaM2Ds1hJItkvguri15FO+83YR9+D0UnxYyKNXfclbtb8eNuOLGTPrg
lNbHWYcyr6FEnJ1YugASHfVGZyIbtMWwbyB4APv4/5OOobx3rCwCsha+P5fZfXvClRWqLpdEkjro
8rx5pKB0Yx91cROMTgwkKgssBQ1UjP6qu9K6MS7SSzIT2DqrrkF0l/A3cTAxVz2XS3YksWVPfIh+
3rYRx0ndHnevqb+suV3pEAayauSvKHZQh6yQ6g5rScHGmeptgYWPcTO43g2VZuh0LDGrPDj3sd3q
K107hfEL0Izzp4nzC1HNbaIFHxgMin+pHm663r1YRo9hH1KVRLSFqsx/7dUdi5oPNAo+8SFU6bn9
3hJF4qkFCVo+lK/yGtCheontkB/oOaIFFoyWnjh21cdKjbQkFFdHvc4N0b7Ae3cxIVGqGNRdZgA/
PdCdHBCdKm1fu26eLUOVrq78MS1+5nyQLrTMmf4JH7SCwulWbgadKDS/1XYTN77B0DC5Pgmk2/Tq
cWwSysiqU0m82ofxKrA/PcAoguD1Ba/V91oOAN4AbxNanfBAbptxTDr4zDWi5unXQWGNUXYbi4jn
QVMv9h0iu+JafXzU+z6ZVkCq6qJMilp3uTK5QMohdgUyd32cvbKNtZS60O6aKo/oP08NeTZtLEbD
zdl4DqXd+jLXW3kF8oS6+8OmO1o2dpotUJwNeZjkV8Zq/AsYJuWw17DaHeTeIomx2QBNxz9Jnqu/
2+s8cZCb714a/b7sj4NFfNTIeGG9bgRVBFZFuiEmyNzbDz/6Jwra5lV94rXB5ZedN6VX/iReiTQG
uv4He2K0K5S0OtKh/bRshdJszWvKyC6z9k7OXx5UYWaorrBJeLlBjeYFjIWdINAgL3Sr4LRolFZz
O7Q+ohqtbLSIvo/6kXYR6dLlaRQrnp1nrxtzqoclMLLNLM7+5c6Oa2OJORraUt3h3YxFCY0XwW70
7UPi433mDD2e05lCrzxjcT7awXfGJjsv4KDMcPf0a+zrqMGLHrpFu4Qdsl3tHvv+NWLIpnYy9wPL
lWFcFWTFwfR/qFLfkIPqy+fiA2cqGd5P4y322uGLGOHbuSNNt5kwyQG8Dq4vxPBgFiGxWTd5gQG2
+apcec9ealh7mFSuhzjjBsT7w/baiImD3tH9DGDthMs8MbSlbg4gC8YYNgaiAInR4YBAXmJ1lURV
C1w8Y6cHryLArLlXWKGJ4OWIGon5V3hLsBUyNGBtfPdmnl9XpteoXrfTnrkZzLJbCx6L0XG9V4jF
JIZNDi0CDbnjAmDP/iz24TMyPfjRmusCjOwwSR2UQHJ/AstHEaymzzA2dN7WdXcL/FYqseVKHTc/
neTPsne0OEgXZQZfBRxEWNL9b2mMl7l0XQxQ+kJFP+FI/LoLiqh1n3Q89rxSL1iQZLZJ3jeTTg1s
n6PNlxUEIfMKqKSVW4Sih3BR5l/1OcuGVjSHKe6EIwafbUR7nBD+IHKpfXXbkzj1360Eo8cComAe
juOXjyjh0ifxWfPd0E+FMATNIJ2YeXKStdpxGC1pQ4Eh5oR4u903we/8wNGwZI5EUdQFzIPGKakp
UPUut+g3rLV5rX7md6naQtP+dbx8hc4vbKvsuCgIniZVXzfGhGcSLec8s/rD/EoDNIsCJYGoYP+G
Eju2gJuBUlA+fgSqnM/lTiyRneE34Ft5b6IRFWWmYaqMa8XYFDY+m/F+kYx3F/junowXuq3bKI51
t/HOGQmDS2bvXR/3SoxA7DXyaA+4n557iBKwEoGYUUXGgI5C2DqawAle3Ha2LTgQ+6JuNir0o6Qb
vduHSgIy/4oam9OO2KX/2jMhdamfEx+wDiuiuZ3jvMvvO1DuNnSREAjrnFvfuDW73WHP2My1beEf
BcVvXdm/AhSbo5G4h3+jIA01x8dn8z//8zs9WhmUwTJwc4KbSF+dM2WCwfNwwvljKWvyF7d6U255
9j+3ncOZ4DJSkjzkHwo5JAP8ZqJMRTCgjD2Qf4pyEkcpqrW/AmJGYefXGQn7xuCaMQ1Bqlys4jUg
V9U7BLcGS3+zJ2OGt/B5Tz5QB8+ynedKVN+OTA6H5tN+rcxBTy4tXeAlvpQo4lmQs4fnlys6t2P+
jY83kv/iaqeZ5K8JAbDGxZzX2D1n0OBRlYtmpzSOHZbGyxTxGLl40a6+akjj3D3xYAKH0BDWVsnj
UbEyzH+ZTPmZDioZyImLlx8cyECQDSW1KPLglJfM5/j5Tb/yDQNzYa8Wq0Qvzwj2bWFA4JYR0dPB
S6fyzCXiJ3H/hFoxKgfUVjKVW5HFgSCTWCo8abEA/PT1LHrbcindm4UAAvEaQMmgR9xxj7O2sLm6
pl7pEWr2Se0j52wXvsili85hGTQzfs8h0HDPdj/hUxBmQs1PbYYexv5xDt2NmJEaNHAWKbYH2551
r9howBw54MymjqBSIZ4JTLYSdrgpwE3evksx2okJkOmaW+fyky4yatWso27qfKly5ljOjZ74JoZO
pI7nGbAcroyMUdYEiF+OClidGFA9kJYC5Lge06ivKu/eK65xJyofFLIXuGLuFacVyxEsRjMQOB+H
nBrfQROx0oDg90oNd7YPw6ZENXq8hV4fxgz5PM0JzSiwFZ+EZP8IE12Ucu7uhBI908OjGoKMXEiN
eyzjeSqYzBnJjxYsXRsoP25tvz1/zmIrxDDWyZsmdX9DIHv8TTGniZYIOs2mwQsdZkHx/g9lrqnm
gG377qO0OEd4RXxgnBZN8324epeAOGWqCCCxEieRMJNOXVLLKzs8zduAwGD3KhwA4IHeU4sdg3Fj
LWDDt1PnCw8NaIya/F+pl/TqStIY8BtoTR8zu67lGOpMyC7FaQQhH0GMd4iAXVSn9VUyhCp+VLwZ
o0fNVLkiqzhPTi0SIjcayW1dhlnFfBy4ECGPv4G2ivtT3Ug1nTYBb2RZ1avcCICG64JhiCIIGYKG
N7SFxumSZK/zVh6i5T6XPFIWHRvWMtvNd+hoBLGPli5hn1OAUNMnR9j8UWSxPN8XjxPXH06A2yB6
0gSBOY8j1lfTiN9771GYyqhW/kfpxPF8S7TV9QJKG6DHRaMkejdnUYAa4wmPsKEsKoMCqNILnRqT
QnlkO2m3nYdY0TFdG3hBj2CcULDUIQIncyNRunOoHHRoZYNi8eLpRokM2YvXZMq1L9t5BT0ljyLZ
bl6VhTN4y6AxE4SsK7Mgop45LC1Dn/tpjtK3pYK8ptD+qg8YcSB/kLtkbc2P7q0H9XfmSdksgXtg
+ENeZWf4DZrnrCxGCC3hgXqmal5FoOIR7jg9ie78sfGvUNwb3AgosCydfZe9hGFgQpyf3sY5ckLg
pT7m3qxjZdKQvMEbboBOKIVQd3Cl+XI+H2FugmGSFuQcabI9ZXYC32nbeGhvQF5DVdb501Q2qM8Q
M8oudkmfDCl39k3c3deX8YQA4wqVy05DuCQ3fVE6bnoSsXBEusIHuLzE9hXTn4ePizTJDSYK4t+P
8jLnBraYi0Z/Fr1IY9+H3byqG8osBvdKQqf8b5CfagOjAsPhWZg5dEnNiW5zn0tp10BiesVuC3qb
HUBVDMdyCWIwIKU7tO0wClP0XuND8BX6l1AtOwQ2xPNKxcJRcqpepoRAqHgQbsw+dzlPQyX5qT1g
/H6sZx3tXh78kh9pw6mmg1xKvMkMtEUPSgxYpxB+cNXo2rIIKZDR6SuZgAIceE3woorKDXMEmz5Q
uFeCDnH3CH8/MS2eWQyMj2avBJYJ1zN6Iz38b2hRJ/xc1NMsu+BCUs0DTP495QwZDcOBwnLcfbaP
wWWL33iWY02DFm/Ns3RUKlZMxKQ/W++1w21KvBHIoonY1YwnWtoQyBceruInzKdfF3UwqD8OMGqb
fE3r3Vkua6+c1BlyYz+YP47WF49cX6EqlR+3eLxD6YD0RHY3r3FqXdHFHoVtc7ZV+Axal0pQXxxv
HIbttc1xrXkh0UQwephKD+0wb7ShwccIzEzGi33EQ6APP1xW6Wr+FB7mNmZLtzpMMwkZ5U9fcl0r
Qs9shjqIRa29yYq4FhRNd5nwEOawFhjl3MlYx2wqhcRY/jAlAyab8w1307hPqDPK5EboFiz6oJlX
VtxoGkEcppC/oG0KCbwSupK34liMnfkE30SyG5O055G6QlO4jvKN23cZuf87olXP3PJtM9tNlCab
pkX64J+AzAaPqJV9lF4xJIYPAhHiTtQqYdXQmVjIFOlCvLbKL1nxKQ/rxxQ9S5XQB75Y7jR9Bnwk
tcucad2l5lIPr+PQctsasoGroiJx3zskG3ZO5dq+1t+64j8YkopUZGzHyN0yram2KtYYfs5hkBKD
L4SktXnYe6T+mDPvyDskVoa0yW3Ksru1j9UVqZw4sv6EuXlclEvwTY57RT/XrXewTHJ/9Ml8eetf
6u2iXUCeea2y4yD1ceKdfT7MZaOzyDouivOiLV2lsFCX1dVQIMK4+md4UOVAjxkzdntro/zlbEhX
frJdcgbJHRqfO9reRIWEEIZ82+X0u4AMnHIwRVaQtRfyCnaXuw4fYqtgNZwF7LqIEqGTZ9yz5/GQ
mDKMrcZJj+TBwDkkljLEhnJ2hyGfRdWCXKFvf1KHYyzcJiZ7qeUl3o5w6BluLGAEelqAbX5VcQYg
EGxsG49tTY3uGTh+mkJloGDfq2sa7bn7dALce85P/9SX6eeIMaogZ8RWPUUxW1WoOxhH0qn6lw5f
5why9sb0ioMu9NQBK2xpwRassQSwzSly6wYKt22BO92Xv4nPCzcSdaSjWFO2h5dtWNLZhXlpcZ1Q
EbKDsSwFbk465+1SuIZl10OEh5cINUmLbvsCUSg0g3iuq3dIW/vvw+O+2lXXA3ipx76qaC5an+k2
fEIBplnYeXbL29tfe8BpPk3WvePfdPIQaDsjjwzjBZawkfd3GwT1NDF17vo34PJcm3ylP4QRO67x
+qTo5TukE1KEMCwkzVlaI2I9SyOV9cEYW5U5kdngDgE1Dbdr9UyiNkFEF9+dcBdhXjECeyt5CNXU
dI3ArnSP0Um/KLn8IsHx+UVazeDxUvk3QqE3mYRt7jK5RJ6+Psgv/bujzYNAU8QejiUogwxap21H
9xcxp0+VLaTdgDzeSXAvZevn0h0PM53DI7MuJ7INN4k732pIVKQiMT9QSYhb9qhkMlTzZqKEmJWI
9/7gO9gUPnNBQobFP0UZG4cFuh3CcujHIXjPKtHP1OEW4eGbWDXKWHRQCtWhjfCh69Cb5WSU0NMq
Jgt+vrUtPNQbGeDpHNeSBxaCNQLzsDgTBKp0wculRGVduvZh6AttIbfjap+R3B7hhyCpIlkwuACu
bbqJQFg8WkDRYq0+ocAQ5sH+SyqRvBPAjnqfVv4GGg9l/XAGc9CSkv+92/BXB35uUNk5lJULpPQU
mxDwA+oBWGVurlpU19SD9brIbesfG+oIe8Ma+zHoVJU7JiIeFPdzWgrYyGnw0ngPbTtjnCHjml7y
5WlCgEnk+tv0gg5f3f183smRJZxo4wWPZeiOBg5/5ELc6V5YLbauGpDXAYEO1OyuMI0JPY08HeTY
qwhARTdPx770mojOLC+MCjF9+qvPa6osfDu3veEn30qeOfTG7KKFEsOWygbWhs2UeOsLmTDnE3JI
TjOMAFxEPykZQroo3Lrp8MLqzCqQnaU8ZPDOIJ1mFF5h/ItYQ5BVKUbLhnbIWL2o5PpOKnaqGooa
G+3BiOBolZPDzbMeR6j2JfcfKVbUQqV3fpiYQB1+wsXsG6/al2FrgMVgnDMLtSsSGcFxHKH/+xWP
iTuPh0bQhDkBHxSKRhWY3FcQEcr93+GffHOS3MPKphb7T42gqSv6Qsi2cZJXuNF8d+NNcGpfFJyx
9nk71oQzulwmdle8VCzOqMspkx9mx5L0/ihl1AoQZosJJBsYvgBwkThX31ieAL30/ffhtHUzZMxq
PFm0VNxpg7G2yHKdL1f/Wt9ykE0hjvFFQ74e82LS0JnXIy4vqJ/tCjwogWQD7E8iLWeZbatuQpKH
hBejHhCWaaI3qT3m9YOTi2JwcgU2HLAp0QNpNU3DMEnsuLutQajM6lT43E85PIbdJY8DXlak4JpL
FM7kmC3vkY1LgocZ5A++LRG7JzvYN3kkJ81jRaIyPjbozw4xEErOeuHdTnlNkIDmF5OjH1qo/Zbq
maaWggHnK+hCcJKxtWexphijvCa5uhUx0F/pnlzkZGCj1t0MzQXcf8V3bsgJ5gMT2PJkhF/YTApC
3sVvNjOt4QpPNxZ8mgC1Ky6dAAJwqlfIhDqnD3S4/tRIAiA0yUF2SG1Vb59ROzC2CgKNIklNp45P
jZ/g5MgAgYdfT6sC+cdO9Z9XVaMdDn5ccdSZip3v3jEy2KjOlAg+6CmN42rbAz+8N497Gh0SGFYB
Bkli+dafRY+4eChg8FKWAxnS81/ivwDoSy+oYQjSQHRk7nkL3WvhvBXUA59zltmaFB77Ek1B0srh
x9Gf0jabHWZD4hExGrfx+pASpml15f0wOx1bqElPGTOAKvA4k/DwkjP/gaqF6Vm9u9aJUb1er2hA
33ZoxThp66yofx0kYdfljXFE9raHx7iUrVEiKOMHVepqsrA5Y4XimEkOcphaB6Nr5kxOpDYFO+Bn
4agAwXkPTqWvHun9m3FXVn9zMc/0yjVTQG0HAvg2/0QdNLHMtv1RyAOcPizDHbUTaYdlmLfD4tPs
h9p89BHrYIi7Hyfo0RrspBGiGPXYYsQ98m2AZ0M2UQsVyd6Yk/MkiCz+/0UU2OQUMSTbXsOU4w/E
NlgxAtGNbuDjJLRboiIxBsT6Ksg+Zi9VnaYzjVhIdQArv02EEhkkOsXbfY7cpo/NpI5U0eUWvr09
HbDNgvJlLy8/7RaRWT0/uqcMjBpPLikaj/qcDCJdh84xlNh892BF5Ntu5vAn3Hzt7hjejL1geAe8
bUoVdMnp7d93Bi5UAjJMtOmZAt6dAiRmx+mKJazzTW9RbQzEvQnr0MvLR+9qzl2F2z3V0lDgfrB/
MwqmZX6tRqCoNqUIruFIvqiMzYx1PUKT+qZyDHEBynvT+5oaPsvkCeCLCjS14GUZtAHI3jndJnbV
cLNQ+biWwIVnk05pL16u0VI7GEDi8J7k5CsL9mw7GEaTNzbUZFEyIo0YfzWIpIQLVbl93P337tFc
om8QJWdgbanUc4HwDcAkXc49n9KaxFnm6Q3ejowOL3D3uUr6t/mg9OA04T0FdZjyr9dfYxax/je2
HNqhjuHRg1g8rYUFLcmEv5l+OfEFR3ZKZIqzbcgm4e/l4QGx/BWiojeeOfsKBB1soR8qWjHHVTRe
JFogwPhJaFgy2/Fi3FAUmcfYNq71dS4OqXEsIroWYXBpSegujH+geERFb+xfkVXCxBUgXx8RoftP
oVFjM3CSX05K646mPgj2FxSHThyLQGyFrUyKPPXSDpyIB/zXbjXy9L6bVu7FvEi0UjJLJ8XUtAiz
PDWifLDdWp5nPn9F/XItPQD0Jcml/mT/TTq+lZaf3c+RiqGOq+ztMO0jQP4HjRcuv67RzVMGxj1i
v77FrcBpuTWeMfEn6k/1rLbCtTDj03gi7BV85niF0L7Z2xhCNReYCiiPZQooosy8Sm6DtcCbiXYg
0kRTAm1jymVIb+u8vmsyI8eTHSR++iZjfFGQf+pZe+pynMu3y8WoG0W4h7LqwnuF3C3miq32fr1k
LLsBhieMRgZrLK9evqYiZUv0NerLxPnr08Hn4t7dDkPxcUbkTkHXObeLc4rm8EZi8IJTxlnoylmJ
XAbijxdwbM1PfmwSGVfOan9pDtSIUdkUdQ9CyJrvCevf58AgJSo0cOzQScIPux9YVwkW4ZHiIu+B
P9YqQhGiMriCoQ1APTwRYU2Dv4mQ/Nt3eVu8iCiycLIy7pClJf+jV1aNWpvdOFlCm3LnriYxTXgQ
j9kOxiMfYNmZkaZbqKWvYko2gYWOhnqSsoeulbyOJK2Zz9vAKNRtu/j0Z+rdlnSdrpMQkJPOpvvr
O6vuLI42wmxoRQkPxK14JX5wMivr+OoQOFteGn4Ukz553b6KHWX4ZUHD/HFszC5Sp3hDL2C4ipE3
Q7zf8/UMWGm3O5AOrVe7y/rkC9f4mxm/m7udA3z7Pt9HFwIzANkKPJTFE+CFSDNBmTCLhEAzMhap
Gve0Koh8XPSW7ZpOupUbGcfcddVu2FtqNmcY5geGJ6SUWqWqXdZJTXkjALV9zQCL2xzKDmdL4Gf2
ppXitXztXqF9roqraIYQnfM3nW4sMz6obhZE41iMcmsvJficnXM4bDVlQiIG/G5MnIV7sv0g9WbT
nlymqb0w1yAQ828li+fhLcQUiFTXfZFTCbg20XOK7Juwj9k5B+ZKJKvcOsW5w6KC44M7cO/T1RgZ
xUCW3h+8Ai3DppiRIvyMilrR6BgR4mXRXnXq0IydPOeC4AQANEqvg9tf6XKBYyqgEJ+X5f28Bu80
T75ByMA6Jhlv7E9ZLDxBk8itB+e1wN4HfcFGq5TgM2aKUQplZuPotHh3FCpOOImXFCaemECRtRVl
S8i8f1rG9qZMKnuelYzCw9B5t3lKoysijWvNZMs+Pn2brGnT+zn+LSTm2UKW7Xv6T6K/Vai/61su
8hqsa8WJ95asAZBzjQjCx2pvyo7ZwnmZ86vf78rm9o8QHeSMM3o2NOTbZmEliWmMTClSdKk35qqd
zupCJdohn7sGR3+Qbsuh/U1kqGAu6K188PeuCwRwmFcl0x3tiR3+5AdHgJHM0OpyufwCbBG8IQzW
+s00++NSzbC8He0JvEsoFwqDX+JkHh69oqa2bMZ8g5+bBK/P2X6KZgIhm3F/3nf+p2LBz9yHBgJI
Fw5EU/NoeobWMo8Xik5u/VvqTapNld2WfCGYPkJIr5uBNFww1jKXK7HnZFU5XfhjwUo6bsSCtzdp
MwoenuDvepJGNj3Fcxnhnj+LIWNaFLCLfZKnaeFSs29k1v1PsOS6TSBCCwSeSb1FJAq6U9UAVLTH
vm1tmmexJVyfoeH8IhfCHzIP/nAvTSwqyP4E2q0Li1F4poZvrprxGc8hLOkkaptD+EwRAFp37KTM
NE0HTOR14B5bAEXOjq/cTqgLKT7473W2NqSyLs5iadHL+9Ta7T4y+zjCJWUVvBAOVQW8dFAFWmnV
jWeohZ3p3fzYosgE+N3QkRV5uIxoNbQ8HWOA9unEofi1EEBDibXkUZlnwIVlQnML4AskJPJSqsya
1DvaYXT91L0vBmqBKpHFKj+frw8CcfUbpytjrXIn5TaHsSjEIRGuxfSFF9YIOWc9mpHftUDINBDe
0r3WLNcCoo/0wK0y8YftTOcTwIuyuycHALxT3Dwh2512OI/zEli2ZBMMAohl/+gQotaLcaPJQUbi
sWG5FeIPbtoEpqk/PcSJ0S+VFcyEUSIlWU5hHQHDwfWMBoFU3bDCWOLTvBcp05TJlpoWQ9WGY+Wf
D/eIw9gYavFwZYI8fS5po6knGqJkEYYCl/rUPY8QnNvUL8HT2xh2Ze5KNH3qmHAXEqJrDB/we9kV
ln9QwCpEE1GKwn7U3TJ/HdNXomzbftHdFHMIOv4Fu2jFAef49bczFb1+hmQIsB1z90as9OczIc7u
0SaehnJCzrf2wauZaWOCmR1cfTBlXfEVHhc1KSrkTTUK//W+js6kybbNQkMDX61lm9tNtftDOC0d
6JHLrtSgHwl4Suo948ZJMi2iGgwGwKiFbjJXN7GHrYlazfECRjH24UjOItR12aKJUh0vEEFI6Par
AbJcS2CB/Y4QdwQhyp+0zwNZvRfTg63GmQ/l0P5ktS693eVcz31HTzqKxoK9vnjwFlv0JxsCEha2
Lb0rsNFZMyAompWsiNjYNxqwlB/f2pBbcYPlTbJXnaFcoIZZ8xSfYQPRcaOizFy0Zbs7POXvg3Hq
TROcyDnCgsJxiL3VOicm65vZcUcV9g4ZpZtCfCVUsDilnwQarZVCkuSCSIK1OdsjfULgfq93yeZC
QzsTRA/w+Enj0fwOQFSK1/RRvCd6/vufCp3WRzZs3W7X70tkFPAANyxLo4ZXjVgUEq0rFuL22/ef
yOabETZDQ6Lqdl+ilmcxBSBbNodfFaKCZohFqmL0hfzVbvhcyBTkuE22mjNgR01WEPlw1zQ0h07l
N09AGrOWqigYP648HShJ1a9iZrCMXNLPANQISLHoDSZXRhEyJ0N88o/ipwqWisiEO4nbC0/Lyvz1
wE1IxN9np+hLTFW86NY6QGGeZ7mAUCc7Rb7NkaKOoVr7VfSFXpVPsTQF/9sTg3sKZceshlh1eMGL
wIAGCnZZH7+DkMLY7KZvIcxz2SN6cu5uE0cGdG7ARsO89VXSTWMP5Ko8vsuof2XpoeFSYLIa2aUP
8tKXhwaLcu9IEldRbYpUz2paoXY35tl3kZWR+jchE561yXtD1j6PY8Forc2ipYOmp02SmMQkUb4O
a1iR/RhpGSLg3v7k9202CfR8CJktyi4hjIt5vGDxCdk4EnbPZjVxOySZL8zi+7fDpBzls+0lxcDk
s0TuHyHSb76xO8n/O4i03KRXmAElByozG2E02Ud2c6UfGjpvLDEAs3nwgpze4xUzV8ZuyS5vkUtP
+1BsHyLfO165mynwQws4IrqujLFkhTW5SNjldFS1SCPfpFP14OSseacOZ4zIedQ2Ymo5KDM2jm3S
fr5C7zYrIG8EFRonRZfAB9lEF94LrAz/z0+SBlwJwFVr8vdNUJ07/P29blqVZlDZvMzBu0kGxXLd
KlTEknCTNCaNh2RDgbLfDsw87a2pKqhPY2dRij4oPxWzHy0nJ5uFmkxwh8/uhJwEF2qMtwasaY80
PaqNy8kBXzp0nghuy2ITwOlelIMYicqfMFU2hD6CFy/ZxpZzjAPN3m03R7TG0VP7dtb2FoRRnSwg
afVHhPjd4+QYgI5PseiuyWIaOwywcCGdq+s6rwXIYXv5zQv0vwrnB4uC0BAgQgqbMuN3aACb1637
N4ES0jng+T64alTDDO1hzszZSRJU1hzZdpV/cd0Ie7I+b3lw08RvduBuiCdueI6I/B/S1u20hqFl
5XPSi1/hNu2EsNfgIRDpljwrzampAtymajk/WBkb5b/eRK8CtqZTWZN894M7jo9IHlOZkBnVfHAW
izgdBcpgxknaViIL4qPa2HfS7ZWc/iiuL+M65qlrgV9jfnkT2PoWHLXlxHXQ1XvZ0He09H2OG86i
TvjN6+htcD+tFkxSi5a0Slcgo9IFAvcWadUl4OgpFgO28QGf1F6poPPZRAj8PfsWf4UgJTJJVayw
W1x2l9gkqoJS038cLA+YsRA7fSNPb/yrJYHTDDoMG/D2QmB92OydcZRzU6S5b06jGD9ax4Y3VXEQ
2xNJ75+uxjuRy19gSr81nIAyLFQ9hYMpE+5v3X6lDouJRLlJR28PtSnNtT+C223cz/vPU1wrEFgY
7bZWe9d0ClO+dxUR3tfk+cW3Nl4HKpdEGUvgNJlct0Q8zdCGSGgBVYZx5awjG1e+0cpZmr0IWXwQ
wEljAaWsiKEbaD+AJpCsiC/16P3MluI3A+yrF6Ohf0Sep7BQxanbDFwpThyTY6YLtUWKYHz00qp8
iiowaAxLKEP7cg1oL/rk6J3XgRuqwpjEIzOfYinZOajXnNyhs+2K9Vd5l+tlQd9L05Pl4nGQaR4o
Fz81OqMtvjEa1BTew/zlZ4OczYgzAqqx3cIPtg6+Kp6zWNAf8XVgoV0lwSrZydoLiPrp/v9olXts
uwLqqV21iYvvf1vA3JGQPQ8qTkxZijPP1Iu7QwKK2KYxjHvPNOsGW/mGyJXR3RDD7AbLxdULaI+p
0lqh/0olsv3rYAvG4mJe1ZOtrLEt3P/ycC921vGkamZ0D1p6of01yg5KiFYrZX38EY7EZIgH1ilW
iHfH5Ju9xCsDcbvEGnl/u7XM2+ZabtCBQjEmOgDAqKret/UGIM21BWvI/DU9By9pAZ2iYfuLF9z7
/+/UYUMUvcNYyKxUMXch3FWU2su5q/MMGBIavw+WeO0x21RvDHmRCnai6vhA1ghUx2W23wzYuPCf
E8EzJYPlWRp3mglk0FOdEsV/nS6UhVNguEUU0sZKXg6hI7DUHr7rD1uXWPiIfRpWdTozHgPweCkk
K/GHgbqetbUCDvTFtUZtowmX1ezG6kVEQGCTPUL5nMWupG2oQKt2CbLzMGbn3kIiB7t9q0sRaD2J
vJKeSivQC+CE1QpxQwCEVlNE4yPdsv5RfT5qPO6nmStGiLjL2TzkqUeL2wf6Cchp/lMhWst/Yz2P
DDEjJg3kjuuACNd5cB2mVlcQLlJ8Yf17AYKTtvwoLIFblPJlmZ0xwDkKBxcHGLA6DgvR3PFc2N6x
moTBJZBeQdywcQn6NBaFI7maz0e71tiZ1lObyt5WrXRBHsfakS2QCfS7kOuLWiX5f9NQ0fB9ab43
6WdVjsGeHPMFwXfmC8yZSBxW9ynKP3Tz8F/mjQiMSeAH4Nckwc1QKIuP0E3H+uY0eQGnHdL0Uef1
r168U5zWzD4IH7KhdWArOkyHC+zREM6MrK59bOpFk9CRYIUPQUQAcDA7mzFx9v4grYa/lEy/nqoM
0QSnRi0Z0ZnbFI7/u79tQe89bICavdG06j69d4yKxypaB74u0T6sPBSep7sVkwFHyzkW6iaSHXw1
3AB37YbGtUrt3q3tUmBpOX5375GpIGEejs7zv+/5vp6MXt8CJZfammTAnC9Xzg+dowC1/IDINzcB
ALqFD8Owww31FdopqS0oQD8ZLsXlBsryqoFKlfFE+8B/aHtGSAGsCRTP8cOxGaAmUZtYOo6Nr5OE
py/FXCEbxx2FLahvmvdeuA9q37pa/TcA6XpFp2poPWwWwOwp1dFxGq2FtpcSedoz5yImng2DBdKS
7adhEPq7zAyEhzH1PAfFxjtWUiI24MVhRuhAykGjbg6LLrsWCGv09oJfM0DGea3RV7FqP0hh9tpk
Z6Umg9rZJbsekLYclnWiGA/vEhD79QmUmUfqwOK+eZhoS+ACpyiN2aaHMc2FQsD6zGgFB8CXFJ5Y
++0uuawDQLtihYu0yTdrKonRiqo308Zzs+jhmkvz8iJLxVTjY62sKJITW2b4efYWfSIh98Wmca6A
4TIVxAXK0YAJ9WVHc5yhmNrDBQTDOEtEzMXWAmjLLe0OfT4d2l5d9V946EHhR5lcSLlZFSbilZ/1
UIMRFArPP3AVTCPwzxj3/W858ze5gMxnRX9yiwVA8qZZh61WIQJJe06GY5Vj+eQAsMAnpld0xgIa
evdf2AlpejohXL6919AVbJu6dk/F+tOlFBaSny/kLQJXPClogmzPHqCAGyHHkdxWgnlrLIRe6GYH
jJR3w1UzMdTZs/s1CwuLm2ZQjBeMz6TjtRVssqCX4+mkuo9nW8y+MXB6EFR2HnQMpezBHlK+aAgs
YJrUN99a4VQKH3pocabbVey9w4UlqdJzSaSL735ZlMP7BacmmxZ1k5gdOSLHxhyZ8N8W7GEhZe1x
ud/G8rjjMz2OwLGLxlM1JNjJuBsNtmADgmcvIUufif8JfDONJL2Uk4rCqTwoxrM8GmvvcE1BxJyU
ebZ6lGQBHH8tY41dSEV6F3bf4i88aMfAfsyHXH+sNJzR4KSHbtkOUk3lWInjeAx1BVvulV8PmAb6
RDXi4vf4257t6DSRunDonDXlVgMGFKuEh8YeObqH+wZlaSOg8uqGpTDiTKNFT9zUO8rQ4tfLmDPf
1Gn64uxBWhHlTnqlE6/a0ncJryAsN00jsbq4Z1MTRCaCRrm7HAqLgvz/cZbR0Z4tGLqDhb2HT2NO
GlMmXKbVndoahn12HegyiJeB/gijCtw1PJJEMyxDWJuj4gl05/sNLKd6EuQJwhRCHkSSm5rm82Uu
pLizmwB+APqQv/pzaMr6O7IPQr1osHlz9ZCounDBoaPpq4PL5ps7ZmdCw/fkIvvW/z7IGcMHjrol
E3xby8i/rfzaWuQBiZZm0vGAfllm5oo+AMoMlhXvtvdfsKWwUQWEL8huoWLUBgII4OW7P1txgljO
ShEYsfgthT1TIcChbW7fr8cN0bVMpIgfoVT4HgmSuq1aAp1o93k+PgPn5w1fG7cK1226k62JOHgH
ExGlRAYhb32J1wqH2NBMHrPthlytEBhLRxzELp9iAv4S3jpV3tjY3yoWcwUXKDQ0/SvC3yN9w+0c
PVF/MadF08MD0Y81x2T8QfkWLY25zgN7Y5tpRwIwCVUDNkBMB5a1WCoT6tc9TJZc6pHmK+KyCtE2
i/1lcZIhTk9SZrOA85xcFtzybOGhz2oVa9fp+N+q/idFag6NVjX3iZmkm1ThZRcQx/l7g+L2gg1Y
3CDK3zNWI+w8lk3s5aG3chqv8qxq9pj7HoI8vzq6Sf6IHrusQVtVN2IXJXu08mtXFNDwPQ3euH2S
1wPK7slnVKNFb5+6gSKB/TnFzMS33R+zFxLYY7Aqxn/xiKmNNJs+oq+tMKQeC4eJUGHce+LfQk5G
kk/vskuq3fnifBGUT5mZio/rE7givYzGb6Xbz1HPKIY8nC5aa27uBpZpQhHa18Z2aOTjEhZWzXOi
JXA0gP/6rqVBE2RNw2Gf4yVUP3395NP2itU5iIvHMrF7tk2W8HTV+IRLtX2G5JNpsFlrnEJJfABp
O09TuYrXzdWau27mpg/Cl3gtYu1JEUkdUJTXuA/GYSfZOJeG4GDuJIWeIvp/dAYwv4IejWYidm0T
ZRF9XbisVsfwPqSJtEI/sYo39TM+NDffQ+41mKWU83m4XrMH4K7fovX0r/TluZ9bYD/H7mLFKh/t
7gZv5abFn7Y7VMqWRuiVT91vjjy9ZvKAkRY5QTJlrSIhggd27q6UfQPY34VDSrEzH8DZlQP0rgml
spcUtBesl4S2Ks7Y7GiY//MbXjDh00TCtKdnNEfJjHSM8B/Mm/H5xvSCiLY9rkYGiExPhr/dumq3
UcZgwOApZcn9KpaYtgSNLRkXGZCUI8scFZuJ3JgCuvEOOf9NoBh91Y9+dTuZ1oDWhyCECtvFiYvX
+C26rupM8vzAybbODj6E/0nIUX+ot88IzccN9f2eJ7irlxFqVlZFXC4Hu1zcGKEnEDYYAVo8Q8KD
TWlwF4iWzLHxW2VuVZyiIlucvk+wcmB4SfD8vdaOsS3u7GQOHE/XVKbfoD/HVx4otQvYUso7ansr
V3pOHS/6Ob5gWIXIPLJSjcVwhqfFW++dAvVtTj919lh1eOBfTlJ8T8iaWP7kSMj7DPz7d/e8XJbj
bbDJNQ0OFqG5gjd1NMpuw2FnSNNK32RL6SqqXDOFt/A2nBplKwNaZJcwGJofx0R26NuQN2uTyE+O
Rv+2whFP76txhrcSZHKsgNY5dha137vbvjRWtS7/A/ide1hhLry5XQoCVlEOGNna9pOz5vmwucTX
HNCeGIyAJKslSnwok16DSHj6RhRrfwCQnwTo4AhCtv7ChzehCHg05XeAmIOh4jU3wsl7rMyigrRK
z5piiNx9iSCroOZ5c6aKuL5pvm4rzi6Oqsj8H7NGe1uhxU5SajOumTVogsFnwAOXYIU4Yg6lj0sL
+M+H9/YBucXkeCsiiknoVbl6q78stDh6ZH/aDc/JFXdGklfsiO+QKBoHwdMnLyocv0UkFfmcFKIt
RJcnjyW5LgtnliTrdceVZYp65gWvmJkLbp1cyB927WYaYJABGCTh0B0ZggugaKFq3aj36rKd3/0W
0wzS18Y9dENRU/y7y7gqai0ZumN8Zg9pwoWV79epN5wkYgyQaG0KMtHBjusnhvek+McD3it3NW0f
IIPCOtbIs0/cq2eIyivDVJRLv8YfTU2fy3DGE4nPpZPSRhfUbC4d5Rgcgr+sM/Zai8HreZAL56s1
AlyDuZMrgWpqero5UEnGCSpDnHaAekuvw08HPOlCdBhUloUoO3taXYZYJ43yFKPPEEarP3BNQBRd
8lo7NEDZQfVmH2XHjznfphpVSP6K9/Kii9IA7PQ9pTGWiqN+5OuElE0nX0/gJqgKPhjxvK1sAUVL
q66fU5SXVjb51S57s5gr7Ak1ymGNhxYf5YLTLUsqBgHiEm2ivypR1frOTYMy4O1HErKx2S96mVm9
Ad8pmh7itFoH5aFOJK0BoJLixKSSlGtQ2ii8RwDL09Cysk6UGBsCze69qZue9EnlJtL1qhRKkURp
6dzzdNClqddfP0Z8RqtMy/a0dICp6Bt80PKrJh1rxb4fqfkd+BOSbL8vZVsFWt0QLoSMMuh/8dfW
HNs+lkr0708LOSot8IWmt71HoJbSf7Nqw/Xv5Wnq1HUanBna9kVMamQW5WHpflnmoEa+Bkb+nYFU
vT4jfluPmIyn+EjtGhoC/vCwMqEt1JOfuFf+DVJ83SNWaAwiAwv4mRxNL/Uo4wnQ6o6Ic9L1KEXB
SnOBo0m6AhvhBXke0b9L+wFQ0/yDy4eKsjAcCUcmn1ASXo7Wyumbm8+opPbq3Jfy+GSBOkZm8OIm
H76dWEhm7loqreCZaLNJjKtL2dwJXGgNuLJEUxbomCMOdbdQbeVHxrrMpBmfuINMiCzbotzMqdfA
d6ohufOf7QV6OlwfibcUxkzf9bHr1cThCVNuBjaJKxCyKbvAqcBiNODaZD5TXQmoQpcb71j/TbJ7
Lq8wpd3pPNaRuOU3HT6TGaZtQOn3faYMEE4JeIzoNbR3CEXVlsXtRDJr6FzqNWRvqwC4lXlwMzcM
NZ12TJ2Pq5i73+pXCR17QZSsb41IGNMLhHxFDABWqEtxn3FUQL3l9Y09tgeT5/apYZoGYvlYAZPk
KtrDzp6zq0ADuYZ8RBFms8uJkkZeTU7YbXt0pLZkMe0esCRIAEgfSD9h5sc3Lwy5bH0AzWiMdlsC
9hotDxPoQzsoykql0H1t7IP3PdYoT78leETjshj5re/TjeABT1O2PmyL/steJ2i3OKDkCI0wi6rI
7dZiYkG7kNY2wlbeaZWzDJtdpxwziV5080xyKFe7RMqNfXI4/mFkFFwNt25oV/QPfzOXIDnf6lZK
Kzh2ng2335BBr/cZJTgALIp8huijMKBXgIMfxC7twyYvra1v/rFsHvi6y/eJ2hUaQkZoIw5IMV78
aVWsBJUto2A7SoqdzD5Shed4I08eslCQvfvj8ugu7YfO5qpSYFUDjlf18N1OGmm+4KhPVbLeRSHD
Ny7xYpDO8HUgQZkwKXQDBplqbvNcxExNSg3dZxpTfd6xI88we2Cf8y1Xd75umsoqFMVbz3BeoQzj
dQia2FxknUF/Xe893gGBZKr7fm16d25PQcCOXLo5X5vHt0jblg5p2k5XRTvczjnMnm0c1Lk5kBA1
v/WzS8CFoGmC5ab0YZ7VoGQWP6tRERi5vtuU4E0d9AFsJ/0Ef9uHxUKzDT1O7SdWd55ouoKDd5f8
m7R9OY8+P0t4Gk4vAFIL8bgOlu8E001vmxz8ne4Ddw/4Ubq4tvq6/AVF1qSxKYUghhNG6YxZ3v1B
dfBJOCT/bmFBOGwSrsgA0t9BQvHcIFE1GLWtBie1lt7TXeDSYReF7AIr3vX1L9AtVfHWW5RxiOfx
JdWpwgf6oiKwTRlZdRpceSDlnlKXEwwpsiR6kFaTns7sOJZjqlS+yDAZVk++7vbRKrtoyRQVLLIE
bfdJKujRtNxOj1zle7vRRlKpnHgxM//zQfBK8aTcLkMndugY+YLSUXTpwY1ndfpV/ghURwXmry0P
sRjzmFE3mEdEorFtqPnM1BxQ7dBopwrRHzBO+aNWcJqR/C1+EUH4dzCOIK+XRpXtZth8C5iGmVIi
La83ACiU19XdQxDsj9a/pgEh6ps2uuPcMnDoo4cHQJhWYSem2aPWSeXxttW/JJi7jkYjxTgVr7xB
axrZkt28FsPWsrk2BM7Rq6uC7jCBGp4BrW3hm0ClDzcqXP6SzY8nfeGRB4y4n/3nJdkvmH8aSc3t
7bLcCZ0jZ4WY600TuGUoA+dqPzObjaxyJx84MicdANybmP9uK1Jbe8GKuTWEaKbpqSEp6+J9hBfz
iKNoZ7jOUAT/GrlcLgjbSHIJKyUg9a4qe1R+E0HCXGLADeV92wjTw4OCSns3XINeAmzDZHyQWEQR
bij1kPqNnvG0zQiai6ZQLtpZVMvbXjcBPIqN4JsTPpUIt4xtw2EXbcAOGz8ztjfRdB1nqS4f1LnB
GIxqaxgRUqzW71B9jriND/37UmsbMrfpwkXK4SvVuGVGYT79fRs0NSVQlIU/iXZZcugVgP90AxkB
jlj2LqCyFWMmwNYAKC9PNVX8khrZcgZ37DkM4WHyBbZH0s1NJY+WMg5o/aOnoDdWFvQc0OtlED7f
RUbMFWXKZHmqq3qt2wPcUQucV4LwcaETiimkXTNqJoI/NlbVp1dVN/Y0k5bGrriscocc7lG4+9y4
xihcS8nGMKJMrIKfkoUtN/1W0a7j2u7AJKpkzqBNULMMeVVddG+d8tYs1ZwUaZvB+wQ1C1N6duXL
k7xelTQxlxPgZXIi3hxVu0YCdtFTW94xoULCxNjIGa+0KoQf/wl4fxQtg6SJR6t1BfhTqD18vLI3
G5o1UdoT38Nf1Dg76cGRkzPldaGN5hjUGGbLAiDApBQhVYo5cCB8rXxHgeMrsrdVmYVeaWGZO/GG
IjcoCwWav2m6cd8e3VkRbyeYKO8grpWXCCHlxeaJrhISW+ow7XwbuvwDAiAeb5VNqEYM/mncVIHI
650Y/jqV0J1p5IFc57GfuB+lYObs86oJlAnAsg7ij9+wsiMJb6WDns/zQGA/DcTGBYicxiWWH8Hz
aAOKRSVQuD8+sqK6YF/MeZwtwGJ7sOw5Q/qlc53l3yp8kl7knjso7y7Vfe8q4mJMpn4dzaDcdisy
dGJQYb4L2U467WrKD4Pa4lh5f5WbJmBmDcjIQti6eC6aMIGc+Km64b++hxOcB8IxX3XGdRaJJSU8
vowv84q1ILRQrt6BoVVfezrRmmUIOM7UVd81w0OUiyPbz0Zh/9eWW+Nca5TUf2b6PIZiEztO86wV
/iFHqHH9x6kqb4G2hALW8XOaiJI7ZthaL0LdrEPH6XWS3QeItHi/KDqKvwbtAsyGZKL8ntZcUAgA
5Dr8xuWfLk96se66s180ZVsGbgoQLw+89EwOG9eRv4edkJh1ixfAAU58YI+QmUdfJbTOt6tuoLG/
J7c6aad53HN1ai8aCyKXZDQb2jOz/egz8AiFVFOpcNYL7+HHl8Y8Rzsa/OTu6qsoVILG2MasIPa3
xQw1L8RDIWl8PCSEp7x6aZPPPETFOWt1hqf87DpOiXnUwQprZvNvE5UP8MF9wQPJhl2+sXSPypl2
iqPfNq0R4QJtGuakkL4gG/8PS161KUT1uGneXt9DLHvVEzpuxTr5pinPHKS3VZC8U0ss7UAUkaKY
Bw0ySnhkiX38ah2JQJuI25C1fobb2EkD9Wh/cR956MXgnhqElgGR7jT6Rgm9qhgcmrGVb1E1Udqn
cvunrDf5tmQUkpu8vo9lXvr76g4pPmXKT4pUTBsH1l7y92/MPIH+JA1zblyR1c2Zdr8hNrppmVX4
f1evvl0a85An2OhJxiRtvCMBpq7iEudWeWQPl2aDrvxccVfbaxarK/e0obZVNYPZ/uHE6EPgjVpB
DcCB80OjKsVvOyrrhujyfj3zdna5IUJMhjC2S8iIge5h0o7l8mvWRuMcJWzJH2v/J9iJ0kj2tq9x
5z8MY62Gcedsg4+CPbCkJKaEoEzpqVorKgIyrQWHkexFpkLKJOuF5mjNgl+qYCYjKfp2C+F7a0Bo
oNsT5lUPayV6Ma7eY5sSBFdJG/5kbalMTZm03qr8pHVBsohGRebTZfA7jFFBk1xkVL1n1bF15Bir
geypW18RYUQV5BE+fcIVG1qQvqQd8S084j71I76DAdBMp99iaSOvYS6l71pZ/QoxKwWlmgXqCpGA
jvj09u9iucLZ8TFdd2AyqfS5gwtXY8Am5gi/em1ly1+qxtKEFBsf2vzc7mZbZCgdiw99UtdqP+sD
P2a5zHbPFFaLyZN98v8+24kjANB9LkMtGJbLWwVkCBJ13ETUoFDqUmmfMhCli7RqX0wipMWAh9el
9uKFOcMtDYp0u9KESnmT80ytbmoDahr43F7pW9Z/u3eaX3WdS7n1UvgVrxZtaD5v7jmzUYutD+CX
x91nXXaQyIN2UxbvD6SsRpMJW72MwvDQ9pFHnaFKIzQw1vhNQ0/9dGWrS5EgKYPTocldsF9zp9pT
jdQ5RFzq6JX4b7cHPfSbezU0r3ycM+Wr9slIWBCI1H5cJMWfHVnDLmEL/WGBhFAHsUm8+EE4XkfF
5Um7wfZx/3ZlOjJ8ZGM3fP5UfHwZigNlC7l7NhdFsi3uFOe7aguzLlIhB+BM5uo+o0K5UwuHWhyw
jDcPdQnUHUZybfxHD3llNxupLnmoGiMS/49ZVetyeddA/qsx1ZBEhWba/flgH11+xW7Rtcyv4p73
m42iTSES/jB5gV9AzG9QnlLm05MgVXzHiHezpsuXbXYc/J1++IUxeAqgoXah7gjITAGJSjlXdy/3
j2GhRw0ahaGuawId9ULKv9zeRL0joeuHYmgZOPmsJrBlieXqkk7nPINHsXhyGO8hBiHF/X+H14wF
XbClE1QOe/90FaH2n/fnLO1MYK1Gfi2hfkMDtrLTToEXoKiTDIc8NCM0caSPSv9BsDLdtHme9JMi
kNg3TJk6Ky7r4kMhVROfoBqfkEReqcY381+JbiyUSWfY+MOdMCDUqledv58uF7m59LSglUvyJecc
3tVy0fIRwCaED3Suaw4hLaEu0FCdwEB64+hvRSk92OA3pMAtN7apt06oGD7Ldve6TtLnLCA8p3UT
DVlkp5/wgxG5mjHiHxQYc8shQaFs68EIgI1OqwohUnPt9jAoycAgRlR38W34E76gWaJjmXr4p2CD
G5q87JXGkJMnPAHziGwKVoP/xT55Mtn6P7xLLaZ0aBpkyHJW+DlN0K+38SEHELkra7rMziMYBRRE
yoE+AuZkBRkcScxHy8GOBltGmEYlZr5YTyl+3hKXCsP+bJRznEoDyTaE1OGXCwEPKqswg1YvXK/u
IH6l14JM3BcLoMjSUEAOmoO3egiZoNwDeVlmbUKTHO3W8+aUn2NzZmKyxzkmVG5tAakdZdD/tJf6
CvTCuDA7Z2ksSKwIE/HJrWm9BsZC3LjK0MA1LX7oyEOXZNCP9TweWYNat3lPLwi/dI78Ji5bv4x/
o0d0XyXChvquAjbs6VfAEe6iDE3euhqADkTw2ac4pGwoCTsL0xFpOX/YU4bHgqrO4NhWhqWhCgUl
jc1231RpPu2mZeLrI9c7bAzI2h0JpFWhlWXApYnw1SW5iM4e0BwfwHAKBN4I9Ti5wXOcL1nDgwx6
vo4wXNsRpcWZ8AoLGptK66mONFrcwbxZQ/MJxda5SeKnNOxjLoS6gCZQuHG2EiJgo1co/VMaJF4U
t1ajoxpQ4ilOCNId+lMMH/9NLmboDnf3pfdpIjqafIV0y4Yx2Xdqk3aOHmjYB8LVLp2Q8YNoOhxg
9Qn15DUAY/IjLozaKdMEJ/0TdltD4CQJVGkqgwlE5aqMROqRyJ5GgYMtpYCRVoC7bvoD1JzpipEs
MGFwwmNuIvkIzS19pJFZZhqyJJTC5F8o20SHf4z14+zRaEQSjcX+asvK69j96nTUKY9InZUGgz+T
TomlswkLxwm/EQbOM/ImtoU7BzeyIeo7NbJiBY6cEmJtDzvm2xquYIUBRWUaHRAYWPUQFp7sPOuT
7GSBA6boAfiFoTkYX+UI+eOD2JfSKmj3oKhPzgM9F5ApFdgmM1OfPG1jD+XMa41K+gHewesUzXSI
ZMeNKJu/ZZtQ4qpeJ/EJtEURL7UWD5Y1RZySDIWxVcz39t2PJTXfGyNlibBljkySfLOe2gSYnIvb
DJOlDe4sswmkXdCMM6N7S/mBpwDAwiQ3ynsbXgcwr7Pbdw++Bfct4bislKMw/CIKjnQ/Tiu3nDk3
ISJdu33jM5EwHcD5C9WTFZ+DpI3oVU06fWEia60w8ItSSjpqxFdgIIynyrVGK8RPaifwTYKS34yO
MmAMCiXkNmiKGny0ftsl0XKgibW4heQz9DhveitNAMgy8K04a3uzEsq2Y4CDEWaO5CgEDjSE3eKM
wqikeNZiCd8VT8eTWU9IR60a8rGchtDRYWBkyOdAR2TXD1T/bOobrm1IWLF/cRI9oos+B4XVMLt+
1kMZYQLeix34rD6wTjyVFt+7NBI81FuRrlqMmeXVmyMbdGeK1MOKmanVLA/nX/Q4wgFbf+8p4W37
gCzpDRlXlZERDfcQhz1nhEQg4TpJeuxhMhXl74ynRFbcDJcRsPkA4C6XSQycrOOwsHAbauSQ/6Ob
d/f9jVQtNEr652Pg9IM4C0jKW7lXy2CRxpkPePWfdkieKSbumBBKWamLA/KNmfv1zPLJiB6AxKnJ
YfeU8ScEvGM7hf3qHcGofUrPeD0m3xkLMHZu0u51MrqQZ05FSMtjDtiDBSJT5FEO/BGRsK0S7Pmd
gDG//2Gf5DeguoXjX7gzP+VnGzOHptDYOeucQ4yO5rQImw/gPPxeh6OOcAf0zmQOcUI5HXdW1jtp
y1sViDbNQWH7FKAjkxxafrY/6Dgx8f/fybWkD6boCzo1BJKuwiGOduraKtjEoU5IA8nheCJNQIuZ
u9lAKu7IT5HdYFLLi/HMVO31ubAO8+mMVbgFnta8UFAZ2zWkCnNAZh5dHep0n+cfR6Ue/K1Wj8QH
Hub5M2afpK1J5CY5m+3cfC0yDsmWTpXW+DjENSsTy7QCTTz13LXdMOSp6bJALuB2oD/bjUpwhUNG
LEXpB0Vi07tnoPbRbxvRxCkF04cDGb3MU0OUZT2sB8nK1XtyLKPj0eBRuqhgrSWnDNM68YU9PmM4
ra1GXxZAMeUUpXcKLO48x6hXYXqYqsnMDGA0yEGdzccANm4fM+sA9+663sby5n+NrlqQHvyS0n8e
Hz7pe7TOryZEGfQ27PUIuxHydeH4W6qGJMXGNqHMRgyjZSDPPTBGBrdNADaDKIcj9oZ01njc0gbk
Js2d3iL2eIG8i10Hwhj0CHITqQ1Ojreq/mCmxgI4PBYsI+Umn+pXncFwiYLhcnooQlAccSa05Oq9
ZzmDlnhMfQBuFqGSqJphg4Vo14QVo7CEcHorRowj6gjCHhjQJeV83hCc+BINAJ3zVJV6sPApD+Fk
yZ1xVzM+UGxn1Y7MppO1w/McbjwyLuFMwEkhGcSpi6TzKCBPOs+AUkjOHkl59J5n4BPjJBgJOQAg
OU78+1ZPb8LQfT3vKDRAG9ezAVcuaSTMEZR8+I2nAhZ7XC90HrXhM6C76jmRZzhStWk9eIZiCXo+
3oX3JQrptHYyq3atv8g=
`protect end_protected
