`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
SZa+pTIQshybUXK0L6tPoH4Qj51upt9OZvviC09Y3+WQ4+syLFpVrjv6Oym7ZorEP59RKXms5DMy
HXq/UoR4HLfzhT+8MXcxJntSaQrvdeBl04vSmITSmX4aT9Zqzl4F5wwl11EnQ4TTMADR9nt3cj9L
NP7IuzzzAkSd+ijeNWPM01UXfoudDcRmNr5f9khcMwpBdOCA0iqyqujwxSlPzu9cJIzgSWAPhvDl
sO56flKNnq5TJ9F76JeDmg4n6tEoDn7QrjkV5r5nwCjdzL4Nmx9k1XbCEMerDpJKBXcl8CUG5weu
DTtLiKQiSlCogT003kp/KZupItDUxzZ6gdczbw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="9qAoyWhr61ehcOOrPH1ic8ll1rCtC/Loq63kRSP/fDs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11296)
`protect data_block
p9BTtFoVlk5xvPYdhXCjZbfTOD041EA7zcrimr2jVOW/bLvgtKh7iaD0DMtQSj01wzV9JlKsgwYA
Br66BCAqQays14Jdl7B75s/3a/TPbZnABv4P31z8x9NkSyUKzb1ecx2XYUkZIksN1ipV+acsQJj5
Da7WOlr5zau/5VAeoe4N37J/HJJtCL2L2QuNRFfV9NG1FbSCjV35wTnC+vVkF0SGcUJW2xwUDUq8
cEXcmQGastpCutlAPxmnEp054KFsK+LlV9OzOED462U46rhlYNxEBPhlFnEOnJSIIjBCyHjl21se
5kZNrljtc0NJ6hKZNLKEUJlCo4E2oQ0LyvbebfdOqb93PaZpHa52geZZJEQxZEpeqjJDpVS3hR8j
8sXzK6B5GXiDXz9WnLzU46CBAkC814rGJ7HpNKHW8rhNO4XoG6bdn46bpp7Jj3RkcLisjFiPcu1b
RkVpG5s+hPpXTksASML2EGp/Ld346JLIau/gUE6PfDCWBxzO3nPxluRllS7XD+7wCBuqd5QTliAM
arsBfSC0dz/CQ9htbdFtjdB+6kUK3vLvQElhhM30yKh5qYXI5BUerX2KyVWkewacE8vE0XHn85zY
S+73aJhhYdWhxo4KCCZUfGYGPNLmXt5X748UeumB7jgdoMiXPPIg2X6RK+TZrWamdxJkUIHqiL0N
U+yOrU7cG1v5X8TxdMrV6YxXSIbXj0sNtHFhVYg5RIH/01K0ZGGUtNWMEWhhY9l4hOGngNOt8vL2
1kaWobRDuOSuErxe5Ta+b2HFwtzuqKEv1S4UhWbOz11u8wjrDLgcBiMRdbpt0Tvz1n+s7qqfWsdq
WRNvzM3i9tw8zCuS8xj4d4Z+8KuFRnO63AGINR/e2zAObAwmPeU4A2T162KfVWtdK6WuewqVnBxA
lD5PQzTmtVUvI1GLNYL8F1aBWqSc3CuUiJUUoB0JjfbliPaGsSm0izWiiqStSXuek9xhK7UBQ8Cp
bl2uylUYV49WZ/UNpZn3AZ3saErxjeBHIE3LtCiNhJyQuzljYXX5xZwWieKzCrWxBEDtRqqIJOHb
001OSkAEXkClHEGWAXcQv7jKYQ016Z/ojeFE+8LbzkvCv9+xd9SLTdwfyms9usZM1yQlq4DOyKcB
IdEF04c5C7c1GzFtkW0Ht2V2nyuf+fYqND7sYcrPFanRfxyTwnyfgtii9ur/UDK41DNkw5oeiubt
KlUTGEFWKnbEAGAOyrSmG2CMoky28vo6S2Mpypf1Dw8IIvUpcGlzsajc/GYvzERm4sMQKFGIkzWr
Be5VPmYMYC+0seUGNkWTkcfaJStGRThxkauKGnZqQ1yNqGcm99cP6qpP+0wDKfkiT1Kr+6JzRUXK
o1c4b167HGRGb4+xsnAeglQMHIhmnjEB/4fF303zFc5dqTqVlHD3Cdj5rus5dPeNMXscUvNub89T
VOOIW4OHvKQlGpi5iANUA1aB3oyMs4QuFOr4S+udgMw8CX+7fYL+1VanyTlyQdJRF6PS44rtqvxB
Pxw47U3hYFpXgDwVo9abko7FFU2glwCjte1FVCEcznsg5lI7wGAiclzo0fJ6lglrX6/68Z5d3nOL
CNyVwJv+56WduxOPOMi54Xo4kCKOxpbEz0MtunfEFlXARiDGCX3cVexd/LGB8mwY+44KdLHePq37
MOMfpkySV5PCRk4ijuGgjMZ887gaB1ug7KYxzWtKbiDl/pVQR1j1qRO1Gd8rACLfDQCrjPAhimKx
rwGOFG4LihnBAPnk8Hs9LxNbWvYvKJpK4VW+ryKTQFt83/rdcNGjj6Oh8EX0nDQSFFtIhiyVkBMK
OzMa6cgnJaPtUdCg+N2HF4cGLIpTUDMEkEIa8ceKbTK2ggNipNgQSMl0iPHEZeA/EctFhENzgsnK
XqjEcxJ9mRh4cSjFJ6Nvle+qrkMFTkrd3jESYcZBYxFxjTG907hcY0BSxxVieOsP96MLonbWylhw
1v45NmQRvwxvGOvrtob85cT+hNn2UQ0Q7jJVxBXEHz+LBUpL7wgb1N9IG+CVBmUG6OHenN6FXq0a
KGWp0uFQOfCDqSd+G73GId6JCqn5ddruNJpohgM70j9B9OgoHR35BU014VengwsOP8R0QxNXlw1Z
qYpp1n7BlQ5sTnbi1WN+N1VzHqzCwQj8+9LGa9JRI0UemdoCiTHXjqifGN8G29Yph21fn9wIeqbb
GUNGpXHu3CaAPHc1BDbG9t3tkvmgP/QdUSsIci0ab/hXO2uSUtT6iIlG8ZFFmN5aH3sDyLq8fqsi
PVJL8wx7xZGpSnfCVQX+FwxZBvBwMooSpNoLU5UuFMOVuUGmsfycdL0UFvaSJvTJdUEgOGrOmPrC
Np4dv9iGveN18lm+rzksNEy1BQVeItP1nkg4qf5J+EFWyVCjlCf1W9dE8/D2mce4EpeXd9J5EFLn
gN8jlG62ML8mJCohkFvIu8T3sZ2/51sKVdU/T12+3RStvm5Z8lNCQlFkUSoLgB1+emfymgwylgpl
yxI0C/FL+hbxAjt3SU7yfc0P+GbBvDsqZChcGqtf+pDhqDZ3QfM2ZboTHFgg9CQ1r66LgajBJE0J
QjNNrkznj8wstkqm+AAmCm0Gg1xLrpg7/5LdfK4xaufTc8jwwgGZenmbp5xQjITlUOz5dic7KUSc
0sMcfK8dtmnGE5JAHdTsr9yxEV1J5+yb7MHfzSg95XcXkPBmTZ2vRMH0/yTBtbC/hahqApP+pKn0
h1vajRmb/ePuHGLtOtN+3BVFHaJ2KCT6ZRGf8EaxE+OTssuQr2RBEm2hFO9Aj7oJUySfD2vobev6
YaH7D7i8rp9zFD0gfWqPyxcYvVbB1R06Azq0gEnsnXCZTCB39h84TNHfSVwJHsxzYQWhIQw3QIw9
3k+ZmvP1ihI3vlKBa7aY/6d++R4hDmcbpXfOfFufx9g8ZiG86SsT1UYhtT4II57B3MISiFVUHXi6
gYJf6IST9jztBm8PmLzOClkE1I1hYfUtiVZADx+WWbfFgqpuHczMJiacmCdN9Y4v7qV85KeKjAxH
SSxBQxWZNRgxwnWxh/0y1YGqX5Te8GCISrfV+paMm+adiO4CZGWSa6QdxP7m8NT4+DmdVNirVybB
vU6ggabp/CGQH88AVPW9eaWOZQKvWqSMNCp3fZogBGadc3eg4rJxyBZyBTaJLoIeVCMI2bv6D25b
GiN8iOSMmaBDpW8GLr+Fi98BYb6hUp8Ki0VscBseUdZ51yqw58zQJpSZK832U4EAQm+3tKuXOuxI
dUPlGp0qaW8yZRNDPV5/qpCu/y8hCm09x0+ZyHOyKrBO697UjPfpNR8Co0PsPbsbpQfANMMh+7RI
oF+s5DcQc6Z53NWQQ5P9IbqLYh9PybZn8+MPfzHMRpwFd4HBYjeNTPaalle15IM8GlqMcvZTdaRk
hMXiaXcFP0fXWwA0qKEnQeciYy6a+CDgHEunnXWrU6TlgDQz6JREf338w9C72iVav7avdilfKRCT
8EdL0knqF+rb9Z9sLTvZuvO6VMS3qR8WbtzW1MUIz2WqdbseMfhfLhzdyWYKJ24Q62z3hQVX4nlk
8/2XcJnVFd/z+hQ+ajgx0t2OlxR073gS2aZFcEsTbuTraTs+6RjB601hDP8y0uhoZW1SdbMwZOsL
rwkm9fPbD3FXgeDOd5KUdzOEnPnALTnnCbiu+O+2dwGJeTy32SvT0yhwg5rTK8IXpsRKz10pbuHf
IvwxgNgXALtJ+Oscw8Il5wb+9octZWWCKiuLmtvXSOaGI6laozwaKghyDeaoxXLhwNdVQkshhsT/
XyV7a7ShDOUmYX+owqPVJoTP3bCZWKnNmJW9733KdsOmrLd+Ungt81jOLXMEzlFC33/IFGhJxuG9
+sRHTQMrEbMuyFxBzRu1X8zjUu5iKNswyjrmMT7BrSQqE3cCYHdSzYLeKVF6GVA4/AeoiRqbEE57
NFRxecGtCkmFuq5L8sK+nEvpgp0haj6BPKvzZM6fZE0SBEJo3IG+IIWUcdPSkgrdF1edW626XwIX
LPMJ9MxXdpzqJlnkA8C7Vr3Z1VIpJoc7XNAu4DdStRQkdb4X2YM7CvqmtidItn3o7ntp5ckj24OL
87bwglrEdsyKlhlttDviKeITICXvmSBDizkLONf9VXPQGjVOI2M8zDTVA0au/k3uWAYv3OkWmHrB
H6VpHLwJ8+nMtirqn6pl9Blj2EJZmwhStkRV5GA1o1aledplvf9mmRnm+QB7WAaCG0f+/Ha66o+w
JZDyzhgdHRZAX1hTiJ7xnDangeiPofFrMtvnWJZ0b0dRa71b7YbwI14Uh38Lz3dKRVlRhOa1tuq3
6WfSKN0Ml5LQYPwypgDYHExsDpw9lTfdt307GKDjgmOVXnx++k2Q1HdGcNaozmyAAqQ9yvaaGT5e
yWixebmZcR8O9CWddmahwwx1zgFITL9jPbgaePSQaZQTGTklNOYwsFAxDiiJmxoOOscLhRW/D3Kw
yPiKMysMMjr+KQek8ePuXbH2HdYJScUL1bKvUJ1w+X8J1Cxr0pwoXWq35XAeufiVL79EoFOCTt25
p0Qad+sVftHnePXos0HahMtt7pQ1VkrDgGaXsLcDGhCXaxHDqrth6T7+f5B5rc3JKSWPUEAJto4c
h4loL030BjuXpDXu3uwMjK62g6KPV/Vmfq+FAS+GWpog61zTJ9xRsq8fddSYAec3NGikWWenDO9R
XusWTL0KeupLfYTdt4GuMqymzhyRUceW93v/auGAwAOoWPn0GPZagy0WeG9HUpdvtgCWs7CrDa35
AUIS0wgYpdCg86N1RGL4hSimyh2u8C19BeBZ3v6s3YbJnNwA4pXmPEcihUwy0eabpevkrNwXzbvl
axsDrqraw3j9Cj1hnV4gTn+b7BMQhP2i4a6fw4ldEX044fYKDAqIUMxwVSLCs3VD5ij0Oivc3txT
vKSOxrTxnWnUuAqaBvx9hKtV6Bw5Qci8h1pDX/qATJhbajmlRL8taYREEDGJIsGGm7FrAf7kl5q9
0RIk7iqgdDGVJZapQSbmyjJGikOQfEag32Q5lpJ9OIIGtuzMij6dwsilviquOoV0FA3x+YhGeK/4
kwfW9qk6vVaSWIb+QppNh9cmxx2/Xt5w9Sl+qdscceMZf/CocsP2suzthpXJi/TLaQSQhdBduq3T
gr3ug8GB+GfpWFsEDLWaRKVlfoRlOhWlp5Q5wwqltmfEGbLKx0JO0jpZfY4IPTRPOIDOZMuX1ISS
8d9URyUl36p0ukuxbsuLdDFQ+Efsr30jVavbsjfDZeOP3/FrdMTKKhFsNQT8pu3waT25k/AN4ibA
oBmP1XPPDmiP85V9wtoF/Gbqk2cdSVCbWIR0xiCsaUbmizXrT4VLvt/7hc0KmFq96TqeIN7fmv8L
zuldKi99hAimmT/F7KZ7LCWa4NpI2XKh41tNe35VsE2aT4HUkS95yzh/Q5+kOpl/+6psoKPjV0ed
aNDj0DXWW47hKpJ/Is+caVsfhM6KsqpfiqfgNcEB3GaUkwK0Or7m3tv9PE92GVHjUtpMuNAUj6wN
fkRpu/4Accs3zXLnpF5otsAI1jgSYYB4W6+k2ENKfzp4ucHLCsGky1fimtL02qdNqJUzuf1/sYID
xZUpfaNlOf29sNb+JPiVNhXygaSN+0owZ2xwPHJWpQG8ILK2Nx8fEIrIbSdJ/PrFTWKqESdFP6QH
kov/Cqx43KHQwmc0pS50yQh7Mo5+aDiziSjAspp7Y6/055EXTNzG1aTu45S+hb1wyKfLeixj4AHw
3j1WbBYyfbEcKbIqVD5drYnl7HuzDnIPoTpQ4Oc2FQ7KJcZEqnZa3q/7mpJdYOvQw1qjJhEnxijv
ieU/ArJYP8BUS/8nYWnMI7yn4+hUyJE2sfrxFKS1mgwqLJG4HjOQu2BC573It6AJdomqeCZtEcER
XG69P8yTY0FwthhNXaimuMMSUFqXSqE/ftfmdq8TpYMUcUnV4cNhMzk5OHPme4pZ0zg6UaaDhX5W
8fp1Y/U0sDLdkNcSlzHXJh7FXhRoDEMVbeEHU5UNq89o83lkbevairoB4DYrQWGPR5AtG1GGOE6N
X0jCKbt/aUrkk/0h/wxcXL2z40ugtcRfDWd/TQKroyZ0U1hPIaXheGmlutt1KcL0QYVF8qgwPcCg
d0s6mLokEiSEDI5zbsvK9QqIxqZhmVgtZ0HDAODPmtkWRyL0PKefINggKzWSMkleBETWEMJQJNG4
wnYs0LI8ec6SOm1yOIzh1NLynLoK7eH1CVegomnc7j1b8Fwn7gIP4a+gm9w5bzrnTCdT49zjejiB
isExXcXsy+Vek4qsN7RQ4HT4kNcnf2zYTuR6KzrmR+lYS5JsM0B7ej94cywUJ5ZHm8XErfGIZmq1
jNcuaWyE1Pd5lzD2CjcomUE4gKq2Wh9M9w/4bpi8Ti/E+owN+WQ+TrwUSfzU0VHKECViuTOhq3xw
D9vKRA+myUsJ6ozT1ReNMEpMEeKrf4QswRwbvHgNYXedpZpnVxoHol8RRFxe8Thc2cfY4hnarGhk
G+iUOrbQFQe8gjr/pCEdh/CLC+2Vfx+zARjp7LUnpvnk1rmPpPHomV89igJbgvwtSo0uFDnEmsSS
PDKgOqfPKwR/4IJ6HGgogBXn1NIGMscZRrigIJ1ztKTApNjyY8JOphX8n9KnxItMurldTLMhPYR8
1idl1BDfiVvUvcePQAqrldyJD2Yr66Ij9GAbPM97B5q0rIESaj6UehQsty7RQJBav2rMSix2hUlE
OrCmpIWKjrFzf+4W9DjmWNl8+jtUIX9E8jn8HvWUe5WA3iI9CA6Tr06Uxt74C3qWX6LGdceDvk3V
FGuGzyIZU3hMqeEjbRg3nP2DmnywFpg8RnnWtw1K5GyNVA9zbZVksSEgbTqn3gklJvbTPW+ai4RD
L0T7eVtyL6Wzg5peb6xqDwHVkCKcHtWmS6az8eQb4qp+pEXwXQB8q2/3fSc0gZ1N0fTcTV4K5c4f
VNbkRUnwPWiFtjsVrhcenJ+GhiPBd2DWH+cOetUsFZMxUyx4Pa3zCheQfYXKKAOiRVJ59sQBU4Qs
YjQXHKVLfTEbU1hvvxIJQNMAe0RN5gush9CiQ+97GvQGaz84Y3MNo+1rRV/mcaFB8apTnTHziKAw
DQHp3EDTyqjNsNpGWRbZh+u8g2+pj1jJIDyRwQRMlctyzG3JkXeeIbrPo4v2cuGxKkN2Fyhcqy52
3L5QGnZosGD+jB51SaQ1QvtGSsx+7aiWxyFIaoRom90osyxAUMZojnRtO5nYsczCXt09MpjtLPc9
IWLpxEt03MUTlJxTGTx6NVT2d5lraV27AlR7L4gFVN2eGfzBkV+jgHBWShayjJjk3nLavCQ/prGv
eHEYztaY5MmI44240O4TGG3R+aYSgZo6nE79Fx7IacElIVPFK6d74Dl7ovQGRG6zzT2ailtjoYJv
O9k77KQEhi+gr1PCNkaowfJBP/I86nCtdj5rLidGPlJfky+HadbbvP6b99n75AKEOWZHNvfP6qHj
zZs48ciAx1QDR5LpxzDJmnpKLvZ+WoL/65r7gwYMTWN2A4CwNhJM95FlsWZC5RG+IvNC8zpb4nRh
hrzEA+w1eukD5V1kgS7hBxqxcw33iAF+R6w5wUMCsfxmyq7fV/a30Vj3RJlc8JdHdYeq3rMFedOK
65DQeQOPWhBoSSJ2xN+tLlzMjMPc/DdeYzLKvciAYMOgZohYkmeYsYnkE4/Y7+WsqDzzjnHoQZXd
qy+a1dxaDo7/lrdMs6WoA4XZnPxQy+XnQ/13LvCPJnhE7363i8hNgBzi/LvpCUoQTu+uOCx9Ru7h
vt7sKGgMLqHhsS58c/Si+DrAiMuAsTUbP7gH3fOhUDagiPW7qJof40DSe6j/iR1fwUWIffo1SbCQ
LWBqaekjthGpa3JIDeEA7xAK1teSwE5TAO1c8/8mR8HKsrNGzFAXGn1C7JaTXzyKCI6VUqbXEwDq
Z576LhaulWYlseFCqQA3iqJQdSUXh3rYQt5Zyi7dcIpQZdT/rSlGhOTuSFbzdCU6yiAkbvV1f4Mr
qcdHu2HduBOtJ7tu7O5kE+mg96c9HwPFFwJTrLMr14Hk+Ky9zcA68Kwjp6Jk0utvAUDb5s6HurmQ
Y5KWI1oEc/5c66GQGSeB1VVcT4xj0YlTA6xtqDP4GcBEfGiDPQmm+KBdQ3zs+qOs4Cx9uTDssapH
fFB/ohOhthxb5V0pCkA/Jz20CcmQ7hJgIURpxkSdiqqscDM1iIU04tlygs8eCdSFCoS+0dbEEICy
yg5tVl8gowVQSQK3BnM6OQsxrwau5ktcK/9BF7RZwJUHKdX4U4HCpl4vo1dNXk8maBIIQ837sybG
BlYFpjuTJaUaRSNkklZCTAjlqdiieKPP74TZ/f0LSFZ+WSvgDlRt5yoUTVr7AIz4uLZ0R6byQw9I
WMdwevDrvdOf7cuuZnndYCDoiFjcH+LUXhExZm/ZvqfxIsH8oULWwhWyeBG9UesMYHsu3vlhIV3h
o2g5JTW0/9Et61q3JxiPa8PqQqSliPyp5tAgGG7VSOZ6mbrnMC2cJiCUYaFBH+wDVpYzOKugc3Ct
MOxFNPjN/5IVNNT1kfRD99J3r+Nr8wrQSTK+bEPUWJoOGICnXfejnEAC/YrkfTVyMSrTQ8QCNlHm
d0YOdlDJShoY3lmUGybImYonB9F0f3orKM2RV4ubHY+92RfcmgmkysvYrMXGBjrR//XB1m7IOWmK
CYgB9HUqB5tu3/fqfEBNlYxiDU1pWwYFlj2RQZkkTpgPYDkWtPfktBcPdv96HIG9A+myIpfCnSzH
VkAXRkjYBznq0ZxSLBFdVH3vnG+bHAzciPUtDSSsAKKW2diqiAZzX8JkLWaJf5lHoXTt+htpofJO
XC8WNc5sHfbpsYUFU0O2sxqAwfxuHSJbfiz89No75pyQQOCXlQ5IFhzo4gf9oRTIraivCM9SJ2Fr
+KiVBhC9bcIN7wJdtPxv99JxZT1hiav/dr7/IGYw2sBLUgvhiXaPkURCv8CoZWzX2cpcKu8Jo61F
tK3HDwp6n5BSN0fo4Qcmo+tDpmKM7eu51s78AK17Tw1VGAZRy9SSP3G+HeVAOpjqb5L5TcG21RhE
6hVydSpHetJt5QOdX3bBPpqjdiZ/HabyrCePYy/9748Tpgsi0VfVpqRBtL/4qbI4lipr5+06rKzl
03GYRdKq1Ygn7XffFzuQUwyUxAF+xNcYyW4R3P9ycAtZwG3fjFTjtFHmuAgBeAVQ5Y0II2bM09VJ
WCY0RzD5eca/FddATkartSv2NZ20tDsk6Kmt3u529lCnJsBYZrBqL61DaYwcVM/wgqd8+XZA30Xy
LpAOO4KQAo9JNQrKzP1Yrd3v7kA532rfiAJUKwAfZlsKKn3EbOh0t/QrTqNab3ffgNKCH8Tt6JhY
Rzy2ldESLGf1kRNxnQHQNwzIdkFp7So3ND53J4dcUU4pBEk6Cksv7yV9cQshK9TgfZhec5KCG6Vy
TeNsksONdwPIpoN6qM8WxzNO9QPL6VeqVjbMWllZUkbrPf/HDthCvWJ6GSM46zJuDsNzLFTFaEo5
gmHs093Fwx151N9p7+X+U8/eDR4oQyTUgpqQbery8IzEypJeMF/Wp2kgKtdMrerrZh4E+6w3ZwH7
rIzLT6d11o0ibi+Oxt603pCGWVCcaptDJn7d83eZMZbsoTlX+uXxkGke5LASMhMvMVwDxILmkwIP
+w7032T1KhmkT/A4/IOVqxfSjZ1mUmIZfi/KmCxdoImUAAIMHS/DNEGv1e3UbBr8DIsY1L296mcv
nDdt1qM7sT4tYYbqPcXjs8CQ4H5mXH2z1fy3k4tyjuLvqRHVd5m2LBDaWf1sNPqkrMtwVhD9yhar
WB1e8xD16a5Rgf37WV1kz4EPWV1gpA0Lu/9TvQeJvesM0qGwZh+apDic5kEMME1FBRNZB3bejrVj
voHQD/ZcBkO6wU00yEglCvRyJEhJ2dbRM6i7E6A4uwA/ViJiITt+G6q9RIkQcwlwyR7tuxQc89m3
FknBUeqSA+VWUqvLI38/d6nMJ/XrNzJhIMFiwFp4H1JjyLzGNF5PMjwdxEt2zl24OGufTqkLg9Bm
9Wk4T2khtdhbSx03jDctHB73PjBlA5UoRXxioFvNxOd4lkSftgZ8l0DYl4E8b0Y2JWoltmfLsLA+
CQ1HEG48lLmnn0gFGdAA4uXCyDe7Bxq+TKcT77vUaOr/Jvguz/z57L9dFDHfqaUs9at9aIdAaPX/
yXx412MRoSQfh9ye5gwvs1JQ0XW18HSTDEzt1VZRGhhN8eeCKRtaT4tgfYq9RmsId7Nd94fazlqv
1l6RCZiiQK/N4Ez2VLo5zMD5jDygiQlfk4w3BDR84EGHSPswWJIQBYtobYaNcwUGPpLo7oSHSWka
+PvqN/En7+jckmQn7mVFFloesN1twaIIX7bYpZmUEMM4WYR/neL/OZnbcdUdxka48Asjmzu7hzEO
L82JSIRITovJjk6/sble+dUn+42C75AxvoQEcv9fpoJrb0I606/Ofyz40o/1EEB+PVcMVGSZo8QY
YdhJULS4PyJGLlIcSzmcCgWeAfx9drQ+hKrJqiEhYoqO7/ETgh/TdmyWuYifrRJjOlXsE2wcSgmV
/x6v/JR2RuLpbbcHXemb63TSxjwDjfNRNSBiQGyu49pnGg3dwBP9GiL+d9VxYYn57K0ewija45mO
D5VxDP3Tou5Oy0ocDRbERB3aWuoeAk10Q9yA4COlO1pfr9TKL6ey/euNI7stxSd1ypiEamc2/TbW
NIAgIQTXFlapB5Yq2fmt0oCQDE94TbnNwy90EbQRruRNPoFLx/2cAubB4ioO025eNzfq40S7PBGY
NlPe3DDNKynqevYASN0/gKoEaBwmP8gBEg7e9raXodsNt9nAwL2Iv2C2f/FYHwXnCsIDPMfwX+a9
PPhUQpiH2oJXJtC2wonSgWYWnw/iTSbcD01gyOppZLnSWlglf6+mOqknWYcr9pIgXUuzj77DWEht
TXN3bBa8DBGlLXXmMw7diSaAlsdQ7X155o5/bEB5qsZ289kyFHSDmnWGjh/oOAcT1PgLN3/mSHTv
HbdULi3LfdqEDrYGX6/Qx3E+qfoBigu4VAUmVvY2vePkJXJIKnewIXs7I5E83RHsgHrpY7ZQYD8C
CAmhIh9+7lF5D+jaezfmqp6c/HYU3fmsPxjQNQwh2/qPj0BHGa7ZpmI+VVgJHBHMRBI3Q9aletuC
BoJri0Bj7LSCXoV6EqGdkUhrTTiFIPhUAUHMRjU8RHDhcv4xGFL0ITp9fKCOirXwnoY6pIoXFfy/
nN/+QQecc+1+jh4gY2wiHQFRZaFRL/X2GJVS3KABXvo45U+MhjXesQ+CePTUfjA8beWbeSEH0HEC
gfMnkheGZtVDPv9m3SUHIbZA6WZkA/q+lnbsdwq4VJeHpg0Vj8kYTaHBdmeTXSPqfNvbPceWdsFA
cGcG2DyDY7lcdxjDDnIbU3uQl1lcWluyDEdEzbs/dLQ51Qtj9vxDrYjPkvXRwjvbc76GfgdvdPMa
SpJWFjhd1a7ZmFwRvO/asXwqy4Xn1LPSu5vIEmkpwSL5rZAl0WudfzJCMja+CI75pmT5s4rSU5QX
+q9XpMv228Ho7zfkNbd38+dij+02alp8Tj8uV+/oAM58WrR2oYcd0RfSQW258zOsxNyt7nmqjmWm
OY67WeaRuhma/KAC2mz797w4CZS4myt7EOndU2vS+QWiskIgEagaDG2lYyLOo9S1qJ0nMFVrKkWi
qKQ9mIiCFQgHcGuSKs6N6IBw15oEGYh6gJuSnnlbLexY3EXrgw4iFkwpVK0phrFyLArxoKDBbm8R
bLqBIYTu18eyygn898NftjiBIysLy3RpeVapG+kDtT0oO84SXq1d0ZDOrl9yagFjuD4l1QSws3/d
GgDYXtIJv2zSUDKKUuHUh0Ocf9GIZ/QX0kplEHIRqAvoq0thfCN1AJGMxcn/h5F0/jXV1yH7zs5l
BiBctA7PcCOid0gRM92klRD8ZCPX6Oe/fBXnBVv3jJott/EK8M1wvG+UkYbSZEWFcVavRQROD7/b
t6MAXdv1OTvt2LdTTZ507Z8XXa19rm5DM9QThPPLIlnXZFQ9boNM2+jPwHNmqu1ezAd/O9d0h6PP
fEel92jfrEOAXD2+JnsVpg0lE9PMGBfT4rfdHWkx+TLERZy5vUEpvzM3EO2+ic5d7LKTary3kFRS
DyJvF1BTYum4q4L9DBzTewvOWfC4ysYF/q3L169mksGQKXbUHqMrKMxPMo8tnXSDBuqOw9CwN3C3
595nX1nUyFjCq+NdAWE3OZg8FDL+3KBz1sWgQA3wP26U2CXlEGBcRXqbk8s5r8LeI9Cxvwsssn8Y
gqtX5SyaReXhm327mX+G5eyx2okP3jt1yvCU2MUuyrlT1X8kR2YO8FWWJiomCxeTyd31OZAx10L9
KbCGbOf5YTckKYmXb6wuUB+a/XeEQQcyHjUtHMlG34IWLYPsW6frXvs9IwGS0HemHfFPii06r2HA
LHErrplgH6f/WhHZvCmUYZh6ShgOK79GrIyu9sfcUqRj3R4QxiDU6wB8cbXiWBEu++tDFP3e4d6n
sUw8TM0DtjWLFn7B1rN6pSr4t0XSsCaD943sqaWtxJP7kRABeUo4A5qSNgGvbB7Kk/w805VMHqut
MZIPPeKKARHAW5FMeGQbpGeIrrEr9d4IFRgsC7ALFaZwagMzN8LMERz0bkZxUjVbXdaaNGYUlWia
gvk1WGR7VCyyJ+WJ5cxA3Wsf3doObeEvDNZqSWC8ZhaSbSTm1ZRtGPUCLKPOhXoH3PbE4vw1wpdX
4/NBVPJO46WE5tGtxmnw4KoDGMHWfCuJzWxuazxG6KaYLKsZxVhtut808dH+RsNcjqGKTuaqWtht
NPe1nXVFWim80jq0Ww1eIP4SWoCg1uzfITVqu1B5LWqydj4IhSIklLNGP5LPmy6j8GSn9vDRtaSw
3Aj9OxAy56b9r5BkXhnCmyjIWye2wTo3O3j+/yIX0xisz1WW90s6YGoKt2Ou6vYjaLVwtOkPMF1y
3f/QfF1YVu1DPzDUFp/XYW23tZw1F4TItxYMiKfrVuHyAR83g5nXESW1lwpDgQ0WoBloPQ2dtnDi
80eySmYnvVhnpSXw39trxSd6pUL4G8n1NZOKeL1a24lHbmEYIYyTYva9nhN2iigYfnG9gMltFYVI
MXfPKOGwicHA/XMm+jrGFY3hHeYIqUKUYrgZ0HK9E4+hz/7idEootJIzz5bFJv0GzbAAhzkfAgv6
GGEeUNsLXR/d7bPiEG5Msvy4ik0VxzlMWhJEsIh8U+X4agSIEZLUEp4B67mOLfUuHy/lFtSXw3BA
zDhtIg+vp7QwJefBclguMSk2AXRY+bbQuTPgFnCdKtmjXFZz5hyHyPQ4wz4jAIFOxGYDq6pM13UT
2ldzRRbRbGMijh0rjXDUafUlr3ErRjkgl4OGnq1ZFaXcaLsMVLLcRTzCPnM3pCQXqDTEyjsnC808
HkikCPe/ZtAJLRc+bSv4pxaqg73aUPbcKGyjURQqbwuKElY62DCDMkeitE1rAvxm3Si7BJkBrKqj
v8KiV8O8D/4aDwAsy14oa5gHUOD9oe3JjHF+qIAFwcs2fBIL1eKv4n4AVvrAn9uf2jimQy9QFOls
koaEwKGJ7G3afxUOaU4MOfWatyalCZGZX/IsFi+dWnpatKTX7994Agd1uPIHscrrtZpq8KVIXoM4
rlgm6Aiwot/t4zJOSfbompHt/CImqicxoaE1lmUJ5tuyOrt6MQimS0/K5Gi4n0CRx6Xjvltjl+TL
2IP6GyMU5gm4Ix2Pcp4RmReOxgijaM2rvGuDvykaSP0S0Em+DRUCIRjkjBHk1BeL9bhIrO61HpJs
SQ4fTCI2I2OCC/e+c7oDJLLCTkADlojuSQdZm5Xfr+ybPRig+GE5NM8rkCKSCdhAVyqKCZhsiqGa
DV+1xTyil0NK9GVIvQwYW+AWJwaCCl18IaxbieHTxmVqRKYsvQg2scwRS7vTkb4HF+O9Cr0OfW7P
CFBzrQ0WkFbaO5wgx5+OERaBPhwAvSAkY7IMKQ7Sjqw+RKuzHTphF9Q6A8LswzAV0jaKpZg++MMX
in5sV0GLqvMcs9qRGBzd8F9OMOoPOq8zHLUq7WrBRcQrCvozt05qRhduy8JCRCJrdBcrPUCUtI1u
wDeqX3WTUtZCWT7dCDdzT9h0UPky9177bNVVkpZK8tc8+2Sxg+xZRQ55OVxxlWiNS3c1YSpTUrGh
P3DUEHzUObZaTLcfffz0AsimgRClkXpp2a+sE/Ibq+MDzACWlGFst2wKtrqXkedFaxvI28XZ4vK8
E0ec4860EnJ/9xhi+xE80rUgoc63cvw3GbObtxoa3/dnv07JtpLDvIk6l93gqpkSQFXG0Y5fTtNW
nWJisSzpJ/W53guXnAB25gDq3TWo2Lc+4Q3RgvgFnuG5opavz+mGNtG8i3QmHAiVrwttfrD6Thwu
xjmb+FnxY3ywDVki3MgUBRFPKc+sPOlKQou2CcOe8skz82wIdsusMWBCZcVYVCxzM4bVdgqIALaP
SJii3sYhMaMLJDnDX5pMYMyhWfWtNFMuwp9Z0WsSrpe9vMT+JL9ydTXYHEtlHMsOgovMW9OEiCqI
Y+mpLEvLWsH+DgpOsLF2nmu88L5ukpk65iSSFKV4zM7v3mmBqi4NbnMfMxbIINAd2dati9MBdE7O
IZd31n1qjFrlHEfM5ImrqF4dcIQ0gi0hNFKprB4zyoCwpwwoul8066+rMFXvD+dOHn/SPcT8z8pu
CKC57NzvIWmxICYY3i/3aU35Z5Ort9AwZUAsixomI/3vALs89JHyAIOKynC9rKH7MEHCV7sGr0fE
ukxQZHTNm+9gi6aPAUZDNy1iVOt6hgj0QEiLVfE5iaFWDJD+UZUPqSQ1TYTS96Sp1BfHn3+/zFR8
MAXnBy6ob2TXlt41+GPMa1AoHVp+ksjoga9lP5wcGmBxBFeiV8XvhJP0HaeFdYM2GpG+hIKa4kK0
Bz3MvA2DutJCdA==
`protect end_protected
