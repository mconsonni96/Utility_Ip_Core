`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
j3U1D9a1cKi+drP7tPKAN6Ovc/cbXWoDG/QIbwa5QnW7ska29c7cmSpJFjvZlaaBi8F1pLIPLT0C
z93LSbReA8h67vGd8pYqT0Z1Cm4VjxubJ+DGn7OwIWOELpFCdOMgDUoQyOk0rqjgabFgsSr/rJd5
gxzEu/oi7HMWFaNpvJc+5Frio9rD3UZl8vZ7GSopnjs3T2B1H1+PA7fdmDGb6AeEfQks5Jzur0xU
ouiUr9ujEJBjdSPyn4UCuL3zduk64ihiWqWxD22wnq6I7qIuRokc/UyokAkQLvEoQyV/xFli/Bhv
DW+mMW0gv83FGE9/7p9/XHBDGemkgunRRl2Dww==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="j1I6XEPez/ci/FrmIyaZDDaR0iEuMw3SHAt1EioWq9o="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11264)
`protect data_block
bjFuX/vNmkR9394VEJBVBrN5+yx97sWk3mtRXh8ehXvtWLFR/N5JQ/2R+NuMzKKKaoepsLpi995H
Krz8pUhmHdkWQi4LsbWVz62XNa4xCHvgenUBiJFqkm0JaS3JOC99P+4KWwiRZHJ4YGbFxOJB5kqe
JuD9cGQJsXaU+riDdaSXMBUVnGIw2SId9knEan3TIP6LgBvf9TVRo5ccI/nBKiwRFBOuH0sIRQ9S
mm/Z7LW4cAZiGn1u+v5BOQ0aTfxS9WfdD3q5KG2ajqJtTzWiM2jfcP7IzwZvMxNSTF0A0wI2yKRE
WAaCz0fF2quIhTSxzjzLJhKnGyjfzM9nuRNUC0ujQTxVhK8HnNvdEJJBS2iDltdqmSbc2VKLdyD0
Q4qscx3E03AI7VZBAXjQ8tS73yCCxAsVHL7fLyDsoc7lE0sCp/dHsH6hN50qW/Xm2wuynw9MzIUV
vHhA+aXCxFoAoRyplwbwc4Jaei2irhsB8qMOvRgI9GmrJsKI+8O2Rv/fGKt9B7DbvKv0nZkSY462
/xod0IgOlyblnO3bgfUEWmQjRhiZYOOM0LJf5/OSqYjFMPuBUoWLZOG0qPYO7v5VptrOtM2qCh1n
TD4N2GEeV85z5Hwq5pbvFaRU1gpDbi46OkcqQPL/ObTxD+h5ZyhSz47GvXLpy8385cPFEdYjx2OI
AwXLzfxjrGOKhoFJWWL50/wCCdN8anEUIzijJ8oK/xNxRxCzuptaBj72B4zq7JYdORNuZLt7uDN6
2VPbindOUKY3jiICyYtbT/xULeZ3tK5qY+RLINpuFZHdazqxNS7cNFv1V3jPPibmdnJugYiEeFv9
veD+rCXjwrNpJOp/QcZpS4nMLOWAydeLOujNqndTsPwXka4GAV0lcyFQmxxDI2bacja/Q2eU/e0s
uWqbtFhaVeKSLlx/84twMAgRCj7/JXq62yIBAjFCLOowY7jQgaDL0zsA9/VsHTcS5DGmbzKsM5/h
jlZEB11gccNwKg4Kmxz6jkGdczxSrdXmvWkjPvGDBSmKnXs4LxSN3nVxjpRkXoSCCYCJLeBYP+4h
fbPg1P2xSNSburvQdYJW3SseuGd6CGgh5tGArBybAaEn+os0TruslrRdUSxSdzxBJ6Hjwu3SXL0i
dkwrjJSylYxgUY7hPX87cIxVxTl40QlpWmgsLD8cWq5AgKk5TK4ATqVcAsf2TtGtR7WbjDjoJHSq
hQayS7elTBRdcFJoHGCl1IGLaJCAgSlDv05u+2U2UjCRWAvJrq5eS4iLFmtzEvXHNsla5+dODrSF
aCFkl4RAZ09OImANDE7kQDpfLHX8JrZB/Db4m84DTtMoiFg/4fogw8leFnmruteb2mpyil8FwFGX
qCtzoJLQsonB1PhpOVjnH0QJZ4At2DzPJRrDUX4VMrAwUyWDJJ6i4RYXZqkkwQmDKvYUH1OdKXzE
tuXz2WEdkVu6dCNASvtcUbhDfbuKx+uoUkBOgvQmQBK+yIyiU6K0ZSL2LLtfnPiokjBN1czY7/Gn
C1GC9NdbhhCER/t0tnRceQqW23LC6XyZcvt2sqdtoqfIUGrPrpRvQxdN9PuOdqZzTeV8vT00F6G7
Rddr9DWwW+6NBL+P8ooSal0ESto0GYlZynWHRhIAjvJS9ZcGInKMqsEup6tQnLDWSwt8sIplnCja
AFCtd0z2g7PaRlcVt45bilkYl8wxWxSxdaT2QYKJT9CGKvhHntUbpbsftHkuXcJYPg6FaDEE+Jba
mHSUshAg4sBjTVlmNnbhpLib5CYDbWCvTwO4QM0DPBlYsncc7m4VtfrTTdxKb+ub7cmphxS04H8Y
+nI0FcSAH2+sC4WeiCzedC87zhO4sDTAy7lnO/+XNKqn5LUCMSB6td4rbtIauNN7w42BqbtqtLii
t5TS6SvKRjDAkInNFApT3/W45hwvXZ+4NOgXxvKC9algGJ1gUY5r2d9B1o8+oxcZBD2wOyt3s2ig
rm+at9S2zQJSmykcXy7hPj3FeXLMSccFtdrGu35Zhb7Hl089bNTSHi5lLKfr5nSHUbQdm3qFG25y
JYZ8ke4yxF6A9kV+QJbwCOYtYY5Xa4w+0XvYzy90ceNIwISBakoltry/cFQnlsJyO6sb+zYdxdUd
UJoPDTAILStjCSdvNmRLRUv8/bJ6MYqstYHy93jvWGzZ22TD3F3iEjjBFQYrjg4FwLRaYmA9Qdc1
u4tzcoxq/OHBHV8+bD7ALGuPwQqitTMVT/m36fs5EtN7jvJTkSrcJQYJ2Bup8Wp9TgrHYG35q6HH
oORgnrKTK7ayZx/yZae31GFw5VfKXn863Q0ApxU+HqCOOx4Yx9ycJ3NtIdQfXaqjB868hE/EcylY
7qdYF8PP3ykKo0FQnbMIBc/IhmNv4oE1aTIS/+eZY0dJaaesjzswuAHggMuso4ujhauSky0jgbFX
tPQoAGEO1Hl4gWMCjYDS1d+BpjWoplFSIiqFUFqLpuLJZ3B1zkDvGb84Y5zb1mJBI2ByGsiFemaX
RFbbpYyXBVFCj3ZKbm07X/L76bHBjh+JhHY0VU4ztIwJ9GqRxX61wmmBhtEIsN1j52b62/JsVOeG
dR8A/6I3YZQoMSI7Atij8JCSuDxeU5kCQwRFA9vd8fEwcmBmnmnI7jfai7qmlynnbwrpH9fk/tcj
HsV6YPbBEok8LwuNWVGrIwz+XANhZcHHdokyFIi2d5J3hC8AnhI1T2zxoBZedTJwxQ5ciQXVRZpH
DPdin+EKeM5RMKXGSqDGwA04B5YbYfyt6cvXawouc9iH96C0eIp4aHchxJQ4b0IRn+dpwE8wY9Z8
w5z5oXxcio6TSFbdUKlXWF/MH1bOsLRBDcQUeTnEjoVAzNBUnk+bGPhrFRn6pllb0zgUxqshS0nO
VfCz8UWRD6Zi1xrOO0wDyy8nBaRCH+eYsLt8w7z4SlWj7kGZadeNkCExiKWtovex1GDcatCjM3Bb
HxO8MyHJ58JssQtnynvVnitQFiyjxOyG53pWO1Gia3yC4JsYSfweZsG1rqGHPzbjkLAVlu+raS6T
DkPJDipGUO1VUyG8bl/KSQbYV1A2qt8BFC5bMSR1B3Q8NaBkRbgcS9TVqZEctMwM91EoulzhY0V+
8t1GDzST81YHDTLBPC7vpOFatY6yT7YSVokkkweMWteYSGoqTYIDn1YeIbCLX9OJiksRO4VSSPeu
1ozbmu5A/YU7d9cU6Gs0ZFhx1Q/s7+58RjUQWbssoMD918H2oiFKRbU5IKSSEd+riVnMXZcxb4tD
M1oawGaqujpRjM/1XAW1ue+9FZT0k8/ErQvgR1RL8Ra82wgwCt/Ba5trpAbqfzqALTmA63sgFN74
6bwl05pVgt/0bemWfgBqBNx2t9uvwjYBd4sZjXoyqnr+cLcso0lZLqhsJZ2HhxGvPqhYLTZTGHLk
T2XpWlYZuH7xaCsyY/A1CDHrduLaA+6suA+KSyLvelwOHYr9LLVIrK2bGhvtguY3mAjGAyF5GIjl
tbiprW8CVEnySZA3VUdrm7IIA3GjaIeJGL74mE07uQqoO4VXu6CpRWK9OS/GTPfHXy9Dn5cQe3uK
CeV5K24sDtKhsg8E/GSA2aCpMvp5E7JFFDCKw2hXj1N7b1O/TGBQdjwnT7LOVmTNmCMvrfU6rpQu
sZtfvPsUp8NJ0JUAvTXkI+RGbjXB7sXIBDdENGShMmrGlC33oqaqxms2/+dwxqSjT9Ua6v+qXHDq
w2q6cucTS8I1S0AqlstGCy+kS5fQketZB4dJ3BACJCRJBEx0NJPBRuCNL8DnU43Y1oPM1CtxPYpE
ZAtFjC/YLKWffM4IcsU8yB3iY/DEgM5Xd6feCfOeYdFb/5MvYcmcFoSHQ+snecFfqzQy8kpVLXts
D0AFh0WhbccLB3dnm5zrulRLPMD6CqVLOoEW2neo6JsDgHlf4qkhMGIWBn80SpWcqkGU55oWGgkq
b27OXyaQp36mEGEKZ+IAClaGxVc+ilIKz58sERjmA5ahSsyuDnFSBmuAcF6Sg66rk3IxgRheUNHp
xhzVXuxB3M9AyQnMDSO6O/Fl4BiP4o5nkMBmwVrasvptR4zo+AKKxJhTyP6/JnaynV/L2rgeuo5u
u5wADhrwe+WpUbZDYnn3ggB3/8hscUfPrq+L2Fw9p0OZj+mznRp8f78PgLB83M3wWueqNxVRW/nJ
1es7bYFGSRmlXPaftSaDwTiej6tFeHh9yumPDvle4PkFJ5seCSqWoLpvwIkzIaKyNzGTeMpxASf5
uTF33JEETHhyZtEgIxIf5fVbmGHZ1QjWjN98Qz66jabO53QsiUlrOvSo0lmVTqOAmC86OsLRT6ul
BWaLeWpsg9WsO9HTg5r9K83ehtbDS8SvJ5N28DIT/dRyJN7smqS60ZtzBAy1je8gv0QwvH2ijqV3
OWy0f/jkP3vpQJhrpWXsQ4cSQIsSEZk0AJCyC95EU0L8EMZuBha1lRjDkrEDlsTd0Y33NRsPraGy
rYrEm97XEQtREkpAxzntZcaB/7uEjczDQwQ2dEejjpudAtLM4jYHqMGfNlm/0ZWV6maz03p/Mb/p
mfj59bg4BQXPOvEee2kIqHmzThLE9shecmiB43483iqpHSjhCw2EalpCTOW1T5IEmKNKN4gGpNEw
A1Dz41wionlHwI8jzJD0NGzNJjBZCVS1gk1UYPm/AY9oDenYVGkz1bilyRZPxxdr6oDqWUWp1AW4
yCKJefNI1j6k4/OxoBSd7mjxt9fqd8/0bRIyPz55BRKApGB3Ridt/+K0sIe9S1m6+2H7jKXdiVFv
Nfqj36SRw31bKBddYX7zSOGStaSqOZoDtddDHETUvZpOslsHaj/RgZvA42kN5W3OMOf2dJ+xV5jY
lTGGAZiwf8y/+RBK1W/FpfvIKmcey5Elu2E5Bo9HC5gYfoMPji7RN9n8p3+/mxNY28hvWKpf2W5l
D0euwA7x7hqWGmF6hALmBobpXVcSEAtzuyhLPuHriC9d3V/xJ7tw2flyFR7XYNhu8LtxxNP6sq0g
RMdC0lH3Q2mPyIR9k8pqjw6OShTc6dfb4e63nQxJ62rrdC0qWLiCnRbZWWDAqWL9JRXVVqWUcWtS
PssXz3BZPjPNCAjnHQCtT92DD3tPQaXwIdQBtHsyMUX9xOxLjSnFjdCzOhy3GIGeNuOdimslecEp
zttgmJ1EamVp40I9hAcxLLVKG7srfx05hR8x2OouzxDqRtjTxG6fLWE98pgmalgsNQeysE3ym+k1
kfxrd4nlB8B7jyKzYX/2bClNwIPJSJ6wACtwhfV6BK5Xq1OMX7u/3O0Q47+Nx0wL4un8LlJA05+O
DtX99nM7kaZHqMaze6DxTAA17dglofkgRwZGy4MEgd5lV7HCpXrIFQktR4cBvp0rNsoocSpk25fZ
ZApGSwxgiCQhG16yVRckz8CKLhdJY+CC+zC3fNrAwlkulys6KVF6e4NfFCkQqc0Tki0kBS6iBcs+
c5upUtyevNEvA8H+S5ahXn+atIAiELW8QRMPBHLCyOCgDmey+LwEOQVIIuIDoo4UgedlbJqpIozv
Vf6QGRcnnyFx2rizK0SEOnk600u6HBSbsC012pLwJBiy5/BJXQAjefg8vPI5aRBVoMfnaHwndfJD
abPofJYLsb49QROD+6foEHLE5dPLr4aA4qeaTviU4axUjX89x8dBQ1zJxoqifC9NqEiy/eZM0vf/
jjNyId0823W6ywkhp4IWToP1/sxlyfCbhTHcTTMGuANEhAiAxB8MoFROib0mW2rX2Zx9Ovmh4CEG
i9+e0YFjGEmQQOIQo/LzZGD6A6jxc9dTHZgjB6FpcMMbNr0yC0h+wCCEzmaRIXsxmFGLku8f8QKC
8Xfe4FHNA4BOY3G+kqUrVd3MblwHelTBMjihfQNDxrQLUCRIFEMPnCtENUaSpD2/pos39ow7l4IG
7G4a2IWM/ir7maGF9ggHgLbA7j3I7M2TRcfF5E3qTlgPgKaU9gUyec6xxii4YhSyTpqF21/sficN
hVQFTDiBojNfFngmRB+/8lQm7GWKp5wsIMP7EF9gzxRoej+WXZrzWpWMirAlYClkNBCpnWNa8mnU
ALwob0A5ald2Vo9ifF1CyqBmq1Jwuo53kVnjbko0rD6h8yPIe1yc99QGdyfWpKgpg+qREEBTbhB9
HfvU9zuTSW04O8hO8L9wvDtfYO6KPLJAtjDMgZIqRmcpJpkuZFmiMnZvtWx9yx/XnB2fsIsHklDB
toOr+wZi3OnYjoY/0KNAqn0z8VKHb0avaMDCaYmndwBywnNBRaRt7OxgbWn5sHkaGZkD2V1i3rq0
kDQC9gWQXoOvIAO7hPjfYMK+XL02R+G49TZGksVg9t4UiFMqc0+RylWnAi3V1d4nDmiVEbW8G4lj
ixUDU3Nuzj88D6wAJnhV5WwWViW9++Os4sImtxK+SHTwH/T+4qipISlW3d2Y1dYy1umvX6ilDTvm
lTDmqJKDo4aRYvCwuusQ5t8qd+S2+ONJIALnn7aqmhCZD45DIvyg2jbO/3GBa3WBBCliN6mGNYFl
0EsvjB8ugV2p9HsAKWjsEepeqjkvfpnikOeNj1baWOjLufmeiR8trfisTuiTTsikgLIwPuNUPEGw
hAXlT69+emIpHgSzLkj/D0fQQDql5O+qFpbEse25iQa5UZcLxd4DpSr9XQIU4c9wAjH35E3MpQN5
LFMK4n1Rn36oNbhcPykOuSE4iH9xWIr8V6kk+cfRuPcX/hZsGlaGQj7gzaMDXW0Wd7pyM2Aj3J8/
vyQm1A4IuV7EWpeMD4nBrHjbhiQ0QnHvVtvHfGzTKTLqQ5v4Ug+vXEI4+4l2y2OfwFoC8USpG+IC
YWX/JAiXYOrAwhHWf8u6J60SFTctsMTUAHsy0kFS5GTEBzV2tbp2HA/z0boABdcoEG1ckjz4F5Ct
+3y0od2B+X9droGe8tw7+EVAUnrKDvwPPcr9kq02v8pMU/jKoU76swDViQ9LnvQX4wiggR4rAMvp
te6KMhaozRY+GId7jvqectm37zCfE6abFzbMwbt0AqzxY6NC/t2MaYQgsIB0gaZZiylkiyHtT2jv
CsZHSLh4jpTV8BpSR854UGPhlthC3rgsYypD/0onHVJXfRri0fnYSgiJrhPQqXbX1SbsPy/3fGX+
/NkrLvaGaf+lmbUw72yF6lRmGNIdaKBYIw+s/fEFI6zJ1V+8yP5HI3a6GOlSOjVigpZwzr5Nbi0R
FlwDoPrxyUCOjN+ITXvP6PQzbOc887NJ0MMUZ/UW9EbyCr1eplm/lNHEMMH6EzBMV3I35PMiTvz6
FF2D0u7OhTRJIhUdu7cOO0hX27mo5Y0Y/c8FIAWXNExUyQYCC6It63/XbQdytgqkhpywfQ7KgkYR
3Q/asHyyT602o17AskvOMRkcJCdVbc+ZMhK+aC/gsU2aS7EIw1EjV4KN41kfHpZ44U9V4ISt8ppC
5OPSHWz27NO2kEXz5x4FJBuw2B4hpEwcxGQsxn9ZgLnRPSckCBfbCzjtlQSuIeLyBAqWFuA46H7Z
jYmh4g4S83zMIYcA5L7F1xnXgD0rKzedb28PZ3RGVwI+y3l2Gc66aVBDi55e53PXJb8gDvFOliDD
ZQ7TnHBGtLZIdnUV1hky/UegpE4s/PUYvZYZotDkz7zxnc53rkx5q6B3TdmRBzmj32iGlBdV4yfv
KvbfOL6Uu4BWBP58Jixm/lMc7JlHUkR1oUP7Ao1xCID+SPQk35pchxs+ERlSUgpdYJNPNL3L9M41
2Qnf+4RR2YEE4tGEj4O4J6r4FdYcnobmaRlYweWx2QzheFklFrjWBYKo53Beo6+9j6JP4C8fsgLZ
t61++CNSuH54J7Lfxt7RuUFKwO+mp944tZEzYH9Sw0kI3a/6yS+qISIHD9zBM3EVW20mjWZTSQHL
Dwgk0lfgNaIEsHRlJEKEEoW/78UzcUE4H6dqT0HQWQVZIsk6ZTLwhUjlXCiiUqCc+/Ep7fUGATQw
6/HM3Bj6XWUe7fyyxLbfC+m1G0YmoUOFfBz4fm1bSxAk1Kfru/KS8OKeh+K7Z6q67gQy1yKlZW69
cwGnRzMhE8p9MbQhe07RV7h+aGMSPanaxEygt9Uvc1CIT3PZ0cu33rmoPn3zZyi+vcFqFjfxhhz8
C7ERO5RzhLlHwF2b/v+mczyKwK9A9kEHJ9ncofUuVRdZaXdI5W2FpZKyv8Rl77C36O9R/jURTotK
GNG/E9uyvfqhSzAiv2xiXZ82rOPJ37yd1dKsurHjYLg13V/4+mpvDZIZByVIA3j7vwZVV+qgkAsg
RqGAseaIZ8sx2/6l4eTEi6Q4vbmovuiDhyrzkEocIdUhsPjqkJ4g/Q3gWAz7zoshNsIn9qwz9ZSh
dHzg1CnmwVOCncMRymy9Y6ez2teVmgSgm9TIRzmDxqpdStMsPpIu1hmVw1BCH7V4b6j9Q1qp5CS0
w7jPlWWoc+SYDIEsY7u5A1efVfZQhwM4M2ru0NzPYXKcc0E0ctq9swDKJuiRb5Gt3Ge9ihh/nfnz
59J35Fz8UNLBFYB0XT4FhQLYYREQ1k+OPjxxb2dswcH8kt1gwY786ae+KRTGcS4P3SSiElaE1ABm
tFfy0gku9zS0uvSAeugDruMAxHWURpETNbciQGusYW00JTDWVX9uWZw/jgQe19qO14/NSjdg8DwK
pbUSa78r/0UaH/6kPUiohrnXBXoEwmr486wkOFBcZ7xJgEaWkvvfRwncgNDFsjZJOQ31SAXdNYAE
DhM5ajrcoucyp1vkkJpqdL5NoppCb+LFS8rsOulTUJsmKj2mNlqfTujUi4jA6G1i37965i3hTXOy
UHRGn2UkQD4jCqOJ1RBtJS6E24+xpjB4AXpMqVXdbCRN40O1PW15A1nDzfP7B0aBa0yfzEjNN8tw
jOACvHH5QyiUiAArewUww/9ivYaire7IpXxSZMk2BWPNbb+zeLubT5nYGkB41SAlGAKSBfRjk22J
wNiVvwdNIb2M9f/7nQsuxiQGBk/cxcnnkbv+v8PTCJfcsXXCydaAP/5lZnfrZhZNulFsTkvl80G8
PXthprqaL215neDzN6XtuDfA2el2o0tcmEpHSFaoj6KhD6urbCckM7OFEobpf6oOi5380D3G3kHf
mrfaZG45EJSqTndq/syqlellKbDK96FRUDOuc3oVqWatib2d+hU2/WJQcG/gDvsKva4Vi6m2v7OX
QFz1mo/JPobxWNX5WqUVrCjX21D8xhVqpv8JJeynxVa+uLibsd5d3gDJTWA3rkfiNcntc57fUav0
htQDL94rFK2AfGtgdxfT7nm5mstWoUvdS17Aj2OyWgvbJ4YB0faie2EhBW1lqCrWeb0tnvE4j9Ew
SNKt8ju1R6it0TGLyHb5m+J9WdiJiUrYeoQsWl+GXj7g76fnqt4Phmp33VhdcGSYQYS32nqJnkGq
IaNKXK85xiMQjYkwmFBY45QYN4ZJe/Lttz9PKkC9r0N1si/zmJ1L4rR3YOzvWrS74RNDsGozfoSZ
UL7kcxeWvE9o7ijWNUfR70ZsP0ft6J7XvXPxSwEjod2MRvzDfcGbhB0qXJPIsqlR63hDnZIeMxFK
L7tyq7tdpcd8Sh1dXizWLExPhpXauFXeppJWWhvSmx+/IXtulOmqfMMvKyPGfEGQ/XW531ljr6iy
vVPvYViqvG+zOSmunm+eKQLyeuRwvDjF/QJJpqvC+Ek9q8XgiG56uPJQlH5oJ8hg2WXSAXWvU25W
rQnql6FYrKXHJZV51WLwZchXZQBGkjV70ene7noyhUW7yRU1sxBAXB9E08QQFwEs6XBmIpXmBbrw
gNEo5mj2aM0NuU0+tjbz4nk13H3Nb7YtQh4NaVuUuxbWlkE0NHG49Pz56MOrgBCvNs/me+HSjEX6
qDWIa7y8NK+HfWZnvY0PZRbB0dDX8iRPbZrOTcfehfgTpfY/66/ph0g8jnUyXyhUALACuk5sCykS
NUstlSIz9giUQPRR5qQNzHNxSFCyoRSUdNC6W4NrLbRB5h9R/SVW6DI7Aa1/UUdY193ek8hHVgY6
8TIog/ED8YYcasHiwrwOItkp1HXcquc0oeEiXUyzgc63zgVTvBH8NL4hsOKPBySDdxHFj6XboMo1
kNBRwZ6jBGs7KhQ0TvSwJT7jVTXxqLdrXrPeJD837UaKfs6zGn1EmFZWRRDlTLO/whkUtAEs15lT
RP4yS5+0APFaYPZu+lEWPZmtk/YOpxtBjeD97ONB7Ar4vnO5ZoPjVO5v6wnu87jYW3u8/bndHX+Z
tP/NpwRC/gEW0wuTduM2Orky3hi487myOj8U0GkIvGeQj/3NiN2Y8E3uTkT9cAUrf29U//1b3sA1
bCvvSOmUbLfew5BQxjKWCSJdyoSak+w/Urk7N1mrxAPfLvIF4gnAY/p8O3nrozbv5lh50kOkdt1f
Bf1e1H+kn3G/qP+wpEL/gLmzIZHClHPdG4E8+YiAVtKtGDa/W6yUhue00Xtpya6CnAQo/9UYhsFG
O9a/4WuqyNA9CiCXslw8Wos6xN18iiJt75ZVL+NMqlqc56jQ60U80pplorZ1p5aP9eQDjnW/++zE
6OLSAjBnH+RzqSuB4pVbtmTbZ7gMOvouIDJ5B3uSgF0GWKhqn+UOwa+/rsqH/vpVNGvw9bAmM6dl
6iSZ7kpJm8jpMPvPaBTn9birdfF5HTE6M9UzADc6kVRgOo4+PPsgdq1r/fZZMcffuJ7/sr14kNdO
1XMRebJDT3FCZU+0TXmVUhXbC+H5J3+fbaGgtH2TGkRb71As4OctyroAIXl0oyY4dXCsu+2FqpxG
Qc4BY9qF9m5sgUW+ZDuYrRx99cZGZRieKLfHE4FXbXiyjNkx6BFVLDR7t59jOJCJFEPQte889Idk
U/AlLwM7ucH42nUH5U1iyJ8Twns1dI2OiczMXqLjvdmHWg0SBTSJwnyfvS8Hp0p+pfcmgGPL7D41
yUtGN0hiROFeITYtcqSLMWYUD3I3uFikqqhWcf66RDT8LFRhg9E0uZUa1HvyQfT9Oet7BfM3fyQK
t3DXjJFlpy/IAIdP8ItyBuiqRDHR75SJohB9eZRrXiuRFHAYFAEaM0XGORtuh2gCI9JxR18rpQbv
HbpQNBn+cfx9cHgrKsWKHPBwsd1P40v/DSQFjFnIbxT4hRPG4dLrEQLrI9WlaiJixwnjEvmI8Pb3
jd/xqqZNj2h18TNS/UuMmLuQBVZI9UuFyh/O0dZWeKlskUX4BuiHxiYQhpbKTilTSPPHsktMMFXe
nFH+6j2UVplJmc5rq/LuwF9Yn2qhFHk06HQ9DEWLUBzzKwJQ/2A3okxn+px/8lv+FEkgasNsYplz
+oR0VEo8TLEeaLOjn67Tc6TgPSQYkui+fShvcrqfOs81iam0Sw8WDUogkfNBMnQjmRdfvFCYYgKU
shmyAuGZFu/ikVFG+++MknuG9FRahgeGXwCSMxGa2WxarNwFKQfiAY/zd1TbgIBCRog0JB4W/MWH
iSo4sF1X6HVbl1uuH8umYN/g/5gH2lLPEcwFHRf90uTLqD3/381+DbedIUq5mUgbNE4G/jcoYBUv
KiAagHDHLNjI1l07IH1hnvB6/ouLOpDQ1Z12gwcwAdCH2sSdOVnJfNqbYTUSrkw02N8WN6FPaZbk
R/K6N6wa5ZsknvJa0NpIAE/RMuTyemn+DbLQHMshqf9k/SyUedTYXzZk+FO81vea2vc+/+bk+lDY
2i3RJzCoM0TLaR6mHS5JNIP0CuYL2BIJs6fz7C85ESIAPewZSFJHd/j3kZCcLFq5yzAJuLl1igVt
aL1/RR7n0k4Xxp0+VP0lpiDXH7W+lUy+zDSppzQSScIp6ABXxWmk7TBRSCYYeZ/FG3tGhv5TOySj
SiVM9YHvP1KDeYlo45tGMfpzHX0PqRAJkWBpVK2IOBPyo23rvFUm+Nsj+ykqivF3THnXN0qK0bmX
d7WwVfYrjRcm5W3sHC4jz84JLHCbazCp4mCU1ezsN1Uy2l88CMb0WyhOzdtJQMZG2rIBifp3g4rR
UQPVEXeuqYfBNl4pCXK2wwgqjNDFlE7oYv+MzLmBfuoFIfhs66l9c4L9y7xaCkHpEHRp4x4sBEG6
LHwoslpceei7YLppGb3itNq6myMDXJl0Sf4R7KBzXyJkY2W8EFLVpXI9+oOmtOuvsltY/TLN+2JI
qKz8ltCOS82Bw09C5A05WPBbnSnxirWVq4+NvxctZVIlzltPMivcruTlfFTIkSiWJwkkxvvNy6MB
cyB59cI66gz2GLmBOmCJDStXsMDxzSoWT4DdaqGD9IMhpsx1Hwotrhc1dStPaq+To/g/iunw+5/7
DoaqaZJ9yxPqKAdko7LS/F2Ba+CK6uJoMmXs5y7S0uzoTAg/IZgfqrH68wTpWzMI2UotlwN/6GI2
k7G2uR3FQR7bmjSvRgye6vVw0i9N0VSafB5a7pYUOHuAZv+Z5cEZgFnCdqPv/KAWtfh8Ct+pTylF
0Xe5FVCUOc2+b8aYq/z9P4P8X5b50Vr9S5WRhANcSHgE6FdMRKViR7awmSEhQ820BmLyIUiS0WCC
mlen7ascVMErqb/NxycL1HF8tFg9WS/k1Hxzui22vNpaBTFPZzty8E7xPx99dSKVp/0EKF+6Y+on
a3+wH8/d1RY1KLeEScaGbc+FmfUpobWlOBcM7ca4gUhzShNAvsbhz99gxLmHQXhyGyQZDuae4xAu
iRoZfcHXdOG8/TcBS+xUNhQ0biGPPQbL7YOxc+gZvj5m39SJszIB0UAHk1/tcOLcKm9B3hAMd8Jz
yeO9lOoTVUflzvIAOSPr26eNSDk4O0mHAWuiD7h1cn3gtP/JvtHVM6zD3LwFk4N+xY+RSTGwj/Og
4isULQrHRpQRBKJonllGMoupPSVlOBLRLlXybJxtZwnq9sZcgqxACMVzABVwRsCxLWTIc7NeQQkM
I2yz3CBrvJaxGzGh+Huxgh88yRDsbUzlTHy2o50Q/T3z73WT741HdIWHMPonMK3EQAIVZ1HiVil8
8wDEFm04y09cfRrQSOkz3kUPUrhT83aTPkySRM3HvURNasvfGy+QN1808foymprbSbyWykd67aCW
XdNLSpixjR9SgexCRhxLSAmUz4JgcAFjy5Sj/do/57hvOrkAPnxsQEb03Wh2v5Kk4nd2c/N2IQ0j
kQ2s2gINc4rbhiKLMqI9co3DnKK0P7UVqM39+WTGIZ3ykn4YWFc6oY2ak+LTggipv+OSTtBIaQFW
lChi2BbJiFCFBsAgOWAXJD84dzE1xaE8oD+ReBJR0szX0bUIET1zhewp257zljX9nHuavWuWl60N
OdwJfQtnVuILILXoA5quo9A/faLUgthkRDhT2I30u2j57mQaXPP5J4eWgmjfTJaWHZCRota4wkde
c8auGDW/zelrNTseoEEoI7DR039XmXvrVbtF5t0whLotg/oqEGjDoKxO4tjbwxtq34zjCIGKQEo5
rwgO6ceIKHUxOSdv9UfEunG6OM7cl6Xha56Bb3fT/zHOHFTiWVbM1I6rTNEoiGIl0E0JFicgj8CX
/g/PMbI3J83mkzHjFKZgk5DEja1pjQ2c4KRLqCHElz6SoxLJgljZyXmoiQcRrKiSeXpm1evCxbTj
NC6MDAnNcWmJtxDg2KmatVl3/qnoZP3ZGXMWq0TbpZqcG57e/2abGfFtfxdAF2UGEaKgTo2/10mz
fHRcW/SE8Gc2onE0ShUF9iBpDxlRSfR7RkQabL+icI+cwTGK+ekCwJK33+NqJ3Lrt15XuIZBsHTu
8LxWMUYpbaAVB+Sm/DXFSXXAPpGGeXSpCOkVQ0o5U1+rRENk9+5R43S2TCMXxFV1vVCqFxjQVU5c
ymFQCXGG+VXC7HWz7N2WRddQTqwR+LEOIumWGZE8QT7deo3OX6a8/gMnFSOTDD7JDzXJHkbKePVO
NeVL24FOPAqeeW+mfAWBcd8+VSwMQija0dDTf1FwbALW1tStmvaHzsODtJ5yeMzWJ8asIQ7tBMKs
+gZNqVcMC9aXIAYfaEZ4sqNREKvFvZCaoEQufsAQpX6BblHyMq9oMqakWzggOkyhSxj0eLOB+QE+
eBW873ZDT0BKSERErmm7jW0/JG8YIh5XWPQEeCFErPIgtAMn6TTiX5iVmHtlN3F92H+X/K1yk5tA
A2F6GAVHV50xlQjGux7JduT16z5jqhp0XrTASHy135pMKCOjfnHN5LebVfy1w9tdoozbdYYfPJjh
ladxdqGN9D5GrbvPgtBYCN2duSsNDjFWyk2wKFnTjAT1wkHS10jzjn0yQocrJ7TpImz/mQe66nOe
FOi1X4MFSHEpv1Q78rMw3TVxtWAsrMYh5HLLKbhuH/mQe62x7MNYaAtBtoFqmPAT+9Di17Pbqgdu
C2tzo+fX7tyLq41N3acoORzw7SuEhWAJAtx4fQAgXTkKUqHYAibI4pIj9T3OChkV3cmGUMzXVMv+
OqPXLQ8kFGCPfqRYwvZeQ8e8K5Zsy+slGz0RVlCEe/BYs2VReOQaE5lvLrPPwFesv1sce9beQXeJ
Ws60tKH3eOlmVnBZAJHqOFSg+flo70GcKRRg+4RNOaLqzJnD3WoXrf/TxADxmyz39h5YHsFBDLu4
yHjrEB2cvNdFsMft7xXDZfKUH37OvgZqsqVu87xQXdB5Uxci3dCnSKUNSxPzQsp8JaUtp/Kj1gew
JJilunj34v4YxaFmXixfTrRDTG5Ed39ZRSftnnBU+Yt2mnhO8mLammUbmWfWKY3RjGq2Oqu8Ko4x
YGKabSPr8VRSiXKGbqd8sK56Tnhe7tXtH6S9TGCQRWfMdk8bJ6SL2Ca9y+L2oj1amj2nZUTIcJEg
RogADkFQZBhKYOjg348cPaF3r8sTM+fTzhN+FJmkfsSTVFR1+H5NHY8IQ9kHmL2zqqUZOLPWrDwf
6Z4fzYJXo1Ew3HZLbKicLEIlS7eNnA89xw35nxaQRxtG4lyfAJvwn18956kwpbMSibw+BRwRU9sO
P5EZXKzml443jr+VvIOPFZvKoSfdvT/fGOCBC6WKb22F0rA=
`protect end_protected
