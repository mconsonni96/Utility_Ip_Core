`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
G7jqE50vHS8lRZ+WtZpRNVTZa6O9SyPx4JizO/DQi30/jFYzjRKurWtvlO6SgJjSp0yHJYPkdkBe
n3Drs2rOw6UqRRijnLV/gKUgGs7w9gUwsnc23FgIWUc+b0EcfCzHqQO9qz+RaZqoAqy9ejXX3qyk
1jg7D9Acouu/fj2HuUlGfn3Erg/EOVSVGMsFt8pR12RA0KhKtuqr75V6NGpnBcsVJJbnv6NoJlJ0
br9a1XKfGWGlliwWxaqvSs5HkVfPFf0rzqX2pDs418St1NFmLKO9UUuvp0wy27QBUMzLOAZ2abM9
r272II84pUpj9xxnQbFjU3aYd5xdLJlGWzGVkA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="pW819Z8I0g4Zpz6wdlnLgh+mgS3yTlkxIWMsgNCIl1Q="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19936)
`protect data_block
kJDd2PpILystqNZ4J2VnfgDinK4d95WTAOU/tLwgEfE1VXEbSJ3C0QKF/bMsKoWebte7YunwqwkI
Fsf3hSF7X/sUff502yvKWWnFKGnEO63mthQhzzHbtLlJMM5DKebD4PJQesRNDbuh6oVP4pecBMgl
19Jv6iv7WgyMgyn6snIYmx6GhNYmgb7aABTjmbeHbLDh/BY8xQm0s1U1d76ILR5aNZKcsiJbQ3Uz
Cuxd/WdlCwiq2tU689Dx8Lh7V8x+PnYWEBJAMSwK7cnZ6QYUGWtjFYNSYpSsbg+ziK70K5/SVTF5
7wZLjnV1N7Vk+A+/8riwQ3K/VQ6vXSg0WhsAhPPgq761Asw1EsSFYNyppB+le+/Q/XOkD6BXj6Sv
sXzqrov1Qk1hCcC2OdtUHRDgETh4+f3qyxS5OxY58A6xwHqOvfU+Lk2dGJhooO1M8N8ObSChfZ69
qm1SBSqX/Wn1LpA9PRStPLJSe34v95InzadjuP5sAa5dsMycnx+Idzk5EKW/p4NG3RkTg8wThRTF
umxkBroSDg1HR2vP3i9ntoDf9RoIHUJ7Xkz8vYXa2U3rZStnTknMj9f8LrSoMskNHWvjGb0wwbSG
sgKJngS+C6uftPUbHsOcK1tw+HUiO8Ad2B8hhG3S/E/9AaZzF1mYQx4Zv57Q3aVm28kxzlxCPLa8
W0f+CV/bWBEb8SygRDWg4j8OyNhBFn2WgwtgfFfu4s2f48YE3Jse+n2L92NjRda1iZ7DxdVoFe7U
E3R0WOn+cOvbBEZSnpT8cN6IC6tEvPyLmycjPMPsv5MfVpWRzTni3M/kd5wrXXzAni5iIfpdMwiM
bpuzlZrCOWCP4Q2RvS8YcB9J7VyPJLSaYonDpDxBfmmZDBt0NtxF0UmE8IRTx+ejdH1i7WpCKYF5
OHznB/FDMfYb6PX5qWhBfghXl8pyfYqa8fELZELVKYu4b4UzI/8k0/at9coIiuEBd4d4tWhK7zQ/
qIvOshEs5CiuqyW5etOP9sfd/U4/OQX++DrmPPhMIF+9c3GsSGNa1wWMabRlMEaRXR89YXffMk87
qGiAK5IJS2HNjwxUBmcw3kQP8AIg4V5AfC3HllR6yHmOkbIZfS2KVu8M3jCPqjCvdEBVHAfqSSlq
rPilJF7/rJnnvHagZnU7MEFCuXAorpktEp3mYB7OT+cSU7r7kynU6WR+roF6HY51hY57dHvnu/2c
m9GpfkF0EQjwGwNLThcmvQtjyp81zw7AaKkJe8wc2gpE6hLqJR8rwrgLZxR5qiPYR/dIjdVcHg70
/IXsbDAAc86LjAO0yHynbSRJj4uEkC7O4oxKJR1we0MQujm0d4riOlPgfk6F5Ie7PRseDIgG1NDW
THDmkJjJF848c5A8GqpkGiUcc06xQV8n1PoJP7BWShJrawNz+UU1PshT+ax1yQnvLUzLp2cjtnEE
TXPV6s3m20iaRC1kSn1OhSpIF/ZhuEU7ll0sbWd+7Q0s9D9rOHa73mNSNkF/+1Gj6lqgoU1vAjyc
Jcv7jrCfVYxT+/nt/eVPtShjBUILZ5UukF++KK35Sb6Cz/NBJUMKXUwC975crxHZcSZiSbL8zO4O
D0eJD+S/TcRZfhllHNxEVin/D5MqTS1GuX2yRofpUgTaGW2cBi6QZu63VQkwypv9X8aAjfjRqkHK
vE7MnLDrqMxdAqXsf4+Kvi35DlfxED9oBR9AVo8/Y2L5o6OcQCBkRwnh2qdTfzgHDa62VXY+JEC+
Thjv4NE+ghftdrUukHa4m35gIpc17LpNHbdH5HILdRaC4LUS1JEAbJdCDflmV2UFr+INHOjXraUs
/qbUcdTtkkSpIZXLb9VJWT/E4QhDZ4c4XzhBzE3tf7bgXvVfmLHssbyxc8EhKwzM/GtBU/dG9IFs
oizwg8aielcOacOugXvbo4zc7b5P+Q/U/KvZj2+khUBeCSsd64/JP7BOutMywgXdnpmqJUs5DnHW
82RYz1ccjwRHTCjvFn1Rpro9pGvSmX4MyI7dwLHJ1AGPW352AMqLo3AXyLEU9sIWdgKtyUXSXyR8
PMAZ38fODPhzlGylrrl8Aoqf2FGHRuInND6pBg5uPJ4y5XsvRqNGFJjdtUb8i9S3ZoErF+Q824ZQ
ydidmZp9R8zSSRu0T5JQ16Dv8p4liuMdZ0Ce4OT7tFf1ugAj/W6PaEBg9/twwdc+MErnYFawWfLl
1Yq+37VzLTJIjGJBKKH7eoVko3BX7A9+sV6r4zoVXEKYf9lQOFb6PPOkhRqtr7KnYt0dnFuQ1HSi
kQsHjov/ZIcOmsL7VEdeboFHJXgzBgjjEqC+NAW8cNzLXCTIEdeEJLHL3CIkgO1GFY5gPYlDGQzE
sm7iDAWoJsCifoO+nNptzdELyluKkAOmJlhVcw4yfftS4Cwos3wEbI497NXyz8Ac+GoiKwuuOQUv
x2XFZ+IqubvUvxPFoPUv8vGRVQdOfmO+8ml8H4OJ7xg3+tkhLAUmRn/109giAzroSbnALX40EviP
zer3vjNzdekdfGAiMqPZmLpYhHCHoIZ9vbs1O+QmJlqlTW/PHI+jaww58fYWbZqnUZXfmLdYeZNM
Pg84ww02osmFzg1EMAqhJ3bWU31neylOcswE/iVy7JNntZ2V4KjnulsYj0JKzfRdT+ZKPiyIMkC+
z3bmD7Eo9Tv9Nt0737/JTtAI6F5PNiIKK3fM6sP5Q442MmfipPhGrqQj7PjO3ldx2Wv2Rw6ReBQ3
DPowXN1sI1D8RbzPVBN3pqtZ4nvZ6SmFRbhs7RoOs2QXesMhwQ1d+56kECwqwDItr3C0qF499XPd
jCsCd9EpN5M33cXbKH2pfbE+Ht7d9kEiU1E+vALNDi7oxXeEIGNkkSOESxtSw89Lnb44BgazB7Op
CqgkIV2rfqCD6YqMOaf092Y55Dgj7HDJBbwjL04kRM6wodzcDSs5CEjkN4Yf/zsj/nEd+JNJS6YJ
Uw224ud+IWWJuydhwFEnv4lcmzOJv84GIhVsePJqMSbkYPkB5g48uF0ISbMOG5epw6JC5UdZzYpt
0LwPS8Q/jWJ3k73g6K3IMiUbx8HwPiD3EwIpK7yyBvNyBwKCHtUD2CQZ53+6wSjKowA2JlS+irkW
OCDyA8oI3Ur9St28ycMgSIxKAJQjMAf+NxxSg//De9ovyCJfCl/TvF1tq4l1nGKDZFAmH2gSL2R0
Jq7bYa9OllL6Gy6lF3vOAX3lgSXMLBTKDVPTPeee8VQIXRIKQD7YDVDUUgF1bYcxHoRH28NAYbgx
AVVIImMQsp2jpnqA4gs4BzUXET/KxHE73Q1B6d3NCk0gRLESEisWqXkyaBvIuy+Rd+nP0aWNrrja
B8DpUCtp+1tHt2TAeAwb0PcDSsRRwDTw8I8+eydSQxYPvuEabQ8RBSZrGbHrXigArBHg1LxTCAP0
DJ8DyOD5XU/A65wEPLcXyqtZKKLb23EgMAAncMIXXTA+gZ6bBVKqOUSYN09CEbQ9hKgq6JkDRbFI
U4w+AxWK4/79NRwSMvVeKJ34WWfTkq0YYif+dWT1YsqsXBCrH/FTm8Txy3TDlH4EW1Qiaa60ScIy
/hVCvXFnPbnSK0s0PhuKnPJWeSVloSDLeT7Smoc3YiTX50mJob2bdrAOZQFEogQGEOzZGRKDrQeD
PBSeIiBGAXHhZWX/FcwzgRPzZKBwj6FKJE/0eXXTD1zxmFyjQW8g3A9EBVdLYHIOaKjVt+ffBK5a
nV5CjYmwDdZCRMKt6oYGQ82ou7I30bxvRil+FdvqzaFoLb6Sjbx5ty10ScJlih7tXSbTdcdfULIR
ymYU1zo4sGIZBJiZR76Ng0PvcmdV95FSpMfNKsNBiuK/GU2/6Y1/nOyHDpaiwuBE8RF9OY3pgsdq
WzsU6wRGG6DbohXn91l6gBax84vI4arekU4mEarIs3X7JBs2t7pKh5E6fFTiqmrfIYnSYcWNyJZr
z+NvEdwCRZYva7L7xf+7ksk8Y6+fPk/M1eFpaZs5b8O1Kane+zlH3NZmLsQSaZ1wOi76dkQ6/o/e
HTVrhRvRHspCc/p7a3USl9VqyZWpWkAs/dgzHq/DBwjN71XyJHTnm5vDaafcAJD+P/R9L97Dd/W3
O+6cfgjRCsqYh4hqv7l+70S1MhpUj67AXJIWNWlSMPYe4Yymw+82TR9cV0xX7brXAR9B6K5oyKdB
zmIv04Ym5QULamEHrbo8e70aXqD+qdnekTlJ0UQIaMTZMIzSYrXWA45Mc8mhz0jHjApNRpwYMV9c
yz5I7AnNwwiqTi82Hn6nfD6bnttRkoUxvNF3Ho3udqqLAh2xVSu6jDXPyG7rHqP9aBPSoGXrxvkF
d8YeuFt4jxCsFHOpc1/eY2ks8CdtH2CR8xrMQipYXa5qHMmZf9iWXq1LJXSGl/s+7pAe+SjnS1mH
x75mUsIxzEdqBP5u72ZHr4fqVWoyqS6H6BwccZk8/uNv4A8Vmjcg7klSwkYjlYnaS1cu4fmW5BC0
0rLL7QDyZCShUh1CFcrZBpYZac5vIZouhxTpcmd7O+hCF4IswXEH4d7J+HuH1ZT6TYaglJxMuEb1
Pb7zqByCyNklMfSWOqce/mc/SlP+eV7VLgYZjtIHl2M1llbn3/FUc3cUeS/x26iQqSiKxDf8D67q
1c4OVHdwMixpVYIIPD8ZFNW03dtpd8ZSMbjvd/1KzAUorQYJGkF0QhMkS2M/k4i+Q938x3b7CX2b
FLQmCLhBO2dbfLgh2V6G9Rd4TIleWfBSfUxfGbz/+r4s2QVpBvaPRDpUi3YozDw0jjdRrpqWbzkO
eO/BYEZEXTd3f5HPu9fBjekyKpZhuxLu34VN/8cHMLbeHL09hOVSVmsWySEAyDrsK+fHs1m6ULTH
NCMKCW4NEgd5KV9kf6qSuuvtTfpa4Q2dbtu5KvHd/7hPQR51X34odCPe01dhP5zBeXUJ8pQdi+gW
B81BUZwPO0/p8YIg81D7KpN4z9ULsdEixc16TtOy1yXhSr4e0lXgcUMnSglCWwrK2vQZPgNY/htm
yCVw2L9hTQ+9H13M3Htky69j32z+S9g+JxBCmRJtECPJgbRzH1aFNcw3RshMzjfwA7a21UGT5Fw2
OgoxV0nDeFHzzCP1Fw5PBx0NSRF9dcKCI35+7uVZLy0CzmgsRmr607iG8kuPIypT2fY9/1yrjDX6
KZ5Sm7Wa4scoitmquw7RAnwJTMINYvm2+HbwUTJSSy8zQL7uQP7ca4gFnHqKDsDLzNoRJZqWDAuX
+XwCwSWLzrO9i8bFo8QO2cpn7X+f2dEgim94tyNZulDK76FEwYrJEqjF5Vy0PcHLrgFd0ySb42x6
SwVZKgDxMBCziGOuTKfuylFQ2PdvRrVD8fo3+hA0QLN6jKoLhVhaNCAyjNb9et4Onvdt4PsfwUMJ
kbV3pBWG8IZJjls97Gq/fVmSm+KKGwpUSeldBXV5Xe8QJ+o3GtMMJZef6EyqWt5qM1GF0i9kR6Mn
ugW5CZjiZijILH4BWPcLT89i/VSaojGslF5PE/GSO7W1VqjEKgLfol21J2URzD1TqrJlVOqLztHg
qadQt7AypNu8lPk+Urx6/Jv+mate9uYpDueYCdcB7ed0TY/UTLIU5kKRD1DBIj9NUjQuMt77zKL6
F0myV4OwZGYpi8ybxnWml8d7pWieswghL6+uE41c2ZKrSUl2uRXOU3DaFNGMQrITvDfX/m/F5fNh
AyzSxtfXmezOKnYmZq5rWLhqrsvmi+h1IwxteCaAWoboWwq1o9EpRaBMyolfgC7H3bq93/uZ4Gd0
ml7EkvZWzuJQ4JqRXt8GPxRzcctlPfAuhySnCheATclAGFWIoClBEG0j6GHAVF0T5jlws9IrULHe
nVAN5mJE3USYrwUbcmA+llqVTSF6K/6PZdl8xMRvB5c9rJaiI2nhsE8Rbay3Dfr6cJtPCi4fB3C4
6dLsLrnQ4iyZse1JXqFyNvRwT0HrYTLPa5Rem/vumQ/TnIWjA9ycdCXPy2quav6m6TpmbbrEeA/s
AoGYEM3tto5WiCifSxfS3ZmPigJSO6S7KFkbr6W5JXp4aS4sYFpMe/FVNa6lIaJw16UrPuuAxF+t
w5BTHLg2zqebHF3kPZPhDxh0EMxqIRl54MIK+Qcfwm3NDEtOnKN1DlirrxQweVR4sPpsIvfgfM/a
n3iORU5P6XPFCGwmko7hb6/MI4vqovXuSRfHkmRYKb0VK/uzFevXfOLLEDezPwwltS02K7XwDJbH
eYcazjZqgdVQ3KhVeAzlyEn3TSdq+Y6c7BM6Xbs8VgfmWN6+P9bFMjl+oRW3WWXs8XIQOOwiecKf
Kl1lofOpZpaAwyB2GcX4PULbLp+2q95kDbt4ZuspjIXKOTm97ouFzM6zDSBC6kDiLC+C4Bm7/TYU
FJ8ysyoIX1MoY3mnZsV5+PLcRUjih5ijN6xFnW3eXYomgi0f5hqIKKLnWo0a/fHA3vb4ef9aPf5f
+Go8mcKdxo4IbRvM5fbUH1HYEzOF1j6x9ZZokduUSBzY8BcwieOJRMp0PLCN+MirURuWjItKGkpI
fbNWnlpKktHqxExW0aXfUWSipDy7iwvzQy065AgVvgx2zlvAl0MJZAEtxvKJ0mb2zmdftFarehN9
OkGD/NGndop+Dq/CxJ3hkqLAyF26Jd2no1hckfS1MhFGC/cTawoe2G7EEsQ6uUzhr1U9CXZXnxS/
qLugx0e+1Hj14q92+GHpnM+RXFDRs70bd5klhUj+NTYLqoWX8FUbR58IDarqhGPNbC+6XulT+hUN
YgghWkIu6FA7z+j0gFwj3RVyBhOy/Iqv89HKwxc32JCpRjbh64RIEy2ZplS1yBzxbp7kYsjOAHSq
z9HNR+PHwI5SK3R/TQ/6387XF0gWaWH9nPgHLSfeU5SNtOQhAka2yOpikh+MDiuHajs1cPy2gWZm
5mxqX7uONAa2T4lY79zlBRTWX4l0AIc7GRqfgTuwKgPTxY5t/slvBkAgJxoXHjW1MwoKtZAiTNjc
ii31vyy9QR0MJ13ATkVDNOeUtan9KAFw2U/8OMyEuXprfv0haxZKUAM38umuWVYEMDuVnk6iii04
b0gtuLjQwwGUiCzTakf0kfQySgySbEWFyye7DDaiPM5plG8B15OSo8Pnjml9ji3TW3gAgJHfHZVZ
kUnxGzEiXvSBkTG+PHnJwCll4mtQ8F2Bb/SeqreQ36r/qnR1Bs/SNmyHAzgW0E29cAhsIfeeIE2N
H3qJuIZeFXMMM89Z4xE7S5lIbbvtlKYpnQSFzYfaI8awKB5modqguhV4+aVYXwzLwkUhFon5k7et
iTKFsDaq4p3/QJiRFcTxV563jKF99M2/KwIuYRWtla6SakIMWThCw04nZzwsxa4V+QPg/Akc/nhG
hDs3IFL6xakMv7CkRjP0CSOkGuL2F9t2FRJZSVyQNRHkZ9lsD1EJ2AQzlwLtQU0h4S4VqgvvQEsY
tLoWJbRIjAQaBmSPT7mpU42HXNeVMc30o8u9VrcBEo4GcOtudIbLH36bRjLj3epTVEUzr5o4pKrQ
4jJndacxTCmOqwmMBcxOOUt/bvVFN0ubypUWRpO2nGck9CwoRVKeHZnD4a3IATFQpSMU8l9kM8cE
+8YSRaKZ27NN2FYkJE1EnPyvsvd4XApJln+dACX2wGYMGNdjKv48akocaH6baO9gL5BM1dce13Yj
3kLBLN7ksLNbJ/ZdAvsyMYWCCYk9StDG6b1BJXThUZT4uE2lxFTbQzvW9iRg77i3OcWRqCigLOJ5
8uh896/BGnydiPiSBYPWIhf/bYNsoBExvPA/CGCsX4ckEaN+BjfPPZFyl3nO/g1Ruv5LUAH3moXc
Rz4pEvD7FfZGCs4CzPZo+Neq+uTz35H7qVarFAV9rbmmOlRzx7ivEgQyqprDqDQ4A4pBYVP3XTzf
+sINTHlBdadKkL1her6VMoAic/SzNwI3f2vBI1mVT5J1dBG/Uxo4yhvn1jIyYuiPrwAWZgSSPyxI
3NliXCEZ3mkebOP/FoZUi+nlvcHM70HVpQXSd3qPW75ncjH9vA65bpHZz1Fixeq1VqeBV+vbtJXx
YRYwh7oVkJP10dSUmepILaDRWmH26v0N/q/s/D8X3+uI09SoMyVcgTnahkvEIi/YTsn3jVgTBaZA
H7TDDhAgF747U3YRkzCvTAgP6VHqxuVsHKFf3QtPolil8tN5NyeEn5qAvnOVtGbBwfnaxNDDHhXP
VC9QjsWsC+nolbKoXmc+i8xU63tkLPgW6r+CIZR2uoHkpNDFTLIv+INKlL1UtHjNGM7RhDVUWvuK
kSxEq8MmSnn80T2Wlt0GYo/mbk4VDjt8ys8vI8nvvgEZPyh526qGpZVEgshchi84cWAjY90JwiL2
Y0MwiMi/ZLksNEYgV39YRUScZdXz/IXpQLJ0Ye8Stl+a4kRJYVkdGWRzpc2SuYP041+KapDUPdZN
4yj7ihwcTIuEWxI4HPFHc0wxuyMCn/eRrzMKvQ9rQwGuUOWcsDdyiGcFzEqMui/E5QSeFqtokRLe
EGnrzyP3ecFDjLNw114dm68BsQK+p/qDh3hLLpeum3oZjOw+rsPFojrU3YOWUP6NjbvxCE0IwNG7
YjU552xtHMvRjS551rJ8ir2N0oo+kRPp5NgSeFdfCR39i++lp9M331lpPeRxpwvy2KxqUgZuSipn
cItjAXZ0OHZOm45WnWqYqmQ7A2H7Dwwx0fHPoW7qJgpajDoiI7fvws/H4AZ8wSzXoFtrBiD94zeY
/k+Cm1iXdNHrX3bb5dwSM/MD7yNGPJqufEPSxCkVwasmDRyvBP0k6q1/q4DT4oI4eEntKR8WEkca
9oUdkERYpyeJG2Ke2FUh8EgSqpAszTcSoOK51STh1a39KQXHS90V2yl1EkAHnwEwqT7gPTrcJQN2
9Wxv4SlMSYJipyrLDXOSO9FaHfUR8hsR6L5ZzQgF3mB0cgW/Kua1sYzZJrPevEn0S274lujgFRrC
TQVwUR0Iir4f6/GOkfpJYR5eLp8ph6DqgYm+uCs6P7rBEiCj9zstvlVpS5IijC8h0sq4spRyFvcB
/QZVXvzAm6PMx5h5dHg+hQycPARsT81fgyGM/eBhtyq9MRMCaz7W5Xn/whjiqEPzUwS1od767uwr
cqiPkB/GMSxi9NUYr8Qt/DoY873E43ORJ83hX7qzj0B6V9Njszt8uj9aBm75V5HosW1bClCazGB8
QyPLmLK8d6gd9u1Yfj0EMGp3oQZfqajcUhc97xreNqUdcYLfDqbdQ5bnSkL0zBV3qS7r+IrMXrKk
FirK8g9ckNlPYWCXJTfKg7GhaSJ86fNI6K/H614pifdz4U5kDdzTW0AXhNqxBNDtX8V50HujJk0l
aAXMXXYP+S+EGCN7i8iP6kK2DVDlJ00wsVS1tNtFnhAEuFb7UXJk4BMVb98s4KJE8EebuYLZaLf0
YLE43GZnzZWnW43WBc9AzMKHBGvO1IKCGEzgd/Y2A/Q/Xbqu9ijH01uPKmvq7+Uq0FKOSRxlvo3d
Fb46U0uIf78feqQcIJ4QLC7CnMifaDQk/POvnYZ0bD2NBgtgpONRznDCQmX0ehgLNhORHBlI8i1f
OCom/PzH4tLl/qjmywSVivUQTzVomqV8dH+c/ykIDZXzHuOWEUo0Gh/pIsKcgNwzHmjVSxc/09Eh
fqNAR06LLqqZaADJtLxgEzZYHxhXNJUAGt6q8S77oisVyuZ2GaZgtgJasRm9i1cBZqV8HYGrQw51
EnAA6DC6i6XR8myDbCKbbuSpsQRtSBU4xu4vGRr7W6uF+FaaOhjqBAwjaMWn1k1nJcyua7CsHFZj
h2R1OZD9wUuOLqSSOQamEh10QPFl8H+uKGXtTej/6lmRQWE7MH+pqAGlbc9CR5Nby6psISp7blEy
ExLLroU9nilH8BN9EFl6sJWQkCuocdbUCkT1L8a1encCSgLRqGwkXcWX8jf+XggiDZ52NJYJjaav
bwDjy5wccWgdgoJde0djMzg7GDccPF27HkuGBYGQEohD9yl+RwLiuVPx7GAS+cdqlsC1qIj9msZg
kRJhgkg6O7hv5lTAf+JIs+6FaD5D5rtUlCH9WK2/yc1AwEC9g2k9KNRbt5iFHJeIl6dYwitDUU5/
82sKPhcyJPD85ccIErmRBet2L1GE9c5ZvyjGtylQYL3Nh/BoOZ81fwXoqE1hPwIutcU16pd7aBY9
iJy1sTeJvZfBdiBtw6mA7ZCL4zpUl8B3Xp5tFvfaz34fHkbKQJsnWYxj63wCRzgyS4F3XCLeXLu7
R/w2JzNV0gf5XD05oowKC2A2QxP60FQO5bGnrlRa9EwVA+dkwvpjD23wqp2PCkZDX8QePZAJ7m98
AkogbYZ08IErNO8Bt1q9jNxYHDdL2RBM+tYr97qj7aks2Bm1oaKcn6tYheSdYIlSYK26hSjMdmaw
L74RbDUAJ9XZxOPA2EDM9JaftMNylBNWxWIPFUnJz1QIeWjUzEZ8fmGrAMK4RqM4Djsj6yfiUyeq
vsL4TTt/UVLbYd51Vf/onnEjZCL8+eny8uzU1DRjS/trA4mT1eYDUn65CIEANXZcGEOBEVjoi1CM
alioTQ33HcCepW/dnLATH6l3nYlMNuwn8++cEbeRRhyVH5OLlPP+lUs/HRdL4BPJLMQonZt5yRfI
2Lp3exxzxezGvqNlXCMvO+LRw9lAIHpTCFdODF0PzVRTsnIIrYqJAawDuoIRmTrheE5LVrOLiOS+
ZUyvPdZ1KgqS8JnibBwWenad3PZaF9SZjSDZ9EUmSvOXTojxfLLZgPaBljddjVgIy62HP7QYt8hb
QeZKyhVpMksn9RDefNr5AwkAXUjJsijxY7y7Nt5JMx3ghLTbKecmtKtBjc/3hxS30tlruNBx3Qka
6VLH2G7aAroCGPu1BiihT1vqDVvKixxVLjVYixqrTLcY3lIwu36H3X9pR1lZkOY7yFFV/vKe1pt7
GLIq6Fw6XPhvwxs4oP6ZDOogpvG203/FfdLCeCwBMOlFBjJplTHixVuDfI0a6o1NJlqddlI/RuhN
LnJRvyoONXwHkL9fCcJuBdmITzZi6BKt50QO/rrOZ32LOSOozAyC+Uf7sy2rvebzVfy/wWJ9eD+a
RA0SvpoZ3xxvLndAps8B0jDvmiOT79ZJsZFlO1JpnwemYjpOyuC9ZhFukhwrwkbeXSM28+HPy9ZB
cEaFmS4W8fDtlI2u3GJV7TtPqjuX+6vFxjRdatpLbbbfiu6iKTy3FzgbL2lDQiD/09T+n2ZDaNRX
8niRRtADKDPYn7vrQSqevi2UYK2x12MJVJF/5UR7lOM3ZnOSN/nltItQAoSpsWHo3Q+wLVJs2Mzg
rsmXmIsEkGX8dzHs1Pa5E2CXSF5n4OvazzzMIGjrev6R5K8u3RSKwS927FJpX9/hIpCayN1806JO
a1N8hRlGT0hsBD2mUN9/FCUdDlmuxzfDk9dekBjraXveAcnZy9HsaSJS4SmUHhgasO9sN1l5TfPG
SWYLK27fSW+Jzc+Pwb/ccXpx7pv2Gd3NodPZykBuQf/H/8AnEcvlQrdBVQ/fF3nv2j31Ya/46CB2
BfqGcGHgL/vKYL3Jhn1x6qs8vd4V5JjtVS4W8zCrreemSCmZKoBM1OjlEW22SjXPPgivCI/0qEnn
1nlGOZUiEUzz5/Ua4oPH6IRGvyemNBq/9xhVv1SGRDH3bxxz35B8bbsyph98J5fn8oJayThR/+is
7SD0g7OAggm7hi0GfLCWq+TAgpxyLRAfWqzmK1+QCLfQhPCoA2gbH+6FEE9MWN2YVj3/udTMBL9U
N/X2odiFUcgOX367vwEeOWnxNPI/1mY2I8NGiYHfScg9B/cjB/8fI2IlH6iWMUbC/fwUy4RuZh7z
bW1Kmphj0Hqc7TTNEFuVTqqqkbwc+/q3n7dUn/I9yAAGnF3c9orhsG3SeJxdWyOqcKKWB6Njqggo
lId7I81bu8TamiJMfv59cuPztJdLLKS0mEpqZ9evWORn28U8R5Vwcu5FAw0leI0Iqdwo+zjNPx2i
IFn1ekHjmMKt1eBjFn5z/3j3BL2cq5rNIoT/rboRnK6S0DDxtkEUXxEcm8kFQw7q9AAMHFyav3Lp
m8dBk3CGd7MKnGE9fN39RJRgsc5s2UbOHpLY0TQ1XYRwkjaA0DRVKExZIOUPBPi9UWpmHBctfz0s
803h6VtBryND2nTmYp1tYm6ctIrzQQRl0xcYI1DLE7uxMrlUzOkc5lBHKMeq+67AvJ9Oe1nR308X
WF5al/b/K1805pHtatDVMDQkdzHjZX1vAg1k5FmYnzdDUaFWcr8S3gE7WHwGsXNQcQkI2OBX2tpg
NgLBHNLZFpQ4GOWXfLaihG7ku2LuwKuwux+Fv7EKFTp1y7oihE6qZ42PGNnHGp4ZrobjH8eCZdgj
zvJcioidcxdCUfpxKOWllyc24HWFz68N3VfK9Y+bE8tq6Dbf6TX1sX30rKJGJUzewEY8g/nrB/Fe
Lbd883ipoG+k6fKQ+RuW3cME+K5iM7mrK+BvE5xeVc/QY89Uc9nf4PYFY/ecmF0WR2d2MI2Rq4Wu
kwf8eezVT/ed+q3Bw8QQmgWhjIaudyHyrd3lRL8MdrTyZvCyu0XuYarb4cp7u51PoIx+zl9JpkrD
pBTYKxuo0/CTciQY7zwgWhj1PAdIx+w18QF1srwuC8BBgfPdxEE1bsNU4PXBcs/9tbBsCuRMgWdi
Df23I1pM4B8wnoYoc8TlLSsC5p67JtHT1w168rrD998FEulrqpHTVVFGB3PFrFaURWzejP8OHcq8
P9RrllBKWb+datbOEGWs+Cs5OpzutOmPjAHP2QxxP/5yOTX20NornYCqKfhp1E4Amm2sCU9IrgKL
+NwAaSyiI6FeDy1JcCF22FOsqyxzc2ya/Ry0WBbWqRcqdWhq9qTEBXRrp33PoJcfG3c7POHNaaXV
GsSkKTGOV4m4edm0Kz1HjDCpaY9bS+vxYyeobZmDIxuuyrjVRgYdvT//o+9efJrUZNrTmOdn5/aG
JBV2k03o/aRlijh4GT/koMdPpjIoOOBvSjxbXSZdLEqDSRM+jF+vIdE+mZ2z5MnZG2i7Xzf89k0v
u8MjvSoZI6PppuH1OAaqLgAgWrELHNX3nkdayJ9FoolvN9pzfYbQrATcS5T+O6l/AzfMXnqVEPhZ
Cfrsv9tUy5vdLqrmjcUTXJzeIs7sMjDAodZ1gaFL2laFgXBeXFMl+TY3vkPgvM+8/3uRMJE3BLmF
oY7YIlbpXwrSYeaMjc+LnEv7+uJsOUR40vvPnw3jCZUksKcI78fC17d6SJxTndgoh4bdCZA6h0Kh
Da/pBAlI3dfzZNAU2PDtDab5DcLQV8flBq1Q/EN3fBj+aZyvGX0Mkjr78DSxf4fje5LwtrtoAU0s
l10RBlPXK4Lu4G8l3NiLQ080ZKWK/nPwhk87AHW37M7BYWNG2GSQOpFSTphgrxmdha38uGp42pwT
Pp4zITLf16mYhTl2+tJzjF+ChxKCUi0xznK8bx32AmYOQbccwFhSQDnsJUDECTYlzuHGqReAqzII
F3cB9swTjwXGG3hHPoCGYVd73V0iHJVflFE7OWqtHcI13b5jUNO/OL2+SntZbtD3zgS7U4U3VFFR
LR032qR+PQWuVhLIu+jEDZQYP+6Pa9ESc8nDSRnpKBgCuPmKaWGkQEfPDl3C/5PIIrbTXecyALsk
Idu2di47bVBM4DN87gvdthsN+Xd38ob7G8FeZ6qTtO/445C0HjETNk+uivMyFEONIaeyJX1tkgMj
znZ6gC1VKDtFzV8kwBgMSfEiX7qlII1PSnZD/nYy/mXhv3nNKFWL2Aw7m+rIUOKbnJv1JGyQvrcV
ltveiyNSCWAD72VN1UUZ554l4+HJ6Y6wzd7O8Sttyn9538gDZ8XLoIAFGauDbf35MxbEfoyP5bjE
iWRuo13eBtHxyjaK6/RPdp3Iluy/sN4kHqQA5I/eJldH41LAXIAwKn6dJ27M7z9F4YRYBofet6vm
uU3eRR5GjOoxcErUjlnXjMvMYEYOgbCZh5w9940pnMb8nkicciExJsczQJDBwbg2RkZb+96weXSc
EHvmZuqWMKWzmXx8N//7nJVsxfIwO5iH0DZTkKh72B5Q4fFx2BppVvnaoMzAiSrnTK/HVrhMvHy3
rgK7CNOFPZ0Nmz2Y4FPGblGBS8f7lz5YKvyID13gmKcEsG1MwKOlqzI5uECIfdz0UuSHikDv31aB
T2E0loPEDg1irD4l48tyzu5/4ojE5eslU3r8RYYMOrgoetqfoq4NCSVrGcwATcAGQwtSTzjCeSTb
S2NtGWxxct6UfKkZ0Namir3J42fhH0tJoJLaEIUecEIeGWvyHr737MqBGUa2Ox5oQa/3/kfl20dM
e8RODDnIc3K92GfMoSTLti9ej3nvxaS+mz5jkC/cSwzmRfJeOeHkMoFfVFsLuX2wMcQU/Ph2+nPx
ay9DgL5zHL8sTnqUJBqtQXWX6iq7yb+OTzQZ4Jvk8WA1T3/8/J4boRdhYYWnsHNx1eaB40fojcNY
gNvGfgP/GdKVsteMFvl00K21Jzd138tHQIEdvvjn6ZZobVPZwtlmXR8fBYnnAjdxY+0C8SbPXXUh
P63qJxVdu7ePb7JDMVrYYvSTNau5kYunaYkvUMoZ503ElxDxNq17o58Tpu9tNRB/nRKHJaI5DSBq
uNkw3ttNQSmQOwpOrho2K6BF+Fa5kb7GRxDTWw5pqf/B5ALTj4P/7uC00hE4g9dtYxmY5VfdapsU
o2SgRLXtv67TBVhVMeTwP1Jm0F7pE3Lm5Xiznq9XE8CsnqVQo/AcpQdJn1w+Ttza0t8GWmACBYH9
PTb1zhgtrw6r2W0KwBuPXrJRkf2lrYjNoL/4AgerqipOlV1zFQJQQMDKKJyrqodUWIAsFvnXyuft
FeladYKJshrmPd9vgW4OqA6lqGHmxDI13231td1YHdc6AZKsSfLi9fqk7qI7QMeM84gfz8LT41Mp
n4zfyXhwjMT98s1m2GlM7XdggNwdjmdhgsNrx5qk/Sb7wIijd90XyEOyJMu+CtwnIB90EN9cLih4
r62nSpK4tmkc1w39wxFElosVhMwW/jgeHXs6xNCc1fsaiFLZZa8Oc9qDY5CU7HGf4AoOVq3XtPyx
SeszR4DAU49yt9i6bmngm2miFJmfzwP0fAEZz1GCxNsxee26poJOOqfxAyxnWCRT+Gh83t3PLajb
I3Yf0BgmLQy63ei4Mm63GgGYbbppcQiFPhOMJ2dOO/1HKdMe460DVZttDSYFY2hK55jtYQw/xWWp
plDtCGMOsF/W77jn5rAPugjFAeplMHK3KRVcApeETzy848WaXZN2zU8S6vW8Pm96IfyppnfljbIa
zDvCu6csTwa/ENj7EyPVcF40roLcLSX/FNlCBqi6JCKC3cYPXNMbuQPmnb8gCLxD8ZLwtZgI64Br
uTWDkOhxNrrftYL1WoDVDuFtskJAaIa5A5Ry9w9jWGFh8NYY0PcO861t0ktMLPu+xAMIdpdP14xL
Ikxkrulay69AeG19+1MezrIyTxN6j5Q94YbOk7UA7e4ySLr+kI1LHJAKii1o1/7o+Xm9ogMbcTwJ
Jdccv6iw0qvpo6Ks3NNJY+zy9mjS0wemy9PUzFN4h10UxA/SzqBAzDCzcFKmhND+HZpUAf9rBDDj
izZJrjbrIQ3Rm0d6CX6xGVI2+dc624aM9UPjAkRNzkgveabPkRGqRM0997bIbBex6d6nX4UdMTa+
8UKYCFWjMc/dJTiB5FvaFz5x0ulkqJB88zOO14mzfOvifklhEzLZOXGUR3iULT01RJVVRlXjAEwi
ZFdQOBfzIvnGD7q87MLKufidQy8tX2vFAOA/Ya2m2chE7/zgQB3cLFrAZ9h2N8ZenSQsVL91FExm
Ry/SMD/I0/SENB3DUSfYLoTm221lG+n0353SPwD7+3hDRNCX3EgpYZKK7JpJQah67OrGWyWJseUa
2sh26M/RITOg473lro2gVlFV6cgiVT9M7WEpnX44JZH09s42io1Z3HOLnKDRfYxh8BskvDx5/NEJ
kQfx/nrMpM8agm9ueZVPCSWjbIDIuhgXvm5zGYdvO9J3+BXz82Q5sqDBohMXXEDBX18tyBqxc0te
iRkcDYz7xJto0y5DX3/fdMV/6tpX2xDEYsSTRFcW20hBHX4YkX4D4Go7qWSdqqFZ80cUmfMuXSAn
IzBB2viDbqJpn48oSHadwgJBOwMKqsYBU3ROQfLH4Ziz0R3KL5pYJGTn/ghP08sDX1ENiJyC/Fqr
jS2OOB8tUpM93U6ikwEkkhkmrbuBySG77vIECyb3EfBJylfiGPLc8uQc4BQBR94fMjyurZF+lq7Y
kqMB9z2tKEyy9aWczfNx3PMcr924qKMhImUINErv7RI/l1odprKMf+ejtf1QEtIBvHGcElEKf+sj
nL2NE20JRCzySr0aXHxinFpihAdUcrET00j3y8CrRPbSmRBK+6IHSr5MCoEXg8n2z8noV/Ly23wj
1qeshu9A2VmIG50rlaJjpfcxalPQNO1mge1qrQwaWf1x1WeqSSFeVRejCyIu0VbIS0WtFklx93A2
4JqfQTo5ZkriKuU6MrodTs5TuJyu2RdRzN3C1q6BNO+q3FAEppiLxG8TVchgYm+vqLGn205wChXi
nEi9bxObBcZdzS1rspLq07zsrhYgMVDoUskYKg99tzXUhRBVaHT/6+++W4esXkOiR4mvSX6qHFCn
eZnDtWV4OpD9j3zjXAXDBSU+938iLeVi4Wuav1PXTDBwtigO8zDOnVdArBAcrISIfUAapS7SnXXV
OaQDGIHfETawJotHBDuCL4grAMNtUSXF3HaFJQ6lz3Va105zeCXnSgUeU+N+tYPcJhOcSptYyPKM
uFuZz7n8a2CN+BTe7BnDnyMFMPJ0QBqMzZsbLnwHgQJ/eZG2hfDfKewmbLYd+FfGhAqsVpPkaFZX
QCYgvDiP5yhVqel/l6O50wRXdEiCM6irRFI67/9pQMmKMUA9BKP3H3qA5v6S+x2URQxp0KgC0VYM
1teaiIbjPCsHMXLUapJFlaWJOgXl1aISurdPGzoZPddZ6nZRyDYGDVEkrFhFxpSgb+BOujXFtZUF
kaj5zlO4DuYW5XIkmlMb3FPbusfNe/zW8nG+p3k5FpMHc/V1nUymRpvdKDQWEpk9NN24PVGVFCEY
nbL3M0aCXKzuvimmNXWiTyMAUeJSyAECo85Skidi49XYiRzEwczEzrQZ1E5vUJwZH7tby8H6++P7
0vzOnOALIW5bpYOimeK1ZHPkMxEEh+w5qBR+fxHDXuOiww0HxzPlp7ompJ2/zzY487W9YXfwh0mI
qnXBMgA1Hx/oGSoGb06Xo8Mr5bFSU4YO4bjBw0jpHi42CpEMDTnd54aUh0gHAiu5ogPYXpjUGzK1
3HF1ERWX2LE0AJ0dzrQZDi5jD0/fWU9Swo7HzHynOMHD8I7Zv8soaUPXICAPgn+5LobVF0+uqWK2
/cU2Ct8RyDfLXIq4H+O/rYD7/P8gRlXlpJQghpuNui7bbV50mlgEE2iMbv/YH2fqxAMj68x+tcVp
YE8F8pPZ1f1gMminOqLCxDk6jGElhXk5BzUrtNCdh1RxSu1ulaSxLm6/gxpiXECukywZpq97yYr5
1+zip8sd9wQe/QuBSgTgSojKqpARMZE5Wh4UuoSSdEUMM0BxZd3Alp3/2+UL3q0EyE14beKScB4e
uPcPS1LaIYYNCzrHesh+mIHO8fBeGbiMT1F5O8ChAK+m/F24/LPNqppfSP0Ir7VCJtmnGFZHIj3m
Gcx57v4xMJHlo68T14kCUe9hNdLi0+vScnzR1pVGDsanvLhw3tVB2LCEcVaH/CaR9A8qJRO6M7No
OdQ8ALDuZsoWfL7qZ70ESbQ6avTEJZMW0964YNIVYuLZLqpaLC/2wpbhP6zi8ory1jOQBTsthZZC
ULGmg8xgpXYYF9EJ4LFFPYvR+PF8ZUGZrrhUXNlBp4l6Tayg67firHsBwcr2vjUS2+hWC7cgcIQi
dBLkCEWzNFf63k9hh360knGm+w21vXAwfLE4Vgxu0B83JhBPu+IECOri20d3mqE93z/NvB5Du1AJ
9hgHN9f9a4+9wFovTJLe5BrXRIp80WApMOBLCzsMJ4va+CgOgZT2YqxUQTx2aN0f7QnzgXmqDNl5
s7oYR6Rv1OPFQkuG9pjJs7VUa/+eyp1eoW3B01RM30SN+6lWC6JcCZpCK5J40w+wALZI2ZTG25NY
m9aJGUO/HCDpGd9tfDnXt58aSW1n77w4O5JknYAsH5BzgxNc+rxp5CbeaT89xpiZDzi6SicB86VD
PTRmjGvFykbDE62bLJCsyNXs0HSC8z3wPMqhmAbC3JuitEXCzXPpUjKoAGGfXhXD5vmyvxvH08ee
WMKDMRHgIpZb3omNBV4F2r/TYjubno6UddeQu4cPOx7Dw7k1T9tEHDN6YCsQZk8fRgARAJwtZ+z6
y2KFnjbNezg2srCikP+D6t0oqjJwPklxsufP6Z7CdIojlzxtYA3aLHv56WT3EUtfnnwNMDm3tpTj
z/WkWtktgv94vewFxpfg68uueogectm0n3KYxIKgoScv/YJdxH5QWfhszcCc87XHOVDpnDe1rt2u
DkGa/bIij/H4uqRImMQ9RIR70YPcAO7P5Qv4u4/vexJri5NQ35npCpmHZqfRltUpfDFnaeSDpO4T
81SlJc1D1Pa4URJNBs/GxB/yJTeCgJOJ0OpsXue32Gaphiu95Amc1ZNpkjJPi2BC+XIFRxN3u3jw
fBc9Lq9i6WGY4B7bQuGb1+XiyjOH0k9xmNgseuOX+BFQT6pK5lQz3SpNcJno54cM89uDD32ZPVY0
ycurzJbFzDvu/P+QNf1paWEURa+ep6lOC0C1BIb9ytDFHvl5QsQfArtr8KnmGWYuLowqDTbOkRim
PRCMyf1JlJyhAjzGcobvtR4eg54tNQHogS1HZJAxI8OU3str5j+xRsDFaFhrF/R4moHkUCzoNoel
v7twvFWoieLwnqdLO4YTgahjmstodaYCYC3pfbNbnuNUe5m2Sgpv3yXEvyCzbDTccijzN9E3SRDx
Bcfglbn49Y2paWz0tQxX0/XpZF+hnRncZL0HqLrIqJE251oOH2pahi4T7HN2PYHVYD27hqrIHlMa
cnfUFdK16TLrPci2VcO3YvGv3RetQRD4WomdemdanRl+v/oLgzbMKXnCNJx1i9cWea5HvACOppIY
HWE7sRiE6/34dNaouh64WJYjMXYFU0wptbnu/D/wny9QyxyQxgQlfGavO0ZLl0ZrrV+Szh0K/sl7
9XWCvrwDjNaFr485w5kbT2EXgAD5ZW1KPFuW4AGXLahyDYDvXYZQ+LmId35SK0BgwLcRhbnc7ueg
rpNyH+q4uQ+RQjO1BL1BpTywm9ZCea0MV3+/jt0UPCdtB0uHq7RZCItCuFia1WzAucOAnacx3sSj
s9fryDSvg7aRZpv4jToO4xKVFWKjW2rhm11e4pPybg6TdimsSaqBwlypzPKhBmEECdFGGyySM3fd
JzLoIM42I2AK/XERHdcCIdENqRpv4/d4LtMDSHNAtXtAksmT/B8ukawlnJU1NiQbyLDwcNHyEdRM
JBQ8FB3oRLxX8kTfoDrO5Asa8f0chc+Hb157LJq3xKqMZTnNEY2QgJGojVgU2DXTa0SwWWWAr8KC
2ROUo21H0UUIa1Ak5xHm/9MTzR01VuALIEsF5N7LbIu/g3h+AznNBl1Zwr+ollML1tV2LOQrAVjL
QJQxgKTevDkSMYOj7WlSzDqVIeTJ7B0iJjRZCrE9b6kTCGs02GqOs6O76Njy0m8/ryTgTwCGAbia
NGge2zu4NIuFI1WotZnASfIGgjk2gQBmiEU+moo313oJrrdS+V25lh+VBz+QWFoMyq4+LTVrHJ/e
hO4DGFQ1RiUeH2UYdsFl8gEOkcB3FpLNuAKPamtiXivUTP0X3eqcOMk9GhaAbFOjBfGzz7zadN8r
vKDGMPeiDGF13Uwdb8K8Lw5heA3SIs8U3pFajsKg5Z4fY+HRw1u8VNFgthl6FAbAQNxLN4SYpSpl
oFr9I0sR/lebfvszHViBdqrz6HOqVDDU1golewztpadanstP6E9cEZVyu1oF6gpUsspUr+1icumL
230AvhV2k5VS7FuNzaCTiboZJ+pOevlscz564sVjUrqSEmMETGTbMKGQ+bhSpObkJJWMwaXJgacf
g5iMn/aLQsIdkZ2F+Qq95CQxfGEz/iwTuNyKhxwk5AxgM0xN4MyxLmkcGbEKvx9STWvDJFuZqnwO
e0bnOBs55GFDxZvApxrihC1NnM9azHbJUQ5oGFaIv9qf3Qu0bzBp2nP4NrF65ypg5R3tIW4Brzsq
i97snKWvQDDU0e7T+DnJDKg/rx5tDMEUPg6KJmXWzxitP4X8Sv1JjZ5L6ZqSNz8WhtNLR7BtPJt2
H1Tcw1D9gL5mXAePdQpiYQmt+l2mzsyXasEt7HSHuU/urKM0/+P3PBWHvlNfxvDpFBN5R41r3+ii
hqmMcM4WKD8745NxXnA2qocUijHleObmFN+oypImTo3NM76OycCKMHgs+Iu7GI9DaeBBLJ5mJl40
ZR2jzAarBXI9wXi+vAOZ37os7miWqAUySVGcRfeAWCE7ezYYnOvKoNdETiAkEQyE83oQoz8Qeie7
JLzUtrLCFfQZbumLYpDYsqfmtXJNWNgz3MV3zUja80J2YzZLAz5q2BjBoaLSjF0JMuuKyyY7cQAS
liWB6f0CUFgbuOW9VtwAV6ItHxuVpaftI3RfyXoITWW5kRoYPZVIxrxsngnRNCuzKD9vxnNjLInC
Yll27Ja+P4VFPSsXZtoJk0RwNQ+ZyrZDhNmRgjvSRk6W3w5tXgIv3p5tHBF5JncoxHnhjE+B6olf
FMZT6UiQcqQ3eIoozdFQcnocnaJDihiej4HGom9Ns/458Ze7X7Vd3tMuyAW3VV2mwinX7Yg7To3z
w4iLCu60pFqJxcwNv6EppYDP4nCcr0GkYIOMxi8pi81eE90YoNCTgbBigXDXvkwuwHI35epQPYMz
A5+y/vgtTsXg0FV8zM+4wpV2Q5eJZmMFbLiHgm1RXvXVuUhw04yi6RhHvNem2sMVdyPM4X8iyb1K
sAqqRpPv1ClyCN42EMjjgxBtdn6qbmffizzsQHYwQ6s7l9h90tHpRt8W2h4sX6/IWPq2obz/epMU
CGqN+DuBS/fI1aafZ+xjPJrR9FuLr6tg4noogho5vttLtnxv+th5MQuOj9dzE3n9cKtggkKeXcae
NSZPF40y6ge3bLANtAlOeh+OZsbnzhFlCPpkY1AnKn+YlecLx5orAlLKHF+kuiEzuNIMgmuktinG
0sGZjIZnzwoiC7lkqokjDVWTUkaScTh0vTTXQbTIqaQn4WWWLJLu14JbjyhhMpN0rSzSFGsYuBaG
9hcvD/dKyFagQpatU8wSezr6TT7cmZwvXOwTcSDey50m3jfLjoUzmdntmhOqtJvAr9xo/7T1eyZf
K6uy3sO1S7I/pTsEwy1eBec4dA/YmWfKgvdu/6R36ktKyqunFktWXIWupTC0WKEJM1ZTkSddXtdW
CMQqn8mQopxEl/DGcSc1eNGDbiY1EkHYHzVwWnhRTgUUXTgJKQuUXtNqSZvJ4xmbmAomn9HAqQTL
zaXb8+rcSEXpED3mOetr6IK89IVBzkvDRCwb4RdI4tL8XB4+UEUDr5QEyjxVKwsELbWqsP3XD6cF
DivbphVIHF2c951XQZ2X8uhjfMCxKl33Vk3BZZZxWzDEEd8euRetsTSYX2WWcue+45A/TR+iFkK0
NaS/y9rkq5D88BnzojPpZEyG1PzaKQDY+8WHPSbwhkA2Au9mUmbofyGi4YqOGiERd7g0r1vbzyAj
E0HZ3kU8vmrZ3eLV61MMDgBbQC00CVbBlgo5te9m8DrNfqXvj3zuyMgUEpC6FuzJP19YSVXkpzvB
P3birSfujQRoeOOIswr+BrQk2M3c/tBmptk01e5xzU6ang9EHIWfQODb1J/J+hLmkvQSBOvS9RU/
zFIulgoxz+efYwKgHNxckHo66CTaM446EDvGMOhWZ7XJ9inIKZ8P4XwZYGHh2Befuoh33j/QztEN
5+riC5c5A+hF9G2ukalxCItJQnmTsQt4Pg7gvuX1o0TqePPnJtm6Pg/9bSvV8A0S9m22tixoRwRf
MhZyPBFmqWHmWPYBIHRrCXIYTsSNaTczKxhOWEb3L/qif+w0aromVcWQ2B/ECPAWEuVedaoP5eNv
Ajolqns56v2x7OPjv0rDDiHUhIl1Y+mt1xc5oX+PxCwY1e2bOvAK+d/f3l0c3WnWiHhEyM/7C2P/
PcmHJKOFuctGuI9zn7BqyZF+NQF4HwcxwM6XIhuan0WfCwGamz8lTBZFn9TejNKhr8Bhapu7Kgvk
PxO9OluqUASrbAyHCPuXX4OaxBr0/0zM6CsgF+LmkLYGGYCwaSuVQ+qsm2awPtxMJNcXqmZU/drq
z/q879YWpslPaRxl7EtTu8mvN3mRH7MEseSibnrcKukYY0ycdtevSuDiywuaREc1stmgD4ut6QPv
ObkIomEiKFye7X8rRL7RoYFypU15cKUfzzch557wWgUbzRHY+mkDeFRqWDtVRNkmBaDXfI7GHNH8
28DSQ4uIwzbG3SVTJ8gzbnKfkHUc79B720VmXBLWU2WYLeBc7O1Fo7uGwomA6ydcooyiiWW8djwJ
fEX7Z1ZfeDqKwyeZHmgjni1dkWPE/TN06wvSi+aBfgneY+0MheeHJ8lLOvGhTsbKeG1g9JyRlTSQ
ov1bvBXX8+UT0CDStu1IrOSWfn40VDsnpyGxrPUGKoOGIjrfhvY61eJYXZ+YqksvSEhULu3/KEqy
moy+IzsO5IB+rXdA50zmeIlDh0aZd2WDdu8fSPy3PxqYc9aXJkCcVCsOdi3r+suOR85uLm7Aiz4P
MVZc4CkHCJKCg6pfftgyetupFqDkiMDWod59nXXy9BMmA/dgEAKwPmpytayfvOZ3EG/PU8Ki6Ols
Z8pVGDds+LL0mZfbVOOuIH/8rRvWhLjSnr+5NNvVbZYr7vo/5xrVzJGsl4lXIEtscP60nr+JF1ks
Aq44+5v0kmsHrXQtQRSggUN4H1d359O0EdeE50g/NWtaTADYKfPRkcEj3c1eP/oYNvxITe1s/xyo
J1VhDgn05itKRP5AdW7iL961mmMcK5RWkv5LBEo1wRzovchoB/+jWadRHKm8q287nG6T0Y0su+yw
BoT6cvLvz2xPUoWnyaToXzMrfpl29hpVJCPclmJgIZvM50ltHKgnYsbCyZ1x3zJ4FwDJhKC+wAuR
Fl16DkP0azer7L7cHKWhL+md/u97NRUROKXcBR00AWJqfMlS5xqJdNcQhqQMk/MICujwgyhq5nJc
ULdcPvXzwqoIp9bjrw7yIXnSDrecvF8eNfYgoivcHeeu2wlgYLU2wSAIXH00sj8z/gTRZ1maKeWk
PgN5CjpSUOMqZa3tOLgDCrhkD8rjYFU/vXUH5/pNH98TzvxFaJaLZKc/cRhN4xdFxTjOqj+50Msd
vCLAIDgS6Gkw4W1euwwjq2hDMIhQOiLmS0Q6Ue1BVfCFrkLDzsX81TzYG3N0Mlje5qGGcosVKmlJ
egy5jc8bFzXxCsXgo7FlRuO8wBdOm8btnpGzYhJIfgHeGC1V8rj0ATcQ0Xsb4BaeOnk67AQ2S4Zn
aoBXHeCSjR2+6yUpkqt6X7BscdKIzGb/++gQHELk2LEWyKHdlSDIhFSAMC+tIf/oLp7RVL2cNohz
PfY7IIYqz1PpKT2HrYUwMre7xBV8c/7y5BTQEGTJu/dv8poMeIBlGMriCYXrcHNHa1fXlM1u5dn/
Usi0K6uxKRIsD+OGQamXUovebbBsYpEEzXWNGU/XqWgNec2wD1PvwoJS+00Tx/2kwsuFegLRzuB8
oXN58P+N92/J/ByeYYb4ShUwA+yMS1gICaUija8GIXckronn0+xRI0HGXgD9sLUxzLLHtPQFjbdX
RXgdZfUkrRWBr7e8LRTGLCSm5WxzFy05TiImVsJqWVKrrAUiSLan1f69XAYcsQ8UDCvV/apU5xce
x4snQhglECVODKic44Vx9/NVN+4BYc74gkpY3C3BNxQw1h9Ak/Dat4OQqC0djUL3i0HU2Uiu/Wzw
ZZYrZuQHxQ7h+U8RX+TYf7NEAPF2Sb/XTgu4/WbCO/elNqbnKudI44Z+3OVFd/tGnhXO14jUGKeB
6didFCK5BBceYtRi2pOhc/julEXD8GVsQ1SkSy2rFlZDrkPqGDtI223U/bQZOuQ1XhgUB+MVXPT3
y+9ott3OKj2EkDLegCILXU087QyJ3ruyFG+nR3pyNEdbwV+g170OI3yAWYIZ3H4JQVQB67RgHtEl
dxFjCCBeHeeneg1/BphoOTcQVewT40Uu4Xw+k0f9CE6tURCQomncSpj8uiSv8s6PM5/LJp9aSBgR
8pMA1Hq7ucHDbwTqFSsMdidkxcxmJaXiViKDbMlTqojmgQ3Uw3l0OnY/P+G6mUq6q3MeTkYHx8gW
CNO1BCotaTOosWho4AJcThQ53FcUOmPrssuszdgV01eH/4wZ8cXubnjfQ0NYek3M62JzX1Svqjsr
ZX3LqotXi7e97zo2FpbumRTPD6cHkUr01FTH8YW727HPa8087LLAISarZx/ZenWft65sCaI8qNj1
rkCVWHK1F4rrtzsHxAaGwZOszcmbH8aOAdcQZ8cbS5BuLBPqsDzHSRyXORuoH1r5IW6mnYE8pjPy
LlTuYNEj8b+PXqJaum25+EXzCaexr6sZE9uwEgWO3jpyoqg9qtzpAI/eklmGU2sGL+6+PpbDY69+
+J0zUUEqDUismVq4njjbC1pY+B2oXpJ/c6dP/a8izZ6tRGXwi0L/IyPLyitaQ/XBdA4fHTpSEW+K
jLUKCJ+8jPR4YosEYsGYwwmKfjkYaxvXr1wJCCnt5+OyVUsEviXWrUw1SNK/E7Hy7MsM//M2XlAF
7QcOr/skekXo8B/Us64K/n5zo8N9IO75whNxQY858WS4VY7d0E+oZQnOibw7vBwmGQWHV7qT56Bt
ZFQKXvalC+d3vcarN/u8H6PFGUHyfHpQOy9CvIi07+oKps05473s7NYliYzenf+lrLvo4Svfg3p6
HUzgfFCUjebIGe5kdmF84xhSu3LfXgDQf2ZqzQeamLfDDabk0yEzWajuBDydcOset6mY9soebNpb
uMydpzBkkBj8i5uZQvOUtxT7jK7OGTjMut35zVgbeuyGWtADGsfPdxaLuZ2FQwmbuMoBwe6cvEZF
J2DX2ZT3hWnOI5vSVW/5DGB7FkfwNEnY6K6KZamMIKQBbc+PLykJjv4vdAtVg3ohikscHXLyLYUD
895axUK0t1hDRy7fTAGKbbxCIC9MReiTPM5JyvMjtSUg5V+8BX0pfA9wJSt02hF7uI+BC+oXFuBE
2KA2SNnO2s9W4LIqV7rzxGO5/P24lVHQ4vve5lU2bzwyF9tLK3tIf6VY2OwA7ptBHbJyzDjeRWhB
1a3LldwLLwm4DRQJ8m0nUIE5ClG4c/clJogE3C+gesz1+/+mwsWNNJEnNh6uATk1vHtAJoqGZ9ZN
DihGkdGVPrPmDo1KiqmMRSlyujZFpV9NsECTiBtVi2yNkZ46Pp/aTj9TTxJwkQs9Hymkuk2xAm4T
BoNvnwgS0ue8x9hY8oNavKTeY2/1uBkn3hRgTn7uUoRZi8YMtig9FBnbeqxH7s3BCpBrIv2TNFsJ
DNZdXraIYkUrc/dNfTwfDo9ykttF0VC8h7neaTUlxxI8s/jWxmbXSo0Z1CW6G4WguVmIwYDqDGlK
Zv1NgoRfaMdGjWv5ZTiXJNGWo/4MJZtSnM9+wKp5/+KySOpf/ioCaVAVjvAGwd3QlNrSRfVCG+AR
g9qGxJ1yhE1N1aNXfN7KomXdi9ZThwinYCduvme1T/ucJYbFXEKGV/oDIc4ZE6/5pN5O8d0Z+OUO
jMX6lPT1Oi/h6b/X6UzxP/8SkVSv/y9LXkBc9rKKNuoc4Hc7zaRZqhBfWVKEdX6sc2Imdc35Nwde
Q8oaxuXvCVy5AHLPo8nkQQyTaAOlJRY+GrjWotybPiRMmnz5rIQlcCYZB4/lga2mZbG9S+B+6/CL
+5k8oIlaQC4rpm6gzzoHQK9FDMsrohyYDAuuJ9eVTe7fFBpdicEFald6jGyd6+1zSSpVjeqMtL+3
aHeMJy98oXrqhBrzVzqeNvS9COLdn5m8C6XklHrYRc9McbAVoR4yS7XOe7B3jlTc17zMavGWj8aU
eIecOv1lbionmfZkepsdPd3nL/DyYZ5WuWPe5yW28Vsd+YFcUwqU0+EQE5XJ00PeA2iLFkE/sbLA
tufpzS4JcAqj/gOZ3b4jLSx5MgPp4VDaLgqO2ZN325BNdMb701Os77i3K8eeZ1vC/Ck7CAsgsMAi
inSIZhFtRSYWZS/bGOMUpvgT7UzwumDfiPierOGbpKTv3TFayjx65BwAkZp+2d4MD7nlvQM++kvu
hQsxGQa70rZVTrKVv/XmBEQAAX7//IhCk/GmZq8OvOvtN21X1xNQ9jptpw==
`protect end_protected
