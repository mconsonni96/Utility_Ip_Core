`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
X4z82Sc41qTzyn7uzAI+4t++YWPhHPZKEqWmzzy53FZeNL2qeX0+KtreAZKWjUxTZzu45u/Z+ZNm
X8LNyfqGyAn3kx0AZlsPYnAdE7MYK7zQG3Bn5S0Ew3vbMorZvVwzk8j2T7ySay4hSEQZR7kqa748
haL/QYLCX4gRv7qaZv/BqoQvD+TqOWz7l9ecD5g62WhjwdL8FRZsEhMPSofwWNGcK9NFoLB1GfMN
cDghYSmV/YIXh7FIQCeqztGOeJWgiVETD75NTmTGZTDkdHpbobV4kkoybCnKFAN6cfJpXcnEzG+9
eu6XVl9rj99PR2JPZpMvE+C/RDBarLFpwpmk+w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="TY5j4Mc7qDE/bs+R8Vfhz7Uc3rlJ7xkBmiNjqh5U5AM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 83056)
`protect data_block
4PI0gSjy8FdPu6zWO+7P7OWdG+fdzYxp9O2QOWxSLnRSSFdy91LgPiFtQj7aUArGHokzwRcObOrl
8YyKm46OPEJ/SwuYh8QMoQHMOp1/cJYrDykDqEK/SnE7oCa+VdbKUvh+TubRxS/BdMOtV0rUTyeK
WIHgmMh0/KVl06E8M3Ica2t/lwilOT8gbevK2oqcGZR/FSgC5vCcYJweg2tuJD/9bKc51TTRPLQ9
48dG8DtY4XJSFDgBM4dj0jQSzEk5vdhsAyKDLkk6Y6qzO6GT5tvo/1JAcJInE/L2GoEeEo5ugHjy
tBekDDYDUWzwzA3ts8X0+NgFIqCVj6g5EUn6WKDme3rO7+TVTCCavKQtuqkyU4Z5vL2rWKAurB2t
KwCvHljlszQ/JaHF6ynMSnPm/D+5hR2yHnsrUctfCv+rwUUxlIbnCY3Eo05Ftn6b3lCxIUekfTmG
nFrjjs64+xwXrNUopMkVIZ1dYyZbEFGVXlml0ocgrdigXLbt3yJ2bmwuIpE0hXZRiVPkMTjIqPFe
ghYQ4AGpN2181eJyHpWmiSDL0qZ+yOTMTy9Sh+auF8ypeGkQ3otpG0dv7K8VmXUIPmAvadSFgBg6
CC3/xYhAK4qZWpjE+IsdLt7QcVIaiRI1pVi8RnKqxB2ghEDEQ9EoRrciaKPw3ZFi0qM7mwjI0Pnt
8jWq0PAGoIvJHiUJjelxBtSsdEgZ9ShWrSnU44ZTqfFyFEnNn8rjBngxf06bwXGEvsmY2j2yQtxx
TY3Tjt4ugI+qNIcrwFIsamoQl3A+8WoNobK307Zz2eQtjIFhJyiGXNUdi1UJ8kwbcenBWaVZNRe6
0ojcWxLdBkesTZk66YT2wWReeb8pTo8471xSvrVjMq/yJo8ktpeQgewSHEp4mVkXztbOg1rP6v22
Ou9nL8txnJkdmY1+Y3UbpOvK4H3jkGFFCSVa4AXVxScPbHBDemT7deaRHofUuPQyGJLLZsF75/re
zxUi89gVQ/fmYDwxK5Oy/+SqmSi/xo9DjnIJjg0oIhkF7A4UpBfBB1tbbzVxKH5bB+PGaaaAZciK
HehcK17gQijKTvof/mYP+4aaGszIkMahxR0EUPn70Ql/IQMgEsrUb8sS/QoJPR99FhvVZCzXPUeb
Vyi7ifs3Lz56HFBYCeLfrwatgMyR60wPEFCqIzTvY+fJl7HeWm/VYhMXz1rz+dYIEFo9YuukrUst
g+tUT0u/bkYSQg1EjTwEgC4PkCbwa9zuyd8cF0JapIE3FfqWT8LixqykKTAVqNn/3d4kCXomfzCK
aFwH7/4OHfKhq/VPTZb+1W2G9F6zsOeL+cMBLfw1zRCT/Rzpry1jklrjiuz368BTE8JFZ8iFYGYG
3K/qz1mzmwpyn6FGayMBM1QlUT4mlrq1iXwpo60DX3uWOiw4Yu0OB4+hOgoKJHNWcRoVaZFs+m1f
VeKw8DvsTdtZrj2xjKmjuMBrnmzym5cviRzzDJcPcMM5SZng7+AGUtLPYP4q+Nj1VhyrqNXN+WFq
LX0XQAIiOeEFpkRsswrKWBhsI8qSCw7Ox0fFsVIL7rvZqC4wH7fddEhoBmLVJxYprf87ncveJIjB
cqet2TX66J8cazfBPAZkDW2yBaT0/NmMbduJsXZnVVey+1fc+zVGZf3uvWhkgjZ3ucAL9BirGBAp
Tfetu4JIY18K2bicz5E9K0YqMSvCCe7JFF5KUAe2xk8RoK879cxqH29uwfwAWU8DiinDrHVxKo8a
mIBsT3k+h81ej7MbDvUGmgh3EpJO0x2CUXUwNRSNPfslC4BCMfyYVMvbGR15xRMf+gdlX3WQ7230
TRt7SOr+IlqPxLVnmISwxZo5jNb21cHKtKs1ZmajKhcABGRVWE4/1qFXDIvkKHGoNIcgY2d8/zNY
LNCy6PLidRM3TUNRTCG4zy+/BG3BynHBzGwpnPx3FgPPYxyTVKu9T+/svz52Zbiax9ov4CqFRdvP
we82Nd9Wbr5MAHtUDEkHwRRn2HCiz2q8wSIOzK9bN9FXw9WWt+iaMqTgpOpalxwMG6/sLnIWdLKH
Xzl3ih/nwNARirr3esUA0NLZamrKb6vk9UmqykFZfLAGMiRz+A1U7WnW7rAkxNTy/n5UdpDbqFxn
ZSYKkjt4RGiYCmRupd3zOhZgKSsufo1A42ExsMW513qXwVM1wZT0Rleslf2kyg1ZVih1gDvRNDOn
o+i6iAMMOWGpO2qCdglzUrGuMHxMLMYAsbp2UzfOE8MW3QL6/dzq6kER19UwPGfHSJp/KLnjr5y1
5CK1grq8bH9C8vp2AbUIuucK07jEQ8Jks1OPZ4C9jXO9qREvWEHaspTHMv+4WrM6ju+uDaad81ev
wp/kjidUO4LWybXrt0ngPCr+Ik12OL+ktcVvikuAeklMQvakevtfFPN783VuJwy5UHbKhk21d+h1
Gk5/cd+k4BAVKc51L3xbRHNwqWIBdPTpgpzSMRhiAM5uywgcG3OAyOALwSOKSknYYfQ7dsahcRUp
cRKskJb9xyp2fGL7/1oRtGET7i9S8JWx0OBSy9728hRZ/t/FXXmHToGd7C5dSIYocZ4JfygUe7lL
nwp6i/0VlbUjfURHVH520dH4pigN8a4SzlGXuwHDlEn935DBsH/zJ2VC9uVe6KLcFFSFrv18ky+Z
EArlhulGcRZlFjepnbxbUkD0CHYL4RxQFIZ8XegwGrhAu9cPdvxnmQUyQKYg4Iwp2S/huudEsZxY
auti3/wBnsuRF1Yq1eV4wcRkE+BXKWgxIXwwjgK8Eh95gbQXVdLSatt4vsARfLPD+IK8nDk/JNAO
vnNA+mxNBv4q+afZVmFPaXV6ib8L8ezM+qCJHyvHEZ+nlrWriMMto3FDiVFlHuJBggKR9knL6hhN
OaSbn1zyS2BKjxjeehF95VFL3fKZ4CDcLZx8u4aF4UQbolObalZXDS9z0Q24RJuUeZql53mXvUC5
z4x8v/Y1Nu6oYTvMNC6T4HB5DlOU2hkqUu/epKSwjJMJntIBQtz1OxGRg49pOleZzKjB/bvIUaAn
jXYsDqE89jfYxWdLRYb2Sm/02k6wbA4ihxdbuSpjJ2dKJOVJikdnKKRbnNuxLD/6sR+vHvKelvZd
l5t1IzJzNUpMhEXQV+Ja8Gp3c3qOYP7rMMy0nLMvXnbwS878GBxwAU4CpHvHnG9ejC81J1ol94Rf
HPKCIGZzXf62k8/KeRIeMwMC+XfqOkwfSVueRLXDyV/yCmMPqYSzA7cENM0aGrDY5AH2TYR6/ZAu
k4vEZIBH+nKxLVBizJ7PcZ1X84GlWbZhkS+ID7sFLZkUaQUosVS0Om+Qrfpob4FxsAeqzbdytpUd
ho8z1cUpBRw54vjgpu2gmC4YLYetp7sPqYZl+3PgfXNUJp8ZVm19kZ+3rs6z0PjYKVZQxpdQcFY4
RGmthDgcEOzCTMOg9GdYubWzM4yHEH4peJMbG5myP4RuI8phbqO+BsfED06zuH/Mid+omlZIUc2h
9nTm9mI0suyx4u9FbRvloO4xUDWBehnLaOoD/FxJsk/ykmKLNAk8suZMLL51ohCDm4ZojYfpNGm/
cFEUYCNxoRniZA+L5NEPknFyOrkB8mvAyizZT6aTfN40q9HV+iq9jzeWipvuxbfoYouC48Rrooru
rZDUUn8buTH7XQYcmQWdodHa9Q/nWOUDm+kIZqMN5PQG+Opl6BaBbZjLwrEOuPmEFvOaQd1xsNxN
e/Bldb+jFTlaa+MP6ZOdXRMY0Es/meiwD3BfrObM3XkDULjAOxr9BqUAp0e3fGjcVUc0Nm+C/xrz
zhbjsYrrHK792YAPnxAq+pMiKNL/cV2C/Po1qxAgm2cC1wfMFcJzQEd63sV/FObNF11O7tJaA31W
w+tR1kH2qih0A0mf6ixzPuzi9h4Ech+ugaw/kov8PTm8MaL0X1SrMfqFXNXUDheSL4h1wA70v+8P
qKEWDKuM5Gn2Ib6LlO9zVf5DtaDH1thl451DEHy1+lfmk2ANb4Bv8/3CpxROYyai1ENb7tnOysyX
Fb0vBQpmG5go820nuu7BXXtILL151zPHvsWMXtXLuC3x1xNCjy0cQN5Epptb22xsW9aFn10EIVyp
rXico1T2PjVDwUtGXWddP3nkfFOO3eqrNQ+GAvjkFyx7GTh9xzn5FZNxnLtKjaPxdwNX2/tX+aR3
MZs2eMfd3QceQ4uaaIdDe3mIYg3Gx2MPRCVDo7MXb0a70tlY0NSvDzQG23366swnPupYGo/8SZZ9
3uYcMZoHEH0UU9DYj0y+Saa0Lvx1UynW1b91wougFtMisuvdsY7XnoUKOdJc1lvfl9iiO1sC9gs3
BvVqp30gXGwDcXQEBPdJtfrurc97MAUuyJT2JS7Aaluop0jNTUZOM9NNijXrd5bAdpceFLJzIRj/
tLP1SJLmM9icQiQ0nnBhQXMFliOT73T89vj1S2Clrz3lSP/jO4QHxCnefQH9AN0Or1sGweG2ieBG
K9k+By/WxdjThwU4gGF05wnEaSBfXkXlfFI8P5fXoxyQYXyyIo/iYF5LwhUjnvGhm/UtwbSQocVA
w0buSpS1ADgUgCXzt7DlQCns2ChnnQpu3lsNDRsJ6OVBoWdYbStHXp0YXRickSqQ8LWst4qjN1Hg
jMDTtJ8x5zaCs8iXwR6d5V+X2rjlVXId7JNBAohK0JEpbieKzqlT2bJaUgwQU2NLkCHbvgb4msYa
ckknShufCF7OCQL3ijQCBYmUD534r1JQus8BYmuanPfkHxeCUpqUxLPSzQW3zHHFB5EhlmFcYkYf
nD70OQLF3672pVLlfKa9C2PaiSVJzNQ88/51nRH3OE3eJqRC6YnAQ0LYNpTkzHWqT5bLlq64mPAz
BnOpuhn0015KLn1WjEYb4rkeKp8qOeZtjz5Tn0+7GjUJwpjPLFT+JfxOSMt/ep6BBhDEftpZTzjk
giD+IoQLcn2Ul8E9XsMnhzgQp3tmv6nTEbDGwcIxkxicd1lrWzgeTQpRgS4VepVB/jThO/Lsh4L1
V0h+5afg8pxv/eZaiVmqsLlXa+C+dt/ULlnX3G+Mj9LrcdvgK8zNwZA14zDylVCjYmqtZnOwJEym
BMwrSx1sYy+Tlg0um9FP+926m+1SglqYh0rGYoTMdnQyHXlNneRXzuNEO0UogjZV+TPZHbVXt51L
80ryybVe/v35NLXdhKYaGSMuc6Z6fRfM9oKq2RQ0S04d+bfa8UaxDD4K8RhfiTstUD7oXluAq7MG
LWmETIsad02mhlTB0DQTdjHGdag4UjQEA8kDFvnsKqFucycKE35rnToJjdqxt20xB7Lky2Qcc19R
TZ3WX9d5jTt0ntJJDSZfXBHIYubf2qQMA8Kp9/XqezShx5kHdMcYQdSV9PxrIjzU6KcnhdrR4mjr
LfyADEra9ShOIADSVYagvm9d0qpsH4rxnGT1QhUDM1/NPenWGbjG/93KS9EVgAGiy8U5boc3LHXO
jrZyDYJqH4YpZQerO1KAGv9RvtoLFoqlwc9TeDnvxiOlj777vQrpBhUBvFcZXsTv1J5hU+OHdDnl
x8MkG3omz0ks5gl7OrI3NiEliAna14DJc/7wlzeQIwxYA16L2rX240ONlEOOV8l5oVLU1Uf07e5Q
d3GixwuioYPwcuk4E6m/dyHG1bCGmjrcZJX7rZkTCYypSK3ZN4jlEsg1MPFKjoipbAwSgxOopAHN
t1GcQ6VeSALGypWjh2UhcwGWgUDBuG2uj05WcksVEE/CXd+NHGRUilxgFRsSWbCeNioABOvbWc9g
ZgEgtqppphyW0xuw00BHPLXdQm//fTc3ogLq20EOEcni83KOrevJQ5s/9gaSbsEU3fDYdCUL92+Q
CJxtXaQZXTcYhgGMVBUmXs3RVt+4mC1ospmyyAkSwu/amvUz/XFfu20Bo9E9XiBGEjhDhysGbGsT
QLupY2SCHIcLKjx0mgv8d2MvYbypP/GDbPgqLsV5heRcKNKJhIxWQTClJMxytnxM73+x7kpcMV0O
23/JVwEII8czbBU68oxMrAeYTEFYGkLxQvqtC8HTZDmHgWmVDmiyU408BKdGcjSZwGzTXwv3pKqD
rkBAz345URjq2UsMo549j889sUNDdBzwlx0pngbyiMT+G9kaaEWjBVExx0MaRDiVmKpAPuwvvI41
IrW79yK8ozbFUazDUj6zX78CBc9jcne1p4hSeK7mr2Zn2vBoiAIRviszEpUURLKUB1EPI+jzB/Z/
3g4lXm0kOfVHiCDYZeqXtwZzVnqg8i4eAGl1Y2tXZ1p9MTLNK7b8y6hImylsXM6maNOkPIerHPD8
LJDezT0aZ4HPjOE08Pew4EHpWFZwYzCgF6v50JiuSsgsDJ+I7ky7uGd7+LY2ElUYfrAl08C6bO8r
ZDeAyAHKnbhQZDAyTsZ12E2lgYMwh2e4mbQkVNLRS4hAzDow3xgbJyvA+XJdR+A8yEqs2TGnkqRE
nlC2D5sR6ZqJW8KvUgOYCJZ6/LNDw/9T8Hy77fJ5A7AooOrT3G9PpCb3Pu91FkiPBBME701EXwtb
vTDUHwZWa3xQ9EpqtRbbOVALj0E2BvToHEZ7K9KCofPAnidrZp1NsFURfLLVqP0CeGoHKMZyh8m5
T8O/NG91bMdCKWQCgtnbVv2d9vZNcJT8+K+5VlpocgxGiBd9xS3fwBuCN+E6m0A1cVPACfDBG5FE
QNybG5qmbUF1LPrhdgpN9frd17bdk9aVSBpa3waQpxMYHjvyUO7AVuSOQQJpMMot2aOuaFyOHicx
bV7OHvSvDZXX+fTf9qjtfgiBYSaDc5fkeI664IAdW51LwZURq40Wr0NxtCv5iJct8B5rZ1fW+HI6
gyKFCkFPJEodWGU7yCqY4l3Veo1E7Hz9+MPSAhOm8uVpmv4BD28uotQsnodQiUYTpN7H7yQWQAap
4NyoWaRt6/4UlJUEMIBlaaTmeEyZysI6YFFCMnSrp+Jo4ZSLxRxlQRr2l9bd17I361ihKyUhw4Iw
k1Dw851hTaM7o6z+42ycoXJ5FttvArnc3iRjYqLfzlE10hszYkrrNCiu2wtVN0yFwB2Wm5Qm6fao
TelTymsAubZJAjlIqxZZkSdJX5iqKyeXT8jDH7p/a2cKzxfgFTKb27eu44dQJXB8ZVUStc2lkRPf
FfzYQjXo3WdQeI5k9pUVivzWhGulQVHd3ZhGU2C1VhnLu+VF6+bbqoMoP/Cz1iyUWZoI0LXUvEyr
iBgk67cuOQ2P67xhbwN6lcsaFzkAnL9+LtB4H1QNaDCNaAoQkUPMX0+EYhBFVIb6DgzbL3Avn8l/
mDVAbLnHRt8BOa8ONkbkoqtrftq+sxyYlEFt65PiVqbIdka8ujZWLVcSYECyEHNjHmaXx+c8ajhO
72q/YrUtf1FyS9Ixf11vDLkBrSjGEZcdSeNbis5W8TPCThOxLGolF3E2nkm6PQ3WEM5bOqbdTjko
Bqq+yIS/cugvFi8ezIurwOso+ZGGJG4X30478EAXHRNbneANCwl/TRp4wg+Trtz9myR/7biGE70x
Cv3nRvAY8bz7UXfuoK4aay7YTLQ68152bqux0hyhew9nNenZfk+wf1hbdMVWHgRqTWltIAvwIhJ9
2aSx5rWh92nW5w7gg2r5/ZZ8oZqa0pHLrMXjohevHvRavdz8NrUQoSqxOrgZ6HSFoj/2qzqaAlUU
kb15ht0H9r1W+DkywxfuLT/Gs9p3fOR9z8rp6tE269OIPeNGfsWs+TwUKi768qzcQ10u2YeLBT6m
GSOCpvTNHw/C1QfS8qDZzlL6FvpTkWcLdfZbYDf4e43M8vR0VLTY19cSPQbfUrU54bxz0geUn5/2
INHmlYi6QRogxcj5P3J1nvztcifvG/fXZsaH5B9qqtFp1yJs7+bjENPjCCgBlPjZQwH5p/dAcphS
q8Fore7y6HfAweKVVH40rNdg6Culv+KU75dfVlxqcMXqg+/O+z2UmxcarAUHJ/5uf2LapSdEGaxt
MY8ZTgvwbnRfICYJwq031HBR9aL0sNNX6s4f/XM8ztZMBSidnEzRriC7xEc4y28FZSCaRE/Y3VSW
9fs8bUcaLY1Bth/L8tI1t7ncIgPRbafUTXUydYhlwqjcV/0xGGWbWKRpyUtHqgoxzca6ihYwrwMT
v4E49P/AyKxTq8/Ne8q05DMkR4p6mpdeyPGEOMvy0J9T/9lpX3JVabemzHTLwOybPpIKKQ0yK3sH
vEgQfYoWgiK4XsmwG2nx0yiJPZTc3+RNcQpkB1KCQMwozrQFlq0Y/WkfippZizd7A96SViKhGLwe
L+z018AWQxmtCi32nQB+f5sG2nZoH68so06wgOFGxQidl92fKqLodgoSqcL9Wc2krVNWetzCQqxp
WhkCh6SAJyX+57YUjOXJZpRmE39TgMPOBbPGzROI1+/ZqHyd6cRVRGc5i9+orb/m3x7XhYT3WLiK
iAao0VQUxij29NkfTqOI0S2aSj/J1amZSgpPRk6wfGxiRmqn4I/65KesotdKSsL/C+OaZQ/GDxw5
odZuo4Gzt3DWCisENYi7TLS4gUbTDRCm3z6dtMPjkE8RtLqMwych5NKaaBx3nPoDk0C+K4vHczr+
PBXT1mlQ4XKO1U1p8pZO5Lz5Mnr11FPgaJ+iKUZHxzNngWZ7DqTBU9esZWaj/+96mPbknbIxd05p
ABGwx+R120VnM+6z6TE6SIvr/Ngn/22A2bMIRqB2DOBJcX6I0Rg1cesP0UdBIAd8k5RjoZNKZ9Uv
Et5CpI65wHylQ6Zf4O47gNBJyJypChn1+pa0Wgcwrn9wvzFGLf70HhIwH9BOlVCKoQrIyQzVfOKq
dHcWiLXx9Px7vDLjkgtOTITaPc+NmhwjnS8KfjCDNyVM+2Yg5QJiDIXkDiNKNLWm/vOwjvOoOAW5
FE/+JF6OZqm4u/99bZ5+lwDAoTB+RxN08ZR/3QgBKspcsRvukAgAw0Mz/cZYuPXpQ9iV+ozWVBm8
2R0X0dES8BW6MRqSKPkgh98fJ5pHmn0wGo27swmoMLn1UoySZGfbblCsfzNqYFSQtUOno2WlzZYT
mpfcQ59J1+gU0lIAVI7VbPBPex7inNhWlfZim4RAOeu/b/qTJtCSiMWn7QNVQHNim8BHffhWqRqZ
jILP53NkAkDpCbOK9x7/dIt5YNsjrLt5TfmdiHMxk86DhDNzLzf6A5dw62InrLVucHneAsOOvkI+
YErxT9f//duPS4KjPFSxG7COr1rqMOyk2zYQ+Wmwkd1F2ds37ZCOn2YOZvZJGuFEoiBn5KksEcO2
NBkI2GH3v42whK6gAM4gpbhw2WYNg2YA5OofKMsJKDKBNQt2iQEMDK6jC0uP7pKIQryLRP5P4TFw
BLl8CSx5aKvupshN0CpHWWIDuEL0/uiINAG3iCv41K9zyU9JPlYzU2GpT3Hd0rGkt8+1ReQM3iX3
uTXMmr5GCgawkHEX05HNEkhWE4ss1gqEkJdTSIju9sYU5gu3g/FUzh4jXlkUWJhmBIcA7fk51RCc
ip/oq7plE6ycmxmcu9rQrGF8UZ33rRm2G1MW/sZnuwyH85Ey5aIHF9kZPNUTQYciq6zvO4VjNaQx
tNErN3GogyRtopFlpNwM2ydtSDm49WJ0zpCvHDpQlrtQ2eW5swUOwbem8VwfZr/TxMBo3Ke2lBci
L1Edm95q3KWbWp1sY3Lyq5Jvy82FSk5vnBPuDdApMgiO1swtMV3tmCK+dp/N3OYDaBrglAclIEr8
oy8sdZehgWtPybqrO/HnpqKsQaYXTmDLO6somhuiHZajwXJKimrXYmOMBpysLU6mNthvwjaPPpFS
dW8GHVuFv1XVL4aoaZ6Myq4O7T/eSyD3FGs2zVvhmMTjxmgS+EUIOe3LMaJ7DQkAU/6oYh/Rfmoo
8374UhZOWRM8N/Nbfdhv4m8qQyWUK6G8U+bYVYFgk6UvL1XSkrYsYc2n2XRcFVVR9ga/Uy3EOzB8
bxbQhvrbHgoMWAsjfWpwHjQCNaNFMIOW/jv+UdMAN+ld533Fo70ejHoeFGpourcQVd8ylWVpdwgI
AbgPzToUfGg+6FTeemHB60RocxRK2NTb74YFNK8hnhRe2zO6nwlUcgHh9+t6sIK42ki/F71kJxIB
H54N88MVSbhmNsv1FlI+pZmLdmEajBALSF6gbPqrUQdixuPltxZVi+WDTKNXOciJRiGl8ZqjSpYJ
BI4n2Nm94i6bf6AGdwIc+KiTWfT8jfsACT1pqdAKY3LB9P2Ha+EQgIOClgDT5JbFN9P/aXFd0t1A
GsyJ/u1NWP6ZhocU0mMYxOPHcjZgA+hH+3KPmBbpE6S9GPmOys8DlqkhwyPwgYreI+BmaG1EsKf0
PJZVd1G1B/2wlBUQlpiIT7LWZPxpSp8RlXU4u8HzlJENtreMZNXegNsB0eloBgL8u20RJUAGJpbS
gcq+UhY9VPKevg1VMOxjQRgG69j0lGfi6E68giH1IWzLHmownroifqSShL37T43LyBCv6jV2C+i8
1PNgC3gEYgT0w61hUzJg/kTeP7MxYgkGR23TRQvHQxy5BFdjmA17wKHY7Kh471ZfOsEsgZgNXO4U
YeexfKzFQyukNrNxRQe+8Avh+1oln8a/dPyEOMNMs9Kk8qQ2/C4Tmce3Dbod0GNJkoE6wXmEjEBB
VU2SesN+2BWKg0u+UlDKM8av1mPTtB5Dux/aD0znKixqhw35a3Dg9RqyvkqVI33zLxmOoOI11FyZ
s00K8hnJx0uaXW7usuaENoyXDwDMORQSt3m8/KsaF5OyxKklQYD9XhH2PsA2W2g34zLAoqiZKDuZ
dKwZanfTNwr/TeROiQIHmjh32CvTcPPDW0Lzb3DRk6rYFRdwAArnEzshzhxPAhs0VRm5xHhgkcAU
6tszvKotD/QYNU0S9YSz8pxtlkg6Rpptjh1lImnwcBKO+1jBfggbHJ9ZQELBBPFRUtdBEJfUX/QY
RAxSIFF5a6XFMj7pLgOGRPIRJb1FJqewwQXGoY7Eu7z8VNt1zf+Mnirhif0AZDpqTKPvjf4h0VUL
GXWUv2ExUL1ac7Dxw1/BkBpgJxAxfz+qz6y7gsBOB7eVQPUBhj+35AUFK2znkQdATBFgYVYZiwqW
9wpeI+bk+gpW1axafXfUNOI2jKP19IWsKlJ6c1X1CFWTv616TNSFKTCa/C5fmsNIIA7OY6kyenn1
0ua7yxksE0d+fa46eziRPsy0GaqGl5R+2/ucJ7yPrD8mJo3BEtL5YWvpDyaRssobwaiJAUrwKl0m
0bfb822sGOMsQ3LJf8P4whbPJNOAcDs4WRp8KmVetkDA/sI9S4f4KEewUt296vrMJo/PaNtnH4WV
RKJ6J4g8l6GQGzn0q72Ja8WZUjNaAYgIsjdK5KvWgnLxadgSnb0lYTv3E8OiNETg3z+VeTaCNPLY
S4P5Wtdmv238FueAelWrOqmZqOZlr3VgFhr0t6Cue9w57P1jr0uRgE4fS+gD8mh8JO1eFXIFOQAu
3vYsCgpQgoiP5SKRvpAjFY1tA9bgmywgjImH6mek28CvbikOdedBEik6NEi+MsCuImEPSJdCQCdh
2/LanUZdBm3pZcxL+kTb2czEW/qUcC0iqLXbzWjtnEcp0kOnA8pSwpft7uWjp+lB4fkiYAH3J9IR
q7CxdNQLcJix/C0nerxKRCqTWVMNGXeLTzXSLVIVLDmbIlWoYuYRTEpF9T5qQ359M00M39+emHhb
W+o3a0z2CHxHhTML5vjmnHQkGAioMvmdiJMLzRHQ4pe4ebsbuDGiNvIYx/1hgskbK6XZVEfIqU4n
K7zhWa/bICKiD4FSiZRXJxcs0NvuX2cqGcWDkJ64sU7AuWXN1WKNQaOStsZ9D0Erf3h677j3b8xe
IMV+6CUuDGfbCSFn+Eb7iL9NfdXgBUpjQRgu7qYDk+0an4yApCz+Ac1RY+Exka3GVoWRT5JoSeK8
3CnI75Xx0xpkkAde5O98fgLY/QVvKG96eDfJQCqL6irRI3mt51k4FgzEY5hPq9Av3rLdXzTvC4S/
mfWJpZHQXRmMx12yRS38vd+iO0y2Dbr0ZTsoREyl5CgRQkWrqhlox+qz4rf6U696flbeaVraZmiL
nnHwHg69OE9Y+bP2bsYvj0uaq4AEim5UNbw3nnlFIACTH1eK9kKeuPey21cUztB2mMOk4L4KTiaf
GT2rM9RBWkptpvPcnfZUk4yxMpDB3vGTZ9RC4SyDKhuX5KSmp9SdYq1oP4ZV8FAwZOxrOWnCYXW5
9AMrykaHkWJLcZsz/EVhjbcNBorJevMv3GBAcTxRSGwlw8L//l7eQQoSi0c+Bs1p4bX4DcHvfg77
eQpE1fkNGt8KCFWoADx8s5waVQ7mGarIg8w4w/xvOnLnbeY3urBhNbNuUO4oaZN8Zd5mJWiOGw6a
MuDQ6eE0obvyXS+OMSU0HBs4dj1hS/pxsTQWeDLTlsWYMeZoDL16GdPe7esCPqcyfFJdHLI0zr+J
1FYXpCCajTX+5kBZIybCxfa8286VtIXWePHGfqbbGBRE3xfiNgrra4zdy2Q/FTIK3lAGUqFZV7p6
wOo9ZHSdwCR518RHgz+nuo9NF0Z+HrOxgF84H9I7LLbl4hvm+jlvNm7d4m7VACQpWOpnLfowFzMt
B9AQHN6CK9+OlsHO9Hjv9NM9/xACPsCt5n/Mg2FBDUMo6pGIFpt1vpecr7osGGmtAah69Vgggz13
xyFCZpMN0Y0gf7lZVfMzzwCCLeWm3dXu8T6SW/Iv1rNuo1NI0eyThp8262ZR0NVclsqZNeQeiO+b
3wW8B0v/IIcPtbAA066F70ctoEeEpZKX5K92oOpzFkdukiOMzBrdfmY0o7Mgn9O27eJhUqT9B0yv
2hSm7MjQ9ZzPFzwnPuMMZEEBQL8n4grQ4EYAqNKG1srtH5ji9Ew8WlExW04EVB+g8NMb4q740A6o
KjwTKb1VsrxG0iqyYBDxE9NnAvn+ePLzhS51ifqkANofEbE8qZG8OZb8o6ycQiIYq5oipQdRpSYy
BbAFowFnzyfW2ztgdMZJcrYNmiZgjyXeCXivpOkZnbW3NCDIpD2biUYJn8w8QcCczUGvWFQXmCPS
fPQ6qpQQS5Z99EHyfbI/YHxnVdlj1CXmS1anZ3c7ePuTA7VJLbPIfRIkHHFFiUqkCitmUUaVjDxL
XaQMV5s+9aXiqeERLnsbTnOoITkWbcuTmz9DYnAKJ2oKHp6JFcWonXq9sio0MD5nbzJjiHWnIJZA
W91yp6gXKgxdDuO5YXtqYcGhbWhpfRn7KT5oHc5QpLdB/KoOXzuki8IKM0idXHkpsSTOZLV3NDnV
zDburst/n0vXJet8cUAXTste1rawg9YDLOPiDbt6kE01NQ8mPvx+8Ik96YVLmS9djBbTH5Uaaxql
CRksk4PKorS4sxV0nHkzJinOoFYFCLqmHqkNfW7xdtixBeY1Xdm+l7g0Mf1QjZ6FgTFwu1Q7s24l
tLP4tTc2nMJ8/UamdXVxGkHkcW9sLQWhf32oN0yuzsGgWbCsikz2vO0X0QfKIdP9Y155HcYqEZ0S
AGO6nnjOtr/uYZBKPEBfTJ0xrQJLRpATjasBh5cW8jY6Q4jBUFlkIqCv0JUCIccmV2hC1S9m3l2z
lVc4xQaqu4ao0QGNW4t9GCwPXaZTGiDXVHMYP5frXGlJic9NE9+mPs892rgq6XqpLYcUkr3NGj9B
0omCu20qjFwWYyLa///fOH7KvOB9BUglcRdVm14nKOGH1M4RnowjGlIkjlfw8JVxDdwdyKlYhqaj
/Y3zM1D+587kVKPZhnFHtL7i5REVGM7O/SS984XNOCdC7Y6g9981ZeOanKsl4oP37wlhcdA0o4fK
XNdXJl2voJhJfydjRjLTQ4tl0Di4Kc9F9H+Pe3rKBq+YgkazaDHhZYy7cnb57VabjPmwiPUdYmDt
oeJc0L0TM9vWVHtTF4GAIrfkh8Digy8y6TMVXFvXsBtRPa45GPoGrR1gUJHQaFnFCMyCq3ZhvTqz
bKR06kO7Hx39M7Dp5ZiwQKD1bB8jyM+JpFqBxwRMcr/INRjNtO6LCBxpJDdRaITlEyyWqSVxyKAl
vnGXvBBT4y9wAnMMmI7ZYTLUX8R/8lRX+iazRXktBnkpyy8qVgWQ2m0NPp2jSzCUfvJSCL5mRCPi
bK1smOhEvIYgVBR3WLwBD8rt4do2S8waugyJo0XgOZxR41hgF6vjEPZTwggisWugrxsJlFE0oXx8
JzOKnNXLhgMmNVogKxgGi24EAWjIEXCie1Wv0a5ZgCluf9giDo+IwMDOvTzYFTdm5D3EakwmD+Ry
pJyAem3sGFg93SwuK82rLJAntn1uKA+Ck4Gt1vGID6KlsRiSc74WA1pXvlpy3ICJB1SLBxc8yJM6
8KAOGzaIjzYS/LCwBdDIhk4/phskNXFLVdBRqns04jScj5Ott5z8WtovXtWhV0wns6InZEvvVF3t
BY0BWan6ZIVV2PfavsMN4IbFVkMlOU6rue8WnZexPEZLpxfB8UdMxf0X4k0OlCAFYdIrAqxAji4q
MUjnyzO7q6m9QBvQVodHnHwBffaB8w+vYzObuLiow5fw9TEmyakf8KnaBGbyygr6YDttM3dQUn/f
jbeG9TnpTxZUgoSBYjAzlg1WjFxEm3QWCr0xQhuLI8MgOyktEFT85ZQoiAVEabmP2uFsDV09/3Ry
dinGPkC3qpUq3oxjY3uXXq20/Y0eSmaEegrct98gY2dnHbC5+zr5E041KfvBbt56paZFAPHXtR5S
nTo138d/tlNlQldYrL0C3OeBDFdt+55bloPMdqk3k05kE7emEyEKV/GNvZowpWI30RQkJ7nD0VFP
7m4CHEfz6B9tDTRGibnbuPditIU55Tcw0u/SkjOfh4bmhhc7XBVskAlXKwShi+7gnQp7BcNOkMfq
ZGfrhAYflpaEPlejiB5iZrnnpnbN+cZE3+qychNxOFlXdsVtDAEY1wn0QUq4Y/3lCl8ApnrQsfdp
DMdtUtJhNUdeKQchJ0lmyJJ6ketMhX8yFK+HrSYlywTIiAv8uPS9N/tK8y5dlvhcD4AJZqSbCkvN
9+Dveg0IKeJOLbpUL55wnwvz1ChoHtyFvGgnVm7Do5cC5vgsqRvOdfZjS1AjbIiDXZkUdDhkyTlm
Bcf6vXFneGJrmUfzcU1Mq4+hUjSoxyd2DCcgY7Oad0iYl1TH6Zp2cK2faZwpC8jJzd1hq36qz0yX
HFJT876FMY9YvENdM9mqbuXY6Aymguaw+ueg+HeCvBT4MmtlHryGXos4sjd4t9Jj4p8h5B/gi/LO
Gg7JbhJ8ge7+P2voJftXZ/UtDb9xG6MxPqHp+VyJtavfm9dPvHknFi7AF+ELiJnToN/PIyiFv5jS
3h905InIAsGeygjforxblYVApxceD6ARSN51da+2QteiY1qILLO0/TxNELzWBYJ6hOxyRNFEvODp
2mMWA2BvRIYCX6gzeABdlsHl5BvT+Ds4IgFErHEVkwTT+iEm0BBVgJa1PYW317n2YO0aBq8pT2kI
VwU4/q8YEU/layqoxN/t7ul9w4QwEK9UEB50m52uIvMPHb4wVV50rK27uCqXglyYQLxCO1fshfg3
Tk7urOOvliFO4rP9lOYYEey5y5tL0fR8bCwtfknzVnTFvEmJgaz5J/FInD0fqLCQuw9bbg60MXvA
YaFpTng7cGpBfVr2OJeP32xE6PyQE7Z+fyB20rXuKe6+xviaFqHd6Pax+kuRfzDFm2rheoNk1Y96
7aS2n5wGEu4q81QvvHuhlPlOO6r55a+odCoMqYAhvvvX0pR6zABRH/pateqY/fWDDMgjkYcNkYY0
Kl91X2wTyh+PPkvtEyLclCNr+3eSQrcy7q8se3UNHV/JSyaPWHQ8h8BTiB2GdzsqnZcJEHeY7XFd
yzFmuIDdRwvtYEf3bhVzN/HE/MWqvzEhuL2dA3A/O988YF7MnQVY75w+vg4ghzGOyAV7fytUPhn6
Yj7dNDo0g3MJqlZlLHaIPlm70PdFBR+BvYtNeEZiJWOumlaBEEik9QIIcH8nTKmx5LKnH9A+xB+n
mg/LhPajEZ8Wuy3ODRaYe0fGaMWMXzFjn2GplzckwTEKHbzT7kuAhbEkp6ccjchqXHIWUf8IZ/Ox
URrgMDm2Ji3I/EQnfSt6TBriI3eoX+UlvCXEZWsDtWrx0270Vl8jV2zX1aKJigM2nUwxY2ciNWlj
gOfLD7CWEQJ+uW5VQeNLaR2soGKOJS2bkA8Vla/qeZDKYznwjGwUzNpoXbTRUhqjbrV63XqOm2rH
spV8VADABo97NJHvVTntskJ1CuNiTU8lcO8lK25RWfUjKzmtJPNpoeks5YnG4YTO0A7G3IXJV7zv
koL0RPz38WnEFPNV+bYrg5D/LdrHBO4sgTSRJZL+feLfzkgL92iPooNJELG6hqXFPMgBLKn/DNA/
9taHp8oYEv/WA3luj1tdONUJ0MAiAkZtbQq/gPoj2FISd/gCfhhxv5UkE/A6qkkr2sUeoGmapTMI
CaBXLYMAg17n1NJj3H3Ia3ZUoK7fp+K4h7cSzzh87YZIoNOR7ekbAbOMrOX7FWKQI7KBOpCcx3w0
McuhEB5eYXHwDfmDL2aBx0ELh6Pbo9Vt0bfUtjFXt3sa0QZoTc9RcvRwC+4ywik6Jh4PcVs1lHcU
B5lXlFPhB74cM4Qb/M6TgvdqUNzfnSfLVk/AFS1/CzzB6uOPmKuw34IjgYp/Yki7Yvkdfd2XfGSf
Fc86JSrh0Uh3GQj1v+1f4k9Adaut1S7CmW1aDgRm/5GeTiTPoFFjjIYB4j14/LezazHT461F5WA/
sXOJ+InBf+dU7XQZkyxq95lyd1Z7wudtAlc6BU3iQk6C0yGmt1eBxRM1knSkv6fOR1uryb2fRgWF
Wz++JqR6cSK1Uz712iFy0mxSs13zMlG03FoDo4BJ9xMPgx8/QZkI0kzEBSljBNDbWRtP1fzhlqZS
452RV8iznT87e2g7wsEtJQJBov6xT+6MEhjssortEo5Iqznk4WXVvex/ZV8xxXKyezXVOuMgMcq0
/J6dFe7GNZAFBmPy9KAhCbuu+x+wjUqz8WkVQJiC0sdJj5bMUiWJb5SYE2zyc7iy2oQ4mKc/yBG/
TX/A+/h4OTC88WpRloN2Eu4XFJ1W3rKhCNX904+XxrZM7GNGwGuL6w/mlH96QD+0NhyZ5RXnC3Br
oyVefnCu18tGf6fkbJzRZntrNFFtbwxQ6awvw9ttNHttUPEl/F450ODzHTseCuIfO3hu2Bawu58G
12ivlppbKP0eoD6oM1DBf3EUXHtCGKgm+WEDPQFulbB+4wVMHCfwnsUrwtG/LVwHrG1g50C7d3qf
Jp9R6KbyLsGk2c9KyDSWZaKANHSG2wbvp1umbDkIgXls0+1AN3Ehb1pG0thq1CFqucMZt+l8/YRS
/fSwRA/sqfJU39EoUl/4aPo7609/c7IAAtqL3sJfW1oDekkXzSRUc/X1ZEcxFiNGhaYT8PQISxBQ
duN7TPFs9pSquZr+pPDPcjdC2wrSQt55jYm5AeCM2Pc3+kB2Mc7Ib0EPPWIvt9HWu4OhhPB/wCRE
XPXhpK8S4Yo4fQ3p2CS16rZSTfFZfrmH7UWv8cvU4JE/OJ1iCUas2rwbZDRxHUmweuk2G3Re0sF7
O2eq1DuhEmNjtMkrAp8IbeNtsZ1CS2EdLrDePsc45T/cUcl3nHUHdsnaHEn+KXjxojr2KUzBmAb/
IiuXbXZwMehltofgOTlhlJDgPGuNSAE8ANYfJwVu/ROXr11FVOA0TklIkCCWotoEn760aJNs6zOO
5hjameZloZzVRpJ4G87Hz82GAnrV59fIUZn6DH88YP52qrnMaATdJWNhqCSCUAHsc1qlLbzxVk1j
U1/Nz+2m7jEE+H82Q6k/+OYnaxlwRs01c4fiW7ZnTn88/qfIHUV3a2KSw3TqB0hNMKnWDJFBWblF
vl23lEA6HqlhFid2DaTfikAmwlWGK5fcjkobFCAc1sTjmNBN4Pns128z/TVq8Ndza22ooGkKyFYY
eFaGOjtcREZLMXLn36Ld5T+iIvmsdU3QhdTqu616O0WoTpI8w/aQg8Zai1ABmih4//Jb1abor2zK
cCeI0bYD17JlFX9Ybaroi8fMTq0j94Jk40FotD/S+LTknM9QcG5Sp1oQ0cO10GWzL0hndp+CHb9u
ObrIP27MFhwylurTK5Hpm3+rqSmC04jA5AOpTN6wQMB/Z8VWmtpHhBNpI3oZExkYxuRrHO817iys
0yACg8ltP3Hg7yxocOXY8Xc4JcWxhYUeMjZamlRfHx4z5MV5ZZOS/Zjb/voSWweMCC0qabChkxq4
cOtPr890intfKXgJIiKvWXMOcBmcLJtUfA8gQI5hw0b0jBoawaos3qV1MmrIWEOXqOsZNu3lmaA8
pbPD+QFCDKcldabVMwy/buM44aSPSS+6yd4kX6LAqu+8RDxin5U4BI8gEIzJTlE/pgfhwnn3KYcC
jPF5zKR+9Y57YsVF9yAxEH5CDy0gxeWch0BAU6bzBlyXMi09x9L5RQoN20Ti60Cqsa/Qz1crJOCX
QFsELBQwlSeddeYkopHVTfXqkcwACrSgq05wnQcsa5qPcwuQZ9/tyCth8L+vIAL5cPPmkJ+IcPOi
YBmhhd1wdkZ9py45TVd0A+KxTv0BhPSuADAWH4s4qjYqRauKK4a2h5nDVNSW4PXKj6IeGyxhqhC0
WUQb2lp3Euy9gwpZ2tVQ1GD4fdG9c6Zf1aFAmoRbEWrT0L0DXyN838uzmTiAFc/VNMzuyvMcbZ83
AjF/2OBbx5H5/dgVpfLgGMv2Xf1VCSjsborC/5UZ2g3aEnPrYdP84sxFJspCUGNEH7WYMh7CsGiT
cBFXlU3dw+3hHPdhDLYyA19EIYIQO/KH1NYnEte8GUWetTroDxM501D3K4a9LzC6d5gBJZ2OOVXS
DgKE1gDU5jRyNRRmxB4xSWSGo+IzbWytAmTgdLNae7OlBE+4ZlsTBYlfu5DR2otHCs8HrsDU9NfM
LDVsXO1f4dtbiwjRadJBRPlQbzZl9XskEUpOgJ/lCC9EfO7NLJJor4VvO7hjw0xZ9AVAGUplPRv7
gZM6WNLcv7Y2tDPuGo5Q2c+DVJAnb0TxqEztNEcraP/65e2+lvpfjVTHEQ56ArQH0ggGmIKwY6Vo
l1WTESrcmSTeHVSQ1fHo4fe7/gnSSXFX0Ij7zhSTxiJ+wduQvPeUI8Mz53KR/La+UG/lnonEI7+h
LhyLlVU105GEs9hOoPeIGieDocRC2MoQEdYaGbyKaPyM5f1C6ScOwIDsU81KVnSRz5XRrgTm2SwA
dizgoGzfoNE0l6q65/YwA9NIBW4oCW2oitfG3i+eZCzQJNVabQRHC2ezBOVb4kGzp9f2+OYNDT0i
ewUvT6twltX3Mzc+HiOrNVeAfmIPfuMj7IcNg4UNArgqZm79TsL8YOGBMFXEZlkGIvQ6Q9Kwem1r
53apZaoIegRhU3VF+EZw2+TIzjQCZM6lQCjxjR5MskFtdnzOJyb7PyAwORMQJtrrte5Hm73OXDtC
K3oRNuPliTGF3AST2P4+X5MjhqpeTZ5aEOpRcYheYrUg9RGtuAiTqqwXBnwh52Q1lKoRula5e+UJ
cSiNhByofHNmtmDk1TfFRewU2g/gF/7jgQavJ1BTNwFMKZhLs2wPHUJjVPcjfnwdZ41js/oUstxc
kEhk3jT+3QaSVL80cCwBzlQzNoGt00luUhvVW4ILsakgqfMglSwXH7COwi7C44GrEQeqyuGNf63r
A7vrqabb2HscOhKGOogVsZy0LUrLPcNICHr2TuhIytETXAW4ccnPSjqlk1BoETlWxsS0/sKs8/FC
rIrbYdWy/aYt4eiirDS1Z1KNwo1td7QTBT7Zj4GEEyiVQOcv7CdLANi7nm1Il5pLGhkOr11pLbCW
yLR6NEYzFMl17lhLgID5Wfuy3kjHvtm+Db+BKa7HWgkR2peFKUDyO7qnm/vDpClVGNlaMyd8i8LN
zMD0zhk/J4APCYgWjVpxETYLM0bPpyNLB8174rHY30IF8yuurp7HSxgR/y0TiXrlw/0Bq9VCP47S
VSWn3dXW9ZKjpK5YiEe54AAtPoOnpLaUjJ17UqB8frGBrN36+Ie6jFxbB7lggRmkoQF4+5baiqar
d8M7wfijBnpuXiyCF36eQIBqmJR1Y5rgpMqw8NVYOFLSsmE2K1Ynzb26tFW+SCLkh8BLhRLC8pAE
fbOoFjKWQ0mRNoqsiLeMLL2MgBswKjysALaIG1V4azqvYEl3FsMdTDc2SbgxE3V3UeO4ZKojhsMc
OxUCu0elxUVq6Q20p+YcrDsT78fEzqyzI2Xr+xi6yvY1Vqz9RX9gFTUVjltKoepauAHK6VDrY7pO
g08i5/YEwlsPlidl9cC2IthA6lOXe8NNNQYZlOiGSGkCdkxK6cTAZIUJ1XLOINrTUPJfzqKEjWBx
jCgL08pXFOZwO5dpSLz6FlIvtkuFeyQ1CetmeG4VAB2xkvJpmwLCKwztd+ZYzcXpIizRq2KntCYc
7oVBj4HEbqFv7KlD7oii5UidgIgzj7r4aQ7TZuNNnsRKaSaCgGcxnm5dTLzHgBNKXHRy+1jl0RAj
qr53t+I4c7AyYh0PC45a2JieJERmO72ZaUt985XTORF0FTdr3hOvS6+5PGJq4suoObp9Z33X9dPr
TkLo4X2c12v8dP+E376tVzDRn7BSB4tqreeRAPwUcud2jtCJnLTGb1VSjwfEvGQlBTAz2OSeV8ti
46N7PvwjRWq58VAf8/qkUIhWELkNgQh7/96OmGrP2MPLrlGVO6GCTmLrXVw9RmnqvsOGmgR5jaDj
RQ61sQDqojV2Bt04ccwAbKWNTcN3krUgiyPKXB33UhYGFJ/rA+Btmu/zuyePoL+xVbPjxIUpV9/H
3eNbs7+5x3YJ92wiNZB++qCkvKEBVrd8SXYcY5Ejt370jYQuvwUkUfAZ0StP66LX9e+KwII4Oe2I
NmO/4XCK0oQvuAh/JfJSlzIzEZZyqIXuJw7Zo6NhVoalrJiEJILyWcjj5U79UdyYUPdbMBnaJXDS
ehh/r3JPM/BlBjKEc+r+Xs9pS4dCHk3DUJEA2Gxy+WRJ0lqm45sRxClvA843ZOBkCzTouTbyfQ02
NmFiftoH18JU9BXryoUjU0GR3lF7+EH5Kn0xAVYxmwFJiSDBE/diJEZcQCTCUzdJi/NoRXoJYTs0
CzfYCywJPHYuGjAM3SGbFOOCQMjVxZkj+GD4xdyNSKrE4fq+uKoex8RwbTjzxmQ9Xas0c9Dsbrfq
wPchw+0eKoNg8WhjKeeyHLystJ0IYeeyNP+2aOy9QiZbNnB+DRJZNoLCWyhNkRY0JUdcL9yhlnjY
vPULd6LHil68X8SJebLedhyzIviTdz/V/fIOwYo0693M5Bc8hRWyqQ2d67iRt5QSdNtC6mU7K+vy
rHV18hD2FVqsYZS5r36feVVnSNHYGhVfpiWLqo8irnpF/Ml1WYC4XA1gM57t5/RFPWLyNSZ0jrrZ
JhsheHyxs/qXAtQpOamlufd+B100Uixtr28OzSh4IT/JuoeYEBcn3X4DbrJEdwahgUVl2WEjqXAc
HwODpre1A6O8E1u/Dp9Zx59BJsEHXU1PliqLngpK862pXsh4+P6uk3zbEc7mT/zeZ1+SET8wPkFX
pzdp4dgkLNwc/A+sg5zkYEkEgqFYtROQMpNwWDi9OzVtFYvBVuM7KtQVhpWG4c17lEJ33arzp7D6
SxP+J7Iu1ECBiHb7ol0TkR6MfJ7A3ExNNJjdBUXioOOiAnPxiUh7/sB7+TZ8aF4K//hox9vFjkVe
+LrTQSUJY1TorGaXMCN4C0lZ0gbj/KJhGiJlLm1oT8hgRCGSF4o0QEPqwyIUnPkd07gy5hZHM4S5
bGlHIeSNhUC174hdIN9gNe57D9U+Q/bLYtZZQsTxeUb9Pxq+trGkxXduikGTiWB+L2WyBEjnPFz7
q0kGz6Xk2Daq5mp/h+jMO8Uic8iO1nMpNcmr6WpJPbc94oigVKIukEGT6lNMkLk4nT3jfsInCML9
pGlcixxFfoP+vVeGiRXzkKi4zoqJKWGkRqbNg0OwsV5fvzgHTXnn1Dlr5rjhOxIAf+q5MMEh+J5N
oP0IRrmlKsR08Ij08Qj7KYfFkZua9ouCmY+Zk1a3moWFx6Gfe3f3T1CjwRxjvtNLZPTEnFqb3Ml+
6eCA1sscHq0xR0EBhr2KdvK1av3bXpzYLm2uzK6fQKO/MgBw5JlrqTvg1+tpjzq7VrI05F2pXU7T
3Befk8qfz/Jzr8s33Q5AreWzyqt/wS4R6M3GhsEX4EsNZBjIGfz2wHT66zD8mJB7sD4ZwiLhBIJc
nAgbtLk1W667BM5kHUtHjYu2eiOf8Ga1obbbXNFYZVd7KR3MevlPRmT0Hu5WCUS9McsZDmFvkSma
Q1XKyGPZ5qwDJ2z/EuMkzcnIGd8k42H3v5TxWNskk0HgN3G+4j5O4eAGQTeuVsFklTThg11CT6/W
aameVV5tP3hfvLgMjhajkOXJZk1YLCmMPAWVm56CnRxsqZwJeb4ZOLyFhthQjcrRg/Bkcrm99bmr
ZyxtdmXzd8wQkYEHFxMLl3sKKUkRVNqLivHgA3tFgP6oS21dPFXe7uT7mYDfOG2DPDYEXcEb97PC
K8bI5IVKstmPkJjETajAvrb7dpqdE+6yFX1g+9eN1y+IQK1XrWdjSKnrOnzQArjnlsc37ZMYJfjO
UHwFnr1XXP/OEgokf3YHYOIpphY6FicTlOPIE5n+3zprWfeNRqTCEavntPZHBCPBpDZpsBfHku4l
qKzmq93jj0ABdsNJVe6E1xNpBzUR1hPmHF7vMxp2fRaq1jGOOR8ssMtTs76csgNo+YUnSM6ZSBeJ
YV29TQLD4O+APNT5tMKh0+KW3Fbf0Ej9cgQW9zKTqI222q7QfDHUJhZb9mVZK5P2QppqOK5+7Pgs
YRuDnknKKsQCjNOMgPcQh6LCiEEPAklKQKD5z+1GwW+LqHlMBWsHWagyedEd1+jDFEurgHz6BVMz
e0L+mmBF1YTf0CVvgWT3byaR8eRaTYDQgpICPxZJRvJVXumujmXc6kSk20RCBo/plINtLzdQxRPV
fcOjWj0TeccgtxJavzaQ48jz59gQY9M05KX0Cb2kYyMjTB0r33/CVddhZlF08rXfrzkpr61f6o/V
I/dSzGrTRurIQ7nLt+DkIWVe8K3QJQb56832cPh54RYDyYUKzHknKddVYsZMIdP3SWzQh7i9MoQt
moy8gSfYrHAf6i1bqXUbP9k5Nw4wOHkeUBSlkQIKvlg9xp/MHTb413c6T9ZEzS+DjmAnmg6WF+5Z
8zNHckkX71AOSg6NxoS9Th8kweBPqlZbK54oviNtBH0ZQon3Fvmt5Ox1TF746C6iU+eTtoCzYQmV
lmIIiFFL/E2wxBWnF4slFCDRM01V6r4q9wCfiZpRoP5Ylz6tmbP8hgFILKlqlxoLlbnmwSAlvcyI
Btrf/Fl7BpsPln9WuT3WTA5ucBC/FGkGkgRlfW6VubCtQYT48vMNT5tcylgrEsVuM4dL6op6491y
HEg4Di1Vz4eOXdqqNaFMBS3bsOqFAa7ugA9LkHhN4s11G2jD8dH/OpkrNiR9FpvwVTa1UE5nhXk0
UJ4VMhzJj5Z2ZUmHsi/AlBQuGDNwEgM4K1D4/CnqkXw6XlehPj8tJVLy5qeCCyO1R9wXfJ9zXkRW
051ffIwJ3O+S84ZywC38Qg8ybm41JzYTFi7gnSmXXfwgtBbImJey1wDyX5BOkB+qbVXEYtFV5wnt
WdCNW+aNyip33oC9cF4gNv/kTI8rVOlY9ie/nEnv5MErBd4kcqUo9h1eTK6E9LcJExBo5kLFx2Y8
yBAkDpHQyyBb8Cdxu8tRuwA7AA/1Jyj4Ph1ePHEqOiFhC+akyG3meWZOusY2wRwHkgD/oat2UXBe
hC/bOcOB2UzSvRUnVl7nqh9Y05ZRSAWAwHilXgx98V2yIR/I2ZdJoHukQbpSCEDABaBtRySRahJD
cxsMzS+PXsg35WpMX6zZecdRLtfCxGCekTadGL/DJ+rwIUdFi+FXTiyv7cDL6NraVncBh0wOEtKQ
vVE6z2WCPjdFrRolzhp3vQcG336AQG3/wbHAnmtRtyHdRMphxEa/mBAb/4wodTHPEgm7I10uqxPc
ZvbYvJX8J8cC/gAB7TeaiAZ5E2ThVtZkJnVojP2I89T+g9ZBk9Qy9OjQlx9oQeQrRb1StIOH3O9C
mqujj04CSb1L4t2WpLO4R8C/hw6DrGgf7kqfEiyPDWhY+yVFtqNv8lUeL1AVP5q0uWJ7dkwueKdt
g3ROL9RjQrumUBkWM38argR5TdAPo+DKgJL7Sy1XglEXsWKcTkd+IIWjXel4gbbATjEEo/AjRvkI
JpYnBcTB4ngDgJgyGrt6qtSRzwp3WCx87sOib0FVxVtwKomu4LwBhQv/ifY9vac/8oNS+8A9bTr5
g/uZUGGn1QuGlqOjj/j6YGwCIb86hpxv+RdbBqnvOjloTANokiVQOIQ7RYL2o6t7AJ+6ndlcXfqs
RtVgsLTjox0eettR9HIPQmiYa6xJyt5c3tF7u2f6QfKHibntrVd+/GoTouuLqrqXTccSbHKjRhKV
9EN84HIvgR8QU/51C0072YZPANPlCj2yJ7wAXypSFGsSdvoS/DjEq1Z0HI2FB+4Ro2cAg1EdtSZ7
vMKiUdvyonwANx0+t85J1ufchSA9i9YMFsiX0n9CAKPjn2vAvG4pyS54Vr1bQl1kd5z8tCb2cmyJ
FD05NZ5JnAZ3p1H0o+eqfOt2Fo3CS468eGOVjMlwuq+irz7GM3B6ec3RowDYtohi7XWQ5fgN+CIB
J7HeX+vIyS5mms24xwTFS1q4KVyocloTkGUNoliWB3V0gvtY/In4ErVZ7T8lunTsvprXYBQM5Asm
WL8LEVEpi/6BMYfysIC0+cyXzb2Yn/PPQ8S9+i+OqNtPb1DmmpPEsyQxMVLUfVxZlLRU0nF1eOdv
DfjTfKOud50LTnqVvJmDzppfZRpnHYGv+krJREejCmaCLjZzIuCKvPTLx088L2VyUANGGFOMnYFc
kwllBH6PYRKTkL91JJwIHbHX+RSOyShzgwPln79qYdrOuhfoHWEMJ8oBxcxaIS82xut81joh8me7
Y0tIY2UXdzjtF6suI/iEVjKh54csXwC+79G60rknlJsdcTANVmZwYzBmWDMTFWzzrSPnlaghjyXY
2a3/Oe0wErzPOWg/Zapjjn4GEfuorPcugOmQkmKLMBee+TAbV5pbDKqnsPHVqymPvDvTVC+4qtJ/
rVUFukRGpzCdN8BasrNeASeO6/ygyf3vyjs8+MccSp1rEWbXfN9ng/rayG6GoelsYBqL0fabx8EL
YIbtYn8eRzYplU0nIXuiFwun35gyZQXNanz27uTAiYZum0s7T9FtQ89s9Iz7mg07EbzS5dodRArJ
4GnxfpfRCJWCLX6y5IGC7Xs/ub8CmYE4NxdbeJCy51G00Acn8k3RYBS9pUX9mdXbMsWCyp2WsSQf
hMm30xj+L8kACZfmXDc7P4TEexU6gkafh6iHvGig9b+u5NTfaVBwG2WY0bgoFskIE+Z/k0k2dOuW
03cpuUftc+t76v0OLGNv4RXCvJamCH+eowNpSAS5rdfRpRHy8lyJZlhDenwrcpKLteY3D3UTvaNi
WmubwR586tyU59uJjuS6OIFWjbBRx2U9qikvwB2QyHlBsfGXSt2KA1n1Tvr8KV95PXpCx/uHBd1W
/PAXAsAMAl7GG5D/8+UYiuYUwVOYelHklylz8rdSjOKuywBSSPipu1afwmayKv3nSUFthZREgMf4
qpxOv6p7PaBcL3e0uFGIwW1+zFKAOX+f/ZbDNbpqZXIy6sSkBczoA2FVNN/FuV3skjo8kbl6f7rj
+QUgrbpRjjUzYzS1AEYoWEoJ6oNg2Lfkww/W/HZYSt/eMKOTt5Iac1ZZlUlymAasIQzLzfVBUykR
V0oKtwJ4ROkNtFkQ9nbYDTiRn91hOuCRQ0m5fZ7BoKUGEtQN6/wbhgoCsRuV/uIEUkS6gsqEJm7/
yNzsa/5RSUfpd7pf82g2xoOu3bN+yqKJJzqx2wYsw2Shk+GK9cWsotZ70WNpAT1nU58+Lr27NlUf
qIcY/xNKjhnIbrJA1Ubezm0aa/QnvwTfzFgvC/bZUInc3Hj/dg8BUQ4yQWdWQKW/0C07hQAyVj9G
/H8EiPQmg/DTUlSEmeos2VRBuf5E0ta/AuCrdbjVG8zEs1AsVzBlso0RlaTuumgWJqx25NfVbQFb
rhxnMgnhV3izOy49VEZ4UiYAkV37WzZXVjAfaBpc6QAFkwihKz7RQuSDuRi2XBjFr9l1zfGXM3Bo
fzW+Bl2LPgZUcu5uXEHFzfUcdnW0t7jw5SZkHyxf8PfMrkeabanaVwTvgWZ+5t51++Rttfyhq8je
YPfCaoRz3wzTJa/eqGvwbC32Df1rMdWNb3YfoEyXck5hZ6cptUXRImxOsrbZXSOPTal+hORYrkq5
6L3/VwPmgYrZaqqbdEyDFzEyOJJ2EaAUaYHMEkHPFvUfOceZgind4NJ5QkIgz16y6DOtKlGvxQQf
ebfJv+PTjPAJHW0DLCtdt6IlrvhkfFRk9DLbAb6urLbWomjHof0ssmm/R0s7ukt8AdVxsPl1ieHE
nRWMsn4jYuJOzEio9vc2I9rMqDBAKBKPMbY4d5uhW54+I3KA93bgvnaXbCnPPtJS45mIUU123KW5
WLLbY+Soor+zCvmdcrt8qb0B1V2lzFguz1mvrFcU3EAbbyzPQ0QH7pEhWSrDEF/bO2HSE8vT41TP
unZgCUYc3s+uXz3VGOpGTuyJnCvGOGBZx99jBOhpe5yTmsz99i4H+HAXUYsemB1FlGYyqPe6nvCM
eTfXCzVRH8axDfV2I+L11vCwvkiNmwr1CGU881WeXulj/qrs2J1kOF8mieNW1FDrPU90KLbhjv1j
FMbjsbp6UoepWzN7KpZi4vg5CX91jaWc4E7lfWCAJeLWzzLSA+Z7xDIOEoqb4+mM+myKHVSnMSyq
hcFLbOdA5o41uIehmJjXc2zyxTU1SmRCbMpGpiRhoH57wYTSMXQDp4q7gF3NsPJ8Molx43xaj0ws
iIY8ot7obA1Pt58mmreaFicB3AM4/mOKid1QHSv9jTbDa/J3Jt5jOsm/jBuNoPZt1hzvpfLnptwK
W0+lnbpbTju3ificlztFMOnyHgBl9vqJ6+/8//Ecsz3wHmWQObp4dh53NVAU/1fp1emejgPrDYNS
ot86M8cWeZKPa04pbRNOviMnSSJI+lAuxUDSPad2MLnGWAdt3MCn46s1aY0aHIrtSLWubK3FBdTm
QooydMpYQRbx90mJwjdzAeEVhFH+23/YdBeAgG7VwY4BsjPSbZV5B98/DFDdoAwS9JbThcHCXfO2
GAO7OjcrbIsI4cMQPY6UBYEeaG8199CekFnjK8R4fyh+8O4JmfUjcyqQZMmTXBTjEJq4HMe5orBc
ioKgfiTa58Mm7mB9Q73VQWZgguLodN/CUuWPzEFniRa8YGpAy0Vt5WOH4J5wNqpXpMowmUcb2PHX
GIM4R6IDGF2cWturzEgGZ73FAv70HadQLAgRTQtfliXA+/JIAqi2z5JCN+11iPb9E9IYfCi+U5D5
hLYgYttSiw1A8aZcor0hxNk3gdE5EekbhIS7MHEfg3x6+uYBGh5hs5xt6EodR9gSECWtge49z2Qk
eHPinEEduwg1IWGMgJ2v05ZuUnfa+UBll5zZSDFcmO2zaX4Q+DLpHqLzr2EpQmxM04rn2mnBIKED
IKVFkcpIeAb9uOln9X9bei9Es9zPJX1rNXpKY5cRsMHwPjJl54rXzqsQGrnHaJi1iypeWSbzUU3S
plrKx5XGTYC2Aw/Atl9MOsRrvQ/O+NMwcYBjyW7wZdjG32Axstkeh9CqESL7MlLzxdoTSXTAEUOk
jFgOcn08WFE61IkZlqBobEUCqeRpwiBAHoz6kOr/K3b/i9Vl8W2SZG2GTYsmzhZ+gV4FkINIl564
w72jrEt0oGqFlB91/ilVXEmugVruzKB5FzW0vlCCWvJQztQGmrisENqAmT3V/6Qg4pA5e826t+r0
U+dw2KM2QewOnoh88YUpc27Y+O7Z3AYKWLxb0KH84AW2aGhqzk9akMhNjxd1MN5DGBDkuj7j0m1Q
x297pGWA2Un+j2yJ9989tqPj4IPMLeCQRac1Gq7VT0hgltD8BzDTQ5d5wxKp0Idjs4WFeuB74KII
LFfd84tp6wMVn8Z+ZCGJp9UAjLZdW4tcFu1eIBhyQ295MkjrplwRrNhAx/k7oHOch+HD6+7J75Z0
WEa5UXDjzU/WdnNpmXD0h+73QbyB2U37/oe+N6Sfn3NIDDJ5OAyTc5fFIZSuRU62T1ADOaTcR7gP
C0CeNo611M2Hbu3rbcUChx26y6IXGPDjSkW5TaMyxjDDXwsh2gSCPNXKhD+ESZa+J1ZXCa7h1wPO
qdpsuB5HU96hedJzZ9UgZ3iEZG5aMOE7LJb8bQ3dytbV+n8DAnFn5NT6H2fvh0LS0kA24rTc/LHY
oaEOraaB93GHcy+hrFgNIkaRwxtnj/D2dA9oOWQ4AbWnJzURy+jODeY2sDNiODfmAjVvzK5Flgmb
dnkPNPoA0Gv8Lgx32K1ZDnj1TPqsRL97/F/Qfcv5DBJ4WXHG4ULJWiralKyW+md0sutbXUnNj9SU
r5UR23dWRjkuds8By0QAv96PANakfD+DMmdDzzFHjUoKzpqorfmxupFGK5O5E4kbJIsDmLquXeF4
WQsxlRB8UnoPllctCY7jKoWPCOOjs9R+hvVrXrX/q5XK4x65HffUWULRlaDrWZxksCRArq5g2eYG
3aY7ntQ9+rZwYcYu2Glx0RFgpgLmqvnbLCadJe6nT/r1Dov1qh02TxDrc5NwmJL00z5ZUKbhsLtv
8wyG/kgkNtM+phCIu6AJ2IamEXopqMguSmDGaDqo8c+BtdBdyJVedIETNEm31UqVYf5JgHnvhb+q
WNJ3sOzY9okbzflOVW/cV0JTHsZOqvBWNMIn0RuJb7aKACMvEtxgidFhwz69vBurR8GfDOv93Xp3
jEnECFhBY2hWG+srckSgLRQ4xrYt+WdHiZs6cEnNqE/sTso4vgtoB9vsLHGJEylssGrVc4IxBVBs
YpJWI2uB4ltonvp33EpCy5zkowXITCP/CV2jaBI9m2dm7+x685nO82NWWg4Te2HRq8+1B1yw1HxV
R8E1ZLUGZuFfNRVjrnR5GA7iyFzIQ3jveVf5ON+LTTzF4sigK/tolIJu81KIJhFqi9P895HCbEMz
dxO8fbxz5VfZNAUV1L4gZAYzo0G7pJByiU5xYhf+BQ4B2D4pN+dvIXqxZhDNIq6NPrlX/u2xp+IE
YwTTFk1WPqRe6tbf7J33LEfSA9uRKh+jV7rzqy6dYK+ynHuxYqG6aisCDiYV+6HnzRGEJ6STC3zG
bgbM7IcCY+CP148p5T0wDLfrtE85IIi8IgAvBUGOrq1QHezFY5Lei3xbhDzm3FTbhgmViL1pMdkO
GVYFfrIgr3C4tXPGDOgLpB3g37JAoxknJKmkdiE8pItkXcEYkeoeSbnyE8ezRDNebdGSybYFNgHC
q7lOKZGcEDHO1BCieDMjt8qmXWU1iZXBRD36HZwmu8+vC+7DbM89aQXVhoLZ/S0ihEvMCPITFR9u
gzmEnxZ1RFKhxEKwHaKgNhcYK6lxyugJOClIUYtO5grx6NxaLe5oLoQPsRjS+YBj8JdciX4TR2PV
yBuI5DlaLOWs5FuhiWxBR53y2gruOBXtPM/QcJoOfOsZJsNyomV3H0JpDtrVPpoWGKQdVFeDzLjW
PzxVbDCLkKajUgQ57HSNOmwQVZF3BJiGee/KxYfY0rHsi+BesQZIAXRlSA6Ch9YWqM7ZM83gwVoL
BA5IVorTXlYhogxXjAN+qKcNhvHp4emLGJ/lENiHE3oNgyQBfCBd+E1SOnFdtuGNZpgO7yuZmawq
Yf2HffeD4QpOr0rkK0avAc9NFD3E6oORi5+WiIbT1ZrX5Wjwla9pGPRezxPv/elFR5/OGrzPMEjt
Pj2RdG0UB/Stus4y6ciYB6VsTPg4ty6fGkh9w+1kIv86mL0gKtx6jhxqb+spUS+CDzdh/vvdse7U
DSGJk6d1m575xVRAAdwk4Uat+3cb00YmkWrl9VzjmLGCZt9KFH9o++edx5s/QtvhUgSTQf62sB60
g6rBQ93qeXuICiLn1dn883pTsLmMqYy6XvKVzE3zHVoxEGRSP9lehYmjtu5VsxekC0Z8n62d5LJH
Uhb7Eg6NqFljUvuaBIUqaRnX5g9OwIdpPZGd6byui9yNY7kKvvIeEo/MtEBRAe/hHUWlsm+o2iK8
v+mDcJ4jmawJRtu1aGC1YSt/dHVsrST4oNp2NokS49C88n81fKM40xVhFyFVFBihEJROMUEa7eXj
TlbahyJcckZm/oGlZQzqk4RSSRc2Au2pZrd++8076W7k5AvSTvHpS4L7AiIqsALvlrIrz/fk8xNN
OVeqef0zp834s0aWsJH/Ca2SY+sJdX8JAP+vO/V67wTgqW2n1J1CygJemCXj4/bYawUk/NGSOL4C
oPgd4fTGFKFuzhzThm03eZdzwENBbBgGrz5Ilg+mEJyuK7KjEbZY9DY2l4GdgDaWei072QJ0bTHR
GvdHW4Q+mOga2ufNrVDddrngJDlxmlqsDjupdky69/69MA7Ss7618nhlagB1SylVLPyOOtB2n/F9
k/ANfdz3y4bge8Q+bhVC9hax3e8JpKcbro6pzbPg0moluVwNsX2dXavhhNaWJoxHzD1Pkt8mzugx
FPZPx/ha27dgT0kk7J4e/XlRiKyMeKy00FA2RKFvVAIdHOJwWSkEm//Nnx5ReugXbpiO8J4+J0M+
wXeJC40YlO7y+Gyzb1OqiS3dAxLKsEoawfBYEPIitmwyR9mU7KTr0qlF+Vjcn3fz8ArH94lcUBwS
KhX+tZaL/OqqRrHfNrDTmMiJLmZD5JM3TvcuhBVJwfONYKhtO6MqwSlW/s/tpNeQOOTDNkbtCSlq
LEIRVHH2/qWNWLlo5RIK3LgeKDAPsdVOGNOxPjFrbnBaeVy5oURrsii8dqNtVRLYupd7JfmSlF3w
aCcFdBrOmoxpYGGask5EUcHjDFeRrfEpmF8DsoaF60OsOWCzaIA68ApPZ9TuD+2i9J7gTIQDr/F/
bqQz/OFWN85VbrwVRAAZG7CF67A6UpFR0KD0GM0PYkm1GOty1MEmBcuWM5K+PjtU0wr8YRGpYFXs
R61qb1Inq6/rQ2xj05454rVxeVK5REb7iZ34+w3WN2dCiSlQCVQnsKTdHKN+GkMjsJZNHF4FijB5
l+9LLx9BURDzSN1dWbitvgGwyTP0f5/DJD4h6gobJRGbmHiRZk5YRfXaNaIEcMf8449gQT0Q/oM7
JhE/dC3L9ziEF5g0pqSXyjKPwJ/eugRNFCRNpvZYwTSzkvquFAuzQZsvJkcUOthxpO9mlcJT14Dg
EjmEYPdMRCOws9lTBHd291JaberDGMbLS8z6xuZkMf5kUUBEmmYS88GBc+3Ag4HekvptdsC2wsVg
y/Jj/cHeRgyeLTSYJJjw5yMT1JR18Kxovk4c3uHTY/uA0tABpBoofli4xo94US3wF9dEaiQtRjFI
p4VPNOXZV2sPDvjPgMa8bQ2RmCrohw7krOXHNPONHrOn2WplnDiLCsMnvxM5PigQm/O1ERsYsbQ/
swSVZgk47rcwo857xy1PKVzMwmHCC/4rIVm41xUyf+MqMXBuzxJQZmMs8XEpWzp8ywWDS2+dQwnX
EKWpWzvrAvmBezC7UZe314qHTr2xgid8eEeHRTWpNuihhCuoT9OJzgPy+ipA/pB1SmhQYDVbGfD9
0wXYDHecLvb+bXRnnEbjTylP5gSEIRc81fsnSz18jsxdFeHvaAZ2H3xiDy2ch2FBKg69KJkotX1U
PCyP0Jb+nat/Q9j+SOBtDFYAzlHyXD8wFF1rv2C68Y9IkQPf4+ElkbmUldxFnkMlP2xq2wmBmEgP
1J2W+Uq01NOnsz3OyfRalhg/pNE7wtFr/cAM3nAuSCyHMm/3uf8lqfcyIx3ZU0YlBPcY780MArqd
TQ/6TLNfYadoVI7J+98LaTs77JlXQ7ZsCu7kPkeeuwRJhDAFXDXtuviu69Ya67WGs4E9Y4ih7lgn
qZf5sPeVG+8Z73YAxEqpkgsBZgnl0+QM2llIm5uJOllAnRCVsq6cu0ARy6umg5lnVEc4vweHoYWs
2ejpbB61ftBZR0Fve3wd2TzFvifEuhbzm4cvBOtrZSFqQ08am0S4ARCPT+vKQN4HTtvOg0rMSSvl
sZWd4YOH9DdEkBfnyGNrVYFst6oD0QUZ9pRrUMnrC+J6GhRlEFpLBz6shaZ6+6cgLMwIxzx/sqfj
2ofYWNbkB453hr+Gkjxa1K5JzaSrOIRRYitoVjS2GSgttiqK29zFnnujjn1k7eu0noSN5Sq5cDee
C4FtKsS0Xx4dJMaB3Cp5TpBaEt9jIH3unM7NpWhBjJFaDb85JJKTe85NDth0fBVFZuoP41BGDrHX
HWSBv1QfQWQSW+Pbj5AYU7snk2pxQffkMadv3kB9Ai6LSUu0+ymctg6yVc/Z9w/imQYD9MFBmrZb
LMSkg7QSp4RtbiQHPv1FuQKIVlp4r1hU+TncblalUkRP+tRsIEQ39WMyzFOvCEE5EIDoR+ucSqo6
ZrGHbeK0NN30eBWj9MAqGTvkRYMKxHSzxM9gYurcPmw7hWopzuLBOIbuImLTMua9vCU+//yHOQuX
dLZkkjHjWX7uhaY7Uu1wN463C0xwHb+4x+0pv2izKuJH+p4vFqdaHsh+SeldqDFp37vv+M/6SSxw
LXkaJzlV4BWr7Ns79xipKlkL33nFkFc8UiFby5dI34Gzc0MftXv+jSleoSyPIkHOw7bSkV9AZlDQ
+aB/blGDUgVwjUqxpJXtt/poNub3XSLRmgq8+aRyVekUtaHQuSuMgb2j+ykjG6YlKdFA4ciXFFbl
Rk1kELikJN23TRVqaf/B84SFLbsIidS2V29DMbQqz+e+mYf+WaQzj/dJcbB+mBK3e2b3/+UIWl41
hGLmBI3Uf8DziVJLTFpbAX8LbsjTu8ibbPPXqQHsk5yNxDiGmE2SPTvurbQaxx3akrHpkrvQMZ/X
kIIQoC98wFE+gdPTC9qCFbGWnowyEnYtU97IyIwaVpgtpS/Ru7CgZ6r767slWizWVvJyZB1+oFtg
SNb6RzayIGG06frtWUXg8UjwZF8PdSRylZ3kWEdJvobv6HolA8LFMWn8RTEYI2KtD5KSKYwa61Gx
0lNO/pZy5+8KGRdd52tCnvBW57cDAnZBGyUZVv7UJKzCzJNqvEBBfPBmDh2EJ2DeaSEQBLRzzZPc
ryIKlWbsxYRF8qjhakQFJJCv2XlgrfXHUy05RHM3DpLtllyzUGfIj9wShfPAsbkR+AyCvZQRH158
hBM9+bjwq2ShFA1XuVzOcnKxrmITi+jo1F456Uc9PRWXL+A7hYyBxmPtuONf1FR6GrRU3dBLIdTx
vKIulTdoKtS0JACjn+0HMSm/8lGWxajIj7aYcJDImt2dTHCf+nH16fM8v8/1hfCNGjfN+I7ukWxM
oeG5TNPJDYqb14DJOiOz2nKgKkaccRwHw/zg+ZS3GBvKtNDqIgY1AHIedFqGGGnhgUT7kuhN5HK2
ikRW2BMgyqySWYIuD6DUV3ZFUcK/MYJ+gFQmmMlbTvkyALUZt9n7NnKMGArCbwLNs9vydMWlnhLx
rjZeEISDMjuQYOaTfG8aZEJq89Dp4Eqa+HepPaMPbB/w+t0al/6w6nR5K4imTdP3WtjNAK2JVwrn
2jjn5OUxWSehtfKqhiyKLgAvkws4mzviarN1TF9Pm2OpzOb9N6yJeXgMCQldn9ttKWLCtk0ht5aj
G8rH2m4M8WmEYEkLacZgdlfmQ8mfQLG/6J7aYxO4Nly+lw5zn7E4wX8NM4DHfc9g6Bv1NVokounc
qNhYZd8KM9M5pGBxGAKXdz4tPah5QZmKpXM0XRpWbM5CWEuGI0bXvbOXqne8L4DGP0kPmmc/5ZD0
iyKqyuilZiuY6Xm/N5tV3tIJ6Xj2ezVRzQzDUOkubJ6x9GtuwBn5S1O5x3JHkICgAUtr6Yxd8CPH
bOZ+Q+XDDLNoQPvtSZ1AoxxHGTdtGeKgmtjwX5Y5t44LXRKEADUkCDh1NDFa+V4cU/2wV7r5tlJ6
FmgFSprUqcMefpBR/qKoN0CjfJYnZC6K8C6MY/n0RmNIZWN1hx9G5/xKMLTdFtsVnEsxrxPLgQgX
OjKxEAiFl81ecE1/JDJuKsTwH7zHBopJtX4N8NOQdURh+2NiMi9udXPhX/Qxmv+VhIATGHXrPbJx
p2PUM4nEQwNf1wjvEoCliYL/aaVpAYx3iQ1Z+WQZ5lTCkOljoHuMX2AYP0McWfqJ1OecInaXC3ow
yzoZA7fnlvAqYDcQ7vR22IYh7UDNRq30fO5OeuMlqVHIo8jz1A43M23PKdGSYbeOJmNw4EYeNPfe
nVWqDIQACeR0wr9jhM3D4o0ety+W9o45hXTQLHisKVB7Y2LMy0mFpSfqqoQSr29qILrQ/50we24S
MGnQo8iEAoxXP2RXcqssXGHyxkFocAh3Ja5+xSIYSzowbir+81mFBhuVEhiodICc3+IOUgFkw7k8
wrjAnzSLWDYJPVnEuzoJi6WZ7P1vA8vx4Qqwnk9v8x/s8IS0z3/YErOEuANMqjKcr166WbvH/Juf
mpeUi9DCU3mSrmOUWBD+lc/ba013ZQU8eXH9MU0MNpDnzfziLUNAKCKGmNaXd4HrDH07FVeVKDqi
cYDyQ6Oy6o1Ol7gO/7orHiZnw+HO5SxcnMl2tJkNTk2uEPfDA1AppIB2hs3ueIssKFhgQtUHMR4i
aNJpvaozXYY8NKI9ldj/dpnCEXy0PeyVKUocJeNGcxHvfATx3fDDcoAJDRYUGVU3MiZgjSVaby6X
uva3+DjDQrtyheptBx6ryli/Iztzir/ZHwTKJ056Ao6XxYy8yALu+0sspae/BDwmRQ2qpgt5Fwwu
VKocpcuTyriVy1xl7STTTZll+mMmWTVwoHOlPofTJe823UV/pCLDTwefGI5XDNIeK1IGbdYr5Cr1
yVmCSiRHejh5MdhLd9UGOgd4VVNm8xWfsHz45NsW4dP7LOjSmrLPzz8Xa2n3kWvPmdI9a4QTOgx4
Nexs78aJG4WFIF8e8U3MBL1g3PpxRzXESo4wDhZRZwZo5Od+mIWqGwSvNlf9ZAIDASAbiIli2+wS
PAutQMQjTBmbEZSz2mKvwe2p9EX5j+8xcPwcGw0UUm+7B2TvOnDeihcWfYeCGjmUqIXhoXiYYyps
VLm7GqmLkFB6kfUEvmTm2Gv+vd8mtH4AeqOq9qQjGBU1meuOtBPIaekktSLDMP/ARcuvIT7KAKDK
klTY5gBMrWjnArSmJErB5SsofA3spS6RhncSAtkYU4OXPWHGw6LVdlmadLHNe0bZ+zcCu9/deu7M
azzojN4vJJg7Hri0ntsr7ddCwFz5i6pyYk5nvyM5z6kVgMdJiov0vliJGD9AT7zkHEhSkwC/4oy4
XQE0wZtNiVLQzC//MueTzDQVT9OFGLqQ/XzAU/hlVDRMFWYzVhkLgP3JIM35DGWNha1nE8QQyGYh
Duqr2XP33J4ZfnclbeHKN3Ps0uLC6gXDY3cYVtG/iMCJjvLjJjEmDYjjXTPH/OEzfA5bf1v7P1+u
wywlv2jc6Vc9+w++56gBylDOVILBfeuzDRd+CQ/I8PyXdngHztYKJovt2ze6qCkWVrGex/DYKcTb
NaqNoIDgc+Uq+so5PVzhFc9au8jpfq8eWG3eBpgWD0pioYtyLMGjpWFl91iLGswmWNCzrojSsfzY
W3MRbaijg0kkHPdRO5BOsFtIYEjUruRlDY7iL7LP6b4GhVEDCTkV+grLNJGjAgUQRUgrpYFeD+Op
mi4o8YVZL2rzJrEjZAkOGg3hNmnGtPedzMouzLbIX54fpDTgnRCXvtVJjLHY39oZNwJjxSaRQddO
YRsv6mrKtSV/kB33PA3HkUMkgT7AvIedJkQxpBdqj6hwAIB1/xiK7M58M0/S10QIGVVrFSDYJRD2
ecWk/9YZGRGrLjChQlIYtB/sVTyUmM0RRV1eD5ASOaxOnUnVCDQ6eXoPpjGbYKiAUTn3DRou1TRq
01sGH4vdhgrJ9TsLTpqpxt72LNBNBp7nt4d3uOhkEeYiVzxHZVBvgEfFQCnMONytR0G9jVDTstnF
AFGBhv3bOo9RSICBNYqWnQcpF+BIIPcxr8JlO0oQhLk6JayKBMJwGZK/NhsPmvjmjqSfmJ4VxD/e
ZLuwK86FUvR+oXgy5uiNFsUc50cq1hzZXeA5Lr9/lkbpyXk6NnrBKIVU862jRRns+ytc647YuRzE
s8gY5oJa6fzdijn+zCo7/u130f3fbq76P0vOTnRrsR3oX7n+j9KvfMym5yVJnJS+c3j9gmUZwzPI
C2BXmGTD8QOIE1Sv6HejjG+9Q+rqDCPV/goeGqOjal5z8gZwCXqABEPPOwW+6M4x21eiIG7K6CIb
QERhhyDmpK0eWdQHFslJ1K9Rywh8am3jnupHMwXCxwZUhuIvrt9PQMopcUEQrodRoS2VsK/iJcMn
LtM1Nb8bgQG2IxJXS+78I5ZB70S0b1q8xdhKTfbqCFqKrh17OYh34f2krUyMl4SxPYRKLuYFhthY
k7WqSi+0lgeOvaGnUMA9VDjQClgACQUoiiFUG3XMvDx43n+LiFFhW8EcReIQxoBDYnzy1FcAUPPf
kCuOO53oPUPeo2mL9S/jaVmMc9Vpho1/6JLSryF13EiJdySfqfdN3220HRs3IQvCqBlgJpz4+WpQ
qJNRXwIuQq85xgM+8pKUSOdq2ct9CJ2mGg1izgiuzVVVg1p5QclJihcrlpIJtroFh/1OXNTlK55Z
uQjVb5cWhFOunzpZN3qqFjCriZcqF4FzsAFttmdeZpXcRThCTDFscudkudxUVPsDzmyAO0phmoSC
E6+MUAdxQSfKZon2MoR+FeAZVjJQ/xgKPqcQcQUr6J7Gg9+f+au5VJ0Euqs8ewN5vW699iom1Zxu
S0+wW1i44HWBCFapTv1nrkzVwxKkU6WvBiwYaj8tp33ke29LH06JXl7dZ0iB3tA6KgsGgw5dkTpK
bDsBcVBpUE4bZyO+5YD+gr3KXhMC08wKX7AowAk+si1ZUwJ1f1WkfmvS5bMF8BMY5jewDi9qCfN6
XMuX1D31Gm+GtCRa+bai39vRcekOLB/Uuv6Gk0hVIuh2xCtHk+mwzLynn4TNZFKL8hSwS/ULsEeq
zTDsq9SHNqAwSpgGDVo9jEiw2dFzBfORNdz+ExNGML/PU7OeWProG07K+zlBwe3nqfUUOpwR8Ldb
KquUBYg7bH5Nr7R3/UELb7TWSl4qB9k5cLuTsmEoUOA4Jf6dCNV3bdyUMvRm37MuVqDXLbNdpwzb
hQfm6rKUhNgNwZdrdOPBeY7j+YoZAajthvvYCBniSJqSPhSiDCY8l7gXxyRvnzZ3oRMJPlu/nYq+
Moxwf+VULd5RfABF6QZgaDsSC3b13ORfMI1n+rbYHs47grSMvBJ5pCvPl3Gj+t09n3G4s03Cdctd
CYM+eT+/9g6B8cSAsamV83lgX4vTqU9eUy3WVb369JcXrMJqzuvCnVlOXut9clB+Sx6CV+uf8kis
7h0s/Vr6s3ht9JGobPVDxmJ2wLN/cmafa60QU9sk1WPs8XeaNDiQ7QAaJcbSkW+Nh26tX0QD8rkh
FQ+yezNyupfqyqow3RFH0PlNA55RhJkr1zlzXEPTHFk0u+Vzcbq5eg78lSak+IsRECRzpCTXDC8g
0LrKeqLoFzWdN1hN6dZ2F1fwI+rqARRsuQMZPbaJiuB3ULxJfXDcRBfo15fKO/YggwJs1NzUF5Si
xWVZBHHV/iJBfwUq32DUsj1ilpReoIXAfGFGvTwgwn2L0HJa4sqMUz1wXAya9/fALUnoPdL7J8ya
iiFZYhY17vvFnV/SNRjce3WdA9tMu8/3xv2VPhTG6Bd18GVQ6sd1Pu3Cl65xY3L725lW0W134/Sa
VGPtBdLURekbsD0MJttSKlbrfTgKzGImiye5906w+i312SZog6ud3iqWhV6zf78umbkDBKUY8q2Z
kbJGpd+W3TNz+JmIL0I7v+0TIckAJneHrlh1dyMl4LS8ld92uOrrHQPKLCN8E+GsyDdoTvNyWjbr
qHpr9WUef+W8jepidLL6a3uepESaWkzHNF1zGCvqyEN5hGrXPpT8QvndwD7Pcc48zymPCVzzspnb
Xh5kFWZnoYiDl7079pUvDe+ByYtIjM4ZzJPNpwub59DZzzgQjWnYczoZDy4NO7Olj0j+gnc0hMll
6EWb+/J0kCaMW9CfYdbeS0aepRN6JZY1PSezoCsAGorholQrNoTQ1zOmWeNCHHVboKZzDldJ1dCY
Sdn7AoGJH1UA3xJ5wJBQ+wEhcrMcKMOmmPuiwFD6QN08/5FuQB7d2JCwfoidbE7eaoJ40ekbqRqK
bJuOFYjjnGxq9x2QOzDNyyxtcZhyzFIzBsWMq61QkqAYn+N0gTj6yA+G3TSpaGFsPpcScp8F050h
hdWj9yN92W4unRrDZiAgYDu8aLs9dQIUJMz03U/3/kphMO5qWZefj06Qd9Lu7eX7EJTTf4/QliN7
I9n+dbPjB0tEm6ifi80vPTrkVLeuCk9FARZ7A23pG8RWgBrl9EVImMuGXKAvoSj6ZjqnqeBq2bf8
cPWFpIHBCt1OUZ/sSOp7U4u7IsqA4nNg64a2hGjakkZURcKOZAjSQ7C0j32j4KWpeOrwqU1rdAQA
fEuV6HY+bDxUvOY6/PBWKgxFADvJifORuewtmBjEVhDi81lEDhYaCZ7/EQrAWDcxBK5NpXrAb/tx
9riUB45qMnCD90P/+ZOXLbZhF5oyl3tcHMvrvWultO1SNqXoPEVycl6jdHNTs4Ukmg6VqN/vhOza
9KY2SY/oHjhg5rFPC33vuXUJur0ldghmB9f9hcAsaKFZeZUZXWNI+sA6Sj+4/GvSSdYyK4IfyVTX
GfQX/8uK1+S4VvTOWKG63bnIGvYr9RrBOqfdQmRBQINr7gS1+hYM08YurUJf0vJtXCACOH6IyZsb
5s91Erg09OiR2x5luWTmPWVpe/uilykJWhtAU37er9h6+W1WJ61YyX34F74Yii5zHyvT6Vo3C+co
bjxokI8O5pNsjIDP5LNVPepeIpoeDAabNDI/eH6t+2qsF+dW2MJ34JNky/Bh/GGufMqwFav+sgsj
YBFT6uvqNNOf6Z6+XroRmLqBbeAZ4jbt0zDeUJA/+f3ODx7X4d/RCNlTKAyw/A9hxldmU0icq/B+
fwNG9/bB38A/NLxv0Yp34h1YEce2w1y+qAu9Xw+UH2Zr2dN3nRL1bpUnnMEo+h4XZOyEJrBenEb9
2rVdLdS9u9fQ85FAL3mCY5vcdXimXEt2hXUqaz5GoohTLeQMUQfaGWc8UrhC9eLoxDA83hQl8HGY
CjMaeEm2TORMS8m7I6LeNes2SABk3Yv+NQ3BYMwr4vXIIpF0djYVTZVtTYakXFIejU8OPKwl/NHe
ddGUr18EUR36/D14rLJ68AStYYMlpIwrlwTf3ldsOlaevxFN+2qzCYTJd09GuQGH9DA7cYnUAFvm
CnfTMkBwulx9bVPJb6WOKPNGxhG2Jw18ZQfDeaJQUiCu8QFuuHC/qTw9wbytCHRvuIt4Zx7YRy4G
fO3RRLdMklleT8rZJGxE5h1esgZmyW+iNw9FEdN65DwJ75L45FGsCtNPEvXPfbBymURzafDJB6w5
Rcwg0wJSHd4e9rZLD0IA5bi2CEhrR9lpX6SM2zN9Nzc7cDY3oo/AQe0WMmRHi5Fdrnx8blfrnWl+
gGFjiRkb7NyD01sEPRf/6nWXSGkH5UJy3zv4hLqBocWoA1AIy/8yhYiTj6/oaz21NzsVvaI76HId
WMQI50emRxQhiq/BT13jKJlUb4xwVCJpYLS4qCOATmG58IhzbG4OhNX/VrLsS5vi114v/AV6JJOk
qJBSB5GMoRHK51z4e4OPVghCOmAHO9MRCXtVzrAwxI09Ckj1F/WgQCF9KZIEJWPJzwZGBpsoEQ+Q
K+Ay1pQKs4vwl3+KLB2IkPFwdlKs1cjzDcRIVj6gngQjX/XrP7D3UyXBr5OKTYVG8cNJh5ttPZ78
83lYjckzKuj9bxCgpVRc5V4SLDGCIRR7MvPdY5bKt1Npfu/B8D7lchl/XptMixCUUNcOxveXeyef
nJ8056OsQAD0JKysvK1K2Tvd0bDNxtd7i2UUrNHJ7YjfV6BV01CWY0K9fSEEaEgdqWH1oPwQz31w
Vd4yUhrklVGUSQ83Bgt2H3ZEtzvl8XXG17L1pMz4bp1x6BvwyAni+VoW/MBLDkey0zSr3rC3V3Na
MdT26EME5cor2wmHCezU4pZ+CkWnGIrftJwIzZXLeLv2FkNxH+1O3CTpzA0rOY+UxmpexIThn5rj
85LeFzwB2PYmvUlFgx2Fc92365L3UZG9YRJP+ql+OMnBWEmBji+CKBifeZG50xDDlDT+UDNAwnzO
r9Dk99aJEHsQDPRqNODxwTggr4QtENQVPy0pzvsSTxXLlYRPyUFHGSxlYTCEWtC1TPDX5sJa0CN6
/I4J23/s4H3C5mFDRLrwfSQfD1FB90HiVsQvj7g2DFulJ/Z8OAnTMYOPxrRIbDsM8uTOGA6r2iZg
UV/GmUXazOdLntAKjPqwyPz25poLa+Y4oT1LrbJVmPd6PvW686JIQbPziwIn2wLtK3NIfA5grnyf
bLuwmpSztLmcbLdq7XVcSmMuWROv2Hi1dNd3Cl3Js59wX0/2qj2j4oyEKgptQD7bo1LhigrK+D/H
YFe0OSx3teeD/fltZjRzMFk+bN6nr0JThS7yzGiJB/zZ9iI84C697iwsiO461UA+6aBdYEVV+j7I
ZND/IMwepzBjeq2WHJo4kMM6D5QIy1vecDdhgX2YNuMwnwN+ZCyksygq9M9hBSUaqyF7C9wHb65U
824HbuIdHEcVo5MzekIZqEJIkuC8J/dOlM85mVoy6Lvx+FK0i0tT69kDiTJeoyYcD1r+IcqTVeVx
zoPQzJfnTQEpBKbqGSnXPrDbxqPs32qDfiN30kSXvmk+BXVr7NpfyxSpWG7q+s16LhzPjN/ukb0o
v/RT4yzcM25XWyI6WsCxdyyp7qQLl3m1RFwLFyWklJ0TfRCMX0gsibiNpOhPzukn/cy6rbSX3PjG
BiqeUW4BBwiavqAyN2xYg5tXkdHKfS4mYPneTBuxmcj69ZVoaS1f7FBzJOLyrybAWi8tNF9gSPWg
sf7oWS4rrkKmyiAh+daIzcnJDCTge9aLAce5z95t10dYvNqBtg4cumE4Bs/rNZd62AsLSN8+RSMb
XcA+RaCre7pN8X3B+GZhKh9ZNV5znNT7tBEVemyJtr4AM5HVHSgIybVCYnlC1xa4+l8s0VQ3eRLj
F+qvAnt14eMDGaPG1RocxCsVxKaC5tJBreN1b+JPhP1/1/1ajiNL2HB3BWJOzL+OKJXq/VsHebq0
CyV3WmAfCSgirEORY5tRajhvwbfZNt3jHq/xhDij6ZxYisgWc/g0L/lsJIjoxLysro/Uc4WRY9mY
J0TpQo6Hvv8LU+B4YTPaerFXJf4V0cBQXuthZ4IKG+grzeza3mMBBxJQVFQSMwXf2Tm3JtXjOhT3
ksfDmiqof6N5O0Sm/YbbsslQKtKLgZppgQVLHAde48qVC4o3OQvqETzPhXWA07cpN1E9uq/+a9My
iX+HbeFrmgn1bUx+L/g3dryFUVEraQHQg8NwXFn58NcbUshcrmTESlwqKcBKNmdG009u8/qSG1BQ
HCN64K67Q9Phf1MRxOJjSLfC55BPzBOpmO0up7KkMD4MwNva5S/xHKtY1ZIynYLN/ReoDDhB7nv2
JnHpzBaLVIXuUlVKN7myQuFqYrmlTdNxBQycZHSK7H1mCcihYSDK5l2GV5PiGvtp0qlEnFLGNqc4
UcLWV6N1VR4ELLM0ruvjUKhPzupy/VhRRyNY+yjaS4bNb6ZPfXa5XCRc3kPkNdL5T62xi2Z5meli
fPot8YMzzl9HVLvKS2WePW+le6zXYeg77CLdKjAptFCrAo82BvTwhz2eqtKwZ+6RQKv3LZxggGTg
koW2zWgnalNwu4Dl3vrVJPdv84BInVgPvBf3bKnm9xzde0IsJyJu6J8LVcuOlClffE7VXbFYS1tU
kXtYGHnmpkpWPOmVxPQWFrwO6MImvvSyL+jWJaFhzEFsmOUsdk2KqtT3zm6TikvJuWU6nhQ+DNwn
FSgrxA12mKujz6N6zC4ZHuW76HqykJ/lNbdx+9QpxMexmC9xr28/kWM/I/f+AyD7YV6Cdh8T8MHU
7gYjQ/pK5pK/+8t/wlXKVkue120Dkn7pcWhiiFOaxM0kPZnv3VJ6grLrSkkkghC0R0x98WtCTgO2
flyIn3cZS3Yu4JqLuJFDalex5E4rIE/Sy5nGoLyU9/T1WFx6Xk+whcFRrWc6+WmzIwrhuDuFgWDF
Izaib7EUSdzy8GXYdRaCl/Pz1FaOjQTdWtYAt2myEXvWY6gy8yVmB4AETrRaSg25AMHrSyv+gICq
NeVsxP7h1s4AgOXBxYDleLHvFrfvIAh4n3v5/sM3Ou2yb7rGAFsguErvvmqhUBhQp+4RSX6akWmx
/9hCpXq0npG11NoyIFI7F91Mffv/poeUXoeyMqfM+aT+Re3G/D3cHWX5OjdWXIfgOwiKRT6Lj9O5
cfqDxSnAmNRMAxYIpjW/YrTDWsyC5UX2V/t1/fdKZIEBZiPl8PQqvZgW2FBzL7YwTx/BuoKs5t0L
hJdLUOAT4mOg3LooUQSEH9Yassfhd9DK8dWrAWBtSgGjzUq2gDGQUy2hgXitVHkxrL8egvsdRsvL
c+9WQSd2Pgr075d6obRlRib5j4iWEnfTI2GkVhJl+YsSb/CjKzphLF8ocA76/JrJn0etD18XndbS
9W3J46nSDH7yZ+vnFDhC/iObkvl1fJYTtnwvGnqVHyQTCMMXMMY8V0QuaqUZeawN7ODqubGq0rMH
a94XnHchEUxmKWn88V/PbknNOPp98xDQb4CclJKPVJx+CWABOCNE/zJ4xfSNLoAzxmHAqpp6AfNs
ee3EjbNDyj4EaKrUUsw2twcv2wCoLConplX0FcN0Ud6yvorYa67/ZghWQnhzqp0di6hkH2x2qzve
3avyJNCDYg7MzJtT+n84//fGy4bUtNElL1PBVvCpiQSctyMSE8gZkI6+wM0xJua5YtxZ5UuYbHI6
oY0JrhyUgzwafzdB5sDz28njaDoHI0YmPUnDnMF4WJS4J3zeqhiRGI37Vv6GYQDBHE4+e4cn64d0
KAnmeb64Y3nmWDP+0KgaKmbNIkz7qk/ia/GC7QoTl+sIJ2EWd9slkgLoWDIbIAEkQFS4OhmVH6Y+
5OeuEomq3XrBaewLFupdbDuW5/eyIwN9oxziyyxHT3Zvyw6Myw7Fqx4Urrk8G2zzpy1Q1ItYFpOI
HBhcWgRPEXchIAMFgQOsPYCgHBcgxSiurXLWwqU3HdX8a6YzLXuiqGG+iWh407XgD1/HZ5vQB4YW
miFUBWmB0m4kbTVUiXHARZN/M5JogeY3mPf8mLcg6QPD8vvuVGPhz2Tg337BS+d3OPaeqDYhnOOo
wFVhc+fc8N/WqG4A3B+LL/nxZ9To3aAuQP7MAoSis7lavNRM/AyU2s6P6F3e7mO3OmTIuD5gA9to
769AgERMzJM2cyqiS5SuVf8a1FauyMFJxh6rQlPaopV/iLAK41IMGtoRIJQpv4uaKCwi9M/qLeLO
/uZoFfL3roH+aKY+gcer0MEiTpzTvIF5mIAKpUX362J7Os5gwGMVTYd4+eWR2kJvrSMuF+6U7gtM
p4liQdOjl5hrXBjl5h53OmuXapriZBspEpLWlC7XVJzlvlboIbWHVVZkpquvfJdKAI9vpr/0ZvGQ
pskkDQSFYTiDxoYZMoA8tw/pBHntoyn81kcX/v2k+5FZlCQTBX6+1z7VfMvpmSeH6NpR2HOapy8i
tV1hSmSoCjBdSf0eithre9avJ/KG09HzH6mLe7t2/hRlJ3XoUOacQqszPH8aiEuOKLMIqCqFwMNw
e938NbctCTjRNZwxl6lH1jLuJeyokbcEwsn4Vo123rcPdOQfsStJ+S1AqRoHCWS+wfZ5AoJBRWEc
PVrKoeCzxGwJDkFf/woZ7cE9d+ZK4K79yS8/6KJAg+GvaoI+A/XRbfrXXCLuEAOq+FSiX04HkIbH
2EqRkJmmDteiP/js0uzu/bg73XHPSHKk8RVAfXUnyHe6CaEaZsw5gBT3c5ILtjWCxciX4bYaV3nD
tBS8M+rUR6aNwH5nRoQEjpAhbGcgA/p/JzL/hxDzW6CmLTLS1EWORdzx+zoec0j7M6/Ez7/oPL3k
Eaw3jqEWGUiTdqgkTPEQYrjCTcSHjJRUkL0RnAlq3AyvbdO8hIbDwzh6I9tJ+rodTKjE6i2VQAgw
Xyhp96SQBjFnXIhH0XgyQ/8ISjAetGfHTAId/F4oRfn+MuYz1FkxWotjCj+UUTv8L0PInM/euzvT
GXzyOGLwiEFT2Uh1LZz7/oe58M64R+3aObs+5rVoagvTHFaJuR78HBapfX4fGpYlNOfhEslyd5OX
psAQfvUFg3WrP8eIV24tqXMFpSkMhuo4fkePJDegs7eRqXCyVkisNeZAnJDkfYJzgfAvP8OUa8ON
6bnILkKJzsGmL2P8d8Z/rR+xVSKL/Wpn3bjxX4/j/D+Z76YNe370ZUGAycYLRjIDVR+4bZ0rXA8J
XBelhD51GNt5apBDAXimkUlyRrCF1cD3YxBdGGpfSGJDI+dC1ACq7prBbcsjPpTVUYKYlTQLqo7d
h9LkrWpzaSSRLLVqOLsPjWNe1wf1i5npotZUIEr64knvOrJJb6CDFq36urVyix1nKSL07wWw/HzZ
jRQiJQDf5nFf1RKS9VQ+ySbb/Ije2mjVXDsq8NoY3GshgNtJnv87Ui3sfTbVa6dvVSQ+t4iICbl0
2IEAMYdCkfdslzhXACYwjHXgS4DI6jakzszAlYka4mi2FuHy3Q4aE1O2KX1JCocHQGfMeiMdDI6u
LlAT+o0Hxh9MXQHMY0WOmIe690BI+zf465RQW1kuz2VfR6nnKC1QBsNiNGoyIrAZL+Lr1MklqAa8
e3K2V7Ol/1IkNGI7SxmZ246aLFtj8m8Tl3Qi7DGCz7Fx7Xv6oWOT+/teZw1FvTCQRpXOQO+9gpDA
5Ew1z6EklNhKdv5LQ3/OZes4K3D5B46x6xVxhg2JK4y+Q4ifrOABzlkVImkORFo6a72HBmebyJ92
h5oWT7Hq0xPjNyqam5AYA98ILbjR2eNZcClFEcLAHTjODxJW15FKVg8RYQXfHFrd/+L9ggjiFrP1
3YdE4pBmfSXo8XReSkf7J8aA6oNOII3KCAuE2CYm/a6r84xqbi+rw64T/X2PSRGFU7uNc9LqjjWf
oq0mII9adRSL7JlyBeMwv6tOM0Yz3BLJXaxpKcdVlgK4AUnah3uLoYVn9sJ0Kfc+KcaXXrHweaho
OfdWv16gcJsKS5xtGptH2n0L6c0tR2U2yDVgC15pQGydmQyd8NfxBcXBJG0SNz8tdAjJisOpq1uo
tQ2q5VEW9IutjwkcYm/0Eicqgz1ip9/OUwiwTgnwb87w5F/cvzB9Q/w5BIBZhSW47Nb/MTxwUhFz
PdpjoZzjGqjPdw6SoAYk5psEiwQM1cyrA0ZwzAuL6fiRHcgZM2W8yEWbT84ZCXlwR86NNfi7AEMs
LL58GkjaC1gkNDw86jF4glHY7MvbU7hfTgYfUYt4AQdS81GkpcpmJgl9wQubkITbP1xa3p7E6Yx+
AvJRnvD81WvZPo5pGBRXE5StkUjR+GvPDpo2EhnPR1ClygO9oDyZ0nVH1ptlrR08DcjI5gZW57C2
dcawoJkjAM5cvAYz65KNqWxGoycnUNYxYBXcRoSKDmF0uSs4yEvSGh8fbbzdG7RG+pOkHol/t4Rr
9gE6EWyw3thWFAAs4WgIlkZniFQuzkHX04Oc/J8R5Ue7osljrPYUZ2KNnXKPnsLj7faVWXZNl4nA
fZXSWX7EkmTjqYgHYrUxNmyp7jemPLBcf9cO/zOWQ1ZcA3jposnC/eqKycvjtJuSueht89uSY5OR
FD1i729gdzOaOT0aZnNiS00q6T2CZxYq+OczZWiZefuq25ssYdNHgoDTjYMc7k9EY2cb3IYyqrHX
33+mGLKP/c0ZISpUEMe9apmWkiW6L2HecR1vnArhv3nMWQ8tl9lasSrw4tO9j/ptHcyIVI0oY1BR
+0XtUemMBC7//ZYx3s4mMqACxRVXXGf4WVSN1LO/iVRYvJBBnVYvnwjfwpcSjXtTTh6HYg+wzTFO
6hRtVvKiKpk0c4U+WvOlPbH5F9xo9VgL3pcJp24rERtLbA8D/VqelVPNURO+0tMH71+sxpUWhuPr
SYKgXIC8ZJL3VkxXCoceCNoMo+xKog9fOGhhtaLNBxMqNk7pPc7UIR42rgUDFfgy7JPv2pigSEGj
T86ms0pFsmBmrPkUeglpDavwdFO7LKK8FnPdkhDtd/YH3RAMt4djbTWcz5JpM+dnlf5E+nXnGZp7
VlUkAKB526K/ZS3CoAExTn9qqPiN8J1fvf3SLihaBVj3SlqgQduNSseNWkdmuLMPnv5GN8YuHg+O
9HFc1rYwO6Co0x9dDdsj6r+rH9tUpM0ISl1MXeZjlvhZEdj0ubSeaizyO3TmJCqc/9I456HCtjB3
v56jFPKWsGD9wHsLUV6cCp45gQlR+Hj15tcKpcWgmHP2skoIyjusbXT8gY+5acbCFesKRyac/nUK
VpoP1CtYsUmHuLN0FD8zyxxigqFZC+lste7DIoG9jVBmqBb5xKJRbUi8vg8bw0E+OinLh4CUR/a9
t2EIqTAtv/NHJHfcEEcNP12gzVudcnwUN8B9crE6nqVeDuPOoWJJVt9sW67RI9rVgW3f/VS4YlG1
sAlhbiwxQdxliRqO0HziwV+IP31G8gMFL4JbXR4d652bzP18OO6cG4iZD1qyZBqrx+imMcx/lZeV
ObuTuEvwXjVngwHGU6Sy/1FOBw+DZ2LdOhLDjtbDTVyf703TTezzFalqUfyWeaNbBK/EBWDwbBTD
sh2fRfdA17aSGonsT4OiJLIgk587lZMu0bOUxmPrfaD5B3u6wg66Lir/fthsq/G1GBxCkBcR6kdE
a2JXfyvooAlp6lLp1CgXneH2rvI3trPVHTT6SntNkksee52OKSMt4EXrWOaWchocUDvibBKXSJD6
etRO+Vf1KxZDShe90lhjCR75whaucVSFMVXEOXy38tbQSHTDJajHrhq7YKSuJBV+GECscP7Bpnf+
aQFqJA8rVWQwaFFh7QmI0UV/doYxxeUL+KJJE2FeyxSTF3ruLUugixexxXFQFyG/iUM4ogbJNLjH
sq91gEwQwi3JhykMDNWRbP6Vaswtcvh/6BQhvqYKqTXddRavnwQNc+xUxoHwX6jnatARp067J0Mm
etgvCndnr9pBsY8SKFUZKE+XYJ5F5gp8Uz/+4bKMzf/I0iJh4Jga49iMZoC+GFcmEEPHmlqR6ZlZ
kWsuH7wOdx3peXIrU+eJpVhRHOf0O1IxUT319WIz6kAvPeEZ6qKVhaoktQaz6FHdBd1G9MfGSs2X
PzkKay1/3OV6B8UN8MlNrm6MzVt654DRzeM+BykcvHuDwaSpHp6EBD4UnMqobD9NnHddltGYPrIF
RJ2+F0uyOMr6HYGLCK06YUp4h/jcaWADs50YJWpjqvtpy33FnjkP9AJxdMhaAw1EoyjAwRPasDj5
RXHC1WL4B8tW5r8fzhO6hcglupJdD59sVmLDONy3lvOuzboVt7CJbbmUYe6pn0J/KGWZ79WlA64F
ILn+/QD9oBLqCO88UtxtB0BVHxNiTuCcRdlnV8mTbs8txD9N4GbuvWUZf2UrAa+AfAK0+YITM9zF
O136wBm0e4EgryD44xpSDR+/rkVHvzDaFMhI9CrkmPyGGUX1wbJ8n+vY65ZFlU8vGvOXtuHRFsw0
5pDuN6EUaUlQHSnMCpL/B/WiC5IjNBV1JpNwVjWlgczYrZZpLF2+1FUSIl1dDUGZI9Zf3Sa7PksH
IO0gq736ztOXfCCVNTTuogj+P1mewHOOSbuno+/fvGhwe7AjZvljPc/gcTvR54+9/XmNreLoiLEd
rTQECu3IA1+jRexbjnxVLVIGkLBRB7sFVMn7dZ1WnGNifzNs0oWKSEl5czR7DFR/gslqVKxvt2vv
rhfcnWfBXmk3hZ03UNu7kvJXQFUEXZ5d60hnpW1xS8s4tlHT1BtnXk0Jihn87AvgN+RmSOQtjoUX
pSA6GGIL2GUepO8HAReOOglYB6fkvCoZUMhchCwiT2ly2r0TS44mjYT1aoly1KqU2PtDsLojzPZV
9Lxpc8pVUA0gKlzBrEi8ZgMjDJcse824XefBit3BIovH0VcPRpiTQRTt34IivwLSruvrhwPq/IeV
mCDCaKKTwFRLk1PzQc6a9e/5M6Ia8sj082nWfYy8w4qQ9NexMkgeWpYoHU0iDKY0mXOgAYLJ8IED
jVcwkzWwmSn8xzAQEPoXgZ5Z+SgPnqsywIwVdo6KHU+jISYQiFA0HsYHNVvvhp9T39OR8g6fznAV
yoo3mf6yTJsuW0XTnSViqVqkzXQn8HCMV0zCmA6UNEYT9CufdEC2cKUbTKdePU2vTpzd5sXMZipy
HO6GP7u4ecXIRYEIyprMRfu5WsBNicqxIg+xIEO1qfIDflYF7iqf6QJlALdWMUvT87H6o9L68Jot
NhSMU8Osagn53lvkJQZKuNA3tJrJsrfstz3L5nKHVDQa4LlNVusNHlpnGF7n6u8JFtQ8kewhxUEx
pzz/hf0kYld6ZIggGCcBcVreLf1aL0PzOAphOuEo1VhnLKhAP0SrrvFV/qBps6pyVAmwHFOoocOF
kv30TF2cGv2lNTZzf9/oDxmGcdGLSoYhpAOp98S6TDjvrL8yIxHrpCR9RGFtdHDG+vAWRriru9AS
bUmHx22yW3ogF+m7Vv6/ElnaXQ04IVMXvD5pp1tnOPK96kb+9stmO7NUwTWVPEsdvkKJCWxQSBtO
wIGSgbUH34ur+VKeHEzX6vv0vNde77/goH6MGfo12cHfNHyj2LHyAf2EmtmrCnCu9xdh7WG3HvG6
buynKWavYHPSBG/vdi+8EZtqmjTGPq47xtZXKGkbBmeII0odF6pUPF50vBSzMm423B32fyCWs1kt
c3UPesrG0TM1DjAYaGrsZW+WmXCn60YuvnwcJYz8A/gqldZzuX5suZKVCH/iqHGR3XzkmcebvFpw
nZE97Bd2kwYFCXZ2wcouQXAR0nc6FGebim8QtXDRQLQoIsIOYMdgosToeH4lb4vHTqv+UJVK9ILW
n71PKk2ynx2Kh5atn6DOZjoDJXSRKxlV9HC8HuQfAYkLoV0taMOE1YXMFubCbnkIKb/nMV9CXRiR
HAr6A+y2DD0VG5549W/je3VpEsKTwG6zRldbsIi0sWPrIpCszfnU+hzJFnQa8AIfM/vGmZr0ktMz
rCJ8MdElgEa90LKQ6/Bxj6vpDd+Lj1fld8wHMp7t01Wy68mRYBfxummswz6Y6iwfvbto3S5zIWtC
RqoPCgvIEufD3QnE1VIR75bKWBqzw8ehgmtemT1CfZSkiLJ7QwcGYJp7fcHHeWZYmSwvkTlxnFa0
3joNRNwdhPz9F2AFKLZVu2aXzNHG5WqDUswy0qsIENXT/UIf9RYUyojlc77zFlNm7cyiDoR75XLX
r25jdL/HQXlt6eK3yFBZrjgJJWFapkYWYontd1WVfqDC1oWYc96D9ioJtTUCvK9KV75pIFEsDXGs
ALuonCEa/HNIslq8A/GbXO5M8oA+luue92kFFdNvhziw9QnNt5lMOtCAWJ2kX8FZMLkcxgwK4nV/
WwBUXlNJFkhcCUJO8V8fD6Jp6gQhZVLztwsmWuvliYeANg4sOIhD3HVV4CsG7bjg1O3HqtR1zV8/
+j6+4RYWBpJE5m7h2xvuSz9Q3caNKMVHDLA8f2QHgr2OrOGQT7ywxD5Rctg73XckPtglCTK1OHlU
5tgYTYHcxcY3bvvKbogUfTVPPC7yEZi4bZaM7GLnEQjXBdOa+o3GmZEjgfW6kIZeh8Dc6n4iQtFz
BwxINzr6AjbE2yCkqMPWvRuXe/IpVB1W1R+9xsvHC42y+jco8WNZihwcIbqnneAD8LuO1zoTbqYf
ZWgIWHhf10Eb/cvi8MZzyYh5BmJUnEchGf4sd6XpefglCkmUDpDyTFB0857MwNd8fxRaAlzpseNT
dWCpAnhUFCpEknNah68qTyEzWqVDRi88NDXLE3oGII/nz8g6Lcoaw98qJef68IJdE8kvbFh1yrXs
SgiF77mPAmrzZVdjpe4Lpcz+FjbudjbPS8gn1vszpIlJgkDMZqIQw2sA2Lzjspwy+/PVdzMhzp6l
T99MHiyPy/+g25mXh17Vg18olsnBdJ2RlDxHX5j2dmosIPLqnKSC4F/1lRZoUOJr8FSUbJ4T6lqJ
rpQL917IGVGgz3dNFXKane6+/akAFpHht3sE7mNUVZKjrDJsT+gDJ0/IoCJ54UhOdzpCf0DKjU1z
6ok+1BTiNIP+2RTDcBqRYfA/Oey7yR9s4N4mSyPaIgLKQTV08fN2DxzKfX2Y2O6wQN/IqkZPVx1d
914FuxX97BNkinjwfv9lcBs6R6tVn2FfYg1/7f1W5u4xfkx6fmYpvbPy5dur0nuHlP3KBcS4A96+
FJDo8l27xV+RytQKrTTAWmNm0RLjHFs2d4B+cLaxDLBaihLR34LD5gcivps9npDg0yV1If0mJE1n
1aQAsCCzEDkokUUSbGRFG4tgY6m1MjJs4OA6ZY84T0Zd9t7xQOoK2WTfNwgLwLjRxgWS6fw2+jwN
LhPkKM/C+kCtzK964U/wurkSGZenKWMqzHIQUJV3xRhZHXVMySwqFY8kjpfqF0VWvCJ0m+O3Aa2f
kHaarfcrl91eww9TjuekFHqEQB1Z2Jp6sRKcFvGwIxda6a/Ujc7bj2e25WaDY64mIBgSXzs1wZD3
+fOSV77/tQ8YixJHNrf1jIrfr327n/kHPhT7G9d53yZ8X3i/xBYZ9VdRue1+e5Q5V6eCh/3CIbn3
ix7ddN34Ar/w0snQv75Aec8sFvlrh86vVU0WsivoHri/BPit3hQmuGixbPR2IavYU+WsSFRkJ37p
7sm8DrQhzFA4ilGx0z6vn0DsUPPFE5L6S4AfE+vBbLVq3nNktmE+7+DtFhNRQ2yq58t0vgw1VEos
XIN3WUYfPgK36CToyMgUhIINzYjDj/8XFr9rsY4VuZi1mtIT0FssPHq9JmLo3JjHW6PvdP36uoZb
yBt9nHAAeTYGPzhITkblSU8bhstTDhZRKhF144A3gWaVJNKTfj2n2FdJUGWb5Ou0Klsozta1UpII
32UokNjo+cGHRQlJ9tpR3GFfFnsANk5ayQFZaRqEvHRoFNNHXva9b2cZOi5Lx6MOvOT298V5WEXu
maeWWZUk217UcfI17+bSokuJXk6jTns5nndah56Maolt0jHptbUBoegIFxO81uz3TEuLBicGEJ+L
HVw9H3opS8CLThWk9GKzItOQIANLSGKB5gEvkbSA8LnL7Ye82uxzqYBUz389XUHqoYG3XsUrdMLH
w3nO9iQxA0L3Q74vz93jmiAPq6ge8Yy94P3rAMAUphwhPSfAUQusrawe+ez1/FwMYSwL4ZZSafrS
AV9SEhJoAsRQmWnmF75F8/eL45E8LsM9IfkbPBfv4GoNn9Cef5iSqOskS8zNsJfcNGSZxrFLSOGs
9MMwy+IlSCbD+9oIbOdu7y8vQdMJe8Vg8KNteljnvMx1K2niDRIw32E52GdixGOOzpAHzB8fb/JA
9JzE7Oe6WP10IK4+/AmL1T2OfZsEvLfSg6eaEb1Xo9qFOZ9QnGzXf7BY55u28M8hJ8gl0bt2awO0
O8EBicbbHqE5MhLwzIAmkIIa0Lr/DuHxBW59Dhjw2OHfAu8AkXIlpBZiaAtC7E7RN+zvJZOkoCwY
MCCdE5HIrCi8aosq1sJ3PKr2xmWsE9pgdyc+KfJ3fFR3SFnnzOpvcoFOItLK6100m0GlV2c6P77p
2/PzaHlQot80M5NmM2+OkNz4mIr62yYxybNkkSz1BzcaXu+crWRc1lLkEkvY0WkDp7VBgiYqD2Iz
4j5ScaEZnj5lLUCsaS2e8kpeHfekCIrI22Ip7NKbrWIua1dXicP1XNfjRBIBnV4dNKqk+/RKewRg
QjhVWFTrQFrdc8Mu/CMxpCJephqRt1GhkL+MVwgTpzb4tmHT3Z7rfddm3kMkcq7o4xoTWW9DcXCo
Nj1Tz9QrMHHR+7qIBnfGr7kt0or3yv8HT0eL8lyMgdyZ/6BiH9ENr3fnGmS8fCLmeuJmR8VZLKFZ
YFupm1AQxMOM6BBFwP4axbuomSb8MhSYPmuSsOt00OUmRiq8eKXKqnyIv5dKGryNWKoYbbFPurgg
nq4lhE8Gyj5g2CzX6VOoD0tm5DnxdMp21S+EHIoWfeLL/UKPnn2RCnzL+7TRMgCAdVC/O+wKSnL/
wpIIzF4uyL849F31q5mDrxngrO98LS08C7FL0KBOw8PkNx7fP/ZcwrJpkbxKzZ0TZevClUeTX9ps
rmgwkBCdpCeM99ADdP6wvaVprk1rktVZf1q4dojvlrLi4PMxcC/0pJjZ90yk6qVScPivrCWRrfEl
IilMbm3noZQDBhBy3qoNhdyMB5r1oyKonT/Nhs1Uq9DVKLsAMJo2ERfG6Md7N/VCjbNmvhWdlwAF
7WSx1NY/ElPb4OQkupO2s/2bcXp5rfa7H+7Zn3xJNhHViaqIdEQDWFnFZOOvXScRpnOhOUeWOxSC
HFQ//PFl23HmAFlunDjXE8+ElUJQs1HyZl0bVHy/e0gZ481pM6tZcJHTrD1T2E6vjXkGu3DggXR5
587rvey4oOj7171a7mpVAt2IzC9WRbbx7hZ8NNeeoSjhJCc4e5a2RH2vYUV7fIplJZanfoCUqPeZ
XwxDfhUius2i+y/d2vVuRNfWMDnobA7cCTdpG1l2K346v9ElW7L3z6Lx0ZJBLhfZYkGbjLOZzuzI
Z5zQbiL96RBbcvWByTv49C8dm1wtMjIkoKkMP5NJPFJbGCuZGsrPncCOtDcJMuR9seqz/BAGn6gG
8kH3FaVSI/gJv+WURP0YBvTPjRjxOF8LS45q9pwT0mSixqZ/vKMGJqAorLKrprkHGlT6vPU+PNxA
Y282kK+5JhJ3aHLNrfUG+gu32KxJUzn+rHH+/SF5qUMGC+ypYygzwmkDLty5MmCY4F+8w9RSobN8
oES/lfMX0clP5D1ynGAXLUNbfqCMHgDWRdouUvXfEHsNkSVm4PNhW2dQzCpZP0oVCHBElWdZPnMB
kfDKO7h0JHLdYe2dY67ZoKXiokLISPYxbrkEutGE2f4KV1kDG7rI8Ab49w4ARZ455iGoYeRvPpr+
lzQ/YFc6z0hNBzlIPrMT0Bz8DEOLeZGoqn52o86ncCC/8NMkp/FZMuA187gqqQsgGttDIDWgXGS5
R2/UeKYMs8hTWpxgubWr9HjisuSiBx+OwPNBbk2jvxWl7RqkUNOdJ8Ukgc83cIeSuxZoHYru1pFF
xS5NjpzBizjWBHlo39XtbHBvs3Cokgy3pz1DszgB8W7yYZh5eLiNRZjneclemEwgr9FRs/A1Qet/
sKDyhJ4ZktXZJ5L1NIAKGOHlip57trLJhvDttNHoGT2+DMNNgJ8rjCubL4owQM22V33ZJyl7SWiH
ERqo7C7fXl1uJ+nA5wj9dTg0acgpQSQJ5sRKYF3uTXCRGhbL3fPvdr2gPeoZvJPebpNlUnBrRSqR
424kNNBdnlV62mzj3PTQPDCFFK1DGUVQFHkDEZfKlIzoqsscKEFMl0yuG/15jHdHQ5ae/FG6R9PH
GaCOkRChpf+MeMxJA52A3jsOdKpL/YhwT4JAlGwNEa9hAgTo3SAxWZ5au3FiZNrGnjICp5m1rrQ0
0RDAoZ9uhciqGqDCN7fXMJ7dinV+3h1D7tnWPrc6X46TvWxpjgCRAMqP53BZQv606eyPeJjofeu6
tWbb/1IZje4NvWFfojKIA/P/Fms6K3nd47jwYNgGnJnhGldxWEhEcRUk75P9Y2dql/Iyx29V7eFo
8xAx1uRhJwG+tLe1337HULFrpjmoL/S7ErQht8DNVL2mllrOzUKLSXQ6ORq6BTWMP5kZTm5suOe7
q0OYh0o1dHZIxJAZbZUcxGB+RI2RwhTc/TzBtqYFRipc+QWr4QG3o/BVnfwsrQWlAKW+shO6lpnE
7tmofU1u7r0uevMgoI1lJFXnYigXdZnqBxRV2Iut6E09iZxCssTk9qf2V/U411GKav/HpgCvnxrr
SX2U1eJOQGbwxHGcEMDmmhhGODejIUtrJ4T/bIzkGjtuzTfct27Ztm53m4FHrw4kNgJQntba0cHd
4nf3b+0lI589h0d7VpcfCw2LGIAY29QsO8+V73FqmfIjKF4kQB2g+sRNvl6L81+KnqEV0z+74M4Y
newxSAgayyZ5PLRxFXjUZIlZpbR8d+0id/bGPo7w+REXP9SNIs/NElmXTFVc4Qd2aZhYkeyfoBlg
aqZ7lC8V9XHnMFUInwOaWN52QbX9qgveqxHHzh5aG1HAzuu7UxKl5h9iiTqu6vyxC1+Hb+UO2FKu
oCg0Y0iGMx/iAaTbPHBzD76ySWdxUmziB/q7ph2EQlm/niG09fIn+T2oMYaXo5OaO9dZOUuVGspz
9cEeQ09k9ICZS5ucYM1wodJownUs0vbk3JVWi0xBgtAmIkgEQoSRX1iuMKlFM8i/++irkV/3n0XP
DzJVfy7bm32MhJPHN/9omKaekbow7Gq3xGVSEYvcUm7dxBZ+dcM0VB49O53pNJzOSDo8zwbpuVSy
k78OatEZ0CU/kAurkFlQWObDu0f88yoZN/ozNbX49zkmL2OhKvIBlvurb1Sqm6xOBufgQIPTL/XM
p4TFNY1Tw6skSHzcgZ1WXtLUF8OfGymHLcE5hdn8FXKsHT8OrXxHCOK/TwcQUR6qSIcOooodzRZn
iyqoorxj9roAT59LdTTyyrq/YhgcfogfmUoXWXRJ7MKDKngek2IetXOdruFk+ln+fBXjaC0dMDBa
1s8bJiTLfu0JDUuSU8wHmOAo1FkMxpgdlHSDoaZia86pDlvreJqgo+SCA2tYm8XP/jKsDdV88889
SBWuraEDZL/huIzL7gauwuihRexg1F0IvESFi+ZsMmQ320LrWttMNhQpfb4Yy2zwY5kM9/DVLMBz
ALlbz0ZW73GuRuUpXFNrAqe1oasv6htEMfVSachERk+KqCwpYxcgnx1NhydpK/TPRq/cgzFwu9W6
hiDv9BGWa4N7weQCIH2HZ8rQGWiQrmq/votyvpnDkIReUt3k6FTJOedKR7B3T/kEd46sNbCD5UZx
awOcmeDQ9jgARQQ83Cpce76cVabsp3LQPT5yuDBxJQ4ojw+dSDr3xWcxnQFIHxfAYs8f6BDTh42C
57UFF6Dcpy8za41dRgRw9VnEGwqYLZkKMuXGcbaTSgjF7NL0ES21cP3AyuBXyg16aZreSUxwGAEK
0wTTxQDY3XTQXSk0ZD7NxrkQM71kEBNp2YWffrEu9fXNl1nG2gR2K7Sm36vpPBBrHEVbiWXlUwvT
2rszES+0ainO1mvLDykiHd0vNEHso/GlK4Uy5eflD/sCkn2OKqbmDr4d+X07Mb5kXLBSlJYDO5qf
WCrogjzSOY+y2ZBMPRE71/EL4bLu5Gr43wpn/ko7zZ84/HlpDbguW+E0lBjfIATHi0OM7iamJgVG
hkyfK6wA3gMFvnAvqiPy5BO/sIqUrswG47wFDiuNdtcSuq20lU1bDLKrEgqgstxZ94wRguA5M9ha
DDep+E0HaaZoU37MEJ97rBlFzJ0zM/Z/jN+IcXCRBwt5QGS+70GdNpuC61hxxzimQLbuycR9kXbE
ll+SZ3XWzrUhtQzyAP16ixUuFk+Oy/LsI9YsxheovwSg4aiK+4fjrQ5UlU3xQ8YSNWQtJTKzigqr
mQv4W2NuECWA2V+RARZkzf80zAsooHjDksBdCGmqtl53dL/JcIY5kOTja+dHuJ09/m4zmG3qJJBX
Ibf1DC2FmR9SnQiR1nMnYHzVwDTCk3iTS4/BFo8b2fHNYk/4kN3LRLMK4dedRnknbTl3FgIAgmkR
loTUlHj2IzFuNigbrHG3y7aA42sVr0Xyo3J7VPVEzIVbSTy9RYLbrmqOpw7AjlBgkQ7eil1DJHpo
VHkEMWbYbohlSs7szmc6Comty4xXSMOiSXsDYvrsoRJhtgBLtKxa4+6yAKkwwGYJryZVI9xrKVeJ
tIA6sc36tQniA5yTxfa3/825xgypiV+qFT/F1vFwKsjTVxOrOJi+y2/sybiNQGwxWgg0aii3RXBb
kESrz19TAx7p4eXeAfvC9DlUcrGPIfAgIpgBdu7j2I0F3LoHqj0YNCdsWU+yfSqaVEiZtiIcBnLj
/2242LHt+ok27jex7iXaeS3DukNlUmkTOoigH96ynrc+nB60vEkRtjQxmom5+r1XEfeAvRRm6Bc0
ITaU0cWmMhsaCXsbJX4fp3NYRgXqjQ5BNFmv/e9NtenPvGd69CWKYgqetfdP4v8oHwrCoBuSEFWB
ssWzOzE3kPHj9rlG+YeNnG2zuEQYK8UL8RcSqonoVzE3w63NgcsgMnvH7BhYvG8fXMdFhn8Kihon
LuQRA17yHAyTSOyLRPQbVEjZTAxn/M+28H/YPzbHlxCyNIyB7vHX01sNTbECw6MhBhCveSAqs/IM
HiZNCklJY/w61XhMAcGf/x+P+QEddu6LWjSeJts9Ev5Qa0Mi2n+dX0WKPWaYKp4/o1WR32Z8BQbp
64uhEkDHacIwVJeMnTaw1XNQ2NBPaWbflbhC0yNnpKSIH3wWJwd2XVJS8jiqLQHtgreQAs18zndl
dYW+QelfCOy0Rc9Hi/DdIXVObN5+OabppAf1a9zgtiDL5kS59MjqszxN1SvVE+CFKKtFs1sBm2oR
dZJshdcHahptQ/I+dB1e4KsiwIdxWR2jBF4JjbtJRNsZw7+jQU1NGIclPsUe9UsutKDov2VCIp7R
740Euus0L1j2eyfnsTFNZpZNMehmLsSlFIecig9ZWrPTdLPZSV2PRw8l/mIzCnT9SPGWfblI+N2s
xsFOHVNCP8neKr2NyatFMHRb1Gx/2gIXKPeiByyjgdxvCqi30btum0ObHW+q7DuuhYPV0smMrbgd
CdSo86yxhkzEEJPEW4DG2QNeK38VMMiqagF2yDiK/Eiht6pjakZISknpoCXKL8U7kaOYrZ3zEhr9
1ExS49CPHOnQjkF48PSUv/G32+QQZY5JTOIjy9X9eX18I8RmehqZlXCnYyWGKttDQmmCIP+ZsDMI
vGvAD/A7/+Py0ZsCKe81iFO3dJug27vUpdvUO3StBzakIf1ZhE0x0J0tpaYshVLo3p6hl5L0KWZi
DWvFLK6CcKhqGUWnYJtLAlFgPDHA6HELvwy71JEarxYHC2cZ6r3RHKaQ9xPMz5atRar7Odnap78L
lFdFT1/nJhDUmSqCJfjIDXmH1XlqCpbIRbIBhtAXNoaWTL2u2NK3lRDbv/9ebqa5WNC52jDA60lt
aub1pJz5XZH7oskeS6hs5VvfyZwWGPxJEFphPfKAHqwHOu+sIHeTAkKI4tVxIQ6xzRuTxQHQkS4r
Jc7hiE0b/bz9ltFFm5l6H/TIly+VjJ35uC1VG+NC5bb2+AQX2cpF7FbAZz96I3Xyw2abhibfIGdX
aHlrbbaSWIXJ3syCb8ag2jeQdIHpCOa+h8YnR1WmDLlgsYA0eKy1Xmy94VIPtEIuKLkbhWWqTZOy
P+7y+1q2W+FebwGaB3zTVot7c0Lyzy/wafWtrydCwg71D8MfRWy8SDyAJza489+k7fKLgHJ7G4R2
khAaonDrpKOLyzRcY2W6AzkBAWAgSd1T1FOqjrlOmFqknhcxcid0sUXPk2XO5aGNdqSfmnT3ShtI
G9pWnT9GBn5OOvTNyGHAlaeSkLIEUm3kFON+WionN8a6tsUWw57zz2lqM/zneqHEZOsHRrUwP1Rr
UMFK7VdHEH59TjzFTBXqJcYdf3Fdphfn2GnoxKsP1FPWokrlRTHDjXA0QvuWxl4Wa+blXQFYqsd8
xNPFLYb6PFRqkbqSX5m9qoBV+Lk8GPSbI6sMzXo/F2iujPWjke3waK1Dbw03PvT6L5fuX56Poiwa
sQaWZhDYGw94Vs4ZY0o57DXwZYJGOQvP/71rB+DJlhBDkRTTgFSDr0pKrl29LOjdjCqFuRDggcN3
Cz7wkXDVDFbmEI+oC1q560H0DY/a62aV6SDoWxhmB1LQc7I1j0lftHqf31IOOq8lwSuLucfu+Kv2
hG9VfYNNqsYqUNQCLiB+8mXLEZL87MJevuqMChPkMYa3zydmaljw0uZ5eDnmPv6dXIHB/1jEd83t
kq3EdJbcxL+MOYVk/bpWZ1lqvByAUSP/+5WAOSRqBX5uWhm5/WbxLjXdNW0Ih0RTIlOHWePsnSq3
yKZUsuUrVFAV8pE5+Va2t5EZDfunxWCGpyZyUl9n+0lPxdvlnpd7NVpDouqzvwv+l5P8ni4nWywu
3vCFSsk+A6pARz2HAbqf8eqUuzS8+BjO0Cw/598s6tS+mqlALqQM8GclYp26+rJXx/uZB/gfGY5O
9b0vl2nT/XUDxsS/HIHcjJHFXANZdK+TnK9JhAjWO2FxSF6nBruC2BOCsql3+IivbnwIxlCqtUkj
ZDnXIHw4aqvE5ze3ZfQ/ODPKLcd2wHvz8r0byQxzQSSZDJswvezLCbCIwJ4Sm5x2uaP07xbp7sb+
9uTkuT/KEmX4HnwMDbObuWkvy0Ujcwww0ePwe876rarUj27nMMnzorcRP1KhJV5U0Ul+7CwueTDN
aRqu0xFXp1K0E+30HVWPuNU1+rhZ8gtcEV2sa6648fzYHMmBmEkQ43GppfZY4aTlN2tEWeTPBNeS
9sO4EbR6DbJUjt+m9xuYmBQOhvalJX6T/fKF1C5ZHJAmyCGbMeo/tqaq0yTNNlaGsvZa//ZUMaX5
M1MMY3VL9glqjgOmHSZ7haZkjPVpWSvAMqzOxrkAnrscY1pRz1ouXU45IEIyoT1/wa5KPPPFRUZe
TnDdfuU0BPPl5QCG9sGcqMQPjIB+tpU4bo9yATD+lHyg8BTzXj5myPyAHpf+4b0aYPHoXHHPT1qH
3EYsiAzwtjcBZQirnD8t93W23wp+U2vrgpYaQRh8pjQgG0OS3H064YNAXWhn4dsMNPmaKlPjLgME
5bnKuDpEDn9ZxlTrnhrpD40vztNBdQhn+SyHDEb6s5pKQmeQPn24eNDddbKSPl1lEb60AYQ+0JxH
X3+tFl7dIjbwAcW7JicTDsLGEdG3oKP4WXmLmTML9Bd4k0t6UFFrUclBlCmrYaDBH2ae81RkXwzR
F4cmdqHqMh1XsaXYkxU5I2/PZO2nVV99Sbz7Zy890z1bC5QupnCNhyWyO5u5lRcyRyzlBBcNVfR3
oJUjKjHRRLW/q8BlZjYvpZrJt+Z5LlFd760As6zdzIRYquuoW17EA2Fu0RzXP1PdNbk00qNqHp72
SRaB72WcKZyVDc2LTO214bpTfPYk2ehqA5+gMj4UcnL1ZQGnQMOEeAHWqzKPZUkYFIEW91oYCXCE
H0Zzar6u1zF0oxbUZOmSYnKJ3ms4o70YJI8QSuQKzRBQmm2zPmxLsCVZTrjR/suOCEoQLhdWD3Xf
sigdaDoRrD5X4lju4dyubMiZDvVSw5+sQO4lNR+FQ+3ItShrGsW9Zq29rfjOHk8omAmR8T0i1ADT
M/cVl/BIyqGHViRtI+ZKq+ZTddU1bGrooXpaMKS10mIJgsOf7kJHMJeJKn172efyYP+5CDnBRBf9
/e7n68+rYCWVKa3hiCgEqQITxMpdfmI/FqdP/G/wXEG5GD2vBTO858wnEauDYd03/YriXIk3N45u
gbGGI+1jfGaMY6Kqn3nYVqW60qgjD0Menn3aA46fUR7Et6hjijD8fkPynXfC5JrixRXUjZf2z4gp
I2Oqyfb0CTVL3L5zsxikKUpf55NfMB2z7yYTDVeoNg+7M9Bw1WWCrl7dgTm54Mm9JDqEqOIbmkDO
/qElP+LsaOVi5WGchx/dPUse681cQkWjbd4UNOCcarhTEyLdlrdlbQaxxT/h5pk7VtF6iL7uZKSd
WBCrwIc/shT0iPDK5oKcnGmNAl/ELvKnDobekeRF4DN2oToxKxYBak5bQ6GV9ZkGc12DWjifHzUh
FVtdOLe9b1Fl7h3xJ+99/NKM897qttXpYQgbXjxWwZsN/uou8rpDbQiJZ03tSOcR0v2s9zOQzjo/
UvK3v7OGxJ2x3d8NZNoJJgc5x9dnukEkA6wBmzBcLJpGkhxtRzFT7X0U3grtLTacbrm9GmbMoWFb
6incw4PWwL3oytAFAGniKaCD67QHb9iO7vtF4ZmE92v5aPXGEt7wX9st0fKNwSPnuscwVIvWqYnd
BZaFh0QIjOfBScV/3JVZ7H0YYWcyyVQst8Gv6ydUj0vwlM2MWqvkc/bWZa622RHT10rQb3kF49V+
0oioREg/1/0yAx0puvMd2FBVT2gjs03zXYhrk6YJA567oGhTb/OnVgFpx+FsRB1AyO8Aa/dWNIGi
2cGDyvlCrT7B+fWlwsSmX2ooC2klUF9Sf/s5Rj5tr1dNON9MSCNOwYSIg5f0rBFoVJ4IQsV1U1T1
fHjlUfxTJoC3nggOc6pDq00acRNRuy45dbZKduOPx80LE3I3b9Dhyh0MPLdH2p5cWB/+tS32cBY7
qCC5/cI6UAwoXQAO0ZYooKdeNuh+TCEp+mqd5UyBegRwadCUAa0xWvdnoPcVoEaTCq2WDd6Z2OqE
veGeM5wv27bLLodaWiA3y/1KQYnr5shkMxeNknQYWuomJeYPaLTw1H+l95qCqjCZE1cfci2xHSbq
eYM6afzy5uJwHgZ5jN6v0ehhBPfTf3/d0Fq32GkqJwtMKHPtSDImDROojXOkD7gJucJTEgTuE/Ui
8skpzV2TGk8pix/w0EPgb+v7xytjwTxouaoDf4ri/SXDK5vo87s+GLAErEAgYMdnTxFMw0K0RN5f
Ben4yEQOHr2e8u59MpHA2FCw48pJup7EBfAdRBZe+Jmn/YGV1GxiAeX915xDFShqQ/vpPsP/TbmI
KTr6tR+nKMQ8VH/i2j+SphjYmUGB1cyuiQQ162nI+qv7z/7qRtJMhFlWIdoqdM9yzXee+PwZpiOB
CLA76VxMVmjCDA6pqcOewl4sCGNieDJjUGA5RuFux8GvWZT/AUnYyUSXCbrYVEEKXtNTaHgu6/Em
JCLgJaTOZWPsL138KFObxySIQKfHOvAYUHCBovghjj1sFodtz7Kis3sR3LB1UhPrazNeAYbFuwyC
EUwD5loeKUs7ykmHK4ZOpIOsCqDBTjebpwL2onF/gBe61a4MPFAUVfAyRGEWVzfbjE0XKHbH806P
P16Xlyl85TMLDcVU2PO4tYfxkahXtuM4Y2GknFDKvVq95vvsdCE5PPNrocgV91VCWdW5DRgIwl8y
pUgqyHitP8/aul7Zv02QWJG8bF9d6aixwupgPahECKjFSBp70IM8KExWMRIA2FI1MYTLiF4sz0cq
+22Sdgfb9Cu1Yzs8v0++irNc49axkS/ZqgQSZDc2Qc+ihZtacNEX8Br5KJbukatxd7xZ+r2koj7B
GD0M9GQa3uhWTm7ZDT4PCqmGSHWkuo0HmvUeCS1/+0M/cU2ftsqRLa6Jqhyoc0a3CKNviw3GfPHB
hQ7I3b8ULV5GBtyLiibdquI1znuPuQ+cLqHa52BH0/KOPC9fZpOSIeuMRB+pIOHmCMu1T6KoFHYd
hmJs1UH5/yJ5XJkycE18FmWEL07yakc4JIjE8S1JBiMJG1ucExwdsMUmaY99MWOBNBFW3hzNfKoa
x/s2NNTO7vwpJd2/Ry+yzEJimvax00ArzZps3PiMpBLjD8gNEjXM8YrxoDrdXIhDAO9F38Cbk1BQ
JnkqFoXKTY3/xYcX0k74nKgLsEJx2JdDdEpV8hAis4Qld9hJzNGu1GWXDDi1Am+H+UGT7rIbetTe
jt6tJHVBrwCY3tg67bKegOXO8ZcQ3vZ5158FRIEiFJQUGaSjY/cCu/2TQ+AcnvNM1GV387jJWam1
clB9zaL5WyuxUqem0t6SqBi5tNKDO6ETG3JBVlru3wO2BIXXY2Z4UKf3ECCvrWywMaPAh26h93zO
4qeBgGfITnxe7eg/+FMxvLyIaaij6uQjUac4ldKpgmi0V/rPJJoP2Gm9CYorJkMpqtrkkqt8gi0p
ftWI82v8NaxW59HJsTK3iPxIXcDmSmdz2xkt2RZv4Ct4n+NceFTI3klqBGa9ciYqMO2G8J9QItYf
68ODLHBpRCJx6ttR87yG2QOAEThBNRpc4YKgapGqPxayEw2eRMSX5R4fb5I+B355KJyd9jZVIMWd
6xjGtmyv1rEfea/rN+zBMl9qjDkfcd9L6QbK3LEezseDSg4m0wwRileswah3E6zwDY78j2sqiHEN
KJBcvbXlJ4qa7DbthDketzPQUvOPK6J5rkDMDxTFsTfoKEfBV46pX4Y5LLt4nHG3M3L3U/yemfY4
uyj3YjkRkh37WaxBrUw3xsmEkbFXWiJDzS3wsGolq4ziOKau+rcgb7NYXvwd0bN3g7k3GZHVTPev
mT1dg/mOQCGHmQLfAyF4tvLyg3qkBhpjB7fDjevR9drv0diSdeUeLhc3irq4pCTYc5NXMEOcAU19
uZz/grIswmWMiriCp6Xm/rJOQWHS5b9w5A5ox/IpdClW0oMbqk7guNa/ML5nhy/B/phzjBcLipgM
fHLmfzSDH4wNPNDTeF3hGnGhFB8RwKWjEuyPrl1HGppg5mFyhMmmWXUCmHehZN9StxmLg+uF1fe1
IlfSckPlR5mO98nW8Ar9x5wnwUVhJdRbU1iIjCLIIYwcUzfMH0s1DT5NvPvMt7hqVDf2NGJgj5Ym
myRgDF9mazsE/puwwMa9QpNV8F2dgYHkscAT1lMQ1ZIhaYbfeb1Jo+cfF9KPfQxH+c//qMOow9Y2
7AeR5Lu34o5J9Q66LCxW/oXj5HZw9ppw2+QWUnVVAg9lMUG+5Iq9DlLf3Cr57dO8ZmXCBOWZpHDs
ZvQdWwZQyHCPgSqNkpNLEvqlI2YzqL2NDK1l7eQGhf354TCFS64dojVhHsBhhYjlDIQqi6pDQO0s
kjXqGzFLAsfuBkw4LuTsqC95BcbAoDvIzJwvJ/ijn4YcB8qRc9nz0Z1pyNvpuoTMw051lWxvYX1o
jiuAoQUihejOh81byqqJk6dWSJc7a1AZnPKkSS37Kk9dag3G//MQLVLRzkKW78DQHLyIwPh4wpzD
cMaWzCoEGpNsL8pChiccFWosggWOkGe1ZKvIA+a3ed4zB4b2E+Nw/FqFRfz0Pky4cjrhvtHz3yTz
6zodFETCUEfGIQMgjlwOEtCRZhaXZhrHQmr458YqyAU8p48qro2v9rwWlvygdjEE+ilsS//eZxL5
4VgG2pBg2jjP+a1SlkqREmvOxs71LXsWX+tWtzf2y2sTvM2g/EOVTLLdIPU3b7AFNPWWHIjoQ9tW
jhlkVPsQg3s+EqhRkSU0M5mvcJ8Tb77zvonuyYwKtyYh5JF9UW4EnPYtpe4I8TDbz7GFzWBlKvTD
v4aW6HAnIRK+5/JCd+zV8shZlF9p+suiPLVPq9SbItfpxX493w6qBbWZtvTJv6Yi6CsG0+kHsxSr
fbjUXpZPkfMkmtM0pObgWJqyeeFlGUBUssx+ygDiMjzyPFQDryUR0fRUQ5rlelV6/1OQmkYmDvgE
WeeLiRJrmHwEopezBvO8LUvOeuhdtyZzPh7RlVFrryENq83uwZwUdhZbqvrNm4/t+n/Fj7ujip3d
YBkLjtYmfoVyaJH7erliNkErxWKUjDey+zuvJ3FAVvbuZfZIWoAXNg/WYPXkF8pBHQnMMwA/kDJt
JzFCezFZ+fZN+XdfDAr7JDDKyT2uHpBF/OMh3dBuo9Q9k8t+bkNPTwSm4seoKZMz1P8upa1MQVUl
EBd92Ccp26T7zmnUPBUOIYh9xI72wbRuLwqTMfeiqqtllQBR5RRBrcilQRJBSePzyDfqf0KDhrty
JGqDj6JOwjRJpvyiN/DZvirRMZNvQdKCR1cOiAY7wRW/LbfhbEGt91nu6Dl9OrEZGUtEbG2Q96zp
V9zZhkYudwO8EbzzcuJsB5Sw4g0L0N72f+mpOe1yGFX+c4w9xI1erc3x1sqeXzkAk8kqwNGsB36g
SYv8jY2lysCw2d5lvpopovPsF3lt7lvqCP2ctKaJN4eG2q7iwm55tcSymTikXyhlAC7eYs3OqCV0
2havaNn9SRpDDKJmNePLfOb9XjV9l2A3ltTm+Tffe0SFHVODLk1QKSp4ZXTkJ3uwEIRwxJIqBRpH
Kcl700AxLaNUIWOZK4ZzVYzRHDX5ccuB343dWB6LY8f+DHIAOiPGFqMEkybJhHrgDEtkRiukkh8S
m5/+07mOg/K+dACGeFEHaJ1JvAsPdnM9uKaHIl33skKhzDwlM9O5523esclBsbNtqSUkb3lkn4Io
RwfVw3wiP0438pDeoxmq6bwFwRUWZRzV4rm7mdOdOYSgog4UgPCGeON2HIgz/2YxDaFzj7NKatLe
PQ1sHVz62NstHLVVOxN6OcQ4MteKN00+zL7d/j2EOJ5pvFBcoO81qmzW6WAHwgW/1aUnhxix2fLy
X+czF1L16j1iuRQ2cTEKOTyzqDKQQvzXWBBEwLdaPvOhSx4HXbonyiuvlI99rxUIbEpEiffP8C3n
t4+9391NMT+1lvLTlk7I5+/9FIRxlkxTtc9x5HCX3hnEfTC6hV6A4vbb/wGjd/qH+W5uShhcs/uM
oq8bC49KHLuwiTWcAMQv/aYmgQKIdONqOR5LL+SYg1oCJJ6degOyAHjCQIyUt9lBI1ydnF+tnAd+
g/teeWhnUuGB43SYF7wuVF4kMoO2b10ESoGkRGnesDgj6T5miH0nb0njDRoPl4gJlPG1lKlooGUX
d4mMQzIY0zsFQz1UvrnG7jSiSFk50wArjx66OzClcLOyPTCqD+MIzIT8H59c3EFIm5JXs87/JwIq
cW2Nc4yYVpel6e43ju9dwoL7sf3jfWJXNcPkaay6e3zTDtDVZ7Hzup3ARuwWrhSjS/pqA2iNoDLL
lbyru+9SA/NVO/VeZeykchCTBpbe3CMMEc6Du1ZIDI3TP6k9A8MC0O65QVpVVZm5s32h007ev4Dw
5iP5DDbVTxBiQYoGJc6boex8Y02kVouEkTp/LRekfVRk/KgJBzikpwTjqcdnpbDu0Yrn/V91sFHP
MOHYckbxaADmlZtc+3AR7PL+VROU0aXXbC70N1lNIgSRkY+p8x7GBwiqbWAOGiekNb2ZxsN4nKuE
Ca8LwuU9CMcX6yaPlfYStsZdb18VlXQ2AV25oxyPZYOKmNuxD8i+JWeJYIcM5tMnKG94pWvY1eFz
X6eMAo6ayXdwFqd2sT08TUXGisxE5ypzSOACokgswUc0u2CBXUaYymFWdZImJbCnhVJ0CZe6feSV
GvfiBWiwUNXgnmB/Mh50meSUulAEia8w86wel8Ge23mNQ5a1lgRglUw1eeguNKBD3h772H57UWqn
69YYkucdA+ESbM3796AYiw/ercKmCXVtXaJtQydzegbrtLSOizpdt4l2qxmgzYRn/AfLfKbx5+BK
arbpBfJxSezXnh7pFcRMTxqp0CphnfAsHBdT1YlxXsZ0FbcchPxldro3w6xW8VNlC62jFA7tVPoV
/6W6pv0/K9qzvY3X7osO0zumbnKqri8YWQcr6rmyEnXxau9Cf9IG4N4UxuHSJtf9AaZ70GDuptOQ
p4I0xvIsoozqO9SZ/I6b2ba3XxfMzJn4HbekRE690kcEva1V/8dSp2Sz0QLkK90oKX6aSh941ZIK
YsujZrVyYxXIIg4alF3j1wmvvkXE4ptREvTsNi6OU3NiPiGxjj3cG6qJBtwiR6ACsRYpglWyPP+7
Kg4PbsKfobNSD7YD+AhyZ7IJ1AdAw5Upui6PpkwkNJhi2AP6ODLnrn9kfqL5zPSiUDUm3tsXxkF+
SzCM61j9xjtfDsC0FRvMmdsSkpCmlURGaz+Lv9GdYiv8nReB4IpCP73/rxegvuDgYbmJRpIF8aLm
SMFNQJVmfufmukipuWA7t+f9mleJmS63OkCoqXnV5MLTQmi1G27khPXMx/0LiZbcj/Tlt+RMT3YD
DwaDw+qE7v2dGcsA4nR21v+XHuT4uyXKhzJa9kRyUh2NLEp8+ptHr8o8aVdmlN74CoO/Maqd8GN5
4h4CUVn1gQNx53iUDLm8C6RgZHZa78IyM3vFlht/Jv/hJW+04jk07HOpQFTLLyA3AnWQXgcqss9e
JUYKC7K2mr2ahVMn03Qu/rSq5tnG+vPaBrG9SFCujVYN+soRmGG/WfKATg5k7BWInn9DSLozraCY
jKTV+O93VWNxALz50LTIhK2ksxy7xjMkQeeIYK7CSvuzcB9uLOLCUFSxdugk5x0Q/T3vIZXtf6Tu
2InDcSs3OhvWDD413vMndySqk1liDdY8AE2bB7gKRvn70w8gSWEQYH9JbRDCkLmcfta+TIK1XjZ7
lfs9tel4s9M5ciarKCBzNT3MwwSwzxDRbildBN/BRHYhuKC/msaoVc8lF652/vfvfToaU8SnkmRR
xe5slUmxmH9lp2BW4aWtD6QjcrZjy5918elA5WjLGA9GecIg91qyEjfEK+4M2oKqbAElzOB6Qdaj
h3nA8sxOy6Z1wC/W13wIzSJ3XXu+Xgwe+gLE7Tg9yWg5gPFU91fDedOs3QPfbhTiisqVBU2QqJFs
HRX9FpK1NgepUWbE1QmSf7GwI8ZYYcsb0no/pUgsQeQCmKNHSOyY0xiFzab77JZJmMwo3oJdtxAY
DR1dz7qQUUWvK00MpKLHkpGXDaUYZbpV0x79t+xcMGed8fdrHG6vUsyhbTJe0yI8weqjfrAEzCdT
53gwhySCuegNgP5p8qGb7ItKA75LU1UVcP2IceOCLhtuSj/RwAFq5YQ/mF105m4VQWES4kftClGE
z80cJgj6Gcx2N3/POYG+9nrGZJtWPYWs8Kh/cbNuq06ioxc4mDgBpmrhF2eypZx5rA3/M3yOPfHZ
ozFnXNoFeOgvUZZvUdVD6k4RKhFxgNJN+Jhx5sxjebluy/IZBYwjmylxEvz0bKhs+IF27Qns8TgV
bll0rXI1ooFZOH7+g4cL0rCKX90AEzn1soii6Nor/n1dqdid1ZYIy0/jmfCTY8CT8BdLpjOUmIY2
E7Z17chBJc4FOK9GcUbu44v3Vd/vXv1GY4TJm3SyvrDsVUWqZSC2XKG4pDTTgqD8sh+4+FX2EP6P
9mTT4Wvlaizgap7diRmSxwGvIU7B+97uaZy5wUIIOPhUBt31gBOkwP3uNTZuJtkX6qi43yQiwzYD
TJXZvsUBN8tHY2Tdb3MjxKuGdcymgdvvdO4RO9nFK7ghPCJ4MtaTwJUOsFS8jaQyJagxvNs+9Q0V
D3Ton3VBLN+KRX23UuyExzIotTTpiw0wvpg1APhYTjJV0EMWPloFAwqF7oQk03Oh2O1jhgrWB74t
ETMXQGMKzNEYNYLWUp/PkNsNdN4HYRj2cfpR4GZIN4HlpN++TFka9OMbB3ga2VqhWU3X+tevz4RB
sf4aJKYCpQTVp61NH6RTlLPSM/aNgWlk9G8GXYbsg/bW1RrOAzS9ovn0fz/hmSgi4xRee7NjMW9V
8oyQEOVxn4rIOzTYbkGcX2d3elnfUYR93ZWARiNc9UjISJlhVKnUFNc0j58vAieLZzoI9q6CtKeB
AwT5S7bi8tMPM6RhJqz5/b6avIYSbftRkWInByW56zOsW5LfAt/GML5ZAsyOSIG+srZ0Yi0AfeSv
aQKlHfFC3zEzIMtKTA0NGGRsk7NHbj+ZQuuRVBDYD3FKYXLkNr82TJelAWADpRr0u3S4z8ubRV1g
zA8iEXJXuO81h6KdXgiVmzlUvKuesP3z5BKerPSxNae+VlftaNkUZSgVNBiBLEFnv1JjxvHiGdT8
qjrGauL8Smidi8mTyuTg7V/azJfkyupxT9lss89Cd2WrR0BC3TNWblnoy20lEfB6yvGOMDv9ZgJl
Q2KQ5XIGzsLTxN5BnKlM1Q50FsEtKzgAkUKUqwCqFt6gNWz0pE+HOY0inPybmDnN9ZKDPxgPf3HR
ujKOjS87EUGNl4P0IFe06w/5p5wEIYPwtS4701NyU4bvn1avqHEsKckKZlDTxfMMvaYxsNQCu8tB
ESmpBLd8eh+RaD4eQ151SC8go1X1NazkNBkDdZj19pEnA20xq1Idj6KyiUwN/QU3cR7ggeiMUVos
WZuEKjLn1W1zp1v+ovqi/XeMsqhYwBUnQ99SIJNFBcMIc5UKLP8kCehgYl1vS/3AUtOLCRc3drvL
9ae+CQn84N9pkIxkRy9RjGVp7Un2MfVcpAzbdv8up/uJOGyFF9Mw+6ZuJzOXoHkH1ICHY24pgYOk
G5Ren3QeTA1EFhIL6ATgDad0NtP1N/EJXplLBWaAAQAv6tTxfAue29KblRWBTupzXP3jXxAwvr9R
iPJydpEY4NQFZVOwH2yyZa4rhO/G4EFXIxYBtTofpQShdnR6aqj6QlD5dEPqFNJwVlYhjMIf+EZr
vvcTCSi95MpYsSDwNItLbv4muV6/wNNCVdWExJTKsUpoUSbyHiukNhURlrWpr2GwBmqI52hcHgNl
s38dxvaLQ314s8dnLfumZzXFO9gmL9hqY2+ESgjpzPptG2UNOmH1reW3TK+8wMtIjU+F+nc+Qdtf
fEKnfnplCbloXpkiyGFevFg4sYeNJyHuVLzgdrWr6O+SlfhTMNz3qOyvdG850f5bpa9HixjyLGxK
t9kSPehYHlZqO8TvpdQ+/IuhdyYkprB0u8QS1WvbXLC3r1jP+UTaiwFAJ6s64ip2NJBwU/XvI1eN
+7fTjBLiZfJ3gmUpk9JRln5uDhYN3N9vnnUgnyfjvljM7kRroE8mEl8NjXxn3NdL+0hfUJMZmQJU
Wm6ZUjaq3z+a8oS2luG61p7leuMXN7sdZoDeN+3OBCgy/wQYYjbDB3jB9m6/vwL1XFzzNX47MSru
xIUNgOws2edowJHf1BQhp1r/4FXi0DRazQvL98O+ibfIWq4K1G5rHYM3M+sA6xikhelQvYU3QLpN
nlQNbBiZArXKaVqvq1hbGC6hN8N3o9yWTJprMXrgm+0uY7mBSvqBtGL1OiC4gWtqYE/1zNp7z3jR
682+FI4e7aMeKGCn+koxOePND3D1dcnivuQTXdzKMXR9Yq6ajPPvNumiIzVWjJQvxzVg5wyQmC0P
oKbKzjjPWQ2wNiEnqDMzieZ7XPENaTHwYzZFESGJOCvsU4+qc4LLBODxObqTSGgKNxacYZHq1Pqq
jSHrf5sq1zCuFc5dJ8iuvsGAKHYX0PxQupnWPXj7Kpcdym0SBrLYC/cewa6NJFh10D4pb8GjCPW8
5bpmCu5mvsCSKMjjuMLb5TiMBZUm5dxsP+n/WCm04pDFkJzU+WAc1s8Ytcyvw5/dRVyb4u5c2+Pz
CDjCBMSTdvyWC0O5/UrON682MAuRmh0wM/8QMkQX7sNwRBo6BdqWDVVTosI5P6x1DybFqdF+B5FU
cwlvfuNlekN3RNgL5VvoxtiNbxqFmys+R9nwsUxVzZbGwZQmo2O4g9K17/hdhTd7mPL70aXq0kCC
u59RPpfzOIqG4jX/MlaXJN4mWwbvTUj5RFmsNjOdSm5TF8Ix1qChgSTJEppdWWXcNccgdKnKdUk5
XT5EzmQ4zUJKv57omgHfO5BaGGiF1nLWaePDJ1EX1dUXIQDCADSRJxTfGXoJcr5Z4isgdTpeOxYE
Lf7or3bsQQ4AkChNS6APjVKx0dbEPO9XZLegMq2B+QsBGd1reSEJGSiYoejrYHxuQJwz0bA8ObUo
jMAwoR69COQFo8Q1tp9unOZtdxlD9W6frzd3xpej/uj0zI1q1Doqy9uXOqjmrhhNZmu5Jj7dY3BF
fSvx+rohaU/XezKK2+8jVyPGbAymyu1FuFwETpxPynTFHrDEgJZ56LQf6tfyLe2TejEZU2RkK8dm
4KNffGiLBNAJqNGc/Vi+G0CgcGD/WOfFKOjLeHzm8V41xsMyG6xbl8MdysShk+U3m28JTlQLPRki
PCt/ncIeVAYZsRYeNEs+L+0+HpWddfonOJouYqO7b8/zO8CQWDjbsn6H1218O44bNcequQu23iZL
UwVtltt0vdKDC1dMQ78UkMMhFFWcTt8Kmr1JgAz3b3e8zVI3wLpkaodHkQk73+KM+fZxOVGZeNu/
D7VUd9NLf9oLDNZtXXJg1gi2ZWGAR9wM+RG+Qifjn/GhZsYgsTI5564zzLc2ni9EaWiOHSZog3nk
QNtcGO5tTBkSvkUiSYZlnYrAA6QnKEa9klGRO22DqFBw/w6Ioq3Xuf15ego0umx0+9SAwVciMaL6
7jdySTFQiPSzGFRS4gpluJQhLeg86RxLnJ9KlUixZjvxksqhFCTY9c6tXOgajHrWOjFs7clWZjZn
dbCS86ayb9RPYmOZwpBPw2OK9tLOONd5ciKph51geEqv+bQHQEDUsj0MmJ3SfA9UttbzRJy9UVGL
+VpsPVPizSX20gNnuZb4XpSUbjSNUlLuq2viVn5oAXgtaD8goCr3CD4NtPOUIWz2L8Yrqwm/hMji
Y9Nw0ZVmOdKLReZypWtDstr9rueZdWdT8m9AyFMhmGDH9BDk7+iW1qCrDuyhYpkCjSiQZCKW8+Re
krvE8//fHxNe2vTUZLSYY/18fosqYA2k92Ka9Sjg8PmzZeEwjI0UIDlG7cI2H/830ywckxsTgY6D
iz1lmUVgl7DsVJHm7TdAL4oL2UQAia817w5yUFGiNuGSXIlq4J80ZECID1wfYvkf41LlPZK8vb2o
p7ZWbSO3MMDXvlch+0YTpZaRCAqrBAZFouMWJghaBgz/BDgD2IHz8YkoXvW39GsNzMhPqaBgHezH
u4NOvr1XITCABtUSxC8qz0D6CClAnZEXT2SCZW0ONVtRDw44hUyF6JV8r26hsX/Un+BAVFuWk0JU
2/rj7LH/EuCTPrhEj+vAhPsXJ0z5Vg20IgGg6cJGDEx+BzI7xA6obJ7GaZRT29PnYe9sAe4e70Ud
4dmgQzDRSYd3+Wu1OoxEOYC7Om4u6TtPpUhTV/2K/Bu+d3SjCRZOQ5Kq9Wg8fStmwK7upbXwdSYt
ZodfKPlsmzl58pkg8nf+NvHrzoiK33LPKRA102z7ZFDrwRXN24WrI90JrSAVveADzRkYGA4FnRZe
+l75cZ8RQ9tCDgjVHsoByn1qm4jJfbJs95gUsX/mNN5/H8Vh9onAIIfXWgnuUSSpGxag7xuTvwwP
70BCblEjI3Bmbe0d/ugJP7pFecUhumtQjh7ZhOgKE4mI1hFlyDZbmb+obT8qdVFrIbXLfgvPW6ta
y5gs7DIsLkZ9FSwmiAFTYRFKr3VYZ+bEzINWinAxrM8rOJVnwWMm+mNwv2q1+RL7odJC4blGuZ7T
Hjq2EyXTgRcg+tnzrdC/vJpVccbRH8uy5n3yAe8KIvPLocgkdLwVqRRZWrH8QRF7n1CLv2bxORET
sFb2i7/6Q3IQ5UtLJaqW7e3QiK/EqtAGD3DPyJ5HS99muILk4ZlqmhtgnwPv71pFos9s/WjiaSnT
Tmzp0ylIyD6BEtAGoItr/E3y0uDg+LeB+DKrJ/h/LeS11iSQcX48bw/2qpsMiVI4KSmPnQRSy3hL
Zbx4jODBP5aAePaTgQb9YGTdcxstEKNyCWKpHPcM3W/adD2F1xNoKKuJMYZsKaEdTlhwtcaYnqDi
0FJnd7F12gDWnLsbhpvozhpgdyBvOqxKD2F0eEhaqX+94iNhFJKq5gAcp+WtQbdXJTdZKFPWkOUW
tLLRxiM1T6tDzcpWHGf5v7iEr4LGnzjU1ouX90VrnWgqE5Z9gZ0ZzCZS8lhLfgH4NTei8CDjwaU2
XhIsQ0PyzMZKBWguF1fviY3LCeMStp5jj7hDz7wGCJLF9iMlbAtD7jrF7E/tgljZvplatmAF1ysF
ZimQNJMxfV8ogNXUiW9nwEG7qqjcMXRzllXWVIvVsjM5+yrc2CC716AV6sPjsTdbCL1gM7bHZC4R
UtRwUC8ntUnkn4LBFn90g4HwOQcgUq16mcN3MClbueVf4rdBzFPIqbNQ63pQpm/pM/yMZYAzws0j
Q/2lS/TpBDB+NMEKKed4ofo+hfTWJzhxWhnnGMPWZEGRzGpFBh8pDhVzBoZgH0wd/LVaCMQR/Mfp
AxleW9TS+jvIXQWgKJEfkbUC+Y9lynpxFe13r8BhFkba34XEvfX8AI8eAocFHdnl7YuolCuaU7nV
RKJpv3a5GYZcCSzLPWc+ghGgOWVb9FaqtM1Q0xWpl+fQjwrgwgXpa8CIBm7vDjgTT2YniqmBHEXD
9V/Q/AlzRUzeFOQ4Zy3W43z/+V4SHfTZR/G22qCffSbzAfuBjVw2iwoN7hIbupygWIn6Z7D4tyin
mwSvxjSVeLadS/IqegeQ8fx+gwVWgjtwfhVwlBG7ng+izeQihv+iItB5NUKDrljbWOVa7H+ut+rV
a5olnC4zFEOQR04fWO4BNrPM0lO0NZU4zntzeesjHm5mZXrQOwF7DC1TlPCCZ7vNTzr7v4yo4NXY
+XQw+57vZ2HJf0W7A6kv7KbqzTuQnEykH/IcxrEvBQ6oGZHXeG31BGNggqhgEKYscm5gDDId+IPl
u8v3JxDlVgKrutjndghDXZ3k9Z6lyYZhLvx7HQ4KMcZR18vWl5BP259rFMcTFH50m+VlSduafutu
xhZU/93ZlPt26PtlC+iJrdL7ucXGLGFH7V8DOt5O9l5fpvcSBVd6JuTaBTvzclCB78I+zk+wmaN6
nmcGS5hOnOhI5jPtErSvpAARV7xEv9BvxV7cHkenAQuxX7vFeo9h2LvQBnWpF6OXLywFJuah/kxp
pIEeW6rwehwC3hdtfrZ1j3jFX32NAgMe9wQpfFy5T7wfw6ksscu9Ab1lBWvrqxUrWZO+EzjT52FV
iIKo4x2SOp/KuveDW8nVLNpZMygtTaWwhrT9xhI7mzVRi/iaq2YKP4WRXglkFt1PnHtoVKmJkmDg
coyNt6GI1Q9mdRp4oy4sGSrgBhQwqI+FWLhLERLirzd5sq4HlflgLun+u6CNI8GiWn5xCjtegIs6
gaE7bL9Sn/3QmUiQgL2EZF8YNHtGRTuCc4mAk2rf3J8SEWo1l1GmPvay8en6eCck4qX7LqoK4Rj4
3t4N1qfLMqGJckJ6L9JiV8sdZ7lAx4Aq7pmg8t5pMEndloODP2iIqLNj6+dk9Wtjm35Oi16qT+sc
mlaQW8Kv9/d+fE17tgj/jeExxltOkHHvOZVYzbjnOZ5UJ2BnSNONfM6tXvS24K5fP0FI1cqM6sm4
ujD8dvVTvhOjSmSNVA8m0XzK1aC0Dd5fQKToJr0NaI3dYq0+QXpNld0TyRpbtcg8SlNMlqDFLQ+h
2SIYM8meMOg6nNHP6BqlSO7BMhvcSMOspWqOmlbcsGM2FOFNe8GbOBAwQE7BiOivZQ7j1Xxyx006
jkKEPawP9I+HwOWax96ZT8oQax7fSYAhdQKH4LHTCCsyPT0JOnNLpFL70XuYzljhtkb7wqPVnqJ8
eKreXjmyBiFKpomfr/4nzNLF4zysR+4zT4CpdcOLNfkQQ96QuVtrVe8B5jnzibqUA3UZm3UOzYGU
s+xxxabddCOy/kSbB0MgSfp7aIXoQC/tljNKRw9z5OY4zGhvDH7bh/703Hay3BHN35LHcpmqNfB0
E6Xl0triyZTfaH+g/Gqv9UhL5sTcqtMsChy5UWIDSl6dNsPsjrRtM7O6bITjQ8UDwyeL6vOGycJb
1q4XIbVqv+KJffhj9sDYEjiiw7jAXkJPNpSk8WlJKIwCPDvgnWaJxGaLxAuerOgIUUWTgPkKHRZX
6lDiAnZRA+lOYEE9Oj3mDlfnlyn9uU6fNlCJh3kAJXtvGKMaC+OyfyPfpRCxGxMcYj59vo7Glurw
+YNz1zIAwvocirm5UzECAFvq0dIwaQ3Qf1Wp2LoEAd9D+EBbhGa4GxNGtvLwHCxKJJNnt86Dit52
tD8kvxfKWVEarL1EFtjbmBfbK2/5KIijDADcKULv0hWNTvRp0nAIJYDPfz5180lGg1X6Vz2U8ElW
PStPHi5sA9k9o9icUtgBYhQ/2A+IT9zMdU5DTZb6fNriEPPp+JHDjG7XxsnaTNSW3tDtrUnbAiGl
46dtXpx+eDc/lD90l37djeV3g9bQRWkM5eDOVIj317mdxVSpoo6/rSV9rZO5425aWkY4sRYDxMAi
7QGF4QzSCo7+Ohubo6hb15zmqPa0nxw/aWhHrfsL0Xgqb36WBCw1GBRbZ2zEUEJ0isPwE6ll9w71
Mfay4mzlhT1qsuAEVwl6iuvrJa28KbZKYl5a0OWLhWriWYFgtMXo5q32icPR6+MHOfF0LwO8ExCt
C3XtFxZxCjtR2phURaDUb2/guprMmR2YLHWwmIvhk2pZ8uH3Cq7agsC0csv/NGrEScr+2pPYoTFC
HjsuPdE+mgXSoqF/XZA9AKDvDv/pjHrnyG61a2kil9tsQk4KwIMM+4rwWBoj/n4KZ+Gi3g1QHckH
pBEJPl8Ub6xgcdwXe3zheW9tpEIoq4gDoAUfHZdDHtTUE8W2VI3kj65d00wpJmT6vUhBWpMAqyZk
BH7qwx5RLYyppbyWwzUztaYt0SU4U7en8b05NxkmANV4+3ilYCfH5hXxlhUoXMmhp9odGwjGSDlg
6fxx1sHwsoL+w/R7wtyR7H4EBPcMvFlXmkyWEtKMpwf9XmknBYmlEUZgAFpRcXWgNHEZloI1AGDU
+ZVhmT7T5we+fJu7aqIiiTGlKcQRKdh38z+PwNjG3H+/R7M587EPm4cNzo+CNbWWo0jlSE8DLG86
P+6b+HEk+cmFf2TIOo7uYUp6UQpfFHe0su6Byx/9Mp4UWBheM4zw+aj2+w7XvDMN+CtkiQyywmXp
7XM6G0hiXChwPBPymL03LLYXs/EOeCc3AgMpKfXrATnzGG/3YaeA2kw0/y7atT/iGk/XUNBemhaR
Ahgu/7krqwPP4R8A9SOLQbLmpLpEKE5jGvMNx9ms+4wa+S2A1Lchs/eu1FNtx3B9L8qfQDmve8IS
wfSJatu67EbNrRrEpFe8AdkN+KiEkR+B8+SVVnwMjE0bAdj70wzLQu41miKiU5HT1+k1JwmMg3WZ
8jlMSUGKnoyPcZVrAh7XTqG0O1eopm3QMRTss+tk5Y3yDdlOOTvsYfpPRZNQS6acq6JRIHyMJfHE
sLwtcuQI4+4SPvRafGIz0PbVJNAcmqfEBuk+I6oiBPn1PiDiDPwsl2E2sK6zuq0qNHlbBSG4v360
2Sc+H2+vi5hfR85Sj6uDi4vIdNY4vGfUnMblhwsjQFhTkF0fVUbPqYpTZaCYRuFGEa325Qi6iSaE
2FGE1fQztloWP17B5gIN7IY3Oi+n74CYZ65Y3sYB7tb7bQ9VCj7M7dZRWSE6s+TwxCCtUScKsdD/
ARuljXti/n87QKPYo2ggsdA9swlTxQgRg9nQdH3C7sUZqueDH9h6yLoapWWrEl692f3ep+10GkjI
ggfJ+fIVomutTNZc7ubfa5koyboBRnjNzx3ShXTCk1EzNpQuuT6+aKNt3SpMvEzJcvYJh43vkcoS
LcGrlBiojosCRqDJmSax+T6iVIRns01Ubyz6LOfalFidLSJKhOPjGp3MZgpzvIQ3KHPsdfAPC55x
Nl3FoSV+dYRrZVmYfB6VWZlnE/74mNKZO65Do30TJqdeYawUBFrwpf3RjDiGnZCMaZYuIrrNGzgV
WW85XKBJH+hg8g7CyAa8A7dIVVHwm38EbC/vxe2laPsZlRUDqY+SeorW/fhZ3hnXADlt0fnLfup5
kK58iCAFqHOMEfN+Gym/jRsuX3IOL9JR30QZTngBVA76P/VV9C9OGEnOqLyos5qBc2Q1GlkqtEhL
fE6MTjh1w4HEuUVfqAejglqOYZAAQzitgO5ql1pT8tSn51pUwuobOtjG2di61nHs+2T6vwg/ALuO
Ehp4eu0QfgKj5wKyy1Ahs/5ctrJ571+wtsZUMZJCoGJBggyDopbnT3VGYyLk/w5PSUUQf9IA45EZ
Ik2XVG05fNVjrZBSzMNYGdpHdO/GH4LBQlzUPPJITsRnZJahKydCf6IiAJEEwbiQpzXolAVx9x4s
yoB+lXHG9aA8csyd2elzwH6kAPWkP3kiqw9tTAQ1E5if1gQvLLRHweYBJKoKAHcIvFzp/AYfdVbv
BjRA/7m2rY4kVv75cVIEfGzfJ0Rt0RTmG5h6Juyf3aLJPQjA9xN9P0Q2FGg8HmtHdV0fMqEx7u1m
5tNNfVsas67Ubz0v6aIVMGCWyXM85NAmqmHm0lZu+uGoZlTufqSNhzmAv9UZYu0JWpWrkbSA9KWS
wvmRv2jjQlyc2MV9c5ZKHnc6/HZnTdSnuHxOt3FeUoJMK7/8mbYqiHVB44OQ2/Yq0cz/FC9aHABa
BC6Iwz/0/9eX6HaxPA+2xvQLlZroUXtQEweFxh6Ww//trGbZQPnfms5Ir06tw/ALhX47ktxBMEK4
s1jvHSOU19gJqtjGZYG6vkkPso9TRzJxc0rtVpF58da4tIx091nEYBylN4GGLRODFYiryA9gsXLT
3Qmy/txtUweh0n0p5BH7HmyUSAJrsEdDsFUtkF3Rbb1Mu9m2P0ZKWTeKlGSorv0nVqPWeiwCy6f4
qnzxq269Iu4+5UUbGGy7GeRKOgdOx1aTENR5GxmRooKOhxYmFj5E0PQwd6U3Wut7cH1PKZTC2o71
CZfeTXF3Osuw2Nj2LGIR+VGdY0un1/kn35sm7hQbYFtjRpySvltLYBA8LS5RMVOPvtkrElYhFlba
Z3JuoR0k+uqoDiBYij9gzTFxHruU/VgE72PIgFlPe6CIROtB4WSn1YVa67Je93LCw+2HRsrxN9oA
VJXQ/6k4m8cPwPWHSKzA3TQbjkvUBlaCPNOCbESL1ZKCy6xYBRnQaDsKXnzrn7d7AHUM0iRs9XYl
SXqLACCxq/ik7FTpCwzSYSkxFUDDMa6OXms/D+9lu0Clu0ml5i0PpV68zJpS9CJnYlBGActzeBtn
stbaTvkk2PGfIZF9ayMCq7BP8nyl2viGS4uqD5hAw/X1JASwYVqUZrQ9KmgKmJfm/owkT7wMPa8b
ooV8Cc2Bi2je3x68Qee2YhLNjrjH8RYURCOXO/I86XxiuPI5ArLEcOjIi6Z8x+nnREU6rcCoNPqH
HKLBDahXqdIdRSY7+VcL89Tgjslih2TK5dJW33x/ROfnNrM7xyiSp/ULzPAeqTFKVF2WRnbxWeZJ
+qglooHC6+jSHoYYJC7p70naJq/TiTXTdA75B94Dvv18e/t0sG9GheB9VouEOEgfxHkSQ14UYWDx
cpO2C4Ivzz1soeY0Jgb1Xj4ebcocQzIDNasf30K9aC0AWE+ywAhX8u97e/HaYky2DulJ2KMnvkJw
Hz9UE5Xeap1BjBxGGqr2inJjS60IPtwk6Z1IoA2NGTRczbpv9IgHHuYgUaPnWIDbjWi/Mo/HFRzy
5LWfpGdzRqJrFE++NyyIohSAJAE7gdRrfJ0KjYnveVPkxIcaH7SHcynGYJdF3A59yS5qft8Qbikc
hbJK4ca3qPwNJ1Itb8GQezPyqnEpmOVoO8kjsl8QsiEU17ZMDx4FQo3OEDkAYyFrvcJhGmjMoH1b
zzH9jheDVIBa6rwJBWaoNy9YWQsfxDLkRNMzkiQ9naAUPOg7vlVnmUHgtRmyk5Hdq4rk/4piLCrn
yESgmxJJkg7sym1SRhnVIID6+wzS+lVoSTQzdriTgdkjXLxrNO8dZCDIVT8csTlUh6TAzYef1NjD
TDrGacdUGqKm/zP1lYc1XCS94SqwxfmeuskJ+HuvAYYCNN9BIOhuBEtKIQZiVRjnAdgZbCPeyDit
NiI3d7bKpA8zPomr8E+iE7/6GYHyRxF9dpMn8N6U3Z30viJx9gJrry3aO3TvKJJ2sR2Cur+/Xgom
zl4MGVNkK76vAHC7vPbIwULVFeM0nYTbzFIiEQ+azKDqlih49zYGRn23nnMlfnNYNlKM7dNQoKXF
+HgaDoh8tJYqoVTbY07sybmqAjHAcOsHkr+g6bWi3U/aUdKsr1EUWbfiwWPoAqz2t7nQOMY354RN
rv+kYfFewG+9unhonZd2DYLZfAzPU0+Zx+zT3pIGGkRqxNz6RduvOlYOdE/vmo5gPb9XRvtI4eCn
yqpWIGYaZF3WEW4tZW2GzxzGsMEhAyyAjVlJk1KTWQxyVvF/tyAe8tNB6wrw1eA9Vd3A7bBuMz0p
DIiV1nJWwqSfn2VNdvMWVWFDyhelzxzfCSA2RNKjT5R0Z57rxmIEnWgtqrZqnGNRHipNVUbIahXh
ilpD/I98AUmIqZqsJRwTyBDkNd2UKMBY5MU8J0a3v79QQZ+2FRv5PlFOhVyxjcXCqRiqoBZZ4q00
wCGbkIGNIDpgVyOjYQOWqouan1qo0iEf7bGgDR0KEHZCnt2ZbOChUJcfS4f25W6aDoiLO3fhJB+r
boco1y4/9lEHUWIGZxd5SUbAz/m59boKKYwN4WY581QsawezuCvOqk+AaVVH8jcwLZB8CPhTg0DZ
7P/nH3jW6fdqZUYD3WUhCGx38eGL4qmLCGr+Vb+aRpxurVTfqr5p9UeuxU+CsviROZYgsq938zQ1
pxZVEfGIWthxLwqKAJRqFWtj2yOpyHYOtPCly4XFl9NSZN6fYKnxzl7OX3cm59cqN7R3VoCp2m8S
fJ40KTebP2+1yVFNyPsmAeM87z511oc6sVvkBDIUZ1QBOZJZbN9qAbRf9yAOuzo0h5VnRvOU8yJ0
n4jdTgw7t54l1M/zHyQvcg6qxQ9TurF7eyWs5bGQY98BnULjrFNsKytzSvlspRaH7NVWaUOfk1ZA
s5mIXebH/s5QmnBVb7W7Pi80uk08nNDUHGaWcoWKcELddercA1txdS105tP24zilXjYEaphYocqd
aKPQVORF8c/v3xcJhw971FxSYR0iZJjGSe+p3lAs1XGUYKpaUNqK8SbcU84l7L3w8GqQWeJrjqM1
81sDGDdByHxgpNob11SgHhTxshKiWa4ScmCw+5PzMr9t8AsQpYR0NFyHjFP1aVNdxmDCRBsEce1v
sVjrsvgQQytkDWI0ncnSfOlSJLBm83cy3AR+xVq0nC9g84DTv7CZ9sQUBzN+ACFQXUhORcTgu/BU
bjvyPPPSOvx1U7dh2Yd2UYo418VZepnCoyLGoU/Zy7k0tBgGj0T85TMh4WkDFRzFBJaC2SsjhcdU
DA7tzmVbYOG7PxiwtpC3VDJeAIAoDeAaoAnc9vKA3xACPyoUgqDNGdJyg5cQYwXgp+Q3WQ4FBwtY
QA6Sz9qCWK10WnFmbCHO+b+csbzLcgNQQfd6v+rVYnClLmMG7x+YXzQtaRQOjLbvqDNX5o0eX2gI
smx7hjwej3A6+SAPYz2G2dqGqroGXM+MdQA4UXbZFhhSXkT25tJ+s6HO5TPW10FKkgsankJlkkAI
DkXQIWo6mea6mebOoXETperqGdtldYbtcdv7ToOWSsqRA+SwNBgWUD86OKcCJUhf4NfI+ErQ6BqQ
Ak2RrFMfb/QM8dDW+w6Uez+ODHTiQ8zkVPnsrzwGksnDYN1RlzpY64nxpmxkRW0Xx5zUW5y6nSXj
/2DkpJ6vpWuiErMhufmk+44Gztpzqw5ov+t8VH0NKh2pDbJPRvrUgrW7i7OcX82A6D7R5MH2KszW
R2fLEm0AY0WxpA2VHMrtQ0CXuhqIBujZmfkBDcwNZn7qx3UsLgohwGacx6KqYVAfLgvXib1+anDO
eovNXt+eb3r/jjdBgbCHSu9I+G9H+HaZUE6rgBnQw7EoeNJpHwlj09b8XY0LvMmyARflvQq8u9ZR
MMR1djP2KnMnVnMTsCVHDCj8PhNcM/px6Y0bq+Tv+AahJH16iiQQ1zefxOsJnpBFQBfQjSMZQIs3
xH5yBxo3yZt/hfdMHcQAhwyEKvuF1wHti0cy7gZNGdQPMR1H2ZXqoN9Md/NcgTvFbRUCz2Y8Zj6x
kpm5ntxyXxrbUyH+9QBeVKCuV0OR2a9WVNunRr6Dep9P7vRDeGBAYUC8IQB4Xas34q6BvyPE5T7l
HPwdVX4Dqjv1Zx/nTta3ZfuBlsq1H/TWd9MtwsXXDfrjywYGE1fReax7IutZA7P70+yb0L74rL8B
h2se0XGNq2iDAeGC45RaNoFQY8KHM6RatF3W8MqxDdBYc4hXYplDmjLLThpzs0fJOtRu1jQ49569
rBC/AwPyqZsrDMdMg+bespWpLpYYPmlIfaAsYvKGfNpCwyT55LRUA0baOxWTsPVuXMsrm2j5MVu8
ykiKag6DZ228TO/ir7I9o48ceOTfr2Ia1WkkfJi7yHcR7fWBbGGiBRcIXB8HMgNNHJkzefJJ8Uyi
3fty6cD1nMgcyN462C+tlVYuIfiC8Xz9fVj0M1E6jF487gWA1y0f5gOfq0SjdHuBS/lBdbzF5En7
NQgrdgi+R0r5ObH45o6nzbE5uA6Nb0EhpjgLFxnfCBlWBlf4FPhPCmiY5P+KPvSwnvq9S4604drq
/L8zDiP3Sr1vTQb7o7b4BUVcJuTw++nk4qE0PmmFXUzmXG0zAXo8RcR4khf5q5CTgzzF5pQ2glMz
FfWK+7IJYs71kUdHIkYTDwFwSruSo55nFsfm20cH3ETCmv1+OIToHsbg1ciMh39HfSPKXuuvXGDF
/DZPcfvAX1Y8yyaHJDqjGIIY98445fk/goFf6l01po9LDvyykQWVN/sLyaD6am/5EirK6REch4fD
O3PK0Hwk7adBakDr0htzj6r2D8cTi0pXWtjEoYNb0FdxhDo9LK5AR1d1uju0VIParEd80U9+nIXX
yvqinazMgv1ykNxRBEAXR1+hUMR1EEYkNzZw1/2+njhI4fUrZ29ZKpXQXTyrz4Ln7PskDFdto/Gj
syrHQI40ZUVEMwnUQOeNJ4GQHl63/owxCLMVIMNrQQ1gUEa7I17S8LxRevGEyHIXQxQIh+PxLf9s
EecpeHD9kcCYg+5Zkmv7CpGgs3aiIsrUnmT+8B7/OOeKHqw6qvXBjahCLiAbuXJ4GBs3EwoQMMnK
fOo+DoVtFgW9KTc5lU1XHbazt5Zy07ehKr1sIbbHPFw07bcoWmI/VCJmsgzMPrmNrzwuLfQgcyTa
9eACBnib7FHHpUvmn4+D+YiT+z68h1T4uSSwukg3MRrFzxInxT0xUZfG9MGb107B+kfNUwRNMvnA
z0Lhpn3eKK+7j9bUjGIfTNwWrIdzZzz/69f6luJDDlZGrSO0hPtDuTs2QsNVTT8n3roR59ZC8SIl
5snrf2R6kbfRq4kGAg6o0U1VIP+Li4nlu/Gzi6Z0TFQeA2PNi4PFHy2vNWj9l6qZSBje995osg1C
O9EIoLTjy3fIQZHT9iQu+uiWRDBaB00JtjloBIQET+sU25Ni4cV6BWImuxY387VcbF8sUoLubEN6
uJWgq3ly4S6LQBllzveC3FQfmy8ubqUWOZFIZJAG3flfWv7wts3KyudtmtGUyF0dBfw5JUlMbYfF
N3g6kmLneBnCRxKJQxpOFqoBWUcSH71aYMlMNTmywfG/ppaW+RsVbtNhJXxP1gm72NOKMkFNpnyu
2z/3Lo5xDuP9kLH2qn58ZTDiCZy+xy8wqJEfjbwNKCXOR4wb1a+26e6gTwK4UsIOzRNYnhEefD5+
YFAZ8dUl3nhiutGbv9sB2dLtjHtWNWga7/fJb3Qgn9NAiVZ/23a4pDZ/PbnYoBM5S5MJIkE4MsoX
QeSM5nXgzbYUN7vviRovG0izgeO+nF5Cz6fb96rsUNbNON0DWycFL1HmoJO13ZpL+fYXR1PHTuxS
YQGRaDuEAQpscaFzPisUFvTxp4AzCjtsojQQNRrBrzh1XsFOb2A7v6HZq0pM9R+MRjuwvOqq8TqT
qZJJlfvRdTqchz1CH3YS+iupxNRfzPASR+rMvTpJpN1GlKG86Wy46xooyV4r5DY69YsRdJH/oxGH
LiHKYmMsiJDnk6wyenzK6r15dDQwwt51Ei0N0M3w7Y4SbYVEhIDGbsVrbBkU9fzKTX6g0OPf3AZB
yWZNZ+dtqUAzqJCLO3/kKUIHMvXuJKwt0Olk/IhnQb57KFLIAuZYZPjfZM+1WgaR01v1q9MoWhth
jlJfppOB2VodkuoZNkinliDzR9t2KFJclcadN6jyhdyKRx3G9vl7XnURScMFDesQlS6z047SqvWR
9cKHBcuhP7MpfKQCqV/tnnfXaLMo4iAlt98c/XY9Exaa25t3QQHWHWfkRALHbnTm9IN9TbeuwTbV
IuHgGtD5TOvWbIToIk4YfZUUFGu6H5vf6HGhoe3rOd8sWGsqcTBkfmgzW8z/v78S10t7sGu1whA1
aM5BQjGcA+Le+mZeaYEC1x34FDTIBfarpcTPqcp+v7sj1I4AXNM2LNXP6wmmY67Q7urFcf0mjeFZ
qPCWs27jnnm+nicQIYiIl5GBkXxVuENXeBFATjRAgBhMRA/JS9Ufzb9uW1/00e0ubssxay5T/7N4
pwyc6KdE8V7UAX5HoRoNSxG1mzFU3nv2GJ2clTBjA3U+2FHrnzao7Q/U77ifI/fMVpKFVmAjN7Wo
fwRJxvzyQXSAJ2+1gaACj8jNXwlEweYF3r55Ku3hJV+r9JdRfUvrXJbURY63fqtY2mpt8V9pR4bp
FAx7gm5cDt4mamKV8EEovctXwZsFT1hKrBPSNqhQIZ7zKUPQ94NErZgStJivLyJJqhFWBxMA1L7V
NLMrfL20fV9kPzEULhI93iKQUHxwTOB7L7M1+y0cIwv7ts4wiryE4RcfLr4J79/ZqG9JvyHhOY9I
FoygTq5WI/bq4pMVV+aOb8bZ0SZDa8yeZ+wxEYR84MVDfGmCRRdN3kEgsJpH0IHaIO1aFNXQJpER
FaV/8FkriBoLThmyUhi2kEPCI3V2t1v43fuxr97Otn3jlyl3FZ7YKZ7OKuno5LVh6a7IK0N8kUAY
Kgw63P1CUoWvJyQhB5vYRcGqtIvFdQUITfXv5Ulp0xfqvv/9Sl01AJ3Pf6ZgvidnAbBg6gkzNSjp
ZVK4bgoEX7H6ZtUV85/9VJC2JP/74Y8QikBU24gu2D22bI6+KIWNe2Z+nxtlsDbITXtyPDgxBkOW
UbzPwOAq2HjANhqbwPRz5HyeLvm/1bvNpgn/W5AxH0tMn2pxcf/DS5hR+I1p+arHzXeDQ+Fp+kqw
UDczihZG0ARI6w1CjQa6SfGiISIN39JCefc44we5Xo0JtKwM1Mf1KbmCynjvdQTJpZRY0Jz84t4d
bAckkqBaxatI8WiEv3gFGfT7naTrczl4oh0z/agpvdpbHIk/jF8hvJEhnb2EfT2HKc6mFNYNto9t
4Qp0U5SzUhRhKFUegzxMiQ/4y9etWcdYR4UBnauypwbLLU9CZ5w09/cJl97PMWML7PAmwprSfKA6
5cjhX0wYVaEBz0o43cuyRRYMJAxnqf5FelXDuUCbRWAkV4yeoCWn2RjgzvGvesIn+SlMsVjSD3D0
n93higpTZRluJSncvOvqWkC6h5d5kUrFWbNZq/qVaxdGesWXSd/ihUSqsnr3oVFiaWzM3iJavDY5
RWaz/TvQ72T5psc4u+ZcmPySE8AdqxEbNfZl2artEon+EPSAKEIcHbRZhs7tHgCWRRgv1is35gI4
AYfcE+QZAxMCUhmMTL3yXz6AU8AGxrHXE0Kpi0t2QBKlrOXwIP6kfSc9Rp7Rg2AZy8bDqlLYxDDP
jLAt1ZqPYrmdHza10rTH4UazSu5FvAoOrsvSg53S3CHptaVaYgcZM1avujDM9gkFM575fjyTk16z
uVNSeRFBjd+2/E6eyXlKIY3aNMHGDBgrf5m11syAU/hnDyNBy/rkZImbA4NB3yktdjRRYNVuidcR
GIqmtyRpp7QYVI9/qsv0QTbem18OsJJJmC2ESSatzEwb/AKrOa/7bqOEd6oAU6wa/4wninA+1sxO
3f54PvjBN3k4KdOjaPtYjDjMPzFSqYlFLUdLMyX5jnwxrP6Wz7x1LqAjJpp4lzD/rUKtY9/ttMna
GstIKIgiHVemo2nB4sm0+OQ1RhdvQz/yGsnnXia7bbora7umQmMmRXv57Mq7EJ9lLhxxzXILVMqs
DBm63FZ/acW0z5rQF3VMUBayg9Cr2RN8/COTdxVl7q29LdPgopewTiqBo2gwy+9AAlYfOyhElomA
Qkn+5FBWNp2V02FIPqw8R7+dSxj/dAB977mJ9cJ86y8qNtO6YuBikC+whdGZQ+Wd+IJuoFAo2MJK
lgfL2NC358pzRYFmF9ZtsMRQ2VUOhEn6G0rCpF7Djq+pHT483czvHZAz2OcUDAcve5u13ApyOxQR
g4iYQaPc1LxIa7SUm6AaYW4R5BY5O6Kw9vJ+tSS2sJmNy/OQUox3ToXBN3qLpmjyCwZuVgV2bBuA
i6/SQ4zwW+BnOb+PgD7u9Q6XQVVBZpx6IFILXQAUGrWWPVPPkLXCZGU1h3xjIWP9DbzFK4qICJUY
UoMVDDy/MZCdZ9SKoD8q8AGVlbALwamSSvwvt2WLSjqwqh+zjZFoZy4lrhziCp4Lap2LlOlcRVjl
I6ixJZg3q3VXhmz5Hy7Hidd5oZd2NgubNFujTh0RfuGOLiwMdjHn1aieXSYnbBQcIWSJduIkCqRE
N/4NMQ/Nnz50AQv6xhjNXHSKucZTnEk80+4PaztWvYmM3/USkrwb288L1OBS+jbph3BtcpER/rsu
amN/rAp2XsBp8yyT7sUM+MQUYpbs4o9uM7CKchJVr492iVJrV692dNyp/GxvTnxuNOu4wHr08Xsv
YLnBevX1H5tVNCZaml1nds7KXx0E6ZfEJSP2NR2U1uCwlznjw9UvEmywcWnhgTTcE041hF2djqjQ
zoRpTW4iH3VTruIveGtjn7+FnfAEdHmakfpvHwEzJ4sFEhT1Gxyk6ebgMyYeU/ATbKulehrAYa5V
sLubG32D5fjg76YMcf6sTunopUF7NsPprjysPy+JsKhWS/TMQuN8b6C+9BrZydrpkKnp+5APop1u
iU4dKK8lj9szRfZzYNTIDs0+4aW+kQ3auOqaeWi0LuMF9K5+dAtejCNGiqVARFMnPbgW53Zl8lz9
wULz7xGNOsSxm+4iQ8Os9+xRyhoXctcgemGhuSwz8bONpAwlno1Ii7FgOt1FWlxJ6vNYfdOk6eEp
m+TGJrfb1Z1QHXuM9fd5EFczlLoP6EJZNRHFx3BLYxtWQNiTWU13CATDVuLi4q+B4Pigbu+w22aQ
zwSaKXy+2bxjSJcoM553YiPIV1Opr/Tgg4o75ckYMaSyMFb3eHmYYpbPn5qPNT9HhRbPxgTIBsc8
DfT6BvdVCxnaf30Hnfn/rerBYDe61ZfumGjUFo8+y81YbOgcuUiE93fIOzCv7Mi0vQ+8MgyFOG+s
v5NVTIyGaIICC/ckjGRH56faSirCa/gU+2PE6HaiZX80Z0NfU6T0xy2GgPs9x/Ap0fLRNG+Ufuj7
JKppLms9BM5ZfG+FG9E7dysoiM/w24OkCJvx+v8HwjSJwCikhKYvZGifCfx5X2Cy1G4IOplHYXtk
2Z3qqAlu2gNYcdMtIoGBnpM/wuLYG7qJ4FBL+2hTZ1tT5M5NAOVqgCobuDpLsnvrKfjxtjW+C/80
BHK5s7RWe054q2fXHE2jGxdrruZFPbOfUo/WCXt/Ky9PGqPILvCKFNIEUhZCjPVWLBTuM+gRInXZ
IH5Lvn95UvoJsYg8UIw3hhDczC+4ub1GVGAkGNDEd9/pQHNGb+H3T+x6/fHxeA35Po99z/8oDpO3
KJbkT63ga6DLETCbiYSbGs5V8JsFk19ZQkmwWaSAkphCmYSh69qvl2y4kESXK73iB3lbzIZJtIUN
cLn8ShytA/NmKOS+xj32Qerr/7Hwxbv+pfPZ3lWxF0F94CFyMlw+1nyuNUCCwEgEuQe/ORC56XpN
REpckb6HtnA4C+dPESIwotV6YIAr23GiadiBszFixmfC9RWvJx6iEZrR6zVC7n/Jxj9wctn5vL4M
IuX/eRbOkPsIhuqxidjhcQA7JMaFSs+0d6Pd+npDEG1NgDe53wQq97xYquQYMj/irvwQP0wpF2ao
ph1gtsnlukgVII1m4VsIvV9VHHZFBUrWASaiicA2pAgGmgNT6JT06yjUtX/h2F0zhNvh9v++y6iu
1J3z7Srdi0JhfIzOF61odsw/t9ItxfDbTOKPeOFLzNgsglGcZhX9VrjSKi/Nvnd4er/q1B9IcuMd
+dAQpWQrTfMdOzaoKT4VnlzaxfHZru6S0Xd50HbMkKF895SZTp+U6TrNkrH58dKU3EMAZ4JHWimM
7H16JoVclEiVfjMsXBoLgEd2o6usjrJpcASoOdXGJt6fPpkCSGe1YtzM65/dF570pQa/L6flBkks
wgS9T1FZc+/j+61qLjpfsD9vjfRUG/eswgh/78uhDVfkJsUOeUhpqLI0PTtvg8e3QbZ6PgVUk1i9
+O+cLLjzxqYVBoqX6Y1KksP9E0ut5kISYIKBEiYlysmZRrqqH3hKF3uzVumaFjIXeUiFCeFTbW9X
sQgvzKYeyvnO89UNZA2OumiL/z/5M0XDqqAXqLIcAZ0s7v3wF/88a8oIHQT0hRUoT3WNYo5HyisJ
F/MbGr2Cy+qzu4aBnj3SD+y31MN/GsrTgyRUlvXzMh6EDIvevtMjNJfIQ1zh80lnV1VjtudjVhE2
BkMNNWG/qYfDYg1CZbX5wCO0cM4jlyObFkwDYUxf60Nyh+i4rlLiITF16abqZk8lFb2NxSmEGNu1
4XvA6lYqfHcqahQH8Z+0xlYnT4mnd2vrPUYRUEfOmAAFGHiiaYASpGmL5okQs/Db3jYhgm3fjTpE
Cgzf7+EoWZZZR1P8/+6+NAvgPJK1GnYiiLw2Za5LB9pDsV8QttdFHN2cZvHobBmr4+j1Ba/QJo5z
c69R6I+3NonAwpRgoMr4UgKOKLdwPZugmSHV2ihjt3w6uZcfQLbCwis8fg26qSDAuOAKIzcGybuw
jfUn4uX25n0P/MlpdTHGM40CZAoKGPqgmfrMyFrR5WHP15Tln1lXzACIMCcaLcr9JJQtZ4aSFRu1
yP0mMT1X9tPe9n4uhNBkC6+Rsmy0dd6AS9q/vYGD5+480Ctx8pV+RMRSsz9SX3rL0XqvB71vReVK
YQ0vcTTwk8lH89uIxyP02XN9SDAEtcRdzVihkxzSmWoymRR/x+kFFSpICNFxh92zbGxurkkZ0loe
nazauc31R1J3B/kvmwJEfYgt4RWiSrZOiU4YS6Nv7iFrF+o1ah7sJKAMtFk0r2f03WBRZmF+so2z
CbqXONyuC2eJUOl/ERLVD28MkyFZuF6cJhanEq9qYMpczrgnu0U3qPhFeGSR31P1tRIlCnbVDWrn
bwBQo9KMWS8Unwf8K8VD1DZX62781qnZBJvwy9HA1IDM+1DYNglFEHJx3hNC2asmrodY59FU/oZq
0IMfQrc3JstihETE69yh6c1PxKj9EJNyapweUU1VGn7yniMWseolzfVMOcvV+e/tlllueVLAsgf2
FQUdqndweX9T642+dxxum8iqSxWNzeHrYT76TZnGFT+9n/rUE5WNT9XGcFlBjf1iBsn/nl3ZaxEo
9AfcX9uxjWujIfvgg8IVREDSnEx5dMZ9z0fFfAsHJ/EDuch2kYZmuZN9awZ/e4MZQLzqdqOPhMYJ
xZuGMh4s7sLFKv4VxjrYMkITEYynN7yj+4auRmr2FUzEt/ITkeyivHLq6IhhEl14SPbKl9Uuw2p1
fk1osu3vf3F7ebijguB1uHho1Bov32ae8XkAO/OLtvQgn3/tuE4bSBVZ3Zx9Adh6RBt2QvW0m8o0
hA92XtKWB04kVi0jTahaICW8nSJoLf+MvOHQhdEhdKv+0us/IIfv9KIkZbNLcKFmy6XXPYns9qK0
07EIkOO/hJJHb737qIXeg360Ictcg3ByB7zJWJOGIMGPMJ5mY382Sj3NeqEZvQEOAY7VW44njXpr
1ytmYzSJ2+oZ6DHP9dEqhAqfmunuWf4IcRk++PRI2TlbgCJDB0W9cmlVC9CQLXYAIGmz6U4FgwIG
XEjs7pggECvnCPc2R6tPbx1yfZEoRbft7d1FKZN+HLg/r/GyN6xNtmWGM0wQoqqPIo/g9ctEw9ip
QgnVYqfCMKZKnfGtQl77sGOY2rEmizzxHAMplQ162H7fq9Dc4E/8iW5Qd8GX8+JQBC3xmytJ862C
f66JvzDMQUgWoQGhVVSVb/VYFXBHVELpBV/wDsIDe4jjuAdtTdf61+ebvxwBJOM4P3hllMwqIrvf
sAQFVRbgzZIjoGepylJd4aRzlVRkG8E0N/EbeAwXnMHkFHjo8gyLm9fAE7JyAGQu4QEzvj1+dHRf
tyA8yjZFOyO1EptIOecmgDHrEzfpgUYwqEvWgMJlOpO+Wbu0QPm3zJBC6Z6kHkZRXU3vAzrC7Gwj
OXF8iEBFsVsj40I8q05wJISovpFXtTgLQM/sGYearYzi1UHhsNPrHRh0+817FycDUMT4c1lHHTFg
1L7LqjmRSt+vpR8M/+mo2sfWcWrKuBZ/4qnGcnSWpXS0nln+od2Q2aHraDx8Ax4MWt3Uf8W3bP1p
PT+IlXXpEm8MGw6isuwxivPXRYMzQgoCtswatiDTBw184I5+b3JOpWf7AHfYmxvbWtyLarAsUzqR
8oxcf/dsQR87e2RSJy9aO7d2UOlY9BozvtEeq5KpXAxrKL7m8jYUDgodIkh5ABg/OivNN/x4v8kJ
iB4MbUjQrMlx6Q1hZR5uugAhRPddvo6OTJoIYC/acKn4bGLKfAH6yJ+xoo070nyzix8h+MAURqFC
yMD9dAxre4CesC24+knXHUm4nGrN5iLMUHZu5Vyh3YNLggpeS+BglfpfM4i4gPEUx9k6SuXZAenY
lIWyVBUPBc9HzP/J9YiKfCzqcc9YIDVJyLaHRemRzA5Monnv7R+AfVwIzr29nKttdM25mNBmFFDA
EZPYskOzEcWrx6dUz6SxMhGyMufa7bs7qxsIoizWZDhJroRR2/6FQyhAZx5J/H2Drsz033//JNss
klT6RSQeHxFTX8CyShWkGD78oaFr2JTR19Kk02k63Yx6yv9Ltmu/EBoNfLYFD2R+bQ/hIu93rw/Y
IvCFurxRrjYxc6ueoZzQWS2jt/UwN+YvAz8Z/bURcRfxvzauYauhOQ9jcoPQQqU2VbZEwSZ0mXtu
L/scIxPGP9A6qPLqRlvKm224Ogu5YhgMUHopGbSiPx6el5hCdP7WJUvWwI+Pyz+LTw2qg5BqJjMT
wJxJ+VtbakFTjdd4EYFP4GF7NpcQKMjfJL1FuMPhC7OkVB8h9/4HScN/1f5c9lDPArF+bHw0tq0c
7skO1vL2pU+yQDbHoB39k8gTbRN2RRtGtXk3HZNk3jssLUBkmqBI6roQQ1CuABl3gvEOsoEViK7t
LtVZWuRldkaYhxmpe4q00r55PknOWHsIBXg3bXz7Et9I84EAtA8ALUVKhuZ2CHTILSGhlBqBrNa9
SQOyVIxyVLI58HuFdC0iGkZSp8MnBJ7rG9YR5/ZtfG4fuPoOymKYRuTA35Mr+7UtBc7Yb6wqOASu
22zLI3d3/EMimVBaue5aS5Gb0AXeotS+4BuV7zL6naguOm6x5i2eqsiAujj2TzrbnEH/1Qw8JC44
JgIT02EC/tDX5U729HEEO1BCzbz614KLWwjpnffWmLScB+T90J/rbA66auzBOY9LAH+8MaO5DETQ
AMjBJM8bI/uWcHgAeV2HxmmeKBqYNyWmIsVqRIQJAAlZN/XNEJ3Be6vJqbH/hS2eEGoffnZhzdLe
1ffcf7sWHjGTuHN3vSAVeuDTJhriBviFEXK32VjFlu9QklnfbwGzkdTwfqfTc98K+JYDN+Ck/m88
uFa+oIPFBn2T1nYcCTMtsalTn7fvQ9E+o1BP6fAi4KN9673rC22n4SVvwLlkTntIh/PyhKruTPyF
n953QyMjfVwi+3geAfb4TkZbYFa7A+QPWQNGCrtiIzmAdFyYnauYCNHNQP4LfrhMaNLZ9+4xDflp
bMtf3WNzdn7abTYW6G4MLvXnklkFevChcbEUUJJ3yzUXe2Ue8T0+1j0tT+2pEGAqwxhF8cc1b/y7
Xo9P7NWNiF9VWCnmWr0XDNeYSW4HNiwIrIlRHbVzqkwXAvDk13M0QExHeARYnqc2jXJFiEYdaF6h
M7nmQRLxxrFX2ZlzW06B1l3TjoK6FnYzaAuq1pf5N0g9IPUQ8fIleOXyqEbBldv9GiJMHaJywwca
Jcfeam60TcwqaiSH0PkaMJtEFZfx7IrvfPBrdLoewXWAjtvvN7TFuBi6MB85BTwv8EU1kOYOy+IK
Y3dl7tVo+wJgRogYZAmClOy0JAbT9NubIGWCn3qS1BiAM1jW7bZOyZI2oXgVn7jXQXNe6lZDkTjR
+j/C6UPrGBWtYxT6ntpDYqy4e4V9ks05hKwtNWozE12yKZAM+j+fmzDV3TV0FfVF3S6U7Mkg932Q
tDcJ5NiCyrScsBCRl4pQYiYyoYOJjU282WRBdUg6/tKtMvuQ4tyk85z4WwR1aHKF+kQgO6wsd65R
cmvEL7NrUGiVWTkrhhFW0EoPBRhbeFWOhLwbgXSeLjbtE+IicnL/GVjkghgFI4kuKTjPC3yxjbTc
o9aZD8gui1g41NegTA8PRJx/iZeTChMypunAD4eJFHhm4+Gi1b9b7rWk1DoKWRee/m15I5zTHLFt
MixduTzhtfjXexf9eNQAzPtDefjrkXzY9yFnJiAgqDmHDETLOH2Ko9udjQRBVkCZt3z9PU/+k6//
oeL5Qf8HP+nUE1srpRKZXx3dOhTRmDbHlaSgcxsZ2kEDXHnJdstyJHtvho6CiqaFCVjGW448HJKL
2I9sq5H4/ltlkzKpqyUP6vO6DYMQZZpuvsxjcRECe7YGsZJOwQWz42dhDrVdP7lIpb7WJPapbBMq
TzZ5fGHnAiS6zaedzOeUj17Rr+QL0OOPRZp32BJcB/vj52en5anCozy2BnhhC//p9McjA3QbLOGn
hvVivvgCGgsJ0YFM9j6mDTwcr6K67NM4qaMsxf+1NH5Z7Pj67UtQmKDmn3zzZ0nBUO9OofaVnEG3
309VvhVvknHRQDcX8N3Nb2bKMTeEp27Jj9zlXjRZpjH8hpBcj2/hfeRhWHbQgiDKJrX/H8tB+Kbv
Wij5IqRQEro2aeIW9wF1j5yLNUAcEufvuu+0D/DT/ERCsxRaNYpSEGB+oyVVANbf0iB5Qq+/6U8o
eOYT2ASpzZag8swjjnxVUY/aQohEZEVpq9RebleJ+PKjnpQ6866q4t5XgXgvI1QXqrnLUeSMiNvy
PIY0PF1Uz5fQVGQPEE2Cb8uJ5o35HG0WEogm4aHxXdrUeI4R61QAp3qlrdYjDquBDmFTrjf37/CI
g7+X6Ha/OGodw7u7B5Io0opBoJZpJkDgbjBNNlSbGsQK4YFSw8A5QJWSZ6HKBKlwygz4rnOqNP3W
iaYxozqYyy4zKuiBT1yTSYDILyHC4/hUOdsQW1z3rinqL1BbWakFpcZ885CdergXZjCCabD1se5I
rUm7PhC7dueqfmwLMKtfQbJUhlqfCDelOcjtCZ6LVrfJ6GTyaI7iIRzBAm1rpca5bKfUTGq73HYm
0sxJcqjMIWmJBLrVg0axJxBZU5ZfPMYKIKOjKHvRl5z90CO5Xn8OAZ7JzP0cG5i2Em77qNRiwiSl
EQs6XYN9EHCyn5Ir1qsG2ggrvYKPasEyyKq6Y1H8v/VO/x+xVaRqkFvayLUvH7G5COrhWVDndipo
WA8QKXF/n2TzQXT0fljbm9a0nLGjCVVAb86ktoP8fHbdB7FvADejjtIXdK342xcpABRFdAFXPtbF
stgCBg4R3zoQpPaL/s/Wy2RtclrZmlpFpxqATm9nGGMHNtskrqlEQR8J5tuL7sgQxa9uLA6znZLW
/3aDnoAcn+u3bVKxt8akX7h88fI1Aa18x8yvVAe4WPaCmxb7RKAbRto+CBiCtyB0QTCfjJSGR7/g
efzj5PlgH79Tfmpi/Cu85bOSBQ5CVMTTN0PVA9eVdTyV+fchsOy5XjuFG76LZklNifqT2DfKE6uu
Lh1THR0lUVfcu7HJ1ICX+Q2bH8VtbvqofU5Gz9hGuHgtMdU3vir7C5O+OlNbv0/mYBViYl5UC2w9
QNAwbKVzTc9ZI+vQQpvdr7t9p2IPm1YEkM57qpfcHa+l8tSfHZ3ZULbT9BZT6Bxcab8iqjERtgNO
HijByil3L2rKaNKovB3VIJ0dPvQQH/zUnzTLFAH+febb5td+3OoxQX2cFJk1M5xues2kxVMRgeGk
Vhf09VBtywUc0Jcik/qkMZNgMK/HT4tnTcarpKzrUJwraTJCYZswBS4FV+uvUR/5B4+O7HzbWQTI
/6YqXAXpX+H10CF17nBcQUIuLKdWgaEenCbvQZfK6qVZsOQrOgXbvxiZaTLV6QNrxR+eGharSwIF
CzCvqA0YZyQMROflhED1Ey4IGZanEx4bu92MbfWi7ZhOCrg0G4f1HbYAMt3Ny3HSElbcx3K7FQFU
vbgQFq5C8greID/hN2KHVpuN61qwYUE5lCBgMY+HbMKmEO6PbN2z4PlA+/bByG6rQeJoP3xaUJvV
w5wYVxXOipKrkcsQjJ7o/xbc5/Sn5RiEE7C5UhI+a5KZOPDJLvTg/h0H48sJB46tyy0jkmBHl3Uv
zM/EZ97WwLqwEr/oYkCgwPuY5gBo5+wgnOUqGKaM5VgjyD7Q7Up9vFDYTjNI+77e8Fwl01kYa0FI
e6dbaZWXUijsNlCDdrWUBnGSvft1bQD44rONiiI3U92fEN7n7ldpQlR2kOAfAWhgwCPPInX5J9Sv
roYDyT7VFXwMNohcTFtItGMDOWVAi+T4ncSU+gsgdO/Y2Y/9qTn4NYK3EUj8Uzo33nP3CNsmcYuC
bONgWOH+HKZCj7Zo5BKTDzmNSiJ89flnpay9e8EqYlUPNNSyiXSv0W/LduLRL2iHDuQkVAytMYL1
D70i9RTTq1VtrO5tv3tLRSDK0wl1i5bGN8OfGJvQ+wp9qDmrkZJK6hak80+xlZ5x0uhLhNmw3dWM
uWDNTT9mqwxgQ+abCY4yYUXHwPhY9B+IU2Ots/grPR2ON8BEnmrfiPIXqLuwKZhZi/07mCybnUrM
HtCNLL8DbEOYLQfaRAhtJrIeiiXkrYL5J+2VA4slYv0qpi+G6zVrDpQW9UVpQHzKlrBIvguIA1rr
j5zWG8PcFTJKvyLsNA4yG44yJp1CJyO3e65dEv4xnVPhf3ab1qktTKJdz3/vAwfvWXswDVKLtuaC
T2yzrmBPquKL3jL6Fu8MFwvNEtB4s/GzpFGUObrzLy2mDcv7HM9SKD/bVUXkbvzqNGNcBEEDJNws
y457u/EIu8t/r7yXJWuD+LsdrHOHbTZSWg8cXBYqm70RkcNiMFlCfrGOLkGA3QseChyQfOLr7ruy
Ja11i4lLjJA5vuozHiBQFsyvfzr9DxxXkggbohXjBVnM1D1HM3moX8vPUBI4Ypyg1dhigYjRNoHu
8uGM63DykdrGM6z7SmvzBile3d9f5biOamMtD4Q4lZ2c0/sn9SKXP3zNhYPWZVLBSUk8a16e0Yb2
CufJAjw18T3D8EF51J97UCtEchh/d4W5a82M908rIVNvsoSGHSpdymn+BM9SDvhOD+u2mPBfRHQz
vmQqEBJ68G3yY0QiP4J3ARmAk8gm3YDiTqOhxBa/m5PqxB4Y3pI08/RObyLO+LHc/+iARWAzYofu
nByt6AdvEZl5YFB4JCy4sXxwYXKKqufe8JzXlZO6v3+sab914P2YJ14a8SfBXERIcwOysRTTW4Ki
xTeOQ7zBFNtuw6w9lBtXtGhrV4HlIJh9puJviXIZEhont9HSKd308G8c7q1jCHw+UA8NEMsHUjJd
lssqtNwBclx5+8Z66MpQl6Rf2a2Odw6d1sWaxq9PMNs16YyUZm82ZLrwGko+928HV2Z4o74QSxVC
pqfYI/TsZBdVQdJ9QOMPt1kjUx8ZQVSsefX4ExnO2giXrNxrf7qN7px/31IFH1jrd+MEE5MTSoaf
VPmYfZeGRxYGsKHXNiSzq1VNZDCid0ZMNw0ApECokZkRacA52z88h6gXqBIPf2hfup4PSlefe8BJ
dKMoRlhMnzgQBlRelrqlH2NmyMRFIEIS1WXcq2ZWONQYa7ffRLFx1u4mVnLBvMh/QotijO1xIdj9
W5LHSbnI2elnL918tN5JEVGWUqMrodOyqHKlBivkWZyH29RBskTRa6o29glxTDxBoLta7lr9UAHs
K0h+xY12bOg21AvjEzs2R4sjp8TOkrCp0rEGeP/TU4vZalIet1qWtbzTqkYu7RtmOmr7yLG82W5F
IiFYUENYagAG+yQu1qBmrnsqbDflK/uWXtOLJ+09rwxNi5UK/3lzvnmx0LIY1g2tPoUc+lgxAtud
GLUVAMDKVjxH7z9KwB/grgGP4obhsMD8vb/PXGbADRhsw1FkxBxLwZ2Lh7qzoEf675Wo+2Lgh4VB
JCGbiZjuwocbzft2Yig4AgsxDuNmu8xXj1sO5Fc/IWiV7Xs5nQWGByVkw+8VBiGU08H+pmtAAl+E
bWxhfiBn8p3kOoDnyf7oQAiCgTDCMCxEO+nVIjCOMkTg5Dt2aE+Nufz0n/MgYDBYt9+8RRhTa2E4
LwQRVLCffYhpyr3KCUL3g4pYkpz/n6hNWFHDkeKYyh7s/DMrPC9jQ4TNS/xpaolLU/ZRRobFb3QW
P60wmHc8Kr1pM9Q5fYxk0o+/x6h5EnjblCi7dM4vAa31qpjpqo1AVMXNergpXe4jcFCWJLmJmgCo
SqIPHSDVUyTLD1mvUPHIcOAFiBzD/OcvzA5q6KITPBngjOZ5Zay5vNAv13oSX1zvPf3Z3xEVgIfT
JzvHNOLVVBAsvMwfqpPt1joHapMAeW0tQ8ybjm22G1vdh8AZjGAyDVl2Ft4+MdsMQbi+9ZqKlh53
YBBchzFiJ2flXOD+Pk85ODjEarmBljLFvINhjgKkR1H7pxwplaK4DDdVOBa9qHVsT6a5wQOnv2VX
RFkChaM64AEZmEfa45ViPN+xi2eQZ2axK+aq8W7ExbScvORXivxlSuTfMO4WCx+y9zlBaZs/qOyS
rQGm6429+eq/OjjbvTkA0CTux9xHFB494/4mJfI8Pk5tuaHGD2tKjqIEI2akwr2s18NjISVOLOP3
rjUB39LrYKwKcmDzEZLXaBT5LqI3qoT9+ErZq2pK3EWXCvGn9qzcV5NGCaVV0Wl8M0EYARb6mgZo
SdZDeAlVKpfkjVFr27mKZrBQ8cBoEGezH4CIO08GxP9HNUBnweFYSEpgQsY31LzTRoEwLtHFODMz
1eciwAcJTKZUmNgZY0i/FIrccn2Ak8v7yqQhdcUCIaOy1uWXDxIOAGWDg8v1A3IPoBeneDOQ2ZDg
PQyoHOCykWoZWgE0AR9+PGmR/Dp9zKREjEJoevclICjdcdebGQBPpmWp9H50USceRSuiinCDBjhG
Llt/7HzCi6lW+wi7jNd3Vs32VxT2rvu0hqgjyiSUj8Gw+PfsFjeM1OSwyUhfTq9yYFKzLnPbzIlV
WqEY1S+Ssh7ronhto+zPTPw2H6fCC28pE4HE4bb6ekt1jpevlkR+R//g3ggwvYbiuyi4lXJGS1d2
682HKLx/+t+GxN770e92cdUkurkNTGnhfYyfM+njhnq/Xt2LaGGpNMrWdzsuBN2ZVNz0bZ0KcP0m
DdYQxFYwcpl1RBPSBzs6BFGVZJPbtni0tCuKz4hOxLxtgwKhTQoNO3K3zmK5NaJKfDLT+z9++Lcr
ZlrfcIg307C8Omz6vh+ZjM8jqX5qqZOQmNgZjaEjZ8tz7Zwx/u1acQdPk8GRHooOylREeXyERS/n
btnVZcV2KUJXRMUiIJNrkkYVymnjgD0uFRyjwckLY2ZuZOi+y/MRmOq/PaTjd0cN3Jb3N1FNtxUS
Fk10O0bIHFu/Eagi8JUcw05TCBLu6WQVsROzEy5Gys+Yhnh6IeK/tujWFjeSNdazs7/aybYb/wcf
mACPF5KxOhY604yyosVE8nKICX0QEoc4o9oRYH9OmRGI2zE9Op4EyJtl3kT05rOuESYsuaVte0tf
6rFgrCyTfx97MHntseGp/uL/yRuMZg8BZeAw8zhpS6WT5yKpFGqHR3B3qAlvakQu7r05LspupMqk
hsr+H+k3ezDdhckQJj/+XUXs0Zo3LeGTp6iMZrNnW8oBwJLfqBulsz4QfJAV6T5RHzxswQ1DpDz+
/Obf0a0auVKLBR8CWltCH+jBKRVOd1U574we5m+F6B3mIUZvWMRxZRKNmILJ66vo09nuz4AY6ky6
HH2jn+P/pEAz0eIJUA9rEqlMnBXq2rFqFFuFAsJ5pMBa8s8HT2qqlo2+lGfCEZzJtJVM8HRe+Tph
ZMyjS4UWuEkpP/cNqc2rx6lQoh834zhDFHOoZA4xIb2bdMMQQoxHoITpn4rGAceBhEXNjfRvjOTF
920ogEW4guYPstafy2XQn/NcktiC8/Qk7uh8IUMNL/wyB84nEmVkrgi7Voz7rHmEjye8E/QI42yH
l41Tb0KdnN4LIhNwExvphHs1k0Fs/rwyaTIJDeU99erIyb2RTeGOvxzw6KvMpuBj2UNmtynwpoaZ
fUWSOvdENymFNknb9+KXBUz4ENhljDYVvmCDkAoE1I41vrGs69v5figSuX0HlR6MnPSX/KLvS3lk
W0rkDaM2x7n11ghEgHt2wsPbUntrmCGtqhEBjv/jZ3AmmvNpfUn0+V7kMipl8FGAN3SWMHs4FdhB
7NJ7hfepKyUYQrt0bR00n4ENCby4mUJEJRzuo+8CbOo2J4LLLOa4Vhv9EpSKvUvWuQavd94WIq6L
VlUjgzr+4oM1H2WQa5R92xxuU+t6Xlf4qLR/HEZmJsQIAh/O2+LsB3OtKQyepe8mXdMdRIV2O2Bh
QJBTgQjwLFtAmmEw1M/TWwQQxhIMi9u0gWcDfWH3NSqehO68cWhNuk3MqKNiU9kJ8f9fUD0pQXQk
9TjDy18b1+mY+G7fQRzG4sRemYQaW+KOvXxMSmyNpKGwf4zCuL/VhcbxbEnRFWK2zcJybb63wCHK
iM2UEz6T1ojLMgWmrQL1i7qiQp8Iy0hCol+gHOp7FzY5nEnGwigpOnVI+fg7bLHFlZGcM0V1akrL
mc7BUA43CVwieUWmgeZunw+NTVar56idu+9aw4UxqNntAOY0WoU/KVpkM57J/T9MRlCkPGR4LBxu
sMf0IkNoQoX1gE2w1eQEJ8Kr9yFiPVJb/1UWaFIliZRSv+7NNzHGCjpnH7ienikInklUm1Kkdt0w
vnR8Tcx4DMQ72HyXdGKwtF8zvbPkAHUfkyhBwXE/dO2O5C1exdOI1yXHKKReVYcKw2kb9dhW4APm
rWMeciPykCVTY8bspZX2CTDgcTf/dWTp4BG3VgTYsRMdKCPqVrOBvpDjq9GU1/K1vD15iV2IyzpX
ktU41FBgtPZFhgoXHzzqaMNpccVUd1lgwAdmz08ciyapubTGxdlLT1JpNdgIJljXRyxZeS+PeMY6
FymsIVjvFXOQFdbSPV7bhpBHlIQM1y2LMlTNXNv3jMwNTu6jc6cquTe/pubJrJCOci7FZEqKuWQx
3UNgicBhIzQYIa8H1Vgt04MBbN3udjfL+7Bb8YMBpdtwFC1Eu3ScPSZdeSVJOQ05hHRVyWcXS2pD
tvm9aDxHA587shLfu65TGea1H4OnwE/fVhlvwv7FRjXekkj0g+IQKmRdv/Kb0Dp0MG2e/ASlNeRU
iaqODijSky/J1WiahLKu5XvkFYaPHVjkY4DyNy9kPHB+2sQOyGwQ2J1yJTRHuZadb4M7VMDqxML5
0YgGZtVk+LjzMR/h6ltjKoUYOb2skWXNm6Vr3mHBbru7RrBLbSbFHFf5C/Xwa4abrwBLqmfn2GJo
mMtNVmYBa5x8UzmevOvhnYiYFxFKqR5n6LJbahlO+vehjyjyjShq94IS1Uf8S2ftlRrWC7hdS14J
koDfzifCs5alCfqQoLi37SgoNxuJxR1ieANszoEDM0BF+28AR2yM0lAV6lGgsjZgP3NH7BXRcRxs
GCuIMfLRTQHXBNPFykvoIKgdKy6NcVK0rFTn0KgN9RkIi6ypLsgtPgfXRE5nVNQrUTQIcVSFjfor
T4pJYWjZmj0D04j3uj9w4D4nzGuq6x7FGIS7zN5NzJMIauSaaZFkEudNAB6dc3FK5XC6dNdsv9EZ
YmVrsYi+VvC0UvuLVEHxDrhl427GGzWgVLnB7UbPpufoJnXTbTjMTeZAd288hhYKSDUFEwTXD3t/
Kkmmfvozfbha5yuv+Lw8Ns834uis0hjDJ1Z/eKaaB86cR3OBEmq1uoTSZVK1sXf3bRzzGgUujpIR
nMlvh+Xr6h9614CZsiFDCQrwqymvnQyjqhZSRpWgxPr803FWHOgKJ6o5mvWMXrSC3YJuPO+6/w4m
EwxT+iApflD10rWgSCMNAKcuYDfHgNuC2u4Nu+oiBcQ68nXBamnf2fU5qFobevKkmsguGnI9a17N
5WJdpFw5QPIJVzS9jHVUMbBLcLhK3lqeNRHeglvZDFINX+a0DfDuM8SdMWUCqXkK6snbqlubeye5
/1iy3FSlRrMQeOH/LooVacE04yXSkCyfgbSE5bS9TGmc3FRP97/r83fBuM3YN9lVzwTatHziEcUJ
+Z7fltzhXbAG2CsNIQu8XYFUH9RazLVyxAjXNeCALKOYEYUsHuoHfTfTyL2j3mw7wzvMmaRGW1Up
nDvL2OxN5LF7E9kvjUQiMTTFQwS+GYvri8qlFzf8EomyDg/ZjVA32FQYian2EoCL086sbOmlUvl1
TLRekHXHM3gMJOOfq2avGFkJu0TMRsXJ+XYSQeR/yQvxC4BAUJCd2B/fPFvlhOx798RnFc9g0UqG
u/n/C4qHZC86GAIbri//EgRxReqT1jgs2LjqtLsYi4rRWwDewV0hzbB39n7emuaAFFmZyzswNhNG
yfK8cstPOazzgKU1ZJ+oNI4v05IOM9z8wrrcV2/DHD0cobZl6WPvoDPsxD5U7k8RUW1RoWnREw47
AUWy7k7K5XgPuph63ypd+PVoF6GrV4Ny97BQo/DsxO4tx74UhoMJ85lr6VwJx45ZxEm7STlHf0nW
lgVDwbeEubnHFgHQ7/axeGVb0TDsTp1LPgQKQsltRjNqYfLU5Er8VWykmNxVF1sk+9QSxgFYPO9j
JfNVuj3SogIdZontbwvtxkABTsER84IiHyju7vzZ+7Jak+2yHTCXZztIgPou1xYAGJYtaoei/BLN
NzGKrcmX03u9oYFEDtFUG1/jPWXV7Z9jQGkZQk0KYRlqGogoVSP428VMH+FLRhnaHpJ5QbfYu+i3
y+6LevOuNukGPxvczSCvnz51paiALC8UPsysCRNhAuIhDgT3sQOjLuYRlQOivaXrvth1r8tjiQkx
sVKRW42Q+5+N3LFtNzZbgoRDsTT5ZhrEodxWlEdyofG1nd1cQ6I/qob8BX1D7JLbq/s5xGEbiCG4
GNwDZc/hC6uNWasZBOcPH8WjUscIiS7Q2FhGrW/ZNMPvcK8X+Pvu0bAzTtfNkURHEDmKW+A20aDC
wp/EhmHD18kykq2v1lZLRa9sxBLYKUrvyqJpzLnKu4/vxN+1sCd6fxWpCqWDwUWpwTuwMWvCKkX0
NHSVR8fzn4Mk8KJXSswE366b81rGqiYJtIW6r15Sp901NxqQRedtfhXHa/fLbExNRu0nK8qkBzNH
KmznW0ksqkBsmwvNNgHZuJNNtI4OdhG/GqF/EhX7WSZBhb0DmXPTLrPfcDqsDNz8eqqntmx90Eux
CpdBZHTJ8C5HGiFjZGy9+95G8gqwzVUc3F7ZjpNg3QMCTqowp3OqIPs6mHKcZs7Vn88+w+r+3vgw
Rw0ZtQ16CvKnUKgIYzq6J1nlhm2yB5hzMmSUgXjfJpQeSkrWKVwuLqEuZdC4HdD/x0/jpKTX5EAF
2qfCK2WxbOLT71v+veWT6aL7paEOQ6dFP/YEfb9KR1BKGRE/XF2whHJK3s+Wydmp0iMen793JTyh
4ZQRZEqdq74Cd78RSyV1Hx4eTOMl/7XEtfXkAFOnqArV1vquwrDloobqfi0JX+gwZAJ0/FI05GmS
bqXN3t5fXONqBTJXAPFPuabSIq7JMUR0X35lxtWEcyCpyil2KE50Qde8aPt9NBu5hN+kOGNp9XNQ
4wYW2Qran6tbzkrzgPadiwSoUqzqjKQ2TJG/K8avCz4PYVQM4EVx8asyqjGagmd58aVJOqQ3Z5gm
3nkhcWpgxdtrX4qhVRT876++Kda6XBFds2HCHJaeL8iZ5LFHQJNoo3EC55taePbDY74ZjPtfJTZw
Pb8bqmblhgVfxhOCaMNi4mpUT6GmIRqezWPP4CcsyUy2IvphlOK9il9VnDAeC+nr/mI/WbHOkqiz
s54L58hIrrvYHbYJTyPDrF4lkP1Kkwq+naY3e2139JKaDgkCm68jFsvl/tzKvDBDXxRsFI6cyQ0i
tsQsaQJkonNJQQKbUku8j5+6NQNan8JThio6GnK7a2Zd0HT/4aPPUTTsunkYZRDW/iyPysNNmddg
XgCAyLsUHfcmqKHmJEy3qcmGEF7LKM6eBDgxSRa8kkcFcz1Ze1N0x80vg8oTEmv45niQ+rMaQIP3
jxOK62eDUmPyYe9yiKievy2cJdRfJSdBrkbr6pibNmk+1DvKsZ2YNPS5LZZFb1M5jYT6E7oKrkhG
OzMi2zFqfRA9qxwOP/lH1jX/F/1VGFIrp/dK8cctH0euFWpY5AiN7L7sG+WSqn7cxrNzhWgJs6ZP
hxLx296hPZ5q3Avs7rs1yqEd00f79glvcwlJGn0dH8q+h94c26qcprPJ7G7PWmdUv9EwNQ+1WZSU
wDfACg/jlyYobOzcwaka6oT1v5lpHN2yXq0CRe7Rt95tEgxm0jmKaUklBkibB4O6/IFy5U2rvuCG
QyP78RIVx4CFhH5jdX7qfPUzXHQL666JYXX4n0siB19MDQ/oyOwgxdcMgVo+wu/d72WGZIKrHTo9
SzTXwsfCXZ8BYLLmcFXNPR+hN5qC3r4u/6xarWptIxoNh7QdoLE4Z6jU2pQBb+0eVpta4F8QEL/W
E1cj2qnAjZvmlRoQlmUucXAq8ubMomreWu7z7XmsIYdmfH+kWfy0aw2tjzVfLCpWN9CXFWJzOsz8
3T8MyGqkwyjTZOIL+gmesjljti6nzv85HUbznoPkUm/LKvvCxTVEwuMRUgsbxl8dKDABM2Ofscpm
4RZKJZ6yKvVRbg0MAb3mr0naTq5Pt+FoIdiqA3J1raAbomv9FCGIWN+xS+zFRvaYiVEoCp9eN5ko
CTKFV0iqeWes9tDd+pnuR/40EDyEgcm5in2NAGwwozsNx1JAe/zYEPaeOxsWBTdvdPCr6BX4XooT
0cHjGtElw9g+RYkbbh4yvCrDyAnZ9lLoFHiXmZCBlgYgz7z94Ypop8kgW9Okxn8m5E+70ofxRGxv
YEQEZspf1ZZhIXT5AwkSlwmv+EqlDjBkCOVywn6tZk7fiIZ9soRlP7fBF09Brw0V4qd9Q06xdKls
30cHL60DBXFWVmv2zbGyq8uBM2YNQpbNDyIP5iR8Xpm8gcZwb9Eacw1Eli/TPmQvnoyWr06XUWI8
qwswUa+xCAdHbKL1ZI+LEJ+3MWQR+Yk+5eTqS5EPrzrctSO1O0yNMcFRZ58b3pQgEwqwrimGM4v/
zDqzoGdcdINgJv3UJNDOf9uC/abH9FgSngfqXzIcZPb8rRKbaOdXdvt2PQbzFQyz4lsnDuIDvkqO
pl559o2hAEmwgZMDXR8fTVCZOFv85hPyM7kXNpsdyRd2cuCE2xFTGairvoc2Yuf/Pz3dXZW3/8NP
02xn35TbNVRS/vajT2mLBAuCSxkdYxsTvs8w/uJUdN7ydf1BEFh0E3i7MTmH9al41y3OWuIrVav9
gFs0YPhl1KwR9Z5kuZMxbhDPwOzoi1hRe4Z9V2fc7a9jtdmlJYCbel42SP5crp9qXgF2XO0eBhAU
HsK2MB2yYMfgDQOl44YvvJtWqrbEn22Xz64v4xJ9dEvn18Ec3WpXB523pm2kHNDejQ5AUIBxlb8x
txmlFxdqNVJTTg2xs1K3KZOxQU8053iskCYmgvai7LZHfxKXENuLlxL4OWjljk/abZVaNOh+/Y5v
eSQcZyU04F2XRrxlyUIahYH1tuRvXvoz/hcJNMBYJbC6oatX02c5VgLFEL2vt8BUaIH1iMR4ox0k
zlwctKohIOL+3AQJhsTHbIe6pJyeMkpZcy510Kpf1p3W4cHzGAaIJAuaVeCnNjdXOJqcm6W4+xsY
wiXDj0MUqDy0sBc2e3wHDXEjiLQMMRR49LK7STWSA4rgNbNdGxWbY6WdyKMLOF0kOIrSXr2eWE/8
vHry+LsTOA7Zus3/GVhrhw5PwZBO2e0NLv/2GX/EBxBRGl27qWms3Bil/O6Ka0joXYzuod1azJji
eqG+zgxQCBsEZPOGW/dhk6IAbArVAPkGpf5MxrZNi5iJYlZrE9GPwXhTruJXDTrkUz8yEIVJYzxe
l7E5kysirgts0uixhDAHNHzKd3/JKgUz7dBzmo8G7mgKyhMS1TZ2KcGf5Px9BC3EVAVNYe1A6i9g
q6YAnjLrFOcojRkCDIzwhOm4k2KsOuHhHlife8sxY/Wwy2hfsKohB+C28giwwE8USzwlynuvDVvH
CdHrGo5GhKctRUenLOFwmo+tfEuhcxqICgTFcsEkfnX8Hn7RpiuBdwCPmyTwvsxgsVuVaVtSQe98
qN5v3j9vn0HiUD+3J5waLldher7+hLOZ3lWbNfYLHwPDBhZhrXGVtZKuLrNUokSR6NpsUnqsXGyF
qPL4zSM3jpniUw2JF9+8ibbx7PwYIiHgKMeWHqzR5zJ8vOuJR9tECP9VxWV+sgAaKsx5ZD4/XVt0
UjKRHXDTRW84jITzCwtFMwC/Avng3Nb4eH1/ankSqGE7mLtfSTkTrNspSV1BZfDYm1Hhd0nrTeD/
dX4QoUYkrfivrUNvFJ+QT492fGPo5IWebLTn//B223D7IpDOdN4oX8fbLVqgSWVs1HR6o1kibOTx
/NkJHpUppkdXrQiaWZlhC/gV9OwPAmMSgWIPwJseUZMRWj/tjxDPH9FpIwYe1GawNLxqtRyAQlVV
MfMLuMs9NkuO8gFvimxgvvKT9gV123fqFWj1hO+/y4F1RM0RIaGGywF25CkNMc9x7T4d5EEegBoh
0UE8vpyBY4IWlZKktQyfVoEJZr1pU5HgTx9202aA6/PiV6NKblraW4BcHNps6q2ZtiVJPKbmIVEN
uXN0Wjr9sa45TTL+M7DJtNvVCitHtwAKUupFdUbk5v8KvBzi0RDrAzyPQPiBdV8RvODMezmIzaEQ
QfveTU6jnH/d6rBW0luihZxbmrtmiBc4MmYjaNvlmLvQFI5O9RDVORxj/b/gOJelqzxEf4WbSgQm
/xcKZdjMhNZpRvzuEmHJugfdEr2kYPiTmp7CbT4uEmdM07qCBTrQfo+8tPCWWPgB7bp8fVW/Gavb
Can7c5Uxh1vMUMvWgaiZHydeeQROeyJj2yXvyqwJU7QowXMEmLZvU9Ks3lCt998HelHZeFLK/FNI
mzBToGnuhehAnQcYHYvGxOHTAu1xS2hMGJ0Gknzhs+1/musmihVAX/muK6HARHePj3SCA8G6FVRC
Exw64ItURAus1b1PGKNURTxereqfX7oXtLTSRfxfuzEdSB0p05MumQ3bE0qsoJDT/euQkaViaLuv
7Rc1Jw/SOF5DUl2mzHFe97nzTKKCYAxac9GrKrjVEinnmTzV9HmtF17yMBAT03/4G8oSJnWFPgxd
XzylvPDCI6P43W3A4JEP1l8+bvwxq36ChEXxv7o6ipiPuFNySnJDrDhbaCO1GASPy9lUwt6Z9f9K
suvBto6qpikRETP1hHatGBVRbeqEG/gtn+ZPCdvxIASaDJ+I7AXFHfzeKhRD51qvJh5rqHnmJF57
5AwChMstLydCG2eZSQGS0vIjiLS9W1NCP7kC81WR3+Nm/0ctfDQgx45FyodKirnrooUQLEKauOxO
hxNKLwpM6ZPcxMDQZuz6IrrUDrDuIZ7INwjH55KWkoBJg3XbrR0qQ7GfZl/m+k7rl5XLWvl+23zi
JAOFvuxcJSPkYwV6k+puEq9etU6XCj7EHUjaGmkkftP1q3w8yACiqbruJLSyi2vdFhS8QYS21d7T
BDWjsTbjs6j2bhvknT/7wnu5CcLhCh0RzctMrsjYEKCFyEBSh6PbQFIQFON4PrzZ7rmzmQFl0hzH
xbxWQgOE+CpgKxlVVNB+QSGcM3vyXLni+VehAfLiJ23YCguKWca2RkQfKWnqp0cfO3zW6r+QFUkR
KiyYG45rjEUgFUlHI4tqOlV0bwf8H9l05CLdvvEDGvE8sFqvB843YXuaaZ/WKFbPzCM9wnvzMBWK
hBiSVDljPImmiNpt6IJxqbYTD1hZZ1/fistW7fZWcPZzTrmyROhRCGYcH5p+0ZkGKUCbvp2vWnVs
3jVH2qoEQyJm+4lIsF3X8XD+5oFEfhutgXz4JV245nkLq+EV2bi4SwU4dxCr6tck3ax+fi1NxpGq
k4SXytaUpxWIVk8yJReHB9ieJ3TSwKPQf9gDeDZCYf6r/Vwy9i0ORiQnv3dsIyAOOb1IQKmxj01Y
1uTEw9FLi4yr7XgtqU1J1gfjCQ3jZ60lgDmEX5IiL71qtA7nwR8hO4F9JkQv2NUDeGducZ2T7X/6
a+5UYowmYNT3dn7HjGhD+1uIfvAFBaopLy3EHIjQL6ZhrmIBBcGjc7PjeYojh+PNRqaIbdGnm7LR
WL7Ken8JV+MBk7wGJhNLBD0eIyDXnYKCuctDRvPicXmYK5UYX+lfcDjjEvYfVq3Va0frORz0LksF
4yxjPVRp6g/YaruxwIk+UJO0a9ZVGankqY3PjZ9h+P2S854jTqaKs5JK4K6jc4WpNjPa7ksGux86
29/aX3sD/OEUDH2DiIvXcLFQNDGxv5OYmI4Tw2RXirPMu3YK2+3+2tEESpG+HGx8wUORPyhBXlcs
AEhe96+QuaJsegbwsXJTd4RHpZfG49g73I36xGI5JqH7QNFdT5bRNBWKtNJem2sk3kIMCdaoFQeW
/nRkPcuxv1lLb9d17YHPQNM/dQgLAmmcH3gNHO6zy9jj6NodzIkQn6XfjyMEznlgXV76nR70Muka
wkoU8ue0KjePXHssXRhIy9NNkob5zfkSx31bnQbt8DfqRoVfGtomsrC+R9HcJ3V3RQ22WfFYEP3S
nUS+u4Ob/m8wsflaUr88sfk1r3GF4qlIRl60ttiW71KCM3U38uTWFC/5qRBOGw+IXzQIeCqLGeb8
gxIwTc6gWMU+5zY9PzInQ3wVJZt2zcpChC6IixVw21PH/e0aA8Rmo4euiz5By22gw8g1P03oVio9
Vt8Z6MP3XSpHDlXoQ2W74UcfnlkfeBgBGZwnP0O1403nZtCtAXHmccO3jZw1rqyRzsC8djIuUYsY
hnkbEH6KhjPwraMMDqUjpqSpIHKJjQkjL0KgPAi/CmfcuKJlwtFng2mDg5kRN3AWqVLqslTV0Paq
lkUCLYw/4pMLax8L5nHkktJDQSdz9SiHaiB+HkUY1yQ3IODoN32MLonAxLKuu34ouNr9bkGbmHWa
i8uVus/+M5FumZ5VhEnSG/mMr3aiwcsLL9icIHpfxNyjgag9ps/K1JPqg8CnZtpEUuY5KqXu6Rpl
y863l6/oGGvq9shg2uIiopjeu4TngmP4ETmIviSy54dCRHq5PyrVY5OkqsEtSVOeT0QXVnOQoVj+
DTNWx+fugKFuk+fYz/eSBU76oxnRRgoTsOGxYPTEfSDXoOZtLLlFcQ3WiN3gU+2XHJdWS98OZXOo
9PUh7S8y5NMQC5Qi+L0aHsDSBgCFF3FrvsGrDWV0T0OsRUPQXlx61VLGwAMZLaHE51lWmyKuzgrP
kpqE5NXAVNx/PZCHMvAhM1wPsAT1IJne94Xz5MmaS+uwfXSDaRuQBooNlIed3vKiVi4dxtezlo09
tU1joYkYLAuCTOG++luNp5ajjJDiY5FulFweKVPslvEPNmiQDfUEYeT4i35NoFd7bJKKn6yQTHGD
8h1lVx8aDodj5dDulFylGjkfX3jAiLzSWyOXEQOr/sYe7mF9wOQp9qri095U5s2/1O4nBUtNVgfx
tGau2D4yaaTVbDjkQOp8UqvO/csh2Bt5zKfh54XKjKbRzfg1UKGW1OWa6v8SFOIv1zw/GsItdJzr
belluAkACIjHxxQgb47gilYiGKSDZQHNTWbUIYKkVDC40KNUsiIumKgCMk2TkpmIypjgsLrwg13E
S+QnWk7DTnJq4oI3/VNpkEJFSidgTrljNHYCr4hV+c/EEl7EZlUHY5TjptUODlScLx6CfzEGEKCK
6ISBZSwi9VwqmgF0G0lSuj6u0EWGbPatHBOaBBtq/+yHor4nv0MxhovXO4T7KouUVtWvAKn8uZ8k
mp40cMIDp2mc60P5QjdpCR66oad198jU5YnUvK1NhLyYsySmzFEVWZ9XAB3MUqS0c2MR+tlAFHQm
yieto4dTspE+5zKS9oc5Cskeo3BeiKK0Q5MjGTGhQs5lLBk0kKXvWx8D89hylcGTuv+8S9inifAU
z6LAcrA4b0mMHcCbHTgdv6O3PX6nyf9L7e/IYnGkBoTppLZoF5rI9CO7pMS+j0culzJTFswcm4iS
LsVnUcXLOoPrI8mPP8E3HpGGWiHCBEAaOHhAthHGfLE1A1QS/VNr2Y+g8nn+po8fiurnILursNuX
1OMyWm1nmk/khmRfvt7k8bSjjyAVS3auVTIkdWrEsK/r4KDaNk6T/xStYA0TC1sE1VWixSeX5WGl
kMCNB/YVNYN1OKGhy21cMd/0E0Z+WOhOhs7pM/K1pjTcC6oPxnNweK2J+Em+BEbL5ztjvxtx76QQ
FJ4oW0bMRHTR5EQTfwCrXgTWMXXcY8S0dVCnKNvOufisJEg6BFmmSKw0jEYsE/uI3rpNi/6H0Ap9
XW9m/OdrEQra2nBIDHUWQe65HegiRxXqRH+YYBkot78IehXJ8xllw4LDUHBO2LF04RY5zNdOXvaD
dFKXUjIJehBhJsxEL6d8P5EOQ8qTtkZUi5qhS+6kpiAythd9RmkvClSy2WRHTsu5ozeIsH6ODcCl
urpKmNtP2twwxZIvF1bcHCKjokNFVdA0Au1ftn8R30Y4fuHMc3D02EqVUZNNnICWad0ALBQ1/7OT
UUZsq98JqdMzge5R/9PxyDpxc4ObqvlcPrAszoj6zy7tiJEcoxVjtllU9lvieye3KAWzTbf7ZQu4
5zgMm9ntNrljBDsatwy0rFGlO6OnVQgTggaZSpjES7L2TAVpsi+DeekRU+57ifU6Ymf77iRALDiw
YYB+mm0u9+VRka/9zsPvpIOVrlyFmoHbctcJv7w9zKNEIhaqbsShoRk+T4kjRC1Z93qNwVKrerPJ
01uA/TwMLEXVxNQA9UXpgufALbxHt/hWJyI94/26cIpO1ld1AAZzOJV/mv5hjYUmfUZPNYiR25YM
20bb4z7vs3Do2sZ5pyG1kEvGgMWXyxX9HV8AP0cYLpRBGrW/wZqU5A/uRL+To8rPiyiTWak86Ax4
RtbzZvoymZNMtkq1EXTxJl+eliTiwfqTIUJ8Tjk15Hgd6UdTMkJxaz2V0YxKmfj4tCDfJyZvj4L2
hRexC5wWdkjvvO6Te3Tbfhcv2YY7Dn4LRpF1dI24OeFvDbRW1H9wwDLNufV5BFnKcq/0cUBGm9Ce
2JXJpbCRa80XK1hghiAGCYiEn3Co+87vwVMFf2uNt2Zb29yEzpW6dm8KBthcDOUCnHcXQWu7LsfN
T+p3t4C+PHo8oRrE+t0TTPod2szTs1+W7fiqCzPHIt5GHMh1oaAUbeK4VpTr451fCX8g6k0+cUNm
Z9veFxRsbYbSQNKww5ta5k0MXdptnX7VRTF0bgISxMULGehr+TwNbdhNF4W9uIUsj8W0CIfkVmR0
9VMU9tE8Agg2YWd/kLlkcQ7O5dpjioo8oHoaHaupGmfLFOEFan/KPI1TeFlarqILvVtDhBXJXlD8
mZ1hfFkGARYRJTFgkIEJlgC4NK4tSdYfHT0/aipizFHgU8OFnarQLtJ0ePMAY26UCgWbUdvSjouL
vsML3GnTppE4Pr66p9mIBtTjRwQFr7RD1S7UwArNC7PBzeQLK4rrLDqUbCPYbVEOdcv6aj9dHybg
TLSLhT0mXhfBNF8BitXfe+R5vLuzNe+tz5WZVrBDF6/UnaKyB0anwqnyty996L7+PDReYH+8O3wX
w6AEnTdpjBMs4LSBxNASdCxMnrR9Ybsd3ei0dK3znDhD6WJ8tNtbEla+u25TuB5XdDDXF41gJeIB
0kwM5I94Lcmp5FScEcB+UnBeE4BiTLAcWRSR1twksjydO4+g4uhQB6GoXn8Cb5jVaQI6Yv79zQDN
2EE/cqQJJuX8X3/n6hsillRQql8XX4EU9aBVnjjCmB5tkn6lLqY3dlhCVO6EPCKMIgMYWaByCbn/
hrNV2a9SE3u4EBLC3MDkPXcP0WHueB1goqUkv2vGeZGMj/a0M2q9DeAMGL78yCTVxjCIbYKUZYtX
gose+B/gRNKwpNQz7mj+75Qe3Kw8IAjP59Ue+tY2QRS0r9idRNnpHpL7SOkxQG1PGfbzSvdLWC1q
cf9WBum5wzTR5Q4oK54FuhLF6UhyWUbz1TCMVJJmpwlvzqq5BImB8k92BfWLMwtRuhrhE8AL9vP5
uaJ8aYJh/JAx8eSMfgRJ6jc/2zWSvrG7hb1T7OQiNJ66z+D/4OAOLmi6rXLAZi7sqFXTo5AmFYNo
2ImYb+2Wgpo6eDuN1faMB6mUSKmXSOsX1+f7VUwU+VjEGfGkwkQBD50sz+ybdOw6HJ7/ipgQAxzD
5jLsF/YXfP3gYHW4CH8fbDsl81fzWYMVGGJ3AedwiLs9jTT39Y8OgVjU5A1aSb9umNKx8/4tGIi/
bpimY+MeZrV24Pco9/i2pf5cn97kQQfFAQDU5AAnH7Zs08SIAC5eAKKk6JwfuxHkrb1xiIfD6Wab
POuqSBdWI2AnL2lFcPf24QQ0jV7H7Xe/gSxQEikbFWzNUlAjiO6KMwstAKW4a0tX9ptxnUsPPv9Q
pIip1Hftin7MCP8ODSHzHDPUk/9J4rzbshiXlwdiVsNi9lUeu7k3M8REgSesNsZo6ROdEToI0Hdp
+w0BB+0b/RxjXfMmk3ijiKKVN2ash7b9eP2TqhR8rxoq6fZZanidv8VdVygIpeDlXAjMG7Kgoe6Z
fvsPNYiZrN01fHaXmYgylMSZufv7f3hb5bZ8z403TpEUBgRlwPOD0jBqRhnKM6B3rGgE8WFhm5OQ
kWcP1qKI4e5YVb+hRZDKTRJcHzse4vOH2KuA2IQVz2k2b9AwBr1b0tZOQTHgw1ZDeaM8S8sCfLkz
ceWlexzX2wgbrKPVr5GJFht8ufPxAfVym61G5q8B46jWjaEIGh6P8DJLGihXRi/LkkzjVTK1XV/T
iqEKHPwhcSOd7+kLC/OV4yhubSfmRt0FX/lmdIjWKMKyyI+UDRO5oYDDLDwW+Y4JzrVwoa+p6Dxv
MTxnGx3V6t3oJrZGU7x0mI9OWYWf9Q292uKap1IjaVvIJ2T742AsU1FhZVo2e09D6AMGrl94XyPo
WRHMiX2+mDxiGB51TcibyuRSkzcX/nak+pMu3H0yBcjeZ5+OFW6Jod5yatct6gWOzaG8NJmbZVY/
NK7fDHhE1yHVYRcC/QLD2m+qtqSXrXiUB+7ASHk9B8bmWvRPytIeYLxf0p7WId4CCpXyWlB+agc7
MzKwX2K3yW0gPwSdaNqNk1N3xyNWwPcirDqPYxpk2lwx+jOuINAVQAEnEXP6LCp+ZwO06Q4ybuky
Aa9B+//7IKkxXBH2kbp6KpWAk5cQ2MEyllUQ0FU5ALk2+JJfYAngyn1UOpkS2yUOi+39/kz/h73c
75Mrp/oG9GHcG8Xk3hljTMdRk729t+Krj5VSc2bgkhhRjKRZuyJ/NZpYeibBruP4+Urv7D6SRAIG
nRqtTQucOq6wLfeNQmLUQ71eOFHNLoPiOP8ip4bxV1Bht/GZSS/yKXgHZJ1RZ2c8tyFxikvTpp3r
r5dcnJnkUTYjLNcDMFUHPTY0tEKiF1aUzK+FScS6gDM7E+TuEn1aM7Ox5yS2lBThvGu0/t8zHhwe
UUAX0tIcLQvizIsXtGdjEKtVd02gZu8SK6HEzQtLemBRaoktwiu8oRvHzUxAjnnak03bk0OyFpig
LCUKlTnnlA==
`protect end_protected
