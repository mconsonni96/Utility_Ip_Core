`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Li0RCxpIiMDl6+DqoCQ2cgVoL2FGciTEOdr63ZcHr2IbDmdvt5o0FtZ97oB4zes2iijDKTD1lV7z
wHi5t6kTxvMrahxkJ4uQ8Wo0B6q5p02t5auznSlQEm9WF8w7fy5O8fxzx89xo/2ODFm30gTKeor7
gai5Z76nWpkBaD2aLLKrqpDtCQPk/yNDODxprpSx/a3mhdhM3YnTELhqkGkWMos+JfIhI727ssqD
VGsY7dsLOnHszC6RQuzm9vjKRohr046gnNu+F5JCjIl/CH/gqyiHiMXl84CPtEVf6XjqEIS8kPlw
2YKtshvdGg4zLctJFZD8qYA+XPqqMWo8euXkLg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="aNsevbQjq/3+lB1/tTrUl18AFsaUwIfPPr1E1LIIb3c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25168)
`protect data_block
w+NMyaMIaBAyjhcu4BdKvWz5NzdWl5Bp/pDq2lM/EWCXf1Mz7uWonWuLuuEjNEsUb3r/ttONBl6E
avZg9uyVxRLpD3F8uqZnloJYqvs3uED9esTIrU3eDcvDe5nTeaZSz0uS7rZywwFvIZmTabzYC60D
c8Rio/MeDgS/WUzPiY8mgiz4qA0wCVn81DkmfDCCzwrvxGUfHd2BIaA8ACD3J8aApEyzDdpaNitZ
klW/nr7UTORZe7W6pyS/0kq7oBTlL6JbJ3h9puDGklBZQVfgmYVvFX1vmzwEM8YIFhUCoXk5HwCO
wdPxAXjoVw8ARfzEnF8TkoNoPwH6VfnOije1/KX+oshpcpS9HItM9Z5xvahy9Dg65hontry3pQ8U
c/LxWIj8LjHCxLxdPgU1Wc/PK74K7oLbZw8K49gFdELtlnuDrgHdfUkqRonlxHJ64DU/4bqSvnyA
opq/SqnQr8VHCONlZq9NChLy5v6LzPYO7gJujlcjh8rO160bLAhTW6kiZTDlK7W8y7nVT3Lq9OGV
RT990Ve00QWdeC5PbNTi6N6zcc/FpVKQdweo2gssBsPvTWL14lG6/TXh0zRUjjA26f1/iGPlQMK4
O8aVRa48hxvhvALX9tyy19Euc2AoE8W91qeB/F9dTgkOTfRuBxrJMgVzrjKKJaF+P5w3ghjn8TbZ
a5x7I4LwAl9WFjNfkfxnDvRiiViWux3Rmd9VKtlPAVLXWakD8afyHiYpfL4JEQ2sdJa2XgsBn/YO
AsmRP/pbeF+wkDVlE5B684/J/GPRq6LIDaE6yEPZGIO/TrPtdKlYKh1rcvCzlX5y2pyEDy9qSJP6
0Re/PyvBZlPFVx4onEt6k8HVQoR8PJacBbiOsM5UBWgc89FwkDN2v6NuPkVGqC9YbgXJndOnNR4C
xw9gTW/QR8KnD5ZfX2aFvI6zkrhseutTBKnZCYPtuRDUVXSxfZimFvjIRta943BT/1SyAt1qJLb+
VFqWC46AvMTFdyFm2FIltl8J9ulepJmBLTv8sZ7VI65+SKb8bbyBOwrGvA2Ze8jmLVKYDLROV2aB
9mF2V1s1UPKP/3V+iG17sQQv5egZGY+QvuHUqNgvO6N+7TfXXyIOAttetxA3nnCObFhrFH9uf3Bt
NjHcjYqT0L4Wpg5mDfYILhnLQ9yGyemZuN2eb2qghMmTgYf2vdFow+SCcy9gFeKetNV0BfMLagns
2CF1cCePECX2Jxci1WbFG92tlSLVynAuBoFCTqMh2tp+wLyEKSgvPgK4hwXn3vqOqEWTbYMOYpn2
tySA2tDM5baGaakFflG8npTBRIchEddDFAO6CL70TeagkT9+D9KbUk0TyISzil+r8LjTOmEwbLyG
5EySYFLqJtqMAVAy+PAfGYatDaU75f4wk6ELDKMWGefpHAupRrow2atCMthhWKzaykkS5U8Jpf2N
tKfFCF10T/b1YwDqdC8gQ64ewtQBfOuyK943D8aWJHC2Po+Gl209e+rFr5vkGh3nZYyhnCq8RGXQ
dDbzqIEbftx7msPeVJK8ZpM3hyXr77yb1qQa0cDC3zfWWfVlPFvvAmKHNp8oA8kaLVPnFDs9C690
H1jAq10/HY7Id+H9iMXRLR2jj38BpdkxyfNjDDTFtGuZrb8EwrUJwKrmGYXEmypY2GT79pWuQtQ2
7Xpcyy/JGygnLXqkNl1izI7n/dFlPHmT7NQ7gEMA6cwbBBRVY8mp7beVFE7f2koFvpqHvlvYBeQB
vX0TomoWZV+SAwDIZItZXyG/nNBQZ4GOL5g29iAGRD9KX3Mp6Z7BI5Dr4Jsa1m2RlCSlQz9G/vKS
RAq+t2ZX4f9MKcKmh+lvV2StyN7cpZ3m0cHDMmV/ldBajTeXozJf31P4gvef3tNV+oQOa2vosI3C
pSUdNBH5P+Yww5X+VRuq5vb9rTKmWWCUJEXbhDhAH7t0sinUIB53/47CZrrsKvjtrSGcgHXsCWny
K3yfeTfjC65CCms65/FsM3+5XyuhUET/I+8dFhpI1kZnZ9OR7jE5P8rmdbR+4BwJ4P80/1GLYZfW
f2xAP/anhm0IPvJKx4P9tgyCEkFpuQumEtBejrFzeEVKo9M8TXWzNFMTYk/cvP79PXXc2uUu0bHw
2jBOJGE2Em4T5clDPyfs8KzyQ7KNM6I8QOqcmg4PtWkjNKH3tBSBmqHbGTFtTKdmHCDGpDNAxK/C
6PZ+uVppEIojh4GvMmJO11mBuFbfY/H9kbH6EQmrYTdUmSA3SYEVV2t4QPxPmipIOSALuy1QSXGy
yG3mHPaiFeNaxmSP460Ta2XToXFL1jtylrDlqIj032WrLOjxPgsDobaTPSoflj2NYITQScHOpDLC
6gXORj2vcyKtIE/KpXIDofVv/YSUzMlM2owCFveptxwUjVdYkdTbTqc2QRzYBTLPZwVlqi2qVZA2
N7qHT1/64ON7cdntbTnjgjE2KLVjKStXqgT1MQTF/Y6m0YD1NxrzmMZIpjfB+yttJRAtPwTlR9y/
K093B4QnCgUpf4Osvx/wHniBToEur9K5ly6JE92h+8J3NvVdZz+afUVHkMDLVlcMpou3QgjsYdQ6
iE3g6ibBifeyjaM1ZIjv9LdBZMq+AVEoBUfIIjUdLL696VbnxEGH6+j4hPWydGaO8vfmvkVS8bEQ
bKAXsUzHLk8SeO5hr9QdsK1sAEW4RnzfhGPNYDm8/SgOcFmfv/LpuDajNoR+lpyaf/zcJXFiRjmi
XMpRF3sHRmn1z0wEsflH4Q5sp5vEOKlVsRZEaZFmPGclmp1Rgptfm3I5zdWDJZo6QR0mmxfCnNFr
zuVYwnuwueqVxwKGSzGpViIzUTtiJh2l9DKdWA0Ht9fsEmHwfZREOTUJ4XyBBo81FST8TUo56V+4
Nxxrg968WuX5osLQJ0dPxX053NxT36ba5FEtO+FQfoZYBnV4obrFeDlOAQy3k+9GM5/MaU5Z7u+7
HRuJGiRH/UPDAzpYyXFrsFm8AqiRW96v1f8ZKipkCMZwMU4R1sG6dS0JJUXBjPL+on34mo+QH+PG
WZdCwszkxlg27bL5BxblisD28v9ZZimM1e3L25LDLyuffJ2APhj+bK4Agpa17Mi51O+dc0CDvykg
g5kcZidLg4mCCfxVZHchgOIbsamXQw/E6nnEuq4oNLFCuI/9LmYPALH7R3dBn12NnXil07jgS8wp
RD0qnjFFjnO29k8h16/LceoVW2sd+PBoqb9MjgdV/rZJ61+qWxUST9to2Ns1FbcpVPoIGDRXFRYl
km5fDNVkZdJ5n4zAi0+TJOkVe/K86doB3j77IA+xNSa9Bt1CSw/7La5Yg7NPvre48XKmulNLoWUE
5qcdg6lO0YBWet9yuG/bFEyj1Ha9oKidchjIm+pZFRUAgEKRf84MUpSEqAualbMrzKJotqzHnE+e
9bgszZzVvii2xP8FPCgo9+PVNxqKWGJRUU17p3ergxyeIfkLzq08/laGSaaU0hCIIglKH/ahgfON
l3YL8PVNkp/UMsoftA1oCmPSFbDpgn9KDIdmxVSy0y6cJC2JY24XZJLwTImny9tF8Mv56fThTHtb
aAt1DIrTn4iAqS1LEhkCZ2BOKG7h29y7PUwb51yJmWMdizWBtbR+MQiiJjAsBtJ4wRgWzc3gLsvc
JMKUgjGkK9v441a2TrAkykLCh6TqKqRYnIlDm16gMC08QGjxeXT5Mm3CYLPc6SB1EulYDgi6iCrH
mToJhD8SvHXxwjm6kzkPd3KtEsMXKJrraWZaQvK038HwszXQyEhvu7RetJyRr0kZEXK7AP2XDKpJ
4dOmqyyZJor3fLPw3wNS2gyqFXslnMZ/d91guTfUMNwU56LM5IPrV3kSxqAgK/qacX4qoMduXud9
4JSzheT+gzI9IGyYBvLlIAm9bydVn6cmd/FNbUpcuaQ0ECWFH3DNM5l65oJTjcPCP6s6A4xUOjml
ZnbRgOKoB4NXb3HxYFI8uy4iG5on7nlJ2qgfkvuiZGIkAeFgGv1E1EkB9XR2Bhhd1meCH4ecaQOH
eBGj/jIm6WWYGhkAxUx0oGn4gdlf4vC7Zr2z3SB2l59QEXK6+XtVj8GkDaKMsCsyH/2G8gxfDE9N
TLiYD51A0d4dOq5HdXuJlq7rAZAWRRJxyVwVaPQWhSi19N0w7wpms3LFxj8V9EJ37mo0lEIHac8M
i0Ja4+peVAf9/nzisDZ7GPnBnYweptPrbs4RW2QWeRSEF7zVmoGq++PEkYei+G7FUO5ZBkifQi73
yTuL1i2jahdYSjrOQj5GLbxbDyOzeRN+j/svnD56k90LfXAwnufiAOu5E/sKdrXoUkt5wkxb3H36
wyArqXIBVoPDfOgbz4ipC2hMsq5Q+89msvKxPz+syq31EXeGtKN3kvDYsRNpCmHMd9oiCk0wQsl+
ZdK4Id8B/cUFlI3Lcl9/Pd95x3q1Nrtl5d+WtiqHrTyWaFBNEssDKnKsznY1/zMMT62//EJvBD/f
TUJ4G+3rVnCjIQwDqJRpj+yFXgg0ubKXqD9SmA7jB+JWzNvB6AYdalIi+60JYEJ7oL0+R1MSNXHA
5rt14//Tanzil/Wkl57xx59xVxBgJMAK/gIT21dXUAIzBsqQ+AD6QJ9TPftVt6cswRpfCbFT2p2p
fEfcKQ9pZb+znWpCyEEmCwerITWaIUpg7OJe/eXWeO6lNZc17VSehkj0vo9+zGGPlnuQ6lWAAo6Z
z2MgFEnEV67GSufxUqft7Mgr5+OHFybZzzmj/lrIktCIrfXeIxuxfJXk/P0En0Wn0mjWx4QeJJGX
CeqguxCDR6wjDhQ8hi5reUq1WOD/hHfrLQf7DQiV8IsbZ+2mSDSe34mjr3pR3Z0fM5zdZb8b3D0+
tbDBPyaLT5Y5C7c4s+9/731/YBmfjJoRaVcjsSneNy5U+AzgVGizouyNfzHXca/yWAWMxYyqGyCd
eWNkEYVPxkO2ha/fIg7sb/RWj4LtSz8kle6FumIxbKQPSA38aVRkmO81hWP3tH+JVXLo4GONmM2/
sTXaJ65ITGKZFid4qTAyQEGlFdhZ/VcaW//lCV8skk2Iw9PTY0KLYYafUzhPIbXsmO1ntwoQra6L
U35eo6LcgmCHTv6WPitzm2X1oHu5GPw5qjdlJP4BHGCqL0/FEYGifckTA8NOwHgacmVgXdFh5xFi
1zh+EuYHeXJ6kM0uSlU1D/n0M3AKpzfBvITzJ0bArmGC+/gw174HspHjl2tEcW3kYRWpWG/JMhvx
HH7EDXcapOx9Rj1gkidhjWvesdIw2MfmBo+FK8byeLwvgo6NcQWfjBlhguemDH2iJztCwlABSKbi
uRNMPuYQjLfWdHavo+6WO+Iv4frd0QVPiB7/+P33SbStXStGD0iAxbwQmOxOG0Ts4hhnm/VYMpbu
7X/C2PNS8TAeTq2KWzrxq+kevArb52CGKR3Ykl6hLoUdrAidIcdAtYqBktMaYcNMVrJE7AItLuo4
+o0xeFYvk2Rk/xPVePZ01rOQ9cBwpMjQUcB5MIdP61s6oqbbaSi3WDWtJGLjgmaKWKRins5WvUZf
SOM4F7XxC8p2Sjb6RKGIPSYk4LKft+jCkdQesBy2MTnpYgePWjSlHl5qNVq+eD7pBjCp6Mmnm9Af
DyMGpqjh8aA9q6UzKZRYED9kFuEy0zCZMbY1TY+cW8ND6LpJ+AOZXIsWCOG25LfoOmcJQr3IiB3Q
HeBDtfpgu8t4/3Z+8zfNjBVN0GidiLDBE2iZQbSPbHEHmXHlZxzvn0aXDFkCoB1MJyAO6M1xV+2I
CkgwbXYyddnvMuLwmYHb7Mim6qBb2X3MG9IdJrtVNAAsII+8IAPtHZXkk+tUQ30+n6W1vxY0lTo2
PXxCdDp+gZCjWbwDm4VDlXJpWBT/UDZ1S3dXQo6QKQm4mZjIdNVYcBIZEC82f7wqf0OD+a3uqxGb
QdtWHPWunV4fxfQ3NK68BiLsCnMAbSF3jnkJkTHk/zfoZtdTl1toqvM8TxOqGrVknuhVl81FWXVq
Usz8ywb/WmR3/ci1NYPV2qQJMsLQ0y4m0LuLPPPICSt1ggGsYV4y39NcMM6ui7lpNydWQp0DMplL
8SsouK0D9VGmaHeLBIdcHdi3KkVuQGFCPdbiPHToOvLswsiiaddsVPREqlBrGuC/8CpHdapN9PRT
3qOOkdsOH9bGFOmI80+yEGFB+znRY08qhwA+mzz6VTjEEbQ0oA9fn2o8mHJ50Z7Pf6sIl6O6+pLy
ILsDRZv2IWpWt2/ifbekCrygJHetlQlDCZIYEviDs7fm192Nqyzx89vpZBn9KAEQGZac26K2jpHz
ncbg8MVSA5AEW6pHQ45CSuGtZft/NFaiBgFIMTyDN4iqr80jzWuDI6J8cJtwviWl4eftvZoa+MMd
zPen+httXwNp22w2Ad6QA6tBNE7HI9QIAqBqa2nDdyj6pF6HytfKaiYfLGl42ha3F1EfnhXUDWES
b4xjqY7MXycoXs6nRWVMlzb2eFJUkti/1b8xOwDi3t5wob4NEQ8xk4kKIF+0E/xWqDMLZaLnx150
TypHGWUvBDz7Gx17P2AtIgDOJ/vB3HjR+WJ5yot84DuaOAboCdrFYtTrQFjNieFTHjX0P8aZ83XV
9GHyeeRvcTKTelhv+0BKQgGPeA/ZDFFz+G5iRJzTePaUNgYkXdoaG660i7XJnvVaCr+SLVk/+52b
GABHNRAymbP7MjuSsPiG9eEOwDSZb8kEWTOhmG+B08ZtuTirqwydGRYHGjssu0O/nguhIJ36op/A
9cjte60qLovYXmSM4KK1oNGTDHnVJoo/AluAEI3/3Qk9zOmOEo5HOmZsCl22fMgCpqyO2esuoXCx
jdBUtguZ4Rcus6k5TKgn7MYhXoTRlTqn8AitciVFJNK2h/tTe3z4SMNt2rqyPoukRhqp0t9j5rUf
NKQ22GwZ0PT7+PjOwNapxvU5qmSM+HGNlw6T0akvIyoeqhAeWKQmuRw1yfZcYSFVPvyHiGKoQMKK
1dSSNCUR+p5JNOkpisfYLC65QCMKJ+tFzYVztB5/8f4STajPLxQCEX05eOleLHThBHpUCkTDU7cb
7uBgqoh67t5yTzkZJr3shArcq65K49MZhUUHPJLM+ThuL5h+vvGsdKyOtfvNkgigBHjbJiW0ak1Z
piIl55BHP+jNUsw1yVzNHTbOHFfN4K3SZuT6zAhnTg6Qg6/p3JFzZFFriQD7Ym0KkBAF3SAhs4xf
D+ViW08wKw2Isp8nncu6OTPGnf9IM2SO4zsp2JhwKjSgNcLsAWbW5qg4nWNap0L+2h5nnamtwdKy
hjArePHaa8eDguELJS+fnJT6gThzHCyqSq0NV3EyDIoyruzHT76f6ZQ+tdx2/ZvsvwzHqAtO0Av2
KAmU0r/k1/J6KqJ8e9OXT42avH2oJPtzF9VXy5H+6ktgNIQPSr4FNanZisEmDupd1AOQzi4UjUwk
lTwaHOPMDaarWnAmYf3pT+ewfBArNyL4eH9Qq2DYWPfls/ficJtg1UttHjKD5S34VOtcRMU3St4l
vhaxXXiW9KpbcVXj89fhCXqprv2rvWzCeM0C954kDr1lE53SBgoWtMC5bLRwkhDOTqkIiWljs0W4
X3ViCtWIqZYf0Jho8bvtU2uE0apk76o7v/DxBdMa5o3TYlGyAy7+3BpdIoIM5Q6MgbGTnKn6bUy8
xxRDPIFiDW6eDga8A2UIzUWEoHGBnBf6v+T4U3VQ0l5XPAF3mH4d+LGAhckjtpj1N0CsCwo6+fd0
Z8K5qDPlBUUsX4KmDgz8/RuEsiHuDc7y230/l1VTaftVRkOMvOO17Mke+i6k0m2Vb3G2iVjerZJa
GnhM7qPs2i+p2oaelbOlD15uY0JqcRTMsA2Zyzk+kIjAGLQkKbt5FOvvYd5k1NVK3UMZaH6Kvxs9
0GKuISC/lzp+XHpNBIBPQm97iMT9r+ooSaqx/604PYk/ECPzyIu3oRWLAt5+xez3FVlqfpuuGNSn
MgPQPw37UMogcn0Od4RGKT/QVCk2EmgJn0JnjIaouhmEjFmXfYhS6e0lFG4QFXFY2MaPFeHN9l5i
jiphTXqJSPKk6McxevirEuRHboGlG1ZJglEqlwZPTtiVxHK0AJnUXAATf6mWMPTFKqjTTTEJomFC
cHGxTF0S8QHTawkJLmslCl79/DUQ0jCuCQZ1bk5AV0HQiak3iiQpAKBAZ1mMaxvIoqeQwZwQaSy6
uhXh7ntAC6mtFxsnjmUbRVrebp9hOjqSXjOmrzSqEbOB0o486UmxH5Jau3RqBVSBupyGwUtdsF2R
jdkOQULCjCNYR9Hnpbd9eL3whvXtza9O2/9NsSticXy8uA3c5QdDBuBBjxfyh6hG2FNuHunMrMoj
Q4C/zxq6zAUsgXUARjQV3xSXrV3uQdrDGaXcy//amWMCQ203b9nD0lYgd0CzoQqUQBIVFhohh4Eb
aUzHxIvl/S5xjlqvYtIz51A5u3XRYN7svAEr2dIGrvFilMJti2fao548Ljxyxp3bQw2bZZ8KcS8A
q5EBZDYobStGedZ+LZXJ2TEfUbzhIXBCBE/QElyFTwMd8WnwDCtg8pAv4Qi4jujIbt89kaFQIdNt
ckfaEiSJGToNET5WPXHBJ3nGhffb1U+ZwzXhj6qFw8FeCcO892zz0mUFOteMcpEhCEJiuDGOGjld
t4wU5oP/R+lXe1mTN+40o6e0nrnPwz2X9hu2ewbT74gBQiE1+XqDbVIYopyGqS0w4FdH8OGMjJXk
s0QIt4eEuCm58S6rKoaUGkRW3xGCF0RdAyM2nki8JIpLmDLG6rzMBfg44gFNhGNHoffl+d6YBzDL
VsTAG1+gf532wkGil4IizcyAzf5kQM8eVAcYMlpEzZE+M8WBEtL+jrNEpx0KXevLKbD++h1xdcfX
pJbDCkEFVVbAILV4SgoLO1IHtzi10w7jYOTzU/rpw3K4XuJvh95Yb8mknMpklZW3SBTTY6SewqKY
JX+kwnqbrZVdP07IcGs9PCOb4azYOyfBKmyUF3WxxgEg++d77DPJ2Mygw6vSolrHesJtlnvCgVp1
lnJPrL0sQIcWlr9ifwOufSu5ONCXzMEYPG4JJfXKFxpGH3DlKuXFFzY84QwvnBnJ2bvR6pXEsid2
qRH/UR+ueG10XtJz/MoAW39/whHOL4DJy46ZM33FspQyBGC5G6AbNnVkQ7+7Awi5/DWfzxV4eScF
lAnDFPa58jZh3PH6eo+ilB+Ixq02toIOdPfDntXKCYFBLYbRxMYp+skNmSGbD5myupb6FL79P+/w
3PCdcKfuX21p6I0EmSlo3EfpcI++qfFMCsdPo388yp6odiaQoOhZmTgAMhXFncccULFWfyoDb+p0
e7M58oJED8KT4uqMLwX6YOgMeIwl7osnyPYv7juX6lu3QxWhot6y4OacgdE9CxO4H3KTaCPZSn5l
S9LE/eXrWGktI8W3vNg4nrym1G+YevGcBsK9vJgqTJ/tuWkQD/yXDC5nFwUABWAgWNBHOU3SV/R+
p35000FmHTiNlw9AGQghX6sDgZrgrplLasw7YbMDKFKCaxL4AmbeM95DSQxtSEt4tdHnCY532XeW
Sgvt+JgdyEKlWeUdxADntc6QEVifCWqQjCEOWINWvZt2mEADrIGIH7UVBBu1R18RULiOlspCkaCM
SsPbK+vCRtY1Q1CeaGp5OA8H/tC6ZtFJcKMFmv6NGGxfmkHr3mFdU0DDbiX7yyRbyYicf2XOUSrI
xvEVon63r7B2FTGzuEVDQSq6BZTVTDLzORN9LWk5MdxtB2qTU4bPsfZ68XMtSJj+l+Vg6QXlEsqX
p57AQoeqXdsCbhmTfmYc8O7k1xVosvZmCKLwnyBFqv905afRSDAhdic1i6zhS0DGPmAt2LmigAoF
DkAlPRuHVOGDLp0iFHVDPZF26RqVU0OUdCf2QATt/68p0BsIBsmaOPp/SNEztfUr15jt+uL8gVpJ
ctRcB10/agJ4iP37maAjhnSE26RCV0qKJNRjp5tTIAHrOkWBtQWuydNAzKGUj8zmCK8i55AWGwqF
04OodTI88LbiROt5ysYumJ0M0J0bx/lrdnzDqN6nNua/K06p/p/zrB8/EZ7Gh7MZnOxuMRTFPUSl
Ulopem/3uiYiVzj9HxFwGGiDthHvLlFSG/4I6o2d4bC128PwdvhnQhrteXjFUJWwMHSby4ZMAqKA
w/vsbnEZ7149jKK3QWTwuUJteXhvie5YEiu8EZWuRc4cBPLxNbGym9W8ln6IJL/oPjV/AO06Nifm
5571skpvKwkKih+yQIDeQEaH6DWvSbesWFTAfiiyUHvoSbLpx5NZBMjDYfdUSUXQT4FbBR/gdyjR
y1KUHNSaXya35DV0v6kYg9sA6gIAq3+ma6XgQmtlDROSdzUfl3D5635Tzw29aLBelxtj0BlCcpH8
9KkhC/yPxSQ47hq3YJMFSpn+kg2ucendpT/GehOMth0YnGW7G0VWepPRTd87U4/23b5/SnFsD8/x
p8PSlVaCfVaGamqdcyUFSS0bWnUDXbsI7jF8dejCcwKoCa4UP9jvLrwDDEejFSMW4al7u/5hD1lZ
08Wu9TTqb4rNmtT+wn38gXN1mYRoKW8ty5WGEWQv6ajQaomT8/990k7KP/XVO6RUzd2ul98ZD11O
y2aiiczge44qNx+KkXnKQpmvEbgo/H+vgXNiKlqyEYI0pihpLqOyDvWauih9NEzQS9OTm5skCFGI
AITVAA8wKQmW+A7PD4UP2/4wf6HLYyJ2IQGu8emHxXaYSa7yLUY8byK0TElpnpkCpmPh+r8bkUVL
0CDWm+wyxGz1i1mEuJviLc27v4rOTHhmV5PUh7VB77kn7Vpp4drWPfoVS+A0+/TfHv/cRwzOL05H
uZK8cogZWiAB+6FNDVr29FtTYKNu3PxQX+lfw/QJ3ox+IzAjv/J3lXBj9mjrygHYkFpnnKldfr9x
pLnZ+pWpgansoNOmczjzpUwRUfH3vzev+a09EyhFcyCN31RWbQW4Y3KeN/UkfJ/XbmmnLp0MFjZw
YE1m7gTPS5eIIXus9NA1jvJOK5QgT7WMSfLdCEC5rkeUfgSfsvLjpl8iKmkc1eVnIdVb04LFH2MW
WlGqgpKZwv+LTNc1x9lr6oe405UaHmyODE3eCW6AyXd7UwNYeb+2rC2moNE5/KHl/2xVzIvYX/9k
pWxxRfKAul7pdHsqqav8Ow8ltLDuSSH93BTFBy/eCj3g1bjYM/yuYSuFPv7iBsFIH7mDlCuBQuOE
aNjB1vZtZsMcOlePzUKhvYYVK4HGEPL4WkuNaJsgVFowwI09xkrCnEajiJkLWFe18uc6Dxp/00Zs
DOF3T8BZpA8naxA0BII8Tk62OiBDE20osSoUYKj2LqA/mpKdcSisqsMysGWGYEBDJGxbKqyghzve
xIGrHCk9Rbft9pTntAIgwboxqSTYD3fExS5G5KzmtX20AsR2BWLPmhcvpO/JukNxr7qoAk8FpPRk
QrRlcxps6EI4u142xEahzU/gIKgB4iFDFAyaxr4Nf/7OEZ0bP1dDC6mChjLdYqgrficBEe96TKbC
4rI1XPO6WL5sBKxCCzEGpnP0XaQRHhbrZAAF1mYyvtacDmGe5rnbdnsk8F1pQdL+bdfSW7ol4jvk
AJpTEAQ0PqoaTtLbOQ0aUTW3NXpuu2Mke+rv3XrCXb17OLJUlD4WyQuX8fgXXIQK0jUktHw74DZz
oRk8hrlTPE0O+zj+zzuM7jLa2kobXSVSFh8+kfy/zgKgrtq/Mb1Dklf6jzvZqe1JZ8RFX1jEJyB+
NNOocvP4RPHaMxzfG+8g5z7ht2gXFqrLX0DotAwB+Gr51/CQMtUhQX4bpfHL2sBUQrszdkg8Ek35
VbVQyCkpTqGH0YDN0bboLMcRK2tJmVdYQEZqIyh0E6rnvCj71GZJ5uKYYsg1gIxB6au9xoeD1kQm
QUrTerpdgF8FZcNWAyQI3Ytox1jLvN/30qmbDfpOM2RLcDXtMF3aDGzlPUaPvSv6YyLuY1Sz0IFu
szMjDreWKSWfhS06edtuXd7VqACKrQPv/UVuL9jT9gJiXaMIFQrtAqMehkLvfD8XDMKNHI0hLKpF
3tipY4tm10NeUIe7yM4dgG63/6NTP3JOhF0qFeUdxDqKb4pezthDOdYtgBVGxrU8sRpnYHN/vmTc
uiWOBNK8M/2ujPJWQD+r28Yqhw3Yzc8eWC5C6HwWKhFz/xGKf7nkR4Fvol4kzF9gliYrQFi2d00k
0jtVJmZDrUy1lZTM1xZtCxhUD7eTQzS6vPSytbjsg4kKjcd+ZZb3WDI1MCOPDt4NwUUzpX1sNjfF
D8mpb46AcIB/rkYzO91PR7jCXbWL47yPylwPtj7rRBSfB3Nd1RaJwXHtsp7UqUyuDwPTb95TXlZj
0vsInQNZ4zmiWsZKDXLUWTPD4IzReIxz5Gttyn1+gzx0NWhJSe4wrHPClkdnpZw8M0M2QOwARwNp
G9Hkq5kVbRhamH6tq0nYseVc8Qgy+Drdvx/AXDA4DEvv/x5jg1rmVbdDHFJIFhET0ZA4YYuDaWLe
xHtFP+GvpkJD0Y2Ds7V+FgONVMhJ2DVYnNuBw/CIBTchLop0EbtLWfNrWLq7BRQfW9X3iQUbg1xY
HlmslSdaXBMJ762i/3c8fPQo3Le//OaG3G1tHfGEMthoVe0Kfnqqde6C12B3SUKzm6rVwcQU0F43
zwerwSCXBrsqVI1TR2MBzsAGhsJDVDy+/smUJXDtW0U7RKvo85SEdyRM47eOVrvl9sAIjCUS1fQi
bJBFsfzZpc9ujovESt7zC9EPXrDFj92xqvleuyOYdZW8MqcyTCAMjJbtMaFj1Uqiysb0fNjESRI/
Y+xhjrXGD7LRmuDSaMpussOtnNc26nWd2rCbpuMHmM8ARynJ5LwZd04kji54VrQllPnI4OoVrRus
tvX6V7IADjDLtuZOGFbXDc2F79meby7xJDNr6fKchyYBHcP0L7XWRMxLe2RLhELjvHDKB9qjohl7
Jkb72bomXIAL+cvxYOFhqbKJZ+ennUpvhW+hoZHZ5JsillfHH2u0QE+wrQeIA/x0ZsLhEkrx7NyL
uXGQI7z+jaL32RuPjf1e9Batnq2jW/8X3E/3kuSuZl+FAn/myP5ETdN6Qb9awARXbZYlG3B78Nhu
qIxLGv23T6MiHLwYxh4bR4SDIcE58GcrZCST/kV1AE5O3K9BkMz99bHlKHa+yEX3j2JXV5ZWYHvh
sxxL3gK1zsMrk7k/iFt4noNeBIICe704aAcLTZuT1Shtf2s20xpx+40+V+qUpPSjI5g/UTVzcsEU
IowgQfq9aBG0aWGSLN18tadAnKdB/xYVpf76PMDbpEg61DIjjSEJHD1azmam5KQyHutwqN89r4iN
qZkomimVKeHfDjY/VXvuKsx9hgDEAvUOrejjafWoxaf5Oyc5UWmlHEv0XTE4iaoO2+5/boIEqpRC
rbYwWEO4Jj/FbWpbbQpb4xZsdPynh6wFlD8121oE02KHQO0/EJzhzDsiFpeU6htgxUaoXvhlPo66
uvhQY2iqn5uflmGDZQFFAaQmdkjipcFw980cfoPU3FvesQIVIGeUunRYwjBf6M3eLoWs3sCaSZpC
KgletE6WXbmV7V7UOqf9yI3K+Rz+uq/2WItYyAOVO4WfXsQhpz3QJuY20OUftARcfSi9DYvB6sx2
YJPWPQtV2xMRlJaK3xuOfHPC7wdp5u8H1DRlACrc70VT8GMp2e0/fRwPQuB7+jrJvC8cp+2c4dRX
i8Jzj0+pqOkB0ZnANMRixmNw01wQYG0ZoE5XXvep8P3ZvYvlb/bMq5JE7ZATQk7goUcs2aGlvLem
eb20uKkKI9e1lMGDuIkJKbFQ0xUVdjo/tCxnE5HkXgrNaN74ROXwdg9aGg4TMvbCrnqnZjsGeGVD
ilYANKkDZbh51R3vw9q/irzZpmpCGR5fMKbEQatKCD5BpRrobgOBR5fJINOSj4rQfJ80AUH1sw8v
/ExAnU/dcXDFKUaTIO3rkSG4qhjNIDoSOgb6ovkO1ay0WXvA7aG8gdTXyRk12db9G3jSCrjgTvZY
jJjaemlU9ZSvxzXkJE+MN7Z06+poWk3wsFEwHh7SJV8WTmjtsw6LTu5CvpyV1bty2Zwfx52D6iJn
wPa5Br4BAO+SQ7g5Dq/DxfAvP5LGKR+Wf8ymq5Dj6sajPzAAZB1EEh8HfcPcvkK54UU3j2eLlKoY
CLnytN0cxwjWFR5T9YtZjpEIqlG/b4H+IUYlYSFRHSU4id94SNoWhuOxuL2eyuG+ktusjjQeQisB
wt7C4gej6t0tolSOYCP9KVuycZhnasGUNvnFkBuUG4SxqrvShhQZ0sTREOXTmHZxNgUeU0sUYhQT
dzgFetqcU1LykfbjcHF3iC6t3oPXY0Sb6rWHHKe3OSZr0ehF7CkPOj27NOlLSEGtdQOwhVHA9gv8
FDgEU2lo/8gpla5JeNinSzLhFDtzY4XJ58xryeh8zHjJk3MQHkFWkpa6JDblDIESaRMcEPfZh5Eh
N3Z9gYXhCKtH7P0kLpX6TGWjhffBA9Oq3Sl3cGUEInwwGK3ms0TyNCal/TxltJyYVeMUZSPuEche
iDdGn0TP/+chB6cHktM3/zNBQpkFa38GpiPQTCagWHeKuJK1b4cpo/buITwfNZk0e8c+x72pRswI
KyhLBklT0VUEoAOr8ZgBfT+VlSrqKASYL/RLOXj9r6w/QNHAsar+9pfsNupGXQ8za0YqPTJHC8F2
JD1QdfJbM8KZO2i71Fk0TG3CAqcyjsw68CpHzUynspKyXU8g1Tb/erPvzLxnBa4JdQtED4QgDAJB
ltSPRvhJUP1TgsOpnRkVHPP/NBbtXIVm/u5lD/CMSpvMSb7F/GhOxerQFcoK1Gz1OI17Dk9scwp6
nwidhbfusS8clwjX5BiRtT1AfoPPtaYsDLWjD2tXLJ+b8k0iLp+J/uRSx+05ITfZrGBw7wQDX3uE
qgoNjyOkoycLper33a69YcsjE6dt7/tILTsr9HFBc1mACZwuFKdLnwoRM1BDhn1CozbHs4Ch2MOI
OMRLeosMQDzhfBSbTXYNFpvF+vbFYJ7fKmqNrGb5+oJL1N65ExsYzV60AUQvUG++g8+dn8b9S6sa
19/Jr+GH4nYL8J2ShgIhTggZxm60/+H2fT5VTuW7RpSzvjU8c2LHJvRaNqRfIjIXy3w7RQcYa/Fm
nus6iQQM3gQE8x18TNdddtNFHw/bsTk0r3Z0Hyfjl5nETPoNXEvodgfiC0U2JXC9JmlxNlNc3mVp
lz589KA+PrjIjXuQhiUVASBJVP9QZ428XPH7d06OdfwAlIyzQvzz02OyoIBp5lMNn/ahjqT11N/H
V1Ege54OLY5NbJZkuiOEPbiOm6WznX3ISqlePmcO2Sq5k5oNNZBKSnxF9Qzg0XlibQrC1IUTUL7U
W2xJ1MKd4z9MBJX6wS2VAuQgzRBL1u4dYY+nGf/geakFSpsEgdOv3gGr/OVsXDZ9ysJsytoqIZBm
PxHVXe6n52EAr4kI6/8Ys7vVgt7Put5U89TWO0q9sgyhoxd/+vGH9sPLw8xUEsKg0gqCsz+eDt+f
lQBA2Ql7y+Thk+m9XiwXFyKlLbTeaBgvH5rT7JfY52tfGIipcoExvAUiqjxmU6m70RTSOOgIp7kk
Psa9IimZrPRZ+mTeUdXbz/FYmCHNDE9x5WcHpjvr4P1SzIDfSD+8qLDayMdnfu6KH0pKUpL8AECJ
GMyaZdMPQNPMPj4KgPTJ+z2/vyoFqcBfeQEdOX0FZvZLm7u9SmTwtkhu4FSdjKL8ehnZhQSVgpPP
wOHv1jJ5mAP6GyAJefJE1qpK3vgbW6nOHpEhJuNgo9CwrhvZ5ORMYCkPXiBkN5ef8yHn9RK7plfH
Cft/LtfiTiKUdVrZYWiMHXfhwlg4JYN8Qk7ouWl6PlnmPZ88JJSpyy28XK1ITGEM60oTk7nSd6ms
kgFRa+HTtb/vOu90WFE5dAr4uRoODnb6yQ+IuYWyS/4CZXDQ+a81MCOhS57qyXhSF0VWgaaW4Alf
8dXzD/Q+wq9TZE1rwgs/dAaZ0n5whiiD3gBAzKjznhGQqXbSDlPPjVoHL70rXTyFIA30GpAeWmqB
kIoGVEfhpi85quL11MAoVzcZhpP3EWUEcUCJRlnojfjk/yYpucr9aRntpgbkRZlnRYf8SucOGdql
B0FsZoi8n6uTlcBMENYEnxmchkTxgSOVuNP8veCE/x5ULsZE6Fjjpg2C7+BQQro1heZwykjy0gr5
q4Lab9TjoTPmP0r1gemu48UCLR9Y2FiY++zd8+NKB49gqk0KHito6XSMJ+d3Uh8CRuRjbYEmEasB
0miDkNUtC+7Rcwb68BcDIcoiX7OmYB/Az0hCY14kp+bry2Nss6gL3k8BLSc+8+T+pnSXqqY+W4Ei
QZhA+bsMcXGQefVJrGYv5K/GJQOijUuefwYmTHeyNpb5HzBAlwE+UFt2aPHflJZUsdeQ3sUMx+RW
eixekTUCBgmMFW64picAh8oI8FmoUh1SxYNCjSo+YsXQ15NgEVRJh3eWRacNlUEdBb700+40WYlF
T6mJ2TKGF9g1bHi8J8sD/184q/d9Z/PoAc7aXq5dO3nrI/QSDCsUavplclOvdHGB/N6pupd26E2V
uQVGQjIY2TeUwCoG41SJMuhXRP1TZpNYs4rSHZNsPWS/hEQZGabwxPn9kqDlEChFb/MztEsCja86
giIRWAXISTKAiTUnORLRPRAMg7vj9wudiWLBGcrafqMBRMSUH+92YGOxGarS+fUsKK7bjMSSFE9N
xuz7Bvv1gDAPkn3QJz/LcSjI4JyBrZLTBXe5GNoTy4aO9/mCydQLt3k20mHaLuNtW7uuCxHIhjyd
+cqTaAnUMhi36r8a28RybDFxUdKx3uJDsxMX1b1u6sMbtaLaNNLE5WmZ/PSpMHLP9IpvSJ2CgZh3
o7N0FKspW1EmENjW6HsVRL0FTxjjKql3jWhHQ5knL7WeEmbmG1hzcVqZfZbr9FNLXoHKhdAnzJyG
j2F8CZVdIe7f1Tq4b2n67q7XcZTg1oNK8A46RZdo9EpCSN9NjrzB8bIadliG4jwRan0mJI2CfRa4
7Jtk1Zc5rR+Jcf2bKK7/zOjVxR70BQPQ5jqsPE+siGuv1/8Xwdddjr30PUEhqFfCp7wP9ch0YHow
sUmRCX39Sq85i0twGCPG0IeQw1+mOUX7jnHPC+/AHUQDhxLVU5lKs+ejKldDMFwePnmQ94z9qyXw
JuTepitQ526orRSO3fmXoMbS1H6/TGhSnfiP5KGqXLZXt/okjrKMR7dvl9hv9Br/PKP5HtiSivX8
ihWek8hUXaOjPNYg6yPr3dzV3PEPc0pfPu6RXLlV5McaxA1fTiHgmGqttb1m3a2cxfmJG5uAeQ1d
Ki6LDlB6FQU99sTpq8ga7EwBVO7X6FwO9w7Z9F67+HGsXRYUG/qRDML23l474VN03pSUWXuWXQVJ
Z9Wf4QfN3TbHDWMHOrQkEt0OS3oZO3Fiqpko5/knWRwyQmTOs0d5PTduZ2AYVLRZ0oyfvI0pKp2b
e9TNnSmxEbB9vQ+dPgWDgV8MBao/1iETmbsWzlnOa4AUQfNTZrtpvfxZ4Srr8o243tTygEFKf8uI
Q+kRge3ND77b1uIv8hF6CVliZ7gahO8Mln73riiNF46HECH7rsycUOb5d07vergPgaLsw5GNz70x
WQVkCRFOYpYVy0vxqKKJJehaev7RBbWLspf81i5FcOYn28o4m+HM9HIOY7qM1d5l767kqC/3cjzS
wW+YFjfCXQ9d1+SeEx06MHb67Co/s0SArLNfPkMTBxnaEI5DE2dYQMJwwrRWfeA2ewttUjpoUMZi
F4BWdeQhaTp4l6uVM35vXcCZb49lSKKY5f7rLfJpZVZpTsXvIrYJPAC42aJ73TCixUU+vjuynKlH
S4Zk15slecyy3iIUXZshRvaAXunLLcvbsKUkPgj0nO0Gp+mJdJCkGQOhYaE522vi/SmqROiJr7Vw
dF2a3owWEpdPmiwG6MNwEUYKSL5nu3tYpr86TnuvB7wUoHx4xMJcLyP1cCwXiks6TadrIWtTTU3h
1TGg+5VFGzq4sLEH76Qvo28N4E8hRE7kMgmDiMCN5RRWg0sFnBJQ3J64cGCxGvRN3WOxYXi7iCPY
QL9BjbsbymNKo4E/y/1HnJyen5zBid56hjW2RBBY7X8UOiTMSSXkF42e2vDlJHEixGzW0UBcN+WU
sM4cS195VoOB1fcCsS4Qx3cyNgj54X5DpEUCSkC40l4ZCcMYHtH7hWFozxUl1HLySkoU8u8UfH2V
acpucnIQksAIP1mB1rfRKsWRYDmQdKPKeQfSe1OehrDvRqz49Sw03v8Zcf3tPYm4CMXmGW3X2qyT
+2jJfogKe+o9VQEwDDJJdM1jdmyim2yVij+/upak1OVeFs1sn97P+5pigbv6O2gaMuL6tbgX6IB/
DXNV2qzdIPIkCQt9Md+uXMpFqyrj5j/eU+fhLM8mJbNLX4FZDbXapOHZylrkFwFv00uSRjayyrHr
UgLYabwTDxPab0+WFhZt5H6Yqz18gwkFNnFBHpAGq+76XJ5uYGODCmuHqNayWUEtWzI4jUciYIyK
03NMWJMrYbTfAfAbopVYmSrgFm1fI1rWIZLeYAHJ/7oDxIGcOViSIzrfyBmhwoJ56VBwd3VlRHDZ
2BvMssTMsA2qXiwWKMnp6cRiAojsy20iFKMC44RuZonpRt7N6ZFLjl81CvFQN3xUOVTqbtcnCGF7
h3ifatyGQAlQ/B90uslStAlXGYK+sWi6Gvhw3l3/rRSuNryArnk4dMbh1Vv4PrZqLXu+FFOHFUIy
9DL7hIYm/3SKabTsu8IE8J3tKp0wcmcSNUOLDUzJ55kYPC0ec/C6O5t37exFSC61cdX5I+y2/Q24
wRCEj1syj+5whwX/hKgE7pyv0bjGJWFUtGH/3E387acvx6yXiy1eTBNFhS4LpXYSRwQN8L2nAJVg
dYuOJ+HcHCCn4V64di+JG0ePquoTJG0u7v1s3yNGs5NhX0U6tMSQU8IauemyKw45rNDEeaJOw9qS
HX8+vQ+OKmj8mikf0IATcJiPpq3rmqLBGPXfO6day9LakmDDxshKyCoa6L8a67zboeqVBfttL1NU
CjMfB6QKfZDY+kYXAKyoUFsf8Cc5uzqS6kL50he4O+b8GmzO0rkHpFjNofzEoceqwKM0MtlBweit
NOeURbQdRai2j/gAluIO0q2c/+bqJQywEd8L5SOwNHXtZ9O8r1UTcPN19u+sbNVMmk4dKdMToWvH
Pq6kck7O3dElDidNJiHUxlBoTH/s6b5TCsa0B0McEu2KFu+SGTtfdmNmMJMid7EDBE0LVkxLiNh3
jR5GBWfhNZkGYexFUFkLmJiBwgzXKWVTG/eNuiXIsc8QngPgaSkSp7r0aNXGboy6pHAhUpAY+Sv9
nsX1o62Wg2jYHVo0NVz67zI395hmvJqMaXL29GHw59ZZECR/XZbfc6UGeZvKrpwxApl1PqKT+/ap
GsiwTPw683az+06iUJcBPpTi39iOEBQ8Hu1iuvGIBhGJLq4omkWPnzH2Gv3pd7BlxEoLTv4wtVD0
Pe/cvDv9WwYxx5pZ4mJ/kXDtVbempDkbRg3wiHN61K0j/Ul3bGtVmT1nx4irEyPcQEsfsICPQd7Y
ehMX/TIqJBa71m/4WAuMNDhWRcTk5vYOOS20gsKnDkVqiu4RguYxXdgEz+5bGdTGABW2At5bSxiS
ATQOFsIxo77d4o7iCT4TmkHKGFMxVva1Yecd36EWpmxWZb2syIYblXU4wXCld9SyvsD1lUdJlTWt
04BkipsrhrHqOR0Fbj5oq2j98AqkwiMHv4eztiY57z1sfGkVTprQCpmZUMgMc9M847RnY0DyUEps
tGmh5aY2IjUGk/O/WZnwke7fUipTLwPZq7vIb8xwhfi90b/eVsEPjMywU29NRU4JFH1XdDrrLoJP
T5QxkFdWZCu7oAzD7TMorXipgD68eBFrPC4VmSiOeJOswCNX7ty0OaHCG+pIcW/8t0bFdL8aVaG6
Mln8oWkBVtNpmB+2BL42H41Jw2S7iBTquR4hfpC0fUCiq+5bQ7g6SiH5ry+Rjsm6WCedfZWQN9vI
vUstK3rodMkZZL52+gQjMYZeB34fqDbSHTRjuxBgq6k7wQBC2GHF+liI7LNMWPGcFz5yomdtqNVq
PVeA+m0Fd85JC5IsWQohSWsJRie+QO4DLEswcD2BEQpdmNC2mbCeApYWTE1MlsXQOKacEVDiTngX
clUN9bCSlPC6OFM04dvkm5M0ZbXiXNsm85YXmEwvvlMfzaFGDIUGf7FtpKj26y4tBezEi/wXr4At
CiRvnOQTXbA6t8B2IGLLZS7eRhrFIGz7U1HkW5vrYSJ27HwOXlfHkmCyG9CCJmZ9/hX27/BQ4sr8
yyWFWlQG9ndpQkO4tb5PG2cAD9+en3NbZCOdLkF36CDUfOUxnCn335QXE8TslLVHmoM31DGY8z9a
yCNFckbYGaMSdR9TH7fqRiNXKUmoVtmOWWb8oztIolzyXxROS2+PzzFZz4ZKLJhJpN3dASxTo5FO
kgLYu3NzlmjB/YVfW3bZ9/wMt8LWwbcBhWbMTOxyGnWxh21q8XBHTxRCoRPebiCLyz227uZEUqOO
6+4irLIS9W5/sVyf4loDT/w8liotj6ZBjck87g6QJ7eLis6u/b+wJupzEXk2vLzIyFT2CyrkE55M
BaImWIBTA6j4WquLmjVXrt0kv/tqVq9ICf+QtTqYJas7LCuYhjKjSamKJcgP/zdq+L14nmYY5hPP
9v3Zs9kUFUMwcKOAHDfJgXn0/59IFtgfWhMUhwFgDHMTtkvbEv1A+fYVm/kimumZm0mkXX62fpnZ
YMpT2gmeQVDAn8Sozen6fFs2D3jH6I8pZApZXtrHoKsv3OtejTedpmwh8kHP6JoF8Bt+y/p0fD0j
j+KTjZLxaZLW4nHPqKOHUMIKPPE5R0WtWlGFH8Anm2AaWhJn4sYuKYRx99hCNGVyS1d4xeGp17mc
EDuS8E/NaUQJ4IiA32v+x7q9Fej+xIsLkeKFzsr7CpguItT0o3s38pjMHF7JatC4wgqFb9pjZN49
xxF9Ygjn/yhTGBiG7wCeiSOKfaZDBnhzVCCizAzgDR55x/izMqFTieJNt3exDbHFH6OYVFMzIson
kv0lTlqO7USutUG1Vy1vhyVY6tzh9B4sqVwV42uulTW/ghyVbZe+XeK1Al1dR9K2Nu4fz8SeElC3
6BNudMxTbOEKajVvmruiI1EYF2tODyk7mB3+tkVXxg4Qt1KIabetsgqt60m+jFdG1H3MLi1SwzBU
U+qP7aLR0BCLQMrd5Au9SgAuibV4yfCPCWkyhQK9eSfB8Jrm7mOJnoC4L60x36Yu00b7SiZkYGoX
3QfHw+Y2PVMU4Yr5+MqgLdkXi3MAu7IrP6g+JI9EMmpBzg/uxOKCbO2ZEdNJ4oiACbUGySXoiFwr
4JViBOrkmZGYYsgj2enws8kdABC4h4Qe+7EiplIn1jFcZALK28AAtjS8fS7KhUe//65e6BjXr+CV
V2ErHzxadddyQ4fi1ZzZ95oNZszNCnwa+JBFv+T/3Yuhw0iyBVQnytZJtg1bb3wG3zYOlTDIC2lG
9j1sA6Gq0fNYhhP0OHxoz7ADlZf7BZhWT7nN/xY+2tYOXX2YtIbvSwP1ai9t9MH+kbyGpzWFE9Hw
LqAvrIgiIKcj8p+287Ef1oCvXjKEJXofZ0lwMpKun0/C3L2aqsKYTd1GPLqSc4NrZ7pshcrqq9I/
+RDcUvuniEt2Wq32/Rs9mLkG8oA447MdvL5iqwnti6w7IBmnYZhAmi4Q/LJ3NpD+u5JpvEE79l2c
2uSkUsjCjRXaXg5MWRDDPMZHEwg/4UQ2ImFIYizC5IW++mOH5Jv9D+nc5m47keQqlinZiF29Rea3
W8gtJr21brsI7UA0MLoMeigwtpohGMpBc4BRLOz6l5AyQMOsiFbMWXy5BJz70Q8e3qk5sEGrXGmG
loJcuARRs/syUwMVmL9zd5qoVsB+d4ZRNfsXqTtqQz5xDW9mwmYziGmL5sh5ItFJvjayHZ7KnFQL
9RtOLCJk+/XeM4wjwO5upemaie1LDTyrQx95v40KkbS4/fCeQnDqWj5LuEW8t+UYnLIS9qrkqUED
jE0chLhpSDrvK1NWZGgM5957C5z9MwpT9DWN3RPO7nwy7ncoFfAtD0MPcvPJsGtDfioyGd19wn6e
X8e2aVB+HMk6Ni0ghDB9FfRepOBtq/zOYGmhyugRvOvtgbG6gJqSgg+Q7FFmbqKmdl2Q+/IBQOcu
gwfQtwT1zwCXe5lK2binVL6CG6/GfFfP86G8rxLHrVL4jUEVrNruT0o1brRKMVCkitOMf4sN1zEi
WPmhRRcDV6S8hCXOplJhnwoamvmCgBRVHPAahbomh3myOuX6ZLZ1U9FuF7WqdxPCtvLemQ3C4xxa
DZelf98BxHZGWpAnx1gumDcA2bfYHKcLe/mjmmA345Qh9K7qCUYKsKTKryYh/P/Fms1n1j1J+VlC
5Ebu6p1SAVTVPDIytHHvjaNUESbDE63iW8kuaVTjLw3NiFa6IqNZIDaqZ4nkPDWtTacgqXDpK1TI
b3NMqgYaR7u8iZhd74pB4zllxu8quamt0JfUhHLohbeVUs1XZN8PjZHVM9SgSctG5yN70oJ3/SaF
ZNrxVWYvHI88OLvi1OsXMUSPxFV1pqjQ7qBzn6f05SEg0plDvx5YHFgWEg1OqD9nOHKameKkJDHd
b6iKxsh6DehfcQQ9MMK++/j1tm1ADb6LgVAQbXNnVlsMlBQ2nF8vOfFvLG1Eq+X7WHwoV/Sbow1H
0dPalb/8xcgeo6RP9NW3vjWVrHJmbjlVFh82/Bbow8lRhbRzh/WHAOzMT47fAGQqh3DzxHm5r7gz
Wt6Ee8PUnzZ7TUDY8elMI4l5XGf252kCvo2xfH2Elg0GcVhm3w/vVyHitzDcC/CaS+eckdDptVHy
pIAcP7wLp8VyL9v+iG/nIZDH0BZTQBSHUyDtbIzSWnJvUd7N2527VB/4LEjMswf/fwQVJRD/+MIo
mn9ZxAuCddP4odYDYXWSSfp2U2YchLaQ443MDr+kfh6teyUYCJDb52MoZa6gi7qNqNH0xTOXUyA8
g0p1NZdcNplP6DxnUspcHfIuYJN2iimwV+sfhc5m31heiKXKI6qGT/RywU56PI7IX6rxcK0pREtD
v2zlK8zAi104R8FNDPnJafNzXvvniHWK6/F4btSo0isXMwySxEALjT6AQ9lzLdSQyjpiap3ZZ/jo
fValiO5iIhpN2+lsduEt5hEooaEbdnALQqcOhD5Ln5XjlTYRO69MVj/XXdLipGFfF/vWA4nisIc4
ZXcABp4LQC6ONa9jb6QmrkQWey2X/ACaLdR2VXxklhES8fDkPWWdI8EMZvvyG+JIilDAMTAxQWRQ
YAsR8UbZJI2WOGpxAD9yVl7eugY7nHlTnrBUohl3mABMhPZSpOiXudE46y19RWObn/xQJB1Mo9P5
4P7krPJeKJLkf56n9rTbs/Rlikvnv3bO4W2qKORvi04/lYV9y5Xn7pDkvJC9s6YpOozwB0z/yIcW
2z4InDGvIO+tuAC6N5F1BhUKlNCzmFNW+s69or/vX8pjnTvXzMXXJNgAKKKk5tNRMtZ+ORP7DLQc
7JagV2NJkc6c4J0wBdo3TE7kqDQYTlHnb3a8h3zFFumLvQNqcxB0RJOq6n3htbYLp/6gQgJzAYif
fKJk6Kw7t5fZttv7VxWO2FOGAAXFt1k9PS+ewukN0gBj81WEJAspe/vQISekzCXQ/ABD2bRjrPT2
ozILqh+7kfHFNTtcfiCwwix7Y0+U6ZKUp8bU8YKR2rzixV5At0OR6NjT9epsti4SEE7aH9ornVUR
3ERcD9zaOEEhnKX4P5OfzYtV6IsrL1kmvNx+Zbr7RG873XLMD0j/uUVa1XDktQ+7+0S2L8qjtm+Y
XCOiFBPVUd/cC/dcQbtLf3CySKB7lk6H7zQnVsnSt0IhmHohrD/L8to8b6gz8UpDek9uhZ7QRNr1
0AqMIZ8ffad9dy2gTbrWpzWZZF9hUXPkSDzdINnC97Wy/4QZ25PAnoJvBfJ5rubcXSXXHPdqvSij
oziYDjDkMmtgaxzi1Cbo7ctA/yzl728JHBwGEjJn3KP2ERvZaJNXYGrs3Og8BM8qXu7lPhlHLiM5
QdCAb7zvNL1Bjh6/SJcuznQ28t5lhHCBdFJ/TcmdAqlUBID5mxk3nRkhas0hLl27l87ehqADRwL6
5MKNQTEFVIGkENbAyfa9J2noMh46GwgA1ExtAhF7LPOXf21aQK7Edr+C8S1nAl8xE93xT6d4JJnh
sOI3M31hUVyDUZoqp16oPi+LcsQSAR3r62z+GJPIJ8uSxWN0MZMhLoHrdIrhgMtPO7PmwFwOlZ+A
N20cCtgPKjJlvkGz1IAwd5oAKzViREnyfUTDb9co4n8y8P1x7Z+B49XcMf8ystumgl5SnGdtxQAq
gKK+7Wj+MvS3O43QserNT+enDQlvzUF56VCLtlyQp1xByx3gpJntBJrOsEsNqtGf7U/TcP/mZer2
SluP2C1iJA0eky2j3zkrbHHxPv2dFgPPJ+4FkpfN3M+f8ur0Tco6gMWvmGkakMvs8a/nfiosF1al
BRsCv62lq8MTLKqNQkE3d/5wS7Oc4RO7bu4+3uyO6YVivIHWqDNDUu392yzq90k7YwDcrgF+Ny8v
8cyzLNqjigXv0OUmcvch8SIzN3SvFzxMa3ZcWpg5En9HGms+UUtdEi4lhjeSXtKQTZGcmtNPV3ko
tTcPXzBDXEpoLJIrwyN8IsuytS3oK1LvrpdrN5DpnvzbjO2sRvDexkByxd6ec8YkZy+7iWoHhnFD
p/GpL3Z1Kmk/X2/vRRwhIQmx1tqtyBkqeFlZOfC+dqVYjWEGGWD0b6CtPB3ynVGdQ1M298anC4Uh
Y3lpTYAVqXbrm9BFrllMK5pmLihGmLcyhwh4aXgT7UEqAWjJf1r8BWZl6IoJoB9c2qZ/I+74O8t4
oGiteCDJ/upbYV9yjMd0PVptVCxE2NUGAvKPtBkHOoVA0b7O6VqS5rjcEQkPoQ8u9QEYqd3XTxcU
cjMZe/y9KGSbFB1kpbUFkH0FP+IY7tA1GVDYVn1KQzosw48sTgHxsBkbeSxbJzSufah98aSx8vx+
PnWdnYCQbqlhpoWgID3SmPcPDh5eC573z2HdA8MSxUH9To3/7blRIWGm4EowNNwADVrFMOC2zRqo
xofJqxd97nMM0/jEl0UyaSaCnpT1cILxw+5od1clx+G1vmhvBP3H70mt2OC9TP9YV4CNYFEKB9Bd
3QD9VJNvLAHPwFwmQw+vBao0O+H9kuezGcekmlBcOIr+jNhE7Xg/iEd3IK58VpO+F8xgrpBov9sh
4iIGzkvHHm39gwvneklkkjzotO0LSXjcd6eKDUa1jkgw+HD4pqQxfMIEqBDdb6/WUqMCaicYXSP5
sNx3W3pIL+qYtfjXLlcQz+RIo4Y9OURAR06nZ5Nu5tsQzJYxA4keIaXzuDy7Q34zrdBryDs/dsPb
hMNEXfoI0z5rUOqM1wrcnUKqo/79e/0IKi6WUI/zh0/tbOdOuv9j/x/ntj139rSnwdzfcTey9oGl
uiYXixkSggqatJ+11ErsrV0xmeY9k/koiV4ErjFOrblhXBpmRPUPVzSMaHhxAaNWqqZ2V8q3Y8qc
+WlsVutpEo0D3qAVFNH6cAnak+uNODqijMaksIBXr6E8HDioEOP0uPPRU15iTyS2cNq+5GaorxdK
Oi9ZAA/VJClDrfNbgGWnXZzfUakdJaKf14I4sKK/EAdsGWKocJi4n6pNSjaF9lfkkGNHxQ1w5ybo
A8zuDwh1UTLF8MDxUloV7qGMEo56Ju93TrY+yjY/ip3+GSxXZ2xOHQX9M6w8kJQ7E+mgU4+dl9VF
qeGn5J9D4Ea7GQ87yUWSkh3bVbP9ylKUA8gYYLUh80lHDq8xyIO5GKZzwQs7JNV6HQk1/vrTmasN
HLAQjAJEaMp3nYpRhBD/dliJvXhCyB45W7ofDtvXTxs+fbMboYuyf44tjEjCNF5/uurUgp07eja2
bkCVnxkagjFvsA4T9svNZ8zp0ae1TZRvOwvWZsYAA9Nw59owN2+ueTNB7t5FdZ6hBc4mzFZmQeud
pwG0w3Y5bNawU6PJUAQwrh3qs3hSpFb2mwK7xF8fcdNq2HbtO5YdFeB9ROEwxudPlASZWkHqgGCJ
KyvhE/sXDi7CljwYe0Oj3+9y5GKEmHrPgFewWKFos3gvV3KqIaCZMlb4jUbPsljb6uIH3dr8C3ac
UbNuOjWGt4Fxfbf5fxa9phMFScopOAD4Ok7xb6ePHnOXpCxkdNR138Mryd8q0wdCGCGKXRtttY+h
jpkgsa0zoRD6wjHKEemVO+oGwvrCwsTicnB9g15lkWsk/GyvJkp35tVYjISWqoEaXiLAaeHhwYhF
jaRkPfmUTH18ZSF9sfSsuYZcqE2e0SInyz6PG/fRfs0FnuQQG9lJTH1ncVJ8QN08qBGRwyUQznxi
ltcPaeGLoBaBP95Hh4eJ9egcqTy15/5D8tRzptZJ1tslrGCEmy7BXl9IL/U9qoW0BwfoVWh8V91V
OZk8kfttGv1swK6c1l/BV7aOr7rxj/5TMtWkx6d/zbISWl3aF9dSPPcCIRR6ctc3c/GlkE1GI6Xx
gW5xkGCsa/tLNs06xe5NYtDh5wFyXquMy++vpnWUSlqxx4XxTnWHmEmQaLlFBTGNHShXvsbNj4kg
9ynfsr/bI52wAt55a0Q/quVwb0ympvDAz9JVJaCZHSIJo79q5qA3WxFiUjeYgr8Yt5HFLIJAaCOC
9qfxWLINep6CEWtZevTvCk+NziwgpCl/QU4gj65McXdQZ3IbF/wI9Ay8QC7JWLR22MkgXI2mbgKF
2BwhnmD8wXudD+IRb09ey2gw56j7jvhRW6upViGe6UY77zeMtlOaMSrVJB78DAbW/slg+tDdCwBr
0p1pAciAxCEEtR2KTX7sDVMHXgkKLjZEogc2qZ8DsADbWVOrRgXo2aXPIaWDcGhjsghBU6IAFtwf
V8mFqJ9AiARdyn7tJimOxyZ1JJydeK2/ji4tnmG2s1n/9MFX8NY8xwvyzA1WEXlwuy/N79rnDIzq
4jsN09vv+bDXrB+SGZH+cuD0NJYwaYG396Wts3TFL9ln357/WnYfXyGC1eWjzArYA46vjPyW/RHo
4G6AmupszZZx1Kj49JEuI8UWnOdDLAerRIbYOpc8LgKAmgrTZi9gKnssx6F1JJCTRFKtVwCPwQ/C
vmSUkvx+dzRHSdsQ0aOG1FWyvJyv0nIcPCcndWaC3wOzuX8Hd0tkn8Y/b/zYOE1kqX/t4h0Sms1p
aJKDQU5sM4efAXrTfv4GpazyUATfaWSrDIJmgzqO3qkORG2VnFa0g9ENw+utgTnZJT02wJZ1P6RF
Fd/jIFdCpXJdbF4LMhMcmQHDyEmG78LERcHTZuKtZeXxcyojN72Nrgisu+bDOgyAczVL9lz0MDKx
JYmtWRbLamUbt5ZhMjgBp1REt2bpROYE79VIsekTKP9Tu5Su4HhpvAQPY7IH+wecjWge51UTpgWn
6xV5jlZ6e+pou3oHExYsiZkJHCkgU5aV6HbXM3fcLNAbpzVZadUwdtkHlHbjySLRsE1myCePL+Zy
4jQHYpE+JnA86IB/VwkPA6GkJsYlO2Csms1m4Pz9A2HVo5o6KgSAFZTbAvz+w3rDbyK04fVkM9MV
O9FtCwQlBodVNXwrn/YW5434ZczA7Z3onNI8IX14Pg887218Rcelc8tYKT3NfIRWKx1OHkaYLzPM
r5EB/GxVDt/4aU6UEDQdshNCvVeqRm8PRnLsNTtB30edmAEAVmYQ9BmTA4JkHr0bNhR7ybfYs00r
o/y68bks1cWdSeoLgNNzggt8K2EBd9qU/uB0chymyHtwX2K5iAi7xk22m4ZtmzENtXnV0yivYa8H
PSKrr1zNw+Sf545Ay8BJcWEp8aIzkA2YfAZtbjEZItIGsaHab2G0Y9RZoZJzpXjetPOa/5C6MzeH
7gHWlzwZNZvaQ5mkKUqB/L0IuXaaJNxnC1m3ggL60GsakRU97k/ECKkBByJLm1hj6gtmEk2jTbgj
TGWpCL60BEhiCf00B+RMikGJjggeQnB+1NdbGWVRJiXBeyBdkZ9O3HD7pI42AO4NCx5cJlAUhH+Y
0sowfwRBXqVW5nCqI5s1VLSL2Act6VEJ+apmXlTm/vc07P6RsRkDcgOE+FKJ4Z85gqF4Rj7KoSsZ
bHUa8LjZSbnR22kVBKwiE9ndzQy7+XGt5X2NZDVoj8E6tXvilJwZhc//KaY6nKrZg/9nASbf4jbI
zaR3mzom0TawxpJa01oqPCvDwoiCWErhiQV3deE9BobxHGPjHi2gzWmak86VJ14Y4XK66fzVll2m
MbNvnu4XqS+4T+X0mEdI7zsIgIEDm7xa9s5WeusqBZqiZIPDcQxo8Hk1WOuRpAnVmdStMYll7x1H
niCAiglmaddxTpPoKgEJjk3LRMEXl5C/AeZC/Mf2bhH2HZOiqb9wq5eSpM16JtsHht195Yi9eA1i
feYllQh/jdS8LaN9FAZ/RJctEyrx4DgjhQjAv1b8mDyhKe8X2BL1muDsboQUUIyD9cgVAaZ/3013
Rv8AQkCrNhyBxOU+VYpVNZwqH2agIHIybYknNt5ON/iP11E0u6UoWCoGj8xa7vNTobKzkDvHeecR
beXAaCFhhJsJ1prN08qFkCw8uwZFZckJlGxbg3r7hRvPh2HwyYke9tfz/IajHmfybNM9mZ+qXrlR
3qp01ZfMU+foHrFxK+3VcgbixoWyytraiaO/XdTUh7GpSP7PSk4qbTr3DXWNY5z0xY0/ExRLnYUl
j8O5MiG6dGH1b66WRMJ8ijGUxLDxADJFq+4C5MBLds3VN9U48DOS8ERv7QUqoSm9zaQHKbojjsO6
y0H/ZKZyGrUHSqXgXuBfdXhLHhDHwObS4Qb4ur1A+91yLL5ocTH54v9Lmv6lASGAyflrx5+S4oxB
YCeBYGSMBBUGt9mCOBO7edhGVsvHp4WXvZqeIkjWCz5xfVit0Xhtm33zVYM9J54DwHBlcl/LtkR9
sNhJN2ohXC9PYFxZhNoM96rU1Dpp9+kwHK0E1Jh8YmJbEg1p5gL/FBGQg4kozxX3Pub0snKzMK4K
tKIRES8oVxnjvUTlLFKrJoFpQdZDhUpHw0yNif+oY6TMZAbbEkj+pQepHMQpJwzPKBUnQqkb/8RE
eTXu0dLsZMIVvKRRgUhIKT4pe67Qa6FjbdJiiSSsYrdVSReJ2tjL37s/7mwY7x0Kgp9xa6so4CsM
WoZRHvNd/wtSXncyKMLjfoAILWWbviWcjydQdvF5VfGrasYnuW0d4Nf2Eoc8b5GSWQrnxvO61A3b
Ug+x5FO69rIfXCI4wCXJSxMKo+EvLIKdhF3nWh/tkvGRmNtMH1EfMDy++Q3KtP8dZafZxTmHctvj
xQpg6QS19pJZ0dHwCP0IzmovJNhafdyCwdTrUlSJxZt0KKjB6YtasTlH3XfzKA9MHoDVIw9LjVWq
QL98+RZB7duklHhHrPBfNyOqVlXAc0xUtkp9ZuNX6NACsUPFbtYrPQvZVhbapdVaWquvxin+jcdJ
d4Jp/r2yVktdw/vuHUeOYDy+pH5TElFUZscmNFI4qIxSEqo6vyoUi52j5ZMgdJwAp1zmcgPevSPW
NYbhm4pbqu/L+2tvOav3a4WwKUmz6uL6fE/Fgcjop78Y9tza7LnejrGiJSX14vJa06+c1WQ3EGZI
l+a4UYQkdtnYUDcXru+RSFZBe5PxrD8AFX/5tQuI8KIeLxIyx1dYNZWMnTzjdHSdqm03SKupw6LG
TrisflJhm02unA1viRlbz157jlFwkUTBfKW3CGaDR+KpDx3M6JbZ8mcUPXimOq/U7dS4MqewP8Ha
P4EwdZHjTZWKiCyWwGNcpfayn4Sh/m5yu4tEqe3cFBC3uOg0jSFOPIJFZrNJBes4K+gfbvM9/j9r
43YWShkAqYKOYfKPCIiGap9+Y6dXucLrEsWdhNqGRv0Z0yZltA9UFDceFnDeXawpK2C8Rhpz5RTt
Vp4tqucM7tikmdzZQEv4IzwteEoMZ6bvVOQgpXZkRtiFhCnZxg6ke1YfFqgxNtFSgy9lcPnRMP0v
McyOwM5JIhs6yEpgvZhDX6hyL4Q1CPXxogARnvcqncGwfKc4VucY+b7UbhZ4a8kpu0bqZ2iRderT
NUFumLuSmfvvmvl7d/59ZAx1fmiqqMXzFkBKRAKnuh5YXjPd6AE9ZizRqxQZJvTjOTDTOvVF1YGo
6i59Ye7muFdFGMvEcJSTYkRKhSTJ9t52LqQ9mKVUWuovruxh/YXI9vwsSAnXB3jO0ILYHoRvM3ch
zYhVd4Pjsz9L02+nD3SJpCSbslhYUWGO1XbTw9rFWqL3c61k97S9jzsOIdctuFzKZjuI3+/nhADQ
q6Kd90tfYCHh8l/qZUKEldX2lewpeu4wxseKGIVPGVEgGhDd9fK4brqxNU/fsLeKGKGLdoE8kke2
6z9Qkv3TMGrQmQ8WeObsSghmNnQVuncJ+r1aGGZ3oagrTfhBy6LxnX2R2x8Pon6zZ6XfSe+Xfd4d
CLe/RboM/gr2stpljQJtSkSqOL1yEZ4e4CBugClOy7SIYnDKhXYS6Bh308DK/Rz5F48gHp0K/eEX
IyNi9W2vphtkgxN9vWtZI6HbE7zKUIgQq/q4cskVUzM3cNtfzplpOvuOknPwMc8fV8wKIdSO0HDG
CbZTnYc6XPHXGa3McB2oAskRnYWPeuAW5LpUZfp1GbxbWbUmHmTqeZy/WF8CXW5Rfc1cluiCxyvU
OGRIhh7M7XkmH+/S4QNXBZ7fjgWfjs1SfBsBXnE79CqbC/V1qYtio9PuTo+mtacrs7p/YEiro1uC
9bjZLpNnlUitg3XKeRbgsG5FSAgsv6byZAHzAvcMQfQBoxjpehok6ZJMqmNtyB/fe9yAtKxZY06I
eNCnmxqjypZHuX0pFFAJl1JNgiloyyviqcvB1pUwEFArcAzQ02yVAZypUS6rzip2yoCHaKzGhyy8
mY0AOJm5IYFWWClwwD5XSImTYjZEw10n24Sx/GLnjOoBxjuyZw28nouKvJnfWGMjuAN/CyTOtDhO
fRGxD2fnPg0p3CVPyLl14G3SkwZ1+2wvgVnEbDRIfQ4+6FDHUC+ZfRnOazLV5BE8RJrWqLRjJmWU
uQDYDfWRbLkmL5huBdaCCF9cpqAPdpb9KE0R9/Zy7Gp0p21GUcFMa4GSA2thzxKxdZ9UZUfdHLnE
B/NQAEYaqLnZ6RZk/s8QbpPjeP0pB4LRW+RqlHxWfJOxuVYlRwsoBk4FF9Rl/b55ZIO3KE1WGDkP
LujVV6oeRXQRJuiG8iX1pVswBOadmhFhZFROQlbmZTWLH8y+7wdtr4TZPp1EAZua+t6pxYrLz7Kh
SOgqUqkY1IIj3ca1TbTU5tYwG31dXXp2cIZ0QBbOTeEs3dFz1Z0YxvAWJ/WiuevJFD5zu5vZvWEV
3zYHV+gtB42g8Hsr508lzHU0EusFhUFIfmVdc9NqnZeRgOmVWKUuQcXv+0QP6+U/E99Wo5aEJu9s
MqRS3BJDzPRP4IPF4OIj6bb2CDjb8a2/QKexOnzOWHL6VbvkK6HrlusEpTkl4EocJzK+soe16xwX
FagmSmUz2MlaV/fQ9Yqy04vugxAr8n9RYq0VQ2TIDsQNFwaxhWV7u06D4k2wauR8KMJ4+m6AN3li
miKnh5TahHZD3r64eQ8mThI+g71he90+K/PC3J8jSiNRAZwNw/mEGk85N5CD47dg4X67up/3qExN
HicfJ2EaYbgGrkw0HoySsnvDzjTGhcNfCOumLEn8aky+abYVuQ61oL860RnhRnIcOkL0nNWHPiAe
HzE2llb4ZHCiPAMMhtzQcaJF6wfUK09ftvCrvewFUxKQPTvVceIZUq1pF6Ko2pUJJVi/G0EUAcga
FBj3Iu/DxfEG8+o2EugDw+vQUx9UJXNGq310Y5KvXyCRg5EtxDjSas5lu4gTNdCnPMwi4IanAPjw
x64jC6vtMIoRfv43fP3r24Xw2rNtIRdg9fG0Bb+9wQZRV0Hd57mZqjkTe+3TJHT7yCBKVTuK034S
XtKsrYh4GcqFpWFWNaRM2+ATBZnarKt96z7hDagqTDK2QjMF7P/FUqJtO7sgzyQUBfGNsAYaVXcY
w4IQUonNTR8g3/VlmI/rzHxc1n904ZDT3NtK6Zkdun09jnezvwU5LEobUbgkrhY5x8hXLJu0zvct
Gd/AxiEdHGiqK5ycyn2qxQtOvJXFx6mULf4eTqvsb0Wuzkg5lLV4yEPafwoFp5GIBVGm8BuranxX
9OtFkM+v+NGy098upWXn2JqowRjGAuhdy77DTW9H0WvpnH8+iCQ64OSugVY35dGOpFIPfEQgjU1k
Cr8M5cxMy7dzmJ4inpHcLZPDuB/dBBj5xn8Pe2OnJCmjlJy5HK8sIexYZBqP7IUVz1THlrGji73d
5IUpy/u2hFwtckueAeVqWLClcTQ0TjyAkL2C2jaVfQmxHvbtUE00IRuBu0J9P9SeZ8p0oOs8ZMeh
IqZsXOXklo9DqTrxUmbyAlhi6oN/Dc7i/TLPud+XKLPa/LlAJLyXHNk4vVyRw08zzq9MId/jDHrF
mViYDB8hGWgitHmX+cRLvdDR0c3eG68I7IrrMzelecwcPqrO6lT5M1t0rBuRBIYg4xKQmSxshxCd
qE/RmxA/dPI+O6J/jbLHiFW0Vsrzm21wWLpB7UgqugoWHkPv6HL0oe6PEHzVAr9lxBx69Lrg9stt
5n5Hm8LqXZH32U4S8HmKXXtLsO1jrgRzRXJ5kQPUrt1agmTE6h2dkYcjch/Hxz6+OWdZVx7z70dE
VsLWp0RPsdrdqNVM8o5dEhM9i7G48XTRodLTmttSTyCDg/fwEedqPnex/5uUY9vLiD5O56k9yMEz
UlifOLiAXVZb8ApkVW9Glu+Fzxzlt5whgN4+GhKNK5M9AXOXb0DCwzrHHE4tVEAo1N+CUsa48gxF
xIPaigXQNM+qXrrPgAdqHMSLMYv5OJIGpULkF9tCxcNJdu1n1OKrEEYebbYJ1iMQXjdVmfBRZYMc
RBdGcmxaDTIbof1UnstzOfqIDbYmn0oRAtU17r5aDN+1WgHiM1EDQEgybmzcXHyNWd4x8if4sCqa
Zz9osiZHexhzJT+OmkNg50dpEr7dGFSNoy/8tYSVl93IKCN/I3yGgYWcsVHhsDkDa4Sofus/eSUi
RBPdt0McYztO4Hq9KbssRJC0DaCaVzoAnXEL3111/+Ab4JzVyaq5v+GEDdm6KnLcDWkN0eowEOFU
atwlKxz3vw4UU1nH1PPSQZXF+uKuNmeMfwW4kal76bf/n5iMYJMQf6sH+iuw3g0nI12vCQOc+APb
EPqGr+sMBAbt3tFeK8vITpy4XZG3DRrm/SMc06V8TQ==
`protect end_protected
