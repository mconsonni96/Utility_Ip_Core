-------------------------------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------------------------------------
--                                                                                                                     --
--  __/\\\\\\\\\\\\\\\__/\\\\\\\\\\\\\\\__/\\\\\\\\\\\\_____/\\\\\\\\\\\__/\\\\\\\\\\\\\\\__/\\\_____________          --
--   _\///////\\\/////__\/\\\///////////__\/\\\////////\\\__\/////\\\///__\/\\\///////////__\/\\\_____________         --
--    _______\/\\\_______\/\\\_____________\/\\\______\//\\\_____\/\\\_____\/\\\_____________\/\\\_____________        --
--     _______\/\\\_______\/\\\\\\\\\\\_____\/\\\_______\/\\\_____\/\\\_____\/\\\\\\\\\\\_____\/\\\_____________       --
--      _______\/\\\_______\/\\\///////______\/\\\_______\/\\\_____\/\\\_____\/\\\///////______\/\\\_____________      --
--       _______\/\\\_______\/\\\_____________\/\\\_______\/\\\_____\/\\\_____\/\\\_____________\/\\\_____________     --
--        _______\/\\\_______\/\\\_____________\/\\\_______/\\\______\/\\\_____\/\\\_____________\/\\\_____________	   --
--         _______\/\\\_______\/\\\\\\\\\\\\\\\_\/\\\\\\\\\\\\/____/\\\\\\\\\\\_\/\\\\\\\\\\\\\\\_\/\\\\\\\\\\\\\\\_   --
--          _______\///________\///////////////__\////////////_____\///////////__\///////////////__\///////////////__  --
--                                                                                                                     --
-------------------------------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------------------------------------



--------------------------BRIEF MODULE DESCRIPTION -----------------------------
--! \file
--! \brief This is the testbench of the *CoarseExtensionCore*. In the following figure we see the result of the simulation.
--! \image html wave.png  [Waveform image]
--------------------------------------------------------------------------------



----------------------------- LIBRARY DECLARATION ------------------------------

------------ IEEE LIBRARY -----------
--! Standard IEEE library
library IEEE;
	--! Standard Logic Vector library
	use IEEE.STD_LOGIC_1164.all;
	--! Numeric library
	use IEEE.NUMERIC_STD.ALL;
--	--! Math operation over real number (not for implementation)
--	--use IEEE.MATH_REAL.all;
------------------------------------

-- ------------ STD LIBRARY -----------
-- --! Standard
-- library STD;
-- 	--! Textual Input/Output (only in simulation)
-- 	use STD.textio.all;
-- ------------------------------------


-- ---------- XILINX LIBRARY ----------
-- --! Xilinx Unisim library
-- library UNISIM;
-- 	--! Xilinx Unisim VComponent library
-- 	use UNISIM.VComponents.all;
--
-- --! \brief Xilinx Parametric Macro library
-- --! \details To be correctly used in Vivado write auto_detect_xpm into tcl console.
-- library xpm;
-- 	--! Xilinx Parametric Macro VComponent library
-- 	use xpm.vcomponents.all;
-- ------------------------------------


------------ LOCAL LIBRARY ---------
-- --! Internal Library
-- library work;
--	--! CoarseExtensionCore Local Package
--	use work.LocalPackage_CEC.all;
------------ LOCAL LIBRARY ---------
--! Project defined libary
library work;
--! TreeComparator local package
	use work.LocalPackage_TC.all;
------------------------------------
------------------------------------

--------------------------------------------------------------------------------






ENTITY tb_CEC IS
END tb_CEC;

ARCHITECTURE Behavioral OF tb_CEC IS

	--------------------------- CONSTANT NON IN PACKAGE ------------------------

	---------------- Timing -------------------
	constant	CLK_TDC_PERIOD 	: time := 2.4 ns;								--! Period of the TDC testing clock
	constant	CLK_SYS_PERIOD 	: time := 10 ns;								--! Period of the system testing clock

	constant	RESET_WAIT 	: time := 100*CLK_TDC_PERIOD;						--! Time for which the reset is '1'

	constant	VALID_WAIT 	: time := 10*CLK_TDC_PERIOD;						--! Time between 2 valids
	--------------------------------------------


	----------------  Coasre Counter --------------
	constant	CEC_VS_CTD_COUNTER	:	STRING(1 To 3)				:= "CEC";		--! CEC coarse counter generated by the internal CoarseExtensionCore, CTD coarse counter came from external CoarseTreeDistribution

	constant	CEC_COARSE_CNT_INIT	:	NATURAL						:= 0;									--! Initialization Value of the Internal Coarse Counter in CoarseExtensionCore
	constant	BIT_COARSE			:	POSITIVE	RANGE 1 TO 32	:= 8;									--! Bit Dimension of the Coarse part of the Timestamp
	----------------------------------------------

	------------- Uncalibrated Dimension --------
	----- Uncalibrated -----
	constant	BIT_SUB_INT			:	POSITIVE	RANGE	2	TO	16	:=	8;								--! Number of Bit of SubInterpolated TDL
	constant	BIT_UNCALIBRATED	:	POSITIVE	RANGE	2	TO	16	:=	8;								--! Number of Bit of Uncalibrated_TDL (Default, Equal to BIT_SUB_INT)
	------------------------

	-------- BeltBus -------
	constant	BIT_FID					:	POSITIVE     := 4;												--! Function ID of the Belt Bus, 0 = OVERFLOW Coarse, 1 = MEASURE, If BIT_FID = 0 the belt bus is removed and it is a standard axi4 stream
	------------------------
	----------------------------------------------

	--------------- xpm_fifo_async ---------------
	constant	FIFO_MEMORY_TYPE	:	STRING							:=	"distributed";      		--! Type of FIFO; "auto", "block", or "distributed";
	constant	RELATED_CLOCKS		:	INTEGER	RANGE	0	TO	1		:=	0;							--! Specifies if the wr_clk (s00_uncalibTDC_aclk) and rd_clk (m00_uncalibSYS_aclk) are related, if 1 clk_TDC and clk_SYS are locked
	constant	FIFO_WRITE_DEPTH	:	INTEGER	RANGE	16	TO	4194304	:=	64;           				--! FIFO Depth, Power of 2
	constant	CDC_SYNC_STAGES		:	INTEGER	RANGE	2	TO	8		:=	4;							--! Cross Domain Clock Synch Stages: specifies the number of synchronization stages on the CDC path. It must be < 5 if *FIFO_WRITE_DEPTH = 16*
	----------------------------------------------

	--------------  Tree Comparator --------------

	------ Stage 0 -----
	constant MAX_NUM_BIT_EQ_PIPELINE_STAGE0		: 	POSITIVE 	RANGE 1 TO 32   := 4;				--! Blocks of bits of the inputs that we want to compare in the first stage (Equality comparison)
	--------------------

	-- Others Stages ---
	constant MAX_INPUT_ENGINE_PIPELINE	:	TC_POSITIVE_ARRAY_TYPE := (2,2,2,2);								--! Select the max number of inputs for the AND gates in the second stage of the TreeComparator
	----------------------------------------------
	----------------------------------------------------------------------------





	---------------------- COMPONENTS DECLARATION (DUT) -------------------------

	----- CoarseExtensionCore -----
	--! \brief The CoarseExtensionCore is the Device Under Test
	COMPONENT CoarseExtensionCore
		generic (

			----------------  Coarse Counter --------------
			CEC_VS_CTD_COUNTER	:	STRING						:= "CEC";			-- CEC coarse counter generated by the internal CoarseExtensionCore, CTD coarse counter came from external CoarseTreeDistribution

			CEC_COARSE_CNT_INIT	:	NATURAL						:= 0;				-- Initialization Value of the Internal Coarse Counter in CoarseExtensionCore
			BIT_COARSE			:	POSITIVE	RANGE 1 TO 32	:= 16;				-- Bit of Coarse Counter
			----------------------------------------------

			------------- Uncalibrated Dimension --------
			----- Uncalibrated -----
			BIT_SUB_INT			:	POSITIVE	RANGE	2	TO	16	:=	10;			-- Number of Bit of SubInterpolated TDL
			BIT_UNCALIBRATED	:	POSITIVE	RANGE	2	TO	16	:=	10;			-- Number of Bit of Uncalibrated_TDL (Default, Equal to BIT_SUB_INT)
			------------------------

			-------- BeltBus -------
			BIT_FID					:	NATURAL 	:=	1;							-- Function ID of the Belt Bus, 0 = OVERFLOW Coarse, 1 = MEASURE, If BIT_FID = 0 the belt bus is removed and it is a standard axi4 stream
			------------------------
			----------------------------------------------

			--------------- xpm_fifo_async ---------------
			FIFO_MEMORY_TYPE	:	STRING							:=	"distributed";      		-- Type of FIFO; "auto", "block", or "distributed";
			RELATED_CLOCKS		:	INTEGER	RANGE	0	TO	1		:=	0;									-- If 1 clk_TDC and clk_SYS are locked
			FIFO_WRITE_DEPTH	:	INTEGER	RANGE	16	TO	4194304	:=	16;           -- FIFO Depth, Power of 2
			CDC_SYNC_STAGES		:	INTEGER	RANGE	2	TO	8		:=	4;										-- Cross Domain Clock Synch Stages
			----------------------------------------------



			--------------  Tree Comparator --------------

			------ Stage 0 -----
			MAX_NUM_BIT_EQ_PIPELINE_STAGE0		: 	POSITIVE 	RANGE 1 TO 32   := 4;				-- Blocks of bits of the inputs that we want to compare in the first stage (Equality comparison)
			--------------------

			-- Others Stages ---
			MAX_INPUT_ENGINE_PIPELINE	:	TC_POSITIVE_ARRAY_TYPE := (2, 2)		-- Select the max number of input per stage, the EQ stage must have 2 inputs
			--------------------
			----------------------------------------------




		);
		port(
			------------------ Reset/Clock ---------------
			--------- Reset --------
			reset_SYS   :	IN    STD_LOGIC;																		-- Asynchronous system reset active high
			reset_TDC	:	IN    STD_LOGIC;
			------------------------

			--------- Clocks -------
			clk_TDC     :	IN    STD_LOGIC;		 																-- Sampling clock at clk_TDC
			clk_SYS     :	IN    STD_LOGIC;		 																-- Sampling clock at clk_TDC
			------------------------
			----------------------------------------------

			--- CTD External Coarse Count (CNT) Value ----
			CoarseCounter_CTD	:	IN	STD_LOGIC_VECTOR(BIT_COARSE-1 downto 0);									-- Value of the External Coarse Counter come from CTD
			---------------------------------------------

			-------------------- Data ------------------
			-----  Decoded TDL ----
			subint_tvalid	: IN	STD_LOGIC;																	-- Valid of the SubInterpolated TDL
			subint_tdata	: IN	STD_LOGIC_VECTOR(1 + BIT_SUB_INT-1 downto 0);						-- Decoded Subinterpolated TDL (Default, Equal to BIT_UNCALIBRATED)
			------------------------

			---  Uncalibrated TDL --
			uncalib_tvalid	: OUT	STD_LOGIC;																	-- Valid of Decoded of TDL with pipeline of Coarse Counter
			uncalib_tdata	: OUT	STD_LOGIC_VECTOR(BIT_FID + BIT_COARSE + BIT_UNCALIBRATED-1 downto 0)		-- Data from Coarse Counter pipelined | Decoded of TDLs sub-interpolated => |COARSE|SUB_INT|
			------------------------
			-------------------------------------------




		);
	END COMPONENT;
	-----------------------------------------------


	----------------------------------------------------------------------------



	---------------------------- SIGNAL DECLARATION ----------------------------

	------------------ Reset/Clock ---------------
	--------- Reset --------
	signal	reset_TDC, reset_SYS   :	STD_LOGIC;																								--! Asyncronous system reset active '1'
	------------------------

	--------- Clocks -------
	signal	clk_TDC, clk_SYS     :	STD_LOGIC	:=	'1'; 																					--! Sampling clock at clk_TDC or at clk_SYS
	------------------------
	----------------------------------------------


	----- External Coarse Count (CNT) Value ------
	signal	CoarseCounter_CTD	:	STD_LOGIC_VECTOR(BIT_COARSE-1 downto 0);													--! Value of the External Coarse Counter
	---------------------------------------------

	-------------------- Data ------------------
	-----  Decoded TDL ----
	signal	subint_tvalid	: STD_LOGIC	:=	'0';																					--! Valid of the SubInterpolated TDL
	signal	subint_tdata	: STD_LOGIC_VECTOR(1 + BIT_SUB_INT-1 downto 0):=	(Others => '0');							--! Decoded Subinterpolated TDL (Default, Equal to BIT_UNCALIBRATED)
	------------------------

	---  Uncalibrated TDL --
	signal	uncalib_tvalid	:	STD_LOGIC;																					--! Valid of Decoded of TDL with pipeline of Coarse Counter
	signal	uncalib_tdata	:	STD_LOGIC_VECTOR(BIT_FID + BIT_COARSE + BIT_UNCALIBRATED-1 downto 0) ;						--! Data from Coarse Counter pipelined | Decoded of TDLs sub-interpolated => |COARSE|SUB_INT|
	------------------------
	-------------------------------------------

	----------------------------------------------------------------------------


BEGIN




	--------------------- COMPONENTS DUT INSTANTIATIONS -----------------------


	----- CoarseExtensionCore -----
	--! \brief Instantiation of the Device Under Test
	dut_CoarseExtensionCore	:	CoarseExtensionCore
		generic map(

			----------------  Coarse Counter --------------
			CEC_VS_CTD_COUNTER		=> CEC_VS_CTD_COUNTER,
			CEC_COARSE_CNT_INIT 	=> CEC_COARSE_CNT_INIT,
			BIT_COARSE				=> BIT_COARSE,
			----------------------------------------------

			------------- Uncalibrated Dimension --------
			----- Uncalibrated -----
			BIT_SUB_INT				=> BIT_SUB_INT,
			BIT_UNCALIBRATED		=> BIT_UNCALIBRATED,
			------------------------

			-------- BeltBus -------
			BIT_FID					=> BIT_FID,
			------------------------
			----------------------------------------------
			--------------- xpm_fifo_async ---------------
			FIFO_MEMORY_TYPE	=>	FIFO_MEMORY_TYPE,
			RELATED_CLOCKS		=>	RELATED_CLOCKS,
			FIFO_WRITE_DEPTH	=>	FIFO_WRITE_DEPTH,
			CDC_SYNC_STAGES		=>	CDC_SYNC_STAGES,
			----------------------------------------------
			-------------  Tree Comparator --------------

			------ Stage 0 -----
			MAX_NUM_BIT_EQ_PIPELINE_STAGE0 			=> MAX_NUM_BIT_EQ_PIPELINE_STAGE0,
			--------------------
			-- Others Stages ---
			MAX_INPUT_ENGINE_PIPELINE			=>	MAX_INPUT_ENGINE_PIPELINE
			--------------------

			----------------------------------------------


		)
		port map(

			--------- Reset --------
			reset_SYS   => 	reset_SYS,																		-- Asynchronous system reset active high
			reset_TDC	=>	reset_TDC,
			------------------------

			--------- Clocks -------
			clk_TDC	=> 	clk_TDC,		 																-- Sampling clock at clk_TDC
			clk_SYS => 	clk_SYS, 																-- Sampling clock at clk_TDC
			------------------------

			--- CTD External Coarse Count (CNT) Value ----
			CoarseCounter_CTD  =>  CoarseCounter_CTD,

			-------------------- Data ------------------
			-----  Decoded TDL ----
			subint_tvalid	=> subint_tvalid,
			subint_tdata	=> subint_tdata,
			------------------------

			---  Uncalibrated TDL --
			uncalib_tvalid	=> uncalib_tvalid,
			uncalib_tdata   => uncalib_tdata
			------------------------
			-------------------------------------------
		);
	---------------------------------
	-----------------------------------------------


	-----------------------------------------------------------------------------


	--------------------------------- PROCESS ----------------------------------


	-- ------ Clock Process --------
	-- clk_process :process
	-- begin
	-- 	clk <= '0';
	-- 	wait for CLK_PERIOD/2;
	-- 	clk <= '1';
	-- 	wait for CLK_PERIOD/2;
	-- end process;
	-- ----------------------------
	clk_TDC	<=	not	clk_TDC	after	 CLK_TDC_PERIOD/2;
	clk_SYS	<=	not	clk_SYS	after	 CLK_SYS_PERIOD/2;


	----- Reset Process --------
	sim_process :process
	begin
		reset_TDC <= '1';
		reset_SYS <= '1';
		wait for RESET_WAIT;

		reset_TDC <= '0';
		reset_SYS <= '0';
		wait for RESET_WAIT;

		for i in 0 to 1 loop

			subint_tvalid										<= '1';
			subint_tdata(1 + BIT_SUB_INT-1 downto BIT_SUB_INT)	<=	"1";
			subint_tdata(BIT_SUB_INT-1 downto 0)				<=	std_logic_vector(to_unsigned(2*i,BIT_SUB_INT));
			wait for CLK_TDC_PERIOD;
			subint_tdata(1 + BIT_SUB_INT-1 downto BIT_SUB_INT)	<=	"0";
			subint_tdata(BIT_SUB_INT-1 downto 0)				<=	std_logic_vector(to_unsigned(2*i+1,BIT_SUB_INT));
			wait for CLK_TDC_PERIOD;

			subint_tvalid	<= '1';
			subint_tdata(1 + BIT_SUB_INT-1 downto BIT_SUB_INT)	<=	"1";
			subint_tdata(BIT_SUB_INT-1 downto 0)				<=	std_logic_vector(to_unsigned(2*i+3,BIT_SUB_INT));
			wait for CLK_TDC_PERIOD;
			subint_tdata(1 + BIT_SUB_INT-1 downto BIT_SUB_INT)	<=	"0";
			subint_tdata(BIT_SUB_INT-1 downto 0)				<=	std_logic_vector(to_unsigned(2*i+4,BIT_SUB_INT));
			wait for CLK_TDC_PERIOD;



			subint_tvalid	<= '1';
			subint_tdata(1 + BIT_SUB_INT-1 downto BIT_SUB_INT)	<=	"1";
			subint_tdata(BIT_SUB_INT-1 downto 0)				<=	std_logic_vector(to_unsigned(2*i+5,BIT_SUB_INT));
			wait for CLK_TDC_PERIOD;
			subint_tdata(1 + BIT_SUB_INT-1 downto BIT_SUB_INT)	<=	"0";
			subint_tdata(BIT_SUB_INT-1 downto 0)				<=	std_logic_vector(to_unsigned(2*i+6,BIT_SUB_INT));
			wait for CLK_TDC_PERIOD;



			subint_tvalid	<= '0';
			wait for 20*VALID_WAIT-CLK_TDC_PERIOD;

		end loop;


		wait;

	end process;
	----------------------------

	----------------------------------------------------------------------------









END Behavioral;
