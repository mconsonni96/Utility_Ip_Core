`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ZBHfG8anCg0qr6eOwRLKOO7yxjcsN2FoKAwTDFDG5C2bLGKXmnykhjTbTL4OotrBf+2c2Nqzar5r
+NCpyUyhmYOWZJx1tJCmQluyXOdS0RbVaBhcs9bx9TNvuKvQa7cgV/UTPXZB/8TIi6dkAddfY9Ki
lK110Hhq82z9pugW2BBmbmDlFrkz2+iYSDwbVnc3Ib0r9BEdm2thtfYWnS3VwxfInO4LnmQoOlkI
NHwu3P4uIfmVjP0/x2GkNJLVe5E9X8XSWfzdzGwfl8NbpC+LjafEVHEy9bcVOdqRXHNg0ifOC1GN
3zPD7Inl3F+jUgzE/RcgeUGaSMV3e9hVDYuCZA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="aadqdnIUlsP6flpKfJ516EVCdUfvmjlkXC+d9CJBOGE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 83056)
`protect data_block
KKx/DW5uXfzaR7Eru/IIp5ZAuq6EweT3y92CSy5P+AxDvxMDQ8maHnFQP0Qb3IjOJVhg8BaR164c
80uG9+YfISdLbsdiubtyF04jGBU4nyld2bfMM26VdJXijccgHJoD8Y+76NIRbZekN00W4ud7+TTt
QG5MHWKoAwhRITH5wmgcIpk4ZhnNCF2YHeiAAmdkf6Y26fCUC+5TJ8bD0FVy8hD0jYoje6juLnjk
ireUeSR4a8I/qzZcYMGRyniDKNaG/BbnOVIYq7yVr+aAwqPJCzcNja9T591xwXag/cEGk3KlQTJw
Y1w0iQr/EUPIkPPdt5vGGt9ESDxrvqDH73GRYgZUHoKi8cjupydFZPDX59qllNe/Pi8b6LLYp4ck
JYocl80FuGUxIMx5JPjFsXr3Gk84lZu7Ru88WzzUMvV1KcUP0n6sK5xadjrIGRHjcpUdVvH/AmFZ
OD0K7dEXDHngyXe2n48el4eCX5D3rXZZtQOEuaQVbnLlmmFzIwQER7ZRVhNkBtQd9LrlxfVnXNsP
/x0UHhqRZp1cOIr9SAyDrcIw7HwG33Hif8f2PD8xcWxAuQmJt2anVVsi8asAd6MPqznjh9N1vzdV
G2TOLct7fYBYArzzszsH3zifqQYfynWWXeZat16tsQMCvk+yg8YOu/lDTKvQleMrPh2jWJwnWtRt
E5kTHLduuIXi0HvhWX9NG94iuERA6xUOz6NBE80nQQ1nU+uAEnoDiJmuppaMa2Qa1OfOhuq/RqNU
mYicuRfeFP5FEwI/AYR+xVMv8cJr/PpNmYTvusUK2bJWGW0ei8eOti9ugAlDUJnMF1ilR1RubczV
eqPR+f2W1+s1ev0dW2+Hx2bk6o4nnrrSwknblpOn1u6Y93XT2ysJVU/FZoLB06YKPovAuOIF3DAV
zTy9aIS8jQ3R9vKpZqnHmF8ad6ncVt4EaXwouRa+DNjMBcAMkdRoxCA3GgQGvgw31TJR90SAUlxl
q9RA6OlfM1zoE+NjNsJ8reWMqsKOSq9v3/xLhzoeA1XYSpFfiDiq03mT2QKGMkclOSt5ye/DceXg
6hgsrjq6VPVXTZJ6g2g54oGkViv1RfdbPgqK4v9PfkCqJGDnwPIPDE0rt/G3sZr7EbqtzPbekwx8
+TsQCpfmacUGHbKsdanIBYUVXoYeknM8TXPYGl538ruLyPSg3/U7AEZFvlDJIkkT0LUFxVfMixj3
YhWYIxzIlAtJu+mYEImq4VvaPcvh7+0WIEcLmLiMlDhGc+bOQmDAaqndh5ySt5wbTX2ZzooYpYzK
Gdl36ShsBwYn00AO5EbAnJHSpU0JTdIyS8usEeLBrglW6+K5Ho4d0VGq7NLdNUykVt0axOgE0TGE
fV+ejVcNULHJPZ8Rs9ho/IFLasx+0S2wq2QqhoSNkiWpzzNUZjGqIUEdJdaU++7ihlgfXiGuNmun
IhyigRdF5x3coWMC23OVQUd5l6iJrKTn4Xu1lcVcpVie0TwSf+VwOY0GH/Vz2S59CgsZg4JgBb0Y
3JA4rXOtHlHTyikzo642nJZZwZWZhd1XmajpkSZjYRp2rq758DeGc3CMILhwJ6VwE4wRiQz0R7Ue
Dfjx7uN9FmJUo09LNC1bYK5Am+7SPgbxs7yTv8luFaL2/UyWX5eSOXh9s080rVsh4KJOBPKTzyWg
vGJtsTAsFkWCx/3u1N84llEYiyQ3Ri7a80LYXg9Ei0WY/8IhapqC3h5APmSBwmT1NdMzuOv+PTBQ
sLan+hhKFK521IQGWpgxfKyJCsSL2YiHmQ7697M7S/lRWys9WSY2kC9PKWqCH9bsoPWAjfPmxD0A
F10unX8dxiPaDM78+3a6mugSxUjkCLklK/J1nmTY+NRJddIdTil1MwTtnJ38B7Rfuderxd+jy+qQ
q9tFhdSXJhAayJMPPQyvu0jmPtiiM61zXrrod5yNepiFOK0gpp8PnmVzvNlQKXtT2o4z1EDk5jZk
3RBf/Ab07j8a9Xsrv4f0qB+RdERdSOYJB7w2IrVs7T/dA/r9R5NCMwfFTeL49uZAvfvvbpr0T/9U
ruHBSr99XuvsxmvjF0HSCHZQOmJ+oh5rmY4PeWhRFseGBlpEnW7Tz5iILGh+scfNDpZj/qLJjE8N
p9ZvsTpr89XP2mr/c1cJ3oQjK2vk/sfObfJ29alPZgciYfqLmMWDyTsX/vzIndgdsBwohj7Gagot
rgqpKfX47NHp4cqI4m2cJE8hzPVXMWUbC1HcbOcxZYP7azYFPfq9Zo7X0rdsMl9RvUcHOl+XdrOS
w1I+qSzACG4/RLVINP2KQ0Lgh2a9CLKPy+8dSORIir5p8cyZYZ6Rj8shlM69tIV/HquGUFExQpbK
eLToP92nipaJ1HK46v+lu2EWnjXQIoMEiO3zuldmcMG+RX/VqEYo7QfTvdte2qvLxOVXt/4UFNxQ
BnLLzeSsaQynlv88EMRh4tD38+FKi4s3Hgw5OkwlyCAwnIfGuR3Trda71SVjClH5nyvID1noUa71
fhKYmz/iQPiAXAsErQxRiPE8zTXAWlaxKKc33r854+WwWSxIYlWybYH/CSh+TmVDYPpsVOXmizQh
2QoWmL/jcfl8gIXJ98X6Rmgfj0BeJ57Nf1j0hrSq3DLph7nPiaTBEw3NIYnKp6K18e5/PJYB/pHm
Jd/fOIuB+/WlUboG5E5Od6MBFfrOsWEJuc47QSF1W7x6oerDOrZ+Mf2s9NnJNbBSqxJl+07KSbi4
Hi9S+FRs6KfNmgl9OGbC9DgKqeU3eb1+iBHYKjTlsCUV5usJZ58vvFBZ//jjtD0whOwjg7cLbBO/
mSZDw5B7wzcRyLAns+DekE3Kn7go2FXvnZMPaJC5dUPzaJoEhj7TRVFRMOCSo7pWWlNKZLVvU/Vv
QdCG93lKN7j0TEvRMhqbG3Ccco3SVqa+33/gEbU1uYWC359CU2bG3rZnHuHUgEyoQfdfb/2qTf3G
IJHNPR077FvrNal/KQ4RIAg+VVTjHinH/dlf8O+3V3NpMeEfFs86YZyDrBVVFeKzXPKrtY49DD1f
TSKvl75Y8QrKZniOl0LIM4LeCVgFtzHXX1W3bKVAyDyZ9duOWidUSCsOJnvvPY0Ga7wvIgE6Vl4z
RVp5+CuRJgJYmCBUssFkamfqNgYldEbtj5VxmGOkCBlGkDV3i4Q1UdivtMIkstxGVAaR56fJvCKf
L58eKSgnHsWo6sB8BThOi2eCLvywShk8sm4GO6x59GilxyTTJ2zD3K4uBpmPH3FD+nSEy7sO+pNv
BXgXkh/krwdcKEcdf6vCrosmhl7MLosuxsCYNo5bi+21UgmQnxUkUUDlppnZB3BJm+2oe+8T14RG
Aai5x4mv3g6qzZG1EAaHs2Wa7t0fwQAIG9nR0/Y7N6iUKCMeArhfIwdSFz5ije+n70o/Q+LQBRuI
GcD3J/Dk/DgpJYay/ri0jJOh5C5O8jPw+KTshnAZAFpVCF8UTePjkO1vkq+WyVSa+IAuJgr9DJG/
CJQVtzLG8bM1kmIUEX9RWF0kCRqpkUgXxZsigJa8d8g7Qv8fI+QJKe2qO4/Zde4q+sphyI3ML5kB
wexYotX6cCNmmNAqqXYLt6gb8mbYU24fxT2Vaev1YTJ5Kd8URpm3Dm3lthxhkUfB7dcZskcfjbXU
uiDrQFF/9KJaamiZn8WUkA7TjCNIxXP7mek5qI6AHjRFdYBPAg53E4b9HQ1i/ekcOO1Opt9pATbB
UrtHJ8XSqDB75QJX17GbuvS5qVbBBE9qb/3fu3a7Z6XpclFcyQ9xyvrl74dECeZryXrIvkgr00AA
Ffs0uX5AJXLkw2VHolWC6QaDjycakkPhkHVbtFKwuNDS2uiEwk81r3wPRe1NaOdCylXqY7O2azRn
Dm9P/Cc631WrcAeZYT7qoZULZEY0heZbnJkGhJlLf4AM1aOnwVheUxwmGxYfvVg7Rz6QaxfLeBtx
nG2n1EyBqCYQg+bVqFb0OFzRMvsUSC+pv17s63z1J1i1HCrWhWdelNau6e5FrS7ntBNv8sfxPEZ1
rQbWT0126xavJZscymmMKeuxD0OF959TE5zL11i5Y00XoxU+dEyVTT7f7jBnumKRBBx+gBCjiAe7
ys9sCrHBr9y0ghfjY593JHBYPhtHTXSR/BtXv2WmTZZhuaXNCv9yNOUhfExilIu8EHB0D3KcPezP
LXO4NvkP8ZkKzrOLvgqOOWgceXPv5rx3qtOBrG1rLxhy3xT6forGIKKJF39YfTX5uRQbqzSIqXpO
/jfoUcXwZdVnYGAzKCTtoJi2jaeIGavQdsXis04K7mpYgn3eEhgiWzbxJ+oO7Yir128zYQcA8RNC
0imjfk161LmusXVRBAnUfpXjqEmThp+M8iRsrL9EnIwoJ9H3XtJYlpn3oewYJk4jpKbB7pLVPeQZ
F6HGaANNNw1ZYxoDgNRb5djCR+txCOe8iibgyf3SwzwyHxPYLaxasI5n+ZwKd4W9Zu0lImzOXe7u
bNLPspUObVm5wUIPd+3D6iD5PmBQUo1/yqFZLj885vEPoUheg0yr29OmOK0eZRZbT2HwZJl5Nlyp
reb7WzrrxKSIAq1BS5XcU8iKznF1SkOOYJkxwbs3L6zs1sOg/OFE3kbhsXDGw2Ql4KrQhXorv+rN
qA9JscofhrcVPgPGryxXPqQ3Os807GyhJ95OHH1fJF0+BdXOytO86Vwnhr8RmMJvc3eKRZeJ2L6e
gIzom3dy6dnBLsLiHfFZby5dUhevWE2uHMmUTs3yy49xplfjyFESJr92NuhfyhHrnhs8cc+XmoOa
lRb1DD3Ktg/X1kght4BeQ81eZSiTZnYXzIoYc+whDT41JBLb7KtBC0IjfFhifjMHN1FQXud/7B7y
NgQPAb2cNkwi6yYpHmWCDKt73Ad+Nj/TT1xf1GEmrRWyjWSQeiNZUWDoD3Bqi9ANwiRBFjns+4fE
DueuF+SL65i2/yxlmsXVqG0jj1fxJ96UnHqifmGNacLir+S2wH4WIKKn23zrD5iojSvWINasTH7w
hBxCfVSyEEVBJV0Zwf2FiQLCdvUPyyJR4qIGM2O2cWFMnuSYcuIVtT6JoBd8xzViPyRdN7ntdPa6
qR3MeIUF7SmLWlH8TJE4wAl5Vb3sfTX0vhC38R7cQcTv+JZM22meMTxXz+RU0PeAT4ubQK3oT3QL
jb/YxKFO32Y3bTiAEZ7EsrLmZL4Im1Q6zSqJQzzrripBp3XqxoQ3Rsu5AVisabv9GMWD/nOBBMRd
yMP7QOPJqUfRiU1g1/ZXaSd6xa4wwhtuz2ZB+pwLpfRXg8Y35PHx+wHBsq7NLrqs2feCYW/xqEIR
oxR48vZEcYXGRNvWIgt/9SulWgC1XQTP3Z3LBj4I78sDuSL3aQHapW7Orq/tK1g/MsMwv+dgzFOc
X7ASTqDg0B1J3jqCIExD3wa4bO8Ar7zeDQq0afMc9RG9wunWL9sILNgxQmHBQLl01VxUX1B6a473
zPGtVJOQWzxfrX6flxp9tJRmWBnOEAdGREAtKiQYVF7tu0osTXaTwLd/3ilGbr4bq0QnDU3hNhJN
uAlC4AIabVTcDxBYJt5GpGNigp/IMr9HwTX2Kbbcull0njPIaL7EPtpVRP+58B/3ND3fdmpFjp5V
PNnFVC99gMbbK4QIIUVWHODG8w4viGXkGjHUEhC1+EVSac/1CBPpJu/QUUkanD4job0+L0JwQVav
gj3bytIJXSa5Uphzaif2sn+P9sM0E56l+cPjo50gBnNI0I6S+JKx2vVKSItCTqzEp9rcyXd7IDRN
1+Hr/d52+pY5oMhgzWhk5jcO33i0ZToGpFtRwQID0962et7fjkGQ6EsKXfsNu5byO7nECluXRk86
81Dut17oy+Gqq+5SWUw9/o4phz2LyTOLRXklUsKmi+avOvm9iy9WSBhLXm9UMEF2NlhUGY+hbmzf
pkIoe3G2kuQ1uBjylcNje9gJFstfcsEJxoBVz3Nk9t+zol8hCaYyZLeIRjuStD4XsGiq189xmtgl
ZV8VI5OJ6qbUMs4sX7yM6XFTvfna8zljiAoBC5LgYxhFyZhhmU+284nhvHPOcYeKJE3OYrUrJMv2
/DTqmpYd05B/9O4GKIg40PiCK6nKnYCWYRTq8QS2rx/DYllGz/keqG+CGS5HG8rn8MnPl+O0xs3D
La2Bpad/8I2DLo4kniCw1hkjb2o7BSCjQMP2b9bR7062bLebiOw3WeV4ne+vLM1y2L5KQbYNZYB7
hRSOqi3LPBYrvc8PXBdS50//qQg4cKy62eGwHhO3JmTmmysv/Xwa1+gwv65DqjjIF+7urAV7ZcTF
H0x/ODgfqWD27I2GZVuQxuZ1cxmmnswj2tG/5QchO+dym+TrMlrtXq39HwhJk8FbsGGOV8+fsKR6
3jGVkDKmWLfWLzLtQ3NgQFdHMNNqsyreQ8E8pPWGSh2qlNST6gbRhQh456sb33zkab3mrTXmVQMJ
eVCBpZcMxgKYnr6TYAQDQ5w63PELHsJj4D5JV0htJVYakSMXD5NID/lRqS4e2/VmvoT/myCASXkn
z/Rfb1tj0lAtEiVO0ipWGBlIDlE8ETmtJJhChDTnUG3acq7P16htIbzLoLz0tG1askRN0mLJsVNY
xnwku6ubm0RXi9ChCyks293mjBruFu87ZkXW+eWNbRpu/O4gdpknGXC6ZVtH1WKyyOACCoy7VS4B
JbUPKQueGDocuJWiT7qdL0i9DtQ21b/sOSdqENTzlBo0P86tJEyEiDguAQm7jF71qMmHizmVdGJL
xdh8YuV+A0m3pmqS7wzCTSyxz3YrvfTjMn2f/XoA2UmHJWNrCqCVItZHGNeiP2JqogdEKwAgcJNo
TXLYeEOfMjOTsGb5BJIL04Kgqv8dMCSUjh7m2EFVt9mI7vrQ+JVgRj9zdouGqEFcWUZLXb+YG119
mTsL9pDNbn3dLdeUg7yvmi+AnWxVk4YpGt/jYdTskIxzExYVSBbD+dRaw93kqhmBMBQjSiUHhx9B
yRRJeqs94390u1rV4B/9l3f7BtFXhD3l/xqVLB5h1InXPohOELwe98biR1xLw+VPpK8IpMUdy2Yq
aF9W6qZ032FFIMbK5D1eDgYLBX0UD+kznTFmaYsfFckgxCzZy0lquCF2IJTiGeEpDEt7QlL2KkjW
6fqvHn+WdQg23qVKEWfCLKCj9YCu7bxU1uK9PZ6tQXhYUgEMIue7T/U+50wyXtIduAt0D1SYm2nM
FgeuxyzN0gHPaWplUpYNxiPjvcSc9IqgXNYMvY16SMiVa+rHVV4e8471W2Q9NZ79aYkqe0g+VtQm
dzhCPTmWqNvd7BBCC1T7nd4jzPRHB5CVhNaGozjsdYEXxW/rv2Of3mjMHfIj7FT70iBTDQ5pOaIS
7J3U+tLfx7WnlJtOaRKQiSuhCy8EqYjMj9D2BHyvvaI2qxCCl+FmgLtUBv6glkp81Q4yF0K2GkgQ
sl3YSjQObTok0M7Dga2ga/eR2EVqWmfEAo5MOYqAts/qYegCsKOc4XuccrE1/fHvgS3iyw9GK3am
6HU+z6nKuxdRiDkBKi4Qsa4WpxvmV6rfFBqwWAiijPVlHbhR/BvQFpfgVFTpzAoKHbb/BYgNQzMp
CGYonfKUu3q0nFoLw8AJ3SPvEbePtpzv+bR04zkZeOtNyykuamOiOdxta8h8y45IhCIslpuPCWLe
jHMvfpclEWAVm3vXmI8bq+DmtGdyyOvOqWWlkeoxvstKg3jwY/lPpngDMaVS92uj/v4nEpagxsGo
hCQ/QG+sut0n5JACkFVUR36Pp2bgEJz9ek13CJ2YBZRrXIiy6yRXQqOjeszfagUYVsHmmryZMU02
BgNYxIXU+EGL857gx+cUUfNh5oa2a0enbRaWsPR/Nb8SYssdasZ/vvkBs0KSvEOXTBjrlPdSaT+4
oEY43YmQG0liXZ88X0R5Nm+hGwIhr5nuTp8SKyVg5JIIjAjZJPDx0qOX2vjoNHpKkDkPVIwACgZR
AdstYoJo3vU3szKJy9SKvXepMtyyM5GqVAhDq2mSVFPflkq+GwnGaHZ3E29ebxgIES9Cr8kQx+pE
GLhyPXRKDCpw05oLDPSvSGeuYZMwQweM0txiSSEQ4PxEGhKB03i1Ybw2sEJTCkVsIFVeCFZRF7id
XM/M4BD8ILEtPo4fbXa81/tumQqMtZpJ8mR+gRslWZfd8i9o1rQzqqT32tbCsTMbyDyNqtO9sslU
TalVgG+1Bfg5VKo1hSbEeBybwclGU/7AWpMl6s+E1KRjUQzLRKkLslx2/ENrn43tbs1+MNSmCQSE
bASWKSEc2+ysshxY21Di9HfY1QI8ePb4w6V5niwoIT3mSBSmMTrl23IAYvMTVjOrcT7Qr5GmUNRb
aTPkP4YCA6pmdN9TzcBCdmCvijS+LDvZHKpqSrE7SayFrds8DRtIPlwUqthNYKesGWkkaW2DCbVl
9vV1Xz+ivJwJO39SN0LwquW64P3S7byPzLftYGiYWZ3BB38c9vjJvO5DeotY0XLgTiOoWXrHhGpB
2/lzDjvEdeNGsD5BvhVcWAAk8G9/RVlhIBwijHejT3djNRliw/+T1HH37yDxusJ0cq/c4uxpgjho
CptNHQSLIsic8FjDo2CvIWs6nRz+piTAliOao4POOUFTa0pPNz7e7i7MbGai/QPxqQw6CMvZ830Q
IN3P7PKYQiCyR87B9cgdoGZI8ennGWz0qP49YKrKv8nD/cr4pt1rgTQlZBM1FcHV9j8fQNnalJkf
ra3zu1670noPTpYoJvB22i403N84ZRKvPW3r5Exi9wkqvkxofvVDIpnatRQFq/SmlEcq5VCQIAW6
8aJdA1QNXWVp30lHndnKjAiNkCQ+uC9MlhU5sde2+TGg0tHog4n/N8mLS2ereJhohj8rCkVvRtn8
4Pg8I3GHw6uM9cc+Hoq89xpr78fCkbuejiYauBk/ONZ8ItLQT7zemlfnXLwj/WjufU4NvaaeKCA6
42L9HbHN8Z+rrN0DKMW4w4Zb/cpVQT2SI60LO8C4w6cFNciOzwfZD0QvMrEZPkoW86+9r/4QUSFG
fnZfDX8sT+ET6BEabQNJy7AsPxqe4gDUZX9BkqoNzIZw8L+mQ9/4vWGNMzsReyKbM31TX1dcSYSF
NBjUltzXb7kDjOaiblS1P/FBaoG0z6pgx4E0/zSJeHQfeUzPf+QqmjmBaktyN/M67Z0wU8AV99/u
ZnAWOVw2faeXZyBUyJ+14R4j9Wggl1DcKCqwoZ4SPCpG/smw82UWUVPzWQXEDa3sWidre2U3xKFQ
FCcJnM0XG2Y7m8INf/7AB5iHQ+DYmmnJnsD29SmQOtjcWYynAH5eJNRH7Vh/boV8GobyuW2EFIwT
GGCIrU7692o4is8B44zsAH/vYZSe1qkzcvy3BRzh3FUH8UDvgYJWoOil6GiDKsS2NEfxfoOTuusU
C1sXn/FMyZwlO1wTF+MTQuHkG6478JGOVY9RjAlmpXzGsYCw6I+bH/O9AzJ4+xah888kH5FUPVqv
M8SPUg+PDHI9fcg0FiP78A5fP9xX5a5m8yomjsSEDhdds7dGzD2Ko4B7qx1VW4KP9Lm1deFOlGwq
Jd5B2IzmdhL2+H7Av8xXuVBR9XliDI49vBRDXeTH3r5i4kic42RErBo9uRlDZv0KqPcytHbLnuVJ
cZJkqK68tGjWMd8A1mDdZBcJU8p22YuerY+9UAbp009xq0In7xI54Vt21s9bRwAyxnlgx6yrboSs
x1s6Ao6sBfPxfO/0EITjQH7nT8utJiLg2bkSvc9wZ352NY+LmhgdwDRZv+DePztlTdZ3+4pZwd9x
iWcTNCN6zX7H+EwaVZtMABCDUEOdoa1W3cHMXjIfVpXb5Gge9TuBDOWStC93fus4HZXRWFdleWbn
nPMXF6PhJ1TOZVi8dI+VyLcPW6Ue5du4z+1QBGXRDO6omRSk/x7j7DZkCR0SX3Jyjcj0o+igjxaf
GQnWCoKjkfi8aOXCSbGSLDlgZ3gi18hYyL4GfxuWQMlGVZAF7AyKU7Cqec6lg5Hp+/uInQsnQ7/Y
PnYihev3SWOvRbp/GHLa2wAVdrtSlJXF+b8fTpf6rMUUbjyxa+ZsnxOljhPu5l/Z8ZGw53mdFBVM
kKb5PBuj4vbShR3tVxgNkwIT2bec9xtwkaRc32xDrHejhtRsAdz+ZJYh0JPFoA3izn9d2qQKNnf4
4detkHldlBAI3i4HLCE/rm+z+gpNuL8LWG3c2+2yU+1miv6O2lMqSPEMU2IhDvBOq+XhlTn5LF36
U90QFQcHkfm5EfK+J5vhjfrDpc21bPlxPyztvlt0Z02mzI2/7a9r++wmFxbE7+WoI7T6cpyPGDpN
4+6IrPGjgFstGgq8+9KcXzlQl0BvtCxCim+q6F4iuyD7/luy1nh2KE603rvX9FVqP16cLhB6bPt8
0y6XlMn6xBzGmcaGDM1yxLpY5j4tBkY+qvf2X7ybx0clM/v7q94gssjuOQ9/l2HNggbD8Ajspfc1
AmQWRJdeBIK42tCU3g1z7uzmVllTW9RSiaW0nksllDHFW83lzvaEOJVsNP6fk2/MqVtXgZhbWGqy
8RKrK8p7Ta6eDtwTXf85h59TQamQ+47hLAzaeuCjmwNVaxmT+VfAXXQpxOI764RngW99cvVfsEEf
T+LObMC2LPa6I4CMtKuHaB9ppcpjJJOVN6A6YEf3tbta+e6O1JM4REeEl3ph31YAHynHLDj56Pst
O1QgCddGI+iN9XhXrHVmc3YgkRy87hQIskrtIIyEEejAcTyeUif3ux7olYWabAJ97tWCqFTojCB8
I5//E1hsKg1WcM1z0KBtCm7faMS1L0Jvhs3VucLnEFl2913DZCp0t2RmZKC5/5Qo4wK7Wza5aiO7
JR8Q89fe7MkPDSpyBVRkgyriIKmGvDEdiA9at6KaNhZGGyXbtmYKvHhyokXJdZEyAiIyMPA0XLnt
qGKtRODstVJ4zdXA+pcwbM1+kiRHtS5yK2MZ1rP3Gyh1HoSmqv0ooIq0Aiy4zgKeAmryDrWF7+Hv
KEZXyZ5VW6tAsJIKrtif30ng6vNK3RBRL/uJqNeB2qc4RwXdNNplU+Ao53V0D22cHm957J4KsE50
9x41jBZKW/KIjv83e14EZDnB6Hf/CMxIlhNnDcaa64LEMUavoC6Tjg3ZPGZhHpu6OFLUOsPXy2Mw
vLkQYNTLqgjmkMbxl1v8uUbJkRQSIO9xnWAqxWYLH0EmpHUYPzqHzLh35+y/oTJ6GrM/oNKEjVjD
AtvONaVhPiltLPWM5AN1rTH+FspkemDcF02UVUkvfAspUU9RxudOwRUk4LSdlEV2U54CLPan98Ox
vK8ZIKRHZ07ygmvDj7FFqyZI5iJgKX1/HDipICdW9lreCAtEl6N5u0d1cZuuHq7QPUskWq4Q01fw
cm5e/uRoXa+uHffU2qE+8nvjUeDMhYPn6Wq21TrSChtq9VoI2LNqibh8bTI+/OoIUOQtOjIYjCCy
amBih54sUUOrwBOqlS2yILjaLhMcBZSR21B2AXyOhotF1KhrsT44xchHlcusNBrS6s/d2DjMOJnU
ZY3CzGCGsYPY9fwhiHXYlSoGRRuLQPnsfPKkekUQc1Szolim6OzqlDCDrf3iZrqRbrGLgFqMP/G3
qta+pmNSvaBMzS4yCTFRatMs69ZoGmGlQx5y4wwN4Qf8DvE2VopJdH3lzWfFCpWL997MlOWVb5+I
+CRCZkbYFkwatO7a2rPpo1uQgVGs6e2Sxm5G5tY3HGeti3bPtAB6Ql8ToH/4gu/fXECXhiXhkObT
kcNXcWzvh3UStZ/fpfOBsmJfS11wLnb39MecRrjiEixb7AknfHzZKY6krzjFHbLm4N57kwQ7JYkh
rA5ZzL1QMTwOEJ+z/nEwKcrDuHltwSqzwaNgCbS6tUqk8iNJdeVOL4z8Od2VcqTxT8tPszgjrSh+
EA5MAJs77ONzjW+6vSdlW6HuwE0JhJJfcYeFnV7u3RPmaUp0zBNKKzmWw6OmE+M3oEwq2xY1iKED
DBoVHa47DblD4PS1aaoQR+VZHNV+WTbvNGUIsbVWl68jufELo0bv4RX6J8mtLXSSKFuDZ7+OQwhj
Jqq+eFZgmmN7SfNbA9DLmwaOAKb59oDRx6nJp9fxB7TkEFD+cD32r8LxHqN7MsaBSFLPBRUJlqWh
GS9TSe3sJv2CMlU7gsWEMqgjwJ39pv9swxRT9xDQWsKJu2geMIJ7tcjeXHyXz4iy5s8mLqV6cevj
y+xBvOmfvTfYC8M9mJTs8nhQE2VxmO11UlJF603FxyL9JPHMUvufEzdBoioBT/WBU41XWWRq4xFD
6pLMTrjLlNtFPaMi/L3Fa20WEMiZbtpoucGs92SNFCOqaMsrE4Qnuu9v35owgbYKGxA87PPFGooj
CSUKnkDsuK1BvviKQEws5Gcit1gJdG02QkcwVv8vicspiRc5kqXFF01/fAHLZmuDdAHZ7EKZHPSO
dLlvVkV4kJjRm2WzeHmtalign53FLoIHe3kO0ineRD0+MenrEHmTsnu4R02vaE1rLN7fCKubM4ic
Mc9wxl/fukMxaZjbVSx09XSlQi1KFN+Ze1e2lnEJ3xYegJHUwfKJg/XxlMT+cjPuPgnJJVbqA1gl
1qH+9oSrzcyvEABK/gZ2uvaWN8CdQaPJHnaHtBsc2lBPXsY2U13MTMO7iGg5zm6FwPgW50xovz5P
OaEmpefy9B9LCm9/JODkHHbZrHGdz4PacB3f5IcJRezTstH4XKMNabZY6dT4PalrddiW11JrgHet
I+pooCYqliuABE6QhCYJs8s6noUJ73VNurZrtfpvI9YQjKqcBxBZYHJ7WEhy0p6l3TZQGdiL3frp
CbUKnAw0++ulkV9PeB15WN78/4+qFKld2hEHmOaVD0QDN6PKvAkbMGel9oaqJtmc4syDlXfsDzh9
5/YxRi8VolwD61CBflQXXpUrfeMX82x8qvkXTo9OHiSpKY0WsaKntWXGlOsXNULQgJKd/qeav66g
MbJy9YX+GTAWrMUdxlQ8hbZW19umZ257KDOFmK1ZeWaogd4s2M3GGgx2CGFHjz86VVJLMlR+b+Np
7uCB8eEDYzszWBqeaHRKKKJOFAcC/jkmsPwkLoJYGWyMVcEqQozzzSCsaHvIgBFHbc2cXMASbyDR
iyud4DBEERk2zoByoMhUNNWD8N/Mi6PlPKTbcvfI6i0kg3a50ZBbyLbjvfOl7+ciRe32HiXo62v1
Kv8+eBhmCC59Z04U2i/fWY0yymXUwKHDFFXnHey5l7oihhuxbKNRGzKRznPJWG0QqkMBID4XGhcQ
nARff3rNSPGSJHBmrm9c4nlRQYNAMx84kyqi8JWMxWkTTpPpj3idkiP7t/N9KBQQh2gJ3zf+nhYb
pn+P+y/MOhTP6HkBb9JTTAaCxW02+4Ff15ivd+n1XjlSpDEYy4rqM2So2CPwr/XbJ3VD0YyDZeHe
TO1PK9VroU8BRH9IkB3/R7JZoGtSN5nGl5VyP7zL9XIpvXJXkG65sWNuIXTdMOkDzjwhDCcJDlKX
I2mQIaFVyci1NtsVkEWt8dJDUIMRNlkc6MLsuSvkQbeAKGmygfbM+wM7ZPmp8po+0DhX7DjxfGcu
flVvliFrYExwVUyO7UIFXl0iCX9gfjYPKjjhYCrrXA8sqh+BzDSy9drHJwM9mFh/YfHXPNhmiAkU
8cBn9kTnfhnY9kOeCK+agMp1T2mtqaKfOkQ1Rmv+ri/en7pr/d4MlJ0UT83HPALZ8vf/mT2voAwN
CR3CA4Nrsc7jjU0ztFbpX0DPXHDgMSDPcJTIz6IIjewIvQoKQnt/nOTrXJvrgTwGXWZCDwvpoXxD
cUw0JmznZlGrbjxKOYIuuN33GNVbTmlBcAhGdSCRALiXTVJtASIAPPClLZKGeKhvful2BI4SgZuk
+/f6FumEN+YAmt6vIYHLdZl1D/JhOEGzzIgONhu2RkBEKVE/koMXAAq/fysmyNkO27DXBpht+tdb
RU9hRCXjL2y1FPdnDvNbFTwwVb9X/v56JcFOwKzglSSiRBl+YSdNucrz5zJZJkeYj7pjuO3TaEZR
QrhKiLN1yvznvYhSadrTWwJpq2v5MTqDZjS9SdPfOoxhSyBjcdJqVbvL3/0jDYsNJFGLlqBwfS9m
28AXG1gjUFGsCikyzc7KNG4/d/rpCGLP7MKw9wFZiIUH62dYSn7j6Dixz6kJff8cU49z1M/RptYp
xJvFsCBTHvW5DhSncLCKCoJgNkOQTbmkx1x9SMnDfwBtPgDQvZJUjAv6Lr7PHB9XMwbWPJ83DHy3
iJHPnLBucn9Zt4JMuAJ9jrZ+Sv0f1+en4dphS8jUVziXa27r8lzyu7T1vK43sZqxoC9zeNgbqHPC
FMfA6FQubGLyz3Nnc9KOANCeJVebALpJDTcUwQbYVlaQ0zeD203MNZYFwJo5nc+nVJFIRqW9BzVc
Nh2Kv1BsUIReO0LrGwusGPrISDvzIqZZ+CT1u0eoA3Ufq/7CN87l93deBYGaVht6EYx1HUV0RCTZ
D6TgY2P5jKv3LwW07XsQd2mWS4hf81wMmUafq7Ynmm0Zr6GE57uMapPVRsecnjvhxXW+GNc3MI3E
yrifiwR/7MYWgoGwOrHJNW3GtsPvguLpm6bsv/+8T0qVftS1MTxA+HIGY25zh/Q/vGywGxsemYx+
8fWP7Ja6AMRV4I46B9kmX+HEqEUOAKy0shV0N2RP2xA+sZ+ynNnJzAJivPYAUwo8Q/5ijI+yCtuT
rcM6VR4aUBHIV6zeXVWB0qDXdA2Ntfp/fERlhasJ5UJJIkR0FqlCZqAQYHoRbeQ62DYJZgXhFpc8
HUYSxm33Mi7b9/vlyUo9ZVKk5/el7OOnQoZGQa27Kl0uJABrS7m2Jr8T33tF3NJpKTrTm8zY9zt8
VVtuqn22Um23AXg5/3M0Mg5E0kOsUo/zG28C6UdLTJ2XSt9t+JpMVDklNaCezDKA7FJm6DYXIsyQ
EzL0WOt5fCSBO2Ozy/jiFSf7iPFpQTTyF6upsNoFVQUECQbkHwCbefzkD6g9lGVus0W0WLwQGwKQ
Ej9BjW35RIxNkenrbt28ljpaLpVmrxZi+j9MqNFWs/V1ea0Bm6Qsxh6mjlow3K2DynCKyVLcaEXE
56XRNxYV7iWnkkrn/xCJ0A6GkWgZ2Gedu0c7ECv9OD1WhMotDFG7t8FFdiPycD7i1bQ96K5+BCt0
kmke5xsyvcHa1Kb1YRFVc85mnL4XtFVVaGuTms35vZwX2yso1gpn7k6jgnNXckjHmmAOS7TTVMoG
YmZNhVKESrd1Uj7RY05gnaE6mbOq2xHrAaZXonDP0F80/hFdyJrRxD/EcXC7FoNUB7lApcNJiTU6
Agu/gWu0Nzc/ihZ23JwJri8PNCDOBQapt/Y88jeRaSu+TPdWAx5hR7KaB5nD6EZ1U83Zwi2m2MRt
Z3hhinb0/TlpUxOPmo6s0kLvnsRgErzAyAK8tGUM7fsCx/EWSVMF6CsCdwMlIxZQ5yFNle5jDbuw
X2Cy91qkp4f7m/7y9Wc959CoKgusx3TR3V7KX14/MBnQ+tBBvRK/9MsSziS38lwarI230c+BG5T9
IWP8PBAHiAaYtXI2xRRzzfmtMeXMA+jr5SOaH4wEJio1Lj1F2e99cACiFR0Kx0Po59oNec+PAyzF
QVPB9ZhLQ380YzpopHt/pfvIhKiljbdqxLCmE4UZ2CYPBnppE4xVLapnJbjoCEoFycyySjmFe3aq
WXvHM8tMFaiZ9lC7BHrb7ycqH3dWJDmR4FQV3P4OhonVhlX3sU5wbR8+5dWvfrpf0mqCqxSbu8rM
E7VSLbbED1AHRbDSwykcOw0MS251dt5lmJNJleoV5KRyPDpE6t3nL4wUgltY4M1eMWrShXF17miO
EXSPV42tVLEC3p1QOYCpzmoMYh4SexJmU464crmL5LIjt2qjbARiKEeOzwIgu4anxNRczjZ9qfs5
qZzdSsVuttipx0lOYYiwd+0eJdZO/MXp9cAm4c3F2yknFwg0s0s+WVTFrDDDV5V0Ennm5bcsIq33
ql4vtKpSA8T0Q7TPrWhlb4KFZdpdOYrIJVWXbe93BhBKvloqL+EEJKmY0UtVKwfi/qp2KRFuYfTE
fv2vRIs+k9hxBa7bXQt3uk05gXfn6LbaIUbGf4O5JpW9NsJ1jD67G7NBbnIKqirvfHoGjCX6LP/F
X+OTTfo8cG1h1UpOQ/V08O7Rb3YHBwSHWkZiepKDbpTZ3RWNLIRpQ2dOfPp5VvZAbGoXrPiKShbY
ZLLNatrmFRn5ASIMjTHMXDU5bRJ1AbsA8YzfH0FPrzNEXlQg9w3GnjD+D2vkQCurcN++PdF4+WkT
kOeVRQ/EtNqIAACXnQfg7H0L+KstaQ68/OzOGfmf29z6h6eFcML59XA4MuNpJKY/V8mH34r6nIiP
WK9jcWL6Sea75bfZUnQ1kZPE69FM/pgLCavRd/pyxHCYHnNkZOcM21l7tzv48PDK8yBebZhVm7M0
vDvlVy9T+MUvKdwVvifDn9dS4y9oXS5rUh2cT6OAAfFd+A4ax1eVDYcZ9eLk2k4j6G0zZs9epAm+
e7BzS/IcfoHUGEDpvgra210IxEWE6UcigS6iKUJL1FqMQm5SLq4y8MlmiTXmDTwHOUBns7o0RIah
cWibOv9tm5kk9M2cm8v7LVo5ygBG1SOIQmE/+Kdv/nV3yogu4Xk9v94+KWWYbQg2i1NgPyCYLjpB
w0pf/rq5UE3VdWN1KA4f7uXqisxdOedOLikWwIfI/hNaRiGCQHv4ayLZC9BMgjjDIoLKRFkJQcah
Os1JA/bANxFiLQ2g/9JKppvVLJ0KzyvTzRjpnZAPywtOhH2RvC1Q39+cy6vMFBwdB4bv0/Zfvh23
wYKxk50/SWC/2VzzjYfC0t/yhgm04wAIvyg12tCv8HNR+abgEubMBwtUa/v9HzH7ez7Q8/F0ya3g
pz7oA2r3I47AFQeh+1i9yeDaYISfdWqiVjuJ8+zu3lGJsSrXGT3eLIsG2dE+8hHyJ8LCPT9Khp5R
bebNFi9fo49dwYuHRb0lKORD10U2lZqyyhB37UY8cQAOJV+3NGf2UuFpVbWldlZCVbv/ddPPXM6n
8Q0H+zhIL9rL2eHxaltqA9/k+XP+kcSW+0PJ9yv46Lf93pptgSR3A4pLsmuNcRraBjQaC0xZ2Pqa
3qWgNffmEuPmTe2VakWVKPx+ALasxh1zMYuiHLrtxquKOUTgw4OE7Aj6FAo23KThGQW0EGdHrQWx
CJrj2fMWA99ddL/j2LQv+PbyUal6SLn2bkGZqOQim7bZ6h8AUJUONKk/kbx/o3fsoTvm7W340PZO
d+486A9UKlvbc0eN3gRChC589r6de1dYDh3Pl0WhymciKVJgKDgEKrWHPZ/wKoenkcnqMUdE2Xcz
yTKSqM3tC7I9jDGs6M7BdLbz9W7hAPpsKF0OyvBOoqZh3yKpn4vxaUqcN2wKxn0AlUNDsY1J4y1P
hbk4NL3x4Abbj86dSl8hLGrBLCXatyxus2E0bnE3nwU0OU9wcAxekpXs/dtuG0JwoxdS7FKsCTwH
kZVRmNyGI/ykcAlL/mvRPmc3USQyjBfUts9xW5vxhncTVgdeveqTAYxeg5UHq3J6KItoPvuvQGDv
1kVz5ot5KstRB0f5DFNc0FgeAUEu190p8B447DLDDd5aj1jA3Stw8xh3wQd+EIziSg3E/h/1/3og
5e8YhRaAFTU7zqfngz3r5+k8t85/yzhbwNwy+V9yqIc+OuOJS/DHEuWy87wIl9BJgWUS9SHy8ZO5
Z3o6pPZue+j3By/9rmDuFqt0wDbMHzRMfqDeAb/Qm3tEeefI3KtdZDBSCVpQMV9qsW4e+IrN9Het
0J1iS5P/2OmOxSv14BJUlp0Y3eBuLss72L5TxEmUAfDCYVzGNjB2BjFiluvR6UpP3A0xg2nfHbKt
8eYJ0RJQweDMYCt0tgXA5q0omiPoERfS/b5tb/zB107WnWcRn3jM2AtFAC80iuOWEYb8Hxckosqr
ljGPIupA30sNIcLIt3QzAztXS0G0ZcujHybIgWgzA5SkankfsqhL/Lm4aGKsG3x3iX9NB+FXsybe
M+SvaS0ofVRFvgTjs5XJcJG4qsIsNNUBgZn/ztXO8fWtZp7GGvXszJAS3grSupnzcJ4Ehp/21vzq
FsHLSrBEK9EnN0bfkgCkOl5ZGSreTQgKZZcRGeo1MmgOfADA5fPEQlKj4eGTdZOsb0JHIJQAwxJh
mhVtlv7BkVlpdR8HcckVJt8dQv8r722m8LhGoHpxqkGUb7+f34ZaxugplMrj7wEUfKjt0i+iXhIH
4qKFkwfmT4ZL2T7/bAqCZ+awQz2rs9OH3h7x0Icz4ve4aPWd7/55Lh369jkS7FnOUjZlo+1E5dHV
Pl/0ohDdNpwYd6Mz5PVANZIasHxp/NeCdS43uIAUeCX2kdq1sXAjYtxbwOnFGi9295tmO34KsYUl
LPu81R9xYPI7jnmKWYPsf+F7cziPu/a3HyotYctQxr3IpfAozxaagiRoM2NA46kAyOFGy2jYzkCY
CBKQrwoROJ+iZ/qF15Y7RTjvWeSzEsZJDNww+pY/N2ZTficaxMB2eudFumsDjLc+tJHYfYtTpWU+
S08pN+d510FpYNKPjAY6HgNINu5XTWwWW/yUoqDWZE58pxjNEC799AGuwbooE67FNrmDQgSmNTEl
dc3Mp+ln3Fa6xQPIqwPN+q5JQ8s9XVyy+yCsc4W2BBxreIKeb4x4y9dKBwoedYoTWZ4l9k38+uev
MHFU3vnae8l4FZM9BOkJZ8wF58u8pqwMzQ/gq4kqA2JrozXYbC6aDzCG5i0Ietc7iLerPjKW8b55
FlTNULSN97JEj8rdijmDtZJqyYCK8XErSJyKDtCtI7qQuF+/LDjgBWlDr+KVvcY6LRJSXpjfx/bG
LfDyrwZXim8uVTby+16jSkMKVLryqE4ZUJXBXPeone4OBKRnD/9VrqOL1GcnQQW40Xkhu+3ZIhI8
vzZK9LhAZR7uG4p5WnmR3dcqxLQMGiHiID5IzqZeC8mGif3yKovLCUd7eCfKDk57L3G8WPWBC5SK
8dWkTt2AK36eviMyg2A9vhSy3AbDWNWakluleL45FN1IEw/57pHczz4muMHDdA/Jw+7LE+IF1i0j
qstgvICFxHGmyuHXKUZxKOl2SQUKXkzOb/C3o0mUkvwZMCrF13DzSUTQA6xRRwSMWPU3pATKvDQ1
9sR6sorM6PowXYMzD1ZDPhqKqfkgIg3Irrl6w7I/iWFKTpS0rU1LW/YhD250BkfsHLeAaATtol8q
fZVoq+cwXbK5cwwJj2FeecxN7h2+wIr/BpAcYWpovKbTCK+v+2MSsaOVJdbUebN0y7cJa/YlJP4u
L8v3SVjudhpYRBCTFpOR4vLnRODA8i/Qy/yKvsQrIJwV0ihTUvEZmnaH78CH4DS0yXV9AdLuutwN
tiVlsH/zbsOvZPB73seo/6hlpx8DC73lg68O7kotBqRNkdVbXltcAdyPB/8ZBzAoFZCjgpRvFwnl
WgmhjLG06ET3CRgFzNn11TxXsLCRqb5ymet9yobx2lwmxUKqJtMH6LV9q9UXLoI4aaLgVp7ZB+yK
uw3qlTmzHoHak6Nsm8NEW4L5IOfD3Wc/ofYSFF2kmkB7VTIFKCpvxAoIIiHsnaF/rx2exwmulUb/
SwvgIuxfB+HjevbvLT0OBvU94Z6t2XxgB5p+tywFfR8hQYbSVxANA+kWI1tuieLdkmhM3xd+6ak0
kf/5AN2uAdwCqSmossQoeK+T+k/ilmqp3eKEKEbXTyINgMFXZo0kwOlPLQKTPE7rYDuLNEOmILtC
ChwopfjI/j1Ni7gQLWXSCHLjHbZBHLtoxkchkg912mKk7Sozk7Jha3yAGauGdQ+gz/3zEicvainL
yb0rAErlkrQp3hxBS00c5PQcHp+K66d9e4f5I1bsabniDdVLp/X+nNgd4Oo+egHtFC8bAAEVyVtB
Jc24+WdKJBxaTaxChGZnWonoX66RBDiWH42+NwINAF22R/ree38bVnxGCzslUn8Iq9zzEWMx/SfP
5MZ63H+PsvyptVdY3A2DSP9813oIG+6kBcrJQYxDWj3T0FocKwR5YHm00jNvwVAadq52KgK7UGxw
kR9E56EiraUPIob3AT1HRnXp1iLXnvMXXN+uWlQArAFi1l15RwklNAmSKpfqOhOXprFDXVhfB7fL
byom7xWqVDHSkiLjSsKwOZR2QGOCFSG3AVAdpjHECemvdGTeB6Qmbht460LrtbFKEc+TArQmJ1L9
AfA08D5y+GUOuW45cqNBJiN6c3lLqt3ftSj/+YpyVfzYULGbCwSaL42nBM+qxjv8npameYhU8sLJ
5QSjy7puBgHO8kWE0bLsJq7CVlW3Biu/8CkauSoDESrW4UqnVKL6WwI6LgHlORT4Vk9oFDk1yS2A
ljOYfjryyTa0+8D3Q6E8szwMzAmWogcjazwDGOp6C9heN97rKDCixXZt+QtUm/BiOWktqHFnw0YY
BikTflckaRZ8b/iyigRwaEBVf63smNR8rFA6J3bkPEgkZgsEbQAV10XXjI6bPMXeDAs5eAvHaAlk
N6Ve4jJr0HziIW+Z1671oTQLhygZ+ABarta4WULuoGmLywd2GYjSF1P7VjvOCvPXYg9j57Yh5Jug
MtpXhg33HqGaVS+R4MauoDZ3VxYNxxSofByLUOFsX229la2wow/+0zxguqirsWZlLobxopNSDmF1
CVg2Cf2UkXufldhH6s0E9T+ylL+VAXvlONIOR6G2QzODH3cgG2GkwyoYvcUqDnoYoKCdvG0Cjc0Y
w3YLE2J5HiGqYguCvUOjk1/81VFPI7T3Or61WwRCO5kLkZRFHie36njmR/bnIqSv3xsjyr5ehbwD
x28L7ML3ONPDc1GcxjSYiBm97x/8sAjGYHsVrbqBqz0yL7kE1NPMaGPyrSqilW2gBHLJUEf/+nNc
6ZmIhrjdS16pno+kChduKqgMZJj1FaRcWfvCrrFGsF44H6vU10n87dwYrTop1UcZoJFgzcJ1snMP
poJFPziWJlPnPEp6xlC5MGsNGCLv9KMH6BQcSKPBw1zFy28NnA+xN6zWeiQKrZ6bYl2XJlWXXC4/
/Aa2AoP+DfLcJzZwmCVxXqrii+RPKqDWmWRtRezPyo0ptx1jb8PDm/Mf0YPGtF2ChbRa1WlfagJf
+Kna3+CiWliuBxF0Cw/2+HC2JShFiaWIDsg0pBdh0ixrPoQqydLfd9ldi84ET6M7Z0yGJ1gpRKjU
ofACpXShqy0lx2MMUYDvCgTMLiVsq3Dt+FH5L8AZxUBEFb/QfD1cFe67P6AczCsZjxyXfxwK6F+i
MKPw6OFvpYi01UXKAnb0PIFlREvTZ9xIT0tq6TTPfNa9ivlyi+vbqJ/fvCmcujTGWH8CUn6r6e8J
fpxAWbYNcq98t2cOxuAOTVx9ETXLTXC8B6WU0GTNQoadnXPyWchbtjkqmQ17B8TKn6FyOpcuJmEE
xzMkLGFn71Ymh7CPG6goZkGmmVIj3fc3laWGXvrBgfjcPwBqsggll7jqQQjb81OiNVHO3m/Ozdi4
bbCti96M78jjZob6ogzpM5sb8e1OnZ6br/uVmxhRDMHb2cu59xrT3r3HMseJo2KHMP3TpEme1V+d
XdiW7pc0av9ee4A0VIQBHW91Rk6NfVL8ZtSGIKxn26jRDKN2e/F5RDHbvKMQAfxUjQrrzT61uKfz
LduGB5Lr1GEhj8bAHQrdp5drcnubGaEeoGBDmagEEC3LwEeg67+EVglohbZcSutPC+TcPJkr3eon
FTcQ7NjEG42CokqL7/Ux0FEitm3ulun7vBuO0DkZvQ1tdpuHkf1+9VQDv7Qf0fTcVFHcidu0vNwW
r+LZiOlIB9zrJxpJ4uc46vooDSaFc2xmw+DJOxIMnw76aiejbkd8gMp7yvqrWmxoo2wkdDgDLIEj
5oFlKKzoyyX+P6G8o3hl3IROp3Vox2dxTyxrTIGI5b2eE+zemWnA3tTg+bcwNWVRudZVwT9Ut1re
DuiebHuYqStu47rxPauMEQ+DoPPXiu2PvdDenS/J+aGGKBWwDLAFPr4ZkO/89oomSF3eMAJtZPnY
kulWzY68tBPvZzUryLeK53/J/YLD/UkKDPSMRveOpYrO1R9D5f5y6rFPdDifdomhsy9RopYXWyEM
6ASrlFk35N1kdmdb10nA/wP+aYh1Zh4Fu3ua2q2HkFNtSoiBGVbnuV5d1tOw0TNtuXFqv7xKz4rR
rdLmRy1yN0r3nw3GtWcjz4ccuoPaDVzsJWkc27i9/lRpnvUoeEnvNtQTkkijF3dif/3Aw5Ud6McF
nBzX7WhxayxiCF3wBwAFSSXJ0IXB/NJmro0awlo5nbealr8hiucW7VdIJg8HnSjKwQwCpLercRfI
U93bTBao2Thvg3QQ704wdqiNEg0T9O8IX7aX2xYWTjBNTSwURp9F7reReSi91FSeYz9XUnt/asri
XbgPG2+YCNc1SDBlq0PeTIX4ZPLgSEtxiUYiTDEsQeYihyKYpor7sLjHzQxAN1mTT/yAnfXUFyen
Ry0Qjxqfn9ccVbViqUYdi7sI1CQXPzWqOD02+yqd7RJS/Jz/53Okur9e4uLjg5pHiqDWfvtF2YU8
HSLkk2b8eo8diXo3hoy9abagXIJWG+0OhwLfGl+aQ8pnewHszvX9KmUpK/7BriqW4MxYmtrqlrSP
Y9yPjKbBB6wKnHVet92ACz3YcsnasgMmbYl5WC1tcNplzoQ6gunxfNWC3FBfEH4/MbpJrojuF4iY
bz0H3LcohhA0t2C8bpNwhBW/GF6KSKH/z7lTSOlz/FZiEzqkK17M2/3qMRB6rGVGVs048tvHPG53
JFJzOQHmUFu55ePPKSpwtPy7aGuPyKhBwWZ4Npzr3uftPDiPHGuezGlAG/vGLXNDipjRapDSSHlc
8gJCyqIpGx9iY+DN6qMy0Tm/zCEXty4c3Fe6/q9PhiUEnid5JDpT18AQ7dakfe7w/2vnxueD56OJ
KY5vQb8IGxXTrWt2kmxA9PFCVPLV7NOiXrCfzIVRVVPFWeH7k4kwMjHENWblc5qSw7lv0DwL2Eva
Lkxuhz9G0Tq6COZY7hxloAxehh7UHigSZ9DF/ipXL2j73LLP5LILRzD5OrGgD7PYptWUibEW1dR6
8L+L6QKJJaaHzSLPzCEEFq2ZJouOlItTsmQkh86J/M1DxnbAUPP3ofTHwE/0XNKa4e3dSk7MW7gb
lpHPza/AUEsNrs2qDKoiPf/+iQIpLu2IvPuqqRkkHjuhOzJ9Z6qxTrxdSWOxWkcjlp75M7iFZdAl
dsIVpe8nfIbKF/anWTvemfUZp59Fl2/kjVJLO7qpBX9Tno6elt5BJmdLUr984vb9CNoA/pLNdNlW
Hd/H6WproGJoK+D0uRJiJZvYLtlNA4/+l34qOum3aBHwnxslCsGVYLAOmiKuV3Se5tJGQ/26ZNsI
us/+bpnE7imKqYICw+3RiiW+3Pc6uR4pjc1o6gIxGUl9MyreNVBtMK9d9SIsRIoG9Qd4y8KHy849
DpQvUm3Krek4GHmdTEqJ33DNBL0yIszcwtYAJUig3wBg/DhlzJVZbKkGLS8hbnGwsKdN6Np2/5mn
p6JvkKeG+V6JDAiSk3ZEa0l+fmRBXiq9H4a9EUSgDIkk5sqcVvsB0awPeF6chOQBuc+eXpuvEyY4
wM6eNxLhPnIy0NuUcYRuXlE2eawJRl9LxkcqhrtQdhg7sup0WS/SJcx3hgSIS2HWOhqqOaN7wiNZ
8P+zhKfBwSTFiW29SDkGnR/bycUVIl4+48dhOXdZywh0LR3FEdL5FuO77qWNub0yjd6HNr9LsCUm
2EPq+TncX6AQUrs5M1Xlhny2maHC4lEGO3ZMadGyHmehoDYNf1s/3BvGyyNfD70H0yqTX/4Xpkr2
KG/BZ5slcfB6Bd2WBtI25kDwMrF3vJ3F5cGe+V+QOphE/A+wnKN3Lxbt5oXfyfVbMRjgKKVKaLPa
rVtyqhYVnmYKa63DGCepEkJxhvdBdFRE8t2uttbcbjLYT9+62quAm0GKGBJIUiINRRwCXPH65sS1
o5tIwFow2So/ZR6QPSW6bAvQH5HF2izGm/lBcRhy18Oeby4nzYNmo73elSlv0DoxQNFBK0XHNqwW
J4F9ojizao4wQjMFJkP+P+n3gJRHDPYcFswpFRKx0F+Zg/CO5m04fCaFM/pYoVWEUrKImygMQ6Mq
Urgx4A007Rftaph0rlVf/CaCOfugx4Idq2TP8gHAr3x77hq0NUfzbDnCovBZLOUHMq9QWuzy9a2y
B/JBiFSL9VqvPoAhrcPOnHR6xZia+LIZraESMIJD/LUHygIcdDBBO0d+gcRh2UKzlA6lC3ofZy26
RvR1oTpEiBEzxlSy8rHPdgFkucxi8HZgiZnpukm2fQBk+O+MrYGpsAN2Ygtaily8lzMFpTtM/ANJ
vflpHkdYozXSTd014JziNhw25QBgrpr1SBwugsHAKQxgbAQ3xipUMkT7krKrH4UpVgW9g4aJxyZq
Lw+Qg/iVOfLKAcRtqDkHB5s5RiPnjopNndTjN96yaKKUzI7Bk/jOq/T92SS1hUpiPhKPQQhUOoNn
t4TQSIlZH3MbqmSdz8+RDAHX7IrhbSJRh3GZGlLnUUeUq7tgLAzxyENLGbS6XnSGXunnudN4jQJ9
r7clLtGZVJQZ78GZBbQKIkI+RpptG3EAjd9aQ5PTW5WxiS+a+Ycjkl+2hy3JDLBbs4g1UAbDre6E
pwEIrcg97+oKA3LLpSE5DRhWBDI0Q9FVLTQkwQ4Xj5T8Z1faDaLjiVhpPeKxF5k43n+ziIFsoSX/
/ybutO7nhiLAaxUG1m2qSHCtxEHiG2VsPL539H8BM8hisQ1aR6e6gvBJzfrsjC5NwAvSMInpwAF5
j8zUuYb6pftnDw+Xz2BuUtURm2WbHywZHfUXCYGri6nsGICsTkven3+B7UcJyJQD8dMZgI/WXfpi
/qkq2e1kQAe3ZcMfsm0h/Nj8M7VXTWfMb8RcfX9bmqV6i9RQPwsKxej4b2lP1i53DCXwRGpJVZI8
L/UpDLy/N4LlWFXHBuIbWHTFyS1DTW+QgT0ijrCkMX4+SeQR3lqjRuCdDnTSUS7LBH0q1/XafNPn
CNIPGai3fBa+PMxK+wR8TCtpbh0K/tR4XV4Q5jMdDGcTtfWGKhLu1SquuAmDLV/o1YR2rj7AtyHf
RF/Zeq6olHhzkPNbaf72E8xEs7jqrTz7vSW7cZqj8oCQ7VlcK0phqbTE+I+9k7FjmLWTv+IUdYPc
R9XUlXLlqWSuDch6UsDTqhW63PYsOrPf3Rip8x7bxVf5usFZ6ZwtFiPEk+YDpRi+rUhL2pKPS8gb
3fRJhVOH7V3MiysStcyQx3zrnj/K431FmwGNBThyosyvPMVK4nLxp4D0F9Xd+BvOJyQyMe2iQKIr
jcFCN3Vn3qtckf+y0MxdqJdP7b6YYafLpS91k39+8YdtOTljQvJdEbPYYzvOeEpTFy6lH9VvVm5b
zbQ+f+Z1KXoqBkzQus5OwsKcSdc1IZs74AoVztrcvakuJRD9BOOdQbWaiyPNhVeEJlkQaH83g8k4
xdVXr1O/l1GTan8vKmw084x/lTChlHdlAdYy1VzY4ylu4yn8ODD/zi9Ns2Y1Kb5JDX8c6R3fyQQc
hqODSVrR+OfPqjEip7egYO1ObyT9vVTM4y6lZ6CLVWeQhBo44cM9pyOwAEk6v/9ejupfi3n02ocz
kdhmRbdxwAYfMuvvg7aIq74Cg4txROaoK0pJwZ2i96qAmRKWOCMeGintoceH5Rv92KFBw8yudIBS
CVFVBIBGoj1QbEGCbfpDKHttrD9Df4+AOB8D9w1qN8Bnp8ydBq+byuxAgP4FK6LCPTl14DeHqfOW
Se8CVnCI61CY4eClf3RZ8t2u/4fbfm/AhSaYOjuNg0kfH5DaDwYi4AVYtM28vIanlh77YwD4kZX4
wUZT0aT72Sv8PqfsajIXf6p13k//yWOUt5OMGHROdIsJS00NlYcbLfLRbypOiQzKubXQSAp7uetx
A7txFWQv/qTsXduTnDgn4rrjv7i85Mlv+Iby52JKhXe1sORtoaYrBaGcAunSTY5Y92G5PlgGYkMD
gQ/GiFZ2ROl2AdhFsnhZRsvIBJtgeRDoIMnoWt6cq0/oIUtfltYGkh/+2WLYG3o0XPtBckgi0mYB
NjmvpSk+GCwOXlCa+Smif5au2NEXSe7dowDW3LCwrtvVJNgL0qnqHyc40VRRiudZ5Sfins5lVdUc
hmV9s9kmX2e8csnd4/SuuKVa1rHK5BYl9rXxqL8EKUsX3I4mwsF6tf3XDgNlFPgnrYz5DxcHTmKX
YevtjBJtE5L4G/tm1ObL4GsWtk5GMIY8bsMxGMUSDTYX3edKeGMhxHK/9qkFFD4MSohtHkfQzWmN
4o24rrFPMMRginy6jLhJhexEvCkrJEvZPxMxyfoHRQLessfpFJCpBfKhJxdmU4W87uH45f98AMQM
Ty6QjMMYTV2mshZEk2bsSZ3OHCgDthL79DSVJj4fqOoeflyNHOwZjVXtGHwUzTYgTHgSr+U5U+oo
DUa46T6D5zf0JE5bOVDBgiQNJOlw+Lhrr++RdPBldji+ACn04ix8nXUl/PjbOt72f+3cocFRdhsl
o8Hmo49UnYC/xGWUpB/t/J9gArBjxwiTeZBATJhwQsVRVlHb8hKWntrPj5D+XP/d+P32T7z+AZ3f
zAyMfjO+H6MawTfdCriCnKRgMF+3YyYKPmfBsQUD405bWORlQeln9vW++dd8Ahmbr390OrY8IZCb
o+JZPhUXBovqtoLr0kQsw+T++uUYqLEeeqLATSyuCmpCAGqlMnYo3kpchRW1cS+JprfZd5CXPImm
CKuUij+i1zV+YF58e6ax5++z/CEqMTPMYm4NsXrXtVsRgyMB41MbBdra0kMFsvqUKP82xjNNr6a0
eidTuL1Yrvl38K+jbKUwGc+BOnrBGpK4YvzHz0bB/4n8+96BHY1kYeaZ7Xvs5c5Of0gz48lYNAbd
183nPY8eTJumuUAzsBrxc+tR5x5+4FerO4c1jrcrk65GKTFpBDyn5YjqNMRXhvWQv5MavX8mf5jY
51iKJwfH1FZFOSwgyq82nj/slZbJNv07InJJIL1ADZNBrgF6l1xUEG/9geb6I8QfDIK4RRPxqU8W
5TjDY3xM7prLmfdkZld5Up9Z6p/LCSpjuMYA/oQVXIhivKnzAkTa6ha6gf8wkxkSkAJVP/t/BYWi
JWnD3y9gsJvJ+GqBepyapmOrb60nWp8rO5/I4Z+qZfoZb0LZerg9XasQ8rQk17M2s28Z4yV8/pl3
1jeEpwOhU6Bhg2xuM9VBD4+QgEw0MiDExho+hC54c9o1qOYi7xcnszo+S8V3gIU/8CxkQxxfvEl1
s4o6tqr3McWp6wFW74yrG+Y0QXlyJatpd229WWen3VLUsQptnK2QPiw/H3T0YTPEMZ6nnxQs5mkG
GQCRBHG/xfjm3Wb8pwnIpwUS54raWe7WLysp9bSDTG5stnntAbF4lzr95PvIfyU7ZKAEQNVP6e4t
qvI5wGkBuJjdX2jMqNYMeAn7cDNCy4QSjA6+VcKpf1YU8AdpE2uw7aWi731MwDUEm5scqXDrk3TU
TRe3HoBxbYGiFTCuRR+/eOmdUHXdMGJkMoa5rH2efMQeAM3JSJsnMYg/6ivTa04Fbwn67jnTAIuE
W13ZN5pQ88kSCL//lvysqry3/8em5defuNRemfImkABT3tQdPGHdMhRhxEzA+2H3fp3Krepe1WtF
cLedMDsJv1t+8GHuh5xcS7td89Dr0q/FWa3i+Q+vn+X0DtQ0fOxl4N+WsmUMKsV3gqM9UJhF94ba
t7WCObQlwwNhx5yj/6CWC+qjZ7zRReqDu86lKkBw615hH+OoPF1PVFDPxed3gHX7obsBdtFK7EdZ
LPh/b9cDhjuryskpgeoapjeyXAQMkErmXfg9TJoWLwsl14UeTMbTLjbAkWUpV0olShR4/ziZGKwg
fBW5wiGv9eGL7DwGk1728f78XFxzMbt66ji20zUw3bWyPbq6pPQZceT6fGo3gcVel0owpguK2J8m
ItSSRhF9baNKaK4ADRB8BlfiPsCduY5BRdcPk6THcXaYzQcNJxmrUmGazAjvGT6GXq2roPqN1Wxn
VotdcSaj8VrZYg+IHe3zugXB+Euk1JtJTcQF9FT4YT+e3ljRdSc2+ljf6nAdXpwMi9s8r7Zg16yS
+LY2T+x7uLTfexNJpQPBbAkbYHh2MwrfGbsj6iKQmSvx24nwhcvsp5+SlE5PnUBq1IudnrSQ4HwU
mCYH16k7EsUpyoWYfC9oO+Dt4Eogh4TfgQnPw5M+mKaS7VYwH1cEX66Sn7hY3MvQ9OSln95cCOyO
SJypcwnTrF44/IzT5zoe0WtWLs6KD6mSiBlO6b6PYYVmM+/SLYsuBpthQNpC/7cku6H2aeQQqvXs
u5RRybFaliizOUhtyc7PaSBkarQlRRqdXXjSqm2EuOy1UP9zlwnWYDlabfoTO+UHOoXlM+PZ6FB9
L2A41NYhS1YpGhFwf6YAxz10cOQWepOMcJShxnn37kH6XbX74VLDmsxx2JIYflr+SXAiPEmo90Z5
pbIN+AKeC/3wEj5m1MUCRSBzMPG84sVSVq0NDf0ljax0IkZNjOT8PKur9FSp3LleRrGLaPef5/mP
bqjO7LkihCTNDJIBWnNhnmgXFAGRg+6V5X75cLxIm99rz4+e6ld6dBURw3lJGimXgpYudDN2PaPJ
8g3HcIsk4asdm/jA27MhtCUOwGbu+5QsE2+FB/r5LcL+vaOMqVuAt6x1BuGm/DoF0ONdD6Bx1xGU
7i+Rlce1t3mz0wfKi7OZIYahSZKOHe45PPx/SX+o8xCvevFK17/BLj7aEK4U29zA8hmXtrVVg4HP
QLvIEnd+s6Gtfspal3i2T68vIWTk/iPNS+oSUT6FTsK69N+GwQ3QEIADPUJifrIQkurjn08ShjsK
4xJUhbl+p9aUFJkpjZivEKdCpHJkToZV5lNzM46KpEzg1uEykzdhT/DaP5QysdClLDHv8Dc/gvd3
vO5vMQ1A795LGUmxt0W6S7nj/60eziPO2Iwkzlr1jtuIumWCB1ZMLxBUTxmGx2qeqcoPmmkIoHC0
hSAHn3hDJmgBGkUVUfseIakWjhKztkJywxiSaNKFkkypleetqwIHHZB7chrrChr+0QzK/Ct08QOh
sQgqYBBl9D/qpiHCagzx4L8P4Rjpiv448773LcquI6XNVNVe7eQRYNut4SCYl05DgvgiSrn/AWAH
/mURn8aKEZ6MGOFFd+6YekVTtJVP1Nvfxs0fs994dPq3w5VQ2WjyGf8MrJhYHkbVRC803aUE08L3
FlqTmLgYi2jifdrbok9WROpwTc4KNgWyiSoMZ0eo5cSsftuPdKGF8+YzpS9bubadzk+Kc9QNlB67
RTcBUP+Z68s4n0ffo4bFgOKJAmwXDAGNLuzO5fT+b7RGaCrNq52MFN7lWDYdUBIfxU4lKKCT5fyC
7sJD9ZvtprSOjw7SBVK+sPipKha4PlESS+MgrYMMBbt2uGMhO6GY2muGZ4V2nUOW/Z+ICaJt2mXs
HHjvpRFS56HnvH6EfTVbj8NDCyLlP5rCMzpGnPNBKRrd4EyRcmHepaTkEvqa+Jm0sKYkNUgVAWg3
FG9QGsT2RknZdagQY8g4Jm1OxhGI8Mk+3HQf3Hh25l7EV259ZyI862e7w6Ym+rW8dnA2fqpLsJ8n
P83gxjcxWRzC93tbRPRvKABEA1LD6YVaVRVlehSU57ur3SjNEbZ/19ykWRdmYIxfxbCOSz26ZVNv
PRom23qxs5YpySgpNqboh9C3R711wPddwaBjoxOxIAEkCn1X340efNeMuFAbyUcNAlgeHuSLx0jB
jmcwZQrbzpzdCFGI2s9HJGVUiVoX67loWp4bW3cnexWkv+uWWZelRlFdwSHiJ8cyPPrwcBlgGwEa
rDXv4G8mvvnzkVOviOUlroT3vizxCH+Jen3BTzyseDfKJoa1fQaZ/0L4SaCtDxjq1FICOnV/ON/j
yd80ykxap8CtbT8yySb+8Z39h4OT2n4boD2rabvQ4g/DmgO1QUB/MS8JqarntWeuDiRQtQMeH99m
vBIAIyg5s7XDozaQkKTXW5TNxqn2LQ3JhLX5j6ZCt7QCdX0VyuCcWw9jMw18BHWJzWvRs0j0axuw
sapu1ZHcvs1oNUQeGn8Ot8ttmORfmKhfxTMswDRtNUztuFsWB77ReK4QaBkAB4drj6NpAlUUdFER
tor6GzoeA91fbbJYyNuMLLas0BJlMF5O5bycQ40xtvT0bxmlJRFaSIMfC66HodMh5/yQFXRbapVR
kA4ABkc/9WQEQ42k/dcY9HE+4pFCrqe5K2nHBZLdTfGqtL6S/bosybw1CwBuHVEov8S6IZLkuCOV
zeEs5k3J/jX76rXny2q5wvmR1Ptp4OgUjXgXXYgEBtznLH0QajqX7yox0yxoADIB2L7RHwA0z1Zh
/SeDatfe4JNoAFy7hTns+CxMAV+6r9q6uQ0MDgXGkjegLxq6qEVshAGcRTQnCGCmrblfEt7LIS0U
0fH0tuLLqA+UgVikf4G+xHwnkMlblPioJ+ypEojXFg/fx5hjWRfRU2MjPP7skOtMfX5zybv+hdHB
nw2NlcE4fi0vx1N5ARwbsdV6i4LQ8BkxXOzwi6RXdMe//lmnuMrMf8drTlFpV8MJLZQEuMp6tQq5
RHVScsrY+h64bOR/Nli1tiNGcVah1Rpz6fYZqmknNQvmPfEyKyY4K7FIK1h4tl4SqhBrGMygGtEY
KbISAXbpdadZyAiSloF4wVhD9xOebvhartiCksFw/PbQmnzJo4bp7Tm5Gljqkr7hNqW6Bu2RMvhq
wTBjClAQdrLR4pdYDsdDo8hMz9SAL18T+xwiTi4wm7dYgMyXyyDRR0pspDuiUqKN8hXdTotMTPN+
Z7tapr8+QAQtan2GNVGHM2MkDuFwSMKH2dx8Fr1dLbGL03YZoHhmd5dlCInfNk1TO0wKkrZ3AHKo
6DpW68vh+i+VpH6tUjgatXMMLVCGhtYTmVr6vH5xHm0jivJm/BF1BggflEHPiI07+wXSSG9MdYBQ
xFkQTv/o/5NRt17ONwcoel8air5KZ+fMUSekubq1NGYaWSqfmygrvgF4txeU/uQrtUR3Erje5TVF
5r2WI5J67xEH5d/KyNWrwa45eHOA3NqxclnzBOsrKVK9nYsIye3Mf5sifzkEJdfHvh2NGr3gC02x
LUC7QQLDm4hjPrM2DG0aXJsvfaBzqZ+2yYOVbB5dy9kvtu9HJ7gE7Sv8TgshS+B13w2s0aoMS0BC
mirodQJx748mBJiRj9FHPV/Y+UovK27RNE0olaqW2OvqyYBoX9oz6cQZ9Ech13dlDn+w/nihk071
p3mYbj60hTUE+BU+OWUNTUuwNB/wJDYq3//blmw2rydZhHPHukD31ZLAOFvOjwfjeUzN2zbydecQ
4/J0O5RFROUB+fDthcz6g/eHlEgfJz34d/EOKfOfmgzT0HCzBA80q65o/Fx1LAxz1LeGz5IWwv4i
0CevNwTqqQ07s/0kfvPzJ0OeNcOyCs0YYcOzg7Nv/RS94MBoyuTmZbjt815+WLYwKrWl6QCasAgc
/6SnpOCPCiwCVYKcWOCWW50IQrnbdKKr62Drio65F/kKZHjajr0cyzLgo2q1yLEFovj1ElFLfEY8
N300nhTCRD8CI8wZwkyrdzRfUR5CoBMhI8AxzfE4NGRXQffI31xyYdxSO1TItxCtdjAjkgY0C4qw
Sqg0rfOzU7V0x53eoo3oE7Fg0+Jzn4V5OCl/vmry21+e0YCHFDp8Pod6NobJqojPb59yBClEuwQC
BoP2lnsa9jaO3Z+Xmc8/i+nlR/4ZE5dFQC85N50qT8mHk2veS94r7osIluAQOkrcO+8MGBi4Tfpw
J6vX8T1usUc+9vX92Jp5tYZCBm8CwSnq6jidDHpjGF99GVmDizeP6eOHUzrK1bnLliIIbjMAKLOo
gaRkqMKVTSoAA7557FIOkeEHV5C+GFp1R2rTkiyM+mwL4npDiYErdJAcWB/UgCcIxFK8XwNuG0tG
GbMFYyLkTx9Bl5MH1BTJyeMIa/VgLLeOzQ7eoOL8PKVlS6vX7M8aY+dDcR0x95QswP8HGb70vK4t
2dUapJ9vh8106HJth2oHG+9yhtr0A/joE6GUOGNebMOyUInOzeLop8WBR4xpz/BdSyy+tX909nKk
bnXn5zLZ+BxAiLe/DrjJG2ixpUN1/kDMmncYxHsFtxbwh03vkN1wp999imlk1kdgm2iEx22GmaXC
c0OrpTHENH496OQSDuCYwoGLy7SqMEI4GS4z/8OEsDBux1ERCK55KDsnL3ptHz1SCRTsFGh0jUrB
EfyzlaKY6lLRB4wZND5fo3d7Mb+ItqyTsOepBBbshSD2yFLauTGwbvGQeLPU8Qbb5Et4Gn7TvHS5
sowEaEZyqkFrXFYWFvgeNXAqmhWo5pytDI8wKX9hQHdI2CWlhh4OIiGTswkJrNNkU5dG0Cn3ao4f
erOHfZ1xkdzwdy2AaOtp0B9rc7ZdrOnxY/MzlEcc7RQuyJtoEOj0WIkRMqnwVNnfE8TckP4ZMMNN
NbdMmcacsE1YkFRV/6NB6KqiVESslj6FBbvFqJZpwnwX3ywOBYNHcWH9HXHxOE2DJbobR8HvpKLe
PqZ/Lw3rjFEQrikjSrjJyUPgKUXBK6wTN05BKhTkNfzYPaO4Qg+TW4oaRWBwXbQoUlczwtsyksfk
5FgQXnTS7dW+WMqjILF+9Pcb+XB9rQVOI4ObcY3vuP1J0Yj56U/sn2tiMDZMwD6b8Of06yDH1YPf
UJDyL40UdhrJAqoLtI1Cnb0/nlLVj06n7cXDYhLrlNPG7c6efeV8IoUpn76B5SXMBXEFchWSFksg
3LolEAi9c91auZH0RQ4k8aHVrsuiWQGhxcQ8lpK6IkeHSYIeyIObZKrciuXVQN5GWu81em6p4p25
VxDBFeUXMsg9tsdpAeTNPWzdI+4dAEkAN3IAmTpO9Yuv6gpf6ckKLuPvVNQ2g73ufln9LHxPq4H+
K0+5xKWHfoaP4QLqhEOI9ErPp/ZwJxa/LIktaDUnx4XqfEKlKoCqHH8+OgMLNLUiy/75rZDy7qBx
EdLDHyDBsj1Vtuf9Q5TsO7TL7bk9kTIPwadmibiqGIr2YTKWF4ZOgbNZJobppCE31hpo+dEPS41V
4PUs9m3LYX9BUjDlmR11qvNZ8UNvM1M3glXCxlQX0NQEZv4tbKYzd9U5Ku/2TUAR2qTlz2mLjjjT
R+XxUfTkGnMQ0swfxP2FllGi3EinXTy+jhAnSVbPXLOiVnwccJTl098mf416yYPIxwGg4x6L0uU3
NZ2tXjZu1RNsCV0T7JC9RIVyKSdJsVloaYuG3RNCMDrMd3U+YB78q/A0oeSvdvoPC0SScBitVsAT
m+B7gELlodCtNlLQg2SDzCvmYbFPFz3Mjv3VNiK7OYcMyijtUQ6o4S5qgRVVkWvKz8Um00no70x9
v4OAH3GI3L3TJKO0+3B7bGtOx0NCP1H3o3Zilt6EK51+5rYtH1WXoHJftgiiDgt3acPW4BKnKZP4
o0iduEum+Bv84JxLJZgBworNidBUiVRDgGh0j4xn57rMkqNbCCBqJ3OlB8fW/5ye2ecsnMdad95X
hkaoxrsgbWBiTbQcQYFAq2tCVFTTFbf6k2jTjCRQw6rkn1OVsqY6XRAaC1QBJgR/fFXR8jnf9Kj9
1itxyIJ9atUgz2ltkb2f+AXSMJPgnuuGpOKm6j9Js36yL5bEb73wlKi3Rs9f3c2zGHxqggGgsOi0
34Nh/OFd8TW9C54TI6EDDgAvw2C+5IV92CWjDl5D9JNVOXPTnhA0VAbNFwb2xcwUYZEtmTicj2qq
3Aa+C67w6vk+twpGu+dmt+l9pCoMAirTJPZjIjXY7HxmzSxM+aja1A27pAH6JZWLh+j/1tsEUX9H
uHBjSmcc5efKFGR3aE9yViqvo6NbiAGeCFaaMr02Kah4Bk/eV2M0Wr1mO5znJ20CfFrTbRfV/K8P
Pf4Q2WpNME15Neqv+g7MZCCaeoRsc+0Ida6QC8R07XWrz2+d30FG7r6nfRBKvqsohBPoQabGvqBz
wYT6ru1PatfppX7ZHBWyNBU5fUzZ4OTD4OZ85+kKpJ0dObQI+r4j2T3FFzmLZj9kMUOPi93NMkQ2
i4mmbeIwGFM/OvOlADZe87p0u2FqCo4I5M935dXlPbok3yE4iPlc68G56NNXnA1SwU7LrgGEqApl
bzTWi9AUHZfqrxXq3OS5AUmuTEcDtlsnAkF4g3X+T/80i+0JPE15EWdGaoro7mBp8e1W2n5F5XaZ
SYiAM9DkCGnKY90lvSHKPDYG0osWYMS7QbfurJiAoxPv4vj0dVDy86TX5wzib1Y14+dAE4h610wN
DgdrwDhdTlKFw5SJSxpZnIFO4+pe3MPgyNYvZmtZRltr/FMFt3mgYy8T1C2d1Zv083vJ6+FxTCHc
L8mRSmnkSi56WQWj3LJiFLxQVWfOiPkbTb0WmxhHzCsGwSRx69AcEVK3DJGD8IRcq3z8ZIfQ7X1A
udPvR7bSSzj5zgR8d9xGBJgeZMc8IbmxMLMOD9tyCVKV8/9HrWzgigyGksG+PjeN/v18umAOgrV2
yMq5UWyHH0qcI1FxHSpjQT/zPOWg2gLnA0DHwnEc2rBtc1IpODfItNA09kOUpbS6wUDhFeAVEbeW
A9djm7bvnfc0/iTO5BK6VBaCnHnEM1eGOU/vt9stbPDPckBUxrqDpwIkiIVH7KU4zg+t7g9bwnKz
eb4j+OfW+tC+KeJJvBwumv3PBTRA/Ak7xhXlubg9n1+pwWvGIuQz5hAdo4Iou79YUNNGTLrFbKFc
w/X19saP4MFH3fhrUMzYFdiFyU50pyhoJbCePY44VNd5bif3yHwpEJvtfoZpNy9iKrVCdQKIFrFy
pHi3ffEgtKA3tpYk9icIHpGv3l+ub0Ivc9NlyfN1ERNJlKlXmGiHsUHRJp9GG3JecbD/zLobAsEb
eBHeBywxoAcw7xeq4mu0OVedtqr0q3FWaIloKGBZOiaQ6S+L2oiF3LyjIynunBOqOeCHxJ4Azzpm
A6sViPtbVXL/l8EsIr336i/dtnec2isWMINwHeEk2gKoCDxQfryxydYjYfiwTT6oX6WjfvllWJBR
eN57I6qkk8iUI9hSpvflQ2Al+0ViOae0+A3dCtNmTvxDzGGFdnVM95iqnZ/5m+7op/y5kvjGarFq
fG/BXIKpTKZwtXKTI5lMd2EjOnRM80gu/dGBJjzGDMTEZt0iBt8jwff9ovGi9MbadsUETVfEVo74
p1vh/tPdhb8PFAo+x1JiSSeiWEs2cb3BzeUBcHzi09I0J1mTkBzTdTSuAnjyj1zLoP1wWTmTuB1L
GpnqlZod6eStPfsKYIuL6u0bspy8N91Pbf8jrjfsJu35Spmmss1ocrq7cjmHs3fExSVd4PmF8Oaw
qWtcIeWPJ7TTypfISAkkvYOCuwaOMsNEJG2PCMflsIYABrn77ebI8ETsu4lM4q8UThshaLms5dy6
1kBkK0FRa6mFv1uAwU6ijG2BJME753Xjuxhe3+zpvXJ6tlujKTd1Ynp8GuTYzgRO1PfJ3vYvLxXd
p6E4tJBptQoQyqs+rwU0u+8bnwQTK7vIOJGeXvk77EYu2yhsoWnNsT6wlOsUDb75qpJI3j54thd2
8bT5FQElJOQJXiIFKu1Sne0/ubh8horJg20ZGUqH9XXdQewkwdX7WqYmsJme76R9vZxcRvg2SR1j
eGkulOMzyJEW/4i7a08mS/y3e4MprWwhbwron4IpN2+MzV54Xinsj3Gi4dWN6tzSNLCvUbHhgI6/
YglGHtRdvPtyXUwzdN+Nh5djmGmOTCRPuXRiZpy1D00u59vXJPv7P7v/iQv1L13YYmzFUl8toPJn
gamgv46WoYp/gUoR57rDx/wcqu1RnXDemJi555Ke+HWWcbdFTCsMdCDgf/SRBBTRJeSB5isYRqmh
qf+LW02tYNT33z16Gj96b+DixRnFaDBEDxWeMFOYcxSYrlUrXXRWPjdkh+6b3pUG9lllVO7jJe39
oFDKpNioLcoBr7vCi0TnaaNlVxWfbNCNmr4loljYgOu4vphKEzhvC7wVOF1sOz9LsnmZVDBku0TD
AEAFzui5YA7M9GMD/l2QkluojGlZMqTsjjiXp6eYhjQ1CT4cewlHDf4MIh/ePhYIbAAyl9z8+T/o
7mpq1J4CsJM0m60i8y2GjpraJF+DcONWeOn1VTFfkCSwaHFza/iElKv2gR4Hfjn2PFCYTTZzxMwf
1Khcr4nj+KbuZkFqJmCZYgFSfg0GEJ9PBQqMxY17VwxO+F14Zy/3Z4MxqWz8WFo+gXB5p34j9N7d
d2ZE1q3vCqjm9YyIt0Ot0Zs0auwc1Lde22f+bKt8ZtVHsa3oxdGoPP+euQYEDERq34d8+jQneGgG
7V7uw/Gt7a5U4pgLcZUVVnJFF7Ab9NVH/q4rPxb4WupEtyH4kped8AVvb7CO4Abh6KQaG+hXboWk
DAQpK/v1Zf641SoNLN9pUVspM+U+ILcSGumPfUsXkfobo+g6lZ24WOV1J3ls/I4Xs1j64B3+oOmf
WvNQIbdI94MDIPcp7stlJGUZd6K8L/N0fLao7Ia4rxBTfuXvKtJhlSGMPsPNppbeefZDa5xIjx2E
AdsLSZz9C1UfP1uGACg0s1Ka/qmr42SuEH9O9ojLN69/tNBg4R/txYa9tKTZb6AXbK8c7Y9HujPz
ManO3dEydVL0/Fr3mRzttVUj5hNXbapeqxlKWyNYRNPhqp53XdD8lIkwpL9tAa6EkZjfaTtbQHSI
Pxn44HVdZPq+P4nagakOCwXKZRhlbA2F/C4QGKXn45Bqyhz1BHh7lUpXQydYm9IKDxP6kmd3s5/I
InESvc+7PYf5Ft1Og/jk7W1slJvA78wZaLxixdRDJj6DVjkZyvnUPdFs8xyuSuKneCpwj+Wi2fmj
Ytsf9u1bTclyIp89OP4sqGqoW9rVuoMPk2BSw05tJhVuLoChv3chrxMIqvZ9RIiN7USO0Ij/OIBE
0YHQfNW+HNQodZTMq7P7fggFZiAPr6Bvqnh+i8BvTjtEbAFUQ43kYSuRHCLv9VwfI06Zj/K50j5b
rjDOOqfVIcTCI9OaPqsqnIDSyptJsanuaJDwD6IQqacf/2dXFuNgkCXfx6M3B7GIF4mkdVMwLjFY
hUI4U4vVR2tyR+6NFlCpgsqUGTt906y3sHVCOaBkPb3NBIH5gFSIIR0fj648s++mX37/OUYMk6CJ
frM9IyqCDTZggd4mq7hx+s39HgAnq14PpgbUAqlQxZ4azE70eE+f/mf0satXEjDDsPZcTBIH1rD9
5XTu7K9IfZ5EdJTgsLBPE5k638w2VLGPsmh0eWd5nMC7PYhVKOzzppULiCJpxvl6vK3N/pM8fRUs
/kP75qZ4a7WUJQvFapsuTD9j2afE8MzKB0G+hUjAJHQKGESXBFOiEkbQjrNKMSvyYmjBjMH9ldEI
cBxi2gv6fb9ppkEF6JJqJcJzajjyoF0FDnSZClPsDWIz77SoQuxymtUOdYZ5TttQ0C52TEYq/mcq
7T4sOMhP2f7EhZssRP03VhV589ukOOcJrG5kaIlztppcs8Glj5iC4U/5FOb+9BVEN2yPazjqfXRU
hZd3Ut10Kyj3Y4tbmGYL0yVggd6R3z4BqIGZJB4HjDouS9r5jcp/8N8zc/Z0pe9P/EmXhf5Fov5g
jZ9gmAQexU6031ufBU1hy8oqGodsJTew8VRnSTVqvEdSt22hoe9LVjPyHxv+O45B6dng/x7syt5O
D0Oww2VXB3H/YYasCDbtATHvANWiVsDJ8ksOFK5F9cOdrCdENlrqYa1jypIthaepsURU244zA45i
fNwb8QRiQjKSOHktUCeS5rvo76zZ88suJ2rL3sBdtVcwX9y5aujnGBpkRl4Iyu+dkBqCDaqIbsEa
AS3GB/hT0o3bYZLYaR7krHtJSyCAbxKttmYMJH3GaOermEuXyz08WSZuZophIDLrIMZtkOjGEoyC
RuTWR3deTctU1X5BBRvGNk0ueCLV0uCDxBJQnrw405/g3vkyhhXkBQ3TlkGclFYsfO23XqOOxAR5
fqj7tBUjqowkR/63wQJ1e4bTF4cEPUakCKahis2VtGNS1INIo5OZKYEMqJ6TrUX1KAYjtxOGQVc3
3lGnN2vZmT2Z2PRslaolPQsSePELPrDKmiJvk6fF8iItdU6CSI31E2guGhO8bcDIcOH/YFvQMnDv
Gqo7lwneGnBSCqFDMzHSz+aLBSnH4OD7G5uInS1iREEzgvscpRAtMdoKggnv5j5n9moXCWfuV9JV
dO4s1N05rHdhArZ2thANFcxJWnCNVE3HG65tJfHhTXkFP2AeeXJGAcHBE+mWPENxrDbPMNb4HqLs
WV2tjeiWMC5IlXrkj4i/9KAJdXrs42+MS1mkGsMPIR8Q2GJfliU0wywrdjlmLd3K5RuUfBWJmxTX
G1zvl1oFkFL0jBwHKXun+92sUkuCk1fpDSlUIC3HZ/4yc+FTDdhE0jc0BIP0gUY5bCv/ZbSS9mCQ
KfZlHvyBb6Go0celXvInBIkADPX/BEjCoP5peKVIQS71yDxTdzidbzIkOiooKFM5oXJFr6ci3maq
JZ2LVb1Hxd82SHifpBj5D+PDZ5N8UxM+Hh3GzsvRALlvMiMMZ00K0Ysd1xi6o5pT9AlWnKOF+eEW
z6GpAzFg3BMx6PLZpVgDnvk26xcx31gPI2q1ylA5BX3+zaYVaMFiDoxGYVpVIRMtnxrI2tynQo08
/OUa47XCGVJGqwEKmfMI9G9qasponO93iumnxIU2BakXBn92bOssmkDfrOKUWg1kzjUsI8j+RYFD
Glfdycy97YQh0r1D53SlpW2ST1kw6NzFMM4EnA9YehZWijqjWCfLofcSFlpJY2M4+DMwbFQSBkAJ
vHqfmxTEm2DVNdBFfPwdXGB9Md6+1+uMcz2J02lpjQc7F5IkfpEL2cRkN+65i9X3U9bJNqD0bq55
liVTZ35GGrdI7bW2bbdfcNoqLcJ+FUzF29D5NlAfurF+CMhf5uvkidn7vYXZnculqvZOAgMqw2/e
FOQaQX/dhlfYGXuXwnpsHh6UN09um4uPriYK43Qh/tETzLvzoD4bDjksPE1380EnoqrXHUsfzlN1
eeSe6/oORCGfrBFyt6uo35HUsWrtbcYX7p/WQoRFgmXi1bA/vFnGtmNG3fN1RlAUTV61pGsLh6vj
cwVNbkYkuslzKUvPABiMWuSOxE76bhu/Pi57wTULbZ6qemR3bcIGWrgLLHwi3cEz+oyNtSGB6Lu2
Vx7X12a33csNrzBys1SS5DeTQT14N2hJyxnrFoOynY0JpV7Y/H4iOsZu1KuFytDmdcgkM3jxi36Q
7qfmSf7qAVBLEZRBlmliPosUBkpwyCH8IvwM+0zt4uD5SN4iKBUS5CPwFI5hWhgldVKsdDdEPkjv
RVEy6aDsOLAQXWTthPtcYeuQJhbjAk0S7wkmFFHt/fbMegG+DMB/EVBGeMi1wjOk6a8gIcA+B6g0
1XAcS2QCMYe5lCnz79vW4nr/EgqbpbW/OXOIDuJGUnomk4sKrgXrZBqZ6rCxaZcIRngNHtCNpb9q
hOskWUI/qVuKcEhiVULnbpz5D4+z95IJr9LZuJe0RA2TLE+X8PNgh4991E1SKVrXEZxgdWqMK7RX
7hSgj3Y749/6oGk8s6GA/iwjSC+4WWkO8+QNAw7+fhi96k5hhTk5MeObajOm3Q0yc5fbRilMVZ3R
GquCwCiJJpnZByUfyxNTGSrY2Er4ReTj6vAZyXhysuGZvuvdwOjY+eAIUvqOoI8OZ0tfvzVfk1/p
uhHTiiwR4RUkCJQwGawXzCOxOaNbcmEx6C0Vy00nUfIX51NfCwaeBGf96tnzBMyMDJReAzUoG64C
IpfId8Go2A0dr9g2zS3mghTZ6Ie5kGgCIqyqj34/1y3m/faEgSCEDYWO+YrXJBRGrGn+cBqJvizL
/LKDRO60NmwZnLXnskKjziDXv/EsinCCbE9wsc+94S3JMQchlCQkhSAiaolnI5OlHuYv7qx//dTm
pamLLqCAQ001E6uo55iyKMjdci70lGgemqagIyqS+hzU3zabDI2feSZYAN5ojc+l1CTpf4BhiXde
QW5N2Rv5y0ozb7fcF/dt4oLcLt68F36yYZC0VqrAxFrXlVyRp6vHYf5ogYTF6Du92OXzOBPBQX0w
bwteWJ5zyBFPTqZoxt10otM4lvMqm8pjxA7kJG2Kz3d1t6TaNlDP21WGwTO6ktUoWhiRSUp1o/dM
81E/dYXrORzZFP0WUec3V7cBsyPZyrbYBVc+yWk+K2KfZQCWW6tt5WY4ZbCJbAzwemux62eUmf+T
Eirg+UROFS59SWh0nQDIRdYXUtq2iS1Qqg4sHPkG/LxtHURePsBYI1Z62u9d1pjxiYgwLy0vxFPv
IIQI1d/Wm8Xl9xpXbk2+FtmxNI+DgXhPKMnEsZpE8kHcCMHLImzJaYWamhwL9tTDMlL3Wq3C8qAV
KACMgpFMPePIBaVJWxsFakAo84b7BswTCxPW5S3tuxbZTx255BKrj+V5c0z/R+j6UhJF7St87p5u
y731VP+tQBM4GXG0vW5wDrQwymF2HKBp03y7VSOXZBOVvJg/+s8T5i7W0V+Fs0mUuqQ9lqOXMLvJ
HuRugE8GhhSNCU5JVaYUqEIH0VuZjLQ0M6R65lWvM7FJG9yh7lvza6Ov9BrNhxUdgk+m0bsNjtzk
tTPAmAfB/o5ZLEEtuF7q6lEmLqV3jf1AWrKF4gijFeLq7PUTM3skWjDHoOb7+G76zLwdnKSasLXt
F6vE/PEhh5ULxSGM2z9iahvjMfDaaQA/4UxxzjEUd7nM2t9FH94JUdudpiSQm614sIog8jkbRWQm
9fBtf+BHuJmRuhzurTXi5Zr7XdxHPKkg+ANSfS/3ZjkSVdJ6aC6x74DW0rzC5Sx3ikE89GhyIIA2
bxvZwNnSZlO5fMg7ae3GTHKNrobW9g4Q6Mb4ALoMV3CdZZpecVZ+3qhzNRJQi/Yw+HzctlHKFDWX
YmxhmGgKP2/jCfn4lU9/5Z48RdRVpdSZwuUrXLFTwAdLVaoGbG1LnuZrkLd35HmeZZw3N7TXyRzD
lU2NISBm7ISZN8h7LmKY0jJPPnqlw693to+EQU2GQw4vbsVuKl2AreV6L1mJOw1vf2HC5mf/BsnS
MX0m+sv/1cXs8InIWKEsUKqJUYoNeTIFHRjmOSuhTaKH97vAfVLSsjC9uIkmeaQq2jdUpSSy+vIJ
qahRA1twQMH5s6rcyRt62RUwmYS372WesIgpLCJDS9Txt0bBzK2cmC/xbVA8D9YANKQfFxg3HOcq
Ll6eqbyM54WdxxQBN0b/sryV2eJyhoxoqX/CW/oyANSgWa9JlQeYH+oaiVMkQoWit/o70NSNYQoP
N0B/5LVMtfUygod4SdkyfhKqs54tB8SO1C03c9c3dyoHL7mYS4cHiIuDvCuak/dGBLSIQ5SVao4D
npGf6QBPEvnblY25JJZPnyj0tTd6ognaO1x5tzSVfBmNNDIAk7twNjbvur2y1jl+NQncScrEghH4
ElxmOtZAy1kLgFabiCC3iowLLaJV0jjeqceDuMFz2y21RsXdHhNhLsR8XaFLIH5yzUYvA/Fc52RU
6VWiR74nyE3/goCpNcYwnmjMQ3xcfCnQlJqzOmNF5kPgeIUjLzQyyg/l/u7AU0BIQrn2poB7/BlL
if1er2h7uAwUmCDkd/JaszzNDmZuYnoTlp1ullujjdK3Qdl+BFDWeJHSSdVQTjgD819vO04mRHlC
kLYLFJdWWCFvAAu2kZCop4umNiCTL6/tzvGWJ7bwOyyZCR85E64VrmGqYcaJalO9vLI2iA2H79Xi
ThjmXbi5Xw5uQknfe3cOiOxedxkt5LfUvGI5mFfC6suB6w66HfZTpIRIr9dPbf8gGYIR47yp0lh1
BZV/YcMlNCR96Ffl8L4i1PpTAEMPPInPpW30RHVBiV0DBndNzPa053aNc0fSiU8i0SD3IZOBjRNM
wYGH9jowo7bVfc4V1x75QY1EsZYYun2gx551NiqaixKa8TjZjsjFb3SbllJgulBn2hsew7lDlxHD
FGrH/ELBnisn+9o7K9BIFJ/d/H+98HkOPb0L0YNkbfcL2XmMr3VTzIgzMa+9acAP/61YnxfSQK6G
SbeKF/lwdkBwVneZYMorQ81aB/vLdULyzTKz/PwfGF8f/R1zh7w3ozc9e8zvapqMu6WkeE9ata4D
gvDjWb37dxGFze78OQk5dkrUCPeQeRC5799kZ24cJy71ww5KOyGLFLnV/lsdPdGzgVJwOFcffd5t
anCgACzkjrGe7aqVKZHiZK/P7AH4YGn9kk4ueja+DZZNXYuc4yt+QmYAgIzw/Cdf7Ky/AbD0ICFE
8gQ0aXoalo+lBuPbPqs7VINxj1k04eepEKQ8FPw2zE3bQHG1oin3yXCHckgBeMIkcp0hOMJrNr9u
PYJmrCquJkqXRIiIeqNvaet1eqbqkuzXe5ZcsR0tA3PPtYs2dMWRH0MnAMLi9VBgO3MQFusCBzvK
VFm7GqfDC+zAhRmWyuENwcs/OHNTxcoMRetM+j9kyJYlDXDTM4TTJ7gM3rVHOlYat0QvuxcoAkoh
wPe5rhib3c8MGouMORbvk2JHLS7hXC43NPABmBxXXPnzJur+V2lhVJrL1+0zGGkRG07fkmoUbzUa
DiPTeyFIgQ7Rn8KkIc121+mzFGfV8VkWnyUeDSgEIIcHjfAc4xq75KkSZ3exmFxPMsBfjmDMnBe/
93ldENBHc4hPmfaMhSgb0s+Re3TZ2AOTftmA6AHtd63KezPj1uM2b2BeVpi1RcHrcRmyrBc+vGVd
4bMwyfoKzYdOQtsOPAVhajCDDeFmb82qSw38DsNnviMaBjrz/KVQfWGv90S9F6+L/0JMky1BvNGI
NGBxGK823/B4saG7XqX1UMOoK9OuZE9gpSQx9Qbo8H9px4eVn5DVfnajcDf9bjDXy5kFw1vWnVZy
paakTXlcGbF8xr9umZQdZjd8FlcL+jbmwOdagn/xGtOYLbRzzsDcYJ8E7/3EbuRipdBXOp/T0xe5
AZxkXRAZLM1pbx0L2Ar+n8sg4a4vGkovbSNDJLtosCa6ihZSGtZsIiNq1rgAsxCh2KiMHdxvm55S
TWrXQnPilXSJ1A90On/nZtEyIFRHkQqQMtBnOErhnYRXoO8+fL0hh8taw4F5o6Igj6vtcIJ0DH0s
73XqTen9S5BJhbdIUUK7A+LpapzDGzkd0v21OZbYmqmqsy+3lOwLBaD3o9FyOlkGa2q6dXpMqBbb
Rq/GmX4VROjdyWmbvSWAcn3jsEdzuOErBTAjmeR4PZU0hqwKTsxkPKz7U7Z0aBIrwwhtZXAP+uKw
yL3XVWIhcMeVZU2jerQzhYktT7XvRvllw6ZTAijaPwFrRJM1GwFoWGnRpjs12uCSTEeiWe1QyTKV
rDi7AacZ6aCdKsFcnfvWh5ppt/v4qcDrx655srPAKMmylCVVxSdEkn5w8J/2MiBNQj510HW5wh/R
bL+l4B4vsps7+HcvRKqKcEXpSEpoaFW3QihNmPxcqCdqqApqcKECZ9NzlZfmgC3QhP2Lim0rWH+m
tjilVAxEQOwIPFNIULwxZn9Jb6M+L2cvUmpwA9Yc9TmsmNd9fYi/YuhN5sKuXNrYfGtxq95DSORP
JUs6PUybwaSTjCg+DOv5y24Q6y8lHtz+7aaF0NNyoFVlG9AFDGAA1IhXJrIV5YUuQr8dxcJTOBCF
77eB5Ywqw1k6nbLv4Icvk+7BXbU5yl0KN3enVFaeO4dUDYTHO4YjPGH/vgCMJOUIPvBh+0B0fXqe
udpK2uZ/9PQZ4SDurjC7m+N6SlC6WYoCA7R5pQR654lM7CmRLRt0q2lEeDxW1xE0osHdsRuc3OjY
Cn40uXyLMuqsojthj9w7JVA/gkOyQOMU+5vxs9CtWqGTjpni83xze4QAvZkqT0sUrGnEEL9ZSvv8
qImsfP1im4+WHSfSrzxqnPpnUFho0thaE4HB8Bv/OK7/GBSHwk8szCBRncphxlSGm/r5WGVAzyPX
VAB0fjZuy3ITcyGRX0Y5i6bKoZ3yspWOgpyR4QuFipcFoNZddAgr3Zo1+jwOXxapBc70RKsUFKW2
R7ylllExr4Mu7vO1yFu9/LJ8+ABDqnzqZY7lW/BfPsCAPK1xn4poDIN1ZLD4ZCNS4Qzf7ud3yaXf
U0B4arYyWnS4Kc6Vd6Rdb5H0ZQQ9mi106BQjcP7EwhZDLzpU5uV9O/Vr4NR6gIIP9MSp1xWjdZ+6
2865u15qsav9YSEMdl+Uvbd9PyGaEAJNXj5kxfADOoaCkE0ko2ZrqbqWCFG3zXgPnkejLA/4e7x/
ZuKWpwId6WIN0+YUSLi7/auwDpHjgCSPDJZPxdO/JddlEBzTaAhfSxilAChAxmn+cMEHoEhozdu0
xej1jfrvm7GqRp0zZELy8qwhoIYmQYn5oThb+4fuFy8zLc4AsxZmF9XrqoZhyzQpabH7PlonEMwG
DUon0GQurm75qh7W4nFzw6dCezqGLsiwzTkVek/ulLYlSKf6zEx2hsa/9DTsrc26ehv6iNvV9kIO
lpe18SZnXPvp8feUb6rbBkdqjaopA0Zgv7aPpJRNi2B6YaclWNNT+wm7CfiapoJkiNZVD++Z4F+u
vnkasfrUjI0ct+hhT7n8FybRfXnkXX8sQqaOIfhUnoXiwWev87VnNKyV/gM93CIK4g6VyNPq2s3s
O/2xkERn2fcOI6rAL+kMvGb+hz2t+f+S5sWDaEejhXNY/CBkc76oeA6Bc/cXldcmVhtL+DANqfkI
BPqNf//37Z2LS2dvR4eDFdEQRV6CubtcUW5seiNw8BiseFji8dUSnLKmxXMViQeXqAAEfJiMVd28
Kmtq5lqMYlJDaeE9aUOFzqRYzo6T//QQ1tRkOd1Kshe4HkKr6LCK8d+bseohBUrpNGFaP5FHPlZg
9A92gvAkf+GIDM14xEUn8l8WjWXXW3XnvpJY+0B88ZW4LzM7Y2l9PqrfxwVTTQ8fn7QqXavdwQRt
RmVPyYJbuJe3xVpjEz623J+eybbHwxksgnnFjEmdRbHmAiNLxsuXykIA07pPaMRTvOK9sTffMvIU
fkPKFYH79wlqC9vVJZoWlJUjC1njcY0mm1/iqk6oneOuHYKz+JqW3QThPwfX7RowLn/SuRlXW/+B
XuKM0GfJfKh48l5dD+oDgCUGjiQrT0EFeAUKkf0p/RmoRNzkg6Ex62hVCfFdsbH9gk2PaVUjs7xe
wKvEIe/+6ucPmulRRVEaeblrwcOAWeiJHGd0CCVMtZUtfof9DF6TIsYEzyJH0NeOK7Z4+lvKrOZW
4JsQ2KFA2GfitpU2zR6fHYE+5GEMMyPUYMJ8GW7fOuV6uWLN/Fpn1VE4ZsYNQPjbgzM4r+Q4DTTL
EqgwMTniyWDvuWkOCGNI04HLqJLeF2DjaTAHnzYQEf+/nY8Yk39Eo7C9HVMLRNZRUbfkZJldv56e
Fx3fstH1LX0lCc/y40+m7Eh1lnpufMX1x2m1WJw5yQ0MCDMJOxvjU9gDvYnwSk3+LwKRKO6hvPNH
aP2Jsu39y4sm/T+bDWfuEeHChQxJMtxmcWyxVGOLt4LUV6yeux1d1fIt0fCvIyNIDmjKk+a6HxMF
dp/iAQDBnhNpon1hGsdzkMfFmgmPhXI5Yq3jl/RK6wyvYrsLApSzaJcTC7O0UdKAsWdK8hX1ZE6G
KHLa0+pMGtoFSfdMSzYG+4CS1vqq7Vy05SOHUpy1CbsIYaD4wOeB/m0y/QXM74AB62QmucHMUo/9
Rq0NnfkyquepxtmqNAfhUEef61CG6Ct3v4T4DpSzGRVg0pndjRSq7pQHwqNxsMnn6oewCnOeVd9b
dr4vE0ipDVAU4FGvwx0jNmNIHqGQBo93ODOci0LdPVCC5cNKi9pYajm442hl9Qzv+spFuBRoZb46
IhhsazsvAEZdMOcR6P3fxv7bK86MmW+6OMzFn6zyUYnMaYmmKUc7BQxXCJ8KBB01ov+GK3eWJYBJ
T8wo13N0/h4DOAC9aoUhoXW512PjIRe7ZPLIrAXVZpn9benvdK/+7n0XpBLDw/j7XvrQ9XOk/XVp
NkpGhGabCT73Wjb2EWhRWQiOA2rVBpFKlb6aiHXivoADnTYZSG55W4CRdRreLqJDZx/O1XARb3M2
NsiSf4rdaOukV02ox8B2Mk9NDsuqBMsTSVTAqVtmzrjFKP68WrNd0uXAuiAu8ZOE8ZxW/M2ICiM0
ekwoqnOni/5W7CObbb8A95dE26EBT4/N1uxnf4XcMCVu/HiBJvpMS2j5uKPQPRTQSKaqieWn3f3G
Ut9wmJv2AjqkIVVqCAZBM/Ap0wuWw4mmwKiGvbq6Pp2puK9fjhgOfA5XA7r7lpvbuQh8PIJzPgs3
X1ku9ZsxyzejgHXNHHPC8Lv2pgK3aWUe2p91esQKKuRgpepcxw4KX4YGwop5DFhYanIfZJbR+fnT
BdyzElRps3XFOe+N3UvBn0y6UCwbGWbhbPN+4T4qqDlfypH3jErI2MFozWx1ExT4V9vUlGLfPIeh
SDp8JwIzH9aAySmR22CGSLD+qDV1rBeYKG1qzIsqhgck7gPSNVUK9moMllzno6x2p0ahb4Y3Yulc
h1rXq6hRhjvWVbdhCc/Bm5IHCGi/p8ioEUbniKEHHLv4twXT/+oxwl+mxtggqehAOduV7f1/k682
dW1JDewfhpggt/tg3rDywooE1De5Sjj8PRbSxt5d5quVLkBE3ihzpXNBc7jdZHY63E2RMzlv+GYg
CJMW1xGNtMFl19Gx+qk+FKiXFWWHhAmJy0+L4gUAHpOdOfSd8nphBN6yD04+1fXVl9FCdm7/7EYo
AKli6N/5pTp3xSmko8sAg6X0+MhAsod+eYx7Xw7D1O5etoM96olQLvxg7kWYREC9s+IHd1RtT+Lc
BTq6XUr2pm86x2hYEsFc6frbTmafRFTSxE3gbc0ZH0xUPlaXQZcHPnGAt9QE5Xu/daSpVfsHRe/n
Mh82Y/t6Uytyr0cJ0GDX+AgVrd3bCA+ZiWjzZtLr+Trq7uvKhK3OMMeBjyb689URJqXD8ot67OxZ
IwtKjbc89RbdtHp8e8bozXWN/9rdB8BbWJTBLpNgCz9EzF7PYZEvRN5HUf+g0Rk6Rd+kCwX2P1bc
XWn+WouGangz7kf0D+2uP53c5M9sP7Jr5tnEDq1MCxXlCD/1dDWELUHVHOT87zFe8egKAZHeN+qy
aYoAmS4ecPjV40TVJfw3tuhj+Y7njpBD5kNOW4yNHn5HRbRtDno5eXUJz3Vi0tHXr7MLy/zpOZe1
oCfFwHyZCYA6V7hn1va3M0Q1p3+ZxIl6j3/jzDoTomcMy5R4t05uwvMDNGrobIjYHLdrPFXtpM7h
+mRc9HZ9X55Eocz0tb+mZZJsabbCrREyo9/sXZ0tMgK51qkGDF8cQTkoH3vaMPipVC2ApoeXzv7+
YiYN1up5hAFw7AkOwpZXG4Fg3yXo45S360SxahmJT2KVF9fkerhgRPsTq4TroY79qCbzldxbNd8k
hHc+zK2KRN1N12iv5NfRj2Dd+i5xr6AcboztufgXFJryUIIsdsJVJZbf/sDVq4ulvX+od5UOXELP
YSpJ7MQ780YBp0t4DH74j3HOVLiHOPZGFa8bIMvi6K2a8+GzYqj9M/GtqbV4GxnXLXZdVPFwZgir
mfBFfauP447nFdgKEVfVMxFYyjKUWmzZRjYceO4oz/TQtxdOwa2jmM0A2trRtvCB+cS8pgj9IVea
u5Gp6p7FCzlUB1hbxD8tRcZ1WBOAWexevl+MM+eiI/+Hmn8FSZmMZYi3svxyxzHje4ecMRnErK/3
Qra2pu7v9sId+5n7MljxlI0HMno+qULdCxeOmsQgvPSulncQIJDPuZpNJAqa42yTcqCwm+AtInCG
Ow3O6sQKBAcLmGxJzMvqhvXP/1twh9KEghqkCqK1r1W7TFRDFf8QClbxh9bvPQyl83fRhAPF1eEj
qPYpPe5QO9Wrxcw8QNu6rMeIMCZW28k4lggQC8IzU4pWhQBX6qUeK0JpgwWc4f5Q2DoHTwOQOj6T
I35H9wHBQIAqPI/ivH1oeI263szbsn++pIXi/56e/XFFY+6CAD5PVAQmhOZHPnS/cGFByAtOdgKj
i3fzCuTFy6/4g8AVWnb7NcdCLL5x9YFiTNkwB0YxtXk2Ioz/EVhXOcTmnIByJxoLRPDbWpS9vB6c
4OVia5HdW1dhxhW/I1xigi4q6+2hV4B1PfH5VcagIpcfymy2y+embdK0k+eeiiDJbe4k7wapD5qR
uVZHo3Ww10FA+Mq8Wq3jKhVliWV9DvBA/sgW1llMrG5AagZHsoZdB7maOZa9uLknh45P4ZlP9l8y
4e3pw/kpKJ4SDCL6Vquzsw/VEyFhQZxEEcKcmFWItUkGKAG9e0r8shvPF1ck+Zbxh3v90U3hqQhu
TjkYQHdW+0y0WocWKsHBi1dAh13hCIVNPqHnR3a69rBq15b2uEHrn+zNB7Ixl8dajIv4nQ3bL92D
5X6wk5/0EM8kV0QcaRTXFdbMZyk9FL+AKkBBgZUQQmtQK9rtm/OBR8qf+5dDoE1HTZSoZd8gA6fm
neEzvyoFomBQbyXC+6+IgX2RzOfmg8iBY6ohHAu3qHEJijy0326O6Y0DWw+ISiPrUJQat7E05A8Y
aUzyEFCIjF7B44ezMR6MQ4A7tMQW7KJNVmxKLhTo6C0q1hocs7WmkUKFZur1+nzUszP6gaUmn5l8
BvIwRx9vdXzoqBjrrtcCwVNsrqLSjkHXvF4so4ivvWpmeb3oXqeqTXjp9UsMMCqUl0eqAjf6LVx6
h9X+ZNADaLCHagH5A3WP+7i8ir4ZRRKGh3v3mEEEqU0MRPtS8VceHpXM0d68XKFYMUiyBUpRQxht
uqV3WdltwDGipgr82g0l2thCpOIruMOzZG7wJE90IaayVEu0FTBiXBCSj2KBXZXIkLEvZ6PsDP3v
UxLtozTwRqtmAkqJewjA2uLSUtcoeXctF894N26TDZJoHNfcIBBbHRhoP0qyR0mkTMr1r3/onLMJ
HPuegBqkPrpSeNfQUM8AZd1FAX+VXapUp7crLnlzySTN2/AtVbn2lISNBABL+pkM/AIurZ+DNfCO
pIauLopCJUZDaGLY6X8D+DljbXDOFLSNtIDej8URgkmQZw4n3dtrkkFpNopxJTLsztUvWVbafKr/
x9ts2GoixdqtDMZXPOT9h9SyDyerl1oribrKSg9VaEyUad4lYxnvHiedWNfjaOJrGyDtbEv08YvS
U4tPKtPPy/+VkriKV9ML2grZGqBOvUj/JPCziA7+rS/ax2eEKPN/oUWzTsqir6/w79ZqYZKpemy+
iSAits5ce2erTvGI9V8+r1Svmh0DxbSetWZ4QAYoF9PlQYCopII5fvqqchdJB31p4A3mkghToMZK
Rv6bEPK1LNofnyzJttMal9emP9+LbSwjYxl8PhNaOfRGHEf8FgG66kiParPd/Yc1KKmD+0fPVaiZ
R3HDyUxw5YdQkCG3ssJLp+cqAxEGFTOatt5C5VxKDob33mXd8tByhse109G/Q6/W1fJF90l/pywV
VO85wI7px86QJu1eCw/q9JglW9qyjzuTCWZjvW3MnFUohEZM6eD1O3Ge7Kb14eBx0FtAMHRvv117
3EBS4rtFaKVxWMTJsqB8EjXSmX4yy04OW5zwA6jU9tk1su51rKM3Emren/wH6yiWRTfW2ljgZwSR
/O559iRcrY1njCVq6Qww6T6PHj/YYd3ot9bu9HPvg/FLcKmqJ1aPpM/lqNGzxEm7+Er0tpiIwl4T
tJCju40M3YCnrgmCDjD85TtAho8d7hTyBKOZG1zU1K3okaITg7HFBYE6ZH1sc+Ltkn43bD7OqEb6
H1RzihM+Q5+vrggSGDGZia63nzwvOBpLau4ge5cBkw+pZ5tdROZJ1KWpaOIfd+yeamCXvXYmrVW0
TfOvydDCXakCUY0T9FMCSW1uf6zc7NQjUc12uJ6e+0zx1/cPoaZokuvoACgUCFwHJIERta3h3ZbR
bleVjmxzu+SIdWO8lQI+k7PiyDgMDz2Jp6vJe/ZA/52mVKxqo44iF3QeEV9zB+8bzxyzCXajh8TZ
LGfc3z0l3V4MG9fvYn44JWrtpsRDJ7TPjeUInBeVaPz/EsZF5SGFgDI2059SP0qvqPjPN5wxApqO
Mdp89W8bQs+/jraS8c9yL7AM0toucSOcp9ncXrEA1mEcB/zRZmEDKgSc1bMCkdPpIhJxQu75BEof
UNFme+2wS2mQwRYgM6Mpatk2mdhhrGL+QpwgYmrDeyDe2rdNWovA7H0TR3fVytxzrKzWwzw/XgGl
uryrL7CQ3QQUIS75agv7UJtHrHujUOO1lE2VAmzxk3UWaNKVyi4QGSt62ZV9ypbDRpuZyXfkl2Gm
Mk32yZS/DwTeGcSkJaMMc9eeUbinpWVSRgjrDFHYSnYLrHRx1xJ4seKn4KIK8Egxdrx3UGgi2o+Z
Mlvq2+qKRtR6JtcsuONFuiIwqRjBiF6oEOM/0pZwRgF6PZxGmg1/+8jZaFL/hJTaNw5BEqGp5XZX
bVC+6IupuIhMDKLd9CSQ5QMNbIsdzh4T2OKr3VBpVRjifk634cT0WJYasFqGsgg2kFYZ2EyY5d73
TcCW7/08TCwwxTMV6Hq662r/u8owufZFdiLEqBOmZlv6qXK1FThsPod0E0tgPRoTVdHhA38ZKKal
7ZoGY4bnZgh5ttoS4D5Zp9SP2KgrpH7kNGLq5xKB14jtosnn6UYazcWF1GgS0Kaydp+Q26NQzg87
mYqNjvUdvpxmWPKi3h/8zeKLCQBKiKR3CqoTXHkhuhN55jStzDi9hQaULS8aEXgJ1CF15+ZlfF0m
G7Y/y7fJTNAQzdFbge8XRGP7Hs52pjC4LaFvGHCWMr9H9g9lHK8BMN/ItOlwgB26vK0691pEdzvg
Z65qMvgVt84eK/FXnTk4IRJHSrWKqNZ0rvC+gCTObtQeJFPWPGFYfUZMvZD8jg+2VIIYGpm+BjCO
RRCk9Clrl82WwEh0vDCtSsClnmH8xXDlKVw0M0kOKCe9TY0afAe6XBpzNPj6396HEdN08zbCbB2Z
zytWq6BHZ3z46X160lUH4lzvNaRWf9hnxWP0t0Qo4sqeQaMpiKYcKtsJ53tNNBgMm6F8BxCHDJ8o
qkGuHDStsp3os9ty8WLXV+hOUBpHSVA+3HVXteWEBD8+fjkwJRqimwMi0xlc2rxtjknMqvfoaW3W
UFsMQJhI+tmBjxoofRmJMNlpHoHhUCicnNtr5MMxe8yAWcVIQKKqc4uz735tdpqqCH0PBwQZRtSU
O387+sFU91R9K4Oq2XtQ+G2ZASZScb5kbOCbx0gX59oD0/K8U2jacon8NBU+Qry6mqWvB4LBpMs8
LMR4TJh7uqdV3Giy0xSZJAaVk5lw2nIQvE8ChA95oPG1gxotWJMX1nBNv2dcZencJ80LNuIyqbL5
MIPKWCDJCJHwgks3Gf9u8my4nB6JpiMdKsdFSZH/tUYAf8fwsl5Di1MczmtvXHyWD8/rYh6E2Elj
Y6ERdwUb1eR4O5fBqusu+jLq5R4B3j5kioPfpG0GK8zxfSTXyXnq4iW4gVO9O7mbTMfI0/0yUt1n
8zDphhAX/0NV1YBtBgkKUSsGurBsQGGQWjYcp/70U698smAqu8f6svF4mVMibobIstD8dq3oH0kE
4eN81lM7x0LJ3U3EK1vqeeptNoXl+1ER/tuCof3SJPH58u6qQAXh6X6xhrWIbI2VRdWMpEyHSIZx
x9BvJrZn6jIXDN7lOijthplOClKRbMoDGNwYDDTmOQnNxKlYMDtbeW3gYAAnWmYNt65tWcgTdQu7
iR1byJJCdYJm4Y8SuvVu11JA4wUTQdVIL39b1h3f+GE0gAiMpA9yJWryzrGQrAPyCnsrqa5pRK9D
ou5tovsMSPq0+hzBK76BhW3UMapK6n1RwKcNTZ/MlLD+uwtvYG0MlQo2irCxvlTnPqRgfRixzStV
y6iCHWcFPZaSJFzqk64lk3kHhkShHLeiMzKZqbd+jCf7EhKxapTj/DF4QyyjTAH/QpUt/qFSjYLO
p9pWVTh1DQCG2lY4R7dv2GwfRk8nJlvWwp2RlByp7i/Vyf6QWMrqcdQN4qmI9zFK+enKp+0rBlTp
nafCW0WZY8JEaBVnhWDtO4tenwiOe0e3RfEBoCpicb8gUAw+NMoZpgNr7VaaQHgUW+XroY9eid7W
NAcp0J2frCZCWBt2MYLwNn12uUnuS9T6RCOT04tuSuRRz8uf2eLmZRX7sxVuCCD93uVDXziiOa68
c8w85N+BYjvoJUpe5PGQ82/essQ8Hc4VZLr+b/QkhIIBsRjwp5WxZZgGKEZnJdhVq3xf7HYk1F86
MN0AGcE3BwiIiAjYOvyDKCHkrc+IA58hCx65faJGnYFHZd3D+Km3GRzdpEu8t3QeYtDkwQTLgdwR
KT/cRUlH6NHxCAvY7J/PzUhLZB0Zv4P8ZwHwmSe4/TmvFCBNgat9WERsoqyTNrsWG70AUIjQf4Qw
eWzatrm/QMLdBAfIzkElar938IIoZ50aBBGzUX5FZBDO+4l2q+N2XBqS2H2LmKhCZWJVP2mntj4t
K7P7ZTGXMbj9F8QFZQ+ycqdLraLIbaCplYdU5oTeA9Zd43QbiC7Xv+sNEngsmX/N5vwcvP1qmlP6
sh5IdBFUtleJhGNaSxukzuERWrt16UosiJVRUv2LrV+0ix9jTeBbCZDSwDn9u4YTvsQudrFnMNfy
2ypEtg6D3VMzCBk5BvRJO8Mfm07DojayJyvs8CBZp9EY7NpEeWIZugAtDiOnA+7fwHf2jWRgc7km
FwjOilbqDpbi8MjV0ObN9pd0oLpIrKnANPxK5JuvsJAoqmSWIhjxYxg3Lr6zlkejFX/+yjmVM5TL
krK6rVPbFopZKAutWqv/1zRhzA++Bp9Bs7au5FGhp+nOH5sc7+0R/1yKNhNJ2H6w7qctzzeKWJGt
rc0bj9crb4ogZg1mIN86uXiGu6V0NqC+NJ8Q30+a/d45gcCqUBz8Xy6aeUnqTrEHa6++KJcLimuE
JmptlCd1eKaSy3pJc9Nc8XwBMEFdS2lg5iYpgAHSyXZ2A7O4R3QvwoQ5hy8QOvC58VJCEQUZyHe3
Y/VreTepWyoVviX6RWZ85HFgO1zxoqLHc6kHAsQnVk3BDVh7d+WpZBRJMf/6xyDPvCndm2svIjZr
/HvVyC7+C9KVoQBCLL76TlRtCsIEGH6tnH75Nwu8LMEnkx+gZ9VOuY/vJ8SJQ/nBeoidtF6+gxvv
BQYU3CltL1GWB2/ug+qqDUY51qnDXlpQEXdJhuOOuryJs9DrhVRH/7J+lpkaan6wHQCeEu0H81Il
q5bHpqkU9nEr6zAIq5zwJwoAEL5ie8eppvbRFRni/jDV+oRFyo4rQ+gBL/UtE+Vg9Figr1ZHb6Hx
uzEX1fZzYLOd2Vg4gYYN4SdRdZBRb+J3/AddXcyV8ZlTPXtagzGxVrj/qmoqqTN86bZF6kxtSAuR
kRuOEfYoAke8S/W2+CvEYL7A9+ckI8I4MMLPI3vxzKQm7zdPMmcFEBBC9v4t8Ka79/U86oDrXC+9
37TXeYiJUp9PKwax6B/1ps1cHzlsQSQFMTIWiaNGvwOtRMCqzX82YYnrMsx520Ecbjzuu9gAhCmW
5h/xXxSyBh194exoaLKHQJXZlODBTja7OTZp1J1MGZFsdMZjCA66nEVLXQoiUxH8CRNyeK03P8lZ
oX2msafhesulEWTAE/uiayWQADj0N/MAx1FSCBxa3b3Cl02TQQa6im81N9PY2P1lPs3ejhMhPpnU
99zej/Hr34GHT/eWwhA0EtUnqPJT2wct8LHUX74U7I/hqYKhrlmBR+qUdBukXwx19/yImFz5gMte
OridBuR88r5DcVPqpoWQQNaALshnrhZJJCGbTim0023YdL/4roXIEbVpd0/DEqFJ3k7U/j6rFnjv
DEv9uPPcVaQAkgxqK/JO7vIB5ADQO6xQKsDp+N5pNrG9DRqZQEJoGDJswoyFU53UCnQtfJ0TWAWb
YA9nUWX3oqvq9liEIYD53/pAEWJXFDpat0bW4ByNOn15MhyhAwMGA0+Lz10Xw8UtpFs87yzH+ez+
kAwthyZLkzl5oWIUyfs3aGVZpjJo80SLiUeJn1jGwGA2BNmo9FEG58rQVylBos1tAJyDluJUBX0+
f8WkGn/0Chr9LI6n6c7xERNAkMsxle5nBpneF7OOZoizGzoS1FyGJ7kGPTvHLxsqhqi/9ZthlIf+
gCCjFXM+z/8EhKlghhfAh3kSsEKME+hiqo7lpT/2HE5mGJHhaXbaE+t8KiXA5Repbn23G2knPC8K
e81ve+KTqY3+otuGgltdHDybNg1Qrty0HgIC3riszaNXkmoV8S4HKfynVJXl3LIoSGZ9ufCEwJZw
qxiMCVYLMnmAKJkv1e5rl5Pm932Y7kzo9o3UAbRUk+QCAy2bq5EDWpC+J/JUcUsp1ch3SLAYUsoD
D2R/snwOy/ZT/ZeWHpxKIHFVEXhdjfV/ns2pwPaEYC88bd/KdP6nEMjMejv6ZEPFYiTCiN97Cmco
HlGNUPt+zycskSNuQ3oSr5Ux0g/qQUgW9UII1XiyH++7mK8Dt9zD9mqgL4oCI3TS9emfjix4VOlu
6ZVv0rqGBLfV6U3Zzet/gz1H1hQ31xTbN/lwqm66GModGmL+r7SPAhWvT1N1NFu+Cp8AQLVLbzhl
5rbJbzd+u0rG8x8JPNRfF1lVO9kql6Gz+K2g057mRX55AlqZSjhmJ83LDVPKcuvJrhbaCe6Qcv0G
5JiJi+i2QlNwR0+5R2peNOzkTOK1CnW58+C+lXFx35LFK/8K+7Z35hiho8UmbblJCpJ2V0lgshjB
HFKFVGT1RSHzMm1GiARC+2/cEdZNE46CNO5kLwoqMUsMw+UW4Vy+N2jFYpGQlWUwfQXZiRsXjGKO
9yzAyNKgVXKZwobzqXyEvV1QsgBDb6sHJDKYsckrc6sHG1yiZ0SwioTZ+B4eQrzJ4zHB8AtL01iW
0HT2hTUG7MIXykNEHb57aJzI2nb/gUTVfCcnaV2yhAmIzFlhhqT05lGcj6M7RCXEHB5jF5lfhkrp
ZBAi+NudcGymFyOeFcDW34DcCnGpFplyKvfyAwbe4hVHLpBqPhaUYuSn8A2hZWz3ipwE395vRN6I
ldcEGKb2eZPRKKXMbtJWQWp6DBjI5neVDZD7alLSkwxNukscIrF+5vGh1YfWWDY2pUn/vbfPap67
mKGsR9RpRXN/MYb9lzF7qu3FXurcVwSmrVYp+YgNYORMtogzYpEs3hMUdRPY6TjydyxMmVKZGIGk
CpHa9360xW9Vl2KB0szZ0sJSoyp61mDk1BYxBfakaifikRmsmBinVqvWlcZdIHT/aGOeE9ENm46X
ljPaIWFFyhMGWLq9Xt4VQ2dThWd3ND58xPWR0MgPBUhEsKlknadWmKbxlz/mkWdYsicor3D/4z0g
hc1ESPy6ufXHgaGRb4cL17qno3UZktRdt8WQPor4nT/nMO3eMTUZ8YL5SfuZQBKGfyt0D7nNBgKV
xJpGcp2iaqza2dWGJdrMqBDN1tDJvC3zB4S5e9oGxvqAXGFZkPAUSIOfxqO1XQ/JCg60YLn9f/Wm
plq+RwwRas5FtfFw3qMw41fjohHzEstNJZQy8a2zkvBFPKg1QzTutCRI6OnCj+USOoRZ5tW9CjbS
02URHEpYKShJKd/NciU2xaFK74YMwJsK2K9RaaGkS8cSjDINp55p+BRHHEURj+yNjko2Q9ufigP9
zwzJ7Y30YAx8ldLXCNlXKzQjkC11viVe6uWttob/twnyH7oyOBmZKWHN/NUP4dmsDb6ZHm47kX+j
Uvishmk9JVn2USrXBMi1ORZPDJXaAY4s1ep98Aahc2EOpBapjA+b9jzf1E0Pzu3X9dX5rzzo+6Q0
wgPs/b4fDC6vnSK5wQAma0YD0QEuM4dzLdOmhY4eA+20xxPaR7vbIbZKyzT/gPjuMNLsp+UtLda1
E2d8U4fYZ0nevEyKOGqC3qCxdoNkgimlNkFBmmYXcRTraeLKuWCY8ITT1IXsPSiFHJT2dA6mVG7F
drqMC8Ih4b09LOC4mKKk+Hut1QrmkuII+VvafvEnWWPdqurcrvfLanDy5FtUFTa/+CXkiULm1a5h
oV/S/L6ZlGsY0jNRON/YW9yzQxnTkZ4bNgLuwbo6XYwPAJa7y3O9Gm/jVWVk7550HA41WeY36uBF
wOo3j7IMT1ALih3xFL2/2yUQWYz9h5Hh6T/kuGEcPb13I3QA+kQmyLbP1Ap1ho1b6i3kqeoMoZkw
0EY84JRWiAL0cQ3UyD0vtY9IKlyqNB+W4fEudnXDlDfU25wfVI7rQeW52hC6C4jg7atiyotQm4hS
jQupjW54sNrD1w+gmXN+deXtzt2DRza8XDFptFY/1COokwlmaHECJnTWXjWxDG9KWCYN3jiBpdnA
CSwgOwK7urJJNgkqd7ZTHS4SaZVhvrfoInLKZlCrqoNq2NPfRO+GrWV+UwrQpSp8E75AueskGFIO
+5S4uwM2iNmsCorj3D8yuTALTx1UtS1R8gdouujwFeD4MxCYM39HmxnPcPyuAKQypvSXHYPEn1ln
UQVoh2MznKau9invuk1Y2Hux2K/g/1sSLGg4xxu8usGQlmTAYIXOfZAopPmsAEBfHe7LH4AX/w3F
n2fOllN4SLasbeBPQSupJZY4lsB0hdy9sIEl/mD4qxMrrul64+rUnDjC+98rzuiZmqZGkiZ6HgmQ
1TP3vUKCPkOf0kaPhp7QmC4SE+ZHY/LjfIfqISpWXtaO/S4GG8PBnJKVO2UMq9RLKLW1Z1mUUkmk
CoLatd7Cr1J+jlXmaIyCqpP4XJ+e9cHv0tWuRnij10URDgyQ4ZiaGQ6g2JBNJwj0t4qorhfpOyvu
OiO3Khp4BS2k1igDw+FrkYXpNWDByNYZfAL+IPhPjwToHH2Y1/fVGmmDdXny3CmwqvBB6LSW76ot
vESzD3y4ETNCivXj9M2XUhE/9JewSZ/kL/NSceXsG2FDLu2T+qFODzJZYLBK132PqGyVKT1OiDtW
HuWR/CEPtckZyULtZQ8bNaDzGv4nZvrz+b7hRK1A/7K1GUayoxuOyc7cfwjWndUsV68IJORVdmkr
bEeS2ISWbPaeNG1LTuYrJYWyGaKOe4JqrygsPG1WILq5u3ViNlRzWBzbLVnaJJ3v7bJXljYG5dwY
JOPmqug4UANkVyD9nq6ZmWCOfNEZTkFgtIsMKfHk/jVRuz3Pml6WhpmoR55F+jxHKx1IzUQVnJU0
Xj1wVYpsVM4SrpeDf8fj0dGZgyrDsBGQSgCR6SFo+0Q1IkqOYviNI3ohHq4A4m+NGuMdytftI3pK
oaBXTVSb2Iq5Y1+ZAbo+y/ciEYXWNsSVbMDUxvub87nLwxDo9HnFs3yrr1zu6+oy+ull94oE06TU
PaoryqPvAaNsqDtGG2T3w+Jaht9nqHme1vao43RG6yACg7CwmU52jy9GA8lr6aQkedi8rBI2LCm9
7liWHxsLEnfszvYN2P/bSfo82f/cvOLHcnm85e9TgLgBz8uiXch0ds0ASXRmjU2hqcNosHbWH7Nf
ZelKxXc/YvmOX29MuOynx1U3IThejrDCXktoN1cdHDIox09BTKIZFFn2E7+wXChEOuUE1SMqiCaa
4r0EIU9/fIi5DeBxqxTxHGd3avj6RbZjlHtGS4qk6+g7laxLDI2jbb69MxPsPelUSvG1rYPLwGuV
vAS+CQ6zs3eReBMp/GwopdAypiOgDO9y8tZiHkOrriheZ7xJ7m3fxNLS6hvL0WzfDoerCYZe3tOt
iL5hvX7Dlj1a5tKGfeXOlPChcCti041yUp/CR374RdlaLRyEoBt1lT08745Qji7OrGQ1L7CJaZpI
oTUWHO3ci2iYS57Y/bQWfWKrjuMSSKgQ3sf+njA6O8HEbuZnbfXl9+mORPF9Yb+rs2y+/x99BLnu
XvDEmtQ7zUXmjuusrrG7oKe71QtEhPjk7JwS9LGbX75ft5pzvYtUZFUv+9pc7dNvDMz5ExD5oSOd
KJgwYKXb6MMK2apsG1WcVqXrNte0K8yQ46t52LaQUwTv1C7SJANv3mvUzOdQ51zgO3bz7qf5+Y1q
roOsvzcISXpsCet7PCbOGCI3yy//NG3YhVACOBzPHb3xKBruTbRpu63q5q0TEwYVg9MNzSHH6F2A
+7+p7xZN+fGJtr2Fxw1lFHXAmAOHN98s5VYNkSKZW/iKPzXgTqe1dqNDd2tTMZXLuBek/cl4QBDO
KhUjiNljuWHDu/yddSwZfgkrgsV4J4vCzksDZ0SAIBnMvE8mRIZ2oEfsi51hZhAgO8gruqsu1lW5
mRDuzP2Uq/U70AAe37oViDhYJ48deIVC3pIeD8fc1NrgbdDphIRVowNgWrzRLv/6QfNII2jLFI0B
8mLFHSFqpsp5eUoXjjNT7frpggMxS9UVtW5yKrW54qZ2Ss4NIIhGSNtFyBvG21yZIx0/bNviOu+M
r6WUMjYedanobhwuTNcGTvHZixyl7etnQ67Ek4yL5H0OwGOrTKP5nuHX9mo7uHn0kLbE9OZ+EYbc
VztYUwY1wsjmDvAMiA/vd1zXKOp3zBTsF+WvUEVF+P1Ov7cDcCq8wvRxb9f00Pw0JiXlps8RtduS
X42cw7KAXTltO98SQbqbQVkwIITM+zXAFVsnFLoO9o1ZuNqjidugRwx3JMCEpXMuH+7rhLIx+sk9
YgYxqerN0wibuRYdjNwyLZB4CmnuHxnULwvJe19AEzbB2Swymxn7E3BsGlQ7aSy0uUO37Fa7RAcU
a+iqIOIDaYWST9fkxTETj/YBeBiJ0chOIrSvO2e4hG8dubZXQHjVZvPo2tcxnjXn8KZIyvriIeq0
kerHZZgB/9XSujE4p9eJ+l5Guk7MeVN6kHbJbZ/gc0AdCl4W/M6nW5UFpECgC55mDVoWl13aYx86
q1WKknR1PPM2DjvA4fy1BViZE1LdNutgBo3CQC6EkyMEMM8HhzHA1xrQge3DT08igH/mh5dpW6/C
6hsf2ZD0pFPanDvm0jzKd23PV0cmksGynYzFcUdejT6jPNuw+68rJ7nMpK2tySnOxmDXzE3Aw4YX
gu8Bz6DrOWva9gs0eiS3RiXoghqZWowvXWPsoQTIcmNZYkz8HIdqwekAO4Mu/dE7pGNs3VKhlYnd
mmbx+s9gz46sQBE/Md6t/MWDB2qdusAnzRBwoOmVgS5syRGWidN1Jf3ZjgMez78R1u4Ma/7DmBAf
zTBa2wqFSfvq8jHw/W+VFX307QR+vcawGdC8kPORQTBaXM44u7ySV0zRQXcPsaNQdUCmOjvM2PZQ
hDyYcBU24gr+AprREEK8EJLNijuSRTe89gkrvRd6dAb9Gmub/oEVZiIKTFpXZ72phmqviVS3Y27c
Wa0neGaUZ2BtiKaXaSyisXsXpaNDMvkEAZLkOWKaH11izCmRERPUHf/whiV6EEjQSrNaujeRXWJN
4IDsXquQC7jenanxwKUtERlQYJGLB6oo6jJEKcQyZRtDH+Mle9WRGRVnPeonoygyZZr7VIA9aPW3
Fvn+i7KwTatYf3lFvrI6US2xhqV8onVGrvrp3uLYlgiM6Ohzryol5ToDXXxcmP59o7z+cISxnTzB
AR7I/FRBekUX8Llc7NhPVQa76nvsKpqgsGmyW6jfw8Xbv/AJz3op/FjUAlFiBC9ilgGhHZA2We8S
sVPWwIQfiO01ikqv+l0q40HKCjp0QyGmZA0sTU3kudfjiRCMAm3JuFlrwg9TOzbquBGaev6CaVEp
CCaQ5uhMoIERjOiGfM9e+yiA5W0nm9gwCDoVPuGczLBqnnOAkyHsN6l8w8KZ9pqdpt+B4Wm99/QA
lE83/cC741kSEFNZiZBT1XUwutIhXoduPYH+ImCy8kW2YbGObm8/dH1N/JZeiVfuu4mTfTTpqEE1
opayFJot/byWDRHIeOWAj8KouoJtr5qdFaYj8GJXWMg8tUFBniqWBGnEH7+DF4nQST0FI6A2DP7l
CmkWJMkvjYz7tVeYVauuFLLuLAAwaVWc6wdOehv8x3ISwViLtehe/XiQ8Bf8tRoP7CgSKXiaNYjp
KyfflaUJRhu9uW+l3roYcJ43wffSRfr9m++zVuXbnL8Z9YBCB8lhBfNNHtGEp8JUoCSXSQo1qSId
wIOD0W8fqkrsHb5hyuTqFMbrtMiXfZkRSUdYidap3rVdndJqi7ZRkBwoWYPvOItseTyE1Oa+5bn4
KzYJEZieci2va/IH4RMyrzvM5qQEeBckg7vkYAG95RsTkpbXEbmDcdKmqcKCN3NTqG+29+XMTOv5
5i4GYlSRAeKeP3bved8xOZDGyJGihMxzrFmvjhj89Rozfaom0E5mbnqn+PJrWRy/luQbNdMkFzxm
iLUnOY6xUdwqWo3XZppo/6qE4xuw5JrU4VxHgBYXygEZ8/BCD/sAVMKObS60Zd9x7JL/VHvvuipU
CTlHfJQpZB5BrE5Hpi0GUmLOm8IB2lzqR/LH03Gksuk/FALyX49VEMf49K1FkdsRFGf0vKOvmBG2
xVpVVYDZbEWJQ73kmk0DOByvOteAA+E3SGk5s8nAIAipAR+R+xzoqCZUXuVNkJt9kSzsWdHVjCwi
k3CCHgjbC7cwdvgI/OzOx5Fcl8xFtXyLT8T1F8pYJz6yIY4e2FDoFaQ6xn1ONrhJpsE01oRH/lq1
sd8IdHyhHsuQL0G1wUdPxfKUw48vHw0jXwYmIp7bo3negj64lPCtbgY4ak+wj/C8AFVPJdFWQThr
LKgxm8MYZOIKKYBhCAWNCNcaZBbGO/+KOW/KQmb3PR6jmPPHP03OvBXDWqv0JugloLJzZ/KdDNdH
UzxGRaO/oGvkFDZ8R7BqCLsRsICuMLhzOevAmP2DzzZxqpY2PR4TQBVn/3bLreyERHRc4/ZQmLJL
K+V40+Y0mmda4ZD9b4VyjjpUMufaHMJ7F8y5NtT3WHh9+w5/eKgkm1YknRrEyIomKtVQY+wEdTFL
IYZsegtSJMcj7SqShBROiszlhU/ESpQMb4R7Zz4qb+5QUPbXccC7aejo8cneCw4q7Jckmdvn8Izk
2oy7M8Nh3WYrMmKPlofMWhBwA18ROIWXJwbyNvQ/Nqik6lkAC4bxgq2hauPyeqxuEH1kjB/HN627
1alE2TnPMgQdZrNA4GO2qLPEglvLyHP2ZcWwo/SpeAtByJmVKrI1bE1Ms8RDoqTwuh7vRgar1taG
6qJvoiyT1beC9jTeTwPzRU/mC6jOj9xMG6ffiNkfTpbswezgVfT1TA4R1ZyFbmq5/7ZugGbO0JAX
6DyYXfqCaAJQZhXmHR6zvuBs6YA6h0mqQ4f1WY3fXVXt115CVqzYx+cDHf8M41irXIV9RH0Pj6XV
G+p0wi0bCueWJPcU4KbtExjlkqq+4My+KWb/viXs++qZKKnHcSHzjNN4qvcJdwfBwB2rPkh4W5UF
//ImzRwamZpPgNX3X6J56BM93HTmGZpcYaSXBccnF59hyFkH02/7nOptM41L1FEFgVlwQoRKLarx
/outJq3AqcXq/Bjoh9GMwyVky1fXvKFt6w0MN9eKM9fOgmKcNyXUTvod3GqgVabznJBTc6rfY2R4
k2xi3Vwpb3iQFtsYs6HcdgIGoogn9sW86nHHTMiq1/+d6jWBVkzwSin/3DjFxXf6pHEdnBSaeLUE
JLFspbSJ/rS4x43sB91XjkkphojCv5YeNyIjeKwqzpJp5M780I7lCoJdQtWE2UVzRXpBwr9Yrdsq
pQoOiJoOCGlwUTA83TmYbWz7ajfk5qsw4E/AjqmFbCwGO8mKX5djWbmu+mCCsEPWHfegt0UrC5fc
beE+rKEy76yW4SGHwpBgYaRrnhbPL4jonvxrp0jFuImVe5vx+51LsyRF8i/MAFEbeQtDR44Q1LSp
igY2VT39v/pZKbmA6wT2IxF2tBRT+4NfnJh0lw/e0MhgauKBWgGE5ZbcSmZkw+3a13wwHQqFm0OA
k9pvwS4mxdjhFIxHMUeOMsxyIiiGKUm/3UwmH6WykdMP+MyrDtOo2ngQ4kdYK3l9Bo/FO07GcE8N
baOtYlkYvVSMkO2cWK1FDPfQKXPfZL1AhQeUXovKZLEBerFMZeGLsP8koIYbuysHZl2YUtTNptD9
Q5lC9rjFHhqVa5/Fm+NQIJx0mhWq6kO8zNn5Rqmx6PaEpED3EF6PFZr+mvIujbF+fGXkt0y9AlUV
6hpTO0R/92wKUR7V7wtwy8CdcwA9+0YIEfKsK25+h67IPRN9UzcNMcWNxqRiui0nF6bnwmMJrjeP
HVkHB4Anr8wUvJtA8tB00/nWWWCFPBY+UBXb3TyeEYj0Bp5ebFaJwr/MliPejiIwN+FmlzOPxM2x
eStk7HhKu8MiJBgh1rH9+rdmZ2GwIN9PRGAorPDB2Io64mqHuCQCHKjL5npxlvTnZAbIz/eu+nfw
ajD/1E2Myhy0cCAIjd4fO/oRb/idTRRfLh00tNhVgj71cNypBloGchpJAbzl2K7pFs4sImG7OKaw
dqX8uCdSnI4v8ANeikDm0DZF5kiJa1/M6kfXFDOVmihhBdbVq33gGVCCx9YpzXFJQlJ9VGPectdP
VpiG9J5wF8IXXuRoxS6+x0cVvJYSUeLcar5Fziii/MX6YhjorOXaIfCFOUhJqhMILdkbZtiesqIm
c20btXfPS2TovRgU/+C52J97bpEWeUh4adMW5oCeNAq7Z0P6eATk6oh+4eAuEOmpPJClJgV8JIyT
DGYIkisK9ImQoIXygEQmfPo8Mwl1fQNQU/tzCmJINLdZMaaUdqXt3sncrAe8RKEvjVwaC+TwB1mr
zDHj4YyUTngMAooH8ztVySyJprttcZyPpaTNc/i7ONeJhKAcYxANBPca28RUfZxhm33ACNR9Aj48
2/8v69wStPMZ26lP3S2zHmS+KBCt3MUB76cd8+sssRNYIBn/yJ8Hzxt/iu+XgRF3hnODOdZqwL8l
Da3PAm598G9v9roRDXUrCDlo5MsO4r+z55VmElrC3NSzjxkbgQ686jpSpgIjX47AdxOv0dNlVRY0
poaVlF+U5kMSD29givfgu3lNu3P1XdNp1BTln1P5KRG8Y9v9Wns5ad3IwsfoIgtGYlJ0EuOlhR0n
G425o63FiO3Lnjb0KMjU3dBtPIswaO2sEdOij5jTMY9YWW8Js2EddfamdEvsdVIBVd+KjS/noVG2
0nFj7fEu9MYeD9+VnKlfHKEM7qS73jmMmZ97EimTlCZyZChUWOTfRIO2YlIyBJj/2HPlACfxBes5
U/cixlcMQeTtypHgwQyPbfvAVNrGybqa4otXaOqHLcd5FAN5YQ8c/2Hk9oEgqwUCMpUzWx4p3xoC
qsyLRWN5+a2w53aOlyhysVFTb2QF8HDIS3105V1DGyZAFfN1yWAJ3+v93CwsbjUvVyigNOqZBLRk
wKi7tdNhB5FcQEDVUIVZpzACeHZC+PJKA+CFd53Of+iHWjoJWFBpf/jSV7BHUHC6vghKEoEG0Q4+
kcBl1zzoYTiUyyxG69s2240lmLgpeyL832MJPbKkBcBx0/NL4R2FkAH/Z1ZN1QCDLNndkspAhIqx
9mAAOfRt69saaJ2vbhdgl1zuJ9LP6P2Fox2Un9QSV70t6eqs7fad2ryGTKBKIZZXdx8muRpPgEJm
Xeu285K4lbwDW28NNcdotChqvRefwzDkgqT9MIQWVL0lf6hMyvmLlAi3sVUcTH5LCdTF9S/Qe6nd
F11GO8TgX1uGPj4QoFNarRq5LjeFKcLiW+ahGdkTdEjZVjzH+c6uAKz6dJlmHqY/BAd6quabOHO3
CJcLJljuUgBF7RYwTpuyjJJxjuD+nOKrcim0VVEBHwAsNFuok64nmgBB/nJVJmOtg2U4/GtNKWAA
dloV7nNoLfioXCEjqFSN2s1zGTyJt98AD8sjWIKp07Vx67xvAHXgF7TA7ysvKc9Sw8DOWqtfG4hp
sHtZZuAO2J4czFAUm9lLBDgONd6reBejylVD0jgG0IuUV5LQpugwBcBdwNoRMoQLIxfM013VmdFO
LjMNctoFGZuesP4iNwMA+CKzzXd5wUhpAFGD1p69+fuphUlyUmsK70xQL/mwuwHZPLNqBBxSYFSD
/Mm1ScKCNkAmTDepk1XhPH+P+SjdQx6n0HChYk//sXa/ZZzdx7fVmMCi1XS3Ju3T3UcMA/5bAjGR
K/1YsGlQdeEeBS3kiXIdyehqKphllfXCaqz/S4bQyfqlUlJcOtavaOXaF1gBVJ4sxrdchfQQLwiW
y+HLZC6yqzQX6iHmcdD7bzoeSzTnNQ46QmLANFjafIwMhb7nnnpm/m4+JTxsEpcbbe4+TzSsbm5U
vxSPHhis0hLMReKXTIts3UbEEISe4d+a/qBO8q52n+IyCO9Vxrdbm9/BF4jfImmNdIGk6gr9cxkC
HgjTyK9nQopsM4fnfYqm47XBA3Vj9UfmRYFYDavXeP4nXBhYYJ26VmuTLC06k+ODPtmPc/s4qzjz
LkO8QxZnazHEFrhz5LUJ0WMuIDNm17mbcZdhl+riGpOUW/rUEhkK7fYI5DaybXV25dqixIujNKHr
n0d66kGKSE5Gl8+1PvzkWRMPbSMXaxVWUI0zfzvji1P0IWHhC7zB39IZ/ItdDODQXdw1OvgAnmk4
j3g9xWhldWyy5WWqz/Oa6n8mKvn0NHqzpFCDLOznZVH0yA6UmTC4nu6HIkaSsEJ+Mc+35hMdkyLs
GTDyb8wUJuATNdrKJkHr3r9UCE+hSGA18kV43Mk8hKgH0Yr1nlaTZYsm22ovh0jo66gDIuD5EPDW
QsgQ3n5x9RakkGoQJ6QxjM/wve27WE9/ZtbXs/bTL8C/Sf2ey9TA1JPeMWa+1cWG3W3Hj/COGG6A
bup1JYZKo/FdZOUvJwkSroNted6UzvqgjoLQ12WEUFpqUgy1dGBJfXsDXe6KDrDzWNjzC4q8ru48
MnPIAHghlj2c2BoROFrv1TAA/xRiBxEpU14JsQnePuuocRbto5x2S+owI64TLfNM501k4koTXMR7
p6jDn6ppZZCyvjpnoQm+OHJzmhcaosmzVgZpSjVsUMhi+06QbqbK2Bkax6tbjDGqzY311kYmyUPj
9ZAZsjQVSJiMaR+CKeeUAPpQC8BiA4kRbaGtSwGS1tQkpkOkGy+JgIsms9NS2nndOAL3WxGOgM1v
502r0pEGcgTNHpM/dfnP5gQU420fPzXuwrcKOhvPZPWsmIi8/3EllfrGK0d+nrGHgC4wGCLKDyWU
kUG12h4iT+6sYdrJU4I58OxAnKugbGhFPfuHvUclEKdBw6Lwz7fOoRUkMcdpkBLsQsINqN2boHXS
ZfW0M+2+igms7XujNCQ89WhqMTYXev1goR0Q2cbSQhaBZnj3iKdPoBFkewaGmP0fvd4Z9KJGrN5j
r/torm5ipKcLk0fxaXBAv/hBfuRF1q3NGM3BFp8h7RDiM236/aHPiSpTEvU2yBqIP39sDQNLIPXu
iSMirwEcAyZS5WgChS61WOwXeEC8dfOazKYdC0t24JHyrdAvb3YlSTB4bavxzbh6mpiILn318YGk
k42G5tGTB5zIIb1UFpIQP9usuNAzgcHC5i6jCb5huagAkCOVVtTa2+iLG0F9qGNmEShRkUkG3lex
M8PgL3i7767ph+yymuQXqUbgYAhwnIg+fyFKvz5RyYnHmoRV6/Xoc1fctjtgU0fSUnhG/Pr1t4U+
P5y0vGtPw4FwygaCN3kDcJK3CVtb/oig1AXWshW26EAAQxsCx5driSs7BTeJMLn5ljU81IvJYi6Q
zHHSXdYtXvZSo195BrXFVGUt6fIxsLqxwHsQTmmY+kn04o4t9xc8fiTALtLHI2vfiI0pMkAyeEJ4
WN/UbTh0PSy1ymvBp9UvJ9QAubLMFH8BrbafhHybS+Np1xBm10SuJNBIdeDPZLaeKy1iQkQzqsh0
cIx43YUt1VMsppKCGBhcq+suQglzzrBVLVaL8zV8DZOq9JQqJFPMlq0nc7aq7sc7ogmt9xSKf7nK
mHeT1E54JrHOLGIRafN6eAWgqihO9wIH62C2kmh870mldV8/zsXpCq1PethdMfoOs/qUW2CGoIVM
vz7HtI0OeOEIOgUpQWqiVxEeYDT7BwOW69dIW2EmDx5DMjziNITQpA/+41xJyQSD5PEp4klvx9J9
wHyQSiGv7AV1fbOZpSqokH0yX5X0doFkhCmeQEUi5lWBZPNo+xxSdJsmC+ZZutAtF0WoZySd7VXq
gPo1XYkrZldty3tdhSV+tVMFw0vN7PUd9d0LeBLJ7SUeaukjG85IisiMW5ksF9IUmi8ZO9wXNrC+
TqwVPkJAZqJdhayBGYgH3jSOZq3LVWn1uSsGJyt/bQ/mUmsl4H5T3H9H1n//CRFbVqVOwWbYbnHC
EeBZqkQAFOtFoDv/YKfhlu2IA4CGz5hbNtMr/CFmcuq4GCJkW7Sls1dyQdBSLf7bgOrrey+ybtne
LuDmFpk6b0VqKEW1jREQEVFZprcw4MrAVzvwLfL2qztjM9XxDoFoSMujC/eGLLQJd2Up+aHBypN9
np/d9GhRATljS/Uemx44okwOR7E0pySB/sPrIBXkcadNskHH/by3n4bxZbopK9LmBUWl7LPfxa+1
pes13FMUCqblrDOnc3+VBaZZQH2/5/zU4UfdHFuZZTRnUKw9xmLXmivpn3oTkXlV4V7aSUlXrIXE
qSl2fAGXJq7JTSgtNkjUoyM+aSIaa3rT+V5ZRpbgAYzFTvPWTvfsxYew1QDvWIh1Oll7pyvmHfn6
XbF/+qIOpxVQj3ELSHig4x4ae8qiDfiD6sPQSXIzfxXcEkA2GqyGc4mxh8O+r0ZhpmK5SHZziVp4
HanV4qX/SZbQP/9RLa9X8/QC9sjApe5DCQfNoNrkWb7LStS9lbuCf/NRD3+Yrp+RChSWH6uQitmV
4KXtdcSbwUm/q6ZuFAnvf79dtoBb0m7ubXDl/skei+RAOOENzeuZlyonwn0f+k6CFpeypZyT8Q3t
ihHSdmrB/ixuBFGoiCjRJIMUX1JuW3vNxtwhd/om6m7nX7jn5r4IMuGzmWvPGvEkma9F5JnogHUB
nUApEny8JEPeyjQw6dePyY+OHCZ/yWlRPkUN06CJma8b+2H7EANTP8m4soxnThQRxN8/CJLGwl8Z
JFNL7S3gjzngS1BrCHx8ZwvPUGMH+A6PZLqiK8CnluGb3V7XgWwHCWjAmqr3VmPNIzUXmvLYJjXO
hlgyTz7f4GUr+ca5jCjJ0Y4I8HmotpzPN3PHpeEYcefnw/MP52D9qt5i0xiAGC0b49vwSgtVzB47
eT72ftNPAzlgeNQST1cp0GFlGIGUrdl2qRZasSSBMb+z6eDuWwpr1Yih9kP9VOIVYS2ejEerITJP
wyI8Cu14gVHtYzyZ/hqPRO5AtYnq4KipmRyOP4NqZqJOy4VRiIeTk72yQozUIt7ijqNuB7Sq+hs8
JL/MfoCg6YO8sSP9WT6KkP+hJ3OeaA3vQa8E+n5Rv1s4tAYBR5eXvHeU0XKXuphBT+QIgXH2ZGfM
x4PS7zH5WK2uIgniTluV0l/7jCbqJX4SCi4hdaIVCTPyjKZqokrNr/Q8dEeqCRw+Qh0O2X3NLhMo
Aj9y78qOCoCyYgjLrZB67QUJeiVO2cZ8kHJ/XvqGjj5uMTxKX+NdKFzfA10Hl2V8cSp1C2IHdhk7
Tt9ZRsJFjMX7blOGPBrToUmzbx9OPpSy2uL4J2+xdCo2p6I1mIEsfv0kqlNTDnoOM9D28TpF4N6S
k7HzBQjDWrHFOU6FupIsOGuOj804JS9tFgYxHj1Kn0WPVorN8XMX4AKNsfUZjVpsYOpZjl5/oyuX
3GFN5DLCvZ16Q79S+ULVQFcFmLb1OVLHZtCMMEPA3YXGIQ3/Yx+V289Oe+F+lCM7DOv7FijZPHiw
q6itDyRhzc2he02poJhpPbcwG/haaUx8QMzwwsJoJuyYtFEQz3EJ+nT2yoMjgROGzTsgg82lyWKQ
DkJ3uVzjYV0mkZsEILCilEcx6KYjkcB1YwUO0R0osxc2SN4eO4cpT2brHQV+jK5MtERu5Z94k4b2
8tB/NvBHyGz7rqds6NC+Gbiw3l4579DtTa+tvm1Oomrh83p012Qj+vtpel0L0u6aZciST2jcnwba
2G1X4tuljLEYsVuw+Jav4rHuCIkG3EOXcWFpmIECtf5JKA3xgzqIrwO5kt2PxQeRWwB2moiZmWvw
Nf3bllhSScZxQw/r5hy8fFQX2NYQ3lpfrLpR+4gzEjcf5D9y4Os1in4f738I5hwyFTUBnjylQueK
6LmU6ry5zUOOdehS6YX9dz7D+fOlI9mwXLcjgb6EaFz95PsrFbxDXvmZDCl5NYMzlJ7E6Ma2UT2/
jUqVCkRPGTdSN+xWBPZoZpgN2SLk+CsMC0BsxW+EGwfnm5X7PvoJnZZgMsza4GNG58g+ywwlCWmE
UV9UafwImctrRJfLnhuDZx7M/TXvUqixxVYqo1JqRJ2WcE+nFImvUJcHKxlNJIG/ZYxyinCmQ4Qg
AFdZaZPIuA5QxVXeNu5kUq71pwXsF/sZt1wHiktsOUzszQqfdUzo58HiSROZv5VyFb8AQYy01aOE
uBrnmNv8wTQhdI5G6M12GDZRZgJ5+YSIF4sye0trukS9rJcqVKLasSc+usQUpVxrz+cHSevM70CA
YzF549GKsicqH8f+l10p8DRAsDzj+t0aJbMTpIyUA/3yjb/dTvsg/jTrXJCDS55WDUNDYpoKiP9b
Gh5gnus5SpZNx6BUvIXJUXkYUzRa8nejv+YTm90uB5Zrbb1F8Oc/Qrqnt33uDJHtbQd2wrVe2ll+
wguOrXQoBUejFi+PnH2nYWMZMLXVXKq1dy0YK38YjUlcxFnmYkGaAz7z60cENajRuPMyCyg7czjy
wW6JtSXIK87PMon6ei/rvs155hY9C5A9UuD1lsrjHUAUXduJ9MzmqXACuFXXlcU8xptCEkMcFqmD
X8vth9lPunym7hjYtdkiZI8m+hAAYrTQycMuk1EJO1QBYoTXXChiJoFzUSJJu6s2s2vH9V1E2cQ7
HX6PVAe2hlguaj5etULGR7RSOo8sEK5Y/Z0bc+t/uFUGlxjuPHUPc7qpnBPWekAoUAUWf/R/S4PZ
OTtGepYIR0aVkVH0imC8yD/hQr7aikLnE6habgBDvsl96LFpO0Nt1m+JVlVs1FAI+8xzJEH/XhSW
E2DmtRpNJWE7QUiHHhNCxyRdBo7QYCxdDQByNy/4EaInV+mgYAQ+ysn+JRf8/I9U9sol9GQt3NOC
ANGx5BGEpA3/5a5CQoZaEYz704oGfnY8+2xKPtPJZnJ41T7TPQjFDmVADtSpTTqKaLp+Kyc0C87v
v8owfc+sthYHO4cx3saK+CpALMakpbrlXX2RTv+SlcZeXDaa+wTlmHyOTVqO8eJsr+yNkLLjaqMU
tmaQFTC+seErAV8rsdFNhZRtcLYIddfrTGe8uPMaKQ7rQl1+3phqv8blz+D2AdJIYeaWrNK6wYzc
2C4GLQtXacZdAANwNks8JSMZ2fg0l9vc9iw5+kfTmREzPaQhNPsHcZcZuhXKXK2q+F3u9X/XyEWE
+lYjZfi4s9a5S9rOhcO0JLRhZge29pxbCiVcPrhaPmOhkZsvimCZtAfJ1FS107AEiUl76PeD73hA
xUyPRuxTmkvlW5diHqkDXbY//hPfGCk0+QxND6uzSp3avwrrxyQaZ1+I2E7ueWnhCE8J7bFEufGu
ZigoL+iUqEkJUFpjix5nHj+x7fZpf80SFbkgnmoDV2m2BaNxnATA0x2jiIzTLrfvlGp7isliz4Pe
wmgE2iQTCj5KIbDdmYhFWAHtXGWm0LpaRiGQiYx8UJQtHfUKUl7d2WpsjsXckTSLYwKeboBuBZLK
5tH6/3WGk2ZgUDkNqtE51Pu8oem72s6qNcbv86+MpWtW42vI3+fpeRyKyNl6EcXelykJ/grbBx4y
cloZrV1V7fqfLcoEsLXPjydNFEiuV22+e0BqprA+Z1SLvH2QQUmSkU2plticeu8Hbre08eoBZHtY
z0C4YAVidZKkR0PkaPYoQ1k5XzIJ3YO+Q0R3NojG0fDLZHz1N2J7YSril7KWehajVoF6KXsjqDcW
7lo91VyGr0gpELprTrGxUuzY8VLdPjJMyHGMgYoP/7s9yxQbhdDTeYzcpQeHszF75oi4/cLLTBx/
R/7ZqAZwgTUAuXmFBZ+7Z6cabCjV0XU/o5g/Z1I2gHr0nh9deJyefo+JoXxixk1aJVJGnkSFqh4h
aYfhL1er42QgghPCu6RzOvRP1joPYpD/TMUnw75dFWLvEbVJMcExniREGiV+4dKjokgtzHk3A1Y6
MlDmJCgyzMAjDTN0IpZwZb4/+VYtHGzMWOUmTfgtgO9JTpwNcu8kI5DuS/1CaN6jw1cddb8/42qM
ZuKJZg+uaEHDHpb7aNpeKbG6e+nh5sVUcidhZydkgwD2YxhDqv0Lmsx6AKRZ3oAesIM8AnR0FrkF
LmROlFN3u5w6zxbaMnnqhhAbi7q3qEzBJYdQ/EZtFl+YyK9drktVFoZFe1coR4q2zcaw+hjUBmoS
sC6FprVOc8qLuBx7rmUJXu9+y7Q0FHFPT4J3cTBbmz2pmGkBvh07rvu0YJ5Wgp66I9Tqki9yGWEG
AFMqCXRsS9lbCyybxNAVLeZS+r9h8rtJyF5QZ6X3ZYk7VXN8UfZtuTkg45o4K4hjfJzS+AZ23k8G
PWvGCGMpPRo/gmIwsLEWMU3xiNI59rh6mpmR0TClqQUlV6cvqIvgzPQ++60thI2YQiApyR7jcupu
MYJUQu8hbKma36gakLodtZSiTpBEVfUapXECQpbqOFRZGacwxxOcQRvYt1+arsCYEM1nnYNx4/WH
nC82gN1DeoBxxFNPTshut/JSiAXOJwV4B39rwG6U64XJ0AQxVpeWBYEh7NK/58UuGh+opRBWNK5L
a9lyuar4Z++N9u3k56qsgxwknBopSP6+KGXN0aUWwtwvzIFxm9SFccdReiZzq3y1wLGmMmzbbz/s
tBoOjYf5q7461DcCr7f/DD2EAMSAAQ3uFuSY3McaPOMOEL9XrnLH6YRfsWPpYrYxA+yRlWdIDdCn
KfMS5LD+c+QLiR36hAHsIRMQNPItyNk1pqTTaXCyFhlkHhqE3givBZq4MVldmoobwZ7EWBgVsxgf
rsatHRtKVSWj5UqvqPASesMbemXRFt3cmUQP+YyDgs2gBQEKxgHxIf4pe3jIwNrNN363MKMHit0k
C3Sx/c55bhnb33Cn2NTUOzhxmMoRATYTsLNBrNtmBByc5Hvm4JxR7d6i9Pl+UiEGzELDIfoCGqq+
Sfqxdq/NEHi9D/1BXzv/wvTf0ZvOWPwMVeu3Zs5B5aHEgVAjVUPSout25IXKf8ClGklAk1X6C650
twaTnq6clcTErf7oK7WAOyMdyEnl7GhGdPS9Ib/cWiDON2OraN9hmVJfvJb6H940A3JqrArJyZeV
bx0JQRD3io66Tmy2EjZL+dj4y5fveJH4V5d1M5QbPH0oNnOsbtqC0BXapcBg4L/8QJsrhOM68rYu
qksVNtPaZFuc2nzv6eJyvPcltNT0i2gDFCVuEQNUSIXvqfNghad300kZ/lTgDO40/2b8ZoimmdUI
MVmgujNizJPRwNEs2ovDSYMceI+zW2gTRw8KLcnNxQWlWNOmTQAhvjGGpSF8WdOEUWk+dhvAPquZ
agVE5k0yXR2I6OhsZv6NTrUvrGMTVQ2mzxahuSfs8xFCztaLA0jXi14jPOmROMk+PqqsgRS0g6qU
8/HttPHtAw4J61xBaWxS57a2bVoUGIpUocu39TqhXHacYG+QhDGZO2SeQkFisOPyqeZcRJEtKmf4
qWU3T1/wmvs8PQvEIo9KWmU1KoJWxHXXiXDDaSHK4HDZ9hAKytD+2BAV30GeOgFAEebqKukD+OTl
hxrCV6PBC4ErAauxyOUKcCXekTMpYfrXfuRaCXujdq9YoVWx2UYLUiWH1YaPeSQiXxFCLnh9Rq/u
A7t+6nbqSfZmtB+yevwNGLGxXQaeh53Pcs9MIkLLg0q1pLKJ7ydkYkxga28E1BU+p4uHPoz0sY9u
Rd0qAHICK5VPGvbVG8jh392LEzDZ3xh7BEHpveG4vnPIbRl9vxv/Y+w+hX61ilQiCf48DPE4t2Wq
2CohMQDmWh0fUuDtjXAjCNfKQ83ts126avbtuDzk/jvwwBk5zC3xwZS9rHZEtP3+XCA2BdVaT/H8
d968kZNDHfdQlAfUhVHtlulu4ENWJsWJ8DgkJvtOvEMxi7ntxeSFxyivKCzCLxgleBoR/pleqgMM
H/n8O+CZrRQS12KQcK7PHNmek95EhU35Cb8ldIdpsPYBpFiKzzX+DvUFwNPR6/kuwBEhJDYGYqHS
ny1Xsw+08Ef+V4Q+Z/yXxsB+3M4vOouHZbtSG73OceQHBpZqKOPM7h+3ow9Ax6+lQWKkJk4DX66S
YbvUj+nymnDzlU8pkHiAU3ijuMb7uP6knRtby8epbw6W4g+5akb/PIE15f8E+LVkDMouugK4wx0F
nOsLNNQN1FSqS65baU0zt0lP8LZ5Dk4gOwYoO0AWYhMR5ofdmMlsIbAR5ZC3qP/1Jb+pvsqq3UfM
9Ch0dmQSIEL1Slp18ml6pk4Iqx8HGOpLQQSylQQSaJARhWJe1zrbAhC8OBeuYXylJqOQ3AjO/bsJ
vyTED0gNPxcQiSwUgFxLn1QJHBrIB1t3B5PZN0H09k+2zMsErkYup9nxluWrdkopEaPMKbtxN1At
U3KodxJL2x0Zm7H1Al4UBcM1yRaFW5A5yr1wgGv8nT5LefkUJQy+Zq/BUWQaAfMUXaqKM6EGlDxc
dBJL8gLsv3RB2RYRgdOnM1B+OMLSOi7eA9PoqBNPdYoikqGuiF6FdhY4nLTeVz4lnOWqlrd5vy9t
nzBe+DH97iTZilZfPdWNwfGlVWsF1md2nXprpf9GUG/dJ4svTbmrAYm0CbAe7YoSNFEqhniNn8cG
nvjTaF6HyaG6Lip8kEBUpCVKQ3C+yWsvizTJ+5Mycd8NpF5hFvtBJAhL1ScGKjz2EVtEZSSBxbEV
N8UQYHB2SBPALbFjMjpI3VpvjBm50NtYFj9viiVByFxKqDV0oh2S6A2QdqE+x6qouISSs8FvtqMs
qr81Io4cGyX5rKVL95KZURg+AcC+zBJrRWcD7wXNK1RNl9WYEBXLhrao+xO1LpbTpOSgKeItp3vE
hw3kyemfqxyyFCF76cagkCpaBAzAUqHBcKS+2IDKt+kq+VBEzHNWOvm+ekTUXP+C1WQ9veo2XKxw
XHfnqMbNmtdnsLfWhoiZxROkGaAkgpA68qHr/Xr5LC2kNVU8AdiWLIiRMIfmwwCJ1an0Z0OvpyGV
G9Nnbo82Fnxnwo7esN0dMujgHk70CCbIjCxD3fxrQzPrD03xmVXJf/1fhZir8Yy7Yjwl3RnUEyrh
ldmmsakTb2z43knV2ukmEVAKP8ZYtOS4U6cVJ1/1HQj0FeyYJQiuthHhe64w9pqaZnsHEbUX7+aM
8b1DbSzuOGb8zkE1pVRHgDqQug5GajBmWKJqRlgP9XHZL4Gp+zVPsRpPiELcAaaA6XiQATaP3Fj1
hWlcdeJ4I1Uz+vKcElcZY54ZD8tYi3aH7Fmyc/mSHgIIaDb+U7E9xP+Iwgg2uA0YVcWhgUWjuauU
apDUqkpdi0OcTQXxgMBd+RFZbPkcCu2C2OUMicYMXf1I4tBycTsKuhPDFpcv1xdkIGal8j0Z6P7r
7viNZpGRKsgGhGMimFaSypVDqSN3aO06qPpSYh4vANUQjaWvZpNRJMx+i3iErutsacKx1V1pw3+9
RVqGEYx+CYCtWZ+vFHfdhaQ4a3C7xVZQaQhYvRzUXDArbwfNrtiwKcZi446iTmBoJYCWdqtmfWjK
KXP/0G4IQjhbFnJegbkKTDGGVgC/NAQYFqNPdiD32aR+xULvyz1+BpvE7Xd5SAXpUXIP4vVfIe1p
YKG7ZIGKsGhuHQPcEZNud1A+1nf8+UqmgTpmXHGfgygIS1E3wFZ0MfR7xREpXwb1+Ln4nqCmqikE
tg4o0O+920fQQIlIGy3XIYaeZTQglIQAURFVIVAITpjygrooEeQi5c89bh7m1CZsfpyC+jtFedjx
EWd+x/WIvNt4kT24f6ykrgDUOPSKBj29rneEi1g+UOGV8giJTAJLN6wHJdntj0QVijf0YWXP851e
bGn/NLC2jfGE7DNmOM1n2FDQ1k4+mM1iCL88WLIU3pAFwDJ69gEVn8LMQMoCzz7EqtLBCWplxIKD
vSLtYDpH+kbcekXtxFz7aVMo7rD/kWGo8M/Lp9KzKKOwqjhKkBIMtauKs7QppGcHR2QNt5h0K5Wx
jbbjWTSbHAapFEajwwLVeFM+U1hZB0MQGxpMg9Dr7j0cnwA8Z7YlcXvzoUPpEFASUOKVcEq1tsGP
zLo3CxpS3pcg4oI9euSQNZrnJz0UtsPlCYwTL5a4lgro0RmWBGVXvvWw7qdLgNXsYgaTy6K6hkqt
N30OHKDF2iFT22ObYZvXC5rjCdldVwAe9WxKMclNifvl7YXiI4jWWMiYl6NweZ6GvK9MCtOEOQdf
/Duz2PnqvFIstM2LGX+IAhp1tpB9RO78eLWDmt6kot5eo68Ro+SRnZVy63S/AzoPgeccV0LoTjJw
wXXbw8gtDyL5keAFDpKlLsCQs8Qms0bNrsD7r6XV/N9afVij3m6MnduxNArEzQq7b2JioRfTl/0d
6Wb7m0ua25+tgpmn9BP4vmBDgvrPWB4hdGzE0GnPRgP7/Gd6QRlkREr+9/klu6vQapSRkyZx/X1/
J8qUjw82ja+MmQCFUgJE6R4DQSTVhA3vK+Ta2YaxIAUT8MFhTAuvT4pAsDz7QOTJ94SbUQbRwxfw
aVygAHc8VhbbIEV4EgbvGeq/sQHhE7Rn1c/H9ayMRAAmdxj6ZsCPa/tQNxwUpwNr5+ycNxJ7QyX9
3D8qMCCoZrveHjrb9SbAyHm8fOKMi1F4oNSPjxQrbwRZCtzXJSJGvm5BGtn583igWL8snc0L+QmI
zFInQCn/pQf8p7dntTnJ9hnlyvCDv8fJFmRiyIpteKYujwRSdpR91PGUqr0NnvMNLUATEUzt14Qe
Pgu+xcdiR+iHby1nru0UpnPN2Gz+O/CNAVvqEOMx20/sL0QMMY/kp2QrykQQKuDqdMIfwrQe7Yqf
YCAEB2WWoic/VneZ/nVhOjS01GPY2t6dyw1uPHr+WfCp120mLB5x0VBDnX1mUzvIjobgOig+wExj
yxFMyz6sYxvs216rlqblWpRh6WqaOCxdCOiktO3LHULC2PeoeEd4BjWAAUc35UqEkJ2rtE+VD7u2
9pjYuFPIom1xec9idprkNKDSck6hhQ87gXXN9h+W9bYbmx2QwhgmfpO3LndEgwzRxU9Aho0XCbeu
tcQfmwM4+Rv038vN/stKIwNXOy7NyjpBAweWMWGFtxIHewYpUO9etelgI64Dpp/NeNCBvFlL3pIX
s2lmg78+h8AGilS0gRlpepmke4os5RyMd8L0o5ARD8RVPDlbvsliIEXxydGwZqlOafixKinmCb8n
qPXAfzv8ak7zbopqbVDrFFOVbnY8T+VeUw2hSNX5jxVYLBNJ1pkVpxBUMTP4/+mrLykrf8fa7XN9
rDR13WhyAZy8B3FTR3z0ZzvcHD68gh9a1ip9+mBQshHmwQqb8vhMZNKlO1mpyqTslJ3yMsbPyULn
l2EERGBE3h58kkVbHk/Tlqq5pHIlU73Do1ZebO8cNXfRts72ZVhC8oMXrKiwAg23Pke8aMiUX7pa
vCI8SQYsQzV/9tYifnU9r+yFhca/7YmgLALkwl3Sgh2AFcFVIKJ292RZD/fj4lL6MN6uevk+WGBy
/FFMbSkSwkYDyh9kA5KiDmXN+T5FvVAOvoAxu39p8L0+V2+UMc2kOGTq9jG9dC5P+nt1cWUsHw7Z
ufXElmI63jfETigA8ISATQeYBGAPP7uDc49PhgzqNPaTkeqJhQycANG/lgTQpSMxLRVVg4Fg2X1a
Ycv46VG8upyF++Uf1SB+3cCnxVSB+OAf6pBa066VuemEmaFMhhl2dQbYwSFzk/f6A20BWjgps8+0
zn/HmftYwhDBNN7tYzadKRBsIRvdLSGp2mLdTXPbjy7uIqmb36rpjHqzcW3yGGba4HbyoDU6UKV/
GtkPBLo7Q5yHR+ekg4OinFn9M8SpJFJLwAHjL5JbBUt6kMaWNI5cLat+sE7s6XmdlkAPZzkO5obw
UpFX1HM1i0ByXwdGsOrITzp1jHzeO9s9DYJsAFdSPTH7mZDwSXtvhH7QnqXm+0cr4+q6ysLpv+y9
vpxXyUKBChr7x1aT18H36Wx6938bCLUkU3NjioCpngBAv6eeR9qEIrBn3bNx7uaJiSmB+8isV+s/
qDeByVyl08I6AiSFv8Y9FXWHF/y0UUM9enM8piW3PeJOd8su41y7pPSWr/ee+WYnphAXY6KQsAOE
TO3T19X88Q6zAeP0z8ztPesxmJ8pEuQ3uKhhyQqmEq8kQu7S5ehbhcp42eHZ8YGT8j0WA8ssJt9o
PoBIXGELAAX2em6u8fCBjEc6z1B/ceBYhaZIKw370e2eMDM57vZ3Lq+fVUbA1sfbo2kjBlghdO39
Tn2LEtIoQ+ws8/jFl2sxfXzhW1ZuA9YIVTNpo1qDG/FcBAl1t+q72e9gvKepCHo1Pv8ddz4kGy+C
hcuYlR7hvTrsYsaFZwmGrz/yTuQ3T3k5P6pdl8O1X1KxLYF5py1hRUMBGw7t7rQy4yj/RLtB8d68
gM6EQUs1wsO21rw3oUKS/RqZNDueQWxwQHTdy/mSRZfGEjR/fI06PGvlEiSBav0xEBfISiz8pjGo
woDKfDDUFi6cp1BRpZZnRVvMPF2QC2Z+3VwPvi5u/qZJLQcIrrJAigPMoYfQHBDNTNeLA2ICpgOL
G4NMDWjM81bl8ChVdSKABihChwEmwk3+3l2BcbCBr2UC9xyX6pmau3WAD6CKN3gYJYEifUI/qyjS
YqUTwwBdlq4Ml5v84WxZ7gGwZh0wx9nvmTMqrYQnqfsZrlpYF2TiXXK8fdCf9VEpA5NVBX/PvoVr
5MTaoP9AASXe4Vr5n9GmnhxHGWk+d3N1fNvTOxe5I/cg88jiBMX8XilfV5CzK6o+rk2G4oMtVlYq
w0N05f5HqG62U9k9yBGRGlIJMrLF0BuLEfQmUtdUUH1jpmf7YfXDJjnnk9/cApHbxZITNfFhQrBd
7Bd/8jmI0hAgtI/v3ROsnmE8p2ooKYOnkZJ4kUtyl1HmB8hc7uaYxfH0CeejjpMDujh7TED7o8SB
Kwj8+kO0VHwYA/I6HRFXAipx/aAQbr8wZsB1wDn8wjjW/HRVBYybxmkTCzbBlHviHtarbOrY1BPj
PTzIn1efak/w116QJIjBSMEaEBmVLArbYNEHlwf73KihnozM67kq/pNlWQoxHjgTufIdDLtq2DSd
lLwc/Gdm1ZhDFtCLRp6OA+MHc0fNOgskNLtcmITLdgasN1/+9i9DmXcpHPwil6m/AUIpwv87qjBr
uq56+jct1OUYkXYGkyGEkdfc2x8WUOR0kqlPQkq3BQbvlmB5pKhCyxwwOsUWbZWF4aL/c2h+RjcX
t9f8F3vDzu3qYwDADn2K2+3qblWZoUluDQrFUhsVOyHsSJs3pFH5+5ASDN0eTSkw6qYaObxL67v0
qFBNVgAWgvU3wzrJC/MyHY5WKXCawFREY5O5i9cxxATT3X6lGE6sQa52rjFnT5wnVwTrhvj2ZlYp
Pu974tqjZ6S9WgGQQcyQmurSRX0htVE2cNLjr0U/jNkIJTv/JCSJm2KZdvTNKyn1KmWKtfO4Yvxf
6yeOVZ8zl8GtzDgGVls/C34l+grBmUcVmCte6rdmKsWOsRouytCeb0jc46JEuLAEJ18N8LanS3HJ
gWUwpnl0DG/a23KD2PEXG/tNpiybpbBCITrxq4FY9j48UBubu1TzksUF55kX5ufQXcGLFQ7/wC4k
y/WbmuEL69Rrgfygi7XBp9HSw0SrMoSOur6F/lNNQnHYNZDwswlScKe5/Nb5Tb9tRTdWJK7tBVUC
LDOFEDvVBafH9AUIUfcVZFr2m56qKsRAjvKY6EA3Od4uVFFy3EAQWdKDFMkUCNS/+ucQp9Hq28R/
QyrVuLsh+NiCfVBi10HduEkzWARR3CRRcPcLt0ffVSwSckUqBDnd9v30TZr4bsOFOelzkoSJJV+M
l/g2yikTW0HeQXEPxBi/wvGqS9cOnAV4iDAxXJf+TbQg+7L98DmnLndHIJlptNhjJ86hXKZmgYto
UYkvZrP+ql7XyBGb8KjuBIWwPMM3V6hfLfPagZS4SF1yyFjURQmT6d0PhAvohpzhj++zWIk5QNg8
OsqcKyfr9XX15dFPuzzb81i6zz1oUH5E7/M1kXE3D8+Zf4i4FsjczdNpZpAp48JeZzRuHD78STos
PaMjycvhwjGILxeByQxGfffGSR08EdvcWosmgXqef0yRCrpp0fvDzY4z4dopk6PF9tn33J5r+4WZ
6GTnjuclVMQz55OsUKpO2YI7uFAj3hS1nkWykdyXWDrF4qijFmotp4k9VnDuHuwaSilmsfABvthL
CRuahsHfyrYjfPjsGneCh/QXLR2nvBTKfO8p9pvnLc7wrSjDihhsSy/YE0FeFWPkvCCxQyI/ZEFl
oxMAkTea7wxdOiOM1DT5yTUQc91G8Dj+JxsGH7ddpIbbAwJXtlCmXluU9Ok0oyJ1ffRd4BdAzaep
j33ofpoXO+87PoZL+Q80pbwzxEGnT2l+xIEh7BvKpmRSvTtIuh+z3n7v1dvVLKYVvH31LMAcnwLz
rcwoG1W7QjfmdgScFWUvEsbfKOY4qtKwY8rlEKt+u74EmDpMaqIxalAf/coqSQ7D1fV+QFDkIoLZ
lG70M8FcLQUK57X7WGR25gnoTnJ7zG2kNw5tZLweI+pkHDrht07PRy8/kbXp03lC20Cra0K/XIC1
iVMTK/zsn8opzbUmHDuhzOXr+QWUdr0SOE3qvsv2zn8TNptvOE8Fw2DQR+Xzes5P5wsYbOW9d2MC
V2o5MailzI80qG2f9Evgm2O9s8MW1fR1sAWJyCCwDrLNaefEbjxWglnGLWvJaAeb58zOtPUYQw9c
iY0h/FBBdKbIKvcklNPbSo5Ap+N9+2dYX6dZW11h23hM9wUBcU8F97pXAoOhBZ7dCHnGssgWZCz2
/+vio/pMRntBW+v7gEjJWY1bYZ9Bt5pBKU1g6PSCi/YR4nHNLyWP9OsJVryfa1DfarJzHlmtfqjv
ZAqXHFPK//BerLIp/mBhsuew7CqKlPpIu1e79rz6ZT8NXw5gCZEJ1RtiDMSVyMpt0YQSO1BJdTCe
0kPOT9Rapy89MLjb6q/tQeWPqe8kKDqtPoNk9KY3DVy1X3Ak4meCtvmJzVGaWguoSJyU21rX0GTi
Y4n3+6HJO2g16ulvRGoFFlkgijYMLI7a0kr+XY70oEFHyyEqSo32Taq7d6o8hA+AExcOFJxUP65z
qByok013zCcD2RzAY+Plerf6GKNWdQ+3LB/bgcWERUg251QzCqwASR0eIXf2YWQdQbQCl1vLdeXw
o2vRRYwtexIZraOEO0poQUnqsq7qruElDgVS0XAJ/y4IHWsi7OFhgGsqc0EAAsIpImZi+PYMutZY
pTLx2CNupvUGlIhKtcjlsBf+/fd8zJ0aO7XysPPSldm+Nu+t0a6GDSlZpph8PEhy6OHx7nrDZF7k
3fz/q60tOTremYOUgannHE46XCGyqhAHjtZgggng5GinyQWFjHC6n0wQlSAnrK9EiYE2lldMQ49R
OEOBSAj9by3o0GO2hQk9fRfan3dEjX79BdZiPlDp3RHl00BuulLTgBSTLhkVCCwjp2UAAJB5P+g+
5PhFWhTn9tbUM7RhU94GdAeSvUI+qi0nH+fKEfjQKU9FPOoZO9NVkMyWkUnU3sXg6YAlgYmt02NG
kB6A+6bBiV/m+jUb7KY6dgK/K4t9fF4Pl3PJ1fs7mofg3gP/IiD7jinwGz0ZsxsCcd3zYJdKVFb7
wPN8y3orWmF7mvUbwPXlQKrJmmWh/jqnmo3CsJxdLoizzyXQiHpy8EB75LKWVLQwaW+vseDWO7Y6
uQWjic//VKED2lPBCCoZ/TccDahGbDaeqKk5dPtOw+qic74qYV2AIZ6YTsvwu+GjfT9HIgI6aPq+
iLKwIZ3MoYQWYi6yDii6taXXZZDe+FeC6P5Cyv/iFZYT7W5YhfvyCvui/zIdkZFBrCHlmKUf38AJ
GOVH4wrApnQqBQew9tpxLW9BzQydGaaNG0jKbWGKRZEPkZv2QjhzxTaAQzWr6CTBjJo6B5rQPSOn
8aYsgwYzDCZ7JcPER6cnnHP1WoXoIF5634LUjU3pIo2L7Mk9QXTdlBtZbtZS8gFN0D6paMard+dI
PdsI6ysCD6z1+se8LfM00O6eoRLevso/5oJjR6qOeHPkN6C5S0L612zYarjrbdwIRuOIdKh3Q4N1
qBW/8OLEOZmIQp3c5ZH3vG7KkoOAKkCt9N4TI28SQyyw8WdzwCnHmku2MyaUG6OpoPyI7uGbuxvl
2LE5IgoSw/g9aSQBywGxnzukh+E88elxMOJ3UrRDOkYn8KuTrClbBvRnMKip7/hReJTMAZsCiuB/
sECmb7KWCCCbmAHKVpl6ujQIjxa4k315FvjHn8h93N2yjiCMUOeIWHs7Z9bSXnGKnr+E0XVKY7Ps
VBZpgqiISdaLkK7I+n+IPHT7OVSZMbUBhsuicX2k2DKNEEYD6y/JhUZGPS6aLRplKkPxqmGp9CEG
I0TbpAVYwBNqnvDGRosoaO/Ain2V5xadWX51tlXCrE1e0iUznjWmJerCwQTWTPe/8l+EXcqmL04g
OFFMNX2s9o0P4VqVDeouDR+n4NuaDTCxffFFfpalusBnIKlLTGXt9Nx/8wQv+2GuZjVDZVrbdAFg
1LoHL/5TE6m+Yal8jWeSzmFyDkrek/UaGD7/P+HBjqR3HVShCBC7oI5N4lCnXcDzptlQm0wbqv+M
DxHCeQeEZaCWR/gNiBC8hmbFwChs6kysuPChkPrWoslbMeHW7Ec8JK/zsyRjzs8gm9s5j55av5PH
aSBTjomtPmkdacpe1BkJwrE4qDwdo4vazInyK4inXwT83PNz0XmcA6V8ybPJZsvN4zitcHz7ICot
FTL0IRrRw0cOZJlQdKLJS6CzIxKfHFtsohZlYQ5XrGVYOixTl70fojXLYxTCc2Fu+cJdzjmz/W8H
Iiuw4pqnOnvdF3QE0LXyzJyf2A6+cvcpuatnxo0C5EFfC3tgoaEOOIsOTEZcT7Z7i7tpuD71Otso
SlxeAr7yZO0XSPJwF7UWo3Nne5xQ2Q76NBY3oD5OmZA4omB2IAX9jWC06ds6tmr9tt7x8qbza6jU
jHxtR15F2GjeW4izSIcq07zTK2YyjynUwPiAwZo5NNCZcqs1GNcAoFNHXVXbOXopubZeFdhI2PqV
y8taTs9a3UV+m+6gJtTpe6XnudhjNhSDXWDII1+8KbNSa/FbPb0LKJJxS/Phu8alCMvDLl7cI6ch
QQOT1ZMwixTghJSsogwVOsC5AAv+k9BIWzy20YFZi4H8dueX8wRA5SdSKCnRNnr3EFtUuj4d/X96
kt+r3yaYCTCrAOoT8SjR1hGdbkU1iwCl83kB9EagaLulVHmz1T0GQk5UjbQ38YLA4jqSA102UNMM
yXaKGGXjl258QyL4u9R8moAQpZ1Sr+DxQl/2iHRFTePHJhpS0SCYebb/pYlLUmrOhY/0t2j89Ig3
9LlcbMkD6gw8kVaPHqVUTGIvNlU3RiBUcLYJWhqJySgu8ubp09EjoJs6FSZKXEgNpu7iChyUxrRX
T8vCX12c73UOtpifGD/K4cbI4Szb/zQYc7WzIkaRYvmk/4CTD23D2eY0170J1IhmZuVZ7tyh2si0
JohpHP9a9Po8b9otoe964PYqrKYVJhzpReIjfm4DC1c7/tC+lD++7K0t4E8C19dSCTjNPCwmtTtn
teH1dr54Fpu38mTFyV2FU+Ucswfc+s+uA6/IVIiLJM6R+dNHG0z6aMzWaDlsjhZFL/6vOomirH35
677EUv00DpFmhOBAJxdfEl0LwM0h/AflsPKWqObLelbAmqijkDXxMFoKrEErj4azOyqG8b4EKHjd
359/7OiSGJkbHPsBQqRD1Man22cne/Ie0GWrkw+P7NxCuuUFugYmPT/vZxb33JGcI1nZxt1rL8m4
ytKRyApx1OFs1cUcaiBZQrTUOK5vQNGX1FkXmJmBuCr3L8k7o3Mq701zS2yGfIhhwCfxJACAsKSO
HKz77t6S5u0Bn5FBDaYdYKPlh6v32iigJs8HfoubEm++t6l2ZHm+vQ2ZdUsZUCfjEToVmP7gpwHv
mnitp/CcXaPoUd/CzO58QgzFmBgwFIxqZt+b7fGwvBJvBVBxjHj8Hl9h3wUoY4DaisxdVWrjG27w
8k/322dfMSlEAcEgVIILE5zoMTedsNDl2PuS4C4nU+lOTTy0xtuT/YQWjozMcXziZzpFwdI4mGdi
UY6OhbKz75uGYQ30E/3UGDqUhJm3egfrLyhW1bDzpXZHMHPH8ohZrOVG+r9FrgeHGWzjkU/GKh+J
alK/u7/V0oMPs4fLGOxCQ0cOajtyMYlXlBEOEhVCnCsk7CgjII6ME5qRBjlvR8vjwge6AlahmkFj
OgSoO/37z8eTXLNWsSbJp2+JL2YHUYbkLkrhhkk0AYDjrijDpEQ54VjUUV9xlMgF1G+Yip+9GQ83
Hyv63Js0ZAXk6D3GD3kOEvr0diWqoG39w1zVer0tkntuBlJJqjQy4yuZ/2DvZRDlvejTcJUlf9kb
DMXiVk+H7j4m9QKwCzUNO8XoLn4eukQ6MGomnyXtZcBMXd2Cijr47aP2SpdUk8/fWtNvtvSxDy5b
IaCxalcmhz+Yss6zlZUfUrlx78/vbBVD/mh2Gn0EjF/m0/TBBQJjvLbP50nTRRNQQR4tsjUgorDI
XycC5WPe7BLGyf+HesACFPlHrRdp8sIRrMLV/qTI7MpNItcQjtlg8E3iJ5C+JgLadVeHPaMin2bt
OvuZ35dLCDysE7Vf+/W4yX6d1jrbRex8cwZmTCy/QyZ/4ExZ+kg50RNplmSIzNuPqPAZt/+Y/YPB
DCh4Rlbx4b80KGCbEwqozqIsk76BG5NQ8hDKm1NYT/Ss5FVb20AM2yBjQ/WRZCvgt0CgcOlyihuL
90shCpKQE/xC2dIlIXb1HW0pQb4qN8NL96bpS70NitLKg5Y8rzXa0EBLKUBOl0OgptnLrSUvCO4q
cjehl6HSeHDnsgy3x3a038XGlq7iMfRmqUvIX9K5YcRocxSrn4GCxojNCmYTGIKzs9asxcHY7Qrl
58A1+cInjXjf43ivJgQPf0dqtZYdk/67OSFtd7yYbWvsi70FdwwepG15wVP3HZM1Ms8e2G7SWilu
BndVAh7oNBl1EJZa044eWz4nf/+pgLwEHYyHMYrswSzOxpG+2EdZ2HSxA7HD6oY+g+gi2l42zLHM
sYWIf+8SKMP+TEF9w8Auy7LCiyYWZsES+3xBMb//Xq7HGk2PhLl9AmmTjvCSxb5h3Vxik+et4Bew
gZmfXraTNtzGbOUUxkELC69Tv+T6/xH35AacdyCQcjx91+WGmz09a1vEX0Hvps848CDuTPPzgmMk
hDYpdCmPMjgd+2q78tr8Qjn0W62fIxP2H1aLR6GHaeqdxWS3p1EtkLlrRwDTRB0mVZVwgr+LnLDj
QT53Hg+7OKaSLkePooRKSRDuH2Ib/q6/X+M/1rtfgzbquvqijSoG+2W94tJjuOUG8dW3zk7Kkvs/
+wVC8+ywwvmPJvushrHHg/Sr2uFuza+nwzv44EmRnS8PVdK+pKxffDwQ1Ornw0jnAry559RFnPK0
Et0RlOy5R7Q4mxytn3mjlLS8dwZ0doFeyEa7vBSyccUHnzCPusJJOrGU3GVQAtrg7Ijsa1xbxlHa
NOKbQcQVbSDtg5qAcLCi9v7huBxx6p+4mnwK/d+owpCnLNX7slsHvL1Pe9H7Gx9Uht1BMgSRrIU/
fKPU2gZt9nr+b4BgYAyQ/QhBUPuqHryD8gsU7eFmruuIwuTFBqcmqo7ingNlHMMeyLfmoAyOGETy
7chNhRn8vITpXlPyk3NxBmhNUAThvBaEETeGqkvuEO5Ey6Vmz/RJA3yehBI7uPkU/hePb4fGKybK
NRveGf4lXp3+Z6w6D+so8zWvTLQLAzorE4KlP6FNTWhlAHWdmjvIgRoiMiWMR93dDw9d43hKqklf
MnpBY6Bv/GCvypHCk9m+1+YF1NGswZnzIsbhL3AdPW2oxSJJX9J6K48+/ZXYw0zVMrcpuCW4M3zq
ZJEan/YS5Eh9U5JFAoUfnoJJ7BimMFOeNJDNRqMS2kJAjmsGXVYaTJ7I83YMUcARsYfCx2ul06Ei
gV4wYToZml3HpnzIkkIw5aRdgtHBq9b3le/JzIsa3/ewctVwBtE1CmxX5lw8VOTg01a4nOXXYzZV
oCbcOoitl5pZ25MaQHpVol5AUcRgf1NNmZs8jGRspFtLNRSI+GN+IDw5ipzmK5nUAYCB4nuvrbS5
dv4k4vBIvlUdS+4yuvQClVC/k6ugI+tVuUmiZztyZM5PFxuMrvmzxF7gPtzQZzi1ILb/ViL3BvgU
YU42FZmoQXrbmJsuSB7/q6YZzMaCQ6VYe3RBK29tu2D2J8/mPNImSWjzrxW73bdhmXY6cPKswffZ
+784fetyT41Bou0CCWfuodYTJUy5O5tU8mWKO0/8ya7yTU/LQWkxKjwP8KpYuylk/eljETqIfoVk
klStJ/YK9FqPJYQuyaf8lFI4jz0Sy/m2m21Ma3iuB9UsVfaLpfto3wABmYNljKrYjRhEUgM0c2EU
TFmbBbDBl4ghq8PiJQ3zdDqzn1j5FtqEKkT7f/uM9brp9s6tgguKAEysYHMGocThjekEfcHKYaDN
HF5HYycGWTtTd4gKVI3ZDqu2fYKyG3m0lu3e3o24nw6LTP2Exvcqbmaeah8QUwoamlAUyhV74ZUX
V27xvjQVTcTNXGQbj9VDL4t316HB4Ya5SCYoajMHVFlJRS7YnoT4uKkqhmiAFaEyd2LzNoZoPt3Y
8y3xd628ov0DyouRk/ToTM5WAY+d123uBwy2iphStr4o3VYosV8YJvycNJAm7dMOCsiENC1jUV++
s17VeoCwUOJl1VrF9x4FfRYw1TLFVK0GfwhEgWOZIEKz64tCFPSwyGTz87s73GxsnCA5cbsxK0IC
hzjx5NvSEqmcaz7UOPus+afNlozIfTVkylliX+SPqNgdJTQegRmT+5rRWLCpWrNFmt9aDwOlz3Yh
RiegERCNgqDGjwFeGuOsg3H57ZBX8I+QVN0sNfn56j4ISoipk9lMG6R+Nwhu1+wdOYm12Aq5P8go
d8URnuv51xcmsixFR5enWPbQuTeP+9UVZJPiISzpbUwMrJ5qw2gmAKJ1xqEtQf+Vap4ghQemynSx
/g+q45otOvZLE21HR8QOIJwqhGorLJsSqCxedKW6wAgq9WCL7+UKqBnscjk69L3jh1rTQ1eiGNrk
fwJJgjCHD1FjSclObg1STPtO4yxl+WuHAwFl/J3mUNk3joXc3HT2fkufAU2oiLf6T4vBdCbtR+RC
JkMq6KelssMH4FT922URlq6Bp4EEr3kU4Mfv68oSEZqW0X+ghKmBQ8G8nTPOLIwlB4McADq6Iy3F
2Fj65iOopqp90hEV8uH6g8/CXwKQeYiFZ3nxgLqfJ5Af47Ey6n0kwcmIHrbbUvDwHrELPOJ1dwlu
D+ZklJi9LwKsvlfPhG582Gwb7yNafo6xb8AF+3/S2cp5epxiAp7CDoXuEsW+0GJ0CAJHZv61e0PO
MAjWz4lK4tEztsQqOkewpVTzbrZkODbhY2/hUOdQnEOuArSHDzS2w1dOPZq3tu+Wj5Ift+MfbA3b
LuFF5eLAWSvp26Ws9JXDDLa9HbzoxhZUPEAMXjAS+SG8k7tacySa+NDYp5LJgDgzSS2sEtFleazb
W7DsEhXyLC5eQgiVrFNF9Qmc+v9aIfly8ZgWFydLTTxR10PVeR8t6R3nFMHXtdrb+LhFkr5Z0O38
ReYYAxGlM20UD9S1X5wZsjtv98giCLYGQoUjLVwx+lVH9kEZ30/ctsptSNEmJCYixxQIxuQh8X9N
KM+POh6exy/HZbMc6g4iBLpiLSyx7zWWs9v8gUllGD5oc6/jK+6ge1VmjiNSpMAQz/u233Sbdx2e
HXa2owCCwGagxJZ3Pn7Kxkaqj5BdzIXq1THEaj+mTTuybaFubuOxLvJxgWNq37uVPfiv0YqnfPEf
7jzPAIHd3BeTkbFZxCTrJeIGkPfmPclkwfPVQH+aVEpTT4V7F6kO+4ywSm7g2nnOguHTW3CTu5uo
llJpu3nkEDSjJ5nTshOa6PqI7LC0UK6PGNYOdj0wQx13uG6vByxl7rGnZIBdogaALHckrUTXjc28
ZEBlgd2rIdumMLqTO7lxaQOt5a/WWZUBF/ZWPDkUuxFnzTYJQjq2ZNisim+pDdzIqKKxUf/XyKPu
tZhZ9cHV9Rfm8uNpF3LIog2GdK/qPk7YkZqz3neu/5yQ7HJELM7xwTOddkfocAwUztcJ2aosUV7P
iaTYiRwq91lTnh/Z3nesdAOKDzB0XqWJyDxqQFy+LIgrfQFZak10NvvFDKySFpBRkyLCXfq6b4ll
1sdj9TEtCez2ooIIB0GL0tTCa7Bw4FipQf5n/QBP7if5WyNIsu7wtlBfEgPCzX7zCB/vH4F2WdEt
IrgHd9R0zRaIoaPRq2APUGHi2MaZcmeUnRpQAz3g1iJ4XOdQuRB05nsrUgdLjmOiWZutQrOMyg3V
srVqyReIA9D1rsGzN54gsEARZWy+2NJKIrdk7nGzopCIjsw3s1cERyDh1Z/Oqn4z+91rq8WZ2GMo
Ci5rf9kmOI7cqIxrOjHW0bjXoYPVerUoiccfkn5BsKYRjAPk6y3D/mDz5etaa2mzFciop1IaCby9
+cH578UOAHekInjyBhauLRKQjPSxr8YdKWKjTDjuPB8ZnlnytCuEo1A38v0t/mS28rwWg+AV//lc
gtTA+u34NDZCLPml5dQaqFpZPnwT4JYOKxcECvrPnxO/snDmOZpu5T3E4lArprff2eIXEZS6bVa/
DX6iJnRgUPqenOiY7L7b8c4ff+c7CibiM/AeIsd2K/koNBNwdclay4/htoW4VlbiucpCEBwRKdB2
9oADXJ4i5u4dQBlStBSjg2x8vtjDuLKFKYXNRxDDjb+eCcnPzI2bGszVNS1K19nQlgrYmQjdhxic
piEguucRzyMl4ucfC0YhWsx2sBwUklCz5utudkjdUS50OvxLe3nl6/WhNZz1kwNLdjMSN3U+EE7Z
Fu5s0VvV/Lu7ylakdXAXXt/lsDOxP79rlPnAxNtUewvwrmMThg7PHrg4V7oec7VvWv9AlgQCVDbT
iWyuUY5pc8ypJ2K/KiLyqNWtquuGpMehkzbAVzf96diBk7osZnF+tZI4X/3ukYGt5rFE2UUMHkts
KKWoMB3XmVzwscHRZjw6I4EcZXKxQvvMZA8k82Xw06QwSDHcsaD2okiELxo8DKQmcl9Rwa544W77
2dY7RUKvgPISPdvAEYU+cMgBohLy9ECteVbyEfJswmjNc+34w2KjGYbQMgAXYKN4HCD9PrXiAV4M
ayT+fsmLW7bqMFLEEUH0Mild4IfF65X0nkCAI/KOejx9UCA5UFRY6Rm8fVT8t6Kne4pHdWJiRJd7
qlcGFlDktYTR8uZpfYQQ4z6IkA3Cf6uGjN14iUk6/ewWhtpHiqNMDFVz6dhUV0e3GF6/S4wAHned
teQe7QVczf1FSGjp2SEBJ1ji01PXsCXbJ7nosTbLToNKnMZs6Xb7vHZEjyBjx5ycuOGo6wxi5OuA
TmDqEba0iwwGqyLjnuhHFg8wEHNcjR3MWF5KO9vm7UrTEqTlH7krhe1DY4rd6I1SlDabQ6KGjeTM
cDj2XykMhh1x0uHa95lon1zlj1M6hmur1rAs9WqR5bvE/F8/KBesapp3UDY8apwW/3wkksaefNsC
hig43uXVA4tuTxpS7mbjahVcGzwWbCa1BRJRwuz8+i8N/Bk/mUEM7IeFs//zc5CBIOhx2L8B0S+I
MvP8aG6FphnotcobhPLsSaxwZiQKEp8wC5HXnfw1gdNpC64b429e5WRbTzxjX5FwtYesYt8jsRlX
4+XfjaHTTcP3vAYFRjrEUIiv22RGsyiTv/kYO7rIAdbre5pFHMoYaSUeC6l2CgcOftQGLbS5vogD
P69Ygr88+tCdfTdzEWEsky1t6ST2jSfXKORbfeydZWwMquJkGg+zJlf6blPo3sCkKmc27SqVA26y
c6NJinSoRmQ9SIq38PDDr6UabtaYj0URclNFgV8NBGwrur7GzGe+EYUur/zZcDN/2ugfhTNRUGNw
mntrKnrLgTQseG5x9WUgXpARYfACSPAcAh35QuW9LQSV9wN76np+53XmACZeau9hoi9F5wXTZvb/
EgPuRcX/P+OrntswivY8+ANjUOkaUS6ePw9D1lpx7XJ2wSc8yCpeoK7HqFBdNryUESV8DNii0B3z
NEfzE1kF8WtMprG5r3uyxeLx4bngpc5JwYpdNNmhxZzTVArB3/2aqZm+YsfWwFa2HAO8qKrJws/x
Wm/S9lpap7Gyg98KCJSYcDMinq+WC7AIHRZOcB6wUF6Yt4WGud3cJhFcLEuZawCUfJFyRZ0dXZqz
jkn8kgJqejV67F7xApPq4BfFxoZrDofGk6sPHmbce9HHgFtjNVhd/h5ulZga/qKMmbcJft3qd8AI
ZNBPS3uN1PZc9eGhvP5XflHakk1goBz6Qm1dPXStvshXcEUnCUuaBT4lMXAndEiPxqQHCnh3Z3NE
i7/e7VsvrpkLq4Wc+BxVK3sDPfAgTs9ABAtlRS7sA6bJCb7Y/KOlQ2Swgyg7HqFRCQGko86c6MS0
zsD8P8dlzMAzcB5s5A6Ai3LW+FAJCG+Iqm+AgzM9P1oDP9mQf4EDKk92s6SR4KLCpnBh/4zZZU3J
4d8yv5CGUEk+iac2xV6bURPhlBlCP0F+/rzUK1JwW7+WzqYpl0N27VyGv2BNCBenixs/Xkll/02x
jDaNd7r3RyX8/mwtdh20zID17r/Ep4whGLCMFlDGCMB6hUJsfw2glkoDbmp07YRsDtMh9A0kfyMx
K93GU3BxYme1jZU7xVaJTRZA5ygdvoYlRd3afQ+XWQZ7j2PKLkD94Mz/53pwQesdC51fTvXJNNKF
KaaXJkgsboyCM6Gq7KBqaG4XbwBQXcfDJ7FY55eMMp5NrG6mFppCXRdtpmP1WRfjHWOiVvyx5QVC
Bx6syLRWYJO+GQR995TIkqkvtmF3d8DeZoVFtY4X4b0ZE/Zd7vGtHCOBChkHIfDbJtaZEdSHt3ox
1C0sfvKz7p2raJi72OgJjb0sA5OB3hTG0Xj2zNwP3aHl6b3p/ABdmZX8WQfUGIaJPkHWlKtmzka0
zaeGWXIkOMy9hXNUQAvSFDo7+JL/m/5s9Ce0LihJ04dgCvvb7fH0IBApVPdIKPYHGUtsOeF20tvt
UFexzj1E7JXjJ312fsebyCbA+zrov1ow1XPtdiDkucIZpfo/yYoER+CzACzIabdDE5YyqcZJhNmc
nnQExFlZ0Z6d9zUPynePcXJeBU8Xq3hpJ/Ukpp/qs6D7+H+Ds/HKjaZOBvKlRt0T+X4ULHriS3uT
Q6WgVHM6trSeHgbEBuYUAXuA32pLcydP77/ibxxxr/4z/NvYqwcZd5A++50VyLYWchcR0n2C2DAQ
8wd1nU9wsJPSucJCobAqoSUClARO6EanDNVAH5H/SSTY9jEGprssf/vWIRD2PUgOZlKW61e5AT5J
UFHdW4zj3u5/fdY1rP+aoNOhk3fo42pBrkC/8uedO6bPlNiqcbwMPG7pgYyN7f0XQ2y/zF2/pBUC
eej/a21wc1xn0YOYcbhM9o04UGm4LoEF0/BBJwoTg2ts+lGqyqQeWkxjI6Qw/SOUYajmuSdmJg5h
uZYC+UUzlup2cyLcMLQmcXRS3UEmeXpqC+6DdJeH79qGEOVcUuoy0SlS3gr7SIf7pNOiDMupFr2i
xCjDo3XgqL0/CAX3TYMdEeXqxngvYeI+fel6MboOPdjpHdE7zEM+9ALW5PzR3Rv4Qqxn+WEWZWMz
SrtqLX04mQeqrpQ/sxA5Y+jcCH9gcU8ykC4YbLr+Yroys9MB5lsi4NCJUPWASYiPLUHtjshKBJN6
Qb4c+BDctcOmTfX0lS1dxr6I2HTIPftwzY74e/nmrvuwHUyNps8o+klvo3bwFgd17iW9N3wP0D8P
puJO85f3v9O8TUazOoRMMcgBwvPrYUxP7kVOmvRS5z2nFWDC6zvdWTFFpMhyqDXa74lcT1GpSkqH
JWr3FZo2jYH7aumvBZtsZ1l6DEwp5w6p7hPc3RxlLBeTA6nZhBAGrfzk7/ci9t+A79Ehe2EjEbZk
wlIe9QshglqZBGtjNCcS5ZTOnCXn2NDKyALUFOAiFFwDtj+c1z7VRkKVy5mK0bpi+1z8e4de49wd
1vv6TvPw/tac0v+5NThnMaadEYSLGlB+XUZ6aS39T7kpnvzL9yXY71dhP3GyVG82Wt85cWD1ILPk
/gtIJAtZ92i96sQeTLQp60hmXtuLTpxnZk4aMK7C/Hu7GBHHzqWDM/S+qyo3dXhycf1ZpL5RSH8u
x/yYUA5RlLTMICrbCfnslNK7a3B9l1S3FVfSWUlRrgeHCUFKnFiO7C8NiSE4xFqvijSZu8q7cPnP
u98N15QW/dbmKxX1sBAwWGjhSurWDPG9IZmQEN5QS2locBoHAmLsOqJ2YV0EDgeXu9pgeZ+Ip36T
iReVitYsfuDxJ87ML1lEtNr7hVrDWjlmig407T/LZt873OOsyCpyBMsE+5G2edKMkXDyvPathx0/
9JGlX1JpPOorNqvF8Zj/GmEzxFgrVraJ9nsD/Pv2iarWUrxo5beDodjplfUVHZ/ZcH8X7nF8VKsR
ADrJPucnBYNRALpN/CxDEgJzZCeO3YNoRYGbbLoNnd909Edp9Iyl0BFliD0KZFGjT+6vaB03S8y9
pL6mjFS7Y7vWfDf/5mjsTKsP1LoGMzo/DiCC2J1Kttqhf6rH+WxpPb5EHC6QJUgl3d814vRc9LA1
tdx7vbAv7phLA4LY+BoP3HlRPDG8eGtZ+bN6PcGxSIx9zyzVmab7jhTr2PjzxRmggFE+fJK/CCMG
x5b3P0xvsjV0cdMGpeqbWLX34L8NEf92TJ8aFflL5pXT9SixVoz0IqY5evDZFCWBxh1YHHs+eCJ+
2F8KxC+CeZHPqhUuKbSgjf3kIGngmOxbsfQHXdmzYpoaWXQyDdZj9flyxUhnJZSPP0DxQcjGM0XI
JyjdvGib58shejGddRGPEaCB2FlOflJHOnbvigzjrc1RQ5g2kvfxxyf5MwZi6UUINUKyqTLnVp8G
XYoGPLYQwCStDNEHdCzBUzZJd2aypKX5kw+5+roBPmDM5bdrsaDdL/73228fROWq908Ti7ffusVK
swYhJmlc96qtqreezMhe+h60bmrow68HlAo5ITDUGUf80tfYPiyFBkfewithiQM5jZGHCITrwV2p
tP9dptNRSA8Ntp1zQXQ1Amjep9A8apXbnW44zDLF4XoKJ9eSdjNHyX+Hu9ZBmxox4qgIm+Rr84PC
t3O9pmHe4ugQ510UvcxeBhTFogmbhsdb6KsjZoWY2BKySE6JlQ2ZqEsVsV/Qm13hQ2YmMzvTdlfi
dzVvOUAEgkcEqyjYPE4aupckOt2/8jQ5KScfgvuOgYHEa31OXd+XdKg+2ERSiSqnLPSZH9eIdMik
DtTEIysKo8vhWwN34JcGO3HXVSQsddLmaXfbAzS3Wo3cmc1QuzU0h+gRcM6wKyFkiyg3UsYOExl+
qfMK5SrsF9AQZ8Gy9UZdbWbKv3Up0W7ZcZcfWrF69ye6ecgt2floxBB2f6dvEf2w2XCpgly2NUCy
Tmz5nL8e7I9Az+F025lHlFGv36NaO48dmPxHfXShTceO6zDb4N6DhpJCa4jIMV0FHghai4WAvpeN
hJjnOPlAU3bqWkSYu4O99JwfjL+BgA535QtUbMMBwkbOhx/RAnsIKO45oQPK286DcejlRBK6aRtI
wRk0p5t0BnYSMJQPPKY/owOTbXhl7l1Yiu96zvGnPJhItzXZDBQ1O18x605UF0ERiHZgAB2j0+E2
ZFpj7T7ME1MZMgKYkddgBk6AKGT9ddTnlBvNXfajPRTtDdO8flNlLHq9O/fZXa7sS+QeFwaPAiE0
Zcatb+ICs9CgAPM+98yjQZnXkuue4fGnTIQ+FM2K36GziFRo/MMgIgNRwVDyEtNTG7JGB0WzO7uE
1cY4t/M0UhaWZMW+Zwp8uueHaXggQsQ42itkymKVON7yVasoyr8oVzJ3Y8U79p//usNtnKAuZpAp
uwzSre+NpBP19DRL9syiKni1yptV1L1VtTSJFV7FeEzx8N4fde/rcwW0PZizW2KASNNmqvLHOXwL
C9UEXp43vV0+4DW6CCSgmYIoaqO42Cxps1SfBdfVDeKGIqEVgsXTMO3taU4f6Xe3kqqNRpKycGwp
Ctzo3AlR/cl54xHoktLvT3wJMxva7Fn7pgGN8TSLAZxtOAjd01sJutrTzRwRjBErKFmm9VCNRs0y
ouANxFMlUru9QlyvnbDYHmxMyEJ3KMGKVoi5OjnOWw5H8pM4N50+2igmyRftvESmQT70wqMY4WJo
kKnY2I/I15+UudnHpaQmmDhZ9aA5VLMNHf89iubI/+fHI9F35XRo98SjT2vla1te5VDCX5srqz5D
Uji5EQq7SoXEZzUFyURL5SN/P59dAJEi4r6SvkC16NLP6NxAf7P0zq8wQ2irV156VlpPr0yGkK/N
9ThGch3sqvfUJHQcL+YDjJNLynk0Q88FEPahDRduvRyciL3LpXOFuYUpajStqV5OH+0id48Bjr/P
qZs/fyMg5LGfza2AY7vGIc1U/oYyQuEM9Lq/DB9npZwf5FFK7lP9Tp2nYgWqvaJK1ReZLSgzZHIg
Prim49IlRwXuaDqfOnFFMoImeZtm+cuc7Rf99CvOivKUJvfTCUrRwWtjCKOpQ1HckI6XYDqDqea3
RO7uPveX4RHChfsTKQY+e2xxk5KTXG12AKN3SFxvzvcRFtYfE4hk672zRlLf+EA8SMfFV8Rw3Nv+
gtsOPMqo6yvTjfFYyod52WXrFC/YANwNEEV96wCvbKoMeDcrL57m4sRRuAqLj2xffUDm09MD/uBj
TcEBf/wWQwHgplbrRsBFO9GlwIkVFS4cDg72Ao7ETBuA+2FCMs7RiGbAp+5navNaUEegou94XkVT
lFo06dA+aV/IgrywXNofTqO0YxZORU05GRX6oJWEP2SpNhPL0cYULVWLM2Xm1MWmz6fivir2Cach
c+Vt8lK6YXGZCzh9nEHUXy/bm2FED7a4TrH27oZc4vNSIMJRWOibYrBtdnpvXamwk46Y9MVGzaqW
M+MCEWjHck6blD4/pqVItpezjrWrY0wt5OaYTXMfvGQWRnUY2Gr7HZ53Jkau7jiATa/sHvqAjho1
L8MAUnEcgfaKp2YrhQF49lVBUAIl1XI8anINd8avazDMTW74xvAt5m8VwwagqX6OWk+Oxm+Em6w/
JXfdEJFW+fls4ZdX73Z+TX8y7z37b9sPSYWHJ8XhTUVoSfxSR7nWCWMjIgD0WYrLfZYEULctKr6l
odgduO5ly7NqkkuJcOG9TzQ/JqTMzgBY0KeOfnMKxWNMhGu4Y4BiNSN+toKpoyMWePyu1SXzVTRs
YLFTDVM4Jkuregul3YR+8/bi8l7U9vq7SX/hjQnmt+0HhlVBPSrSDl0AiNyI2QcrX7CewEMCTiwc
R9RaVjmGNsmlbqftBrh9+Cy/kNClPpoabjcTMUGgq0cHXBooQxwJFS/z/SFFNnMTeSge4cKJGClE
WzieOnmallRhB1SHFnYi9cHth5L5kAI8Kdu1t3i5Q2Krz5M+EDlTPi1UzGBvsIs5GyUbWRmhTiQX
Q7m4IfR2jCj48s0fgn46LPm5R42XMzooptdDr4Xw1i76moruAqoq4d3ryYkOCk1TUu4n5+qtONQk
Oo0FWl2Ky/0ddYymUFvF4kZhiw0h35tmmIIQctNJ4X0iaOaX3wPRdJrYuZloI/Ee5FjbShUges+w
JabY8q2yEJE3b9ZhFe/S8fF6iWhKNGUyQqS9z46HRtOKOyvp6iZllgiCUD1U7CvQYBL94/gAr6gr
umCpf6fDwt85MFPI7brZKNbCe9Y9Gd438ZxDcka4AwCeuCE/w7M7yN3l5e4c7afV7mPwh818hojZ
ovE3UcULBaLyWds5r+LsljpxqMDkxXE39FMzRLh2VLF3zgV/cnBL292t+6bwcOq2FxzPd7Abqya9
sbAJHW73/GJsEPoefsBEQHI6GESD0kf2KjhQh1QFsdrGstpsVR6bej57CaHEC+eRkh0oQb+0L6wH
LkqDSckDXFbKNet/kOA9K62yh+ha+eymyM36u5DTzCEF9c/LTsN20lNG6pIZC3m5lR7ZYMjX6G7v
taUhzW2UJmcG4jDHqPc8aMm1mgIhXq/N4u7y3M7/eksxpOMYWHanPY+RsVJHAPEDusBFxBObbRdg
ljTb/YI0oCGK2DP0NImHmShY/DdcbKujQ0wrRJyErPrZv1wMs6m8EtTdrP+sj389Hl7SojKl7WPV
ZNGixxVsnETEFVsXl39TzWg+bEMFh8nO8DHWlKiv2hgE8At2vVxF/iemj6O1LjXDLmFgMH2fVztW
7Qhh/IhEgCfxXYtcf/9tHkQsEHcThutbSPUPecG/8go6z/RVYHgUnZrTGuyRxFyZsPJqaJ/bMYcM
wCICDNNp4l1kzHuE/D1PCJbQMpROj8ACaNjeDRgzXkOiGA3yqItxDk6eKv2pI8xYAnHvT7Cfhk94
fVa7u8Ma2z/UcYkSg32xhizu9vA9y0ksEpzqZaTudiwaZNtGJIeqmVPf8xkPoOWd5zUkA4XN/yEn
zCeqagJ22a+SVoQZGBZj1KbaUJ+zWuPBrMQDb4SsZtyhCIas3aE6ATm0PN9JkbsC5eSPj1lgOMxt
NDvqC3tcoHhtPkFZaL6nZweiAisDDsQjwXkwDAEoYiRyZXO3760JXUG6RbXso9ykBnm2a9chCtMl
2MYvv97+x0W89kZjyBrSyPVeQE7aoHTMZnly7OiU0WYfcCXlZ1RkYFfGZ5mMlnMdYIpknVp6/oy/
6Hc/LNNtKFPFfLXpyr/KenKdHMIyKfLcekc/5o1E3hE/l9CHhh8hGLNuszad9Mi3Df9oRHtqtm9i
xnMzusGs7sPgbQNyPWu0LIQwjisW8KohfgWXlNaLOIL32jJEI1AFuRu6r15+QxioRDL3KBVeIZrG
4kgzCRkjW0qieipglgTE2d4dWhGojKbTGXcaVMIKFu4QuVeXjet3m44tAegoLXfBusHug/2kIfqH
74/Snzu5Ol8SpI2seawuLlALsJxJ7mzWkCfRMYFd723Ca4CZtmnlBW4ET1nF8STKuzk/z4NFycAz
uDUT6q0bEgeDGWeytM4m6hu0mTsTbEVTKUdHlELlCTfFpFannYCSqf/utzV4b37eIJQobCrZHpsp
IQwlUbEq8vWjqPcsqVSYrwBHTtVgxT+rLsclzkV8jY1XpX+eiIvK6+bZw2S7bjZEJmfapoU9yGs/
S56/IRktpwtHnhQr75kPTLwYWPTAUppx+PjmsCy5tZEbETfWXe/OxtXwrQXzih5zbqjkOtSS5VAK
FcUafU5h3fKymnfQL2pn4tSXkximu+YOCn/i5o70v+OVJOsJrqLT4DHjmvQRAA70YLNmiXOMhYtI
NX+I03o5Wk4lIS1lobDeLWYpb6SATkh4lUWWZSe1eojUNef2Vm5AmJK9isPVfvF3LIFVT+9XrNAn
rGrybSv2PI9HIz79Te2i15J2kt9mOP8fHRzh1tOGHW6V5mmpT45mbr9wLPeISdPcx7dsFoLhEEuh
mCYcjZrccGku/QvV2SBbKxB04ZdwIfnU8FMkSEluXcbRVTWuXlFdCfwHuIN+kM8ymxEZCs0xJfWv
E05mTsr+P1ca8yTU4Ka+CIws0wnQWKosoUOumsBfh6E6hnqQrhxA3Z/GEexgLjQnHOoaeMCPz9Q+
SUeGf+QBQwL4a4QoLbvsEb8g+/qACNjtFSw16PZcFG6WuzH97Xv/fN65K8E1yGrxXQu6ViDFnWi5
ecRV54EnRWtKGC8QUyCUrWF3m+dh0Ji1v1dyMFy3RkSiyZD/bDvr/5MAZpM3eBrsyHgwN3GQoJQv
vxkfAgYK4V2lVzmK62b+3+A3ITWfegfgrXOCQUbZSMrg17V0ZHTyMSyxKymN88aJFRSf9IJ6X6qB
di5SxMwmXnwLw7QoPfYIdc5Nv7IraWdPQjCBd1DJPsCwbFPluB527EmjUPo2jPBhE9egltuUWEID
VBOrXFckzp6s2HhFPPTT8zsbj5ZL2a2LLD3ectF7IKdF5BlqDM2Z5wLI0lvUnnL/shF1dzBJEbGS
oV9ORnkfRFs+SSzD25X70KdtaEglT84tEQSKpyeIxTCjsgSlkwBphY6FLfiwNqFXhFJ8lA2cL2Xd
DwjNP03Xv7RP8unKf2CiKIa32hdeBb2UhDy9WJj+adtn6tzY44INpRwTTprG7yX3mscBv+2E/R8g
yNnRBXPu3m2SNA9RC+2ZAvRfYk/ZzF0Fyziv45SmhKArUrCtQqibA0cDVQYt5ZXdxbgXlVi0XclZ
ZuUGm+YPp+FxVBUIOh0IRKPeBGLBHPurhcuMF1DG8OA3FfhVch/+e4AByAc5snJoa+Hgw0/gFeT6
BhyWl4xTnkYKWYzFJO9fPIHI5o2JM4q3xpkx+eF90oSVuKKEJsX6pM//qxyPkVeXqVbkhzrfZqOk
jCmNcAPudKiswr1msMurv38qWISuwxFIKOJsXmwnZAX4mF2Ypf2YeJHX7AMMuHEp/Re2cqM2tRPi
r3ykETl7JImdMs51zaasKnhAhYz6/neTqCF+YtdnjgILDPd45D6Lv2mNY6j3B5k69jcqCvsCKSBs
lBL3qNhtpLlMrSUxw2nRGxrRgDBDsbip+UUr8xSt5IXuThKgOVRyQ5rw9jhJCJRjN5fZvzaAxTPc
jUUuUYbqLfTiSIYoM+eogEyzF+p9g0T1Ex9Ap+t95SkggFxlv096mJ5yF2sY7G3DK19xxMMuOwEU
wnAo+deDLCspNKSzFkWIjKW51mbcs6fDHU5Rs0csHgvWdsxsOfF7+8x4P7LepbV7gRKcZSNOy39s
gHrEphTDDOTVTz0G/AthDHjkfejff5oXyNnXFIzHDd9jKzY1W8zkAsQtyPagotc9jd6vlfCKeJzi
tw2Xe+ETru58g5+Kby40QvjQgBA3P6AtUJNgbja0vCYGx17dEwsdXLA0xqrPZtIiRt1SR84SaSbs
DS3XMg9vEOp3kZ+Sbf5msiEuAOfFT+i5yi+ITiLTefF97ClzbeWnQs7vwRlVEc+GbvOgvUEJ0tqy
H286hfaPYEJE97oKyY3VVksLmY8xxJaLbxLeSK0qZKo+hKJMnNZQMFyyxGFD7QKcbq1O1UrhT6SY
HOjznFA1Fe5KzPPA4G98uQMA+PKEsYOUW781CI9Z60DnSHqMy+QIPkpI8klUKyo4keguBN8pwH/A
SBzdJQU4t36LHhu+uVtVyv+qUk0vO2A1E/mAKI4FatPhzo5ZjWHzyJ1Xm0PG8wRRTf6TwUowh6vo
wPDT/c/I21ukrbp03L3Jf2PFoRw6V8ybV0gheQ6/EmoAVxQOpmtiXorJDiyGjCd6zuL+U10FUwIQ
zISmiedh3Q/j+jMpepvfWyoR73MYeRXJPbJW5QkMaWBDJy9VRcOq9fMhQcQv9CrL/z/j9sJrU0FH
4ZhKRNxuM3zr4Vtxq+nXPI21hkjw+T1y9vDqv+U/oZyhMzl/iR3KtoeTm5H32DoiqdyapccYqi04
WPnuriFKScZ71wwBerOAjwihTTt+8T+S1mK96Qx78KvdYn73ykkVM8cgIRQNC8iQEmK3wumMuroV
fzTUsXi5Kf+Kve02RLs/BRY2vY46XI+a+CwLVAkhDFofl/glNbXWDlPu0jrshgm0uxqVuieAmUVE
Iu7QomUf9OLWg7Q84D+giB1he4ko4dSaVSeM5ztdvBEejxc4NGb375tYQ4W34gqUHe0a4zAgXIFN
/6S3JMTDmwbn7xI+L4Thn+cOYlE3brBeON3dY8+UOW2H/cy7iNOdkyf7AxeEulA/fWSgqrqpmrHi
yzaG3Ry1c/o/vs31QhU2TyNk6GqYFv2aNHr9tJB5p2bQeigMDgr1Ss2jHrVGUSA++87U1EpkKbCm
KWx+wxLyChLS1GdXubCsJBKDWkWGCbztY00nEoJnBQDOVAG4BMCAxvs0U6dbCqgxnGivZfpKUFm6
Tl4iLkhcek3JPtbbutk2flmk+O46cY2ovlVFbeMbqK45NU0duvA9nfHrMSUamicGD+HcpYchlqTP
4RMVvZ6D7X8h3oWW+Qm87FX/zEa21Vr6wgU4w+sITLkn44F2wAw9mMwjyHA0nXkWD0wXNNxcrjnL
AFCp9u52AkhUJpWEzIFDPcHBvtzRikf2L762IaK1Ne2LG9VBeujUe/UVcjrG8xgkl+Knbi/Gwp3w
zdUSG+U5bd4y9Cwsj8v4Aqe8ZpoGQK9ufWiiD+I7KGGqP7RJsgQTbnr251S0yw7YrtxXhXl7SC/a
KBnD6buKmP4P9MTEfieIeQN/UUP5KHlDT6zVXa9BID7iPPYW+wemnvQQxvx+qBdTlYqBvWFI47PI
nQZXNGbxJR8LMdSAUp4wciXEOUtMXfZ1FfwxmIVKcK1sTzA5dW+BAcTaq7bpodhdxwZuvclMRFZT
pI4paLu09JhGz+NtZPVHiNTUkqJbHkjp2o/BFJ7a4R7yrzv195Np+np255r11cbig/yQYbdLLyVw
GjgBOc7JCU3viOBdR+h0F/miszJ9SyfK2S2BPVmx385V0JgKxgyNB/VZb+b/tawmqTGMTiXsoWPd
NmfdjFMBgKAIKVqboY3HlfV5m9QPdv/VNUvFhRY66PQKQP1V68qFJNA5hxjdAYEpEgBknNlQm8vQ
mGXZ2W6jfMCyEM4pXw1Sk6udqhN/vRrpQBO1pNxUji+M4LiensZkJiRolTGvvG0S5MjRGIncTxfU
Ql2PtDvUBnkRnShAS3K54CiDaZs85FhkV8GRHbynYffTpUjJ2UCzBXrZbkMOVVbWlR+KzrWyirG6
a6Ga77HBPkc2DMuZlfIR1Vqud5qfl2qXEIx3dai0hYkYeDgJVvas0GJFrzM9V+Z72zEwLDhV3mdv
8xW1dIFjzl2NPYcuPBq3sDqr/cz2OgqMx1XuyKTm6IhYiTZ3HlBVIm86MJ/VSd0L3z3WK4TbpFkt
YvEPd79qcd6R6FJUIBm/YxJd8DzoJPngkYjoDKP+VZkXdatmGfy6UZwJ8gTIMVQrdXIVONoNvizF
RLzDnPKMX/6zVpcrcOUhU1W1dDvhqHhk+19/UrIk0f6LRSlIDPaZtYZFmrT56jzjLSbeX/+xRQ/r
N2kADCsKHRyfkrxuRqNKVEjYIjLpmXAEHZDpxUs16WdIjQXhcuuGUhBQbSylYsCy6liOT716JY6e
f2DI6RhCssE6waFoLii94XZZIYRxpKMZHpPsFvTdBDnaYxwr52lRVkAeHlser0A7NE81+CTG9Ir1
6AZcITo/JAuvur9xdCchMe7deZyGV+oKjpMMaYdC0ctAWTRTJ0eZtVrMZyPMO/cgPxkbfIXi26Se
hx0cY2Di8PBBq4CRNEKOTW3ShdyTMA+OZnTvafhQ67R83vLh/Is5OCEr8gBFSayIbHLwZLhqfX+K
ulQt2Muc2kG6naUjMnADJjz/CRJeeh2Txlln/qC3/Lzp5mJ3wOJ1puNfwCNHUEYVVwVUTsnp4l+r
D0htFDGT+ddiTYd8RYSFDfJROBZyv7l9dTxLAghuT0JEwZ/th9/K44zOwoRj/S7jQJf+T1Oxb3Pb
xDhsMUx3TMEzseG1OrcsAQVxEKoa4zCRo/4M+5nRFlhwzJmzVm2k66vJyNeAVAdOO2Z+thtFcVo7
idELdL/H+DNFPwuTE7Cf+nGi2VqdCZs6JTqB/qvUNUZLEzGtuFJ69Q44HHblfLCiuIEu4J8Y39pi
2i8vEBr6rvBLbfpjQr2NCKSNc7/ma3ClC7s22GO3OesrccvvU3jo5G3eNpMN9EuhR2Dybcy92Ack
k2w+qZ/gK1XwJdLuoxOb82SRENPGCVdyJXm8reZH8ycRzLe0ca46HZ8JWO2Qyzc/pS8GYd1Lm4Jc
O7qdj9yZQMrCOkRQXbA8wZw25urJS6tnNxiSLBk6pBu3/YR8X9i5o4YqByAzLWUdn9fmiRe83ROq
clVVQdK6+qV9QVyTY+tvkXXkeeXrNZefU62ewE/A7VjBzXtr8tqaiPWBqw1uvS/BffbgrhsrK1M4
lgRyWn1QIJ7bc0zynOKMiY+DCt0pTzqmEHLj69IbMVEi0D2Hk9nSfDa7qXJPvSzzrH1UlnBRGlrE
sqy9W9okMViuowHmAIJuvY5DAObY01Jkoa+3AKXntmYNI00Q4uCbfP0Km/PqSdDFStZXDePhSVo9
Uo9NoTAE/psuz/WOWWpqXSFaN1DoPhcm7SSHN0B/Gloh5fGft6M0d0pJ+VZvDRD2LZh15ZelY/8P
WvYdFI4S3Qsv7i5o6qSmS5zJRTZLNGRYEL/FE9HVTjPaECoSMTqPyt1CEi64Ag1DPtsZ0K/uB4tn
90B7U54AWt5+dWZH0c2NvEKJyaTAOUkaM0fssb6tQYQVtKC2U4Cczn6o2ilaSthbb7VLL1iFt/wo
+9SNGZ/9ZeZpO8xLeyGxIQwMj80ccdhHIMTZlAm0oMgJGzR4cZ+hveJRrz0l/XKugwF9QtFZxykC
qJZNlBEnYcszlWYDrYwezMl92ih2u69PeGfxGAiq28hYWX37iyy6yIS0sT0GSU5a/797aMnuCpOK
Nw/v24+Zk/w3/7sum1GeLxWQEgUMH7YgzeRu8JPdstfXtzahcnVYqCvYnFUM8yN3Pki0v5KaF8a/
kMDNlo0p5W1XCE8z7tsXztSNCKvkF7qWsdRHWy1j1JkMefokixiT1TSqp2d3w4FlpKHWfmAW4HhA
BeqxWfRgfQN4RR0wTgDAsHfPPmcuYCttW29lswOtyANnrw2QAqKzciI2IXlx7n4Y7mwxIzwRSlaw
p0LVMHuVC7T/mdf9VNOdY/fhA6EM+vxU4AGpv/SBCDhHSuQN9YYY+zUGGcAjPQEoPlWwtEHnKKkY
6b3iLplgzpoE9nPI7MJXwrL2J4gpYVNQiFoUHl1qhl32WXET8a5nvzZ8cuhlN0fy2za6zS8AFsL6
cC4i72lfkZuQZpp+FT3jh1kdyofsLeuTUwgWtHFK69vfGTja1sgBbSzpiWC1UUetgoJ6z8rUzxW/
OPcbwidPNcmN9WUzBeEHNOUGF75rm7s2M4cPbgm0v/PxwaWKp1Qkf0LdtSsxlI1p5Or/zayeVMrS
c/pcArYxOjpP/DZ6wzIS0psrbMTr7q7MCIgL8rEuAd5oR5Vkf4IXU2gUn+/1hnw/rpSWK1DSD0ok
7gOzSZVbFVXmsxLkOT3efXRJ++XHUQ/sbV14T1pp9iJqZI6FCdAHZr1FstCVIlOnZz89TGtkFj1b
hBFq45dNfPJqXNI31JDOFV6NAN5OfmXemba9e9sP0g40YCfLLUm5QLmmF8/3YoKn58aunwyvU8Fz
7dcr+B1Kkc9Eyd7Y6IkIYPD9cJFyytG2QmC34GLw0MMehcGx/JqUhFcvM+wRVGR0fHxINMj353Hf
dIc623U2sRyjHmktRR388hy8DZa5A4JMwE3Nkbo6jsmDTmQ/F4+lteCrRGkh0F/HDwJMY5yDKxbC
9z8/EuJLDoNFpJ8g4Y7z6AGtIDqtq3/NwmdH6DN2dMsudy6tK+cOrRyQmP9jOr3gPjL31fJzP9rI
pRh8vgxedOQqbLuqyxLFAHBaS+PXYVKVeOo3IM+fHHmxJBiPAf1HKBSBxMrigKyzuvW9O9OgFoxt
kGXarP5v45A5VMN61LQ9HOUVYW2Yl4J/2U0lVel+EY9m5Q5mDtiFe2XK0FNISiL6atyVjh3IaeH1
ZMmpBN/SwIb0r8n6LhOPVvvKRAk7uamUIFdFpxoYJOiMGzJa7FN7HXgprAK5Th9peUGxMygt0jD1
Kn56bS9lRnSlnm/vwqDxcagd8RP8tn1T36jghr/4pu0k3e7mSUIM9svJECrOjfy5J7EvcfWid5uq
RZ6lZd8e3ZS62uJxqAZk9jndOJqu8KCkv3ejlcrCQTY318uMjuxsiTq/HOLCYlTk2IIcUHXyb9A7
G9owDZlukt3JZRRMZgkEcGNw8l+9CchVHXSZA2r173fjP657Up9MFe0hHG3TMNm5MoQDVXbJa3Vj
dzIEbaOXS3gsp7JvAPgjoKXYiC0HE8Tw/1+AMxtyRchiCvW7zDAKm9KRz1XlRBZrFnUymTLqHaCx
Eaf4JHK/UreM6TsBAq1xT1EOVYSlrpr1ya5yFtGqrcPf9khV3BF5+6V2LWk/dk+afbCB3dPz0JNS
y6b18v137f6ckSuNcPZ375x72YKfy4jV/yMMGsQIBYHGWMYQ+pdTj/weXZA3yKN8a73XxdrdruCV
yW6+zJQLzvwFawW50jRBWwwAjtnkRJLWzOFOBbSn6ePYmOks2sMx3Qe4KoGkzHayJtZyVLaDP3Rj
izrUEi1yOcWJxqN4YSA88gcMhb1XFAD+/SOyK5xlQjnRRfADdlez1vmPhgfyHBjOSOL+V8a5YoPF
P43Hv9xHQbEqB/prtcCE7Bi0vPL2sSnx0HAH1PMqDFRi3Ey7HXOhvNSDI9ASJyeVithtA7CTfWfN
XuTRTMxmha2z8DqZqYgfSVlJ6RpNNI4WW7jaxIf89Z+lnrMJWBnLab7c2chLEwvCjzmjy4+e2jVf
fpONLUAqrQ4KhRB40dAE9lpzk5Q+CGH1QIP9gaQ8hPjCFBUvy02DHZLjY/KeXZuSip6Juo4ISkIO
X3y5xY+2tFiC5tUNEIO10f4uYNgvD/Zc2KYd7IAna4DD1sG9lVLI1dnIoxUa7hRq+UTdCusTNR/W
fa/ZmdaQjbaNlvpLsQc9HG1AR3Er9l1Ony7MLrg441LiL+owtMAHkiLb2WfLFmRoWnuFeA+OtpGb
egK+Qo1b6mS3JYkl6lKs8gIXfiHQNt1uQypl1j3XnuewiWpFgc6oDL4NMhXI6CLe2mWBOfQ3hzlz
URD0tTX6jltkyoEY6w9z6tRbU3K6HRC1+FHlnHTPC5B8+MlFgNSlyUmZiEA3dssTe+1SHJXvXHiH
q+Y6Kxa9mC7x9Uqs8+vcP07Gu7u8+c2UOkBdor7bR21o/MD2YlPGmwy2f6N3w6m67mFJhXxaoqwd
/M+BhvVfE+8VQXY34kuxEVrbJGbSVPAIQw6dXenA6b2UAJIJ5KLJWTQ9EJQGbXlmoH8BySrSn3MM
rFWWyd44bOaMXx0c/CQ3Bifz/Cr2aSZPgJapR70m7qjepgRkQDjHUI9xzE9VmaW9wIxbobk/GHp5
hvIJZXx5978VJbkEcV+Nt5cyIIB+N7zP+vOI9dEYZTG1YFqCconlTOT3b9wWTQlaxZFdl6WIQqgm
cBIfwdycq3eJWzQrP3dn4lF3XUglfkV3PU8YS8cLrIS0CHLF2yEXGJNaU2LQtKOqw8Rng7AdjwfC
0khkOD4g3uXXZYtsiJdagkh2fXDHsy+6nLHy0NItRUpffE3IfPxSRLYQfbqFEHiWA2l0MeOhR/lQ
LNck9z4JipafdNkMYYDU/yeifNDUEvha3NPevukQYXCDx6bprxlcc9AbSvL41MlOepBBJM/ObxOJ
T4y8/uI9XtGhWF55K5dK8mmg4sbKwPBFl8H5O3tC8XgkSsjT1T1thk6io1EJ5bI/bOKj5wZfeCxE
5TTo9HMoSDwNqyxopnu6/6P2oayQgJkYw5R2wfA0Ab7McJGt66852mXMDAOwYKhIGzSMgP93tFY9
MSSewYM9kZnVNce8Zu26sH7PufO73TIj+qOlRUJfgeZynHBjbMZahDpccc0pR8Cj+4OMRaJKnUQi
xuJgLTzQqoyc6cX2NN3tKNXSMDxr2Lvucaup9Z0FV0NXxQ6ITSRCaYI3qulsjPTJLR1Z7qp9YGgi
cVrW95a91WO+lyXX6bE9stgIa8mdUZlh4LaJ3BwRSOwKm8f9FLfVAMtTBej4Eds4hfTfp8ETWOpF
x8xGODFH34EP3FqXP1ITpz4wm4ocY4EXLW6eAlb02Hv8DVkORe4jeIOl6VddZrvfVFMqO2B9NHPP
GYMSxfOIGD6tu0RUFrzd+7YvMjF0N/xLFHPLVpAzWZb2/rrDf1e84cwZYVWB4EipgfVUjAyan1bY
VkLQJ+s1b+lzgDmz3pTFQ4Ize/FALuwm/iPn3LeIK6wMx3Crgg6qOeN+iJbApHJe/KIC4mNwAC3w
i4nXKBVpSL4gT5CExDDBvcyNZnGv+dT8XXKRN/Gu4qkniLtixQLUrCmpKxosSNCjltO3zHUXKIik
7iOnNAcDgWd1Az/QdwphQz2e3wwn1pz/On+bPHdyBIupKzXEvfEe2rSuX+Zq9F6/Gcf+udHtZOTO
eKf6TDPylcKzs/8Uh1ZiuLWCf7OGdY9cQs05F0M1FaGPV+pljIPimV4iEZ0G0OLMKabLt7pr5gYl
5rhld+iXSbbQz9E0mArUydz01oNM/IEEkwuioJ75md2D0NDaPToWgofbYDgzkPpQPU960AfAPB+5
JOA6zqp0cYpX4SRKpEDv695VhfQpA3GUYBCx8Ewgrqm2TVsoti9gU/49ytAfw4NZpjWQoiG8osei
zk/fVgMG8l0D7vjDQnifilTXkuje+YPsow9JBjz5gY2xAxPqqlZY+VSA/4dZfLKTZWs/oRToppo8
mdqNIdL8LayMcX7qv/oeu32j8QOjbr0TgV6HRHkWKZMXp9/POGJC10Dhs1gpXftYD1UKZzEbarO3
H5vu9DnVUru0QzYH5YqqkLUey9VjWjaA8kgNk+KSUdhnuisKszyN9F80FoXu3CnDju6iIJA/k0ev
9lkN12ObJnua2ODAanLK0fzJgoszm0GRSl5Z0A0Aw17Ro7cGmtEnxaqUcltPBODPbuHqgjQQFm0t
hDoHiXQQ1QFb/vZ8QH3q7uNNoczgCYsnwlNQMurLU6XbReu6N1LsPKBAEjWj4Dljtp9XXEgi6i72
suWTgvoyChOzQJugnP4CVLLMhl34CfSGZqrka/ofp9wRysapwvOVsBnrPhYn/DvyFmbSm9cYSXAk
Y/PVQb5dIvJ827JS/xjxcZFxkAoIgFioNnjzWHwGEEe/qEKNXFGBrXY99BzR8c1cN1HfSdOHRSer
eIiR5U+hYhVTDVjk0l2MCvhlC5M8dQvlrJeiYToVfhGsjKbHG40Bl/BAYWOaMQhIHMfKyTFwOe5p
ROAvLYPsxSgFkEDbbTyUlKVGL7gkyxi150OONA3UxbwrBcgM5++x91hVuk7kccgzlGyFyTV1Jqd0
xXA1imHq15eRTkL2qNlKYOYwRzaO9tV16c06hKJmOJ1SAPHICG7gQ+z5T18PlGUYD6bvmOy/AFo1
WpQeEBLq16nQmxi71lsl4rwfUs+MSt2CHchQ7tfUGoZYxuUBfivRIkpUY1i+WfPLjp3xWSKeDdhM
1vQjdaNUVRRVGxUaaU2BNxT3b+c0nACLPuNRSbRS8/wX0KFIKRIsPLEzUiBif2KyP7GKe/pZfM+x
AxtOs9SbhqiW/g1s5eJtWsBt4xCj1KGwzFjpaSeG7BzMekxISh4VErvEu7n3V6wvYJBNsEc+1jKf
o7qBb/hlJjLfm99oZyfW+3KSEcO8DA3lF0oylu1BqOv1AD/22Hjarc7Iz8CsT6C7hms7gp8KVNtr
1nMkrgDsjifjjt4q8UlzVEj9+oJ9Gy4qS0UTSYaod/F1Xw00AIliVNV9PsRZlQhiJr3HaWnW5WTo
UKmS29F0OzOkYzXvPLbzA4X84LZNvoWsXq1BX6HUGzzNk8ELXPBV28P1yV9ogtq7pSlWf70zBFFI
StpTBp1PoXUjT9ixflluWa8N9CVnkgTELCNJslsJ9jUzccjM7as4dOn+Wit+N/qe46we5UahDlLE
j0djDaiKREu+HP1sCB2R435z1xvKAxA2cp8wzG7hGfIyULzCGGWt8rR8OCgote9fIMp7+ySDMvL0
xwO2ZEFDAVXhUZlDmGBYg9WMdcKTEOANfLp/uBvWLEQ1BuhyFo1ztcGwjA/iaeI9AsOz/6a3djJ5
9Nzjk+SE9mmd6SpA5JEz3iAnGt38KF6GB2c6EoQ+13++XzqevnUcuoTp/9C1A5kCG4zfGR6OorKR
9KeEWIo4xeAQIvmZHlcp+SK0VPVK4uM411g2Z38YNQjPZeDWyp4Y0MKpch55XqWNs+mfvZkyOhC1
OCGmec4RzGyTuQWynL+EYR5TPdZ+zI0x0yHnxCjayMz5egcsYObZZAHiBwi/To73QQqs1tCVrv5T
uMFxvVsZBaW/MRIslFllSJ/I2DxG0UR4mZ/4B6ae03tHbljP8lqPTMKHyZEKfrZGzTrtRoPTyzR0
c2x0HOt//GPHVzdh9KnMm5qDr1N9w4aJxZFLkKKmq4/5u49aHynM9+nz62Hffw+32ohD7yFsjDz+
cLWsaB+2iLnsKSkWasGyZWkH3X/5peaaI5aKbGq4txIxUajttcKG0XRo69+0/c/RhfjpfjsO66UA
1GISodAjp6gRlugRh2OCfUDIIG0wOTDNsISXz7SAG1rKUJ0BTRMfX0dEVZWhIZa2YJBJNMQhNLlg
4Lg90B/YEQMJDrCjppmGPlXv2ZRB5zFfNXN7sdKfbyP/Im8QwOBoJ0c9p1l2HkBG2ICuViTd0DWt
IdP92di5fe2onFb03NDV2a4IEi1xt+L8zdMY4jM64vrEbQl6S+YWdSWMhiR6HA8eKR7L2A/QuF2j
c2c1FXXACKL4Rc1TnbZAyycwHlPZWdpU8wpsrXyLdoaAGz5JGxLJckLQhhAY0wTnJMoZVv0HQpVF
pYDlXQyhRJXXjMI0ma/UTqDB0xCz5NgXe02Usx9WzKoOVnefh5mOIrQSAlKcE3guFOwGoMmxWNfP
XXcErj+aLU/Ipc4y+PSW34AUMW5Xl/4a2UrNgWB2AEhFmgJbkKIQAw1ZBeS2dtTPHIkTJzvvbwh0
1wEL0bKl6ZBU+LqmNybJGTFEwkRoTiqgVq0Rt5f/HyRBL9VAAUQtT9xb6eCdr0oU5bK+YBDDB9mO
FC387fT/Pjfkvd5TqhsiCRbNjw1C+Lq085KMeatpUaTK+6ty86CF/VOGBkaAcl3Ka/ELFV77kQgv
kPcSZ4DC3CoAmbk/IlbZZYXsyPZtHWzr53Ys8gstY5jlRH2F9/oQthqpVnJ7MfTr/kmEoMPATs+2
ONTo0vuSP8dRBU2nY59BR9bEIlVBDL6jYseYV55WppAmu/WbbLHD2481Ao6/AHXpurI7PAl/x3s7
dJMmPcjsbHCUCsmHVYwKgru2C8XlmtK3CY2MKqPS8j7KJdFRq+KjdOvsgbFUGnkns0ZyqeAL3KxJ
eIefxEJpRGigBdWIrUuEfHyXsXesj2h+dM1N4cFzxCgWP1TyZRAuxUNOZT7Ct2U5gYGkKa6Ic/xw
OngTSzoKcZSm/TXsOLWRb5wMBcmj8LSo3mZHHCk8JvGMbC61nksotZivNmVnlLw1nUkj9swZJpf6
9s1UgJ+7iVhqgmlIsxwU0iaWaFWnlZHF1pqWchIypPj1qGV0k2o3YsIWtaoun/m9bgH6UODkRTz6
uVf/qzijMz3d+SjJOO+8Lk8qbnjA6OtnVteW4hCDpRZovjyzC7jrqZ/a53FsMQktIFmXKkTJ7yek
eW+WRZtaD8bn3UFy+P33jOui3nC8i5y+f24sz5vM1jE8+pL0zHJdJ1ql8LOUZ6P1xwrxKGbvdMPT
QomN/sONZWKI1/yZA0hU8rAOLv/m9qro0bvZaqTsHa2weOX8AvG8VIBLRYSLWfp/rfS8MUTMYi2l
zCBJx8NwxW2kG9Z+eYRsnp6rYPv9mkK30h+3QRoSbz5nYosXGenyKK4gFpHixXqfFeVNHeYXWF+i
6RkbqG12sIxWbvYc2X4dLVSlmTgORkh9r6/p9Ghf4vBCm/75ZVE1z/7XkIrUxX+oH61+pPPGJCTL
7wDhbgDX2z4qrzQ31hRtDmdXEkinYCb8poFEygGfXgEhVAxOuzp6cX7n4JwnFCYI+4o4pjHqPPXI
R1i5e8IwcyWzdpKflU1vg1m2HtxbQE1b6cLD+7t7vDpWmg8a69DfN1zwDoisMDSJUCjy+FEd+Djt
nC/AcaWRr15nk4fbu7v+QKrMn1wsubd1OaOVfdKgqmf7+ErTeEGUDRAh0ug7ftEuJm8FeulWyC3b
JvIa9BmbBP8A/b3/n64wuI3vvTm68npXnd3wJpLONZJrfuJ2/zcHihnQEyEpVyLr9N741pLgRCY2
rxZdTPJk/eHROsB52bvT9WMSRvP4Q3gLpGKtP+fgAdXtChTXqpsme7SRBj5d6ON8k/j6INxbB16n
5VRS55r4JYjH0/MieHJy2f30EM2Ii1m78/GxtlVxta3QmiiviAsnrjT9BMHjpvWH33LwHW63l7ck
C8F0gM8cB4dHFkKo7LAfuSWrVAxfg5pyGEvzqBZhkvywEwJEf6b2HIwAnDqvxLiNjBdXw88sVN8z
Rmus6DkcTu5o6zwF+65kzj16xcplfBlTUeFKnH6s3WKX08O1dHkCOV8l92swQsciIMW+BxkAEgQq
A62l/Z80oaomIVk8d+IyNCQQWRU0XhYpydIgf+uC+ziZTnVUy9bzcOgCv7WMl/vwH7HPAmEH2TvI
/zxvNqSHmlgvOxSHnlhx78rnJ38KA+G4tto5CCTFzX2ovWbOAcryJ37PAZmhl6kVmAm7BpuxmTL0
+BrchQh4M0Ki16JfyjoorgQZYpmSjLey+/e/mNWYZ03OOOmafJS2gkFB6s3MTlFq3oEJLrhj4Jjb
qV88Cp4pSJ60ct508sQ/v1C5KTcLEfwm7EEFXJ+2/CUm2adraUvzkH0+eeStuaQhapJZZ+4fwTYW
qkQCPyseJ7nKCgLApLCim1B5MRBGHERbyCyWGpG/nitJhdWxECp27JeXltfhKq/wCFSetcM1hp3e
JtuH4nEWEBufs2Fygh77DI0aHQKpI4dE+Fx84ziXUqBA3ZIb4jKvzyWx82gaS+7n2fHQDyt2ie0H
NflxUEcEOEJHhG3rnNE6RXLoqXJCnMlwJDwkDDDtPyIfKf4r4eSyZ8zLjXXDFuYPh+w1/hQxLGi0
L0VJgFuROc8x+yuUB8jhmHonV/yshCKqIqeg63JXX/oJoGNN28z+YZVI+2h1H4EVxilYFK3gWT31
AancZA3OVXMF6CviwtZSE6nE9e+b6VqhJ6th9po3p4f521VlUnz1Q0kWDLhaqhqbWtUIL/+j0pp6
mpDJN5Qp0+pJHCpJDbvXGSBHDnS6HX88K9IiAhipYzPHrcav+CrzcQMRC50d/NfzvM8eHLxX5Rnf
b/eWooRB8NTJkbxqItvh+B2c7RTU93Dg2bJQ5F0DFgh3DuIf4AUS1CS0cFtcW7U/FRbsRBhSaDfS
Hvm1gVNsEHTyrmiomy5FAx32ge8B+4eRTtXz5XyGFe+xk158hOmh14RI6gzkH9EYN18d3oKGr8v/
P/vCJPU1q3ss6MBhXJQkxJi76DuwvpE+DMduWjgaaHHcYYIp0hn2XSRgxm7TOcesQuL9NE6kvAus
3PbXPoC+QNMrvSxtBKyyxEEJ9i+A23/CW2Ofee+AkxRdHmh/hUqf2aJ1LISaakjYRO6I4STJPYPK
WnW8I2mN8/6eiIPFHEVMHRJfGNU3AL9boZyPbWuqLsWuMRs5doSS9Mzaywh8lBHAF01F/yGIJO9B
95JQa7RxbSa26MA2koArULGxLysxMQ5Q9mUzT09ayS4UtBJHytsEmAiD0l1nLQi4O5goEvODKZxB
yoMX1WV367t+2hhh5tXSV6btYGQl4avN7lvIs7UHtz6cE5ZsyLGN7Cb7lDSTscpT7uQHOWkMffUE
XbYlsny4JPIcbI18qnvJbVRRmtYwsB6jP1gkr0u2Gp7TzZcoopg0DVMhIsGxId3bvAQ4sI12gACx
H/7j0/6SRcNnwBjyohMY1G2OLEFkDWyLz3qnQgrE7U1gYzvpcQ7ORM9RJc6mu0bGweXXlnrUJ76O
IEEcjKrjhaGiz82cZzTx6WNEcpCfX9IKlDkT/r6bVm8Hzgn0JwKFj0wPP/3wPhTXe81vSpfnO/0A
YjAolrntwA==
`protect end_protected
