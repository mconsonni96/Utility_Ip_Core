`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
VKdXCOhNdYvb01pN+yybKPEvVi8D0BdMO5vMANfQTgLY69Mq59FJ/mFDy4TlJiJ+Mb0yJtQLPN+X
ADXUoV3z9rInlNn7O9j7DfiatWd//kl2fc5klhX8UGGfSFNITSPks+lfcTZstLmB8f0kT+FxFpQR
uyD4y+UCKNxIC94qxqctl/Wc/C++/NyTlluww3JwnywIvewPDMUehQTaZ7oL0GiIZGoDCr7F4Qwo
LOZrBOZcG/IjomcyY+ei/Y8Qg/VRjxHIDXYIfoIG1UasfnK/KUlEbrpe+eWj8SLTyVC2EvQmv52e
k+E8GdlGbksJWZTCUWv5dNg2Dvsr9njziXq72g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Ntqf2VwY0hveKXnqxPyNmeutAvBIUpT/duu4y9NmuFo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15456)
`protect data_block
f6Z/H5X2tFvkSUyDM1EU2RFvDVdJRyJEcgb/cxwW6dMCvNkOUKUBPTs8TxaeJFEe5md3iAlapaaR
4usS01A9GuCfqdiaCRuOu19bFgvjoOjUP86rvOnBw3gWLErxqvOoDb3zBzAcJt3cn2x9J5deUAna
f9DlsMNuseu1lSM/6gTzbsC77M1j1UHsEPkILLhPKXh6Rcje45CR3YlZS4YeNsAEEwvWjSfWoIlE
CIsoBB7acL+A3WunE929mJ1v6SEeysd+/5lBWfTFOEOLeKmyp5iseF3so+NyvouEh2IkWYEGnYGE
RJdN3KqXfYZk+A6O9mStCBFn1j/dnErVHsylYeAKAp+f4ka+ttZqIqb2xvBFc9TK98rxrPrEvYKK
Fgwc1i1Vc4gKF04754zXlAz3eGXamjQLoufCYe3zPQ2PeMfzJDX3J901azCRs8w0luh4nRrDEkD1
Dy5RxQC8pmLrHj+if4zVLE3SpLouGx8e03IngbLaJ5e+M203S8qPCUX9OClwvE/PfRwtQq158vCN
GKDpPe/i++imENZdB8A6KJcB4cJBxGs09NezpKCzceR23vVLWBG/MMh7G5Q4ycHurtL3XLFJCxb3
Y1Foqp75y9SynjT1zi54/MLdF6eciaKca7tguO0diMPpIJO03Q89yyHSW1PYJxYNXTKYjHt0MrCv
G2nfbFaT/YP2R4tryP6efIvBCfVwg5UPyB5jIMPs6qG2BRjPdHf6GnhLOFZZkeDQULFZUYiCktDT
isELFyNvM+1XOWpH8GZyvnTYvJorHwl8aqHa13L6go+gt/g3rssDTCjUKvVNUC+zmWH3xVXCfQ3M
EIabYNXQdmQxR9BFMBCHd+RNr+LzG9c4aSucKo+is2QR1HhNGde9MKmaXZcTaFwUJvOC7Az7xlV6
MCl6FKsJ/ZEepDxI93A7SKbf00NUzIttY1L7g5UbPdC/irH/7YVJ3f1agjrF4qNFnkZWRic0zBZ9
fj6n/UIRBdBy0DAuqDfQ2+a/t1V6xeIUPDZg4bvgohz+9vs5P2rFlvTlpz+3QwJufzH0rQaMwcrA
1aMpvbz1Ua1usw7L7Sx1F5FmCKJqphhTWnGr4qi8qS5Wrf0hR1uvJrQ2xe8AI9pNKgyX+l1ZwFlE
sCAO/wxEazWX1AXhnH2kWkGhXge3atFYZuqxlRWHtrnsDbuBFGDlsToxFYaeywxOG3owKV6k/aG3
7jL8yLPIp7pWVHeRbF1tfHf6w7wcv4wtWEP3+WI6UHAnEhWtdnB8jbRbWk/TAdNJLtgPU0b6ZoqZ
aLWpEoLC/W9qivc9Vfm2QK0E/SjO8vTpUl/BMVPirQq8mLznNuVho+QcD6HRq4X4fxzx5+PcWcB7
xYU2ZLOixlwPjkFWSkFC+ruZsp3PFBozfimii7kNKWDqhiqN98BAn1iZ7kqhKlWKwmA2Wxx7/P05
3WAt1wxFGAMGy5Y0zmF6dToZcZVJzxlEQ62cRuGbhldpiqbDQPQr2ePAAO+NqEc0MJxqqNpGqWxu
EaWf0ZXi7JQ8GJbt7Nk12kKQpSpli60h/QxEKH/7GhqK/uNaKxqjgDl4iGZHxzVF+8NDRwCTnyUe
z7jofjDdFBo5QDl/mrPdIJKq5rU7iHp9LQnYtacfdOVcHzS/G7f2bpiv1JXueL+lpOypJ2rPhlsn
ZZcZLJaCeOtWkdMMTscG2v1cdErYz/M1aoAIFbrpIwvLQR5onNftX8Dp5kmV4TTY0jsOem/bORAl
m4yMD0Svn0LihoEOsm6/Mt5OZZB3GzYMM6aGACr1UAUymcoeyQl5L0kpPs6FD5NpXrepB7rzs1iX
TnNa7V4EeZPoDmhL27x67LhXdnQG0r8gp+DTP6jiZ6/0Cs20WrmJ3TCmf6KjvfiG3WNbpvDt0K7F
UEXhOMyH11zqfIvhO+QTXV/Mzzdur7NCzC6il7fFHaqlAApp4juOTDNPAD3iVYfK8U8LZmbRgGJi
yAdAjE4uD8evhAQ1cJl1a6yC/5EkXxeXew9F9NhxXONSse4p5yIpcOJfGiLDotEyesRvjZvnM9st
54+IW/YfUSHgSzu/z9bhdCJp7gjSGUJZxq8O8IYbAHYSsQu8qEoPFZJWa0QVVCxYwcYOmCTBfGnW
3xBTSbpOQ+faBShTDmTNpwSETlviqBB85B7qWUzNjwU3O7IL7uLm7/508JNnnGH4l9iDqbD0onxX
IVsc1Zac0oCU+p/507pbRPaziCu+ceoIc4JkIyn7pVkGrx+Zvr3F/fvON40kRUSiAVx4juhZsNJp
bmYvajFT9a7ysLy4CE66znMISBmKCgqQmuNJqZkwZ1ElWDU3H3qTRzOgT/YMGXkI/gA4XaV8KQgG
pgkHC/OuQet3Onl+hCKugHg/g81G/5Ch8I14ftsS8JKDGEU24/Lrn6J1dzjRkITS4ez+Ppr5t2pC
eFQojDZA460/ihD3vzAGbbE5nRztJ2hNW+T2N5hmLOwdVgRBkGThKArZDEjBEDSr8BpeSg+8FmIN
Y0XC2o7uvDTfQX/RG1miFg8qDYeWtTuStSIZ6f8xXxECicY4AjGVQyKmI4Gp+6o6QtP0W4opciuB
pkLy+AecyOK/XLESx6uT+UzC2xR3vHeD0QLw2cP3ZRxIGkQIvQqdnrowUt+3hllRJvUj4zguaOCI
cMH10Q4JaIbS2e9v9SUMFPbVPTRa0YLl1mYTtci2kG5tMFzlY03RK1srQU9xxvY+CD5UKsRLvFC6
hp/2HqMIYkwDCOMdiNdc+tMSxv5FRiyhlTWp8xgmEIT0DkT/0bk0TUM8S3Ni3jK8n6ShTOwCbJpe
sQIwWylj4Mn75yejxWgTsrWaTETNjFbgZxN5XD6eggecccXsl/6QWQBtTD/JWlGokBDa/V6Q9jdP
Q0c53668IvOun6SV/fKkn0UlVrGxhIFMSnAehQaqSfqfwB0Oo8GArET3Ic186Y3NWYbUSpTAi3YM
bRWuBSvc2knvP+IK8S3CbZKsVeJi180n3MLtMhK9Wr4zDjGJLohk2K/FUhJNsf/0DolOHeeJCt4Y
6UJ6qnglobG/h3UgKVzMuNGA4E2kaT+S3a9YUtcpf4WgDe/jvAeS0JiMCs+YgbiSVor2RxVV+F80
93bkETfRMa/Z+EIWGi5Vj0IG7aKJh9jSgtdC9EKS8/uysWW5Hdt+HlaEIHKH9q7Qzfxfy8M4fp+b
ri88dWHblCzKjvFrms6dTbsyx0bwES4bN+RHrF/VBUg6nTTSdB0US581V/HW2UYK0mrACqAqUpGU
ylxIyIFtymsiSOfXDQqoVG752tRUR0WDDkgzFWWfCpXyJKnC4st6sRcGIl34xHGO3BvTd5ncuNsN
D/cRofv90gygT82pP22UXp0cuwxwqpD3/dIznIC3kXx+yr2wwZEwV/70hHyRDBt76NSwxLjCJaLk
FWBFWLqaEv6DD32pWoOc7AwN7g46ETr6uBuIbrnz4egsAErtNXqVRs72uze2UQ3OvzBr4nXyhOVS
oSpXCAZPjm5/eFZMOGfi1UjEJstOell9+qOen3uQKHaQ+2jQAX1rya+OCnAhOqZ6Cwhp3Oy8nXXA
kJHzdXjVSs9ZJgcXZ2lajHGPO3Jr4uPYnxbiwT8xsM2woDu7m4bzMZuw+M40Cp5txKZzI3WNRdDU
mZcbzaYXxjKslVU6GKZHs9bkb7MZMC79TRqQmkL0OmShnI91Qyha8Hq9sUiBihwXSie3ST4Epzpf
Ub+jAIOLisUfOCO3KO9m8VfyabR1eEPWYvBGIUBOrNOVwnsKThuP6vi8vyMyeDdxjUB9m6aoUY1r
SGM+ED9Gz/sn97HY+1TDISX95rXnQtNY7NMJB44Zg0vhX82sxzAZA/qWzTm+baiRB5+wiyxlNC3t
ETsacu8MULJ71I6pf/jjc3W3QAAfcu45y2lHuxR9N+lknGCeqhbPIGFp3JUQ8q/AO7RCPrTX/Dto
f2TttJZRyRpHzg+d2HULE2Ok0xhsrc/xe+fLWQKzeO+EvgwKFt67xTL+RoF2D+ayt5sOm6aTiZa4
YmgDx5jNVh1LHPAqyQy+LUDkBEk7Xm0++yBn6BtOT2+UECK9wqbOLCjjKeBDeYIm3oMT0xC+54aF
gvKjDX6dBeL25NQxyDe0twGwz6u7CNXmjo7bO1Dx9FKijg+lNiUYgddzM31AuWb6DzmD0/oJhF8V
apabNY7CoQ4fpRduZ7Jye1fI0jRNAXeqPn4ruFpfcMZt0pefPaaIlo3iGl3QU3kT6azmBfXHFr16
lkoRpo0Heran/91QBZFstmKJ/SafDpKmp6jhVuE3YYyMX3nvyuyANgIUhq/xOWQy14KcKstddIfn
TCqhlwx8eZRiKIjNVZvUCJOI+gOzKg7ffANzARm+rlCjGP79lcq2fimhSH0h6PWB9xtUpXpjX1aU
5j2E7DB8WsscT5MX7CpU3HaFVKsYH1HECjld6GWBHB28en+WLEwdepX4R5NqtE2wN5WvDkmKGJI8
ex5K6iETyt4rJyHUFGrKlAhK+EwJtIB+lkIvTgcjGf0zIheI1FEVWDY4t1fUXaVrHDP49PeFaGD3
ox13grHWeDsmD0QBlYkPPKc3Qg7Gjvgdl5CkGs5srS4a9kaJYasMttd4NA6Yy68+M7Qz3et5sl5d
tXByn51RLabGiw46065tFZLwc6Mhea1/lyN/L7oWhr7JxPG30TZKJTg58NGxzCQl84dzVDLN8Z54
+KOXHS7vgY+BdxQLK4wJ2vxCzCZBtSnslj9Lt+FSmpGWaYvcVgkSLu2HtvaAwdzBRuJ+GGr0DAz5
ic09L1FpDDc+rR4sxrYdry1kOX6byXWGi4YgkldSJ4ilFgX1nOJsynQ58oWCUcP0r7xrA04yN29E
lPtwzwT/UprSlU7Nar5rS/83sVlwXmNjN2V3SHSDY7kAhXyGwg24yBDm+KId4WyZwgjgKH3/R9SM
ch2aA49NG5OaODe41mz9tn0ptcrSlC7i8V3UIDrOvT9KK96dTJvfCuI8u6hQa/3lFHIZfbXyAoj7
D769xEA+F/rdyT+dENwvqGJLQ9YOD491Rj9KSiMV/+dxbn6asD3t9AxIqc7lY/tzATIwMA6GO4pF
FfMMCH88N3T1hf+ItIS4efs9yjwqpeQ8Yj/dqe7cNntEkKV5KsOXYEiXqdF2FI5oiwkJHBjAZ2JB
xFxgeKHpALhADK8EfQLTHgGVPnXsTIIXDpEQT0V4iCKQiIvS1g9NkiTBehMKR1Vu9rVDBCrnlLId
msPnsAXtKW4OvXglrPZJ9doP2ZEh1ItKdRATFtWCSLdH/YllgTibePFl/zSy5KpbskW4vP89z/p+
df0sZNrlbhq6nI0HAdNj/1gk9ZUyNQ3/b45qgrVpRZFNmQ6DK+mlSvL1vm2FQFVZIY9kfUJHnyxH
86UGgDRxHStxECR/lSiwMdK48trbHesNpGa/pzFwrhrFoKwBMTP+K2Mfgi9Zq0AQW/RSi+htTgES
VrrIGwtv+IkPSAHu07VOVW4AcVahaJFjDnqZpsZuMEqe1Z1wBE4tdPcpG5uyUvZ+p6mGgDaNRAFi
qcDAIs+8QxDYyroRl6V/kVGvXWzjcLDokFFOh2dyy5LVYscoYv/AueslM3pLJX2gTFytgJWkL0X/
FZYh7pWWiXvxLrhwqa+ON/NMX+cyd0FZr0eigJKXCwQgkRnz/mmbAsBvfhc1l2536zngILh4zB5B
K+KelfNoXmy2HOKjFjp9qg/9g8Z0rlVbM+VVDNRye+mKlMQGFHA6Tqdf9xZPYKcjJ9dMos+Jg6RP
ECEd1aCujkQSs2+RrI4UgEV8fp+DEfl5udj359K3dbnE4g/j49cGSfq9aEaN8H1NOo5OXRTqXbYs
/eh41nNxYKHe3TN962yaFsOKKDTUh4NrC6J9+Tr9SAO6rNvh/oGq9PoNr95rriE4Q8Gu45XAQdzL
cv5SBiKPi7r5EJuBsnaJFAd9CjijH5Eol0PpNnNjY6QOFS/5cvRbNFx/vOiP0BSjIQQo8fLOntJe
oidLFZ8kPe+h3CHKV1wbcoHVYfB8NniM13AgJs1h1rImqmcXJmQ6FiRR2sQcWFeheqvyC/nVMGGj
d4wg3dovClNiVhKEPXuVWr37OAo2gn6+Mzhv7L0DNzKf3bTdqrX0OQNc4z6TocKfdeDq2nDSN+fx
x3qJNGjPKCvhZQWi4ZgyhNZpnHhiprCvvimbykUaB8fAhALmrSy6/gUCdg35hW4KzEL27BtmAScU
9u9qeSZ62bgZlX/RTaJrwnffWT4LwBzY/B4JmUaBoyjUNUBtXokgcyvJvoVuTWTLS8KXVaDnmD+Z
ZJpZuCj0cE8JQHBMsuJr8IADR5IK8fXyx461fsQIO+CoHUk3Ukjinz1KTi6ST9nzmsRDi0WTZbOU
fTDPye/7H+yf5gKwOGgaiOZM5Xp2a2JmSLClboHahtOerVebD/hCMklGeshV/Tdl3VFDgZRjVBZI
2Hk78WrX7eEtMG6sigE1TecVh/crKj21apmJVKV45AMMypXfLFGmkMMfijHjNDeiM1hGNMh5pE7j
0oxYfNUbbejXvnPDLQWZuPUj632+PwSkhbiioL6yHObOraq/kls27FaFBc+X+hwdfHO5WHg3BcGm
cfa3tBT7FMEoH2JrkfFvYA8xUZdKoDohknW1ro0qZhWcMuA24O9N7DmjEl2243i2KP9il60AGh04
JCTIxCQf6klymdGGKsHwYk/YBDmPwuWogJm/t0hnj+yJZ11jqXP+kS0vqtdACyWpDmRp6r+lYJZP
pqUqdANBsgxEqWej4ns3gcjb/W5gLzp6reg8hdZM7S5Hl+FuYlv2elQfhg0+nwzJd295O7WNtcRm
iHA0sjaHelBlVol6zYqBYFJypudlYgjpCUs8Ji6VbiWPcFsGWKLAdnC157jVwvisOtbbZNvLGo93
m3FT5JdRu9p3xk41UoAgJEBNTPFwp/G+w0ShTyHEuWSnnpiXh38ug1GsnET8Z9ipnrJPLycS6NbW
trt9VlDANqCzWXvNq3S8BGCrBWxjPTdLxoB3papsCyj3UPl+Vf4TLKTXob2uLObh+oUkWr80LRuX
1Qzl8vJ1hboI09/MnuH9RJ7iuIKzfkdbQk2YdwjW/a/uIw9fC80BZY9+o0x/Ssg/NveAIBPuopqr
TDbn7bEHkwTXK8/zqmTbGyVxTbihHxzMp1qpKr3Cxj3pcu1pCTmCJd9wpvoY2wMtOdFzRlCt6azj
aMhnjxSUNOTrAH1j1vgpNcKnY3hgbkgk6zXXWgBPXhrvb0MBgyftt90xcIhvA5glZKcgBjfIy3zH
wYwHTi+Py59H5cVzGv92gAm1N+HPUtJ+ThLwwGMT/GuL2+gA/UwoyplIWR1cxfmj8Tgkij+I6RLG
1wylRAIcepataLGzA0P0zCwzNqKTJlNymZCLjXNM/H4GBvjhogVm544UNliV+AhCMnJqnfnPjcvU
A5BQKyOMKeTeqIk58QpSiDGmmspWRLPuih3UzETK/AY7Labl1UvHOZH3ARifbvqBhz37Ec/qwEGK
8D2/i8OqlZNUdJlky+bO0TOHF26pP7vxxduoOZOzYyz7IbP3kLbNu+icMTFKz5LXgLWCvsLgkNq9
qkdlgQWrTiJq275+uOSTl26JkTP6nJxfmBmmFaz4udP5SDJfnLRzwmYTHAJThAwgzMjgneApcUG2
2q2rpXpowz6N4lIFITZi51FKyqRSXUQzNlpq6dXoTOYeQeGU3rfECeveMsi92Oeps90eWPnyGFa1
adAez9M1E/ClKDM99kYDZ7tzOpC2NT/zo5KMQpZqP/5xMm2yhWs838EcQRrafqNGJRS5IpPeWfzi
fSP1pI12Mp84P+vW+aU5U/p/TFXZ6STqE0NavPgS6yLLZ1fx6O+vN1XEq1qLYw6xJFVQcTvQGmMD
YjSpkzapLefFKeZ8Q6tGthjqLhyLd9CzFpzgik3iAi+HxoXmAW1KVs2F1eHDoL/dOrkvMTxlvjiA
/8GzBLndUQdrXNL4QjbR017DLa0MHsKDNgOweRD8xdT5OTYc14jorjPEUbt3gyNplLLi1YOkmW5x
4ROC6rvcZR0d0C2gGK7dA0LLGdR4ncY/DHgmxxB/oWIo+nxe420Qg/AxhVfq9T2C7o0jz3h/ujtH
jJ2XeOaG3/VXI2gx4kU8A1uem3cSpYnpx3F5KY7qTnSUQEIls6raJhRaCtW79RKwhTukCQBzeDM5
EUuhEIqYnWXXQYLqGMSMIdCXEDn79+cTudfA7VdDtcLYzUY4ohEPBNbUMVxC8koU8qqAHK1rnKaO
NGnD2/da9fQmLjHLp3ho0Z7M/MpQV1lVj68R1eDFLL0mDj4ex3q4VJjsQs0X+jiEPurV39ge7Xf0
/Ao0PK0zTyw/s1QDh1EHWoYF/FLJ3JMpYHxhA/WfM5lb/xPoKDr20yt9MJ1D6V8yH0hay76lz0l3
pdGsjFOUzTjiKC2BzQwpUUy2+943Tc0BGczrB95qH3jUCwtjAIQfEP8zpo4c+zEXfj1iir2CjYPZ
lwGgCq86Jgtk5zYVHgliJzsBfbm87KiEBH6DlXSLIUGQWD48OCgYx6IGN1oEQtVKfyOGs4uI1/3u
SDnXaOnws1lzOrHGVT6PsMiVJse02f/kT56eZqk93rNGntYwv4x6eRLpp/gTJehxAY26I9w/9o3c
JkHaPnBVCQP2Gmv1A4B0qwALJOhcNZ0ZTGKKsSjqAWamAfriVrroq9Qes66HLclTiaQ3fMRw59d9
+Jqar15sEyHWxjSJeB+eOD0Fgu+3sImGx2tyb9sy923CN7xCETGpnO0GQ0drenaS/7MJLnrcQgQ6
b4Q+uMP4tDEoFxcbZHGjzBRKR5PsQGBoS4vWDpEVVZt5MYuLMsXWAm6avmyz33pd3jOZw4oQkgqK
YdjdNTmr3LvLEv8accxFAor04IhjtCMLqkkWcFRMN7u01k8CIC0upG25y8SRj0deXEfhucbdV35h
WzZk7Omusr8Oa2Uy62I/DWelCzFvBrqr4wM2NveO+AvRgABcxPAxj1Qn9F1dNoccfXvv4cFjpt2P
bRKgQThZ7Gr6AsTC6skyrz2h3zEZzHIOjFkmDfnjMjZ8f8qW0FiQ1WD3F2XlKD5dHEyUJ8MFVdUP
1FwcwjsNWGqfesEY74QXlJEtdJjV+mJL4WejVvbbI/J/oNEYZu0qgDlQJjjtkwl3xChwE2rygMx9
lo7mDn78tjkIexEeKeGK9fO8ylb+J1zcKet5pSBbDpQ4U53FP46XEs7Ol3b3lA7YltApW5m69Z2Y
wK6NMZxfQSyxcJW/mNq5fBLCoHljL2Sh/ZTjJza8/1L2O3RFJ3NCNS57L4XPWpG5WdoS272IFEps
a/S0ZmaCYeGyXrvJwYJOc//Px2toyQukb92SOdEJpk16HWUATprQyPkrIvR4NKDgTqRLoY/vllqT
+l4kODMhU1JH73WX/ME/mZByFuEX0Y42bKqLcejDYLDhiExUMsM4QQTmKpF8I8IzItl7uwZSK79G
rWD4tNRiUjSD3TZHSPRzsb6QsEx9ZiGWLKjvYQ8gguIFTG+qLBvmNrYvTDILaMIh39ZHxasBJRvR
EU7vZtpcZzo9GyIqRSQ8+RuJ+9qDLOoQbzqXTml8KhSRQjx8xOl8CzW63XeQQTh2LKtdcGDraGi9
97ShN86VZ7P6N1kXNlYoKu2HrrRiJF0WqNirD4y4QKTz+sRd4sOXmhnSpU3RR4baTP2z9I4ZldXm
zCGNVNZV/Az5eiailCThLGwhze1VW44aX9WOnGBi1a8JR5qTF4eqYY0SYXL9DRYdDPsK50+FddTO
vl2h+lSVfnT8BwGDgYPaYZzuDaWWzUyO+k3vj7vx8fZ5WgcEwjmcrY56dXYUy+/y4A9qYZLfP0dT
7dL13apSJFQnpwhvxT6aL2II93Yw6v8f+hrPnp3S6pb5bpZ5wzikuHQKKUdm0DVdaWfRT6L2OC6r
85J+DkFK6GFfINa1IuDdjsclNEV2x2y5LYffIab9FZ8Hq6ZLk45IUUqaJTkPSqYQZvURu8ZLNOtB
/uEomDU40+CSCd5zF5U3nTACbyEBblwImlTPvchzZYR3lQwsaBP6CMKPzj2KaulktmUkGL0sU2An
Oxtx3vb91cDXfLE0Hzf/L+w16/OhUwcrH9NAtNaMSOPB2vIu62UNuuhtfuUZBzAegESiEEgfj9zF
mPMseX8sKMkIsKFFopzzxg2yF3iN4rUNV/aeYXz/5K2V1Q5lIizHLwx4+uaxMNDjoSJPPFzD2Y25
1b+g4P6xfW3/lAgV8+lKnQsNbbYEWNlFsZITf8F8vDBqqHPw9aokRKxwqm0r/fus6Vu+l1sCccPj
dZ9S8NCPkdA+ePhmHedyhsVxO4wqw9PeoHSaB7zz+ksAqjQ5UD+uJWnDfEdVoyvSsdc/QEPyoXtS
jwEvEhdck0zo4CV26qlBPHL5dPK2HebYdFnuzD/139FF+fyFeCYz4bbnrincvUFtki8IEtiDh53d
uKjI4lfMwtGBKcmCio5zaB+Z06zJzwy3KSGqz9V/l26Hip/7SIgt3lDs17MXuP2sTgtkpDwSxpSH
re88Fbhwb/gJMK+64B898POYLu7bc/YSr9NUwTRBfSpfnSr+3e1erKDOrmKC+FIT6g415m2gpYYU
0sBuymgkg7weeca49d9RJDRKJkZvowRqPM26vHeraIuiPnb6T9IBsxqe2ZKvvmxC9EuQW3GMBwoL
WyWgSOr2mUoYZomG3Yq4Ma0vM98tMzqzjvaVPokbN94r5w3d08DW7sDgbM0pxRmlWSgUUF2xWKMF
dV0uQiX8lQsVdtO5UAxm+Pzq7gALHQP6AIPtEYHdmkbJoNbsstovjsW85EyIS1DB37Ba5VV8dOd9
B1sUn1nSepF8UwvLDOd5vGSOPEwcwt3AO+2o7flhWKIni9B7Am8BJlSQZ50ze0lDhzF1woj3RCGb
qun1TUQAbnGkeKSJmNiZ3KOsql4YRhSh3fFUv+yUmEwpcahH81XuY1FH6z5Bbe+PSaGDhEMNykkg
l5QnqWs0/433bDvMx2ttMAFgwhVUaBg7UAcZbbKl+kDJRC00AH+iyJKAX2dkGbU34i+CzQEsNOWv
x5bE2jOMvWdDZ0jUWe34XSsXxZzZ1fJcCsYAGHtAC24m/ePw147c48wgYLaoahC7oc+Pu/aBhP5O
v3cXbn7ARK6YtDHlGzW7ZnZWKP5at8KaWv5mz25AGew81OO1Xs3VrZy1sKnWz6aii++2RowIUHJp
HNlELKClVoirmRDEM+NpX+F0n88FF2fuP00tBthhCvx1Kel04W3xMtXNO7YlPZvXCg+EhTPYPbDp
PSiKz2jGQBQjI3aQ2+BzKRENo55Wv9XmvhFsBmOg/hH57uef1+nv1agMsj3rn9i/iJ9gRWlHKFCe
mnSg+KNBPEBmviZmyPLcecwLTsq469bVJdf7paRT7Q2/+1rZBKq/wfYvol22ycOkMtRZ+QTrbafV
sIAQPsoIc0kIzozs46UmX+ksZkSlQKbkZCyVdM+BPLn7eCENm7ppIGsdJ4KPkb3kR1be+ad3mrpU
ZKXmC0RZrbnN/mkkx7TguqYJ/0eBL+jo6ynl18OWO8qgvkQ5BmQeDPzBFFekF9UcwyK0STWQ0iah
H6g01BBKJDFU22cEhgM7tD21IZyWv8N7ykAnIOLdsVhAdPeoQPCCiY4q5Vg/S5CfI9eGrQ8riXeX
fViyzkjE0AYdTo89TX0rL+IDGbAAh/6b0+n4G9R6FM4rP9XHBoRfvhrsd6ttzdoGGM0KDYY75+/s
xEhjQdjrRG/WsKpVWfa+AF5Mzy/x31KxJ7YqR9XXa8/zakX9vbv4exk0pik4JrqkoZuVLmpSHYdC
ynEfW6mHsc2YU7/ivmFx36LLXrC6Vou63b5FqfJAoxOORg8zfgwu3XfMkPnU6VC1byCEneo8/IM4
t29XURqg12n26ESqinfNCd5msjNQ7EIRctWTTW8LwT6sm59BuVRzafi4GuGPQswbSY5DUIRXlOxx
IfDLiwGL9aT7brm/LuoU2NE0MXZOyiXXzEiot695FLybEMRWWcURoxo5CTrk/avC8aIdf2wRerlO
HQ6Sl0ubl4L5RvvqGlOG9nFfruxC2RjRh/Nf5x9ixGb2YaaOjAgcfmhIIOr2vv+RfxeNuCUyRaog
pVhDcKOPp8rO34GA/WsuPe+6IMoDGtLM40x2U6K/KQwgKhr3gjopaIgAreArH74o+yTQOwh3B7Ix
TXWj3Qj5MYvzy2J0Mp90KzvhVD43IxuPdTzGPXZ8YOHgtjm3N6yelqIdREl1HvzXnnceAamyHuOi
J/sgeAzWpRDpyupxoS1qQEv3Zg4yk7wFVf8NQPOh2ZQH6gk6rWz/FBsP+bt/QtvtGYj+EXqcJXFc
FDS2IXvwBhCquaJGjdeZ1ZG8qQ/svqGRiBhsn5nYuyKkJ7T//I9Od3GXJXo0QhDI6poiuY/VaMGY
cZvcshlocdWusooz37xwcPhPoHhAuUaNZng3ci/GqQ3AEVfxAkzHimZ1/2Mg6etIeTpJV1YQary0
yXJBVYx6wWZPEGuBk0SJkHl7oenDrqKA7HT0gIh+GDOKHBmbbdzcQM1gQNlD8lP50VtOsGFjQoC5
sO4xDqhvzpeDgCqXYPN4ab9tRIg3hFttK4iaEMQEP4p0UNEl4YYKB7oDI3l3AHZ5vqSk7zZaJxB7
CGpfGupVNbxfhigAip12XgyeUaGzLEiZijZiUD60wp7q8m0SYvDYJZNVbVKTaO1tWrE29mtZYMrP
2aQt4LMSFZOyiGtju04Pj/hWXbtvt89YzLnmz3xEeLzouV6DeTCG3Rg5maTGO1+KXreCywXKLaam
mE1WT5pd4FnWODA5tS2ZE38nQn51Qt3vtk8s7Hnm9+wb/T9QvL2KdYY/XX5ODeIpUbj5u3+ooW6x
IrGBYqzdfBQiD8MUkMNqU+XEaVE9yjw7fD2lDzKgj6b/HzxlGDFbLlJ4xkdbB076tinfRSbXKan2
5HgiJF6wRueY/zfyKy7ovqAglhiU+OPRuVAAz+I7+rqa2li9gthPwHGaX5m5FHoUbYeHkWigGFAe
1uA4SQ0w3g2uAegUwsfPm3hqNudc5Fthu0QKlpYWLxBlhhF5emO39KeJckbbycvNpUeIrfswzYco
vCi4J2U2eiOWjISo0b+ul4mnSPlmn45X3+Vig8qzz0mSVAlmiGaJkTeXAH0DU8EwZt+vPRchTFYL
y4c3w1Vopvd1VkN0rLWTRQ4mBSo3m0rdh7QkpgOucpygBL7ziKKFWv7KO/5I5pW04/HnulBivoCM
xX3YFyBwlgD+009iM03BudvPIzjG+xdecOSVKM9AKTvAD1SSiS7cFUqq0S0XkMJ21P2XX3rLs+pE
oV4Sx/2TjQ0SFwBSBhHbh3nJTOuMOabwETia2XR6aiMuSCB8IUbrwV7/PiFWtDAkppnCevcK6nIT
DWvHDLpxQOm+l6CAD5YBd5Gjkzg9ADzMNlmZWEtuqIZ8Y2a2Fpevns9As6QhO/C9kY0BGV9YMOwO
Ekr3HR0UiyO+VW9iOCU+sDT4nSKQOWsoEy5Oq2dw9SxKjLymGBsUXbGQcU/MgcUyS1Nz6MTZEFeX
A2gWisWxn/lhg2uYTiduCjCvdq5Br04YAN2dRPyQTiJZyWenS4XZQ2L/gT1Km8QPEQX/JExnNQs8
CJKWUkWeohDyuH01+7Z8qC8g3CCo+v/+8Z+vncR/4Bdw5U0C2AJ0JzOUF5eQESgx8bIPuS45a0xV
GzV74F84ZRo8BzjzlcQyh/mAubeoG3SAoHh3bEVfMk6sedYnLwMWuMj2h95eGEnn92K+0bu+6Q6N
VlLDQYViHHYPB3LGfbaInxbawxEppB7g8F21DqV5n/GpzfGhFO3MnY9AYMDMsvjrYLapz5EXrGgj
qu0SR0bqgAPnEMNMbOobjs7IJK1GBPMIwDvc2CQ7tSnJOjoLmO38Qa8tkSCaW/j5b0q9YkqRdznF
lODYvFMpL9ywYMO5mwkdtl3SOns0ESw8b7o8kvkUE+H+1tJCqBkwHjEMelmo5qy7TF4+cAGMmTIb
qWA3FKPB0vnWdz8kpgc24W4Z9cREhBz6kkjPtzqYAGMLQiqLT4NDrVhfSj59IieaNL+WbostB4/+
t4MULxYswY6BMkPLvT0uN0jjIL0ac5ZGf+NHOzFwJ8bKaNUacSEMJthsKFrC9dlK9VQpY7gMLt5n
bFDVSWfYP/2Dx24ovuMuFuESgEmgN2+bU1tOG3BVUmbsnZ+/Fi25bYhAglKttdwgiFjWPLrJES3C
Ib7KCJzTsziIcjbHbah2avpgha/EcR/nagTVLYQQD7PGfJpVZRNVcJuLSxZ9Sy+lOh/LiXBFX26w
8EvPGCH7Riq4e196nHb/pKWTmsPhkrQGk0pp7IeSyQ/MHaihVUJFSfloBEqyyf1arJedXrUZhtMh
/6Wktq8f8GbD+0u22YjfXisnayrwzdKjfxbCe1Aa8qhKjkaWO+LC9+9B5vC4kf+gYfhTXVM+SWef
e3HqraS1SDcK++LvcrAbJhMOIJcyOVnVi3kYYsHDl21GKuPnZBEhg5wGSMjtz6VFJrJJLUN+Lk8c
ZFhyDFGNqNA76fGY5gWecaSrGJcr6NNKbrbjVdGbVGaN9FH2ENlx/qEYA2vLexUrvECLsouJSmdf
eocmt0KgzCF1PP4GylxiKy7Hj4NwB3e5IYttA7RvXc6nnGJRsmoy1TtXfuV21jIWp1ukDLEhr0pQ
4HILMbPREFjOoypP9XaVDjd8aDlN/WhcvQ5c8I7Zo7vhDlKkEXziioaGoraehu/ygxvSuLGLi+NW
3HDbkPXn7TOMggpOV3NhjmiXlV8SM1Tl7DPJPscS3+kM9nXYvJYfuvETm5y1JtjuGoJnGveE9NcR
mPB7v7Cqg0rhWA2Un4iAc8l9LLilNvLSvSSfotyc6Fgqql2Czp0lcFvm5y1n6jUcgVlvnJoAwRZE
RN+NAFCQ0eninKyzova/T9kSEk8x6uL+vX139o+N8nyE6hZH9+JKStXs7xI5PsafAGEyFwdjyTSN
e0pqhD2NbiCKTVTdhFzj2vUIbAYCdcL8k+i1S2bCbYqTmC8GQIZCdFQAp0pZt/xoBOYATKbIN6aS
65sL0ZAsg94wMmQFRiL5rrgBbCiKiRSE7q4/AleCIkIg8J3qifTeJURufSpeTP/Nq6P3K2M//K8k
SMredypSM0RhEb4rZngRQj1hz0MbMNOCXMYDvayC47HC2RwyK5NRbHavbCzB0zCZm47yfid9LeDX
nQ8ox1PQF/SbzO9lelMGepPmb5+tZ0W2aZ/CwbZUGw+gQjfnrBT8npD09A4fF5YKOh99ZJKa/gPY
wq+anY1eIV+LgieBYiyWSs0TXFCpOyzSK7Lq9cPhToU5O2diMrKssgd742ACSCir64zD+sZH/unq
a+3oFtO2bF3db88GGLrNn8RPhZ44Jd5Ro4nEGTMMS39EozpwIMY4MF0poJIz60vnhaCll3FRlMSK
HM5Ck6/22VgVsHePYibMVhQUIOsIz1wWTstLfDGRam6ooC4bIXeqS7py6+PWc6S+pGpWWgJG1qpm
47CULokjMRPxlCg7nueJUbZRyEq0MTqjgi6mYHYHN65VqrnLVsYqXE+4JQJeYf617B/O/4xMdEzB
pRygKh665cLUzKVnXyiERTldovjj9pOtq3xescDxOz1OHxl7hrIr4nV3O/Y5TrOZJRDnKEa3cUv8
xBC9qZY/9wnZ9O8A6OAMngEoVU1HAkk6yarPWz+aepq5bzfM5s7eDcbUrpo6QVfQ5Dh/TxoY/4/g
p4IzJZ7/JTgKGconfBP2/bc2VTW+atS1PPraSEUAgGe6kqBeKoD24aKNIBBW/Cfrz2rflW8cJEE3
OvWI029/gkqtKqEOB6zg9tlakljQU7rkTlDuzkfdtmzpikI9jTCuS+TWvCxQt6rRAaHOyir21gY8
xjc0muU2AJqYZcFaoi1GCOKVturH/3zMokrmPWVegMnFRkuh6alDb7TCgsIA8miKLjuuLbrbIkNg
w788gdIEEDGoDpnYoS4R++BC/YbN6JmiuMMVWEYIIp98BX3wxXCgImdzr59W5ZmrOdSok0nvUoI6
YL6CXdmS4xW06Pnhdi+UvPEOCu2JiAcLWbeUo1l8bzx9v8W7MOfCItgZ+kbiiQr9T0MLfPGnYvnr
g3nfeGy2Zvl2bjxGO/tbWk/WJDJf00syvZL6bKXVLWwuq/ZEjlg6meSo19COfjDKl1e7ZFtGARuP
4W7g5eIRcjBxD+dtVl2AS1yXKeGoS1Jkyvm1RrccLddvRD5MueTQb0WYPUHK4CWY9vNSIIG0VbnZ
oxUZHNjGQhxXnEnS0F4n8PV6VaEcQfpARKykpYY9a2Zej4TX5KeBD2QVHBYNTqzP/MLX+rNuwG1F
QBJX7ZA9DJ+7FWCy3BPIkxz4aTN4S8Cw1qZDhGeLDNhs6IQfahquGLNWwUUWZ22vMZKhnhAwevTA
qI1QIkG0XCsClY8uXbZHt/BvR6VaE41uN0c2tStNvQtmBByCTRO+3mOmdweZtHGewonXwkmR/fCN
c8YvNmaoKpogIUH//KdLXuHUqMDvYvvWE6kn4zCv0rDjy6NajzqQH/gHNnXeV6ZwIUFqpxjhXWdT
VYtsHBVoGKRk5tys2TfPvt4lJIDZg+8552CqwkB/paZZUmSo+87qW+4Fin5Ap4fXB/IsYKSLH+da
266s/faP44mgZ00El086sLp/daRl2/TYxV0SnZET0F5UD1f7p29q9l2nlWTlSYll5/gw2auhmEBl
I1hVwBtvmxvUC0exxlOrioQTCu4V0HLCiUxlYZZLdZwXoiKjCx7lGim2fbVNlyvli8tduj7OIph7
XEc5CiQWvKP0gjqvVQQ9coIScdNTQtci7OsrYnIFSFCBapXN2wKvolm05LWcBSrvq7+/tefy4F19
QEUrtBZ7VzkJVdFUZd3wQb/eXqLYD0csrlSQQfP5Tgb/tMhCSxvY7Byu+rGnmfKSYiQrRYaQ1LRq
gUtGV5TPO/DCauustKi0a8BxyoYQUXUWhKIzimANlcPV+EL+VMioX6lq4pLtvCHifhAomVAIbRPT
o3Lp+sK8IfU8xPyxLR3c/RJE3vCpOzoIwnXAUcGNyCC01ObonrZvxh71LA5vGeCu+Yc92m5aoUd0
JMZBzs+zSG2CKgaIgzOJdOKMPnBv0MJUs5g/Lxs4ROxDCmZc42n51G5kOVklm9cvbJ4P9s9tanMG
dXU4xnoLyqa3ZY+QZEh1sv5fNvZpr782LlRWwMfVJj/zU83faDhMjUX/oVPoE17gIJIxZm9dVGIT
lkaJbvnWmjUREIKsCR8/4zW0klYeuOSrEW7zccPf0Z4mvtR19IKC6doF/ccD9YhabUMiowsP3MPC
bU3jGpyr44cciuvj+xbOLqp0yENYNMpo8QATnA247T7wzzoTl49datuHNcGuS8jEuZHyQeYCGidJ
kabY0NYMOw99IuEyMRTVq0xU3dnLvK3bS8RYtzG8TvsEVwWCkL0WS0ImRm2wlnid0GOQjmZPEIpE
cKHIOsUOKG11yT8VCV5zBR0V3pKBuEXvk1kMiPIFj4K2HyCGekThfBkcCsZspa9y2xaG8r4W4BYB
Bw47bSV6ENUaCYXSRkQq7Zkh0chEOcBbPQm49eTPjt+wu4zhMmzy73PtOVKgds7iwnZRriy2R0Zc
I0ZG2TTN5tYSWnsWhAKpiDoPL9qpKWzb1K4ij0Qo0gbtAo2pDRy5kFY1ECy6Y2bRFzbWcK2el3hc
BFWC4/vIFkge+IeWutfQBEkGpBWf+w68zt1tHddVQjwbFND4VAf8HbIwPvX7p1lU1++gzfFjEIOB
gucYmO7sHNs6a5YYMs89W9DZ6U9uun4rbpkdFI6uM8ZXSMQywgeC3vf/u0aExqcao8YUmhoiybmq
XclJijPxYU80fAwFoEias4J533bIJ2omDFkxhRjq4Ar4vKPlsd5Hj7jg7zBsTa35+eKilSh/28+g
lYMSeGBY3KGntvhVwlriy04HS4VhIgq+tW3O1gIjCLjWdYJQ7wUm3HGCRu037z3ASuSrqvbGYd0I
FB4B1JGEMh9x3NfVvyKTB2Q1F/a7FFiFI8ojK1GMFr4H0EUaRF9Nu92NO9PTo6/a9elnPwpE77f2
3D/jRcnQmWMMDwQ0NxGbajXcG+ZlgV1HmXjJKviZXjNYG5JO5LaHydmztcIg2Bmsy1qrhLH+4z5j
uSh5ZEsUuWFdqC0iTzXALHIQ0s8qg9mR6XZ4bHChxmzj8sd5Biux0riD6HnFLB2Nq5ibMSukLUlc
QILg8gTHACTxLFywcOeOsDcc8fzxZq87Dnku4j9PKqh9ZQ/PBZyeVB8ZeDwnZChMpgJmbHDNOouE
x8zNgRuLvuz6PJKdH8XxNo8h+QFSl5m7tn0AF4llrQB80h1x5R2zmSDDR5JGZyiaWPKQqpqpU7bD
MPebtxD92rAO2aSiO+879E1zWkh6N39ekITkZZZPWXwrBkJTQ1NIKfLCf1ysSvkVaI5z2Yl2pTWj
EoKDtwki0hJsTPYjsiu1qSPfVFb4hT2OlL8RssK3NLoGNfvTnoNlKGPCwNg52RH0at2mXH51/9G6
52oyvBGwD2Fa+1pU+tji6LoIOQQ5jAz09++phRd07dBE0k70JVU9olsstoWegttCCynJQUrRAiOq
E+wJSFlmgzbUEGIdnmkuaJ55HbI+PP/YfR87JiNggmD3ArePuxyhFZcVOgszp+VxVmUUPEjybVwM
AGdlSOffYoEJ+GlvFAPfw+X61/JbqDIiYB2x49R1rqVRSjfk5/GAz6fr4FZFeQNrX5L0wADk7j6V
apgZE8F7uT41OOvh2dELlUYdCteHU0KY7cogaayl8obEufS7AA7dF1x2a/b9KbpZ472W/vIK5KE4
KnepR6xWiMl8yVRbZoJpY6X3E6ng1KTx0kp3Cavq+ooUGnI0bjKZnYkDIEF+d2C1/6YsLiwSJWsq
CRU8E9i2gWpVj7X51KLIyoDrTO6DDRJVHgzo1YwS7EMqhZl3B44PHSoKnbkfm9ePZB6RBB5SpBXQ
ElQTmhQrmowukB9AX/mijwT0D0+Z4+YetOcmhPykdZ++Lp/eFbg8E6fJGqHQ6qRlSe3sIGOcOHlj
ZAGZxMYAGjzZ/ZAK6K6hMcxv8j1RxH9h5WvfwuaB2U+z6IUbcDOBFKw+ADPfBJGY7MgHz7/7f7SS
mOT4HcsL0PZpQCd88oONysw67YtkL5WWWYaaj811We48vJGYZMG8xCcLMg53m9ZC4Cb4cbbV2mY2
o/i3orKuybRQpO1lVTQbTpb1HxRr40uCutvjyDnMEl5/J6OGC/oECqxo2aqlxbJ/5dXoeocp0boE
eijI8aR1ktVXaQtMD0MPIeBNhOrpctQVMMMebP56gFvL0q9LLo5tpHHJSZQjOhJB281o+TzLJhRU
aNq/E/R+9s+IiEGeQX6HjIhjxztJxFPbEiimr16kjI5LN13M4YzdoTENcSpD281Hj6EMaoQn2vn4
S9ME+13Yh9p+mJZDO9VrD4aSguGWfi8xP/HpgMxfaYht31t4SndtH1so0ai2i0X8EMvMGoo3efvG
+gNwVHWmq3ibkAE7KYCkJC6hMtor1WigD2i5DbaeCCXl0Tz1Py5hYkvp2Kb0CP+WW1h4IpxlC/8d
UTGra0P2+evlsWun2ZLKjvU4dWxkpsDR2JMqWBaVIbJINCjwB85fnjfix/6BBLBt9GXW91Fe7D8H
fLm4vzDduRKlz82dDONuMq31vvopfa+dTCPQy/xXvmXddGPys+cMcnf+QoaaQgXGff6rzQRtgdt/
6Z7NkuON11tNIPBE0gh4aRnhfroZHSd0HBlkLMKfx7SCvTFCVnT72YRegz+7Gtlrk2kDphVpEUMP
ltqal5DxbZSWMpTaEgB/HmtsrPONqJT2d0YV5YLT2IpfoQ1LlrQ6ZwDrJPdQZUwtNoT2nwCfkFB9
RVwSkAF5idQtct1mBeZUA6cjaDhdvC1xwPMZT3GJ5NNH7RboeWBXUhUcQ16p5M8aFu0g2Q6ia0DH
RK3PDgdAIESAGiC/WPDOerH5Ertc9ugRg8G8x0aYHm3qhma3lten4jI0svJEQYn7ZY9MTbNWnSJg
y5bIPZeJDTYUGNo8HRVd9bIuhYN4UUfGq+hO1OtFM7xRRsrEN2LexoFBFtTXqGccZLYcF7tacKPE
KBnWVVR63jkvNPxc0v7TSErAuc54c5kgfzohi1DIiT/CDKPYhuMhL0XSvNsKm7HEkHlCJPr5Wfke
9h+1KsjyNbSrh6jLMRvlHV2Do2Ac7aziW7g8RFE8lWbj2wznnWoA2Uq9U1WP33lGkgGDnyTPXCBU
xxXuKbkS4843N8bi6F3WBQi819WeNNNpzAokzAnj1RaA2bxhF4RmTP/+R2DKSma/Z4MRqC9KHqKU
4c+7iXisx/WVynIz2Qpnpc7VRExISiix07JPh9POB7Qq5G02mkGVdCocsqSoc9vwg23zuoxIMQGS
O+DEHmvO2ybMoMu7UNkim+B2DG+bHvzywbY4Vv3P7dwRzeD6XZQLdj4MM/pY2SCh0bTEYGVJjhZe
YcW4XQVUmrcL
`protect end_protected
