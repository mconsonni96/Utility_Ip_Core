`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
mZ3O9q2JUMfAXl2Q/tfaUkCXOAU5/mXfqxB7mf8tyeGjg5GWhLyvyqxgZ/NW2bNnoAmTEXn74G4O
2nlDOtjMtgBizUzbn3apOFj/Q/zdoDL+7jrD2F8vM4ur4YFInxKIs9zh9HX3QthKZo7skWkhrFjP
AH9LO7qTXE2WetFO8lEsOuDzCt2TfF8ekeQ/CCxfcBmqsvhIXrNhENxsFlqwIq0rGlpHxIYEAK+U
ht9FC/B/AALTJmFzonmLpmP0gO/ua5qaySCULH8KqyF4Fzu7G/C9FUl3670VNEZnZ23AVwDez97r
TYrFNhnANAS6kfUNIdzWLxo0D1ezSSEBT5llng==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="XqDpdysxbvcZmxbrRltgj+Bpj6p8DIR61YH2Tp7kWh4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14640)
`protect data_block
C6ewaQwOHqmWoW3nFIzn8yEF3hRWY59Rq17H2bW8J6L1DKNS4VCMv7caKdWV6XnRhYuunD8o63n2
5m1q+RyIhG+DMtGO66Hxaw4dl3lzYnCB+3ovzCfApi52AlAE99JHpkQyNEt2POYS7DG0+1hgw5lw
CEBUtWwKJYQ1F/BNSg56bQt/mV6vZHvojVf4tqAf7m4NFT5pzWcnmctx5/6tLoVzUzdyqUhNxYXm
Af/P4KAS7vcznFXqp9/PhlPVPUzkec+MG5lWMT0UOyeIF1C8KqQpL3kNkm9vaTdTl7IslvIxLm7w
D0ISfBiqI4LBSPIcDYG8ffM2inMVZOUzvdLe7HTQcCSZ3YgOgUU+zULhek8I0ePqJbU64Q1YFitY
CFqZCEWjRV3bad7yKyRd/HMQnSzyEdP09RBKbzFgXBn0+G4UgPVkbMcX0zrQMWdob3sSCbea3jH+
0w5urng/VZ9Em+YikLK2kyhxLfO/zpKO0kRlC+nNkvY4ljOS5R4S9dHovfFGUa/kzxOY+6/M8Z3D
oToE3IGnPzkY6pedpGK4v31YNW2W7NqnuB3jpIo3FH1Pb3e4QSZPUb19noEJIkGbV06Yj8egaDot
lneKkH1auy7bxNNz/IjltERA2L2U2iJ3/fYH0BD6fA/Pv7R9kArxY1x86Yb3dbe0pq4QihVs4suV
3Xe3yqcE3y8jiYlXNCC+xAdZMRYWXPVbLuw1mWKPTmINX2UjpUhw0O29Lz4MhP9D5+MDymAsSX55
dVI+UXxWONLNxXrnnSA//B3QbyXEjn0sz9213oI7UHvdn1YYfQbcEjJcKUPC3VNSMwj6cV2nB/L/
H0a3qVZPCKqe1l9K54PmjmCY7KycmR+aY/gXLL56FL9URw/EPOfi8udx3CZ8RKgura/vM4Mh0rtZ
D8LpFxh/+uT7vauBTwscOCayea4NAvxXeeaymS6EA6rwTM2TruN+tLAt49Mi8J72VZiahWCX0UZ+
dZ3dR/aJvof0I5F4wRqCjL5DID/UUjC8k5QpHnxYrYfY7SWl0h9LwROqWRpT+hyMw6bo3xb6JMUM
04Lgu6cOesx2GWldeLBQWrQYlAehl6JnTDGpREACJV8K2KtO+Qt6JpCN4e7Mbv5pm+rv/LpjL9/K
0T4OruggD0CqjKDWZDLFUpompvHo4GGWdwmfmLrjtqlHoejRAhcv/PHmGDZTULho6x00fL6dsBK8
H596RdjSOuxgmkQy2xGLn1bxjhDtAC6TGS0BYtR0kc5FbcZWemgNHIYF78x2GAGTlE7Ux8W1CGyF
S7Ex0TlP4wQR8tawSOFO3Aw+NQEGhtGuVSD9Pw63lj5NhPpQujMer4mqPLTgrzBW1gTRZgAh9T6B
lHRVnX59bIY0ETGQcfRWWMT62RHqunzCfXUXadgWKkDjGJOajlEwqQYBv55+CQpb6XCkE3Pi6q6N
XMyCBiSoUsAAJzg+euaEdE3uwpnKbK/JKtS9izBmlBSi1wf2+OVfvHkKxGoYTtg+hc9mdoVFmDJC
QAsdlfrc+5EJYcZaPw2uu2pqlv5ur4tfH4qYGnJDTDQypA9Mo6flCSLsLIncj0tOnANU515K7E7H
IM0JO28k8FCwzoQgZn/k7a7epYVV4Noj+TVTgeYpRQ7/RLr2gxiQIztUheOh95IFpdfv0xOjx4uP
Ip1jk3wtRKpRtzYcxFhuVYFIVylbXyh4L20kRWe/5HdTfQHPfIda56GyKvFKbtilbzeAI2Timr3A
ZymB3elSNb0sfUdJP46JuAgPPI9FrK/zNiMiU9WyiO6S7nxYsnFU3hg+z0v9gfAp/obAs4foDag2
8GS5f3KPrbc9EkAN8AiilB1xEOGAd0332RQvMHRprF1lhMMkmSG8MpjWsW2lVZ6gWvCWnpk82buL
VEreqKpiFrTUIFkvlv0E6172kQxDRm+YRnpHxR+C5SK97i6l59wLCVATjVfCKg0YPBax5nxd9/xF
j1sBJqQi1TTFZhNjstuhXc8JuxeFikHuUyKXWvOUznR9z31+/GGYUte2I4B3VE7lFphq5XPpch2R
yu5B3xWt7tpQoN9z99DqiF423D4IDgcIUgXS0gZrhHVXX61DB7/Vex/a7Ux/IoOD2pCN2F14MypB
kMHAwrsT/wF4P6bAaZOAQMBe/quTdX1tJzMk4j36p+SDwaTgWUtJtQnzvsvrRo1zF45LqDCw2rf3
dwIMzwRPfh6oaBCjF+iwPY1myLEoMuUZavWXelQrI3zY1brX14QvjPt83/+X/lElEgLNKLH+aR77
chAWniiwa8xI/LrQHEoBXBOa5/Ua3MAEawpZ8xS3DdU56/SZk7x74oB6Iwvuagrwr7v7nWgyi8SG
/xb2YDEtl9vk1ODxpehIrxUwpWBBrAE3tXw/Dcbqx5T6NHrydO8zbxDfo54TM3DiakgvJfgOmDSB
Uw5fTsRSTtk4/QgUa3RC5e4QDO1Zf9B0KJgrRnCo8tsBKJ93xlxS5ZlchAAbh6jTn92NmAUgyS9S
kVz7yZzYV4zwrtqEXxUq2tvTu1s50SrPXAsIp+UynquvxH6f0cRwiQO4IlwcR4aRaOtnYf4mSL+V
1EmdwKDLVkGPNBU9E+IGoFM3kCsTmJQjYvzkwusgo+mdHo7nljOIifsycbIRhXdMq06r8g1bo9nj
D3DGrWBa6JUEqoR3NzNSQPtjGTKFcjW7lMUS7PL/XBv7rn8CidX9KLXlxotTkGnmXSKti58cJDDr
x5MNT9V4XecqG8xWb84VfkAvywBmiWbCaO9B/IlDQ4kiydkfqVLHplgvWw2t0v8eST/kj+15V7xi
yDrkcR9HPtd8KahgUiFeOogQyeVD4ziuIpY0XsIK4N+vRkNe4jPqT7hO8aAXKX2Wtz4D7b8cN9IJ
vyvW0WrkIiT79qB/ICvboGdGDunYNegQxucoQZFOxpQ8qUOztBXD3YNLvUmSteCoa3+vjVxV/zLe
t7pgb0lKdV33U3sHUScLfod+5wMODia1dBjHDrQIhVywpSjEAuc++JiMFGoN7eIogknFURz4ggFk
HmkiV2LQCSRlnJ+V27AmwhQQCqmeRL2naijAw6KPY/XiaSNErQURynLDDf01OyXhB7dfVl7WLK+7
5B27n4gjBcPnh6xMQRCHiwZ79k1yYphwlUEtYoDjybQDgKQWd+CcYG7Rw3JNSmbaoi0vZbmAkZJ4
Vn2Asb1BjU2Kn6ci5bcKxQWM3utjgqUEWvH33s+WBzruiwRCvhTHuDUpWnB8pHqt9PeHeFRvpoPL
mE1HmN9WMUuYrXGMVilfmW4/YVWCVAFhX0SO5nlqXcPXoBDbzC1/5r3LYFcwqWYZNVbZgVGh/5dp
G8n4EO9FWAqWwgiiPUJiwYUr7KIMeVHmML0NzCbbAKca+XQwXClQT4r2MseNZzl5U6wO6opVsL1X
+DRYQfQYfW11P2+jgR5qshb92N/K5Zqedy2Df0R/azcxtgCOyY4JuncDRoVZt8r3Qf1Zv23dHGD5
kNif1blPF/5KlBYfggavTrb6zcbSKC11WKNw64B4ickR78V+3oTLYeUGlyLpocUsWCoCVoLS2iyl
+Xq8Jw3TSk1HPGohD9lCHAebH905ri0ilCSePDD9GSy0i8mPDRL8lwqyrFwjlt4aPAL4IHO9P0nz
mMb0E/UUSd8qajObjkm029kNSQXEyblFLsrYPxiiWnSAa7EEngBu6XQMgNB89p5lw6fUDwS4lJ0a
lrUNJnQuBluqRAXLdqvt//m81P8U4UnpSUSfAVb4EO4yBrDppgjYQJZmC5c4t5uLON1rXm44DAmU
SpeoRCtaJsdQbiT/PI5J4d7u8A9RBAxMbwVcF8eXhDFLO9OBDnakTTY8K1jJ95oAfTpm0NTVG6JN
uhmfNAeMG9WgFcdt7z6IMpg0EKqE4GTgWzeSTyVFDLjt/QmJS7BVSZ53dmu3X+RSRpy24hoZEhu3
PLQ8Z2gNs9hvkWf0xLqqWRq1pQJ7q6rV7CZBrRH576DoUgQYJluGPZHzDTSS/KrBISVu3+UrXeW2
zFcH7VfyZegfaP5R/QLRa1gcxLHJocrQ/NTc2217Vx75Hc7bbNvpUbpigf/moCEKQiu2AJqyADve
tElGqtXKn9f8zWwG5rIbOiOJzTxHhgkEGb6wGh71G8UYgoDUj2wuyLl+9TyZ4e8G/mrQdispudeA
8iul2gPRZoaHr/3SfyMoWfFuisY9lF+NeIFV4ret7U1dZJW2C6TG66xR/HE8keDZYau4vgdts8vV
A9cPhCLffaoSVSY5nt4bjg6/gFKeCuqHg5tvm858TVXP7/A7M/r2QlXoHmrqnc9NJVaYlDY9Kf13
iOQlJ02gNsBPPu/l9X4oCYxyDx21+oDEsLwkIJalWyPav1PgAaum8j4TEZbpP3tWSMeFBm1cWJXs
zSg7GjuozqYbSXj7QesCWj1b31Sa1q6swhiyZ25cK2NxxQ7nHW/eMX8YT3yOIEEsvfnq7pmVZJDN
x7VadOVX13BaxF81ueqWj8TgEq0wJblgK83Ky1avKCOPUPuIImrSS0eAJDoIa83j+TYt6XnaB5q0
FsRd8a8NgAUtLI7OMXOd54GfujqML/fGZEL9mdK3k8cENzYZH3WAbUoNm9TDbfD3v+l7jiKySVkZ
JSUNpLX4gaSTZX9WU46p0IPNSEh7yuDMTsHesrlenqqvQ/hN3vZaxMltSv61In0MBJsvVxzQdWgL
QUbaOPoI3RG0aEXpBPfaKXRlA9PZUjHlzpcq0eGFucZH+apYXu71EkfmHV1FfXSlAKG6DzbD42A/
TzAlDdfBARyYXOg1aHtVvo80+dIbpZHL7g9zfO3ZGIi8kZKBHsSLuOXITpT1a8lVDG/Z6lCJv9wA
r7eZcTpUncG/wivAPYZBNBxSAAHO1e7g4XbdVoLq/uu9gYOciD3M35iERDl0OU8MgV+ypkxg0K5A
0+PdHI1bkHtH/DNcvEMNZs/UvWs2TzW1ntWBaDWcMF1NIs5NAsr5KhVUzuJvFGjdfrm0RUzoWoV7
7V5tcPmrLGSRmWED72HcnIat9sQQc3/JRzRiCA3UfNIGLPnhXhBFl+E5iroiZSsITQmctrpAHfta
BS7k+AebORTrpMshyWlpaNMRB+moug/0SBj83FqX8N/cVvj1D8bg0mePXAyo/YnuLc7SeZvCwMcB
R7EnJXF2hUrUO2POR4ZmhykiJq4u3UXLYb2wNEqEBgjlpKV1Hl2mwYrpQb5UGadadh24taernoL7
2AKbTwrq1odSa1SSwn1bqOxEz0+y3ahBkqEiGEdwz7c0r7vA4Z+XMlRs/a2vh40pJ44EKX+w3nVN
adsiucNbpaLqNeCJPrAwzcSaderPNDOV0ZErWq2F73575+JSXiqfNcjEZPogAajs2wX/a4hxZzXM
1soBCR+GxCT5vfdfQKp/CsA745u4sByOe7BtzaqC8rO2bWylKPFor0gfK76fcvFrJPT/lfFgPCET
SuDKRVQmvmEkd9gxPxVeyDSxFRZMfrVCprbmK80wHcIrWMBLlaL/ws0FZrqfqRt5wBv4pZ+QFTHz
Ob9UWYv4kzhF15pBvFHJAkEkHR6zFpT8VOROJcIzyZoiatnQ1IfUNtm1UvOVwZxae6EfLxb7YCKw
kRfSb9DsDV8WVyDkrq8Qz7da+lzmJIMVjLhnrxxuJ2D2TZVlFo2jfiGpIlG7wFTQ09swGxIfjPSG
kQ3xUrboU35FhA/2gGg/DsBg8NeYYKcvhYBA5AoB+lzllZdcv0lMs2vz+I0cidFCde5wjQ7EHY1i
BY7kTn5vRf/TlYNzCgClZNksOoUzXj/WGrIpPE1RWKopB0YHdUxIFEsCmfuBWB+a9Ym0nYvdhp6r
RpvrJTmiF0yo22xRPJ5Msyk8ykDRTEvbe7gHi+4t3DgEDQRoR+Ww9cz3dEDq8lV+56svZ7UHVHII
5T5+imNG9gdbYHJtwJIK76bS/ELgZrlPmzbRHT0Wg4HCCVJMwMqLbXqHuKXMMBCRJllXCQRDCuek
N8tW6vrSs4oSzZ/d03McqIdjXWfP1Jq041i80GLhJaOuSbEWm+dgGpocm76yVD9XmmN6afuOrJ99
mdlx2yJDpkQ+NYjUggHy5xi0FIpp3J4DvYP39vrThBTXdmZ4wlLRFQtb/3fBRq4q1X+GcddotGue
9mvTZbj/683gzaFO3si2WCOpb+MY39ZTuCfYHZCeGSLlFb6/Sa/jQsvezSB5LAJfR3okCTG6MXFx
hFPWq3TK/3iTUhMHqEnvpnP6rmsAWkE0rOce9XRNIupsWNwYXWrKjpk/4gDKIv7biZH/3uYZnm3J
aO6mZEevn5WngxZh6F1qReM2ifbbG1YX2hjjXc/2mKjz1Lr1W4FzRNOFPnta/d2JFgjd3b2qcMTK
1IED5VYowfv84LSxou808/06YHxmADGNHLWKL7RwGmp8lLra09/YdUaE7koxWJak1WILP/tvrn4B
+pMrCm1zgIlyJlrrpvIYjg7uscfesnSD6cTM7QbmBUlC9vlH3GYRmysO3gDKPhX0ZUWPUrbdERBj
tKwelz0gRx3KXH8JYc4ncOy/R01F0ka1+68DY6WsCalrmNltV8ENeqqIBUUlxCmjtWT7nfzR7xZ4
Jb+CY8B6u5dtHRoIxdAEKftmXWfXj6ONd1D2pq95rQdRbGBPTdwxtkUsxgL36DZ4MUMTqUXPw8KP
9ZMDsKADHvrGd8n3sgfG5rlCWLm2yk3Rc1+7/suIrb3voqm0ThXIHRLq+/mjjgx4OZqRLHlz99Br
ePlFY1raRSTfRATuzgZeQ2fbpAzieD9HRpXt2YOPQz09QRkAeKMtvjAfOu6GxQC8R3AsPdVlC8/V
hCF1nFrNbT5ZOqC/XL6QkQm+MkhU08FbOMsBLpTAn91Wdbw/3X/Xux5tszlJmRDYsOFi6y2fpaxw
HMw/5y+FO35i+334NPzydX22423T1MjpMXGu1ce0JlXNkOjA/2igLudvrVeGdgfZg4Ov/C4SJC5w
rJxmVKnAE7IZyF3HcRidjgBQEOep+lGHKwv0mZZQsLMfIYYgU054vJLaGKtZZxxMgj99jJ+YLGw/
wcyT0anliINlg/QvG2+TS1b1jjMjZ0ZrJVT/hReOv+HdmCGx9oUmScuCWNSXpmKDyGn5PV/CAX6A
jFvAlO7D04ZUbVWkiq71tll0Xc6i6rWvUsxs6seEq0Bn0kem71OQ+Mc8bCiK1hW1cwhz8ff8TUpV
cO4nYmGdVUlxuWKDFzfveXsF8PRjkSP3WBC/zuT0sxpQfNF2A70wH4AHojMmq1ahEjrlZPU1kIda
loOTOgVaTze7c8KGEjS0B4ulQuk0GyKGp5EDIsmzaRnCrnwhHIR7T6it0S/RdA+GVFqgMc7nprpj
c1weJJUfFo2CaCRdWibKl5qRbXhpAfBfW/6DbaD8sPxxycL8cagw78C4aF2mYb0Jb4CkfQcrLJov
ELuk3gPqeYOpxaZPqiYExolXM9V0xdoj6Yq0gW7qorR95s5yW8vucdaFZzdltqzYqSL11wRyAd7i
+YmHKy75WDY5VgYAMHkQCxfIRUPXH68EloY4eG2kKTir59cF/HG3bYANJKQ+5KSF0KxJp81ZfkMM
U25uWAC4/dpyMGLLa4XVXYeN5qmME+uqj2n/0efdfio4J57nO29h4xffY+I457bbhMAJUpy54fYA
nFfKJWF8Jjl+dvM+fs1mUooJ3qovi1qFVnksQuZ28675/ogIsidt2YVU69BRaZS6uo0uUZiIl3Zl
mkbTgEGC6BMv3mon2penZUpy/Ttc+XMsDNtS1ZZa7pe3pBfs5mjvrgETy1pN+Sz/4Aplyi3MnPQO
ZNOEAZg7vXWUP9PCFdDomVF5CWK0GmFauLb9OMh2VNKTbohpQiYr6QcQoT4KlTWv/XXML0BW6vja
DJ9vi6Xq5rlZkkzaw2P8tRYOuo9f7VedGFe1lj6P7VU2YmltLrk8u2QtE7N7rZ1iHWSp6LdFmBEB
U1J4ra1CN2gQrmJijv4C77NFzdxH1JBdldCJ+UUGIW1nBSZASzvRaUSSnfe3Trx1ZF4xNmyuA/u8
tVkZF8imf2R1VZl9r/lBGQlvTDcFfE37hCwIks2E8Owku9T8TIQpWIL8iCwIPdW2yF8we+pqEiU6
LKy0mZ8DqQ0JAmgDwedvXwybIb5PnNGk3a+ulpeItM8WEVSUd8nES980HUjU4RCPbv0v0UEu+I0y
WlvWnJbjW4vCW3urK6LeVlTMwAvJoiZ1v2wNQqeyxznQN0kXAj6o8S3P09P+wVpoILZ1ntYMlkHz
pnyvEoDyFmU1lOZDeXVum8YBDytNxJ4O986rZ+LRR0l/FSyMGEfUnjUq8M7psc1NzPMpPsS7//tS
xefUphXrHvrMQ7cJ3Um7IxKqnHB19dVlpTa2Chg2us6gQuPI7ye1yVjE8NTbY9j48HlK4+60216n
T4xKmKNH7qsRxIXMVChk3M5FkHA+0g7Fn9CJ+ggjLDvO4b8gHO8etlVR4hq5QPMTkh8A75Zmx59t
2FA6OXJdaybbDKU5azXFJuqRxbXuXX1sHK5ZTYg4jTx/bjwFIahZmPg9GQ8I8sEkPGoCeHgxUwBP
YV1o0xUKazAyajBhd58q34EEt+9Cd1TnAIkmbvOPuNjP7QYkEzyJTMxcqGjS0+cIlMEzPXHBdf4o
ykpLV6l/oahsSTE47eMuvowAsBP0M35Jf+ISLhBWkyyLJ49fRDbjD1vLZTkWXKgVRA69sVO+Ivwc
CJVA86SEHbY9MoK3WtmfzHXS7FkLVF2mzqGnkgz1/JjJKk2NKFH5tpJZKiFAc64uTv4Caji7OnFS
CAzYib0fao+eZwh0oEroBJ/anCjQc1iTUveokju/e0mfKOqoGUEjRp/HsTPUByhTL14fbNnjgVqV
sznBIDVgQ4M8N5OnZnLXczMQGsTEskFr/bU6WLMfxujTV/loXgMjU2e4Qh54e3yrD2w/r1W5bKMO
FeB6ghf12Z6mQmdSsvpNc+ly1QpRDMt7gqzfMpGuwLlnoRYGvimc8268a2H2RkMC00uVUsLtFx0U
JEWaIOUnPfghhxrNwP/ZrnWYHCJ82ROXZcOwolpV6+wkYsompt/bEszxrmrNM7aBR2sfPmZnrMib
4qQayoLXdJOBi2usZN1V+njcGs3AeHB0U8i1k8tJouDFhsl1zMN4WVGsKfDsi5iVgLCkWg+auh2E
D0awfDR+/JjOaF9bRm39/1dCh6grQg1meWD4qXBumHbBj9FDkuORLlF4qSlI4DUPurUAdRnEmvue
3oFhBtUwGJJZXHU1ueMzfxSiWdY2KqO87cLVvnbUH6M5ILP1iSUWq+6jlbAXRpel2wngZ/Ik0TpW
JUxNkTlwrqIEu0LKwFZD5yHOYMVjSdBOPLWDu4HXTCE6hdC5mANb3XlyPEVZZ1g3V6mRX5HSwe2L
FhJolTxZL1WfmJ+WTl14gChP7/OclPDamUdlCycS5Nf0wIXEMoH/3qX9zGuam5PsBHjTm4qScROu
FZ0Z8Q5SHEvnmAKvpzbVYYpDtgjkjrRHT+KiVaRbFJxTVDCMFCg0fSLtoKKznndHDnyV5zLGk2mS
h15+6r46JsIrAROZgfrYEuGfKlrw6gmuFjLXO44S9lIPSFlmOccG/vdcaL2lbJF+ZPivbIWkwrII
D02qnQWMN+KBy++LnqvJgeVCe2g9XmN1DnqXj9AbDLrjv5q06ocQBUPRpgaBMrrTUW6ujkWvp6AD
nE6Z+RF9YMVpbN2Ur8AXKbkANBTMuz5WJdDGbvPeU7pLYwBIscGzkK/f3Xio82UxMYwPqHYMwxZq
pYfqPrvUFwYk1rokloAj+WNfOd0xZaetgGsh3C3ObxW5O0VVAeEpXXh+Q/LntTRCvEwKo/ZLg7fA
nm6JVckZjfefL/JDZwuWhLyzkuS8uEpcfaU9i9f3aYHXpLwAq7DIClU3GKyBUa5VjIFDY271AMin
IWqNqXmBDEg9ImUaEBrURt10fpQtVh//Qh3cCTya2IfWPvEGzryhE9J2/nB3x7LqEVqXDpPlEciS
jVCJnFSYV0DghUEZ55OwjKs02sqAmTJAowNmaMW5vzTTTt6D5ZxZWkYIh84pmQ0ph1sUcHWqG05/
xYy4CJwCuBO2lLcqsLbr+tFox9S1VZsmoLzgDZ+7qeZBoHf9DGnhsfpFdDdjw5Glkgqn6K3zLvn1
N1mY8aA0+CyfC6DH/hW31Tt/jxDZPYxjDDTbDb2AN5c8rPPrZCWaK1JNU4Yby98PWI/u1D5Ha/V1
H0i9x1WE73KOrvzSR78N5HQFU20ACuYgyi55wcD3UQU/pNDmw+m+BRDPGX/4MucPkDyx5n14rR9Y
G2aEjgHNZMVGM3irRp+T8YW0LUQtcYWdYRVJjRT0P6LkX/Es9Il9NFxNVlfXGBoHz7QCnDQoKUx+
UAWVLr9Xd6rPgYb+T7u4on20MxuiVJKokp6YoBhZSxXUHhWimnDcqggdXoC2Qw3UW2hqvQsqH+sg
H1b0euW6LXkuT62Hi0ULDxV/dYQP4Bm4Hpx8CcGzigRP81rq74O3xHKNwg3Xc1k/eXlIORr6NuYI
c9Uk7IkIpnaiCVnsgRwkBO4xs9S1l1A7ZV7mX5aHOtdWfumSpYja+f8tNKN/zJvn3Z8LU3dS+yXZ
BrxqJ7XRLg78VdcNS38IPhbyYEDXpGZRCXfezgRnhIhR2gwKBte7S00w/hCOMS/UGIrRUpQ0FATU
3bHM7LEJGxGglQRgWODp2Hs/SNPTEsJxJ5WUfTHukvL2sn92Ajunzb/qe+z7uxSqexkZhKVI0qja
KeQWb3+GPTaC/j2oZvFXj55l+AByjJoI9pjP8xF+jov77ime3uj2aH0mBUKR/HMka9V02CTTLAjn
Ao7PIcR2ZZict0LH57DLqUQVAf5kseojr/+wrtriZXcMjvOL6RRvFZ+mz+GdGVIf2cIzNHOqkAxE
qDYWmSe6W7Se+vXimOeV5oq3lPd/nkbVS+/g3HI57IU1b1xnajcmycTWS1I8o554t6tYG4RO6vnb
7tgII4cmflspY9ZLaQ0Sun3Diml2Sd6IFfuvEVi3pnC3trZ2ICrWV7StpoJF0TIffqXgdCl9epDs
D2zABK0ABR6b+Z4wikU7stN8CjoYSvHTWjNeiWdeOEorl+bAlmCAIo+bK6jOPlu9d6RevWFJYspS
4jh9AYnZb1KI23XUI0529xLB0LV0uBnN64PVaxqLdVMa6bS2y0IDsIP1JRknx5QsOXSd85Tlz9pe
R1CD5tAz9O/KnJuqJuotUP35G7HwbikVMxSyl09U+MZ142g7ELx9IAHIf00257iKYw8SNcvdG0hc
JoVDhptdd8XgRtpWp/SE9cfxazUsi6BqPx6Cjuwec8M9zeOsHKRb3rx6INoDqxBYnaJMl9PDk1gp
RbQdpTQ7A7DO3cHpwnXsDMIT0NyhANMvJmu1lYuuEvk4BYth7gpywJf+139AqC9S+/bDDk7O+SZ2
nF4jpsWNpv4Tmlbal8mA1wXKS8uGc0i/5/kcwJ1nX8HPZfYl8RTKo5qFqPg3JHCfm2/hP4uYYygP
e/5Sm1t96xQ2GU8DaofiTSHL2S/spn1wqYk5kj1p+nZ+00Zmg90fFq6BaTJXeLomuJIWur+691HG
FW6hJd6eAxYKwPzCykYopXF8rXbzlCFXAxBeL05ztC6QlyUgd4K7zUodG7dVnj5tFoM9hrZ76GLy
qCUnc/lcdQoGGGNU4KM5mNBS9ARmsiJKC2AQYdsbeCY5DiyILGH+Bs8BwN/I+xU4VKVT0V6lA/Mz
Ot98Ow/H9UVZUQRT0Wi8DpvkJ5uIrkBeJ0FdQAdIhcGitpsQkKcQBs+LeGoTzhy+Rc5OiY6keEZy
eH7N5eJKGGEiqIDe8yBAa4MZ5g0Ehm3fqblAr3rYxAHG7g+TAZrvGOuxz+rk6PanESOViuUvzGnS
/YTR1qEbxzwL4zptwCLW5k/w0zafUpKwWa3s/8uCrENnqYBNUjIJoiJB/m2Vss2HtMQJ6/2Ek4oA
hBd6JBZcqZdlcNpIiP9Uks4H3tc7aQ/iOJEQa7c4rsGgEJ/i9MzVyICFI67NbTUuTmByHJRq1L3n
hAk3yqHnzc4BfEArZgcroamuYkUm/F+jkBXOahD2eXgROW/3Y66slqRNxWiQ+9DA2IxKfyZminx0
nAcno31CC45JRxEA07qTzTf1scDSF3VGUCuxGBhgYc+3T2lxl/Mdx8cp+7yO7vyo0lda7359u0rI
nG9LFxZ81ZDyCSq62WF2K8XydDdM17hlCubMrXraH32toCuyA53uLtSskRcvWL09/uCqkRnxEom3
iuRlsbsX1vPVFdH1JVlBhITjOBG/ANUAbRpS8J4Uk4jghPyuiM8QSmCYVJ7zB1cduxqqM1WWCXue
dB1r2Rmux6GEgGaGJW7x41ZJCY3QE7I8rSrDWhZsZAEsuTuwi7VuYsb89Zl+NDT8KcOnaKkWm3fy
S8g928MBPf0ZdbUNP/PhXpoq6p7locsmiyGSy1W/j1akL6Hc5Zz7QTGObfySbQ+tKm+vwoeJ2Q5I
KVliXZwXSB8U0mkK+wUtt7pbv1iSFbGOcXtkAKbkOZHVGeMxjZNbCbtD4LHqd4XU7U60tqKbtrVD
QNlVWlAEJjmgejFYHzzYxCv9Hhg0pVl5MZX1JWWyVUDz7bW0fx0pRFuf+iSccm3sp8i6bpl8rpRq
BGFhpF4IsL7n8yvYQkXD5LdpanxTfBGF+e0T9mB9293GvwBQU4mUD6rX56BAxor/bQ/fJD+4ZOHu
MBO7TV3Wxrs1WgDntqTrsYgb2ftkfxyeI67cmtAHDgAsNAXszHredd997XUjR3xXYa4hzWJ3NXxP
WeG92NgLebM0SSWBJG6oWTB+kNDLIkAdepsdH9dGaa22tzl2dJ8BFJOgDp789ww4CD754qP72fKq
ujZItqGA6h1mi4PyTy3CTRylzy5N4MCTyeeJK01gsiS36u0gNJQoXTkU2S+1gnop2A9J5Rkwg2bJ
5GLLMybgKnXZbw3I5LxuFpSXGwOGNJyy/DaIzjZSGGts+xl/zvB7R1oUN6dqbmW8TS6NLZQ88V8k
IqgBj57jjo5G2je0IcsFe/gSXCRV/9pd0i5R2reRVb/BhKF6SIRZheXBR/U5JM7SmXvOhAF+TETz
HT2Nxgm58q/jG/RTW0YgzDYu7o7c4HhKgYwBPK2l51F61il9MHQk9L/zxgr4eXXi+RI/KrXxtjl0
MafbprawqGr1df7moMN9iUjsYX4dXyVcNLCcmL+o4rawPOYyH/vTqwVW+rhgErBMjRdNCAFTPC6I
95ccPQX9bKe3i34U0PNCACudmPuQC5hLU/tSv+FTtplXyHTEdr193istdm7bjYUU42V5unu9+Nez
D/3uinooh3TeaYaDxSur7xIeeurV3pgAV0KICaesXPB9P2EpwGwO6t7kXWKRhoPje9f2UknYDvL8
T8pNRbCT2ymstBv2TcapqYk7JemplYpIWcf2HYXUQ/fIYCRydY0bZ5gYqnT+PpD1Pa1iVqMKyPc7
jatU0R9JkiAwnO48Htr0oNpZn3B/EVzQ1y9bGeKoqeE/GzJNdAaHonrapjZgUeSaPDGWj4g9Cd6h
rd/EeXznvErQVls3mi0OGZu07/+CPqMxY4nTMgkXR34Qq/kmp7VsIATtw26nwL/nFCDQ066s1DPg
9sZxFk8CaJdTDMO4NFpN6baa//o5ctfm1/pNweFhhRVJFw/j0qHdXqMLgi6QiI3UjPMkyQUr0M3R
GxTQlC01zVIvbcs9DM0hmfwNKoqX9/x6nD+YDxSjp/APNz99aFR/AJYwcnIbyiYe3PUKZMNQNXHB
t2Ik3fVnSb4aqhhKCptekAfscFioo/E66I2HPuwoudbcNorcueBzG4aDSOaBqCc/BQJf4DmcIf8C
qvn6BQGMas5Z5rnKs1/cXoBDP0F2R2+pdKeXukuEnN7+gsdIo7hm0t0dk8fj6W2y0o5LWpbzSSY0
cIMAlz403GMk8OdQ9xzqYwNQeulHbHE+etJ0rUcPdrBj7NQHsaN0X5oKCWLHKIqjg4AzeKmmg7UW
aYFnWX4kJaJFZl/1kSRAerSh7X6DHAjoW3DHjQnLSicTpgrB5daDEO8j6lxyQ2cNFb06EB0RwKjV
yoqEUgghItpLIiZJ/Zb0uLDrvem+6jaf9R29LexQ6uLY5jOiXtO4F17xZ70CG/jaFCoss/Om1Q+N
o4MsM6/0ZhPEjt7gGpgNqCq8bsG8baGvG9FJdYo860oidjaIZDftBkPh+w6BGyxgRIFsYPTT1WnZ
itNZZlH+aQQgaQ9G1y/vE5bgpJknCcUvwMTy1XplHD/uwxXLUxRZ0O3+zefjalttXWhU8sILB2RE
JBYXWm/InlYDnWBdD6QdfyoMm1ynZEchxxZRMKgemStqJJlIizD+RYGW5bGUMxykuqJXXOlbBPAG
v7raj5LwcRqjclFiFHqGCmbhH8FYF3BLho4ni0tWPRtqkyoA93DXg9n3sP+ZKI2BUMyLsFpjV9hh
MvthuXQj9n4CRlvvaNUXvPUYWAx3ZuCfg2yi4K8VFeSIA8KW0IBxY/raqpYienDEHzYFjEzMmwsl
KLjG3Uq2NBooDp0e4J+c2mlQSdceF5TN3+buBRYCtO/cFl3ZO2hERfftvh/07fA4i1GQHLb08elT
7YMkclpiFesrGNQmDs4EyTYBRpYuPixIpVAQiHMpn/Bkm51iW+DcgTKX5pDS3eJ1HbsK9H5t1vsV
39H64NpF5G+O1fNmTyL7QPlsWTK7xupva29jPo6m8Z8BQ865lHU0ueNkeRVBVAxyu+4OfPOq825R
jCq5oDNm7XUXqX2FD6cLa/MWcf7uAGcQnRVKXuJwPqrlwEe8bh+v/4YG5JjKj/wmcCUJwH2V3/GD
mOHJxueNk/R1w2tTkzZar1vm8zN1lV4TwnzdMyckuP3/fJqF/RsVg+bbPQVYCiF5c2X2AQiCwxi9
6Vfok2BklIcfmfA/4wb6e4Gu9IafgISFHlSmiBLL/92KxQIh6h+cQwwxc0ebKGiFGlL9TCZuDzHX
sZqdhPt8nRfaFwHY6OqRXGaDNCr6m89DiGCGKC1iNqrpQhFt1nAIFVsq86DCL1/UKqvYqZns1c5s
djsymdHrP+0Mnql88wNaeGT1MtrODwg7ruNCaRFz3R1B3+lsWeUO9MqAtVztnCzLYQtN4JHwd/iS
2LMdwMmY/GHeCxzLqkktm95ClAp+vRn1c6QiAfYwvJuxscFYSJA2KCcrz/9JcicduTggQPKIU2l9
9hunmCvd12tACBUX1A7ghwFRERt4vKbAGs0/ONdJ6DgYu9D5YEkvs07hw506OPBm7zYowsHSfZbT
uwlfKLCeji1HOavBnrWkaiPQ5dOGfrMBhO8z/CElUC1veZMw/5c1H/4nYWbGTb1YEtnJH9l3TweQ
XRgM0GD0DcOBK0irEHY6JMJy6MKjufQVtI8hiy5A7ibnnewhbUVEjVDr6OFZrz/h+7d5oVZqopMW
nDU8L55UTyrbmVoVEgLN6Fa5J2XX28aF9msXPndea6AUC23elZ/IhUQmwLkuCzF3Y8VcHn+gbnmT
Z2KWDycC4xzdhhRjAAYnctcv5aU9xjLtdm8iT0eRNTvoZ84Ae4Ftvf1LlU4vIBI1QB6pJt6+fmS/
hNp8GKf/rd7pemEedAaWxR46lgy5B71nJ0sGmbgyo/4E6M2WRa90bAI86dUmgIQLKnPaJt7zrd/Y
oyxDkX6fV0U7TtbLjjHYnJx59ClrTG7Yv6Nw0FP2u3m0Cgy6itNihLc2OFTMJV0ARFqBDc1Ktz8J
hu4dRrbN4Yox6k17HqkdEP27sr8LtcLZpRbDevNt/hhPBcHFYpU/j8+H6HK1atftyGhbgz49xbM3
nCDETDyGmb/abUv3uXeLZOsmo4Mt649gVL1qZp+arfYLD08YMTe2YI+JXxd8o1ngsm9TVx8q501t
citD+f7NPhRj6Fa2YsJ2+R9DL2Y9K48aGCfvQRuJLD//QlKLGI1aqcbDm5J8TEplCtRdn/by/gGH
6/fWhDXKrBzyEUtmqioUJbSspMtBTU+gb56KL4zgv3V4gqNufOpL5KMj3xg/LzTIxC+p0dFyn/3y
vs6DuC3UjDx9Gsvtd0jx2CdWP+krRdIBgVU9YkhYXdt6tp/y/Tj/+e8EWAQu5dnRVsk04dd6/3Js
sS6Dwbqs9ZOctRdr5qTJdILvZ/n+yK4gTtZPik7o3RMF/LzYrUhDpO+3AgIslVS/IbF/V39uMCpF
C4YqD6jUlLWHpyGtQIiT4nXYjVWJ3x7adzbBx5s+4FP6TaHzG/GvOlxcKvap98VDvnKI8N+76GaS
jwyHqUlVRkyrpFAxA+vXQFYqgqpmgKrMT4vXbyod48/j7wUZpdAhTBwpm/MeVsRDkpy9YC6J0rWe
wlbAMcvsk4hoAbOx6y4bsdhI2LWaGODHoCIUP9YcaAAf097PXWcidbKUAwr9oOb8mzyaa4VY3tBe
W3P/I1s1UlZR6SYcM4NACjiwwpHVubVxgpAYaHsgFuXLd2FObbpiZ1vp0KF14iX5kMxsk8eHizIE
z5QqMu01lwfGfMDCzFsdEV43TOaVPTNKjv6/D6MV/y/Kqv+vNKU1uLXP1kNhd/s8c36OlghiJtZV
1Vm1epX1fYJ5AMnI9edTIA9KQgaFG4bLb+JX+1H64vz0Nv5iO7m+cLtekliAA02s78odG4LQxrtq
uJCpDdcLWpM86pSdb6bJk99swamp3CExJmxDW2iHebjwFDFe+6Vdrvh1r8y3uHD7Q2Yc2sgmiPQ9
H1yr3rnFJ+uugcH+cvffsjJHGT4pVw26Hrb8v0MxhMj6OMBrYlDrAfIfxCIikqwuBekQUtXrB8Vn
PhFE3zKTx0Lp/raD/9TRCXBA2ERATOhgyiSiEFxQjlU7DzIPCsqF6VY638uH3ZHQAtd+IPX3co6J
Z0MgqMdINMLt39zk6/KjS/leaWjuB/+gavRefiwsKpV3tnUvaZxfZ8xs3qoXMRaX+zyG6R3KeGOG
aaMMz8BdnxyJgNx7QQ+bJEM4o+vScr3OIcXa2g0wET7F0XpyP08BaIYpjFFNTuwhaSJNlC8C6gl9
f2vNBHKHnlQyB4vlG8srfp9C5+gP20uHpp6FCc86LBGagCDUhXbwi/IZMXfY2R9mmPnfhaBVSUZI
3m00EeWfkXoZIOCkIKhLjrD5q3btytxG5c1/qQ7tVBtIbDYL9yspdrLOf6v5gYAze07ircgT0yQe
VwjVBDtccWp5sJ9cjkasnXoKIrOM8upmwdT4+cIBtZTFnld8VzA+sU3GRDx+BNfSufNrVDEWdqz5
r8dajBaqS2rPtOFDEJKzEPGx9es7umk7Af2d9OcL5Z5PdCBHklP7qViSepzMB5O8u5mgHnmxzi+W
EIUKDzi/Z1MPxviAGajj6Z/fBsOGn2z0uP05ssyrGnojYg9uROqaiQl2QF5Z/B4bRHyd4wOz/ODk
LgKAkVsaMWp10Tvuszv3xAjcygYRbutgohHcSsuP84WIpAd82U4iz1W7iGPShvajiBkNMIEiuyqi
tfOeaHGQ2JT/RLWYxj7Rxv8SDXa+fsV+QmOnkM6uOVnfbma/dN6K/524IjorClUbkQvWxT/g/mm2
zp7N5pEnW9f8E0SEafzkp5BaNq2cT91JAhU9u1SKyDbSUs0eMVfZPDlKqRE8zs2MPYmihQtDtS5g
Y498kH+0Vd9HAPrw1guC38BNo+NIpqocjqqfYdQIpSsMT1kByFBTZAV0h8I4mq5CLT0EIidlsMP7
ElL7g0nfvfDVYDQLlyR+JuG9G74WXXKE7FLODIVo57nSRvc+tD1XAar6Q1RPMsIo27YZgaGu33Nc
tD9cwGiFIMoQNWlVEfSkGNrIotjt5vYz11JNS2hCCFIsoy639EINpZevFf6Oo4sB6+kbJG+cl71g
hl82ryvLSIqtV8YmvS0uP7ujPDiVBAS6XMK5fdhW3XNMH0rsYQr0EvFTsh0o4ypk2gV2ehZ589fB
tr2/x851qxIfLEJm7tMUobsnXVxk1ArXmoNKTA5VqJNsTGBuebmIyKN9f4Wc3Oav74hW7gmAX7ls
flS8yrEdRmVKKVZkEUa6mxLrSoD5p/aNOZue2tA/J3uB+Afc0n65UnnzZ5FtCRXOz1hvvwL+/tjF
9wkiJN5wgCMiFkHbhkEAZ3DKg5t22ynPnObbpzxrmETyLyrGz3V28qggmaQ/k4mos4JlN+X1reiL
bLjy8Cm0jnF2I78dQibqdsjXRQ0HgqcpX3yoloqGNYtSn4u8icyPPZ8w9g8LcnwGNMX4SFdnx5W9
dsntrqi4GkW6i3zgejOEsZN6I5PvBFCVrHjQh7tr7p6BYwYXxpQqLldQ7SKxrMcorYEHVdYspC51
0G9B03ieIVc4J17kvjvYczw80NpiXftHzIvEgUFciDIhhWAniEx4+SuusYl3PxB9gaw7BNoCLGbd
FHCmKo/lEO79XkVcxHu4EVxpHqTBLkkx2c82kx3+coJ+o3o0aR3njaWf2nNis2lcM4hC3yA6ch7Y
xPoOedpbot1HRvZqUkqfvSxOg3/t/kCm1zrL0mhdgUp2DLmNyuqWf5Vp+GXe7iyWXeumNTji2a31
DsBTpajN7TEVFZ2B8YF9ZYBs7vB8Xa7w94oT+cam/hQAxKegOY5jVIFv5dodek8BBBlT+eGezMZq
SHcdHiTFBrLxiY/m0tu6H2EEezRljnxidYGmVtgupxLZKW4OubSQWjGLJyv3M0DrAI6x1d3zYAAx
R1nO7T0fXa3pmysEAPNdmMuplMSrkR8d9wDIBNuUIo6BVi6S7SLeReQsiPH2lT3CCKJq1JzRKZAe
rVIdoH1d6/bzn+MFmli6gSNvWInwR39oyoYQ/QT37T6tT85vQQz9PCeMQ0P8kcRxvrfCAEXaTmIv
r6KDZ7UKnyycNQUdt69ZdzyAc22M8M46+NNxmsATL9jd/0QrkoW1qqYM11+rbK5zgYtDM6/v8pnK
fpgGe90XTlLQaR+yfclbzwFsUP0d6OU94IjkOVwF5NanpQsj4/ZAdbRm80OoXSSpJKCDYb0o2a8t
IPyKWFBo2uzTxpfE0JIp/pEGIj1fR5bP8J5qcPqYdWpf6H917Xbwukfl/aXI6YmYs2NTkdBayh+0
/mPjeDLxjUQTqfHjsTT6PkBqZNZxys9SHdci1MIHxCNLN2aEGL9yezyYxV1r/kJTsW65gpzOTskm
TqfTRK7h9WFoR9gpo7TIdL+nzF5NC+GpOCfKUhD60tBRlhCryhbk6vaiKIq8n2IUyBgy+WHNaLHV
ofvtjG9kC+JFeb6FC6KRL+IYb53SUZ+ZWrCP4twVaT4d268xINtT71D10XaZ0QgS+5zzmfObgFy5
irNibS0KeM6RKERmFUf9twjrzazUiO80xAXV2NgEjcfVEL9gsxdhYixxpcjawHOVfchpq9k60uSf
U7y5Uu0Jxi4iBuOuIZFsvE3KAfcHWXgzqHcLCt6k905hIzQZ11IK/OfOXCUAJRBv
`protect end_protected
