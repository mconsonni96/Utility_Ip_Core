`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
U1HO8y/eAErPcw2a8/vazMAmb0C6BmqcAQwdECC1Argzr5FmZucJXduWooCR/56mCMq3ITPfXn/g
7/hCOxw++pzrI7bTiP1cFx+pJXvBiRzPu1c9Xz+0S04odYxGA36/dRRFq8GJWOKxmOfvBmyHECD4
CCd3wamhf1GOlMukCVXTtMbzbX9Ie0TFtLVrCqORSpJwOj0YTWDnMSThyFdy8Pbi2KRP4ZZSBKWn
gOuIRrpvacbpuTJLBbhhEpMi+xT3PMVAiqti93edzm0eIR/sm19viAXVLIopt4m0B8wmW/dCUHdz
nGH1fc4xPYPkOLIGhwbl4VzCRLYSKEuUKbVzUw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="qYBX3G+QhY1uXIki80YFCvvQG6cjY8vo+yluvCeZtEk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14640)
`protect data_block
hP79jbmEkgxKxo8/CIL9pJSAwdM2hY6Vj4P65ncxbAoSoJjn3HNfliyxDmqWOduifoBzNxKAnFH3
yKm2F3Rud71bUc/4ZCCiqyFoJ5gUYe0whWEsMsdQIlQW9k9vjIXji5WLzk0OYoEmLqC4Y66Q/NrL
IYQhbYylrTj8LZKaAAT0t9dSuknozAMkB5rqVXhoaLvUKKHQFUHMY4/xMPGAj2xbOQMHHxfNPHzv
iHzfEJlmMbsN4aiCDNJ6sH2svwbG4xmuHW9bAveEPl9ozpaIAFWhAzP/r9me6AZq84N9i9/vPQ+Y
1baCQasmcTvgchKjfMjnWhRBUE1+46yzR4jagUkjknp0W6BJKhGclGOJxi7uUzekAe5Yobh3ZRMU
LZDac/hnRSttVyOEoGLAZZHwYfHFsBbYoHX1QbHNJU9tDvjlJLZrhGGmflt8sU/tZU81bl11MPwo
RQxNCZ3as3jO/IzvRNaQWCCTsgELfUA++EAnaCbJQBJd5p6MbQ5ikuDEL1KWGLlRDVuimzirl1sz
i4DoMXOAuc5BZF6dzlC5BwcdsmPEKSSCVNFm55N3pLJcMMk5mH+yYEeRvh7yOK/zEOtNxvLHTwJq
zF3xdbaFXmV9ndK2yzFt3lxuAoH0W4cVACg01dUfPYYjeuBICX9Lt2qN4uzF931Uv0vlQcNCa0HJ
boeuQsfR6dvLIYcGnhgqLoUwArwocEvBI/lpwWnfI2rue2grmERr9G0E3z+9pgYTaJdLdYc34wwG
28HOEupJXMVsVeJx+UCqlTivLwlqQOC/YuwKuqJkGJ6jyYyLVUDYpLbD3PWGc2fAyRCiiw23EdvI
AqDYrGUCWRe70GJ21T06ohtVmn/oXxQwjPUTmT0+kmGtlg6TLjgPwxwivoArHjvGV4xBl7/ntouO
VuuZpWh0yXg2deP3cETRq0CcgSwF4aNvFVWh6rqwTWv3D8rC3H9NahfkO+hd7Tmq4Vi/tkt2NtBc
d6tqJFvl7DiY1Eky9KWUkLFtQ2IgAy3IlY9ylSuBl90hmhgZGoYkuv6NIPLpk4Bph5QIdlZbiXV+
SOa8uiiIeUXd2FiX4UcKguZWS5iJ2HeBvl0/lxUxJT8809JoE7dFCq9SAcCbfo/5aOcSNs4B1krt
aG/tDSQuRdi4qHwGNfGc7C43UAOFNTkcppNGP1iU7g2Wkqs7rtnClBpoY2PlscrOzpssvq8Klb72
t8n8duzLz13rpROcjsbC3ZfkUWwt1GYyZUO/CzS/qfaXmTY68Ooz4B4hlvd2Tne+7J2BB9AeW4//
iLamuQeQRf1DTBvbLeVMoqIogLJqjXQMNiqlIs/zJUzxJKqLqIwH4mjechdBq1faNEel8xPZVkbM
XrhczV0yrj4d3YV7dywZk7/CDT33RwBvcF2wFDeeWmKDZAQnm2hqOpx/RpVQ4bFcLhiMT4n2m4OV
3w3BybYlsQQvCQX1fRpZmzePAP3eDA1uOHQXA0F6B2kGjcsKXw7oAEieAYOEX4lWMYxUW8diWWeF
sn4s/3EHqi5JubNCGbsjCuzAWslfrKYv6Fg5StF84jN2s1KOja2dSP71ieRaOWblFEdXp7/DRtYQ
g/3sOQ7DbjBbhrrAm/ivnjSFuofjuHrp70kvJmE8n7RvePFUzbCBiyV3HkHk4neModET7/8uKOXj
Jd8g6bmdXTkieqP6RV+iAd3k0enCt+s8+Kjsc2uqc71jMxUyTOPGEv7hOC9KspF1LsJUls7gW7sC
5iSt8F+QZzlyi43/2+m40p/VmBnBrThcnolQuOBNI823YGnpvgqukr4uQ1Wk3WdHDcMHj7gkNTs8
lvtH0RTS+JedcRz+516gAXjUMzw7QmcK2F+7/mW1y6wdIQJhCKCMy8NJB8S8zS7Gdi5yix9PASxm
UhXiX0HnFGfri/IeDAvT4EULbBQ746+Xohb6O/1foB3wsWuTrTm2EVJYTBFBqEZKb6PUFpExyxpB
Z1TvVOflM6EWKrEYL4EJBZ47O8BKZyE2ztzSR7BLFxHaSCnWox7zvr+duj/bbkF7e3CfEKFv/FZ9
fiGxREJyg9exZW/loeQaP3flUwrwBZbPBf9H3FLqUSQMzbWRmpyWuqr55ldxwevl0V4jHLDyA5rZ
6o2obHA513dpupkWNvY3b6pKhxpSX65XPEAioYFLe+uiqXj/BM1tFFyY/KyT9voYl5k1KHgEXEwa
ha9XSFCT6i/NrK03brzVMfb1j+Y0urPRbagz1kgjS+4mOq4FPL7TFwKCIsEUlhULwq4f9N4JTTkg
/QcSkPXUuoW/QybGSAE2qNr8QGlpixclDy+HGM2LrHaVHq6gOswATe7+pmKq0R7K5aw4rNDsRpZA
p4JCYqBkjSK4HI+sG2D9n1UeYmfWCGleXG8vmvZq2FNFt0qIlzgLJpS3bQsDCK3hmfd8eKjtRLdE
TYu3gSqEvspwMWAf5KMafdhoBxyZeWCS0wVF126YxjIwhIBxG45VI8Wn18KK/707hYgmINtgnEZU
F8QBo7EI3OTywX+bcDP4HbZ+RWtVWWXZT1w4BPvEAr7Yzz7JoL2aSixHMxTag9CYZX/4ZqHq1eOR
ePdjBRVcI5VXdDRx3NcTWkPOeR6V+gmmkqEW5aIYok9tM2s53Ez7P4MeUDJ+otoIesIBUqkS6TdB
9QNwT4HLfcSj89tnbfcyI1mz4ogSEOlMOb6NjHvhiwZSH9ZbtqpB6khV6c6W89qJoKKVkdXSpWLR
v2HwgrvGzQ66FTeo/q5HTBb1JqjTei3SWzX2KE/GTxuqiJjSNTBzwnvjWfpFRIq75fkYvbSG5UFN
XMpkmUBrP3sQDxdV0vIZVyq+p0zJOE85d/YHjN2hjuqkb0oZvbbIXkUByYYuTd4Dmj0t7wibxadr
BkWA5IEpSnMSbomLo8PgC18ZgRIMlpXOWYS5jiWTYBAl5sBukj7FsCOSQLhWyiAhriXgh2hj2NDm
Ayc/223C3bPuSbQhVXEMdBduw3xMYg/EUFxWijksSvb3ufPenURRoOkJlvN6+oFuapt22kCVaEzH
6Htxz4kjAqM6IHHWuLECOYFX+QqQ+Ateq/F0fQCfp+lkaIH0q/Pesrk3/vtYa2dKgqCI0wVbxtjU
Iw53gRlKOqrbpvxnyH/KQPzreBiTtsMCxcFdrYdonK21J01NNnKLOAUxvluWUS5kxzzWsCI0gBA1
VROcCFsHaje3K4mbF9BJbffRrNVUNoyNyG5FS5V7l2cT2aJpdahD3LzUpGlFjVqx0hLRxBq8/Rl0
albFFPrw+z+/qIdTlcWrQkvMJ02Byv58AqWCXeSoMP5WCRJSqZFiueaMPSnvotcJwUk1zr0QpmUi
r4Is4kJ8Czr8s5TEDgykCtdy02qtZVGb54wZGYRetI9Xg2NXckN4Eo2cSVBtMhAyZN6UYmSr4mOl
IRyZVzE+wbZiq/MBD5lvKsoqi6RxkRK5aq4dQKBRt6/TkEMD8UtkxwX3Ir0DtTpe8WzfQ40ef8oK
tx5dAW5hg46co3O3Wlob0EMiOj849mZ+E3DnQ9I30NwmWb1xSgsV/FHRrufPZn2BBQ+7xtwvs+95
vWGRpGILw4SLeQpPcXu6LJ1efNXzbedMXY9rlQdr+Nvb+fWDy5Ji0Dk2jQ96eTV2DVnnbFSkh1bV
NFcJSBhePUX6NdM8t5TFyv3sbGz+V7/fNPL01wym45JD2p6GjLoB6gyRYa9q+pVq4i9CNEplDJKO
8IaSRV0y4/Gx32xFM0XSGwKNjHpbdUt2ckKAI2WRsYNMSc2pWAl+cIbHIcWe3v5qHrfsA7gWvn1X
hp4Ew3USHNp0Z24qpo6q4yf75kkcD9eov7oGTxA77jJEKiv9pe6gAIT8dtEXY3Es/Dz6sqNxdGup
FaM24rzWpZjcYQR5NQYJl9F+9xJ92/KKCNUBkD4Z/S37ARFEwLNg6bcS7k0d0p3IFZqiFR68W0rX
rwxKZo+Evvch7jjUr0Voo6Q6jwG3oPeLg6lhVhsBOdswfwjdXIx1MoLxQ7w6tOLR0kUfme5M9IPY
DnzpA5BFDa81BHYsluA2OEonf9WR64zFYJj2k1NQLCNldvwVsEzNMo3G+nvTgNvjDUHCKGRxexJZ
5wEdwgpHn8kqfrJbwoQYpNd7DzmG9GV4JoDqORvuXGYvSmzgy4oBk9S8DdpUA2VLJRx3aMO3hSDw
Q5y9JBLh8h+uEL0di8ZruZvT0VN6wHfZlbZ0lJ/DvvpZYV+pUGOhMXDi6DQk0shE6pxU4wxF6V/9
C/h6KKNYLIGfJH1nSxIAPErxj8mqAhzlGgEdviUtxl8voXaHfS13HEEBE3GstrokwlBp3JzbBAke
RVKTv3tkLVMAGd0Pv+CktEWpdVB8zf99E2MPXlnjUNKAp3p6YjsqUH1zIIY9sthSvW9T3Jw/87lk
gEUa5AikjVnVMRxtKzSHyXgWEO3VwBynak2ooz5jLijhnIQ5rWFEYYnGYkNUUnqOzYycI3mDzya1
OUggdrGYDFpxHQFH5oCKkXzvUB84GOxkoj+A4W4iCF4drbG+/3ZMLXCrsaJVIZPisyOGlx3ro1SO
Z8+Uy1GqQ54ocblND/+Qy09HKJdzYvKAwU5CdWLv1WXxPxeUhHxoRbjqVFWrB2c1+C9zuFXudYaB
jE4dfASN40cJYqnZ4gMX90gxLrcCyMSrTtXdj71YuQwsrzQ/I/TaESGjIQBGeXyEs2uF5fPcrceW
NoO2vHyuB5T/zf6A2cZ+qvhng0ym4CvMNgUbdLt2fdAsUEcX2MwkA8bZXBPSGLRRtpBEssWUaC1W
Ggy1yvzWaffhOQSxgfZG+68uMBf4r9w5u9RK102Vx/LMdweuoDYnfvTs9CCGL9sPMl7TixB0gKOA
LrCUgRG84yc5wwPxsrMPr3LSrSGNxgHUDxjXphW+aayNHx93MtSx7DuyUNy16wGnIVFcR7L5jjIl
dnQw42thoymxUCb8b04Q6Mxxfr3vxpwzv902APPG8R8R7nHNUcPejqwaN+2YufD6GfMmt34DeKrl
YJCpneWfdMpIsp0Jw5sp3DExf90oFCNQAessH99U5R/A6L/PPQ0EFWBHjGp0ET7Ar+7WoZaEcYV/
DE4uYSCGcRAtAJ3O3395zYsdswiXZtw1kOS7K2z/2Rz2DRKzlHDvJvReaO6m2vsDQrGaE09fzSSt
Y0gQp9IVsPUvZzynBH5EzD0r5EzBLNkk4pekB33myGbOSvSEnObsE4T6/x/YawSz5ZgMvbmHJd48
0qqKdjccYdNUHuQJ4shrnSir2XK2kzqv0x8HUTWlFmo4GGG56TZVJ81gmGLpu1EmvJL0aYp7BQSk
89/zcfkaetrBAUy4mXn+o7+i62YqN7VmpaOZhMrWDDMnGEYM9IPv+1tlVUmx4w1RTbidUv7KpTsZ
lFFI2wh48hBUP8VuJzzIYV40ka/3MLvHH5GWuo+wf6iKd5pE+Vo6mTnjB0FwFAqz2koiBJjdVyeQ
8+0Tkc7C7ZQ25QSCFEIOS0/98/AFjDHgEjvahzhNUKVV4CTEzRQI340+PEd9nc/vEQgFssLvEkBl
N2SNtbym/568R7q/oQRpBbJpOIfMrDhmFjnPDbb37OJH0qHRP6z747A/1J0hfzpiD3Gn1W9ndiMu
8UfK8lDbNFeNWEUq8J7Oh3w/AapoeWqtHTpsv9ZodYA0uqjyML/e9ZB6x69l9TcuyNIYOxwC3/61
J1q99P2+GSsPhmmoXDq2EkHaN1QBtVI3Kp21ZedR856gYTF07+EyyZcX4oHaTIdPAb488Tn4aHWe
bMWhlNGki6GDMQQ7XTiIGMR5x85aH//tP9UoMKcTd1DrJwDIfyPnPCY4cfLc/5xyfD78DVi2TlFk
KXzxbnfge27OAC0V8EjZ2KPdvVMVURQ79ZN7hImDFXAez+Szv3E8XkuaeymKt1rsQ8IYynkTJNRv
CgB+v2LYm9lA61X2elhFdU7yd6LlREhWIOCCmZAUGUX9R04Xx4z/NgrUOMzlsAvwEfGvFaftMRC+
F2Jg2j5EVtbhEW1ZJRVa3Pt0dB3KLpzcHd/6AzB9tMO4k7kwGKOPzSRwff9htKSypA4Tq6UJiGTO
PdYbpCgTtkEPwWES53u7hIGeAPaJ3zSIkWn+6tayUMjU+Yu/gsD5X2+g9ADHMTKbLw4A5iRtMpP9
hGvhu1ss/ZAEIpqmt9e88hhhG/NUd9MIoEnUo5Nxpj99laL5fMZlUlyiHcsmtb80oMwR1VVlQ/g3
IYxznUnLKMVd8zjG8Qu+yXB64qjn51Ot2fJkKPeHUwonczzSrAoYRIBffsrm5WQ9ovDIFKh41O8P
MkwJDB7PyF7pudNzkq/99slceVc3wppF6YXbeH83rM4WqMtsDsrdfbv5XwMYASvQ6pvui9hGUqz3
5HtzXNF+HT+kuI3UkYaHdiLDQcl8H+qe3cxUMuQMAs5wBLH3EskHmLa2qsYnP5KjMDKkpaI+aN1T
A9eAsSZFlmBf23EpJdK8lgho4CLjN6/86K8TGyKnFxz/q4sjfI9LyrvF/kE14wcr9Pu4+w3J+P4i
E/DW/NLGwl3vL+Pqq6YE/zI1AnkXBwXGZ1shGreOVVl4qySbhxZwx7v/y36zd6c96JXoEdXyGbsw
ta8ZBa6qgscosPqmiKugyhMQwi/1+i17TrUKMk8UlmmD34ArP8IvQpR80AzjF/EpGbXRjmugFJ92
zV+a5ncMraZFhAeSbzRKEZKqN9DZjQPN4vbtbIz0blzOqKRzjhwh937JtfhCFLlZqoITaxQlYQyG
OOrHvh2x/8gjM0Z/u+kc52HWS7dPYLMLD3hKa9iKRz6PngoaZe4TU1T/4PfRiyGetXZajzkd8tSP
h9bu3U5t/bDFE8xJLWjmLqjkWnhFHJbfgHV8QX0MdJ8HCPaVjjfVOzZDqk2x2N6y9dTGX5NP5Eaw
liKWbePJtZ+NAOuoVuF8Ka77gyE/jUcWxVR3GJ1xACQBe3CSDkY0Q6/iNdPezBKi+MvXp3CfgA8u
2pBXVKGBjVLkbFVKgPpQe3hWlUbBrZ4/Rr7vGdIgZxI8c2f76NOyUmySOP/MqjGrH4lY8v+n/Tmk
kvpUNu2ORSPwXeHhkuhfZFaUvYadjjhWI3HZ44mOZ5kglg1ohb25yiCIdNMP9olMODMA3FQvE/UK
kGXwVDxwXq3kPxeeoVIX6hyMsj6TTr3UcRtn9LdZvnP//cBdguS5RolNRRy+N8n+nQFr/8WUlDDA
A79Z8xpSouZI1WD1rG4UiDxthqA9xaRQfMbcxOr6pNGFN/1Fj5yjJ6ajNYVYTNJl5kOVVnBNJrXS
OcSPFywzSK5N+NMG5YlN9KPNowlYihPuKHcrawxYr17Vy0TQ+Q5zoUzbjowsjhUYiA9slvWe8oMl
tDOUdgyBRHqfNxGqsmZgbtooAHZQiEQVyyXRJ7rr1DdQtIDvFZuNfCoC8U8ENVYi8zJApv5hZhF6
QCenEQcyr9Tuauf3yZaFxFvHXBr9+YUzSk0QB0oSQd2YSrD3JaCxsUzqkDiXa920wU70fcM3vMmX
bfbKIPijK12NmMVSBZErGMS+8SY8kjaYYFiveLCxhkPdwkVXV5LEK/aqLHLNw7jTiP9dOtbnpodD
2y8SNJ575bWo2WPbIzPoVcGQ9TAs1oFuWFl//UL02iQ7XM2osBik7aXyta/Btsci5koZEVpAJRrz
TsFqeRKx+8u8GnP2M1dYjqnoIzyrKGR54rLaxl4RUeMePQ6OelHmBswN0eSqkU+KY2BwROl0CiLC
LlHwbq8ouYUIH3qVy4tinhG1jWG3QIXVvRGPr6QybTuGawpAf+K3Ri61FAnKBnVXPynO2spZsR0P
jD4IN3vuSn5rrU6lylZP4ibUBu9a207zNOqEoTIT3aHRi9WWMD5wCFOm1dMmAboqgKusoNnKObEI
SWlf3Kxyw5W/wUrYo28QEozkk3vGtcjCAK6WwrDumyYshGosEeYvtmWJRzN2/DzrMTki3UTtIHCN
DabC+xX24JIHFmArxu2Y/zhJgYJ4EDOVzy/7aha1bYurbZs84pGihQrSL75xgqaWEj21FHU3CMQS
v7PWmhuLkqnfvLjnk+EV/zmBqVAoukmwn/BIuMrIfhvc8GJZsc/VVaiDkaneDEKezzzzQgCgv4c7
7BkXL4rvqZLHQ1ufqoO0/an98hP5sqeYQ4s+S0Yj1GxlwLJOBilN6poWP0xWdXiSfYiJC354TMOq
HmZ2rlDsV6Ng9OF00I8nSHotH4K+XI5v/lDY0k7XZp/y4rRC8PIDkpNY3XKhCgZDSwLNrdWLfHjY
9mPJdzq26sksZJamwoFxNlDxD/qg+vExC3h4NLL40qC3a/Ck7O2dp6PwYbbI4hQu1aGzTyhXAMsY
/t0Su0IOeyDZi8ZACLegisAFlqFtwKJ9DvvQYw+Jagl7ne9X3+CovedfKzK5jW7OF4fOk1JmNc/4
1XYciTPosekrRboaDBzho82owq80+yhIyI2f6/XHu4I8vATw/jYztvyT6QHuSyGJlZFoLdIN2I60
F/ThGgNTuw+XsaAezJisAjWGm0JdeuObRhW+k/0zIdCeeFcPyjZhfL7cdGNZ+rEQ2LbguUalcVWm
/RTsn2tZHWLlkuS0mrTiqkUaqTbgGBI166hiSsKzfOOxm4OVUbgCo9d1GTS2wW0M5sHCxZbEKf5l
ByOu3kxxhBMi3gQJtdhnT+1o2j2OlcuoaRMRcUfqTkYA++3tuWsLrj54V736ZEdOZVKAn500yGR3
+BbWEwa+mLCFeMfv6TnoCCe+18qh2dWqP0NEr3jTlWnJu8yV1udh+kTOwr0ydm2F7HVikjy9GpSL
7gn+OucbE+5WVwSxSOSrwcNRLTDAoozo7uH/v/dCAGeycwkOTW1iQIX6FgGYf/1JvA8IoW7szyAs
VBwitg9c760BV+b7pwUNoKBMG3hLdKHf241sZlCtLyk8bsiw7A23dJIllcDVnK5NTJA/0zyvvsns
ndI7LJIdi6EgRABlZ8h4CPffAO9vOkH9MwdYl0fQE6JdknrSLJazZn4El0p+6pmDM2blEB/GT2Rb
v+ucN3wf6R3SDVEKWZ7gGADSq0pBaSMtqtQNwbdbEtV8PAY1Whqba40LtdZs+uNq74cNvNzMQ/nT
8pr/xPz5hVhhDnCx5sjnnxNlgBpJFJ2tvIYa/k0eF7j68S3LVryMoLK3jmK47TgxJge1drPRLR4Y
21DBbehz/3iV1cx5cYKtWxv5mUi5wSPqr07o20YKHYlfPZE2wfEK+LSQDHqarEXyLhp44sUjQlT2
upVw6JDaqBn/HEvoE1Ymf+idHD2Nr7DGUd1a0l/RMKgzuxHx0hHjoCfVSRebNllIAUzxopM1Z5br
G/GlCR0TRJBFBZYWBXU+SDvGPLk0vtMp+zTTNXC2qHTVJ7ImDcPjRQ+RJzwG1WS3VXdojVHW0mdP
HTk4+fK1UXtFQxryeWaCrwEFukXEqauWO7GHnS6MhCiytE1cG0AS9rNZ7sHxeeLw+4iQaM0zyRtf
g+ZII5xQfAJzIVig4KJBAy6Dxkgt6JaPlRYK+RYZU6k4ax5Gkl6PVw8WbtXqGh7lNn3t2iytvge0
xBDMzbWKWKpHD1cdvW2iDRibQn8ebyL8ln1sflfn0bp+yNflEgMealTTnNn2bpAE8UfLQY+MSSVI
IeDBPzPV8L/FhfdC8AGr/+S57NhIU6Pk8PQUohKGv6EWPcSeDJylUwp/l/nRixsvejfz9jwgxZXT
NpTx6TiCNdElFW4Mlu4GVLY0Y4KAMcspMUT5SmCROs0kTl+Y23Jw05eF5zOlVnmGyM8YBPUlFJJy
YwHtd+QV+Mtk27lq8IKCuq3eDWvVWHJjjo06k0X7idU9YK58Cc4T8gAVPZGN3f7K3WkJR40+gzIV
pV6VsGaefDvY1yQ57s1BTmgIvpUU5mfzIkDYtrANDhkwtsL7WU0rFEuxbm7gHleoAVbMvGvsJwtw
Zvg2nMJQkNsGLoSo+EgxDni2j+qXmMSk9YGn856RSUoHRD5LkusBiH6k3HAGo2mE+pVHJDDViaoF
2ipNu+2k9pM4VeKuGrecdogPq5d/psocGQXe/cDci5ZqTWX7U7Ud2JKNdRnFlNlN3OB8h+2ZP8x+
lTjr6OrS/TjS6qQOgWRHdN5eHIP+ND9Hhg67FNKmvrGnpwDqqnoIitUEtA0vUb81qJt5ew261zKn
Bc/nPxqFVe1AHoAJLqN/EZPk33Xm+49morIh8rV9cDnvdkEuZaGulFJoXl5eP5T1Y+l3NtZ7qWIc
7AFvd+q8y5YoRwZUkPfOhmhTLCdIY+VxkmMWQb5AF994eDo1DsU1EYkoLfzX7kiFMP08Cf5w1nUN
vqhqF6+c2qt/yQZQxrsyvCBZpNkCrlciIFVF0KaNu1mHQ7tWQ7El3d2dc3iembNF/AZKHBNbtMbC
IZd6YVy3yj+qtzSKF4n7AGbGsGOl6c6xZdyScI3k2ZqGtSiyWaHNYe3A9xUVSdvoFv2+w/qTpMvQ
Rg7pfgiCRyZPyLI9STORDjuQ5t9ATYJdblF3b3+oOXt3YP4e8mx7+yArpF2cSAZQkhGgSKLA0m0y
2t3rJzCFy88Way/aGP5fLlLHvXzvN3eSUKUYzBa92aS9300USK6FoVHl1w3xcDi7RbLr/ePokGOY
QmBTL0OWiBzutWfZmw5xXMb3WZ7wahhoDQNf6lLAeP+s7IkNTYdUJZnj8/Nwi5sF2a/fMhFGOU2l
WpYwUETetr3v7X4/xHrNbw+dnk4ljEpSvSkv/+RdXt+eiwXlk5Zzuat08JWTVngHPANEqaMhjA3A
Wj1tdYa8AXyOPI9BLwBqcqwI3RKAmaO87FaO3nr8tSNgb4vvup5Vg3ayQgB1MJuyib3hCA2LxpXr
2sZOq8XizX5CMClaT4RG2M3rI9CXg1eQ02kC1eM4tnV1zb0ijiWSv4lZeUe6sFpj8VL/HXER8OQd
BXp1mgxgE/i3X4kffmVmLFkFD9SeBVEMtaOurdkRotNRiVKGVLWLXiyc96P4DvBS9GlJ7bVfQaJZ
ZEHdNq0wfE+HjOFaUIfK/SxtfVdGFoZBUGtQUdVKTHprMijufAFYFzV6NMrv3AfCI34KzQKEhi9k
K3VQU7HZ3p7xgILhcqM2DIDrO3mzGQyupdQ0wDJjKyT0iGaYz1Yw3iUUSjwAbXFnmumfUTjyJyoX
TCF8Xxzob282IcR9KmUjHy3612QIZCew9pZXqgarbr/M0G29lvn5B8Ddp5Kc3SJz6azCkZGKh8Ml
SkwGnHr/Rj69PPxoWY4A+h83mZsIFQa9R52Fk/k29jsAf9TorbG0kfK2/1h2aoo++XZnXXAaM4TS
dC+Kw5wW0jtbA1IUGZSF9rRlGty/Jm6zhLGeFX8MRFN7/HBnQTGm3lNA6xGEto1oDmbhr2mdXFDT
5jvf84I7VdKiZqghcDzSXDngfgNfJly688VTbjjJfW8QgxheLkFbwooXvyLUr6MS2hDxsNxoIRuB
XjUi7AP6sh4xryW+VMKoPksri4zhsmohqGDN8h/V2P7ntH1r92/0LHkYT2cHDRb8Hcs2TQDMehsD
FF4q0QNEnCzeryAQ3vJhkyliEMMP1IrLmhB30a5hwPozNZY0bqXQP5ZsW9/5JJALGE/vWaoFtMd/
NhmLPKjJM/ZPgv0Ys0eI7ys9ainxvCq5jl9fnEYq9HRGq3tc4fFDAI/IKxiy3gDDb5QMw9nAajBH
1qy9DikXRLqY2EInScUKUpNyO4VH5zIUTWtGwHjnW1bpmpx0/099o0jsLvJRstyBkecznBgVqsS5
bdiXWojFhtt4NllY2SwcNCAoiXum+iNjXsTKWaDeraSvnDdSPtxV2+oxz0vkisXkdyO1fN7tj4rr
qMenKrymjjsbazJNrbxFft5EW0BhzRnv4gdHmY/NS2y/Vz3h0SQUc6BrO8dLbCquJonYPMgSvTHO
hOhar74SVPbqcs2lfccJPxlhTwgHq4S/itfQ8zLFrSCZs/wAVKkrbLt1lNRgWYW1AFvIMtr1on26
bh76H5HpHOAb3+p4NrS2Zfj5ks1fvgV9cv0SaGrkZERd35x7sCiK7hqqdLanbI1ust7ySed2fVtf
8uvEJl1QG5MP+1g8jDFEoFlyupJl99sMDs70ay849EqLv9m6sVU0Jtq4BElm8oPd+rn0dbhRdXKQ
0ajhzTEJlZUlLooSukccLIP3UDICGid/ImiPAyujP5UL2uTXrzaW08TUtDF+GgZUSB8MCl0FnaVo
XTaFge4LXxQ2RXM6EaZtg9o5FMuAxWafxWHLFHgH7rWbqe3w6x0SaMN5kAvjEHrVTyxy/12GvhGR
Laf5nC5GO46cL8dmTs+f9o9SfS6nkpFZQ3V4cAtA1BvVA1kFRHD+V1X9sqJ71O/droSgjr7VwJnu
mbiC1EzIuNfokgH0uCWHhMkTd/JZpz51j1auUVMM47JMZEy12y63acqmFRS4LGvU8mpYW+aBbCI1
FwiUvFHF8Zgg0RCGHFHGvYRsPBLaPbUlCTrPWhYLn1x6IQdMS99JwNsFClEuGHdM/Gz7c1eukhtz
z2da2vLUz5bHciWoxp4N7ypnLFVXcQL2jGZ7wCQcxHBG5PAEBL+MQ26Pti/UCzaYF7D5uOB3X0hJ
gsKTOFROtADCyYLMFLlP/A3KOvdFuGjTfN0EB9jkovLS1MPKBGZsbdvFzPDliwFatHl8FErwaiWg
ZiwCL5btljY8WYLd2quAltFofJDwq2ZBve/gvVhFn8o0vrVhzI1b8RSyc/JPv+s0H9FCJD5Opn2l
2X4Lqw8zq0zQGJ2uYsPf9sCylz3Z1M0qSPVo223hO1qsng+fkRm0DCCsxP1eQsa8HeZxG1i3yJnL
6o6asfpKE8IB4COWkQIYdSqtA+N5d+G1fUgipNkmF2dEqkCKHFl1Cn65vsjx0RrBxWwodEPGyE3j
ZiaVyGw4RtRP+TqSwslpBfv8KiUPdEquvrWjLum7dydYO1PxS6YaXTHiaoFg7j9+kw8Qg8Tzq3zX
m+JYaEMVNr38/hnmLlrs0w/ZX7Rfw3C7AlvczbCQYvG9vQkDxFhh1+Qy9TSvNLcSktju6xXPRLxt
YwHRypHRGjIpxyl1TTsZOCAb7xklsZSs6mHgcB6wPuthpPi31em7dprJ9VNAfy8hlMfL+kc70Yfo
pSTGmw7qp9bwWb1/nLbPRQTJcw69eKGPnZ4iD7snmdxSwxPIaYv08wg6FL+qzS/MlpclyooAMvUi
NbS06wFyzrDUWM5l+XK9O99qnh2aiRDspuZ7Rp7uVfC4OSWawD7PC2df7sgGmwvM1mK0fyi5YTpp
4d5mLsbSAPYZaRlWrOLTD/vxhO9nK6AbaDPfYFdLJlAjg75lVVOa68xlJoP0zl/p2NRyn3Hsaeap
ovCSxMYK4CaqzFXCbKo4mdAJ5wUgEFy6qGLs2uaD15qL3nbAwcpJWASrUMDpe3BGcJiNT1EyNWEl
ncdJS3TAMGLMNJbR4uVH6D10EbSxoXpv2DoVzDMT9pkMBzvI5PFw1poTDGDWMerHb1qKhK6Y04TE
vlMCq+hMvSEhbcUFJxqmhbLLDCAPSfV2AG4Yi2NcKMZcqM1YaLv1GXEcunZh5hleT5e8rkJr1KhZ
lQApFAK0kmNAaI52pg72bGSSStAJqNdEZt23DacoST+j2FdQAcb8p6aTZZaQvc8feYi5WbqtZWjW
BqVAYg1oN9sytF+1dQotWomychu6toJdXbZYBQK1qqvd1PzLrSA/jT9vUD4Ysp/JxdBilKTIBKwU
qT/q+Z4LE8AtZY5PcPISYMqkKjsScpnBNC/QTaLuZjhinN3bSFtgVfnWqVNMaxiB75LeV23UIuNc
LD7OLuGZTug0OAQWnOF0D6d5l9eHdvi4bOtAFGdMtP/lxp0K40+gWpVZd+sjVAvuWn4jr2jltadV
3bODhUzZav2hngbR1OMWlMGf4hJ4K1WZFNRRdTYzQqMY9CFuPHKAf4uEvFWmg7ViGRqtMT+Hdhjh
LaWAM5MoNgd4kSTdXMiZFqeVDgSWe4mo+iCeorx1R3leCR4OuS3gvzKf78/hMY3j0bO4utl86nKQ
Gyni806Q1B+xGnYvZ7pQuHX0tqBb6K0ieCBC+4QjdRrARTOUOYR0QYwLTCzdtQYObpkQKzabskZw
T3T9Joa/654EetKkwPcoqXbPRy4ukIyk26qNPe4zYU0sHyJeTJ8SGE+m3vjgFTL6KTCngXbv3FAF
XbB0GTNgmtcXSEIJu9mWKpKog0U9oHTOH9w0sDjiJj13IysejVUzJRjwJ1aIRtQJwLnZqaD03PYW
oiO23uQGDfy+FzRggOmdGOG/gO36pXHgkJ8v7E3aVFkIFwtG6EmFjivzZJHzoC4NR3eNUZ5B4L0r
HanXR1ZA0H8QFJ0vcWs1Aku9BAYN4VaYSmnelmYQWHEWbjlb5vTq+GeImCqGwj22baaBxLciHEHq
JwHF0TmjCactQYW/4dJT4jrSocPc6PFfsZ2NKjtMqSxD0ybFinSQl3mlxr0mwACrKuToGbWKlZRv
AgNxrnZEF2EUjBDxViwSQEHp+Rfqj+94F+jMhCzBObxhCJPH0T/Gm4AtLJgcmfv0WM/rE8OV8HwT
a+q/6gUjMpVvyj6tsaBJLCfDBQwomlSUBZE7udVGqenS4frjTByv0EwHKT6vihQAZvSv42vJup0d
dWAZIg3iRrm+rS0c8uN6sW8YYeZy00TFOX4MM/DxIF1w7vT8gIipZ9S3WzVxThUo+9L9/XDUsG8w
AfGRCUbASaxp0Vwm6yRIa/Iw2ZOWmyKxE3nZTaO8CBRA7tyZl/lWlIkv7SyC3I/oNOrEo/YVSGoR
LpQOxYME4hQifkWMmxjDufHWA8Oo1/ZNVjoLJjK3vHIxGH/goS1DlXZn4b8zTX8lrW3tzcd9igXi
ReS8myxyW4NmRttpAYQAJI0jyTIrqaIApCxolUxIMcb998FDXZqmAm/L+uonn+mEI5lU/XD6KClh
qfB+uS7gu4ByRpF3vD/HAs7Y5Hn+AMX9uu0tWCxUx0aaydUYDTox5RsbNa205m4LnxBpUH4JNflQ
A3wT+LJV17lSjxhEt/Y/m/74of2OY4RoED4hffKrby8rxmeKls9U6ICgv7kkiVhjJi2Uov1ADuVe
gquHWo4HtaDkWScbGchbW5PPunMcC+i22PUFF53JVHmPH7mrSrxUjYookHaLiqpoBKV50DA3S+6m
LH9ZwB+3VOMcIV3hq8d+n115q2JFwNDT0mHy+9AHpNBBHdStPFqv/kr22SQNLVODFZ5S25F47G2M
tpWcCSJC04CUCLxQwN4a7xEut8Z+V9JlUUf0oMeO8w2opFfwssR1bS+vFvPZq9y9WZpMHQssCIFx
UgS83T1aKzjusqK2C237tKTHfz7v5shj2MplM/Yn1KfObKyi/0L20V7AWYoe9o6wgQ8LaDlyZEPV
ob6M3ILQoKsrh86YpiuPG17L0Q+NGNwFYv4A7CkBJLstSwzvNrge/KG9F3swoNj6oyTatWCqxKiK
UpkF/fmsnl9bXxrsS95Xomd06fRZXny3i+zRsD6UUvqWsOiXrs3A3/vewnGcvZ4bRNQ5ZPCrLWi/
UGGwflXnUy9Zgl6FZvhXrM0upiEHM9w6+SyCmLs5HoQu804ukrmGysWDIDxAF8dhNr1jCKITlcig
41ZSQL57JTsQcgR9IMwMTddVLyvf4PxyhInNXu3UWiw2DqJ1ZFIZj2vQ4ogH5ZZkwzPZ275fmXW1
ThB2SrX8FQr4Y2y4eeB0u+zrmTlIYDcJlaW7AyahN4XTshVM3qtDVlKK0tVgyo55WGsCALV6S6rk
jwaEzfqKs2VdadoKEgzXmYTWPnBa1nGngz+rr7duZfJAixFEkSDq7pJh9kQvZ4609m3zMBx1iOzH
r0v8FDaKiaWQLODiX645//4k4FsQlhY+RAQ4jK65qOTk0B1yGoVdJNgCuosWJPYSd2aLjYSt8Y9w
aOyy/O0qyDFDpslkXv3MZpoz21RUJmkviA9eYebqtDVwc56vX9LRdLPnPVyftl17x9mkaGFcLZVI
W5U7NreLNrbEdbnQ/CVaFhffNdVJfA7dP+U0MTZh9zCl8VPTt/oZ+EwvRatqLjqaIEWCOVDYsJhQ
MiWXlGDeR+oFyV0sNcaDl+3Dg+bMayEu2pHYWnUV9v7bELOZZvqJbciW76JNxQIAbZWtgX2yDXzR
oyHs3/ydbzrnSXHsfLkhmIJLIg6itpUxTFt9dkEbsPaAyhOX7XXBPqXI3jJiifv+Yk3yJK08iaDh
fjN7qbPQE6/3Si1o626/EwrXnozymdad+uKPeRJh38nFzTp4Jev+PGTGypD5NJycAlkJFh6ZboCR
tzRd6CmQiZ8YGatiG411MfdBwrPbp61kBKrSqAK4JW/W1IYTcqZV/VvlDRcfQGnZuLQ514sSvI3T
y7eEZOikr3czl2ESjpv+OwMcKQDFeP0gqJJKzS4c4P2Q/J0Koyoy+ue41ZqYgVETRieM7GQ4M+7e
2w5T72/8lG8du90YtLhc/BJFSiDY9WfAEGPK4xNN/BS2DFHVGgCi+3fdP4TJC01n8QfkHR8Ys1HO
Ial0vMcMLmt/cFW8k/TWTIslU2plv7uw1mgeN+3yYa3LEedpUQHj88OTm2eFdiP09NALQQlF5YVa
fq/0yTg4s3vYc8IiL9Y8Wa8s9dN5OKqbJX4RdbRR0CsVDWuJ3z3w81jNmGM4/B6z/4EXJLgd3UBq
U/md2vR1vZlDDEtm0fAHd7LRu4/hFONz/koNFhb3YfTSB470ouJwLRfxZ+Tf0MoSSLx5fSBIGLpY
VM23DWe57PDzeMIgoR3chsOlqvtaAJ3FzmdLPgXk0pHQ/o6XRzScSZD+dB7XodzewRut52+O/R33
DQDiIJV5MFVvnz7IiqLjlB4NKN5Pyh6DBYGcrq8kzXAbYFlh27EXjPl1r/xD+U0eg4xm4ZbFst19
VM1onL6w+ZZnzFMSNwAvSzTIWMRiLZ3crT8qFObbz7agJ5pJH/XVpNpxsXdUtWDD8LFwy7GmFZYu
6hbSnzswesPBRUTksg4b5cA89kMrv1hu10TMsFVVDoykJiHK6rU/Wr/ksmUmvvOf9pJBUZ4Crtms
aueKNav/trkikAAiSUDSenBkN7jP0i7GFe3RI4yQWJWLCWXR2vWemB8xzBnxQygcz1BJur3Rd5WM
pWjuTCnugVqPrSBQHH+1rGBbvo8gRgAcLIkyBU8o1n/rAnpZWCdrp9YL6VZg/3Hxe476O6unwtHo
xDyvLR96Ev+Kq7SzeYOGGNv7vU9CvEQc5y/cihluHEiF2CWO1D14XFP+k8uhON7sVK5cI0L45DRr
G6DgTjWEd1blEFjHin+c+ka9CtAVPl41jAvgmBytno6poTzXeNDclxCaSkJyt9+Q42cF8QaIUJ8A
xfLfhXR5dMrtB398GiqwwiM244M5ucCZ33LG7hruzAFe+JMcrFYUI6hUQUV/FOgg6Eipn3G19K59
QBkj3i88lVm4m32ONZeTsa5dxyJYPOnwqbxJmrbLcOFV/T0k6qy1N9wE9lxzz5sjXWSdtR0ioWDm
SxnjQEZ5TYPfO3abzW1BS3tHKb4haiBD/f9UfPKOUSdyxNGGDFywTNdQh3x5VbDD/LzXru0WfK8z
AZQvlfCJX+pc04KfeXNjmDeGrLwQWz//Ujn9JB8/R2/dUmq0jaYDsJuj46LAMzJJTXYuCHk6hDGx
oNk/Jvd4UKgVLUlSX5CeUjlVAJpvPcO+XIlXnkJOuWfSvdNTPnEZmS5ezzDzQj0aHf/cU1MfXTb7
Q8vWSBbg6l4wS5/lXdqfPAX2jAvm3de80lCsr9YpKnWajsNwQYvQ0Rj49p1kNdqJIKyE0RsK2Ppp
Yk2SQdEhxRQXFqLRhcRuDizhMPZB4PLgNldkX+2aRGHShqUZyp+7qSY5nLeb7lgcUJVYkpg1GdCw
56jZv8b6GyTWYbt9X4ueiyKlCziu3zptUsGsuWzqalxKbfkpvOizLHHhiihDwAKYRHhjF9tnsnxw
LsBVshgiAdudifSV9+XmCijs5zHUKJKmqOgnOahZNJ//L5y5l7WPOfuHdQ08Z0RU9pFlFiIPcfkl
Pzl7CjipMwVdvm8bfe7nw9y2FgoDxjYKWDn7pLzHCPpIzPVg/fATNmdgmirq2YAoC0wR/YXNe+mo
8IT+AxGyT7BAnofwnlwAL+dxTWMcsWw7R6K3k8UGy4CrdRbek1iIhRBscFSt7VYh3TDGmaQ8URVs
PsrQHmQ9EEci7/Wov9npGF9FH4c1luAEWInBYVvlSxt261ENzBUaI3OZ77qdmWDKVVj3cuVsH9VA
IAnDrsWOsllqGoTIxz/sJLGpgIJ4XDCcML7WVXjhHAR82Gw5eOO6zEZoHbALi7qkP/9b6uuAoypj
ZD4EnfAr3vYIqsI7nBWFFaLRkZ0TSyXRU/qjJTLGDcsbKijdhgr7E/dcrRp6jwoJSqnmKlmA0cSk
onYG+8cwRF6ZySqdSW3kcuvwPYqWVS+gh3ZhGJKe2te51WiHWqhO2JHePw1KuJLELfn/CAoEgaZZ
qNXAGf9WQ0e2dWz/EWvU+LzacWA1yjm6kGv0XZghMCB+lSennozY91IA1fHNqS4GvGp+q5rrEKp/
dG5QFFnuBeyzLJOV+le6O2hM3z2me0MYa9VMdOI+HVGHOJ4MGME+ESf6w+HHyinClNJKiXkmiOve
JJSG6dkjRNzkrz+Ub+D57NObZwaXcGz2UTwIFKIHWA3WAlvOtHg4KsZiCDsTRbodAzbDnoz610/m
vZ/PF7FGCMY8nDS4DrznQ//SyEqOQ9u7DI/VJ6GSOHfX7S4Nk8Qtw0rTsmZ/ubfIIxYAerdu4qPO
KtWfzXDj2v4W42QyeF8H1XRTYaNCiX1S0aVvp1aGPdmLDJUu2XhtGS/P+PjPnrg4i/YWJuSTgEgX
8/iZ9RVkKmi9q5RI8ZKv9FswmZZAhoIWADS/oy9zLcNoJaFgPzq2TzG5yJisnirLVHX4Fl71mQ3P
UzajU4lPM5D4Zbsm2g5rZHDy+tBFkt38xOHdXnju1lQjt9U8xePSaIu/RruA2MuOFPuDijGdAu8t
BklunC7UQWNMmHlfGt23DpD+s8zAx4q1Gt9iRLa1e28MUdpLAZD3MNrNQZpTXVu1FqTmypytQG41
zRWrwIGC9Tq4g4yW1KE8lLZxYG9Q8moLLd86UrsX8tos8WpG3BBHyVr3MXHBKZXMpV4fZjal/NxD
7Fs1PmkLVkUOZ30ipCgB4jpoZKw6z9ImDteB90eGAnI9IJd6AkDg3XT+XOVAeh1RC506/QXt/3EX
jP9sBr3Yats+nSbO7x9d+vLeb/c/iJbh2fHxYHTJ/L98Jny/SNwfH1hNHzXMDlFC4DZIitM3lx4F
NHM1vHeKTObAF0+Dl0WaresdEqGZVzpDeUqsE4fBZHOisKc1ad7zd+QcBFy1edPCE6EYoxgF9Lde
3PMUtEHFx+NGsqdgXaH+qkLQjOYcWQLu6X0bpKGiTFLW5p28DzVK0pRmSlgPYk8z
`protect end_protected
