`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
C0wQikoZEcTSWwtm/eBxwTXxuCLMvQ7+RZorZ2lg1plnpHks/mUPKClLdXKZtroY3/Sd/CN53JTI
WHDLr519ATyzudRQ3hB2aY+OQf2T2xwb7kODoH2vcUPbuxYu9xsgJjfOHKH6qluQu5RrGWuA/hyZ
I3OsFP+tVtZgSJ4BrDeCxK+AGZ5DpBMDmbzf1RUgnLvzuF2xumYRZPcXM/OchWzEt1XuJycjDF4j
UFnSyw8wPhsGj35gwu93Hc23pD029mO6CS77z+f5RLJC7huZJt/BYkiDWqm6II4yxe42ySIZ+0CL
7lJKRaVKnnV34R8Twt69YymLyLnDDvy8qXY4Kw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="P49CiquQ+Gye4xCTNd1kSaLzvtnjx2mkcswcUnl1mbw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10736)
`protect data_block
yYV+u2lXX1gMhairtewwtkU4NSmoeb6n9XQbvfyvrKGi93txxo+R2FPLq5bTv9s7023YRfDsHLDI
6cr4lbEO0q4Dum1LjHurFYHGt4ZafkBsjKsK3XfMVLr0HLq9STWA24Pdx7UvkOJrcFoltf1bKsUj
MLwXatpU6MBfcgjeKYcC+ydDp+etBIlLfNk98bgAhaJG+zQrZmRTII2ZGNG7pRhxqx6ylTEJmiUt
QpyIlYPGISt6mFnRGJSSh0RCujn3+x746LPiJqgC3XqLaKZSqpLWym4NPVFIl/sVWlIojhtzvJ8M
Kw1y+Bjkrt+5QCpi9A7fuu35X9D1tIRAdSR1F6BIntptT50sigAlBQUrMKXBOoXKCvZ1lSgQs09s
MGi0gfWXqg4B9C91dDY94UnPffHWBCGnmH4gWwbTuho8RGqYVvzpHG3+OsiUU0lWpgjuZfieO8aN
G3MgB1XO6zE1O6uQGTOgCxB4di1lTEUFd9uYrOLR5MHgkwYuQNt2czlGCX89ipETSOlbefeR7vrq
MlbPGTZkYQFIkhboVqpXG0SyyjQJ6HL5zBJCim4loPw0QnvRxsmM6X9ZNLAtmc3SQ9vGDyaFW9tY
qPRYFIej/bxBQwkBWktK01h3BacPH7DO4lV392tVyKTKis456HA5noSNC+v+S44IKZuKkHChOl+T
Osn9Q2w+s79fOuGZYsXY7S7115ujg+erSEJXAXGV+t0yFhZHPpZqfHtUpntdo3tPzybyRwVtkq/N
5w1XRC1Xv/HIOnGK2Gzw3xEMmMmdcOpJ2STwRzC1bZja/atkT9h4JBwB6SzXWQP4pViBt5yU430O
eDx5ymfIAj/VAUhE2wwVwn3WrW2pUd1v3HEEp5AdOxwB3bCwWYIpGFj2ILvOp6uv7Dat429dmqOA
wCVqi0IUPq7YhYl1hHVDghO4A472E65Q6ciGWj+/p6dy9kB/h9PoZ4cYnmyMF0mLIS0q2Tzv5MKT
cH8YZKwGHdHiZnCLpJgbVinlsV2/Soir3K7T8uEUoEbNJLFowzOcOKXxS64H4/ZfXtw83OIsyDiz
QBbtADwbB3aoja2eHRaicf306NxNat44oBw4I4RbUqmkA3PwFpd/SMV8SZ4qQTjp+P5cAzqEF3wp
HfhGUjCAvnHNGNPW6PV0BA+WPy33KzEOIWaWX/DSYhP9oA1BgUnkG+CCoLwvC4vv1AgjPrsKcV/6
YApuBL1GjBJKqpO4IAHB7I/S1RNL7K+lwjh+uH/x/d9IWt+/sVikMm3tS2Z894UWMx4n6+SBqrxk
kEMrFgK5vvxEvuedxT3JyNu7FePreNMf1isE4FYqKLms8w+/KEmzzaI8QORxvuLgT6CfWCCmFAja
Iw7zNjIalFYm9YGuAmox+714KCSydZBOzL2RbCkO9Bi58OL6DSWG7BuLKLmqblhbVNAFzbYLF2M1
U81dcyXJPuNsnDdv/nF4inzusJgL9tz36BzsRdMnkrM/7UFcGhV3OPAMQ6WO8IX4260sh4ZGByj4
jttQLL4Ze1hXU9UlLjNhlLi6UxYpZGA3juJ1e/NByD65QEVHoxLMg3c0is5K7v61XBV9qVhnh5zz
PS68YhK75Pc+9LbQ3jSXvKOOluQv+Qzcdeh2mi8O6QnTRct+MaDtaPvI6usF/XI7yABppIss57D4
Kzv56dVCb7psFDc0mWdtRUrKFtDmZCiMQRnCvQMoiDYxY+Bg4loQ5HSX3sZJyDK8xyyBssX41ATV
WXG5p5Mz5LN0vGg1Fjtfdcy7lpn03EmjqkoIbag5djwvXgVUWrWeyvsV5dVz2/CqGPcHzGKMZ2sb
Ofx3VOGsdjvUUiJ/kK9w2GmU+izAlNtdL1RpzvLplGle+8fp+9gv+oRiXv6FKkpP3WkUJOxazxdw
B4LcKYDHyD/OcDyeiwCItki6o7KHe5KtzYXK0wqTs2ICJql+Y0nOzkxg1Sw/J9w3b/oC3coHqajG
UoDC1AqZaItf9pmjzKj3sFnLqsqAChN9OiOSBEWNoHxz6ME3otLdpr0SLio77cTt25dK42jxMV40
KvIXfG01lGiE8xvhUjwWUtXDfQJ/wDkOcb7Qj2vHlpee7nMQsqMkI2E88P6CnRggzGgFmwCV5AbJ
hXYpwTbgoxEfRV0D2Fghkzgd3UgvEy977snd2ufUoKzDD6BNyCCpNm2B6cxWeph3qI3cMgoUiuNi
V2x06uWgctX+BLAv9lcJuFyvBzEKPCvV1k4pgD6T5mlg2e9xlrYbg5lw1XFVkhKhU3TYZ5O4ZlMD
4R0msejGRDbgOjeZ3ID7BOOpsSJBUBnEwhaC47zT72hzJwA2MTBD8KIXlW6Dh0mo24ynsOfj+JXP
eC3lR3DBdW0qWRR8rRF6CyskAdIDng4GZ0zQHM1bxvSXAUwY4rXTGfRosdMWqc1hZpE9pCQeSqWC
6+p37sIePOKPFTnLLb67LzraurVwXAVccOqpDyHtrgjgQDqsdDS3ZcUzQwniJEjQRJ6aE384FfmV
dYd2H9B+k5/u8RwdGLYSuY2mdbUNXeRoZLCwyBgIuqZfpN/+0EnUmpt2t41DFpqnHCflb/ea2q12
DXqbZftJ0YvZKtcq2/jRMA6d015aysZpsta2HV9r+z1cHEOnCJ5AXtxiKCENQGu8XFAeZILOCWrn
izZU20zCep0xKfLk2hVq1bqfZzizGgp8TWXaeWatDhIMyzNKsclNt9GLMxqIXm8umAUN9RRk3ttn
CgNtamOTDp+7ljVjHdiyFF6OlToMw/lCcuKeBc0m2TJURgJCWb3be463pTvDfAUlPMupM9FACS0e
bi76+CsXru9YkHDRwrR2+KawNgLd7Lgqh6g7MEYzFaGWpg1TJ68ExgQTEBjgAWeIigjVnN3nkoeN
jeuz32EVKoNk/r+IntoRnMLD6VygOKcRaVpxwhRhUeC1skhXZR7/55e16Jz91lyV7TxvfvDmsIBX
fpi+uXTxbTayyOWezU75S8H8VfUZK66RzxPnppGaTfXYo/h1xSn39cHGDonKFAqQiqbXX+3VwI+O
PwAfluUPWgrhkLf4xsZckFZg2dJLQYGYyS9vQhGxgOl7uUkdmvAnWsMnbU329RNcjWsBG+qI+KTJ
PBCIX+rkrVH2ephOmrLaT/cr5QGvQRvLnMZB8dDq5KFxkOsnPRvzX6c+sBO6nbb0QkRngsPywHW/
n0LVmoYy5N/x4vbET4N25qiXRDbV/SItiob5sOeMxNyzygfDxvZmGQPskSqPi6YlthMzf667RSIh
8h/9etZezoRbQu8EDwOrv9b65z+O9UsFbzqqRORaozwSJCzlvrLVZG0gb+WD70VJN8bFTLXDRY/t
8d4d097IBQCws2QFcp1+5vw78DobnOv8ikqRhbk+zDMwiTGzO67Oen/Qmqnu3R0nNo5jFFR06eFK
xQzd8OS5Lo9fj7pIipFrz/sKFMXbqEmOjhfG+FG6Qr4INJAZXLduBcA5kqv9NlT8JvKqF8ZbmrO9
iWmxrpYjdoaiXgCoXTPYSTplV6p8RvdJhi6ZaSJRfZAMCaWYthXqANTQJo7y8cg+OwIpWclGDm0Z
qeaDOKqHHtMPuJIQfrIBiJooQrHmWLjfQOFIcWE2uVY/E7MIv/VIXay5O/RV86a8iS2u28rxZROx
lcGT+L522iGponH8toBmrBOFeTO0LYY2n+ood06uHRycyFp4lJsf14o8fs84JoHgTKiuI9ZaLcgi
MYT9Ujt16tuudUiLcQHbIun9aHlxH+7HaNedvPGXq4s/xapRartOC7C/uqx8+dE8Jap1oO9AwZu8
N+Tq19epN8RtsgGBVgRcwg795ymBfnWh2kvDQH77rHiS0YjUFBV3fk2DnrajqSP/eScJo0ElQGai
bKYZBEUuZTA5FlfmC1vCfIbyLqlpVB+Z0r4aeQ37mMbCUbgCOK0GTHRih+JU3X3FF5J3jos0vVtT
UTi6tSwwSTk9PRIuWf2BdBOu4L8Gm8dfXt4kWOX5AY9a/8V+2Fy64CN+5/7WBql54ga3mHRefzFd
fiF7rxnFHQEpmPQsdWbzALgYweI8oVa5IBlOoLBhue4dfl525ta4igIrkkgCPsB16Fl02AL7ay4T
aU33Mg42V+2NqTCc8pMGvR5rFyxuVIpl7BdaYUt6CE6VPlcSwfTKeZ9UOKNfIZMxKy3mSr1dIo98
cLQ+M3Lj8YD6z8OU46X7zGv02qPBvxfJ1IYTiz+kG+56zusHCEnSjyOk0caxS8OZHM2pV8p/JWOn
OY5ESulBvXP2TMOiVSSUNjCSmvnO6klwhwmoRltLxZt/RS6MyipCHLFflZOaLAQdEx+BvugQbIJD
6ZjV383K6Q6qw7CrdbxMcle7NYfZw+rdT/gHfWY1JoUILYxIEqJ3DzDPVHseIzqYh4Fk4fBpFTgr
2xXWCTa907tA35u0ZhH/ffi7MnmYuJvV2zHkMFGweAJ9w2FVn773/GBC5+OV6RCbGPKbwW8Zj5m6
zRKBc3xDK9MXghZvK3uVnE692sBIo7mcC7wnjWAc2t/MhKxfj7q+haGdzlBYTVdJyl4OCtUVtIoJ
766ap78ifZzhiYLOc/JIlV0mpbJ2dhqY9RhimEqmgGgP6rY0M8MR9WkA1+qQOw8L5OT0pEltRHkr
ljSsCcaQnwyDZIyG6emaZ0rZY7oBHoh39rARgzr36eH/LBoPAu2GUCM6vd91a+AFKl/r4UXkXoNu
oW02T6mqnwBgJfamFMkEvd0R4XxZceF0CTNt75O8vbX1NMMCqnizqWyCxbQs6kTQkuSvx4kJQID6
1T5NUAEL5lL05zrIlFpY8NvoQAl/dOw7So6ql2YYC8yWwaX1PikaE2DWAKNK47bRPLsKlTLuaul1
dVUYUYx4sTdlsHXe1n2yJ2wokfdPIecoOJkVLwKSG8DN/0hyzQWp0oUt3YVxBtsJL/755RmoMsKG
zW+YaYiRonWMQEeTN5+OJRA6Izacic46kIMPJzDp2+xUx1z52CD9hwl+xjM6NHRWrw5VzpBRiI4/
Jrk0DANCSVdjNozDB0w4pLE58uDWkFKGkK9OUWL8mjgFZhBTw15nwhOeJtHvHM8ew/eMQhTRmhGK
u1WTj+PRk8WZqjRJ6Vum/N5y+DJosqrIgYYEy5JXTMABltNsss0T30Cydz1ojXA2Pz/t1F7NxCGo
ru2F8tjkaP02/50yag/SAFy6uKkQClobl2/TequuCtrUlNLMhgYTPORBtH+7Y34giynj4pNZpFJ3
6mA1h2O1I9M4YDlxgm0BXpVuI4Fe0pGOc+c/adClg1vImr3yWkobYFSKtFRtBUZohcuT7xpE9NF1
EuFHHGo3kEMsNK4s9p/58JkVKKO5+DnRsmlOxwBEDyz4Y68mdYlY8t8jEtlsPn4/1Vgn5IxriVd9
SonRfhE1ob6n0gnmvMyptMQQwQuO5mKFbCHOQz3OUZCf/+NHPMKv0Z/EwuJnM6TolVqmFh3C7oGF
8f4vKnk5tYXAK7BgGQArxXzv2LoZmj0L7YRQN0X9Xbq2sE0Cly815V4s8rqRnvBO4rTVLc1UOPXB
fZvVMv8dcnmnF4y2jSSANEesgsAbPvKF7Jw7sfqo+khBkD7fnvI6UDX3cfIcXX2wXpa4jraZLIQm
MgKmivJ8A13xsZoNfafDefG8pod+/MtW9TszdL+bvX41dEs3HFWgfSbRtR7w6SUAa4C3PGnnXX6W
x3q0XkxhHZ9ZImPsxpkp5di+oXbUoeT2qL2qrigRipCO2Od8dlJ5BAXf8miWDoVNniUZfyqq9YFS
T7Xv23i+PWojt6lMkSVdD4aNXqtrHJ9DFJ3VpPuOxmqZV5e00EQYOqxLUqEJ4bGV4SymTl/1h4aS
tC44AKX1x+tyH039orql6wbHLqaG1YCWM5HvxvaY0QBlaWDERz8YZqzw5Cr7yCxevK7AyFs7kJys
LZDVYUaCo3xQzSAMWXv19VVR+TUdrzk2o0TXg3LVu5yKQjGvmztuA03SV2GDJbDZOJJ1NaDOlYJh
EYSmtjaQ5a7sdDEMe+iqUWAWjMKVRx7Z/9XioOOKdBAsjv54R/3esr0uNH3prH8RSuTr5wjIdC8h
5xJS9DeXK39w12fxa76oNVtI7fDJGw+BG2HqDvBi8b0GYcLIJ8DPuxy8tFCFz/yjOZo9eoU9ovDV
PTutGqRJQV0jWwx54D3ohAMVqm/OWkqBr75d/XORkIKhmcEdFd7RQOeIqY2WX5fLzzjo1+eKj3E7
Wh8ttpQIF1N7f80gxaHLQeeIywpnjbLK0DAVL6seIK+Q2ziQbL2pxN1QI/fyHpU72FdyBBUdIb9U
brxgb+i41btV5ge+Jgk9iLWNYFsgY15AGxvWz99k20orlkEePDJxuH2B3lePmg+X0J+6TMJbZrPt
0hig9x5iQcZwckTq8RSz9GHajnVpdNhYik6pLtvw98z+YO72Na2O3UFNLHcOuKOFZGdz/60eyqYu
wKKSx2DX1d+6IvgGIrknwz54qZZv7nLt0T1oE8XqqgngZUBpAHytoxiMmcgPgXz2Mf9KcgtoXEBb
Rs/kiqOtyTl96LoXI0mkLma+lSe7U4W/z97gYQ+vPc7lJVTnoLKRLMAGy8vhpDfFlxhMqzBYrGrd
IOm0PL5+HkDrRH15In2Q0DxpTLcfbblx/J4As8QrVLtLpMbyG24xpAN2bnxdIClKIMD547Fo5Sdx
w6r36oyZatG4gyyYoc1CglcLONiGFnYSUsB8d6LWF4PmQhDdGq+Wb4xXDC8uu4RN0NvXjuNOtrsc
qBpu+go6HaEzOwzIPLGSbtpPODUnI2SQuINyTrqCZXco3es3/WllaSQ9tgAzE5DhzuthETfAPlWm
7Z1tgI3iLYagiLrp52Prc2n8ftDEUek3ab86rmsbofCrsK6FjQFVmUVquNl7Ypz+i+Qvd024B8uY
ApFkX5pgrzXpCKd/iurHr9y/SeOQPzBPuzR3saTgkCdi+aOhBdxygC2rDG5eZrO1af4KrWQsgdro
jBwT3F6CSgfJ+trY8tfCNlFfAxHZd1o2kptiCEXU1nH1Gn9x0eq9bX995peGmeYb926Kc9f9/HYq
EU/VqnEL/JA/oLUTV4TuWkKYLak4xszu3reed1P6DnBIEfDU7O2TCFT6WBvcJpteLTH4PkBOAULz
Us0UM4LT9Fep3lRe574aLqDY5pKoyxyl+dmmblCKE8XkVZeHZYWrjQ2YN+FSix9p6y3oxMNOu/Ob
6rP2QbDTWPr9/C24RzECw9VOrBA7PykozQp+0VstN2Uy+cXUeNPNu/73cGF2oqYgEnGsS9Su9chk
WaE3Fc4wlOmagGlB+OQEaGtLiqzM2xpLqnmsekvpnpDfJTBe4+kQ0dBGUovypbfteyDQzd66TvcK
z+IK+nlE6TprPo2kntOpAjEQWl+YpW24UVlyG4ARnvDBWceNV1W3qJrfPMm4QMGhE3Ts7a0CpgA3
g+6n2kCKIPocSyTeHZ/5SdwmfOlMrEoZ4CLjvak6zuRNnlIfTzyyamVh1OZE8dKwddiIOvBjP8hw
hHlQBzK+FXNY55Zzi7NjOQcM4LO5/Cd5Gs7Kvaj5KKlJjnuoPKX89BFXE+YrUwrj6OlNtmz3pZqy
gvjWq++ks5u25Mw0qJ+VRJ5lguRSQTlnR/zgl/e8ObSByWAr1/v/Z31ZSByxNt/ZPhFQFGI8cZTp
9HnK4gR80b6nCofoFRqBl20uvCU1CIpQu5nhjFB7Y5DCiv/lw/i7wFy4dLQYvgd5tZxr9zXYpoeX
jHg9aCCpoY6tF2uBHR6nvESIJeNfCxuc8ytGEXkTMj9m0kySvb24XMvwf/VHJkvXz6j1ak5GB1bj
CmTWVulIwmZdh8EwVVEygoNDEWaHHfnehe4vATrOVEu5l6DtpT0cqy0RdalQsqxnnEt/G3aDiGiC
Gmn3qOJwELKfhLTy/MQBHu5uJIYxkE4mKlpPbaxmhcJquNTKdu7WFDjsxeCLySnB45jnyjK1PNPG
LnaZ4y7muIJRqaDnRRs4dNGqgXvNFSVI5FNO0iYzF/6zoQwPHRkuBTCDdlzk83ApFmPym7GxiW1K
/+ybVcGSMmPBM6CDpLASZfH2PWCZTjddd8NxI1CbVAQQW34XcC8stqtqKocUbzC79o2HVVQGgUQI
LR2Zb7BP/FiiWitNgYvsHkFxE2QnCyFN3UJFnt13rwa1GffnMwRvCeMc8VtW3Zy5WL0UgAaKFBnt
ExyDLwVK+OQbC7ZGms1Iqdi83Evbfr4I+sg6AAaebHJV952/gTAU/Afrg4mggfD/y99vRKLjH+8B
gtGCIDea490ygExdYzFyLvM+o5x9ccg9PPKGbR+cBARX9v0Nul5sq5OHsmGafviUEWET185yNmOb
YhKLyZ70XXhNfIafT/MtfZ2m4C/wKGdZsNrY5/G/Dwmx9Xv9lpeCJ26O3TsZP9DisUz4RJHa4MlG
/CrHzySolef8DfTIo87s11ruO9tl9rqsCi3Arpn+n7Y8VtyCj8FX7JTzUfmvxhIOHu2DoAVoMGOS
fVjORmB5X5LmcIsm5XPFfSKV3cs73wm1WjqEtfEe2mlvApCexxPQZRvYOBfuIp6q7eX4rhEFduQQ
P9el+G5SDaG2kDdsEcf2vTjL44BWRI3N4AeUDNWRJ5MYWnzopISnXvHl7K4tGffwfgT2ddWS+tbe
xv9b3QJWmOVZoDr59wZIdNyVBOX8425E2OAn9zbvcCbQyuDv59AaNhasPYxPx2ltKrbHf7gdcgop
fkZ0jOe/S8ArQg9HZVNHGknQPcHZmdBtBTIhUzM8rr9/ziuIvhPZ5w4KySowaBLzAJrT2Mp4q9wf
fYbwVX3QPwDBHQBc+cB6ZGa877ktTfoWR4E199sy54n+1F7silbdzDVdrZRkDQDcEnFUReCSzRr6
IxMUs8IZAUsBEX5otB0sAY01XLiGSBd7lTNqQvKIPjNwGU8fxS7hzugCcd3phf7OWwxbEUjtolxm
NVpJEykuZv5ZO2npktNWBY68kH74YAETCKQSDpiratitFLedlPtKTaaF18mN0iEi8QCwKfhLP5HI
bFclNmFAwsyAU+IZxlbLz8QcYnPuyBMQQDithbsWkYoroEsi9k83oayyqJVnAZ32AZXpah4JmXrG
z2/n2vnbYAc+BSzvv/AJlrvzoVbl8dUcKemC12xqvnOT8tFZx8N//954gHJ44yiPR6dzm/V0Jd8J
8XjmFYnzNhD3eWhxufNxU7UuPXD0vPGEw6Cwhyh2RVigC9ZQWmsOZ7+GZWzAg6SsEcHBpM5ZboGC
e5zVgXE4GCle2AT7VsdcSmG0hDO3JBkLjYcGUOYOfvdgy1WqFMKe8N3eBCo+pq/0Ws95QFy1iNQN
k03pkxWF280hNQ+5d3zv34vvBtzMWaYqRX2GsnRb4hUVwieJFn00N4uwqhdUWcPmUSxjJVLgJ7FP
DcekskwjsaUVusuNKmX0YC5O4sQyXZi4gTAJlWwwwSlZf8EzY4YBPmVxgZz9XEu80UTSv4P9jSxm
4uHwm4WZ67H71Cz6nT4OkpzDBA+gMEMaNtXCau3Wp1xhpEc8p72iIu3tEmgNhe0CAeg96gqW1j+t
OAGwWi5XY9I4EicejBqhjW3pZl280oUQ9ZmH1SwpMee5hHACPtUL7gtQe8zUyAGtXxa/dYq83OJu
sRdI+t21Pz+E8Yemst9Bq+Mjp+A2uA87kvskun1v9M72nK+b3GBzeW3R/2Cxc6ld8pYvzRj84w21
VDD8W/PkzWYOx5eBQCrfr8/tplTFwJ3CZxMRQQH63wzYvkwSnUPiZoPxkdxDIuV++m8BW9SASOh9
Nr/AU32L7yaKyVJHPYybws6EhuX0QJRSD9WnAwFEnSf8V8PDDxFtiP5pShhGzvfBSdgZdZTau8rN
AYSUNyJ9ZCf2dy9IKcfwLmqRwxt5r++bLgA/2j5zYA2ncUrwd/W7YMOCE2iRZ/tmaotoq0eQKGDk
XY3t3yvfJWBtUn4o4F/sp4Xail4mhcoHQOp4so4Zm0kZ9aVwF7L4dCrKBSgkuy/7DasmeH/TRya6
PHWW6vveAGDRzCUbkG0/zJr48ScRhwSuRhQ5z70XrLqSqf0uLWoaoYRVPDeB9sSFRTYvXlNsQRT1
eywdrLVgtaaTHZcuK+YHxMnkqpUebYYraDpStFNL2rCMuqnSUJFe9UM81cvWX13KvxgyS5+YPqXC
ChnAVfxTu8t0unZ1TyDqnadfKpq+kDl+uDjuV9z4eyRVKA+e33yNRHTWteszgxZgImGszCjv1qpZ
BdUjgxp+tAX3hEe1edN2zxjdtFKCqtWvCAYJCCSkxeynrOum3hY2AJTThlAhSeXZhytus8bk+XK9
KRRJ0mCmYlAhZFqabz4O5tA8UyPvrMG4ERPVqfYTzz5KUM9ObUUSBQQOOLxBQzLewtfXuQgZkhE4
2itief9HeIuWKPLYyiMXNA6sDKamcQhzM+xbTgCcmZmrSRFr7Nro0p20zoKV3H3mBm2eIHmVPnao
sYYNsRXT091eMxp7oxIK3rlgiU2Ha7bsDvgavOs6bDCpGoubpOSl+Lb5denit3ZLwxIAlJvXjUyO
JU13yp8NcQhF8/cyRsKitGeHKOZcVaYMDBPvEME5qAxwxT3u5RLIobewxBPsmKMTSwBpi0e/vBEd
l2sBiA7PJinEfG8Dr1ZckD83SW0nUwB+AHvWxxcS2pG2LksJ9/H+W3U7IdzW2YsFSwc29Da8k1ZZ
8U2oxGnw8RjGCYF8LvEW29mhqIDPzIyIP4Wxk7Y03EUpVWhpQY/pMPp2b92QcsdQS3Ge/I9KRMhx
TdxVunHWZTT7cwedZyFBcV9P/iujqdj9EbZ44ook7JQF132P+c1h32Vl6JZ0c5RIbkWL653G0IWt
f+QeO4q68L9to3lRE4M7T8lX0hECm2CDLoHDNx6laF91FK/ZTo6k9cb0palJfGGna32UtWPJuHyE
bUohcbcWk+734MX+ZSgjD9sEshJ87UBrwLvw/BeP1u+XvtTdvO0ewEJcFRhr0UgoOdRlcG3sbcqF
mMgurOmYx8GfGzqPh7Bb4BxTkaqd1d5AwER4hyipxS1Ud5hHmu16RKly8yPzhYecj5mNlVURvhwq
UONNef96ChlH+akfFWAXZU43+EZ0PgpIc8XR/GiPuNEvSIgzthbWQdcaHH8rpxnNC8GpFSD008Xi
uQG/9oXeFD6aMy7aeRnjJRI13ROWXlnCzwJCuV6gzLc7wPhBswm+JROtCE7JaE8zedh4z7LUEfAL
PUMT3Z2SikZTXmttF8monEkKg7xh2/nfN/IBFqs1mGSzpYjPa+IqZav2ZZHsG/fPzdfL7Na/yNpz
z1cb4snx2vCThJo4PJ2XZP+tUdzBJcruB4r2yghZDiKZfV9y/kbjabXTampTD5tp4ISG6+T+5HR9
H3l+YPm5T4Nay0trVouGTCFkGh4HfQpPfr8urd3t9kLh21ZiWkQ7JvwP58ny6JrupzE5cJT1BZs9
PcFdYL06W8mhWjKseq1MyR/2MRoWlTCR+DNsRUqJLno0k+KVXKLVIxcewQgtvT2ryk1NZ2jNZi/L
wlW6CXcN8233TN/V8Uv5r4P8jBsnULOWkvqSD2w4IkQVQtjJV7p2vB5+DXwaHqgS0OrAHmuDoAdJ
zCYNwlGtSGHPqKoQpOeBQG4UknofoXI9MZEf+gOGvYUEycQG3qkQJe/tiVQ3lsgcCY93Z0cFjJBO
C7aXbsF7ZquYVwm6R+3EwtKB5Sozq6113+KjVw3qduVjVjIzqiJiCHSOl2nw6nVJ0v8Mta+DPWKe
Km0PMRlmB1fQ2VKl6+wzVozSaZcO/DSpQuLMDqmR96jlvpveDXM2JAb2ArnyCXg/nI46axIVc5qN
+lsfV2azU0xjkH+7fluaNC0F5eDtLY+/SDLIsxeUhzkHGFcz//IxsYIMbJFtmEvfw/Maek7Sml/v
o1Drk4dEBYKRvpbHyoGS5NblucYTG9VbTBdvvYwGgTXMZGkr1D9SbWzBpoCco1Obhbv/B0p3sVR4
n0sWBrJkxkfN6tDVn/Mfkm9ZMeywGbHEDbZWECehEGJf4NjCkIn9GvdZnlsAcI6dvHWUOUXjJa5r
vOp68XvNSV7OgMPsjeN9KQto3LAmURXbQ1im0KqVHpebzmaj2Hr1nvYdRvr4AKDYMbuP0yeo69W1
VaEWxSqJAVKlQLyOb+VUNSqvgNNKPTE2GCw7Y6FwNFQ+O656FxIEt+Wg40fzb+G9q2cVaC8T0H0q
CqKMBRKp/jJTNuFAqFdQs7qdvGVzrsOvL0mXXJFWqiTm1rkE2EQzeWZbXKEl/fEebs0TYBA9O8T3
tlCNBvvLAJixjeio/kWsLLKhR3r3nLRGj49zpxw29eOcKNjfC+hrnyToyyto3jAeB+lW6PE4IBlK
nP/4XlGqVWV7JUQ/3J5CaaAOrSbDVaCbX8OKYXStSLz81UGGmF8x7FbVKvZNXCuJUso7GHfvb+bU
L2/AIIPFybL2D7+SUBtuXPkueHWTLGFwgK7IpF5ml94/nmcNwlUtUK6oK1Cfb2S9v3DvZyFctCp0
o/qwHwT45fbSKxfhAF00oXbUCUs/nZlcYg6UgMa6hq5UNgZWXYk7t7Q3/8vUG/LpRXv1aoD6yeMF
IudUwnG39uupBqIAVLMLlw98cNRCxhYOARbZi5/fkU0x0JiDpIBIJBCvmNlhmvSKyhecKdpsFQtd
anaCPanEB4nS5pCS3Dzb4onFeYPZPNmFNEnEjIdKr30UcdQ6Vih10wiE+pBa1mEPi3j57R3i5H0o
PIujNXVEIvrSlIlsqspMdnS6lqPOYXPiy4na4VzRS7aFZ3DPFgfWR/j8d4PTKcVP/f8bnGLoBVXx
Z3N+qUAPBeqPq64GIlfc2aorpHy6oWBOtSubWUlUvYd2ijofLyGVEgUxFoRPRRTWgCkWApQ0+CSY
5nziB5FHWTDLJgf1p5b824aeOCcrKQCQ8sALz55Htlu1y57ssvMxEhBlDBL4nFhdHiPsfuXOMuOc
OJ1JOGmjUuLMlNIerbgLVg8mAMt8fLDWvl4LuuT2KU/nTwk29StiyD6JFDECeE4QChCbWdPboeN2
OXnJ8pFM3PljLid42oT0OE/d1c2oCyJSWZPErmSvQD9HCUTAS+sC47iSqUIK1ty6SR3AkCTAUShE
gn9mU8hw8u+HmJM/6eON9Mhl/E9uUzlybi1lQwdnvPKMPUDxG0d/4mapBJFQ0O1/lURHVtgjlbHC
r5T8qpgL9JNXIsFyR4QPKg30Nbpyq7LrKZqCGNeZ1nqYDq4RS3jJmPf/XHZOsL1+jwaU/TEZ+fQT
Pva+gc97CeBfEGGEuotZpPv1PHCpHM5IlKMe/YXn/bIrS+jJ3U8aqfkRFOGHjF8q8AlkmXLz9Pz3
+E8dOPS/LtJKLvLYcxGBaG9DJSJC+RhZUgND3I4yk0P57DyZ7lVWHhUxsciBxf4CyYIUqz+T7tjk
VWBjFsIzuQZgVWhLN8hPsV3v/eMhid0BZoRP/wSJiNv9HYTohhy2MGTWn3DpDukl3PY+Z1yJphDZ
jEKEqaVE9Bsi0p/o+YsFN8fgPH+V8JxG/jxJlXG0HVDtCdNV4qSGFwF8bUq6AnAMQcxlSnDMfCQI
AtuhK41iHTFrnEWsK/+HXqKVjKw1AX7YMvtILraFeC8MQgvgE7S0ldXxCF7ytCi9P4hIKP8Mvhd/
TsHCPo+Yh+Wp4Fde5ueXrvfG81hIo5RTYQRPcGQe2aK0Bp7phEefTBucc3v44Z5TP3vfmUg85o4r
xL6q2AqUghzEGdXO0SGXPT59m/6vxXKO+nyh0SQV/z0o0InCgWdYqgYB63LHeE2wjHGMn2sVBfO0
jp/6z5oHmEOYEp2xl6Yr0APfEKbWJNK/myuCmoWp1+fTIzjmFTjdIst5rxXcM+1jBdxK6XcF1y4J
Fwbf7R1wLX8VB2ozlgjiKQKnjBmc1TK67/te7azRcxbGEtAR4G6uwphA1IB6YZKd5cidUZBG+32t
7wm2MY0bJwfrVfbwk87Ik1wiVanEFQHLOHD1E13Pr64hkeHSHz2+AMF3HmGpgKUyrad3VxP2sJsZ
e+d39VoU3NvO6LAowcXOFH94OSUJ1+7YdVE6QDo3bp1FvnBhv2rc5hq1UBYYVRwkN1LOSv2Yio1l
tWGF8gpYpo7E9Noc56UQ89tbp6u4kte/WLq8gZnw1XKfIFv/8kAFtfbkrgE3Uw1C2Ku/I4JXkPJn
JQt41bF+e4SGtZIOOzX8nnkQFEJ6JWRaEMj9knOlGWT83gUV5Sf2AWvjNXeNLkH+W6fynqmlD7vw
7zZo3RXlNxPOd4pvG483EvywA58=
`protect end_protected
