`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
UrCbPXy7e1Bhe2BnYFa3R7+OuchA1GgOZYdPGF2R5EOzQC9j0/lkPPz72Z9dIYdQ46i3JfKLbVTJ
AYdsH+dlobPjJjQ+aUZ5JgDn81pF/sCmuGiZp+/Mk9L7V855tUjkIcTxWpi5t8FtgPiSli4doB40
sD4qHluhEBlo5lbkRkHNfadXmX8kcGuXH0Wd0L2Y1GvV3LKaVZzQe9enjlLT10R8bgwKoWLeO7C8
oKqgjg1mW1Y11CYMcD+ULZ8wO0Jfo7/cpKY5CQ36hi98rLCJcvZUO6MBflm8VIBQBhfkChd0PaCB
rXkp1JZUgR+sGH1OYJr3zv6LpQy39bQ37fpKoA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="oYZsuMfcuMInU1LxjoIH6gM6kDHGcAbdoPlyKlLlr5c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15456)
`protect data_block
NQaxYow12m+f6HhjTM9QN+qTA736rgU5mhvNIIFCLIgKjaYB33BdZlKyFPxBqZ9+BpM5SOR/u5Hk
H6VejsN+xFicJbiZhQ08yIgELMHzcdXcLVifOTM9bR1jHJgQi4u4Be6nyWIkJVoHiNF3XGTe5C5L
R1yB4keqw3lYm6DxOtiXquLSjgrflf0tveqTVtkChhucG/04ydmc3z3OD9BhnlUiOIWBXIQ0MqQl
tlxVyLhCLZApscu0A01QtOUTJJ0vIDdct5jURFyXCLwP4AKsl0b0Yn9UJCIlc+ZPpdddVDsUOh1h
gOb3K5PWV01G9k0+3j0JkFhut7z/57D7tMlcNg4ODCKeTe94m9Ws8LjQRc95mi9R9/tzLn4+nl4D
Vy45aN7A5Ib9k6RAA92lH4Cv+P/wxCmZrW/C4tJCVrOoHTKWy4W9g9jeJk/SJGjPwgGcVu9UnBW3
tWHyjVMswhjViCqH0Za9Blqbh0ak2OqpJ8zG8Hx+gez4dSO3OjDO962Go2YD1Wr5hy1TtIjPLT4D
8y54szs4bpZTAwU1fHw1Mt+SPBJ57hr7m3uWVWa1sOtDmKyNPcIVj8YhzHIerNTqDHXxtY/7p/W2
eDowkpJKoBtArJoE/awIGEHPVn1XvPIQvtXuFx0YDTCTqZ0xfL30hkYKtHyYjSg+JGtuo6Olt0aA
+czl/YdaRgm7dzxwCRBtLfFub1DY+NeHBqaa7ePROLkonCYfrzUH9V7pnXAUaWChwGkRHxUkxCAf
ipjW0yCyGiSx7t54Z70opHt8dnbX0xdVG6sbM+ygoxflyJBXiJ5+Y3EV5msE0EQfUL7SwFIobqrL
V7uuWyuDHFaDXFaXN4xUCRGAuSxDh4OzrNfdV9jtGoEzSfCkNEHzfwfXcrnZ06zx6i8qjPTkITcn
eQ0q/gBSCPtyii6E+ee7W8LF1Ar9t9C/xL5u/vOnqLVrs6d+bgbBjjxId20i2eciE5Q0m3lOHXgG
YtT2CO+5a9qJdaHeJzDC7/uztLet4rIvJqD72p/zjKhWZgdGWIcXElDJraIRdIeXZkgBQ1QrIVaG
DPBuReMmz++EEr8XNNhk2HKi7hMQb2BGu5b0F9gSgw8facZOmzxw/rctT5G6O2Z/5M4Cj4dBog5p
GKqe4o9SB4tQBsE73n0E7e2x7fMvl1/FzsU14nouHakvaVAkK7lTbdb5yu++vxzNsIBaPjV/9JvK
YYiCr/mJd2NI5HscpcGTOW7wfCdgwdOIhn4MrzukMRrqaddXAHUpAJdmJDreJzRgWCOcSc//WHUH
V6hd9DOeth3mJ4YumH/qi2lU9lPgxeba/J/SxulPPF2ROp07G71PvKVs5Q5F5cQEY/l52JiZOTiX
4WNYbSOCYMP91syxc0kUgCLr9MXpIWwU33l+U/C0Gf0RQk7h/csJ2634B5WT3p1Ef6FqF00wxRvx
2mFnP250T5rm6wSSUEcIny61OOiXauYdB8tcJJXos8G5Mq/NsMVsDGkKo3SIZItwxyoDrDf2SbyN
x/9nElz0RIns/cBBBrdZqVPzKOE3Vd7YjQ1OqzaPlENMH5df7QlhaBwaJdAnn1oXDh/IEZvSGMrU
GHtx/Y6B+gpvnoiyG32iOTYfQq6RByf1+SyaYxTanrQM6Yn/MSRyEUnkcJelU6FBeatFGcm2J8nG
/DdpG16huP433cj/aT1KgxrxYj73YkoT+l+lci/gYLCP/tbe1+x2lpQDZTwGwDb/L4bZ07MDSZ1s
lHZ6JThM9Z/WEH7jaX33tvTWI8wC/2VqP/6DvO+a1eFY2ebf1M7zNDUH96bu3QAAj7DOyH3UTtua
VQMwDALwypNFz4Ax/tjz3VDTVCre2tP8JOqtVQT4ZQ1eE7CV9bRrDZKxPkm1bhSZqL/4S0up/CWQ
AHCP4SvUHXzsJKJ69e7AoJvJLQK7ViR8ZJZsUCzUGYuelVe80hhWfvC0T1YnifJ+AdLHKtpAcz0x
FAx+GOX+zaePyDkIOTCWiY/gEKt9b6/7ts5jgUdOYQxL9LigglMs+3zfhT52TbhrtbaCBg+maE3+
L4icDHeLi/9M0S7VQxZw8HSHgCYF5YTtffDfvnNTBVRLMRcPFBfbA65dDth7sNFW9cyFInnnqko1
a6ZL5OiLXZpOg/xZ1gVpr7xzyqFktHoqYRU9KAeanRarodW+rBppI1lQp1kUb8pe3KtZT2wph53A
GhQJBclE3oUNVp2smThmNJiut7x34GyR2hp54UssUmqBm3SjKR/N7Dkh0vlJ+RU1iOFbTl2vi1Lt
06nqecRXzAVRiNQBctqYUEzyfjHoopmO3uz+m8Kg5u4lKhNjiOUSagzl1LnsKwRyEeG+gDp7cGxE
oJnCsUSpyQ61paZ5Wr6O1OhC6qG0Q7UKMXWlxQXNh9VRD6KK5/5cTnnco8HyCtt8kWm5W3kF6Qn5
HhgCIKgHY0PtgMEJWLJHV2VcmCJ8zUzjrto3zV+sJ5UE8DOB2PHrGn7mv4MEJxLYTZ9x+cC+wedx
c31s6NssLf8dpY6+Um9uW7CXVG69uNKZKhKW+HIkXmn5N/NZDq71ZBs/qnhRkYlnWQ4dsdxACkdZ
24CFGe4Qc5lDj2Bqncjq+vHAInD87Hg931zkfLK+9m+iV6cF6AzuQQmR1orZHeF4Vx31RURPfItx
swop4vc1tnW9VTbm/CmawELxzO93OoiVlztxx83DLjt7R6SugF3vfP3m+YmNfK+Yi6ikVvUysZFT
1dEGtLI9Fj9bMt9WsqhrgwL1L81//y1jIj6BzM0PH4K8uG0oI1qBF+fFvEVCd9upGYdgYZh47FMS
3nwUV/RcJj949a3yTRdpcELccakIcxCXY+2sJevrDiA8R3vF5qUn95koqdaks/MwCtTFLDml92G1
lBaZGnRe7Mn8J/SsMagtLHJLi7C7PmrwCi8zzAwmxVMBy1+/QKL34xIAcE0qiSx7mu2azPgNREF9
xcQAvL9reZISjeFiPjzZU2IZ2la5lOboW9JhvtDzXb8N/eGD2HPiDGGCcWxlc/zbj343wLexB80z
ifuMfaALNZK0etE4AYYdLOuDrMP/lldbmjBH5jtdngMUcX1LplaDuXX5dMtlanniT/nP1R47iqri
OQQeHDAGM+E2lS7r8+BPd1EwXl8ZirLU3GtTJysSdL03qupCdfQsfWOLZEAb8NmW6a6/zmQqEVMs
JZt3Vsnnt5Rm/ecmQL8pqURxktnmMPpHjJi3fFsJ+ushp19G4LXHoktqYWxR6mrpwHrBHX6LwpPZ
s5Kk/OcfWvrmgRDhxlare24DPncXuo0i71o1qCh1xFCE1Z56VJq2SHIXuaHjY9T/b9Gns8HdZel3
F14E76Dvve+d9ZzPUBHsy0QETwAxPCY3ypOhdA6R8kMQuqO+Yrm+qw9uRrx7J6pdlvv3h1DAIsCR
G2BvSE3WID1JQw3GSe7FHUC+lGZ6WpNSoxazzcxsNG5TTK7NHL+HUuliRNwiCTSD0JplfjphKBE0
7isAYcWe9RV8wYup8R4/q+vZ1YLj5W4yqFloDZnl+piO/T4gEnB8gfDpp7sQ18qfu65V8RJs2SvZ
r0mAzq9fay/LDzowfAkSUnTtG1itX+vsf6/NTfLDix9TlDWpfbMrQ3AHZDkJsMcVmbSk+gM2/C2B
NiB83//bGhTieO1ry9iRvB9spijjKaiYFoo2LHbJyKZXD0VbFcu55R+lg/GTpP4NGZU0ngLrJEuy
YFQLg78f7rzaBvLSBWLyp+DjUFXELPq9a0Ch/zyP7j5Fz+WnvprCArglCLzJyD5IzAc/1iPbCAqB
CRvmBBgCmGcjQv+YBM/DQFExK3oOyPHe/RyIOI98OdBTem7dafNwdUoW0RKkffZtczZsFDqsnmZL
Xm304ziILoAT41xnjDi+MCQ4V098KmZJdOmUDbalQKgmr+TV8Kzzm5fDQQkHU8U2QkNZGlfsJiZM
ZiygSkOAzD2QhEhx+FVkswYItEAXd9s3djHVFDy/E5uSf88xQSPS82YpBfRQ/j4gEwu5CYPGZ10l
nquxiFJ62q1ZP2qyLg9UI6X5oo5gDrjQCFuiZJdknz5K/EqPgutvOrq17C3x522879jjZ67ZgRns
f8AQbaDJEpk1hcugJXL2zvd2uXhjlRFoX4WZBx2Fbd4/Apm9Z6ZvmoMvR65s0KkIPRBLUCDo+BkN
yMoZhd5SLAzBLMMhRf14lxORp0y0F/1C8mV2nRbftFPin0/HcgPW3DhTYsZzDCj+XscFIVs/9xFs
+Ac0eCLtvdooUC3JkKtuDf5Jg+tsjnNoqQjeSHia5dyNS56qhH6G649n9QMZ3YWSdNXY6DQKNEZG
a37+Di/IUlKafUn0a8RfwIUHO72UtxGxt+i2ptLR6MCXGunoFJJlg5Mf018B1EXACl6S+U56f82C
qpz0m3fiyr0XfZzabhTZqTIdJks04Q/l4k1x93fWsa8lJIuyHoVY+XcjW+IOejxz+/0qVoM/627H
T7bznGTZNTigd1HJhUsHRrGTN5WZr7yb9z0njA1B4bEmNAyFd9YHrVaNNiwxoI4qJ2fQyXJUWbVA
Hlb5DGjpfTbm93z3AleKzz5/tY9mG5ieROYUERgGf4p0CWD4Pi4uMUW/hyWqQFDNzL4+dYUzdV/Q
SNBSjIDk9PhROfpqzk5kfweQYPUh/PFGrinaFikrLy8zePQVRaFo1u+XOxTzcGdK5K+8fhtsnL8V
fW8gEKnbL/l69K6MaXEavcndJls/UV74bbyUeD38b1Ay9YF6meGgzH9ZBY9kDe5ggms/WD/ADCnM
BBXAG3w/Ud8t/jnnl3jMQ54ePw/g87V7A4b4vfIQDkElnKnIeT20gQRp6xGEmMdZi4Zym2c165p2
Z5gmGPd5oecQp+HxB08R20305o7tQ0/TOZIgAJztjO6Vg922so4UiI9SzaGYVYuTV6slplRMVODa
gzkSuiZfvBQDn0L6973kkxYd2bdpAzpzpkbcZbKA2uUVTpoxBFOkmAdpgLrJHFt1PtUxyC0BRERY
jWmHcKlhuUYGpte7velQYPQ/pXlbJU3LhGB/156N40LMv2rUJ9HXfkFiZoCgo+kJtSKyElmO3Sn+
Y1D9okEGI7PqeJoLF+DOLH/AVze2pJCiXjMvEGONTkfDj1X02CTyMZHnTbQ6F0AUXSYj2wOALTRS
HNl9cFABbjTSP4QoQsRQHBKYpxh6Nma10jos11mrn902suvq7QaEK5u4ngOeCWkvsFiJtuUB4SYQ
2EGWVB8TrmiosO2FWoY8jSLVlDpQqpoyKvRskMVFD0OGp/nVjC8hfnNUl+UuPEGfl/yL1MRaCZSp
+7unQ+LA4pddiRx7f57DXwiJBUG1VILL7vwMJXAs4T8GZfXmCJuM/AEBhxjRh0Ih8ppt32OCyE2x
Ot48cLSXqD+yOvIN3Wdwz1ZrCpitk64LkUovzercVHIeuXBwZ5QLVJ3Wth0crYZXNtJt8F7Zm5Pl
2ex+UyvRk4eU60+z4Fb6S5DgV6ZJeSs28U7f3E/doe9t9fbsnV54VmI1o/JsBjcz1y2DfLgBNtpV
U+XFpz0BTCnqO9rl685OxRqw0a6FldEFM6pAQZiDBgMvfSe0dnun6Fo6ITsc4uVuZGJt4QRrQtlt
ByM5lsiuPlY8W+CaIAqvsOCWg16xjaKPX2L+RjRcUVBYQxOv67B6uXlvVWARIphvjEuzL1pkzfAv
DiqSnizhZRdZ710YQKsiGDl/xB99xnfXiH9ThIizguMiqcOhWB9Bhd62n9Ere9913C9iJx/utGhW
/T/IC2RG8jdI++4JzZbMhbEzjK7S42uJJyiuvvy1C2w7wHLU2OC5Ktt/gLDgH/QF0Eeul9zUTYLK
qAWbcgSQw0whQ/ITmC1Zqgiy6f59wcB/Vt72fKVNtLrAoAJS3ftxEwOqCFt8cBDEHok3EuJL/a0P
liIpCOlGbJqIESmBxvU91iGgj5HiFOaQXUI4q5ekzdujvWkXr8J2eYRojSFtHK9Phg5UHzxUxsVW
h2lwTG13KyVyCBLrI6q7WspvFI/CLMdM+biOMsOkyMNcFqmKaZN+d8SbyP6OPqXoASPn1W/Rv9nb
NRhzGpum/N5yISGrO+WaD1Fe1+A0p8Qdc5ow5Ww2JpI8phHoYpAwIAMFKW0W9q3Dq7hWyf1Zs52N
RRfuyV86T5iRkVD8ADiAZwq+OKMK+RGlA5JbzAa7xHJgTaA+qGqPMyFURMXOqMRn+4PKv8e5GV6B
9VmFgRCJEd3Gjw52cbuTVliCvml+njPnAQm6WQJOcTfY74sUMDHPyrZ5EmUNXtPF0q1NgnNipRxO
FUV3zroLxyRSfbEajycJrkTpKis+y2FHWR4SgsW/26/VUEjP4VJBI3O7k17a4YVM/y7nk+BifWW2
hup7BJtBlvVHy9aEV5yptiT1JGCMH6AYmhpeVkPUtN7ZlAXLiYCcfHJJZ/AkgnGc7xajxi3FXE4+
KTEvGa30jnC38IVJ06nKMlqtZ9AVowKKJ7EQlPKgC2JcztXe5QvS1ZNDM3/ZmRhB2YpoBQRvv+80
+LyfGON6NrxCGm/o7HV/Oxqn/0FXOr7zxbgFpM7/NNmSi2JtRazlIUzfrJMH+oLaJEmZQo2aR9AI
9XWi7Hk4Dcz3T0bJvNPa9MZ/mt8NPvT4dbOzMTo/ph/8fnarT3zdeExTs3XnCn0xMjPcj0saEJMv
Qvqh7+cN2xmZ8chH0xy2x5cm1zZjIe26FEiW9seRgsz5+nC1AIrc9835GatB4J9sJQDqlYIWh+VD
t45kkJDxQdeaCwLQX0m/PHxNsLqnr88f/wqIsUdmaY8IksGxEQMSTrBUottlCRHtHYnk6DkQeuas
OfgmazjcgrGcCwjlbPtZyH5nIP6ptoISH5Q/0CKGTPVqeYtv8Qfdf9J8cgpNW580fUTXQROoPg7H
lUQUzSoq16kaEiutSfD+RmbI1sEbdD5h8iVAa1GGx2zlk39HpwBf4LIjgvdMtFQYfB/IcBfEj7iR
xvaW8dkBilfVb+w1gkhy7ZvvLONpNgeUDFn2EIDr2Ta6Wj6bEdKctPsJo0Vun5vyXE1lbIT+VjLN
smBvcO/EqXjgCH1FW2IreEGZ4XTl8efi7aOYNrDOtUbR3DxfGdpdLanvOPegap2XicD+Jh7hkLNy
AdRacXQgzGF/hAUhAYxhGt45opwu1/BuDvShjNpFx4s91k+yJwCdyTs3jC5i3N5gosjwcNMY+iL9
loaGSb9RVAj6ZndjMzvfi6RFUJ8Wv+L3NK9ST9jtGMuWGZDPTaJUNkFAVkNIal8cvADfhiw73r28
ALniS+idiHC5D7IWgnfZfs7srFfsRXPsDWYuOME6iNLmiCdK2W1Bxez/BtGN4GVcOw5ilnuV8lQP
e579w/F0bGBDgCmybtXnXn/T2Cfbt8A0YIC6pMJgst+j4PsL5k6tTf4FrVkX+bNPDuhy/h1LOXju
NQqKd93y2gC12exGr3nZuoi68IyTrE42GZjVTAzBDEPVqQkIghUIK+f9DBV2IBTerrcMLUcBBGjX
orxB7ZHfoXcDnJaNzKGzkTLR1XDuy3tGkFlJEr0myDRGQy1d/MGbyIcvkC4RiDOoUXJLXZmzdOVz
yYIDpz0rxMZCEQmO05pjjDp7f6VD2TgXIZOocyJYnf5kWE0D3RSNAjoctQmZ6fcS+/+eEt4bIuHR
UpAbMvo0fWEDKyDKcNNICR/lMpENknYvIEvxjIiAPK/f3PYLePreCEaC4bhbOjnU7wN2o3Ub9opd
K4jTr1OXZieSEz6YhG26On8RajgOKHrnXFqU52hCCArnaYpRSBlmer46Uc15KWWJ3dPDCWf5d3nk
5mNMGdNLtzYAcWWZGKQHhHEYvBR8Z+Y4rYX7tVVcoyVys7cikwN5x0Ypsg+laTCRDiK87slPe1yq
MCHy0AvK6Bf8SHX41siQKeaYFB84x+zg942eaKurmNe0XLhW9+9rGGIRIVuCzN1uhgshB90qrVtn
ExMEMNt79tweInGd27PcIOYXZSY0DIZDi8X8UWobIJh976Kla6RXZE3JB1S3/H3pLrMOcePwI7Cu
+3xauaPFLo0lhOGurqUjmb281qei+aClWP/1VJiL3wg1N2h9EHxQ+SYclVm8EnSEqJ8ZrLjTr3Xp
fMKjw9eEIDhpKr2lLpWo5RoN/OgPZH4ojwfSGGZydqyDk7brutzYC5kBOGphDLUg0xQVLAryo39K
HhII9R9vfy9vLeUJMhczfVaApDD08tl9ON3vftUg+nfXcz7S2tgiJ4HX0SmmsF8/jIjrEE67zzQN
JRHnmDV+apKPa1tDBrvF1RrSGQgNncM6lKK5CofiQzUMR0S0lsCjlj8y5MupUcGA//qd4tdebOhx
CkCCfAIeu3ZAKSAlqIUp66tgO3WmQ8C31SRc/W1OoWMw4nmOYLbYSoQ36do50aiizqv6joehfTsd
YOKB5izDXfKLp6IGILwGbs72Oibbq3NTZfwFexZ4mBwvFcfqel6M39TblZ/DDsvqwHUMtv7k8iZ6
wfWBv44MNAg2vZwg1t8/acdTbXhiJOqXS5zhegaSiqFeF9q5Y3zEIPmiNGjJSJbJCe7VWWG4NBD6
SpoikeylFCuCkdmN8RZVmB9w9m8p4bX8wYT0F2A40NLDzn5liDx4+4uoPQ7uS49pvidXuZuRKx/I
eM3+2urrRa7rtFj96uPytj1tYLeLZrsllLW9wrYce8scU1xfecfuj23IOdN8gGmVycruEHBG8Rwn
oJplkqfG/9Lhjqfr6ykaVtz3vV68WWabZ6tZl4J7WL2SfNV6mV8/1Atl1SEiNUp68enhNxU3TBvu
2UVwjP0M6LvAHc+jHo/8ZcCVX+lOFJooole/sgVEuMtVzOTEKPOiVt3qLx6icOkNPllG8iwB7R1f
DEh8mmu+i44IYa6uODnjP9mJ/sNEPpeLeqyV2XHZUamJ2YkUJpLDZ7GqeJ0n41/Rt2vfLQtd69+s
jGw5jHZF8lN9FSWym38N9tppz5iZpiCh98abLmpPB6N+nAmzA5JukONEnoI24lnjXuxoTPXYsKaa
OfvoM7e4CtOHliVEsTZ+R/P7lbc/t+lnuB4bHpzIVrK/raYwPHEDh/moXqHsyZLQ50jFBpMyco+4
xWNd9odq1LxHpNMh9blEI+68UwW0FOtCxWKt9HtVgF21wZA940wBJCkCWmVy16oHTHH/zHILAjS+
dGdAdUJAFixKT7jPdkmPQa1JLtSh+6VrPk8kDBluH0Lem+Q/iGPhZrkJmPVLgH4P9PmRRKj7m/9/
7Jc0pdAnCQYOrsM2JuS2ilfpLNtzMosNP2sx13QRqkW9l4+Kwj7UW2Pka/pY7Qh5MwaVs+ylyLgg
JaDywiAXlt4A6dOEAaQvLAalfCzJDOjyhu7B+ecsZd3SLv+Nx5KUIqWCsNbvsrtNvYgZG2N4pehM
y015t2Zzys/C0mwtlzVieEKmIcLjplusLXpfNgIancCkUtRB3mgTZmnsLjAs+5KD36swsepU3uJy
CaswCMY8rrnOcYwBCqaQWHHQ2h/cttj6NkmJ6qO5es49L26N5EHRCGHispcPLureZ7uNvtdvzv0K
GNjj0ZDffIzJWN66TSBLbK68dNBUcyz2kcul7qVQQTdJOwsfy8Pm7zvXfiysZto1zM3jSVl5LsrU
xXhLEWPHZpNKtllcEUapmDOm4lggOAlS35Hdfea8vySwliI+cCI+9Bwgm/xO34CwPVDdHCHzliKa
HTRM8Tro4EOKDW3obZ/vzPXKguyNKkJffPi4FpqSf1kqPQYSvb6Fz8xqhHPvENrCZSYj7EPngr+F
enZSfwWK4yAUy7ceKA2i76+bwCZ1mqNHnRbrCUlM/zUdH2exnK/jWJ+VKh2/Rg52hMxJ9/1vcOSr
VpthOSH9p6Q/gwzbhF9vkADOgNGTJm7derDauhBlcrv5FOjJag2kzxkkPSW8jQnpdcm4rqJsRrku
vmEK6/JCSKHDWXTktdwkbj5wMnaKo8Nsr46cLOKfVWeq8HksG1c+Suh6J/cPMI8H85KFsdESlIjT
rBPT0/XDNy9qOWWyo2+jR8jtzN503p0nAJoj0z/2WuwMSm2ylVSNFLXCsEizqp63QwlqZ0z+0ux8
4S/6RaQrE2YelegnZ9vf2qDu7XWDLeD4vYx/R/K3p9IDsQyyNG4YztPW7XkvtMRKr5r/BgFSlw/u
sxYXLBlOXcxrkyCVFqfRPH67wkDOZbIZOQCcKUFM/9/HItquFAylzDrYOpu1uDLFFi+zpHjGuzjY
BR3TE3AE5n3cfvobV4cMaDyJxmGlfk7P1Jb9n3vzr4esrUM/w6h/DDDfOJ1ZmelxrgMysgVdvPxB
Bjkg4KCQXU9gtfdkw8A1ZH+f/GeJHBce1UqIjhyU+jIti+Gjs42+EJb5nW3bP5s+ldtuh7I1yF4I
QvmRslDaCkJTAXwmalcC1G577QYEYiSTcbpF9dr5fzvTKCJS9CChGUgtIITMKihWYqBLkqsbmSYg
3FphIJQGx/QbFPFv+PpAS8h1pbpJvCwjiAvoTcHc4zeGaqdkaHmmwRD/KK9Bm2w4qAzzPLFuYlIl
Pmp2E/YZQ1tTvnupuawpQ84MAEslf45aJ751yBpBPlhQq+kOiD1SCKGqWN9VoYxxm80Y/PvZspnt
5VD6lrFK9SYazovNDUzNQpj8hk/n6hKpc50284H3T+ord00Ms8UjqordjbQ47INjILOwa8tDD5xq
xnS+/mfyKSz59MU1/hhVn1BSI8tWdDjGXOgz+n9YAaYdNqD70L2yEQSeK/95wYb97e1uPtcXrPrS
Vpnm98Gwqxas2aCbmV+7dhewMAefMopwkSUEljyfGElApGQwID291Ay7dCvt2lhKtMFar/ElpyzB
EMU6pisR1YBfDmqGN9gCjdVyfBlEYsTdOU8bNaZ7XqhQRKZoV1wNqCdE7DuPl1F7haX3yhxuqMh5
qxLoYLnWquUmWkQ8GM+qg9capgCC+kTGVGBqJfldPLkqnEwwS/4fBMNyXSqQe+JRXDEiL0n8tP/B
p3RpKGYG1EXK8DGIl7VLdilgnQlR/zSL0Z5cwPk58JncaYa3YfZp66KGxw1CXiCnSeULAHWT31cD
DBhch+LXw1vIHbhAi5TDj8cHEaG8rBknkIlns5zV/Tu/nOizRfLqJO3VMqrUL48c0IAvYRj923Q5
3WGh+PdAOD9DVTjbXcai6aQLAGg+TBxWRV5otDuEyKqktS8N+AoJ/voG1DkqMtOL5dilYxokN/VG
qki72KeYyUjP8J9fztxUu4vTTgJMwPuQNXKfSF2iLuLA1W6IqPSt9ZfjQmete66fuV/QOe16gCe8
X1AZ3vjv7Rgvb20GhIO5JWAG5e/MuwVRMUiOSdrcpRwnYMiDSfPfv7fTkcsoVR6fyGRzH01nvQBS
Ela63G49EQftnA+70QSPtzWjYQJZQZNEiV4Wo7a7QaZxowcwq2vqz+I3fxpKWtXEGSgahURBp4Qe
NzzfhnAZyRpfBrAGJEJeDucOMoWh0K4brxlAA6nTwFtVKyjAxVM7h+LYZbu7mrmK//ifHzDjKhnO
5Ec/2svsHzWTcrUz1iGvtvvcuWgHqCJZ26QQ2LAGHf3aL7IOG+U4Owlc1nQnzN2OPEeMd+1vY4hF
lVM11Z+oVDaQUFVzjS88RGZ0k5Ji367aHs4q4iczdVxuzb+VmrBikM73k5yneHeKjSbs+mEid+Z8
TvCLQ77qFKff7C2AEYhzI8xm4TN1Z3BklrYpdona6eJVX6DsxjerxtLkZgjeTJhph4/OAK3gQMkE
eLJNMJdK1G6oD58sv6p3PhwfLWcbYC7+LQjU1NJJUHQTdtnJDc0+J1Ou+Wpolb1NsPKM+OqhNNrW
0E3jBiw6jTPqUDPU24xhu8Hmn0fGoJfP0ftYfz+tT8cr/HctzK6DZwSuGl28t8pAZIcQSkiONJqL
tN3IipGqQU7SV3+DwM8heAj4nSZp3m39cHenfUP0pQU9zKZHLpiXXrhrJyAtVlRKuYvtmaLSuiBH
RE3TgaEVcppNCdNbsEVlAaWBdpZHBghCSSyOvVGzxPPJRj7WSZhq5u1j3evwEcTlImKFEqNpB7jM
9wa8TLsVIzH5DxzXCpcYZiyM66/jTTiW48Bsztj0DVZSw3hoUrk1IWIcluyr3dIQre/5dMgyGOiK
Hb+btrVI76mO8l6UQxWSRs02emXyzDpXhRisv4zewSNgfge0Bo77D7gE4ZQegD3QNhz1MNvpd9Yx
Zg09SJTF43fepcT85wrnD/zlqljBjsVRFNRCVsfd9hgwlxrhcVj1033D4dE0tTm3CuWoEA9iRssR
nK5/4YmeejW0GoEcXze3+VPMQ4dPU/VSlACQ6qP4TTy/fQ59lwiKvg8OBDWjK9HQlpftUZuzEzOb
vmfd8PSeRa6J37S5K0DkCibPIu64yTte8cx3lEHbOh/NjfcIBq7LrQ5+Zt3xl0l+9KLVdAtSqThi
aGTyB3w3AT5/Xht4MpKb0R/m7jT3R6aIEFCR9FIJwV+K0dC0S6WjWBA5ehJ+HYf6NLH3LRYDnrLr
bVMiiorNj2LgVm05xIWM7/KWeDgcIOiiJpWQH9BTVWg/rWwGELuYLPBcpMVJi2g3u1DBlyHNPtOE
5Ny28+etFS2iYlKWExakcDWFD1JZ1gTBer65hJieOvsZGYQQTb6Qm1uZekltWd9N0wjUlNcHGBI2
raSKYqPRZ2G57hGd4EySM2xglL44jFjREMmru+zqyODw4MSNzee7mgBsDYdoDrB+nHdEdy71TwyT
Jcq0YqVvQW7ukFn/8OnVqK+0Z89fx5RjsCuV4GkQCbByXv83GTJ2IB2xxRzri9zhMwaXm+RXmiPa
mleVZ0/ZVsXg/vid2Bbv2IjuZhoWEJKtXY6Lv1/eHyYx56H7iohoK9XQbp5p7c7QoCLy//ykE7j1
ap9o9hP/2SOJrdaVM5YrkbtNyeXiuw4bxrTdVeYrBC62m1zh7qsMIJ9QI6EIhpEzSD5+WrlRIbXk
savNtR5bnqbV0dqXjKmkesyNzRpdt6g6APTHzs5NcmDbhdQkLckxvmBkAMidItZBrpPLftwmMExV
dCzGAwOSjiPrv4qw0fzavSJ3IhmrTuIxdqXssCkEJ7bwxx3GLyuUk5hsUPRMl97HIFd5vmf8SxiS
zJ9bDyXV9PNeJuDYQhMpluyjdLIo2MYVJvENX9rdyWXN9J4ZeppnAwYpERSHMBeTiVuqLfu4qunb
kppAsjP7lhPyg9ol0V8urWhJEpFmOlZxkiROPU7llZGiSmxXWV87pwrtCGzbEXBKuqhVCz4G7DRC
4CtsYfCoWP7WlS0Uw5omtAOtipvWiW2aLbK3D1f/eGyApwvsOpKp07ZXuLiFaw6grlLwaokCxlji
PLJELJ5bk2USILBsObKBlR2ZpUTaof2ZWX97854NlgQHmfP63IxSVFlDR3wUKi9XWTauLEmEALhO
3qbCLNt/VOnxsrDxxO+Gc9HG5Yk5aPFEp5tnbPgxRKdp+iBuCRb31XoJ94dqRI28Mzbhj3VS2jQH
Y6M8ZjwdMJKbvJWCzoF+qfhppexwkV8teTXBONs3S6LXIWlAY7f3Ox+TfLhsCTAVMp8+s55eVU5D
+uY/6RMVYIHsZHYpLi88hpoMlmjyQBqhFCqMg14Pi2QUWZQ11q09kGxriXqFZJJCxkgH33WfxuBG
I2UeYUV+OkpP0z9jqsurqjpe1QBp+JF3yMqp2mp1YNXBI4GE4AJ1RcmrhXmyEmpvQ14Odg2vSMt2
KV1HRED998s1mKs4vbQNfbUUMfznL4Vdh8wevKUkWz7uKOytbxp2utfr0CCxDQq4GtMMuFv76MwW
NPkvx8wOpv3T6MR29F/gyA2xNYoPy5m7mv6UEBORjAlwWVj8kkmY85JulAz8xKHRSw/ZMJovZSRa
clyLOgFplJMdXVnXCKv+LvIlbSW89FPJFe0Kx5AgE1QNS+8SN8Sf1Vvrg4JtZitCU2cq6YSzv6TN
P5iCZaMrWvu/GpR+zjzzedJ78vDWs4cteqKQX1lvd094z9rVpwBewsVhpWOWy1PT/ioWhygU509X
JCIBIycjnLqjbkbfUhQuMVO21SANmDXHe8K3ckVsQwO6dciesXehham/vXk+xzJcq1siFb4OZpi0
7k8PPwJU0xhK4MCq6n1wRyhLXAj7Hxzl34QWV1QFtPLVtjomYDUPZp9YSUjRgHKoZqLHduIIUGiE
seWuUp0FPC/vQFmaYKz2OLfYBQdzucnjr4Iyh+6NE5RIMCglo/eZCZC0QI/0Iiqo0nHq7kQRDNjc
d48cUwZ+IG71gclBk8626caHdjPRQRA/BkdTAd3aS0m/UPK/igIUEGsBm2nBLAqh4GQv6sAS2XmA
Sh8X9eRn11TQFBD7xOerx30vMZ3aKt5yrfnZIko4TGaK5BZVEhaGkRF0McdgLGKdi+utZAWikB51
5lhPtI4tPDEWScq4tUqhrs8FjKWY6kl78SccoaEWLuMuLJcSaSsIG3qWTNwf+EpmG50g9wa6eGwS
f/S3KjhJBHIFB1SFBy/5HDN+HLptmo5sG3et+SjWGpNsoFcri5qhWcXlU+m9tZXa+MUsJD1tJeWK
7DM/0laXRDAsGRyDOEmkiDBBFfsa7u6drLoEucH1cVhnerFyKyoFekBVBZiP2VxMj9lZZ7CAGG7T
4yO1HQoVvomZ+YunymB1O0l58GkljImA9CoXjsFMio/ZlhmoItrf9otM3YfAviXfg6YNGGfKWpPX
ekyyptySxSbq0E1rAPbSCI2bCQWb4duLBD4rPrOyggtyQkZ+q834M65pstPUHbSH29/cVawvrskM
fsvp4y1yJF7nQotWczXDjaYPuYhvNv0U89mj755BUef/FYYxvzwK5LGzJNCVagP5DUmhxSAAQLwp
SLIiJoXu6nmLAw11amRhl+UEgqTBUVgsPlf1LrwEw1WF59mIeRvMjy3L3y/i5LTqpUxPN7Tgp49M
volCUMwf6g11lgWWf6jmQaPelQQctF1V2Vb44tagJR73IC6hFmWibNs86WIq+nl4gGjUcJ3RYErk
Y4LM2fEm62PD3kvx99A0/HD34aOoRInOpEfMv7lLplVLTXEM9/n89AOEEZXBNcRGYsZ2gQr2jnQD
lExMwTEfyhMeJxyFGstHET0FgRTV3+vadyCI1t4NTBIY4n9Pw9PYbv246F5SMGBPT+8lK8PtplAx
GpE1Iutm8Oy2HHLIXW4JwdbCCIVrol+vfOUsWFKYO+EWEd+tKhTUzST3w3qV+gOmM2i781+/O8PG
AnqxXVaV7ko1CHR34j6IPLv4cUaqiJqQJnHY1j65YxbUMzAT6KdjifbZZ901XS88ABJK2mZIGwv9
fLCxhM56hGR0d6hh3nezQLc0Znx1ydLq0g1fJeesr6XACCD4v7k1gkbICOPzYmCRqsyDeBAwSXOH
CpuTvYY9T8bM+yUkXnyh+CyQlv5qkIl+hSj8gl5kpmjzIUTirOGJ+YjYi59NM4xuTCRtWcazcBOB
/ANY0isnDQoQPkxAplaGwJbhEOfA/N7uiNmTPRm3LVFptMHx+pxEAgsUs1zU144KQf0sZX5P02el
w3vSWaFywZKdwXNM6WxpXS2clebA+Ecs71cngesdOee7IJuXUjTVdzH26yyWTufY7kmIOrfWrWib
9lM6tKnvlvZVpsaqm4L1VRqZ551wt3HWyKRXrfj4jAqCeB3/Z2IbxcULmVfG7HsWCoTtqrYPihUa
/PbxrqiduW8mhG2J8JPDAjTEnNuOxWnFRqy7Q7KMt4NvGa4M5bzzhEo7ALg10v8nS+YqSvDpAcyS
8Z+RXU6E8HyGJ3LByvXutwgDa2pLLOLWIXMmQjcxCSyVgSvtojiQvtrYBMbxef2PuyDnx0qXxKma
6fvqJChKFwJ428sH+TWVN5lbpUA39pAmUX65H3BCdcHFwMs+L1fuWRA+IeJJZtEQjFsdIUDoy2Mo
WsYPdru9rT8JevbCNycKRUWQq736c5slJ+35MaTTwYkR9JhHwMisJma+hcCMIJdjoc5sYYYMZke8
XMKjvpkQ92HcXZx1IkB1S2oKIvvBO6Z9RYsvw+xQaPDUq0UeZTr2+D6oarMcAABxVIY4LUAtR/e+
H+VQpuBzsx5DU5wbOW5ATMZ2hN0F7kTZwvP4YHhLxsDBuZfCSfCQk8Za1ouyT6zC0LMSLKicKN28
4Xp/7ux95BYZpVZHMv0i7zSeVNdmMZeayK+P8V/NsqlV7nGMZH/+SHtn0o1UyUPSK+Amw/x4KggB
vEPwkSRF/Ipqi9UcOZmk9ablylX9+6V/ntQPbsw/rBGjLlFzCupld4/4taSSIy+IknwBeVlvB9+J
aghO0zMmRSqZTHC/wok/VL0V9Om4kKZdz4o8QGl01dSU5rKNRPBQeFfqlvwb+X1KKzt7+NP/j/TD
WEC0PhKeJVxpZb2BioZJpxpXHXaqI6mxxnsDSiB/jojyz6rK1iqYeGaY9aItuUInUOvHENxn08T5
oxJPQKtOTJeHBekDpRqKxh4SQBPvkTQK792HywK5I3IWEjhfDDtFJlxO4UrEOqTzpI87VQjcuYUW
rH34EqVVrJJkmhhgyzmth3ev5qtAYKZSFVR/quW9KLHu8rOP1Ks9y1/sr6aCXL5hOXytGXxOdhUS
TNs775Bf/5mgQB1rozW6nZoa4zs7BFaRtGNSvOvAdHk5FefG1L+x4XF3RYxV/ZKDkRzNBEuvGeUs
NRCb/7Y6DId1vtlC8yhbVXVWhhyCnu0p0DYTedx677ctRrJq5ThN96VnxRGAOKc3wjciB307TBTB
Q6uNIrTey560BDcg1e9vuGVA+Wd8xJEMKmoaPeTBTVq4CM4nGtmwhX+gARf6CWM9iHUy2OHd9wcp
Th8QAoyb9oKnuOfWGA8JiuLjE3w+9O7e6a9ZuPrqKLJX4XalSr18UAKkviKUGexAtVdgvVKBZzFI
AvDYFoHriN8Th+ygnYNtPE5IrpSbhqnzOHfbNhCyXcFSXt0nxvYj7D5unaq87msnoRRUGPuVKykP
D05G5ze55Ra3Q1nIJYX44Gjrt9GUdcNXuwuo36CIw0rqLjq3NkDFl0QrS22fpW1FJX3dVHN3o78C
C2WNITb6qKjN+uqwAaL4TNpciJkBbfMrwcif0cfLIclO0tUzxKyTxoft/LOmAwZKf+LKmm+8buaZ
eYc/f2WYQnZ1UklQHEGkDkzpClwJQV0v8Z9Jickcr4ujudFKF12JY7AB4dT2ptyKgIpWPsd3u/mZ
88QxlrP7Ys1Z+uuj7ky4tQgD73hYdFcn1h0b0GvmNhk0Awv45wwqSuZSFCYln/zrNR3ZSICW64r2
dOd9mCYEMCYM3w3r1brAtazmDnUloVNUz6fbxMzitKVitd73qQbaWlla9Q4CZIkJVzQkOX+GTawB
zQK6B34mV83aZMnemSkuC3/HRoiWs7bX5dsDrzCyRi+JESzBSxMQKRSeSJFup/rzK09hgMdVqXjQ
ayq/4sq+UBZKoaCUzZ3f6E/pMid+mxpzND8/n1Gix8WCrSGcB1QYwQ/zrypqsrSdgryeckKmM29F
+jj6wYh2qgA6ccouSQf+LBH0btEqcRwE7TEv6ugJ7bzdCt8rD0pM1Oldtb6DRW+6Bli9/Idl7F3y
kXWLZapy3nsQihYzENDH0acY28GwJSnbD6n77+6gr1SZPpIkL97nHeGdfqjo3KNZEt3o0RHOUr6z
uv9aPDrtUTwjA8Mtbx8cQ2WwvdX0f4LfrN6tk8iw9+reUa5iYKFG4hNDtEDD70T15Mj5qch7UeSN
XIKMrLkCdoGrMw4V3ddzeDgYEM4zSUyQhDd2QS+32VM3OgNRTo6BRWjfh0kU9Uv7TDSPZj9ahnIr
gTt9Ol2GGXM1pKIRMLh8G1QI2kjO7+M1Ypf+nmJ22Q2gcITXOfsSbOKivxfsUzI2CfSyXpoivXpy
LeNmpRzUzHHdzjiZJkbWzEmsHTswM/YTRFUwfaoz1wn9FudJod2PsY8+eaFaxGzxCAPrxYpNL0A3
VWC3YXUShT5LuE1CH7K1hTzJtfEUS6SwtCuhdqf4KG+aqsHzrCsAjOP8Yo5UvNQDFDdsBBNZjulV
Cz1xvQTplq/ehdofaV52N1kn1HzuE+akAwnsjKBHgEvN0Cp2f2N8L1IWSGTqumyAcwnnG4yH3CVm
4nj+e5N5KOIIZ1fLHY9JaePHrfFlWiNOIrYcQ1TakDPUMSPMGA7oxtfGySjMs68/DWlnw4fFe0BF
FFreo7nuNbAy9guF5UJTFKwFrHWpk7eYQbWRSdN1oZdTIaUCaOVF+AZ5Xx+hy0v0JhbXIGr+R80j
uROcFgMmhJlcErMqGy+9Rvq+Nnk58Z2TGwUiqqYcyclqb0zC7Og4/Km1CDDpqOaGUlNGqGgSyD4e
UNhPRMjtOKqHvU3dGr/NJbtXqzGFSQN5V38Xurfl+WH9IfAh2tlUubmFTo1PzJtHzFl7d71S7+dJ
pbezWQJcy8kKD2O2AD5fDuLeTRm16YxKo4zwcpQOFcO3z4yntLBPFFcPxKohKvcACoJsmOwaXepv
9PpbjHu8+vJnnVkmqvvb1Hzz32KFYsXutRZHV/qjcvJz3vUt90AqAecdsfNeDeBtSgZtRbkKIfiz
9o8TUAyVcdQA4Yb4oWnNOgK2H1IgLUzGPSwA7ZdTiujx/omZlz8Gnbh2MoKqadEO2tjtPFPNK2Pr
MJGDh3th8IINQY7nJKy1V9tdUyZmE1mLEfcwTVTuhArJaAvU1dRP/ZOjDV96RQiKz52HxmZIP0VY
H0BJgeQZ2WY0XZ3fZfx9rTRLEu192XfPozDWXVYZ4Wc9HIVqroS+IDQ6TGJD2wADtT9WmB3g92Wy
tWob+B61LaMjxIs62OsOrsl+B7KFYPUu5Ax6Amr+fX4GEVXJVhyQk7AVQeBAUzSWSbHETJ9nYDWw
qXpLYL4nKwvnem5cJoj8rn1qR/+H8u7TF/W5vLE/+rsCMZpNGdmWH7+iqPFPy+OZFvD/JJQUrCOn
sTn6t9fVVNRoqgQk2YtIpNkKqMcUSBPWPdKtk08/zbvmHnMqmafDD0Ih0oneEmcSUYjvlRL9ZTZB
9kG1zN5w6ahYd3x8odBT9xs+ZwLy1r/9IIBdflnwPhl0cEW/ChmaFWKpO8A0QRoCpEOpxTGwklm4
vDQmgEIuoSlNZl2fzWhf1i9EuRwza904M3SY2EAboQEbfR0Jw1fxmTkW8hlrT3JPphebY1it5zO/
h5tG238e62dKXI/kU41LyEUBZ4TpRzgaFcERlJ66qiZM57t7jqyI+1JigU63US5djoTb7sCTjrM5
URhiOhKv0fX5PbX3GXI7zD/naFMpZztcQg8uZOiG6RreneUsF2qvv7gS9J1i30eVS+yveCeXH7M6
BUM23MlubHMwC+zT7O8D+IKs89YBjlQ6xA8T20r3H/lPDbbQtnt9fFcvIBGu4U56JyA/pxIettkd
IODWP+a/TOvcZuRrocKH+2RW9H/8ToLcGWCRll7ThSndzih62SfKCFUuMZbl+pnWZk9esOvpE+ZH
TFaX9cpzL0vRQJ9lcli+rmHQi4oqJtNfjeUezFQ09cft2oQsfemdUeGwrcRPh80LThBTYHRpnnQn
2eM+RU+LRj+/IskUVSFrN4p8clW7vVvT7CPBgeszxX6CDIvYfK5JOxRhG0ECQDHtovJjQHGsg5Rl
50xx5sLBhKWZNakMLKBWhabOnQPTkgJdMKPC5Osi+u26BPAQyDFrsQHQ/avak72GGCySoZjDHtoq
Lh2sQZjIeVmNUkf18YlJF5Rc+j+IuoY2VGrO0u5pKjbjhts6Q76moFK5+vf+o+Rt8iy21g44zT5a
1CdglGFGCnX6l1sOzMCbqW6rtpHqZD5WOXAoKhvbQAaof4aOTijNHdIPmnItxeoTOUGr0vy/w41b
o+moZqruVVvBxQpK0QXuET6liePmx/fm/ndebunxemusjFHu90B8cXFwWBUMNYfRE/XrqapjlPoz
6MSuzrS59n3MvD9E1mgFJCbRpUgr9dPpSGDY8LPPm+4IxGOqEaQeps0OxqotsNY+AtwTls/oDdje
cIW5XJ6mpKVNUDWRwSk9yueMifVZZK9iiHsQvNMU1Im7XRP2O7btR16Su/lunlDSGOd3Ygmp7SKv
f6StFR52jWQi8Oce6pHSdefcl2UhgR5HcikWJ/RY2WHfxjM0j/kBqyxr4hhj63qKtjt1EyQ06GCU
Y5Uoq6bY7JbvRbamyCZ4uYkHbIoyBq59QlCuwDiPCbOql2zSjCNCi4UNGUw8S0yw+20aSRAk/WqR
cWY5jjwbBI8th6IhKEdfNTIueo2rBhKpc6Mgt54MhoemZxTVN5PtoYP7cAEnTv5xeUqXgIxwfKdM
ZFc/mt4jxU5tcLDBk0vglD6SG/5pw/nYBpX3NGZG46thiuhLEUCLJTgepEOKVjT2UgqlYo+N6Ncc
9lIOAi3KgIU6nX8QCQMFRE5hLc75YuhxynhN+DQ4ndLQXk5Khv7KPnu3wY0wmJ3VbIo/W6bkgcCQ
yssyQHTt/lTUs5X8o3XsQsrr8+hE1L1e7KESfzEFMmRbOIARJaYaRk3ZvaYBcQyUAhRjF//yBB6t
FACzPmWCi34O
`protect end_protected
