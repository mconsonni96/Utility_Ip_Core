`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
mQ4XxBmPtIavtsjyBcuwjmp5JYqhcJLSux2qfaQybdLHb6+u4XJb9Z13KFdHfw2qc5RW29mXqBjH
McpB3CdPxbHyAuKqJ0xPwp2k1Hh27aZ3N81QcmeMDmB1gApWdFZZ+q7Rj+C1BCafOvvFV94be5Mz
rIEqoSD4EmtNok2aFe8B39VocHQ7x83Gm2AMYYqNqtMweMXoipyPxHoh66hDa3FJPApThALTzbCk
5lt0hbFleZBo8DUbH1+jAEImV528k7wO90Cr0VVRFLWKtHN7QXIU8O4TL3DnHH++z0wjvYv+vabU
r/YfPNUtcoSQGflmcg3Hivluqx4ApAtLXJLHBQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="v1KjhHvTFnZsAPf738Zuyl63lKrN9ezGpFbzO1wmPcY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12816)
`protect data_block
8B8test31qeEfgVbHiFDasDBiteKafNl8UF6h2EFj0G3wwVoPFIDjSWBo5/tnebxgwLM3zS8rni/
yEQKD8OTFxyk4Z7aTHD4IhqaYhPIxF/bLkw/yeZm8fa1WnCwLhayO9/ZoQXG2YX3PLPxD3M+JLYg
+N/6CMFtRww+y/5tcLMbXjJtHq19QLaMcW9kSe+gDRZGTnlDlXsrbZqydGBxWX7bjyh9ywlmHWPJ
FpZFe2dXA1/m+X32DAVhgeGsm8slSlr/iWKXDjAHsY8IuniTJZCNZTs/XGlJDrgPWPS2HRwbWs36
OwIcxy7BMyxVDEhHt7rhSL8VDHgatkJZ9edhbvqRCpSv8XvcKc3VH/A+Xmfmi4Q4dO1ka+B00wcl
/QbKk2H2VhcjZpj1FaqwZ7wPHMyJcFh6veLnbOsx+ySheI5rsWvMtUFTrSK5YZaOkuPTjg8K6ZZ2
80TCx1njeWxB4fbYUawvDyO/FtmMq/5y1gAsZ1CK/VDzK+cd8E29XTmOr0QCZljXmEw5moha4De/
y8t+zS/bkIpoIUzUSe9PbEkq98uXDSyqAGJwTWAeHkFz+i+VUX9i+Raq9BtAJsTuyziXKioEIEG4
yaEvMcLKW1s1uzUx0+hueP5yEkluTmZUb1a7nXuwFxt1GVuRywePnvPj8uXYyOIu2iI2wOn/ytI6
SJIZ8TbuDCwJBusqTY2QMiW/TTNI32s1gr4/jGHhUalvv6CNEwCNtAKtYAU8kvWGxl2UxYg2wXbS
xK9zNILFIpOQ00TG6Anvf3D0vR+roA07JCwk7pfmUpBgW/d5bfo31hgrRRNb1F6p7yN4AAfnQXeq
k1EqwiEk2c+ODmGN5QUVJ0QwS/fhMHTv94LzHcgBiGJWkXnlRYN4DfbRBhK+isz95GBkE6mTNl4j
H/mb9fJ9rQeR3ydWVCBzZ//BDzhizVflp44qad7REwvU9UAO5H7Aagtl/kPmz2o6PzZ+9NrX4TG1
SFiPXwSURQToQtA6VDAO3r0uUmYrO8AbF8UDVukICiIKDZ68BdmCpwqcn0ftq+YdHYHImP5UWI8y
zEZZ8QTB18LUpKvPBmNPuFL8DM1h9s5I8CcWE/IgAoy3rnXKeKln2yN+eaDMxUfn3WMpxr9GUAH1
bTsw6qXLMYxuQcHpdFUEE10oL4Uyp4398Fwjqfp/HNf1/tODdhVMkXfdwPaRkM/GvM/4ZuNujLXA
1mbVo3k1xJ6J0I9IQGbXCuptoj8z6I7MnT9tlyezd7UIs1O3HloZkZI6jz8XujvQWBQ2xJpZ1fXn
pwK0niUgaxImNBLFr1RZ5nzrhPiI0rZl66d4INQ1EOPGLLUWnrzsViBpxFCHfHY+j4Qc2cMDkEpJ
ApZUwu/wZGSoxrc6gcXd7ilHob4GsY+GAsRoQWB8+typnCXxlxibD4lIMkoWsz8PdWeboJfQWpTN
3J+tIqbBNYeRx8K2vNW0vM4RxH8zB4yYqtsNFpLDTXfeqyMZG1kVMtYBYtyAUQhCwVTNfcBrC0j5
0bAbA6rOyvGkcl2Aw8ECBxt58XZ2EHxMI+1sPBkl1PRDqiVzAe7ONYPmDX1At1ssBbq0WFpFpTy0
Lom3Jmc3Rrl3/1pb+8SXjuLbvWjYfHGePLgpEU1o+UtGErLoJatYoOfwaaRr+wO6hjCLGhNiTIrg
L8ifSn7gnYmME00lUon4LrJ4lb3U483VjKDivOCYcnQOYmUVdO/AB/SOtJjcc+qXT608A3SkW9dK
V1qAF92c2BkynRXY6ss7vlVOJY/jk0ESi9FqSeQPuooYZLyzjT256IoQn2GDf0Kp+ebBp3YKnk0M
wmQE6D7UGkCUs3SSNQZUwNPxS9hZEs1yApM9Vpnu0fLNbQFMrzONttx3UEH8KL/pB6gWCSCYTxbA
w9H2inEph1zTnBGW/TiuCqdyro6mHhMu+G8wpZXnF7DQ/kwgGWfFaieb7xpJfH17eQVtNYA7dTXt
UwevaksEEE3VnEUITo5KnZBG+5U4rv5l3cXCwTLtOvEgqitfyO6QVrE2CsV42CWXRkdOZ10heurW
Z8NrgIdxiE/zY2xAKUq/0hKYChdOHJ1of6w4fYj9ZYVxhe0B+acx0tgruamLRMIjLSxm3+5Y7LcK
hXz6sc5Wu8p6vldtVGP6MuR0Hc8cr1JcKgIf0FK46S3t5cVNdIBXLuhjAU/dNxIx8dC52AzThq27
vpgnumdDWHKoL2yX9BeoSPvl85G/+pJQI20gLz8HjyW4BTJmgt5G2zWx8A1TWe94Q8d7vUTVz2wM
WKo0in2x3CkSMCjAO369SRtpP1zledfQ+MvRpGeOnQFVoGZQ2O+6Lo7o7bc3UbqmRenqzxnnvqf5
AbWoFwIMsev3dsRAyfeKV4hAwiKEoRnQ8RZHiGKzBkzMZ5wkqax00Uu0yeMuR7hhOJ/I39BF4tiw
/ukChZkSgz6wQeeW1irxc5N8lrTwDTqYVyzoweV6QoiPfhZ2st4MAEXumdRd4Ehi2hY/lP078jjU
xUOwWUti9O97EjHlac8ovmJxQOQSkT5lbhpykt2h+H4D3/1maqVRBv/bv3xf8KgG844DMFiPTmMC
taV9SWm3vsiT36jayTaUA0iP9/Q69qpIg50jjB2a7PIOvBp12Q/Awai1TtAF61v6xNpu5VDB+07t
cK1+8YDoEhx8MWuAnZ3EeHChI9pJ9h1DpbzAyWwjJFmJGdhKJy/g/1bLhvdLrhH/+Kex1h0ZERvH
GtElS9sYsU0fYzIl7GTsgSJ8Hini12ue7FN9/ap3tDLgY6cVlZ4Ah6uq/ymDaip180yFwQrfJIQ6
bCsYr7hPOAZJjdEctABGaq8/xJn1RORe1bhpmLMpVlz4raOqGH1Ndv8pIjBqPHqj5PFmO+m+GTvF
qxdhZhAsBg3GySjw0tCPbSUxNeN7jPRywP6kAgqSRAoRh+uxljEwSqk5hsP020FcUmVfjobCfmIc
Pg2uO/SyjcxwgV0Zr0Q62rtNVHdGtFBHbAE349Xd5hVGDUbTT3ecJ8tzHyWx+zUucMeqjXAJdv5e
yr5hbwTZOyrTrg6JOydqevjZA76XLrzIsA3OeVQ75azlyOSy/X3Cs5kftVgqoByYzWQKZhiZ27yN
ViVTrdmf/d9r1N+zRdLh7fTWp8yclCx24Y0thz30Bch0DCFlQV4uN+wTmjsb+O9Qh4hqmEzemSWU
9+ijLQe9nLScHP0vjfREE1WPxwuIMdukX0iEtiuJ/1CNpZPkTgNIrtr0Fpj6TnXNZQL/LX+/Wxhg
33CPc9WOc/2VvX3RSKiEh3XwOSDWa3SSyIaiLcaYVt+hpZfldHdbxP1LaY8FsepYtZRVxLpbEjn4
HOah7y4hD33APARra6j8W3fmItyMveylGOhYD6DWrJpVCfTr5GMeo2HM1c2HlXzTpz8pULMj0RxQ
+jo93Zy4NsHBqwqmqlOeyVDya5ix0tkybz3ecLgo+E+ofZ1j6biAk9B/GuRBDMzIHAR+wP1xZOU+
mBWjVvSdUblAxowYYWcUVEU6NKuXE6269VaRD/70ujWelYbozitbDtwq10ny8CI2OEDVjnW3v5eF
CI3qKoS1Obm/+J22acbbRxMSPYkM5ugYKFt/G7f0lWGRWqNSrdd5Sj/rIGtWgAVzWSIQ88ivtXmS
1Xhgui8T01nJl6uE7bcttJLkDF31rpisbmOrY3C+veI1RGkbNrpWhzDaLLYOHqQx7/PDyfgjlT+Q
TJmk706JbHK5I+EN1TUwZVjdLqQDhaXzbCcyFxsR3zN12fFHGY6XTxaXMquVO/wsuqoVQB8Tscu1
ZRwyBEBIgQ6OHcZc7br9EzEJLvTVaIeYA2Z/u4Yv4ErOJoIptIJYaWEIN/y+fYqKHh26ZQDKUiVM
eVL7NGCKu+0sZPBcXwAwXTZjDLYlloLQI2xfTLzdiLGsHhrmZt9CJ+6e+7jg9YIva0pbyvA9fL8R
dTQuHwQ948bSdy3DnKqhwkAdVuKhu73iViHS9niLZ84FRjlBmFNk40uNAKcP6zrMbH9EvAY03C4B
kAD8cnn39GmfZjzFzFNa0XEX768+t3il875B3Yl1E4vdc6M6YIV15csAIXgELwtdVWHGnTgUBcxF
xOVGZ8l4velXE6tagZhPgka44dQ2wx/wyHocuI4dkoT0PbBjd0Yii29UhcwDMubEcizPW5/XMWru
XhVWuPyKbnKCB+JOduZuU0Uv743mporC6mmc0YRqH0lqzRTogzHLW4wwoC4lMU9ITw/QEULpzwlF
zMXLSUdTg7YaVRMdMjSWAtZmE+QIMPaj4YCEdSYLpDKQC7ttXP3HEaoU3Ly932k1LWOoaSFai9Lc
LJj5J6udpKkdZ7/YJsNGctWcYQqxtccaGtYk7sljjeehF5K1GEA4fEucRGQQSCxVwLRqZOWRhPjb
5w42P9QN1zhB15/Ht4bTb8yNnP/NOsN8VdiEqFGsrJzu6iwOphZCfj3xJAy6iyGtyvXisbNAYzDp
DwosxPhY/5YaI/Fxx6aPBE47HdNRkq8ua019FetJcy0fuwq0bBqsgwW0qx38atKAP9u+146DZtKF
kh39KSFxY+LRlFcGTM5/ogxHNkrDGrEExVVLIIsATFzCCMlioOHqJC3tF+0repPfP4RNlTvyOMUQ
qdy+uTX9yt2f4FKQoLewuvIdKot1t1f52U3rtx0/RE1OI65hcgbelPtwHFGn+fgyF5tbKc4LZkVp
eqVeGWIbRXvoBgy0tmukI3Jtq92YKYXgRe8584+oGMFXYqqBXQekQSJx/TzihAhVnw0QZ7yDAfdM
8EAp8fy6p5KiyXSV/RXrmX5B5dDA+hIxvRlhc4XYXITvWo5wc5qXPf9r1A3cfrkS5L1xCQFuj166
VtWCqrWBSF5NJdAXaq5y3XisgaUnl3ZupC+9th4APPfouMn4QFmM649FVZ+1ZPLgSfCKD93xtCD2
G3StpBA1H14+dgFV3IZiCUDfh+uKMHRHmOXOMqGu0+iVsMcpX6fdDu2eL42u0EwDcrzeMGLn7baY
sX8qxl8tZneaR0/vfEAht/fsTKAJUPPm1sH81lUJm72gsI3KMoNEnDmB3yVsvMBw/7GtFYU20suD
xQ8xEMdYhoJSwOtmIMyFz12+le8o3cW8dohmsOtWFlB+4W209iuDRQz+V3oclubWFksg5nFamYBH
bbx0jwXvGnEFIlOIsvXDRtUIPOd6qk9nKIviQMCxbkqy0Fd0T60i0w6W8iZ6xNvdyTdAPdVSm9RO
CD6eefEIyNUa//0uH8ZduOuWgDWhtUlj3J4+oh5FvHD5pEa8nsQB4J0kWY0LyYfksp7UwDmCstx1
XlhNj4tPnlUKIh7BoE5oBxc5oEkFM6M5KvByEeRLg34Al53ZGUdKKGkEqLrWKq1Ug1ocU2ZdsyXh
82DNMSoXqM/imzqOFKkNuohYrWD5Q6aFIo5DGA3hn5zwL7nI3z9/f+f7QFKrSuFCndgG+uUjmFaa
SpwPJ4SvBo/uCVq0SWrKfLg2kg1uoOvbRWv01bOC18vsG/Ou4X5ti4Q6+YlVneYgma8Jn0jPOiwt
7o+8FBEKDsC0qlOgPifEsOFN8FSHXbeqm1/0MGbYp408OKTQIO5ONGMsam89f102RZePNHHp5PEv
abqUXE1/GrRw08eMQi3v8hasAuBbZMwxQmjtHKd8ZGwNwJcs8ijPKvqxu+yar9XZIiD1bqMEAOP6
4ycVQSrnKt1rSiBC2nqOuJAQsC5bGsxZuaZldC/LEzRwW0GE5hVRqSpDKGrzx/LCHgr+103cDKaJ
mCCRsqgBD/f9jy4AmdhAi0nUVHHsrrzW6qQgfbQt1NWntc/o66z8FB4SMNQBY96E81fiOBgsdi0D
FpPhMSTTbGmZXjM6nd8xtt4p9e6Ai1GPfGKB9UJMaTygzZ0G8uvWcXECZef1dr0j92f98iJ2WRVm
Kyxwz5GLnxG8UQZfLGbONQKVt30r3gZfjAzbpY139kztCxfO4LVaaa9IvHR7BG/lMENlDzySqQZZ
DMNgpgB+Ace6nb6UV6uykPzjaH9a0rStktBQCzPiyl9aoLU+woyv6ler/sC+4UWctpUUNi7ucIes
bQsKnc5k5hPGk5B0INjZpIYu6GKYCBIJ8OEvQBbDvUMq1DSV1ba3N4Ls5YlcGhENtWFODCGtlYks
XPCLamEtuXQu5ijDMxdDtSJoYRxJ+/X89t4wp+YCt4pDe1sl+GiNIoFaWCe8UuZsh6kc/jJ2vqWC
4z8Ij5gLxmv1bui1bQX3d/w7fERLI+ovwX9cDVJfnOv0ueYYiLuu6CGod3e/Xqkbe0zNScCLh8/N
VAcY62pKWJWIZCvxzMRg8yEWtaFgEpz4QTxdab4FY/DUQXqUuEpC3aHLh/gCeYhEMp+yfuzfB7QJ
Ei4ONhXywOm30G1Fl5MUZVIhiYhQw9avDdbqiq5i96dzeKRDYrCPTWEpsOT0buiBsj/+twG2QlGb
fGNYBrOwdf184CzcQazRgaOY1R6XRL36776OO013lNkHFLVE0QiEFD2S0BFnqZdhhdzxe6Qp94qs
n1riz2KaN+hvWjffDmeAk5Vzo8GCEtHnir7wK7ko2rTByoKNV9SWgs8klH2pSh72vBTVzxbNpPD6
cQ5raCuY6De4T7dael+1+GaPwLooPjJBML3FJB0ARAaqg9de8hU1yGNrb2e/a+oTJHzi9BforZqO
SU++6yP0IfSyDbyDmos6zHirbHTmPFh0UQj492lUIWL/Pt2xlqEYuXUqmbzi/MHa6E7Ihpf4ONBB
r7hzUca+2yDZG04iJApgQdmaddZNWOIquKrrZUzpaUQB7B0HbIEL4YFQoioaAXhH5WkWJnXouiz4
c7BZC2D9qIUg/3njDTSepLUEovIM85DBQFDhzH2n0icDkARm3sX4AXV4kj4MXaCmn0P+1C88Ycpo
Oe/R9N8nPjCSqDGYP+IL9mM77FTWas1urolP40qwt4OEwRGHATBT3In5I1gepbRxLYyZibwL5wRe
K6Em17IU1xKOpxj6PgzQVC/3h7rRmBl3/d/c/NOe3Pszhdag5sZ9j15xQ8CRPMZCNOKUtSrphPMl
GQ9oenXsWb6tvor5tIJ7xwmOhBpCZa6AyIDmm2Dty4lTI1mJ+iodob2YkSrDfcKdCL8BIQcNX+0u
si4HpESupQM98geBZj/XBdCtiDf37tYCsWR3M391YhxZTKGkVN3GXrMv5IzJQH04laH7cJ8/Ma9K
vgjhfJdyZam5zMdaVoVUbGcDhZvnYIzAeShPSFcJiAgcN5agdKdQ11b7W7o+owhk3hfZIQIZR9Wf
uiulSCjVXCwNv7TYl+a7BH4J9c6IXE96V13ckuSGCmHat6ffJj7cAKWpAIz/ztuecota6LM+GbcX
bx6ADybi5LpI2/0tQVf4R49W0mpHfPbQLNd4y2JPw4d2ptdVQwrzDskpRtKe7seyJAwyd6+jwsr4
J19cnDleXWikcKAZ+saPi9JMYlzhMUfBwLCUT0PwXpex8CVQci0zYIWKscl2/pnQw9O7Ur1Rz3cG
LBgGKdBGG07vv36P4wEsyuCagf00UKrk5VxS2kK4QqacWYexzh8Eq54dZlqPol6r6kOsnTOjgsHH
GoRsv5Xp5HHMnvT+uBWJwqgB4CKPl1wGbplsIeRnF77HkKvnfJbxB8WRotW3byRh6xcyiMK10241
BijOregNuZrOJCquN2e/C2iZ5pXcnZ8FUXlsLW3Yr0T7TIPfThD7KdJrQt/LXAApcgZ7MItz1cGX
HztCCj0jfiHtclmAZjLCGgAt/Top3Ib3lMc2nlHwqrSwQhBGy6fZdsQn2NfY5T/xIdy/Xdr/0AXe
aD5D0//p2oIXgJ1rKMFUcnjKhnHNSZkR8LnUnhRFkaHqDd8AzskXDy4X32DmJLUbe6UilovtMA4S
S5gQqQmWuqh6qNKHBljW1wflxzRK0D+oQKI6d+ztTsWN/oQcsL1zQKQit/78NIlxFRqtJH96Nf2t
1hz2uxdLs5J6voy/C1kLFGY3jbN3igvnOqd4dueYe0MADZVhrIsjYd53ThvdslL2cvRTT60nI0sf
I92pWq24ZLrPGy/IO/9lh7wgDwZ5QjsD5FYBxiTvlt+prz9DzHTlO7nDkrKN4YhQs64C5AsKSWS3
KIVU5EetL2qzGUd87e5IZintQ0sNk2eUdOrnBe4vbkYAZY8Fom6cGd1cvuRiH3YoI/Y1cJEpV86R
2vS4tqZdafe21HtggJw+MVN71+5MMQCCXnye0nqJL12Sww0GnbwPN87wF4O/67AhTouLrDpvFuWM
4yxqxnbMR/DDhsqBPho/K+3fyGsi74V6wHBzsOe0t0AF6UztO4sNjymhAM2dMU2fpBXjFt4DLrQo
4BlR7n9kgBrpOkqFrdCT6KLqmhKcQPS2641WEi6OHHpDvLPyk2G+CP/hhaZm4Y9HVqDqdtyoBub3
cHKshuE85rib7IaFSiy/GElTEFt+yv+Qqc//uewlKM61aQ59+JfUAahGr+lsgM+u9Vku1br+iYez
flF2Gq04iAXmb4sMmrse81GGqzEpfb9dd4C1zEaoKIA+9cp0fljMWUNvDiFnHwwqnTnxNsWqKZND
Dym/9dsMtvd4Mj3RGhjMl9R3XzLqq2h8UiuwtcvxKoHeMJMminjbtDjoVddwaMaBCJLtdknL6dNI
GrhLvlXyDZTu0DKDNe9ExgTq5rpk1+HmFxDUZRREEejbfF5TOtnBr6OfXQSGGXFGbCmiOxNA+ugo
nwKXetXoLks8Ju8c9+ZSnFz4G09e9tT+nq029810ja7TTGy0hhs8nO+mc0Ookgk5KS5O9lMe+9el
S1T1JMOMwXYkj9liZakgTp+9fLNDIXgu/epLwc85idvISDXnGpYlMyz5cwYxg7nTcnYa2a75KSao
1SWTvHsTDY07/b4Zx/IU63AMxEYlSIco2vT6gWzxq09ttJ9/6i0vJrp+/zG6heOZTGxcuKHBVHBt
O4vq6sLHtccgm3WoKuinne4LFSeOBROHKnGMT8PRqslWp2OcWhElA4ei4+aAAPCJieaftApRH/P7
Y+9FwWaWJQue2kPpsDh9sMVAZZbWEQ6/NSQL8GSMBKIbLd9fMKDqXEMhhgqBkklfvsCcP2AOg1Qf
I0D5g7PjHFbt/XWP/Nw9J6CD9WRx3wDRXDaQJWH84JhGmTQf6ozF1J2ZGKuTCUKSvSfVh4kBFWs3
L3aROKx7esYCBmXasma0oYlgUoSrkYPhoiOQUlAdXEE2TALAUy+TUMh1h8ZiErfSzdHYKmX+ixus
7EPn+/ilXamomuJPEbXQm/6Y2qsxooMQmzpLEcCiuqUT28kmXEhoUe8xwAtvg2Grdx9De8IaN20+
EkyDYEVGJcTzL0/2vObSYUWXW1Hub9ibPe4D79hqLVASSPL75V0xhBhFvI34DDZo5YhAGNl3jHqH
QPza81O5/rP0h5hUzzE7QUkCas09UDdxsKvetdjdaUsrTSr827yObIvJGBKzX/EkKamd07VSqwIs
uJ1ZbhJvxNtMeJctCMGYdysVxotuYl/VuUAybQsFo/g6eUsjMhhqdNWu7vTNknsR1mtUXQzHRRgW
O50jKztHH8jzM3M9EyWAQ7OXmgG+DI3LodRfBYhsJ1zNijKGhD7zpAZ+x4NmhgMSPt+RDVmOE6i0
rtl321OBBk6VS5HO2od8Ml7ZqtmQuuovxjX7U9mNqthKlQF1mSkEyy+smHX4T+j6WrPXCuRFu0NZ
vfNaEHYsRzfSHFjA7E1W8Nymg80XFtWdfwt13SI0o5YTjg0UU+rN3XatJwoQ5W5Z3VTMZtiGwx+x
vM5whx1mxPECy1iDQ0RvP2HFjeAr74jDpSEe9r/5MHy+s2kkVdX9WARxMFVN0N2Fi3TFV1vpI0iO
pWEXfxczkI349lHG0V4Apj6rNBsKcqWonrNRM8LbYLmuR5XrfRoY2yA3ShyM5GlSo6I1gFJir/tG
GA8fFwVJoMqE33W/VW/MX1+pLACSdJMWed+1qZCU0cLpWTqo72gaFdbi0Q1qv8vfwD3a++Kn3SwE
At9XxqzZ+XOQ4I4F/YZLRjQHD2OSW+rZ3p5aqQexS4pDjG5K0QKiwcNLBx6/s+I8jh0I32350Xja
K0cbgJoqJJYOrs0NYDW0sRYLInos+PYVvDWuhyn/JavboRtcNA4uoYFKktNNX3llLidYGsKfAdVF
c8V48QPZc5/24zgmOFwJrlIVmrL4ynSwmPBHpw9hOnWJbWXic6wiEvRo3nXg/PRYV17uRoQQ4JiD
TbfiXInX10O/GHx2VDCahi+x6qXJ6z/9FdGlEf5FEB6hw8RlKwhR25X58FCLlhziXP4lZotRDEtO
ap8zMzwrlpqUh//KVBJ0l4PiOErlllkyvJ32B/EG1jwsCoTP6ImODOWawlnE1mn0wk/aaK1U/kEQ
0MslLT3bYQiZxtE8KTE8W86PhQRa0HxyLlrkg38um43hZf52vKcNaZZSXgNzdhVIvSq7uXOanEWt
N9ZBetPgIg+FY0VETxGoWlY+mTHzC/WN2d7jpu9PAnIFDJXVv0fHhcya1qO1mHZyLTPntSnTO++7
xNKGHWfRs8l5jsRfbooJUY4NHx9J6jI2qH3qKhuOEIwWl48wrMki3oFJ331MyyV6tRsKsCyp6TD2
2IOMFDSbEleDENGyY/KLyrEndhY2V9iIIUbSGilDPFuaReM7y8lOKIoyAOwhiz0cEHNDr4U3YiBq
ZnoQ4aFNnDFh/4HKmVvIxbSfIF5mGbsl39MELZqk1lqldUrQ6nZA0J6+ZDDK1iwC51B2g9fJcb6k
R4tWTdzjXX1vcvf7WAXE5hqPoRMqk4xi3GwtwoB3pEj2dZk3gvvoEYIYqLuyTSXis1/2Q1HgtpZm
0dXt61jGafgyGJFuCOlXo0Rp5xFcHzBHGs52RBFEIWiBH+AeaHF0NCYThwcOyiYW/940y0SoE/4y
AD2Bde5YwVDlGQhFC4NphJ9laNc2msS+6Rp2KLUxzVQEFYlCLbMNCeTVIgIxp6lcvODkgz7YIrC+
22uyd7yDTFf2ToaZM0kD/18E5KXXfTuPZ3pZk+PX+sjxTBO8ElG5bdJ+aVidF+9t+o5xh01l6V5V
PzSUF2PyrB56AGBbS/32CIvF/I5x+Z/qF+J79ABLJiejX9uAV5PljDmsH8RSgGqtPRWx7f4Naz9t
3PefG3f1YI+0Hfqj604A4MFy5pLqlLXJPn7481/xnbu9N6NcFOJKDF2a/DmUX0rqfzOy5FWulVZl
hnLu3BZDbyTXLNKTg+c8pZ0ogDtZ+4LM3BxCH8lsZoFHU92W1UPJFVYYgSHqt/7T0rTv4sitSmVu
hIw14EdDlm1EKhU9HwiP3wT85ve1ntDSJoXZNGBlGtwfx+oaxjEEKadaNhlBp+tb4DDv51S4EAH6
OpcRFn3QpPuSec8ptMcytgoQDMx48HSrjyeQGJer+AiVQtUqqka9/jmD0FFIDF8+M/3I7WFaKWAe
yJ/D8xgBWXKXv1YpYyO7T4HdBO/FcsCtN9RmDpIqpz5j2yv3mqsDDK0OGQuStlvVvN9BQyzpt8Hh
/9+zSLgK6mmf2jO2KBsokP8fcOMUYG3BRzPwWybOKGFOoC4iQX5inzJY2ioE8sGs/3EUoNbmAHcU
+jduwaZLSgusJ4/3hCaH0/PZzqgVTkLlCSz292P9HYTfOLotNcQaok3i+Cogj67MsV1WaoZaZAih
Uu4dZOlsWdRIpLGjTAEClhOT2zIQeNw+oUDS8xvyY17T7Hbe1xdVAqXMebkLnwThNG9+aN48X09o
WKMM+t90n3r05FF2beb2NIGn3J4122GM3VwoxTqWPAU81/qkFzAuY2j1Ow9ERRFhWgEL5aTtV3oJ
VpBsBdzLxhQ+qmS+GNev0ZKUTwfNieSaTqcTr0riFvYh19JKj2JfwNhi9JA2qcnz4t0a0cwf9qH+
/HQCnbt6qjCwugla1cDcUOi5gUTfcoM9MlMqUrctClzoQHpFUokkR22C3jrUPH2jUkNx/3ikzXWM
EUng04jVrLe2Wd65NVMEP6feDNyNqWAIYu9gDusLcKcrsXXoyqqjPr15ANe2nQRi31C2o4emdSAQ
4yti8aQMKzW390rx7nyG1JzAu7EiIK1bhBMVxide5dX8dIeiom2z0NwWCkXGVqh1/FOv478N49XW
UV7Nv+hvC7YlTrdn5OCcJdwsphjkSclFXmO7nI/pMJiOjGWiDsrElU5h7YwC1q/eti9ti5OSzkdl
r5h1ET7DrhTHCuu30RMXTcs/qVMxJZvFjL8mVrC9qziWs7uU+TaZKrmbLR8uG3sdR1L0Hr9HcM6p
K0JS4GmDBC+DnOXTKsdCIGzl8HpJ9l1V2gP2rfs6agtf3ZOXN93+2RNvHvn2rnfRGt5ghJp6GjfT
tCwWaJxX+m5+4nfoPKGKJeAsgs+dhHHWScW7IyWvL0pJo3jplyswaunvclMBFoJn/Z2Ac8nzj57L
8pDukVKxZuPpyo11DcbMY9AeMUFExoYHsqbibZAdzZAt1jCBmVJyB5NxkaAAOS+Pn9+vx8bNilcV
yZpuXl+oEiweEC9oHVCH0dmOie4Alv/4PZm+hzCdE4sq95slIWQ7P5JsIJK/zWRds8X2NutcudX8
S+gkZm027D1JUds1DNBv5GMQrYd5PTJWD0DmEeHR5Ou6kvQnbsrdkmjMD49ShkGdo7YIs774uion
Qa4TyUhOEQtJkjh7ZHaVball3zQenjqtq6FBHZbLg+AU9osHYMO+PQR3+aDuYDrmcFsyw662wWSE
RbMBx/S1b0MFCxTgOvnem9dVEaGfka3XQbIrMzjyTghc9bQUUtjU5s8smCpGlbhNYAEtvT5sbPL6
IcDlkvOTCr0kZiUBedRJTnR+TQz96BYsZR1abayWA3vZVH+rCYG43fjll2TTDUAGiy+kWRZLTMbZ
ZO20MifvBETGC3ZlynRsP/48m4UThxpHc+MQc1mDDN5wFxVMYdmpuPMAc4gHZyVKjDXDrCbySmPR
6zCH13y7s12c0q2+xclOXs/VPPyDVe8Szr/Mt85BORkuMH6OUTCHYukwVzvksFj+RzzKFu3vrvMy
/bB8YPtLh57knoaHgqnV7TPajZ8TWCt/Fqy+0tRfnzaClbCReYlZknboNtpt5R0d5nZtZ1/5hiCz
6rmYTyvk+vQfD1l3sRTVdyx9NS35svztw5f1FDhxLOWy1aXax0Ic3IVuOpYpM8Xs/BXBFIlINMH4
0ZF1Mpam2PCq/Duwfn1Fg7Ukaf0571YpqGLz93GzJ0jjfFPo82676n1sa7aLzuW2JRgqypiFUkkj
acU9cbp1dCRTI/li8K9pjz+H9E0FKfngCaHMPjt35Ohu4aj1GeEE6f0t1JhXm7xEVBuFw1W+qLIJ
HnTitxk8QoOWXeITXfC2x/G1H3IvXuf6kH5MD7x38KSvGkQakJRoDnPToKJo9Y2eU5uy1/1+OocL
JqfKA7XL/K9okBdVlHr1FLY7cwYJbK+3nvoO/e/B6xp/6szo44yeC5V/0Im/QVEg+ENKMiB3XKta
SbJv7r6CSoVwMZyZEhs8PKm/pbUHmVgJjWg1jvCvcy+AvzNp+sGR6bzZoVcAoWjuEZu8wa9oLtlA
CYxQb6T2H8sEtjKT6pRtD/dfSpmD36/9TJZSxhOikJgworbxClJgRRd+qTWIdBh+vDmE418rApMY
vAc5+GvTlKOXcgV993tAoxwfAVJJqshEp3D1ZWDMU2wKmNCSG4NEI6saO68d26CV2yn5xlgvFBbn
sk1nvnoR9njjIbEzf0EmVc0oLgk3mxUXDsySOgKp2PDvzG/u1r+7ULFgCcYTn4feEhG9Lbc+f9xQ
aVVr7C5texRnnRAxZvMFemqhljVYLk0bYAg9a5+mEgQAD79iuLG8BjLzGtlwS61L5uq/luohhyzf
oKVjQ+++7A4N0zZm+n22KkNk2wFGc6ccBzqk0fz0tkoxsw+exbkE1DblfWwlVJMMDvt/oOmFJs/y
DozPP4gsnV0gDckDQc5YT8Nlexvj3JGL8pJMHAdLK60a99BDz4A+UZmV/+H/CbYCqQNgvWHndbtd
k57LhSraUuptcVYwsy69rs4IXrdD5RRySFcUXWEutW3FHgC5WRS45YJID9miLavuZYoqbR+0jjEC
pUklNbKETKMZEHzL9Txxe/agFyyYtRqj3Ne4V2Y3bL0CHb25p2Ws/4xnbMtGg1VZsekzcYaiAbfZ
DWqJu6+xGeuWYYRiGhhRKMH+LKGAEOKBNCalZOeHihFms3FEk2YiIYH+GSErj8izbkQsnOj0n5by
2g5BhhjlaI7J9+0X9cb+lYNK8kdTazyqaQxu6eMDu9fswx9zKBdQ3tsp52S9QGK3oHcA0mHLYn8S
dzcp7xKg5+KG1KhoUZ3tuc+zzKcZZ3WW65enSs9r0VBcsDq73Dt/o2kFG8YsMq7kLLbHHDhtYz3Y
CHqBWwGMrpTaQ934f+KsfMIBOKJzzLL4a0eSZeib456gbHrnjZDUd+9EqPKNt7Tb3Ph4W1jlZTCm
3Vdvg3cBgPlr8NPtmq/vrd9oReFodOz1X1OcIGgzpcVwemycXe2pK5P1s1Ktje0UqDAnrQARpT3p
soOcna1BG9pyRSRzyXB1ujSbltmgupDBvfYDZtSooAqQsV+arWGY/AWwfmcIGCbtFLVAo7X8rCzS
cNbWDGu7qGracalys1s1Q9FkIfH+zKNmG1rx83xemvzFUya9Qt9+Cr9m5ciaWq/R/GCUKn3zwlKZ
lnq3ZUN7yOqFPu3zXSaxqi4SUL06S4AMNQPBHpdESxUaBB3yCWJrxTyTc776jEqCh9T2kZJUiQqL
3OdeyMJm51sz3dyQTOTiNFeya9EEn4Ly2ex/kU8LwO8TFGUevtWLTPM8uvM5SgJyQpQ73JCJ53mu
J+2L9LuoNZK6eHLxTFXceAajVArMDtqAZtu2ALXEH2Mqy/NMOT4l1K+LRBflQdsdhFfzsrMqg5PV
u26WndUkiETbblvSgjRVZTBUV0V8VAImnU6vXcjk+Eb5bOvY2/+0PpfApqxvtlRvXfP5FzPVfsq1
PgCQgZkB5P1DdB4i9cC0Ale5TyhDpx/Dv7ix9plwFJJJn2fV7jnz7Cfg1xgE/dvNvhsZcsVHwK/W
DvjNGNPdSB+Bh1iCaPLbDvE/d7L7kUbfohGDezc71QNj8ZNlx07R1ncRrjVeX9hcJrv+GoZkUL2s
MbTX1nv4AYJXBEV1VLUU/RDB/xasdlzkS872cR5fsmV1nc1qXTOtsGizkpOpkaz+PJFVMIycPXbs
RS/jc/RxL/cVxSztd3GUiNg4NCx7GB/y+gLc8I+Om6qRxI5ipgKHq1o0YjqG2Hlq6b8jlYYQNhmO
9G6HLce181eYwRQR264u1Q+atpQKKolXndTg3w+wxLuDtwxlK5LDSa8xKz4BwueZSxwS/gfClftS
HtE4H6RpBDfFD0tF7qfYxYTnTTihLoQWlnzJ+4vbDYBSy6F5QctnBilopg9HhVOqinRHCyEy0EgF
GpaxweuqPcFuJpmIvSVf4eGQxDW30ze3FD3KHXjD5nfMiZtZndEWlNNi92P0potPzQfYP/iv8mgP
w9m/JnrRU93H8978rB9WNfVz4G4eFV25Yk6BvdaC5DzI6EwX1yERVMEhTFbvCz4RtN7ZUtaIZpui
Bqw0a1I1Lr1NNhUTEfGEoY7NUh8En3l/AznuiV7iCYgJbKT1Oefvv379rHiF/o15ZBIcXyXPdzqs
auGZffnKQ4o2OUiPwmuaVbgmy99x4eduQdb6zMv3teRpfkvIKsBPXm2D/O/2IBCOsE4+L/uB7Aac
76DDnxD0XMY2E0rh275GHGzTuKPvjWuK2IBdjOlVz9fnZCXC8fz/thAnRWkXegZoG0N4zIdy0d5U
PT0upynUhRdewQl2LcxFd3lY1uwALAcgIwIF0a/c8/KDzL0WK2Xe9P6jR88XTTEvXkLGUgvx+AE9
bisFo511qFbfhUu+MXh+aQ7+Vgg/ieVavedOGZcrVOxJadT2snKkRiaO8peuLDo4V7JmcKDQzmT8
t3/7elxPTQhmbaE31BUsLd6lNkhiv0lQaEJNakWuv2K9bPewdD6haA0PKKjL9XEuuXBQrOOEnc9N
dPVU807QvkSgrYj7SPlcE91WfnkpIyMoDbOSk0SgtvBvq8OiNVXu1wMRqSqP+0d4ewUkWeQUwwka
E3qMXmNhQWMacwNuETnN+eCXj4x1ogPk87FviFYIFvzPVtoYk/+aFFqFPu3srk4Mg7Xcg1NNuT2V
kZahi6oY2FqeQAm0P9ssPqW3GVDnqvlzITU7D4d0SXBfI1Ojt0omon8JMSR3fHfRvP12KNEv+oEU
5AfjADxCpm3s0GQ88jUgaYhpnY9o0VjynzDWNARpULLQtqD62keCSCCYef76owgy9MHIa5/lk2Cu
ajZoY7agsGfsg989kY01DCcsONGuqyK1kiz27OVHMemDafVarDA4MwmWnnJOfqdI2D35AEPqGtZX
woCC7WpkEycYv03F24p2Yj2Fpnw0FPaPgQMyxn+m8WgMxpibXtzXNY2bcM56aE9V30JZV+yz2Dsw
ZmZCfp9JaNLxT20wPWnx1iUuZGusB0eL+5bo+dXUkjup7B7E2JjelULDFF8TS+VBl3+pBp44cSv1
helcpAArIG71yD8dfgbeS+myAc5utozZObD5b2nZulmxuSswC8zU7n2P4woTXb+0dg5lraZPhwpM
HiDCpsaBf8uyFg/kOPOIjblRxh3Luu9Zi4jQSm5xfyP8ydjbCHXOmcf2EUfGul2y4l4hImMqZUBM
tNx9gNVJViye+UgPTsxAmhvqJGg5zcxDFYa48/F3IAgt9UoPppyJfR9WdIJb49CnZkZmBrwu8bjr
LXomi8k4CCbsrz46iEYyh4Rl8xy1ewpxq9wVBknwGh/G6uxpcsoBcXH5IPZA5OR5nifs/jH+wjTL
V/rlN0v479A9vn6W+1ikTtrSI104M49pUPxdq/yAZ5cA0Jwxo0ZF5Hze4UqkrxDJUHUlWYfuLARV
sIGvD00L1dGvt4JTlwPinxC1p2wCYJe528UU3kGH1g80rvQNY6PlgObTTM+0m5hF
`protect end_protected
