`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
DzvvE59hnIK8w5kybb8px57uro/8xzigyWIzAg6fh8AZyXgRonVzQAzAwdL53D06Zv04Z2l3NCw5
eBE6DVjnHQkIML/9QI0vgNrVJppxZ2h5hmVEduW7oC3BimunuETCCScgYy9QpibBEUYWqFdF9IwM
CgA8QxzqO++6jon2KSe+hoWxhbhozQ9q1upIaoP9xSUqDr3XVKk7t1uZzF6V1bHeFRvjKDAeMJWN
XDNDZF2z153IpO1AGTYhG/pS+N+IlIYzEKYC82F1lAtVab2zsWhTYry+HQp8QuC2LpmeTD4O0ZIu
XAmjIWPJJErRjLXxqGlSs0FG1i6Gd1wtRIiPFw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="KUdMUWC+dh8S1uCCIKcBkJkCmnrJzTbindwjDg4Ey4c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30112)
`protect data_block
TNHU6MwREGsF5VUJQFtdsrLCFGr6pWIkp2Wd2pwhDNLtQ8BNolFrPs3PG92CyJn59jqm4nvw1Sxd
EA3Q4Dj/gISiJWFSst78934mzEIo8G/PAGhmSSOUcURfre95eYX0b2SZKRL82zxK2Cc5bRNVq/Gw
RbyAEYTdNyyvTNy+bUXuTA7CnbCcku/Va3SMA7oWmschdDBoSwS9GAWBSsSXTge3zXfViZSbMhJt
nRnW+67JwSlUbNWn50T9/zoykkP4Z86MArdfshs+MB/2D9+tgJl18gIiXh2dGlD8AUb6lqMXPdqK
Zn6rz6flqqp93BHVl80wiFj7WiJmdQW38ao8i2m2SrJiDj0M3O9e5ML5EFu0ekRhYxyKp1KAzrDT
dY+2t11xr78bS4V4N3wN8zkOGn1Q6dfjRwvnOIcWywioU0CDIYfzjZcAD/9mPAHGXNPgJVNc3Mgh
lwzwTBXWO/5Fmndt4rh9HEZVmu6+sQUA3qlh52Oa9KQppKYCuOlyZ9J3T5dW4dz9n8MtR0EwBJ5x
k+6yFoOVKask2aKiecTzGa3VqwCGKaNdH1lWoiZaQ1aaWhFK8NgcAocP19lk4GKMvMUDJrIbr0ae
u1PGkDCg9NfVizEciv/iq5C3JJqNnpwmRkL7M4M10wSzCIqQE1upxGFz9k/TBcwLkMzY5hODxszE
DLSfme9C2ZXLVD/MerS7vSdlAOG0Bv44FbE/rlp426aFm/fqa2/2gc3EkVbDt/VRjWTbqqWIU8gp
LMO5lalss5zmc7Tj2YbFOSBVyGDx0oxRb9ZvGFHHtH/WK9crvsRUB0XrbgB7ugXwTB62YSuORERK
PUxPK860aFy5RYRSuGarcT7u/67rBiklOEfu1W1FjVa/kPShsqYCPkJ2SJI0Xp2HklHOJp5cxT6U
zB2i9l/1DaPwYMKY7HstPWZ+OeZ2D8Fz1fonWg04hws+xxUlqwrJfFbtUzm6LvFhxYzBpx8Ncudd
YxahehfY5keUSs9pDFi5ZRPOKe7b0qZUmgGIFq4TcLHervJQnek+uOpm5oZz/VtJNbtV6G6bF4nm
j0fvdd/gDpzlpZXEbMVj7auhNdSDvek4utSHfdxq/Wu08JwtCUfDHlyhTJwAzk/5pA0+8Bmc7m5G
SyWbONyHNV3s0dFy7V8SbSZMtPNA5EJo8iymS7DS84EygGSjci7lKkw2RFcozQRpyPoqhPalkR2z
0Yis+pAfAd8c15VZdFOK8JSiS+vCTNDoSAjgPZROveCZvOpxQZ/7NY31ZuSyBz0owYTkJ8mEzGd/
MmUTEcQsJSoZToyOaaeLh+AfOqI5QgyscdgOmOBiRE/0zGVoiH7FFWYKRJFp2LuT4rdSsBJo9khK
3+qT4rht3Ooohu3YwsOpQZdN9TtYZlIXSPJFEPithHlG8L/jGOOZZ1g0nGRjnirdtezTUswuRywo
JkZjv0Cn3JTsw2Dzlae8ejxgQlE38UCA948WAL0V7PGG+kCmxnzC9PbU8hi8Qh2OnvQohDHxeT/Z
8Rd/w2dJ0LhsD6PGdjAQavwgrmRh0WHUr3kuB9z2zl+D3narabcbceIulP1RPx3vvmCXWsXlwfuD
QBbNmSRbC8cMM0xPbvczCLc28IW14Vg7DYWtxxzLOGYQcg0yRahlIF1Nz71dxtZdvi5f0U0eAoFI
iA9k/7oO7GiGoPrJBg6Bgt7etjd+v66DjHsuwJ6mth0RVOw/vwk4BRTVyANQVKx1brj77BdT0jPw
OjLRiTycy3Z+j89m8OUj4CajszNeQtAT4B1DfTNN5J40vbp+IEUT/sPTgU/NdlZjZ3ENkB7fmfAa
YCJvG7F4MWmSaD4Ka8JTbP53ODV+k1ADcnMTNAjfqUaotpcESuCUy0Lip4B9yScEk2LAcRBn0er4
sGroQcdg78vsaSD37cpSsSsKdtTUte0rDMcRGYB/97HCHHWC9rooYZvYYHfgbkqDvVfXWmP2FjeZ
7XEpp3ZEFyO7Zy2J58oXMc/8ZPqvFtp2glOYHTfORdD26OeZ/LQHG9oyju3bRMI3L5T9bTjEDVdX
c9wUumVJN5xNEn4rvo/wHf1TgDDi1nNMggU0/eINxb9Uy1pouybbfqILfwGLGH2GfDe/g1NVfdHL
N4N7SZ7ECfZNlAr1PwOtAlmeLycb6nFVEQIpKGJR6Ya1qfh2yE6WK8CAu/3+ugXqqTn+xeYkqYkD
pDX3D8zWNfgStzNvMBNCWdXgjquDjH5SmIdCwVSJJM921Eo10k9/2nN+KiqJMUCyUSrkI8OMgcaM
yg3bVx3HiEFpTJWky+QZHDx2OGLYJdzzOwpeFO47YQJ6B9b+R2HA5dLNeObkHxUgwP7YpWRKNYFN
bQuAfCLGxddIvB7S6v5xafR3ZPPNpGIP9QGWC5TVOUUwFW8PjGOZYpvzDn+SmrOPAjadDD1QaYV1
1U44IYPCzIrXx89sEOvoKRTsoVyCkUKjFrJX1uylNyXVMtFT5hPRHuOaKxwho4KwhD5/mTVZ07PQ
gUXt9Fx0Dm4etTmwRosO8/BatjSvz5Jo6zaNLvDTlaG3hj/WYbjrAnd5tmdnP9BIgPWYOw2l4Off
aoePjssN2skuKkJ6HM1cBiSlnXjWOi7d7pupz2cywJTj/q0iiSOVSUxncSRz0An3AsmKqdMDsjNX
56jGirSjQQDl6gSwAMruWu54UuF7btVxMXRSGLh8yZcXLbp5uv3zekRPK9/ZLrVxXPGR9a+kG4rc
Aw16louObNmeUGqhncnoLv/+mNHvjtgKgnMQNIx7Q1+aV1JjuHwsR8EGfNHoo1BrvbI87AHIt5it
V69Ne1X0DxKqEDHqdkeg7gVfXtTYvZvpHoIx938INawPS9n8RuQjMWzcOBA6sR7QAlAlz+bGqLEr
0DtVjI0db7Qse6DyN7z+KrU9F1WOZ8NpJ49p5hacBpV3kihfrDPl64gliCvKEOJGZMZEk2Hfk3ty
Fue3x1jOIqXTI2vYpZ5Or2zipLAHIBRbvqz+6S2bHNsmX7Qhedt5lDgIy/2iB5+YJp1hbtRWnpvK
GrDQBldRDm60naD1aWcCdsF+A0apb+ekjAcelOLzRi6Im51Y+QmGMRnHoPyG8tIPUjtLkkwB23Lu
LkFFoJMcXrwOjBKxR73THek1K/D+iGaqjs1P2d+bnPW3fa8UeFdMDuhU6MFVu9v3Mig376Pe8BBc
GnOkpf0HZc+N8vLkbummgn3wsgQPSIpm7Ru9UFSow39Al01zafRiF/VOP/KhfTKDmZvpyLCGcSaa
/JgnckZgb6DLn977VNveBt5XDErDEdcucThLqlig6xTuZcG4xUq1OKU/lgdlJZVabcbE4CsKPfKV
fJxUMNDiPnki8UN4El3pxjb7LbF9RN/GnRrQCHuDDnaE8PGCA6ldXLMSRChp7cQNWy4Qaqo4UksR
TR7F0ceGBjrEKNXb7FybIej1X8Hk8Cvv+OofLhrntANtyMds+ap/ft8nHGRPos7pllYayLqVe6F5
9Nf+yj4LnnziiKQgcIbkiEXV0yeiBW0jq1E3Hl31OQysQaHGZYc42nS011oKCzsL1GzzSdirbc8Z
wpHPj4LK3Q5mSN/CXXFeY8s9n1J72NZMSoZA42li3Yeg5EvYI6u54g9iHbB0CJXSlzZ/kOoTFOyM
CVnyJBRlTG68QXt4SlT1HCH0gPTRZPG61YBKdyGHC8HgP2U1cfvRu4C4bVSGZcmFkukKwStuyZvc
7Bu0JKI9GstN+vDW0+Sz/oCwgIh7drrzvu6JZZvvuqBBe3b3iQQPMfGB0Sm6XI4wx6tQe1g175Ot
axLj4cdTLHHToHZzwpFIB5l8ipP5Wx2HYsFAIdVRT3tp7Ed7Q12OpEUZKl1h1ZNxNTLFBX05OMgg
S7mD8p2dQxLsue6EDBkBvG2+WS0eGmuqclAYPwApwiATIcm4i0CZlaJDctR8lqCm9Y1C1KKbH/Ym
PoB4VHTMSug58YGeIyB/HxmMWf1IiKUuO5s+OgKrp/W0jq18R4wFkChEN5cXBq7Jch3Z1tBCYnwG
Hcxow2UcG4HDQxGcwK1ca6ivRklIb7uhELGWmCWa8yLFTRWDuOsgHSFcDHEThR6S7KTonTP+NEvR
S+Bis9+ZRY6pabNeL2QhgrIbXIS4JfPKt0BER7Isbonm/peTA65vmrvl3AhTXrfTmcfu2m4nl+ck
BMHYkOcudQH+iIvRmZ4R+EHlyaUO+ApE0rjRQdIViupYB1MdVsFGf0lpFNCTFoc8DFmSypZc45Vc
VATtdeMIRLzx4Ra8JX7bxkagDWyPb1hyYGIaXUomwM7XTUUF9H92Mh+66hHjXVazxaUCQYvffUwN
8IbajEF9clLScBlRFGqfDYdos0QbWr9kiY4Zl+AdpjYnhwD2ASkIqKlahRCwKOybah9Q4wd9AZlC
dDxTTrWalV3R+fghlwrou4MBmMNz89uGK6SoTcgLF06kXmcLj5lK+W8AVHStGIxWEuibuydFyCar
sou6Q480pAYIlsOAWMRuv5eR9iDhu3nmMxK5eMUzOP74MaYG21CXcS78kfSqeMSR8Desq3ISA8+y
9lNusNKGv5M86Socvx98mpwC6hqmp6HiCQSZ/bmlJXZVHX2phTS8am5YhgdTZLwWgvhyOvlRRq4Z
AXegxLmcNnDgpnwoMLI7w1TXie2hdvf/hXON4rpEfdKSssbOVYDWTqQKvEJYMkB6wHwlYyERplDi
7UTyfTFNdxfKFfPRstVbDLNS2WJR9cDC6C5BZ1kFgIlY9QgjsTdMU5s879eKYtJjw1uEFNeFuJnI
0NfVg0XmXPXJtUOxn14mTdUQqqIWQlpb+I/T3EB3noDK70Hg5lohX7sczZOlZtykzVW3liSDvKNY
se4s21meSM77XieHWQSP5lhoJ4xgLakG7273eQBp8CqCxlJiGhhtzpBP7j+GPkyGhzMnhgzIoEcl
NBRd2pDhEyeLMBMICa0egZ3nNggLVRfo8qhazXjdR5A//e7dGkhURH0fD8Tdmr5nwF/oIaafppnh
76s2r0wms4IVrQu4VI8BXWyDN8gn9ql/SocsYm7CFp9G8mTQLs16rvvuXchTvpU+eboFNinZb/4B
SPtd6D4hCZepZtXXNw1QRxHvhUEh8/Pt0livZAOtydMFO3O2OFlw5pOvZzLvnjI+s24DU5aw0rRu
s8+jc3SwCocdv54nMzviTngoY5NKhYUfvJ+TRW20ysklfdwN8YEr4QnGB7OKViZ184pqXJm7iR7/
vSrL4vSB4khIHySueNekBMi7P4tvldJPXkotDqL/GXS4E/aS72nXoyw3rss0gp38kJQg1nygqhBb
kJ4hc/LGdSZ6YvY/lFE3TJ5ofFdJH5BP0HCGj2PIp3neY9V/9Odk/XiKuzs+D7kpIeZU0qcooSCn
+4FAPKriQq2FDMG/69tRV56CmNNfkUy8wsl3VVOci42hU2j5YirvcH31Y569HK7rdMil1TwwUBy9
3j+03h68dzOPkg0j/S0ohYV+MwYfxp9NKYaShuaLEgrWfVYCQ8KvkeHUP+NTwEtWxp8uc1XvYLgj
V29NO1WMhEH8xJQ2884LFT83qVz/HOM1ziv8wGw3IcXn/NeeY6T2RD09eGD0zOxDm5JqQfnWdgrZ
4x8j3GPf1+O2LOn4+tPxqjW8BgkDa8EuBgv/fcGLfn5zVoOqJ8ow1lVDkCZRluhl+sN3mZn6q5zo
Z6QEiQe8kEpmyQSVYHDqPygSZBE84M3lwb/+NhtUuseHQ4W2maMwVWk0OW2csH5jzyrCRxc/TBMQ
pZfqF5lU4Ps7Aas2FGizTjpaWlCPzBBlk8hiMmLJmzp3RQmTSso9maza/WewUNUG4waH955Cgj91
lxIImO+5J4Ha0lxw4c6VFEsBx0wCTOSb5wL6luYSyZSjNSdNVdEay+Hs2P5ELZJguJYB68xhvyg+
RVUEw6Pp9r/lx7HW5ah5JF8vlwiVAnkzYqe+JKZ2b/sDx52p9W7yG7z3xfkYhB7x9hd30SZqq6eF
aDvGZyx/s0RC94I3xMpACinOtAnwVLaVjmW9XKGavSZ7qkDsTzyCmDhkAAmmUqpijG8MW/ZDdYn2
VTz2yXo/0Zecx1FWtqn4Mo0djFKFY5eBPnW9mQddJngWJRL92BprM3vKR4xYmXa+HtIWMd4w6Qse
zkFpc4FU2htkoaQoiIed54T/1iIOOiGKGP6K3EWNKxV5NKapNgwDKos7I7TKLUwN/NBRmQnSJy71
gHI+arvrHu+ZhJS98mI+UAKcV23boWwGaiY3Bj80LWdEWOBdO7SsxuOxOuCw7IuBpfsgzeWRgz5L
0nNf3u1XuQNP3KXyyYX8+qps07hrVJTmJT9DoOJdfVZK83BrKc/+I51MOJHoqAPVwwjxmLPmhaAS
5Ng0dMigXi/iZGjf7Yk2MrKQLWCZq7PcseQogaT6IVbXkb4TcZ8orrRfMjpuRXQZDzb3kNK72TmI
/7kOmsdL7cmKSZ/mgGjPz+HAkv1qIHT7KHCBZ5OMiFTWxjOGILnOSGmgZch5+i9s4RONRJ/SzWBH
4LAfmRoFZkWO0PU9nBZE01A5jhFnKv4sza0mag3jT6ix4Nf6YRbsi17FDPJPlrKzcpBq5W6VslFb
CQGXlcxNDAzohY9IPkfv+owiIaBuF00I9wAeUSA12MmIYpKxGjQKkOUgj579rNpZBEaWkhl9MJNv
xlS43TkUnYoLoyLDql+b9+l+BFwT6OuMXE3sizVQdSln3b4H6MW2khiOcDevDvAH6sBxGguZysWx
yfv1J3G7M5seaqgFjVjWcSC/GoNFCPSG9LUWE0Vwn4xpySuIswJJn56wb+2Vku9KbOtOVNyawxqY
IFn+BRIVHpPd8i/1onZrJqUUBfDYgoBhuLI9xzJ467Q7aj4STS2Lo20tpfXjD2+X33ahm9FXy5Ra
AN/gH+Keb9yBIL6caY80xCn2E9c5nBiTAeI6Cnjf5/luXel8wnbpCWB6pRsppvYqV9TZVfNji4ek
sS17GhsUGkdjGGo/ZaRvLj9LkWQ5L0+nNW029x4vVcPy8O48DkOfF7GLwc2M8pNHSzYquI+8dZRv
yqOZ2pcd8hDX174LCzWJdmhQLP31qOXITMmuhDVc70bQaqXOmZHY8cfwXvGybGyGXRMQUqB7Zb1u
xH9H9TSIjeCoYrQoROTddtxD76DCvv6yXs+bkl0/sRs8zEmnugHH0cbdHxUJmGrqOQTX6pQttGcF
CILadY14Qqh8xXV4ecTJB/9OMNRNaoZWcvxXtuL/PlRtCYZgO0bbsQkUW7/ZdhYEfchnS1smO4LV
RmB3WVjUMoujeTha+EPn+qqcRsz3ZHY7yfUuZ4A7D9UdadVuHd+LkE9PNmd82YXbrFnLe3YVaCkI
EmEFPMKMHiVduHSj7DaSQG0wSNmnBoTUv5VqJLraciIcNZ8hiyhjLkGzpDMq6SzNt1Mw6hb5C7CY
t2aiaeN0X7raEdmn88JDkZSc1wv2J0Nlm3MkckEcK/EOMY/H8MXHnWF+Nf75iOghVnGSI/PJ5n+k
YHlF+0QEcmDLbk5aricmGF3n1/BrYqHA+xwZEacnliQoBJk1aTzbzpzDRSW4hsRXFgvuQzrnTINY
OfuQDTq8uHUD0oBSjXc6qDWFU6a0Sq5IiQtsNIBJ6IiS+hFk4l1Qm0bnmf1Rgpual1BAI7UOJBaX
fjqPkuBYesgI6n2mGhriBnvNmke40sTl6DhBXofI11rotzXVy2eJhqsmjsgAeySn34akDC4QmT2N
b4QjyGbzzushC/kc6Xz4wuj/JIs1+C3uX2F9ktV28lI2aT7y7lbspkFvGOosuK999xaXlLJod+Iw
ICdM9KLvd8lvQceUuE2kZAiBmkcXFq3CHkrSgq2CVJS3Sf2TW75Lk2rhuvbc9p6kK023JVANS4/+
RzVv3w1SuPauzPoCPfozQk/QXdxojgStEAs6qLZ4czPS0DUd73eAyUpQnNnp8B7WQEaNI7S+6vlT
VrzlNlSPYjKm7VQggYDsffy5UGkCyQaEoa+/blXQLp3P2UWSxlwQNyLe9pYzJTXfxJCpOHkMG+uc
L/imrAMVOF+Z+ihmBHKW5uxHZg4QZ1bQUChhz1G5oZiRk2J1ITs/SAahmqbkgo0Ir12wrAv83AV6
IDlNqHw+DFZ66V8Oqo43kCWn7FMtddcjA5O8XuQ9Pi6x83h/nQUKZHv32SJjUEcX8B7BvOKhhuA4
NOutoKmRX1uIH8upcXMQ+398JUjPHHNOaJ93ltodIBrtJe9OBtFv64jnosb9feXE3FlHFAa9jwVx
n2tjSZ44Dnzq6Ye/+2lBjcjF+yEVHMQPAZLDeKhF7togdHFaBtF0FTEcClW2Hb3WtWpwXG6Y6je5
/LSVOQLL2hOB6Dw3FVonI22LUs0BrtUPOFpOx8UJ7OP5GrxEZvJ2nTfrIvmZqJyehrNkOKfG8eiJ
urm076GyLw0Aqa4W0csooaAvkpbBmG4s0WXewva841uSj49w4JDcxoO1gIECp+lE4g52TkmcXllC
wHfnQDfdaOYXieW5v5LgbnWxr3ZlVBrwdhXI2iDOVJ4fH30Z8/FqnZT2sbW7op5te8y8VoZW9ujW
QlzTsh3KvU8Ul1HXj6qXJRlsPphvsVgZAxMquzigVylylE0Lj9Ono8IyX4wR4B1rkyntxEp4IYty
uQ9SdKk/fDomhccowu8Ynjkrxv3EB5Dg7D3Xb8nxci8JlJDk7xYLreYFzohuJRsfu6gYPKohR8Ph
5LW5+pqxFq9LUcUpPYzjh1/vvK4JJOXLeStrO3YZDU4oUipvGuj0YSUCVo6psbaPi06DIruu96eG
0pXdamk/o8QAo9q1e6qknrUvJrBoBcXSU4IvX2Irq//YFEB/ogi2IeapUQqYDNvKm7IjV4RYE05+
6imQku9OWqZiFCjUOdSHsTMrUGFa3kYlAo5p2npGZlW8eAQSCRXmU89nwu0lJLdEg71mrmU0/VPJ
gRgFhaR5K/hicTCrYxixcxK9ObqWmXJkvj1ohSiJEVZp4CUEGecAkg3E+LciYQTv3RGHp2GnXYLd
IGiHmQGkS7+UuljDOOXf4repl3uGBm8oJCM/rPaXS9PONV9cF8t04Tvb4o5WXU98E2VQ462eQF1W
EtTKLEr9S8tC3suLJUwTBpwSzFS9ZquPbj7xv6hJTkkHEi7omqf/e3KywKVgvgU0eFJN5odNxh0s
vMp21Q7l6aowfRaYeo0n7xbOLY7Z4ox1vD0RR8Uz4RBGHXhM4NuP/A5dVqg9iWvWCDLlKdf46YwT
FT7Pwdo5MRJwa9xk0aBrhh0ezkDEqnP+lmGFEp5rNOD+1xrif1Vgukkl6w7TYkIFd+Dm+sxWrvvF
VKGcTrRoqFg8Nb680iWHSzCpts7dndKfjbHop8Z1xwnsDBuIpGHBdT7tEkqwzZ2WSMY1dMEtPF7o
xWmayvQBF6m91slegXgHwiearxoEauZzkAUM7QBh0urHPPIrWDt4JiPLE3yDGW2VR1Y6cAwWDKXs
LYGj88m3MI4DYZeQYouHNRLO7mqmH+cIvvG0Ky+lUk5vYzmfUCQiYikzNFjHP/HTwjNGhMCaQP1L
meP/tCGfKYKnY7xlPJThfOdwOUvkTaK/+sF6daydPKwy92Ig2H2prU2i8KBeumy2dibKufd36hUQ
WHOxXaBNY3ToaAuapsNiygMsUt3oJbeoSeBBe3S7R2u2kOmCTdbXSdfK1IFyvXNJr2WKaplBU6rr
7TnOSCuTg8LwMCJnEv4YvofK5p/4VbzYMdQjjqFWSxoCP+TVKC/qUTgsb1d0RPELiChGFSQFkuOt
nlDVBEnBGA42mhkXuhDqKdUQAA+pZcw139NC2kaShZBT4RCeknfNar04i7HnFLZLYc9PeksAOLPG
foYXgYOnBUCG+JKVmywJKjsA1jnDFyLekHAVIxQlhwsVVe4FmTHNKMLNUCOprjO0DHCHbv7mAo4x
xC+QjPQea/rM/gwwRYLyjfVMirAHVBsInmulCXteHYT3QUX/uYIMaumShzk9n0yWjHLH7t2vwasP
3R0k6dV+aFVX4ODIwzHtHi/iFivmgyE+8SXwyffiSzYlfr7PYl9cLkfsCZPenmcb1nO9MxfJcuy0
a126lEx1MLPIH//G/Zr4GAC3z6SvJY91ZGyGEq5LayVV832mp6ups4WefLdkK3CcQhqSAtZQP8F+
eE08Udq0T+z1ZEqilay3Mn8HZ0Kb0zYHj1QrEp20YU162rGBVuSiQzZXBd6N7D3eXZc45a2qlGhP
dF1kb86vwUm7MuDfrqCrAGiHGRJIEXIk/Ttj0SGopUPKWBIG3WhdCwr8X3DAqZ7gwU1t1plqUFTI
csuZkQNrjqjMZJFv0Rd5/sAtSHd1OBOh8jAPcLVzi+PKDAsOP2C6klF+zgFWPcQfWdeFxOc374Z2
pfEz/WSFLpq0nRUUYjw6PrHvhUmYfW4kc3j3uJKuo79cUuCDEplTWh5tb1/HbR0XWYPnCWVI0mD9
vuMY7RDrjU6/pteTRckyb9YxdVSNWTZgras2LVsUF5MKzM6E4BWm3abVOsZKBgkbkmtll3EFt2d+
LWCdGKVmkSVtQW4B5cXKQbbXZOIuQCxHxfsGqoe/fA6LqdWaZRH2rL+z6m73nEPsNkYhiD83uQVQ
6gYARWeW3r6mvDxaIwuWorqF3Aax2sF9jlLFjizKkXsZEfMxM99tRky94HfVw+CGuGPQf0f8wx0W
6IMQde+IiGNcNkRB2SI0aHW72lOGM2G5I03V2iwmEAkIedLDSISRVBQP1PuEw1bVBRSV4N/5vqda
leNuV8F12WWdWrBDQJNfzxEqcfaTEctwudrUf8gBHzvJbdekUBayC2i1eko4Z3AUTMkO3+onv7nb
Opt1NaitdIOL00ivsKv42fu5HFc8nT1ezGk2ymxuizjIhqmURAzzb4gnWqjEXk+pOoYNfkOUrjVW
diHHla7XxfGFarwtwcfXuo+PheOGYrYUCPq5QZR/oRoEdgwoilNzNXRMWNNRgxmH/0MJSHfxlX8N
qcem4np8iRFPciI0AChIaK9mH4Cz0cW16q05omlYwKjiP3Px39uPsTYR/2xLCLTCxpZnQD0u0Voc
CD025NRKZkS/yCxF1KIK65YM0SKSYEcOLOTmF/eITsnO/zFITbq2EUs1MWo8N+qQvMiP7up/cpgB
cqUZhBSCoZx/nRAJOYtf/mn1RiHzY4ZSiK9RRauPMjrRIbp8P4egyCkkh2v59j0fxDUE3bYWBTQ1
7ehisxuryxVSLgDWBy5B+kCb0wHp4mpBxd6a1AjkDuUoLS53I2fKerBvEEJ90ehnSbC5PRv9rRl5
SYvi+xrmgIEEFz3LXkEmvO4OkrM1YwR9MsOHCd4nbJoZixUy+TxRyA5SIXZP6Fsr/3fUTjofmCiy
BeOP7C+i7kcxrBaijCmfpaF9RPeQwEAMjcpDNeFqVJRXukJL+ptGnIEkaFd/VQvU5FjfqNRsKNIs
/j3OTDIXW71PbuLHiXiGtrY+545tEnGrZcEieuanC54uumqBFHgNajoN3cAlmQRC68XeXXulXzx0
g1S06VKu3gTmB61TPgpIymlAy+YwgrsVjgM2q8Q2RJOKVDek+VyUhVRqpx+MMD7eOmjqrdMG3MrW
mlCXNDHCKFQNVoqOAZEfYEVE+i/wAZAUf5Lt2A1x9yH19jWKoAbM9UVm7EGCAYoZeZjwrkCsr+bf
YNdXfNZHAfSv//Cpq0RSGKEK9zx2JFIDbxtUBhrjO+zb2ZB0SdjMlanCLPlolcJ4OJkvBWwjG5JF
UM99z0PSB9LsDErVUV3t61QmKxRm7lVwzJFqs8jYySWbkbhaL2lpdGyhUFrSt/1Y6MjKyxrD+bbu
TppoipYu8GLGTxOLQkkC3CfPlo3qNE25yCBRFRvCsE0K7PeTj3DggoTvoJ9zBzl3yeDp8mFm/IC1
NZaoi9tZrbXKVmlRxwuONaxuJcCWoAtK5I4DVzcYkCUMOxj1B+pQqj8/XsgW2EJFwUdml5Rbd/Yj
nyenaQ6f9s3zaV934i7irvKkG3bw0yH11DyXuwPhIqzYE15JgVN8/8k8hogNLGfovns8Q3QW7Qcw
4NOcgjLyCzf/TCEU3MTv3ufSUE0rsbh0ereDEIufDMOQQlXFatMHvTIBuaR9nD4E//FTbals+Uzw
Q5QFti/y2ZqVEE0zg7yDDyWvnBAhp1KTI9JQuGwr7u7nRjX1L/yP3IXqaOGg6Sl14ZBeK/cZfvTe
zU7crY3EMuUxequnzMQvq+iqrWJGESzbOMZ6KNktN3c5hfLOwiD9JdEzo3ZOx/kOZNvYwwl84Uut
tgm8hhypvwuSL1SJqF7/54DoMmlCWCaUe/ecjUn1Y8W1lOQ4gozmbsKMF0fN6pTZzr7QGgPAYwhg
HLWpQQ9o6xN9pK+z/94d0X6jbmdj5luJmnrytUNAF28Z3H5he+XvrrMiBWiUmlVfZzj0U8BUV5sR
T+1+dPFetHB2JSQeS8F96GZcSW4gv/wTtmB8nl7ID2LUPDwK5nWnH9XuWh+H1a3atxpGFs17tIwt
9EpsKSCEj8EPiC8oYdmpPHUR/GKVAX1tyBWOiin8dZpn2Uxlfo2D6mVozmj4ZlI7aFzTSsLPpMT2
bxu8rUu2PJDDfDqNei19wby03tcLyAPfK/gqQwWYCifdQsDjHnb1rJsnGhqSxjshrnnqw0LBdMQU
8hLZhMh2O5xnYuXnI/fSO+4mPJ3TKzilPfMr3NFLLv1I/DVYpvV2fkFCxa2uZtTV76DGe9qUEXW7
t9G6L8Um01u4FwlGdP1fTbtrYnkQ0DiXEgmMNkkUOJ6RAIwN780DkjLJcfTKeahZZ6dABnJRXn3m
pTNyWQw+SnUWU8B6auung2Yi8TyECacUFKjy9gRBYIJO+n8k2oRcKDon41V0W2PdobUE3xELaZsl
5YTWPSmc9oWmIQJb76R5lX9GreWyLr+tfmRuyWs5HnKDTYqnq+dzCnUiZf+AqG0jSG2KtFCItkNX
sYrjPfC0/pmRyCPMdFeTswfxGWwQWplfgrVqX0f4Hi3ej+INIHC4GkHmWV+w2QkMjHcMIVIEtd96
/oQ7jfpsa5X5t6yKTe85N5hK0zA/rs22UCTtuc1cu/9cyF4rnoRBxYq4cXaKJgaJ4nDkCED9z3Yr
wOsoDLBK5nvCWoz5D++W2eNGV0kmV8NumNrqRHv0G8NaX/AY9qfCkxFnY1QgEeeujt77Nsdh4xn1
U3WW78hNpT0DFQ75LF/mMFUsyfuwV6vT7GGGkm6QVa9QhikfC8Rz3vC98oOQIH+8/N15vntkstlW
2iTQzUVkxs3XDzUD2btPFi6IXQJY/P6YrBJ9HGOH2N5B40Sq6WNUHMcL+fY3ikXFDrFRvw5SZJAo
yvfzz2fqZvhSuEqEEFbnsgErlwMwo5Hl1P8bOSooNU3g667bLfBiVMRYnVsnfu9RmZLDmesfdxwI
YQ4AB2x2hbxfLQaRgmqK0cqjnlbgJxVdVoOveIpfdvHVCiF4THsTlwM/40MURYovzEV8em1CyiLx
UbEbrScQtsgmLy0VE2QHQb4c2jJLLyZKMGdWfgOdSTCW412QfSr8P8Y0LtWvDzv2mfWqd0Gr/6oG
fkkiO2BWYC7NcrXl182WJxuaUgA/1ufMx8I04NpyymPxKB0sgMs61tYA3Fi6F37lY0ndyZzC3GyL
9JAeQ/N4NRT5CGrVdxl17F0PtICV8I1IVs/9VAlvqPLw54w565ip3xKvvwCV7N7NnngO8fJFT3R+
7FdRJSQ8dzfnA9XXkIqBttZl2d/KXrlm2/7iXKMUaGBn7rdFCVG7pdYVeBamDKLAWTfNhb+NTXaT
YpXuJlip5uQKYj37fY6DSRuTBKz8EzbOxx5fvp8557a30G85EKqircdF6xGTxrk+dd/J069PJElA
gnRJaEAd0S9RWBP/5bPOouE1Ay62nQOS+8k3hzJrgyvxPpvvvLhyeScApZSlMxK71vWKXmrTAg7T
sDJ7fYohNW6jK8IdRaSQdn7YjFLfmbofA7y3uOSjbD9guce5FpELnKdBEGx7mGYRVM/5RuRAKn76
2gFOt4chyICQD1kB8C6e///l7ey12cGjMAagFOkJtzxduHhRY/2Td0+uAGifAMXcc58P298cSYu8
+92kcQbETh4aTW3+vdsoOZ3gxb5aBoYH3jg5AiANrMsfq5tkvOnmcNpgk5HRrp54IWNb6IGxyEk6
h5JKKeWmcdwQHJkZI46VYKHNYwL+Ec2AvHX31vgyKs9qIUWCtFKmmNqAufw7meYCPH8HdHsOEwVe
PoWdd/MxfSeBAb/hpTTLvaIwACNaV82qxSGrAnoHPtc7G3BYJNBL7eFF+Ml6cI6uo1AmFmLESqkW
EY5JN1oRxiLdlDaELrU4x4KKjSXgHxYpbd8VJlrg1oZhzo84MOgwjJIqLh3C8F358NlnIjT43Iok
VBcnPURaLCtD3ZnOrj1BNT3kqdqbjbTcN+fIk/S9vPn29A1AO7JqAv5KtmwhAg7L0LLkYXLnp29C
F5S1jjjTa5z+IhOxnD6GXiRoF4M29EvuEE8sJ2lQzSwHZEc/wvjfq3R6QgRgR+rY8wc99CYnb0ps
UmF0IwhsiEFuWSr7vHQ1ikkykknSy7KZqrLYS3HPMK0R0lAyNluEMXw3g+KDwsg4E3/M/Dp8JRgA
rsJb1iABNjxrkyfl9M8EjqKC+bUmUdftJWJjk3dPHmM/hNCVH07SRvByXGoL5B4ZbL9COBZYbMoV
NKZzsaP4NqfGXujHjbTGOBStj1etDvAOi+j7SFuOaG3fsNIrQ5UNhNFGBohyzrlEQNjyf8FAU8/e
V3JPk3oyDtTVQiZPm8RXnLejmyVC874bJcgosCc41GqZIZQePXQEDVZRjgQXNQwMfcQD3mKcp2xE
cnydhzJ/qfzvkAUUKCqxpNQUWHP+KIQB45MPZ61JSPMmvs7UPJlo1gEXo6JwjIO+oFHBCZTsQ/aI
QIlx0eFbjIbYvUn6+sVxVAoIdlbQKz42dWXtlsLMiJvNwfgzBA8iP/OsYOmZLVlKgJWe962N2Hf3
dWiNMGB7rqLKHSzwn8iyPydQm51VQHb457dfeBlQWLNt5SgaIyR8Ci3UrN/Sdj4uEoXGkPxnUwDH
CrmsqfiR0LwWZstVRJlJJNNFkbIp6xF6meQ2q9KY5cF/wJEz7sii2WuCAtp/Ml/5M1/rwh0AR+Vw
j/m5uCN52gYmLo6JZS8TePjDg9IIc7gvZ3tYRS5JsJYHBrgOyK3ye9SKe2Qn/kOjs7czNMH3xTvb
ccmW6tHqtaTMCQwW08/GmWRNU6CARj/BXRCn60TO7ijGyyM4s6c3V5ze1TL8ZulyZGXv78m/WuaI
gF1vWMlzxQzlC1kF1DrgT2T3KWrWOXXFt/YF8UrbsXbZuCIdmZbQtQlS+7toureTCWs4HiAQOSww
JYVVVf7TfnRFIFloXKBJxp04SoHNy4e4Xt3QDpIHPaf45+ER7UMwsFJoMIjCNRzMivYMcR/xcrx/
fRZyzOsiiZ/tSMxt83EpBCJ0LCScSnejGPpJAxmBtpYXFpBm+CrvdltusfdeYQWnDkWSwgh173+7
gbd0wYuDwTovVI36uvwyLxAyJ9ApAnuwsNisENaqmefJZ/ivY++8jPFCbYx0IZruXfCvgGDwyYyM
ePuFFggeJRP08Ntwat0kYBHWtKjH9D6b9JiYBiC2CyLBTa2dCwYvYnuPnkqTsztg/2eL7KTY7b9X
ZmBauRpHcKmH6ckt+Yps6SXvLLtnJg5XoR/beCamoZ3jta8HHqbiN4f9ZWBpDn6FGTivhxYMdjsr
+gyiLavILV0AYvdkUtFcbVXKrIu+EPzX9whGMRE4dx++e24Psg0KXs1DeL7Lh3ExI6KH3Rp+De4V
JaJm/4gB8VvVAVImZldAVpeLEMkVosbk6YoobMxaPd8oS4a1uggTIk1c5RbI+tzwppvQlhMUAlzg
QU0yOHhsSLiC5TveXXn1/Wy9JbgeiW2Diimu7ufdhuh6pzz2WyiB7PUBTzP+3Uv8Y1aJ7NTw7f4B
gH7ybVOv00gNa8IdSD3xlOnQ2pNRKokzBpxUhzm7GzF0EzLa6I4NnkVhcRqVUXx8MeAbkjhQm829
7SAINRj5OEyqpB42y4W9cogt/mb+EKaq6UpP6S6pjYWydUKNuj4Hfojwcf4cu9DMA1H/B09ruO9H
yI8As7wpkoiX2oEvxnlnBgrC7p3ygJKz52U0VoDRxpYGP8IeXIKSBIigmcH76ZjTjjm53cCQuDBY
DAc/q2qNIBtX+Qjh0oVkENCV93xRN32BnMsGVqq0rEqiXZ1KOCmC1fPNHryM0HQTTy60AtgKrOt/
KUhV2EIJvIZPBHS8uCKYm039/D5LWEDwm3u3NJiywv55nK96oNVk/hZ8pSzoA/z3vfqZxtJpFF1C
uSQLD32rREvRYM/YkVTmVLlqYgOQ3NCmh4lzSXP9AkgYbtnAzJHCoiCfFAIorWnq5iUMUuorUZkA
KeCHb35lQoontRWuUknmpVeMfa2sTa37PiyEvoZdhLWt/9K/lWgpczbZr1ZHUFdXxtssmZeFudQ0
3L7zQ3y+Kg0TblGTeYOWCDtLHDubbt14MhkAGM3d4Q2SE/rjGbGA0uZb2bGiMN4kATKjeVp/pWlY
XlodrvC8QmKQcXP69jaVv4IVUm1wDt0wXG8WHrtabIAVPd2SW5q9wUehApVezHJf59ZBGZ44LSUI
dHkhYBagUHdcGtUPuF/zIqUiZVVCHUmPWLsLkDEM9tleddaabt5TCF1LhLjDuNjXnP3RA54zIZCx
mLS4RwuDsMG4RnWDJLzq2TysfhEOxMxxYxPc3YEjajDUVC3LzUxo4czSuJRU0TFxRrAWL6B1HfUe
hs4Cg24rpu+UtZYh1TtqawRwV8FjxLvkRKPbmubTs5UHq+rnBulrurBnwrZ7ptGneUw2P7Ez0nZs
0o2JWQMW3KoBGGWkikQaAJ32TRGBqheGwNk7ezcDM0qTFhNA/mR547h94i1YsEVWqCTmnCKkXZAg
ajfmli6JSWSXeeU9hszt1OGVSbHqa/hxVRtcPPsoqJye1WuRY1gDKyjRxczMQZE4sYALAwO0PHW1
BYingjBfzAoTbZ0ZFsmHmdxgGvq2pLYpfudZ1XGy14VjE34eHaAY5UpLj5XD82BjzJM17xgxZ3yQ
s70D8QlYXiYY3f9NLLktfH5qQph65bMDrHVfYNDMFJPJfkOWoLSc4G/1McaKaVnAFpIomZL5zQ2g
gK9vjdb+505vwAInb6hWGVVwkGUdaHAuHcTb0KSHMaPmScxrESBWWT7wyih0ElDkA3/KHSnV1KPE
K7xjORbs4wFboPw4KYFmOnpvA8UNt9Rx/tHUiKHrysdi9jZDfKQzH30lQergi34EbPra5jR6EphC
Wezw4UlZJQBKI0OGZF2p6gyY29BB3goAaR8n0mdb/FScJ8Fejk71SWG1ahXMwrG2zeZmWYOv5pjv
jEM6IgTopv2y+B0tRO5UvAEbmi7iQDuOsMnG+8W0aGda/CwPTdnESdNY+mbko0wFU/hHi5NmV6wK
uBCvw+5AyM845XnFUVjA+cuNQovfeCIv/srrG9cr4k/DG/LViV0yGcySZyydm1UGC7JyCvgk8Ifr
X1K5gpJLAPNVVBBp9x9RL2iX6XIXmyRMevFZMyw+aX4IFpDxFTOjaXvRKV5I0xDax6Zrf5Ets5Gp
Xzd72Io9PZAgXcFBRprunZMjRh6gMQLFSNCXsLUnXXtn1Ao9ER+2FHBZ1M95/MuazueWyEctW2jp
FxR4twiM4njpy8kVvY8K3NfWASNSzvMA5rcA+IntGYWGT6K7v5494mTzAaslcJDk1zJGkleo/z5/
feERGWQDPnf2Qs3PuHOyTI3Em+teoCt8T/G8UKJ/BKEFIGiCdxh6JB2+0vRBQ+Mo0T6C5CgSKiQ2
bCGGtfHlbLE2j8CpVLvxW8hmFuwvvqH5RZDfPUfkbzfob+Q4z4epNihX7nJH0y0oPqWUVJa12Y+p
dmahscDX1Cuuc/lN5rtFvzbEFUBLv3iwppFgDQkKD+8SEWwFlgNulytv8qYuRq6vU2DbTJG1CwPj
MWS3cGJyA+DBpjkCLq1ohwcBWbutNlaWJt0mk9Er7eQ2FulyykQSjUVIA38nhAStvt+BjeslqFKG
SLGfUimbZ06gd+k6fg+0ONg4+HQV6xv3t/UmUdKjkGDRhFaveI5cQ/Cgu8u0jcTnHRdKfnFc8m7s
oclGc4bY9D5viR0lKazpHBUnvaL3o905ipyu4Y38Cahgz0esfBEj2zC1q+LRVz9k0ySQlTnvYyE5
eyf+HQC+h1DKP7lMfcQBGbkh2Tx24rZb8h2YxoxUR8sKDbH0kY69pTraYqu8hRfBSZcuzIJO+kVh
WAUYwwvx+3qMQvF6j59M4a6QpSLElTClaIUrWIdxcLOCrvvTP4xdfz4AA4KGdCrhHXi6SU73G1rS
ZyU/3uH5q6w1HcAbNMVWOtzTMiFlkwET3xU7O3qXq0NfZpiegsgasOov5+10bpXaDoMSlZmyCa+7
DNhVdZpLQFzPNVYh19d9LbxDT+2+xPyyrKkDVapPp7csNjqwhPTZLkzQuQctASbQXsz9DhFSKn9P
ebc7TokyXZQMkrUEA+orzkW0X65VGAh9HkVj4btimRdm7Te3QGWr9N1QK+5BG3226YQLOwO+Mw/x
+/v3ju7pf8sveNw8Xi31qfloIk43s07S0y4RERQmIxAdV6DGBsFCUYxP1r2scctEqhkEazLS1Zgy
08i2s/AWbOvcL9nfOxFthdSA2dgu3Q55esljnBSCHPAArTuQMZKWZPkDD6BpHQb2UyWCMnpqwe/X
FxRzdZ0JhqzGJmP1HURq1irdCEBoMWEH85HOjmnGFyCcbZIXPhRo2fRfn446NO4zLhfloPFk3aaN
fXOc+/iEyscjbggGxys2YpU86sBLcZ3cyh/WCReFrM8N/XmMZN9xE5K+WhP9j014I3j70AN+mHZW
Nt+Ve+Ct4NEDbbPJAnVpc/5+0rJ3wwYg8LhWCWbOoaVk+c6jPA7hJgQ3s4X4yaIBq2acSvVE8a4n
S0byZ/DIpFBxe8QsG5GNuDoCgOP1VcgBwlV9ZTrUdN1nzC2XkmSyBEh9trUCMXSwpc5L6GiuwYBB
bRtfLKsqSQ6o2Hs6eWbZHTXHOPASnaWSX7tGJozJa87vCGNQBaEHdXY3Jo+f6oK4Obb9mykVJTYy
Q/rVPDmj5M3MT/t3W8t17A66t3OYUio/IniuPNTewD8AND29JZvWZTClFqsKOTOROMYTAq2G1Y8o
0l8LYxuffAFsq7/i5OA6b/xiWLc3obfmD7LB1GE6Q3kw4wpF/h2zYpU/xiOIE+wjtlrf8giAp+lQ
P2o/IOB7FSNG8kdVBhR1SGQtuZmOOmIMOBw0KqIw0BVyXz7AXDCJ9YrvpFN2mZxeJXqU6Jzh8hyd
ZVyU+hR6UB4eoG48qXE7vOuc/2V9bc45xfghk5f2QjODWh8noGUiIZl/7mtJ0hGLPm9a0hBAcS7Q
ANIqdWrsOpssMuK7im3YtKZBz/CNK6K5gtFeDDW06JFEQR6T0j2aoPjGa1bo3zCRN5usuIxNlZwA
AZGuDz5K8I8+gPPokK4hzI8RBUKlkspdjNsI3ZrylM0tHEGn+ums5DxO6miklbUaxEUl0J2uakoG
6Bk+zYDSX8hk23Gt/x8qTD7rIMr4j/hF+WnyhbgkUGLvcN5HInIHmP7CGuXwWIrtDZweM/pOKIXC
tA+tBHEEkhAfPA+vOvT7TMVy/4g+NWvTzIP1vL8VmB3geVxd+Tl9FOBkqfRIFh0wmMIzcVs6uQPn
5dc9duQvyrDlv0fWDWa1HiF+sdck310F0PemH1XYuOI+8fMB2b1jLAG7Zq9uwD1JMqRDX+eKyBcF
IjT6eRnOnNZzfljSDFGflbhLbQ9PVPnojOrLwtRCkGAHQkBLtpaJu0KZN1Jxd86QYXfgTA8505on
gkvo079byCfTWePsfteLAyQAh2kgWh1CL88au/6rpMIBWT5G/RpbtuG2yQXcvx06bxVggmXGIu7t
vcliof8TBoBT0XMFW1amXS2mjcaQg+I6pU0XEV2VFHBWRzHWHKH1GSQp2yhEb1q5oqa9rG+1SoKV
rVl+ynVUhe/TF2BFr/bwKrhxfaY10oA93P0xRWvGa3zjpSU8shpO2hCbZYcekag0koiHGfSJpdK7
hFBuNH2fk+SLCBwKTMFzYlaMlQPj3FUs24ZW5A7oDFwjUPYt1js0pXWFju8GbrRaBe1QsrCfOCg4
Ydf/2YRrwTyYSEUfW2mv+hDJwJ5eBsOq4knBi08gkTDTvpNTgcoCcLZs450mZQf+qUOvapZGHGCm
gGny0zKa/hZQDJXnWFkxdpNEP82NqN1gMmUueaoSykuwHxpwiORWsPKnql0An6FpMsdpx9maZ4gS
Y5KqY5jLA7Rcg2zBRzjVM00W/e3YAO7iQp7nTsTMtPPAWcsLvOFWHDuGX1zX8S311hc426BSJ7+w
PmvayTIUgDGPWJV1ifaXMElWN5q486UmOEgt4Qe4ZQlEEe3WK0S0aA+Krdhw9sSeEW3iBLhW8CZk
OxCFQXL0KwttOQkbQ47N6wRdBa92fESqTThUMO/ZqGohY92f+uH6rdU7OhE3IglAwU4Vi6iJp1D0
s2TFo8JxDTElHdUfuHFsHTPKIpaBfJRJG4o/mh992sII3CJyLrgjmiUEGHxkMqLWynKXETS53VA2
bXk9cdaPD1PUImoCgMi2zTHIAq5D7+tXGijLRcIlyyF4pEgA4M/1bKfN1/k7iWM5P85fWr/b2YBW
YVe5BIu4wgrU25/xhm4+OI3YsO19LW7j2DdSyd6TXj5mkBDAgcklLhYLOcKwBTWvwrWC6C+nwJZC
RiOP2Qhwz+NVPKrcMXn0qDdYRilreuge34MSAOI7xikASILYg35zYz3BsAaemHkjZoY1QdGESXMv
TJVJHQwP4N/r80dk5H4NAbKQri03Jaqk6+AYdA1P0r5LchjBMZu2wrWW+3DUEbZ6WUxMBH3e5YO1
///LBFuwv85qfP4l4lEzYCPq4SGPW0qpkLZvQIxM85j+DmcyxArr2H4C1TFWgT3KRmAsCt0L2LNU
D9ll1tGMj3VHGajtK8ZPRQuPXhIpFDwyNqvwyytYiG14tT9t23wvY0i+Bdqz7oiu8YscF5pXaOxg
Qj4x2OV+NxVGNZ0P/I8UWFftuDcPT8KRNeI4wa/nUzxmpcScO/bYvMRlqECHD6wYRBOEu9ahcJBn
+ZXQBzu/cmAn9ky9dWjSl0qV4wM2Y3YVnrvo/zTeYaepO1iBunFXW18i9QpSoTOYgHDBVOlGC3ex
UNqc82Un24bkO337EI1MxafcmVZowaOgobWW4AR1aechkwNz89VZvA2tbcr/sC1rkIUFrJ3WZ6eI
dhH1zLgphyrbGtb9WPgzBfenJ5uq62v+orTsbsU2twtVMebiyTrRuZ1MxWiz7b0M2/3zsOq5HmRT
ct6pdTqdOJnHlzX6VpnB2QT2QY6Z1uDHNw2aJK+zWjfB/hg8TUYr2+jCY1sExZZzGat/8TfHP3Sj
nkcaBl1TjutdOJ+VVBETNoPUsRipwTpbygXEy9C7/qz2bL++OjrIQaEytGI6zPci8wa7+POH9sdj
onA/4pUyEaENwAHpguufE5c/Lpo1D0oidT9+dc/KIZQEFT8FpngsUv69ynXvXaqzG37JQ0y7PQiY
KU7IqJHeUq/8d8IiYXl2PVPy8CeARqYvnxUtQUQP1v0k2RosJBy02sGjvQ4FISJC39sX1hLRgQjX
NY2C1u6Ds5zbDN+HtW6aG9dkjHBk1pdmShR4S3HFs/W14GyOryJJ9AofQHz06PGw6O2KxCFtJ/kU
XxBtEjd9gm/Kf4mxBchQTBXHmLBQB9lXwl2W1ZJ7yLV8aVmJQTigPM2jhoqvPu7iF+7v+QxpgqHr
R22Z3iQuXGL5g1XDBvBACnzmp5J63SC1YoT9GZgNMhSuuP2rgkA4bUGOa3PfWhme255dTIk1JmCa
nEV+1lxxH04763iV0t4K2V9O4D/akNtoGNRsP/KL4QrLtBZG256VuIgBZv92OGTIy+hBMNbe3Q/H
HJHoJq9/xMI8Kn9o0NFip3VD8J8dtalF38fsMH5CTCP9I/LicE+7kyLiwY4H26N9FXs3n3Ac+X/j
F2m+Sdt47S+pCyaQnjQxo+2CXAsYAPITOorzvyI8KYUhAen826iO3HzCDXbEQoDFmkrmgdB3uROi
C5Xm/EYtyIc+6f9ft6kzRRPUWYhNncJT4OvIh+5fy83nrwhkPNrm9+MKrW5JfqaJbPo8CYRq0nA/
fUCCp9/zPHJlaIavwUs9QUD0p1MDQPCrnm2je0KDx4/Rz7gGWVoTWg6pbCbRlzwRdlh3VPG4CgZB
SqIFWdogYu3eCqS4l5bV7t8BusjUPB/J6frdW1/s5ERs2G3otftbDJMJqiiwlRZYlA2YZm7rwalb
jP29dAiSO2HpPrxzx10cK6xFLAilqnmqKwfNdWs1fHBSZFzQ+63srBWm9niQrZ17kuChsSKHU7gb
XfoCg0aEydjr300uGgnO8JBs+THv+rUPU7NLlmADBqsKuECNYna83ZNBHy1lzPbx/aVjyiP8N+bB
VljCPuWYb3HlDsx3S3BPqRvl3LL4NookGUh901W0cH7efuzMz0Ubb9flqrGXOTCWJ4bmIP/7LyNM
SECSF0phekNLTB9vVvlnMlieU9KHvtnKSHQ8H5IJ/a9OLZ4z1W7aAQH7KugLquPHhAPNgNUFUP4z
U+UcavV27I9y8nDSffkq54WxxKL+83RRGAAzFCw8C370Mn2hepDKTQ2dbeF+rbkEgab76iBEsdNT
FGzVCHBskJsH9mkaGBkYawl5xLT5v5Tu7XvDavMOsoIWky/3OZGDKLSiLj06cXbvKxt0ZKSSqv0Y
mlzvKUzCkdc5tiF3bASZvEbglE1d+mx/ZzJ/ovrZF7ZHRtV56sAwSgh/8l+VmLxGja/hRzYr0/3b
2Vg9COBNkQOs3tBKF4PwPOe8UD1nmdcHo1Jvmb0AHuIbEVw+BgZQbLjn2o5xnfYrtoDCI7XNG9HC
uh1f1dxtgrBDxSZmFaPZ1YQ4PMDJXvb4UWqXqXh+MAalGT4dZNRR588rl+fp1oHb1VpxhjmT4q5r
QEl5h2l/kWGzY0rCMhZD/vG0FxHoKvQXjvb2tednjjPtxbFFU3TyrBNkcZ7vuv/4F4ojP80m3ls8
jj7ku3utr4aBJuC6PXmXdIIYf7zHT5IM903VUS0uT2NnkXdfTTn3JzHe/2BHGNkr6RowGv2IvQU7
F6ilpf6cLlE/onsEPZkHRQdcVOW8XLfeMeWgUgsw09S1TRAcbtR5wD01V+kNMnZFbP7EqAVi9iEZ
yk8MrQOUyYE2cev6R01mkiUTyQj8LaOV0caHhFOM0FnXTjCXpATBitRBgVAJ1kPt7LYX7U1d3g6S
y9j5PrRBWK0L7vx98Jb4OQR1xy+AvXJihi6A/ug0V7yg1pe+AQBhqvKjoeH+fFDXVss6bS7+cyo6
xjWU77UbJOuKZJikedELhOBAP10T29ttd3QXXsZuvar5VHcgss/YYPzRhlCQOXBRpNh/MUrp9yFO
P9kEbO3f9DNBuBP+ElEQTQRiBMk3vcICYSqj+wVgKyz2IWpfR9KhgYCnBcunXz33aZxA7m/JvWqW
MSCV0y6sspnjNPhdN79xfHaN3WkWGWBC9T+0CpvxGGCFq+ZpbDfynPUFmBGGeuEzD3ijzvt2RDZx
40Lgto3vTTIjQA0ixRwT8C4VQW1TfEuYsCDoC42uQrc6yldzPAkGxykh0kXOtYzWkH6XItn63tR+
zdrjZ2bycApBjZUSfaJtObmXvJxYVJVHsQp/vrnDTzxmmSOeQUgMi1uqhLTfJPsjWO+3G+5+rL9T
VCQ7kHFdXfqo5/dZpfYdvuEbA4g+xBw2lkCzjmrz/WBId+LPTaSx300JhWWaX2jbWOosgGpWKOU1
owB3xPExW/zJPVVxGu5QDe/AoxB1B9mz7MZWSELNzARQQb2T+VFrE1EaEO9n6sNugOlKqVFH1o2M
nhW+EeY7xkiPLGw4URLQlYXpaFiN2qlRwUO7nMUTGlNrZ6BKkGfCxsBVB9b9ak8S91j572vyH97S
kg6Xc9hR+2jQ5aIK2frg5/Gadlbg/gW1MY+dOjiPHpATj2s31F9LjKTQcMUKF5XaxygNwNO0+5L7
f1RCdcuLyhc88cVOv7OXeXgnfl4QdemgxjaTHJ4vwEg6aHQadFVh343HvEJ1qWcl3T2E2Uv5FZw+
F6ErXSzGxcF1JyIi29tkPAk6CcIcWIIMxhEkZuGu8kGK4qNP2jdNrX/mvToUJ4h9fFT3RM9N7nKX
VdgW6shzjWptH+MifbxSQ1TZz4T1Y/cPshkIqaN18cUpFPiYngEJs/+olkUA3clrEOc2H1ZJ9p6W
E6kwIA7PCnNeatx6VlN0Bd6QKuVEbgaxUTSANsg+64eGLlqtWxYm+tYgSJfSJ6DDT2XwOIg9+bkw
pG691T/r1FZcMjlY0j7wuYPBVFmztsp9BvQ0LoPLeQIwVcjQszY1s7saJMjx3jje8ECdYdTg0hAw
a3eTbzdrkMp2i5/zXqGKsxI+C+TrcOLSS6c++6NTp8rsr7+X85NWLNQXGwrU3ytPU2IS+MdlsOsm
FIkLV6PRTHtwlECUQQ6yCWjlSeJMmGTBaz3N2IqMZe2wdMNFW2SbamO8wWVHsA3BdB3CUTxbTbaX
FI/U29W0WM+IEnT2dE64HeszO5Q///c0/7MVa6tDFsR9BcTbOPVW8W4Tygmt6vF8DtKhnfpJGgYI
VDEHOCp1daR5CrGnpXjwJA8npgSnm6SfkW4Xmes/ulS3wPZdsIUzihzd7r2RN0LtO/ojQs9JVrTP
T7dIycLK9LgqjWJ36vPyzO9t+v+Kxqab1IKk1vfuNPOFhU2hf1y2U+Y+lUO428xN5hm5ZWI8uvhO
590ebtcDLtiSHpb6QL50ALXx8INNTv+RlRVHP5LTmPvaxMvxZKMPwOcwr8W1U72acxSQRTHgiI3D
aXF2nB5ZO15zSSKT0YvT7ddA43dGck3l5T0G+COBjgDLmem+3K1y6GLv93dw2T5nXrYTpSXPb4v2
BdGt7jQK1VuEQ6ZsecshYV2AV8B6ijaRi05dNKfArIEwrJY/QeFIYKHU1/GtSEXHLwNtOwZXKzL/
325bWCaxX0zVRw4kfbq6rugKlzYcPnGQ5v/z4EtbDD4nDfmaRLphR0cBsRPqBUIE6hXEbm81bYEH
ZbKMWSMwvNckTBP7sO39itVKABe4lumj0KKiX3BNFya7ptfddgpyBR14Awlbw6LfI9S6mXbT0SMo
AAvFw4zqmfGMReNbsIvwZaqDHv5YQwfvFN/VlReNDOL/nJzdZoVkQhyww1IK9/qxHkbzswX6gCdz
YPhAK7Y/rigqp2xGMinO/KXr+2Nn2DAOKqbl2vFt4Yhfk9k/Bba9YckNWDtKq/VwuUHvBeU6VYUB
EsH44Cd97kvgQndvgdQZP/P8hrdakGRhEgkdTJNYLr3lh9HjxB9hNVSmYwqoa628J4bio0WxVd5e
DvazZWfMaKdt8U7779QKLSaRbTg0c4x5MYSJzWGx8uVUUrjAYsdr2/TJY9wYwsXpy3T9VYoIOi5n
D66MOcZADh18GVI8Q57M1vnv3ZoN0PQPhRGcVGhZ5bmIwCZ6Ffe1IkJJo9jNztKRmbJVpN0ey14d
KnNnaCIqzd9uqdwyCKfRw84J1ucbF6J5SVLCGVPHCKfkBwmMpFVOis/jNneebyqfSUlrqHWcfios
UzUzGBrdqxgwlZI9Qoz+nBE2JlPtk8EvoaOtMCvRCktZX8xnJD8Jji4eUdqTtNGqlTVlFtPLyyQG
OgJm8j5dKQnrKhkf66KkcKKlufgCQjLIcHKu02HEFJdFFUNCsLNew0haQOi3KaooafCVApAA6rOy
5LHDXAnBpGvMX5WIt9TIlcmOQ/k+qyCXIxyHmd4aiGTQHen503lj95fy+RgvXYA9vu9WKFHZbGxR
OSKFy4+1z737KZh2hgmF3byq/AKyaeck16xk3bylHgyVaLVVG0vvy48mUqBHIEp6BhtC2RA22NSf
UO1o2YDUhiEQnat5KL/pFqpRFtdilR0VU9vr/fGAGEWmq18itwUfZhCFV9pBPDkK2yHvf/63H4ai
r3iqR/L5q5HOjfh2I+ph9/z26Y6jGsb8XcRcFeZIXvBev1TFPduxU5U6dQzjR6pX3aBsP/bftBtX
MIpLDhYk9sCixrpVnrcwJXGM24Wrb7la06jrPludhG5HFKwXQ5vEHL2PxLfmNxm5vI3R4QPN9ZAU
pE5OoXd5DYeJ/B7VkYL9mukcP78rs+M/SQxCvAwaAYAE6InOm5INImuQ2M3hebhkDZzDa/1w4Zac
StH1rpYCRdIM1F01kjvOLjR1hlG4dxDHA+WBtjsHr3lxZRHjJU4y1/uc4Cu0twsun4+CzUeWumtk
ix3kSIPj15o4jyYGx5+67mvk8WLrKtgbdmp+B6gZuXP31rCtU4iPs08EEODmcmL6wmhoSRRINOyx
+rXW2L3AcIxxeIi9PMPabKEcuQP1uqC6EY36z8qpg5jJbrpF9gB2YdEWu+y5PCjUMG0MCxBxBmtE
dDM1cIVqzm2AwNJod0O7JdrJe0AUm2+I6PxavWetJ4Ysbqx0Njc3JSXH+5vsZPz6llRTZCB++XzL
DXrfKq5xVklUs6fquEZiyKu/9Zu7Dfy/IWlhJ5m6aJUNZKoc6S94AiMTeJjGLV99TYJg4jaXQ53a
DgYUq3U1aGVHs2o6UNM855U4aMvPfTxOcs9e701R+wWsxmXtEetAfTm4YlmAomxSMrYg6s8Q+8pq
/TeX4jR4hO8HBFVlkNl470NM0zFCayTzPrITexq34ayxc9RpuMnMKkTDnGg3S4zTSjmubrNCgqqw
CoASEBNT59jgkTbXZwRKU3WDAJD3F3eYRzLQAWkUTlMKTGYBNQy04pSLlFJ8BvgW/Dz0p9gdIJAR
RUvwwGeaMfPlP/iqSTzm2sMmb5GIJqvlIIS1F3m61pka43QjjFW8aSo7tb1u1LtaG2S1PRxzBOB8
RGl6Ddp2VKJogYhxzPvplnjriYHnaApQRHClSOfU81Os1UAz7hRCuySR82VDSwOF/xBYsrpV/tat
P49Eyw4l+vOZyefjLGB8RqoqymFJ55FpI4gbDcMbRsWz1HK9tujc39dneRufOrfv6l0OoTS/fvbw
w9812tprRaMuOfpoSPyQA/uktqr8N+KubgOZYKlmd80zwxCH9nHo95KNIUIrIMrYX21L/DBQk0gG
j5Pk0YS/HV7q7qjF5R5oBgMa3ZAcjAPa+uxpJZKd01VAPjIuT5RO0AnvdG7C0TPbI37Bc0N6cODW
LFfBn3zG0zTM3QfTTur7qd7myO2PmkkubK5yhY5CWoBeiDpAH8r1kqqduCENM9RJppnxot/HXa4k
rKYsM2TDSxbC5LY+6WjuZutGDkTINftFAbFMEI3yXLzSO9hf2xm+idh42M6q4bQNCD0iuqoj3vX9
MfvBkaw4NgoqpJhJvoVPKyrwAMwVckI1K0Ps6tktb0dBTQRwsmC3wV3FOfBGI3ipHbKLYGGL4rTG
ABQfN1R5AWQAgy22256CgRCXEC7LuiLgGJeYRiwpknNxuytyPC5jktOANwbMt9KKqlFsaQV6qlu6
BCwdfNCDhqTzb8+HBViOx28o3G6m3XCOUeN+GpxakEMuO/HDWNa01Je4avx3e90iu1YO+iHJfHxQ
sU3crH3npsjRKqRB/WDXYiLR5G1OruGDQLYPZcL67O/ps6ek50xrIh6GksPmOJ+D4XgFh1Cbso0E
7DbrMRiX/OWrcU4coqPeAi6xwYs49WIyKvM0ZAUalqFyETqUzxcKbipKNoHPwRMLFOrHIfktesWZ
QwjFerjM0WNd8kfwtOhz+xHCDLZjCnnb2izRS3sllXTi+Rvjyvvb7dgAR2KKlSPKm8ukIP1PMDOp
t93tIGo1HDeE9IX8hPqQdmUbNohcBxz5mKcRK77bLUhre2rqy4h6y0OuItHuaDhwhDvz1NIcn61I
Gssb7HWPYvD299l7kJAkBo0tMlNm8IIetGIQM/d34LQjXrNDF7i/GJv+HYRDU0d9pjgfD/eqjzJB
2rhtNkZqRegoy9dXsP/KvCkyf/aF59okw+LPUdHkAKY5M9bYdPxYxHVYGBdcq19/pg/K08VIehlT
CL6x2A4lhF5PnGYABykSfRa65YMylQaUWaK4yVWiNU/vEvjWAZHXgw5DN91d5K2w8B8FVk1rJrGj
K6T0N87ITLW9F/vpAP9v5ymln2c24MB/lYNKdS1mEUadK8Cshel37Re+enT2UASUV82IhrNTcqw5
TnXzfGRxfqUoA/e7VtiKUsiIst4/MQF5z2aNSDXLwWHxA5zwe63MTTye28LuGZRiYdn+TGeaxhT4
iqDkC7re5jgMgqC7VohFaE+qxW5TcnwY8Dwn3EzW0ETO2eX8H+X2LkChmkxRSw2an3/sH92MW178
FjLAW0wFGQXH5NA4/fH9KecoaC7RPaHmWIcJICWPnjxs7UuzrgWbUDAQIc3PH0lhBB+Ek9RTBNuT
QRKbR/mQWF3NzSPll9a7fPxPL76/eT1gwevmpNs/yqEVrvdAylXf92QykRiJ5+rx9jI5vLlWHEAq
Fd7l5fNmUDzNr0M9SEgfEcyQqL5FPNf1DoNO4GGz2EpLV8hSlW3rJwDxQlcUh47BdB3g6U4zViTI
lLef82bg9MIZezB41TxTu4qq1vagexs69faCpxP7EwcGBDqmzq4mUqGbWh5srSeFC0Ef9dERIlt1
lURGEOkBWFsOe/50CABBtN/wlIwrAFJcVzkESL0Av+pqFXsW0wY/Hw+ThQF86RdDaQkq8av52F2A
31oosE65bQDfNOIrB95YSdgNcKpqSuzgzbJs/bVnZUm/rPjBHxYxWixXS2SrZEhzEeUHZyUHnX0R
a/a46jVpUcETmYXRSzGHMOoLYtCbgq1kkbOhyORcbmiwYYISlGveuXI68ZhS+E9Hg5LwOrM5zhqM
Sb5aJLDERbkWiYy4IScTFygcJCC2JwlRuibCAVftcjCfkAFH6iear4h4G8SwDEQQezdWgOkGl5xu
X/O42HID8LwBrzyn8Q0C/h+fLZqbXKnTJ2OJjngiZ/lwqMQrv8WPP7aBzuOVGFuIYWCGdB4HNSIo
2Uyp/Y3wvU6KY4B18U6oC7lDzg5EIGYZz94rBhjJxEVH/x/3fBaQDV4sGfeM/YxQpYLKtQ0S5F2e
tf1Yb0zhMVF8p6JcH+dWV/4Q2ax1uHiDWEXfQAoCYqG9MlGCj4Iw3RyJjp1ps02cR1l1dWXMJ+Dx
95mr92L9VP2RMmnvNP3MJyWGG5q+mKzxIyn+ztNBDS4heFqbSg9nVwmhvUc7vlON+6ld3gKX9X6f
D7jJSeXziwso5aMdlFjPIP+F/sEd8pBHJgmF+y4M53uMluSWRqXXIBEZ/ONBr0azT0YSbfKHdJAc
A0hUmhUAD5BGL1ZSsf5DSOgqATXg4XH8p1z4qKFWmUb4lKNqA6k2+2Xz/GALYAkSOlULYz0CQos6
1RRGbjC9tC/elsXLeyPTurDF33LjMLq/dSonxuiTWKw8PNzXI9X3K6HBVK+wLpjFcNg5KWKx07aS
BoJgH/Mrqeq4KVIF9RJiyTDJezJJqpAsKPzJ/u8b+w+7Okdhlg+OCmWqDNVAoFJkz2xoA3dCVuNB
PH0C02uDxByyCBkqJic/JWGoR3jZuGd9JGuEc0IprNOXq2MIfjpnAWy6GRR3U4UYUY10GQQ1da0e
Ly/CThgNPmG7SjyITk2mZiuAPhd76hfqVUGunF8He/P4xdhBVqZxCG+j2SbzQiLNNNMKKTk4O1mn
u39gO7fuJKpvdY/jfi9Oa2TaDZRcD56lX3APCBjnPeAo/r70FJJ5VCU+7MCFnfHpH9dReOdLZWQB
YLK6t0Ijn0p+J/wtmsbHFxjDcNjwURGf2kWnudmwmVj6+2xbGOP9XMZ48ojySgSlNaM/tyAITyGF
2B7/HhfVOZnBI/8FXsJewkJU/IUVtQeWJk/bDapSUz42oDOMSubu6bryhKlTP5CW35yfLiyT4qvL
Adt+sPXrsQ732VlGcTeoNl85GwdYRUnNgNCSY76S8N6zGwlT5LLwgSr3oBb2oOHgb9wNr+4iYp4T
se8AC9B6zxbpjIJ4+igqGZQERwtrhC3y6PMpdc/iwyFi+mjXQbZnayRVoD7QX9Yo8eoZyYEFzW5i
k6POFDX/B92b9KBqOXpxhpIQrPlkXv4G6f4wStdNXzK6zpQ971RBRxHZvu9AjErw4vfu8cSh53Pk
p5tXSN7TTxPiPTp7/XdNT7IKOBrpw+3+sEKKJnsw5Fnyf8Zrrn5atMmRNt2wsMLMRCVFNMY/s/lY
tMn2OXnSEBUw6Fch4vDqckFkgSBmMNrXL/nXgVu0WWbfiblvCpe4vy3ImGko24Stoakb+Gg12Gz7
VWKxfCQwF5vHZvWt6edtJlfNrorYdQJLN7jXANf94KpKafmdTzYZV3AvK1mYrdsMSTykJhzTgKOn
RlbnsjuOkKdo8BO6/ZzGapRWV6WYwhgOsamG8n10QK1FANL8BLy/6Pzp5gHx55u/R/3GthW07AzM
OgFNTiAXJurW95N2dNWaj4g0MwzveHT8w6Cd28Fq1R6IXqHev+AUjL0SyOm57/dPvedgn2pTBusk
i1vzJpbVb5CZAZVmIGPWZZWSuczaNMf33IKmdWJLGuT6tyZI3QeR2sdwf2nySpa+/ZGyiOynpdFp
TmEegBYQkVl6u33xNEuGiGXohKNsnS34txjAO71JT8KkI8O03RaHf35NCVHzHliicUIypSGK4dTs
3Nb0BVtZ3e0OHichAo7bBOsPh6EXPcZVed90wIGA5C0cSwl6cziHWMJjy0w0LwIzG+DUcf8BTcjJ
iPC9MN2xU3/4Aqz6Py8alBDY0oRK6AnHxFGly8AjS5XOE9sNEYR1jh0dCoUkxaZ8cabpSC7K0+XI
fBHjNhXz1P9R/eyOPHDCo3BdoT+/hwPtWBcLOu9M/pFImrZraTOlWLtBa0ksPrQt1ibard2fP6j3
ko2Jo8LV8EVHHLCRcmQgnwbdD296Qy6PqADM3l57G2KEmOWu/wofnsR/+q4mCD4ehpJBNI2Z5S7V
i+rswYHSXt/KdGLHnMQiirlCNFgsjkUsm32BYODb+1nRAZaAKX9tx4zF2EJnhSiA8dDDKvs0Pz2J
peIrvUj3YhsWta8248RaB3TRcgQy3VQLRiNiJY6YmxkbJDYxKrmI28zRQ07MHPQ6uELbQStJwFMT
bD2I5A5z9iEhgfNUPIx8qunb/dt2c7J1P2GvONLM/SuPL4TAYbCBBmb5CL8TZKMLEnuAQWVrY+IP
ROTJaLRkUQISkbD0REZVwcWcub3NKagj7UqHgvgsWKsTEXrFqORtaGPKyoZCqp8mCIZpeDmBbLPR
KhsnPDoUinEllvZfl/f2URRRFgQG3oH7CAjT30+ycP4NcmQweHzZ421kol0lE0Vdt7r4bvPU9a+4
DlQjtnFirACZ+9SNhkNhUjXHFprM4SPv0ZC2ua07TA3kn3jfbeDT7ZCH6Nw3ziaYVn7ocuxu1DBe
0lUZZpyoJ99kkBBnmDQlpUXa4gvJIuxL4F68sTDoob7fFrRHs/4+lg89dMwF/fj+QbGFcdkplTTR
m3+jmcETxgcQVu5CglF3jtB4pwmySzlrhF7BMi3Ltg+o4gMiq0vl4sH3Lr85QhlTBiC+s5P3YZRp
TXkoLrmdnXqYJdAlzwuAY/QGfahRglrCFJU/mIPt1XFPUGUHICPfPM3rOy7dElYRvz3/36FtCXV+
+fAVLAN2JxLPXtyKoHZkclnwG17ecFpTBMZmbYkKmmSDUPFS2ro3qvmhHQs52WH5/1tAP4cIWlux
cBm/3gRUzidMrbFs/u7vdj4XCnjEytBI8ywePAzk/c6I9qQhokbxa3FDX2NE4eqrVAkSuPQgDw8C
yn/JhxDgzq43l1Yxh+a3z8HRSiEmOtxYc4LnwkSFNKmnlvOC5hxoGkAJebjLemaWqTDPvIwks53V
1vZ3xYOjJrcUFeuz7XnuWfaS4w44iaZn9b8OxKM/jb9MCzE1denSvwwDFeWRFbrPr32biMwSl+QE
ASlxS6fK4l2zsfPZOhQf3/OA8ehJdpjdrIJ96Jy+gDmYo1VSpICgF0aex4KBMweYXHJYGLTVLUBP
+5HpccK9JPfBsr1dA0R9YM4i1EpD7DXKnuwaf14JnvPB8lpfSQbYnrJ9jn/AXBtQj4HqdaihGfeo
mboJNexWYghiUHiKgZAjdR1bueYOC/uYLsUDwGAeGHjRrI5ioICSqt8cw6iVG8Q8vlZfwHrK2zvd
76HVZFnPaETFXaErpjU1aDYmtBET48Hm+bipqMSpICl40qSc5EO0sLTi5Q9cUXj7zw/5U7DzfF/v
4oNzXahS24n85BNFJmeCdJ39fhgyfN10HxSSD6IVIE2/iCpb389Ou3DzJewl/c8uo/o620ZBNr41
EESMb6/iXPtHpxq9kb9ONZv2JzBpuHxNaMwwkJtO/Ij8B1e5CdrbFnbz3oMyyAsWReeFzRUjC17t
BDZ4Z1OI7QJ1XB1TZhmd5P73HxkSFRdJUZJQ6Tt1Horxnq/x/pm/EvOQTaNDgvMSHDXCKhhQT+Oa
TdmxaYfZZP8+LtgFyqSw/xcHOM077x8vOF97v4N1eUUFbKbcifKC2sH1k0Hb29u+eNmhg7rE5/hY
UUF180P3yTTF2eBovwCbg/lqs4C1tw0nN8k5p8Y6k48stibxXHTjpG/n62bCvFt0XUnnwVZPGM2s
GpTOiEqxm7iHIKFs2J4qXkRy1w1cHZn8cTtQQnJjDTrvg9voU4+wSejHlq8ZmGOc/cw7yvDIzgxK
JZc0uEDN9p66YeQQkG0UqrOXhniHxXaVrmSy3wNidsd2BTMz4COtkFde9SkSbBGUTZm/DTSNJ/vv
s/cdIZMr6B+YUiLyIVLOdmuW+AfD3GtY/IICt0NuwI56IPfLkzp/A3hRHTM7TiT3ijcdSpKSlrx5
f2l/LhLwhgZg93ciCNtfDfGKYYD9OG2pTUmv7maYcnwMyc0vhnDxKVCtcQyWXjfV/CoaJakshgRp
SJdOfFvWABEgD2tUc+gpZ03inJ1U2bEHVaHZKnHolvF0UfV+4MkN9ZYRawN+ykiewZDeffdziSqO
i8gJ39MPAFzfHQnnHPQ8snmFr84xOx+T+wJpOGRB7aVrGyaFdjBdHA6deH3X2Uk3nKk0ORkI3vlg
YJKQ/SbWxyagZV58Nk9gxvAw0/fm4CqMmoTcB5LYnTQCtwcdu3T//J2t7OJQ9+cmtuGuKZnnxaeP
EKTz/VY8rQlUGPtzFFB+qkjOgXAWXSgcdjNuqseea1t5J9sVfhFauI0gB8auA3KL8J71zBrxEber
MhcA+Ap4eiPWylUbBMw4iCgMbXJVATwQNs3yMSewmw7pxr5gIPSOUCM5v0MqTmn+uXRLDBmDEDOG
MsRJRMCnfXO9PAzTo0D076RbDX6HvakCklfyEecJN46/xnwTjAFRxNW+vT8wUtl9cxCtLfWpaEjD
4fwF6IPKumILC9b4qvm7JLGR8TLtiJa8nsyfRhuKCWPiYU6m6zz/Ytvq+VXuoiFePGyZoq4X/w5l
QZsdcQzQs4Tg3uGrD2dmADxUEA/QZ/EvMTV2H+iWAiayBuV2LWgDc1gz4IarHOTZqN4lUwiferH5
S9G/Fq9/33bvguJ4V3fCM/yzS/lHJvNpwN8W0iYSSbw0o7xuox/ljNDBYHqCkMwVo2pTmEGZqcJb
IwqlMRQlhXR/cJdjFXRAGmDHZlUMhmulrVBfE0PWbSpxzwtEd++BZJondFZUQLJ/fgDpQmjucZB9
xXfNNWci/P3iw1S8dl+95hgFhkG/PQXc8IfV68XQgKegbZVDOdlPxy6aFiWd6QPJBoMe37f6ylVA
mQ8P/DbrIYuq94zakJityFHJEbGHCO4DmXm4Bb762ghAm3GkLmkPXNihLZzC+etXvUiyHG2BfdOn
/kH+mCPnAYD+trSkWgojyuyk+Y0wNknWmAiszQCXnloNthxHVbJluvFKoQBoPDwJuTKV6ApM0BnI
Y32rrm+nuo9DOwyav1pyL6P1gSBjW4Bu6zCPXOneZkGhiUL9SV0dzRMDCdmBt2EXIsZfXEnuCa1z
0NZ/mL8G8FC3jw2aU7X2af+cJoSlR1aWJFUS353pgHi4Ps/lVzUSQCz1az9FfhvOq76MqBtet5Bg
qekmynFdoULb8YWAI/Xh9+YVsguXa3EZGPg3awb7q2rWnfxpIjvJxQ/Yd6l5YEht/v6xHqmwKuGS
2mYb+yQ6Few9+YIJ2GxVdFo6KPh5X4AYT1Nnv/t9wr214C65DX42007uAshRAvi7gNt8enOT2ntj
OJBO0zOs+Yg4ZL9SCGHVsXpe9YWM9bVO6CSDinIz3vV1niZjrawruR3IGLGQJM/zBFeolNZyIz5T
0BZAL/MzElQ0FVpqv8STxBDyfAvJZ7jDq4IMW79TFs8D8xVopgl82WXYzLzy6PCYp4OzlNSnoY2R
E9mZ9KK6nq1+lMpBP48tcbRD8BFKuiR1kHlbqcvEcImfOwQHMvDAhmYDcnxgz7gCjxLlABSqqW5p
c7Wv/1LAisuOIilvNwBM/+O3kAXlD+Fs3t/7G/gatS7PiDHgldrvWsd1WlunhOzSc89+FJocJdMt
cfgBDX62nZrTKJ008YpOzyKAJ7ytgdd17MXavFXe7ZXBApJHaP9rIZTNgOU8P0IxJ2n8ymF/jS/3
K3CcGIAPGwAJREm1DjVOx7FUbBbIczu8gUixbqGp2PAk+gLURJ1ebviM9gpCdtJQpT11qKpYxoUv
hZVGWHj6uImozATJnxhhOvhXIYJLcCxOcRT7qR7GS176jDXN9LIbd1nI7ErVTrsLvDeAX1SqYwgL
YpFT/TVpd4NFmyLbP1LZioIdFA6NZFsr2//P5ioRJ2refDRHXoOgX0Quhbr8vfzFyMokFvEd2r7k
CWrGa8YjHI0Dh1LYDW8h3juI2+5Ug9Rj8ZovvrRuz4rz2cuor11TdBzcS3nIG9hahMUSnCaX/63h
iOgbY8v1F6RelPNAfsnFJdVOmuGZ9wpp+j6nTy6UqKYemUVd7JNPU3kEFUqjmEAWW0P5AxzrX+F3
oPe18X/cFJJwsHFoiObVMCGeP0bD9r8TmPiZoz17bZ9zC1cpxAHvaHWtB8YlgZ/2pB7IdAUGo3bD
9NaqaK9+HCQOuu9nu91rOt2xDGkTYpvOvKmPKXpkpQ+xI8/gVpqJWJYIa14AsI3niNwfPM0V4lk4
CKbHw3M5rfZzdvDtx0lghqDk1v2oYOLfj2AynlZSI3/RkuVChgnLsZHEOAgC07bGkw9RcZQ0LB+N
81hvcgh6TryIUdPG9zf9PPW9YRf5FHgXmbmI05gNHlAtlYUzeeB+gr3d3RqPUTVFgmN7VrsFE/L4
SFJkqbOKmxNzUQgCn5XQXKHBSY7BLC2MZznnb6XEeyiEEjS5zEO5NHPdpR6DUrm8iMHeIiqnPMGC
TNIGxBi9xWFzJjS9azaENTBw0LJi3LFP2B/D3JwgsmO9XwghnEE8XvfvTY+bIcJLCMDAPjrFha4m
dRO78tXpjUcy6O5Xkxk/q5MuqhChIfTlLNDHG9fKQ0a79I8eJUYYR5+srx4wlpfQovYst7Mjx68N
XPKgqUtPS/OCUbbCHBiANAiD1CnJ3j87tU9qDV+rIZ0aQxZkxfmc8ycV840LsxJhkR3dizb65xWy
rT4VzRYdeofJA8DCXyYNtR+TTGUFsnYsLWaaU1kM0AtWs9y7tGjxnhJ1pMPMBDsfxQ9oV/+bMATi
ZN8f8573/76QxWOm3ChvgFm6TiCPdRhsiqnMmwjgrimWzV/dRp/WBqV/IyT5IiPpMBBxhkgB/4qt
J/ogPiFc4Y9n6NaeQiUx/Htmf31XPMsIgZHGShecb+FxGRrwTCk2YOhXphqBePYxY+WYhH28pekq
xthtXHXDhuf/p5yFWzYaWvE9fi14qRJD9IYqIZfIj7VLI0Px7YOeVZYWM4Y9tKqQxy9GxvPMn+QQ
C6PS8ABkdMxIRYOWkDmLs+J/vNeS5k0iXseFg7QMpyeNVkbzGAYUbB/jSJ9+KIJhbMm+G8S8eCv3
gVyRTuCIlxQjIHtc8wv6Zock9Ma24ClLnsj4RV4X9bQJXc7UdiXVzjbgLKohajgtkkkIIWW7V2Ep
adP2dkF4doyQWYo12ruQ5eeDe777Li1gFDNxjqc8gBcw7mgj1LmFUaIMvCk65/gJGgMkiOMzUFuY
ey0fsfnt721gLoOFcb+rBPCXOn9PxJDV4rHinBpfLY83Dnhcc9wjnU4T7LYmdZKchwaZB3GSqWEl
MOQRPCr6hsoQTqPBPs/51jvWnpvgcjLTIq0HnWQkVqvWsfH1tWM8mIJhHQCnOosJcQ293Hgv8tv6
cA+1Iq88gzORekW6cd+6D/ea8aZz2J8JN9HWwz21SpYmS7raBRjUy4a8C0WrNwOM39dLgRaImYPY
DgRxRrCzXm5BAsss4oD60jWWQbQjLqR+jEXEio4/GOIausJMlLtQGvwqlwVHOn6Lty3ZC76pJaTP
Ylu8qJ7QlGPL05iQupCOY35nv+NgJlomIJom9rBXEf0elp7/pDyEnC/6NcdHuIkT1xjiiByOPRlI
3fJr0g10/UT4Oe1bp3tC9P4n9YaYVU20bxpLKpiKdK6zVfmrsBpxjJZYozGY7bWNvvq6997YTw8a
qkp14C1xhKhHm9uNtzYGtnSBH/6H6DGmp4YN3ESw3AFNxujwm6d6K9dDpvpfWuRvHlc0zyDSGzy9
UIM8Tre/bkM6Cob6GIOZf3eRDfucqOYwpKwKXdns1e/wtB0mhAdB8dhhNYLd/f8ugLRf8et9r6DH
r6iGFtZhcC16pGbLyMgs3naIw9zYsm9unRlM+0uYMgdZKxZGcBIqpyd1b5rsqPKv805pRErecHZJ
k8R2hqytq/B90RmumTbzxrbqx0dlaV6QmFFb1zALL2+L9uh5FiRIcE31JDoxR9SrgnwwxeE5brdF
F199UPEN6i2DizOo89/pVMa6U8fftdQshWTdmGb33KEa2uq9XsFNF1700d5f2xQRTTIMWusWu4yz
KdeKV26bREocg/EVWKLh6WWDpB9gzZBDlyvGSjqAY6ZA2/OkKR5vldHT/gUhx8xErHrKG0fQ/Q3Z
DPJhVKgLEsGzKgRx150BOjTv4Ct5yL+hmNcAsaH3dh6KObzsn5+ayzhd6qA/murxsEaZXXxvfzyK
sj7uk7itburiBTsNXbdzyco5/gwN2Jzw5QGfdSRCNbfyrkwdyAZfWDZJZe8SWmEK+szWlAnE8Vvx
mIQfnPl1vmVbhx9FsV+0O56CdkBBBLYxPfDTUK8E0DgtQhDrspVlu+1IWLqt2fVRffMtS5m3jE6G
6gnqs486c0EsbYzIaHZvbQSiOFCBiJ3OCdERv2UaT7zK1xEdw0a50nDtG364fX0j+ACwWCaAkGz3
nJQqnZ5ufxmaZd/pWmEnug4IxyholODo5cQpm6L3aRyhpS8oboBL8lWXpZZIT02alYZ5LY57jTxK
4NjslzvmUe8aiFDqddqwpTTPh5d4mZaD4v4oxv4oLtHAv/ysB0M6vkMdZ6Bv6oKwKbEDynn4bOu1
EczHuM2odlbpIsOVDYA2OxwN9EnQrIl1NB1ezSoDB6LiPfueOnPB9MnD2hEx3jKbdX9c5i9znBk9
NuwE8o+u9NCasOQdVmBxyZNJbKZ9H9+ZN3IndrUnTjByPiS9XB9EVWc97Rrx3HenGAoo/awck0jz
txt+idUaQY8Qg3RyY1XvbrCxzakgfUnwEBwWKnJ8NLS/9q/cUEBa2mFbEM6P8jyKPshVMdZY/Lm3
blR5UtADHZLvGxjnq9655jvj33ReU+tqGeaSAvOTNfznqCK5y09LUjUiLokbn7zWEDjgWChsCSW0
13cGuKIz1QL7IRFZh+4J3oOITWyh21G1EiZ3Bb+TAe9aaiSaFf4Uu6JW2gbNGgPLC6lQjel1un2f
iuMNsnOUC6LyeT1Xny4B108M0TnCtskTProuIy5MwVWP89GPQCROrboJap9nH8Jx4ELsqMpAbMEV
6zgHT7iCm+2jqb6hNh5a5zwje/Ed0dY2YiK6BF+8nKpl0zTzDiQ1FZeAtTbvIa3an0aiD9iicDmA
IXlmi/omar0UWmiMk8hFb/dl5WlhN0cVXPqpKKOcGau2GaYh1L5DI5Tw4UT6Z2OxGlWYqVnnZHCO
iMGdc3UCTJ57n1kA+POMGBS92Sdh95O3oTKjEeuMyqceU4WbXAvHl676idUQbdCo6Di3x5HoGv3h
Y4kus4rej7ppD8UN9aYEQxQyTLpSh4tuMV+9VQ8vCBlyHVL33KzWsloPvvbCnP6nPC8y3mxAcnZD
2LOWDjS1zmfMUiK9T+6wAWZa4EhdxZabw6cT1JeIZbelAGhwbyksIy4GyY5QzLCS4Cxxj55xBTzV
zzBZAFEqrhTi0QLjmyORqz75fOWWiAYgZ3ePg9N2WqzrlsXhyTb6Qker82+ILPyrK5Lms+eM0mbf
t/JDsRQJnXLBin83iobekV/ZDddTlxQdoV5ES8HM7Vssz8a8GtY36ygScruCuLjiFAIaX0Nm7b7y
SUXDqTVm+zQVcEqxpEQUxhJ3smNDrS8fV5tPUVjoo+gIIGiW2G43KVgFT0ASL5uUAoSCHOkJ5nZO
BSTjLAmO1X8NaEakjOMXkaWRZE2NfF7J2ccUhu07L+y3PA5iLn2/vSInUonaByH+1r2i226qnFyc
ug7TlWIDO5uWH0IQrGh5E1AHgU3m52ABSeAAA48f9h9G9Zzty6HtjWPu4hgslnUL6QzFJm908r+Y
oqSqGaKNKN+VTIbetufFERojBhxq+NBepWprVjbFep1TBHnk/AruuFXfRgAcedRzMdfgnwMbU1tV
nJnEHoSsuHQ7/dL32g7KNUMMctGMJs5y85+KOjcMmSyh+RvfkxiHLAzP/8UamLZzonD9u1ogYiAv
VZEGmzzK8rFB2iEShH0g/eYySXii5W2nPMW8atGmKXclS2B7yEOSQYOYmj+n3yyJHo8uhvWZD7ih
d7XAuCnDtTrj3ggpBA6BewbLLE5UcHtkfigGBQUylu4LHxjRQ3+ETIIVnnFGkIe4wLCPLdtviv1f
3sfRWilioJfXHv5eiTLfbJrpp/8EyP81dP2zWwQIjaRhTOq5CWvCuTcNV+JZoMal6rpwuF546Q2o
4iOYpcdNiDez6K4IjRtZ8wS5e1TqxtA/YM0IZgrW9yJD7PTkrAm1G9X4GyeuRHOdcWpnrb4lGWFj
kOX2WSs3FK1FiqHXEAPeTOqINvR93vzzn2xcHOSGeprZ/uu9Jjs5MOlaNPhDh9PityUTTTJ5sjYz
O2V+QiOmHH+W9yea3ml+4NRsnW3yCWhXJfL/dE8pkEfR6DBZy2fq9fONgw9gtbe5hp8QyGKdem/u
YPkRZVw4jXuknFHLbTkh3bvhUAHyT1gMwkRm6yK9oyoY+iriY0Xb9dzojTI3kmidTxBPkp/lhCTu
PHFlCcDiIbi7V46FK9dP8VwunKHxEJ6M46cCxi3KGMeTtTeO3t7bAcbunuER3j9dQz6QHNDOYMYu
nzpaLvQI8Nm9Hau383kGaHxC3kYWLxKjoUjgLDQJJGAefuBu+ldd435rbGCOW5219gQ5/szdNiEJ
MWM6zj9HYiR3w9ZUUq24/DDVxoUxO14TsS+dn6HLHYCkHL9y37kXSR2IF8uILOB1UA3fkDKEXbiR
glLy3v2VFbq8OJjwlMHIsHJInMtna/SL2/e6T+DNHa5VSWhHSPe+o+G1/SSA/Rox34lMZmlKaHJl
Lf8oj8dgQ+Dyp0rIfuoEzYspx5MkQO5F8v86rQL9GmQCSDyJb3sG6d7wY+HhOkeRHBgNkEVTo1U1
tF1xpJ6S0tbnTmTuhChD2EPomrCi+J0RjSKXud5rvPrGp0Iu4p6fXkDvm7aVbVy6qtvfx30C56vD
MKdPgIFJvCIgUdJVE3/cRw==
`protect end_protected
