`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
gM/mn+bG/XkHEwIqSUryWKz4U4Q1pIEsj/RomspninCcpB8084X0HLUfzXz7uT6UP3g35H565ilC
x3J2ua8P9qo8ci4MGtXMID5FwgyL7P+sX4ZaQy2dztDzCnqmgDvQx+OVkZc6OF+R1dBA9o10yXuN
7HpexHh9ozZC82EUVIbfI2CQACwAP8fqy+Wvg9xo0JSSpl19rAMePdajXlHmalbcVu7DYYFXB1RZ
0y5UKav+qKKVaw0vEEGAGD9jw1HTQ+g6WTMqFKoeudaeGnr6k281FUQE03tB2GRyfD1EWZrpgfUS
F1eGqYJMEPWK0jNtzT9HfBY1VFx/AO1LSppK0A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="PWyGfOUYr4AcY1AAC0QKW9vPx3OBd4K5mMORsIqjjzc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 183456)
`protect data_block
O0E4tGQOqtp1wGpqI+zF+TVYnePYuDMRfJE5Akx618w7yVfGJqaNEEC0oBM6NTqpzU4t8aCQyAe5
VwWd4blfO/rrLxUdUE43QBjZ87Xu8uKdwFpWEA6yMGc/4A+z4rAcUPcmCjcHCCDcHPG3DQhs3oLe
Pyr1Xr3+Pp+DpFmQp1e0tlHmcECaM2j9feMNd34GXDHzSskBwkyPFatMkMbAChyjAplY19Ljepu9
IGmwj1BX1VjnpDfcw4eykq7f1WkXaGFuCQoPbfDsQWVrZAytDszPXXFR7Y9HXOPxL//FaEO2ED6v
8YQfsPLaWdy/l30flGIcjn3szh9zuma/1wae16uzbERuDonErq0g4D3vBHBPqNvSnyxBeMdHRFtp
KVSZ6Ufus6B3ssll/tMEiB5jsGyO2N/gCxWQ75zD3H122Lnz6FTlsjma0sjpErBi51ZTWhf2iuGH
liwev5hQygrU2R0QdjTXtpcpFMjLNWOfo+0W7Th22de82TwDg4u1EKLYTy/N9PDHOY+7rovAbXp8
LAOoJ81C90PytCiJKmu7efK6BN/AhhxS6rbJfodetiYFBHKoXldA8keYnxCFal/TFR56vTV7/59k
r/MrzEse212Ji5nKY4uF9CnDf0jjX0ttRSUotzz/klYdHDTyfpjFIhDSZWEKZSj+6sfQuWOefG5v
MLNBIlkM9woVbYNNJ7p2tmykyI1Avk3YfBDlZvk4aYzMsDDAttbdTiXTZdsbm4fTy2EJa34080Dj
elWuxLoeqvLUQOKRsP0cfc+Y7F+lBLQWbUv3SRffyXBDsbzQWBoSK98AxdMWatAMauDodKJ9C+DL
afZEJ4DNkS4oZgIlRTfW21ySUK8nB/W5N9rc2TrtmBih4ccDowVpYFEwcqdoMIu8Xpwe6JU/wIT1
G0QARukWLavasts4G9Z/Ou3VzE0U1ZBTHGMOfd13rtSSryK+NmpsDMFiDXjDCYm6hc9M8pViEo42
krvbHiN9bLSqVlAy4ALF8ptqg9uMGqjzcmslm1Orr6mkZYyr3RWRCzXRSC3jnJEPeLCSmxrqkQ6H
oITdvxSveEdRQIeq/XBoneyD/7JgJKEDP7wtXqGKOR5UqQRehp/ifu+RlOWoLczu1YtrcpHCbzgl
/+o5w4ia3DQ6xEhgp6y+l9QJjOvupLy2Yceinj//FCDbnSVuwfS0yCzFh+dEaobaR6z6pmsPejIw
+MbU4hgI6razwQIPeN9XL90SKD/xKamPSqH3EiQi+Kugb02PUemaRq5reN63igo9X/cVBH31f4wi
SlN58/S1DucLIHM2xsBv1V88B4WuUGgR16X1ysxR6jtpmzDqUR8DZ+rRQXc4XSZmiVsLlzrq7Qm0
+YKw4Xw7/A/SSeqrT47WC46RTRip+D/aUhpwB/vVAzMxm2wjFznylKk10R1bkfnJ1/esK/jbWbWu
pd9UqXbqN7T1m9CghcTRVQ78mexr6jlWk0u7WXL5dFNmo3/EHvoibLGWM3nQXIbcTrGRQc6hhrZU
RAEts/Q5DjDP3eOvg3Nv0m9gFmlII4CIpfIhiPtzqkCMGuJmEUSmLWvBBPiMLmkrm+w4xu3DtPRN
2KC3EH2A9e8B7lqIOYPG29p2ZGJdb2n4PLcqYpO/WqdRJB4si57TBn3K5dH2IGDUM3DVOjxBwkH/
c+IdPpScpcTfkGy7F66tOfzV3ilWdqXAO5LowOC1TBIzfidul3fPEGjlTHhnZt9Zzwr3aB/Btvd0
vtnoK1lQ8BKXq+m4fY5dYAvIqvbcstdEdA+ii3e7AdQBchCAhnrnQB+pQK5V9u38rMKTz4qv3MJ+
36rl5xxfGoGI8XtDSDsec+15NlfSA0ChKZGAAfzRUl6JOM3yWdEVQwZJXwuBxy/zylhc57IvJGiZ
1f6Tak8dSm/q+WPJ7Pj/YAn4tVqsivCk5+LT/XTzYr+cKDFA127IQBsUYu/QMVXKqKQKgERyoVP+
5TsjVCQbVJMCfK//EBzzsNjpVnr2xNF7DE68Kzm0lUQlhg1pKkJxVQR5uPqu4KsShmiOcHwALOzF
AiO53C1jnZinb6k0OjLEU4+ciVP/urdiWavgCgj4VDlwr/awttJyKFJ88a7De/WXSJ/Eiroiip+B
Qa0R3yRH1gjevufSqiTrpXC5B8XmFDL9I6311lHqVJ9QKe+AejGifO6vMgYpQegvRpvZCwwHKQ3B
PL4R6sfafV8eY1uuVmrgVZKxadWL1YpvdqoxOOAMaq9SADOWLEOx2Jz3HBqn8XE/85KhbceArFuv
y7KNxXqCbpG1NLkfrvckk7QSmfaaA3Vi0Hq+QdPVDd5NmK4Y1PhJdsFIy9wRbBGbgEDRCmDina0y
Zw3a+TjFiFBKCSTgt9QqU7k5ZcWOjNSs1A/zT4ygryBg9BI8IQsN/0DGkxEZvEfXvRmwBPg5rP1V
VEc5q/+CjKtPYjzxWv85tH2x/hHW9zUOcNvj8z2wZe6zajN9fMWzIQ5sLtr42fX4R1sDWhzB0ZS6
fQnGRksZIiOJe2uX6DQvu+vomoHG4xv8i4Xk3sDFVFRUeRmFqv0uc/pBOLN3GBcbormAUBFYyO/v
i9VFrspURpG8WdTl24ViAVtgRKCfW9QmRZeBXyuX+2i13+bfsMVDT+NRCgL/GBrxAxsHeGi53RxG
YlBo4YKK7jyzoFpSSWfAcCp7SCY1oXtUJN9BBlKS9EFN+H8q+uJPqvsvDP5IAnKl+bKHvcy10kZ0
ZxTYbZCbmH/YswOnPdJ/EF0XcKy9p+Ck6gsY2Gh8y6uReAUijG2gjKXKZRQTI9S3CIqqzfISNZJR
tIvD6uN0ZUKFrFGYBsuHvmASGyq44AjCT6/xGWfa/0HyZwfDEPJc2qOQs59CMi3SYlPGzoaXRKSm
eQRgjs0qzhmhsb9P9cGv4R5dXuCjH2vChDT62mPW/LZLLtnq71dxWIkU5r7LVBZtt2+Ju3sC/2Io
sZBe1hmXcToUJiFGFdCoEbBxOGgYSXdpZNUnn/O/5NKcRE2QxkI0iopAoxr4QrVor8sdyQLV4vA8
WRyLahnCKCIvgDLoXh5VVkQIuPxLBtW3xM2fVutLt3rqWVkmKeFMjR9jq66DDPq6nIUF6tEtdSyV
wDGsMRM5DiKJ/kMOLCYzynx0/ExShsgMOCorYki2yJXbX/iQOuY8u9/nih0UqsuAXJCsaurQVhsC
wyLz4mVbAf3ICcJhRmn9tY9gDUbs5VHQC+gzqnmFVkuTiY4Ifh/5EuIJAvAwZ5vSAYAUzr3bhCM6
hMOW+b1GyuITgi1dUUHznqkivd8cApHLYQCedqRMd0GsHxACjWmaUgROc5uj02Qqsebv8CzjTt90
d0u72+VtTcbh1fImEe8tZvDJEllNHfK6znLmA9vwxv/nekAy5nup8sQKWHuqtUF4tjrZXkBerdZV
XaTEuuiReWhzW26xIbyFjYzI5FSRx+ra3vBhDFdAA6AYocea4ptNtelDU7xdRZfpw0QYr6JT7SzT
dq0of7ikyodN/YUSJtmVMQBfDKu3gyirOwOUlGfADN8JkbXjeaHtR+CORy1cdidRgVd0JFV/H3PN
X4dyW+3YRxbRbKUWLAgjIe6f2l3KUZDpmlCafDMGA4Gh0uNX/mtwSQvjSfRnNMJI2qYe3AjcjQRs
ZzeiapYKTioALElVFxkOrANL0eIr1frkfWM2WGdgvs44J8uCOkfZS6Uc8SAcxgJdGOl2jNAzWFCe
6I6O6mtr8xhaI4A28GCVqI9hhgx2Fd7ywy7GXrSoybqhesl2Of2LYPaVNY+Za+pN9jDeGicjCqqa
GXNZZWRKZJdz9DgGCzZ/5JAqUjph2ZaeWU5Fm+1a5lcAqSW9jv3fvtDtSPUqyhmh5PEOn61SOlHq
CumlX+Y6Muif33hXOU+aC556BOGWH5T59ENGymRVvBoBtkYIqOjLUAx7anshMUliirQxIeJLhluq
B1gzc4fzuP4TZVOxGbfpUgK8jKZQmPTgVUrm2zK3A2Ozm7PZA1/bQlBlvkw6wYUlysfFOTeAPAyT
tuR1RRfRdFtaeX0LDkW1aHjw3z3t8Ig9sbNnjI01zatCbHBdr9hOLWsV973OrO8fvGZXeMrYaivL
fBb8K0LzHyWI9LrZVhZKcZWRgf1UNTJGOfHEhdrGydOIetInZtmBcHu27+QSwlNf1SQZzx8V+q5w
hxiTChhwOIVh8ZwKwYg0N4RpNubbvgIuW3AxEPl88hS5qrs35fB3BsbeSBRYeJ0KmkIEOBIhZGyc
W5oLlUB80Xoxax4qqa4lkMBeEU9CMKalrnzcly/0da/SsVt0je8T6APNOGkO6tWlCMq9bcwaDquD
dc7O4O9f4tuTpNCM9uLAUP7vc97w3XmMMduwSMiKLaUBaQB/G9sXHNa2ezydMvu067pfWE4YVSwF
eZ7xCLEGz/DHBgR6Flw9214gCRLcccYBdzMZGLkAxYiFxo3LK6SFnpfDHsQdoRbdk8sv1b2kmEjL
L9O9QiwOcnSvxNMyNgR2a7jwAw9gcDoHBi9gwq8hkw4wM9fdphrrcghLkFWg3W+yXMgKgD3P22dq
AClFkOzpOVf9hPEZ30j6IRHjuvylDNKBaxbm5qqkT/pdWEvzgnIHNni7D7kwycchg5KjLaoeqMD+
nZg3HJh7aL/WhDXlAH+EgH07jtXkLWqfN4Pn2bVvV+0DF1jSt0bdf2IP2ASWatg+mDvON3EgUcau
rgNGzna+StGyDgaa7cEnoh7U48ZeRnPsymGZi/esG36bqWN56dSIg3E7aa0G0n6O6gdfe5rGKK/D
8BkNYb+qHzmtFFbPAwwKE5ZgsUUrSfvHFZPg08vphzW/tTVOEjvqDu6O3mFsOQeRcSOcTb8NqEfd
PWjac9ZYuk2M0crsDUgSJawlm2sK9k72s2kPEFblmh51pKIwjR76m0Mt/9v2kA7mjb+F1/ulvl6A
BZPhPV+q06NXtKP1Icou7/vFyFGgA4O4lCc4AK0iPfAw0BmtlC1zhPlwU53rjHCPcUOG/j9MQHms
gn1F6SIpr1cr5pgj/0rrw/4cmU+fGU+cBuPTQwYMs+uHgRg3PKN1CeBMmgPvv9Q7Cp69XURhqWkA
+VGIOp+8H5zE7GmoqcCFcBwHwqcM9PaneO83DGxFe0RlWVJT4rnTVN1tGFfjZqxlS5GVJgPMs+Tg
I1ZogSuJi3nU3yfp77UAuufSc1fiPl3nZaXVgFdATeQ+myCtQTJDSWlCUL8XDfTYmMBYf2PvLIK6
KmIHN2vLGihuwxCFHI2jgESDKOK8HfsagOnuMJvE0XKQhMNPyhlI4qxyN8aok/KeRwMiIEw8Y9SC
IF7kPqUAoUrm9kkSPU/yO8DpwIBkXZD2YsJbytBtC/O3NvF3SdWsb2D5S1BpvqOBJNuyjrdEVKWz
jtyjkMAYIPgPytcQ/gfA50R5Q1WI8dycd/v3NPrJBa73ZJeuzb+vTtPbIojMSRpBCvSZjaSvU+ih
71E3Oj0fQMr7ouDDP03e2Y2JHYt1ix9XK1vLQ0zvpmkSbWqK5e1fh+KAzDbRIcXZq9QfiNKnetat
/rjfHJqN029KyRiU12+RsEV6YEuN9GvW52R2X6H1WzyQDnYRpoFWbnUpgkb9hcbh6wbKg95ryrTH
m1tCJPstzYyJkhkaDK5OvTlkgTzS6D8VFdOLS2jIsQHhHWdT1iBSEKJH2M/8foS5RRc9vVbSpLOc
SVd+0Zb1YM4FTHUI8llNQY2H0TLeg1QpwKeR/m0YMP1Hs82TjzVxHNLdZ0CZxO09/V8Uq9k3qfD+
avkJ/LYfnC20rSqzM/DyhZHu2e324XhN9X1QQxgePg06gZbutoZcN3xVp961gDsbIFCr9x1MUGIV
Jb583uuU9fOJPK+5/CDPtGsm8nu0jo9MbeT0gjswc52wXerX9whE53XNhie+JM7AffB7auSZ/6Ax
5i81DAJo18qpwjn1zxTuo1Vk1kmlsKjwExV31vHlTRqSptu8Z5Yk5c1N9rO95ZtQkzmkhH7uMsCj
hFbgjuIVpit8NaZd4mJKWweYnCSUTEvVra3OWZnHsBV4qL6OwzLnSpAJMY+IYbnes5ZahPtiM+VL
kjQ6ArSTc+Z0XYVxf4Fij+6il63Q5FxMr+Iwg8t2QparBDQVjuQTe/OkFj3hsHbMd0MFk68VS19g
p25O8p9qotYAZr/S7DQ+qNX8951sAGOCBPbkwLN7kauX8GyI4ImY6nAD7IvAHSYUvOIN4DToI+0e
43u1B9VFJkMq28NXCi3ZlyCZwKkOrzHPEExgH2eQEGb1bXL+6/DwqAs76LMDSHJN+a/711ouKeEB
+0wZnQsvtVC5sTbJCQfR/anMYVyGS6gJRuOI8NOQowt85HXee2TQjh5qTJYy3FGxmdaop6d6rhDB
lMI6FM7kn1MKBzrLGXsM4WdI7RnDpbZ8+ve3OPYs4VRrDrgedyWW8JZhQOImaRRFDJoV8MsqgdvM
cFAmeYJ0jxyYqWDcn3eofQsTucdQhZYnVLGH52BJhNp20DJJbFxJ2qaEXbpku1Ud6b2sFh1B4K7b
vPlUpH94o598QyhBLxXRoKpYi4nBZ96LURcfAVj9wVm6WJU9C60sU2QnwxZqExXm5K8shzB/XJWt
ggb+E/vHvzfwEMRyuv0rsy8ptnf8yUTMo17FIJ/XYnqVWglWOTZmgQveeVSQVDvjTJk1BqjqbH5E
bm2MoVXRAHxpkj5445+MijsM+xxrnsj2ht2RuSUpp5WHxzs+jh6gH11giFdVAbmU2ZWbma1Ky2SE
hjXhpTVbGAWR1Fl5gZIotqLlUHVbErn2AoGlPjA8hsYs9jaN5pbXSzIzQ/3sntd43bLhChrfMHao
/hdNinUZGHlsds38MRB9BqbTKwdKkKdBLKjy/Kp7PqH4fL5JVRv8UHpufnwk6xu3Oe9yunnFi36p
eooONImXpcsaFpJqToeBILmrfjITP3bJB2vYK9QHhbkUVaeBudq55nOaiBrSHSIgMQk0P0sXoyVc
QZ0arq9b0TIUDBSWjR0VTF0L02NJuYlmGGpZhNZvxu/TdhbNTZoTxRLSUN0aOIDR6JFIh4o8Jrjo
GN09fr/LhzsJeUJOxe31Ksjli+Xk8Gq2J/9buU2HpD8TFyfaFnTfoPUfdwI25FXk8b5jVzCnGMc2
FEcDB5ifVGTPfSRInR0LRKstnpO3SbtXwJEacTwnYPBItFcV0f/44VbtByrMqNaR4HCRn5vkDLf6
YRg7VcuaOKDFspdjiHZQaXBC0cQrltfYCwi2EZROtPXCA1liaIAISpXcGE/DsmyTt9XrrYr9GYiH
N2nb+eUprDPnMDKW1bKrJMrTQ2Ti8PVmnQQ2iqxPr/4bujusK/ZFy/9bMVMS2aenJ+jw9fnvzoYJ
BqidKYpjzPAwJlgy3em/dibD3Gfr5lKSlKlzEL0GGV+mWYop1uQAxc64nAAix5RwDT3/6uMyMb/E
bu81UeTgGvmU76XTNLa2tExFI3cXMy2kwGneuinq+paUpb611ncmLfnaQkwnb1E+xy/MhTiuNm8Z
7ma/u3ULxWIDKAieBk0IeFQiD9cXhtYUw806HqPR6/8XWKDk80eYPBGKhZ4yQLud89+Mi/7IKOzz
YEY5WxdQyWrjs2v/w6cX7HXCwRpKpolvRE+MixRXkAPoFWsPjCez3OC/7q4EZAKEWWM1IY4viF59
99y+KWT9lPpNFKKc2WIGKr8075EYG+xg69JhL5+/WvIY/llmYS/5eOgJVLUTOIdEaQEjrmpTQwQ5
o1neJuWv7B21NksjrrW5f1PA/4VznmLH667lYYBcxKSAY+eyk+L/fkD15LrFzI50cffKcLydjn0j
pZqyWybMSFzi87A+VxPwqYPAl1T3LGwUiZCybRU0/nd9vkmc9l3Ja4MtqL2aqT4nCARc7qWdyJo3
LkSek6oYBNJSqFV8D3iL2m/7x2O4lQ4bSN3goe4cFWMRhe7M6gR0kpyNEaP/dpqci092/LI7jJ3p
RwgT577kzjD+QVt1fiP3ORtXeRymFaye0IUG+cDHTrfhKqU2+bmzZmBMXZvirErSBmEOY2f3hstg
jDMMudgDdtwhN/fgyrSJIcf6hptvIb/5m6R5DPuqXH5mpoOT35QsceSXVhGYLjqZyVEkv8DegPO3
cMDy0qX55aii6LE8Ych9HQmdl2FyCpiJZpjkEw9xookVI1NQM7YULZNikDkm2JtZdKkM8L9aEBo0
AaxhDBeRAEtrpsXFFw3NWKX6zOBTQsIZaSPGFCKSaUen9lviM5eIHGP/XW49qWRvwUEaswZySOCL
z7xY/PZxkEPXBcQyOTmXhP32DHVcKxHuBrZgNCz65Y43IMIJ3mYMMVUk2JYJCIgjV+2NE/y9SK4y
VBDFXbVwydJ2/ZgSqJ/gUrhhkACu2CX+nJ8ixVzT9j1S756l6D+gtI/ffhXXIQNQEb3HGWMLpGL5
f+cvAL2515pNRFmuabndUrDh0j9iRLVMqnLl5rTpCQb0HT6222U8YdytUPy1mhCxxZEug1usXFqn
j9kMIcxqu/iRAGPD3cLoJ3RK6rvWeLd2dKIJPTmxE5JPBmGe+LCmFCVv5N8X+XzRIkOeIANJFZt0
EkOcurigr402CKqdiH6c8eeNL+NeGZncmLEOHYG+COgj3lrYfJfpujbsmyVbYH/MUj3X2To39BZG
DfC9eoOIVg8PlTIcmWgDA/jmidUJ/P+6HrPIswPUn5e1mMeRI6YxmFVnl7CbSRKyFUaXuLLuMuFU
AQA3TcuhnOqygedA08F+XUEQaSd385XTxGw3oBmw2Lzr9QGHbeqB7TFgr+BiCTBmL4b93BXMX5xZ
AOZX1XNTrrISaJgtTR64otapikK6zN9yQuYSrKL2QC8EIsfzmEdu4xzJijll0KOeT/Rcf6AjUnMU
0jBNXmSE+XZy+S0FFBjU7HJMbZMCTrbov+IUDfY83uSHEDVXwMnKbYUThA6LUpnegGFZobV2sIgB
1e4+BoiK2GEW1PiRGW+s1c1e0TBEYf8v3j9vIkSiOongsAkNMXgdHnwRXLGREQwkq0ibuWjSySMx
37qCFSyaInqZtuACCA4fpWlx6EqaBzla0kV7JW4QJxH1k8R6jVKmC4ZQggadoqydL6nhvnO2YaoQ
Y/gWNNvn9SPSPrumVOU/DaYy/zproeMstyFx9fZLQYVj1pg10RYyRwHD2CGnwgJVtDOuLcm1RT5y
ibYA7ADUWZdvNde8zlyyCJVyW3No/M+ijsf/TiMm+6iPti5BJ5Pr5FEM4NtstjDGkyH7wJAaljQd
a54MeBt94/zRoI8C4c1akBkezsGF+jvHihH5caJaEYCHqLT3vR6+Y9CApHLN8UVJGqtj6euNmlYz
3nt1KBCWDdrAWsWpJvqLFAXogyOgdMeact6+xVzWS/76tyf6I9cRCBaQQeCSkAOHlux399NpZX57
BPF18tVmcxaBPFzplVYW4/RBQNRSSGohbaaQBarPxxMlau4/+WF1KHk4EN9LAcdJCydtAAi28NAI
lRlabBdsF+ZML8dAXYZzgpzom62KP5kS4eh5swm12iBdz+JEe0bcFBPxWSPD/EjD0IFX9WqmCR/W
Ux7a9ghU+dVavd++WstwLoxO3WkHI+yGp/BcsD/o38SVIXzct3RylIoAjXgDwMeGn5c1kIF8Mteq
8JV8WdowtyksPynZLjDpGSERzjpV4/4FBDzBDapuCf9PN1oD73eP216G3cvGJodvI+6CYz+3f1q+
cK2hQrKr17W8WkjU5y6nWpY7PpKPqICX5yBntYbqYNoQM3QoSHiH4P23lKcDbuh5QIh9x8UBprZX
W3NlO11rE4UgIgNmTEhrA+XvkXQK5ckeBo9BDzFer3J7N04KcHZmYJNRjDa1nlXV9T734LCrgmQt
lwVkZUM/yPIsgHHcLzrTPNvpXQTLlh6pekZ4JtfIIOgFTK97L2G4acwF8XPjkkDKi8nBCPDAs2dc
+iLrEj582wfiqaBbHEPR+Y+ApZm6/jCKC+HJnsrcxqDpLA9kZBTbBszc+QvmqnkcYmND3hVgD7lB
ytM/6uSUwb6hlFXzC8yrPe8eQ0/CNMWn1LuF1DX9Xio2TDltLfcq35ZmIWpOh7yaqplO9oR9UjwW
9PFUbLc9ShEhgYM0X+YlLcksFiRAVxzlLWsuATjkSiHL3M3Ze/mnCydBbN5QM2ZRy+RGYO0CqJSt
EBnmUumLullbESPIFc0/sjKX7liY808WBChyU448a9kVTvhLq0tgsSDrtwjqwMN2jmmFrYAlhfDO
reE9QAVjFe7ubMDGt+T86Bo9piQIJPQwsVMY1hZM2vIyJWovnqZ+Iac+Rv29/wEerQiR4j6hNuBN
Co6jOaR+8t+RguKlzGROiLgLFIcgisLn9aIqF/YbUXD/051oA41bLGv103EWvbGYCYVpNPAlH3+Y
dJaHS+HOJlTu26fZzpfxzzxBmiYPglV2eztP4ReYYaLR2DNrQa7X9gGP1mPWvYq7dZWCkUn6CfoE
nURvJ2PTRjgIPne2Aw6gK3q9FUU/TY/F2v5LgmR/F7CDedtgG5LGRVhOGcRS0I5SifUVMzqYw5dl
qyXd2cdg0bYWWd+VpA6MdF9vu7HQilnoTjRZBpvC8GFdIS/0VZibjQJNR05/PhV0Bsa3iLWso14W
RZQtmIyw+yfWQo+phccwUsS2lDXiOnSJr6fVrUaOwfK3cIf0S1Wvpt9J2TzH7meNGj93YIGc0RoK
9rHifdE5fT5BAYNU4bbu+oVQEEeQZz1H1cjKKkvAeJ8HgqxzIkyrOUUlx8d0+EqQ6X/rr6Nu3nY0
Vh0XXTwf3GN+iemOSq2xOXd4f+Gm2er0jX3/OReVX8gApsXBot2EG2/fUHdNLaS3MVhiOC5+wFDD
HrCZLToaQgby5YqhktAdsWGAlVG9kmxXqnh/oJFuth2iaMmVW2A34ANwiDCfccJ2OajO/1XOI/9O
w5JLuoq+//ZdTMaSkH1DRciQfZYKjGOwL2jhAR9K6372PnpEIPiIr7ZIRLn4pYWKQ17EJCEMnc/g
4FVHOBzo7Bicg0kdVQEHJntWWAO1SOMMn8XOO8f1XMpkBiGVijAtsN0FK4vhkvhTgrPPvJViTA/W
0KDN9MPLKLsCvJ1IkxOzQC7ObQYZtws8rVGsLsWD4/dYKE41rnfDX85lEOlHes9FMc98xm+mFPfm
q7y7rBxMrIzLcY26wHaG9L3/mGzvwH5n9wVSnbDdX+b3MKXD9Y1PjzZbxsHNNd2HktiIKSmVF5CM
HLUX8NIs7qOfcfjJLY6Z5h66K4AJ9O4WkGT4Qc03KGceaNHWm5LsK/aAft3X5W58kL0AZAdnpej0
iFiRREKwANnrM2RSvy58lHR5rsoV3OMATX42xjKMAvrfr9RNDqpoVgYecuxpDGkFT2gKVz/3FbEL
Xg0LOHKxds3k0CVbKxnEbIANpcbYcZIVNhER7JJq3aDfnqIIIIy/0m+ZpYwx8usXnFS+KbFN/dzF
xIYJE75uU5Fcp+5r8dZ9+Uj7n36bjwSfcirU19v1E5cU77f9CuV+NZaL3YRd4ehwoKCGC7PwMwW6
AEYqtEOljzkJa+1JCXYE69CxVcb9RBXRs0cQuvdB/7qM5e0ZZw60is09UANlWKQuRN/zk8SbRbpy
yaP5eHZ2cg4HWwdtHieGeSL55YovRKc2CBG8c6+N7qP1qQ6ckXBwtriUHcNHm3vJSA+0t0BH1YzT
ymzDqU8Ds1wEFoNMZrmBvuXAhLgWAmw0CLoBDjYBcOJIcWgKl+fB6ZYWa67WyZE4ZFOP88swwqap
URzj8OVGsdayZkt9YuurysdpDNfhO7J3aeeEw3x4D735HYcgK3IzNTQJOKjOrkDW1nItX2eEP7xY
M37Vl7A0VLGM45a2Wc0eyG5k+tdf7xNzUCMwHN7T2Qeou9we97n0T6WjuKx8SXZfk423hcxKU6Zp
xo7+NiLsd/lJ58103+URT9EoXIPbh6NDxWnbaCf2dIKEwaXQH9WEUu94xdbuoBDk+gclhrXcaoYJ
y/6V9iR0SFDTQf7SOj+8efNGUSq2EmLs2ldpizItJY6Wo2IpbSgZOxexr5oOC6eygJcb/QsPfbVF
3ntJpoxXDvkmE15hegdk89P4nUlrsDiI5OBLSsimOregsG71kDWBX6d11ZgnQ8F9jKMLBivIB3hD
eYSaF+UuiKhCEoLRPAdIRxtZR8vzJ0yoayJFfr++LLIer3Yr0YqStGmKllMSlOBBJnZzLDzdU8nx
5jr/jaGfrjLQdUQD9kIj07b9Yi9m/j5HZCu5aA2rEdU1BXxMSIIf8cQtoQlBb6ub0gyKUcaE9c4E
O7oglFrb6yYFeJDdrIP504EZJPn20/P2Qj3tNdEx/0CfznsvGqvaJqu80ttZBy6pc83EZGd/ztFk
Nc2gVMoNEc++VQbgEBRNemPrxOTll0/hwTIXPTQMk2CmNBjv4YhxNjms9PhFRLwNY2yHiG8i1Jrn
+0lUErjVD2H/PVIBbWVTc/Bajz626jrzKQ4/U9JQI4GWVtLWUDxvhrTRT4AlkpVAfD8e3hR284ur
5LNYKd28agVrKfL4KgtUn6WlWKYkQ7z9pJ+8tSUagXcID7WKejLWyIVu8lQVS10HiRVU5BjagBb0
A9NUGJ5wnsKFPwOBASnbys5ZtsJFUZsFba9XGot+mgBmdGVerWjgt2nwkcdrYByza0WBA1vQ6pnZ
G0GlE9AGg5drC55YtSBffVE9wLsd72uYCsoGrvXZcnhGDukh46D90DXNLcwC0nyrfE7Fs0qaD6uB
1Yszf1sN4uQolOr5yAGTrUQiFGKAlTZsI5fnYTcrOM+DIdboi9kINwCIN+RzNp2aN+eM12+OBfsv
kiqCFOiQX6ic1mCTnSLFoFBWfUMwWauubaplItooKkRujySDLDX+CCjjV4RwtBRFAzsV5qR4Tp/P
utbiUNsUbhr1hWkJGm80cTuhsxpDoXMHZL5jUf6OHkwqIpj1U4QV+wYiF+0ck1KnGN/vouNUzl3o
K5J9OSUdJwphMH3hBgYa+LdC3dFD1n/2/cKhdjZDGu8cVWKJmmuz5hwNmD/9hwyKycZxB0SaVU5R
cBX97g06Un8Euplg42uQrDbYinTHbZKVWFzaP6BMRCNcSZhwcEyeFk7tj3v8/tvqS58VUFsUdOLB
BnQoqOOWWK0UUfevdtoIfWEPmZXqhs/HFumTkxXE24zVzPuqKzxWAKRNgwL1PllnKYWp61C/08WH
uIIO9MdSAcjt7qXmZVrxk0S+nC4BXmEXeFYUWIJrA8i34WzmOfSFhX4enq73cfYE/U9FdfTljE3+
PeyAqWNj1BUZyjrXPsmH4o+kl/mf5qMGPBaN9wSr8zawCZOBdMftIn6B812I89uTCylNBaNJKJyh
XxrCLjvbVonUjhSFahj+ulEsbjmNYAs8gI7AFP5dLrsV4n2oirmubFsbmP4330pWw1h/fp01LqXW
FtYuLGHueEeHbnVeRrDRhdJuObZZbQnRgktiAwTQ40C3B2GojJ/2HM9i0yo/XQNgB6sGQ8yK5EAe
71LeLuwOvw86Ewg2cmiOwkAsoTq+yaBANVQPaRu1CrEe1kUAZyhLs7Mz/UQA6vLLfTV7Ccg3gmNN
x/qzPC6iRHWbB7jBSgGnIPvOR9iim9aBs4LzUfvisUzIHls0ES9vG9d65v41Ij6z9IR9jbMaiMCX
6NKkgDMvvW+vzBxhv4JComkZ0rSpBxlqefWQPs+U/xIgR21EE035jiyU84yt/jDAT8PdJ1pAMth1
3ZbU3iBdgAwW3B0hB7TIxfuNIJDKzs1HNEh1B91jSpSqVCU7r8DDvtc2mS4+1LC/OuUy0oNR/rX8
xO9BOzT5v/ctPac8TSm3Z+U+H755F4COLa0hrCqjCF8JS6QnKdQo/DdeSMQdPNurgHTARdAVBwVM
nnUI5LtJ6DqMGxPOTM6QUpJFFoG44xmS9J9Jk3bU6MeMnhWJCobbXSDMchwWyR4q79/Ts0iSlKf+
nh1ec9nVrhucDzGpDgg7U8oIFqKrmrmKJ9Fmca3UHJzaNtV4quwMm0P7xJzmJ6+xTWsj8Fi4HUN0
wt0Soqc/E6yY4nYadBz8zDY2RwdoiwMVghy6w1BUld6HrPdMrdygI21Yn1GsR6rTDtnF+pWA6tME
sUN4fGhjlYDLKsHz8ScGapb4rp6rIQUA17Rqo/7qa3TJ6+bCgawk6cm4JD6ERzhZEWwaJELAR8s1
+a/TF/7uDXZB9i9iEU1IfFXFPB7bPrSgKG+gWheulGh5TkFsEN6pqK40wC+RPB4XfrV7BsF4+yGU
u2E3kAKwxSg8m4wQdnZXJ4MyCPYl3poXJF6us4ivUYyonRwxRZ3NLmzi2j+KH5w+/NHQa/rWeBN1
TJYRmB28BoYbpTBQMhhELMeB1D3EPoNh/eivFjjTMF+kMS01ZLlmj7Yw8ogHi8omIb6kWVSeoDWO
ETNp7HJoH22z8b3eFN0POhm6HHpLf7P5/qhCNOWExdTQwLCzutYxvNZdVLvYzkGAAGh+MVat8zgP
oQGPQcB2U2MmkO2q8SRCnTnLBJ3bR5Dvr42ynYwu3QfCvNuAM+qMFIL9+YtmOnMCtxuXjJCZiDTt
QSsgadBzj5q6d8KyrX3kaVLQiF/c1wqO7leLfMAg2UPk5ovgm5cDrJvrpy6YnFEzxenUwHUqHn1z
+vHLT4gr7btZmbgrlcekwab1LhgLhbv4PQFQ226vWWU5IPrXarS4IRt6oyxV1nTkvLo+T0oVcuzx
LYcZUkbuzISz0IjNl6bYsRo4ZMWbu8Qizdp0t6TbBuO7fqhG9vBcbgYttSoeQpAk5g7QwtpXubf3
uFr7dTfSlsESgsKfFxGXBCjELZ6D4sEY/qgE3QUvEUg/VKWeVeTxgO6a59pjabSj2/D0qXQKaBdN
HrOSPhOiL0MoTwlOqFgiDEKbKpSOgMqsSnMUKEcSGe5h3+SgVKY4luePuA2FPvEelkIw8JaokpPj
eqy8Ro1zzEOjoyWrjFc/LleLX5/m98bv/RjCpS0t3h5Q594GbV4rVVzAw3C2bp8gd9qp0Y5bz3c2
q7l5dI91df0/PdYVoXozLTQAEkV5+EOFwJ5mWK6hOm+XIg4/tCQ8GzkJ5HV65iZk9qrwKpU2Srw6
An4HXPc1/NuDM6QkFx+jxlpDIu6j44YaQ9hXqiitrr40KbEmZHXoMMe6nU+vZZ+aocQh/9PifXvX
PDRegzIM4PepZukLaGEiw5H9/6HIk2sRdJhI09XqWYaCVM/+vRz6ALbnDL+7iOIEx38RI/GRWTqT
VC78CDlZ3Ptp776AdCG1wnqWErD864Hc0CcDVfbw13oKBmihw5xslEwb5YuUrN1DA5bmuadDxgzH
kU3tnVgos8gvyVWmwNX92AaC1FTpsOGNkJ8MblzkXF7GM7ONLoaAtDdpGwveCtB7wpWxf/HMMqZF
2ZBEH//m2yWjqVF494PaAviFYLRoENUt297q0tNQ//42oPMA04pBOMd6+gDislWH44UtEzZRuSvL
3cpi4ppLjEMOKicRnTaD0Pop9vlw2aaWTvsP3OdGaufe0fFLSlYqVQG0hcgOvtmeEmepPkWmyC1L
sAi7QLbJatTBbc+LoyXRHMggUhnacj6DKRt+syOnFe54PKZ2oelA2xMf/+B6BQf/YQCYjOC/X+Bj
w4wzzgMbkqkfzCdMZQfvkPm/dFUvboxLIuoVnQO8q5kLiQxTqbUa1xGH9e95aAk/N92XaWNir5h1
lc/e+CNwD33Cpnfci/asrYzb8Nje65aQ8ZyMtpRnHR616deq5rznyLfTF5NX6AaRP8etCWelOiP/
zD/xaZzq942039SwBYQ/rCxgH0yQa70ZcaGg7u7L8IIypnqxU38bYWbmB58HtF2yDdz7cgcs2uw1
rkj8NrqX8UjGcnpPeGTdQaiT3QwVmeOQsm5HE26bsuRrqejkdHLjkgwji/5rJtbutVWTDEQHF0+u
IKiKj+6tqjeU0JplBK9tGp/OHCjaQRiYxgXSZnrB0Na7TTATdZusfiBqW949dGjCPbuKYjTVfGg9
mcnlW5v97Eb6D44id/QviZpKwsEuwWQ1eM4tjB5URMTjr5hABwRiNBUDJfZ4RWzlVx/aWWQU9J8i
dG3KxhFzjdY2WHxxYHrLKNSV9avSb9jP9sLMZK1rtwjDlVZBPYd1MZ+wPWmcWjDawjG/yFNCnCwv
VK8mq+mDt8ei2GNLFl3nOkLSyoqknSMJBuTl0795en5dRzyH9xMS2Mq7rSSAfTdOLJYXMJbADGXL
vKaqOjyeVdOL1p0vX0vncErPGF6EmPbbJ9yv/Nh5noloYYpjxIQcPWNQhbTBEl2msV8JJHCcXiOm
7H3c5Oxuv/ArbKlWkF7b6P9Dm/mmbXzDeqluasL8AUDeo1+Dd6j891TCLytc/M8lgNeSkSXnBEjK
a8pYmLx7e6J1mahCFcwV1sfIhF2iXrvUUA1D8GN/cybz28y1z48kRP+GxcleAfeFuujVsDBlbwox
hMFenHmUJxgnWlNQQaAfpvBK1TVBwsuWANAO/d737+Y5+pgAq6+tYijyt3Ln7GZ16bq9OZyG1kYk
4JUqcSnApLzNPpyECtEeuQoLbEP7fUwjlHlnm85jC5A6ULqKjC1Qn5R/4H/ak7TgbMJ9Qvo6Q6NT
6GXqTQRwMrScTBNZmKNSBsEi0lLQ1vsKblmwdsdn9GIBm7d3PLbDyktjAC/iP6LzPi+v3z4O+Hz8
hqoazYBL1VcArAiMti1Kxl6DgfhNLMmWZ9VO+HDCOM97RkTfWEXnniHzxZCx8kek+Pqq/D9hLDyV
CCoXNsP9jKiuwzujKJVg8FlPxNDsc6tkE8N40yumj2VyligF2/Lbv5Ud1EMU9TIeSVWrdxFvxwqN
AcVShPIDsIZQn8/x4a6GKs3l1uZR4IYDHhCwy3ERYKfqI341+o/hUh6Ydr6y6JhS6qGQlPnVcAty
go86J2ZOQENqY1HzuuTsPOaCk5Qv1ADY/N5gmCKqZRIgeNQqYxv5hEAuOk5drOEODJrLREecSdjt
y5zEnyW2uF4zz+7hYLd5CrBlWVKQGAL5M2n9/oQfuRv/FKvgQ3sLr3xZRH7Y9ZGkuj+NoD987mm/
nWV8g2ArHcramTWEnGRReANyBjayJi/5+7Ot/6jRlOm/zBuFbKePxsUS+6Gi+xV3ijS9KrHWlPSd
CrGwI8nfQnvEGTJHF4QALPwM7FHqX4Nnun5QLnXIOk42vV9K2BHqVm0TK608ARMUGHiUFZ6KO8lR
obade9WbttpWQOt62vzaTgOZDpZoXWLSItwfLRlTanbSQH2UwqNHLdV2GSCy2wACi+flISlJlXJp
Y4a++fR7sxyXnrTAq5VWK5ilVfRh83Yr9h3kjy8NF8n4QUdsxG0TQaDV9xD8EmnOi8EmvmhISdU0
uTvIUIpEz042ITlZbAZCKCpTCVIDs+mf8dV1IJsZ4tOpU4vJkHh9MWmKc3F11iYZ8TGU4WP5e2zw
2iqCzIU1YyY9McvvmzXkGGb1RPBFGcaRsIf8udZLTMZB4B0b53Q4XMZomx2CYS5kic5bLp5LJBdp
KV+hy+irbpwIQyIpg4uQukA2orTf+79pKVJKlFai9YQtp5DndsdQlAaIUsnLuYuoazkvhBPRCs9L
MRxWqrhN3nfrklnk/0Ouy3zVLL2p2t8yoh6/HAChSSoeG+PBEsQuSEpeK+8s7tfi8hgRWbZPM0BA
hBroXzV55gzTPbdvB8phKWGV2jp6abZoyWLQyxo8UziZdK/S3br11CJovkcr+TiZUH8ZWftcSY1F
Kk3jdBLPDnDkpOZcPp+TIwqmTD+4JXlABRZ2gaD0xW2F84uBnHoHR6YEotR6ltXggspM37UZ2hvf
C5jqdSIfXIzl0prSmtYJt9P7JVy2cY9Q2I8soSBawWMkZkHzfuIBbkcu/zAVN+rTmmYguf76Y5Mb
7kuuRCAV6D7foQS12z3QWBmcJyPVbs7cuSzk4Gwy4/nLJPHgbwUT+hSBrCCTJRz45Lc+g4rbvay4
lwf0hrgzwXoY2iOiyPAsTCiXcSFv8VVp9XrBt2e/AAEkV4Yp4sBiUsAfiOK7RYquJ9071I9P8na5
pB/RNBl/wawBeEF/EEqk52lQ+Qi5hw6NTsW6SXNvU56GlloWfAdPUjpC/lZoer/L8nJeeOZiRlR2
kFzBwkApYGxKpAms2q4kftcHDfx/a2TZ5rpaGcNCnyY5YD7vR+ICU6kWttcJrkRkctOb5N5sMPQb
+mLc45wPpxHGnlO7NhXUHqtIl50oGMfEu7Rh+PRoKBbIynjPRTk9PmjfnoA2LGmOH/AMzHQowqd4
MNS1s2SYjKmt+Gav6xCSbEQmDkuL/MN/8hU636eNm+dWTnNxIguFjuNUregVGJD4kUyK+mD5n6Db
QK8o3vqOZxnHUjbXYGzED2iD9pvLGl8F4xdVxaQMsZqVa/nnayop7P2lnwiU9cZ19UeCThDH3V6v
YtMZJSYG2f9zgPmMcnlR6+udSuEd4vRBN+b1YR5baIu4K58NK9zLhQcyz+y2i6slyGGusBEBzTdG
ddz7IjSYlFQEUiup/J1xxP7As384ytKZtDrgfVHRIhz3VOc98ofA4jBIShNdPSeGu31W2QlSF2xT
hnM5CxqvuAK5HfCTvC7ByNRC3viY+OMN7IiDOlPYF5tXyFz+7x2IlEVCJU9oMN+RIUGOFZ/sU7sk
cjko9fcvzmdgG7Loo3zqIfnUfCcDwy5hdk3PP3Cg6LE3waVh1Ju76ySkJICaiXiUEfmyENeAfnRH
nDnCfsH7IfFZAkMxYXJ+chbbiCRHYqsIl9cy6ifKDW/gbVf7ee/d25QBFpWweFeqBJqXKPtfWlcz
nOjIHTxyoKp3mspWvvcgHSq8umt55XijTW/UikWVK7Q/SVOxtHgnSgU8w1/FLG8I8CVSU3h8sQvz
lYGT2YHoW1F1L70CsJI9HY1hz8wHMylFMwR41rXD2nIYzziKWi2uZlVMMbsRy1035CcjfKnfbCCI
xWxi9MaO0cRlUbkVJkZ/sjmkigK0xiWyHQReq7C/7xSILjZl2en2B/p2cqUtP8hj2qJWo4mReNpG
R6YlF7tugrhY0MhCw/XFVC+d2t9Kbk2aE8pMk46BxFvjM3XTT6RS/vZn+VTQ/5jo/xCGO4gMJajQ
pgOwoJzNw+DeZYUC3K1bU72X3NrTTU9hnVbBh7ek1LIpED+dtoqqhJKIi0QFzOzqREkDhnxGWRfs
QqwmwPQp4qlS6c1yfaemr58fdhT1epwjMXw1s4RS3jB5LO7xlp9bLtcVDR9RRY+E/0G8oQUHRx00
K80LLPn7/us6UD7wA9jnG9utMdHUsoGRrkSadXmPR6PJz2QKVXqFALARLuuAdp+H/nAftHtaM5f2
nyCwTonWjUDE5rqmlQCzGcYDRuIhNM6YhoSA49HvgTYVcdu1j3T+SzeFbtMe5dwje5mAIZsrN8q4
cmWU2YoZX3ArtJAB3PlOn9y2L+lB+A+pQlWpsHt7VIrh7GicRo18fPr4tWtrS7PEDbUeNFx5agiu
QpQXkqKecvMeuUzJixhApThAvZOqre773H2hoIB4Trn9AXXDdT/1EKgjxj3/Hk6DeOfR4apZFLZX
WYvCpMtrP3JJxw89E2ISgASO7FLqUr9I9G0h4WpyuDmpjjWNXgfkhzP5pUCkWoYahOhx+JXFTaiD
i0Q71BVYXqyaLtwjH2q/9TN/ruFFyFFIBAfA9tHZ2C/PGSbXe0Q/EV4vVxZnasISFv5+SUlpDn8N
v14Cw+6RcH9LSUJM11s782zRZp2yYFEX5Z8ezCrOSUu5AVrgP27uBFjS/l5vVhgym9hClgIL+NB6
kIEnJwu0vSDcvs8ZDj8cHJySICqT81GZSSa5Mx1AA+OYaTN4lo7Uh841pwJhlm2BKjQ1Sl3vM1fM
ndaTEA1QCEiwByqRYwTI7SojLW5uPQOjMJn6E4677kxmydcFzw3YrtxuT+shLmr51zax1li9XQf0
FKyAT4y0JHftuceMEfc/6FfPkWRGuvaT8tT05wJ0Ujej0EMIIPGT6xE8/3v0OvLX1yjDxjrTN3ym
z9gu9iSDHUhinyNhSGCPPJLfEMXHTt5tw8OfOrnAQ7RKLFznlhmJFQsnnHi3TMuKxufrDLLN99oK
1u8kV7fFWQv/SvPJ/TClNUNM23CWT/IlH5OGffZKP8QNYR2RFGVxTIt/ngaZbjPuMgV7fV2K9ycT
QWD0L0M6n7N9zwOwnjegiQKT8JmxuG/ZWhLTKlAL/DBRYxfqXGjiqgIh56+dN4N19kFABmGsHZco
a/55/SMnBmXbc/Gnu0SKXbyyjcSAWQJriJA99BFB/gnBPc9KjnepGH2c6pCUa5arpZ/gNvIkO428
3Dn7cW01gGGDAAQBLQ8hPCEjxtrtqesTvB1nODYkbMF1h4DBgtwbrltExD1rX+TcRzjz06c2AP4u
2/POddrGr6hQpGz2OyE97ag95erxs86k7JnPSWn2JbAPZXpKSLEp+KZiVC+FjOZLQhZdIyajoZxW
wQkKIXq4+I8yXeaILsHzE36FxIBi6yw5cexW2fX4dqTgwJAbrEFkGXNcSb/EfA0OIjRqd20lvIC3
G5fZoQVFVtx0NBapWIAfuDLCXxKZ27p1aEboY/Dt7TBcfrWmxV4LNNf4zs1GHLx7rBL13znPdiIY
eaEyRbFDceKxHWD58JvkjmMa98OBFiFL2soD8lL12nd3/f2gbNW1FwzbWamc7uElaqIX2CNX8ir2
j4w8C3Sdmq9RtjcEjpl3nRdVTdugmvFEXSSPs29wi2IW9a1U0xsBtBav6WMVh3HZL2JUKocBPYNA
6Kdizc2QDevQj1ylr9pb0+nBNTbvwQ/XjHCUf4MltfvNyQWtFroxHb0KU7IX+YCu6JILizuCrtZz
P3sLJnjvny3l5Elk+R3fvGajZmEOYeEjxBOSwMmO42+mg8gbTmGR8Pkk16mye94/xdzcMTUighSm
4sUFMVH4H4Ky/JjM49URe8aAd8oXnlZPcgqbm3EOCAcpviunp54+WiS5jSXJkxC7rTixmbEwJeJ2
xUS1/vRj4dj7Mn0q69KTNh9mbTQAhiisbTaZAycOYIV1Dorbdm7NkNsUiMP++q+epeZhcc6Kx6m6
n7fzd4vyBwh57jp7amodyptl37vEdNjN4m1z7ATl6Wp6iG3ZWioO8qCoPhKfuXf8tC23tZcTGD+4
pP2HCZhkV6Yr8Wl4pg64f5JW4e0PHhbcQyx2uAvjaNsMIfUVWrVo2Zh/bN3udtzGiCNLG5mScGuJ
2Ew5RkhmR5iCMqySFIpAxOiY8qqNiO7xSMS+yaDc6PAmEbjjECxgUWl84RYLRkz7ns8sRRMt4Qwg
px1zoAiDdijFouHwpbdByr+yo+PPFoYgiVyfwicDzdghk9jGoq4OLjfYuZFsu49EEg4hxp6FwNbZ
+F0YtAffiRpNpWiouaFPVhDmg1i4scS27DLBie4avQzK7A5RBcOL+rbA2eAS2x3yEIHbxvkLU2mm
w+FRQxDjNGUXE5mGsmJelFeYu0/coVcXEUvktBPtXkqsyVSJSYj4u1m2jtN1D5moRhauX96pwbyV
Du2DljgDlDKrSMf0pX/JJyeoj3NEufKCVrsnvaNP+6eHxtnZ3X3pB+YKQ3SQroKDWqHDWUk7IQWi
w5x21fmjJsRJSy9jEbTX9vclUXP9mSsT5w8g0sOQ54F3dLUuBrsA20O7fI2gGbOssXBV9unOjQ73
vsYB59qCcrBJGSRMl41mCvQv7HmV3fk8TSr/5kqkKMzZpMOFrHiNdoQ5gJAW+GmKGDRMzzzZAGFA
pEwIaQdQFrUO4O97imuchGOvnmAtjDsgMuC2lG0ZoifAykZJ5RiomQGLutNJuL/3hmvQZweGOTq9
xYXy+n7eIqiEXYSchfIl4m5pw38QrkAe+CqIycBtjUoRNKiWiabifFE3cq5RUZlu3IcLr+x6Jlty
pzXWdkg8dhNwbO3d67rm+1si0xYMGPP5CzNszq/MTMgqGuXzVNsphWcGBM6FkU1mgynUZvJkyRiN
8UbHMidV+NuDcwzfnLU6U6NyQGUJHcebo8tvQ4JZ3vgrj0iRMe7Wp7OhMtxSVAOpoo5zcV0oOyi1
MQbrOPb5biDvaqs1zElAzsN+BWo3vm/evTMU7jxNbuMzhyefhJy/BmJ2Zj7Uxh2DksRP4N7j5cZa
K35ToXjJOZ4advhMinY+58kr0F8FWe0yUHlyknopH+CF72HTyzTLKKSGEgV8FYZQUUAOerNk3FzQ
BOoENlcS4LCJ9oSWovtniLiShq6+WKD8ORLQG0KiNKsy3D5fGWK9tpvV0Lm4o+uQ/Z28OTWHvEC6
vTWMtiKsSeLXkk4tHdNBLTD0MXH1Is1K6TmJf+7FG+l1rtyKNlRG8Gl9KmreBsFJ4uNlXpSRqODm
pakfo+ONqbv1DC6F29SvVUYiszRLr0Tm7LguZDjhMIphM0yA+Gp98JhximQVPj7i5Efj1QIVqul5
0C9FgVa2aSBtK5lWREX6SUFxZuUj0/Pyc4UxxkBSJ/tvbL4ydQ+trGvIc7yrQtjmHsx0a3ShcSrS
Jga7CBCAigWgLrb0exzzHGFoHyS8lyoB5OQFjHzu/+3KyEI90o1LJbtZa730BwKRV2yYilKd5IUL
T3dy0+8Meq6Hr0aZl375oadgrN7d/ZveJ4zV05uu2jEBtvC5yL1VW58DvH+zhVQpcLWC/4SZd/eB
cxRIxjmeEI1ykz/G/qI0j7jvSDh9Yu5bm/yvnXWGt+5q3BIiSEWR4vRZusCE/ih7WqgxNhj+8LR5
12Ku/NXNU/LbjV95wz94h2rYtk82giGEtgDJwpuypYLCOnIluzCvRitnPCLtM/veG1FC0qxcw+En
HQRZCVAPDFL+qJjlf6ZlL0VN2dfCGKVGrn3TSfboSULzra9IELNZ+LP4FXjwAhMRoNYlTC1dubzK
+aefJ+mRspI0mHMlTrXNb7GbXoo6f+twJOk/rv5VVjwQtWEwfxHeEsIN+ejdQ35HJJvLHXF9Ytyr
Uma/xuAkZHBSih3fObL5HZwWSAti2ORHXupqjFmeUt+9mSRm9AKLWvn8HdFYoIgR7jmZGXVk86SJ
p2dq3JlJxUeW4zj9wBmt087w8y7w0eqvpeqHTjU7jQHMrvO7kU6jYCxTRs6HLolUlNmGTKZ+6mMy
8Q9xUUU5URT3aeV5AVi6qUZizGSroMs4aJlooe6XyPNGz/eOUEKqU3L2jAdxOE5iwaYcKlc9fKo/
VyWnEUijbPIDYEqhbw8S5/ey7mHPZlmrPYp1mtDR6/78tFWnt1iXCnxoDJW4N7uNDpNOTY+MxAuN
9J+TpmlynWkJDphQW9wTmvpXeCV78hzS4SAtrQLAm6Vi/JvKkdfRF9G0q16WKoejz+f5nC9DRETp
jAzJBxtZ9jfW5hh4Vbnc8SwBLNraSsDqRKFS5lfP3aewHWE9sbPF6cWRnAn6AUA4dL5wcxJC/qrz
pBnOs50ryiYV6L1QahGNl8yOukVVy8IV/1KQbdmuSxrEjpAKI/AdCJ6ArE9QSfHVr6pZClRgZ8jC
Rk0jlHPdpyILIyd8BHcPqIqE0vaXFLnJpqk3QDSIcuimacxDyDqF8+JQUYDb4CW3VjDXQjfgUC3V
ZVdtQi2Es+jediHqw1PXx2K5kFiJhUeCxzC+abY9l3y9W7fGCkAdu/Tnz/6nbEnvR/AJWKMPri6F
dep0TEMxsxViZqobKvUvjJHrGw4+568zUv60wy1L44JoUhINvTw61kZ0owvzAJE+4sJsi+xA2vkn
NRu+vmyAu3icSMBsurXqXZdcSeBoeSkU68pKnZSpDxrIaI4zhGU+X87NO4xImhjhVDWb6JawBTdB
KFIQ4ovrT/Sh4YR7sKVXhvTQicEZh25K82wryqnYRTJSBOB5zs8aaSW7RR/9DHJTTRzUmGt4L+Ss
WsTMmhfRWZ+DWYehEq3a/h3dFwjxVWf5eLyhCxP8IP3pbOIgZynkbty6HJD4fFv5LHeSSQfPQZOl
8mrRmmtz/xntwkDYFji3mAREUZ+7itdOqjTDii0fmZ/j2PeIwGPdKdQ2j3Dhd81kFjjMOvffqau7
E/jMYOO8zhXnB+sP6BVPfeznns4bx6TUj9ozG046QRaWoB+rt7eBl0JesY1ZfoPT04Wm0E0mYosQ
0GZxkrfLzCqKk4v8CPhYp4/X4RMzZxwXLOoyhsgMuZCGJ5+IinayhUvDcISXSvPRl0MQDjDIoRqS
vO8nGJobbHgxDgWLAZZ1ijo5Ffs366zXTRNmGg3YazxVmwaeIQPw5Ru0ut4XEOf+X6PaocAEEmkF
LnS/qn4Vk79YpArJYPYCkfwYkATiUiyhav/zMC/M9aAz8FZINyp5YRcodUw4Mhd5aU2skitT539Y
8g9/G5Oo1y7PXEkFfGoGw7w8cL+c/0rpWyDzX1lpJmFShBFA308lfcbgTlW4W1HPW5adU69nOuYv
BzXfz8vSubGsrwxnrKmE7NXSgrJ2p7La7BPS5C9BI2nHB4A7D6/pzeOBw/kiR4+3e5nyS/ca2y0j
nfdtzZvbwJyyo9ykYU3bsX1ZgBLQnZKup/54o2hJYPWZhO/vq4gULTsCDZ8JX9Kirpg3GTFHE/BY
I9Bw1tyaKffU1WBFzOwlZtrZeEh1e7N4eznGZLvMNDd7XdnWA2Xa3XOed6qYx20clyVZy9+E1n+4
haKuwL6eXeRuWWTUQMQuhNMRX5Pzoj3uo+BJhgcJjbZy9HQcG5HDNh6Rvvl7e2ZxHPW9bhbHUrnY
SshmpEpNpt6MWLlQsTGKYz7ynR+I94Zea2W39pH/Jp0UC1tYGhgs58ITtU8+xgryegGjdDlZFOnC
p4pBoDZqAOucy9pw3c7XxD288mIga9rvTMzjmkfG+knAh7osootqbhil57IOmPRj8SSB0R7IMqHe
09sr7lqHncotcSrk6SH+GftKlGlSdBX/SEzCdQO1Kaz0X55dK/nBlOUNtyKYFv3YWFeSJzHFdb8Y
/pJXeybUTz7EZkZeIuXcIEq6BecqReE1jvf9p6RQ7a1tmx+4DSRtNvzecg1ya4VeewYx1i+3QAiF
j9yRQRSgc2cC37B4dH//Uxte4/w3cmEsfdKCM0Jl0D4CjV1QJTxQnGoGvADK2WKeG5qVf+WXdBeF
n97bxTCIEtHoSEGg/xkQiGLgY5RZEuEq2hTSrscwyVu3NMDIVMh9BSiZ40bR8QlnTQcxOJShmxXg
OT+yY9hGvrmz31SwnFd3zugf4sW29VI74WalJmplaB8cBPoG1WCeTdsMaoOFXAN/zag3v4gSgMG4
O1drIrRxXj7H3t8cbO45cfm15+O4MyX1ytHU5qg9d3+XMEDRRq5WK4fj1o3Pax/g72xbeKRzkrOv
S3rSy09AgjLx/t6/ZpG+d/ybqh/Yrdgn7NQGm+5ZwjSVarezbnyFtdeHmi5S5h97BBO8SGwYViw3
jlmyTIXTkE52Ax+3cV70bYRUl4DwF8LFmGEno6BJuqNzXUkhZQzmW2zwU92mjnEYEJ7S1l+WKtKf
H5OaI1WLqy1XqLtc00qy/Q/bIfej4dCdwSR7ZzLwTuCqe4WExK2fL8YXqXwIz31OoUdZ8mtOebBF
LqnMo7D/97LsOQeMrhYsUVHEkIYk05AxWr6/bAERlXD4rbZ8QJOk4X8qgQU9nUlepC3+GWmlMV1w
Xe8D0ioFehLWE6mbA5vNsX9kg1kFAZ18KEU8UCbyE6SyBdhyaRozwHhMxrF88McqVwTL+bfxZ01S
lT+htz8656r9pWWtEngCjxVfyFfjRBo6mmZinAL14PFbhoOhz6U+Cc5Y/FffoUkiFHdoQWgxDOLm
FOpntAqfMIDZUf+hzceC64gj2Xndkgh3IVF/oGXUGDhzVRhsm5kSZwmwza3m7uQp0bWhMuEBTPAT
OOxM/i1SuTg/6XlXt2H0RtH4X5vQpjzkCC4tGGbD3ESDxBKlImzoIR1c8o08P4peY2VEVzDB1oJ/
Uujw1TIiTAVCs9SzMenEqXjrbehp6y3pi9YiuUJKH7mjJ0Is/sQloVvsfzguZQDiypk3QhG0Pcw0
U5bBUNkg22VAODJSoS8eRsqaRd4yEiAQk9FxiL4rtSJGoqyH+xuZvQf8FQoMCwjcIo4nKX4sgRG1
KOKkbfl3GATbQUzbfsedl3KQ2bNPSQjfHEYliV5o3nUxQlHK2QI25Ls5FVxXp9pBJhc4Cwi4ModU
23h9eV9ScNCeEKo7Es1e1MQN8R1MfwVR2vWU4zq/riINJpjZA4RSJW/r0i0V8m1599OP3+oMyATp
HL2K6oNi8VIs4vIzcoRxNSY+Qktph5Bdvl+A+R0/kBL7XiiU6anH52+OC5VBzw/F0knjVlgWCPwz
lyJnn//ZtwdOcv4bez0DNEI885/Sz0+UZabR9bZbmnmRx6fouR2lol+EAwnh5YSf7poohV1xu0As
qXmP/UV34LjwI3DiwsS3m1O0hkrnl1++5ewqV83FaQ+W+N/1NkkEtjcQduJG4bcA1lJaWZyPD7V2
CDjpoTPmWnhpW96E+kt85z/FxI2pvTXBCMhPfKFxy1CNGl6fvbBjbRyW6U43CBRj+L3aosQdkB3/
FTzvbSkCJtrF267/nNYU1Xor6uh6nRJoYH9leGMIHN1vHYA3y2p2WQ9pc3NaoEsVD2goQ5osccid
PRMsKkadkfiTKPPtXd31oGHXn6jNrqW/+G9mIi+D7nLvMVtK/V0GWF4dNEi9NW4CBVrnVM+2hy2R
nUeI0a/KLk0RylEfPfQfmBJEUGVVrZWUfRq4Rl7X6jRlSZa1zYnLh+0jIuUOnCQI77w5/vMN7RmD
PmuTHnJJMmp0DXdbgKncMb6za/ZHBtHYRkZdUfGGE4e9XrLlWJFxmSx2TpjU8Y92jAOJRKK/5yxn
R25GXMTA8svpmkZBgT3kXtNMHx6JxVUGit3giSbaKVmB3H7qrVYgQtJ05m+7j2L8SU877VssVudi
+Qt8yNRCyI2UjAK9vyTyZOGCrHEpMTJgGzvxDc8i3k30lmYwt9yisI+Tj6eWPDtQY+/Iy040NlpI
LLmyo13XShSfGzYgryPCU+uclOWDhgHIh5eu8ZCFnPKkl0sgcHsQCzBViaUNCPiqXowM/Vd0BOrz
Hp7Xd72gfyNQN9cp+54Z77d6D9Vnods7KGzUm9s7h56aKXu7KM+fh8s4a4+Xj650QcFQ5XlBE5P0
Xle+1EKGSicsFQrUSDhyy2PvDFhWQuQ74n2hRrbyqgxueRDCkH3/LFkZMd1VwNynGIAJDWTZVjIQ
JGns7rl3bDaAo77pwrq7mwJVvjbfLscD4DKL3ndWej3gZ+KN+Vskjzp9g4zM9lPAk/VHIBUx6gsB
6cMtnTzBiukbd6UzATNYdFImx+FxFrFVi6+ek1ofQpgPIuzZlgIJfn3amBmEs82brsb7s/RXv0sV
TmJBFFRUrHZZe3isdV4OP9HJi4Mq53xlht+pL34b77xw4YUy/G5OKt4CnGeJUMT+ci7N1hkfJUoK
lEzgpwXZeHXyfUpJJnVGhtc51gZa4teseg86jPUf1+tKcdymdY2ZoNQaKvqETAmnbRpYtMMF96D/
1dV+MP5xzyvtPK0aNm/NI9vGwIkPUCK+IlHjtQxfL3Oc0qTXJtGEB1u/DTMIxwQiref3dxRZe/Tm
A66bMHjGCaVEoQuZNza0Qb8gmLpDRcjrDlG0tIvN2rJ/66A/LGWLm9chIQOfBnY2akl2n4FKJ4fi
sBdZ3tSD8XtyOKsHX8FUbIzTNZy+BF5qla98GBIybU9oHcdBZ3IFETr8H96tLc64j6dbaUkbT/qZ
3T2wABHUrgdFjw2fd9g6FPPJ4Tecrr6xwf7HWq1S9OZoKs/EUNZPHD6Vwj5lN2xNuPzt97T/C5HX
ejph4wEP6789dplzPM4F9MC0xYhEAB9yDuMANxbzdOvuDtiT16kJzOSvxxvavqz/xRPrQF0GqJIs
mVNtfbnzRWqax8LEEglMkk+4aoIJQFTcxoJafKsPlShzw2aFUXAbYAVTTmeeFz2iBANXojRnu3EJ
SXI3K2gx8ZYH3RwJxopxMwuZce/BslInJGWZ+9/RYphvqTGa8qBhskNsfXTBj2Ivjvd10I809pWK
WZsK971WUd1EDjzFsmvIFlRIopf6nP3QZ/seiQVuQF/JBDNA9WcFic7orHmgp8G5K8HfQ6BVbOXn
Gk6yPm0gNun042BmqFfYgcIE/ftuB6CS0H9/OYO4V2jMDygCSUWyb1pUKjLzz1XIiBlmUKUn4CPI
2Bx1bVyHnIfkX683jxpB556gd8Ub1EeZeblan3hhrf+QCu89HYdozA0CVd4A2JZ/6KtqffWQ9y1P
3ktofsqlMX20gAgfmBueLWhQfE52z441RtyAEMf7wklp2TfCF+djLb/Lgrus90Kf+8DySin8nKJj
7Ak9pOX9bMEpV22MCCy5mXduVAde+bnVYMML2pDt+kxLqBmo/KTHxiTRrzVsU8ww6iT0r1FZe8VF
CQ8x1ZGrii+Y2ee2bcaQdHK6QymFrVW/cMIPbMdMw6757ufeZRMZH1XPns4RqM4Nrt+rOJL7dR5q
jHf6TACuxO2B7F+wfzA/sBSnt1oVtgXgEJ3lhBO968X37hqLq/1nRK36Gw+4vGcKuT+kzowDYvg1
mZJv86gi9BnVaO4PuJwkw53dYhMcN4xe9Z3w/3M71/owKjumc3hA5EsW5hFbRu2x9NaqTHosLxjb
2WwheXYBi4ObZC0c8T9cjeKG8FauM2WIqu2QlVKGm95gD2qngbhkUTwBYq5rjpPmpIzd55f2ODhS
dpNck16xHDUfB7VF77n0MFy5ofWNCL8CPLZuM5RB2XS5aAtILMc44HnZfQjQSVuXxcGJWl4yJ8QH
qGCnC1VcXkN2LLibFmLEGc5eIUEo7OChLzUJuC+TeZxYmA54JnELnIUdFeDb4FlaYbUV3q2s25fi
7ikzmIAwnzBVwgg+QmMY+rh0xGwlwt0ll/AbGy0m21g60II3C05Le+iYPvXG2eXbZgR8AFTzD9S4
o1Pl+ZL+dv+RvpMlN/kkYV7hWxIiiVIMNkhAM5VXNIGEuJAwKTjHv4K//BgmYL+1zEE65lYNN0nU
p9Zbv8EwjSLJFxJ9J2hHWFA8wzBTott6eNYNza8ovmuSFn3Xp8bo8SWH9PWNUoVZWIspxaOZFjAQ
E5Q1foLLkzRA5VoBY1x0oCaktcbk1E6bcZ/LBaB0svfjKFdjrnm6ada6E5jyFJtFtKvK+N4yKmg/
Im/q3yiVwqLVuH4osIwm1MgevLRF+BY3Ow6qVlQt9idwsI7CP5nNF1/CJO23w+9ZtQCapJRyc/3h
UuAhLdoVt2TXs0cVMIQLgY7MNNAj49yLU/6MfJkNsv9E/Dxu+JyfTGQTA4mYrzQa3ZQ6Lca++eOT
uFefElprcLCzMnQ5Xj++nLaCGZ56NI2yHCcdCuOU54ipW2Emjlid3s9YenHY9zRZVd7c26VKebD8
Il0uLIkrz0EGMw7OT641a1zbpOylV6ROyqPQqzXqmbkI2EmCcUP2NzjARIO3GGEYbTorZVEzxZZs
ZO4p3OzvSYYh6czs+AnNcQggw/i2EFbSNcvpcZ+mXphvolXzA4ceT1wHGC45r3pIzan+gS6ok6OK
OFEmKbMuwZu2E8Iwpd8lHeh2oTScIyPhmnECKzt2ezuwzulPa3YbTfDOvRQPR25Fdb7QaIL/aZ6e
h2CnAXK2d682IrltgR4JFbLxiB0xWBW6lcZ7UpaVag+I3gFFt6euVFhlE+sczksKnLnU7NrLXb5T
hSc1GqAZBPe1I7Zoit51yFtlsyq3GNMpFAEs99//Ww0V5fq7j1pf7e8pKPzDrIzu6IAx6XTK98l4
tBPfA6Bgm109Vjl6vTuCBzCZzWjEAnPgaF+HvFheWOc/0A85+WHUpVyytLhVzMTazdzSvP252bVh
EEtDuIrrddc2KEf/eOivh4Vvl1ghBmUYNJqf32x7xYCiq2DuMzc3z8aabXhrJk18N8pu0bJf6IkZ
chRlkiGbAiRyixeeiBRiJd9dkiWl2wxQAObF0ML3ppVZxgDanMVVjvA38N7vflaj0ZO352MpjzKT
1Tykaek57T9FbZUs6QW5WygflExAcubKsDrwyUxGT19b4v10LDTrap/b6cN1WEADy5MaIv1dVp3w
LtYoKDRA+PcTpNStVzsHh9Sx3HF761Ogrv/ZAcmTyoTO3Fovp3QAL9C8ILoS3CTlk/AfqfvQ8eqG
rPcK+z+TIc4NflnfSTN3CrXUIGBIMaQ9hHzuOGKZVIP3cieHVyUTOYez90iHMR0hfJoRQ4rN8IzH
oyEOK8yrZf0QcecwMzEGOK72eN4FelKIfO00xTLhb1NuMGvYFm/CDSbrzF9LtaCV2ZtoW+Ig//ZJ
oKNXGC+deFgpNm/jYb9Dx/NCJCXK4tc+AW7xfSwdcAm+jUT+a2uWQzH3HLi8NOPVv2OQrIRhuvrC
5qHj+5HftqlBcwedwzVGn4KtHZzRyp0aLFGaBbISCy6/1JJxeB5uoETHNHzIz4QLGEzoUTMAnMPx
4s/Xe8dUHWiA0ywmaCD2k84vb91usEFa5LnJSi1tRg6WrTkERORJ1up/U7rr0ew0H7kq68JIKrKu
ecJCDCqHdYSsugRkEUSmF6MWRd7bmzFxsm7EMimORotGVSyFyRg2BDwFgxDAkVSnraOFHIWvKDBe
q5hsjiqnGmbwZO8a8L5LHeoXZmCAuW18mM5ygsvboR4/qGOpIGMIQwETeVeLYJhwPZivp0xo+m4W
c9ZOFRrhdOlWszPcsXAh2VWPo2vHNxxtCS4zlNRwrJPGdmTcv+Fqw7s2Hypv4yvwV6qAEIvOCdar
QG40vXYB/ZceS4CyQH7b5sbr+xK5Fp+IyKDWMJLba+vSSXVcvOQQKKZmaCs/xzAgj+IBSWPq0ulw
O8p6IMGk2bjVomvopBjbI6qm+NR4iJcRqeVeW94zmUrJsm1Bo4MNmjvdJK2jO+zYLJSFZqZFtR6Y
U112Bn+hQMTjEEA08rMYorPXtDVxYsbdOUomxK+RZosBCvKbcg8c/eFdOW693frGVPVJwjRqSuc1
28JBNb7tI2jEeaMl5ugNlI5V93BPBWSiAehAnlTxaRQTaHax13cNhEVXv2e+xvojsVNXux6e9o3b
TZ2K2TqFomX8MkA7XIPgh2mXz3Hg2M8HDXRpjrVduaXQNDrAD9IOJo8+z8yUdtOPyrtquSZevprX
eGcjjEYpuCIw1n2mB5Ly4Hbcf7A+rCq5yFpVi1r6pHn3G7LPdiZZdVvVsroD2Dtx4R2ua0Ys/gYR
lyHyIiAvdszCscgT62pzoBOqwo0Q3BLPEg0TozAXUCyfOPeK50Q4riwXSk99iEDavMBvTrtKZ/xW
Yr2gpy5yXvKTO7/gfQxClBCj4AGbmmukUBy7HiX6AAl+xMauh0vinfwerWtZ4HevNfBft8vJevVo
gEE8MevEBirAf0wbgxH+kHFvyIhbX5zNT3s2w/6HtARLVDM4s9GQnipknBS55YmRVV8/B51BfkJ+
QjhCNEFw5j7IIQSYx2dGIbjZWMeqfzi0OK6bSlyISzeqOgabJo/RAmOMqV66/Pf09qvx1rQgfSzg
JPIMv0d5MLTFBA+JOLgu1+2RSOmo46rtbdJOL94mFqJD5000MNfUxQjUhIw2JuHV2kBiVbtWPAuB
gMQa+EBeLTt5meDMxwjn7pRZiA3XDzmQrXtMLzOfH2fxsTHDq4jrxdYq28Kje1kPVD9+w9Fs2y+y
XiAmc5iU0bxFm63ZSRtH8y9ykjJYnosWpQSLuS9KkTvY8iHswhZT9Oyk8GMSEFajd6DNUZkFqyv8
D5lvuR2xEnFtii120DxjndjqlvHys6mykiLQ+AwnnSLR6zC1kRTq1y4prOR9qMcuO8eSkxYVGAi6
CalsbM03mnFH6IMLg297q1J1VaB4DzMMSAaBi5DiqO2wlwFsZjSgHlxvAsasKKRYqt8XFxSuUaW0
/Fw23vl8s37z2etTWK2rYYpEvxUZwFAweyX5Sxyjc2hzO0Ada022yzp1uV7ki3tjrk2bbOFr+2VE
wY6RYLJAVCfNzV7YOrgGIsM75jR1BNj3qKsX3N8WejeydzFAejDilhmLDblfnBwotk+EE5C7VStr
uyH9TVrU/Tvb16iJPqQfqecjWDO1zB8zswKDvm8N3kAbNdSJYdyNl3kT6MXYrJTD537uwPJ5AYGR
ZYEJ8R7Do33sQ9ffG6xBla5ss+Xo7Q9zBY6WrKVv6NLYuVwj5SF1NNwjoCyrWuHVqA5cbIxG/CK4
xiSZPJEw+qh3fuqB6aLfAyTrKHknjuAbf/uf1ckoGkQMuO8K365Tjdd01G7XEO24jFiWGbC5rndW
Qoy92uLOdKJu+2v0+HHwg3RauUWyAWLEUypPUlgVWvFQCc8CnPMX6K75FJcfMp1683iUR68b94Is
6D7Y60wpXXQKYSb3toilCmjrD+KR3JOLh3/P//qh2OXDsEYbJVJa0rnu/NUyopcKYsXgSG+m7paj
Qi+geju9NWzgIqput3jcG1V3gYcd6N7KRnnFqSNAcq5r84PK/pwmkVLfgPvG5Gg8DKzg5ruapqK1
65fUZyilWtd6jpJpIikWCSyi6rNeVLNy/pdS5pkVwqipocdGVx5Ll5JnRQfZjGVP6VjcjCDOe1b9
CgD8F65Pqy5SbExO9UZnHYT5zpyJAKawFnFR/00e2sZYyW2uPn33xRL7NVR/MNL2tANAL6Pjh0DL
LENEHYj9r3Ac8f60mMraSvsrjBNrly9+2VbvIJlTDWT2+F/IHYYPnEFMeHrMa+eL42VBNaJ+13Uq
uCWnoKf3Ym/CdJ/vYncjLnYCEPUm89eUvZ3J+DpK38mQgGKNbY9TzHm7dy4X07AKZ9Ih9hfsZ4hU
Jh3LJbs3jv/4WNzeTseaFk7XPAyOuYqvzMRvxR4TBn0RQ9qzCDtuJe/XGYtCkppfBZNwdC3Xg/MK
5TmeU99+5XpBgL8bWl9iSXjnHzFuEBbptIr4Uup8b2xrPK0SCQQWJPlkGLgwF/X/RA6S63rkvMdv
k9O6gq973Vp6ET15/gYR0lKQpROJx92cyTE4cDMl+o0i/UgF7RfhcSI2FPhPStLbkz6QdfdjyK1l
1k9uzOWwSg+07/9R6qXakaKQBMeJcF9A4n+LGUuPN93qSR12BdLJCgNeBRsqgVApmfZ/FYZfdFhx
Gi9g69txUXvKeVXrY42OMnRfLEiRXS8hJ7dTaZcu2svuEGHiL0zM6Y2puCsFTlb1S77bYSzf3+9/
d+WaR+6p7fgVNp+td46rACbYqQ2agmBvNQ9dpsVipkTEBHX+3jh/3IUeQrUpWTED8MRcnt33zlMD
nY2vuAEB8Bsax0s81vtQC+W4OcDUTQMvJmSobR7v17zxmpUquae1aVT89zpa9Z6Obdl43oom0l7W
z0zQjgJjUM/v32xmrSiWAfRoAwkTCa+f+7KPPUHecuj6A67QErRCJkX5g18eUuwPdKzALGAbiIjD
4aHGKOgq8wzcgUDc9jJug9l/I8MRU6KO5Um0Icd6puA0JQMOF1EXS/pn4bhQD+bu+GSWcrwSuLVX
V38GI+gI2Xg7ftwcSSbl1jQabXix2H00/PY8pU9I9dfXVxUsKn4paxo3G/a1Ey8GqrlNEcaOW/bf
tdhCF+CRhJ1Tlb7xeLQqjazOvcHsSruIZFlu7lms3FxDq/NyIEnPl7wcEd70IMzPXDEUnzbWCb6g
2pdlo70XAohOlopu8zrFfC791xPKvZqfWhjyPUYukAQKnvmxzoB2EHqDA8soVUR6z+IJtZYdEU2s
g5c2HriR1t2vSdhyk1jRaoYYXRcUWinjTjy79HPW54/WbIBU0ffnsXr7HMpJE+Om46xZtagf2Iq4
yUW0fuE9WKmSHYTymPRC+Uy9GML+Tf0Lsm4rfcMqenve8LAT7d2Mnf2SyW2V+4e7QkZ4O/ePigSQ
CgAVuNXA7KCI2M0AF1KQiDMe3a79591MPQ2nZK3EArwquwJLyUFWUDML/CDfw4eRJzdpnwawocED
Rcs94QNVlX+LIioTzWD2JlH9fv99dKRUv3Rz4lphI4KDuN+6S7S5VH0aYwOfutP4wQ7LBStrjl4e
UjH/KJvXnBxlIQKZs6ZHrZ2U0G0N3WDPy+zyzTn/nv1bgpiFAeeShMplFu14uP3ezNc4325edZCn
pQplO6hMGNWZXBBja9bSobS+M7+MIwk3dJye3AJ6NCegD07YWi2Te+KDeyT2l4WgZtbRIhzZ2TnQ
qqaiONVSLTgMGFqBj0gwMPttRZd/wd0Cn8RlmnoBA6U4/uBPdv+YJuypUh6Xa0N6uMHSgwhr/HbQ
CFZ9ZCBm2ShnkohJfweo8FOR1uOy9w7wV/w0OykznFPmQnuW7emhVQFVwjD1xilL9NltYSAVEAbi
PBvcS3PlLn9Q3G1RzGjqaNNX3oVa+VKG1hpc42/hXY3fOqITyHvYvpTTOMgS18ECsSZXn3zP7iJ4
WqsQDjDLtN6aUaXCy4te8ZwkqWCPQKSHtm1A2pnLtblfTSpQrDHtaA2T7wklKGuW7YwGvwwazKgp
JaivOszqjmRLcrPeqLq2IaTU8mwhW+ekUUqQrSLUDCTm1HcUNcKWb4gkhTXt2ZccTKQAOjwe+qWJ
Cn9QM/PaiB9g4yrOX6+DrTduMxacC7hrJUHFN9sSHdSpKMEVafY4ePbPRSTXIq8dSwARY+rhJUuI
7bHO6OSVP5Rbfir5KzfsbBqk1LQjQG8ZPKwRQwOcBhTfYfOOjYmW/Qq/AdZO/W2BAnPeo2SgUbHS
WEwNZ3Hh1qOgJwlOTDVebDOyPWA2TIh5RnJzS4n4O2TRguOiIeqBwRXHyJjgI2uFb6P0Zn8Hy1/G
+k72DGwOnZ8QZ6Xvn6sSzzVZYF5Du0QHqwY+D2MwlA49pK5eWOY5ptImRBbrXHWU5U7vU+P8r0dh
0WOOEcxgCLDf8tHu2UxQ3PJji4snRIxDnFozCy0BYJve1RGQAhuapdsRB4Liit75DRmDxGhz9XRk
p7tshljnBmXBvbPV+8xRUuZocUhPUbrbsblyZfzvQ5rAe7qPldBkERZsvOvlj3OdWfSVLpiEWdfZ
4BzwohYVJQZyVpeApLOOIlESXe+SikZmsS8PvxfvstGFPnZYAxS6zpSLs9JpYf5T+YLZ3PXU3aKi
PgfJVliaeSMIMjRQMYYEefSno3lgLqTOZoCKQqzWsP349fwaX7nWVjOmibrE8t/u7sD7wMESI5bi
QTgvgxC6clahdVn/pE4BpBctMeA4aIZXKrEbUmSimqsMEMi6Fk6rFWj3KwPfbd5Hk/UsM5gVvqwC
O8E5go3eDj0mJwTB+3znrM0drjnfLXRAA6/qg84HyaLDdCPk6ehx9O/4TeYKU52PYnLsYjRk75xy
OPlu/X6TZScGoPfGT+cMC6O5GQTDNJlCkDDJ+M0nD4t9jY1VIngYgkb2OVe8YqZUT8jhhNplRxEy
uIsJvOtfxD7AAdUZS7XErLQbu+tLgTilfKnmWKLAU4JF8Tg5BDCoIw1f63oH0wOB7Z8WpRFLwsdI
I7iqN0cedAdw3bQq5cB9idB6/NI8FCYC6u+sPk3mLD8Gr1vHCb/jrNRnJEotKdJrRSYrNDqICTMN
jojhkBJztKOI4jHbmO6uEnV9PFfu9UYOhEfksetp2gA1HqLIPRz5X1Afz8FRXvPX/TJhX10CK2Po
CdWycfShrPyovRLCy5aHCmDVLmTK7xpdUDGmxg1WSuU9sNriekwElgqhwg8Yg2vXQxrqFFMmRKkp
2lB4/LqFxnc22iseSp+dku4Fb2Lw2J/Hrzpm5CCdnOtjUsiNBU3FSAhmgdVhlbDbaGBDJH/N9S2j
F8LNKPmAaWcnt3N29oYFkQ0dfVNtNBjNJumG6Pm5SK4I+DdIQiiSad6NZzg9EB4y1a355/HGGURX
o3YeKlPBTpFqSL1OTdEaabRptcX5ZHlHQBb5nvTZe3Toc9uQPd7UklGupVpOzhG2+OrQDt6Q9V6S
i3imHzrodl2K3nFqo3jFeSSUtQS5p3IEK2FP3YIU0mWZ0F8ag8fyD+fRRQh6z8b4mS+CyEYwxSF+
RmajetMZ9NuvFM3BqprALM97qIEzEU8zUePDlP+Y7tBgqCJde9cypfM4skRafBCylRlTnTuKAcHh
n4s9gV1R/8+1X+k7LVm6ju3rPCzSpx0QTjeNYyBf4VpVNWhQ6DhvV6ef5p/JaHbYVChDHG/n/BEV
BspZw9f0VxWd90qKXRmyohQ+Kd3jsdagc8xdDpUcHaU6yRgQt8vJf+5pdhPZKT/9ZkoKEh1QJNtR
PPol3p1AMuJac7/1k69bW16+2PuKK++s6hf8fBYqUheeohaUAEngYPFfYj10+tIkQUgABRs+gW/B
1TyOBBLTwoYSuVdCBbDsGy+S53H0Y9fbmdDn5MqSGu09DY24O+fcQrvyigKD6Kur55T/z7/rh1YX
sGlFSKMAIQyMce9IVkw5/iKt4VXEgCXNScXAbcUVlQJIVKPFJtISP0Tq6SHk/YU8/WJy86GPcvYY
6vBQEA2+/CuWRbtHBBXar6k6+tpgqb+NrN+keY3VzdSAOgx6X1MASRU2+Hx1/EkwtRn3oGvZiW35
1FLPEZZlnxvEJ8ELFsehSR/2097GAARkYv/15QqxJRk67XatUFwOMfC8o0ELKM/hNKjkQQ+cDEj7
1c/RFPG58gBTP2LKcLOML1sqs9tIFa9nwLRTmg+ysORDYQOxSKC9XhcNcr634uKfT+CeYivgLGRJ
lP4Gzb8qhLeldbMQKAmPP7lb5rhUPwTb6N8t8IYrgQ7QTXEmBAehW1v4z6VMvYklVim2yzy4fPt5
krW7HFQvzOuj9ps515h3hZU0qMg6AbtP1tqGmR0yopk2NKvFiKOam4Pd2wt5Mrl2i6gbNdc/tyPx
SPCT2tcSJhVKlIGeJhGxPlovMhf0hQ901rv1IdVOZIl00s4iDSmggvASWuSbECeM25+zD0wbNeHE
6rW5K1anz7rdUlapowpQzoLAMzpap5SusXMcZ0VbVZxV4L9z4k8Rb5B1DDYBg0CYV7q36GIrGsii
6GVCkK/Mfx7M5r7Ucw4ZyoAs5LxsgfavwfAaj+seUW0HQ633mJwIskAK33wIieOJvlzo8XsOxcLt
bBy5gMLXOaxeGJa/2tZH7gfFF59qpJfuxHn27ftrfKHDd28KOmYENBpLLULoWOHXRCmt+0lA+Dtv
uL0uk0Z/+kwoGumSq8QA7Nid8uX0bf2gla+8PSd5N/jXuebcPPdJyPIcLK7LPcsq3teUDMb66Ae0
gu/PdLzVu9yMGwgnOESoRhxifSWRQzDNK6lOcnBM2I1Sfm+75tQEVH8qoFpD0lGy5WkgrdrKd1cR
sVi551pa2w13WdqCfg0K+a13bOlHAFuYdhaTbL0mce+YS17j0ABTUnDj5Sh70eLpUP/RlSKDF53H
kM0yeT1xL7haj1ZXWR3SzJQSXqo8VTDp1I9fZ5v+P5x7bHxj7His3oMlgwg6+9Xzm9xeXPbACWL+
+FTWrYtLi2kKjRlBqJbZN0ATceZEk+deEDGfi+YodymssgQz03j8WPUrqCmpvJFBP4OSOX0X5Aj5
iootHd+5nOnTIRJEJF6Z7cF/gXJXtB2gVi6MPsGF5asMON7ZTYAxxZKFsJkYWvkZYBJCVC3anxPw
H9NN0kDQZ0S579hszXi8G19/2jirMPj3puSkxD/z6io6H0bhU33HpefHv4PSPtczv0z4QTWvk6PW
7UNP3DHydZZDsx8K+niU/6IjHXECYaK8mOKUGcfNtS5iZxqIB4YMf+J8hG2vZgxK4Bo6hkmpaF25
QGOyZNoyEHbaJrru5L2rggRriEb62RK+Wo54MrdnN8oq91NxGN6+HkcY8V7cccXOSWf4/ASA/yqT
vDPBOFs5wR8mgM0poqDefb5dbjcfP7Mpt6Jg/S71jZwhxlxClFuFQPbY7x8cLbdCgStV6HHGzFKY
Upt6WWNoF3n/m6z69jFNE+IpYCmABak3ZyMTnHCOmimuj+9bb0phFmsGzoIFlMwaUpo4OWUaPL/D
n1aA/KBY3VXfv46oJC1WQvjtPu6YcPdcHb9bKI5KYjKIMv+y0mb0E9I91k8DsBJm8gqPrTB70DEG
Q5iM1YBW8twT3ZYQbJrtJmLxpWqO2ddYFvl9wBwZypWhA3H7Rqlrp70TmaoO3IerjQ06TU/GBOVD
eeNZja+Vbw9DVVaBkJYlOUKwvYCtUnxuhFJ2RDRihOM0Q22OUU0FEXln4Z0MqtbwXZD925LywVp4
sTNPC0bsy37PJG4JnkvMddZ7wy7nZmXghN5Cw4b4DDNOAw/Kkkg0ZKEWsZPN3WgqtYa12LcrOnpi
LPG104+CUPJX5d7U7wBiBI1TS98HVkpLcx8Edb9FkBc1/dHQKTtGB4G+z0gDQytP7vMWiH+YknPL
0D7R1Zk8TG05zxm2wCl05WxoZjcjofaWZ7CheQhO/p4IkvrUtsYFpzy5GIAEWJaGImdbS9VqBJGv
+jVKAuDN0xsgx+JbOan8it3V8B8+w9rPw0yD6a3ZFNZ8NUpTLaMRaijZiM+ptBPO13FlxDmt26IY
YuElYQvfP7XLLHEmSRP0EMp47vO+Eq6rZpC1/rrIF4fydjhrhPjlpAcoRGCDes2ZJcopgnfr8TJq
lRiZZPZVeszcEgqq5ilGOk66FlTzKGwauUFwOI6lnwzzqDXs5wFDiTqg7o0s0gTowgx2FN+ixbrZ
V0epraJStL11LnHCbXR0NMe+aIL9FmXrXSsn+52AFnjm6Jks9Emmej34C4c1OLvtENvsR7+1O9Rk
MYCjVEzcmCft5dCXeSn8NThb8qOfW2LOZQp8J7rSNxI9LsVzmrJ3l4+ZZXrkFPKrh1k2oecfqsXO
DwK0j8iiUZ9TDkcXVCn5jRqcBo4SYMQHB0uufSV2ajQH+Y+aeCDQJgB3tYhxdGUchUciaRmYsm1G
TcXe5f2YshtHNf65h7f2/XmQBDt3FVRUov7TihcwvMmWOyiFJwjtxUuuOlo+KvmXXGmqN7CWTCt2
hDgpKRv5PPBPBhb7eZIss1OkN/kiPCL04ssy8jKZ2p0s4Pl8/EDiO/i7yPQJwStRjTSgWodnvaai
WiT9nQE5NU2LdmlrIuWmkhdYBtVJtoUsiuFjPxQKZcnhgS4xQ2+VGhXFNiNUPks9tqxJ6T7ixRWl
riFEAtJrXpGwQTbHiqMKi1cUBN3FvjRy57/Yi6A0h1SgPz1i97WzRbIURmUDvInS6OHEljmNXh16
IvmwS60PmhrABExqXQPol0QlTeB/rht8N6MubWe+cxRIV6xUNzh9HjBOTZAO7dyCvqT0tlya5SLl
TTR4BGM+3jTA/qsiZ/MkwPt+xudbRL1liHvQi/sTlwBDwvCsLpm8OLfO/N2v49bK2StfpUTOoXaC
nrchRmPOTSrZflg7G6nOksyDIK21u0eGjhJGmYPoQrkmYHSUFajf5qGtzFbSiAokhQIURVxRtED3
F5AF3KQngH1MnjgWupEDTfPlUAtAOh7eDjBszIV6J0t+emuO1yEKvVVAOpCkZcPn1BOtAFr/ROr1
kaLGB/40vUorp+oaQujrZOoHxFszcfvV9huOq5Od0Mb5RTPTdIQ1DUzkSRDMp5A75biJaBAV4XLb
RPx4ZMqlUzm58l0N7u6UatXzNkhoJA24+TW8qTuww/5icJV4/T+3a/cnztscpt19y0ZDGfYImBNQ
A0UIm8yXDppJDtINL8XYufQ5eRqky8hpoW//5RhBWF6f+SroBtce9M1w6aD2C7wX1ML50iXzk01W
JP9JSGE2McdcyWqiwrAE6inI6lkAgPXT/axOY0FkVcMs8ftHHn/gwaeeWPr9guEINVgDItmz4Kym
yfceD8gEFJdbXDsYYCZMdzJ1XvBz5wvCCnRo01euHluFJmCEJSxP4v+FSY1gynmzJ33e0yN0UOSF
yncibt9UUoldNNH62xMEuhkC+wnLvB1W3J5DxiPRpGwf7lj1/VuMvkyZ9PMgteo1ZKQSrI3WDKjz
G/hUf2L433qEhp07lJ5Ft3Ej+IYRVr4Sg/hRBwa56nAe0gMbf7tJP1i36bKekBa7HNdHEcwRWuxT
m282ziQRa+OhZsAyV+g2hXC5hOQ8zpZRuHLzt2jA9OpVnKLor596t44OmPgfszbDLiOxrXo+VjTu
4UWBn3LXFmBAXoyc0QLyEs5GeRPJRsQp5lGgMD8337fk4jSkR469C/gxQEjGBklsJshe43jU4dAr
Y8B1EdHtjGvrEtPHFMvn3GsV7jvn5kuIjFDaHYQl1eyLUIkw/EaYBGDf2rRKlJwaaLw277hfDgDy
J5ivwpr74i2cvSNYugfS2z4Onqh2Y4yb36qFYGqmmbdOioGY0WcVEzFc6l/SAyPBHv7N32AxKk93
jHul+C0XcepRIPUAwBhWhS5mWU/rIb4AKrhDWfOy6aRkpninUVo16YKrWCD56QKGkCIcMTneiYec
pA8kNoUMw68Y6VFt85PBFmU/VX0KQnxPbpU8re0un5VehEVX3HU+n25Hdtx6X6F+9n5NrZUYveUb
eRB1/ULBLlM3054XdoWEXgmjAqllAPM+xgmffCHwMSSni2XZfvHNS6A7Mv8reEWI3wMN/QkLec5P
XLICWfEHfuP6xjC1JylPk3s+zDCEtEGubPNFnioFbBa4536PrlHOJK/Ylz3i9ZLuSij69WZHNlV0
eD3KgOnwi/XaBTxLHrjWuRQA+TbGFTJF0ZCvjk2i4GHD0aGdRxR9TxNilqFsjBn2z9Q6gcXoFJFi
5OSp8IXSDIJTM8j0q8tr2lLpMV9mJ/Ej62CZdD/ukPz5odYk0EYDF7jiXOAFJVZpl3HjNB203gmQ
ZPihmSzsyuaCzydME1p/imVCKn+vr7/wHJZFbRr707tper9xY6cDYG7Ta1kWmLvVwgxFV4jRXeZU
VrmZi6muk96uwS1eTsdsknPhS3DKGNkgAJxzqbfXZ4SH8LHjyzeUdW23zrAAeOunYX14Q4slVcM5
Vx6NPFSa2A4cDnkP2zN3R6aS1XxWx+cTPGn7AbtSvYF84rtW4wv207Quv/f1zfRp7nDe56xutN+X
a0VR2uwtBVpjUUApofHHCmHT09Khlvu7twPwxc/yCXGquEvwn1YgbEJwGHm+uEmDrYq0+VH0lyl8
GN5RJpLpygzFBeUXqp6vEou9ffe8VKvwPn1lh0r1RZ8jed1nrc/ueiU6JroF0+PHbQ9e44DGzrLd
G24sDml2Hv+iWyPxspaYzig5GHb1amEfLMqt6E8KADMGrHl6h3al0tOW1OqPUEc1/LKw2efBzOru
J4eiVBpbpZkudR14JlPv6/ev53TMgR7JSY5quKQrErjFFlYbKoMiutiC0qmG2fo8LCDtt4yZOzvV
rlo4Kiyypg+thypGzdwIlXp0Ukgp4Ra5Ght/PyFyrVI6q4527ox8zhfCSdJsLVuo8vprDo4biyx3
Q/TzyO+tpw1RlU7Mu25cirSp4z1LyuNnJWKitCJdZSEsdTOMx7lbWKKibbBj//TuMCpKbPOyPo/G
tjOkOWcNH7jiUZ3vYNy4IzBtk0CdA+5iQW1x+2xQCFagDjFiZeNrA7KxYvABrjrniZ+BfUCAmcTp
u7YbZmdesiLs9RXU2gYLCuEAFNdmhdQ4J3iqE3mU1+SJ3r8QJ9ExjaUwaLW6K1QqfJb7p0yK11Fj
bS0bu08F64v6tbWBVFjdwNRmUANYx6WdaaZNv60aH3PxCMNcB2erNJpzrF7fQ7TFiGhnyA+CCHZz
RMqmlTpBXBmezrqm/PIHLdU4bIPoEkUO4jEfczjwng7XfOkkGJfUJQj/QdlrGeBD9u2q2vLhdjBD
fdrftopJG4CI8KPEL9fpAHDKyklh8KFVVOwK+iyESwAIN31ohGtCjzxc2QIGRbbAs3Byf2cc++L4
HASlRA47zUPXjJKl619+G4g+fm3RXwF0fB5crYfvaq6kNx7bqVcvdIKjHWadPnaK/K8Fmii2OfNa
eNY3RnBZRF3riHHy/R7/iGLaW3kjohgYFVFq/9dK+AqyR1pVgNqPA8qcoAXsTfcEYfjX7QDmyGZZ
fGuIoupyEA73YWgJnpmnZ4aAiRgCSnBv6WL6Jrdo+AN+8TMV6ypiiUGuTv+LGq1huOesjHNhoV5k
Q5y+t9KeKDIKjYhndfWgXj5W9AUR/0DGMBPT9872PmyeEoE6A8/4iCc/C7Dy4dOu4llakqldwcT7
C1soJ+VaOCfmAIGfGpEgnm3JY9KJwRckGH4acroGkv74mdudqvBh0aW85ndgbyOMr8tZujpjaVXj
MgltHBtMsILt717BBwAB4BWH3uDKPIdi7Q5AJYOoNcbyA61qBN7xznMa+yy+p3imwJZhb4siXYah
INgU3xegnrRy0ED/xZ/FIJoMabVeLMTSdmVo8P+oaMzQWx6nDM7Qch81zZs4ZbCts4ceoUaWXmpF
dioYh1vFIG3XnT+UjYI5p35JNRYFyRYqP1AB+iU4AQc5n0pOCR1fit1C6jXTIQC4LriwOygjPndC
jSx2a3PXb4SfrFi0z6ZV8JreOvB5w6MIlMLW7j7AA+pbDtGSb4jc9t22jOcTK9FkR1zQSboMPW7F
g092ZYMqehSrDPxEEbXjE+IBubO8tcAc7ysi+kgeqAWQZdAyRhMLoQ0YMwnlAG0YATkDZmMb5lc2
Z8RCUv2W04kUw8yxQwAnC1uYSEX0sSI8XhFWH/SyGVF8a3AcszNEYIUx/BfZjPHLlRLRRam9l8wT
8HKglETeiH4nyI9Pzd4DHgaIi8EN9My8FsAwXzcjE9wDYSZCUN7AWPx9vPbsY3yrNFdhmivQiXec
g+VWxYI0u6CzfDA/klVZQFJMXlGwwvo0sall3UqruSdQjMAz+h8hyEl686zgs75DapRlrH30TLLl
ypNUPz2CU3wUxavLOk8MBsllA/lvZWjtZtoEdqjcnz7jJAOzs096+icOMkytSz9p9JN+P2QrCsQT
fDihcRSDx/n48dcKx2vmh2LWJb2qXA99aRc079HMjV0yZoCLRqEX8TKA+BsFe7O9uIjDm4H2vtcG
uxX0SutuyGSMTigBtS4TKLdF2pXRMz9MEB17B7C03GkM8qFyZJpWK1XygdRZ3TMAbiV2RHFxt77A
f/tTd8Rz4sjPYDSI1W/XPwvCBz1E+plGNAoTJOoMoDuR4s0weYAEeoTIbUeRfAx5ublpx2RLr4XK
w+CsexBqz16NCbP+xDoDLTqzYENr2/o4euPHB4ElT3X5qE+tiAVBBAu5utFNcfuDtqX6SFMzo6uU
3mEGFnEvSErmAZqfi9DB9ciyVRCOF6EJFT1/GTTj7dyKTo90TT2eVuPGhOLnuUoUv8E9RQfmoG9e
qNqz8BCEMmGYpjQjFT6i1oN9yw/orcpPoDuy/C4fb7a/APolAjH49T6RqwheHd6tXGAnVxupS9uz
5Z0AbP+Oek55e3142uuUhF+jEs7AX3Ygm89R4RKurQEvBSBGi2k4LracN047GThza44Mh4RGwga7
EQxPywaphEwG4BwttLubvYSCyQ4OyYghnKmc6nkkVg8P9v7iq0IjreG76H8LNrUOrRVWUCaWoj7m
UGNO6kVf5K0nzXlJ9b84h/NDI/1UUMyBUSc2s6XlgVYhQ8M4ki0HmErbWIqrMGLhUL2Tbu3UD6Ph
EYh1b05vetNBk4XEGtsCFp60eCwctpkeDqCJPx4XmlEi2gXmepd2DBY2TZzYLNxPpUffegNJIsap
tztKO2F2tAVxjatQ1SDd0Z746Evpd+8lP9uF6Q52k7HQqZNaFk7Z+Ixtcy5X1M4AzOHbGrDk/3+R
HWDe1s9pUSy1F6ZsOuUdqKtzslZ6Q33ErBlIdW4rMA1A7xfKZ5juKrrIaySwv5ePUnHvRlbXwfT4
0KqViypquFQFCE1uYrnVTIk89Z5vCP00QxzHj/ppUldPYELZ6CoabU3Rq/riQn8w9ZVZ3uCTCuym
6e10r/ER24eOOtNXICOgQ+6mY2xWBC3n0DNwGVklospFeb+T3L1Lt+HqVRqHRXr0MRGJ/4HXtDnD
0d05eyFqQp+vYC4t3GNO9F5X1Xvoxxz8L3ea7oUDOZ3e7HBIWHtp0C7X7nuvJNrzDFgAr/K4g4hB
M8VezL5m4q63VhMCvP60gzauq1snNsDcDrL1Zr2y4+xrLwuWgfIE0lp/yC1EyCciIy/Q5A6ZZzi5
HOQo35w7Mi+4o09bAL2w+8L0BafCjbt//eEAA9oW0J5c3QBDWUZS2DgThLpUeLrwd/a3HjLHfS8U
2KhKnYV4+ulfv+XxDZtZQCRqGdTDLGWPPpo2SlpBxu1nJbyrJqOR1cN+Jmui2O9Fp5PRZk8pzXZs
eKLqVhcNi5HY2C3sBfFNP8OWNtr8s5QA1qU2GKiLKhdmLcRvgIydpnfqdyJnK8yBqWeS6/Kf98pR
i+2td1+wb6bULIHRDpYgVf7yoU/Bt0Hk8SdVohKgtWIdkh2TeWvcMM4ksJ1PdWFbdmE2jvmLLVd4
vj6lU8F4EFZghHx6LES6fXo11FJQb+18CHvz7Blq2zNEDgXT8HMn8gKvj5t89Jmo78iYYju96q5B
PWhzZi64HodVUj4NdgW9MVhCzoxZqpYwsN1cnLNvFvav5YIjwNQf6QWFMke5Bv/lJa+H5mUBmLOo
UcoDTcghIjLbtVYl1xHJ/gwUWQv0n2U5sBAGPhUMlY5Xst6xYVxuGGUX4Cz6xsLcIe/RZSJTBjkx
TqAlczQEKk0ZS8MxoJntmrrjXzPlvDXWgDMvRVVSRfLoLtZifkE2XyziuDco3LcWMkpU92QdSUxC
FVditUWAmVZm1MvvvYI4DVy/wG3jq4Fv92lVkRt0D/FvZgw8RC1e8QFe5fhbZ4Wa4MDMdc2oiK9I
iDwbI758viJMImMSjHuaRLUFk23KwMYtSokS5GS43Tl+J2KNm4tXnLx0ERRZuqOtYtM6vHR31DJA
flhAi/Kqwc57Ad8RpUcFnM0BSMZ6G6gURXIQwNZsfuwtVY8ufQi7KS00sEa2yePvDCrARI0nyedx
JhiaCl94nthHeTMZ6GlRirA8FRPSbPrfXK3xbAqmMqGHchbAh635rvhlE+5D7ErmHXGR35HjQKEP
F5M5YyAaYRU8uEUY0oaK4iuVPw9YrMLHJcXum8QsBOLh/AzmSGGm+pkBRYWSGaZshpjNGLubbjJa
R4iSkEXtB0fGxmxJOum9r7tLr9uvisH6FRJnrBFDuA+9e57vHniN77VIc77KzKI7yaiXag6VDfJp
5+zcaXeg9p5Lr8xDTMkQ7ciP8GoY6SZphDhaNrRv25lPtwJdXDJobhenHrdzlhSUU4P2Vy1/Z095
UUDuMC3SWQVlbNcSFZSoDzHIR6pSnszuUmP3CRBWk5RNaES+afNj/Me6AkDwAq/xoZC2ejnogzIo
wlGSfjj0XQXGNeuOq/XI5Ho5113zSdbXnWw9VDiYe5/DLfc3ybUVS9L02jMAQu6Jia4L+QWGE0zo
Y0LK6gyt4fQ21vt0oeLkwrIyeTyqfMONAjL4bvqdg5cNSbixIuioKAe11TE0MpWAWVBjOThU0twR
khc4QKNXKBtE3IS430WWh0C3JYq7sFeWD7QhTmxQBnnYcg5CX9TVZR+ob3Io030z9w6VcqWxZlFq
oypg9vX52DfkX3WlhgxDFC3q9EGAmMwvvwtoKS5cP0UNlbtb2MibyEFotBo8OApy2LH8f6PLjZ+t
qr2C9yR/R2kSVmljIuUImrFpVBW/Qj9TP8aGGnfEAPsU1qNwx7gEm+Za1LcbsEpvo+CWCoZRvXo/
ypxz3+0myUYZeHPBiJn/a66fUpU6v0nhgOOnViJKIeXqW+HcbhrCIZTU7nUUZWLQH5wFrsviHpRs
BIB1qpA6TLghlGuz6gbOGxpzk9jcGxRVk67h5qM/fCS2Unr4rc30fc1JCM3bRX3N6mfUylGW107J
bYe8GZ/JJgwxH8ubNw46ey9V28bq2edQXsV1hg6u+eZRCFH+LpaMBeZCtbr5gb3Htm1QTgGDccgo
HD6PJ3bpw6Ms+Ksl2m93tWY/N6GvQ5PF3EJyfa+idFCEaPOELYFAyTKWxeW2a+ymbTCVC5RXtsi9
9XZP5D6MMrAfPH5LJXLiGkU3jdxyksUBO+8ujiWu5q+Uaog1/darg+f0NuEV60aJLiZROQFFsHcj
zLB3qGNi9RF59M/F+RPzLxfX/BBaoIVV0rahKLPUSaVECAUdRO2zTyjMRvk4r0oqNBzZKmYDo6TT
Wjd3KEUKO9v/kJnwN/wdBmAfrM8Jjm3Xwwt16Z/om/AZ2BGZW5M3up3OGR3Z6fIlXArfWBhdWyki
BFxiQPpFmdcDE/J8F7Idfr42ey1gYGyJpuam5AgxaqoHA75E8AwFQqdVkMNTZeCqy2Y3NP0LWzo/
9B861TFDwmLiOZjOf9ebmI8nKzG6TOPvDymx9C0qWeR8btHQeK9uIGbEfW5d46VgqI9VYZvErOzX
rducxJAeJYNYAdueP+ck+Xh/A59PJ0jBIlzYgSw6lcThMrjRexXEi28U8Gs4EDCLwoGdHCr6TQxr
AbsMzyX+dQIIfUmoaehVldX8nru5VFpp9StaUFyzTw1QdQs8UIq+O96jVMaRHHZLVhBjkogrchYF
ow3QIR5YsLK+5FLOyloX/3f5yREK6HTHb5OHn8o56rCmhC6yqoDnBXj9sfe/y3wethaZi8Fs8jcx
8HXSUvon28T7hGLMeUHO31yWUxygJR+t5WI9zucXgtZuBTE2Urd1WNeXMiFKC9XWZaqJb2DH1I+b
ob8wRr5DtqiV8IAxbpHGemtOYw6qkcd8a5pNExGqntjQZABQeqzE1s6QiYL1N9urqPIO1jc+nhqR
ENZpXYFMt0v4tpnlItuWI7t/Rw+DSmQd5/K2B7JuKWXBakG2sq3MUznYjafTmDG/fMU9qkPSA1ZH
lEMqcUUH8DQBkCHST8idELOQU13iGv8S+zXoV4T2+lcYCf7ceYCAi72ZfJOYZHc4pJBCySgr0pDq
EZGUzZfiLmNimqjaqsvnA1yWfw9H3n2CBWSJjlhKfSc7vwoy7h28qf8apELaOS2NH8JFgD1yIYFA
DxQjN4pbIXg7JZT4F2QNVUdZL4xxk1OmVeorw7l2/d/ClLJ2hiVfAK9PGYPVcpGsqLkSqlqoA/Fs
f8rZqoxdIJw009Rfg2g/0nRNBi5uc/GKDTjkfAYh12qonkwpB9mdf0LpONw73Vn+TQOcwF019TkE
Zm4VPP1Cub655CWuJ2dUz+n0BKJb3OEX08Imo1wo9pphjXgLhiz8nQd6SxZjnD6qSs46rS/u6w9y
BiwPliJ/ma6vPc5FhO9nYrwNel4EOcsnZB5c2K0ANYKKlx1F46BnN+dNZg+zyKNgnkysg0tRqDGU
ReTcTtSajHRCt73mg1/LrNNSVXVMkewxOzZe4uwRfAAIfUUn/aDKbexLIIIvvcNyZjpa51/FQRhe
e0Fr3yGoU1jUM2i3LsZWHjVaktdJWz7Pdt2V9FyutysMF8fK63YmdYnvZGcYB3wFM46PTgqfrRoN
PJ+zLlnGfZfLbtjrd/QbYjSz7lxFfh6BLrk/EvK/sb26ro2JiHH1nuuEBZM8Pgib79q64Q8ZZ/dq
gtNfYKbeBigpuPotEjSI6Dy1m3kLx7gnaFTSspzbB7lSSl/vmtcWleORzjG/KAbA52OSkIu6fXVw
nz5Onxij6NmVyzn29G/Fdl5jI4o9P6KKEU/VLCRXUavhQU9818pN+laaOpui8vHrQQHstIz0nBJr
sH9wrceHrNLWiwuvBbt88Qm5B4HbwTuqMThBJcpuCfSw9p5DKQGG5GZ9qBE0rSMKJo9SOKteTe7W
T6tGuQ08c/Dw8USoohf8r+cUwMlVkKOmPab0z6gevlJXTO+hjQm8Sus1rlFZei3pVVZVg8srQDUt
QQq8NM2zGQ3jw/lmmyees5mbtt1izq4Vjp2zx6FJM4Z0IZGxOFHlzD5XmUbJjQcm9g62sFN0aOKH
1Ic8DiH5wu4DPoPwMNiPVgQEPZUFARWzMryd7Qc1/EeAvipQh4y5Wm/je0MCBXKXzj5F8dX9Gk5F
8O6GypBErxmY8wB0iKWhMYdyDjvOSUWiDCxCqFhC9P/16wQ99/PrNu1dKTivCoK4Ky139ZZWzjR1
fyifEIp7gQSogXUmWSuI/dovPIFVRc6jDxPOVPGedsLu/KVyn19E1z1t8NqqbRboC1I0jfR50f8G
QHjjIrDP1Isq2JWW7kvurqOcln1a9yyIvvvKV0ANpGtIyn0r5tMR2So19DuNeXoHvbRdcqpotVZC
4NGkSxc1UTnKG6u8xt0aLpoNuIbwr/Hkfam1J/pU75rBCpTOx4j1vY8/+kShYRlgpv6XZrErB0Dt
0FFQO0DNIZSNRBob8yugQNo23PbnaBqy9zQ01yu0DMWJLfYWQhOWEcFK1yiz4KujOaJyLnGQ+DrB
GudyGLzYFANYP1rJjzW3bqXGeEWJ2CB22DO21FcJ3MXZFLJDAhDx/Gba3jNZU/xElAoptzcRdzFA
rtu96eLCtZMma9cjXFciUm0fO5JsQZf1iam1JFZWQttK4vtXHeRxwv0pvzliDNnzD6yuyTW8Ds5g
Jh4etBq2zFC8KOv48BlVF4OdfnJOe+NeeCKzIzukTttmKlaonXf4+ag8cOuElK3EfWsjMV7I6Zw/
4bO6oiS8xFNWRUCvDCkA9FUaHrV2hn6W7wnZGIQ3z3CjNDKfbKqEX67rNKlvEJ1ShYUR3VAlJXNn
QcumpPUDb591Bks7kO3hp8gQ12iGA35zEw8vDmG5M6EmbZlMS1oDl8sr0EESvB0E6S8POMM+RO2a
NTpKrq6Y2jcs3xCY1ps4ea/+CT+tW7HNQZE+2/mIg/ijzycw8N5yJSYVX1LQeWy1VK8KMGYXiQL3
+u3lVjEyhwpIvMQY1SBOziJXxULyLTIozagl0YcqesGMOGHmZpwQQqeNDb77Cbvzu9k4dX5D3M0z
SUWteoUFjaRyJUCE+VMmXdM+Czsqjf3TO4gmUyWkMhwynt5sjzl6Zzqw+9xf6nW9Qm1mhnNC1Jge
SVLHy/GVRfYeIdSfJuzyA24/Gf3zq3YytcZl/hnKzC2idJ8DZoTYpFgEdjFGavDS0CFsoUJhQjBD
uQfZMXMqyfEnhSDJ90hST75vK3291HLo7TFoCzme2q9Yrlrh+TPZr/DfEhdZJBQijsrhuwVLqXqk
z5d6Pabr1lBzXuJAwjkgk7RjhXVCPqiODTK2mEnvJnE9uO0oTtr176ZCwQniov+It/SBBk8xan1Q
R6efZ5F3k7kseO06uYL2trV26OTmvZXX4XR+0D9Gj1eyczNntmf9eoIr5mj6E9oq9YUvVXcT3q1j
aHPsRu9/onXBC6rZ2mze5f0qoJNgipf3+C+XVqXEJxjGWdElRUuE59y/xzo91/wqQ5e1DFfx5l70
U0eh4Rt9pvaXTohOCYNdcCQlMtpaoFqPNhXOHdm53iUedj4TP2li31ry0BiGRSfSxoC7SRBtiD1T
p0QE2R9XgmxMJD1rx8mp5lNeZaNAp7RCoCPT1qK2QwfRjLmUxvq7uvgaFcj/vPlfs42iinelMRmn
zyA0/gIl9KRgP16Ucqd4M5LAxNRxFxRx64KBp+SWTgc1hBt8wF71ZKPmK7jvZxQaJcHwvQ+FWIs6
19MrTDj2/0Wi9Fn01w7E6uS2zbF0vtPcOfpVvnI6VcN4fzlvRpARqoYGdpsc48QrMTJg8Nen9wIO
OBjr6JAo3ATV2/Flu9JCUACyxFrAGZ0d8jbvcdndeG+6DRhQUQNJ25H3z2sj3nqJsVRJvlBeZoYB
fotgSEI/tVV3z0nEF85hA7/0HhzwiMCENs+L76Zox9KEy+7G00UlKCYcqgJwTvrmd/Z0MdPc1F7R
D4RCcRGq6VK+5froRgZ3j7QUQ4ww52j/zgwxdluA8HnEVOXA15EOYbiAm77WWcrRWWl+ut9TWQWM
bvIvKURFqu3JgVpDGDo2l6MsqhGuZd3PQjb6BS2g9ST65SMkBWrp+7MMaFnDVqpPWftqZebRC0Vm
jtwpBNkYLtjyU/cudY4b+pt9qXvs+2LDOsqhr1QNXcbOBT09ujw8r0Ch5SKBTxXHednVwsBei7Gu
0p/IBn9S2RroAiKLTpclNNjsVE5IV7rqQGHGxt35oJXcafe7+1kR2p+xrfddR8ICMxua2G8csLlQ
yF/bSBFJI6nQju1hwUqIqZATOA87lG+zspbvZUf1CB1CtCGx9FoyPrHjpi7vsXPIcWFAL9aBtbxy
hqk2XZq3zMfV+8JfXq9FpmhKVtNLI3TCqvGzWYGyxsm1vudm3DU13sx+r3y+G4cEC8sXffmCzrsY
T4WOOrsWNQ701l/rqNnENazTWsJIvF4hpB9r11qaUjsDf8WyA8Wp+njEF7c09FsOTXMSD/24g/q+
Lwxg0fx34WyYZzxXmRmipufcKFPbw0a/otYjixFkKAvXC1cRgZxpgBuFZo+5jBFqOcN0I9rsYgfD
I55dAv05IwVXQAu4HR8/h05atoW+HmvsIw3aVvn0rz1IzqrHOAfAGqzHt//S8rI9FeakZS85qOMH
jtyzPnreTtwDai8DhV6C4p0/LDsrOI5Ds3+QWL19HvSoUaJFX+IEsxXV+Tew0BrHg9h0jqSpTad9
ksxUreDZixjKZoVyiS/M2mJRn7mVZM0sXl4vl7IVrgxCIQTuoqIPCqXXsjxvqdI9fV90yUKR4rwx
IKigXzOHTkpKNynKk/rpQBf149a9iqRn3q4NaV886C8JsnypXaeLUgKz1y8m6ARYLQZEBKc4kEzV
baw3Hd/5ZLz+u9ysqxphsoxkTcoVZLjKTa+hNl22zf7gg+RV7m9+frDT5qbu4Pa6VlE3fc/OzxjM
K3rgEaVDIXAdF0SotQnTint7dfyvsTGS37FH49euOSHZhnnWGhTdYbZkY4a/tOYMGV9ZZT09QBQz
eOPPEA5CuCV0h87BVMHt4awjYtM7aSyvo7gviQ9FOUxd40Cd/K/7zIKteaGNbva45+W+GVNyggGK
6HeGpAOVFk70vqm6z9w0OAMlHcANaTvHRfn/h3MaVjJmy/KOEUG3rKpi7F2/Cz63n3rUuWB73iFC
1jPic7j3XpXaK8omS0cBmpNq3Z9dooOGaEC23MYVQc6nAobQOg6Fxc1P1sp8Lfy9BU4Y+JnT330y
O85LMZeingkEpx04VmTP3tucrUrrK+LKkUv7RZk+CyGekQSWjyJViNEscDOx+wcFEbd6pEUJGaSS
nc7ipXTbpfVUMQ15dB8UB2D7OfWfVWPtPQet/mBp/oKUibitDyV9JMDp9dlpAk4H5Tt/dm7h51ZS
HNqjGYIB+NZAgkRiVVNzN1AbK2IU9v77CnaTqvG+j4rSvecWLTJtFPLRCdr3zOURIYZZ0RCAwewR
pG1B1+Ufz1JgovfswRllWwrGXehJ1n1t9PYiixhTK0b3Gw/lO1pz5/zMvlaTD42KPe1xmYUJDp1V
Pi+hjAuiqgoA0Vxg2XA4jGMFtyxwaEnfC3Y+VmwR1AMUfyit5VtzQONG5En03LHM8x0B/W3Dgvg/
juHxN2HvyxBDLPO5WhAbilvGYZVX8JblVECjzJ2tgTiOphochWbaFsLFYG8iURtXoY7pyIIdm0xP
syYOTKlwbU7uwxB7CcPTndgRLoH7uXFHasEUQhfOnTpmlQxkBu6Alh+j4H4tL38rgatBVGOBssAf
GgTVx1xrrA0qc6NMU8RvPVByiWzCr1vlAeI/9hwNlI+6J0AfK++5LgsUXX89pauPhXRqwJ5rWMZh
Rk3otlpNhR3UwuWoOLFyfOdmxShH1O1OwF5Q72q297YbZRy7lo48TErgEhucYsWu69wZJJZtBg8K
t9uiQ0AUXqziTMUDMYrl0Mg02Y+JoBOVGqKTnocjqHHSCRa24B2iXJuoOZJ1o2rHySJ5gU0Mw8XF
rWv4/2eWVbJ7pxXaY8ker/MvCjnj/a/yq8dWUPIbtAsNGzE7Sx388PkHXAynXg/XAzjk0hK+xxUV
+9Xqbjp/AZNDAAkWgw3zFFcykRNf57nhA1ianp+bTzFJptQT7QSTBgkNrYN+j2i5lqHHLihKrwlV
B7Y+1DfLzo1hrKilmPJDZ6CdHYV96Nw7tn1sp4ezxQtTAJY6ef14/LDH950OQSdMmOVvZMaSAi8D
7B2HWwF7lXEIe0eE2dEayerTpMMvBUQI58K4X0x7fOooEkt9O0H8AedCyIUPYlCq4aKTera3SL7X
CWVoxvalr/YgAcnvcVHtxWz2JN9D2KmXbNnqcPd0pRJxVdZP3d4lU3PJlCd3Gnhjcra4xHoIYKkb
XuwVMMs+aAaacTz2FF4Fit7+2eybMZGuYLkgMGPiXYKM9TuJ6CVILT5CAsQUPJY8RsBEOy74s/0e
4oz6PGWTsNJKPX4LrCL0gt9DSQJfkxIVB3XUaAcEdJDr839ZmF2M9cIhQPIhbSCYX1FBhqEAL46D
4Ws1shLujVidfVuC33N/LOri82uQYs5jcTXUnbuYWyxc+Jdao/Wkq49yDmp8gJb5PlxnNgRTHSod
poL4ZgRMkYVKQ/xQT4qmRIw3uGzjIzxtqfj+qvQTm52BPAcBQMbuXRZ9ndYhONrYTtQPJLfJIVA7
NC0m7bT5yzOwJGs03Cr26yOOF42KPCXBH2ucE0PJZDK8iRgJOmsUslTj2/Xh6Yl7Uvr854obgt9o
Evbr8woXQgoDIY8MZ0hE6W0ur0DMA/fjvIVdDGV4KgQtYYzSg+KopfDKJ4EyCT2WpkKxCzwIOWYL
Zkuk1aXXk3vNao26AvdJAVcUQwhv7ljoXDOqWubmQBi50LK8sNGyFQ5yxSB0Xd+6/5aGXJ8NK0o7
fMPoFpC4BQrnXy9QoiI8eQrEgRDv6aWXV6z63YvJse3TsDMS36hVrvNGNy83zQSV8R275D+6RxY+
mZPT0UKXLGxu9wqiwe0VEM0iXBk9EVQ0UKW3zfLldveEH90Q6MunrWsYgYCBWw5M6Qwh6nbTHGxc
t6DGOV3jxz+xo3gRBgF82Tg2G4bPkyKLYkcc9wFzFrODphD+GDClMKdQzAGkcUT7iJupdVKH1sd8
4RJkK1BZD0qe/giGU66ojCBw/9fZ5GSyD2ORcXMCo9TiuIAI9X8CkUBON/0uaOBvIXsweyxZaoWq
tmb+044BESJuuJcCOzBvrNZUt6+FUqsxuc2iBFsCUGYSpXhhdvA3P8V1RAXDdWzZ/9KWts7MbRsU
9LQV+QdSzf8mYX06dX/vJ2zWHioplqdEnsxN90nQ8C8x2EDARbHQgpxcbPqARU76rgrPRlORQUDG
Zlov75Oww6IpY82ZNb77aW1HisMgG5p+QNgi6Rl/2fDKH8jWRIaog14F9YmRlSdbMfAkwYqDv+ul
9XLXW2OPNxoV8uBgdsZquXur6iJb8T0Yanwh6MFCUD9yktZPpyBRW1NdTihMM+nrv+HXpNvna3UU
YehnARu7C15rBFySCahrYXqc4Kaya7hV1zk6z6buYCdVv0+DItg4JVj2ZFnegQ2PAbF1afoBBybu
HLdsFbNT0fYwooeuKoi6qXEbighvXLJQbdf+I4TH32smcLcwUjYS6/nw4FyMIiX75nerftw5d2MW
MdTFQPWKWPQ98XXmB3YaJVINGk+qzYrgUsgL0MBazLZ1OpHXe/A6hy2uOLALTCidUTUvnUwlHiMQ
700cMaEHZwOeNAHsmJ2lpAN143UtKL+CLY+7U0VdeRym3Ngg3aLMgd4aa5TBD7TmcDz+vaTU+u/W
gzEhtskyf2ztOodunXI9KdiJcZLhZPpULhWLoeccJd5QdQWsU51AAeMIevHGNGjV96m4CdbNJw8m
CvdhAZ/YF+S16eNzVowAbmEASKNxrnfbQlXStslg1vUW9uD8yohfVhFA/UDE2YhgTaYEPSvPSv7j
tjTZP4czHCYLTE7UCPSy8HDAdZS7UHoSDylW7f0hJxt2t4j6yyDkCGnICv8gTmOe1ZmoGeW503OD
Nf+nrCSFS2gu9NyUctGp9kCnRN6sHsMTAfW5R5/wykOx/nDha8vxMKSGB0EN3AkX3CxLOF3DrqjK
PO12TdrRjtqkRkYubUR/Dao021V05O57hPV+upOmDTQNCSb3H8F2Dypi3IWQLeYrYcs67Jkuozpf
vV4Ef8YNdGcFSBY7TlOLj2p0QmL43ywVyQcr2kOBemQmAUve7wQfOxHsNvZPgRnFpGi11pn2y6xA
bS+mDA+0XK+ehou1MAmbLZykeq4JfxAAx7EbkVkycrOW2HgGH3SvGQAjni2FbT5V89VLkTY2j+fi
JZwOQFYQYCP+5y1uaDXa7KXSZw4zi8/2Z/1FFoGKG8+52sL/dOXaoSdxT2+oJEUhjiqm0GsZ+o4A
ww789E9F5D032e/gQDUvWQBs21M6NDE3B/qu5c/zKLYT+Ydbk3YEa25a1G6qYCQ27TAw6kFZVx4c
oNleRZImu/PL2VaI+36DDC2GvG5aRQuKdUvi/rNQk42QGwpU2GXAmDAG2iKkeWYh97tRsjui+dgO
gniVSDamQe15TAjd4R8KDkUoZlI50MBg2oJUap+93y7GwtT0I9lOMCSnNkvSj+Ud6Jy+opD+vywo
qCqzKqYHJ5OzV2K7uqylbVs8T2JUcoYAudJCMXp6d5BXTuqUYh8GghKef4bQULSxARE7qTSir6j5
WeGIhqU4EbxXIVKQEXJrC5opbT02qzrWev7BRL36Gn+71GVk25SsJ26moeSausIpqR3GrFhMn5X7
auSvxItu5UL6maVhmZRYdEl2h4e9x4NYf8u3MAasVeEc0vb+v1a8GTizssbPjI03ULWlbzjZYoY2
yMhqvkXHQWA3UXgyqQzLRs3qf+BQkZ+eWBu8nubItH6SRGSDrYQSAYhEw7mOe6A/9IqN/yeaqFyG
cGeaa6rmB2A9geVc8lO2VNanDaYc1T3NIbrdcr1MryuHHJk1imKzlp2eIU+YsR/yxKDtpSvlYdJN
+sXqq8HbZksK2wbRuIn3x6ZyaTnLsE2USkhyXjcdlUGMXv+eEuEgH0Oep/vZ6Grx0qoroAGvbDg3
BJMEcA5nPbOFl98q0SMqUo3EyMh+rza6bBELBZd3/ci1AL3w+ewfXg6Z/YRfNttkcyxaKJWF7fLO
3uKcag7K8gre+NZnceCvHX52k1Im7BJFKdq3dwA7LFIYWeazH2chPvb9c6QZrMFx1LODO08750Se
z2ZKU5YINSf472a79UjZbyLpJDmA3z9MI4Wjy6Don23oQWZfYEbUXBqHPgtlVAAYncHdv38rh75D
/xGsU9kndQyEHD6ATPegCsp/l2i7PReE+u4xm/nqtIqvvN7B3Jm95oBDeK48mRtv+WNJop7q81W8
y3/AoIT32JJuI3jI5olehzuheDT/sxXYF0tycx5DITZk64nH4HxPggFVTB1ML8ON8txCqx9E2lD4
NLCk8OgUmeJ7KbmJRlpvnlbN+CYUyz2/MrdCj/UrjfK2tx625e+fI4NuPtyGGTj1buBY3jMPidBD
HL3drBsY8lBknS9csTCDZz7DB/HHOSo0uB0GFB9fMi1y/CXKeSx/uDjIpjxvgDALxpdHaHhVpIDX
Fwt0eNZeJNPYpeN+ZWWAnW0M+FI8BybN/9ojo9q7trPxFJ/kaDe15T5ZDjuIODSGzkJEKruTeM6u
4RIuZg85INLuwhNVCMXF5I2pSIX8Tt1gAhtHVpRAK9l1c7bjDpzGwWmR3hhbqCv+nkTRhojl37VW
hKHv2al0FyDr+wgvSt4jc2I0W4lj08hjXR+GnFXqS49jEmWwr1BXD6vs/U8kOh5iIkNjMLoT/SWc
xJ+1t0XnA0xHOXiFOWgBghl8/3QGFkM4M99EA0LmIGV0D9r28ikYtc01gbk1G5X35brBamxL/RFV
Zg7X+RfZk4pC5IJNLOS7RK64PR+CGFNGxa+o5xOY2rDyrqEhRPZdD7mnTQt004QTpyuOFLna0067
ILRszzkn2EIIcKEVz/sSi0lwW7Ift3LZGEKG8y+xgLY2zmiNTFh6h06t3wRLHGj3PMwGh6Duj8kF
Fy1VMQiSPywZbNrK6MIWdMnuUVAqPxbzpwyxLi4bD1Xo89GtUwLK7FmqbckxA0fsE1qbJJtIDQvC
zzSgxoBqd7Y6YtZS3QqVK8aFQ+Ak57z6v4EBBB9MDQ19b6kEmTQGM9oOgF++sJo5vzJ2ag8+4aG2
mzbhjTEWu5AAkNOrQ5oa8KHwQPatva3k/27gdb+Ju5av4BQMe+tsF2wN89vTy1LocPwYW93nfK/1
3E49k0v3VzlBm0tlZy3EMrK8rLMZUKR1k3wM3O49LiVt4s4WJOVEcqZt673kAIL/Twm/Co1kMYrU
pDkEA7d9xZWJJcg3fmrnP5P3OeR8iLqu6AJo2tEflhY1TjO/cNy82xTBnNKQJbXZ1vpD6Khi+Jgh
UMzAcNrIDB6bV/Aj13vFAv6G/b9ZwZZC9uXt68ja0lqBqFzGXeEJaIjLn9F7dUoXvDCuECK8UE5y
gZA2svTf22aLhKoptsbA5Xm3UXsr8ZRiMv4PjLjcv2miWn4/VTP3pAZaDAeFFBsVTRcx92HFxRnK
niFzY/MahCHMk7V9ooVWU8FTz42F+N3InAsOUdpAC80PfYpblaTGYkGLz8oM67OiK+mYdFHXeIZb
jxQgd6nQyfwfBYGnDZLr2t1aSiTbaolySOrzoVXVID1Ukeq7XJ15YITBolOuG1CrLA5+1PRdCGTM
qoQ+CBdl+rKL9bft6r51/0trs5FDla33uHo82GLpYwLQlS8x6NZEMovajXGGe3k8pGyCnZrSBp0e
T013yEoshN3SRn193QGYKk7e+dhaVI+SJoy6D8poSUv7FSO2kegMUOy4709GqVvhWOFzDeOpex/s
Zkv5SZPGQslgNCBqPQTcqsignJxNbYA4F0ezc7tcaXCOyFQgHyZwfbg1JejZ+6gaw9JGn7bRBVmf
WkVY5kLaqLf6xq4TLFkKZ4MC7vzxaXwVE/v7PEQE/0s/9nWIK1ed0gdKyfbw68ZqkkRa/eCLIYTt
HmHfN9M5ndJMIXv8lexM2XKUefoG1dymcjabps5ak+54Iu3XvXaohCfqobaf+fWZyq//ABgUT1bj
yS1J4zPx0YvY7I13/n34xcg01le8ymitXcfoenDS7nIXSMpYhX02rS0n485Bv2Hsf8LlR3sHErH0
ZCyeG2ft9HXfblwFeJ+klf6qjsp3z2SzxIFBBXAhAdvv2HhF8pfjrMST9widPYV7nQe4r/f9FfPZ
ZKgASPLtOOWztZmZjzE5B/O5ZK/rKJKhBqE0vYaf08iOfMSqt44ifAKJIFwAYVin7AiB2fIHIkvP
0OfwrZJc7gjGjW9gQIB/abvuH781sThddGXpsy7WKOw0RCI0PciC548GJKVmlVBQK6SbMkBgbI8P
nOLdHeuqJKhsdrsCND2gDPLrajZOnW24ozPfS598ug5+O0df/2yZvMRVBejQUnLLF3Kbhk72cEyk
2tqPpBVx/+llMli5H1Kn9OeybmJMFrc1xJty9RDgfoWy/5g3itwg+XNJAM1+Ycz6fgjon2Ej579p
4F+zuNc6pV1xRz5t3+CSdkSSQgplZ/CrYUewS+aUF2mKLeOw3o+12k6ZPcRMmirB3s8JqS+jFXyT
oGrvRL74kHDn1egFQvYblgj8nB2P4aLb4u4pc/oXP66tZ42TLQFtxJan8usgBYRn0YRH/SwX8Vys
Fa//6Vj/jhmcdyEgiSDZ/4uoBmNk2pVvYq4AvnBBLxJmax+lOpowzVSJRzwZ0v+HmJ9BC/EfaUHq
yLtYQtPZvk+qOxWbLpOw1DxxP6E+zyAD4zGVTpq8XUhKh0+h9etgD3UaHIEqxz25L2+zyxph3X/u
sNuD+mdqFMrXi0AjtrOEMj+fUGVF4IRr25/kQBX7XZk1iH88MXp48ep+yAfmYEz0qqMh876HJr4B
4uXECCJi2MNow0f1nPMzYCcbMGsjD8P2JVvXLy1CIyQDlOOeBS5Frnp8lDFXhJNV3eFMUd5uOhbe
rVfgTdShY/p8iV4MS04vGmftieO5lanfKbiFOK48n6/6MHu7zvVSqLx31jBxtYf5T6n2l86DIVS7
vsu3zS0BzbkOjb6Cgco7SVKraiQIdMkw3dWw3FZmDEUna5W7Wc0JI52bOL9wlp92WdvMwLLDsAo9
huPx1FZfMIj4O/CnLUZ2I/TubETkVoAzchBDSlQKLnu1XKAnc7sd1BZjt9fX5TJdXPz0uZK0dYZF
nYHQbAOJM7fdVyC4xJFiDxaC81HWXMXFn0W818kreOz1waKy/5cCad2lP3+apnkj/0/Z7kkxssmC
2A8WJoDuGwQEvHC3TaYx52XaR3D7KxWwzbh6kljjbM33rHSY5ositBzCp3IL81/uvJ45fkvvIetW
uXMFv73NoJJU9U6Y+xc1KIZcfABWeZEfBCQO0eLFMzDJ7usmvDMUNsPcMjxLY85gLo1YYNWx+2Z+
NKPgui11DzELGib3KEJxRaghxQOZ8BqnT5F1iI87CQoV2TGhCQeygRawcmIft8ofTWYeFO2gTGIH
JSpmEPa78ozol0OtBeLjDmvYvhF2c/ysUU/sLIZsgk33RKdtgkdqBI5E8/cPIGmnijVb2M9lCkAF
q1j9nVDgPI32UivMeFz3v/nbDjjILvj0tsyKEJ8AbDg/DF8KH089LXlJnoyH73SKrVgfsSVzfPo6
W1RgdaMkIgSuRWFEnA5uOj17fk4Cr3TFZoiTNutb4akyU/RHBH3o8qzaa286tFWZocVChnijumqq
imjlCvFfOw7+Tv5uwXgD84ThMkHbgaLR8/eiDI3Rbvn5uFHifa9or1g2FCxN3ARVHHN9K4DLaO2a
nx9093is4fPZGSLb/qXjaocyzP3eAhiEpzywDU5R/ZJJR7AM31gXieZqcwbYxLcggWQSsPkqKgTV
cXDp9vOKpaB/WXOHcEFRzxPsZR14qdS+cSrcL/2fYV8IJ/95BMakrMMv2htDv5ZnYwDfAgxrL9xK
HYul4W1F7r20ubBqBn6sGvxBS6R9H4rE1YfjhrcXjYu8BQ5YSLbcUdBjKw8PzrbXHHy2YgNn2swA
lV6dAdq0HXz54+hxihgwhqnZiibo+nSE4PueL8w7Pvj9Pvqu8p91tute6TI4MTOOGGzVxcLsMKK1
3i9obQ3bjlRxCA7ASmDt0ot0tklAsCtt9lSi8m7LHB3nIfHh2c0xSfwXyVPt+y3sd4Gk8F6ZlZyk
jaSj6WbW8mtxI01/RHILsmQZhiCV4zGjXkYZzBIrardcYeWgvn7x8mnG5k9shCoqBgnCdmkWHMQt
zEJOW/3lpVf+Oyp31oLenuG1g/N3A3rim6FQAy6Gi56PYD3HZoDqRF/6P45NLrh8jXCQ5nmgllVR
/kmEoIB0EdKB60RspXHlbjrXXZAyIxv+BodZbYsd3z6IM7DOomy+JzzkktC1JFtDLy5zdga6FD65
KIgJUQza9CdadQSv5mWQZKDasiE1xujlu8aVz5TRtSmzwS6jNgyAcw6kF+S3b3bv/RTuAW/k6twe
NJnbz5GAe48/KLTLJ6O8DOaU2hUYdgNf6W0Ao0E5Rdg7Idv5S8ZB2EyJxRDyJroQy+ufweY3CfMx
hM1bvQD4VNGqiCIOsclIavdTKRUG9LRPazYGCk30RvR+PggHDZCKbQgLT+D7kk7gZ/RHGcha1Kb1
7CAkQy6FvY51gTfPFxVcgZsCR4j+I0gDbnUQjRie+Ryi00ezW8HSdEktgD/knOJrEsUjSDONjRUB
DacEPE3zvbL+gK2oBLZYC6IUTvMZhXtNnKUBGzWADv2lranymUY/FOJW3gT+gfzLcvvB+4ZSi1qs
ySfRP6ecj2QbM74cqBxJZp4CyZeeDGRw8E6Z7TZhO3OU/iK4YqemOarbBJPHCxri15kYA8XuNuU2
rpumUH2RJn8ZE6MqJSW8kuvq74QxZwV9e4r57Y26iSikr9Jk4vvsX9DAo4sJrSnKYk0Emcy/zKY5
fCih9kxgZs96yjn74gcVecdudAbpfNJQhDUFaZd9H60/G927ZXvg6jOUGdhjEtJbxkEvCes5mD+V
w/aAiDM/H5P27x/kXHGRDo8Vn2kU7iAMOteIDYHYZ19DTfYp31Zck1/MpkIiuOJ9uIoboI9/sm0x
A3vP2tjGBCHrsDNzcI5fVHmsZDdSiO8sDoZDeaXUeFuXp20urEpRQpNOJfvx9ERFuOw7+8h7Pu0w
DCy6bLT5HwWCDEC9CAUwPrd+dQa0I8kCb8+MgcNeEayC99wnz40bTQPdQoYA7phOmpD4VsiFlApS
vE6KCTlKPox26VqJlN0Jjv0YHCtLbPg8a+90CNdymgrZxjJyaTI5iray6TYmW67Lq6aLVwYfySQL
QhuuVTYl1VrExoiTyWHzt8ajD5Ls/4Rvd4OFCqDh5SCSBJ9wouOL657mUdSFeXuFaUHeSy4Lx6mz
VKFtsPFZgNE1/jDzvi7UgnebhLbyutva+yM+7iPkOWJNZ2iI6daSazykfybWuNjKn8EuAFUVuoGm
cpWccjdCk6qI23kpZPPFY4xuMXMa2VzBxxePqPpcJRhepdM+OFPMMthBGMIpzHWqfWrcD/WorEVK
alO//EbUSmdu/Qbovkg3I7Jr/YsQme/9LG3Xmv8O2Hj6Ghh+D9h1xcSCNGA8PLdHqBfQtK1t33rP
os7lDYVBS/6mbq93FrJhDwP8fTZpMxJC06iUrR3QiRzE42RszLWvlp01po0rqbSQl6mx1Z0bvNXX
Xwbi+kpjUBa+jw62zL5XIAA01+OMxD11cFiKjERrg2HUehK6THTrrCDr2bZ5neq87rJaXJDqDG2p
bM4dgZo05xDC3Mj4JpvIfoy6i3G7VRsC5jpCEHDmdzS7iOqhGHWyhsD6xVQyimr8MT/Ikb/H6/xb
X71jgInutoN0s2xsIfHg1GPEEnNJ+WwGvO0stjZYyDOIQr9TxgBROG+gYVnF3CenomtHNIzPjl/v
QEVTt/zVZKLEAemn3hkLj1n1enQfeAb/6CINnfy2WBkRQCL/uCW4JeMCr0zsbZ+IQiEpFDQZsft/
X3sDRjdTfWpk72hVveNTkxbC/Q3oIIn87YgO9XNkSf9cv/ib7OaLStiOUgQdiNw37PVtd91WKKcQ
5g5XXWb08bcYzB5m9b9jbqco4KBwvK88WWRZkFjiRD/lC6d4twYMbJ59xrSJyTtyBdH1iOz60WAQ
8UkUqWwZKrhVkhI3JbECDejaDW5Og347omYGCXBeSWXh7A0PRtAzatlkKDllIGC7tVWL2SnKvnK3
oZ6GkXxrNJV8G0pKCUwecOzF4D9mYUVWIYsRK5V69QmoucuewQ+Q/Rsrwws1NWSmc1LIEOOHjaZ7
+HTDkdWeGJmsIOS+CuOsLFBGGw2wQz9P5N6QBH2a2oICHortLdcHGw9f8TwHoAGtgyYbmTRv5IfA
ZXbtk24CRUdNs63i0bMuJMwPMkHjglA05otMgI+O80BvxBIMlenATXS0eUt0cMrsUKSrnVHb9g2h
dwqMZIDMaUQehY4grw/HNXpdxNUXi/49JAots28IVst7I7WdyHTLNyJKZ9F5t95n8Cb1IOmea2k3
NWH+FIFsxXGSp8Uzl5E3aNWdwJLiJpUSvHeQionCCIX4Nzgh3thscqzsXT/Y+QHUVyCaG8VHpg2W
+b8P5LNJz+Dph49Fx3HmHuGXq0WZdibV/xlclCtJI0hc5Hnt9G2v3YAAdPPOdybO9kpYkMjedbh6
IYOqBiiQRvY9fk5LBVo8u9sdQKMEagGTwpwIAI6HJQUUJtgwZUpL3/tPErr1KyZxUb6X/Y/Ia36D
TnlxLocEmOio+zyzoSL6d92yn9QL8RQEppPGApFN5J2GE/SLqD6HWyDN6JZaBl+d/3rOR8iYDb2m
47gN0DlIx/b1GG8pP3DuGXWmlCk/6zryD9YuAFWXlZs650NjmgQBUEgByfQz/7lHCykZJD4W9022
/q31888nMKZoWIUpxMp48wPfB2B0WwHn+kDP3jJtIlUdhcS5WbZuLMyeVjmFQdar9dPYFSfRPfKZ
N5c7gEwOwFbuAqTJQfC+phSRdA5FG5oPckGndhYnQIGj/4LFC6LqwDeXL/FPHySNA759jLW2Cip1
P/49wwYNnT5knVzEB6/ITuUs4IapTieV/qiwFV667nIJglu5zH7o+orUCJL7neV9nyUmLwiIFSNO
0vvulh0NvjVyxZwSCuOQvBxNzNqR8vUsTdNlgTUbtFYz9oh+bEoZB/qnB5sFBQtqrTHAVpDkG39T
Sacewy3Gtw8Zw09lMU+fx3MxTCNaQGImr4v13Bi0t8Qcg8LcX+YFNcKUYvDDgtwVGf09nCpQ+0vP
rReNdZ8n9PNYzKSooSTIwp8Rnitj/8gCNM1L9CTx2lEPALRiJvsUWnVIS79UB4x9wuv9h69hzfyB
XJWBbwldz1uKa2daKWRB56FaLwEx60JeIIWJhAxGU4XZEFbxGoin4XW5vIqBM98gBgSOSDW/TrKc
CiHG6yBDQLIJIn9B1o2MW2F8QY7ckEvNeFyVZiWMgcNLkVEy3ZgNSmzzRCGhzon0LyLMw8FbjCfK
hhAJ4RFA8gNrWLxxm30sI9pSXZ3UqoHhodEa49tgPmI7jgQK73bXvOnt0rRjoCMiFi9tz5CWTEgH
A7uaOxtWcmjdbxJLND+YfCiuquvKkzU8/iHV6XAlFCj1tlIR9M8N+dV6xUc9J80EQbep9344cgl8
ndThknc1xfqR/HOrRLIx9nRkVzFRIwOySaYI9lWzTCHXyccNndP1wSXJzVEbzPtFUQLgAoH5VPk6
sycBoCILAH9LUNmIwn9BdePIce5UHjDTkfIjBB45hpaSWisNU96T7XiI2+k8Zg1dxkmSa1M6AW9e
pla5MLTNnoqGNy832naelkhseV8v7HD4wQoOFUdMDBMD2vY6z2RW4lrRNh0FcV6hS2y1NtwBnKnV
3+EImSkkrhr4fbZkHOQzRn0gkS/a0jFz+Ukbj+1JcF3vKZl4DJsIWMRLeXKvdnX55YJnD2Fcfw8Z
KX1DdCZT6+l7ImwLhZJhzMAiov39HH+dihSZnSjA3EiFMuSTIsOxCnfJiIW6Y4sTWRlDiErWTNHO
E62FBCnSHASISje8gG704JVxaNsy4P2iaLB3jlh8Y/bnRYHEFXRJ9ZcIutHAAaJ6I6Rk3b3GEYFN
R5rwvgC3J2IskDP1sS+3Cm3UKhPSaCC7SlGd4Zf1mvAVHHychXjy9AsmeFEVtWv/sx0FBfu6ILN/
gbDAm/AV9u+jw2KQNZ4CkIe5Lr9szAHKaYj4XmkDBR7WP+Z5hdpLALs9LTGN9eECG+XmO/gN44Bx
CXzxKR9ME8ayg+cjARmveI2WXhLtU0pMmd1M/w4ZU1TFCS/eB7GpfTRVNKCRQ2+sznSgxXyvqequ
5VRXEdQZzb5EsXyOF56O3x7qidhWQQfHnqEaapNfrh0zmnhj2wpc8LVHBQb1TcvglcFbAv07mBtO
e1/QzJixxaZtWa+bDShfNYPl94bwlvXRPbAom+VmD13aOYi0hUttHCSyDY+D3MoYImUekeg/GnKa
4TMizTMefmjSu9BtTkPPXDwVuHVBaU4yTqFG+7D81DPuH2qg8BnBkm14GGfb+6cZ/SpEjmVvXnIZ
k2VZbrLBaCx57xI1U9oM/sSMo6o3B7e2azhKqh+CSvjP99I1urA6XYkrpxo3LH/VTkNRRQZbV1OF
QA8FLeeLXggMi7UNwfrF/tjrsIRwEo5s1NdE5MwbrCRH9AaJ4zbIFxWRbgbQ9bNdHAnm2C41gEDK
NQ8LKVbaRzXbXT9mj47c8N6i2AzWtQaj4ypGu2O2DKYrAhyWXe0GxIus0tipIU+V2csDEoQwJRdJ
x8GcY28jFIbNA4oBZU2kuQHGvmXicZdVpUdDhaIlZxOlWLUlAjuLSkntV8/cQQHZV2gjttmY772D
FZwE+gcBTfSEwl8Rhheg3tj503h2WWphSD6DNkCVaUG7KbtBWcIyIVI7YXmoga6eORvPm/uXmJR9
/5RhuB+dImEE2ltHmPdfG90A3dMOvIreryTBQzfAKu2qBLZbC1kYkhV58oIwVbEnu6XL2rvku53l
VxDxVCtojs4pn+NTnD/7Y/2oc7/ciYR4KeJNZklvrb4+AY6MJEV8Qbd/SUdEPohn4SvU8vGNvXvw
XBRlGwxF5WBT+ddHa5VV8sMxKJT6yb8ed4i73AZkOlwevnyNcHUNVOtV8bzI1vymGrxPDhKmvMWF
Rhd/hsrDs6nEoNDDSXMV11vJnn2k8i3LHW5u3xugfFNfqnVjfGcx8nO6FvDOMHoq/Rlh8kKlcutl
xaKQraafBeK+DBDhKrUOQ8hkL7oCf7vDQr7M7QvjMh0d/iAb3YvNPEpnTB7s1z2IU1Jdkd0KlTPP
zHSmgHbNsb/aatYv3bCNR4Jez8QlJ5KshxShxQrkrTXNmmU5zxLHsrrdOUtkb/bKFqAoOwHuf27c
KcoRg3R2T6PPCfXrN0DIp4ZWW64Z6d/tuopdfwIe9U573JLIcICVkeAoB7cgAquOvE5cck2bphzd
1e+kfspm0HScvxlZP0afA4csNIiP9w+7jOzmd+wis+7iBWM9xCGkMTOjl4Arr7iyQUS7RY804yPU
+VJTvos2+SpeIiohbpGoE49VgCtCMBD5SeiE0Pjk6cFbUzezsqnLje7mURVkMUG+ASlNq9uAIKuJ
LDYngCB35odl1VUI2cPrdr6Hp3xbA6HSSQlJYc66Tz2BIzo5JpDNLWlEykmxGyV1SMJxER/Rq6o5
VNgaNT/sg3766StFjtMLXQR5iN+i6CCNMG/mmi6MzmqLKN19mC07LiNBpdTyoTQH2sFW+tBtMf+6
Sa5F4B17EYgssNCSJa6Nd2H8ZODbpesvvywsrAOm2phrC85dCy1dK2e/oO8BIl0kQn+4345rPlKJ
FDXdoZWDOGS9Sz/a+m5XUAoVPRPcA/CAvqcKtGs+zURgfNWqQVxh3tX/++OVh66aQ/g2By2wc8HL
LJevIo4nb1nfA/MM7lbQMeas19MajOlbaq7JGRZ7zhdqBjEkwoDDuWIa1ILBPWhtj9Ncsdl5DqUp
feb9wFz322deVSt3C5sFAIl+jvt3dh8O9m9CX4RLImo58/wLAt3JZJfv6XTuVC/ot04u1UPGIpU2
2p4zV2Dk1CNXPbI0A0zd06ommBYMR1QkAL7OGcZot+osHuFzz2FAu+XuY96dD9ADYK3P+Kx7Ylv5
tScGqSGtfRAZVdT64NTD/aOdaVO9AI7VziBoWcPHNxkC6v6H/kKWspVUAcHJudR7NmyffNxA09mV
2j1fu5PmocHKxNk1a9JNzuLenjY0voaGdcrAUt4ot3ORSEpszonQGne141I9sghflbANzAuIjMog
rLj3z9gjtzgq6UKR78hRrN502CEHkulIHi1wq/Xb2wyVxv0TjaUsaMvCt8K1paRzJWFz0q/jDnAD
FDlChbWCHkecOnNKiisB2/mldtHHNBik20xru+HkBdeEu9rPv+ATdCwNfZ9Kb9NF7dXCxM2t/y0N
X9+7Vbt4W36VXd9wkGnBcdQTZoM/4O1qKBHjWzXCDoiR8RF5dEpbXT9jzLDyLDIwjo9GUFuLOq54
ftyq+r5e3Fw4OptohvbCqDY5f6xMlOkpn6FrrYQeuJ0Y/48sRMbTSOUToP6nN/5hi+JMY0QBMUSZ
m0/wzFT/7HO8ZZNXAE36azofeNgIM3/zP9xj/FQUw9/hV+4Tjb062kRnUX47S0DU2E5xfAMUd8WH
85wDktfz2O8vhwQuEVmoYME7WDCTxhyNqiqJaZOnsk4HW0EAie2dHyxzk6t2Cm6nN4FXD5mhTsNb
jophfTSE4IVDB0RZQzukrhJHGbHJqzS2E9gUyBKihf7ms8hhjPK967oRYl6mFv2GxlY+sglLavn6
NvLiMSUr8R+xlf1MpjrnyTOid23mcaqXyJSJwlb5umN0RBIkCJUYBzj+dcqjNyt54gP6VyN7x2EU
a6sJ9aBBKb53kyE+fNv/e/UFCSre/kbzbRgBGpRBqwnq7p3rkSuwt37ExnO5FZWBZSoUilWU2P+b
jjxI7IQyUnde8NqOcitNuOapDvdgHqtvr+ubIrsnUD+jP9xWLmPF3aFd8MVyN9UtCU4NI7craNsi
VQOtqOJQARD1cdoM5YigWpM7ldYZ08Rl5XpwTkcFQQNiQJkv1O73Rxe5o7ge+JApKBkmypQOzywP
cIcikl0g+fFzhuan5pyXzk3/WnhUf4z6gls52XXZcvBIypyRKySOGl7OMzDClVnLEKM9LEVpa5gk
HfgMnxDTATKzXtSyTsKwhL1WkQpuxTbpgWSdVcbwapvkZRhlDCK3vBWEj/Y3uIGUmppKi26vSUGG
uEC2sJCjP4imdLSHyC2Edlvc1+7W3CUtefkV9kn0RevlrMvASNFHi+yU5vnJ/AqP14hEBBBENU6t
j+SsfqT/zSTwC638MRLwbvviW8sWo5Q93m1FRoP4V5xyWHox0lnO7gvdaFQWZ7aIAbWQBr97nvsf
OcvWHNWn/7shN5dK2Lx5ppAjnG86RCKVO1OBSJ1p5L3oxA+bb6ZUgzG0UWw0E3Xbdksn+6JE5cA0
Yj1HOQHX7DmrwG0a84WvTNcpfrx3DxomI8aDQ6G5ZpBkKFYnPofeEkinKGRo7zX/JORVG8q0xgVP
OdgLhseFsCahf0qJn3PLwuPtzGTBYrJjHiNEtkNbMzt5DuNIXgo4kAb6jhA3pkd4tOyPr8sSTquO
ff5l+z8459G0yVLVQUS750lLpIt43U2XEIAAlhAUAblnLHJOMmaA+66kY5/Bla8H61KaCHoGiAph
SIB05M0yf4QzwqiqgaVN/7xMHGBSwagRcGORgO7c0aZHzOWbtwojiZt+sUPln/8FlN2IeQRmWRyp
Lqp93qCBLdMd7jws9vonYNzAk3qyZTgJPkGCMk7iJSSTZLHsqawv+AteJn4ltiIZG51MupJXNN79
+h+QT4vRbLjLPSI3iEDUxqILbrV3MbENkazmkN6AV2VGlXL5AwE1vxchiCCPB/aNYa5Wsyqfzpwy
fnl/Wn+G0IANK2Mjgfdw2teuUCdu+4eMcwKoX0nb9+VMlxgKIXj5Y2xIIQwEmLkuLZkqnmiofWeD
w844RjibyTdA/w6CVvOYRUjCQ0gd5WL+G+E7mI1mGyL8SNiP2cerTKZsfUM2Q0vpquC3DM+pokl3
ubt176Ch4VzA7xuRxCoY0XjK5x/5JMn0UaPgSVMuHUatbY1EAchQ2UV12dMicYq0D+TeJcjj8/fy
mPyyCTwI+GSiwCeadWIZ/hFS2vWqjCG0JwtLA/WpVDzxKhmvPx0gIZrUgc9WiWkMdyyQoxeEVYX7
vAuzidTq7BzX9Pu9pFqqxbKXIniznmdCoiz8qFWbk2TGzFIBblznwqt8QczeMIIXWf7Amr7qCZeo
tJcjoE0Ylfb0CAKNl+6diFn+tgCa4sH0Fma4WMt169LjN/+pEpd9F8HUQgZ/OUf0BF/HodaCTedq
556w5WXFkcpYKk3BKqV3d8CU5sMay62iIwdAAj53z+0LogrfmX/kNqFDDEcfvG9zoIxq7kmkQV06
/F0DnpQO8iYOWZmWQnMSkEGmVZIFKtzu49w4MPzlK7X+68nVyvJCEsUUzLcT1Ew5j6uiba4HX1nm
VmJ50snP4YkLiStIsQggSN6HwN/xKs0QEEMBzdHThCf1e6vp6HzzxBMvLOD+KwHQau0+BvWsqhTF
OMslgG7D8BHforDYCjjpZO5+cFvAfVhjYZWioJPOUmxDk2tk8taS0QJzBH0jDQMi4cWqCxVJuk3f
hE/5Nr41MGiNvoMd/WGhjr+/Q6ZLHuZsYFlTXtf1XO9toNe42Op2VuhuQUud2X+6tbUsJn6dElKu
j5WlULZxfO6K48ZWDeC3pmwmlONaUsMa9GYV4HWl5oOkg+RUkW/FLDV+eeInNzelEUkKvb64M74I
B8Wk2SFMeAXNQisi4hM2Xq5I1JA9EnEj4Dy+8lJ9TTpX5tJ+ume5bdtZ43etWwnS1d9xjgho0Wqn
gcLdOBd2afdwm9bQH1eYvIwxa0QAb6bc3ZzPHkJDyD49F+W8KTljW6SHoAkVUcNEYgOVH1zxxkVB
ELnmHLznm0rsx/rko9eHn/JuTkSM1+icqtf3RS2Sj2kzBc6nkLuqd7inWGxRpG8XBqCVntlJEfpA
I7QoEBraHVXTVjk952PwbiAvwse+irBEyphVajLNLOfPjM94SzNiIJQfDEBmNSP5BSIRE0jN4TLS
s10MATPlS6gGVYJ4QAyPLSP6ghmd2xMxNdFC4oDOZ8YUwjvp5E8SqBWrC0mXZ1v5IbKJNkHMnvAC
KlEBIcQQsZA/BxoXYZ7HeStovdz81vWUkPMBBl4QDaXbSp8mxkd6esubmq+GyqZzsDfkfglr2i6k
9p87ybzBdwUNfCO+IC7OEE4gI0F3TmgH+ljcqu2S7RbLOzefuik0hP6p6pcsFA3W8/UNAIZq+G2t
QDubC21/YdsOXrlKtHUh6YavcFrGN5g3jP2DgUOY7rgA/0AwE9XnNnVI1IIdSbiLcMfriEvMJGF7
tvvZTIqy/n6GK2jJhk7vEYlMQw7xnTAwI4pYGK25WBIaniXsjJ6bcl4Fq7gmsi9DOr4/+jBKpSNx
ywjE1m3eXiy185OyXyGzwYOozb/O6maO6r6kTYcmYkI5xprPaCTMegQgL3rnhO3cGlLogxx2scXk
RLR6sDF4nQtCuCHbfjQd9o5e9tBSV11B3gsQTUrtv/TShS+Swiue5SSzRXGsp0M/mAMZ2RTadOjS
2JQ6g4YROdGSSa0v3V6RdEWqSAGJpRwlu1iTsRjjKIZvPcZ/ZStRq8/BVkaUtr8cAhyELrZ453xy
z1wO44Ozdnl+vYIjZDOMRzmfvP4ulmYPOj5g8SBvY8/HnN6OvY99O3K3ooiSfSP03XmNP82b2Iun
LIbE8JGN8U82Zq+qxbA2kjcGH9U1z20cqVQb5DiG/Gq6ttSn8OMgCcnWzEcQnmNdDZ39VTBrjicX
rFFzAJDthUr1Eg7gx00ajm6D60KT9S3yH4kSaaKk5nJQfkwVVtxLq/KNCf4SgjoyUW9ppOmPkDi8
YeRMtz6WxR+yrn95aHrMq45l0XeEqjOqleooHNSKhvvoTGc4w/559ItUaqA07LDmqfGIdEUDErci
9Ak8nQQFjvrr7eA3TryOQhVyKO0iiAdxzv5fcS8kEeaz48luATR+Z/2vNmPQ7l2HLzvZ3boR9tQX
Vlq7hm08KvlfUDJ+Dpz8oxUu/JyXvY2gKuZNRcysNGKIuF4R2/qjyFTXfQpFUgDHdo/c4MhDg3DZ
z7BEiHs5JFBuUszTP7Z8AW4/VuNxpf/ZKCZ8kmhRtIoJTJFaey1IzYHGliUCb7Fvi1yaJunf84e8
3dKoNJ7J8Mf78TA1MWpsbVKsr5/wgVZOfAsrUG7JDq7ebJKQANBzxUB6uSdmu+iLkGQzuXRMESGT
ls9JcATfyEYzx5gNvbAwigj30dVZtqVwqJUKnPNNzie18GAS5rjm96GH7VXd5/QypnLulEJUanJF
Eu4YkVXWm0Dupc2SKy7q7zubWeGOrhmCI7YhRQBmF//O60m3bq4JNqJb+eVGhQdQqy78cIbFFEjv
TfHarkJ2XeD2MTwpn9V0/WYg4TCnRqE0JoM2eziPHorlhRlZWQNbuZOQ5r5rRvQVDAA0AGMML9Fm
cd6Q+eirG7KdhePuYBV2x7RUFjm4Gzxf2WF/nrcyfqbvK3EQl1b5k6sNN+R2B/xq2QBqI2tij8bc
pwXqSme4xJqS00aZbsG7fcCVWVgjZM6FnHQpypFnrgYG9kuXjrBQyBePqBBiM7eGwD4YYGX/ynV0
pfCYtmG/SsW249V2HSxGCFgjqyVHXX0vuCLr7+eA9+XL8atu2EQrDIgz6ta74LPaE5PaOgnXdIGr
EnwndJS1/Aoxlg1cK8gSKIPw1kYYfjSL73zvkwxMssTTGeEDrifgyozY3fnBGPPNIolNfPdrICc7
NaY9qN7Tgr+mM3HcHRK2SlWzlH5kySsARPkp7KoUS3CcRkGTpP0KjQypGOjSw0UqOCIyb+FDW6dO
nAFrEg3Jm/rKdzoBO44A3g5uoKq8M6JkbYTg8CS0mBePSgdkMvtSCN1xL1Bv4z8Caqg9ErjDPvfy
7rtWKiO3b5EeNcmcYXqqNpQLRoifCdydXjjKTqBW2h14fkh9IwaDuTHVbkvPcGnmIKog+rFatlUS
ZmzQdkTrIQhioQ0ycPVf95dzQVHPSPvb5HUF4H/QOz4LZ8Vpyc4G5lRDMkXVeUb8xWXlo3CuHr0l
QAquWjkvjf628/AX6IqHcRwqChqUWH/izFv6UU3VeMLuYgUs7RMBV+yHxzheCQRGYiK5f7J1ot9K
QMZPVo2haN8G07Xa6tjU2FK2sfACatOR+JF13eYK3qZc+628g6cRJvslIPXblUkpq8BNp+s6s30e
gmcUD9RK+po2tMQufvNaiqSJj0RsvLvpLXlg9v1P6vTdJC8p4CmfarJUXOh9wQmtKmUqi9cce9wo
4cX4h3APSPJojXsuQ606vTV1pHNYf+VyLcxagA+jB5/t3mW+uQ8R0GAesIxOYnwqzDo+vTQtG48J
+FOIlqFkGE2cnQ96ioc+f8PEUwEWRRoZ9ST1TzTwJckPTtTFOu+Yx7DG3Uy3WS61o2GaYYXAvh4O
SKjOXVSg/Elh8HEc1kDvwyLjQjQ12MauDKk29dvIvsz4cO/iN5KY476Xp9Q3QViZtWmSSBjwfepx
kwnzMLGV5srOeRqBJ4LIPVoPmxMvVTaG2f7254FJFwO7XoSK/FGm3YM36NKP2OtfGN/NEf1oFoYU
fvHDXXeQMTqWoBvblf7mq04pvKnIFZUl71JqJwSAY8UpMLu2BRJHR27YJeI/G75jVB0QtUXP5ntY
HTGj0DGbs32sn896d/BFMEKlhHp2lC2DoOI1nhaNLvbEwlMNr4t4qkhTNMLERksoFkTHON4gZUT2
90DQKTdeVf6eGcrhzRtRlJUSiwfMiPG4Bo5HmKSqZRtofBi3AmboVd+D4H+8UKtHdgukBBfoz04e
usUKNBBnIWVQ44YSGYkywv3kDONbs5/b3IP0BD4iSIo/OldDrYF2XkBOG+ALsxnVjPOtBUO8BOdl
KLaXIc41aAU5yZvydUq2CS7ibujvW0+TneK3WOIzdrXgXo8tMuNm0AZtzTQlhYc+Hjt2USrRVchY
raqmZxgT4WbWXWpdvfTZdJokJUskQVdUUbFNDvGhDbxIj99iSY7xaoMi655gdIF/Yb/Cf8VDxTGN
ykZDjb0j3CjynpQrKMGoKMDThLyJMB8NzOm5t+J28xDXfIcwjAw3DxbLlptuN2ikqeXNAzsf7K4h
jMq1JjuwYIdXawbSAk9x5fuUK5WMNj18aaiE+Wi3e4xzgeFwGlwgqj9bZC9C90tyend5JJVgfQPw
MpNM2aev3qP6BQUeb4ZlhExwJQQifSoJpkAN0CldhgfT4UxrZlUkoMP4PqnEEXXTsAICwtG0gj9y
vEYbf3Ad5fm0hScJNdDBWxC9XAplHhi9WRlT2u5Pk4oDWY3alUEEhRTQT/7+btV0ZXdQ8vSDN5Rv
IMIa6hgg4BJZoEIL3zHgZhpclcvcdAcylM6RG+eAvF03eV4WB7bGzhXavZoRUr6Gz7u63n7D6Xsx
QI9bTF9j1GSbzZoXICxF1uvm+EKq0Fyh5dWeUhgf4eaSjlfZOs3fHYHF5dAPUdCGOJ4YhzLoiKpF
8c8+0zBIadE67as7YHFLYXP8kzwdRYGW+x0dMG+LzpQUxKTFUdIBE4D8+Al4bCq2V8pPfhkIxDQu
9A+4ZU6ufhyQpyJpDLhvNzU1LNt+Gz8EL05SOzrFbSv8afDPs2vgjWb4Eq55tQQrJj5I1M22MG91
IBlfEa3CaIvuzR/ZDQC1Y8T/Al1roXcrGn5I8zl0k7S3EAP0N6f+6H7e6G4xJ8IVFGpj6lpoL5Rx
PgIRuiPZDpvatoW4/MAlVUEDbSrnFXVlP6iKuaBYCTV/hHZB3V3IMWEk/uxfFS5gSe72Xfa1ZOEw
dS8EvGcuwCwRndHfPFoPCfK77VZMSaKPFd8mT06KvRZYCHfWstNsoSIDVU0Qa1KDss5TqO5BmGtI
RS1MmpIbJCIMfH8AHbhNhP2agmfrqAo2QrK9ly2nB8HFhZkZVdEjH1w6CMQguFMqy8UAHhCfOSeE
6UMSqPh5fkeOifDUh29FZ3X3LbOLte1BipHWNUIONogefMJKkEiqM/Ba7D4ybmBLd5xKVSdY+G6d
mhxkl4DIM5O/ECXhZCSVxqswLRIJsas0aCtZ0CXpVUiSVjtG/w16zfKNUZYadweKO3/gFQHiFI6h
sVNeuxNOPsIpNKnbzklqKLp6zvIpP3thT/XNAcDm3I2El7gxIBivlR3V4Oa/MK5oVgspBzBuEkJV
6utTHXiETlZPqO2SlTaockgzXS3CZr/O5nDq/0j7ZxPsbkIOav/fjVa+IYf0VOrhB7OPkrZGsqYI
wydV4hJ0qcPICL4uijmr1VUsaF7Lw9i8iIrx4foNBS6dTkLMBkQM7jpjBvMSJ781HgfLJwHjTJ25
ua5jZ/M1TCbE/cVR4UWs4vq4/QVlk/MOFpO3SxtiHYlyI23Kx19rb7ctEqxfja5c4uO0MDhATVHw
5nt5fDKb4YjW+Whup26otFvYBg2uiLSN98CZDoFCjiNrJ9CcjS0D7kgzs8hcG9V3tW1eZoszJSTo
LQoxruvu+QRF1qJlJHeUFL5RtmrLjHaXnuIagc+5ZNgbnjG/qfHidIWaKpTf6oNBsyem3phKUqD/
Dnb1p0JO5KO4cnUnwL/ODDS8dWVCRshc/tXuybLePkWTWzrLw2mDeZ6W75e84TnW3tZEFLwZtrec
B+E/ciH1d3cvaBcnP8TSueO/lcY7RwoRsV+5BIExa/rfmIsXxTAB4l0lXX/Q3R3Ijd4CQZv7q0IP
PTjvCJDlCO/hqp+BkLoO9N+zBAwPY+y91LLsI3r1I0IidfJbO/c7lRCdDZOiCFo4q2lbR57ahr4N
hRKDcQWj1hjTDNf8a8xXUBo8AxjiURKyKRlzco6hjevQ73a/n9Hm67HnXpskEX++vb6UOwCa1i9V
1R6O7YgVvYBXOTjSj7sBJpDELM7/YtCa9QNZXKWoNBIIMVmhNokJgyVHbNAM50OzyLrirJWC5Xmk
yJApqb2o5DN3LCgGD7tTaJI5DmdScQjRx8vPCszHqoTDrFeCjqbvJohEpqQo1R+06x3MZxrBIg+a
nqNDdalA/15C6IjyF43V/UHRz3or4FdCLn9axZ4QpTKWdkLTm6F2WWZf8sIpeeDlcThI0vl1NFHJ
Ja6lHDSoT5BZwiZDtKA0LQjgWyYk6jr8X8m7FzAjnA070EFQFchZ7Se7/U7WbrGxMa1HvCPunTGN
XfQDflTThmICwUW4NHdN/xOFaZP8v/xDN/07fqqxijrKpkI4WKkEHK/oxvdmrKz0yCP80usa1Jd4
8XP0XY9VnjR7wwab31bg2Uhj0S+ZEHBHDwcbwDTu3I7xXYplG19/rFRSrwjpoCy9q3oD11UUJ5Pw
dV5utlGU3fkMQAJ53cY1EUGeEyoOdgSlyWUBrJXVqIaJ9OQ+GS96oAMLv6TmQ1Ss2xW2MVOsVIZx
TsETkzRI2EdCJ8qdtAtEJzoIlesgOY+v/lGg+sk3Fmg0XBsgE6zOUiCl9nWhbvxvFOy31WDvraC7
0gNlQwYb7AsOVmZoGNn3xJVBtL/xRsdlVeAMgl8ZG+yJTEZ6Z7D+BAqwC2qpIJeYgImlCOflyWxC
20NX5aRmIs9xsn4PrRBdPZqBcP5PiU/m5Pxek7UeeVaipDQpgykXcoitFO28OgWKqyCHuP+g7W9V
x87v2IVRjAcoousgxK1/cnjTtJbxc2h/sQko8vzksGWk2dyAHKCnDcKR20zWed0v2tfNAPIqsCHW
+8fLpgUoTMF/0h/E5scATdUkaSbw64rkMXAYmh4qN4uYsK3vRoK9iTxfgbxj3IxV+e/fUuPA0ELw
IgsIcqej5pxv+DZ3effxmlfaXwMkZctOrR6ygM9tRT3AtFHZ4cibJNwhcNFKVeP8yiqq/l5tkUgh
M0366DvGQTDjzxTMcfYnmx6EU1TuHBJHFc1JzZWBAqxL0euAyuh+xseDKI4fiu8ibPtz3JReQu5u
DDiqTZnRV/SH5QZLDax2XHIMPbivG8/+0kPMRRpJgb9erJq4Vu4wGDuCaytbMJOd1fQXEnjRVPCc
8SRvOGGmvbABSVxMtA+o+9zpcUo1/q7Q2rDnGZ4gBxYbawxPomGvaOQAwFZwil1xy9u5BAmO48f+
lNU1C8u9fQA7zhv2W7P8nCMY/IyyxXFDIgqwttqHZnxAURC1F0Ay12sz4+Qs6uMeFwwwfZdOk3Wy
Xu2nAJg7JEZDcfcbF5tqZ9Cw9HEKDEq+Lv3ZyMufxr00oQWUTKynkE0l7PDRiSidjvnJq1OlbbjY
grO4D9dTf5sQoj702qWdA2gLfhx1K2vDOd7q9wU+0FNyo5EbTR0nQC43Z6etBxPMOKWfKHGyS1VF
pvwn2UbDG9vSksSdkNrKm4jvXe9/ayTfKUchwVujDOSe6WqhfUVNofaEb5phARrKdumXCTxXIQup
7s3dTyRi6918/N+KO4n0zBUrsUseT02D6Ys50fbXbBglYfmrgylj6Sd50MGp7xZbj/N5XVTqmg2t
uel4afKr+n1B8KQqN9jOxyVnedyVW/gUShUrqUEl9Gf+4r6Qv2V1W7GFFRm35dJOJYZ3bDaT4db2
sLxcWRo8amopFFywp7mv8+Vok0D7TVTMf3O+8yX7Gr/j3pt7VkvFdCswrHr4U6l6iFHKPCE+Zm3M
1AYbGeGSU7BQDeBtreqjqARMOaSr3f46v+Slj94h+PAWD8dE1PopuGUS2gq+eyU0PwXMb8AmJEyg
f+ikwQL6qcD+LaI5svXIfPYVxIM4bqDzl/6A0Fd6ID1XDVOivw+VdDLWTPri+1iKLTSBQQGIZKam
VSP3kf0GCi+CQnnxUPHjGuQBt1DpAlloQJjmam6/0B0Uw9RekRwRAU9X0bgskyiGxnfO1Ml6kWiV
sgKIDVBRAkspo65OWyfZxmXkhkisfps/bYDfebQGSTb97u51DFLhpl33SN4XudYXyZO+4Ni95tRL
PJtlCtnlj3g8g3yZlvHUSdPjBjoCUt4DUCRrEVplD0IiBu5+NpqvjMlt9KY/Jt8/9+ssr6paqzXd
Q+G/GcAdhE012sgRB+hiG32aLOvV9YPymbC4KCIZcd9l8fgPelM3NnSn3g7wJNvfeA5HxDSCKXpP
ngaiPSXsdMxMAJMpgUZsyV/x+gP6vp8OFWbBbeWiRSMg2CjmCcFGRqPFEVBn8fVT1/dcouxtZkzQ
JG2nlIGh00JuorIJijl0z4c6r+rdB+NDTIEkNxARs0oyvlhiqJsl42NdM39T6vzsp1T/VVZ3oWls
8l9B8Ftsd4TvYRwOU/PFjvDfUfvA0jmoIHwlDyxohKDpI6yJmV4Z0wvGEgDFHMkbSk2+QmrD8ZQh
t19vs+d+NTW+UYPJExBantWfjUClZj1dPc+eb7dIPMYWtgfuGeRWaMPErHTZg7wLbDDfswHrUNJo
+LCMQ4YI+akhpgXfNbR+CKszH5IUYmy1P2woyjdero3AECyVocr1DrvZvM+vhRsWvNvsElNo6d52
acv44h/3NPHFL5VonZ4Rb0pUztXOdXFJ637kcHUyUMaVOvzcO4Gd2E6837TSHzY0FvPkOt6y1HDk
rRXrpKJT3u0zuvy0ef92us7meezo68VT8iqw1ps3RzpFDi1DN6nNfEScti//VILpTuJk3AP/oGcE
/Lkc0ahMBQw7/Xf05WJ84RyNFdpxzaACgM2v1SOwWfybKvTltUreqjCeQHqmvhPlJH648gZpAYxc
5lft7h4wx4di4MGTy9JF+QffnjUXrEhDS7ipbOPoFo3dNE7lwLPEh+Pjx7CpyltCT2TLrRt+lWO+
EVVyYL05tk8Or/Vnze59MQuYV2z9sc0ca3TMjrOL7RtVWbCDSjemxX8bC896r6OrEdktbzZjL+/I
/EDM1lwO20tNdzvhxm1qC2SDe2iVpG+62UQJQY5DCmRvh9XIl28/TxsQKul4+AShm3NuwK2kisEN
Arxwz6IhMAZONFbac5X2JidqOru0WkECt+BBzrQuXCxx382KEMkrSuEehkQq6nJXvnc2nCfzOU3/
Vk0YyvMoaUaUOrzhqKXnKD9ued9AEgkuDuhRHu9O9sGS4CIu8QEq+/KOJn5HAHpyyLQCBXBcSjBY
Zi15PWsBtysiLy1NMlTcU0C4nmV/uzd+OEnZHjSEbJDN/qaTZRlp038jTdwwttBCCmQnkXEytSrM
vOq9QaIddSnMvkNsbxuboh0JUMtuVZqGdPbPsv9ijxdinLDtRW0edGirwLvXfKewq6/nF3G4QdGE
YxXbM3v/m1lcEYeMG5BI4t1RKQx6kcRA7KQl2XpmCaEo7BdaTU66BlmjpM+v6InVmWFXM4fhqUQ5
ztNuBKmLgD2x7eQfcg0M84PGVLZdXJ1uko6MJVUER8LTC8r1UEPZujLVJlTpUyBgQIn9l+mvO4r+
6JFBqPGFAdX0623zmPrGbsE/Uv5fhoxupVO5c634sl7kdYru5PozatmryyK54vYZ7ssvS9SBFZ7w
YL9MrisPiwF2XeNOLI+S8Ae/NyND8Zko8BZHaIe936varpIll0je6ZTn5Ibv8/e4v0UvYS/4j8tq
Yw6AZ/Gcac1GIiqCdn6XgL6La6QM9KXF3mj04IK1ylMZl69y4lXwZLzBcCKfdkF/mvTVZP+oty/h
pR9Zz7DepscztrCqcENN9F75qefcJjhY6M89C/MTkHSFKh2tnx1MldPWZwtvyH9R1Apm7HYzrzYV
rwICDrmo1wmSupOfGHjWLifLmVgr6Ijdo/kyxqTqPKKyuNcbxq8Tdse9+NnL1slKlUvD42NdnxcY
sR/MqapcfEgMA+Mgwc1IXNCVsA6TD/28RcqVSAFhoZk4Lg8vhkbUiAEmY7Y+WaYj/YJspIb5yWim
yj/9qCuy7EpcEcb1zUDno0PBCWbSRdJkAhUCNd0ya2tqmeuRCAdDq2ILyU+QIWYjX25LofwgeNFB
z5U+KgNMhdbfobtucvda4YuyEz1NLXHngDP5oRTD/JdHC/AdQddWMRrSJdcqe0SP5M/att4Ls8rZ
vhChWIzHk4PyJtVHzMDHLhXEj2XQA2o0w0cpXC0Ak9Xk7gDgw7AT2zZkMv2OkWJCu16A6fA0R0A0
+IX7EGHS3jtuDK1X2x9V8SZsjKloJruA9MftKmnpRSNtj1EIa9P546OB6SPNGbYOI4PdaVPzvGdl
8oLjOJWDOe3QTpoKJdEM93YI2Dl5cnDQjsDh8PPrdA8k/kfZzc2u6K5fgn9QtQnnwtJ1tY4IrOnG
3TCZh4P9yVXzxOyqUFnYhzLzdmHlPjHah8UgEmNgU/K5VDUUyKBeE3DEAoijtwpfUXTuNHJjHPHC
fNSgywgRu4TiI18OvLTrFDi9ZUTuXuoGeWo8Xja/sWEbAN229OuJP9rY9nulyQk+OzpKJ1rRmrX6
WDjLe/9FV4KoGZbUzZI6jU+YsxIMnSSsDt67KYlvukG5utKOLUu0Eb/hKB09rPoT5bkcL+xhUGAe
dAa5KM0CNRVKHFo9cPiqsX5UsPmap+8P2cl1nkExM3kG/DYz83eKSdvTsromz7b7b7Ao7CCX2b/q
BbN0zscjbFUWgcyspZ5SHoI046cUDbXWa/c65WJGddLwApUD/Ir8tRLhv5Gu26T2/cpQOcpgI1Gu
rq3ClpwPtQzVR1mbyUKutOd/Ctb+imZEjWi1agf5K4E2iJ5rm5/IMg5mxFsTBrTmafea8ukxmTGq
AFTVDuM4CTZxFPOZKki7YFDHWS1YdudplMFNAm1jKcW+Pv4XKPYpKux3BLG6J9apgFPnc0P2lD35
74G3YMvRW7usvijoVU/1SYROUr/6AKypbqSRqDbRHN3wi+pdcIDC7AhglTrNukNH5AyHu9tlxGpH
1v+XecCzoSU8o6OgzbuWhTZBYVgtv0EBEKl4CAx6RdVGQVj7m8Zx2Ni0LWrTu6dA2WIhwbXC4xiW
gTlNM17zEDZ7rPoei7Vv9tChbjqPw/kvZBjxSVZHLBKfNcnqHJeJcXHmwGjPZ8rKBT8UMnGlXP2h
NcX3Q/jIqVLqzgKcjUQQP6DHz8Mc1TtTWmwJJz06WyT/vw8/C5KUqYgYnhBgiQrCPeqnZQRNYOJl
vPtPV8f1UravpkELqM0nK5rvU19L6WF6DEIndrOj7ntaHNso+946pAX4TGrRYBCOUdom3MH23f9b
i2nDWZQEDg8yoQq44vKyLQMot0hwKx2SaTKeZnCPzhSmtvePjUa25sU1fWsjLvtA5B+RLgvWlOWZ
5QjQQZrdrUcd01f6lGUWiecU+SupPbhtClFmMhl/zQ6QIu4JIY+3zs2dyywdwVSZIguMbxD4PSCR
wEz4d+ZTvTLyoXmP5PNWlyxz4qILNlsh6rNZnyX408cWk41HiEE1ZwXo7kEX/UxyCXU917AdWc47
+hZT1WPrnovPr1fUa1vqWb+sgfqP98o272QHs9Rb9IdZ0dyP+l2yxo4IfP3Y2dx3cj+E6rj+UrL9
NZ3H/Q4BiDfLY/0Fck5QRYRXbAJW9OmClZySBpquEPPZHipseJ/Cw7jqWHrQIYIbj98om118nh/E
lRmVftVdqITNQLmf9vDsr1QhLluL2mHebaI8H8picSUPk6QHKRforUBQfeke4ACwEKAvbbNYnvtP
jzHZgIldXn6k8bhkfErQhM/bBRgJdeIb4LcU9XIKUT9HDOMcoI5bYw/1fYKTXdijSpfKZQ7ulBXI
5mp5QKsQHbETC2PGjhtNQtf4jXG7cjR3MJtD2WIh3QHkbuVmjB2hdGa6gaQ1tJto8XpOtI42yzXL
02XyVC6yqiqOQyCs4UsthMf5CvpmshRDp2ejRvNLi88wK58zK8ioopQ3BuXLy1/wCe8v4NCVY27H
AlKaKGhCt14I8fmEaIAyb+ORgX7LiPNY5IeWqgql3URSo97bFxOLM6mEY7yVTKMfrcFajONRYs3N
3inwjIaOneEAgXfsBnFFbR7N9Krg+5T29qOUpvpWVRlFTcjHe60Q77+kZs3h/htam8gG6PUMfl+b
HsUohbu5NSU+C/LwwsmAIbBylWzW7hhy6P3yXTGdfsCIqPrEQ6yL4/G7y5akwkzJWVb+vFN3hep1
3lW3P0bIhlh3Z9QzN+m+Ux/PT8+dx8F3Jrpi7yHdpOKc9IxEKh00HNiIL5+KilCP+SsTWiKVzfBQ
22p73LzBrEmaNNfDeDiYPsDH8zCnfYXeAe3S7vvBUgdTeHzniJryKiPFvSAqcDBQI8qf54swZVi6
T3stG2hTVkfjcRc9l+ljO0x2xaVohJetSSaORFJqoSkvFQWiWlKEFyFogMI/VwMU7/n1fkJC+dO4
n4PbDvPW2jHK3zaPrCproMYJCKHGWKorIEIypMVpjdQLzCV3adQ26JB4aXMNZ3hVHcsvb/gB4QDU
y87SG88zIbd7T5Qie/aBlKTvuYFcmMBiEG4U5mW4eNQgK5+hID+wWl3D4sVsSPk69FEsWWgk9Ux7
fVGZz7EPTpvicXg+bi6RYJIJWnzWJEqr6F7xl+KvlK+Vn0T/oiZEDARXRVC/gPeuJS1AumXNsmOp
c0EUsGc20AM+gm2ySQ5bmiQjgtrGeehCYdfIS/NzjCKJ2x5BSL4M3ff4rFYIpTohZK9B8mbwYgxT
fmB8Gg8krmmbBEyljsTd/r4ozq4s6MqYe3AytjXMKj4+fcHXG6OTkXXJGD0/SB3KBMUVjAzkFBAx
Flplg2ApT2BFZWbjQ8Dmthw7bhp5B8f0NLRK6TohFbO6lud0UbuQSNIpdJw0OtN8eD90PQaZECSB
2OaA5QIzgGHXa0U32q8NDjmZniD5hNtaeBFZAOLgPSYYL1SrD/9TFwz4GkB7X0QHwsUSsguUaZc/
cx8ulAejH1E5L4Xs3tdszYrfSktBODIaR+kj4U6VECn8o8JFwRPkxZ622uvEcCHt3SooDjrRrLZS
Edj5pdOin9kmqmkFfzbO7KN9g/zxfLPn1JCkjxkEa6zc0N4KDPe0cgigP2/C8LPvTcGdnfwjshUy
uqL77Ebeq6U70otitR4iZiK8tkURfjmiFmjJigJDbViwcbv8SW32swKa07dnqtqc7mjHWDTWIIEn
bfVwdgwDldfIZouZn/wLrpr253Zb8mLf+hizq0pJ5B5REPzjLMTsMjMWSozXZsv9ZrH9YqgwBfgB
JWND/2X+AkyYjRVJyP9dasZQp7ZSP1pcFf5fWThiz/yEFl1+ks3qu2MN/RIpHdH3+cOOlGWCgpxx
Rk2IPedUCjsLK2USHDaATQ1MaaCR1CoUxxS1Hy4lJhMMxu9wreQMj3gWr8PBU5yba6uIGXHcDDRE
oUYUC5LM86awn0PAN7nGaEodGpR7n7olYqvKQRTNxl+oC2Y1a4V3wVVOPGRCyNZ6/IDGA9nyPdhp
jML7s18HUu2IMPKk1x7NvG5qOLRAZoEd2auSzBC+KB9W6gleIaEIqWPGuo2GSZzoN3g1Nv/zGEj9
/sTTPe6CxYKqq3fzVf+KHcbZAA1o0u7hwXlmoWyucmwFCz7IB+p69P17AxieM9M3cJydx31fDLNi
OD70Fzn9WmgKm/Q+dykakNhXqb3vCUxNzPG3A/Wct1+Vrh5XgzuWtd6XssehS/6K5vdscQKcVsCg
4ilUy18NMJwhd6bQdrC+RYJnivCFj9GQ6aV93uPn6HUdUTu/NvaxLVkMjxrD4gvoquOqr6RZHIRa
JlwDhEDgxlVLz5OQY8XpXebQbXi9gypWNUfSNjnA0Dnike/A+1bII0QYuxokT8mPRdepyacIMPsJ
0qxr91DguJjgdmnfiAiwDW0AgFQRzYp2pxbu1pzNvf/o/juerJDO0J8aifuUTCXsfKcx9F57VLJ6
zCEpmseHfzYELyP8DWSOFzuZbM8Tt9uFKKdcwFP6qN1kxsq+Fuc6Ox6sf39W72mkG82D7pvXztmd
04f2F3S1iS+GAfwxpO1OMSYXxcdATKjcVwRJhFBL0+yMCrjRC6CvKMEFRE5XO88p+/+nVS4cx9rg
Dz7qX00mDg2szVWSZ0VpTW5ZjMSD3VEYyYP80rOEfiJIF9kxN6DDsERtAQLTFl8PxJ+T/MamE5rj
3f+uYIBk8+yxG/WUm2IXamU/gbBeJxHcw45gex+HzTV2fV1yHiNsRaxxjst1oaH/PVQxdGDThsQA
5j3kcZhJ+CwzmkzQV4m82ruuvAgreJ+jSOQ8lndNvjHAvzQ1pwkAzB1C2t6Pxv2AZNOuIzSgbDeA
seX7YeNa0nB2K/kI81hmqLP7il1MSb2K6oftpDWN/9CTWoBc2ZAy/qLedkj5tZthBlM/8KRXqcL0
64XtC1PLdppY25Sjdgqd7gNWAwfjr+HPKSB38+tHJOmO5CpKbQT28X1wMzsqlMomxyKtfjTGfIzj
SN+D2cZHU+IKAlwgiPTrqH3w8BhDYBB3Z0kzUoVRjmQHdyyUVDENGsibSck27aG9H7XZOEBrYgMm
sCLGFPYXWSOzjFzEdd5pp6v64ic1jc9mM7KcNdX2UYQ/cNhDZZvPfvHoNq2mxe+SaVLX21K1382H
d1r88ElRuev+I7R/Bs4/5JWbpflmPAy4rym4EGAPWrpuBM/Kd8IDqtOPT4qThZZ3Fr7GAzUSXzl9
CnMYX47gx+UF3c2NObsVLH1w1FCgWGVqL9Tb3Pqh4O8t3SYy1w+JyKZ19rZG4LgXRPh6IoiWO4cg
5oZNzfc5GMtXZOUlfhSk1xVuJPr7Ydn9VGp57GlPzAElqoB1YEYeQWkqCvBos2mO5HrmKfJPPyIE
eC+GuoJDmcFnT/sqPxkE7e89P1BdmGI6Aao+2oZ9pwlwY1+DPaP8GUpjGb0h23i1PIRCjBJJWJXS
WwvMaflBntaJR57TLbDdMw2IP9JlIT16+dwNW1TZFiYngw6/C0dyWJ1KOR9azfURgfKfF4mvyePV
HqdRobMpEIAntxwPZ6jFEigSvPcRqIRzG8lsauWVuJbFVal3V/UTp1Q3507bM434hhv9pRlC7jUU
QtzgocLKkWo4GcAaXApyySrHHPAwbzGHqutKmTAX79tCJXlXBQQmGPBZqcMaNb4X4l8T4bBb9at1
/ohUcmCg3lawHOI43gO0wUTSY9apjBGM72J37JNUsxmKTdWorxLepyj4ruEfA7UjHrL2w8UUwAUG
4bdgaZw6DcR6tW0+x8scdmgOLZaEH8gMjM6hRSUvimTQCQehsE+Coqwh/f4W+ggnUNeDUUfgXRWW
SEOqNPPJBQziuaYMB5ASIb6Kd9Omn51sm6VHhcbCabWbqe97URZxnr5q36K00qoBcRFa+Wd2HzHN
EzOss4eJFwwfS95Xl8r3QY5P6YZQ0+vpHYgrITRrPQhA1dQFQOVifDZUS0tu2nDgsPkW4G1qjJu3
m+odtXEggXjlziILMl3/UAaUqTDrb7rT9FSBnuk05yVycmeLQyC4BJjXeiebqDqeL6f0DMjiPlLj
Y8RxNi5gL/mL5JQFMLmNfDiJMYLHKVRXer6TfaUjBe8bsg820VYcLrLj5ACY8p0Y5HRy2mb1DdU9
/OtRF66Z75rXh1dzeP9REmqtGh/tBzSOZ5WWnci+OF9ocBdbHW8e1Jl7RFj4hwJdsYRWRCa2jdvF
B/BrrW0CdX0dRAY8qFnQm5AlCAiRqgc4SgbPYjPIRmYtwTF3EZPb0byYc2bnK1A732NfP9C056ZW
EsHmU1by5i+Eenip6qu+v63/YJthXYLqEgfmzPE7s/SYuVRB4jXK3CcOCp5oq0LJTBUYZvdA2NHk
ESn5i1/NWlpslYuG00uUP/lvRxFvZBgGz8bves22AzIB1sgrPTerMiKogM+zgbJ9+aXz1rU1TaR3
8d//lPPSrkgGog+iWuG17Ie/VfM/hUPbjvG2OSFU9hHIAexF9ZHEGD6miVl004rHxDMDxY2sck3n
wuNl/TXOcUhPdZn6VdOE79reNBxf+8oCKS95o/EFGrjVYDHMxr+BFHyu2GqBV+PmDV/tpG/DpnEc
asnqDI7tpiSUzjWBxTHDrx2WvnafvV+9fnU/M5QdoSYPV3UYPjKjqSi2G1rlU9XfxfHBJG9DrMZw
oCBLrcbTG+8yy22vX6wic8pFh82qUZRyl/KUAXpXm+ulxFugh2b3Db1cp+xz2HsKacrrD92pgrqb
lJiAvxLk7h/Hj6apmk/3BsE60A+EyfAhXpXhvfxnzYfUTz1l1ejyjYLoCy2TmxfJGPdaeTz3VXt2
OBqCqNcAwT/4iCZWDfk74G81jQ/ShQNihk9QP18NxfkpT+dbx/pcR5pxwV8QG3fl4ASUQUIgb1C4
XdhcvSZx4MdvycKhTCDmlixwCTxwnJSfEoMFfnd/Zwhc/Qh90BUDCoS1abZJk+D6EJH61mry/Zej
Lg6QoEcN07iFjgH4JWaNTJym0x9Fx+K+LVvtPWeap01XjZMZy5GzPRCb+SqVZNQu6UwRqRAF18kV
ELt6U3Qua18uyrrlJOLDZGMnb42P5m4U+lkoheKjuvOr7W+27w+oQal+WuOGQmx6lOyNqj1gL2ms
IbAJaFAVEkx/eQOwxY0krMDkrBDfWBwsJivmRQuEScv9T6d3HXaxdDgCD/xVcIfmdmFPV5jUEaNg
qvklvBi3yEIyUZW/fMycxKyfNWuydXblExwSsybUyXsgAkQOcJxxssWpONjWvfRAqeupnU4wLdqO
XzhHEV+4SwYPGa3xIjt6PzBDStENsgW9J0GsjfCqt24pkrOLdZi9rKat5W22Fs/yevubmfwIjh1S
oqmOmc73gEbby/DZDEqOT+n7QAmocX45c6jedezPgKZh0G/6t8T+kuJGo4wzbZX88BsjQ6RxQDD/
c51E4zo2ERCyL7TsaGnCItARPw2SoTqxAydgFeTVSB7XRUhmV+HUmYd87DRGvUVZRFGF3j4jQMiT
qKK98Qet+saoSnJqlN7dy/yM9PRCq45Rl89NZHmc7lsV+aVYrLcecwlv8594af8/NpHYyAKeiVOS
JVMfssRPcgRtEVl2Bt0z//zbA09ZTmgDq6FlxjBHfH2a6H8AzqEylmch64b43aIuZ6fLpNKbf5yd
qh1wOtyCfEsbeR/WqRPhcusa7+24kaKP0Iasxf5sjpdJBdxv9hrarVMaKBerWFCavRsU918ejAq1
Jza4m6nTkdr+xncMqenzFupW6FRWvuqWr9iHVTN4k5PIQHPnvLYge8q75Iqk3NbqC8l9O/ciNDV7
tGmXW9+NHCjHotx1fmg9LT2QuOzqx/zl5XwGR03lCXRzfgUYBtLtQR5hqhGd9f5vtXB5r7DtnjIo
4ukR2FUU+BbQvB/RBdVrAV8iDb2VPduMdO8KMdTvFV2n4cdEjXxHu9SrXwaFVajGbPgsRLC0Qonc
7T5AC9a0vW61FSJGYHjL0jODVJ3zAwNzX7y/HKTlSx1FqJk3g2hvb8mCiKxWiEXwx7tT0MaQ3CBJ
BmhTpuXk9RiUWxqu/pDcwIksx3RlK86sE2vGeFiTewgi+hE6k5efc3bLtxt+U7EU9DJ95S/N5r9C
INCAafdbPy6nK7MI6cKcANH32FgmVxL8ODA4xEYuqZBYQUPlJrKCbiGhuiBQtLvdP+Kzoy1HaZTR
vKifsDbzUSrW5TdsF+obKQDB5/qxE6kvC9c4aM0ttvQunp1kOz8yl0sV+W9FUVNTdTQtIkZOr3T9
IrmbEDZb2AUGfgF55VW52ZH0OuBR7fKIVgxVLajqSkJqPxqyjDUAFlqKKnvp2hcywwJzLlD+N8ty
whRb+TQBIhhAhbQBB1lTrpCSUGHgBEmAv4FyzMO0n2xNuw//6wqy8zm6Lf9eVUTZ50epYF/heOVd
i1+AUNmdXJq2sva0hJf8+q2PAvFHqpskFor0q/Xgi2v8Lj8gSqXjYZ06zmQm3c0cgpTIneIDtYBS
MXqBkpnffYakYY73hEXdhkbnOnZCEmoyasa3cDSsrgdDMyfvPooZ1JtyRUxtOH7IFwQmlH6nt0Yn
piCdWfsiUqO95LYFIFM1D1ucWHrofOhfnn9gdW2IRZir9n/K15622SyKDXfwb7yqXBkJYK7e5n5P
kkkJdGoN5NwGwIA7efAhpvXXkegXkxXTI4EeyDlfOcOP990S9yR9uhD/xqSoButlnFvwG3Smp+p/
50CcQYL4odDz4pf4YCIIVneNXUhFPLc+gPL/kge5KsmzfhxdI61ZzhHLCjbohim0wAwdOYLJ4r0v
bJS5zOvWJ3VbQCwI38opLwF+utLnI8ec8+7e4s6rXjiNTrVA2adZg6Gui8tLNOTvxs7pbriiWXAz
3jVxxLfcviCMxbaW+VfT3n+C68O0U/Mv1munDDbOv55S0uqO6+LmR/Np/fBV1ciGR46Je4jZRrUb
twK7zNW1Y+/HA6jggtrOZI7To8+Zqp0NCZ2RTP37fkk31l/g7ye6YcVFdk2Wh5c0DxMbH6fHhgZt
feJ3IVjfwZIriZL4IJZ6ix4TRtkIDc+g5gBKHVa/OsH+4BWUO5MJ/6BbT1TzqMB0MdR2YOoxQB2Y
ggVkhNWdoVS6QJlOngdIEnks0S3RaOELLHgmGS6IkyC/1Bs1wVGtxz9T7wSHK01JM7ITbjSVQTHZ
+AtAwxATR/PJsSdu/qmyoiW6AIws7gkfEDFd6RKsGaQlZYHcggls53jy7yUvQ+wbuCqF+hWy1VNA
1VEkQp5mlutjZ2KG94ovP4YqGo0lgF/rZmKMCPavRYJb1zjQ5AwGZu+yeyxBv3oOv3erABZzazyv
80PD051oTeM91AFwBLGRc6BEK1xDz78pr7QDgK90VpfAJME64S6C3YRBKVmVQWV52zYVGWLBIwa4
9R+lQep/+OuoUHgfbdO4CVSCdmAqJnYXOtSs8zZzEJjyQT9ZrZULw5r6V9nRS3QfcYK8AnOlMeqs
KK/Ejg0y/fpBCuFNTpvnzueI9Oovq7hKYXpgSeQcs1szH9CtFdF9bRIXnIYNuN8C2+hgNZXMm/In
cqklhvNxXicAjpzRhB6JbuvizHoAGDhlTADP2RhGkAIeGeGP3mhNEWhZl24MTcpU5qwIgCVIC/Y0
6d4yxdc6d3mhhZp9fZ88C+w4lnW5r6MY4BOPf4PP7O6lobjU6b9NcHFxG/vPs7e3sUD6k0n+FORx
szc2oikgyIhvijt3TXYfxhTZ5VB3o5GjqwWTWnEXbsMZ9ki10NYGKpPRZjNB1HjujtRsR97FHpM3
OXySHT+Q4ohj/wftJOjY8NRWZeREaPUDfzekZvJ6ps2yw9sZxNwuLaTRrqNbjBrJ06vMvgY3K45P
oQbAw8s6MLuqzhShMk28dbqBeGTZxZcRP7m49/0C+KSRUuDWSlEu8lJwQxcnVQn2O40J5H8XOsbF
GN1XJlcPw5EcI+ojb2Awyt9Ago8OWNFSP0mfyYL9zU835zGxD+7HYLgjjibeRyEiEZMUL7GOujxB
FP0WEFyZFES6RccJNSlEZ5rePbjLPacYJN8q5wWE+0v9hee+LMHXp64A17yAxDxu1dEsq6luUjbJ
F1uIqlgPthqyiOHlCl2QE6pxWPv3tsZZ1xu61rVofyUc2prMrbDiouC28Dj4tyRveTPQQdgGgLxo
zTz3hka7Qm9ZUykwI1AAW9TAqhHPDfESVVueBhdQkWlnsIHiroEoa/cexN5zM8Qbic/7vgSt35Ay
PRwX8zvF9w8dsYygqlaiO1ggJQV8tiaLB4Lomefp6RiNgEIADpuXdt8tdhsDAU9+YC+MNfWOjoEa
JTvW+hIZU3RcWk8NqMlPm/2h1vOxyxIAuiP57h4EpPVzXJglLz1ZFhF74OyMp8iCnzeOX6acLbrM
4N48lOMKol1213ObSsc7D4Wl+Z9e0W/YYB8iafc2t+5I06OqIVvafKYSP7pR90RmYGbcqY50Zx3K
xI39vevn1nCoMd5uYuISVbs2GKF0oNHwppuL6fHJlA4so9i/Eb9jTIPR/3/FYnH4E523FpJOiGXX
nX6kC8C9QA2R8E08eLLx/To+fa6H+KcnjvvI+tByf59YqDkaeyYaC/eVV5gVz5riDXPs+4H8/vfP
fN2vLdOjRQ5/3F4crZlvLb/zZwZwNUn4tu1SnfcpbuKq/ap2xjEkz3HZY7iwIEvDMLmcRRLnOyEo
fE3ShPJtJGV1tNwomqJAemlMbA7UDS8LJyCRcx+uckpF9H5/e6sDDSQQ2kqyDTQdvrV29oBxuMzR
iZtOdk1GvFfiAFXev6sjajUhxtS/4ARHXg9RlfMQs69sA/GluImpzHb7p7UHCYijmrq1YuMhjPcJ
lOUPu6jFqDqgVaUqQud8nPAD/ZiuCg9TgyUrXO59jbazrVObiBGdpSdpcgeFRNR9veLDIg4ZzMQ2
NE5QdlpRmCHEwxRCw9C8eAhwktocBprOLHyytmPLOHUsC5rW0uLPYDgjD0XQgLhuEyRcEsLUmhJQ
fng2bvQqUCKfR2+QZiGiIVfIW55p2E7UaWLim2dcMT8IVVNJ4WkI5MDlHcrelKwqW+ZGvX/RbsgI
YYhYP0Av6u16fD24cYElQVIXsZE9MAgpaZmxDJtPBKp50SH+FuaWe6bVBxUU9+rRWoDPb68HEjeU
CLnwF1rtkCaiYcdlFfW4CEj2aSU5NnVWz4sXeoVAXuTymidWS1G9xiOTGg8/2A2ENfS9VW6yBTHK
2dbmWBqS6UeDirE4JR/wHk2TcfANYOwWbVGADR2ese14+TzmvhPvZuvgEjyKi0tq2Zq4hAcKIFu9
VMBbyb4lNyXs2/+ycxp/0vhQesfz9mJIjnvu0YyWuyCbOkM2nkrFEutbYQWNLsAFmJ0NLIEWOT1u
TkXQwXN5GdYFYB/niMTk9/2Jcgv8Yg/bISQle+1ltW1oD3M+ZYUjBCkS+TiCWt6WHrB1ZtJpoXsg
tNQamY1mDxcGUPm2OefMJymmY2V5J9XaoldgMsp7MWlPBbbVXwZOOSAaWfg3IBnGee1p8Eyiyl93
+YPsFgyBd5Dt3BAjI0aC4sr7WWxc8xvccQYHf5Y6sTZQlmAB6+YzRFqsNxUHWqucixLKr9LfWDtw
3R7Mc8FVMxAPHod8T9vNEmyZbd7kwtDJQSTZ11QY2fH8U/MNLMCX3utN6KMnOW6rNyRIEpveWvr4
XVhsaMolMHlDjJ6KvShJCkbi2bmsEYFNhiNnh/CuV8JyffrzyZ2A4X98rwF1bgOSfVyZc+pQ3xcl
Kyd9TayHzvjUv6gdxFHGzXT+IUKfWywL7wzFGVVSt/T/LvEyHzRccrZ56EiypAurEsoP8SVx+63/
oIScsbUdg0roioFpo5O12iAb2SSHTbOTfisFJ9Vjrgv7IU/4zbeTwjYdy7Os+2VnIICWrKwoc5DF
Loq0Aja1OuMtdAiLppIk+clLsC+nzYpSFEFPi1DBON0I7Jdabh1CLyFXqnWfcdp5K81MH6yd+wZu
HzZDw8XtS+/lOKP6elzCw/mHnE6+vz4rb6ZMiZQysRiAtcAEdYsyZevziv0sAgwPwY5AAO9vy0oV
NLptBZp+1tczCf5TGegbMXrpgU1iJSpwe9jMsaV8//Cedhf0+P49bWoJAF6WNvC3hYcItPDEU8MJ
ZZBRfuio/3RC1WounXw2pqFBmWPzZW5diJgIDdpr6hi8uJVwTqztgLXGmgSmbnspEB/kVHyQ2I5o
mNTxg13wCS9bDnPxLRk1VUHjTcvHDd1SizYv2QE4GpI5CVIRZxRiv7lefQA1/QYCigl3GeoAOlad
6g0zTHXP6dPeRfpbyIXHeZ5bIIrUHve0fjsK6yEMZikENgggEaXxmw5cOJFbP3eZZEiUJjLBotOk
urb/VslXS2hPwN4ox7IXE0qZqsnXEsU50jR6kyTC0zRwz1mjeDOmHA6XIwGH4gy3GJHhNMRO968X
MKk/5YnP1rMjfVLyzCpXIFzUoNVcAyYKXcrz+miXKJFKad6RC/lF3SjvJ/0CwdrGMbaauMVShJjl
UAouaaHeqk3rg1SK7bXcfUgkwYjZ1lI+ZAiHAXDZwX8pDQBYMkuqpyFgc0SqC0KK+3/scs7pb/00
sMBiA5cLYP2kftVoqTcsDjqSLWLYvG6hrAT3K7iNQX+mwHJrPwuy+9FHZ6nXCNMCFiriM51ISP2b
HLuTzfGzrCDdjXil1UFVtn9gljHilSxZs6doL6SR7gixc8cZSVF0yDXWXwiFJVWYgIANTmu91cY3
O/p7spwPr20T/OpE6P5vRJY/Jo57hVzJcH6kj8XhAhszS7L0uxGlz7AyJNQ94sN9i/HhEulmkSve
OOck+nfIzVohtNI/oqckFYpT6vwiHLfOAXvlrsEFPeqtz0NUPokBw6g8m6VoS241/Bi/mrEQpm8G
2LABCRig0uYZmBYqZmnEgNOHRKoCxgj91OUEZV5NyFCgXMVau49DQotv9ZG3ghhmgA8kyh3yqfEn
rgdjAyf5A9Ykixb+Fqv+wPRAEFdkoFw9G90+WKhvKn3pyvb+iE5PDSqJuWq7hdN2FouKoMasPcpE
y4FV8ltw7sKWzL3YtSFbxa7Czonvo6PDUoqKWcrqDxaVbk6laIF55RlXtfq/KpEe4G7kHsCgrN3K
6uYeya3PKD4JeXFHxG2xDJU+SUzAEht0sN4YkNfH+y4HqvDRuWtyVJ1RA8xZNvF+8ruq+DOc68ma
WU6iUg3g5Q9ge75IFnQfB/2Cs/BVExPCReeSVg7PeELoTuGpgivR4xCV/2x3drKThx1ZdTebc2RG
NzEaYlFEy9Cn8F4Xr+O0RU7gZM76RCMepRRPwgFv+lUrwnVd3fl2UqbH9GC5dYGQ8aqxJo7ZX3ij
JjJh2veoyfCEEIyxd9FDtEresF6z4OkIfLimNYbyQ4zGgC9oUXURp3vgTMg1rTL+9iwhFtnQCTUR
zMHSh9mL5BQWFGCEeySi+qUzDniAXo54z1qVIvFTn8ZSP3N67LLNnTaKPgxoutQOumaedeuXYkq2
J3b5kb7IiAtuM7pTtZU7LMjQNN8vG/KoRbMAPn3jied0v2eD3PtBg5qr7AdmDhB4QoJWfTPDZcuS
3fADKcx3pAzzz/xQhMH2tpC5W8IN8se/X0d2IjxDvQTJOl2gglZwMerZKUjq4GdclI13H+6w7M/W
hV5DaDGxZN+Brh4Lw+5YwCioK/wBcxBJ/yjiu3CH1SrjOuq6BXWeXSw/icRj3XfNiQR6xwAjbCBS
nblvBP/MLOe9XXjjR5653QlSIykilOYfK9m8iNkPvV3g9AXDEOmiK3BPUfwtDeWe7RuLaKrVMC8S
pULRSp2ynEMvCuTikSzd7OJiTdVhXnh7E0UE1CXVLFpFPbxktCqotm2759DMpxKhbjs/Q9OGrJuh
9eEnjkuXap/YjcrynXFFycXeiMEUHN+biR+x+bVxvLF89leGLeEQxE4bsMTWK/ttlG5YXeu+7PHl
TcXCzY4m5omIH9I4J7BKP0sCk2OxnFdDCGMHxoy3kuqGFLl5Vwjz2qaCGv9X/zqwk44dMLphit+N
qrlBrxqLyWoa1UkphlqHISAiSF4H4q7UgszFervO8Tf59x63IdgYde8Mw0KesxNuli3fBQmMB+et
qjFvuK74A89AP1c2NEmp6ITRNs3b0by1j7wxxcya78MlmuSRBxgHuFNQx4xPLmqQr05ojlb6+zQ+
C9UmAytvprgyRPtKDO/Wmf28USl95kERLQsOl9Ao+kn1zqaLmUyvaH7/nqhk69ulPr/yUAZ9mpsP
6MuNMIvbJ65k6Qz7VagD2vd2MvX0ao+WOPvyeBYzfpVauZGZxdPDp5G0xYnCHFgR4+1dLlsqn1AK
Laf91LaynhoimjDc3Z+a/+lDnlw14gUzKWid6/L2X9odbgGhDmG5kg4wJg80NavXFCPCa7NV/Lux
SWEaByEaOs66sPCLw5/BEE77vRlGxJI2vR2gXb3eIDkw0+F0itC3Raj6ohRG5Fnc8WFbkjQmqW3z
UVNAepdaLw/efMOiq+WRi+FK793exzG2/1Uw1x9Tjk1Ptt+vqk6n+utj2KVRqY2WvqPDPb9K0wIx
f0Q0UUsuu9tcaLvp9DEHCk0HhLrhkMQhfEsQkoOivYk35KpgcuQOfnzutGxhaZgUa1FB7FoqBqFX
+bKLMclgXKSbYt8KkB6PqccUpSYOiwNI/ZJ8BiF2Rm4JtSxZl7236Noh2jKcxTjQRr3lHY52QRbI
BW/Z+iebUERNiy3ahCjS9O6jIoxaBMIywk6WVv0uu64R1tW/bHFNDx449ddbdf506lbwduZ3I32c
jWIz++KtBpPhgQtTAWp2es65EiSjfZi4CTCFYD4znH6tb9P1BnGVYKreAQbr3b+/CWswfKVYAqqj
Gsn8dn0hexvQGEYFkEOfXRKv5two/3du/SpvORWOIF7CpgIE9n2HISl5tAPTRzD82EbASmD9KkJZ
Hct8IYHUC4UU1tiRcu6dJwkQgu57iCHOfVx+Oau5FHwPw9SRzar2w4c/iPz4ySUSkKyv7/pjMIkY
UTIhh2zSDnY/wPj6L7yG2xv1MX3BKXFP8rnJikafL1x3Guu65LnOs9pqDDjGwDXvR5n7cne9VDLu
SyDJGTNoCgEvo7cMms7E88T41cLH+PxqEf5M5Yb1XwK1np7H9dpJQ2Z0BdKMCf/bMgjH7v+c3pNv
qIqEZg8WeD/jmG2RqZLhbeHdQgaLz22lkrt5R7svUpg60d19VPYIm/oCEoojcQ3L17tgvZCYInQe
HmfpmMaAkqXNGwaAjfBh8HgYFHXU1jJ0Yf5bssnaTrrzneMh3M6CrzFQflaQiYhMKwvC+j6xtp+8
f/D1lFbE9zI6aHuVDuamrf55hISHtI+mYcev76nEQHcRX093BHLh3d65GzA5IvxmG6wVYGwM7ybo
qDuNqocEOqk/2HnrNkrfOG1uJ+aigvdyJVYefEb7LFWw133kNrgoOQFFYFKgFCATm5q4xsLYI8MP
1OUNTpt9USgTbjg3Jx9P/w+fEUafo8/9xEdUa2MS8MLowlQwoxmKK9dRV+o7sM/6iQOIeZtds9AV
PQPCp9NIP+z+nZUkSiDyDlZqGPoqzCvX4d08eQx06Ctn1r/Hshj80lZvm4Bsw0nnP8kX98b45YYr
kHY7Z6C+qFXB0ohCQ87jL+yzCmY/R1PqzJYY5wcVQGzsVO09Mr6M6z7k540hNRdUmY6HKAO+k/4E
nbPuOwxs5xqiOXzyjNehBznjAzoVXxkFhRJtpao8PvwRJ/4P4V8nCSmC0Ugx+dlYVuli/hXbIYGX
HB1tIcTJHhi0kpyNLbkOKnA6Zn78Cf1kq1HMBocLHpdzV5TN5U037I0btZkAG+OB0qWZjyPkJp/0
u6Axb98mg84mdh+atWxFfH2tTLJpLdPowPSSBhnGZk6nIjsueyYcMTvTCDmwVMazTNUgs8yM0rDW
EGkWhih4fVM+IS9DfPtfOu288bwG1IXnjVwv6iNvkuCJZz0G8qX5VVNKclbQxJsU4+dZa6Q/OWeW
M0/oN9aeVaXE2Nx6Bm4Hl2kunfLQJ1CrP6sjAXhlHBeoDkidDeyysWv1hVi9ZeTwWHwzZU2SJgyh
55zz8656SIG49i1LfSymUIEm8/AQLuCk80uSQXb66tcWywqkgzf7K4HonlwiSdXUqbbbiwbyZO+R
pEumpAkf/D5iVdfajIA39k9rlFsF9zEJxgR2hV2lekjraNDtEu7ok/StvEMMs9I7iUGv+MBg/66k
ipZHzqlfzUQESy5/Wgqgdox21xiuWgOBow0xiFi7SZFEgdrI4yHqn73BnziG3uANmTrYtgZV3+J7
zf9j+HAAhakBCgi1UNFJLR/u8caGgTmQw5ZRy1/Xu59MkDt+onN7Y2BR/VxHE1qaL/lH2Tw875St
L605TIx1uhwtfG2xvg9oBo6NscBvLOgXw3GTCl/EwkRYzeMDLfxgOGVXtiHWOveTrveikoJ6g2lH
ztRsR+WTBSjG7DUnwzIqAXagUCi1k6iXUQ0jd8yMonYrhepQ9M+z7X+vm+dZMCNGJyeJcwGfie1h
UwPdgknX8Edn665pxo4OzHUqw+c+g+5+HPDFvxrfKkatYv/CyIv2ZKYXd07XngsGA22wY7IV+UhW
wIqSvFsPD8JPedcsYFa8B54UAHU4kASCGCnD3iu8eHN6XCoz1cBXCVDhDwnYwk7wNAFFzodIY1o7
wtAfrsyO0T6H3joT5/LeY65suyj0NCY/JcMIiToBLpLHX2Htb3APfu/cAs+MbquEWr8YPMDbHDdP
fmn1CUaj4j4GMOBydIzw/av3b+WEC/kurXXSqhfpg8K9DeBVr6VnCJW0FJn1ToYQTFu6ZRp/UOLt
pNuSI1qAJLZfXaTV+zgDfT06df9ekoQM/CYmVUv7f50YzZGkOq+ib92+z2DyZRKWc8bBQRKK86Nz
5QPPdZHwGsqPchws5UnynGgG8aCWPO4v+b8zoagyr6Vgd7SPRXAPnEWqVLfUpzr3H+S0vNDN6Izf
mteGjUw4HAbfppb32/XeJjO6oGU8Pn7ltU7SmAYbFdshDFrvvwbBajkHPlBv3UC/m0gymJLov/+j
W4luTvmsdEH8Im+MwJsoPNiM74bQaM5muZ6S340j3g1nrOIlNAH0zl3ePTjwcb51OPwR/pjOcwsC
twakMjqo3ICyCPP7IsrHHXwDIqw1kDg8TARHErCUs68DLxBPY/nIYO4RnrczSywUJGdnkFJtm+CC
JcsiFLPnPD29O9JtLLbonS8S7qrJEC9btOs7XV9/wI/vgTYW0ZiyjvJ2scyVy8hJzXUxmDt7EyzD
iIOsl8ufeFs7ITva/kBcPfdYruPYcpIvZR7EfArg0hJKoXV4JJZMhweRhyMOxPak908fByTWHsn5
hDgIKRaAaQLr+AwkISUZrXwDHXU3gWcUtkHw7uOfctRA0bLEMEdcmfuj3Tgc66v8YBG/aaoQHA84
zUrerZftsIBFGi4b21h343mHClPZIZGV1gMQYpvZG0qHjougEXGfyvEwDCF483JdJbz7/j3UDHR0
81KX1cb/Q6Zfbgkj6V7lBlKWTulst5sJmpfJLCkbcaS6FBlTJBYKW0zSuMbXzIwz/yRzzrV2RtQN
lEtvW9BOg+yjpj7CobppyR6YXZ0Cz6qocQLOzsALJkgnXn2J2nyl/7ef1Q38KS5qPZEI69wN50l3
jDwn38gZzY8s7KNqGz0YmeCg/fHIuA8Hfzslr3gz/0WJc2hpfP8FoahW8hNdhImRn/KfvVRfaR+y
YLZuIrvFa0bfaRxPUmy/fmzQG9qmqsAERz7rfuB7Gd8DprvnyJSgXyjNmnwar9rETrpZQEufTWAo
MwtB1/5we0gptK9oHbMXlulh6sfFUbf1tgU4p14dOaYTp9NRiII7RX7m/bDCnrJZI+8EPNHbTeAA
u8qWcpsSnqVfkWSdn6YJHML5Ad9UzgIe3IdquJTNDS+9/U7DoZ8fzhz9lKCy3GbhwrUmfjCb/Dcv
/8IKT0KI2X9hwDxCx87TJWtND1JOxEKCKoyzjakUB2np1bEomZotkRDhzbnrEpQhtmqg5sC2wOMU
4yEnFjKPx/0opts6m0qpw2Mj4JrNGZLUibE1Ceo4V/RrxxERZr3KaIlFkRSG8rbDNk2kMmKezXVF
//ZfwF1jT2p4kZXnGiDJBr2Ove+DWhKUz2oY5TtQeYevlUOG4MKWSW3u2t2vcvOZQPbTaV6mxmrp
m57klmdwdaUUxoBzXUI9sfrgoFjAFgXWpsU85mclubhpAMdVuZ5NiytRgcM3iIms3nagZoYRoqCc
i/Kt33yaGjY6O2ylKI5HJ0GU/ymHKLX6aloh1wJD0UCaxYo92OWuAf87CeDIMltzkebmtkgXwzCu
osp6g4pz17MwbK/TOnl8z3xlABUTSfoVnfiZdReBeMrB241sAhTlMaasVvIWwEBvyMLNIyTxM5j0
T5fmmNnc6Pps+nIbhhjRs4E6O5jxIHZM36dyDjCDU4AeQcs+OOXg6ezbJj0r701DFn/Go1ZQUeAt
HuRSaZwumhvLgqYXqfgTvalG1Od2axoPu9hi2D4YZoS7jM5td4f650OZBTS4UNYzN8X33D4QeFgv
0NzFvo5qj8fm8whRnMloHVk2ORWDGnvTZbE9g4GNYC/Tq1muJWtRBEZt82wDtfnX0OGEr15CO8T2
edGYj/yft3/lXy+FVE7iiyPIgHH1tqi7lRRT7tO5LmKGz6iWulMnkf1d7MA8tVszUxPdvAeGpCiM
F6adW+LFxWGIvjx5ZQsuDG0quwpfgDNF8RCqwB37bB7roIfKugcTZ2aw5lhSoaXaVskclinFPT4u
jrjuRie/5h5zbS4SWRavr7vOFZmo8OzGzL4HOOfTCuk4sRDVX9gncrWfeOrqu8TCwEuMUimy/xI3
cVaWQWDBxh84xhnhAA75KPbNkeoysh0GkN2mC4NDpv+zA50zs0QL0DbEPkLZ050XX9VnKSa33ajX
wmv6OYg9ScLm+ugr3NAUVl6QpOQH4d039YmMTpIyaWnORz8lUkCLWoNs8b47sTeDGBrD/Wv/BEdR
nJdCVseGYrtQb/LclOMQcZkdV+tqQACwBN83lMcyzbN9xAtFS02pWQCmLueBPFdK3Jlp4mRBx4xp
MV9PinahZY4msR+9kwb9W6ZOaUSzOxvDHWd0O23zgj5uiUheQUOaN5v7KT+ZN/0+CU0xePvqb4vm
ymE6G11xzEXOqwfLWMaLU0ajYyb7bPCB/4ADwvolQMTeVK1jLXwK7VOvfcT6wyjTDVRMWCl8WwK8
tdmY3HD4KOgu2qdNYh2lc6WA94zTeAMOWrcwb5lNN2geo2VUhZryrigSvIkDYyw1gKsyfKdfDWWw
nVZ+IwaF/aoxW58U8ILwiOWHWCmajwQ4OuheG8wQesV1SjXlmttWIW8HdqyCSqaUZSiX+6HExBqt
1FYOZHyyWHgzvyStLjxHdhlPXYW9TFk9I7wF3/fevpnhGLTtpQvQShJjhoQXBwwBeYs1mq+B4CQW
pCDvgBWUo4TCJ7NjItXZ5avTW7Zi5223KnN+uam4vDzENnllqUEAam3W0e9G7dAEJOnKTIDFWxeY
jO2JrpMWHUkka6U9Y2AyNYtPlprmeSRDPv1SMj2xFaEb4mCJ3Tus7YtaKrEk5lGzWZRXETCm+V25
z9AXXMLKZjEKaFgoEZqkjawal0lSZLs21ZE26tr7ANICk+jO+z1lMw8bOfHOrcr1TmwP8NN8BZKK
M37PEk37VuT1IojRVRioITVWxCrv8ch9XeSHtlubjFcqIqjgbmUl9XnVcjrZxCzCBLXV7iV9WgvR
bqIcuY50UzVcjYdkdPM2d7O9H19sj6Mt+2or+9nzdVT7/6i0g/Gxx7xnQZF1yBspAs3kIWmVDSrj
6kt+ePzP2hjRvGKP9Q5AaMqQYFTZoYgJ6JP+NIY/46BBQaF6mhAHh+Oj5ysz7qdvnoj3D3kjwSdv
GE1fjPJjVPP2LnAYj/bIyBwHY1Wss/NfF9d/DAsZ0OBgQt/aNKzfQHaFQ5erhhQ+fZlU1LoWroLw
LVVSuvHqlYCGsTdbgNAjUVgUNuGqBTOYrLVlz4D8IvPndz0HeIJhy5soicNbY9LwQKfrgqMMsqGF
F9ftcEhdKVvJpdvqAKewhdQ3w+d6Tdrr9qLBdTY+VZ8RCvGukSMhzNMcLp4y9MPrpAcNa+pMu/4S
FGjyLrA/b4LTZfg71hGU6Tnk+FEhjmSpW+B3ghvYEayCV9B60GTQVniuhWy3INwiTumFQFkDRRFc
15/Qt7sepVn4dylpW4DMkzahMhSXLP0lcUc+tn0+NeR6wSwipV5PjHohrzQJMKcjwq9g2lzjmsMA
OVcUbInntV8xQmGUcgJ12Umjkr48ezp827agpTFq8/8PQAv3qNxh2AuSrkUJ4Rwyy8MgNGd/o64J
Vv+MMRFoauxtJokFpeZ83sUoT0O1D1EATA4aOYwhxBZ6juFfMoEz310qObSg148EKwhPzZsXtBUw
ijH8JjLO8BOhQ+lmkPbLU18fbfZMqr1/XFqCtdYCYnCdybMXpvmWeb1tHtxrowDbD04cjGE4ZDLG
5jXFJ+Qm/yi8tuvxmSxk0rjtmQaGCmfcvShkKKPjDB8/8XXS7qSU0bRNZceo7FLw0NknfRlvjz+6
jNZnRVDf/yscKkl3y1XnhGOO2hNgOwG6Pwyn2jR16NWlc/1xGlPulbP2w0fS6hAjNQBwCIGcq5s6
tBnhOirXlWk/ozmXGvK38hC8FDmT8jfL0N1J7hStZgAO663yDAneFiQSYoODmPoZNvQiJ6mt51mZ
1cp3qsvCD6oVb3TV+tg0lcSo1wzV9tlLg9yHWYJDltZx+ZvnvgLyV+Uh1a/mnR5CJE3B5jIVtXty
FJJdQdsgSAxwEm54WON/NuYov22cqRLTpN8Zfx3bCQ2e1jaKRTiFUux33Gy9kxUqXVoPYIfE+w0K
2clBv3JSfN+OM31ri/LdpuTizAWqN1TM01DrcSHHQDSbZ6Fj83aj+HLPNGh/496u0tkS2ADxrUii
dRZkEBCiLaDufz1mAqdO2iG+dXDa1hU9+3HyQ3+ZiUdNzzEAoOQ+gZTu7V8f9x2vrDVuPyoxDPYB
rwKadwGrWEb6+ebmpxiG9qIu+AJIVAZVrssF5SbAxixnf52YFxssm0akaQEi9V1z3gqDzgAxa7py
a45xfyPmMs/BkfEcS3Vwm7vZSeslkyVDQUYDeEl8EnQH4Ef81izH8Af5p9Kt54Y5Za7fAH+f+07x
4+uo3JDCMEnlHLdNb8yJJN3i9VLKZttWzj6ehBklI/Ll7Ob/7+5Y8eiTT7gCDFrc2LkUcWh1ruBZ
b+9j9FsJHknoocKkq/4kKhmrQ2/wWNapQ6e/JX6JSbHM4t72nH7vEdFxUfyz/AG7mwPDpMGabIVY
OPYE16Q9wV+GQjQrgSy55/cyQLnghCJYxhHHxSTnAR/vgkHVthtYi6UjdWLYAac1V6u7/7cT+wmi
N5sNFg9zjZkzBIL5P2ujZez7D23owy5mHssWUwEdPO80SlPJbH+SbeGRxtgxcb+0Vpj1dBEP9935
5XyWZ6BgfgrYwKeCJnoR6eiZOmPtrQtTakJiMsa6FYkxZMTLvCScB9YQ+SeTMXyjDaGzUQTqt6wP
RE//5AyJeF4fZNlIXMZtduCo69krmYOmdqyJbXsXHBXO/K8J7ngFnNLrz/kQZ84kDu8KpzIvh+cB
fdYpDUPVybdwZmapvQwKzP73mJdcmGKjrq/TqUiEcmg4QZcsodgIgcKtARNgUCGaDr6jUklzPMIH
ZyZ7y9owzcHq719WvWm6dZCme5qOmRfQKC8eh3jW0th8p/brsXFB2Csh7tx5QmG+kYOzHgsCxgNi
W9jgOn/ETAjj+AqVgJMYSQaArwUo9UXBEjZlX9ZttpoLxFy642oDb6mHe5FowHf+xhrTPsFGnsch
3ZYTFmNF+NyxWwSsmV5iu//rvOKdZ30L/boqGnUyk+FekylJG3aQqe59N4G1Q87CcXF/Y+bYuKgI
hsXVnefoCrqRhVuOlseb/rkgcXgVYPt/rdCTVeXrqOtFHQ0q8Jv8aHvdETrvLeppYNZuavllRZ1I
tpvhwVa/WjLKjtRdAI6oO1OtRfbg2qo2/Qk8eGYAEpjar/91PKZpAsDKJc0V2yrje/HajwTAe1rX
mPfZbSP/4C8XzwPLYyoMZGV7ATCcRXy0ul0YMenjX9XWjkbI6bqTuiKdiGLbKlEHhv0UcQXoSwT1
YkNa2wp5+fkLss6W3z96LYn8cI7L7vJ4fpiAtJ6oFRQJwi8gvG532DjrUZUVkz3+E9/8knSPUu1f
+Y4N4sAIdN61KXlZt1NdgBoHfJCNadyLkkQan45hGSn1xDrXi2CHE2WlXU0vBRsySB/NxSlNmHki
9cO9PduW5EdPKVimUgksy4ntK57LpNocgBi/diPn21KN2XPn18B7D4nzPpOsUulDay1KRcGKOljZ
b/h0LzMf/oCmptqADJ16rKXesFxqEBK3Up3op67fNkczdOTSfwYjqthPu5Q8JyPAQvrCZ9SnZH0p
Ev2QsmZZ1hdS7wWzzaauUQf6ZWC9ljo5rrPfvvefgBnQ+HQiypV29QdtuFuc75ZHZXrZHIKhnTpR
JyGH70ujTZ8i11iIjCNIvMVGJjdXdpAkENIV6KhMGB6E8BrCtB0BtR8nfhWGudm1sioESKLRFXOo
JbWABwHvHIpXtEESwKFFmZT2jhYR4Y8zsNSePOi4Px0VbtnKTeUfkJmWjZEb9Tl75RJ4KNEYsquU
mLgBwK/y0wRkuSRybp5n1/BMn4NSkRCNZCs1QgnBItXDt/knwOa+l9kVZr0uGrB7UPu8/L1FA5nC
59NePD8DAzikY2Kmc8Md1sSTGC41hOkpGhZiZR+Q42wZ8GO30shkd6OONHVSnocq0uF/0sl2lm8L
QVf7jXtcQcfswBHV90BB2QwBCEn8CiuzChueDX7ErtMXl6zl0D4vK6mO8fBLyajYxG+oEgLie8Mu
bJt+9qPfQdhQOLTAKSCFsoXCNymM7hw2+bPv/kOyLzvwYfkPtKYT+Jsfxv4KZcHCtALpmohQq5W8
TX1zmoHqh86kjkhtUtrQtTHCVW4O0MgGoifJgtHSdtiZWTB5wKyRcoc+bTjiSmq/2DyOAu2NSMmf
7a4x8S13HXUx4vMC28Y9JKnC/ySVMYOhXNWTmgOQK8d0M7XQG0OREbFVNrcwmJ50luYFkqLTrdto
FRdeeh59YH51onv01jKGbdHV7n0KVxQ/dLXLBtqxN3YbHTcrleuJpLhWj9K9hoXTGQ45CvLJl25P
d4GlFH/cmNVMW5ambS72cj3Y63x5EUKCMtyMqQVRXu5s0dmZrnjhp6cHDoEAhRtDTJOsaY9YWnvA
mL3rkl7lOcRqLdz0hhybQejf0CRMu+fA+U++8GTutrnxy1sKranQNCLvhVPGBOUQIoDB1Fve6KxC
M27CEsmSumhnoUqpSbRk/d4bq7/IYEudsFt82rsjoRaWcRLXlnHeWBVvaPofYv4W2PbBCK9ko85f
KJtdr40czrlaaguX1j+DeXIEftgd0MEPCk4lAJ6rzuu9+zyTRZE9DODjhLfJL8nW9KviWCCYbHvX
e0aQOuRVbkAtEoeBOBWvEDwA5VKKp4h4hyG3hn8QAQSiq5pm4z6ejGuUDqJtpK88A0f7eWF5MQ+o
JWeyuqAEh2YYXdxpc/Wn8CQuTovOF2kY9dlhqPAjmAwluEestjBT9amqNmjWgFnXQXxnXzz3JRuf
2ONMymXFg+eYLRESMzQzX9gciQRvPQN+BTnlSCh7ST6Pc78GR4Lz3ms43rLfBYyvTlWrwfaINhB3
txLYfr9zHZTxfrwaGDC+lRub5PDvHXo5jQ9XlqDyK+ZZJXyIHZbaDvuzcje8XtCBDwWn3Fb/chM6
uRbMUmEl5QN1ceJMozFE4sHHk2pk2avjIkx74UaU8j1ZDcsC7LiUlSQTlafu0B3eNxAiRwMx9MM3
qXgSyY+SxPVs65OBr5o/rrEo59r+Na4B55ZUUf2svYwj5fBZEAC2YkSCaOaROxTX1i+8oOQvRAQr
wTVeMQ8qheVe7RWmljjZCLjw2vXl85FIXv+TCqMajD/KoF3mIniOekeUlNoQJASkWbPTaJEvl1lg
Hjz0PeCekfzBT0Wv4bZhObD+lGpfe64MpPdkUXcpbkXVddrndAOaK7S5Zb+b/o7MC/2XVGL7yDGO
N4zYv6FibWT+D0tuOR0oz2aA2ducUc7hFR3Ap9iWC8phTOanU95yRZA+UDey/wKxA7eqIICuhC47
j/BBcXhKAk8fIpRF3fKkdsiBKxSOLmS6ApahAnxjgZ/XGAC/aE9Dj5D/+frWSYV7G7mJgInHeyhF
nWtTtXr1DxLAR2tlPTT4aJJfXMW1cfprPi7OqbWtSOu7lx8NrjTufFR8IcWji+jX2vacdjm+C+Ui
xy6Fh/vQ/vFXkpenGHXdhjWqlnArqDHRdmzDYylBWmNZjCWzBnby2mi5RKWQSFYFKVOvUVTfTp9y
TlQjyKxq1tHYR1irFfprMY8PTLzDq8uWna9M/VwvuFnKq699a4RRPRbCX2daoE2CjK/f7/P9N/6p
L3tgynJ4b0pet51GHp0WP4zR/ha6hk4OxxxUJ557e/DzFFJdY4LS+W0P9eajb3AoVoGGW3208jZP
dcL543DyaIIeQwwnazAFVhbM/9Z5cixE6G9S1Y7XkNZmErX5tGJvLAgRcTrkCUW5frgEdG/pQLh0
vhiWWjnlr1Acx5iBKQJmhKXifWLIvNbzOZfZOw3H3cd+5UrfBEtkTHWnyf/GcIf2vQeD+z+AQISp
vtlwT//Eu0GEGBjQKgtpHiPfLGZm9cTyuYxDfkIn4p+NSXeU83vp7sQr3ZsPsBuFDDeYtwslCKog
N1oau1FlMYHkg7ASpBFgHqIw8VaqQDyzKZRwwakBs9bo+R6Bxtzs0GQM3eoVk3iyWQbkdXfM8kts
lbHDySgBvg2+Q325ww6yeAyUVO49dLQ0UW5Fj/pXYTSni8hMCf+DlXOUl4o23QM1cvCnDA63Xu36
LdqurDUT6cx6tNqf0tE46oymiTHd0FB67mahMTBeq4ginO0P5LNwQ7PluTjxZEYZgbVPTLafYTSN
EtgdZmz5pmow1xbPsTP2KW7IOKsfdXLLg3Uyy/FMSuasNaFT91IqTCv/+TuQ2N/GsuyUuLWGNVUs
HP9fyFVs/cEbvTjOl2pC/ryg1AWJxngwfKJdgNPOuWEKRC2l/eolLIWIGo/l6ctGfOyK836ihsGe
RTO22KgKjRl454B6crnpK2k6WPQJz1D8cAxkM9LmExlSWNT7EhU8Imqj1CwTjHFOVGSylYBXQHl3
OGNsowpaiJZp14AWTQhuB55U3iCHfV+gWSHUILo4x7eUdPyyWE9O9T0HZqys1yfyy0kPCXS4vz/l
NlVDcXkBQr1yQaSvaT7Kal0ELA/59DY+8gthkEHgyYxdY76UZxQTjr90tYq4uX7r0B1zzoeM1n7a
FQp1rvK1o81+7Z1iHVKwhkoE1P2Z0vZ7DN7m/IswM2Yz4Ny9gJjgHIHMp8Xd+NbuUmSATZctnAGs
tT6qK7NeFeycUzM/Dv3vlzQYt1ms5ULcmr0p04xkzrlOZtDIyffoCeGPFof1qpnHjVR5hNyC/LXQ
jTPhlDZjPYDY6/DbX8YPKsUAiTYftG3jVFBNIPCBBwJuT8RvYhHnsEG2JLUFG7gpgRqhiTz+psLG
VZKsjeJN6gIzWgyHUBR7ibEnUGvshGAmblYCpzliy030s/2HBp3u+lsB7uCAV4PTnzXej/S50WUF
NE/u/9pnNrC+UwUPxcR3lzUVQU/lgo/VydI4eHvmEJn3ElV6dbIgBo1B+5AiSgX2qyKPIlwhmhLH
+b6COc9g2GxdJESSffCo8+ayzVNedXpG8krMUxk4OYbUpiv40wGjNjTFsY9+YQd4c/ZOfTVId2lL
xqMhXMU9fjena8L25Ew3X0BPFd+PyaU0mi4zOOUpxu10ACtwUi60bOOiWDoi4qbUFMO2JzeHjlgU
EDHdwN8RBo/DSSVWUP937dGNf+9BD3XbcKacldspZzXmCExeal7v1i9Bs/7Sar8HsRALZl3p1Ekb
mnfeLRRBG/8IzzpfpV1Y2W2/wHb7Il7Z/yDCmLgI3RdSVvatbmgGD8xziOJCQA1cDjA1UjpjYw/J
mYM1ALC5xyUgUrnbUTRH0NYfldGeGXfLylvejy2ByyBrbsCShXUGO0pkZd+NfZHr2YfwQVVVBZe3
/oBTQZwi9gNo+5Me2Gu5nBd58u1OhEeaq9yCLTk72CjSZQ0iVG5IRhr/q7J+SaSfHTdHuS4AFEdC
NmUqFKHcFEauPDQlZSyhDCPY6nzkNuUNoJiOn+dbG2JxuWxKs/mvBs4efBr/wVgQCDomFwnfpIYm
Y0mcbYE2auY+5+DroF0DLEN7EpM+6NT1EZ8qE76a0xavl6SJPc3QPL3asj8kcN/5I16JQWV7Bgzu
K80IaJbPdK6KFZu4d84H2mgLcVlEnUQQmRwE4cXR7CMZsdh3LmPyR+NxKNf+n+NXdLUJHPv4vWmp
7EZKXvvKrGzDOUoqGqEBed0MWKrPdtwhM57kdr11tWwgWZaeFBnkygoclrr+lZ1TH9DIQHthA1Kb
dKFk4CHCTTKBLefOZV+S8yIEhesKpCmlVG4h/AXSOjT+bgbeIQSR1YqdS4fUpcTjqlV6+ERP0ogx
eiV4Of0TXNOe1RtuyPRvdiZcaOctjUN5QHGTQELHrytF6EvKtia6wmPBi0cErxWA6OBIMO6npfl5
Rx/ms8/K5G8OV7wC60zrZwYDn7onjO2HV0X4Ac1tk9quTsghHWqYqA+xA7noi1OX0+DEU5pfAo0J
6DOaUzuYwylujs2OzYoPp1Q8OIUGjxl5S/eDmEuYLICBRz+z74c2CXoMp+cBZXYxWF9rVZ1J62Wo
4pDdFQI37804sAk7waVPYMyOsVqkrQ2vpbzdlECShv/tA7DFPC9we4ETTjhnX7arzrPoyl6JNKQt
9QYZEBNnrzCS+9UlLaXfsPY6xCkZkWLqzBvtGzxiB+mOIFF6+ZV3XgV7W0ibL4GcGgOLXyLQBnaI
eLWT+suDqriWZNCYGTegIp3xuGZ2vmG0imUe0w4o9aCY6ol4gNmVQbTyfZRZOXQDcmbFoeA8FTOY
+2Ua6I2o5W7di7O84V7i0xxRS7q9SzaM0LcUbJb7+rbjSCrFaI96+ClfdLkuZ/8e8U6YKrcv7iGG
XAM5KZ+CwxeAywxQH4g18qc/LpUDitUfi/NSpT40DmB1/+Fi2opE3MZn1rC/ThyH51g70d6f6qIY
ngHBdQg9Az238RrPH1JEW55Pk+5OmFoOkq7NWFSfeXZ5zgJeBwDx9c1nxo8swufQ9rrLm6eUzKng
OfImKI4RUUiiCGqPvXZAvqh6pgkE5ayKHFsHdbp9oHe/8ZwM4M5bvM7afua2IYH/vdSIA5h7xCMR
F1M2TI9pMTIHGKZuDpTU9LXYn0EE76TQlKN0w+Gc+V077tFJZhllhQuenNyBjW1U+QQJcVnx0WeB
io6DpFevejMqKGO0Zv9qi0FXkJAgwvXYeTi/4nx/b4BL35gKN7/Nxr7SZT7IiP9uhwYQEQdPdkPi
P5IeRaJjJjw9zt5Uz+I9ptAvlK1AFXjJBV76XvUL6N3jgYUi2Mm6EooEnjXNQ1QTV/jDUEXKnknA
hlFXdg8iI0H3mfEDbpGA+x4FbRKeh4OaZKz0yfKTC91d0rTw+HtaiktTC/wJF2P0DpAMSN57kEx8
iJQELtTfSVBiSRzTmblPUCz08qWMGjCAhbmU6GUtWdzWUu2f9i18dO6DDa69ksDZV3PczQNTzrie
eOsr7qTE2h5AW6d1h5AbzlAGUb4Wb/8Dt6eJey6zfn9wSlkuxu+ZO7wBRa6+A11JAu2c94tvnCpZ
wbJIXVQXV+1c8bQQKVRm2ZAPwc+vBMXrEhkwDwOmSTL/NIyTeEW1UO8UKXkYWgZABqzoQWLRiZhT
RanqpOCWUupLQ6OAgWNIwp1hrCw2cdBx2kow1FqZnH6l5nZ8QFIWa1exrmEKJY8xJ5dF+JuE2mT4
M7ZbVNVoOAjfehEu92QlzTg5l4HeWyVfXlhmBMetK9enzLxWWx+rHgH9b9ott9Yjhq46x/x+Ju6S
NSIz78iKJ2MDC7zRPtI2BqlhaLnk+yxP2lkJYjPfpcdi5/7ZxudJxBrGNhOp3JYO6nH//D/s7ek2
r/plsRbbR3QlJCMNxa7vx0AdclrUP12XT39k8uTwXT0eYmb+AOVYW4X5tTmwsTgLrRaDGMUbuWRm
uHPupB0+za2it2mqAYhi+Q2owdt95hmKO7xY6MHtl+x+YRgVfub2bV8waFXa/l0Cvs2qjH+/XJfX
o1aRBkcfZkXPYzSFC3wVRhgTw+Vms5mwUe16x5Kt/LtFxnlJuDgjtOEllKYoWmwMwdd5u4j5U6sX
hPyocwAzrzCMxjNgaXZfvBbs1IDTf7njgCFTESt6JVNUG7uty8AAd9ebybqwVJCuXkUYYsqfigjT
1bTrlrsU0A5hgn8v+5wkHwNkwM3TgJz58y20aMTHeDlewfa+YjDppTSyA/OSW68TxpX1AuoDjDni
ez7Rrva4wcZxya9+ciwkG8u3V8Q3AYkMVRS7nBm0npvv4N+gErfuyI6/qwhvEZIj0CBBlGwskHOB
B2YMPK+BUbQ1mnTcVY5GnMhdZHeyPIeI6ZvbcAHQZVTS3KnaguGvgpkKSrPJ/93ERU+JqabHHSzT
Z0OZjoN5ifzOD3kxiEjqAj29cq8L1lnfr/+NfJtHlQ6z092jo7u+gVFYk15EVRPBLRW9w8ybrxZ5
yiXlZnOKMq24MBpB1t2HO5vvJ7mFKrpLsEJtR1FtizQd8xpq0ydn0k+z+1IuP5j1XdvIyvcdqnja
sasgyyIAClh929ia3f43pIu5hjsA0q4weynk53/Qa/GIBBKJKvLFrnM2yxD8sVJM4Xyz5yYG1PJ+
Zyeyq3DCPLPV7eRNvS7v3hU9Fya2VVlnyI/yEkySBO9lSNluQZgtSFtXKv5FQ3z6ycr2f8JPmyOW
e4xcrHu2OO0Q8kb7Go/ylbKqOZthGH+KoTiIEmhXaFbeoXOzm19tQubea7SQpM6WplJ7If7owe1T
Je97AKRJlOU1Q9VfnSIQDewJVedml0GPdiYAfGs9504doPzOsHGYuvDbuJENudjk1NNVShqC4HwA
/FS+PhrW2QX2xV+y84i9c2tsGxG+X+obWJioe/yIGY75ATxM9bD6oESTMHS9POZatz2jNo9rGxTv
Ddf67ba0uJ7/xaZ3+0R5vyJPKLVpjdg7ws1I+SSueyacLe3HZ/1T6eDLNpp/0VcEP5kHJKfy3DQA
rGITsHORcxi5t15rJW7R+0JVGLL/j7bdh77lj55993X0d2FJYPy53LlY5Cs5G79IQIHXUMQhZW8n
WENaPgtCksrLV/ZM3hk8R8QXB7DeUO76Ct1rPouo3FtW7rjGkFwFrCRhhpN+fZ2o84pmwJaJ7FzR
7geT0KcmQjMa1uNq8tPalW+nsRRT5mUVhGTKXnHqIo++0SIFMMqMOKAtIjbU1UJz7XET0viEMdTX
1VF8rB7mfApzhescr0pR5oyQBB44OFFKMmgEuuMnXwGuT3HZUHNzz9cJfjUfKcpz7H+GnMMW+NEG
8CP8C3/IEFQU1TbiRc5qs1/CKryuwr6HkDE0lTYRcj/1R6q7Galuhh/XXPqFR6rh0fA7vHqVKwj1
4OUcJEA/LyJJQyzJXTc04pUl9k6l7W124Sae6ZNnEqJxVwKg2p+nzw6QEgKYCXuwW/FpKpWo6B9c
LftO/5HVv5Xei5uX3li/LjhVjqFEKPPRS2TXsOwjlL7mCOsHvoCAuyrRKPEEci/Q4D1iO2P5hvbw
aebAy6rDM4QfoVkETO75fPA4WSwUAB1cbtm2rDBhqMSVBvAtCUSXjxyJVYhA4Jh5FdKR9pulCi5Z
8gVu4hgpuS30ihkyc/Ypig1pTcgdebmhg0bFb28dCHKu65LqjN1mC5YO6MYDkMMEoQQwlAGoxd4z
LA2PfL5g2YSSeXO8fIx8yOfBH/U0XSFRPjPXxJetq+LGCmGKk0StcFpCYupiJbVQzuXjwVkbmaTB
yzkHYJ38yb8lmq8Q/847Iy8LSQTDSetv7JF9HxOHOaKiqxdjMOygfJdVG7njLW+F/Ane9Fz3dgk/
rnmHIi1KZ+iDZmy2LqOAWpD5Hy1WnsltHYk9NI+7HNYVXIStdlwpMMJ7G7drEOVAgpkVrdJ2ZpSX
u52W8YMI9hdmFeifSN0FyYcSHZ/EqHG0tQKtdPDABdGHFIF3BrDkvqncutspehwQbNNaUdcUVzSP
xIsgygAIbulSqTYy4kbG5HToEAwLLZAp66Ndses5Vgty8bzrbGZp4NgfEh68Czfq1fpQZRGM7g6U
Sp2UA0dY8A8kRfAmeywtV5tZh/LFfLDe8A9FBxtCeW14W6hus8YlVdmBU+o0YGuaEZLGp4q/KlIZ
bBdhVZPjk9yTlQXtdUUyLrrK/we9oG/c/TjkealAvZms2frr6AYaSmtXI+ua6zPEMIRPt0j6QAy+
siAFZXT94zlBCZlAFMRiMQlz5yaNZt8PtXN3SPXEn66ELhj+3K5huN7KQWnfkXltdg7xEKNsxL3y
PgL6bVSSRm/EAYy8EtbWDJ8QbI13H1zt53nS9ahFZIamt6DK/0UnCZyHOweZXjD+Gkt/8zNFrGAv
SgoZgGNkAqksrgq1FsNbcBeBDpnS7DH4pJqDh21SK9Zq4GNTG8zr7AfVPAzTFrYRzY90XZm3/dyJ
WQjP3S5Fq1I+HwpZDVhfwJpn1MaoYQs3Oihwj1XtptR02XS8zdv6Rcf7ORKd0Ts+bDnxQ8s6PAX7
3yoO/0F8PeMpeVqwbGhd1Uj20VOuNPVpT42H9oLiokkq+fdGIegavJSbt3LK0mKh2ptws5zpdYL5
hPxayztGHnaC8ylXgTrRRG0O6hcUQ06vvu59FZpE72ohVj7qkRqkqJzm7/KMcJEiDJnQWUXmEq+6
mXL6G85UyExkNtk8x7bS+q08bCbUCcXAbh1CBAehkQsmP8jyVBDGji3sivkqn65C3HvSVClo6qNC
BuNZKiTF6DYoyg1oXAtxqkRsm+AnGcHf8abFWzAb7+io+uEcsqz1w/Stvgo7B+ZIpCttTqdtgYAd
H3yIHGAHDsGyiJ151IdEvAJwScu5VcwTKtCDBCRUrId+lsU2Cn/ggehCvFstkOb7dZEgQkd/xD9T
dCq4rU6y4emJ1uu1uPZBYhgDGVBSmULnCMsha07JZvrd113VaHbZWv45fskJn8ytWzfXvLepplr/
nixb3ZaydoDSHhAcX3cM+bofk+jQwEmf6tTLzFZXftdBg76Ul8Wznn3G6BwYyOJJDdCbG0jTuGEh
ZIeRZtB2Bn43vFgdfXk1TvQyHyU+HSgavttQ66ERvvOQhoVR0+Yxx2NNVBNcXbi6VuZg2I5rWWas
7oFq9ibnyZ2HWOS56iWxqRGqc8FVRNQmpg12NRaHmAYao2nV62ySMM8wcGZp5/N0Dt0E+iMJH4gi
aarMBe+wqjRhoXgQL6VkKE/8dpQAJJqy8G1/bOpbKKXZ6WuxGAi87GerVAZ0VuVnYAT0zNBm4Tfq
wEGMfTlw3hVWZ3IpogCK/pmbAshltO+GE3TVHUWxOrlDVEPXVLjHtVsyNUwO4gv+kTBElNMmuVbi
yS16bXT0fIOAeBGhI1SFn0R5LMHrdctMZZI7AigVW7cpABocBLN0iI+xNZfLJTSfDrYaAstr8Y1C
iFZ0jcU53mbYCCZwAuLHNkU2FhoOubG7BhhyllvCymMFKzmg2nEutwTw6S0VBO4AWqEqAqTjKY2C
z82xFY5xNCshcOy6Z+rLkpknmwWeh6arUsIlxd/UK9N9NGIyESvN0mZMWOOjQ8SQpBzIvmSzR34r
6r+vdMqG6tiGIEnKnGzrYgy+bs9D6M6SKd4i1WUbTulB0wFwH9ZpBrVy6Fe1/UlI/isBt5B+uyUK
63Upr4wwFgynPQq2wziSWOqKfGV5PevrIX7pPio0bbH8ocL6fKV/jpMI2LA2nrBaUU3OeDrPDckL
gHvTe2VOa2shAkR4o2aFkbTSBphBNtxRoWP8Nw8A8Z9mge8Zf0hWqHzBYkA0vs8BIlYV77s11WNw
SIxfs1XDcUjylpy0COCl0WWmhcZo5+a79gzqbP/PIenG6vecRul2L8rCiezkSAgUUpvffs9A8qY9
vAxwznwfH8gYJpea2CJHrdvJMZeYtkM8iJz4/n8+utt+rrucoZ5suW6u0sH9qQkJCYCMjBEIWoMU
syHijSwC7HTmVXOChNOM06mBc79STzPPFzf5rUaHPI2nLP0Vuy50oIHBfKzR4ysm+bXUO2y4pc2L
RhA/+2P6yWTrcB71vgk1wTB2M6akhwPKPZ/NeoUCjnYZW/iGvVcNie5YjyZoX3nU1fypgPHeRVte
ZTeikdnM2M0W0AxCQ26Fsl5iBR0AUXsHCZlBNnuYP1LCnfumCgRcQHykSWesB1kbT8HzuFLA6IjA
alMKAZdHbGpUfd4ehlKA89B4t85ecjRknSjeHDfpFVTTDPEJ+ZCWRTVx6IVsHcMS3P0UjyQOFRDJ
9S8v98UyZcv0xxagFNtCfX7CNDa5eqGAz3Cx/hWr0++2YQYIz8uBdJlcbwN6g6kLigeuuTW67VFO
aj0ZBQH/qvKyVIUNcV86N8vOc1Nk/Mmj/CvO91YmDWZL9ovEKGVxPrhl4jaJnSqXs5luUKA5F+R4
OqycvWib8dY8bvJqeAJKHiAQJllV2EVtufmobvlhQiBYVukVSIIGofYgw2Lm2s1Nz5JhrTSrc7zC
oD2BtQ8kGZsnDvo36kbmDStrE7E3/RdNxXg3yu1TFJZ3H4iunHIlT1eApcoENVcKXE3NMp/srJ3N
NLzbJmSOhhqQprCwjZgpXb9l+BM2jhwLi4ujspNSHUZgIQvtCQa0c55us+FL/sD16TVsWsnQSngF
8nwVPbJtznMzRgSfRTcy+Z5WlhhWJXCq6PNad39h8UaEGPToADNxfTiN6NDFUz2gMOxP39vcZpia
2F8AXbi+XDYKO6GvxxnpVYBwxWr8pB6kTH+1HS98mYHgpRnuaHRIThMQFVcrZoPe6xOh2YeIBUsd
HGcjsnHA/VhpA5Em/9bEtspNGiyRwyI/Gs1jHtOMPJVAIektenlgkEzLNk/rzYzNNM7TrOo5lBti
3TyHi3KYMS8jdeVYgnpSXHcGCmQ/SuSoIs+jwBNnT8PDO5rpvyq6Yp9KCrl+tCg0DJUYolKm+ID7
L8CV4sCuUJlgzhJ/S+4XrP+drW2wURYw55yNQB6LQFwxsgBw24wuzH3vMkhUkOSVGEIhOVnCVrxF
xKCBCnEZx24ojMyYJ39Qbm7AuJ98C7FonSO5mNJGHTJqyfhouh5AWAnsgPf3hrucoJw7LuN72KlF
IZt8XEvRjyTCXj/6ieqmYzmuDVrqoT8re4pqJmx9ZZALoyIsYuQscEQ5LYH/Ga4nK/XMgtrQv/qT
qw1tgBMBCSbcnZFTOIMqDesHKyW1ePQ5y7NEVLSMVUNHxrl/rZErOM4ZxmKsN96/THAaLuGgI31C
b+0cM906uXh17UyZFzoDLkcgS2HEl89XrD2ttgQqXvCPqXEzFojP5oGp1QMS/Z5XWG31iRxVLoK9
njftZokg/Awf19sS5nUFTPr6XTtn4WeEyYWvZ48yWxEoIucNmrqgElHRcc4Q3e8O0eUZgMR9KGCn
zfOEiPM1BvSlO2OQEsiAf1DHg/9iM8gLEdIwXl8dZPl38IMLB0XBhR0FqbsFc44/MbC8lKduetjU
E4nJrPteeRtw+TyF8NWi/FR4C/DtmoQVM5T1y4UduuNvtaVqEUe2+LRj4TNKE5snhBrSAhd3VRno
+cJ6z4zlhRx85E4s9/qnUV97IR83BV23RCktFn+ro0nTgykV8e2lcTUAByUX3VZ217mXXHFsBQNw
+W2DNbN2+VlOl4niPCAQshl0lQ4qv32xQhuizaDdaoSetUumxp5Xjbc1V9VlTCRT3p4KF7szSsCo
8r5J6n86u+sPR70rRu1xFnNEZ3p/YdJzR//UHo2rxHlJbR/u3hPx0emkpLkO6vrMeX4i+SROVxMq
1oM+2mo3rm4y5nMwAvOiaZmB7XA/h3oC15TKJdbrAj45x0slyyXBq1YF+auKKAoUnm3ttMw3yaxB
kzl2VJVqBS6Ma0xebeSB07qe3FNVUJyXUVnb8V2GkYOJdGuHpyUzDAK5TD8xNhN7HQBknk78ZsAN
QMEzXoLt/fFge1b1maw2wiObS49TRePGKt9Lk7kkR9jPB4croKW9qnrSu4MJlQ020dTVTrNKa9KP
9QAquc63/S+KHzj9W18wZeNiGd/08pSDuItJCE2IMDP6hPUr5xIAz5/Bl4R4vA3qrIinIp4ISpDN
6Ctih+uVA+zcxIMNG3Hs7NjNWge6vvQ+CvlWZndqIPhXy7r7A3qj1NCpbAHXx6ERt1KkUQlzyjhN
c+K714wV6rvJG3mI9UbpGcwLllO5q44j4OyjhX8rdjrrHRmi59kh0xViMK7WGQ+dJv1Ti+pt9A7i
PVHLELMMv1DQCi/M8kmLTpkbSd5M8I6vXjx6S7eCp706eAWrjD13FTAq4DeCAYavmXHlwE9Bw905
2bPyw2Qmb2wviRXvcRcfh/Z5Mcr6XgWm/eSHbqpwrPQcAZ13Y03LSQLmbqCfp5wpQwJkTLNEUL+B
pRjOEWKFE1TzrcCTyQPqmjrtRFbtgXMjSdTeufHCLzTW0g/tt1aFvW278IvkE2Q80Wqa4av9QSje
gOHXQKKa5dlbHQ1GaJWqRrZkOapW0ywONrgTR/GnYz+qyaFn2veNEsUJVZ9/z/xpRxKmfMREeU6F
M11ZTJ9nnPVT2b1kwXzqCtjsEfWVCZNYGv+EJONRA6mID4NG8mw4M9+YFdUiMIryMQiDf1CJAFoj
103BdewHsy/C3B40lSXIUJD1FRi6uxUxBGu4UZ4MpF5V0hNCpoTx5u4ePNcVUF9Qr69ifxEcHS/t
ZtJbt0rYVPJxXUsRR3cPS9jl3GrbqMaLS6usSXpkYAB8bvzmR32TO9bhHXO6oiF/Yvnw27nCO16l
q+lW2r68huIxQaKgHKa54aij+QEPUzERD5d9KdQ1Cxzws1Xp6Tfu6z/aLytH4d8cwNYMnC+Y6+V5
0A/Q/fmqeTC/mhfqAR0q4Skg+Bak1iUxXxI5FuG66dUTVfj3qT2y0mzImfHJC+mE/WXXebjbgSMu
nalGmmYnn1Otopa5fKVAkjpUp5W5E1y/pn3gEHxI1iROPRLixazsTti5EJNuIWY7uLV10EN9WWi2
Rz/kkWG5NzMgZ6MyBn/4tFjE5qJVQeKLXPNDcGr4SFTo71q4jN4nGf/tNhv1sUE/Uzebx5CrnA6J
/ZI9azLoNmMLgKtolT9EvcUeDF40MTly9CdkEDmW0+EuGLJrKIrUjB/6QPp4aNcThfnutGBxSIWg
cOJCoX15NY80m/AtkXUZTu5u6CyP8BMiWlP0pXAv4Ga+nqPIYNj+g21UefsemOmOMjxa9dPBqLNY
KpLD1fdJ28BNSZBCyUiNq5QMBR3wydh5X5mVFGLQO+bR8pBCw2qJvq4ZUo3TwqQgEs251Q9v1Fjh
bksgDbGANNXvhC/zlh089XdWvODPxo0t6qr69S3C8jBGrVgLDCn5mb8WYXXu7+Y0HrjMJeebkSAb
La6IG5yIp7KtfaQijBHGvQMd+RF//DlO8a5eQgHevNOttL7LQdjHi1UNyjk9o4oi8iVzF575dDvK
K/iTfDZMXbgj4d9gP35QHR+HpJO4fTkbWwIozGbzdbUaHPr3RO3ri3PEF3UgBT3lamcaLlnoT90G
TR9YqYkkuO8etf9LWd4r4HFEM6JJRyVmvr1JajheG21oG9yVdLwYfF9c3uj+0XMFasmkeSnDfU0G
85Lsbs2fTk4Bv2Gp2ThEFxOZmxHGYlHHzbPv49LqSI6FdBJbHqCAEFXXZQ29EXHFc+rFc9ZwChbE
VOlofd+yZPPAREvoeeKeyzoJVqUOhFv9Wu4l1nUS7IMu1fX8PNHIALAXzfzZnsm7Wf9SLV/6Nwgk
shzQQTxVz0ae2xFdEsfcOVVOPnOyaHPhPhIDT6K/cTLKvE8kPMizRM1QwnT31YHf/CUNVNspL9Oy
AqwT1dOKfeYi2ANfVLDsnn1ygRvfFajtec28SQS4hMbMZX3mB+di+N/b4Vk2b+yVAvDU2o0XdlJa
mfHwbcQ8E4pBDwKDUCM6P7KHsNqX2ZWqzm9WsLE218YLXW9bLLoJOhXLZ28o2IST/3fTxswAIS6F
5xl/IFTuzon7Vj7tpMQetlqsintjkUZjJjBMtiNBg1D/8nyIkBoaA7t8r8r0GIdpUmoDUNmqX30m
5xyf38n57asoPz7jyZN8cNnsyfRqjfM2Ia0VMpfMUjrS+sEeT5eHFSYGxoxaqTjg8WyCcmPFRKwv
CNe7+6E8MoI3lPkyqoZJmG4Cv5YLq61xnggDS4wrp/Sr7ZP3nRq0bBIJQi4QjId8UXey2AHGXQkc
xntIAlVs8RmZlFKtM9htAZDnfzNnUsp+uR5AeqV7zzotGDBvmaZbmoTmlX8t2RLXlA0y0bbb3BCE
dby6FYcu6s6C5xNLybpKs5w8BGge5tbbfXgaROztUE2olw0I4AXV7TC6Bl2BWFVoufIgWxUAiYBq
Z0S4Z5HC89BSmawRJm8PA2pHpWbHCQqoZvHvch4EGaNW9MI/dQjO1EIwrpl4mYIlGtRGkjXMUrHW
fzZQ8UYZ/79w2iupfcjkUrHrw2XvUJZQDb9lCAVISN1OoyUawr6BFwplAuKOGipz4ByX70F8lNkk
hsxepCTkrxhVa0METqYftEi+p9hcT2Cec+IbX+tqoDrt6Rp9KPVo4ARAeovC8DUwNtUml9/rzsvZ
PsW7qxkBklt9Q8mf2wJ1iMqi7e5h5rhh8/Z+UyG5R8KgeQW8cBrBAHeSCI3Qtmx0Zo34WPyoeqYr
LeEhYV7+fYbLNfb2IgbdCBINAIdc2jxO1SbWdTCOIq7mS2K0EliW+yJmAEg5+/lIWoqbkIilbiCW
mzphR9EscErSLYiO2kD6AOLF4l3r4CMEd0uh+027zAwG/PEkIOlpyfq5VJdmSHGXUICYeqYA4Bpq
qzfGpgS1j3v+eFE/yZva9xsxR1nUti2OTNWAax1gQFivm2u8hFILagsAa0/MDI4p/RIRH+qmmtI+
rotRXM/f8o6UkjhpyByzI2vSXfhooWBwyTqRDdu9Huo0fudxXVxh+gJC0FFoVOPWNekNYFejyXc6
GnpwHuM+Ke/mBu36QbQiiZSpRSsV2A7az750g5RFWaJ4ri6vYFpDYxQVY43rcC1WjbVIMAql0NwS
rLJudEFXKgdpQFNgHZ1HW539NA9SMxdiMfg3sLhLM0eOGhQtkx0nOEg08fTVHvfK+6f9P0SktqZu
m3DVNOH2SxW97Wl5/1/KCnNg3te1iMp4xhwm0XsY+g83RWMy7XhOil9dTmKmZEdhebTkpG0L+EH9
4mSJL8gR3w9ClVpZ+oGvIKEqChHletdq57FJ5jcdyzv5vL12Ekf6OfLMauerNHhJwPhpuMjY+Y8f
Bof/0qdbdIeekIKREcOPS1f6kBG4RytUZ1P2Un/0z5CkWvJ5mtTumb85Kv+c1n5pkqrs/H8Tj0Pu
PA3bHrlqAmLwCVHBYIqEj13CuEr5mh8ioZitkn0xu0PzRoa2Wj+We8UWon/dj0SixJdRL2rP+meN
WLjPiJu60LNlIP492GMCsKkrlvuA9O1v2jVR1Aa46mPGjFOQz46KynF0X3Bhk1BCgswwmF4evP5r
s0Fg2a7PT2ZqGo6lLn4rwiYjX3gyu/NTkoEiXyPlWIkuxMzPcn3ZP3Yja3obuGP98vZWtsLp6046
Jpe9KTQokPmmKSLIy9WyvPRYoUucoKIG4BpTR1ngCpkrQj22C0clQ8FLhljNrueo10aSwhEAxack
/+LPSl5Z07sijZ+/84GDmBVgrbmtvgdH9apHD5h8jpvy5zp4cka846F0/fSgb5jRQgMVi2dPAAju
kM2jycTtysoTviPh//Qs2Y7c94HcxLxjpjYedU73Osvglfdgz9hbbaUw52VTrSsXHMdSkvLy84y2
D3t7zXobHprD/XOWzMQvDoFiRU/ut9wdZQ7OgjR6/QtCRo0LNpN+a6r+/JpJ4VLy0ra60/epgtsS
08A9hHtTxYcrhWRHKP7dT/uTjyAPV7lU8ufw7r+68w8rxSpcQQozKFLQwGxCEL2wVGlcAoGY8+Dl
k8DcvNO+k+VUwQbMgkdU6C+8euAi9isZeHSbcgumzQzdyRGQcHOmW0FJ3H4qSQunWqXP0x5YP1ns
dGY4ctQ8YhfvJhLIxx69w7m6QZecEJvUA5egY2AcO8vQFQMat2zudOY2MECYx+BzMUIUOSOFUI2O
3LzDPYgONkQmrTGsygC+9ZhX66TafaiCnec+gV/f+yu9UroBuVrqC7nr95uuiVWHsvcqD03VwhCG
JxAmKg7GbdMUbBUE7ep9J6luXZRwBD3CTYfbj6PUVyuMPkrZWEY/Kzc0i91kz3Z+tGuXscMLCx4v
lKObtXLaim/vnywP8pDc6pTocZRry6EQ25kxtpyIOpHo95J2oKaUE233IfoI5/yHJa69ECdvUHNM
vqJ1K0hJnZhMNyS4rmL6cgNZWsC+JInaqnWq7JFAo6o0cDqVWBUGssyQAOos9rNTFH8BJssYH//p
ulvQtSmBSWWcaQvPQEFz+tIgTFYaHRbp5EPhsG75mim7/D0GkA+osGAlHbrjb15zkuumOPV9950D
hNkWyRmYd0YS5DZRcuQ0nho4HLekf8VEj0WWCgZyaxyr34sMR+fol/Pxs2ST8PG35XpqJ3yeJ1fc
jEpTy+gILrXL+1ELTkz03K09+Cm/gz/Z1O+FjbNY8FSeJtPVUmxEmr8orIILzFttWsPTkX0Mz8Dp
3A5cxZeRQohMc1FLNF9XMMz4Rl6q/edyhiqrmKoVuJV1lUGlLSUsxg1P7lDCOeMECBWZOGfMmE7I
E+/uaA3/jjYkzYhVoUIiOOXC7DF4SjLooDT5vVee2+6X0ulVD5fmV7BTj6kxVUuDPOSuuOZyF19Z
pdicfJWRv9REVhV6Q39oNKfXl+mTNDbGjyMgMYmHW++Xj28vHM3NNrbgWKi1iuSqfSioIh7yExCa
O7fTu0XNIT2Tn+AIExuzG2+k9W1S2vF3g3QBEUQqSQnvWmKE7DHWhKHUSHW7Vy4QEVynq32ywD2G
gk795Ffijo7QJHsaVy039HXA0LaqYIwrq5CCA4AzpQQ3RwrCeVFakB/rCAytxV/StsB+AXz7ie5V
X9OTEWqekEQNOWJWElY8VzwYjvKzaGRRa6hR1CXEoZvWZ+e2HO+2p/QzijPI/mRxJlhPK7Zv+ktw
iEvEcXqCy2LbJyV3yx7J5hFQpgb2a/v0Y7enlWdvwKlEkozCqc29DLNmlme1uQtYQl+g2MgRF37E
QCyJxPtf1DzlyOUZge/xtMAMItjy8ylXFtxKHRmlxKBgOfLU/Y9AS8nMP5uHZgQf6qsGRTJbr02q
usG2jEAC4JB7CMI8/1cSelW4iwS/TZdlj6WAn4DvAMfbwCIeyDnuuS+mQ5BCVnzC0AO/+SvkrhyI
DP2j1ittXs1QHtSGfvHF8mniWw6gXej3JT6Tw+89HUpP+MHI5qerWGDTiYwKC8s65t2knpL4gTAh
5O4X0WF+JRmsxoe/g2q2qiqyULwvTpxi/MlA04LklAt8KBcQkt4MeHHpfs3mKyfV4jTYgudYnYzg
XSJo8xUM3v8RS1S8nlTQJm5uwiZdaacMx3DBBKXnQlNq0iXAr5ldIFNaUK2ThX3SqcQO3/joEj3P
aW9f0t1aDiOhV8VtEwZye5c0YoqZ/iNXiBpuuh4pkjshoTNFWdTZK2SJykyKp0YI/rlQ/iRp/rDa
GFCV8RQ4HequPml+svHdhZaX1XlwaDNW8z+P9COfox70w1sW3P9mPifdT5U7uvxGFk3TP/wEB3Pz
cGqBDTijPHyCymnp1L4GlO00x9GsSR36ZMt1rNg9snZ3z/TBnbJHQWTh6Y80+9OkWBUJ0EcU+1Ec
m/jo4ZIIZn7K8e+d1RxJ2iAryhls+tqJWZjaY5jvTJlD/n0P/H2bfds+dUA+tZKeP/pCkzSts/0G
KqDUWXqajsI7xWTp7ueIGfW82BNMgULMA9FATHR3GQ5qpW/Vahe8rVUyYXcoyKsYJ9WmhTenVAW9
5HG98iVB3qAsXOsyRAviPy3EzyUEkBTfmndSYIfmYyCbNLeOHUWdqT5gTl+eBAThuZbSe0Q2UoFF
ZnukXIoM5OprqNBt/quhul5FKIJkRxHglWju8xuMNqNl/Z/bM8sIPhiVnIDZWcxiwVjK633XiPdN
W6AA8DX7vjwI4WNDpv2hxINuKORhWlPbj51jHLQSq0S5IQj9m5rUtPKgyYk4mmWy2onCiv1zbtiA
Zo5EeVK5eGmvUjJPdJM3oodjztufLAtvgiI6LakfDb1DBDZJSTL/gsdckaRmHlry31kkdYw9lwpA
72+kKsRjdKmJyfc3vLVT335SuuYQK3xioXur9nStTlZmt9Wv1GdKTwRWrRcfTfxvt5/vhW3FImr/
WGaSziM+1KtJ/GJxmvFK8+FdZEoE4RP5b6fGbhnkAwUbpPrC+29g+hL6pZ1ynjSjwopNLKYfHbe1
sHkWz6gjn8lig5heiLQzbj8tkrfPg+H2CdBfNGb0tihWxU+DZdsbspUdmWcdlc+jkfHkfTEY+7xs
SReWjxLy53tMrhSouRXI2oy2ZEIZVC+zMz7rtpf56w+jIOq0sjInOZ+m6yhIPi8CeNdN1x9E4lvs
NQRiivncs+rpHw15oQJVCysjdNwdOm6tssvxF2Rkg920k4Xf5hBQtUFZ79NvHD1aHrFasekaYZIr
Zy3tnGZVhp0u76UnAfrHTYX49RJ1nH4GCmv0vGz5UsURZlVz+KAj0MvHcFQriGeiK83xresEGntr
9V4UUbjSyPvp9aAgFk8d2SGqAtha66bhXv1Z6MOCnEvPlyY6/Bp6B0kxM28acSSG7goRlt2yIRD2
Zk67rJHBBvmVR4hn/Ikuy6y2LW4R5AmyoOhIdnYCIejMz4wiTCOoYKWGyZAW9r5xkaQXtnwuEXkV
njQRDT/SbrY1jK20KS0mKwlLkv1GFKQg6msNdRY4swc4JPaf8JmL+UgHuGpUKmwkSlJLT+CCCBd4
j/JlObjTyABATGAN3EM+rCUpp9VQfjpC98F/5FzatB9uuZO/9u5dQoS2kN77EHFuSoNGGpNeupcq
2VvkDIif0tRhLrEkrnfY456rbKT073BkgTIc6xeiQIg7JiPyug1D5KTvw62LkxcSo4acWNUlW8wt
MNYwTuQ0cBfQu2vQEIp8RSMum3uw2S9CONJuYVFkr3rEeUE0wLghuTnxanhhRgbHOOMT+A91mZFU
+j1E3VkNuTl/KNucX0mzaGHt2rGagbIb4acTFJFYv1r0mRInEeIO5vYgg2bTYi6leJ3yeaKaajBN
ukO7jW4kuVztI/r2oaiOaTpQYEUH+9nyI3xVVhcEq7SxXIwjvYBZCRzbCNUAgf4ok7gwTDnaXJll
nWY8CxO6haUjWCZyIpjBQusvDfPaM3xrKnO2s1A09XyVQGEqOsg87y+2u8CR0AvYHag9O3WNWJrD
ArZ0z8sqcZez6PoClAgeROc8KfW6km852HUJ9+/31y3MR9OPCXLuXrzEuybxh6dZEE/lUu/+f0/f
AzVmqnJMKHNhakWNaskxuRRZMo2Ag5Y14bSUTJqOWbB+m07IRTKhmN7sU9vdu0tNkq/+BnYqG3qo
M36UGxs8bfok74pWzQtlrlMPhqMzZrDyV0YIMdb2EE1LQWy6MRbbw+WLjyAp0vhc03qneRNFKRN1
J141Hq2vS5sAByNQ4XzFRRfBYQCBQjnV829UB8esclIHkSuYB1ARWU2b/vQ9BpWktiHhAZQGeJN8
cjJxPWGySK9o0OY5XjeNri7z67NW2Xwx65rqyqAv78kjf+LHsBX242IEpBL+xVNDEX6821ZLHksT
2KOiQiuIzIMdqbjZw3zlJO3pexmSnlRhT+ChptFyDYXACPuP91RE/mxgkpLZCBMAE2pR9ZcaeVyf
uQ9rJTta+wBDmRfybSGvd+vPNwlKmsgV0Pf7DSZeYpL0m/jlytFFlAf8R+F4fiYfBpoM4kD2HEbX
6WzADlXGEa5tk2Uin8T8XAsu5qwpnsfr8ZE5O/kpsf1VTC/42stOsL9PK+Ilbdm+Jfm/Dm9uk6A4
yd8sEkAfOAW+A2P3Eywjb9JguBOexut4zfMtaudbhTUAWIr1fW+xDf7fr6c5j3eQpq5yqwuUn1zc
TMBZ/59Ak5ufDG5TgmV7iw+wyGfUIZiLNtnqFbxf/EssKPLS5Evf8UEYIigbD2xi1NkF7DCYEtgV
jBVtjE4GU4areZnndetDSc2GSSpEuAXIm5HJS4q4Ja3XNemGLy2psuZnvoerV4XgfRXGbEgJ3IQS
hcmtkoZA7NS5yDNVQZNBGizEWu/IITkeb5Ms3gD7hRyF37qAcXQGJLdZlTU23nco2ofrstC6J6bY
45K5f9KGpqBmZdPWTD/MBPS7HkTyzAtEKUG3+XcQVxK5wuT1H6qTKzziqcjx2KZqyaztQuap8aSL
Tb7jcUzBLqXtwmiH+PC2Y/pPAxFZCCyxzkUaG36imbTm8jUXXn4CiEOHk5iLEznklOICCsS7UY6T
HzlEa8CzO1Ukkw5hVR7kn30h/39RT4AOLSlMwVnEdehf6IWx3D4MqnC0+dV//VWwBj0ansIDs5Kp
fC49HY3f2ykre6PQ6z4A44u9a6UZBmMCwsFZH3KlM21FBSmXo1FsOaCuKSoFveCHP4Dbg7WKH7gQ
7wMiC3hPF/mJxADK/pOcqvtA6ifFQzOpeBRWOsJN0i+NQC8Qbp27MsftlIDRp0ihp0w1Kd2vZ0Ds
JOqKoo7NrsGUemBdASKbnhMD2YxjQl+GbFR+q8T4f1aUz3OMBqP95Ra4u3ys/AURN41sT+5zsxNw
5B2e3+tbLndhyu87HSqhk1ZXAugIMbcw6dqMFkX9ybVrm9JY+X6ZoS0pK62KKl6YaCofUIAkwt3P
5cU2HGp1SIOgf/NCfDAZqcxeVM4s5gaNKLxLYN0a4fthcFlqbWXpW1Yvm0mAqMLFDAMCsl2bRqNh
ngkq7zYnX4cr7DI/d/l4cg3MifIHb1BJSVOXoQcWhWl6aizle8veNqIFUB2lh1DiMLcNd21Fsawh
bNjLHSl36L0lttFeHIWXwC40QiHMY9ShMQanpDlH3ihDMXLqVGs481vrkPhi/Y7NYEtg+mu8eZ2A
bVmHG08y+5JIkGdBJgxqh154qXdltjeTnXxccsbBZ2ht9SpnLmagfXVuaT9gfvkyI9pVRt3WcY72
LbUb/rysT3bB9BwqqBaOsFkkSx+M4Bm8b4aY93h7DEhay+GHujwdf3HO0ASXFP3FGaa63V0rjZgv
KC4p8gN6l9q8pPuFb/kNJRKQnHC4vFLsOyPJbWKEUgq06Z/CAvmnqcuuW4oESxCxoXchPwqj2Kuf
lY9mV9ccrGGH0c5xyBBV2xafeklmoDmPC98CGNFoWZIGw0ULWpNWSPEHg/uhNC7zmP7xU6K4SqDb
21tuzww2QwqIvvEClvPHJC41/Kc5NVRzAhPimXRVjEoewRXrvqgLqG+RMyS/H1S31ZHQVGwGzhz5
stvTKDJsUHXYv6GgSa5db9ezR84KfRt5SNWaNKCBOokLvBOao/jk2btQjzCL+KGcj8bwJw/LRccP
xP3ySg+GcpsFu//S5kYchm4xy8l7J9KWL/tCpT/+NEjLnFRXsc38jlPUmCKgbiOAKp7DMVd+1KhL
HNHQyjfwwriXxUAfvuZN/+4PhiuxMGEW3MmGZ1kt4xjGDG3w9QM4l2+TCw8HGW294KIrywdP/muh
2TgBEzkzTY8bJ+SSZdgI3WrlBAu6QZ1dz2xeawKBjOGRgZ4iljfC333N7OBPIX4E6ZSCRVs6HBwu
CA6j4hX+B5Bx9AkrfkiBMmeKRkhCOGedKTBXOFmRkzbKFZutosdP7LVJzaETf9kjIVPgAA9AgJfn
uenYISyXIG/vPAQaNnyFtjoLP1aoVoVCi/oDX3K8tUGL/N9F5FtiC3t8T+9/nQIykVxCMC08W03Y
WMQAbqfh4xMSa9+xy+Fa0TS+2jAO26cxOHGNvsNqXJVmnb8MwH7zekwwsTpK4SpNum4J5082eysf
kuCVWEAC+YVsIHEg+ICrABfG4LrmWo3576tKlX2rObM4xYxoLYJ/5Ms3PVE++Cw+zLYY3PBSL8Sq
+KM8WJ9mSFCvdcsSoADn83zC56c5VlO1CrkqoPsPUSGLAQAMWvwgSN6vrfjZu2ssvjKsdRXcCpC8
7+Wk6SKbRKg+fWpv/Hdb9yuXu7lpH8MrxKCvrwr1z4YQJ8Noa6iKE6RAUJzqS6GLkQELEKK8MaZl
L/3fMiWyVQOP0cs5AJVGcAq3/4R0QwFZzI4dSfpKXsi4am8uaQAeWhVGYpcKSN65Gq+ilHz9NcrB
lgfCtQL5VG9nJ0dCchY3lncapY0OY+nWcvqie9EcgDGD9c6mP5WXWoMPFEcu16/bFfMJPCeobTm7
iFH1jt9jT9wTKuyaUnfDdrj9M/S2WCAqlhChmOr4QtjjjnI2IDWQcrnUgs+kaJimaYL5vD+cdc5v
KVvwVnaoF/fY8Na9I1NJcPJ9zGaTFNA3zap61veSZ4VZZ5zgiZcILEMLcz6/+2fCUEjlxRIgTyqD
1qMI0qK5VYg2kTX1y/vf+n/6V+govJhlHh8LShM6RYpuTGW7M+EJPLlZfFiQuMwyWvzqgsd11hud
jn/Mmz2Hqp+WwImNt9sD7z36L+EAc6HuxRk5tM+qbKYwPTRjXcefZ3ho6ijw7TDuyraARoBBHsb7
IX6DHXI+KCKsAztXGH8evcJa/lAdV3tnbELHtJIbqflCozQdWNaB5izGsxewvcEhKKkos0To3kM0
3sCPrGo/lOsc5O/2meDeTtGiwhd49BwVRfLXJH49J1hCIne5gjpEh8DCFn7N8QpLHZHew9KiH0fH
R5gA1ln7+HHaQdRkQgywZELdp8IYIUliFiz3lEh3U6OSrr6eaim6W4NL4H3S5wmOQbphIvrm+ieQ
2+UADY+4yjh3h6EbulWGB2xXB0Am7lRKvuHY+zcellwRnMMxlhweoDInOh1yp/LSZvCmxMZYWHA5
g0m201KGARxRvkpfDUEPDSiSK8qkncNtJfgfjPpjSjFhDeMR+23GApBTGaKFPiNdI0xzYX/Mr2tL
4ekVuv2Y7tPHWeLuA0kfFoI0Ly8JD07n+/WVppOtW4JzmWkfeGao7SRipAMOCKcXynk34QgNkeL/
3OSaFSjBBosutSUGKB6CLtMgZiBhxjiv7y93hLHlKQrOft8FjeYnl7iIhkFRP7RmjS355SU9aY/Y
Pd0QUurumI8dJX3po0FZVOpmlj9lfQHh6H5t4nQbS3r2XyPRi5bNksOxVwsvz3nVRybvhQWi6gp2
Y0S7KVsfxzgsbflKyfkcT4DCkRHugiHxjlQj6Xi2C5UlLCkd3dVZ4ujbmc6N1P2XgMZjVhqcXFZg
YEuV8e4vtJOFFFFgRSgjB47ZFPNpuUKZA6Hz45fxmMg+qdCWibz8kS97t23LaJ9LseB0iQcVvId4
+QXBk+vvzc/uq5CroHSVl7vDpc4epqElMlXmHognhdYUW9TushAq8nBk+u7joPypFnP0DcakhKQC
tjii+gDcuH5p0qfKhLYL80mmcd8XtJV3qPIWLq7GClhwzE0amXUQfxmDR8cFQapYoBgwGo2ixl/u
OhlbfFetIl43tIrbKtmLcd/kpY6qETMd3Bsbak0tqepP3A+p8ZYmhJHb1cPS+KIKK19B0e+OIu2O
pkT5dhQCy1UuOz2OJ41fH+2mKiTxfTGK0AUVKXzMfMCYgtPiFw2qA+5vMfMJtDz1681PT70eG0vL
wjVN4zzMadCEWk6RVvJm315X8KZbA2U7F9SKzXzcYbtvjxAaGPWl9/TBuSAl2afPxdr/IHe2mVg5
WxB8PuoPJpiBs9QmeMfJatrb2pxlF8BTm1RnkzS9jOdAvXEBuZOo3Uiqnk4XOzTS+PLZ5kakLkGl
nyYV8nSfwfhMaCteRMeLRvoXm9QcamjYHNNWh9xwpK1ErC5r1c8c4xJtVTLTTR2myG40yNpMp70D
S0XD+UodHI9dOxo9gzFOfrvuCeEwUfo6DHQPK0QAsNf20aQLCo5p7DnyzxToaVfGwxO9eHcb0Z+W
Q7nhLvXImqsLczJHBm7DeM7PU+wUEPPttpcFnkgO8dyQZdUZxMqXzCMsX5I7OU7buxqHJgBE9IHF
F71UWIOyo1XF1dF7w5L32of0PazJUQNRFn2fEZVDcqVb99+o08/vPm21q7qEtld4lNUbzvEpqUwe
SdK3Up3d/RrLPyPeYMS4gXLh/JAWu8ePu2OYCShTu7Gc0HBKoKOhFz3ULdeZd5whBvNJFCYY9kGS
B49hu1DpElnoGl2tJyNVNSOSyYX+BLwTzi8SDdF/mWBryinOsaZLIuo+kpQqVneQRRYUeFjsxH3I
96W7kRBYjgYtbb5SS6F6iPuImSqp3hwBQkSOaY92x09rkxxFqAPCUVbAJMBcn68/TKrdcdznyj63
ZL5BWDThd8oeEMb/7yTKZXES48eJyc9PneHPFT/vySf+g5yVPya0rS2QqPguqVmWVEALRNqso13s
N2Kf8K9aJu/XFcJnWpe0mB21qijgDfnu/MJnRoZCqmepqrPbRyX6vRjhUb/TQoEztMdXwZb5r3dN
f7ET9WBe9vWfzI/yYeXo3JRUGqLX8thEKXJZRoHryiUHbbmL/tm7BN9nqPa7SV4B0YUHmy1V8Kqu
6eiOrW7ohS1/Lb+tHXVNxZz7F8au8HQaEJ4rcUNPXYPiOJbx638MHgCToULI+dZQ7w7YzfaZMdj8
yUxisKpLQFY+Eu9XUudImlQejGfrOUT9TnFnuVkOBApz7S6X0rpxcBi7RtKIN9YQYeT9UQMviWej
hDXks+WykeEmoD8S5iljOlkmlOEhYNp02NjighWv/uBDY3q7SA16laSFD0p02vWI1clbyNQ/qif1
rHVnFv+hmoCUPWahr7BZ1yLv3fxqDyKsAoTsG1Y7/iSJ1xC/UmHfJ9R61IQN57d/1GM6vlE0R8f0
dhh/YqA9RpnNGsTeqmHgR0ZAmLtGPp0Cgid3G/4XOSpIWKoacE3wd5r/BP0O8c+wkr8Tli0bSuWg
0dtCGvGcrq1/Y/5Zs1ZeGlGwPkTvn96nZZ+TEyCXn/EB4mXNAVrrVwGA32Dvy/Kha1Reci4VNHaW
Qz9o0hqqYvqp6IU0ZmxK90Dj+3E/+t2bcK1E0RSmOC7gmnwZ6TYP4+I8h8C2IXWC7PhkSOamHwvb
c2wlBvneuJhMWEwHhVqIX+iqyT1uWj59+WKm3e8eHeh90+ti3BOW722w1/ONLW67yvUoH1uUY7Io
bg64pCBw8EvDu2LJF0C+oeahTCEmdBqLLEDSOm0tF/VKG98xfsywY8BVR4SoQIqit6IaUUjtErW+
XiCU1ID/Ebp21+xpSwbhmxZpyAuthDL2Ro9COj3eXFAgs2lh+3yCo81qDFn4h3+KtQOU5a1c9p/f
SHMJ+3aeLfYECmE1ryLMZqg5TGwqQhRhPwpwI6GyNHNnmA4FVSa0/3fszoP/JrXcBJ6Y3gXI9Ynn
cv1LBhv2fJKCNyLhaEt374nDwjIse3tUyyFg4m7COnkzX7EArUMkb+jZSKu6mvb+p0hRsgLPA9Rt
rcAQjuXKacIjYQM7gEMxj7/MC/Pc51tGV7rykFKY79xTeMNgA9nXId5KSTA3lu3Uz18EfbPOX7PU
01TdLdEDFmXHbpe8LwiCvG+pKs0tMSQWFfm0Ys5BfIbQ1CL1vHnC6K9S8qqZalQXXQYvHIy8mWpf
hFfqQobkP7zgbUOQcIkhcUq1x3J08us/l7KvjOV067ZK9dBCVufVtrGelokt/xnvTCmY3iOy5zF6
Bwkm0AwamgugtoaCDP5NNkSi9pe4b3/cHdtZj1JIIZPXAt+td3EK2YzVMofvVhr4cIB0iiZ/kHwW
ZmIlZ79jt/s7eGoaOgZRZvbnwl8MvYIF8XwNjFmPEaHUpc9x4hGGeI332Kuzz7Rw2fqKZTzRlVGd
0EmtUdHi79wLJk1MxFHwtiPBTlw3Qe+tGsgn+cb73Kqv/PDOlDu5DSDBx0VFptANvwT7DzQdkz1J
RZB3paIyRxhR2DKz68/ZDx1WrKTqKRpU/CUaNo2QZN3AADJ22nd5INouK8iy3gFxEyogXhAkIKoU
g8KIHWrw79/mavEI5IZ5jaoqE8FsccLkSrEuNIugIwBaNqhH+4z2aDuGaZw4fG2Au/3DCzzjvA1Y
wOwbPaUeZFbt/XKLqsDPRziEgKXMMfvIt4kEqs5awlmSnpSao97RSTUXllp88EBwnZXxTDrviTvV
IwMwI2E9xNWqBcdAwE9HAYKD7wtBvEnGgJhkoxNjphpeLmguJPPPNwmWmnjx371uQG9B0fkyeEhB
qclGYVJqVdbYPYJuAfv1L2s/TCT6MtG7e/IrQsaUgrOxtfHn6/xHyex8BDBtryUsiW0EJzaTdEu9
XKtEV3yn/OdKLSgwC1UAlWx8iK33n2sNUEPqJiAvCwXGo+7C8x02E09h6GiU3ktq+p0xmQDjcjal
ytaJNwMhM4Iyyp3Us5iyrQEc5MDTW9B3nEIVNZGqBWwAbueeGSxgNXKs/bXWmy1lGIkvi0nhl9UB
ABS4z+Hs6IFj0mHBsgUGJsDHPHdWYu1vZcRRn8nVFTc4MFYlrQ143R2lLeY5ShJ/hgg0OFZCew2u
GjMZOZ6DyeMWJlZvZHVA2E8819n6OSYsZXrzFG6Ey0PB59LzGzh2LLwAAIYMOf80UkrPIZH2MWmo
YlU93hMWPkEa3g7FLiYM6LKaGPK2sKZ0wkMAzYBWaBeHvuVJ8WpBmcUwlyePmUBXGZ5oULFjA7Yk
3T46YlGaTr1bBntn85t3zH84+AsbmZhCTZpcNq1KcPPJ25zD5yLN3LVJFGQdnyJHQpA9zFgbcwft
A1M0zF1BVpRheCVIdTSbssP0hK/R5+OigIRKj3YuBIfNcjvbJ6X3Yqa0JZp4p2IS7zu4Z7Dw4gp0
zev1jHywc86keOuhtORpoCwmSofUo969o8m9oPs7aRkhqzZlERvgVblVIJnE408185O8Pb6wE2cn
a76E5WCITM76AQIKYNdDPPvnxOn5CNgGJgZQBpeAOwznXbEXqGRDf05zuHi6NCtuzrVghaYbx28+
AkkdztZYTeZwIib5TZj6ckvPseJ5UFmcA9p17zFnhXeD+lY1Md2U9XP0V12WVagjRIe6X45m86AD
y/RcqncWlEcFZZG7Y0hx20aKR1YpdonWVpY/B+MsxCwLqmM4hpumscCOmCa59819NZQwPg5W9nRX
YwWZK6m3JzE8ap1ic+6swGcjQHssMz3dtJSQdCj85Wo8nAH9HoIaODLEz4dr5dE0FruYRIHXAdOc
t7kYnSvR1ngBNPVJ56Vb1kFkpAq5Vy65Kx22QFz+smh0Q9G4orAzqLEpzVZR40okyywlmiAqKquX
KmP6m3Tim7woojQqEGVThli0e7RNVbBfRDjicSEc5wCN7OT0GMyxd4ZjzWcmE7mh4i24ikLsO0ME
dS4c7u8AXM6Jgj287vB5A3xXLNUp/D8ozj0Pu+ImG8L+FZbhguWG/AaX9lAhF8OBM/2Eao9R3esy
0KOhn9G5dHyBnEyOWpJRYFzbw2RZMAUMPKF75d6xsVyx2P46FsH9T+bwvqAsWtM74qAKX8Bv5NkP
/SWKwrEttLhb5vf1XCn1EEKF7rYyWzQV/UXkcCLBd2ziLkIEbagn3VFt0QJZmBvQvlfuAwUTVSU1
eC8gsy6+WXlF2u/uW5VOL7O+kSyY6KcMKNbVVsr64Vxf/z7eMmlcDVtvoI3eVfIQGQLIPpn7Z9rz
XiPDotq/riCLrPb8IplyD7XLSHLnqHBuAyjMNMcUJbXDbs5qIMzkC0SNFvYenZSqw2qZHfekFYKU
i+aP+2cShCk9yE1E7t0CioXAjwSPP6mVJrG0fRFpACMukmprbSqMDl5Mba+0oVry21GJ5cHF5FcZ
85De5IGVuiZrPZ0PImzzRAkX8ALHwHZLxGQka5+UIItgd+jEqT6p1bUoZAriXgOXMFheCBZOs9IY
e9HdCMj0kG2qznQM5vWSNDxPv3wX/ODX/f1EDrMnWXTPq+qlM7bIDJ8t3ltquW0/xewmG5pIVTNj
8RgkPevxlQCq8Q7GK58U8OTmX69lA8lNzIuA6G6XeOo0aWtOuLfPZ0sv33E+E8m5s+BrdWKDU4gn
OZGRXyzpWHzNLpbUuZzWzrXiUdg6zQF4yaTFTLV3U59qATJXA0e+g94plYWGqPuLvWBHS2gLYoyT
hM6GMyE7SdqzBU3OYhl8xWqQpEqgwRYVbmrXFKnV28ch9zkQ38ZmypwzadMDv3q5whnCb56uMB2q
BFDbHwFjJb580hnJa88ZAXjlRjufa+v4nDi+ZiHK/adJDChrHZZVVuNTLPxWXVzx9nzszLMnYphN
EfbIr6SLIsth7R4+nCMFKkctYkZ+4qIe6lJYJ0yggmcdZLafx9x2cPI/zXDLbO2ngO32QHaccsC8
dVkLbOpLKEAlz7nrPgcHJlYfEjzv/iHi2ak/RSujI/IVyWsDv66z0Covpiv4D1U5pp9xZQZTgISR
paGmSLcGqRZ8zsl0pJmaF8ePELi/vZcxVOnZlC5RT8lXB+VvDp8l+2StS8h5ga1u3qxvnWoYPL4r
QM/0cm0UymG1Nqb1N/Zy+RJZ39xIAPwECBjqEeANvcYdCRPAelltGX84z4szRAO0egFrVfPTUMXt
FjueT454YX1darlO6QJUtvt+szSfTrn4C1zvyhmBTAx1/uCPwOQ45UBG2LGCGfOjhgwOTF8IsaXL
Ad2KV0oMw+jIkpkb9AycORztkHp/fO3CiVN4Jihs5kcvpJ9R4MVUWpMndAQYzUOz3r9EdGVyKfuy
6OLo36Z6fb2672djnNO7uIa5An4qON/4tqodShzCRYE/kW4jXQZrks122XcVa0WHFo4Loaf1yWHv
mo/1srHg9jF7wULMqeltVoy1n4JgKIWElWo0rIYahwoXmFnczg8jfPJWCLEfLmv8lCo/D93ND23B
HbgqlGLT3OCxnJEIlhaDLt5DurZkVAPRnyhbzW4IizBShjmIsbycvPtorwHSjLA5Co/lCaU1a9Xy
IwQ6dEzsLxs1KR6tRoUVpvtQlDK9ab1Jxe3WWHAd/4ow787+PpVKZnb5vj1tiCVXq1Yu837xEPmR
a9NdpmH7uWMYemtrdrwBZAoaFSqFezmmIRopVcnM3vQRS4BrT2NHeLKWp/KJSyXwtYyu8MDYidOw
PmgF5gOWQbln0g1BJ3GiWI3ijLAxIfSueCCYdEchizQSJmi5yk3iFs5uW4pPbeVDDmGxSaHhsuW6
IlXwwjGzCwv1S6oH0hJifRW4PdllfTD+KkG6B63tBwmufhvzMD+n+zvxXb7gS7iiLDfLuPACwEk1
R5wwvicCQ3yPJ/xZktz2UbOQmWgxarGvaYyh1npvNsXXhfSLOWKL0x0MmDq5r4zYOkRrC0RaYGSR
7EfpNq91qRWj69KSLy4IW5tI08U5AEu1ef+AQBCk2R9d+OETJPpa3cducF5bRsiUVbYLe0KsHW7L
QYlIAtdhJKwRXWrv5RzBT41GaVAspazIfFfdMCV9om9qv8Sg8r25Ga3ncH7pwbwiUzI8J0hDd4jr
VfxZHIkBl0DY8OiFlrIoP97yMxpYSkLEXwQDPll+bwEKHEyIBwv3ZUqDvJKHxH532cMDguv03iJ+
WDdtuBVREoqn/qFQve5tvKOSBq67037m+haFMiqduTDfNtBEP7x5m4Cq6udA/hXacP1rkDrmCyqc
C9lKxh8tNE8CxBHHcL6GyblS+nd6mC07mO0tmAdp5MEABFPs2FKtMyGfvMMXJpzw0ksSva64P6ER
n0w1Gs3SJUR6pcSwTDwJOZnH6+T2GJOadW6TetjoFkf/hvgQ+rra0Ec/RbLPwTjdk/0e8y9UdaUs
ewfaB59pAp5cdbGScsQzZmOOkXElcy8E6SI4HuJfmuG8mUVa7e81Gd6Q1fROH5ritiT4jD96hUOx
94YlH5GMRD4EBthQyrPKHeB01Yrq1+jSUYVl3Qny9WBNfmEZh3yywegs+q4UsR2lVuvWz4u8JMVO
2oDpfyPrYvqmxj4jTJHVymkCFdCrk252iWmPt+6p1/1GUf0Vt3pW7iRF5MqVNzmI/uN614nBmD+k
p7+MBIOo0tSzOzYkE1dmvdW1WwSfR74diII0iMrTcZDeANMzQEOlJQU6kuf4AGPNH451uDT3XpZb
So5fUPoXWGYR+hOtFWqtoy1PUdgzrNl1swCBEE+U21tKPMHKVlzOHyxg6e9u6KSzgYZ+0vTHlfke
q9iJCRUDssI5CZLm4m464BU4UO6YUdi61B7Q6PQT33qEwub63DZ7hGPvwKBEdxiF4bgJbUrSF+md
aJQIX0997KH7uPqlbVjsSNuBgmklZ4fey7ECFUVxvD0gmkXRZtQHJISqPDmZi1iF9gUjtSelN/Ol
qQz/ifFxcPzU4OUnwqeF+QHi4oWuTW7rdq3u2zFSI8IRKA6+VgCT7vnKUbaNUZa2Xb0SK0/Z6K+W
5c9JXZuPicWN3G9UKSECpNnq9DJmCfXn3jR24uwFCp0GE4udOeyRZTtoAFTMBAStCLPaI7kM8FU1
vT4sVeSbEZm7dqbu6eLGrvhV+qYj5W1vjvrzgEVUSt1RxfTfh96cPvbigYeVVIqMdh3AHYiOrajU
1V/YtgD4PIWe+6SFEif0VxPLsOhgEOUt6zh6kYpz1C8yG9+yea1jPfACyGZ3DrTxyYE0SUk8hEUp
zrfzTrmZ9IR/UlA7QOwaV/65H/Imy6gZJysoPf6Z2v4QGC9cYSGQBzLzbnmaA/TaRsIwaT0KvFB0
X9RbhTm5AWDmi5zsVemXeBy8sZbtnEDUVCWJrm9Xge26AZlMBCu2YFOxSL+khPHGcIQJTgyYmI19
CLCbqYeJHpYMvWlHnFDnv04po3WSa5/mfRGNA5smZtp5BYQyn3uF1f+yJYuCEGctqvJUO5a39y+H
nzQPIZvK3QFIzMgZR4C6gGwbQ4hfkfNDyNL2Mf9+oEDZzZI7ccQLJNlToV7qg5h+vygoW8ae8V/1
BOgyQFav+J9Mmon2qRaeD1sA1nC/40k6gK6cRJqZrvUvV3/8R4rDOjvcnEkc5THJWCX0BNDUWQue
ZuT4A8gzEtQmlG3o94kYRt5EprDcoCViSbklzSpjikiP+gpgJnG+d/HNiycCWgfiaYt/tdguKi4T
F9Htz0qWQy/wSmWpXHqztwfotz48vIKjuGlDopT0BEC98183cQIQLgrazurmi/s7ayRnmYzecdLz
ggrXDhZP3COANtwuqE6Iw+/djWX0Mzwjx/l9Yam8dHeHWoNDH9sP3NB3SsoGY4q0gy4heI3vB18E
uMw/Z3RmTi7k+s5Dz/XAUxPhgLBN4GjgDpMhzw1bWylMIOIxp026MoYdtYuoVXwAieVsERXnlYCo
HtgEvzZdps8vLbzlI7epTEbylL2wCVxEFkJmpN98TvFYLC9F25su+vPIfy/nly1/S4EoUn9dMO3r
cRZtjQ0UwSN/rXElFUB8f75CJSUrr9loZ/qSphC77basaJXeVG7QwTUWZwAspGEc0M1UeVKevvUW
Fdv4tKaFB9Y6o1ykdG4ZGP1K8sE7NnUwATQMRr1gBLKdPuvEdWubnAOxBTz6FcV0JcbvS0Yq+D9M
wlZAxCdKoAIPf/K1dt/E8KJ22NSZPDHJ9pv1UXCygedq5FfbsvNVzPDSkiZFNsPdmnMK1pCMt11V
/CTfAI2q+07PS0Bt2/IheRikEfScB2oHdwmw/m/2f+dGmDy6srykvym4SWeb4ZfAEuZgOe1DKHU1
pz+GNsukRKcH8pXJCF72lOCpI98D/TVY38lX3CxvVGtTfe0TrPDvd/CelEXkfXLB5w+k93BLC4Wf
izYfKPwcjGOw7+x7jQ/dxsjcPY8oI8onlW8/IDxeGc94kQaas4AV/iS17lskv68LcPrlaAw7cltX
MrA5uNKQAAjuv8gVtezAMnnhxXf2NnfzvO+LDyFJNlOFDnJTuY4KtQQCd2wvhFyjlMFsGsvM2x08
o4WXuCQW+Ay8SvXItb/+Zfyj6iV0931NJ/OwlMdEeWmYmlKYuSCU8kcibztyfdFZjdfNV/4n0SR7
EqO6DwmpZNxueZdWAp9gTywB6gNYITVyRyXeRXeo3OCJY54cTaN0p37tnHpWGavBp55rqaAs36sQ
Ivo39bAtc/Vcu4Iemz/h8LUdEco/n/YxfZTtuMrc3hl5rVPjiJF5vSA2JZTQSZL+Utx3CQLZSIyj
0GIpjjivL8Yfl2SsSx/w9/VtZjKkcb/ebyYZ78Rlb30ozcu+l41SzDgmPOa5mothACvYycSceZQs
3wqihLnF3Rpzs/ZNAWyNGhc/HMkyK2ib4x7tIyb9d7hthKMvWWbxauVLzc2MfcNvv9v7VkWwv4W6
yiEv+0LYTd9i24huwPeWURlZYwkY74WjsBjRCsNW/iI2jfqp0p7hgP12QedYbd7FyV/8n+PKKwqX
0C69NeKV08HGErC9T5J0lGXi7OGmmtlGnpTtDIDnkrdrQvFFubzAIeoxVwXiBcYlsyhsQEOzyogc
Q/5LOOOezfEDrvqwhU74VfrsBx9qCwiCgara7yW29t8gO2HFucMryaXK5034wYPmuKeX+U/8aiSt
+XiD/dlVC9uJHh0a0+tGyls8CN4HeKEaPnZb1x1yuV69rYRiX+CcUZp3hjrV+U1z3wwZaHluKX0c
ym86O/PVyu7588NYKNr95xWUQU+UX+ybfYHEKdfPZYNDZ+IIz++aYoMjzGk6QO3PrxNOd+I69FWy
XukPG9mPJ5tP1U+OD9POprDqyg/7CAjEg/Q3Mioc9yBC8bN6oV/Czvp8Cm/bhNkStiH2Zf84KD45
b0UNHyyqD2/89kBbj6JCDpjMK6G5OsOsHQv+vTbFpH/nuJCu8u7GksaiV5ZwLuc7Gr+nPb+O+Wk/
V+EJqAg9rWlnk6gbyBr5mGmlORGON5FBFaVdLeB2ogdnRREsYvAQa3vWs1G6YgD9OMrqRwpf52YQ
PHVH2GDoMz259xYTpURe+FrnTJyocGNnZ0W0StOhwux/gqA4M+upIs1/xAZ486SmlcyHtbJOWx5J
swnGnAbbo3Puv9VLVTV/14kGDpSS0kkpLdsofGtHM5rgSmGY/CKwEpAFxYmXhAQ6Nz2RY7kjVrBo
GV4N8baMRACDhfydI8RgO48QVn/umi0bkzRDS1KNqIyyamcMq0wX/C0WbHCkqQmbYML1jcuqlP44
i9+tAfec7Xp2AzSrmQlFF+vuOSI5sM9H71rCqzY/ZuX8jgHW7+u87NYEykyWkCsFe9lU1AuQyI9J
/hiM5x7rjA0cSBFqsjewZozITj7f5LSovAIgfPZ8BXBFmhZsk1y8E2ZhQoUZcqHrXch0vAV8YeQ1
bm05BdIWqkX8GpOIiO9hKFxiCkJWRbSp/Yv2m1bxClaLVOUVyam6gyZO810PjTuBGUi0w/CKWLJp
uIxOmpbmKk3MrfEpSV8tUQb3fFPcU4FbCVNKGUKof5pzQAZPuHZS+NBgv++PEATMxUamupfG/yr3
EKrBjfHMukoAdTMfl5GrSiboV9ITd/U/j03T+KuaRW0sPcFNfi+7bQopsfAbl3uVnxaCxxId3113
bRQWCeCOS3r889f5dHs6A91Z68wt3frN7KsXKZH3grFSxhAFDWMOPZrLEmcclffG9Av7fBZUV+oN
MHp5/hbvOZJCrgE8YVZ1+qD52iua3B9T3ycz7Wp9hiEusQ1wBgRYZ4QoLq93WaakI+XX6gIch7AA
y1DVU+P2uZm5+L2hs7ym+ye9/h8ym+LuI7F0ZMYt4qUdvgWWTo784beCiKApszyUA7aAje1GO7j9
5yZ+gAeVM/NbjKecWdK1+zvRxgRt8yzU0ej2Iup9SmKtBb7SQdEPtIFUTrN3CIvZy34Z7jUjbvq2
zZModn8mGnMSvQxTK4SQTitk0gsRWtz9mFSI/0VgP7IQtxFkSbXh+WKwmhGV9abun4bSlN/f8lp0
nZhrozk8ucGTR7Fy+OYZAaXfB5WJuEV4XFbbWo3V9TJTKe9QlUedIIb7Up/5aQmMt5qkhwPevGr4
Jfyp2rx5ZhbB/sJ7B2DFTp/G/pYjxEIvLtgkY+7CxEu6v6/dGopcZF9xdsfqVA8eAkDamnhHkKZg
IimSL3VCUGXpNwePGW399Z1ckRS2fZTrNQ9yyeqe0tvaZ1MwLZR3u0Hm+OaUt3TfkSx/3F+mXFxq
La+RVAoOekGy3eysWXlFFgmzbUZi8UFL50ZNckKj7ws29ED3MQI9U1NWqDMdJECoSEHSiewCKkAu
Mh4ZqnoQCd7WEKOAgJqezjavxsoxdzQG7yM2ImaTT+gih0NiprqyF+PSPE8p/pbZ7ytw+KqgCJ7o
1usZ+zFvzfJpwvEdqkW7J5+Onvx8iHJmTfj5p2mcBQYSK2XvN1ro6ochNMGzDm9+vZ/TaxQf9P+Z
ytCKaGVyQYL30zk4ysNIwvs5IwG7lrq/zw2s7am6WnIaosXdPRMb35tPVdpwWFB5bJWuuY3qTr0f
b4QDstxgGe42Il1615jwhvs7BGYugtfMKn89LhMBuVR+nUwH7EVfZqs/Ajs0eDOeU6W7GBg6Idup
tsi9GgvK+zcF7xvHtxC/GCSoZQKHKzKouV9Bz6snKMhWk84soAPEIAP+3WfhsN2QUgTlv6XCUSkR
x9cWXhYtEO14Q0ZR+Q4lrBO0QRudGnen0XJvhHFyn3jnZRnyFbKpuVDJ+adXqpgaWuhrrKDOqkb8
ga5U2Ub8xwDVfdRQiEK+1D8wT8woN1gmDZbRiJXroY9V1W3bnbMti5asYPmYtTIE94AksQ1oTt8X
HlT+iumUepm8/kKqu8OAD7wiH1VNDZUSb/vAydKQodOo1i2MW4xAhP4C2xXt+nLFzFTVDTeFCRbk
PIhw+oVzvIjsiMvUeMMkHTnlERQCyRhW+itkjmM4cvz2FscYnvx3G78j38VY5a5QwUXC15X90kb2
pQij+E8G0MaeaYg0BJ8E/bSLCIwdmshkw1zCgMqyhM6EHaMLvBKc5DkBWCR3j3AhNutbwFZbFcli
dAnk2vhXmVOG7VX4geP6Dg6QmPUvtoTrH7jJR8tYWq1XGa2w5lF6cUyEHMY2d1UAZSqQDgVqD83v
zFSzdSo1POCAk/o/2iaYeYKsosR5kJMHVzHDgO9JHZuspQMjv7OXv7YlFfNKVh1Y3oPxd6T9L88L
5TwLerYKLb2w+GVy5+pzGlTS6h21MSp+8tKY6sjdmsMlkiOtXJBQuJ0KCHa7fZCdxC+1m8lr9m2n
DQqtkjPxYhFxSQKZlnts9EC8iF4f5+F9vHBPUXmZhDTzzgX9U+F6cNN4hBdcc/6TY4dbg7lOwFm7
DMj4Z33OIku/TlSFFi61rD871pOTDhtWQTgag0QKMYAMa5cfdrFnUmEkkb93ZQ32GkBhoDsz4bhQ
pEAsvV9WkDrCTJoyAWaZuB+4ilpaonnbTJubLuUyxgqFi9zNRNiGpG++OeOjrLHqr5HPYUmKwfAL
wj9NySwnMrQFSifibG5Kq5dh5sVMf/tgPFQ+KGOTc33IfmsRBsc+zl5yr7x2XfF2TUF+4UkOKZGz
bV2sOwtBcbpUCsBRQbFd+EN0M0J3pTZdznTKD8FPFy8TWxkU1X8n2nX4c6KlBcyjy/KacGBviC74
Me9e59uLKs5gQ/e793r7XkXnreBwjmDM85NuFvMc5U3TaopCdXRQn7g0psiBSK/W5//eUDM33MZx
wgBl7hQyrb2K0BG2o+NCXlEyHnk78SPk8mzEuEfcwjAmoD6Atmuj/HgfcOjg3rmRMssVmmrLXP1e
8VXGlqeQQBeGCE7Z6ZIgUgGXEaMnUw/HDAa3ttekZrld/JSNqWax+lP8tQjtkhBG2yPXG45RqVmL
RrOIL4kR9OwLOCDhOAg0MkEIsvNm9XA2Wd6J6tlZVtGedsshj0X/TeYoSo2yh4sgFZglJbbKig5W
dd63UU9WW6DWMlQzHpbq0Mjc0MI//Jb3aQhvJ9eSfgykZXL0iOaZ0qOkeXBuRTbFKQ4PmVwwlunt
xoSvQiQIDEPFbaNcwHA6dz25K7Kf/kupGBqW2H58MIkyVaY3Rj3535Q001X4t+JC20g0wkTAzWhV
T1jAvEiDrIga8zs3vZPcfERaDne7uSgzY37XU8wZNNcKahYrjnT2huH2kdFhP1TTnoPx4VtzR8+v
1tGH0OCMo9r+OfOcSvbicIS/wbdEWBQjjRBH2TTWZg4mzU85WhjTwp4YnIOLYpVDL5ttoASN7v77
cR6vey9hod2slokzr6XDyUxjk6MCeE39uVet9MnE134f7CTe6cKkacD4RcJYRgnVz2QQpBWwme2M
+V7pOeTjrhO4T6cOuy2HhRHY5j35d2tkKVQFrYGNnUdvrsYXQN6/2RXgWMZftPEVFIyBO4hTs9a6
d++0MRhqn3M9hn9nIvSuT84tFfefGTv00eDX5kqDcpUQ82hrbuIX0JBF0LASE1PH9mrIzNOHLbcA
z+wVDnXwemYBJh5z3BPpOcg3YOYoNVnq75qfapSlGWI6m0zRqNpnCCQgKHucStD5MDZh0fBuDbTI
c8gARxpsEar7a3nbjs8J4rrYPeYj9g5TSwAg0TGi/f5mrdymWIfp/1wP89ZFjFV5sJKGmBrfk0R2
rAz4hq/lwo2gH0WZjKR8hDJFPCJgP8uyJDl/AmMdcVZrcS7byjthQL/xvXYaODdzRrMX8yjeta/Y
c4G/ugpy5kFTRhVLSdQnQLKGKytG5NyACScFR6n2CFvGhOe80g1H0H3b7brrleASa73/HWoCSx9W
JOaqx0sLpTbnrtLRjJNwhoZDbD/RZfTVj4JxXBhUMQlQYnPm6XQkBVkbNagyxKfD8lmrTUc22zHm
TWPe5y9ulm0ugJNvCRoxzpqaoqtdNIANNNUrtLil52CWkdYw2DbkmqqPc3Kgz9jQVawwnX1nKWWc
OenPL3emOCVCtuaOax3cRcDxxAsOx5RTRBF+YSr212UeGjCmqOEoA30k6FZTboUMTyPiiiZc2/3M
Ob02reUJrSI75Uq4z/3pKqGmCW5WASNPd3LnLWbVGwKKXZSvcNRdqCdaATZ6TPyStfF2+CVJ1Ph3
n0+5Ov9pCFQcrIEwjNRxwUHzz5AVkG2EO1YPkcEWGXYLzqi7MECt9gOHFuXwmLBHlVpC+8kmtC/l
iLurvM+UFHA1LBM9ICEzKvp6E1WU1eNGkKj1U4xc+AYNkmqkQ08ZoqamyFyLKgROTWK47V7bWd8o
aAKgH8JJ+3mUtUbjnxUTKXdt19QxNIJtzcP35UpEh20arPix6B3OdoAryjFM5QCJfMQHwEzhDByS
gp4Wg5QhCIKP9khx/0F4JCjaAJ3y9vYj5O6MjV6AuPkZBylfd1xgFmb5yDaPOVLTKH3VNOcQOrH/
y4Nc3it2suYhQIMX9n7rE876nSKCzkz9UScGtswQK+32+LDko/wVoOJlSJYT3G81gwCxWVMEpgpG
3eTTc8G+emtynjscOg2aEozAc7zHLSAaWDvYtUmd8Ul1PNDn8G2k6TD3RRz1Osl0wlxbgaZ9+sS3
RCI4AR1FTmDtBeyUEVGUTfw95t70mBtZWtoewPot1e8xeXpaVJeVK1/e35hoFCdDz89s1ZZGo+P7
ZVISuy9/Id16zg2iziInMYlkDCdyDgHOROy2JLgkuinKl6YvFF9mt4sXFfHWIAt/VqNRtACtBhA9
LAzZASUAxDUYNJc6yXIx16CsI8zfcONxnJYh7Vv0sGTHE3qH9l1cy9cJb3u81GtqSrxUq8d0h8Tp
dgrg4bgxioK4a3S5l6YcLaGMmCt5DpUYiMEHdvBbAxjtuqbi+wL6+fKCHuewYPoBJz11Q8Qb3UI1
UmumK5PxGgtnrWXY2tskhS2vOolALr8rkCqfDASyzgn58y3uDKt8+NaaE/BGxOfgv1gsjIC0y7eg
kT0hryuqP48HN3xaLThK7JYlDe6kLDbEDhLEzR+xAWl+dtFwcSCqAiCUfuoPxIXLQJITd/bYlrRB
T9NBXSyvnaQZDmn9AqMX1Nvf4YAUt3khu3CdQdDCcCHydq1TLnSraBrV0TAeVy2ZZRlzn5c8RWmX
2LRcXWexPIZGOk6y/SIkg97YaXBskHLuej5Qg5sYy5u0r7amhThNSdMqhgw9jWrH7hui69glB7oG
V4LqEru8yW13RoSOe0wjYuYJ8hmUW60rFZhTodnsoZ2DrYTz0QF9ia0jnWqPm0QkEym4wW0hFMQM
uXcFbOU3GjqaHR3jCU6CSkNnwMY0VvU6Iil9+iLy6lTHUm7x5D3ykTy6KX9ti0aHjKuRaW2vSoga
msU836VyFHrE9nWdENh+jqivUBGH7+9Ue75ryCIXKecJWOCLlvRNrYL5Y9k9zbvdTNDI/ijbYFTn
CKg3AtW9N+eOItBVDCypsx55ojFA9a5RYFeMleFDOtuDEFOAUpYZgn0n1ByDAkNhsXaans6M1F6L
NISHtRIvqAakdcImMRGTYg7yLoGjSe1AeqdduGIMrbI6SHr9+f+U+rVRMEafdvBQYwWCg1DTMljL
uRoHvsrcVvgNpPlHcWa8Na7OKKDhmgGP1CocLij8z4N7kqB7aWkAn/02Ai7Lj7K5M+XCIj3xm887
yMAzAjBHyilytbCYbRgdvvzULljYADOcnv3XIzHeo076fHY3YPWSyywLL7yok3d2vjA2OdgrLNAa
SPrloMtCUHLL6cul9CcTsm5nw0LUhu9SAJiSjMippGELNXe6S2MoK/w0+PJbj0Z/Q38DRwi8M6Xz
VadsLBQnv/IDvnLZJFQ8/5+EbmNl1G1ZK5WxLWTp8U5JveSlLMsIz9/2hKKRzffOjWp/DuOwVuSv
OR0pC2Ok+9zzXxqMH5tOhnTUMFrFv8/WLSnCmKppNazW1MzmHc+XR6mk0UB2tKhLXE4HGzQO+6el
kSOEdPU26t7DEuiik2+UvGBCEzWDRpB2JEHYePNsTets8Qd8ZgnVNH+LRvS6NkC++wCH+VRlOcUQ
du6PIX3fc1UVuk+L0pw93FRqRlROYiH0ptQYX+Q6e+zMS2dT9YWLJlitqSv98R3a7FcK9rjo2s5r
zVFdpcrivFC22mTQlZ4EeKhNQtY+qhQ1YuoApwUoTLL+6gBj9O97IslqZdBYcGOSmY1sgI57fBMn
v3vb+OkXLFAiJXamZ2ohOxnCkvykGb0H8Qcr0udl0kPiWMYV7jtRqFkZRa0TFvTIOToSCvtiKo+J
KHK5E/THczcxridk7uvP4v/YvESpudcLmp1abdYm88IV5TpKr3tlbnZPgzObvb8pRI4FJWSTRsPi
M+NIl9OpfPx5fjcsAvy2AWz5rfzF4syZvu0rQIJRa+CRwh+sAW2D8a0VzE2aAuV9poZXr5T2Ps8l
UTIZ9VVCBYtQQ7HxzqNDIe/H/hTlW7YUeznWCIqg6impMre65TgCHbqFreUAQg3FFxAuksrcfY7t
6VSCzT7+iTjJr12Nb4LB98yowOLye9kGOezmX+2RTVV/a6rcC4Frssd5rCZRMu+XlXmrcqjATLPi
w29neHMWMHNbH+JxAnbPaX8HunbD7QWZnNgb1RxdYVn1DdAo7YWcy0kp8/neqgYmmGl79DAMR8Ou
R8BVUQJqPACsGRi0IK9xVNAedZRXSSqx9mlTIuj1Gq5J4M/ZwNI53cRWLOHK1qk7gGN1matvZWCf
s3nFCM0qZ9+aM2p4QsZkAKwk7Tig6Sjylx//HAC3mzhN7re+Wo0wF3rdZqbmui61pIRRlHSR/qn+
I7nP4fF26k+YHvZd8TYjebRGoyfKegEAHufmBSF6nhwk5c2LPzWaxKvK1bOpm6vfZKnYuSqkVZ1v
XHg+gLtDhqLoeBtvGjWUSOr9Y+cL0Ps+Gn4lvlrmfPVb80M3nRqkwGRi34rTp7gr4l5jqpI7Fjoy
lOkM97px5gBKtkErOkcdTK5xn7ng3lgHOMrDzRv6enMXmILzdCsg3CCeEULKuLsAekHnO/jE6/Hh
cNGyHrPf+F5PFgVjovuYz3KKjra1JWPjGVA0i9CTcPzn40ej4fsBjEwQkn8cOqbAWEPx0LryI4eK
rZbDqmaAQVt4uP33xMD9VgwyN/IBOOG1OzKwoywyiYYBacAPRRDo5aZmQUSY1qa3L3mdotixbsci
oa2cd+twKw5iaYbTePQzNQMGiXKZtYlz/S6nPOKmz1EpHGmYzm/jHs3KMY357mXiMtPEBtOBoFD2
o5jzx5q/lI9UHBJEBEAxL7vxsV2vVFR8eFQ5zwDVdHtJKG+Mkzugv99OwLq6AP13yPBC0JRs+LY5
QmnVi8457MY+Mp9gcLmQXt8WrIMKBrXYivy+yvDapE2dJc+xmZ/vE263vuKQR9cTULbBLm3LCHWC
VYrvoMJvPrEuixmDUa4cO8Uu6Z4xt9i20vxc14Yw/hSNo9SrcwhXgovDjU7A4yUue6d11uwaOIoX
klT/FVbKeSd9KUMpGetp9YfJ5yi9x2zJ74SdAXGpI+Y47OXyQuQV96Z/CtMi4PniSLqv5bp7mUjs
EU6BODQz0RLSoNHFVU9QUxkNPMdB9PQn2cxjzMgsi+2ZJLv9VguNQVb7L1LLl/jK1l6v2kQDn1/5
TfkQuj6s9B4OgvG5uaxsGqCucWxG3TKLX5wNq8o3Q8BDcBrDxkkDV0MVKy7Cr6wb+rZa+IzlFRgH
dk6OaSmuaAeb9FoyYezCBO+ytqxTPzgdW+sldVm5mu16fb/jm+LeScSkdZal5aIk3qHnU6QjeAAB
NmEP316wFVuCYP/Q+JOXDLdSrpjadYqv9RPBiwfXdfeGqRZ0cENxCyI15vZ9nEpNl8IOlQ+k12LI
YUWERTddKkTeu5DrCBqBaynGXzp1L0gU7H5ioLQokK3E4qk9eV5wRF5SnJSBBaqPQ0hcFRCGOVzJ
DP9vsmWijsA3KHSG7Yp2WPiShHErZ4F3QMQQYb/gApF+j6V1/CvIUeud7uXWRFfjO0QhkvQIN+in
/iBv9oAD0400iLKXvsMr77JOSA5roYfESovYZQlULNXQSOQEfejcsodFHDIb8xUUyQ7+gibN72DW
AgcfbqHtQ+1PIVP/oQ3DcWF/+jrlvyRiDMPOjuA9YAwZDlEgXX0FmGkKoPHSHDphzASHSX/r/pV+
xbqhIfIt8t79bF3Y/3dRwv5hZz8wIhU0tSvneHfuRaJLA3XZpPvZ6YiPzjtsi9Smbwh30TqQZ/8a
NJpaWi+mXytQ6d0PSYOqXuhmt+mMH2LK8hC0gYlVoHcRd9Oo98pJBoy8ks7byiuw6QAbO8ECUQ3u
Q3YSvg4gCh0yvLoYZm7x2vySOjNouKBM9/kt4oZgXm9mfYd1x9Pn9CDbhcCR/sov+VTKIKDCfqfL
bD/ruS0h9NfdFa4OnB94Mj/NJJ9y59qGnjdAfLIOqngWKct+7udQzL8EORzi42bZfMrqOLlpeULl
x9HNeHlfQCP13NVzPD8pEdhF+xsCpddpFq+cys8zvPSQM+O6ZfiuRA+l8yxMeCosKl7zlwIBvS98
uyvHq2XLjGlHyxQFGaUe+MgQOqZyjQ9k2Os18P0zOVHVPdJlah33u8PyvyvdIZ7gIRXEMA1rUJF9
JV3jMwOz+uvZvvwjoLtEg65aQ5dCVff07KHAXs/YxzpAFALZAJPqJ2g6LbY+0f7nge2HPEsALNoK
Z0MIAjNA5rd/kl0IbTlgAgGPL0gZU01bl4toSXl1rdOkE5BBh8GmYlAX39oYSphUveNrIFg1gB+W
CeUwqI3EOhKMRtNRykKPzzjaUn9SIWipsr2jDg8QBMWvB63IQGdcP89iPoekgwHQDm9kHJPT01NO
55xv0S8YRkxOXAqWgVnGQ0QH9vg4OISy70b+NkxATWvDWt5wjgo449NC+ZYhdWnPkHl+qQAlvRoV
uCvYzjNPDc6TfCfoarEhsf8Wsd72dnMuBtvQJf9p0vIDq2mw60JRq/iZFZaKCeThcT5RM+EEFcq+
l9DlsC8TagWsbKophA5kEwwDcHeAnk5cnQsrQ9t1AOlbCHVcoDE+9TwKYUKugcPQFViJZEPxeHWG
kvu43RB/qMwwelmBe864ASgtSqGlMrVI0h1VNWLsLpWP8jcjairsUXcrj/EN2FNKtHVP5e9or1Pa
E5a5/4FGToVjem1RGhWYo0ri0j7eeDxZ8Zk8BlArvUOR05B5Dq5p/tC8feq5OOTfBqzRdr1MkNrO
ms7Zu8ITGMFmyzY3aMyHUhFJtPMTfy7IvznegOxSHX0pdj/lVPh4TEnWXluNywqqjL3mZnbdfjYj
oX3l9XwBK4GULa1n1NMv7zyVgM65dPm9Fta/6QlVm1gHaO0nz9HpVPri1uCUVfgThFvp/WTuTnM5
R6Fp2CTDO+ruDetWDHAjim8HU8Rbor3rKyVIIlSSMndu0ERlhLltZewF3Xd5r7kUc9LtYY4NH/5t
tI4VEnHRQWgsVx2uzvXJUsOiYwbZVQs1ZoDboBui5d1xq3FxuwE1vTNRZQRSt2rgnMV01l08s4Y/
XImFO4IyY/XbD4tbBViLPOWS8Rb3O42aVGSvXhflG5L/Ierj+Y4WM9Cr48jnzddgMghav41V1y80
N1iEUgVvyWsAgqdg5uGlpXGpT+0hxY6sjp+96CiqpqDIOK+lHAIxOG/cLMiOXbGXhfq6O4FU6Puy
eOe54O34dHYPWCsHhrmBZoO9c3aEbZVG3YRXQEnw/nNYI4abXSzSlNmFB4rt24FbiZGp+dQc0o+M
ZpEWOP0T5a2qDAXbwqwe8IgDD4pdzJnk8pxZu1kzEit7O9gwMfssKPpWWSvszX8qkucMyRA4D/AK
uY8UU1gJlP6fxMDtmKgVKnlrZw6I3T7QKAOUZxabpS67VbKIWaY1rdKPqHViRBmiVFReelxzvYg2
27FJ9JJ/3dapmMeMwaqkFJK8SrL/k9ug6NRlq6jLtqlDArakRj2NP1jNz9j/Dlm4fpV5DUpq6+8w
Fcrj3uEWEznSQ0vGZmrqxZ/vFSdkaafoCYpf5qSy08j4P3vKXlP7rbqTWoa7o03wJSeNnJE0YTqA
PjfjQ0ctQw+6UFsgmh9v/dpMhQhhgXaDkpWLddEyJOubndYN9Lrzufte8UOiWpLwOGpvCxIcElIS
Ns43hS+4ASPDqgBn++Z+sEKWWH6d1CmmHESFu2ejkOXgRWITuRrHy2yrhIoHukSlTr9k/eLoJRNw
x7O+Ufqs9dORxBNQ4RwhD8a5TyxHNmxD0gdxR3xGcyBs2VCAPYDnHlVBe2o2VmFdR1c3YVPpmVyX
BumoZvB1XvK8hnCgbpeV0h9WgRtMP9jTFr9C5AJCBQCJjnOMXAXObrgjEQBTTj7UMf0HzroIqwdI
xYeKaGLVJrHCEsbKR+dDAtm99D6titYkssguScUId0Yb8DS9chB7wZ9QiO/bTEky0zR4WBpe/GlX
OCvO1NX2/3tUmb4QqfQ9hQrRj4nksfhPu65Y4RGk2G3Udit9pDbGDz9E9rZoTUhmIssZCJWwcETp
lAQPm1MjF2PlYW2b+4CKwqWafeV2OKerPnDy6OPk0MnRXNAMXqR+9V+z89AYjJj3LM7itmCcQxW7
3Lp8Y7fjXNcekEBnXpDB424NnLepKTU4nYX/+TclTUYmkBAhMzSBHUgF7c9haZfqptSvsmNlEh63
dt0FK0nRTcXMKynXeINmBdc4xn45xreXWqDW1za4t6igL+wUDbdaREFYVyLJORZXD0FLHAofBRO0
bAhp8Sl6kOZbehJ0afHbx7mVfQcSTcT8xaleeeKTnNL9dEb0eDtFyQfuJtIuy69UCpdUFpgsCD9E
bP5ki7XGdoYI3PSPgq3xE1dPAdvC5HfaapmXlHhJcKbD8kRWkXp2FIrXY5gcBf2vFXTov8kZzh59
g5/gBUZ0t1C9B+gkx51Opz2Qq0w06XlIvcRHRYK7qkr+AhSOsQ1BfMtF0nk4gyebC0qST+ezykTo
3AlZzwI/M+ljUgUd6HSlXMZ7+f7G7q9Dr6vUwmN6Lvhi5NAB4BfcaR5QHkpHPUo7ComvABJ4foGy
3k9OBlvCMdq43g+xXMixd29jjspK39Wvp/2uxYnHR3zfrqFWj3YhxFhfdDw1R+QtURSZ6L/xYuoz
zmjHDoCV9uVyQD1wIWUPzuSsZhfKDvFAk+5nSJlPVs1t2EoHv3ISIgR7O1Q0CyschdXG744uJAmM
Eb1LlJAyL+Kt5JaGuYOrvIjPRGmsc/axEbsJSGT19oeoP27yGuiD0QBhsQ41iU5MPAW9qcQtIf2Z
z+3rS4cJGYyR/baU/oOLnoMNpi016EoZ4XCHmM2drXaCpf85oB+dPI7ny4cMeM+oY7TmEvtOZgyK
7UV5H2zHWM1vBboER5nVCzJC3Bqj7+Wws2EQPLk2ySjgksrvM/b8L+XpkOd8lErBkuCcAKBZ6Hr2
yUzffLTnRYS7EwSxAh5vcaX4dKnkD1MsRQAUd8M8Pt/3a7PkAF1z7D7zCWn/RGttO2BZYEO4SEng
JwVQdtEOK2HIXNvUQBzwF+AD62yN5g6GNgtE0r1xyF+ZlaT/gNd4VsacBitv0513NTTECNOHXbB2
EwsGc888uv+tlfUTYgAwI1HKDWTjJnJ1DO0sl+QFOGY7SsSJmEQ0ZPtlVantJMIpIYgfTc9ECxsN
R8dY6EsP80MFcq8K1vYRwpASDJsrqL3VKkbcOEDQJ7NXVCFll6MfKit5nwQkr9qLI25EAz3Z61RX
mQ/RBBS/X87j5VymJMbRPgyV1wJKUQW66RZUTM0o8Fb2uJLJcnyWHDz9JOaiLPPKhJTuHY+KOg9w
5VHpda3sThVcoxVL605m3NI9bClJPrM4oPF+YFSScozdQEg4fQrXylGswkUThufPLf7KKPRyt7zI
y/QFjJWbxYYMLtdaMNhaCCRjlLFFWydFQnRfq9ph/eUabMjLb4wCkkdrnTp4ZxVYNPvG07cswY11
WiKrHKrT42kZq4y7T474ijuhqada3aX8wGeGiFuFq94LcKlrUMsx7Ob4imGlba3uJvYPdV/Yk0VP
/T40afoE1upY0wEF71E/OMfOq5C/xizrm2d2v4u7edB7de8szk7PzLittQ2x04LWp+ofkNYj85CM
AwoEg3NVn4GO7Q/xBgMzlNma7jyjGZ3b2CfFXpZuvI1NyVUeUiEQ7a9YD1Zz8A7Mmq2t6BDqlOCX
31Pl6xtoFM5OAJrQ1+69eIAkV7OW3m2SYMfE/UxQ4v8rArufHIpKDspQn1FYGprnvMYIfW09hmvb
N6gJ5DXaKGigXTJm5ml5jiesk+ua/gl6ugmjcFcnp9+HYw6XcIRGF+QhGO4QMmDJtB6PJ/mbvsv1
ekn+tbZAK3VnvLYRpjAF+hKxvqlAR5838MTNimD1tN9fIBG91AIBVxaPHKZjCmSuATfXOe2x/QHJ
KQ83/+Uw/d4UM7Vw49He8EdtXCcGWazmEgM+bANJQ3Mv2KaNBhe9YtTs9hT2xCTfknNiaB/H27tD
/F+YMYBeQ6qh8EfAo+HEFzXc5Rf9PS5a8bn3w2hcUqLWXttwMzMF80Kq4Yf+RSp+CuNgVnXQSfui
VATUDlaSaKdwu/9LENh7rFBFfZVRM7h+/ZbYxm4rbGfAz5hY7Tww+Zuo1sQX1l0lZ5iKVJL4kR9l
YE2UCDtX4akvhsOa8mNRCJe4gqeyKBoI+wsJoQSVUU75Sv6InNf8DIC2gr+sCnS+qWGe6GvE4WyC
h0BkDdkfEybmF+AaK6oGLQPTpAqNPoBl6gjTEQjTSdHfqKk2Bg97gjBfsLH43SFVWhHupU7+Sy1/
3tbkNNaXg0gINTWL3PA+LaWuXzroRQLj4l1E7Gd0/rr4skrhZLZfjVtffU2uI0YLHFJoHYwdNF/3
RZWswab62qIGkDSxujlUmBgW3t9oU1z5DoOiZhSlClI6E/ag2d86WyYJTRH0Vy1U2aDr8uOrcLOn
WVwlJ+AdEj5nSN+SdDokayiDG/hNQ/BjsMuMFeNClSy1ukEKJ3QKVQz32PPuRFuH0SvZIJNB5w5e
zpN7aFJMtfsVNquNKMmEJMNdVo4oy5jWPj5RvoaWQcFXAs3dr3yVZlo1e2coj09tn5zZIWrW4pl9
JQqVJrTG1SZuUQpW8svKtbNBKWgJJquXUjC0ZOZgcFH5STCYslTViYIvtIngcfNRmRDIy7i6l6rn
DBXOop6JoL4uA0KF92003OtTTndSnZF028BId6GHdS3BezFWtpU78+PYv3Jj3hcm+mgYPD8tDSTX
TrL+woSERxeDtn658po4fpSwlo096l3B2kiq+vrTEBSJZLc9PnN0yVY6nx1n1VK2JwWbgrGSNZoI
Pey88FndtqSCgZVyeMZ5jEtGE4vFIU6MH80fjV2BQQpknK4D7p8ni87/tiQwcfLipj75zzPTBD+z
RD2LJI6oDK70d2pFfxdyDx3B2ibtjdjYQkOLArrjq/JYRGSrqLHUiyFKXXEXsDYf+Adc3vRCdDjG
/Uk13hnK31oaEykxOUZyTGxHNgeg46LtgEKLLA9CNAP/PIJu9NMPI3hx2WnxEMvnZh9twVijgQ52
xnvBX1Hdr0EEjBH+uXY2tQ0JJcE3yIZKdxS6A/bqamPrrTPH0xHxtzQSpNkayQDBT6ZaVRtAkC8s
IVZbb/Bpa8hVfIY6ngDz1Dz29ALb9zImy8FeS9vwm9KCZ4hh5nta6zYUYV92Y26FIh7mfEVqd0Eg
Z29XCZsrFhBA++iWk27vJ9DHMaQ+VYmuSI/RSVWZ8INyBlr539evB968KQZRKiI1puWKsiUtghRf
1IgXfKD0p1r0QKBSPntgJ22bUP0E5jbHrAGed28k6SdiS6FoSVXsdBKsE5fZg3fjjKuMEGkHNUMS
3g4MoXYG33LUsr0vt0j/HqQNnoaz5mP0BFcruqHBJykmqbpIBqEoKn3OMHWkIYNGslaqicXKZ4qy
HQT6HjXo8BwPi7xny61B3CtY251iZyZt8staB/qCYOCgH26W3tIOgFNIeeTRowwEe3yE+3pCYiYe
nkdQy5UNrVICB5SOgyP4iag2qdPKEHuwV8VFp9tw1I/psJB2XRapIW/KDP9rmED/FG2dBpEbL22C
ik0K0Fzvkpu2qF/2OCwuWmz9cMVH5r38qHA0JYbSA0wBR65ItK/2LjmRRbuAtGc38qTg78b14QlX
1KrQMlB7pK9hQi3Rk7jntTHv7avY8nBOVqc0oXv+X0+a/+m+yoih+fdqZYSz/sAygm2aZeMlnDGg
9Wbjowka2Qez50aK7my4qfb2NUW3vm87Xgx+PyaijCaQULlazvf3OpEhbmCENc06zdIlNBrZUNjq
wdqUj7mO6slFZMsCGaFOoBOHBDgawHZUUfVkAErR2hzr3U80SZ+i0v3k3DjYpAOPZY0urlML1sC2
k/d6po0E+KXP/8fPxloG+57IlxlbNi50eTuYzOEb66imkk01pPXcmHuf5Uddse6RGC87ft0BdfPC
9OyK33hR1UazPM1ykh5hiZiC2D0rGMm72FJLYN6Bp4x6zBvPjKy8Y8TiKZC+f6Oz8POg8zgHEOxa
0MhiyX4iJhfpZouCdWPTk07V0A85tNXuUrYGQOm6KwShSTZDMj6RWCvbfmrZC2YfiVSAoCc1u3Kt
+jNh8ZKZ8t2FPmzkVEaOPtqoJswO9jo0sa/+OVTyjTv/ST8ww2J/CiFO5gLQI4mB+VuKNdr0k99I
/WyeohdzYzWO7NiDEaR4jViXw80U4kXucprn8VVjLPIqjvQtc/CH29sZUuTDEea/3joqqSw+Hw/O
P/F7FTD8zIZ2xa3sqlW0O0zIJq3FtU8m/5M3K/EJ1NZtOm7Ycj1PuleeUHEj7apopCW8/uPqc3en
eEagp9fxoD6TE+cimJEf/yJrBjuUhMHCfst7dbfsH3/h6fwJ2fRr/gfr4+911QQJaJHdBF441+wd
ID6hxd/MZ2VKQjeKdcmhY1evOuPNfMI7S9XlA/aDk/TzTr9e9IFJ+hUW2qUWS7n+wdpTHm8y7Zgq
u5S5X+Qo+nrU1XvnaHD7zg40YPe8+d/vav49id7s0OIEXUYzqaSe/EIs9h3tk7w8AEwENr42vlOt
70egLgyMccPFCnpk8Fkj6Pov/WXr6+O9iCmlYUEoSuW6pIiZmqjbhXTM3aq6RSjYQXUUqcYyViNN
/po+dyrG0e/DF2IW9Nk05kQZGQcHiMaNJ4W6yQ4iBdJeDDlEqCNReMI3c5JS1XNa72DkVYcDc2xV
CSPQv+EvdSqEiKe830ZqWHngLtBrDJgXGCMOJrLpcQ5z+z5ILdptHkVv7swYv5ZGMPsM5iLt2+4r
1T4wB64ZFuVbwS5Kt/Iu6y7SphfCugIIx3ym4iFeXBr5RrxopW9CUcjKmxhl7t3JvlwVCnrpn3ID
sA57rW5B3MCbHfKrNhzFe3YrA0lweIv7uyIA0RgN+LMXc6asZrtpFedm+rrqI050fu7YPKTXhET6
NSPVmWltwrSkvDKVK+ZWbarDjBSu5hcEUFcig2Yn55TXsZpejcwadQTp6jqsrvkpveannM6f3RZ1
c3McEjZH+0MsM6gG1h8TA+0+DYMJugt4b6HAJT1pYHzsePJOIDtVu/X2mK5jjbQYSNA/c52o3hti
3pe1zvxmZbF7aUJKdms2zY6T8JSli/4KfHVRNsQ9bYefrxFvBA+HwiT7WgKe/NyuGKGDjMp273b5
ZdTxqp54Cq8cRdu7rMxlH34yp5xqf5D6zqCn9rWzLjPuNx0eP2dVnsc2nDVz7BgZXtEjEt80Gpvg
RCR8KPKNZ2YbQJOhF8yeWwnbxnrLZwJDntKCjH3nlEE+o7KNHpdPp/KdRTOrF+vjLEePF85F1TP7
t+TiO0Y4oByL1RoZuOimOZoOMCO8i/PI2yZgp+FG0M53PPQ5mBQxHd5aqtuimI3xDcdRC5zsEJ9s
aB8pyfHfb3m+FTf/5/YuiOv/8EkbLq2DfTz5L2DGdH7l9w50F0dcTZAFCtJ/jIHd0w5Aw2/VgQax
P99uqgdVBs55CbXglZDNHo6XN0YXYC6EnMAO4HIMNfM4T08XxGV6k8p4zzuGTlLlXf5cZnMDuAJL
a9ktjDzg9Dw9OFI0UmK5dyWvENsaQxkQMwrM/mTIT6NTYg+pw6brnNyWhJNYNjxKC8KpuXmusulH
Reca1XxJB4gN2ZCWNUohL30/X9KnJPbJC09sSIZF/GCpkRd2L4msbYHTJdjKh3k4cFyooAJatqh1
yn2SzJIOiy76+lMVEEXuHhY7YJR+LdwU5oXp7Y+O8/YtnGbQG83VHMeOGj7WCCgl4rPvHaQtzLf0
ClJr9+nv6oS0L4ltK3ZbuQOlvqnF0cN4iCbIpdlJhnUEf2SZdUruC9tsiSLVtNEwfr+PCOof2otJ
irLAhXbN6EYwXpcjNzBthgIfM3hqknFLWKvRcCYLCYDd7+bhfdG54jNIKBPZ+xyEWb745Yb8xuAb
phdlSpWWagEv0CLcFdDEklnO/lKikYx6crICA4RI2rCO27+nyHLN+92JWC/j1kJOt3+EZrSNhm6K
pv4DlM7pF7mKupfiFrjgAwq/v03zhwd6AbEnlDuV3QtUjLW2kjFQwwNXLwY4r/WKOO/o+f2SNCaD
rCiCChTuhfSPPd4FQRul/UEQ0hjVQ8paAMhKviO7DZUsFERPR7U4NH6iyS+2rB/U/5uQQ3bx6suA
GAP3hF5zu9gLuSdCBHxTQ/nDHzMkrd5cJHl3v4dAdkw+kKFX46mkUcMjzDqUkA7q6icCY+8a1ypM
/s0PmxcTDVWnwFzAdJM46rYXuAdJRtolTXCoZ751FQ6QLm5GjfqB5F6nvQo32jtEEzv6R8oJtQ0R
awUQPlM3dMok7C78n6SWkz0sPNN1qxYBLvlN4ETYefdgaUxqBYGsR+OValNokUj4On/gDav5hZNP
LA265s+L2/HSIe9i9VaSis87HEwKt2B56dIMY60VJE8ADBcFYhDMUwwsUin22wlxsRp12RPpuc4O
QfnuMgdOr1V9adspOH4OaX9i8y3TrCWJNTQPI+hhGWrwD6HXCrfk9UUgyUyBLXwzkM35pSTDli7H
e4D+Aa9b6Ckc1ZjpVFmJCBf1IapssKeXB78+XeafNacx8ssunUgMMDET+8o+RCAsDBlH7kPbcnPr
isbnR24J/X+sX6denMTwOxUhhZa+6i/sMwPls9LrrKzmrICTyT9G+3pnl1cSc6k7qem75Ks5vcZD
qb2Lre54PK9wG5liciCN488nMuP5czEAjOg3ASv6oOcPY/YOA/ufpnrzERuWS9YdEa1ubx8/yEUb
8gDZ1BRRQ6lOxBhjvyI0xLTpb7z6/TXSLc6K16S2yITmsZWZX6YbULumbnhh6zJEwBpj3QQsXWKj
Dm4U83rSHtXN5caIc/izxpu36SYD1/W/t19cGNCDYw1O4L7Od3g2Ku1+77OrSPXVj6I6IahJzZ1n
3bCnEYKKNVLT1Rkie5Wx8M+56b64F3vNNDDS1L6AuDI5yHMmSRC2zLsjc1w2nrJRcLeaNVJZbyf8
HwKhhIIQMGKjpz9xqLr8/NaW6qsBNnImjJfQnf7WUwmUFg1diIpHFyfSPfvdVjaF4HO8rMzR8BXL
U4zHTwRU2iupo9GBJdpueDao12RygVFwNhdkAzTefeGU7lI2dgV6T5VNDy8vnrTR/QAe89RFiQ7L
7YWv2f4wa+ja/wV96nldduRbPrylW2QbuDadyGBWNxaAXD/Mw0gpLy3slDkE2dbdo9JUdbNzw/71
oQHzcmpNDTAlhWKJcIitI/13hB775CMoZ8quIslItzXeQ8paUN6b6NlkCTrkvgdVMYKEENH1nMUP
cCy/O3KFEBL3A1oxzuIq8e+FmbiFiQyh3vqcc6cll6MBhf1AkhGR/zT7z2KL4dmLXjSjhopLEIJe
ohCC3bFyIH0NeIFCYg0UjvgvEmkG1HndbUdBiXOa0G6eJxmW2DwoI19fPH7ptK4G7g2nvIVMbFm+
K0cUOwcy7+SS6kR2IDidzIDRAVl/aBRkZoTzM6YabeMXexnhHa6iE+0SX3X/Q8800Aj435SVVK5N
UWB0YurQSGA/y8YVVajx+Q3AOcFrNN36gOJeopfLy0sPJsuT0sh//wODbUOw2ZG+DoyKu4B/2iIU
zlDAuuO/zUvQLJRi9WWRS8EIIw2p/dSDUdG8c/k9j11m90k7Q73k8j5x4CrluTWA1C4zFsRejo4c
aoX0pnMzQJEPYDZUo0TrfxlO1w9N7D0aZz3WjZO31ALeZbJ1oO/lY7qGo3l0uSBUXq8LXS2T1PoF
Kb/deMuX9CaYm3K9eZ6qfwEthHoYQ0JaxyaqHQVy0m1sO8kxF7f1HtsOvCqhRA8ck1YPMissB6tO
7wC9NM8UXX5IbAprr3zLaOv9epfITwBQh4q/W7BpSybgywct0AWlGzbx/3KVMpjdc9PaYOPneY56
/lyPmh/PgBVp4VHBGuWucizOxx4uy7qZEHarW/oYcn9SYBkYzgRiKmXgLfK626wbnCKza7hNSN6D
7ST5hooA/boGDZhLfXknkYcBPPKVZIiXJdJ4ZuilaNsdB//dIHoR5TZVM3xYxnm+YnjUuMvBpNO6
1bObW+0c8EyKsmBNErcB/GJk1PQHS92B0f8gor1lzVr9TvBSXqsZW/Fm7arjvQ6yMkj2I1bt4awT
pSHLg0uRNYR3fYrQWwdiXyC8jCdWadnJYA439qQ2xfpCCfQjKx1V8CkDdC+kanTO3ME2aM0xrflF
h5Keb3jobvQhja5w5s6JxhhbfVbwtVE6IkVQCD801S73eoSzniWp+ecSsqdUwxncSSD7G56hCnhW
MI7KMnZd0kmRUJYKrBqIaTxG0OJnor7hu//Ti14U3p0yiPW9frqFhpV0xHwKXjNlFmd1MnC9Fu9i
p4iJ9uUNENw0frA+jVwEXS5G7Tg6BAmA3N2ssj02Hp3MliFFjsjQ3mqTZRwj9l5fv80y9S/p/70j
+ulr5cot4AIXEvP5BjmIob3ToXXBXD3UwtIHTpOtrZf70vKi5ifeBAcN+ST3Nau0cg5PSCg9mixA
EhjWZ7O0doqrgx5weMRWJ38GxwrihdIxFKgq2P5G/q3f+Xuz9cZSQ0qbOXEfNr4koFNbRVR3HKrY
cf8bnLoQd9RHHNd9PBFu1BTVWS+r50QMKgpKgHx3NnvcJMmZtRZxGDdfcgRl5c7qOAf98HXSHOlQ
YGsl+NuXgkQYCurFx1Fs0xzPzPaMI0EjMApSl3hN5kvnDPdwAwfcyPsze31lftRGcIJ8tl88X6pR
HStb23LwmY2yy3VqrB7zyAikz9hhTM59IInFPucaxcK9Dkeq54iJFPl59/hByNbetBVFnGxVN8Nm
ME8pl+NgEvPYOsU/T2s6BnGUlZohFOIqKpwhDfFHXvkFHvT/D3Xk/+nIhbErLJ+N5LOXlmYb57Dy
q942uKED1T+m8Zy8NpKoPiUFg0O1rNj2rF0yuYh6tH3nuVntlRmh5DV8Rbte7AakIgLcjhysajes
oK+bVp+ZpN+/llOGlbY4LkVe4MA0DN7+MraPrC63WfKY8SEui6mdXZCYTgfAsk0151tSl5kU5RK7
pIzJcUiGBLfldtTU06ybnJkcLk1eHSbAel03GJnZxjpqPRLbzr6QON6HzxiVyvyvEH8ZNGtJDeIN
rbuwSZsXhibxGqK4/jKAsvG4OSzM1KqCXLMXZN+ZIbRjnhfeAv3r0ZSXZ6yXzMFPsWN8xblrN9hb
nzWkuV2cqU6pZ8NzOqpdKRKEy1orNPQBwpSM0tslH/gncULFgMdcmajnL+Vewd0/xFA+DPpoR8SL
GMcsNy5WXiQoseABsiyKu1dbmIoVg8oSlEgiSh34yNGO8/PcNKbv/kX5QJS6Hk78iz7s0133+wax
QAzVopJR8SD2va8IJBs7ebEmwObP9OrzWfjWXnYpTHcVrPFbXyxJwLgJ7LoKYnZ+pklEFrJncLQC
cQel5FCEt1DNBXGtNz7y9nmuCUmYRaUEpuCTcwYPbyQgjrMrUWSPqfxDMNObJJkPzxdPBC97zcOE
8bG2IjrUcGAS8UinpJa8La2S6umZgs+20D7PnDoMOmV0laxtOjmxUvw+4q8XB4kq9vsoFSL8UNZQ
klemKpigULTvzhIVyFfspuoQfc/bcW14zKGu0W6zC6JfL+enUPPasO8wn5nyiJhZXT5moeVXa9FC
jmsZ5PiASzmpmcVuY4PjEImd/b2d3nicmD6MmnVmvLKFlSsXBLFoP1qR7BY6z44WWuEfAl7YRpP7
YNoriA+RX6XUTaW9J4+YKCv7vI2mPUdkanzFrpA42YMVdYLrHSGv7vtjLIYyILHmuCdlCFtVXdCz
kRb5NIXMg6ywc3Jm8GhMORFuMbJcml0e3DAiKOg71t5+ukMgfegCJ2fl/3BP2ObKvxPYOzdgzOvx
UrO6NA0PuLQNTDAmR4A+1gHGoXdrj+t9Nv7czQKT9vCnRtOKE7r9RzWWMDldGOe2wgO7IixyoY1T
x29t2ZfqiYuZ8quXl99o8++W37x/bEWA9f71bqDS0W1QSxUzpirXNqGp9xbYaA5dt3AbK01A8x6w
u6fTfxOdeZ2qvlShA8xkyBZ5baCFDc57d7LA4esSr//rmhTBrRfuA9qnjQt437LX4PSDBm6+zwkx
T4YoYQHLPv0RBAiUg1jateYfaFRSI3I6F/F+DozybOwnhU83QOb2KVzDR8Kdg6Bki9NcajdyoWIr
BLm7sEfTkSM/AjOeZZ1gieoF7OgO48Vrg1V578CGBoeZyXJlbQtAHJ4QEHhqZohdqhyfYhrEHAq8
pF/Geis2unuIoNe1dcqADhtA8xub8cKqfKYi+wqzKeMK45vAy/9kO1M5crqdYzLtZPWBRX8BA9uT
/9wJcmGP1a5e4qzKf8G+WI8Cl2OAaNCJIdezt0R4cpVBHErRty2XD4EpIiArjcESFCOKEPDreZ3l
/Zy5tnS0EXsPiUgoZaZ+VDhEf6Psk9Rc7ch75xzO2vEht9CWGNkYpueKFTmJA42BbX+q6QZigYIg
V3yFPaN6Vv+lWFulrguv0rJ0RIJoZ/nRITnp63MMl6WXHT4il3mPZVAeWdUMYZd+oB+IlfaUSYRy
1tzELRdb1CmuDGA2hmE+uXLuDaHMciF1qbLKvGuaQsLrsqjXOM76Xu3sGRAeXFbIZVZlKvcV8HCZ
/kZsLpnyRYdrW2cowMqIs7dCfNlyWK/odPy+uBWLk43qCV+Xq+4U+9XXd1TfWHX1bSoACm7yciy4
i5+mWM8QOXZUnXo9+7Jdl+TD/6I682MN7aew3Py9eIvUUTyjTnKBppQbXg/efFpERgakGkeh/xBA
IHkBi9tIvh7QafmuFc9kmlDMG8q+fpLYXaoymEHn/V/u1ny4TEmv/G1R1+JaG+iJnaaNUZbbdyT0
v5gPKCRx8QxgC4nj8FqfvlbaztNXQaqJSjMNGZz4aUlGT481WWd5KsOk+KJyPYK7lPjqu80kAXD2
/ZVntgw2Ylww7awhu15/338tUFKJ/ynK27bMGRrZ2nJxUoIDMIyvxlPzyMLR8FgQwcrikqJqUPru
hjtVCVtsCL6sfY4uVao9QmnMRlwl3DPibvJks24JxKrSIMH4sdx0X54IUkE4debRmFSY57eDoX2a
CfnAJgtFli6uH8t3q6FjdipmoG8Qg4RXBrR2ZZ/RwvVfi/3piyiI8rRw9F7kx3AxWsnhASBolvIZ
nLNXleYrjW4OrLSeEmCeWFDxCu8IJhuC1OkZoTjNhWvjheK9n+PhbJIN7P32rWSbtlankNlEERsq
Qlb3dXfl4vtu7w8B2WWX+pRe1YbIDtCxuRw84pjqQWSV/dooSstqKFeFqG8glE4HGcNKR+BIoEf2
WPVIqe2ARMa0Cb0pQva5FIE7pfYgNFMrgmBVx09igUqTHJFL2zpC5SfijKt1pn67ulg+FvS93qN2
JUB7p/GVXZCnITmS6/3LmRJs8Tqd098l8ilVvzN5yXizje17NLZKIcQAx4hz5NZDbQlbNYklciZC
oSLHs92PCYAtM3Owh6QFmFByX/w3pCWRg9OaNlj7evtiTyOPh0KBst3i7ea5vXOo1vwc4/aTxrF1
Yo6uZ6FSbP/JC6c0gKRMJv0Fv31soZgmR9k1T/SoL3nVM11Xgh8F6qSbwZUUDBN5M95nld5kVWKN
fiesI6fYBE7/zNztB6YkJ5NUAqHsq6hG1UzjUHNdAr+9xVaR2ysMte0Iceum7pvYx79whRssJj+e
XYXpk2b/0QqGL02IKdP2vhxSHsNl+Ch9/ViIfEWtjFYWd33KcmHkCSAJqVF7nE6wYlLhPzbE/cQ0
5TdAuQCohEiFrxutLji08cMqkG7jQBmd1K+S4pkI6O3xYI8yrz6b8Wz+g0E6XNmzWpgAgcifhuTg
4UoBy2BUjBCe7xDoqHGu9bjZ/oalqnbZjFinGnMfAC5Mn5IOy7xtpewjktWaCLrL6dRxCOBvBYvL
kslKj3BqIwgUAUY8cMLJa68lbLdr2orS37oWczavDX02jafeUnU76HVAq8EPMOKuVTWlGgaQatTN
+h1VzkJaBkiONmwx50Rw4Nnxq6fxSHjim5F+odwLlCgpwswNsR6R55oJCN5UZkzj+2mBxQZGS98+
ZXPw+MyCJqjaZX9iqzWFhUKl4/AZLtKCSsBfsyoWokP0mhj9svdUVrmZUDgfvewIWos9eC3dEEYO
jxNBC1XR5VsdJDQoCMmGk4g4U2XVnRDqmUdPq1R8PmiuZQXhmRYWsf8Z2+Kg383ReQWoTTd0F9xi
Om6jZrV+tqOgddJMoCamAz+Y3i/4N4/g489ZVi64Xj6qirr8fRslOO5OpRrKMU9wakhmaw56vDG1
qgSoifPwoLxXqDXpWJtftVv3RV2Cq+LT8lZ/RtTc7lYTSYqysILrtIBLzpvG+rI4PHH8Qs8noJCo
v+2hvUlEzeEdBA7Yng0rZdPGjrCs7xKOosVY0ap+tcIX9gQNlI1ADamY3IrM8t3QuIt7XCjUHNma
1kKM97eOw0VHdbyzcu7Y4DpYTQ4dQHxwM0jbn+cCSyb3FIHQMwXiQdBJAY5WhDGMR6nVXPtj5Nbd
ykdKUISXUy5dJUqEN01aKEH5j5NR4lKpAuuuOzX+6GWz7gHuPm0vyNoipE+T0UHJt1gowE55dk98
VEpDE6z8xNKruq+NnGiEzaFul/6HTu2BX8qVrEuTN8EzzZVpg+Rplsb4LVZPfSrpu7Tx6dqyN7pl
X+uxpJ0AF9cSy4CAg0ZG0JRmrV43RTVSuGEdEKGAeTkZb46eep6U3fsNKfWTuD1GegCK0WnG1LpT
80oC7lFXYGnqu0DF9nrXVW34/HeqcVHd4WoNgaHwO67LAitVbwXfOFNqzk93OPCBjiEZy3oCFGo+
mIJ+IU9XvIiypuzjsEIGboQSmDk+TKoJJMubYaoHmSSC/yAREN7kZ2DVBg149L1ShzIIhuC/kDZ0
gQsfwELbkxPRbQdR2hj29TW36odpLXepW7A6xUAoIbWcVD/eEKl0+uG100zUYZr2s/u9GerPvyz4
rCGrLnhTBeZ3TKQEbwQEtfVYcZG3vTR9Il06ZHdhyJjd6CKiAhffbWQ6TF2gfDEMVU3UjJ7i5NC9
tjWYixPSr6frLcPeGK7R6x/JaWFgetohJgV1ClJy1PirUZI8O+zU/KgJVpT36osgz5MEa3eboabQ
XAozqxGNu1kmdEHhZDngD/NEiQfvCmYsXCLLRDAdopuepyzgE5Am5KKqV5Ouu0n4/RXgQYOk5dlZ
at11m+wK5fyvbTiB33n7A/olN+MJmKg+6DwAO6d9k7mo6v/QGMrM+NakzQJ20JKcq8TbFoh8grYz
PjcO84l0J0kYrGBOkbm8qcUvSTN2MygxoWU2gifRuqnFtu6n2Cd06YKemkIzf+eHzU260H1H747K
E7gZQvWoFq9AVxsKgNpWPc7qQEIO4cIpPcj3/qn0NLI5TUM6BQhGzABvNo+grWB2cBejiB5CdIZj
BmlOJ4h/zn1Y+SJk294f07CXOUP5PhQy4VnrWwF9DBxoIHzw1TM/rQC6G7hj4TyR0IPVCeXDDL04
1PaAQ60ot3d/WBbdjr1RBL5PDuWThcXYhWe7nhYzFXw2tSH/jCreZVaNt5fTfvwu3jGnOCEHYFb6
7Qm131yQfQfb8AexxoQqsGrZOBOgOuJAPwkp55m1/rGy4gt7YFRg5/p1hln9vZ1r5ROQBilsYvib
kUA3qrCFLngaCIkg2bBRs5GkzmOvrsaLtZ0EF/0zFYrbqOryAd3BtcsuGEW68+5/CeTeNISixfrr
kV2+D5lTPligZKNMW5/alBYOorpqSSXX2DtksQXxiT/fYl82X/HSxbQFGcvab+Zc3D+jXqNDqsjw
5AHoQqDQi6R5sfT/QhWl137bMiYeql1cNmKkuC9TkjZgzWytturVOv0d/BxypGc0BMcf/1hUvcNa
mS9xA4hKXeobOlZWoD7E47qjeW+SmIcygfBt42yDmKjaf5fIJ20ixPOtv0Crq4p2pDRusQpbJdCA
oqkNOw8OwmPDRz+ThAm8xEpsgpU98FtqmnKTb4sp0rvObKBmlhXblqUR5MXFFAPOqFb7kQVCMpP7
9IivEYfwfzKeuxIjOq25w6SHc1oytUSatl7Wine063/WxV0zWL9MvV9D5Ls8juxGOOLj35tOWvlg
24T99yl7tjGFeQZJGIylmz8L30WgBxSnOouClpHDszFGTzZzM0mX0CZGjGq694tV+UzEDPj1c4Wd
NdRsUrd22iNRToAKElIpIi/cPocY+l8YMH4NK72KaqFmMBVlJZb+v7YNnak7A+Q6Opop1UJeetfe
iFjNnrcZAns2GIa9KLMX/jF/Tl17pfniodtH8kgpn34z10z7LTo4ay9fQYU51MkTg3Qx2bL6+dqI
aBNebjLHSor0mCdvQ6PxN2F9fSW3O0fpf8GaB5Hd3nrGBNJD8bIpFaPO2RTx1pedvA+gmJWrGI2t
6SaAkyvgMb2f21KRbMS4xF8mOTece/19AX4Q6Zk17axfjp8vT8BrZNxc2cOl3GW5CbKGL0xRWeXN
00RgzJg3rfEgcs3GPXFY0mcxTbYi2hDi0ZNh0xV2ne/UkWeyv7MxPSVXA1yAHcgabxvcYCxPzBiw
thnpxJLPfXxc99sFqiTsenbfH+l8VWAnMBTOyzdgTSa175T+a4wVWcvf7AzM0EqLaFK+FTZv7TD3
FTyrG/bTP6xHEc0+RKw0cRiFaCwpHKmqahOfM4ZCcJ8SaFRGW3aRa6m0WbaMk3N8joc+blBJ78Bf
TenAtzAwEHQBWzhq/cyooZ/UU4IvcYZeG9WVfdPhJrx89CGWu5ZCBbjkjd+hEhrnLjkPgZiHoZ8p
Ciiig52xwCmDWb8ICaZyOYiHzejZNkjIBuzUqvvSJv/sG4Haho9ksUMMTho/UZQyqGfQ2ppbZDZJ
uIUMmSoaJvukIbvtgDMmMzcgH6IysjuFJjUivh3quL9AFnhjUU3QD8RZrrBfVO2XWz+IMrv72zxk
/vtatIIK4PGnvIQ4trPGnhlYXS8WtKwXbjjFIoX/CwetPE/nHfT+xiVgj9Ys07THo+uAZA6tUriN
70qRrAr0le8qZB4R/tkaQUdPnThK1D3iPt4lcccM9BUk+eYx2NmtxYMIEuZIaPXPQ485wFB3iLvy
of5GpkkW+53ejCfYyhSfbXNVwWC7CDBCiiA7gXmenwik8jCY6FZ56UDLAh8vAfrjFxZUfl6okgVA
tFElocw/9IKZAZ6oE+R3MJfRIAUgyZLUn+KJccALDhPyx3cJ+3LSPpIdf2nSzMdKSEk6GXKL7T1x
i6DmxmimiDcOM75qSaw5g6kTFjzUiIETgS26jG91dyRg2cFZe2igfJceKWElkFQSpSfgOAvduu7t
KkXE79QugDGJNeje38WNMy/qUSIsvl+a5uE50BAsz/3z382seL2r3t8fSGEhh1Wzp6F/P4uGj+rI
Yri+saBhnUSGwlO6P+q+CM3pf2GChoSrsOE+ng6PUO8irs8zfsNOQaTSq4SahCO5AOiaYUHeBLdu
azlh1xeDldNKOeB5KUlja1zOQdJQvw4wbDHJi7jOF/hLCE5jG7eaz4iM6skl5F4/sj1PBmf7WeMM
OaAA+TJWPHk9uDYlPxM3xpIuahAoSDOi4ytQ/kC+4yaSRca+cmmblYexwOu2JSC36/+I0o8iaXv3
Z5HqBqUA2NfZ2pEHsoWSFbHWTNnozVXyfkBFgUYijgaKbX929aLP2m4WbbIjmGKOFFl5lB1tQkv0
HRZOwS2zYfu9EKW3gymg2YeUCryHBG5MZZJbTXYwcQoZb9szWObuIUIT/cmdOW14xhMFtcIzkkem
7/F0W56PNq+EEPuJHXZjtD4dQjYIZDvKhIUf9wkQnrRkSS8/uqQL/emT0LUL38/qlOk8DIqw22Ap
IYgwxC0T4jMCAyN3gdUoYgqSfal+Oi4OiwbAbhvl9EwT+yNITpPNcgNrB2WV7KpghE5TxHxPlNgO
nPq9PSjBlOExjEOFK/GrdLmCdDRsPz/LbSGGdpKzC8g72Kzn9iO6nPMHMlW27QzEN1GAhBekgvS6
naTT10ILfspPdtV97YlF68qa4dVZxFxVrf0sUvM4Gf3qP97lTplgnTvM1iQkqf66UtTIA+3CIojl
DdW2/zkvkEqrNMJtCGh5wS2sqmMZOKNxxf+GdlNmv1cAqEEGpJSLzmVxvCr8WZg1Weyhtlw6ST3/
XgH8ocBrQr+kXQjGQoLlEFxh8faY98HLBPLHTCyW2Wh0VKgE8YZ1YW5Z7f/RLadrJ9ItlNU7iKDw
61+kaiX4b1hJVeOepfS0HI1KULITZ6O7X3PzgZcTwDTE+wpYuq5Fk4iJnp6mQTbfEoGnzSW5THE0
tipHoLIfaFhKLD0f4hDDHcUicRvm47LaUIsrf7zDu6bLVKvW2ClA8BCGj+P2LRONsA78vrNrssc/
rV9N8svV8ZP7x+yvBxhj5Sv7Tw83Knql6Jw6B7IWwYYQPFmt1WJImL7j4wISPWNRB6uHm2MzZEeh
ASYi1gM09qj1W1UripDkF3s/ZU4tQNpLrJqdY2B3q3LyFkMv514Nd+EgiWJT+yPF+Lw84Xxqo5aF
/LbHjWAl83jWQX2TckhLwkcLNrNTzcYtwMdM9j5P23Spd2jleoVTrchMmeYkYSfrz61RRbwmLQb7
mpppJf/1egMblb9iFOC82lcm/RUBhGnVEd1mL3bzbkdi1Ct13Jx9O5aLcWBVJunRNWoxNHHZzmLM
hvhnCcPzlbbZiwtLecbBlwhF01isGZy4NL/c7U5SJjOUuvK6oF7CaVE75PwDbko+FS2acezBCjhF
W6csrXz68tkSkvIQYHAjgvXewEoDXIwG0PbNcHV37E0GBsXCUKY9kknFqjsHEquxZwuqzNI+o1XC
aEzl1NTuSZXTYGs1STeJzW6zwq0WDujzmf+rXWrOF8PvGnuf7i4MrT6KWv0YmUV1/Y92Cq9FgLgo
zhZHdoeSa49uxip7Obw5XgrNA8/I47oI0W7lOLF5Q3tfkYTelbMbhSuDe5jklRU6ysMiFWGIdxUu
ynxAecDILACwLdZzYBcNBXpeaK8lnvjGtrTZSh4VA06jTCo178vXBrLQe39duo83qIcQEFq7xV9W
gjjsH2l5NxdsP8AY91AJwSEHy6QIbieR4VIPfmUXsiPxu74AVcZIWqVQI7aX1f3lvuI5z1S1A7WF
gXF3yOEbAw26mT7Dmfaw35V+2DXgVDKcWVId/5W6p8d4q7WO+Oelvtl0e7cbmnhBHbmfMPBdi6wO
VOOl1+8czfP/1ksKYLUatrwkwwyJh97E9uECV0y6ciCo0bEE46yYPQaXQz9u+35a9JEsWf0sfvwc
99ue7lyrm0w/SuUnMH3f7hrgL62wSPm7V0QkicwqXo9Occ3THp1meW4L3FDnytW5LmH4df8AVOtS
K0EmL/pMmNd3Nb9TwMPzDWMRCEGceoV6PynLl24UO4gAyUAaahg+rJcywzxEHHKi7IGL1TQ0edne
bMNw9frgR7iQK64e4gZjxF3IZE0yIX4ZpHch6IpQC9MfX0JMxuXKhmx3O6S6EgS0++raz3kuxI6w
cM1G2c9Kjzf/DAujEuwzxviOFYkzvjg4s0IRMENou0MB4U6dLNp9BlfjcyFvem94BNFajm1Dtk3y
SXNgjjRWkaBIcsyAipdGkFk1emxoKGGtxP+8sJUcYaT/UazU6ND0MLrd0mBzYZlFiSXQIQM4feEd
FONQErbwyqpNy/PP/Lzy/GXdoqaNUcsngJrTYE6OC4NdmOpgOdjEH+qtDrm4JAdHQ4gsjbD3d/XD
ek4LqYLjBa3R2+XGb3fMezhU927itEUOf9OGM/aIQPpsgQXuppkeTRp+8RvlEnGxdQOG1yzOIoou
gXXZcYQiz52IdcgxFghvy4zH6UIk3aPmZGJDcdfVy2r33SYEM57m+FPIM9teoiG13GgOvMMlZ7AX
gz8wmperNZsONoArydSozpvRWL2sIGSnvtpo8LP7xyYCzIB4qh0Fzr97r8Fkb66FwoNNxC0KDCsN
aoqWHV+93jguapUHlB6r3CtqYsIrbAxaC2hkHDkeX93zuiWnH+i2QzG4S0609GmAXVdsf8b43zUQ
fXCvA1drmgThweA00mol/I7myusCIzGBQymRM9xjfLa0Ndk8kF3lE2eIj/6Y3wAORrgTc0ChLftt
fOr6aHm5FrgkfPeB+pmPz9vw0HMpTQWoaDExjTvPN2jZ8rb932KyFl4ExdfLtc3/VEXgCbrU1pAX
XdnA5XaDVTg8o56DCKgsTAUazXhtL7//b5zRvLpY1TYuEJQ7k2hitAgOhxUY0o7bLMqr1gF0v/jm
RcHkPpGlakIDOuDC0gXcIXYDrUcKt1eOkehm91sznI+FrG3WYJGP9Tl61eS6AA32dpwmL+IP4McK
6bASmtCt9uKvuj3yhZXSfGldB09IAjO5N+5M7Sa14GFceTqMhe2S+rKUt5gFKFEtkwRcYjGrj7fG
MtulbC8AlYKbwHkNfpjSbrmp1+Yo9ijFnrVz9Xvfftx2q/2dBhGHGUoxpTsDROmZ9a6L1QxiEjiL
EclCxEJTwxwHXzoU6nDqvuWUuw1ZFFww2DAAvPvH42sXbDLguigYnRJFQmcel4Dav0HC/XCQFj8U
rg7WKAkWKm2k6qYsGR+mX5Ekdtx4lTpt/no+AnpQAj0P40GAGRjTHWCVjspJpfZlHXHWDJ8L6CWQ
rEcdcDWAvT8pTRkZj7cb2oy8We7rKvnzk3bX6ErkSKsf6yFVoJk/gXNAzhQg23r2WNUbJcX9u/0p
z7RKTTw7zI2y/1jZB1S/pacZWQ2g7fKYigUAe6aMANCbK5jyQn/mpI6YDH8+87Elyl8zQOX2WZ3b
TSIGqLHxkhpFADrWmt8DFfxWamzIfp7wqlstT8R6Pw3pCNJ3T55uLB+06TsZnk/mOuVwLS0FC7IW
Vw42w5BZpcEUOyW5MBFnxJ870Muqk+70KfhQABKEU46+sjmdiL6KXfh4MCguBsuEy35F99tE3/A5
iVEoy92wC7BJFrn4bRhbDx+bW9woGqN1y6ojOl7/jH9vRJ53d5A/pes06iOPQWyt+nRaJyMYjpM5
1ZeiIzPBcP+r2qlsBHrO/PPWml869cwmlRAwptvfvWWW9GphrH5pnGBtLjwKKE2I2G3D4rBEH+SU
k2HiruTXo2Bzs6vjKKV3wZHNdu7WnMl7bWjrXhUHeoRVYUJENQKHxcNrl08zWgnxnSAnIwRfPh9b
2+ti2o314A6Y3zUqtsJve+1rdkpWu43UhKFVoRd4UXKA/dsFKHbixEj1rYmXadg7zWIWo/DfB/cm
gocBrroS5Jz74Wwiq8M5ufily92j1UbvGNT49sHOwzd3omSVL865Xbwog0u9sPYSGNRic58spWpK
mBIm3hf6dscd2RxR9h85Kj2nmYF9gaHzs+RA46qQkcVo6lYU5rWY2Ik99dB9krRSt9Z2HB3OiBgh
Uk+eE0uYMud/ss7nweCaRJ8up4mDK/XkIx9W8rFfujNjZkhti9hefcBb/zSL7Q/lHKGCf/pMuWmw
RPUgPhZ+fflA8XvPr4GSNDZOmwvASqMz2s73+BGHZmH96riOpyxFG4Pmb1GBVUiUiJkvQzHD+HQ6
vQCC2oy05I/Mub0EYuNb53NPJm03QaAS8mxoqMLHoek4WTsMD4Yrpq4NSgXUXpLKRMPDpp5atLsA
nlHftTqP9/xMJmJy/8FMtc+/NqgXAoZ0069XIfVcXrX16akWyxTHrmerIMH/ODC0r8kYlYV36vBc
ofXcyVkTh6sh/yTZ2hyVIY1k7kKpBORZRzQnhk5oelpdAzpWGct+u5IdaweYaBzqSInPO/tVoNpn
+jG7qXpYIiZN7xY+nq8uBSa6iLsgD/0VMtlssj8mljIf17ukrhyZd3PludiTYDNk7Ux/DQyq1xHE
OwFOql2hrBOOOb4Py6nEHy+mT87rtbDQ4HMujUXKZ5jPXqZJiAPEEpmY+J5mOgygCsHHuu11QB/j
qkYbkekVfcfytdKG0vgOnDeatEtmOLUst+BDVYUgSCoVwVbalXTiixdcBRtDCV/M87oNewKhuL3N
1YYCXNkl5xHw9COmQipjUJYkjJa79VqRshYaoYPgg8FlSB0cpwpC+MPzZAiJyFGKpp4UGx4O5Q6e
sWBijoz5FEi4wCBGu30YeGYluc2lIFyjTTW27ZPPAw2uHjc/OiWq/oLkHb8pm1xiB+CepjQRRzib
0aSlhGKBsnL9dfDFfPknakxGp13sNfS2YBfFB3VD0CM3MRx72tVqO9R0NPW7d9ajiuEB1TkT1AZW
XcInELJOdrjvg+FqbDTvk3UFGtrkSdJwg/uB5b0HwgKg1UB9qxJI8AS+6k9ireIIoOK7xCFcA/M1
7CghF62meO+sd8teMqllbHwypPtUy8fOFGIGb4vEeonx+IySr1xjrttkbR5pXTzNkw+5NnV0ef8M
oLU5IFu9W7F7FpjQnlADlR+WSquCO0X6GVddkIQqiIWE5WQzoUF6LbmhtXc/xlXZueSbsxMfEUCV
lYHKCdrokAPvsZWQ7vcJuta0+dwRjKOHwwuhZVeKTJG0ATbTVuWM8zVNqh+OXtTMg3Vf1zOwe3h2
Z6dcDdsPb3fj5298I15FV8X7KWtclMm8w8saAqa82GK+xFrXFm+UZlPgXATDZPCkpJyaekKsvzht
jEAT8SrpV25rS31m7sBJHy9cdLuU1H3rdEnabTxZofDhWy1EWUnDqOnzpHN9Mjvfgb3AfbnUnWuM
EUGiZWsrWYA66ZeINpGJD5WDSEZ71u0oUxCGe1035X9sczWLTwiFZesqS3Aml61JzSK2Sze9M1ew
XApXN4sY8t0PzPBZVse/yoPIa09Le7R8t2hPSmlkE6XSe1Xtrtc6rTQmSLWfE0VjZ53jZeCB7fF0
HrZ6YOoiet6GmOfWhQxrLAAYRVUsmnoHHhypOqWsE55HwVZgbpHGn/laOVYIm183XceoK3Z6aYTM
1Sor99Vv2RnZs5wfP/CEt44MJYKBJa3cOmmD/W/0o06SXUYsikqabhsWhSJOeQi0m8Y2Rof+ykks
/QHDnXbJ+1GjmlmsJNcf6vmiigSjGmQcS8PvPFxf6+9Wdro6nV3wcSEaQwwSAmgs5l2ttl5o3oGM
pViWTKez9gplVWxXEboSyC2+dFnW+yKlfc5lznvaCSgDsQYRKVi+NaEvLFZB+8F87YVi+kv5p5TM
c2pRZftX5SSSjDmIzct7gfKiULoCkWbPatdy4wvKd0q7HxoNZOBcSaXhFkTJTaTXd6T2CYDgowCa
mBIyfQHT75nmaG4gYr95rqEK1H+o0ywo5Bk1KFjlwaxQoQ5jAEQ4Qw2E4O6VDQPvnFnbG0nQaQy2
U75UzVAdXBfGHJeYNPc/DYKxlekyC6z2gOlranJXdroysK93Tk4Snm/p0hFgxQJlGG2fBieF2FIi
xjvrB67bxYIdtUJeV/WnCg5+QodccOqWjoSFzn8V7XaHMw7FXpWu4ZTXznSHOrvu/06khCp35OYv
W8gjEoE0GjSl+u5Iqv6uVEBXyCxyM0d+02I8Lhgk1mnoHfSTEXMB2cuEe89gwOy3Sfn82YgGFYvG
bKtM+PoaOL7UEa28e5+7z58tijh7pkjKf3w98hL+s+DVJdcE5xUnWrMkYse8B7gIIBfXFZJDorTH
tpL3bhQSbNMGh2zlvQGli6jfpT1i/S9fpeEp5aY8SivL8iyECreVcshWNB0liCQbLAAY54Fh9ZwW
bEAdTsaBlgRAEohdoX1ZjkVCe7QTg/Fdocmador9Eo1aGhIZH4xd3267OLlW+lyXURsb00a8d0Kc
YsQnkq3DH2rUNJjLInCc1qU7Uzx1Z1nn/z6+kV4rgf4FpB65aBNy6B+Obg1I8Ghbds3U4kEGCjBH
B2tpp27AKb02yndZx42H3zo+rb9ZNKONf8uzjNOdoWD01bXrGekys6X8csBlzcrOBNAAQr8+yEx/
C+V3FaeK5UPoxZ07+QDKC6RhmPUhIgCjIGLkcIKCuOqKu45hv1X85dRPh8XjS1L3j+VMwB8OKICv
PmTS75xv6pp3eB9QbmY2YZ3WzPdhUBKrkrZECk3oWB10QMp9XUdwy3rPUHHCepakX59Xo/6ESdAG
Vuz0X20PmHZsifJ8YOkOy9a4gaU2oxUvYL4XFDlLjQkRcDMe0gtmD3VfGefxreIsd0RxMWuDO7n7
u8i9kpILFphhGzJ5R8R0yDmTK8QJXoPBAybtxzU/dB9AuSZSAvVmQ6RbTrbmk7Q9xnlzxvWSs2hw
ozIHSUQJJAowbQoBNC7SFw8OX/E76iA54BthKF/BZjTGtu8jg8YwsQ8RI6ByUo3eGx0hz9n3qik8
xylu+63MKqGfNl9kadVdoJEt4TjmvC6LS2rzhPffUuRdVO/hbsfUtnNwFUSdAaGYPgtg4uJ8v99w
ag85RGtER2DplYu8aLJ17PEJrFmtm0pN/2g+7Ku3UoeNoMf5fWluPVPGbQZyvo59RgOE65sJtj5j
67K5geO4Vq77A4K5DhXwuOx0DU+0TmkDCzw9Ce8Wyo3316m7yH5fSzU6iKP8zil3yn7sW/5xXtPX
wg1mNf0HLQgEgn4MgwDbb25dkX03pm8EWTs/glkAqoqwPfzr1TjQScHl07/ZzNJJT85vOvefwhNr
xoCGTdafHk3MopkX8Vu19FKR7tW/04zSE7WsJpo88JYFgjyr8vg2Hl09lvSEM5BSX4RBGNIy8zxo
69EMFjC/9ZNuqyI6RP9AWNpC0Revdlw8TOtPXD1DJmXQedrWMesd21gGhcmmuf8amQCYQW0xWKch
AMHO76uaoKsr3OnBUaA9k8ehkTdTlakQoYV8ao9z2pHFicWPOxQyR9eU9cF40uiISvyGhTL4An0U
yA7W3Xt7307ujfq8u7Nm1BunR7bdCsW7ksYzja0KZzRLkCTfq1JhhKsk66tcCfDvOgmltvqR/z0s
gkf6MCIbNEyL8ue/Wyl7DQsAACilD2lCMTCpystbWasA/aKmYcGozlDkQ9LXGgbdGbk5qQrdREAI
XXc+zHrM8stN06IGXGaw1ExOXJUl5sA8D21/p9DvLRDQtYfL+d39KZzJBD6I6XY0SZThzml0A5Ru
phltSWtu1mrSZipCt8nzLgdBash5MFigliQjP+p8rdE1AKVKSdg6TgGwVdv7bqQIG8qJcvc47DFN
yiG/2n3VPM+KNQa1tqtVVWgMp+JbVMSdear0LS3Y7ICVqHk/IG4VLxWlrvB3UTJsDv/bZP1tzDKz
FBE/WCXrx5BeautXlWBm2gOrfll9RDGBf4i5uZhNce+BuPDExyYgDmcYxrE/wkIjJweRUjAmwNnh
gtZ6Uj5a0oqZBWu9eDk38JSKS5or7c776FmRkm8se8Q3krI6uOM4OSkQLQBBkz+kL343OXPSTxsz
9904Asvzr7geVAVnr5yFb/eoViyxbr5X1TRuao7nxGAfii79o9cIjXFasBV7PwfObfhjW6moDYkM
KMbf4tC4dRYgRqrAVhrUny/D/f0ZFekPAU/NRw7jmnunzHl6/nK/rpmagJElWbN82PVhYb5AZLoV
ZYez+6oOAPs8W0RUIaDmMCDn8BQskuR7fLr4H1+2lG+VqxT9SBbN1apsuCddBxQ+VLT2oU5ZV3Iy
STn0xH+vmRnkU1P13keFVjf+ZLNrdtFXWeTF+ZHHSCPeXjpTr76tsKueqwmzNgdN7mFXXjexJ5EI
B7seUZLHDHMoKzNMtezi7tEdL33bzq7PEsWNIKsnDB2Hfe8LZW+ybPqRiHazbOZkUufLDRbWPBSd
xtTD0PbhkorPJoq/SM6hHRyz0K9RjtKVPJPdpnrNMCxFkbcdA1GjA5mzKwD+GZ8jUcF2xeOExVts
4r3zsB5lrItMPXfptoN2cHfpcgMujOYMSGpwxuZJx9FDyn1CKi/npD7cCPwnns1NaRw12m/v7y+Z
OG6GTnL2IV4PEzGY1CYZ+lzyhNBnvmqfzr3lJtOmwXwqNm32x3R0YVW5gWtjK0lSl6GYYvfThO7B
FGwFF85YjqpttuCUchOZw8RZjgdalc6KSQY6YpydB30Kc76x16Z8cjVObW9pqcQZJlWnqOAmASgP
3C1eA7N3JGAV9pYLLAiEzccCpi505SF9KDBfX3lTXGsllbRdPYyL0/8wBYNFAstnB7U3GyMLaCHR
pxh+K0fkQIjzYXemg1ucxaPlCna7lOKQFCvG9z8jHxHAr0thqTW8J72dEASVrJ5uP2XeL3XOnM0r
N0moKp7ON8AcX66fLJvHl0brWkNG/DAEMI8w3yLI8wwaUYBt/WCavLs4ifc3kjwTVxbltGi/U+I7
gQiXfw8mJUgc4FrXgFSXMG8ggYlSgGjA4uUR+OFH9+cQjqP78R9nm9UfUG7K+giFRblalwb+Mccg
koQYN+AEaUcBTtPt+MIbtdZ2mNvP/EXaJGdUoHmYpQGr5O2o+fDz/oSEnfckkmKmAv8aU35/1Aat
CcuqeAVtW2+88rr3YBFm36DIxLVhgkzDNttrvwGV5gzV7/umb9GQJk2xqMvdCQDJ8ZhFbB8ZRwbJ
21pWv4D+k5OfNjCq3G7clblMIErQB9uC52TUFQo5AB3n2xL/2iKmY4xcgdG+6fSjH9HssmdHnqfF
Ohjt/VFkercK0MnPvVJCaZX0U7loDIca5uif3NMAntoUz4OmE7L6bDM4O8hjJSCRne2LRTvFEYbP
quQUcyE+LMrEUo5d6z4MUUAM7gsBg8Z/4BcOZ6dA0pb71TY3Zz5XlMULQeLA7avQYNVmZSV9HxiT
q6P97X3Af7k2IIR1Y0fcmgxrRFbfwXNZAWP72OnAouhKemsOjP6tmgF9tpAyjORssw+2bQv7PNdl
TniC+Zfn59zt1VES74ySzNObdfJNs16c41dL9+7wMaJ+z31NqDIUuCOKXXLTcV768JpJNOehZ7gO
HcLW1FmDtXmBxFc1alVxE8zxJwl/XqQczBzqFaJBLgkGS1F/6NVDzh2Hn5SBPCxvIlZlqGNJLQ3r
IJ1uYRgJU08K+vI8vDSykCzsC0FT4k4Vy+dC46eWmBz+MIK0vO3rleLN3cueBPvgl3rPsJ4bodbm
0gh79jwSimYruP4CG+n0owX1vucJR4lFYpg+7neBQkQwe9WHNrpi83JEktc/c8f1TDUUX9EzKGpL
InBpifDt9cOxU/ocmfCg/xPnA7hF5K3fNE10VcWHBsAJWaQEYh0eSzpCu/wjbD9RLAe455dP1kJi
9T7k4p0ELihJtxsxCF8CL+j+pyDDjRHHuwxXbotFMOFEvYBLXlMmnGJHntEQeDPTK8tOTm2GYGhx
efDJmJHUVgLiLnIKzqO8WCj6/Y0okWp8aVx7Ag5Xkzw0jcGXrAOgP3wgrwGvgJfsu3CWDLmBloDM
e1v5KOs27x4vsitEqwB9a6uDgTnV6cvXRQKk6VlEBV3fzJTWjQBjTijw4JuuURpOA5NMFWWV7D3s
R7nBivcsraig3SGMqayDEaoDDKZ/DRFV67u6lzDdxgAseX3ajEuat94HrRpA5OHMxteaxLEYNJ1q
8fOdI6AQVwRI9X+bNU+YdVMU0EdoOCvqFc9DW95RNanoJiIjI0rlAAd4fVW3QBp7Gv8LTkQW1zNJ
TnGqbkwl6tzhln1nAwm0h3CS0oU5DS5OaU8hVIuPFbVlnsGRhXj3a8L0DxEeFdO8sXj3xm8nOTOe
VNnemw5jNnNQZA9a14VA4LftVlbVQPgwflZmG3ufqz1aK6eYOiz5Cm8P0GU/3BwsxDrvM+TCWaj3
B6Tj7bms7TPhSj/sO/jEOx01Oo9sWm9pX/7HZoIHn3JgT984UQxV+Jfq4CeuZAWNoQtBROfKev9H
pS2r7uDWJE11OTPBkKAvuQ0UGMvdw6E84aXFRs4v3A8b8f8fDEuLNPsZflkM4HqUFUtuz23TH3JK
If1Exdjcmxr348uX8I1U8FUCmkK33zzWCZnf9OF1h41zNVNuIJ2kzErF4OFbY7a+MEYWDv9d245V
OXYwsjBkcmZU+KNr9C8ehZiRORBbal4xAn/ZeSPxPakQL1YhzuzHc3g/1psTYqofKLgGVQXwT1iF
k6Sk1Y8qFU795UdJlEY4Z7amPZlHkH+YQp96o6RlZzn7DRqoG8G9Nhj+ms3BuJ5e9g9VzDNE3xWk
ONJJFuhwX6dbKbpBRLdg2znWQLvb+QKDYc9n10kVlMnpNsIVskqKWdA9KipYdm0N8UGqafZYEUMS
f1lxL0dXm0SAZtB1Hr0wVH0pSp9JXXBNmdkCMaKj2CC8Pp8A2ydU5ufV80ZA9Y40ql8Ba9DlLkrU
KMX/xHVsvkPSHxPHMu2v+WqDXxjsF4UkQNj+8BljLQc9X2aPZRCA1aefVTCe1vTsqvXMfLgEzPj6
XHNIRC/PPlO8QMQ2aBR695P4aJWSB/IKym+mvkXJ3iJD11H/tiekw1keFvnJkhzSJq6E/y2cGlXc
soACMFoVGjJCsVgWdk40e8xPuR4Pr9OoqnPYljOIGwuRcjfxjd+4V+ej/k5p5PJzUdPZKxiAU7CD
BptK9yFNbTWGrMb9Z3NhNu2b1Idd4Md6VYl2ORyuCj9LwRAO6CUiyCGI/j7WR4TTsyI60rxIhg/n
5iR1MkQZ4nlkwiXLmNhV1Lyb7kw667+BE5OL/KL64EhvmvCmNG9aTI6QXjlI4rk9sDJXF5fTym3t
75/nQOzq0GTri6sojzonT4Ncire/4GHx3mTNEu/B44+V4dxNNCQtflQpTdBwhLhjMzsXJxCL6OMC
yog39XkcZy5dgxQxDmOKdobw/XUelfSZ+oB01zHdxVmJq9MtRoxezHDsn+huCLAC4DbEQZ2jrRa8
RqxnK+9QbLA07uhLAhZLKyLE2G7e09SQ3kJKg1cJQGSeFhKGt1tWcezRvL7X2w6iz1Cfr5AntZ8D
AY/U8E0lPHXC7h8+8F1ALEIK4RWcbjck3UCFb7r8J5jfNvp5A0/6Mg0VRJ0kVwqfM3UwsoXN8ZmT
UuKMScUI9zjXJLVl1VxdlrWklqZtrixL9AWyyry7/2HxgTx4LY4/zqcYacR7vbQvce3rNFXg3UI3
dfwEH2kedAePedvEGERL4JGxGvAcKl2/sI244ZiueepsipU89f/Azuh2HLUTs97FsrAQ5b9/Y4Hs
FYB0j1QZjLNid4xVjpH9Bb7I3BZ2leo6d8ZjgbejfuSvHCbeB892LsckEovTepUKMkgK1vbsU79Q
8cXyu/hIpdLXcdCbqdqBgeV87ury4L0d/WyNHsxcwa1Kcp7c2lfDI+v7Mj0M80mF18xsAkdmn/Hd
wArv20lfzb9U5FsSpXf9cj3pCwA7bRWHzkqauvjShdozg8aN7KQQVbnTJXS2VTnaOR/DvGbmohYT
VngdYPUPRXSgLngh+Aez79TYLizQsSgb2YFFuJutAWVC9O9GOeLcd2yfOwGXH/ZMGfs/oUSu3f9Y
gjlxeXEk1ouZVG/F/dS3TM2JQFiAPROwu3gjqvADAns1uo9T+odKjRkUS/jH7VGJc9Rn3mxySNGt
i3/IuT6zTNzVPZ6E0r9Bm7R/GM+8GXQHEoR5DLdac8NetRNcBjPTvWWmeau7TP7ySd/4q3GLhz8Z
6ODMHAUAA/AQOeJrYzCy13OwS2fpTdQWeyNS2nVG0KMFV2S8ev5xtW+VykUXxtXB4EscME892+fV
ug5MEvMzSRuVmKZNbPdn0jpalHvEmBaV1ythm367t6C+rK2f6ywXrWlMiI8ajDF13w3SuGm/8823
h1MJJ/+5MuRKJDRM/5I1VZQ3Ewct5WcKrr8wXMtX4IP2Kv8Lr6PCJGpEMw9EuDywPid93nuXFc9m
e8OxWhZcpaM+zAtK9Wh/Yug3gMva8fFDgWxrugj1bq+5pHwz+eLM8detLwyFRNlI4TeEAf67SJ9q
L1sRuKERAt0T8TRFbTj6AaOq6njztAl15IHbB4wKgKlJgrB+RWKWW4uQoiKAidOXeED9lX6RMGy8
OZ5+rzl9Zm2WrOQ20Y59xTaNmEqpbC7QNjz74X3zZvB9PoFPHKs45nPoS7TuKzLc2hNYWNXCElya
J6VzEKLHA8kgYmFIM4d2q0ksinc30bd5bTBPc/mMCAFPGDVKsQTee0kOWDB6oKju3a2PBPkHEwfj
ZcJCpQWC4W7tDQ0fUHNaR/ZBAPukeJymtEtd0C/2cdg1OLZtlqHJxNfmbto/33m0i5VOSXTLjFZN
5Z7nKLRWOVyWmtScOB3c+MdK8HVruB8hHHObWqXLL5qkSg6u3fFfftfMzTsqIusH5VKXXVLVpHCI
PglpZ1IS2xvtqeNSKeyvr9DarIYPDWNoAjmViGSxdathqceDD6blaisvlEZKc1/yZufVAlDb0Q/M
5Y1FkaFw7Md+og9PUfyCLDd4KJYkeDWCwr+aksadFwRlJvBFfLaPsRbu7Xu/RP26Hc7GAjyMN/Gd
tCyvYJlUp26YTL5U2rcps+drTraVN7jYLZFTtMB4EM7gmAveVAG7Af8KsACAWi2Jq7F6YjX/e1EI
zPcq3IMcS4VG5PhuN4GWgMriRoeoZKSoz3RRSk7DkrXGqd70CIk7y/XQhZ7afILcYJNAfKEFXCGP
FSm7Xj09vL62LCDC8xqm1qNaQS3OU2IB5G2YIoJfbXiKcRJKtE2j8oBeXWWp7bVqSjm9U1DkGWkJ
KMOpREIIVEX1XTsjGWDaX5AcvVyWzNEHeFvG+9wGaBuZ0A+Prmp60efYTjCWYaJAqg0i5Fi8bLU8
plZFGW7VtpmTq+M+Q01gHdDk0ECo0BeQoN/TIWWQNvbEPR6c4E50cvxH+Q3qZr6toXmHIFJlihi8
rZEr2gN/BwWzWt7T+oevOg2oxHOCpR/A/mdui21goUtMrSNe2YZBFjnTFBkvVSGoVkNrKZ45HIQz
aJw3g1HXI81VY+aqyEa9i8llEdHXuze1UGlaft1EZSPRaTwEBjVK4WS4DQIarBIyDnDK719TDkTm
WkF+jsy3102suBW3E6U+aMR1CfrjnTl9sRt9VhHPsw3+jvxYVNkEP+n7TmG8N1PA0zppROoO4Y8w
954P/qShQvppUUN+1eDZ6ax1kBCwojmgqxMi8s5ZvvX3pdnuvjWae3hEtX2L4vTRC7ttU2yPNC9q
ZJfFzX4YsMJfPEnFHkevEP/vJj6zrQ2bFLgoPpVErh+v6m82RumQpGlo+rrxzfvCIdKKeshtTw3j
I2WdaeX47ZkDMoBOBJDzFOJO4TVQAcGABUeDqeFpav+6jVSHb2Y4LtPoHenohqC+rsUTyHfZLgFO
OKWChY3qsjl4IICdIWpyLgB56HK3pQkRI+XAwMHQViMl+kq5UjSDixDfmmCcNJXST4HVX4E6ow3p
c/15deeb0QsRxypPAqScpskoSz1w131dc2hGZ1+nloLk3MRgLGAplQM7oy9fwkO7q0ynA4cO4IlU
6CdshMB+hHXKTLdQ152DZqvVFkDSJFfE7OcG15XbeE3iWz6NmghH/NspFpBFTvzBMaW/tIBcUEsB
e8BiHzW1A4JWusUDwWz6Slu6bBIKNVcwLaBQuxDxfIyTgy/cUrkL1G+yV3CpgHKZTMk+6ly6lCEr
dT9eRyQCGmDIq8n3FQwsvtXqiMM45BMVp6mqd6lrgTFMKxe1QWJzKZtD6YPw0M/OUk3z0VtkVTBi
guRy51ZbKU6oQUTvElNr5hcYDUUMVl+NVDe8KXOhTdn4Ry24MnFVAW1sMc1UkiGSsPQeEUSb2bQQ
UdUR+mdb1FtmVtvdTMcO/o+GU1SVRiMqQlFpK4mixs1HCin38QR40ANYzE2RAPU3pTAKPWH8XbBp
qLgnIiXmXVYn2XxL2why7xJwTJdYYOaZcsRIPSYuVb5QMyrZsM0P39RKppDK6+Rl+qy8JIqkIPfd
25dKjYghnBRlIOYl+r0LyM/OilEeVF+MuABsN21Kd6zv/Kf4O9TfH32RFXXuV66A3BcyDUDgFMfB
6qq8GAAqVBJVBEWOsdO46P4b3Bk3KY1Z/WRUYG4TInSWduCwUvVjCa7zRTn6m7bBE0xXcYfxhIOT
0vTXtuESd3+LZ1jb6DXHzZnvF2QB1/xQNCIOidOXA7HbUSMHK3vWGp2K2cISkxoJz1THAlBes89D
oCZ4cikxRLSXWn4+JkYxfnocPP+nGaNc4HRmke0hediFM2oNYnBf2XdIHEgvO7eF07/IxVCcyqZf
szWYcEGuKVKnHCr3v9B3tK3ZA+pT4MBA54D68+VTl++CmjpwDvpQIzpBXJ118wr2/fsrrpTHdQNV
Sa/ojrnMkQO3nZebe/w+Sa40zLDnaKWY/prYiLMjGZvwqWJdj1BhNvcKd5zk12U0t6npoFgTffqn
tia4FO1lBUvEZvfULhdWKgKkkyUgZUbqPRKDWinqk2r8e4ZFtsviyUo6m19WStIaiCkLOTCRVvaE
7VZDcHYVxFFY7A+Gs4GE3imoHksEtN6LgAnT8/iYjarhY7D6q9ERSSp+nzflh8IPY+CBCgbXw6+f
e6CmZYr6VHUQJtc8DiPddC1FGUjGUXoCXoWwh1w/W3jU0QimDAVwWPLjLuPDvuxSd59cln/vCKQf
24xco6u+b8+lwsk1LRoIvTikETN3nVaQTTrGfDPrz2uIc/9tBnOMxiPnh+6afI5IIq+6dQ4GGMXU
dU2K2IAFxj4tmqwFxz5W1kKhzPSr3SUqzesAgbRaGmVDEv10P8AffSoOcZsGEmLxyuQGJP9/tidg
UE+hMvl+gIKjmVkbdcxHbkqsWtV66EPU+DqoYci38AKR/HWEZsDHGq+jDgJpPn8/82w7Y6G8x8Kf
GBa+xxLQOmWsxYvqaK3CL6SJFfnvhPWZHijrLPzqJ/UtkaX49/ivIp/wBzWodLJCelyLytc/dz7F
2miATDOq+CZWAI3isyOdqFbvmGBX4oW+R9Ce5ktkihKR18YStuzO2Fibka+1LwTY4m+VCLxN6/s1
edgalhzBfbw5dPRvRBxOvuDNMrjFGQHQbtQWtLo+/AA6beRPvjn9/ujAcrOo0JP86igd1ifLSoaj
PngtPckuCv4nxOi3U86riJPaByL1eXI5ASzziiGpU0+t1bGoogiu0pfTMVR8QNQD5rgazoDiUr01
sfuUEc1jdMqPStpEanGPF2J+SgaSQc3fWjdRn0TZRcHbMC8Wrpnbhp85nK0SoEoyq/m44jTVV3K6
Io78JGXOLMMrZpxv4hgb09fWjuFB0+bT3bBz6S6tiiTCF2q1g27IC42Ad3H1rc2B+xwPiYBE3TP6
P/ths8ezOPg3qj6+UXJtrI5qj4eq6W58tochNMEbIlXICMmtRnFk1tZ5S+mVjIoT+ZtpJ27gfrUk
tQg/rvT0RaY+M109AtZHbqgBi6szSy+/sfE9h64dHZQxTcAbH53t+3UnIneAHksTqKzTjPJZa/hJ
gV9gSijl18I3eFwNuClrm3sNnpgAlh4/KZXESPf/LcUziMvu5QG65uSrULr/+EQb+o676M1dCjBP
317MuFm3HHMmNZmAIb6uu6z13OXAUsHvlmU0rpBggymJEdEFb3EQA+fKGW7xVoEZsFTOXHo3OjWl
qyqKOZ6WmmUK8/WSmYtGrzK4K7T4aV7t9/+B7h2jVmx6+zUh8rRfqa6MsDxi38DNqFX2lolvRtLH
ZacirHcOQM30BP9RP8rBYKJ6R0jXqkVr20TMqLDOzHYHQLIXRhGmdupBrhFyzz9c+hVHUG9qGf7P
ubH6IGSZ9NrEIAt1UGChUWEKlHY/G2ciCUa23qYQ4y8jw09wVl0wYG/Ee4RHo5a3JcxD7qBG1OBB
4ruJ+PuT/aCGNeHyuxs8FCJnpKoQok1wVpKitJzDVsL5+JktYAs07Z29gVOlF/Yq/0EDJqLShWdd
7CdG6MiiqV01vf+h34UEinROxWVKmJlunCsEePxiuWeTD0ZotGVNvp/ufrUWwhweOK0wr6SIJovt
bDscoLVEadIQKTnhE5+ghFu5zwRKcdWRyuDagganzsJ3SWtRKIvgdM5L2yhQjv4T7rPwmVeBL6MM
2qupbssqU0BrakLbqamXcnToOMIQQP4o1mfE2GWA8BGEfqRoTixuHWB/q3KCEQGAt4iMtacQUAle
57JC4VCXaGeoxy8ZFhUjNXS/0DzRQEBbB04Z9Ig8Gd5029peJEExZPGTVHSSMkBLf99ULD/fctYR
/+TlHp3PbqbegKbB2jQt8QLP+KW/TJv9WA/eIzzkrWrVOhia3BymFYXgWyx916e/afgOvnDguukC
PDYRrPIkmc7dRmydZcwlat0x4xROHDf888ktNyltuPP/qV64J/YTAyeETvAEOluzOVBbd+FAwtrp
Nqbxsc0CdVPeTSq2Rn+VwwSRm15QS1opaMhmUmB480bjKg5ZUEycHhAyCbznMrWwK8W6ekfgtswH
vb5dPrUusjOwm8O01n1eindcfCNxpY1prfeLpURBagDAlnhp4PB/Hl32JAen7+TZ/5mW15jw1rwq
Ct4pBWvHTwPX7z8HD9ciT1mDn3T61MH433l018XBIAnjShmZ8fYcJg1IPjXSTHL3q8OdSkhmzATZ
KHKiiBjF9s9CRWAXlKROxtPa5xnb/k1kB6gItcXu1apmKwjtlwk6KnLEpM0jjh7KFkfTycAr0UF0
TepenseBK1Gl2NTJET35ldkyq1kiKahWSDeJFmN4gI7OaoRA0oogfUpZGzjcQ6iy24ZGjcplJPMI
1hf2p7b+POIk2fWZf1VRtS4CIcBgCr5C6cNURXaHnoH5c1/huPexlA55Kud6CJMJHsn1hGNntetX
cpT+DjlHeioFrWsHc3sO6N8d+X+euzvuNyvFsRhkrq8UL5KWunCpSIOzChln9s1IwFbpyvKhAJzT
fvKp8WPP/KLiFSOOCfwIpTlyrvcuFCknBXQYxt1i0g0I/dwihbmwMs9mldXSHtZ4uelujVAuYicw
HwxELlPLE9huTyx/dPabFyUTlrhONvztGOQ8W23SJHvOHsR0ceBgOUYd3njDYX3lkQ2pouko5Tfw
AGhfBdLEFoun4tain97/ZDBgfWZ1MUi0Jjj0ZgyDav2/V2z47eBU0gNIjPvJiRrs4Dtkt2+9UOrO
bqB15K8sNAE5fESHdBYQOcroZNgKsei0ryWShQTLMLw+sVAahZbzxcQmPueiXPlczWSyLDKVsU4k
u+ROadNGYpRwBC6IARXudTrGK48a6I+3vm/NRPzHp6Nd7GPJUFhU2P4D6ny22sRl/xj47mVU34rK
wP0PROPu21hmsB/ql9iXCpGNOq90iKwefN9wz2qXdr2pC/QSk7EUbsrFouZApdkytu45dmIX8MV6
tcvabe+l5/HS1BcLPpPjuVogkjVS07f8Oj3Eob95jQhWn+ueWTowmeUWrd3nuNhrO1cAT8MMBHe0
pjT09MAzXunFHZNKYtyA1FPYXzOVfgRujbRW9r4z3obcw6nglLfM/Y/aNDYKMl3xbOaMaO2ADlEV
5RqZy6JmBr68KJZiEcZVA2Nx61aPFmnS0FGAmWc9jWhc7sgo0UpAtaSoKc1s0JzUxNQ2VKs2KKsF
qNdFL9ebeqau4JxpYmdLWtssDIkeT2NMy9AUlaUxlk1i6aUdJsv2CF/iLj/SkdeqqneQdYYijqwm
e5AYOdYYBMwEuuEKh8f2Vx1c8DjTy3AoA1Nxz9CCSlaiVhdeuUnnz6T5yBALrLhze93BS3rpQkm4
rnR/QEBxDqDHnMYQi0ray6nPlRfhknSB0Vhq5CHMn4A4roSil5oy3s79qbF0k7IJo8cPwxsKWaln
x991bJIR5vEUq7WPX88UHc3gbdl43fdEEizDtnw84/+gK5mNx60/ef0hTv1jSQVCkDQOmYP3px6s
EHd2C3P3cyOj2iQRPuXJ/FVSt33hHy6uzJ83fnAERu3FKW4MYQ1DhLVcK2TPnIvKjj3KToax5ajC
i/ajHVV2QFSYlanro4+I3Ayb8xWctSiZgVZ/RiqfN1Zd5GE8LlLqUZYqs0aHzjy5dRnHZFgsf7Jn
4g/nbxleSf9tLrK2b6n7aoUxfUmo4Uge1+46OKeJtjDHr8sBHY6xPLvH49cII+i2yjZot34JS1zR
oBVZ9Z/MPsxZVRK/UKx5NtyNrY5LZrRvcwMrP2v4StrrOJbS4RyoXzeOzl6l/Apj1lnX3h+c5cmN
uCwYFDJP3DLmqYvaiBDwtwLVQt9dIjK5/msZjouP+VCppoe2rDHdi9jCh1XNHwsWvWhmNTymDoUg
hg2HaxpsUfXrYZqUPRFCkAB/Jfb4jPTj6UqBdFoBk5EtQ9ZxMydo0pDOVCabl8u14t3F4H1R5lvN
Bb8sVmtLekDxzoeJ1tgHzCPZnLucvYaHUnr5yq9FxN/fq5Yr7dDzPr8dQJNjZzc/0oLT8ZnAqzxw
l/aAKEp9Tx91lV+VU19C0ofYNWYZrH3qIa4/276khedkILdIpkdZIDaB5w+c6j/Eoj7i4QVEbBP0
xcKAtj3015G8vFavh9KPtomGyuKe1HKOFgCCeCjcHbELxZZkkddlHW9YuLQMq6hnGhpoWXfbqrEP
dNYCdjGsVFV0NqficJoL/09e7nxOcSk5iaUPHAya0t4HMuCEXDvO75eb3xNVIKiFOCWETd9cQjuE
Czc++wcGk6vYWxJcZ3HvjHRvjB9+o3hD1Ok/4Oy8qeOm3uhCIDMEUL7tpsgGqvuJn6APhQJpAeQE
y9z8UybJcVfeA+B97DFeh82ceQkMCDDj2e7rO6TPf+h99M7EZ+M4tYdn3E/sqLjpHSpbAZxoBis8
Z/Lp/3MmHuoHTEcyqdAhzzUkFsQA1/oTuRdOiDh0aV9NoU7bf7ymQfvpIGjRU1rjULXTl6aLXv7/
cxIN/dZ2tfZtXsl9k6reA5fzVcyrr6PzGtclJXHr+6cHhws1v1ci2bI6Uf3qvE0fsgjh2Caumvsf
mWAas0kmal3Rsm3RnIbWe8HRYrqsNtLY0O2qb36HUjya2AxUGR7laKLZugSE6eGI+Cry+2tqaST8
kg7d42YKXYSg+IaxMvik3GVR6qD6pGObYpCija2kc7/lW8nHy8jhkI+5FjldstUgvfVpZPNyMb2X
YY7Y/jqu6JPRD0DZlGaGdDlyv58vip+r+W8it3WDvgY6zDaUEk/KAkbwQfLbaHiuEJNSI9DjCvW/
GRFgVUUZGcfqJ8b0PMmsonGxQDaSUO7qFwVT6OtRH2CHlNpHXkPQxH1WCH2YrDvURC9GNQq4I7LD
yvwayALszrWKcvyBdllRK42wvaUfVBTFjGYkUIrOrZnhiPAh5bZUOKhTp2xIMGqQZ0Qmq/LAJ8SO
yu59HCr/CZXMhvxFUubfHoNt80hRZRxF+EtTmenzvCWGxYm9t9r9bRy6yZCAdcLbilfWWl/MUiU5
ivV8V+v2rFC0DxbE0Yx/E/kqAtb+Go4nTkMgb6U0uJSKg3pz8ljQCG0RhTJtUxgxBF3OmJ+dpULk
3+lA0vpoB0qG4js6uaM70v6tXJvUCL3U4QPhXeoIkFQUB3FyJkR1FDax5oKGMz4ga3b4P3RxtcTC
VklC318OgcPHcNGo7J/qs3PNZG5AxjK3P6zs1uclsYCMUaQovVofRY/+2Ry+5UnT+OnQWcdsLMjJ
8WnmOQF7zlgk/SbhdPgTJwV5UM9IrsapmfCJKrxL7Pf9gZ6FS6TPB9gYf/i6eg26olR6LcDxV6Hm
UodVQhfluTASwQbCUq42Fy3VVDv4nVrhGW4ioia99CwjfFwSrMOjZI9g8dBeZ4IyRNprvyqOMq5z
sK9rCX0TZAsUB0rv+gmrrPlf7FZZ2OrkhX8ssKA7uDhY02lJvvIH0VzPF4F/5YUd5B1tJ/05sSxg
1gRx2uHnrdBZYqlI1xESpH3u+NXsyZYL8vO3VKzKPGytG29x4ixMTSpxVDRyE/Cjz1/AkeR+AYhu
R0BQ7jg9mqYWhiOX+Y11evhcv6U7Q2cN884u73J7XADDMIBwf4EKY7qMv58Z/DaZmoIBcxd3vwok
tFq5TgIIBM8JJcBwK1i+ojF/qsRPpK3Erbh7npbcJ3YHt43SHTCl0Qw9RSAB8FRWCM7A1nE2KNlx
FiRkEHOYNBdkZOh3ur4Kb2LjN/e4zmGEVE/w1sSK3j8jCflUCRHpz4t98YQCHFQJTQxSYHX6g6+0
J+BErB8yzP/zWZc+0B83+xjTdLLdQZ0uRynbfOUmdgaD2a2NJm/eLRylOhFa6JvhLAT3mEkDHDO+
4F9lzuXeHvAjmKe7g6bb3Qx3mVEG33uFlvPTHcGBl3RtBgtxDBvabCa9MGKY24zzVA14Lufr6k7H
vrAMACWy9YEEgd5TUrjkVB8LGfBwJ19nR9FoVmKSgwlLgZMrdcLWFLH/cgAuBu3aZFEcTy9NPw1S
J/UL0ARLiO8k3Ebfg4M/r/fzF+bp3vptfvKi9Su0L1SUSF2xKv3rM2hHRSu8a6tyP3ny4QvnBQT3
WC7rrdF5Gc674bnfzkybOGnd3Pk9bAt08LiDktqmtiuRcG1ib1xhI7jAf9unOqNMtkGqb4t+S94m
p7+uvVZqUO3qPj8Pz0axmCge+jm/fF4/PKI1Gg8wXSu7bv8YAQRQo6JZ+GtSIVRKDG7kyWEJwJZ+
+3Z68gK8EnAff9zTHipluyIvXaNU5erczNFeLgddto6flOAB/U8pXKJZimA13PHN0sc6ime+C8qb
jqgNiDXV6emXDlhofmbFELlMbdH+kPzhxTBcKDjwEMnd1wA3KEi9NFovQfSplBI2iQ+oFb2rW8g9
JhN6+fQS1NAWRuqkwpgXO1KKiWCT6m8fRHF6j3YA/4poact3hwnm8tYc24NVoJLBpzqBfpy4t0do
an1NGXfjmT5e+vMY1glboH2Wuz1/GduiXAOO4wQzQcBadTyxQF7B82r0pBVfmphSP1h449Q+vlTg
AKKVfnYeAGAjXhCQWilF/rd5S/W3fgBlgXzJwtMce2mpoYv05z8nkSwpfsjefFQwrbz6GyzLW60w
XhRd5+Gz8HC6/3+c6tQL3Ie+5cmdgdGVxFKVbcYc/6s7j6gn3S/82oZ/Gkkq8R03yKyE5xSD5Umk
kRjyIt/eFhuZkjpHhpPA8jzfR6Ng7mzKkCuLpG1Mqg2GdFDfxrzat5aAfbvD8idVjUDWNUoXVRb8
VwAadEz9LwyYBUpuRpEqznwaE8O9xp3LWKUwQBUB5FlfnkIwbF40Rl1P41pUbabaSE5QVuTxmc0l
T+QFl1rGxyJJgYMBHm2h/uC5GSWaoHoDUEDd8JNIk1GompDAF3vi+Tz2P4meM4VIemNgAdJxhME6
B6iuNkB7rbq3ht7o45GhLh933OBWztf4ebZ7UqQ8TGlwX1hb8cvFvPunllXM4p+ZOBpy2Kg84uW6
O/Uzr2r6SY8hPyP/FjMu8ZJauPXzdN1CSJfNQ/ehxfPU/7Exfg+wij5+fAZQd7Xhn9QTA01FIg37
0YqWC/HoYs0S7YegBNo9uPKrykB400zirrjgC5DIaYeCkVmJv/3HX5jTCgvn0VzQ5i235m6karDG
+XjGSwe594mEOLujRCVRtoN/F4XwwDSe5nhFdSKZI6xRfb+WSVB3QSj5fWFU1SlY7VSxlIzcmtEP
Kt0eqcb/lJsjaQK0ulMC7hGWH1Ir76kssCIoqyFKpMHlATMcqLSaK68z4j0n7Jef/vhoKONDnjBY
sVk3r4/2EF2O25XA6ETtaf3ku6K0jHjXi+l1PyGyNDi9c5IdQtSFKORByocdXbKYhpht9EdV/T3B
V/Y4qjJaAB+rMWl67wvKX+oG+yzDJ1HC6OPw8olRR9O+stb3UqN3BxZTGODA2n2TKxB0wE8Sav9D
Z1Ub5GFs29IQZunqL3MpzZ3mmMdwhlka90XbaZXzLR52icpIdzJPPRw5Hci0iusDhjrjT4Mc+CIQ
dwxIy5b7K6M/ix2luy4I8q0RO6ayQWLAtVqtwoTizRzRRrsSJWDwte1am4qJBei7tXOm2L/ZNPp0
q97IZ6Q3dFR/BsLBslRh1qNUoZvYO/gN1mpTnF2LMTFkchtVg4+sgtvQyC7ZeeRmd7SpTDy5q81S
vSIeXGudiVmN3gqIhv+wzGVePalxMsr6ZfQbAjHA9f2fd3L7Ab+sIsgrQKe5KzDa+fri/DIT1xIl
i6NNYz1tJrdpAtuM8wCeLcFC0qWCd/mqtqglDWUR+EffIGgt6OnDwSBQodxqdlIBUctNutHo3kcv
pjME13Xq3H3q74GkmA5Jd+w/B9LvpmZ9I/6WObhypNIoSWIfuHznpSYE4wLfAQb8xVZDVk9f2zyL
X+rgP27vr5fNNOVjZNZmCsrzYhBlgc4CXdEAhwGjNYsAZDJ0okBHtryqBfmwUEMbRf578sDZXb7j
1ldvgLZbJLF47NtzfouUpeg+8mcbhWIEnZgN1ypjXvLX2UW/iPb18hn0dL5ljbaaXt6FT05b8XHl
O+5L6fhQK28ctEm5rP3mfLlXj/As9icZ5XxuBitBKxuVO6Oco8uibafQhuaiT+QRjZYi6vTOPE0c
8zMVT0uS9AhsQFHhbcjUOHVSPh63YUWTSUOtWXYSJpNrlP+n3tjn1tC8ATTiyCVsKcIPhxkVMPVi
VtEZU9CK1ugTEnVHJbCby1MPQIQ2B41VHv8p5e06hOsCNGk6afIFpD6aaSbJE+kWyaYLf9jXZNT6
3Ug2uZckO1hVgEZta2qxy0VoZD9CSPUZMW8oXDIrCSjyLzSNXB2FAiy+X1Dyqf0yULL4m0gH66cU
I2tbSYKYK7lL6VVYBp2kmE4w98THHibxiksI147lnYsjNaKKSnYT/t9TboilL+mXEOBv6fXoOaQb
03uvzrDn7KFMnJHPyz7ELzAYk47FUDdyYNE1hPpyPYuxnIZNQuGQPFnVu11iFrtZuCX0tYSTm2XR
D8y3PnB9a6B4Du1qTvRNXAr6hL2VLqh7tkbSkq0sUPu7317fXuFR7X5bTQOt01xfyBUICKqkVJ2c
MKNHKrj6NhDLqI1cJZFTjj+LolsKwRO1t6XXhJHjg4SAL85IGQQFCUTRXXbRBSG3KXmCD/pTXUPD
JsxoLGJi26x7ri4+u5bwE/sRAtHYESZj1KltgZE3DfnkdVL2TeaTax5kwVT1K5uPDKLR6pmxJA5K
HQFkbuixQqnEnr0fSoXTqSQ+NJi2YI+6o5yCnoHcEfc5VXZ+r3fY7KNPdVplV/krWos//NuR7EIA
+SDbrgOr3O82Kl2Kh9leAUyPaeZUe9q9Y8S8DhvKomaekAG90NEeDfWtjkfVrylEaiDgf1hEvgfn
ZEtGTOJXKkfQBCWsqJO5fTpWY4b7v79uELmon6ImRoaUmwZqcibL9Vd4YfBk92I3bUBtfMzifDRU
rTfQy8amv9Az64R0Z8zWZqlaFThK1VsFeY6wsGEJXG+6jV71LLWgep4y1n7zfknTwfOVLMfhI++8
wvbqvhAARDjV/Q1KEJxIVjh0YAQNyHtBvVRlBuQ2Z0SaRQqZPf0chdl0VneiFefrhNUcAGHrfw3w
RAgydX9KzOxwGOm/IDk9D/lkrexF1tVGetBsUHivr5ADnxuDkSbzB2T/0eRJRh5VcvpXTsvhz/Pi
6CfvN5x9Bp5/Jk8h+9ObyYqnC1dhmn1rmtfb52SHQqQWjPhkc6Mdz1iFnuK3sj2c/VuppF9SKDTA
JYdzveGkGTtbfT2lHGRY5lyDGD4UwlsTzPBkrRb+5m7YB//Wjj1A9GsOmIOS3d2cMe+5+odt2lmN
S2lG+tn41yVoznMSIpmTAOYlo5Lzm6JRLvuXl0d5FsFwD6u3rrdDw5ap+jiHwOqWuhhdtGJG5dmR
0PZTJfeHEWwgYpnvadui28aHypgas2wH03VSCNnP0E09lhqn/5eSrZxAPkljP9sjy2jRWOrjTTdZ
dP47yAyZOUFMJmSlKwIAZ7frCuR9Rby3nbIM7tb5W2ZFKi7IWM/iL3/8A3JouJ12h+87P9VxAcNk
Nrsn7He8luBFh6sjhp2TfO+hRVTaLMGKWm4KIG0qgXQEt2MeCGvrIGyBzS9wF34e9JhquN2I+Cwk
eOTVFg6UvKnqC+t6T+KZYR7D4POLaGU2xb8DmdFR78ZqdTvIIsiBfDxqeU+FU+CHPQSlYPPdWqnU
GJz/Ppfk/Pozee4z+hFGOIF71LSe0WAHXckV00Vr4jEDmemyl7n6jkabSiF/O5iuQjGJE0S+JyFJ
UFfWdFWFEq5i8bC+JXI9Jng2rtcygfgXb1zPyNaZirUex98EX/wuqpMdfUxpuUbua6LOT1nfnQZ9
wSs/VP5QG2d8fAKO8KNPBVboPZCY83AptfQEEAOkBE6yiCiraWRQ6TlQEqJ/LDpd8EJoD1hhw9za
40zmiCqq53yv58J4/9EoPUq7H3LeKr6JXv78ieZIatabNputcBOi6MWlORmtB6yEuCrwt/O/eAn1
bPzEC3a2eo0qQeZ1MV/lOIyRQWxpEozoH2eQqyNin+WZEYS3aVaENr5eHzODxJTasTDFjPu9Ywz5
UdraBWbJu0CqBgzSMKRJuHl7aVckFeNFGWv5oleA8QciuFOUFBW5Za6otjgYRIrKwsahFKvD4siu
/oIcOhEnMfXXqxuHLW9TG6+3u4iaCG9tPxO6ximQQCnATmflwabPNpQOzLeHcr32fj57I3Z1NPAe
tNVpDHOedTUJV39mYYivSbl+LXd2+EnJmkWo1oNd2T9ITT8UqmdcrlFCQNCunPYyRCioyAa/doGo
IvStlfdcw7WyZJ/SgaBBxD862LBJ4mdaOFIvHpZt2pop2IQpvxSkgXyfbRIA/w8AGIVRSi2ghOGb
7VVb+WkqCV4orFMPLydf9/ofW5PQSpVUpN2s4WRuNJvn/dAT83S7ii7v9UHqsAYRRSGzldWJAgXL
7p+mIK/usqw6p+lSuchBDTtTxvi0zEm53AEkfh2RaTeBL5lqNr4oTcXYByoollXVhKI+7lTKaoAU
tuxR0c6kNFnlizB6Adpe2YCPbY20zlQae5tpWPPewzFc67+bT0vVbe7/mhVyCzc/eucxG0wkYLb6
Pbajfgep1CioW+bAOwT3H/CMAumNI9YjcsDOhsXdwK75zyoCPFuSosfVTZgR7eJKdPvk8/CeoYiY
Fz2QDQ8wNbBhFQfx8WyvInub7wPPBrPILacDKOv7dX2LHvIjHnLO7NrDNkiZMXzk2lhgFZqS9iTj
hh7L2eqf/ZB8yAooxwrbnFWn51vZkYof/ozutqsQR+/WCycVp5KaYXrpR14SImQ1x/Ol21oPOwYt
/TdjpDsXAcXtobGI0n8xFn08O3LlfTyZl4bXsGu3ta9AFf7DX6nB6/nAvCSjdGSJZ3yX96FC2TNk
yVtPfJ7nRoRrzUWb4aXlVP4jdlTa4uD0LPFAszpcoS60wTExOT0LbWYF4yXjS5tsCHHBF4YHb0V/
pvq/D5eDqkCAXmT/oj5J5GpmCvygMhv5pI0YPa0URT2SZit36B39Lu9eGtWgkn2gozRPZRTMSaQ2
Ea00gYHIomxnWkaE/+ERolFzZAZv7FMA+B6NhFbElrQGNCJ3fs6r5Wp8g8I7MafWsKStpZyT/rn4
hBTtWZHfehm72JJoaFkRU4kKjTvWyeUYMPLzr202vLCOp2ezpKLPrcdSXL/oJDNJcDUNTD0Fv0K5
bzrGOz2cFnmVh+81hdHrBXM29TRN/QPK3oyIX8X3kDefbZOz8GUb085+meXlELGy3pb194cGQNyQ
jSamhc6JOGMJCE2K4qoWz5EqCv5EAlquIYRrm/vYRwM/s0Ecb72AbpvL/oNIQyI/3i1hxP3Ansi/
EDKOO/qe1ysu+qGo0Nuz3w4v/Hj4df9PDfmToOpXS89HkLgP/PFSnfZRNVQtjA3nWERtQ15v8ZJh
uIQmzIMOedrR5cXA74FbTkdkUyoWBV4WlbcGVeuy+eqBVagzjbFB+JLquwnKhb1RrtMh5WYaVxHa
kjGdOKHPGvMsad6VVqU89+ucukgS/vDoaKBaboXEo+65wNwZofRcfpVGDwUyeKNLhPS344TspVJr
7WB7yYnW7s3LlZ7pvuiEUTkgvzulFdziIJ5lOM4FtEhLdf6Yt1HTQQVim6C7S73Zw3F2y9E08qEB
CFjQQMCGc8xxuV/j99MwXp9rnBoAvXa5u7JsWtGIKADp1LF1fox0lAvW3wb7IXK0RlESEOyBVlvs
7McPaNfCJF2hRY4AT8jd1ZeCthVbPPhhKjko/7B3pOi3IFtrPra5bUJH3DqSE94u2AYELM8iUipt
gdr2RuZkNSoFbSuNVfX7ZygqhdNfZqpkPd86tY44EBh8bXXXU0COFfuJny4zFLHyMI4XOQJbPxHy
ZKwMdcCSt9RUMbSRgw8lh0+9IPC2Qk5EThPqUdMqa1l0xlsPVmkpgoHi+Xh4ZAaweB+d9nTe2Rx8
gcDjaFChFaNaV7Tot4ZnF4E+jm60IwjWrM9HpTSMQH5OSuVqiPt+MpUBG6k0gL0EP+axqrAl4kUp
SnU79x8BTCwEQ0bGcK/caWbGBUWzr5gyrZCQovqdDCwkfgDV9kxz+HE86ZfO2bREmyz1BzRskX8z
AwLB0RTXY/8mjHNmcQNF6+b+1ZjvzxWlEAORYBngfksWaM8YPSUiegm6Px2YQ7Kvxa32L8D5uEz+
x286ydWXAZ38uQxbwOG3a5VsIhjtm1gtShd8nK9RAYeRPlzrR08QGoIgmrniDAq8SulRvDI4sR13
+0DKkd2Q/FeGpJTxPX4Eh0D6J3gyUqpCJ7oGPXQL0mqvKFjNUNIPAUNqjtjGkhgD95RQOI7oQHdP
FNL9WXDk/hB4Ado+7e40/3f96GlodpKN6OQqrMCOb2g1Lg1vlJ1AmSpz8cR9eo0qm8t7IIEDYUZ2
LuLzQJ8JULWMU8trnv6WwGZUqnzfnhar5EmnugSbQzn20MldcGWpq83YCH2MiI38NmAPUSkr5Zat
ydTktwZO7UKCb7GWYxhiDWFwkQEuujnGQeClF8WpO8ZEQFcv0+lcDKV7EUeJGKJg1di1iioU3fdH
wUVO0fwyEaJiLcOXyxtwJLqQrXqijK0+uadZ0vfuzpwOJGoZ4U/YMFW5QtVt8f+vzF6kbzBGHVjm
sffHgcTKEL/f/r6LsAsxIRUQ7FxzNYy1S40Nqqc6iuk/aeeYhCxD3I6XMDelxjJG8PjGL9tlgBZR
oMQ+65Xwf4g5EjOp2x+qBNHUTPrwXgLQ5l/s5g1cN1qJgPnokZuW2kwYNnTlFPvBtAQbHvIlQCsH
ogrqrIej5yFJf+jy68XAOL7HtNgO0Ut7gm9yCVoiROL83RQMYtnfzmGxKDdfUsk73O43mom8ZyTD
PO10/mSqqlgZFYxl3FrAWdbAMq43UKY/uoD5MGWkKGymVY3ZqLRjZISzqJjx8ljLpoLWLkCnrSvp
nmc2gqd2/fxinxTAd+uSHbLifXyYNhP0maZR29fdpZYd/ZQ97UlArDzWjZTlT4NBjP95LvE+X427
1oMLlqfwbd6DhsQw1W3rHXhhwDCgFtFfrZHb7Ad9L7FM+E2fPwD3tgv5pDpZMrMhqQDPGFIV27YN
sdADoHwGAYNAmh2gNp/ap98iWuyjgmHL5J/HDcmMIWjmvFU8JnQVp3t49kihSt/aeOVtcGJI36F3
YzyBrjchCpkTfoAfZIC8qpZcR3Yd5ddDd2rD2hxbojMj2YtoZjxGE7vcSwffSbprgzIMGkFIlOsp
ZQ6SDxOs+ei8yOpFzq+bR1b5yqoeUCLJQKNzVWsDksdFrDCSwztk7UkosjgGR9qwQKtg+ceHDgPc
F8cYej/3zt4UDz3um4+CNjaX6vngqQMnbThPO8IT4uMGYP7+1Kt5Szs9pNsZ5TwTDWupfKlo89r3
3ItWYfXQxUlpeE8m91Zfo9wULk0NDol3/3ycs/AnTCJ5bKvT8iYt/nwUXINlYAVUC4kG3huf3Jn9
tNMv0fyBK4b8TVpHdorUqy7QB7o5tIlL1W7OBVCFwoaE5BnVZfll8nQXaMk/fDSZsSV6D+7zaCzx
PbhtMms7Z+BHXJ/2/V2gF9uGwCp9Hks0raE8H1zbyfoVT00PRGfIOOJNfRCeqFXvfggLyp/zQlZ0
iBZbFgkwH3xPEWm/HzgwXGVDLb405FjZ9KXcxjMtCaMIjQh5XxKfmgwVK6hmhwRmVI7m1Ofteiv6
NIBBf1jWrY/o8+4QZ6PvTemFvbcuKLrEqAI+YiH0dF273lVnTe4YF7a/PNpksqAIaoZwR7d/L6Fh
Pxa0Ro6VBH3GOxA6MOg2INv9Bf1KV34nPv4J69G0xFv27yuyjiSswIOdejKzMh4bNVZ7rVKKt3am
SI8kfBoe8g5fWzlFMxYNpjM/dClfGgm1MRzmUWsjzVKRlnsiEnkjmgB8bycAPpMDJhPZtuXDCuHO
y96MlajypB/iHFM3vsk6RSrLz17RJoZHE05Tpn+ASrB/K8cKpsF7+ZNRVXgQQH0XvhD34euZ19s/
M/ETfV0nrVZXAqP8eQvFkdCAFJejNFKLkWtHaVMLEz6QpCbzpzeHGqkE+pfs1BgGMG5JLK61cmPJ
3xvxEZaCg3OjwSPEK7NpQBT88SAXJYD0nRQ1SROjmwKrWLy7sI3LTIJ0UkyY2G1vRVWZ5LjIN7BX
s6kU34jXWjqjsQscH9ES0DWt+2EZfPH2OhsEau9neta/7hUj2/G5rvgIP6PA6FsFZtOv72XClwXT
R18iYxnezmJAqsdXGBGszxuLeGttPPKhF2IMcuIF3tzDjXA8tVQmDung7iXbnog1ArnwTpVH20FP
Y0VRwhXl6P2EibUyfBgIzUAOcupWPxLWIgXUuMAx53OUofWQC6Zd8VHU/qiqCGNR+lhSK7bAgx5s
lab+XJMRT8wxIGSYesnDfVeK23JtD1LNHemET1JkxK2QQlQsD/Sw+tX/moFyhQ9qUDx7Ae1Mrptl
eQfXhaCcTzyiyQs1OTLIJ5btmzdk8kDiEOiVDIf6QJCo7iNcKb9gU5R81s0AM9RK5S/UtYte1KG6
pA8Y8SavcBHif7qtQys13sQ3Tzb/Gkw+dvdFflTW2og01DNvpQm9BCuxPgqSmUlfU9dUaEhDSU2V
o591wjLvYjSJVg8Lal0qZ82Mip7ZVbbD6o037x/YDPpUEK9yrSa6h88RGj1ZFHfT9j5RJESzVh3H
YwmOCrP/2ViJJAP84AMLON0oHJvDijPxOlNRk3jo5vX16aD4gCdXP0WSRLMdITtYhC7qWvGIZe6C
3jAkvnigL855CfSNxIiPNgfTrd8AGsSeraEXpWXQzQgo2oAof4+NGgLrYj5XO+8UNRwdR0VnNFIG
RVm4kf2xD+SGwJxH4dxLBhBdQILo8MNzxpIXhsEoxDoC4HG4VbI7OQ+3r4dRdrt/Fq9ICgW3uO44
OYFST85ObN/4RVH/WCxvxehtWoKLOUDdBJ+WDMlaQ+0ew1BdanTpQ30XZLXUq6KZespThHtyJURP
UxvoGnJnk/AXHuhKeKsF5xgX6kONhk2kMHOj8LTKiOFQCZIBdhrtgXm1/TdSHFgB05/bxJzkPO6l
IJXnTFnmSprPqVAa1xRT507ihRM8fVL3aNV4iHmt4j0o/Lc48rX2zkKx2/QSyPEF73S9n0H/J+rA
Q/vUYlW2n6+mSs4PY5jk1wvdzuSM9gbAKus1IEwhQejiVZINVbN8u+XycZBFzu24zY+toSVyzSNh
GaDtndka4OPDz2OGVcpAJuIy8MkzwA4bIDABGYXwuruiZL2IjTHoPBZ2yZli+A3G5VSdngPjmE4Q
h7z3s6BtdYnwXkLP3yUBNF2ukWMhKozPmjQpSBRzx0SRO/lWEGtolg925BR/kS2MmKhOCPqX+Bv+
binLI12oAYVa8/autwv98S0NuPzug8uEZpv6XMZzpZDumOp3JOLgVDDh6rXCmhdsxTsr4AMkURK5
PSButEAWnVxsyILm3QkCsoY9+PGiBgjS8mq1MsButxD2SwmDaxDgU4t6BnZw8V87geavdrPGfc7C
dhexM4E5EZb2K2N7zfWF+3WYCeN/IUzOAFbOlO8tRSusVEYIVvklsdaoghRebbYLjpGD3fNqFPM/
MuGpjSKkeaPVsSmveEiu0vnfTn3pdlW0Ddg7F1oZOCyKXIiBQUVZJWVOyDYwDZDh0lMh7jSdFde0
NVtD525bwxgnHHFwFUQmWvIcwESevM8rV9Uqb3MKkBgedt2JqAhjWtxBIe8JpQi0YMF78OHU7Tm2
z5aavrm+YwliBI7R7mSHks1eMOdTnrkiT+IkBgfBZLyaUh6F8PC26yolu7MKMZ10M9XMxplwB9qd
8zK4dvYnpaKm5LwQjvhGRI4frau/JK0XpEXdLuY3/QMuC6seySAL9w9KpxRxh5sgvj1xskXdTSkq
tSjO1RWZpY8M2ctZImnK1YUTHPDRlFfwSp0/dclVmDWq+oUdI70jjAMlIp/ZoTr2lVYqkCdIGIqO
kPfYPDOMBNiU+X2xQn3xRF8D5/DUAz8bmlM/EVHN2OyNGFXL6CiTeWYftcBq1Ze81wRnjlUd+Qf/
Wdh9Cnk9H/cgrMG5EPIB4TAO9fazUz4r8mASxC3jrWsmiR0qmj1IDvI5YNabmJQ86xBNe63oX3H7
QN/lBxT2emONdtrKAB0hJXTiUUWc+Bhod+l9ZsnE8Gva3cYKgiBt1hoePHH7SN0Vm+v5BvWCt6aw
sNhPeLXNVJPi86KXJ85gUD5vTvWmXjPULuFx637UcqzmuUIo/dPoLa0NbG1JzUb0DzzUczSNpKxo
soPCiD/Za1F23P0AnrC1FwYzKJmQ6lrNWCS9NRwrVH2t50eXO3z8UDaXnAvZ3JruqjFE+66lpfVd
fcHGf3VEFZ33EIHdoTfG1hcQuwKTidb/4/St3n3Bt9EGtmh/beJ97AQv3OZATjRP7dzn2N/X8nwb
/3eUU3bRT3B4Q4W4BPDveF+dzuT62qlCjhUhdp2vi0sqo8y5crJcv+y9bLQxlmD/cUldtULVF/rq
bRBsk29shECOKKotKcrSF5dRjbqlIjrQNh2cyGAl8i4CIEINI0u4F45sFlMlRjm7TdMTIahydISG
DifIdZdzFNE4bDe8Jc6WgTYFkA6hE5OUn2BnweiTj2CH+Gx+P6fFlCGqoRy2q1VLj/G+OZ7yeSml
OSbzO9wdFQ2Xw52Lg/6Ou9saLGxzmlFJIuO5sfMgjVz2GjlqitW1Tota780VTdS0PFxUdrV55cFS
mMPAq/b3L7H8XV58j1+CU1cnHb0Wqtbr5tHtrlNMnzIZTrxgslWhJLNribsI24XuE9JjO8oADjCd
2Av798WpCPJA9Q6tGFR9WaUDeG0YQX4gbqvcMir5DV5VGTT19hI0R/GQ4mfpZf5OSHEt3VrFEExd
CZkLmzWy4983c8JC0JVe+CxX5Ru3QOc0HrA8/Jael3UTPbr1t2JLu7jVqABtA1VuhXL2XMQH+Tkg
yGDqkDVSnmjHXOx+8wxeOIIo9VGJnJKg3oe0CiA8TuRgzBVUi4Fo8iHUYAJh+dMwHZxltEO7y99v
n8pXVIQ2pPBpoN+xavSQyjb59uxhZzLxc7HC0tpp20/L8Cbs6GD5hRjP3TrTapLLWH4CXzIOfwtf
48B+0LwMn6AmTatMuvbowDXifOAXUekZKJ6GTlsbRoBaNX50opI5G19yMleiiHhigPWSL8tm6EMy
xrVPzFQm7wPiXWkAmcM1JBLcQdqcKYIotV9dFULhF/75dJBtor+R6g6yDDBNhPR4jWLQ8rV9m8L6
GVfdILSXicvREc4TqoKD3sj14i2FPKv+lOGotij+TcSt/tZU3JNdsP6++d+91sJtEzRvvOSxy5l7
mk39Jh6K5owXJ8z3dK92p22VHJTRYhUb1c//OiC47KBu/AnJ4yrTB7tV+c/o1swACMCPLm1BHKdk
qvUBxVZEIVpIitaVOtAoZ6lxt6pNmphKWzcyZN57V4NJuHbKx4onS8RKiNHLNTRJgPII9UtQpH/5
iQPn67AOC3y1giuGcgKgM1amftROOS1WsLwo16MtST1tUNWdX3Td+1bnL8biafFD7gi/w5BEiVb4
MDaoTzlAWfG230qSPP6G18lmcrQG8/f7MjyMqMyKKFgQHft+uGcx/tcypEwKPql8DGXfbJTha9v6
01PFfzvVqAE3Z7Nk7Um5bjM5Bv2Y9lVTp6OeNF7pTN2eCKaE4lbWoA4yW/b50f6ctvt+SgJDQlLA
XpSnQlWYMqaH4xfHldvG00ERYHzIywDSqIU9geyUj8BrU56FPbKBXF6KkXt1LU2GibjvK0i+7J7f
joGZHtXQM7hxBM+JZFNtBoM95YaHHLz7ca6t+8nRn/D8F5SwXZM6kZ3wA3skY6RDtbkM6kjXNuZb
cfewGDtEQ2cRiuGz3jEdbgJD8kFU4bvgQmnPEsn7vNCTLS9wVZqNwLoTWb02uvlVcDLLOF6W9cUt
8RjJmKkIylMYA8SqdW4jVJTAUaX+TxB0xyWzoz1P//pWRtH6N5ajbrhXxSOwa2hAO2foYRK8FIwP
B039rtfB+aA5HmYYGKzpLTraRMk0hGE4bHis2SDpTy4rOHPSt8c8teWi+RZTt2sKc4gkOIen7D/0
0bD4Ir5VHdqFLwvmQutqznzfL62/9OxKOoDIjEH8D6PmdY4HAbxASNU9lRqGP3GkplaIo/srLtem
bK5kLCu0u8PYKLsGlSBgtnK6ZYjM3mp9iyOu4z6mUv/JSn5DnZcBrwm4kBBA9hSRFshaCpFkB1Ce
njx5T5F5uBwzOUKk3lnaRxshX38xDNweyOYi+DwMdvJPrvUjc7Bslgw7S+DFOuWsIu7q5Zx/Yuyz
Bf5fsJq8q5kx541XdGDy+ChXoj+7s4Dirv5g3w1qCRU29piQ4BHxDkqHKwyCQ/elQXMIjKlU2DoO
YJTAxbqxlCUwJ5MGjUdHX+WhhuO6DCXx6ILK/0wQv127BgGJyOFL7d5MDemd4PQe6xdZjZ46gYmw
2a8+npjzvT6spk48XkMMVEwKdAebQ7wm5bLrmqqsTpnidSouPTDip7rXBQ7pPc9rSW56WW3GNk3T
8Tbb9kcoiWDWfCdIoBA4A5P33rf/iAOMW9ZqCXQ75NVbYpTImHrRFTs2IahR9Q7Fh70tTu/vWmpX
iHzEXJrxxMtXrjCxRzSEDGIh/UKlFbumX/uqjmthgSEnpbLSAFZMK+KBqYcR6sSjYQ9BJuKBeQiA
35oKOiZPD1tZxm35UcXE53hFwdrtu+4Od5Rw2JadANIrobW0yDtsWDKulhylbmLuPNYM8naBlQ7/
MYdG4Wys3S3GsNqlYQ76Gmd7kG6wYNDmvdKjzbpabCh5Ybo+2z0OS6EBC59a+XY9M7UQpPqebq7u
d7SooZcjUpHrn3cFNkHG/vw8zok8t+U7l4IxAXFa29LclrGy0yM6lMBffxqZ3SZuhLCoYg2MJXfT
SB6oUFphoI3UIH4sLUdmr8K05ScRXbxB8Nz3yZll5kvERuVvqJg3YaC9uADzWsynW0qtjtP3eSol
6scUIzL5wDUOllV2ZwA1XbqzLOUhS9r8+EEaAioy5DmLhJaxO6EgEYuc+uSR9zefCZJW6LxzSmi6
qgMZrFnrKPe8RjnwT+6qzJ1bnE2MoLbExKdezPeEqRbBgDV1PbvRf9GlGmIA61kAof0RkRlVp816
tyKtkbEQnoJVG/BlvOrz+rW6y+tIp7c6HGLjdlpSL6tvWEnK0+/WHqg0n5eeFQIOUqk/eMjse0A9
WEw7tAGY2K4hBkNBSS/J4TU4tjQknLplidbpuYpnNEEK0kJGKtFdZ/r4JPQKnwF65mIJAYebfxZn
K1jxmGvxb5MZAV5Ecw9TJDayAumyQwNLcota2bT5BsX8aOi8cTcFZiz7h6VWDifxwXvSNr64elhr
taG2wrX+etGzkNDEg1QgPsk8/BwdQXIzoKV6UV9vqF47Yih3dN0Fld7hRgnoaM+tguw+x73m/MCX
KfrWZ4S+8CyHJL6XyS3Azqky07i+XwcvEAYS9WjvHL2ildTqnFrvGb9aGhv2BGYPdNjB6Y0IjDvQ
ZWYeV78AnHOAOn/qA74TigOhBNIgx5qWbTVCUUB918zvwEva2txPVSTsaxDaeJGHu9E68aUZfzf+
sLA4zkolTHZ9c6Ah4tovoDo1Z6psnsQKnEhi3XEIaC98e8+W01jzI1I/1gNnkbii/b598Nxl9sGW
wH1LzdR1qcpfd9upq0jyOnjcJO/G+u0H1y7VOKZNby4SpZiadM5Slyr76I7NFXkAjmB5zrKamt2o
DXR/0j6jg8ftWytSgCIuJcA9MVK0eIoGG7JK+U/VqUoSN+OvrR5ync84zaj+MIDXxsSCSeLLaCF8
0folz+7YwzLJHFgE8qYmpdL0C8UlUT2ijl4Iot56Tr35ObxV4NbaI3jPidjG+9ZITlw0kg4k57Er
2sUK5c9hYyuVoD9k9W2CD8RKqnBiAAgZg4IPeEe3O6xPScbknQbGmyvCGdU+SsrhFK+B+lOzoWto
CxBaEWcqG3FeVui9Kfcakq+RpJS1vgdK77Pxw26Y4akZj4Nq6DbVQNiJgn6VL6SJfVFmqmaHo+gp
czMRmg7ctMM1k8/4wUHNGHodprKpfNdM507K/45bEVNsUL4Q/zP1qOgSizgoApZInb8p79AFR9Wr
xpUX5R1Dp+lKB0yTdkv1jYERCKo3pkzjBjiV3DsY6vup9h6c44bDkf4kyE0Zvguhyw3WUQaxuYEJ
LNjxWewQ5yaAiOuWm5X4gAkMrEZBit0GYHWUfn0Ly0wafXvrnOEVEHtAUVHaD5WCAQWBN4PwPH5G
TGTnKgYFrj9pZKzP1aQQ9cJLBHkuPws5atTeVob+5BkRxt+6p8X4EZfEg1VgLDrV3SyyGjsgOmng
DD95jfwtq9wwd+aFFWkwem3f0bgXmVh9fuHQXN+ggmLUQeZmnm3TJACdUJRt6l+SzdRpDCrAbXYH
4FeOv987fgHbR7ttf2v9fwDmHOUThRJzy+0AfCoQFYWn46Dk39AMUXEpnh7o2EbGtmGnEU1nWY/f
1bU9YV7Bm9SCwfCGeHtf1qfCiPJCM/qhM8TsT2V1fDj/GA7i5w7MoFyq5r8S3IeVt0hXl5SRqHZt
Yq2MQO8l8pVpEw5AAUsqqg2XHwB8bPnhfXBS/C+87v/jmjfpzhIh6BSACesmR53FCpkuXzO3mNSX
P1tJO4XQBnKTBGWcwjI+j637wrhXA5byEViCf3zmeWwioEIlOELv7/vsjrGAQ0InCm4Ki0RkBruZ
ilbkHZ8hL66jRcUrFkUc62rYgl0LPNoVWxRNjPGoSCFbGO7NfuBkvrYPWgyZg6eXX1qbSeUkYkZp
8Vt85QlZwPd3tWsUbUId5/cif0m42k45G1MO3UZKR/BAAoh3em7ex/9bdf4Wj4vIKQn2JkwM29nm
X8w3uh6KyQw2wSNaL0REx4OTUCh+d9RW/mlZ6QzLP2//wQDky0OVQuiQdoEnPZkvdfy6xscZodlY
xwijPZUtj+kQqPZFBuNcRTPz8S4M2TsuPXp5TWyW08pgSrUZPOmFXVHY1OFTwpC8Z5SJV1zt0EbC
7l9jvPl0X6zykjgGTQcSNiTmDnN4q5f2o0sXvFZ3x/Qi4d7xHWO59P3FufI5ZJRoO+8DcrqQxvFa
HgNMlNxFCkTHhi8V/m/Ha80xFH9nWBJcjde2wI+f3uVRDFvxyyRahnW2J/ln+Ctb64BDfyVkcmxO
J76Th1fDW54FNJhJlaezSlV3QdchukCGTAfKiAWmkbldunkCkFuTsCuJtOhg3p3Vx1VUHsUtQeEh
ZhqsmZUzhYCNJ6CcYfNkFDBai93nbGnov/SjGmPAokFFo443u/mOmQqKnXyX/vYVRZMLOq8kdSJ5
IHl/K+LHUmKKaRLs9g0gcSG0YnPfbsXWX3ep5cH7McHVrSFzgm72n0qydqchzY7D8zskUaExI7Oc
hlIsxNID9s8ZFr1t23MXiqYCXf7/3KUJb9xJAMINFbLEYxGKG/yk1QlprCD5CFrNm42TQ3Ms0MF5
mXLKtWY7kD+cqZOvx99w/dWTM8d/5O1O+2MsGRwOZsg9ZzP3th0c/krDwl5hlC8l69i2VCkJeVGj
9B9o36aer1QGFBOSgUnKcMfSPDK1PgeAzjRPkPqNDUHdYyb2XptZJN+d2O9Q4EuEDsG7ldfch30R
dcMBLjXPEL4+mb0EG8tNAcNjdjpx12OniDMlyVAijltcuzOF1E/osET8zYTP7uDQcjvKUbNDVceN
MCQdbwIfgd8U++XTdR8mbZ378FzKF1x5zaEoLZQW86P8UsN8xJGOvJHP3PnJjNkq7x9YSVas2YgP
4p6cG9Fqn76lAvDtRooikci4CuidnOqC7wNIGIFLDAneQXmrYZkvAcPb6p7ptNkv+DVlwCmXh09n
g2jFMyKehgdRl9FdydOlpOziaQepKt521xFZCVPmiyhNCPNsjH2H0Llo4SzfvG/v3992OiceJSYv
hBDDI2jKMhL/ciIXARtgCPxhPTgeos2BLmzXMyhAQSphvViNngPsjWfdlL1A71fSKyJ1oa+NPgau
u4QBMqjJRmphgH+oUsKWS0DKtJ1ix1tQ6oWZ0R5Da+66xQiEfKLF5Jpqq9gjTfleRnKLBtKgxC65
7IC2EqVikR0OnGlOVBQRbEC5DAPEga0FvYWPUVQkxZhY9ga9KMz6opJLanfTn2ahMy2DkhJVSnjX
6wMK2Rfn0HiojF6G1A1kkul0iNS4tsGaA1A6kBMdCpLT6RiT1ywQ3uMcu+RAp986xqqo42R8iOPJ
MHrxOQSuveqK1Yyex4b300iWTYwIzfHh4b8ulY3XigVM17Qk8aPCjzKluzch0QYPlBozQAxE4AuE
WsxfudZATkNqZ5iQlbnXEgPRrrdl8fTbtoH0B5h6GQef3HwP2xqvx8/3j9aBjTQ3USrptM2UgMxM
7p6U2326Bk5uAksdAJUHjX8z1dvr966d2V0CbRCMsXKcITdwMUvG05t9NMK/FMLFzNjf5njdBUS5
zK+VVAobx3TSkN+9tkBO3WKYCTouNmL9O8MKSWJKm2s1PxxgOd6uebVWehLm7wwVcYSJAA6y8UBe
xRToEEFykWz1nSOLyfgSC2sdsYkcx9mPl7BEze41RBz/vB5mw+C8VrilJC7vJISHoRW4MbgSWsjO
8YkAzO3TuwVlJsCApAigr2vEkwryZPxtI7Kp0nWOtaseUjZ7JKC06NVIn41XfanO29vhB4NPyaiK
XBrnt1IRsr3qAwpazdGmhTbESZacDT/SybBtA5LQnPNP1h8gZzFYfLYooxsqM71Y24dgOybastMm
SsYCZntPSusObrP7EikTt2ANPjQ0Ofvq+TGr/mnnpAmxCyLZwDwhUDAJRoxn7PzL07F41MObOpLU
qpGTYjfRzDtIkEhBiU766/rBsu6I0VjqHIylTyvmsehElH4mGzlIWn7e1hWWXUQ49BqimyDrPhTD
/rs4G09E6f5OzikfdGyjiN8kT0FURurrCOZ3mdn9wno2uK7eOYWIAV0rllp/J9ErZRbPTY0BlKOD
vIkeCe4WbpNGl2vRbHZmc778VHIrx7B7msBY9kaW49Cp4V1+RtD7eIXI6IVfUHKnrGw3ikKi6WSl
RBpWLuIshuJl3nrMadvrEiIFYN0U5wyZWEzLmN/kS1w8nRA3lSW8GD4M7zsNrT8WRSkwZX4zp3/D
/wdP4A6csFSkjahhJzbyVi6MzLhtCXshtPcUq5YBtIAoCRYAEgd4+OHsmovTk1HL4fMHQidWS/+e
tjoYcL4/YKtEThoVjceIOeUzpF3X6Vl6JOzQ4GMxqUj/0xh6O1p/Ik1nfINdtODsDJVShrseam2E
8YL49P+Q5ttFkPlq3dH2gySIhOJfbL5VdAEZ4oYwOJS/jSzQYnIQFXi2yznEYmifuPW8WH8B9YUF
rd4lPTgieTa73BQg+DI99rjpTv8J3LwkRcRQBbmBagXlYa0hIy7zDPaQtge2WEQ8PBePQ4FQTXnw
M6iSwDPraSPU+hY4+GPuBD9bEOQzgh2tawQrVx6mZrr6Vskxakqyz/s+O7JhmNQaI8Q1WXYDKcZM
3S3Ays49jdYFVFaUkibnqXj+SAStP/MQ8c9DIeR1nNFhMUWUXkbBWIWrJNIh2xcaJYoVPs5W22rn
lpfylaTxMrC5w6B3M/9EJiqelkKzrFzuxEWpjvQJ4uWe4FfnjZ2Pa7IXEt5dhTkB0hhRJ/hl+rE5
VIV6t43BxyyTLHKNUoOdHZSQXxQ2qEP193lMAlNAxl6WDvzUza8z6L1m1TpWIlXdf27Q2xqJbL2L
cA9VQwLwySO2bNfe1Ka1i2g3ryru7cqlwNMslXKXJ+5MEbw0xnJ62nb6mOn3TyZXEA5UlXtoHRAp
BWrHhFdJq3vMWep66wub4hSaH/62S0GB4QqwJ0739zzde9Y7SvlnYu6FdxFVF6It64Wvn8Zo4wlT
U/NfZ3zbNRn/xdHFsciqRmgD8gp3qqngYazlaha7wA5TIzawUw0rvIx1g/8dyuIWQIAUgP4jyJZa
iiAs2dt1KGM6g1JDLntCzqwO8/Pn8C4nTX5knKVK+BHPangG1alKgnif9IDWqu7CqMNfhzkZ8pc2
3a6p+btUHE5GMNcNMH9l5MmUMUrEig5CszGs7U0a2OdzdGXCmb4R1QPTFoUyrtHBHDyw1bfz93Q6
I0UrPsjlmYIhp9vSQ7dQCA5oGGOlY91W3GsBE6/Sl6+olUf/BpfGcD5OcPQtdKQtcULrvLUbl0Ey
LaVHWYdjAReW7aFWKgda4a+ZL3cENGYP/G+3ZQ+pVeYJfzy8sY3FV9TVpg0vG+VWdEgBmDvhVd2u
9MMKkCpzR3NfZxefSOcCYqrMSZ6c40lmRwXgHzTPdobOAK1ths3v6eJFAVvgBWtPzRP/ilN2b0dR
q32sMS5Zkekgst5o8thjJOHxDbm2K07liHffwbfVhCMhENjdoT1dD3+hHr451STbsasElG9ATviB
KqrUMZGE16ksDWOt05IYlWJBnz817CROd9bFtsG6d2WyGyt6/tmQ4tGldcXQ8akzFw9f6Wpe4SvX
R+SV5QI6k57k79r7HB005HF9AYqLJQhrLPxHs9BiNBNnnZQ6rVYEQj3hnFuJjIWYmo1qGiJ2ITU4
OwBJAMTWldpfl5yss2Jq3pKpVgZvj3wo2cUicysmNE9pQnZ6SMyy0F90YJsk5fcxpjcTxkibjdk9
IANs5qohM3lNoBflgl1Z3dmYJ51fPUNMX/GPNBLnnN4r0VvjId6S6oAjQbbl67UUjTknzOLt6yg9
NsAf1km2kUE9nbjU0Ku6VqCDpSwSUeSVFTnu46ulISp1EmEZQNLVFS85dPF9WCcWiL6uTxj9xu43
1i9UQGnrJWdtEF324an2Avh5Gp7kOil1SRBJrX9eNuwxE39yx0Owp6QOKnZTx8pykzQpmWxpt8Q0
qquaMh1tuC3oivHSdjmxrlkb37i6O9Sy0iD3NPnkIBrdMuWzyZcfk4exoZIL1iX/VGqna95HbRZH
IdwOpWuLMfl8puVPyaxcjq6uab0YnvBu0LSX3xg2PBntF5BvgCXnoK0dzsoFGsHp0m0BlTd7trYT
5EYLLyH16O+bpJcMMYoIJU6mNN5IOydQ4I8tHRaNMUTKIP7iBBm6QIFE8IGDxRTLnoLXW7CZ7aS+
B2hRgW6VVhazIdYGR41DKfoHD68vtHR7KayFzTMVN1MDG9lxXfMSWwMXa8Glp1KjeRqGbnSYHlpA
tQq/dpoZXY17jBKHuLPTPKh8urjfUNuc8Jv7WwUf1U0JxQdRvKUe7Y7ut+fO1G3yR4EIcykzTAaS
w9ErArajaBVGHr4ji4Hvd7C1sdX76+SVbu+0hNfhbHXEED+q6mm6N5QVK4WVELbTictxPJnBS4Jn
ukVkoEPTEZznmKzdXeg4GunQpvXPFjvRBIh1bh896ktnKnoROGa0ZphQyZpGYkceHfuMAbipuiM2
klSM7Dvz2eAFjzzkTdo9Q50YgC7/Ne5MhHcQTxC1ahhEh4OVpYf3Z0q4It3jbpkkKYPh+mivxGb8
ICk/DSow7xsCrLEgaSZaTVhD71CPsQxei5UeNtecqHs4tvw52hv0FmV/D4CTBKSo9V0tdBWnUd6g
SKIGN/zzYS8JOh/A4GFNLJ2Ho8tKoF/5KRsW7cTtiuS+P6xTI3thTJT0y6o/dkB75qyEz33D+Na0
blMbNNai2zhUauYaBjuTakHkcf3HMipg3HwMNSF8Wl+Y/vUb56iwtSXbxc2+bEL/ekZH9Zbzd72z
RylxGsLX4+/aAbg5X77emQXF1ccoVxyLuYWfVCS8HjGrpHbafJsMogC+LVyK1uJqyfcmT4jvO7Hz
yxv3ihJvxEKP+1K7SevR3TjXX1mxoqHbUyVw87UJH7fOaBi3jU1gnXT5oj32ZVTR+jj5EFjZw1Xe
X/jkkJ4HqWqf8I0ZlsU6WEslcnZ0YaSFV05Gdp3MlnIAkWo74kkyuMV7j7yD57ab7qs5irZ058qM
ie6F2nGpUW8heQXNA66ehQFHNW7dG7B7BMtle7/gzOb4oWZnpQWzv6FUwk1BKTS7OYlVOsV1B/MT
MRboQIqcWuMdYTneH2i3CqxMhOhS4I6KZ9aOB+oSCE3gyfVL8mBrlPTxbcdJsJIQOJdPjbaQli3H
SqnvGQTGQG3sjX4j+k4lz6O8FvF+u85Xj5aOsIrK+MLt8amfnnKyaQWlciQwltedR2sBGx+siLqF
q2Wh6pi6JfCgshkNbGl0fa1MWqiQcr7bb9N5o9YXwapspox/4mwNlphO5tLuvJhn72rMyAh9OfTj
brbauL7rGrVdZQiuak42B5seBfIHSPgYnYcOiDYAWI+QgdbOBjXBPoJRqlCwfG1B1NWvzuSe7ZSE
QehPAITrBIoe2XlWNBm/vH+7eztDrGbCAKFZvSptgK51LwRdRYS0X6feE13TIHFBnFkYpYegDI1x
Mi05TPAowBhi2W72hda4s6urXkGi0E4wLwO5xpAaRE1ZC5wZGgTfAQbLd7kK2MAouZgZH/Xydj/g
TTua9VcFgHg2k2UaAf08UA9jHtYHCHBsPlng/RuuTHt971qSH5vA5deqTo4jE1eKNbUORqaqnTiO
pRhslFzjFOTl/mpZjB7I+SZa9+wCyd4l6gUIQOT6E1403eJ1XovQRxz9C4ZAE+o07I/wx6Z+KB13
2ndKVh9WQjoao6YoRuzyRAY9nxXkpBaBYpTXPrxVkqeAAxhvSpN30bKNTLukxZIL3LzTJTQmLEOY
uhwIfMDhsvSdCKPOg11gDj6DFMWmToEW+PA9Fm9KuE/KyBb2lIIOaJ0aBWdu3bpydU1syovjpny7
yyw70sWsBNNYZf9JY1DeGzdo3twPz0jTbbjx6OBlQltZVQu/TNbrcG71xSTgDSFqZqJ+7NIoemt0
S3NohlFTC93JBB36i3O/0O0nIfJ1IaKzWoHysaoNVvJTtpZf797ECWwZzHADyDyhukgtvYFHgpKd
D6Bztp8CFQmPs63VflrWzeySCncRHYws3xrENoe6DHDZUQYXy0VG1LlBWnrCupBKB0GrTuf8ct9/
li3u1eyrMR8MFJdppggbaqzDXBIRTplPc0c3JMN+XR2JEWJFS0ueY8zHn40ql+A/3sm+DToYkafq
QdtlBFTdf0LmEQfWBT32WH1eGhOd6kQiFXCg4pfN8dADEg4dsHQEz7g9t/1xNzZjfzbE1uyNcTBZ
SQMkbqzPvvkgt2sf0fY2j1mGhYr8OO05Ya+WloiesjLFrIG5oePiNb+fmU2BtHp9PQrydWsBoVfc
la9ZeeC5dHukb2DV5dQ5y/icVjqrZPAgTPwKWJKwAFPMOPYXsGwHVEvJPi6G9SjmbV+T6ucYXOx1
Ce46tLIhgJNnCTHVpnGEMAHD44uDXSl2nRdBOyWWobKHXh2tZ9NUed9WJvbO6N28OZTHBUT3fF5M
EQpX9dED5nsDUQH43zbAHtcfyW/mzT2qvLvV8YyP+0iMKKG4auYyHBB1xJEkoT9wz18sHjgJfn4w
xk34HetpbMkcnFPay3lLmQywASUdC27J/M4plP8CFO6EdzaUHpoMpMUkiEdRRJymatxsyNLM4ua3
16dJDWTuUfyrKbHttAtk+KwQiVQcNomDXdBWQ1qoYRAqLix3CKZ5lo3EFb1eYP1Km/sWq5/TKW2c
UFc7Qw9Oc5w8pBvAepKXV5NWXwNGk3eLhRzHU2HAbOov9n/Iy8xvpY7HAYUl9IyMrTJzKvybQ3g3
ROzTXvRXH3Di4qTISGPF/VDWElHIQ2X7HJ9GB04m+1QZgEWYBXHT6x2rG/RxUMhbEwIwJVrPaPCx
fkRDaKWyvqetNga2P+aU5HXpfl/bnVYVaBDCbCREfM5LcNOHpOgpOBHRjjoLsdZuRBnVAqBbipN6
U39EEJS9uF5f7XbL7lJC43Ib1pkoKzyQxCEvc6C9bXF06mNU9nwoRQc1noIf+3qcC37qlkM3yxoh
DxUPo15wKAHZxKLf1zixxMjjjnkx87REdgbZO9YYAH16CN8NRRkJrFRd+r7ogHP8N2KjFsz46S3W
rcBXTYLp4WR2V/zZwpUMk2bToTpVEnjm6JOBbh+/W2bT/+aLUupHvm+Z2WpTl3Bnls7PqyWfToPa
2ansTbqBa4BnIqL7ykL0MYMqSHXO8Br7ROgeaEypeXvMHVv74X/yofMprxOUuSadTUTacUzD+V40
91POXKwUMp+L++hauBcuF61bWoWlUiFtyAlUcRyXmL5phr08IUhWyMfRdhr9o7G1isPlm8R4MjVj
TRripDY+eH1K/+cV502DxjLq/rrOPHxGEMxZMiEPuRcIHzgDq5Y1XH30RPOyLpuslfEkAmyG4XZp
zboiCmCBe6+oPvv32y9hyGIZihyVLQ7RJ9PSElmUQ+loo/JQKqamqCXnBx2Adlb3iF3nHkvwH6gj
UMmkDvl+JrOsF4AXFGU+baa3DXBHfn5avaAbSNxSVXjnFVixCOP9Ac/ajVCASWs2FV6CeDgTR550
TkUPpEIFXASzU/LNTVYwXdQErzZodJIY2K5j8faJNVDG2HLuGez+tQhMEzg7ekno3vpCJVFvMaKK
OZ2cvZlxpk17x1m0cHIoZRmnDav0wYQ1sTuNRG+uk0IMNTeoL+7a5SvoiulgAX5Aa2VuGMw7IYVU
OdDwNbVZ2KJJfsS8/ClqH678F5W1PD/dC0JyZrPLzmqWjNL0eiWKul+nWlEBaYLmYvSt10PkWviw
OYRmS5JbLaOJlEYYIswvduPIHO8CMvsn62AJlY++oL2PEnoDbVuSE6xaCqxLvjYcD9S9aizWfd5i
xSjEAT5IGIlIO0zZvDHQsJ+sIxfZDP2WAcBieWCITPO+SraeuHKgl6urPj5XkziJtAFd0IJ9Cwuf
F5O+tVJSdBvxGIAZ0WQNgcaaPdyZyrxucly0OYmdj8nYWK+wThqCGOwZpSefLLJEScwdaeANIwCW
CUbhbSlrPbsDQ+v1nw9scuQEwgxys8lfl0OiV0qwNHvebs5vt737J7Bed8GmvOLmlD1nInFW+xHK
WNrnKJhUccA/ydqaw9JmglbiATmOTCIPB7q0aco+fZFMeJ2yuNkGxabh8JWTmhAQEV3nX0tm8c7g
sFQgW2O2WvEXjmqaS0GfMSPsMqjvxUTYq3SYMG1PGG/njSkYHtCs+1rifxeIfpzDqZetGWaIoODx
YYjryWH6CL6Obwca/cxd+ZUeK2swI/qgXL/irJiCrGVqbRPL0I9VM8OqI+dG13u8AWPDhbsUaWpF
6ybq77eRc7aQy358NwYNK535K+7HIxx9od5RmVDbWgY3qEjL7iMPQFKtV02zMbw3DDkdMYW+Dd+w
xR6bLkzJoPBi5Dyqmcx8fIhTsaLzCo4q9WT8ZtRLAgnvCWUviNE9hi9bOlcG0dqAYTe7gFCAaSzc
/Dx3trUG9Otb8nsraeEN1/V3JBRdsFebskab3JVtkuCyJSznAuY2Uv48Kq3k50rI4cpqfppitqOn
0Ineu/a2/M09R0tvAcWzrEPCD/SL1EVajSrMeEsW3N87wJqDm1ndAmdzBxnRxnoaMwozwl3wQJFv
vBtvcFje0PLTxPu5TQDM14niLHttPvRpjrhG8sR/ONW4piSsw2u+PO2DLkWxbdATf1r9MT4y9p3r
T9+Te1CehxcWJtJCBQ3cxG5vxykAFFrMs02lwnAx5YAWYsxOLqtqmTjSc+iEk1UJPiMKPP8EAvja
/yfddPRLLBkPQ3wwOsTHKn4koxKk8gYWHKkw32ph6iC6w9dy8BJ7pgxYr7UwabWHGsUWd5ZtmaHe
IcfJp75QY6y3uXDZwumQHWR1sBfxouAZVz7CEd5z6zusj5qiIQvTOWCrpG2hPnAEtkSxg+9Dg6sB
nC2cJRm3pI+xgwr8hFRYprcCpckUsAnrDrkwMpneAb3gQONX3gP/8avthWQi7sKTb+aHhHyRWMGC
iZCu25IKtU+GEnHjKOdt6HLzvuJfAp/Uxxm55gDWR4F/IGaY68Q8XuDS+j+gV6MBkJW2QhCDLOlD
N+CmXMKj9FrXHVsFKZTXmsvbUYzR+aqfWw5dzAWvkZBGqfWkq/uJWu+KDDpg7Dn49TJeFN07Dw0w
rkU8Oqxzt/mpnAR6wVUuijebuBC5tUl9k51bQE8UgOeufk417Y3OW57weYrFAk7BVDdQcThf5FXC
vYrLP35MJ1HMCjXNVsZSjNGzswZdl9Ne1Wipwhp38VzX22PtpAnoaTq52ZeCuefEUluLxEPqRm+j
vJsY5JnFIm2/2Z63gq00Zfu3sbD4c41nY3jHLVV9KYK8gn2TqPymQqw2GH9dyMu2hESUkUMR6XQP
aVhGFQBDSTb4vqj0lwAv4HJn3Tl6xrDgQUemdjRBtEUkJpHX6T7q5t+4A5a8F78H0Juila2Q+KJM
MKRrlUUH/tvMzo5rgExQ8sVPcVc4ZmGtFLsq06s2dme1GvBsiKP93jqBgIxrmmsQkjEsw/j/YaVa
ZTxZYyrwNpE9BYBTnLRaNrGuXUB+FpA1/gyBFuwRZY7exIAS3Dr3oJ/kjCGE9u9/OECA1EO7ulu0
aLsP1lhI5PHUmp+d8EOvm0VGs+bsRV6BZkRMITpD6Jm21fFyJ5RmzCd3UmdYMi8volulIu+ZbxhM
KGP1K0jfmbhUToWrvlAU+hZhjtCwg8SuO6t6kT/EbpOSM11fNkMQ23/8MheIkOv1MZLciZr2mMv8
mq8pkDfNU6czppko67g+Fa+0Ep+upF9Pk/6s9kZdMXeLfupoDDefSjp4cq9vmH1hQEmSCOypb17A
77Atqg82zuBwyTiOVQEb6nOPdpN7cM66+u8C9tFSnTWa+ehq4Sap/m/7akLcaqSns6GVDldoB5rL
+PUJ05A3g2nsr/1tKj9HWqnkNkFAcRAvt2MgqqHVUbu8hpxls1oMRWJ8RstGWSEHZCh0Ffq+mW7C
wL+rmGlzA+sVDmSfnoAmUWgMn6xsZgYF1Z0QfI1d8RKO3NDKRljV0YLXK/z5yJ5zV66gDA+3LqAV
2pSibfe/kFalTsy1U0R91gUyXAk9Ow+tQm0Lut+MABZHuy/f8lkDrNWKPcTeNKXJp1b9SFOKTpdd
wfOfpiMW4mD7XaEe2tzifgdl+zQAVoNs7w/qw5x7vSZcoWfR3HzBtVQioURIRypHORTig6hxF0f4
2z0JHWa30fNK9qq8TbeEZggcxN84y+ITgcgu7aMJfvVj8McdeGk4WjILcYbSVQzy83cO3I2wW+LN
B5SVqyQf/jirCSvHcf6HH+aTZfTKwGAov4n4GYRvvUWihIDE186s1h+WUN7pZI5tkKVNZsq2p1sx
Zccpw/HeRcXws3eawsYVnyqGZZtEHKUXj0ot26r3AvHBwzRqJRah7+CsVisyIa6XHvpDy4PsBf8z
ZHwTRVk82k5CnP1MsaoJADK5axj+ZM554PEJanxwFSBuceNfeAhQWNap6UVh5w0rxXitEqPkzF7Y
+PCcZJ7d6jPQfwIZSZ74AGDWr5LcAc6oSK/wJbZ7M22tYbXKQoyip4qejICVHKp29rawgzCrPu59
iJbbs2Roqs0ogoQ3CG51rxk+nKioh1oUHxYiQ32ppiSPHZI18pQgz4clfXIGVqextrdx1ILAEAxa
cQNgHxNE2UPZpiwTVJmnNPJBufom2Q8qUwpYf3Y4jCvNwUj5D3jwGnZp4kNZZ1tPkJ/llj1m2GXy
VeVf1SUYrIN8UsGVDEwlkVFD30s6vtA9y8IKnSlmBPZz/+m3LVbY6bA3IC63HczG2DL3lSvJpDmF
djkFV/UGiW62mV3zSWLe5Gb6asN+7sA1DKgOMyn13Vej34c2PbTuH846hedr9FZF8goWNOyT+CzI
0qV32SWxt228Jrgv1MShF3Af2qc7Vb5De1tXzCRmCi1b/STX/1wfGuXCUHXze/2ZCCl30J684n8y
p1qgL4MWi4ztZPIhTEpeIpUYdhP7P9pzDIzOyucSCUubF+4Ccb7x4AuRJLak0KG7G+UxSombcyW9
04ZsYwE3wPPI9uNQ1tj0qnR9LFMwxYUOR+ak0x9pTJ8x0eQQ72PfBw9cVd/lH1Ll6IQVlojvkXnT
hJIuF//2Fzoux4iCLNS34acvH7x6c4AlneJ4+cl78jSlNpD1ttzaq+5WFfrIwoZJK8XDQLWYNvUo
BSGrHKDBeXGL4Fov6NNWac3lPxYUJlxEH7tp4rN5SHHoHr4KMVffm2fcwSZiXAemXXAjZ5zS7LnM
u6869FaHcSi3JVuGiXJXb/+xK1koCgkN1JeApT5fywR7ucKRQu263Djek/hC//ln+QALdTA3kNjt
fQ84TO/llPJu/8KnEgr2nDLO5yySFU5RXFUHytm88phSL5Md2DBl8VvjH7W3pZ8Mdk1nIpZeYjfw
JlyaF7EWa9SccnX7OW95S5eMRj7y8noVTPTrGneRSmCR0PPiCqq2kJUrwE+glu9TCa3VHwB5Aaq7
O606AnECm0kzcDPuFPqMsVU0AuN8JoRglSUpaKj6q/77H2xYkEMqmy0lCliWrO5bXZ0+cBqV8OtX
jz//vy5g80DoJDXEDGRYuToGlWNZJHu4vlVgoxJcL5arDda7kzZoeZD2CISjElrayyzgP8qbcUXO
jtskNkJ6bj9meNQlqKGFGbA65OV317O9zctrZbfi3O6uu0UTG+M9bA8jYAW4KB8Qyxzd+1smEPcj
ZK5EMMILe26ozkmvfraSkL+WtPz5jIQJA6tMbx3nUncyrhuY6+NbRx0PnCRGR7RFDv8AlDluMoTu
tNPAWQoqclL5oNM6kDfRu4MdYvYzamomBu7bydsshmJ+2/AldlarQQQqKSOFS9w8gPjCbXaYUyCx
Tx0gQyVu7R3Z/6uzwUyEDkmjiCbAiPBn2rc/L7CjciSUo8c6dy9t1LIA7KdkFumBVv5q3hBVTZYh
BFn5fiSSqxhqOfx0WIQUY+y0Mg574OjwbDvVFyy8+TNeJM+nIK1qgYQ8TfXg2ixSbf2VWXF8OWJx
waAFKDy2FTmh3+wEKeR8nEyeq4CvfNq4lKlzpZCBbJrOvDHTEfAvfmEGQVBQXPK+WaFFRHN8L+JF
8iOWT+Uz9qNpAPesK0vAvMNf2w74CnDcsmbCr/E1D8sSPrihjmF/33Y3eoFp1mRE4dHBY2hfBQDI
8JuH0DGyIwX+BJAhkU/8XzC3mHf16UP0NzDBNlby2i+acGJESp77AkhleuhP1Z8izdvhMe1OCTPM
m4V8BBEt1PmJ/b2RbajAYOYdGBxDAY2IXEH8lO4ixP6ifZ5E+vOc3i08CaP/K5Q97nhS5DqSy/WW
cpSPhvUCsE+Xhg5oMs9UHxRV8ksfqHL8tfpH45FPanAnAKl7w7kkvUrEvVtiOactwdgEk0em4lJq
y6u6frwhZDakdu3sf7Vwo8+VGEc/bbhU6XbOcxWS3xqJ7xwsZ7stRpWRjxwFhc9KfnPYQXNmDnRN
/30Ax0vFPkAdNA/faSev2nEiTPaK9iwqCYSPdVnzFLsojawBFoWrP2iApAidkt11ofWF8Lwy1MNz
TUMRtlZEx1Ag9f7ul0N8ncbXLvh1cxmSJlcfyN5i4Tx8wc+Hbz44/tjmHMJ4mW9R+Ab84Jf75dFV
9fLT8dX5tmlndYRvnHn+5wFQVO5z3TjjUOG3T4gyxT0wFrf3C9rjgHGM0SR+fXnV0APGSrLWCaxN
tI7apZZpY9hn22obLD3eOAMRFLoEaTBlds9IucNlpUOtJn1oJTmKeiHxGkNYb6FfLKTwaWVCm0E/
6hj/hEOuH172rVZ690VQBBEsYYhjPE03pv3Mqo0lTpuKoB57Fqykm98xu0ma3epRgjOst/DSYaw+
X+x1QkZiFy6cLNXOa8HDyhhhTvY16bZv4eXjvvqwVQPDDJIK0jpvhvP1aF68uJganFw/efpz6rpa
dYC4Ko+yyze+rTjqRj0TNCXhxuEFwwUoq7tiYMHI537NHvFad7hKiqssEttnkJBPPJjoiMbTJWmH
XiZzSlXAifN/5C4HcYwoxP/+aXnOEaeEjSDIqPjVr7GS2IzRCGcte9i+jGQ9Ed250z4EfGTWy2mt
V+kmAyiLpb0n92J0vYd97jpsMs74SoIXjuv91CFNCzw+CwC148Utj40cRYoGoIgRlmpNJdKP3ZEt
KeXDvLluvqM/MuDyxlPuHwwVfYOa5J1yBKamOfsvBe56M5L8JiHt7dk8FY66gIGXXQNKB/gqvpN6
ouxXRn0C7um4hSqmnK7OCNNW+TmrS8o6g8QgoxGgd40vmeKevebI7Gc122ShvLQBoz3fXG5YNOFe
zii8Fe8bJ80jJHw5ydNeMSJGlCS6iJwopbczk+9ado0gEvgZQ4oX46Bmnp/4Abrg8gUQQM2wCxAY
3NsdlNIqg32kWp0zLkIzJn/pKH4dph2VPdNENzE/anRMNYm1jGs5nUbQOSuqkPJr2DfWYyFCTGKA
7uIoujyqzCKMmTNBfwQI0RootPeKdS36bi+7jsEQNdHbT2xvPnUpbNf4zFjGPSa8zyQvfxMtuwIj
ShE46oXb+6lIKvY/FGYLC9xPF7YOu0f/6tDRKveiG0uupDKBFL9xBIr6U+A00wAzDWPaxQJzdc7m
TmDrJyMFoTDO9464CrdigArI23Du5qvBpZBXgBQvpSE0RHXEUb45XCfVgCFYq30nSltdRuOhGcU0
YaEPSGW92XLmvyjXgq8M+YiguWDGn4hSlpjh8FT6zrAKBM5PY8JwnUxNGC7XBDSU6r9nPS0soc71
EKjEMe4/hVUGxx5gYlsi3vDF0HKGmjsmX6kH5DrgNuAKyZ5ty1QUo6WSYRwvbRcEd3O+QeatNnlI
1ZMis7akJZojqTi+TJlLYZloPuN6viagK09fpVTwXTs53tr+AzhPY4QBZUqf5cg4NR7pZLvQbjhL
JCYzMkOKsXyEttNX52uQ8DqLY+2Haesu9+pHUugZFDuSd11iS8iKJc2/wkrK5dcLRE30JnZ4/C0i
iPkomrkhgnQYYOcDLJ3WQl/FBPyKpU5DYbznwKoLoGoH1U1tCOzXntoLyeiiT9vBuXlvZpTocCJ6
bF6FACLlwkXF8b3/mmBiuSRtrok/uiYb/uJlmvfzWnRbcfDBoXQ04HqLkS09sIYywP0VYHAPQJkb
Zf4/aW1gLXyuyPWgT57WMwXNnmNKYB5744CgB1HulBLpo6hWKGn8NDJxlykOPjBv1J9nZBUFj7wj
T7/V90S/UIhGRo3D6adEMJ+9s5uzdTDzoav31fZve/ay/bXF7huzpREGVwezaNcaRZIr6gV+0JPW
FZKdvITs6U/dtt/xQmJVdCpBFzM5LfkJ7dMJNjv/xy5zUKNJPLIGFAQfLXLPEK6HudL7+NEX6o7s
U2okJ10/RuLy3tG/LkuVUeYz+GetUxO9ffnVd1aR2xncgplEkdkwWlPf7B1KDgWAbC1DzggliUMJ
dMknCt9i2h/xwtEAGc3BDyOab3YopdFtwVj8fdZz+Pxor37L0T6w5Dx8rY4J62m16bjQ/A8/oUaB
LCn/oBAEZSs9Z2nvALrt2UP8bQ3fQdJs/xQDd5jPaefnXpjVMJHZPD54BPeZE1vM7+H+/eXfaHTD
nEymq4IzVwaUKDZt2ayTV54HzdlcWELj84XXbXiyjDjGRyjAfxzIu6VM4TrswWPTJNzs7KDgUTfS
c89WQH/mieLXtNaRRtZcLpOXvrA2/6tWoLQ5/hRDvwiytBvD1v/vC4023BgbW2ZChGhNFubXoRkV
dUh99LB2O3RjtEV2SjJrmGd3SYSeYmzxdogemRdwZ4LQSK4VYaxIHL5mWQusrj+435vHW9ot5Ujg
0eNVbaYpn8tB7rtzzhhO4hqt2O28IGLRfhK6LVqbrqU/ikp2uRcAuXdZNti6o5SY6L7Xmdkl97Y3
AlD5aeMLZ/dsJ307L2vGV6oQ5b9aebZJfZb56yHSE+xi6latRqnQaBGu0zpuJRbtUZSweyhbiqbI
Dw9++nyQbsc5504bHofW5wLfv64HrGR4s5Y4VrLhMJRdqIzQ/eDQ2UZ6WGZi2YJgV+3aUdPUkSxi
21IpKvsXAUkzESnhwldqbQCIfqfgx4qxbiJ22th2bnLgpPgEW7DwqCWVjp3BP3cyDP5qTthxUsiS
HBRIHbZHHlT1XOJEFlYttNowmsPKOKoiACvr6WN8k8mDK72GqfunXtuXNJpGCemwHeQuwrKVWcLO
YaArFI3YaxAeorEt6cxbtmjki2Mom6z0nX2su5vFrm0ymC6QaZ9kV1M+zbJ8c9VCQtL4HOORPKT1
w28OoyY/wnEG4fj8zg7S4jMeuQpmSlGThDr5DQ37Cq100Pa19WECloZuJyBi5JjJGP8yf+50jVJa
vU6WCOarYOPDQdJ4u/epcIu6VfJ4K/z6hXMf0pRPDwrgqdarD68/hTCt9Fd3toAQhGt1pZsfggW2
K/b8XrrvK6W1Tb03gV8QOtCRjHnug6S7eJtnlzm0xhZaykxzlsu6Oj3bHn6j/o+HZ9zqbFFxotMz
q6yX0UBWvIOUTnVfw/en7m4HbqO2Z0W8gyclVx6yUFzHguyewbCcN6UABiwzF951y0O9v4XD6a9W
940cJw0iCcLcrtkLIjnXOlAV2GWVWwEQR00m/Q4PukEQpAmTUQeV1738PXzloIb8GqDMjtuamlAh
NXr1QikrjZWruWSAOjQiYZ8qBe05vgCWf8vuNI1yK8Uqn0+sGBtR3y2UNldLjBvn5P+U0VdIsliG
ipbBy5CpzRtu6VU0aMIp8ihTReSCEQX4ebqbnNFVIOHwScRcY/FKQ0uYd4J8MlDUceNUhLvYDCCJ
GyGaltafdGRCw6APz/6Ok9gwRcMtQecZbiXqkdvmH//xxuDDYvuMuFeZ3yoS/c32JCyPXhp+d9oY
+Wqe1ni1UuId18FxSbcv+e5xetbI/oYg29hbHnjro1JK5li7tSTNkODRI66Mnfnp8qnmiejFLNI+
FlCiwdPrSKCiDdGajPYqdUIVzXuKjKxKHJ6aKcLSWCHwmUhOAfIdLz+NKpMtwOkEUgGOISVtgnC/
Nlpblr/S3EO/a0mB6mG7f14so5a/uVovxkfDEGZ+72f/5X2Eb0riFGoUF9i7WztPO1M0xww8cRPc
UAbozGWyKC6n+yJq7wvmAwSBkbysSrRKSXS3RXcIoN+nk/PFLhb6ScjMYVHBT8jpiKfQtz8S/edM
mCe1GQn1Zm5539HBxZ+tj5RpYYrRCdZEp6f3uokNG/kZZU6Y0ucFtlWYQ0j+KJ8DqHqT6uoRtao2
F+f7HvYbCewRx/ccEhCINYs3/TUBOSacOxrhky/2kNibpraVHxSAWRoLVx/lhGS0n6Ca91GZ9VlT
/lWzby8cZOa7pxwe3yorZ6eOHeu0DrqYXCPOlBpudg5PbtIT6QE90rvmAfgTqJNN64RwzeniUQc5
sHDox5OyK3EoAXehFC9gyvz07wFFDEoeO4Ji04Vy3JUYWnS9HGPsDzHNfM9bAeMjEGIlvfNvXKFi
tzzGQNE8OtgfXmJWO1ImOOl4Lfae2Uz8Aa4l2chot/HFDsuoOwRtFECu6OyNdDhF4sLt1qKQgJMQ
2ysy0uk74ICeiwKVHRAEJfKkvYhtYM1nRS6Xqz1VqkOOW4Hg3IQVDuygo/RnmhkVHy5szxfYZEzc
mduOJqbXvm3kXpyVJG5sciMmb8nJQpRZ5Oln2GoJcpV+DFJkjJP0SeOoytzgirlvius9gRdL66gC
cieJL3n5fY38YP5cDGPfLIw4bp27WKxWmBG7pSXjCLdghf7ewEO7L/2+38DAe2zN2bbHxSJmsKg9
yOBCHgcX6f4/1Muvrr4BPBEto1I6PghDENZYxfEtXT4QzWo2xhi+a+XxQN1kgtZbWoY29xsGhKfe
QqTjk5n8Ord4vqkN14QjQ1gnPLhXb0rjW/Uj9r360IRuO25anBkN251GmurjygrU0LOud2zrkWhU
IPLrdChbKxYJD59D42nSkLKoJIyXHUGHhZ5l9wlRYCN331j4Er/x2gI3GhdO9fzR40Do+L9pHXn2
eGP7fDx4EaLhqiQr3oafD4GpDOtWIPBNASMR+drpaniut5L0PaJZz4rURuHasHKD2IXyK+xb4qPp
jSjZqbieFliKFQUvSRP3BaXEwOFUhHqQfT2f9lQI3NZRVVa9E2KRwFepn7kAGXZ5zcenCKesAIhf
LvsMLqqctxjXKkbcMgzJrsp8uHtCU8vzeU4+22I9Iznx/1XeVeEcDaEJJyNBMOK3IeDMIJf/eRne
eyV3zHByiLcYy1McUKDtvP669ho5pSTKV5SiLYZKhTvEHB0n7TfeZp81CPppDRL+BwXVtZCJ1TWy
evPoYmIYqZ5NFosvriWtjA/EK5/x5C7oeRaJU1Qh026nn3dJ9RTCO0dgMPS2iOA6Rfb7XmckNq56
0brwG5oyNg+cdzGhD9IQttTtuAeCM58IAd0+uqciXj0+tYhlv1SDJZVldi2K6aXIs3BxmAlYuQAY
JxsnXxnBd3ej9PmoshackTLN6LmYuZOFo1CfjjtXdTVPoMDHJgHjAdnf93un0ZjoWc2qkkorf12Z
Kw2RVvJBDhVR1jjiWyR/LFYn9uxtzx1iIeOWHtLQkjUmkcDHwH0Z4LvHe7TveT3sxwzVpa1ikWno
TruvaxFm/uoHxEQkjk5gfHPSPUP4nD1oFJuv9PMOte6GNaBmQbth/PKuTyxLe8CoGSo6tkIAIBTm
QoZ+OPGzk0b3rBAbrYQ1/e84KHUCWRjbs0oObbycUHdIceOHfsRjk+6rm9w95CsL++WasBMmB6w5
KgAkvWAyBb+mrbsyOzjEr64P9WNzZcWC0yTLi6JLRhCoN1LXC6IVd9uuajJR3Jx1vjKAkZWXlGwI
IrJ4+nxIyuobtXzX2rVec+5cMLs15LXziju95eUowzpAXVPlCXaPt6UPAI/RZORJQXxFTV0u6RtU
OBjgVS6+k9uZIy9wrBoCxh8cJ9N2/2AzB5EpA8sx3OD4Hjw3snqSwAf1L6y/a/eXD1W/ogdZ3ZAG
saUN8zYkzqKx82ERq4anYwGwWoKFkjqHNbQtpXEe6AW4v4cSdCYQMdgCS+g5R5o3ND6zR2qnii1f
1/40z1t8NQs1q17V3wRctWTg4BtoaG1o8RfucmrcVIgUqiwxp3t8UftyWS3IAOXxK3OPEFnsZCxO
63NDJ2XI5XJx7z2J96RJec/mY7/X1iCdTP9bevJoIjCCQN1FKjstl/O69GCW+bOT+PvhS9pJHPxf
E3+X6aXZNGNgt4mDUHttVNA0Ul9PuFIKBLSwBbBu5xA602JIK6NBNcnSo517FtyqlnjCfBqZCoax
l1jHDWDhEqk/Ry5FJ8OfSXASO8vDzxIqqwXgI2GEij08bQ1Fu261ZuhFcBhiBOvyyDKbPu1QA3rU
vk7bwgH5Pud3T4rcQ03/pOgSeEMuB319LS8y7h7nodtudGDomJEGL2xH+b89vRrrXqnvbPu0+I+b
oBdyl+QJvpP4MRcQNR8AMbovE6RnBgcSonouAUNKzU7FKG5NjJQ1h3LREeiCPhMPTYqhDuhGNBMI
yIBa6TGQvUqViME80XFV46uact5kOhzx1hGDQ+Xw2vQpJJmaww5b125roUd+LA4CvZDWchZKiiQX
aIpvHFbuSgPTY7sNUDmIN9pUknAuSNz1LaHTamUf6IUhRK5Ctyjue0xPvx2XtcG0yqwODHgX7zXd
c5p6XPljOprKXH+qp23yuraZiXWkC66AjwsEimGhPBgN9s8ph4C6tE2guJyWYKnFC23I6jbCrqBE
RUj0RIpDfBUii5BtNVwIHq/5ob5guaocXFmKIeRINOaZqK9ayr2gFVxWnTL1bgZTnSCkZ0jEApps
fcoeC4fiE14XL4GVjlhMMwP1yVO+cZDqECvRK7BGVOojX+vmoNPRzDdfNHhapOoaW11hKLP2NA2m
jpDv4q7AVpkbwjt01WzqF+wpXVkt9S6IP8Bitw7DU+1LxL5brR7Cfz5wbqfzq1JVNn03TXfDd/bA
OMDCdr3Uk01VCVALSUQKKomBzhZezxFHHOwF/9zC2j6CWnD04jNznzWUVIxwqmSpjAcPwVy/dBYQ
doFSNknM2+YXJKrkz22CBUnk5zIe6wNzjl+5QaQ/6vn8FRa/RbQiOrDxf8Jggzd4HFHXFdrtDQWd
VlvuhZrhMClyY0IiAws1DYKZLa+dnqKmhaDJIetYAHKPcZ2DJKnZd3uz8dZWzHqaSw30VHHypdMB
T9gwG9YwNaP7Vuq+uus3ldqu/Z578KDPoYAWDJ0p1CLzt5oDTyoInO8DSHm/0gE8Zz3VIDm94/FX
XzbGYLAsOogplad7AfUTBFRX0tNXps7IM3Br0mFO7IV6d+S5psSCoXytk++AfLTwkDMDq9JWQ5x3
sNnSHzUzwWC7jmSFTsfF4Jy4ooi/B1VO4b5SVz0X4dB107RNHkrgHsMaPKJjQ8gykDZ8S1jvcwz5
O0Pa43twncgltwWBaVBHWTf1r3IsX2bOvgwKc19ZNG4JVJWJJi1J/AUZWdSA21Yy/odeJSAbHvgP
LtdDdLJbZCwRQFzaHkok/6VJPyQ0p2vjX9LNtkGfu4LgelnIbICduge4Ewc2nliB0WWn2bBL8OcA
rQ5zygfTCL1VH8Y/Smt7s5VABWdCZ6fA593PULevbdGP9bZfjwYbpCxoQ9S728DslfzxM5R3wLjX
dOMr8Vpv1LaT2q2pHyl0UD4872+fAVrRh2zxSrJB8NPGcgcXmfIFWCcWhdceb283hSlckNTNzYXk
C8k6WEfvLzIZ1AVWg8J+zHoH5KAmF+eu6NIx0VlQb8WFYLF4kEdHXnUeCq0f9TKw35Yqc4msV+8c
qpLlz+Xz9QWBNIOKJRC0cJXN96o80DXmiN98n5WeF2XQRxzKCGKqeOt1ZoGm/oG+cPikfLpmq5x5
qcGjMniJUWJ2I8eOV8X0tithAqICPAiKO7Hv5BYpCMXjYLXS2SMI2/no5tddDZBe0ZFptd5iRZc2
sESu7DAgGwKmcGRW4AXuaLkQxw8FnAX28b0LK/Hz72z7yfbsxZ/aWpfyxfSuk4/bV0TCfDHCoojN
7MFE5/e75zM9IwcAkO7DjI3H0FcSa5qvVE7ODBdzVV2xO13SLFqsQDbsCInDzgrR9Y75Oj0Ko2Vl
20Inwm3zAoA8QONMizKjrpZi2CFVG7ZQHxjQzSSZ3VpgYoyxCXaDIzrIi4vXn752LthzwngUTKrA
KsgiDHacauKz5KJ57i+0Eo5qPblH/w6V8EXyuJRqjtzsjMMZSVN6BfwRXzU3YO7MCSqmRE28dPXs
dQT4EtFWMFoIXMDSI7DGgM2onY73HWghr2gt2uTTsl4YpNiXB6wQ/Hnt+/TunTqzxRdgJ0U0PUxh
SJzI+D4krTzLX81RCmv40T2KFym1Ki0u0+cjp55TCQ7PwrqrDRftH88Umd8h/2f4Zlzg1Pw8moQS
JaM+JTvVVs+4L0JCqLwn/iQ+jGBrvjDOzfdfkacBDrxwk0SBWq5ls30lF2CXdZwOT97xq+v2BI6L
eBB+S1gvvoZcweTcHNMWb1OrjLAsBCvv7olBEq1NhHrJwt0lh0Qf9idCtaD0Im1x0OAuG9F4APo5
NYSk0HoPji3MLHba8NBSf0hmUpFRMf5oETxLJ4cyIzQ97syiC1lH+MScZX/+SPEVCjOz3zkQNMVW
4hRBbr9bHfHznQqxqJWftPC+buWnHPVrP8F/TKyHoB6qAC+zoAbs2L5extNQy5fgZB4BhJ5zVLTU
I2vseezf6CmG2PUgqOz3/GGDfMG9t4GnPIGd9KcwfL1vjPLePr6ZMci6qIKZvo9lUmy520NeUzoS
umfPgC7LrvxoL4DQIWteyuU1WxB8ljwrDsFxcSjgbmKv5qH1Vf3Zho+cVXkdvRzP1g/6ue1mZnHs
5h4d/ZrZ0ZNIyJ4FiD6FEpsv+bZIcsSm59PdckJSoQ1zFYljgyLp7dvjuNT1NAueXdgjEOJd7sZr
buNpKd1s62OS4pMFAmIXF5u0x+GAkxTgmOnowQKCQT9a+jI5z/GasgNU9/UORao5V7CfSaNCXQYI
UeBhXKxkdVEjuZIPPv/QivH1irOLQGC1Z5xBd3iG64lgkHqHOOvvZL8G8FyZZqGG3XMxhPUGkPyi
HDw6R3Ig/MpGyxqtLauqpI6hp9XuslqCpcV1zPotb8SmECvMK1lwQ59TU9yy7+Z9/OJDAm5Dlj/s
mzKCIiRp7BSr53hi4GECmOSlu9oP6gfaXL1ar729MFyrHZYPl5t2DZg0Nt3cceVt1cU0A7f+sroA
X476r3+TSP8UvZsZLlCsolv+NNAawYaeSdF3ro4rjKSnaeSS9MJdr4gA2qzklK7WNh0qjn4bktcO
81Rl0cpmrieU0fyGSvMci1gJsnEg+W3aYAQQAhULg/BHHaq/ll9WEmW2K/v2b2Ug9BoironTpow0
VfYEex2MUsXbCT9UOe4RehbU5dd5gsHHofCLFR5XvkcnwRDcooPRrnPVg5lt6y0EaLsAfF6A4ZbG
2HUHs+DoexiZG/NY4KOjjDUKks9Y42AQVudA0xfBva6hBscvNmO+YeJEol6Zi7AJuCzNy5mgSHzu
i5eRdltW6DAf/KD0XR/hX85sFNu4OoQLcKn4q+tepYk+gPVv96iACVQOL0CxksZrjTZKHXjCoH9q
ySoKDW/Vck3vDhxU3cQ0pygeKgcPHrx/FPAC1zYdwGGGiQ6TXsPdmXkS+4x23rT90gN1tcDVMmsg
F2579V/2cg1H83XzgjDh0C8RxKNhMJi9WBvF+ssBK0RysgDUyWggxP8/7hU7z/S4cVvdaVIjyCQs
cjMtBRmy5HqrNhgtP2TVs8utQAi1r1JLY8SXNWGuEN5WJ6kI/S/YfvhEOcA585ZDLbYxga4qWn1o
fOKyztKKZUNEiMk9x0Vq6V91xcP05eFfmAgInLpXuRm8xOetYelZTB9dQ+7/1jOmkGDEDfiM2BwE
TJi7cu6Kxjl1ikpcHGTe4ge3ghjKnrc24u5t/Ke3VQGozLkr8FR/oIVzgxoRFeLhLGAxP9WdE01n
VkjAPgwiUt+mAg9nZVUYC1DdZm9cWOPHQInSSPQM9267ekDnsJKKQTy9S07xXviPGD7o/BekKprK
7cw8wKID2/sj47h0OLOJXCeeznrGaYe0t6QU4WzuKo/lUYZnhzFWQqOK/avesguW9yAelg8htP3m
yMits4iRGzQEA04s3cd9Mb3oTMjpVm3+lVzMhaG9tJKyIm24dpXSAOVPeoWrRQIr6p9HNtae+ab6
RnuEXAMoLGBIr2d8kss1Ro9oydztQdFIuYjx296R7MlauLZhDiIdWVbRkWlx+/CRdBNTurY+gm3N
KfXrowuW65Es1I0wTT7n5qzz/+D/QYcp/x1AOmI8lyui32CatjfeuujaPoGqsCA/cEybu/9ztn9A
ADDxk6WK2q+JYbNqojFl1EoImeyAFskfUfUXlDGT8ryW3JqejhUatrkvShmGYEPlDjQM83KSyk3C
CPmmD+QygGGHbrGbx3I1fW8a3u5M/63t/RrEQC38xWOmx78sKkvOMkABeVt+DAW1cV9g5EC1hmu9
psfNBhIxrvrQXFp4Br9IQO0UsykLwcU8cmvIHdOZyfqqrdQaMS1WQGvabwV+giTI4BKblOrl/gsV
/f2FCKsmAnXJHV2k/45taIllwouHsoir1BblwyFEtIYu94Qy7YHiWhW2AKxA+m+ZJjmjqUya96YC
qn1/OJLCh1nLLOvXOasX6gDNpNjmwLtUOGDIeYhfgRdBS5hG6Cx5iUv4GhpVUo2UXwCd+usRhZmS
BRALy6KC8XtFQKaJP+KhkNnqcCpnOWbMmxCxxyRZBWuq66nD4Rxlc+GI6Ua/+RqA7H3zdGQPZMsk
W7gLMJbyn++08ELFe8b1ltkHWEes8iCWnW/BL+wqhBCeU1I7mG/ptEJ9+VkDRL+3gsGTJJq8FiEu
NWO1f60p7NKoxAl6rJJu/5NA5dzp6ivZ7A2IRoNnmhneaeCO6MtZGR4AonB/ubPmoSQhqM0Y0I/T
didL6lJ0nZ6vs2eRLnW8UHuH9Ezf03GiL7yT2Oc9evIa9I/REb9f84sSrnkYYFMG3KZD2GIYiCZg
b4gXcN5zbgy2vcKlTgn8YiGYxH+gWIM049gz3/Nxw4H3WY10cyGQs6pFJAgU/18U9C08OuYshDsa
ePqIHXwMudJkBr7UlJy5rVYdmMSDEv2U6AaEWStDwPjO5Fl6AHs1PMAipAzqGo7insqVLm1uhUp8
CoVP/T3mMmUegUix6f3V9kzaah7DKJCrigUOonuUyfYR9Tudv8pThT4zlU1qo/pd/OLjV2BRGRJB
N9Jto9bKMGLfWbD38MYMG0ottHh5v4cMjK9A+v77J/81Jwu87gZGZ6Mcpy5lgYwZwkgKk3/bG3Y1
nU0AGrAyRUHxYzzSoA82ZVnmvpz8oYstmj6GH6saBWB7Jx/xl3BEewjhCNN+VGdkEc4VRgoKl59C
UjombMdgCT8HsbQNezc22pKtNbN5l0/0horc9mD3mB+Q/2ysXVj2xjhAIpq5XhCYtEp5ScmzPdE7
88UvDXNyXd8W43uVLBdWgGPKqTBf71uMlLsqkBzFnh1rN1Q6MEIjQJVl/8uo4o+7u9i7UR6QtkLW
FBwyhfhvWisi9H0F8KizlHGXExarRImZSfp5FijjPU88H+cMOveorh1mDrpFlAIvTUcJ3PX5t1ec
TMfDjHlt9HQqmlTFFDrF2TdJ3s9WMbJxZ4E8lSKSOL5X4BzI2qWRBrInFShfZxlrWqNqTI5+ap3z
bZWI27N7+RqdmxwctbhXf9x47QJ/toZ3oLCle5xJQDPfpKwxbOCwASyGx1hzRGfudK6CXQfHpyMI
7xxRGuHPIyLWRilge3CDwJOwqFCJqfg/VH9XR9rQWoRThGdnJFgex6co3RexDfwrF5iDbjl4G45j
7DpqehgJamQ453sLyoNhWvuX+MUFoitQQkUjSjTRQfmS1Y6x3AKtVZt0A6fIVGYOh1RcGWdVYI81
xZU5L3NL96iX8muiU5wGuf/oQpXf2NSuQjarKLqSGkcsLj1//bFbVEbZzJvx4RV5ALyDExUZMBJk
G3XTUDNzyhIUs43J97qjBv3VkX+Wy+fK4QgBrZ3nhc3NYIapj9k9TQiUfftbudO20Zo5rtKN/e4b
D3RUHhTwciTd+wz6j0vjdu4DJTlmb0g/BGMJsKHfeun39bzs4adlCT/lDsnrn63DbuvLqX2DQCKH
IgC2lBgKIxMj5FVEua4x9JBglATyE9OGmNJOjFwJ35nb9Ca397ph7/6wen6IpoiwMA2f4/A1M1j8
FP5hxiypIiW17+D2pB5ONXSuhTLGbZ/HdDGximQnyj7QIKRDqJvwIo/+zXcvCuehm3QY9oZHvMIN
0nIhPzGgUiVeZ9VRg36W25GftDqRDLOsnIbEcFrNdNfkuOWU/lAzgDNhpiCzWt284uzhRM95cmob
lDwKcef5RicvB4c8/OK2uoOe/0MjLZotU/JUZ7x5pPrHR8gf0G6m6Bk+Pp1/Zb7pMoOmWD4Rwkf1
Lbd7pvAMEGGVkSlF37CzLPPTy98B6JiYlrpF4hLWyrKDSYSg/OeqjkwOZLfAuE4bQj0O72BiuH3l
rA8HTbdh6LJon9LrGRlFpUXAy4TuEEDV8RdLk7kTlwDTCGA3KMoeAl8a07DJdeWmPDTC6OkDsaJg
e4Fo9bHugry9wxZB64sKfXkmLD9DXttyFtEeHMTEvIy79i0J3XCRwbiuBwSXUs2cKQnt4uBWWG8H
IcyKOejnFoTlptxb0MAPR7cAC2kZlgXGTgiCaunV/m6dYftucJFf4tuhkijUOacVlM39peGqbys3
9yY5LiyQzZOaCEZscnUvv6s17mjuxhzMaFSh/UYHDrAuqt+kAMnz4ijXIJ1MXd6MyaWVDDZd2a4g
uFeVkmxHcmq28juD+WvKXUfSTuZB5ScwnxScJcj+oVaGAFaWHX6DB7O39owJ7/VIqxds1tQRns0Y
GNE2PuF2ohoVDuc9EFq8BfZNZXx+bsuheRzPK3U9FZLqmuoi2GvPm28hpEFP4hibis8y9Z8vcJp7
SPcqqFblLbbtglu3X3iCFWvrQa25uKjVTDy/cZ+iGCIObzQ+tD9NQxwJOqHQ/FoJGMK74PzpCzwc
ejeYqWLECW2OEstyTtn0NH8U8wurq/h6xrP7fqlMZLmHp8Rh8k0l8VR73urgWKgUY56aEMpeTF7S
YMF+BUpf/lwAn8AJ9APz96J7xCrKsJBY1y2+W7+ylTI2LmXCwrWqw6D511lEI7feJuvhjmDMpmjR
nddmcDdU9+NUNVUq5b9+l0RK+eM9db9tqMFACThjoKlN2arikG9kNIDsLhdzN9NNX7Fk6WrgvIZz
L+LwzytNlwm/5+ZKBPnnh2chDDkJktUoNbEo/FTMUD8TlyLkq3TfeSz43sRQ3AHsUCkoTHcv36Zy
cMAxMceyMsbLkh9SQ2TLVPHa6lBZvsUxc9shtFJicGdSZY5BuOkaS4i5c6hqXN6NrL4YT9GUV3RQ
z9jp44XgeeyhiM1Ymdiw+o3AJ8FjLrnWbRE3YygbFh9rvexhzHHdxwFNFyHgoEKsSS41HVQ5Mt36
xMKo+yWaCUw9kHTbLdORU1KRb6grvUsKNcEqbQUtvNejx4Ag10BuF1zcjHcrFHMuYU7sgIT0LTK0
SZ0GZJmmSmI6UdUdYLgTP3hKKUc6ArX0IpuJ/p3EBO7I2Wc8tyk4I60LMD5rivMj5hnYJPFBbg3v
ccqNALAgKnPKcC5a09D7RAeHxobdf3F5HeVmnMAdqbWIH8Om9sawLgaDcSzrGakGMiUxdVry7Y4n
CwU0N+BgCDi7DcE2QWweQ0TpfjEJq8px7mQUcepNP4+zjUod/aX0LlF4vTB35pCJ9lnkeM1cF38B
MeY2UIA0sttQSVoAVnpzFKK6VmLFHMI8C7aXYS04uK2IbjfmrZPSzsVieH8jOiKn7k8LwtXswTZx
g+mQJtLeiktNoQKmdLuN8tzuez7CRi6sv/Zwuf959ltG591jprPfKb+DUDnW0RIQfu6tYCUBTptt
Sbds0jJf0TvR57UFZUaYi5FGxpeusEeikJZoiuGryMeD3e4sXOGI6LAV4XqB2FCWr/telpJkTan9
ejAsR3iomBosuklgFVzBHOEPrG1ZCSUd1ahxMWQtEyiib0KPE55GNGlk8pMftI9xC/uk5WGz8OUd
Plqnqb+Mku4a0YOajfidCQOy/zIhVzEBPZc6lmhy28rAYKJlZYkVi3QO8ZsPSF5hXFiuBpOhMFhO
DXC3BjM0iB7X/JwZX7NI/PQvQIIHSKsmdzzvnKKiU/fIm7+CfPt3eI2YEWooLHik8B0sp3wJNfo9
kxHPqNsX9C/+ejsvTe8r4iHAppuK7mS4/aVnvCTcblnT3V9QgMkPgKA/yV43TAMQL1ipJr1YrDyo
+pzuBLoJL5O2fpK+B9/Yx7lQ5soZSRs4RdemrGKEtL7dfbkocEFgubGuD7izOrVsjLmpvljA6TY2
nC1Xc4bZ0EK7dXvwd9eGER4tVdYfS1JwgtSkDFdBGZ5d1iJMSn7N/ZAaK5Pk0Uh4Q0T+rscYt/PP
8q09yzOQQPWE4CX594KbdVErFF4GQE0/6jVMKIVZTo+NqxfXE4DRvSl6CpPBM5404ZWHVtGKY8sU
ogNsGBr7WNusw4hd7mLKvSaxbyxoKffX/uCzO+hTm44AfQWcoXLVh7YDy5qT6w/qn2Ajij47ABYV
M1QMFGfgGwoPDa46xG6IjQjTLT2Ga/VC8tkv8penvp5JGm4gan4CySEDtZ2tH75jd5HlFf3lDqfD
kEiTfqd8pG5vH3LKp33T7QPwnc8Y3C+b14Ze8SIveJ3pp+w7mGWb4H5tJ99/mOjoxGJISlnW0okN
bUTasw1Kfk46yVq/RDw5Qr7NlI8QEkRAo6FbKneggUGKpBFsI/uDEjL3emHtaqdYR3utzaMNdL5T
8f/WpynzYHm8lj+6i8LXP0xxQGk9/dYzXbdTS3I5CH9Cy0SQKZij9pW08G9S1/QkPn9f/h+IKp1q
4ZLhU3jOha3TkJ2LZfc0o0fkn4/SnqOfdwj87ejcJ+HbESqw13IyAfYhUjoL3b0R7mP/P52jmp5C
DvqxY6y+4QGapuhDqL6Yb1F3EOnvhYgT5/mTUAC1SoA3swe8n84BknS7Q3va9qVzuhjTn0w9KGNZ
KaDRSKyZr0qCxINV1ydM++SHS1tZ+562d/Hl4qj+OQA8T0OAZ7FrlSRsshcFoEhGVQNVPSX2EqHp
dZL7yWosML6gI6pTIVnTOcAkaP+iVKbV20SXitN6jjiYkQmV3cTHSrxxkCM/bXC9s8wOoEj/sXAX
VGNHHhvufcTxdD/Qs1LcKRySu6rXsJdj1pNwC9ecaYD5iuAtYU6wBa3zpqPyECy8FVAqd/QGvynR
YSPkT2A2fqx1ln/FVb9z+W+f9fj18ecpe834AEC/C/XzxAecDtzhelhl0X6+TgCzfa0B+hQIasQ3
FSYSNzANcbPJxobDHmHJ3KCbDJWl9cx9wWGRMRFkvTdvJHdWUZXNVb2tw0jUseAAUAd2ehqVBz1C
U/SnULVqAG5uS2xAiZRdEW25quX3/JZfKZuGXhCNZZPAP3okwoIkginwyew8oRfIDOENcLliiLtx
c8m8lg4JXaFI8sGxDbcz2vOkqT1Z6nHZWLvqt927j2BAVtxwnjBtVc4Rtsrps5YFiO5LSFqngS8R
7w1awmn3M2fFFiBHwZ7J8cGDLFuLDeJpAizXpOBzNHsBjNkeUzWzvPguP08iNrNJShqQagU11u8P
Z48jHVg5qmy6ZxaQYapTb7jxsbwJZlNVHZDZBsx7hwlCEpWYr6gTCsqFdZ6pH98wlUwWlY/csnyV
ibW+iCzxsUEzlq7/HfJH3vnCgTgvrx2naPTpL5Rtj9ewu61jnrbJOBwC2tiEwbUVPoCadgmptqcL
9RK6fjlhK+MFQ1BDrRMNGLjS+vQ0gJR91kHbYe9dTYj/DsPAcqnt4oRmDeHMrMRx1/CXEpEqqziq
LbeV0MWgXB1wx8c7ykc3YWJ4FiOgEKuMwmpG9MNzVe+t3jgCqZ4FwXep9rhDuInhhyOhuoUZ6E/8
ghWFTyaCpUKSxThmhwjwcqXBcx/6HjTASLoKiS9+uQhY0+9rT0l3np8NtKsGX+OhFET7eVoCBEtr
AoP7XF9Z+UtqoiB3l+qZtWNNelGJ1JSnQaGHu1UWaYeo+Yk4KclQDbSTT45/UfImyjSYLX7FXcEP
GwFzaR+0nS4S5goH/JwTnIVAlDQoLjtIpnf4nIHzmlDgBqfZpb0sb8k2XY9mIG/6b+F6cF56iN0F
saAkd7Mp7fWqxAjBbNGGhaR00Px+ALPpgP5UJkOyn/XyGJ9r43Uq+EAWCaHJkpO/cvaQ6NyHXR7I
NorRAqELp416HgvxJ1blxyooglyBy/xcEaEbZs2T/wX4S5c6dmQOmWs9OSdh5O3Al7rxfsFF4MyL
Kvme2gXPwFJZhElm/jGAS3N8JZ3zw5YzLCwU64c2fpaKHDYPUD9cLxKvhF8JvnJ4Xqp+GkHGut62
eBlx3YIbWi0t/uAEPufmJVmuUzPCwTv6Xd5qjgY5QA3z9h4d3/j1NWjym5MU/W6O3/NWFdvQUftu
NDQhRXC9ghB3c9T0gADB8IbPGDORmxFcTLzkUaZQZtoGPwK/dhIvRSgW+w61DJgpz8klJDV3pOQW
xO8fX8gga6ynsVM3d87fYg5xXcEAVZiiY0tyiRkPnkvZmNbCHuOcaIgJsJhlgldy1xtvrB8MV+Qz
ez+O+5CS32nXCgweKmaLoV4MHa400/kpRR95uKAl5xGM6SPEmPzBP0q4NAovHWfLzHcOs41+IHvf
IaBQnqIpFbwzOZ/W7eJyjcYr8NjM0noaN4+LFx/h0SlidZB/m1CPtg45a/KZnNhieqi/cbpaRm5i
Vpy0dSdGxjDcBNdJ2x57X+hMrN+pcOnEFukXGYgGKwJYmcCoLek4tmhaU6X/bHqPGCkBWVIqozPV
qwy5wZ1/l04y0XOA3RV9I6l9Rg7Xs1q+3NtHPVhQm+mbaluo41FCCgDeb8ArdnRnGQwaIB/sOLyv
SsGjofVSU3Ksx2HnLC1YKscKWAmFhh3UN8MwPAnrIEWE8pv4M59N9OR/WFtGgUqAtw8XQ97laaMK
026XwXl1gjgOuKx3Fd19WqR1B8MIbBqwxd2zDryM3qQPYq5btlMIgOQiebyWG081QBHo0j2ldD7z
XsZzXufdrRxzuZK+LA7hRB89PSEIuyzQmN7x4iaXr0OFW0W6vz7hxQXu7p+M443qdvhWue8/wVb9
fDsEJkJzPAvQ9W70WdDZVqnoFaOuLyUUuu4/qmJTKkXEblwQSw6ti+A5FrMdJ0dxInPq31f42XTP
5lg39mF4xkhi7Wf92HUkIc25ksu35bjAn4oy02q9Q8axLFj3yOoKQc3S0cxv4omrfQ26XLIxdMtN
MEw4F1gTB//YEgC8p92UGd4UoopeLi+3bk+lOiiLmWckLvkURtzXbOpua2WzE8RwSMDZnjJLhPmA
uhrJWsp4UI02bvDcPBGdytSxg+5IeaBtUeNkLDvhsc+WIaer3tdioB4gDm0S5+Sm+BprInplSIfZ
5AosWA8bINfm3F45/cboWeOFtdns2BLhjCsZosqAZrkH9VQVIii/1eXZ3/25AR/Z1WTnFk0fmJsj
kGe/lqinddEk9j+Nv8mHv+Fng8VuopeKx7cpPwlfs615O2btZ7rOfeYq5IT0bTeOc5fQNR97V9uJ
de4J57fjqkSAqmvUNIZfQgwNo6thTWudeRmrZJHBBpynjPtR2Fy8FiDCYvR+y9BUI7cRMNiEZXBc
lUXbE9YHj+Uj2y3MT0A0jstGcGnVuc8ton99Yz78ZHExJUZuzKoMq9VrxUOiB/tAVI29D5QsnalE
LSwqx/dPsQ0gQLCVT9yG9VydzvSSO3Yj1ANovFG9HUWDnLjcTIBL4enNs/xS8wDxnuOpUeTJOFjx
KLCNVrws5r+d9ZcBByrUp5VPXK60mRNNnHrWl9cWfpXFEGfkt/g3Vb7iJTHAkICQzdsqi4qg8BYU
3R/UIGnxxBJGS59eEFEYRdMIzhAoCckMCofmlkSEL4MwSjXbaUs2iunBOgviFcbdiI9H0knZe3NC
kEP+ymjK4hVSUNrmjSNQmww/JeCmLvDFQ2F7v7aCcIIelbdwHtyU62kC3tsSxWnFVKw9ffUddyMk
iwJ3NfZul+HiaTuueOculN4rgMdUHLI0fViI4TQF2e9FTae8806ndhU51LrFilUV7IKlrFDFpJZo
RVq8RntolE1wxPqbCPzz0SDHxg9Jb+HCRXJY/RDMq5zHSCAzcahugROIJJHlmst7kTt1SVI8lgr4
WwjLJAiuiGiA3ZSffMqvDTnQqFc68lvJa5+FV/yqZMJ5Emq2N8gP84fX59KzC8HWLLIvGGwW7Wtc
6WQfVjuO1RXNCLRtoyAVF1hDL2DesiMJNvjSv51DOcrVZZC9mdTqMos1VrTUj6hJnuYBs2ZpnjjZ
LJrVOv0yZ5iiveoVBdubPu0ZZxy1gz7nGjqdw7pGvpYvvNUZFc5zqr6dJQO+VSjo9ylV3C1fnf7X
RdqemlJ4ruW4vv1s/5idHbGXdtqS0P7RQi/0bIMM2Yv/v9J+dZ0PutqSHa2reqK3UffeE+2wJ+DF
DiGGwOAA28ID8tQNtUlx+qJz9Oi6X0KQxyGfvfgHFiECCb9V3xX+RH2/V1Cfi03YdALhAEmaGm/z
vWYcU4wcaAjx4m4VyFiSo0XFuNAm/9WV2YnceVmxzZNqt+R7ORLEkmcd/bRJxovg76bpWIyuRm9t
f0Q+rN+Exox2ndbiMAkWedl0nGol/Db+cL67Zxr0DAHh5bz/RqhA71hXEyTpNXI4sbV+JQJlkQvG
qEZKa37OJaN82VCX57GPjXx8dMiy9FA2UChG+WpnZTU7g4W29otaWYaxFSYdjw4vpLdb2PATAQWA
7QxH7cSyTVoQLW+r61hPf+0GVKsZmBEzXpeJgePoMG/RpvTrxYZylP6ncF70ptF+PwcoFus3A111
PORhCsbNfH5GabjxqeSnrhMMdgwl9rJ9fzY8NkZos8EtOPzHvk+u4lF98mCUXrNuXbuQwlxL5hPw
mfmXhu9IcASP4XOkQE/xGN51WqQS7h0ERz4sfcmRZ88PKAcuA+gSxC++kxCoLkhkzrBUhM5SyHHr
VwJUpqBbDKIP4uvdkegd7yN1Cox2bQnQEkag5YAxwAwph82uAHqNjfUucqmJ9z3+kGPovpDqDoTH
GlSbLps0uywTSraP5gNiU6beyR6tiMQptNXvEknjkOz8dIneSyWi8b4bVRTnenBjPv4NbRcFF4Fl
EkTVUM30EEvfIe8XR+FTTxEMOwJvXpYSpbXsraI7hcORsr483kLAqV7hqIwnNOpxmP0awzI/yYM0
rDUa7ue8ofpXr4lcHUpUXWi5yTMH4ZeZrRcOvLLtMswufs4w9yNAb/uS8BMMb21TXNEREETrswhA
fMYK79vVnWdMhWsOt/79LlqAmFvDDtsJ7J1DHGKZbLif7BqCT0/iUWULZIdeb+Ttz+lZxTh/fCcp
m3UZGjshyMdBcxwX7SFF3YEFeqv1lYSjFXRvfO4Tu8glA3JlNob/FphcBCzrynyyi+IY24olXd8p
2HbyEfmBm3Z2yEvFXS62Fwbd3P3X09QwWscGvBakqt2CHIWjFf+ikOXElXvj7T3coIcEODevlbL0
DtQMb/IzYMUhrtg3ZPxjfDMptDHYjtou82XZWU2jX3Yd/tpSs1B5/oKsd+aoAPKxWDGG2SRdKdsq
/zNb4b+n5ISAFLrBsxe6ipeGxdX6qiNnKEwccr92M08ZXJZ9k+8p1gmxLFMceTsA7T/aBWWXPIjF
BLG4jPJ723plfpg4KJyP9FdrH9p5x3iYkYduJv+4AKICCE4OFA0QYYqk5Pu+E+c3Vt7nA6r84I0/
1Sb/Dq8wM9Rbwt6OrKSIGMJZ4V9Ctb6q9RF7Z8ydZRhrF2j7SP2Wv6r6awIQW0D5Iv8B9h73I6Wt
6eH8pCyZNkqKupnYXaW5OmEKmjS5hYjkpJvD7lPj+HQXw9JF3l7QBYiZExUk1sWUJY4jJR1md7ei
Tgdcw4ny/ci5crbirBkMPztFJDDnE+1yQNP+piOTV0j7lfq39j0fxve3ty2IsPBH7/jcVY+vhczS
x8+MqSgNZPhhFJvxFRJy5aotI+3n9HYDQK1vAzhFl/u0yNGytV4gkxBNR2hmYCstMfFYZGy5+6uS
2gjxShsU6D9VGUOzXqyFq0ffLl2/gL6lExGCrXNQwJOsfO4ziYA8pUEqUSnBP0dtd2fHjCjd2ZCU
rNXbdaO3WkjMYJHVHIiOvbJ00/0GnHXUFG8DluRjz8a4y2tyejsI6TkhliJfYz26a2rzDHUmGFbk
AUsXCHZTdnXnXh506j5PR+fR/2R2GqVFeM1ESfbEDk92RTDcZVhGqRbet0uDv4cY+yrMMMrElRgj
ZVSSgLxh76mgaSmyH98LD+Kj+k98/mrNJTeUe8EzXXEvUANrM+/cqz75h54VUluf8JpZF5UyceJ5
+18Qm0tZ+HUFrxAXwETCyZXWO8PQhbWtUm7KmaqNGwIwQvzeQ5VHO5YOzO7hrDwyCCKS5nVG9jlH
Dm2F62RF0EpYVKgfrTaNT7+xW2RffHUXfMW3ONAqSTLsGtkdi0SXVzRTrkMVFwgy9uu/l7yeL5Y6
C0GgOFmgw6aFdgoYmyhpl/YECfyC0ePFFlkjqoPwaqta9I6O94gdadRZYyKLiBAwUCe8jzOq6WoH
O5Lb52fhMPrf4vCFSXdRTQe6kYMm/JHxSBLt373xmF1I/3z7lVSs9uQuXTJYP7HkfmD4cGo2LA98
r/q/7OhAPqihy8tQmuUMhyKEqMKskYxc6jEDlbkR06/uiUBMqo9ZQrtr6QAyhnX+w7AoIRhH6rLE
kT5b5Xu1ZytdhBsFSWCcyekNooo+knjGjI7cBycLBKwYIaA/SyOHg+lO6dqIGfOEijzaX6QcQNqy
5Fo69L415fb7ep7JDXBxvXiBdesFOCWK7nWBB6RZViGU4zwcpGS7c+YTqPIvgq5QQQrjNJ10emJ2
HmtdQok3t/dsR+WKWe7KbIdwZlLyHzH41iXSz6kCxJC5x4wZXD43hGUv1dKai5ZF60tOmeysSPNK
L4p/hCHbcyiEc72N9FLR0sEyXhHVBJTYSIgCn0bdW4jpHzW5ybjM0sZPkwBs0A4bKkQU3hnUipAb
7zcVg+VW94LGqb7yz/GD75u61fiwMpszBdMKC6fEn2bG1xCTW9eEeyV0IlvKkuYvdm4pAPRzjEq0
6oOxcX4mOf1aq7F5xANTMjaq5UpAFPKwyv/IuFDjiMsEt4BJkPpCuvw1uxjM6V1k17bxHhfM1gJR
gJGQolnptIMb+7lY+IxGkChqf/Bv8drggqAZUTOLSMrbbzIpXB7dhRwnKD1MsfP0arA+7v/QqAm9
D+bLA7+s93zSPbZqZgwSIj/w/6tLDV4cqi/cNIToJSWuXUnScWS41NLsqGDk/ET550tBwCP2e8Pc
LEIsS3yNJ5u9ZgWN3mvdqmqbdYAOL/eUd09KDTo1JV3QpRgNu5vmLG5jf5dMKRKpwxzfPjB3SkYk
CuuoDxMKXw3kDH1oN2rvsGCw+I5HkJ5kAYo4rPgDTEUVcQfbKHR4keuhM8+HD4B/lSKFCguCbI1j
x0trwztQOaPtD2hgn7MIVh5q33sTwUC4F/oHsUr9l5lFY1zINP0vz9ahswApF3Wu5Uva3xElHofR
/tbS6f8hItzdBS7pmlH7KIv+jrRm2l8vIgzw3iyk+veeFXTRQOMOE85VqWKEKDRRvcffU9tKKlOU
TX6HXrbpynzusO9gSHWf1y18A8622emo9bKfbDXcvwHnLyvT382QNptH2BUhL4egULqTc/p5osYa
ipGC6xWRnrawdxb7mKdkYXVdP3VcaySkyj6qY0Ga/iMD7p75r7aOE13b8JEeUW2/FoTCCEG2/+H0
XIkDfaEWDcWIZ6pe9GkVVeMug/v2jsTis4JJsMHWj07Erlfbht0DorJ8C4p0qzNdb6gT9+DoUAWz
uhc4wKz9WqfB22vSy/Qv6wK7oqRdr+RfpS+UHooxBNbzUIkcq5S0rzp+0OzbkoouCuVRBD0csWmo
7UWKGWnymGs4fwbOxIQwn3IQDsBmbdFLM39vBPgJgXlIIOZZDOsWi02UZT0FpVG+I43SyojYE4IB
a1wQHJ/bEKuQvjvT9map2MwkKrEQQq9+5m9E96hHPF3aAwst2Vd/SZoneQHwP+v0mLevWGroxC74
06ydcIOeRSLYhVraPMFfdhiNn55EUKKbim3vxL6jA8xTg2kBHOJ1uNcqVMljsoKKr6ro/zY0f5Vz
BGS4IvEv9hhVuMho55TRZoJIygjsWYR5/cHuCArPmErWOO8xsojTfmtcXOqjvTJjQRfqNyoqrmO0
o/Hi9PMrVaN2xVDJokj0rSCH104/LVpZTgxYXsqHCXBy6lfIrbPrSu69wZe52rs3sPwTvAmDjftc
YJRn9rQNum6agNDGfgYbX7fcxR1QMRKX0E+vz0SZ5Zq2MdM0oL15ZqVitSqixiA0yKttjc7TCQ7s
Smo8I73/QYMJ+/BuZG4gQxSMsPi1UI1rhk7LbLSy8AjUikRAVAQgC1IXDdpe1AaS6oTO5IhfcRF8
gGBttv3XAWZ45PrjPqn1QgRciHomKSOjWuF+J8bEoeTjFUiuPq/NEZyI2GIxLcA1iPIqm/VrRHj4
kr5yaHRVtU+wWb/Me2d7+Zi1l7alpt/WYHLjmDEjjwKbixGNPjDzNBSrAgykC0Wqmo6QWvveRSAV
qrFJhUPHlC8FrQxjOapQM+Lm9R4YE80aH9JGxOrBaCEWy25g3iThstfgp1T1X+xf58ofmTnONBri
OASCe6o3CbWP1QaQONcrqwDgaDHwt9+4ue6lUyHdsVVkcUu6exbsgUOZC0WkKA3wqUClDKgTnib6
3jv6iPQ37vo7gcr6LSJwhVGiQR9EboaMoal8kx+vI/gqBDTPyBew9f0beQVns2advT+L6aAV1g5Z
D8k6tHJRAF2fiEYyliD0OQK0NJJvC1VxeVqg0WwYBGohboAVntZF8pizuEcUQLxB0rIEAZ9gGa0g
vq+hDRvNjLJT9vn48dCAbY63Uy4m2bNydPM2ucX+P624ur+bvlQcmGg5tX9EwNztwynpOktmrYf4
AQM9f4Uzs5/aFPORPQQ1ObBu7M8ay6HXvJUU4vhWjic6m+G60NfWWrBHdqOA2lprDwiesm9ZZvLk
aCvJNCoOCca89CzR654rNpxXRcfnsNE/phlwH+dGUpaLLNWnrO1MAVqOWfxLrS6mQDueeGKFP7EH
p2+yYUZpgFZ0vA4nbGEfB5rF4YtGHqC8VRsmNhU9fnwzBt/FWbYQvdYWKUU9gqHTFqdj3Xklku0b
JSztyTYgPY73+KLzNt6ayHbPI/sOi08zsljW9RTQvdHRafO3YTmVghvVjVr65loguY7D5pPGaN/k
/2b1fjIpSDTuILY5co/ib1SEjTc1CbaPqaZshN71MahRflqNOq5SG5NwAcuHryyMwDdF5WOKeonc
nH8VObQc+edV9EoBnZJWRo+ZRXO8WYO2B0Pr+kwpnJZCqkht5LmpdR5ciVgwXPW3XVnzjBRVI9Ev
u+Cl20O71p7F2b+jhmMg+sGwQUnTGY/SDMgVMT0Zb7J+BMRIdKVf7GYjwT5AUUHv3jQbC+lwPFFd
Nk7hbWMiDxAmd8WPvjYPYgr0HnEjxmK4GrHRenCYDJxKobyQrlF6j7Fboo4IYFB/uZgpaInxnVha
Dq640aZSI0kWQjfpbtnc9JGmQ8u0kS3MTHFa2cEsWb7nh9cyqH/MDVrB3XvTe7/KaKlAIForYuYU
LL2gKcE4+PxiUzTqbSGY6sTU7l2QjnXE2HOWjgipq/FU6QAbpb21+iF2dxIiCjcI++2FWkLyDP7i
JHlgruGP6OO5BA1Cv+CwcweklhElmNEP3glCDVERl4SFysEi/CkbzPSR5Y4on7WSL+wPVTgxravV
QhSqiHwt8nlcFSVS1xKfCYRp+ORWWc8wqjAtn7f4y7DeHDMuN8Npf6IbtgeWWn+5oxWHG8fQD1F6
BbjVXW9Hv555JC8J21icRwkOmiw3EpzqbQASjtK1m3kamoPsZo9yg2Wj8DbIO+bRn2WXsBZpOvPn
jUs0xLFTUBf/LZixoFDgM8DUngCWT9mIH1APfMurKyx+4ldh+P0HIYor/25gVQwc1186TIbCHb6G
lzj0ZS9Sk9aqAubLXpkLklUP9+xjSAGeNUtH9fMl3cezIFqA7RYz+8JmEJcKhipm7C3GSSbRpTfy
3VRrC6XV2Qz/RlToMJ3duPL9+TNLj3o4lGXWxaR5IGNR80FSmZ1/Re5st/DYoObeOybvHp7rS+hu
bg4DZPg6e6mOQ4r+EaMSs4A4ScnLuJfbUd1g087ZWSSMuGcNniVfyBxfKh+K8rlQcRipcsDIEGj/
oo6rwcL8bCV/9r7a9ofqsFJfzCeZ+OoethDVVU+afm7sVZnt7rszJHaVj+qmgtBSjV9C2e3BsuBX
/Zdn9IFjfX0S57oqDNlxlp4XnWxgZHOga4DltDO/00jmQWJ0IgJeSG/Zlo88QWgylx52LB5HO1a9
RA2b2tG4LVJvktNI8iHFhmo7clTxMm4jW5w9fmeS+Db85jIvIUesN2dMs+smdfILiSZXKnye2BjH
HhpC/rrUKqztaZb/gmvI1J+xC4v2XUxrELD1w+6i5+Czyq9BNcT7YJpo41+0bP+4+wy4l1rIa/J5
zvvA7GRWn370LfLCBciSqOUaozn24RzNNQ1cqq39zgJYdeo1rhDnl7IiiwLvyLLmvhR0YpFkhUzn
Ou+WChs4zCeNwYtm3NqXd6C2oIvWtcebaq3qg9rhEx3JInuSfknxOLcUtz5YWjE4sT+83ksxSp8q
o04pZE9h26QbvpfwEDWJYkQyAnlZvqxdzsKWT44wDCraEpIFc3xauC/fHJ2cH9dj4ilztRrHTcn/
4bn0rvj0dXFetS05S1nGwkgHuN/shmUotj8WYfavMaSXJvK4cm6hVdTDxHIqerhqQRiWq7mkz3LP
pQ5U+xuheu5OK02BtU4jUKPoxR6PchyKm1bFFcp60CV5eZF0SUkRF10xtCqV7BWg1UlIPYtVhZSA
bappN2yKT/K/LAjnYWwWPp816gAQh42d5LeI3TfA0Ya/rTTM27zVyEsXL2oPgwRVvTnzLlovkKCH
fd/q9e3n6ow8kJZtAVFyoLGliS5QaNjx+pdB2ON5Al8+Glw1CkzqF+gvpmJU3RGVk7sORYKPRUWY
OlsaswhGyCI0TFme5TsucjnQEMt/KfxazqLCHK7YVJNGSEsxWNS2EQ27ozlbNP3zpOet/NcluUjD
8WdnJ9LIR3jpTRdy2DnB774+DUn0luNcehSIA7266fdAjR93XiqJwCOQzWH1hvtYeAQpMDD1MYZK
cAT0Yen4LfEBI+y4SFNOb2q5ddUgIF2TL+/U1c2bvhZ74sQrf70j+LDBS+GScUzBwDiW6d6vxlKu
IGdKnRdSqZUJ4PSfmLNfWlpo7JR32oxxaoMXL+9Bhe6MOX2Y7qVDMhvBt+JMBYfUXRKiowm4zN+A
z5XEYCsg9hdCEUHvBBWPRSqUUp/7sOHHJrEaLZd+8hp56/gMR0n8Enf6L2iDF9GUXZzekGmJP1+g
Z9ZeqN8EoO3cESwf8kKe9ncVozfqpmsjC73W1sm6gCAONjhrA+TrCjHAa8U6zcyED9wytBzKiDS2
krtVR1FHDoHX9wVTrAxnRWTZNo8AAgn8ep3JaSEls5Y9FFpXJbbU4MIKp0hlhtAlX3M9wtg7TpMZ
S7xx3SW2qoe7H+y6dKVnCl46DTwiJuf5/vJHl54XIadqta5H6i55K4X4I8CR7sD0sx1dHkdwQS9H
vJRvxxm82/nqoYaHoYYtM1ACjLvnc2mHHlng/1+Pua1Fr4z2bT3VElRxLoVrMcyZGNwbnBS2gRGj
PQhXO+j8FJl4+j1hoYkDHWb8wAEmhCzJ3B1wrXLBkVzfP0Ie6cg4xf6BIt+/NUt0+50kQcwohRdI
ZSztxHLV10i/H1bX0bjSpNCaOQzRcSpvQ/runnWdUcuMoKHumWI4U7jsWclqWGJJbq72TOcB5Lb3
coFcAbeEr3ZuObSxllfdTlYeH3dc17UZ9c9uec6cGXF4dC37W3mnG87822Qw50/VnSOTB1e9w8zt
5gCX8Ob9EO/cc0YHftFCcivsIZPxfW9QU1PlCm+0G15TmwsU5ZkqhKxwXJWgwYhtnXRB700KfeH4
jo2Wk1VPn3KYCnADyEvDDEhLJQIfTKRcEZmewprz2FMybV6ipxFzCCNhmvS0HGRqEGuuXegUUuy5
QD+/HPIxXWghmfY1KwkxoC7kAen+8CGljAXz6W0aLw/8TgVM7ld6KbkMi0z+5r6sm3wP19l/PyRz
aDwr8LGgy23PqkQH6FMesu8ilOYUq/+0ba+1pe589LzSPHKi3FvHHgYQO8S8sj0Vh/13ycZqTn/+
gGjs2nQfhY0oWU+zrdFrstZWR+ZCuWljaUSnG25tNmR15FKk3NM0uI0ncLfOxia/1JTUPimHYbAM
uaC51YEqLe0DSFANE7Ws68ASw3BGKvJzybmk8HQanxvLIoUcFoS/2iXhYbJJqC3sebsjH+XehDOn
0vr15wZheJJkyxcJc7r61Tlw+y83yYIMWlX4lBMf1Z54z7ugOpUXrBP/936ra+JFl6yDyWMJOOta
jxiLhpDQudbqlTnSKXBFcwIMiiRApfIrh5wG3VfBda/FEM5NA7eGocZz2iv8BbpLgvfSXCj/D4cH
5+N1pdThyZuVHTdbkdwl3saD42Ux8WTZSONhBBuT8SAxl97ZI1uNoDdOM5ynFY/YMT9qkRnepCZ8
QG0jvj7lLBQi67s0usHFc1COPegGhiBmJ00/A9YZ5FIJkI7dumOkoyl+fZBfiYX8sgxr1/KPmej8
hbfYyge1TeyDfbK9T/pYw9rEzjVkM45FdAyCCm5qVkyGFEC4oE6xl/oQTzkPM+elFHU3SfeCNjOH
pGxwLNH29s1lmUmctWdGb85lxOtGXUIAivqNUxB8dvincoio242o9qsc+i3BVs3Wqpm/WzZ7Rvk3
1rh0qZ1OyQA7qtcR8Vk90vgEcz1biqhkTW6bUWv/DvkIWtRlh9qdhxEnNLYxK++DLpXvArIRvzs9
YuNCUYgUMeaFF1IDRsZSrGJTe8PPlpPKqF7S1Ui6Bi2P7TqjQLDymWJgEh2N0PBSw0ChlzMMqdiT
eI4kC+GS4pUMI9KEnR9dRYw7njlO91QEGhdgXu6sq0RQTj9KqDHZIGvcYLkzOlylKCLT/3mr7Xez
YPjXrTFtyA+kyuZKFKvaZqKWUPekJw/kwFZdo5Rq/bDJGHfiq6yE1ewUE/u2SM87v/zSA51RY8lM
Q4DjGiQRzVAwuxF20D0BT9lDtmGGvh9YEwkPfx+J6PQYGIpQOWJ8R5aNxDGLOa/O6B+QkPwOLfs2
jC+6P6OLk8W0ai3gCrYsW16gIYub4sGrgrqT5ZDzxXEowCa33xoMBD3MK9ivHewfrFmmlY26lGKe
wUtpPm2Ddy2Fi7nTaZ2YuBFh7ePm+cZIPjihoyAi6lkJC9MYAthefGF+OXZHw/KxODR2/5xJvVss
e40bmo0PKHM7iGFh7dk6kGSrjcE7x/PP0Ecud0BC0te/1+uqOQTcSsVl+cW/Wo38tZgz5VXqrlOt
ebmarauY9GJ9Dt0ixaMRnaMyAWT/iQo7JlrfjEg8ymgSegoyzNwgEsmRsBRlW1rCACUAbNPWeifQ
PPYMKGG2fwKEZutDZczMn3Ag+lLrJ3Dfk/wSLaPDp9EQFroCM4QHJlRLzPMJsgAhMUpNZ28YWuOt
/hGBQp26trL5ag7LhMnR6lD9ttCDk3oqeuM70+heW9n6IkKAm4z37uheVR79sCsuJI59MvrHNVM9
dAWxa+kOacqYE5DI9vMbE1EREHDY7SfBvgsN8lSkocQhAqmw80aKxZd6LmWRXOUoaqtsYLVzVkeI
r1PDnRhuL+w+yqmQZZ5gN2FXSftktKsJFY2Xj3ybds4qgcU4AzlVSKsmBsFiHLHoYnZLgFmuf959
4MFZPlkzVE1cTBgnQ5e72gW6FrOZFbvZ6iYhp7OoL8bQn0up4ERzJKBPjKqv+n7329EC1mXU94Yx
XSB9LajQT2NS6pPqEBetWSk3LnPZhf2++mpfpyLdZitSytt9rekcvCoJSangglJGQPyLI/4ngjSz
QlCw1S3RCJjXFNtr6gLvvWh72nd2tFnHCG7edOqHxGDJNTuAxCp5zvkQDugPRlJlLq5/MjYCb/4k
zkPqaGj5ZySgNKzoJHcnQ+7SZXFp4NwBQsU5NrqlihMyWPyDJ8qHt7BUaRyMUvN6hVTEClan0eDB
ukYNxJGW5V2Cd+Z4tGCY2dyUzSo4MkExC7ti4Ytnr3B0kmFt3viWI+vEQ2U+LCKyh/rr0W9i3XfD
8gZGZdcMRXl1j23m+7+5mvBVekLyjXf+01eOcn3f+eb3vFxLXSng9kIMmdgpxo56IXbCB8Bzf8tp
dAQWVGuZ7wioAH90O6om9faFS2XMy7zy8GHgxwICL/5z2F2EUscq0DHFkXx2AOBS9/S7BAtRTzQH
ANkIlQoms/fKS2JD3qpW0CHryl7GN0ShAXbwtpc2pnlhDivt+aZUEQGGAf2nZ40RIauVXSlz+Pru
jHlEK1pUtPYukPu4oF6ibCKEgfMeqqRRI9nXBc3Rp/9K+AEnRff4GbaW5POgJ7wNwzN61TsxvBNY
7Hi4VQECPIOcTlmIMxCN1FEZETGSycUCo3NIRAGwGw//jrVU1dstBylvGvA4McOOyPiOVNWJO54+
LzIUSjGxmhw2nOqqsRmsRcVvmx4AbsOZ1YGEW0xLYY0R2Yv8Z53Q1DUqMwxjv9GgV7+/MyARCadn
WVX8yaMFhh0Ydqqtsm5k1nU1WxouuymllCVFEVHC8ER/qioaTbZZv199Af+to5FOoQl+j4/J9Ak2
417WKhY6oUPvY1L5hdWDGRC0pCr7cPxBdyo6yQKa/he94tF7bupVxAHEb7yliasmrQsZCtG8+ClX
hU7H/Y1e7AWRw1vmPmR3hUDDdTjxOlRD02sjIwpCQgxy6RqI4yfIMYjpsCAJ3tosodoRrC/NizpC
NZRhIK3z7eKfVvnzTY3X8jbA1brqcff+tadAJD+W+Ugyl+wnNIgc5PHYRGu4x/J8gEsXsd20XpJ9
RCh8UgTfk0wGSKn2AUsoCREiyzwMr/o7e5mxXFcI5D04uIqMm3t5IfdslgtGwREfoB4PSzhBHGPD
lx4FknSjCKOki53k+KH9A2N8QREMu85WOZYNqlIftYwRsgiWgqcV9aaqNVmK1I+6Q6EzHnO3VS0L
vhFGofzcPIMsCLe+bDO+lPkfE5V50ZWE1fT/W1vbg5SqwTQt8xoPV8W8YryYLzUYOw3WarW3JV9D
SDYaWG4pdA+KSOV7AQCzlaKZjB06zhGrMQUe1JHeJ2/8tUihF0i4BtR7ZRGkcGnBKJMMe2M2pu6M
3ud4TUbia90YkBM1GfrY8oWeCFveb8eO0gXga6dwng5LfKbyMF/gI8wA2X3PPoJ8sGt3PLPgNi11
NaVUxCrcD7dFwAffUf7uEqF4cksHiJkReOtJn2k7v8ifCr7v8NTUxnwfAkuf3joLKjxX2GiXdh+G
bzRrGDxkvwc8uSbacw7BVl7wkWubSjTLKPYziv+2xzCP1H/OCFmGUCHRQf0uSSImt7vM+5W5CzAL
AEFhAZGrzoeH7foTLnby1gCqixlGPJNlNH6vflXzSKEQHkg4pV9Z+f0WEci3F8jI2n1JSsVVnMkw
ejn8K+ti8ybtD4ILOhbDa21aLolcqbOV0+0EPhEKtRS9MjLMXxDD22WWMTwdZ65CuiHxxvCNK8pf
2rQvUL13+UqH+bB0rqD5FZYXaAzXuwSLWPF90k2zPNQnjObiJFSjivOGE1v3AaFBEHIGyD7TK9b0
SoLPNQA3OGuPQTpOZh8lzQRwdvvfC3iWsBTuNLjjqtVdkfwMIAfOMC4sbChdgGlUxNJnqhLsnQLZ
aArRSvLqYFF4TfRibvF3fFcOOyR/I/3ZBDS9OBmYGiY7x9GWJPNIgq9L9/CwZHsTwWPjd2TlsJCs
hh3epM9GPh+1uN/PlikVzBIZ5SIFo4WVl5xVQjY168SmQr3mIRUsVC0F/Gjsy9TI9ppDIZcgXtJ7
nq4vhd0VirmD6BJwwuhcJK/MnCWYdXwVz23SmSvbit8QC+ZI0flSA91Cqxbwdki5YNVQCV7SPTdP
ldLQB4M2dDdoibHWXiNznvcWpP8P2JlCIyrMWX4K5edgiac/44B87l+iStngJLJMwlCV5t2xqEiX
zA5g2jagSiS7XJcotkjN0lFCr/1y5PDChrPcB6D6PNB/PGGXARUHv0osWXKvzfdJEP+AJHvVGG5k
WxOVfcJi33izxYQf1ymUe2tZkfV22pcOvNRw1fiT66rPGGMTig16daeQ/Ak/pdhPN0wVuhZKncqQ
6YuOiqStcnnf0AnXe8kxgd69trhj+i/MMcKvysoIR05H/ANcdhLVDPndrlbiReipsfWs9VQGYgEQ
ARzhJmK1Ivigl0FpfrrhOZ087Rw+fRbNBTtPXHcw42WWcOi7gybcFQ9MP5xOBvu4AbG8GN2Azaab
NLvQ9bok9f3VVGAJ/GRKZBx2FuiRDbllimZUFEjs2W7XkhbkrZ6EjNi6YeJlM+G2jQnuw9aueBAI
wsfFFglDRWHknvxWoIdnBkeT3YHYlGRAY980tJRYedzvoMpPETOjAUI+BOD4wrOaQ6o+t+raRnDl
S32cEY5ww4Pukm9P1O601EEG0ZjOCPMZbqWCSxE43Aal9iF66CYEzap9hLb6c08XRIjqieYHgfrj
/HTVqVsMXt/cPHWB7E4n87OcZMkQbdAx+T1O8CahxqpfYK4c61FgZ/MNa8NGQ+qj5/g5dRCfkomb
l8OVlSSzAYrpBcvgA1KwaU5EWOpaaIVs/9RbWEUNZElHsrLsFapxVT6rGLbeF/XLH73UF/RDPTPV
KIZA/XyBkJJ21CzJvQmy4F4XadLqSUVEpalIlzaSHls3DV194mnaGjgGwnjAl1mwu/4M/YJ00ncQ
mwV6OU/s2arap1aOhlb55XPOd2Ltz86ztZZ+9ed40clfNUt0V68tgC+i+zx0a7LDa0aR52+H+D+G
LlZ4utjZzMZpMU2XLDsatniAqqAzgOdSgSg1yI6XTFTST9e2xo5DSIF0xHZzZbpkI1bP/cURUA4X
P9tRhP2hSheAiQSwzkCXdJx6LRL6gjB0HYtguQqWxgQM/RosopovcigY30PnIQlsI09ksfoHDfKO
zceuPjypU2Fh3i7WJqrKxjLkGnC6GaK7EnhTm2ItjWHYwu+3+PE4ce9kjU0Rj5nZy23rJaSUDlLA
ZqAgK0eFADjxkcu13YcckAgSsDKw611fW3X0Atxbem5b0NduAm1rIoIle7OSW+Kl6+XPSRcDTk42
5HRB+fjG0rGr3wM8UlMbQuVTubIth3V6nvvF0R86VyoSO5elD9GkUn/zp7tw05R3rTyOwI7KqZ69
QhFPIt85slBKfqROigot2CaZDxg+hsZoJk23Lk5a1Ys66lw02NO3FCQubfQez6maf3brZxhk9FYN
kbLIKnF5xZX5yyTi+5bwt77nGsN2nXdhWa/kCAqdDOd2ZZQVmdiF7bmEyOjp/V5gewwGIjeMzlvc
XaCu5cDZC1t/DwiTTQP0TNBUJW47pS9uD6KKL8YxdGTKls4jQaHN6lv/RWatxgQoqkiOMmP2yXZ5
+BwKiAH4ifERd/CNCvANTpsaiYx3SMcAH7nkznuGLoeHBsFEaWGE0stIV9Xvc8EnW3UzEoXBI4up
bpJ1HDKSFVynTQfYF8qtu6vRVxgAK3scjbhDnDGiq9GdC4j+apahf1boBKZb9JPQcp+bQJqlf2fV
Bq8A8KE9ogq7DuDQCIe3odiPK3BHDaahYAX/9UgzA2SuAyVFeDeAEsV0BG/b7mY4bF3v+Uf8+rWg
dOYFGM5r4If8JCkGam87C5wW1S7+5cyX2l4sr682n/k2KkFkAzn8ie/TJMN/Hsu37P9pyXLf0fHQ
3HcqgGyV97Sho2Pwr1LgA7vKB7aIlaO5kOQlVn5AJ7FwABWDoFR5L4TdsymSZoXcQV90Ik8Ryfq5
cjETV57Y2RaM7usV02sqZBHW5B7FR+k2yzSJJ9Y8vuJzwW/jU6vZLhHcG1cYwp8/b2ESNWLhZ+9O
PS2jUVE6xZE84v5mvhhd42lhd/EBujsGTd6GBdcxNmGlxywXQ7+sYR+XJOyUOmXNhe9wFknAhWFR
85SVkhok7EP72aaAbA3BIBs8DRHfwfM/Oez+dAhGsHBzyf1BEvTGE0IhQrrwU5hlxKLPzgx+9voj
yDL4/Z2OeBDxcGvJQKXnfjTYIXOBNoE0/BW9ImQO/3f+Zs5YExqW7Fwn19s9C1DVDmrSj6I4gq1M
au+7nmq8j15ASBghpH6+JWuFnwsfiZdqiYdZGHFY9izsSSTsVDCMJFHt52sXw96nt6aDR4Jlq9S9
oI1AB9qLzDVD3RyOTsJQC3MH8LCINmZCJ48mCf6+w7LqixxkgRenHM0Jd+uZ+zziJIBQDLcyOfJL
uH7aEi7ECjMZpsJEi75ZcOhaQILsHDiwnSEf4BA0o6i/bOx5shZjvDDceKQqquye+2lK50zRwhAe
RRChimD3GBXb4Lt91av8B4S5z6OasGqjzNKY0FwabpZpAgc+HXUI3Uw1WyHQoPx1i0cVaFB9rmiG
6aX3OOoJA3QTbNp39//mdmEOnCpaThsVFJ5xiQD1KUJYccVQbewwIrbec7HuACE2p0gJmLsTku+d
hq62wJWDRnTgHD2hxUUNbe63BwZk8u2QoOy9pbZvTJlnQIDc8Mu4hGym6uMarMULgaIU8KRjJbXF
Z8LNy9lttts21U8PHKYkUReF5ZPeTLa/UGp+m0CAt25hvl+cfNyK0q/AQdApqbauceXowD5xdFMq
P2+eEoERFjg2cgsROOxTiuxZWcPJq1wD28CYAEQcP1TXUFRWp6w4xyw6K2k+KHduAIuWVJGUiQGj
JOzj9nONN6lqudQYPyR0fF8VpiimecoWZLFwyEFvLWyQYFlqBz7+WhnFocW237D8W6PGjaC0QnY5
mrF/YV+rI7uapfIIhsv8V08bW/WbiMAz+cZMytQYgFFiHhG9yuZSq2t2DIugCnPKOv+8dYyCQX7A
/DKvr01XtideyeuRAETk02uuHFPdsj94CIT2/pTlgatkHyCbpfGS3ibCqlwjFAz4zbP2n/QuOoz4
JTue94qSla3YAsXlxemsk3TPYTnAVC2LGZyQ5OepgvD7wQBucaHF+HP92KWQCxckcesSiagYSlzk
HdJmMZCUa7zl9sZZ/CCRceC+qk8h9/SyBVsV+EHZywGY2G8Fqn6WMFaFGkbZowNeLq8n6HoqyXPe
jninS87i9hPLoMxlTI6JYRDxAMcqTJN+cMvFBmjCN5wKfgGUJdRknWEWEdwrTdmKuMqQsBk5Lr4r
cQpdQYs0kQ3szZd+CgsdzVwOUCZO5h8oMeYAJX4ZespukmsoAxhm3sbfm1zZ+jXlVRNniyZQl3f3
9herUnwfCQ+Wv4o3Lb4sciIgotHehHofdLpjJpoRm7GEO5WqCFb6QnDQ6y+Hc6PRdqtdHnbE80AQ
SbGjVbh9fUglnrP+MpUMYxxvzPzlwy//k6u/wjEXoywayXZ525FLWwXE7BUGgnuwwEOiV6BnIyL/
Fp/yFZ9GX+J0bA6/16028rikoJaHx0f6ffvS45ZZNXkPrW5hL354Y8w6i+EXth5AcQG5mdy2ULKE
7XPyGwlXC3774uAABoo0oNR9Q18UD2gHw9ZxDXlaX01Vinvwkbb8nJxuo3MMBACyiQNCEo0G0ksi
0ArkuyhgbsNDWxU2xuIVw2nlmuGpK3knq4HuI9Aa6DdoeglSSZLDkcgIATOtyFFqSf6wrq256k8P
fdLLXJJMONUePAaEQce9vBotzjV4nde0aNDdEJWgherXNqj0eVsUE1ubCcQeOC/4SqAZsq3B+N0X
tDHdnIauKCA/plpjDFDhx2yCxUVdRQmi0tL2mLWkmOWYN3FOA3m1jXmU+XW21fRoe9pii5PRodIP
JGqBDIetqHGMCCwijAbfH+BTWIbNXQ0yj5aNlP0ETCdzgwbdCv9X4pDGpnh0VHs3IyX/mWfgexI/
R6FudocOYbZeD36dv3HN86BAppmkqoACFgBOMg9Nsu5biqHRWUDHGgC/88BHfKX5oaUBFMqGQBRA
5fMaRep27spF7S3CoR2uqJfruG1w17o55jC/stZivVo+H8hmS4Ml8Hhpz+8YGoYPKVdgoFfFJBnv
Nb6yzcuCDbvPptcolavlO3CzSIJx3BULYNxAdiawRIsgo8Y+/RGaO+CUZAuEtfPEd2rmA/6PVMCs
0Sv6lh60+zAMjyf1vOybyU19l5qYOm3vo4/iHolL8BcWW6qn4dJ9yFRoyvMUDOV4+FhiWGQZzK46
sspH9AAHKPFCRI+rIcoDg/PgcYzghfpbbhTze115wSVEEDAANXYm5kVtymaThGTTzh3cYHbgkWdP
dgU0Hcd0MPKP3CO9/4cvds0IbEmZgyugj7GG1JTZEHcUDtqeDm5A6jDqbhOnv+KHUZWm9VH0aBMB
c4jk1uFWsrIpFDhjwUZOKF2v0QuYpHUo64lVuLHj3tSk329NjF1wz16C1FuWzOQjVI4TSpuLz1vm
v58Wz4YLK6UwSWSVgvBQznu8ZMapA86yZCyx+sWPmgHvg7Pior9NxpuPWl7PQB53JkMybWotRBY8
xKKm/2sxHVDxlKEIMcFTjp+XUP8sD56ODdfuEYOKVGE0qEBRfgJTfJdu8reoJiwtzgfsgpzyjir9
lT6gm9lpRPQ0gn+jsC+yhNaXStxAiJY57q4z7zhT15XJBD0GDGpgZETUGa50Nsuansp/c1souAS3
B/JfM2+EKCLBR3IR9zKQpH1+dWy+ASHhOCRYWD8hVnB+kZtw4wqLg8F85+RAVOsfb2pt/jZlfjZM
N7wQMU/PMvoXS7HOnSv/y/TWoIL6+FFvHPke6mD7oc1Mu3zhzPVb76HWkCQ+nmXl09joKcDRV7aL
/4JdBvBYC9YWT4Pig/YNpUFdjpzwU5bqKjVomyVdV3bce5bj0VCefNeG5R8Cz742nw7P2U2wMAas
CrlBMmf1D0aIev9d/tiiqM7wQsqyK0px/zMZgGdYxGcddO7kVvxD55U4UHds9QxgrfJa9LohXdey
8JYnfwv0JqgwO6vMoE1aVce4GvMxs9OjezQjLtBnKXQpAiB9bm90PiyXen8+lWYxAdxL8XQmfpdI
AdIVWZRDH49RcI88j1Q0j06H895/50KLbDOrm6iCyk+bAnbalM+Iyg8ZMuwL1eqKY5jVKTFFSN6w
i9xVXFaYMp8vetsTtZbnRmrg/T1n3gdw3EvsAI7cHy8SuqvTqLuuyVene6KE30pEWrK8X4aA3sTd
dZlZ/zHiUAyg71InHkM88zgGrqH9cKxcZb8tA97K14i1yEmH7b2tBAjS+j0SWolhApGnnZmUKU4a
5tLGSW/4izTPC4MB8qETMoOKndKHrmE5V3PgUU0uPmO7PgCBBe9H+hTCSLPXwk/65AE1QK5NtcEL
PpMnTFvD4hWuloPvTFB5XMSeQYuKnLMKNnIoUAy2SExjocrS8L6G3fG9ALkffiyWxFNa/veNV1On
VJ/5MjQ0kwEjm0phBkBw8tzYHAB/G9Iqeginmi+5dHVTOHmPrdlxsUAbso2FdJoUVb/6iJuszuTC
VznvZB05K+aI1D3pis9ZeYFcEdB81t+t7y6jaS6Bts/wVuyHeImI27XFcj9l/fi3SKCMBxpuhMP7
eesDjS+2leJxlMIfhP2YI4MQVETg+cdPqkRvBAVVqPLmwCcVW1Ro3QVckDkK75IWownHPoQwHkbN
O7fLef7wvrQp5TabU9dIz+c+oAip3HLHDvfKzSjGuZJPOixn+wYX6JFveET7IIe/KCKP+af7l0uW
jLxNe7w6L7HwWYZjOAolcocW24W+9lsU4ZPW4Su44V1fcBzIup01PP8T0DTwQvtv8JAOxeYWR8t6
qvY3dgwxB7AVBV1bFyBOvV6gZv7ZRj802B3DFa77uYpqa/fNtOc3R1VUSBQLmq5bzBCi3glCSwAd
Ord96EmlWU+ZmcPfOtcW++19w6+UTX5Tzz+fwCK5X/H4asbryXxWH9SzrFSl7incmpW7Wq5QuQQo
vly5g9SHlprX+Nk8Q1chcSRHHyU6Fq2Yu2IRRt2nwsfh47sbYGkozz9p66CI7pDIORaNbGwKFDIV
wpdcQdzD5TUaKWnIFu2w3Sa9yBUhFj68YzEggEFqWLnVUVqEMGnqVu+jZ3sTcL+XeRtdjq3oRHi7
tLMW2oJ1ecG7rG8AbDfO8fIGMr+xENaLmZ5/hJAlOVDmzp8yZW2rd3fAJlzThWS6jmPlowJXsiSD
s8+1c3ZJFo3vDAvdrMbOm2jBMoVYyT7D7VYSb/RmEkOJqynvB8q9pKoZQQyaGn0lYPHYr3XgvYIs
LA+K8JJiNUgzCA5bdfr1O3ZQvxPm+s9tIoVmQSmPX/toVwadaKJ9ZjGHSrHftrwRHLRzCuNMWBDb
fsY9YqaEBrH/oxFzh6FIxaPcuTrUchaF7RRIvmxb0N4MVHKa7KpRGOD8BgOWtISwRedsX3yc8Vyj
maWdG21cVrZ7dPIYMYEM6D0tSHDIsqJRkZwww1/OOm3RKkOteH+PXsIiakz2IzOB3fqJF0s8pITB
wPBPTgTWOd4QJ9T/rM2FkVFu0Dalt4W3wA+dsTVjmjjnFkD5pIE+m+GqsWD5KCxdlYH6xejoUITm
yF0YjbbZFPMvWzvaIJlMBNvntqnIsY7n5O34y1dANRf9hdPHR6nk+jv/oI1JyjF7+mffDjr74BNU
9+iRyHPv11wX2Ni0akpURCE0H+vbfbJMZ8QOj3t7gS1s7Rp79ng9l6tOJj9uxegSKoWVfzOQBxrP
xf4orAQkReXppOqEytrZ2z/WzxMyWPC5LnSSYm4jeuCyPiGFsiRpQsZCh6FiF9EEnz3ezlEFVC0j
6hnVlKS48uzUb5fKqY7+jnC1KX5UKJhdTSdP5k6WT0203fbW5mLCg/GVmjlHcr2nZfgQuauaEm98
KJAzDlGok2Yigfj8iCPlfnUNMHA3sgdPdDnvgTvadQpwk4HFTVaNfwEgT77Mhlg7QWLC1BoUxEy+
hwqeOPKA8lnkECgThlviUxQJcyzOmRG/ZUFezGG0G1dFnhClkcH8O+3yIQODbHQhYJuBU78c6ccl
KkNskcHZgFv6v69/hdjuw1XWB5NMuvy18Bm48d1FG9B6rSlRpiiuVg86SQKGX+TLVz/7TM0imks7
l9dodgG76XnkyL62qccolB81UOAEaL5EmSzUezp6x243irbgy5jQ7cWssUJFDT+Kn4/ngYh/3PUw
WT4IapS1HthSwn6GRSY4UlZKm63IHIzz0TE1xTPpgaWHP77OADWk+ZQs4QP7be5PozwSJ/dFuncT
8Lfhk7EcTRtOVucXZRMIWLzX8E6XBBa89kUVEvz8tXPpG+V7/MFhLEX5f7vAPyrGtxgd0ypgvGCN
54MjVG42SJLahuW6q4rWE92ZAq3lvRd9CnfxJXlTUAZKf/7u29IUBn2MSc5dVw4lL5iu3Rehisao
hKktZiluTMXMb36wh1Ekf1it1zC8SFW0hUUv0AWP3BTsJ7xCL+NVy026ee2Om5vzlhGi3vssCdom
cHkSMtvKuWdws71pATx0833JrlnPg610a0jjy/1wWhpI0nzvKy/kvrgPDWn4aL1snUK245g3xde9
WUhqOBY2GAhkLoFMwM87chfDFInuVh/cDEToDt8CmA/RumjnTH8aN10KyPVP7NVz8OfHeypgu1xe
Gc9tmTT80xckp5IF3NAzOLr5Ke8RboOee1wX+fgQfXnAbF/2CGLenAI9vWiSiWXZMAyjGegIcZrW
HDyH5v/U3E4DrzYjOULk5piSXWMAYejFrPsPKsNuBmnol2I/EddP3GhNovy9bccDDQHBcVG8bZy7
O0hgauDakZrCmPlV+YfLnPkBfuqrw/uPAaWSVB8Du0zAlQYV0kzn2aRD4G7u3hgvw/DiOybmzZmN
i8ryMHvvq/z78IxbsfUv5JtlXcGECFrSG3ZljTXbeg32WS0MO/7r6XyR9UbJHf4vjCnUSA9Nqn+q
OxmvIJzukutZgQu1XfgVInTAXtwGr4stnlPsNCRhPLSDYpD9L9bqUW2NmQ/Hthfs6A+eQEv2VabC
m6njKOLBgsqrmYojsDzdGFRPB9R8RtA8bY/YMlNx5EPL94XRoaLM0K/F7as6UfL7028/U3IMClXt
ebOc59nac+h9NmrSjDLHgH/uQ4JfsE1M5tu2mhSelXtwnngdT98KdZM+PuIoggDeu7Qx4Ws6/KmS
mF3/ZOph5PnaTZ7fjbAVja5NaQrucorcHcFn/8HLpGKABLniavLh0HZyf1E2qDE8w5Kay8i6BM0f
wljlFh01RckKbn8e+GoBDb0484ndzyhI6KZgBM+Q
`protect end_protected
