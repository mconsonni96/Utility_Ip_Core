`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
s4IkugzpiA7YbJa/Gvj8mF4lf5G2DKAKv7AOThTYK4BmsRCBbMFxkIrzKGt7gOZxQVQ9Zs22o3Qt
t1OYxI6tM5tqiXH8SOHzOGiEDErIY8my/xMLu8rLua4LiikvZCwVM+KMHQHuFWwEOKw98SkbsmDX
akQO7HIBO3bacgILdJKS+xuIy5iMzEfwz+u7ObOSdAHI9xwsLqhsL/11FB/m/IPXMDGD6CsA5GMM
1PFfZfNCDFq+DousdnB7HpmIVZdkyuYzlAtFYjAfWMYtrYuDN0En2AgIMqg805TrR0EHBssJ9Kfv
iJpkiojOFT5t1c5FOZFZ/XltLqks2NCK7sSC2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="AocdVr2byY25L5s/GqR0yJkU5xGXFesVxVFAO5N9es8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13184)
`protect data_block
ulRk4nTmeZNXy3tXSEz36xPAAKXmjk6xUH2lwa4Aigr740echtgL54Y949VNI+GkZD0pxSIZ72Ns
tgq+kuxR949rEFRX1GMfUNQ8P+Hg2y0gWuQUNRbXk2Kl47uMA7bEx11nH7GG1nsrkMVQkxYx0B+O
1mHM9UtGIPuLFuMBfvJCiPHzy4eeSt/jr4m6IxJeLXYaIURvuvGcEg/ztqBSl05MLhQD0xA1VyBd
LENZevrTn7p8e6wwh80BUT8mcVZIVUtcDPc+MR0/Ta8o8zWPactfJHy1wXZah4hsvZAWonvrlqsl
0EKIBpF7hcynIzZtqnZypfRNS5s6WS4CF05aMHuUxRIJBYoMSJ+j5A05t4l1mBXbayTK+LSNRQoU
ubPHpKonbNNQCUj+KS7LPcF4/H/u3PORTFofqEqmsnB30fOB1HH6EHwbKQNHgNp7c19JlsDrCh9T
YwtsgBELUaeGL/RrVgBFyK/qtuof2uxt0VWUX7h2niDXyt5mskfKcF2HjRQYpk+fQY75Yh2tGqR2
5F0hnfyqx7QnfAzDiKMIGM1EuloiGdxhkSL9VHV/T7YvBPtejoomPE/WAFnEgPQfLq+BZ59srFbd
79iAQp/NgUxICOBnL4ugLBKlHTpEbF5QQmc9YW1BlwnPbq0W+JAkczVYu8LgCoTNRM9Zef/TYe0P
x9nES/NH5O1u2j5Ul6ojtjCGEoatbZ75MhfJlVpn+vf6gqvee8PPqHPpt7mdpk4eJW3ZzXOFsYBK
94xoIpAs5lsCZ2memSccutlyTk1MO5j8Hj4/Ydx1RJw7xNhoUDMJgk/a4Ekn36RD4I5kQ/lBP6QV
qsxBMe588ukGNgnhh61BYiM6GdC0AAgtJzIb2N++9ffafsHM9x4Wzk7t47gok5JFLjOzceN8v+1P
4rkw2jucam3tTKeKQddW5wWVfTcMg/muf9KpPUH5PIocV85gaYnVahE4aYlJObA2/Q5B1tnj/qQi
2DDtCRDDVgypRwO9729Q/7A1VSd5RaQkkiWUPiZQwcBWTCq7N/wNpx33FCVti+ixU1Ah7P0SdeID
GKPokMOv5RdKoXqbajtX2h2x3BWkBkwfS4dT/fl37AZfl5tMTKJKbUb87tMwzr8Yy7bMUWRoXoPv
x2BB/AwBSXmEeHZJ0dgoAXKCT/r/9Kb4Cmdm0xNwjYypzwt2bY/4czrC4w0AigHt4HN4uKOSh9T0
1pxmq7Wq/BX1ZzeSGcOR4D8UlN8DBUo0To6SBvm/zfD1joHKPRyRX0uN/kqQL/v1pttF9V4eqLVj
hV3I9g3IK8Tfd4OeGv/nBSseUEj/Od9gkxAYF98zYqFYid8X9Bxy8j0sIEZF1ktDiZBW8GdULxKN
iwuqyZmx+79DPgODTxNh3GK67IhI0AjaoihxXrom00zf7RiRpOhhCWLI5oHB/mYbNschqKq7hNeY
cWvhvRKnYQGAzThmURKvIpKM6HT9XHKWMtsNW7OV9gppY2xY1c+/JVBPmgMfG2TS7WDc8nILV8wf
HaL6gLCs7TfJpTx1tDLQiAJTaUpuqf0ogD4b2KJmq7HlAVV/zod/rtIgc95fylkRv+KpojTA4syh
CuRhT+R+bh9uObcebnMvJKwpCAMrSyIaZJ6X0UmUc53haBST6NQ2SdQFAwzPUvY6i1zaTDyouGzW
uZQYbgMd0xL0Ktozh5DrqMVQEIAfsevUJUIkETwHHLUleFRPPZfu2T3v8SEl5Z8A3h1HC9x0yb1X
lnxBNgjbHp2DIleR1Yl0V0wdLpGWFAX34kA41a4fi4aI43lP8JSZBXL1Ww6zGSb3mO6eHgJ9RIU5
WmY4vv3XexfeCW/R/H4y4JEZJLfxgVAlUgOuYg2JpcGtQVTm5eQKu3teEJ359HFRCPU7fthi6A+k
116nZhEoy7rCfhcqPzRF6Jztw19g74X4GCge51WpiHdk/SbvhkMJGsVEj2aytg7xc0fdJyyyHKDp
2ZyacXGHeEreHeHfwXS/Q64pQQpAa4hKXb8bSj3iQHj6ekfQNbFOI42Of0p7Z3A84RLT7MDduZbf
HQLXQf6Pqg9A8f5G6FhIG/a33YMdlnVpRe7/N7oMQJ8LZfHTCAVZ6CTpiUVTEt9A4CfsYo84PQJP
8oGFe6UIe56GctR2qyYAKB+WrY91en8kOzG6u3uXbJpacBjKEOKBFqMIQbDAhd25g5XcS9Au7v7G
12qM+uX//UKhBQpGmuz97PAyDSgdOcZpVYRE3sASUcuTI0vQDMKNX7NzL6/4MlGtlQrgNxJ6eMm1
GHXMaWg+57YL1DNd/Mxj9u2M5wXKC4Mf6JeLrJZDo2TsHhRVUm2hrMNyeP8yxCZ/OtjF3mN+TD0r
NuI4Eb0l65b9vMzJOb0CL5VUUO7HbgClJSTyaHg74SefgZMlxnqBy4+MDpeAnRpuISh2MpKdKsaH
iq7C/daig5MLEg7JlhYF+ukyNWpA7PaRW/ksnMOC//NdSnYvpWx67VVOulEF8dKwiBkp+vClsTkT
1cOu51px52UIzGtSG9JUw6clum6/7SJ0cvnj81xG9df2fasN2fMxC27ygodFu9JWsxZCxA/6/WYg
Pw4QElEtlZUNr6FGY3hUV4dJGUTuz6qNVPv0OBwExfwSJYYYEwr5AbX0oNlJ9gLjdS7BEUjiR3Qz
HXwm9ppXgbgMrFm126Uxr9uEu2ndZ4lR0Ysvmh8t+BRdCk/JzkK4DPQntRS8jZwIOwFlHiKYSOQB
a3ZPLON/IqYEdSeP6odjajwQywgX3C7NoK0Yy4t6aHzzlCBqLECnSozHKjw9bMZ7Ym0OJ1dUuOrq
vj8lPZQ1tYl+oGfN24nvvG2SMbSKNCEM/SB7P0PMqp9CzmVVmWMSNUyLN2jIN/8r3TkxSSfvp/CT
/1nM6zg7LdJLQlOt5j2JZ3u7/Vy2e8yxarsIJvsqO5wEyI2M3X01x/8Cr16l/X2Vudiv3HQ5JxVe
qWwUlvKKHd1an8IU9yzRfiWF05xe4eipWf0M9L8shQpgwZtAtMy1UTigdFM7CoY3TCeLkBnQITIZ
KaKTizUIoXEbAFHMe2asp5L/C61oVLPurgXY8/5qyC7Efh8oka5CQ9NwYZhx74QwLdSO2k8TMMIr
VG/wP/s9tgfx5p78q/v3MxprZJ3iYg2Ydw2OP7C9wIZkrWlu3olT8DpA//qStUoOVUcu9WrIruZK
IFl45sECvTPEq7vXNvU2Gv/JZuf+eZQJc7RwhBHoejTEBOkLnRdFgHSQpr348anMUPJDbwabkgds
n2KbXOzUeNP4bjEESn5Ct89fTuTqCzUYfF3KRa39vHpOmd+4uhQELDp80qDVxJIDH4LXqIzLKcDZ
N6GNc/nSQhfWzGsp7ptatoCMc4MtvQZByRdmejOPdobnVASbovh6XdnAZ1hZ3gplZi9hobn8Bgqv
l83Eie1DqXLeg8QlNRcdLAsK8VXUEPJeMJGHQdhihNqnVWKjpeIBRSflR38rQ8SZx1IBPgwMO+yc
9/seV0bB1l5iwb3HOHQCj1S8ZxjI+mJV0DG8aRnQe94/kY49eALTDkedOswY/3ZigVedF5Zu+UTS
EriEd6QLbY7cjpU1eIbrfh38qaj7xyJsTCNutD+40YCvqdTg6eGAEJPn+0GtpnuBvInfH5CKiMzc
xdjJ6F/+csdmF9fvC4YicE9XGAASlzagRO+IrUa7zLku7kWZg17nRAiCgnMxCOvc+bYl8kz2i7li
4COChJd+dpBJZr/NWgufkKczrdtgPXwg7QIBT1ERC9NwDUJI+YeYj/PoRdPua7K3m9ueap6UZt8r
gfnip6vxZNlun+paOBru7k8/TcQAMbH27oyrdKKokisJfOnH95m8H6Yc9gfB0Q27OVdwzuxFWuOf
m4vKW6iQ7zqsOMowa2pUYtGzxHQdMbgjO4kuUqLVtKfavNIrY7HUcp8eMPc/A4oIr0NviUN1cxxp
02FF50K0iLunADqHKms4w5Ong756Ssj9GtMN+px9ElpynxKJj6hh6tVUYdf2DqEQiAlATcAhMhiX
RLjuJtf4wPJ8TvD60CifP1IZhKFgRaeVKdtg6OKLPZA4T43aCngLHvJSyTmn7lSQat8cl8rYF1l/
R4QROzFCqnGjpDH75PhnpikwDMI8FYbtugNgSErNo2SYe7h+VKOzTOAKDpO4FKvOkqlMimZFKksJ
7qsPXZiaytdrrj7O8M8djNfSAgCYAgc2WqARgkBEQ1SKuwkH4pQsNsnrCbj91hBbHJy3Yzpa7rmp
2qiOOG5W+QCN55EDfW0vnOpVLV84tFdmMseOw37irhaBCV/DLHG/L4pwYdT6IRrjJ7caEDZOHDbP
qfZ2o+zPOmg6sVTUoXmWcEwVNkpJx6jeGzFWU7ny7Tp2u803JhCjwyH/MT9PGDGJS2XJiFlphP54
XxI9SD5Ew7ATLHntY8fZ0yeW5XebGvRU/1/Q1+SkP+zj15dyXvgzd5lH05/mCeGdH6nj2FLkrhqZ
Evcn9ZtCtoz4s6vbFWMCPvbO7xpVKYTK8oewzPcmuBanL2dbgvhHZWkhj/L7qGNTq5IpDeDOPFwq
zbGlBW3TcZcpmnmaQKQw9XYXgl859COqQQUdehhATvp03J//ptjJKPXCQtghXdOywFycWcSxOJlT
3ONeFvY0B8jkw6vfO3nH7BedlM134An29Lw03ZLtTZCibyElKLCbf1VTcghKlAXJGboBNQFPXNcf
wCfJHW4mgFH6OSr7OOTkgetlA1HBqCV2MYD1NLn1weX70LGOO6scDwbFlcJV4Z9tCjpNX5zgwFMs
++eru7pbQlDvgGo7MkjAb4W0zcdVznk5oq8sBciedyC/iV8B14D79eZC8IsBCcjG7ZXOgbKVoIVo
8WNQ/lu/je6ERDH7FYh1sk/MG5YyY5AY6473k3ht0bbruKtVJc9rvhGSXe45oEn+1HWV/4kxV5L/
ZOiP098w+bVSXzwK8Oaxq3is7I06c1wh1hRijhbc/nTTtAXGKa7o2jRX+yRW7RkSGVTD9fF7lYPi
nkSQQFhOMbtKlo88P9fx4SQ7yKdb8g6NBNRCqfFfNb8tQNymbC77MOp4ZN5ajZySdHxjvRnF0lwM
UAx5QE0lpTPmo0tGo7pMxTuTlYEQ6oCLImNHZm5Rp7pR9+aCbtf+8wdQeHERSehMYw+S7uK0I2kD
OoeDQtA9L6gs34A3YP58nnq7gJlKMipHa44w9PNyfBU/Fi+wQVCVdkMu9jukkGKx04VjWpISV3O8
GC/zCoQi/r8UGhHLKAAKltx0M381ydSU0qM115XNlHSHLPNy46G4xD2U1C2RJVpRJtvQ/iAI7jv1
BC2bzzrbNSIrFx06R1j2r8tpiidIrYZ79TOFgHyMTZl9sHokrbrmxJkdlgFUHVZ7QDmr5qW94SNU
ve6vEZ1ytaTbUI0pBG/wkVV+oDM25IDcs4d1gARmOs0WrIf4jq+A4KgW1qD2AY/VHBdnszez70PF
cu4bb7O9qQiOf4SBnqXTxbn7zLodgS+C1waFd1ZPKiiNWZjqotR+trVd1r/EkIzvR+IVppTsqctI
aCmYztYjByoCCLArLpdXaMr7akca+qxLKJ46VYTmhIA6+7VzE5gmPvirBz7BHdqzGHjqP4K0GlML
SYKcQsDHdCqLOmP8B2fVRTFFtSaEAUVDsUPDWufFbHf8dhB+hrXfWxx7s/pfeUc06F/BaZy0Ywui
DOJSQ1lFeEcVsVlN9I0M0HrAtXmI2eSHXrRVVcEbvxPe+8Rd+exxBmWUwiL7N8JTZCBhrB8NQbYp
za1fb6zV6EETtGaBqXqHG5kl6sA5e+2jMJfSpEq1WYz+I8px/uGoSsEuOqly1+PRma+CdNFrfEqi
j478kNwLARct1tOynZ5g2SBY9QKuERQyiGiz2iZKzsJU6d2/cSPhrvQXUnuEzGe+SjekygDug7+d
Kj3Y9Qt5PyTj6IYsaIIT42jJaiNGAxy7X8YkdygbWgidts4KLKsjyhd1VGzsuax2/R56TInz1JzS
OzvJbTi3K6cbUHrLPWYT1HR4vEWCzfpt5KDrkDjCVCRSbDGccQu/enPWLRzD9KJ4S+CtWdLMBvFX
P9u2fDqkpFEX2dIT+FC1Pjt4KidbM+tBVQ4/I3eNj+5V5Brvlxk6QEWOtYP/bqDayZ8SnVZUE3EA
wQOCIIYR8OPxVe+ujuDAk7dgrnvSwDwlk8F8cjvWYvls0OnB2PnEyPguqPE8dSXNJD26I/cWlXck
AkHu8s+HOL7YTfHEoMWyRA9UKlI7hIark2BX0QPqw9ob5EHTB9AJDL9kBIZmwv9FRiMNgoYSrEbD
mXSMnDR9VFTPRq5W29p/wNZ3Aq9lZp5f/TycLau0oXpc7gIrxtRqI7VjeX+Ga6gMBCdNHifEOiMf
vcr6BHZs+qnCtmpgH+deffAO9T3sQdsEaR+IqPsBk0znBEuwGcwya4JSd+HrVgJRAV+Bw64wPAwe
HxRu1WIBcAxFPcG+24e+M3X9mzIxMvb3VfH0GAbeDR4UiPT1zDNRDSSWk0pYKGuFTtC+EEflkv++
Pso9GWgRNvqTHRUZe/9RI01u1IYQl00x4tjv8d4VJp6E5qUj+f3jR68JbTsLyXWJZJYpCWHr2EeW
PlqzJSLxcZcsSJLRWHQlWoYsnFs/STbbD81DtvE3h94DT3zVapXOKB59zNwUpqDUY3MAzC+xUc4S
8M7jy9lW2uT9dUEaERrKIPCbqhZj5Xhc3IgFW7YxSPbe82wAHsX/NaZDVBx9fj8QiBTzjDDyyfy8
hclqJ3QYmiAUwkVUY9swuIn7QmRtzuF1ECCKwn2GeNf7FfC1IeCnsgBf8L1Ln2RXWdNWhu1+AmKK
V59r8jN7EtYcAIGvUWaAdGpDlpw0ahDR9zzIxEXMsCVMlv4sUhv4suUR6++1nSSz2ttGE0R5v2uw
eM6yCqJAFeYPfCafA+k4xz67rMZit/BMklUIST+iuOuuu8ad7OZiyVc6SryfOoSciebJXU5P6dSD
ZIcQj+1E+Mf7Mv1VFKpbJJWHWLfLThSgEb9C0Va0rej/G1UzXgUi5oVFoA4Vq7ojlIJZKmiZ0RLB
Mo+jGISblEKKsEOZsYXpecGrT12kGcOTDTCBE23XIczKYjfPeAnXhzlca40NIcQ+j/vC/YmYw2Yh
jxRZQMwstgkouEnVVo19+ugzwtof+Uj0f9+5YXJuJL8zJjUIkKFsldwF15wSzuZ60NwuNhBXC1gD
ES8puXdVtOSGX0qzsqH4VK046GL4trFyt8P5ATXZba8vCBSzqALEVij2P24BqG2gs0LFf5EdSz/H
ljityggh86zuzNWvBG9zKHOJBYVKStexBydOyxw5s6jS5BX5STEQMtXeJVJu4cCSEb/GSzDZw9Wr
HGfHS0uhoEOIsVvxep3EFuIZfYcxN1Rm9RFUtwccBBtXxY3Gf4AuEr7lnMx2gNo8ElCXf2anekGs
mzD06Ro9XlUeZCgxhWAdX8CY+YR730XVbT9E/WshZEQwVE+DbiZZyakwhD9MqBTmAR+eFKGs6rKV
S5/ccmSk3wYee5vhMCOYkWVJQj2kuSsdcYJ1Vyoy3YOhtlENRDi0BzVt4SO6TAa7BWtyYCEtcNvU
K083x/MIdMazjxOq7++UaRDatig/YCoH3Q6L1Ylu27vdQg0lWTD/0ef3dPTMf6t8nbDGKDF6v5E5
X/WGXkMeAjfb2tLpYF7bOCyRxNVNXkY6ChGKGGAzrt5DTDxNL1NdjHlOC6r+Dc/AuXY2YCcp0KtH
L2lw1OhthaOsrzpc2pGj2AMLmDiOrS4MKiaoqQQaeNGnl7Fdxqf299h3FRomidbqWrHwuMoOw3N4
Co8PVKG4QktvqmqdpPHyKBgf3sL6zvvyB1OAp33OpWambpZZlItLv5FbGER9Hc0U7dg6L4zmu6T6
GrqDdoq8YergTH17YNouQ6UdqFcI9hcWqEUSLeFOQNT81fxs9sV8sf+5jlsdaoa66PfuCuZAhQ1E
T7g6jpUmPy22k3/UL/A+Jlqh01DzP3TCo6mhxVlx4J//d0V1WtFF9iy0t1Y4Jh5vVygjyhmvQdl+
LiaDlQiVFexxl7JIiqStefbV6JhVu17bUS3qKZ6spw4/iZcRrZXIsW3tJT3PHtOKV7yx58K0/YZf
rT1Vext/Dm2cEc0ovHmON+DnTo54PfG0W4l6TbBKDSCAC6TQfRvVIer4esz70seTPXyY1Nz2Whr7
zssJxWa7PfrWWrCQ5Ugmax9UUBNUYS6e1/grd1AjkMAFdTsN+94IuWxVVcDBe4VxNtIqxUUwYu4/
e/qVy8kFfZ+a/FxbiCCmOn82hR9xV7v/q/nzbAiQ6/JGBStdKG+mPR4OvS3S19jNbbq0PCBvAh4u
J8XrD7ZVfvUO4VGYbiFWw4xhskG/2qAal6UsXkVfWDRmX2XD47q/K76L4VSingcUQwHW3xPrQhhB
hMPoEMIV4IMx3NsVmhFPXJDXkmcFco/8XLrRHqlvodDxOBZhdWyUpgIXjQCp/0O7S/0f/eF72HZY
KNNS6BQXzZ3IzzHw2SUy3pBGSnh0ayLZNCw6jxtW9g+jAYQzpSuD0B4ayUvsst8r6NaABNc/K5zH
i8B5umCGKhWYze5/F9UgDmnpAS2deUDhMzEf5zNUwXsxis5HTwTWDYA6DmtUqG2ujHkQb1yscCg0
YoxQjnQCvkvNJWv0xPj3JmLud6kE4LUvXXCj4IpZpS9V5Yhn5ARfY8cudkWrb4rUWDdysn0klzWL
koukq7UtniX+BoFRzksHOs3fzJj2nVanAuNDzezAddJEzi34INqBKyFqUjDm4Gqu/S/NlfBGZhuH
QDV8rgr0B0uXlJrPNW/TGayMuUoAzlklUCLlv4HxP3WoyDURkhKePxF/S3tZY3I6bVhyrljirIgJ
mWaLRfHEhuYUq528kkKrpx4VZMWlzCaBQYgwOZTaj+VktasqDccxSbpXRxxbGEm3vaceD7lWOeE2
fNrHDOGCv5XOOX31aQqS0CbaKQ+rminzFnEMAXhvC5VmVIv6EHyYo3JAZJGCk1y6FUSEK8tienYg
GyvRf6bdzuBwBTaIwVs9KNpztU7xHqa/95LXTxByKhuXbEeE8svElZPS6EsUTx8mRXHLO028HR0F
m+6TJLGNBF0TYuDXj/ycdE27y7bZ1Vvg75GKvwbuCUWhSppuUzZcJgsrUXcAhhDQGE2bw0oNsiaZ
i2HV8m/Jnb3dn7T5iNaof/mXKSBQieTJU1EWHSFbFNLE1NC1gcXogzv0hvkETVjEsqJ21cU1sURh
GPQowxYkq9H8x8hDCtzzRzJIFP3CWwHY9r8gN6fxMFfnMomQdOCg5ThdPMIT/3Omqh5ZLo/jz8yr
wS1bN9+H/lXtLkmCYxSmKcopwUTUIeQ4KTCPqwuNmFFWbYpMtO2uo7s+SFzRuZvXlLUExpIWJV4f
A//kmv01pwpNMxHaxhsu04ZXTxRVKMtTCzMrkJsEZkKfrTVF3pmilfL2d1W41Xxar69L02P0AmVO
zgAWdSPVdWdeIRzQGZOPEKRui8iSKXwdiY692ZeOBboWJbAtMfFus9l8H8+d79gaxgjEwCFotKqq
YmfyNX7ywD70d8N4LPwkj10+lXCI7lQPdoz0UvdG5O6ufCVCsuyw3ZcfQsYEVbFPHGcQlBYBXo/V
9HVI5mm9tx0+s7CGnILzlRe5yyyRFJSuNj6XvvbPC6m/TPzcRZS6BVm4xwMI3h/4xBnhXPFoQF5m
5mmtcOqmtuaNkRrxKUyStvwGGiVbQUt0PqjY5C4Z7Ufj0bo+ZaxP3ZDvpaT8ZzBQpdB/3Lak+HEt
LzSXDKzRuPFb1o5iM+uPWGDmh8XqpIof5II41PLFvtNqi3Cl6s5QHjy3yDix+qIj9G8r+mZq7hKO
0RP7OlbvyuP0wH8P4eGa8xpqAd0zTc4rDIMdYU1p/ICWml+PzmdAQii2wJFWmTzAlClV1BMt3bA0
mmejpF1ErUDFWYicpra7w3O101lpwUfdmNRadg4/ds4R6vcXByDSnUm09NTQ+DCD4gGZSGVpoOcF
uPuOodb/IZy9CBaiwilEN6I1DYVslNNRDheVgjiTDY86Ako79saptu+1+P8z70Q0w0rD38Z+m8ZM
EjmWOQ1Hi8JSIvDINrAB2Tgi8gyfyrMZpERB1u8qgB/+1yMBnxIPf8KJDNrFyMkjPge1GtDsWYiJ
jSjEXJHfrwThqr0Y1Qsg2p4OXy+b3WTSEf2NCBBD/dGm3oGrJJnWSHuvb+Z3PUSXlGDQ8TS3872K
radiKRRKXJMFbc/bZ8959kszs3swRL+yAS/xt6/oS+2rwThGu8HGQFS6P3BG9YAmWIlwBvRa68fW
nMeiX+fYizuttyJhkkwEvGUbV1b3DTJB3aSU/3aybgI0f3uVIcdvOu+wD1+9u1kk9nCxaZXlkh5l
q+McJHO+KF+w2lOcR4vDMco06mXzi/6Nr8iZ+IZXdFDeNtm4ol9cfRiCnSP//yu0QX8mE1Umc02C
pBasxBs3E7AQF4PCFGsSqYTWaAp1Vr4kLsqhhkThB0/Nln8w59RrKsyRBZg1SzV7mgBuIQvXoKqg
1JVXaWLMySNjlLqte+dL3CjJGw+Gvg+s0oT7hZc+AkviR3lcTK2HUUVwErVSjK9PTDnIRa9BhoZp
2QdmdOKZiTbp9xSJ3CzlF80XDDKOuv8dFznxmc9eIx93AX19y6QHUHIsGOOzCC7X9S/KDNCB+QlE
T+Wu1Cywk3FFKTXacbBj8gPVsLBmLP5pPnVOGDeyLfo4+IX9RZplkp7jDs2iTWl+bOsBFf8UE3BF
TqAtQVNdKn/drVvPdOBInYyximU0K0Pz57NnDbFDmaG5ODrOuetgmjofi5uwxfnyfu3AEtcdRjDA
lGAV5PQ/SNLC77twVBGQK/UtGqVbfmK8EyjMlZyCupWTWbn+Gz1n+yAabdv8L4yLGVn61pezM6tL
2YEJRvZX3h5n6UngUdOBVCy7tIOI/9U8qLsMGdLGnLiWK6dPiTvU2K3I0g8aoSrezZDJBEJj9Amb
f7gluKnua5tCUlRxdxtxSs+N7G74eFMMwKPjA61aqTZZ2oe9pX4vwOEMIPZa6te3sZ1pwDcZgeh1
0oyUCp9o3TboHylMfvW+KiVX4hypbKJsauH8sEU5eo6vaE7xIwKnnOG4oO/cjGqz2jtVArNQsnJu
9DGExTaGKHufOltYe3uavAZoQ3VGvIZ/pUKs8JrNld0iI9fII8wLI75N7lRFKexTbEBWWxqemhAL
iEymZQoFvv3XB47kpBYHLrqKLyXItJcNqQFKsVjTkQkoPtNwXIcGvwAad9ejDbOUR9kshdGEHkyb
Vm/J+QLe+4A8PHC0YIy4Rc0zUrWMrC7Sib9eVyoK+FKYiUC0zXS7wwNe4/jYc2Tk4BJ4/3sdaVAv
98kcQHY1I0KqXXyaMvP/jSMU9ZT5KVOFmPdR8Va4ZojCeuC/SH3WHEnNL3rCRqxT0OkZDPQbmwPF
xIv9OWNrA/7VVlNT9UXiT6wWk0I3fSGBlMz66il/VUMpQAKL9L9qafnBjk8hmyvWipoOEWkOAvRu
Z3wQmLkP+oUkvZd6qLrtB4kiymLygNZ/qhqbk9GsXzVzavZ9NyQaBlxNB+drmETMJUlCCf+SCOD/
wdxT/0Cwf4LsUUq5PHearyzD705Z9QmPgRlcR6RMa2GBKTN2nN8NNtFehRUCjuUDY3fALTk+152a
HpveF6VWdXfytucc0iuItuXYpVWqp36ctWxicOHf04XzK+3IF3UREbFqrz/Iq+RMOT9n4OBnOmhW
UNHav/tVPyge94DNyrtAUHfRjx2H75XpJUKGcXcphlBTD0YG0YD0nJrbgeYKo5yTH2brJHU44eOb
rOh6nCE1A56H8Zx8IJic3lQ06sGJSwAoSt4rVWu7LmBIQ5+WYcAFeHJCRhu4Hfj0UpYEr6N/iVYs
3hcUt1RM0u+XPEtaRpTcBTRhBbBXjvsO8vpMO05Y21NgH+g5SYCVvW3F+EgTeDUngDn8NXMS7RZj
eLnwU+5ShHmSJLDSWfJnt8wSiSPOTobmI4iWx38UUTWO3/0nPT9zImQtaizC5fF1ZCuaT3nLsl3l
JnItcQkhyqNtBQSmfS74961754DBzdrU+7X1EQJTdeA4gqE5P1W1Cw1yJzOyvIhJxQk/YykrKVK9
ns9/y5oNIzjnqKWlJsITCFgBLLwbgWVga0itrLTR+1QXHNAD1hWHrLu/yCEzPyr162rokMjLLDEU
CLmjGcUQrCC49fK27518XFuHo9kujtIvTs2xVdGMKx1YqRA8EBWfuGYHWlXfqYcSvmzhIEznycOy
jcoQZeFOuqEtYMNqwYPBuwk4auERY/2+HKEuOkP+IyZy/CoObpVSaXfNpoVlYEfRdtosTm5okQqM
FR7TAkElQ/MOlbT+hqVtF26juAlGIV84K6NS/0X8VmPVSMKWi/dRazlzN66f9Y6iq0c5FLHzWDZp
pfmy3NeHcjU/T89CpfcTK5559rD3VLQRLbd1/pmMhemrjgWsGDo3zV5woAukI1QSgGaFMzfFV1+W
l3RBKnFKwzXbtyUA+Rsab/GVs9x4/w1O5G/ZzFUM3zyfnQI+UyoRkhfpKn5WF06KhBrFg+zndCDA
1tFr7KArD4lqp85/0V7EnDI9D7mXkbIp0+5f7aZMkb51wHxAQrVZii4/SLgbrYEJ3pfphBEyWO5v
BincHyK8ascvrPfZU116V+wbGE7mZxuFECpOQCaQtX4l9y49Tg80oRvDgk/LzgS3/uPnmsXnLQpf
tsoyG/oLHe6m1UM6wZ6hH6j+rkSjanQjqsxSGxQxPG+ThR3gcLOUjTYqW09nrPt/4mFkLpDKySN7
jRjpI6rvYg848o43+rOGJVEI4/Wa8PetXImhP+gV9fcdvS3bO8g7z4EPUplrAZGzuuueVChiuXxS
XBMHKyD69bkOju0g+ZNQbQkDLW4cgmz6g5lsCFkyLgWC0YRcEJpomeRhTC0GH5J8YxanT81KGOnR
w9inTz3QgOmkGFJG+m0DmaenjzeZkoNy8mwwgz1wHVLs/uMZGvqIwR3OKsX+gRRE+xW5UyjRTA0/
QXktBLSIpQZ9f5xEuaVBUmdeCVIXsrA4Au7z+8nvMePXZyq0TjaeyjBoXVNj2QC3sTDmeaaiXBmy
A6b5ORjsY2c/sdk5uzOa7nMOHMCjkUkO7nJ5LYY9cULr05EKnImOg3WI3FZsQMjilHpzdCyBAqa+
4weW6bCEgct8LdcdWBA02LnhixXtqdUmR6Ku8hPVDg/NEXl2MJS+sMtAlUT0l4vznfW9EsMYHxhV
UB6QeeynKHp4SfqwAZYydAF0mz4/Z6lY9mdCcJaKWLxntJHbjEMlcDVqNl43MSNRAb60pOMuU+Ei
jonKh+O3aslNnJd4lTCj7BTaRGnQuFfULYIs2sy3zdtVQ0vgDeGBVFAuhHsTtyWfZQkTP/4xuzQ8
emMmnDeOwqcNm2ag4prv2oCVTs/wwgSXmiqpI6iiM7sAw1n5du43aui07iKQeAAgYipdsvaxdVs8
8PtbcX4Aub4ClTbuKU4LAnSxGI5L63Re1h+ksTpEc+Zt0ao++qsUZsIsAC7e91767sFyTDGAYdlq
0u7vf7uRVZccinre6wMuhP3vloHhhIm2XIy0yEELU/BqT8a3fltV5NnU2OcS+oz5wvA6YNJKm3+d
WVgTAtefQXxIDOCm1NW7c1IYSFpeYQb46j0sypLDwbPLNNVmBhfQWuQdoxsZparDd9NBJZEalpHW
Nh5xgEQDEscqf9LhFZ1HngCPq/IuBT4IFdIe939yS24cKX/MdstCttWmaeeetYWCZEYyoVH63bxk
S1MV+FptdzBmoSZ0ANawJLQthiFChDPwoarj8G7j4vBHKiaCny3FHYhM/Lt+95Km5UJf1xIVV+7G
CuTOLz+iByfzruHmdqhFMUkxo4soKn1reEElHwulvPyIL0qytdvOl9vxxMZvUNGjdpmS6bju2ouB
dR2Dmr7ELsyJm3HySfJWwwKL358qtm5LglloWYjth0H0DRW6tClAmh3m9AuJWua1Drm80WfgE7Ru
l9Sgv45hCKb4Rx/vjuwugWwMk/qwfI75mH5LjuOvFfaEdQEKubfDWmtd+OZxHJ4derIhulDbbZC6
MzhKyOrqg2Agj23YJSmA18hxX8K2c762puOcJ4UcJkZteghhP/vkoI7Em82jFPunXlX/784GwnH/
A7Mr7fAyQNMju1XJd3sf+Up+G7JPakVPTzTkcHjspDmiHjpUnUYEp1Ucc9hIk8CcJ5rFsdOWOVHm
ZpYJ4HJU0zIZitw81IgKzwwWcVEGqjec8Ct1/Ci/rjA1UjTOyPaMqs1K4bhzZH+EFvNAvXONhXTQ
ZpZWBd3dLL4lNk/GWhyCF7bOTeTt2RviOSqEo73pJaCAqrx52sUjXJ1N+6TGR2qf3C4m72/5o1pZ
7WKoKE0FjRtnBjYqkP2uf1K6ukOAAIuXYySGRxGfcfSXISXKIrcJ/LomVJzIiQG4OEFbBrbGhrPo
FTNNfaK9op4f2WkWM6HYKPN5ixWFb2xqzymai9fGnUdSz9cb8QHx7O7wtid0LdF3pcJp+XibRusV
CF8pB+PCxFlE1OmiFlTpGPTim8H2wvf03OIJVv2Myxsg0EXtMFE5085D3lVPEanDvjdxWrBhQXm+
ZzSZT3R4ouB9V66WOzhiMGPMX/Nbxocz1CYMp6QE9SxxqDAgNW5NHOheg5xLbIb3pk3IiUzVo/Dl
8BP11aGb0WQUH0vjAS6+Phma9bQ0HaxFJLRpeKxwGUYAUuUsVR0pkoZd5/2lNVqSq4xYhLLyYXe6
zQlyosi57ngx/LjYIRqMPlVOPQpQRbnvxulWig3rYYKWPJVvKcaus4g3HC2IBfop3Kq6QuupIAIN
IOYOPilnhNrDm+Wl8TTlhKsgc2W9aAmMfexsT5kLPXODuVg7DYRxj04op/CZ+A2jXFabkNHam+ES
mtohkPmMF/mDLXt+aqowKzhVsXQ+BOtI2RnBXWmCo2rW8yHCdOPxubKwBj3+Em3786wpZxp5n0+x
BbydzfJJagDhr89I9rtyqgYBoa4QIP7R4GN2/IcnKy0YvvEj2Vn6wjlQ35eG+WuBy1AdXk/xXUdS
8uG3QUJGOnfCmYCszbKIvIAVThaEXIII48ZwcZvzXIFoQ24yJxAirfLpORxRiJxmocz3lGGbzSZK
6+QYLqT26gYWPZ9MLm907n1Ud71RW+yRsCMsqTmJrbAgPd7bTGa3m5M9iGmAMxwAIhibQ3FnD4Sz
gbrWbCi3b6AVJknrluBZm2o+CniZypjuLwUXQ2wubI+PdKWGh0mRN8TiMNmtskC6U9yuhjzAfv0c
wm+3QhpUbpC+H1thRPefXv/NXdr/SLN8r1Nl0JcBwSbnL2gjbSI7IDGSRAdeZMspDCL0bWe44Zyx
qeQ0AF+jd3XcAoPQr57+hT542dWZKmDUXJdLrufgNPf9Rb2ALrlWFsEdXhdub2+9///jUwOp1XWr
NijFhJKDZqeXo03rsgtS41sZ2OMtSYjl7K8jzYEm2F76nk1h9sRod38o81yxpy7XoGivtG15npPm
m/HVrI1Eq/J+fJ1MP6AYTVzGa37RlNATPzNpPzO4jqdYUouDB+yxpGDOhVKlYU9OXtFVZKeHoSYO
SUF500SBgm4ooxra30nWcbzP11rAT9EpBme92g4XfwA7bsATzq6smT6K+3mDZ3pCUZgqlD/vv12t
JLDLMvJTT2RMAfwIyuXsOB4y2pv8rWn1CeI1MRiQDtS+sylC+GL9P4PtRmjdnE6Hsj9ODG1xpDkN
kHms8bUw4qrrT/+rJ5JsQfD/jmbvjAiET2qWgLoSwTeaX8gavfa1GRuo0hKu3WPAlSrnIWBIEnZn
O57pSOWN/xXBaqi2ie6T/BxUIGEjOCQCJimR/biXxIYZFYFMF2owN4xNZOFXCKryUQbDvNVAKb4W
EuJftcoHA/It3v43Jwlwou7yyI+jBeocT3b5dOW2Uy/RqMVM969cI8DmS0cIpQ4idx2ERFwP/5Ad
gOJ2TN94PrO+Wkl7XGjDB0sCpYIp4DhenIsIaBNrJxKaIOOkKinQKNemr7Y0PSf1NMh90jUlrSW6
ul5UHDQa0lzz9ONGk3t2HI+Ei72wCONQfPYXgVWFkZnR4zoI7Mjtz+bt2Pz3hupHydm4ekUJJrV3
VPgxl4XYYDd5N2dV5AxeJNgSN/n9rl8qj1CNceMKGscLI8WmgJgU0M/KbL6CHqay0byeHwS2tNED
3szc/GnCcPxlZJeqIQ5pR/lQthwDj009iFGo5laWgGIpvOMJZPiIFPCT3eMjLg1l4KX+hND27x/j
q1iL+mPG+f3uxCxLjABh0NK4o63RkOQxRkcSjwnIcw5OYWF/WFGHGR/tE7n9dmxv3u+lkIPa59r5
ZaAHv6ybqRLm/+xepIvv8HPSEvYDtLL1pVuyNLrGTx2XxCTCJBqmgMG7PD7qBhHh/YXEoS6TvBnP
OFJIJvlGJ0xaX09iE39LyrNrmWwZtmGVCwdVLYEZQulXC+M71qchMwd/Hv9Kvcuu1XB28ZL4H/Fc
o9QeKwrjDox/eFyvylYxP96cd9aVcVa1gEMAUUl8qC2HHTE+27BQgajbtuORJ0sI9tcyJMowU3qE
Ou+IKnoxY5Qpee1Mkc6mGm4niu9vtYTPxhO52q6sT4xt5sI1o25D2zvAzkdqROFhwBSF9hdmG1kP
6qGD7z8PILEjyK1vwKiufbWcSRdcO50Qn1e3Lhv4P8ebH3lp5qORTHyyD+2wqsgj35RNscUA1S5r
vsIUe2L5VOE11UG4ZQX1QC6DJrWhxLTavRUqv6mNoYL5PgLPaGsMIx6MK1HVeahHbMkR0tbrGGCD
Q1eD6R/S5H9kWBWs9JYl7u8iWAwy11NqJLvbmB6S5EXBgFZnv4RQ2YRRsv4AYvs2fBEEp/Jallua
chpfuRtIlcVq03SW3D6c8MQQtF1VWPJN234h6MiRqM/sdatQqdVmkLZ0uWg5IjetnJ/YD0qYMvoG
QZAEaS5Js7TPbbcaYkWypbFQef7tvQMTHG2NnwZcuM+s+muMihVQKa1WQbjCu1/bMOQ8Dlu8oPkl
SZmELs2gLUnp9sGu0XP+YNOjbDSDTLBJ1SLSCeitTgIvKb5RjLFx1dn0iAIjpxDle7Va+PUjBxp2
i43ty9rG6QYmUAmeIGs/nlXa941Cxs6Oa6MgKpxWHFds9T1Jc4aAR6JD9q/+4P5bQ4QfDi3y5lY3
RIyU8KTBwy7VdHQnz8EnNPwMb8yZQk9kX0pQB2Us2ugbyM6IYKzQoLdzqCoDGWcyxEvTHeBKj74k
tZXiQKWuXou31YYRxVxC6DDBt10pbY6K5NpwbGX0SiP4rmKR6kurqlmfaXty8evC8+ULcF/jwz/W
gTJB8DV6sQS/0sUmtkMEHAU9284WciKJICkSliVRuDsDu//og9IvbtD1Rc5r7Q4gBJBIbEi4fIPD
7FNd62zR6/FuIjwm2w9Ne25J2JxAOjPZ17Do7G7+f4VC/dKN8TjUVHCjKbFuSB+gwlsOsqSjirm3
/AcD/vOV7/eq5hbxhY+hR6w=
`protect end_protected
