`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
X8wsoMgjeLYkTIc4iS8F+6yUXEMoqLxlZHiEgUIpYy5STdFjgLKaNhTcLBWpDPukG8ZBGLC9WLIW
khwFiuUc8gWqmUZpa2YQwaX3DOid8tqB6/SyYNInfQHWk8ghj7oI5V1SUxbOCdNSeXIN7Va8Ay/k
qLQWn9ZhcDRaRIxM7K8piVxcSEj56UvQLk01ayQUAjvZEM3Ln7dWtKTgrLrLkRo6NYe+93Z0AXpn
xzFmpYiCujRs3xdo52c+rgcimYMjHOB8j9tLUjNsd/rhMhUlZEceshEZ5e9ZirmgkihZ982WN5wb
HXF8Bx34pmQw87w2ti3q+rBSoUjiXg6rjkhgHQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="s1teZGT5UMH2m+YZUi3BH1TO3k+IyJZvM52EBAFOXCM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7648)
`protect data_block
Tuwntw+Sq5M9QjXh3ZAMThVj6Ke2/6Y57+XedeOh+td2jNfAFZMLv2E+Cpi4J/dXIQ/QldsOIpqh
DutcV6UfSsS4SQIfR/+6C4hUjYS6ktKgt+gzeqNnvqus7nzzmfU5qsTyk188kNSMdW5QwZ4+hWNL
4/njEm1vv1E6nf+ydIqp09jVzP3oh9tA9ER40D4VSR48hu+3veWL5nVuPjYYDb5/jq2W+CqpkLlR
Fj6mKmU2JCog4gPxm+RJd4KFX/RZWaOmyOQMwlo1HRrbApspmVKFeHVY/J6fv5OPRoGh0/CZvtTD
/C2+QZHw0CDMvGqeRoMkSLZ4C3UNDd4go8MHYxp2X+fqApbeLIfHWHn82udzShP2E7nR9TEn9cdd
pIgNzhf2csPVymaKKaZQtxJZ6n4reZJw4a++2iPiyu3z+aTAY0PD4vGQCp+Ydy4GsdIQaixXibYQ
ThVv0/SMz+QX9CBWKfftKAtBPVxByruenQPOS3z5T+HAYuHW23LrNETQIT7VFU76SUnxwd7KoIJ3
F7Fz0DTM334GykvDW4hDxjuZ4JPaisdDoVuBHmH4Q5ofUJQzCD99rKaCFokMUflUughbJb3eXau4
cRjYOQnnYNk1kRIUxlv8+muYwV3S1/6CRZxZaJ6aGxISD+JxctzFtEi3JimkZJE76cPqDlqGsRPi
oTBUX2vX63X0BqowjUY3prWSnk0BWHXHINnQbymJ4u/HShZqlLMgE/wd47GTxMg8ll0XL30kQWyj
SfnOOMU72Teym3g+cOKVPLfsN5ynoc4JGTKjVSYWXIc80kqv+hpGgaCZ2v+QzjweP3ETkH43cI5F
beHVyMEBFuQBHmic0a+pOUx5Us3WCZ0X2oLMV91McTLiQWdQ0XjS0LW8DSvQWoXI8IGSBNcQye3V
pf1rQc9pylX2C7LrCtOtYZeHID9HcW6Xfn/hDWzSGCMbwoCbeBKx95x4XlRd0nRq7cL9ITMm4QHm
8CXJWlf8XkgIvvTCHJJv8O1PlpeSKUQK7fNfP63JkwIFUk6h6IPDc7k4O5sUf4OOLM4ZaEGx/T2o
T/WiEe2CTv+GEf8KqkZl+E3iuNim2EkwI5K/qpk1qmK17PH2fbxXtrHEMg30RjR9YDgoycc6qe+x
kgG547taswjN0OFpcUnhozDWx7Y1dEIJRmBUxjfV/mp49pDxX32ACFJ51XMO4EvsvMrfXCOT2JF8
ncm707M/NDLkW32nZt0ajj0+bDQ74iUhxsX8iGWXZsFGHupb0IEOu2G0CKG9mfzadcWEDRUI9FbI
ihC3ldzqXYmvkZt1XX6uwShVW/trKjFKKuUpJwbIJYJsD6oOQMKsbu/+3pNenKgD2l+XXQ75KbQN
SKrbudZ2UY+ZCq5A+4Z+mHuqiU0O49yBHpFhz5BI63YNiGQTzGErVuYyyGKpZdb7TOXTdD1KbNKc
OlwILlWDnMlZ/niCV3SIcrHyJ9RZhQrGW8nhWYHZo6CWeq1iyAL+uHEyKRagy7Em5ku0L8e6iQLU
H3kCk4cXy32FY6bOwp/ZHcmZFZUsnqagZM6uGssA7lyGu4zLb8KUalhDsRJm7jZEyVy9bngStdgr
c9VB3SbHAhlJFSh+k+aLWaL1O7rMJZU0810OCmFD1MuKOGn4bVpQ99QpjEZQfCbVC3GRKKj4WjNO
IXCCDPzzTrGqa7eHPiHdOB9ghNGwoaMgBflmH3dG6azEfJwKV6g3PyffUwYAAeve15pO8RrFwWvi
g+/yapN4jsg80WOT89LwEh+EIlbhy3zQinF499TVEmqMhbkyWAtkh3hTGMSgkbfbvBd8Book75rN
zZTcQL8kk0d3LLf94R5icNu+gZjnmwQ4O6rmwoh6ihpwaRxWBA5Tf989Wi+X7wmjfcCiI8AILJBx
0GrWFqZguEiYUcUB2/cFCOQ8egeMZKgiZhP/J+GhG0o+wF3Op5p1k3zQH4w+D3ywQbY83CMDwM4B
tXvy04N0UtjhE+2e4w5F5wdHLxLwaraCJ5Tk+MMycRpuiOFlVxH8ZOOrFofOet1NtKk9MDLSFyz9
TqRZMgya7okuTbVIHpz7BqNKu16zbtVS+gHvWQmaTaqMFXKcalx50VdvczJpKjAOqUahjf7v2F3j
nc/mR/bnBeNalFgXE7LPYg6ekcHG9R/vGO9kAiWeMaB4JJrJ5TwYYCHmfJafJxHWetKNV97UoZpK
e//yt5gll0xScE88MBb37Vuj+tWamBtvnJfnz5nPGara7NhgfnnwWafMy/NVmvJsHBLalXnAPYS2
z2ILmES4ZmOT82462uHava9yRg1zzfmfmpkWH2PVcq0VekO8bvoHMWu8b8N2P3hXO6KzprGMlY2j
0+UuY5jcadK6xTG7TV724lYMcBXoULEJ8nhard8Nj9yesO7Li4XgPAC8Cx6lkUbJHFTwqSmqpecz
BLEAL60C8lpOuDo7bQHqC7/hbEbhsDUT9WnNbw70BawHN0sDL7oTDK9xAW4DmuwCr/g5YNtQR4gB
9b8TVa0nYiswma7kCTBVPhRV16MsXJe6mcf3xpgnBaw2mEV+77jT6LDMNnVvr2JqtZhxWwDopLnv
7bXyGj7ognJlJhudSZNKHIzyhHA92WHTAf/5JyPX+mTPkXchw87k4pQZaQFd4KGY4sbnEFVA+z+e
A17/DN6SgRj+6dCWrfOIutkTbYiHpdRiDvihC+S8RTVqQyIubwSPc5S9UWKMn4HIfB7/vQh+aH95
GZv/SUQmRDs7PruqFxb5ntP7i2LWv48sYXT6gQC8TZMYCGao+gSk1E2kyaiZW/FdQJm2WeluYB0Q
hnFI390XOjBeULwLHgIua7ZiSRGHtjuMIYSeZkxx87M97OE3YRhRD6Bfq3DH5NmFb5GOLT1wlgzQ
rm7n21NhfF0OrCOuh6sCwy2AoreICycyma3Gxr4EFMgsik5yDRs8LEDELzrOAKnfgM96fgZS9a/B
czKV4IbFOHvkSH19IgVenojRJLsUhh92EwcYRdOnPh64w9xzRjaiKvPqAe+Wl4QwpUD7v0iIkqhG
G8G5jNlAvTIAlqcf3NUU/Nivqqvcae4nFCHlruoUhtRngeliwPJLhfRO+z/kSnglB7hMwlrrNVlY
P1f2D0WBVwUiez+q4+TXEkaDpWJ+dD6EXYfYpOX9o6RzlqQuCP/CqRdQKR1+2sSzBVWTq2aLQNog
fj/lkWkG6LpHKyDwThgZxgOPIYgfn1qRWnxfdeelMlaNZu8AiQoR1xcTYHF57wRKHkaCQctBjI21
2PxBczXLbY4DExGYLWaP1EiwLtUUSS2QdV/HZ1GC7om8czpNQN1+ghLQsn65FTu81x6zcEI5qVbg
6umPFlCqhpDLVduuxU1akf8w3AcMaKsrvvDjRAcccF6uW2moHZXJshLkdYt6T7OKGu4yxWipl5fz
HuQlFb3LpuZq9jICKQdZ+m9nC6tltzUeNiuuJenl/DUuJvexXVJJf8S70bH+OjpIdo+bMbI/8nf5
ilFnCWdj4azf66RQrwMzEoWOnySpJh0t2HMhBUsz4MUuUYM9mn1LkZ9TEnqgkOyIwuleYT7paGTU
xfPTh6di81HViegDcqVcxOewI9g04LDHyClkZzci1DJA0lex7UjgCo9bajOaCD2KIKKgboYVba7S
3obPGTKswuu00iFw5UTV3t0eXiv8TCFuVq+n8Qta/0n+NZySuKyumuD4DP0xXC0ultiEwU30eiss
4ZlBrplkfnBuQMTjdo5dVxa/UTr+wu5EEcavNvZ/lSSsRCB7MD6EBOM0lltyCfpwdHa8HBThm/As
qWPSLKiQFEFPBbZg/+G+nr3VpDmas9BeSJtrtAEHgAXv+h22FWtHopOzxx5aH2q909MHL2jUxdp8
MU1/Wt1wnYOletIWkNF6uuG2hdtjbVRThX0mih3pgU+HRGBbAKJRZyX2quSOtcRzilGRQGnpG2xL
2689W72UsYEKvhcINd3lCNFk3QV1h9+ELeTR31SYlmOkP7pkwTnaQet7GCuu1D/KQ30VMAaoXwyz
93hCtMUmVLmXJ2d7mfDgmY9vmxBLsYEr7mYmeO0oyJj7T5bnhcF1BKkHZgRZI2xeJXQMkUmijdS6
9rO4yIgvEbupCVlxr+znxCA6GA9oP++WZw6wLHihUyzvB0qoWrTaOpvKZMaYvBiJAYT2GyjSZFp9
CHqYn8asJySeFoeRM5DvaCpaBZcYxbDnCD5XmfXJl0s087J5Uob3XQ6Yelj/xcx04pF0xzFIcEg/
9ge8NEPG/omhUoHA2RkW61sUCkpQz7+i7XOURUEbMfZOLV9JMsuM0jWt3zlA0GKVOyYKOQUnxmmV
oiwv/5MZy7C01npn60ptQGqXO9iOwp7y8LUd79tCjivrFXHS6xfitR99xgTjeglVI8pcTs3JGlbz
VUDGyaFjbEC1+Cr6PDq5fjKr48F88SprcE1e1u3cXAshifJaP2V2Dy9OPmb+nJrutXYVva1cFvCZ
2xSvEf0Z+4WT80zvVL8CnXXhazQw4B1JbHPVRR3270qj/wembrOKA5/OJxCFWLcQ8PgYh+l0qdT2
Mxup7xgQHYFWboZkmw1LBzwarH1aI1JPuRx8tuko8zxi1XujXVlGPsx8+C9ev/JjCj+7pZaN/+pI
bLR4zdAzu7mm0NYP/7G/sshDj9Q1jB8kkSBDNnZ25UwvPOM6LVTpAE2iu5i56+FSC9JpDt0DiepW
NC99vvx0GzDUJIWcnMzQThmwVc2uQiUdkujFBnY+spynLAKDOqcTK+ruqwJYA5zEmsnyGzezt3rI
aYAV+lhj3XXYtv0J4VpLEgkL7A1mUUihg5UtglcjFBIJwlVpzbXujnjZOk3UQrXYJdwNI4hkyNt+
VGK3TmNf31rby3yEjk8K2lFEvH4VxIFAeMuoagi/QVBiYfmLJHzDYrTCsrgMw2/aaQz4WmBiTJ20
RzyxkjALhuH2MAflbwBfp9mtPvahVficjMyIa6L9QzOYGyijNIXS8Q9mYfHgsisW2VEfEALrpkJd
Dotzqypf3sFXzt8idCDFIeCvmqyJv+Ov1QpD5ebtOivxUU1jay+oTw6+yUJ8HZilgXul3QP0uANd
7KkUgGjKqb2xqQ3bjPk7SdQ95xICeJxzbUQdXi92jFmBAlJH/Fgajb8M336sLyCGMO22PSRnl3Cp
xzwil8B/Bnt0OMvF6nGwdSWsEpfq8iQCfdgjs9qctngW5lFSvX4LoOQih5RZDGdlfZ1KOZQCtENv
w+BEeW2RoyC4g7YSHotqkPkFj4Ko+CSFZMJpUyy7HSD+65I4JOWYR1VZ33hbwfjuppKR1KMl8RDG
x/PxrCEkcvqRk0c2OP47qGuviyGntAPIF0ebLCu4n2EuknfdrgiutDRNtJKrzPwWUfLD2VTNqAGc
zd73vaNcJag60wb6JJveJY8WEBhDCC/ABO/sysjrjOjhUifl3cSxQHalxfC7DoBSdDQuALqZNo+4
DHQ1ZF50X+wWBHomsYekyWWevt6O9FpU/qV0rg76vRAwwFTBQ/TN3hCo+C5/2rKR8Esoda2slRvf
8AMtCwvKmvPTTPKbCX473vTlcanmXDBR3zlh/rIr5LosqLmifFSIqicWxFCyVE3a+KZ0+Rm9RVJo
K55JZPqObZo90wNgbW3FS+x2LuI1r7gWrOEM5Pf+Bw8TmT61Yh5sBdX9BAH+wCXMdC9wu7DkDwqz
Rxpc48Of7O7NQ4jcZDzzUmB96my0SVDf5xzawcQ4z6LI8CT5fzVzDiTuOkCJ/hLINQpvbetkrGop
KNHy7sXQDo+n4OXsAqPFkU16Aviy8OkE4hVNiyefR6MTQoj+nBkRXacX1cYJN5hPhj5BZB+I4FRM
CPu3k5js1eU4/Wv85Kv6DJ1CHSCR7BmDsthdhq3XJ1zIxs2q52tBIbcTE3VJT0gwXWGrJbJbtgzC
9rLLsqheeBB7TiaTRjwYG8VRqKLqVLJOe5xsPmqs0fZMPdLqTGGvklIlB2fxdBiHyQE7cVd0fJmr
WKhLNlqCZQHUmSJsDb/6anK5gjTUT1mjzv4nD/TV9aEMyI3wVWbhIOdpxGwcJD/1VjF0mM25C2OT
9WByAVFRqRiQ2iGjD9cd5JnajC75ahJI2sz8EKhWS5gzQpEi7pPcrrgRFPSAHrZAQCrqsHW9ywBI
t7w+NvJqFf/1BdP98G9cOctgs0msN9dSxVapfWRI3Dg/T3vj5gnVYuf/xmtjRK4c47VbkMP8T1nm
XTmlOaUPeNfnQO+Vi9xHH49A5ivyL4eOjGAB203pzud+MTull0yGeLv/6B+PgciBTEx4OeVMFusf
ekrEp4mr+dRnxxd7pwR9JNZv07Nv0EyF5tmw6FTEa3E42uHsCB0gwU0D75P8V+qhAoeTlA1e0AS9
eu+I4t1lOhscU7M9iineHDEOzKRO4n3UCFIJNhXHyEWoozhvrz2roPxsyYKE9eNkMg7xMj1iDt8+
CzBkAShuXWDT1oGEf/4xDBxCF5K51AbDiem/8A58eiO0f1ltNQv2D0/+SQZPBiBst3dxFb2CmoFu
fr7X2WXlQ3sCSFbth5ZuEZ4xfKI75DHuJ2HS+ieImA8NuSq7VnQup1lIobRAw75CfZhlEYfD27MY
wE7tCraiyy+ANSzBH99oi4W4t8kaE+nzZps/OkmHmLu5zxZ9HATri8XRC9N9CDD/pzZpRdXe6ub/
/YvHIMbRSTOKaVCxsN0FgYi12pPHjPc1sy0tYHCKxRjNQLIkGcr0SJL533D84Y66oEA/9cw7K9Q/
renXLochCLLxFOBjzx097qvQ6BN2LXSEbw/E7IhP1TKoNjYy0ONY3RfnrPhxxcucyFCi6ZesDG3i
4YFo+RKsUBiqnucd1EFrFfoFl26FfMqeModUPZcsOoNJmOffOv9yieabBS8FgoRgRdfU+0kOji3Z
bMUtzRJHE2dNl43QUVTlwZ3SFA0QAAYI0bArIy6BAGdEbJBq0sMfrV+giq4PGcwsMonyyDp2K8zZ
eKJx02DjUHCW3knp3aQelRY6x30jjsIMY7bSn3jtJfzilH6jkg74Zxi2lA1fStso4Y0oTRLv9ydo
TdLdyLl0J1iOlTV3nSu/U/aOkKgBQ86IBkLoyynp0yWxl3spIO1rdfIMKE+ORwnU55AWuGS0jkQ4
hEYf40pWs69uLxZp83DSaoWWJA8yJBMdM4dVXvFLfQYOlLWE8LjFgM4RSmlFGsJ0cGM74WhGYRAk
fN4VSEbKgwUkalrV7NRhtBOJT4AZelroXKM7DiXGgD5SolW6qkl2BbRKRGvE4LRZDvp8uBPPtDa7
p6DbnWl+XHB3FcZOchSeS95VhjPX8Kh7vPAmSU4sk+sCxk84yRjaVC4TKr1wDeYalGafG0wrpsxQ
l9EDmtbLQWpKrecQ47pud13pBdcSegtwrWvba0Apz2kU41Uu1WwqpbciyYX4Pfjilpmb6MIAvTfe
8rtDD3HU9ieinbGISgu4vY83GfKQBPa4XaVC/Pq5h5qJdwVzE9zql1daxGfgKKYlCWo8+eKBTdGN
DvEYYStpEovpavr/gocLkqwMaDIbfZJrFGHpD6aMjDpPSfsnDRdIvzZNM4F+qrv2m/phrxy60YAK
eY6T2mn2nWYnHeZlhHNys7Rr264tJvnxKQpBjUda6pLJHH/Kkm7sp87FUvqk1qH8QxKnl6LHNQV9
iHzZShC+E/KWLJHpjG90lMjFYd54aiOFsqW1YOFVIR1VzFJMIKqAQa446qYUwLbGJG0/fBhDCfbV
9vxacKKwjoRdAGv8y61EADKOZmIkKKSPkCHjPZChgH+lSi992VE0Khcq5oLdOOK2fpjm3oxt7Ud5
A6ANBN/9Jr/RTGJCXtT2z6Q9UVRJGi9PCVSlg+1cLhkrZnKTJYDz/f0gGhccRzrg0jSiv2mzaIkY
oWeqYZCR3wEA3/5PocKrt+tjwgHkIZSuLydkds5dUXO9qL3ETc5k9lLJqcFyfCB+vrG2aG4lOgZf
mGZ61wz8PADvxLvkem8FrJYC+BnxMZwzDzi+jV3QEcV++ubH23cveoeAnwKjO78ZrsjvkC8+qqfL
V0OLWOHGdqmbfOeHHKZrRyBTEnDpHjsZme9hnK7xQ8/QKh9pV7es+PSCkLmFiVLhGmcxW6M0gDFk
syYVXtReHw9vdQoKleojE+icIPddoXxn5IOAroBCT3+77YOH0n6BJwzFYk9pTkLkbQJrVR8z73S4
KdlHre5HgW9ne9OqiDeR1YuQywYKLuhWaN0AfFWRCxW7oN0zEt3Wjh7KpHXvybQu7/0MEYaejeks
10fktHWHUEysi7Sj/hUdwqSKTq+VXKzfj6SLRvxxEq+SdKvNTqvB1U1Xnj/0uZ77nIlW7tNYAvdC
ayhN1Hv4JEoIW417yRlzTPi9aB8bPN4KPK10mNhcBH0g/EyO3GNcJhESlOm2pXie5fKKPUTJdeFi
qep1v8HUlth5XagzQPRL6KVK4mPq6XG5n5viAaX5Sg0CUhYg7kAJuQB9cYrUljQYEa44BhP9qiEi
tylPNntETvu2j0Pd/AYugzn6GwWwug5a3++NXKmNbmYYYmYcnNqustJEuB3iX9H7nIepJehbJunq
vceM5w8FFfZoPc0l+mGbMpImtMpq9AbTc7+lyulPEf/nXcnUjoy0qfWMb3s7CB5zZUAbTBSVwqmM
3Orij7ezaL0Ybv/yt9TA3LD6COypf/LwMnmV1eyrRkL1Xzu0D3LOEkrMIB9MHvmJsjlMMAgxdpBi
wZLnS5GnS2su2VEw/Wx4Uaz0CPlBdJcjFL3nSqPXIB+e2O8k4Ez/7jeAZ2ujvtvoXwWRxunyruLk
Mj4+krgV68IazjyQbtptvdbCuqTzzuYj18M4S8k3wyCMttUHlGNUjo+EvySooMvOAVigcx1wXQF5
jIZRwibBF5KyCielQ/V2nd17cR6pAS/ctHSRGwRfyXq3BWh0sU8pxVb8HbC3Yrmoew3t2JX0iPLU
lIg0w5s3ZWt04+E7YbtQ3yDNORFDvsqa46/aB8gqnIHh3aKZ8EzA0O9K8m8MFQ/rubBIhOli2zn/
U89PwLiN9MLkSlT9qP8Cya6yxxMDpIKJoLxfFPKZGlAMScRi94qx8/SKGpPEWzP8TH2wbW4wTbKn
IY6nfiw64TS1DnCkhbSgL6QUvN2OFvHlyTgNAQghJpFHwO3bV5R0cthkZyKQMHWbZyHJ/MOU4/TY
20Uk6AfVpSdwrmfLTFqXErjh1Gphk0QgoQ/6MYAtc5eeVmA7bZHFlHQTDNckuggRJ/J6d+Vfh9dd
F4iqYK5HZgppnnYoFr2hFQSgEgkR53YEYpmnOGb1Dxtw+FhISPib2emQP0E7Xhb6KC3kOjZR9t/w
kBNZiWk9q8zZJlHhRXktbbmBw6K/AbLWst7U/DRW2yBV6MpQZqghE5I6imYmp/+aLtzC0fcqGGBs
pvjP7qIvv0jfoga/rr6oa8SUXU8kfm9tqkis/JGX8LhfTLRadXCOiejbbx7CwEdOHakEmRqDXQlq
DDozB/928I0SSwz4dM2g4Ksb5w0GgSMNbbQbGTXs8b3tbaEny3WoBM7Kgkz5hK9Rcj+G8b9GK+nG
8IihOCKaV+5SXxb15r3tFcqNxDZhtIbiArZ0LJC+Udm91vx+XUwJy4EC5osi8bqThO4CFWmzqLHF
nXvz6S9nmvAc+zN8xEVLGLdPv07kbtGMccAJkpVZCmQ0fW6ZDXOY/EJfLCYPgxa4U0vYz/milSa8
iBRvwyvoSPkcRa/wLmIVkuJxdurWWZsJ9hXWsIAgSHD4ezpPF/jLcAa6q3wuSz+y1+9lYXctXjOm
FeWo8ehz7JiHFKk6di2elxlUp82Epx69jBFSBqyj6KlOO8YPIVXxG9dd1mLy4IxNFEwzSjt7DuBD
3fyhQe8HbH0lRpWsEWTrBI9GuxYrdU4DlAOqcyl5DQXKUbiFA1Q37YISwDaGyP43Rtvx9aaPutzN
JJILXtsBE2GaFh2xhsFj8H/D+3+NdMpKm8vGg549GS6RZpHaVVFfIbr0gLl7QfGVJE+RSDbeFvbd
7lENYzUfsspl6n5Hcc0BSScO+u7U9kEQFwqni600F5tbe7vTD/ohJ0KPOayZP9G4zwWWIIUjtB/n
we5RjngazgRLklDey+Ho4d9FKGgrLeAnDzC5Wnu4KZTDDgijz/ZGkX3ylnNwP6jQKSoB+q490tql
EW6gAR5oH4Drdg==
`protect end_protected
