`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
IcYwklQOp7BXpFZQ+a+DpFzvxb1PNTdkN39cYcF8uEBbCRcKzJ6oRuXGj+tbapIAxW6ZTcHsQl3e
jWUfYFS7cfekwnaNsTesfHLZswUha1oUwD7Go2myjubvYoY3gw2UbtOdNQWNcOFGx8UwS5Fk0sVc
oX42bcLYxAV6QQ32la0zQwxtZU4QqNY2pa5XoyusubH3t/F5pxaFr2ZRmjTXhIEtUrGsSBfJLqPA
I4P4BQIWtZzzp8YMUR4FXmq4NsGRnKszishv2UVQyhWNo/7idfZ3qd3n65uNxn9mWsjlikd+7xYj
tVn4oP5x47hX6X8a7+oE9/4gHgXoCKtxGqDD1A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="zPStMZlM0NUEB9i6UNXBjnjQ3ZT0Gu7YHgvOzDQgAtI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 171568)
`protect data_block
fUYf+NJ2WV4A64NUxG265PrICXf/nIuMhvx2zc+kdNcjwrRf1EiWsvgONOzEaP9K9g0TPl0Z2oPi
Bt6trSaZdTdawyW/NgBLGoL3t2cDuEcGkWo8XmsxtcKQ/GoSoYGWJM1DyvQnTGXLS4RC+NAR6OOE
CGHhPuKH7a2hHeWS7qN6pMyFIuVvUTvD7EVP3QFelry6g2rUeYSIrDiUfeaNUr1SOJETGe+mbbuy
L7s+G5uaLpgO2Vn3Bze80X5I2ysrxOnu+TCGY7fgjJuN65sLF/A6mTn+hL6Lb7WaYsTMBT1hksyU
+4nj9EA04J5tSiyUb7r9Idyg0oJDOi6ND48hFdGDbltMfshJmaOI/IpNwQlwBypzvdbqrT+OpeQp
DlsxYeTqSSUkJWWaXUv7lK8BaPq/HA8M8RiRQ9DYRPNXYsiMLDMj0xna8weVn0ExpEuE22YjfaiG
k9T7vKB0rXlaEAwM74eOX7+wbkp/qQ+BeaY8aXkLqMP9RbPgKNO34LzfjqMnQ5EOexbZsxk9XjPL
R7Nrm+2gvLb6nj7qppZQ+wz6e5X3GJcpMsPSwUOQ7kUEV2UZp4UXa5+ZsaszMZJEuMeBbm3nEb/1
GKVgyTF5Sv5gG/Q6qK/7IIKk9OpXWvKGsJVcia/W8HqA4igdQHOELojLronrPc0aSsEvc/iQiznH
JtV+AVimbjxb73g0OcuUMyM8wHu3Lm/tyhehdbN+v/P3mKah2saGJabmi0QHF3ftv4Hnkf9HytGx
/JYlBrE+3Yo793ZbTooeiqqMJmZFvaJLtF2wDmsywv0irqKp63SpmYJmd5TlicaLTCSX8HWW4AS6
ei0sEDoYQb4tFVc7OD44LPhIZEYTpOW7rUKU4uHVI2K21dVRJLJNSLL6e3XGof+Gf0cwOA5aYMbi
NX94GXnp0NtrCb3NVBc4S1roJ1czCfv+rvhG0RyezPzwhuJpeje9mb0s1kbjLlNBObjGfMvUKioA
paSMKeTdo+SiB19oKTph4xsqaRT9MFVFQGG8PgwxW9j9eEB2GgIvSz6bMno0Utmh8/SBLgiDCF+I
yCU6PBw8xPkEQjxgx/78s8Y3FO/0+SHnbbgxPKNl9JwuA3MOk5db1pcNufNBCFx9VxWVYNCf7yE0
VyQhJsXW22jryPexT9Mc6rluW7As2nrqihmmRMOZV2NCtAFGsLIWa/7SnEB6m51xrC84WOrVEAs8
lzs6mKPF4Y9K+CbnrjtYff8O1RlsospUGbf7Fg5Z5VwL0/7BCf3XDmvUvxXAbW2TFAaavvd0ac3y
+P+hRCcPeELE0s3LZVzWlDfTrH0hb4DOasnGp+uENRpboffa/dWYGF7gyLeFeO4q5KyIQc8Ub8Vd
WVO7d4/3cqRK/9RVr5tTNmlvgyfBO8caKe5UotuWQknWZLd3OdXHHpIDO3ASA5HWk+vz/FZXiVxf
ml4w/THsEMDxAaaSfMjNTmClDg3+H7E8L7l7PlV8Y6zK/ZGMiCmQmXMN+5PTvexrp+m1QozFmbpZ
DhBelRiywNyJj6RzOvpUtr77+/GRc46gC/rzlFwUAFmO/qa4eNkGGsGrhqmV1weXegaYPUAts7fw
xuZlpF6DkXoWzrvpvZKSvIU6TOy8sv5CYaG3QORuopMKbJAuVqQ21Inn2VFW38Xi5Evwj+aFHgcn
xdY7mbkSOBwnCEbYbtk0QCGVIVTjBjgOBRY/i1jXmcyM7MXa6z4voIWv+EyOxkAsMzdUnMPj9x3Q
Y4i5HDkgriXtGoYR8ZGkgikKC/nabA6/PiXSAWTJS17tzKjR5o2q0zZdcg39p1l9kpMqZsR5lKsJ
Lv+iy10VVyfteJGVu8gjJ0ERVQMQ7YdhokIYSUOnzmZqrCvb40hABmLUB7upx/uhYbcoPOve7xPU
hl+uo5RS5uy1ExeMBS8nlpFRJbF6Jdpt7DWQMx+I21j5x2TCFTt/c8ZNJK4rmlLCrpuvE6dGWA67
ddK8IcLvM/3D+mtC3p/sjx6aREqd9XYP2/WJE3GY71KXXxl9fzXheACEz/vKRhje3FLQwjavcXBV
0D+hsrEwttzUoDQ8AV3a03J7CuZrx1qMstuJTeyXBdJp//QMqkeC60U0BTnE1XHLfjGt4hxousOk
BFmcdndJP+J5GxT6t8k/ovjfaYHfvFpoyFfK8tZTTbgER1q/YJ1Lgm2+SxSX6UIs27d0YYBHq8Yj
0LECVmkH2gILDBOGIjLGhLa5tTxRezXCDHsl0RUankxRrqi9Ruco4UpPaGjloQyZPB53eNK2mP5P
uIJ2spfI9YJlmmidIDlHmF/aKFllhE+i4LuWMRv1X1Myq8ojTh0BjcXl19ivMeiv7aTL7J/QWD+R
osUx5XaY+9kJHBmDAcJLppZekrPYhwwCzH5tH0OprHi2Gc9LqPJv4nX0Gu1CpqkMSW/V/q6u+yr3
r2aPNeQFoRrshV6Jsn8tZT3bMuKcUc6ub7RBrqHm/Zzh3FkJP54WO0IRM47DP5EBpuLsrnbN6fVg
SdT43/vlc+Ohq7pglZxVQ+g/7Q+j4wRWbBo974TjlfKdWqfAaabELZcLKkcrcdrhY8LkXn+sGqQ0
2d46W6yw573LXoFkSDarzdW38dDDrxhQB+Bja1fvRwMeBpkkEK5djeLgVtc7tcIxAaLjEYx5PGdC
7MUyDnz76JJxGQVDAqdQl8/u6ukH742OOtZPFdaexL5G4qSw7Iako7t7E6AhQdEJz4Hhoeae8BS3
vzbI58J6f/OxKXDPgmbUUjQ1SuQIO8waObysNEjBi8X9POViewuELxFCuHQ0PPSq5w0YrwvjALx7
eQ1IqyrPdJnZzecz9KAHFJthlS9ImGev9OxfbECMEzUXCUFM7rB2tXDmmohK4KsHujA+chV4//UM
/ja2NIjBqMSPOWIsJoL/RvFueHdvBWl8FzP3nzGTCmKViCzneTlOAuJa0ZgWig3T5QbjI2Q/2Yyk
y3wLjbvKe3pv3FJyrvLLLbXclWV2bDjbya7X0z7QZioESvRNDAZhcWGxtAr04WWONqE8ny5LaEw6
0toGTxwziLAvjCNoQZZh4Fo45vYO41dOzr/MAdzYOTTzCLFobsoKTc7k2ZaA0QonsqWGNKbPZsYm
tW8HfDellS4tqfo/cQZcXjJ+F5syV3dMk2OpvknGtVF4iMC187+NbajDP4Mi6rMfdOmXuwmBYcEI
uIwe+ZuEdLVh3dhY83vFZCULjHzEUFxaOVl9x7W9iyVNX53w4JqhebJ0F1YkCUu2ijdkYTmzklD0
q6TIj8cLQK8dtFylKZGsB/VBDlX98aboVzRdqzs2+JYIemKi8UQBdow4RS/WNyrChvuRjaYicyYK
H9+dAJ9qdpSGmO+ypVCBfarR3ewgqQGwgsRRfIlHzuQGbcYcZAj3Dj9tAAw/1Qt00P5Px4cY3gtW
Hga2otfwX2/t4bYfc73PhhtX+NAdYFppktHoMlNL3O+HSdePsh/bVa747OveEi1h8aVLYQuPWEv7
vapgnS7rD+svuEs6cJ5lDmY+ljKvNu9LKYERyX71cvIEuF4hhE41te23aZHM/stFhPlZbx+fUaA5
x+gXPDiCEQ1xIoeltshHX0g/xV/s9K6Hw/T93BdLhn1HohVhhr1lgu9AVstcxrfY8jOFg9Nyi/jc
EWaUrBiyYIlLUAPOYNX8D5/uyIueYOxwfRqcKjZV3MjIa6HyjEM8zsHh8iAOZsQO3Qm/8LeC1RnJ
EhMGpWGEuNqKU5RvUBC6l9mmfGYTLyvjJjEFXgMS6hhPx0W0j3gWk0SLWlQGyQqktXqu/tkDy5H7
Lbylf4ATq/Wd+zlOUCZXeT21mnKSo1WD5O8MRF9AlSOTOgqPRh2xZeK7qB0xTmZiAmMjVW1pLMum
DaEC1dtY7qINkBOJ3Q5ReDC/X44a/ej+Y1J9ftLCwkrXDF1PUK+qXU/1ObMRsRxF65coCMsNwCCM
Aq1C5/FEJgpNUfMd8UsUtXHJ0tK33k3Prhrrbs/lCCwyrEnYh7Ns6BFqhcFhQNakValO5nRMSOQK
O3N6J1UmVaWXIITpkgrRaKAl1Z9y3vVduXBPyAl0bbeaswEoK5bokmSH0NnKyshcERurU0xhITkB
RLLGMcZWBXqHunQdrNv71mK0Cx/4U3autvOqWPDB/oh0l2CcdUfIao5UEtzdd/fwulbBxhBGXL23
aCJr7cJu8Ul1VdFsRScPjs/y7ur5H524FJLR/Hon1MmoDk3elVfjMN3DsKfGwMh/VDAMvktR+zg6
zRsZpp1jOOcefumZhgvUk4ibGCIC1n7VdYqT1qDFZQY+fW2wrUs7PrWT6JZGJpqrUD1Dgh29JFPI
NzT54VZHKaiKpm5QU8zLqbp9ap24Ho8kYqmEJWP+4oheYxsLYi0tAF1n/H1g+zHUiLrupQSPASZD
kHqSJMOUNh5b6s7rfTiX+LOZWZaTkKUWCeK9jLabzjnhCBOi/bUI63XofH/+xYLxwfETBg8pVlrS
6Gtmx4Kz+8JOM6OUTiNHRjKtTQDo6nmzHAAXzvXIVdtOfNobCm8Vid/6gIus7Lm9/KLk0chDAzZ5
MOH5YItvrh/uV6YkVTRhz0mOzPyvTKIy+9Klr+pbDjKgDBpRV0as/kno42glJqhVHlEWduT/InFU
rt4BZTzaMEsPgv1GsOQA5/a07nX27HaaR+fCuWsGw/Fym1DsLSKWclJquhgKiI4RyhVfLctB1tpe
I50Ffl4y9MDEvaEovmQ4mX4LcH5HZj8UG8mrNsSOHMRPkESMMNVkjQwOsGCQHAnN+VEGX/cZ+Pch
cJEI0n085PfX+mHIHDiWIFBr0YCtlfTWJb5iz94R83SMdlQfHxCrMKoMLhbmfY49IX5i+NJpKYj+
ZZhcsQqBPyUKKuZ5kelieqK04MHf7pvJkP4rka1ccBW8WstoA4SLb+Qgz/NiTifwtjn8ukhu549K
0ibrTLkUuf7LL6U5+X+Lz0jmRZ6nYS5NrUksfcIa/JPJp5ZTUoKvK2CqTSxlVoNyiqUlro74+QoD
xjq6JMPF/RZvwCySw13o5op6QsTtwLvgBXaI3gCELCL/S8NfRC1xXSGIMw0xsVw7PfGQay8g9dvz
yCo44w3jUgeOGRHS2LE+KafK6QLGiE1hGM84KVz1YShSVk/7MxQiJ3cRjlJQk95Fx14sKycWy6RR
EsGxXLhpmm+T2Vp3Asf3R5tM80CHXctkH5giGEXQS2IVcNfcZoNS7Vzj4hTMrIRA2Br9nzYjo40z
mYiPVXywL2WOaPrbL4zdL8FBYztGqVJX7rhPxPnKRczbdxiP97vgloXMD0/KsrwfPTN9Nm7uWg1a
L+51ShvmWxk4MaY36RX8cmjNiOuePiD7u2dddk+m55nZGtGizxi1L5nTCFTMWFM1CuodYU4tANcJ
pnXcfNOMfsnGt2YoMrrokagouFVk8tSmdRpVIcq3K62/AO+l6Y2pZqhenYwgxcLehLKr3e2ejTHL
W9zTTCAMPjjMXs7/VKM43lOkzbjkgooyn65Zj72n3kB029oc6+hkG0Np192vZ4r1h588JhFWhBiQ
uTING2X41ZisGw5ZgG+lI6eC1Px5roIsHWszMDd83tK53lTncPFxfuVugCFfqIivMTF7f3GgWAF1
oSxy9A7xEG3G9aa2+/uhIcow3Izeqz4hF9BdpMbPIMafk2YrzlA/ZHWNckOwCBBfObYpWvrXZjqL
/Mrt+xh18tsKg4BSIqXv4vG8F7kRqYq8q/tvCY0caNdWSv2XAARttnLGY8oPSFjYadmbAGSYdUb+
CgThhxVX9FnmtrTweEwn4rB8MtxzInpT6vMDLdjHvoYWImHCfKfPbpaEWzvKF3gci7i8X4yypKXj
mrYOGYaP9xd1cjIsBm2/yu6VWdF0k4qCPZjci1o0+BsVAw8PD3ySREAi5fmI8+l+0Op7DyWA9Ef4
eMGBXR7Xh51hHvfX9l8NclAIn7g299UDGmKygXlBHFY2QZ9q0z3omW1SSdZhg2QvlEmNq7+vjUTq
A6GFP8jl389Tj73C4e/9rQO9bVQtTvlUXqqDQksfrOHSx5bBpLRu/vh0Quvpky1LRxlClLFVnMjP
aEJ1oL3CRxodOacDJjdcadOeu4Y7kL6XVuLn1xk0/htF0XS7YADsJFiUgeOgfmupmXzbXrNCWd1h
BAQ6KV2pEl/cosjk0KdweRXLUtIHrBTPLmHDAHXvdeJn6OhFiSsnsPn9idoKenAEd2zZk3iFzOe3
FZipvjOlHEedLtJwmnK0hs9Yl3n7Gxn+o1oOLa64ZQdWC1DJddWRq9C5NFhA+ASUePSspYP27jNT
XdWeDGT0GGQbYI802gpJDVlOjskFeVtXkYbSBiYtwitI8/LFuTYHBlJWQNI0rqnFF1WodmS49/jR
riIBFGtrYa2Z55XdPmXuwHkx2hdoy01DoML5WkNbEdiay7GrpqVl9GmODVnPFVY6yhnqh/0b5WwD
priwi4QB0H+o7UTgMLOMY3fYvaXOCfZZM+qg9P+/dt8kOUgAlLNlG71o1DZEpdqsgBot4vxdN4L1
wVXkDUbFFBp+JnHUcrrTTLOJSXoT3xlwkPSkTA7LRfFpP3w20BKE8P74LQcrrVS9v2lfoMek1sOF
J0JECj/imGyUFBBMT97WyZHdPsQJSETKSyH1+PwULYRuvBdM7QqMph1zATTeJum8XQLDDF0/33pt
izk+JorPR3p5wRFRt9RJS7PABaQ8WkcfcAZejmt2VJ2Snfb3lrgFFNcsn4pWhyhZwRWV0BDFbR9s
D1AL+QKHcEZg6YnktC9iOqrEGjCS6WIx7MuM3X3z2ipBRtgzEXlMwVbLgNdXBxxB1HxmGo5SxX6R
pqR+ubvAZ3JbjP0ZNpslkps5ARWmn4XBLQA+fsLR9yvlowra/lgjAA5lUA2e6PI3oqirnxJPnahn
xrOW/F4SgJgzHlUhUao9xKqMjxsQApqOvZ+DI0KZBKb2BPK+xKbCRWf5FKkzKxF4ObGGxvwxmY89
KRiI9f4a/8immz08b9emUB4FA3N2BkGorFtr207t6QNQhDLkQIpdUGf+1mHaMI09iHUGIpYsO02/
4KzKLMSP6vVWnFiH8PJzajvDshlrs+YKuqWBtRRCglE4jItoWZEgjpSvZIkW7rIu/iLDKcL2hbIa
rlnrzvJauAozVh1V1Uh0faqw4QLvkJstJkQlLzSzkSTvU7nXbTRnl2EkwlY8cgSfWzTo+1LkPol/
WhfD235NhtEbQxIU8iCD0fTMScqe3FdgHqVaZhcdB7naWum+dqL/A9d5s0ZsEMEIWlGDQxuHqIRf
5aZIa3dR015v2mBkhUc6FNgfYhFhnM62ArGvWQNeqH21qBpgxoaj0oPK7H6sLmUABj394vMiVwBZ
bH+ZVFgNSUbIbNhN24vAe5ArScHaXVOR5wuh0CHduH4Z0xcBsMyQfGU7EuJRxmZS9w1zpDhMiXOw
wvZvfRjAB6x1sHaMOmoMeGALTsaNVBH5WybWMORgzCagyxZAq8CXzhbKiIKmIV1PnkeRecqrB6xC
7ZWHI/rsmvIFT8mZXhw7HG7WOqEQLki9qvKhcbRCuJbbSub0c2DmJKEVvamb3hjNHqYwIjDQjFGx
6OjCOlfJCfMtNZUISh3yhd1AVETnUpoIDd5LL8YZNxsj9fZ5n4trYlJOaj161arHpjmMNgZtv7l8
WCm6AmezP2JvgupSF6FTY92pQsuOMRp0MHSgW6iagg4oasdiQtIwBjmNgyFi4RaLvyyUnmiO92Fl
OqwKMhDOKhh6tKT7iDkjNsVMQ6Jd+78KU54xWjSNTy7bSvhwuW5FlEa3yLwkcU+9FhNiXFLmny3o
uqTbFT6zNc4DhnxKNtEkTsqKk/vJNHrWpuZndToUx/Nz5ggqlls+EJrX4YSaeapgCq9FQ73tXrdn
X/y1jC6mOZnFEb1ND5jPgAmo2tXIVS2rn6IIvBNjsfvpFM6D8Kt/j2Ki2UI42cZfUj72uJNdXuwH
e4U0O2H71dZfZ7NUjiC4/NzAhehp2Y8PEnITkp4q97s6iH2MpyDpMb4lnc3OqQYMHYx0BJeoqqOV
bmOju+AFQUJCBJOqypv5Cc9w8uZvAReRPv+1s3Qo/qP3d/0vsT40Wah9Jw8uI+q9bTBiHrx6V0OZ
8Ka+j4Pqx8VyBj7j99MZsA1nGPKtbHA6EW2HDA6Fioq1D3woIqws3Ry+mYH5vgOq/DWsy+R/uopI
OEX7Ircu4KANEf18CSu/ThS+yOQPakNW4Yno2O2iX8GV/YznSZk27ZMrOeXOBfKnTAKRVZsHjAVj
LEY5mf95P620okyZ64FrbMUcU8gUNrysZQdQcYB8Sjxpg71RvOx1o6XjpPTMNWBWzhNgj1Crpk8R
BhIUDbrptpLZhJa1MDk27aCaSbTnZMOIQTRBF+AvUzvs1Dz37kk4Kwds6dC8eU+zJHzLEkgToWun
BTJi4YFZZT0Ko3ACtitHylJXQCfva5qhzyLWXvJrWBXyEXJH/bG4FIgGGNplEzW42zDFBrtd8j6Q
TIDbqwatF0ZX/paM3up/9ovA2Sd9Np4tAgq80u4GLwCitBJ1Es3mB+tkZhw8ctGiVz1ZIhipXIpB
ns8WTnJkg/c+vHkwEnP7hfqgFuO4WBKv5sVB0/SZlWtvfBo0+HV6R9980629D0ZyGTDvYXisAq3H
3FgoL1CqNBZEa9n3VN1lyfTlemleGB8MPRYLbOdAfbq1dDT8AqJVKjPCWqnGkcLvfD4XEaFF8aUj
EGUsqF/1rFPeMNcK4KEVuopjylR10yYbq9Tr94sCtgKNhNwX6ItI1rjKpFvHRdlJ7d/X3W2PeT8k
BwSWnR6xnWM5c4T+zbAmxSny/NcpCyMa5kJI2hib8oQSN6azhDuem+RdDQGvOoVo835tH+p+DajD
X4/HY3FALCJvmX64XIHuigdcE5iTO3F2iHFxsC+QJ7B32UUld+tbhZy5hekfUqATkAyXGgwYDCWk
wRxyFMUlUUUklst0GsAuFJxUrDBibzF8xet4ZXMXTWH7iHF57xJjRrUATy/y+Cqj47QMCd0k255j
7QIFchO+1ARZyox6Jx1bWBruv+4OE9RUlrtRJZIL+MtG08j7JQlaBn3uvrlqQpLvbedB/2zBQUHV
B91AgE5LE5dVHl5aQC1dZg+TplrzGOy68CsP1ablvtGy5nYZnmXA/zO3pi/5MYkh5VXLCHKSBNjM
U43MvTO9eMJetKemxXKxQBdVbhSk/lfmk+KQvBx07rsQgG190WXDdJT+wlpS7tv0zAVa1NZpy2Mm
+B/2IA0C+v+6/qtSYCsmrOVVUvuMEaQA6RZkOWX8coKGRu/Iz5n2jyP4l1kSlNkdb3ttyMpJ6HpT
DmiioGlNKW1Q2cT6QJ8UFAqPtdxd9xuh9ngguq96HfZluSo5ZD5NXkO8GgAdy4DpCxlyfyzhKcVO
W7FDtI+o392FEMsLGXsmkolnLzyRRGaCgDM8jKV+iWvaXhI7OzMbUx8AFBL143iSFtaOvGEROVzk
71gNQ22mNWjhoCWC8741u72vqFfh+y9mUM6AcWqCIUwCSYWbQzU/xbe0aAKCnssoNPYtYVLA8cd+
vjN6pPQtzVBZGt0Rf3VmtPMCPCfdV9o6lBl0R4a4iaoyCTQuACOJm/P3IeQbSjPKen1AVkWKNsli
5DADGimAp6TVVLnfr+ZMlVgIwW1thpgPkYL6aQ5CUmyk5SfsJqy9tdHyluClINvFrlPnuH8voNiX
GMguAV3mpEZPaq34eV8lbSio0UQ/OhcMuBCS/xItVFTuJY9VewFznVdEENCnriH9Yntc57LiTa3i
gzol2GpS77636vbQSKMMJ+Oysmu1A8L/cw9C/P/dg3rX7mreFYBZwoLISQ8bHEjtcUc4zUqBPBb1
FdlT4F0e91fSCDBcxHuaXuZnfn+X9MxA+W6F/NnAQaGf86uGDXXPrFrrs0wZY3AKxHuw46TQA0N1
rM8PEa2bYgIW7UIxIF0FJ4U6RFTNgbdz/cdXGy4qvqHGbX7/yc27irZIr9JmU3dKIG+VnXMel3VQ
UXcWmB28tPbBzgjHfTTiixKCPzr3rdBCQGS7UikeFJxsDkL/nMEqNXYgaq8mmZ/gwud8UjbjMoVv
g8TfATQTvExmizKjDQymjxsQmppXmadCXEUzmS4hEXxuykCi2HFnhT0U6svAU8WqvJiunm5LQT7D
78yqchhj7MRqfzVz7esYpfixrS93t0gMDdyKewWr8W7tMZ5Pt3pASBshka1UJsl3ULqWFFyxF2Yx
Vr2bQeyZ7ni8CKoZqqUto9KBUX3ah8dSy+WL/uoD5muLvNBYMoTsZaZnY2+/Tc1izP6A+QAOcwFD
uQg6WohmmF+O7CGmX7THVvfmX1Ikof2boefhGHjD3PZ4hDzfPxAvwC7HojiLS08Hz5bZboSsNn5U
rapnr4Te+5tvdkMbtBkBQ7LJDjdTy1sDpYMOAq8dlLt09jXei7uo88jtWbcxh4DKFGHVyBtJs+44
cTWKHZgowc0RG7FDI9g0MEMOYafwgjpoXjJhLgaZwvk9f564tkj2BTB1n7zQYwiibU+j4N0QViBZ
NWCqpJJbTMHkvPoWNdOQMNz5ZWKWtmD1TC8d6dFdTp3Uy1x48LTg6Cw6GmlpZL7Nx6skStGjAYpt
5bLk+7dNfZxUzFPtTA93lVG4jFbVk3XbXlPYzBGtYaXuY27OxhomofL2NjnCJohEevK62hgCTW1h
Gk57C3jDPR3px+8IVc34h2guwGj0pEjPJ4cSoQwEdI2jZjuoPHrHTQrvSMO1bEBNdqlNDd9f3O+N
oNIFIL9l5Q1oS/UpxRggukIVhxi6Z7PaynBrMvp5i6oNnPNqNVlVBvfC3Zj+wtWP93j6sk8lSzIl
QOAYOhVSY+7WqbiNJwuB9QBrWBmlxCaNe4Dr0qQGN0Q4RrexlqJUJWo0WdPjE95PNjGTveNshwfw
5QmBxtuAHGq/PbzmxLZVhoykym40mkhq8uthdxgIMNCpnCHrVll9DXbXvsPiSnJhOHfAI2seykC5
88E1EIqSDhOiVIWqcakQggbIsUkPzVe466FydPvgTmIoIFZCCqPVMfzsChPzeeIoxK2sZm9jhFCe
oawfqysURIQpLavp2IAs4zbgIfT9soY6NXvZb8Jf9PsVFhLxbU/PdMz3feCz4jN5n6G7C852kame
oJ6MK+FdbHJ+n/dQRh37GbfBHv5kwetD3P/Z8s7DAbalE/N97oK7jlmFn1q2gI4x1S/M8Qw6KTF5
o+xVnhk91htkFIUdxsGK+Rwcak6KtxlPD+T3b2/gQGU8nWOLq41JJ6kz5KU3g5vAKMYvla54a54Q
BzO9HPVUpfe2SfqrFcG3m5I3H0Ds8tudhL0wXbMQUvfNoDqvRERg6CX+Pz9HlIGymSMkzO1c/ysS
7yMOOupwSizqyau8EJQyYv5qRpZjmv2H1GK9lYkJ64ptfLRu7GoNC1NKFdOi6XMWQJzHsLZwEQSk
N6i4Qny7fHqnJhtrFQKm+vTHrDV4swJFy+tY2zQPllCOEF1DJhxO4zL/U5v3z4HKn9Piv9U1AQ4J
LRdoPnOU45Q9ld2V7K666LuGZWqJ1td5w6CXnnDr5zAz8Wz8n0XZVP482PJeXDjN87nwwI5GONoy
ycc4utQYnhUAUv3s5PybEYqvFoHAKXHYTKwhy3+sUYesLj5ZONdQO8ih/PtGvG/XZCq2tO9qeb6t
DmUNQLqp3aj6rWyW0l9xc2fd7SX8nDL4SGLQEcfU5sIJUDwOIjZlDYc39KMI8dHij1uqUarbdkrr
ygpNW7StsaWDLjuhbIWbYCyfoUSxAP8/EHmuc4PSUmiZjAyzxb5ux9JLxDHSu1xO9ZR6pxtE7VzY
fEtyiBKwSt6e03dAaljeMgguASbC0ItAkS68hWg5MCtubZttyqlimiPLkniID/yEhZoZ0NKSCtol
QxwEtDU2Ggkntbc+O3oaSdRBoKImrpp40maDkrRgBMDZ3UJfmykqdJZq+mW3lciv8TbR9YrlxL5W
7Oo3HoaiqaFbDgpuMXasqDHmYvXBf95b7FCenm5dBt37iWn3zsQbJmed7CUF11Cn0Cs25Rdh5MOn
8oTWQKfYiH0UOfgdEpDlfeEy3EjWtsDiO3UWPfK2weWOGo6Jcv/h0DtdxQWUxH+tc0ZTykQMDhAi
WJ/VXJX4ESa/nBGcKmpacvHhdLO/5Yq75bVFAX80CM94zp/uTtvWJFFEPemNz1jsUzpUDzdPbMn/
RfZaLcygnlvuSSl3UHKwN4zUHBCNE1D7BZ/rzU+PaR67YArgA8ueDKR/8RkX8N3JfZQ8qK4rE9rd
Cm8Uudd/FqP9f8dTResFDxyNXvDU+0NgLxO8YQGCjJCQ3Y3vnD/rFI5NM50yMImRHUyoS92h+YnE
y1FlmTRf1eFgGspUb2t+NM9hH9tJjjf2BOMPDT/9f7Z0xSZTFxaIiSg5oKx2/lp+lexRACccr1ZU
9EqVv3H7vGoO1WHT9um+aoeijNmXvFf5jMGooeKn2VgZBBBEzo/oO9uMU/HhgpCfeXYmTDJqoqJT
aqdBSPJ4pJ31sAjymlAwjn3TUusz6+/h4ES9MjcixX81raqHLOztLVCs5tjewUwfl3W4RnZ0cFO4
oSbiVTkQUbvCfBEsDXsGoqVi10cLQ2Vh6Of1n08dXXCN5HGzRbSVfZdfsA90GAMV6LL1qlsDPACy
ejXH2ZTvkT5PwPYjmSrPlGNpyStirMfVe/aNfLha++hs/geBeZujhz9HLkhUH9saViiRc7QPjFkZ
W9cDNObT928jSpIAhBfDpeRPsXkl7XYy8uKAES1tuDomcBjEsQai4U9yo/b/i6RFWS4KI6K4lib3
nboPcQPbmbhDtjZ85C8g+QV9pr+rBr9hUpy4CHSKzZz3wcHL9pNoSspS6RuMifjK0QbWezsf2g6c
V4AshD0urFuSwSGBR9MWQi0PokEzlnl+q9Upz+fr/0b4I5di8sU9X08ubCLW34Iyag3kxeygO1UA
J0Z1E8waZuPwtsrKUGJQHOgcp9jVil0f+6ksBxzZGcOpkcRjobhr8jHj5W1Nrf3pq2xBq1hLhTzp
pc5mHUKBGzKh3KDaOiQ7DhFU8FWyD0hkAWd0tuRBV/yEToPtRVJ7NAN/B5ziLx8CJXavpDxRdE4Y
4QyB5h0kHWwuVNoyQGmDyNAykCYvWF3rfOfwtOIVu1foE6d/w3AVgFgjfp102vI51vHVrQtJL2Nb
WBX3DCOq+4Lb42L2bQHtMCOFkggXbZgV9LxbksyOcOL1/6xw8Wsf9v+DF4btJKGR02a2ijuPVxWu
A3l09crCu4UUY8/RdWRBdZGtPz9cIhclP7YIk8rX5IknwmmuuObKYH/UNj3AWXgLpuT/st5uonVY
sC3tViYBehg2ONnSm0ZMjar1M24j8SZg7/gyFU53Dcvhn36CN4QvMjbBVGpCZI5x6phkFPvSKENB
BKEfBdKM1LAz5NXIImV6LfP0Kx4w+2yNzNFO4MVv+QNVyqGsCCdCpIfkBQIuuHISzlqN2ZJmIBSE
DSyuMAPGlFN+qYv9O2rNgbh2bbntidCGZnYcfC+EbFx24KxJ0QIlEQ2VnWw1JTSPt3r3jqdN6t0f
Zl1fZqKSETK3reJB43j5O6CE441C4DiOaPxZw7i0rLhC+R86sPre3iBzWYMrFB1X2yVImdYUhSyv
/ujiVTx8UlZ9y4X90fPVC9gVpnwOjVSyU4k7Zur5sVWOWwwsahvsQq0fMCyJ/oyYDRwJelXJYBGW
miyyir9ansjqsFhrX0uAv21GmA6e/U5r8jsfpnHqMxd1lanR8MzC0MsD1Hq8EaubM0QGNaz2gUOG
buELaP9ifFnOKomSilnj4pXlJKRBeIIgaj9o7jyWhXkCbnKiWR8FhAYFJmlvAk1UFvEC+wk904Yq
5v/1DCQX1Jl4Bsrz0VjDrh/eVa+BfX70MpzOwMCXmpPIxIcOS9/Vo6eO3UzUohJqkmRH2x2WR5M8
mRF+2W0YqqyueswkDl/sE1tRmuCOtPuMN5hGMEc/bRQvfkKs6wjgBs6bHVqvBuRoqcRIRUBWP+U1
dN4nFcuG5xnF9Dv3Nvc3HAiz0OujWq1a3dvyzk9SHI7zxTShzw8If4nw8w4Iew2oZ+L07R1EzYsk
p94iiUCOQJJXsSget2sLYReJhMhwc38hyjgzKWWfpxV35JJsmL/JxWIgZKiiALk2rHQ8tlIeGr0q
7NlhQXEG8CnPW88D7dK5oPJgoRk/fUC07pMc/JshkAlxvWZ3s6p/F+5bZtbEiJHP6hm+Ub5i7Vcw
Gif6WuXytuEckQ7cNSGguUx252Q4pnsRwIjF/YGKgm2Lsedf+YTQtgwBQ1H4H9Yj6QcA2KstwDvP
tnSs+XQizv0etpJB322qi89Gmqm/IzzH6TLU7uIGNXTbMrmIY7AQFvXRSwj+fLcn+l/h0dJ/KKEz
KxJ9L70YSMmv1S54qVlB0iMHhZsq0AolldjcOUiBf9ZRYMxh1naeD47Kj1YMvdDzlqdJpQskrSBO
JQzzq4li69yQPkCT5W4Oe1qJYVf9SsntZOkjWh5ztAWU2ZSVEnqRAHKiVIIOgqzYyj1CvFsLrEs9
BfTFwY/PnAejKEuI42nsXjyCDHlQySos+Qyn1K5rAOWkWVcy6iDDS+uUZHiv8BuPH5VmFTKCIPCL
g2n2Rl7k0cZk4J6tYWplEzef7YV8ZpnJPRNnUXPvheCk1cJ5BJHPDQUdFAiYRGVB07V91ZmS4z5B
TM9vp54BqFhKp7I+sSoRqJ5nMcHX+PDuWnouVKuYEPDl6kOnELjckYEilhkqa9ZJBSgSyNGlLSM7
mGUvcMGcoR9NXKp8SGItXNHcCSgxubgFz1ZRFZbzCA/g4s1nzq4TvnhYgI6oeq5Uwhul51q8iypT
5/7Ifi2WDPBgL51HBSzu1+bMo43yyXzsTzwZHZaJxXj9uPJqnsYUin+cg4J28qnOcP/42BdI5XMg
wPfytBTmd7h3NPmJ6kx/OqZIggSjr2A9tiIuoKPVmWUjrU13zBQHme7Rq0oUEOpSrsbocmZHD0cQ
0cHDo9oASlSfS/96uRH+06PunkzeTrlEUSYIEbH3RP6ankih9pqUSLwxcbtomdvS2g66bIKU/Mwj
b9RTNa83NH8j/zYik3ahWAIwWMzpEG7cTeH71559Afwcg8+yjhHWrSZWzbJ4bFAR47FxHPjykYp7
y0jxIwehBrPn1NWD7XViOhjUrKCCE1Ip4EA0ii2H0UPEd2IlBd6H9RKfL1ScLretDX17YwAoGS8q
AawvRKIus6DwqpnTFP3z0Os1sZz1dvGotW1e9CRN55dcI0fEAfdl5bBRDiqfrk38dE1H4G95z97k
uS6KC9Mv7IE4ymoQPFkmW1Qt5DUyvI/xu4p4WF6dGXjd6HJYFv7/l3FBV/7cWwNGNhCM9qXyod5F
/G7rX5ROhh0ln/bbChQE/Z9ZFZY+8GY1x6hVsRewtOJcJANGEoqbyELb1ZTqTv6hgjTH2lkmYzM5
j7PZDj/leKKvDBYihsPBjCz3hj1TohKBAv7EC/UisZz1A07Fqg/axxzw7jKNIB/MF8laDKC1e6kT
ltD3FGRhinJE0oJIeQrlSPvyMFr2M4cfa1SnzeOuFNS/dd6gZHrViqAt5V9vOBnK1maASpYBfw56
iSBpL7UDLXsJcJ9N/Nq/Vo7dvt1kww/xayU8NvuoMnbuTYP8UPDn5l4ig0PuWZHT2tf+8V4/AnOt
stzvtHXgiX+E1gAYxdJRiGZLVNNERUq/mq9Tv+ypeCQ8HCcHUVqEHLmo19yt/55ULZj16pt6GTrJ
R5amUl/3zx3z+9f4SMp3iW2ZZgiGbw8YzE/igsW0PiRtpxYJY3bsCcBQomyyeCVFHti9VSdreuGu
KjwBpEvPfamzFrrSdMzPNUZttbSTQOipT5jYZyKXOuYdk5i2NfbePWX/YlZSarKbAYazROkhu5Bh
LZRgVk18pK+gQP29rI4s9oIpdv3TYGnLxs5KhCjQpUb9OvuJVFqwbjZT4C7Pn7W2ZJaIgKaCVYKO
VfiYYyPdsXnp0jzM4SKsDiGWF73bg+T7zthiK5YxzrWy11pEi0HPvYdOpcAIQDG6v+0RP1cuNOvy
5Lal4zPWvWjMld/HXhls5ycNiYx7Lcr8UlhMZnwNzriTJlxbt6YfO4UfgnJGNAz/4sjd+Cv/e9y8
DKYY4cxr1eYkxkYRUfgpt6McJJvsKCUHU6ErHOpVks5kZzMkg6CQxMQJIO79lPU8BoWOMLb/cqL1
rD6+K6PZePS6a56U4NmB0fvL5TVW4cuRXRBYuBit3nJT4LjU0LPWCjv820saosPmTMGnRoLtuEtO
5E4Pf3bM8ivtqTYRF0nDShINKvLzpZTThbJEK9BEe/LQtXqf53LAMM8488ijoQxhke9jFVcu5GHA
MK/SnYSn/33eO1nFKLR+M6iCzv1fs3GU5vqapvjZFJY7d65FVe8FtE67OpRMVs/6h1ULcI4FCp7r
PCr5B1qF1K5DKa4UiMz/c3zCBHZrtXxEmFuJP7Yd/PcPnziE+7knMpD/EWDSci8eD2Xi/wJAQ0cm
OhbMuUlbB256wFUgCumr0JdETiF/gAbncj2sUa0y4xUNMFb1S81lLpHYoJUw5sXRadxxy3D+ITLx
/AbZgCgWMcXxZjN14u2w0YW2t3CjQTJcdxkHZOclWixMBiJQhju0pLA9W1s2uEhD9f8c20t4UODI
MXTX4afBReQT4ohQXKpiLYfTHehFvvrfRJgb0ZOKk+SnMGZMVcsy4FleIx3Gjp4a1RzHn8E43IIS
r8PQwAKD8uqBjcQoNnHlxBiGf6M7/cha9Blb8MlnmdWh++5srju0pDmfGWdetfBD8YaNmi38wqQu
+ILeUzmsFq63328d44Fx/NfKqJiDjY5p2fq8VBIFaxo80JCVRmZvr6PupGlMQ+O3QbVxpciRITWg
QuoNayRAF7BZz4f3SiysEvds7ChjI8g7JweOYfjDcRoA+b8XIl4I4ZZo3w1XqDDRPNrrWvx4T1+0
53gWccw/YLuqr2LfHorYhKHoYb1hDBD36vZoGmquKbK9uLSQbPt8crncvjCfwxq1FRMCzZKsUEUe
/aZ4l9lNCRrivenMsBP2bAQN2iU3s/kZzEd5guEhPErozscsFULIcZHjczth803wupP/cD6ZaWwP
SlZePJgjjmBsBGb8uv6NwydgltcTMathv4GnrKEmsjVS+SssIb4wHWSTl8W7ArTkgPyagC8RP4oR
DB7gH+YtW3N+VSzj9RpbpCsQO3OW8ODUEOrRY5yJoPpwF00RSg6Uo2bddyLVKQcWcIKSbOlmnlo/
1mcmrHNP/GsNKVhtP6r8xks3kSzzIRoDMxRHdL/CXv4SM6LGdT1VHF4JBZCKt1Qy0vje/JHU5VhZ
Rq+FT0CyqeTVl56ulvveDK7NivNb/2HgzZjy03XvqPcdzqEu3N+JcZ2oW0AIyZ5SOmalY+EcfEfN
FpigTh9+N/AwiNV0ySY7MMbAO/3gfRtVox7mV5+lk5o+GJrTh1hpfAicsfrV73+DMbb4BfwILaMR
pCRbi0gOvy4bb4xsz5Zbbpk05Q1q5dakt4OMT9/dEtxXOt3nttKXwIp954xCVvcBJ0NG1UfrA/Oh
yGtP9uYtTQssLl8kmkHRje0JWfxLwJBn7FX4JNFhrXWe6t50wN9x+Km1Jm9MUiIyMhl0beZr29ri
l9TGE3K0xg6D8pO8G1l8HHXLtKPgc3xRpD9NUg76g+5Ay94zdzD9KH4rx86/r5AqQuHzlbbzKvZY
oaXH4tpqoPm9LzQaoQ9zZX2KAqtiI4ta7+N7B7bpsjasMzkn6SrudiCSJK5A6ny96Ch8FsXKJWce
6RZJEnd/UfOFOBA95j8VEdrF93jzSL6FcAQmVtawvRtgzvlsmsgtNfJ0P6s0zmZLm6cGOw0V3E/Z
wQFzYMYmZlNmTpABkajO2oX67CakSrXQAz+oqauVB8ta2+gRjqXIMlnsMNWGLFwoekpkEF6bef1l
K4YRQiniVGIJZx7QN6yd5rfsmLPMAh3hqMX4qqYDmTh53ffmm8o2S4T1AP2xvFkhGodyQD68iuoH
HzWhvA6/Qa1YFGa7WfXkY2eEnEQApKoPqhmGfVWCavR88ioFtq4zQiEah3byTVohjfTAxQM8tELu
YqSWH4IUYh9hqYmCEojPXcbIHtmb2M88Wvj7GXyvuXGfN/YsEoF60uy66QTdN3tes6/qNp/QSMbZ
ms2bWvmkeYvqeHO2ZCTlkV1en249YgJmPW9OKoi32dSuVxQ6ehJweJxEPp4E6EWGM+305fMhkxsZ
zB/EvU7U7TuH0I66KFMRIALa8vuNEwmDqMSInF8J+kNjbK2XKE/IaeVQArRWemJfA00A0nrYDeT2
AhLzb9tI7X6peMPntyqX6WZhsNnwr8p6jXe0apCJH1bF1sFQ67ue81BI+kZvwB7J+YINt9eHTdPS
JefaibxERyGqcLIJa9Et5SIH1MbKvle9vkO74Z5220cNTcGvYk8b6TODaPj+BD5510ipcNlmosVZ
jeGWHaSEkA7zh01Ji+/RNCcaOLV1WVapxyAEX1cg8tPJe+UbQBNQX+8xq8aqJ7PlTcObt+Tvu/uw
a5DYtURFJ1Yilq41fkkHQJw05JSvPXkAG2c+6mSqwkX/dLl9idpGuAuRUr/xCZo5ZH3h41KQCzf2
WT6olyyEawnGSYRrhSWeGkef6HU29bG6Ub5WBonrct6SY9ECsVQBoKn7jITpHGjG5IXFxnh+0euz
BIf4B0JHMrf1EP5IcTUr5QMMCE2oRLMxH5LfjWanmSg/K9VyON5S+ECI+gpIAxr7XbbWXSykZup1
scbKWY3A2cr6NxwHFTEx8v6Qcb30UnwplooVUgYkZA7q9OP3+bqdUuIy1Qp5H11v/HvD+XC9L2CY
EOm3gtLwOhqCYuRQuHqlJXM5LQegcSz+peQNugPmhUZFKMv77G8rRmHsPbFDa9dYEW9MvBvkqP1x
yQQUdhRXGUvRiiHZHW53ghxtWibo9u4sKTDpq9g9Z2ENbhGAJdF+i04I7e/KdgU7UpR0TfEi+G3B
fNmcaY2UtYAhAKWiYeDznUJZasaIi5jQgRpRit+sWRd+ERAN2K+DxalOLi/gt3ZzOcNPLKJig2AY
I6ImglvctIRE2RCIc+qe5fWdd7eJYxHhrC11Myq1LCzpzcnKwn6gN/QGQ2480b++C5UxFNPHmOPR
siZdGGwqFPzzQMiD3IBuoGk6uScAJGtaOfs+rkkSPXuAs9kA6V161707kn5GpesE+feaDo4zW5xY
kUzh/IHCG+0kBSb22FFSsI6XYTRRd/Bo6z+jFUNjwwlrD6O0a9JjfORkU7worNvO2PbZALon2vvI
Q0rmHKzNCqje3FCqthe+sFucYRrLgy2Alzrutjx1iEXWq2k+CT13OgxESzah4nYMfq/l+JiMpP/e
H6wTFcwWbXeJ7OI+RzrVMHYLP6VidaawNMXME8DUYbWkXzEpQF9Id8OHctdJ2CByRT/niwGowTtv
6EBmtv16ecQ8kJoA9mK0fZ1jdAKm5tk7n+utJ+aEdG4PGOHQSPDd7ZtSfsJWF7nn/PJ1qI7qPWiE
sTUFTaN/3Hh3AzRY91GRupuRgdh2SoCMsq6y3MbB3Bc1tb2/I8Cs+GYn4h03Bgz1/NKDYtDaQoCe
mIG2JYtofZAhR+Z2o53SCMwYuG0wd7KAkWdqvxUn64WttnwJg3j7smnXlC07ZK2YusUvfbns5gDf
YsA9H0PKLERxtaMeSMmRozM+OWOX6q2OI2x1ouj3/rLCBc8+mznSxY7WclAT5iiQaJFp/5tNRqZb
EJX1EfIRickulqe5CwO6cKOUelyakTp6AnFOKX6xt+IQ7557PBpRY+p2rlbOkmyKzETkDcQr1OX6
9NvBRR0v/zM/l+BtiSUJNCFYrhwQMfL4yQMJ7QXFKGGl6GxF8z7c0GaX4OQ9ZcngSy9DbW7lRLjw
hqt/uxgLvWALJlY4yZUHXt4oTD+d/QdNbjaNmh96vioKFHQ/9n1yybC3a5fGp37HKpmCw01sOGqT
C/1Pis1q2RNEFBVu1y6hpHXB4I10nujc0I2Zi2djdi4Jg1TvLDW0I3BACsVyLqelrSyszpGhhy7r
wHq/8Yi+mfuq2JuwOQqGQJz+bo2TaAWciZnBT5nCIplClQ0bDPdfZLsSui4norYyUzanrYRtip6S
JPZkZid7E0bnMi2I6BiXBPrDrSc3HJI/V4ziM/Upur2oBWry4RDa2VJvGyjwsfeHULhse0jj8HGr
OEMS1N+eXAN5lc+6gEZFqvmIMpe7DBeq2VaR1rd0FLvd3mS6HsJx66tNw/wyk+gc+YhXUYa8PGeZ
TEi2hCxhTDEen56uQzs0JUQxz++/Oc9ypBQH0omtZPwNypckg89JGlxo+6BlG7cYRh1TjJhHLWSL
0kTHLhuUBqRGFCxzGLlr4JB7BTnQ/dO8bG9gHIinQEUy7oJS6ujfVg1wYJ4D1YNgDXkrhUeZKtKq
ZKgP0+B4nRMIsZg7DFQXMI6Pw8AKnpRiQ5rNeJ39eDt38NOBMkhOH8QOhUKGPbTGbG6U+bZY5OSa
6+jhb8HxkTfcv+wRRj85legfUKvsJ9pg1I9mBw7SqA53o491AJlZ6MirYT4PtsRsubk7fYiKiuqW
c1GGvMkknkV8jYdo1/7ItHhp/zDfhAHAG0tKeDVTyfpROlLGDO8qldGxesQxZ57U+jgrmaUy7Fg6
lrLqnRD2rfRJAxvhpQv21rcf+zsNnaTtlm6rj0KEmgO3Qu53XLsQ63YnNk+pJjWIFj8OoHRs5tt4
h9j1QaN9JlD6mhZNYOSVxPxXZ3T3LIVNCxjQBaMQAhcJEuqe4mBrRa2710bgDudQgeDCT1pB+JHb
r5VQ4LK659BJx0vFb0EOSHUWUzQ5Rqhl0ZyMOzR8Hp/qVRlIT2L57KHQqLhXuZ0ZSdUKfpbCiBhQ
5EUfqCgtgvU5KIWG6e5mdei0yOFHdduUVZ5j1ojuZ88JtZXfbFdqv0oiXUdOMnGO5ewvnAubatYa
NFg5CtCXjnXTjFYJnMTWaEzH0WThci3azZIbjl7RVOFAlDDyQUl9vkXhUMWm9sTHOWwKW//ZaONd
OYhfEQhlFEhhIS2O3MV4It0EwyARwHOVzKSzaRP/1e0dS8xiZsfNsHO1WM5j0EiSc35g7pLbQOUe
HTLoTYHU5MsaHmnIV0lwFp6yWpy50GkZhMrXoBO638ojW04dX/2s61Qg8Pvii136+0ruRSSM951l
iXcHVuaTmvRa5WBdELRN2fOlj+Zqe0+ePcjjkXfpkIgYIdeR5f1oCLPHVL2iKLUmAcb4fVWylpSs
O4Lfd273P+K3J5WlMPjSFTQTs6+dknFUpH8jkW+57ozOUgMUlHGmGX9A6GxoeBXGjJiF42RmvO8L
cD1XSAtjbdx7rWnUDqHv/inu5pSGlujOfJChtxeT0CqfpfjNxT15d1Z2BgfgjJ+nFrKkW8sCaMCc
gSvG2qFomB4Dnpuv3UVjQeqnOfON1WfiuswtmJ8WxIma5Xdy6vTt2AznC4PW9H/NkXqhZUUzHC2P
7xEpS4d8MwgQWXSAKUjeBgWnnu3dORLbV9QozOj3+pYDGphgiWXBBgNZrwh0Ja1PkRRbjVFNuyn0
kMpmAQIJWbuj3aVWs9xBC+RKQ1BH9ndEodpBsIAe/eoRKVoyO8SuRlwO3S0EWeoYSPBMd6hmBhu+
4pN5DBx0MS9nL/2mN0tBeprEKXhlWBUs6ha+QhwPpdz8b3LYGdnsyqxlAb0aJG8MKuJaQmjLOtw5
UUgUsvDMCbIrE1+mEhZdBXIEpdCyEp2LeVfd3+SyUliA0TXnoSYUwbgANRnMUNiKTiRR5J/OvWfd
U+T+gmts9HE34kqChu91LXTZwYBq8VQUj4TQ9hGoQlcV4LddcJLY1LRaxvTbeg6VF8DqUo0IY0Ev
dgRlQuJGaDxJaxyxXncXR5mGPSg3U16+4K0+lVzOOZ7WcyowhYhUFs/f4uL20oZ4yH8zgE0VQ8fU
E4vkcob/HY2CrL2mGxZO0ZTQeFCpKFC56qA07U/bOK+E5s0WRp02MJUaLSsJbt2W7XO7M7HNo3XG
voDxvPexg8SOIPZemhgNtLhfSdBnDuhRwUEeK9Md13xYmIcMfp9WQbi/1CpZ9i8ierinmXdfcQie
j3F8Bqk+oZllCJ1EAIcppAaBrskIb7I9IXBl1NXjwFeOL4wwAORsfPZQ6qKNO8zpd/8oiC08BRrt
blzAQk6ujOgExiZqVg0bCe72mGGMZYdkHkXoACAuooDnLY0ScBJRaypHC+V4LS1mSOj7noOd3cNB
rkyYE7tqvRpkdLBCBwymPBVGTIbikW6BRZPrqA0Tv8nZNAx5fv6Kjsz95q8DuWeuFnV57My6pBcL
V9Jij/3BVx4DO0qVX2M5NPJqwOriKKPETEVA3NGi1DcLhuMu6ilHuwb6G4zphNuvWVSbaIug3Mgp
I1yHgwpuqufVJtejq4iT7aWwUMEaZgXTehujJvSGjWdVrFr5YdgS81bX9JoDpFMEerx9oGPEIUSj
DYWffdWioI5YtSx8wsN39wUm9GkSHCWtxxAVAbNvRbDmDqYRijFtCWMN1MZz/2g8OgMe7kMPUzkZ
o9dzwQMHqcrBeOU/KX9UvorLWDv2a6+TjqdFqL8MZzC6nn7ruUVrKGTTSO3J8LvycpVGTwT/xUnn
JpqwzoOkpoUCSoM0utvb73HiOZKX/5JXNYLAXMoZjrO+p4kyEulwc/YeLqPo7itw1QBr4oyjKdeB
XO7dnd1bcpBcOercPByZ6OFJUHSzpbjknkwoaRo/Il1GNLhv5/w9pCw9u1d/2m7hfUCG6/Azk0OT
BU4rXzEO4atev/BAD/NnpvDP4/2dGGU/vynIe818Z/t1XlB6tM+4BznqE4MXo5pQEITJmmb2vv7s
iy/4zJl8C9aNRQyrQyiQ7U+k0tpB33VqPshrvM4MxVa3i2OXCXjnhmfUIRhZpc2nbmOU19hCfRFs
wuT8Qfo2tUk/y+hluW9NEDflp1eNMLkMpdadOlcVNql77eDz133T0odg3YvvyxEpV5PfiOHMOtQU
XFujDUpskwHNqx6D3u1IWL7tTsTH3z5daXkhYCScLO86T5ZfESZuCBaFmgrb0iV5fhpojGg1CuJf
XGlXt+/6d7MuWZqI0z6nW+3tCuZSk+D1hdLYAg2e5qbexepeCUaRfLnNOG84jWkm/7KL5fFVYotb
JF1Imk4SJjQ4Tp7ovx+RfhKYBhxrH2F79LOXMrIk81trXXiOz1nNG97ZUHczVnwcy+kRTN4byzax
8SFiIy3/62HJbNdSIKKiWfG/SehzmFD4UaEKiKp5p+j8z/2NrWkHKyxLvO/PJyzz5dA1Ke8a3WOA
LSSpQdoP7jhl2zS8HEDkL5F8Ht0girhQMOcclI6vR64e8dzGRPu5SbY8VMyYhoPdX+KjT2eG9/nJ
9rshHUamUqA4kBjR26BHyrlxKjBQwLApXrgP6AFNZwmu5m2813WWPJOXOR9eKIxqIi0l0t7kP+Sm
f1qwK89BBhc5yLt+WWcWry33ngZj48Oq8apYlOrejOhiNJpdMd4ibPEhBgh/AL1AVa0NmqiRCCDU
c5twUu1/DE/O5sAfBxqYofDA3iCzQ38FJVGxD0nRUheCt/F3YLUm5kvBTAvDZkATuRFXVxadIY2M
j6bVYvE0bZ9/AEE0lGFt1wWg0Lq1qb25F1aEkXrJ7ODmUa24ybMVS1T48fpp7cSSc2Bi3Tmqb29J
SmQRsO+sKYoI3DABqiSmlwqBoVyqm5ticlsl4/5SrMA+McWG9rkCQ9tthnhhgMmKH+7kftIUU1k7
mM7rpg3ss8vo4roi8f9Q0E2NXkxCc+nn6k+fqQe+t+5uvmb3J8Th7AsgJsygzi3h2d6TDVG/1zUU
BtNrBPUsBC8J96Jb1KiBUd/rghTemt6YIuX0fj6GO5MKWrN+JF1rlwxYuz/i1ttJ+1oy+OUmZ/MY
HfEnH2S6SQ2pcP9GVgVoopAxG30/jGP/qIFAhhDjeDr4XIICvqrKHile0SEblzmxtKcX3LLBuxk1
Wzqp7uutnroPXU4K0Il0nZIbDM74jHtm8E3x8Led8eU9OLTJYTcNRFTQuzWSzc1U9zKJsui9BBO5
IpVxMXOZm1J5gGV/qw4xagA3H1QNjVz+5Zyla9RfY68PKJuYRXbZLzO0AiWum6Ud0TpVX6V4OwW0
/oNjDDNBtVBUQ1dIgSsLkBDKcmtOjTNTMz5Tdm2e4Gp5CeblS3PeVUKFwO+6VfuqBgEDitZ3CLDY
he1B4/bgBFJGC0VqAbqve2XewCmummnk1JCqD9z5SW2/glczfaA5VQnO/tgXSeLVHwpYFxrvinDp
zRdcfllvgI/VCZoANlRWTjfKZ1pCdADE7pMRSd+JxXH31m+FKnh0lXhZPQTvWItkE6jx7K7hABnK
KAZurp4yhUbMjN3JSvTywezuHEW2dgFc5mzJj+neNo/bBc1WDwe5u+6we8u7QoW1Hp6kYl4ED1dw
uM9EJAMgw3FXqoPdEFsPp6PTeAdocmkqDOCiQxj75BnIC35alJXiOFYycfj22bdxkgz+FpsaQFry
a0r8JBRv9Lf3/ncuUg7hjnE4cWbZS9/p9dyVq4hbFSq9hdgqjpE+JBZnGTDZ1JswPkOFw5E0NoiH
ApjV6QTndZHEtroHoUBJfMI+f7WfFmSHYoPnLjmxkShc4Wa1l3kIxSdXO5viiwQKMewhngkPKlHd
zoAr2YIA/XoOyK6aiLbt24kEJ4NH8lScJWxcmecGAy5927BrUS4CQHmemg2y59RUj9wwCHiEIVpU
0PW4ZTKXZAy/kpG5OAhjgAVx3R5h7ew9j8xq4gj+rWXoUR2gSqj4m6AMEsTTkr7mAE/J1xcNMEbh
wIMBJm7IrI8FpKITYjZDG7PTJNn+1wq3AjHWfP1Z7QnB8/zJr1fIlGMLEKuRIUOt2knxzVoqCHC0
36xJ91aIQhmic7rdiVIDDZmgMqaH0LeEI9M2cf3FTP6ht6AVxH/NAusK+DMuFi/16S2t7NKKBpeY
0UdFkC2nXGkueja3Pc0DkzV9fcbDU+PfOk/vcrvW+7YNbANMDV2DrKnLd4uZd/697KXpBt+iYNMt
tOLnDQURP7jC/CbAkYkWqhmkz3vmh9LCBbFYpL9fW0z2Y6Dro4B+QsOT9aSNgbohMjItlRP1Pzyr
BeOjH6vCwMMN1YqMAlxBo0oeQ90Wsvlw0QPezVHWByn3PIfuRsWflkaYyuHyvtkNdPId80P/pfW1
xgd+HZ/XXyxAp+jVOV9qjf1xC825BEc0S3Ku9gYjWxln8I8ubepPTz8k1TRUaBFpFmL2ctTPFNl2
oCDYQGkLt8YUDLqT9m92bD4zyk23LIz2GuUkPJ+qQkqrqqH+Jxekawri2vG5X/LUCz21ySdj3lo7
YRNu2smpggusHwDM1ux5GJw1SnfGuYUj1678ynZ3N7tbaKwrUzWBnT+Prp0FnhvWq/6uMxhNN9qZ
0Th0UtwX66i73s1yJguCdBR2DDsXuk0Fs7ZxMOpRrcmRWt8M59DVA29XSM6Q86dffGEHqIHBCOaG
6NTRwP+h8q+QYALPyDclDcCU3bstmOC2tVSQYF7KC78iHDCreMEbKiBNSmZejQR2AbTfen0OKwQ3
61uGDTdksxbKUOJn74l9cGEOqGzVYElfx4RziDDo2wVEDMsBq3IYB8JX347jM+i88jqSoN0Gd1KW
vtOCF4x4BNFeR5fGfAOVWCyU6FKPFXm1bcUu7t4Zyz3/gX2RQkXiYJ2wkE2CQwK0ixWw8RQ22AgU
kjDHmLVHOeLVJqczTh5NL/ozEBvRVJOSaQnY6q6KGrCaVZibZi5Q8PNcNyy/aZSFfu7gQaQC/ifj
LEC5gSyGTbMUzjQBEOM0YrvRSEJupI+8X6ON5eOEj3oElVRzZWG+Dz8C2gNcpMSYXiPM9zFnuqTI
q0Vko3h0z2tIqQqn6y+HZWkG0eoF1jjrMT3rw5HSiR3CNPdpBetIOCEok7eOvy6hvKu9JsawCyi3
F3AHde0i6mx/d7V/BZlEehRGxeFPuMXuTEV1e0asYOAB0/z0LiarryVDrRTAEYRr9qjXn3EuExrc
BGEvCVrqXPSnJhzxSNJjLJGB7RQpFv/W0ZNSXMUeWzFfyc7N3GdGRsH+EpkZaREe8TSAWiTAbn31
DpRVWWSgiyEnd9Zfn61TPlb2ZtgBv55/WMQUBoTQAJHYQUL1DZV5sUljyJijCJpknQCO8KA2WpWU
vrImjIC2+XZ14M29rZE0VUChTWCyjRtQIjgeLf81VlEo860opEg3teu1Skwsf6EoJkbLlTyIIYYJ
qmVQYOho6wPGGL4Q2KTg5z19x+w41kU7L9Bdq3n5sXU6c1JRXM4DE7059k6nEpuw2AUvJfMdWCFg
YJjV78oAmplohZ50e2iVdcdyiD7h5r0fX4WtmRhsfMgtINeJGztaknEeCeeThWff7wtPpc0mhPLq
TyqaCDOghyxZKGnrDE3bPEzD7KuK5HBkj4if2UhMi8hYBqGeI1Hx8f2CNBGWTqUDBSPBC+IFfI5W
WoKSD9SYGou1dc79cyHwv0r7o8gGgIBL9KFhrLgMP2Q0xeg1mpZvudiDcdMvxLCVz7+YNOUWySef
UkfAYmA/yIZQ+dHPWn0FhJLHnT5JpaiHe3l5re/hzJwNfIbqROfjFVP7GGW6DYOuwPbSyxJYGJqk
yp7UXM6W4eBUGC3uluYNFSRMQ4ghr/pcKZANai6rs3TxpYLfLfKeyYJhe/vGGfpVONgHF71Ihf0d
Bc5AvnXFQtM6eMcADXA1LItlq3Iaj7l43qdwlU00Mkjy021DKb13Y0xFClQmh6VIgF3NOyfl77to
K2nfeThN3AbHWNbqfBvGN0PjtXLDl6vc4Y2T3eQ1D4YLsCD2gsSeKhZ69fh6Ku+1ey2uyJZHdMAR
H2ezn9AhM/tqXG82r+nDuiMTSeIa27+3RwD1/MTML3pMfCR8vA6ehtBPULbia1qJ2aG7um7Q/ZlR
eZgM8wRk58+AQkdDCZleowLbFrqMdSQTSs77KHCTLjGRRxvmgtpHtVpUUKpOW3K5mb11nqO6DGJc
3FZ6FhCi9UEhaNkACdN8nwOgSe/4E/dlJypxkPapSwnwBcEqv1vbqpG/RL7/WojX6Addpo7ttcs6
ekginqo/gZrBBzZO9JK8HhGAdC0mvq99BdV85+ifu9lB5lIJxgHCHVuHIdMLoMG/TJgygHY6ht7Y
LgCUwnN8DWL4ktEX3flsWXXM7iGLqUvyxt+u1t0yEmxK9o+FkGGblYj827RLzI79JEz4+SCdpy01
UO5cJqr6cN/6IvA7tziLN/RODcf3OrPsi/jFfgRWOST6J1IqGZqSHK11dtbLG4WbXsZvJSDsYFvS
+2W+scwez7tpRH392pYPy8HwQhEL/qhhkdpVE3G5i9rEpjPHmUhiQykfwQfk0CI/0GEVnYMkqBfI
bV/PPEdngfOEKYSXGB9TJsAhPBrDyf8Skwf8QJCcjGtTIpY7eHIOPHMwR0w0/rEgyWNXcm8x6I/b
baFEtcxBwFzansW1EHRL62+3G/Z9i6C2gR7rGKJFxQ990IQwWP8MpdfgrQfMj6XpRIV/KR+BZn5E
ZuqGWoqoTSLr5zkYKhx35V53eNPMl7gWn2qdW/f+/hB7vtiSta/weUB8jQuwWSZ3BceUZkyZJl0W
Z7XGcznaiU2RJAbQ2HyklerKwDTBoNl1jIsZfluBFQ3va6MdPPnLsflWlr5J0JCfShK4ldYIzmcC
dOu/VpZrPt3pqEK/F4gTM4u6sHebuNRceSnfZfgxPyO/a7Mek27tC8KmZV/3/3WYy/qp7wnLTRbi
dgJi8a6p51C+ay1FOwI7oGTqEsj8mfoL5SEP5Z/plOPP//aVljBkgLwscPMSk/YqqC4MSGledm+4
/I6yBq846rMQ6a81XzhRzzZKRjrOeKdsmxK2pB1B3WnhRDDUkyhBmWPfQBTDAOJy5RZ0rHXQ5hk5
NNOKK92UDVBoz3avmfVF08oxqqO9rvDOLIVvwAbjF07u6jTURL8zcDJU3DuObQYk8pBN7lnz5UM7
mNGebbVfqKVdGVII8OjYM4HkGqXytwQN6jcbpCt3OEQ2tCwES8tZ2hD4zUt5DKKx8al9uwCzTsqG
MEV5B5kyE5NYpCOt/SXvs2Ta4hTejhgnmviRl4QszMlUuSy7bLSrlGz79J1Qpaa5L9O9m6/55RP7
QvGX8NtZZBwV7Y8oAlBbLrUf7p6YFsCOfKN/yMaWBj6D/z6z1azlauqZ0eZmfshxG8jaY3SEFHrZ
85zDiNfvqJu4N3kxaps1rl/pWjOMiCQ33eu5w4qoIllbSbbW+UIwhqzaZv8JVvz54IT3ZOQEB9zS
YmYqt+/MXWs0XDm4BjflOsCeijbCMOdlYTjoyjNTxYeG9HLU+fxysPE9h+4bvaRSgWRnA4VeA76d
0S4gtgr8+h+HtxPYL0rwLN3PV7EclCMD5FlG9v2yvfr7ZCBP8j1t/61mgCsek+F5SlDhfqiSfdpt
xwt4gL91m1+gXmvQpSA4tokgboLoCVPjhFS8UiFYCYyZFJoc8aTivlPxTmbYVmLLv+7TBhLO2ueX
nPa+TsO3ZJPfzI8RXy6XgZktPO0tZusMC3Ds6tEjuxOCFurjwg4vDFpI84v/YBXufQP5GjnyrxRl
/nhu9giD1P9/M5wOLwSC1xJ80/wwPqkk67uD/Vn7PbMcme3vHWtpbDkbLadjJajlBc6G1sT2I1GG
IVMe+6AbkWQAh+rhEra3qah3hbYwFDuDOZNfvzzaQpyQm5eI2O+sq/TI7Q2sX11hN4pIK1psK7SZ
NFLKdzKAIHiIKw9CfE9Mufojsl99B2JRMqcp+kKTdzRMV4+Eu4if+1iQjBdxIKvGplfYQi7AapkF
fT7DD89FtVKdRs/soUxJYNay207JqM+ppUqQI0TL6gvqK9EU1VyTUniEfZA9zdrAKZMWEY+girS1
CwApHzZ+cWURJw1uImDuckkB3RZxI1c9fv+LSj7DqWj6CCzWRKz6XL9iw+NjsDISfFU2gZSJrDfE
CfMH/PIM66ZeQAXgR0qb+Z1PcVfTtm2UGkA2O5V8SUZftqi5UG1rfEtcXSZJSdViaFby3WruBH5R
KSuX3IZXj0FH5aHx6XTEZ7/b6t+Rb3kW68zoMjsni4rTeNyDksoskw9F01w3IY5LX4MSfuoiTdMB
SXeCEvy0rW9v9N1SHLz+dE5H2IzpXG1yJBWAKurhALdissV25GURA2y/EzGBQVQuiWVOQfLyAQHh
fej466YtU9Nfaqkl8u4nDOxff21N1BrYKFoyrDy5wZA1rqVSfVwhCg6LCu4xloPrZggkVS0nSttC
gGWblRxi4BTe7HCRyVtsFYeE/WUVsd7bQD5scWX1MI7GRjpXbPr4FkQhB37mpPfK9uWpiScTRHDX
iKQEjgAVf0a0i0FFKNLitJgRgNJSm7CSSazbI1mgw6lrntaLUbf4ACkUGTDR9igWlPTmpxNHG2rY
OtbE9QmAIBHZ7mYGJz2FAsr2BEEp1s3UWcTAtbYN36sjALtrFDBgBSbuLXBC5v5Qtc5MB3CK9cJG
TvFi20q+AppwJINsC4d1PSKWiirgKsn+j1DOeO05kwEcvXpjZK7nHjL/Ga4X+BbErG9U+RrMMq7J
laq11JF10Q2/PtiskCrDIFWtVn6EA7l5mvB8TvZGju6j2BYT6GSHkAmZuBhl9jmqiIxM8x+euy3E
ORkGGTMe+Z+23h0lofOy1bnOhpgDmYmFEWtJv9lUlaX3UOfhPt/GnQTKEzU+gm7JuNEHWhDIlbUJ
6iRcyd/jeYgdUwAi01sMkhXSFXwmhYqFwAc9M5Pr7dmF+Zc0uE/TStMywzbTRgJ3URLqqO64p5Fo
azSvzHu+ahpnYMEma3fLPsNsA3WnRNcP3hlqUHsZ8q3d6p4xRwPiX6TFhz/9QpB/tIxUmyhpdhsu
EIYB2UeH84Qbi7rU/5H98lACflPVJgju8qrBV4za49/JYyO3i7lUrWnz3oE1OYHG0a7sYj3fG1lD
fgY0LSlKmxoY3Uxok0sxTSbYnicaRiRI5kAb22wAapssjsow+HgpFctHe/7RmRgLlbnElrkxrqRx
ObNUNmDrkblNCfWbwR55/j3yF68/HJ4mv7/xzl+HiQigq3gVL/5Mue/SyO+YpL0kwIBhYURzmZD0
WnXpPEMus6FBWiDBz1tG9abhBXzHczpAgoQ48FPCcdAwb8nnho4fEwclG5qYDrVSUqgK5VcncRUZ
ccixYk+/f5jmHjZgMZg8RKe1WJdOZkJfRbFy7cnf4F+CpkCk1+7FMw/xsC90vaMUDNJh1dGLxxPL
yttbt3pyP1eu4+xYtCE9rQqdCr1DKhgDDXxoQ8UM0EcIeVkm41J0zchnZuemFmoBK50hg+Fr3kXn
4tY7xY5Je3aMDVoSGujc/uofGFvXl3IdT0kEMCPt/FdcAAxQ7eW7oFDngAPNXMpawIYwpeBjQKdw
kvN1R9FoPjOjMkrK18HEcOIQDE8q8vcG2il1nO+Z1pCoUt+H1OfzwkrBx3w8w27sBMABY0VHcScO
QCj3+HeHWgfr7dF+feu/T1wZnAFkxJzCUe6MVmauX170oKLT/QLz4MhRMD4c0vor+OfuwfwjO3p2
ejnUu1FIR9GQzIdy/hY7TycOlqWnBPBtJzsWID8GSOwNSUkJM5+96OSWb7la3InRGY+CYumndp8d
6LEe/BXtrCRm0hJiatDawFXXVWljOx0bkYwNEf//xj5AhHi8JgAPQf5hgrMmQSQTKKEaPKKmTbzB
WH7WXZG9npDPQoHuww649qEepRCfMLxsbZjzb2c4CZ/ZkjB7Jsu6LjuPzvp4vHsDt6sflzf8ILXi
K+FTbdieP6kSRmUymfumCysLa/kxSrEXQsUIm6ufqSm219iUt2WtJyiTKlLiytE6gX9zBD7wnuBn
enoz2q/oS+4LsI2wXj6ydPm6Ja9cbkGnByZ+GOQRu3pNN//SWpyfP8lgvIbQpExPT6GxrcrluYsD
V9UVUhnciUbC+zW7dbytV1O/Lq1zy6xpgtzLqM6geNPs2fP9qdbtq5EKmK1TegUFU6dWdcQRoYSv
umJMr/LGKKgevgcnyEZF6o/NtRgFayCuxfA3UzcQW9C2o5VSCJAh+SxEO4Z8VqYIsyQIGUNPxTAM
5uVnarPaOYMWvfCuGE1atuf/RJI6MfJ85FxfTTpwJIr084fJvyadk8rQ9T8RmN/z5McYmq9VpuIf
ILlXeUqUGT+mTtMlh3Z5HfqhKt55dg8bIb8CeBj0kgA1fBzaPW1V5Z9v8LAg5L1rBprGcr+2RqyT
8F8EGctlZVwm0Fyx7Iv2Z1fbTXAWe7bO9K0P67i8sJs6mY6fkLNRl7k3C3grEAUbJ5ZVkj0drkxf
/1fi7IURDe8Y++j6jLSzTZKcDAZ1J8JXGPJDEPs2V2UMU5kduH5NiJiC0k/e1BDLqkD8vk6NKA1C
mlGnfXr3NtMgCcryIAnTha+XeVbwNRyRUXxU9HJokOkiBjoCc9gw49fCBSxAPIkZ37LOlR7uGlYa
Dc6wSkKfuiBISl5zDacgCNoEnShzhSWO8fyjtTRhY6p7Xb7EYpztqrXhbfPwknHHA42zk3KkqTux
tzZEJAn23G98R1/qbAtRxS+UHG0nQS835ODwVzTFCQugeaQerdbEJSP+joQWHgISV8CPfYL0qeBQ
nNKqOM+1fsOulHlkIHoMK5v2k2OyKPBYF+tOBcxAS30Sgd+7Zohp/7li1HIWKhhpd2Ivg4DPeqy/
tESjn6JlucmiBtFkHxDbz3ebbl5g8wmKc1En7VOh5xEhImT3u2cPIuuPutjv7tMSXZDAtKR7d8Rk
wB+2z/A7opSe1YNmUWblq+iQBkiwtgdNLLc8p97xLa6T+5TF93dEd2FDNi0jsxN6kJJlu7MD96C3
NKpm6WRuHTnhrZF52bcu1e7yvz7P8ZjhUZ6IIoWs8mSPf3kkojDR/jD7uzaGuIt3ATKw9FSKywu4
wNwx/gjjizwc/cYZ2kn3MHmG22NSbuUk8jkXFqotq3Y18MTklUQtuNabdP+pO3xod8D2qEaRukvS
NEHRN847y+waTosE9gyPJAXfNkuRivMJyRqYnLo1wPFIv393q4PuCFdzG0AU4on5E/zpD9Vc9WKd
WvqCWLKPuQ/Rloz+95NblwThdE7Jt5nmSXCCbrzQH8eEk2zfNzb2q1w6ktCR8qfQ6b8FdTuyOIyK
NnFrUZCbZ9B/E54FhekWk1QAnp2tyx++JbVFAleNTsIw0uCAWk+oKUMLCYxL1czbsptjE+MuYBUk
p4cnquGvMEofLGxZ4GWogEI9jo8ECJnE+MHUY671HcnssnNJBcL0a41I2QgqZLC41nDkHVJHFBsH
g/kb3ex+rTmdTrj6rK/yijyshiSs4dOTq34VNF5nf1ieelpU1zgYYHYSomxumWPSISrUPJAtrSut
SNmNS2UvNCX+inTCaS/jDF6QuJ4xe98Y+0e0uyOa1qeWwbD9cGBNQSsnr6++KgwxMPfqbcnRU/+O
dIhlv5/XXavEO6U/dbacGWGIYbBuvuV+Nzu9BkUOKBPH8OuMAX90LtxXURUAXSijaDehjhcR2Wm+
XugnnsGWIRDtuK0ouLQ9YQkG61o5RTRh4G1FeFsxv88lbbyTyu8HJEbIt2cjbb9hUl6dzUBXB348
06rXzTHy6ffTtoG8kJ9tg7RjVxru66b90Wx4xsavxCkOyC3elk/A+MmNgLdLKh7mGy+Hs5PzDCxO
cZlqu/vvEmNGADC6uf5F3tMd+Yvvbtdh0/amHabHAA5nFlB3FihACPRoc9vtpdnUVQHpGxLgcN5L
aWPb3NbEa8iGmsa6YGYZ9q2sv6noxLlHMX6/CJjbQHwOHdeIX1e/9S0ArYjSH8RWRI1UUUUiwgea
OmTYCpgOcUUC6+RYYAITsf1X6P6xE5WmnirZCczAFAHKIpBsOfHOuHgchabVeNwNsN1FJtwjbUnO
VrXnIh7MG5Nsr8Qgsn9/sepAkEveZ6uptPflg7uMu+FqcPUo8RlNYqn17DXBEfkcf4CILYJwXQu0
p+KMiylgy/6I/Mq8L8su8EduMnlxov7zN3oSqw6jCWr5DY6MLBrNtKdrLpNw60tPu7+f7NcbgkMH
/k408v1EiwQMs8eeRI/pTA8x9Z0jWTCV3p5u5Ls3hRXQzfyOiZzb1gTCuzuz9HvFnqdc8AUV3E/G
lYkcPnU5LZ42RUxX7GM2gevzl0zFeE7BdGfNNihnARMOsQd6bvokuIG8tne06Fnp97kH/wfqync8
BOwU8ADlanDtF+uKHcTw2220ehw+mFU5K4ULuVAIA6ffaeF3WPJdNTfiNYltnqqHdaNaPCvJeY69
mClneoss70zsFGj3OoFCBAE752dKk5rfk66+ItDaLFHMvRaIO0SVGTAwDx1YMwyy52epfqxH/DY4
siPmXT0Fg6GaxR3YVqux6l2tFfGIKiufAamfSRhTLcn6TKpZTkYhLyEqzI3k3S8DdCEpMksT9m8l
BtmIy5U/bvRJ4xeUnjKPJhNo23aHTz1w61JoqSkvkIwvYDZDwy/dfZZopp4ZSe8U+HmhJliFNrOS
PyPiG/zRMYSynWBc92cGZQhU4GEiEJaHw9O0miFz30jnqNW6sDcIS5O8FntUktMdqjVb3c5AE72f
2lH68qw34omn2oDSO3SfPBccLOt+GlLdPta/qQL9oeBr2OHiLNZMpsPv05919oaXU6Hk5idLY9OZ
/POFG2xx/kQh2wkeWvdjDAiX9motKq3p19pHgPg3MtQlmE9q5kPHO9j+KZe1I1TkczypSb3B9LEP
x59UH7OzO9tS8kzIui0+OJ43+yH6J6wl585mrdnIMvrfbqeSk8KGE9gCsdjRa8unSqu1F/OPcdA0
tnj0JG3hiFaWNlalF/DExhZ2wkHjkLypiwY6hv1KKr04mSnvIWOd8SH/TsBKSk+D1WR8FLBaR5Mc
Kc1PaE/T97n0o5r8hCPin57P3JIBjeNk1p289BFFLTSwpv40F7o4JwGqBArAhvrRxAadZiSz7upq
SjoKNyhWpX3nndBzkgbVVIcqNTueI6Rd4/d5piy0JRVo36hnBJw9rOZQE+6dKCUm6G2EICAL7d8a
PlHmVxZg795EPDOTWdMPsduLEobZd1aXi0sqmswoGIy/7whETVQgzkAgl1Cj3UdcL1/iyRMpHQZf
aAsmd2rpbMsToLI/unReqpfwceM42dhucXD7T3a3VIw6FEwpzfNLEs1fCdNHPVLPWL/IlP2wLyLo
BKkdpUEP0E3UACXcl0KIlb0VBOzZComAGef9au4EtoO/erWhWOnEo0JWv6CIcqmX1fopOISGBwid
hU4A/VSiiZ7tzH5D0vJUI5vwd0Nu5Pzaw7fEbXFE2KD+u6Rlanr1G8RJvqR3F3qYZWOhjCOou+47
jxSfLruP5rdT6/b/svvtu4uy067EJJqjPxDLu+jdTh+zgB+MFFGBxntK/JiW08Azp+rJnnnAENz4
w/WDkk2s754PixwyIl/skbRUN165cSAR6AnjYfQ35Ct6tGf17ClVjfKbBcGkp7r8ZRZgMmHnUnNr
V8FPF2IHpmspd/z+acgNrZbPJhMzyhAieBl0pSJ+B7DaAUERFABXYK1SbBrjduhLB7dQnWTOlycX
5U1DNw1DYT8yFA00Ykq6zhi0B6VFHVm3nM39OAUMBJyWaUDs2Ng0AieAKv2OioYsD/DpyvT0Wjc1
dFBb73YKHxlj2q+ul8rAyLS8/MaUFSFhPQOQwFyaW69Jeq+uYYfTmnQR9DPIbyZ9bUPZNbATfdMj
it8JajfinM9ugCI7jjaZhNEV98GQTUeBv6p0uBqou9RiV/Qh/hStpUl1f7w4ZWBEYss0n/4fOG8C
NABxOLGtfbfQfkz9bhetdyTWzp6sC/WTnVNpT2QGqDrfIR4weGEw3yuLuYdl7cLScsnAr8mj5sYa
afDVs0V3Ny+EtPNXgCBjdgXKwOwjUGOg7PjcYo6BF0AwaAfkjZUUMRDdqWLvFHS8ZcqzWpio8Q7n
zu+56WkzdFWWvWIBEdQUwhB/4HSuTZENAmtlJ/k0eHoHweFJU1oa9fy5KDq8oK1SH3T2TUF7ITRH
DvAklLmhi2zkE5s8zIPfGPQuSe/unmDTRLPtps5CeaDajtVK+ihB7SL/+YpvlUImqWJdW9SPWmg5
evkHirufK5WwnFpogj8P4E7m5fEDT0qoJkSqlqfQU7jzeQg4Wd+P63HCOdmx8ZHuWQwvrPn/W43/
EGJgvlDITs3NGEWTT1PHNJrN7fkgXCPR3lD/+i85WQdO1VTRR58jkKN6TGxOzPQ1i/iEU/5nyFWQ
h1r+6nqTlekF4UJlYwluruYls06iTVHa+zpdZO64f4Beyb2Jz0dzvb66ryw0fFn6cK7eiUH9A008
QdGtqewsSk3fhW0cJeA8ogyYFBMnsvZ+FlccvZi+7sqjZag/gaJtDSPNWmKcCeOV5VFV97fnW5X8
A0UfKEG06symsmonZaVzv6L4o/isYuiENeKwF1d67EEY9prTPs9nZC17RwrqfZFd/OIcwTSk86OV
8pHNjtpnbmHgKL+0c4TL6dr+SOc6EDFF4qObrOB6SLEnqAk5tiBJd2ggbgduYQD81w6KNQRSyGWv
vbmb+mqkR+g95mPDZCjlNLKQwl3WrJAuW4ekx7gJmvM1SY8BuZcN9A+j7531KTehDlTpnxcT+NPS
1zGfl8/HuGOERoJCMdtk5vdQB2LTAz9lQU+ILHWuasZRfAppbSisM6Q6zC1reLAnOeNBHXaqN6K+
IwR04rfVCqqVLpgC1h7X2TG7yfwKVXxwXM2kCu8nu4VEORiuCSzQzprGNvN0Ic5vesD6V/poR4DL
aWFxVGhudd2RnBXtiWgAGTxAa3/tDwvuGxUiIVkUYHHC1EqPOVjZoje25iXHwF7MhS4xERG+r4hV
z2PU6CdsJ20+dsfWMvzhyBMHw/7JpDb+T6wgIGo09zsKv+bmKRuFaj3nYiH+MWVCyFMW1iKiwYpA
/Xt5HtLed7b1A7noym7ZB4wTXplngDn9PyElLx4Zk4hXL1XkefOrM8r8nj1PWN39adESn+Q2gCHx
xq8tUsGuCmmTemUUOTuEK+SwpE2X5qkDNYNybxkfIKIuYSarxWpUn6Anl4SwP4WliLDCEsogh+9I
rzjtsj5LOh0276eBFiiqhmGEZIDLs/STY8sArnmlfZsn7ageaMX/8sV4i0jhKY2m0YVTOrgFDZRL
JpwXw5z+Cl+BW6jBAImH2SZwTV1NdiROTS4jZZuYgSayXvbDPbJ9SfEliAumB37zk7WKfsN1dtyC
lRQWNbLgZHQzMuajNpWA5MLBxOP47Ix6TapeYP7je0+ltHGWiq0RhI94cMaOMN3KQgikn2EY2Tdn
ZcBahTWPDGtD5EMIdYnQkBtV2veBhmz8KeW2g+1sn8iES0OcUBIGMIzOPJA0+RkFAZJ/DBB9uec9
KHQwElGI34Cy8MnLp8Me0UfOzBxPlTaUZYwPP0Osnc2LtEarsHV9W5Lm/k/GMldmYV612Euz7rNd
9NjLKQ/6KsddFy1/o4EF8/LjkoJes7idzRPrvt6JwN+R8xW56WluxdaPJUD8HWYLLXES3ixp8T0z
soc4meVHnPB8nGzHGAfclz49fmR78pgRLhr01G2xuSbxHsPSmoZ3wfjUhM0PwaEUrYmQsI+X0tFv
Uv34OUgd4H7AEcSO8TYqsDPC6RqOAl54lI5RvC9QkGZNLaP9lOh6SnXDpjG3ZoijbOvd9Yd4EQ8X
vflx3ylZvEQxw7iEW/pi6iOvJEdrLkjyA43CaY1YH7dh7Cm4NIrGVbldn2jIYGDxg5NkpIkwKMeJ
XbYV/L46B8lUFRQ2ztHPzfvBVhQISwptCpRAVhhbPALYn6SV4JlscfHLKktpPkIQfld91lhEu7ls
KEPwRik4fmvPcveyv9Pi9imQySSv1sEo7s7gxrlc6PEEy+ylLJ++6zUv2OUDpynYRiwit2bde/i7
4cB5IqPzL8wDutCQdHzQ9UyHUyPwMNLwJciH5AcD+jxIUmbtbLWLXX4hWYEEMff6FYaYswzEFBkH
8V/zo0VuppbJF5XGAw6QRaD8DlnNWATkehOoe98viAeTX/Dj2eJDIIchigoR4xsT7CkGR440Sd6N
kw5IZQ5RAjDvlKB1jJegbFdvT4thACdxQvipsycBd/N/rmEFPCJ7xuWR/N5C3BagiMwSRU4Jyu0H
gC9D9gOoLJlS0mmzGipO+420Ta/X7RHvd2HujXd8OWNlreQ6GtGQA0lTS42fsX9FWlbjY5KHLpfh
XDYV+KEQC0NN1/24LQozBV3kMZFzRqUGbaYmvaCqZuZ7UB11T9eKWO1AiHsGf9O0JFt+YkNpAka4
sAQqS5AmaC4bfIYVuNSz/WmFRaugUZ/X5ctRq6LBjpArbA0rX2rshJCIxZhDN9ZTuvkZcEmvLB8F
8d+8u2xGaz7bwemR0Q4yMFUScgezYjzquSd0iOWiheHC+45MJiP1bS2B1ncC9CZToNVyhDu1QUZh
pLhIWURWfbsiTlJrWk1wOIWgBRErspRI/+NbBI6NMWoctqzfahASAnKviZYeLpI5uTokojjQfFYp
FD+tokJvmahqES8oQvjyQCHz+0vnNvxkEDReSwWUOKLaGOY5fj2EDknUAmPWVq9OLNs4q++8nXqh
O0klt5XcwwFJp5WOvUwA5jaANQurZIlJ8/0W+0NdcgLRa22t1vemdPx+yl058PXhdil8PpHaJoo/
JIlqWcXBb0OhG+eOojdUrmbwa90FsRTU5HnCdvIUSilbccwQ24lMI6wt+Uq/ztiLE8OshsB/iQ8y
j7h7Pud6Ne8FLS2u//ouVZJc1htsedGyVK8AouZ7NMoyv5KFTDoiImWfOvQsGsOWSxQqVVDD5/98
7diGXjVwQl2RKB3HGK3hguQ+OZlg9JBNAc4b4SeC8ddHiEz25JGfxscIjRfQgPVW1dOIOQkZVCmi
TMi7YYfe6OJ7JQcMxSeVVMeMVfpqZRxuxW9fQCX/4EA4cS/qK3rKcMKiROKbZ9+TDnhgN2LU8PcD
LVHLZTLz5jhIcT6vTqArFyZnI8q5S7HKDDXxIs6PakdWptNlUyIkcCO7d8GiGUqsfw6LRLp1IGHw
zzj9j983wPNm2AdCCWU++nzftX+pT3HyW0Z5I7nWce1j/vReo0R/UEtlQDfWHfMY24WCKz58qrK+
/eQUY7YGhCMt0RZDzJTUiCwCFhHhtApL4niO3SNiUGILkFyx6i16I2lUgrIzldvw1VA3rRjZO0R9
FPvCsu3LT15RZQxz9EBCaSfM273oOvagoq1fVMJMBwSdz51sPLcvHdvH8SjowoA2Ntp4AaLRkmX9
4EMXMMpbDJ0BlB+2JYEGZw++opVJmIJR9RQ/VnjKuN/030RRG2Ry17z0ssCzkmG8utUKrww0zldP
df+xxDH6Pm07DNYT7t6cy8lS2ppSeA+T2Ov+W+QWg75+T7lSnmJTEdhI+J2YvJlky9jwM7sRK5tc
BP3NiOP7LVXP3aPpiklK4rVeRhRgfx3cqRr7Jfg5oD7iC5j4P3w3eVLPz2gh/xJ+aNXNRQdaR9nj
y8R+qajQgbncuT0CXa0YQ35KrE+dj1+4me3hm4BJsd47zwPIHOPmRy3N3GOR3HM0QdLzeSa/X0v7
nqSQAuPWooeuOd+Cs3S+1HMxGNhZyzLuCPofxcgyLUhdO6lS3ixNQ/0a+LLGEy7lDBtDBzp9DPTB
ZDC6pRTWbrqtUqHyI/IggE4QhgOoCCttWAsF21hgysCW4WOOIGzyl/wzL/mDPYhOgvnvM/Sx9g5r
aL9ISpUNsiLQ2Y8lexXot9Bohl8Am8toMcnbqUezlfwg18jpt+BwQ5vRQJT0ZDIHD7OVvq0pOeJg
WJoHYZkDfmmAlKHzANHkGchjOhnZ1F4J+oYnUb/PjtFGLxv9f5/bSXqsje5ZeTRYJOWHvzSDlYCR
C3x2Sk1i3AiWO4zSSE3G+6M2tJSCbx+iJafzt+zyrbDDR5zARWX0Ci9OoHRr1edzTao0AuPMzhZ1
QN3GfvAfsAEDK0hPszvEglc+n8A6Si28KZ6LbZ05HqYHNPY+MuHtvnqs+TmQu5Q3cKTnd5uW6Qw8
fuZiGSEze3TObLCDYTzft88/Maa3xCkieVwMpdzac4tH6vjglD3iHDKMH/AwN3yPTNFLjw5MVZJx
Yhpa56E+EmY0AfWSY3zE2CwkUEMqHFiVeENV4fs3dvHfL4aE1giL1NG41bGygrBBVQq8J/wZfKb5
gtfUAFyQT3VZikJ7h1OuicW+0b9hN9w+y7J8yPKnXD8D7Ub+DpY+/ckTlhBW3F2toHvYtwfTphWD
I8zDhH0fpQrE/UoJK65M7Iiov7CjW2xHvJ0j35w67aWn52UDEUjeySoH1h7Ketlz0AaJ+f1y9CgS
DVt9PhMkXHLvkqqPDfSG5N76Ls3uDREUyV65/GEbGLCanfgHxVD2cQWdy4+vz56osHRjWsKdnZxp
tJTjCGXWsfsv5n29dYgHHpdyXmNNVnbFuLjfaLFXXevHrPu/jhK/Fuvun1YR9Hk3gHWlRCmIaR7u
j8P+QFNxO4rwZbokB7LhJgAOEd9PWfoj8Gwx1zRLSfPj9QOwy6shz7lao22MOD9YdNIvKr37fLGR
tMJhAqNt74CI7ActYNh1tmfZq3FeGeAZgPVGBAQtO7VsDjtnCMueGDWxkQVXOjjOx3clTsC3rEop
hawcaTA7YcqS4hnB4HasWilgyxJ5se/BfC86jUMSMBxO9dzBONRQBGV+pzl5K30EqMaadkXZuX/7
n6OO7e/LBrXpGKhvdMZTyv0fM/b6sxZnOzIZSaMpQWtM5ovPFGkbtQ1RtxD+xhVUUp9ZStdO0gBW
wdnmGuBBBs4EqpfpNCAqICLwBdDmiP3YKp2WWjF6lBaNjhlr6xWJ68WtJAJhYQ50hQsN4+qL1I58
lrPjh/UX2+r+Q4nNfnG0W8mxXd8Lm1+Bf2wbP4JLuB60SFzRvM5DECmzO4vaj1spVeO4xrfB+EiG
2O8/Ib43XujX1L0ivaUdagCwQuIE16/vSvhB2jbGjgELJf1vKkuk39v9gqg+Ne+fKpmcOBkehXXH
nX08kUIxz6bJQH5VSh9V1ecNNmvcIzCiiz7KulOgny9z6V5MenTqT8UlVjJGVbJIPbchFnvV1lk5
zogJIF+6K56s/6ReVjb/k1TwlNon/DDimtFvKxFWGjTWCwZqmenJ+qtVADcbKv8bgQC0RDSFdL21
X8KsF+vjfo9MGpO+KvNhaAcIJyX7RBMsMwFr2hnCZ6vjC08wWC/pQCoygewSI48QFj8LTZ1MxUzS
KF1Jdz8elZ+HH+Qybn6PdKD+3Rg4l61yBxDaChvpBuoO8zj3bcTxHDA6U1Tu0/7s0bnSrV7Bc8gC
owPCe2YLm6WCyTCoo2Ff/0XHfA4lrS5lW9vokRKuqhXT/+dVkmggrH+Tb6piO7hu1i4Yfcc28hz8
s6Jt6kfBSjt7G8fENTOXm3WlZNIzf1oaiwkH2O8Q01vAerAolbA9eXuJvWO1FeAezFd3ODsz4KPY
5251xG2fuRuv9beA8mYjG3X3Ig3CMWvNh6Sr24c42c7yYRAZtD1Dq5Da/JIDwLIEQlFDNGlyclsz
dUWeT0LjowGpPX9BFUEaSdiUrzH9iQj3WZiyu7c1FAtuRYYrzbSjGzE0Je0/9OvuqAMHyGVLmYoU
7ukduArolCr6h1Gc7ku7rNF8XoyD1GnCFl5hzQDhRfzFYHbK0Ftnt3ol+xTJaXLibSkBMupnvkib
1hYi28fWeaCT/LSYQXwiyumgYdlO2B4yD/uIettHTpo2v79nr7I2xfhIwjPFp5JanI09euBnVgbZ
PiJvqE4FZ6Nxjflk/Cz4s3L4uzL1NzyKU3YTId+PdtMaZmT0hZM3fCvo1a6RVrodl+Oj+D3mkHA3
ibLkvheoZqCSutvRTGDoFPmgAdouSI2xF1NkHd7Dqd9YGsUu+oc0VMG1I2taO9pHD+aSAZtk5k7+
G6zOYxDJXc9b/RbdvDNWpA+1oP8HMzfl26smy2W0oqMvPpGv8oeAsyHyxHmtRpdrzbpAQTx5zc76
8MYDY7RKbS8q5pkJe0oAIvS5cNEHYtZcEy5Jjw+8f4+HPSuoNcBHxNew21RZmcV94jgwyiurldby
BLWuTyfnl6TQ0oO9pyjcRqKpiaJOX3b7NZhxT5OsOrl6S2PX/aJ+xa2HJDNKZnxFqMZr7Bzs5MnL
LZwlDdsjs+YVpXxAym0At9lTv0K5zr7j/bQrP+/qwjvFfUn4prHk/mCNzwfLXEuWX6wC2OIexMnh
QlvIWEz5Gq4znalaC/zjSXmWzpOdv+LxQT5e4Tj+Tb/g4OqlEXMoRVfh1TaFHNu/7ycluguVUcS5
3r2he8vEFnrBLGWOZRnEaNix1TV85RJirfhRGs61yTu3BccYi+JcQ3rMipZttfLKGc/V2m9ybaCz
H+7kQA4HTw54C04svhifEQqiRu6db1XsddYpdDDViO/mcUJGwMVFFp1Y3VRBS6XXNjDBuEUMp6c7
jD1/mtqFnvsNJFwCSFVIX9n/1vun7xIpyBvIu0yx4ZyNPFOrX/9bVcsRYLrdlqSvXU1FsEWzwE7J
0FCf3lVv5sZWlNYfWA7sFgGZTAxlSCdCCKzGjzwlPOr5Llte1ktQLGWxjOs6WGV84qbIzq88ZL8r
oVy2MU94r73hoTUS4nRpbd6+9lVr9hEMDFMcW0lYOgkFzRHoAW0M8Py5G0nSZnL5VPgVa+8W0H2s
9G0pVAntZKdi+zAm1QmGAJPvFPIra/Gvt0PIBGwKPkmP1YjjxmTG3tTycqMAXFNmR7R/unQTz7QD
mlQs51fptuKBleOn1U07/sVDTo2jD/dtfVHehyv/TcUWK2cpnj6+TrWkZg7bwY+tyIQLca4yXJkl
xje/C8B5jxf+25f7MQ3uwiaFRdn5V9eFqKhFS3/dsUuIOmYWcDcpdVxEHtMP/orHVS6dX1z5RcwT
Skpf32MxlczZexzT8aDD4lchoqXduYiVqfXciMsVuR902Y8c/n52toNbHuZS9epFGq3BPyATPquO
Uk7OtrFVM3o/g3QFQaUhBeeMusFnOXkG3IYBGqdiMIFjPI4cFEo5GwFkuD7AsVnM6FxuIwr2B2ez
crXGYKDAums+kUPMBWByWmSJDaofKWvV/q3JIrQKLz8mzkl5ynEzhjaNhqhISS9WJ9kXDvbDiZZP
FVFrRbLm5FjFrn0PsuaARS8pcldX3mVKEzEAwLacuidoyusfqaBgsA7uNKh8n8LzWKgMpDPS03L9
TZcuWJqaz3y5Nd5lucc1avqqWdDMy7YxbVuDdhiozzMs/je/OWM5F8L1g6tX7uJuKEczBmXsr/Q2
b0w6LL53EMmd2g2nB81vYaHhGjeOruobgUAqL6kTvz+U/imgtZpUfkA5abn/jSEvibp6S2pUm/6K
JT8SxeVUzGL7OlC8UXaPC1LmAQyWQ0AzESLzi4nGGdyEp62ry9NvvGWuVmvwq2hVKcM3MKeEhoHc
eT6XQ/cFjb41DQXxYKNsV6pcKnev//wKccH9ihjFaysJ0QLzIAboUhtI3UoSt320u+X+IPb5CsQz
jIFA662+gJBMnqUH1XnOEq+0vik8StCD/Q6dvmfLny3mcL0LJPxkW0Cus3J2rlximj+GfMUpzKQi
nzeiDsUeLbPK9OYJSKwv/g4y6+3+QEAs16hkXFfWcTiSvFsvA0B2rvMXuZZ8g66UOUAKAsoel5wM
SQFdhii2a2/tm5F+upgVDWeJ3HPTtTPLxzYKWaa1IjK0o0PhLJuwQbE47rqpOPQqtBfxTPCw7fTi
ZfyRqJTmMHmLcuhHwa1TQwHt9nERx4zbXCB+cWsYWrfo/lmGPpFf1US1oZzxLFMzFH/qn8B4r6A0
rhxoHbNSUS2A1cEvbtejliBmOwYnyYUCJtWCYQmMMI2XfwpS2HtkXPraIY758a1hEqjhu34Us0Z2
OvQ7Qf57ubX7/j3O3Nvs4Eu4lAfOp5bh9n86O5EcFoKDOjXlX9GNOOZSE6y5fQVnzLEmsOVKuL5v
HvSSv3VYWE2EBkh54Nw9s8Tke19GCN9tDBVwTjkOjREa8zCGziAFpCzaEyDkJeI2DcJFuwwST/Fb
FRZvigsvl8nP6fC9fhuCnPkyxRq2NXJ+ejIGXLj2f9X7PdocwVV/+9M3z9Ucv3QBZAi6sDys6Fsc
+F2KJKF5TL5f4JXeiM83QF5ku10GZTL13MfiybMIx6i9Pz5jUODkyMWC1QWXdXeYI6ABUNgAfiGg
xc7NWXUfg0Sn5vtj8MuIosFTml6yCcwh2zvfzI/cTJ8VfSkxrlr1rSnoeo0GyqPsQJHMnWWWw/Lb
8CDst7c/27LFHfBFnWMOatk5I4Cy084CCUiMtFLr52kDB4KlZ0wLrGmdW6UzXNUGYd+aVSBdWz9g
F5Ih9IBZ9RLKXNl5d7+f9xxKyUgyFOELP3uDUIRsYlfe+mSAio/uSckFusQNHh54vt6f315IlKaE
7kADTPo3KOXsoTCQBTjkqfBLYZNTaLuxN83gXDk/hH4+zLXKVed1uNKfF2tjZYaRn390xuQwXBDe
KazJdbk9KjWZiYEGUNaxC0xp6xnIDqFjckC5PrPaRPvQEdFtjC+U3cUeV8+0UotdqTLzcND/YyvB
gXbD97uk0s1Rq0CZk3UW0n4nk2wR8ff0bqlHWOgxrVgS/s9LREcnktxcialQqKHEGSXhvhUFdn/T
bSE8iL5rvnZI5DVWbnhIar/ZtB4jjhJgf9wnD05v4aD9eb84+x46ogvvlX3tvIEpmSrH0UT683wF
0aNr3yXMrklXY7Kh8oOi9avp6JPKi2jJzF2eC4jrBizGPsesE+B9d4Wj9TCUq5T7BKufbzjVk4za
LmxYvy0V1cDVRZI8IyqCTouQGHd670X2fFM8gZ69B3UHqPVEAkI4xiiTw5mgeFcZ1Ik4IXk69nLp
Og450vFyUsPYL8Ejyc+OGdcJ840O8vuT2dhhSIHD3wXvHwEMhDvQqTq6yF74b8diuL3FJunAoSpz
caENCkCWFbUWiD9zLMZpihkXMdeAD7lzhRiDV0IRsPuFk6/HJlqRqR0ICQxR7AqQzXP8hDF4z6aM
jJE5mcGaAN1S2oLY3fawJJ17bjIG4xGSYq8abFoBJ/1jf2Y62SJ276siye92VZZsb79ChStg/vah
XK4IR3FKaYvwiPX/sRNUZBSc1l1EZ2ITZvfc0EIYpoE5NBPO7CuPUdYytMzFegEIwKM5df4oyVS4
0gPJCswYwMmI6G++bITeZ8d4DsaZOJEEmLJZCjjhUXlAUm2Rq3/u2DaHgscehDFd7bZt1Q6L6iJb
5D28cPAnBDdXsNM626MQ7Qmr5tIY2BzLifkGt2WSqnOX/MucCwMzQ2tR1B8Cb1Zw3/wjCOylLCH7
WTX45K/aoDQmVgtLPArlTY9K8ke27j2LPo+cxhxACoFPiO42LY4Pa6P/5/DEmZVaD2iY2MVnTsSU
6qBiad+wlYI6tXvJ7tu4Fg9D10sVp4/ugqMA/MPp+UyKsdCGUy0Wn4dv6J3t2/f4ME+OchRfWj3h
G5Hd3f+g+05COhOuzs5MZN9m6hZRTfnSg1TpJU+qYdKYQE0bc2jFGQGXgbZNILDMKX9PHbVezqcj
jpVq7RdR4rJuwbypFGRe7PIvorwflBD83esHAsubHqWSnPdKrZEG8d/OMw83t9GW43Bdw/gFoSMs
9Bqet1D5RrzYl4M+YZABKs2mYviQlt7tFgiDqVX183TZdtwr5SvttLWrqxr91kTO7ffAOLIcWv+J
kF+JVs6NtdTPhzUA06QCL1F5rGPQKDYB5ILhrg59gMGHN3wGrYqhzdjb9zav6X0/AQFwuqlExEMJ
HjPsFneN5piefbXRRa4KqM/94gZWe5SwwD11dnKBnaiIUh+QhLwGdI/leBQlytX6aCs157gKJ/FP
mR8eitanRn8FYDAQWOEhzavsd6YSKRZms56nkJ0Y6Nl95RzwucOW/RX16tfEfiRCW5D8Yeam4uQv
w3GVFSEcE3KW6bBmL9UE8tSrIXlmdn6W1BhAd07McPpYiPt5Qwsv46/lP9/cUEPPk2lBMWe1yeMg
B6/RjdG9IKt9f4emNcrLui241T38Z+GC7d+5CF/z9TM2e1wFL+PSDe9cQbuarGUqQUVCO63lZsMy
rX4CRgGWa3ty8CSqpfOh4WLm0O5Pxy4BgULDJAahz/9YNjbfc+Cx4uAWgkmEG3dxaK7+mYjR83is
0SH80WonECCVCr5yx2/LB5YOr64NS7YH7Hwal4fC1r+hJAYXC4A2QoAE0EEagFUda0KCM8exntgI
DyWvLF2nXqPz5LqOUIdfDNKkHkRA94lxrgyl34cA/VqbX6eVsa9/etr1pNBACX9aJLXoXQKC1VNq
5PUfX2bYbRFUM4F371FADepyXu7cxdvA3iQdsGBxtT7gFh/fiSBvpPHXuCutGlDX+ZzMoT9Tte44
18RulyB8ruPFMV6S0Mf9UfhDkVV6foxsQMseIhl7XxzDbr+GuD6segbFQ93mR10ZhVwTgf4xCzKT
2Jb+J8pVCEyHVpfLdJyiEKllXbsLUZwi6OAOclOmegto0+7/htOpfZLCUHaFihwbv859VNEvRDgL
2mVr+EJZAQBz+Cl49aUEiPg89nIpzCK4nRd7Ao6Hzi0uClpeQyLtkwQzYUMdhWB5bGRf+HcSYSvO
XpBqsPvjCpAiRLDoy+GgzCPiDroochHFQjv7Sv+a7Nq4jFd6JCCHUmw0cDOsSxmBflCgRvwaBef6
r9ZJIIYue48YN8lihFQa9Zl4+F8ZDzI99Qb6nMz8gvX2iY7stgBoHy8t6ZjG47AHBRXGvF7rZSw1
pNEGCRIz4FPjTVhku3hHpnsBsLKQ12ZeHyBSw15W2BjKTdWxZ/3ju+te7koo/zd7zz+2KCxO3mY+
uvRZ5hCj56zReBXFmNZIgCsFDgwL9i2Oa0u5vdM/pDIru9DPIqN57fokSP2rbfBNOVSXt+2wjisG
+CbR+bpolsyqlTZezvKgdNg6rqqYfPiDI7AvKsUO0o6a/AVfY0Lu4/GAcamhP9aWNm6Y0GFmXnZB
6l18xU0/dknDUQe8LVryedDhjAGiCYnm4XXy6UQPsUWKYLZVIM0M1iMWqxiYLXjkV286Lxbqy3xD
5NoDFmDWSYWmhtdgYM8AaEe6KzkYv1qZH2eGEhEWgsZ66JSvwtl+pAfZBnLUji6CW+8vZVn5ehDS
Zpspvkne4oKWzfzUE7k4ngRbOegK8BKycSph5xwwfeVTDsgt6YQWrRnswuuCIELMjmNkEQr8BKAZ
sgeF6TYbCmWwlJWjAfooq9MJig6KcsdLGtwR5NOHtMj99prhdZuvN36eHVkKcsYsgMHjtbDc6HX4
tGUJRVZRld5FGA323O/zapPh5vKglJwRfPF4OQUrhD40ajoqFlFnDGF7ZyjprDcItWyxB6FTNn4U
GVECmuouIM9UjW2kJu1DWqMV4PpwedWOULfZx+eF71aIc6Jbp3Ylpr+EsBLJQvamEjcSYxJlBG+Z
9aJiqcwhu9qknaNfYqCItkKMXOebPVS/HF40UH+qhH4Wn139YMIfQ94sO5DaDUli2WM5lVBX7ZYe
ZnEgcpYIegbFc945NahLMSCibtoMCV39HpHw9ZKb8shFKGyyDlCYrT1SI/Fuo7LVNG01NGvgdWLW
O1yHIL6r3vMA3VWKMK5BK29vF31OjucfdKVyhib0A6+/7NWSYpH8htK1YOFZ2XkNb/WLMTgbwdfe
1u5ODLIU+7PEn3RiRcIK4F23gvWW63BTP/L15/zpLk5B0MvVamiFipA8VSAlcAIdIh0qecyo8Cuu
hFVYNrgii22PEXUjZk2Ft8VqBS77Vua2CyommYRwhrShlXs+yh9+puUBkjgO9HY71bFiYbqVnb5z
7uuJvTv3Ijs+mbaeCypSNheBU70IKAt7uZqsaSeIaoteGniiVo7+07s9b8Ta2Vgi7iaq7eobWBGB
dAp5Qo/4BL8mTHTb5S1fRNT5rtP7sA2WjY/L0XDOIGQwz/hxro13Gddjz8C9zCL1Spwf+4SUG6F2
y2MqKTfVfayxQW9Qo3bJyzFsFQ3LMN+igCyyTJEWaqfzENw7H7V5wIABX+xtvl+iz48IIIMj7pbp
DvcBMSptR9gL3yBtnhJc5Vw4a5YkJh2mNNPLOVVD/aqwpNA5Fq8mHbVVN5/INO6laHPohXPoV67J
s8xEz7w8lS122MJlmPnxAr01rlQmDeMap0Eu12uhIICDNpm8P++pwhdPQ/+GYyVu+2i5nl0IoPXe
1kvlup0Ro5DF40HVsdvPUxPYovNLbCT3l6yNfwwVut7lmCuTpKxaOWlQQve090+E6an5eJ9gtLfI
ibGTf8nhEaw8dOC4BOflnUH4t+JYdClv7HCzZRlHLfekz8Me2mHIe/BAu05f+KyoqsMxNTsYY81s
5i8UmueWeDHMoKNeHgWVhZm4xZNvX/HI0FWMBgSA2ZKgHizzIkJbgfBOdHrVtUx6VEmZYs6Md9iV
VD1O/05oVGFy+DVKLySOnk//LvMNvV5LhxOqoQKX5QVHUofY44QHqE7Yg+GLVXh8BQTUbCKOXjMv
gHcVWGsCX1Kzl4xS52ADlf9ctcMnmXA/Vcnm85Ad/rWD3aBk6AMfg71N8U++NLhNRRJp9R6FEJnf
K0oxJfMwrrTwELoHcckWO9zhxiIZSpN7mGLMMfXSrvIxiKNhINZ7f2h+RJf8AIoAnKTADD3JYjd6
aSRxU3+LSqTPPh42tkalxCm8EWDJ7oPT8oYZjGDp3ciVX5cgeGBPT418pJ8U3qkiWsvL9S+mzSrt
Wqwh2NuCEmMbVbc++esFov4G2s0X+YTLZEmcuWcTrCGTHuIKvAp0z5LRX3mV/g0ooSzbYlTUaHCf
cGFlmZTkjd+ynHCnLg9cNWbr6TaSUk4No1/bFkz+fMCp4eCo60xBZadtC+gYDAHVlkKuDiG0LnaW
wgEyuKHywT0QbJsVk7w/6Wvtlk5aHtLTU273flfPBcE69xe/Dd3QpJSDf08qIY1ehlhxG/vFpTNv
HPtbfXXtM7VstqVcWWqnPWVlFDdwqTC/t3xpQG9EWIU+oBaqtD0Q86xX2gCHPg9OQjvjysh6UwJU
V8KurYwVI4wwP8DvFwdsuwJfYIxpVsiPLargxTM42sHGM8CVQc9nC6rz54Yse38kfV85KcnKBpyG
gQZ+VoS531/TzBDjMbB3SVDdW9mbzmOxPYYbotdp1YdvPs+r6QzEZ2T1GJFlw3juJnLlnn5QGd6B
IGRghJS1RQ70i7gHN+gM9pJM2CR7DOFni+ne+ZiOESHvtOThRbNftLosVLc57yNRR6WTg/GmLDQ7
GhP0BPAgXuJLKMxqfxNZu6RQaJq/oq5BurUStbwSxnoLhLgu+xJdAE1EsEOpBCsVxWdsNnTlnvKh
9erCSMli7EcPSp2pgMWM0UjQkiCeLoGYgeXCuQ6Iy/URONdXVGTTXOAHsPJbqh6ILSZIlQSgTm2i
H5QSgfgowAgjRReBETpkGu+SpjyRwQICmaunXov0BzIpKkQ4ovpmhJ3M9IId5bGzyCi6STyTWGnN
bl4zw5KIG33txp1LIfmr19ljvNpIquhhnodLXS/Tvnd9qWlS7THe/bJyW4J2dY5hI5ABKaNYYZ2j
11/W70oF+YSW8OczR94yoIKVaf5J3y53YYJbB4V1gyB5+DPMAEm7vg3EoP5UbpY2jK9cc9Mg9+i3
+MYft5h4jWHPWtV5zSHwWPp+IS9DzQIeh0di/rqi48Bmr1etjScYrmJQs0KzHIA1qEUY8hntDFW5
pxAw5Cw2znygadB1+1fns/WApNBkM5vxi8fjYvG2/2+QPIz75Q+0qQJGc4mSgnwEEJU3UjJRfPda
Mbn+dIpUrQ+QA+HuzW3eahP2oLOVjUv+eVuAEPQF/BDIa4p1CZZRRAGi2XvG1T16D3dQFp4XVXk9
6XhCsriRC6ntxSbi+vc4JzA6kFpI6hCmi0728zPRzc/EoXl1DN2G0/2nSe9cMzu+ieoljlWUjuEy
ojWxhIUVNCrorJNSwhlvp/QniuKZ3Zjj+N1a7PCImCP3sDfW82qCfhZ7ItW8uXO7skHx+9p/iCzo
vlTH4u3mgwFqAQMP9gp+dFS539uqz2GfEYVlLmgHtsRyGnsla0JX0I4uYErwt96Uo2k61Qc/kY2f
Qq7czX3DpkJOb3OLuon92CJf954vzxo5Zmfp2YMbHqtA/vf1wetMjC5ZQ1GXOXbkenRPXcti/vFM
iqbUvCJgqjK018TEeEbrMEbWzSmIBkbVDVs85xaBvto5iFYVRh2H9fLknsKO/QyZxhTwLZhjhniC
ttKX0oqc8BOczfBCGihffAiwBkSCZx8sYw4Z1pCJAnZOLn9LDsfAvKmNAllUuuAhS5OqFytunjLj
eBglsbAV6O05rHCXRJzoY+aD7wJWz677Y6oJD7oHGbp/ZVzMzPH9GU6K43iOMQNhFKeIHr570xq5
wIkpcUZUaFXUge3l1T0SMK6DUmd254DFWIXX7XTuqyaU0ndY39NV64uorTzmxmrAxOB1yTV+R1Ti
hC4CTV56v74PoW+q1JoLof8zH9E+K4gQygRUlVVDbybOmDvNLyve9kBRfNZlZD+IcbnQMzjmTkbd
V0pFmURPHfmQvJtNZhHJfKk7oatWVeJ1056VpEda9fd75EPVbNBYhNHPnyFbLTtFjjnynZ0Omcpj
ZufVldxiZeO1NXYJuEqVRY5qNypc/z0OZqpL5u78NIOK9Pu1fH+2dR5QrRvG4NVGWDkCRk+MdF4O
63qTi5Rak6DF3tYwA1efIzzWG81JDmeyyfjGtsqtLWfsfkm0jqTxMrkXEZynxWKVhc0xE8o3mMs+
CFtKcqRxQNmf2Hu8rzJv85GcErxab/ceT8N4dbVjkFkVrYhCACGFElTUEIMiERSmgWuNT8CHx/Tv
vwspRQF1Pd9+5zXrge2dDEdJdCoWbm31+rbCAvDIxlSG16xPaLWjOrtzGJTVWaTSTgnm2AyA36Ba
MFDqrJVw8x5k1XbBi5W1pcOXLTz0oEPXZpWhRqNodrwi76/6RjjRrzeW0fHVld/YKbVgY1ZgI/PN
446x6E3ES19PJv0X+WewkpyEIq6zfLwZ4AZ4d7r0RiIx/PgFUbhWVFCexy52WSZFrBBrCxg5W97+
p67J8Tk5sLgyMSoae434GXZxkhgjQ2w7LBi1mJjGLSJEXTjTXBNhouR0L42Tz8ldZo69lBsfshG5
G+Cnm98qlDgTupXtahaPoZTkyVA8UOJdLfcX+Xl7YjkxDs/WnbkvdZf/NIdVtycdcszztcnYprUN
BkhWgQPySWmiDojxQ2Mnc5IvX4kLAi4YDBk/eYgA2rqd1yC6jKjz16+P4dCTo4/XyzzB7kV9KdSS
lWmBj+aXxIF2ipCeKNUZ93KDZDilehkdHBBgd66tie9Hm63l2ppbOr7EVGDpBLqY5Fu/C31DMhpF
XgRJFnf19Uk0w26/6rkn4VPQdmauoOd4GipqVjuX4GCkANGT3RE/Gbp7aID9VYBsPtn3aNA9iBem
kr+EbDLoXVz11IuxLyttIDj7Fq4H3D84mkzhLzc82Q4AVpuAt4qYliguGp3sWAs2pFmFDvBXUHNz
godvoCjJ+3sOFPjWODprQpu7RRMh19TzmmXsIaYUlwT/rjVxwfBaJe+n+cOjmXO+HzPK2YXOcoSI
ev3IoyNfc9SDZ8Lq6pO3re2tyqVuJ7D6raH44bFKp02osLBCexbuZ93ytAKongQc05JsU7+BYkQe
XzptR5JXVTzErbmFvQJ0iG6HvRTrcIFqBYYMGFV69RK+yjJM6uiiH/QLd+0717Xj8dFrNUnIr6SV
/w/98hVYknA3rTUtEW4SyYd2lXonhhqvSlr4HzO/kKYcW6jdMq2gLT6keaeyYb4heDRcUh4bzVCb
5oTBxiJA6FTqBo22ac8JqJvd29hRm0XZIgUWSsMUwGUbHiqUXmPpad7qGlRapbEVlD2n9M2u47eH
dHJ6oJA2h5FMjYkIqBucPXlRV9FC5lSDoBOshYDx/BAyQQ36qD41LxEgnAKcRzmsBptdJo0F0LfF
t0zqzasmZtFtHQ439F0v/o6atWPW4KZcasEV3yym2aLC4Qx+L21darib0xl/T5ODQcBcC4LVpibS
BwWbzAvbm0n/ggxAZyWt2MzofQZ+gfqBDy9HxogctwNjEPtONAFjBv41O6NyDZqoIbynSEgqTne1
Negqi0h7Jg2Yxx2lr3OuCFGAtlVoXSry4O3f/3TIzwsVhQYqPTMNwjrJa6AT4+tikcUzwCdkIi18
QvHNyfYje5fcfwQxTBCHDaWz1Xj5opAvSmUWZW/70rp0BFpklu+2QmJ1ilj8pG35uoM+7gUCjB13
VFuleL3ClI7qPfKC45hM59dyMtDMi1Yop0qRbFBt3fezATh12umi8/cNtUdCoNiGcAIYZhwTMOFB
c1U5fmRgc1VCsn8d9R6Wce4g6ekkIxfGeVUOOBGYX9hwoM9LWx7JwVXJh1MW2do4xczHRDDEuyWo
NcswZs+LvKd1QWcwSiS/wRe8NRzPV4vm1eh4ilb2CeAJa+rmHcQCCUW7wYZ18a4s8Ge7KXluaHnd
im4gMrqVqUlxC+7/z6jUSHXWR/PLhexvxUy2li/Lklvi8sR17arkUSngXMvrQoXoTENqiEOmBYwE
0QZ5OYpz1Fj2HgncAdAfC8TnC3VIPnEqYf3XsZ4//N6EIE1WaNMVyR/uMCjPmm22EL4odxTkSq45
TZbFyd7EU1dr5YQHsfIDfhd4C4y7Rq6DlMtShoHB5DdJvVT9ZUsMRXKFeX+Yy6TTu4KdJYC+Wdzt
ZsBbhIh41ha4L6dAdENrAf5GoZWFFhm0quqMAXdp04II20yEX2KXV9E94QFDwL5IR/7vIzIG8nrg
1GfltabIXW/LGcdqlc/2fYM8XOYLi/g6uKcJDIPcvdb6LBzvF7SFrZ+I/dWmHnsnNvoX6DxepXVG
6khYyyxLztzbqx6Bu4KmBat/IQ6+DgpEmXp94CGPgO8aQL8xJtFC3+VEAbtEus2gAf0ezGrk2DOP
++ZWzLkneUfSK51ZungbsgjCcwlL0z9G9HABK0jjyiLTAIAPAhm0dZPrG6rtJHzocH6fDu/TrVyS
4PF4ny5AwnHerVdckviMm8+uts6jUvoRnXgHKwjRXgOYChnGKhhksuobo6i4RZ0EUO8qzii1DIE8
3q5BH2WW2I4WoCWZ+h8E1Bt5wcCfqdVVs9TnnZQthQA70UlJYi0JxNJ1/M7Cqlywpyk3OZ6hATTj
jWnROjl27AQG7mMdNHyQb/9VHVEJ9X+YsuYxXu0C7GG0UDzpdPjqZ0MF3CChz3FK/5/R8y/KZIsd
oxFHktWFWuwgL2ucmoBQ9pj5WfmCwO8lBSs/yFhKtuFKy77V7Oed/IDNEzlIB55pteh+R3yZfEO/
BJXEpHWv9Kffmgcchfoe3HmxWyXIo+o+G1HQYGSIJ1dtN+79HwKX5Ss9NgK0z2R9l24tzW1Pay3g
TWU/j36CxfDcs+DOrbBZaJ+3MKCH8YTfC0EZ5/947vKbPnmg+onD0zxpZ7xDeRsyOoSIdlvcHa9d
nr7rvKCslE80OL+cdSrs6sxKG2riXWipoIvM0gfv5nU4HABCdQIaqWdC0wxaQ59L63XTCIQ4E0AL
fC1mIUCAOyNJ7d0B96HJdgdyjWnEjrE9UD3FgeIEnZjKLVW8SS1cUoIBgTkdpjqkTNGG0ODbKAMm
sbc9+hIVVKb6EYlONpB79/FWjKEqyG3X7D7V014Pl5Hl8FZyB+bEJFlWmHJCQO9mpxPSqpE44v/7
WlSPNzFDcVsVbN3wRShsncnDvmhgAnFWh+fzPjfkXxr5jlTDy+VohgVfBKCECmELJEyPBVw+icTi
qQSI6epQVXxq2kdxkuMbvDzyln7ycew0Jyw7iAfI2yV6YjXftGpUm08wx5i0PAOwglazPz795MUg
DRXiyU/Qtt0E55J299cGyroQHG1xAiR6Xxw/5q1JJKJ2hbLyPG9MJ+1Yg8v58YDzo00G9CeZR0T/
hHIPYvZgi+djTRu5AC0TbVSjFSQC9UYmQi7Jpkc/pYkRnSJYsfXV1+xWTWuro06Xxq0gXGNg4fGS
4dK8qDI5YHG2G17hPb/+8ghgLEiUfm+0WH2fP+55Ap9+HVl++G4LNuvJoJyw6WzNKO/uNSmoIScy
Km5J4r7rHUF0lnOvd+M6HtLI/B//ViSpW2uLUQ9nfy14h2iRADiwcHuArZag+OGVu70bfb6W/oqT
7JEasfhP+bvuWw0RoqKKcCsSIovkPs+ZSeAlaTRGYJ6mYzyxbcoqt4rwhfZjvBypDPbeS60j1J3W
bua0oKIsyss5C8QcCiyrUXe//P7xyuPS9YVPbIKytbAasN7eoxYcDs4zZUoD6A4plLCfjYbLst02
CLWU0I6RxKZ2E+IAmpTFKwyetGLZ1wbZwvdJsGOh8lhxdFX8K/nn60D36wwzuL78RaUe9QU2QSdZ
ehB7e5taa2vFNn1CtRSi7C4mjKXEPm1b0T0tpJraCJsWabm+PBLb/1iBtPKn6JnsSWVCnozOj7VU
kBPTIHSluYlwKMBBSTP4kx8WJEzZP2ooHua4Q4JS+hH1Dvm31rrjo03IstJAQ464xL7Y0umY3DHU
SPaMOVw/j+zb2HpiksQ+XVQpcKcL7L4ZreGkLYmoAe8DwhlHAbS44UgnoIRfYT3+YY4ugg6VjP9I
HgaoZxMFDTYjkqUTtiwrJ8K0JFDXO3igPNeKKe5fj9R0FF+lUv0rSO6o31qdi6vJ9f1NuxGGMrQt
BOngM/cLvNoxmHjj7s4pQgZbkuR8gL9tkGaeNG5iX7wPSjNDjOUMUkBJLr2pynMP+8vlRpyVYe3F
vadWL5uP/Y4gdeJ3EgA5/GdJMo2BGyVhd9j5zTAaYAYa+JASEMCgmTPhPQ/yHcwkNuXAgzh8ooYj
v7LVNmMoAJMdKSruuLhmgPf/08tPmvVubKQ83C5hZ/BqwUzsEpy7mzmHpPiKTHwfJ11k5DvGpDBq
zfHZ92Q4Cjf7tubWrn56NBXolroOTxgtKeVwzWQ37UEnb+9cvFiOlY7bqhGF3bVkxI1PmLXCzcJy
GhcP/B9jtqBA4TGk0peIfVKl+0d9wLgd/Tn5eyDYL6lNb3Wnuog+9q5Kk46BHBMLAMPyLK+k/Mct
le2051t66U/U0eVirIEkrad3Y3s3Wa2zJMqS+wrSUUeeIHQe232FLl3rxKfx8n33Vmt7GTI2ph3z
ZUxF8t/nSAGznPahJIUs7fMA8hMevAGPeL4IXe01HVZdq7KURzR/1cNgfKg0vkoBsgCg5Sfflxby
C/qkxgfcXHkQGutNGC/OrbICtfLdCsjUeMUgzO7eUUNZutY+yu3Mh9yRyEShtzoPjbWFx782VlKR
cYB0DQAHrsXUlz4ChCWyxpjOVkNXqJlWUw0iM7tYmyKcsu9ae93jX0hcXRf8ZKrhOYhTrA9LfIjz
vaaAPnQur6FTL/o37IvSMN9XHfKwLO0Ths2fEds0tX/vr7jf7eP/m2CKd/fN+AhV+1BOnZgRYIRX
mq9zbbU0+trq2W6OFwilUX6LGSImmkJs3Ygan6NQz/S2ELl0cvu1DVl5ZlbbXBqwPIwBb/n6SW4+
x28Q2wi72hbn/UOHu4fHjdpxPgMIom5an+QZGNG1B530nakdwWoVwHz35Q9S4rvUHOOmGRSvi2bm
karjQqT7CD2Udyq8M2AT6Yf4gMZusTDyo8BYnnmHuZQnbcefYOc62Xel+510lpkC9opY6nY6Ro65
QfK/xsNMvodnmAy/zoNy9r6ge2HHZoXD+SVBV0mcSJbUK7YxZDklSby8uz7DoEjGob+Ud+aQT/mF
SCaUHNxRUbFPJzhiDEt8TGjFhwDnEcs3sGZpHGhWosHRsKu1GuGcZTR2eXYbF6GlSByAXLHiLQFQ
NyugOCwmpGdoCbgUTs6bXL9Gzeg4fGbog43xD671qfej3ozdCHMbj12D+Y6funHFBJVW7Gp10fVG
j5+6qWV1WOQ6kbxgjZHBiC+piPPIf8qCs92KmBjeq++yfyEi6yZLU3riRvOAPK0zCiRRa7z7SN/F
YYimKGjwgGxtQYisRukTV+BHOOiNO/lnCYn9f+D+Ohzhm9MsCoMvxaXY2OFvMzOOuOKj6liMmsmg
1UIyffKaJqcRkMfH6/N5PeVAglT+BGIBNWNL9wUcw4uX2/CcrtnQM2rz+p1vbLrNNjw0UtBTIY8d
8crrAZxNfCkAG2UejGB5MdbseS9sEPa/0E1VwX93vMUAWOPI9AaQGoPvp4NTVs5IAdfPJM70JEnO
WfFwwF7q9AUBUw2bYj6GyAhKfOSOQMTtmm5EsJurTgev4D/DTF1nOJvuA7yDtT7vnjvDxosDJW4M
SOX516j7j1SmAJnOZudY6ftrNu6lcrzoNjTEIbPmjMs0vECVumo1L0sP6YduyHCTAKefUN3iQRbT
L9UljQazYllSqkOJio4L3ccED+79ly9bFiS2YLAwNTdeIRgrmjIVjNCejAiS1yRKDkhGcnmOtFLw
mRyQsCiqlc26gNFqRN9hq7gnjmvIBIT4hSNZpaMN/kA8oHDpo1juWFM/25QW007fPxFlz61WR93P
7cR0acFwexDY6y+WDz1Ql7tXTFWaWPYMpRUXirJNfac99kIMO2LZlszKTSSmXtF68MBP/5hUkQC7
Yt4xNaD0p//7TwiJl3JtDHylbhJJy0tuic6L67BFUnGV+iAp9nq2IskkHbGQHiiO8bmckQFQqrtV
H+l7Bx1rr8EPcopItkOTXXBeOcAebMygqjgRh1oCvq3HVjGlrhBRGPpvx/onBgfSYytw41vuhKIJ
UhA00QVhKitgjMq0RHzXys/aoyofGdftYGGAQNgfWya8T4s2oMfLpc6JAgiyDo6gcO/V5nQDtghN
/lWnvH8NkKUfwiWRlil9xP8ncn7iytL80gGuyUrQsQ9718hNO/MHkN/raNyPgJBmcmAvDq/kPujl
pOvpE1qKADEjE9PK2MrFx9A4BD4FvdHjHoucGI2nQ52MYSdiV14dqWSbJ/ToW3ed99b0gF/5FS1X
EvIwUStSk4PGYnTIUAoNYpF1dWVw/RXg2mdMpxudd4TAJAo/08eVE1rzwNKb/nLqMozSb2wle168
LUgMKi63AgompfHOI7KrCY+LAg/c1nBxr2XcxK5EwG24YS4WbDZWtvIo5C2hp68ojlnl//daagZX
4vgC4qZedCFDZ6gETXl3pwZ7GL0SasEBmkczPd8W1nL+r/CccYLuG8PLUdzynAxUpSckcNM1l2TL
oPeBUMm4FZwuU5vbw+hp13X1CVvqxe2Bpevvv/6HDAysYXj6Y0nfK7b2gmFbXQ5YIM+UrjL8rqgg
CB1mD4TiuhcBPo0k0fvIuKBrMrVn7O6D5WJXO0O7yA3oYkFVm3h3QUhad0u4j+1EkVIrN3M/Y16/
7+uqKcHeh7PYrZe/Ss7rJLrg4ZAg8rljCikBpupCeAHJLetIjJG+ay6DdymHxTYXii74CByPlImw
SNYp6xiVUc6eUZ06oGdzeyVIFI7FNsLdXgt/77KtcJuJp6aZzqeQifaDpmmBOgpUZvz+xrSp6yTL
DYPcjfP6xMKsYtQn6tvjQsiLp4KMeG3TxQyF39yYY4uf5Nsd68N08VmSpuayw+qbzOWb+rCzedRh
rig/zSRkvEdDWUJA/ZqFrLoJHl1jerpcqJ8WZVj1OE7+CRCEDNKe13m/JCC3jr5eEgrRWm2IXqmz
PbWy9WBDXXU0s9oX/TYE+7Lo+BC26AQDa9mooIVW+rvexpwlGV8oCGe5IwrZf65BzRe5HgWzNcCD
Fm+/axTVbqW0SNvElG24dyEPNH+nTmQWvaj7er2Sj8549xsMphr5aoJchDCAg339zp4x8KAN8tpY
Lf5SfEqUv5VQqAsp4YS474NUGBdL7wINKjoCb9mdiEdm05vpSyggexQ7DxYH4oRzvqWO1Nsp2OwT
I/DJdSNsTUmbuHQICkFOw+r0TbbkPgK7ZHVbE5UASExxjnporQbSGQyumqcVzJmlb/bKTGePkugy
UgTW3dc4q7LhX3QAzsKsmseYETV1SxBteA2ULgm5sKlN+bBe96Ut/5F2Ar6O7/32YnlI+XjmpjED
Ew9AFhTZXRPU6NShV+xUZ/eGkghW2xvEmb0JnFmSz7kublxxVhlEzeCcZCb+AxU3CA/UmxMQOAnY
SuddvNCHvMqqgfp/oyRNe/UQdoYHI7dEwrNeogu0ce8CZ4cgOEompjug/3ViJn8/MSII+YD4Rdbg
t2r8bfPvMd22mbH/IWTRYEArX74SF33SC5Kio9095fxCJ74uJEWWNcFBPoRdo2GZcI/MFglTLi7P
CMq6q15B9nKVsHfm3QIv9sD6DGrz7GpoA//iHp418aZONPTIo/kQfHbQlzh3TupO8hE4dHNdIriy
TLxTmtC/f4f7dU+x2HNPrzWdO9diEIM8KNwu9pypd1ta3C2I1gxA1TlhgNf8WQfkbj7Nk94Gx3Zr
pEMtph1/fRm0Z7SJkNaVYc7efltp7OIIvVHyO8BzLyTu0AHl1cxhAPUE7nM/BdyP+vUerXhlJkda
jVbu7/QElC4IITaqfMTfXO3EhzGr1Ac9x8Pg7ZeO4uHwn48HwXQkSc/onrZqvpdVHyfa5PzlpkFt
vLUig7OoYzm9F92SU8aD/5q6MN2P7AayQjnl+y/lnypMDVptv8gYNqBV+qE3NtvwtGC2wuNFbQqS
cqFghwgESr/fODMvjBxagdPzzf8jHMDv3E8DnpSLU2STIe1L/TBosCBOXiKCukNamcIdgv4nfyqm
AzG9eTaTN5dYki7kS3tD9y2ZC2Xi5RUr9Axlriajyl4KDHQqk6krqZtU48XifOZMhQMGQHkxbOvb
SiZJocFsWkRVRvuweHheokqt261PlwYP3W+VyaMDALGcm+REdKwfbdADDTVEj8up5cOY/AyFvkaR
EZCKw3flhPG8UAefqSNCnWOYVi+dYSeMCe2IqUcxSb64iO8F8PCcaZuzJWQeEo//owuLkT1BKjdW
lAZ3MSB/EPnOZreUeLHhk3V3See3VbSozfpPFFHX6eQBBsXHeZC+87pWoDgcd3UdTV8n/zX0P0Z3
gT3uuiUFQw6ozZy3/u3JC6e9j6/khP7asMxn9ZVG7N/xaBn0LWmJ9XD2TCjfEM6Yidl4jbdtcSGR
qOhsYlmnLqUr6ozC4Y3HVX5zXRD4pPyZ7PR7u0emtAjEEv4HRDjLvk4nWaEwF2wpxddKPH4xkQvk
Ju5QnMnRi/2hRz/BOUEsnXqh6Xmv3a1BDQkWxW4mIOXfoNnBZ10OrEz/sQjet5QBgLrwzKdGy4nm
y076kRnIjZwsaoQueqp4x0f6QJqmw4wU7LBjoYn0Zwqdg2CFEfp06dG/VA8tEu3rmJ/uDAMHV45V
1OXo/ZyJJCfiFba0/evu9TyDtNllv0R2aKGCeOiJhVkwHzaqrNxLttumK7IEP1PZn28YSgvvHGqA
o80G9zTndxlmW/vtzNo/EofA70pXH6XpxkxTVUg3dsl4W9kQ+Tlc8fL+rWOE68wVRZNBhEoxpB/U
3Ubs+N9bn5D/4JpZyrBO5SlERakYqjb+MKezkrdv7U9rOLCxXlzxiyB8YdpQYrHhfLnEqUNN6Bmy
HUOD2y4ajutRgs+HCNggS+lOxb4ZJL/i9Jl5x+jOwKTNrQlYowX1g6aWoTmr0f11wDVqUTJtq6s3
XOfSGkCVCCODBftt8ipJfDfpXSxtTzVyAaNPxd8IP+V2zN4PuBJKS6HHWKgVJB7Nj1WKfdfgnbQz
bc+ipmN0/81w4+YSsoP23lq2rYh08M4yx3p1WcbXSPc3XrbgwdcKa7hNcDHntI9lynW2Od9nSRaj
ROxaJzr1GxYp47IWjX/KeNqz/aZvAWvw9O2HUIspkEA3+IHYVpEDyyDqFahO96JCUEybgKoB/VE1
sEu/50zJOYogYIU5NdvrfwQ0uf2I7DU68STXvOsuF8gy1vx2MlBwXmOBbC+Je2A5iyX9zdIABDvF
u0JEnFCAJ5sXQCq0xh9J+zFqN/Dp9SfV2CtROHeZ/K4NDlKRbS/nFH7td/0DNnXNFIYX7UaFiAH8
kNrPok3JcbIahhP3yakIb4JQnxuZZZG8CgU48XF+mfR5oNkmGs27YeiH4TGXSKedJm3qPAlQl9a4
ijHP0zYJKC5VopL2L0vmR648MWm9RWjUwnKpqNtWhq5SJdTdJFjOJQQ2xifI82c2+4m+lzNMp381
vlY3rpNZ5P+R21yxdRl0TCbmn4eYW93QAcOqjk6L6FK+5Q+yacX5+HF0ZwA/csAOX7QUbFgi/bdJ
t7oFdtEpj+6lnNY+BGVoDuskY4bRrnvmTOtmBjl/um1cz2G7XbG/CWbM8JQULBX1Qlvwy9B4fixe
cuLI37ILMFmNULRcKm6RLQA2D30+YZ2t7YbDReLeU7t2rRP7ypsOi0AxU6+1D9XHAA4svlPSMKt0
UHGxWhezRpXD9F1c3kvenOCZNmUH8Bs0/JPofkzFqJ/bi6UKkXSDlqLmc2sCFmjX5JkD9t8GFPRb
oDjJznn8X3LQFoQV9Zuk+YxsSN8joaXgMWR6gPf78TkK8YC7xBvhJ+RnLhOj2Jx+Sdcq5+ufFBcc
HpDALC93U87ePlGF2JCaBmssG8yesgdIh1tVXPdXQhO/5raHrkGYbnN905zXllQxO91EMfdM3nR8
1lh5h4IRuqfYLPRqNlxHVrEm4+XPCzRwY8ZF4PGm3CMC4DicIXjTQVMLJskhwqRPUmGzZEkhoiD1
SR1XIKXDH03DlqOlGSAapqsRm5Bq3osdupUj6hRi/S82ZpuUfYi6SvHJKPe5K1ibLuX1mM8Ac5do
aEoburnCz43r5D4psCC562bqWr0A/joMZXcKfgAv7+4UyKvHz4AfmWx0MqzxzmEI0dn0xF/zol1/
BQBPnQVi2pTz65n0ivxq+FGjzurdCejJii1MPbWtE/YlPbFiFUzw8zAG/uTROQrjHV5DX0WbzlMC
3TeyZVig3WqApzHyDh5csMNCOlcuhy6volN4ENvy1TWpqyVd88iUUv5ybOJ6SIr+JSDtiUOzaAxU
cGwLlgwOI9GdEzbcMD8E7rur4qL0BIi3fhsY2HcNVmNt9rhnAU+xR2crGOaq5KJKlKSYBOyP1tP1
NUEKg3GWSaOf1o6vcehvWuEN31xocpTRboic559qf+qyRGpgauKiVm51mwi5lu0jyDAocKT6X+RI
nxepfQQ5L5k+x61l5PVtuPTfgHJsRjp8SMyTSi6QM0SjE8isp/OgvBB0dTb62LoDGxlWi4ow94j3
42fVPSdPNbtje6jBMS3csS+fK+aJpE3Fw1otuIN9o8PEddQDvy+RYOHCqOtf81QipV8Ev3aEOdYN
fvVmUFLHx3TwyGmD5o2P2TnoT/XsHvXw1wJBvaR/rbB0ERxr1B6c34ePFC/merimQO60rSvSQ/+Y
+OTSNWBHq/w9JcUj3wbkaRHDp6HUuyjjB49UU9Nqa15AUa7scGNPXkjQhcsAuHViDr/kAyAPFNxJ
YFtXMa3jzzWsqLpQ4VKiB/8BT9cIOUKCxyEOt+OwGYhflOfQciSSA1bIGs+KY2b0urxf5UcSGIBw
5JLvb0VyMpjJQ7mhyfor9oUc11MktWksa7R+FQgeoSM6lEaDjbOWFnFVJXcHUT665vhnMq4hi3mm
GoVSvljeNWoGopgXdyITQKM5wiMtE1X21u9lpVcDMjTurF9WCIuicLjWI15O+DXPpcAZaEIdwMoE
YjyMsPhk2v9w88BXLFyaPyuwxu0XHUOnBiwecDb2/csKJzosMSUAw5ANdmYQPez1j7xslscxYSdt
Dxcmdht2KI2Qxn07LkyNxVAsWc/Q/ODWF84bkLRv6Rksl/4xx3n6jtcGNFnkJ8IWDmq4rl9i6RpL
9z7UhDoqJRGY/A5qOCckP4o2ksefCwtrTlHED1+d1WdV0YEqZpGfvu2e6NYOBFNbVaOISRbObx52
ICrOcLY+p+zE0Xny/j+gobT7GdbV1qqBRm0nLF4h+jS2e0Fq6tK/qZ2vZdnq3uHPjrFJLBOFMM8M
or14WDZMjBT3IsOB2v/cU+Qyulk2B1Cco+rzrIyCjhWgssfNrrFfpWfr6k0GEGt46y6nwYf5RtK5
SVDnhm2Fu6D+xmF3KAB4AQuRXOVWl+79T167SYRYpqBxFxJ0zaOk/gnU40OWzDZbIoUhYBdnamt3
ER7lFV7ipktAwot7Lz300dy1UJbvjoUeGJuwx1bY9vREHM9jYSatNzea5R0YVKdola47Y4lXxMBF
26RbJhUlQaaM/btF098X/HIDHOZauVIgl14XYxCeNUS5g2X1bU6c3tumd0JDVYSGazzxNKA51VbR
BXQsx/+K5bp1cEEaQK1BpuIpOGOxI6C0d2Wf9J+yKJkk6zLwZW1BOZyXFzL7S0u2giDBrBzSU3JO
sxBiacKW6iRtDndjDd+06hgM7FMrHrLr8FdQWwDcI1uAWpxGebDC2vAC4LA81pv1FyLWROWzcXbI
NQyq20savpUfWV4TTGV1J3U+U3+nx+73MXKBf2l2tFO8dDAodcYailFqUX6EInMqsErZKWtAMRJW
qyqDsKBkj5g1ycvQTKAVNcy0kiDrlH+BNlgrm5Gb5MutC5nj7Fql9s8l+n89jDFssrRoewBFeNRL
8NNzommyLp53KO14xr0AfmltX7gRk5lcDV0O9q12BApxHIaAr2kJdYPWjO7GYoRak+rEZAMhpIuT
VQjBIPoyzolP5GLMXFo+ArFFB9XL9xKwiZ4DNBxy9G5+IBY32HYPewU+m+rgvZWcQP4wM2+oJ4JN
JaqWrarCLWfMpXoT4UYbh+EncPmEcKHMcbCnwQdmHmzmhzLeIfKEbp3RBs0ELKXQWHHKU+n9/MEX
AZTyw4HFqLp9nbJ7NOeQharSIaYT3nelIgCiQP800JYTFgdUNoEInWXJBzgO7PgoaTni8a3N4gRk
dOkblE/p0KMHXAhbkbALnNlYvhT/o6BG7ihZAMkzGI02GxSIwGx1aEY1qmgy7UsHuIacDfLMeIpm
qkNcprFvVJXMRMfK0N6ODAWblslURT9RrJTPLnGcFeygeei8IHTZptFFDbMH7wl4782RqIEok/j8
mWeQlH+bIfqid8xnRhD8v7wVVbOVRnWNOU4hvb3AiKZ2ZPdjeEMvas0aVD7WKcXACuOFrIqpa57M
ywqaXM90y23EdSpTTpgga60wXFvjAdVd9sijQ56urDGtJ9rt5rrek6e3pO/yfJscvvg5J7vvCHEG
aYbddjUKbhsV3O3BoC5reF5I6uOOpC2TcYQBwQL1GsgayTrkV9/gRf9wa8SOt1MnfvR4oFOSDyOQ
st+oglpp9F7x1Hd3ZC8eh71W35tLBhUCJj9fB1CErlHyfqMKVkPB1KpmF4cKKW4Fr1HPjEDpgeHF
ve7ObIvGBxzRrRNls8YSQlMDUT17oNQnC3QqIj+eWXQbGb2pwHlf895IqxMPIcVyLOGaBfDXBiVT
mKHf6AQW18Cox46fjhcdO934Pv9ou6DOUvVCyemHeAFE7gCiExTDtVrjzK4EOY3ko2RzyxYhE+jo
Xfzpo3dPeAGeR8Cml5yiawWpQJJTykg67/F42s099ytOIbeAV7eWVPJ+lEXp2fM2q3SqlImulju4
5zrvKMBq4iQPgp5LoEOfjYoiuKrqNqeyIv7LytDAeZk0WXqLZMt6CrSWMN18TdGCIYjxalQNAS5Z
PiIkDAg1+RJtOjENN9np389UmbW5DwUJJ4IxwYOBNO8/EHVYRYNPUNUEmrrinJBxK53ytU53DrH0
tP6agbgDbusWhOdGdv2DxW5xpRR7xNgQmOFHTTFenO5jbU7ET7mhtyjeeZvMwt07aGirXJaIudwN
RzqJdZVAAz5R52dx+wnM7scyX433ju+7CBCm7r9/HE4wIXQA824amY1s6SHSTcgs3eHKFKzPzXGS
a5KO8JJydEXAF7Zm6StRq/spsnn9cMkE/hQ4TPwBpD/1YKgZee9yirCqqKZpTxnZPZf3p/2dtAGX
FNsYnHG3iXb8K0MLObbIjx/V/JsBrKttlcGh/TreOenkGLTuuXVpaRdUEx+Yyn/XnG6uB4SNoW8H
looMrOQdzKJ16AVp6Dr0yiKRgkN3gAMFcpgcqLqz5TrI+7rdD0lEOgARCmWs+n6fy2KHZdKYIC7Z
CI9fffY/DmtlHaD38+HyKkoxlj9XqGuWt6HBKm0lb3vcJ/y4kONYJdWTSS5hJcx7RBWPbihBo/cR
rM1lwa1gG0r0r8Uth75FyCsWLc+Qa6/U22r9pEiORgTzgWpoZ08ZyxGLsL8YS4U7hCPRckm/G9dX
kPG6gbMj1QjgY586IMNhWdTqTVadpgsVkZJdfOp9bdlyrNBcAEBrTzhXEGhDm21Muip8J7sKRv1M
NUQhIUQ5vE9ZKQjc/RYtw0Q+raJ5s57aU2vx5RxeV/JlXT/arIeeEqrfZl3XhtWHCGZLKYXEdmpB
xjEZ4fimfoWLurokVylHbyPlDhznBB2y+y2CQ97OUnMmF9ie9FDuz/4AbqQ+1wD7I+Ls20cWSNv8
l5doitkYrpV3qGalnh/T1UYclSfmf7jHCKcSZYaLOna7cURBqdByac7iWwc88dqqSoT12p46G6Ow
Jtkf6/d9/AH5m+fg2ROnPgjguj6RszVCe/my47c5y+w14QFFphShNGWkDwv/bfylfJyGUyxbGDf9
qCXtg+F5rLJ6HdU/dp2WaGp7A062FdWnRNeGlkuz0Hj8kx9JG6DNyhDCZ6RqnHNWBN8fMSDdl21b
/R+6BZPEprl80dD750k+khEvLgIA6iYTkgKfaJAZM+AW5IGIJvVqAtLqdxxBBoqrncOn3IHK6WLC
5mqwBX0uOgtwjHwUM8We1nugEvuRie0+X/3/URarkOksjZQ1H/VLDcdaWdLb+L1ntfUvGM9p0lTt
NeDmX2hDaW6jHOyGnjkxdhlxmuqShBXDB5NwSV3CHZhzufEp54iJbmnqdNddaOFCY2KCyEqGyvPc
ze040cerolpSb+2M+PwgS+hWq+Hns8TSYQcBKSyjfVcRlJvegSl6/AIX4u0vCBoEXccC1n0qnIN2
pD8/K5L9S6Gav6cZi5ymXJ4v5fPUPxFpDUFSJ6O22oN1nSylQvsyKYd/R1HtG9CLcRs7IokpNSx3
K9Z+lOG72Dp/PdSbbtHFcNhrlGN9PuC5+0Kbtf4RP2EibC4yDeZC8fipmh7IXgsxgGp4qd93iwEh
AfDPQ8G4mygN+95NAvu2yH+ub8zwkuCwuwMBDuJzB4QLP9DEQTzjhaPUPIyFY1a6dH7/1gawYUgI
Nu5AUxoU2A7TUlq3CER+K68eW9fX4H/Im71bCA/N/NeHiY+4KYur75z0Mk4vOWhu3AJ1NLsU6fjl
xEensulg1jhkNmf1TE5n06n5tJaj/gNfde3AuOCACSk8c/nJ6DhUPAXvTkj/ZufSygac0iA3XvWe
e8/tnfau9pP0oHeg/pl80vxLmq4in294BKpDuwrluobZFX10L7YMw1jp9iQiNUNXKrtGx2ehQy6P
gaTWQMBFYXfnttIaJB43kIJ4yI0c2cAAbZ11RCR9Bu+WT7o/7PriLIT/n/VOzVXJ3j6JO8pPQ2II
odGvbEJRxadVPCJH/i8l/CXukV70OW5sVY2SgX4r4OQ0ermpTBr6Yh+SojQ1S0ugWBLL/qNW8Xxw
Ex0mdFydPnYnKyrSQcCLQVRzGt452YuPAyNMaL/3mbyEpCEc4FJiCsZpqNa2YZ4/Xa9usV/jxoEw
HstiXP95IQp5LGNgiLCn9WCdHaO2kXtiWBEeuxJeAtl3J4wmJUo27shHZ+kwRzLsQGbwQA5V8lSB
GEMcxvtw/Ip8qux/dXSNgoEFT2OJQzfT8fx9d59kqZb3v0RttWn1c3Tya7rylaHAqPGUJtiXbyVv
KXJwxEnfs+HysBpLTKFFXiSUEkcsodku/dMu+dwRc33YoHWOtenrKdVpyyXrGvK62ezKxO1Yrrrw
NjNXhSRPpvOUgt/hW0irBnhdWdOoug7drMCclMUPsfie7Zov/6mCn+48KhcTlb9hPyGfiiP7ox6W
n7n7d6/nUZO+ruDIrD335W8KM9IbKZ3zwnyRVGVoGI5qij20n5lZqxmsl2wAUOhDCBJ8B9g2pYb9
vX1yyXzxSnwVF//A5vmDGl5xxqpCq0ozyZnWOm6IrRuilzobd/bhlbbIcMQkp3D4GYcmZolcoewi
J+8UicLJJr4uJsHYoDwneuouOxRItvu0ozHzHJ2qpzp6akkGMnEEF79MyESanHDNtJNauN/d68sb
uMhU2nzNRC0Zv1OjmKJQTlKN3mafhwunboCRRj5UEeUuajdeZQcrVAylMczTj0Mb88pbm0/1A8W1
c5jjcLbtW8klHCZjUA+QdNpLBoFk0cSsyQNvT2EAaYY6dEgf5GZKVOjR4SYqSXbO32ZdFc1JGCy/
H45YEeR+U8Z5paYXtyGXHrRy1XiVi9N5mZa44tn9TUqvXl62BitxXsEubrwoz+/XtJ4ijgzsuL7X
sOarv73e26NCzzypwjhrNkrwiWXsOpajQkt1mbopa4gQnUTBsZ5isSqoPrUha5nZfAn0zo2ChIwY
r9w/idY4UCnFjNu+qQCGDYwdv8ZB1RFQJ5mE0IqJ2RhNgmO4QUJar84rsonaN7WQ3DPRHVlZ3GUB
O6rmO33qNBqO3qAVKvr4yTFTuSzT4SBSJHhEmpH9qTIhkspdheXOHml1G9jXotCcilGOycGfYnW2
L+ScrhAD0aQY16BWOOzjTFdEdsJ8MlbXEDq+qsABX2y/OYhn/fiWrEcd0bkdOlv5d68t7BKsEBRv
EBpbfq03bEItkoyrbJaDQ9yq0Dy6rKhwgAqaIqKrf+vXpvuAGetujiYwDP+UnVaF5vpatFgki1fV
ETTpMTE9bQ+VA8NYcKeaG/z/34V51nDa6WIYzCK2J+BuumA2hhFaZmqKQCGPgiuPBnVUHJcdKd2r
dGHcosK2zHTkLTUWlJ5QBC8/zcStJ/1R1zYI2xeOWnIWi9CHFgrtQX/e1/tg16MWYv9JhXNINYix
XK4+OyWppyFe95xGh1zLfrJw//mkjfC4RP2GWQ2PRerUhWzJR2LW35pFRiKnGrkdzB2JxPQHApDJ
ToGI6L+mdqpPboZYDBAGuo6+XvQzM4ZdTa+XjD2r2MPZ7w3UfYc26z/GCxMIt/8qzJhoboUk3/1i
WTMzin6I8ATk4YyDyChZo6Ck1nABlhNoVwbi5txdw4ToZAvPPMRT6qG6FX5ngR+6nKDLO3j7umO2
zro2yXRlBJazAge3TA1rUqtgDZyhSF9BiU1ahnyMPQ6VfI7J8gZ4UXokN0Ri5zkieU9TpefjmGhA
AkvdU+xX06oTzHxWPyoDpssVaXYNtDjjjZ/aH903jWle/cpKCSbrdYFrAGnO+LRgiG4QJnlzgjk+
3o6OmXMfISku8U2nHDV5SKZXwaLQ2gAZg11GHwc9+PJQVtZMRMCK3ynbOBqjCOuAL+SH93aoyauD
oUroE6GQqmRe7I5C7fughfigJ+LYEw1KKLedBhYzs0ed0QTspYsqgFcuXLZ5HWR/g5GYiOTWEmWg
IogbK6yIMzoZtdT4BWp+ZpMuwwiW0njvQhf0VXVprNCUVYnDZx+l/eXRlqeYcsIjsDDsy4fa4kJT
+F9wWvXG63FWMZ7NX0VIRQj9H6iGZTWyVaHkRMsMuE3ZfxIt4wC1DUlqxwPuyahQG4qStw1eV3n1
podILR/SjOSyiy3UK2sFhbTfQnThcMZFlnraW0ShN8RHEFX+jfdsdBspLBlk9LeEZnP+fDeuGG32
c565NjNr+9v8Yhxcjy/88MZMyF4V7vnaJ/f5y4WWdwSXyJ1W/xdsG6zEguC5bakJeKruI1y48sY4
OqN6R56GnT5R6gaBiWh8vj243jttrF5Qir094zZ5VYLGSFrxCBV7cxyCqBmWrK2G1+jD5WXVFhWp
BR9fYvg6zLumXjVZcQRztbiAepqE675zjy0uTeW/KcFeDoSAA02Pj3mYVVfWaGEdlBNXCFg5aGAx
6uMJBya08s8AeUPVonaWFJgGiEEW1N/yGmn5lS/QEO7tHSNoEpIMNg1iUxxv026mpa+0oFVXwRTZ
u4d2JSx7tmP91sFA4Z1F22pFTFGEke6x7hLkTh2KH9ClIIGA2k5a4xcr+tH0zGk0TuLpSmBh09eS
0cbQS5Qo4NGfRG/JUZq6I7cw1xtM5/jxUSfdb8FK/K2oE2Zbl+BqYT5FQZVHihGDk0icNuxmWoe9
gUu5KOluQEwbgh13YdbuZKALa09ZoQuhYpSlGMFvmlBMLmv0yuiK960pG4D6v2oqHhNdz3IjOOuy
aan0wHwvMg8MDFa9vD8ImmYrY4+VHHfvT6rtzmzIC6A71vqQmQuOCKcmdfCgK21FY0ZKN1ZOPINh
jmhn3fnj2MI4QMKLz4Dsm84wxQcgGLRR3TL2jJHxPmkRF5U5D4I1+oPvATcTAJTCf4UK/JAQNTq4
ue7xSijn/+zvzJOZASOevxxnCJxBo8LOHSq1GR5DPcMKwSE+teqbIjFB2eMpYdyrWHaZ7P1cxxYA
JlbzL+4BWVIZwlI0lY5Sd/q+8MdLL2XCfMK5KRNKchA/Z18UcDanya9mkTxp765SzgMTQAp0XUlB
cbDerBw5FZW4zj7HFowP9R0eH+V33odcSxBV7BwoQllDRsexf3PuBD0ejEccgX99V5cKMbDqOlYp
bD/utssHkaLRF/xdqYHfKB80P/78As0XR0jlg+q3giZBGdy4dqHE6KlZfaFljA6Ah5hMi3dM6s8H
Yj1BuLbqxKKHD608fi5ANCMslg9Vs3sAHNISUOetl8c6uKAW/SLFnXQW3PiJPTm+dXpL9Pj+s5m2
QB8ugypLsW5kbIq+ua1XK/c8tRkSDrDfkjsM9oC7jBQa9VGH+HiTPwTZ8Z2ltAV7NaMHVPV9FiDI
z4MaXKag0tigLGy4zJI3KZi3I/e4ENHfMuh+NLJazLd06z8ZZLyEHftaP2ZQk/U9+i3C40GK1Uyo
m36mLRMRJa5uWI+FE3sRaPhAwmD250eT8nPdvvTqjtmIfvXpVVxH9OvTvYlQskPnAB1ppYSVpVpH
CGg0ocmdWgZr9LhGY0tLiA596MB1RVt7onsC3fumtpFaXSrSrxRF0NOLX28gxMaptdM3pJRaTzOd
ugKKZOe1uCyr0iHdtIlu7nbn2thNrY+i87jMTUo2T6UDMzPKXeYbsWbscQ5aRjUIMDcEEl1emvj5
eR0AG0BRyNo/KOu6sy8CEoE9ZgjOEhTP1pOKc/xFzJsn0irXiuSDTMhLBY1dZ9O/uetKH23IbgDI
B/KaIJPpQFCWq2r6kDtO6F+3qURcoGCK7jpm1Mq5p7Mu7gR5FqqdA+2obxmx5P8AuiMm1MdXvdWQ
w6NTDuF7iJJl67MQyP1/iKNKxEPg3TmLEHxGxn0sSAXljCYpbpDYycCiOXjpT5/zj110r1bLfKD6
uTDqD+sm0Hantqo10lMNcLVipBB09hTyb+Q71IK8CD6tyd+//9/XatXwgWhjcu6T/GRxCMLpRPnN
5WWvNDz6nZ9yKd8VJv3AyJwYKqPPR8yVnFK6rNSEKVgY5OSulXCDBn5gMElR7sfKfRiTjfXobGr4
djXShm9NL4Kb7AXqDWe7htrERB7pGgggg6K4HF1CCaNRxqsxVwUXWwUkHPM7OLkS4IT78UXH/Gm5
VFgebV2lzQUFq3cmOR6FVR2Q95GQVvk2ks6uGpXyPF3OovYrnOZxZ6ARzQglpnrnZEo6wVCBLzRb
6LrNxxd09ZkzmdtoBwfZMCKIQ/7/NDdwUMKDyP0/Xq0W+xWmFQE0+fWeCAjPd6g/OQ1LXIrneumn
pCBl9/Yta++DgqRclLsEvVibmfqdA14JFy6FcjqagqgYzgDDzU4mc1qhQ7RPEYnL7x/4+3dAxKnz
FECUj8pgM4yYJnx5pk289nYdSQwnafhJpDQ3bd+ucFUqo43m6bxRjv3O57dKBtJSP8lqjxCH0GAc
+/1zm4FJH7sUPyBm4gaW9sHQJLTcIrqQgKhyG2Iq5dE5sqkkMmCUG25gTkb3V+xOLnRq1XmYsOYh
RiKQh/SoENBwRaxafcQt+z8sjjyaUmZMhG6ZuEDTHvoIa5+yoDp/LcEa+QGv458NbLXtd5jdHRB3
EPq3Xiyo1b+7lA1jD4NHBU0u47f4EnF+AHrUEFnxf6+JW+YUXFxUFe9A5OV2bXfqs6pdTPKbm69c
ba9z2zYyiEhXuIrIP9bjtJxCf5nWzSYsUER78RZY2lTTbIhyt6mDoEGpV6FldSoEfQBuOFbeUfQ1
Kn9j7vaZRSdNanNzWq0PVe4bPsKtvQ4WH+MwpWoMePJXOncLtgHn/Qf0+M4h5FaswsIdWeeAkbun
Gt8DFN+h63qWYdCMphVwmzP6A5dM0cjpFBdjmwhxn5n0ChrpyUbaAM+reEP2VLrSLWXMmAU5aZwM
zAeks31vNoBHo1mSGAzNwYiUZc56D9DwPtql0k7ewgAnFPr0lZ5D4cSFqKPDZMveknFOtg7v1chv
GPlz+oeUYPAYbQGU0XTMru2Djw92Z0R5HdMtkrIFflmZh/UMz/LzJbOlw8Zxc0BunqEQcwLCO7MW
e/Hw2HC/bZU5DVgCldnb/enoa07Ppvi89iIg80HMIogkDcHb6Ye0tQ9EG7b5qwwS83Qk1SdB7eyQ
R4nX7iqI1DYvhlfw4d9zXXRpQdhr1AauCQG1QN9QHaqOJqnzcY5sPMckhAkNuMuPaUPcDs01pF+m
uaBuJPuZHhwjcz2EQCei2vJbnAnotdZpJS0P/r9KiU9zG3W5l0tJ+KW4fsl07/0jRoaNWLqNpEUr
yB2vuzki/HNwsNlIHDkH/zaPxrqw7jhLDWbboD9C0xQ1nfszNkl2P6raWhLCysJ1WVwAI98w9RYK
OhQGWI9d5A9TZNpZEOYeypecktHz7WmmVgrtIrgZ8Jx25qQATPf/d/asFOoQ6imY5DFH622CPAGI
FMnBkzpqyhoiQpRalPkVbN6t6MCZS1/pqRP6CWvqxmOvNiiWnbSSsTRZ9BKHP+bW3wOo5sNBZTtk
aEml3xuNZfpBRbL+RlNun2T2enbRNHm9rwtDyNMu82F7lGm7jgXidLA1dS8tzmCzCRJjtGTsqYoh
9OMiBREicxwVW/yeqo3OD/38A+GKfSyTQWReKoYCGCwCxNDAkYCitstsMB3DPuPAx7AWsYXgZTWc
AZvUStXhHn/hCl5vM0ROFmMq52C/uEDbXr+2l90hbvNuy+Sa+Ow0MGIrFfpwRvjy3+TmCYkBp1c6
G33vumq269hfNZr3OL/s1lqsFcQUnVKfzg+5nVXkCfg3Dc+eeKjgmMfFTXMSU8XWGYRRZOOU0naO
LVonlCrSQBtaL1FsKSvfQ0+8zPJWJO7YgGi22jWEC3MVj0OHwyliNy0o29Dcpaozy4EnuXDJTERK
YCDkJhAAtOCHUIKVrP3Eza7NmG/o1yWY+lXMulBREoXjhDK1SYXboMv0RLjqUNtCoEeINvYzCe8/
AbrnLuIeP0FngmBVsXPcewlDL3TWimQ6qO/0PaclbJzg0IzcjV4qogU1VaJXKaFSR2SqQ5qlEet9
vxUHtNWzkVlzMlvOQLl+1aoGq3Nw06I0q0WgMng6vCxyLZinuubSx7lZmUpNogdE4WcYBIzUX7Ot
29wcXKZ0UXhkIXzhL/YkN1BeyBe75R8z6T//NQ/OpJ4T+87g3O3lrSag1gBYxM084b9W6eMQhxGI
qVAHZFoMJE8iiKvllAPU8ZfVMNrcKu2UnY/gT+5VkhvKMh9G+wpsduZM8uXFaYr0kU9DYGz2oMTe
9m/DBxK412agKyEloUjs6fgzegpAot9EJ7oylv/QDA/IFO8MURnJ4tSLdtJivmWxIyWvvb1XKoEV
+O7AVKTqSQvYQLK1FSOORbZCKGoOdrjqZ262wDKokIdKcTMrmw42DpUAeU55xOEj4NsJ6JzgbupM
3CKyAiV+T3eM40oEXuVTRj7ZxN1wH4GgMqmYwVSeVipZxuN3gAfoQMMLSsByGErd1U9RjjrZ0q8v
IilJRUkO7hLQ5N500QqFZmpCKiSacqTf+6rKtORLT5TvqgWCUD9Pc7nuFvz4+idGV5YMAsPF5LG0
Gpz0LC9iYhJirC18rTkWh3KJfz2i3ECI7e3NQ5d8HrznOihwxcl4s8ieD84z8tWazK9S+A3ioL4q
z1vSLYLKfVylE4i/mV+S7gSmIqXJi7YErr0qdjlzVk1aqysPnzHHRRIS5KnjZJEejsQRA20TcETF
NA2AhFRvvJRzgPXt2qF8M+IMPK3K/c8g1o2DZb4re9ivL56iv8pUdS6Szwd6Io5DCPIG3tWII/hT
Iz+dwvHOyI5tznTaXg/cwUmBNUJNHyKWkfjp7KgU+5u+eTphbA3SRaZblSxQyk4zvGHFKVFS4OFP
6feyTMydVqxD4tNLvHx9USfE3DZHkL2uHLgplO1mUuBNGg945NFIzcX0AfTOZauWGkf6H3PKEFyq
MP+9OQJYYXCCy1gU27gTbUbYrid923H87/KoE6Cbg7+hMWg86YBIOSJtejhpAY4rGf4Pmt+aRo22
KVzw6D00UaeAIJyHXnigEfUq7qeMy98TbfCPCmNB1f7Jd1R3yXA22tjrE1LZCbR2QaLs7Gi337mP
aWqs+oMCYbqsoaKaPxyKijVqtIh6R7gXLD4iFdFvNky2iQJixo4Px0JTyYjoJF9Ct5bwPu3t64JA
EVIC1PtXDISSWToHEYMSykGWPMr1f7oz2Pfhcho4fgZu9AXK+3YIfeEx5LYcx8q77zNZUexwnI83
h1yOCkbNIBMUqaWzyqgoZd6FuEqp7hOv0wldpP9hO6pEF1h1OaZDAoGZ2eltXcF2aGwd/QPhciYE
1wQJYzLGSZaLNba8ddo3utBqvsqsbjFdvAF0XPN7bNHkV4MtIPNeUmY4V490HXJTFqFkcRV5JwxG
4gWOjceH8D9O5i5uzvi1TgYnZ7U5r0PFsmC/+Gm8u/6GdMT57aQQnbep76G6YMMnpaW+qnyD+C2E
EDHwAt/8r9xefemtdVO/OjGMK0jqm9YoLG6WFAdmG+wIg2Zu7aaynjuSrbay6IQZeK+++Jwm4Azu
1bZxBxQE0imKGaPDnATKjrAS2OGjFZmX4MkEriZyD4wUAfVLsZsUJZcEchsWoHJJO7WPHo/97ssR
in3Ev+xRUWBYc4k5mAYgaMSDzNXgfxyTpdHk+dQqfTPHb7plvL7z1Tos7XGQHQhIA0QkxWW3GnhA
m7J3qj3vgZPAOFz90Wzx8Kj6M/VkHi2BNeSbVa0dIRUVlI3kpfM2UAx35O/cArLQ9wDVgv/XoBFO
4KVU4mVRulnxbrY0zJ2WqEdYzwGE20JBVINBnU5P5Q+lqPw6JzII+3dGsFPKilUna+v1vAjTxJqQ
JBnn4+21l/US46C8Wev7V0Qa+/H88vdmQ7BFzdI7zhSVDf5hjI78KbcpPq7QbUDbmXhlkY/PfwPG
tAKsSXqZFn1NTmGnHeRGFWkdavKo+aOlbU0cbmEmE0q3CNGSZjsF1spaETBBEsJZ7K9oObErODNR
zoDeYzDQZjs9EScpanOBDYA7fUpeJHcKB/LBFJPPcdo/mXThYYKb9kXhxaw8yFx7rD68sg/BPjXI
NJxmZ8lO01sTKnP8zCjFmjhW579z6WbR4I8RRHVbwngJ0Dz+HKbtHkk3fzTFxM+X1ySw95zXAgaD
qIzer5FKU5wA+QRxLhfaOqHgH0x7oNqBzQ9APEiEJUQjDNkSXLftHYmooIUJXlXKvHm12VG4+fJu
YaBQZwc6s4TX9niB6C/OnLFP8D78FJCHH+C1FmfHfMMPepDxC+LtZ5L0yETm2ORBMQ+TgU7ziZrR
hB6A1R7hJwIFX897S4ZOy8S6QOux7r2/2ja/mKHAAH1WFHLVUgrgWhgLD8vrITqXDg8SBNlrWRTx
2gMRELL61xpw4Ll9qisTxsvbK1IQNfD3r9h87CSlYruljnFFuXsuDq6uVrfJjxhAjJKHNJkNAmzB
9oxfR0BS7uRM4C+YKxHPqGArjU0fN6FM/3VFuVhWr6Kj/nNFoXhSdQvXaM052bqeUuINrHeiBKYq
wrxC5TfI9ZW60X5nqBGRQBggXt9qIgf4dfP6iXqwQZMCNexI6TBnVBOIr39OCBXfyS3tCimC1Tuq
8uCUsvC2JmC7vaFvTvIZeq0OQwDS3z3AFocN/Qi1fuD7rbiuhwHflcJxrxH2aS2hedrIN/OFegkR
58GgzyYtSxGJDbAuXNgfym9kVjapQPdichVkfSyCM5A5uIbXyljezzVy7n7vN6/xp3IqkspLcxi5
t0chyJ5v+vBK865f/MjEb6iT5NlZMmuJep9CyrFTfhaFoRdzWznuL56SdqzYpzG0YPLcaHQQHWUT
Lmkx9Vr4PD7i67PhUfwjRaca1g4mMOV87902Z4MPNAP4w6SEIoQyDsUD5WEuUPkji185/95tdCL9
/LpWsVhUaOFe+XvGOtlw17aN1QN7XWo8o87YwC/GFFVWlpHMfmtSKvJtvnU/DrrUdCrmzWn1pRSj
0Knt/dZlAYGXvEak83wwrOFtlwQpnemkn5K8oXXWj9S0W6jiWRaHaaIM4xItf8Zp8p6SbfMSJEmP
A3zMzByqB+EfTm3Ajs165A1cP4N3CMJDHYRJIyUQ3UvWTupaCOxdVoEiclzcqJ2yh7gSJe5+eA5O
nxPZXmRKJXNo6vN/m8ay64gS08Hlsp1RSxxZRYsdikU6zIxtkZai0cudeDYSybt05dgN88IZwIft
9d2ZR3kn/Or4suOa4tBBdn2XKmlPmWPJa9UrUE0+yS0iafoq0hgNmflUE1mC+oNeS2F88oemVW/+
Heh6QMBHy/2bZskWTUi5J/yLLsKLapwJuPOvh03lNmTdU+BVl11LsP4Z5lbO7TDi6mTmfN0c2B7G
H06ceciSATVd6eivJcISuyO+M5D1ao2fCOWafa5M59UEWwsaWDNmM7tbo+u42F86oVUTCpUcbdPZ
58a9cI2jtsDDtgatzR032VFj1NkgRERwO5dJoHPZE63TSuextPZ5+SUhRbMaVQc4vYznr9fxwhRQ
FSW44h8Hc7ufr1BUQPwCfOQ9OLvA26dQtZPYvnVdrH0O51ya/alQ4AzTvj95I12IKDxXv4gs9IK9
pm7wfiAYC2GnofE0lPOFys9rRBhAodClIYxw7GXZ9fqhooGus9O45UVHRoNNueOvtsoVlihp4tFl
XuTFZVEuiIzCLBOL+Z03FrZvh/m44dVDCwAit9fwcTB+Vy6eIOf11ezo2FBpUiwVHTe8x+Rx73BD
upQiNQlPewwUe4HHcC+B5e+EUMKaJaTgQFGaQ2p0U8f+zVeS+ANVhURmHWf5asnZm27HP21RDU68
PISAJiieCJr9YV07qY2TJS77hBKkqO5oq9a9bG254crKlBdVDrC8eSVNwa+D4bQ7carQH3D9HYWT
S8ZovB1jVPAXqVAze+i+EzKfnM8w/rVH1wHBIueBOPwVQpMI+dPl6JS5pYB6whsf3d2MeE5a6sfV
De7HU8Ec3KuTbjqoAsgh/bRVK16R23Q63UQFZlx3LCn9ynQU17dzCU85ctODJfUH5bH+x6rxosOK
B9855hpNt/VScH4gU3YocX4435h71ujvoTmBpMIR/C9DbSwB+0+qmZS+SzzTNtprZ3ikGgCiIbHt
gggPcdDy9seRl2Yfm96YlMy+ln1ldWRmPFm4w06XZEqE9yzobzVE26zGwU/YM1E0sM2cEAscC2ov
K0E5oQwUbdt0G3IJ+yEOG0Kt38ufQtUuqe+QDZg5U3Zwsh6pk44fM8J8vaaBopwBZNHlj6s3/BAf
VLXCdliipAT43OPA10fKUEYa+CDDR0ckN6iy7dzEJe4hMx4FqDAlWtrfciYPVxxjBSs04y/om4Al
U4u+vK+LHn1U0Nm/w+fDvt0G27AI6L8UiE4glLCQqduN53muB1DSkGgN/wYswL8ymO7IlcdLfTqf
R3j3IsUTwFgGb9z0meZfJUM+IsKvaIGpefMMxRNjEVatugOdGqYU/7oLHnW5eOpnRJqc76ZI/pgh
MriBkzyjOF3w+gwES+f9Uad8u50TGQfdSFrrI3+mG5hLzHK6zP0XmO5lbdxCiUC6iJX5xzDO2bTe
b20k4SCaycvtvTR7ViiqHRwQwn1EVkOsqcuCwETCd4uuB18iIrpxxwHoyhjDehEJNxKGzSd3tGOa
Nc/zz5JRQCHs+Y3elkhCaKM0yLAwuaQ9R39jzsJ0oQfD0FlIc9fZnZepczts9xFk0vnYoTy0owo+
NM//uSYk9Tia6+zukwvfnKQH8e1Od/k28J1rJd6he73XSpEJqLr9wS6agBBpA6NnUsD9+Evkiq/w
P6hvMvAqeIJSZP+pRkS2264pQLxEPA5oExeta8IUbGqWi3dau/HQYF7rXuWxNZsb7ufaoeC6M5jh
YCL1xjXPIiPcIJ2r5m7uzsEc/6I9euzgACXrf3qb113S8t3oyhKiTv6Jq1tTxPEL/Roexoi2tqZT
meVL5FA1YZG/L+GvvWf4+K8ao+m8N8RVf91tYlPDz5QCUsvB1VZdiN952PJc0Tbu+LwOgoUYILJa
7ibAS6KhIhsjUahT4sl5Vggvh89az/pOh59Jl6uCYFJTI7Tjla/LAhQhea76DobuJ/64iRsO9Aaa
VG7R6CZ58Ml0yx8xVCASL08wNNnVXMPofIHotK8ga+E9tg1uIqhaqpnb+zZ5KzNgz8hV3nAZmeUd
mSwmNr+jlupyldYRsVGfsDDvT9lGEkNWPsWPKg9sz4ZilfgR2geXp/xvcmIOvwAWuWm+9cSFlpQR
ksgiiy4LeRG5M9Bi0X97bRj/uEmlcLBJZR/LdHh2QeKiF7wCoGBuaaOPg+itagc5lei1QBMTMPok
mbB9x8E8dKsrRlLGoWqNHVLjiYmhd3uwrvIqu2NyMz8SB6ns9rRYiyRE7QkszOOKbwqXm+mmh51L
9+u3PleSsngXddEslTAc8dOdDG2I4F2U2IuTotVUB5dhk6FtydSitt/cRBOTFRSn0/mM8I6GC81T
p+XlnDrgZYPDfIWndTVZkd2YLuBOs7rcCf5T/I/FkzjinjkMtlgqpgagBy9eZm1UTPOVWGoVVWD7
LajXjbpcrGpFqlK5Rf9bObSuzPiDSPZUt/Xfk+bx60Uu+DSBTw0XajtQ+PcdRlWoISdJ3udBT5MK
cqLxeSOVFlQCXpbdcEUjZ/aVA0mjselRrLwvKNW+Y+1z5RTe3NSKU257sfeXyL8miDdELHlocyuI
Ipj+0lnmfNXXUnne15ofs+2ZoBSG7B+2r8yMvfpF4uj99g4PmKBiRQn8f44C+7Kke0tq82ivaMVc
+99wk8wRJClb5LZs/6G4uImzVcbj+eeuuU4qmRnC3LJfjCvtqKagInrTM3cDbU1RJPnr59dOiaGn
xrAodrp2jvwf6gBh/hZiC8s5hAo9nIfrQ6cFBmTralDRizNbbcnsSk848mYFs+X6S7gEzCZYJBGl
ctLzOfrJnb4vOC546w3Tg451UVP9mfO0QInKSFuMWFChjxw8I5B4e76Q1B0rU4ez72yqKGNmAPIE
p22CV8isGuz3B9SJpzn9k+eFMt9UjSknOTmptOcvkYOw/jXs0XpMdfJlUhRgm6XbAJB97VbYYgdc
g12RgdkTbsGNB/Q51qdgVJf9+TGM0MY1SsQJtOR62TtAQ6AiwLDYFzMHs3zgUS/uoSpwpr8vL1iD
1pu3oqcykM9rqcxCUmsvdwu8/g6l2GMHwQHCHE1cSuoxkAkTWBBGIE2+3tTn3+3wYQ5MRNG77Kzw
CbX2/zbvoOz+r4oaPb8y5dGhI9W05cOw9i6eBROZzO4HCQkiGaoDM0+QYq9FMmD0mSWR1HsKY+Ot
PTbS1DG7iNIGT4ZzkDVN16S7a1SKJ4AhbXzSZaW98WbAVcZStSj+Cygj8RbmF7pFFh7Ys0sYLgfO
27rV1TtmpF8blJstmtutRCL7UtGytXJrWriX3yIqbjypHejxNwi/vtGIeHsvb18M3ljoEpwTQbjO
tLbAF0dbQXsC+GeLM4ji8uBY7Dk1ONvijEUR1n7Hd7oEmN6foADBa3Xv7ZdOixEcCHMMb+FqOkRX
4+5qAgLfdmxkmKz6PEFdjeEKYYtNrtqYg3XqtoPS+6v9bGthC770KBrGX6IanuM3nSuw4X9pfE+W
rQ0zVuJgfKgySPh4YlKgEcJYwiEpMw0UmTIX4VHvOzXk3vltbI4fMHz3JkNvc+0Y4782cX3WaL2u
WkW7DkcDabUMh/WGES3lpagnOOpKx3YLiDt1SPHFxnY0t/bSrXYFQsyI7eZGvynMDD/i9V4Ce6CV
z0aZzC4FD+t96EAiSTiDVgcqJoCcaY3zGUPlj1MxU2CeWZnnGkHPSMaCyC/nQLeJvImY1qigTwlD
ZIGPdg0KuvtiyfEBG4Q4lNELv9McPMUanKzDMZYApSwFj8YH56McvpmFUEmiaG6f1yUhW3DBaGtS
TeaixihIa5bsKpq7Wk0Ljq5E1i492oUwIWzOOTFIBfcKxMl107v0vh8vbj+lOmhZFanDN0rWcpNE
kO7LjhKKz1oj9fofzrKzOLDEdB2VZfqvHi7O0EuLJqflLlYC5SuCuNTZc8IFXJxUOPwlrBfoUxba
wCd7khhF/9Qn+3YXVGmTNQTO31MSodhyUcKOaj2dq5ZYxhAlRTsqYMyIC51+e1tEPhCPRXWbvOVE
kbblC+2CU7faCbl/OcYaloJUMWv5LtWiVlhKc1VRwOVK3+5KPsfBoc2S3PIvuGKTEOnPYTQANZ/Z
Z68mR5LhCIKb+DamiWcsOz6ulzfTnPy09bfRA9thMDZsyzOW4NAN/za+o7Ulk6C1XZnIfaGSO8nK
gsfLSR2fSxv4eK1ZpTs9cr5McyzsnWeoqJx5xEQFcaDc0jZnHu4Mc9hhVad3cBnEknyArdfHArpL
q3+POW5DDPheoVOrppIRZhWLyj68IH8Xw+wnmx7003IpailreM+IK+imxXFsvcqTvYEwdRofkCvO
3hd46w8PrKEXkj06mfMbt6+gE8KDd9+ek4L4c2KKIhsnW26ht745AhSZQSb1QRfThN8dusEyGZDo
ePijj8OYJ+XhK2XjcPT8S/fzcfYAYrueV761sqSBB3PZzlVS1CTaq7azcNJ+o+VO2OjesAVfyhOM
7uCTlsr1oMaP/EPisEi3sFGDe6DbpmLbNbg8/ObnL6hCcczSOFCt7wDdwBVYENA8uoWDm3m4o9rC
gNhRAihOYBy+qLbA8Vzv3Qyw+HfrN8WEVnMaPZNskXnPGTrO6ViX8vKIWTs0VaS0YLyiNwK0K8q6
5ZC+Mp8WinNBWm5t40DMvsCGGyUk2HhgVXo4xKYIUeV6KAJaZ0SMWK6KXZmyfuMhenlvaHHKL/vw
dP5DqQeGMS7iai3+aW9FE3cD2A1Qpi6Ycvr2Ha/AtidYBVI6bJsBPbOp6dBZ1MjRLkjAc198/4Q1
nmqw/kdSddIFgjE06EqI78wiDEFYwqtblrz7r+6avaz9MDtiFmZvhFlNk7/jB+S6n8CDyhCOCQdn
RhSswAaToPfHyFAuix1AXR3+90auszcOTptAHUChwhYN+/Nww3WsnzsmgiLJqXVjof6rB7xPX4yx
Qxdtd6m2uLWmLHQvFtCsWm4878loHBpTdRuuDitMcT4T1qvVOrC2AgwmPsrk3RG2CcBBp9dFmclx
zVVx3jqo0agdrYA2lutBClypMR505CcXyWUOzx06jHh2WG8rU0V8CPCKtwMSR9gGLneoQ+uorDqF
q28hed3z2waYWXopOlAnjcPpJLlgKrP3EEscNAiCNxqOE6+iEs7LA/5U50+9sMrrlmUqbcIBIroH
CamaSefkTv/U48Sjh9cQxCOm9i7LJXKhv7LG2Gb8p/vVm8TUYtjABvrcCiajQeWsjimDTSsnSdFo
qH9RmfmhoJsCQde29QHJk3UqNoNxkc8KijUzaZ8jwI+5+uz2hT69bJ+M1vZZVkny9ZkOUBb8SANr
SA/pLRnwXVv6CSuWgLqaa9Yx2ELep8cBxpWrk+bcysietgNSHsgUD3LmBql7wKxS+1ONYi6suMYY
Lax6KkNt0qIfm5XYjt77ge83Zl+o2aMT92vcmJZSyYtIciiPIH8bEUXdkQsFueFa/HQQDSOGASR6
f9ULT4vAJkOnvPftu3uxtA52NpbuoBmnQd+jCdS4+fDcWEDEGvAEwTHtKUaeA1PdI1s3+CF53DPb
RhUnKbcgIOuay6363UaS0gtSWD+tFioy63/u89BNfjKh7tehzM1Mezg7urtOZDffBukFkT9NUeMV
baVt6DV15aVX0uwNZGeWkiO+b/nzc63//w7w0KXeeV9mnqQT1+p0Pgsj9oERU7ifZTPQJ4QhqT0r
+sj/x8nXIQJq4Rm76e+Z9KO/I+sEtFRE5QHdmzTGtsu4m+xgYFmMhjXuf+aC7BC8jMoppE0LSDBs
foYezoiJTYu4SAwoqaOVQeMexR80wulJr55Xu1vD04O7OMhRRBlvlamTUknJLZZgDvtbBdJ7bKUv
r+wFb+pSNOlBd3REEAATZpD9aIv++beWL6Cz+qncwmMpJwpQyPcfKVMjU5P8GqG9WF5jzW7ldc1F
CyHAPZ4LcvYT4r+cnrmbm6sTwVaHi5mlUwv4XaLy23xKc+9Fl5d7iAo7pas84I3kPHJX6VAA1wV9
Lg4LDtyo8xpl0wZ0UFipNaaOFoXmQoXI6moUMvo8lIiAwN2EMQ9y0bJjbCxD2xyakd2+ZKyCfwDh
y5c9om8b5TyOV/W+EQ2yuWukIbWGeLqz6eUCro7p6NOpZYRoZwWpnMraCD64ksnfvLSGUiz6+pKh
d1fVhLB17HcjFFcJEIJcOCHQ+4DksOY8BUXhiI69v9EiriYmI4mwKDNzY11PloVKB5edAN4bhlxN
49bXAue0UdvH7R05vMpEeBS+Dp1x/eMNdZpfTHDJN40exFuBCZ1ZG+ovxlX5GXzl9pqMVELh0goI
T1Hwdt0higXu+g+N2QRQWQxOLw1c9Fhh3NCe6oBkKXpbWXhO2bTCa57G227U2CnA22n7bSCDMBuD
CvcPtiUfCtTirCTFhadAsRxyCMVm0XUX0t4eZWHr9eAfT+xmVt2MvJXgXIc3Z1SxI6lsUQckVivh
/3g/mtx1/cZwgXOmDLqv/umb3lDGru/azQIEJa60EKkHpRO0UbQZYiS3eoPUExtxqUVh8GCzDHjO
MHgEELfLTzOkwdJtlPmZntxMJRNY58KVePnWi6N6MgF0fMrBjK+wehiIRBYjjyR1t7KbEys0FyO4
crHBPsPlXB15J56P+fx61Ez+TumvkqoCB9mDPO/4aHwFMEHIySq9tGjFBbiBrceDXA6aQZyaFs6o
kGudRURi5kZVoArcJ1bK6T26disexi1eqOYd5Jtv3gN/z0KIOPtb2sM8gfQnR020nYQsHfubWNMF
1rB3GFQYFXmbnw92xGD+V2rwR1NlgEw2A+f7NcHgu+6JxvJnQvcYR3cNznv/ruSaBSYF5axbhECq
/TXK5QjOtFzIITBd6kvZPuU6QmNrMKPlYshC7ZFDKT866/KfUz2IIFmwjr2BFYt+l9Y+R0dzlmMU
Mudh3A8ppkJn9YYm20YCoYvew9LEGTskv3Ee6HUd5s8LnnnWxYyDU5cRZ0tvsI/oeN9z2HbbD/KH
xlV/R2uYI+KIFP4MVNA3JW+bvJ4HijgZtuM0d4+Vh+2FeYv6iiQfAw/COZJpxol65IRrd1xeRjen
mGCHzK0drY2RRHgLCTX7MvXx2JmZU7HTNFWiNU7YOy5CLpUCgiCpUKeDd8H+u9MX0VM25lpY/l6W
OuY0En9BHiNh04XsufzfnH6Q3JKizDRqQbb/bJLQy3IB+3bRMCplQHVBsi4C4h4F3RAglct2CJH6
djra/Uz5+nsN4qu1uscf0/QVi1+ncL9uV0Yj99p+OSSG1w+k1fn/j/jGfYZIAAcSFdQRAAptiWzL
4esqpyNxMVMnOBCM4lvx3VrIWg4jvxYVxkt3IgjUwI5m8UB7qot9ll0ekmVHRmiD/DlMyjLkubBZ
UpUj4ybMAmwDjZiYKn8P64cZ2+RDm2Jg2vkuKEb9OfzenrKg1p7j7F/ZNOA1yJAhLj41lSSZt/Y5
mKd7SdFDbEfoMyuInWGRFANFoHNCeuVDNpSDnSy/QUUXo3e7Ilk7YH4ar2MRYMmWC5kcRcmBQveg
SemVDq2Xz5G0rqrdDyTNbBo4JOuuuQR+ISYsu1EFB1eyDz86O/bgHUQxJAtKlfyGHkanokut10au
OlIPr83zy1R9jeoqoQX8rkBrWWSRmRNNQxRN9GlPTZEWB/TWJOrQXjSFhx6nljaJ1Womz6lECNp2
W4vtHNjA7YLWUYWtf2OL8BddXR1S6+hj3je95X9A/+0O5lwWHf/t7+a4CbPvDQ6ruye0+8Kup3ik
jONyCZHHNs3rgMbqazPjqsdMqmIXWLnunIEaJi/TszV1GD3ZJ/hswjM8wB/qPMZ1qivg5HiE2K1B
kPCfe38d1JgZNdJgYdqcdAR5p7En5RDEeQUClkrmL9rsuBN5+Hm4jGlr91biXJ2S7f8JgzNuDq2F
b21XhyAx1ek2qwZKEz1d8ZEQuJ6i6CX6pAwV7zvdSda0+0Y1/kvXAQM5HS539btA/dfhDXNPDi9G
d13eJpoQOYppB2Mbc1S4/xay42QN5NUpFgd76fjdgMXLuyh2e2Gz1qWehc/Sjkhbu3IKge84TkTf
7+FZMaq2xzkOrHYnwEgNiSWf4by/Z/AzQnzUwl+QHS0u4UKt3a3sYlDEMlftpfx/rMjARTXgynRh
YJm1Dlq5tvTnmdxmoARTKHJ5V0QCJ9eNNLQ5hYKGg2FXflk+GzRtFeCD5efaG4pH5hHHrt9t4o7S
ZSqwEmZBICVzYj3ZnmpS7/MCSVRE+1QSllt+ebeFS49hWnXuJvNO77XcXbY9dNbBotvaZWpHfYbR
KgFrMuMxcIImmPFvs2O63/oAgQqhc++Xlu7EtePG4q27hcHUakhQv/3Xv1wo8WIIq3nh03Ktu+Y7
pEFWaSQ2QVa+3KK/dMtCu5S+7egK12tEmOiqhC7KK/xGQUTTd8HBfeRWDlU2NI5oehVS2KdsS+6y
k/ex/iXM7h894U5oJytQxLAtAbik6IvBaU2hWJHsf85MU+qTafWPbvyq6Ibq8Bq32OKyuAseEA0E
GPwcRJdsKuy3Yr1DcPQagdDmtDvi7nAsBpsV5H+yYIpzrPU1zsGlAUuiJQs1qVETjy+1WZv73Roc
hLssRx89YODa0KOcneLWEBxrOaaC8Pwai57enSJV7OmN4r/cnTcEsL5lWsPwoRcwKYdOfwuPPL2J
4QbMz7cKUHdgYS46CmKg5/S2tPpzeLDQB1hyzn35YjwICjAc2d6EgaKD+hKcRgWN74dYe3JeUG3G
PsTVg1zeO9Xku1oljEEKOgVORnpOI9wlNALY+06B4wSRGmUJL2fY/k88F4sjTWzFOgKqPrIl2Zi4
XC/wz+lyWpjv6H6bYlst8G+I4aHIxka2ODZi9AJSsL6UtMWavJW9V9c2QLg7OVX6gJmx7iFpUTf5
ZTojD7BVjaFoPF0e3O0y21sNwAdORomz/hr3km/XH/QUygp79xcxlU+MVkPDVT9T2+iHLPeiLXKw
KZz7gACTIq5+4xL/tidVJf5oWOmt+k7rd1OqGsub3N3M7g9E6f3IPQ62hTeh2Z79dYB2nEIK3xYJ
nY9B3q0/uW9ZV+NXxP7ufUi/SIf5IKg9XKecj/Owm2teF8OGSPkAZr03JTC6hh3RX1UZm02Gkg4c
bnawp9qnuI60elGuKlJVELy/D4y8RLISw8AfowjdOTG/tQ8x88iM/qq5/p+dUN2P8AilkewNqYVr
1T+OZRC9nVChxzz9vh+Pd1SKrhgN/CKtn60lqe0DFNiN8lIdoLXFExarxdXEjmrKBKjiGr+W/vxS
lUbY6QUeeeH11E01Vaj8/mFGTxxIkO/AEyT6mbobhTIJt7jKKGlMxB+AIybFOnbhLysJ73KvOYfh
gJ5LLY+qcxlwCAGN9PuPv+sCG3r+IQ9vRNxL+KNsBaquEOo388Hmwyks3brGvBBCfEpeT2mrzHfo
4+p4NfxNSCzGJeGI5f/Y7U4vglQna160yV5I0jJlhDH/9SiZybuc/Ah1imTqgINhRCGBjnqpqnu5
EnpbW7r3rTjPbgBLGnk21qYAxTNdRcyutVLM2EuP8J6pvw0bGxJmihAdyxTgNlW8qqnJsPvdrWhd
LhPhOjEKxx08iVUMnHfomyZCTRl+5hRVtSc6GKJV8kbX0Un0Q1nUq/nIRJQLfqpMYAdsvZ3vFIC8
3ntJC3Jh8Io0HcnA9ovVFvVqLx3D2dX2KGCqmS0LMWDPPm82dPQQDuC+4nCJsEtG1BbWXCOpLkvg
yRyb2pVlzsU1AjneyDa1iPXepEUHhvh83wH9sjsY8OWb8xGfIyDgWu96Uz1zoMIfbEBDknijaznh
qz2C+W/lyr3sIw4/EOP46qmvME5cxTLI8GGS/QCaGRxMBlYafS6E/vvPFy0v4Lr1XGDCriQTHEic
CM1K0i/cqwRe5ctKRIMZnZ6k9GBFWO81E9wHyvx3YV6nJJklE5xTtgppannyJBDydq8nYSFspJA8
UsdPY6Pt5pfXlQi9Z1cPlBxMwkeOBY05KVJFseKwb7WkZk9soYp6NIMsC9ZWalNH5ZKNUb/lZKTM
vrNEdFa2LUg2RztatwK87NB2CV3yoVza1lilY8iJnFdus2rvMnnQQwS2J9M9jehdrRmUg0TlJZvJ
pl01cxEU3xhCHI0/fdnU4hihxEdp2cwutw1YX3Lc/h6RV36NjH6v9gMt6NQPu0XfNNuUONte6u0B
81n+QZJQkpZgYi+3PuADHeHkU28Wk5RONdSAETAamgSjJdo91oFjeG+YF/wWkDVnT8fiRJIeQBav
Zhi8OcZjuqf9yv2UdAG4gY3xaucysOHcT/7I3YAO6iDWO6v4u3uDkeJ05u3kgau3mcklZWDCbfMY
csqDH/wvB+epwcpuuOY5y5bHSHqR+7o54lD/P/0VxNTBMvYxUjlJ0kRzuXjLS+kDt5TMNtlJ5uE1
ZbpOQcFb5N84O6nOn1bw+RwrEKz/UaFs5eGIee/0guXN6Vz0YdbrJo0Pd8NU/via9D5gprzWLUlL
uzrX65xiEHv205xp4RH3QBuYSpFxyvsZGjYVzlIlj4lONUw4Jd0LwUx/Ydy+kiUp+xzd+m/v2t4S
m8EMOw8ngRdEl6TG1YaCjtUMmdVfPmrI0mANWI/aU26FtQ0Z9ESg55AHPGV4HP0P6ItUQx9ngJ/w
BTN7GLufCECrROp7MoVRpBrLOt1HBRYi4bxY53oaDWG37EQTmQRuRiTJF48u4BjBBZ/h+OU3Flc8
t829rXlgWjvGPotmHW8HbCZL+xWjuYlhp/sCltqsjQB1K5ENHng5d2m2BXVgitXKEJeHtciME4sy
NZTfj/O8aRFkQPGFwFgI2xco95ab67Nv2sDw/fNOqxFjwY5NQ10dWufK4i1LNKhcbPNeM+6CS3s5
GNypARxghrvef1KySdET6QY9vJm2HQcCoi7aCT0OKZtkZYWV2d6j6O8Mi05n8qnhaC6lhaHdZp9d
7ChlBKkU4LJSCuk9Qe7l0CB+ZlhT/U48dSXpUU/IXsFwiTP59nhHeh9TldipW4PIGK6CfCbBAHzf
rHEBlqIY0U7k+jSnbjOy5JcM7DJ035N4zEASlTawiqp7H6TXvfEv3NbICuz6G+0vVGstcp/Qj35I
HULzxgRQknTlXggAEl/6kKLQNI3ZOcVkg3VwklWU7McGI1dedV9e9Zqf/Ms8BlmoS2Lrz/Dz9UHA
9wPwnxa6w5BBwqMUkuF2v0Du0y+N4Q5MzZYCaeLjfRcBGALAr8N6884+ceUQOZOroM7Ca8BCGgK+
dqXHQM78y/m9PkcWs1Ov+3PdlmkUp6Kw0VNijIFVF0S6pNEQ0NzKXpuYf28GfbYQ5vqoU3GazsZ3
6E3TKynoiKH+D+LfPeUpA2KQLgrA++GtiJzQRAqKqj6M1u7OAcyhYkJOjSGqP+/oW1betwB6l0eS
1MY+3wgS0KiHo7XiuGYP0hWoZwtSS2ednRlz9QcEZ3deoaN49a/CpntoIBcBiEWNDwUoaoyzYMaw
sP38TO6LiDD0IVbUs4eysFBQKOhEY3jSotujVqGEGfq+TmCqHwaQgjihMUqlHsV2cthgbZ5QyMUu
2qHXJpRSAPpe0q4Oyfae3EooEjlqQvAEVDV5+fHcdQfsjbz1xEjIphCaOS7u0S2Vi/TkQz+BDwQp
kFtWcdfFQ6VGejpz0REUN4sKwMq8QaYwK9UajCEa8ibKVi/49lnDTv16BchhKMRrT3u7gsoUNrNq
E+wiKolGZZgfh0z1kpyuFCKaFYlLq7R0AZIK0BwD1HDU1fqs8l0N8uz7eITuQGruIQ2TI1I80Igh
twSYTC/IuVMShqphOvMssLzaOj314mCCquQdEJKON/BLCvEcVahv67QWVHhq10Nm2hGwI9J6GxUc
SWF0Vg+KHuGItKnQCNyRLEF1LHrZZanKTqaZEy1cBfFdb39vit5YjX0OZ1VXlbubgbXIVXiGoy4x
0KolpL8ObH04V4I24fnoiXrFlEXrWVgerp8cUWZC8HTcc5Bu8DZ14JcfiKCLm5yWetL0VSxp7vq5
lUM51xrwgmLWiS3IcVU9/R0ms9woI7lar7e4zeXnhSp0YcAlmhBHnfB8gKLohs6sITGabklDVIWp
V2ayy/wOxFHYhNuUywNoIzBUcthdz7Lw4mjwo3AXHcJyaqUC9fryxbe+ywXkrYfRMdkbPAP6EjgC
MwEKMVuFD7Ts0AobvZV2j+Kw2kVa5bjIWzNkyH829tMxdYmvFcVZ266KJnzJq8oPKYxB+hhd9VD+
WNvseCRKUdKUVTg8V1H0mxYjU5vC7g/+jEmV/L9zHMRfnQyw0HAWsikUKNVKRvUAvsAG8LK+jNVx
nXlV5BMQ2eKgkJ+9uUrYuc0eE3/bkbccQfVvGXmlZOC6ysYbZkXZkWXdRn6EtCW/fOIm/ZBQjNwB
hLiNbjZ36Sr2uQX6tE5HtatRIsbsZyjCruC4xZ/GXfLiX9zjB3imiv8A1dHQI4X9ohx1rV06sYVB
SKgxfwDcUVXohl6XXiRVIy/WZtWORX4m8KNWNPLHlRmHIFxKWZa8ZjcKOmoseg0eEX0dLJWTPZ/r
1AlWAgWH/4X4oYifZPbOWX+ht4V49cr/jlfhAtGOgsBGC3kv+wUHqB4uieIMC3d10PZaffw6woc+
mX/UklmVMRWaSCokTAky5iqdWEPV5BQ/BA6StLOE8AQOnI0+rgcr7jfCeLnIqcjxdcdsItIOcDHe
xl5TodmNDQ9F9C7sZg5oFr6ZIv2eU2Gy1twxJJT4ya3Z3dYpfUP5jkwIKJ06Wz6SYEGHXnqPks1C
gac/QjuSqwllZjFGUfAv3TZ2m812cWqSsAOIVZrA/2vTHeTmF3IkFFY1IPpY0RdcGmEHDSzAkISq
A1EsZ5K1gHAIFCCGEjZD+4pqPBsE8OazrN0GRZXt7hUO57sxZOBdzJSLdEjHA3rtjnahulNP8WKM
QtenQ5cgrjwsuksEyDO7hPh23iaIKz+ZukF8NMszmQydXX+0dFBipMZkkLaOOqQaPClVSzfiniOA
1ZUowNiwgo/bE3AoTqzcpJqz7kCc3LIaZRUrcK6Z+hGcrg7bDCkjfOFLhEUgtkoVeCYI8610Z01E
uhcN5+TLieBSCkvdZFK/VPhAm/goAHyJcRTTryv+KwGv4N3Gj63gSLQTFDnsgnqtmYxnwBjfh6mk
ufn2key35HI4p3EGyzyuuLIlLDzAHzKIJkt2skHkjvmREbm5TV0JzQGqdTMp2JnG9l3viORgL2qp
U8mLeA1nyR9FiFUHrhs/xX9MwYBPtjDZBhnoFvxGA1glWD+4yrn1M3PXEBvyIQFTma8R3aM8I8rL
vZ7zz6eaBp4K77oM8pAXmvROZzjGb015uevPdgAK3bZeRKDvrCTJEaBlY3OyJ65k94Jc4kYkCk9T
ZVEPZL5P109Er4CUaQPw5QdvAgFLAuV10hdQqWdRB/cVtLr8uJYzhqOLazSY5Ti/Ma2h3z6b1rrx
YJjZvqiS0L1HuhI/X2bxdJXLevsVixMLL+H0A24As1OjtpsyF028lZCIZhY+W0tIvK2wVCrotDMS
c6ZFwc/JsJbVLUwZR2wbyqtAURVvpuNbQzc4xq2VzIeMxP6Srik8ry7h48tzLBi8zQuEZhWrDVRQ
BUGkCqttSYYlU0B3AOi+44jUocabIhLshToowJWD2p2iGWh0zdMdgH3jEfI5GWAPa3nkmVemz7LU
2fIdhjhiDkQ9chT5HrtCS7O80olh3Arh4t8h4NdwNJLWGmJIMszzCG0mkI60VPvb2yks7ubA0eyI
4eBktkNOJtyXd8kWIePwqPkhG2GNK7mSEV3FLRc4YfmZhivSinJCoewBoNoyyetsX8tV7eoE5WzZ
75JrMiP5m191cRqixR502mTrokMTGvWH9+HMst4B59en0dSj1x951OycMrZnBc1bD7Ob6VgucNgz
pBxX1oBWj95VwzgHh4gUBKUZ/O8316qTIj8M9ju3VuSQKIySfItLO6QSzzGE2xDKKOIk53mWaNLM
aL3aYHHWTtThMfX8EOO8yHpS4QSmPiS8rkTZNnZpItVUKTngXAwAeha/sPSSSYPFEY+0d8bN4rrT
XFJYrhQghgAdCGtdw4UQLZhYLrguOKwI90eq/lc/tABvP3sVGPtql/YmpqO92evb+g2SiAuz1I6M
+IdT//3PmeJRjVhTfWwRMyBKZpMxcwEeugATYn0zOu3/98qQAmGuyI7IK8Wy+ugjpNFJKwAszna5
ELDQgYRYb45kwSts3tRqJ9Ep5zE0PCui2WHiXcfuRQSbuRt6ybobIxsqDg2VBAzzv6Mc4ekT8yQ0
JBg2VtMj4bwxa8NYJbz1Slz4R00GOW27TuR+dxLv1b9K/iri04MUaFkRrw26lq1kPkv03iOWmtP4
ctVwkZPXjAiZXNczJQ0k7ts2BTzaXGPyuUUvjIIkp/N3gnvx82J6wCyEAmlINFFd9v32IAEFZkpg
edb/Hxl0k301kNOEVvQYchbFp//hdxxp8BWjTf8B0txLGdlZjWS6YMpUZqHvsuK4KsWCiGnDjmPr
p0Al9QVBo4I0FjDx+SoY7berQAUZynQPQBb6HndJp4ll1BPIB8BqNepoou1KatHuhDud7u2NEARr
V2ltrKLjoe10eaKp7UJE6igZ1nra2h/8BSvRWBpcrXk9ndLwwLRke7dHtLEMTfpl6xnJ/rB3ftS8
SDkzZ0mFBehigIgJL4Vla8dKuhQeYO/B/8oaN7ECUaN7t86O1IrKDXbf6PaFZcN0Fn7xZmtTnXEU
1Lc7ltYIbK2WogQWJ6OBJz6viEa71QObeu8b2k+tQAVmAYqhMOyU+Ync4zSN/+10yss7E6OP6ZNZ
zFhhdGxFzuCEs/YZlCx3h25P9VnVrONQSdCc11ZzCom+fLC7PYAhRuhwlL6ubJBGf6fcYH/BPEVs
zl3TyTNoO3yl6n/YRlN/B48IzOgc3IDc7kvHNxqiDJg/bONJPloXIDmFK3/MmlczonhpMOdmQ7Uh
muJOgPRhafghBaQ+SLF7DeOFAsNdiQkY+81ns1Km6akiyIBHGZgH2HEAt2dzEFoUd2m7eGmqXZYW
f82Mzn6TrxMl33YyYCpY521yz0ZBnte2aWZdUQLqPEQX60yq/U97vjL22HIvh103a9MX9ZKMykNO
jCWdCO3+GcnqaBrAVlNzp4fvpOsFMLnhx9Z8TYVMS9P77zXR17Bhazv7tUjA3LuzXKMkQRIqpGtW
epuzT+N3nqNhR5l7GS6lb1arnuB/0mCIM+j5BalWNKu1Ie3TwreGfsOBqNgf60xSt8/P178xXddB
Szbw8EqhmeT/bB/DoOQjjVxT8YGs3lNxSAfgRReBlfFTVRjprTSvqhfL0OhlWWAk7Bf2D5LNue4h
jiOlCibvrtDQAOlLunheHSAdXtVMCe7MW1A/yFXyace+NaG6BFtnvyBMEbjRiF7A72DDOdC7nYyR
1feAe2hy48UD77/1rYY2oCHi8Qf5ySkSA2H2AW1k/w0UUzNXkgrVSMFnxhLVrTsao1Wyn2EmBlP2
1fZINrk/XWtKj2jSQk//7MMNlOLECGXJeD8I8pv6sApGHYou9H6epCImFuV/GxYWbJCaj08gVL0M
HCl8HevWuPOJNm7lsPSdsBMG7tHaBm/kWBQPgm6WDtS3Z2uSiSEjxMhcz2dI6OJvSR4+wZ+WuvAO
EoTyUL+Sy5QaXjZDEr949TlzSQ9kpWEQ43ulzlZQhTHGp1ZXjlNPDHhAq67uEP8lQvvhgOCP8DFk
RoSYKOiC2yG8fZ8T6sQKpxjjXQvBGLUG1+tNeptaoirHToGrAJHtJ2lG/MNWbpKNS1aoZpt7RL8J
U6wovsD6RF44/gcyENBUNbTVO8qprV6qSMK0e9AtZKaegjGc240rPT2ELp9rrMCVXjMdnyefr6Av
4thOjXPnjQ2dryifwKNTtkEEMdsvmEbLkTn5L1jBGML5rjrAG1EGp9Mvr4enVz4iXJ9LOcFF4GDC
1A0JjYhQQxJe4zn7ET1Anj2YTfPdmFXmT9meClBXDiZN1T+j8if6+0eK7nXsOKanZ2IAhW1wdwlb
cF5wCxLwOCfgZpBSIhwU7p4mz+W0PFIbj7cR/t3s9x7/NR8PPWzYu7GMJLFS7vPbUijEDywNEE9L
AhlGeXQdEBM/JOr9DwMypQeLNEsf7qY+rd16lfCj/LGDjUZMKLP9HyFjm+JaMXPxqSRboAXHxKGS
cD6YKua2NRYVsn5fQgyp15Qu3Fb8lKFQrAN39ABXoG7wE+UtTaLNiw2tmGn7hknfyJ6PxqpiysYW
xdQBIORbssoYh3GqZOIJzFbWQ/VPSOQm/AP8wJoRyulAPtizz6pCp+T99stqxsZ6W7xRF1ifyc5g
C+hm9ggYnqUZalM+e6j7HScTcA7iJd6hLu89X3XgNAfXAJZ5REKau0uLdZI43PCAcsMF+PShxFg4
3ywuQeoy/GwzCEkmDyUWB4kpYAzSToSqmXi+EvrD0b3Lwc6zVUqvw7uYTpI9NV7WrV5IsX5afi4J
AhegI6o3dTOS2cFhs6K97y7RRJ53UjYXLeXLYTbidzj56AO6QIvdF4wrryfs4xG6q16PwzgsOQjA
d5Z58YpbjUxAEXxskwiKjY3t6rWeo4AMIVYQAINLFaOaj0ifXJbEmd9Mb7K19+at7coS9Re33DKu
w4aJCAAzAO+tz8YPWKIYwgnE2KDdey+s2aWQzLNw3E1fFD4pQMR4oGOuXp0R/Eh696C2ltqQQSUR
ObQQdlgWft1t5ol5ZDvqzwOaixuoLhvajIs9mIg/LylBBxfzmPle94Rq1poU5ArDaf8/jZmQzpSh
8/mKi2IAc79gA4xNl7/3+HpWluDQ246CATh4g2+YHd9NMjeHDm/OtQNxWqKIeQGUiwCycfMK/D9e
b70D4tcXwnARmwhQHotkFdeQTf3XZATPqxnbV5lKY5IuxeCd9dZ2mv7YIUiB3S1Lzrl6SqcSGyaL
UQgOKjfKLLaKMO8mvVMluE3KMyatO6PaGyHwOpCHSrSY8V9DCmvv/r3ego6yN98/GvWp6VhnddQU
+vLH+a53U0zzqKpg/06b+eSvhD/8ibIJ6xFulbyKMhVUaL+gXOfteoyHJSDtZ7nhZbhDRtJqnIQt
NJk8Lkbpq9PPMMoM48b5NysAGR+TD6me6pscf3IWQPDs4ZzNOuX3hrsa6UucK5GIEAX/LCXXUimX
t5sGf2ByIAyw/OJULEHGVBzLtkiPiG0ur6bRysAxSn8bubZtIYcMz3TxfHu55NxIXxDT+GqESOQK
IeN+aHi+VXFywNvoTsjjuC/A+6fGKolmmfatiYnX6powG4G3weQMyhw+uoaYoqnDtDvbt/DS2Vhi
pkqD+k1s6xDTBeiLuV1BW9FB/zetmC+RGhNMTIuz1p3t8j09EyTwWi0XkCM9KmBu3XC2nwCF9ph2
fLafl6N2MQbLu/iPmxkqkc6O0PZp1dPd9y96iVApcCv8wUqaROPy+GPz51ESqQGrsZob3mNxtJYB
mIj1qJTT9PChLg7KRPznauaS8CG1EeW9ieO/a4df/cLWHOB+4/5y9wpLNOcu3CFYiqk4eYmA8LmX
iZ5latRS2M3n6UHI6Egk/uF7JHGsp3iKDR+yYWqMZCdA2r9KCLjhOFTIg/orJktEC5ZODThmPhAU
h/gaurZrwrJQGZl4YoEv06R9D4BUXbaQ7oI1OquBQCsVa7Crszeiyr3WoxUuQSbNPtHCtiSA9Qhk
EeeaAnP9sr48aAqPAXDT0/nlIPgk8LeR7vbIsexnPVYHInhg3tOYtDTmHMMnFh/6smJDcT4Y0Z69
8iOKsb9GcZMi9b4zaF0AOgBapP3uft9++4PZrCSieNvd407EHwbtfaIJdBT+6DxgRVdeXcKCZTpK
9vRqVlBWYiitdwLBdxB6Kzmlmd5qvCYYwgMQg8QXVOc/N3bVNkfFJ/RIqVJUA4xCxmIHi+8HK9Ru
aUsWZETOguBO/9RKZWVUemD0jfjOFqB0REwOHPWXwyFRBp4ki3puS7oS7Ieb2lyW3aa0mf2hWce2
VNHDF4gVKsGHveEZU7S22tCnxymax8sE6EUEwG9yNeut+3/mpVOXhVezmGnaI0sAJuNmqtkMz8NV
+kT0BFi6UywDiQGxJU1r7tzf0MwTr7z5SSkLisFHMWmf+uQiqxbYgCekh6I/C+B0TpxEUltnK9sE
ICHSl0Vr8/7/jmz0/zNzAVBQ0unbSlTzcVHDY890XJnjwbmKYKuQLFkRrrviNrsZ80eoM21o7soz
WYlpmK/2lY3hPlUnBEIzFAoGiE0PUM12SAwG81I1OLmykJiYHP8r+cpn/a4/oTZ0bVslihVSL3LH
c95yBE8+J6svqDF+eGzADgTaOQs25YPWeqe0ZF5IcpYGfb4gLCuBxt/sTmti7bhT66n5y+pTpjCp
rYPLsf9rCYHTGUOyDEce/I2hJGxkfZDBLxtzNT4iNdHJ1FmTdv0za6OuW2/bpancoEi8aAkCFQ1Y
wZd/dGN/FJkciJoZ/VtiLzlHkT79n9d1aEiaiFxUzGxtHiJE4mriFdK5X9M0ruR42ya3l7+cVU+z
R6PFj1E9RZ5uuHumwF3SIsls68HQs9MiOSV7t/Hbao5vnSqvl5toUeG154kMF3M4iOtgIRCLVxYF
+oh5QSBiisIYG0RgIQHd39ocaC5oWiKmLWhryhUR4lsaF4Dx2ZyFKG3KwIs5sRoAIbFWrsu++zOO
6bFSEAmJoX7I6jWK5EAPdKM71v1DLr7xHZL13OxvL0sb2rJgb02fp2MmtlhN27W+9vHJzNxltj3o
6oQSqXxpDt8UPAGS226661nqwlp9NVWR/iz3xdZH8mXn+UvkPd8HBTLRhfYvYNcF0IHbs+m/KCXR
tljhF3vlMbwDRTbVynY9GNlnitY9kiztnJrv1vnLO5arNa7uRrF2anoiTneKjVDAvKc+dQdKYtsN
OkuDbt0pTk5GTFbYPj+Kg3yRrUTSMgjhNGOeHIvpMjEOWrsB3JIsu6AOjFg4DPXvQgbvRNTklzyS
azEe9MK6IaWbXKKG8An6b1cRrcbN60thX8R7WRG4lxnGiPmcIf/wq8i+Z94nvU8Nn4irvytbadwx
ZFUv8z7Cs5W/JNxwUlMJAxzvrouWfYO9QAZuQpWvFlGoMF1tf0axg+lb2Ce2iMPZDUtgdvZIHkcN
lHFPhUgEiSOEJiIY6p/bVWJwqqCu1OSL0FIzTMBNw/QZhS5i2NJdcLd72AqYQfNdLsz+CLCutn9d
6pF7ZPs2w1cMG+TD/N61ekex6jMrqv85gpufZtsSO//j+oa6YTUg3Q8CmLkT/FNl2/rQVSVpRqnU
rXnFSJELu3j5VDwiZKpwjJzx99UoBHQrrYWbvzuKH7Os7r38EeGjGlou0DL2xv4t+KVTlvjDK75L
f6KvV2uTHSXyOOD2E4K1YrJl39C7r/o7aTrQP4krYZg89NMKA3Du1X8+06urE04go4K5aPtxeNF3
ksbY7JhRi+V+E47PueELvHO39JEZ5Bdw0mdiPpQlIbLpMJc/BXhwy3JOxAUZtFOqYrv04d3kg5ff
PQAeOL4MpovDaydq/jMW5VD87t5SNVI84UhnBDt1JSXKzkva6CzXhju64ESyoEo9Ayjtam4DeLfH
Y+4zgjDxjkF3Xu7zhdI9FRdfl+/HggLDUmokjBIsW9cNS4iDJ+OtPGLgKawmF5+hzqpqmeU5MGr1
w834yJDMa3SKAhr0BpK4327m7ut4wwU25DyzK4N7ByILt56pbxMcYecoy84n9RJzNVP8LjpcxT+x
WnJrRbCydC32NgJnW2uq3oK4ZfbNfENGlfwD9Aj3QKjV1W355sFRYZzcXRRa0DP8RfZU0GzFr51v
/G4VFmSOdSJTD+i9/XwKPFoNTEbh8XApH5v1FrGf/0HOlbZxiQrn2FwxS0rIA9AqAT9wUL5e7irQ
4OiQXEW7nN05CTFEyjrcik2TEwrBki2clTMWe9QUu33mX05I/ZlGRmOD4XAFI6Cma4ELOYRm4XnN
m7YRJYVZq809DdW4nlXmzmkF7hhGye/CIax8T6ibWfQdVHEz/2+VOcPU3B5Xxns8vAd8QVZDPPZb
m4Q4l7sHn1V8KR0LphnYV0cqCbRbGF3ceLTvVZJ40TAyEPK56shKQon5nlO+b4XiRNIE/MKIRJsN
qbByefpsi7lcDKZz/kxVCpIXoBcUYaRctpogPKWL/SUrnwSA6C2pxWBRk8o6hZAqzF2gEwcLWgaP
vssWaZm7UCurKEexLXNURqwFwrwYXxhRgoOymEDiKG0QPt+I6jxp/L0EC0HeEffC3g8GK4MEaMqe
KIn1iIlS60gqqS2ZRZ7o3y20e4T/Ssb3RRBHB6pm9IQ9sF8d11wWxk1lv6qHJEXhbmHGG2M47XUi
YTT39QQzAQAt8CgovKQ/uwXSEsq0SNlt5c5BwPvSwQ7GACGEId7QQ6ojHxN9HGoKxxfU3+XHRxqs
yF/JszFG9uR+7NBhaE2AE8Moe8It/VxBvSgaSYp/peg1wzUG9YglYAFI2NmxID3TAf6nPv4uq1eA
XEjxgwfc92OLdtXRWcx8NSdALi5ZugyuVrqHxoByYptSnDZOYTg0RMb2uBGjIoDM1qXr3LgyuqUI
GolW5mzovzMJGZRGBjTB1viLjJQo+NfkVkRgrJzEuknVnDdlJqy73rXEIL00PJ8Eh6PvLDGN+oHt
1L0ubCATGDn/lYnnnREW4QcT2/olcxGOOdluxfO8njTqWy2c1X1AfW19DZ41hJc1tonKU2VdAWic
6kKK/WVcw4ufi5BRAWCTWKa8XzelYPnFMXfDCaSXnWCq9klRvtka8FC/Y/4O2+C6ZHEC/YBWTWAL
5t4F2d8mz+sWhdxozwJEFbF285+98TVsTfHh9eKhg96RrEbHKBQmLT3YIw0lqzqeog9q3951jGCr
GlsrVhdTNEvlPbf87q/Lz1LZ2Mm0JdWRWPg4LmjRGcTw+oJsyAEuFM0jwyUxbHGd2wPxRcMkHpLT
ZPUTDl0YeCfRBDtWW0ytXU/JFhSexB/gmJSdWRf86P42p4jFUbLPW1P5ZWxQOHBZTcJHhznJMmBv
9HCiJn1IlHjZ+60EgdBZ3UV2N2B2Jyzqn4rrEqlrmVQ/G3L2gzh0FVQNzPP0o3ZfprijX+eWwXBl
/Ul11USXWKIzCRuxrQdswf3r0n2e7uiMsrmgF9wdLfBuiZ2szQy0ZyKFsjGment0WIIfvTPjyK/z
PwSsOLQETuSd+EUXv73FRrCJI4TnkJpnAQrh2550blVsCHm6xSSN8hF9sqUvq4Y2aghxRmJZM1In
EnflZYet1LUlUdB6fhMlld8ydQFP+7BFwpHJVKhVWpgbMxDMrNVHLSDWm6T17yz898xtAKJ54ycx
OhR3KfsxO9+gDXtlXmRvpMZ3rIjPt2Afbi2IPsNHiLg7XlUOOhV/MnPdajkwD0JoYJhr5oeaz7/l
e4ASe8Ah63VsBhWDJV2z4QIbP4GX8/MCj4Lc1hkhIKuPOwujGRr/3wmHr3ET6R9bo4DcMOSwo6R4
24fuU4fRp++G3M5/JPpP89S2TuT2mswZzbP1V41VjNKIn/vseeWhRfNwxYSZfEwbecbVpwGVFxcC
f/ZyRYzKBH1JoXA45dAaI+V0efNcfN7EvpyYErN6hvSmiat5VPWvOVsonBqVe+13OHhLuynUkoAK
gJac41IgkmH63woCYEBbOOLIlFi/NSEpgob6Rd79TPoNH1ovaOPQYqpekrBDrn92/SLVq2ubonq2
xkwSqEWzIVw0kpZ9tzMeQakX3tVTQ4jwARSYOaw8LuoH2qD17O+RpSpDRufmNQcId4XFqitRzhdj
SYlWcVZUd15qi5qWRSjVOR23urHGlg9I4QY5rnKdOgQAG6rseYBxGK+tM6+6XZTIhOIOdqFKx9Zm
w80PrCdITpXGj4z4vUvGi45o/DUADw38PiwgUPoVp2uzQszEpAV/zuz+DR9M0XqUFT3SVAq45Os8
lABhR7kFNcRigylnb5ixbhZZdD0ujMeEy65/E8Q6qn0Cve/bvV4l9nG3ODeKpGBBsIUiYy1nihzB
zNAZ2Svn9oLGmSBdeWi8SwvCPSxkEtVE6s0hm/DwrmKC1PkCet6svET+X3mSgKc4Eh2QxA0I7yXE
8IPg6WjeKM3dM33OnFj15sbde6fptDWDRsUp+aVrB1NzSO607mrGboihM9C8I2wTnkAxbcD0sROR
G9R0dYXzwW1ALST4uFxKj2QIXawuWIzXcdAyP2l1NiQG8BWgiQVwHGSoIMwBmuaBnTdKjweS9RjE
BvtSKyCQG2AaM4RFzRH2n4rwazMjJKGauHmjxMsfdmLMwEBS34mJzaz87mZIXgaOwsLtHQZm5Z91
d7jC49s1qhFPSKTysetPKcQHMHPIzcupWJBrLUkkDq0h8N9+XJSOBhWM0MLbDCiZSbFuc6ksvpqZ
zRRcKTOVexAZLMPgmlXTTu4elSZGZQVgNuE2k9SCRX/imv/9a7aQm+dAMYjQIAV4rZU2s/+OrVLz
drCgGZArGE5k961Z6WxKlfLjX3i92TqSbqWEGwfAv1stH9JhiZpnCcZ0A2CCPOJFGaelNV0w2+zh
3ZhFj43gQohbIp0lMoKM2yOfxPS1oa2XGMlzCjh+HXRoapWiQ7DK6HDJkyNHcH44kf6A+Zpjg24P
1kyf0O/Un3H9c04w9W/AcLfid+9+1EcDoxD+ENg9eweyZMoojPAs0+C9vdkXRW3JL+r6xsLSrsek
YLghNMsJEpkXcUNAJwEimPCZ82fXeg1H2tDvjYPxSxx5hPo5MXxQ0/nyrFSJg/Tv4r82s+sLldD6
mea44wAsjlgN9SgUCa52LeFc2xp+LpoQSMi00acNmAVlg1OBaqiM7/fXhLzIL1l+P4GF7CaLV23c
nDZwt1xq7n4/5+EiS6jzcsxqRh+CsgqKkvYxjeBUYMRG1LHS52K1tRrvFIM+8uG/LMTckjqCyH1N
hNf4XDIyEMwZQJVWPUFVMLYKPuxn+eJsSlO+u4+kBFKaWZeHp8bPl09IMKJWKf+NmvXEPQM8K864
neJEiHlxInxXPM2hSbqpyBWWFh766dJ/ePVNRktCeUtAVe7JraPewdZfRJPS3uPp7N0EA0vTecBn
mKwPjzWJU0Ls6O3jAjyu7a2QJbP+g8pHp5vgyihpcemD7M83/4V4LWiJvHNTzl2yBwKQP9I5LGj6
tc7ZjZ65F+e9gVPMD2P5xFgDoPEm+le010NrYJOKtJV1myVUpg/TkvOiUF+E9R2eGsRJ3YuddGOh
EXcW3Qt/utTr42qZjchyJ+GXR6bg0DcZgU62dTS9s0bWbX7ZMZC9abI9jYoIuySOdCcbvZ/3ZGwY
3sHUenWKKcXRJ9/+6WX1UG7JhZuYz+c2kJM2ad5lpKvhgPSwL0toVSF0J/28r1ku6eSNlNDSzESe
lbr9cwfaeFoRzrDL5AMxnGxOPGMKa3ThNYhFajayf7Rr8VoJIH9XJcd2iA14ojF1urZlt9rAg12d
wxpypIVOLpcTQc+eOAjAqsoQS5frpIC1b8d1ntqQAtQnxjsLH9C5ZrpoM1EZcHchVZJIb3eHpkn0
Syp6diOBy091yIEscd4NfWvItyCOMXJH3fzlBVT/XPlJu9QD6oC8EmabE5lwFcUpdFlVhYqrDtKE
KHP6S0Vmn51w3F5HRd4ZkusuCTOfoGFnYYlE7JgZ6ZQb/Wgy57Q/dCYg+1zWH8ojRf6pGBf4LxPb
m+jCW1adwDGC+epu+K7VPRWv+sx998a7QiEdRdaAtp0aAng8pmNxW3ihG7HUA6gGcqSFwIkkMo3n
ZWZH1eqgF0ZqdokcVYuUcBpgVOIZUvWZpiT/zjwW+uNWluQkpbrhmRREGoH3KhMhrdkH6y0EwW7G
uPUQc8BVAcbhKqa8BHiSZr8MzDC0FgQo8aDOmwKp24ktbFaQ8dqwVNkoVzdMWRlNCU35totU4aGS
/WndZx9Z1VEeTnS4HTLhKy2v1EnWVxcWUMBDDObX4iCdtnI8V4SXQcOE1xudVmvawT512s4tzihr
q5YD0pw92G3f9v/jtfvXp7TJYbo7gx/XQzrfedSqhIw5GIftIiBoJv9iF1DEacxeOI3RgshxRz+b
zBKAm8YMQJgkdlX7iFrs7KYM08VO4lZ0F+6BIISaQPw/xqJRSc7lAlcfdjiIbI0BahUaMZ12Lz/+
fG7WeBDRB5Lc7+l4LIqMq0xvuVqYFgp+saGWThjGvI/vmNnSthi5wB2d9iKdBGyZ+19DEbS6yQ9P
GoLEwz4s3d1Tic1oxDhqLMw5pTLgwXp3PCAnAYjiCcmasIUJDVC5aT4jQ8FT3nJDVjdqbrvKTMcN
HPrfmgZsCtkmcOA+jZvO6PmVPFh+vf3aYcyhUxlyuku+bYUrmyRHvByh1DTVAvD5ivcZeWmzuHBf
XcHX/bj9R3DU93divj/dLhXrztB5Ywomb/4OiZ8uqKV8/Ip5yxVkS1Jkj5RWMfCywDGsLRnkPBbL
mZ4AqrUb8emG4/UqeMeRMpLCjMDNqeJ7eIS0WMWAbJDEC/U1bJEEIRxZgkRiCXum/SlcHO2hFWSQ
DHmcGo9ouwq0zgmeeCeN3v32nL3n4COsPynaUSnOHtmiVMbMfyQwJAtzvhMr9ixvhPTEvKRAt1PX
51iad5xKCOgs/2npQ6TZ/QpufD+gF1y4VwAQct0xYnivnE9B/bNoy4o25PIe+0bE/3/SWFnEA1+l
Y0eC1ytc1LmbNxd9uPCY6s3UJ6g/7K+FKlN8Q1tME9xGSqqY9vQEpHDFz79ic4nhstsiHU2kpgaT
jLhAMcxfQlrNYxHaSL+wAaRHYsJEuKSPuIPZMDtWsbHvZIZPpMjSYuprFbqjf/xDxSdhbA5aB06A
VC1eJ3XwMfdhn/8E1xxAYlSNYgucckX4ioBq5I2e83PUHSO6HiPtj2D6X4CgbWEPFJTMgaRDssWa
MUzBg7D59XBy/diFVg96PSKKNtacr5SDaPpEtl7v6ItRXfXMq+sRUYAMwmjRj7gdNeEwb6RWD09N
dU6aUYlz9nyurFw1WR6NHMng8vV4Jjd/rdMDFDM0uPCOCrk40nbBtwCXKielTafsVjKuT+Nhrk2s
R3ZXPNqqbk21kTKRariT0+lZfaTZuX4+lAv8PQiOxaeXMsf6MPWGq9OLXDc+zYm5zFHkMo+5HjBE
9twXu0j7i4y74QYFZD8Dr527gG3QXfCo74CaCmoIrzKwWFp97Ik26CrNcedsxakUzPFWDWLhxXSG
fUs1fufJBZgRPO7IwHPAmttiXZ/zFDaaJLtsTJ/x0LOl3+c4C9AW3hGJtlQk9mzxXfY329bJRQGW
nwSq5h4pSIVXA55M/MpOh9jPyOtPaXFVbYGhEGz+sKANrDEtOJ+rx6agIyRBSbef1QHRlxsWvOnv
AaptVRP40c0pT2QWap2ovIAP4h6MTSC+RVobfV6AozClIyrp73mTCZ/rwyxMIdTNSbTM2mmp3jbU
fh34fBxwiFKbR8u3YDlBmmqPci0n8TM+GRE/JgmFnhwRU23XA9T02kH06VvJ+I3XtkutAum9Rgs6
yH7v40LzEBSL5wafNJBBFdAWe1vIHDv/AuWWs1e43aI99BYtR0S9mWdZaR+HSNk78JBEzoyOmatS
4EPNZsFkf5gSnx2uhdZW5br6qkTstWK6sdedhmpxJ421kzxkSZSjTAsKm/m5xGMRmKxfmWC1QUcO
locdytbVCE+OMm14Y83vDTI5N66bzErH1hMC/9PSlVmcribbsOSDVtCUi2bVwi9QGzPZRMwu57/E
dM0cgi63NKTDvU+EgwV/KoT5KDaHntA6r2aeU9ggci+YHlUGJmMk42ldY+qq1CU23LcnzIJ6RByh
jSv7ZjOpwCmQvZ7M3O8gCrSy1jnJjUDqAxtwCGbDMUMG100H0iLXHfRiq2fjLOAuPf44zF8BSCtl
NWENy/RhnAqMBKUhRM6zqih3JPnPenM3FqBv3fC/DYbymjeaBoy6LCO3hvBgAZ+ocEZy9sLdi0rs
juc0R/KXXjs27C3f3yEx5/0maKFYVLiuidJQDetY4+tS0dgle7LWXUIkOvy3SqXTbvbvSFtyzqw9
OsEJPpM7qltoWn0ajwPrNv+JEChh5na5BiTsZMux/bZFUfPoKngGkhDfvT5lqbhVpgZ5bCl5EDz8
hNmNBsXalYXsYCz7QGksncZqFCN4zcPf42hm6soKH3NzO4WbMRqonOOKBVIxbSuGxwTJbZGUD0zE
J3s+O4o72lZlMQt/AMQV313K2MAcjXxNaYclcOvMPFSG0BUrOTiJfwqg5UFh9b2GK92Hnhm+pBOa
cFhsisAfrO8psK9OrKZ5LgzYVNaXXvWxEsifSw7gm5SLjgxg3Y9/rIRa5/fWs9yS3yP56HCtnq0s
UDinfSg6dC9zk72TT+EXb5NiAzDsppPZAanfxF3Phxl/VFChAfQkpHBKm/dx5e10ZLCiBqbcljXy
JbZ+AF/k+e+enM7fTLzANU2Cm3CqnIEkdzuVx3aJUEClfC360MICOF4DuOPx044xMVD29Qol52PG
ja1A+Xw6fEBLxt0pKZGQxbSV3J4NSI11jcBJg1BdYLeteyms+l11l41NbBcONTBEpNIxAXDWR6M5
gwrFmfiBENzv4QOF3sywnugaYTm3J0o6hjWTMERA41AlQvAGmE9z51iWhNMKMiNRWEMwuekr1yl4
0sLj/EnZjuMqkJVH5o0LwbLvntwXyrmN2s6TBGmEEvKA+i70i3DjN2iEGf/fmNI9DWh5muv3mMFk
k6vchpykrzz00WSjifELA3HrjwNBvNB0fhiHMzJY4QRCwwlPDAhUXzrpQm0VHVYa4Btl96blHyaj
nsHkJHnXwOe8iZ839yvYOl6k51JemgBx0Dl7+bTa/efC/AmPw0fIo+5It+ymoiwApusw52kM8B+L
UYAsddoyDlZ7gpS4fiGF2FHBKCmcWWYnhHhTyH+/UCy7QiOIZbiKgZ31a5CtHyK4TFH+RmEUhNuQ
ccvEH7MGH65bfMfEKScorNwYlWEz3Kl6v+xOWa4eko0M2RO9k+8XPT5EHY3JzD1K3vZJ2h76i6b9
/tT8ctO90ZrzIDPtw/zdldYFRc90rgFeRn0f8LMUuGyp+6d/kBU/7t58NzvgS8O+Y/5MIk3CEiXk
PTYde6LwGGyJzTRFv+VgA+2Q+2U12XOXZ4kM4IVpgFZ79bO38D/UGt2VpJUcKeLQXe6zenvgG05E
IqkhjPqXbulmzEZAx/l8cg0M5E1T+gqBES1iOUh1tglAVjNsTcRMQdgyLhjUbvQPQGHHM5KlwruZ
DlfoUdt93cfmiZAVw01rT6QUKfLLf3x5GYZCac9Saxxjq0QQbiB0uhYmIm43XXWYx7Y9HEhOY8GL
2lJGHisbf19nzOSgTketYaRqL3pVs0IA4adQj8C+wvxF7J02pZ3aiOKd+rmeH13jdG8zIzTZ8AmO
7tv4AW0StybDwY6SohschDMPLl34IbGHuYZ+zJdJh1zkuEhajP4mEW1ipO66RuE7Nrf+9NAkX8vd
QfT/MUJR3fon8IRiX4TBHmEMY4WPoP2Zscb/4YYlyYqC+9R2wgDtl9PKk1aqbjpQUXog9ajuIKLy
PHrrTZYKU0wqJ4+UwByoVKH84dJ7nj+C7/wn0RpdVscZbfJrDOdWg6j7v+iv/PjbbkeZ7OcunMhW
sEUqY2rt6dMVa9/VJSSDnuUQGqGoY0GeL2PconGoWUnwf9BRIsHC1SL2/DyhyG92Q4jOZfMUSYf2
sU0noIFOJWPDWM12+ohUoFgsb7Ht0Hl2HQOMUBGKI1po1+/xayD9yyjTQGqpsEuZopVpjwesFaQT
ep7UKtI/hFQtQCMr6THX50u8WAXrKhoETCHY/9sDBKHnlMGnWCouk+XjRcQBDjJ7pAwel5bUHz1s
HHgt4Xv9or5TlsaZnpA6uH+Dxb1qLjb6PGhK5nPsybVHogqyfm/y/Q5NtOB4KBagSYqdwjXy0mKi
zUic778beXh2ziNou9Ob8YbtWqj6QMWbtst4bcfr37mF9FXJT03gwBBwf3cb3QoOMOqz4L8FSnra
4IysYoZLbLKjdnAgnMItQktKRoaeepCP7l9IA3+bJQvyD1/vVmWvoMc3uBMdzyQgYTfZM5b1okKA
8CGxW4/C5M64Y5sWsK3RhW5Nfgr+K3OhWer8z60Fcy2ymd4zIc/pZAKFKC3KoJU+L9CFl/HsRDku
gg4hHGC2GoXWyp9QWyNuK9jWlSTo/HDHIse60YnHFFV8hf+vhkBwCvHuU24D93Mr5ldhNZMpq8dI
AVxQxYeikSNGsNqrvHTpgQtt2BxTNb7TmhPbI8v3s6cgczkKIm35tI0/emLljVbA9mLrT4VyLX5Z
U0ZYAT2EvtndBsd/1IJTbE0JiHENu1TqFTeLgftsMy8neJumeQ2DcKiKjWi2XeZSJ5uT+hweVFLi
kTkAegR7COSQVqGe7OW+1blBpGCnNSVJzJ11zl/28yRR4ZaFKWTj57oh+1oWPicvcwvUdm9qfwpL
baen7BZl2GMqRt1kYdD5L4CwictCOXNThb4js+h2qYSne7Cmhkv77Cs78MfExHGOfFfckJTC5m6w
OBaxEtFQHkY33CLbFaicUB1T+Z8Rr55ZzYugz8r/EF8/L7GjjYpSvV1OQNW7QoAayGVwf+Dujtr8
M9PbQPA4HgvLlm3A4dmS2rg942+UOZLShOzezQz3GO3B2YWgDyQ87f/51nOfXhYb+bTdsopRv1Nt
PxcEqOae+TwwM06YgMruxeyL0wvwySYM/DSXrY6SqACzzNJdXzAEXsosJ/AknkGk37SRNwB/snA2
4ebI1mQiGzBftLoY14SdOaxW8ZrOfLtMek1lls1XJWLueOsEeqABZAoH55LSTsNTbKUa2/bSkmOx
/hUvudFGFJSeUOAxZZhVtRojdRolQpyYNVwUYnfXo9NvygCsp1SoHS2L8HmCzqsaElTtcdTDyRw4
EUqxdSduQd6/zPHumCGIzBH5CsapizAzwWsVxwcMkAXdA/XrKra4aE/3uWaiM7VnqJ56UQ5Qs6t1
b26QvgCiqV1JZCVUJYOUvWLHF1tPb++eiNVvqQdsx5YXqUBF6R/CQlZrWglPTz4lk5NsC2mQFFIw
QG0dZqHRmfdNvDKDFxviS3XPiXZWTjzTUoBtIsBOBoMXZW+nGFyJJ9BMSwP0xrVxvbHOYut2NMes
As15BAbO2PHuQZzzejLxcmIloy7WdLccFLHULB+czTLFNNtDmKed74+zBji+RKSiaGwJCmWs4TlG
pXHQR6FTHPmAKdguFYcY5cBkaYGb6d56POdh9gCvPwrmsttBYLFj/hg8/tLBofLVGU060QuG0HMr
+vNI/O0aGVYrfwT+5y9WiuBJqL+fJgmdTnmuWz+7jRQpKyryDwN9LobPqNmYDrPIOUTQnIIPUEkO
maCFtQiG7TmVE6ud4/nQppDQ1854aVJ0CHdv/JnhxkCL/BLytYP55Cq05tlHu0GxJnc7Nl3PosaH
hgX2EnsknuxoobeHk3y9erCZGncKl0RxnnK2BdeCvrgvrPHZ005GvQhJQHmnZMNwWsDFOl/GuFTb
zVJQzF3lEjbq6qGb1tFZvR+h9WO+57Iqj50+GRad2kQ3jlM0lGTERT4lpxW34KoJ6LUOsxBw69R2
fBylVwoAmG+SQG2l9k87ZLQNw7ymM+MjP4MwHqU8DLLqDX8TrUe5o4ipyj/zEz02GHTdEYmih+On
AfbUDpIi7y4v6Mx15Bp6tD8Rdp6a6uUbR3QOEor2FY2aAH6g91a6F1QMUAHn+T7eaZCTdhxk6IQL
kCdgiQC/jgfo/kWx4fTavI6kFyyD5GwUbmIqjf8atkyU1QOoVHB4JAr7FGHGgisfI3AQIErRHEum
+w3i/GfEHxYA1IpGlNjFrFs7BhawHUxTTXgGodvQji4e6sAPi+ccIOVU2jtJquXPrK8l1eSW4KUw
vIHBBApB3uLvYIP6UvYjPx0hYuvk6hedYhGiDoJtEpG11xck1rJ1LP+em8B/IR5p3cnms/MwQdeZ
p/gIWEG4s6jd1I//6+Nw4wZfj8Zl9qeeevbLhK6ypCODFHFmW8uJihgJUM4+hTQXTM+hou8gq7SH
f/U/HBAcrOqpqvOeA+KAQ+hFFd3q8vcsvMCJzFHyXLrpDEfnY3hUCKV078LrrCYBQosDW+m4/kUK
a9zSjP4FBzCrDhYZI5UU0NHJvbh72f9MEUBKIBaSn2FZa8zQ7whzAg4PK6V/CiLVRNn2juME8htI
eMfgb8GH0fhj6QoNM2tovuhKka1gENeKl8PjRNCjwPo1HNkGrOwFw6vyAWA/77nhU6hMVG4b3rCj
YguTWbpFwM/k7GR68y5Dzmyqh0jadcXPbhuuIQFdEcsgxnmuo/fc2fefC6zURJQ8PwVQKys9OpAh
rZxIHZKAl2lSSAfNGhm5BtCGWT5JQcl6qX+l+ZyeT+JSbcvmNpXeh7Dswdob5fQ1Yi7C4WjBTIdR
3oTUiEydQoNtfIs5fZFu5ecIdzbOjIXbpWEoKz2aGC4TIObeRaVv+2gPpyIw9ynmc/dHretX/L8Q
mTyu7TnScrHeOFN7cc4IIvT7g3lLoh1YMOoAr3nLvJYpYKON4nbhOlqizfXhob8JeccXS6q1Gc6m
XKEHS/XurlLlXb7C/ft5Y7yZvoSAuM7BGC0MzXQX70Hw8l03hq05NliGxVR6D1bjPjCuUMawwA9k
T6ScajeRikLJAlxMiOMJS+jI1udGsGOAwsKo+sILbPqUOL2OgxfWwIVeb9qwzI+rhlnoS3RtZr2B
rn9VoBgQro0OZjX5SH0toAd6Qaa/I6V1GrE7Mxp3HW3pQCk0siQJBcZ2tA3P+iC1R2IDiCKGhukO
/2jtfC043Gqukh3WG8qfGOZOEr8R0LfngiJUPtBSLkRM3/EO3hyu3KspeS52hW/ATZCB2qMOwdM4
iEt5GPVZIsUu1Iran8sGSHBdsc7yAwN84bMNG38hDS9LVEjX/xMcSIZBxgyICfQpMHGCa0ETkdmH
pgFQyosKx1cNLobiHmGcFzTEpEJzDjifKQ1GibOpSWJfCAEof8Hw7DbxjEbmuRHD3Gu97R37/cQY
lFZG994F9XuLvQb+HDTrhasO77gwDnVMvHlyGhsCGiMXkr2QXX2mI9HFKjofDdJKRVNB4VWY6Dhm
rECU35jU3pud/pQO6EkFqT/Ap7Y4x46T6OmuwOHat68+jvTnodJS6oBoj1MJtCB+hadA9IbdxQvO
nQuxxy7fP6vwcuY6gV5VB50OZYR5sm1G+Kil2oMyZ69ktCJBYxUQPrDTHAOsw0YRPbfRMn/SiVvm
rp0sVQzIGXOkZ2FYn9OOtp0iEkqLf+O0MYyqfF7T2jjDo39jiTDW/sSDHpfGqVOiTeBemwdq92RW
KmNpzQt1yy+lAum3fHwy4RDVGB+gMQsUyAgQHZTdxVJXpLPCYZt4RIP3MtayibODFOrBwc7iojue
jUji2yZNO84H0/ZseTgL2scTdm/LvYrBjzWqD9jvos7PqrDmUrIPRXAVrQkmhF4DpTwytp1KeMND
qcUOVXOpZlNW/ENhm0329wyMqf26P9nnB8hTqsS33z5kjjPgxY/iCnbZM6iFyJmpsWx2I7QjSJ3E
mvrdAN7ohtvJV7i9mw+6l0H9F5UacrbtkozLAtmxSoZaVlLzb8TlWk+LZu+0TEyMsnud8Kemr+pl
BiUZ/nwqCT2Yo+bqfdgRRmH0zhWITyFS/GjG+7oSupbDUmLwY4hqGd3ShjsjBAkCG4/WeXlDksZe
DccjSdki42Y/vt018LawuMODGibGlTeWx5zT1uqlMG18cVBW+tq+i0afKYOMCMAAywnDC1czc1pl
VKVp9bjn3H9oG8GGPdCZLd71cgjH5BJdLIqSMlX+xCXoGcOXbcfYr+l7y2/KqoOmYpjKiT0zWrzm
eT42DL6qMKZSqjxGlofPlozlxoj0ie4Vk48zPi2+Bfq0BLAe4J6PGt1xd5JoyxZ/OLMCd8Ylqrxb
0zyhdWCcpxLTECp6fK36CLItgSIG1U1Y8M9l1ujN0mURJiJY7t9fVcB3RxSg8inEeWm7eTTVsKDO
0yXlaRp7w42lYX/byj3HYntoBmcA3FD9b5W8asFukeWO5QIY5FJxCamw09RY62ARtVX2VQAOvGYH
kOAYMfa1pE/rX3prDoYS7iANmxeJWO8ENMX2/8xxhKWHNGVNH6f/EaczGGso4xA3OQyouuvdNFXy
Y8pbR3RsrnvAcrytkAjc0eIF9C9zU9gE9yUWtc+lQD69jhW80qifXHkKOoeRaGQ0ihHOhH8fbCUN
dTAeiAMBsv860vudWLFd15NiGuuPl+THIRug3KfM8jFitnOLeLiL5aD/jyk2/hGXBvYK+jXBaxNy
g6JxP7nd7TaZ34szSORNkmgsJU7alzvlt2tgK1sTaTNOOnoGPNGnHsabo/a/AqcY617Fz/3dkobF
Lo41Jil7OTjCXGvV36t0iMYQiIo8vF842s37DdWuvysLHvF0LfVSd9KCEvsT2UDCO0uJM6fWpz/l
7HhrP6ZR4FTTSwBBNBF+hfpV6pTqZnCLJfCCSkdACkwKRYUA4NHI7LpNyeA/hdiN6cJRfQPzHo8b
1sIi9hPk/x4UYJlNt5EL3d6+1kTqHhW9BANhoi1W/Pob18+6EbxvFM5iV8u0DR2tSAbczAhUVIIV
uLMV61pKABGgKED3/Lpae6RDIjdvdhKa6VvLPB/QClFF81vh9WvlkeiCbNSSwGroIJbUlzWRU1iI
S5UPW7V7984u76pTyIhal6BcJunBaK75Z0wd2KQrkd9ZBcG4SHvoWe2QvnSNGst2G/xfpYnF8PCE
yHXdvnmxnbtbNzUI7csyT0Asvora0WApWn1V6bFOpgwb6KQNkV8ENP4WbaoaAR6NY2bc3ZHlPIWO
ZMRIMWhTJ2W7QRTfsG2M34y1W11ciu1R078wApofRwPQL51tCCmpRP0xB4QJL5Uot6E1Cf2scqHC
+R3LmPBtIvEaNiOsFBzWMkMAauIxzvKZgRaCgW+NHgQ75ZYcjnvkUr8NdQvCc/LJIG8bYYohFmgL
9pfniprXcXE615PosjRZ0vrbV2I3SIeNhWSgd8vbMrLyHy6mMWnvg3DpeNdc1Ufr2M7g7D9oUBSh
Vj2Wy2pTpoeEtFfaxxPwcg6RYwvahqD+VUbGHejODyllqnstUWOKXYZt6X50ud8xGVSfNB/OI0Pq
EL6Fe79rnlUxPenkbIF1N1GqRC0YuyPWTYCAQNgdq2NKlEhNNhgNJwMsDlnljwJBmsQ3NRsAvO7O
BLCkYNec9frs5jeo4AceEJGFZ4TZ4+sC3WikVw8v4Zi6BkSi9MWo/HsyTcmnnHdFjyjOwv+v779f
Ue/dmThKa5OunRQisj0WR1K2HkwIR8d4y0catuy9USJ4h963G5N5gHET1dB1zhhxaQxAB02PXdBo
/OaoEefRYsgKK/Ug83uy463cKexiKPFotSU3ZnV/d8zq3+FeZDjjmtuA/vSCP0vhFNS9I7MwSTRS
quPt/gdZY4f0xmSjNc5PhfjGfR03x68DsJ9yi17jLi5f3rOITGWzceRij40XSLLGNRM5DPISdZiV
/7gzdwceIjz98+YEHnHafHl5VOXlw7/3zo0fEFU7F5t3oBBkdwf+B42RQNdt+mlAzr2Mh68Sgn3m
rmM2Ph4CpxqIhNMDhsPcFjEIaxgYpm71DOUOeVaLagxN8aFi+yzvRIknBG1N1gzaPOPEThH29m0Z
SU+a3JmLXqHk9IwjayNCQVfSlXvzusroHZ45m1ymfzzIKOXFLPmlEfn7nm/S+vGjYv/pC74AklTM
M1uFzPqk72gV6Vxs2dQH3KipRnfmYfiZH4rb5Eb22suMtIA9Kd/zE47KSBX5ocnXJaYzlnROl1B8
D3YEnBbzoyoJDOOt8xs4JOlKJxiaBogKyJF51uIYDYijGl+7B1k/o+/A4ZFsV0dFlAg29sCh5Sl1
kD+5iI+PzZXLvD7QWTSAQWs1WOrTI7XUz1bP72mDoJ5J1BSMSATtxmF6octFKo46eMHvlvNwDy4j
M2bEvMxrBjGS10xBGoQYf/HID60uF+SAwu9ym1DBsRZHp3+cPUunq4IlzjGmiX7lCNyfoB/oMqnj
HdwKf+G7O5HmC50bx7INrE+eDhEz2XDsXxwd6iSPX59RWwGqLCBNfEMVcDrzFFgQe38+zcJLMOsi
N8H7DBQJ58aFXlAAhBEAhbYy9FdMwmWrc0y0sZFWPI586hjJsF0bdlRPOhaNw4LgITMNjZj5mn1c
jYZuehqaX6ASdcDAjL9AO/GP+R3XEgAp4kTQfPo2XAFDfq4GQulNOGMkzy+obQpMkWX8nBy9LN1a
LwpQQE4vdqA8fZLNu4UaCjrYKvSYM+MOEzlkbvNsiDuHLAFVD6HhgJZvyRqooI94Q/DdQDp5cWYO
wWFfkoiWxcOX/Ek8ibQL8wDIdR+ZIb1y5PtEUn++N7/SJKDijZVvu3V14duhmEEGWoEUhItJehNF
TaRSlKSb2Vi3x7HJRFXjGzh9jdufVL0ukpEhMrIc7Dp0ZyMAYlcneL6gNomnoXIA2YJyC80/E7ju
1UGdXCX1bCirNMSMAGWzG+pIvbFAdR3XPsV4G6lAjrn/xYn2EcOgw9vMGPARxFRSyeyLj3KP5HEJ
ci56sRzmPOC2KXSxqhMx76FV1DL0ejI2Tmfm5lIKpA/K+MTbBgkJdN/fEEfV+rzn7ym4edSOBFgy
Y75r5IeBCBGlLWdQ86dQ6jZS+xeEGUp+E+YncdSk19nUzhRgqwAdg/7auG+JpZzQw4WOVnTeRu7s
GledltAFx8H+nfakftc5RI56plhUTV321Z6qfCalVoQvo/4x18dmIhpzd4WtTH7dKZeerivcBMvp
04Kh015BxMoZ02cmSLTvYeOQOQChuG8dBwPJpbEcYCbl4CKPvG0+CzrwsArukSc07Ql2aS2gI54p
ggBlDtd8CrhWmQpH7JuesXDbe+u2xUaTptrvjMhZQTchYd3+tgtzSiLeJ0wQmhXQ8WWcN+53hI14
Ln8huEg+e1XIsGFsbcg9eFSKkTL93ur0xtUaUkcrEttZ03whqzGq79bpdpIMtUeqZQWwRwVLh8KG
AJTk0mS+LzckYnax8xaykyUZSHiaNaUoKwcMM3RWaDVRktvjQ+klTmLY6c1BB6BjuO+4J9FeZkHR
1AxzPd1ER87jUpILBpD6BH+TbWUAAFjbaiZgteHzsOqr7t1JgSqz2H+oErYfRDBteYaMdMfBPlBL
7/Ab8ikJZlWyQhzomGSIEBwbfU2DLmVUWO+YMeRowCG4FJBPVb04pRJj99gx1MOUvUO+YROz9DEH
AoJmf6HcXFV2nh3eEVQBf4jhD9f//SrCLHFBTgxDByqEqkvGsTu/c2dP7JTczQpTK3CKlBWMll0k
ZjjZyHQlNnTCCTECDiyNuJK+WqwIBodh7yHNNWc/dVagnotlqwyy2VyZLfOKYyOPdC5lczhHnjOV
Y2KA2oms4L3Zmu896rWz11GHaQu8WVrMnF6LxlZTrMIDW3QiTQ2yAbNZhkgV7DGP3B4V7fUSO7zY
J4YrPBanh+PuTa2FuzFpv1KPhgj6niMs4NPrbEmmAIjGmPOWuRzWLV2mF1ncOrjeS8nmgj5UVUgZ
aU/K0jjrSBPufLBs89i3BEFOg8z6I15KaaxC/A7YDysoCRZxMqY3mN7jujy/GMvpKzEf4s7p2sjO
dX62TfeCmsXt8ZWBOI/vf973Yy+xpLjDeOsgEtxNDQiy7JNLqTT8oY3VKpBknyOuwa9QXkFi4Vjm
3pnAucjzyibMGLj7z/wpm8aXOBzyM0+6xwAbziF/Ygmp8gbf9s8VCCurPkjvJhhHJD7fdTNh+sV1
KpioGFD/H5E1usymESCIBHDrLYosQin73dlwtTpH5yrrHskqCQKm7ed594bb/2mcDxTyCUkRJjf1
4BDKH3DPvXZqIScjYQ8g7PPivzPeuVyTD8nHgD9tr0Kcclnbiz07YQRxse8zXswAM+A9n9MjVh68
5iospsXb42bSFKqYO884rOiBSy0gI8v8shLXLtkyDBD4tkPUtS6ru3sqtDR/OM3C5v7HxByf3uCm
YalMehdIbcvFaTdYZNbZS2/5nn+efApGRSbECpeC5rTvDKkqcocGrGW/+bt7+kWNLlEq2bBQsexK
MUKZianZMYXI45HriZYiUCWqgleHx9ZhavnStaFp1255oIVFrWuHNMwH4iIbFSvkyOkdramWl4sG
eKHQrBMt6hUWnmH8MI22oRKYAjgNEZ3OMPOYbJhDbNOA37FW0Kpv0gXqhXxwTyEYG2vbkohWzTIM
t1LN7pbiWoUCMNbWxXVub50EgCWez27lTMwKVFIJpFSgBlF0/J8SFJQUtsrJf/5qm9+0/3r0ZFo+
dHQvA74Pfy4BeP5eWoRpgvAG4EDWF+Lv+RKJuIxrGKhJL6Dy5TMiM+GefTrgxF/BcAq47igb2bqd
MZUyJYL7LsUn0jI5NtWl1h2UWLpWN3vGmwsSiuCWlJWl8yg5rbNRUNvNJE8074R80tjPZBcroTdf
YlY9NuR9njhlPWpxIuyrv84hRaLHwNH/akfScG+nytnwAsisSITdUtz/JwQ1LYPDzZ5bo8qeMLZL
Go6wKldXJhbVrnnd97A01tM4/K01CsBJGYAEzo9kdmb0q9pd7OUj6IkLey9pQuJL1qLHc+BLAHAK
BKSJqlnkXdqkujRjNqKlWoI+77IrWSQxvRH0CWgB3PWfL1bEKSXwhXpgnRosg4U/aQ073MoHfuQo
B8d6DKZ5zuPG6pm13VrQvGVq4Vp2+wLNXrGct6N7Oj9+9+fG+ddanL5hNESUXJ72XJGoOE4WS+vE
XS920X0toGfQ5+eWEKo/1W7iow5ej3kuSvI9q6I/kH0j62yy6LnDHSj9nyk1nmJX+SH7zl3t4aLf
Ufc7MT9htvkn3j+I+p+bKOaK7wQWy2JkJtv6Hz8N7egFGbl1WnCTtxPE3V4InVNerRUuWqdk/Dnb
qV7Gc/sN0FmophskVkzwkiJgziY8+RFAJzFQzmXNt1TfpjbW7Fn9ucCcS04ez0oKCjCLg+gaTJ6v
ZVHwTnddgmI97Oyn/pbwDmpT4FdPkORPsy3JAT7ys7jI5z8MaxiG4zuGwzfHXwD5G9gHXKEVQdNS
scbA6OogkDnflvhZB8z7K+EawS4VhXCVlQ7aRgw1yVtKy4370+xsA4yLkA0gRrMmTTmIBocva/q9
LoC/DpS3WOc6aN24cvOBnGS4sZSfBbOQyeHGPHECz9NACmUQOvz2mz78PKVGQq7ndnJEu71Q+GUA
i8HkZEtoZs45tCwAeWZFDnbLS31IxSCwobwhbEurTtTXWeHG1jms5O/0CQT0SpDha7Q5fPZlouPi
XQqGnKdhwjKK2HADPmT6kfa8ZhoEuQ4AFxFBnEyGdlaWRZQbheyNB/NCDPSP5D1pOmdD8KG5ooY5
ryOAkBO1FLLyYQ3emlk5LbesstuCkGurPMMJUNCdX1Zr3GkikmtrxVumKf07dosdfYsi/hXJ8iaL
ZmKTPr2HWXqaWCkBhQ9kkHteKIJ9mht7or7LzF1SoC6Ntsef2zi8oHKTzBjeX5VjgGMHjfN+f9kX
VisdW8ofxJCaN+AF6TlBwMJIzFIkyaact19FvFtGNVyC4+EwkagNuEipTFyQ/i6zhk59qdn6BWdx
SrwrWi132TV2RyxX4CiOYzZX3yIASY5dXnYQhNFoeGDPK38TtawXGES62rDQweUOHjTAnbC7UiWB
MUTK1iCXYvsQ1Rw1C4fOe/f0NTUnQO52U0PnoeSTPA5a+leKkG5PYGvc9/oppmV19EywGc/Pts+E
NZHVyqgitAgrAN0EGjFXedFGfuZobWHXcmPNT9SK/AwAGx7KdXF6DurPDWKb8+aoxgVbuZrKLjsu
Ey9mY9yNqZpVZHa5pXtnI7mG7GcpUPKn1L8WvTV/wulq3NB2kRNOW9+7Raz/gAtHuBHlxEV/1kH7
hi2AKEtEriwypVjYRTSBxeInCinhks/Mxf6pFih5SOphgMO00amSEMiO4vUbFVcybZyPSkIit+Oj
8IQMuF2DpMnD1k164aALqrTgu1bygQr7SGny6YV9aKOCb9HWXyY1aoukG7aurdYSrRT53GTF1Git
ysqgDf38R2e9b+SW4+sZG7Pxzuet1e7sL5eyL7JzqMi3cfQl/FNewV6PcfhRy1a8CVb2pFF29sMs
IiNqs0+uBLlVz6NSrmP9+INLymxuKD0sc4tZ2yPaJaENAFOgAwyyV1iGJ3qG1dt2FPra2aE3Y3QI
Yl7d8Al3HUzpzcqR3u9DBNPtBShglX0qmjjGAxSv2L/u1L1ULKH0Tsb2mBXXgSvTPQFaDtc9Rp0e
FiXH+IcUP68LCEcqT0gPtb4c8hgUJS5gPrplrCYktsJ0aW3jfsP4xBy4UyJa9WgiVlzD+GF+4T3Z
BO5YZ40xOTV9PItPk+ztqmep5r5vib9/Ry2LAaSNY2VIIBAdEXR9MOaTxg2KrcrbzCVEE97OC1KD
BiZtqCtoM6qnUpqoBOy5p1VErRB2hoZ6LWLP1jPs9nwnDyDq/VJmsqwVXnGtJDgQrWWT3frt1jRi
5yaKq2AZhtDcpe919iIYrDyisVow9WYcPhV98EWXJAKn5g4SmqotjVDKbBEzmzbHjA7czfqe8u0v
GelodmxF5BhHBlR0WgjvAnukD/kFr66L5GT9OgF5AN9uHDujQjzssWfWDrpwpqsRek1zBIQsa/B2
QxLNHZEfJymZhXQqQHIAPddiFAx03nH5b1m0S3ubXKyQr+VLNyUV97+CzxrtphEnXb/Sf4YmSCM8
WSj9386RN5wj8zEaSKcTcOVUMhKuXj9N8cKR9bxzjXx/USUSmYsRw3JWAjBhujQ8GYZldQOn1CEz
3rCc1z2sfb8bMCxB/eF227GKHqpyg3kjLZ+STMRTeo2FjPOdnlZC7dOSjpNM5axJKPW40jSgMHoO
pisSR12b7T68EE5LLyp34qMMxBS5FMyEgo3B+e09T1wQSXxaZFUXBAg/wuK2iPhl0Tg3ehZ0bL/T
dSgwxbJ/KnAAApQ342OYxtDGEvGxPlp0H62oOTwxvidErPznAQMPnMq9NUbcLM10pGU6wJ0QR195
U8haKjW4Opqgtty9GsuKXPMBsu9qIsYcPemHjsNT9H85SXGoQ+skO6wy7EO+trsMThqVxdC2mC5O
jzT3u0PQtdGYuLkPqDbvXbf2EP78YwX29BDU2qnXuXjO4i2aGO0oof84+XAkURnt1zb9PWqEix/h
daJAgtw11/QbGssf6h4lEOE1C1C+VsE6dPHiljX9pfFUMSlx+LeZ8pU0zBnUbJLzmsfrrKaZRc8K
Uo9cnYsv3GNt7ebdoIS7SKCWR1CGkKYiYwqzMEIRl43kgfHDh1LxSiMMCpQ4k5uLRDJ3MghsTM7V
VW0IlgoUwCJm+SCrw2uXCA7xvLlBXmWANAmgOhNzOhUeIQRHMB9XMP+x7+CUHcYRi2JOInSA/uBp
ied4N6AGoqyUAAQcEogAVxT00h4oUeJxNR+h36y0nYGBhZaD0n6LVAQdDVQGIVpPbSk2ri+JU/RO
44OEG1khRkpo43k9WRgHBasSFtor+zCpX2bMOmArhCLT14TYzUEV9pn+tgirMcq55lR/M/t4znuX
/K+i/ehTGVqn5nxXVbOcN5w5+L3zfy4jZ3pQcA0CAGVgqRhfVm9Bz8uri8bkJRLdP2eWv4nVkTV6
PFoNRjpK/yQ8xufOU9K2JnOxgcxrqAyICFVk1XeKzAOhNIeKArqaaDnNArYMCT5joRxuvFeDSmbb
NbbcE3zaJig70Y/TV6XvlralQBzevadfzK6YkEy0YaLMwN/z3XWJef2iddt53pY+2ZRcD6ihepbR
Iy8jDB5+T8IHUruThL2c2QtTRWNs1aP4nsJiNUmWhZOTFZ1azBmuRYYZiO30dL9qHdMUd0FoANjG
8DDCU3XvtDWK0sE8eeO04w43N3n1h9fMyf86j7BSxcLsWzDdbka4O9ONm54SuE6SM17phmWPIS8i
PU3njJgl+dafXXAUS/Zm8paW/Pvx3G+vhLRygaIoSW8ren3zy5JBmXfTrMy6mlWf/802r5pyL3R7
0Q7nOsXeONB0UZXGKCgu+OeR5qjGPy+ciMh0NxT1HzzrGlSN4RU8R4StuAb70tMqCY4t+RfUb0hx
xmixD/Igo5KvQk9l3tVCfuPlhrT6fDfCp2mp7/bjGeIkxeWFVYvLI8DaPQiWAl/l+6K08ZHF4jCW
d+iVvZImoKTCjg367uQCKNICHjuqKjBM4xnkVbQt+AAfPA3bpavyb39bMDhcr9kO5rQAQRVjFAK2
ZKqJYAI/CPhCGE4I2q0F/IxG7UbUwU1MoU+bLXtlKMUMALOd4xp8Sdru4X8f8xHO6vHzYIzLuK81
8fFw8gNGyUIViKSfaCMO2nLp0l+KL23N7GnHdWBooJqnMh/+OE8JdgRXkDkqCvot8Iy1WIbujU3H
s21AwiZaS+1aaDMYV7WtAuGSRkNeZVj2ZOtYxP5+cOvifI3kPA9umGpFT7Te/yV7mHQye3cqgaYl
+8BUNfTUbSDLv8i8lCuhdiOs4nK3DZBQ6LcTcqq2E9eVRkIFYyc23mzulP+Q9HOQUypiF4+SKR/1
1iLBKwVCXbgFVRy7NTcUOLfZnEqP24pE3274A9noKlJIjunbgwy/9c4WByZHNeMvcS9ncIPfWD6O
OFBYERyXm/ps3IZYl4mVmgkA9MhJEJCc2QaF20q614J2lZ+An4hYoFwXjyKa9VADOCQJpuBtWnsD
ZREJ4pKqs+R4Dc/Eoa6oKsLunmXf/Lb5ieLwcgHPjB5KjF0PeNbmavZPa+QDwLU9qNFLH0cvaWRv
nVrALESffb44jyCcimxg76pYA3Pz6xdNcFwJDpYmffF20vQs4N5ELE0eLG8oIGgBMd9h6obUeo8V
hOHWPpsVyIHRlwniITqx0BRDzd85pEx5XlKYUbsiexzor6ySLiXTeNAu6MM2bq2R8QlJpWAQlpai
Jm5Rp3+hYefnpwFgP3ZCng4QOMoko+MCVtg1WHhzNlsMmr1ORPEH+MEzjogSbhREPnZ7MUzYlDFo
tNFYbmo3WzEexIx/j5onlnigrQYZn0bNMd8p2CH1/mcYKozqvgWRXgwzI1w93J8Hu59os/qwhZq2
p1MMxpBYDcQOpnSIq2QYR++0pFYTekAOM/FkkN0qisFJ9MgFyK7USWRpy2vHs5X3nEGQ/TqF4FlS
bhH/qTjvOFUldPu8pfPwHyZaoUPsUFFGW00OCP8iag+MLEdCSTZb2bAQ5ihp/0jwmWm64/N4ShWx
yYhPPo+LGtrwHSUGVdZ9FZFNDDCazQNV4bQ2ljPqPJcnQ8UQwdkTZaPpXtAgX/+Xu5oCq7z+1Hhy
zmxem9XjQA1ZtEa9vrUL1pUtFlT+x4uJs83Y60VdZgzShka/IoxXihSXykS7dtH80QqE1izCirqF
SUqAYMxvFTNIUwx427IMKq68jdy9H4g8XTm+9FSu1TPifZmT7GhVad10m50vulsgXXR9e3xEhs1k
w+9yKy4jtfz+/of3NxlAkJSfJBsx9+VD9acN9eIGxGt0sFV6FgORmGD11iUqm5pylCrUKUla5Gwt
G5u9BmtXJr6JjUJdG8pwLAD+XJFxMNI89dQy57sU9Pa1b446R+FZNmvYz8FllHKoBhkz5xzqIn0T
DmPVzynHRZFMLY6it80Mnnf5ijZoZucxJK6ETlu42yz3wkvWae3XIlJaJkX1yk69C7Q9wEzif9il
f7QRTfwWeVyrmkjeYN8POO+YPaJF5x4oHef4fMmTX/TEO94P17UzsID17agT/r1BTsz1PbDFf7Xo
l+y+oPZAvPikM9DtW4rsz9UOag6hWEO5cs7Df/M1/I0Q09Ce8AYRQlv5T9iQ1cbYv4xIiPLAT83a
+DS+vvZyhlmYTuwnqDYho/HH7PBCYmKKbX9tl/zSodsO8f/v8Iih226sxIOu9aCYSi3tbGIxptBL
QIOyUkDeLs/j4fbfnXSlFkcul/0Rfs8QYHvfURwAOcLIXeTeBHGkKGEznvduAI+SxCBrwI1UT/xN
sMzqV8/jN4VJhAT4Hi0Fn0OBJaDEKtaZeE7hMw+XjhDIoEz09ZSFbc5zm2ywL37idJTrmNqJZZLI
mSAZ0+FcNciaeVjsyPRlZmIe5MFkGSxaFXv284KbozWjEMutTB/2+0LpA6W6+lPQxhc72rDVNpUw
oanWW2SpvVq/d9k8RcpEH2ZA1vUFJXToAZj/JoaRvKvBfkZ9k2dLr/NVeKYqMNeN2IcKnYG+wo+B
PNBkrSvdddPRJfho4MNfjRNj33EQH+QGtqUXiqwqBkl15ZRd3w+Ic1vCyRDRHTRiOsTCSYx+Fxg+
RNWlN9C1u3SogrwEQLOeC2JDI4tCis0+oMktCor6gBGR0jddagzyLyb0aUuxqO3mKiRHQXKkFRbi
lzEPS6PrJXrWiLqBpb5qLo4NVgddVPMPrAD7TayER6DeFg1CtZwXA1R9DkYq9qrvWER4fWpVNK9a
QCaFa5532YCGLaqsiA2SXpGEjB7rDtWSKScJqFfRcuzjPe4E3rbP/6UsqsXQem7oNwmNZyc67MHF
amKGGF2AzCP7zjA1ODww4ZyH4PbPEEJo7kglLfH8nVMPYRMi33N73blzOYbkUkjuylJxCCAPbU3+
dad79e4g0VAuEJvOEmxM5Y88myekEiq/hXtxCoJxnZBNkFinhr8/oRZxiwJntxH8R5vT5o9syd7c
jqc0LFTpXkclys222wmkdOLKeY0IlBTQ4gaBo128IjN0YGjWFzAXKohzASlOQPO9rylx1w4I3ydp
KQ4MnI7itabVlrjzyR8r2MmF6TaDzi1+kUgNPspuiM9JAmyEkCl2f5F0D8U5tN8TdMhe8ghTczge
PJDmO0xUSrRqqGPc9d09KsY/9LfZggGtFveIuS9ouUEGdbRi/lyEQ2fLlDtXITCcbK5WyeATT3Hn
9aOOsv/VUNYWFaTeAZekX7TTuSAe7bc/9tpoWMGEFCGzK+xYrcgphylv12GEgIMyZRwQftDvLP9y
xr8E93JXvMfcNEVT6ZIi9q4sgJwpFqHPsN0064BekmgQZxKyepbBHebt/0h0aAG2wfFoQ3RQLdAx
22FAVUAffvUNAiEgvr4A34OtCvu2WglL6hkLjInT9zMzsffdfVpoRtGrrgY0um9dG3VohSsMvDqt
1lZLJ03F1Dv0Fte77iSyIOa0rRQbZMDaYCABesFUAKwdNYdr7K8rull+o6JMX/FMQPE4h5HRVWEm
OAGetw5ThAGeALppa6rPYVYJZ1Vej+DqAaaHtgNMBlIt/WMJ6919xJfPFCeSuBMthGmqE5MIBXIZ
unPle42seCQtDw1ABmLHNKQkWDjPxa6MXHAGKQ/6H9w+KxpTmp3t9IIPI/nFMENSm04YqI8D1QoZ
xBXnQaD/7UmZJ5OdyajOHhpDCPwI4wzouTWZ3NZcTSVno1MSf9rh1mnJrhV78yc7r9CCmcxIXZrZ
nMUvandhMRI0viNSAp/39rGkbByDadXNCHdtd//kFM2YtlyQ4QEfhFBzroSPB3+FQqPSyJezmMUO
VH9vot2Vi7Hgavt++dM/iYv8ro95hZRwiFqKMCr0yLbOj/FksOn94Yls+A5Nj5ATouXMEY3OkmPT
rDbICLSbkdsruPutHpDaPNYHYB45n1eILCMs1wDi+5fr5RZp6nlx5VF1i9Vvj0Ubx2Qrd7z1rxgj
Iv/+UcaLxBDICqUeQ8MbP24xNsF3jU6jm4KwE9uzNCxeihjlvAt/rIX8Q4/hGIhvCJW4qWnK5c1g
61x8fyd7Jqyygv9gVjhKTuSYkwMNlytjtxpGc/eC2OTXP/qCY3Y/GxuB+9gdB6EyvRggBt9JFMnE
siFI4dYUjIg/qmW6XBvVm0Ibx/OlrvAOuobCsT+JkndbsU+Gn/6ZkNgcQk90UtIIZa2rCU0SZyNT
C0KvT9pp9e1DxXVnLtzt0ZcQyvcyGhMMcbf/9UMFa4eeGsVqbYtxTmwmBAoR1Pot5qlPG+Ix8jSd
PmGzRheN6nk/e7hn/+Rr+Eowdj2IPb0OI7rKDSB2pSxkqfcj+nnDA9fsrIG6aFDkYYwjeBreY2Tf
CrTvc4gekA5Ordlv/y5SIzeUb6xDsNKTZaF8Qwb85crNGkWJE/pKJBXJVKTVwvinmruLWwpgRiLy
5u+UEQ/W9Vu82tVLasIEO3gEMFr+vF8vhLPNofgYa/D2hi6e04mmfPxbi4G+h7dGRQWF575nTi5x
LMv15nMWygLqHfNztE3orfFkCI3KK8+udWLBKA4y8u9ELZOkLI+kygFda5wXnvqlcmMeGD9B5+rw
8lRfa1qeTSuRky0nNy81p4NGxTKG06tQPcv7dSU2V7fpiR80oqyhwjFXHPKhzOJTDdihryx7oDSv
WhB6reqOYyW/dopy/A83YW26mxY3gdOGlKJbYANOT9OS4pZKdYIseJhcojaVf/EFnO5iFcFUHwVL
6YPJCJOLmgvIwB9JEZX58EN+e0o7C46pijj0L5mv14kjB6XZHLys5Fh2wFk6BSL2NDy5T036mAAH
9EamOXSpPUGkTTryB0eUXgcmyp7nQjpmd5cDtUR+1TXWIqLK8mgAs+jjodq6tue6jG6WpOdko4BF
tn2Qsl3oXIEkPGVjvLRTNYLdE8Q6MGiio8ZTfmcJBkctK0GV+eJNMeInCFezaGbXulg+4SI1SseB
jhlilgSPEhffCpVdoMYWTbtrvINEWlH0YSdhsvPBcvl3C3aJtG9HaGM43RREnDdiqKnnK4mQ+CjS
wyJlaTnl8HmZd2Qj+iYXBb8/7QPdaA8CyJ0ziuvswDT5Bs8zNq2OAzcmvgpg1Lbpic+x++Wb6MYX
4I4fFwWxSn3p7Rjly7Pn95xxfoF/MqRXk0HHZk9bhRtkIUzr2rlmDFhOndAuulRpZiXoJKGfQG2Y
CHj26BX7+0WvPgE5NUujUa+WcpBbS9YbMwtHWtq8oOBjMOarhZ+6vmxe9iln0ydp5NEbiPD9sQrL
BQdZQK+sOtdWo24nHwFkrxAMtqx7wZ/AQn03LOKJWDrurriEGyT2qJiPf045d4txpyM66l+1f5G+
TDW3s1cuH9gwMzttMF7G2NYnvaYK/XIWGT38GlU3bkIZfJY0GEzoYB64+wPEzbsUjs4H8OJDUwoE
u31Znd1jqBPXzre5rVCqzx1ATtK8mbAea4UOYBQf9AyAB/sWufHfCyd654erQWs88ztJgt13O0xK
3K4P1N3KXteBzX7l/IE/+87hvM0xXQoH/sAujM0cA2C9zFoEA4zjTM8I0aYCYDz46isBAi7C6nHi
BmzHIw2+OtfOaOWRz8cDk+AoSJYXlHUoXnPirVQlQNjemwQ7MV0Ox8CZ2MXhZ53OTmxYnqAXTO/B
XOjWhmzzxJ6ArZzzWNvMHOjACqwvybD5qefWLCuzdhVTK9/mKH1YuNHMrijPjmRbmBy9JaBGg59s
a0NvJqaGsRZzbCtExlltMaNRPOi+XYme0HgPYluJt3TWBOPRze+uwz7KA0Nefc4Ht/m1gDxPdqmA
yBEA+mMVGyOc+L2BXIolMdh5eYVRapSUJ7KopbDGh/67MvDW0yAztpXft/21CQ09z80HCagSXpdz
9FxqhMHJiX1VZZg28/2ehTr4ZZyOzZpFZqh7QbrKqsHonTOMcRYnCGwrNzWjdAF45o9fKMFCPKzX
4l9liPz2gO4d7WuW6Jb+yccdSGM3O8Nk4uRdr4OKoNGpAO4t00vkPFmcPi7QcKZcWqaxnE9EcVZT
gIX8LF2LfZ60AsUiBypC2vKh5oxdp5L1ypGU1Y3A1S2l8wOKW8LwQR5j3+S6UaqA8uFLVW2m/qV1
rVMlh7630nbY2WhzhWTR+lqCMDdpXjLBbPD58puCuxrU3lGcr+V7B+Big/JmuhJEGASGXBoIYEIm
aajWfEMC3FpG7dM0c6O9UrYb4/fIbaewcB+gB+Y/4rxQP3uyTVQlImnqoA+jjmvjcvYlLDELFSFk
prFaOFJydmnBBuNd5fUR7LJLC2pRbV/5sHzGXPh2pZMytJPF5LVqX+QhS6zq9Fw+LAuSBgP8W3XI
0bqOjTMF8XqEpqM7JnQNUBciur6AyauYVJHxD+MRh41Zn2v3FBEPoqRIQ1fG9x9hLMkDwd5+7cDi
+hbTWfpmF6MfdughJ0Bo1j8ujk7xyGlb3wFartnVgyyWaibCOloueqTaFlgWxUJuoY6RgZwKznls
3D0Ggz/6HnJx9SPLR+bXNZY+D1Fst/U30wlkFFU94EEapTbFLVOh/KRu+/wGqe4hT+LWpppCIE/E
NJIFmoZ37Aqf4Yxjh0qkFsoqsgd4K1GdhID0F/Bq7IOP5c2+5Xa0jGAnxL/40A5ENlUPa6UouJ2N
6EHPLMXkjbc/8C9DTRuVfCF8fxLliKMMGuqLW0kdEWHjmweFUjGboocn2KdVb+HMkmjrNqnGe0hI
sFH7M5oApw/dbha+D5x0sBr7nDtNJSqKKHvqFUj1NOvnuh5DeU2JksPUuF5WVLMGfLemOTDusGZh
lh5B+zpgQD8bbAfKyNpVP4h5eEKDG4L7nyVtsVk8TTPrXD0pySBksMQva2mJ4PNnssckniNrRmdf
ZBqD62aEczlxt09fmhDNm7RIKrrO5R5FOiWkpy+LN2hTeAkYNx5YNnROKB38z+8/2hYl9PnW6BlS
tnYfENP04CGc+QW9yES87j3NSsOCenXYPdVMYxhR7UDFFcT1M53f/g3QUkb/3QkbQEYFJ+kaW6B2
fQ3N0rm+4zLzJP4AadkNSKRiQUY0R11cDh17P+4kK7AhaXqGWbbM13kXHeO2RRuW+swpXjFj29dD
R0ZHA6iO3+4sEBiNbOw0AXVrqVpn8QnH2OmsaJ4GQDEuvtZZ61Km+JuDD9vMgappyGr9XbWBAMRd
NS+9Dflolp4lxRxk2sWy/Zjrw/cthkew/whN9uurF3wUcevAadsokNcyy4OM/YBjbVBI3OE1IeW7
uNSER6KKw1vjEjvSW0dBgg3+oQSBQQvNYAKt1O/b3VpeOM/24drZgKUzEHhsaWiJoFH5440zkcFl
xhS8Dgy7jwNK7Kpc6a6i6BaBhuu3g3W+Huh+6ijEVs9IrNXzAE93aRJP0F3Z9838WstZL6drHbQx
vm11DCpNbyNv5DnPQWUSMkleUHgm3QIhzgfxAe9WzucxESjffLUDGCI2RmzGBya2hI0EcIwzI8/X
WLM9q390nb0XHhxklucwQltkFrDmPYYQer7dQ9+BdrK5lySA1svwP16UxK2hcgFjqm4KI/KTT0bV
Yb0RcH0AN3cth5FrIb69udKh4/yTT93tnqJWLHQdO5AMREaeOuVowPM6/lpdJCcsXVr8wcLcOntg
qZtH5Lml2EbEIhTVem84rDUVyrcZ/zv4WrBkyKLsZw7+5sD0Qm7018bFRTGjG/aH97gTSof3/0GC
AU4vJ4kcKg5HD20YZWpvfY4R2041otzRbraFxqNjwNLU7p3WrErjtuKpbDGdyiN9MNYBye0mkSJH
jl5PaCb24f3QqtiXkn4RhkTMozqmpLyp/yNlldIw4jH0xy06DVRd/VoD4VKdXi9fQyjoQZNMnc5L
okcbic4DMtDuVmAszcveQfDkxsojE/JX2rj6m5iSUqFyotJSZrAdoQHxhnmsnsUf4qM2/FgGORPv
N/+r0vEinPGOtcUcy38j5oXk4qeMpSLsoHtu1KGz6RK5P0+hs4hU1v7IEIeAX/MbXl2TkbSgK1Cz
MVEU284bSo8EUvKdOcmupI649ky91DtOvqDD+jvbhQQOF/DLSvHNTz6Xf1W2AthRt03UIFObNFH4
xtg1K9uBvjJjp+k/gqN8nShZwgO0X0IzUWlBuov9Psu7aGk1DVlD5kFil50ErtZHdhRP3RjkT5ki
yW7zDCcP8E2uvk4r4Cxea4MiYxVF9+S7rzyoeoeXVELyeVEjscXAMoSFnn1wCgrisFFWF7IuZt9R
LdnTlCcIUUctP8vDFFE8J/5B2hldGOZPTv21qcU85ktuXXGflLaE2Q4+YFvGFyOpcOHxKfZ+qF1E
UN5Tw7WZGBDT35wxasv7NIE1zXqgMtMilSK9i3y2pL6LAU31mMdSVCXsPrvz6tvcOBmhX8LO7s8G
t5RO9Z7F667I7GHLreB9Y3yE+CD2AnAozMPaj2zFvSL13uv4YAQDs/i2LxU+BGwctWmLZDeMd6Oo
pnEIX1PEhuY5wZJs2fIZZHNgNV+0j6g35ejq9YG7VUc0vS+MIWtRB5MeLEkn8oVZvfunfGp+EH4z
2f/LwCt6WqlNhl2BdmDTve+k1C7589ciBWNrulAqN/s1VC29tkcUQ4jutJx/+M0PUgFUt2p+k7ea
F+TSfYkmE1zFeu+KJ8WOHxLPLRqEvB2Lj69FnZevDXzgRqokGXBGaeXy8MMF4HwBebXaEoQu8Lpz
y8QGbh0mzkUWz8zIPWmZKLbUPkuJSQaCBLBhM3SnsaSgDwojw+V9O4D24lhBV27iQCn0+0kV2+xR
19eubQ0tHrLY+MyQHSUn8cniDZColu36ahFGI6iuyfB/z96cJChQzrweUXZkXU9/gNX6TMB3N9Zv
ta0C26Yhc/5xUlBChan+KWbaPa0Y2+/+QaZEczpVmspcARaLy6uVmDVU0GyJFZvy01ff6TsnRVfY
8DEIOUG5gFsUb0UuoGsat8wUZmEQT3QKcryWb7U0rqudMkoD2ZCH3C6M6Jd0XcjMVIs/fnNxKuPG
BfFpW6Ps7SK7JzhgA2PjCvVPUUsQsaI3YCXgVDo+h+MOxC5BB31FP6sYFtKhFtNEBeeUh61T5CyE
OICfnUTPTkBhTf71XjgCdQvaio+knnT5hQQitTe/9eGHYmlDsKlvX/1Lo3gST4EktmYblM7B+DLy
QHeGNEi/RMzK0HD/sDG6D+bLmuaQPogynTy3WOBtsYdLyKJvuqplqmHYim9YMD59rM6haixttFFZ
0pEnVtVMNQS+iYh9VnhQxrnu4MhK4m7jSvEdYYfsXoiCnbtJIIEXTsYXeiXCFR/maZWI0tz4jLtJ
fdGctBh4zj9KMRU2weSephM3DhIGgGrfVDhNdF+q1fJQm/Y5SyC7G+7Cjog7lCc05tmBW0nXbyh7
FbKSSliBZleHsZ7mY4IA4hg9nGF3+tSdkLkddfPsE7ChZGHeQibO1zEo6XRhsoBRDA2AgG/fvTuD
McMZzdHiFbru/g+lGC3BgrFyfvkLupqfZaOjsxtohPY+kMZ6DZ8G7/H/0Nw+PYz7z2fg9Mz8nCnR
gBCPSMIfaLko/bgdIIMvDMkvwNQvt/HWnkdpa81nMLeQF0TNFaG9sADVmgHtiUU1xGFJ2tcNDLxz
EEnuHTSRKCTk69XsK8GL1F9vMVQY5oYyrc6aX6QYhALQMC9LmL5akxSsBhi02GBl+gt5RkZHUSEy
7y0n+833jepRki6xnYLmorpaVIWnNM63XxeiDSyEKuKN96b4EQB45UXNKaXbv6OCV3ITIXbrJUtk
Dxnj4yr9/y4G+fxg3rKr4KlHZDQxUfb3pXHXF9hHOl01um8yj8HNXyHUGgbl7z8zYyKspRwVTOZr
D2syTT73vqh02FcsPiki8Ywo1T5EHCGo1/4Jjl8XPbCvdVVEhPwjtVoTpVIzQwW2vxL3mcFasnfd
4ZG0Mww3xuSfrafSA3v6EWGnxMABs4P6f5ZhEeG+rJHZFN/SQDgReY/wksTM33gEdk7fBSlG8Kfh
v6LZsq3p/2QrH1WeIW7qQIQf9z91iU0Y577Hdwz8UMW4yzwKARfH7BvMRvlM4RQzZ7c+Dq0NHu6S
GFaQtDOgXr715JvwAfV/v6j2ZMK+RX/LW7gIqbt1TvTNsUi4mD6OY7cBKMtgdo0Ug82HamIVWloU
/KahrI+W8QVnJioF/S72aGmVBI4r8iTKT1QHxwebVV114uIeI9nWmwOc/C1X2sal57DHIlZEWPwB
3n4C4/FO9+WvxNkj1YeB0cgjvF6ODtiqYk6PIiDydNjffZr+mfz+O2NiJWPxYOZpP5rzkLoE/fN9
/Z+P4LmUSUiyCgWyL/b1HkE0yRnNHL6Z5bLR9g0MCrklU/yOCfjRNeKzgah4c+75TmiiHbwAEDoo
DQUsobtEU4ZWzOPcvxaoLXBSpxTSV8O/raWMiZ4sgEAwuDvKAbeoCSVnbKd0LnH555IsBhakFV1d
16aQR4j9vrEc2sDqzh9ounbBTOZGKLiZBKNEr8BNlzEkS8SAD9PJdxlj3mi4JM8/VhU1SK8fXkcb
t0Umb4DCe31ZI/isknfwMZPwwcnBjb1Wj1NSDX7SHDQ1Og8DRsu6vfsCQceK1jK5SvjFwC5mnE74
idfYAFgXUR6FEU4Qdx0Bl9dCnS6SwXJpNUP+BxJo3wRTKETa1J4b8yiDCmAVbBQFlq8CbmALDAtq
tya6tGfhDux1YcQO8tWba6Z90zk0HVqCyWfkQz7JLdVi3wNH5UN8SQ1zN6Nd0TpF4KmJyrj10An5
aoEl/SpLGJwhFgl7t0Tq1EOqGdo4ghcrpfqpl/ZWoGK9J5fwxuIxa+A0x4PSPXu1Fq0/KAU6vrvt
RSwY8vjMWHNeBRoDYGCK3ZxPGLga82ZVAcN7u3MNAwIRU9dEXJC25lsJp+Ymg+AKOA0F2u7jccs6
6gdRoGWHS2BqP7K+uiTTTXhbeloja0SoVyGS2BHRtcKLeokNN4uCKZDAkENvIxWstqLf+AweFp0h
t/1+9YiW9kI0nTrg8F39CEGSPvO3HoVQnEYH9xJ1dR2b6kDyUZPTeEu675AjdF9IuOwQ1bImkCzG
/6yDQ0ffNroE95Me9hjZ/w3SNQeK63lcBk/DY7OdDL3gHp4uOG3m37mHrh7zOAEQnXyranY5lGTb
qjm9lh4eFXG+N7ofTuJs3aYDHsorLdF2ERPUXj76YEcU18FZsr9W8pUQ87BET1fp5SBu8OavkK/H
XmrP4chyG2O3jj8nPtYGB3P8StkxRJjDn639BR3It+z4AofO1H0dLZg1wwcZFUlAtPyp0rH0eEQ0
HiEkGd3YBsJzQsaUKAhxAD86QiRpRajrIE2JiF8Bs3y2yFnEdfOfPFykS5F/XM678RoYT3tSoBts
qXYEKM2jHg6NZprv/z/nMwgBa2wqpQVnrm6n2s71lzJc9YXkWeLjx9rNjt+NzJPfdSvYEMSRHXHK
63Rqn+659uzAmL8rt59WWKAng1R7CWccb+REO+MQnWs2ze2dpXWlm7/C5bCWi1Aa5LjwRUJxHb5i
NYQn2n2CT+KeHtZms26KNfQxMUW6GYjJUhQJEw/fOAUjFW9dDVuafdAaYFTlps7s/jV3QpAAgS2G
+4kiyxWWZOCOtQfi38xt60Punx+Cc0P/rGp2pJJiZO2HowVzSJOPUn7iu1mUyA0i+tU/UTTtzavR
8uNLFX0PO7BCvDI03pDrpKF6yYO9UD2hGBEKPgQnbDvQ8bpwqw/2N3tCy31LWy4uk+VstU07gFJG
uiXOhUgob/VZRDnx8PddaYjfjoseKVamWv4w3PfaaJfKR1hOZsu3NOFQaWgnCRYtWScswbgdRgxx
EunATzjMrCVqcbJ+Nwlj9/jTBCNt8G4PEI4fzs/E6G3wyqDOT/zFa2v75edrbQmc/zRxTfZTH4sy
y5FVjjZGjUyl7Gh2tjRRVyxY+dWZ5/tcybW8cGLSsZ2q2qnD0jBz9LnFFonQsQo63f2UUMn34ymd
shOSnopGCOMfu8N1dDxz0aVrj9Adb+ErAc1t/iFnvMd9tbO5o817e/Kl/uVJJ6bBQftFN1EIAgn7
7XQcgUEcxF1VV6OOJCpz8TWzLbVpKKNN4rkkvitIe7wuvBIb7Xm6pLKLgAputGXGt3GdJKOxeAUF
gyI1ceiYvgcj/iK1zoJ7Gr1OHsYE5+WdNPx5t9GswBVMbs8vAtt26VUxPlBekdKde2BK6EGscgTJ
ZkCJnIL5ES5pyo9cvcxFdacsjCwb6bYvtOv9bVl2C+C9GAnV9TPzvmyL0sFPRtEGXqAbTix1VKcp
G4z80OlTYcGDVxytVL8OvoRrJPGew5LJSciO4VE1IH+iTkSj7T1wHD6NWyBMoNl6ePMtN7y8i24V
QOpwYxZUzJUcPTaN8FLVyph35fXu0Nar/xz9gDcLPi91E3uTLqVrS2XqanqmKK6HhRz5DdDSxClK
A16MNw8VGsSezLoAVWmmWkYNg5R78Wpv0yIGE78kCborwsnhBPNx6/0zIyRO0lHRtPsmrbcZINqr
oXevRz/0DeT5RiqX1rB1gUNiQ2N1UGSxSeHrNfmxirvkFjbYtdcdv3EjtGdaTdXO8dIgF8q5qfEN
u48KSbgXflxN8u9iBFnCV83J6OjvG8ado50Am+hMVfdIdDBg0/zeG7rHusLc9+romvPge/hoMfzX
9jBeNiIdakoTyrMDfnhZBVav/pvavR3TUva4fJrWDzU+CFzLDYRQtKlWv4RsS57jkuRBvi+CMZll
+FFyWDNdxFvyPJKWUv2BarZC4oq3HRHvWuU0qSESp3THGUGSZ5h0RrVis47d3W2nlmCdFg5d5tJv
It3ZlWDbcv9cn4PlKUVsGJP0KAPQqKdaESqKG639K+bShdahYbom57V7KzZgQdGze90DEBukmbwI
j1My/6biBvUoqjVbqx7ldsKSHLzuDqhyDE3JWD+CGFtdH04PuXSh/asT6+gSbyaBK4z8VjD7NW4j
8am1ic1oAke164ig4oLlwY+zZ4dd7yrQVMz7kDdMvNTgL8U3GnIdH4xzHk4liorS0VvGlbC3kcqP
/H8pga/DDZumpweC+gvFIlEuZrw8hwhPgSO2L7zP7uppo/Gp8Yamd8S+tOTODcpruyH2PT6KbNE5
XYE8g8pUDsfPq0y9SE31y9iLpeqcpYOJqdpWLR6NYKjlKHFXHiRDFYwN0pXAPP6c+C9NLnCSi+VD
TJ7AjXS5bg4KBcQCwwcvoYavxVsDaNyzXnAQYKXDpRER5nbSdj8mpBWpjyw9jG56tyP+a6Hfhtku
JYRqlY0CIytyuHdGFJGsqUvsEfeQiObrUHJCx8LPmcMx0vJIlDoWI73nStLt/cL06T7V5TcedGX4
3tZvu48PqvZRaXeIEjd9dlYX6n1LzL4yI8p6gAWLc6gQsKNOHqKJ2QaVExqxqNxIxOa8SMJd3Fqa
CaHBfDlPWYt5hJX1upaAoiZcMO0NbUWPJkJZjts5Nk6zzHRncs9Yo38wuOeo+Rb9/pMXCuy5d3Pw
sRyjawn3AvevbsFntixgSbe0HKctICIfoKLkscFDyP7DBzS9Rl6VX9tHHkk4dpRUJ/PdQJM6MlLl
2w2d5PvxTnxVpFZIZFZiAc08VQUFQseyPY3NvQvvODRfXLKYFVbw+UeSEhLOeXSOfLmgZvDBG1Q/
CSeZsBJiLxyzNgOpqaoKomh7yuS86AeUFnWL/CJZTrIPj00HUtbP1FzTDThEfJ3DXRCwq/ZgXL6E
YQdMZjIi1/MtTdvzE9fnagMODjHIwsqNBjD5HIgWnVqr5bkZ9YTsD0JPiTDDk36fqqUZqhkq1f0N
D4PKS2OS3GGrNnOjK38KvNm2yys2p5cIHCAZFNRU+/+9eaLs77DR2pteLVjeKwxHmhf0aTdFeaP9
D0jz1RzokzC/4gMAFBrE47iNiYxUhbjQGOyld3HaPz00y0L9qWqqfYyPrPt+Ku5+vquJMZrbpjo7
KU5XqNNi3Re0H/b1FOOZHCJRP13CsTsa6YRzwEr2572CyF5xNzAZRcQVZO/rS8ehYT7O8k1cdcQ/
6dOEOaOuy7BXpKTp7lQow2Lowc9APy6F9VQCYW06jJEyKj3oX4rrRimgEyZ6AumgD0HH5wGkclPQ
vVLU67b9pzq9P7s1grSbyVTxpXMPxPdjHYdK9O/RnHsPk/a7TNbGgMpNdSi5P/fNitV8ABaDXHKN
V4UhwyiWPuxt5AhcKjPbuTABL/5E58YHvAgsXzsgFhumoFT0NNh1moEk6pT+47CyZxVo0+FE3hQq
68s1J9ck9aIW40n/0AaPm74fwaSi3Vp7AMKS0n3pjtYDOE8CD7K+TD23XgkELGzI0CQ3SFAquVl+
3KmAUaSeuXYfiVGDCPD9B9EIvRhyP0cC5dr/S27S86jnV3a8qUWfPALaqgoZ5c1XJoMCu/PPamCF
k+xvPai9ULdxs4KyjHy44DIb+X7IaWkXEbtAo0CrIM7KRiAUpmBGv6/Bq3Bo+GG3/v0OnjWxCkWz
BzIph+UpdNJ0rFmsKoMszGv97MA81IZDlHXY3SpqXE18NHzrfQ0jdX3MebXrEffCCMSim8NmALqY
Z4yMUhoDfnaYILfLh8QBHdQF1FGaCUX5Ggrypk02cjRyPOU+rkoB2JJA9qdiQUqCjJzNmgXbebu+
zsWuH/hgWf5x/rkr3vLpdhQzIDsLnUH8OdGdpS1d2cM/h8oPKxCuHSr0HykGrDAq/qAFxIIyn7e+
iDO/Uo25FuWuGLntCqlxvgSUS5EH0Fe4i+WPCoNThlx5WKvzsO/BjyCJGYyFqeR5r5ckxbOtpEBY
E9TBYhQ0hpRk651THcLTuBI3pxvieMvf834emyc89ZWMxnpfHn4wmqi5CLsqT1AmApL+JagbRHHT
XhEYmnPKm7ANZNe7pTGBqwDiVzw60401inLlWV0z9AdLnjf3kjCU2PoFBC9lywVlVyrrznXxLUvn
GppwCACB6+YQDVsGsGtZ3HC0F/8vjUJ8ufAPImK6FY933LfXbbBgMzscbxugPfyM7RGoiYjCpmrx
63OgtnzBnDmXCNmFBdnIO1k4kA7RTOBkdAo1/LfzgBcBOYz0TdIpLlm1o66L5cvjMKhU+oce5KEd
yYXNF60ffIrvJ6FgKCetiW4If/7FgdV00LXmyqbXTXEFMLbgcmhVtdLpzpzGJu/W12stlt+QwItw
gS0OXllENvX45G5TZOJO82QRHnlQ/TqRQRcwPvrr4+qkkZ/kVZDeYWcWz2pztOqFh7n/BR5NT7ey
VPdIZybNOthpT7V9n4ECa1kKPFfDzdttcSNht8Cq/2/JkmxXy8UGPXxZdLVgYcrTMEjONGKk1E2k
cLW5J5hGBZdfz/YuVx8cwrlkvA39cJeQJbtIA6Lkr+jIV+me3yrxnEDlm6S9Qj+vHG4GEZujaBTy
Ngko/PUwtPBcTRwegiamK3sgAw77UU8MHEMUccnPaiM4uyyx0Eci5JqHzHj71Vx5mPbwLBDe1Uvv
uf0Tq6EEcu0AThP4nT8qjZiRRS2lfMCvOyzvMw4swQnt1ByrI8/dbAfN11ZxHtOszAsGElW0f38v
f/1dbvKDaB2nJGPqbAVAsOetV9N97eoUtVAUnYMrjPHuukQNmyYiiHuCdjMtxQSYce/DmimrAtpq
gUJdGhM5Bvd3zzlTS2SzCMQdoLoO1am7kVbstijiSfZ4R8bTVpgKEE+ydwTgp4kvLoCoRyk+rkhG
ETsGJ9B2mF88mcCQo34m0c+FEFRyqqIvXWsNhGPwQepEF4hNOb+mVBLC7jwAmHcO1t1rHrwdNP2H
YEVCyrU/P68GkXvjAfjUNW07wfz3gR+D58L+Davqv1Mty5GS8JbctlUlfjnfqRreCL/JIDJmvn06
sViti7j25l9XKlbb0t5Jk/clRV2eb0a5q8n06d80dVYd77QaRuJXru3dhDrG5lBBc4NJLI/y62Sk
cKPAj7i9tJUCgZNkO0r4pLElY0mmOkyGb4xOjDGHCGoadIyfgYkJ7yk8QvCC/eAsPBIu+TkM+Zl6
fbJnwys2P8SPSJ7bgIgilW247PBXn2W7nsFCzfcc8E2ZwFxOx2MxbTCYCHLMEr5qpiYWbrZ6qhbi
tlzF/aRb/SzyiX6K3aMUxxg43/LlwAk1rlg+TcvWbrBF+wr3JIkD4biOwSg1kgUUIFbbpbsaVTlu
W1eIuqwPe7hT2dWG2nPltV4mb7qa4NyR8s0/SszsKCC8/hSP/zrFLWlTiVN4ZdSrSfR/m3iWAPnG
3hwBhCShqqWkwMhnNdLBybRHKFPVNoMH3u1fJVt+pX5rvfIcqutceiNBHnF6vREQFP00HPJqmazq
htLGWT51JDTsccQx0mtscDqyet05CR/5FlF0f8AOdPINvdKWI6jhX0ZryiWeL4iMtYsNBwiRR2wc
BDbk++eFPvZNtTLq21ghykBEm91jkgj79+OER60ePw6vyeuJ+M7vLqsJVdK7g/x8nxsaPZMctX21
C4yOefmgqvVMx52cei9U05sJYDPIFC/MjqZ8v0BOm7oJBPKENygkzw9U0hBf7q+shJNgvlzD9Pn7
VBWcw72JH/VxZZNO98PW8RkAavTWBz77RZ7+o4DHMegUgHZW1IaBXtvujhOupnYPbefXAIS/vYpp
+txNDFHbRBqTyaDMOrc/JyZv9U4wcHa37bZidOJF+5Ar5yP3D3OQy2tXTgfd14YwYCN6Kj5oCrgl
dOg3Dr0pnOMvKYKWrHqy5Zrd1otKf90mgB0p6pZnjXCaspEZikSPVJziNu2W1G2SG0cvCNstZqYv
gVwq1tGR8xOOd3uP3fQWb4VSoYS4Q5sGgKDxHmTIosGGX9URUiRQSyiWtXnM1ZYXYxC5Q3xdQls9
Ge7vmecJJLEd9Y/IKdXun0Usagr2b3Q0+Ulo3ySAY0O6gHokvGrLTLDV1pAtw94cOwk2UoXGQbtM
zv0FEkeJlhz0cS/sVnqV2OVw3MapRtek+JlWmbb534y9FXs7SqYjdgO3UJ7rhXjOoqxL2IcaTLVW
Fs36oDA7Cxm8rlcwGERtA0Zj3JrAjsP/kDvDEKtyBaGv5tkwhkRg/rlV3Yo89wdpeH2bdabVQKIC
rRXmNXEGb1YSlfkBFwxz6QLIRIxZOmGRLoYpriBYbypr/DaZ67SUe4/YtAF0Z8+K3XuDmZphR4CS
C2dLyII+nFsedeE5eml8x6yUheBJJ0rSIg+HaqMSe1idsj9P2p9TIruLMp68r3hjHwZytZvSehPF
mukywMNq6mc/I8Iwe3vW0DCrQ5mpWXHV8py2lbOG3mz/vtkpnDpFYNwrYuaXlqrAV14rNm23R3C/
oheBvLhbPb+C8kpviiRoslQez/G/2EXzgst3S4vFPXHUTZaaGglSdKwo5WhYRZ6utGXhji5xMDo/
P6SYHylVgNs69hwYTiao7XBPkyKZevxNaL5Kce9YRdZUu9vMLp/5nny+wyT6MDA/97kMBq+Jv34A
i+0tJgdjMtjShh1LEyR0HboT1SyXA30Yl4GKZefxfTH4SioRLZMusYNOVKOz64l5Ro3t+yNcu9wz
Q92ooHYSoWlFiRLBUXY18/fOVQvWyPKCaKsQ0tmZRdsP5YhtVtkvYoJviID7EA+vSj40boWOqOtL
etSlZwT/SRzlU/FnC3ibXfEKbkTNO1k//E4B4ranG3fCYIkML2TGPg/qLN+WZpQe1/apc/yCmI9/
qQaSfqtsYonoKNXMCFTDCtyycE2BLtb6jylSMDXhb+bqTnjOnyEs2Vx5w7+Sd3NKOCI2xfzO3J/h
M6w0pY5n88r/qlwr9WLKoeuzNH6WwDLpYoHXi6IH9uOdFPG+Wg5htJJ3244FZwpSHzA3Id6dbh+O
rIJw2wffGQCQWL9oDg3uiNL0TNYLK5Xv4zQrnImR1MMdMVsSPltZveZ4XHx/ubFjXp9cRewcGLWg
b2r4QBa3Hw+75F4qU6kzOFSs90VwQN8nqoptuIloLdbvLqvmzQFrJcQ8tgPxZwLBNiWj8yPXSGk2
uHiQ43iHw+857/cu0+N6PJCDvDJ82oa0P+d2s+xhPpkHTrtMyFx5M6yx2+FN4dkSs1tOn8XlM6Qq
GnxIZz+h9Tp1zI1owUvWpqofhV16J6rA0/sTv5xXtLUC/+dIm73uyka3uIBkgsehoNrv3Gisskm6
qw4M+OjYsfGKTlRTlyPWLVGRr+IdE7pIx7+G+++/EmzwYpdy7U0NbBFplCasAKs95jaa2d1Hh9ox
Te+lA8LG2tsLJTK3ujp1JC9zyi2kv/BB7fFMzhoRBD3UTzAZS+7D29q0F5+o+CTNx1tmEPh9n9g0
hPxoeSh4vqvXGk/QWc572m5wkSNd20aJa3ziU27G7S2Gkan2EExNLof0Rd76joZO/SKNET3XrMBg
6207evHS2c4sGCFZPa2bUcfbcfdSG2OwIrJsx6UVdLGnfAg6uiEt3j2KQCHR5GVjsMzybRX8l8W4
nYhLDVhMM3H113OBTKK2RteiAsoA7pPta/JYOOTtPJjqid53WI+jS5x2nm3o6vZp0FCa5CBX3qZC
bd1uQEzz2KwDP0UTlqUDQG39b+RHQNuZXdjnUpzQe4rVoYbk8cNN9LD0/727aqWM0D8lTjnQEFBW
zQiIoevR0Xh0usS39etIW6WAg5h2WTKb1spxDKUbGdtQ45sRAfWOcDAOcrCf3+tnSGgccKgkGoM7
vsEBoABp2xUBeBuKwe5B06vEZD242sQXPzfYGTEWi38hL5RMZNWAzygBzWqpr5N7aOuPz3xVpnma
bSCki5OMLxcaq9LKwF94WFMbysAW/IceWw4Hm4ZgtgiRuq9j9QLfR4PAuBTgVO0LBtVLU+A6uX24
EI2rFzzrkMhwG3BYSWMzksSD81R6+kP/SopShQvlCt29qOwRGjFa5EJF27JO6kXJfCzlXH6gxWvX
L4tImPnhauS0q2/2AclNMHqVuRRSpyNsd2woqf+XkkbXezN5M80SYfwpGDMb9+1mroXm2rkId2da
wuJWyydHtmbeGt0QCGHv6NV8XK+aftb5TfWJgmemnzHfa54Tbp3Me6CgUzT38wry20c9EDXVbk4u
eSeh4INuOP2rvOpiG+QX61vUPtkls7a9/t5BBsHjb3wHdSdhcX9BIklOjiklvqhZb1UsUfZFEdYS
AacEnMBxXindALRj9QKWilqT+04PwKNOh5vnj05d9vUPnAnK6TRLmROS6tmJn8K6msF3Lg/GMTvB
W+D6rs2L6lBYXJ9X9LKTVwvZ9qJp8h69kgYiY1i0K0lJDDyR1e86OZ43sZDH7lLiYoJwZ//B101m
TxytMnAsMHyt2YGs8SZIxOL+UCFemIFjz5HGjTZp5eAYWsIyop0Xi8MPcnrV7a5lIglUbAcctOHP
45gLuTgRwGTGq5A4dARzs2i9R5KzmB3tSy9YEf8UqvJ0rnu1vBMHUHBUZbiWuNKBjUDaRecVWAnw
Q/Ze64C+X5LH+w3j7/knGbXeiy+6bHM4/izdYi8zrjPVepibv5nUC9odyYXU3ApsyNmb0esya3xq
IMh0Ei+AaZ48bubjboaJUgktyzPgLSVbYFTSE/mB2g438d/VDlKKnyPvg7e+RiTfLh4HAJQ150uH
E/3qRC43iDdcExZ1o+iP4pLUmZMbJE79tSBMhka2kWOS+0Q+Dt7Wux3/vqd4W+RgCITP2RoJo+wY
wK+EzSx9i5XsopnewSCtNrtqwn1QfCqJOzPW3UwypzApwO8/J3RXToK/Zd61LGOhH2YIHKGAAjt+
BnTUhHtUDiHPtr/qA6H4SVWVRNGG4eTiygBQ/tYRDWfRBrlKnDWW4W7YKrVVLyGjEA0lkafRH9Ih
aQxBiPHrpWU8P+fwuK3BMntrdDCELlZzhVQ7yQC7pHPZ/HEuDhWprW8L3ZjTOXrjXsaMxwSWdKNS
XCu/wQM+t2ni20oQOnc3FebO/GIZDABS49fUxEdh+Z/Zyz/0Q+8+0gtql2M8DMmgLSza9+SZGkRx
vyov31wsczF4wMwiPAY5usQTixf4jPZgDDtd3goizG8mZB4arnzqDlJUCDdGysOskQpKVJxEbN9s
YEOJYLUNZOc/Y1jkFMNqIqPKJYL66hBmyGH3bhoxNuBUgejJtf00jqQAMKxOmbMD4DKgVnCasEcZ
4tP8+gjXMVZbBuMJjrqccc/TwgW+t7kF/vN8nJ5JzA23X/9GdjPv22JedQknXarYTqOhjxmsJA9R
3/HM9Kw5nlgdkPfEhKXXy7pQtIUrDW7eBXsSXts2Uk5o96d6PY0Zuf7ddLFq+TBsu4d07RqRS5cH
RdCtcXAuDzec+WtKWInH6fOV4Vf8UmfsRJ5SUmuDussvsTXtY3/962ritVtA+dBIffDL9laWkjvN
Imav7PZ809DGG6crtEf0RW0rucly7/nsybN4GgeNUDfZx4hLdbvJsq+QbD0eXnQAIB1EaQ8fZHK1
d+jKJnQxw1L3iAAYJtr9YKxgScRhW58IhuAkVTXqWzToHeejOEcxQZP48ohxUQoVvGToMfYlYAi2
Uen/b8hvs12JRazePdSjEcKRTfzTO79ov8VjOPb1jfka/+PkEps1/U4tMOo9DhWPmz8YdZzpqQ4E
Q1y3zI824/d4ipCSckAwzjwJ96jhAryToiirQGcfB2RgsMd1YWUF1hvEBg926wYtwrICT5GnTx2c
Sxid23zNcCTOjj+Bxubc2Aeyl1YXF+b6kvE5IC17sBB4hWZJKbr60HbBJg/nAjTk/XgHqqSOYJFP
2E43G9dZBGh93zzrOGnXSMoq7xOloaFVfalA6StlFufCNWU4SJzCDi33Nx+Qj/81OrmD5HQLlDMG
Oi0vFhnuya8T3FohoqkldZvOh9+PAlSnDgatrQt4AtO+SPoOAjUn9nFXKNkoHCJa2Zhz3NFLolpK
1cfyP9qpf9ukABrRJKisz1FvRWtMvl4wwNN+NAbhSVw0NuaGH/3HJ1MIeUEWNhl+U7O/vK4mMrEA
kA9/kss81bqU8Yk3TWHkSa8E9/2jzVL0Hb+YPjR4pVEE07AcozsBYtMsA5ZJ0sdmZbvzMBMeW1sx
TEagAFrMYsQzPx/q7Wn17RSby206UKJRK4YG9CuXblSg0QTvYXhoO0o4HLEDTjfC2AMnfnuSl2kW
SbffV+Ea/To1I+9G6LrzAXBxPTVTiXS4i3zLaEjMNBvp3TZ00+ov8OUQiBvqPaVh4w9PV13tj2Sd
4F5JkDmBof0F0SOgmCJl02957NJ9xv/87sOuuH4KMTEJUgtE7OE6eskJJZbxwARHchosfdTeeGLX
76run2KEAAQaga51i1AK43O6/bsBMZWkg54TCxCJwrIp6qxLGm+O5Oq3xny9ncrZ2znSYE02zSWV
z/BE69nr/tpZHOCRRX0Xw33qOYgiLL8b1u/kQAVqDCC3uP2JmLAaQTSnVO10KmAY7g3bHyrIZULs
nLJ/2v60o98CrL+BfnPQJXc/jUM/r1gZLXUDK8mCpzZJbBZ8BJm6fdCTcO3kgBh1GoM7m1IlbyKO
d533qOzRYYNpILjsO9zMCDFxHOTmT8W7vXVtiOG1ar8uvxtPdtsQA2aMrc721h40JRNyHfkaMJZu
E8evqg4hH9v6hqVGHubF3Ei0KhNW/ZH36v4ZeknY3fR+Tsbbz22XU3xQumphaIgNkhoWVi88qQh1
ZxVMT7gb0hfwFWjoKTaxa1/VppkUQH8Ba56HC4Xe1ay7uHXpiRZSx0G3kfJjuuWsrfbf7896X064
3fXfxLcAwSySowkcspY7KHbn1jO07x6mcrlCBdhNro0T/RB6L1Kky0DU5N3ASneAV6NoONfVqFv0
mYlxMNBt7xRGpaYx+s5QvWBobpJfaHm+vQOoMkOa/jCnohXbdVBg1UOm1i91nHdOgLQDGbGiL+Y0
C5EE/AGKw76mxZE9aXn9OB9ypNb3GkF61qRscpfBmG7TAGF3/iF1Bc04jBUs/XZVA6Y/cjSeQdM5
gsOtTa029Yq2pteqzmvrIeAnU3Ixm7eHkp//WQ5o0NhU5q0wyr7KvZONFN3ynSmfqoENSYnYZp6T
XgKNO71Od50oHzAP0kNu71EVqhe8U2iSzrt6kmIKGwx+r6hnOsPeiPeMso5/yIbMX+5WSGAM6Ypm
8oc9Gzz+6cHVjnku7Wuo23bDu2m4otYITCpjfR+0pQVZaFmOMqN2YCkwjrPSkpucltP0VpmfjdTF
201fZYD5AtzGeomwV7NTbgvAplZh3vWUBFrnkoLxuv65qho4/VDRCrkVnyiX5DDruicL9z1bu68P
SkC2+tPsBhcsVhnoj+kRugD8Md74bgTNaNrSC43/pZ2er+A8WTx+DCtIL3475RJojH9wOFK0cy3s
lY46kU5lkL+ReQ7ptk2Cncvy3QOHSGYJtQ78VFb/lQnxuIyCxTN5Ddi4D0K1WxYedsbUwSs0bfsh
d1pEVCIlO7muL81vnXoLm6u0P3bOGkjc6MiATA6OjoqPyJPAiQbJrcquDjWlgusY/N0uw95Hgxc1
yG0usIVgPRf2Xb1MwMWcTOcJWmR1fQiMNN3YmUV1Vjl44v0skyEviiTcj9QG/bGwjX1EJncbj1z8
2JmoIwvdJkxzxGKxzQ0ZlqFrOjMAZihlwfer/nnVnVS4EsRiRhRpUHpRuGjlERknzwCfRMZWFn0U
h7CQTwvd2rx7LSQFJTZEfb/wJfXanWn8YF4M8WuBEY0oSkjGcBluzqdpsMc/mayTRm8bq+nAm71h
dyV6n+dmC9KW5PW6grndjroYYGXtpx9/0jvYPWA3gj7/EXWPoS1Xs+m6B23zCgldfs28v6Fcyu0l
LHIqxQGC2xqqNRb4RHzc20XE4UBbB+wxJGmr0EdSV5oBfK+ACbONwqsSnJk3vQr1REao2gvwvbY/
MAjZ6SipHPCJaD4+bonbf1PEbIScgkEX35nK7WbjbSSP/E+fh28mFqFqgX5KYJm1RVAfl/b8z7Bp
0EtWA7g+phtKeD3i7nF3CkqorUskDJWvtGF4gy9Fsb3E6VyJl+jYD/GbGcbb+BxVXB4V2ySxe70u
hdRdVeHQoK9JTIXv1dO6dfRn5TUl3QsTD9nLq4aBStxqTmkjRTZTJi2D1rny9pJYepp6Fxz1GO4f
bAzHuoj+sTUVYyx0Fr3+SVoAo1S1g2rIroZChrChm/MikL7oFrC5VyM27sLPetdNLMtMPs9RlgYf
9ovahh6Uk7uK2WOLBNif900apJ2ptuRZZMe6UR7BiOWteWQZda/c4aECyoOJZf97If3ASnfinGEC
8ku+no0VZsbDiumLHGd61n9A6CMi+8kKd4D7TgilAt7JRekcAJLIR+QfttHc1zrwEL2Yz2cA6atz
lyPYCh3p30D+PuYwvon9PsPdNVsvg1G7jVAIxIKSl4GAn7SBopy/Runp8HvwWyMThYExndalVNts
NXCxAe0eB9CKMLmbqxvawmsUwP/RGLF5DLBP0dZgEhZoG0mFnJun1N9wB0FRjuI5XwCIkZNTAjNT
t1ALtAMMbv/HR/PxrkicRYYyi17pjuTkK9gSQ9KaRSHnS2UDVIda3ofPiEVo2L5RzszEGOjn2eAi
Q8cs1p36MpAJ9n2ko0pFw5MKDFGy6J2lMyLOYFX0kUahwJtqxGXz4FftkPjotbJSaawTZ7LVg9+x
9GPe3E3kCzYCHEMaYSWbkO1LXJ1cJXd9YH1MJ8optq5MJYBAv2yDmTchGoXjK9hW9U+2dfyZIrqD
8gK/g0ALbvNVFsQnI7ipRMDn6BqpfJrJxlzM+MYjPhXUSbH1D0wEWOQO+ePJzAl4YQLX7P/NCQWM
Y+HaCeJNmZ7lUYdf1R3YuXqNtMYSUm87m9R9uohiTMuRgSXgOBjvAz8h+D8IrwkvCj3sXl6B4fbr
fQZWYK5S6OdpotFVJFIdXY6xDKCs2QrraXOXFOCnXSIurXM/O3ZisPV+k4dLW4knVN68xKUBtIzS
LBWW3/abjnnkSfvWGTGNfRvQOXw2JVqZAAvFfwTHO3sPfr0eNCconDs6OqBwHmuRxWIWT6A/JZj/
xnqlbiM3f7RZKGi62YB75C3ExHzINtwpqC3QgTSnvalBs1KP+SGVwlKsd9ShYGpg09cFN5YwoAvL
sjpkG/awauaY9ea8QcDvrweX4k667I0zgWkIpXrIaEXBeaCqx95IkYR7GkugB6avoimqIUNs1rVT
NDR45gd29qr5wvAjOZZydA3n/67UP2DCGGJzxyKbW+4rwg6VlVo0CBzLAc1j32vjK0f0HGMNBo59
DbiV2FLDzDvwMhlAoOgfRxi5XqFWQE5JJ6/L08DwJ5udA71EQK+KIijAzNYomlVraTReb9o9N0m/
GhyTv1rpsBB0a5Y8BjBnA40vXVcizIFlzLsRW7KJNb5ZOXePzGRlcPEG65aO3S/VOM5yUYYw5k0a
lL6DxQTYqsXACqi20aoKwgKuQ3SrMB2WaVl/8rTApDZKP+LrC49GwQ7IEEvUFfIo25t1yfAV3qf1
oZQBH5BkRSb06o/J66HAwtXJGrElweJaKwAyKJFQh2fkOItnffXkkvaXnQRYUElKIxBkOUJhtNxN
BUcD8gTGsytoBSmDccB+I884MfviEI5/bYnAxLfQtqMSW9GktGzbN71+PsHUt97chAiaxUiPwEVP
hkKPpHrkEQEj3thbQUJqvWVYYhARV0LPtyON9lCuYdQ0Dl9YAeC91dJwUAzMJ0Oco02vklW6Wmv/
KfTtdnN2C4qZo0j6+SXhQegvw8fBb4PmXORYrYlpYyBkXGVPGsj64Jz15vy1QZ7CGuh6DWTrrG9/
Eo9rlTgvb7BgUpp+Rh82egTKJbPVNsFXkpVNTHvT6w+8MF+ld/giOoQpdGjG1eLmd74p2c3PwSwB
bctXzXXmxvoxCrgOWAkMJsyT1ESQCPrEXLnM6m36kiXgYpBH72mj5HHiXhCOnsW0AW0YcpZI4Dfy
r0VpaPTmjVX+nkV+ZwTiUFlJQNaSVvHnSkrbYV35NnSRqdys2hnFn5O8w0lfQO7NsV+lJUM5mn7w
zwb70GPQzSwCFYnzty/98+8s/9oGd7QLrBYNP7OQh6lc48161u8Q/4JUQai+8G5kFg6TJ+oNpI5u
ONR8wEzUNPat5zbLkoT1GbRfvgJHT1c2bCZjFxhKfgzfBfFe3kBnw+7x7ZJWf/nl/8WlzKXlm3II
hdeggHA+61yBRWCSLh+CHdH+72Nl/73V9Da8vhRXai+N0tUYDh7xM3ypPgPo2nC5gpOSKVJPZ7TE
n392TLHyXdl2O1iw9kPIxXVPpqXOtLkZbtYukcAau9r/PnJ72K6aZ1lJlK9F/4fgYJfc+ZCFDuMx
WE2nZjX2tbrjT1ttA/WYMIndaa4Ap9GwXh8i9lEUM/k+2XVZFA/NmEp2YZaJvGUMCtfe4pSYmwTz
5B3oZQEMi/Tp/p0AxaNElodN2gpH0dXHGc38cobrqpEXe7cS8eZHCeWQXIi7ygidy+VDt9+4fNJF
z4Fn7eR58z1Oq9j1PeMVgqohMP/g7bW91NvXXbzqxYakRKWe2pObLkgjocimraCvOhi+WZFIUsa5
BkOgpFoKswk03UHJm+daYq0pbJ1WzNuW2FdehnpTahOsJJYzCRl2RH7LVnOavTBBEz5QOySme7bn
f20fGg7wjGjH9O2D46up09xUN9Xgbc15jBJM6qq3oCmH3b6voh0nPEdKp9iKLGOP+ohFmwPTLiXg
ox/byPb6ExjNaXx1MoVuuEy5NQvP9hLTugLR8xY92eaRLM/w38ya+3n01ycgjasKCqXZdbyQvu10
Ib5khU7nDikvA4SbnG4Gd/q/s/Hnsfp0saf2tsbGHjDOf0pPxhZhGUJvrZFBnIbhfLh1YZxjP3bS
D530qE/pQK4IuKnktskyl28x6P6GmqHrOgoYHv9239HX5xnSTkNOfkEnEHeP7FojGAwmtTswOKY5
HFUmEpaxxJ+uhTlQ8GSsTDmWDLwVMVJpAx17+4QTvyYieFEf7sxBtoCYQ/9DqbTzspYkH8xai1Xk
NVmvCYv91zNLb7sWlV02zS9HYaXkYboQyP9yZUWCZia8DADx/aqnm7+384BodGTAwHlpW0IiFYRK
vwpl37an4cunK0XhlwzV4qeSD71MN7gHXJ/d8L9Oo1Ed5NwUcAHocmIW0wtCQY43OA0TFtjTQpWV
DWc4nEWf/23yQC0/0bk2P/307DCzdGDSD9xkt9RChplfqiZ5dJB7+e2H7W7v4yrZPjGZ5RZjyeH7
MA3p+MS6Hlt3ANpLabxudW0YebMBPn5gpW3p8Zo5RY/jnj1x7qzr+TrAmSUtQ4j+LqAaxnKRHyRi
taLMejRCXOR9vL4bebEF2Vk9ky9y+oROwjYpJgmrGgorwhucNaC5epXP2oNKei60Fem7Srznk+L1
W4RYQmviTUukGiAcn3mmQSS1g+7r77hfmuBhXMVWOpvtXiHewx2EfdfN4ldry+OayAFJ7MzHnivl
1jS849madYjqBIwW6r9iOgQHLsFRy6UlT/wX+Q1Xf6KjHne/rdj29pouOGi8HhqdoFIlk+wma8y4
fo/fc3bPl+m5xfBCUzopwrRB3SyHIwfTwualiQNUKuV34BhPNvRGXFtw+Jj2tMZ+D+ms2iXiDkw7
hAkeo+95cZyd1/rSKhjsocB8dTOKTSIhzVEWmfPNLgIp0nyj3k/OFW08hmcZ1BT2YkYgjuiMOjGA
+PqlGqeiZkWPhpnDdZR6L8GbA2vi5oCjowA32HIPoCvEwEjyseF102OL0vdUBkepkzRQKS4+Kx2Y
THklmTcLpEKbzz6eXszbBFyfSw4kebDWKQlEw7Fb56Aav7iCKDu3xQq2NYKG09xS1N2nxaz/GlVl
5usW5CJe2uFIc8MvBf2pyFVeUF0sT+1l46BvN+26zFJjaY+tr6PJ1iExwxLbGhk5t7aBgayZuTRw
UxErLxMGThyi1cPkyUtYFv+MBirgLW+xVhOt+vgTfaeiWth/t3DN/3chPHY2eBLK+JnA4qItDtDO
NCOF5VJaRo5eswMTA/37zYoQceVHoLJJ0GBEx56qdvjjlpPxhlAwSsE09nm0Px6AIfxTJWoOKtdR
8G8lwCkAxFAHKRraeztLhq+pashQB7gj0ZQkMQm4bLn1KxQk3EiO8qNtlBdJtkV7pyObnz3pNZL9
k1fKOxerOS7AVc+wofksUoQQYlvFWLC4s7ZKjWSPoQ2JpJqZ/DfcXX6Afi/ylJmvSSm0O7XU5Mv7
2ddLMrR9xBFNEgWfaTSzhrfK0qh+jHCC/1Cdsa23RdVuZ9lLvgfzqQNE0sIj22gSB9J0dPbW7ts5
iJnbCX9MtbX872jOaB3XmfkNMs1mHO4By0E8sY24WcOt5yHfAZITW+LZwyLSEqfL0RmrIntigYcz
bXVDr6iiI8n5JW4cyNL7ioL21AK5JvIzZH1jWaUykI7itFAsz05wTHR0nkc8BC5zi1v3CDL5uhlA
ukPtG8uXGIczl48srkRpttk81Gq8cF0Vjq6XQAN4HrVy8/cZkKE7xu8fXR0xgehmdLIUJq9DEhYd
ozUKtqPJG578JB6gg8IrEHunC4gwYWE8ZcPR28/F/k6MZqEkiKnaRjfhnJNd61Co0IW4tWzw13x0
4PMcnEf6Y+jQqi2O31etexmtGDRflmqZE5tPKt83LvDC4RRRt7HV/6e5wC/eVmHRMjqFWOZp3fx2
F0FYrV6QS4UaPssZMOO3LkVxFzlA4Jyc8kNxNAIF3/dhZ5i4bVLR4kAsOHWnJxJmBXKaoReqIkFf
6SM2/mRwbBeWRUueEU2OCBrbeYrtiUXEhH99UTOPKYUs+2WFSQOlvspsvpV4UGlmJuXWWO40pBPM
s1q/gMtweGPRSQIALBEbXVaWEXxACBX/AsJmqX94vZ6G9hqeB+NyAfbOCMsIoBX5vHfm5+/6EvA2
97R4DCAe47IkkZYhRmMGAFeKS+qEv2uXFdiDor0IrJL2skDe/ZsmnGMx7l4puJpLgi9x8B2VNWp+
vupaBf4+JRIJSbH36yKKe03OvgkRIuudRlNwxRCsaVZfCTkReI1+XJ5wXCnqEFV0ke4RWewfvRmH
waGsJjrsntutJ6doqtf7Fqt3Jq4oA2LfHZZnBANI2mPOtp+4hZpJmaSqExouKRhdlM1nYREkkvww
tC6SorsJHuz4kiWo/1ywnH935DKx9JCsfRytTqCnQakMaUfinEF5M6t/I+vZMYS87XeMhY+lBgN2
X5kphZjaeS2dL5TE3SHGq8dKviHTfJrqQAMp5CT0ra+4knUOiQypb2gSf2XJbXjPyXksrX2+xUdE
9U6a+xMvRBJFcElXJofhi8wZxq+xnekUffEQtttcVIfIsNhMbzLFxFS35UlwV/2flBVih92ceEKa
fgpHF2KAj1vvTzYJJEgUwK+nKScNyQsYqVuFEHb3TVTS5ejLO7vMVrkt9anRmoMDUX4T9vJpAvzc
fxV42cswLcOH7/uYZzZYhNjVtXaQ15GTH1vA3tvCeB+o8tLrWYDRfL1xK6aLnAJLCQNane2yP2Ji
Mra38yygoBv3PnD1nPnXFrsSwXUefQrpFejcPWCJVr5GkN0URKrV6jMxjhZq0kU2Jl/8F6MA1GBx
3Be5iE4FMjJwmwVSdLqmj+rO5oNw7Aq7+lueJkmqEIeR3tKa5u4Nu39yRtynEINfl+QL2cNr1ALH
UP7pZYrnwC53wfTgejOth0koniOz5k9aHtquc1WYoq1aPt8JvUwIQLTIMV5zbo9oBjnN91bNV668
2WxnTLekk3rQFy6wkEg+YbYh03tDK/4FdpXJw8hefZqTMl12vikZFrPxVaXAVgaysbbal26vkXH+
lL/d83XuafFJYf0Aficzg9X7/o/mtQon2j8/NYygs8fOGzG+eRycVVhurIynpRvvXQ5oi+pKh+9w
2gO/Dx5Lye0R3uz7sfOfPVmkGVEBa193B9Sbp6X+xQFpKUbYFCei7VC8JrWOW41PaWnTwmDlMw6g
Y3BQbEYdWH32HAucS2DDm7IycTAw0HDFaqciQvDYX+1HXxxB42Cs/4pduMx9cHVErYoNpC4T8WKs
VWx2QESdGqMZ7REtXtCgce65tLKaX5Xc/IaWBpBaDYGt9bYCnH5K+hAp7VHEt1sRPa1/+g1Bi7NY
uwZ8J3ShX0iE1vP9Sai2VPd9LBLONDBdEUmGfBOaXUMduNFQQ6yIGWPIqJKgIwGySyPiVaMbiJ0L
CZ0eKN9kKM8lvo94hedq3eUukmEVG5Adfzj8hl3EHUBCTt+t0VL3jDnsD+lRtTa1GlfGxdhJKEnr
QwmMAEzswPKQeDAf5uQ8e16sTtu3HCleSGMDurmNZSMufhWdaIaP8uRFMjxfe1ApZGs/efSWwE7I
jH2HKOi/PVBPukkdQGiL8i6TcZFdbAwQXCBjI6oRY9Ofvb/L4I3LBZmyMGyHMnwN3rxz7GJqWlnD
79akvVb1OEs0AwqgRpNpShybK6J93hSMoM5daybDJDW1PWlvPaMXjQgCt7VDYFib+yZzjsdPPn2z
ZJURg6GPGZsOAEN5ghrQKgEgWgL3xNmYPgMqP7/ma9CTEwzEq0LJeeqBaLYGmTd5FXy/vLUn16Wj
YfAy0OUrv4m62tgC7CMyZNP1deykcPXa9LgVok47FunnTbzHJtvH4fjHxpQpnDjlBHa7Q6hAxOFn
ildbaW6Q67VXOvd8iOqxEEfL3WTClsZK6taYVO67YtFOxUGQ3H8kWvqNIbBkEJWKHdExOHoehnhG
2cUL61boI3dXJaKeHUX5TBmGYonAvaC94iF1OcsNMnaT+5EcDgqKJdDrcGy3Lt37RKw/B8qK6NJn
sE1lbhgKF8k1b/ddzZWg6lraKCzS/0wRdosMSu9Qe+ZaaUClsj0IpeYdDyR+uSn/Sq8OJITLLq5e
XznbRGz3h6+zyikZ8pNiZ0ynp7o6BQT67Q2nZkwx0d39vqrtTUWAhsYWJKJLXZa55/N8wHdSVTGS
S5VpHj3quLNmE8GMbIruaugFSN3YF8wZfNJqTWbU7QPenNcLA0+3Ykja/y1P84l0KuNUlayAAKK8
+PwIAKlFOnuvVV+boAvj4RwjqkQPBRF+7e2geVJJD2ITB99cf6LiYLVPgyZfVxPeTEDwfZ+wix6V
7BlchLJfNi+fDO2rpgjOKG8X7z0wA8c589OmTFRqpe48/R20SZHtsNi1Cf5qScL2kurR7HxImzh6
+IBZlzO1McJanr5UaZmWeRKyIj1P3Knvn2B4q8yFlAeYpGXHGgOi1bShkwSYXxmeU66W6bR9ElQK
SvsIz8oEuzlfuR89/kNAn2Q6/4qtvnvlcs82MJ+wq61cf4fAOzS+1lvr9Sbvi1dhMMkEpIDOOpTv
Z2mvyNYyoHRj0ylSJzcJIw0GlyUrjM53Cpbvc3vwH//+10gGZsC1i3qDUDWvGNKEAjBccbhgwiFk
Y8phtRYlOHlwhiLKFBqq2e8tAZAkmBHkHDj+aKIY+F0ZC4YhAu7x+KTub7WMdxO5UW50uE7kQmPZ
VxS9wwKZbqiQgko0SuI3Tun7muJjWvzhcalfFjFHvoYTue6QyV4w3skJ1tTk/6aaU4iH8H1Umkh5
/aZMEzk6XDRVWhToa6JMFHTCAxbj/xaC2piJwdNU0VMVnZQidto74HSEX80lSc1bmsff1C3ggHNw
2AZWnD2JE0KfljkttZGedAWnDUpgYknFmjwfaCIGBcNfk8OgRe8LVWSGPmOqbFAAo4xN1UYhHcga
avHcYT6Ntpwwmiow/J3OXOGwIRQdCrFO3w6fTBN+XWFvyrRiVHupb4t/R5O7EDws+jmPmY7WKIEJ
RvGrXli7ymFVctjj2gtFaeZVimkzPAarrTKgrlhfRrOtDJaIUomWt3Z5AgLqvTHYUfpj0U83akYy
kbCYwpwzIAZ1kZH3lwNNG5NhxbB1LPau7MZDhb4YMFaJTgEIYxSxx1uUarszjw43dHxsNXgB1bAs
C7qlMs1sn6jjCZgZzC2Sce2C72mwl1MODMtlHf5Ww8IRaqtAkCDST8oDMZGD5iWkNp99sngRi3/Z
s+EBvss+zCydW3UtbE33kbPckmy3rzMkrB5EezZFRDEKl5RqYEoE9Nq9Bq68QDVYs33Fjc+EDJkF
WMN+eB1NWvFYBlNMm3PoOcT2WseZMTBMDRVYfgSKbR6thcqj+Rvu1INlK+ZWpyD/KIBHwSAiq/mg
ruRQyt8mx/NWuQOsEkRKWBb5x1BotvhumajK1Vm/wOD9JefOdNV0kFLDJqKY422mhjeMN8aMct1n
6OTQUzTutlihmzA3LOsWP8Vmdc8hOTWGy3Bo7W1sXrXv6Fnbrs85/cwoJIE7Tn0XjAzFvu0r6hKg
7ZQnOMoll8jW8ANpEQa6V/bPkxQSqBF4ONZ/ueJ8ZScojbzJ9hP7/vnY28JOg7WVxzPBhIX+e8Te
HOSTDgFy0JuECTPpTtmJHyT9tKruWewLCnDNBDI3y8LIgnEFGV+lawj8WArA3UDA1XCTV+j1ohlz
x9zV/sdDa4TX9ydJXYTBa4DGKNweAns6F5IflJAK4OoL60ZAZcUFdJmooLk97o8PBDWmiuUjd4XJ
mbrtUyGCssS6cHvCdC/Ncd/M90ofmvQqwRtP9TUBLcHBxFryPakNpJHLhptZnT15uwssDVZnRR0c
KgEn4/rcdMHZ+VQI0UAbi2eVW7dSwbM5EQpb74cUvrBDm+iPg6v9/jxtMHnk5Lb/BTaZAx0x7K6t
B7HW5YZpXbUCbo4eAYywzuu0uVWqxQgRIU9R+wva/WApIdz/BtXPHW7TofHwLcTuyiRXr5uDTcal
DH0DmfmxD2L1lqPvj6Oxj26BcP8EmHErwjrl1aNISA2RUxtj+EUC7qL8tnBX5f7QyyhOPq1hQCUt
leHf5gr/7ANvjV6VJDX9yUrqLwu5S8W0LyjtuJb8aSIF5QA0pTWREEO9SP/cFUl5ItjWP0gn4SrT
tdTlYPpsnZftwJM8kszBpGN5apKeZvaXHUoOjTsJJbSfkJrtOnif+S872YSn8J2ddRUFrjyPKQNf
QvOEE9GAlpm2ldQuyG1TzeIkW+jcWzrayZJQ14ap887Nn43Pcfo6e16GtgDB2wUei9r+SK8rVDIP
wxaYM7rkx3YLOV+HC45/2mC4jSksaSplc7CavlWy6bD1wW6FMfQL1R+EEbU9+ahhl/QZtdINrNjz
SIAnfqJ8gQ3T014fm0tsdQwcR02s39Y8Du0YEo0k+jIQga4ZsaJORMtImq/wslFAW/zmthtzI/xw
M45jbU480D5Vs8xQlJe/+c4ZkgSMXOtdl8HjJjCYFwqJdQ9kuts4mYNoBWY/5lJSievxQG+GWhdP
qHBJMec9FpAELLS7DnUUbzq86VnPzFu/V0pz+YhsxpnYb2MW3i/vI+8W62aUAmge5DNEPC80yC3g
VCxRyC7cqkEhGTnVilgF576OPvLTBUDMMFeUn0e7K2hyvJheCnrMPxCOzjiS9JkFb3KRXlKWaqAj
4UWp8ONNtftakWUBPXh62a1qGavxOHFDxzhoSy+oSWnYRrxG3khuSoiSdfyn/VF80/o18R36U+Pq
q5SxM8oIrliIO67vSx2Ru/xpRP9+O4TyVehVNqG2r+nTc4wpTH29/PmoQ5NSimVzDCDmzl+BRAvC
CAoXOr2WhIX2coL/NROygheIjYt9KhMhHBTaXhR6ir6sShO2DGctk+fvf/xjZmz+kaRKsAc0Y888
KDW/VNVWaz870I4O6xajZLxpYUIdTv9ZEUuSKF5nw9O+kViU2qeKtiXLQNPmCcs3YfrXkvvpEWMf
tA0jfjKpbSicTDWzcIE9fPhtXfRcVXEm3e2GOWrDInjLcxaOuFeNmI6B0aZUXXPBaAw0ha75CZ8A
FV60wj8x8lC2KL/52hOkSSJgX1jTT8jPJpNE+bhWDcRVIJK+B/5oxWkpFfeALZfHPQZFZyhBbmqk
uGAeyGe2sZA6enawXYOmfuF0asfspdKvaCPrybMqPFsTztqwReY6izFk6zg+hdHO1pnoq68f8BcU
kj+gDM3HdXAoGTfUS354orjmgOwvszFG18Inph8rXhGssstKmTR/dYCoN3GRolkmRzG7/ruR6z5Y
vMdp/p8Uy7Xzu9DjPmbynCtFICtv8+98SjcpvtItmFqbbYc5+XwCTvuKZJry6BvHKpkM4Om6/jWr
4buicoJ5EG1sWjI4HXfZLX2aYRScO/ZFno3SGmdxRhXmuN+ph4ZMQ4UKs6qA6s/SFbzVW6WxiwpA
GVqOsae/ra4Y5O5gZY3aQii4wI6hoQCf5CZsaWzBCM2PWirYaCWLThq+JfeV2pznUt+/5yTRW8X2
3zQxYyr2oSt/NOwn2KNRGEvuz3OpoC17Tynaua4NIrMOTNHTJEPwkAHTC0DUeKEYc8m0ZXtOlZgL
eI4u1tHTaWCGkWRmyrGK/LG51WEkKUrDOyOMm9GabB0upIRyhuR8u8FUFWmqlwJpVuoHfZB+eO5/
QSkfwNZANeRUaKxunSOFbR6poBmCUeV5Oh+iRA3HO2oESnSjJs+2B3LjK/UX8t+GHYWF2rK4DSwd
Db7iDF2u8tfVvgZCzVQ2HNPWbcwnt4Wkcj/R9XK5MlWKC/5ygrypGi4UMM27xCaz8BRvSPL1vkG1
BH2wjmN9c1iDgxgGy4Sfj19vyh8MeKdeZlePO9xncwe70fFqKYJ4I44byp3Cnlk31f8Zs3pSnMaV
vglZInnOwBl5EPuahb7g76K7OEd0spezvYs/HkvaLy3su4bGA3Tcjy0s9vSN6dpO4bdEm5YAD95z
CEGavyYBt9vZyxUqF+nKg7OnGCJ9NE5VuFS5FfQJUGxY7qcLQgqgoBjbnjvJxpNkQZX7YWq85IAe
Bxi/r9n0aSMe9kOMST+p3FJXdlX/riBEX7h7cS6qw0LYE51kdbc1luWVJdsYKrecSTQvyTEdb8By
0Ru03I68hSBB6/CRUuwfnZkJD4jKhxYCrMJUdLPj4Zs5sOsIXIJ4/LNN4UpoApt8AJ2n3sJh+0ze
Zy9w8ZZ/wvvepCZ+IwlyVhuQ46EerEn7iIfvD01+TQzoj7NRTcU5h0ROMYppvEInK/Rv2A4b/6M/
pSQw+XrVLEYiaKdVvayCyPxYtouWCW8hBIAlpAZvjNdyBLh7SODNsHNP6z/HD80UVMa60kq9FRUt
iUoQM0tLjspLLQScTNWgrhsZuX+MVq6CJOXwq2DiNxsPDLi1OtRY5m6cvcgTiF4v+g+x7xQKBrhw
IGwdCqn7fvupesohJPQUbXuDXv+H4wRuJzrougT3OU4RlWPUVokTKxOZxTETrGkv+kMYtEP7g2ke
+LdtTo1JGsiW7vNh7V/5fmZYcSmLa+7b6IjVnHX8azGGPbV37gaeoWJB15JAhOUBqooXZbzc7GDY
ita/3Y2hFHymOc9sJn4QdXoeCoKNhINs4hOIYmiM9BE1JKvfjlhJMRkadr9o4MiGKAZa14QdAtky
XnbwQrGVIiAVOO1W1QLv6cWSdB+1feVQ+K37g4c8xTaR765euj2GFsFkiigY/j9q61pv7IbgZW9I
F5DrIcdYfnzioCcBPyXEA1rovvEefuYm2F6eR42Cat+JnK889Yp4y9Gp6zz2aQGmYxLosQslIyY0
llmlXXwXWKJGZG0S4qrFauzXbxrJkTOTZMJ8o2zdbXSmaWPxwLWD9uRZ+ojuMdbnCx+pAEzx1Ri2
vgVMHIhFPnKGhG+pRcxsOKVleZ/YNcmeBp8QM9EQ6XMhTxPSmzPhBhuuXDPEJjZKGNJ+sh2aAjfE
Ma57hUmrKFn2ScnyjtxHIzxcHrpMRP7Nrtfmn3ZkcO7KxQhMuODXqosy5Tjz2QuJE3v9TeQExiwa
MqkYnAzrxzMlabExxNuD4mus/OianvxG7MgZOZCH59qKIq3Nzr/pqOWv93FXnDyv/jglC6N02XbZ
NqUrmCgiWB1kOHzKv+WGnKVY1g/zuWGyw8GbmVNjUHAmtKHIBECfykvr0SjZCp2LBeS7mJzEtfNd
UAekWp4YuRYO8UU92bhVOWmKAoBvjUCFsZE8jasIU+fF5t36jL5tkCCtPJWQDQvVUlG6SxsTKSMo
t1MZe8UR65lN2f1WHMzm3igb4eZrUh6c+5c530IywfO6j9b7G2Lw45+nHfHerxUnAFHq0dSbE0xM
Besl8PLOBrcWyrelY+bEXCky9mknhP5UtSP0gkxc98o6A/BdFESrShtv8qDkK+a2IaxJp0D1wtyf
rrHKc1QQFWDmf9ZxbWb7oGi6d2slEHui67l8kBGdlgdomMNt6umiWe7FYM33wIHWAwZxAeHmUDVP
fJyzlMuhCFdv+Z1uyTDLsMIbnQHLtHtxrQBPZxAo6EmluENutryf+qK+MAKcxeCfmHcu0I7hbzOh
SfVsC5fE090+ML13Lv6q+UFATX5w1bhZ6Nlx4a86wBuOHSloGodnGHw3btD7LFJTEwjersyCJ4dt
fsohrzfn6fJVOt4DIYpNcMnK2RgkioNTPP0nEm1nRQ0JXGMc+pQ6x9imrN7WPk6IrcenTFGrA9Fd
0far67NUVq3dkpsJy35XjJVnaRHMmNJ7jIT9HA1JMETa+4KOW38gaKov5JS6OTuTntjqCUjs+1uL
ngVv/jY6elQPI0NMJ9nqUlCcDtcuED6pAIAKZKAI1rLjaAJ2zE7ytEpRz6JcWaazE9TUCNDjxaB9
NvvoFqyfIo33hqSbxb+DWKeImdav2se7mD5hD+zDD6fUywknsDYDwj1TfGDbQqr+ThCg5EZnQxHY
4x+InFhjNbH3rNRMHTsPMZSWWEsTlp+sNaloPHkxo7XW1jO4DCzakzusTtEEwqkFa+NLZ/SklhTE
qhZVbDj2m80q3SqXpjbwYtQqLbMINbRARA6GzfG8ZBhnRJxJ/6XxmsOBvj6R/DCLVMRrnJAE1wFG
oWNKYqC9vvgo6F0vCUUlFwJR+lNPwLZajVr2pv2W0OTkeKOSNmrmvK/rXYyzMitL5U9IDeD5Jpmb
w3gBpnjxZttto2Sl+wQrQR3QunR9bmRA7NjeM8gFKN07BI98NdJeG7qgtgDZfUdzbsqDwC1vKJDi
QuM+ehndPi1vBi6DcERa6++haRNmTpimMkrqWICHrBpXTAlHBlEch/4H5KzAOHx5r1iAW35AgCHN
J+bsffsa1gIuxFr/yntBJ5bSLIOPEBdrnIHSmSPJxg0DYJVNP2ndIyskyOOojZsAdRz/ahL3Y9ez
N9HVr31lRnTmGdCnjTdcm/fkmtRdikH2JdyDcZdqAM7j+eMZRVxCfZyMEYIlGIB3Yrj12FStLE8E
gEaK8D8f2wDWvVkT21BL0tFgzi0FNmZCW6SBSg/notmMp9GfL07aI1qTTd1dFPexGpf6WYfPXd+x
1SEfHiX5TweHDeEfevCiS9Xtuz7ejO9en3MEbvErpxKawWz3EQCkaP8HPeusp5nSMD1EZ97XloFx
T93nxseYvmpnUvIsRcSlnTkfHWow8UUH5uE0PSj63qV938DCiMLnMEI/sEqXYiLLvGCFB7CHzF+Q
eQhIgHtTgR6ToZ4MXStOkqHnea0I2C6iY+itfq6QYm9PWxUQMCjsgzvxsSwkVs9rC6T0eBcHs/UA
ff/k3xQ8WvbgEKDCBIDrcUF/ZdqAPkT5QuoB84VboMh3maYmU31wE0zXgUTT3yLSuYtNzNlYwpPT
gY95rflt90io5x2VS9xTSq7IbiX+RS8m8cPBdG8JFhOAVgPtqXK9jD3H93nkf5OTI5I5nh2vMrAS
fyzdc9MBgyVrKZ+A2fOWXCgVGn7Ux4SMydLLQAMkyNz0w92jXDmZHtDDsQVCwikPbKOFGdYvPuV0
DxX2I82Jok6YEulRT8SpAoIhoA1FH7h39FH0z2D0lGnHAR3GZh5FdrfKj9hqbmpoWo5Byn1fmMe8
AbZaDajKBFovqCH4a978snr1GfAXMTHZcZGoZ4FOVlqlMpJG30fMs9HxJj/akBIg9icLCxC9Uhsz
62UeXdBh/UVJBi2aXv/XCveyfqg0QzX/n7qkM3q5ZBrqrW6V5P4alOgQ4EvHRlSe+f8ifPR85Yqi
Dte/A6qG5FPLCHl9gbL1yIxszXdmFt+1GgsSuOkllRSYDFNpaiMtQAfRFf/CCCXjwGNUMGKDGQDY
reDFP79s5t97infs09tOUqXC3caq1xf1LSED9SYw0lXQ7MrIR8tZs2ZCES9cE4lFxKQ5BML69cwA
47uGHe7IviimO5Cn2OuVdqNuCUp78Rt/N1iUIN8eaED7bmNt6GaVYFt/fR1wcAwyK8c/3O8zGPMZ
7YKFgipQz4DklToZrE/ceF43QkkRecE97YeWkj5s7GCX9hh7HZoZqhJFqqb+oLPgF5kdrtpe7le4
bbIKJpLyXPmB3pFcOZOtO8gZS1dlGuMdBeGQ85uichds8FY5oJ1l/L/A4n6luaG5bVYmvvvE6shJ
DfqK7n7Hl8bkEC/qHvJejOXgi2uC5XCF/rIVpZh/vmfiLNQIDs/PNVHyPZ3rFmIjEZaPRByURQd7
iC638Fl4jTV4VbolcY0V7bHO6m9pQuKySMDeMKqwQICyh0dzWhb6MZwK8TWUiGj3s6dLYyOqbDna
yuGqX1zFU35A7GQ9jAfKBtfYQLuDdzaDje1eivH9JGPwILhwLGCLz62ggj/wcPta5dpKN8WP5Lw3
sMTpJ2YnETlcv+EbtbACjPgXY9++MzTCnAisce/RRWr2UjSiMLxdNHzTzLuWcAAHxrAFL+HhICKg
nW3QB+cvEWNFZizQahetdZ/V6fiqUYjEuSkB+A0UZ7r0zU5mnBmr1XKeuwuiXtV+q8pV7aZXjM3E
D/qE37iAiN81tiRKevalqeTZDazU/0/Fy7bdoU1xG2jlmLl9L7zL+JML23UCiAA8bpuvqEJUqjZZ
laVrpgIqq/IMzVSnqf0NE47Utv2SgNfvnehhZe8t/uRoWJhYqlqV5461ACk1by9JQznF6hOA4jfd
BL/rPrp/uv/tRfXLIY5X8nF1ssfe5EdgRLJU/CEdCuOCNCLmMSVa4zxl+fHhSgKlZJAe6/qlnc3f
bE5LI+E5SYqBTyFM7RzexOIah3uxcm6MZd5INe8KhvO4zZrYXT5OrZ0nZNMBLrxXc06DrDL+LqBF
JYpZVVaYAlkm2SCaJILu8gK/HIEs0eioADkX3mEdf/33cQsoMrTscfeKe7NNuBbqUVaepxZuMI0c
pX3uOoxECQQ6JE4Cg5pXD1aj/fcm89ZG783brcZKmMxU0Y1Ys9GUE1Qgte6flJlA1Mj/PyuDI0cb
OebLkWlvYfY+v1YgDSDmfYN8ZA7kanwhEeatcme/E0YZoS8KJAOZhOr1ctUXd812uiSPB0Agg4sC
ByIOWexWWlZnd5oBIANPTzy7JBhB9wpJMi/uwJE1W4SyUpAwPXaIPe4xECnmGD/EhhvSxudpcZkX
DO85/de6AV9tiv7MfBeeq97V6X74u3x2APbJciLMvg3aaLnYG/Jy374OSQI4Q9ZSgMvKCbw1K2vM
rdU9mrVpZNIga4wpY4PK+5J6hf3OsOKNOuH9NvzDlGfEGRSzGbnSyCwK2NIHqpGhtCKqd07G7Sba
HX1MdiO+xN0xi0bDDNCoIrM21SWrL8AxCDI5YqtGFkv5zC3IEpJ4LdPZhuNxAFGTQ5zPWt3r+nx1
9jxIHq1ozTzahCQHXV4/AUp8u63E3uTWN81MNmDNpiwmZSsJnQoCS9EbGhpWiBIk3h+s1spaLAnx
nnsq511T+760Mid7f8E9KWoXvh8Zke9X5loJbxUfSvzSRlG9A5oWPQSDKtCviwnr8v/hAa2Kvt7o
E3O/oCy0Wt/fa22cLhN3FauzVQgLLwwH0Tf2vML38BdMV6XIxTn9TcxsDm5N6jWh1iZvyerSCYNV
cJTMAH0ah3wcxW7mWkw79ifWZrb9wkcT/5qUUspGxHYWYBP1FnZ1GTBfc6fkLqCVO7jntP92dOCy
mkmXIEgHXZlMy5/MuO/CNuzcCKu2h4UEJb0WtLZhfzi7+gSDEp57vjTTDsVk57KnxNUTLQWAeUKn
eY6woO5A8jCW8gvMILpNP9zYnBVGdMdeCVT37C3XkoO0LnQe/UJEjMOHxzhfOc3IwzsGhGDwqasd
RNH4Z9H5nCwkf22Ft9yH4AdGKEZb9/QQRfg60V+R26SJoH9iMIDVbE+4jyhntHAD00toovdnZl8u
Ci/ihyagi4ZUkYvw1dTN/jIcu3AaR59KjBWspyw7HvJqapuv3t0qRTvG5B0/8v0HbQp9g/bUOb6r
Skdjiaw3m7grYt6EqITzOC0DWXg4o3eSFA3y+YdMz3TO7vfpW5eHxif7Mvzvj5b7PUA37inifud1
SPEb/dtmz1YbMbnXZKytnpUU7rila9AN3M3nhiTSYw/G6CsgIZcCa2ENX2exiZx6gCd2OYk57pfS
0BB8NJ2tEe2ufNopus6fKOrkIm6maAkGZVhYtGwrQY4QzzeKoN3q8nCSJ76fjxiz/LqOszCAsx82
+FMUhSQliGtZfe9rvvI/bwxyy7RCsMHiLf/bexJLMH1Nnbn+nbNWT2H+30BGYrs24DltzHUP2A5G
PK27H07zgQTQ5SrcnXCUNbt5ysLx8BmGZBJ4adCJN/eE7OD2T0pxLkjERWp+zzOPTaKUq77TRopA
nOTiXuQ/jQTlAXWCZ4MLYolM3Jv81Gq80uugCtuL6ppIYP/vVtNQMIbgmxUr14wkxlJr1aBiNnxF
4+TolW2YbcVmTUBt86P+KhJwgXm941ZPZ2wLfYzLRGgn5l+je5tWUPq+kptubJxLI5LxotbDTiO1
ppNImsM8YsE5JN2gH8kzaVDwyg5lQm4BEgGD+EhZeprzO1UCW3HPiJ8Uc1B9ozHxIWfu1Qato5ve
WxFiH8vLT6+DoI8AMGH5Q8ouBW3SvGRCTCgSR8rqFobi5h9iUoWEeoTTy7zJXc/WlAUIv9RNYCUE
DS4WxHrLeTW1ymDw3/yHbD3ZkVnY5wCfHaeM3JcGFz8nJDUPRrdT1673HMthGJRXE+5jVJmXK7t2
Y8ZdUVZyv88/HXjBTTW8tKYjucemINcQg1AB2k0BCWxnFsv7UXzZV6ErTLzUN417uAe62jmW0XV7
3J2wDnjZodm7AcG/5TubgIAQU18trtQH5mSKZA1U7P6CwBnF1KEfDNSM6wMWIyAUN1F5mMKKBf+V
H86Nmr8RBKxjdDuy2eSOjh/zWD/UhkPXWABlNEosMLD7o408mOmbW8mMsP3mUg9VhInAB7yRAzBF
2FUKEH/rZv+qHGOxdqGjlvQrl/d3V7dCjibU0dX/lMWdxLcS4oECHRZI/TqDd9uUWz6EVRJKih0K
uril6Ca/Tm+kcumXDyWkl5sOAV3RiFAilclh4QmkUwbA2l7m1roV0vwDXtEpbRAlKdzznRwMrasY
mg3/tuw/NjuvEE/9NHcxWsa1ZSyi2flWP3ROELaKBzBftqpH10wEs1vbRc6rQxcW9H4bn8a//7mq
aScFltCF5y0WBIsvI2nlJkc1P+uv3NFaYkd3UWhkOaA+F9pECzuidExOS2EsF4niLSmz8fr/jLHo
SBXHSGnVCfYdRBX1P4Oza/CbpZ38tMAVGtS2nbTpyHHrqdmXEqmLaadzGakyFa4YZe6siAj2iKZs
GpqRqhXztwMw/w2ukqerQHt083fxQPuIogiLaM5AGYKH+tT9L1TtzBgYw9ENAENUt+kYMgsZxyKn
UODy64+CfvHfj5lJYitH4a69gtSAARyk1bLfL10+WZyPXxt6WQvixsctmFSezmJCtPCLigZYfJrM
CZxW9y/m9ZCxi0IjQ2zWl7LZtvkTl75IN2z80gFHOQqOAMbdIf73QDYb+nbRGnvy6wjcuSt05BgH
HdKUsttGWPWomj8i++fiPSnKvQSv+d5V4I6UuXpRPEp7pWhRDZ7PFUvnXG5Y92He3QHfS0+uB4n9
nyKRsr3JCb7zatVrpj+nRu809e3TuoErxOhmsFZqdI+zu9jAnNyrng1XmwVyBgyKrds5QjSuDewI
z6uLlQ8jGxUPBGWlUn5A+lAOWw/1lPLNJnIGuvP4PysyE1/cmtIkp2cL7D5tV9DcviP1Psu9/hEa
JInbDzKhtysNJuc+obpSRAp99yZPgNy+P59Z+PFCsXlV7CQYqvpz7xiGPsn2y7+TDouXLiXqq9eZ
Dp+0BU/ZWyGiCuzC65yVC86YjR3K78y08Cl57Jx25M+i7NxO7f/uXeE2QMKolBLTa48G0oDF5bcs
Wt6j/Orp5RIVz99knHCTQFs+yEpp343FCrjVJLv4slrfZW6wgzgMsqq+d4XyAjfw8cXoMmLCup46
YHIOXGQhgKb7tP23Dz0/+B1cRcEPZpmYuygfrgYQ5/atG902gJZv3Mo14zirDe2PVwBJekuQXHYz
ctBW+brgA2zQUsiZB/f5k7fW5eKXXQi2A6ucj5i5hTuypI7jdYFA5q6RNDkHo2iyXg2rGp8O7fbr
QOqrOZyhd8xoMx1LTtA8ittbeprUUUsc7SZc7CghZfxjSqAUeAmhEmgHjOtinww2F4zcMH79jDC2
xO3mvwfaQT+n4TV4XOhZqtcU4Ock1rU53MSZCxrRyzDGCRE79tsv9G8qZFwvNTE/d5VXqXjkM2Ep
0PJh2JLrn7j6TQth9M1RfOyh+T5UOM4pVBhQIPjV15T4Bb9TAykcr1vf/cN5FvFkrltGaLa8j+RE
IPiiddSKNInFhuNr0iNGcL+zXBhEFMczRAJKShwyKMpAnHhz2loAK73oD91bJO8uX1836KgfdA4j
JE64efg8iOA/tvUMAFBPi40/UP0Oau+Qql+qSn3b5XX/dvgecZ13vnF0aSL3Vs7vWfPwgRdymnPN
Snp5ZbQHUMe3Qk2Be+ZieUT3vK+Egk05eep6E/ahlO/G5wv7ml4kRZ+7r+GKNT1KUpFTUlw4deya
tl5SYGGWtsVI8Q5i1MAAd4ZwFDiMO2mJuneHtx8FIN2NM3/y4pKMR3IRnqRvVz2UZu76rio3zcj+
Cx7ae6CJ7RN68hYAdJhgo065fxomPl5R8XCSH34ycItEoABlCv5oQXdMKJwvKyz3CsTNS2VZNqqZ
o+ROBaJsxArAJgPm9DLpkzexTwfwrwe4SpRQjm06wpoAniY/GKsGUdHjeuGImEuL9rUIJMwPyDj8
CGX9OHXUINCyFhLjr1QVz+R3dEZ7RfmrbQHim6psFaHthU1y1rcuJyiM5q3iaHcGowLfkQ/lXPGW
gvL4EwK+W42XZK8xLMohVQjHbbfoN5GYRBKpPVKzBKdco3NXizdgQxrGHvDEtTN904Gw/sXFiuJA
pkSYWAAIlcL4hWgAJLWUKb/1+5hpXKupk8xiXIsae//bRww4sW2jc9MRMS+CTMVwKiFNOXujkeKv
/gx+nDnB79Uk1UxYuj/tKP12ssOAwwJ3FBBRBvP0KMI4wfVeF41w5DoShQuhv3KhZInkVG3H6hWc
Y/oOShGnzSljLnkttE+ewwEsUEVBG5QXotAxHh2xlh0TngzoufEydU1dtqs7Uw/ukL57P9WRPrUT
Uge0u1/0sQ60KpfZmZpV5GC8o9Zowpt+KWaAtT+T/37djJxwgUVk1mPejBCs8u87QH9w/FeClJyk
KznRnJtVmA3GKwAJtrtkkf4qPr0JZ0851YOkSNwsufoVNNtRb1qyTuXAqCb50NfuRvmZqYPJJLBX
j71ZKRzAbE+nIDgrdoWGV+DQauOxeyNy+AjeiuTWAJ9/eypzXE/1kLqULpg94nY94mseP8pfJW+B
0uE6u4+Vhgt9wb2eAvNKFmlLa4y5nQT4sVKupy/NhLrEFtACpTqsvLPHA1x78LISUBrwBok+efM7
MVyWxwZK7gI1NshU76R5Q7FC6mGqDQz3D+G4qwXAxN+NZavjpvj6+QovYejsIMRrm0hLQgx1Sno/
8GXWPKfm2V813mjG2FH3h3bupb+8zsI5pmvx+mHul+647iHwTBENnBHDPAf14gpZllc2lx94E8G5
vxlhY5VM/ZdZKkswULg2Sj+63TrSIlV75ZZi+ACEu7rquuU+yxww4/+zCmZI5r0j9ZbvvOyNaDb7
m1iE5oYz0/MF6BXUw+JXoNsPnK3YK4VPhWeYhayaNiXp8nrCJK+8RFeeGhUm1HO+OdIHpd34xTZq
X9pfJuWn4+Cc1uMpwyf65hzNYdO01JcQWn4DU0e/Q+Z+lSMoG4b7kgVWZEHYLEX3YHBoS+mye9ds
nu1uwV073dmXQrsUULLTS9PYsqpMowqMbtFaVZepGyRRPB6IkIDIU1wpqwKNlp1MIZjND0Idztvk
5iSIQ5lnz6FTzAKxKXv8JlNEuNBi1R0Kjy4jAm9+yElKwG3f62/gTUb3nrNSxMeY8nNPR9S/qIiL
bOJIB1JgR2mYUulH6QWCLy95CYFcZNEIWH3HjyjP3hQQKSmnrNV7iC8jAr0ArMd02A9sQtvTR+O9
UU7qTfBI3e5FHsrBEmaggl+xMcvNU+mhCllCFcsViCQ/a+BWrByzf2RBTGjLyJJcY2JQIwdZe8yE
2mXgFnzvuUvzQgTfGmFgEHi6J7mKwYQW5qN3Usi9Ity1mo8JobbfpN3BiAxI8R9mgRSysbMuQowj
8fgWCQDIRdfxA285f+EmkvyxpVj2zNthPDFKXKzY4f4Lhs+bKToU+i5ZAxblrr5C5sAt9McC52Aj
a3W7TQ6im0rEBU4oWjuYmB5cxL5zdV8sIdSgAsOzjdLlkL8H3IgCaDoTxXegufle3y8GE0LWiBN6
Zo23sGZ2G/zN4AVaOW8dmjPZi1tuAqglZWU/EuQRieadTXC6+dowwQ47rn+uCUdknHd7Nt7jXH2N
kchC5SNL/AujOxfh1j7DH/BiXPOSB53phaztR3X/7WgNfC3nJAKQMdnjoLHo4xO6eo4o7wd7BCe4
NWqbwkJ8PImLpwk2kTXjW3ZBcp7l6yYJEAOjHk+n0K0dmGjIMEAY05M03lxFwRb88oAuLpXqCLXy
Td8NxVbWq9ZpwyCoW1aKNGzbuFL02QAzTdrxbV2kx9xllSBA6kTlc8SZKTIr/iRUpIjWkF0GxUx8
3NyK/40rsHkmjvXNYXHlWCD9USy88Jqf8GdF4FH7tQE+RHY5MAXHgVY13fbu19DqbVusBzV5yiH9
w2EpMxsTuXW9sXiYgqFbwgbbc4WpKC9APEHDcswiTqyhA+IRlcDUxUDl5lVvaG8FC4h/K3LeAVYd
GS+FjCsL/izDzgKaHMPh5PisuyHgfew6aijt0yxhCesdf2DBJy9EfBdtwXha17a1qxJrKbpUTs+O
jo0y57d00+SXWJyKZZQiQSrPFsxe3h548ew1dAzX/d+cU36WP7Em18iTDBw1GFzYc0OBiv+aXrIN
mJf9atclWVQ5Fvt+MzzjvjHDpHlxu/zkPgL58o+G1j3pVBC/cfeF2Qi/7FDmiFvOEUerfWbm36F+
LXAMu9+ulSl84Wr+i2HxJJ2YRlXn3ga+Xad+Lph0o3NBkmIweg8cbZBRXeG5M+jPtgpNFMTWxClQ
N7Wi0idcPy99WX+4EQrn646h9h/ubsjt2vebyu/gTekhCE1nnoB4O+jRrQ0mnrMrP30jvVqcL6Lg
a/6NDXqrcpOuzurHZSJIrv4UBcKnVpEdfNk/1MLPd69Yx4ZQKB4r/j7pD9dA9ugbQhSloR43miv0
o3pB07yVcETl0UhwJvnsR5JxF4JLYrrDCk/ohtBxIPADbiugYGXEylof49JONAaMnRzahsUIYK51
OPT6YSf5k7pa3lIhm6LJ02AjOq/4b0F+g8pi13JZkQ1IxzBnbd7gcWSR3GFeJ6WLXdfFcah6AVmO
9cR8gdqV0BlmyJZtuTSBxd23uaqrBIog117N5RitSffthyaloKeisOR7w8QegYfmRMGEbNm5yfjp
0KTVM7oQ33U4i1UEuubJ/oa+amNj9NccJdjnBEYwtKCNGqpEp7G9iXZiyjCAocA9CjfsIMMKRMc+
mOdmvxc+Vs3uKQmrzSslzzDbIcD4h0sPcaBtNtcy6LjL2vsDYKz+cVylo48IN6Uo6RWZJcaCfeqT
w5GD2/tM0vuOY0u/Iuo3zZbwHAZ1OnS333tr+7Tm9znFeCrirCbH8wX0SfvPcJNCGXDDF0FUcXLY
PB/nAFYMirwTfuTSoLC/NEnWGg56QY0nLvMP6SLtAAAcvTBGhI/w4hyaq5hkoQEwYGiaSe9wxqS7
311ntN1oq967zgcrQ1IBZeLUEV10p6Bm7UTCQDUAtUJidO+zMxmh7SZGHEU3bD3A4qJCniAap6FU
XnPA0npb7K8H8rD4NI/XLFT9U6+gYOjPf0KfkjicDu92tooysG0/+xEI0HNaOcX4KdvXLE+HeiIO
gGAoJ3gmIwdTucoh5Rq20foBW9nd5TZFGtNN5zSkXZJdkX9PrXXHC3+kQ2ERv+oste1JVRXZqCmt
KyGOkwXVQHbkyXBgS7zoLbgZUlu3ERrHJgJNa5rzrxeSkVCRZ6n0qqTEswY8T5zj5slQ+97cBP9H
HSb7L8vtDB++zK0dML2uHIt/p0wOK0SUEHCsYEMNDuW8DoqO/h6Hz5maiApDa/Q4rsq5hx60ZCu8
WZ/K/GOTWIBD0dXF19os+Gez8OAgklOv9o9jrvN95Iv+IkPMHmLG//FeFWcvRTaO5VkctVz6ygnw
0pPOdbr4vskP4Pt7faOPK9SMikKDilKxJZQawPeHIcLiNKaYLCCsCe3BUM2lsHOofjB+SeYOZ/7O
8FHIy13g5AuoKkhEzzuHYzlhIkgdHaPX01XPo8I4smFu0Udn6Yn/UwE/fAT0DyrVprwvZyOI54/w
RrWmjewFt58vDx6FoLz+3xQZ993CgVwoZmasDA+7JzpLjvV23aC3MV4gwA5epfVOxIgMW2YW1XjM
Ad0joSPkOKHVdN3fRnurV+bn51LZ60pRbFjjhzSJ+J7pE2NCIY3dZWKUJMOSZpArC3wOEd2o0ZHX
7KG7HKcwR3ugQK20iChC/tKms6dSAd3rubH7CJafAbrO3ed94YeIsXC2/iIeNXIYhXz2BcyFIyhF
e+b4IPuCsFZw04n8Tney6UKi2+bywaSZL6HB5ze3NyMTRBq//QH8uhR+zEg502isWahLwpdY9Y7k
bStfZsnAFkyTu8PslmGFvNDDE8e728UazMVuqzUJBkffmC/TOemHvmBji21rK6FECLei6OGLNwDN
i/SaQkZEEpIv2QHN02kZMsFLh26ohsRO185GxWN0G1Q9OB2Y4ky/KoaNfWkQ8r7DywlEz31fnpNq
KIWRmNcQ4uo+q6QBksj4S1hg0EJqTDjP0oO9OYl7RfZ3cLuFs7v1QhpzoD6DuTGTk92Gp3pFtoEy
K7XHfTs41dmJhWHqGqoK99xZ2SRSOWlBrjYVf+QK2dvLp0dCuISrduvl00hMADCzOG2hjX03hYCh
rh6VUsGWuqd8In649x1EviIuyDV5xwg01Pd5korBTk4u6OUuHPb3GcOLWieca2yZsN3iUpMxlzjr
BIaKUFIoz6pPC3q6pT29ZpEr06tMVRne3gHdNRLXl8oQbA3q/UIdVO18o/hV7z5VXfU8o8clGHvF
ydlpaQS9wWmxcRrjhbjQ8eu6BI7SI7n97pUMZkDBY+uNwykbt2wlaRUp0/De6NioEjMJt3+UMSAn
kpzjZKVFi4NE5dC3Y7afGvR/8nWqDs7hGwmtVDFA3qFZpJD9tPTZhaCMhyM+0jc3PhquEDQjT2R4
06yPrZbYGu/dFyqgdfrklaP4RjxtvH0+1vAlS5TaNtWeflztmUrcZi6XmvAscZsY7icF0x80v2oz
Vmj/rpl9QS5Nxtn57+Y31cgGN7RbpyZxlPwUGntbJ3QZAdxA56DP15e6QjaW7HXibuvPMdMb3Gvy
s5GMwRB2ZXpgHMnyvoRO51BKFAEDgsDJ/0MfNNWJdpn5viexg+Sx15/8WUi3ZKPO58qqIgz/BnBT
gjR0g8X8q9vXqcSjj2+fRdu8t/NqQQUoOpbCFYTclgaW3DRN/AQtZW71r2EMBam3M6OR4p4imimL
52ue7cR3bGHfbhVPOTEQErzhSZ2urtAW7m1m0o5+MRURAdsv0SKW1DkCrME3Kyy+ygg4awrTe50G
1sjqkJJX79cpKesZ8gGV228hKUcSiV8MkPIpLtUae6O9tclMR2ShQRap76/Esq6nj3ypZ+o+RvRj
Jqcl00az7dsLwuPFYsPkT8UICh5YX7wH3XH9AdtISEOuVAeY5A8dWayrE0J49AK2ch/o31/fHfHU
0NQ/wD5RkHNUqI+2tAvMHg04dk3PCE6NKWaPvH0dkhPFwItqvgeZSRAB218yeCVncj48t8LAJ4e5
mnMb997yhCum6/cjL1Nl0LUEB+3Z6NWIjJfvYEUned9tASqFK9rd7wU1Oj0k4H4VtWRlxQiODmua
+JTdj5wq3o04Oe5YXWVHCvytKKHegBxgwvKE8y5hMlhUNrEkuqBAG+Qj/Omb7yJ29gNmcbK6+pOr
lTuu0jGwc5yBgFOJHylm3WscrLjAX+uw9YoxRyvtU+eUbJLc5W442HEVHH45v+NS0m8gjRip3i3l
h72QpJEr/ajBAAT64PsOLLg3cFpYLyKyW9UaWwEcW7SGlQr+/HOU8K8imJRyK/oIB9Ipnja04x+J
XeFwzQYwRsd5SThzEVgxM1fOKcLKO6igtcv7ESw5FXn4Bc1DJ4MMRlM+V7MP6R70+B+zescJKRek
u4lRDAutkJo25Ltv+UYk9ou6Y/muHqxQG/eUpWV7C2uh0uSV80koNipVfUP3cE3x8YzuTyMvKNBx
YuiCQIzO6sRrV+v2knkgxXDS/46KqsqSzgLlczT8OcIVY9awLRspz72qfnGUfQAzAGqdeJQMtfG7
64G6rJs3lsWIPx+cc4Vm4g5LD5ES0EAEr0tQ6FAOMaMyqlgph2P3H3SYCnSXcZTdcvx/yFJdsX/E
4fTVXNfYwPLVBdEryU33Wqmaf1uO9JZTZUtMWMwGk8sw557GzLrR3GB1QNRyyuCscU9vIK9LIXjz
/6biQe5/ijtrLkFzwYQpQtykWvEmij0zkdi89ViebFdAHAEssVl6xnf3VKIUBJ9AUtqsIVPn+Qud
+i+zR+wknebRffpT5x0X/myDANtgGPnrHx27+LWviTkqB+So3x2Ioi5WpBAOF9Tt1CbRZ0kJrsWX
0DvVEQJN97urqCx1HiZ67EwOT3Iguu8OnHE/zaaOCsltQzNp2oblKq3dmZoG7eGss2Oxx0T+4ckR
kNJfArFSXlA54nSc/S0xP0BqWIUfp9MQsOmWHNCZhapiMeCqamkY69fO/nwxKG8Bjs75k0Eu4wOx
58QKGUfwWZB1RcWAaw/EwP29AfthbT0UGi0qN+OFZRLObch754Cl3zxVw87wm8kZwtKBwbkMoDwL
Rv7/YHgEHkcZQLKtWkYigfWlQwOG+TZPwIYlAvWUPDft6UbZBv6SQVcI4sPAC1StQ47aPqWNhkSc
AcSHGmLZJdCFikLg/KWpwxu0ue0r1x3SeZGH18KadVhD5SIwlkAb4PmV12F9GZ4kh8jxvX+RjMn9
fxpVP4UKAglDGOe8EybOLghGaEUKe2Z3eHYZs7wIBVtKQ+blzkkFS73zgszQ0AO+HezSSMzDEcKQ
DzHULiK7slvZRBYkJAYL7Vy0X+RvVIZ1mjfQHZJ0aLMD1i3EMTlaGPNYpnEjIlnW5uunvncGXcoU
TRh0hREfDko10gcI58a9szaRk9UcoASOxlgQWDev8HtFf43pcLWcH6wwTHlTRuoSdZZF6us9Bq8W
j0H9wOvAP9BpQi4fYdiEHZ6NoxHyYhzZ/MJWtO0po+wP1t+ejs6kjlmfQ+vgkrBOkuxG4k0qDyF+
eT9Uc2FYP180rQP0cOVWN6t5HjuVWCDtO88zXBElMBatu++Ll8ODySPv/BtnkvTmqw953OJRhMB0
8aqftT34jZPW5ER1HSXZAPBpDxSn+wzZOyxF/xUnj5SqOln8vYvs3y2CRPIRKc46Pk2ntnMdKWYO
jUSoFIqTHIYXgKptqqYLdwrYIy1yjTB6SjyZsnlyo34iHifuxkL/s4FQvvjC8S312wAMD9/56BYI
wS+hHwm46AGlfIMzAFndjF+ZbVeryY0SYZc+3t1DDYwMm/+qaUMbArdvDHlbUhzZlKFBY1V0OiYg
N/K5viPKI6SoXrfLSNv7NGA4zUrl9BMNKTBoJ6rzVKwGqzYWkYcNDa5+5ZLEoHXa7fK24lwlF7Rb
c/SxWGBEK3ihKIXMyh10jlEz7C9ZNDMU8cc0Zm0YeFPQMNBfnASLhg/+uL//5cNKBOknXUiOiuu1
Qtva0mUZfdw8NVYH1keHEK161dJzShmJbVNTl/WCKa/8lQlPVmFx1eCEMgNtxnXHVOZ3vs0Udvgh
TfDcYKAlrLc7+2TT3M6Q+WTzvQlu2qXvZSeeLX71iGl6B2dIHdFZLY2ofMiNorwL+uxtoOlZmkYl
8fn0SimLpDusjT5gbliR6T43wI+zQsrDOlxhQF5GN4q7q3fb/ZbddY7C3s0026ZWS7nTLkFZchQW
6M2d59Wd0UbZAIJ9G5GVBoDCuD9oKEueFNcJmAKkqJ9g1PdKIqSlF55nHqC/jbO3mGKIwhKozM4E
ph9KIgK4YE1dmIHSSv8mKQIACok5f9/Zx1WzOmoBdOPQNZL0srIJrsFOO9BN3jO+3pdodmaZ6/IJ
yzXOxcGbKzJ79UAE1V6tgUhBchue5vQk0ZlvuC5pJMOPA4jHZw0LuDi06D0dbDSm0TE6O+6CZFkW
36NkxUK0edICBzH+FICuBFpmYQBwOcXDAPb/XsrjH4aDUftAlY0bwRiQohlcXLE4sUD1ueJTNdW2
SYaz+kbVjmIUKjN/ne7oYjFMGLBuZHiKiXor6W20rK8Y7GtqAKeJyP+nn9ML36MgaUhgtrMS3Czf
dngmdC8f8qjdsNZG0z8JiK72zwyRYeemwNMJ2mVkHZpWVFHzKfBY/TZs/LaUFLeB2isQCE4KAbto
7qySCTxb+Oah1LAENxjrLpCiYLiCTS4ZavIAidNfbO8AUIhddhri5ymxRV9nEkRz6oFOo+T5rJTG
AmaO0mDP9gm3sad3197smOy28ymn+Jxw7ATECAOtjnYAl/Fn8mH8y/9IHbGOgMhaYnBdEG7GaLps
VFSWIEXlKXTE5Y9TW/w0BVbdcAtiKsSV5xOJX4odFRqqWNw4o5W874eutKbVu06MXsJHs7m46sJL
PhD3pasatprLiQ1QnvaILfHOFRliFpSh/VG1fy2x4SjMi7l6ghVX7KbQyg0NFUep3r4G5q+gE0HA
fayZCGrXtXPECxRF7ZjbBze70oEGby80rHg8CghDlXBg07rqOR44X8WNoMurz00NQKgHMl9Zt+yd
tF7RUxcv2UFh2tPrCBxv8mGUKQMUJHoBSVaZPO7y0iDvaJm12gF79cyHiRlKXvSS6N0ciUYnU9PT
5PIUKXgUzeevMMtd4Ot/NqRREdewRgNiy48T/3AXD/ZSqgp0FeLFY+0sfVAutkFyHGAmXJgW+tOh
tNIw3+gGRbiTcdoBh+jc6Tql4e/9oTQLVcX1XoCa/fB2/Ma5r9s2lh9LcyHbMb2ukOoWdS9Ie/O/
xTUML8fqIefDdiA0ooan78k9BmwagWo6I5nUgk+bzsemTJFGUD87MNp43HIGDF9tPzkL6zgqR9Gh
fWgryIR4zXa42WHBPkqBahlZ/JgSmu8QU0DCTPbxOaUhjzXZb09V0wAotlsNB+tiKPN0/YO4+q5f
v7WoafIjX1/OHn2hk3rsrtfQrycbfexnbBsfZC2flT2k11myXWJnXAFB0lUoi+P4myzaq8g07+sK
Oz8/Sk6NXkh4K1G8Z/zoHBFkhL9G+EgYnxh/VvZm8lckSA8qrdPSih3+HKPIfYky271GCbScvWFc
2vou5FVsj80Zr9r3YW6idzJY1ZhLQbSIpZRa25CcHgvq00cBhmqw0PTA2bmkidx5c8M3S7hJev0s
xvQSfFl1J+a4owiGy96Db+Ixa9oKMTk89uGCJWcKQm2pEcoiE5ZBntAnUkn+CXfLP2fSCDOL3tBU
zdGE3DPlNsqsKLdgn9SxbR4lop+wuLmyEwmHK97G7/oL0PyUmMakri8+AxR4epzRo456Kz32SEeN
tYEdMmk5GHtJolSdWP83J6T7KQcw9/CoQFGgwXOqJEp/7KvS5ZTE2hF0pgfMhJJGW+bTlRWmgL5b
zhvWzDJWTd8SfETUQ3fYeYW8VckZy6Eyy42cX0RPh6l7c8OARQVpVC+RkgmaubM/lFvYJt3wtqRf
oPcqfU1UwqbHafurmnIUAQk0h0R8N0gQ726RnA7qtd7ELF0lIYCd0/mXcP/G4arhPc2RQKb7wk63
NOjny4MXqIUz6zG/MfaJxo990ERUSjdVIUNX6GB7ffQjjwXdzzuVEA4P04U3+bmpAeVkE2D8qn9U
Se4y0F/JNH7hYlJVt0Q+cQqhlKAXCQr+BwVTYGspHk7fVyaomWv9k4Kl5EFffmMKjJGsfXczQVdI
IKVM+3sx7WAC81fWBxJXHbtK2rbWsozYfWPoYpIXqxn9Moh5ub5X7PFSF9oFgGVIrxB41ZFICOfJ
tvhqLi9NhVIsnkoqVLUv3nUj4YeU3mCuEaGoqcSQM5iKUR/8lhkCWTFXfk43MQsbodqFCaHxuPuB
+uYWkbkIvLEj4VSLJ7BgHDha/OwKqW96uiqsMyvDw2VKdPwXDWVnjUtkv7huxoqTb5OXg/kF1Tv+
MCyJBSGcZHpSAOdPm32GGhkwCaN3BA/iS9ZgMF+ltFCXx/eypqZ+guokDKCcaZyWGM++q7GKA5ck
188HHBbMntmtWPDuqkgZ/DlirCu+JRVra3if7OJxEbd/4mWqMk2Jiig2Mzyuo+X27QSiOPsic+6m
KThJoJlnVb09Z2rV5ioJNqg7v9gOBLF0id8N+MIw4S2EbvQwlvgkeO2Nv44/BQ1QgvwGtfM0rNjP
ZEXxpq/Tzz2BxDD3BaGO6IT0KV5ON5uRxdN8iFXEoZzG1YyvV4EGNhil40SpDZeweZhZ53zkrnMf
TnrNlCUpzhMzmNkU1aqIQmLvNbvbORIOc8Gd6cZv36EQgJMgii9gpnp0+bzI/mhNqwksMKSwEBz2
FuEgUUS659oepMetRe05+LJr5LmA2/vueb297ZB2qI5iP0W16UyDKywbdw1BiWQqzFLoyZqgAdSy
jb4VBA3V0/qWZss3evr7FvECAfg5XmfVI3H2lysQ83OMnxlAhyg48zaRY9T+X/1CZKBX/dqLmuyk
MwDF3eAsXIiEduD5IJeido4MP7Lx838d+WVOVM8/yYOiZxWcTVQYiI/Yr5OxEtN80j+M3RtjEbt3
V+9BWxRAw/tc44w7g3NAPbSOWWgeJyohOYR9QuQOGjIlxHem48LLborJb6XsNjgu/u/MjLaFs99M
Hct+dl0H7S+pCtGpq+NHJpMiuMPJdQ5o7hGkSdK8x0xHPZkT/HYcSUEKFmBL7ZO6F8xPItueLfAn
LUpTuqh2F1u5GttdWPSKWERqQdKJqwIN54wjkymFxCJTuLlQWS+yMxrkM6mR+GxzhefgriuChuVE
ZR6H/wPswP8MbCKxByZUezLDm3ada0N2KaVXPdEntITQUYQr8NBNok1dGga/mzZU+loVmhfEIpMu
bcr+DZ3tJZdEMDO4caGdi0CrKDqIgT/iFGg5132o49iG2CvyyqCcGNSuUnNtDv2Q+Vf69UWrNBsS
7s345UZHqgLMEFsmBhJK173JCSo6PdjxEaiTtA+M2z8vVc1Q3Dk0AaFfIK0BOuYzZjVrxR/v21ho
ILti7tMwekWmg3/UIukGWyzzBd4OrmIlvvP4dXHBfrUcQOFx6GLvKg4ZlM+i2ylT7e4dVnvbBkA5
oMH86QQ5x1ehi+kROcZLlehvYPS7kVQb9h6XbVvZo3wURhWp0zXWATafMDzVQCQBX8VHQ/m6mO99
2InoREP75yIW4m9HLVgfl1UqfYWoYpeZEQ0Qv2qhUMcBdQiKjcTGja0sibvqSLvJTRbl+Wr4Srie
aRlKI0GyrSgw7uHOYMa+1aBKJoeZmQOetd5nZMk8S6VEk0cGD27hiv/cPX8eFTdf0lnHPNonEx2M
WeB/Xz/hAZK0EVZKlq+Da337/IaEu5MzcAkSn6ZLiNN5ifItnZMIBkefItokM2f/kMs9+N2xQ57V
WHTqGhaZGC7/DuLpioVsOnctVdEs0FZdlh025LVAVYcnuhKjFfvdaVOo+v2rXeHqWLNEmyq2X86A
LMLgcKI4Tn+KOcFnMzNj4kjEGp+1TrwzD27bt0X9hc56/shCnQE7skRGIblldAbppYaOG5rT9tJl
HvoIWSiO2AvfzH67QJfpf+sm6rJ4uGmWM/fPyFmhMS4TuutcBA0eZq1bP/mbhRpWU0DhqI3iaHcZ
YGmaInUNVzT/yT3PEEUMw8ijGLCwGqEa0I+YULJy2eauW+tONi1SAYWvWuVuAQdHkhFAz9XRUwuF
tnLKijLJ6RbHNNkBTN6tsuf1RIbSthPz1R5CSMezlYcAeHWWxbTW3l68jbLhe+Rf7GBq+ZajfN5p
c8yg6RfNuGvW4hbW6GOaYNKoEzeXMQR4dNhYO1IZAIKSGHjIkB/fN2hr/MwMQhvCCWS4YAICYn71
FEFLmpvmHVMQExUWG4IHZXgBf5njbIwGu2xeDyRbEu1NQ1KbItr+Uc96Z+iR34UhIngdVsl19cPE
XH7eBRHNe1tiHhOeRF82eMq34UFn5fn99a3uoQ5UlqSfDDfa9Dw95/XKV8i7RJwh15AN+xObCDre
F/R8A4oJ+RHTl5Z52Uyc/lyZlaVni0uAH2aHOaQ78WtRHbPasCHuNSpN3EESoQz2tkzm1xnvk6ab
xEbSzpTdhNgQ7A9cwM/e1ow49zg98YY2R/OM69woBmKKE/oNnXy4Eo3/gN3L+5BifRYjSwCvBV+K
nhevXfnRbuyiLx177gjNlOLDwwX7/JQsqeSzU9/fI0dmk2yK/Ss6BosF0DFZ+TohZzcSSQWfW6jI
WKVGDnl8ROdqzTGrBUDZUghcFOyiQ/NvuoUPkm3wGDQbI3FbrW3WHbpImwgVvv9mNIHoHo/Xmk+d
O4xlxvJpufZFphJlC7EInsQ1MnyOiG8B3obNWpsbPio+qzgXYB1xoTpzt/E4PXRfz5HJUiQ6IXHK
Bjo5F3ezMJ0o4VDrgwIPrRMCXuxkTsCat9RjwIZheridsX4Yipi+JKNpOu23doNMgX05eoLcCR1N
jes/jYhTorkupw7HG1rSoqzdpbFa7drHliXpLju/Jj99gk2fF0cB+ReEZ9bN9oeWasVh1LYEiiMH
8r+8n2HuyMt5PFQ5JA64pUMgAGMs7Zq+dJh9lc7sqcxQFx0zLLBqwF1mbPnNl9xhZTvOrd9NLB59
000ttFDgGjsXMmwR/PqEL/DvnOD3+v4g2S5ENVQ4roA59CPCOOrDo3oNvFOM7g26CWNGFrU3JOzr
nCAd1CJdjRS/84dD8G6U+s/ckJJ8zlezY1pHVS6bZAwfRWtpmYlr3p3HK/NEok4qc6kEYu7WQWv8
UqWD9Dqwl7t60sP7PuxQxdj71qg23SvAXQBtdmFgY5cqCPMx8RgTGFDwLC0fekjNfju5MChNMr9O
OMUCYMenWuEHRIRWx1sgpPfCYmJFdQrV/DBCUaAKK9sOK3KlqsmDZgM/ItecAyO8J+3l10M4EGkM
Xo4hhdD8HXYIhDsaaWuavjWfCBhOrliUBULx5JXRSkQpwMoLxXOhBTo4Q7dUTv8CT86W4y/OqhXI
6/+muj12Z6dNITLtzv9fxyGrtRW4M/S/zQq+GCSEZhsnm3JR3NPYYvsJsjwTCJiSYFhxqNQxViHO
MdH34keGjpJmM1X2+dlrVCt3bdTyWodL6Os2lnPTe0UbrD6ZpUTbMWCTLnYqh/P3Rai0q4XcpIbP
VCbqw6opjOUabt4D+bJd4hsGlRneEqyjSJyScCnCa+p7rSj72wiOYvfknqaO39XRdbuZvBMKusaF
9tHhRdUbLUPIXiqkYX009OdNqvq50Cjm1N7eO+N+UEcRWzj7tb028wz/3GtwXqHbJP35B9NBtnol
Mnva7wvfKljFYKC96WKEsTbxubFyUjIS5jwrS9CwVy5TGrTyOKxxk5/sIxglNWdASqFbaLyL5mYR
Q2XWS0jS3fMSVde3T/17pQPuRPdlwTqtiTPge6gA8uLzcpBoyIpSzQndLO5n56IW2x/HUnsNbvPn
sgKj5K3D3hZKb9byHmRUZatOnN1m70mcYpr432xwVHTsNqrON8EF8jh95gvR1W9O13K0Nk5nt8v2
axLc86IchPty8OpNz3DNPM7YQV9lyrYfqxgQtDcG0OUfyygafSVXNWPx4KfltG6AfwzrJdJylsWx
V+J0I9W39mlFtVAq0PtDjkYGBAHDhBtiPYDbOHHXVNU8iLnr3v6b4/LLHem8EFLSHe3xzD5QY8G7
/JQhgGhOuT8nBB/MlrdXhQE/ZzUx2MQb/5xdHHRr+n2HRJS5ZYrB6nV5IHYF8PqQqQNNW/pQNVqs
kpTWbRDjwfa8PXrY4FsKJtEGvqFskoiVY34bdfcvd9xFIkpV/fWUaHGufHUIER8Buz2l6wgpsf93
NvtTfIsgb2CuLd8GHIbGjMFs/2RL04v9h73o+H0Q/5q9CaZ4g4clzGzQfdosmDTnGDhLrC5zukl4
FLyj45agY4GN/wOpuP26PtH/qhJ4hamySDHi2TFStiJ0ta75W8eR7Pp2Lfe1XP0zd7M7K6wf4Tj+
EzcejlOBrEiyHAiX8CzBfaFvIgAFsHh5cu5hr6N0zImTyCoW2haCHEaprRa74Qt6xhNs/8XCJjzb
Fug78LA7tkb2vYOBsYRMBE9pDtL85m/dIJx1DqAwbHj14FquAlNMEiy3DbPm/kms7YNgc6HIK4c+
pR4JjWicXVnUP0IsZdhN3x5hwvhcU+0ddktCYIkgt7vMHn7k1/jyxH/yCC2XqZzv1rkim5Zo/tn6
LqU4QfrkIT5sJ/9GOuWoCYgKxjgvELd67br1uD0Nrkq0rGX4BmXd350cRWsSB6w46QV+yWEaiF8X
B0gyb8dcDMhYzWm2Dv2HHx26r1Mg6eV1BZhkRuK8ncZW0iWa6fzaBqIByefzIrXzlOrvq7/rN3mL
Qfqu4ZP/Nns1CsfzpwVUKMepNJ4bWVtSsD05wdkOofkO0MWbjKwpJN7G4G2vaayrqMOa7uTG+yY2
zJAwXmV8iYtvT5FAvww4Z8PkFHXiAiM+KVZDmy5XdYZKh3Az5plcrkUugpXo301SyXgGuuOLZAcn
ERTRwoEkYh2fycBQPgcQ01QDKo3x3EXNLYv8w6HOJDBWfQIjQLmXJtedjGISpWsPyVWS+ja6Vm5k
ZaVuFraKqR4a3duX/a6IPl2cMXU9LBqtcMY8ZKatvycPEhfUjuZVZObQ3AOfAxMNL4ePb1C6edUy
cQxu/u3X0AjsioDXXlXCi5Tj7+28ndf794NPumDb1hqVPWfr272+u87P3reA/deFkBI9Obzn9wzm
gumXZEhD8UT3bO4Ql4BBLeu53Ch/Ntic2pwZi6lFq8AGK+Xnr/TXcamySdGfU2x4zbtrEb/uKgoP
aJCPLBPO8LZr6FPQLPIhv2PeeykkhtMVXjCsyj8ObHT9jtimDfynhaZ7gdtudPD//suUZko91I/k
q05akEnFORVz2M7M7wh3qMW/J0Q9MRj2widfLJTa8fwwFGelt29J26jtIfy+Mh+03BFS21Ibl8Ih
EcV0Ko3Mmq/yi0YSQnefpc6K+hNtnEvDzrYnR5RLOx1z/20LQeJBOX8bVpuLW5gBPWmzWmGJizeW
+boxlR8DKHc/lFzpmkZTsfcOGmrSL6zB3vadjJ3i+vqumBOD6tZ0nAjvm4KHP31TeI16mpsnQxVD
704L35qy5Hrn+fDf2CVARJ3q+IyMT02rIE/W6SFj0e2e8a1wDIxqHTh7khh2NP856Tp5QOD27NxK
xT83mHL+4GLMKSQSwPzL1U6YRycxfjXkwmx0JyKmksSQR3PvQryiTPwUeLzNIsFLB8vyKgSro2Xj
a1BAlAL69/MLTpan+EbGnpfnoy0QADIHja0KPF1DUg9qPnpQ+eMH/IMsbkl/D76C2HvZcp9b7OYG
mEUEhY/TkMPwFF1vsfDf3wzvGDvfI3r24bXcoyeLMzsUYnsPMWTUxzI5oM5Z+AOEvN+8dzN3Fwi/
ZLHd1koeqON8VNygu36LFS9MUPCXDqQJCuAFL7ivSnkT/o54SrVLemRhJoFJSCgbubIiiMr3vw0a
vIyliOWFHPyVJFXrnX2KohbBAbu+9gaBANYj25z1+2cJDQHodPGI/DXIQalDN1QdbZ6RKrRcKsib
YuAVU4Z8rbFp1li52gKLsij7UqxQ8vHA5T/3HJFDBRIxDgSRlQnTJb+AqAu9lW0ol0bZfpoETbpc
6qR/W0iKuVjLIRphmhzDMRxsbW90Uoqi20f5VM+9yqOoA+VpH5cYzUYQ4He+EtOXiWA9xhPYZpzi
aIw+tkKMUrBwjmeUIEhRX+sUhBkg7Y/iaj4MngWTN0YYogzC45vePGpf+XR4FyWupemzjjGNbgXs
GTQ5MVmp/PCzIXFyXeiOAv9OI7BF/nrCV0hGZuPTgy2IeVSJfsObPDlukQ1hC4okzEYZU2cvysxm
TsVovWdZSQu4sPybE+uZUPyTIgyRsAX/YorIG3BuufU9Wwc5Q52JCmJj81uf7MR+vN+csvYt5Cxy
fER74ekrDYD78rqkhYy6BiwRLBivgKPmicdmmKAoFaFje7fjrk4Ph9nYD/niVRpFpDsvXTLHxdhr
KW55TGFFIn+tR0ny6QsOmoemTGviddBLM5CR+CW5TJEzkuTBQFfF/uT22P0PQbAyqbxTQfcQWhVq
yg/x1hH//DcrILPGPlEb/H8zNUeGfh4oZUbmBI79qB58rHtDSoC98Kse2GZNU2YK838lKGnU2M2m
Nc4jbIVk4BLfIyHM32U0piI9wOpkg8xKAimkoTOX7iE8GnTjxQs/S7Kxt/pUwpDJkYxczj5liNtX
fKeeYecg/vLlbRAYMOrYCSRGPLRw0G/mKTM7NpR5aTq6+89KjGTo5lcyFWf9ehnTiqGcIrSClOdc
dct20LZX1gNjfj+QQSfcNTAtpZbvmeSDMXJ2GNlYzdVcLU23B/9/QBucj6Y4/8JqP0qK4D6ARipH
eI2Hfiy+NjQmW+wDf+Q3KX1zvdPWDlr4ya4ysbmtFQ9WUCoVYexH7on6jsx0+blz+AfeWZ/5SO+n
hrQlO/7aizDovAVxN51SFbsMuFFueRmr7i2r2wzUvOnYMLigWw3WabeWTIOpP3HlbyZC6t1fKDFN
U2I94GFIIYchkrKye5rhHA0s1pyMetoH7ndWtNtz9Abu1HofbNqplpHnnIw7OnhqS1FEigKjAtXs
DMxlUfW1IxsqvUwaPDAa/okUB9izu9TKX/ggysKOHL1Whlef99Y/B01vPkFf6jz8fH3dTQmzPpaM
IcspJs7PnRtW7KfhM9VW3iKqdaAeFnfr62oD/pqoJ9CLEd6mvMRQzVzQiRnnhc4Qw5IzPfkUm1iC
4N6lMj6/p/H478o57u3NkoE61OzLQCipN2NrPszBhjz9+eP3PSRsEgtlm1iJfOM+GXbf6ZjOJt0Y
za9JWmtQPABGFhHuJbfmKksmULouAWJV153xsseoMeMpFE0WGdqHoE63CWfuYbeRUWbh5Ok50uex
bjYiVEahjZYaREf0TrKD4bugDxVEIaZOUBhQ59J3g2IkLcFfv39H2Wugi+JXPRJ5gaCWIu8s0XTu
td1YOJHYGIHqohSaVqBUpRTJ242P84mvmRNusVinCymtEM4pamph4WDNH22ngl6Yz+XCeOwxggWX
vIA2s0SVtdNuHC4Yc/qPJ+kKGkmoPPoLbpnXw+fXw4KPx+xTHLiGSfixtHr8cfSlLS18qjfrVQPb
a62HqGrdvZfQ9yc2QtykGuV75K9U4mRSqnzNc93wfVrBxcniaMPa6UCQkZlYUdOkm4UAejDvoKIw
2gSDylfhyQusj24C5Ot4Km6DyPJQOYrHi0AKWNIoSXp1B42gOul2e0AqnvE/NAzeWbVGdKlgZ4Z8
4hQ3eBTlArzkkCxchcWju9RgzcKEtVbkeGn+3yYvR0lVEP65zkq0CHY4kCQ762nam2IIsnqmc68t
fXUn9T4EgoLr0jr65H+v1zlV794rOlmpRMlyCjQsNBwTfhl9X7rrTnkk3FaRiCcIVfrXRWOUGiMk
sm/Zk0YrogafItUbl4IpID7K6piOQYwMaA0J7Lj/pDG4J7WeR5ecvxJBU05cCiaD6H4ntPHACOpP
lRtwR6YdGiaWSamL1rlZcEUxcihjfb8qz18MdOrLhGPSIzSUh6Z1A2ZQXLYRc0L9uZOchzKgC7U3
xfMD0SenO7/RQmYHknzeaL6LPkmieMcEiLFh0KHjZ11dbwudZw1sza+05rrDPnfN/CUoWOZ08OBQ
5W8caBblBINq/c3dcU79MpN8FNbe/5jgVrxQNFoLbNV0LyEDP6lHK0ADV5+AqZx2twxZhym1kmg1
ymp0C+DhtPsN1f5j682JX5uYX+yn/8NCMDmlyumtlFkxzdMLjXJf/A7oEa+2mfUS375tlaGElG7w
e/Pwm9qo0qZlEGHuur3AS74U7rs28LHhvfy2i0xfVZZjT6pJFOFkNKGyP78z4x+MFMbrJ7V18z4x
inD4CHxiLxQQYuoJHBTg9ig0Tt6FVvAH/Can03hZdO+eh/j82W9dnJxSmRVrbHgaBPVOjc+slk/N
kSBB+OW4kCMEX1XFfhOTqV0wcNtzwOC2tNKor34nrszkhb96fzOl1Y9UnIHV7P2FfEQZ80CN3FF0
3XEgC9xCMCwDmRou1XePP2I+Ol/7DJB5zZsihu94WmO+imCpxXhu7OuahPpG8H8nd35L9wSnexRU
HhrOeq4Ubb/5+gN2of7OCMP0RZRZt5FAz9dejMLDzCne/QDT8tveJVLnzZxrdNeZTPFuixTvSA/a
T19GXZYxL/HZzoaMXO+9UUPGYuERQrvce7Z4HjozL2VgqGls9go+6h5yGH5jT1EtcYH70A1YmsY/
YujTe77WizHII/7yvX+S/ngEtjvlJNCFoVLLTDYZkxuiw2+RfP/Hq27dtwiyviu53wqVdb8PZbbU
39WI6Losll6jfbtu2j+aIL1Lz+Te2yaL1wvJID1tEWxt8CFa9fHawZjbxTbAstszbBbLYRciiOQE
AX1xxbTX0mGLIBzKwIDSvbygw88levlxfgoepViP66Sl8IQt2ZXw/yPaJA0nVhR8f+zmQwotEs32
24A0BYeCFnk6qiRVEy/8mxR7oWLNdXjHKB+pvaeE91xf0l8VKZ3ZbjE2CLTeZcU2Fxft2YwgzFKQ
YKn49Vch0F4iWqEVMdgYTAT6MY4zVh2rJ37DxA7f4yhctMD1SbXf/zSj8Yc0ezoxf+NZ6FvvSidO
msXdR+OaSCLjex5BlJInQ5PoNqa7z8jqy7CIMxNXRUsRSPzdukicTIOsTq8bNFp7jO/iKcIn56gc
DPHxwgk6M/0VqpXDWI6SRu7kBy30NdX8uiP8xS1Myik/2ZOpY/eIomeKG9UZD5Ijxu2ltwpw0jB+
faFEjVl99LD8Jwr2Mf0693/zimyEDJWq/WpedfjJx9Ww+QWcd09OAcE12OYmQm0OGjE5oZIbNUC8
XUIVizqQLMVDCut6GpLTEZ6YGL4YAbfULM6UrBsaK17lsy2DHs4UXtTQVRxvekBW5a/1ywmTEkgW
7idq4pMIG0weBKVqCoSEy8PQk4HnRyh617HIn5g1V1Pg89TB1E9Pvq0+TssHm8M/zk6eqEIyDW4N
DNBgSWO9blX3aaSk1QQ7SAktYpQSuESoOUtNn6+21tZNqsvx7NADoGiP7srJU1sBTKEAy1O3oR8A
x2wJML/zSnHv/9ze8ExDtEbG9f2/6h7WjciQeoPzzFOoXTY+GpkmHMqfI6Y4P6XDkT3C3caWGxLZ
iQHxSHQYOL/9vHQsPbaA0+xTHTCpuAqqnzbE1jvsERycCOoZS11fF2gJs4Mt+KZnn65Un1cs+zIE
Bm7+iprlFsQmyu6rJS+82kVg++pZnszG4G2SwJ1AUn4hw015XJXicjdUpVHjiVQTkFdxnNZCLutM
8d1tcyAbtoc2TeGcvXMjKzyeLSbOkQLyB6KERXJH219+GxMtNTG8LfKDTi2CfTreqx7DiyfJycMw
0K89V1of+XAm43haUVv6bXIeCI2r3Tyg2oBe/TiX0M2wJE1pq//koqcSKcG1kHxk4PrsgkWO6NDI
x8zLRz9xKSumn3jDJOS1OgEjeiXcYVrm3ZgSXkkpRbEW9S/tbvsW5QffylbDDmfCBkh/ndjbovuh
VqwaXnrLk62RfjveqB6mBABXlnLuhtYl8oBeTps2H0INwcOEAZfg5mibfZOehJUgH/KAjHy2k6bN
wIxKoOZ+gKkIk2yAd6tYnGEdAGdZZcqa/58vzIzVHS4aam0x6R0mSyGFPfB2JLiGGGTbDn2zwIHR
3KJBOb/+U/R3u3XnjoTeKmZSZ0wruI24j9QItjjkhSLdpc0v7bpId7B/+cX8J6T+FRgdmub2UAT1
L5ngN1lLdyNlgscjC6DsNCxTLsIgTpG01pzsEbphp3JB6JKCgpEe+q7+AF7MkMgPa02PSpUc4WXx
2MTE1MA628hNE1LGx1MBXvW4uvtnk+sljQDDH6mDXYI4Wth57KNJrMQ1NfhI6XV8DuoLOQBRkrH+
osSWkBt7CY1KbXjAnMIsFNKL1z85TSXvVrjU1h2g7l212ErXjUcftSEKAM1di8HqkyxGHfwW8519
jC88UyfmDw5Gsxp+GkOtG/DEWh1rfajQfs/y7nZFS5BPNtCDiK639mbJ+U4kUCs2kS6Hq/AhfucI
DAomUommnCgpSkgLq2N4VkAjxaenQwmn+Jm9ys8Rii60+qmSUfUCG2m/WlKJbe4h3HJzvLiAuaxU
yBLYwDiGPPQvNLeAVVUBUOgovoVuWggeiL9v46tIZFRuLf3ah1GP6f/P+isezLXC4wSEMaLJYmlO
TMOXod+TUpFbkb/gMtunqbzmHLq1Zj2hSDktJc4AbVfw5YeMtyhRV6eXt1026mG2zmN5tHYTt92D
FKbuEZfN7rbJFrj5lnJ8pQoMqxVinR+HezG/LljnehVFoNsNYHCAmC+lZoi/7o9lkl+K6bVD+TXh
mzz4VKaS3/ieaPAQApmKnVXELXUfSUYJgOnjkd3NS+XjXT5OZVmkjXzlf4KilWJKlmwi2K6P6Gkv
XgtzvXwGKFPiosb1eQQ6aSTbQnc0AVgAkOYP+tVCMTFkoozKggD36S0eX1Efnh5skn+wJ/ECbfif
Qz20rvdUY59cUMzly9BSgtYc2vXA2RmLsKnLTYOBwI+3+9v1VubdhP4veSbFNjquVDW//1VEgwXJ
hLCC5J4JUq34Qy3m9upQm4RfyH9LgufeqJfeKQ9OWA8mYvs5ZTZU7TEoamp04MEhgtnFxY+hJfQn
xWUz69q677A1+Za/j/P3llehtWYG2Ndv8KxYOcAHYM85ilzXvIlsv+soRcHvA4p56OFW7MffImtQ
ojkH/SWgEeXdVwUtBJSEjDoWwNZwSt+C9APEQSQtrAOfygbh7CdaK1B6kQsgfQyibSmbz+RlEHrM
I1+b3sgpAkhAfhZFetfFuMUHWp4Ly8emvAp4/4y2jlHDpXtnMqNzBQHyaT6TrOxSktBDuFhtYG2r
6S8H/3afSbArtC9eHhC1pfUB2fH3YzNlxjutyU4IMRVNWWIzDqm60DhTknbCVLwl5ZUoweB3OwUO
4rKaE1NZTniid3oK1uUaUkeJbfIIin0tUowdcu8rZ3wgh14rAKztfhI7JnsPa6CjTOofIFOxXJzw
gtPJRJjLFndTZtIYabQR/7gktLlfQPpbQpboUZABmelnX9iCrcbytCoOScb0ZvyziIm9kzsvs30g
XrjMnj6tR94G30oCDMHi283pxGw+Y72Lo3M126EQ0cTMU44uDiwieS50F0c/J9W34wdmadsUig3P
q/ccrBFJ9AFngmbr4jtrjIj5Vx3Jxpww/KXdDV99+A6oJBPOULLl/2DBNns79sYOxXpgOsB/OfS7
SLrswVdUAOKixICEBf/HZDF0im++AP54O9+UJGiDMtkAsYGZU0Ef3tCtwuV9rscJwmCIzSCY3UBS
wxQ0JqQto40zTdhHJdBJzakKGcDk6UC4E9h9bAOmGyMJzFfEt5QRTKhGefw0GS23cY+tlVuQgMYP
jmOTx3WN5nxYG1xam66ymBqwb8lN7ZQZW+hWfb3DpG7/wT1ms2uLEO8UQLk2zs6B0+AEV2MGOrH1
JrCZYPLtS/tVkMwv+PoHK3p1UKergewA2MXCL6rvCKVxY36uFSQf0brOazTeYZ6OYk1SxWOcsoVV
KjORUqgdLfExaqbFh9DPxmctFWNBj7/8u8jT53fzVRDHFJ0Bu0v/bVwbvz8ogLaYoRdiJq3O6XRg
mqtM9XbADjzxQ0eUPnBMGbV5Tq+yAjX4IHfI31e5GFQVIgE1nBh6ahFagsmCgrl51Kbn+wXh4WBw
MU2h2KOtp6iSss5GRB4OLE9xWy1ZtaNkUHHaAzBAzISHskEHEP1JjCkQ2r21wFMOI3ho0lQ28b3X
iw2cLKY50nFQ6PqP89AwP50965z4aX8mTC1+7p2Bmf9fi0B0bGfj7Gdlioy/Br18pYZGUSt1sdzx
jRz3ya8WQxBsVROfSfMC2rrVsfkzj2CWTg2I5ouUpjpEoO/6R7Cm6/1ZtTuA4OuGsKYIHPkhIAkg
YDe73JGBs/ncFpkjHizEujGvr3ySWsaPyFUKQYV1NHUvMbS+XUmgVO3gAkMoxnaEeSI86ci/qsga
Z2UoPprXGAtx/qe9IBKFWA8nVObXhcIgFLQ+ch8TaRbxJXRvrTibjkoTay277Q9vH3GqhzRoaPgY
4YHlk/ft3BJ2d/Uq96rGXO/cp12Q7tlOXRm9PWkTKU73Utldp3ANjeHNS58shlEhCHA9/G8BIYlS
e7rX86orIfOJPLn4cgSnpAOJfeTGhmpBfAB73cdZ3/DZR9GzQ21JmO87AFzDtSI2sM5kTnV3GXat
GqRDa5/TBmhYuykf4n/xX0g5JIX9vGn0BK37xrg8lapgD+5g0ovxU1Sth1+oQs6OivI2Mdndaju9
uVq99Ys1p5OvxuzHeDJUwAq3R7rL0WBqssVJ/HGfnVEUa5TkkHkXo9uxnilu7CtZfmsPWeNVvjx5
P7KHh3KHPFBU88HH00eyM+Ybw/195Z+sRqSh9gN78i3/8oNh8E0GuNYWno3H7FWLA+QlvtUNe/lR
/uOUgdF8yLEPXf+pYednZI4CrbAeNMi1hYjTugdVuz7skWJsNGirmdvVp4kjirHr3alnrQe9T5lF
hUh6S8IRUUvRVOrP7NtQiGxo+zt1xfHvqNsnz+9NYkAw5TshQLAK9zhdhInGlLmnlSoUMf/xKkDU
B0rPDDqbbgor0T/kcEosrn1azWqRLhenpXCfSRMIGkIR1Ie12mLkbodCb7XArJ21274+GAH5NyCk
NPevvoBovvO7J/8y9BZq49l0U0eNYGhHqbSqF4i8VSjzOY4y13z3kLdVObDFCgpbPLs8GJ6b1v6r
6ZBnM5y0MA2E2EG5W5hPeZwg5WkW7/3QMgzbCC4OJGYMdJ4lHsSoVzc66Rrw0DgPhqjqXqf61dg1
XHfuJC4eS9CXfeBnG+F0g8++BjHRHXFyvcXnwfF3J3b/gX4RD+2pKd2ybURmY8B0ZxxXoENLRmMU
C4ABRQ7PL3J00SmHtBTX9Fuua8mDKqlxDST2rU9GexomVwjGL4pqPJUopeni9EoJoMOSaRSeUzCi
KX69KHNFyX2851JUn2eX/OqlwhlucHQFRi0KqgfvJkFLLano9rT151GP35dxzxKZwhP4QldCB351
/Gz+nBTSmr/ZRxUjuCFsW7C9EQ/9KFPULjB8VK1DTQZsf+81DqQrQ8TE6SZM72ZlJI6Dhdd6hdrl
4wXHWwvQRVxUpqEmiEh0/lACVpdrQ5dwAWnhO7kuZXRMr3xVDfEpwfHbWtRz9fIM9/XEVpaBy82M
g5GuUs66EjgwBaVwCPcjMGE/JJVqOpGwi65T2FMg3R56lfS2vZoPu1PeTECg8q5wqK+MrM/CXVV0
owmjqC2qUKQyUJbVe6urIAu9lGuZV7EPtFhxWW9RVFvhuV/7eagE5to0H4me2uAOgPJSeRiiuOE8
UQ82LldOAMdg2jv6Va0pwuryH8nvZU00NVugACY7F0n4EGwNXeEpIub98SWDTVD/nreqerUsS4+t
0Sds0LIIUx6gY/zt77Ot8/6/+7yoO0KLdKkpdPej6SrA9KHyEOU3inQM2/TjiUOkhG5Fxi1OBEt/
BPgmCouHetSjpt5kscGjvjoCe/BtwFhGG7ah1rQ13bk4mVde7+cqxXatfHNPP/CaqnNvkLWfPwCc
2Oy+Zn4CrJ//CxbulqEPUAfSySwevOyZ4KLmLSvefvBn17rtQvu0WgCfvzljjMBWg8Z4mNDbgBqX
S2rM+dK1+M18+Z24epB/gm4wWwtyHGndIbKxrHJz3ckM0QhF2OSI+oWhwN9QDqeiUYR9rlBT8sIA
CNbhNl+Cne50sXhg468jBpWCLK6P+Heittm6VRaJg5mUvv89ifupiiuhgizqIahvtEPlK/8nV9SL
A/+oz2kTWy6ZkKpH/jpc3+V3QnzWMxXILTGxxyhVtACPoOdz/fTDJlVjeJz6aPwSyaioy9EQS0ls
95C5BAVnJLevS6inCiOD7lwh4gbYL3yXMLykoSXY36WjU84sqwWyU+hr3uyFUXseXs3jVMME6j4K
ppP9kju3zBZOmGDS1otwaXIPewOns58R2ZhEmVGzjxyN15qQIWURs3Z/gs/4odGaV+ybe0I1E4Vj
BmPYEUZmDILRU/InAjlp3/5UNbbzjjex/C9V5+dJ5XQ/+6c4BjE0iNKYH1A+T7I8TiEf0y2vTUgR
bvpTkrj8rq9sfyJqg/ZKvSR4UqNrGBz1PRosZYtpVzCJZXmgDwcsqEZfeRGCJkgyghaqJIdRiMBt
WSQaX8eG9cFHIVfokOjfv3dfWQqXpazOEKwwUwO5w8U8dBpWwkPMNRLSv7pYXD7KheYIaR0QAxFM
3lQYp5NmTimMkc8hqwTxuqhFiDJ9pFP3eX5b8HpPPdjs9LPuftCbhnWCnjv3dz42YKvQb8PRoBxk
94jh9XHF3JqML4X/Ato7POtuhIV9RjeBwgAXWzjlbUOn6GGAwAplykIFAH2Nuoh95Hw5p2VObIgK
/FXd2FQ5IAAahEsAODeFjnJc41Xuc4w3exqkPjtR8K5P9AqBJjQ3d34nMBcTbIQzQozrORq/RCkN
RleEn4SvgDA8RkOaBJBifYbV0sXGmM9Kxhg8lfKVFpzaPucHLpJdlSTksedC9jSLfFEDEJ/IloCN
itapX6Dm9HEqzoOuFp1rcPSupRPh2IIOxHdR4KjtdvnpdPaDrw9O1s4s4uhVVfiirw2stHuTIcPw
NQmeSKI9dec/AK8oozyqqs2zJfKAzvBIq4RUzL92KUZy8HO4wt4iwCelfkH4VsVNfXBlTrEefxXb
ru5lPqicKd8+Fo8Lr/QSY2eupbsDq+5bBL0jC0RD4WgWKyy79W7RWCqfyrIalsnLD/ys6gttGlQ7
o/A3jFjVgMpoI5BqhZvmyiShzqZRx/04KheR9ZzxkXijqU2tMVItOoA9ItPoy3GCH6R8kT9aAl5c
hSUAM4ypdZShJqswLTZO2zK2qp4jUsz3OtpOf3gHHy142xg5/BIt9ozmB3noL0LpYmsjS/MDjmxD
7pwsayeIIASQz//0fq783sUh4XudjE2Jq06+VTmstvLmHnkSjP8mChyMCN/svcjXu7pd1VVgd8RQ
2Ct2iO0MsMSeJNBv+0KSSVirjEPpXGqbX1v+LlZbSwKXdB1qtiD+6zj0V1mLSPLw/FkjoAA5Frvs
S78GXzYtPQ+Qb2Xp/he9yiKK/HvFWnk/btJ9kq3Kx4krqr4PRPpnSsJYKUy2BthUL/f40k2Gu7DY
3UxxLFPmKZ5dUa8l4tgnmj+w1Ma2wNINOq2522Bcfibbe4ycBdJ5DFPiS1912gmlg6T5ihQly+uZ
A65s3FW+CIyki0sc1+f+UwTM1xdbx8oIJeaVqgjJV/CTjh6M+iM+h6pa9hFFBsJEk9sEaVt22ndo
Pyn5IBibA3qrcAYStMSy1asVn+gcYOe/UuHwNz00FZ5v65Qpr3qiHZyDIX/nql63A/futqyJOO7o
tWaeDESTdsDXBXxTGLUhRw5vm+ASE6LL+pJJCLO+HBl2wi9KXNerCvhtnFI7whkesk6GUMyfZUqk
BL1N/qpqgta2B6QLY7A1I+3/6qu1LCdZPn5cGyRF1TW9FKCJGhF+adQ4zoyW8MgKSPiZzD9h3jkM
j5Lzb+AfDtKibF83B2/jzVvVhlAWWYCu/gzLWT3JFMB9MtFUFRPTIjHm0LbwfFqb43SS9/pjGs5v
d5NQGb0KbtsmP0sV7yAEYWguL0x9X3P3Kf3tG5rqx/Q13uvg3tux6ENUAwHqopdRe80DYFJwq0vX
76YLo4IHZR2ZQtE74b2KZz5KaBrBG2TJMhm/KaFOAPPgie1JKwNDr4o7S2yNDtd/ptwojVNKHerj
iYrlhL5SkJZxc4PJkhJyRro4iGsOgpLWymapwzd4mdYs994qYYvymeAF2Q1r4yVA7DBoDO3jWbi6
8mB+7+Jstm5WaH5ovoi9ny/oMtZUQPVqY3Suq5gnDyiqfkpFD6enQRQKAxtNxcHJluU2hly0n6vI
fK1MxwadM433e+EkkbMnfWLwpI5Zdwn5waKvVvfY70MHwtZkuEkIQ90IYxbFwJor2BRCYxUnrFLG
adFHmrwVtM9jigwhjqmKlG4I1zN3ez04Gv7Xic0AGL8Y5zQ/OBemKkMIw1t6KJo/bkkaxMBvTGO/
atIM2r0YBD0EtgZku/ZOnAMKfo2iOuaRQia3LcICeVDDZms/3NiR3MI5nBQaF0hedoRJsoxbkx3X
VpimG+umBiOVw7voCS6rQI/zOdj5pVGFK2QLntxlqY0aN+VSu85MJPp5c7J5H9Kkp1YHVeokoyHu
GSzVK0Gh+L1349YDLPqNHx7iHXJVouDFc5rW+xagMzCAQCzPANZXh78pGEn1/quNiHfY+vi9lJhe
P/698nIl8DJt0x7xtVqd/rVmJEh0xI6d10MGZjXVk9RqRoqT7mKuYcN7wwtujG37I+g80ej+v+6x
nWAPke3U/lKlE7/poG4vJzmiOkN75QvuE2muUw2vYqkT0zh3LyYKWbbVLpFGlZdYvFuZL25xC0DI
mlKFdb5QuZy3rN2ijNd3F75vEqYvHygdz3TLiGr2tn+rOumtLBwonKNXPHGUh2tq2btSrL6HtcMm
lpabZOQ07d/rN/IzjwHzrK/5Mif26gkU6wEENMo5QqHxAQQKZeKah6DOZR2ICktGXkwTwjkhzqZm
zFXWsVOZlY+tlT21j87tlDeK0K6F9YVnCWcWd66ldIt02VDJklrkg4xMhBkiM5SpZ+yE8AV/Shg3
7nmUW7vylJGupyqNwGiYkmU7XlaMGasMOQ5v4L0BzHXeyaohdTsj42becZybo1j1AEK1QY7AaU7W
SOc37WhHRVlF+cz8KlJ1h7G0i8iRn4ndpaqUfvl6L+pQquh6dP5fChrkI2ZFBQKsuW43abJ2xd7b
K2b5m5C3BzthENTA5K/RbHqAPwOLb44rzLVEyRfLP0IZ+Abo4/5GhX8guolvdo7r0wqnSFjxlN0B
25IfDmp05Hc0Lyib2wTzEoPcKRSsLcE8T/RIcX/xwRlQvVH1XyrLfLIOBoYpCbRojZ3YnE3qxYX+
4xcL6nraKcHfSFn33fzZ9L857g/vS2fYZg2yJKjVa3Ccqz2HcaAhBrHTlPfTpS9MZrwEm+rQYDZi
hAderJuaTYlxxpCEE5k1L8NoJRVXG/24PfY6gMGyOPUlHJfGSX+X2ONnxqGQLdsaoad3tIeDRIzI
m4lZ68VNXUNYrtsQw2et4yrRcEOPdX8eoWZ7LvZHz1QcBwEIW/wNZ5yV/78MAb79miRpggAagAsz
Wwq2CayjgHtKEY/OfSvGZKpD/a9Kcv3hDKNu2bO72ZoHt3WoSHt3lYHRGNG/fKlNtajiERI2bJ+s
jBhia6lbEZiytoxxwF2KjWfjbqrpsLJKqZBXaxsIXq+pTJ/BXqvMz5swyl4XCP7dWvJ8AQbHkykz
0VajQAL/vgVSyTMjEimCAP/q15nPZqWhEZt30whdaikZZM5+6G/xl+ns3p54iB1VJ+wzMtuGjAO1
A/kJHNNbWqdYh3tEakD+tO6954yOCDegPgDFBN+Fxz4cA7r+xL25Zt1AHhXmj9UMIjz2CZZvfFgQ
1PzwOSkaCqCS1MbEhQoKBRhomrEcz7f9N9zPMCCRJlK1STBwlNJlOsrA5xFrBYWoYV/gb4+prNOF
+uh7EH4Nu0INl/F4782S8nlbmudJ/tBSbR3Zf7xhMla/LWrRI4Az4FQcD4Q+a2CVbDYVeJglcvT4
g6NpMkMuM/1pFY1fbwWRK+BBoIfitKV11qnZ5XPrTe6TooBEwW+CZxTo2jgh4tVLdX1m0iklIt43
vQcuEg1HxYq/Faqxywl6PAW5hB92nLHF3+mu7k3MDBz+zUMbqxI1ls54/eNG5zjCO+IubEKMFZP7
bBHfVYb6FEMxOQs8SPALCARJguS9MCdqar+57S2uYNyrHqFfsckuHTu6APGc7YdQNaTO/IK/NshE
62oq5wKbE1EwBcsHBAyhDHKTWFSBqqeqPCfRgIayCuV1rmqQ1sRnKQ3/YvGblU2/u1niZU/BSwdZ
FLlX69fMjRVPtvH0gwQ1uajCbL4XTK1DwlyYbu5OwF6eAu13FgtyQy9oiGH0kIAJKnCWRTWZlleE
Jv/Fmu5wU5Mcq1N+0qKHhXOlclH6zeRx2DJaKg19Hh4zawNNGogthL5Y7Zm2LdzeZBDT8gs3WM6F
IJoIXF9DwO1gGFwedtgWOxwdlTkKCWoFHpnWjO9v+dV9zkgMPgQymyLqUKB/E1/bp8K+t8+XTOAZ
a+nVYTVyoTCUJqN1suMWjU/0KVeTgZz8/3K6Y4fJMHacWvyCkYNqWS10fUzxO4cresnm8guAhd5a
0ZROJq4AAJeky/mMeSZ2D7slbXLb58wQ/IyOIK9ULfmYt7GxIGhZjQk7US6cJGGl8xY1s4KwI9x3
/Xzdj16pyHOfO1xU2g+Hk3zGw+gu/1RHtjp+8At9CU/SfG6MGUNXW8XjxPdyFo58l8Nwk/crItIZ
vPjGpXaAa6waPFW8W1FvTrHBysAlcZwR/wwmh8aNyhxco7NaVgdjyhMgieh/shtovBTFm0aVNot9
3Be6w+QR9Yxe8cvJT8fKlUBXWwZW1C7XugGO0ByGrFpZANXoTbVi8GYiALn29k7Br/aLPzXJxEVf
ZlUINy4JGQR+8wh1Hy7La+lUawM6XYlaBqinQnauD8IXQG8DPY8rRmOtrTbIbgPZSFRidrZuqI2P
vT+pM06DKUuTfiaFUrFXHYWT4j5ZiSfn4xAArKxCa2HjC+enwMcLSLNi4gDemcli7s+GMoFYiKwo
WHrsdXzVlw7ozQ9qhSjdz1QlCuJIajO+BPpnjEKANaGlUTi3FpTGeeyYgO98uNubgiSTluIYzEf0
7nJvIJzPU039cQAXTMTT1QF0jAq82dKQKtgjAxjsF8OdjrId5h9Px5asfvUSbGu2BFo8Xdused9m
ilHPSsSVtpNoLUxS8Ja/nRz6BR/n6D5QoK5wHJUTitDxWRjUmkYC0HhYOjXZYCOw9Y8lL/HkpEZK
BUrLk25FWEgmDVZYDRDAKXk4qa1VX96EZgxs/Edr6TfpRMGgmqYsgEP30xRUUJ/nCAOzoDPkgz2B
Piajnre+3csU5VUmGYQGnDvS9/Gcib9PxsswKCeFyswJ25492YG6/OVKO+vQsVEjcHdYxqxau2CA
jLShNh6odch9uWeOxrvB7C6IlUytCM/LQG0eC4Ctj4u6+YKtGnUvcpSh1D0oO2T41MAIv2JizkRC
shivNSJv6OoxO7mlBpyg+V5IP4wbrSjjmA8kyEuFGcsUIpHR1e3dlBD3TBcqz3iaDGKBz+AkE7uj
cryV4vQbByl8wNYZkC/LWGpPZ/JX2RQ1haaDqHrns7CYYcjlBnTXY67R5oyPpM9S43qIZDqiXYVo
pUcCSPrPSZoM8Y43T0mydxFollyG8Ud6sPreNg2IqbyL3i7N3M6Ro4n0Lmku76YjGPCAWZK1pttb
hUmPz4ukTOCtCEEJA4Y2qT2Bpvxqzqm1Qawqt6wCp2CdgXqCU02VAFUM9rq958HhkmxcDeLSMp4n
9mGdN/Q1T7S2NvK4t8jdstfXLFXNOjJKQUFlghdsZXe5XZrDK5iew9AIZjto+mlQfj82woEaIRgi
9zF33rUELDlMlCOlnS2xPReaE5/6lYhyQoDv8PNUynyknY1Wlmxf0/zjtaB09xJSxb1Wax/Rivah
eO+lKe9D/4u99dazWMbPxYTxgoVnSzegNIxcVBkfCJ2bwCk1kSs5fJqKQc+XZ/0eyXgKP5zQt8Ho
9XXfVHlHOzBvStPh5n4vgLtDV0EfMbrjGjLm51SinyKcuNfnIaUeXJ3ImTlXO7OPlKkVVHYa2llx
DO/VRbOu9EO7eEt2rwy3BnlNye2RI75SYu9BfAvRWqfPjMkTpfNyaseRHHVhMGCS21jiFPj+VC4U
WRRrd9zbYi8SJ5sJR+eZmP8+F6Bcny/CajD+oiR8cqbYpXOVjO/aF9xAhp2zBWbpB6fTejOEOfz+
gY4cJ/Tk2He6kQcboxDjvXI0niShq5FJj8ghuhIs0fKVtSwujGpCPxpkg+VAZLP/4IGn+XBHg3yV
HyV0LP6+nIP2/fjRELS/VjJtP9IAubbp65A9gM3R+sK0MUFHgY/0DL0UrX9GU4Ya9gWK3MvgeSSw
0DG0DNa/ESth4J5ROu4W0+SJ5vITym2UQU2Q6xpDUGxOdf+9kr9G1RRNXkaH9ukIL8MTgdKthUO0
6XImgRt3dJNKF2Qc1/l7MLIJgssSxD1ASYrWwgSwwXv2kXvZeBFinOpGQvoP0Y0MjBKUgyhf25l6
fGkPFsaTqbDl90gKA5UrV/TOBVnDeu4jDtkN0EYCtipx5wSGw4ACpimQU++UY43JKeAwfHxo4eZo
6LPsGnqPTJCz7AQy9GbOA5JaH4jFw3WuRQUKUaumEpDizjWplPdLW2wScJGxccwzPT4v8cXJYVqe
km3kQL051FCPmAgCW2oeK0skj19cVFM843Y2E7W83SZe/aurQl3Tu/ef++6//B1yA7gSperOFmWG
yHHpdbK0ZX51WA+1IhXRQVnP5hYUK5nNjNZ6VQ1shn1JD48j4riQaLpcXPleQnAb9mXmXZYXYMI/
xF/+7CAismDIavmWMNCxln0Gz9bVs/ZbQqH9f67HqE0PmISbX6nyNttJgTN9yS3GxbKfO7Sq8FFY
TplTTlDSYuaHJUqN0VkF47QJzdxFdi6gboo//6z5WyEZb9KYJdL90WxDRogmp90N9Jw+u/XHhqxs
aNeVEiM93ZODm+hM9PhI/oJlYCEZGlFw+8mVt5fKh77GrHy8YRaIGgjIbzUCzWGbPDtQLMBOlTLo
+Tl9UhbZnmPsHJ2+ODdOfiQ46nOwa+ljVFWLy61nHQzsCdNE6q2UqD/sAS4Ch3Endikt4azzSH8O
pH4La+ClHv99oPRMi4shx9tlG4NHJYhvj8OXE2W9wmuYFlIMZaLJAx/8nm7Mvv297gXfyj2eg18O
RRj/uJl+c+OcNj3ZmT+yK1mGoixqdgF/X/QYLmB3OcP1RGFJsFxl/v2+7wg/ZByPy67zPbS0NbpE
bkEH19NCnMRDqFnl2AzMo3WdgAkVfWXV/xFOxJgBcVples5sUxunM5z6Xbn7fHZPmmXn+LYGC7Gm
NArvLvaEi7AxPGxvznJAp7EFSenH8Xk6v4FDNUs6HI1q4LF23Kcc0O6otScZ3t6YNGB4zqDOmKyc
SwAN/3joWEmw8pjxocOzXvRMf72aaGpKNboVNN7j/hkLFLiyih+VFhjL387P1dW0ksaFdKKwTZ1F
u6FZMLtRLJHuBSNJW/DVGpwoQ5GQALf5yU5UOr8215Ki1ARaBcPS9M3ylGxsIkmM2vlcn28IGOyI
baIysrTCZQcqMAEJWwLC2Vo+u9yxjwturoeqkZCIdN6JjopfK+1bYUJNLB4n/Vf0eWgR8NGHVrrT
E1pyrEZtWZUFxnjUQmOe3PMU2A2l7la9nwF7lBfLlesGMbP8B3q7SAIzecn/osA5OBhii4X6BUdF
P6Q90YElutc2feds5U8EaLPaPU95prORi7JeIPrBFYR5h8nUfmTpyvvMzKU9G3x2F6t+mJ6PUDjs
Jz5O8+ox5OuQ7aTUW6CIQkZDdqUNg0jTtzBSh3yj8RJYhxPKi8J3BI1HHOTvAEyj4tQxsHM3yvfT
dmxKedh8KvGK8wuWlPCwVDI/Qg7qbp4HrQ9CVIpnzWFddttrTyO2R3UrlVEAq6yQL1vOj0A5Jyyx
2hAdkbf8+tMGyWzFKforWDW9UjfDCAENA2eDc0Ql2ClBFsLH8+IqhtBEdmjZ4T9k5awh809MBwB/
/aJcri5SNNh1x570bfuvYISTWqZMrCru5zDUaB3cbfPB+L1maFsO1JSiPoiI86r83GUY+Oa68D2P
sKRwBGzo+TJL5QNEE6lisKtXg2AoWXva1lKoUqrLR7IpJvgyMCNYUmEIOp5mBgtvSuurGqGFc6ky
AKnGNTT1DklCJ/ODrVVThpYwxXzQSjwyo2wA4FW58ZRULPqZG5hr9jtjo1r7ZFlexsHxsAx3D+nv
2w6k3tnYofRHGFdF2B47PM3E0ZRIltt7rPQf8UMFcF5fWD5QwZLCCiL7FmI4HK+vY4MMbOpexFPu
1yNJDDzo8o5MvwYZ4JYq3b6O3JgZM2GhLG2GtFFKwurgW0jFvxF1AGNxsljpB5G/9wFtGxH5LLwr
oVwvWVf1Rp+yan8CH57wb3+T7inyf7N1YAgUnCQ3fzHPk2f4DLijGNL52tiWMOxqQjEHbCGejKBv
+h6ZMMp30jzcIK2q5kaEJo9AkKqP4J2NinBBehnswKj1sUvsGJrVG+R+FijxoH4PkVXXTRrvGGzU
NONHmauHoeo66RvuZMzVomE/EJnYSg7CVldrGibHCAeB+Fuc+QRnvvLlTBD5kGcmbDUK9ye1PsCQ
4ZwbAZQG8NQblDjwD15aZAt5GX+yKRaPsH3d10GQVI9DtN118aT2nxiWfcAagOaRTZXdBZ0AezrA
dKz99TfOgwLcBMp8yMQR7/6p96UWMXyRnNHgSrtWXfXsPuEt5AtyCP88Wyt+YA9qwu9mfRLQHhnh
JDkYqmu7Bz2sANooKipS/PxBmcJgADP1NN6HaF3TIjDNcP8wc0Xf0dR71f+Od/G12EtNZUukH7Ve
/o13xSYAUu32WmamUmgq7AoJFN27xq7sFvyPy9leSoBL9pMIlq0DsYv7V+uox5Wk8gokmUAoaroh
xgIkOjTQ1D3dTGVrO1uSAms8J9IXE4hLhSMt2vRHjBnYLL+yTMfR0aLxHuxn/6k57wgFDj+bbYHp
BBFfOr2Nay/ISuL/duuyn54GWzB31RJTU2fBAXdmN6EmJmA5jXkr3Mh4ruw0/az25C9PMeI8GJtK
loZpf28WYDMb8XjQORW95uP5A2T59F86pSMi9Whb6hEWeFC6gIGQNCu0A1zZlp8gn2FE4are1NJe
eQJsPjfWN1JOMy3n8NEvwSHQm3SXilKKx/iaxJljZCVw17W0HidcOdNQ/PFEvg9yRLKGmnQel0pi
UUhdp2hUbOnF4adqy3L6vkH5x2r6IQ8V3LPUdIBC7aokt0Mf7+0YWuc4dAlG5yGWFhLpI8xjYNb4
5xlNy435lgZDVpQJvcba50/Y+PaRMGQSIaVQMpKGjxr3gapTK80SQtmxDsEmvNyeosqPXLE4XEz/
ZgDOyntb0rvXndO63XUi4xgyDA7unUPRYipozZz+2SY0TwcUqNt7eYOkZiN4zr9WT3nRVdtXWu3K
Ac+fMzU6/WlaIf3T/Vu3r6n/lk6TqVmye7kpC+j9YZXHHggBL/Dwwev8tohXlt4n0n2gIRWnBWaC
3+TlDjT2nTkpe4LP6x/s7tuS32Oa2okVFKv7mSPs2FE/z3YkrbsEwOwpA/bnvs6yh31/S8Z6LEC1
hENL7d96sWZk0z8LVO7FxiuoEBpQzBsN2ZzVinoTr4Qm92ihi8q0A2XZyKsD5/04RYMThSnOL0nX
WYbkrZVHUWe/x4r98Yorbv9Je9DJIYLvCd5rSdvHvOyZt3DoDipF/6q2PPhdqaJFpouN4FPd5c3Z
JmsnrpHZGEc4JMj+JZ7rMnY6ZDGD5En6O9xXJtZOroQUJzvEFh6o9yA1HD7Lqm4qPWGRwO38gfRw
Fu2WTecRHZtAJpyOx6hUcycuSYIeeMVF4wYm5alpXPKMja05QfRDk1aBzxd9e6tk60tMU6szFERy
6eZQZg24nQQ1KoRGPQv2imfHrMBAaU4+CEO8qA0t5/qjGf41nLaYuGvfC5geOI04+U/k6msGaKT9
SfZ5zr1DnEuo+4XFn2En7RqgT3GCgkHmplwPdk3pn8U/nxradNAedq3edeBDx+P3uGRMmrApeFIj
/xQyUgB8Vwoe4SdStOpBjo6FUL7OY/1EfQ3NJFPl9MgvWTgnGc7pGIdWNuHUEomjJ1VkvVlGKcRR
uxtObssV9YGoS8qNDX7mXe1/6mL3pZgRcrIp5aDeLWUVL+/cQqKP2AuFpt8oD1QuNaXJ5FcAPmEh
DQ9JL2m/khc3d17HI9MxnLLqubRigbwItW+LKI3nLLXvUkhQVlc3kMhzdXxjBNtMH2iT5NhKLlbd
J/ctFP6k+jiMhRqNCj4kZd5etgGigWpHA9I8Ic4sd/PPMWitHCNSOwgqQtDtk8uYGBAho6NvfzLQ
U2nD9ZUd+Tu6lU58M4NNDzuKUC3/rK2k/akc2DwzPUmH1qzDtlatDWzvM+9mtlxOhyCw0e9BBZwO
p01qjR02+DFdpHt2Cs6IN1PEkVzFONpcw1eQrw27gv5paLh5PuHM1sYynouSMMwDcO6RtIYk+uND
ukh/aaghZvxu9Qa58qNKytckkkv0yP6Ij1Ig43OBGXh+gzACugkhVnGC4n3maCf6Vhy27TCZ4WRC
54qNzDUF3VEWX0yvdVTFbS1M1bJes39qA3Fw5m+kUED01xAherVHfIFQx0DvmL14HjQft/KjFrWc
/YLjgxjDlFx5smcoaiOG6mmzai0hXwj3qG9yi2UaYTM4/ZqcQFdbPnvwj1Jcm6bQ/UyLnikDbgPA
tXkc4HU6IPRGdTabwRiTW3FWDhC4U+b2tRRV9EYYtRyriHnnaKDYRfm1m7gbIHdGN4Dd/nAdWssX
mvK7A6tU3sssSff6dVUtquDdgAWgUKHO1JoWx+DJf/2TXQzARmcaqwJf/eqYl1FeCU5p7iBHSL+O
IAcrBYzeO2DhvYHRyg7sO0rr0MX0O7lrMdV1Shy3Mkm1TJVMooR1stu73a6rsjZ/DJDV1+N8uPce
Z/Vq4D5qCaIQYSrKkWJ64ggpa+PnsnatnuMDSV6RdJWi8dYyyijOyy/EkoRaNXTYgyHNLDl8iWy/
btnsk8LaJO3bgtB+bfZEr57/cDy4yATE4chdamXhoMuvMR0sCyLR7ujrHmXcI7hwbCf9dj955JiG
46xzyqF+qeo6wUWwPvMB3kmbmwaxWiNeZUhWCZ5oz/xjvtDV5zLBXua/Tt60U0wjLEYqRc4KV4qR
OmJ0PXhGNL2zdHH5nIqNgtJM43dQFaL7tlOPR25FS1D4hfVQjW2ZMXC/e/l9COouCXDek5UGxDRX
wIxx6nucTmYFwJZxvOX4kCyYyEFf/bHlpW7UWJXzA5oB+NOFT3j3/IEAUtMGfah0D4iZ/ZGS27fc
GWAVhkeXX+5AGfYmGxCLMuYCaDcO4RIqeLgGYf4mpQ9uMR0GjaOoKovynisOCGcNqNjKj1YO0q4O
H1uMtQzLT01ZSPIKRuQAMvAd9Cp0BOuAuPdIIi2Q+R3gVZUN1vAPUhcxHvokqmY/GhHYGkBYwXg5
OmUMbkpny9cxdgOdyIf8Se0VOTTuWd7/KjIRlFxr5i8C/meOTV3ZAPasUJDeAYxS00rVfRgkK0Sb
STXSo5GAum1Iz2c7QEAgYNDGAOqpRx9BZiSSea2Wou0r7ljrqz2jpolC1EG9hOQ1l9GDrjXne88d
4ZpgQqGK/M2Cd3/UqI9TZ2iGqWbtGSNmu77HH8QVVGYdc8FcDslOiAtle9x9T0FKZ8nyEK2VoOQN
ZBD7iOYtOBqUR7YXhDLyOculEvgQqJnY4ARWJD9GIwYevWJsprT/rb1RcxsU+Q+eMQ32Ot+tD2dz
nYD3gUdwcGt1t3vnTRWlqGd3xh1bW1W5fAL4gLyOXyX07Zjr1cscFSn85ONH+x+nV85z0tj0xk+I
sXvYhr7ZjbIsPVrfJ37znqYXymRsuslUAZZqBI48B22f7yAvlLaokwd3RdVrg7lu1vCoMInNBKSv
Kffwx70dk3oDO8Rzdlv0JQllqbz74qhgJzbHF/HuS1t5MUGBjcqXWKKijyuxNPBXRoG7hKvicSZz
5QhgHd5NlQFX432TwvgXLzdbHZdyEMbtQcZZ4132BDT407WF6YNk3I7gBwuNmKl7IllXh/movGss
mdQvjtuNkxteFoDKOgWxp77kmt72Rtcdv3ZnogMkykwwzdppQEVtw6Dp3uNZQIdDDMLY1gxOOYX7
YTlXdkZRyuptJlCs6+CELYav0X6JPzDRfjMolb25Cg8nPXfSBmWiFGLnNbV8Uyz5jy0w0UkM9XkY
fwBwfLiDMM85FiEDzVlIrqBeXKO852Q8+O0jS7T5a6nEX26hPTwRWPPv8NWHz7vA+Xvvdlvfsatc
EWt+mq9cycBZYnW//2CJxKx8YwsgetpSe6NrMe6eDnE9jMObgHtLp/G62SxAjHjIFLxfwxoQyjIt
nKKA/UonoM0AwZhW/HbFR/qk1zpg0S481AqYS2oqtju1rw1ceGM12QHIsQm6yNChw+LnwM8K54Bc
MJG7xPsHzzg5ku4xVtEoBcyyERo6c2Rj6OSsCH3SKXB3q0nfRGKvWCGsTubVjIlCG3ap63+Gy1SU
5addEhtG6kTR1HkKNFJ7TX1Nhi31sX+dl6mFl49dAkRN/2H4JkyzXwFbL8UyQWXewfkXM0vC7dJ9
czEMCrhGKZOTUVO0LIAERCKazfVzyyUO0zqkFEr3h9B3gosIuAgVT1yYnvfot5UZrGICKbzsPtfG
Cm+uajPLKqiyuhBY60JV2K9bgk14JpADsT3KbF50yUTQ0TZ2Xb+Lovy3r+sobJ11idPfCbHzvrW5
3aj1DPWWvgNfcZ5a2eE0hj354BAVlnNjVJXRWIBlsnr6fBad5kRZ2mC382lFvAtoHTHNZubABJkg
uf6ZaNHejeOJBmudpBuvax6a/rd0g2mnVhdTaFQ0C/IzTx1H9O7fM6s/DMJ/eVq1/EY2OrRc9NZX
Gpu37wdYV098pHDeu6KPzcRGFl0BYWqAPN/rum9SFTDbsEAEPrfq4mfMvhCAj2xJYLXkZvlcgGff
sVw3QlBnXUMva3M06hrkUm/DGB/VwBuGvQ8o9NPbSVt4kDojWVoH7owuBkGBKa5dZCbYffUd5NK3
aadIcL+1v2IkGXFE5nv0cI2gnXF832lLqvEE2cQEeLvqPmwrhlPzEQKZFkIX14ajFqQQlQ/d7xyL
b80Y6GTV5TRqt3h3ytjOtw6Q8Er5nfqAMp3SavR/kTjDbSASNSuDc4sKbf/EKk4jnO2tYEkq8DST
RCKe/DcHslywb+23WZZCmRyMqHoVZtGKBOyi/VhAn6rkF7urhbRiK2UTFNFbSgsbObUTT4OpkGfm
4ZDKAMvcgI37lbwugE5AXxO56bDDppT51O81kP/IvoiDRgf9q4lpsaP07Nr0HPYmQ6srjcD0mPgK
EvJMarJ/5Uk4y31F/EdkVBMlAt16bbl1wKttTKsKLupYpNPTA+UQKvRF3bRvEBa/F6TKeOb3ObuL
RgszocvO2bgU+IxZHGfM7u2d0nxouZBqUckwEs0pUMinJecOtbGVnwcB+2RRD7VOR+eUTF7bcrl9
dFyMSWgipfzsiGiPvPYht2GfUfWBsq2yYXR2ZNWN0La6L5WqqtYV2egUWLYDxf5MHw00qzWncb+M
CbOrKRvZiSkli3VNO8NM7fJF4HQc9nxQ/n1Ok4ov8krs+RAdFffWFMgW4Z5/TcGuwQgRLvxiodAU
o4Z7qQ4wmsAXLbkSG2oVTsa3x78Xru26zzgMhGS+biJhBOBHrf0P4ybRUA3ZV9tYLMd4XS3XyPVv
NcXAjAIqtwNyB7Id//x/DaoFwsUCTer9o0GqTDqjFpMsNPHQXD9STkYNmbATLgwAghr/awMeJMRb
gU10vrKghW4RWKlmysXSkk+QoDCkty19jKKEWcU8PfGkKsOYI6hS4JAvHzW2GbGPa1gGeM7txiEv
AQd5aMogS5Y4wzDrH6TTNTQP32cTr6EIOzZQB9oZ8+fVPFeZ9DacDvIkto1rpX3FOGe2vQfuvm9p
M0Im5jlM9QcBGhBLXaDxnvChiJmJxtN5P6BnOr6nudgpfCj0cqFT2uROjedyvjIOa3UHsdbA7U4U
nUg8h094si3VWQdeaeXszQ1JhmGv9p7XKuq55snVFf43hA1mVfrQQEOH+MbdOPrLdOEmbHV4A1ay
TGDXq+04UVQAKyndLcKzT+4/Hrwo8g23fy0Pb42zj5b2yo1d+NJ9i9CKRsV/uPksYjprVGCjsNTn
RkdQ045oHgDQAtsPgEYl5pz3NVrYXSvjlotw4h/k0d7zDoVcagL31mJP7pn+mlMsbZSVTB+fD5Qy
9oMGeVXgCWwfGut1jC3Iffiq+VSwjXxq3Dbn18QNPDVCMRzrF4UbEMucYc67kIUBrPezdXL6kTC2
Zo4qbJZS7OnuMu1XyZX5UdH+QEN3aecUBXq2V4kFegASGz4Nn+CHvDhxM2pTzANDdUGVTkReCd14
YhxdZPdc0oss52IvdICMoC4+g8UTCwYBDG8HFq6syb+zSPpVGEEUt98oSQi4/eIsgL/9ZieV1ThE
Bg7aP64ajXpjBZJWwq+pcjIEBs0dKS2ly7tN2EJwe0DUWilr528JDeJyl3afgK5Ai1I9LIEWSos9
htwL/m0cmp01dMMjBX3hWZG1koXssZRy8UWfKDVIGp5A6lk59Od+YWIVYvjVSccIi73orPybU3PD
YJ4Fo5MIQ7bF8uZFC0laxeDnAUiEM9vRceBRDqdgBbKhL7Jf9l2QJmKYnL/Z4l/EvNTKuEItFuMf
VfD7B8DBuaUIywXjbYVxwq3s6g8e2AvCm20BxuhjapCrbSSYS3b8ZYxh0YP+ztQ1IKV4v5OGy2Bg
mrpxxpdqpt9cyLcSpSVe0TYvQIL70Rw+6wZzI5rbDJEmx/FX3tBIu7oGcO23if66TSXZ5GTsvCPn
/Gi8e9ypSeX9fN1RBLYOF7l+nrDjdmk54ICWJHqcFNn7WElaYSTZI7che6gYfyMVv9QdIijjeOrt
35naavL8dJrJmMDyhn6lA/+yFo4rx2f5Us03N8iwiGm4zsUWaONpcVyWizaZrao/hoqxSAiSpcq+
hMurVYTEEOzDB2ar0ut6vF+53SaInGw+SX+Zm9gnwdd5cQtc9JMNVcBnyloI4EecU52qGznWOYQ2
hKilUFIyxsK9cWmgvP6vHKf5v+pL0gjBiCeXtRLFaIi6tUO0JKEuzD+hj27gxs+l5mSwPgf5/D7j
IHTttexhqrAt4Crkx3K8xyewvK2FJKqOvoqhI2YJd4ySQtrzrt8M5KhGT/Pq8PKslAuqJv5rkNDA
w3T/eDDETHdX80Xw9dlI2OQX2AXtwIRj1WNS/FqkWCvaV1n1vwKFyJ1YaZwYm8AsSHMBG+cse/8K
UgQBpmVEgO1baoQrsR5bDo5GA2RJLdVJBXJECx4wAb3L+g1YNVmEzzl78Uhv0KU1LpOOsHRXoWhE
7CtrL+eikqlxhlcVA/9CWz1YFtikOs097mhmqS3NEBmC/AhlMlye/e401az/5h7j2GGxhlvQxwhC
cXSsiCmZFyoAYp7i6rneNzQ1ln2I9aKoiXQVXh2Ti9eALN03g7+VUC6T+lGuIWwvOzgyFGKjTUAy
nRr9Docb8NtuoUkTlm1yFwdr5iZ4bYoziHStlTt0U4p53hq7r+vRLjZrGpq7yMyvKHhROaoEX14m
N1T4qYNURG9RJ7OneI9oT86hNTYp+C4wiAx6zDgwH3BexKoJpPKTlTGE5e0DOF+SkkvhFN+nwh0l
VRWee2u5LS1vr9LOQaaYGZVUVOVL/M1wNA7Mt0StyQmTQrZfQPAPIs4x8gYfyGAqsz5pOWGFIvrv
NafLhovqY+phUUE74lmEFaduxd5uSNhnQvuqbATi7Y5Qiz0WTfPI4C19scA6Wl8dCwZUhekuMWBc
k3I0oQRpU2t+73RVFEe6RGDgF9QtJdIMJeaosdJiYhrpqA8v/Z5PTSDgBYjJ4OuHGfNQ0URDUfoh
KUDcuQYElgWONCWkz773CCnlObBJap0vedvttL464YhoZSiumzkL/guaxK+hJeKmkEHL6E029opX
hSUa+Sfbw5fTJdEEU/k1rX6wC+29Cax0Rfo9sb1j2B7tGf0odUY88B/IY5WvpsW7cuijCOOM7VDQ
4kpkZDlHDqDF/4qOuTIcNh0E1ZDVfpLcMJJjWy+HbVKNEzJJdcgQCjxAX6RNGRwgIdc2cAaYhRYj
fZYwsjriiiTgGpktxSoZreipvmivCSeQbODoV9OcsVAzUvfBJgvzy+mXAN8Ct1GA/hby4C/DTTcf
KKmIL1BYiZoY/GvoJkoKmIBfwp+SmR/4eF5DUnSgRpD7DTrFHOhZh/onhT0D1l9mKogFO5sYDNcH
KiaAxnALfbbRBEM1JRn9/tUQg41UbGEqU7e+Lpgd9TzjreOKsmT9NfV8+B/420nTS2mkQEOlE6Ay
kiWdvTIl0atQZi93++/CRHMxz5P5fmHPO4P1PZM7p2/yVriUzl3xZZQwMVtoRjGaU2izwi2Aso1g
bISsUM+Ln89Umh0a8OYEEl56NjKjR09Ljf4pmwlo27wFgDJGnVO7ChxSIMS1GNwXDX7Z6o9ehn2W
vtyH+zMwgua/B8T8AyWBWXLCWtVNxe0ENUA7P+0o3tbGLAl2YLa593Hy3ys8y9aouPL4cAbLHLYh
ex+SYOxfb+rDUPDMx95JfJkKa615B0+5bVAPDeEPl2ilv+T4iv7cwhnEQotM5REGdPo1o6GvaqaP
xu163vOkcWuiBBSV1p0KoH9yhxHwMUGOf2gZ7CJwKJ6gQz+Z8ETYauJk/P2TW5lDpopYlVleUs2Z
ZDzf+4iJANCLabf1943CfP4e1Cn2wx6MgNvoXYWfokrzXH7kif8lRz8ZFanwJhIZHvxdFySQQxsA
ox3nVGse/KvXKTzMPoDKiY5qFd3k1XH45zxGq7DDaZXF/Djyrs55zSxhptFNKBhq2Ryq85pQ3Tt7
h0NsXaZ1hctN139NOVKA1HZ8dCMdyy446lxijl3xQf7n1wwvYLlV1FN8WJGc+09ghk8m+aB1dWkf
cc5a6w7qBO2VRpcbf7Mv/4CDTz2x83yvtmxNjpEAUK7vgaXaGkrlVvg2Zwm/cacxI8APgBn06f0a
OVYXo0Q2haRqzmxqDemFQzsG9XplUih7U3CYQ4cwRnSlPHh3I1e8VtnfVz4q7iUQ1Uk9IjdLfpZ1
ZW9rBB4RjPVlPp7yLkD+bazluwY413Sdvadc5qNosug+jsiEcmDd1rEDk5qKq8I38nk/q6/i8SlG
QtG/yKUXVZ0gbMrahze3vZz4muKX5owA/CdrvZOzY1W5EwcuniZYnYzT/iEKVXXxGB1Uk2W1RGm+
Vmet30CWMxADWYLvud7Q96POlYM69O8+NK/xm5PZvKBV9M1+oiuGNi9GlHdAaaNibE5zefhvP0CF
fvxohysZ8E02FtCfxlYiF6kqukBXAm8+gOr7aYrRlqUbrvViEu9lPMR2bFJiPTnU/vxibczwiCHd
uN7I8W1ZX73SCRosdUdlP+E9G6OadGvGitLrF1mrLdjk33tpVenTDNkdCuE7e42FUUw96CBxrwei
lbHGjQbtQYP2Kqh2qr5w68OCdypYhkWWy0NXsLWLeMRcIW7G0Yzi4GrHvYtTFA/obV5KOMlRDCmL
GAUQ2wh52V2bImcqzdQbNIVNH/tbZhNbvxQhwG3/jUI/gZhnPXQma0jIP1FFmNS9sEsXOZVQgEzr
umbZHOG4812BCT8yVe7wUvIUqWtpDbK/o1B/Z+XAuWWZcMSl6899fBdtkNIrKiDV+t2GovoApVgU
SmiQ0/JmX14lP3/3eFA6YUSV0diGc9GQL7s7g0PwCYtkD8n+OYE+CLp0s8JgXrmaEklJQ4f4budR
pD8zScwUaLmByKPoKDvBdFZeDTiR+KTfRJtJ6YPzpR0wuxzz4Qg6XBQc7FLI5xIHcMdcTfLykeGp
leyKbxOBqIhfJQs9tPh+Wniiwhntz2wBFgm7mKqtYPJfYTK5KFdkPfg+94hr5tlTtwMa7risY43x
AIp40yp/0deNx9DRWVVZ31269eE77LW+sYloIsFMzt/JysVIQOH4wRcIe171j0qwEiay1CqIHc0D
LpFSzkXXT8RiypRz5GLn6RGt/Wj6kKIyuMjWRQ1YQ97D6Ipy78EvlF75SHWS7r4jbYWK3w76aN3o
Xwcyd2Ct3M15awopNGZ1U+eKs9MT14vdLFxdyG8EEFcEZHbzOKRF94k2xFRm5r2uHA1YQYjOEJHU
KCkzUWMTK+Kt5t17k9YzA9ymjr+Q/0VQoxJfsgzhbfA2xpYQ2YSCFg2pu21Sr/K39sYMDv/lp86N
RwU2iLbVL9YpeRdaLMo3GNda3f8CxS7eMtcoTnzRcuDqbzhUxyL9BfGgi8PRKu3iYzo//+rUC8Gg
YgRf9hjXnIHCHfYQJIkyZ/KRi5OH4OQB6mHXPSLwKpXykz5ztECS4/MJtp5cWjs+ofar8RToj9zT
98C5up7dir/H4tCEPnGRAY1o1AJs11wxKJHYFmqgBux+Gfnn5VR1ExKVjEDU2iRe+pqDqOqEzOgY
geuxBD4TslnYdbNauIzjH29CfQ14IKBQPEuf0djdkkOyPOpJR9Rtyf3HuYPmHGujM8QZErorC4GT
Kfps6Zpkflo5qzGxWrz6GllJpt0ui1helD14I0Y+m67Sc9WezoJmMFtPYOTb5gDkbQs5SUKeJiTn
T15o1d05sfsXtsTuF9U6iRi2jWtFqtMD1w6AyQVtMh3284/PLi6GPPyia3dvYWfkOuYIe7KOfz83
K5E+vaAdm5/EJftR/G0iCoHIw7NNyOpNKiz2ePK17RPEy+G/BGENp46sp3ozlaw5b9qvEFU2D7vg
RuWFKAbiS3gkBoNa9p/fegfh2WHBB+Rj7Fgm7t8p/wpJvUn0bXnaCA5cT590xZyOUMkOaL1uNVRC
PDT8IB9I2EaAlxh2rvumGCPB67OqWomfGRsKzU3+CBfJJOweBWBjphYAC403C4lA9Et9vPkVOQcu
RPqo53QTix4n2U2fXMEDddJTczsmIZ51vYWzgYU02Zi5eyK2qUIW3myvfXGz1aqnm9Pzs8KrdM/4
Gdxh6vEBUeRZeHx6pK7NjbPoVD1EUT1HACWO5OvU1/INLo2vv08yiYURHgjmyZpKEPnRYRalvnwq
3th3pW6bpgQdZTo7GpE79Y9I9pWei8GRimResT5+1APcRy54GyhrhgkxemfB4DWuJkmCbvcXxZrh
yBMX4nZ4R/POWtfx16Nb+jNHY+Xu+L4raFjXjdKSmnDFgtw+z1M4uJgPwJ45/b07szLaq3cGtfPB
jN90hbnCt6NlGBTqUHWBOrGpOBHb4VhR3caME1CW2/S8SbDPvFM8hcTK3oe+v8wrKecR/dnskPqv
RuJDMICnOVhCc7eMGbFSf+7k0hwL1CScldy5Fj6YMOfqufhvEwxQCJ9f5FuVnfxqqe8/N0iygVAL
jF9KTSQHTCa4YEuxnW6rstaekXeE6g3woj4UsanLKjYDElMI0zX01DHDt4wlF9Onrjl3wK0xU+DF
uXDQb5TnF8CapEbdvKPHNs2N9FPfURiKSbu2EEs1iLf2e8eGLxzQTmEyO3YNaZpuppZBC2RnYb9m
nsEUWU2zVb3YdCoUwJap1sn3+54n8hPrN2QWJSH4glQhJY1C02u6E8XfvndBwEluu5S8aliYnLiV
wJeGvbgrPv9fh7WWAi92trD0ZtfYJKMex/Bi7FXD1+1akqw54RniQB32C6QM2RFXtiKk0EAWR6Cc
um/xQjuw6Dte6G+Y9zsiVRIyvSWQQ0qBw/az0jyTqjm3aniec+bsQcaSedxhE28zgraRERSOQddy
lk66cfFRFGO86begh9RFo0DSdxZ0+6amMomL/O96xcoJWB9ZVUU5bWS2hCWqcjOJf/47r9fLyZxf
lokVDe3RkGtycackO4at8+ZpoCAlKTNSb3LqqGeJ33AqN4nDn/7xiHgxeNXNqyIyS5byB0Dfs1Ac
q2k+hMgDGQplkPW7R890NzfXY1DsSEHBOadMEBWdM6tMJAMlGT3vNdUrFAxQLft8MkxZVCHbNxhX
WhFDfTcEwJG69d0Ecb3aj7uKNbh//8hdHxscF0MyhRAf9/rBGVCQDohnS8w1cDsmny9JucnTJKxj
RAxafPSfbUfZCYOGIkkJILXC90fh1r/DmcRgg66MRGJ+QoHP+xyimYfqxYU5UaiHvGN8vqWuHUTB
LJbXY2BeM94fIQb0m8wLhgYvJrWY5RTIfwNdoHWxb09FCqYBZKQGLTz4n9sDMZ7oTiNz1HTDb+2z
iZPdig79W3xfkbxXktm8nH3g+5ixXgPD8XVzAsnPYzUl221PiiEZnpHz9QSJcGUfsIDmghDEcOmh
3oZeet07ptMAdvrjQ2S4jsH492UX+xofYMz++ne5wDsEeSJOsi6DQgRTfd+6iVfPTnxg+Sm4kyLa
VTOuGtS5nJOL/ej6K6N03aJroIJlFF4w19zk1XhXf8sVdW9TcK/YB8kGkLgw6C2LDN06r+O2+A0u
bNmuBTgzx2f9M5fVmsgw8hbjqYCpLm9oYoZx+RhJ2KcQY0ETAnJJIRkt2lgX5mrj2MHSgQUcXeru
xkIgKXZqC/dMX+5bMTGxDduk9l4l2UqQLFjLtm/1MpQWDkgemy/zl9De1MexJ++cOaxUr/jCG+gt
DWljpEqIo4aCBCX6AZeKehcULz1vTzAqKhzd0KSu4On2ClLxgOuiFZFqRDihLiOOo3+l/X6oHcsG
2Ibp73rHO7lxwYWdCJWj6G15eH3dbh3ivDykWQyyN7UCd+93VBgfTiBjaR+5kbN/ToESmiP0NyiI
hKjModrKY3O7ssiOPe3X4oT7O8gpxafHdkNOmP65yARL3Y/Q6O9Ff0a1kJodL5FAyfSpESxl5Bur
SXJ8F1Wa+9h+2ayx4e7fFqWtHhXzhlymZggJgBrnCzSvssjkrKmkuF/No8qlCnmq435uytf26Ay+
q7xFsLJ0aaqieeiqYGHR9wyJddvI8ETI82syDMeAPQIPdw+TIB0vSVoeP9CxUUMlJSFEVnuBMJ+P
F6lKBoQLhytcRn0Fixy2U0ounjcJeLZwF+2d0CQcOfya6uscGzKaSGoOrrrHoo4n6Qpvkd87hNjC
Xnf445b8IX2egQQFxELrDZ0peh5yf1uWH3uE4WLoYa7xU85ZMkMU+k5/DDIyF4Eu0qd4KHnoJElq
It28AAN/OzRuqtRkdgHNh/duGjfxDe3F5k3/tESD+/bE6oxLOW+wT9uYUHdSCN0oE91jsx+9rJbX
TXt2N1iwH2aoSl024d5RoB24v7i1nGHD6upHwOabAJgEEtTKMJlo+x/S1tT+90N+OxjOTrCVkFKY
R9Msf3Y/Uvj/6Skg04ouCE9YMtsOr2EcKikvyahpBFbayKURl42yxgquc+nRTzx9WQzrnI533h5C
0lqZwZL1t/ST7EEWFIKW2t49weV505vqCrZnzrDDr3/Wn4j7SA9oV03477j3fImD9N2gPTnitXXt
ta2DiLmDSbcrptcCmeTDVLioZwUH/B/I9vGRIajiR8zF5YBcKcIpcNF71z1NR+v0Bc4OwHaBsc93
PXXyV5d5A/wW0dp/yj89TpLz7cCWsqNu7qevD0xR4xzDsk3A/olIf+pfCm/vO5C5TguW8wbvekpU
1K4MhhGIIN+oJI6yt1AfBlWe0NyeqvVMqSlRR+j2Ve4AxA5D0QMG69H8gI4sl01zQ9g5PRS4sWVU
530bi1+EVnDZDDpM73wC3KBPI7QYyNzogeQX+h4+1zLoRdlukFCzGEk1CH72GFFLllRgT0xCr8CT
fTQvEZr0tuohTEVmsywAWqkiqgfQ+1dLntik5kNyZptgANElbkH0G1fB36CYPNeAEeN38NBgTi4w
uTC5gNe1AMyo3mNwdadLpVsRn5mG12R1tZzgL7YB2gRl+tTtAw6hcJnMtI78l9nZKV1fKxYIUprZ
t5P31el2ma+PhXY48wwfsl1ZXIAxwTwqsClDjhmcIoekMOmgY4Y1xn2Uk3eNGV6nHBBeKvGy9WVr
z2F9UDPuKEiZIJzBBS/z922Z99ET7w+az4xLkDGRwD4yDj4nHIcgf+qIBhvs9SHRdiWruxP0i1CQ
+lJUMEiq+l51SV3uQaQK6QKYUaQYg3EarNYgs7hwnc4n3Jr/FrU+kaaiELxG7N8OeX/GDO1+65bu
1OgA4SVKb5BrDoov3Ek04JPaCp9ff/z3jsn9YX5IvUlG21AmPUH7X3xTpY82xYAEE90fZgB2wPkV
oD9H03Y9B+o7WyPJGUKxUK8y3CPD0Zhy0wDI5WSGmjL04t9AzONub+upLKP8JZ/LgjSsN4l5+K78
QTA1+IdoYOL8pT16uekYa0A/tcx9ICu6WUKyAIhpzshB+0yGbe8aOgCp7SPjkT3YuEqMPeY2S72l
6SoraRRPzGl81UMnfsRMjR/IXJfkABUYV+iDmsPoaYULyQcUTMln0uVWxISPctBZ1BA557zdfXNX
qfh2Z8YgFrW2DxQtTW0AKmBFn3+eRVs0pEGi2EPEKuVA/o+IQEKFJ/Qyi3TaoFi9nG3ojcO+7Hh2
rbZQqYyb+UA5usvgqKOC62D7QUszmsN06Ui/Zez5boKWGX6wInwGzgg2NVKwMaLIZ6oLkmE/EvwL
5IjslZJW1NflXByiWx7rSs7EUXoN+fFrEghjhdR9iRooh7cz8SNzXnVP8u99w1kfeNgifH5tWU4J
1XVhPJ79Yk8pQfU0gRyUjZjPtiw3JALBLp1KCJs51P5AilJiQDlGMOr4WczjESGq6TGmC2vC8CNd
O0c4RV215HKwk5Jr2dQDGwgPgXXOXKyoTAIOHLNTytYDpUae/adHTiSrfYbaDqpK5uHJM+PfeS/u
v5TmgoIG2M+7jfPbz6NNk96F8PJiA1ACv2GUNtM51f0XRO5n4fS15z/FfJR7SI0Y80OFt+0HAaln
C0YZVIz4OkDYls1Io6W7y0LEWlVcrlLLyWvLnJy+lB4JwRB1//3PF25tXrcKFdzWRxxXmv8Ublv/
wvh0gZjfEOTFMntdwkNNx8NvZrtdR/mdiQfaAjEM410hT5IoslfyIoBepQyl9v1JvEzasNOp6aj6
PXxtaqli8W3tYUxXE71CP3tBIZ4bUcVC5QFku5qcVB8lnYD+oDE4zV0qDREjEAB1IUCH1RGpvwl6
pGq7TNVEfJ9LCPsGwhAAWlbkYMvUWFCZvsF68FrjC2REDV77LpumjosbjdTw0MK6sw58zJDoninw
44XT9bmNaf83Gjl/Mgzloq8qtNukFQ0l3J5V2iLJlnjdv1y8f0SJawbvSu8MnEDp/QpEkGuUGuOo
hYuMYWKPHz6V4eucUYbMPoEUdum8akOy36VfrHgWhEMEbLCI9JfndAREj73GtkmvtgSFh4M9MbZ7
VGLUKAULP6eHn9RR87ZTSAfQHXBZzae8nsVtSMp+jcJLVT7KvoKHG5K7SZ8/eXjY6RUM9lohcpg7
HcFvWlGuWXsIB7+eBdpBDpepcPU/52XXqfB2KltmiMrjKhYFvYeiqpEHujTiSnC4US221P1F0fB0
33AeTCY+5P/7N8lrqtTa19uT6O+fZ48/4V3L2uX9ynRznMdL0qrRS0l66oQRoV1dC91OA3PMUGGN
DSaFMzqh7VtC5tYAfEyr3KoDWGhnqPYvJsQfXZgQHEzHq/YTxj4awgIvjKNGX+/i4I5B+uHwDM0v
ao6/bVApDE1+295xbobFJqyMGR4C9jExpzIapsFV2JsDzb4l8nVeD1CpDztrL/tPzqH3ivwkDiS9
AuMiNwMJVZ6OEotayAo+/dOW2iSuiqJnQlTE3kzuJkaP7qZQlkuSa3pUIshwUW82S7h0hwpwW8zy
WXBUrJkd+aT/vhK2lNkwBbmcBI5D4h7ZoaEC2XhMewCXWXqYz3wy/YDJoB44mJXlbUEnsb/yU7h8
dmaLE7bjkam24qSR0G/M1dO+inqviBNXTnOpbJtjaqWF/j41P0hQvHr7ETUW+yrztMjB63Moruh5
rYIf2vZyoQDZi7/I41A51CrPEjRu9zt1+4n51DoqK1gzAfSAIDlAvdBLK0xx1W7hY3DJrPF6xMDD
oF/5vZxt6qQK9oHtXCkSrM4CQylzaywXMSQCi4S7XQgetem8Ye3aFxNzmHJ+u/snJ1AFGtkBTFIa
CR8PeX1Zjel+p9KCH3qdbCUEUEri3QVrVRzvfXZorSUmxOSl8EpiZt+LCHjuhMWH0uo1tTh16wjq
8+YTb2uZNiqY4AUS8rStKdId7glZvLXUzmHtFECbUm3wNLb/PjziwT/jgULu5CuuM60G1+R9rOwz
NfOM0yu8NnaJSaCpjahkycLZC+krgVLTnkGvakoFv7yBacISlhbPMt0kErXdw5ug/r6i94o74wE0
dRrT9LPz3Tj5pN6Xl7RS0RqQpdocea6lgM+iP4cUhzNqOh53jDlo4FvQRkhqVI5wJVJToIB647aD
jLzaIO3ecpXgPok4qEU217yL4Rg3B5O3nyVJIlMDj14v8mVVbJwW/Uh7R7TZ0W80W291AiVGO101
LWHx0MMhb/UNUg4n0dvYX+gd5b/l7RfopKDtvi24Bo/DgnJDy16S4iJUe1vdWS3z6OZ1VaifYN4+
hMT8mf8aGuriFuQf08shtTmE0XATsePsHNi7+b/xOm0WxrenCIyMZDf7IO2yvTgJNGseiYUgu+pi
cQjMk5Fb4IOedEGzXh6X4+Xdfqx/WmJtMUGP0nKD/IQylLIrFjEr3Baf0+8ljnptlJpDzjicGJ07
qNV6ZpDjBj872+/iSpXRDBiKeww8mgS6s2zkUzjD7RXLbFhdEVyj4Xi3JMTDyT1i5xlix1BtXJRC
LTcYv+d5kVPuIBsJU7iz7r1bez+yzZcsAog/FLSsEqDg8B41bqhQDIxaqr9wPOxT0nKngrRn85rQ
9r3kjU/ce6qwQxEjkQmnQpzTgZZyf2J3EMPUrwpdIEhywn5zq3tjWWb6XGs/l+FmzM78WFJJyrx3
OFQLjx5+XJdooCtn4Dp6uK3BleyXqk5FOQ1QAfjYnm4IV/TnODCFNwE9Ox+caf8bUST4QfiJF92t
yN3x9n1cshRvqrQfxWJwNKx3WZKEP21anaA1ODb3TuNsCHOdJr27lK4aTSYh06s5GXRCBdQYMIwW
+55Grm9GAwnkUB7pMYA/hiJFMGpEbiOOz0wMmTwbuu2rgRwXNhDv8+kUViZ+GgsrArtzzhWmiqAB
8gXxMJRm7t4Za/CsN2Xjj5CwToWOJyEcwsRafIjuCX7Ketq4NJsiN+wX7Q4HANMRc1eIPHo0Fmne
OomyEEVxgTRPPxLW8qVrB3ziSsu317JnRyKG2GlVczGse0DVlKS91nzWdhG09BBK96Hm4uamS54L
O3Q5nqCfNgnTI/EFman7kDICUtgejILEF7day8c7pyg5U0gm1QlalXk5T/3mV2vWSba19eR44hYH
XHAW4H9dn/Hl/td6HTxTgo95/JF6DmpCQIbK2vnV2GTA2K0rFRglIxR8mGFJYYNWd0ZS95/YLMdI
FmUCVoDPPtzWh2GzdX+CREyrFdUM5cVfFsgLEJZN5qaCaGPkFR5ODQgXtHnzVy+XOwj+shwPoqMQ
S1yG6ZJdj1AuA5kxLnEl+2zimPx3DjWRt67yKBYaZV20auvEXU4UT9tZIjCKGqKQTrY2LTJGln3R
ccMBDItdvg0THAgNFzZuSZFmMniJmm1JHOm2jJlbkhRwrt4Wi6nAk7o9ajCKyNk9EAmtc5lPyMtO
PV5D3MCoGObDNbaOnC57SRypFKGpsPF+3siGFAZ2AmLNAusoQJpS0D8tzqttwfZ9pWMZB5W8x5+P
iz47+8TP0VXQOpUZqKRTwivAEW8D5qOUgmetIqTbW3SSfpEoTDWoLe2Id3UDw0+lm6Nv5+J+bEhR
QvGo2W+KbOxwu4ppK5MX8/slXAmJhrj66NsgcsloDd+JM4e8+WL/D7MDtlnatldzINScMOPM2//F
JLUwzV/SX45TcrkbdJoqGpIZbUAyK6m4s/c4OY+7APBE/3sHCqZ76oboCw479iWssjGzOasGpV80
x7hl4xqTlywmTIBIXu15pdT0e+srZdNBRbnecSSCM3jIhlvEWmMnA03n1GxmfrMd87ZYiOSI2sh5
op5y6jL+COVwS9WMr17SpmkDlYYkvJXfambGMn6049DSuBuo+2idMdxk8LmaaYxFbkxSuuBsgwwD
orV+Bt35GbsbIO/j145NX1DG/G72ZPQQXylSiKsJcyqpdtnVchdWi1aDb2fVy4a+UEbnQS8JDxpq
StbCmqMmeG+GICKSQy7+Nlw/Bp/h10UVmwMnMHQZYwnQsijWd8/b3iO3FbzZG85V1HDfYYv+k7aA
PZ4bRtkNYZ9UMW68LtHmDL7oh2TnjVLtx1P+B1QjsNL8gzOxNWdRM++8hCPKk2iTRzt1EgWjrF3y
X8pqLv5/AvGp2kQjO55FverqvLAtJMQW1BgS1v+Qj/6imu6ZiQ75jD6PyEGrylEFfcIbkSCmZJyE
UMz9xtL0dIZyWTMw4SlbuKdIOBZ9J469fcA8R9N18RhyxKo1z+Oqcvg3DlWu7g09talXiNjE+3OH
jEj8P2NlE8mLgxOsubBT6WLsK9vuDbHYmtRK1QlC38TXFxYLg461Y4aftWDbRlIageDWgYoAGOty
UccWB0CGsPP1NQzZH8gbyrpqzdUVQoGs7UAkgo4/AfoSy8IOlEzqTKCF4OoXJIipmJJ0TJ+20/K9
dooOKJR5HIEgaHUDxwaiD8So8YX0i5C0xV3xxGI8DXz7eC5NbgJCuA3HNfCusw/KZr87d8CgBIeP
2Hp/e6J8vEiwoUsRAosJaMU53QCQMXseyIbN5kugJXE7giil3VVS6ArXM13CKGpgOrJ3KZWuCIOa
vvQAAtNgnqEDA+AELRv/1zlJHCxfgj5Nh+WWz6YvPvyXF7VQDf9RdAbKjQKchFCRWsu5ko7iMjs4
Fd+207OH3sEq+oalBP7X/xhB2lYtUbVasxg03iOEywyXRrBK1l+Tq5FSg8tG5loxdSMLbGSlh2uC
rzmBb9P0pE61iHtZCwxTSZla3yS01PowwqMshJBJy3FPkCre5q/oVUBjbQMyEOWKYNubhXUBuIX4
8iM/prC3R3wN5sKVBQn+N7NfdSGbRO6sumfocnMNC1N0FEoRdD/5sRZYicd+bOR3n25MdZmSlcUy
MppNz2apqC6SW7tMtYlFzDGFKCz68G+En5wQjlHGWuLVO9+/tLsAEZS9zgE6iAD9ByvH0h3zKjHu
prjgs7TZRVMF/fHM5x2bvg5e5NbtoMZ4XSY0twc1AsU1SbjxGZIajM4UcKVeY2DBb4TPxByLtZtf
LQwINHvGv0wtR32uUkPT6NvxVdSbVrhasG96itsoCFnbq36HqkzorS7iXhs98l8iktDCh/JuRiys
LmOnLxAgEWXZTAvbgGAg/A/2TRgPyKJ0ZAlYdALQ1fDL1W5yCxTVkGLBICgOnNfjlxiMcRHrHAqf
cP6sTXKF6ZfzJc1QClfnBG02Ihg9JlXh2p0mrvNQ5wHN1klqszSNEvEG+jJbQrH2aNLZIXC/tF4/
6TovwEmfmL+llBlXhcVmJlsu8KENekMoY549pEDJXYOtMD8NGfMPKhdohAcBupnKKvbfgsjZiuLf
5bUKxXYypRLSIdw62uS08nbRGnY1n1IWL7dW2HoEqZNznQr9gE7yMg5rtcSamLXBzoixuQdllNVC
VuC9rogvF7wDrBMOSiBHf0IOTNQ9JvlALqerP/CftSnb3BbjAu1AeEXhBXc/CiIQ0fHOwz60oxPr
WEARHJUPbX6/o7cQt8EdydxED1SCOB8PjW+V2awucd+shlBOIBzLnP9Vc81QydGqNTIrbMQOdxYk
7syspIQsEts8ydg+FdmdzEsEAr342YgtsJ4vFAPGCa6rnuWqONvifHlvVgl74Qxmu1T5Chmv4ftV
xQAFwpnVrnXwHEVg+dkmm43XRWf4t56VRvBJ3hzCWokzRs37iK17PDVB7F0cp+G4FOPu8nakzASi
KILmxk5X7DN8bwR3sWtpZ3WkjWXydG6sVEygVL8Lp+RfTexE5gksGbkVFZ1bJwVG3u7SIaHqFk/7
TQCM4/ZeiKWp60TgDUdizm/2g1WA1aUoENcK6M5OAIgOO59Ahc2gx17sRaod8pr8wockrr4A/Av6
5YA/KaxQR++/He06aPO/l0sxQfROqhrGe+SUNkK+vQUTa6y2PigiUUPrfx/vVTxz4+3DE8xG7wiD
jXY/008Lk823NzQEd8JNRVdzN9wC8kzo36ndlicCrdBWEFITuedJniaOqJOqZYN+J/WGWAM3Z5GY
43lZY0SeUL4U6haXjCDEWD5UuTpso0MNV/E9hq/7RUSpZuxgI2+IHLeemRqqE7CLU8M2KxhMWhlO
Kq+lgk8dV6Lx6q4f7gya+gdaC5CMMqk1m1NCiB/8g3tA5UpaVy/8lPpJ4R3H4usfiilV9QfYwLR0
Q2teuxZtzGzBKsLGjB83VGvbvdZIyzajWRc3IcLboRNE0WIDIY+GvPGPqLMq4U+0wt+v472pAsjZ
M6doQRkmevg8wZvWx9fl//H3fl1BCGh5ghZGUSRRFUKSCy5zDdzXkkV8QoeyTDhxAUH0tOe/Jqvs
VMSEMH0lhG8TwtQaXdg4LsrzxDgUTh0hrsg7U9sFNnya3X3AM4TDc6D53mie4QjJ99sb0xj2nz43
a7fiLgeAPFrSXMwboi79/c1oeFGAUj5s/rPXNKSfo+IWthWTe+kTj0QAEDjAutrvA8j5iX6OefZ+
iK/05ZExjeNEfQlMWLkzNAZYPSIVkWtvAg8oizxK0hSQnhTklRgRleKeuOKBOHngVQFv121KFU3S
LZTgX87op5ELKdmgGFp0nTdFAz+EpFq+ZbTwDve726QBZTq2K6QCqoPnM52FKN/DuUTWCMk7GCwP
gi+j2KEZDB1SCbtbvL3zqMqt8c5EbYSycFKsjVSfPO+ZSIj4WJ0BHHUXULq9D4f870omg3Wb+xli
B+hl0tAS7gvfyRnfMmKbNDqOiwOTdqDl67PMWiNhmfRL2W+n/NkTZvVijU71DyQ1vK/7W4DfeWQr
J3SAUWIXU59YAVoNXhlyKGERfc+byOkyBm4/1Q5BYfBF3yTmx+VboKWnseA4j0MDXMoRPS3uREDH
2gn98nYzZ0wKkQLZO/IAGIuKx3Yf7V198Qx1C1hCxmOVqahQBTSLyhXvi4P4OOoJlFeiihtEZknc
WmJLJX3HfSXN+K2vYkH7NpB/QKONENhvg3To4P+7Eh5cAWaysHlAPhampRPdH7pAiXZKYCqjRivL
AijQlOw0uRxJOxDu2znidPvreIKmcMhpfTTohgy2GF5zY9zyUvDJCGGUO7f9F0Ms9owuVyz1vgRD
v3i0AKE3Sd0BdIe1rZXSe47E5KKrQxFutzSfd7RWVIn5/bual7CA/U37kFO69I2PDAloKCJUTxW7
nGFSxGNI1rBi1pANaO3nLLYeNHMave849lk/YLWouN9eg1GsORK7dC/YZcYIFf452/907f6jJGz7
aSiZRWT6/LfsZ2Gs++BcqtEKRYXg7qrm/rBU3mFJjw8FvGSK/9zlaZ74IY9cV2Rj82IckNgnB9Is
OQ6SvyckM6cAFarH2xl3zqFKE8mBWmyhjZ2JKr/lYx1o6xb5TQlGZPCr1W8klSQfwlnVBj7KoFOy
3WXqNFFY9Qu7mGlbrktlurNePVr7/GybTvUr4HmNOsWsoNn/WZOjkAZV4mnsHbFycXR99TLe+QpK
ZP+MR0bW3PiL7Fg4dIn9UenxR+Sb9E9NCj9EY36VzBLXf0ZbR57hIFJ4IPqETzKkYtfmcNUximy0
nQp3F/M6M43TI+vQVX7gad1QmHyVoQ8jTWqb9acuDLiaZdTK5WJFXzaRlOi0Z9n/Vniv/D9wuJfC
H2yiZ39jZgT+VplvR5Jiu+Uf2nC28hmLIBvwl4ZTd+3TuDhL1S0yLSvng8ul/1HAHtPowmtIoJHR
ya+eLCG/bRUVVE//EYanmayMluDqsjFp2/DVXX+nRNeinQyniqrRqvU+TWNQIr6EOJHgy7apetKa
Ab6gUnNId0vVUwxuQ2vkoj9GBtkOMA3bEhCYbUQoepVoSHRQOhEbr7XsALnjpXRORUzhW9bIXqHX
JuNKR/MY4lltE8IP0MWPrL9+YHf9fKr3LrfIYnq597nj2GDVjmRh8whteJSUx9o1f5hrWxNpqORX
16hSQ/0TuY8XHqiMJnGN7DYjn945MlKOHmU/Dnnj+rfHg9WtC1o6Km0rWWpb/JwupD+El1KoCT/N
A75dp0a7XjjOGkP+tCL6wNRkAYxSSyaRokgWJafm2t9EvJLCKKiaccxXFPeU6gmKXl7WRn3kawAk
5sbBxTWdX8jurxuQcq7lE+iAhGDu8FWmLdVwutxi//V6Snp+4NejfmVLJ+5BKO5KrbvudVPvEYod
c7QeyVleZgnGQckwQ6yoIe5+He/9jLamt/5afwVavqXjsxgCxnr2VGQoYHQ2fh9pEQh1gFOURAXp
HtKAd1h4dgdhdLHElLT6MJsibBGr6R1abVqOiKzeenLKuEddHmIrOURSuyd1Cfam42QqPwcCRjnC
xDcowztxVhjU7Cu0M5krf5YJrCvSh2sSDiF5AcfMJombMZnlIrgLGF4ZkjJ3t2nIDE26ZOb5aJpv
aI2s68GIgI2VmLWSAx22yfxczjlr6wQlQRymM1+O7afHW+kuGTa7lkSyoO3jll8yI3viXe4vxLvp
I553wK1Q10jJs2wWXcs+X7nU1Znrs7z5icpZPit78tuveWzMFK/eiqb/S+AN5WAIpUT/TTCDXrnc
jvfPi7URIEa0+4CPCb12IA85Q4kUsQODLjWlPGPhVKHfP2g/oYo2N+yvgLy77h82T7aKqb8GXt1e
DZE+rr0ZoXqKJyELJ/q+KK1IIKUN3B+raHX1MxKAIYeWfedCwb0T3pQ3r1I0NyEgqSjJTbMZKy9F
KyIP0WYvkiEY6Z/Fqb6pR1h5MK89EE8z+kuiBhOgB9mU8JdIXvwbrciD9H257ZA52wYyyGB6T60W
qEvnlRaXCEkeSvkRyY5S55S9wTSLpP0TC+17uh29T4i/5kl7baGYz2Vcww1e4+sOav3U2QHv438V
qIAMKIdUq1+pksxPnAFWB/3ulkAASmnMKQsTOnW9aH0E+fTXLUaoChBXzGBovyodwzFKlwSrHuFP
j8uqN3xmBJc5YRuCy9fBY6Dw0e+18oCKjbETsw0KWWBhFundDjhI1QCBKdzNO/wWN5WdY7u4xwYC
ifi9uw/FcHAdyt+B7zKSAWUFzTbQh3Zix1OpFx+vi3mB893shh/yNUDR84tG4xJ78Rwab2xUeAbg
+b9u4IukftslrP14GMPJUL7WUftaKS6nx52eUFqfNXqSx08mwLV35pCaBiY23W1EBcMpjsTDXyrl
gmFjSBPuGRdwkiantnw5Rri7Zw1oV2/tPJop17r7198NYPcsrYbWQN3A/NDTzJaJ3QK4yVl7+bhs
p3B1L1NZ6q9be5RA8UWUzsun5BkCVTjYcOrvWyeRIAwHLW66kHcjH9OMmr044+641/NhlhHeFKW/
hw2HPiu6ot+mfYn85RGLUKkbbgoXONHKXJM++Fg6SaCdpqkTymjjZRbP0iUI/B0m6DMCiwOMMLPf
/c1SxDOEyTK385kY15wzelIoG49Mb2cHmkPg4EB+TWOGWU+8QhS3WdN60J6EVZc2uGTxKeP1IUd0
X1yvFnrUS834Rq5BpGNnaMM/1BA5SLJ5LrWdwVIyOgapt3NUS+b5STcD6Bp2APQUz1ILlkKlUd4Q
wwEI1f54J+WGZnrA9tbWkBy+pEnFpA2sUcg6j/gLQgnjMFPhCvdHx+KO9gDIOYqnWCGjCquj7Vz4
17Fx2Q8eHBQF4kMjGZ9N6D6JHZcaQRi7EA6+7vyGGawJaWRMnp8WXvPK4Ng5Xu5vVL7N3Wk2TgeP
fovB7UP5U7ZhChhym8XfQbfSUf15LjJ5WYzJxiFaJbuaRrPqSgh7KZfXg00BK/kVs47T3uWuVeX9
p7s8QtCF2O5GZPk95ze/PoCfjK/E/jMAtwG0rM6VXM3Yx/UerxU7CIyp2IWLMezTeZyA1IXEzEO9
5+W5vYb77MJwo1Mt9ETRfx1Y+Tw2Fv92qiR7ooel4M+HLhqnS0fB9QntxO0G1zSQttlf6CGNNdUG
bIvT5wDuJ7hGHV/prlcA8I8hw6Gatp4o5vCw1oKc15tTp3gtgpy6sVkt2+r1vXbPrr+Y1NLUR8qc
tqLQ347LdAsE2+k+FQG+5/CSzHcKt1zKeBxWAk5Ft+XDPFHqa3TJrSfmEvn7kCMTNhuJct9s+mbs
Xu0U3ZDVOJYziqQ3UBzVYCOXG8JANlA1SlJeZm1ZQpy1eAS/wVbvi6QfjIVaXj8chYCYEO+ExBnP
c5N+SNyVZKueGeIm1sbJyD480isR5XUKPHwfrHwK2PsykdsQpo10Bkt7Mrf5Wk1Sjyvg46+DJpag
HTxPNYYvuJi3hISxiMsZlTwUqwFc3LxWN3Vp06ymTvXCPZVAKCf9e1nDJ7Dv1GOGTCI7XpzHKnkT
eXBiBjkpRdjY3xyt9wF9U5po9wgBD/h9rG944HTkFlgXYg+9GZaWy8xZVUaGZJTb5QDHtNUQQJBi
OU4aF4ibbEaxIpJAvzjtiUW63M/t5I/7WxEzdGC1GTkI67hvM0nqQ9cw4XNnxNR7jb1Eo7TMrLYV
VF46bY4jORejkTl1bWd+Q/yP04dDHsS4bh4pi8Xf1YvfF1PZ6vJy7DNOUvgaTLMch188GD2V2VZ7
7tDhQ1Dgb1GKV8hiuvScIZGv2cum6mb2zxMaAenlL1eG8ytPxn3zu8gl1O0kKLQnvtPO37m8Ho2L
wp0ePEdFdUfYNAeP+xjWjOwD7J6P5yWHspPN6H0Ic+MhWbvb7uprzh07Z5JAIThjnbdS4y+3ZHrd
4F0vB9K7Dg0y2rLg0ZsPmoPMHh2fI3+aEsGnYBQ4Is7inw8coljRVidAPve4pEFB5eN4DMVX+sBK
8R6/r/JZoBAM/LJPVTayEkuWN1Gfa2e77Rsu5RgFWwNun56ozNffoHLtnvnJP3G7UUXZw3hNlKEo
BwgMyqaUHvllHFPqk0Seu5ajVBWqxPTHPFQ4BuTgmsd+ql6TNGjb12p6t2jvbUQKE4kk8xz0tndK
BYLM+jyZjkMjM0qHwaafoQSexo41FXQrxn6vrdqtUpWWmm2wegpdQ2zsgOxBhgFNhieJ9OKaCamL
I2kNff+xa0yPMX30mHWrevH0BUdf3TubHMbA5jZ+5vgaZmvlEw2k44geCOJ/uI0txEKoew9WyjHX
tyfMk79k6cP2p5smlnGahYKud2bDW5eRISG7hgyub1r/vTEUsF3n84bMg/so0uZar+MKTmjr7WbH
A3sAGkAZHg6faAv1p7n6AvSDTFSN6h16u9hPP0bKIiERdUy5Mm4JR3hbXUlgLIuXcaXIpnsS7CWF
3zZKkzv7ILi6C4GcUUhUAXeL6ldFHDTMJ3gY99d8hvOk7/sf4dBYcjL7mF5fyXJmSwS3B2SOz19Y
CbZVL7Eyd6YW86u2XM6IpG88KgmMGl5a4pz/Q+QTlQvMMMdWonNhiR2/kot4cj4Rsf4nzTzKHZHT
2EtVY8mNo8nGLFEHkM5VSUTHOGSgjSqkglYIZ0RSdALWDGbVDN9qeWoAOg+BFCbjpoDvYIRzG4Zk
qhVn7YDGTe9aA0QntAU4ACAiOI1tfRT4sXN+MggUmUOcxBjdWrMp1a1Utx7XFk7wIckkgNNmxTrO
Hszny0K8qobkNVX9D7J1sXWKefxvDKv/IQn8hTm+90C8e0a3MCsnqyV6h4SUBE42pFSabfkW+Q6t
mgw1sDRaRaoalUGrR8BxbKHap1OrA+ChEAEa/2ZUhp8K4zTjgUSjzybj5KkastYEUAx8qEqPhD4v
bPDv84iPKoEIF/o3qOlJEJYTjDq34fZp6/M4PiBX0CvyiSBBv7KeZfeObxRNZ0Z1xzvVVx0RN5dC
XG7mxe6Zbu3Yt+fznUyzR+U6MkG5H2hdHu4xAZqwp/B4oH0/KKI8d6x8h/4qnmNMUM9DcmAz7N44
e80sGuY6qOcSc9C9bUBBSiV6aaRWNOOHri2PVKe0hFDoVzaZ/uLj9HIXVBXSrmTdj4f5ulntukbK
4+CpnHZhSlvy6wBJK1P168UAgMiQvs0CW4nldDJ4P4E1elzN7CdCUJ2x56b3FIdy2Ttac1YxFOok
z5VeCnyVK9GNpTQtlEiXcpPOK8uGf4W+r7JmtuHhFFeB8zXhYdIFMw6SrOb7DWnSbbzNmC2UJYHu
jZ+HmtP5a5aBJ+a622SkETMPDNISGWHnsX6nQdLh11iLIAtM65Zn758jjE2F9RcBksqj2vr6Scr6
M0ipGGNGlEkBE/SpQM8xSVMPCPnciBOYvdI2NjaxJwNCqWyqFzXURd0yEKvSVk+j6CZZEMWpc0DX
ehoKllGjtP3nG/Nh8MYxF2mqK1LLxUY90K1kd549hGsstgC926K/bXTQL7rwY8t3rqwnMMXVwgTE
vLehDkwnuDTEF8rO7jAlfc2/uHvez5V/AExn6bog9ehGnLmqphhyfOTO51Nqzg+Um0iGXkubcrE/
hPL9ZwXkvIs0pJHqNhiqQaQzt5vyDB45923CRkYiotFHRytjYuDRrlSCeNIX/Jsf3sDTr70KidpJ
NEnTl14KVROG9uwSjm0aADexKc+BXI2tk8CVth0X3MYRehr/K1iy34ZKA1WJcaiToio1TKYLDuRo
WPzogDhIeUnuzQQ4DP1pc1caKi+k77BzzPmU4qGCz8ZbrMfEsqJn7D80zvRBB7Vl67x6Q1+36GNf
6IMQLQa6OR9qgRO0DoF+IBM3n3U1sUXsfHKFMjI5lxvS9bdP9l1MJ5rens2Xb2BXQSeDb8iAP1iu
bDoDQBi+x6UQgQ+y6CgbnVjC6Oa9VeTapcoC04Gvlw3ZuWqV2YlOnRHSXJXys0nRv0Veza0FwczC
mUpFSaGGhh3ILdmEPhC9+XHnfu1tDduWb4gaBo9Pfesjf4VoEeuVIbXX9kJDvtpLKlX/L/ua89FU
f0qVPazDjMEziNAJohsQfCb8IAlzQFYZIxBgjGyXYXkps6M5EGeXhWY6Kgt1nin9qaElCTJnNfyV
8MfGbXkChKDdTEnLocf8VCpunq0JgUfHkTrjvmcqNcK0C8NpR/1V8TSc/20mZUJNyrPdf1u0cxIy
3Mef720NEMPSNKb+kGfrSKPECpmwdoG2ufiEc8ZhCrnDQ7hQHRXb/6MUkDRVp1TVlCgLvtMdRnTK
Q8q9cs3fsvVY++RBnLBwojduwaHBqwiN+Q/tKqe3iy4cvLuIlkGlfq+7HWTm6TONh3YGTMWuBD3n
I/NKxhS5zXebmDGhHeSH9xyS5EJxIeFPhEQUztDeF/9FzB7zv2xaDseBEG+QZbWozIXyWJXUEmDm
sWFx5d3qKEvhpD6RZ4gF5sUU1A0LuiHSwt+yHXzqpzWTB4ZCStLAAQ0cO/8gNSF+EMKGvMW2qxLd
NpSKlM+XgZj/hfkCwwZT+8sDSEZXonm700jTpqg0d6csknD5jMLh+uIiqc+eT66uqamMLoPFfRuN
7Q3tjVQXWBGsAo2LHLZMgwXUvD4oVYuxW3mydCvFSElApfFWAG8xf3ERCN7kL/BmYGtHXobj6j4d
ggsoTZ8n+84gZfDEfvfij8F3w3nhh7ACdlmsRmXpw/jVq3OHZFwk48zKKcvWhqZix2bUQdY5Sbq2
W7oAeOfsWuk42vZ/4qF2Ua/cP2tTq0iq9Myra4NDiaFpYgGTlBX3rw59AVx0uXuYJEOICTGEXoRj
WY19B4hkC9ibZsJPfH3fFS8y8Ph7eZLeAKg4AmXO8XIjv2T7EWLEmIz3tqE/64iyJhkq+2/RyDqY
D5MVLrUOJj/djryBniq7BnvvFxzErIfupgs7UZPKhf+byzsptmdVBjoT6U7YqHaVOeP8ToA+in5e
fJ0Ji45h5VFDXfLfwX/iZEhE+ytEVFrp7SnSD1tb1y33AtvUzdbqBxfjUQ2jQPR7islmFYVnngnq
lYv1+5i+4BUvCGamBjCJqbxwanJC2S3NZs2O2ibobfK1wEYN01DC2S22oTdRtgmKKyJ4MsDJiEEM
f9Xhrm1cjtTc87+lz9SkK7HyVQhpMKA13OOqquPxnDfTbujXphJw7XEQJ2rumsVQ6VVMN503S499
EL+cOrXKMikrukZj3lD2/u8Oxscev+pBNkeJqxsC6W/F5KsGrmoNTZUBLUlXbsn983X0VpaIJdn4
HWbUigQjt62CK+PqVeEtZozogbDl5WhMOqbFpvxpBFO4rV/YI3Bfxpnqng2JcB/uQ4nAAffpyC8+
EAKYE95cypbLcHpcTU2DDbSx46ZwD8yGHakBtR/T2W3S5CoV5DgAJ9N02/a1S6DL1fYXj5FaxkK6
ZEr8wwzSkzcvKGBxA3FL8i4qVGIKqn+Y/1bHz5sOeRUe7V5eF4cc4Yj5mSFP4xqMGtAmyZC/8jpt
K9rfvo6n/I96ZVtYKHYC2NirM6T6eSLYgCxTDSIGGkoScYoYbkWJiLdhknKmYdP9lc1IOlrrReWQ
Nq9dhThwzcxWLi3zEoudHOcg8W0JsZ81+RhBZ0FpF6VtCa70Uv3fWXMVgTSl6t7cdOOSGVPKbOMw
OAilzUlExFB7dkGYl8gQXsy2A4YFEf2uGvRd7tQtoeNfsEh/HsAZ2CKCBLAZURAE8ez7XCK85W1m
V3XcpV0HTUFLBvcm3S6y+KXYS2qvTIG8q4kO7WesgavuYI5XRIVYB0wcsc3nCdBeMaqIiLLSUDSE
Kux8h+uNsJOxX9c2rFXC2w8mgLaOWNAJWkzNk57SBqqwzqK0j7EYvmEs2faYQSmtSMnZcBEPakeG
P9jo4goOSETAPM7VYOA8yu3I6teWaZs4XWkdQiHfSAWlHO81MekHSQB2Ftk1VwgHEcGL4bOJfLa+
u+Yr9pl/3R3V6kt55WFp6omgoSCF4u2J+apNyIUOKewiFApocmAEj1B4i3WUNjiQE+WYfTU9BKYr
VUI4YSuaVGl0qVVD0BFaNVQHOD+N5k0JQ3EByWDG0hJv1VqylJZBuEO0HcA9WKPG5/LfLwh6VR3O
X5/YnRd0C3n7C91ZyqcVTVHHDX7rluxhwnzPvwapPCPj1W0oe1dkypIhnXHvivCFzqVeGz4W6B1O
IN8M5BCVe//xLMrCSPQim6SFhsxh9Z6DN7ywdGxNDP1qnhPfYURlZQ62+4HJqkE4I8NaHXL53Ksa
IsRW7yopcCHZ5Fgbaihotd9PVxyx/52Xkmh5opsMqjFofCoI/pXlpewNMBlA33L7DY3xq68OR3bF
5Fl34AkHaBjWKPkmTKxex6kp/FE887wF4gQSwlPqB2AcaY+5rj5taomEiSnHwfPmxLiljgrIieJ0
4ucWfJTZuNyy+uv9eYvLmGHDHg1M6qHzarJ+bQyYelWC0WvUa7mL+DbfULYH8gXG0qPM9q8WKXQU
GkHSdmDPzlShdoBZ5asjT+BpidV0Op2yP/hGD2SMV7EYAflzg5vA/nXoH9onCtkgKM5hkdqYEYii
bZB7oRxbvsFq5MB32wYFzjjmsIPExXiJDycflsrXR+cnd2f7L86gDUUtmyEv6UUx2YFFHzOYHoem
gLkZm+rviTZgo6KSlzvAhdMSfH/lh/zUmFVdYOPSWqsZeD/FCU474dI16CsjULy/1fKzZYUnO7Vr
8lkKTad35LDz4VlUwgUazJjcMrgMTzIFfWPQKT+SU82tFEG8Ny8YSdNQ62ClDeu5HdrGLQ3D/ZRf
kAv9p1L1YY8/IQatQ86SZ2NBaDoShS5kfB3piFVZNpficKO9V3giNNl7Q8U+0f1axvUr2ktnzk5e
nc4l14qqxYiOCSacHqiXu8D/9PWjnLjzrvPhqqWTU2o6PGfxHABsGSaW0wmur4CMhEXlL+lNqLtL
7zUMrpG7OaRAQ6cu2uHuTe44aIakRDUHWmj5cRlxaBAURLNXyX5TzPZSNqn3W9teKIYw9npj4+YZ
sFVBrrcFGTyxKoFt/Xk1CZrCdfvPYlzff8tKFB4vSTifrrkAFqAhPaWIt1INrUjICeVkHH/AURZl
QpkGXjYbZB/h5ZcCSdZIr1TrqXlKyhckHmkbbyPm54oQd2x65dj94qQMSGAkTzU2E+DwOqwL8kWB
wuS8+k/w7tB7qtmTbwXJnCJgDMzDK57YHY4NXwIgZvqTgT/aDYwaaAdqsaL0kBYeDTUL1cCRRtbw
OYz7JpIIcEAqn0Ik27ICHYEpUjIrRM7PcjJQjTnKcUTPcxzkriruj2lUfmpONm8sS1DwCaPxqTIb
L0d8f3N9zsKeaCtwBKAEuzUFuRDjTWnTeu3wzv5D1af4pczldjhyduYZraqb0ApkBagnFOH8zpoE
BtkbGTKibB2I8UIYkf+UgNhoDycteGa9j0vOrb31G18xyv0fe4tt/VKCi/NKTSGWN83w4t1KaF6t
dJijWEYqV9WiEoCZz4PpLQISgtaEbWkesrgYMQsyCL4xoVZ0IefYvFg4BEWWYLpVVEGczGhRQK49
8Ooo0k6F1yGISj56cwDfoHgeaC7saCEFtvoffujdMLNTHQP52c3YiHHlLTO5vAI6bLexne1JyVz5
cABDGkkhph8o9QfZw46Fjiv7vjoDdf2TyN0ZGQ2HZplYqWK7rYnVRIINcmwMXAFqjKEilYYS5Yex
rR2mtI+8CSi4qq01mGrBzJUnsZYwzCyUUSeyluQLJA+3kWgZT16cjM2cECGsmVsuIlWEM17WBryP
kB5BasH633FT+siKf0r7kzocxsCRwNBpTOEePcXWaX2S3BC6FOPKzfpGr6ydlzkgmmw8m9dRsb16
T6hdoRV0cy8wsbFHvXxrRqoARIs2swXG+bCQ3TVzunXu2EHKaAWpb6pcuzPBJn8MYARNRpHwVchv
e0ZVA+zZ90fZJcTPrX8biP/lfMoZcf7sla7IylC8qeS6kvED/JmOZ0VyNJuoBs91bVoti7SQb4lP
IzZ42fSFvF6wPcmJtg6x+BCEHg+8DBWYU6e5VEOobOItj5a4dGnIfL9tDEANtcMrvPPI37olLkIV
LKbo9mMjpdARThzcoYCIjpdx5WCKU6B0xQIncf1mgQRrTIjUqQxWH2SwgWMbBrdVpNcqQ/MlA7L9
t7Yhj0EnYrJ+MHTrnRuj/lKGtIsDedAyXy8bmSeQzuTkhOUEZLqzSH+Tgo4JkEa9OwDSgcwBQk9S
oUxFTKkfW9xENJs6AdbJtmw6gzz3cbtqGbMeN53xIdSkouY7yaEldmOpCr/EFusfrYUD7YZ+ESQx
g2WNE8sa5l0mLT6FAH2BvvaTUxG4WK+FYPGzfPP/8+8n1/JAgFJwDmz4KRwvbTiqmOGin0+g7W1R
te8Mkv4JP5ybcQihwsI+6pVWLt5YoB0qEoGrsoSD0DhzH86AKECCVT+zOxh8u5rLt7fpB0e58CQO
jdPsugssdtVvnqZA9QOcbLolXdroFsedoF2hNaXaFpMAi09Kvr96XvRa3E9u0dTOFKFSikIcocaP
L5WR/kAvF5cvtDPfTTrqB2sDZr5j2KSqex6P/t9/IT03urwFe6M+Y6liWrkVEU5plfsrL/dRTPlP
pv9s6UdoCzNhBMiCSZGnxITIguRQgLI69KptmbyERp5NHm1TufilXMOMcBgSf7LoEgrTs2ZVYkR2
PzOIrgkh2Q1wPBOgTgnq5VRwRYxUi/C1PfgI7blNGW0JcRpa9Ry5kLi0nGeMORVnKEWCd4sx0aZD
SvHlfaMNAxV8r+UMtJwrAOeoi3S7WFgUuW5iIHild2RCdm8KdRSw/2hmaEbuWF9qPKc6fc1Mm672
TO44LkL7OiaOgcjcKLoxAQox8NtmFDNX6LFvRbp2oqPz7V+ofsS3L0NJ3DhyD2Re3OzP7P13jGEh
WcfhwV8CYsYuyxeUj0I2v0uxobdmUuVMRdopKiIkRYTq6M9wVlSHeMQNv9LBk4mgCSs0whYxgnxZ
xEdViWjFtNowQQmKC9GpcClWdxIM8+ofl3cJAOG9x6MZ8gj4iRNyjy6zaaz1XQAztx62+NIp6E6w
EoQk1FI1kLsjUm6i/nmN6TvPp1T7zzruaGugAh6JGP9wFYfDUKDoVMyCeaoGvnHAyb6DjLZ2zOrd
WjzbVEBu2GfOtrP6OD7S9d2Hh8E8ff6s9dYaqf18pVE4LXQzhWRKRQqhm/PQRqUKZNJZ1Jmqci/C
d9V//aJFiYR37Qeh0rhCB4upq9j8m9Fos0j5og6KilaPNZ9n1FJcYGgTZOLgaAPVaJ4FQ/WtgcJd
Lp4i4qgU/PDszYJDCpNgfHYY8AJEyCkmF59p6VIPAdJUAxwCa/jpUxM5bC4iGFZzaYJoI/qzZrL3
XFyIV2h4/NWX4SKP8dQxe+jFeT05mt+mezcewlGawYS1IBjB1tjXojeSTwiDHOJAAH6XVsWTIrGl
wr5v+65YSICjgAmqbSAz8CWZ2GKBPTSJwinJOqnD8qEYjDsRuJT/oXa6+UAo4T++obwZmvglZ43w
giBMUZGkLEHaJmo7UXHwQmx/mAlQAAkrz0UGEALz4lKvCbI6a8UfWechYJB8wSNyyREBAkQ+d+vU
+ekln2WqbeqwaE/D1rD1ymf7L3vKOCv0GhnysCTyMmZedORLvrTPApC98HYLrP41gGGhY5xs/D40
f0YEjZ7EaD2eF/N27i8HqZxJM9kc0N/xhYDF3UhYISQS5DLOCWNY3usZLH1ZTGkiyaqrY7Iu4mU1
rLf4v48Q/3d4sf3o0r7JQBH1wK9BUjvA0FqNvvtA0KcZLvKlVdMtZ2TDq2QYZupMZdOtKEWsAZWW
gr+6UkWNdwRYHTtj8UIQFzsE5VPkmxX6JQcsO1GG0A4cdiE130A6jSBRV8WQ248Gargla2O9AwOW
JAJFpLM5lZnd1unMsP3z+7vpLgLoXN/qEPeVDorYZWrM8qHdGpdGPaMrbEKStuYUb8OYiU2B/64T
UJW8QrCN5lQlEke/uqUaTRSo7n70FS9gfzTLN8KljqIW8Wl1w+pSKrNUXK4lYTQk/es5uhpuA9U+
NlXa1lQc7R0eCP1wISpUjcdOKSHGmvJfvpjzhQ4SIxTU2JSmr3Btys3fzmzzs0vihErmGMhu2S9T
hcAGFWzYB7rcXATmED7TK2gYfvHlDzlAmrY0ld6Jy2RpRXJt3DpVn5Zb0eol7RNSE81lXpui3m1w
EPMVr9nIpLMgUNd8K3YzOPyvoZwmVXVhx83AjO7VQ3TqUrsLyoZpyEQXfEqE/vd8UEiOwt+YLmay
PwFFQphRKxBOnXmhNceuchSRownR8OQI2qybxLSA8zX+NvKwbGE2IWMuCn0A/vZK0XJ+zhvab32v
q8LWZfxu+caiBcMC0vRE3nlkxdzn4Gy3aqD4DHs4KkdqHkSDPO80InzORya1UpZbNKXmeGBuKzCu
J4rHltMPsxpjgH5nJ7SdtxtzBhJWanqIblvheA1WSk7Q7Wlu0pIwjMLVO9BQUXVO5JrcX8/qvaC7
0RO027OqadVCVwrZZH9BRZ+ZYAw/CftDktj69/8lb8+HZW7FJf0UbinLBJhn9EYMmoiBGSHtBeA+
7nyi3LIw0qKFJjaM9XV12dlnhPO51DbF46oJykcqYdAA+dJvoBZH/EicOeyoY1KqE8bLXQDLQS62
FDqbO9Xg61Urk4Th87ylSN0yvcfIiF526Ss9hhgE2WKU1I+irQkd87GDc5zOMCpP5Ww3J8RxwRgY
c+SkC6UN4Lsjw56L6zNK1x67DAlJ2qck8hOAAzqVIXP3UpBq7fWX1e+EEOfK9d69bJseGWY2AD5m
aPuixg+s3+8eISXEPc4WE/8Zz5B1L94FaEIt860mePA1LeFRpIK/F5+i0g6xd2a4t9ve1i5YdACF
sSE9BkgvVosBHMOMMJHC74zgmwEkARLs1w5hrfISORbWjD7fwTUKXbRQf2y/2mgoqY1MZdeQye6F
8tmACZQCt79L2OtztZwqFUUJqpz3WEUd/hMzcAkSyTstjVffBpJabuBUa3SXMdwnZMJRNwfBfj2n
p1iP/OPrS2HExHRVfruDayp7iaVImDwz/gKQRm0z9DHgp7gmu1A1oW6wh+R1x2vbmJvWcZN+xp22
L+jSwrBx4zvcjfgb7GlwPhpK1IxYfKekkeht7piYsuT1/t+eCXVLR52qWc19hN70fON8VPlmPR7u
fqgJInkS+nbM9+rr2hHPcf6PdPeoKUAv9l8moR0A+c8ZtHpTX4k5NJSw+zjFN3ZxbU2mQ9HtXEMb
62usZP7A7KahGp/uAuB99sKYNo5Y1KUdDiajaaWqWBww2PPOa+NCVgPkPM+nExRThVcGmBRmcVbb
lU0eLNqZfg8McN/PcMR4hFuqkGsNtItp0INha4GPKDwTBqboZBx7j6akqMY4HVpYqu+BgRF9ZJrT
gQT8SMIQVR03VG+w1dpWDbkEsWqSUjk35wjKjjHbyeOpUmKVCT+r+mJOs2qCLmf30mPi8FT0rm5Q
JOBNyqI1lryN5zTvv/p+1tKLEvIe63eOQFvcdPqNf7eyN2zhFZMjMGHZctUlRxYP3et3ofFFliJD
0dh001vzCIYQ9QVKC5gr2XKKxC4EcI8d5N7QZEY41WAVLLmizMgayaHHHJN++WNTFJKhlvqSbcc2
KxKP9qV2vFCrhaVXlYEFfYcnsFWcojJOYri0/+SX4gbnnO+9ffLHEAvonud4FqZefltefKtr0vIn
uAc5e+ZawrrhcLiAw7rTCfkAQIAgZt+CqFvvde+9HpYNsg2n+HG9whl0O4Jn3I+8kF+qm4uw0Xv9
K+msRpDONoVdScBOjGyhugXlTZN9bL2a+SvKXUUkAsqm2E/k5tqDQMQsmdYxDFXAokDryHo1UBDL
v0wLeI5rsgkTqLlH23czHVIC5CUSpgQFq6kqu7RCt/xoG0Ikwzmh+pWN1GHnphYDtbkvHwBAw+q7
JGJLN2W6XnD6hgNjV8YdFpmVW5iBIrWCRur3rWd0+UppFv2gxVrRJbu5pdMoUkUFMjpGyJQfdLF+
Q1Awsb/TuwcE/To6+G7TE+nIZF/nJ2LFmKUtbN4Eure+Cggl+8DF+5r6qLzPvuCzN9IsxMUC4CG3
EtvhjxxSf6V3HPCkIiAh+s3tmSsM83DBHOA8XPv2h6NWDSYUkbyy32w7sEFHUS2L6Jme8MzgMQ0W
KfrtRxcxFuBwrk3rZpwwIgz3QO0NAUnrMMPEzEP8ZkOayBD+Vse/Oh+Gs4c7g9+o3ZnE1ZZtZjwR
d2OlFjgkWA33J3RcuCfTNS+Xg722K7VEELCCPRlXY0z0wrDihhBhIGOqCGgRkmFlm1xUI9CiBmk7
c4yBRbK67CwV29gmLNw94zNtxENci4w8ARUla9kheKmWJucT73HthUi3tIiG0c4hbi6H5bbetpjn
txfDHVkAjq0DkD/icCzTzNTxvJIlDCZQd6bz9sIxF2lZu3RIP7sr4pymAY+KtXgfKTQWFdKK+vgJ
y1dMRz30rlelbBijaQadeqnmTh+J931w5U4SftJKifNwfXoChRtA2enEN7WO5NOdTxD5fvY/uoBd
egeOdRUZpQ7ex0mWTe8kdsdK/QGKPA2lifUnfZtvD7aJKfEEiVPINViIbdExRke9xPkXGQZQ0BZ/
P1czfJJir+BSQbwz3u22l5hO6XgoiwMadAavtgJrdcpN+75zO3DeSNipZa/LME278keLRBRu6+1W
HjPGQYXXmuoeB4pJNUCu2spswj9dL32YQsa6mwIWbAvNSO5PlUi81Yt5hjC8jydBo8fCOQFwbb+g
I7qspkLbDFBHQdC+xgc6zC2h70gHsIPbnqXFOSjuxKpRrxfCCrOZnuEOIujbPNpsqERy65xTjWr5
9nYzjVbZSemIz67Y3vru2kcc+udGkD6XVXEImFE3iNw13exsNtCIENQCNn+MNpBrHoxWDVFzBUGa
NJEl2fye8O0T2Nk0l0BXxwfw/xp3EXf8fQ5fuvHVgziFvXzkFucbPHvUPqpcnQHycrQjpkFYqGui
OTXzOXA7CuZlDKBMkLxDp0lzVmIGprmYY3VO8gG6lHXQW6FzP2KAe5QNwzyLL9Hb+9Q3gjFfhImK
8WJYKuAHi/FwxkdLOq054Dvf82Scs6cVSqMp0bvOJsHTGpy/ay1ka01o3ybV1oXt6FkzjpoY1GVf
lZAOJdcOYjZs95jAbJi3lwTmsszTqD4BbtkLFlMv8TudvztzXp8an7M53Qo4aHXb34mQiM7BWXBR
4qiU96qaDt4eh4f00X0k83+i3YvzH5D9UQOairYT7LGqN4Z2mjLAk0V2cPcMrlvbf+0qLbtHt76z
cuUmoN3vwk7Zxj+I96/u5UNS2VgyjC4MlxltCDmgm4Hn3mbq+efiFc8qeUnHrq36azVszHW3nJVx
SmBSUYcUbzQ0WnZb5iK8/sKsJ4WpPZhAaC7EIorsil314Xv8fUDHTlajER/Y+DsoqgvMX5i21EKN
Fapg9/Fls0w/6tx9XdbZFKBvS2vJzWw7+kFgZ/6tIG2G1Q1/0N+gOJ7EtFyh6wL3gS8DbvuchxlK
TV9QX6prg5khDKIJ/bppXOKu/CE1r4SbGFvgCZ9iePqBNAYyPysoQDnjnQtc4n9k/lM4jsH561S1
As86qUccoNkma+QzaNwYbo0bxIIRN/C2m/KmaiVcFN1WTwCB8lQVq7DyOH1QJpIFIH0HUqOLgYpd
otnUKxJszbzJCMgyCGDAuug7FJAjWboqpu4TS4amClhHJ0jFKjqSdEmB8rBa6w0qE0d6gUOWgm+a
GwCFh594uKO7Cgs2haOZEkkywGxb/uJ3Gd4DqusK4e4iDMp23hcrhCofZvEMlQxidFztSPeVPvCN
6QJNwnbqnv8YxJq05IRUSzk3m5TJbeVDBNum0WBmOjmYeAy2EpyyqKHWOp5ogJpzCljaBjRSwAQ5
dcqJb7AbiSJZqYmly++AdgL8JVCqjZVIXRAlSfYvXn6EvD3P53m4PcYlLRmhAL8zJWByZayMBzhH
GweJwsoBwlNtnZRulbXNG2fd/u76Ey64UM101ijd4/whKH2TmSBIElvRAFLrQXh1LuSnbUAkxcfh
MYAt6aS7ddK0dBY0k8T9lZQRZ1KWoFa47OsMHj6R6J/aD96k5LSc58YquxpUoOOd7zYx0Te4cvLn
HM0tVYXfjVVnXUCZC+iLRwJL1wFHfF58VjXlSLs+m/CbC8rl8ZWvjgtcwRWWXPxDTHD7oNC7wPZv
kr8ZLBLcxWCtc6pBT9InsU17ok4bvUG+nXffTGoGdvqQ9nhzewJgOzAzR7C8AH4c5efwBHXD/lFH
IwZpfLtWXZ7f/1K3Wudxc4z+LA2q/eRvZixI8Reb6sSUiFTjsp4fx9tn856TUQkyJzIu2HzqtY6s
h/tJm/JNHbAi04AuKoNlnxvHUhAPX/8almpS1B2LIIKrHFtlXXq0VVC7KQ9ezh84vArQvwrryTlq
V8QSp3gQrswRUVNc97LW0VfzHyeGC7p+/gVBtnAhYQ2n9RMxKD7RozDbbu0Srcf+GtbzfK8X8J5z
FRmOLx2Zb6JNvfVxx2Bmj8jqEgn6hKTZCEAQJuT0Iqmvh1Pu0BJaUF63qIYbE497VXD6/SkVbVx0
e14Oy9Bxmn/y4pham/e/NSSGQ/2fvy/KwHOSiiwBR/qp46+hvdPW8uSg8FWK9mQ05vqIwso6NaVZ
oYa0FL09mY+8Q1ZZfenldsEHLZPhRid6GpQjCN9c5HztBXUTJEnHcBK5rlWVpb3Ye8CZ7rIW4PYP
t6O2aALMWcSaq+v48M9fcyg/IsLgW9QTs3uFOwTaM5LAkXRBgGfGxAzzKYMNd3yoTADJ3vYdG90O
eDejzK1z5RJdhmKyimDBLpYY6qsOJexDvRHQFVDsEGeTtDBScdDBAS7TAcplQYChwi27lKj6/GyX
AT1+zNJngCEYx6qwbe1bD5zaRejlegeK/MEzn6qbrEwouNRtfYzqRWiWkrjw53Wnvz0Qkkfo1Atl
XMExT3VhLP/vPHSW9YvFsJzOI0Bd+jtEujYBzpidGFdayOfsQTwbtZ/h+69clnNycPnKFfZ/nyHx
H8jqy3935+3eGq4sWPlIIi3gfVJLrORFdghTmUpxVpu74Q8NEMCOkwHBfmEVxR5oW5cC6TXMoYtr
bfFVogVEzLJMU9WMM9O7bhtrTsjsCJ/ORRjekKS4jZtmW4ZkFJM4J4QxMkhsT/dOR1Xxle92ZpfT
aACgpics1onLYN7VofOfO0CLWnLcTKGUHFTvI8SRVxrASJwYii3EArp0Jq5jw8YokHFmSiSKSesO
wCdmapbtVaHnpIoHYnOb9JXUbgBCGk+vbuIH9qjLCGuphYzWI3BGQatGSkVQ36p9RPYgSnRABs4Y
5V7S7VtC+Rez3ODVU1ABrILsLs7RtCKvsJETgmsYIZ4trlWZnAWaaXxe7EsMsnQD2VvlBNWfNEck
BtCqfYGu49MVXaD4SYduFAJCqoOIqgHGJGaPTmzjDHvzxsOFenxqLy7uTe4JDKHu06eyLmPIeETo
IeMZy1X+wlO+hTEKuPsIQAy2U0NZ9ekHUjRckg44uPbAcYKeWVjzzK7muRrj2rilc4i8eYDOrt5N
Uiq9If+or5o4z0iPEfoKkF5ET8CxGw0EC6V+U1Y52oS37EhlQtllw9LcuZa1n7wekn6MdhCta4Ue
euv2ZLE2mkitnJo8VGGwJRYg10Ld9qOjra3QbWWq4dfXTLPRGAPAehLe3ctWPAjbv/65iOuG2fT9
Kz9jewnoJdVNMa1W40J5ic9dyKK00IAUIb0uqEW63VReqlEHZm4EucIGRHDpW7g98R3Zzc7uRcZX
d/3Bl6mSr/a7/43mkLPHhAgCk9AGFuVmbKdSPnmbE2wtidkOZiCzAGZlaQTvP4FI1boF4VHrHsCz
hOD6EnwWnRCR0fx0maMGkNFN7lYfxWHNu7Sp+U9nptDUcsDAu/QDC9c9ag+GKkaYQcKXVHrDJLnW
lMs8pOTy32EYMIBVjZoNloA6lYx5lJxxguzFofRzgLCnwp5fd64JQCqcKPgL9LdSPRYlLt9ED16D
ADS3K5pWjyHDj7wUcQ/ijUoMlHapkOfnnFsJN3YhHBJiJJrmqZYJA/EGQ1VHBdKQND+jbTc3Etki
27OZBUsd+kK1b4bmp2WEEJVQE3xrmdZcLZhR137oYflyRVZiI24ecmeAUNngmRQUBNTg8oLS4zbH
BKeBUrMNyGb97Z3k+jJonvMztuotrZzVyFRlz+IeqsoJrCF41IA9nwEeQn6HpD2hZsB2Viut0Hqf
Chh8jRPXpBwqvrXKWAlyR5zeiJ6yLCfYx/U7yAHTVWbkaZRIVffzUfca/fd9N0kzefrK2E3gzckA
AaJ3UBsn0INJfRzFplJMdxEIBYqeItupdC05p8NlZ0CIg+VsutZGLqpMvPIqlG5r2/y6x1QwxM4Z
H6S8fxLygqYzqMjF2+0qxF9TLE0v2YVhGU5TjWXooYu/vU/Dj2mUzE9LeiXT/AOaGf3XEoM2Ik8G
fAWfSKrQ3J65RNSPS+4mvuhg2qJ1ESQcTonI99QXonX6tIJtOajjRwXVNLu5J+mXzp7Ai4YrxKoV
efszLZwPdgdEFcLlgjfuhiKwMGPsY6bVsgFEksOeZZ4Z5ilHUmmOgG4vbRBYJ0gNMamIypJ388IL
qAPnCEsZD67J7DOpp3tV8Iw0pg1kEbabM+BIhq7uxRL++svhIhbI5l94BGSlCecJlMIllohRo9OP
/DB9GXsmkRv6ZLtfDDozD8JEobFjD71DjIgMFvLiHkv0RQn0hxsQzQiJPMDQTtaAUBVmskrcnaOh
ky7N1u1a8CV2lMNZK2p8sERVBUKWSdpdnRkfs1BhKC77duSv8R9Y/trAwDEEf9J03YlQdNeEIq8M
Bn3QKcz8FHczudceL2OWixW/z7uUWUSMOtGDqVTREt2a1SX5ekoxzKcyjiBpu9YkCblWc8Q0g2mE
7k+tqmtx/TVFuXJM1uUu94f96B2zr7uterGvx4jVrUWqA8CXigt8A2mt5P2VlbOhVmSFvapH1HKb
hkkZvJKGpIPLz6zcQpYnyXQC3m4yMZGrPzYmBdzTO0SojDUyFR9G9TtAb+To4Y1zsa/pZdi04MWp
pkMf9JDZEPf6SxPbiGgre5Gh9Hd0U/wDShN9RdFc/dNcyin0Ccezum8We2/WDbNvCQJg1I/shrJg
lHO7S3FRdQTyy55xmRbZVzdG7QfZCF12EGRw1n6ySbB5ZVOTlZkLDzZ14zIpfQeBsVhkz84+y89j
TaNENUD75OeDTgQtSDYzB/iAh+kNCdAbuqezjBBwaJFOUj84I20xid+30Bc6Grpd+80u3jXIa+73
cV+v8CYy6SDS++zyk6YVY4rZPrU6vr//LyUz9OxQ/MON6v9F4PHn3XB0TVoSaPx8Ngk2/pXy3Lnt
XgmtQv3s+gK9AUPUcQNg6r8pE5i8y34yjCYaA2Wock0v4dXfg52f/TWCFm6jk9CdOwR9ZVjVRCh1
hcRbsyTkyaJSKbC6xJYSYrKIrkS14kaFOYUAKUzzR/iSJXsIGKc08Ov00piYot1NUZJmawsB9LKL
+UY5o2poDLeYb3eyPF9FAU1B4Kro9t8WeZu1Qy2AIpvr9MBRctnVYkzCR6rlc9q/3dUO36Xl7Ce/
PDUeYhZzTUNZxtZR9uMdL67reHmJymV0meVxk9ZtWRegw9lQYIFx+g5HpCMYaceDPckJoc22Xbl1
YHvNFtPCN34qNP93G5acDwtZfpldbz3ndeeWWcvrSX7KDwy/YKfmtDYflVbBeQny7CmIfYwY42Qi
Z3I7H0yOGCmuGfqVBEIX9rAGmWd561EdypJEfwtntmwXu1OwYpdaWkubP2kDYd4tLwHOFStRdTcl
rJm2jCGLnRxVZFk/09oFYarGkv9sMksu1u7rj7J6X7I08nP8B152Zs/jhzaXi+87tHzKYMmAk9Y5
6nGW6xJ0Jmigz6nTGUci4Hhn13Fmy8jjEHgwX/Lk6AO4RJlI4OwMUT3LI2tUsUvfnfOxc36vs3EC
kw+kuJ70xuPrlI4dTDdat/3Od4RZ4ZHVdFgf8RAtb3Gm9Lmgk5g2xLeNydwgDN3yXxWbbzq6pxyB
GT0TgIpty76KYiIIXzgScdpL1zIZrAiNsJB5obwFjejlpN+9jqdevSw1lZ+4g/CpMBsy2EA/J+fb
hejCOt2Lb9sLyCtOeAU3TixHzDk2SCxarzzPQe6IH82Qa8vPb6Mk411sfbUAzXPWIhbWB45donsn
K0KLCAX0/8lXnYsP1gseKtu5pTjJr/XDwzR5p8RBko3PlOoRUQpa0J+v4FQe82Clc/Au/xhlDQ==
`protect end_protected
