`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Fsk2N3yblgt6EjzdCMbheQEQtREVLQqI0MW9WD6epGtOmCKKXJbakU5Y00HuI3p+SD3lura2U/LO
hYvbQ8opYGY7M4W3cWhUPGXnZ0i6yaf08nWCoLbMnw46gpriKL04PQOVFQ0YYEdsl2vW7lBrSaWO
fk0Aq6ZKkxs0W332I6qW0EXXcOp4lELq7VYuayZGQcURwHw62D01WZacGoCWxfJo/eST42YrQokQ
jjqEqRLfQWn751Flw0MgY95fGWp+tEPV1DSl61rTJwbQ/WfvqJDlX4MgDSxYTzNRcIOnRLGqM005
hQVvy4yDpCUfXA860nYQjcXRg25iwK8X9K1VUg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="v2uWQxz6p4fQzVn4xU5XucjO6dwik9hl4LTQwCEOS+8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 672)
`protect data_block
Mfi0mQ8CCc4hcwql4Y10+KWVcy/uvzxFWR5Qe58WR23CwcO1jXxwPfu5OMFTmnJcPuu5w1pEjudc
udOJzBtIrGR6eQDe/R4eCOT4TI6Uew1Bm3Z8L5dik5SffgTVxrn8HEDGUQVGsu6/8R8qnv4S59rX
Ng9yQCRCU3PwrZro5EWiUnPAeWl6WBPaMFZv1guJ1A1uxJrJz0rcg7LMdT2/qn1+rZZwO9CcBSym
/qWtfQyDCJINRsQExVlGY01eA54zKo2fVuhZLtKG9jZpiJNzzGOHs82H0cTwLea8beMWa2sZN2Sz
JNMk/LOnTeSyNYkSnlWbT+O78vcI7phwebjjtHuCDYdsFb3GGT+jLbcCrDUZj1OkXBECaA5X3Q0n
A4hPBc46Bkg2Ad0GdF49dGZp0X5AU3mbZCcPbdsEzUTjGpX4uUK/33I1om+XK7uZ04OFyem6a7SQ
mT2z/aoZQkgFyCDw3iBkYlBjT22G/ftOhrFdDlexzlJjqCP3e1Iwql6902l2rjnE/d6kOJdSxW3W
0QjQHYBp2wpGJ+/H6doI3vh4BUmakW1tmGh1RtIfHi5JR88r71OCa6JfV3Dj/F9cAalClPgDr+Bq
mNZiTL//0btyLhz5vTsq4RU1lQrrNXAj3yA/ND/I7mqZQeqWzkwp+qwiUGbZ/hkWz5f7oeSGFgGr
lHEwtLaxR4NZCbfWuv2GgfWtm3UN0hB2bjA9kGK0hSIyrJ0x9o5+TMI+0EjYSCXzJ3DZNenjfgo4
/gX8XnYkUHcaBHG8gwjFKJGOMhaUGa1WjbfkkUkMGgnbVGSfuUNveSbvJj/dWfdIeHIV5eyXAL0k
eH4bpLbumOE/9D1uWvYC9aZimPwHbgPsxKMnSeTCRs8sKkpmSxXPZI5a5+1q
`protect end_protected
