`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
t0ImIqVFctOEs8b+dLfnbRaVBwlJpQdHPXfO7wqypbLG4naZsd4Ums5ua8Y+SE/RhWXRZ4C3L4LO
Q242Oyd2PknREKyDZqvh3jGdBclcwV0gG6Qdn7by1Geet5tQYqdQthM9qA2YiUDX56Ad3Ia0Bsad
VB8mOVIBqE2Q3nWismiTurvN/rGf3JZQTcMuNOUL+5zZyWgTIXceCurxdSGOeHRnWGEnjsIvDuin
DBIC+5XYntIPEE0k/YeDR3vinrTlbGFNLbmTNhLGmLnhhPaScD/btomRtSZAUs8Nj9fjGD9J5Vs5
W/slOVzK55pxUwLvf6OcDr/UeXWOyiiVtTlIMw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="G7eJrZlKNbqClC1HXsMF5c4SSPZB/RjTB1HjzONK9wc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8624)
`protect data_block
dfQBrT+5jYNc8y3fCHCtZJKKvXdzpmjiFilWD4sUDViPsryhd0qkK/OL7RgbRP3FjfNs3NU2eHnN
0bViouoShjjwnJbDKzti9jQraJRcOEmc/WY+YVrHA527QC4NAKHaQigNJeP9+1FkYdm0h9nyxdB4
NHPN/S4IwNS3AFm4wZCC5d6EV5FcAM1tw5vjHVQ6PNNcb7sTFMQgL/qWxZOF6QKaKgy4WHvsGzLV
Iu3b7Yqt2XwQqhKMyocEyrhdBVGMUcWAN8dMpgILYXDSXyhigT+SCABosfdaudv93TF/O0efe2gC
D/0rWRdWuiSAwOEQgcknnCelRNIK+TZPXneUNsDbmtHFzdgKnmlEqvzQO930V4MT9R0cemfZfUPs
isyk7ve/tVpY8/nSQ6YsdGD/mKkeZTb2F42mrR5PDN+QB6gGJPb3NnevT3QkOZvOWdZTSFWXU+KN
ECnLkAYMT+nX/DyXTYWcIFGdPfMk/DgzB3jQX6Bz6yJ9sNgZIRUeU2ZyXORzfPxHYoMjR2LjrxAM
VuSF8/3+PbfRKfgncnTYwHCkWiKzjNXBTTmaIRAUEXvLTC4oVciMmT9V6iKWlMVrvG951dstWlCP
EhUL9AYRACtCEYL9VSBtJ3swZZ+DNhnphkn0uOZTelF1hsGtH+WsVdN7ncTrDWj34F5wsjOigzLq
1aIwpXX/z9LOZBcPTEhotTCoLOCFOd0xV+Tcoy6qoRIjvCjAjV2UUYDYo9U1oFxwXyhmGERsQJRl
zKjcsLuNMBME0X4M9eT5tCHapXfLP1fuvb/rMZEaCIaAj3m3SxcqDMHl/NKvqc2bkrfe4P1ipHhl
SrsqJ2pkiT3ADR63R+ZlwiLYXixLM92kpqAywTLmazesNQ/HTAs5OQjfRthffQt2J5b/eyD7W06L
6svKbHH4qhb9kS3x+54OqyJBvU+ZTQIkzgAXC6G5qPhbFVSAJzZPs4caYu+I8h56db75AN4k2TMz
h75jWSlVf83R33eoqFgDhLZ/p+EuKQsstkypK7A9oSv4ZDBkraPEJCKMO1KrKi79P3hDkI+Ho+Hs
UE5KaQXFCoQlBzCiQwWWP34tyFldyu/fBYKIkNTQFb1IFc2zXFDOOVQYvR4iyns50Mx9jCK7tDVf
cAukoR30OHB8yLRsu8SZqEtW6AENt6pc1qhI9KTHsDA4+egd88KL4/Rn8ZezaxlyWryBf+xXZICZ
78xCUe+9R4xA1X7hMJDqyJNnzriarR6FyjkA38X9JJX7JoFMttPesMUKmQYlyzHi9QpD5vB0frWY
4UrhlIgEXk7GuuvL1KfSM7BVSJHBm2OGL3dknYMh5mLRZsl2c8l3wg0UZvLT+ahuSGsb9pYVhkzR
+VAvaNwln17MjY7Eu3VQ3tDNRmJrCH/qasldzF+L/2qUF2i7g9UoDE/Xi7niF6ThJ27ImkUYomcP
+HPh/jIVDa5nXTy34xeK0Cn6cNK2XPjHq9vRNMgQLJeHFGEcxvtIOMQRJmRIxKmF49VvOt16uo/E
aM8diIaQxq6VdVvaglj1I08/RBaQutyB8QgdeomkzRqzfcie2SmfIRHYryQzcUKWmTMQulLFrhZj
zVHdk6doi3L4LFp/2hYoCCTvA+g+TgX0Sqf60iqHKy8NH6cQ6AeHhttzyVvVomQOdz3Sxv4lZrbc
0319AgtStJDcvm0Si/R6pYO3gBq23sllB3bPyjgRDcLyPb3Uv0QszAQsplR6tu+Z0KiF4UrYQm9b
pmSXn22xyYxzQwvsLiNqK40A7dA8jXEggnJmSj2QtmsYGcECcpHN5VesaPAaURJaH0i7rBpqVFkx
g8mUcIeC71PwZOP1/l2D/Zzt97f40/ycrAtfcFiz7p81SfKcCPhl+AHdorb3M5e5HKQqE68A95hW
lBHlAkQGYyiEAKBvaWLkcxJASTDrTdD/ZmjAE23j7bbb6fpytmgPP2RmGU3NmpT/GAbBEsCUbbcq
QLDfSKXkx5xSAsqkuSG/TyzBjLv2SWylvWKNRUZFYut9NVg7S2bRK2+dTJ3dcZhPPsRuAq3U1qHi
PVJ8bBCSZPiMVJkbI5rM3yQcaUYAwEJ6Q8yQfeyaW/MJP677SGBQqR7OHZnKXO0MGKzRRvQjZMFK
abXwfS0U6k2Iks/pv+1IeHsQpNVEKUKsMa1ssa2Nc/wWvfEyJ42WwGfBq5V+LGslSgPtk8Dlf8mf
9BQJOdyKKllydu9+PMpLQyosUOztcKyemB5yDripy4sbUZyMw/V6hR6N8LS/V8dZpzrfeLayNyc4
ozfpNaRPO/ktdccuufHSdlkQLhBOAHYokUGAi0AI59VPY3zvVYRhO2mzHXe4bFOluMhJduHHJD58
7+8ZMtEGAlNn0WqBnAG7yGeBYa9qY217vxSrMmF1JISU+D5W0SmM5h8NVgbjwM0IrR79nGPRc9qn
dvhezI+cNz0r6kRmjQkSSB1VSlqKhb2VueefCHhXiKNFrThw3ySI/kinytQs8C627Jo6oidWFvM4
O/amDMzaiiL+31Rgi7oml4NUl+dFwUi0glvMOO0gu2zUgOZJfQve8hwRhirGVXxHP2HWgPsBUQli
fQpIuLhCzH/yDliQ2T4iciopDINCGOdiMlYuxF+SQvmONXVOTytJTD2S3mCaKK+xx5v0PrF/c1Sh
RKwqXDXCn4LZNXzwNdxILx791OvvZBrRYWsKwlxUk+eZvRpcuKaxZaQfNWO+Z5BK1qxTtQUYFj8L
4l0C0IGuQWTefRNU73jfsoELX2Qxl3TV22CpTpYYyWPdItbjmRnXi7kT5kGroIUt/CspwRRdqn/S
0nP4NRwpPX2Cb8BRs8BR4/1lyhigbqpHv9vXbl9jywAhMrjoEjebLtQIrCibtsFTZEWke0YfiD+z
mjyhQnWWrvwPyzzpaKIpBvQzK5rtvEhN0FZ3HZ5yDJKpL+jixMsy9AK2lcxtu2hYoe2DvZpsBXWV
WN6I5dBFi8RcJmSCQ/+IL7iblj9l6dKymmat0c0Ctl2wsmb1WMYYTVdZEHSPUob6+Q+sDefQDqfP
EeobBVYvgO1XQHV6BWlnXM6wZayrBqUEp//tN/OlpEXjjzPjQvFepl03gDwih0zMLYPrE9VuXHPZ
O8pNrZHHryXNJNr/mrN9nu3oAxtq5+qnV2GGIiZ89XCDlg7njI1gTO9k8Brl9ifzsDz1+0Q5WMaT
WSCytMdG/dtJIgJBomIGUWlsMbm2kUlfVpvhXG2K/2QJiY0es7u6qlJbioMnUpSxTCr530kT4IIh
JGJKq9ze4W6Qa7V56ZMko9DTBzFKY2ev7BQ+RJhTxkA9yITXDGEBScySDcJ+0p78Kv0JViKn4lzT
fb/Xk4yLmC2Wqa4deG24pziuCgX2wTsrumfIevjv+rjU4cUqqBF435RkzW0yvTMYqVu47er5wbhL
KtJqwuDDhA1aMhsCRSyMhamoRc7s6MoZ3Ibu0A5KB075dxBo9etSqG5dDbI0Gqk9rwPoWRLdX/VJ
/P9jHv+dDpkJxq/1hKZBTMIZnJ2uh0t0DhQgK2Atcagh0N5R4vEOLMC483/I2z7/ULOZeQtQh0Jg
5jZx+s3CV0COPgZme00yVIU9IVzT8pDMHjTlB/U8Z2434HOUbROQR5JRwMMD5oxbv1+xUKKRWLAd
25l6UWxp22czDk350cUXYxyt3LCFi0/yeJay7lOW3mHMVw81RAgf6owxf47B6uU3cTGClnJUn76x
0cqHPXJeIYCNbL9XpgkPakduSGxngRwZShn8hn6+2l4FgV+20gLIbMGS6px+YVI3fNkZjnbWbbhh
TIdg8vMGAPi6VSNVKd9ugX7QEmExygYhp20ELLJTxvlFXA0ClxG9ZzZoYZ4FgMosnvDSxMRbm7Jp
JSK90jUNsPHfmQrTS6+wYvB/tbkfS2FEyWhyzzQGtfYhjBnwdtjHvbAWlg2GrM+9WPS/bPWl63NC
hpeXh/05rhiUP5C8kjcOcm803UCGsxMRX3uCb2xt6OlcOnPTFMkZ37ydagWiHkaoqY9NUDkNzaQV
PkP/mtSaRXtbZ9krO3UffXzhTvKO0KJRuopVTlzqkrBBnHBRM7At643nXdaLrbUFd6U5Hf8aVGO9
1HcsUn108jpWDzsjGOtxyGDwNZhcralRjde+MbJayA+gT9ZVJJcFzVVcRQ54jK6qeDtvaYyjHEKR
ZuHu3DlOebjGsPaVs7fzwfDBy0OLhSllT5LDmCTJ4dNxTZJl6js6MhMIdhcNw/0BN2DLqHr7z0rM
tNvefym8rGEz3kqvUl6/YB9UN9VKE9lWbXUk/6j9qbpwwjSfOS/uUk4gHzDVpbHk2/hrK5ztQuNn
jTRkJlZU+BzjIBCbnMKTrB2G3dE3F/iOoso7jatXjlKZvGiea6IlTLcJ8fy3aJp5tXn95U6UcO2t
BFQTmnYuENn6jnsqjWX2BJFngelxfAMmED7CrvwuuqTEh39InJKktyu6YmRPZoro0dkhzy+EEHnQ
EXVeKMLZZalI2ezuFxx9vCLdK/BXHzfaiz5KveQK65kIKM9szEWcoYy1TaxQCZAPMzixLDIpo2N/
C5L9RKNGyJjzb8VKaBo/cYxvz5ppWxdblTwsiBYtGGU/dPYUoaAVfTasS7Va+xbfHyo25i8Xgl2s
Ljt9vioTjyscU87+00Zxi4XLmdxvJDTModzlLqjrUQBIXs8RKlOTAStUIPEdWE0uzWbRVZbU1HOU
Rui9l//ht+sUtdidGSDgiXORQCf7QiOGezUWZkxdUPDy0upmTkDhVQnYbc2Y+flhuGXljuJ+Ka5F
J/VGnGyo4dEVkgdNHi08SuvVSy9OUqEw/NTCz5LQGy165zjnPkmJTx36Kjzvk43D963IF3O7pMtA
nqwyqEHU9fwpl3/eG7r6E7C6EI4GhQUoWMfWJnZf0IQXzIQ3ZhE4dAAC6XEpYwvk0yV2g4P/W5Sb
fqyhp5nKzecJT7wz188BD8Y8a0OwE1gQxcWa329epCET+D+c1w1bnxqkFjXl/aAYalSAs7o4piUK
NckZwsOsbjoXonjV1h+OIgEYCMAXbVH0Eo93gHmgAKlo3Xntn/uqI6QeJBgrrFK1I1niPfVRqgf7
4JCQ3kilASJhcYhry4hN4HhLdBsTIyyAaTnPEcFDnCyMaa55GM1GUlV6de7CFb+pEnNgJ/hfHjDF
TiE8qUUPRpG7hzlf2Bekr2LwDk8GQyjxbuO00c1I3VGmII9m+G8JwTsxgJK9ckAf6SO9WBv+zX9F
piB+mSyystW18o9trkIz9niRgB7+hYMod5Gvq+uyHWaPKvOP74uazSZtJRtJXo8IMUhxz5ES0Fxf
rtNSLrh7ueyS2Cam00n6rKH4Y/xOYIcpLTE2wK5BZQu16yTYFOHdoZslYHDnyJjLDJhD6jO5jH37
NN9fYDFl26JZ4CviDadzhWIGb5rq+LiJ3vsT0mSIaUDIES8xyiZxMTRQ66LO8etTcRiF3FJZme1x
3JsZVNmkNeGO08IJrUWqT7WGdIGZnr2oWds+FfYhxW5AuumVIr1+rrdHeEQer1P28ZQLi2GKT/UC
9wx2MjgV7pgyONy3ilo0jditsN1t0UPmf6Mmh5fPaxUMiQL/koaAwl744LswLE5l8K0G8XwYj2ja
Q4MNeOXsKKCLg1WmXhbjFjylzCOc4qPDcdBdGAUy8tMrM/0py29emKHl226bYa4zDqBGASc9AW4d
NeKVokCTXD8b61/lU2eh/uBwjMPj8LksJvmE70PpomxwyjCk6HmGwU2mOxB7OtCOZ0yDUN0nvfl/
vyNW77QWMHgxg83fLLCGvesWDZMGHskLtc3esbLLD1D8TVEMvo4nNzocw+92jXpH5A29pivxf4Un
R4bKCoxejYdoXX1+e6CkcRPoVGqG0iWriJAO9qYlCc1MEKHwj0IkGuzsD+7O48sicEjWD64QFFa5
oFioFkoRRGpxDTaqQMlvihaqwZAdUjgeh/HKpVp4i/c5ELNfQDrJ/HKphNbc7YavX8Ub06Ysba4Q
Z7yEzPpDqoVtw0nJO3JAw22+TOMJlCftWoAnx2pGCOCmuioCgkfQSNwub0V/fMxfet03q9PSiC3n
fxT96w8MgtGoTsF+NHRLF50Jif9g9p18FaZp+6xqRJTESACLpEkk0YIsSayl+jw/SXZiU/DaFS3i
l8XTzp3Fo7Kcdtn9dYs5xJOv+eqd07xCUhE982Y+iq/S7LEYKA1PWeMcgas5JsMRe8GsQ9hN8efu
KPFFgeBAvnLqZrexhiPYpZp/RIx0ekt6ge0NKuxWpmT2YGsAPwBMXvvUcO4A2lk3TojOlNTqPfMH
o++XTP0+bmLOaHconH8ESPDAf0Fkd0FVQnlVGZjvqjQVAefdvoYJ5sNugtYI66ct/JYcjls1zqQc
XIwQRLs8ZAcDj+L4DF+NV0vANbtGoaxJQQM+W9vNAvCfw/KiIvK9t978vjQwWhLMH68Gl0thMMHe
Wxn8k4elAvg5wP0APYPxsj3eqPCIJKmvsrGmCwJ2s4zavQU7m1eVVXShhOEAKvKU9141xWd/fCDF
bvUQLX+GwClP+sEvkC+8LMjM9DJ3JbavY7bAmLi3dWrd+jnI3HIMofZkwwVsHk62Z55s/YDQTOzO
9mSi9ayh9z87Vx2SeMFEyuj/jRh3JiuBN4jGUy0uCCHo0NACZfcaTBqv34tsFHPAjuzhUdV4k92m
xdd+j7zqS56Lv5eLzRuUFWWd8Z3n+/sP5k7s0ZQdv0Qj8fuxzWU9WHjwCSVbocvkvokyXigP4KyY
8ByntV+ueLM14paSNedQfX0sak58T0iPSbdCX6a2qm+CYY9NsnzPo4vpTlv243ejkXrSDGCjMJVs
3BTFfxKtXWoWVcGiPnmulcuuETOGFzVZ2Q676i6LSe1P69giM0TwVdmPgQHAsMHFP8GeHt9d9gM+
4/6/Q3K640rWlCaa40KFLbMPyUwTnMEnFlJXxOq1l9HpHTceJ/fr7w0eyP1r25+gYka1UCs5EZ3W
M4WmPBCJ2LmQ5us9DQkq8nNcPtZ/cPD0iwaj9GINBflIE3RxqqlYR418i1S2EpUTZ0icgqrXBXUE
2aXtIQiVWkHNu53IBZV1GA7j14UwGfc7o094bmJLTa+ph6JBdc/mMeda33K93JeaRcuLJ3CMS6XR
bS/tpsjQ/BnZDUKYeSg5/O7s7YgXMxIu7jGuMbYYub02gVnGM6OUFdPNLeftK3xj8M6ttyXPjRau
r2XIOQlZc3bfXlfSdl6l0qh/Caw2T08m0Rc80ckPxYaoM+Z3Og7mGpORTR3PvxZ9wI/r9i0gvQ4u
qV8cZIRZY9tm33hklPzXAvZgMywCwAMtc6PNUSn0wQ41VvLIFmZRSmpaNxT86ebA599DQMgv4fqG
tbI9sZATGDNyJQp7LkSaucuokcGY2tpcPtNT0joV6wOtaTYxgtGcqGx5wJT6MGHynNGZ838TgfVg
XGDQgH7KQhGNpoKG6vpBLfNw6jGl6GtgXRIOHhVl11+vRkPllpgR5Bi2s12TjJDT0KkzUKmglVQq
vrZhYOeJCyppRqQ21yxM6ewCJNRnX1M3oTx2LYHkkm2/FMtX7b55/isrngogVpEx5Yxfw70e2JyH
cKdtpu+qMCv0twndmIrLhmI9FRV1A4jgb0sHj8uprNhttAzaBSQ8UytYd+Md4JocxOU8zHyJEeFI
rA4knPt5mhG0PoDKD2hhV6jrN/LaRvdF0gy/rVyLEghvZFmm5tU5k5VakY4YV3y88caoug+gcTK9
leMrWF8uhR+2TxsgLwKV7oyWe4Uv4tXu+0qLGdetJEDCOrQkgy32vrjb/u2V8lf92HWfodxSDKVg
wY5AVb/0TbTUoXB2d20AYkOLrgbaCzjiGOf94cciL4FTG1DS3tdZOmGLxuRWmPqrWZCbaKlHVWqb
cY6YePCMGt6Mvm81cLE2z6FlwNmMuGHa9ONse5weHDd7AMnh624/JBjOwwx7UlukIKsl+BMsx8+E
R6pjeldSgJ6baWG05wx0Aek9BjLRWeQ4o2ETCfqGDNBbi97IBtCIgycEW4TTK1zyMJgYYvt5lfp1
M+Q29dKsEGHpHEn+UUzK4Z4aNdiPULB+gvZsvtHG0yp6ftk2fLB4W/yKeFEs4zPlDyM7zEe2eOU5
Vstol8ZLoD1FBVGznbOS/pa2WagMQrSXwLguiKzh3yfqkmggjDYb4DMGJ/B5pUvuSfdeJZYRq80P
zgX5iui4vbaKPsi2gVFRrOzf+kU7iA5I4c/1GIvhH0rCDugSE9q4TGuMxm+T/Wir/pmPbUhepBzl
NNUrhIQvRtmMSfP43zOPyHTJQqTwSE2X2foGGiudVc4/IT9U34pnxDVpWRuXI3RBuW4Ny1kYn+Ta
b2nFhi0tVWHaLfkVzFL2KZ8A8hthKEk/3MfNr8cgWM9wBhkAXwRgQeAAOFRYfH7kmzIV5LvVyt8G
vgeC7baSmW/43qNsiVvaIl3ZemTv0cBCXTcjri+d1zQP8EJEKsQLiN5LfyqWMr3YhL13KvCtMcnl
lH3hLM4G3QLZJ3keo9106lkIVKbpxBA/2qsJ8dnWDLBErqt87OMSL7eUhWZMtNyIGCOJg4Tsrwo+
BQhRmPl1UF0bjPkNyBxJrP7nTFBM0qsmS6X5wuNg/yOcxOqTt7JFykPJKrfyuelMZViNdZfoE8HP
Zekg0r8a2Eve/TobJ1MV0gJOVkmRu1SZa39Pn2JkUC9ogxmc0H2OhPlViShBxutRByOKO2xo/lU7
ZgUtKhTws7soAvgrWcpv7OGO7s0IxzPZu+rlVDI/AD48H/+seFuw9bIdhdCAMaxHkEOT6CP63JIP
z+IZ5UI0PKC17ZGlXMdSWGQluQtRFk4y2Dx5GwZsEqE5eqBIOaS2aBacdeIAZAAuzbhFiyNAtzt9
qhuxf6lncoTBJUT2TJmnTuA8yGDCofPJC8+XCxeI8bdTq3GxkrUVITHkCvymf19FnKFVIxIRwas4
SYROEY+XeV6iC+KAaAWm86gdX6bz2lDcTpF2ZxgJEkBq/1OItp53fzhgfCjDVW0LedcSL9VABCvU
cWWm4Hs4sQSV7f8FzUNDOHBMP8+i3QeX5Ja3snoWXTiaVIzjH1VdyyDt55r9WssAO1zQ4pOowGXQ
vOROetkQ7c93mPTS/zuD6odqyWDYDwURJvI2sXDv22GuORVW5biPaBhy6MsQKhMVIZnv7KvpiTip
sAZl6WpPy+Bu75l8KrTfhxPtNvYn6O4FyPS10NtLqpTzdV5XtRGvO38sYZUeO45t9a2w2kkY0Ly3
7iK1C2HQxO730K/Q1V5evhsbivus+yEoQfNIchGnB8K6vqb2d6c0yIpJl+sqwBNcqvJwExabzL2K
K9778SSDt4AVdfBqQwJHhEYT/BhH4BB+A67L7zBIVeTPZUty6tTa9bLUK5LH2A3lc1Qm6Kbrhm1z
vKIH8lkybGetJvNa3OgF90fHzgOCLe/L+RNdOhXVoKdGQA8dm8BrSphIwWHBxEQlLsc87mjs2B97
2RQeQ3K66nhn0LacC/kxfJjeFdC1hZ4tXDfd3QR1GQYmZPNw+bn785Eqv6cYl5BrJzq2oCChvgZ2
nP8ZDlteKok/t2k6l3EX8V07ZXkt1BJo462+5f2pkrqe/uAhwQN2ezZ3uNDGvn5b8G6M9SZ8AoJl
UkFI/tgLPlWL/YR0HtQ+eHt87Sj1vZ9ngIH0B4RvsvwcQpPjJnOFZ00zVViZAEO92msbl1QMEFz8
k5ObsqeK7Flz0g5ILiDI4k4+f37+k/f9ceS02n+a5QyFXBxGV6pC/QJisHK9Y4ynVlV8GjyV1TU7
dbfDwiKMpf15t3NDEFcL3ZEo17+w/w9XxukKIUko7DeEtwkFhU3C330smpIz1VISQ+OyQNpKKZxT
NAopqFSmCNd+qv2JQZ6vV3PZQvIzwHD/iieNLDdWq9GLz4fAztKo52KxeNKLSHb95If2I3igGDV/
MrFN10uFSidr81MjMVVdygJOl0QiwGBKmc1pMr5SaRuNOE0wf47tDwwAuzXZQ4YJjVt8ho36gAAs
ZvywxT11cnSbWlqBdd34cIwqJhnFeysTRBbdk484Y0k0LqxThkT/x9aY8qlR9ZXOUcxip13h1Qkc
wb1eS6UAKsurZ1qTKTG/RbTjA4ccIS1f93VPpfsAnRiczeYYZn0wUgg6Y4/KoVl6NX0EZMvhtnmn
BJtthrs8WMxR5K/viepgXjXBGaRCa0OycMdfdJylezTVOryFe3P1RI3yNyY+TrIXHINix4tOUftm
qOeJ0g06L3dYqTGqE3DMID6ppDMu5t59UeDaEBkIGgbVWrb64RJh9XnfLlx9HMjMQkCBbxJSC5UK
rxVg/l45NgueBAYnZZcCDmMTslmO1sC++EQxsoujU3/egbtXRr+KP6SEY3SqzeLUeOK6OAMngoLd
tPyIukY0SQp0A5rzyTvnESYK9S5b9rXc8X/thaw9GrpmvIjuMSXdbiqZv9GSH+rtN+qKIERdMaVl
RjJvTcg+J5Ha6zwg0/O+Hy6ycpOth/5mktWDEWNyzs09Dq5NhUnq+8FFkw86UhcJeOu1QPACED5v
M6O+f1XH+HxyUGjIrmyJCdp0XI2d2qrT+f0tzabmW6oo1CAmBwaiOhABsHCzcYNDnGNTDpQeMPg2
kAavcCGjPNOmaKeAxMtJ8prsPFGPsMG0b/yEG5gs/4u2gRU7cSuaIc/28STga4zpMwSWOLnPuykG
Mzxx5k9uZNlI8ZW6gOiEKqVzvheUWQWyY5WFjkH/mvrwSrDh5cVgJQLLxi9wqjZq3S+i4Av7/4XZ
8XHIUTIa6+qDPhxsO2GLG1aoc4g3CZqf7S1fH9Z297QzRS7eBvlY7UKc3ga+fjr3iho0TcxiyhPL
3Pf0opyPBZrQ+KaAo3OterppKIgQA4lCnLee+7HNa4xE+RxB0SFY9PBh8d4/HNy74M3tXklDrHEc
C/DLVaf7hN1AqAZR7nS9ZZyW5pbX6leH9aZshzJHdii2ZLV5uyL5qDdKoBzcghKra7hVKu7N5xjn
lVtbhBBFMzhXHOTUGO9603POJyQj5eEtD3Nk2F8WWzmRcLybLZb19LNhrlC5vAtYfL5EwPuNjy3f
z4RtABU5PcQ5sfndqXVBf+A1jFG6B5/f1NCOyUScj4Aw8i+hre576cJYiagusgg6vywOGBQVlzTJ
d3+wg+ufYBUjJ3D8aTwbn6fjfTcKwTx37jagUaKcLmLNr0q0i1F3SNLBahQVYYQVgnhmsiM4LeTy
ZF3nz9KA1kCJSMCYPOjDJHW4gthPagqnHLxmzrj7eihFuiDVBb8Xm8c3bqXpGRDPHS6nzVlB2Kjh
jw2rjgeG4T4mw07jKKtXCX8yRNDJ5oaEEBbSu6TixShmMCCoewN26eHhsppuw/xrP38y5TMRzAj2
svAqcE82IZoGJdsyG6ni1gKYk8n+kfVbu62gBigzK9Jw8p3EDjluZfAFTzqccEUpc0sXODW2JcmB
mHoxNuWFURsgTrC17/GVtWU=
`protect end_protected
