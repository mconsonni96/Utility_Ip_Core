`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
QbOhK2OgjgAmdhRWRzQ1vjMXycOdby/oK65R0qqsrGChAaELCzvs6Tllnx3K+IXZ6Nr7tdtvqyd2
wBMdpqmfzmnH7mbAHCLdNF4WIehqW4PujF/aiUUcPlUis5Z1iQvdL0pKpbNZfpJK9Yd2OJtTZ5KE
uuj7WvjZWTY+wINbfa3K8MBmT+vefc3GWtSKyFSNnCv1I4AdmIt8/k93rkn7Kdqgs6japXkQ7wYr
SVF/BPPm2oVzZ4jPA4nB1F0cOaX6yB1ruwJNxrx78z28s3QUIEYIoBQ2hTR36lxGQuxQFteevUm+
zL59/JM6JWHT5DtjhBlghunOAzANTabzSGIovw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="m6kpP4uHH5FA0szMz5nGNgaPeVbFCLyH6kj5ArDsP1w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19936)
`protect data_block
+f2WAMHJxJlJN0tjmwElGCboipA7oORjzfyqoQCW3FkBmCwBqOsdsqOu+wnXHQ2ItnfYyNiUd3yA
vTiaUijCWZ+MUeP76m8O4dQ+EuxQQ4eIel8D6v61U/tEdTcC8Prw0vtrNXOmvRMnPnuN4YUc2IVS
aPFrfRW7YQiP4bpS+0Cjaualm0oSylnebluaI6oNMtPdlJ0QWOkUzvpJrYlRVWiN2JWUdltflzr7
dQALrnzHecqieBtpg1vX+bxWM7TUTtSvYFM/84ITNv0xivonq77INTWYncX+tcVEqODiulLIsamT
BhqdLKTWKSB/cyEaQQDSlc7uZWIIaxWuBTwdC6Hk5MGCJLRPpIotO+M4pOnv8e0OKY2S9MoDWAiZ
DNoKBis1MUIl3CmgC0hTJVC4k+W2M20NR/nORGr4WFd/lIFVs0gQXZdgx0uoeNBWwHb2sZTjAf/v
5GxitP7eUoTl4bo+0UG6y5cw3SbcVZvgQS+hHgZqnUIIbu9UNO0Gpl5J+4H53pxElQC1BzGIaMtz
HrYGpIPOyLNOPOYZefCu4C2Tfkl22uNqV7+M5jg6WUZ/eW4S6XRs3IPwdalxiS9do7kS4QO57P3S
dgQtIA8XVXPxVzUK6f83Qf5fFPsBapjsb8ithqvXI21sreCdDNsO4/bnQtu8oQqA/5A0hPUFITcb
eFB0gKD5aZvABma8imDR1svbkH8/jivjhfkADq+xEud19IyxhGbfRiXYkBtHpo/APTAIT1tLCApS
UeYs4BAhFzacOKDQSXizvQZyJcq1Yg2Yete0intoW3/MdNWN7rv6LFtD/fD9EiuFYnqe3OC4jt/5
SRqZTFQApUWcLAgZ1NvP2AWpFg3Fg9/K8H5GmTzAQ15Xy8M5m7S4tjbUOYrGrMnCwvXN8GEX5OWz
Iu1BUtbfpEgc1NUuvtE0PWhsl7+xVrJ4WSlIFl/hMJQS7/Gpyl7YmJAybA+p7uNnFFD2gJKaq2g1
gtjtJbAzziILmHEuhSNTNdWTODq6uTwGaGRcUFN7m55K24oOZOzt87VstOohxanQJeVu9Y139/VL
MxNVBzUKyDA43efzYm7F23HkBnZpOWZvLOTsT7V5OTeb1s0YpYFlvt5Fo2tYPQcYcnPeIoR4RgNg
fk76t4UYXHlPxSUReCi8Ilen/x78jU/yIpJEEOAAI+I3tQry2uwxntQmUGDKl/57AX3QlhX3N79M
xBhIGHXSQGtKEft4C1ML2ggcgHSNpm2tqQcIQyZu9nR7+iN/HbYLuSfbrlwQQMzavIUNG3EZL44O
MFBoFgj2xNLDAsgTFb2f5xIIntQabr0qCV7qsMnf92jtwHilZFkpyW0guQVT0gslRNZTYniQU0du
YWmnkYTwr9w77SqAjvoz94rxRyTMZAx/JSuKpVYpiP4SlfTo9yfdH9y8z0qx0N9Mt9CLGS4pIWpM
AQA4gWRXo5bwvxzc8uHLNI+6GBNSCk+Y7AkfEudCIlcWwdzxmhNfhtzvA6E0/ag4LZ1jbhcqeAfO
HEZGMWv/qgY3JCtuZppo6rFFRGzGvJDERA/pMgjQQSdYmZqNXCGvoThgQ1cUOzLMaH19pRA6h387
OBcrbjPyiD0S30qb/7TtskVJxkFHvnCW1mAdfVr2C9HU8/6r0IcwSkPKr5DPXBy82YxkHQqJVmun
yK0Y4TKDhiAvv3K9Q6+nHcoSvb7407C2X/IOSIifaxm08XEImfW5F+DV+IRCwv8iAHctOK5YDHIr
gX2Ip0D837Acm0k89TNGQx+CJaVIlN3S1Bdp6FY+jV0mJgkKKCAKa0uXkiYfdW+25Dto8dqajood
ICHXrbJcNFXurteK2oiUvJDVTP6UrOALl1b1u55fkynfXw+5j0mt9NPLJtGdDYOblvaeBe0Gji7d
JyQK7Shrf+4Gwlm5mv0wn8pmBoKNEspt7tluzDpqhc4dXpkdcK6Z9cNbksO1XX0HIOvQFp9ppfX/
8uAvFP4a1LbwqQvuhNH02x2m+qZdArGob7j7CKBaCfbVp5fFxDASwsZ8ZuXM9hPW7yz3D1DKtoxp
mwQiw47S908N3mrRUgm9840QPuXR6mtSvE3IiRzWepHtrKxLq5+Llw+ENafZvGNtYY4i/LJpOb0k
rTUYBtFckhMhPplY7monqNnK0i/8VjZVKvVdgXXvrkPPUwC/zYpHL0gTZOgCIxEuhb6oFxiCEKsU
avaLWCSlOC+VTa1rxgSRvepFuuLic7AkYjQhGaEXyI+Et5rHb0F+mkrcy6EhreTymNLz/VOjFcoP
A/B3fBtW6aSZcU/vTwW8H/3BntMsd2UPSM0aKxhWw+ats5oThHL0yJWpjeoFd+UJboNVKLUw1l/S
aspbrhW+0tMYLatXvWgyhOIewLxfBhLlrTe/zjL0wW22RalS05wCmGP30LcsIA/G0U12A6KVNXsF
EOJ2+TsKF2MsNKkWLLMj1Calub8agKPK1ePoswvc+51y8Esb50VWy13r/nslARS2yX+OfhNrcH2u
tgCXqva7ECuMtjW7ztsBUKdT3j8pmpWB3vp1dyZFXeZ/vbE47dCOWo+owBloCDPtbItlhJC8eqLy
9IfzmWocCbKUlVdW/TtGzw2NdbJzDko7mN3+a/2oHDVwDrZl8Wq6xY+d5W5Sh5KUJUi0fAOlp3WS
MMUhBfq9ANwphs+dgQu8JaAxSg9lxfbZ4rLEeznZk3J+78/VsHiLK7eu94lb66EOt1ODZdYECUbW
+j5P7GVEN/9Ep1TkIBMuEzSn9Km1xvqMiFVFA37rbJIFqUHrv9e1kII16tEz4fCjikvWesKbkVR4
DoE8gP2ZxMKnEXPxIG7HW3oz0FP0tBnkFA6JR4G1hdBK6NRVKTefU52jLPLeBeBV5ZqeSqGIhfp0
PAVWzErVKTdZ0O8bsTAfn8P2DlAZyWW84e2U9PNz4lCya6JUCjHvz9TNTgmkqT+5f8/fJiR2wP7X
8qOjzBNYt2lNuKg5Q25KqHFA5sJKF1Deg4q6OFu6rkFY6gEBAewTYw7zcUjsm0bVshY4P5SdAwSZ
EsWyN7fKdv8behYcrgnVM62mUqFW5GXN0c8jR3LHucYWbIFEAIlxbiiDMfE2LHM+Q0cO0tVvBGvs
kn4AA+TMzrvLKV94+D5v7pRaKGGdiNy+EDvuVSDaGI1DUTruVZMfJaFaQMC9JAcVcylFsbujtm2P
w6Q+D+oKwGtZlnu1x2LSu5IkRja5ATzDXaV4ZAj351UHjWrMH9kY+5Dt+RsGezrWkZ4PaDNUHM5c
YYSR7v1rI+aFK+if3IQ42MuqmyeT93JFvZYHCGVgnRvapU1ZeWZCtESocddhaR6C97mV17dq/5X7
Yu8hMFy4MBYkY2A87/IgLk00DPZVXf0udIc1GDqloapb+qZrPEL6x/JEOtHNPR+br1Ao241egCqr
R8rhhjoXgHPgPlKWIQrnfB2aKne5sixnI8KC7HuQMhbMCEFCH0ZSoopz6hi+33uxVczhlldfYnyB
QyztQRzbXIcnGhTwqDAu6yvCyvEUvIAjM1dXoFRO8aCLgHlPf9H1edZOJNldJ3r2Kfa6X/MK6F7+
Ykvlmw16gbmZF71Kmd5AfnIue2xSHxuFHboOu0dktWNA0DZANFgehfDcHmdY2+XWJQJVuNdAG+Ij
0xKUsWNwTCIJaFUkr6TwPJnea8TwoZ8kVcpeDO458iLlCVQrPLfMkNjrmXEd5dCzqC3fXEoIXplO
R7MRPeicTuUBrRyww6NwNAdCX2qYIv1oF4HFjM5dM8UotFLwC7BKNIRJodGUb/nExY7g1kesWr37
7W1Ms/vo7bIsPN3tULU7RZP6xF0l89TdaFC8Q99147Ec5ymnDv72/x8egnBELHqHAqWUdC54fGiL
CbTpxgqrpFf7GbHaSmHrV4UdKDYUSBjxu6uWIzeuAOOPja3ZKVFdLO0XmdUfa7CyI0qUz0SuqRF3
FsNzCHnZUFbzAN3zrZSFZEMA8DV+qsmbhrxNnLrNxnI6tkq1D03paR/4dz5OVLpbRgTiEexfUSfI
pI8W9EFsyT+0Sos8Q2KdlIzgoLk5/6RslDMfV/C3SDJXq/zDrJRleBKEu61hGFoK5g/izSNiZVmo
BKWdHTb0OwzVONPEKIM3pNXclXr5fuCO0HtYVHWYVZ/2WoVcBHXtVnp5TjfrC3uDcABouHt7RyEW
74gjXQLnCPaxwhHt6FQRpgawf9/Ayg+QA/xPVOB/Nv3dcgKEt7eAEteOopZDlCPT3RSU0+ANksWr
U/MXPQ5IXBjle1ctp69HSZzNT6I35OiFtQGyf4PcYWIF1VCn5NyrSuG4gV9cehe0hcPDBo/D1wtz
j7TZb1tCPr/w77jDFgec9p4eBVdSgRSNqArPIC202+h3Wnczkb7K/0fTa0K3peXW3TdxAWcAj5Yw
IfQhmDGop3vKgQMvxjCVvzQaGX7G8RND5x6kJWv26M5DT3R2BaZM3B2f8XGdCyFf/SEHQD2Idc6k
YOHa1Mcc/2D2MOjmYH/h7SuIk8Rs8c8DEoKoQY6jUjrnUwpheO5gCHz3O2C6nGfC+pDRWZGuSJ8G
LYPrzlr3x7niK3EGLIt5CXsPdQyu5ThIto3B7q2u+CVIyuXXeW5YxWOL8wrpo1qA1CVPL4vqIFTd
Xg5XYlXOVxwq8JOsm0WhDB/r75Dzw42p/ubfTBtGQZGDE/46fUWiN5E+1Zb+UzpxO6fqsYVLbXcZ
DQGM6U99CTljiUR6hpmO44V2ntISX+Ftd2nbbzfddFrMdYY+WqalF1vRahgkiz8m6V1I9fLMJkZZ
dvYn4xLXnUIxmYgnQrSN8BPWBXA68EKlhO9uMR78l/8kQsIma2XDy9bDRkJsxJ3KOcPGXu2q3AFH
Oc7QR2i9dUWw4KNRznNsT4lU3xpGw7fRiwi2CXaaoO8Cf50j+UksDsqBsOzxrVvK3cYTDnRZhV//
iYJ+fayVp0FrYlv3wPQ3kJFXk9uLKZCdsqhqCtU5CWYfTENFiLcIjjmCD3TqY/pGLXuX4fs6bIvB
SJGPnk2I/iYCD2ZDU+0lPNawzDGkeONnzP4pXGWWmt04NuQywIRzrTTi8PviUlDO/dq52Umh9dUv
SERu8BsXrK+US7Jayii/irRKpgCcdLHVj+1umVDDk625Q5j2Zb2BNiY1rH8pj179YjtSbROaULLu
yEIJHqwvAcje8HDjzFtOLE1N/S78KdbEYcFp5uCkdyYGlGs/Mu/mw5x0ki3YHda1wFMIZ6u+q+mS
5Zz0py9oGZX1aO1R1izbDdH881Drr0P4wPvQ/1ruFUd3+NuDOS2yJHsOxRJTOVBQvpOueLEg3ZeE
++h3HAmp2LjCcJrDxIPRPL0/BbT0n8pm+PqW7drw703hpqWh7Neglv6LCIjMDF5GJrkGN4MIuvNQ
gLLVWJVht41ge3kQi0lRJhU9HtCKXo/CCxSK2euTuY8zd3VynBopIsRQhF6mw6YUYnV538/Bf46g
JVB0kSqDbvOVAcW8HSSODcE8M1cXI8zGc/xJe3TfiruD8Cdjn4Ua5zmPfA7cz30rRJBvF2qDt3XA
GYqScJkRpRDU4v+a2hRIMPkPXc0ASjsMa0HsJzD7pMLNESpCEM+oPT5NBS3hSo/vejmf4NZb97Ig
JlFldgMq8FiznrLoBkHk+mobZYC1qrvGuXv/ErMiNE/U2D0cUQSJ8HDqS2E44LCbk1dM16zLmNVZ
o758PQWMALH0o0xrMsN3pdCHDh6EIOxf5UdprYFr+XfDx+A4kcKqMXDnUsw8Ilm5Al9A6ubnorxe
oHlgZ+AGE35sJPJUCa3WkvRYSqzvNTHv9GpHIC4tW9fPwVdjf+ahujh2T0o75UjIDI3tvQ2/SfL3
vAUTcq9ErcPQi2IUfLbd6zxzFI2KGl0GWbDLHHW/3aZtqpF/Lx6MeS4KVaDfQbJ0xwuTtfy1SjG3
nN23TZ0VW61TaamlDr7uuFcqTq8uviXKd37CGPBV3VxYbuHlqxOaJyJ38S2RilMP+tW9wwxCUKfn
lLo0oVdSmoWgOwJE1zIMW8yKcvl5icASmcACfKoOETYwCLel3CZ1ojaCRn+l+l2BpUnl2oLdBwcK
M8k7f8UvF1io0ocKs6Px960mwury47CLugEJht7GrSk9YQmzk7kf9g50XMGJ6gIdDbpxIQzahGyk
iBNzByU7r1f4iLUUs6FkA1kdXNwr/Phk3md5aQfwQc20yg0KPpDhooLm1YURoHW8R7bQT20xnV1U
qkYgQIyA+M+xgw8Od8bDshaTTTrZd8M7gPQ0UqaJVCOL1YJQg3NAkeZ2HTBoy/GxodgXioROdpWP
WpGrws6l8aS/mKG1+Bk+MEh0sbyzhUCsYMyrVYWzgN/vmm56NAfuwIcRXChIE+Smb/u1Uy/IUU3V
jB24YN7jV+yGauuJHc+lvhx+A8heYtOAqY7yLhPk5fY72dnOGNQ636HHASi0cf8lbFZvtWAoNnBF
u+yPvjZhUvasvVawElbDy4Rx+7z2+tPHL/RPwPvrK47o77MdSbzq+gqTRI5JM3FhZdCQ8Wdv9wry
tMCZfkLIjP1xHMRv5LbZ2F9NYI10Rb9nRfFo9ZCzwTKRq6P5GsiSrmnFYpcHWk1kl+GFxA9xFp+b
qt20+/UMUQFLbHtgJW4Vz4jR9CTLPxam0QDi0ScgR913cogk4NxLqJ/To3CKU/9nqpHTOOS6Rfk1
zd0Le3g0QpSuqOfUe9bgFzjnFPkbdWY/cxCTGHR1kOXwiaMMlOXpugNGqV6j5plDBW1BGk13Yp6S
kbcsOkSknBCcGcc5PP0ciT5DBRlzXyaCJAz3CgbIB5D3J8CTfhzZpKV3QlPaXiQk4/oae0UlMovv
xHeDaZI6FWHgD463zcdxeWnhRtKgqZFiTXTeUmHEarKFH4wRXbQLNwcE/7E/zUYBH7fqaT0ePlKh
NsTaysb92eyTxqgqSnQbJyffPiOm9GBiNsswO4H6B16c0knZFe5b5hQg0VuQLBJ9QG3TB4lHbgLm
ni/0/ytLcmvF7WodbBiVuezxwegki8p7LuLNCxq2H/m27SE0kEnvdjwm2xPeFNDzSVtECW+1Wy5q
SfuU1U/WXxgMdiI0Ph3Wg0K6m54y43QvEAIhSNC3c5yqB4C304ZK+g/vNY1wasFSyKtJBD3joKG+
ICDU3Jiw3SfMO5JOzT7jbeX0Lf4oUGVjsb0jvZWTjMXWE+Ln/N1Cz+mWy3vduDQE5aTUNcYC0qB3
UpwD18vTGgSnugwfbf/nf405EtZOXQFCZmScsa4QGCdUCJa3oL9qw3mvJUTrsvym9tJuE1CT4Mpu
BOR1XwUcDo7cgTHQ1ExgW9h386zqLjxvjfSethTBt1z+uh35WaoTVsgQlbAvXyx98Aebfr388LFD
IZvcwm4tAHIymxufGF5hO7ijQ3wcQ6qZPxzZ6JISTp+moQeMeYaPz50LRO5Hgjl+8mSo5pqFX1wf
6C8h6t2VG0vT28XnwFknss5yoXhBOyJ8jBmHI4xezX43EnDSmXdhei1tmH3ujmg3I8kRCYgxnzef
rcQ/iA/NUBHENGMQMgvWiy4M4IyI1JeJ9vmI4KJZ3nxXYELOFcTEsobvprymrbA10DaCGSFYQn2V
CPFy1SN8koFlKeTQ7vk8WCqBfia1hreFI7jkGs2xdrCvpLKfYTEQvPf93uN8lYG3ZVLfbuDybMYx
5LL/bJobeb4fpWI0lYdZ7QnTkFbsPiwFu+Ke1j78CiIhk5UQSVNdxhpfXMm+ShoTNWNbY1Up0ATx
iIwPdlTWz0i7RGfIayuRrOGEj2vFJxITmlQgE7WKz9z+t08Ap2Y6uB5DNp3aRWM1z75C1hr9fBIR
A0FVqFUOe8ZUpTIO6faVTc79VMT9RH4A6irUyrcAXSER06b92HA/rmfJlvpCqCeUridniB5WtKR9
t8/bFK+xKj9HYaswMvsZLGB8HXNSGMvJ/0F+qgx42taAI53J6DCKhgHyRm1KNGbypbmx5I0/faCf
SGE2jF+PllZmGw240fPiBUzmTgPK8LtWbpvP+DeegpdGNPN6gwb1S968scg9uy8NxF1DSZR4hd2t
70c4zuxCVOgEXgIeDwaSN/EutcfFO+GQ0P7NQV5K+PYGBPbVALFhxmnzBaSHPztc5Xkt38indNuv
Cs4zo/uwk4X/cC/MyfK14x5KlZaUjeGTrWUeXpsejWOwDaQ54Gz3XuznPrBNZ/OCgbaBr8OEpGir
IV9tutY8lLSsQzip8AWgyGaEsTQIXRe6Hw8YY5WFEyxk2GEbWBUqVhfVT45lH1CBetcK9V/WvkDt
CKJELQZmh7kZz2ZptkfA1WS/r3/CL8qxHPZXmFsU5vm1zHuFTJn9xjfJkhXqxrSf8kQrqyyv6IW9
AdO97EPVE5M3fvTucPxfIgkIfSrMaHbl4Yy6IAIzbSUs3XU3llNFfzzwuVS7bzKz5N1nbIN4GiAG
mHiqgAgvSrUYtJL9BzbVz+xvgV1pYv0mkrnx3h6Kb0+SQFMke+/BfxRcQr7ZMHufOEizHi3Vc0AS
4el7J3VDdS4+xYr32nLr+JhhA76DqYP9UTO/s3rcOVrXCPKud4U3Qh56ffDWlYiJ1Yq8NawcdpSk
RUJTB6vujD99zVKfp4bMzH5Sab0+fdFLPUlh9dslLSe/+SqOvLOp8qmABfoosLdZ1yHY/8NLEKlr
QGPab19SotyleRYnKz7cDEBgEsy2FZ/AhovkJtzmDGNuTGFIZnZwVed7easrVHLZtvNdo+rH2eFU
FqxzKkpbWQNLgftZ1xkNjwap2MzPFZ/vdHczqE/bhEf/9gdB4w9KaWhghkE1gTgn6fZudhDQN/A0
lqCi5SlFIjt3H1EdiKNDoEkSmXg8mXjrMRVpBdIL8/wFZYiyN2SMAiyOrRv+lE5U/IgT3WM7xKnr
kXbN5pKVVyR2HCHn9YmQDndAOCg7XRd3fQkznvqsl8zlZpOnPIZwjcf5qfu+eMOdqUXpfwhQmNmQ
eBPw2Que7wqw4u+iznSkEtsLxZSMr2icEYcc+5sabz0chvGQeyrHCLc3Zr1mB4dSbf/5suhhRgbL
zNEMplMxIA+CbXu6ym4oAgVP8YMZmuQMHFpvWzrBS4E2MbGZ5anFeI7iEGJk8fzVaOvKLcbVm8ho
D9Nn/5WnTUPH1xhGDLglKeU7WOlZjoxU/RwH1ElEjr5VDTIZi8YhpDS+d+NasTMzELJ4PUnbywUb
3Nk3/IK+A0of5NWCSsnRbKIgFSc61l1Y7TyxTjWqitF5TZsCs97uSt/b6UchO08YTrjM9a/fVUNN
kFzdmqvKZ8gdt6o29INglWlNn2NWGd2+thJxLT+pcPzNPQQg17WuPtGvvdt5DyHd4bYzDSSS3P3E
91oKh3MreiY1Wwzq5zZtaBG1Sk2TXvJYCgLN22tyly7G6C4ngj2zh/x7bJL0n5mPk0q8f+gFrSrx
naeBlMs9adPAQg+LiNTjyal4vMIhl4UYcRW2+kxGr1cI8ih0l56JFTDBv+Jj6u5S90A70dYOqekT
CciUNEbSqf8IYP/M18NdV1NBDvv0iMWJ9uEETVYKWlqWCC+7aVWlo6yIWIcHc8pU7vsP9wsH71UX
p0GyxJdjFYbimsLTGJx9ejqJDhyRxw/gx9UisfIDRV50+2+tlg5DoldwW1ra8yRZz94XvM3WxXeY
eFANKQz4HZ8M3JpXTK2hzuB/NWWLvXvX7EMCIk7ntljG9NYd3DWsBYTxZenp2nQ2EbUl1uzmRF7z
bkhoQ7+cTPDztnbxcUtzKYZAT1dWpLy4eXmR+LDAu3M4aUZ4Po/X46JLPWFTkHAKuck0DF8xxM1k
7BzIHc68yvUhcvyC5Gxa1nIPTPFTXJuHFRsntMjVG3NxgFd4uIwiuHsI8sudMALb7VA6GVpI4u89
8GSxYVtFcUGiLAnnJtB711Z2047ZJBJf4Dk6y4AY5ii+qPi9MVjJIQRo4yslN+UvdKmA4hr/1lZn
i0tUINXayVmNsurn6/hi4wJH0bM7Oa1k+UKvcgcp9JgKY05C96sui5Y04fbFEsQqsdaJCaKYBgo1
MgNRRr4dd/zuVmTStilriOQ6KSsdZL+HIMzKcw9tWXGFNkyM3ZQbGJScSdz7eyMoJZ0xaTDR6cR0
I26sZDR9E0GpIO3ADUpb2GA/O9+0ns161dTuIWO7BLtv9ZguKqTvn5JE4xwDH+xe3ODhYyLoe9Cw
wEy8KUqsrEurgNOK34Ivz4kaCTf3KMSKjD+0PspCJp13mulnTlnuWx1yw/twmf1FMAw38ttS5PnC
dYuR5/ykjA9IyoDDMuYZhI6Ze0sVdVmUqqA2pCtIhnvnWiCTWNILFucWFtCNUEfNjfJ/lUgwOmbv
WdOyR+3mJRVTnWusfgijSSSF1Xd8zcM8NKwoFKlfZmuSPkCnm/R6PGORtpkU3MKO2z6OdZ/zvV25
sIu+djgFR90CpnppdYIqPoZ3uPHUOjNPrzPC6bzUYysucc2Fo1qwpWBBnyKcoKTrMOdlVtl9I3Tr
a+h6vxXwRPw7IsqyTNNq9J8wsxXIp9w58uUOL6IfV9GReH8R1PpoMgp+jWK7++aBasfkMpv0jgCP
Xw8TwSNGbbNKP0eJo0gXA+TjPmwhYos1QaiEKkc4kmwcxWv6YstsCndCDNjC32IfDX9G7LjIBwJV
EL9NweYCnnQqpalHBGkEhAjcfBuc+jjQ5+WAbqpi9dPeNL1juIbH9Zq4g6QA6hMlfnQauZcZfcRs
iitqtWVvrMOKuKmB32wZkHnXpVEAvtMZPKeCyYIkW6KjjhDL7/seky3jMvb07wvo/jHtGWQUC2Vx
Nc628chKWHx35UTFvJlT2WoJdlrq/+qMGBLVOh0Ge6Vd57UpJ9IHRdhqWxMJchY6rB0557bWr8Jz
Fa1V7GKlm6HvaBif4CroEXyX2xPYSqGxdOAR1FCgPnvOCZ2jt7Vq+kWeuo50E4i1Ts/drLxMI2d/
yZUbFPgBa+aPd6jKIe8NjoAbCpmJeTTv+fk5cX5ITzFbOE4653EsHWXIud3BzlsVXBqWQY6sDeKW
GRE0ZQW7LiYYB1eiND1EX2xXx+8sJXrpiBnA3EGUc+8iNuDxZfH0KS2wwU/AoPsm/DXBR9KcpHxW
durq/rCsMVf+t1Ha/xJ75PkYleXyxyJfiz01N8TjFJmHXBbYf7jfFd0rnk6XefTBGmNeVp7tRobj
c4sH8TXno0l/qWDtvOAkAnFGIJJSJ2Zp4mDiUknba04maj/3fGdRW5Mmm3H4HVQsbr7HIW8al0SL
Q1EAlC0ekCYIYZm7gn1aovOyoYjB96z/6yRqaOL8o4+p4qqs1Kuoh8ux20nWW67fjVfliOCrH4VL
jMjq2mnM1YnTDFtFYIHRVBXSpS7gfrf/KQJv95ouMLV6bXvAZqyTCRcQirM9YVTD6Hp9+Bi/s27x
Ui7kBglv9qBqvJOO+LhqS4JXn+mAkcRsYixaqQEc6I90MfhhZ3/YhJBSr0Lu9Ni/01wW58w/l6qD
jfFv6Ij98xf6IkL/PQ5U1G+S94njenFdqHIA9hbyc/VSzyJSDPkBhhgfDaKsKXQ6mD8EH4dPYaBA
hbPH7hkV7fSeg1Men0bsUUuz8CVvIo/hKygh9BLC26a/+hXeXknwEGWpnvwufeWpYOUj6W9QUGvP
BS8l5SAIwRV+Yu0fGF+tD0cReREea5+iGhOnsrg4ZhcD4o2s/HlwTiuHsZVZ0GOmo6PnnohDG5yc
Xnfske1lhyc05TC1tru1nPUuJVtwCpUk3/oq5yfMXzQx/Ci9YzT0ha14WrxSCSplFkDQorrDsdSJ
US1VGTYxjeJGIV/R3XUaY7626DelfhZa3QAr8sQhOp9CVdcgn9KqrFOB1r60HJGGV6Q1GXJqvWRT
+wPXGWYXtNM925NkOJUpJaf0zfAdCD3dFL7DbWhFeiO3I63ckJZZdbE6dXPeS9ycpb1IozsqjWZJ
+KXSxXI+YE80G+A2jPVsfOsKkbkOW2vQl/b58i1SjVWiO7zGjaGZ7xDcqsiP+sBfdMxslDiAb8Ek
x1l8ZATV329IRTrvChxHa3t5NSl8UoE9WyQfJ53qKamdvNQv5uCU8HZREsDgW+IQ3XcBfYU5oCpS
nf9yD77yv/LnXKXO9AOJ1dkrc9+5FgzuMMQ3Cdaf9Xs1bo4GS3dy6TGfGuQF5v4N9RpdyktnSs6o
8Is1IOSL9hpYWvanZdmpJ7seMdIMMvOobawlzAFKnbjXmztFG5be9WbLOkFtSIKL/Klt6iNaNKCy
/3mfwXANLG2vPrveJYi+0ULhvGV4YD5i7JTAV9urI2bQzhjhEE3rFq7H2cPdK2Y8WvV6PnxELoCQ
acIRwUd0ZsQEMIMxW0VpDH8GVn4XaWt43/j6HP6AcL6wXU2/IAqVwmu7wpobZXweahzhWGuva/v3
rfd5gefaZ4EyWsHDoZRGINuYPRfYgUR/3betRGZNomma429980CvHGCzjVtikw2Mup+90p2ISXxL
poGEZQmrDANKpLujNtYm6AOqe2YdoZgVhy1bTz9+ZtBkGRth8wBYYrZHkCGwiqXw2VV0vmVyw8ih
PROlih7vm7rSrJSljmFBdkyTKt4+vbWhfFsN+Sk/yRNK+ac71yTRP/MY4nRUV+UAbunc1Ta5djLB
fTXyp0xiPiywe5CL2zUFacIodjfq15u6w/1DG9ZcsRpeXUq7sMU57TV+6+JanufVhxUwxAZqraWl
cX1YSb5v2bCVev4Z3mIRQ/84+Q35hys6ZERyP3XZOMpttbBIo8QFzPoBPzpvMjpI+Jk9ta1vyJLN
h+LePM4P9W4kAD96qHw7sx/FBZSJzsNumGRZfUrWZrbmYmIJ1VTGVdUHp/VmWw3fpb2qGBAk8H6p
wbbp2qsJIpSqIZmAczSjRMd9saquAulcHzPZAFHXc5CG27fea6BxVRlPPKHvLXW0DcE0eXfewkP5
a16153TqNbVNla3hOORmlh9wlzL9ua47IvTpVMNyO4xUci66RgTgM0lZuiRKGf2l0d2QgOtfiL12
QSlfU+9SIjy78yiY226Q9VOYzD5AYD6Ma1GoHIpxUKZmuLCzj/L/mdYBkYobIZwNaEicwI/DS+mx
/8Yy0FQOzvBU6uTKq2IItqKYT1ZJQv7pkcLE66E66JFEUpblK34bnDrY1P8g978IDihasBMYkdq4
+8/NbVs5euHf55pVv79MX1+gbHstkDw+CSan/aDBL0ktKQ1E2CXWJV3tz0f7GPrms9naRNYu8sG+
UihgFCESox/pJBc3mytrenbjTAYXoL5MviH3GsuRHvdATjeX+gPSeypQyTh4bsgOiBHqbpKwEjwc
kJOMJ+czPnT5yP0GaFB52SVSSrirzNMlM/F4t5NMTBxOh2K+MoQjOiZxlcOHQyAvy47rIJDdSEiH
MbF0rize/SwYr6SXMEVZObNp0MWOUz9ze1/J63vSTxXD1AH5jEt8YXmaKXR47yvK/FXWyC3dAYlq
Ue5RyhC0hzAatTitq+pCMNOrFFVq0KefEKCiPm2bps0XklqgSpodMeEqKZxzf9NpWZLVCzGS0cVo
pYSoSaTvItBUDm9ncDmxomF+8q+Xq5lV9I/Vu/olmHsrRsv50YgyBpIbqhJ9fIBI/Okyz2n6XCyW
GXycXhJL8uOUKfMxXBB+8vm8DBoER8g7aw19oUMVm3Hnu33/TIIw/33WSeaX8lkPhxdTphCJ5FAg
1sz1wNBbRMeIe0Z5JuB5Eh12HybyT80HlNOSpEoEyqLkx22kwcc/QXZ24Dtnnuc1Klpy2hwwONf/
0RMnjMRttsGjDUlGSEphlLH84Xd8PY1nJEbuTJX6tv/6Hf6LxHYb9XztR+lK+jXPbu1xD8sLgWNt
90lppR1YVOlc2ZCIqXWyLFLRyxhckPR88ml2SvKPwmdPyxaqv0AoksRMySlRYY+nWeUyoNjOXZ4B
l4K8bQ14HpVwFjwt/chmLkWHzBDlkIbtulur0/FCoTW9QQMY3HnavFe4l9I3RzeIWTLBY99sy96w
zpGLf3IHTZkqFSZ/tKPMhRxM2nLz9CQalags7QxkN8SdFYh14Yo+NrbujHJEGYShQEnp/laLzLzE
HSRsaJNfYEZEBaQaRCAmqi2xWT6DsME/ibLSgAEXoQdXLAY/10eOFEr+iwEFRPST1nCciLgR44lT
YgS5/dufPE1ULrxoCB8PomLupCRQ1Sm4mvXfk+DAvPElug/ayCsyp/wGHKoUenJf13V6M3sxVCa8
qejhfRWt+x6VCM97wmKdXl9JIwMUTK6tXyPKFGB9EhItV75cb1P0XY+whEU4b+XwEextmpzOw+dZ
z1DTMytXKN9cYsR5yTAK9lmN647g87st1cvBBrGJsyrMDmyggEGHaXasbBN16/eOiAoPmOvU9Iex
RhGnQGW/p2upwWEHmx/bZIbmPiZu8ECz27P1mLdUZq6EzV9ItLpafuAAU5moPZ12RfDisbG+4ioP
FXuJEk32FWuE0HSt7gYeGPN+PikqHaygXei2J6gtkCphtI9hNQuNY6WjNlJF4JSkthCjxnMul6c4
YJMyBuL1CJ4Op7E5mGeP2bLCchaLhuiEI+WEzKMjZV4ODKM2iQS5ZCzqNve32e2ccvKYvmx5pmpI
oBSzVJNhZEnWt3n4IImZFrWHoOucVuLVs90yUPkwCEY6KfGJ1r9AM9FF+DYNgaM7EJUlwPFnijbF
mbB1wg8ELQf6wgocXqXXBFPczPL/Q3btyoyq6GC61/XG4K9KvOO/x4dsy6adyokaozS87tYeeqNA
qxSZ/OT1ZRMeB3GuY0FRq/Rv26K0NLBrqYbi0X8SYuAgRuCQ75Z77rW4JYdSkgYFdVNOjQtBXezM
GazevTqXRNs6rYtxhqVd7oYgFvr8fwncdGzrUpVrRbU6KSq6pfWvZjeiEWFE2hqYZq2SyYymI84H
RYnMHDIsvQCTJ3vEjJ+BIv4Gnzf27bjWbMPldWYDo8omRpgEaubXQnARoqzC+AaCiuDT1l2lhc/u
cYXax7Hv6DryFKKzKi2oeTf+4mNRq80C81njdlhJlJ+MzST693pYzeoBZlz2SlZC1MdrerNHmeFx
wiQjeG2cE5DYTDugzJhFB1B/DVqs7b2Yc8MV3jOgJjR/fjBoUH3w5GnBFjtpo/lSawyTxg5tN7ko
2TcwLGhUq3dF1IHkLjRFeI/yCA0nuhzYOkAIodPOWbMNH7S1knMxSl37F/aD+pkDUMKlOwi/Slhw
WLGCZwKuTOHnICsZwcIF6KZIjt9aYI3Qx+NLBXTABCjuC9ljR/1qYALELQtrdus/EHSWvMmLqSI8
kdx2nYo6a7ggoYxoOD+H2Dft2YCzx2iR0eSQVrvcJ5ppz+Xb8Omi7hw1pBXRH/EFaRI8Om0zBn2W
aZkBjFVGuiwF6shN6qR/0TPAS6ViUgLlXGGez3SMqj0z94MLslA5pcSkb0rI6CBKFMi22e4Jldxl
ZKj240K3oudJt0Ln/AR9grorVdCfX1TswXpy+oQ3LwnvOji6LhBmZ9SMNCdAQwTXflSqmbzn4gPf
0QGAjxhaEghMvRvhHEUFEyl56SOMwPayzAODHzgJ69WuRhdgNSJlAUPrRI0jLDJ2gfj4CnOwP0e/
zNxC6Oi/nTRBpxvnimQRVy5pEcD2rlMy8HPmU2aEJz3B1K2JOxDS4Ad8WGM7Wdl5MeJz3C0u2Zco
yQWI7ElOvHtyDmydorpJmwa9PqUdAMNfxTiGKUIQdi8ExfPbNEhAv3f4cUeRB7TO/iSqsbt+eHwp
ItCMKhjQ+FixoAhce46Qf29wdYZ2Qo92SMap+4t0DZ4K9Om/ee23nzCjaCNSzO+86rm6Z1kQHC7b
UChWlJhFZwAJDx6WCaawQtDZ/xjdKNpBAWRIm+hb19TaKdHfyTl67AGBkYrdgJUMv5abRwAQJf3g
wejjpolw9n9szOq8FH65vThcEfNPi67jkL/yYCAMmFtc7Fr+B8CWG1QbEpvcYLUPIJfqiVtvwu/0
eHJesOxAP2ii/iUEbCJjW0ayk8FHkgkC8yQj/Zu+EiAupwbRmqkDms0xzLWOHS6wt6WHO3gbdTCo
3bIzoH2xNOJ76Ru0liSlL9uJLhCGxNkgjg210RpZJxVxIz7DHy4Sol9c7KP70VlNN0bwx7lD/T23
0Qbw2urPLJGP37xw21933OSTm3hyU+hMznaOcVOlSsVyiMF1C5Szh/Ky5jH/v7TlAGUuVT+DpKr1
jiLvy9NJx57a+g5VC+L1iOPNB6SXQr1WVpPgPKhzzH/Fpse88QfQ0j2KBq4ZyujHvFVINckREKJE
t+MsGrK8L2K7afO0lS1ilsZNRlFKbUfcwqniLhfRPDqZIzNCqYVF5DNrzFcQzsxen2tFywptj8/e
pcUKOSvmJvysmvdDWSJMk38KZGTDw2FiOWT0QEYIkf6KX4gLzPRtqyzmEzuS36mqlBA/pm/U2Orv
tTF1UQMAX+thTe77AoEL+um47H/+PUMvH2cAdjVMxwhSug8uGegsfAUleaMl85S7nr3Zx2lVS6N/
WuQ0Fw5OQuMMW18EFuy84nVMGyOTZxW97z8fGFhnOx4tIV4b5psGVlCVD0Wjhr+G4ivx3mIMWFW6
mG3XIPy1SVByM+Zlb4ueWW050aGtUI7LO7RhJzWcYRsHjAkgwg8BZOrYxOjvr1trQ+zfeh6MYrkR
8har5rFAl6gunPSDdn9F38tYtPCbC9f1AuG5na8Teqv0rmtJL5+xNwWpmIerw+VewGype0p/jl1y
WmteBp9SDTTqUBv3OmyltGMkFYMr8YWqZ0LiSWCtZ8WwvR1fMEkVEIX+nun4cxxDDs5/s/6sIbSZ
XFozQNjqDk3yAIvhFElx00r/q6Bxmk3H+NZV/bY3p1RweN+Vjcfa7fTVvq0DbZC961Vuhj3gaH0F
ycurjvhWamZgUATPJAR6UmADJezjYyT1oi+9LnsEx1e4XAnXjHcfwZCIFctbGTUCiv/ovNTWu17V
XDcQ1xvBJYOBQZrphpSemFpS+h2XJCHNQS7fP7DdI2QsOgjtidyn/hh+5KvSZNw8QjWgKFbYqX9f
plvKDrpukxga9NEmxJ7MLKv5UFgpP2nB00/P8Y/gN7CQfEboMDIg1y+ekOH2v5/zRGvcpj+rXP7K
6Wd3E/auStO+OdDtcLcEzlGIx2dNEUcdAlHOGg7pGBY+L7FTRm2pWnnWGrhQUsq3qpNRFwu7v5Ec
X7j3nHofhxXvKKwxJAOFDmnsbl0jvpN1MRJrfILh884yPUPIX/nEHammXE0lhXEbvEt/9ujRq43A
KBfF1ATDJ6MXEmfkPFYE6sciZXpPbh30GS1JjtRwwm75f68MF3s6C/SLvLEjtwNdzdC5x3G67vE2
OvLrKq5Cm/f+xS/Q9Ez6g5BSRt/n7shhzY3wonnSciub3CNzvkR/G4o0bgC74zJhXbq/iT4GXZXj
dUIAX/rid5CBzlCSs6KHbMfF2RLFpwMmZzWGZbBXdAd++hC+pwVOpJtpzEzuEbyn+ONVr2kpnCuF
UOB2WTFl8ra6UD6S89MUxRM9t6ezY6wJzF0ngKRPTvLVZCNY+tMRoDf76Ou3WxhR2x0SFWDOhEfu
raLZ3AOFHgbP52xiOdLzFnpnclVkWoHQDdr7sws0zqOTzmesj/1f7qLeXaJ7Gm14jYoX745qEP15
5TXL03jUPhKghQ2XToJS7e7+NYJVc6aQSzH+77B3sDyZKETienLDKlNwPvbbBLjHrZRwlC9CqqdX
8YWVcK69gXKp7TzI+Ix/zdAk+l0mPNtax2779DshAS/7go5SRrvA+glhP3r0B01smgsmwPgAgVKw
u+Ww3A4SKNao6WHEybv7bW0uWM+LfX503L8z5EHCCq1EJOXD8+FNQAeKRKQJh4rM2/mI6iwkDYIr
MI/2reUueLLOpOMvZvOYx0AtswfpHtUtvfFfE7tFdvLN5UtR7kj10rQEmoabYxmDIfi9VU0d3WV2
OfwaCmMvNbad4eFCBH4qWn8l0w2c8KER2ciYzdi8VsW0FNEFcUUhyrQL6I6nhNKcFN8vT6m8WzHh
2cCl1fCCVZOPWzf8IyNMlk+J6pJPfXGMKEEs3kO7YKaYDeYQRBrbXk3zkAqcj8psYA+XDXa++GSb
KF3SJnHgZlWGnmcDLhREZGf4lNbFPxRadV4q2LzglN5f1vS15GEyVKz8v1pMwyNK8Lb9c1ZUNRgQ
ib3yiXKK9pc14BZ5bnxHHEaRyCihYr4WBX5fKz1ciaWMmQxYrGdL2tw5dmYgCKzz5zAVdKBRGx/C
hQFr7sKZ5YtPXVAEGwDk5HDvv6UuHZ06PncjSXCbuTcfOuoOXT1+A4PgvY3HWstirymhYYIbIu12
BLsgE2HyGAweQjSCnVQoh2OuLzQEhQvQsaA5CnC8u/CRzqOQaS8/2Qrz33nqVkbhgn+zecyqekd9
TYBjg43Z+1sbfFuggHeH4qczhQpbl+x1T55x4rORmAnSQKcES94Ik/sXye0sJVp+oCByix6z6+U5
YTECEiRUqcXrZFL6mWXh6w3boOzzYfblt2ESW1TF52QnBLkXm7zfcq7IDY3SZLGTVUPDolcDSUeY
6MULnZ+bKeI1uvGP6BRBid6yh76SxQXOKAOFf9sR+l7HjXeIRfNoMUBnZC1yOYwOT3D/gzmLmTWw
+xjQPrd+To9KAzlxz8fdGv8zZUeqOpA7ltxcHOH/v/K03B5kWdoc8QlYE9GLJeWHpJyAltIYAiTS
5DtYCqPw17UzyLIuZ/iz4rtD+lI1KPjcrokytr7ITMwxCkU4aphRhGi+1JhyhimSzujNf/crYWZo
qpA1+GCdw3zJ7T4Hyc9uHQDpy3fg/wR8lW99VdG2z7fwESO4G8YcGalNFJVCHlX0UujoZiMOif10
qlG/ymRPYM8TRd5NhVlSk1g+uQe30g3o9dj6BZtD7NRe782I2OF94d+DWhi4vKdqESWpwJofLvlQ
BybilEqe13BVjC9UupUE+zO+9LVqppiwiTK/dQvC5oF9GeFWtcnbVoo4VCWppEApcukn7PetJn7T
z3Ncw76Nle6c3oFRAFhlwJoc6x2FETBUd1xPkRnDZZPXb7XyMgplmmve5DaLqAbffUhSQNnO0BOv
n4PmpyqwnZp/igfXCJz1Y5AKrxKg+t2uL6Do7X15mb6/slu7f8A9aMaJVvYi/GOyajVBUPsZznoX
DnMWKf4ETRuY9WFRUnQ2Yse721H7aJ5iC5O++FjPNroSMRqNLdsaq+OCq0TPP0JdwHxAqni6T/lp
dwk+B/cGtFReUOm0Ih2jJZUGcV9vVwE+cJ/F3MqJXZLEMy9/MK0+1eZdcwlUhiYvxcJRQvAA+hbD
Eka3WEaNCifww/poqvrAGX9NkttnkMYEfVrgNNY165AIaWaP/7gWMBpOFpXDCHJ+hV1Hwx5ER0P8
+Ef+U8FGhftKKVY6NIMqukDSoNXXr1DV2zYjuWMusarWvGdXYUJ1vBq8zZ8jNdTPqwQyCCCTo1Zr
bXzXgyOnTNJkv76xj3G7HoiiSrr47LKu/vqtXuZ35jES0HO1JFph0AUYhoNwNdJdOZDaFqDyLUa/
DJWRP1wdmNpVz4zruE8WY0ScJYkWZ4KWhU25Txe/geBIlUoEY9r53WYkcxp40LkwUQCGtXxgYDjZ
aS5at//dRjiWaI6kGqL87poSG+C1aoYonUc6WwWlI5Ufzd0QzA/rbqqEm5k20Wde3yEyzk+qJuUW
32iC+ViztaUjDJ4mrbu9CcYCCxkauoQ7EVkxfxpPCWLv/rTwf/YxQ6xBPDRWslKaQPtVMI+Ow3eo
LDJPfOia3l+HV+G6fjmIjD6K7HqM+w5GUMyrSXD35VyVG6uUbyXfS2v/kx5Phd5SRDD5gSMHNlHd
pNZjSbiXf44Frm5o1YKTNADcsHDXEEOmdl2JbZmMRg4mLoBPhUbqh3kd8FRzraVgZqwT/TTmRa5R
aAxuiSsRg+7/x+ByWs5Wv2IwKJdUosfGrjsV5gM2gVYA2/0rH91t9Lv4vJ/OLuSTKvZ0H+oCY0E/
dboNVsTpaI793YfsrYhVCXtqzNbs8U+hu5M/CXaraUq/VA76mLfuuD/k2R6UvVSKGXkt0XFfHHr4
9cGRAaZ6rAikOZRw3saIQwfqbjcdy9Xfh8hOQ0JPQb/xnP3C3M3nYmXVp951YwUT2j5bI7Q0HOI8
hkMHDHrVB7PxOmAU3H0aw1EXM8AXX8GuEuLbhkBv3w4T+DDqE7/PPnv3xWb2BW/Gg+lnSCeFZtw8
6OtToeQpldEa2uPWYwNkMIHA7JFw7Qac2t/fBVf+iP4cYtw4b35rlKMX5mvBCWyNkSPKjVVt6MGj
RnCCXJ3Nwa3N3wDJOqUSRoMnA+2AiQ9cr7eNABKlacDinR+Wn1L23HhuVAf9S/GXAwBlv9rq7y4m
hRLV98Ela7ehbTiVz0qtssMnKABU+uKB22UbDW8cUV2KDDVftbmfCN7Q4OmtHoF6BRKckj4xJVpq
i7gmT4mZFWkoj3SC5HybHkVJrX4PLrMJemQuvzQIsB0l5BLHBkYORes3PjsfiusykJICUwRAgQha
uHAoLeT23aZh0A1FbTCnAjPmNwYjMtPnElQMXO6lHRtbuMWxK6NLgV8bTG1xMK2z0PYQMjwREtzj
5dPOLgfytmVAJHeEyDxns4HwxlAx50Q8n9dnRy7Q7z+7FdvGy+xSFoX6Kg/G8krVpBfsnTIWp7jN
DtvhNJuav9vI5RhDyUVMzdflMl2NBtIawJTBWcQ7ecVUdcYtI2Apg6cWTLFNnnkkzgSX3zXegtGj
D55YXL32LIsDJm7wMHJdfRCz4FiwxIf+5//5Js46vTuWU5EOCPt72JCmexMsxWerg6WbDKF+Pexz
okcrZZI/BlhM7qfLYSYITwcW09EfKnBhXZuXXRftlA057VUPRG6CAjrbsMVFLyRMt9kJMDu+0Ecb
sDA9j/FN9JZGY82sZfMl26l2x7qYS0oaPtT+l0UOtkfUEXDsXevlRNkJvrks+G8U4NSJbQhxksg2
mDGm7ca79Tm/JZ0/Z4LMP8fDvX80XStlV21tshZgekYk1ey0HfPp5EgwJoGlbWX/sV6BMNLriJwk
ODkNdgxsQyZwOPTrXlAmoCsjrt1qi4VYVfWbOjCQwcLPB7JUQIhISubOevSbViKQj4KUvnmAcxkb
akcw1sz4bvLDf9uBf91LQ2YwKERLsfX39aLgE/CUGPAsbj0Rqa3I59eWTS6yWtx2ilqJB0jzpNGV
Ixod+8fnQlPVdQpBElWEIZz92oLqFoUvQuSL6dttaXwu4ryRNP3iHBPMxnRWVA6lC/P0GPjALfbz
yoVgGv5PwsJaGmcz6oEfRS3AbzSgsoXRuSzEhOJLh4oHw+9IX3y8/OZ7eOEwSnwpVCrY2Zhl9rlQ
h9nAFfcwJxAE4+eSgvwsa8yRBBP23/sW5mak9kZaKszDVCKqjluGOOrNJQWTGSjxQig78NLJe36q
3midvTVv1apKpARElupPqD9aBtwdMN/vJ7rQh9nDriZctAZhmkvDLIsMj+27y4e8lTooMGIDR7j+
qCMbm7hLTnJoCLpmcGGRBJVlqwWYW+PAdi8feohGOKumVdUupzY2RkyeHEziPk1tPiDvvZCEVwac
J50B2Dk6UHLiJ48U5b44gXUwQ5hB+uTOz6EVqPM2DNqPZIEFlpRM0oSnVsDB6sU2SOvAZtw0SToL
VsK9SL8DAzp+gz+zBavjbFrJfGTN/iPjOn2aGFcfX8p1JeUBO0rj4WHk6ggWGXX4rFd1D9RgY2Nk
3pUdgb2tElnix8E0AQXdnwcAtJXG58WBBVPPYXF7RmTErm9m2s3Di6Kf6V+GcPyV0S0Y6vvB46xj
MYkIlTHqug2pEVsN45X3wmixKbwWGZ8ObF4MyxXb8iF9vwPMP3PX77ZfvGMxgzuWAoo12aA/OiJM
V3dv/4Rs5wb4RtC9wADVqTqDafgKJNY3DXiuwANOT66JXcH9PgNfRdLObe5oe9zYEOOpkBSYcmW4
/1+c7gMtO0nqjtHRj7i4hXjLbchvMCeYpQO1ndAE3CPnt1vZivLsOpYGcaRNbSxUEpMjwiKH6dLV
d9egI/MLoG9AfY6nJKY56t8ZLoRk8p6aReXFEYg15eeFWr/lpZ5D8fmvmraBQRxXfu9+w/AeJvBO
Qsx3pIyPQZYVsiQ59mIK+ThfmvsVc2FNLgm61h/ngz7yWeGrZMU5QK5JPVY4P/r1N0kShprjUb0u
ot6gxWw+a29Oiu9IqQPq7LJlX+hLlrUcZwWWx3eOXqe882ekLj8NchzCpq9ZBKewHjRZtCbScPln
PICW2YUqR7htaGxOsF/PVcaSwNhdusShRlzHL0ZX99xHiZSdHLFcXHY8tyOF3Z2dxMAUHOkSSBBa
vnpbUCDVFm1AZzrVvyGv993WO30zhsGdKaJpi9afkCAEDWXUm8jhPTdaeSvZQzl5GE9jtWrQkY03
a1kSxtiAwr7I2gvIKKmuESKWL6GZ2BGKCbRO5s7XUVreuVkHcXdvT01kWiCFo0q/LEH/2KE0EcRG
PbOaEkPmB+7a9aAGst4FyAamCDLictI2m7kOBqHu3SolGHrlR6FqYYCUZH1QU7bjOZ17XVawiV7v
rlFcFyw4nuCSl0bQdPPbIBy/dO1U/7eIjvmxsNUXH/YbUq5lidoEnJYNuk+cGc98JsIDeifLIbjb
CfURHA/DO00Dhd9fGEzGZe/3StJGa8+nmxES5kPtz7d+DV3w9PdBZbaTDYGjLdCUvYuP2NMyfuLe
jN8f7Yo4AIRovAbWL4PWzAkPlogtpJMg8YL2aDz80f4FLyx8y6UCKWNc9S25GSmSdPbtjPyfYiMA
njdSTem03VTeKm1erzlJgsyrqLUK+eMKodgBlrzzn2eYC+oKzjuz/RkUMwtUaaYpfuHitzMVsuuu
arSImgtz5M+x6RnHQporuYuY1+9SmTObzx+nxzs37VTmFrRKQje85QoaeaJf70hWihJW5XuniG2K
iDtnnCRrXEeMvqPjWo4THXqzPHcb3mh8pJMpY7ENZPlIm9VaBI+H4X0iBV8s/XP9+ATx5s1ngwLe
kV0BTgL9AKNQzLBURzAKnYale2Al6pWm5vziZIcaqJ/8UFTK3GJOZhBYphaEpyI0e8En2qOZeh4C
NxlOyTWQ+4N8JLfG7OzOA0fWn6NjK87IdR8X7PP3BGdMYSGGCct+9V/4HTngZ50qPgW/WnAx8aOq
rLFdJkFmTJ2r/fNbr0cPsOOHuCZGQOMGabhZw2Wu/rYNUGRrVivQXvg05TFClNFiPWiVqcBfnHZa
XTPzNC45lJDuhT7vDwSP5sqVSgSrYe4kAZt4IYfZ8N1rP2vxe4aglymBeYjG2bu4Qd8r+v2wVWo9
v9mlDrK3us1EOsPxPM3V/8U7dn8At4X2PwWJAV5fs/AyRgn/c9iMMdD0UpYkqHnjOxIt+qj3gtD8
9/2FXQQat3/3j2hvUBbWY09hcBVdQy1gxC4C3gUv83yKOYhxqYblYCpSaMFv45/JNOcfJg52bT/K
r0HTmP5sVgjvxJfgmB2Ii7dI2t3xJeRVNjL4SANAXxngHqqTQ9YcooFsb8yyRoTxPoKHWdLtAiYv
qBqOLwZn2PBooZXdGGpjmnLiMeGRfaVw41agTCTcOLHw2OaBRQKYhllzyVGloxwo/LqNYfVOnWCV
hbdRU8m+RwmPK+1wvkAG+LTuboIFuWpisZqj0XU+ZcZdz0p99boqKFBNkUsK8Surn/ps9HPmJ0c6
jtjaVTbDVoQbJMiCoQcRoBLpE7aGgJnw21D/nkedFh0HD8SYcha84jBbbBScOLXqLTS2fNH+9qna
jg6J5Xi/r/lyASS5mYRnBhEkYC9mlUAugefFcz4IO6g0cy8uI0KPiVSa8f0K4dwPR53gjuCYoy28
rBfre9Qg+sSJ6fHsDIIu3P0txmZd9/fdC3RSE93VYXwpgfZV6NqfenUBkq+uLFeKVCNjQNELKBtl
+8+7XnE1tAzs/yhYlxVwsUFdMEEg2XHXB1CMuJpYj8Xh0t6ksR+hG6/oJI0HflbWGp+GT7T4ja+o
bfdOzwUJ32TTazn52K7ZFjEkwvbzkLYIfPbXs4vJPhUelreHfzPXWaxWtWHfRGVrp/Zb3Wb2rdaR
yRdWO99Qmxsk57Mr5lFGR8HPNxlOBPgE10mbeGZ6QTJzAGxIlhOYd87bVCf+w4Ggf4xop2XP3VkW
fwjr5VXtcagrlOHMJgCQivRS5KdEaGJDQN1wcyWA/54WE5vZ2hveznNn+UQvJxicoT4DkU96KgdS
Sja/psK94jgxlTmsF1GdcxEJzswKkg6DT0NWzaVHP8RJ3AW928G8iqbaaHsb3Z6dRAWrvV0xoyw6
d3UYTHG/5QYfMhuDFYepqvJqmg22OZWDQFtt2YWZh92tqbuyggEeyP7VD9kZM1pwY8LZ7Cbk76UM
cvLHHv7dBKxHx+B7qex2dSrYKnQdM7odGeOXjVgqyHouZbQbQgHnAgeA/NSWucEf/xUzCTvBAjby
gZ/LkgInaMuiy48P4AXp0zDeCy6N3jYsJ6dV4aeECh7Yh6DeLQKSZkGR+DN06QB7puQYjP4UsAdm
O04q7QhsDXbDarFOgZuRdENtMvkwIUVOnX6SfznorSaKftuZcVK4nckCXeeX5EOC4AwPJU3l6EKm
jX9BPpluyCWPmaZXsPm5Yly5TakRSMREIwY/2G9B1fkQdTx0udulgGwYWPbyMlkC3G23NJPcAmd6
Uns9nfPZaov9/bEE/IhiJ/jONTcRzAmwFohZCKTIA3Ysx0zbYwugWKgzAVH6UDZHKHHNciAsgCH2
6VslKt8SaS2Lm+ErRUDwDtx6iZdn5eKgzJWkW0zmUs8dQM4oZ8IYkBiCB+fInYUpK3dBxiGsAlUX
WqDzJTnnTzKEnkgTgGhjvtCHiV+TP4RlJPfDA7+4bPX5OBsocfItpIX1rR/UR3ir+bP/IGFp8Zwo
65VfC4gsqnJzuvcbZdnRuDvuCVwui1qeiCApeQ7ooJV2kJHG4MNvhBll4RRVd6GZC8lNQyLO4rAJ
UhTnAcHO7PcExsVoA4UoRyo0Pvy9dCW7kO/YI0AuBYJntKDTcxjZi8F1Kpc19VXRNWZgjFH9JtXf
o5pW/C48sE3IJk89KfuqLTWYIaT4JTX1Jx6nwgbD9zs6XeGYPia/XbUd6yhhCUKMlu3JZPTtLQTa
A4HMfvThBZGN8fJFPHbBR2Ff7wkFtayUuhUoh6xYXE26Oh1vjMctsdYJTVFr/hzxVT22hLdGTwYy
goqAzd12OSa2Jh3BbPvEed/+peJPY+MhTsSpvh5CraWk11a5fJ4q2lEknJBAxeDa7LpkcgGIW5I/
nrbgGaldqvDE8Mlp+HJ1BqdMrFnQpVRBSJdlnjC5eW1NCLy/7U0ZuVgOMYS70bwolgr83qkoaZ01
h2oGvbFfG/NPH+eTJrzl327Jft9MdFJRMPiFiLMsZffcli6/jWwSWS6H2Z6oTIJLv4GslOwxmadD
rfW+X9dFv8/OaPfGrgPU9MYsW/6xfQZ4CcjK7/Kuy9LpaS/5Rz2OJe2z1nPJoCVFQjeJCA01JWPo
MIcnvTzIOuaQ7FAkrdeccbfx7XczI6xPtJoKvaAlz4EBFNx+bt+xrUab0ieqtt/veHet5XHt18p+
VMIZqHER5uDeLSMahpXsIFJdszdV09XDG+Kbr5+9SBdbSDPPGa6EMqOT2qZT9UGl2aNtoFVxiKpk
FTdr+SXPApgtiqgK9FaUEhIjvL42CNZ1JZcYk99e1vHUlOZ55YD0ug9rrs34dVF5PEBTA2ix3jFX
3FZuPXJS4QdB34gGOWesR3AUABlUoxW0k9oMrv1rtdtUQn4vg/oblKM18T6oGKaumxJ6qPHOnPp8
Utel5HGXFBqkeOSvMe2ed8zxdLfNW/wEDZke7mWd34/abKWGD7OmX3QGLzxp5O8i6xdiqdrajFhh
sMw25+mMHa78sVtp1c51UuVpR5CSiSgOj/2GjkMyanNuaKPDvFtgCMm9JFUrPjXn1UQItShWERKR
0eYCPjasgXv394o12olx6zEjglUgTmfbjT55DFgHb7u+YeyM48SGI8DWrBBgkvs9lY7GvXYoGDJi
xlLoiEOpMbDDUHRkFtVN9NoGiBRHZaK2FqHsbxpxNgkpZZlUO8XbONLNTwteIhrWp7zAzEc6kISK
DXOa5AXbC5SsLyfuzPQ/o89bu898FdohafV8Csi9wjciBRT9xdoKKQ4nmC9hRJHUTaGYz1qI9BGv
FAaLBvjFx9KglwOiGCRWYQLqA5YIDBCp/XsFAP7pNLo+CFsgGQNLQ7Gv6Akk+nBROzB0FWYVgdVI
iTvRH1zsXrR047ywj4q8fo4BtDcE+5QVtAsSRWZULvZeDtb7cEsAH19YNc3h9jHUCeNHzMg0Cspd
rQaQW0sjZ6OFzkqSbGbnsNbBsljjLf2JH+TtVJfR5XkZ+3JZYAb5chqSxKB7YmRXoH+fYyeEi++5
08OIBbfhozgtDcSXdeeiazPfXq0+tCJRu3UVSI/0sqlj0PIeyUS5JRsx/Pu9nphwiMFAWn0lOI51
zREXB/cgIWegbXas6+Xnbe+s3Mox2xkO8/iJRCEO+UNva+/dfIvT6jUYZg==
`protect end_protected
