`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
G1MA+0H0sGig4BhpdbjMmYkeAI5jBLx+u9RJ0bHuSk+g6wMzKa+4c1MglVGpeiVOSwonIf9XKN1Z
Z82xiggcRSiPvPDZaNJrB/VnNHfCi/yt23r0qp9UcvRf/aeNGBd2UV8JZ99k+QumnirZyifICh2s
L9QNFrhg/BAA8zxpepsOe726b7FPmfD2Bbje3aJSXaerFQCDdQkicmtp1tN4PVkZ16DmVZU277yq
+wajkUS78MiWlNqvrl9UME0F0SWxkxLOj1rS0z7jsmq41PIz6w9ofM992sLbeNpez29ka4j7CJ1J
fliHh+XYZkwAc7ksHPZzolrALQcUFtGQLPQ58w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="loLbXYRj+Idia56SVq30VOejYU8jDM9spt/28fpAKlY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11872)
`protect data_block
4FD5Qa05COI3YtX4mQXF0kiicsJqjvmXXjB3aaPitc4lHtyBjO0zEIM2w55DJQPwl2W16OzZ2Y+0
Qi/RnnvirxSGpHsybQ1f1o0GnjTS22mtJzP8e+Q3WaUvBLN7sAfEz6Ejqh2wdwfpkcrO6w7NLkAK
H1RxjRl6uRBOxkXHYDTrJQT+lUc2wqjT8jhrSJ4hBQufjib13FVK1pTEfhKx2CoyVKrPN7931Si/
OHucGy8Mjb01HyT4sv9/jt6Qb272OieXPmaQcSJJU7VS4oPPcqRnoYSTXGOR0e4HJyAkBFxFFpps
ZrNG/VcVjZbrA85KGHbzeZcysyZwFv+rT9FViDpTPrejuZQTUfvxzE8jVlkLJJjeBLzAJ3RIYfSb
cULxeTUHkCPAWQNn3B4AapQ1ULLHcX8hgztZj9jCIPjohYNRrB3hNzPb8vOxvxEvCNm2ZsaPrTOT
7pLcu2oQQhM8jmA9UyucVSTtscraBSH9scXO570nJ9nrBbc+WaSHWxi8ZetcYMbB6cDW3gV2d3DG
ef8h4yySm7xry1KP0i/ln6fuBT0DZjBXUifEYK2C8DztN1J+EdtINbAgmRvwlGD9nc2l3aegBY5w
IRY9+81qd7ndsQIU0SfJTXhWRqHQ0rnWeVXEWVuGI025fSV2vcztjKnPQ4gOcYOjvZOS6CAk4S0N
M4TJ5a/RgeDmcjByzIDPUUK1SPxUMIKC0anwujZQVrXWobdwa9fL7/VoeRCzytluX5XdjJnOHYkO
bPbtBsirKl4YICJYDmho/X+1YL7lHO3lYTolFNvnFeJAMoCyFRXZRdz90XtNBd+mVNS4kqp9niFk
cYDGjSbXby9b1lV4ueqmj9kI3mcRph1vEUE+BPtkH8+A4EGrCnxh+fvJGS6/gndCGsQoOFhBw9zd
/2WS3qLfL6gXe4EEQK+CuFH0mTWvKzwQV7v3rOTF2Z8rqxtr3qkzm9WL0ySwfYDFCR5Q17gKj2Tj
nl502de6YqlioV1tOev8bwZrgjMFppD/br+W0bUr8dUTed9k/l9fcDxErVyvikkT+YeBTuI8bZml
60hU8y2CMLrcpIIvkeGPxs00vC33JCdFce+ivHE8UWprpYxizq6RB1Iv6IDgmOsQzzjVEVsMMmlm
dv9WzvfVKxAApBYlvPIr9GJDE/t0UYesIknfkdoOJRThDgToWT9X7/LruPzeZfkUcWr9FfQw1ukh
kb2FbWQiDGPa782RaRdiXHlCKmPEk4QGYOVtyCpVEteYFeYUYlb2F5hrgUIl1TbSGvlPbEHXzYrJ
aUKgbR4iY+3BoA7WNpVIk6t35c7mz90q/5bdYM5Jrt7tLDX+RLP/Q5J/dRuSl99jj/ZRXROvu05k
eK0xCQ+KDowpDvxbKP6e7/QZTwlar6ZrT4gLkK7/reLTtZFqKUBjd+DG5EBQWUu1kz6nvjpRXVeW
54omyKY2cesTonACrbQ9AexRvQnYva6OZ45JaFNeDd6xcfq/wXCX4c0oZTdpn+qbZS5z8Ffoi4yf
6/CTX76pFRam5m2zY6DDr6EPL/IQv8bR+/HXHnC2Q+1INyDWVQrWoE1N163Mwvg/52mvYNmRsMLD
u9rgOVeK1aXzH94PAnZlvvifvjx2QmqISq2wVwdKtCbQiQa6Z7+8H+Y3yta+y7Cytq40oxiD0a4B
YD+pB4xaD3p0vGitw5TMR7MATiKwItJwsqG//I25/zMU1mDU5tl8Cyih6vABhw6N4HBJHWi6C0Ha
Tq1WDN6Zbub8jnravQR/YLwnW9WB2Rn1jxHPfhUs9mFdqKWI5o79SXLUa/WO6MiujX1JlcXmKj+B
inP9KIy0ulgukizJpOewapB6UCqNImx2yvwTTChyyNxNQuhF45ArK8QbAUwbyawsFh3sWWzbc0ZB
0uPJaDh45zcBlV3ES1+NTqOu2vEwYKBD1+4UwKDwDPOG/EZp/2iManJz/hMggrqDn4bgjk9OxWzx
1UomRci152A4LpJQGwUM2HKIY+v17R+RAqpaMFOFD4XT1u82FOEne2gnR3IpogLgMKY9QOJ6N89l
HN3kQI1HRTS5dqR4nDWKGJa5aFkXYZSqMrg9aE3CqUcAmdljX9OOXXqHaeAxZaNhdvXpJPF95GnO
sBln0aXr6mtXB9XXqm5P49jrvr+4QSB6gXGdiZiI9JGFaQ2EIv4xQ3AsvkjWJXPr/lERiwHIyrVp
NWwcfs3LLtQiJpA8xeNrNNDVnvcHu4TN2a38DwKnfRLfPfufA6ywF64naEujg0txmrN81wU1I8Ag
708M06h77BJc7M8vf/OwzuHbyDBQRrNJM71m+JLngoZfoYf/Yrq1V8wVG1zZ5AluyD+QIKOiOksK
TjoSwNt6pKxEtbqL2f+B7VSMdlSP7RjWX/Z4DbLxIi69rkdkHMbxDdB9Sq0WAgb+Je+yjcRrgpmU
ZrVthIcrwYPPQ++EYSKiFg+6Fens5xpjkQDdluRfqBpnc248gss+kxEAoEtyhAEPWgdguEWWFZfJ
LSrk1XbUEF0CT9nSFxnPOQRN92c0dJMIMLL1+J/Omo/+/2KVkc6RcGxFQQXHGUfIMfK5KCsEOT5f
rWk0HUfYsDjldjd9EKvF1LOhgRwr7lZ9/UOAw5pONhl9NRIF9E52r2vh5ho8z5SUdXVLu0g8uAwI
uFxh5ol6WTX5rPMLW6uQvy8si+RVGOG3aoxbhk2dilfrSnq1OFFmSkfYzHXXnSunql3sTEB0rlpu
cWUW1pwgXSkXh1MtBdujH4CQVZpPqQ1Srwh0Dz+p+RgybBb7xc5/llbglIV/4ZM77lsWtf5qZBK/
Nr8MbzjUgPNx4FFyT9Xx/wjUiIuzFhdmXws8E6elu6jKG1drx20qg+BFgiwZ1SrzUJ3MlU1Bo1La
FYRRvVREXL2GCtHSaVZzYgxJESIqQcXxZ8Cg0EMDYvWXhzfg6NQhRZEgsa6kuLv2gVaQgb2NJVv9
WmCq1ziDvuWUbQmMWazHCXAyMLR7G1LjGAH+tgbj1B6ty2NyO00mb7fwrSjz4cHg6ovpx/RzmEzn
VBzGvwkj67abSMePgmWMM10Da46Kwqq/gbl+EyRE80mhp2TOk6HB7M6kv8Eyq98K5eg5t6hegpvr
ojiK4+N4Cs3HOOMgX6kafJ2au5ff0zwmRa6X2Oa7//4mOJGSRpvsRllbD8MXJb/3DtfkyxVmURh9
oRwOeRi8+uycFcdrzpDQz+1GwhegUsFPAs8ku4NdhZVvFxw/F5PTdJcmHl/13YdT/xploxFr9lvC
LFf/2AYuwhQg0JOMbCuXO86K4foDbTJ4ElLHFEIB1qbFiqhdL5Oa8zc4KuuTyf2GabiNk65EESHr
OD8uv3VM2saTqKmtLIb9vglx2233/l4l8opHz/cCABlnwoz2vKh25HTBxfmXPYyQqFIR79CyMZlD
nJjWlGrhuSYtSzQO4Ox+S3u+g0udvCAmpi+QRf5VBmdbPJgghlGvRv55H/VvtLVN6yIxKM/XZzfQ
fjZMR2wBPGD/aFBWc1sCYWeou/fo4ohnXboXssjddUJ69pVKT08/tExi4AW9kWYqUtXANQvhf2mF
ELdK/QFpou5YQeSRKigA2lqp/cDl9jwMskt+cAepmkFcE//fmGR0MLTMeef8WF87nMlr2LNo3Xag
hIZ0tOGNIuOe0cp0/rvq99gpJlAMxPSOOv1cd1PDwjnbI+oef0Xtesoh7LEvZHD2hRNlTos2Ef4I
fbyESsGa0/oA//nZnCBLE5eM2fqYVUsJaAALXG9vOakB3vSNZ7psJpaFvx1ORU0sLHGkh+iT7VvV
KSsyrs4MRloo0G7VlhW5Nof+7qv6iD37oJclFNJl33bbdEWsQoP5p3JQ2dix43uqb7ClLr7Yxfgk
aEmhoI4uJdb3ThBRtpkZ90yCwKWH1nJyxMdtH6mTHC7N62X0Uf+Mbj4SNLVUidMUqKFeY/Xj4/nT
OvS0xa5fENrZoJqmyDt+fJgN106jvlh+d/+VXCa0wFVS8NUNFNwFrrMD5kaDlR9ZPHr8V/CvCE7J
qz2HRols7x6DLvFmUusoTNTy+1N+4Z2lwzUH8w5IYzyd1IhARGHpTIsix7iWYP5C8c88wo6PORp1
TqHaubysMmc6mKmA6/XMj1Q/LMEj7xQoW5ZoSs2Qlfgb8dgQVLvvkoFDmEB0eDXaOxh16lgzlqpP
IVHk/YiwFROxAbl2p1TX2fyuRfcx/Y5IIbpB0BmnHBUyVV9N7cBmt3HRhOX+tYbztGjnEzF9Zadp
r+p+zMXREu4yuIk9aHppHiRKkzUDIPUGv5oSG7JFC9EOUU8fkcVE9ehRsdvi7iognBpYCKUVWiH/
lssrF0MN0glkLcc3ax6KEl3g/5TFkVCxsv5arSoxsR7FWNbCApsj098Ncn+Key1pXsF4vy9QoOuv
UcFznR27B6g4Y3fVcGYbuf6lrqi3y70RrWbOhho++5UgHKajQuW6AAKygdrvYag4YmzOtnlZACiR
ZZhNWaeWqhL/k7+ImSzRPwtfnIrfmn6mwZeC2w5XrQyga+FuOzhCcvtQoL6BYcad8WlcKdQ5xhKK
/OQLYnMu3vIY9+vVgRU+yPO/kxUW+OuF9HRM1Tpqs2JPbzBk8xPVPgVICQeQnEHeKeTMGqM2eBhb
Zgv3J2hvJ8w3Mi1MKWeIkS5hVPAmoLa3PT59kGzfBGolN2imvATyd7/rJ1rxi/czTssY+Xsj/6pc
1V8yR01rUhFhGlMjFoa+CbB6+1smhfrQ7QUmF2E4Q4JG2qWM4HNY3MpVDDkREAggdzlwgrGP2i+j
F2jdxRVq+xAqO8MTeWv3a807DaQuwKfufAGrTdjRk7VpCK7LgCBj7PdtcoPjieRivH9d8QBuFh9I
imguaMXMEaVgvz/0KGJBp80uMKJaxr5W/qXrzpd0j0GfRBb9l+aIoMLsnReKd7ooXaOfLLvq6q37
fTmgLW8OGC3LksD5EHSxeQBIzcjB23Vx3+jwMthnmmmgj1pXBUC1AcKfPFDqIWqQ0L0XuN9wYZuO
JDc8RwavjZUYnSCAY3R+KfRnM0YJy5yX0nI1OC1u9jb8c1rCgb3l4Y4LWU1jPf5zRyMevCKZpRjD
1t9klWort4BkE7mWm0iQO0X8STRfQcJqPfvPBDYP9sV5nEQyxVYRbWfszdDzQZKq7nDMVbo5Fymt
NfIYBUtuQxYFTeOYGKJeKatAvZxtRJhRf98HzTvttn0fo122ThOkMWL+w583H0cKL5zeEqGTUe4x
cp7v4P3xPcCKdULD71XNf8XiEO/wxpQp7ojNw1H/7BttyHUKRLTZmUb7PHRauFLchOlepZurDyjs
+u+JVE4Er8iHjzMFEqj98Xyd23K0uQ516WvsmbxIgoWgBHq7Ww8ac/hutfL0q+78YA3v5boOGqVz
dm0AFnQ8xjUb8eTmudcwSPMJrUwU+oxknigYupJ9rQ0S1iByK3wALQhDMiIAfizHe3rV8JuRQpWa
RcoR6B4uaDEmEtx5t2Nn9Vlm3RXnXOw2R7VlOxfbNTETSqeAOv2mKXLkjJjsWBa5fmaJbQnOB0J9
WUlcpwujYEqx5Dj7+boBczFDFCvJfCJSX5DAeuCmdu5U+JV2M84XGmnU+g2XbBzk7z3lesKNqhQv
NAuTNsblxcAy8IlhZLva1oZcfIgMwtUkFcLyT9kalCBnYUHxLY8gk6EbdMXjRVP18wJNJKf55+Be
CaSH/nzbCzY/WhO+Bo/f9l0FzQ5dHCi5Om9uS39M85wLtvvsaG04tcqtBxzz1Q15nHuOBPwpGvRw
ZPm/KjsTQ1Y+l0D+v84shUC9/Ip7Zy0Iu1HX8Xz13OYlvBipz3XRD1K9fsnXxvExhb6NRbFxdJFX
1GB7zzRsZf5sfUO4Nk/qRI45n046SIUQgaUPBnllPYjfVM74M1E3mRaIhx6VE+f5sO7ZEPd2BT+3
QoDfS1E1IRdvM8r0pMpivnEEKlg9gcxt8wJ1TRwAbOr8/8J399BMOBh1GGDKhLjWngb3qR7FHcYM
BcFkE967DUi6Wmq8faJHTCPUE/CSk8G64ZuipulhSKDBUGpMDflOnV9tdVFbZx0D52EOZIGbE6xU
Ar4TbxYPfe1Rzvl1JdoyDDaCRYQJyF9rU7sdKPKhJGoPnNuUiQRiWIggPfyzrl4/bRUwlYmkP37A
j58uyzS3VPTbXzNi0/5Ifl/NipOL5M4a0yptYNGAxPg0YObWEe2y5r/XVn4qUWqclRtjSbhzENbh
bWJWbKBxV9rzAEALSccHbgIErA5JqqwU/BG0C+h2MIH33e8gzHEvG608MrEZpWN0Jogt0J4BskBM
szsWZsbkIgiOfZCtb2poZp5jkzgUMEnZ9Exn4QAEEI+uqvpLa4rRxNN88rrkvCnjgfd867xh59pQ
xS+SFAgJWVu1wiXIF6ltmoTyrsKcYokuzro7PE6V1ck9F00Q8Li/98bP35UT5eELkFfdhevG7JhO
/60O0Zi1i9BxVXywdyhqllUJVGsIkYSMFiFtXLh41Im/W8LAD4Ksp0Pme08JEpTs4fZF56Q96LtW
a5l2gRj+y0v0akJ7M3TRFgdRFIt4vJ4C8qNNdFEOFmnTtoWY0RNQprJ9/Onc9hoK2hFuJnR0r7eG
nTdXll1M9Xr+5GPsUkBv3yuvcqxcteh8Wev09jPZCzJvEl9DcCLqRkV69iDFDXTaDy5gDbaVl9wu
pFpwr/jchcPkob4RHht2uWDvi6FbY6hTTaBBsqidAQnK8QU3E6A36xAhZwEtvzudkAo71bUDumC0
tvpmOiCK0ipeuHbHykcXtjJCT89hgRbwDNYp7zSenDPZDa8TESi6rahg5tG/dWgSxm2agt14PJbL
fd7bMop/BsdsedqPlbFFVTYebTgUBAggGJlyO5goxj3qNvvrAgnTGLEm2O26+KUc4TCAatbK20QC
c5OfWbeMc8xGW1xtfhRgX7E4p5+Sfzw+9bI4k8XQEsM9lv7U2ECtkqVAKMeIvi3BBxdBhwL9J+w8
P9xBG8Tv3Joc0skN9UYvuZ6q5HrN8ConiEsLMumwD37QsShZJvPc41dnPDA9KpGVebBEXMMeV53B
ra+cCQbrfp+yCotrKbX6dL7m3Km2jUrM6W2TTE2zA1YNDaft/Plvke6+NKPtggKbxVEncK6oWVf8
W7YeywMs5r/Hf2fVcLOEQ9kjlRtFflaQzehsfCHMUqVnjOHZ4eDFWkzXG+kzsVVcWNnoCfM0YuuN
77vm+gRtIR5keiqIEZRIUyA2EE6hWTcPaKPZKAhAQqhacqQ2bKQsLlCUa/tZ8+AlE+oz5QFQRU4x
Q9XPDSg81E8IMKwFUlEhXyiS9vEkYpbaLgNrmIc3VUe7T/DkHSEZRRrC8AbyJ3xblxdS47dyQjED
kggjEeQJA9G8cq25oHpowRMxc1aU/xz79RAYPci1OFpuBqSVVgLW3CWvo/Ubii3/ypQ060hIdJZ6
nOKtbyGPH3xhHj4sHwmdWWi1idwYBngsF/4F6Rm//K9tuaaXllpmNnt3Tzdg/LuTq631/cfX6eKH
J9On90m/RaUo4nERFAK++as7DPbY9jDRb58TPGAo+SNrcc2b+mZ9L+mDjiahuBLEVB0LoEzZYunP
qEHk6sbRHybcCPJH2BXzy+bzYzx8Y7J/m1maOpiVzICa8AbiAlF3mTbFVNN3gC4Rhq81dSrRsHAp
2hYefMVSh9D3Q/FgmAWmtbz/EToZn12JCbb9VL119nX+6qQsKo8ptRRxrIHIT2OumGV/ogBhf0tX
2aPntePy0dnE28KMNhR4vcedY3HWKeBZtpBYmgB9fOWrVZJA83jh/Gwppxk49AShRrrtBw73txOZ
X8pCWHitGTiXYZc3baxkndIbYhP8dCi2qebqyCWSHTTggiyGdaVZ+Sslcp7F8hIS+kktmxFlKN1j
GL9bOzg8JpR0CLtpJZjgPGjLhSt00B0kjY1hRjCYNOiTgbRee54lcFLdDzucOgSi5AB+/+N1e/jL
UfbB1+QWAyp+Vb6X15onG5YCZwtbnj4JM0wIaJWdPCrHww9zYssp8qMuYJumxbOlCRClGoai2DlV
f5Zz8NTezSuSwIuy0FszOnxSXIa3ifkkaPyeY+fmtlW2VIZLT/jtX8w7MSEGb7Ne1xehugLz4yf/
R3VzKCKMUGhjvSpMb1xeqLCmj/RsvHIrg95B+p90WZZOQo9LYA/Oy4Flq07ndTfsPJz5FSMEVs0n
QOPTX+DuSF9S/FF8UYtbkGNKCwNZ37P3s7v8rj71FvbNCtE4xCK7bV8o1NFiK8yDDYAvQeULqAXA
WVZoS/k5WiQrO11+vwLZ1mYoQUjs9ksljB8rRAPUtRYAtTNSn8NKnB8pgT8SeCFeZG5mni+OPRax
vxLCCq6wYJbXy4hDUsTI8Z/x/sfm0HHCYOYMCAhVzTpSEwediX9c3DxNP7iSaIHFiTv9sTjQoheq
r2GKXv9IsOI4wH6KIC8Srog9wN/43re0GE8P5BMKWH+xvBmB+7zo+uWzWFtCWJowFpTUNL4jYo1a
8xgPTN8BO2AlZexo+J3oeyDTUJAoHAsaLb1616ZSjUXES8byxmw1cq8hjOrLZHh21TfSxp+2NWBk
TGmnKweRuKX2rnC0V2DEfpI30y7Fao5J1DoGNFLuQ6o81P1EGnmCwfPAqgamNX/FDKwtE1Hy8Hnu
2U0Gj8QJRQt0SkkhMv44aFgLuiZK1M7QaFguKJWw5idU224yKjmgPCwtQTwAS2+7nyy5k/QlD4DL
Kr4wRMWIGBwaluCzMp4sL75khViv63w5FUgQswMjZo9WPww0ocXOLqqHaMRmbGrlrYIdJM2UdjiE
CH5r0pI+S45Xg1LYu/VV+r+HaOqksUnfMo+1H41VyL5TAKAA+w1+rfQc1x1y4Rr8re2VhMx1Xmtq
0XrD5ttJoZpgb4rlCuZe2VFUH76V5/dCTzUD4RCVhVHeWm6gTmNirHh0V/SRP3NhxGQaBxmCR3C/
EYOPAxQYqYVra+17EIKJ/EmvE3gQGKH5hqzw+oJYD3ZMXPqfq4Gmw4JfjT43JICtsS05Vyp9jGT/
kxqLGxODq8XqxSELYLSHLWvL0JuyxabFlZ6kXk1njq6vsX97Tu3zzOIXRE3gDE51kc0aYgJiMFiD
GHsWoZgMZlMPyVYDQyuRHMrOu9jP85yW5oxImy3Z7G8VFl+WPDoCbjTH2IImfhg5XcGz2xdWEqQ8
W74dFUuo78Sk0oOtXG78umA8jrVHxy7gX87VUGpI9hpo8sUeBnSLGo56AVtzfmuOEginyDrK1hJp
f/qA1XHLEPXdADSRjmOK1yHDOrD0uOdH8Wv6WtxHPdmXrrl8mLjwTPjj9gRnToKxMf2i+MpiS9CI
1i3HRrbdiNsbTGcK3jeF72lav+pWWme/2vf5UFJO/beNvxsiQrL6IYXpSfDNoN3N6Y7NBabFghjH
fOVIoLzObyrM86CQ1Io9jUF3FkYIHrQ1aic5qKN9/pRfzY7rtXuBccSDPTSlrNo9VFdHW4DZ7JOT
BE7D9eZyaoo6y+jNNNnCCGUl8JUOTjoK0iBIkO6+sylDMu7u9R9c+gPt4w4V1ELcx1GhO19C5rIc
kimaBoY/jPmwD4lAAXtucmpXxJkVIPB+BseS01wdRXkhVJ/sv3DwARDfCkbRjn1PhMEG0ATXOGKF
5gJRjz70pdUwS5gkeLBfWeyMWX+bh7qf6eDjLV48txcg5LwsTXuEy5f14mcBP0pu1ufqXpeY0FFh
l2AmJZUZ53HwDAqPOWgJdANrZm3QupnRxm0hmG+c/4qrFYlvzHNa/jurmLDYmZTgF6cMYWuSW3+V
eb12AS5qKC13z+AwArh49ma/VotrOkM9fnPLm4s173TxGbcLSq9ncbxLAjXHr+4nm0YGj4wv5WQ2
KLoSrO97vEcQe1LD9Xy82wStG4GEMyGOvWzUCZwMbt9fMWwtT+pDCQvX1CnpJuXhMTgn08U9aFsl
b10HFSdFB3481WR7EPRzw3J2JneN9UC1yANyUwaHZPDdJltMipVu90nri74Vut7aGNoUf6tPiUhS
qCJm02tBr6WxK3Cs+adWXKMJXD+9qK5asF5DLdaYcwPzHCmmNcmZI2tiuuKGrSlyT7vCblcF3WoJ
fza1Ium6LAlHLqafgZQeVdbDzl/laZIHWjLmcCYH2hNPYGenuCAII1Xaj2wujSRYkJK77PJ4V6Eh
aLU7fL384VY7TwaNJ2CqK+iTvBGWUvPo2XeiN4LAot0PeIY8VcbuU7YH7/ga4GGWX3VSBGYdykR+
U6I4QNR4rBddqc1eUKnUHOtPtrSHNyTqMx8JSIZn7F+eRB7e8UULwCj8lcC8ZVmsUXDH7HI2BW0T
60NWso2Z7wxoSHLrvKMX+UDF2qxuUvKz+1KIgzwyhCwQpBQPFgx/ArgTChTyReu5Bvdh3mfXdEc+
ufDz8D+oZ6XBxvr7pPl5oHlrFWck4eWvKXdm9EGk4BUOvLio8VbKkPckU3TI0KO4axbO4HjFf2pt
xGYtxQ5l39XGSLtit6fkrD9UBkYGZWdCPRCBov8JjY1zBV+qJoyuNqPLW2V/yiAuYPo0kTdhw9Rs
8ZM0YIJ2Fg+AQC38YuUeaV/lz9HUdlaLMA3BOhLrnnofxEOhVNIpULh/tEh6My0nxaH36M5IWViL
S9pN76+rVxXUfxQu41TDZhBkPdP4dSDCqTiWUY10HuvAjDrYI1bdEakRwTm8bHN2u4dBknyxeJgb
jG0DIw+0aBHh4E/IKgD95qLHX7GBCNLni5IvwcwIeCMm3FuNjaXCwHAod+CMt2Cwq2j/97+cBJwk
vb0GTwP2QCHlsnLXIBHx4zDdRR4US5iSXbCToHo5wx4z+deo/t9icy6yNTm2SPOE3vg60MBA5njX
nb/HdVyCRInnD4a7azD5nfdMyq1glrmy1Z7DehvZvDGlpFdn3nGr/3jVPvalY4CXB31LAcQzhO0X
qxZXRQUg7VrEZLSPNgeQcCYQ/ltbta+SsdBeSfpDlF540uG8nLh0+mxSjVSd4ZtUlKNAFbKquBuB
7MwNLjC0EOXAqtVuiMITCHbAWB8D/yzIOmgjRKFVqUuqOD+dtukGW/wtmG8dh1K5lo8B+pWYpzKb
M1FPrHZh0KIbKoDs5zSn80meq1ZplT1yoQW1/qgDrVztedlbdThYdv42WMJfW+jmWX03fbM+URbd
wEgjkl/vLhVoA/WeDNc2pK1ks6CWRlRWQx1TE9mg527rMBFMHy2hPszUtF6PTZu/A39mDCw1RKO4
kWegGvbBlDY2XAFNmUuw3pJXvImdihy3IXuNRxyB3v4L4+7XBWceg65lmZZyje492pS1d7RjaksE
zxLrL8Y8pt6CkolOxp0cg/YSM+J6VYGj48Bulkyh4ys9Q/ykreZOVfq2AD0qonQrrX9wtlQfZEix
4EB1uC92pKwK9cqep0+NYTZsRiHZHdDi3tDo7xqAXdrfTcTnaNZzK4Iklnk1BKl+uVGCY2hZQIsU
VAdTUkUUT1rW7PIQ4iLzndErXQ08vuX31bPKstivqM0A67y96dgEmX0BjyufedGwaSnPwtlnyMD9
WIyHrqODUdv0FisH/7N26GIIlpIEDZhC3kPWQ73PwgbHtOjgTT3Gm7h705rLMLrvkmrHSLgtD4iQ
cbbQmqdMcM4ldpJjVJ1B+Cjr1Cpe5qi5S2OAEphMKEbTsBM0V1Z34Zn8kee4EmqVMqpzl58alz7R
ZyzRLh3RyEAt0EgQn7Divxi5dormIf2mE4VKpWBxSAqXmENgSSk9+MXlNWyby1Ksp2MuVpR4cuJe
PrAhUqr2a5AArtrac/0JMpBwiHchQoXhagiXxpJUveM+U2rrzROXIWLo5sjEhrQGaL3RgvmexGGw
3xPz1UOTaqhcgKgCgMl3xGTb9bBaf4LKoSnCZIms6/4lFylkti6uAcpg08X265Hr3njKyRwBsIho
llGryM11GWS2ZjSfJ9HSCoEQHzgpBVswgDyZObelRvWxCdrwaYw+zsVWNoJNA4+p71eYHsvOV/ao
ZKDQCVO682tEO3e72inYfuOpVkG54QcssS1sQP6L018bb4MKf1t39Ks5giSPzzoDKDJaObUNAZbF
n5fVXR/nxhGIpy58L6UjCiy9rwwYTqMHv84JlWSfn5jgVdMC61kFtULeog0c+Quvg4OHFg/mGxUp
DV91Cz6YnzCQa8uv4dMhlH3eNyLReou79OhZj5vwokIj7RRFMtWcr49PIOCJKOI9hW9+WwpNoZcQ
MPt+uRQHF+/+LdNMa2Xn7Z1NtApBBVnRpochnNnWgp2KnSlqQzaenPMzvZRHR0F9+lJa7tXR9Oaa
q9vvlWJHZ2uzsZKkjsiYyyK5nCGNqimX/HPT4w4KPTkgKHMMg/HUkWpvsiUEob7hDC6akJEZTveM
fJN/QjfutuUX8mCIUwLb3F+cqyWb22VSJYWi0ZlEdn9O06m2JIhQ5AEuTpA3PwSze/40KdXgI9cZ
Tle6fSTIySKyiWwyOW44573iCVXUY6edlRU/RByoofwayOkjhggmPzCW5rEEA5bLALcXJMtvDlTP
YHSadFpLD+GgeMk6N6gsoe+22mYUjKkfXskCjbcYejcNcyPUBnKfsnRjeEJhi7xofYCOwKeOH/tb
MyP9C2BpMy3N6WnSKIpOPF7ojy0gg7nTescsVB6TmLfRDCLTed73QPxVBDCBLBzFPwWK0tSzpnTV
E6CdiSfDQHHbPBw2xJ4pGVP93Ka5mhn5kZQHqGAC1RzTg8C/40mQAEbINiCp9sBMe9bADkh9MYaj
LXnq0RsTKQvUuiR+fJ5ex0pVA6avrD6XTzowt/26z+nns/O969N3zygnI5+2uGBs9sXxhjXqDBjQ
XrSZBSz2Mxn5aq8T8cc5FStfEAVx3DdJuN5H0VL0wYHu4+hmyAh9ISnvOX0tyuSc0MPP+Khf7zxh
Y8N9lAZFYrmogJ1G1TpkrrRGRNYdGBwu7hWvgCbBB8aMmBWtvo51agOr0/tj1MfmOj1SyP6G4Ab6
Rxfd0cTro8yhzL8cW/8EAB2UwuA/UkuSxDUko/DsHwQc4cTE2tFcr3xiW85MEqJYJCbzdx0BxsTC
C6Pq/gNOO8Ak6toP5gbqTEaCKKZ5nP+KBDh34zQZrZGhiimgnLwuT+VKu/eZpUIG9st6jpT4M5uk
kKyw1422zrMmAncUb7knjCSezvHGTrzY9Rf8TFP7p9/8c3QUALdg+Wg89YiL6Jfukwc/LU0a1nH+
yFV0NMVuTuVacSpCRltpQufKrA7qQjUnu0N0zgSJSUtB3qk5xKvz6K9EtNaa/E2Xc0nJYM3b2WD/
pCumWvJKHU/kHPhRj+p0LSZlvPn2gLcDsPuyClbgr3CDfB7eHR7wkkmr6OiKSOs+VbtinObZ3cdg
CQjhiV2ek+tHUQUZte916sHBYJzFUzGksdSJVCx7JLzIsJODd7YhZ1baf5HvpEqhD2om7gEkMT4q
BtZAESHgJroE62dbOPB9eOKoAYlw6zI2dYAKsNYBR7Y9N/kdzf88o/64jlfhlIe57Zw5+0vDWXqM
HEUg12aXyw/2viN7ibn/F+fDL80sq551wLI+SyjUBFTxYaA58ku27nPQekbops2DoadG9Bz3qDBP
iexG11evBLf1vPmHigiSgOZQ4RguhIH/asZ7p8flah9NRHAjhtiKZCyJxPzg52ZOUdoCYjmFd7oM
+ijg+/L6HOC39xynzmcXswPqy87bh1qw190E17zN7lNEgLGOS51FI8ImoRdemarff+WUxb4YbB6A
agLgggXHPMDrFkykMywNQbZ12an1qwjgReRTC96CVaJ/wFiXgQS3QHK1iTM9XsyuSbI9z14JnWSV
kJG7nOmmuZCWUcUZvM/cXkGOsi93itGSfjEgYrPMXztab9aOYPIzSElnREfgKCzbTzGv/mHN0spc
rDkYdpTbsC2iZlVmMjMhpwh/mKO7FV0Wb/Ox3aZVJdNLlGriUsSnkKz0LNnlrqfKbjMxtzNy/pBZ
eXzq0y0zkzcX2ZFMjeLvTihEGX0snT3PNsDVZwknxu/a+YAhIiAsc02bQ5i8WI8/fS6J9guQBPHV
+2g25YRgC00HHuPAECpZx4FyUAOYnq+Qmccgyv9zx5S/WNsbiz0h9RJ4lrXrjY7+tp/R4y9OCXEJ
WYSwZ2FPsbb81mWR0HzKiOany19J7Hs9KJrUkgV2M3EleHuWQMyxmjygT4+DkVPhpMpjezUbBFSs
aRur6JPVL/x2CeBZ78WSDR7Eyh6GSiWouFRH+I1WmsM3zTUfU1mYQ+HL3y7+XqhQOryPbQwj21WR
MS95pjG+OcT1Nhk01pMwNR02F0yvHXzCFdlC1nrryBC/kvZOPUGzHjLJWAlakAmTNU/r4zmHcmwa
jdA1icNAy3ht/rTcR4pVHpdMx8U6uazWfQn3V/pyFHguJmID4GSFuqxdiV8bC85CJR45J7d3yS0f
jzRD08cWNp8t918MEbfBSFmPWHziq20RY8SG1L1FCQ2rS2BEX27Lai4vA08KUvaL1YvKLMOAlwqQ
0dCrnsGsBChRC+X3hbVcG7fWTVbC78XBTo7BHmJWzBNxBH6SvktvokpQZbBaad8uQM2N6H9SGuon
df9YR0r6a/4L58a6wtrKC5b+4HKgbKolBch3sgDge3l5jOCXO4TfIEgNxAUJLI1HPEglU5pRGvpF
zna3mY2z0Iyn3xTgY98EozrEdHfpRYTn/NQgVm/BWqR93F79YPYQVdUatLTZZpXi22GD57pJQ7vf
M1+HUXvdk8mc0IQf1ALXG6APWnMz1RkOtFgbwSBQbARPFzbsU+pIHrDVSsuOe7zJoSpzWf1c3yeH
QALtmJ2RY8QpSsbMfhPPbrH0w10CuBX/R1HJu2JYUZPuEBoCMKnssnYvl3WnP4JMnLDKWHY7Ez2w
DMJ1+ob3QWwcEKbNKLozFiccD4Wf2RosGKGLMrGeJtb655MRGFD6zHjcrodW5+K/Mx3YmhHFgz+O
YL5dh/xVR0FtDzNeP7NNiBGJWaRPf6w9QHMDdfzy1i9jGkkt7y3KfnwImtJvXSF+rwsqdY6RGnSh
vVRILv3+BYnNFyeqXAtqwPFfygUy1Qopfp0tpTmqsUalR4UZo3NcRm0/ZcjD28YtxJFYC0l8ioHZ
kqvHqE5vdS44/cNsXTaKM03yCVmVd8eNbVAgxwWdgmHlFawi8kZu6p7Cgryp/cmzEaIPioIn4sVR
qp5hntR4k9reP2rQkk3Sck4YLriRCy55w1J2lmAzSr/Vr3P+uXTyGx6K6c5ZQen6HIV2SyXVzYCO
6kpGq9PbpZcrI8CGotXVRCW8ujzLZm/Vr59rKy5wjOCMIrvMe7T6jNJMxlxMGHt0ClgO6wR4VUbq
utnCPCtPg9RmXljFRrXp7mTxSgQjuhgKegyoN0KDT3le9zvxxyAHKDgbPb4gi9DCeESOFfsL6Uy1
mZzj+zqXXh6w2DQdKc8nkhY7nPx9+S2/z7g8IbTrHWM03Hy06ZEGrhU5hktG4b7lnELtamon+UEp
oiQFV3iN+ivoEx0QXhXsoNCzMUuyr2a2c18DJP7XsHNCQxEK6H+RTWDkImxQ5yMK3Q/LQ4upUsf3
OHUAtdRcsj4jGDlw7eEWdDKaAGpY7jEwSX3CPkse8OMTxj8ETLAFVSpmpQvApxCYpSKIqO7aDqWC
w/9WMTRAFOdITxk42pgJDxlGkeaZY8wU6DhnLEuc0UmqOpGoSJjVvp9XKAO3E9NKvLNkTJ9Wbbut
KaMffoyL3JXgpoN0gcNu8L8kMVBfTjglS44ne/uQbLasl2PC7JVYqVczgTyFdtGBMo61eRDi+OIs
3RypVgUDBKYM1D+3BkFm6g==
`protect end_protected
