`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
OAjEVo8kw1YfrVvyomRiSpMnHnLcpW/CVMiFuh1fm4NDA11d769zkjPBw2VKVwekMDeYyrLByERn
kRSWYkfhlWheOC7fQfg7B3/8it000PitcR/uMD1HhdbK+5WRRg+wFE4/r5nVNlvvx8RcdjP5CTi5
yVfV/E+UDuVKRgGs11R/XPXD/M5eh7E3YHfrs5Fsl0aRcG7tsPgbDh18oyHKl1sdVy8+rFoZyrKE
6evpEql0cIRX1s8343n0+5d/Ja/M8uUJgEVYRLVUp2f08X7vogrLaAqX3IirJkZE2a8eY3zlByXG
vh2QxuYck0WJlfmrqGpTs49vVWFVYd3RqBX/bw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Kra1ZyBtKX1bFPX6oWcyOWJ7MIQAUv2MCat11TqGcqY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 70544)
`protect data_block
daSm3lRzLJ5iODRmPv+7hpP8dRmGCDaC2ZFw3qSIy15ZAHuiXnlg1GFfBQ3PLRrIwGCJ2lqUWcLE
0jR9ZXcvfPcOZcjQVrvW3S6eLOepqqYikt5/sh+eXHQSc7adZIfO6rQIrnRMWMGPl2ZqQkq+DpdA
7KRKrh30cfFZCXP4rCOjNqnWEXpQimN2cpejuxEX6NPDv0SDrqJiOthUluPIKFwEhXnvEnrG8k+R
tK/oaDMJozrTIXSfz7F5oev6tep4z3+YUS+Mj8NBInAV0uXsLl26Yr131E0s7bKPdaOKofppLF2e
gdarsy6+OCfLwZgE9Dim6LkIvinx3MzYIaLBTll6RXax//L6Vd04aeGEGia9+kDzg/xftEYuLNk4
E7pJ8XmJFL+LMUNVx89gFEzkIeapbg1RNXMGz38HYeWxBAjxpaZOFzO7HzdbCoZuinfM1kQog8Ce
6+qLiZk1vQID6rN9JM3hB1hk7nw3DhN7PKVZkWybFn6Ge/UVaQVlN4fjDcWBLKcRNjy+70N867Da
E1jHcc4EoaNepSN3lVK2YCbK9mwUejkNLLPrzFK7B+cjWciMN2+nPU3BL4eZIwk/sXXpnnNnWEAD
Y7FFfrWbLRyP1baDsyHj9iVOHhER3NXCyl6ztXzyY/F1mlsKfQ26URWUbWO1+gTuOhNUgl/4W7Zi
hmI696EB/2KRHp3JZsAlgAvDY8pumh6j0qZEl2hV88MNVOXQ46kBxjbbujIXEViiZmjkhrkofbuN
ZL6AjrrV0jrQoLn7ROidzZBdUsIXPgmx4soaPZK7g8l4+eTnAdsowST4z9h4R18JWIv8w9EOfb9p
X+tMwOkzaz9EgnmCpEY60P4X37tRMySx1AoiV9EZnQoJKdI5N4bCq5EwkfoAlOCkjTuk6xMdPaP6
IqPezl+lZW8uRNPkpMUPBbkEZnbX2wPKg80IPXRlSEaoI9Nh7jEDi2u6dRMw05E1hOkONOP5ex+Y
Nzke5HvgPEdS4K9igpEcJfPZXajtwAdLw/HXobzWtr7fz/pOy/+KPqukAu2lNopMBvhY4TIpC34U
HvOyGOM62g7RgGrMI2QVRLWBVZueJSNcWvEneAsmwgqFPGl8CpQwfOfP3C3cJXasz0C5nKMdegX5
ta5Yis9I5zHDvnQQ77c697fk4hB4qDo63AIGMfSpoB+kUNNHeOq3FLyhGKREE5C4Hz4QKV2HmLbD
DDrzpxViwrGA/UHH2niGwGWw0fDDRVXbC5QFVrVmEyq6tXwAXQVnWjsQFWvEdBPN580EcZNKbyCb
oKhNNe4V88awPXkNScEWimmX4Pwy375eH3YpNDhoB1d2DhyEc9PaiAG6Til3rCDZ4/V3dkX3DVSs
CDGr+DUFydWjXiTJXYxbTegdAfdn1OT4SNLSWSAB3abScnkFCkcop1mt8MEq8eeAhjA6e/QlUyDl
rp3Cl139eZR7pb/RscZnHdXrz4nbcyjfUkfyvhabVoWOIzbua7DU3cmdKuK6ocE9OOwDgnHElWEf
i8I1icwOOw/+2KDSgIXAZWeBN+03s3sD1MrVTFSk2EYuPNYqqXDS7exooZUYwkOzZ5DId7oOY0KK
v8TdBRqMKmUUU+haVeEhoOGDx1bwYUGUGGglHiLyxEa4b8RZ33oSsA8GqIT7i+5rVpciqAZb/UHs
99kNb+CW8y7CPWvWmJruYP3fqDtzOXRxuH7zK2uecrT2BH2A21DgJPKDc/9A4Fg+PfYWeIs9CeZn
MJqjE1h1+SszWnjR7c0IVedo9QaqAqVtUO1AlKrHDW3WgM/3VUd1AdUMKbXEVAE3d4g1kJR83u2i
S8FiPyHlhYNc9AAvZTR5njLFicu04P5i8Qk38iGtVVD1O3itiAHfvfQo2Ur5FboSofhmRF73iaCd
8GR0J9igDNUf9RQld3YWRSogdoOvgGrTXaUfjpmtgqpUJ4rBPDSzkcWJgBYd0NQ9Jmozd3Np1NCe
Tfi387KyzvzBtp0NzCzePQfSgRXn+VOJohcYS+6x9aVwGMEq38e7TJkhjqN0bYzJkixKEDFzrKG+
QLJ6jk35iJxnyDGy/w0miRHriCDZ3HOne9fGoyY7GtM/h3NB216CHkMgLVjvaUEO7Sm3xMxZNzn7
Z3e5xZKJaplVkHIx+CFq1EWlOlEkMASibATc2QcDlLwL26aBBynx5O7h2ebI50+eddB2F3gg1E2b
BaWgkT0FLMdcWtHhhcQyoFkQvuJ/qIV6THHQrJABbUDzl6NZ5yeWHth5k9pyqQOLyVRjGzxnmotd
1HgbmWOcf3/ME7FM7pHPiqyriTPRcfC/AYWCGMljH2DkEWG4tKnlvxVTmV3AgD4kwSkDiFQ5UMzd
LNq/qjg/8PeDWk2ZMWHgKtC8xZh+hGyJD6imvm3K0lj80wJfSGniQZ7VC+LtJxH5rFoIWUmppo8w
meo5oX3Fw6ZDYWamyThKShX50N4L9dtWB1tRUZBHDcI6s/MFKVFfQJGis+SIPP0KTYbxMDo9KBL6
MTfnTAHaBWUSfi1kQT0frUqVMqEQekmlEq1SJBB7/WOHyu8xkY+8oPaviKzm8uOq91EvSpryz4Yk
hqC9pDPMw0UmByEgZv58cJWlLcTcQuZGgwlOoEX9X7M02WNRXz2MBmdc/89w5INQsroKBvZMRyMs
sBO+Z1U9FgDraBU+Wcycxgsu0VaMsUkcH22EU9WdwfC5oyvyXfhzK8nVNwvkad9a4NhmxjqJb+Hd
r705rrRMDMJPaemZVpjJjxCAgw7x8vYxJ3thM2zwyOFvqJ+lpWuEegMUCEIBm5kpu2hxSsl6Fo8K
444vBF2W+QfE1yCBFXNparslhv3KFWSBbtezgak6BbHWhUdDk4rXg19Em0Lii9JDA6yd8Fecimni
7bBcpcNs+lN6rVI1b4WunUTrJ2ymvaTZHDjuvF1xFtCBaijxftNK6ddPMECPyMVdrd6No2pHKg3H
Eoqucm7Odqmb6cLKPd7BWqZiznmO+u8qZZHKhETQITP7QSOb5SfWi4K2aycNFLeui7OxXtDCcZ+c
Mm2o2UYsgwdsHwrsWibqGRL84JKvIFbyuOPXcuLhknQP5/eG1DVr86nT80W5tyd8FkCL3KeThy6S
xdvs5iVK20hYV44OwMLnQQDwfYowrgSZ3RVYTPQXuy81Ygh2Oouc21UL0+t/5ztD1LoUG6M0Bc2z
AmqW1XFe+won4Wa5hQZDAxqJ7S+fR+GQumlj5PXGW0gMizRHkQ08G9TGvmnA7stFaHbj4mmHy1T4
UT7PyB4BH/Vdod/QsIQr6YV10e2EW2YcWR7PT80GSgLd4Q2IzGr1HOKS4sCOMQIE0Zt9ZbE6nyCt
u602SJF62wS7SDhv0aiUjAREtwvmLoIufJBIY9znSLEimR1V9zPvVZOcyllS/qBcaejHrXKcVues
S5AlJOU0RYI7Sh5SowQB149kWPZOUhDoMFptK+95JAYG1FyGpsBN4ooa/muQRXP1hRkw4gd9BpmN
/VfigOo3vZsyNXr4fzIcwesJ2iaNZT5opbETIHUzZXCxAEpk2e8h3M7aspAZTyfVRBI4pucLPo35
fjkkj+XtW2kty7Rr6N7OJmHhJB7/do3Om3nviOYiPr6YtRMyZn4hPlBU+jGm7547YsDlPAxBJGQP
NESgDmbXLM6Bnb+f/BIjNypDw/rdSOEGrcJZ0NVT9igXk7T1GLTTjnm1+DsqIdIgpEvO/wWl4nNO
mrD4YY0Jf7ZW5o8gfLADHKfRCWYBgtCf+gYrV0B6hhJsFM/JCmYt6ViAhHajFmWTWRby5VMUz63J
UQZG2YaSCMGGhA2eb35CqERJFJcDVxM3p7Cwm5mcAzKYYfm6GLIYjDwd6M19dtMHpMcnVyHnTYR9
8p5ucuoJQOhiJ7xGP4ncusi6wPFbEgZcEFucM8jiPyJ+u0XIlv5S91KlDNHXAQZsCAcyuWWGeuR8
9vzxnUQ+YAjCStL3MRN15OW9VkmqtxocoDTRKBBeJpaB+RjGZ0fQ57W3OhquZqQZEN7NRCnyeNBU
HfdlmCrhy5mZlXPo3hNWbFN3LuBPUbUDELq8yRVC88oh8IUWer0pyL3kZadDDZ+/IhtGMdd/mniC
pykO+XNN+cr1WC7z28X5uKUlseswTXfC6jkWrL5Pb44kI0L3b/BxQBY//ZDN9FXaPyJ96XwBmxNY
Wh6IjHp9HvfUm1mipavdhmbmuyPDJgdkcCm6DIBxBisfeNT7nVVMFxw5D2wWT8YwvYuduTLcFf9M
Wxjfd1b9XyamBHK9AXz7+hrU3Nhd0CmC/otjbZB5skZzPiPq99nPKYya6bzC2yDBB2X56EnkgBxi
WwK207nddY+s8XUhH7yDYjREcUEKe04BC1Uq6uDPP4u2PkJJc/kOkMBX3Jitdn6f/rjeVSaIn83j
MWFjZ97K7UeXfNmFx47KgJPrQ8v4Bst2KNRxZcuYNiPIod4ws93kS0XlqmDbR+FIYKv+U2oVCCMV
1l0nJ9PUjA+iPty8c2EvsI9qZcjjqhm1Qy/s+64A4o8zdXxEFtYt81822ZXsdPXONcwYsLOIFkcL
y45LINJsr5kuyJjDvKFUrWSRN95DRJnwC1vZr6SOtGrxXw/ETtcjdzzh0bgOmkydupVIIBT0e/pv
xRqqgzphF00Aq1faFz25co8cyxdPGuZakU0k4Gea0N0QjQJe956DZmWnxI5/7VWoQTwDegS+YRG7
pQdLgZ1B/7xcIU1bqNUIZ5rKaRBfeIXVlnvWFtllB8MNWZ6U/AvnNdQi5LpyD2CXSjImZgsxVOLo
0n/8noZAFyHlHKD7nW+k9ajoFpY7ayvdahVMrNeDofxk0IuuQU0n5J+IH0N3pAUCjkuD4iMrlejJ
8DyQ8/fqETMsWT2iNNtZZVBzSUjWNCBSgz4F8V4o8rDFh7vbhmrk/iV7yP1qAYrfSd9655BKbok2
hdVs2tJLADXhWLDaMsnheg5AlKVwd33jQmp86MpdFDZjJ/1AsVOKW87JJyebkbmGaOkyZ2WZg71c
7cy6ZUdudHG853VEGgtglILOLS3XULb8REToQjsUDissH1IlV706VY9tgRkGJ7zsLnD/5tnNO8qr
NvzCrUaKS4Sd7CXqNzYn6PaYW627Vhf50xqvsiMnS6RtnxUAmIDZFLoUt9h0xnTl+XevCE3BMNCA
RNmyXJGKa071xuiEPpOmCJHgRU5Eb5iDJkHSiRy5sjPhSsT63gNgDdQdscNUHD1DKncVbdRm7PA9
l5BHFsndkfa/6OIdTpLFqZUtyyptOLiUX9ARZ6bHJ7INkuKNJ47nrazUP48VR+k8bWX+x34mfP2T
+bAMziiMVanngiE1aQAgZFVdkdh6OUL6Qh8nh0sEuAbvaoLCT4zf/og5UDYWK3RM59Q6xX+s44xY
um3qkJZEGmXhnfikLzU8tdg4Qd47dp0Z4Gh8606hedBOZexJCJ0KGSJiGqjsQw9aYrU+MPm6yh9w
j5BzKHZ5kE4GvrkOX8AlYizqgsTcRRPnOxKSWdjLkbFZhhklzy2fNUqAvnaoGroYGD12EEh1CqWQ
H2YpzHFvKXjID/12u99GNtt3ALETuP73znP5Wkzm0SInfctBy/O7Ffr8C0ACuuyWPy1hf+k1IsuH
01KjLO007OESdJTtCeblP2FLO6np9EmhUpoOcg1uj3TXNotU4+1ePMwJwiPlkwy+whzDGv8DiY4G
1Q8ZLqmqJ4zjn2KxfiwDS3RsT5bMGQWV58WSeKWe9w05rXNX67lcwf+7hYIZlPTqAeNaBjFsZ5x0
UtX275V7FKggbo78tq7fo8lelIOL8TnJHKihZdHnskhV98bMt3fCwiN3AmtAY+SBVNL15FXXsfSe
o6FuyIcoM/9L3QkIW7fznAMzOHLluok6JLTdc07cqO6EIWBq7obqcyri/W146tsAGXR/h0eF7OPX
ih6tae2tcPpG6YbEEqfNtUixKI7BQP3FyL2whq35m+rvN3PM/ifx1ri6dW0cau8ZVUZ3qO+kJ7HO
eO7EhHC6a18fpkKx2Vm2S3cNYjryXeHFvURX5OmlocSonJJkIvjZzCelRKlx39aiQNIU1+WasYzK
2klOJTUAfGIQYv4dnKlUVmrw4BnxdQx8h/mgavUX/5c2Xj6NBSXcDlY3z/gZyuVklthxsdcEDrr3
z9wbyq29EUxzxcOA/DMSd2n2zIbBmP2XIqRmxMkqDkVqcNjVebey8xjfrjedjquTE5nGl1taYnOz
rqv+itEdZm6x/H0JnvSg7ZInnOv2+UM7RG1AT5cL07w1Hplt0tG/oEkMkSK5XbQbbTv8IMQMgWXU
6BuVkSXsZjKA0DnG67eMzfpJik6NjiSXIiFnDt0TKm/bK7mxYnLve0hgu1aedpPWfrpV6RxuPWcT
VP6pVtFa0W6apD5HNz5RV1zNLia/BKFc1Fo7deJ9gSIuVT5YYKsXEXHMZg1EsL8lzbA6KaxfgjpC
7r5TGuGQ4mZ6xIbka8m4V7uIoBULBumx8JesBKMbYTZAR0/SYTmTtM2GsLtgT/T23FjHviB2ZDLG
O6RITC3yPf9Ohg5QE1U7XbE7ASiQdN8as7II1yEogFz0wB/ywrHVWTBK8Y8vyOhhL6zILxuHC1KL
u3uXojAt15+JsKAWK2MjTKSngSdGB0jh2zC02PSnJrfg8aTIc9hDCQkDaBU/vW/ZrQgZ/22vqFKg
TOaKUfoUoXyv8lFeOV5DuOJh2xWh63VX9Nbtw7KZk4MRKcZYt4U3k+AlAcQT1oal/lBhaOGmjiJ9
yx0eZUp+uDO8e5u+wt4Ord9wdB7YJe2dGyd+8AY5aBy2Nky17x0cz+noI/dVLlamjPA68GGHoyAS
NJTWAqcmJhDpa59C6C1550CweQVeBd8z+e7o9cxdDp0cG24s+vPQG2f0tdOm5oLXK7DAyUlNv9Db
zaj1wKuzNKsQyhOVRDEP/9riHsi5YgP2QqaUHVcWk8lnAMVaURzn06cpUtlfOihAkDyynwBEdcG+
z10qPP4tLFz5cto9wlK45c39iYUB8wHBp14CcrBzXg0K+CpBY4xIDEVT2IMsNP362TVQH9WjmDx6
r9UIuTcECcajEDb4DwOmBn0r7yCXOST84B/70CgRn1kOu4EE3CYBfH96n+nvJvd8TTWMkGT823N+
h0Y1YsYu6HGVlPxXq+TOIQDfFHxA7wCf47IZqbq8bhx064kgktqhzX1P9wRGY/CjRKH+JGbuIz81
xH7vmG2/kE1R/PGHS/ZlFiYQqxlCSPtiXoPZdT6h1RrqUdQ0qLpF5QYT8xYb4RfpfE09PnS9+H3q
2y7UweihtJhbM940J3pV7gUoCs/ARbk16uMaN2Xym4X8TDyBXS2BsPDwUCvT9ydupuVW/GktYQq/
qVgsH5x9RHfMHzd1+bdPICjoYpxcWEGwKUHKMcGU/0UT7zszD+GFoPa/yemcmo9iGH25dqjpe8gn
tVo9GxZdbGlmLMhcuPgY9GutccFXwV9ukeppyAf8XyyEOUgdGydmKcqTKRJyfzoFTPCv2ChdxHSW
EpTfx7aZJDaxSK0j3NkGssk2TzMrnH3VL4oC2FNg2fpIOcJpof6/zbkPy48f9p1T1dyyDa2ekJRV
2xUDyyKCPSf62+UgDPev6WRXmAAO3ulZMozI4mGVX1Nv0d9AjpDAb5JeEB+pT0Mr9FKPGgpvnU3I
9R9hSc4sXPkf1kUcx8IqCX4oiq5yhxR5v9lYYjwDN0JXSK+2HOVkH33tFIFIyeQfGsZFnRekmcPi
2mPm2V+SsQJyCue2C+wke4aZ1NR47x7CRqia0Gbp/lzfmmjJEgQxANaaIWE21LXE+Xhwv/TO2uzD
PEISc5XthHq8TjMCjJtREzhTQUImWYtwVBy5bSyXSukvLF/sn1sRlK8e50RbNEQr9DzQ5qnAxFos
VMo0qefMcMVuSCrthEO+t015n5V5zrtd11Ww5LyRuFjaT3g9MWYTmS7twDRxwvAAYyvj9t7mIkpH
tOsiK3k1U1MQKm5u9jAM5zI0VWYikj+Gt7LA79r24cm1Ykuq7inJyCo7jGtlCBVY2UpH5+UJWocU
U9fGy0FhtfZEqiGnDr/8LaeGOEQO0WMcoO89qIGFduhJMLeNdifTBmoyvdEx/fuHhwYMPCkj60ru
z9QKuK++23WOl6uy9eRGdD7iBkYZsEhVscWlMhaIfWMlPy5RUpkekWhvwvZmdjk/3sBo5mMAP1aB
H+W2DPPfE3EPczuYUFVa44LZN5hgATdN4Z+17HIzDQ36KmtVD3i4iSewVhuRQUw6GNXMMZkJ+V73
pY3eb3vcC9Xs3jyvYOGz73Xx2/IdYexbX5H4c8T+taHMUX74BT0Jweb2cUpH7gd1iPCntcPGybt2
UvjUsj8RxhFYJHA9upJJWVee4f8MW32WN3Zz7HJ5bjwKzfGyUYdy3vTuIZkhRhL/uLQKY3bJqCcg
hMcsc9w2fxsTBBqv+Em9bJ+xI7gQUIrV3JzOfNmlDdAK7PkDRBr/KrnrNwuLQ9seguqUiPXa0MQG
OqIIxlcDiokOSOPWq3zoxJ0JbbkD90CKtuaPHHk7rCmWb3kMZcVRYWjjWYA5tAvN7i3asKZzTtW1
VMZ1IFIdnyE1R5r3qvLrD2u6PUAo0TW/yZcP0hVm6Cn5/bQcQIdOUf+H/KB1Syof+aeZMRGDgwCo
E5de5q1ts+bCXxIVH4XanltxdkX2lqxISPAzvkULs9DaFgBaiu9UnjvDaEhvEF9lt+zQRcyPZwVP
Yz5TNw9xA63N8CS8WBMSQA7+mMuIefTs6aaspfn91SqJhuQR8DOoT9jfxJHYsE0LJaqTb3lr31a0
XAi0M1DEqDwVPhZ2jkfde5A8zol9Jm+0ZJBuMv6x52wj8d4GztSc+ITyPnK5wgTL9uNyD+MFOzxW
Cr6YnaE35SNYAjoXvGSANKFgecsb3LU+hAKhxJaVEW46x5Vg9HOyPJeaOMkAMLOT7Po4b8oBx4jt
p/ZszL1yI5hZmw+JF2Udmixhv1xMtSAgvX3/jZ81Fztj7zywxg5AJwYJmHfZUY4IukEIPnCtCgiY
cO9eY2/ktgWlNEuYETSmB9dZ0Bv4gU/X1VdF1NzuHSspIx4j7gtZmPz13+9SL+LRpLllQiWaduTb
zENmpwaqx3a570eN0XCaRwRpnkfF1gpf8l5HhJe2RYMQ4Dxk/EzwmV5uSC8cMZNdHiIZBFo2baUc
oJW+8oiwvmBF6/XGHGL0ZkKJG3dkaHH8u4N3dc7A+rfy1Jdry8NtEd937VugPEvm6Gahkp1V42Pc
g18aLuQZxv+J5Sd6fR0hPxD1XC+lG36H2UjhFW/e23j5tA3bditC0EG9lpz0a86qvoFTqFE2IX3s
EXBBoWvUO7N9WC53RDQGaiBd5d52KHtfVn3bQJE982ccqeMbpikeyxymRtStMxqXGhQ31drWgS+a
QO4PplvlFOB5WNkb0K0tSaO6UBFAWwEq/OzJ+LbcNbKKl0vKInZAOPrW+PUOfsL5c12sDs42qkub
/2nuPF1bo58Am4Qkleed1tbfPh35ZTy0hMQZETX4QJ4oppc9U59svOsxhUJZaakE7pGgzdy8ud7F
xmrB+nPe+8h7xgnrR+MhDkPLFzK6BkTBoRM68B1+AIYIrgUuKnDG08rxADG6+yZSsMM7ej+kYkAp
X1xLzJYGbPr47yBmdtpmp6lamtL/phy2mttU/o7tB7GEhjA19Kec6jWhOH7sBSvVCh6H7agtjUVS
T8zYz/1fvEVVvjj+n9ZanwIzW12PaWaQgJwL5tjDzEvRuBorx3GVnl1wFAY0fRZ1PHiHf7p+Mf/P
n/9a6zWv0PStpAbJbjDTcLlZuFVPmilp8ti5fZWNYcYczp20NfCuyvltX3s2xi8X3KN8edUbSlWv
HCUogOM/ItMMw81bzlXqckrJDcJFmJ7taro/13pkByPA0AdUw4nvUpKBILwMO8CLZBT8DpxRPWNK
1qVKNJstZVUIwnaPoL5mUWmoE9sVNkRXYxL6PGaau41x9PDinwNN9BvOSuJm8M+maX/S+Yof3hgg
EOBikYrVdEmBdyEHxHC3KQlVxJnFk8L5HwoibbBbKbnwKoBM4XfebncZkLRZzH+9oyyp2laramzR
styLCieGX2pAJYAMHFhvK9N4eovMsxxUF9GHJSzF4w0E9FiUF/KnFio+T0w6WeWQBBzDPvjThVg1
eOk3g3SFtJLAGOiJzOUNzu7vHZ7d1Q6tU3HG3hWhdyRuWjicbjhnXhlc+SzHNQfBDoe3INFfqwkf
uxXhlcPhbkjBJcez355Lyro+PL3bcZognYGARMNbvxp9mr45Leq5MkMmXKubu3R0j1TMFr5fDodX
wK07UdXsx/kgBUm0mMPJNOgt7Uo5wRrArzvJKqcdjtajHj/b/DKqvuKfu7DFCxvungSAGD/25QBA
aphNpMsm1TMxyKX4yVt4+WkbjxClI4J/OMVi1IkdbEhdsBlm6qKBvhbwZ0t+BZIwmxxj0jUUVkDo
KSDj0crZEDkrl2K928cd7J/Do0HIbm2dslMvO0Vj8LLW7SQmAsfMYBhm/GQhya6ydkflq3nF6i5k
2H3xwnhToNQ7LDKOiDv8s/ZeCsHy6Zs6YIJjScoXxuqpKsQurvSpUtDYjNiA35JDI0eOaWPGsKuS
mFLSsO/igc1eKCxIsqM3Ql2g1HxcsIHMw7MqAjPEHTNn+Mmy1OgXp1bLrhYkTiMHS/PaHsiOnNMg
0nSn7PIf+ZMCDS5fNs0RUTr74zBRUXeoQufTmveFDG0DuXuyKM3CX1zEadtW1udCxqWXWFU8iRLE
ONbFQ06lgbt7Vze7GyV4lD3jg52LK3qHZRSCJy06sge023CXX2C47CsSqNtjCM6mKN7WOLo0yI9O
psZ2csGPUOdT8/StDacU8Lf7bJ2hlLe45MvCHXY45GSKD4X3HH7NkxtKXgbTM+lGDrb+xDuzR7DZ
lE55d5JH5Y/l2VInR1NxTfLFPvh97DCOBB2xj10jJzkYVOqgnBJTiGTMyq9Ye7H4wSDYyskAjN4I
W+WM+I4+QJuBoPBS/URqRcgf+q/DiC6TQq4Y07pDyYZnP1wG1kwUhgFdXuV4PDStuEEBfz/UYYk2
lR1i6LBnFlJpZbNZsEpcJTsBbgkRvenzwZQYBdpBFlVQoKI5VO0hwM3leiqokJo0CGSlWbDM+o0x
t1lekBp8k8nGv9MyPKyB8UM8mihxuWRys4/vKZXszrjpQFw8+SXkSuVvrSz+ZgayeGLY2GKds4Fl
apZuaRcKtxbG9FK67dB0UuiF+QXsDEbgh3WDfi52nepWx3b1ZIr/pwiXU8YWx4xTgdCUUcc/3q/c
SnCyUVhCmholfupBMufTUd8Y6IB89e5SmlTy9ekgvNWh99K7gmzRp7XQZMmEii8/8wdSaN9LSW6z
9UbYDl5pJDKpab1WlpGSH2U+4vvo5Zc15LO9ZoatxxBixWZoymVjjYx8/Zw5hczq7iu3ku40Ad1l
jsxsmwLc5fC3MmbCVohcikzCKmHabEXsaEyU6RzISFN6PBa6RMf794FEgHzIG/ujnKWUR516JEoO
9hitxjbJ0MkB5QzXm2Dbt+qZPjMl/AJuwoXVVTIIy/sMAFZKC8bBKum/YySqDCKBVJj9e50qoDoh
V8UM3orzyC37xY8CcsqZSHYo6+sr/Im1PGfjkQ4pezKOvTsenBIkEc+q7lxv+mP90FnfplB5+j7W
VaI4Dk4qu7p00NeS4NI7MEiKtMSvNcVTT/aXKw+Ga4F8jjkWtp06ZQkRfvZmWacHbPTRf3dOTXWa
2O9Jpof0ceM8KABUPnIi+Kr7xa6/Mrdn4RUwyMkoYLxi6XQeRgEUmmjfgbb0HTxJJ5WP/9KVJkR4
hfW+ENHckmTumbnnanhjnhqPqb4IsTqNHA/cY/We/RoOXd1Ypt0LGKNBOINQA4NEyrX2bOVXa7Pb
yBpn4K6bPN6Pp7a4ac5yxUQLgW/04VPx+J2o3ZoA80q8MM5WWBtEuqoJVUxXqSnv/PG5r4bbWIlF
3QacJ+1TL+Ztk5fMXQklKLptJwfLUPMsx0eUC3Kl8h31O0TgKfflhLQZtGlQXWMiGElgeRgATo1c
nbc2wK/0AwCu5Dik8dgUCO0vnkMuMCXJLSPjfXVT68WGya0T9IXpKSEg12kdWnXb/dDuHTivHYlF
lOiD6NL8pMnOEEI21pDwgSmfhST7Fi2hcAVG9h9omxfGhWU6RCtCXrd94oqfn7EoWGX8Lsm5EjD3
83k/fKeeo155pLRQfGR0l6+I1QFMQChm7JoQcx+5b45slGmsG4WZi18co8dC+HT9AkvhFEZ+y+8t
w+rv6zy6AZ3dzztXPFQvdzBQLpVWCh/3bFVVneGkNOle8kwQDezZZi70NTt6znfBIj41H9rq0GNd
LZfEqJ0qCrUcPf+OT6U2S+YqYBc+ZY0ZS/WnMN33yWm5XQmmiMe6uPmNOBKc4B43J9hkEerD91in
pjGWeCOn4eReJ1ysQDQ65OLwM7WHw1mdlycp2R+9hBIxAO8LgWzeyFdOnCGxA7QMKWrUg515yx+G
Vvvs0ELSPr86RRMWnIBBYqNUFdiqphBO1EkzI1P/yC3tjrVve1SOvo3caFJBmzlXPramvRv1WNto
N8qY8ZndLgAND5zLBOveA5NRz3VoP5LXclPMbzVVtudRwrGs2BcPKfACkV/gfJMn3Kh8Yy0VqfQf
okMAv5+yu3wSuTvt/hTpxemsH5hlINazFAS2wAj0EYcdZMJ7xFbdsHyOTuLW1m76AcBCYVqWH9jc
3JG73j/SCKyN54rh2GaRv6pRMZZu15xD2hNqEAherGfgyyarYEtMcqbf2EWsdauBc75Wcmkssx3b
HgTyYrQ2WjxhZKDBONs+mCdWqZRFt0O8NXXNRPQ+gKWYQtDCpFefdCyEEfxNJRrE4X7FIP0lP+6o
tKAxCWdYisxx/dgPzQ45cKoh0+LIKr/hpURNeR0svdAP0WEKZnQmz4agg+JqxEJ0a5v3eYeDlkdy
8+Caqpzh/2yji+oi60NDax2ke5K5+1bA5L5qljUiPHwlfucb1SdVUz/FMc+mjXHh9ttNDhgYeAy8
BVDD7rdPDMnwtKy9dDas5CTPvgx4/oVV1uMBwry3nxftIs0CXaIgfMKuG6BnUGJ7Gkrcf+MWLech
2ZTL4aQZ7ejBiGqrVLtjBxfMToze+E2OlitMgnzNfdnIFH6mhQpPwWoF+bcAid9B9NgyVY3vQpJy
1nrS/dYk6y9iMBvRi3qoN2fvYxFy2hGCwJd9HvwRh7iTo48YwAt/vvCxlB4UtF0Q+TrKcS7FLiwC
MHQmc5v95NNHkeeMkLTINsuhxBMP3mLhfuDSSVV05S+irKrpBLX/yVXFbEZ2xomCOIbb/+fBjseQ
PRF7PMf5ec+Gtxh0JRWyB96pKNQlE2W8jpoKGPVDQuDNn6z4X2vSc4HUuhyh3iBQ0vhhbfu74goL
NimihlipazZ5uMz1usXinZ0ODKCdC5KLH+iQh7LjWoHyKw1Zcw82EPRF9UnUEXx0GuqDU7YJTV/O
kiV20xMw9cDfG06aLu4nnpiV79Z9O/R3cjZ6wZ65dASv3AJQ+PeOktWVcOA22SOMYJ+1OcR/vmZq
ZuOMUwDqckCapyxZz+o4zzombO1BeBjiyuOQ5seXbpF0Nj0WQhlOjPS4p0wkNDUJZGvAVqeP5wXO
+mTW5KfrfKOM+bVwnFvrU/t9yVNUQYoJOGlXGki2F323CDQrUUDZ6v66mLQLICYDNkD6WfXQwt6e
58sVzRDHXY2QFl4fE9AkIcAAeNoVNoj3kaTweXaL4vzc82sFRYAWGwZDb8PYm5qC4P/FYBbtPqbH
YojBlZdR6n+GTnCBcYmVi38F7ZUOQBq8+w2beTf0Tw0afRrhJA5KM9sR6fVj3SiPG0hFhNpm5PXj
UbSTQaQco93WMy07VOzs2FID3+HwpXTFL4jOBQKjg7MYPXhgpa4ZCtZZlozZggFVWBaniz22WonK
ePkwo8JiC/4wv29bQdigNHbwa8OBtz5quk9j+AbsNs7M82RdZbF4UqHnrfZH+4aq/TGpSXQstoIL
NitplZGtp6Oy2HJwTB85QQ6H8ZLMIrIApbC3KkDh58GdEq25luzgKA77NQE426KhIi+tjWRokDAG
YNqafw8yC81867Lp2DyV0A3h3bSSyLPGwL1707vA/MRC1vaQZ/MPqdUTe0eKXTpgPl7GB0iYz5Rw
SV6y5nvNCP1xdkknN0wrqAHaq6xnGazx6Ynik0ldVzA/xJ3qyLmfBv0hbuli6B9K+1VFgvpHdEMX
N3bJg+706o5HtAQCseGHz2v1H8BBZq4Uge6O987u4DJqvP9w7vfPr08RRYjVmj9gNaampz5DOOzB
QUkc5c96SF8MCOO1MHtTD8SpnqMS0gD2EoDo/DEbwM6wMfrf4Oz9miaSTKGwH9/4s8feSEe4pi1T
klomC8TYmdp3+VyqAWUOXXEP9Sq+1XRyKuQrAZHKSJCouT7yNDp5xN2NpqMmVJp7+45lyt/iyijC
YTLUc8fGMOC+BWpIUzPfZR3icxaJYP6KHVN36duxyqmVz9AbZ6Aj2oIAIXMGX17osn7xAWDip/RP
pjSyfrvwFoxta7svXyJVXTEOyip2DfzYub9SEArv3TwiQ3cc8rl4YfcjnTHONf/AnxHIzq6rmf02
d2BM+/kBcI3p1zt21dA4mPF74wunic3m4WPboJznFLFQcO0sRSzRyfb2UvFnEyaO5wYS0Gjyk+mo
qtqQoIoWS0cHh2vL+lgNC8SnqBg+JQ/dgpfUTRTvmXjJW3FBq9qe+odvFSroLK6pi6NJTAb5NKWg
sjIVv5IUcbBC5P344UZ/03bAbcmqCTHwe141sJrN5Y+xmyhDL/JSc2YAj1KU5958swAwS2iFba/I
6MX8nc62XljqHG41sxOik7oGGFtcikquxSmZrozD/qH9yYet+XzQTbNP+32Sdgszv0fLuhgtr0hV
I7hSx1baZL7Vb28oHsQnbGIu67FX2hEwg2F/mcmqUNgeWsPpYHFeM/WfFOEFlM3upIoif2k/HLdh
13KhIFiKs69yeNwJeOFvnzh4M3hidAyYcw51onxJJvkbMAtjwZD9EoXnsGF/d+ym1x6G01fDrDk+
gtnkDJd9Eg5EDvNiMl4a84bymnhZgWYWzUrNO+Pxc3bVM4lH8nTSxBjZnxONVsfbwfVODD6bOJGJ
4mSR/oMJkutQPug/Y1zcbCkn8HB2Ph0Bb4GUCOln1GSYD8DAQZJp3REBS4dXsvk6CY8sGITWZHoc
01n5Vcb42gcffkjfrKuMoB30BYRfZ2CdWkIaG+9FqS6bp1TzN1TqhBuOQiPz5OfzR2eAM8rn0Xcy
cvlJFMqMDtuKhmqfwQm1b1VTiExV++NJ+tItR6X6LyCcM8DyAfebri08eIySU3iQ3leEmhRIuAAp
moqvfTtEx9LvwC9Z/dP0lyZPvrziw/ePtaUtdsOKD/hNIm+5+9YA63lf1BSIHt/2rTZFQcqQ1yf2
97qKLqoe+Z3+90Og5LbUF3D5q/LgApH7C6MfeD/a436UpuvcQ4rlGkfmITIvFhGmFx9z/z5skLdl
xaKTPYQ0+yfhhdfvXK4IV+AiFQufpYTHgeut5CpNPVXtRMnNS4WS429UWZL8GMuNKufwfcpLZJbe
UCNo+JBXYO7Io/4ajpGhjLalmY+O6SpItZFOdl72G7Kuxr5bnFvGwNsJNc+V4XkPlNhNPKnKH7Eq
qo6IeI/zRmXJFDSqEHjqQ6BoXZqvAHiEOYrebRSgRwXKvNIdUDM7iGgdy/zE3JcAa2thRnq7kH6u
8vQlcd09SZcHTFL+zWWmJEHjpGxsPXkzF0xUF1a9VK0qCHZ1SjWXdN7xxpYaeIKZOPKzra2aET2I
VQUU6Dpj7dbmcGXj64DK32/vgvgpLFxoq4mlCSDKWpCC0SooIf1iUboUyyetPAKCU7DTedfxyW0b
hHeng7S5viSFOv0TolNsCM30c8F08n9M6JiimWV9pFb9oI6/anpnHfGBvnXuBowLSG2BQYs6EXzw
mHbW1AO3oWh6sRrGon/LDbS3zufugL/2lw3et6ajN+3QdG4KYdI3/BpPcsyS6mx0jj4jzRveh/40
R6Qn6CXVZJCT8t41LtKMY65REUb+RrjD0REJA/1Qj6Q//AqFDBXarYgAe55GuXBxlDzu/4+sUCyf
SOZW3Aag2y8QnHxJ4Ftjn6yv0cVxiR0B1sEUxs4tYyhFM2DFTeqe1yvpFvMMRGEE+Ln1s69Ni2b8
SznoFuS2PUmsgmGejDOLijUu7YuoYv6gSmN61vzMfCVYUHYlwW5mXJAhyBRWQ5FN1XLO57xE4N2A
NC+DJVtuS19s9WeDj5M0YxFP901wuUKDV9gE+1r5r06jptDhzk9cIeYN0NiyUYUxnVtsOhUmwhVV
756fu0KY2gzScbnwVZibeT9tiwIAjncPfD8z6tElmuh7BTTIEzaph4EtvcbKrLiOiQzNcGSGQ7yT
XXVaR9geBgXbq3fLnQ2REUa3ImuYC56g1sP/km248jbL4JlpqAYU/joO/8biiMa/wOXxzKKfiOqB
Kl2EgLpPULMkj9uYi2J1+sTaThQxg1wCMvrNjTSyl7RAnggbZUFmIHmmO5yr9q7iH0coPKT5luvU
aKbMBBZLTDyanX/rv18Y9rKZE7P5Wx58X0ZIHJ8Tkn9QcHyLMWUFGEJz4J1f16/H38yzprQCHdw6
WYhwXFd+vgvZHJvgqBPUUIPE4ZDyhLzTHIpfZ5i0jtWfFLxf8sjnzJOwnMyMZGly/nU6Db434KyL
BW/AtBtf1iJi+pU91mRyGRaKK0hsyJ1kZCiZvMZE2j/SvVBbvXojKl1eL9EyKRl/wlaDi8xoqWqs
/RnIoUunTbZDADxF4wSJeNiCl8uxV1W/C5fd/9gnbADcPszRnNJQL1qA7+tT4UvGCa0ydmNXSgOq
5FjpXa8vrNyojahxlLIh+we0KsfTXgOaI7rZBsMY7fom/jYMV/AptsH7/jUKHGLo03yLkyCokkKY
yr6W8S4iHqmFklxVXT/ze/o/a/ehGrplvhkpPwYNiw5UqRx1kNKigWvMM0YkQzmID5pHLzVaw6jx
bK3cyPpK0c+ZWkfsQcj6OA+G1Mp7wJeSqXXvddRRKZDIV25OiamE4Rb4ImNo8pzlUdBUBwzfxEVQ
1j/kEeZcUgHT6ikThF4lZCYBTZHSwt3QWbEUOG1if1okuy6vmWwGrbJy3O+IQoW8cGxXup4HWNPd
PyCICZsAFhSJMg9TUQemwDOXwLzybXQ+lgOkjzms2BggvBVuBWsBKpygeM6pigXFR19mWic4J/3c
u3bjB5oYRF+bADEqt5PCpHWRaNEXxkOY9RswOQdZX7JqMj2M005dOk6aDTNIm37IPCiJlVshMKHP
fR6iO3yo/15CSzoPKnkKD0dLFYXRJtXX/ToIV2xNnFzIknlNvvhacyCz87Us35LHe9am/YC4qJOw
4he5WsFef4/NQlm0/bbmzM0JAw9njsmQOCw9wP7Pjw8hDnDywhEeT0P7Xmt+QLsPz4RcbEjN9HQj
7HQwtKBNSf69flSul+34nINj2vZfQFkT0yj27IXbf48OfuutLZE7W8qp8MqijBtq+7CP61IaIEZ1
RebtDKhM7WNmD8AvAArVfiqRZTpDsWP8q3usD/ZUls2G4nqavjrFOJLTwY95V/K6vXP3TZGhDSlL
Ov+tftpYSX122sjuQZ7GUONcH+s3lC+67cM04ku8BRxh9PN9ru9HWA/mUsrICVxo2Mb7cm+lE3zk
zmXivAQTf38838xx3+1iiOhpweEXnB8vUDlc/t2DdzAYxMdcCHP1pUB6jqkZ0AvT6EAHXyFOS4F9
MBDOM8Vfk9sPCC0U2Qd8xSaf6Bc/dIk1xpJosgHSwOHHOea7FhvkCf/8koXgwkNUNfhCTs6ndxwq
i4lrEHGgGDfktOV4oRtXBq6a2BIXQealoV/sBQk5FgGxF5pAuhENhsxk3faL2IKQWCQUIcwD7sRB
r/ANbXgBxRjKTpePYsH5S746tlDrrJtpZKNAOHkQeo6J4pw2opgwK2i6zqQv/MG09ohjgjxcfbMS
igzFdsd/o/wDdX9+XYthqh6hrGbvH5SATmBYW8/t4TwhzTHcPgmt5IwJMYhm10q8gGvbBqJrra2o
0Zt3FvY5Se/3+oB1T60DE6IVQQCfNk5omsXYZWWx0uzlgWkOLVPEq0jmcgRJRb7cViyANG1Cqpa5
fziUQO9BfTqBpSgqIqE+AAPi2yDAukiOdbyECDM+cv0ixwJwV/qFwpZ027j/f+MwzH49n4Dm1Etq
icKqO9e44DjxmujP79hQ3CUK/l57UdLwd5Fp53H5PDnHsjZX3o1QCvHiyfjzMXfwSEdJGF5Dmg9x
ZoUj2qlvIj5QOIvT6bfrKAMkISJUXxybXLwS5gcC7LUQwdXi4FlTxd0vCjrw7/yiPP0VeRUGrgD9
jHDLdQriqIRun7g+yW4DWDnURA916dHXphZDooc2Iqdje+hL516OSr6/OO+cf1mKEXHKCWOMzruM
WQHkTYDCnxh3iXouKO4V4/FMZ3GgVtkyaEQR02ZKihv8ehzCTHviTVHn57LC59Ar8rd2s0oqQsek
g/5QDeQu56u+EfBkplJOrZ5i5lXkj1UM8JueP0JIN/JQAfrgl/+6zpzd3VrLstOo3Fx7XlW+2NeH
28nKVvKiLvq4l5KgV5fpdh546QIzQfC4GiQh975sRSSOeNP9p+JYJV5ZrHFxRAUhFZM0bnMVGQ+i
8CKO4ZaCuY6oXh6kupVLhrOjcFI+Pl3l/N3sP0r7O1dEMJYNjkJTLY3+MQHBnoP+RJjzuV+Wx6H0
6eM1s6eJcYjcTzqTjvbdQ/WvKWO2mMbNtg71ksX00v+8paykDKQG/I0mFgZA+sdnx5Ht+gVWSMXP
XbeLMeIAHP7kr6syi9uQpti/lUUv0uNSKkCpoXWW9OxSL7ElbphzBYOHRY7jcNYuBiqJyf9qqnYl
h/9A/qlZ8P8zqzuAFix0uCHB9kkNlOJ+eSUgdmSDmcW91mKdk+/L8mJ/qc5PwI39GO2+TVQttT7j
BmrbQoY3KxpmnHRffQDMexTx3VDHTP6as5hnX52gWAEkvopgA7dLmml5Bwt7TIw/c+0elBFtigr+
7xq4ihu/yVMUlLGooZpOv1ZbgSH0WoPUZCozh6bGqGIgJhM3FWznK5M2EI2mRW5vh+JexjgWsI+5
OX0NWHl5ORrvipmrp/DhGtxYILHhgdDZ2tNa3cZwwY6e7Bf0Ao9XL01G6AG17eL1OxuPkHhyODoc
5sgQH9l0V2TXjztPoR4Wqw8ScVaGc3XKYUGtxG50BSaQQWeE4wTt6+mLLT9Y9OVWivhrnWlQ/b5g
hrGsqjsRYdhmn03E3AlhJF2rJlLEJXT0zpTfJYMLpa9qApDwbWN0wYriHsd8rhn6YR2BcByFx+l3
Csv1PWZXCv6QQWXH2g1vQtH9KpmSsf+oWhPhuA9vihhIllOwBxrVy0Ogz0Eq/2KzlLAPbw87U35U
f/VPQUqAdQYSMzQTIUepO2N6LYdkigvm4MsJQV8Xo2ARv4TQzzLnSM1oDful/+UeKN8S2dc7AF+H
28AU21vwNLHec4cSF8iCrUQcj6oORUTV+QyGTtkg3mu+xb8aMLZsBN4RYQn8TeeV292vE4xACxzI
DCANAdd4DVnHGIu7wfaxcRJD2ztD/0/ieHMTqgzq6URkfugbGO7HyG5kdu+ad5Xm5N69ng8b+Z9q
Hzd1kJxwmjnTmTTI6Jhb5DOx0oEh3m6ATR3NeK4ZtbSCpCAe8VigufXJ6kmh/tRRptYVUtZT0sqg
GCQDZoaVIoHzI0BhX7oxYa+I46RjLiTFUMIlyhmv9auWvJt50ErhTNnBKxQGo+VBrZ4DXoTBYxjX
eyceSmLkoVkqsgSGmY4kzelR7b28nRkYEnIO6pgfztMDrJCsxBuaz0DXV9kqb47+bdi3cxMpc0DK
0rWTHpD4jiSDxK6dxWqjngJj24sHAsQdLz/uX7DGs43jnbiODScCI+O04T+6q+a6BhfJJu541G+y
/TitCwJlBvYe0x6ylxC9fEc9/6e60voVjRHhggdd8AZVgJTOEqn9QgUqVpgll5gMAWA6FCacIU/5
ZVHZAHMiBvxsFdO+BSu5v3YeAuYwn74aAwldh3cVt+cTVAf69lKzi4bNGITXnR4DbsMHMCUaudSM
NB6bFOTMd11tn7vAziqhdwaWwxpyCEftulHBcEaT8YVwXp05NSPynCbwP/3WD1dXpokdyTgyXSHv
T3XtYublT6GJjW+v1QDUAUvxcXgPjYM7VC8scrw1g6ObEghzKPa48+vyEbOQlJrmZ5D1YbpP09Oi
LLlHtXT5ToUgiS4+Yti0p6731VqQ4ENoHfNIzbiEZnav6LKEvS2BR1eD16RzQsu9cl5OKCun92/D
9iUFl8Kp70kWe4w4hW86ajiWdUMVeGPV1RMbW1IqxnbZ2miXCmtvKvmhd3+NKRBA3gGpzbRu9dVj
qaG65bARj28Ltvn1t83hPbs0WQoI9EWvdUWlr5jZFcexpw3hE0gYK3Xc7TNNwGoeIyuFBvbrgvQN
bIFuy3fQolGfwRfEqv+ozp+o7p7Ch0h1JztOWJTuk/mP4Qc7fouY9Abnu/DYZPYGOAiB2i9Q8Opa
QEpxSpafE8vzJ/LYedmJ13QrPHSC+30cAB8FxiXHMNWm22m8D36pVnRKiGqaHMFhs72c3EaU8oKO
5jOpw1g1MrlDHRMzJ9eJuIE5ZUz3UmaYz5y2KzM7l3oMoCUwiEyFWFBXlLwO2boMGiTBOfWnh3Uk
i2cp1ZsdnpeHPHk5npoq/0SYI7A0ZChFJbcSQYmToilAzMX63s6aTkjuj8AxMXi0TAHMMKGMuZ8B
GalMLUOLHlXhtrGMbFaHq46KRAIhk7i3eXVXzTWVbgZvSWwURG6O+XNvw/bUWj0S9ogWlDrH5CY0
aG146AisxydmAEJp6rTjc2yt53nMQL/mrYOnOdo6qdu15/HuhOPlIbkS0LDxF4pb/nMZ3GiFSDPz
OkLmG/Qw6zSx6zbxVdWxNH59qR+hAshO9p37cRWpraMDZYy/tW0tVg5jNtkaiTEykyzqA+mqkkrB
yO7fXHstvm9zlAYz5F5WsUwRc5Hf83MfVGoFOrfT3MNzI1oLqM76tHxKtV0B9ywmEh6g2IcPsEva
pN9iR6DzAcevf0+bkMlRRN7nhGmtS7DkH0cQemkWzKM2UopbiVu4SQeYd2NDIm6Fn4E1TpqIsEEc
otW5Txcx9rgef7ia6+CPnBkNbWfuH3g81qCBD/PcaNYNCkmodqnuCR+CtSNQrnIZwiTRGyxxe5jQ
cDuzw+7mk46YUyj/5AsYMOR2b1wIhSKq00O3w4gXyV4Jr9h1rmaQSjMgEH58YnbiSf99Q0z/Wl1Y
Z5EVeHLlBn0VYBuXpF12zvqC6LLDYy6c0ID30MuyV0EwlDU3LUQhhpOX/3drqOHuDFmUTlp9EqTb
pNUGeQnStakgKihyC6x4iE9Qi+1Hn4F/Hp8Xuse6UJ49WKA0nbpYnD8OJZaNFnWBP2Y188fGTZt/
kE2WPONK/I09WAx+KQewNSkJVKAXDaCciV8Tk7HpTWePhCHEGPEnjuDhETH3CRXKfWdxYs4/oZzv
49U2Bvr7Np4UN8olen91wDt3xZCZBfwyemORzwWFyH92fL+KwzeAR2J00gVFUKVX/xprPe2CVMdP
9f9xjDCzgVNYrEAFUr2RF/s9YryYHF+p4NCk/cBvnzCg2X4PTvX9uDT2bwPvcYmDCWQYGQ0WMHs9
+4HtJBF7kdXr/1O4jcuXu68be+1HNGk4/dWa55HbRKRRtJ6Lu0FglRk/kHOxH3RLMOMzt36qTO1L
PNKRg3EDpiKoqIoaFKIAARhuTihI8TfEnrxLYQQlmPi0S9qIM/01RQ6C+WnmXRa/qSofvT8BL5L4
aySb2bfPKZNTlAZvDkE+fooSNb5t5p0MAv2EP6/PRsscebeJqtJLtqCKEHzXor6oj4qEnyIFmtNu
3rf4hL+yhaeoQZxhD3d6uiAva2xkp0GNdiGFRxfb42mWJu2Ra2lKaUL3R+rHP5RYflKC5ZMqoNi1
iAfvVfVj403YlE1qiWJimN2ja1rh0+tCCC+S+rszguP6sg6MFNr/4Y2mCUmMeab1FXu5WIoD1PtS
DANIQb4CflzRDIoUiSdknZef3q0tQccrKrMMceK5gddFzoru6gaQgzEJK2nd1FdIXTeAmC4H9ZDG
VIjZbovCulGRSnSx1Lez426xRigUGnj2VaUmG6QsXifuXofb4Gj2TH+OyOXeaCOTG4b18uFYQD8y
s7vGpIOSWDfgl0Iowx/ZAwHNKO1Gyuz6+TtjQq4iPHX7nyI8FY7LS/XIk4a/01NvY7UFAo2sj68L
znUe48xi9PCQkkLvupDmmpDUPLl/OLfufgzNc7/xO8F5R+sdDPws/JuaZ64Xu7TF6cl/6Y9aj20w
BS3d4mv0WvaChXDbdOlq3olzzjn/mNte/Y5wz7QFQ70/HDgcK9QuULqPdV7LTrRUrI6V55sZ/Fot
0698MxJ9cWocRLQxZt7zfVhvWb27osl+j2c+WrFr0/z5mM52nkYwiv6c16UrmoiwqsmjWjwefIkd
RVEwfjoFZDfn5NnGMkNvRqoMXUvtt29xkC7OfpMFymEltMf6sLrIhLb0omvOytK9F+/tV7k5NQXf
xmzP7F3eF3CTG16kCsD4Ft3/Es49me+2QQQh00SBjEgGiadcVfaodJ4atLVgCHHeSd0JadwPoUko
v9A/3mGjDA8pSrhPIt1tW+IIdgOt/3FHIlHTIFvJRpIk+zKeUdJT21HeKu/jp593ugW8EfCDBluN
+bBaTXGAVuRLsEyKHL/I+fG9/nbWH5yrqVaKI2QPqvxNVCsCxj3b39l5Zedo8lsKmVIcT012QHzc
GGbiT3dlV6Ea35YySb6Pe1HG8Ptso0uG79CqCKcyquC0HrskSjGmf/hzdZ3YHvpdRnoKClPBQuOG
wt8vVS9n5RDbqBJ7XbAVu7BLfOjUlNZuYN239+ebfTPBIphdjj56kZCblTkMqUGZkh+/GNRcVBc8
KVispgjKgMWRPLHIcr+yFiJUjX7UWdazAvqm7G1/MB1jpFfRtRYnxXVUFH841SgzE9xOnkOj7bGU
SgF0tf8Gh/eApb1TJtKkkMXnDz1d9JTJuhQPlCWxU83iJ12fjZxWP/YMIPspNiaVMZe5+lrQZUoU
6DuKAsD0nQQylwIPgSSNnYBzvKsINJ8hqSckEhnDxmfOSXB0OsU1/mtEVnPCsalsKM5+IUm77OPx
n4gk+kyzzpOJP7sKm6caqUdOo+w/0SPpJFq8615th0NH4r6yEXO2XdJVN+v2TwQHDs4z7espxKn7
7qLfB0gr3mAWU8eivnbBobBoSFBO7VUo+z3/u2+hdngl13de8Ab8TstTBIs84u2L9VoAL3gO1es0
qkLAcjs6L6nlcxKaXuLf2LSn0Eup7F65igZ1sVC7pDfQYYZoVIbCD5ElFFnCF5R/Kys+6Y9VxQvC
Jie3abhC+KdD9g4JqAQXEzHRtuiMQvy+NJugs+xu/GJbyBhsbHrI+oszGs0BwyuYO7T/NAp8qEPx
9/M7DTbS+6Os2IxJUARBNBoLLxQmFAFiKJC289Fhrp9CcJreZkozE26D3EbUzG8Ht3xNzfZBvTaN
vucDkFTW0DlxvyCVH4SQAV1qmlHBa4BWIKLurjEUA4SFNj7H6G7Kclz4TRBgkBVE6eePAUqe9nZD
/zrfLc33TNBggGj2Qx3qUz7Eg+iIfg9ex5IkTjunQLiVHus7nSdz3YSi9e4oGX7s9J6to2sOc/7w
Y5f90rXIv/KnQUJ6VYocqotNCkxDqW5rkRDCmQcGGEVsWbtM0Dhk+pTJCguFEweUWAIzONakzDw4
rMEBzwFRoJf1Dk+hklHpRLvxkhKiKUP5My7eFdkQFzGt/jJg0iu+dK9Tg2QUGPEsycnRnUTTOteN
xKQk07cpzPYBlqYH1/pbrmqcEaM4k9A8YDGGfv7LZFkt3r3YTVOi8pg1xU0OPu5jkmu8Rz12w8YA
tg/Mo0OedVMZ6JMLHsR0Tf/jvtGW1/yd2PGds7CzJw8CHaxRhWPT3ysUZfcvDH3ZBIkVT8IUbLc5
5B0iLaUoYv4yVwk4wVnaQ/KdIzbiYGkPzQFgR1Rxe3pdnlbJhI9xiNrU6Rcr9NgYQD7DJmpik6Vn
rBpYLJSAwyyzQScaDSrUL9LExrhowG03G8t2AGZ2T5wsuZvUKyRbDxaRpotkFeXW1SICMTEkRS1h
T+jLJCEkmrsujzAw6KqwQ6vfwCelUAIehDy33QNRp092T8oKKUt4+ft7yfiudpX7B54YNxsqPxsC
0aFSfXftjtvvrrq5F9Y2USJWDv2GsVyy9hwr6CRp+qo3D01LENLkhRAtttXFoEPDhJHsiQR+pVmt
aI0EYWjgwcKZunbKlr4/UtkjsN7yWkT8Y25twYsPL86nFY06rgGPDKNKLMHHE3ralGSAHDpPU161
YPHsAgMpiV104SGAO99ZVgfs9RwZUDnqpRAdvSHT0U322KdWNQKL4khis0hlaqdd1xtJr/O27F6t
ljDcTqCqIXfjFj5RqeJyJ5pX7dGDYJCxXsoKCjUAeWj19hX9zYzYn674frJiBFaxoPh3c5PEekYL
jHS6fco7vyM422JXP/Q3PwWi2fWxFlUyQWowgbm6eeny3jmmKzpVM2jwmjSVB1AtepLLMK1Gr0Tm
9rP+tBWvBtbDD1zjDGkE6zM+XcmxpVuy7Oz0hhz8nsZ+vBOSGuiuRxM5skE0SEyN8YTavQnSGSxV
twlHs3yLP/x62j+gKIzPuKVFjYyMYoSEppieD7ehWABJ8JynbiDHfgpDUmCsWLNmCLziTeQayOJR
hG0soUoRkpfOdSY/aQ9baPkkfdIu3l9Zrf+45xnheFkAgnEbDv4Y4wQHGbDCm4uzgJ9ZPpYQenQX
SWgRjtzCZeaSIVKIeql78xZd5U9gmz6rrex2ItiQ4Mg8KxYRbM2Pvb+auR2fuGoP8/b+JEBstjDy
dlzM6FQ4ymwnaM49GUiQkNKjfpmBEOo7VXb8Nw2E9tVpVCP1DeuC24BOxr21Njaocoo8MsIGnHjQ
hQ5gwQMcSvUebqphBBmV0lN/izMARAUHWHHFSmtbUr4VXlHcV3KqN5v8xVqU/q2qUdu2M6RbnhZ+
PSvMAtdIXskoOJzWxcw5ilvli+shVdQDtCF3Fvzmq9gbDxlbkShkg3CD+LTFnLo+9aYz33/g6cFI
i9cOuOTOc0b2rKpt4ARuhlC3Jid0ZK1SfH8paePWzeSUH7oVkxC4o8jeHMD427TKsnc3q83EuHNp
DfbNwl91ixviXh4rAyTNlr5yng1g5LU7xFuiSVPliunq4ceA4C7CWbGKbFcq2uoGYM1NXaYHatvX
RkISJykQLIbFxYP5NLetfWrCXiyeZEP6iCN2AIEP6zWDaDdbvu9C8+8KhFjgrP1CzZ7CL2lQnGI9
kVgCr64b/GBvFw73TK/zCSBQsZUcAR/mFWcUtgHVGpP7mg7SKwwmLAYhO5d+R8+m4/+8C2Ke6/Bx
LhZq2KbY9TPuBTga5C3Y/NAVDlf676Z6G6kDEF7kTweHbNr5MdJkM2itb+jmvwGH/9MrOd1t/4JF
JTk8O2jCPz+gnrr9f5LFXpMQvwFHKnKNpuMPJx50lEDxdRcFVS8GoETolTXFT2dxhT4rOMxmodeB
k11lVFUeiE/q8sz1BaN2Jrm/rqlW4ZNVU0oS027ZA1QnxjX44Oe6JeohyeB4h+XBCN6k4LM6pa6d
ELdaNTRh+KQB+tgS2Wg/GJTu8XDmBufHIVeOV/nkP5+RtnzGPqY8vXWTrLZ1piSVumeVsFYNEua2
OElTX1psYPd3g6He5W1SmPYZGXpl/iLSpD1aA8oc5ARYuc1SwlsXHhihd2/YsKqZbnIabkzRic+W
EfTjD6O9d30vo1sj4AbnoT3Bt+tIrLFa5ILoRQDsOHZrLnaiYgF1WpHYClbAQzf4spxjAevvfyN5
1VBLB3R/HW+7QSQb6G+gL24PUWSb+WieQd/9p4fvczfP/SoFZUi7aJlGOob/FVCcsqbbUtAyN633
qmF1VpH5HF0wepjbdKmCz8/4BHkymJRj/+b5dWTyGadQKhGdEmvYV4Z+bp80s81wm4S0nf8uTztF
VrnTSQdnWloOZ/fS85mDdcnqcqRcGdu2EJQIKZpCEOnoc6e3xZVjCh/2oescJuCQOQBq+4v/IiBr
CqS0qcOnuMh+k57HfbJco3KW9OL35MDcOa6bUWAhHcGV57XTN7MTuR9wKDSoqS89XjaQqFKbUCzn
Gl1LYFkifPWXpKXsW9lEHU6Kia7lH2DaRIYQRcHBCF63mmSURBXSwzHtBOkrjqiAzOKnejFbJ2cF
JMoPmYYX+E0VPy7GaOyU69SNOy+vKjE0kBzkeJJLC4fonTBq2haFO8+f3JnS3BAv4OaaiVJH5IV/
RU+B2yhBofY0zvxFII7GyVJpr2+K1fvdaHeQ3g2GsRDOLRQ2eTngqpwPkoYYCP5hxLjGYdr9Hds4
2TNzQI8P4PMyc3SZcOkTWpVGeoX64DNvkLbGqK0vEEJ6ObOfqMOM5DUZZh75FkZrXxTvGijCmpOl
kdeo0wzaSsfNcSW9nMSyvyHMD59VJafl1Mv+HI3u62XEgRVa8K26sNFzH+5EVzNQIN5Hm1vf6Dut
pM0S7UXROfziJOtcN6vLT1tBMulSSeea6fmVkqgUidF1l+Gt9+sxHsgz4NijvHf3XXFfFkMy31gE
XJPwksAG1haICXazbehlNX5h1HRgtjhBmXEnaa3eYPM5Ic1GVYfL92hCMas23rxT5X0aTQWi9/fp
GmNcCOvjDCm2UoWSOqt1idpY0YDftQQ2lHgMYf1D6kwVGJ+cTVP+G3XEHhURVuzpByvKPNu8CpeF
oa1/Oakavza+36NS/iZXFeslE4Lq+q41U1xVgUyHsFnD0JIm5Xzrp8m+2TN1OVKpI2giV6ewIuHu
RHYGL8uMbO7YaNJ/WHufYlddh9LqNBGLkL+zjlRnPjN7UPR8iVK0wqeJEkkjxYU0uVezeYQu/Cgk
Bf/r1sjItCFwKZfp3/5fKPr6qsj5FV+w1Lpyin+4PPB9Ko3ES4YGwFcdRTEnh9TyfIHGMy77PRdC
Nh547lNp7kZe0RqMzdIMInyv3w7A8MTsYc20Cf84wqGzzFUvkebG0tkRSVtlFl5xZclJH8nXDHIN
+Fw1oCJkR6fg72+1HOygVmqFvcf0Ahat95uzyPOfsJtOjaFruFQMMfHYC1TK+733vGoMKAV0c/P1
LBNGl3uoL2O01rg4B4oaC+pRtAEdQ7TxpJVFkhi629o/HUM+C0zSp13hnjJpIM5Mq0wNzMS+dzTV
1tlbsWto5grVmo6I5CtwOGMBeDScPaCejvIpLdrw6G0MN7KHvpVEVAgsX2Ucx8NTZhQ0e9nWpDAK
H173zhi2BNY2+ZFnUod2i+9XJO/hz2fVngdFsPy+VVwfqHUY8QsJzOwPn1rcK1byCFiNaJf3qY/b
/DJHHdjfVb25HYJwhWLvAlgbM75wJ2ts8WRHsdvtKCyXKwOkO/iS3ch67aSJPL4Tg9PO6+0VjF0j
EgsO5ib2J9avyNvLSrXfqdRlmuipVuiS9YEEAe+YyxTmQl3FLSJ+B59hGKFFdhte4Ze7VlmN+erR
FGXWiJrx+sZvpSonxffEinEqMKWzQHM/20kfSn7TSp4AZtqK0jZjvYlAhDJ6GN2QPf5iLwpz5jsQ
XGiDx5a8j53d89JR/Fm4tY7EJyRgm2+zzbHKuHF3o7DtpmWMs/0CJClKJICMcQSkLG5rA8tf9YoW
9UjOY0bQn0YwV47hzy+dX5/mw5O7+yskJj36mdvUNpO6xw1b/o8LQSm2JYyXeD3QRMOzhpCsbbtl
rO4sC6obitrm8VDmlLVVWHzjRo/tTJJfj2+bxFl594ZvixUTI0GennlxjGRRcWFdQbVWVZrNZ18U
FRGEyc24pjVn/4jQZnS/dQvrjEXKx8tGTscotao5zH7xuoxFn6y/aaU5HhlbVDTWz7k8iBkfFJ4S
wrupYy/Oenrfb8jQyAQqLW+tnux8gmK068OmN5ebGxG954GMWHuJ7Y40RmRoG9xKtB42miRzenxC
61a83+pvwxyXvKEHRCiX5TUwrsP7/2B089znhjTrRlHJwhpGWroAyZsZ9OYz2X8OzousHvmQTaG9
yJlxCGfRKDiWOhbTuVTMKscON+P4z1Zy9EIFicKIYOfT6rBz2V68HckkTABS78zs9Jr1FzHNqgLG
LyJ3mX4Smyxs5VkLfh1GKhrABdvMI+kBD/OltsyoxM5/omThtAdS6qMHN6IOgzpeoh/DIqrErdm+
uZRnxbiu2NtCdpo7zn9BX4Y4npOj+gkyM49KCqDjTiCJAo6vVjy6Wuj64aUy9L5XLQnOIyw3u5hO
m5P1/HxPA1hDUxr9T8SgRDIVjJhFNhcaxQPWywYooH8L0NwsOkniNOSU6NoDyQQspMxFMh/rmSzW
p8PxVJx9OdctbszZDCuogNNf6MuPyScV4V6roG92yRU1kmYVQryN8Z+h6Z2RyhKewW2a01WbiMi4
3CZMmNEBb9uihV49A8zKgeFAQFjPK83pYyOsWJZOabxZ3kAoDVTghthl9aMhlJR81tE+/pmYte++
csfrtxhnZ4kB91G/y5x6go52ieXAl713+8T6L+vfmEYCimQ5kvC1x7i41Ayk/itJHf/niyDvmnvr
lLoDwZ6diEWveWqsppxud7J6ab2O6k2lMlJDQCK/hohjjqwS8auVud99G/1ckBEN52xm7qJ4Aydv
tRPFUBBVTfREmUwC8+C1MCVx8rB2lsji8CC5OfvcNMrgpOzbu/nk2eGmv12HorpwkAHv6O7DUHWL
OmrN+H4/fwCh8XlhSt/68N6ByTaAOsOdKwRMWlCKHdn5HCyC0UrRos0oELfP/toj5CSpQKfYcMvM
BelXMFrO5tb6RVOKwG09IUhGYtttMQooNmsgsNrXbPaBzLuliWx2LaCG8VXyHAA4+k6ZtLY1WIGP
TiC9DC/LnkIkMuGjrorq7BW5NN7lEMaik8VEZaQJTQzinbFKJblzB+C+VN5KvuvADVErWkmUarbA
NMlzoEMIgK9X5WUUBn2d8rWBlt0EELALmzQ6qnBBfNi8soAht89pZzLGZEFlppFnhM++yVeEE/Xn
JylXE6SmbATwuDint9os8MvJ+ODeYAOMaRjNpD3L0qCcjrYx/HEmkodzmso1svjTTmZt419wSrlr
p8Kcrh/WGFwAUL1qlquV2ICFl5ucCl93OfFcNf6VVl7O7lA2+FO202YS0iyHmEu5LDmHxEbWQ1QS
xBYHR859/dMpPvrJ7AAX0UHTEvaGJZigWCWl/g3ewoP7+ymdCxN0fEPF6HCWiCROhmrp9PA9R0Ic
BwOGaZF3SroAEKdKaEgSlhdcF98uayGf1kwdzYzuuoAeq5Ag8x6+00CcfGVBQ0k06LIdsyYZqVBt
3UUVbBou3E3DIKGi0396AMq9Uzia5c/EPACJS4CJkj8auTybKqlQbLfqv/fK+x4o5E68x5dGwBKB
IdLU1Uk0VPj5R49tc424pAMvztK5gkHcVqDgVOOVFph4lW7jD6i8cIEejbudlNj+rKQJfLYxLLik
o25BfAevqJaOJIMaGLLH3tWp0mvCyMhrQ0HkqnrHp+JrqZBU5GW5QyewdPC1CtumZpXuv6YkF3tN
N5F2+5Sqt+zzhVRBOSwphxfnKoSjIFTr0E+tu+JfyLbqMPs2Ix0hoc+zPO5AUUtjys1afQB5IQl4
7OHIXg2vyUxKxz667eaS6ayanljlhtlcSWle39jQcEIv8X9BnkAceF6ehL7V+bubeML5ZM2jPchB
lExN6NQ3gpsnOtAy9tMkQGDHJAlRZ3MIQT3pEKwNFQVbe549yusr8lKUx/vlSqH5Qd1FyAaP62Nj
mZ8EJBQrPaYAtdJ2YrKQcQEUQyrcnc+g0LaS0wGEkvRmKkbDOcL4lqP6/4I4HEqJ28cceA1GGXAG
Ut530cTj7ys4zmIi2s7gT7Dl6HeZ+oiTeG2UfGv2yH4LpVCukg0RtG4dnFQ2/arKn9i0Q7Qj07kg
sWIqHg/K0uLD6qIJggs2cEkXSOLdzvVrdUKzlFNqN/gzqOz7czqxRll0Bm+4EDdE3BhFURnSqRqV
VoEGz6z81HxHU3FG2+SJNIFg8Zd2beUed538GtVizUiAw2xN0zuHIaJIL1+nHHJ2nJbHobPCwDby
FAaiWaDa7yffZnEk/TIzw/c0YjWnl7RP7I7gudZy71ZhncJBlum0a/gAh2QCOqRpk7sTS6sTvQv2
2+4rkj2qhmIg3FSMTWPpFjAoJhMbqg7MAbkYNiWtLEpXPH6BpJQ+ulhi2QK80eG0lznFdu0vQbEK
Y/1ieReyzuGNmn9hJx1ocd+UgAkRSvm1T7U6XYlIu94w9nCpzOVhQ0lkV6v5LsxTWUOjr3/4HZUl
NoMCAfnMJaw+UwV8pJtnF+2caRqJKwWVhu+I20vzUkcTSQxP0z4Jp3gPw7iEkr2hPgPgVIJ1Iqyo
khKK2A3JlURjFdC4BQl8Uma14JKcqLRfdPkfuUGkAJL9/6Jd1dmh9B4rjJlcWS4POT7i2UwvX/Bu
LzKohmD8VLtxuj2v+h3jqD3w0wVYT+QKfZXVlZ6yp8UDOfg2RLQDOpuAPscj9delsd1Bee7+GkQX
MUhW0o1UF3vv4stDC9pMO51bkp3b9DCof1TiwyGlER73CXIXTrXA57RiYYrWqvzkrXND/Zsv+3+U
edvb3/G69vYXE/V13Whx1TvyPCZCriNBcXMQRtmBzJKo+h8w6g2+z1v2s64e3024YPPIYoES6F1W
pdJMcehEGYvOCxBEQCt/I4SEV4tbwxfevfS495qZlE8czOl42N/2O9W+ZFCV+34f2YcHPwXQrZOI
Z9ZwDehex3iKBHj2PugKQk5yR5H0Za5MMqnkqaGzrlGX3W78yzYiVhQxLsPaxVndNe6OrPjaA517
NtQwTdWm3BILbqD6XOBV4y0N5DTJOURh1OxvOJ8d/iihil44rZ7YfLZw7uE75Fp62gEOhCx8RfFx
whjttkCWNXR6QswogMWVTloj6Ts+xvv7VG0UOlenrkx4dSRVj7RLpW0zpoDKWZ3ebkaXo8TLuK78
QS09XSfxuwGQro8UKM9O0wxZBMsQSHzQgMt2a9PIjPkIaP164bn+1iZ2xfuZyKwdymtd9gSx3a7p
uiTniHMqgVe4EcD3MMqNDv8DVl7ytk5RfJr1F5lb6KDyXSCXnsUlEmpWkkDXvFJZlrx5sSsbDbA/
6AuQF70has1S47SpsUVlOCjPpD0mnaq3VNZym6e9ASnQrNvjgyzisB71qoEdo0gI/eRJTYRqgmxQ
Xrnhy0VLf71VeVb4RF1l9iK820Di6ZGmep5mjkPy8YteOkoDy1M9qzyLa5HB7UAEaJpyDaPUmequ
QRyOswYd4Db2MMYa0FPxL/laNPlAvILkvppHBorPYmAW0a4Oq4wCsA1YYK1rby948u0M+oF4j7Vn
Iiyw1YLCewCuts+rTZqFNjDjwl55dR7QHBbk+8yXQTbGnuO0J+NLKdCoOwrUhV739kIygyea9JlZ
pZop4RefhYZ8p8eDwS+uLIYorRl2PS5cyx1isiDNuhfIltyV8j0Uw19rC/1/ADCMVyrdmGVKDo9f
QH/ILREcf6b5NG74Zo26/SPCzVzki1zFVMUUNZJzuLYvr5ePS+uOQEXBgU6yVIYk3zJWazSqNVLu
XTWjHR37JJJvcfu+0deR/p/FMvnDmiNing9G9Io+xG3Qe12a+QWbocR+/lkk06Hy0tSxsjKU8Sha
ef4R/5A01QeZODcTX0vst/NwL3VUjm+z9Avy5F3PfvpB2q8FmETDXNvYrREtU7aVCzREaJcHNoTW
SC+6AlO2ik+H4YFm2uGccu5lwHVmQbzW/iIwHRAMr1UoXtO0Bl+VmOCofJM67v62y2jRLTAcylwZ
dJtCkr8lT2QI+3Hg+/a3tfYSTNCQwgYU3QltvMYquHXgpYInpuAnK1TRdobeHnxe/jj26QUWddyJ
vgLBukrCsE1x61lqRHjZHuMNQYTlEyeVU+T1eyV0bxJPcGosOzg9BU1iF4LlIsUWziARejtAj9/i
H8CNuL0fKjBOiSJT9d5N8GqdOEAiPfxQ3yjy5Dc8s5/NAbiG49bDLsaRNoTkbG16wBgl8L44qSqG
sPh3QoANpOk+8rLpJGzExtKb/XaZkXSVweBRrtag2fIpHP3JlPWBNvEaMGNLHOaVTSsKbBWmPwC0
KqfMl9H2orm8bkc1Q3EQ+oH7O7lfr3xrnyxaQQy8A3lS4Ywv2qr6SGdlXIqKP5CWREHw112mNJkd
yhZKSt5+ikkGh1Ucbrk+dD3lfIfhIE6viPx2AfS7n6WXK6Uk+oHMSHynRzPIQqEs8f4o+V8EOA6i
8sEwBcIcNN8eOZgqK5Sqg5qjiUDXJB8UAAgGTuZwn4Vn/ozAoqpyQh0JzYROXtlQyfbjQQgPiGxB
6HaftNIWgXgv8POJ1EmrQQjOPeAaKpQXqVCFAeiT7n5xjnHKKnHO2o4BhakXlH6GQBFucziUGuO6
l+tIFjeSCA+wkXBhhIDEeIvStl1/h1raNFpI4mQ9vIr2cFC3S4988wglQdvPoC+beLMOAWmJ1fmS
4w8QIVUSeT6vmGBIpQOQrdlyIr+4HnA2fjg+k9u9xZF6vVNfTrlAQssg18TlwpLMbTGoXIrCn64O
SqoB381HB9mAsIPU8GRjUsUfEh+mlSjmWUCz/DP0nRcgWXS1QM5ty2CgYyExsAt+fAQ62P8Rd3O7
xLEBR10ivaEF44DKTqsg1xXIuc7jBcQzrLZoQN102SuCn1WhldLz3mDQ1Jw31FTcDLNg0vFUyO7p
jkt2n8H5CX/11rVEc/QRBTKCHXJKHIT3HsKZ2Xw3aMrJI4Pw9030ikd2raqtN7a7FkE4L7SNBSJk
nOF7XqJIJpiCwDwihC6rOKfpDedniDBXP5C5oj9uAW5+Olosi8dYaXP7pbxGKKPoJlSROfUynx4Y
LChC9hShC3T1EjK33aMMTy1jvkke7uu9O6KGbxBgyjLIcrZrf376gj8uCa7k+1FXIMJNx0qo79/M
uth0RlI76XtHmKIaqvCSMzwKGfUospmEpO0tCVkJarIpJFmn2aTlKPVjaNgcCdqvgryLO/hXng8y
sepKOBYlXpJldzuAjvoyCLWbj6oi6VFZnMFbpxT1pnO46OUMQDin7ft8Qg/c4N8KiPu8LMWln8ub
9KOkQZpkHAfXwesUgAVWuFRM4pv6sfdgOgth9EUX/0oNhQ0+5XeXczePQmLAiI8dRIekjwaJBKOy
P4OFaXReYB7nU/gp5AYsxU3NG2FB6Z/2lSSf98ayJqUOQ/QQmt4AmCdJ8/QpRLHZDh8mWjOGsJeW
QGC1h54ZBQZejsp4SLKqyF1hxMPdQxT6hqkgme+1RklbddKnUdjUuBbJVM6OJY9z6eorqMEumy2t
MUkyhYr+AnXXZNHGyE9LToQd4cp6F9bDymjmnVpUHVseZXB2s60iMjlF8FtlWbRUsY4RHTGhW5Eb
8whnySm+z6nS0lQYAl1OYFaYLPOfTyhIVt13tPAx7+i2pJ2HWdrE1UiC9NzISjgQIpaVLLSyBKYJ
4Jrbt9tvXFa9i8ngPDt8XMqc8wzxZTQge1J4dawplVF8qeRQ53DsYFuQzRvRBJeVoWxVKezotdWp
SEwbc/105vSuNvRWposqGEgVaccYPz/+Qv5/gWlKcQAPY3jQu4dIYNYEnJplTjV8ipZVYemToWjh
iAqjO5k/gUJD500SQ5NzRkY4oZ2RG+4xy9fLZbpR9FIMWyiulDNSOjtjXhvynj5UAxh47ScqVpSz
FqpOLj+7wxr/o28qk1nXjkDhxZib9K8H69lPKQ/OwEf9GCzYHgfD/Ck56DAAAAARL9UZHS0HDVD7
RW6mMoRGwh0xv5Sbhbm5Fuhn6EFEFtUgKQ1IXZsybFPq/eL8uhFt7zG1Fv6GwgwLMUq8ILWMgQcO
KJ7PTOvQh/94bzTTuW0B/1jr0Dm3xtHUlDzriN7YOhc7zL5+MJhjiwYGqqIqJ2i0MrlGKpL4n9WA
QFGNXSGc1EVENp8bhl0aTS5W11UDBrnfi7G/bDEDv69HNB0Q9fNvm7rwdSIGDi7s8lNZzvWXvl82
/YrNibKK+Yw7oS+blb6LN6D4IijZyT46B/wBfjZQRr52e6WVu771YL+6b+gYmEO4h1vsCSRes56A
+9Pjx9H/5sC5Uxy3Wz03AMjV9ekLxIYZu9INStcQ3XLhs/451RidAV4hrYQhcM8A3CpEEF/yJy3m
ahwqbcEeHqfjSsQl45KKBfML/8liIHgzC9253YI9qjKEkhHvKS6VBh8BCAhoCQXSZDKX5jGCThVo
UyYUb3eZ8AYO9dDw/qrPqWmGcI71zlIJWyx2+K0Dq//HqCXw+drBk22taUTn9orBbsjKxXch+4hB
kHzfoNIWZTvHTCvHyy0jyvYg7Uenl6Hx2pb0hz200X37Dmv6YQAoMGtd4kOPHJjHZu0H5Gl3mXn5
YB+kCTbicHr38aSb99OtYbrnNnL7SfrpR7qhrQ/NaAfHZ6rpF7r672VKJ9lvdnn7ywanANwsJYHz
jE+39LGXFQgBgB/4GliHhiqVWy5JocmBb71FtkOGzKy7tM+ISyfHa8Pj7IHdQ+wHV2jvo2fqzY+c
uc2p+MvjRwUG/e8bGtOYO1iTmI2hQMlT1dw0lpWBs8TZWzY6/JvGuvcjMnpEvKnCZVgoMTXiHx7T
BmQrlCZac4sSsAIvYrW7Jq+ntH45K/d4RSwWHwCi9XpY7hncFnAb1fttIXNTfloS5Qa44NDZUiuv
y7BfFlp8kvO8tgxnvDFA3GoZQiJYqgyZiHIqvi1NTZ1B7VJr76XlBDB/xAYABktBiK6klIzKwVrx
gLXDQcg5q93rLRpQK24KZw9kyxHYuDTJ57n2nUQvStgziZen7OsnYlHYYJcb0fG7GvZQC2XkyMzU
Lz2BUEfVfof0LTaqugo9n2WoWcvfVnHdw+v6L6oKrtXnMI1KYbK9bfB2bt96OFmOgVMXPmPSTlWT
FAnI0iLgnotnM8ixhrGjFtzu0jgvbEK1aDmOeUoQ+sWetAp2d4eHjtgS7ROLDQoGTprB/jhlli6v
sNDpxhENM2qefZHWChm4gEskEfsE431CTDsmutGEVXy4sLtqd+TxChFrJ8kdrj56/JFLhGZnq7CD
YLrRbeaYlaLLaOH/iR/KkY/FE1diWKUxULuAmc0FaNizXUzVe6UF61qKA3lWcUEnTwRq1Mp3FGLB
Kz8y+coXBHuKRRnTI2VSC6+WDjAY53g9WfcxRjyrqP6pqrF54Nk2Ol0C1PecqRLrRCg/9CTIrseL
fzeGn4OcVA2XohjaGwqGgqSEbbn0ROZq7eyedUiPov7jT+qba5/d94maw2n0WYZb0bfa/DmxuVmU
R/A3yPpsH0hgvk/iQB0dbMkUL8JPIN/qx8bEA3grGB+UyMnxKPmFVkqDLisrADB9TmcywoQm1bq+
+4fDcuKN5EXKYKg5QQZRGsSX/xoZ0TN8ce9SeYqPKuwchFtI4bOhlyMiyeS8soRO18a1Ylhb4ViF
bBjpZ/Nc/IoU2WjxHxEOcCZ31neCydMkzAu0+EzRUgRzEoSiiMnNvUhuaW7MLjLDaS+BJvx0Lvvv
Zf8+aXrAu2ZZAYZiHmm7rwRNHHrPxjxeNPoC9rxtKPVw/bLy7RHlC5ofFu8q0hg0RYVqk5/3jSbc
jm2AB0T7cDeDMvBgF9fdCR/i1mxDLDer8sI2tsswXkQSWNBU6Q4l79lBIwyOHjwH5s5aVgFM+xM1
9ujwuN7ZScvhJc3b0HR0UcY9rS205ausNp/jaxl3ziQ4pFG+W2hiLJ9+tUyegfKz6ljtLoRHencc
wjFf5kAgTSvMMFLhY9Bwov0nEGM66kyNHyMVsC0/Ir7vqCTXcJJjQDIzurhBcd25+pn4klxMcsd+
7NS7CGOtwot0wfrx9Eo8QBmR1z3AesbfdLNS/+vYc7U1PiEXLUeZ6CJLD2VLKvQJUXiPqhnMg8Uw
usophrOBCL5EgU6R5qQcclFVx65ystroiZ/5/M5+HE0yv/HL0eenafvkIZsLBhtWdGe/uCR49VMJ
oPWSPmIczirZp2MagGxKUtCtqNp1/HQgUvht4ujr/IaszE64xPhAZSInrTISaaEYH1hYCeW746yv
TgfayEuSfelLL2jwOpebz2GiYgPfb3IX/CyVJ6KHkh25nACQx3srxJfBmYnmpsxOGShjv25C9Aei
XtLGprKcH+tUKOrKzBDgpKM5bfMFoSBb7PUtts2ys32kEz9L7jedCO7C7PMbO+k1DmG5SLAjAZbq
PBNFuuCN/LL8tK65CcyVu91pIPzvbobnRMY02nS4dokcTPrWZXbQz7ASR5U3l6U1tKWOEo8If/Vl
45Y/ODbRB8NHQV3uucvEjipe9MS79SuZdezOXoZMCw0pRRUZ3aR0pPyhM9EnBDNjjURJjjj1G/AV
P4Tn4xjuR1UfhrWEDdeIOHBNaWnRVYGYPXUKIIrmK6fG98g3V93HIohz932aXq8UxeQsf2lespSs
gwmpMhTG4ui6YlFBPaFDJZxjl13qESCumjT/qqisWvmj5C8gROSkOFuIqNqnkMOA6ekdIwIlug39
ZirDxEwzsIx2fshQ4WGDgusvEfM3rPE2yBYCJCjIND6DWa7+Q5O3/EMsZ3NGKM1pJrQ3+n1/bbnH
ytEIDOw0cwcAe3HxeOC0SKrZFLNs2bpFT0PE7LhLUzBuFSdWqFBTEkls/pScyVhNDK5D1riCM7Rj
8Y0UJYFWwatquejuHfZeECKfciSIcRV5z6j4SVh0BMnmodmOtajSMCrfg5X9pd76i4XwcBYZMKi9
9Yh86SN1qCCuTNYM34mtD4DDQ9gxlnmoWtCuldoICWMCPvQB/5N2g8cAYKw7KAkP+oNP/sBmEYbv
6ZLGsDgX7cHcHV3RZp7mkPBb9PRBBh6FjGP3xE6T+bIS4+s8s57gSGPM5oMlQXg69RdefMwcnG5o
wLrJKo+Ltf95snwC1SyM8FjjGkTLOJoPY4SHmkulukqeAe/zDlilh3VTq0oN5a4v8ESLtr5PQeWv
fOFr1nexDKXrj+7QVBG8uX51BaSPZs+flVr7AMLZdnxeYPvUMEKK4ZdJbtVqGTZCPW5V6S3YlFMW
3mGoXf6SPrEgVmshI02PWjIT4zLrmJjoU0d62Zhj1JG/jbRh5BR9M16SotW6FlvXVz4CHURnNT5m
F4HRsnB0Sn16EvwU2F7ycMtwrE2l6cBU0mbTPbj2BjiYfZhd2K6N4SyDZhTt/0xSTVUoLDejkBkU
E/ua0NIOgflb8imy1HLPHxRpegoOyFx7DiG3wK117DSukrpcOOObwbiBw+zoCXIG5/irmbsxv+rd
seR27WMDvgNvyyObaICdjpO/hYDoYx74w57Kd6g6y8VLS7krh0mt79ITAOzYrEivjf3T/G3X6W24
3yvcrc6dABrZTog3RQECi6vT0Fot1E9UCkYEjtqJ1GymQkvfCUd75MWcADQLmHUW/CyeapGsw6/D
mCY57EmihCXw23YPV9y9C0B5UkrAPucGteQ61VW+DYdhtAcXFksskXb9BHdYezCtTKIgjY3JstOz
SmAOndUpcS/dO6Uh4xciPgkYOrjmKsXMG/Nx4aMeTT4M3p8qZ1ZLYg2MUCgMudwgTdpWLwwN2BH9
WqLGnamF0XKe9OdUi9xGQISXp4GnXqBJxB1sGXBOAX2k57HpJjxzkzjLM8+0J/cGGt7rkvCE3aa8
xl0TRdIAf4ssdeU9h6Zs002dUtYt8FOEg5v/XazlsJYYbJ4iMaun5yFulXz9IafdTFPixXorrfnn
8r7D00SU4vKvnEAXXEiVECN89O4IeYYlyPzo95J8mi2thIBh1UqLBwmtu1R43VS+tu7LOaGjAaFE
iPi2xrpkwq1kIvK2WB3M53IHliDmNK2OH5HSU9g2JAfpsw/tfRNgO5MO2JaK8R2kuxvJuuFWHyvy
unYs8Jh0uFwB+Vw+MVQ6j86ePcx7WQnZ70jOLQ5dQcevd2k+HVMLPLITAVBK1kqkXLXby0NmHzSA
RutGKW509a70hhd1R5xH0o2rrrucarYwWb8H6OuXugDZyV71HPaWggXB4qvx/HbyAQUQm3Kotbjj
/zU58LcsmMf/rKGNOQ7njLWnwjRiUqVLaJiiyviJfv/wg4UGOBJP+opiZI7gZvfqE+waI33Il5aX
IOB3K+z46YjGSB2EyU1ZXVbX6I+TtIctthHh03ssSWe44cjHQNhHu+bM0B1v3f9UmK1k0oi4Lmbo
xYvNbmR+de6iyqeWEC/98dv5h6g/bbdfD/bQjCKB6F6BzP7zIXEV8GdqKJFvUpziW9k7SvWaoCAG
sPQshZdXjhaKpNQrpLmTOxggWWXiGuHfVV2CTf0v7S02KUccmo8VbQUdRYYpseuhVfPjWBZWNo58
bzLDBDg/v1A4bv2S7nyL5ebbSOx0IOiIXQJqoRbqyh1Gtsw7zUl2fjcOejFDttXgAdPSfimAZm8G
hjtJTzubhkx8cfWpXmBohZBftsGB2NrHEatUu7YHmvYqrZaqWgJm5k/hLg2NcJQyzwy5YitrvOwZ
r0dzF2K+MSZHeJfLxIy8pf2fGKP/nLSfHtgkP5cE/D2EAir51bYc4gOBWkpI0FBzbNKZxS06FjvV
tjzMGEDi2v4JUYBftWODmEEYsqegaIRx6ydpIJiI6RwAKK64KkN0M15OaBEa+zigJx9buRrfbmxE
xBoT8IiIZF8iVuQcPJ0PC0Ww9uulu+U1zVPMSXnNivj5CPBKgw+iglA/G/JTB9u0YMHfkigJWZgt
9TdeJDpEjigN98TdrGqaMcvhAJbSfU+flxgj++tjZf3ZtVBESy36UcXdZB4pQ9ag2A7f3FwuGRw3
vSUosO3pBRB+gB/5W3WiG1U1pqx4NcEuk4XU8lIBKb805+jsAGZ8VbP2AHFYoN8fLSgzlwR75BAU
ILfw0tjUxkfbK2sT4jc+7Qwu/N2xt2H9rp8Uon6bRv62HfGBzydnzVA66uJu4F95z8C/wIkppJXH
jUxxwj09kdxjOMqM+BKLyZlrkEjPDTeFdTB1JOHrfQMzmTE/rr+7t1UtcljUx4PApkNdjWn6QicM
aR4HnNl5+GWSgk7lzAi+gec7L7VRawq+rmYbnBCdqnvWSCt5Vsz7kY8VH/DWlADA17/WIQrX33W7
eNEP1G6N+7DNrcmbGft4PkXM6PwonNMy+m5S0Suw4OywatBsxnrFoDFG1COv4JyqNwsdv9kqlIeZ
RxW131OEQCXZ0vZMK8vlkX/4LyB/G60UemF51GEXdY2vz+yCS38L4h1tZWgwjdpdFiS0qoaOigGS
lZXXx6pVsXKGG+2IsW7prQ3wvTOAKoVk3gPsHxT5/M3Ee6KDLhtFG69wevHHYkvQx5yjlJyWjAD/
69lQ9IH69Hp5jZERprdRpqsv0eqt//OeI57SshJA/1aHq0REs5WDrHzp4bpBjaxYwYvt1TZIDBT3
hjWl2d0tkR+GSQzDtmNNScH3LKhH9T9IOWVgYNW1sBqb5ldFK8m1nt65Hj9L5MOH583x+NZKnpNN
LF2n1XmCOeqO1l4X3FfVjym+Lo1GpRaFDuSpoJsbqyo1qmjUQX7yaypDrNHlqcfxnWLCzfYFKVmf
o3BQjBVeBP8+ef+0H6h995gzgt6YuhLHFeAPcyK3HfiEnucH0JPtC3kvRxJD/qg7O0a0jJUH5r+F
iGwKPU3HOzLoa1appOZ2nUeKczjbOjefzRvgB6as+N4IPSAbs6EVSXfAjeFXZ6zqrSSgvb55C/AK
1UHshpDfVCPDZYDT5cmN5NxblNBApbV+PPG1LLifvead7aWl1auIxsDJk0gfr+6EkE29iOp5/Ug/
M1OHM6HnwY8DI/V0S13gY/Al3CYJYCrXjb3czl95nXe5MKuosIrXERHj2A+QzikOmrWuuSUc5suC
N8CF9sOtKDBwdC6srFZ4bsNg2iMla7SN+kkD4kRC7kDi8Z2soimXa1I1HfAMZjAPA451MdE+NWDj
4A3UF46bHLysb7r0Htv2qgjXZDRgtwJMDwfVVhqizoTAS+2lm+9r+wISKFD9atDClD2A+pBLEF5j
z2n3inGy7DJP9n6auBm/PDCBsnArw32THEApwKR+orS2wFLqIwZ9353XQKFgYKNRxE5vVg01ZJxJ
5v7k83MCaga2SsOetsYYruAr6mT9Zgw4SKGj+etHOelQWgVe/uitZkTRMQyh3L8suCbd/uyAfGP5
fpS76/zfl1n+0OaPiK60bYZB9LjeFADZCR5Ea91AvK2penTBEUbG2YeXDK5Q5TSQlYWbA81AVcKX
ZD2AccB0Vxfv0u3wfBI2GPJ613W3C+XgBDOvmyoGGnpEZO9OFcdYLo91GshUOTt1lg0Y+vyr/opM
XylY0JbRARiZos/EnvscgmC6UoOgnHvhK8xeP7L4C0wvdA/9nAvhP8qAoG305+g0ALpsssI4Zkz9
hbNYQBt8jVLpxcUpe4vX6MoczEXWDOMMWJsWW/xPI8HUSzCiyUfkTg6pzlNvng4jCZCVbL+XUif5
+tiVBsfgmdsIRD7IgVBnEyysy5Yq8JUt4hIBUFbtQmnNzkYY3ApEIWhUTL1yGbn+9wleXUbv9Jky
kaqe+5Of6wO8BUBWqo4nxRZq5/kmjKevg9p5YgKqHCAcLc2VCVib8auhgNju6toHatnPKjwmz5qN
ap9YTiWnH0GsAGdJMwMc39TByRNFc2IQOdmBNw+avbrlJlLLY1yStqA/buGL4XOq5IODdqp5425w
k3IdU19UuQxxtHtFkYBhPOnl8lH3uDCuQ+S3aYr5Thj3jhOS3D6xXP7v1WsRWCMCVCm28uhqLpAX
KaqIgOi1Sn9jmTDZRXlAXUxLT9eyvCEvNnZvrFACL2JNVG1qX3IPSwP+ABnduh/HUIAscIbL45fz
olqapK/M1coUfXzA9vxN97i8Re6pYvGhTQENGU0pBfA1tXfLNItLuEzcQGCTwjQC/XdMX1zDhHYH
cPTgpECYU7LpzKcDjXFiC+KbWh+OkGPWtZDTUujI8udS73GzE1d0vB/kpHatf/4xuFC6Sx1Dr0Gk
Tu3wXfhqf4LzHAsL7RgVGb7kncs+nkGHHpGHYj7ym1L5rczeoMJavaN7Is4iAuLicGgUbMy0Y9vo
DN2+hsfj6/uludOiVkJ1DC83VUTh4cKUEU3v674QKFxsgYbOnR+a5ZjvPZB/ecHOl0kKwcS1R6lH
QEE6G5mD5gfLI0pvA2o3LzjFsuYABk823ljUWRkwc3bx+qP7957ziV9pJA84x8uXhyUipI88FhNr
lDLlqPcQWTBNgMEJMANMS2pANNekPt4nnTv93haoLqwI5qFMp53pvxY8o1jlauMEpWxTufI96xQg
pE1eWMh31ZDq79WUveF6NhwLj7Vf+qkxtKBqTR8KTP2ZNgpf0y4xQKYdRYjFJYPAuF9pTRd888Io
Tqb6ht4Cfe2a8hDqnt7OuOV/wWjxbTpH3hkEhz7B3RsQ7VjphR0KnXzBvUvmHo+IDR87XFzHuLKE
uzJytD68Ac4OZId1GbZv00+AnFhI//hN7qpMn79YsnN6dHTF70YYet+CrZCRggF8z2hunyZDSxSC
7WN2mW5BGZX2Xq5xfmdnQ46QLOeE1taXlGDryXM92UnBvvFayLn/M0SPjvx5EfShC1+7ATojbr59
wogrF0NTRXhaCKkZC2vL6JPlPzjPaQHANxP1F4xA8aWBFq8hHl3xAPnoHXGfnKU2pj6LftMTFtET
fES3Oq6HIE9xDGjDHLdgt3vu+7Gz4DzuddsxljwhZhlKYGoINULjhRTJ2tq+gN7VGc3WeaEYYKLj
nbbYxuYWR/m7fyRGKAt8Jsc8ORChYN9lX+EPX0iYgkqwHpzQRcZ5FCRmI9sEG8JwOQnXP8Bq+0KL
ArVzW8NuAnY3sI0ADnPL9RHkl5hZEkc78W1ovQD17xfOsriJ1P4MQiIjplq9OBHLL3zR6s3wQC2Z
TRQ9DiDjCVz8/HodRuIRI6v3qYsIv9H4LPezLk+FpJRSNUlpsaX/Paucu+m0KI5xsnyn3bz+kvHX
L5BVoAyDBI5Lk0pVJMqU2i+uuxKhxXaT3luH8SQQYHYYrYJ2bJkj9R7EiVNLXP1+bWaFnOc5PzLh
OC+5ldBJ20CCIYPmN7cotUYvdD0PZfCPt2NALE+zrMDNVxZOx9iad/WvA1mse0qkGZYdFKFYMlJx
QmRukyaq4JPJelRW0KZLZva5/rD4kZ7+T65/Mf8iYKvxfrMfe0DgWVUoMoqX9GOOktq71SwWbLp2
iyVAvClWY9w+QCR/z20uE8yLoNMAqB1YtOM4hF1NizmVqKzYrbOjsqfrgkbzksYtBdVPxMI4Ejy8
acvtWfgSoVycDWZ1FfgHdCd6h2IKClFTonCy8wngWTHk8t3umT7aWZrf3I9/o/JIFfBjUMrm/EMP
o5tm+g2diBCvdnGJma2MxJLx2/9CLJ/x2G3pWhEacHE41RBKyho835tkw8uvnMrHhRwubRFruGtl
Jyz5pS3duHkbc6CykWw3GOSwoMGnXYETnk/fk1inpXFwohF3KI8Ase4kVs7vgs8kOBgaO3cV6777
l8kROBn0mXWJTnHRpASmeYrpeMVQqCdk0vWB1+cDg52QWCrs027yeJSCXuWNoMl0yklzuSw9cL2D
t3HML/sPVFdyNcZ2fs5XrMe6nM/tQueSs4VeceapXv7VCn0/pQzFz47bTr71WfPTxl9IHfTtu3yR
DXmX8TKR6/i2CCjDhiUc2R40K4ho+jPKZPEL4q7L6zmjB50ikrIMdvRbPY3SeE5xyu3tP9So82Cw
gMVcO1BUKeidesfcBKYF/yJvzrDfwbM5l7VoVHzzfxR/hcRyxUM/kAZjWjKRJSeSefYNDpmESPuo
0I9SQiZHWWsdmne7DLKxW5Rut45vdoh++TzOpkSiYxRaL7acQDoT2s8ZfBlknZkqgBQgvju6CthY
gLnRYb0ScMf0t37WdJsDGeHlej2uJ4YrbzytrP0+GST60OOmvV0kIUMYj+9LeRhc6P1HZKGbi8Wo
UXjJMw+po2Qfy/hEdnDZvvKSYfqA2e797UW941lyvNY5YIdhuBsV6nzZ4BQVonviebzVdAztGOYP
kQOdebKn+0Cb1CHS23dfV4WkWHZEk+ZWRyRBrUttHAhuH97qIITqhaHZZn28tBw2M/tXTnW6w/JI
Lpkarwoc3WzYAlzDEUWvt1IH3JWxx62evUf7+zoBAt6v2YRaV+uh4jIa5CgJOfM0zqAAt7tfR9M8
lEaFEFdJGu8874fbYrqJdYLYhzs6SywLDzk6q2wUuV7N2m5E6DyA2iwv44gkMI3h/at5sIeA1CsL
8QYtRNUXyM4Cvi+Km6nPRa3L6pI87ORVAy+AL7sextdMLUqozVRa4wPTgUVkzvPqDmECinGzqv3m
Kidvll172stdG0r+F3tskZCQEEOFWjNOPkZReJzPrdNwxrJZQVZUdPKLMjuDkBUedD9kmhln2cJv
f3+uKr2VW6awuqIosacBnzG9l3w32ZshZPNtkK2RMBS5m3VJS9TrIiXErlQZSpAzn1RY0EaIfHM3
YXPGsII0FS37a1BlqSdkO4rtLCXClM65xELXW8scdN/2heV86oaFjuQsLO7OJpgpDHHsw/06q0Wo
/dWGiJtc0obqXfx6tFt0ST69FpIAlG0D6dM7RtS2/4XX/A5+S5q1O46AN61hkQjiWlK82qJyus2D
vGe94nQQO+yRGy2ztLYhQ9Ry1xwK+ND0ZIxsKZh2xRLjsbjMQlQoR8nGIIj3JU9yXanORerB5Tcg
JhbrvlbDUta9dfCVk9FUZHfm9sNIKHSKRYid4xLBTEfn6/jRUnEM/v0yzg5GJBnkeDhbfSTQX8Zt
1pxPxhhFzEg4ZPddvWDCCewIfi3e35xfaYSGO+7YJk0NQLaSZIYD76+HKANbQrUwPO+GR53wvdaY
IWCwJ8Z9wog3iiAB6Ju+ZUfRjF5/dC8aNnNgpE7PJAwk/j1jszBxYzKk9Fid0iRkCGACpDfAnIeJ
jyZG5XvD5qncacxTD6BkrIe2A5ZwEiZBqLPnp8F4yhj+zuig6lolcyh/OQjtdh51H9dGevlAEFR0
8n8mgl8Pgu6A3aOR/12Sno8neMCZRIxrWifySoLJpBJkGx5z8vT4O1MvCpX/Iu7vCukwEB7y19qx
fpks3iaoq+eGDTyA3e9A2Bq96NKtR7Tni/MSAAwSm76TkXwpY3B5wcaoFJ6rLk6ybSDDnRhKVRKf
rcDDkEXWiCGyx58aCkmLkVT06xW3o5Ae9Nubo1DQNHvmvSdUlByHYchN6LSmdaUfdw/jveF1qvOH
T8tm2tBbP/JjIsIyM7J9ltXIe5L93tMqTk0aWb9CD/beFfioks15eIIPqO1sbUiTmus0o4ibUL1m
Su+sXQu29WJ4EQyff/rTMgRwBWO6Hbtd+jsjAiMbiBuQOWZgJySN4PWI/nEfWwMTZ7GLfGWJVUg5
NoR9ExNL93WpiGghjU1Bv+CesEpWdwcNWzfDKJYAKv7QYlj9Y29ouyIB8Wq6VUd0rjeGZ9hPJ6QD
RINkRBn+1eewZMbcBLQ8sivd9uq5afbcRSehL2IIxOWywN6iSh2evhP3Rv0Q0EcsgYtj6CLnnwfp
xQ+njaN8MALQ0C2Mkun52ayjzzDhqzAaFTRYTQlJ0s5F3KchkCLXT+b9i4QyRsqbPa4CrB8KSmJp
BSCJqgWUtt7cUb0mRg1FB3qWMicoN4m4C+HnJNAdaF7wt5fB7QANTMBf9oBRG5/5stwPBJPRyRIp
FxdrqELMFe5naY/qvgsUHRfM7n2mWFyBe3ivFAg8C3MFL4bkOV43Mt2mjszp4U/6TgLasXZp+nyl
qI1uQ+SuRi2f/6cWZqLeRIpggYGekYXs+W6nVGxgwe1kEMslIbkOMf/Hus+CtSnPKS8n5r/RwZZn
iveenQE45bwdmLbIJbb2ZkX7SHAYNGQnjfyEc2AjH0TqoYSkNb5faggFeCvBb4DHFKrKDBuhqPu+
nkXh9FJp8bERQRQxAS79uf/94bmesuuuexHWzYjkDYgdTXZ8cyMfKP7MSNxQyuOzcvcdfbdVcRJ3
gKBgPHc5nLXTlA6SqgRT0cM4zQuz7OhQgts9sYBgRw4SKM7/19n71W/Qk+E8pv5YbEYDxsNq+x/W
i6BwWTSCB7bWMGLYBKni+gcUzRHE2Jp6SHhsG552gNkxCp5kATdLrddRT/dH1Ub+V34pRV06VFvx
BvZkQhBTjgkM9ouXHiszADl7wZGiFZGFmEn4NuJBfXFiQTrd/oZ/uPq8o0ycR6oQBezBXb9FCG8z
0B5lA8xtn6Y+Y2nxSSusbizB6UCkwk5KRpcPPTwenvDdSyYaiWRsktHmpjUSlvUu011a9CitXGR1
CfKcj9RzKi8MMfMIL04aSqa1ey69iOHEGmH5+s5C2njIziVXf5XzkIfHPiFwJz7iB/SmQ6sp3roR
NRwVppHozHgmDXyidTG06Th8TGe1k52+IAQrJ6qmR98IqQf0oquyJPcOuCyST2ixmtg5I8ajYxxU
m5ZjN7T5hGZU0eMHvr49Q2vH7NWz1ZR+FfKWK3hAJoK5K3mnBvz7HbBEbMkqRE+D4gaEIKLOwCgr
G+yUkaNLK7m4duGtHS/g4n86JMKhjnqg781p1LmVrcA3k/RsJMzE1BF62WkusF1QynICp2MRQmwj
03VO2GFFS+ViGtjydRqaWw3uys/V4/qNTQ8otKK6oPyO9v3UU622zPVHZQ8wbxjzbqjMshEU+e7l
cuUa9zvCkm55rTAJlxTN5CiC7cgGikO52CdXX0mvMnkJMws+yczrXZc84g75pERfq+3aQaIfnMSw
giQpysbafAdk7T9b/WfzM9HjJ9VZAlmU4TXEhiP2L8gcCmGxOxTgs0M8fDQAKQ+QL2+soF2hKe9q
kra0lzo0p5N19ohPI903D6KSsjnbsGNonXtlSLC59ZMk1A/4NogoSkjForHvLzpXKqIcWxIa4Cgb
4OMDnbIzOSEpkIZgk1Mku+PLdaawmN4RWs7PtcP3UuSBf9oKn/DNqQ0I/UXLU1v4zUvuhu1IFew9
xDwLF2rnkwwUrnH+PP20RaaMktkrTSPFe7b0nR3IXM9oiFV/e9hlHmPzq/VB2xLtXITCA+MFE08P
wNVycB0TJ5bKwjgMlShpaIYaatlmv+cSxZf6/HjyqQ7yjFP10B3PDT4Tmr7Dl5q3QZmDelBycHIT
Uq86SIU6oJHzd5PrERzplyVu9djtjhFFn1X3Z1Nsg1LzL7UW244Raac1v9T4wBnH2I9DchNZ/mvH
zQW3/UzdMIe0EN0Zz0gKBDB05dmIj7mMgsL1NAQZs4WiL0qdY3mynbao+Bv72cTH/SvvBpGHIk8L
Em+4ah5SKk8uhxmBRKM/EDCf5XOqmDobOLUQPTgU/wZ3UW9DGddUo/2jnNQ8ccHuwVZbwnGT2Q/Y
5iIqh6onRJldMAdypW/5nALDrjruut8BjP8/5+IDG175DmmcbaRLsPIqRXhPWkJrWnPVeAIKRe8c
gvsGJ0aF5IblJZxSEAxywDBl9B+tZ5+qpBKOG+IlHIKJtnQbG+gOQ/RSGPTl1dW3tItG7mEkPnEp
Lij47k2c5s1Cs2Nn0ODGaRrfgmu6xSlYyFK+wPbHP/QI4qLukr3psC2Sk12TkIk1AEerYlRlR22I
1NejRj7BL+nPKTdzkeg8p1lHk/ffzfgD6Sz4sITbG36svaEs8NRl2foggdSH2ZhJX0oVpu3WHkDV
d+CM6MOYBfC7LILD0le+ruUStuee7RuZ2+NGmV3DyU1bUjoWOlHwOa5+9WWT3z/ljaLnNHH1Buyl
jNV5CzYG5miYvIvP010zxYs/OCeAnywuy+9DGmU8E3/xKbpcLNiDUFDc6NwlIiIKahL8XTis24Iu
quygl1/W5ZI3/eITNbqfHvcP/rW47jyQedPB1S+qKFLcq9dsZA9AMy5xVCnhYqZn87S/UvImKJaH
W1aTzCRcp/Qd2yiUNDd5kJqss4I+XvUSj6jazWPYJmLpp4bTwtkfpE/Bj447MBo27OGCjnNSXNnr
kfHzeUKaiI2Dx8Cptd3d30qQ31/+gfSIGYYvLrqssE5yZs+pHSK6P80q5IWseQkj8Wor/zV2mdWA
mV2sZjZovrb2r+8+fpLWQeL8bsm7qBKlZNL8WXdoDbgtsoxtizp/9dgCcZKWa1kPheXDWL8o3Axe
gc+7mBrd2YcNps+yaIEGZA71VS0uB4Xh8owt3/wRZJgWJd3k3A+iBVI9sjr4jvwBVzgBZbFJWV1b
uu43RrLse9I0Hgb7qySE9Vv8ZQ2Ns0n/BGGWZ+xR1VArWeiWhNM6jnKXmF8S72p1UAYr2kyp/bUD
XWX/OZH1SeZj6JynTgTu0umr5fQbQJia640nF70t8rfZJu0YUhFe6PAlpGbOuADSMooSqZ/6EygG
tbHQfASg+9KK31RC3BlRMxeNCfRlAF1lTkmmKf3cneBjsDzUlaqjtQVFekoEtvrJPeV/M1qQJius
0S5GxXp8/dEsK+iUE6MQY6/DQo+z8bOAfy4XMdrg4qDsuwgDDUPZbexGSN+j5Rzg8xZPVSx1qG6Z
aC14536QjBhpduQSfERc9hEBK463zBurd3nn8gZaWCPzHM7CpNzNaO+43Jt4zrjwSWXCjeQno+Kr
6dVbH/nqh2qqhuZWTsOU+ep2L6sB5rKNHU4co/gzPA5Z3V2FVG74OebsU4vh/iyyEFL81x2v/FLs
lzK34QYAKi8fTdDEG+914PXKZO6jGdpwzQU8/cmA2pz5f5TlxYRycUmapGgdXmOLUw8T9Hfj/uWG
ICQ/B9XaxDXlhuaBtSsodQfCoRRZYT5J8hhM2YkBF3fYgL3FCj0f7LqoRr4Ar1zFObRgJfOtY5xF
zXzDVydpXJGgA4KJ+UVhtUi0ukiarg0AOyImg5TGj0cNJja5CXRF9PSEDJ1Q9x4ihCg797FKALn9
TS/rRul5uLz52j8T1Q82W3/mP3+qI0cxYTIJkH8a4gYzasNrOWQ1b/eKw+sZH1MUCd+QVjPdsNE1
zLjiz9OoU+coTGEVCESMxQ7Fwkr18MFQJyrBwhPl1+tIPgtIkhRGrE31HZf6eK1+8hJXziDfnGyd
M+sopBjsq+/AMeYv4ixy2FpT7hlcGAuvorR4cj6pTKpPQq7mKSdOpZIkKmec5qzXzi/424Xm/E9p
AdLoafEaKuf5Pddno8AI8qPpC/o3MF6ufnZEBSNZ46tXOmVUZEigKaWDhaWGF+GRDtV+XowgdXpY
5LBzzoM0tmk2/a+L6FeT18ugPYa/1AoKgPaM1SIcGzoZJ7/2pmuPzDQ7UXpKyBXOPk/KSOiVAHhA
IAf8D3uO70srn/eNH4O0TLNdPeTFpthBIYYSKe5N1aCdgaxA8Uw0PfdAFwxrdwf34x8k6H/FThan
+K+zuwx0IgKyLJV7p2vozzuEewKw2mcejtnhqPC4gXgUwCyKu223Wf0Zbg6PzEP55aMTSUElwSYq
rXq1no+pQVH1eAOMk45KWpOOmmzq1is/6G+XD6RHF2p4jt8pOUSIHiDEMGFdJvHL9xbS6dNdovd+
vk2drqoQOecOpsTNpp3A0oPJygcpMIQ8Sgz2BzaCoXZ+GLzeh330GXiy1DzxHHbILRCHTcMkw4TC
NlhzvoLD6gMScU7hMzvYtzHkZu1uYkYpUt3Aom5AEY7s7TVRXDV4UpPBcwkNnW0mGZNJLdda8aC+
FxJCySn3UN00KDWC3oZJi+QHtv2LbIzIlGANWKpKErbddAR9fv9ylzF2aoS3Az5tr8oORkq/pZ1O
V1kqP9pd/CmD1beNLw8GuI52VKOiRZioMpEg50xW9vMPFlz1q0NHzfUE1KFExwFcW3IADssM9YqH
9vniEV02D5yYPDOSi5G4pnU1wL/OMdL6PfysThyX7SweYiK7q3HSwk+cXwH5FqR1CS88rWJVbR+N
QBOQn1iCA1vxJAwEA9dv2qghV7Q0w8xrvQHkIPAicaHbM5sYSCvc/dol2wlNqnJZq+UClSPVQsfc
oRbmVqn21I43qVX4tfzlnpHHln1ubx6qoERj8QRoE8Uf/D/qTn9RnDs9aPNZuxGlqyMRb7zfd17+
eW488W0oFFKzxCEzzLyztFijeWyXtJSUm5NsBKiL6YxIK5UeRovDkRCf2N04EST2vb8/Tostr4v8
gYtVlZ8xNbniICeJr38JfNq6WrMLZVzFgop+jt4+cE3BJMjNa0d/xspyKeQ3CvpsG0n4xYKfEYDh
xgXJobPI92mawWTUQGomJ7nErklnIbNLe+HGIMdIaQqWAde7bFTnTQNkXLSP3J1sFWquN8cPtrHb
M/74LcU/RtiP7N5xOvrYuclYJSCV3FObScHfdjc07Tehd7jM0qd1TbutDTG5P5Gg3Tc+MtdDy7ep
66nIln+76jkuhoBFYTsHO024g+I5pRdTJ37eixzOlVq3RKvW8D7O/ob3Sujvp5IlkmORZrrqf8jz
cPkqbB11EFVE1AtaOHn0PKwaXKNFM5fFcNeUE98e4TDQHaEBda8R/FS0KJ1lYJDGw5m8WhaedFRS
27ZwIGzwNeQu9xU6chu8oWxDjJUzbJz72jJNO0mm9TtNBEaSqxh0pVEXE7j7soTIGcmMvUYgrqNI
xqx0ZkWYZdqbcOHeO/0uaD4mc2upxN//oTD5QI5Z/MD+C983iRXC0SfyTMbwp4vTYuUx4EHZKjvW
qOZArhdJMIcziKU+uzFG0YbdwcgptD+zq1hlP5aeTLeBHVjEUFlpD4/EOHAbTYbAyL5AvWNxq2Jx
Q8ph2YyktGllYdjBjO2vWAh899RzAIr/OnLT5jtAOF21G/8rvZyijsG/tC86MqPlle87/TeJIQaD
pCVOIKrj/iSvV+2FVHMf+to8ji74LuNHXKjcD4CPEDKti9m9LIg10mXPgnqzb3g9HJyn8Soye5QW
89KeKu5Q+v/n3wpi62JXBr7ZT8yJlt/NjtzBcsbRqJMv2qKbmYM+5TqbUyy3emDeOlzjrFWIiJ1n
6gbjTcGIV0s1WSkGEHXNmRIs04d2RBfsnbOLwh8X+PkALfSux5C4abyJt/2JfFhKbUnjKUQUwLiO
XxjQx+Ewnz+nn7ubBDblgsSVcfRxhdEMC1EkZz0h343FmM3gDs7ktviDDHIHJtfIBbg+aqnZMLT9
HRnNzOTxLTVsCeVYzwymZPIBWchFoTd7MHKsBwlXqFlV8UdgnHhe2KKtccVbFmHzEMv2OX/CaZIj
uZkkWSjSUrX1WMPorqzMh+sQ4ojctH6q5aF2szxw01LYhSM/IULR5VxsYGndEdrCSa/8k5RBUUac
LQdDuZzm6IQFu/IiPuV32ftjWOerEdLc8zGZxCDhrdixNcmeYwss8ieUGnrttIYvY0CJmvDQfCdo
oRmrWygTSjXjbvvDnfbwmwZ+tw7uMZXh+tKKB6whH43viRY2sxJTizjbgC+AloTbV15dKv10sDoE
ILy0en7o/mZMMaEkZEjFhMTAa2Ne/VHblZbFvnqPBRGVQj3L7kcwQ/cbSQaiPECutuTO4rgKrgHb
BEx1njqOKE6eQqByGvpObvHNbhK9iBWvofEONwXEr/UyOiDgYEBHMlqTvouZF1SrIW6Qb04kAMiC
K5lgLO2iHbUNo4Xz/MxwzTnTp+0zJkCwbnHhJellARXUD/KrT9506XhHp0nwvlnZrJMAbQ57bMpx
p9M64YKvdl/Ium5cpW7WGI3Hbp6nW6nhdtaPJCmF47qFUhSX90Ct2U9KJ4zylvCYF/c9b4KO8806
UoDYFH3uSM2BUW7wJNKa5V7orKp0wYBvehTU7mjHs+qNZy7Wt1hRx5fE1JyvwWaE55HfuaK5TDEb
ZspNWd/QoyY3QSqegOI9pvYZbofoqpzt5elTZPHQgxejTN8GGi5u+u80D0+ByaM4/AVEp6hNGA1D
csOvWVX6uXvwTeRDDuT81mtK9GuDBoI8iM9sIvqdJHXXd87/hd9RzHA03/9iJ2tO0+hJ/Y7KLHi5
JP2kCPubkSPaqiIfx1ltIJCB/HAIZ3LpApdQV/eAdvnM3So45VNLmBqkhYgxAxQCti2UCKXyPSaK
iHR1jGx7jiBSWDmXeeJAnzLeUSYSpkwH/Zj/JVWhpyqBcM8cMjYdbsuO+kgFDa6g1SseXflvdLqE
QIwrroiqjE7hlUUuWJYc+gjvfIW6rTPJcig0SnPzn0L7f7VGU2tOz2Bp/O8/yJiRw4c7bpYrNI0G
wY0c77ZORD/gfrTizgsj+SI6Zxr7jGK05XJCN3vDyctFN97QffbbVbcWl4DuWW7hD27S9PIEdoLY
sXTdtPJFWALt/Xs0vCO7P65yL4D9TBy89NBXCFreL4qK2h4DqDcUJM2T8UXCP6zqZ+uzoCK5GVsC
VCjVu63s4weZ5pEIudqboSfhD9TyhTDZy8H0/IlehOir8uRCUnFOLlVtpxZ7V1B2/cPqFh6FZXDs
jp73ZK4P+jS/anwqYLML6R1yqs2YsUlyQyyPWz3f/Yiks1rC7ZcQFdOvJeonZYMI2xN8Q9FlbZzY
jmfRLk52NyaMPd8GUHB493LlMr6HU4jvypKiwGxImkAaCs0+Rnbxd14DAwQ33lEpKY4zZJtKw4G0
AIDr/DzvFlp9n2Y2KP9wVXcAqZNao8FkPYbjL0sJyE/iNfzX2nFPhHqRCGeDbL2Pq6SO74fIk4zQ
T3FDvBJ76yuiR51jEhaQR+idpx77wIG2LySTLC+/C07YlQWWrTxJW1SEmW3DjE+qb4FzyxHUw5gu
s+fkaVKY+1/P5RwuOkQaxr8G8c2Zr/jHwXTkfNUy5IfdpQLaWWZS6bZuoK0epGPkgJq0Qm+hAjIX
N6nq7SZgMOC8FB287JOULiqrBIdUjKPTv5W6+VAXo7ViTFmxY2ukRPY4LOeszuhe9tzMKNz1ZzXp
KX93hs9Ls+U0pcVli0gOWESuv5q9ufYZxbDgE9SNXLtJzcitiNFWYb14NLLq1KZCJ08mbY9V6xUI
SeGHQghbVRyO7Q9roJ2dXLNiMsZ4JdolghI4yZ5Z4ST1RyFPxW7Ppuz03BovSNFm2tItTWu/6XzG
w3nXpTXvDzyioZT1kujjM26ZJ9RcLKhw3YZNJfpFgE2IKhfgUq9qlf7aoXha7MnR8P+tKdPXG/O2
L1/11pI2cr5p5vgIU5xpyd+NPLST2eBomnsMxT4w8NSRsiDcm3gOEMYLM93+qFb2b9p+to+hBjNC
kjCYcHFBdQB9LSmVHOtrcdS+s0hkRS39fL9saYkUvMaaQy8msXYwB+ziASHYI25zBeOLiAiIAro+
EHJ/9Delbbcj0A/lgvAuBqDVx8rc7RIpiZmwH7/WAsR/9YKZ1fXlh41fMlwB+SPdFaK3RlnNWTOD
ZbYIZOrAnlyWXodArs99+wY5+IIIWbOIfOlRDJvhnjrxu+mv3nw3DaoXCFOvu27ORhbJ0X7gH7eQ
N6GFrszNCuUfYupYi89Oue8qDoSRKd2NT8vVTATBKZH7WOXur46YyhP4PSptR8olf0nNEdwn+kuS
s7cUioAAonFZKPp8asdQpA2QJN+HcRnwpi9T1Vfop8AoUC86whopzXbiKMwEgNp3PZ/B5hB+eRcx
yZyG5xZH4lAllBCT7PrAyhWD15QBcjUg/H/PGoa/BCcsHYyRSuFuD/8nEytjuDHOUgaqza2wcbFY
Ef03xR4BKYxE2Z8LkVI0/RgHdp4UndPUtyLqd1Yn7AWNaNtGqvM0wiEHu5r+2yjYc70Majazz0II
OJ5EzX3YaMY5H+CFLl3VROH4+MfjMXG9y7HTmkvI0zq9LjvutR41MNcZ+SEuLTkJqNiOMVBFmS6R
Jiv5p1AqlRascy31pTS2V5ykx9HRR0chkKy0URug6SrbzFJLzbg+qXw/6APlOrZQPzHRYL2nvxOR
0yTdtvRklkUBkLNw61awNB6yAFowEDQcbrhjH4FJPrW3/9SZSkZyEVV4743+LCwFacB1pf5J2e7g
uKD8q7QM8svnRCjUYHbRSN9jGH7jyN/6uc9vq7BYAzT7jwpbJxpwuTM5audf3WVJ8wxFzH03z0ED
C9VHEnGfeh7mBcD0kERCGMJJHm6l6UvMJFdyHT9fYClz2C9MZlxiA8ybIGySyMMgcutEQx/NbX6W
0i0ulAPwikRxYrMdGC9N0vUoIldgoo/uNyR/6POtv5Q471TbKcfo+4gLFI20SZU5oFEud8Mh32Vw
dF838qlI9B6k9NtHIUAI4RTFSHbYbUZ+msg34ZO7oeo4pyAuNupi2VUleqCuWIBsf33KjBx+jZGE
EaLcSP0MAFciN2CUlaNeDQPyWOr9HVQD64yVpyPHOEHI7XS6eJ61IqSmxP0INjWFsgknnOxL5GvF
8AlMm6+pxzY0/+ldx6i5WPskNORG/P/aX+DtwfbUFZBWPlcjEUvMNqP+ZZuqlNWpdCOmhd/K4FCJ
BwueO4/VJQqwuPYTQG8KJ8ihGtCAd9h9S6esE4Ogw+5NJfFCYO0SdvpbNUZTeFiqmPD5TkAOdJ/u
QF/TMd0eniY2oaAxy9a86m3re78JqD/o7cLSBByHed2oPbYl+onWYt1wAHRJzPWNG6skp/RCM6/Q
tpwcwJ+oYZwoCOKIheEUPgVcqJYWc34g7e0VyBw8A/aoAPCYU5eqdAjii3zhtrGIz7KxGVpv+XNe
S12AI2kuriV1T9S1ZHrrBEqvANYMZrDwkOffLihRn4MKIAAHxaRKZv8MXP0ddZySEpnp8gaqE8dj
EA/WKOtwhT0fa/4IGge5KjxJ6Z93Os6t3Syyefhhy6hpJ9xu/8LhiGAZuHGfCpba37Gfl/VIem+d
7IE4GSUOuB6wPYTFhu9iMj1FiXfQu8JJwZCIf2uSkmLG1xVGvWD9wfcB40eU4MAjKCQwveoPwEzO
sCynR0w1rpkYAaJJ6mOgmJR8W/wG01wzX++4MCZUA6KJLbvsb/7jExGrLegT3yPaMvF4lo+14oL/
uWUBC10ryU2FsJiODtdIPslp1ZGBd470qV3Tpqfa/BoSKluwjUX5OhB+/Ogx450/TnTlxGBWmtCf
QHX8yyRpU++Y3122zntt1pc8T+fSzvtzYfoLPcKA51kLx8YrON/oBPCgPd1Yslf59zMNN5zL582c
U2B3Z24YO6CmIZoIF2X7FxoZHDPa7AlJ7oh6xwRu1h+dCYh7pCvIEAvScOYCtGsHFR9+egk5pmcB
7b66fqMu1/9pDnoljs6KJg1zo69efshNMOJjIeJc13klvGWbDb8Yf8jaLO6WMbPofNs9YSZboM8x
pVaorZkedSTeyo0efkOcdseMuSZ115Cl9sfqfs6BhO9nj3m0tGoNgxP8gWjuc9PUg30BKNha9pnE
xxrzGO5iALbZ42X7zMXDMTt6e1mnR1cOCLva3IjH9hv1dSsKVbBswWHH9/KbAJHN+eO+mK/7fV/y
apqBOQjJxIWI35w2JJQm7akc3H2FCMtqw/pe2hUQDeZNulqOFd5uJuewwZoweMKhZ+GDIa9OWIqp
5ZFtZykX5wsxdT9aeS9aH+WCxi6FtZFYif2fYvYjm68IVK2HlBnRo8zx+pVv+W+ZeOEYWDEoHo4D
zTkxiIVIDBIyRjgRJuh+HKwESd47c5TA5FJ/mNloQbM8MPJPmEy2nSuZe99vuZcggyM2gIM2hI/i
q7OXtlBM/Dx0uGMoQLgcjnCoygKn71fHwfz/GQ6v8Y/CcljBI2+yGO11MeID6ycEXDn8jd72dfEK
ceG3aVgMdGhSE5CfsA8m4gwtGJnw5+imJZUaLbeqEZfXZSWll0xdXDeTLMAeKjfcR/P/jM/UZN9y
Nnqt9ROHLnkU0KTGCQRU5nLE7bnFmfAXiGmzxjWr+ZxDx9cBOe2guD+L9lrxzymOyhohThhY0IHc
NPVYXsisYS/iP9M5U/7c2aKvYftTI2pFX2vc7AJEfbSKIkf3uqjL/MVJSQehVBI0NZPM11XWL+Du
xp6Ep0e5QUIFPR9ja9xuogwr8FB5nNuQKTjGmpHI0jWqfSSPJ+mvNC48yRopOGdQMvvtUv4x0dgv
X7v0I+syq60f5Rd63ty1fvrcS7z9+McAhHnawheYT1t6Jb2rJZHqjlAK9aPQGT8Kk00XtrxfRTf4
UXZn9q/w632ijqYiWfWtS33yE2kX/qTWwxc64eqfUKFb6JvRhCsA9NEZfENo7VBc8nc5rf6p+k4i
aXtqxNmx8/vbaO0x80bjrFNauZt8jO9UyBZU1YPmeffdRUld3OPyfjgvrwQmIHaxGvR6MneZ827/
eXG9WCmFuccnKOk2STEKcAWGEvzSZElD/q9+JtMxwUgHxmXdZLJsFq5PNnySB4gEsA+N87kEJlq4
hZ4QeSaMZtNSv+a6rnVwuoKTPcWYSHeo12R/BdR9o4qWIHe6RSnImB/fwSoyLtyEbsDNb2hbFllR
TlOMlivsUKP7XxmMtjUi7zrBwdWbOr8tcJijycrWoJdPgX9zMGos4TO+6nOGsn0yr8pia0VODIUI
jSK3DFLj7RHo0gCujLObLoSSeeWFNpJr7MMjmBqKK0bfO3geFnvwR/LW++/DnSZLAiEzXLXQOMng
JEJ08j6CDgqDsO2K3zGGBJVzXXdTHes7zzL3U6oGxMiFuvLTdpiioT8j9FMcE/Am2m6twOn36yjd
JCuyC3qmuM7vO+wJ1OfjKy/BDtpzTMT7fFKWBOPDmUfWDGzRVFaM7hLM1wGs+1e7hMQqfEPY/5yz
L9Y5E4yj7264Z4I2pdvetLijrZDnSxPCT1XgimyelR0mTxHpMnalRI4Sv0LEXDfFWSnY3bkzp7l4
Lze7E+yrVzu8UprOzaxf0gGKnqVk2rFhup6tERoEUU9JEAXZvzxfGHg0Ok7NOVQjvVq6IY8N60+N
OkrYI+DJg04IoMF5phXWHFb2vo+o3BSPVzM/H6vV6Pmsh7XIGXLE50zZgrgGnEtR38j8zDjEywHd
WxaG/1Id2+5rw4N/7mWOvVQn0gUHl4nxOI9wCki0aK4FHLVFz6t9rDpJEX2ax00BnK6iRXHJn0On
Q7izW0GxmtwkGfAVCcz4Uy9IDf4bBhVjKLI2gOkgKTnV2p70lct6N8CoWzgt4uC8qqU7C59UidOQ
VDG96Wvepp8q1+Gb0ZiuAePxdqc7umEh9x1MOpuWrTCZiRGc45KDiHqDeJTpoZbF2kmcJjum5L6b
r8TvmFGMOoHjUxzRDl/NeqEQLRA0/JghyoOnXFCsXxBSfwEpMrSSqi/dWBybnUS+MNf1cQMutQq0
4dxu7nbYqzSiz81YUa02FBkuzN+Cd9nM13qZnpSKFSUOSaHNkWqjtmMKDE1OZGnY8qrhdC/zgz4W
IKkEb5895HzTANOtgjVLunLm65vUkpwUN2pUmpaplZu9CCsezOEHMW8jDveomzUansVenO2Y20Qc
2dZaPOV7WI+TQmIRqu9Wlv2TK3OTVohFCwg1sjjoMgEYe4Nynup+aR460rxhqY/21+SPPVn+UJx0
DxvEAkrFFIn3mIc7eRAV+oK3R5wbEhz5Sq2dNlFa/ho4AdBLUhIuSK/addPHz2xUv6p+LcJFh2Sv
MWgGj9T3tsdqkkTabn06ZB0Q3shqt8RB30lB5OCnPNODWHeXP6T7jGggg5XrD6lWSMqZ2JTw1oZ/
y/uLXHthE3NTi2Ed3QF9BeKYWQ2H8sBwByR1WfU6riXlgiCp1OWe+QV4zg/DwS5IsspHB1gEWUkR
ZCNPck0DUTzY/eSiTVUhxjDsDn4j7cwAU1uWy6CVFGCH9kC17+QDBVJ4/PHwjZju61u9IJrN908j
/3bEQLpNM3Sy99Pq5Zuhxac+AhCP2VvhD1TRYk4UV2cqq0emqUgMd1ZuB7hlFuRMRlEOtAZWdEBY
0lfMv85DUpSN5NiNjI4HtlwsmT0EfwmtRpPLI11fL5Q448/2XAsdkofBS0Vrj2siYL5pu082Wr88
ra+en6K/hhrh/XdZJhIiAyaeKfSYfruGp3B/Iizh3MvQ3MqnvYCIOSsxpJNU78lMOxmuijtVd30b
pHknoaTsWBC9TbsAsfIS6qMbwH619i+2oqPZCdJI+eAdD14FIgvWoZ0XMyYtfcmvgg4MjSjU5wA2
c25YkG7LY6z8nIe4iHBoSZA0wSQ9Bpj1Lt2dKRix59ZuMjXz+Mr9AjTy8WGZkdjEJhNRjg++XqHm
Z1lS2NcRsiUu9odzr+n3L4t0eltQOJYt+lW/Be4TLhCdnuuItWkXpM2iQ/9Qcq4sJ4JA6jl9NDNq
2neaBXzbGZT/k7tL/ZO6diHRFk1A02r9CGoyZLRridrGqpe6dJs1W56Vys+0i0mxxQArZ2cISIi0
+WQKKnOJNiEtoqfmsvMJlJi6kaagjrFGcp/aTrd3QYvgCzCqz7g4Q04pbw9gXUDScn1228b53Ju5
FrpiBiOswX8xO9xewmaEgP6ymdRPlK7vbGVnd8wDrAZ86srXzhD8yDNuwl+Q0Ng/RsNzYCCKbaO2
R3viQ+6QiAuy6iDLPaO3HXfdP4Bamgpgra9vPNuMces6KBJ6+nuBHlqDcx18WEU1Ul/dh0gRY5Wa
s5s/HsXyc6s26Vj4WDfR5Y0ei0RcrqNwP277cCkgfiauaVQt0i8Tcw3DiJ2qj8+3l19Dus1CyL5l
7ZukSarnL+uDv/HYSVu0Dw4Dpd2pMbkSQvGwmn8502jH8kNM+q0Ox3trw+GiTb/yrIWqQVRD5j+M
Slvt2ZFNw6qcqRfDE6wu6j3fBFsac3HXwyskKycQkH4WJNGET0gnd60SEAoDSGC/twYdoSE2yZUi
XJzYV7sFuwM1BSJPcM1TOJ20lp3MUprWYAJBV23apfgBv8X1pn6Plf9sXHhCE//wi2bPdv/jW730
Xy1c4k/A5CZRj2YES4vRntkP7go48I2pbVeTnqJVvfXgWN1RB2W+3hEt6jkOfxEn7fsxNLAkgfQ+
71GlExnKYQMtROkJxHG7y1a06SI3WSgRlD9nMnNgnIoO5G9BDnMHHnw2gwDRuEDHW33LT1Mq3OyZ
Iu3hUXOO6rFGQdQv72JRUYGIfw1zf+fadoXs07o9VxIERpz7oOCjvW6BC5U9f+kW47N6BjvGergu
zh/zNQIBS66TfRXoM4aX+rydOw6/oXZoNOdGCyCmjS+ANDaH29w4JHDBRrhMPCU/N/sXSGpyKaVK
YhPefD6AHc1HLJEOR3FK4p2aHubJWIm3iVD8giUrKfIkeGuiBnxLAae0uZZ4E1VZ/5ddbjHp2ShL
SLCnQuNvUsJfiqDbuiCjJE5nI6+GiHgG+pI/SQ6xUi9GFjswMILG7wdJb+NkT8JuIOYAyWWMVtIr
u4O0Lod0KLpEwyV+IsRMYlOOiNyxY+dQxZSnOHEidIpJ+KlG2OlpsphC+xl6HpFV0AWt50+E6tv+
1VrOuA45RKW9wsrw3JirHMPmUQwMQZrrq8iM2Go0R7ZCc222UEf52zwON+iHlh3BJERTM+FD00ZU
jCbR9qVCrYkB43rw1IhR6+azsPihYghTIOKLYw/gJGZhYENmw+1jZlA1J4O6H/Lp6NUjO0qr6+Vs
mhUxXIT6UBXSXCVTZNo9zw3E1o0V1nHsdE8C4mTMzMICaAeyw033YxLqMyoSyxfarRLpv5uLSHxV
Z5PKbn0JnVGJYUlLFerzDOCgZci3tWspK+mvLg4/oTyB6KFPczeQGThUVcwiy5khHrgGNgGSTGaV
9W1HLRZmXVmET6M6WJwO9Qa8wX+l7hER00G5T8R7NewR0O7dw4MOCYROJQEcZU+qoZxmJ/q7MBJ/
B/3nzMqRwZvrUA8BsHDE7F3+xmGbX9oVKV8GYX+5tr2pixAoaFCb2bcwGbJYVytbweGbGXuBvP8j
NKCQuXHmvYFvfRPM65TnUWLHbP3PesUL1ImDxvBocVeB73gMqgLko6lBlsCmtO/hUor3eDf9lL9k
Bj+wUenYlqPLm+2Qz1BybnDEkeXabZ8DJs6oeKTAgQOwRR8NxmlINCtuT224MEho3MABMPbIoSTW
RF8tTOJ0rhGGHBQy/KQm7hQaWFMeUF/+v845e25xFp6ucRQOI33V1E6ggvsIcXVu3RXpHXk2yQDr
EYUWouHd8e9L13/i/wg2JOH4rgGCdS4glc+BhsVsN/qYRbN+m7bT8Bh/wfCMaLabp8vB94P49Vdk
JvK74AhN+HRyk8j/49ZcU7NQbzMT2R51MrN8VcDncljfIraTPXKcGS+YwRuk6/HLmHTYPBzueLUB
nB9dR+lzY5LTlPhrM7PI0lVgT8kISr1q68vK+3vr2YOL58sKuhpMNH7QGSNkemabIRvlaISEWRKF
asFOUB9cICgIuRFuzVHT1RDvn0RIAY+OF4glcV1WdNFOS697r4qSQuFTxfXYLUmmbZtHi7jeEde1
9TDMI30vGU93C5TkE97uunVOY2fNqntx0uxujjkbQjHhJrKCZTPLyMhHtAeMqVbiw3zge00Qnj3h
QJ9QjAy82DpzPlCNt2zyURt3mQutaMwnonvBITymbJ0PTIdUkRhyRiFpnDgv1njasg3W1TgeaRCi
5cqUuS1m9/yB6/xmg6VFZaHxu+lVDWov9GE3QItKYyF75bE4qt1o8WtCsTddoTC+KAQ8bn3GXEC7
XxwiengPneV0VDVDn90KOKzuSJAxdwXYRWb3NVttRuDXauaPEXQeb5EdTybc93+hbr5N0qu3Ft8/
WG6wLeoqmH8TDGKP66JE5+e4dSh8LTIlGv0F8CvoS7ZrOLOcF9gHsrYCE6XURBj+AzpfVaASefYi
yIGYncptYnslv8siK1KQ4cBDAWiGf9gi8SixmAwDZmqUT1DoO0KtSycokSAFWRWb6jqIcLmIw0E7
bTrGNumAr0SH63YXPpBrnXLbXiTExIlRnfOAGyxlPgOAXQFRmazlNGu1kfdtCsqBFjGSAYO/SVgR
Z8nIpTrXjFrfvzH6a2mIGvB13aKt36rfaeXarcKvFH5IK5PJ0ioD+QifqMP7a2527SKE2YVB3z2e
cAH79P0pVkBDlyr8ciMUMHfw1KBOVuoutE1VOxmG5yMFuj34uw5JBueDVeGl8z4dLyTj/NqID9GG
ABefWUTsBXls/ATlG/VWpWOrDNfq5V1qf+sNVGS8Kuvaj86CahrtH24L2kZylQuo+B3O4Srxx7PO
0fjwqDVVsaO7+0Os5wsNKYiDRndSpUMvLSB4eI/AFMGynROSQKAgiOY9+hUIvYZD5u23f3/iG8Rc
qPtn4rF6X2ZtqBHpWzROyGBP4RB3nf9cuWAHowQzZzBM0iltv0fwWLaKsRSjqWcgk7QDs3xybeZL
+lTonCJwQthyGQOXxIX6iM4Itw1HE7ClZWELJHt9CFq2/QJO1sdikaZs/w3+gzV5PtKTUTyE7sRX
YjDzrxQsLczy9+FKddbqRd9WuN2O+KwHKgk1BeIHzaKl6NnQ169CX2vNKBIjlpmnd40+DSMqsKUq
GZZwulhJt8lTqdVIZUjNr3GcXGTh/ky13EdT1Y12ict0IYuJNEDefnPx1JQaKPq5OucOD+E5OJRX
aexunfo9GuGik28lf4uqB842LPLT3g+a39vAvxVpoL6wM3u52o5apxVP2Eoh6TSndGk4WbECmuJQ
H+hNsjt5UzhVn7Lv4ulryQfDSHyt3NWqxc2LCP6klKqQzU2bAGQtZV+PRhqozgm4UJ/Z+k9OJiul
GNO5d9KIc3QiXI24u4vIVhIcSt3GBqH6x2vPmtbQlpM4meV5Ek3bJXZY1XAKth5LTBBVo17aCUdr
uriqDrTW7dwmXbMaiamQ6HurkVhwushDikCMKRkXOPwbG3eOJmn9p6tv/PCCmLZLICpbv4fwA0+n
21A9S7oAk3h9TdKBpCYop3f2oRBy+VS67ZsGbcimpo/NDzvIh0XD6uCeHs+rQpxFqKUO8jx3zHN2
OM+TLznfXSRFBNiKZ1OqG7fBTYXJGJo0LBwJDC/1+1s1SpKRNShaRMYfCURLLRC8IS+pq+3kFHWS
jcCXDCXaZH0rLlSc/xUFbSjZjW4y0b2zpewQC6y9H1Iepz9Z0DftUY/S24c6OXOSUg/I8zMxjfgr
gM2KO77J1eb5vhFoL4lWcEtp4JQtgH6Be89DPMRryTJwKSyHd3X+etsnsb47z43vCK6FbgB++RNd
2MqnB6PDoSVvgzBibSp4sZANvDyRVjhzVnIyrBPuxtuUZxMvE7d+HuMy8vVK1yApUiqpDaWw67qD
7VbJVveILQH/jei0n+eYxmZfqg9pK2PTQeJvuKRXfVSe8YV4ZvzWlHrihT9iqMPwgZhnCEQOuj+V
7JXyUm/bq+OiTmS6I2WYq2AsL9oVkVFXrzgeweQd/RazdJp01Vv515ppvox4IG6+MK+Ryjn7G+S+
uN92gR2Bi9Oo5xOWCqkejCUa6YH33WhWE2buPN84YIksMJktzDRIxlslvdD3aMXkut3mViPYSbKz
3ZfGdYXx7BFiKYvJwcuajuJFtn0rhnDVoIt/4Rynq8rCyv6aDGLcV/0QTL58zTPihtGrOKXHIk8J
ac/P0ZuHjGX8GjCEYZpV3O5zups3FG8uzEov/thrIS02kVc1xKy1SFE1LnNz4X2vhx1BT0r3jlWs
++DOYDl2rXSezFh3aEN+fnSVp8Ke0eHE1eQ/wnUNKnhe8L3o6YOaD5izaI+XjPncc3ElEKnhJKoE
11xpwTlo5Jny/1/bBgEwF18yGc1qGy5t2fdI/XrOO/V70HkltEC4hCnEhN5PWp2AP+dig5KofChO
0Gfo7kP6XxdZKe6hSdJlLOWyqv8qJT7v8hm/vqruicTdBNWYhXzA+7TG3WwsMGk2Vcjs38lCGobG
M8NHDVD/mbnoPG117n9mslG+xJS6UgPdT4xrHedDoE+kGQsIan6h0n9iZFDJmoRHT7TKMYp5K+g4
Eb7J0qTUICauZsZAG8oY0ASFiYr4WSJP8iRrhPeUgc1Gg4OGMRZ33Po8VeEGfNRNFHq2KAcI3+D9
yEdgsQEA7ViduJ3Yf1naUzmuzI7ivwRKbpKSDWiuumuMQgf5rbh3uS2gdr6EdR1rhXxCDlQ4Qvfs
k0BzGbtazeBQ2UhL1hq/6ign0PfFJzUeJBEeWfvGM/Fuy3NAicrbYKQHx2lh3r1f7u/FOGOlIwAJ
xXXpnd5+c7/6z0AuvKB5pORxxzbct+/7LMDqzlncdGuFlOUtQM87a0yVT5vA9o9/Vp0uXR/HC5LD
cgsnjYAcKXxwC6Bb8qZfY3G0v/xpjbh5xzXtL1lovu9J7C3N7NO6JjQv8LZ6dnOtWspC7NqiR0QJ
tCeeP5xxlch1aGtJZ0NykXERDn18L1ipbGJECs6AAsdV1muAycX2xIDnOUeIBlqV5kVzitcBPxfF
NFIY6Jxg/saIDCG0wDFFjVS3IcHCCYYcCZbMwbB2TN94EFANxSrJ5SNN5ozIzICl5SmTcwftdvj+
CEKnqvzf3Timhf6315SgXKcy9J+uKVhDEMNq55rP/is96cXXfRQ0jGQLh6lbwR4xvzpDZnNWyJjp
gZbASW6byzaShB4vjJlF2Qsm5wX33Sw/8dZ6UHY1iHL9spGBJswRHf6kuSz2Cm4XWcHxWKXAAXEv
Fv523JteB7Lpr8jLtDVeZTPAa4fGOjjuggYAojufPYNjyaVkLisPRKYwbjmo804zJ7XFRsLzCGZ1
8IOE0xRDltcavhrJ5TAVhy6vY4/L58oapUmbtTUbsoE4K3+c4ioOBC28aJ0wNA2p+rlyyvYUsP/U
8cdAt/+3cc3fz2HKh5Sv8iL/TeVBoS+OBU0j4oRUun9yIHsGKfITae3YR9J4ejEP3zOwVc1iy3RY
MEGWiEfxUTgQeNC6Z9sIcOu5x0stcgS6C+opWVeWYODbNrPrieDn/RZk2qhcl4kDKBiFRSgOiw+I
KW3yOzRc6DfJQAmqlwXWKc8g1Z/+XGSAy0YqwtIs1d9kb3O3Mf/695hJv7xJcKBxDFz8x9tze1FN
rS2j2XkDy8awNlUihI4kXCorMZOQJIlLc0mj3bLpVbDd87kUt5a6mIp6fB6wt4zvkEDKrNpURX0J
ACBPvxsUUqhP4MlbqrBYKzZKIbEhZ76gTgE4npWFD05G9qXXbe23KROuGdbGsK34wgDh0K9vvg/H
LKk6V+NSVhwM8m42DVMkRrxAF98142pLb61Ft2Iw5VT+X3VafDr6tdil5VL15A5cTZzDD+zrC4yd
2jopS0sI1a7PVFHnt+PjnfwV61LXxA80B6ZUG1peJfcb6yCC8MeLyMZQ3wyzUwxV1XwmD71l75UC
+Kba3tArw5DPdx2trl+h1OL/t2caLl8EGroobDGXDLUqZ97Nh0kbxguciop71LzskIoASCXdbGbC
a452xA1GLGWuuLVC/NvabndvxEgZM/ZUByL0smazzFPF10JrO74ZFsjaCkp0YBn2urRUgEQQ2fiA
94dZTW8ZO9rl37at1pn1TAGeYf90diwCOWKavYC4r/QAfxbfg96pbQeQCz4chsT/GvCmXO6WQpDk
LuQbaCIq+OTBPfVoggvTHKKKueRhtKjFMy65kQMeGHbO1/jk2yPnIAjHUOWDvGWKgKWCSbh/JPQb
maM4XnU+lundNr0vWjKi0c+9yhqAmyvqIOp6WTCuIoiNDl4wWdikI1s959Zup8KVlECylXA63alL
Xhd2SaOY7v+vVofQCEVD9cC1PbSpjGXDDGj6dfl+Bvn+DyNMKf1yljXkJIZrmCFT4ckgSQiAOZOs
6hp6lvaOZBE53/M4LrOPpHelNRffmNAkA5IREZgC4u7XgW3jUP253LIp8fbPh50nZbtLGpqBJy1g
zxmAf6pG7odd3YM0sfHPdEhcP9+jiLJCe4l1y4KbHPzu0YE8pBL+HrhroqvCYNP8Yq40TU9tNMeW
q7z8hSjl+O8vCrP2voDgNOOnUUONydqveHUyIj++W3ge6xOl+GksMtWGRA7FY6XPQb1dzGoFsGOo
oQYGpABW6WT4YlVWSvM2m25qiGXkUPpRByV/KScYVvtJjdDidAGAvKcqIEu7NiB8gzZJTmb1qE0a
IUdXx0m/SBpfz9LGNkvRdwJNDUe0NqMD05jjeunchjen1qgSUHOuz7CGyMi4G7Ul2OPWn1VyrfUF
xJiU0PAEGKWuKylIzYkBYkXb4WCTt9Q81XKkPjOo4dbTg9uRkeyxX26LGnJJtAVEGXzmKTCk/ig0
jlj/0PhB69HQLqcJQpRTm1FWJy/RYyM1RYDXUgDyc7FjokmqO/k1i3UvkNwuHkbcJcvnaEO6uk0T
m72jzxFqX4NJPxZ567Rv3Bhfa96zifQErUl/p8vCclVRTaxgSyerZJBUhoAVu/Vs0U9SOUcuZMzn
VzCKVvz8329rX56xhyVn4uYeg+IZuD2t1WKtYfiupLZ8yT/a8Mbe3CDrNOCeuGqpc1w2yydUqxzE
gSBxRV90JLc/wyU8AfFv9QTJt3dZ6+/MlQCo1juSzQvwGoMQsl82Lp1hKoYetGZfAQtKhB3oqQBC
WKUTY1oNnY0xT9OvZtwj4E26+l+n/wfgDt2HrlImKd/sPhxus6PKORNV3prKJQsUg0atKd+4vPZX
2w7JHsmjTxjpVxx4GVSilf2INvORyBqCDNKvxPT0WCfWDk7Y+K4Dma0qSI6xxZOE7hIr4BScf4E4
scrj2Xk8r/Nb3wRYl1cF4UHT+jsbGpFcTWgjVPJMQqJXc3kTvudEyhj7Mahua0yULNKBpp9m9n06
rBQ5SYcRqwbtZ+4v7EHa5XuYk8vmlwt2YMaMiWZuZjYsz+fT/4SEfyLK5Vl8nWcg/1e7uCWkeIST
evS4eerI/EYBOzCgj8LiimztmtXiVrfCICy1hEuySPx7v3U5oIjliK0vRw1UOsZ/KjhtF7jHY8Py
J3jjVJsvkJuLBTNpYpCduG9Mq9EgeGEU03XDoYqd4an7mVMJWgTX3/BwJBj4sGvj77CMGdgNKFOW
6vWHBYva2M49dDenevIkQqeCvywoLevZGv71EiBvVJRdXEe8526+Umyx2gWLrbontiC19QuhQHhK
35TLdheQasUvSTgqGTLNyBj8oT+9B6RucBalj3VRAHA2oFpn4EndDJknQzn2BRo3vsvvN21HTLHO
o3jQq7KiYnQU9DcMcC8B+j2Og4d3MsZjhDAlvbZ61zhuDORzfz3tsxdeZeWhUVZebvX9xqZWWWzZ
NY875kB+y4e1Sf8S5lrANuQCR+s9ZvkQCZavjH+jVVAfooDfYFKbsl14mu2G3LtaZ5RnaNLoNUME
1T1FgQUBTTzUQpPCNISZagf5ZTTrE+fuaVC7ZJAs58Csu6zpG7I2KCnKdHgnSg+RH4mo9ZLG18l2
6B+5HAYSaz0YP2dzv0Iw1721lMPPgjGUgdi896h91J0yA9KHdQPbJa0xD5ZttPMzcyfCIbISL186
SosjiMK4usydtX2cq4qiQTgzKzB1lQ/WUpaLWHmRXjCUupjrOhicFIzb5KbApHKyZ/QfKxtRM9N9
kFG9ooXEPYh4/mSLbaPky5od+xSEp6oMLy//OEoXEM6ITGMlC/2FdGhIKZFZgCFf5AIXbtnHvM8G
uPoWrxdDmHdKTyBoSwANhf+Oj+UUT9nNqoaeoIKBXo5uMVILPQ1fjkpmObD9odEOW05qFvd6COHP
40AJFWOd0+TOWxHdno0YM6NdeBuHL8v59SpWPsrNpMmrW/VDJ+Nl01ukZxg9Ebq908jN/3q9l79/
lu7GvU4VefDTiYFfMnjcPNYYuXCLxic4ezCAkT+rn/Ne6yYLXIghXPGRXnIEC0o8sevUpI50j4gG
owQoy3JMbiWPxtxc8u5asFwrkR7/w9w+e8tqt0GvYU8U6Yg56xfc413rj1SKjyQ8AJEVEp4qSm+m
MaiPU1bSUHXLMvKMrPRSRSMiKpDQWCDWZKv4ZLE/imIo58dTuUcf9R5H4Wj3G6HTn3q1pQjmChf1
vdVfgIivnGU5mC50uDJbA///vdf9E6KmXkMMyGSGkl/7G/PAKUKlkyf6W/tzzHSzw4/1cKz31Nnf
6dmU3AR41I1ZYt3rbTCQyRuY/R5SZVzgrqgsTqqjTQMkKYfqVc5pETTlYRAV8W0p+AV8PDycJeSl
QHVqtfcc3zSrbmPpWHfP0Z+OSL4a2e8UxbcTnG8MF3KlI4ncPzuDy9GD5aIcGl4Ceq/dhPY7KdeX
/+s6ZtUKQEZzZiOeQefEDjnQBzqFUeqtSWeugZmGXbj8ULqFrLDXFV4E1Nm0NUdZw+D2b80+pm7Q
1v0ENeEOrIGhuXl1Q1ad4sII1dxUUhfTk2zf7H1UuN0fSZDEOTgR7GJh4ZV87SerEeqcElG3kfPj
cSF5v9UFy/sVlhiDVudeuPb/+X0NGX7H7LPhNYI7EkZb3psnxgPWkOdXjIwxGL/1jutzRlPFX+1u
l6STMiGGOoe3MueDD7byXBSQ/BmDWpoBPOUfl0ehmeV9amcxH0cE3D7bGEQH3nE2Z7Ppl1bpkanA
hPc3WbLYevXl9wsodOoJzoNDKNPO9LUL24hHZha+6GPMxiDlz+uzBq9APg4nLmYCTYhFO79uTjKg
9uXCZNgSHdX+5PthG0raZWNq2uebFkkKDC5wmHcCoP7Gi21cz92ZIUrdRtDMIOn082zOd1FvDUVP
t5gtawvkpQxFzK4adz+tc6mQ8tf/Z8BrpWImVcy8co4R85cVvdX+tVdrO8DpX6rN1Cw2gvq3yl0H
zQupZ3JB/N2lQgmLtLpexntewRZZi3/Ft2OhTezW2lM5YRoOD9vwBFga6aWH/4s+Sp0hoPtBkAAb
Ppnf1FNU1ZF+yXn9IqakfU5/zvRCouTl6GpPOWoyteffSKir7UBi5sAzMPvtzsCDtAt/tP4EFQKN
d9zIMZ2MUSvMcbAIvmDuHrtLMhgDJm5UEUdC2+sfYeq7xjqxvKcU1eRMZFX6b2aNaRGPC6PlTFah
3uIepCx5/Pbq09yoMK4pwKSXuP7iCsZ/kd87ZO0hcud8cB0sPP25+MonrZZRHLkDPwR2qi3N0IeL
EoX17Dw4nm5uOqzRqtggEpgpTfpQ96RAps/iqU19TxHolgrC6ojRA7U5OdPCI7jQtQX52r2Rpe5V
2PcUp9j08u/KABvcWszLWNrpfxsMVCjymd86vpm4fTrH5kBp50FdEkj1rmpFaPmy9KmFd76xpEAs
+6WxRTCyKDgrAwfBfHwpHMifpWGvj0c30PJ1CHzxg3c2J2GIn11eh3vxdmG4ObQmqWmZ4HK93OaX
fANmFFwRaIPXg4KzUgDBZjIPOLSqDIxsq5giGO914DkFsfQF4DeeetxLed7Qo+k2GX8R40CxiD+s
fKjfj/fdU35llUWcIURaPCYY/TCsE4gIHfOeluu2Sy1xu192/eGlLn0ILSPcSaPEPgEo9trDySPn
YaLm7oiwtSzaV029ZuOXmGIAABO2Yc70zid0gGtSML9KH9BgwERicKoeHUjIXYcZtU3Nb8cah6Ae
kisD7FeCztKWFXc4h+Vps6MgnrvpRCnq1dbeN6QT2fQXqlucxj5Aif1oKKX8LYWg8Nkw2/tSm7Dq
m+KUJUoLB848C3E5f0SBjTTljLQB7awN488J1jecQwuumUWFzHaE3T4fmXhO4Qavu12Dy0yxgHKw
KaZLYx1LMis/AAR1UiCSAJQeEsHSiO7fSHXYSo9VuQcnZ9acyAN56KKVEsZAuHzMomSXq+nHoCQ3
BqjbPqrCuDi3vOCsPHXT9avJt1InqhdQ3XP32a0GbJ7SI7QoKvuoycsWH+1ywcTUP0mQmFa5EMHk
LKfSVsp0Zl5pO0AXu0xLWrV7wAik1GgQWy5oWEo3TlFArQasKX/b8OIgt0EWqKaIsALZdTPKQpNg
LmUnTvvQAM3kv4gMHH3ufYkPX6KloAxLaWf0i+29TgpdOMJ6KttrCPK9cS7+E+kM8GH/uNbhshez
oq7g+wSTGnXKrNlczBSLTRYhSuM1kLvmeFaUlsfY/5V8m2cMBoUvD7rZlur0I8x13wNfrg7TDGWi
7OvKzolPRIRRb5esGo1pwgjz34ecrIFevlqHPLR6drcjKk7aDvHULQhBPSH6kSpPMsTHqRYtRQ1z
qSgfj20zg/tPWY5FRMNXyw5JVFVs/7Ebo/K1t/5ordBhfseP6HSXjWOk/YhTtJY75eppN3HXTwnr
bgfwsbkk16Lz9RJoaevpObZPVUzJumcfrBzmc9hnW92zgAcJKg7jdFpRMOENQlUpUXW4dx6foVRh
bLmInQvjUgu/PK8ZYEFJ8dwILQulHASa6wm5xg2LRsF93yLDYMzkZtE/Uru3rDFI8dBNbwqLv6+Y
G2a00rr7gFVJH+knxCi3mPN9aYYCgkV/nQZ3jSZlpMaW2qXYlW8dyJY9eZyfD6QBrR6JZjiuxfEg
TMR7ucSTwEpmE5lRsj9RLe2QgdnJP4u9GWvIu6CJuYYAvRRs9KULrLS0UledBz0FBBOsSnF1DFSd
YrWCB1idUTBjc3W67/DR47lrCjPstkvQvJJxzk+wHUNfGexiYDOg8E/RDsKP1WJUTDbIePG3CttX
oXIAaZObmCfV71mgULdkd3DH7GgjTpNXpNClfR2ayhkxtW4yXLtVzoopggI5u6DVbsRNBEgZhQYz
LvLLeSCapGSsOpi+baXTXM8TlYH2hw64nj25+MBsCRcjM71bwbKwnc0SNoHFx5KFcwo2lzU8SLQN
D7A/UJ+SvMzfGBMz3PBYRdMIk5FjgqU0TDrZo/WmV3N7ry5/Hi+ObV5UsOt8DhiT4Bf8JYZc5bS1
Mbd0UKU0zAjf0BO9F26W1rChYEdSWb5sddPnAFFjEYkldAMbFSRxyPOHIFtHJWjENByVbkXwiscg
Pfq1JT4wfaEhbQKK/9PG14MmVsfzPfqbIMAPvS8WkmG/q9Vk09ctErljZUfw7H1uc2OH8QazRJfR
XOqXA1Pkxw4GUzALCFEUDk0bfySSOp+s+4kn8tjPMvqcj2xqTwhaE3+CaeqipExuty6Al9Vs5o5C
b61pX0NBjTZbH86ZMJlQDLx2mLKCu4Q6hM73EJqVeD88Y5SRKTrPQkvv2qrXVx6DMjFbmSRNdhBD
gfL6FuXCTDTXd0PeE/UwSxLV7zsGfoGJT09s49tJUXx0t6+jiiocOAk3DcFXv0/pNTt0ek/13iHB
ZbUbeuaXcty1oJWtoNMMkINLd+oCV6LuLcrCqOP+MYos9P9vuAMPFKMB/3mptitU5gqthd7CJcut
RERIBLGfDbAxp4CfyYjlsfGQaV7jlnokfJlGcwR8CuxW/o9GvXdKUrrNmjpvIRs1BB+a0T1VTXhq
7opL/f6CVNTx3Hg2RAG6hIEAQYyD6RCcu/8IjFaZzGVjzHlhRwJQznQLvwRcOWcjtAVgsRjiI1Ut
des3GLmGJQE5PMs2KnjdP92XYCSWqoFhD+fIbOika7FipTk82tEwGbRB3Rgc11BBpSyP6j4vYX/N
f0oZ7zCO4gZdq2CI9XMOElutNHlQdAD2AKQ36WYyuazcUrwHaYchcdfKjI1A3kWbUnhfBrjJL17E
0IWGa4vSGcQkPc8mOYXBM71nWPH2w7O0JfQUCiRwH+fYnoidvAAlwgxjr3soKct05CgopdIZJh7p
pNua4ZVjmuAqzyb+qV0E8eOwhqiYLGLr+nMpBEEvJPLFI19p2SXQa+uIFZJZhXPG/tIcg+feU0it
zpPLxRiloNAURwsLkf/p3eic8J1NMjON8K1qow7KPW8wUU9lvse5rEcVQ445ILqYT1kUBqowvOD3
29guGJiivImZNGGR2ENhOKABoHg0l/CJtw7EM6+m9zf+/RbpxhAWWuOs2JIKj2qxhrCoBwmRNs5X
K6vp/Z2ZsHmFFqopxYSIlOMQr26DDRM1M8/fSMeQF7oBUWMo7ORxi30icGRKxb+U1c7iVDC+kUbh
aityz7YT89+b/k7rpg+gD65qPC/ytoG+P3rjuiWcCKADbkDy2jhgpr3vWjgsGYo7KfQbwPbIQ35G
WtOW7/CMGe0sUMI7RijgF2aUuBKMj0UG4FSB2sZiek4HsZArOcTYhVAeLmjUnHPs7QVRmG2OqAce
d0EONpx2Tio2YImiLHuAa6kIco9uDjP9IOWEsxF0BipsxXNZuwKsqYt/OrZH62LjIT+McK1HNx1h
NRwjWwWY8ThS9hXcoebBu9ZJV1cx0PSI1gSwIDMW+0/rz8RLmHz6Ic+0WjfmsJY5OF15LWdx4t78
9xCtMrLniIxki1t3NArB+4U+C21+ytcSrgesUttChzqLGsfXmVfxpWl8RRgN3ZJavax13BCPfL1e
/XwNp97wHnPdNzaqdWJYal+HBZ2BbBb5b+djHMwkwkyP4eF8XyzLGkT9gbFoTntReCjgB+MtXCvS
YA0/PP+6ZVGCAIUjRvsRvLUnU7Z14ymsV65ZUNGpzpLqpeUb3IJk+avfiqgGDsS6h4AEdwXA1hWS
USeLd785mDlMl9oZ7xNUkRl7ZXub85nGafwnkqUbN28WH7xWqDY3bw+MtU+xJggn+T3XLTH3aM0/
6ZTQilqQzGWz5ZJBZVI8rNJgZzgY9c/Rd8zDvJsS5HfRVabzlILEgVgiY5ZyEvBFtdLWeTa/ecNe
I7FUcmB9bbMf0MkSLbJBIpRuALf/NlDV29YLkepNwSlA1giPJrDkL0sRwHxCIZ5bVYLdcu/I+SKG
nCmY/OwuP8Qi3hAzIlx5y0KeKqdYFpj4G4pMSUmCuoHs0/n8viw6DzR8RPXNqWhuLq3yPVNh4luu
WRsG4x8bhvQquhvlo7GqvhQWzXQ9zN93K3l63yyRBWXdWyRp7Bq0UGPI1gShUy4Sgf/d06KrcPyM
kHYuE9M38lLlkKS6eVd7KE8p5jJECCf5+ttCrd8IaOdI8KJq2wnjnZjPUVi6Oqzk5WEMbWQLYhgS
egAO2Sm0zyrfTigI0y7JW1NZe8msFa1BAM/8Zz5oWE7uV6CKu7OyFqUkkJFATpvOMHVxci/uZL28
SURfSINTjS8zD+5NmtC7NaFmMANuBaglZtxa23175INgXq57vkSuV3WBaUfqKoXcts68i7rPeMWd
tj4zE1pX4LzJb7q+LNr134JoirakOv7rcR14KkMfzOBHq4pojw/QqIWwqx8NhbxeFTbIUlWG7vv4
IEFUkB7ilXYjFFiljSgS7NdlHdMu1vOSwsfC/cXN/24+Uyt1IPxst4H+2MdQEBz8SdtYrZa3dJK5
cJiYoRsmMYJ2XNBcjNNgF3nddEllL/nDA91mBPgMLDBAi69hcXB839rEL/+UBNLOMgeqh/QX4h8C
X3xlw+Tsr/SHE0ccdPilyT0QVgj+5QOOmOiPCAebDoJ6VXdE1g5ivlVaWNwW4kc1OhKVscatSEsl
g8DeyJQ5wKmtfVrWWp+hs37le80LIuNqwvPQ5yYIB4x5FsSK50Sq5Vk5FnKv47/8A00Ztycpbq1l
NG72IYdDpupOFPAqxDDto8XgFgsFE0jpfufhVOyLv/zunqk5pHhHy5VBCTm6XtCmDT4OZI0xbozH
cq5kYvVyrGnFAeldSUBqLdl9GkMX5U7403qwsBNdw2Lg94RY7KvDiyQ6bAK4cq5b6ENes4OaCkR5
66+aoDq78xhkgeWmV0+VCpOvVBjt9KCo+qWY44Gruuv2X0IT5JTDMGnMAE1tJEcvme+TQo3EK+Tg
T2+pbDzIlRemxi7hqNiPnB1sqSLLA3IyXsj9uVPKTX2YKS9ZUdMQd+OSOH162cEngq1ni4wwWz4X
5ZlkJHGFkn5rPYEqC5cArJEDLt+2wEh2a1Ek/fNX9zMtkqon5IARSy83yN7TyFvdCeeLL+YFIdmZ
ztcpuXrBSvNzfl5loqBB/UlqiZnAXSW83ZOZHb85b957o/+A6Uh0OMYUxVIdLbXizqr2sEAdffWC
xo/X042SF/1SmLFzt8PtovpppS5TF9UD+RaKbok0YXyK3pvkh0wPzEg0sOUH1FvEq8AoqQ+yzDFI
x/Ed4xmujhGu+a44ptDuW9N/3cCmMRcLtMPnm0m71ilNbtD3Yqqq/iokm1V8hZ1UkqqqShEwLulH
juwpvjUiI8htDdI2jxGVgKq8Oh9spf0caTQsBGT0BMeKn6WLy3rc9RLm42qi99Hg3yWOmkmqB4YO
2iWrbg4N+eOkTRjJ7pQB+eisTeZVO9oUActs3ijrCBR1EN5LyR8PEIPM7VXysx+xyVPTyDWqJ1HE
CSA00NHoIBVXStgbVISAP5Nc3t9+20dTTfNH4VJxlEzc4nokcPCyAqqJBhS4Xjn/865x12fgj6lj
1VH7pt7OGEwiD5Df2rgg8yudwOVCiE5voHkCfZuTdP2++iwxP9SnRaugLAnCmWK8rqybCjKV1tWx
upEtTgpL/U8Jol8BBiPRNAicoBIiR/G5OWWaG8Kf/HiD/hsLg2RKJMpI5SRTsYVAeAWOfZBk25RG
E7+6KsI3h1jBfLGB4DZC8ipd/dRykMm+hnxgcjxMrvoPZi+7O1nPutQcmwMY90VwbbgTRFQdt5Bc
RchBcSd8i5IInOfFe10DiF1acBWyV6Cki37FIaIozQl2aRAh8Nt4TttLooLBvCIDXXzt1sNjVCr+
qgT5pEk7l1DB0i2gb1jHUiVEzwiFE5K1tcu4A7eQyTV3gx61dIVWinzpx1PSiVbkw3eDxXcZQa+x
a//MCAxB4PcmdhDPg1YXdRjzVxEdOoKyz2+DifU5cIxFXeoQEgyeZfA2Zd2Z5RYkK2+oZaAfSSur
NCRz6buSpn4+HOAAe8Jof2Ga+7TyIWrZMAbMCeUlGyC+2M71u79QFertxSjOdq04JrXLUz5No/lr
zyamM7Unb4lzs5yDW9w4P9laTFJgB5KJSMZsN4bH1BTZlQBZdJEjKMzXXQ7U2MFt09KLtsSlM3Th
lfe+LKY1XWfDgUv4i0EHDKj4ByHOZoY3Ed7Ow5Gb5aTdylb/MbJO97Lg98+hM3Czxn2CtqpRrliN
ndcE6Sd2lik+wqdEGoDGCQp9yD/Rx9oqjUoShY9Do8acOjT+Kz2JQiYKHiWdBhVPYgGBMlyQs2y3
vuKwsBc/tsy+DUhpOAct8K+QkW8gbQtMtFcOjHZQQAOCQEKSiWkdv1OqhQQgnLkwqtWZZ7kRgH5X
v53lyd4Y7qm59PeXa/npyq8lT1Eh0EEBWGGdotEsmdDKI1HDm9+gdzkYsSnh/1XYtMTzfqUMXXDS
f9BgduSaKEEP6h4gBusiFm9gDeb1wMFPn5qRb8bSe04j3NiqamIzNbrcA849SUBdyBcNgxazaPdh
IQkOyWecxwRpGunm1c2sWC7M6JX56uT+eSemh3+HXsdUMlX0LB92pv46eoyodFM3fcf+6/8cUnsw
klXU4FXj9XSLXJxDsILQuCDNQE7duAa4tPwAPBNmiNobWaUha0KiOdcSO4SmfXaoEfiZfYIlRNEw
t0XmcBJdvQiGEty/bey3NVMDcbY19aluvOwypspcHMPVhh1/NelpwkzE7qJgmt4DXfrh8PI1hvAH
9gdXaIN0J5Rxv3cvP/sLtfp0ZXeBmsVu9RciP5d3reA4eDk1lOB5LvdImo2qBg4F5A6Cm9Dez2gZ
k0LV1iwLAXz219HaDzDvHozRdGGIKND77m0uGJEANJrmi27FY90n55VzNTdYSy7MTs+ZLagBZgp1
5IN4n6cNbJCczRpi3se6rfGpZ0q7oYaVt0vmmzrTcih8PAHWNA7izwXIIt4jOdZ5Ept/fUjuhC/0
zmttgcrgpQQdLNoD/j02PcVJAr6AdnMMIdYIlRFskm2N39jA8ornAvwrtXMpfVque6m7YFsprvGX
Jzdxa6dY3L6JP0ExE1SjlRsIVsMXJ2o1MbQvVHkQ1Kc25G9Jwbma73M1ZlsxoYQEUjiHFfd7iru6
h4A+XjvPraFL/idahz7+kL+HUYS8CkwXfl1mmDs1WiKhYVC6C9/CTJWwMSNqwqpqbLWKE0eL6pAd
wXTOxYWt1CJMQBKUHfDz+KGD+sdi3bhdz+HXNmZECHgcmkSEpkBKd6wDLpA3rqBXD9bAxv/zCWpG
95TWIt+EGEDO4bLp0bVrg3TrDEkqz64gedHg2rQReZRsk6u6PzMTUO9AmozjPXLbMYD9cnvwrkE8
MRL268/r9TkdO/BTF1dhOXnuEcL/t1Vmp1eG7XfjUxazW0q3Fvz7stq7kz8m49gUr8wHqlhpwNtC
o3m7Lx1/dqz73ktsSBz4QiZGek6CbPPeDpxtfR3kB5UOpQG9ELLC3M4omT2+1xAGrvLvBdvjEvwB
dzpv4j6xn9K+wUZHbd4fO7/ChQMY9TWd4u4B7MWHtjNJ1SDD0lUoWgWPtAWiWLfXn9+29LyJBGkS
yRA+jzVJiiXPb8YbaHlAMGcqoQqCr1vgcco6sFMQwhziLoiwrYriGBgnkFaOFDNFOtA7wIs3a5JS
fARg0ZC+182zlUCJBgp2UsKpDirOs0AunMI/A+QyAD4JZba5fWxlPn7c1zQkhaz55occ/1Q+Tow6
voQZz2G9PmxnneyK/CdAVPUh12l02y4N5P2Lb4ZRUy3NaQmruijHP5FMTh53eImPBLwm1cCPZQRM
xPtpTyP2kDajsIZ+n/peXPsjnSCCV+v1yWDUXn2ZuYKuXlexzH8ZwAs4JreZlsUXqw/J09gpscrF
kpl53YTyPKHyf5YtrZLNFiVY2CC2YlFgE9gO7XFKsFBFdNPMiOql7yksjtPT5nfigc14780bhRa7
XVPE7jV6VsiCeznWd6jqo8WDzSKsLfEIfW8FuTLUJyw56BQnGPpri5GOLSLWWc4FDeTHLW2ZeVNb
bjGLsjI0qxM9SIzXOmCojRS8eBISpZypxBxEgI9o+aqjgaxyxITozBq39jrcHdQc34tNPKui0kNA
X8Y+tlB89cQGM4u2T6SOoaadon3llTsMZRPIdg9EvuF8nHOVPrG+2LDxLxHJiX8YVBOi22ufZebp
0ZHcYdN4ynog801uw3NVOKEqL6PJ9IerrWZDFNleUJ8pVVfvudnQ6sQhlhl3KrQMdXrM4YWQzKHt
I24uHJBuYIWj9pbxS/vg80WOcFdQSrSzyfVXZG2jDmrSToB5+DkhGn93/kuAPp8z86YyCeqpvaUz
0WCTsmZMzT44ysDBduzNQ/hfEqRaAUczpfv4y2vRG2TS+R42l/aPU5h1gy45321JMiJNB85K+xL7
N+Rq3RVoh3QcuxYsMJGp8XFMOQPtNDV3I7KxjAV0oJOAa8BjPD0ozfG9x3LvnKSuX9Qm9/zObnEr
oS2gaVvavbiwwmItM8isDLYSwtXjYpI6Ay4cej0K5buO8d+lDUnZelSZrDFLwIETzjPsxdi1yx45
S8yVgwqSjPE0KZaAckDJxp3saub6DQlKvsByIRB0i91gMyeInfgFpmhbQQ0uZJk0uANfwjd7keYX
9G48kA5TDK/H9teQT8jz6+QawwlWTO9oVJonEwoCjhSZYfrZD99iDu6+J2zcd7SciVhlhxeLObEs
GWMV3BaXY2tJyFjNHNebP8uAQG4Q2HM1+G7xa1Qe9laQ0E2CM3yxXfaLLzbAhY79P+Sy9RB+4zNO
qEgJmGMdMZt5UheyOa29l2m2wviHGnqtSddoz18wnTQe4BQTC+J9NLCM9v/vS7LiHdl7lbsIjeUk
c1NzEs3eJkw1JuSwxDQ2UuB6zJ2xO6E14STP45yvdA63HrCiXf7ZpXTwx8oEWhqyPhzjBp7CSCBD
o5L0CX+CaRXW8wLF1amSns7c2IMPD9nA83qaijIlzBb01713C3DDG3uyH8RcRf2tWV1C/ICMRbC6
3cnOt+UWmk4bC2xPwI5PSCCKDkadl0l5Q2QokmF5XqurMYWPDPbka8NGRQwAE6QbNxOYehfbXzD2
fVZ9z/JiVy+UfwDDyiA5bw5YSARMdTMI2u0GidnvarWRZrICtvEGqOjvlCeKo7bqQv/jP8zz1Cv5
Gq07xAim5NsMG+g+uPeId1yoJblJsqM3WRy4Ww7tvzS+pANGgtyUFEscDhUHDgPL9STSff4MIqLi
EFqUI6HAubZ7uWXtP53hSyZS7YXWRoopujC2zZU4RzoMU5rLYy0ZLzLJKcQB2THBEPGH8bIWcJHA
15Q4nzTzFhziOrgfh4RYwaKl077fAUosO5L8EQ/g9YPdh14DkGU5WSzrkRHGHDCGRqqu5RYVBm/P
gJD/OaYgLWRYSc+11pU7lniNrdYVERnDZujayMhJHSXvHJE2MUqc+uyBdBqhR0P5LGc2AQwRtBs3
qthMwfFopqL2RpREJr9xqoKrTSkD15vBT6Hw7ZFQ/Gy8m7fB+4E155vsaer7b0n2CgUhyNMHr3BR
2LVk24cLCLAo1pNJoX9hId3jmXxA8V9CM3qasF8AlMhZB++YtKt0whGja8Is4BgJjo/uvNyi1JWL
sOCLeqGaYl0+o0AutcM3qtJEF48FL/gwBTJHOgc6aus7WpARZJKy6b9U8vel86kAaxYSr9Wh05vS
qsURBQ4kfvrj3E6mQz42gBe4D7ZuYfLL5kJ15BGGPfR+oyTSJKISKRgnyVpvD3hULQ1OwKGoSOdR
Qx8AqnA7L89DTG4Tu6GlT/eXxOXBIxJSw50c4HoEfsZsW9j92rGIjU4oa4MSp2XZYCyc0P7hWpuO
uevTY9YQjo5UZ6flLHZN2OyQP6YJUkngOt7aLwEd6S58rvs75VPaymZWfpEaMVGJ9LVmsIhLOQYm
+olaLvOTvdJ7pYHv0OASGkgShjNWtekeChZcO8lQzwXJup4KvngBI7t/2NVrouNuDoPPHwwCZF64
4RbOnjULRs2zHJQpaMrf+jTqgY6yiY/3mbWihtQRmcU3Geyee3zcEn1cr552Co+LboJQ+dI4gf++
1YP/xM+u3NUaj+sCCI/K0ECxA/OxcaivJkv3HXrEGPfQPxzkyDGIFtJ6aNV9ORYT0GKByTO3Zidf
0tHXN8pgsRh0JCKizP6VH+o4OHDblPhsJPSOj8Zy8R/jAclTZfL1Pmfo3oSMfdtEzRBjNcsMYQJE
KEcGQsDC9L4V21/PGtywnStoMopAibtYP340OWzoIGH7Pe2DvzVVevBdhiaWjRMImjm+Tjhwx/yH
bY1fsNJ9xl5VOOt3Pf7hW7sxwQ9ygOPPhhRpryjGo2ac/21mPdajW3t6lllaSX8pv9NT8Gp+hT0t
BKBmm5p0PG/fv2MR9xYtTwmqBkrtXLN9gZrE74IJU8/M45ftK+FgN7UgtLY+HLxEeGcKXrA0EAj5
IDvEDODbJmc/2koOio0qrTeaptNhPRdgZkOQVPy9zTOjiMo2saKtxGJSRXs1gRR/bgXnn5y1J9kK
g9YzN1fceEYHCrNplHzXDV0/NQpMdG7xzvS5dgGQA1ca2zFIY1W15ei+DO/ES8jWFzhi4eWLP8FN
tWecL9kt2GLTlpD6gXVV7ciNw4UmLcXVp1rYwtfdYVXiRArLNFtccuQOREom1+cNvy91vBHspvyG
1KnsM5hO0edRAUa+q8ICfWCZtQUla7VVU6dTLS1c3mdMjx4FHis6w01BCLD0LI7xvhXP/tgAVMHd
rnLgBfdp2oraKCV1gV6RPJMZ5sSqY3EQ/OHbhyVfITxoz/m0/tCNsRILERoUnOwasgOuhLJjCeFe
zBXYF2c0z4SVQa0xU41VfoY+TpOtnrFKYwzKyotO9m8eD3E6l/S93TpFUJgfLpXGu/5NOgPDJccd
BhEOFzplGKmw9u/zdDXhuAyewBPTJTXAd57IbEXx31GUMMAUmGHe0l4NHS/dSVHcOUmou2dISN1w
c8CKEnEl5UQtgPoEdRE/BcXXCfYABsYK2VqZUajiXgXvlE4MReayUenzBm4+Rm2Y6XnEzSdE+g4T
oasbLHdQ54d0B2Mp+Tn5NzqzjTe+H9JxrQL0oQy5WWDp9eoKZQtwu/HTEW2eGEGlLCh+ebzTGHug
jGdQGZKe07ycnnQF9nQ/HeuQ8JNKi5tPQ42glmLLB3RiUwDSVrMI17bQe6v0xpTZOFi6rodezAQE
6H5DfrL41t5iPl6vxFsBn5D4kvqeFfh0rFRTWQ52djq0guC//t91AIDIRBlk/P2lPT4/XnuPEypE
tP/tLXLfVUZm9bOSQKzQg7IaeSkuXwV0XvibyTmZGAsnrnFEB5W1L8ZCrWTE1DfSMzhZCw5fgx3c
kquBrA7Quf/ne4wa7lnaCoNcRXbwKm82849AL1+yT6m1byOLixA24Fq6wt+pwMIkgMTpWwdRoyUe
veDXUEkRROZBN6yRLYYbuOEv+JxWuOOu4HzWPnrJ8EJPMolCqQXWIkSrpSgIne76Fz9A9WIO0osd
15VR0I3us863o+16+cVRKgj6JhT8sDptLW4ZTFTtFXQxnR+hDjZMg4ri/tJkjgBStRhcCLKfMOAr
NRUD0LjW3SI7dGLbTMeluXSxQPFJWkzwhxiX+g3qAU1nlJzAOwL12PrDxJ1wwQbsW2FkLGFcpxCY
zJ58oAk9MGhWHURRKMoplaVU6n/Olv1udzw8lCiRn8ngbe9DkGQlxE4AJfZlMKh6ePt3EN2vK5nK
PajlcCE+jr1fPZ6WZWTLWaR6NnxthKXNuVH4JLTJMu2OfQxKkRifKM1krwpU9mJWDb9oYJkVUOrX
ziIMS7cQQ3qdDdpi5IC+ruTi1sg5hHK+VsoKlhQy+AhU6xh1SNyaO3CQG2+Sfhis6yYqvUsnjXuO
S0Su2O6luvjpjO5WQg7mLUeT53LqvtagNb9HrmlU80nik+39E6nXkZD8WRa1dNFJ8o33Fy8Psd8g
pdOQFEyoFcjtK6AjDE2sKFeBDfFRfJlCvAqDn6qiYXNYw7h36fiwi2Lom8Tz+RbJ4raYQ/RchrSG
eZ0wpxQXIwwhu4itLp+pZwIuYZmhGSoljZ4CK3U1Sja5o5446BcNq5uc3NyGiYs5QmzLdYX7aeKQ
FulLkBAS7PGhm7E7o998QfFThxlrsN1r7g6BIoiUh/z2B/6ZVgTOt8AEDqmAnZwAO9dpve4p8LHM
x4krdiMtkQ89bU8RTMrzyvpjov6Y1wtdN73Z3+FI8R8+vd8yVGNsFEY/H5KTxXqBqjUmfrI22KDJ
Xs96u9CdHa5ej9u89TUhpqPGy4B358OJDwO9JJRpuUkIuSS5vE9rS62przp6AzKYBfLGpjQF6VEi
jko92w/MAxZbgHDz2aUU/JmczvMgTtRjzvPpYzpTbNLN5rJNK+eHYGgfp71VOPARkK+E12aZMqAm
dNqgrt4mzk70LddAzhyiNZHlC399GhawgEG4/7ICgD/AMlE921s9LX4/STiObiNneFhSRRa4PHy4
PFUQ4EQ2D21cYO8xsCyPsomts4VuELGSdfOEKfvGloj6V6CRtSOGpfEqrJTlztZw6IDAQt38oxOQ
0bi9gx4sAKObJxR1XZxWnqpbmAaw/K8BsGjw3IxfXAiQcPMvVszdSVDXVgqVdVyjkC4BBKPniV6q
wFz2uq0yaU1DWvCd/2s2TGNqBgsbxJ1IbtQSJj9en7n5KtDDwNFR5wsrboonRtBI6/lsVa35tQ6f
n8sEsUTuvqgGvkkn8QoVSefenBETQiGBUd07hIrYYtsvtuLBbl2SdUC78jBJHniRps6uS8q+wq46
v8U6zEU9m33m44Cik7EYOmHzTVpoSV8UN9hrDMb8qxIo01kKAmyySkD1Ci1ddiWg7zu1UK0f+1ZP
3ogHZknkhxQO+y3TrztP/QngLs0LtW3uqvftgojBMWnAPnS1ALLf5sCBoTjMpjuUpN/FRPjSxNDk
yGd6VoPfHyQIdq46B5qukyI+joVze+uSANf1TKeB32ZdC7umaitVTbKre5OBPctghcXKD02NfzIr
BOZqN1iRAbjeAJRCsM1FKLm4M5U5MkVA2fMgRnSa2bwvf82kogtQFPYMmi4g1TWilyceFCitDtic
a2cApWlK+UvwGBlSA5ZW85JzpabDMbkBo0UKY1d3J4o2rBq6WN6OCHXFmZLGizGWblI5fZCu3Nyv
4RtdjV7inN2vSAl4RzTF1DggjMt0sL5/bzID6jaMbseT1DmpgEI4GVAnICpkMb7WnE9fIl4VCUhJ
hrL2eht37xvAXOpfHV/dNeosf+ygDfEWdAFJniay7hsmwOVLKZ/JbSfuCQYd4w+N2b0a24rQtEvd
WPnbCm2G83DTONl7yvnkK+il/cBmFBLbxAQe/QZ1FD1upXIllMkLsoXoWQjeleQo8jDuiFd36kqT
oxTgl9ILngIKe9bMBWryaeS/J08SIKs6GmEAeqjZ3Embo71NGUbYXPbBKLBoIwSP3ZbCp4Bpw57b
N07b0QP/DE/3WdRwUph9AMtl4APBlsMwPGTY3KOH02wxH7Dn7IvgH1jXhU4ddpu27tSSqGeUD7qd
TgMwgmVO3O53MVMlH6M265JRpRg8lfQKStrxSkrUFd22ITkrHz2411rDbACxWxAsIv0Rr6buaK/3
qoKqSj+pi6DWlF6KYsbeBR2IyyQAE/KQo88EbFuRWXZiKtxGICMQoLw4omVtskDCpfCtn7w4IIqF
ENltmwL4Lh0OfdfBBOE2FNsv3QhL3cGLFkEI83RptV2vGv0FjIXpdjr+iu0/Ms2awX0xoR0tsnha
b25d3S7Muj/oKZPG3g3VUnPOgF8aoipzV5aEs7dw5u8nMouBTOzCGu8fJyFNomGK45WTFI32S4Kp
4pvn+KWF7J9H4xYuv+BgsCrmOvtgQFR9ARB/wqlo0HM/v9WvlKbt381cOxADkeMUp3vg7RjdYFjM
n51QpiurYE12O216jQ9LH7eTqElzDeeHQkKAcE+8HChAKCquPm8Mhpo6Q8m4pMRSYDJiLiilYCuz
guAFykkZWlBtMQYZFqSzFTpgiM+uKWBRK3gsAaLPornHeuh8qHmiyUb96C3ennm4Ppdm1e8UufgK
FZb0SG+bCbWAEKaz+9JqEvMnzYOo52nMiyQ5cE5HjEUvx3xyRMKQDsICX6JqbfcKuBbdaVQfteAP
A/GymUAwvdPPBzybbbZQcGoWH7mKaA4xMgbmDFgEU2zr3QgMcQBdVNjIbhrt+SKwqc5LtEBEegd6
T8OXxTWEMpbPmcHarmx0C0SKjWjIYkdlUsqIUP6y2a+C1PoXT/uhs1MxryvM52JArG1H2Rpe1WDF
0Gn8NfuonBXjet6SlMwqS5L7rDAFnRolHqiefeU2RNR3pRe1LiKc2Nao5Z8WxoOVD7IxbArE+rlc
Vz5lApGxbqOFu2Qx8P5F41KSXd1izB57PLS/pwPyYI5FABn8JT+uizbpN4h1S0SafdaMcRur7YuC
56sVwQDl2iCFaAmV3YL50azGPIVAr3KsdkZnf2+5R9rUuzdGe3GLj5YNStxUkgi9DPZHLYwoO9Q1
gNEWb94sxBwdV7Qi6vk/ZdbrTkkV6vN6wj+q4SsPMH9hr7VyHpAWKYoA12CGbP5oFNLPI4i2IsT2
NH3+bwlNkkHzZyIL+HJU6ResnbHax5DFPlD2h0DVzs7C5XD5omXfpQ0XvpfhggSvKPqAwKT/zPlC
SyGQw1Uwnpfn5obsAolzLakRjATmDghJZxDHG/naODuOlz9Nbr4aEyRehJfJ+YvFYukgF0NJozWL
z3aOEuhdtNFDiIjkpt8tYdy/uComTZj9G1WW+xCgytDkzZNXS1k1HYDhw836pAyVk6jW+j5Vf/cY
KuuCV/zCx9a9w5kW23AcY5qa83PQCNqfWIT5ch45AP2ecpjVYZxpUtwb1/MRmJKuj/6SJ4tccgNT
esuM83oRrGcbPNLSRQopO84iKPmVmfEFDV/wLgAXqw3aeyPDG//KkIvU5tnK9xJRxvXh6cpdVLvV
tt1DXkl2eRvDHj0zrFY4e1xDjDCdXR+3DN/4p6cuIJc9HQsQndWBWxL6NvdgE/+0t8lWsPpft38b
zpxlxLdR/DleZJvhASTY+TgS5pS7BG89N7sXF4E2K5ZiGU1NwnVV8H3h98GqKBAFOejjfqEbsyVi
gDrt8jP9o90P/MWZBjrbVbDyc/T6fReR9at8oUNIoRIqbdh9Yj8Yvwf6oHlCWUZZCtnY3z8EDajP
2MQ/sCrfBY6bftSr7iFJIstygLVTJDdtCRVVVh0WoODq+q9RUhp0W/RNvH3FcbNKU28qOmuXSnO7
6+ghqwgAUdYhOH7Fqa9kH6pM07G8Fc64YjxRAtEYQm7Dgm4VBd9r9NMCDt4OPX2EhQ+k/tn5ECcy
buJucxPG4wIkSzOqx4bEs5yV1wudf1rRH4S3K2esekeg7LtZxL3zmOy7rlrNkkkUmsvb43fiP0UT
CNbpGROYOOXOJTPeyke0IXzLmEU3fYhZL16yWK2Cg9Ha4n+ANn27wM/7Ay3Nuhoo7YVMOSeIskHw
d4wIDeLccWVxbdz2JgZUT0fvmoQyfQOsewFXxru7JLedI5Rx+rdOFJXSGer+msPfvpubOP4Vlx3Q
OHxJwsgzts9ZlC+xVsvfLSsr0K7iaz1STalbXrRGK7rJsC09niDmO2LKK9AQtvieds+0uTpqzaz7
dZusJy/fNNpdFYITEtXv5uzZWpR+Yuv/vipoMQ5/84ngvAH1tYRku4acsZDTLGIB5yFGS2ZjlEsA
xgGMaqASV77eqjCRkTLJqMBZ1z6ieJsPi6k/V8y6Y5WsJCGo5lzIPtENCbmJEXc2DYaGY2fBh1Le
tOtKspTM6N3Lw4MxX40fjjVLkAFeonSnB3wqicpwoRHoWRnRA+tebREw6VgXIN0z8UpPF38Y/TJl
GMjdOcwO9sKMiXOYvZ2OpTF83pH/apfOqlsYjc+rNgyr62sfUI7rdMxjyhUOZI0qj2XtJiTCYuL8
amVEleUXqin0Mpy3YcPhLIYSy1OwQ9eY15G/O0moPedmDa2Q2s2TQK0ps37irCIggv323Af26qus
h+k8k65mtZ5rQwp5NddklhXDls93osK9uzdEACIIcaTsyMhlPXK6lWEY2ANjM3h4UemB5yEJtTNm
lfy0q9BZI7FEQZMg1st3M3raqoFvKgyQvIHl9Sr9p1PnLWLMQDzrtJ1vjrlTF32AS+U5RH6PN20M
34KO+ayKn/T8pLfwZfne1HXm0Z5dxifUi25rlxPkB8yK+bBOLoDq1yeCp5OatR6qL4Vq4pWYJcVw
Rtq7Ye17AJ07QEb8sOdh2MuxnQzNx7GdbFjN/pWrjryOC/SdIOpVC91lKWs+T0FvyxlaQJYgu/Cb
MJ35mVGmewmy3mMcYHOmHSC856SvUqrZs6UA93fv/j2dRa/bFMFkFpxPDVOKY/lQOGzcHLV4rz+o
zLz+Z1btTRHyJJcLfUodrYv3vVWsbv6uA2gB43PKqTCWHIfTFvXarZ54lAv+GPYrWUqPHoaICphW
1V03YIYDBOtkhswkUGTbYtz5438POkbzfwWJsDVcL2feincO8oRACPVO6oNzKRm2dUeLaF/kSd9s
AjmyqqwbhpEcfVyE49lsSGUYyl/pzm6hdEyhS+t1UoT+QtEkTXyCbROnJjP8xYb+MzaRzUqFAhlj
DfJrMbPgJG7Rk137aW9yrBxDY7mGK5wA6qM3iySll1BhLxc+kK6iBtlZGowMk1mvwmdmuuQ0rNKQ
O5WKisSTF5fpZA86xiiJ3viIkU88VbuJEgxWnZG4NhV6I6LJvJpd5X723RLyklg4pYnnxjOI0RDI
jZmMe/0gQOqfMcky9khy50XulQhTBtbdMKGPoSNahSpLjAUMNQLB3q3DfRNTeWsgtP1O0BSgHFEf
i7Ek7V4/UqbsxUIoLysuvU7+uDdfmFsuLUEoimwImgXXCfRlx1FeiXZSL/b0aCLClybsNyZM/oei
6P/CYDy/R+p/AF5kPUKw/HLzCxCF+fhGTNHkA2INvn+sf6lteilhVC0OS+JkCwwZ8gK7Z2vHmxbZ
OoyapR2NxrqIZmNl2xPrQwrZTf3RBIPWov3jKeV9d0oLsrZnZZU25Rto3PG3h6zWO2Jbb+6BpAE3
Am7C5zEk7RDzS20EPvnsYBHMcaUm0SMdjtG/Lv8MCRmfHxqQiZRUZ//JQuaUx/YM9kqpaD4aDH5/
HItMDSkv1+68vvWLoMWRtnP1tOHT9eDVLub/73491tkOfO1Y57R4fIOj7OT8I2+MPZMxyyFodDs2
KlZD21a1pEq5ifp+4u2Hx49ejCKE0ieA8SEgvsBWhaOkiYaod3Ioylw5i0KS89tA90RTg7Yc4i9X
rNJACg+M/DE4NXSxW7/4hAZmCxHvMgE26zbFa7fX5VwsxsR6ZDkZWvaeDTzjjOH5o83Lvfplhe8A
AsMx2hha+x9QhZZlYbnPZfKvx1zg4PqnS1HZm3qJ0dbCFfFsyoq2v+SWC2CKcyYa7g8GEDR+JU8V
alWghI1gVJXz7DS87QCJLKzUvSzoJsK9BMjlg6htnzcHIoG4X5ociHTDgj1YxZBzAHoaeFUBSXxB
I9isnA+iW4pyjv167fd+wMK42Japl6dTYq/zfVXoLqer5Zeqkt2T6SmcvWldzUBS1XSwQwJfAQqr
CHUq+j+hg0aqQS4eGahjWybG88dH7aiLXji4Kp9h3/b1EBFacm/98cah+E9DZEfIsoGIBhyQ1rjx
X0h2TRk2pv9ZMvNGIlPx8lXX572bNSDVpiCAGIaEvz1sZfU/w89R+SVMx1bm+jAS0vSllqLpmltM
6Rn2uMrrpHbY3quIU4YdJZfX789l9m+29CCdmT2nTXXN+jqApZu1+GOMoLTyRnKGVKqCS+fGTCd1
9sDpJxFr3ty39EplNV3WimIT6tfoZkqQsF359BXS44mrYfQpnMMj+S6hdoc3qIt77pVqR77I1lS8
i2ndx3umc8qvz4PciOosYjykAQpHL7Pi6q8s42DioGfWT+exsJ3Cj21g3vSglrKER/zbeOTEeCAm
Ln/BedskLSWGeO+mu/v3d5fgDTwi6tJEbIF4KF7hmfS+UP4jQxq5bLT59gDdL7id9BhU0Q84018A
t48RXA/nw2vSVgQrJSXTzI2/k6yocXPcYW1MYhXVyB7kAyM7q2RZW8p37O8mDM0JOUnrCmuYU17P
V8nqmJnUP4wL/mMB/zNW3TW2UdycB1CEz1LH7sHm8ekFhiFW3smsg9TbrIZ16Oao6sGjC9qKksxl
bkyQfl5POhQA35pET2wgxfbxueTUH59meQEdKm0mNqP+mbngdu/9FUcMk0cq/pEg+U9n2k+O5vD/
BpliyR6y2KZAxJokNdTIPbw9PzjS0kO/DD8LOq5nCIXNGk0KTAxegTPDxd0fy6pcMZRnBTl+rnEB
irzry1D3CUHc1Sf9myYL/Za82UE8tZIATc2hx0CqLZu5UwugYaueYX3UhYtWMgCjXWBTJC4QvlM9
n2xT/I+a5PCFhESpbjOP2p1wMHM5jqTv3pCNZSiBu23+9oNT+8VBiu8BKcLqbqH23tSXH11GTxTN
msxM2lt4jD52lrmVCwAYqtlmFcZLj63f2bJGVifLywdDa8mTihB2rVuY+jV/4sxNTPc89GLIGwW3
QWYWiC68PxKO7K+7pPq+Q7qlIIj0jYMWduEIhZEhQgwEDy8pLfW5UqwhQcX4soZJ+c922JODAWZ8
OLFUJnVRldMmfMMSa6Jc/jjNFXFEpOUI6pNnj5Zr4aYHUrz5frn4NkuSN3UHgHkQbs3u1oM1p1Zj
iMqUvONioaLYmYr+bCyfU4OfKCTkwNlyCpL3m4iAKEID6ce7Y/cQuCn+Wd6q8sGiv869uZKkJ974
1le/5s2KN4xMoke40KZss2HxAfvfefJ+4d1wCEqMz4OZIscfewjyEi4O7iPywX35nE1VldBUuc/F
IFClGhVg/Hk/l8dpN5n9wXhrjl5cteonzTIhQBZ3XRLiE/EMk+QQVhAmDxXzowwZo96PpqOicWJB
hStzdDxJyHjVg+/JwK5M+aKU/MhcALmgqSPKeyZy1gYLnGBxAohiOLXs18vgWv7sndSVvC8PJRno
iP6lu2HWp/b+mBURR5Hly1E+b3itcfZcrvecyxMF0t0uNN+DuvpmwwmBBFP/iBa6RM5cZTOfhxsZ
fH01kwxaKcuXeerE2CzNnTjsjy4duXUXpwmcz2ept+Ei4eaiZ0iGvQ7z6/TPvV3H9/836t/CxNT+
INLCm1JspX6hbzB2i1ba9nLvtvAJ/B6z6KNQ+J27OgqBFkG/gejbc3W/3FU4c/XzKHUN6HrThUFD
LOtYWoem5oUQhqL62nE2TkmVdgZcBIdhcfEiEaiF+duW7tnD6kKrLBE2w8eNloW8MmsEhYh7s6Qx
P7aGklq2kPY2RRuClF2xkHaMLeT4mK/BX+g5SsTF2YkksTx7BQLlsIkYjju/gZgyfqyOhcRam+nB
4dHVxCDQSpnhkRkwDkSfzNyx7kf3dKkH+9P0Rufj/KYliO4aeSO6jG+9vV76WWPRDiK3/tGrXLf5
3YPi0lhs2KI9DqQf5+cV9K/AYWlkBOGLMVOMj10XnJNWoOBqJgW7FxOctq0JBGt2jaSGCNW1vk8K
uKtN3KmwdHBhElVHb7Dj448nqB3edpIeO2oHoi1lOwbUrtw1umLIiK7OwqIYt9iZK1E9MLRCgmBk
wQpBi2s5tAg3IiPYPKWHB2qOtb5iDai2PgbtMjlqGh6MiquQ0ruCb8ByGXYYn+5EhfUXGqwKSn8J
+hLOzxFVabWZjmVQ7EntYzTdDi4cCBnwpFPWDbZ5GgWR+9mTQutcbb15LAmHk9+z0aCPW8IYqobd
Pb5XEJkbRTdjXrft8jlTHp5bZXyVMm2Cl7PGQHEN93dUtC+LjZ5dgnekbO5qQOChZ+C9xKGWQ8H4
KVlvRQ6XmilF4Ij5LkW7EMFQAuuAcuPiwUsWsGXRkH1Vq5+DuHWF0hYlDIqy5JtTXoCoSd/8sPI/
lmRp35xdUsuJ5hyKfPt6b6yg7uGYDa9x88tm7ZoHKrbFrGl1x88DxmK2f/jBTzgVVye9OfDlSpAd
BlItti6ESeWW7XaHC+7QbnA8AXEG8Xv1ljCRNB8QA1vRHIv5BUhdV+efY3GP0j0YYoSrHm2er8+R
ppeBUQNAtgRBvHG0ulR9g1S8GCW8zReUgxuMEWxp5SXT7MuOkY6Ni17lRZAfLTgQsElcR1gSo3dG
OHGC9GCKtVdEMQgTbW4xj3PIvyelRaxBHogiwkq/muRp+j5lz0yhCu281/0ARG4kBN00hvBypnOt
s2KlpXBkZZi9+p17WHMst2YnFyBNive317qwpWmTLF43iPO6IhE9Gm0EF63YU1SwBtdSSDkoemmR
O3PPs4HKJ++foTDKWAYlqxRCadjmsvdyBE52HokOGyOzdoxZJqU1Y9Y5Cb/gNxh6qQvxOwUOXv+S
4CxSrthchKLOf7j7MZsAkoigAS6epsY+TBqqEkE35tZIx/Z88OUyPWxfswSt29bKxTuAnJB0oC6g
ptnmef/0XHlqoAdnBjxcJtLWe3AI7cE6BGlvlkAc7kNyHoOBEIpoa1zu7Xb4gdhEIRxsecK9QMAC
9cxdndu5hZV/H0+QrJjvhFtb9yStaz6k18d236LPLahAd83z5aNUyXq6hRZTQI5Nr0PvnxrA1SoY
pZXedrrcEG75EpQ3xwaaq3Kb2XYpZcJ32r8jYEfBNVJGCccoGw06OQxLE709NV8getTuPgd/w1Rx
CackocrI8HnPsKq8jRi4g3hxNS5JloppJK6e4uCN+DsP4+OLGAPURLNSVQ0D31ODmJCwqkXvWRk/
9x1fTcTsr1gwTm89kGRMtFlJdpJgthAgZghRZSgAofy95Whdi084VfKpmwNMHcktjlmy4InI6Yjm
agRdXqhoolMFLcUyQkQPQRzIYW2/+DrosNj7rts9tRs8sgdwwLvPQRRO6wy7yV9BuSa0aLUxRy1H
cwjKLPYIZPaTdc/npNgGSd9oFQd/C//BAU3bw5PUPciN7M7ObkRSW5qBiHkwrBL2BH0QNJ107Dr8
06R2kLdyNTFKAeLkiqgB0CJAmhVp3qMJkJ/QmlX9n3qDuxQcm9CDZOzyFGoAHhRClZcKWGOaehI9
yp5XrOi08Zc6pRR+Xthp16cqg26QWLdbrhBgdyuyw2OzSXLEi5X5mkCuVGuIgoIw4Oew1h0n1DpC
QA0zjkwKyXVxV7nDpvZ1to6mFChwVShtK4/CH20JVXialwXYsPHBGMwG/1ubblYduZzA6i0J4jcY
XwYxtmeEBWKuQL2G2vtr9OB+viXfGqzHEOAPlJpgHMmAuB3y1v5esWVQNAdCx4cH+vuDpuSMzNfs
5UPWmc0X+JeUingUQ64/g82YEFWCmak6dTMsfNTX0eF4C9tut9dxbIbWUc6yzfn74+6I9hI0KYOB
c2WGo76KKGz+aTetqFKPXEmh8rWZt9NXnBni2bolWXjZNvYHjb/B9sDC/jPseL/KVgaKDHGrmD6B
aWedyjrHbxMcjM+fW/SdwYqjOfGfUumDDrERDXnScH1RwFJnkZr1Xke8CqAlmYwr00PBZtibGdwy
4aMt9n9LNgfDcgdjKmGXmLlHDFaImb8jo2yay91gW1ahfvXql6W+YhGOUPE0q/HhJ4hsdxCWBXA6
2UzmVnH4iHb81fZk86K8A4sN7pl46vxyysKRoHS1/8tQ5g+Qk9KRkNeSkaAsI8X3V+GPxYMihZ/h
GdagPUbt2RWqU2VyfJUdSgGoOP13XUy88GaV+9KctvjlK2uKYhrwwTd8yQ93noifX2DMGQ4T/Y10
t0s8HYCBFygkJAMODQxlEVh/LcT84CwZ52loQm1heaR0c6bG7wRa+hdIbOhOyglG5iKoHCiUC1VA
/ysToU7GkaqGJOCa2lgrM1IVVe4iSQq1SQal3oXGz4W571UWvKL8o15S8x4o64yMtrBsXh5VLxHZ
Af6uMjehUVkwdx5oqmn2LMuziMNBIj/BKy0oAFNRYTKbA0z/vrvZOmxQihLo38AnWl59YaxEGyg1
NekC+htMx5l1WDQoRS3PLLoTdFwybIcA7iEXKyuLnhS6j7G9slktM36rvFf8kmissSJOL0Lwd1dz
BNLio7JP6g3bUczw8NrzmYIu9L3bM0/cbnKJbttQRg90X3y8tnFdUtwsgRV51IweFMf/Cw/DW4Tv
XTgvHVE2iG2ziPKoniue0bMAbsCDZuN1A+mFZLnwBgq2sQ90jlJmcB4taqijDHMK5IvbTzIPMhKw
ECeSJgPaIlkVR/ghmApE67nB2ykgizLLCjXGBRtGSqWKBXAIFUQUl4KAlhk9QZb07dzTqQsYJ4Tv
NBkluzdVE5MsPHukO1gYrbPe6IcG6UFIK8tEknER1hjMJgEW8yF8A0wMPE0hR3ZxeqXJLPe8djv0
eSWTHX8FTfOsN3nvoA5Q1C+2+Z3uJL5LDexN8xNtbLP+UEB0PHWtvO9I2DD02ejGzAFlcE+xP51I
nQJsngPo9CXWtbAkjRyu55oqR1y0BMDb+q66oL81KjCx9sFU7meQWIgdew44sM3OKCc2fpRotT9x
iqX0zrOawX5Bvf0MSoDaflKNIoBipS7wTjAa7prL6KBC7JoqErS6kWb/OtFeSLUwnEq/sQqwgETD
K05XGmW//z6LrWPsR1HDhLcW81ow/Qjn7qoF7wCqcoE1Q+HUmEN6hKZJ/g5CS2OuNTYK5DeFxgvN
HPqiV8yNU/SZP2WfpS5elOG3GdcdAizt0gICgYOIWPdWSB2a/gM2EuTh5sgyAPfbu2xDNnlLgePk
W9OcjDk5hw3OHggB7TK5LrmIQeu2RnnB1CzwkY35SoOEBr5BK0Nwp9VzIIWKiIodFtPNbsu0K2P2
WKNCfcIIDl1wvZTnFpJ4VTTcNk5GVHH7CrTzYSjnj1xviKZGAt8TjVAixZFz/ptT5r6T0MWP51on
SRyeMGw5eXxih1iKUYFJd71gJ8IFKTlHVQi/Im4PSjGk43AnmeLlF2t8K95aJ2lk+mYe+J/ApjAJ
8sTYFawMKsXITgAVp57nqDB0IG/Z/FHK6lh9muaZDGVl9SQgYYXPi2V3SpioCunaBQrJyM1ld1tb
5IDfbg8mCmbeC7gsud4bD2ORWTNfFtwvFTZ736vZRgO/4ACGOpRbaiOMBRZle0aboSf6lHU+/S5u
RcK/lu/7iMgEzMZGPek4oWfuz10bzjiMXE3FaEglanQuajGwe0ToLIMrqrZ3EDD04J1QKHfT9NNG
wOcOw8x23UXwk/MX7PtoEs6FNvJbowwIgCExAPHnnCeyYXv7XdQD3E6PTdzBrV7zKllnsTcGyGGH
4C99u1L1bQNaV/GBJ/zpGIIaogrx+e7ZM0aUGmJfqljZPcYouaCD9MtKTTFSNlyTVo3RxEI25Btq
BFcQ3Bj8jclqKF0EIjexWWSFrsLfhr8aEK6DFlDecTjWTn/M0a8SSt9ITxzcnTjoQx36CFphqDre
rO5wwVofDx1j8BXzLsCjTVrt4jYTLJxuzjSafGFR+aFEe63IA+rVdoGzIkKV9YB8lZ6rFOLyQX2W
HfJTg6w+Br7A4OIUUVViBfQzsHWe4KYE+NZ0gqPjQ3J2zun5BXx9LwBXft5Evi1iaQTbS8nrMSug
gTLJQlKZsSk4J01zvi0LuxOhbdaodo6VRRwC8W/ETE4lbNqhR3iS0b+OX7HGJ42U2Vm5+WY4hLiH
Z8p0gXV47FjSghlw7i2vAC2Dcsmta4z32WTJ56bi1DtfHE0NS/QtIc84UGJ3iRK7Bg7nNps/cJAm
S60t/IzIHZk8ssZbPz6vL/c5NeTcgSLczqwBwlTTbM/1jwv1LrcZRpIJ9K96CsBYNNH6lwfkklQ9
ZEU6QWfnZlcg3DKr/rdDDSJLOY6UurK6xxMAdzMf8ZepgPvqrlujZah3ueaXzXbTXfiH5+0dNyIy
zD8PU/XRlfXC+/ae/IBfi4J3uDonduQNU90Gybn9bhSS0/Ard2R/6d9OgVZSCoajoevNfhSGTZtR
fFWCSMBXRq2oBA4O5M/b1tYhyzO6mPv8nwRxo0ldfgDOBXnaJvJ4m/Nx3QUWQFkusPedqg3ZOnM8
NrFLSio1Wl5UyIBXRlRR/xT8N0yMHrXMh+bTOx5dbTQp/QtZEokIuS7vtHsQO0LaHtNXUEUHmHZ4
pJ6Uq4Yrsutv4BHzXsWkX+QoqPssiJOzXUvSMrMAkgEpR6H7N3VpeywudXpc5dDFKH+j58jjJWc+
iEjyHN6lmib4P3epDtDi5Uf7AGiTM2Ez22jMpZHPs5IsRf6t6OcnQ4Sr7OK/OSB8LwBi55495Wfb
jHWeAbkEpG10VrsBGdYLwjkc+6fe72492u1YntNMp2bfZQf17Mpa5rV4mGdbgtIrqOz5bu+5K3GP
7CoF1nhNLWSeUY3OpM1uuUJIfe6RfOLbxsFWfkmazqhKo7wcBD/ukYL/hFFiaYjZ+0mQFKaAlYyA
+FIVZu9vyHtubyqdBcLfN1vb8EX+QwptvicLKaZTQmUSjhOCGGnL6yKwkkyQTaxgNnjo+RK6HpZR
IpO2HFqSnC3Ox+KPt1Zek8Nsmc8v/jxZ0mglDCXJkPM7KBZ8Rv3LsVUMq89FcCox9Xb3cF7gcGxU
PqInJtGGwQ3lhMqKqO6ClPIlHUzboeNp3sn8jTT1PHF4Hxlvq8QfyJfjfmDJuoAdU+MR9dHrx/my
Bi5dXEQyK99n3i6YBiO/+gop0NRX932kO8D/C/ocP3ssg2DyNvchCCp9IJxoRnyjMfCuDKSDx6Mq
2cQaoJOxcLkB0VEgxgruW0GYGCnoeVY9pZk/1xiMgFImk0qXHUx7L/YW+7BBmfBCAgiM2mgsdLXO
GvzwYhrqmVqfD2ivkFpgwcX9UWVUJO75j9CO1pRplldjC5fSAYVcXvvMBoHD25RWv8HKERUNbXzM
YMIsVb9z4GdIsgVNtGEdc0ZWqq6kMVEowoMLSWzPRm2RzuVQ5K4D9YeIdxXrC2HnwJHvreux2HvL
UCgJa27NQvDsWrPEMmZ67CzLHj4UnqwEaNPVwE4i0NbUH+AMHaFJaYz3YLoaea66S5eWsga41dZK
mvPB3UMV6QUtkp7uAjPLQt+FDYXXc4WNG4qGi/eky7mW/wrutF3OMukdsRU+vIfATswkjds0/3Jf
1olkRVfNs6ISFPTTzgXETD6ypwglQD/fWKGyYSMTECitv3zuHoPlrPgfBA5j8rZoMbnx/y5kT80x
2CGQhS+em9/kdEII3VgYyhl+nKFR3pykHuYkByyLMgPi4dhtPER3Nxjy5ETV+hJHiOMGjxRoub2/
tdFXUFacbNifO0ri9B1011UAVjqMyl3ctFuzR1FH38EWLZi8JeVuToBaiERHVsyruAaQ6GzAWw6o
A4JcFcuxwAJqHkionRmAPE7M35FRINOE9w0ILKCiCRbG3KlKpCezGO7r0PyfdeOpm9hKmao6moce
WnOpf2I1ICYbFPWNcRPyYc/A0mPagCk4gxoquncQm9gSFqAzHEEQpzBSUHSw+31/k2bjb0gBShMI
58qbv68Ldznv9zm8uzEu0PGA/UjOw+zJVF3Ovwz7pG2IZcQi+mvtn3nJM4plZWvF5JeO8IX01Bio
t2Q7Qs7vvV3Do3z74+YYeUfDQBFmjd20ttE/NCYAf3REhelI/XhwSxE+ukNNlkh7EbGzusO+lqvQ
797qT4jWuy8Lva615jkHHGSTH++urTqHcLHE+Xsww7gnt6eucfRn5Gx/mjkOAwP/SJ7WTQgiNSWO
qeyfXiHPDyhaQi61bNO5GAx3aCRcTGo2ToW1ha4BUaVaQqdo1cD4pxMsXcs71rtqE3uwo2aV7SZc
N76w3p/OaSQvwdUppR0OYKsda8E89fEb09v7evXdpmPPaBOerfUO7dYB7i4JSDVstjRZGgLL3dJa
Zhx52U74JHmews/NNbtYHCSjSbXAZJrN/wMZiMkSBN6x28yuEmFqABWjmpDOiPA380AkiyqiNONe
c+q3sBOwalrnsyqygd1xa1UlTUPTCamAPmh4oot0OEyrGrBtuEVHk865Uq6D/IWrR64jQ+LQtg93
D4b9+eWqh0sZiFs9DOchgtWVToTT685x3dvYyeYOooX5hbTbMCZxzqnU3qlFb9085XUS1eaIk/QT
dRm40FIitMKhf4ACve3jRrl1wU725peDXk7NXr3quajK5jiK6rxPdvWfqCBIM2asLS9FMfBIKN3Z
5Bjqhz6ilbz4HwW1MckaJ1rLwWEeL7+pXCOBxsY73/peJdF26ykORbh7Fe2A0AeMGCSwkWJYLGgH
4wuQa5X+5nuux8BKzKa71+alvxbfHT3tognSh95289T8gjBPJySw5mJHgRqVOQPfOXKljvqWmS55
YS1O+Iv2KvNdc2fM1xHke5jaVgbCszJmL6IzondhbmXFr2XlUnpPUeUuY6xqcQrGyo5DIYEDBuJK
M8DpniwwPk4+XtSWYSUHC8hr/IgYEMFas6pdFW21jPk1sYyNfZEMUiqySM87J2Wzos5RcozDVAqM
nf7TuVm1RghqHgllp/z7JFkJcbCxt9PmNk+loj6y+RhfSZgSIRm4zbFXR5Er2PTciUA3KZFdPBEK
2EdkYp3/zc3hbhlfpDma2qUsnpFdmXQdwu+eIpYnON65fzdrcSPWdQhlzzRBn72LkzVn/N8WO1bO
pSvA1qZrciEmErjj1ZASemrBaGG+vSnhOE12sjNkqELHu07pHD2yOsullbNcywLLfPSvDtIVxut4
Rqoe5IjmH43tkzlHm9SApOyppojLO421eFWOq0vLPQIwfpN+2fZ95P856hmPjSzPsn/zN12AFwgx
OnMuHPK7EHbm0Y32cMzD9fOZz4QA6QXCR3OWSvIj61l4+tyW7wzegZ80knn7Z8QFUsqKaYWstQWC
iaM6H4E5m5cvbXCiaRSNlmm2ez3ywmwCeM+c5VxBNTux38FEX3eWSw0ZkDuiG7WZK+wyB+4zyqFY
zEYM1BOZsuJ9cauLRVdcwDhY2pJmIgDaaj4/TB6VZanu1phZEnXd8Y+1jPW8DjrKGfc3RPObnse9
Ct43iyg/d814kq8iAYOPf/HcpME75xwt10fkNk0mK03Otr4=
`protect end_protected
