`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
JqM6ZBrk9bayZMi9g6IPKAVgaFXwGKpBfPNUlhQhTnihuR2hL+QQ49q+rYsuqIo6Iz9fd4sfS5Bw
3plVmjavjXmT39McKtSBdino/gU8USEEWDKo2HZSlTuB0PIDXpxckx8QlzTS0FmD50HQ/PX8Whj0
Wehrlnc8mqREf57k0sUGnImo2rAPHuKiSc0NZpX4pu86d5iZ9zGMb+IjKaA9wI97MGxoHyvTQo14
Oo+oITSGpYEdxbeNAyV5aQEORhS50QnFHpnfiSUEXO23bOv2/zWeGp5NQ7Z4QCRxwql3RUNHQvRe
fov8gwaNGcYr7v5gxPjwH/MftGF3qnihFOhksA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="I70omPehL0AmjLVWp0GLlXZHnxi+bDzgR6+OYgEg/7E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 105712)
`protect data_block
FCp8xK/oiwCTukjCbzefyn+Z8iYL9G8xETFCVmHGMC+n2R1RkhxMJOsYYbOYoz25IZg3DkBwZPOh
A8ofmomDEE/yM2BtL8mb8xOLdJfAa7WnyR5v/4vhKcctgQYp1HSj1pxtg3ZAwPTGoq6DUn994loM
gKF8KW4AcVvrTW1JWhvAQOASfCPuQGMIuJ8hPg4hvKXyflP0Uk+3Wz7yy0q3NsdnZOmKCSwnei6V
s5cor3YQE0o+ufZtxs8aV8FgUJ3bCxds4jGXUzf0bHbaHXdJlg+3EqosZehIvK3QxvBzZFxsLpHt
EMAiK/+YkSIyhoh5Bz2bb9y7t26DVWA9HLFnXMgf2cSKoKt25rtctYhpw9qImvBkbBv9nGTR1+Lu
CMPS0TqHk8x+LGFBNf6huF7vhX/5VpZqNm8kK1aRojethLgEM9qBmqsfnT22ZUZ+0eP4Ro8Nn7ME
lUfV3ElF9ImqTCepnYu3rmMxIEZ5Sqwd9ELySdBJFzA8JW+IA4SMjC0rWKv+868mQUu+wmt1+r0m
nOTlV0BuNKlXFZ4n0mzzoiRWBpo3KED7SkKc0OcpIp1yTd85hq6jwYlgJwSLjWdzYDLuEbMx+4Pq
pWoIvS8TKafTzgxgKCugcaXgSZKj2TxVRarn7uqc5eONtoThF55OLhBJUMUDCeB6RI57oNXyXl4C
/L6X/3ooi82Am+n1kKnjiaZ86vsUc7Y2J5irLpU8PhYU+vx3l82qekaK0jdZP0TV/BhwGrL3oWq+
VN2PT+HtZ+jHK4bKsNmbxBB21jeUY2EZ1tm8RvYBtcY2tkV+rEGo0W0hyh3oggXSR7KmMPCGaRPF
2Z2QKgsJE8YCTHAjICg3Epq1dd9AAaioFVnM5k714sm3LYrEHmkcXkT/xvwBQVOqnHVzfn5CLtxp
lRsofLtfH1RSHz/Af0gmz1OaLtKJsRs3BQ2FcGOiA0huFFkq21ZI9JcPZWemjhi0yVDvvwYfLU3r
iCMTdgsKJmbTgrklugfBiaQVRaO64o9PE1pxW9docB2q+pO5qk2s4cOFUfeEe5i+pRWbrZ73wOTy
eOKqGw3V2cZwAOhSlCpGdU5BsBLX08XhNeqCNzTuuaGSK+WdHaObuSoolweJNGIRvFu4o5BNwCSn
Xf6B/Po71BLIgv3EBMfATKnICuMW1XqVh86Ud8EtG3rtbd269O0sKf9yZ86nnhFl3Kw21TM12g5f
9LSI8tidyg8RTrGV9UexiPBYZ5GJmJx08Sp7UD3zrD+6YAe0oMNu1HlOGLloEEQOL1/dUGQthkme
96Jd9b0haxgszOOx3FggvIsX0Ook6Z0o1NExH0JOU2cakFpPbON04GjU/I8RWBCAuxLALiuMomZS
tMJ6xvRChAA3pdWhjqtUicO/WIte/hNCwklBvwnskTACXWAjV9XK0YFOniK56WzuSDOumR6e4lwm
3mW1qS8QMLeGAIvMWVBMncFAGzfjjvb20zNz4X8dodKDIxLFHMrOBjtKdP0NvpjarIAva0VHQnMW
p+PZPXmOWX3iYjVH2sXibd3Da1zZNISpiO2M1FOgz9FRw/wtGH+EUFFvD//oK7KApC79/TYUJs74
G0P1J9aeexT1BNlWLBEbwapk8zI/ZlsfBdYStYAEiggyArUpQa2impZTiWmnWUt1xvk9rmUxED1e
4LHJjX7dcJ8BTHO97DdPrCogNNHWvgjW0f8k1JDz5Bn4Qzv/bLNt4QQ5y0pDKeW1s1NDU37W0OAn
X925yGdSIGdWsFRom+Qkkh4aM1CtfS9VVy+grq9Wrxbp+87YgZ25Glo6K9EVIM7XjTcbsM4/d4f8
oIVW/12/ZSX0HX4c5z5wlRp+F0INfs6k6UAGoAynmz2IPGxEkPLCp7Hkqh4JFjZCb2bc9UotHVbM
1ZLc4zH0+PLw6K68JDcGB4n21B+qNi7h17Uso7XPU1UnSLHLquR+O0qqM8PXuRnwyE9zP4Ve8HSf
STJ0ktzEF5Zh62shzMruw7anvYA0IgepHQOHNsWkxUUf98mtKedOWTb0jKUMEQWWvam0RKeH7d76
vcFgJCcYYEvm9iYoNPzo/pL93MavJs1rUkn2MxvC9JI09H8eL2ItItWce6u2v57mnZ5gt8gLmgyq
E4J2ZeCMYDvIGY+EJyuaLRDSgkXca2cVA0BcUimitYPT8DO4mQAeCBWRpjiAmIx62Go0KGBRMrRa
U5C1bWi+g9EEZq8bctyr8zPhOG0+cUqfdxqrmcFeHBJzLeeA/99oFwztut+4pfBUBN83LE5QBHud
9KK1kwg8Rt9pu+WTr1ryEY3vPfJxORd490Inu6DagR39LKaSCK77kRS+UQBxFLFhBOApQmQcbolh
wZZSiOINeL10cpe3Drlf1kax8X/9Y6N7tI77IvHgPq1Ytx3IjHuG4SOTNEuOiCOaw3kSsTUIqtBc
zNgqhzZYADVP8+ySXpON3LK1eTy0qLjuMmQmPOEbC4JT6/MuvMSynkgyYLGZfGnKXGjVHfUhb1Ik
nqPPqKPxpc8Q9zRCiw+4e/RIN5+WrHwtIl6BWgqB8b1ZShaiKEPPtW9LnIYlJFgnaVbZckxWJseP
dNl9pSZVl664kM/X2+25IC9fY+78pYOLaDL/+IjK5V9EI45NvMW9eBvRz0qjFHScY6PmyAdqwXkV
EtsYlIWP6K0SimKTzoRtrSqB4usPlPezV2WIkb/Sl9KFjnUIaaUQAeRwUJaRD5zHhLrdcR+JXVyW
vPfZWUmsrgkwnwRVEOGU2RcvDE6gd6/BSD5dj/8IXaxiDCbeXgRYfNbFOHc8h1FqUSP0ud7szaJQ
8YXyppswX12FBGdhIP+MNzU95rp/g1y2zXVtiyUMqBwBr59KiaANmMvMnActEUOAfzfizYx9noJ1
7jDAfQtrxTCQgw87bgy3cqE7MOJG5GN20P0wloKamwOQizg9GxIS/6xYjshzLwcXyfHaKOGawysZ
otGwkrYTaYX5PI4pNoTqQ9rSI1ZQP/ZVkUUwGQjUpWFphptRzTC5Vyj5GW2ogy0+O8QT+SZ6seTs
HzXDVK4HjPIlwtONCmvsvgUK1EXQjJTdQuptodckwrJBpNqL3ydhNvFoFOy3HzUDE8qeClf9PGox
9yBxP6fDQtgWVMfAyAr86UJqtHAWbq+BFpqGIK+fzIOkkrapWTWB1Aczi73jiq2Yf3YNP2Dbx9Ac
cz3csblZdo3HNkZQUWmpkVjs/Nj9PorIOxTIwQPZlqweFLUFg0A1W1P1RLgy6GDSHPVN9H9NH4w6
wSNAQlRdC6Y0o3P75OWISrcU6XTfxi7q1IsAA203bjt/HEk71RA5VzS57DP8LeRzDbavERmBKZC2
zsLxfM7ATvczUtM6v5jlP03DMnxEfsPEa9KIo9c/F+sZuAjzQAXkwK5KRsUqsxo2Hk9C58UHQPXy
HdIXUhXWRQaFR2VTJdxvU2kl9Mg2v3k8KSej2fhqxgvJrGUtjd0wlCvH50yGaDYWHCnJvVzPAIz5
HIwtaidcn+m/s28pya+ihTOCifGqgMtoo+L7q1dpu721r1LpF6rUs0ajLvMfClX6bJiLIhmSS6RF
yNyuYjtlRCpuzC+P9mNrKXZkx43AaPuZ3K83RRvnBjM4P1AbJhLh4lAJvweFBox2sgHDUAFOqp6j
3fvoHngHlOW85oKVzsr7xypEMqfhOfDvSrA1GEOY140FjzsG1k1Bpnjb6bbHKWOahYr7qR5xz33/
kAWi3UrkkNkI9g41WLKO2ZWfnt7S65f1U34Ekgi8V6eAEAF7Z5QUqT+lCNpvR7d2xQcK9/db9juq
1fut/A77HsEDm51FmYKlFjv03FNQ30txFh7RHx7oT3hJYveKx5rxx3rxI8eero4iMaufIuAN6OvB
dmzU3pImmIgXao7t123mqwhT0NMo79Qb2zU8xv7xBaeubivSpk1v5+FRrkop4sApLtz0rc6hlz+4
vPofrx6j+feSUklLqV4S64GYJt1J47geDSyuSOpwa2ZG9NNrf3doFpViGu3d4ttQreX3njgaicTd
bxFyE5J2XKajZPIYzv8LdpurXRWvr4xOaMvyf3jAbaaBA/Eb/wxW5WhIjyiQvh8qdKOlzeGXYI5Y
vycRgaThDAxo0D/T7aHp6m5vd7xI8IvatqH9lbwOyyvTX2ldsDnrptELcM0HSSFzVFmeJpAP0sHo
JcQZbV8pS6CY7cWLoc1hwFZlqF20EnzZtqr3suYKoekKJAqO6QQLZMJrSkiReT73Fo3POPcC5TpQ
Go0Yf16zq5EvR/sdtXhQVwidzUovQU4TcU6mV/cG4k25lYGlsGadhwro3rrEJGNPusRa7d2pbqTS
/M1yQT5tk2qlBmxKRGHEx0hYzi9Il41m2/5HxouWGEBuK4BWR6YFm4lhYwosKj4MNeOC2CG1G+Qw
prlLjOcPqo3Dh+x0KgU1ZIfe5bRdkKTwg61naozhBfDwcXjcQIRpjSX5VZy0xIVh8xVh+3nDyOg+
J/0NH0R5g1XPId3CKoVOR3PedxVtFG9C5ikgpni4u7F5z4yH40zkmNasMnj5sfEGnpcxlVQ3syPV
uqpzJJq6mQKHAdI9DvcjAC1Fi6eAAGWmJGsGshO9u9s/D8jombfcaICK7W+oZc83dNC+AGmCyaYe
uJ+2z8H0elJ/pTSpb/2nrmPKdPJXJ1mZYShR6wGnNOSG1IYbmhNco0LwcSO+aEHj7dmGzFHdC8hb
retXEcNjXN0AZcsTXQbxNXpfWJwveyTJJciVHCiy67jkZjnCfOBWahwLYnn7pNmJXadhuECVTNfD
0dTmlFpL1zLD3Z0kegc+aBlU6LLvYbGldLes0Qf4vqUBK/1lC9XMHsoDzk+y2Pg0SfrOC37Z0+yZ
jxdU7GM5+cndXD219vhNIU62wLwAiRvd8cWSXwEsTzGky0so8KUQeicOK/o5VO3M6PKXgZtDtm/O
MP3B1tefTK1PqPmPzqmOxfXzn6LyGcTeKFUOjRzMPkxrF8a+/6NkHQpQC1Izq66yrWC33tFxVCO2
qFjpEgIQtVNeojTSUZO0z29OffIMh4LPyCLNMiJ5FQP1UVW7EoLHjxFk0+BP3vy4W6dzAoSEFANO
0ipea4YffPHAzmF9Cy5CHoGwFwwjb6dOV6KpGWbq3CdpcX2xhni+1tzNtoZY/9e47FWijeLI3DeB
m6sevzsuo3n++VeWb+dGlCOiv1/KZhIXNzA9KQBvAfJTv5MUz3cNiOoRn/qNKU7U65RqDOVPBM1c
HyZ7cg2L28qqUmLOYGjI2U0pGx6f5htItdjpvD9rhhD3jhOV2jkCY8dpAyqNLT/o9C/+AmRWrxnT
yXuc1XKZv6sPxfp5p7oLCaU5j6no9p5EqUi4c+jab489f0/cyNfHgGCKh4T8uaVNsB4dGW5OFCdb
HzEGCFeW3hvAddue2bsMycYWWuJ17ZbTYRAARPHYSmj79GUfUdXisb55QFPLglbtPQTk4W4MGYvd
jqkhJiAiTnLmiGt9ePriyUDjRw/y010tO7n1gDLUCpm+eF+1vLUeX7tMl2M/FfpHY0GmIxAZb9/G
YwWDP/gdBAIqoF5NDO2LpRh77A2BeK1g17PO2aP7/EZGjWhhZ3K682R44pdtNbRHfOM72GXtbNjK
R+8DYlYwNeX2ytFPxXX7z7VQ0GUbDqBch1BBRw93AkmxeN8HqSW9XvAi+R27n+y4oy5D69JfuWdJ
sg7b79Akh0YqADx7+JzpjTpO3FtiIbDwcXfh2LaJhqRyV1ALsOY9YOckqX3UVdKbWcamg5MM8fJu
3yOxT9oZMaQNzS9mbR10csObfw2OKWOq8d6zirugvIPFK6JQWIfU6yi0rDzpU/b0yEJwEt1CVtnh
Xj50qwyxi3r/culRTELmdO7wmaVpWsmdzhJoaNyVuQDnBLUHGBB0ddUTkcMl60zAwUEZn4HvbJdo
xHtyzOdNkClLk1ai2ig9daNerIZbqi8hHVM70I+xNNvnSAKXfw37kykHvjSj5rBp0xMRiSprXrNN
qbDzRjdGGiEj744IBjkfuCd2uIlQgUthlUy1C8nDMf3Y4KkxIayvdeJ2YpzabMhp5QjXdJpyLf3L
bACYu9XbJrqOWGdCZBG3NxMv/ta5mIZKosJi1D4QxC99MaB1IVEIOGA6CwZAvXJG4jrbdPLjhBbv
wdwrJuzi9ADe/vzCSfVBj3svFDdmm+O+lQ+tX5yf3r+1GtssxKrFZPA5r6hxtsSyRG6stMSytiQi
d7LEdrKGXZ5U8WdI2QTLa4YIy1KLbhOaS84NhOVSdJFpAC8SZjS816udSiwieWaBqoyuB1dPFn5E
cBnBZzyfbeHJJbLJQJyLmlSoFMDPvfaNMe4K/SIVdcL/aMxEbrE9eXHROitph5TtvrjEkxw/xnqG
6Em228mYMeSc6FR+9rhqEQ2qar1hBttMji5qAOTuJ6YJxwk7V0EQeekbq9Xe7wGAIPv24w9zQgIE
HdV7uUsj3VaP6MIp8u0EEQp7ZO9NIRBEgwgAlamRvU+u112ibgkM5KY/IRLwqjwkejXv/iD4PkIh
wjC44+cTFkek2RiciPBcpyF6+Rj/1/DHOUlcuoCwopm6KwG2LJTyG7pSgGB7RqJYHR9UhwE/K4uG
c/mex3ZGQ+T3PtTIBH7hftGFp3xNeF1hVr5yv4m4gXQ5yDrQtLkijF4S18m1ZU4GRwGiJEZRe+7/
rMEn3ER8S1ZOIYSC93SOHQLyf+W7HAjU7rESZ6vE4S86PELt9fXLQR30pKh1OMd388wa6p05htLs
aelReuNSYiKMKRQQ7t0ZM4Kif1nNliIi3GJ0OknHhWGq17Dmaf4Gedid5MA0fuNwVyiXvqc7TRMA
Xn+mwmMbaAZH7i1q9I6iPFBMTXhKFQdEIAUBOSm4/tnZumanQr1YtqlWhD60OSEJzCNBqcQqcxMW
2f9tcAAx9+ytIvTu/YX8/JgkzfspQn7As8nl3Y+j3ZfUlfaOvQ2X78Opc6VgrLE22BV1Iw3JnYl3
4zozOcD6gACSJQMzLLgJIo60a6Y6IhYXmVla73y+33QPIQH3Di57bbO52pSABNXh/JU5beg3h62A
/rIG7BGig85UNY4rSyPfG3rwGte5TSZtqcbUVBmxk28zHpSFCWr16Z3aWRPbJxf5Igt/OwoeYYjQ
+BU+V+5bDvQE3wwHrMh4dd2seSBf8LKa3sy21NU16XIQIphSZlIgkk86P1J+oB2t+d53rK4BTgI/
UO9Nwfy0tFQd53RNB9r7Azsdz/+Uimi4SqXGTtZU6sUE5xmPRu8gx/cLWyx/A8DG3fp29Tx7P54i
LiVIvjVgHyh6/fqyXz8lKaPmHFsHpaokL51N8RQxsFpdlLnP9nNaY5OiM+SIlXDNWJvryQOiM3k2
uDsvM2n4qG2doGZAbQFGSH+Fs0F9NnzQNIjIWKpMzSjD00JU3VtSNKtT3VWWoZjjlcAdv4mEuiVD
gl+SFVL9v6Mr6QAszzfFkcmM1bCU2qxbPlfgG8ILFLffwIerytwmr6ae/i/z3hTH48Te5TyrMvCr
ZWd98X+XJlwyeRRU+BO7Agq1jzF6unB6TQLSCRgg5s8KI4PDBH6moxdLBHfWgjEzijzeDgLN/6RY
TPr3CcDBE0aOWXToBxxLBeFf04d3kezSWz/rJsg2RaVe9+w8EuyYYJw9qL6tA3KgoKXInwzl83ZG
1LUEPZ2rtLZL3LYWiiaG3ydSbSb74b5Pqo1MygIq2HVaF/fGGI/QQtD/mHhlMJK92DsJTPP0jWSz
s7FBZwUSuuKxGJCCHLEmTJhZ80PF5takyTlvM6gXHV4lw9YfPxDkgnQPgfSth9osfpVzEWAF/my2
rb2dBRzWDTvVcq/lCIx8/5sJ3s4Si1/ms8de0K/vGQCnePqysn/wb/L47JKRc91wLnV5x3gOrris
SUWmoqG5YeP99DQSIaX49yDqxja4CUGwWq4kb/faBRgorfTiLKmWPH34cgZ794GjZoyrFA1lAwKs
nicrpLc82oeGZlDlV1Mu5TPKZrsF73bspuSybm54bjJ6zvHHspV1IR2I+760VxhoWKqv88AGqBrU
mC4kW4tVpg3a4JYOQrH5inqaEHARUtCKIE9oSn7Uj/qLCpSGSrfYQ5h8HbYgiLVk+pqHmT3Oc3dX
OZS4LQWpUY1XehDyD1+0tFkvHEEMSiiB694CmS31DKvTpHBXKQVQknAjNdqeQS29QnWORvkKynhd
PJtj6O+Tu0uw3exvPnIleChA9qeHwAghZZ6+ZskJddKOeJZ9MUNyBRPQh7vR0tZPsMzkMPJuKstX
DNnD7+sl/S6XVpguuDl8JRNtrwLENd0+5z/uk/bHpAibltzECKb21qbVnWwxGTqu2Us5OCDiiOKl
+VJ1opwpAKe0mRU4ljVDW8KF84FJj0OTW7a9QM375TQVdvHhXBEZ8vFYfntsc1E8naefiuWdZ5jo
cC4TpCQ2grOepa/vbtBRH+v1tvSQE/SMV4q8nIgbDWEWT2U1yPC5t5yEEtW8yJSMjjuxLmBDRCc6
cyTpIhRHeSK1a6JV3ODbMwpOiy8exFmyxMPX6z79sv7OyHeLOtvS4sumoSuH1CVcXq7jzZnaEkcX
9l7rgDejpUUx5XaLOTzBTZtKLhOL2ZovyXwqUUH32Xx5axYfpNBI/s01yfxbvKbYkC3mAh5QCSzj
zvMaIZhmcsSnhvrQkfeTNZ4eAR98THsyUtYA+UDV6LNdC+2anS9W7N038ijeouf603QTW5EF2qCb
XGgzBmBQVHPuH2ynhgV2iuSNmr05rd107ZFFjE27oyGLkd7Bxzlfes35/OdHd1aaK5VoK3ppdlFP
PeYRgtXg0rFVbQMTrA+PXxzdfGwVrL7IPBTokptkw7ZsHXKvPmIaPPreAHXbKIwwCDreTCmDCOHN
O96e3tBRH13FHJskc18WRabwMAUoICrrM93ABYVXwLLMCUuOqlpZu3kkYM4e74UcWjwYodJXIshe
C1UZCkPF6bxsRN/ud1ofCHlaPbOgLov/z7gBMLh5fQsl8VELBabdMivepjod5z9aEHh3mrTYSwsi
epQC1VsEZuGrZ53HRrHAxY9Od3UMr+niyBHkGA7xCe34pLmDFCeAFWq4whzygZiEUbBLuMyAV+Yf
D5FrZH8dfks2RI/WlIYRWIZGFo+tvLXXfbAITIRwNO6hMBeTx3oDizU+QuAlJuj9Fxv+Gm1/thbG
1sCbJQVOp5R0PMhPmemq/5Xji8t4yToKauN6Vkc2ob9p8wxXyUSOb9LTPG5G1fipr22cF5kQWyHq
D4TtWkNVi76Wt2R2z5f/n1gw3HHbo+QW8KaC1f2G4v87gPGvWM7YlluT+//g45MRwf+3mqp7VwFO
MWZidvZCe0pOZZJuhd7NRvW/IS4eHEwnrJj4MdYgcm9t+wryI2wSKG6/YomfZ4Yz0CiNwRaVE8ac
54rDhKva0r2AmJDDckRUsXjpWGEx1wCAYpVuR8MSt2JgjPhg1pnepBnPnpOtzqgduANylPNuych/
6IxSHtM4QBYQaF/bDW2Jw52UpLLj0QlmW7l/TnvHSdBSsO3dYy7kwBVU9vjoqoajBzgubm/IhD1q
amiJ1XUQy5HKdugmThSnt0aMwp36vSp/QPGPuLmMWWomwDlZcYsaheOF/Q2SySVGo5gJi8Jvusgg
aSLWLvS+5prZ48KMJ5s89yUzhTcyM4TB90wt+K5mbPs1qqO+U6cF5houwUhSE1590pV5GuIUEWV9
TLZ9KwmRuhgMrfo/XNvmTTVmGfxP463pVepyGb1EXrjtZvHePckqBCjC9I9KK92F10c3m/dxnjwD
OJPOg9X9zdcDkWnuHp9uIwPYAEslh0ar9Ve2f3FacqwtaJm6IzfaXZALr+WE3/KQeSdc+ba/ipYZ
SnQHk8cI4KYdgqepNeKOHSJsm67T9nS31YQRUUtALjlnej511gBQTezT1OXTKzyC1QaVVuRKbeHA
JFt7IDRWH+VVPqvlzaqEStd8WhHwT63C7N5+mualWMSbfyeK4vfH9+Du6zJbRg0IFFx0qV/aHYSb
xTBViyNeot9wH5YV4ngg7yKG9Yw95FAmtUBT9k7l615PKViyQbWvbx0MrC7OmPG4wx0YnEWxoG0t
pbS5TvXvjofmRkokVTHAUNkVlkCHkH+0C6Ns4eEv2Hh2YRNIw/S0/57sDos+MaT19KLxHbzHxgJF
fdFpKIFcPNd9YDSQ5lusbosLZ+FduGyUuczGWASUmiBavh7ysW8APgbiYUpsu4t+wx6kIo3bAn6u
rQF8z2lMNAehifoWSkmbShU5ZwFcB6UE6yAAPNKFod0OLBXi4sc+fFAQeDLOjAr3czXCy0B1O+Vd
hjvL9+RtLJ4uZ0L/89kz/gzoLn/smtRAhkprmpyHq65M4wzdmzazcaQO0Aa0AbjAX8IEL/W19IZ/
TycDeYRutzo6wd1pNtPo6kLiNahPAih1cuI5Yi1Wfkpl/ODzt9YIx/tedf96XO+FKDfmSgZEJ6Yb
HdKMVoKjMsuxB51VtCX5uAJrRqW5NPb+OpnPYQ6TGnFD9Nl9epD8XoVGJfErS6G8RdvSfpP2BQJL
HdwwY9iLcBVkZRFYODWTFear6OZuuM1ySEZkgX3JbXmltrsNrqKfj7Cqr3hTDfzV0t7N8QZ5Yl+S
vd+tLf3sUbq6iGiMIE1EhaF+zlGcYlu5WiG3R8g/iH7+Va/mMpRXKfWyZ01HAtQI6GgjjpZXeAoP
pr8DV1RCi31Y9EaocrNgkTmN2jUSc4UzEWhAv/gqwk/nG6OjxBLInX4mAtCVinTtcIATIfFLFxwz
wWWrQmqfpML/TTytBo/6rSI5XEnXl/g3tya8GMLmCL19n9H8jGyYgoa+2MfruX7vS3wsUy5Zvqph
Ms8NrYZX+HRwiLAsrWt78sZr50c/PE6S4uQOk9b1Ex0Z+pilPTsbST44psKu+dBjFZl5yMj+3D4E
ajW5a89VhrTSZmjbj+WI/v4dR+dDueHHlWYSEn9Pvbc16uozoQNd6+tVsoWdM7SQMd+Y+ystaBzO
9pVdHGciCJk2B771o4kFgsmMOXJal5UXMOP9B8PiTcURWbYPri/dY4sT/no7ZgIDbDNaQOo+fMLC
pa4YwXcrKJMSjyolR08makhC8gfLPMe+VEygejHI3aetZWHtopNdPwksFGYi32/bSQ+C9Zt8fqBJ
lQMSmnDPXeW1XtcIGDEyLu68nt9WQEINlq9gYKeHXDvEL3wpwhU0vnXJXOCqsE3Yjvf5+p6OJAl1
nAinSeCkrnZb4NZYDUr/yvroUMcCFONfbB1BA00r+NQFP2KHCaTlDXbvF9UgBBzzdnr650fkoU+7
N5swPcIFRdvpBbmRaODJrwy53e55sKykH5+YNlBFwV8aoELN1uyet+Hsdmb87rmJhnjb7WSgMRqj
Br1fSviWtDBAPB8e3nBCyeG+a6NnckFZfP8WjfWva41Khbbo1kZU42DfdLzGNrf3lJXu3SGYTiuS
5Dd0I3CJW9iBRREv0F3Gfejkxb9z9jXLHNHVQjZ/yfICiAPnT8aLNcANl1mjgJ+L8VsruyBbyb16
jx3F5J/HnaYekUEvqV4/MFixNSHytnbprFmcHHBuPEtJpKPUlWA48nJqWft9cvL74JgMuHw8Sr5x
xHpsoKHVH4HkMfMwaiwHf0T9Mk0gxzIaZTF5V9DMtu7TeFM8g8026LcBtMWu2GYLLLF3g8w33+yg
XEITwcCUAmQTFMVvoWwaWVXmMfu4SSXRmAUfIBMmzhTbXD/pZHbj4eONUOSmNEEhkSa7XlmVQ+kf
2W5GWuktW13wve7lOFPT13iP9Az0Sjvqd7aMqWj1pcIeTZSIxZLXyD8yUl4iGMzlcAAhScpY+Hwi
Ux8PfmCLfWgwRHUhaIYqsWECmdZ3z8X3QRv+mR824q3zkH+e/pbFaQaB6NytwkNQEjpJ1431KmPG
pxveD6eXrb1lmV5gxU8asft0MNSi9rj8RirxQHkhyT9kHZinKfFDmk1huf+0Nu/IKP/aLaRRzwI9
htF6zDyK37DABcx4klE8Cb4WSxYaeH4EhlKSXf5/aJCl+8C2PAEBLQQt2YTYdOhHNiosV8sUkG1D
0R8fTQP5Exz6yuve6NnMq6RwphmOAdvlrvIDIy+9Cnt1pkMF5scaWGbp18y2FGcMjBH9SN4QI4Ty
YAO3qxuOA1qY/2G9ApDwJyVlnVrtyaKRJuWZd1fgofH9pYwOhxmXNnSLnnBpwkMeyozrHx0cBD+3
V8g7YHby7noW0CAGdII+WitPIJP4hyp31a4jFEPS4M8BWCo2VMQZLG8n+Ixk1XZGIRCBNkJmMuh9
fykRvQel4wYKfSJJzRat6B3cYu2UIUTWM/JVKXuPWgu1Jg4AIaE874HmTCe5Whts3AgHB+LMxnU2
8iDQUD3B2yGBpzmyj4LlHPqlAi9CB2yRbQ0uyz7FwZp+JVAvg4XZVvltDfe344IHP4HxGSNyxnBK
NDfK72hw62Z4ZJqjqT3cT+1Ut9KP8yhWlj4p3CO7XhFiUoiFAJt3WcAfGiCx+JXAsytTyLHR61hF
us8I+lSVAixcC6YI+Fe1LP1JB26QmpIqDms20HT/sySzdluWxSWOocqc3HXObgXFOJ9EepuSA55h
RLeIFpTsG55S89YZ+hsW2NnQJ3LFoSVqYqroVjm3reKsToMCdbPTK63IXkORL0vD3onBmopMFkzY
gtnyOVaJO9J+kcIpcdCW7OahxKN/Hatku/YUhbAmxZVUNd0vN5o2V4ScF7ZZiyvj/+pYOrw2nHSf
lpvHS5Dq1r+tQiQ3e6lqH/LXnyq0vl3ivgLqRL2Vn8ha7KJw4vhASvdTXsADkADDC8NKFSsNLk1x
embqnmDU0Upq04oY2I6+9ydr9kwMX1VWlA0f2SD84B6ivWqX/hkoFK/MEv15EUxf3CW9SV5RtvKx
8Qd0ZN2qnIn3EIZXZrdG2Kuz13+C8c+oOoCTduxgiGXyiN1cJ6CmmOqhTbt4Z/+4dsFtAlbyM+SH
NTAAE4lU3/3WEDTLiGokozKcBkLqBUJ6hZySri4mIpTNcViCxkIKRftrNuPDD+75eHKCVXfF3N3l
dCqhjIZ110q1mzkCoNC7aXLHDuUGQ2x/csGyqBZcwTW0Mej0tibY54JqwamhKxItZ1hwhXGYFhPn
CC1LXEUaSAlTRBQ7iIMIgy6L0ZwtWhRkhTJz8camjZTUvP6NlAX77+zsdhqGkOmNmU4ohNg2Ue4+
VqMo8FcMKNXeqwx+hm6RTWVfH9r1w0QkIuaRjl9ioxAmCgOskhCG5aO1vNXy3fbbzRmJ3z4+TVp6
z8ebHfuWs1W/j5KkPy8FT3RqUg2Aftn7Udcq+eM4yhIuwIEhwDF/h9+jogPTfj6T9InCTfwQ7Uwa
My1g0sIOOtwiblgHyc9Qo6jfrMT8c/UYyKvTj0ORr7JdK/rLB/DxDT3VsLFXHrKtXSwLMZ8TKcdF
uqNuoq/B0JP0GbkAUz2UJZGNuZ78u82Tt0H7uX0PWhGCDUmlB7DLpvA95QlS5tjmwWNf/ybJXwQV
P1MA6M25/lolpLLZI1nOc4j7gE3zlxIAAjOAcN47j21W0UrxcAyYyoKkvexI+TUY9GCbvnBQ8xJa
tVpmvzsknrXXh/oAAcIsU2qFGESWY972QgqLjyV7nu3PK3R7PUp97uVUL4P15XAHhTwUGyPeeJJj
8dxHGiTqPVVB1gt6JbWTtFOaus6ac9NPimbDMLs+T68RRd9H22yUy9Iv5B6621FSZ8Z9Xs1BJeqW
CYnKwS/xwspzQd1cmbe8fAfkD7ZetE5A0iB9jgUAenlhN4GEpc3Ye4UTxSVPRBMB3XJYGToDPvTl
AiwC5RLFWQY4TPkCTQxIIHxTt4iPZx1aQNgwC30NUw2y+Lp4LGxpXlFXBVKwjhE0R6wo/ncSqOH/
OyKiQzSnQxA9M01RozOy6EMV3EEjNXSdFyonA0/N8eKfRRWEAYEU+v3kQvNa5L7U6Qg43SGGXRMe
myaaIQWzEra8xJy7lx367Dv4EkVJsLS80jx+fGMeWmxSEu32+kvlNoR1PB84jkrKD8/u+8A4bruL
M3iiFQtGuvRYYhVr1ULihCF4rXzwMqLI3r844wkOwdXMNnsZCCalkNTvvQe3F2yD0+20IWSNy9FC
npP+mzzDuPmOEwQXiSkiGmh4Wq06NSyrys7q8HMdTD6LNOURn9VFI4u0+u/h3ouNr+nrDdJsrVXU
8v/0Nq60lPqRk3XQlCQhqvQedmzZJfsGQxYZI2nmpE7lWIhJA0xKhClUwoVQ4ZLqPRMiVBuKxJM4
SqodxFlta3vTosS0dlm2n/409vU7iMJr6PBUnDMNiBlJiUwOyYAJ6CyzIdqQ8cmZ4/ivNR/xMQcS
SwyVlJ573cG0Fi/CDq86J6Jfu5IA8CcVbbsXrIFF8gQmtzGSCxDfLZmgIMAILUBfMqOS04RUl342
C60baltYYFx3/tk2/s5WB3AskWZsr84q9b5zOLQ4gZ7nqqYzXwHQXO3OvdLTRGu72HpaL7JERXsL
uyoBtaXTjCATjd8YWDi+i7C1kg6JBBNKCzfJ+aVTZzl2l7VmzKq7YtSSKyJcih+OkUegDeDyJWW1
tkbqzqcnzOEVg51wkmWwIjkIItkC2mI1anrrCiV85yzf47Q0+oGSrIo1EevAt80/GPjTJpzX8KTP
pn8RS5XkU9cOrQLc9OtHpWng++SHzRp43NYQm/iHd6dQ8jcB3r/30ccJz7O9BanUggEguY+Nm6VY
M3Ja6h2CxWXsVzgfxhkZcLmH3FcEV/OH/vDo+Tcs5obWtn0viIFqAFg6+2QiK902JWAoAUJsecrm
u9Iv1NS0mOWHrxv7vBEvp0ne7whTAbdf99gsab9Tm9EubYnp6v1PYKdYJDSypBsV/BQyDHR99TXF
2bULJiXXmX5mujvh0967/4HRy7uYD/OER2x4oiJKX2DGp3oXiV0S+TBuPQK3x6syLvhDxxS8ZFpZ
FG6Zc6IZv2vaKktZaQ206ddNyfdfKZ9U47z+JQEMjc4JQ9HvULgjZNHJ4/bJ2vhKXWHiLUtnzLX3
L9iLhhWrgSgNbG9yYQPmLOyavz/40vK6QyX5lbbbHOLn8BnvM3iCoSKh1Qyx2YPgKxPGK/EDVNWF
xJI0WUhj5nHY8zq3dEtVUQeWddMZipH5mPQDwgct2sZIEpKzI81el7m3uxsGkE9X2Mj0KeOTsbkZ
C4c1lagF5C14FP4gN/FtghQdaVJKb5QUslgGtbsbvyoJ3YvnPe/u6LQAhkEXGb+Dl/JTgf+mPwrF
wDqS5cWVwKvv3d524K8+xRwUHyrZMsCotU54obzmDJIiK0DFN3dM3uSKD/iZ4kGA0k0t1tmlh+zP
1pa3oemo6yZExOUYPOHG3FfSM/CwF9NimdzRHN4BF2bNgq+ZqvaewHViZ3ZJhfSoSO6ggr5aIegx
hADBePV92h+29rR0Y1nyJOY3GRLhL6++AOgAVHvET5jzRTfzzfAHRtPxsQY0WKWoXd9zEfjVm5oW
bk9ItBimhlAvxPEKOJi9eY/0nwio/t7AjvjSHVwOE0KQXRBLc9lIt5kfMvq/442WEHcq/ETEcGz6
JdYSm2FpT7WtTqTGH1uYXw8hZ2K50/T1XjZ+OJithSYUhAS2trXhlgNVNJN6wH0YuTjdgR0slKND
q7Iq1GMqAytGYE3+12nH/5DL08owdyu+ltykvA8wgBtqkrQ/106B2MErtcKyGtg8G4jAAjtr9/gB
NvuxxwWGyC21/5jrPrVVxfvWqMeetKa3nbd/+iJTeX1wH2ybVI/fD6eh2U53ZpLYd7RIxBcK+5qH
et1LNCBUMH+jZbCkNeEBTgezyp9OT++OGn9HeIYgbZv/h/hx8WF/Ub6HSOIihKlQq1Y72WSuxndF
yBkrB5If8luhgGGz2dEQ9g7tVQS59ENgMb+woyWSCGy2Tj35i5ph3uz86BzF7fFePy/5TRr0II4A
9Qr6qn7OPsGlVe7TX+yR7/p3+sFMhLdYXhW7+HcnYabVbfaR0I0Zkpf4JyGhX9isqflSNaAB83N+
h2DJ6R6MhhNAvGIY5+cysLkrN7TJStGHKJDxRwjHeXA/k6HKIijBq5sXaydmza3Ffc2/0+fCsos4
rJXQDQ+UsIdLfGZVor5SqmqE3mUtAUMoz8IXWy/Deb28eLVIhC0XHeMCfx72MCGK4DmvFnoNj6m+
ZN610iyEpa/fscWXDq3JjMObaFDCsnLG0csilFQaU9x3hnx7l9vyNWsclJWgmzS9YZm+m7ZgcBY3
0fH5rfKrtQOSplMhVzskcIOJmoc2xUJFHjEQIyZDXe4/Z7p8luzv2G7xLDKoqc0yXi/Pdxov31pf
4yEIYuB+Bpsl7RnO0R9YZPP2Nvj66pyH2Byfko9ehGySUBBaqu9L6RZ3O5xNLSYnaiK/kPImTRbg
FXip/tJzRN0N66nfzoaPSn13NdNNiYU+9enTX03yOyGZ6ahn/BvGFYPXGoCaWgcCXGJhmLjcEL3t
ijBEkFPxJflwqrteDlCHVUVXOSt0pXOUzMb6E1s/r81JahZJM0/RDZcGiBGzZDQE/c6XrIiTj9ZI
7PRs5vTLgnNbee4BUXUhsIfr9ihcD6cK77iM5k01XwLSJsQ64GAk+CHMpXeMyf0BIqyqYRt3shAL
suIbXUz4xEP6HzUDd8g9qcLy00Fk1yXkMWc0yiS2QCxn6/erPiKWlLSE4JEjlmawTpDGcVkMUeCI
gCNlJsgwfhu8/nynaaPDK8JMdyKlnT1MsqkuLLW0KygRxO4hcKjHAV68h+PrTA/UNTuFtsaAii4b
FlcS+EwXK5GHlVJbmRBHbAnzNaq4IAxHIoFsEyso249TKaC1Ll6Pyy3+8Ka0NmCGWVdji8rpmqfk
IyqcjP9Sjkk3bD8H1BuuZsCvM1/D4/Y9jniGizdGMEXpHAJKMpWLtCjLdGObGNi6YMkjPAPZ0kHi
6ypHDObio3dSRF6R+AIqz2Hysd34PcZZNZ1jm14UHmXl6DWfPgE8b5SP4k+ykIw0YwPFFYPpffFO
GGqMNM6+ipl5I17Yg7xz2pYu6pBNGS5GLyPICiDpUqGImMnrMdjfOd/og4871odh5KajsJKkIUJa
30o3DDgjU0XZKOyZxiFCBCMJN7pjPZNfrOgRhkY2OHAyEsMg2uwbQFYNo6sz1HnnFT2xwpqAsh89
O10T+lRATOyK9RQPSYUdFFvhM8LBP51M4/BGsA2ebVohU9zB9zB+I1hFzdh/aWPgTlTceV8DtpdV
B1Fi7WQLabiNSZx9WwEdF5EY6bUafy0nnTslTeae90/cE7OySmwJtDwIkwBv7Sl9R3ggHdlWJ7mx
LdLUpI5lCT+H1HMzxxk9mltO2Lzh1SvFj0brwFARsxFc/NtM2+Xe5PtN9PL+yt0guOKEKxuGvJVq
CL+rMIGAYUNaZ1zc62o8M5EnKbwtXwsCD4vtdoQiU5IUjUPPDkzLT7ZOqJuvoFfaz78nFWnOpatx
L/LPbGA4QpkCx5cI8kZnGRfiava6zdJ93wsaM7rpMgUMt/1EUob98oVfWkfy/nqllfApr4vV67Xa
EGYg631lcUwo3haKXgS7eRuzy6wP5s7zR3JEO8NkXRpMQhPhuopZYYi/HObg83F5YmCa+LUMd9ci
AREkHWbgtO2uDrAlhdoyKI7fYzHgQilYGG6qQNr5PnTq0cmQjAI1928pjkp+lU/M41oR3pGwANyH
rQ84jMQdh0XMDwUVKxYae2Sd0IZh8ZMRjNQs8FmlrdKp+CL1Q5vAVnoiUkjL/f9bu5drpt+ZDyk8
1M0gZSnFZ9AsnesqViI0PkqYJvaYO9ptxsMI1ggzsOHdVCrZlmdsaka2WSTiP3mFjm6fZhKLPAeM
1zf7PzdcjxwZta1QJy3gp7ueQbHvC/NTBMp0OdZJhO+TgTNozj6KE56NC0Z0z0SnT9nXdn+KeYlu
yT/jdcvEGsyUuNpWWpXlE/r02sx0i4OcL3gCtnwOls6nqwGvlqL2TtDTFoBCw7GUVDTBdycJ6SS2
cilz0Ss4imT/YBtNqb9KIZIsfnQRYrdotk+5o5W+ff6qY7cgmMBvHPzsb81zLE+vmHYhPm9FiO+K
wkdp+q8XrFPus2/LayIkr83tBKG7FfBxdfNDuBBsYMzXOxvzHYxo2LoxSj1IsbIUic5vFndlgATo
0C0yrU+IFxxOdfNEGjdo/R85UoiSNIR0EqYt2r1Qp5cN4LNJHZcC6LJhmApH4f3TQtBvOBP4Z1YL
PHGjyo993DjOI7EDUUJQLhoEDvyqB31GkI04QaN6gp2/olrO5dsLYmh4INtqcCRHp8IuZl1bGg8C
jdTYKnU1l9ClfvamFC1XExOgaJOUtX8FQEC+MlTd2BQMQ5gb/64Y0QF/uN5SYs+dmNLHyj47lSVX
mO9w1c9KoSC2dBRof88y0HZvh/odCNEC6c5fxJGjeYOTpJBh7jWtVAD2SiVcPdrIGylwf62FuvrR
J+hcIdni5MAQ/UnRQAW0RNlUn+EK55s1wZ2CNnZw0caaShlHGHpxkF5pVkD72KW3UMn0BTO1c33K
35OXrXu+7rxqkbB5aly2msw6RioYwAwAU4q+4Wcn/Gp4/wFpiZ0Bj3TOA7eGds6s7rf2Mr8fEF0N
ItOtFtcDqifwmt/l11Aijw7RNlWCeyrHXVn6jqwd1R783EAOiMi/4AkrwgFMoGiUmvGs6wBXA3nc
KODkQYXoTYqHQR0mkIMno0gZKWX9TI/vkbs00CxHUy/Jf1rxeSF9Ou9AjMkWcjTizstMXFgNu/vn
7HVgVfhmL/eIhEuvPVvo1kiHhvDYp8qWs1mb7NiF/gRWSZdiGUfeTBpHBeyWoNG85uXn+MG3N1s8
Ah3Z6W6McUi4/71NtRdtqNeYZfWIFOliLSchz2a7pCAkwD1XiZwihXfh+DtwC43XEWHgURS8J/YW
zKV94naiOCtaFlwXUfbnSDed5ozxEDRxETqY/7/JPlFokzaQM726SJWZNhs66wYK7cEQp12MErUS
IsFlWXZKGUaRpCt/xu4+ejsnqHxFD11deiHUrMw4Dt6hV4HHfTv2Z2+U2fX84nQNsXTu8nwgA/T0
Jn0oX/qd3bXVtdB8SFvD0uF0M3ZUmv3Ld+QcszNMQ97jQkIL8ou/Fr8fHP2P3ys87MTTTUFkziTM
twMTlEV7DP0M2QnFkY8mU/R1TVHufjDYXeCdcgZhAjDcR/oMgEZ8Ip9QOhe8ue0EQy88BKM/yDf+
H9gnWUDiLDOd4LBQ437wT/+g3mXAGVY7B9ZBmLy88f8GGZegMmK5wQ0VBNhdle0ycWNCMYUTgIFW
prsb7PObeFQ2IRCohc2mNQ1uXPI6IBxAn7PGNferzDk9HXx6//krDrerNAWXi3zkbuRbK76xdo5x
1fkOVR6FYZTLWiBD7lzOpOmbhXxvIFZc1/jxlP3NP2JH9p755ngk1hcAzIIkVeUNaJBGl49eD5z8
kwrUlZ18LLKDQer8NaZLQlK1Rqbm7o7OEKTOKJCUmOfpNmCtLE8P0uTITFh3jPiT/5sIWqZDpRvp
WghrXFh5r+gqcAAS8MM8/UHe6rJ9SpENwTvHD89jvfTIRwFQABiYttuJ5GZM6suuOPo7AIQ2uJOS
rBItRW3/84Q24WDLZbqTif0ICeS8NT3xima2P6kWtR5ve0sK5BNGYrQz2BleXqQ0DZ5Y1F4CefwG
iM0qV7lt4C7YtH2KXm5nJS/Pyw9U1r2cUFvOBUQRdwvWrm4uijK9hc/ibEx3MGqfUjXa8700lXzj
j9QjaYN0Ir5/uNKZ19XIxaPS4I1Xp+02l6HMYLL4Qitt08S6lgrcjdyZ3W5Pl4eBmh2Zjy7lyMOO
Y+mBnZTIU43btztj7mCqslo4WmmYQxa+0IBXLfB8n9xiKtY1WaqT6WdF0GSELUE6iSV4fAkb1lUv
QUKH/7tGbeJNtXRoJLt/c0LkLgl8wJHsuBjD/31d+MVe2Y7cYZLZgCh/IewMMEFyoN9Vlvp/h/af
PfyKGfmYhHOgDtoJi9PGb/AXGxEcuPShBU1be9QRjiXd4p5qFiYgxl879hW7ON07Olnv7lHEsYNp
1bn0gke0scHFXYK0kdoQ/Dx3AkOL+CBIXsrcCIw3j9lZ61dzXUddl3WAvMYX8CT9tKAAqepZ3FFr
JhKvT+LheTUO4XB3UXsaVV2WybUKeTgFhgB6/4pwHlROpcwsSHvLEDHG+jGzU9syTaN8/OWJbZV2
SoIoIUJ+1Z0e10rCSXKQWklaIUXvnCO63haEOGin0YyI6oD3VEJezNTfHt9bFbSBMkQUIckM3QmE
nYZf5IJr9aU8D1ORp8fQO4WfUuiXtdxF7L/Y1DvNeLkbnYmpg5yTlAn8PmuzZoD3c5TEVR6QZbax
1vnZruy7QibeEahV87drElG3EpqICpDlE5o9IsCeyDHJ8gWVPPnGoNFEwYeXVCKXnB+V3BSKpD2/
Wf8hvkkFdH7qMIx7c4+mIjmpirrrDkY3zKXNbodja7H1BZ09m7Te/9EbQ0rgr4lU6DoNK/KXF+3o
Xurj7X3IL79OqW90/AJjS4o3UvN14Kn20X83Z9f5/8q2KCEtkXSHNXGUeb2+I9+tO5cScJWkDauW
DRscu/hJNRMSF4FcQqQy4wV16AwqndDEZO2GlphUWls3n+1CAYx84o94rkaoshWCReHxkS/dwUs1
+oZ9XuwI/x1HmKFPEe9lQTzmZT2TsHPwSI2DPkhzcVNtHym2YmeCRra2dmW6szoghNiCr6cmVwCL
SORJEg4xLBwk+by55WdYrdBuolX1EIkwN7QfB9vAs6r/qi4zHmP2tT/fYhiB/+9hr7a4cv/vl1U4
HVnjRwW85DzLjP8HepEEgONnDj50r2YuIo9FeP7Mf5VsOFnuEzqOP2Z/pDOAUUNd8tQ1tXxnihai
4gAEXBAb2Y5uDY25WScBOWuZmTJrcFALgJYYCesnsAbLNCkbBG0YqigIPflWgzvtPUyAouLr4m5/
nG7afaHiFOMqJgnWzstz3IyLWDH1LlrYJtrt1vtksI8c+nPNHvhzj+MWJAbuQLIXIrqPOn4DEXLS
QjkAgrKf/B76gRbzFf4lRjyurIh+UrAisgL7HaZ8rEuHXt7u05htZMDzcyXAsJfaj58V6rMvxoL4
VN7aBUd3dlP3p5t4Hjk31IRI5LOhHM1pP8phmJ1oZNoEdVr3wxJ20mBx9Mvfhu6YttjS2/2NIX4T
+VCgtNFYCuh0kidu0gnffgoFiaeY7NGPrXDSVS93l3VEmYmFLwjhXB7xBxW5Qp9nfUuYL4XEAe4A
sy3Oj5i8gBfYzxpiivw9Lj68DisHPfLQK0rmie9qkPin0rjluvF9345G4a8sFykqtWe1c7Mu3joL
6If8pibAlwTae9FCM2dmWGXRG6s4cslQ01T3Bk09JecbMFVnMbE2f9dDCmqKORvTdBajpK5YT021
FXsIl+lO7vNzF8CedtVNoeeruzZys22BoZ/ccXlkikEaHpbYJFHXqayo3W79MZ7MSpKbrUYCdmwW
1D3ajbEc0m5TNRIHaUlL9XeDLmIxu0Vb65/E+lCYd3loXewWlYovIKc57jcW0QwQRKqIkhyV9xlp
2YGFQhj40cs3vN5r9ofm9wclHXZHlZLSjm1edkCWL8fSLJQaAXwzCY+scKjL4sORrHIYBMosbIqT
dwMKuNIT+FXz6c7MgCe93YpmiMGU1o8aK6UuNKVKFXXm5d65kuOXqKrLv8qUgKWl4Pcx0nFPzINt
IH562AeXXvg3IyIgXhZ1K4Hh5z1q/nAOpJfhH5aRMvS8lh/G0LfLOLwWjIT/9acmCbLTu4F4IbAE
pK/YAbBbbImghN2Md8wN3azfiR8ye8XNkDyGmQHuuML21kPBTW7XzUn/6pVtsX0ZRZ7Bhxjx+f63
2oyOBrr4iQ8/zW1QbguyPrbhtN2LAVoOibZbunxt14Hf6L+jrArNTiYRjrHqufh1/EbK+dulBi0d
AGyXDPzL3jbhc1ys6+LRInAqAWWXGadK8RjJLGfPwxD3QT5qQPAsewa/9FkzuoEzC0EiCFIX+7HU
htl/iDDjnpYgtaFpN17Lw+lJod/csMAiZY3aaLzvgHctFtZgYg6vssQB5ylH7YfkJjb7GmvTEweU
x0NO23F4wkDk1jtcLlg+nRT4HrQqk15VI3OXuJlR7m/YdTZUNS6zYv0rHCnwDVBkhQN+/2paVnoE
Jor9SlWT54p04dwhBoMQeTArp4AAPBbCRtVrqWSNM79BXCFizbVCjy79Y//+My0m0mtpsmHS78sk
eHdgZ20sEi2iYb3QduEURJLcjM65KBvMNmhrKPc9IBG+2Op4eyfSxA/ErjK7XVrq+0RD0vPR/VUz
z0F2cNFQ3OEcHRjopvXSSfp4A8LCphf8T5VO356TRlUWqcFQLkBrpr7l6HPqWehZkhE0Zx9eIlzJ
IquE/gd//wT75l2Q5lwQbNoWSckfhMvs3J9qGzTUUjKQa3ZoS3p/SasPLL4CIjO3KgG9XaUJh1B/
aTAu5YanyabI2XcC3+GYuRhoXHPPUzRiTkRQnkPOwr5UnocbmWfj0EM9rfg7mE0Jpp+3krIDvZ8F
dApHctpU7lJJRc4GsmdgR9LRAfPEneykx9qHyM7rkUkbCr/kOhJPfS2zDuVQ10XAa2BoEGcFIJEg
l8yDcziF9EHEsnJ9OrOOofydcNkXY+GxptShbkHovJwrVXmMGh41GmHBUoQ1tItNfPf+LjSVgHMH
xU8OFf9/vTuQctrNWW8SqCFLqIqmpx1Km5I/TQh9olhSbdz7sQK/9SVJ67eb/GcKAmlUF2mhcT1f
yAoIZGVEtU1sjcnNhpTguwS+mzdMovz0koLImwjwDtYPb6tbr+3q35+qTYlawFeSDJA7SeazvYCL
NGWeP0EEk5pzW62wvKLi97LKmpNdunW/KZ3e4JFF1euJ+AkvyYYFXpC6E/GxP+T2oFjjOoC8Fg00
/8ZuTou7pBAisyYWoXnSJE0bUuQAwVYFTrYBn8EEX1AEvTFbPhim4LSmJ039e77MdP8MoxZBnxt3
6Be2OIFc41iHClzvpnpvBkmCoBn/gteYw9mSe5EggksFZItUjqSYoVczkQebGLFbFMG4tLQZRJ/i
rworHyMCtyIzqGt3Cm/hK1Ylcd69NINnD5sUBgYjU3PcJgL389nAhdQXizhYhWzFnEDWw59MLNls
eLxVyygDXrFtNOxXn81dCbl3uKy7kN1i9aauPwur8EYF+IvT4eaRAIvAuKDc7fqeuE1nsv9CiB4T
ox0mFH6Fq2wjYkMln9s0coCLzF9U9XL4ExozafE+Pl0Jra+0rXxKjg+7QkrlR/OsBt65eonfcPJo
UTVBqxBnh7pFtL22GRuzmjvLKFpOB+U3++LNxw+CAL7ZaXbKfjsa+AmhXGKcZPuVYxIArTRs7J6O
ZDrbDLgf3sc0z5t4VL3mb1PLxGrhMEJpMmLYH4y6qSQHjD0Wzn5n4XY5N1r10WeLR/RHX61jgiZx
iOvmMcwzUerpR8W3ahkMEDh24qfD25/7ss9qn7SygMIC2q6rBqtBhDYszHv6YropFmWD5KYFi7nh
v0kgOxBjLFxSUYDBhZkVH3sF7cnJXfVhzn6E/EelN7ShMK/bwWhR82zU1SHP4+c+7q5gjcGCkoH3
3eItac199jOSEjaYA4yUfwvr6EDiJa8M4GiX+1Ap+T4kVm+b96sJD50FTfydXnupP7IaqghcA8Pt
Ebt+fXB7JB9X/T+oBn6A1u4x+7T+QCokKrooIC5YzRuDFqOe6WBXF4l7itL8tDaLgCAzcCm4N17a
yujaUiQ1k7osqTdQPJT+EKjg7D1qtJmk5HSXE8bnqYwZp5XczTzy+FD1AX+0/NNZ5SoaLolTNe97
DTZ+Uys0dq6zbCgezliPo6ugm/EhhU0F8N5iID125PJVJnoDPcdPbz1pDC+7/nrl3X9Dq3sE4+eP
Iuu95nZL49nZ6B7SvVQ7cwxlYGuv+S3uph44ehAX9Hww+AkNXdkwtpGS7wXeBZ/R9HbqG5cWplNX
Hc3jF+VXK9P5TG34OYS+6mkEXjAywcc2sQX//E72Dzhhza4qhRWmZTWY5ixyfoKIjhL3eVNr8LEa
KFQYX8VSuV45w5IuxLFeu5TeXevIVFIytGLgE7z3oKq/JIJY3TkzaY1ueHxJtsrK58hvbgNaCiPa
7keYnkn3gRAJqrDqRTXK+w+WoLlgKgX+65JW+dxSQJqHfnRutAxVGrQoiF+J4nEH0CF/wFXFBvvx
t/R8he42cgYKRdRqfI+4qNLZRLu9Ypkw1wBksSuC+1yKavGkrPxEqS89nyu0HHjuOW1kyduJkRmd
gJmsc7GtVkCv5rjKXypugZFb+n/SCT/qol4Jknh47JO1QVp33XIFpr2wI+cweqCU7L/w/NKlClpz
cnvi04DukduCzK8zM2PhF+sN17Xlra/O2qwYA6IvBuEucm1yVi2RrfoYETxiyNzAyB/M+EpowpOX
LpFaohi2wHzJEQd4fKNn/Vjt719WXZIGPkBiNN67Jr6+iq/j94+/c080hUZqoTNmPguuUoiGaEmk
P7C5Q1UuUtSQhO0boB7TCG69ikGZcJ+WPcf8rVGRVsbHC52PHWgyWeA4xoey7lAmaJYJGKLgJzEB
TIGslWdhu2iT83/Yd6bSlusj8Om1z5xTxVJ4h1bVPabM7PtGk+SpostCKrjWz0gRh7ydnhX6XM+H
nhICTHGxXno4E/+2oidQeyBdu3Mba43527MvC7XwZpNtUQHQTn6X0/U31Km650chrYnFteV9fBqo
rn66VXSPpZNPnzyKAFGU/w5RsXb8nCzLd3lDnbIqVQxfdffoFLnJ6UCTRZTDZ1r/rwIt2UAxMtnQ
Y5KH/d/STcGUvfT3Fyk74R3qP7vpSx4WPYF1/MPXuPIEWYh7uYIHOdR4ofzfQi3wMLFnxu6FT9gG
X5ibXBG5T9En9MZTw2rd2jDsThFqY1fXa/+JLFaqFZs68flq79HNO4KbL1WYxSkMSgYgnGUUChpz
z00tJDJcFClHshp88Aet581jr5a5IsO5CETNxyxBv4VevwQTVnpYqkGgFn3v+q3hnas+Y9aCNy4L
SE2vnfdnrBDxELe94dJ97wqsrXPUOAaFTzj2rUPsVz0Z5SEX8wXmWe/rrEmRNttGGmLHZe8QHajt
aRhhfAA1xSKwiaLiyTxg0h2ubJO5P8ZOXu3IuihUq9J3PM25Pyn/7nvx7k1YFXyK4pbInJfUsa21
BY7ZITgFmiVkZljg32HYdSh2nL6hsYpHszWnJRZjuWl3qqxXGbBLDXIpV3l1iCtR5D/Wtm84NLCz
sszfZ1/HhonBHcoBg1PQTA7fSiPYan/rzuGxdnMnsFPmGi7I5MMB9G2AZ0DioR/UqipHR8VQS4hM
x5fprrJlHy0biXZs3rWlQAz6mmJ7HWuyKE6nxMvmfRUfMSs046dhev5eenPLGLyCvsSZfaA88sk5
6ARqvHkV9hTEM0XTTLkNRV8k8nrMYTNKJS5Z09vSMp1SDpYynXtHUkjC52OIhkasauB4daR4A0Am
fgMmtfoMHJAOsVcWGLy6EN6wQgV2JCnjOSCPYffFPCU9e+OrjrgIL54czdFrYlbyW/UGzcwuxtCR
73v0nKBoxbPHoVKAv23NPA0ZGuSBc6HAQs1SYVaoaKn/v1tSh3gtu4Q+vCQxwZmLOyHLlfRaYVY2
3JtSq2PnExn/qUMcShIYBBNUKJ0ovjaZVfupxWQU95LgmRFUm4ckFYE1J9fjzwGE/ExG7fF5h8s8
BMQlb7olx5Nw3Lg6b4sKBZoZCxrjY2C/JJDPfcPn0ZzVK+GobNxVAD8pUlbk8oa/eaxtcYdTltcQ
QVZ28cimyOzoCR5OoBZ/hvQjZa8ldoCmdClCf7WtiZzgzw/6Lp6OPaPE3mXA4kX+dR1X3LTW5PNe
BvhXIVEj9O74JMCDb8CGHAHMlUw7LFBRSfNefLBpl6wH5L67NDojiZfaQPdxLLEJAo+N11FViwVQ
Y2LPJZavthzl9/ieZ7FHBTAlSckUI2P61CHIH/qJj7eOGOEu03bkc8LtMtbfjLHCZxazTFLQi+/8
5LfD6+VCc+PZ6hBYNpgGWyGU2QZoE90ZfE02Z1/xej9VDl2mMhwHDEX3V46E1FfU2FgAjZuRYNmB
9NXRoLo1q4uAw4V7yx1vAwxX3ASFfu8kGOdf1qKmtTkMadnw8GXT2eBXAJOq0SypmfMZgfrEMYXb
AUeLDfhfYlwcvIrElZHRWSO9qnc7XUc85WDunFtIQkLT3NqtVgnXIMoa+YQPRa3+7WB8Fb2Y7Ion
ynS3Hn+oTbmg5/5gt8ETRrx4dGWk5IYqRbCNufZpV9NUrlewM1QDhUR/5xi+ddr/umq2gOddtN8M
viD13VVDwBI2u9TtDF3ktxG+El4I5Ro7drw1+eQrvMWh2pudPBWoI5CWfi+TG10FIoMcvVjBPdrV
45WYcGXAOKxI6WUwVle4kHSYwT5O8wwoQCNtEIN24Sw0AflKKJceocATKoxkIVlGbfruEKYou2BY
mPCYA1CwDXjPZOyqUnWQ+aVS/eDf6SH/hxJlIn6SqyrClN7AaAWYBeKd4v9Yv/D1fKBZmBBw8372
JtAHmwGsegE0OcMBSwv3uh22oL9V9eKApzQK82Os+EBwuV7/KC1R+jcCijlznCRQRwxQPUVLSm9W
wal8v2bskGHJ2ffRursc4u+IExPUIDGLEw4NzhaYhzucxjk8sjtvZ9Zv8zgahHdRykRsGGHlnjgs
X6/vsvi7lPrWB4v98M5w5K/8ZlCuq3Igi3QxRW9va9UDMJa8o64vUuGxOl7fGypPNwMOCB1upSSI
u7GXyjglLwZ+3e9wlkJnG8o2WOgLEHCjdP1z1cEMWEvN/yOBktH14u4gWpDS6rkbfGd+3P3tz5FR
0iBGP/8xkXIMtcBcuXfLuGqY3pHq7eSFnBAuo+y7BF6PBTMtOmCJN/o0PApWtmpq1g34SSsVQ7W0
c0BuOhXnL0HYsfgWC9BZQ5ijXH9Bw/6z8FwOQgzEH9SWJfpokW4ExGooSSVxjxPAu3GOQb3fwATn
qgdjoAXDdLBMYP2JwYk7BHxUX/lm/a6opG0FysdCRi8bpe1IZSFtF5W9nmRqz9V7qs9Bix1lQJYz
7s4Mt3DTL3SS72U3bXSG3zxDXzwX5M4pbGp29YBJHzoT9V3NPBCbnZJVdCw1FW+VoCQitS92UNqk
LjdeVivE/CxvPUraNlCqdAIDeYh6RypY+eUl1L7b86nh+5eRWWvIgnUlAkdAcEvrdRXZOpenYue9
G9jr2+kG+e6o4bEb5kIWLAYRsVmqo5+DWYTDvx5y5FohcwW5Ppb26aUeGfRJ8cyUmkpfIG4MnK71
18yaVLBg8ijJ4QKlkpd0qYF7qbpynT1wBq+ZdUXRJoQK4vjohBrmECJBBQ87UbY0+65Yg+Gyjjy6
C2+FosLKn4ZV6gv6wQu9JRjj5usPq4F0RK6LqUKZdNkriBQYojI9PBwp2wxnoF0W3YXTtHt8w8lc
GDm3+sQB6933zdt1YM/CpMBXPwvwyK6Tub5jbk+tqsLGcOiqUC+UrAg/ZqpuplYfmAPWegj8P7tM
qKqjqvH1TMP7dj3zfpot/8QjUrBfbEJPkxtim1CRZVUstWih6V48hE6rFBn7YGBVHhKLWj8Rl7mN
HNcA1OZ0s3h2EUWmU9lRdNWfj4j0wtAvBVzbz7rXMn+z6SaywJwRQ8BfiJpNHF5LV7EH2+zMHYi+
mu5Bumelh/tcebNzgw1Jt8zgnexPEAJNh9HNaTSi1TnBEVAb/pDXD5WFbnZXCTNl9M5jdI+lhS1G
fKwEuTLADCASk3aefWIolzcwo7INXoZbHgX3IvD/v3QV1z2RHDBZLmvmTyYFP/Omp5fhzQzhSTeh
Jsama5fOECOCS9qr75+5B2olXiaOunSOomFqRTu4UBXcRBxRfgasCGwnw+IXKgecconS1m+MhNje
cjhgHdOwjLlbjIdvha4l3C7HvvzHfSNVt81xozQFXXwZjuiXTmrBIoicnY3h5yd/eZNnzO5c5cQd
y7IDnSGWNrdh6dVufgngQgM5rMYsRGp8peOfqy3RgXDF4C+XcyuaW41yeUHnHcJR0+EfTPhLV4Cg
pIR6LoDKtH+MQ3ja5V3DenZJDT4Enaytjig7ReAW8eh6+PQWKj7+MlU7grIn6kHdmR1KAKLUwL/q
uH+vD88WQc3x7p8BOJgjolzdgcPF5anPITGz/jH47MBTD/ke1T+3r7jHLarJezFe3otGpqZIU3lH
JykupO+Bf9T6KpOqvR328VqZeHDuruiLZSonBh30dYGbLU9lSx6S/cG4+gLAbxaIy1gRiXWbCrpv
VVyn3Em8SP6S187kOkPJA1d+2pbmoOAQBtPDf3VKeTX4Ww2w1lzmFRPgkSuWSu/1qgMmdC+qjUxI
OqCNUr7sIIsanMcc0S1HDY6L7zI3rKCgJkN9Sn2jfRA4zOYaInVW0tzQDw5lQph8ClieeUq4DTp/
BNh/HHbwXKxvg0koNS74z06FCWyXc0Z0ef8683Kue+tuDOA62bOiHvWAqNFLsIYvK7LWKbfh5dLN
wTKx5AB9jmqFxwHwDDQhjHqYA+pID6f7CAFjF804PocNjUQmzCsK1FWa1oWOcwebMOIEfTEaG2Ke
BRblkUgtBRANnHA2tb+TY97K8WvqFCApSm5LZNt2miF5LKO4Vsza8wQ01Sj3hFmhjcPuNp8YTe8v
5F2QM8tc/pfK8xuyTECaGo4Fsz1ML1uPSWI4Mk+eYBRP0lnfye65pMUhB/9B3F3WmEoY4EEW9T6d
aEHcf+opd/4uiab5Gej3ZPiSstXohHvF8SYBBWKOKReyFeM/45IsdfDP94bS9qop2vlnvwfyu/HL
WUUCSMwWbqXsq7zAAKkbDDOvqxuldZpcrukk8XDaNo+JGN6mxPAeFcuoR2iPb/yeC2o5mlc9aDVh
WfXAOE84OOHGrigVUc7A5EF2df0lqv3QgHQycK6gZaLppUhh9cWwethSCAUjGudOyovOD+dhIyiI
eRKW27ZZA8KJAekr5AmX9upx01fnWBKwFs2F5NjqwGtpyiHJwiy7OtiYE/ai6eVE8KoNofCaMreW
cLNeb4BhDgyBxLpTPulhyDLWeJUK+fg5/i9xtgquvwwsSnOZjIZurwCZP76G49s0USBpK23snuMt
ecPFR26PWrGiGJTXiUdovauph607eQrSPoezaDqBNVyZn7UHDICYDPvoWs75uxMdqk4uXl8AavdP
/4gQvJVcE1aUHuH/sIJ8axRfSrcHf411cLT2O6FTUVDNmondK32ePZl2r5OhrUGBG4cQ23ut3Jfm
qAWGT4qs5/rmSzChcq68haNYIGMtPrIwJu0G6V5Vg3tiZD6xYJoXL7R/ZHeZQs/LHarct8A0VjZv
yztJP0yy1q3lIbZvA4txBprsTpj0BjLQckTNUSvSFqAHpJ+rmOaejZqcavO6C+0BZjIgalgDDvm0
wrOGjg12L/1NEEf6CMPyODIl10KhZGFbWu75bAKdXPJU/YoM4KUNk4S0f/UXW06JiFZhe6e6u/ks
dRDrenw/I6K5XVa9eSoY8TssvXEFsb0Ione8aC9yQk9XaOmnJ/azImj8H6O819Z2y3VzLLAvRM5V
5Xu6gqPvD5JXgTj4+NrIFBp35BnKJMxHGVtfETg8N7D+sIU6EALllJ7+zvQl0+MS/PSq4yZcK1d6
SeaiNXW70Cu4BMjeM6RrxsPJZdN5dXbDd8ISl1lUbznQ+yu1XFjl9bxfPJ4kIwyI0OThQVxkWDd4
pb5zHPjjbS3aMVXe7/yIPrH7ZcG7ptqwW0Kjo+9De0UNh5qP6PjKOw/ojT6CSdXnchUeUjKVubod
UBncc5WxbquLpdHFfB1/UE/qW9LOSk01Oz6VqpFmp2AejphUi5Ih2mWkq8OtKAJmX270lCR2HtW/
4LDOiD3OvPaLhS3eYlkEmvc+7WAbR4tEQOUyr6mBy4McddPDrL5FNTDTxuCUNamyxGjmv0AzYYVO
qpkytAaMTl6v8RbYZAJmeatMgIlmY9b8+TYsFOGwulMnCyVFZ+cW9LSfZ4AWV8zFkdJFwZyigBm8
dpVq+mctr+A3kBDucoCCX800u71me1QEA9qG8ObRj9+mOfwevKwtCJofTdER42P6+5LZMudf7nbd
bbQwCKGFhJnK8QWvM6X3ZxfslZlUq9a5sVGwWvUdREpRMDjl4Sma+1E8z08EyVjE/KQ2nQpcgHoq
o3zJr9V+4ZLpIOCIdEtxi4eMHWtdSkntFNYkzr2h6VrGf9vsTVr6/D1IRcvbJuqdpPWojfQlcVGf
lUWA6Rik6Q5a/gQdnoQI+mMlrQfmdxTIrFB+pJvIufJCWFA82d4DGwcb96gTgckK+zlDlAo5Sk9G
AptBDK2UkOQo/GcSaPzRhKEcWgUfXUxhKo/0sHRDFwgCKKBmZGqPQ9WPpxXFB8apWiIYlte9GLJz
AzmA2Ud2Ds89sDHi3EWKS9XU+Fy3NeSnryEW+TO+XfV64c4vb8KCYefPTFPIl/4R3qSsB7XUEJXC
/x5YTUIoBY9eCzXRfo2PUKVAa+aAjqQQtyg5WOUaDQ2r/ZZSSh1NRZXwMp+fUL6ijNbHZrfmn/LR
sHl19HT7q0r7JReyCDSXBNuLv5tZeYSxqsuzt2x85OuQePCjC6yCZ7PIdfRusN778TPIA6U1Jpd2
aEwTkls7tOEiI9EUT7qUv8RYI3zK7qgnvPSAk2D6WXC6IJk4tEG8JTlp6yQa2azbtSButXqRPE+V
YAE8U2GBaXrmkJk3JquFAgjbmeAwcuH00dOsUO+vbwvwX4VVhsMgv6wiN8pW1IY4luefz0+tQXVK
D8qASzetsZEsTlwvR3RlJEXr5gpTLqVgGtAR2CK+fePtf/zFaS2278pEOnQvLz3R2nc0/l6kZYln
f3A8aCGvg2VqpYiybN5OTuFeBIf/FoHGG/tIvIDb2Qs+FgKM6S+6c7qf/eKGJqrYZPHOXX6Y+zbe
4RDR8XLGyJZ7gtXujckqB/Bwa/rpST/wrTqm6UiKrVSKP2YvFNw3wOYHcRynfzGoubtdL/GNFYal
CLnIVt0DlJIllvhEBfj9CQeFnJP8R7huBwF/YSgxzJtKP8E0BXVWi7rbWVTdWP+MAebfXhohP6KO
+9dFrdk6vFijOJvn81z1dxpGAf+GncGbGsV4DpcL6vSJNwMZVjJwB4yMDGVpd3/dDrbsaz3muzPS
8RYV64wJbEsrKteylQRngpr+5LmNZ7j5B5fIEPSpE20MjZMux4Iszb/DBp1kGEgGwN7iQER3olrN
hmPhuifWhli9mmz825BbMEGNJJPIAuWDq5cJ74ZCoHieQoa516EvBjD0HLLAZXbyjj7HoL5TZ8UC
53vOi9GapTD8rslShErFquC07/cqzNqm4wJTZ3qe1bTQmePWxIvJjoqXEkLYZSIeEbcfQTDyAz7v
NkBpPQgpBak5so3EZGW2wQlq50TY5z/NtRgQurBs8skdzXOFXClq++5CkGYjMOzJlzXu7rRSiud8
MHOErkUp0hdB+4HSvm64WXkLZ3GHP8E+i8DLlrM/FKlKl9np1JqkClwnJpzf0BQXezpZb21/MtMs
mdGalkjBhLERjztdZtiWkV8OTrKbaQwr0pkVPhV2hcLHje9PSsPc31UlwbKisG205aUBk6yAJpIN
TOon60X0pLd9dlGFQ6ixLTfdUyhS93kqN14LcegeDTfF9WVdKeSZBzjwPzeyJXui57B4vKVmIU59
qZdhttP5vCZr45hnlK14mNhK/NTbkqXGCdvFpm8TTZy8C2r9udtP9VRd+dTrg/xgSyrPKMlkvqxd
S+HbyuX4hb4DbzoEmGXSCysp15BajfqqOXsC2tgtqzXQiiabVN/6DMXdJ4Ng4q5S896/u4kJxTsl
KRGewxw+XPiFJNnUIUpU+3Z/2/hwbxRWYtcxO7QAbw0U6ueH+K+1PlzscFI51r753t4mMOIeiCaX
RsSyHuCd9SS3OGp6pJE8CURyZKryHGiAag1VOIMhQbxBpPYO+8hko3HKajXBtzcp7ImgIZMfLeWX
6s2ySHEdAwu0KbhycMchK9GD31wMnU0bwMqvxPA79BBK6qO+PoBm4I3yfqks4ag5nYW5NQWz+9t3
JdwUjeW01lEYmTYoAQ+LEJXMhVSnajsyRopHiExB2tKRJIEKRv9BTTbq0E45JzO1KLtuDdZmCjjs
NkRPGPPhHyH8E1ZtYV3EDgAGNa7wezGTNaUqkBJPvI2LZya7eW+SXs5LpOt+623zSIUcwwHh743w
sAkkMEJjf1O8uxsNMsH+w+9h1jvyDOmFjv2pbsOplvOMh2NhuP3r4evpLWMBb9WrSPkUOG+jpk26
KzDOJW2/H9DTAN4Rimm3ZR64JOirS90bDzJAdnqwGQmgkyEiKZQjw3RcRJME491uIXMCnyXwImGb
3FaqlwitMrCVZLz8OXZXxWD01C7eyHpDpsGVgWajRRJj90G+wmMqLFWQ2GY9rmAV7I7h+W2NHnz5
wVUWJ+xT72fVmK6pkWqgRF2UrPPTOAWjiTE1A3VwbAoSYJ+ny3ZyWr3e4cewu4CPPD72cGOkvjjr
v4maMo7Qcw/R1fWC+zG599HSWeltztj87MWV7QhbRZJhrxX/3XWTehbq1YaUgT0fKO/N3/RPh5Yh
XBUZGok0bisadvsY2uS/BFst/n2z9FKkYdb9zMTS0n4+KZa28hPCav4HR/0QM+zRnCp+hGsiEMbQ
xBztwk6bzhpmffZPzLHTIzZmeNsgz5PZB7GZv8jDoDSLmVDL/W9rZauxuVM69EfNtNFVTDaTIwAQ
9/FU1MxmD+E4zcNOQcRieCulu3YYiWo2Xs2eC7dDTwQAgF5J/yAt/VetCnmlVLEZVdHzDDpdgdbW
hZTikkUBbFC+TE8VZ8xtJLtXhfGuSjTC0/OPN619PraQ+HBsNwxmPBKbxhg35Uxv326oIX6DjsGP
+0msrLvMV79rvR9tpQhUvAKFxzUDfCYMmMCplGmMtvCv282N+eKlwThSvyFej4gJcsoQ9VQAA4Hs
7xrBFPo/X7dYjbRF0CvkHDUyk1KSSCFLfbpnZQczvV3QdwnfBRJOEgB8wG+bfiDNAZj6sifBFAV+
oMhPkgS1OtLTt6/LeL4ap0j5e8yZ+nz+1Suxaxzws1XPwpsdgzPf6Ou6o4KIteOE2Z9dhE6BiJP7
BdaQbjF5z0jPFcliCO7BYGaFUZlHK6gTv3X+qfN2UWBW5NzfqiQYukQQJTL3MytHMJzEZUHSUkUd
Uwt7zH8MEmG4SoUfgpcNmz4EH0OhUwgPAhpW0s+JrN3RZoTgPGjZzyjr1HG8MX/fDlBhNlPru32o
vOoVhLJaRLdKdgarhWnpWZwcq7CYUeVv6puaSFrBX4PwBJ/JrjZtGvSNdx21hY2TjJjbEt7/r8Bn
TVWMiA+hwAPrhKf1P3x2ySlnk0K87q0kxsYHhZvISaCUmBQMCgA1RNd+rzrc4RiUtwhqSDNJhuTX
/ZK2NfBLvQfv8fT4PU+7dVhKvfBItO8GfctFyHFIPilkM8xYcr5HaIACBNLxJevSKGmNAqOTvFp6
AKo9hoxhCUY+Rw/eJkWfOQa2CQ/zhYc/cl0dk03OkWCyXCFTy3XuNpgeOFYo1nMV1eCjEL219JBP
DMh+DxB4FlkR8D7mNkeecQuF92hL0N4K40KVoOUIXfNen+rP52HoUyjSTn4WUcQ7HW2yEQ2KmVel
JD+K4IxdUdh+jF06vwAh53v38eNx80w5vbj/Vcw/P642Y+dTkk9rwBDDcWTiB+EKinLnWiRCbvNh
lqp3NyL+YWbp8ho3rv7RI9EweEQX0C948VbqnFTlE4uFHJ3K94MXn3Bfls0qBt5z9uwseZm8FeNj
eB3Dq5HvjWcGpm4bBQoVCiUFUOTmgfSTr3z46LbdgeJkTV5DoOVciQEWL6Ns3AZuV+mhc7i6meBl
mxkgZHmlywomRtW87+MoIIS6JVu2YvYu+7QH2e62AXtRsOyxvrPhnfghSgqYqTS58UNDcQiIIBc+
FT4x05Mzto6vci2gX2ZxhGNwLq0CzGeXABNYa8WQGCdnaNWdPfASIyAX6OSxRrkqkcyIXMEfkW2O
ZHcjHuhpZ2/x7ml5Mv6PfEo79CtuQ2voZqCKZbHInogG3K2BsS5f3oF2+19xWolvP0a1hUsaBHhB
ff8JsKDSOvkHGgfMUkUXbnrrgh43KPNVsCiBi0kOHJF7akFCn2GHSX3uFcljy8EOcGREkbYbBYvH
SbPTY3xMGA8oteDXwbPh/D6j8sCR8LpqWzDPhFwVgM194LESLHmXZaTFSbLhhTMgabUZYj92f7dq
1WHbEyuegxQEB80wac7tkD8q0SkSC7irVQ2a/C0V5I+nruA13v3JjYqkcuvCHkJI+Ro2WQbUud7M
f5b7z54S5FaXenq1+rPWYXOO3W4MPDAz4R5gZ7XO73pMomztuTc/XGJmZnoEsAUPmYJ8+7XJndLt
7IhoeJE/PLs0wyWTXv6LoFO/3xNE8kxD4yJc0jtz0QNzO4rZc7kcWpytCa0IhQwLBHdGZtBNhzsy
BZddeTiCUjq4VGn2wSKcFMfoxQJU24jPhFStdArarfObn/cfHHW2MDsAtZlH/+sEy4qEOn32ZWKS
NfhtMqN9EmjukuN/sZ5Gpy2GFPCbVm2thHrMrgqxXDCXQu5Qb/yRtcJZSN3LbKg9IoNmNT5Ho19O
uj0tEhZJhX/j50DmnkBEa7R53IeBdqAHSOlYJy27dXS6NeqIRUJBDM6uuB0TwYm2VNli0J+VyQ/o
3PJmcJUlUhwi/n9Tg5OTZT6sK1skloEuyllVMiTOMGwykvKWZ0pq3EGXEQPWkK4PM30IqA79QT9h
VrmJveV4u0cqHDivl0I3WiTnwKOrt/dL4euc1NUF9D99UURulE1mwt+IO1O+S0kXwOQn2KR5svAP
cygdjH3odCQaolJvPf/+12HD/RbwX4STenUNyaO+DC1QJeZx26Dt4yzHPyRlwS4vhar1aoUrm5b+
lkAMuBQIHeSV81u1fdsLwZMSkLsIRNSrH5ow+EvgCly+igg8Ej76wtRbYFSudEV7qcWoElK9ZlIB
gMuQw/yEz8sZ4FJGlynkM8Zoq22j6r+mk4bXf0zeHhxTgt/4ePuyqjRIE04ir8ak0RdY57HmARFa
2LdmnmrR78lFhDzyeGZ3SOWNcZ5L4MHQJzy9BdNSAx8gwrmZAINCptnp8g0bMJ2Mi6lUhux3ThJr
fJcSOxL0j8HSFP+Q0hjnSoAg/6PyO9TESj1Z0CM/jsqndcGVNJ1NB5T2/G5Nr0iwLGdhiJdACNWD
434Hx2V5qBDsWsRQ6dUEX4GiWotRazFnH/eHVAi6MXS4NS17fyGOeKpdj3/+yKw6wqQp+zTrSGxT
thywQHBH1+tV9PitbnhQb7U4JVPO7rKXX8VxXg2nbe+puR+oRWroyzdHzXhcgw2za6Pqd0nl4l/C
LOVrQ3wpS8GpCJgyCmXZvBg9KLiEWQuSxh8dt3MW1amODW+6dhCk0UaclOkPI9IokMBm2Jvg+4i4
EqP6cajaAQRMhlf8EpBYqI5Kt7FwDyNi8tOiUGzaf52JXLtNtCHc2aTJ9IGxnVlwZd8yK2Ls9eiG
7qXia5hyj4y6u5etbj/UKvXFRHiCmONeMeh/60bn9f2H1oZmXUDpp46DILRpYus2vCa62lSZ4joz
QqjMpwdaLhkRQ37MKi7Oq1uQVoEAwYnRDLSXY1K8nntxWtDY9uMlYYxMsskZhsptwqGSPm62ikHf
UppgTLUS6f9kouNd2zKIsfSgOjBD88fj0Nr2PuJONJmphAVDMZC8XMhZIc6nDWVfdHf1Q4oOMSdf
TpGErEvkNeY3PJzQL19X+unhMHUrYdD/clAQflh3fCYH5DiN4KDWD68T+xOz4+Wl8dUrtxvf7fYZ
hgPLIr7W2qiAP2T3ojB1AHDgPkURfx81A+6wxlk4NOCu5T//9nTivtqijTWLBi2QsoHv+BdmZ5lm
+HxU6sJWg5j7lIivckSLEuzJ1uT8VXc/CSKuRk6EwSIal3CBFiMIAkL/02G9AK4uRkDj/wKMG69c
yB3lVHiEDjCENuzIGvyoy+to9BwkArOl/M9UtRAquDHJLodNeq41er8Zze7Ti2lvWrvKg0Eszwk1
Bi5tvKvWOHOHjX0jydghbR7ZCG390Ivd0RfWJm9axk+aJbL2b+6brbULqACrh/PMxMZDqIF3kCr/
qjNvdBaOTOyPeWBBLJ8O3jQASeHk17KpctJPbJ6ScgT3nnQVmOXmMJEolq7QVvGZC7hFuS+2HXRg
h+XZlqq/meX2f3oUEhQVJOFaE+4c6gnoVBOdAh6thbQKjp3se677jo4xAIrPFDteDhv3HzvvxO6J
wfGGEaqYh2Vq8D6qqyZrngeJxT9gf0V2QUalYl9lhQISiOl5vaZDPAjoYwGAgqaAh3n+yUasRxu3
EdTSkcAhW3EuGRzypwt6fVdtq+HWk8j1cU3OBUA5q+G9Q2GQy6p4/f3YG+G5Ri0DGiIbWTS4DV9a
YW/pE3WVlxsO8rPTHZBaCdcQxMm+QFUpWSNY2ZbnnA0ohfqcKTgMCvRoeBsGHmwD09kehjFsr/94
5m6ZxUMXFTjX7pItYg7JeqkWsPG4sRcEERAWyb0qyVmsITWrhGDu/Zl1f9qwyPH2DyjqMs/+il5B
G3yDQ6usoVstevxu6xqA0dGi9My7OTpmnGBXKg3OXRdF+gDLpkxEBMpO7IkFsIk5k1kRyPMwRG2T
QNIWbKGqFgUhKsyqwMJA0ZfM+SUX/tlDt0gnC7P6k7/cHirWx3D6zVTPvjfePIvTGxUwl2Cl608f
tHvd5m+qNY3CV5oY9KJ1DrKw8GajRTGdmjyDgWEWrgqZ2HEuKVADIN74+2yAJgDecszA15KgmbFs
rzB8Gn+GNsRwdOtWzEUUW15PVPqd0tki63ILcvmUPNKKZsvv6xYCiEqe/ZIVvYF9FeTFMsAduVuR
LeE89uxawRtup2b4WMBZ8lXGhBddJ/Ix5sZ09WE3WlEmnZYDqW8WFzqKDOmQ3G3nlCkF7GtMIi3Z
NJav2suuZfVFKnyqNYWJcqGEBDYp0bNJeunqOGowO7tkzNsghSHI9aWjBk4ZscZmtfdQBiLHh492
WNNaxvnx+ZTBT9/nENGArlXoJFOZ7ubHrcg6gXVjozh+3c2ERo7y6JAM4rzE+t3XBbeTIsBZOL4A
wOKIQBWViklBKfUZMnPVT7dYCMyqKzoF3lodgiCzwROoWZGj2I60PmCbkxoNJKyVOoipS3Tp45j2
b9yuRcixnCwGO16xLd6LBx9tMgRbbXg3OspJqtx6q51vBxpStEp6+uCMaeaGZGI4nf4JQwXTj1N0
leYeM3ZMNULwkzZealzpjszVxPzB7hU2X7V0f8cEAdMZb9QBKyD5lpjfJLcGr9/xjat8VmSj6I48
jBXIZ25Jruro40WcAcl/kHDZv0dtFB4DwNz4y1ruEtnztAgTk3FHTf7AyBCz3R5nXcxZQzgTSeRV
VoxUNH6c5+QrUb1l1Yv/Qs7zDPjQ7rZC0aodDNt9zbfCmlzxVdIytGATDIsR7wTcs2MUqN5wR2Dh
g9FPjJYoR/Z0e3YfEXRHMXhqUA1Qfj6qCq0bVO5KytVejqQlCTvZ9H30DosUHEzwhZ1G/mC/96j0
oFhLKJkiA5k3TcHSnfdmMgJN9nfj306gpzMWjzAaOCuYXDcgoFwnpdaQOKVjUDm+SN5tSoU1l/4o
jDH+FLYkCUNchKDSuMqgK3RXGJh2I4lbax7jd1a87mIR2G0lr+Xf6j1DuQExfhwpoJe8e2clgVod
tXWFndxfoKxV3EYNPqci0QDwnT+8Q86sDA4dweePTl3FMU68c6xF9TAF7+qeu4th5bh/GFQf5vKI
TKF2uM+tsOGMpdnHDyatIK4nQ5UxSjrNmIgeRBoDMh9bSv6oAOKik+BiWl8f6rwYiFipkfynId+M
ncFlruEr5aO95oJboJmN5NMO2XKq6x1NAi70gGDsULNs4BfbDe7jk4B7dPE85WVAYMiQ2UpLqnvz
AFfxiYzlE9ZwkA06BxCy8aIC2Yr4dI0iyjcNLYSD1pJ60f07umfsf5t8zJjjZrc9LfSH/LHh5Dt+
3MWXjRkQ4GhPVZ5Tr4OEtjG2GbMCJ5P2hn5CVTXS+6BKiCi42Bjhq+CiOGIwBTedkt+/qzqrmTE7
LO19nocR2V10f6vIpHqPVPuNElNnCKNPEHv8VfkMkEjWKFQS/xrmZD4NQZMVuRSsMHwUPoIES+l3
7fd1NzQznkPUFcJr3lU/d7ouLIVzO8y6jx2rNSoc2gOmLrzxkHgCx1oiZWKuXecWM6hTQP60VnwH
y13MQ4q7Z4piKSU6o3NqCUExI5N/H2diXwNu/jmFPXs+BfILPKGyAWvEwlymyNvnhi37arxOIWAV
Hxmg+hTS+BzUC2SXr8Rk5+IP+Bk/kSmoIcCHQbKlTAN+50UigkXAgmW9hDXQJcPPFNX3SdZYsc2s
UXNT/uvwtjuMnaoByWsH87ShKcL5R2EutroPFxheBV0boVApu5fto4foJnuxIBcK8DYMbnR3r7dh
Vl6onqCGNQzMF6JORGWXIoJkg9fEiDedCGyvG6UbHMBCL6ElnM9/Tyz1SsIa5lncpzasNyLECiCs
WNr00olAtL0kTMQy+7EBsyIZq0N5p+095dZfQ7XsRyPJxO+cbAQETg+q/6Ic5Y+CIuCTj4KPJp3H
RPWlvOL27RJLWPvmdny7IJcljD2LoasZj2YmsNRteC4FaLApUN38zH5CvFjITVVkuix3c3Ni0ulM
xG5oI5+keBL4DVNpWqQGA9n92f4nRpI2+Hb/PLaIRTx4YZRlhMyfxtgEhkK/7DrFF19jeFEUSHU5
5w+lcXpgb+T0yhItJJJ7tRPkVP0xwa/iP0piEodk0IduhExBGcaaGmQphSyX9XG+KjSR99LRFk+/
KuZy/GOYXmhd+TjwEW+TSBcjPs8p5M7RrKtqdF5lqJW6ui5wRTcUeuJYaeWnbaEJW5eDsbJUrv7g
INcaJeLS3dAZAIiplOURmg+WrdhW6Qw0Bi71xWbJPggGhzP6SlUbDg8FD6BKm/ki5nNuAr2rqZua
Op7RJ+WyKcxNbbWyboWxITQgSaevwri9aLdhmKC56qNhbEle8uvottJjjUpwRzN2EUYLDWL8UIsH
smQHE5K0eWl6Yu7P7UcsIK8CH5RxA9YfLR5yv5wzrE9q7Ablx+RXILjXoXDowVOiSww0yYrIG0bH
gaIneEZPmnaJbmScoQveCnVD7Zm1lH66s/0XNlpWPxKbiGl1ty9AwNjqYRl+Yy3L1BTPEKddOldn
nfHrVfuVtIMoKjyn1AdVjbq9abjU1k39ZigSUuwR0mRGizIco+L2JEkwRrNfZaOfsvFFqMfMqAuE
7Fgq+bSjeHSlgou8P7uZcdkmdvVptMoTs8JB6G6N12XckWLRml6BZdpu0rpxkrtG6FcWGftz9i9E
wL6UJoZ0vVLuvLMer0jjocqfFtS98YUt3gA8ZeacODzozmvkvhkBk14WWp+AP2X/FO4JiV6hMhxa
BgsNdCT11ISGuwOGjP+dR7/lPgxeazXS19CdMwM608I8iZZ2gbkZvzZhemR6CkTludYgP6GYviu+
oUfzwpdeXT+B0bi1eeDK2FprJcz22SKB7JbZzN9+zt9WF21snwFKk9BLyJyoGtJiCPMFIIB0kl8O
ONcT7kXSA98fFyvCNcv09WMfu9QzG5u08P0p3RnvIsZmYz7ZDCYkUX5bgGWq2ocXWXbjcebLiCXj
GYUIZBZEvoB439z66V4YSCL+vi/V40ELlrErNtJLthXUjqch+nDzZx5vcuY2yIy/9qZfpBOKC00u
hL7Pchr7jfuAVZJGXF66xfR+XKyx4qiOuH8HXaryc9nDIRkAb2XRfYMjR1weW82/4YjX2S+8y0DK
XtmUYiPn3m3nLG5EteP2/XkE+SN1UjPHXFaSxcxmn051zy7leYDoIphuK3z7Eiwu+2VZBZn3zaMz
t0GTep8dsFpAvyi+3EXAbPv5H76jHuoxY37Tmqg4aHu/PY05vmVnNr8fbeZNedNYbFDrhK7gbg80
NYnMLGCXu65bXWA2DNDwXfhwA06iCUTxXrBA/xTB52FnoV7mjTdOUUSRta+UTjlUHWimhk0nSKcu
ZtokICqu5q3MM9vVZGBCutVBArLMkgMfi4H4lKKeId69EEp01w+VEOK0Q9h00yK8ep6gdmvSdET3
FT/6VdsorcqOgKJQbr8SDa3lEb/UkZY/dY+3moECyd64ZgYR4Get613IFvSRY9jai8Xo5Yx7IDbI
qzQ68blVtvw4b1T8W5+y5YlcNvXGRFwZLMDogV5OEq/PKfb7HCyMpq/6RdHNvMFtcjGkz3DEh3H/
KeXwwQa1QQgNZh605Z84BpweeY7fFNhcqK/cHwiW8RsAKJ72is6upCPhGGKD0UAYFy+fTuIMD8lq
58SYnSpnPr85tNfmU3mMd//knpqRJh5UrCWBCVxv5YoGBZ/99wZeef/W9sPxMfloGV1ICJTllnnk
f63j1EWcBMWNWXxDaDy9mVRAY60jsrNClzgcL80bQji5//aECwSDBozzJGLd7MCpTvXPdgI/lbSx
VoVg1vos7Fiv8SzpykntmdgvcNktTCSkKXj3t1wlZSfkPS3sa96kjbkGgBQ8g38W+XYv1EsPhnkX
tA1YCozdbRMXjxuF1uckCgwX05UOxZyIJQ8NSGZsw5xtvX4MwJ0WIl8PcFe4TDQ5/E3H0Q6WCyKQ
dVGSaAIkJn8+18Z3j+0tJXBpjNFA6LPO4fTLaEpHNVvZjmxLhF31gMjY/pWppCfvgs2bzIGi4Dvk
E8tObISSMgLZ6k2EcG9831MEeR/Exto6k+luz6RjtUSWnzXAqbrBZmZvpn4TU0ba6xaM54VgWvLM
C8iyAn5KY3Ww/xVHFxdWk5ZzZ9H2PLoGYXyIEuu1wgEv3omu34DndrF5kTABiGJXZL/H4yvqdaSM
F9F9VorHKrTRKtefCFt7B5isJY4fZxBbk02P1XfOAW2Y+TGnkGVc+gE8yxFcxuSCs6fCFUm/+P7V
t98YM9zj4UvP7Qh3UQSuaOxqjjAxx4Yq/biZTRkFuLZHqvwH0XsXdZmb5ryI9wjbLGSgEJW83Q9g
6pAN6yIgK0QAWoMqpnAnr0jPO7XokNhPZCQCAK/BFOMXyc4DzGE+b+nVAAT1hWymf8EeCoxf+0oQ
QEtRVrVuz5XCrMOiVAbHyqutM57n05qLBjKDVL9vc+592oetnHGQEcaoKtGxTvu/phPBPaO4Ote7
0qxMvaYzINur0EGJ/8lOJlFAJUoIcja1Sd1YeJTmVLCYmM53xLcl4Xp5geT/Rbm5fSSlIfQ3ubIp
Y0ouekp25Fm92BoQZZja3+RnojfQD7gUfVOcLPSxxDOIWD/EXo3j9h9uCFbWfRHvfI/flU8Mt2zu
HjZ6wvwAMLUOE1d/QCpB1tX7T50JCepuPnSgmwoulP2My9u2SbAtrKew+9RMtGxdpn24dZ/J+Jie
7e9GJ15WtQmYAfulAyHoXn484a6854nvS9MMbejDV0Stks5p1Uyw/MnIpaxcnOSb03VaXXfvh6Rm
cSvef5Zl6LzaPlNTnM/NFTIQYEyjZqSkr7ri2k3aI8SeAheZW25qXeZEbZQ4iLpPGlDyipVmvnez
UPrdsvjBnA1eF2su4JCN7ILQRLQ86ITc2hbxexh/A+6AZVut7XAdAmT98M5y/JLYvtf/fOj5MVH7
mJM3Y61Bi5wRCiqCuN7DY0E7Z6yB/NJQmUx/tffIN9jQ/vH+GF1oUDb2a+EBFEJsGA3NLETrkW+m
R3pkTm7v09HkhNgmnaTT7eCmrXoq5J3+D0A05x7c4q9p2FeHOKZRdqWs1APfg1cKCFdnmAd4/OdF
UeV/livZuKU9LT2LMtjOzgHv6MxOBnKyt1fVrGVx4uf5/SyUF2YipSWwEM1ssTwwuYJymerVSq0a
a697mKa6u/r/Xk8VgIbPtBD3w2AxcfwzRdFJaSbR9zDemEjaKrxFwVQL8EeNljHZsfP6NAVY2a6X
pFkb6dYtvm5SjtxXTRsN79SKrOpc5Wh1+vSNZH6aoedsos5+c3sG65MPrIc5XAlNY+MwNclZ70wh
ZKU2bj1GTom4TnwteLwhBjQtSGdMXPO9Ae+yI3SuvNkN+HiHOpToXFnjoRviHNGfdsaJOgszYIjp
G7Fu25v4Czjw0y3OIkrBRSgRSWMARp1PiKBaVgFrD9btaxGKfNEwgN1cTo7YxVdPKqNmWkCmSeGH
wwKr1zvtexQQ+XBgu9hQ4MZB6uNd6rdJ51WYBh3Jxu3aDk8bwNHJKq7PFZkFItZ4G71e/xVnT+7K
0tRFO7FIqwoWEjS+GoN4YNh4ohcZiexnTEtZv22y16bi4Z0cAdlGNwpIAQUFzpqGe4PlS+5DTJSH
fXhRlTFi5kgFTDfVFrSexVs/Gh779qLbdVH1AS9hBnVVjAhnWkS0E1vkbHhl3YLg3c8gXGIGmfDh
5wsxMjj4izF/evrdsplNS/q600WC6jiW3+KnGZ8jApZVpyDuo9xeLSmPXNcD0OO+BItlt0Xhnwb8
KitWGkE+ym6CMcTbWQ94b3MBzd+b+8llL8DxYTPDFb2rftxXlBGxrhwC8KvCuLLqLTqid/z0An/p
BSDwdHEq7xBeffedApCcbrTYKHjanTNNJf1om4GWgEIJdcqQk4BHMyUKP9EwLVTXUUwXhJWXwHJ/
vcyXqLl6nrHtwELNcHBJifljjo+8zN/yMuDhkwGRi9PZC8bJ8vJwsmg96sz8sIaoiORAODxhARuT
DztYOONZyZhxwtx0g0X105R4dILn8HsDQcGv3uLXy9OIxfF1oxyCtKpdwZahMJOCuCcRF1AYPZSN
dIwMNReg/jCf50sTWWP2stZ4UDYuS3F+TDOavL/5QmTqsuf4Ekgd1WTgcpMFr36dWgkASQL+Lt4R
di9xukjHrKiODqtC2DZc7CmLeHmqjD88RJ1HkLHD6aFUd+eP6+r3+1SO/RtNlrD/oDJ6+/cC9WD+
7foQR2OnAOmFSVVdi4dzrcvu90vZLmrydkaHOKnQe5WagoCEgg997aQdKe3LiX5L9mNj7jUkkMB3
tpCJyvDMKjmvHFC7kxxgeijpKwBzAmFjF/2RnA0E6kMgcVc9NvRftO7oYhXoK8NBGTbBHjR/Dx7y
kz7qqKESQcYj2YdqNTmY0UyFAE6VP2yBfcPr723/3Nsj4DjcpGpctwJS4I5/tWsWAvu8vyiKdNFQ
SyrsPSvjYPQ8hb12FBlLtlq+9P7p3iPZzjdmGwbRlqCiQXRGgZXz6zt1CjqlYdOk8lIf1wH9X8QC
LVmBKDOOEaeYY4ZuzxNknDwsX0GA4KAUqVPzEwLG7uKiyg8PSeOEMPj76qQCxZQwc3Bws9uhCBXs
d2s6wS26ZwS78sMPk+Zvx2TB7A0J0yhRkUXsTnyDmgR7cJ2TdH6Z8G2QTtz8phaHeMq+AH1fpd9r
j0ssv7bxgy4z7AdQAyJ4Qt7hvAqGnIQWUCW/khIgbbnMh6MxPSMtOSqikLZM/4Z6blEAOdYPmvKP
2O9TEw8kLnQF7EsKOfBxi0w1rnUx+cWteEajJ+fAt2AaiF9HkQuLx5/BWxaFkHHRvfmAryW6GFa/
OypsH1cmafE3GVwEaKiX82rHphBhiLvIz6WzjFigFxnq/PIJ6FnHeZl1oQ1/DawMY7YKXXEMU89/
u6CyQHhwS2wssDrL21h2RvthRWeXE3q+3HbdGSzeBWuXGaozFcb6BiBjoJ22yi5ngfCBb/Ena6+G
WslBwlHl5ppqycFlFz56IeM2eAtcDkZ1k8evWz4n9zcitejCy5/R4gDLjPoj1rXT5KvRo/7CjAlb
1qjmh8w3AGT4UUJlFX5ibN6dfjuex+uq/gWwv8aTyF0yukolI8bnRJ/+o6k4YGV18kdv4MKHYeTH
vTxXovJ0FBKKtunIl2+vS/qK9B/gZCzH8/Anvn8LLawBhD82B8PV31ppoFdwWhU+/WWVDVJsWIMT
8i0v3S364BIYYECKIAKk1GBIccA+nP6LWOQ7Ga7XC3Gdc++RLcxpzixFJYtkeaByY/7Ccphp9LmF
fHYyaFMDzJlDsHJmFI//g1kZNwoK/2XbUflLv5af8qUxBxBdDO1ubSUQd4lf9IQgkxmDqPSELH7D
ks5rRTY9hQlyGDno5aP5SnL9sYlldzsOay+TwLPYgSVDrkiwEnNUKuHS/1w6/YOqfKH7N2NMlCDn
XAVvg5SAbhqS65toK+2Pl6rXc7tKF0DgF1QrghZ+flYkwwV+genXmNhvVqK22tbX0k1per0Nr9nw
OpbiXlH50y5kzRJWT3sLiyPHz4bknFslzU01lOZULWHJ7ZioYxvedj9AiNlgS/7IpI5ZOxWB3yMf
PRqfAzRXDX9sPEXR0/GX5Y7qxh2YLesEuuXZo9rtJArP0+96JCy6pp5J9ShCiZl7Eu67ewwM6Q5p
pIIBgu72emVpcMbHK/App+B6Gby91TDYufoXJRp/6jpKcwuje+63q4zc614WZQa48tZ1mQuGnacQ
cib6a66D6KJofILQacQPgGdCAIzCcpSv+hqvzOB+KW+Nxtgnn5vun9oRVSZ0Yt29z/muPxUhkABx
M/y0DgL8vGiIWpI5ntJhhJz64EqKTnRwTTS3N1ph4qljRan8Jnd+KiymnvM2nuvtonw6Yhk1CdIP
7nGavd3fkrSlc4lNWTYkRQEkFeg25fNLRx7KuHvT3UCYHVsL9lW9Vleu0z8qDaBAYgov9WdRlnVL
sUAvO0/5HJPAtHJzK7bmO64ziLc5EVIiqCIco9Vu+CWzdiIm2CHPin2Bg+s/aYan36/x86+vgHHz
iPz4h2JEMlrBBo3A8hdj2fgMuG6dEGGx9prnpA4q+njSLbZ6uKMuyuLM8KHcsLwb70cQkoyW71r/
H79tYmYy33sIdauezZCXNH9mju9M4OKQmXFbIXg3lMd+ZvsE6zC+aQRJT5AcUGXDyJBOI1ULVtrK
H29YNSW4tUihbEcXtl0RKsIa/cS62TOz95SA0zgG0NnKF8F2m5xpAfrl3mLRZBHqmwO5lR5Eyp+d
seS207Zt1hikqPhYZ+3kSmjROE61nPXNVJzEq30OYCHmHyO86nU2CBy9nOw7zABgDBBlfLYXwSZI
xpk0hXyl4ZBdAFpJYFsHbzhAJXp/l2BWwpS/ieg2Ha5rP8heYWOmy3wyFhsZLgN9gcv5d1LRHMm/
/pRUwDg7Kn6KeeOUt9rsgcAc3S8a2Kn/7Iwc5Ox0ewplcPZE+mMz8eD922cOLuyKhFBBKvkaVR26
PTjAN37YaA5gtRBeubY4iAklLDR7WquYcP7H4ZNxT4//CYz2zl3OKU2XqUPjYRHV9vlB7GqPtbRo
n8EQiCFedXsaPEKyBTmyghtC8tQuwxCokKzGoaodnAMVOo5KHPMUl0lmm7w9E6VTCykQmc3OgAXY
77ZEehaHnA+Xzx3zvbL1CyOHXYYfH1WPk5jOuPfZxO+wQuJxknBJUgzY8RnISbq3jwk3wyz64ZwY
MdunfG4dA8uQig2G0gfCpwpkOBORjPWUVR5U2aEbEkQy9iXeCMfquX/zXwUSs69l9NEAsz6cbw38
S2x3ZsygLuveb3j4KZ5/B1RQqkR2Pf49vGqXGvjYqYKB9PCa4DGyR9vpHtQcKhtsGeNlalp4ZJ0j
GB4GCfxZl+owPAwiI/8DnLaQYsgZVJrjExKtYLaNnB2vOAUq54lFfNrC5rZbF9y1Z+KCdyT34ZJW
+c7bi3TDK3mtLAmB5inOtbHE/hjxLED4EKls4tvQ4/HoIE4J8oI/ijqH6rn/Cig95sj5GbS65fn2
eizZRDlH4h4fXQC6XS6lSHwYYaOcTJ4pHlOdVVc2EFJ+Umc71gO1jnw4/h10I6A5G/eu1lKX08zh
Jwuku1t0UXyAzEeigDX6FvOBTQWYP5rFAECube8rTu4hMslzNBFw13nGJAm54eGTdEWZOEQWN2j8
+dfzRvpOtMvHgeQcEpmAX4TeNifppFtrKQmeDmmsH222BMAccYVqsSWhicg+B0oZP8OWMgfnR26T
3HD7QLdCFMej06OqJThhCwS+8EgDGgVT7fC8VRzPpCP+yh7wBGlv44wKz0iNnbUjSrGfdPYsQXQU
2umpK5U+UZ+4pILSpLz4PWjS8AkWwp+ufzGHe6gl5REExWTOEd8E9qI2VwfIbfJ9PEIVyzC8luZx
nOvoKGrJtTWkrH8+eacEfmZ9MqC6Jswzo9ziNBkUn2QmMlLIVq2SwqZj21hrkxueUm7HW4igRZUX
A8yFzcYkPM0Z6A+SEopyN8BFh8LBBrIF4E9yE+Wip4lsJ3PrA7gkdEOk+UZLJcHs8cCwrMWselJl
nuw1AUm94bWuiDUZT0TiZlvmlq8XNPso1uwByeAulKLRSqUhQ1p4qPj60i0yXOUeulbLUXcGU7Ov
8485FxJuDJark4xFXP3STWtMvfTHDi9qrfEfw+scpo9mf47UtSww9cNzPJ1hZ5ghTzDJmFALOLwj
xz4SD52W1X4XvtxMZIOidasx3eDKwTd5VoE3y7CYv3iMkUIJsq5govz+HgJ6XE6AYIyfjIQrciTU
+3A0Z983/fkj4S8ZLIsmermvxGePSMtifVpO+vxjXo+h2HtsGyveE9+j5iwQ5vcnBv1FEq7FfkbN
l8UkP+yCpTeeMwM21e/buJLW0yKbCS/kVhGktCBCo8ygUsAOGIP6iDIVQFONGxuKuxbENWkotrRj
NLVN7pt9IIJdHJ6Xpgs/5CQWCY2PF/XUM7ZgmlNvjy8vvzVqCkRe4dvVyOVd+7EJYb5i+9pnQq6g
xAmQUtiWb0YRiXjjB6+zg3Ccy2Wu13B6Rj7XPPUtzjhm+uYuG7yZO9R4OaJbZfZF8YtvzyI3GFsS
Y7GdI2S5wj/Ya7PYvlY9/cshZd5szfYy8nZ/Q5I3LZddQcdo0ryhj1hRxKxRUkNF2J9Sxwez/Eo/
c3jqAA2IIID+aAbj4iT8N7JacQs3As0pUhKDUJO8N2fbAUzU5j21RC/B1kWM77u5qEEw51smiO50
nmmB1YpmbEaOpo8rZJbbGorCl3KsR8ojoW68QRps8NXT+4t4pSBFllUHpPYp/yLdSG5NKJm5k3q1
aNExBfDyAKEm7XCV9h61BGapAPSjytomq9hTVGh9eYb4KJHDDvqKlS8RKOtv1OwQhtg5hSFH2xGB
8cclKqTOwGAlTw0Cr7XSOmFZwksyZPwHVIbBX/THEa5dSK0J2ggOk01n8JlitPtsB2GaMA0gGCny
o7X6a2WQl38b0ZSl4YSb8RNV7p4DnhbeSEiewWqYpQr4Vpbqt+qXeV2v+zF7z7R5CluKCeJwOmKC
3ZeOls/bXnhp7NeE561ZJlsWQu4lBPZstUNiMa8D+qd4z6dbJEcpijVNLMCUufIjcfCfnIRzfEtu
lAvilWkvhBBDxcriAnSDasV4OZ4mExPEBXaRpD17MMYbeOCIftFJ622bMB3hxwTRywvDvai5I/20
8E2/pTLV8hz/HSkbem9XCXR1l4hIrrZqirlL8yAzgiE1dsaIzUR3iOZJBaR/lgv+XzJn80De6mMS
WQoQsjtF2ipuEwkJchpKbZZWTOvkomRMOx3iHHRnxJPIXEgMpxya0664GVpVhkbU2p8rgyq/7pHM
/3ggEcopBmLJPd2ZeQJd06/iWO5pDKhzyNHJbH7iqO7tGYtYoVYJKcndAxlFWlf2spn87HmMfbP2
bIlXbhG/uPC8oloYjjSKx/9Gl7CpGPsUyMNWiQ0N5SjG7w9bzl2uHGNe3apzGtZwDG50RkiAErAG
k2dMPfdvDQpgTRz+gcbPMYhfNI0fdxksDQEMQ1geBsMfD9OCQO2UMNXoTNhHLQ5J3XN6QOrfAoBE
OzDmP8pz2oPicnh/oyer4AS+mjCu9MMVp95IjOABOVxMdmC2ZKXqybU8M0Z32BoXEjQm+OxtGXZb
zK++ffobO9aGuAgjNwIJEC/men37DYRQQ0eSx86+59/KOjZW5A76X5FgSdwBY2hhnL8Noxjcafyh
8RFTx3Fpu7ne4doy3Sejj21k/Hjrde7EdPknSUsfjY+wE8EL0xELCJLFbHU1prOuYkMkvsUtwimJ
botiE4loRcL6OonO1qmTgw8tmAM07ZfcQrYQ2F2inBiXS159sBZTjq0KDcuyL5+YFiedn/lMudor
UnhyD/fsS9LnRQ+7w13tH2Vb55JqfQXSbfYe9T4s4JPGPk8uOIqHxfa54maz6vpDLWavLyGiPTqs
E1REcw3QqGftpdbf/QUhNCjUAgo5raEBDhuhjp2Byc0ToWM/qQatT32kNbSi2DQtD4vpYzUfEvDY
qXSd4rWMKzscGcabwLcHak3ydQWueUB4Fab3GFT7PdNYvE0z4fwondXXasNW6GCutqofAdSLFykC
qFdjiSujpgEPPegOn79+bhmh3oUexY0FJknV7eRPLcYTFc//R2Gx0qDs2S+ksaHKsZjRuMfCT8JH
z7SWeGYI3jZqQECnjLmtSkG7VOpKUDTSJZi9q5p4iMiwgbefOAnqSBafoScU4KyZDAQFWRLaUuKE
BrqplvbBZz4bJUYDzAn1GzFRmmDUFRDVlpw1CTEArNVPbhRkfbsYOtJuWyz+A60+tJYcUTLDgwzg
o1hxchUnPPiSrZJhq7AT+qd9xgvCRYmOj0PIY+DSWOGYmsOz1U0c93YT/H8G1B0JnRqydMBC8zpJ
tIEtU6IZhslNIf5dzC48d3ediOv1J30fluDi+y+0HJc7a6uM6OUoBI+/OyImO20aFhEyrJouYBPS
OZveS0YE5mTztT7rG1HG0nNo9Jm7ZSL1E2yKl9KMv/W/lkjOBkHxSjrN7lRiEbB+KURgwYe3gSJK
0G6Wa9Ip1DxBlJaT49oDcona9SLakgPgbeViS5edGw8id1g8VKN+7NVUq7WpYrQUgBHi2Xbx9YoX
IXZ48SCHF2fR+C1f3am4CR7g+1LahTo5jZ3MuJ/Z4x576JVExZ8O1hjOWCf4lII4ioAfFNbOWGRb
ZreqwTdxBBqEUXQVYyY+C1WfoMZi3bDEM1D9bBA2yoZVSmLV2xbaQ9YeGtXTqztEEElIAhQK0GHg
XqRT4rHMcmocvvk3tqB+/j9JlgYetCSKc49f4okAvoZ8VBvdaDV6baEbE2AqAEz4qkZDa27EN4yy
v2o+0hQWoJ4Ei8fOv6iSHZhmEuVVk7CKGNXD3twcyKu6yWSPuLtYPdyDYUfKl4YU/x4FtyXrRoui
oRzc76SE00P/CRdjTd0rwJGiK9uQhi8V0gb1r2YjG6paFJQ9qkFYVW4BQTdZwdmUd8s94Fcyn0H1
cajofcbJQ209O7NBcMpVmfcH5iD6vBgg6hUe0eE64NenJQnfaMp8+RUlc9vyu1KSZ5BlBtSeUNKE
wtBnFdSnj7DNPHeA63aonGorBmVrLzF6xNHd5GiA6TZ+o7V2WTh/LVI2qGdydLLvmxGS4Ay+WS8A
aJwYTJNxGYxprPMBxgDdkFn1BIAax8wGhfTrzAjBEn1zIIlRz0whI+yrffPn64JxeGLE7v34DRZ4
+7CF00pN9X68JbwKm3uorydbYnpnefClo8hZ3h+wIWaSY1QX+F1eNn5COUvRIFnPAahcXd7GuRt/
6JjlzK83kUApG5I7qBxHapEAOhvBsMSjhYZBFkuZd7yXUyp8iVov9zwAP4xK22cvd510gK2fTQWO
eWX62k1Wb7e0nvWsTX0CIWWk/HqHQ8kZYBCFjKGznrcgqWpwc7r/4C6/wTLTOBrDKixaDZ5efEQ0
93Rr3qODowFxxGo/mQ33LCrhtBQ0ro2mKGLbAt3aW5KXMZ9h6SpP9+/3CXByJv0lkLpOjXTLbGEx
O76RMhkzTsp1zMWfZfs+Q/81Ac9H2Wv7Q+68V7DP3fOi8228QHFW3Y9J2eNKIqonpzLYZ2y2ukWE
Zllc+bRYVD/WnPd3rfH6CrrGtk9LR+9k2V5aWr4h/pqQxIAR5Os5MX5lmrsUDVpJiGGX+/w3RHSA
rP+8qSOzeHKg7P9ypg823QbY8qOjjwB6pC6dFzKKE4G13DGVlgKtgk0aei9SDE0TJkUOdz31IQvb
h01u2M1yi93HIaVlVCFvLY61/Zxeg39a/mmloukYnt0TRyxPTt4C1Ngua3//JrATAduc4pDLgB1g
yP3qEOxJs7oaWRcNOtE4FubpDNbUPBnm2e9BRTNYPWqqwKK4xqA22u2udXX3OXoZAcTD3OZaVbjU
GjtfrbgoB9YW8uuz0NSRkJBkYIunoAYhrAT1hGgVzN4ji1AiiamI8MjqoXW2lEO9H8XP5w/t1NDN
8Ugx9rSfhlFE7xKmKqyZVHzF7DoXVQsA4ZVC6owpG81ls9Rz8JcyABFpGNWpU4llvgPn0Bvd6mNX
8H82fkpcDuHyNEOgk4y2d2MPKBmZSvArSEnt84gPtPc7imaGLYe6Xx+nMOF1UPw5R+XZ45OYXIbo
/TbFzfR/Pftw4rme7WptgHqZ8ED7z9oeAoAlX8BzDvivRSWSQ7tRX/CpCeMw01Oha655cu5g5046
8QHmj4HmOHHS+1J5dejtJxCR1vZLjUxBpYYHieyFPcb6vLewjP/1LywzLCqtBfLQ7K6VKFIbmFAe
RVR5JLutZEEEIJ+8UyB2Yf8dfOguSyqyV0t33Ijva+7Bt09HPflVpzjRm1XwKli3+Y2PB+AvrooB
H7+gpzNHqdj7qgfsnSO9x7XG62Od0QKJ2VirS8kyv/GU7ymcPm0Hcp8NPgnuBi2CKfSAStFz6F1v
REYTbeNLscL4I8RbA2QnrhB6daiP9pVEAO0L4S5lCcNapXtFdJ979hargdlodigkMyEYbNEI4wvA
KGBnuO3CE9sIQujQUlbF6hJyjcmQnU/V0nIXAu8RXaRWo+vbsuXVHyi/vVwv7CsjLDmX3xf1KOT8
Xv0SSu09HpY6sr0B3vCU8uuo+6mF1UCvJJh2sQgJimXzJojt4b8R9tt/hJGiQTO2czB9Ze3qg2Qa
tKzLAOZwP9oQ1cxPyLf1k8OtST2xcsR4KjZHutlnD6TTQHhXc7Ja2T/+qikHbwDZtvXyalHM8UMT
5nt7qDyGs3FzU0rkiC9WAz0WML+VxMASVaQvXvhOEYY+33DqH/vr6IJsaXash9zr3ntdWTVfhvkc
8wzxep2OrtemWDDYDsXckk5F5m9EnSzL8588X3Wcu8hSSuxLg7UixhIq1l5oY0BQbROtoYrjeURF
aK9Bo1CwxsUwoI7ARsrtglYyfG6QioKo5qTin0Nk8Apk6zX9+Ibeb3pCEM0bQRwTZTD0rdyBh+w6
ABlQPZsu1dBxpJ6PW+gx2DHk1OFVD/lAUszeNTd0BwGmASZbeLJHHE30K6tg4tk+7rIHSGn2hgLE
e5NOP9FZ/a50WHyY4uO4gnvi4eSDN8ZFQg+TxTs/e7sDG75C7Nw1ti0QX/cbX/hof4jOxIyI1bd6
7Ak7u/97a5sHMqT1SVm3WLhIjr62QkWtPub1vNzkh4U5lO8Ms/enBo24k9Rr4nw6tWpRAFRibWbh
c9VYgniHToxYAP9+UB9AVFjI9VPAR4oAQxCS2/t6zynXj2AlPx1wboeiBaTtQSk1wuLmBP1YehHR
ijGHVWb43GSum2krE5azacl+x/il//iKk9y9ZuD4avRnIvMpFhbPomy72seselyolIGcwnD21qGb
afdp5l/WER0YjHQM5Ypz8ntg6SUlkqomnncG+55AfVNBwxMkUXI1cvk2LVKxD9yMJ+wiJ1IDVoLN
Wsrf7/3bZQQWsOQqVPT/lzk8AX3MNo+cDEnqTKOlUN5st+N2frPFEvu8GoMhx+oSuVHNYu+NH6Ip
BhV6JpIrB1LdUEISqotP+5JhxvbB+gHfKnZ9nB7ES1lbAiizq/tZRgqBpWnMOnL7inCtGPxFFc9G
UpJjZx5RJXHaPQ/kQctwdor5GjzapjTfTHY+dEdpXwLDU7Ut8Y60xbuZwBvScrR/DYYVDKTTqD61
svFgL/0zYPLZ6Ojh+cY18Da0z4KnhYw/CMrXYGnnjV8l+msBqxBny7X2pANsJQJo9C/gnOxxU7cR
TfnXnEvWkNkH+z0hVNu9XPz72YWyPMeOAECwJs5rsylAqoXXPmLV1p/PhmFFxfvdVTWvIcFgc0vI
YU6rS3d+aQbKhWVaKmHOB3GjSzgyiYlSPxqLSk4nQ8SZPtXtLAqmkK/y+0+lSrHzxinISxJJztMa
1kR8COeHh/Dp45fUa+CwgVnrWnPVFXy4d9fPblcn2H+Rboz9U9iagEfl7DRMa+mirhn55ph2L0YU
MiLzk+kwhNL52EMGj89nD0raUeYPnvnluKqvMlSApTL7Rn/CCUmnEwtOtppha6sKrRUrywtrkPj0
mZhWkznVVcm4pDgbeccFNFdheartztfRq+ggncBYR58hCQRq9v+aXhnjfXKTTTfeacKarYdhqMZt
IfE4kJ5Zi2e27D9fWcerf0XtVqyntZw3wwlq5/rDAerlivfq2UBVtAg8rlV89qWZ8/GYIXazA1ID
1yDNNuw9UtS/vIOPW/1zpF2m6YwxRSJV3VM2vuvtfQQnz34e9sDG++JVJ15u+LT+BT7nahrEX6d/
JWwEG+jmzEe7ck5G3MK9UJiBzVGIy2DPMWg661SgLbMdaoobjMuURqcC7BLF68hDDHSjDtgcuylo
1lUQEyMhrLAaX2lfwy5wgUAKdnQ7PQXxh+jHJ/y/HgWUMSSJTaESkGKaYLX429C7K2grg0uIRFjW
IjXuXNmV9Gu1TMtNQq8ErLPnLKfAS/rU59TYBgQUnFmQvjGgz6mMf0R9gfxFMooI9dk7XT/a2BOY
6cZIm5LJ7Qh6e6s+n6+oCP0p+oBo0VouxnP2yB2cDRvjWDYItKX5nG98bfkzHsSkOgIAChDIlU93
SEw/m9G1JPP6640q7CEb8MXl7cqehC5Xfe6gncZVSvee7X1t3TvqGNIoj3uQsU8ebu+1QtiM8AC1
ZH8iL27CgRJeSZYuK7mAua5ISSAvf+E3rJnVdSZyoW+lqnqi0Vm+TC5TE9ify3kCbjxxs5uEPauC
uEYGCB1n8grlb+9r96Irc5vlRuErURxaNWIKbGKwQ0/0ZTK3HU84xiGTi+ZWVyN/YC3VNOX15vju
gGU3i0pTREVx2ug3r+nDiYiUnW0Q9rjSaPiGTF4whTSCYBMV/XNyRRgOh4aRz+rzS6bC+UHv2gYo
PP2nDZUwGhbzv+QJnVuv7X7o3UZrsWv6/SwtsNbb2In+wP/vbgKOXe6MCJ/WTiZlB60gPxG5huCw
b60vIE7pw7vM7FhdV7mXaQ5FCvp1mOGr8tdLzAwTP9XCNu5W5dv0dUjN8Rj5bIEipg/Fo9v4PkmL
gRylYik6t+/AXNQVcYWvZ6LwxStlc5peVMaSKxiZZQfZYWXSP0VlnS+Ih3hYcSoO5508YDWo1qOf
jif+SvNIzFzfmZvVo4LhrOp1uh5Mqzjq+VLUK8iM/ZMngqeUSbRi6qhOfdSpgtjmKWKrse7NomVB
tsHW5l3/q+PRJqexALLhfmSjAaFJFfN/+r26uASliIJx+t5b+wB47UOhv3AjWxTGHqLGo8BsFbFr
Nwvd0Q3MAlJa3RZWxv+8PCDmkJ5I1Z+JPQUhKJYfr8ViY4hfSG1OxmMdsXlkxu2ELTa45r+AOuI7
AJjZpTNCDywBUoE5VMecVwmw946c46IY0S1n9EOvr0gOoLHOgUUIfmDwcUP/I0UD8/SEn+BGYHzq
vmk1SO5/C7UonfAexSv97ENLJ0EDm+7jYja6kp0Grs5jEuXduC036QdV+jZOihYQKfpX9bWCwoZW
jE5SraRMW+TijWLPcqUvTecLGVFXU2dROMVtGadvE7PPtGDL6sOQRXSD+sxWqtY87n0BKWPPcGV0
Sp5+F3xOhYBQeCzW3cHCdKpZ+tc0ML0dahRqeypC0qoPeMu6DJ/E2WMigEkgvvJl1sbi1m6k0mTq
YKXRa+/HkhiScJdd/j/Hn1SQPHqa19FfBKZ40wgywQ1itC44uWQRNOVu1sbo79SAQhUMYiQRJbts
JE0JTiNCoj4GLubBHDErOMRoiaV3686TVmcNqSKegMe5HlQz2ziLbQdHn4uja2jxQVuSSTgGN4Rm
yfueCBt5fxAiuvN66a//sZSxC3TlI9UfHhjYsywBtNRgbiGN1y7HJviRpk/qo3wY2BJgNC59i7qj
7qyDnvg9iwDQFBJckLgXKQsWyYmw7X3UFCnxWLw2vHrHE3CAFSrnm0S+LvKZU+hlLUL15OE9ASXh
dXcn9/SOrmzNz0FlQMUEN9WjjyA5z3d/wMYriFw41wBF7bcM5a5g2+8oBhxRxkpnMPiznmvPofIa
Sd5/xOslCmWrcjkIAunGd9mh2l/M9YakgsUN8S1Zf5hlG5ZeXuD5KgenYHsNkS6tsPW8M9+x6V3J
nGXdYidnoVHmAJbKpPaZn87DEopQMC4soaA1xn2viCBvB3YiHitIe5pq4x7As5y4L93xNVf0tObn
sBA3fMpiE6snljbaXx12k94YTUZ8oxztmixA7gvyyhP9EHIF7tGA0DlCWSMS2/gx6KDsGSDy7t9N
idbbyImxUfpn0guO4XjVQYsWvzUAZiglfkpUgnbfdX5+ojqfh2UzqdrQ6DgVx+KJt0XCV/4QfiWh
F1n8kvGfBMvt4pRIeLpoH64+wvAHE5zc+GQzU4jnURd+M5NAmuEkah+QR7pFKgETCCi8YhVDJFsv
RbAHl9ro8XUKGAzgF9Tn2ZhksfsCzhIJANvbSypL86f4nkOQJRIFS03Rsb3yypfYy2BOrm2lThGv
VKoFF3C5/+oXQFWcbWCNVMMxW/aXzbul7eMz13VdO9Qb1WJx2eMo+wKrqIY6kU9hHVYoIRE4sOzJ
/J7d7i5NdTxkMR5lw5It7ppguF2gKz8NmklJUAHrUqZQ6GKHUMO4OYGf0Zz31IeAKUcrWgz6Pq1y
33Rx0bHhJ29+IlAD/pdO7Jk+jlTp4oNV+GndZVp0icAoC4oGl9QgxyZg7BNclBsBjcRATuHbcM+F
4X+jm0r2CZHQwANAgBOmXwphcacJcrW7jKG1XGyjkTq9Q3KzZ2hN9L3FOCxv1t+cU3EVMBiQTPE7
aCHllVRYlOsJOfKjTqWdwI9MosFqvSt/jd7VHIuVHFjLioC0od3jjLeE+vbKsCZIxe4NdVsJgm4A
bwIxBpGf+uwlnX6Ll3WJAXI9j+UJDcBJopYHr8mnwnGk6UJ5Lt6XkTXYJhBnT1LDFjDw3lZ7phnq
hKMUxHYxJcR+kNhr2DkhUwFWzcHdH9MgiUf7Nre33cM43EQjel9oz1itF8FLvI73aLcO+OrWTIUd
hWNAyLTf0udZ7ZGoPXaaYzzrW40jtb/t+3jLLCOH2oU8DaTuVmUvfcd1Nyfv93/s4MbSZ9/XjAtk
ycx6ROJIZOa1Z7wFj/mCTlLBZyAqaAbtUtMbS7aAJl7e0VzR9iUsm9OGyilBVUqVtjWYjFYHHpFw
0A1iP1VgcitT7PigxTzIyM7DR2rYqEtwS/i76n2UFNaGSUEaCMRP1948sqoCtyi6GTm+7jfnYloi
Npm3e4e8i7MxFc+ZznudBv2+MgOrZl3fKcM8oCp6vJ5zRi0dZyJILa91B9awwseOI+H09Rw/0EO5
6hZlI8GgtGjjyLdim3fhmaMN/sIpKVRx2QOOWstGLvcCVJhF/Ad7jlPRZPD6oUn3q3KIR5Gfj5me
QokxXKBlGV0F4qC7Qz1J0Xde2nQl7VNk2i1QmOowvjWJ65Cqik7ASCfsp59cHpJ56LlEC3DhInyB
ffe+875BDO7uFGaQ8NV9Derc82UtWz6FkrxzYo53U8VPoRy10e9DbmXxDur4rorS9WuIjFjj/hil
4wqsVmAEgSQeMPRA4NhpGYNYonldHH4oBnj6gjno6b+02VIPnV9dy28trh3/QS2gaHzSdIj44ghh
ZaHADPxbAV0SojR1vLJrrIrPesGRfoQ2LHr8cBkk5X5QbTbUscayX4EZxFAFbiDAtAERp6HAw5Ud
Zv9hddcWb57oODylhke4IHKrL7kkGYi5KSDmh3jspKuZFEryMjjMQZparyTmIAe6RGZp4qrFrYgv
yfNFfPA/v8FHjQlCEIQQTsYUOgG66psQT0ufHrRbvAIgmpihrPO0IP3auymW5kYqveu3kUtRGbZ8
pR2Dj/taYKAc7iUv7ojF/csYaml4fSMSfdMd9AjZqC1JcLE4Y/9yPLf0m+KOK3+T463RmdrdXw/1
w02JbwDdfiMCRf4ZHlag3Y5KBLjbNMKgqWVuVkvuXD7xpegpmlIwOjY2Gj4JAj7koczqyMjIwREO
XTE8h8HwG5vYTXCV7XKpiz85nHDlrea3NGFwKDgZCzrcuZ8F0WI8EeDiUeLOiIztn+Mzxey0ywQq
+RyXYS2AItSHcrPwVuhXyjXaTEXC5oV85/EwJkKBMZR2nuGqcI+gvLqiyPCXA1SxOFavS96zqWvF
GSWgBJa2D5DNZ6yPBzVQncyHrMXhoBYxAUSVxQDRl+okeHOX8Z16ZpdSwTa5hlEXuyBm+HW47X42
+oz95S07gcMDg/tcj1DvAfGchMVKz30ONkYpStUCMMPFHp8TZFOeUeWGSEDP+yD2pngEyjPwNx0s
iNxsjXbwaU+/XmCoWYf0bIPO0Dawi6NNF96btHLeqqiB9AvsC3GiU8fcF0cbD6+3P3IknttmTI3C
YIPMXf7gwOF79ZdT2KevgeFj6qUQgWt7edkbNRJ/6H3Sp+C0G/zvgnh+n/gb0i9ClH4/ZElSCV95
W/9p6h2hcsSefF74fz8ow5kUPZ9EK5zkJgDjrILdZkPkiXUStdN9FhhFiszi48v7M5Rb9gwcyP05
uibfaaqlqMa+74pN4OPaGO/GqqH6Rhh4zHj34G+DXJo+yhIxF9s1Au0u/KbJyGVC7ztu+LVuS4tX
Lr8ShAwmtDryXP509xonbCYLB2GHjBnQ71e7L1FTFoWJODWr6YpyF+KxuycMP7xv+kIu96UdCdcb
gNZYVh8Hdl+bQmLmdK9O/FC706m1g8ZhSHylVG9Pe5GhPeJXrtAyeyugQtA5h0BLwSeKSqsJRbG3
JpbZrqMpCvaVuq/oV8/nTrgY2Y3MCpuB9xuyvcJLWk3RfA9Ec0cRDyzxu+yEJu8Vchi3k9Quw++L
y08QBVBNMDzKouvsbo9OPhV2rf3KNzfB8te5xyqcvUqOdk76X4fmdkszw7fFERjCaTzvztDi54e6
yWUI6OXr/dfPqMXEDOw7jRuSYwjJq8uMwirG8CO5XPDki5J18c7Ts04NOq3JHyIKbCFbkqVL4D/E
9nleieVYYEv/ly3FR+4ktdrkrcW2bXLEEczLz8bV/zw+Ni3hjIKab5ZOdplZrIW7RlNfUR9YNb8J
Vame+82GOd6lk/Y/midCJKqK0v0cuGE5ZjAT39gzi/eVKObTVn6P19iRwOTVOBdzI9RX7WH1Lo80
zNoR5pT0bn5kzP93H8iH693BwDpK+tKi2b5TzNz38v/zTZxM3nbrsqXtiJYuirMYzG+1M3UzaIKh
FJf5CFvP327/j2R0SUPv9mKO1afbHPIDE3F76wx1cTtQRA1YZsbHNsz3LLttCvD2S908lF2ftnaV
H+Kp8pRHBSDE8TnCjNvqXG61lW1Sq0vFBtc4at2OJbgD5QR4qTGfua508OQtNGPIU31+pgYczGOB
yfdsIp/ZhgfpZU1n1/tx4Wff+pqiTSYYnuvvEC/ieL2SPRmHQUVGU3041K0FAltULwSlKavZVibg
qgdNbwcodSMhOLsMHf5a5Bt15jJCN1YifVfjOIEOiIxlGZc1ZpjoLqHOz9kCMC1jmdAsm4fgPe0P
/VK/2rGeUmUhh7x5KhtqTpV/xkhgUhk0AawPB7XKp2rkISiOCNpPNQgWBPR8bqsoKmicTYZqn4LR
u0kYKDdhdX/PlwckllcP8m0PU6w4JIIVaA7LTkbtXs4Aaksr4NbBWSkUZkdPyz0DbxHwPkFiI+Ox
kcGMjTRaebLFkZcsQC2Ys+j/2lg0C/U1RTxxR1Ewa2P42oDy6mbLTU13rONCMOXNvzHwNWXCENjt
kvTJ65H6A/K9Wy9OtcpTEgA7NOJqSc0hOPvPRyYEyrs+aCnonPP+HKvWxdDl7ucyHEE2gP7FxTLi
jKZqZC9kbju1cqpJwqhfp4CxcJ5VXdqJ9PI2YF6r2SjpyfJoNIyTTqGUpKFMgwHPS0XCYl83A7TB
n7UfX5b+XwTv/P+pRTAC1Izxzl/xb1X8GBRT7uwppuUJufO9w44WJY/Vzdl3ArWA0teUPbKgbVgV
eogSTqGoh4DfqD3cDmNCJEggWrzM0xmAEMO1NrebBn/o0tJ6WpZ/P8jYsVH029AeVQczqDKF9Q/B
V36Sp2GnUxgISmcuIjIyiqTW+PjN3mStDFaYxiqPOJVru7nsE7+J7xbhsEgRckfUaW8QmhD1AwxU
/rOZT3rLgDiMfLpf0XAr25Fq5RH9+ZwJ6nYBhBqLQ1ZGu/E4GJppMjjf9DF+t8EwngWG0NOsdEa8
6hqkD+1Je9Z9xXWS20Ijyl27ZC5ohrR5zMtcb6/nqjhhx8ivKmiYJEPdNKO2PAY/2jSeINrjNSSQ
CmpCJvvHHCxJ/zI/S2xneP5JOvhmLEF4GV8O9bvPZHEpgYfh6IBtx6cfC5QzTMkhnfrxNbAShH3u
8sdIAfE0XYxYeKQfb3aSBOwbwNEy3XQZehhcQ1ZN1G7zBgcK3FMf5C2bFTvgJBwMl3FQRODqxPBa
sShw6mbypPFI56MAIvuZ8dO4Q+q7RF3QhXX5hGr8k56P5/HtTNWY5SM4wrieRbBYMhvRsUOKmfem
bgvLCcJXCfnC2VQaBGhyIzEHYLesWc5NdQL5UT/j/xqukY4n4o4bjl1UX9LUKwNpSZtyL6z/UelA
P+XeE0i+6jARcggOp9zdWDKiQdR4F8YO7RCQuAceilboBLFziQ74GCJ7RJhoEaq7WBKNlXKkiANl
Titb89toVAnDSVoCiQ+2I/6mm8mlEwWn1Ukecy6LAUQMGqU7thpDvVQHDWqR/9npUp1y7siNjp5z
Seokj0KcbTojL7C9sCLZTu2YqrNr65I1K2swNYKtFm42K4v0oP3qVrL8ivbgH+bKY/NRWZOkioSu
/+8BCH+kta8C/RXu0OFUAYUUVW5mzbx7/X9skCgPjZKUD37zXN3jpmqZHGeXtlPdBez5RpWQ7k/U
kqc4XroQUAh9XOZYH3mkOb9AgXAnsM+YoYYO6L+wGxBOlU2nD84GkaIgrmQP2TXrCnBTTHuLRk9o
XfZAaUSpUp7GDwsQUCBsyOF6u1UV1ewnb3qjVfhS1aPPVntX5JuP0YioWm1DdJBzw1U3FVIn1Hbr
GjEsBekBiOXrS05tzqOkTlCeb2t5Oly8Za83buOf0WLJGlMHikTIuXwAhkn63wX/FMin94byZk7j
IZkEOg6QvgMAPwY4Y2FD6/VQl0jEA0VvIgUYTc5Ps+MCkQRGCObkFBjKUU5PvwovWVQNmKHGiZ/P
2MPeDPqriJLrnWaD6zJ1L7fk+EU7Xx0Uqm8Fhs1FjaCjBmEO8lmmdvfiM3CZ4b3WS3Y4tYuvqV0b
w1YICFm3XSaceTIOwTk1IFfz79j7wbF1muzT9BbHM+Q95umbsxrCCQiy35moHOCHWV0VjZfOm6Hw
kEFDyL53sYIzXBZNCpSQwi1Chy3ysB+X0nwYrm+xXfpBxzsG7vsxzIYzYpvHEX+hInx3m6tYnLRJ
Vpw7kgto9ZhUgdncUpMd2xR32TkbHP3ynAOM490PbG4LVlzaYYx5THPBzE8uOl1q+J6d72NP/VvZ
RbbVw0/XGmRWbSBy3MtRD5VJ98QBztj1vjOoOhsQAC2QDsD1QtPHcBcjfVAzbK/I8E1okT/Z/YTn
lNgLFZd6fa7c/eqkLvbIjPZYKEMakmq3VseWyshplQIn7rm2AQTMo61imcrKkwxRGY4mQ6kkQPWJ
e1R7dlG8rfIi8YCoXe2ed57c+XBQM8SYXMPG7aJE0P3/QlY7ZxktkG+3kDCldFYvhe56OB3qk9fU
FjNIKfbyNx6tWwiCNTcOKwbky2pz/q2Ib+uSeG17RnowvFuDA/fHH1fXaDIDoBQ3Gqz8+uQK8di0
epmTTVc9Rc0KK3dBuFWIs0B35Xw6pVIth9WV4zV7Vzk+zl4r/8n/rXYUETmq7Zuy0wOFLLDjg1/v
bqPVa+wA04Dmm5zj+lFau0RHWsGdIXYDWZYNu7c1WfPr5+2AaeQmz6gffp12iHI/wQIUFYLhjF1Z
m19404x+nqUTVP0ZPOWYnK8yec9PUk6m41/hvQ1JZ54ZTvo+f4t+kYNlpnbRKVyKN0cYGitxENwt
Zr94twMvcsGjL95/ovfo4a/aj2k8KQGVMOhWxGrNnaQmFy+dM9rrcF3rh2LJMsLKye48Zyt6LdNs
I/NaPPNEL5r5y3/L5kckF6bDIBZYC5VHlzIukXOz3uUQXUQGDnCFx9paDsnKs6D/+f40hudUnDeI
x74HoiA65L6dn8jLedr1v6Q1VBKtgJnFSTrVxQbe2YolZkCHbM0/PBoHA6tvAndmbFCVE8wbqOnC
26BbTsrFtjeyCHKrQpd/0y32/lTSfR70btD29zJ7ugz/gfriCglQb0Rkg/X1muxVmd00jeC5tqv0
cwROhwV9iApa9snma50QrZM4H9q51VuQD+wTbqd9+c/5Iun3XSLZXs0tAeYpeLkmCR3B39xEaAkB
dJsApz2UUD5lh3XiPZ2sLgObmq0MfK5OLxl7FZJFgNNXyFcWA1su19HG5gY7rSvTxiBl6agBfTDU
fr46PGjVasYSyiuF7O0X1U/Vx+NHGijREqLV8g3cif1c5VWF5ike16O/SNMq0pTcJ0ggMD1J8Q+G
zjpNsUe13C0SUl0M2WMRKJLsFGvkbiQkQfTcy/tWg4tUHeXadhLOY6muCGJE/3TgMtXTcvwPtvvt
Lvdv2S1Ql7OHVMGWEq3Md2Vxv5J2iy4vgkwqtai5TZcBcOQnKPaq41hWTE/CmyKgKGQiF+l1TC9M
M7tLOj9il+k5GfvomcwIxsqajYxPJ6PEdmOHw1hVwOHC7gK/01g2Gp0mX1iPLJ7eq5GkwBON7pFy
Fv/wXLoKtaxnmURvy0fHff9peXy5xz64O6UpeXYTWSG/Iinw5EQ5Bbx51p/mkRP+r2Jy2B7h6VYs
bqIFTMmjF2SUa8OPEuHm0vgzbYUSL4j0TFph1e54nw3ueAzNF9210N5naj3j02m8EBiV/2H77fjh
RLdmsPkVZ8+0kWcEiIsU4HBb/xmbYe1A4UNKO+n/0c3gowSSI9VpN6jflLdHCSbGJQrHL/QRRcnZ
zMVDz+gst+vobIieI4OIHeClWGA2Yrlchj3lyjHeM5rZA6hF0ebypDx9tljzYC8OFFh4COUR0yxP
uOt2BQ6kRFJtkCThh4NpjL9oW4LyezAQ2Zo2n+zYkLzmkZXj3UiFC+V+zX1DChM6Rw5CTSRFjZ1A
46h/xdZt8cBpFzZxGRx8bwJHclIX6QaGxf6e0A2muTXL2BwPa8ek/jB69QLHajhwCSsdDyBgQA1b
4oEUfUXopkGD/mZ5R0jN+kfuD3ji95nGu1DfQ1oOmEedselkGNUDibfHmyROp86vBDoBCOLQu259
Jx0/i4d7Kn5jaJ6YwULHAlasjG4YnrwIp4HeorJaL4qK3YAxKWo6oKAiBukqKtfVqcSr91/0OWae
3aWV16gTOtaRH2l30O5Prax5ZOHeDQK40/eMIBSZQZ2HiKoXgrEhV1KOdWhpIYEDv7H1C3ymAvY/
E0xbKD/kXR3h7qJDl5xWOKFJuC8X2v2LSfToA3N4HM4sy4Ca8E7lP6zy62Ul54oICG2OMGLC8ftd
eiXsxTxHhy0MpdxoVShcUfhrDWN/R93pTpS0JRZZlzNDusHq5cxAIYFpe8gdUEXNl+U48xbAtMKJ
54qcH0ZJOzxB8mwxxr9/F45QfSo/HyIujt3YYLG6AJ3CUFcILELHw+7TFB1fmlx/k7K2IvlYY5+p
SCN5xsI4yLKuk8QbBac1aoxw/SDFMRStUDVj/RYlLMaLziSaM7ly2eQMAvCJ6RyQyWKGDQJZo5mU
s21W02/oDHMB+heG6CnxySBedcGxvNkW2y1hEflSZAsXwAJPXM1g4lByD+s80Z8Y9Nnpzt+EvYbF
JoB9XW9dR8N/ZqlWFVDyFLWVXIj6XCYIB+CxlOcuMyVYzcZN5tYx0OmYrl6FkQvGX+kHGQVylxXq
5WUG7+5XEyYVCdikaryXLakKncM9wqwtLgaLTQ9sRrNoPeXprrL3lzvnZpIT5jdNMm5LMl795895
ZPIM5BUq1N8uDaG9VmORk2XTd9Yxp4hg9udLdJ7E5KS73F81pYIeEdOMnIY3CVchFbHZi9fNJgAw
4xaAp7GQI0BcbndfDCEWYwbX77H7Q8SJ72OD/M8r7J4hdlT6QRuzgARicVY6ldO1Dyl+GKBdVk3B
/Rb1Eu4MruJGh1a0xnjwHSb9sk8hD4UzMuTvNFJ/uP/Me5TgH8PJc01Ceqo59XCXF+KyEgraU/tO
ioPSRbwfKpKPKvRiSVJtz0fx2qjQoIZKSlRKg3MhzzOGjPbYhDCTTxj/kL1cfc3TB5vvDkgqlM8C
oCHLXc06xFpyJfwSTfcQ18la3w57UKnHjvtczZytS+XhlLbXPkMzji0O+YBWx//nLpMf7CG6iVfo
7eX5mbZ7+LBtrZ/QfUo0fwWT+2RZzAweBV9omLb7zraFbFtn0KjEugDgZIq4jWs5tj28s8nD009C
UfcsIoSsmIPap9+CNJEBEEx1aoLVWBHFInuR5eMqsjEYSHLW7HIJuSe4R/ahRWxjobpCgpTubOe5
7gEAnO3XI/Kp0HVtDofRKj7JL3tmyrq9lzRODGYrEBYIgjH3duVkeyZw5SO1r23XC83UNZfivrN6
cW4cOHAOCNkJrrl8/W8wdX513AY3aGqxWSNfpPvIiQd0BDP3TJTSiOcwLUip3ozvsb5jQ9HBp+sX
eK+22FicYvUUWcaGkf437Uk3lC/k4eRTohJB2h1PeVxtHr5xVjhlz1PrckBJWD0bHrTu8fEPFOQw
xa5bTKcUxz/UIMZjtw9aAdqdv3YBnW9IVHmCwK07PheD6U0uzmi2q7gL9kHadUJaHgbx/AaVlq85
VaoJrF9l8ybrODWWRKUCtIE4uJiQk8+Q7GCKNhki2pFYcihmXRZGvA3lwnjFjPLIWmYRefmCXwak
q7ISOFoQupBfEHxHhNoBlJxU4A67IM9vMoz1MzagqhV6cPmUX4HgIiPTc0ZsR4tDr7z3evuBiPmj
8/99cKggqiv0tkPTYag9o4/7kx1E994Mbd6QA6Clw/Q+rnac+Bp+jtBDEka3gYuSblZ8zUWg9kHT
ULBYD9XzDbB/VXV7BivvHCRwTLR6FAXPChN/ok4GyZ1H8W1kHMi4ww+nM9eQCl4V6RIB550wDBms
EnwJVxnbBPOFgsOSJQisYIeG8ecyhqjQ23x958EAZwtG1SKxLMgW0QJf80pPxcPxsJ0xcycPvSp9
UswoRNxATA6Su4+j5LZKXfvqpaf5/VCfHAV0YCCFA6K6KsqKVB345azeqMqfKcSNx1KAsnO+UFzV
4UZs0ovCGWrvy7CM7Yrmo/YS7NfBh7K5DDi5XrjmnKo+Ms1o6Jm+PU8AnkDWQWP/TUNg5WciuS8u
gM5nMeldIQF+tXafkzwYQR7MwyUuKlYSGb0/NXwUHJ7dd5SRq0A6zsWT//lQagEgmDALG8Yel3r/
lsF5WpM+oDQ2yK4blYZ8FXmgnIGdYBkrA84dEzVmD3Tl6c5nQ/+N59CPr4vnuqQknSbKctNh7fQj
k2S3DSZzQjSwKAb4/cVGRNpp0Q1mr5E2eftbKEh2J4JUONuYWWGC9B1E3jkhAyntLlS0v/FPQdUo
WPODQ0E6ejrlT8cG66pEzM8CvPIEv5Vsw2ULURssHLdobqvAbSiZy1S1wjLdqmGIEs/r5LT1zzVI
JCkuzbGoHyIKIFpgR5SJ6yGq1G95UOP5pyo+Ptqjn9mgcA84igClzwiWNSrOfTBPAi25jdnIqey0
tjBFE7xl3bt/lDXbLVDPazN+Ji2e0tXZTtrcFOrW/d1TcSN4ynFBJKD+EXdX5CHOW80MzY9VyDWz
a2QFYC6TgnToA+Yos+yi6zPQF/jQiz2BBFv8eYudHTDmvNh5Lcl9yD9DHAWBJ/8bJIDcBO+U3i6g
UfMeTrYFm3noiW+d6e9yFTniV8GZeyNivAEN0rn/TZmBHbG2uUISr2fRHUwK1R5Ela+av37T6nNG
snvN+UxAk2Zr9mVh+X/uaEmQ0sAfeQADUA2aR38BPKFgc75HlI9oBZxmHqcaFFcrKCInT178wbYx
bw8M51SENQ13ymQhE4IkB9NOUWU4KBrqQt46Gasm7U2FW8dSSHcTVkH/aY2NHUdmgWcBzuHHOhog
W3shnYa17vI0tO99pibUhM7uoBqyqIky+lWAUcs8DKvyP/QmBmqqjqWW/Dk+FmIiBOdiI5jAiWT4
q9fHiM6E+pR/7SjFW8mL4uowNDnv1/aR7lXAxSO9T3VrDSc3aIOSwykq0Qo8BqB84vBGZKOBHSAi
rmlqIdH3PYw1PogsOxqwHsPLeloQJfl99ua6582vlfZLryZxPPGYcCxSG22luz+XUC5dxnLX7Ix+
rR806KUVMxaDcmb7s8LOp/vtI0TUPIRUU+/STrAgYIwG5/O9bTgWpKJWOlRU+c5Os8gwFG87MpGA
cxe4DoFY1TZU+Lwt0v/5tcyFAxUTKphk7dVUSLz/M2QMwnO/ffa/5eMVAlDMtuoZhbd44cseTPmh
6HytB56fw1X7QEva+d6yiniyswtKIc4zUXmKdYw2c+dj9XjgDd/alTfOKIMkUPJ7W4z/AnR205BW
FTOEvFa1ScaS87FrTM3lUfeRKgn78q9X60s8Mm2E0nxDyQ2NA9XQ7QvYjFtW1mwJmWF7IfPTX3zb
qQ3s922gvqXMUX71W5iXrUxFwUJv9uqqVmO/COChbSuyS28Muel1WXRSnAsayq3qGfTIVh2O48Zt
y24U46SuvYf7ysQ9SyhTveda4loSHiw+ZIyQG0aR0vpcCq+NzO8jgL2JiFIcXoQ0dp/SIdOrYq19
Oj7CTY9tCpljeSuDJRAYKYoDKXl+GeWCcvZ5N0XUdyyGw7Hidg2Cyaj4ZvqETqqcol1/0GnV8kvY
GY/ct/RUKBDnWJNAaQJsHGrCDUX8iWrQDuFiz3U1u4k+wcYS6z3RIRdxREvonEW4Olc8TZqA+Qur
MMryrlWlOhmT2mFfDHCGWCnJ8OWj2vH359RNJN5f+LGDWbLLHJwZG7C+xozDVFTDsPxqymimBzSE
LMR0YN35dyohoFjpTDmOAMzkTtJdCnl5QUDO6/NrzID5JCNU8z+cYaNprKQZh8IKfvPybGNNQS8d
cZbXJ+Kb3wQAI1qF3IcfQivOUsT76KjLOr0ciEgFhoSf9qfhsm+WSmTyVKLAJ8LdlRlPoiACKvJy
UgW8x5SNwdeRyOA+L+tFrPQqbo92kVbqZkGtARtpDzesQLqigUHYy+jka28Y9NdiW9rpmawUfMgr
7rTNfjFOHn8UEloyYU9ijo8rVRJyiSKpZ40fsgSVQ0bGxhKiZ6qStamykHpHEgt+iTQ9pnOysS/B
R5Dwg0WDO0YbYVEElscOq7+zPfg6957yNhqaUskTPWsL6f1pl4bd5T4dbEAyG2GpYYZnfH1ZLMFI
lAqp7Q6AVooZ9OLBnnStKFJjnj8cVohLMEkO0NQU+BjeS68wUVsXWUxIBGCo8l7DvvvvDHUqUIEU
Ygb3+Kj4rexs1G0FOm8benILJ8mxfvdNByCFskqpiVm+W6r1XjsBKXdrv6wwPJJt5MFUdYE0BbDN
EdKdqVkLIYexHfPu7dG13prePr/3mgSKW1pjco+LvmuOfXYVCkEPFLadWk/eOTE+wna4IM/2WMEq
LZiM81F+H2OrwHGOxyJS4irovYtP/wyKkk+1oO+O5T7VMojMNNpZ22kc/FENsP4kErwdDkJ7uk2E
crHC20TEc1hwfrfh/3fcTEIf9DVOd/qsFkFs2C1AE2pGVJKrCeLYU78uByNt8ybi1hTr+tqTzRyC
qHR75Rwr34WFkHybbEcHne6w0+rsqPt4MOaXgp/SyuiV3zk8TDNYeDFooiXRUNAjIgV9MoMijDna
Wqn23XnuCJaZsdaOlRm55+ihfywbikQQU5A65WV9g6c+3uF8Wf/vLTmps9OmFvZ/6UZuQnuiDH+C
JjTH4YG5zHGa5tU4pQLZ3M7CfOIRmUUTFQsZ8D8afBcRikYSBKCMp6czG5ETRUIrEW9T3RyWamn1
RPni9P4FtNR1gmkNK2kUsBaRaR3jhOU/uUtArpCuJqPMEI2sc/A4vLRL4UweUpj3HRpMCfou+QQl
K+YvkHDzj/yMY8ZEc06Rx+QArc6puZrNUyl6Sjoxj+j0PXRLHIySy35QT90e9LSkLF5YoPnvrNnV
Dn6VGUGgtQumJuf1OhBdUfG5GnxGdJAxIwFwjKgoM+XxRcfZd9C1RmFoQUsFO2EeUNera4SfW6hq
GoltjdmXBOZiynvYWwmz5NZ629WRFVytSW+Kl3BpKqsILwWNFtNGKoOCpz3ePXCA/vNj5VcbX58T
6iChgtWEMgxYX0NFxfMr5X59ys4kQQ/nKn1L3BjO47s9CmkoCcaTla2FtBv2eqIRt94gHe4v3DTG
nqz1pcn6KRNtQmcX9HXCQsdVn2vprCimEqpJER1yUV8U1ZV2boM0q9AbKppWzyvIN88Nxx4W7B2F
DrYGKhBDPh2zKB0Q4gU31uIoEHxM6ewJvi4KnuwB2mc79IEeSR2cesYKa0n1eUuYVtdmVeA3N25F
jjWDAuSIiK/Rcm9+CFihFwWmgy3AUOF5Ae2uCOHjMGB89EhQf2BHzCESFkOLf6EevAqJ8pQVsuPT
QVKEa3j4o7x2xRLEDn8+79z/nIgrrpe51N8gG27wx7PhZrs5Yoy7GBjTmSVgEhiUqvrGh4SO38Qw
CiIChV4NwYkGm5pFnsjj/nCoAyW2pkVUECcdFLqGdl5E7VGtPpfX16lI5nLLdANXToGy4ddZ25Nx
9pZ1emHUARLSmltWfuPJmaIAKgR8rpSHdwhs3aiXQTB5edgzYcY6qwJEFnnVnSPmATUvAFqtOFZO
ldTE+IX2dsVgQtRyoUYS7xK0JVoxwf75GjtmH4xEc3N0zmjJqsrFLoyX8d01cMrnq+xOm9tM/MuY
pgoAUYg3/q12IKeb9lgQc6BDnQQADwqBGx/5OPh8b5wmcKLNydLb31+H1klGSsFUP2BfqbrRt4QL
LOhMZq9M3RWV+uTj7n9zQZ5C57LHEef4EnbgeY8exrTul5zXlPqSASHwVUMwOYJkbzJaxtSuaB26
ayozJMAeh5zax7IUc0xsR9kwOrsqi3+4aESlt14+dOtkpkbLZJTFSDLn08QUbGcgLZLaRAjclcFE
oXLwOrYdL1EzKDdPwzDu7XeYWBuauLS+tkqj0A0GOSiXOn3bIDo+tvKkNI8AW58bm/41TAgj2DQl
fCUbp2aawoiPh2rLJAhmbQAlqq/zFk/VDb6se8Vp+tMEQPbLs5hncQjkHepQ8CCI67yRhcjElzr4
rBFolAfo1zwpem+IyQ9ApxQxQGmhNhQYYIftQ0MtN5e10nra1VgRm0SSrhQh3WqaJ07+np5Ch6DQ
am8ia5lD7SW91MrIozkLP65uzpWJe6eZQ0hJR6mA4bfWYJ+uK9vA3DOpWkkdYsx4VT6gpA29c1TL
DaHyPmwXB8z2YJr5fVSepNr+oO1N5Elpd1rUrzlr9h7cDBpXUAvwfK4UpKxpdCw3GojF1ibt8Ccc
5Yp6ePPOaK0hFAso2tO6tEmmH2KzhC3Rc+RjletM+LsoOjbjbSWjJZ4TY9Qc+Jqe5xLN/uj7Mspm
ZIuWseePUbdbNs1QJU5DGirlVFMY3Q0x+14kNt33sW72vQew7LDAAXIS/yr7Ou++kY47HVQfD0U8
+kjx07b2q+EmEz0qvPlq2H0dR3pCaqrhkVCwKRSJoz+pzWtzdl8mdMx3O9UAmCVifoR9S6TRFAJQ
1wMpzhFn0e2JAMyhRRyzZFvCKQ4l7wPEAweUSArdpWOkVly9bG6Zc5T+Ie+tJatJishGdibbRgim
zWqC9fCyiXNpww9eeVXGGRM4D+yyKGqD8oFZw2tG5j8V1zYTPG14bieyXDSmsoYCYX2KNuac2htN
u2JfGtwwCqC4H/cuMJtFmSbNEPWW2aTLMoS06eoZcpg/xrIsbVsPAlVadt529D68jPrB4GeQxeku
O2wHOjcjbseEtzqFByZ87leRoPT51BsV2zOVbH8pPAYSgsnCJGFdZsf6VqlZb3PzDYW+6obnj3VK
CZ/BZ/VVwD3f3wParkA/9vMYnvsbJHdr+pX3ZLueFO5kfxQl2Jni6Fc+KwEDqYlPKAChhTKc8l7E
EpDS8YEBKBz45szmPwJyBt2naRM+F/9s1crFIxIhBAe2tET+au6QUX/A7RqdM6IrpIm5U+PIalNm
kBkMtXY5/j7NiNB7YMJ1Rwpr+dJ+2qa2igCsmHUq7G/I5DhPCjUjWCqbgv2jDMpTUacUomrp5cTe
P684VdMbh2ua8EjIssoxzZW9OaFyta+gDyTwa1Nh0lt4QH2Fs42moKiCxluKNHbtxyjmxt3K9BwA
3zC1mQ4vM5PqdGSf/KK0NZRSAFFCpUlXRjWCpkpxeux+55AnCTzro4gRUtZXqF/yEcuqHT3abn3S
vFLOzlerxzq7vq5/0N5JzghRd6Ucb7YdYTo+DEXQ/qRXrSJDlwFibPMtULJCqUnJCCuZbS2nR51w
zHIdWCsWM2KIzgti9h7vuHmf7bSgJfYsBkMFcfyJ9QXJ585mXJbh9isJBciBUtCcnfyrl/n6ZoZI
wZwAU8jGypqRlyWuqWgBJp6np5MrG5kPmbxfmWcZEonQfiz3RdeNGwQQcZg4vay1qmNyBsbvr/2q
RMHODIvn1ad+YueCE5a0u7prQ1re3NOpRF1TxptTfxWHWF01lbA4qoh5IpT33ePEexsUhbKWcekn
qcbchCLsJqaBrkY6UG9bDTOcTlv1SYEAqMJGOFVe9YLdlLBEJiFezPxH3nl87aoF7AdElhURb73U
qS8dm/L9R0FCiZRReLtv4U9QnVMab/F9Rh2fjHIN+LxC5ZkKzfE9O4yN4ErscCyoMHKsgEjd/w4O
KoQtLTqs2Y7/pJafdZjVN8UZS/9vKxcoHGpyKqXOFlBON7yLI6lLaqCtGlvdRWjsXscjOFQeQrxF
lqCP2mUDiDN1RiQTmfxCgadtlj14BWM7hmGQITx2p3EcnBiw278NIA1elfknlihbtJhDTZwzx7sm
iQrmsVl75e7yELutH2tIGv3O3RxNHlQ3kq2TgIBj/dysOro8w05BmO9Ag0jJJHUI8TGCdRsVjOJU
ewqmIXAAiOFilQunnmlrZ+AuxAeergewFOk8UHRkkL6zgYf746LjwTVmWZ7HEthP75Om9+o+lZUh
knFGX1cDp2adXagbaWnH+e0urvCxUZdh2K4eLpRyZMXlWCJ+zVSXhAGxpHopUaoLo/0YUs2EYKCp
RwoLgkqBZwp/RXS2g8Z8lBtXqzLeH0AG6IYF+mQlw5A3B+CDcC244WWkHxTZ2+VgzmK8DzCQAgxM
4rVAnRIYSt2N1BVUgEgY0tcXi2izFDi8+ibjLQgNXSc9SMwIM7zPl2BLxqmW0OMj+/iVg1kUN4WA
d2X7lOCC46cfQEAt+Bc8yMr7rEfwIuqQqGSi00LUpNk15nhxJbfqUHktf4xp1rDB9p3kEJ67K44H
eTAcYzCW5/hhnkKvQbrhdLTfgvKN4EcvAVzFp3OHvgEnqA+o17sh7ninv1OFsxC+LcTrqZdBURlW
G9foH0S105vi6gdnqMP1mDu3oJrvO6tA4lIBjNWe3nz9iHuDVvFT4WqER/ZLQ2GAzCBmvEKXi4Ch
t/kUuOsUE9qvWxFDmN9EYK/6ozeqPL3FTpJ8h8GtlgDmxV816pl+SEpC/VWnDP2szJaiBqM/axvC
pEVdZP6pJuVo+Gv5YAyBWFbNUGan/3ohB4W/E5C0+yJrtP/X11uQYnRVXlxvzNQiVlTTo95dphe+
O1GOFHzInZmih8xU3VxyvnZkLmM3A5MqB1Wu2y3t7IhAX7MY3PpdkLTGauZg4og1dBQWZa6NI34g
cJlS6zXLrhyMQM9sI1UwZzm11fAXbWh32jR6pccq9uS+sBYxKw5nM+cUOrtZ1wxXjY+1EmGYg0dD
98FXQSnRn1OuuVGMhL2lC3yCEZ3Wc7b4q1BfojreSBQ6lXbyqFV69cF6kZ2I62cDypHrWfqm1iBr
odYeeC9G8va+vcaVTPziP8cQFml42Z0f69mRh1NJ/X8JzPds6zl2KSzMYDbt680Tvx+osE+2l8GQ
gEefphpGTDw7xKMJJksgzLvo1wL7y/UWCiwN57ZrzXpYDHJeNvzmywWogTZl+lLbvTaLgaRdnfCa
8mLymBiUM/scLBbDA3WItFvIUA23Lm46aHGTZQN04CvyFDwWYA/FilM8QJruiJupLLrgaP0pGzGY
UsVGO5ZFZIFygeTz8BZUY0gw1s2grOYfrWskfZaz1+sUMtqcVkztIsVwXXwzRr1q/iLEDtBr0dTS
BaK1j+qoW/dSbhe91BT7OYVCh3d7jGzbO9JpoMWwY5uwihJJywVzQgYk7GhRaLjGqx8wYtW59cPg
s7weQkacGQTLZIQnh/wk/rXvKxqZ5fddMDeLn6J6rzuOFcyDonaQfFXKz4npXYn1MZ9nrvvCFANp
oHGNzsII3BQQJ7bpkhUTWzts+xxn0gTkAJUXoJBCa3B40xfImMVQgLgB8+vRqzuoezuOwV1+2FmR
twfk5vnDdn7iFQKUbhAPX3at1UaenOQp1qRZ7eXrwkz3b6vPxc1+0mWOKAFtdERMhMTWqPqsXvnL
r8qctqPu9EHvigNsJ161Nzq2mnHvnwULHQUwhjU1OeYvXRwDJRnL6+KJwNltp6qm/V/TJTgzw2aq
wSsAeT+ULwgBJfFssd5KGqn+NJiq1WwEAXA+tXrZelI/3vKQrt1x2kTw6kaMlZH8cLK0pDKOGzwL
mhmHjr24GvxOYQWkcSuKJwOevWYSfpA6wYOLADxY+3d+envp09UwOmztvC8RMfNVpaBwE4+baIRa
4VKu4mp5wgfwjBQJ2zAXlnJ76BXZcyv2NnKG2+s5OS8gSHOKg4TIOwACgAdzMIAEJpkWeFdnfIbf
Lb3l2CWEAg9DRVjIEGgU/z5sbp+K5mRFK4w5/xPJn68Jl8P4vazwrU9hN3rdlNDt4KQsNqoORGqz
Yo1YRQCtNTCA4j/uuBdtubufvxtKr3f65M1Oy3O+It8zDJrubmhIAzpa/uYJ+lXnb6jOn2wQYcAh
nYwqxsremBrJCEGeTrQDAN/V7FYZ+yIN7E+/DUB+6PY7XHnCFx1B2dnXSaU/ML1ViFw3zqq0noTZ
Ggsrt8a/TryA7lypwfx8DGUcI892o3qnsgoUNUAEnH3mfL1X8F1k/3Fmyr/7Cj4BYLrzae5zjffZ
zWq8jO/911mN9Ga3bs2GU4CJB2ss7hba8dWENTBAZ40o93e4SQLhvR4XEDUx6fkC82PxWmcGS/G5
5d1WcxuucPUCA+5hXz1WQF9EJaVzGZoti4Nje+Or2qR8av3N1/0etXXKgf8wIu97p7l1a868Ee73
xzT4YsSYS6wgE2Q7KbhMsRPS27MZHObaI1xHkYEyemhUSvt2qkDTbYs+0z3auGpYpv0IJbAP0Tfj
/qvha/TS9g/O6jwNlYf4KV6r0RFQP3qFLwWQvuTO8yS4sm69R7VvGa0kArPmI85qEMS1wvsWaBHb
/+6Tq8eXvaWdu2AWpQojPRNp/s6mtUZvW4wVtX8VyiOpaYrjHTSFPU/f6xnndDGtGTULC3h4vf97
QPV3OfJ5puuYvuNc24tobGYLUwq4xjCoFdEZcFVhzPE0T4DsSH1QX7H9f0DpebkFMdFsLi2jnMTh
JtnQ1rdfT9GMdL4/KQ57VBqNdyKtYQkyCo4lsEPYfckpHaR94kz8M8ouhT0QqCmMOJVDaOFg/IvB
0BuOCpyjhjY6BedNb3nZJHe81e5vVyXvEJ9eduPkIf7sur0s7MB35BEvU2RP2Rctz1yfRIOTZMcf
FoIozmR0yOLzCAea303FLU+qEyQDSJlPeBbRZt/sCP5BURgmr2j2WaaAeuBBvkEniI8XaZkz7qAP
zWyTHzUh3ngqRTf/kmwqV6/42xr5ZX+/xXwUoSeTrUcckbZa1bi7aCC21JNRZjO6VtOeWuJIXy9i
tgSFHCYUIJsCbvCBf2164bTw2HIdmV10uG08M3I4fpvFES/xkBajixMOYkjnRE/c4cmlkpqYkIJV
kirPeWYP5KycY9+sjiH/zgtr2Pxz1o459gjfQA4iBGhbqbd4rjaf1h1D9jUBlgEvU2tkfoRe+bCo
Tv/8upTEv8KJgrJNLFlQ2RH6yx02N/O73HOBPTPxr0+jPhrAAElFpOXc0T3plHaYWEs9F07JycMS
E1jESozliBztXdok1ZbCgReYJ+l1MoDNYRyw8aPmD51nC3cyeC9HyVO/tuYpfw8tptfx7EzR22JD
7YU6tDGXYk6RT1EYJ361s4E/KRovkbtt7YGi/hX6p8BS6Eyg4pDbFe2+/NWYVJWugyBWQZLxOS0R
XvxC1+ufvh8TwxBIpvgCSDr8NraPuPGug62vBykb5GWFrwjGeA5AdOTLDahERPXMeYJ6j8ovFPVq
/9VSY+9IL4l8VO1uhuDxwu9RvB3OJA30+WLFyeSENSCSDtE3R2pwKHMDqu5s7/n2E9Jfe1t4Hj0U
stALF0lBmFU4SvFS4YieiADX0UUjBIRy2LGWlTSBxrn+HkqUiOAtFUxbS2UXbD+UKYjlmmoE8uGf
ZEys0HjZo2Gwn1u/8Jly3iiKCgqcqaw3QE2PEQBoEGMo6ENvZD46aMYaDP9RMp+lrlD15MGmI9EK
cWUE63FYyo3nBrjMIYSoV58RqG1uIcEnIAwh1D4DHP4raH2amg9//gu49fgK07GnBqCbYVJ/RYZo
PhMtcarmx2lw+HT1YLcU3aTph3LrpjZOf/GOQsQMCN2c2W5Tag+ugMt17blEEJd8G9EsEAijNx3m
e29XgkglYTTlogBZ1lN5IxxjJ7NYkkxvUW1D8+LjvMXM4N8ZeBNvDc4Faq0xMxLHBzYxg/J9HXIZ
quk6qSdtdkJ5FIZNybJHbkimb64Ej4DVDD5cdgEHXOsnqhSkhEBR/SqBdnHgSFLRagTR9aqzcZzv
g5fWJEhJHoeiADOHpTQr7p9n845EIlt8zPNbVr9B5IqdvqpiJG9ifrfDljNWZPs8vbBLiCNL0AUU
xXI3CxfHfcwingrNlAdsgVOLZ+2Af5H1T+vZItmywzUPJAwIXr/TSyBaPw9QbwVIjTEtklB3hjtH
rtFTF9W7G1md9yoSch5WAf1iYTYcHtG+lEp9yp2O0UAN1e3emXk7s56Y+fnVixqEMhFH3hR3Qi2D
Xr2CzU6tMt22pT5z9LihvdmKuIB5XTTMLRRjdOzDYjcKEeHDTYov1Vkup3Oh3TKFwNvR7T/NF7zq
jXi3QYHVWZX7hWcztCUst1z+2hEQyS0S2b6UQajZoM0R+dM1QbGsSkpga5AvD7bMQ+XujbsHu/X/
VREqfv5zm+UziWz2LrJ1rJREhxO5fF2iBX+ln77ffYCCziCg3NZ4Xlrvdj3uhCfz/HuzeeH9d+9S
x1/AjeHmLgh4b3liTzvKN9PtM9pZEwzHu9FZPJHsyp0TxR38hbatJboKS0LMoJeu9WjUjhmT1LXh
kTLMGg3Sf2gW0c0GyB7Zp44gYZmLWoE6R6ih/o5dTtkTleianiIKRsPkPncnRwiZT+jQbfObXxFo
rO/a8OZbJASN4OqSPCz3zj6/o5fSVMLC296c8JchaGuB82huZJ+VWbSPEzCXqopmA9p94V6XBXpX
2J1+py40DHaGFV3bgXUGuPhFJC33H78s2FN6ASHkNkyTU3B+KHXdC+3IN+2r/n4cZhAul/ZxuWLH
ybKZ49R0COAPFAHKPDddyV9xm2JirrePSFNz+kocfY8Syxff8hJkj9bERhipo9TsfMpHQNsrIxHq
RTAgW8NbrG6+HCYhzpmGv9hprhI9BsYUaDpewBQYNL2dF8OthdHwitsASM4ueYTALgH6v3PySW36
8QgMyxN2tvO+uum34MU+1CL8AyAxnAxkK/6BjCiyV40/IVENCXDHWYslz65wTuZoFPCwKN9XmapO
imNdkQdTuoCIFq6XvpO3w6wY8v5iRUXRsL3gNYJ67ysAMvMqL7JZ0IkFDlvESwTI+xBuGdArAY1B
ZmS+l48Ljtb8DqW/lpIb+3RQWlANJkEIFC92H+JRjDniEIL9w+fVyf2prAyqUxRJOTVOglEOEU33
vIzxUGGEhUHITiV43hAhBOCsH1jS9S0VMWK2WXhY9FdVH0LzRXUR9gVAeRTEhFQubHlkFCnSnAh+
FH3AakNjwyG6FzIX3j5TexWgU09wJYmN+ynF5eunTJ+DeJZPEj9av5zRPD6/liRTnYioUDdbx2CQ
iZ1v736cknut3N1T1VDgQ8OHpoL869jycq/fG1eaucoL1Urx5eawrQuHrwuIHaLJlwMPdGFIWoz2
6uR2JKl0JiOU+xFfb8GTcFqUG65+cHuo1x3Cy7VkNxOa3Yofykj77uCPoWW3NlKR7BjFIyAxB9cf
Tu2CzCMxRITG+VTfxIekrR1CQBW0O+Lnjl4kdB7rax3rNUdwbk3HOEl/0DVvUrcGZRqldqHPvW+3
yBe2nnfvXE+KXBG2U0NBb2hg7ldOpMGm0yJY+ze/a2FlOfvFYLj/xqdQfSeZ6GELcFOnbgflEHkP
Ef18ValU9PHsGUK2gP6ibzxAmgEnFOyEqxmw7XDqqpsYAEeEy9zF1QLv1WmUakPjOiNGnRWrwLrn
n3CEq+rof99capk+DOC1WPeair+owIH+OlHJAJz1jRdFH4hg9KHw7H+MeLHYQXsZs2JamGhDDWcl
kqBHH9crQjtMfnpMGPi11jyohm2WsANdqSq6GcxHc8TGOYGPik8RZiFj35ujY4Nif/0FpZTPpWeb
AQ2crAKFebfgKkrwZrGXwB4ZRGr2C02qAqudySOHQ1DM9vQPrvhggWP+JvzSJjZbV3Med3stJRvY
/+yl0KRHiqsJ/hVy3OeywOvmYm/j1CnWNp1dvA1YRfT6NHffDggoMZgO7mGuHqCTuD5DEGTQk7cX
3LGlYKpme/iDIDdmybAeKK08XEpSPpm0Fv0gvir8RKbVgyp6S+EpXAxO2Vtb7V7inr7dqTyaJpG3
P8/EH75Q6h3pU0C/pHgWEqdGYsPbxqEDuq5ut0ihpWsccGiA6T26Br/gTzWw8SQ4R5ZkW00hDcC/
wtceEF9OwcWHOjtlYYyeQfLLPTjtMsIYdzmGeyhYLK8ZqdxnzSKYxtZcwCbeKUhV2r7EnPiT830Y
4muAcMXsKZOXqxSeasv6kFjanYwaeT19VtrQ88uwxRxHLPvSaIMB4Zh2nQ60DvJoq4wDJzIy/TCx
nhXlg2gCwOZbI9Jseluu2RdMpYAUKdwil5TN5MnuSkXnP/7kA7fZ1D2N7H2PZib9ajJTgFn0dr6p
8Ven7iwExyqopO54N9aH6mYMPrzry21YfzsYTKFyjf2ErSJ28WXwItilZx1SLjqeUy/hKiKTZlTN
k24pevG4+Tii+j2wNS8zpF7tIQ+FegAzIAhldiCWRcUGfqJpkiblOanqUWR1m/Q7HTUnjXMLuxnQ
DLW0JJG9JihwvnE/Hr0kNy2yWqbrpG/xY8hyZ88HF3J5HH1fUwLHUn6wBQmjiSKRXK2uAGTFbP2g
4qGRbAQ4cZJxaiQM07y6Ek/RQzkGTNQAyYamTJ5J2/+zHLeTTCqnk9q9xcUsVBdz7Lq/01gOwUu7
Vg5QgfJpAGrn32LnuSymGG2p4c79hEPD/7lYmd5Pf8JPElbb40Yq8FqXcNKGCFxyKoBqXa3rTySV
dXKuAQ8papQPP/KAELiaCS6GR36byh96PVGh8ZavMA6oKPvrUDBuaTcXuf9AcrbgdO5lfyiygbFA
/I7xXqhZZEn/YtoTgGUOcGPueX9sl6a+tr7HmLCCmrBOLNS+FIfjCkcnFY1V2c85sLPkZvdTY8M1
cUff4gbdoELzIViB63X2WX3I80Qhwrgu5SeUaaAATIytwNPoaM1UJcfHC/oipMH8BrPJAc3b0eBd
XN5aa+/5ZUgLV65NNlxu3GjzMCTp1y6O6ggIrpKaBRmaXBNmNNlJjzh7OJJef+nnGU0KuQw3YbFl
75t5fFlnYUyc491PD2yblJnN8w+mynTiXLOv8FxfTQb5+r2NRgNML+tTtpc8iTCOECQ0XCD4Ifl+
ErlFUcp4jLJOY+Jydu0OYRnt6OmjheLRcTddpOY/Ofmvdvl2O0J4CKwAMPS476keIrO38/gllbXR
sD28hhWjR6rLCGDILY34RmDeeKs3WQX3CtB0KnTvXQbjc3pIaQ4rls5GXjmkvuvLKG+xvpKrZ1N5
ts0sWQlYMXkGUWLnGyM9UK1qm5Joy2roehLsSEDzjFQY08J8QUYvb0yyvWVXUshRk3rSqYEKdDzE
m+D+oYLmD5wITsL1XQN+q7nDZmzAjdqpw4x29Bv7QevEiE+k3oGKpJOxdnl+JtANSqKOLgsAqtmQ
3xIdvaiH+7YzHyUSzONSvsGntdQ6oAI49XryMWVD9DOI+HscAx24oDO8x7ub0s/8T7trsZkTIlLg
r/TlL7BSCeyQxMG4QZk9S96WAZ9LAUUG7eUl8Fzo69sAEN34CgvRN5cqR1EMAmqQU7waOdZC7OZV
Ns33SSFAsPrv0UC//jVsObi2ciH0/8Fy6er4NWMvnGp5DjZRPKxmrMFpvBi66SFG5vVkceds3V9g
HMOP044tqluF9XEm0Tru5BQy8CUp5WlsaNTJSqZi0qUuGA1VEwxfj4ecOMNE1do5ignOhp8Ve0U5
26jnTkQS2ctu9ZXMf0BC3M4NxUWnyCbSs2nwp4fMoQqgOq2f2CgHVUy89PmC0ekGIGGdLzDJ0qvH
H6IMf01Bi0x1A4PiLzbsk5TxwnN9f47Un2oKEdruTv7oZ638XyiYTLLHUGmZFUzDHxzn1jBpwWZP
3pFuOHmBhc0Qp94BMkidP2zy3oiTOLOmMNJ5SvTBlZIn37CAMEplsyDHhbWkyKtIDxVUGeosOboh
8HBRahUJA+UpPhiF1Mr5pg+U+FeEcVr0POPyIi4lmyhtxkhfpRTwn68hFBx32QColHjQl+FgqcHJ
CNAhGIhCQCjj6RIGCVZDntK6AJ4SdrbHNLMLcKgqs0p+/+lSWrQ4CSG4r39QTpm/j9pHKuhygHkc
DK/9mHI/2IK/PC2JbkTPejE3Nw3vYWNdzHMgs2/Xbgin++mTEXAkn+e0Edd/HVK6azKYekGRNT42
Fb2B6VuW6kYuVyCejdYqmgL1/fwobNW/vPMEY3voaMQHeA+vHeWfnSo2VeSnT3yC+4jjj6EwK+LH
4XIP2XIz+4tLcoBeiuiTIwSsnFP5dViolwcFfj16XFpVqQEf1zaJIErP09xcVGRQVaQgn5MZpi19
uNtnuPTBDcJQRkykICpm0g5fKLXivtpRN6bdO5fgSybC0zm/DPwbLgTPrcnx/dAsdd69T+Bpq04M
rhbhdxLp0w6sAEkbFXrCzcYAkgglaQ9GWuR9AvgluyN7BRgeGycAV5h8NhW8jDAML927HRD8ZTF8
FB9RbkqlcA3NcpEL1nKwTIj25F/DAkDQ6GINcEm4Nt5Tzuea2Xdkj5LUm+sA/Hsb2BqnFHL/oPvQ
fsYaC6nV3qqWBZxs6RwpQTl8cN2uUVZmDlhStK39jorZSgsvJU6sfpN093oEnEpv6Y05js/AdrLk
Bf/QGdPCgQjySn3X8RjugV5EEGoDkKLV7vjgvQ8Wvt8TsLRmtQ1k/JH0CU1ZsMG4a5CaKytFUupQ
7fbJrQvQB2jBVKEsrB+lF8QtWI4HpfQn7c0CCii0QcXIMDEo+5OasIkq82sWWaPYKE2SeQadaj9L
kuKfrI9kDCKRIH03qFCBYxi6VpVNGD/EbPSPvjA0ed5QWUIRrVg8Iwn/1d4ZzC+OWbjcLyWJLNTx
PzWRBzH0yfCnt0n68wmv+trKelzb0XynFmd1wJiswLXgExbK27xROE51H3JoRTaVh4sessDrAfzi
XfgKiBU5NZQiveh5mujl+F/IANvwJ/aEgabOY5DKGJa03RS+LJLio0eyv2ABX4G+QUgd1TKwRNXN
IiTGCmdFOY4bAWqglGy9PoE/iA6uIdPTcplRkOSAGvq8AU+tTYmPmfKb57j7R3gVq6zvsV0Kwph/
X+uaz28gDCHaOnajN/3pUgIjhsYB0kKBMXqSaoAnl6tuw2YiApp8Vf2k3VsWiValjXl0Iabjb0Cu
LOB+yVl7J7WsxEZgnJbW97EX66G8gDfqL9PNPQRA7hEUPm069gAmqreA5e7s04F+WWFolEfKlsX3
Ffix+kPrMHw7unJ1qUytzmTrzCYMDfbUjlpBDqLfp5J8pVK19WnAqNM1OYHYJinSDbyewdqMj7zh
MqGSaTizWkN+KG+qaO9SAP1tP6vAlD5DQ8QiBMYFUTOHPmifeGaUUep058l1WTL15wNfWN/Dhbt/
OqgWsm9ESzIbZRRrn51c0GJR7ip3yj86SC3cWESCu1I8f90jilF2XFJim/a9RQwTijzTu3yZS3a0
wj4QDiXa7JyXzVWm2JvcNXVXyk35w+PmgXgd6FYDSJN8W9bLypqHrk8G/SAbArbkI+HmH3ItusaR
jHAutX0FghMlzgdpXyQdOHj1Tuv12oC30RFT73fSnAfDSLYJoxE2uP8CFtdE14wl6nMdTOfQInV/
PREUuZ2ygk2M3WOu8s1KdUR3OheynJglH+s/8xaHFcnNLefSAsEiDCUwGjlsieMTjkx5MYySrXSa
a49rwfM6TMUNU0r4e0Cm8Mi5qTnUPfPEX8pbZPCnfJmYiGLj6czcX6HwWw34VMojpPd27GSyQoz5
YHN0HaiL6RxUaAKA320hok6PIFJPZPKCDVaQ4L+nDl3iYb8wkOfySKy9WnHAL+G9WErJmq9NWnA+
60459pUZOoDvGxY9Mpx6w0fC/zp05vz8eRWt51Q24SHcFOz37yN92MmjjyDsKXkfkaUdAXl6rgXE
40aMQ2nKyTJbATqO86nqXDDbLw5Hl4fQV96NQ32tRxHLSrwCrHM/TwdlBV0Z0OBpYCYgXpJ58Tay
3pi0+duCZrl+JAUy28KhIEGnzDnGWyHrdp8qIgN1wtAEFx4Q89SW1Dg+vAeVMtRGpZSC4CGHQf3X
vnPf/pmsb7HoRc0/xtGkVDrwQSI+NKmOM8QyieXsHEZdCB3pnIzxXRHq+ex71xayVgS14Tf+BqwP
K7SzUpVRP6o4iCDj6pwp8XZQE0XJdI59Uq7DXBGQoBzL9UzdUXWER9bjop2oJs0oci4tJoIFZ724
/6kmtTb6py58NJFFl9G8RsqfgZSYTTqtpSncXLL6v/9I5SjzfSzqhqmUcFrpL34Wvs9Pehbj5Jie
dDSxYUKb6sdrfR2Fibs5Ae+RFUlQ6TJnmilTIkUsWRuwI2SvKWHLxP/2VVWEfWGNN0Eof2EY3INp
A5Q51SOulzCOpzyjtOt22WaITfW6yRNOb23f8c8oV97Re90EZE6AFqYCRfq016Ufs0xaT/B3fqHb
1KGiOLQyot0AJP6xf3Zr2EBgxPi8pCO5anRaFoOPplH8xZ0AiTZ0+HMr9isfb2uuJCmzQjcZ5hJI
ZBHO4oioWo9CsB7PG76fhLFe2/AxJAPejqAsCRdLSlmo8Y7u+N6yTPFdgROQT1jZEa5bl9HDPxeP
vA5s7f/pSy42krOmElIUYdJCqg1bgUVeNV+AHsgWbc+tbyUKqKT+G9nhPZif6fdytUbwgwHQKKHQ
Y4fVlmysCJu22Ve93m62Jd5kXUdVORwfmJYhKDZ082OHjJKCSabo1NQZ55GUG3M2snvwdbk7c7yb
oI6Uv3inzKH+iwPIZLiJdFxNqvKueln8hFkfgxArJe8pfbnHnoaCvAoK2FrXTOtR4jV5cuwAXxYT
zn8/KbcKrEgYWfulZH8hY3NULigWdmYN+KihggBAbM7Py2kQ8X9JmtGdVHyJ9GnIRtEPJi/cTZYy
y9+8c1qYPSUoUhTW8weIWFHog/HAJF+6md2ZgTBy3pKJm4qSUn0AgOlTMMfgCTBICcAN11hy0CPr
2Yf7zMWPggYt9XekJBueqUGgb/pl+AHeL7Gf6ge0ddpS3CocL+cMJqEGJoj1BRXMY6q6WAGcT/PV
T3se/EoLM2hacaoLdF1atn0wJ1/vAySfbOCY4xSLxJYdyP4CtHEqSMniY/mFHUveGLB0DFntT513
CW4tyiXue/LAQD2KrLK7B7ssl1e/yxN6WheELKOBwKqnlOE+DjNzX+7xn+1yfj+9dChN08uE9OJ/
Vh9Z41Lop+TpQHUs1hYd7uG1KWHyv2Fb3eq1zBdSHxVRyx3O9TM6EWzIMWOMQiRfpIcyMI8D6BHO
dBkz22NKBZgec8hcE7zK2tArxvjlX43fRnQ7wCjF9oXQ/6l9JmayrradPIup1yD1smeVurIgg3dY
ucP9lKdH6AMt0Dr7+26N/2Uxgq5+QsTzKmxYEF/SmtDRYHNhtc3LCbVduviHiLj4gAwF0yhXegG3
znUpkYZjYnn0tSzMmB+xoH9J6XI4wR9IWD9DX8AyMotFP42Y6yY3QihWKouTi9Omd7DrVd+hfv1z
5LcA1xncuxdkbC5x5QqSmqjxmKtKGALQLM2n18TlZH7imx0WhKSOHsMrQffAyJX7Q8oGy3fgATit
y381k54aYYnPv5QGSsow4+HgpcnA1+BR2BjHs7RNq6qFh58QCImHAWx1jn7OaWkOeLFrpG6ZXJAc
jIPWn13m7yJ6xPOeNjhz0WCWE4GjZthudgfdw5ooPwy9F4I++4qYmSgwgoHt8IPnyWbZbeGD0hnk
L5eqQn9AmebbTN5j4LyLKfzFw+hB82T7a9BMt2BpHBiqmTMnAV3mDPaqV+ojclH84KpCmZCPV5TA
vwu6lp80iXl/2Nn2ic0KEml3G+zILJaOnPlNTJzXVNMeIuKpSl2sZV4w27+Zmd18xOn+OWKID23z
OgAvN9dDknvo9AllQzQzNUPGp1ceLvTBIAWEvCosWE4mO4arL0wjJjFrSVf+eFPE/eYiqhCt0Hh0
aD2mWAao4ijfypFSsWdUruBopHQrAfR7thDpXCd4gxfuWUk9D9ajjBuH0rNUYDSHtElzoewQLruf
+qmhNvZKasghjAGHjkuyhQWXMIlzaLD1d1KUMgCW3yXfFFtE3fifCcMzsGdbBi4EV0fOW8H9wBg2
4J2dDIbiVQ/s8EzRz8jMK0dhcsDgrkXlFmIsRqDZr61yttff82GwTSpguF8g+a+4vqNgQVN9+W7/
XT8LTaLxo+SWK8zos0D9ZxaJO2nCFjgCNG1qufEFJdCaLX/WSYFWTRs8v+vq7kr9mDg8+RMmAraj
QTpuy5onwjCBZUQMljdkdBA/x0p+QKZzcBZvLIonR7dM2FglvweAKRFlOieMNXH3tSn7l/+dL/I2
/0KqcljH0ulJnbr7djEER8nNYL13ojcyW1Wp4veheDmUgokPbQYelpgHgpmZMqNH4ory1JOmSVL7
XjZNHWLQ4yOYvVB5KEINin/GiL0qsoC8p8lDqvG61f0Wasl2cby3Xu1Lx9hG9Typ4dqLZeK0UCnG
heCooPv8pwOMug37RVISAdiE2Rk2857m/aS+5IElln9RDZx7iSYbdNZ84Qh2moIKRYF6mPV0fka5
zUNt+LbysTDBnrk4AZpKDl4zknbQCrGY1d46aOA/LyrTuRk9YxlxEO7+xulP3N4JUpH1BwXvr3oX
P8Ex03DGjCJoUlmeY3qDcZb3j5D+XB2LIN17Jz2aDB78njGDIBoxnLRDnco+XVBLv4nNpn1gzQbq
uuaLF3DIA3WNVJsstO4lgAUTw8+JdBGbMXRfz6extzS6ChRm8dV2JFNpMVFQteybETbPdlB18e3/
78ro9vgo8P5cKRjIZAS1h1scCnwhE1NZLQJDtSkvFqfz6z772tlvhBnn3sZZUnEjK90oQK8COYSd
ZBAtALtGA1ROctDe9Z1K/fwQTBAZUOikj6F5fRd5vny7cY0+Wd9ucyHgConZ5tu4i7OjYlMSIfDU
EIh0LOuY5gqqQkhVXU3BZz5pKVsq9gyokN13pzNc7McsE8846KrN0FuQW3NFbHoatTGORCs6xYvd
G2ileDbfUmfRx7hicK3lYgdZNY6VpgsOakzx5CrOFN4PLukytC+oQL0UXlRxbfUxK9qBg0t82olp
8MYWwe2LTUddFNzN04juOk1rWzquASnQfSm76UZTA8nH3uUL5UNbx7yoVhuzy8YoNWVXZsLYZwjq
sT/BNz279djzW82R1PpAUVR00Tt62lNf5kDwNJcgfCWFEwDk1WgAO2BUBrhhzmgEeFx5WYqS4Zhc
ZxhXieVJC2NKDqbQtMCoQIcBljuZaARFSOQWhnMOzgZ1EUQaHexzZ2gtG/c5PpnChVvMimyAXr05
qdnLnbJ8vgIrapAT+7g/aYIUm75ju7ZeVQrLo4uDpVzd1H338gW526SFeEbU/BGjwm4bGxMz4DB0
ehmndqS5i7Tj8DlqGLuohCgbEYXdnoKNjNhqGbRaTyZnLvCM4xu+PHdK8yIw4zynQA6+92LkWmQK
oH41GWu2e5Q7F63xKHLHiiZSiX2fTPQKmoARvUu3cVXt8NFrlqI13PF2DYQnKfwCqFiyjf3ZgXZt
myXun85nCDELlzQfyqBFKoeLSP4LgfTy4zMqcQqfRiRXFg38BkSR8X3Bck5QfRMaTulY3EfeRFTc
Ol5F679LaAr/3zWLrm6jsBSFlfSaTR9YuNa09QOZKgRWSQ49YmOwXYgDQhNp5hsonxFtMSworCs+
YdD8JLLCqaIg3joOZCvV1gEo6Z6VgWfIfbdHTkj8icRG9RQB1iJWQG1DqzeIEFRNW9m1JlEYSxYo
xuPEBP3XrN+ws9FUW75jM9Vks124tajYqHC8XpxoQ+uj9PC6UPnNyMcoBvEXEUqp3QYoszMYvGYn
lmjcAmSY4ATotCBMWnsn5QukQH8+w5ITyfBx6OyXVGUz3mZOCYlHBdbJUaZuVc3krHFRHmr33cLb
M71wCooY4RIk70HaJYzzWgXRcevhE/KqBPZB6QDYe1ZPOC9Juf7Asepw1IXNTfgx/W9y64Je3Ox4
uZFsPpK9mDlpN9Pjzb+wz7bT+RSJM/wotzU2UiTtuP9A3rjpekLgm+tpZsxIofdK/qiF3qvJNtwq
ebeC3JUAM9If9dPlWukrZGehzRdk9+LbKaMTAWQH5ox1tG09OmKckKHGoPIB97ISR18PfJYaW/rp
c4C+43Yr3VjPREfQi7ZJmuhHqUDNvnAgyO+XZVKqTIX+RfiMN+ZnIzR/+0ctxyRZ8q/oyJYaBwJD
U1Qx+DLkqOj2qZnIJw+t3w/esb0gT4w3+39JhzjxxOUvljT4IWKz1jJLr1arDQFcKooS/Feb9VY/
aT1xpLjPjvAmPrLVr4icng308uI0lCvsAIz7h3jdgSey7UBUZl5lN9W9pr/gLhXZ4POeAC2/Uyf1
Gkj31zAk3diXJI0WnahGucsc9N8UlRjXCYOOCuuePclNtdRqY4sYE+vtnR56FfUkUudxYgpYlUVC
tzGvf9grY8V3vMWILG9kgyB7ID9iGkP00TPWtlBHGkUGySRl3SsXu2BT4QeiJjUmnfXVWO7BOqgv
jHOrWsrQV2wtxv+ci21jMW2ImZdLYWMTPcvmvSfZkBPCcqc1pge5mOvPJc9Nj+fhWCs+FX76koXi
OTyuwHkc4j4f0CxTXcQUyLXU71M34kJKTRdI9Ft+fyYIjefxx9MPu++CdumStFMZ2X10EWr5JfQ4
7BIKT7NSFsJOgNWfd6PtrLwNsjiPNXsyLTHoBJuezGdgUCNMZxMwN75hemffVng7LNKc5WYq/gNL
JXg72WnL+ae0r1chC5NiqxdD06IFkiZ1G87Hdy6xYphfcfhQ53xjI11z6GHssodmtXUiJq+BfbpN
wc7CaKcsSMOsRbNqoiCtsLU3m+FoXXkdj8dvBNXx2LCvnxJYfM4167p+cLYZZ81ubfFIFE2QCL72
XQtjwdHcQwleAV19ofeo24ZHg8vzs+22t6uAIvgz5jfP1nKOvxy1wYftXTAeJ4S7hT/go10ztPwc
q/le45DlQu/T9YUp8FytnHDBV5aTwDHdS5bjDFcnu4jytR/bBA972a/ilbgcpp0hD5cuZvwcDAjJ
V2JjrP8G2HWX4sEL93vebVtD50RhxDaeFgznDnFO/1NuOvKb4ZCzmdTa2xIRBJ/uMaYp7gpkf76f
kHMWOU+qLb6MrstzGyMgC9ZHSqMbvgU5dj+YGiYERDWdOFvjTRoo0Sj+xgVCt/dYTTuBcAvGv21Q
MJT19sKUfY2V+BrHkrK4+SS36Xf/mNqDntOkYwp070iy6oRMnhkD2kzAfmiC/BT2OhTtkGAv1cdP
cRQ6R3rmIdrnzZ25S4+wNWKytDbgP9Dvy9ghPgOi+V/Nkc7LTSSfZ4BeWawGRySQhLMna3DGLAIR
g69H8bSN1L5DdppFCJb8jm4WeYPC3u9QR13eMu7iuLVifmlqjLC2tLgAUhWpcy55FWeNr5H5QufN
Eqmi4cCxPm4PrxMmboDvyFMU3pGpOPc4TItt+qJAyVItottz0riieCF0bFS4lAbtccDPghtn36Q6
Zh50JHOBwH+AcBxHqeTeUp5/aN7t6seA/y6ss8B8ejonzrE/lYlK3xiYV1XXrgRBlAUzFzdVsGHO
io2Krjex18YrXGj5XoVZIx7bbX5aKpglkEPjcL4oZPNpLsmOWQaSZ0FvkiyMbJWekVw+/QPuVbqy
o7x+xFDZIPmZicL47VaKOvXSIUsR+bkbFo5NEl9VScSW3qYAAfrnHD03ipD69FMR/TowtOppJnxB
YAzk41ABbW1kjTIIcU8NuA0zmhimkXGykGVP0DZaTnTAWr8K/mXumb41jxa/yn9toHDoOCADou3d
DAUoCxGD5PNVormqQ0qVYa3f91+YqiCsRkWAqcJJARiTlyiZR7BVcpfXqyzj2O+TmUwR1erwV2DL
QxW7gk9n4VVkd3ZBCBCjHknC4/JYI2+sUUaArWarEizpvLv7BuvJSvL+on8PYjhb67gsHhelyPCE
8gA89Ihie1JwNuRqS8IAhNAnaMT+f8sGzF6rD3vKsop+V46jU7HyNkLlYQu4KIuWsGMEv1JP5j3X
+nLt1ml8IGWsu/sdim7DBF7H5e1afch5mVf+3qhfrwdXXzWaBnSZ0J7V0L9Em/HqYgPnBJvZNYQO
WM+N3wmIsbsRKibvDtJNknqrSXPV6i6yGGTnz3jMgLwOqVbG+I1JFSQWkPQB2L1yxF94myIfHqJF
btFhoiRV/uDlXSBwwTWEl0QmOuZs3UkOjsfCtdMElWE+SlBzAUMJR4TSaaqiDkxYi6Yy5p5Ne/FU
grK8C7sc5FATlxZVOsmvYK605+rup7KN+jG5e4l+1L8IQNvyh8mFziHOS90CZxB77v2lxR0blyPt
v4G77X7SuEKtA0OYFuw1sEjMTKEArfCFoHktj8knmc8umpL5NFZFVicFSlRT+L/TLD3GNC9p1XlL
++fsVumf08/w+HveOq5161dxD08FsCMwjaaw1I5nxv2beebf64YQUL9AnY6i3uShZBL9Bagy0NWP
1bFpGieykxPWL+lhgF1aDfBEFH6i8eTg0Ue446Cbp6JY/RDI5EZi24yMziv6pSSHNyWCgonoVYU4
udvPFpIQ38+X1o9g0VW5zn1u8jSEiSjqMZtyCyQ3R3MVLr45cQm0O3bgB2L6lyO9scUlNWCyKtFl
NTe6nSfN4y1b1po1WHdsTd4adaPBupl8TpIJBo1+gYH6W4M2IZ2q3RnGDYilDnJ3vmDynAzUnmoG
3ztYqdg4jEPiFltUMtSIoDC0fgUFBdHku/WeVXvHFafZgoaEByp/lY8O+8pwhfp+RWm4cDXzq9NR
RRCOV+vGK8XtWtaK1uZeZwICdNFCzQ2gHsi5wXi0rAWinyQp3cuFJOgpjf8yymsY5xbjexM2/Raz
4ALiiJzv8yjjb1B2LZeMj4SLyOZgiVy9UukaiIgtH1sQkf2bJHIChdVivdJeXYvFqb/IxXB4fsZL
jmnXI8BgQR2Q3pHENY03qzmC/w7vLM/IuI8L4PqazhWh647DSPpILrpGTrWzBZ2wwPGfakKPs5HS
NBqoGOGyGQbwpPqZ+RgsFxSwJKW4GDUJrxZOY/Qw0Z/fqF0zu+bVf0CfDH3rYLvu5Oh9IOcqVgpS
0txhT5Ulg4yCVScUnyJBEKDFZujpQR1iXfSNJZ+cdUZDryGZhdoVGRhYBzDtIMq9yLNmB7VmoUzF
7xCB/4mLtEp16cS7VWJz85DIZHXnQwSJVfMwdxiXdVGJaaqj3iC7z/9x6RId+gLFyUNfU/vRcHqc
v1qlM0NnStXKRvjphMrLRZXgcC3kG2iJaW5DbaB/h872nLG4kGhV5/xhLCGcxQp/rHnqKxFDPeR3
YA6/jeUtHGDBLFKYoBcToG/4xDFsrHSGAqT6svomKPRlYCJqrWomeh9x1p/gtd57FD8hG6e/NEuE
bfm61eDdui2ZgnVGo7o0mlqkbFXVwmWaSOfc01vlPT8RkwcPyBJ3SY7iLtSIJ4yVUk+MPfP7Rrno
Urm4BsP7Usu4NTacJMCFQhBR5FCki6Jn6LXJ/x0ayxc6PldcGle7svc/teeD3AFWxwtLPTf3vd+X
vS/gCIHPA01V3cipI6OxSTHcWFUzBENISjT/m5wW9AMKqCGoJyhJKUpadJr8NwDwcMPD2o3iJu9F
02FVA/D9r9Vdg/78uaBYVFYi+W9u5Pd7Jfl8vpKN+bJstUklVHwLz7DbZcgYjdHUiynT154mzq7r
vVMPJqNEBGgV5eWF0huZVHyKHUr/jjljbNS9BmfeQaXT5JpMzJ4/mggbYozO89IIzOhY6ECoPiGD
wXLabUDiRQAimO3npMQhYiT48iATQ71eTEw8eN0LQrSZ7cNzvsW0M92OnsbTket5hWg82tYC8cxe
f+Vtu/+zNK8V6pPdZ5n+Ngze5JCLLxK0yyNhtX2HMWcfOgkpgKOz9hqqO+ORqwivNlmZVQmiBYYZ
FEm/192MaIcVnMaOHdol3uY9/c/dSAyPlpwO3DWnD/O9uUV2chER0ldoVZ4MeeUFfwKFGqJL1Izk
hB2bdbE6scaiLcbY6CyeuS0gNSSwiOUoCu/G2cnnmuRxGWwgYH78iksxGHx/xOImL5NcNh/AEuQw
MJVu/dJzJStEQ7w7AZJL+3UOvb3tiX0B3J8Y8BljgNe0W3G6gQVUFljvZLSTS6mYQfOXfDgwA2Ew
BUOykmJh6BA94pJhyEHPgTW6x/WRI4EXiKGjzqyPJ4Wmv2FkCYhw4ERW+P+5nWLeX9+jIHnVuYuM
gtswlswgsAkcKur+3kbZpHk1G6TEC3zzgwCKXRYsJVYq0tM8q15yTF+LuFKrLHERd9ZgbMqyM9Fv
GfV042D2k71PREy8CnGIz05NlESnmvDdqbqBNrrGJtnLGxGB9WHEHqzYhxZMgtHdhp/WZcicw0Oz
cz+J2q9mTNiY2pPAZgarAymwgzvPMSPIbxtE2/1kF3vnPwi3ssy4y1jujRtKMixkw/FLa++AdI2q
ivJ+O8TkHtm4vNfKJpxC73Fqhcjdk1///XHOTkMi/R4/uZsoOu/rHqkzenLYL4cMGCka+TkyE1PX
INpY8Y53FaPd4lF/wk2/RH5HHg3d1v+JzrKcYINamCzwX4MxUSfvs26YJaIKBzM/Z3lt9EC68Hnz
NdQ79YX9vu6+KB/WvMx2AZ9RPrxrpVxBu8JNaVKX3lj7x2aAbMYXZsnJfinQ1VGe47eRRN7+dVx8
OpfKt2eXZJSfM9mgK5s5VEzz6INF9Jc1Jty+ozQ+TQ5iiaM1DHX/qsAL2aGafA9z4cAjHZsrZi1u
395o5xX2vLBeg5rH+EXZ9UONJfDfZG7jEjNCikO03t2ZkMK8GYoDDoSy/1i3qw8fwEWH5gvtm//d
oMT4oue2osIJLIE1tkXYMPtjhqszagDVpLSQsgWAdmRGrISh65pyGvDx9jDWpHXG64+2sGX8QHLZ
u8/7sNXFIIhHqU7ymOCkWioErm1BlpAdSNLOW25k5G5Nc4XxzPrKY+n50Od0aM9Z7vi2MSYHG41Z
LSkqA4aniC/E3oUOufQVEI/YY8Kx0nAgm+SBMX1rJsidE9Yg6wMnSj0Ooi3oNqskNr2Itslz9Kf6
Kd8qsR0lyU2UrlDxat03cl/YhnzFhCvR641YMRbCoaGUbRLsQL89J/ul0M26em36mxDooMtizzib
trcB1Q4cBN/jtq2qBXGPq4/9UpCg3uMgUs4zGOxRF3fPp651ZioHR3ELWcAC7joyUZL3QxVEyVC7
yo8gC3FePOhGw00Fzbn5MI0ev+6QZi+r7/X9gRk73BA7XwnmXmL4lMWyb+z1Ltw0Gi/ULcXcwwGG
rv9edc2Tuc/YLrcGfpH7AkVGRfQnJktPrNtSIwZQhAdFJ7ByxK3HBhE6BjmliHwToM71JLGfpv2t
iCCPJIctX8hjkS1osrfa08gNiX05r5o9Xk/KdHSyegWjAaAyjya7ZaYwbsR3na5G7Zg6tXUP9llt
1x68lLUflbkyrAj62zCBNh9M8ajhebhgLty5INtOtLmZbEKDVHwVz+HOcKJOU4/0N6qjf4VBACrX
4/d8VWO6wMXHkl/ugPvU9EtbPp19aRiX0JLjTaRa8Jhfetqp2F7KQgrNXZuGzJONURcz6GqJTMAb
drIiIrApS1myjM/5oXn8fnJZ8ASdBt/E3HQUvACyMxOyQ7zqQEvQx61hRPAcDNfwAAU7C51kMC/P
xxkCSZVX7OrzIql0+/mPAEFLvItgZavg/GGI/WI/KWoeJXhtMGl+mx8AIaP9JGbd5lH4p/MvBiLU
mMSf4cxaMkAkl+tFtZu09R4SeVjjSG48L7pL6In0YCjz2eeuooDrVZLCnfLlQ8NqruePpEAMHZDN
5NNAAb37A/c6VPca3FY12IUZE27llJGhICc3zbwfWujMsSlt6OQQVm0I+5jzz2GAyBo83VmPvKXo
HGVskJP2c0Cr6Ob8tTu4QS+SucOAia2xj5sYluqi93U7Sv9ajhz4BK27iIwHylg6X6PRmzmeq8s9
C8EjmQqu3jdjEPpY6p8tz2ufklDdoelTGvUOHJAuLbvjEwRZxQ+Z1K+SPXmfzacPql3muRigSLtn
LgaN2YVMh8NRbQRPhXuSvGgUmeZdNhiqTqiiAZoWh2cnW1mo6pWMrrqAELGAH6uSSm4h/R8VURKY
XJ6ut8IzHCkuoq4LGk1VgW1+exOtRXZRDMGvQYM7uJQy+VOlrLsXMa/J9BN38uCC4XK3T2lX4zPe
dOmK+UUE4xsHVzM10GEBvfWlTCnF80OKepM//7tCqSDFNO6Y9fE4P5Sn8Vy9WvPUYxCq6mtEXZVi
Y0fezhvvxqSbjjmXevm2gjxzqb4Gy9u6tXh0wQL383ly/4TqFZokvCyYb89nUx4alwhe9XBsWg7/
IFvCQp1frsoznqurVQpC1aC4v+FakSkSx71qX2jwVl7caziGHIo1mkS4L0prZ1MEGQLs+SgEWdzY
d7WLPQTMEVB2vXoOUHWRyTl9n6+gAysJoUJrgFxmILEG9UpsuIXxeF8o1Y0NPUVVtkYAIit3R97/
/oVgV5RkjgA9dY7pL/1nl1meh4UVO4ckvhS6/zZ7O1JVKZFR9UCL9nF1yN5ezcKzkJCoPw0XiRG4
6IEKxo4RStJofvzvhZPSP3QUCMwoy9CSGkGE7zJrdbTAQ5gIF53FI0yZRB5hOWu3VUp+HUgrGwv3
kels8B6ickCJNrkyyunpvyKB6RqvA/KF+PicJo5TohJAOCouENPSLGhS2OnnyGEc97Ce+PGkUqbs
L9XKD9HEAsAADRQ6zWgCnDNzCREg93TwTKfLpR6jSZCUT3ap5UjzqH7FJrsbZqHTFtpYWCSzD7gl
QXPZ3hl+rQzfXtxyqzzvM+r+lTqvdPRw01wJgyyC7/+HUHEXxrh33iZiNRtcyznDKQl2PU8htBNm
Yh0GtAz5X5PE0qPDBabMQ5r5KDUgJOYAZOCYGPpvszerKk0NKezmUWzs+/0Ov0uYwwK3/Ls2ehVK
SXXI/jrEj8FsqhpefN/CRnFw68c3MjrwUM1p/xnq0VyLpj6tPK9BaQ5G3DrgklnCVUOEUiV6DIjZ
FmuHvh13idBmk+gNnVq+VHIch8x0s87ujYrziRJ9gU0TKDTRJApHYr0WOiq3IhEo+eXawuJk6igx
AVwUb1OU3ZoxQbIfvjX43XYO+G4dT9QrfjPykFstxEUrIF9rYRVZYB15WEZpHk3aoJ3wkAQx+gAD
v/xy4HMzHUw7NPHxFolxPBrrLA3Pb4rTBBmN67hD7PF6oUZC6rmz7dYN7SBCr2tQcizU/mZ4i5Jt
CSutM9dT08ST7WVkBL7sYZJ2ASZ7jSAPGJo6Mrzz8MaBrMw0Hzf+CpuSdvFoSEiXIT0zerz0T7ep
pLM8Vkw6GSnbMCS82J5rdNIqsClAMUMeY1zXCyze7QbIWi99AkeMPL7pJFcYHEiWFPgLiXiyG+Bc
sCnW6SwhLELvBiegJHrNMvGrfyzRZX/ZFSb3AFbvxFs2mo+9T1JUkvS9EfWDOBKMbvQcVoMwhBYB
3qxsIaVJFvE4d9MtPsqrXk6XFO5U9QKF52kOspxykQ5ufXldFObc3XhUxETMUtHZKO4M+UURyOBG
+9clppsZf7RKDjQL49vqYfUAJLYHFcaVUTd2TGMY6+yDjT/wQ6oGz7JD3YE5bXROSc061B/Dy0aa
iGjas5MKvC1m94tYQ4QOXV/P+SLBg+TXi/dAnYVWutQShg4aaYW6debRy/eU+TYVpudViNPF7Sbt
6TbR/KZdaAGZr2fr78rxuLQleJ7CQbV1QTRocNyCJEOdcoorlVRUCsKL3ANHzVTYcdxpphiGumOm
Z2/dhrvtmjKHnQm86Xw76aw9UiZKGN9jHTAkwnF6aXLHS9vaxTDxKlKkhLkg7IGBcUFI3xhIa9q0
VEkYaoBT1W8uAoxi4pCf/q9rGPOC7I6HGtjbUzlBFa0eyf2uua0RdQqpnVpIYUMjEkpqpJLm4od9
01VqsidhVwTrug2OC8IyR7E+PjRYa+mO9FsK1UhzikD4Y4TnDL8ymi6ZuTMkxXybzEmpOjt3s5LW
Ouit/luJM0Q9PqJNuki5hMKOGM7ng/71m3G/odNGtFrtbhXcIvQFCPDrw7n6H2jVD1F2HMg75O8l
LlikmdWQR+Ua0M2h7+8om/56WjafeGNRobf53pAjUt1c/Urn6+cD7jQUzP9pm5QomCOhpHrYixtk
YQd1mmfntf+JrobeVTcbGRxdkB0lvXJ62wf7jIrfiP5aZneBUeGzDAmmeT+hH2vwG4yq2+IM8gGv
NLRgtQKnO+/ps9RfR4tEaZz0SmSqFheXJsXnXOz9NRNlAE69W0UIRUPN771ZA7wCu3g2+e2ZzxVY
d5IAnig2u7izJbm51Dn4RqiiTXn+1WJrNmf8efgHZi9X0GtZ9TYzqY6R++wDjXmPgaNZS9sNis5M
v5ppXphte/CkBIFyXoU2RBVG0qa+MLBB5iZaHMK/OHoaoRAElREM/qK88GSpzO10BgzzEf4lupop
M5GYlTTxTBBauzhxZNrKma+I2MDeVseP7oN9uOQ8g2HkE3HOqJh06OJyk2O2JZx6Xza16eYvruqQ
M8jlo7hSYWSgExm5yie36BIlUky9vQGDOzLTZ/md/6mspW6CAF30SISmKyJboN9n1X+OEm7Ytymc
2R08kcE76u64/ISaXU8IYdu9wQrPTnaeuf6M3dA+4KHRiTW0V1PTJFR/Zea7HGGO+cDy292VSnxv
JmIZ0ISLeiSC9TFOgb/M18E4mUMPrAO3sscPHC0jmfa4zac5+afWJaKYQ3mMiw0HSyjGfwxAY3hg
EXHXif+xVtP9TNfcKPJ4IKnyG04SnWxSnezcod+JKF2wzafdyo0X+RL7S77gRXk0GRqOXILFYNM3
Yv1DTg6x+ysrSRlXMwx5Np++1UkD6gGHFmTsERX+M5f8JiZp1l8C0GlksfsjHAPi1bUeioX0kFK6
0Nap9mykp12mOjes8p4miGQb86NkvwEoZ9gQk523DjnBMWTMmi5KS21yb2qgr+bQheicHNYLWSpW
R3Y/cY3k0qmlQBbItODEZcZ4NDZ7k/ZmMPWJ9qmZ/Lh/HLsUBG8jdo6qHvGFDNopEaUvNt+s3+SQ
9R4Vk17oam88ozaKoECXXQ2GdXUCPtOr+8Za1gbu7PZh1CCLFTqdVe0OyOPV+DgyU36XHIwhKNG6
LEaoiv3K5qFoRxboHnQrP7fwvDrBnBOjutalLNmSOxkkGw2HbtYPgAO9ZcvEJ6uFhD4p+vTG+C+l
zs2yADhxPwN/biVIYCHUbMM3L+4iUVUZaCE9lmarajW4kD3SELbqkTMmJAbGqRvLpbci3oVYye3J
kJSS7uBupgKvCG7ZzfaT//R7FqHEmhltDMWCM+9mJy48fQZC6a70l84JHWayRbD2NerpguSsGTMN
LVo9uF2aUdFof8ToahbD5NWlqE6mxGeW+ZqoH9lgO6EXmFqmbfbYvdPBZeXavQuDaeccC0PIrBkp
qmpO4cgEY6iJF2qrBcXH4j6/Wy9GtuNJ/F1t6AteGH7YXw3eJTNLPwamlvQH6GilJT0QN6yfUlx7
vrAGJ1QQJQOPmdylqBSRKsKjNRABFtA6qF3FhvHCnPFDJbApdLUI1zxBM4bycXNT6kGYMNJz1c5O
/09MTYnZN2uDWR1tOoq0SPlvfog4vUvOiUlhXivRiLpT8O7hGNOVGEMZesc7b3D6Y+/oK7XDgwmK
t9Hv2wkGmyjiToOIqbN6a4J1Nn8dtdAjzCyDG48hgcJJ18mnEPd5x+o+a4H01bfi9L3A/sMM3jHg
AiiRVYbfay/+pLR5WUzuupvTEHrZUSGl3522SzNlWpyUybK84BUyiyZetrYaZdP1fHSX0VJ14jlM
D6Cko621VYWL5UtVlnUbd6dyTmim6G+qhwm7KgjxMDcdirO+RQ8A5M0073wz4UvMYb9XML+3SVQ5
Oty8cxRZwuoEWwVQ+7tbYWP4mFTrzLRU5lhc5b6QyWeghT+JOa4BvQzM5pcwRkIOvhWHuwRTpe+b
GF9rhot9ENFnmYmVEODD77ATUTksHBAX1a+vMNn2gddnnnFQPbFgvxxni5WpoCbatlQbbBVVg+TN
Ges1358NlX+Vdga/bb0wuPCmAGWFZBHUciOKV7aI8K0mFPsWA/05u87jZsKyOx1+F7hV5hbVNX5l
Q0Ns628t+aFY3z/jg3t+yvYB/F2xxptvJcY0cZHB1qyvlQc7I5unVFhGl6zMAGSFHyTNyg2xg+99
i8qZI2qodxXRRZZxCCaqcUVAXdiiCvHJLJcqnqjxhcOXW4qKUDRvBmZHWilAkaQC56LGZyVRUh2l
kNzEttKAtLf/OW2OJ4HXNTj/mOfz7QsLOMkw4JBKUNeHUlgt400qHow6B/ONV5cGMOqEmaRfJixa
DYHIkeM6SrxDXFzsvR+iR3mWKFIMvm3VkT0DVKcrevwT8iow00Hx5yUfZWpDjoYjRXcp2VGZ0llW
viYlXBrYU9VZxV7lBlmx1f4+m/L8Gs1lbV5qq/+OdCCUSh4HacM9ZY2394zWHNmCHcwlr6wXF+OJ
F9dvELqvFIY6i73mMyYXlIL3Ew2dZ9hIz1Kis+U/c8W60yV0KIaevvhBPBqw0jbLINda1+uQ42sZ
l59PVmj4C7W00Z7+oGLBEz8GudGXsdDxFN5ROwC21TLeqxCNS9wpmVsRJLuLt18YTXGIx2GVwhs8
L6c1ngXR+kZ3qskKh0Kch/uyFUB3Lis0lQM0jrW8Kcu+9fWHxtbLSwSSPvX79V+xReQwzINjklDD
qNFt+J5GW+wArPKli0Cy2ibiCCB0/e76e0/tGo+BuaXikatvvYpwMB0tS2Z3jbfLzCNPul49v/M8
4ks9C3gjw+08Gi4/Ci2UpgfMNr/CproiikQk0PLlt0pJhduXtyun5ITe/+ublCc/BJvrSt11A1KE
SCjvVX+pJoj6NKalMJvk87whWvHn07biqZIfTW046gwseZVS4GqRqhGVes9BZ2opjeqT9dDT6PLp
wagRUOmsq/39D/Qs7z7OyfAl8MAqEL/V0sbj6HQhSj1y4Zdu/4oArzdOzxquvAJVryf3Mz0t32Y7
Q8ctPtyXczdCpOuKNJ+Pagc9+LLylw6qi+omtjsPCJolcxR01To7jXAK3Q5QsTOBvIRr2kQ7whcz
ukUrHMJxr/ieZS3vcR9zeiEi/wwheNcUNdsZWDL3PwWWYyQZ9VDkzVukb0JrnsqcyiEfO3BIbrmu
T5Vdro4JX/b23W8AZw7EtQTSQ9h9Hdm2Bc6AO2neiubk+mUa99Po36El6REndpyWhH8lY3RXVw3S
mnQ71layMN8hMS4AV8zvWIJvfwi1ziZ2Y6mp3b5fhKjs5lAWFToM18VqmZ3vJM8tzLEf45F7EKD1
DzZe1BbdOp0x2+WMi5sNmJKbOXtefU5/khblmtOW1Ue+ur1QPzrOg54yZH5mzIgIP3Dpu+O87qO9
d21xh3FBCYJJKFm5oIlYyJE+hUVTaMAmZD1b0gVyKbMpoM7m589Wb43Jb8L30pFWWc6TEW6kzmJf
dYrtButAdZ9wkYSOC9EB9Zo1lqb4SatXS0oLCnyB9Z6aLAMlV1MFusfS71pp5u7+1+7qurZEhgtI
AuPFFlj1AfSN6QpVA5Ie2mDa46u8u0Jo7SlPsowYll0WHqxDgqRM2/YOcoIhZdOxkUfc+hubQZYp
XF65Ly7q0PhBXiBOPciV6yBscntlG89cwNSf/2mTSEAB9kvZmW0IY3RLcS/zHEt2VXp3lcy5t+0Q
Iq2AXonxatJFL8mj2wsTynHSE7cEflUPLT+yucWm4qC4+/FuqtkoU/EoRIMb7a6Qi0PCiHSk/eC/
M6ga1IqDYSQAdrE4tE3J4laCliL5loqbR2RO/J8Yaii2aV4VWgX6iD5iIRFcc6x4kvubTAgdPz6E
ufLbjTj1h9qHh5he4lsSw7nkgV3tHkzBDHef9wUXUsISHVADIWEe1bNwlk8pLqRxlEjLP/+HdT4O
dtRZXnIgw4TVP2Q8F34QJ6HVjv/cYzAZs5ZEVtkEN3AL5v9CZ+quSNKaU5DpgPHt0xrl43WeWKgg
k1Irjgnu40/On1XDLJKXtKBwUHxVCf4WsBkylz/1GuSiQgAbHCZziirMFSsBB6U7va+pOiR0YoBe
or4hOHz3djfGHFY9I8tfbD8CT8WuJCnlweal+TmY/xNiVGj1hZvOyfxgJMF1W8/IbjmpYcSQpCnR
ACS023kAROJSCEu33ufP2dZ5Peg6z6if5z28L82VWZAhAmm5df5V9qvaczx6kvW169z+iqSzjACX
O6q8V91m9ER4DAHAQ4jKyijSPJVEKGHarbuoX+BVLbS7LZb2BoGAciLwy8WmF0S2J45EaV7LeJzu
PAA8KpjEYOtl2d6GRx7/7HUf+qqTIrjVzjetX6rTaLvtBtS2pdNvetWinu8hr5DNFBssCDkOSs+S
skR2ayJckKtlCs5exdK+tF+CBWZ8TwXd3DGtFr/FTlsVNF0HfTN66KPpOruFnLZGT77t4xMFFFdb
amrNg+UkZorzN3e+XcZE1+J91OY38I1SM/vPmrROjkjzP2x+U2GdYHv+WHwXYDc5pS/MEu4Ipci6
KnYhvNRaGUqA9ce+ty/A2r3omHqCs2pggAb5Hbsa6cjQYoCEcz6oTk3lZPbFHglQt4CGCpBiR7Un
+P7BK2vQgYaaLTTCtl2J4v7iA3k4O3+57vPxTMk2eGSHmTK7NAHIuKJMvUI/5sRQwBf9TuNPVdAi
CdYWcIvXQv8VIzaN4pOFGns5amOfcB+CU2/NjWVDDvnwYa6YP172wZArZ7BQxxSH3JMgl3fHlNJL
mWFFNNFNMa5lncAJix+I0aTQ0d6jspyGk9W7o/F6N4spW+QI+Q/aFwRgVMpNUmnFtIKHVEyQ8H5l
QMF5/U8al/bx/w8aYcqPDBTnMvJFphxRTwy9yymjWEMmJLnxWw3VVKWr7FPADiESYsVpC5nLzZpS
2l1ZjT2rEUFxr64V0/cfP6nP4tS98KHh+hrIlnkIVuzG/Otzc8qII7Emo5mh75UEUhVOrtNegsyN
+AGtzMmpmo8LzOnwDSBq+EIqQwtdMhhXcYG/7ZWLI8j38QcsIsahce4SYZo16lg976T0T0Ggr1nf
/ur0x03iO62f1v+sTW3UolLNnMD3/ylD0hqcN7JSkYWGNjNTCX43cEejKgyLVNp64WJ1N2T+pZJz
XG9XkuPDUse7/5/dW1Gy1tis18M7SZ+V3f82OK/WrsHI1hsm4k3moi8wluFjPQJPKtpqT4JpXJta
OFSfcKKZx68QQb9pzKFtKNmbfrgCghgxa6xobTdNkjT7HAEXame1UcuV5MUJccAhxe6kVdV5jXj0
QGLr8rs6uzUspINJ48wJh/R+HyOk9Q0Zj5WnzYtxl5iF41C4ewaY+HmnIdPItjSFs5R83jRt/4NS
JgMH8Ht/P7L71E7/CKjKpWrfT6nAIHPDhgh7SkD67WxzEg6goeJXaPCe3NwFP3Visw46EFHtpHPx
wVuBXG9Xqt7vnjyKMhM2X4WyEJo9LcoRSPbG23sLDIFU3lfjE+Gl4rA89aSrG5c9ZiRf4h2DwNfy
IkudA2jLf/fQek36+wbkteLqX7YwyRNwnKxVV9yYB+41wIimGBCY1/0aZ/SsTu4jXWVRxtgiWVYy
qeXJYv9RPxc8xkcW/uqZA7ipUv/jgC2dDu7DzFHkyho+IDjuWPd8RGGbbom5yr9G03IO9TBDv4vd
rK4udtTRRWCwzq6YZoT4+KnNuyEC9/QbFC1YGKqavc9Feqt5zSewvz4MixhU9Zeb1GrxKZ4Yd6Hu
30rQ8i4jERVRsi+rpBK03jNG/R1EWNOrUlLR/gJNH9rpQdW5eP1SdaknvNkHWppVUvG8L5ObqK7t
HnjK4IOuYGDVLggdargGcwGj1VkvHpFV2f2JtCBPf8DoNIGtr2jNmsbKKtlD8h1vPg+uSXNz+tNE
bEUB7r6I4YrS6cfxe1Z5mk6zQzD+IwaXl1GOx3v1FhkwzQ3ShsT/i7MTuXAyoOCChgCmH8jxrSUB
6lg2auU/aSslyc+n00L0wh4PsCEmRxSLY9t2XVKor1aDMiVwO/CchOYZE+dWvtJpsxyD8bK1qKkp
07mOhqtED+axz3pXLnVEOhjDGg7rMhUfoNJukpb/tR6yeCS6ikUFLiR7/KjcE5xduHatG9K7JKXL
4QSj9LV4eEiLlrA/lXu4JwFM6Bo4nbqlNgJX2iMh0P9rtSU5yrCnNGknrleKqK/SnjFBaCy+ctOd
8HQlTD9EF1usnZzPfh/mAjJ8wz22tK4lLkbpWPXzr1JLPBPTuFiSWWdB5OvwHCKstzRDvvnYW8xd
09AW3iwTAPLZFOLWk4vjL4KMJSsqbpXyvGQSg0f6W1iQ46PEjbtLHKyx+RtDXuDFq90Qc9FzpseE
HFRrF0vf4kdRBVuG5lb11XiCZfnEclLw5BgoMCV0R1CqnAVQIOd0qW61meLhzmM7k5UpB6uIpqBo
qtYWmqOuMVR9jR4+POjywDzCNEZfBqujReFyeceNKw/6X+fvDNgZx+bWJVo1CvFjGryyFE1WwVK8
IvQjLfpIAePC2/riyLXcVejBdsm3apna8o3iPZChlfuDPJT9tdAHaJkc0d7AWhiSguSfNxucA9Ad
K3Widag2j5MXh7DwxYRX6wQUOtU3JlZz+mOp9Bqv7RADupqH05dx82HxDj8tQynwZ8kTa+83LgEZ
3VQxS8EL1UAeKvMzZvi7hMt/zmz/OlJF1RGro6/W0UOSfZXaHprFH+/FK8Z1AQtSO9wEFdlpl54G
BnTLHHebRDYPawE5xefXW1vj/Vl9bV03ipMWgdWS8eA3svUjb4IpZd59tqMs5HjjHeT+UnuuTgXx
roUZ3EB7M2TTeLSA4vyKXhCfZgfFb8z74cANUcpRO13DDA9FuAvMWZD9GU/8gLV7CA8NwzFp1zRS
mAVxKjnDc8vyd6Sp4Hp/tKNAnVkg3VL3CeLoQyJSbXTfximLha88aY+Ja9ooPMxXZLomePqZkO/h
V7mm4qx8xNiJilis/wMRFC/qTmbO+VOIcFakeRCrNT7LGhyR2MeIjmTDDurQrM4bFjIDi1aM+AR+
VT8fzOvwnk+4Yd4lSa8a8FdnIFbAiB35HGYQxCJfcIY21FIseDCVu3/k4qeFmhkWITdDp5KKrBt5
n9mWiV3zboIQ2xWPgNSiXHHKcvwbmBMb1IDS258xpf8ioDDmCuLhXmdeEzPqNHP0umsUQOt2mxEy
lJ+m1gJLWN5eU3Sauk01cIe7eZvGfwudCVKN4cWCYy/Qbw9txrSv0Z1p3nHFBuvbx2kwW4oewMOZ
AgOdF6bKnTaRpAs4XYctk6IpeoyUW27nvV36SrZMieA3UjxQboxgZG/dt6hA06kUc09emJx2+Npl
GyDQTumbxhBAjb7oMgnQIE5dzXbZNHZyXPf+nxccC9MM9iSu1V8wxd0HEWYpcABkbDhKHdUHWFLv
2m/xHRhClPwcaVIkDpux3xZPTJKSm/hyzw4qs+088t9kwVNCpcQgjejTD8lm98pktMRgCyE0Od3t
F4ZAG6ooFHOLAR3ExQ8mxUAhKZSdrsxS1qlIxN9MZTk8tTldFvQ81pCKfYOjpvmWlD1rfLjb/jCU
ZdvBO9ONJGaw8pD0/5SpEBdCk4H5HDRjbFzDAf2Z8PFTZcYfxiKbDZdae0yRoLDgEbBeP3zUPXZt
AnXS3osHQODuStbfJ8rxOarSOWrjS0nqJ1Xot/pTduTkGTXqpyHACf1VoXmoo2+KFu9vbCDxj4uA
voHVby+6tP3BZZSqe5uo3u9FDM71+qnXVjPpN9cQr/7Zjc5sHMNi2IlhNHP/+cYID25FFOhdIvv1
DWsnB4CZy989M99ZgNFbXNQFSQCvzOkSNwF+FVnebfovkmr/O6oieaUkkaNFXNA+20+zjRt6/vVE
vuX54HvMDzUlvWBU5gF3pSLRkPtgPCgcqo0D5PX7dez4lnxHz9Bf3pBvvLAF6qlHbHYpjz3/7CJb
fPYrwp4ivHvMD3Dse2zkJEpEU1HCPn4ouwhSfpMwyFin5FCRQ6HkZ5ytTGbb+cG3vMo4j8Tben8G
199/PFPL2S+HWHB8Q54pz2d9Wh8OAfkz/EsI6k0dnmK6m+Igl710o71nRIFjQdcHpJvZFB0Q+eMz
iDluePlVYdlyNrflNY8RFZvTWpTvGZoavv4vTHQGeF+ChCzBkbd8ec+ZoFUYXG6o20I9KUfj7PBK
zfQHsdFvLKFZSlRsb8IFXtfBDdQOB1bLn/H7dK98oojlI79SvSk45wfl2j149t5US+1zb9edXzQL
emLSF+Ii6ynoNSb/RwiD+OgZBeOAcC/vkq3jsgJcBYSdGJBMB65sYdJ1sH+eegXdt+AQ1DqP2lxY
wtK7+BU9+zJquheC5L/JSNWiYHM8xQhUW4GG6u3hAH1ADioWzYZa1T4ZKqu3gcbp04eF2q4nb/As
gziIhf37rEazB9g98JGD91H5MbEIzRU1KJcwnJzoAPhsMaE6GPqeDmznUeFCEEi67FuIlSblEBQs
AWkpv9CMfBhqajsu7VfrlkNDl5E3NMgcdoOonSTnCwvv3/oziMxTj2mzh36wtCBTpxRjIPxQpAUF
xV56q4qEpa4TW2Gu3Sjt6VpMwsq6U7VpqDurU/DvqJF22kR1y/4ghEeq6jGGOuVkA5Mr5vBl2ZRn
GBP3PYd6jSc2gsl11HxEyIw5rOcSZjNixHFZfF9UUfIjmAC1PbLfsX3Xl4lIUfzxCbHvR1UfUj7g
D1A2HsiS8gFKZSZme2lLC7GTInnALafUlc1nuB2Vubszwl8btg01QQ7Xe/saCj35nJ1fCm/8+K1E
GWPNOd++L/Rg1dt/GaASV9sWwupwn8k+yDLwjvz8DQSK1tzouXuWTyJjaNdMSXm2flTgFmaKW9F8
k/5f2jxw2l7XTPVvzQ9MrMiYo01iof5CLr4rR1jR1yxO08Wk1tT3Zsnf4O/f47/U68WIko42ieQu
RZWeWvOvinpfYNOI2KifaUIUsAaWmey8tioGVhfT3hDpcxTMtccl6+JoirX9kwP5MZmgTqdiYHEZ
aT6RGQO1b+DCdOOcMBWHsBCStKro11GOQuucbz2Hmujqd8RvGHCyiEGXdhvIjuXTXzbkp4HQ2iLv
AEfrZ9Jdm2GkX+cPWU8EcYor7sjzWOCg3vmQ4bNPEu7vpOmxVa9w1kkuo18TQbi1bd1flx11wX3U
qVA4nXzVkPlfelydtxisC9qCYQGO/jSiEN3Wah+dSGBprQlPtnjFrDTQaBJ7W5Bae8fHVS6bUH+v
g/Id4WpSH5OXV0q/GYH7dQRhtXqu8962jGiINyZWzjERgkR3LLfbi/2IiH24fluvT/q7fKlBxLKo
Kok9pVenw3cnX6FsDY/QMaBJx+/CBVt++I77Qlny61yWRnO+NYdtIN0/VnxEGFkUYYTNcYJYrQ2g
FrMRpYGLCSjCE80nLGmfRhZcV8TJ2/J3Oj/C8qZaOasTS1qC2iDo6QXdRQ04kBSbNFvzlMNZVeaB
9FKZUvSeBh2lbBOWYd6Agyc173GP3Er9LPp0FqFU4uGxT+BVd5Nr93mXJaIWRs52Xvc6uSOMXca4
qdm3jwEBAbopRItXmFLLP/6aBp7/KZirSqTvXoSgjjtPMsw3Ee6tjJPHiHe7CgNF12fqo5sjEi/9
e3nU0yDEC/nfEi8yLL0LM6B662Cen7RxIsTSbmkqloG5zaM/+P0NK5MveZNFveesitiS7rJelYLD
1reWNpj5egBOd/1ruNI+wwNpRNG3d3qSvqoN4mxuKtUsqXlmjKe9C1cipI+VRZAa2lOurfOxdGst
Q2ZG0HcxhclImMYRS5gzUYBR1Gi7Rg5ZxP0lq2Wl2d9Q9ih+e4/syRQYf/tL7ca7jv6yeqkOmXHp
T8sY1glzO2dmRm/kq1giyqUPPrZPMIYaJcZCmMXTUSQeYT4JHzWRNP1EuAjsnvTcInAGO5UykgyS
dD6I6OFd5I6pfP1k6hmSakBnuAl8hcxXs8oqkFddHwgFrqIO78uDfcfnHk1/ZrzSOeABscur1Nq7
o83jS9KCRP4ufay6ZgS86xLP9Y5QcE4SFp1TL1xZOYNqFGpl5DyfFHDnAcwsVUghsyA3HO4uq4d/
7ZSoCEO3SvbzMneamfU2yS8dWkfo/JrYs7Y/nsLpHEXe8ZjPHfZMqIZL1kRG+k975/P7WWgqxKFk
mHcobKUqQKdYFC52EeJH+JV47KPfUXGUWZpg2IArKzxT9ZAZVw1MoithWdSPQyW1V2XZ3o1HZtGe
8e/d20gFxT1q53LbF1lZPhFBTDDlHDB/wugBFyFO+qFwt1PZ67SDNAT5tcH+CwFeNK05AmiGYn1m
4FK3yw9AYbC7XdUMqjp5tJe5DSyXa6kfXRcyWrCgT6rLlT/8cgTgqmxGWpUHQbo8sQel7A+H3NRd
KlLm3ytr/1KlgIoaIKMGSwRtGb1yoVcyJzKFdKsJcWc2EVKqqZGnMiGNQUNo+mv6jdm7zldvvaaf
pGOEpxABdwOyMLm1dZW0yW2qwKUHPTW5FNuoCgl1ZGhckOYJ+5/STR5CnbPXv016w5PFmpHTeqst
c9MZzNIZYZNN4pfrqAiAVmGirGom8Wnh5xHBqayF00zHalYsv7bADNh77V73ROT220CcyS0KgkZp
QSoE9PvLmC8lAAlN1IHhh5tvI6sn/Qg6q715Lw6lr8gbv3vb93+izQrdCrPhkGQ2VJJQ4NNr5/+c
QW0jLkX4Wn814WjRRKM3IA4iWa1cSOTaCmJ4ZA76ZHDQ6IpdjRKO8E7T1WO/6Sxw7tzhli7AURmi
6pyqlGiSfvHEUB8mPFIjDoM1Xu9WlW+N+lwGLr4PkETXDgnVunglOoAZDCC6/1EDZIzrjkmb8X4+
CuTYn1xqXZ6o62mPT955h0YlpCSzGj67UmyfH8kodNrhJcpC1L1hT1GAzeT89lfqzhCtoPTyKInT
cAXtZ9PMh6DkXV4SoUnfbCGCKh9tS55qvRutOCWokGZxkkqceYKSoUukmPqqFUc52gybhHN7dMf0
dFE1+w1Y1a6/H6b+BdjlzImKR2MrXOV7ovih1zcETYOz7qCt19jxZ3bBiuKSutg2y+HdXBAcHmzl
LpcJNmq7EqUZXnR7hKROJuc1OnVqYuaYepHdMHalYlGrYvgKLw9pFZt2Aga3v8alPHrKYI9qWny6
/92MXLO9uCQPeB6edv7tz/XkDK7HHU/7djqd84uxFUzFHpkRSgXRegIoBetscceDE7GOki6fW6yY
Ib/6nt7krChU2M5vJC3B6+6SbWPhv2PpryOzdj+kTnWBwvtaT3PZjL0AvtyAIowoE5KTVVnsihbv
MxlR4ABc0uWLl1eM63cBkdCXhQSJl8/AA+9yNi/fxProYP40AsZl4SjGH8lgHYANcnUDsjQj5o6q
gM0at+8wUDBJo+EVA5+7znIY2zd0R8jR0Qzc7VOEr/MYC0XgOlIYlWZ3cqu71HzNoUgc3YOC8u3E
OYDnWmGCu99Q9i4SwCqXwi5LurfgX1UR5KbLdENGIJoN+mdLr8S0pcFJ9UqXR/vGu7YxQ7dTgKsw
+4CqjwdriY9djJyVoDHjdD9Ou2QPTkQOUixiE8U0sAzzPeM4nWW8x+iHPbQvxgxdCNeFui+lvjDm
ZOQnZVZhTx5BHvd+uEMpU4cN/dwFu7VfQ/eDQ0mA5M2SpvwFEHrQNPwsQmlm6eXOirWqFKaI/g/1
/cGB7M740R5lDzysLNbgE860BOej+GGk4b/mGaUXCFRY5uVsLnWIf7RNK1KzW8Hnfz6nxnpyVtBU
C9FZhTasQsXu9OMGafLxTSbGEPug0xY9F3sds5FF93ofV0W/a/7pRizvQzLTnQToyPzYqAOsciB8
ubOQazM6Ww4GCIKjd+hW5bBZpZXgtxnRHuFQLRmMeK4L6ogTi3pstDOwhPqLmjyZdLiOSSlj0yKv
LBSniLo0uKoQOXZRg4yh1QAaPC0sCSOrJLyJuLNwIfXdPQp5uA9dgKgPQ6ZVrnTtr1GvE3bqo610
fMwrZrBlIVYcE1P25kmpJG/nxhwWt3luc+6HQiWYh7ZuMpmicGUA2gI66s+9WEaxnRtNWlL8dD0g
1ID3TKiBLaV4/n0AngLkRkv9eNoCc6E8p6qMLh2dJHsXQqf1r5iA2MLF7pgon2pSSfCJUN3TiV9v
H4IAmzGXgSPQJ6HhqTtML6GbrdG0yl7SJSJsjXLGlZeuug/7D8XjiX6pGgtQWSg8vqhsH53GdJjz
2+QXY0DxGV2Onf9OZBOPl0PMOboItYCx1ST85XOYX0qY/MpTj4nSkvvu0+vyydoMuFs80kFWqzzZ
82UxfTz9b589OTJCeDiObgq059kxOiPF+a3et5s90GeJ6zvl6zwwSq7OYNs/4i3aVzNapTGqpqE1
+5sujOMGAFpFYI/wM4/tvHiFcpVqPzaVL5xAMVx9so2Zha2/jL8vir/JeUMRNV8SgNu0nB1X9FKe
N2TZEdydz4/9Ph7gBG7/3k4qIqBIBfxbngqHL21cWnp2wZ14Sq42mVB9P9ejKMqm7CFlj8+VsX1m
ONNLrDN0BCm/HoLRdqH82IV7lMG6UbzET1iq05z5QAjKXCjaeVmQ1gMgZHh0Bo8PsSsshhCHTuiu
GZkf6awpvzWlxmh7zHQMT4r7bnXt9dGadqP8enEp+uA4aArI8upqD0bmOQT8tzX6C56zE3At056e
3yx4HlKA6f1MknE/jBn9Qlio7yiNe0riyILcAvKP2GPOBNsJl/GbULzYrkoyePay0J7GkXT3j5qJ
kv9ctMOOjn2V0mhEk/YacsQPMx//lSKaLev2eHcQHjvSb2dQGDPG8BFEsOTaTS7g1vcng4TtVK5s
ij5WhXu7Am0575G/CHfrSQ1tTvtAlK5uzHNtALUb+mR0SBcmwe44RhdQFKEN2Z40Y0/UQMrHvDsO
L5obX5VPuY4qzy6aTsygu90i0P/AbImktT4fihLV8IHGp03i57JxgYaJDKXBJvIyKazzmiicvlRi
aLdJm0yenE+oZ9a6Gl2XZzj5cvMPKfpP0rna2Atxdmlv6HPbd9Xp4RvE8hHO6qL0LqFw0V9WnRMw
IU/m4WJg+SS87mvM2nPV715LxuHQQSHG8IbU/qsA5FRXbGy6sUAMO6UxmUPKEeActs3bzaSpPTUo
78DsmiGvQf38S+8994OHgNJrFb/Mj5C5NFcLi3LF9DDuv+NOD6n84BfHEHqd3sPQk+ZMdV+shIdm
V1KhcrHPrPJRgKTK4geO4iQfUuu9Tfu0btYAV0pSE82tWGrHQieNkKas+1VkpAU5zxBttsyztsjR
OaPsLtbjfWH/K0HQ83q97Y6+/HCD2Zq9vPsyHsyAZb/WIG3XKYHdYPDcUCIc2ZvYR1uz/mpeaeEt
NftVluTFDEJSjSHLhdBhzp58yOjCnZxxKQa4Ht/GH0b84Edgb1OI3fXJ+EN7D6AyZPXQLd0IpsCp
G+dsdbohkFJ2z00K6r1zjAWsPVu0aeVqEF0ZrRiaqbf3tsnfSqd/WCgBIAbU5oNR2+sngZYdV4ej
B1OOh8ouNeOOiSgS4BjOaTV9YhoQheds16TJFRCkM7+7E5BsFn0hHY6ERJlxzx+/1UxdAagF2qqM
5jNLsCOK58olDBjRX1OK+pH0xdw3gLndHMGkjs5duEAFlmGDg5AYSMnv4uz0yjiaUJoiLMf/C1uk
RuHSE9ov7Qn1jab1gbdeC5IH/c2P5MKcOULel5KmzkQ0QQIyna/7zogEz/9nqR86qzycqBp6GatW
Z02kJTo5JAY8gcZHvoJyM0gKTDbo114SXFsVezByeUeY0H4ghx8JC6COKEGsCNKIRt1G2PRaNXqq
uU7uHkcIU58cevyz0c+oakGDhTGJES56Bg8qcvbSLcmjVQvQ9qwmiKaovk9cifGgL4JoyDPIERnp
Wp856+lA/ZLGVSV9R8Ju6y4YUVc39ayx4LIc15TFKQLSlejiNweT8jffngEcgR4/tmpAe6Fbj3Yo
05AM5XkvVsXht+H80QIuvAh7Wjd1uLc15KC0z1MBmdenHbSLLzw68txGUlOeViGKGfi6u0gXp62Z
uVreb4WuuuoFsyVR+ByjjfKsr7g4uFE52pM5pZbmeEOpkFRsW355O3StzKTmrVg4N60phnkeIv8S
XilKBca4btjr17Ardvl7e+iT+9gztFFnTHeytZl7jdya/5IEhp4YU9dRri1YXw/+Y8+AeC3VvSJA
YBJ4Wopz77H1ZwWuqf3loOii/ruomV+pvRoIdM4J/k7e2OJcPj/zvKhSB1FcwtpnawLRAL5pR0N0
LZZmu3i4a++xRIfGcWx70ClKmfzOumoCRphv2S1eCHU+PXqL0UF4DkM+Kh6u4R4fIfNBUeyM6xvq
2hsSA6St8YKs5GlWrmrD6hnPnr3E++CL0iN4rS0ucW8I2c6HPk6azEgt+qbs5NT3Jd9jygQMbuYx
JYj6WDNLthSfFJJbUfAP+z63BgM10hCSSfL+bskcBHMf3T19WQArs5lQKV1/0ejw9hJWa2NDaTqr
uV6J3YwM0SgqDvjv+Ewsx9EAtekT/qLjd4b3NWx8+EVTNO8bsEssEQcg/cmTrK918+CDqhkU8D4W
rC9ob2Nav5OhzjkEWLwFz2g6+u+Opo+FxivyVGTRAvtbX/vjP1Eku3Q5oeNhQk/DYgUPqh6/MhXo
POpu1ldtYuBdK8owmDNIUfw7CmGxcdUPVoEK++My73eTOAHzkOY5ooflms2M/Brrh+0mJrYkoXcW
T6hqym+Ol1jKxAxM0OMvJQcUUjMvQF+DhV8OHdv0tJ4+HTlDnuu2wNcLAmT/PKuVA7WSXUN/SeM/
4H2CjxW/Dpozo7hgSmKyCDOGJFeyut2ffMVRCj+9b1gzjzHKacl+Osd8BOGPujdXZJKiZtD4PxGZ
OCwJGuJGjgiVm1KpJE502qxvTpE53xx0ay5IC0e0FW0Nf7LxjV3RlXvDJhtI4lQmwprsaE+uAR4S
oIjARiELm0tAxjx+AHzwNTwfTqIbXkJg1oUfE+wX/rKRSwKS172pg4aVtzPbfEi9E9e/99Wd2lWf
GvWBnsWY4B5zF41SECW8lR8xv2CC6R8Oa9K/rleuPMa8ed0539v3uF9I6Cz/ifTk2rCCxbMh5tTS
mGjxHiBk2X41LIg41Y2yHblR9fmqsQe4JQQYuoN/Hx2UZCAyoHei004GY4qqAvn/iqijxxaJRjj9
EaQZvZIbiSwk48SxhlyiQvt+EEi98c29qKbLLBcem19QB/gzSXB7wWQYaGlON5/xNX25pn5mfwC8
zFoayp4BjLq5AAaSqlapPlTJ7jtJ9p2vPPdB+anaq/v21TpD+CVvll9L6JqpKp0YyKUnHxhCyRQN
YACvHX8/5eXLDTnc490A3Wx8StHl8iXrCKv1QAtQHjwz+/a5u4XdExCEIcb0YsmstoaQB4JruV6A
SL1mkFcII/nn8Uu/Z6XuHibvmOw+u5JrKaMkgr9qE5rCk77R3wdXMi5gMUvploRs9ripIrdMDsp6
8FXbI+zqo3n+2negewKKRgsHLJ7Frhrr+HYWrloE78HYInXZZSlr/2MALjyP1Te7ukdJioNlNLLE
fM8YJFn3emdJP/BiiOGoHBuQaWYvUJcduEuvSid0XCpje1HfIrXPz9hAcJ+6/iyG7uSe3DXjgkpT
XFtwfIrBbdmTJ0PkVfVyTx42jUrX5stnmFWJkTrxPz2QxCnCkqBLuapm55A4AAvpW+X1dqkJczvE
7UdHlxtzgZesKhuq6Kv8QrelBMT5iQs9K2hgM1jGjOOnA4PrF03NttFAvgaSTp2UJWxU/3jUpJO/
9LZPkPK4ej3EJ8bQyq/zQkf3i63Jq0GydpLLoTFf0nZJ825xIKlFM/YzbdSrNDZeklpx8zT3+I0b
S0cc/c4ToVZS3Nyny/9YIHL/5g4NZlKOYlC4dvkhGHvrBfLlRu7HhWWcZWufkPavsNFBQVrNBLqH
inWC78iOd7T9Roo43zw8xilxRJvO3KtNqxWc4Fgi0KLD1aqBSaZvDSgNFDV9G9AFYWMrQM8LbjJx
wwEy36rBs1yvaYVN6GMtRFpkdyXfOUzVws9C8VMGlI5Yet8FKqU3fKTnl59veS4wYJmR1JyOYoSL
tmumIsZA5nKqq9oHpBHWApB9YZgCnGyUjpGcImdC0QBOdzYkUM2mlYBV9fUiHbc1pfHpJ+o4zWdi
UXU2QXVrWmmGnuKNM556KL/F33WyM/p01Xxz3taDKbDgzZt5mQgXetYrbtyJGRQtoihfUjtc3Qo0
UqeiPKAtHkCjuTrHBLxcwMCP7JGmNZNgFZ2qsY7FMaxcN294Wfiobnpx9MFhvwh0dPJXzedVLtJH
YZXRNGaqFxDZEjR9pfh8P6RAQigjZEIEBda8y+a+58mf6OYV1klfRRm0zfY1hc9u2ZYRRcBLrKb/
wEywukit0ylqo6RW+Bmdjle6mW9HDb/qsBXpX7Z9rQJMM7Au2UQTMOkD8beZvElaE9IeAnICehMs
rEuUyohFjkN7/42FRRI7NL1QKG92opx7bXKDsZgoewU2LjWjfnC9BGfZ0n61kXXVqWberdF8rM5T
f+vdOGaxFnqxucI4Y62Zh44JjHhcbB9THqete4e96p9V7O5VUgOS0ZoNdLm30FZk6Eo91nk/JZNH
ErCujQm9XtZIGfW2OWuhsSDNIr4mydI1ZTYly0EYLqYK97Tlj1UJHz6QlX0Yqt50Ivq6ezpZsIH5
YuWIlEjv5fk3vDmRuk7utFDdt8C22wTGfsmKc5N5wXSihZJynyh/1K0/k2Wp1dvUp02qXOS3hsQL
J7ICFVW6S9ppEY3liS9v6vntGHlZhW2TmTGnvf5/upJlC/p09MzfLdWmWpwb+4RSnhGmlNpdSdSc
KZ2A8ti0GiqbJzrx41r7VNXlz6p/M+Xu+b1A+ZC9lXhIwlfFR4s8I4jlG1RPcH/c4FJHR9xyEyxA
Mb0wmuccgnPjdyIkpRy/WgnAAyO7B3ny0K7KaRr3DVaYQrjJxWf7T0xpZu99iNfRoLb55Tmmq9Ee
TaIw13JyW3jq+C+NmA/0uOfYutOtLBYCOOy+Rwlz3hue/YrLxHwcjdkEEOMHf5mwmjhHxjbsyxZg
isUxS5m2EaKhPZSQKK2QirxOF3NIKKskJepotewgEinmvwAEr8ZqOEC4oBglmPdywKI4ebesvKFE
jGO6vVEm+T5kHrTff+vpv6F+KFDxIQLyIIptdm+UKDU9lP3ydP4EGSHNgMym8vX/7OEM33QXILfB
NLmkOeP+AXeMRGI7C51RUI6gttN8/E1tK8QLMV22efMB5aL6/KjSxstcZt9mGFt59Tc8ZO8x2Dcf
+X/HDC7pV1FQmQRPqMYA8v7EtkyvbRdgoI3g5SQ+YFYp+qtuQ+m4UO2zMIB38k5+8jJOzaM74S3T
q2wRFuMUX5Zgw5l0agqg7sCS5A8CBk0Q3L+X8QJXiu5oaYAvVwSbuRSU5IQRmmI+7UD0liSPPNbz
PzeTxPf/ERG/jx4jHF90SRu+sAOrJ1CUIsdyQ3SqXYPn3mgkBm0TSWw1Y+jhx+EnxLfAW3QoguZ1
D/KqnfMiPulAA6tjdWJuuFQ5u/fLRt9OPbO9uIGNLLxha71XLHP6miFRD5fJPzwb+BHZJAOBWj9Z
K11YeAhhXYnJbN1CzOUgZZ3kURd1se1xskPGZlzgGvfoWLR5tbAtoqUz/1e1jltMiiDwwTnJtkAb
59ELlQGSGiqj/bctUyWZ9O8lfXrK1WxOfdgbE0TgKSCqpSGGNWOQuu9gsYm6FalyjHKOoNHs6mHK
kIltWlxwp6sgyWAfZxEjyNbpxSZGXMsBw7sxuA14xKNj/9vHNKHuBy1x1CiFDXE/i/+o+RHRcjPK
pGo7H13E5KKt0jZhSxoIuLjSY+4GYgYP25aESTfOzcHtevYV1F/HNTzMLsbFa4uak3bsvC6a1ULw
R42DzCKeOMKq9v0QCh39ynDfU0Bh73U39Zp6gGgkjvIORYvnE+kh9NTGqanGPq9nJMII5zFZlvDY
E9lVHkwkl1lL5korObUw8qJHhmI2xnpZnSgaBi0z8wITv6mSzEEggpJyLetcLMTNWdQkFBaoWQH6
3elCCOncGMb8347u0TPI4vh6Rpbhhr/uFgeJAI28YowlKvTR1lwFTIZhOBPLI4Atwnqh+3Pl0nlh
Zk/S5oVIeuVOE8O7L6AtG0k3gjUrilJbjNeQ4xhHDood8ZXb/maMoP9XPTbM5+Ilb/qq3GkYE8Vb
ypDkDWAly68gR85bqBUVNro6iqLzNDT5LD4JCKUdY//KChzyZlh0m+tO773PsbRLOX185DfbdjvW
NzY5dXC3DOJ58mxF72GU05zVx9z6hyIBVF5Bxr8dqc9j8oVAOTShSN4691z7hfvNXsQNf6W0jK7V
zlsCWd+1UUsCV54GgngOXl5l/RB6nCbYj46cevmTtyjDd9sbDDxwNO2sRbOw+uOSdvV2/A45S05i
3I7x9bNy2oYEWo0nEgQii2iJBeVLp8OT4dUxBmiTqJC9eG2m1LwmNz5xcvY6osQEqY2aDuCT9+9x
XhAn1CMt5YcI14vZeIWDVVUGnzX8XkPU5WZuTg201qIbqdZF1oUlDMfBfsI2Xaw2mQUchHZ23jdv
P4GJWBeFASha0YZGa9QXmAxKQzLx/WdfYd82jV/hnPkQtqbp8Cijrr4Y/V+G5PqnxekMa4RBdRg8
bKRdvf7lqzcspxssMlcaykmRfroZwbO+gdOwVT98yB+4Jnez6C3GyXYx1+0S2y6lc4YSNMvo+ff0
3BQZNO/cg/wQbKt6KPFN8huoqxHAxPaa2BrnpIWYHuIux8z7mKC3GukguiYNklUvNup882+OLZDX
Jt1MySilsISy+PUIXxqLs0WYEf+maJRwjZT7+zCAHD1Ak4oRK03AFKO6E45iheGqFGsyfUWqEbga
MI+MOgNMZZqrytT+cpVNdtUdPW6TDPMKwUJJjImJ4wTUhWu+zmrWfNDk0pXEN4cZ2Ee5GZN+KF0h
/zQdXs6IvgGhPbQaXMdJk0dOPLnKC5cIb3YDwFfwnXm6kaMUx803s5CbN5OVMcm243ayTQRDdPWw
xT236JPgdM1yWxxizP/mFqZP1b4cvFkAuVo7AmtOVVktJi4CH0zibOdghRi6T6+PnlTbc4EQ15uW
hGnglfr7HW/bKbShB0bjZh+Y99TCStfJ12veRJHMNvkq2QvEQuR5unoKCD3tSmHWhl+A0UCp80CI
oAaS5o7C2ZyrZNU6NIDBK/H4T0WVZYx9KQSAKBJLqn4pv6EkcrgWK9sudBgYePFTMh8LrgYL0jaV
FwyO1Q/kDLj4M/CyRoxOqp0o1n5JffH8cc4Xxgrgq9Byk4JPfzJjqXVW8QyAOZbC7/txpoNd2P0A
8ZKvfdY/q3ksNfvRfNFJG9tR+aafE98CAiQGM/UcmDABvGNFTcJf2Z1XKqKym+fc9wg/unQWaTJg
x05ign5tv5p4m9eGRss8dReLbIj3WjeGhQi4dVDIGRQ3tT7QlXFrhNU0c/Y2buSlGZRGN81/OFL9
nXXmeziVw4hy3A6p/0DTHNyFC9A0/OB870WSKszB6H56tTib1/TazI2desXE7UHPVkYzBA0MuuQp
6c4UoSrSuhkAa5VMStoe9LNdf0eghz9F3jyn4WwBgYHfp3Dd8DKjtDFJpUwix8q3CaOSRKbWh+1L
VAFFVfwGDFVWiptJW/aJ1Jatat8aBGSwubPWCSNCfitzf/ALZ2zWmvc27xtrbb4xWwT0ByKeMemw
RHc3QuCrqjTjCoDryHzZji8R1/ns67Khh/P4Hu+6ULevR9lLDeliN9zmkwdBNN/CjDsQR49+RcZJ
G4EDDV/lvTun0YzNUYbcvadWG7DEefRY5gRAAqWwSEwzH9hEY2ItcfpMNOv6AthUp2E6x41PTZFR
ZcnUD/WpVspClVGY+0OUn1cis2ftFsXgfU4OxSwmMccwZ7lAB6d9CsOS7pNilFRjZtefU6B/PiFx
9f4hOw/rPS/mJipVU0QNza00WnVm6KIGuqPUc80f5NHbLQdzbGQIfS/TsM9axdzx14kqF2vByQLq
Dg7op6BPeKmG837yDfovYRjXrLkQTOd6ArmkhchnzH2AT/Ar1KbHcLFwoG4oZqs0o0Tjz71t7cew
PUQLT2K4G36pCE5SxiRgQbExudqrf+vDpa/bhEDtxgTKuVLcqru0AWO4ehQvJiVM8jr/DNz1EmiH
xI+FIMZhM0dfeH/lBONNu8psI4y6hE+1Or5JtCz6dnA0dbzSQWfJ6Sc82cnQ2FjQ0YfJm2w7bJZ6
ScvDNT78VNQIRjCKCdTx6+7eG+StSlGup6o+cxSwRHbJP+Eb7oMYFIPkNxkd2N+JzuwkrLskEpnV
gmmWtttYqN9rZbIcPFY/2tE0tneL1ub6S+EQoCcBoCtFU8+QVdLQeli8rfAGrP6iUbQ27LOgSU4h
ZxkLU6bwU+NV7dOPB/sC+mDd9RGGgued8pmD84zA09CpyxZJwc8yyOtpbihD2poPDLa56dzmyHO3
tCsISVdLi9TTbXXoPf9DokBRhJburEK630RTdY9i0h8YxykUEY8poN8QBoav5VVUHUYdmt/fQHg1
3NXgdPEmcsWl7w9oum690T4ozNsgip4gbUaUS3LpTWRdwJ5Kj4kmaflTYM/sbwyAYnPT1mw2KSH1
HKoc7FovIvWPY+cuD+ePfo1nU9y96Ik1FQxlUnKgaOlKfRyj/j59hjBhROpKamtHsLwu+a7z9X2s
I03i2vV4ETHNL6Tej+tvRr/LiO3IysSmN79UP2bzY9PKhrppLRVhCFn9vc5OH1j8Gylv2G6MNG3p
nEAoZcY4oFedYGlT7Ct8BBB0TyzYu2OhLm61VZ+VLaUg9Tjpk+1LbWeQXB6fwNiQPPM7LQRP7O69
uC/AIs8nPWk1V/iQb2IPZqRxmGzOi+/2Gf7dIKWQ1KK7UP+Oxow3qQf8hg/CGva1UaUgdxu5HFtA
CyCJWjvEag6fmGxXzg2t6yADUfL77iP/rjFNex9jyHaYBpRulVE/ReyPaORMoZoWJv/C5brasAEr
C4AT+2d4ZjgPcADCqalRXz76TV1E7f9TjX6ihFjdimnN//Fne/OzMM33Kpz1qe8pzIQI+GCOhiTB
jZXZ5RGe59z2r9T04pQv7Oh7SNldAQsbb7CcexJepL3VKMhAJX+YPorTlu22fhUFne3pymJ/VCLs
xkI9HEdAdiHNwjLhRFFcQOlSHSJN38ivCNtnu+jHnoFrwREkoP+axn63vzV36gn3UiB9J17pb9n8
+2uAS+hfwF6OXzOjze5olIxGbcQQoxfFzU/aN4+54AZyXnzXoUGqQJ67+Jx6G/gDOw3RMlD1EC0t
/5bjOkM8jlmrg3uic3NIwownhtJgQ78MWopfEdEh6Ju9NSar/9T6o21GrWbOOAO/ryFCYAV9st9K
idaZJXUPSyA2lATA7sbl42yBBOrM+XEOdWWazM4H3aOw8D4LRiE/yW204sTcnWO8dgLsvxZv8FYq
kO1ybvbrRpxuk/vcIFPpmKzWPr7gu2O33vUF8Zz47qjOjRyxqldZl8BMA59oSN2hir2Mh7wgE8hp
r4pdKAWSpMgb/ti0lAb1sDj1hYuCm1dO2B++3+nI0fZ0Cr561W/wauaoR/kXEQUfvgxMNZwTBpAl
G3+wwIrGdK9hMBIp57zRo5lzjd3HRQf1qhnKYB+ihavE6B5k+0OoqDsf01dFn4YMipNZn/hD2Hmy
ah1CUxdJtH3QCQ/QZK4YAQpEvGUCPpMvAPbvUUAJQQUvgkpRZO1+b95LIM87ybuy6ZkYQ2bRo42c
6T6DAGMulZG/7ioQ3CAOxv3vYdREEPKeMMRHj9wSMr8mi14wC7ku6HA8Kdi8TcVp2s9/P+sUKb3Q
qMd4BVP8ZOzh3Lqv/mLSnMdGpACqpTxifieyiiomKgYQUMKxhd+Eqzg1sAxROUVkhSExcLQSZRfl
TC9zBt/dYsfyY2Onoa+mS47XToYyVPfkFHc+nS0QMKO7bFYq/guY0/jXPp1T7muo7hn7d+XdZz7Q
kq5QLHOnZft4sQQDcPLywS4TfmFva2ww8CZtsHrYxJZAz28XO/xsp4eX1/cvBAkUHYurIsftasyh
LpIWCE0rX5Mj/SmHo81GZ3Vdsli8wof9nI8sjE90IGseEcQqyxPb1EGsCJc1kL8wXTIhha1vmmdl
bhPe7Y6Rb72JSvLUqu6EpoFyj/z15uw4ZQ+bRFZhQUQtkBukWzbFv/hmguVzlts5LvDjo6Fvd8Uz
KGqvoIwWhVGoXnDtDpY2Wcvt2MCMqeEweWPoUwFuax9RNYs/3kikChrMHax69RM9by2WSG+jiDjM
FluYLE368h5JSq46tgKRAUugn1apZeqa7bjCn2kYZ2vhoA/eKRW1bOC8UP4nhuPomg50LPr0cAdb
zLPwKfO22mZEVBQQYGXOnwgfnpA1J+5Se2H44ykiYtQDZoilJ7bfDPOlc/NtwfHpDQXBYnMhZ3Lp
X3ecq1NZkAKd7+xE3LeYEMrQcE4NUzETiaYOuJjuIAwnl+pUotfV70GwX4Aez89Q6TR3LcBHV8QG
GgHdyhAFwYUWHrhv4zobjZ7HwxJJHh8yoiYNNZxR1tUbYh4E4emeAxhya7sqMTulQ/MxW0lw1GZ2
3Nkc9vnUuc0Gqv55P56lNyWzekVnyaivlSl8Ex7CaSt6cdqm9P1BMgc8eDGoHmWEQg1PZYo+Rzef
1uIPUc9W/REDmKKOHqui5usnhfe7Dwz5tkOd7uCRvjY4KjiwTPPMVwWZUjqQMVA/43pjADsDz3bM
Y7nMzG37vXLsf7l1rNMJxDqpUJa8TATTrRQMZw3FGy0tkwJD6UMs3J/djaciQQynqTUqC9g86i90
Zv7kxJOcnimqUoPt0/HHV4KcF7GHLseq02U9D3YTMFAK9Q+vhfZTStbkatmrTCLk6c8Bce+rwbN5
5FN1XXYzI7GfkZWDmjDYxzkMFTJwEE/CL2rKUEGkEtrUlUyfbShRQV47wdWR+JJwXyI6gcbqV6V/
xOHFJoyjKDirLmNi18JD7u86ZJi9N1S5xKNKr9NItn+kCAl46MfE/xPMcKcq63E3NepOmrHqMOPf
iXsAo/FsLBZl9W5MHB2kJ5sFMTRoM+YE0T1gKT4xi4DyF6lv4D04Jlj8t3M6zNudThJoyA9ihrxC
JkYagDWql4ez7xpkzxPlqyHA5J547VLtt94sMU1pMKrNjgblQYIRwV5c5w8cWVLaxBk1ISDqGIVN
4LcmR605nJDPWZQga4aq5kcAcdKE8ReuEKFYsQjZFeLsOHOOA9vAuaO+ATiA6G+qWVDWaH2ZpoWf
pLUuxX7xKvA7cGkhbC0KFVHNjfrl+RhtC1susSUouPM9zPyDMcHhyiVKTGIDEVIOI34BfdH0sERf
XJhkAJ2diII7R4yir0Y9HccFqVuKEH6BT37tVDTQURfyZ1AFtck8Amyn9sBhFPVbqrfYsUi2QZRw
Ek2N+KXmwTWqo7MchWARzBDGlh0woe54H+acBH+NyUkDoOluoWTSmhwI9UEfBHqiIUf+oCDc+hyz
ftEr8mZ3b+wdEIwRnOR3k8AylodW/UweJ8UOMsxXvneLd7sBBxNMgd/dr3vNenDXYM/79yPHO1RO
mj3NdGZE32B/FnJM99Zm8Y16lU3Syga+JIQo7HlV+j2Jw8cbF8JRu7eAriMDCUSrqAU/eOTARmFN
K9eE30733DL2p4xwoKzfeOMr/EJho97gdVPxr0jn6rYuuYlVLS+9ei997qOHo5+zzbbWxVVTD1AG
YBtU5JTjcsiyxqN3ACpNHimuaXY5qjUCBjAB7KqAAvdUjQU2tj4bTvSoRjHekwf0JAUKvHS3L77/
wCsv5zFr62nEZuB11n04p2DvG+9AKRn4RQEg33W1+zgULR8Kj7xRymkh7HV9tIDooypA6IvaY0d/
7snH8i2Ki3lILGAjPOcjaQcP5+FlG1BEPopgiK8IZ11OGkVMPH0uyjTpaGY9bn1ASh7xZU9GrteT
9C/vfDdR34zCHEUxID25eqj+66mB4hJQ8k9ylyEjmKLIJqE2lv99mwwx0YoZCcBKL9wkSJQAuGqy
T3/Sk52lyO+hYyQZy0oCfgQXF3PIiEcsr0ucAySeVB5dTLMwDCZvFEcrOumiG7Ope842qeCOOFtd
7nxp009bFxMR96vsHBvHPdKbnABgJE7St7N/dsFQm8fDzWgWXbcfTEMZFQl9HTdCkFEU8AO3TL5Y
edauSIptFtJAds7jCp7JgdFw+Vor0K1QFyz6baJrIElRizbXFWvXoqVwH+Davo8Atd9MkYE360f3
MNloxWXeKj+tycGOcmNthWsCbf867NioUMv4IkhpRRgU+30HIkGyl4vSQRBnUf88L8bpL0m0Cb4Q
3OPpVwQS6vl4pRg2TZA0imywd/76eqOHg89KaBE2wN3kj8J7RxWY6OlqmerXA0lAASJOjDLJDPUi
dFwChElJKPyb4XibZRd8e2yZC/1YnYOTYvcM2U5pJUSinK6e4SuSG4F2+iCt/XPpkmQv5NnXhD9a
3HtdzQ6ictCJsLfs6F+M/FVAkJSJn48NZEz+KAIn6bveO3pVMDI/FMBDogrd7wvY5fy6l2oEyzBm
wO10YRjiyu/puDMfMjStu1QGlZDDFriLGVvS6tz08FxQYAjlvtrEa7G3FzN68jopBhBgMOCruPAo
97CcNzW92Y0E/dRCp+WcqItwqBX1BhYSxV1Y2ok0R+pNCjngMabXi9GmkVW5zjbZpttHRFVFVFNM
P1Y5nZ1qaHCxZBJZPqJXA58IN0WqmQO2zh6kIwRCaJ4T2WppqvKz6X54hGxnQIBpoCItFqDbdaJr
9ypB8vmfjTutkP2Utpnxry12qbraIRga++nBhS1pI8GZsHftQ6SEDVH2mlhYzw7PzmUBTQU5cSwr
QPaSocIrfdPMnTl0f1Nr2hri95HDNEfLWiE37GZuYQxbDApICi1KJpNFo6b8ZTzFi2w7DmofD0FB
4WqJPFzMwpXLGswquJ62X2fU1FvJJUBJUa22EdXNyHLg2h+Ov9iprD6hsW69s7ESIkA74bffIvR1
1ETvLzGx6mdF3kQpdfbALpknBimarvxTf9SHpk6I4nijQ7pzNM6ERwOWNWPkkhsjCnJv2YOUR13/
+e048RwjNNOSkDN+HA5LsuJCio8MLAEb3VGbc4H99KZWIeYrVXjFSpdclHFCvz3fE3B7enEnZxRX
BKSC5aWTR2QRjzn4YIQNVcQ84XCHGaTk9CQrx8s3EZ9r4ikRr27MQPe9nyroH0iYdOUy9Zixpf5X
A/tPUEeQnnTywJCc4TUKY1JY0Y1bLP3FRkco22qZqJ1qayK0oFKBdiH3+ElX+KYBGthanvpQ0/lp
tBtaq+4L4E/gdrvDXzZ5Iz3Inu94uL5aTMrIjYqut02FZR2QOTMpcOmw7z3MXRKTJXZIsKLdBpnb
AJ9u1t6SYXgLL01dwNzi0MkVxYh7wk1aPjvbWISzNzJeLVmhqsUVfj2ed3NYEGPFMjREs9zfZmL8
Ts+J2L445y5erA6B02yrNvagFWdvoF3m3oxweEb9bHOX8eikwXnaIgN+9hDVZH649255CbFQOGRm
fGUVJHQFlRwg/HPiqpIBT2OeBMcLrdr8JyV8j421JR68e89GIoRUFyp7qbChbA1EDtOD6iImEvbE
dieRlpH6mihV7wlm/w119/sS/acEao0/LYQyxyngVDs2b/+47ym3kslOMlYJR4TYgoVXhA7Mt90Y
aslHqFdUUGWZE//pSrGKxcTSN9B87qQettYohGXevs//NUQxnNzano8BaJ9dADQPH7WQtVBrIfSO
zESEPctU7H2ZUzkHsxiuTb64X+kBTayGwDmm9UNaGoCl1s40o453L01WYeVeL1mfdnWjDgHwDlLM
MrksI26rMBbErG3wLHf53kqChx+Tgbko06XxCFlzQg1OF2WxAEzD17TbZXY58inhs/R5JWSR70kh
s6oZPg7u/9aUQ/qrkYDqZNrY5EKgu5VDS+nY3G+AfcvjeZgR5rrYqD98E+t3PoHHEury4p9FsodR
xuvfqE+vO1egOCWrWCljFkE5kO1JBUGBPPCJI77b3+hb0H+osEjZc7oji2N6T33jkFfp+TT0Vf7/
JGncgC/obfqEArgtgXs6VkW2nmFyv7vop29vJk0OGuhreP/Y28lhlX2xPbJ9jNgrJohKzlVoTAUh
fFF0rRNbHFDwQ5hBl3ydyEozz7cqr+PN/O9J1d7F5X2uWrP+xdtKu2TXVhdJybRj7bqRSCZXOS+W
Xnv1nfcJ09lp5c+ubfmJSP4X6pANK+DWjLnihcrnzE6AnrSxEWJelkVNNvBUClwCGobUijiSdeSE
+Lp0pbWLJiQnGHLb7iX0bgW5ti3ZQdprXs0r8J3Z1UYLFP+fWBxEBEOLbJLO7ZoV9WGh7cixbb1Z
nLVaeY0RX//0fiJtmSPcQUwwfwfD+47U/t4pRIkWS8OwVqRFDf2gDz0MZR+rLcQcGHdVTJfxIV+w
fwe9rQ1tMV6rnUe/ChqprYblvAkG1sIE/BSve96Wg6oLVq3A8lqIJ5dZ9EpUjWlBrPKdpSG4U9Cl
01yTZaHihnZSmod+rzFj/mOu34k0d5Lj+ErAO/CInbn3JhmL3FIHP1TxJmWA85ttf0bKiTlxctKp
WxYTeaRlPw5ANhyK/bnzAYunQqfwbE/+0q5RbOkq9EVhuj8kbZ4y94QpxTp9tnn78qcIqs4wSzNk
juIUhqloziIyIvogKn16JJC3LKekuswp6rO/RK28d4O3VDnNa8u14fvAvXmVasGjIVHmggM5NA5F
OHxDVkwZdYY/Z7KxRYWYKYcw8ckmq7AM4yD8JVs+fiwhe0i54I0+2TfOmMcbsdFhQ3cpcp8aSQuQ
1KL7jCGDbwKP2iUPskg8IiW61LmfYN+ixxkuCs0X7qpJbOzsdhhi436qf7OA47+Wbg7d2Fe69FZ9
Ss1eQ3ztGruL2utzfO3gAMPtHRdIoR7KZEuNh7HQ0+eEeJew7LoB+hPvsUZoXlQM2lYPzYFkMCVE
5y5n53E+lak3XosqKb61urvTr8qzSaljyZgWRCT2nlAVSWg3r4aAJSkhfzDWQAvuFPHkhG+r8LdS
hCPOOjMczYMukgEB2Lrk3k2PAS0x0eyImvQUz/1ZEm6EL28cGKXc7ypfdB2fsGWUX2M02tqVE/D5
hp268gMOKyOEPOuA/OUkQGUvP7FbWwOst5rVItvftug6d0hviq/pe3QKk/7vSTJ4LQlD5MPxL7I8
aJr+zWKtJESY/LvzmKMUUeG0AnZtRdtlUZfxvphoCrkOFrhmmKY5QctbCY9+yp5vnrTEF5EQzahO
c0m1UlZZlKaJaLS0VybVtbDS7QV7Gqb6vU6rSNlcLaZQgWWKkdlHjZWK31tz0Mzy9rMrTrH5dBO+
jcqrr40NQ/W1joelLutuvcql7JWga0IQ8iXZ0Y/PnFzwVNwN5Y6Pxoyth2eTFfP2l7E4uCbaUQ7m
2Lh1zxi4qa0R3Rn7/lzT47LsbZPYNe2gxRLVrhNhmTC9OQ0Nur9Ej90tKnFFsjJlTaj6n/W10zFw
x0OGnhNiLr0Jb6Ba3XIpTK1ryc2NGeWxxlBjv9co6AywWLvW1D2bfLL7g0WMTG0lIV3gdJ49AS2e
17Pc4uT9XQewYfyK3L60U77c09Pw3Fefu8lJOlEMl+S7likv3XiFdQRpcutYgNSs1p48NsqbRQwp
12D6qItnMVyLf1oxfUKOxrXgK6kPzEIEjrS+v4/hgW1NUS9rp+a1ZRy2pZlWlYqHkRjYFUdLxxhG
h6a11hni7yVBLi3Hu/Wp8GAt3pDRRKXj6InFvRQ7s/pkXiqdTzqf97/KqcbeqrzTi0yXmgo+tnO2
krn0zf9CKI5rQ01+GUYK5smS6otP+D/HQrVfi3Zs0INRvLJdqlnzLQKdC3cqfHuf5Fnhmh/2FOKg
FgRnzhih3/ojgPcB5iSTFnHN2dLoO6BWVQoZf5Wd/eV6tyDdNqHXSlmU4jeHUJAesepSZCgYgC5f
YHG7kVvuZz/X/UsUYrjqWOcFr7YHEnhG3UdG4A8iHv0qT4yQvpICgYtnJ549IdfuHCYJVQSNkaPG
iUj3BdRCMbLdnV6K7HY3vtQy+sDGaL3LnPVWstBfkFHwgaGYdl/NM9Qeeasy2QSrGeMCx1KQt39p
CM+PUK8CLibzzOU7N2CmJzqPAjpbJyrEun13eNHC11VMubZvw3Jfrzx7S9TolNBGdrhExxRlgW7X
67kywJGuZUgQfOkclLSXr6zb6YLN0oVic1t4FF8w+murhfgyoCpO8frx5Kl6yIRileV0MZkzlPYY
ufeY2JmNuwkjqI+XQQpxpouZ/iwvn6wyRfRXcbv7uMcrk4DQ7YifBq1AzYBPPUYFJ5RRXn9BpbUp
5iOD9ViW4fbEtKLVhrLC9/a2SPNudc7+M4xEF8TvhUXK0NUbNsEuaMRSzvONLvW/9J/fkmSteQdT
UMVGIRbmNkBTK9Z5U9e6mYdorgIR3ms+HfxFryIYbISNA4Y//DFqgTOqNTKnLk/qnEcgl87owflX
GnyzliXSFVSRexq7X9VYd8XfKdO4214P3S2AAnHCGlQp1NlYueaii0dq0b+sJJTFXf2afH6OTniA
zU3v6Byq9rN18nowfnxYp4KBnxHYFmmN4wlS6rVMtLMDQXKv8G1gV64JtbTCmbl/Pr0rPPMaOjIz
qNaPxEo7uIYxrEaA32nCAVCA0owkEpwS4rRRQ4wG7X5co3kYQlvYZmYlxx6Ph1pGPUADUVLH+anM
JrV1n/t+fowf2ZTy7bflbjnfb6gwgTtqv0wMR3P7j7PElVNbnBNKLVroCWD2FIAn9rF439bUg7I4
13cMPklIk9cZrpXtsenYZSCmJIooOn739emzIfsuL7zEp0+XbzqCX6HtHo8mCtXjFHrBJT8vO9fR
+0kEtK0Jsom4Xe/ZKyu+WF3Cd82XUlYm/WBU4+beVawDQbe7vgHjUHlUlKDOItY/veyPEYwoSOC2
WT1af2j+C4uA+XWlBYwcViQtYXSzH6Y7MjZQaGKlL+tLEoIknb9kKO4WGhzFmx2PX5Ln9V8vm9Cy
3cIJCL7h15KZReHzWvmmThP3zzVbROQhVwcvS2YONMwBGJ0qqjx0AE7ePJQJDAzLp4q0udRlXXgN
W9vQfztyx6mdaIRWRWp6AmN/Frxr9OYY96+h+TwN87pXGehZJmNSWNM05Nkg2Gyvg4vKxnlntBz7
dostpmN5q6ZCtbdIKnw1u3uRtjtAAF8Soq1EN7C5JMUmoNnIOHweKtTjd5056VAoBFCtQ37cl7la
7a0B4IThQGxfO7V3WhjKlYkh5Ki/fb55f07Ra/Mrqqv1wQKl5uQ9NZpHyC21G54G3eWYG7VZ5zB+
L/gIz+BE0GC4ZCuaUwu3DpdBltSENzfEduB2FhjLygh2eEecz6DZbUaOHgCpc17mU6EveJVcCSYA
efdMqNZTs5J2LRQXd6Qzed3PY5qhwgNyT7i2ta3J6PUkuupWFrvZkTr+vOT/JBN/U9YOtLU9XP1s
y9EqnFjJYCjsR+sCvIdaiVB5AhO/Ns7VTxwVuZBSVzXXODvzUxHAsOdIibrHSm1ffg6jaf1xH13U
iBYehBPIfG7doAN1ic4yRmzX0QhUymjrKygN542LpjZpjOBzPwjgf22KoqnEvGEzOgJrS045Jnve
MHHucZ2H2mBP9DD9q7ZTHNCiWiRradO6x7sPqZU7qW5Tthxhfv7nENTVBAuOlzh2CfihJAntFaiw
jZeMAeZ/ylSjhPGOHQrMKuQPGKn71egIAfC+qjWtynYNw2XGv+l5DL34bDKi07O1rs2oNm3MeWz/
m/FAfAtsVAms27QysJwxpcgXIO274WTG42cd+RGzU2JX3zXdo+74ZqskcXCzDNulUQwtdWfsUbeL
2n5XOFhsrG7SRxCExRZ6FT5pRYN9aGqb/qpiMZLTJIXGnetjjoVc5n3RjsD57xJTunTZ3q3+QmG4
x1tdUCPvPULI9Blc0QmEw+J+73CP3hGBKW2xnRgLqku/Mqqib9wiBW2HV7wyxPjMvpX/khJEwLPx
FhH/7YorpXWrbH9a6msiu3yPwiO9OSxjO4/Iq8OZ/tshiErb3a21iR73Tll8rkfBjI8Ar4PVk4uM
WKIkmU/nTf2TkGnS05o1Za+zMENU7bGwU9S2F9oM1D/yZ8u5jVXM6OE3W1udreOv1FcJHwi5H83h
zP7MhqJw3VECxcELtUyPR3nAMy/yskfZjedsOln0pNWBlLA3Il5noj/Gjl9YWDi2S5OrSFzBE5Cb
6zF67QC/Ymc4L0N780EgDjmVJyH7PV0q7FM8+6mtD7w4UfKym2yXWsSNGZt4MjLRFk4q6F1KASJi
W18ilyjrEq2f68xIwnBubtwHsIcs1sERbqFu3jGWAaq3L4cSfwUNGJKEG5Vh/HlOw9q4ECHkywDI
PdUfpbNwQTZ4rVSwNKVci8ewbbWN78JDmONkqxCBYBO5RSCIMCin7mR3T6muQRpD+nzRuLnNBzVQ
FCH+NJ0jrL6jWA7tN3pK0tOAVLm8nQBMBYJhnWhon2WFLh87Axt0aBm8ZJKd5xL1Mf6ZqPDMP7CO
C0t1ZwRIkGZD4GIdSPj3nn3WVwznMP0+R5lf4eN6xzkf1YWkxiTAL7Bb4WSkcQExZij5Ara5mRfU
kflMIeV4lT78tHk0U940vvjayTDnDEs2p6Cbb7cAICj5SzS1dY3gr3hKo/9PM6NIZQIyt+vnjzU4
XAXLRQkj1phbNu1SgohsZzz1prHbvo+PrL/JgKS5NDueyVJb8w9BCkgrfWeBBn/XI2E5B2am/HZZ
3BhDyMC+IODDXAgh3BB8NvWp6QZZkVB9UpqcD013aVnmYEO/0gp6yizn3Ss7bBa77iMNNs5j5MmU
BpOzTelmS6KLOHGu1ebrI/jEbpJ+FnUDhCaTtw1X3BO4Q2fRufnrCQMcf1gCYXoqqxgqjZlFZWWD
lpnDD2O5SxzV1QnSvtYFaqsk/tq3oEQoOkjmCn4R1dkvFwzdrVAGMNZm68T9LKJfgp9nR+o+W6/Y
pH13P9KAwK8QdFDD96e9/LlwC2i0bqKcH6WuNyKgw0BCkN/rDuucNHHQb/kslny4v7eSSbF/UiYJ
L/xm1XiL4Ix37Jkls4sVJcqCXvK68rt7GrnN/b6bx7sW64u066IyBqO49EuUQKmpWf4VOMxav3/6
deO2FtH7o9rAbhY1UVXoTBxntqUOxMdNrkKSqiO8K1GDHrlEv6oVygkCEU2xgVdTJUy7IzwQZdVc
XCP6xNT9lpKEGOr2SNyUiWk9bdepjagmrfaoGKM9BVRMV+4GSNBxMYuacb8TeAT2eqPi9dmtLAXl
Q9/vejISGY+b9Cdg0Yf9VzYCMy5qcNMgBRg+8gb3P5awhogPnDZ0mOECe0Vo/gadDuyKH2zehOR3
RG8FKCyB6iaj6Ahre3D9xXL6TKr1JFC8bjNUOWTuPHB0UXykqvLFAqWdlMC9rlGACkEWMMSorE2N
f3JxsIroY56IXgpd3QFAJhEikrcSHixBk6KHwc9o8uNelXA6qPUHkysNbatIiZG9Bz9oIBebI0ag
RURWCPzt3lAA6Db9f5FB9fjpk0798vIg0DO7vfZS7OemPPe4kR8eyn5V168VhitzEUUFSF+049fY
I3l12Jiyo/2BhTUu5d6GftvH+6Fhkiw3D7htp/TqO52GEWmafP5U+Mu/6L5aX2PFC9sEACt+4Fof
uXQJ/5oyVEZopbKMv8Ovbue5KnYhOK/tEIavrKqCNFJndz7O/TmOxKh0Xq8/wiCXyFueUCr4+o7b
N0Pw8mFYgJSZfnZxzRhezDe+dlEH94HMoShCsd531vP5EB8U2sOVBjuu1N+mKTfgfii1QfmPxGBg
MQtzwQ7vIyToZ5hoXjqruoVUaT8uUfKIkA7VqL33d+lC+zzuNLu5MWG7hnL1UuL/SFLZtPzTw4AD
f+2E+yzK4dEfkChz97Jfri2ksrnRSClgpIBPQd1npNO3c9GVnMUZOAUvsYHif8UZ3ewZ25nE+wwY
JPy9j+mNSE2DYpLE0HAO2tPeh18hNZoKdv7cgJ8eDB1fkzk0P64CEoFpK5SmuuJ7aLxR9xIecBjU
2nB5GQBbKRakQocSCr3TuPqQDLRs4VwPS4/w9SWKignc/aWPiHK39zJDPdt/dNsjZhsjWJ5p8acD
87xr2G7jlRsIg1Pd2U4hVsDDawkBZBan7yOFJ4rfdq/h7AeMv2At/fmrCB9ew8iu70fc++ZWxG7t
B/HCzE7B/IVzEJfEndHVzs09/lFI9k4MAZ7rsTr/WTPkDn6faGjzTGMw5YOEU03kj9+M1rWLkPh1
0myMwp8inSzszISw4NJbwYGg3W0Xilj9WV7YjAMbzPeTYnl7yrZvtlrBUa6d3szOS12+dl9OlZya
y5o5q+7l9LwwV5ykH3GbjkK/3R8vDRn/qBSmOvoC7yVcrpVVekj/vnqpRsoE2MwCkykns5h4/N4m
L/1P8u9je9MPCj9YsiCRjx+It/sUTH7vlZKHKRrPGKUNh16Ya85mSNcWuWA5DkJRo7NLA/k3AmFp
gmPrbu/14h5GSQMSNWDwbHtN5VmwVgAbkBd5NvI8erobc1XngEGrPdFMz6IhZzytdU1rctRFlMlG
Qabj1YMmoG7mEoPMhraXKAI2yoH1MYOzYvZyCCoZtZACqE96a8oiL+NMEClzbo33FWjkCZtCLboH
WxJuopHCHqoGHUW9/2qCsODqprR2r4jtUn4K2vATpfXx/DENPqShaiCHCNmENOCKbLg7d9nJqkmy
0Q9aFuLHyRNW9Oc50B8iVuRNI4Ywh8mgOCTBpLCVeuTJezJFfRH2MLy4TM6BXMhZ+VHyI5CZObEo
WGT5masmoWkKYR8g6lnDHZpoCsHPE1mW+fVIS3Q3FAYY0dvG3ZBF868nyGsZPwA1Ud32zuMzjmgf
EcRNQNYHOwZCaY2kJN500b68LGZVybTDmcRKAV3WwB13mY0RrNH5IVznJsC/R52IP2zu3ixSgXR0
WUnOsWl44G3yzg2g5YcG/roqmbGn40flGovpqg8dYDc7vbiYYgMpYhR/60moOZ8Jikv3EgebM+pU
fdz5+RHg7ngpolK7yPYDXFIpPte5sZmxvIG22ycqvY7eJWMmFDheDBdO8adxeA2NZ/tGWD2tWdAd
rPHOqGE+imq2d2jVUx0iEmMiTv7caaGqrKz7IfGgncuQhCGltDzBDjsSeIJbAO6WiMfeSvWcnjDl
XC8IojPSdlnPEarULBnYN8+yiePW2SY7xDgK7WTL4TuvUCMOfOIEsfKrGUmgC0ASLktX6dKE/pvN
6xwlMkXZtgdV6ZmcKKEOG07Kp9PQTRCBpUog58w+YDyzQ+ZyucGIu+CHPwymLh7kguvsL64Sfgxa
jYbdAFdLLuQTHZIcDwN+Cd6c13vwG0jZy4n3JoWC8NDuyna7RK7Yw6DpWORKJSDhfzMzrvCk0g1b
kHGHXmInUCX+LJzs5F3ECcO4mQ3p9wAoCBZnS0EgouO4lGT8zhH7Gn73ye3yPsh8C8ybUfmOsccs
Bx1MvoQKlbvUx1rR7n4anbXRId+0dzW4ZwAoy/ICwugqeaIACbHVyH22Xq2VOTuGWfF7MKXIimap
QXsxPhJiZNnPm67kAuQ9zBlKTwRp8QVYHvAAeG6dSd2aFelIbWrwLYq8rLb4cXuauWYzGtNmdGBu
33YVOVLIwfpBwBtDzyHFhw1HTkpmhVI1/1TTLX/E7NVy/7o3vEILIvnSfrJtAQ++ylw7092HgLzN
HeubsR5/vQMPtISeOAXLSVIiJNzdZaa985CvQmq8z8YbX3PurYPNoLPLVcGQ+tWLxV3aoLr2z9h1
kMjmUcZzd8UnaL3PNcHC7YfuGmDtgznaD5Tw9eJOxGOESz4l7j58KcE94uDC866WQ7IUfi2KMoUB
LkXAue56rGUd30OnOrqnYqVYrJyD3vZKRcrX4q96EcPjhcUBgKW5iP2cdxnaqMnzWYfbXAccRTIQ
yundlObHjfR4Kfuu4BMvATxnHOL3Ibg5n+74bqVSOXlFDwlSAsOy5Xueud6SHgdNDIR3hjEI8y4v
aQWnORV5fGrI4QjMm0TRYsnJaENvLv/k/b9AvXQWzFVzRaeOf9wNyre8KIIwYQz7Ux4yynzU7mKA
BF7ER4aS+zdq7Ik6q11X3Ykq/ylC4HX7qUK1NKzczKi2pxTIFvM3qrWPriZNeipASqlWJ6wxNOlz
+5K/WQMnEMEVFb/owsf0+ZivX2CqY1q1ey9sSA7U1grUFjfJmmKKEukA23XMJQWo4v5e7Smzty6a
wEUVsiKX/oLBqa9/BXhlSc4wRFiRpKYVCMxNGjIaUoMQqFYSIe9Q1tVdhL7RCjkQahS10lPnRaXT
0RS5dfEhmM7K57V46XD/s/vr9xaJY5qFKCZRvQrMZUTlUqmxus1+3xxdCqAcN4QmO7pcopf3S4Y5
QCJeayF1a/dONJ9tqpQv+AYHbch/wBK2G2RW/QmCf6zYUA9Al48FSEwHhteSg7wQoRwlhcD2rkDK
4T5sv9z6UlnrYMQBoF0LaHs0YNG5ZRbl3YLY9IDkiyydtm7nMwZuXDxz1gifzfJmZDW9ulVh/h/c
1b3AhTimf/4UL379oYTEaTvgPg1OYIr1/cUw3jAJWghAjJJAdF3ZGwtDYrYVGI+e1Nj0UZtFRG++
gzqe+azxADt7Nbkk48jggfgGqQf9NaWBkhvzUZVFp3oY46ZO8ZZeWDk/kzdlZOPj3Y/4253g6muw
e15xv/5xv0+a64x8jz+NcOrhOYwxDOgmo/M1AOmsVO3p+OitK18PnZSdtbJzIdw+qOHHfsHZy1gE
8t0iCJFvpvwmEZ2m8nF+Qua3gzKIED0olNJnw6BgE7A6/BLbl22YNs6HQEbXNiVh4luIIPmxA86x
BDrhmPbyR/GeL3C7NJ0RbCAfII4dcOuRmMqUilnXx3oj/Ha4UpD2KR34ttDpZP7bcKKti1vN9NNo
IomrWF93e2YcR334MbQQ9vw3k2nr+O5vvoQEmoiYKvhjHGd2SdCzkH+TwWMgE9ZTZ7PCIsSfo+FG
fKIKRQJ4lSs91dl7yVc8YFWJbyT19KYi/jO4JHniGsOqkm8eF2nmy/0PMEvZMy7ewL6TCmI0F05u
qJ/5Y1MES03DcaGEN9Vnrjdm55v0o3QsEX4ag7ZUGaPtm9mc98XM0dXnYkxFBFKxPjn1yyeYIK9V
70+vgX8T3c+b2RFuyTfynrhT6rulNGMnLlIZIAzdLjnPW8uhcoN5mICSTXtw2Ae0SxfoaxksgJqQ
dVuXqgnBRWmsRS1XOf6RIHEN7TjDuGXrNOMuPrA2tJ0Yls67Pm/wibrnq1j2UYYqimkR0bdAxUsU
kXWa1phKMAWAYPA+PoL8g4IbcmdBnOZD4CMddszGZlLLxn//JPNmoMD6soPlNo7K9rn/g7uQyXFa
/CXgOkWFcX+7SzsXNQYQ3i6I1kiJWdxrRS7ruSLedDPwXAYUIqZ5vS+/xiNJw8kq1kbDEVf50hjy
Xluh4ZBFGtykRC1gsmbD2nHQ/VgcCVmj0TSy/nAfdQ+kiPLQSy94QblAqfUInzvab89PngNRqR+V
TCT4nwlrtY9xp5sX/LLgmcC1vxL7d+r/sXcjCrQJFwAa45yV8NMd5k3/LoyPUDdrDtaVPhEH7Dg/
yAIbArhzSfXo1O2rmmmesxQPw6U74yt6DmeTuAi1iaORCTB+TXYA4hxXnijK1rE7nEU0erTv8thk
9VmkMXEB7ZNT/s5Gq3zMZ1/1bS4fgFl0LcrW5HjDn/gdSXNGSKGZyhpjtsbubPpJCdVumtfhEB+H
bxASLezD1qWL2EJnQz54DD0oSEDeykPvpJc3RHz8BBKDMZ/Ld1DiMQmXwv3RKhE3uiaaaR9deDNO
aje1KkxV3JqS4eWLg3GCDx4YPuBSvj1/LxwfjYSK7OioqKcdh9yX/fpXy/S4K8yC/jXNsTlgoiEM
8PvrQ7dlP49fW1xx6tXXui+yg6xEwnHSPExw/5bpyXo99D+irL3KQ2r5tA+zw9Pm5DCiClITOSL4
fd+DBoKBE/oJY6tL8KnKov8JS+rKG7FNi6Ck7pxAjXWwq5WazstZGH2LpA09i4s71KsQrinhw3mf
4DUQuxlICzeqMdK+Hn40NqFXQ52SXN1y6OXWdK3P49KzrrubsrU7XzN4yrVgnQcqfUV3bv0YUT+W
JpcXY8p+vA3ECezLJgyJBob6YSiuSsFX7xaR+EA/mBlDvIIfwzk4kfjq7aD/hujkbL5SlXJgtHqu
IfZabK+lf1+9WVxeR96Azg0DULeAP+s6hm5mh/ljR2Fp8qbagwT1aNTgXb7WyPs3oZ+1wMvGJbp+
FpebdMrOa2wI+F1UilPoGDF91uHxPxk4/9Axq7pIKC/BDUE1DELe3wdvXmCq0oCikNoyUa3DZgel
O71Om/1kU3Q6NJx7myUuEQX+lsrZfnxd73n0Yzs5lfd0OZDMddu76eYRnH2L8JrjLWZBUyRhfLaj
ARaSWnXHK9d4wnGylYK4mK/QO6up7i5wKZU6fPUbSIXBnLFcG49GmOmJ3drRGF5ey9tXWxm8OTxv
SHPNScZERV6zzfnMcfLezZAfPx7D0tLNcW/wGRfGTrUzoVCp7RV9G3QGYWqNKWSjLvGfGGj1eWtk
XroM5+LF8zYgwjfyh5WjVOwhxNGZ8NqAEfx6lZlN9KH/kibqG6InhpXqLhuF7PWLn3qcFaGW3ucd
LTOBR0GaMPpLvo1QXfUI2OD45d7KAJDSrFKfga7hJdQ9fJJFpP+Dk/2jejHh8blZTThA3Ph8whyW
McgGwbvsJBMeDU9VbOkcjxjSOUF0N+Ud6TYTv9bytwcDB8ueylcpdSIWooOaMtIDnZqF9HlUv3jM
TuFjBkFVAcEeO2Hrh1Ao9yYxAvCsPEyJyz1Cxu/zEC0Fpd+Ks4DIbp1ct4RGLO+WOGIWyePJy25f
ptjVw2CYfl+w2Lh4AotaGiNYihS8E1P5uQSVXrITeJNRev3WuO/3MRYfc+HlFS77mxSj0IdXXlTy
x9JBfEqaIU4v8+bs7121FQwhM2tk2mDqvTlJPJUifQ8eWiDW/GzrAUBQRKvD1eZOGasqC1VR7/o9
gWjsRk7wGVWeCC4AzhuixgUOgpdQrlMv5L0ffKvROEFrzsQYgZGTcwWAMIVePlFFb+oP7YCSv2C5
zLgaZ5M4M30k4H6bYRH4zbVlDNCbpR0wyJXRafBmTlWbZuJzKg5twzy6IrwWzp+7Gh3/JSt+dOzt
zFiuV4rn/hBzPIEcN8UvoH6Bn3JJUhdElc4RlE0JvbV1jAzypsPJNu9I41D888S/rGtuThMa5LDJ
ZeD6GMianc6wAO9ocZAgFtiffobb0YOq3Fsq+mJnl+Ly1jdyAUR5wa4Qh9tx18L1BrrlpWWaWBc3
GZUr0YX5TGVIgkDr6qUrsZnpPXKpSCralqkCW7XG+NMr6yOY2tSz5prt2egn+srIc749Lx+8UERJ
dknViX66wKj5nnjm2G6qcWKeTwqvtzV51YAZtxLxYfsD4FZs2465ZZhJC4Djkt5/znHydlty6t6I
F09QL3KSFfS5Ur3i5GLqgdYg8zQjIOMZuFnBOyhmadTkR/QCddPXpRZ12aA+IB9/DCf7WZtB40bk
0kshYmM/Mx+u6A3IsdYxdu4ewztevI8E5KNNj7jGY1TLwELK1b3ofDy4mkHiZU+p2f0c2XXEggQg
9ENHUk3VW12eb2TuXTo8VuimAPgN5XKo8GbbvxCFNfbJoiipix26ZttRyDsCk3zx/NhRyPw/kVFZ
8nN7Ui3rR/mJOzFMtxZWQRFqWYoWOxxZ22JuyB2qRIQxx/t7GIDR6tZvwL6MSsS4DRGwAIEpJTHG
0vXUl1XquUKQEz1vau1bp4NDvpz4RVLi9XU/9OaQf4NBHlYcfR1bMKncStSg0TwMWO68YIyw6McP
l4ZrgyRzZYV4vDst9ZhQi6lQh+QPGqI9OV7NstvuGSjzI4YgUh8ikXY10A75HuvgZaUpMomVte9c
cGlz6P3SqfInraMGqicd7vjd4tPa4sGAK61bMVTmacJx1sWve+OfBxdiUdwa172baSSaPen0fyIg
5642bqXkvs1bOk6ucxirLW54LwmmfIib9Xv+nwR7rCYTQtaV8igBJoBmfKzp6oMOtZvc2u0vk70S
0TyKHiY48/zXxmRX8R6PIP9v0xA/MxchPat5WUaC/5HIZYUrvHtoFMc6fGcgyMJLNURN+Sfmy6vD
iVYtvYusXMWTNbc497fqeza2T37AeOnVIkNrgzZUNeFWwGc/26c7NXPNe/5IQZq+zVj+4pN+rV1m
LgZbD/VAv3uObk50w7AHxuqg4tOjHjb9DBR1KTCkVyUb7v8OhaISLssbNB1KYSFeum4Og9aZQfP6
lHkbs6bW5vYgoQre1nGEZlnVNaVy4zU7D+OPE+q7GNCC9ewFAAadntdTKMDRW/hWbsnU+lxYKaLS
LfSPz1Ak3Nj7uklaBIwQHjJG10f6T1/ugX8CaKbgN36m1vWFKrrt43HkMV6tfBMLXqkb8l9W/qQ2
zI0lq9iQA0YNfUXSZNZIg4852GskhWQ8l7odJfynuxSPja7lGsyAXzOYfl/HH8pTz/IQzz2YIVc/
UdzIvd6XOLcHYut/G44gfMb+nJEXDpYEBWSXOJFItgCnzpLB960IIgDJSBqoY1Pe0b+uGfKxqgz6
H2hfhIticUvGTcSXlqDnI9jvevI8tAOexUd7KLPftWRJ2sV5gs/FUGRyT4q18SeyxtHlOE0w7GSh
wpLq32hEhBR39hGojlGhvxG55MovKJNaILFNVQ7ymMKhL/C1ZnfOaJtoIJrUQorTCHYtv5ziGIXl
KxBXeGX6NdxyODSBqBD9/QhIa9rAOEuJIy2x04PNNhBO2YNH3LgbZZUFWhTxOKA4/5DwnbEdHiLA
HGLDzY4Lgr4fB/JIPWf0MFdruPebG3GulJdAnLYY8dlb5NGSKDo9Ucn/l0cNcft/oqCUBRWLsDHX
R/piq7TNlWlWMDAuEhVObQa40thbKy0Yr/TiY96bZ5uRywFOq9kmRwBU3tKBwJih168pRT1Hsw/b
WJslTK+VgUvJhuMD3hRYCZKjH4+YsmNXIvl6XaATV/hsyeg2j1c9V4JwdFlwT//FOggPRK5s+b22
NDFFXco+s/Z3+eE3kDs+piyZNMTmIvIvUyQ5UZfJ35GJHVy2w75m6XYFp1lBG75IA8ajch4tuCFE
qVRXa43Tjq2p/2kFMmJtG4Coq4XZkZT+JD3cKzQjLmIHRGVq1QV1U7rcim5gX0vXBb6ARGlPguiU
HwmCIx1XIPqO4lMJM8Zq+WWcf/AzkAJS66z82FsHO9866Z6DyYYe1hhs4uPKorzS4yP3d7Gwk0TR
+ykdYCQpAhHaWzGJm00pFypwoQxlRsQiMuYNX3tvixlEAegVhJW6R7QW4qk+vvo4cnEavpILOQF0
PtHJIR6a/fll25SFY/8uHIklN0KccHWnMTp8skEnQ47FqoQb9+Exuh8doY6F4CsdwjzrdyKZypv7
CaE8qadGJ+DZhURYGWv7VirhNsfa29AIQtMedN1hQwHLehGOiOv1rWVNlNZdS14b1iAKx6WR6o7D
gthfHAKfgM54DfXeVhJip9R7BXTFPiyvisICVloRosICbXDlGr9WKvQuZfmQIFT2Y1dOgnCdBnSH
jCFOUr5N5ntS+VCaN1m11ksq4o6GSrFogmnhMMTQxWEDw3o2TkvmCcK/osbgDENaNQMiPz9vWJ6q
FI7C0gFVSNeuRyjA5WqkSWptyr5rpR4liNbdHWu5+RbCfHa6V6ROBDJg42uLCqLHjK4CPSnWPvcI
uXoM1SMB+7XSCQnN5LpKqqUwpv3rQEqbyDV7yg/GC7kMNJrYgzX1bl8Ki+wEyEdb4zWypGktEwJq
J/yMQg1F3HSmR9Ls/c/kIbuE89S2Lvl1twuw1BK2BtOIeW2XlsYcJjkfkKgrH5lgG24MOReNhWUb
O+uqIFDB7hBADS/89kxqQH/+7k6WNo9pknl7JERhP1sApdyTdnE3QVMtRyQEY1H+janrFOnaxoRF
W3jm9Ylks++jiN9kS/eVuzpzShU4Mz3zSfqJ76QYepo96lTgUm6N2XyKKj5C5UhhbLETRZtag4+d
EgibhdS/hekQS3ziIahmM29Zyqe3ytOWGOh1BUScphBtqVKVjra8IzLWrGR6QJp+3rwDnF5fUH7a
5mKBv42Rs2TYtk1smCXcRFvpAys1GnaWN1ILyoOy8I9t37xKd5ri0WPoztg2qaVp1oq1ZndIRRgg
dID144Q6EDquw0DTu2G3AxgCD9oXP3LgR2LndaHKxZHM/eFBtiKts9exIJeBVR90QZM0ua5fuqkC
rc8+0oV89vu4hkoccecMCoizCKLj3cUzctxFDNDf2O6+IxD8ieFToDizIFXpkQKrMaNTrSEKJ36n
zM/pvgIT/NEctw49YlVw6SauXqXx0uGj5fsgHBNuWKAaH6NT7wbsTSqbo8JX3mz/u8egbA4ts+Es
lfD32AmQ+Icu1+KPA5Nkx3xjIlT7x3wO163RCF76InhYk0GXvlqFBzmquh2/ng3tB+LIcIw188Ke
pxe7NkZs7R8Yayx4b7v8ckFe7HfG33n/xRuGK2vPYOWlvy71p09lerLcu2SaBlJPX1WFALEP505Z
+IJO122hjY7iHQryxV39fmzhzWP0tAqlaakm4Jdzq6TBg/ulFP6nZrSXLsGp7fEIz3NvjCdleVlO
bFr/rkyY43lh5pVtNZp9qfPNXD+6kY70GrGPeODs4QbLaMBFb1q0YQ28HQ8P7OvPvs6K8abx8zE5
1xpFLQsnXzL2hbPCL0hIXW1tF6Z5uJjVzQvH2vrH1QbwvuYzr0nnIAhexzPwXIQvzAd64yVtPldv
fZWzZoFt1Ipgq7x7P5V3xi86aK249AmtZjue0gPyA0Vf1yZt3tgzgZK0e4u2KC8KcYZ2P3F9a3PF
csyLiZOAZTtwnIxn/NdrZNhgEg2p1CuwUZvk05AHdOV6AO2tQP53TsSN4CvqH+/b5GUnsnxfIqCd
5BJITQxEUXuf9vU/fsEThIheybNR8puEzgppyRFoCzz1W8W/i+v9gtK1uUa4J5OtRRbL0epctWW8
nioj56iZFZtMRKexZqQWTGCTGSjzLVoPaO2z/4jRpr1Kwk/f7bqV9WI6Ps2Nhsui5gWxDb0x5EXS
nB+HcE31gRwsRne8PtsScTunaBFcb+GadLIrAbvbi84qO5ns7NDjlTXseAFmS1SXJ+Mt9lLxLJux
lQh/KVORvj66dXefdyvJhMGwW4ztsCj8PB2iZLe1i7QYic8CNDB2wkFYor+awKTCSKqLCfEdCo8a
MdoohIX2s4Bq/1Yk2HVFgMS/FUKtwQB0AV4YcAeMRVrL2GabTpyB2Sgqc/sqmu0PvmLInDFvjbI7
gm475TLLYI1tw0NSA7CZROQ0eNBNhDQpVxxSp7lSSFL7oO83AlFRJU/uv1PL8E+X1I8ylpPjMLEN
UUAP4AgknGXpbYo4QjPaO0NP3okGqwfeqP3tNQe/v/gEf8ZAe2ymYYtPEgj7wAccT5h5Nr42IybF
MQS5ofkwJwavT/7XFVlsUL33wZIjzG+R7WWpYzVCeaHK0wnF8UIUZ+Rbt+Uu0GvI8Ej0X5xnWtAj
yWR5t7KIxdUVriMTL9B+5tr6EaRSqZa7CZDtUpnG1lM/GYlD09jMQublulz/7r4Tp8Pni8AOxzaR
C2NfKhwVo7zp6t5pYYd5fQpA3DBxPzptVgvM/aLiM/alYeoSkH6fVadVmMA7yIY8P5rXE0/H8s7/
S7hywspImxwLkhr4y+LaOwfR/A0KFbyjU1nvcGRv7pYxALpNmrg7x/I6Xia46WONUXpi5++UvD41
bZzOaKhc25x09t6WEwJlLBAPdyi7lq7CIzpwwcKhVj+uulnyTokK0Zs7IN56am76cRccId+OSr+n
sfAN5w5Npl7fe7uLfYw1jOgTV0wd6tphTJgvTmQnDYCBd/dkdyF+/oVgEC87jHkQQZY7lZwhO92j
UW/Nb2bUYy/wFTIofXmqO2qImTWXB9yKVAIY41jyt72Rg2uUf+Ai7wW7kRAgHnJXwlaWxuhpZMAx
FgNucNtoSu+RzwnX4QLYoI4Jnq1xPbTVCQbOWfY/6t8c9rA/wV0gkFFKv2RcgChnwVu3DQyNKuWz
MBh/bu30cTV/T+O8Cew0yE2f49/YpFQDFGo+mazvAKOnXGeD+YOWcz8L1iVhEruvHMbmgug0r9C4
XXMJ9yHgw0hX0dOmZC8Gp9pWCej21tVcENCtmuoqqbcpWvFQZqlXIJsM27pcrJgbof4X1i2E2lZ8
hYmMkHrnpbIv7JhQcRZI+Qb9sl1ZWOq6Z0I0fGHffVtrYPIG7bKOnlvdab+t2jJ4iL5y+NVzES3i
hqUgr8n5UHUozsVFIIJVjqFUipgz9JOvfhF+AvgBdlexo/OfpuXGiGbmFS6//KOC6NeP9G/wfdoD
0LvAZapLo8LgvwWX9yP2qBXLJ2grZLOqh4R2ES1LRzGJChu0i7sR6TH9Fsnwg+5IwiHo8+/AZxoq
804Mrtz+HifzcpRb8HcPuUf4MRr/3L4kTBch2yRT4wvbTri1V19j3LHN97NNMQvzth1MAnT063+O
1f5g+OC09n7XNVuHrD89Qcx7O5+mb+4GlaH/i0f64lkwNJBVYd2EAZSsGKBuvZ9J3f5GqvZZ4gdU
+P+AHu+o3MtZRNwUOHB6eh87JO2zhoa2Xcd2EnX5BTu4GI4v0+LYU8gLADalJ9sAu0XuGMZwLbVX
cR/5hxK3YZVNfBp7qvK2M0p0pBCKeUnuYKZVD+ALtKuuZxrxwafEiJc9csEqptVF2wM8nprLoyqm
rVAJI8QLoZ5QUqd5/OKFrfP/0D54qVJdWRlzQWQmpN8lneLb94o8meJ8Vfni//FaQMV7gchJLrQX
DwHsQvAXD9h3OFZ2uwAz7DmuzW5mGygxmsEFbk9qBmaE3nkinaDOzJN9LlTuM90QL3/Z4qA39mNP
h/TQE1hrkDVfoY5JNcmLHjBenIEvUs8sxNW+RtK7oDGaquLA9NS4xHOyIDHqTyZGZaAiEVk+Km2r
wJ5NpnaKvej48SoZvJmTzkGilRU5X2GMMoFKfmsqN2EtlMsVX9RhXmEvh/19F+9TNR/4TPcyOH5n
pwJAngowmc7qwYqfc7vJa1+uKszAwsHxnlPd9tOCX6VSy95WEVhTa6CA+P2sXVhu+lWDL7H9URJc
3wd7eVwZ/98krcG8BMyiLZeLqbuDK0AuOFw9+KN31ZcRTSsApzVo9XCmra/AAcTWOe7lXVa/X2ZM
+BBYCyjMFW9wTFwt3R0qEJl/HmrzugFjN51WX5YJxVSE5Zu2B00C+rTt+fRneErmgBrhfCVuRfK9
tv1l8/atZ1Rfqn7YgrO8Lm+PJcbJRuZLv1VdJlZ1t5FBmwDsNrO2bdLr5HyF8B+BUtGV2UOgLc4H
kbAeiX2IWgkX4h7o1wT589tKAsoqvhW0xSkLQztTqR1Bek7RIeiA59wXARAT0jljjS/5ZqAdOdnI
nveq52N/BAMWTiCTgha1aOQ7mxzjspjbKMF8KHrwyEspDYe9xYWNDXxPFBDFz470O38JS1ozihYk
AFpkNarZqUvjILcsMURfwjwXH3ob4U056Aux/Jx15Q1P6AH0TS3KPjCPfCbfuj6OXAMqaWwsi9Ly
/RgS5/OgKjrgTcOaUG7oqVOlyO/zpdww0P9SUiaV3GFBmy8DKrBgQ8BIMoQJCGmG36POuZaweZlt
H7DKVfPbBaVfOsvQv6v2EtyhM8OHzd5l+mQWdXvJnEvVXY4x9jvhuUqVJwzm1HjidqGG5Je680lG
XZdDzqZjlysrVjO1a+VUabTN5yKNbnowlozK9bc8p3xHj2Ro6ZLLSH/d4iwNsk3/hOjQ1Y5HokgM
18qiL6V0Mzzr8Kl7WxLi+7+2MMeNuicJmKizx7sPnjYjOc9i8Ua+nCvD68o+SOQfwArb8b/47FHZ
ScSWm9iDDgN0maVO34p7t7E3cvL+gqnNzW6uBzUGtbhcJgDPtdlQ0G52bNg4lP8hvbab/bs8a/Iy
tRM+plpg73X7QivK1pik9WyqxH3CAiT2IHrR0fCokQtRk26yrVAORzZxBGWSsp9b7eZFhjfu4bVr
8k6Q4Dgzt+l2852P5ImReX7D2236vX2/zfMhdBgZQGVbM9aum8N5f1VuL4yrd55CtjQ8lEQIx2If
jDDrrgvZUjWM/hDnK0CbxuFrTCL1rtJb8bn/0QptCrcoWu6QO9t8EacZPZKsg1RjnE6EjKTYSMc7
YwtUp1bBujP3/BAN7S/ix59dBM5Dz6ZZR+DVQBVcblteMmqtBZ7/hq1Ok12b5en1leynkT6Ib8yT
XQLMmJxTDblCKnmtV/gIlxnDSihckdUtuFHuT9K/5E0tCbys4GDmfYBq6HBcaFvkiApeDPVqtAYL
PIUFkEGItVSCi4tzi3B6vkKouuP3tj9ODumnN0HA5fFcoXoe0yDCnCrMwJy9tqrgoWIxv+5MBR9Q
vcz2hDJgfGpmwMz6TzXzy78c0k2KztRvjaWPqcW6Q55C5MZbgfnQ5fVE5+RZ34FX2RTnA9Uy4Wkl
aA6qeY79N47D3IgFzwLwjuoqFdq3XdxbL8BX32ChDMprdcndP9d+GnPW4HHw+yDtLbZRfDAAytT8
WNC6wHVI5G/VJByz5aHpJAVpQ199E91z0m5kCBqYyalv4G4M6r6yvj1C3l6/ZnDcaibugchyIaMV
Rsf3SmSrO3QTe9jdpYqoNr79JDVJt0WNq+LtbHHh6J7if95RemTU8gfJrEJm9LCqBs9rtkdYee9u
HJTOWUyF7p+EilfzpqarqW9rxKh0pZkaH5Bz+ODvx6eufsZdEvWlIBVut4L09Z5JdsX3BBdIoyvk
n5JSebxPZaoX5Cb5zD0xaPxOEqdy6Qa1SbuT5IE/3sK0pxAlcAeNUrNo0eBKtjfWPPnQEv40yJvI
nBaipSlgBuhPv1pGfL5Qd/W5laPTCD6nYruSK3ZjWouYmJEHB5CfyLVjg13nrp/AY6fQLIsbvsk3
8GKrJPUDyQW82n6DMm0b4VwR5xClLU5B2Cr7IRAJiNR0JI6ABqHOe1PLkRFEFA/nvxZ0TVk1W5u7
2cG2tWakQae74D+jAduVX5UJATQ9j7c4d264geVNPmeyuakT9g5ao1P2BfwDLVmTRWnxPzWca/0y
CfUO5Hh53ZqrUnzitSqTjviQqX1kHZztXqnsXQFPtzS7MOoOh+tFoBJPhsGD+fjA6kz/9DXPe7Lq
+EJQkCifmCCTFHPUzOYR/soZ4k2x1XYkn4j+5QdESZVF4gPZqz0c23rq+ImY9m0/riQe5fA9VTO4
uabPJtCBqzxAySkOS5E6n0BVBOc6OXi+tMizP+rRnTR0zSu/AXEqW1+OOm3RtLrt5Jm+AtaoVfdQ
xKw3P+pqZb2LjE7mbDFbifojyuQNwqAAjBBbWZE/eUzyCPHEYbYw2M0pye4aU2gCldPucZ3CMnxT
pT4PXBmISHAMD5UFOn2XHwxVofDuK/ujTYYhLnkP5X6dZUi5mLd5TlViGoFrkpd6XuTYk9DUKoFJ
ZyOTpc2tbbZ35V22jhUDyjYQ9PT0nHYBxSKmvNhTCYkrWD0So8QD8PYUhOkYYQ93R9A9egXqe5MU
aeCFnoZ4D/3zVsFNM8ZvJPjQ6eCY+GsGzX3C8kWaRJDaQ5hJypfBRVTZIxFNandZEgq1jlmbJqX6
+jH1B18UtBA814YGX+65JiVLTJMslXRQdQoK9F0/VPAQL95hCbK9P8B+SDmS74gkOD4hUBH/Owpv
phmigjjYb8MnmfO5cfyxI5x7U3zdCLJ5Qy/rGdC+Onvyhfc1lmT/avxlHjsU6TOLYV2HEOalJl5t
6U7DktB6wtKNeTj34bgh+/pvN60zSUC0eo95/RUZSBVZvhLbz4k7Lgo9r4U99VtybQZqxJm+WcZu
ls14FfbvItZK8PVUvDNEkZtjY6Ofd1NLin51wiIJksj0ccLeMMrXJmAo6i/HO11HW0lAx1Wq86as
tVAmMsC4H7Aeb+nNOzj65UmQzAUhO+cRKHfTcyvirv6pUAnMvfLPed4b8+9JlcF+1cCBiH+Wgz5S
6CH9jx3qXnpMgdFWvjUpIWCdcoaZK1xul4BHdz6KoLc3MzFZVlyVnoah7/17ZKYad/X+AZxQTyGp
DOJgOxXCE9lXu9nGqXp88MfHtYJr1lPxEb3Fxj1NaYuuILwEi3sCmi9tm39Dq4PmD5slzy2aMjIg
gQ/PuK+jF8AyZpbDfJL4vQzVmnsgVjg3kgvl/XbVGLHwI5+1fIHoAmP4b2UVK8J9534590LlfYkB
2jODy7yCBvwF+cThDPBZyPFlseu3JIunhH2hQWbw7cgSDS1hAD8fRaoJwCr9aT/e5cihYgWX1M2N
dBXrIDiY3ubODY38eypNr3CU9diAnExdQE7hAic8KLBqHso2C1pzN5IBxEzr5FZR2+aqkbhDxRqd
axa+auUhwrhsfsr5X9lEu4XwYBi19NCS1ZB3YttR7l6zZfDmJA3121U3z8qI8tlmYlCUfLUFqhMt
27b7QkDrK0YFV0zi6JOLKMHvAMNzLbN5MFn4QHY56Ufw7WSXPgD6Yc34o2gmiibBbmNGwUFsX1iD
flxY3wUVvR/yuVPInoSTKTq82+6agrr57k0+PSO2w1jznkbcZPJevsonm6o3xvue9VysATH/ls1H
ncuXCDkq1rkTJUAzwdIsGBw/8unaGuvKQct01OwD4VhSVxXZPmpFryUBNWEVTwOirYlUmCOS5Mwf
D59qI2uxA52rg3qg8oL+FCO+EYaxOgnGnhUtacHmIucbvW/+b6yj8VUsdLieJjIRwhi7fOVrjJCT
PyxCF7QxYlq9VB9cRfWu3qhK40pb80Zro6TnRe3FZlbRK3j8YpIuTIrypkPHz1hGe3wiafAGA4ab
tsR+IRi0E9FmvEhOtwsoh/gi4mt8QoQQ0uh0Id7XRU2YZVoxMfiW4/kNeQOt7VZjTaWL4Id3rsdC
DXf9TApIW/DJPuUbqQShuvIenrj6KCiqWtpJT4+cs/6bVI1XPYTqqXoIM+iR8mAbwvf3NMNz03fO
xa155ARhYq/7pH/o5U72B2Uo7MmMRwH67jnoAGiIbZO3eL/Wpgs56MY0B4KmGudQlTLvfIfAsp9D
K6CsqgyECRZEkDbmL2vAQgJl3fEfq6d34qIgrcvZEe7SCZsWi+ZMqpotTFl3zKZLfEtlYexlj22X
WoJW9mf3KxBFrBIvDNM4E/CwuKlijMO0ZsPiwYxjOlAbr0zhYgLQbJOMAB8+n36svqntJRZZtnod
Hmbw78HOjR9pjFKLr5S5hwl75vEJ+iGkcc5wWevyGJD6v+nZv8nIa9b/g3cRbt+fme+5vjRa/p+R
xRVOV77CoB+CN/KiqCL/0aAfoEbJwLZ23Bhf88jlFnFLApipfbV5qcxbqxBfTGTq59fS8EBI6IOj
avYh4Z2TamlFT/XcUk3s/PGo5SrFKUo7zCzHR5efwNO0aOlPVfFbfKlm+0MhxSbYVyqog8lz0eMb
zi6C7THG5+ecBRpFqhRQ9DdTz8s35HPQ+F8k4E+C/vNZT/swQWwTHJ5xt8ABf7bT4tdSM3Cml4pK
o7a/VdVMrszdQ/xvE1qhGDLWkphZOVNZqdzCHps9Sc5uBhbO2l/HFs4f+pRalKWvdNPhyJ88fcUU
sw93SFE7OjRzDYbBZdImZJwvgR2llIEeovgETrZc5rps9PP5Qz1FyO7A5SCv/T1a2B6nHG7C2XPL
UiIvqvEnoJJApwXlJXSferDZwGoyFgJFEyjp/qX6O8leTSplDw8Jz2tTbm9sUl7dXZjOnb1Vv7Jj
O1tCzg4E35x/OxvWAafxZX+vlLTPT/mDVRmTMLnb25//ekf3FqAJmJyNlNObQbfH46/cJ3AfkNwO
05gXKgfd2oUABQK0tZXmU57cEjutx9mu/z+kHax03FA2kYGPdyBYzMy5Q/yYZ0hYtGto9wN1k9CG
k3wz6B8IGk21VFDy4STHhhm7RI3kv/pnnMqgMYu70aoHEGGcAo5NnYL72n/im0Cfx4xnHNYbrwnZ
kUbmohXO9gKzgkY/GZxiVrui20vXZ13SekBfjtzRLW3s8mU1+xwyE2Alv0wYUJUr8kq/Dx1XWPkC
6vXIOxxIPvdbgALneSXyPusoxbWIXF2NlZjL7pzz/eRBfQxAw9FKH9mM+qxqMY2/N2+DxAtpqZjn
Mo7zRl1aQvKCk6JDsFXgN4J6FgxcZbc0M5GKUG+nTRDzGxPzFBOCVBZjrnnBkBCAhalZz3PAjhg5
5VHQXRBBW0FTPbskpx1PLVJwCXQAihcI8AtoUxlk7uAX/u/7FioHm0Uuqr7YlQ3lu9/VN8GFsNhw
Th2w4gvuBZX3tq8zsXv8B4DrcQo6PjHCvKJCfvkhtK9gnhZmxuNdygY0pJX2Z+sAQk17U7SeKffh
rLLh0Zzx5HFL8oHaSykeCRPGVbbkjC4x6FP3SAMvIiEJLp07AEKhTg+CbMIfham9TQPGSsl8DDxT
S1JZclnLuG4mfbJ3opJjlBautG9GQVSpJSsII0wffkncJH1Fi0QXBbiE3K8uxWieKNNiaMpTd4E7
hDev7fDM+S6GML37tdE63OBKlTS2VApFYVNnn9E8tGpxyQjZHj76i5Md2l9aTU1Li6XTMa0yx1Pb
/HeYeXvX05MPE8bq1669meXT0FpDLmkshCNicLe5CyeRemeCAapY2MmunQ8GbsuWMV1sMdCnE5aU
N81JWk7D2hdfAByJfUHml4hytHTr0KnnLQYCghCIqjwemV041Wbwp92zbbSb8GbplPrGmrYns9tR
vylxbFPU7N5UKR6bfzMCK2DTd3v+3+HGvAUfzsLNxK1eiKMZbSA71dUkpt7fzKXi6SsqGc1HnkBj
UHaratXyKJwFqxbG+KwpkCGTZQrN+JYxci8yIHiHNwhHauzb4GxtbAhAgOg8Y+v4SgcyaMiltVKv
lJ+CcKmVjT2mRWihP6+kelUXuEDe7H9vXQmRxS3+zs9Bg5OiRUhYMWdz+9KhVl/InDaN+VbjNZGn
4LzUd58t7XnQO7S/NHNlvNOfNDxhq07cxEPTNNlpj7msWUo+w+XVH2NvyeO3czAsH8yUziS2wI2I
ncd6QVMGYWTELtS+MfIBTHz57NL4jO2tX3dh6zAcc7p2ZCn+SNz+BfeMNazOBdrVOdrPgeaMdSfO
56bjdFgSZUtfnTN8FX1Sfh03S6XFTPJdMuDPz3htnY4EJkkfmdIKHgfm8hren14U5LLuhurK/IBC
mPZhd112l7u22+g/GWpncJ/H7+HX9KjVrKuMKM1/XydpSg==
`protect end_protected
