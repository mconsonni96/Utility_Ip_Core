`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
G/zJkWYKyYzRjvV28D8WQdwTcW1EspymSGHk87wes2VfTZ6VwYjTsMfyVAlYui4TEhxAvNe/jidp
axtlVJDzaxX9oI+IX89GjDOn572TroGXE9yNq4EOk/YtUke13yGUS1taKpn6WHo0wPxEAKuYtYnd
T0YtLFVh9BOPoJwgDicDX6Mw2QVrAL2ReFU7Dyhg2IzYuSviH0LWaNP4zarg8syUWyYrOiv9TgCw
HGBFMKyF0yC5NzvJsmLMddZUTMbeQ7LTTjyuQFzElQTVD3KAuoCcBTbU17NfIy84gnY7J+Iry47j
E7IrPt/4VXnkPeMzYQzgjxf246igE9A0X8X+ZQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="cVI02/55zpM20oQkc42DB+Fqc+OnsAdVuGA7hwE5nNA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19936)
`protect data_block
pnZl0HgfMR9nnBtd7GVkFwnUcwP3S6Zp74W8DA8OTlHScs/Gb5c5GhTTjerkNau8LkDjXyxXWCTd
vzdRtiSuhYYBFBCIBjU07pLMKPMfPQZywROLvU4FD8A0PBnzY3VntpW+W3xFNMtyUDVrx4VMn8YP
T0GMB5yR8FnOfS6kMa4siNR+HfeDySnAASg172JcoCkpbmf9f7k3juN2Is2Gbnx6Dh/WpMWTXBpD
Cm/T8ILt4ss3mLZPEdiUo7O1LCOS4mvTg7zCE2mVhbOMpGnGqBWf/8zw0l9SE60e7ST4qxVjcUxb
MIIJQ6HJHvzQmWSkFCI1tQoWVWx0uVGerw9bXEO+mdBsmEL91aEM5M5UxQ9toOSJAU48lnumTw+H
X15z6Gwcz+yPlBn+ac4CngHgaa+HgFxKPlqJ3bY5qE/bOJCvvjgFaGUBSgCsqru7ZhG9itP6NdUL
ybte/dxl+ZFuDW82kAST4t4qUaW874SFmZ3qnBAgHZBhNkac9oYR3b5GnlpzoXziu4tiJq+nipb7
GEQB2PGV6g+FbqGe1fykslLMLS8yIR79Jq7lPUsm5/7n28R6y1XMsWtGN/CvvIyYkdCJLgrhnL7B
d0KOyF6bEpszsXGCA1f7VqaXrOijuF0ST83M34Mifw58mTB9AGOh9h4ICZu/8TffZGRjy3c2F7r5
AWQ/CStg8IFb1TEMu6bn1OdMfqSnUgj6cvIrEDzvva+gOHLkrlVxa5nNrjHcnqSNlP6jujdQOVMp
ZMHyYR5CcR78Qa9Bj5Czv8AbSpk1YWMS7ORrudhyGNzEP5xWFysiCFmFU3lo95BCcDGyi4Cw2pdW
HHGx/BX4zpUFJsqOGpWlDvhGPY40owpL7YnNtgoSUZrL+GVg5h8E1Jx0BoinitqtwRI9Tp5rAWDX
l6+GVA6Fjp8vY15Nz6V6jU+3GLK+dYsCuV9AUS1V+RCBfHN5OW7mTK1LMknHLLjEPTLmUIoJTGuQ
BPX6Hun262VbP9584yHrZqYLjqqHpeB99g3fG/qP+RSDh2FIGFZgPCUR4j3G29gqJ7eVBZ1Vriqb
bz6tdGhu3yvMvRW51EZQi62h654H83VynhTSfB7/m9qhg+g/3iFGWZLq6RE8Kykc+UJKa05MMc/o
x55cwzQmF4zLk4e2KAjArUqDqpP9KvSh94I+7lhGBPVpo3jCDYJYAgi1VpylvMcPUqZq7cGO1DpD
MvMnkX+HnaCuAh9fGY5IL9OCPy6nBBNgpnbNeuiuOC97dv5pvJVq26CzMWcxSYhm8b6/wDI6kn50
XHJY9DzuJj9S2J/VfRIe2lKV/9LkurZHb93AxPDguuS6FcmYc5OqxjavoZfL4ndlrjeFYBnxHxUn
nEOgncG5bS5L08zK6ZN2/YcoxscuvNeps4UvNSjNiE5LQKMhVOdFd8Gj07tBY2em8HO/taZLJBH8
kYXBUgauDzBgE6N500F81O6qQ7jERVHdcJZKktDuVM4rMGfrTtoUyccUSQr9W+gFhFcSKsdEMQpe
rH8F3sta/41WbVUJThwJElsdfZqCkNwGf9OQty2yc85ovnNXyj6pjxng84m3eeZbDMwx/sbif3J4
G49Ji/F6ZsWgb54wCVBTQctpooI/rM0R7vH9HEENYpBoePQshYrnSZAl9idEvOJvZw/R3xwHwC+z
lSh0dCazlBZnR0A0v5kv58UBtOKZh/O48aQAH0ZDxWWM2TgPpN03R0Til23B6l9qlFqs6wU+dzvL
V7/keQlSjmbirWRbJrfwLV61EHZh58AqtSW+WpaeU5NOC5RY722eKHtDTIFljFrUq+SKEtmljG50
yaq5CxWk7amUS7NdIALjgLjdwrlN+iocIULHYFcJVVPl9f7i1qjPMgZngUmfAIt1YZevflFMRgry
tKQmVk/ZcJ39gjnDYuFoLKnQCEBkOv+RtQuBoypZMcXisMvmYqYs3hgJql3HFxzqahZI98OgR3NQ
jwvUuF8trkcsqo8BAH/pkmrS4l3ykag6RW8NicgOBrQLQ5+a2VycX0s/9i2EosbdbMbHwsBaAwi4
B1MLnFFe2TtkU9jMdjE01Iy+aR2ZMMiFJDRhZOqLA9EWUTREKwgOeWyzNB6Vtzx7Whti2tRenHV4
VSSUvSGXm8+Ht392ZRooZUugbvMf2Kgc42D5EkqocIWvftskaSUuEvJoihHj8du630bJnunCknFG
Mdpcp0OxdsguPV853TfRpIp8PI5fIDa+mF9NM6jwa9iXaKg8sf3aDqdRAckABPpXbJoEJ5YTWA6V
gi80ItnzTx9+E9tgtY9fRLaEKFEpInu7CzK+9+asI8g0CQJpPLFW+XS3X3Apc7QvdUrNqsXCunwm
TLxpWbi2zojztLtJ17Z7nC4/2eV8opIG0AyUUZI772h1dn1oGpVGk2xBlG3bn5pMVtaEcalDrADD
DyXz/eJHm/LePnkwqktxLkflMvv4ieDu9kPtMHkh+rbIPfvHkBYd+/ZzGZxl6umbksRaERK4/hkW
Y9/m2B/0AnxDG62w5jK9s2uIoVFsfbjzh8yL05uKE1mm0Ru8JdOMzTGRyqadCDluDSgOc9fJ9LEg
xlZZG5QsswC+MpYc79XyEpAt4i5x/W+3S6GbwG9ergrnUnfQ4+v09Co/5E+yPvrKCA8ZPwxo9Dz9
gN4NXSe7O2Ue7UsE98HwG0qP82MhbtgFElQrhXCLrQgx0taG4IOQ3zrJRp00kDoDi3LJ0Af4pE+K
s5NpMCGjAPdkZUKSrNZ7svscgwVMRWDautbKQ8QO9krh8mmuT75mchz9CFjm9Edho2fJ9ADAoF/x
qUhm4vKXBNMUq2Y8u6aEi/XfUoa97nk7H8CgIvflBNPT1X8RIwobccsEBVq1mIupy8o5FuJeI9wb
Wa14UzLoFjKfbAnuiok/xMMNZi4qJu/XSpbiNb4HVXGTTucAgFgC0JLLAJVqe8R4jdJXg+qg0NUi
Cm7/Zod3FvmViYg6bn3XkhkAx2sfRsaFoB1gX3eIk127ITGFySCG3qHfFr/itH2CtDpnx16zVszS
vChwkOEVRMfEUSqxG9YEt8g43Rx31jCUkBqBp3LKIAXKiGnEigfouzHDug8ccGOrYn4PjASFldGC
Rq1b7BDVQFn6GqbsEpb8KXNiHhtoKiwlZYNK9wcYaiwO2sTXIzDjTYGqCL3Q0ct7sxmoDETYdcZK
xFxgrBlWtcaCmKwiX/VyGs4geBVaLLClqKqf7G/7UMKo30Vc681m+sv0ICXW30r6JT1FD7Ux//uO
W3cud2puydBiHCtAUsK/YnAPu5bvxCn45t6l/EiiAGG4LHAMhOKcZJz2cun6zIqy5my0r6NOuYBZ
N+jlfWxUYRDB+1XT3kGQ+pgCh2qfdyH0EF7r8gxPIvtWrn8cV591HoRrK6jqT06zzRxhsXm2Ofvg
5EOK4z6lu19sSoPqCTvK6PjB4o19+xAueR/9e2Q0+FjbAbBW+sSCsxdTLuV+Fa+oki3qXrib1Qa7
L7C3lS3kdb8o8S4b9Opn920uBFiDvGcS/VHXyx8zHeGlWyoaissooD4Zl29c+jhDneeGqZW2roxz
saKwVxcrjEo+yD2amozljYq9dD1HKK0z2nCcahG8otglZQ46By7Y9Jt8ZaE8NiHcSJRck/xUsG2s
v0018MJzyzRCCas7IJXAOhm83m67NFByjuIaJ+AYjxhPC4GRUCE1LmGkHmielfTWD9zFAhGKgIYg
EBcMTQ0exZkLWmT8G4HCTDQH8jZRc48z16hCrqCH0sBPh9s0ULSmWQ9agN9ITV00b87mQxZA5esH
jZDi2TyMwXVMo1SLoQGv8LI1X0sraVVTUK87OTQew/iHRF1lwHkEvWIUTKjRDJqCwNObso6xo2Mo
VaIRw71IvAIctigk/zyz1bEnNBDT8OJ3oiFje8aQJNHp/Dm/K6oUmQaQHEyyn78Lob3BcPja73ac
FNbITd/ACNxbK+BnXM4L80IaN7AZqvMzBrdC+uz9py/6bjDoed+EDkTa+AS1EL3tbPMeTEe212Bq
23SUdTqlEn8WseqqOUbkME0hhDmvIEFhXrOTvEaKmEJMugNRjP0BEPSLq9dtjAO2z5voP8Ycj5GV
FJNqIy9dDf3BhpPrloUa88QGlFTWfZzudvLj2wWAS8TkdxnQ9jJxMFIKBfH5IQHXDE/dXjFetFMg
1zm4oSKtWM4JgZhvtJBHx4kvePfWcPQHcGuc3ShsNaCmpIhZy65UVXDcWT91LRviMZwzUa6ep2Jf
BgRCbhYkZE4nwCojIv8S33+oU7MgrV7+g0FTmYOmVLg6TC1Cvv6M8rn0I+iqFRTVf5y55/nm1Bo4
W1jiU2Qc2aA2aoGUfBb4zhh+dPR4NV0NyGJoO7b3mbavToubQ3g85iB5BvWyBcd0PMg0caC6FeIY
d16t3sSHihG9qsy/wlD9s4I1P3fgbE0k+dJD/ZgH2qsQdkaRwatMNHzEkb1Sv1ZhKMeLz8Pw0z1k
LCVh2W1kp+mF5mDI61HyznpM4GtEL9aY01roQ6VmoRwcdk5pUmod/jYpoR9EytoUENyln4bU/HGK
VtUk2R/6vUctmBZiKGXh6D1c5/zF55gpc0VI6+6iJaIZdp9OvavexWY8486RYCNtdeZYL8t4sD4W
e+zCqLWmpyjrffFQ7A0DvlDWRWlTbhSEW1Xlhih1loPnG8a9U1dIvjXp/ysp4OS2riYCuS0gFDel
uAIZDdeXgelRN7IU2gbGfThIIv+H9NXFh14lCoXdizpnjXff3EqyK+LX9I8QfhrgPeW1LDwGbjPr
bfTiDZlqxcQ/JZ41lhAqwWC7e7knmX1q57u8dl1SM3RslqUDbnzRSEKdH7DOtAU8GX/ZTv6/Hq8W
z0H7gVm3tXgRFg14B5kUt8n/HpDec8AU7RPNexQmYG/4c/3l0P7VbBlmunDMBADBOx02yUTVpp8m
dt+T1yE9q8STp4dzflD3MHAPRpn48vbCQ9JRJOs8kG0fGuItzmuBPSyL4QV3aCTwvbQEEp/JfNy8
yBqR/rfp78NyCa6SiNZZtBPzG9r61FhiQDGRQhWQSfuBG460DxjXTjJsbYL82SFalOlWulIXWqPA
N/C/l1t8/bS0IZi+zayeBT5yUvj46QFXts6wyLnghVEK4mTqZQUCvmSLvw9xTdLd/aUcWV98aUZJ
YVun+dc5aM1x5KPA1Fw+GlTb5/eNu5QvfF+6ZZIbdVn5b/uq8iY+jAz0eYjz/3Ezd7tZ2ZQSaFdJ
Ip+nE2SmRgSJP7veP28AJl5S2cXlvKoRvOkoDuzIxpZvKfv2CFCM7Ql2XLq5E4AT2H7P0ZWzV3vC
H+gadDkypQCczSS3f99CRIAAIlDwx+ffoafcwKRAxhZkrIXvIsLtSGuCWwuxUIO9Q6NUH6eJ0QHG
fOHo4ZSXIvX3g0HeqtIQaSn55HDvTyfUxr3w7fzK5k07s3TnG6NKtuViMkAEPS0oHtISt7PonUfB
P8lBTQIzlwtdULTMMrq8YJeAES3NAU1nYahzOdvDOvy4HMZs5nAn1N0sPvCbqKzTIUz6z89CzjY9
T84Lp9G7hkoLwUvF9z9jykgc53jWWdrae+PwF+8H0fFfeO6jdCUGSk92pdnqxUu1NpseLdztiUvh
Nk/lwDZehHDVIYMFSAOo12km84wA2TrDirEVOaXOXkT8fu80hLGa7BqSZbiBfkrPFYyVvWnhdhp7
gwRuy9ax0gvKzQA+AMChW/pRqXK7oLOz0R/30m5lQbIan8r3UTp97VXggm57kxgJyNPN8MJZAY3p
jFTGE5gLyEVA6Yrso1sbMq5trUwerwc/3viEYMUZZaj7ideQNiBKNjX0KaMSEq2FbRiDqjuUtAKq
kbWJQ9ANPFqiS3mK5u0dtKNw7A1+gZVxT2727UJIlN7FWbuVJXi0YdvyTmj4UQeRNp+KQb3WPhrE
LYCowvm//R/FuUCZf5YtZyT0DxfdHnLV/igLPI5kU7BcHBSObRQdRmKWYO7L4AE8mPbfdcnlDTZW
h7QuIOwMaimYfgRDeTJqTekgcP55rlPz9zres9IJaE+NEdLPkVigoyObErwwd8mxMRBMrq3I1HNq
vkxEa7sKgewwGdvFuhYdtNCLjh/arBfGYKylXgwBzn/n9NdajhFuAUU9mErxv6ujeBj3/Y/pUBIP
xRqXD79yqRTTUifvMo9KO2vT7DPubF0OMqXoFrM6Dzkz5UBJDayIoEpS3SntolqnD8oSShQsm5pw
XgBPUXUHOV1Z7FoAq/Wjy4iWVnJCf7zE3ouYQ8nI0R5/1BZy9XWWIaM1cZGUUC129RHih0CFGT77
3Ao7sTSUFz8+pwPERIsJlnPECMHTKqowULsHVzGIU8ttevoEux36nt+xq1ZM1qNNLpy40cJXeuii
fKmAbkt1uSXTK6Y/xEh46Tstn4kHvo1oygbxO+b9wm5MpqdWeB+naG5xv922DR3Fa+AsuY9pzxdr
0lAYlyUYKDisHmznVj/Bbn+2OT5tcXSgaOY6DFtC3CxwsJ6NEga0GPadc2oxeavg2V3gu38op7s3
943IQeMIKvyX7Ki/SUMbVy709I//V1imi0EKh7kckI4QYaznnBBBF13hEUVdXKnIri/O+Q3BEZOl
D2lioCX2/DAUCN/5r0tYW0ea6VGATunX9FcvKLwvlB2EL3MWJpBLftJSw0AOy3yn5mbE2CtpnZCF
dDkvBV3lcraxGnHpfasnKZyzIN3ZTaRx6jHwfIsBmIDR5m9NXwgczBWiK/l5gD5cW3INxUsB1KrP
8RLqRzhVPw5AKmkw9i8qW34yQL1XKbjzltHeEVP16nGbLdTgeYa1DmT/+Y4tBkEn9i4lv98iyVyX
bZVDa6eo2+SJguLyvHCIPYKMpAvCMLmOboFUPQINa1UMIFsuXHuoZsh7FI8XEsz0hIEss8Mu7RqG
RkwJoYtAaQTwoSXYX0lcyS+rze/Qj71hf8vwFYdIzeIO6EW9pinrdQ9Hj/qAyv4TsKooBVbMkZoC
mRtACRlS20c0v3DrkWjVCZVu5MT0muIDz+bXHzFY1vVbOHPfAtxH4rbYA9yCmyTeoADyxKauhhRM
3qDNpEH4uT0PIG7D+vls40F9HywnHu4zJNRSHObIjBNwGeYksQf2kJyNkNolC8V8jjh9E38tGs3z
ZBkPyCtGBw9q6vBkRsWYUKd+AE6YCTLHKKXaLyl/TkxY+D0JYDB+kpfcq+AjM9FkJPFHfC5H0Vwe
iMuG+AE/8O6zihpr7RI3ludwYPJLy2eRbMo8hM30TSZeBuiop+1ph+GT/J4EO8DBt+6SWGw4r7cF
K1navhYyFH065GTDshcoFd6Pt376iCbCsf8fLeLTG3nSjdrfbA40dKz+IGUTvHLWYSqzxA0rGtVB
zLkrw0Hdf18SGChUuDaNpFeWdN0giI9l+O9ZHf1GYvFxBUClJJ2wlvSGs8Ynnp/ronSaRRMjiOjW
FhfKtB7vEL0e+XAYj+hV0+3VHs0/Q8YhiJ5kNfDeBKnDno+rPiVFS2GkhiAW+kwDPd/ei1a1d7V3
C/thTWG/eAdvYsx2GXfKOapLdYbJUQMYeQv3atD9320ZWDEHGBY6N0/0qu+qx4Lw03OX2JzqNY0e
kvoDeQOtauBS2sECY2ybeQz2LN2SUkuL2igW+hoeaMxICxTXbf/ehOXEr9TA855vOuvsDXof5jOH
7d46L1X+B5UBFI3EjXbrAirAzlQJNqb893ZxGIr++khHWSrWsTKNzHn+Q0Gj8QZ8zs1ZtU2C/VEP
qYyhAeBiUYouvgRNwIguGyBF1kssETHuxXuVgv3zcEVYrjf4MeP8/JpJiwzEdSURtRsLx0zk/zV4
ZZ8CEdzP5g4giMeR3fPu5TCwsP5oxorMc2yPNlQ8zmrs5w18N/u+4wRnByPXO/Yi4f+6+Kwl1qC0
U7YnahDXmGkbG9Ds/V798yrpt0qLfngKujXN4u61+Y1Er/99BaP0egLIvci+mX1wyGOFTomrgRk8
SXQZuWtqxqZppNXJ94Yzdhm+qE/ODGrc1Magx6FpmrWhBl7g/0l85brmbKQyXjV667YnOXHl+UEh
cWQJQoW3EMnuG1VWKvNtd+9Npqzf1JtPB484EkK0NqK0UCKAP/vC6ht0ic9P95PwZ4f/Bx9vLIQx
/1Mbxl5g9gwyeBOuQTyHmLXddgnq4M6LZYu8/9gK2hQybO8FsIRCT8zsW9ICU1l7tgTgj0wxdVkc
Gsnmh+6U7iL4DshJT2VD81Ym9sYq8sG9OV2G6GykmDE5IhKHkZFry2yYZ296BHj1RvC8j+6l7Eoa
/7K/4CBlyBw7WHOhh91lof156oWQIiiPSVd2+KN1ZUV4aIYKAV4RVE7xzgnIsQJJfItxyXwC3dM9
5Q8TN/VgmKBSuSz9x4b1+i7WOxDXEH9XMoKM5ELnJ+d2XJf52EdywUthDzyNoXI7ppO3hslrlWjA
tYPHVbFO9b0c77qPqrKI+bYc6wPEMkZN1obC7v3IU3q1VDjb3g7F87sla1ssmsI7/pEdFJJVzctR
GVzU+YuMEsZAq1WY+xPXk9RM799KbHoCYxV+oiGYzEMLvCx82cn7ioRsTYcCELiv0rbztoDjO9hs
ba5Lk0Kpx5/85sLY/IlI1/X5TNwIf3E3Y4/Arpt4ceMzU1Hndo+plSs/Hhxv/rAVMQCTheydpd0r
36+CpKxK2Gs/gJIbmfWiy4/Ay0J/fwfK+Rtmu2P4PPCQo5xp5TdI38dUwn5blORh+OJHInDr8t+J
7MsbnnPQ+Tn53WfzlBCTVXqVq3RQx8YjfDyHxNIP6j4gYOrZyF1mER7gloioFn2WzUWPjv1GTi/2
/dHymNG+S6FnxarPzEfjWc5q28s7DENBy60iVIIVX7oUj+4p2+wd1Vx9Et3aNWqIbumvCwdS3N5r
GYBjziBdOElKOGigMHlMF7Bj5W2fpr8VEmdlaUuxaZ7egZZbNb42paR98FqfG19i/whxkXBc/i6C
PDLr/1ZpVC2w8gMB7vsUU2cXJQlSf4a6U2ivJR4i0YSnwHXAFsrNTeRet3CPW7prA7UFy6bbU3gK
5fxAB9n8d/qTPPwmVFljI9KqbBp21l5g3CcF6voj64qxQCSUpP2Gqam7BQceKt5vOBY04QDnkOzm
7OcbO+A4GXMgg69Fn8cV6wdReHzlbb6LdeIiqm80yLLanpFHq+iKXZSc4KjMh4JkHYkNkMUcNACl
YmwyAQpZMTzllMOWI+uFi/hcE/hYKZB/lkdrzqrFF1TJjD3P/+e10YlqNWlGihGLPiHry505YMPv
RiF0XO1dAhMmK2dSXwC8Ot44XL3zu+7x+q+3ehjUu0HR5pTLXH51yDbqDbm+ui26PjNbBQxO7b1o
rjoertzB8br++thWHDdJk5W1MouwONpxTvgW3vtLQMth2MA+DVseQ68HLJsu4p17kT5mk/Hn3nB3
Zj2VfU+BMspcFYTEZPW8J5XAXFoGQ4PNf+GwLQob3b65ZYh3wnCEI4PYP0/AXm/1UkZsrrNHJuZt
16V0JZAeXdYSYIHW6tI8NEodZw3abMXISH6fKohbMM4SSHlExpdiEbpySVIYRO0NfGKiMpKo1ZfE
/5aWyL8Qpb0D7ljHDW5eYHY8ASCD021c60apLogl4hk+H1jQbFatMU0qj3HxWElhu5xFFGaPVTGW
PRvBrk76rFPi4oGMI9qf/GhLP7+KkbaYpqk4RJx+Vf7t7UMbJJW433YrNH8v4R5B2oIM1ICU0Uo3
OsQaxMmLgn4qbpxw9LNR6IDd1bYutk1PUmED6O0GvBdaauyneZN+eqhHDZWcW7c6pVaEh+MuCIt6
BI7UbAi+Vd8xY/VIQCtvV2xBTRZh/p1PHsJeRVM424l/fejBHr7dvvFX4KZdsLQ37tOarntIGN8S
QET2HirDhqkIsvdMKLv6yviKm1XHZK4LG/liSCQJuURorMbjam+XdIpMcdo+nTr0Fzwy+08GmphO
kB0nlfVPNo18DdxAKS4zXJ67UgxRHmgmjyQQD5oB4+kJ9SwL/zXTktlyn25dsCU/st3pK/Vxk2n0
7nHz+tUp0gxxXHVLU8bV4AATPXRm0L8mUQPukcqW/tXGAoftzlGIjtK5xKc1vLcDiEpOm6spaCKd
h0FEUx7TN1Kbkq5/0F7uUuXjvGpzVTG4lHgErAFC3LPoau+DHndq3dalfW3pA6Hq1ISqYlKfxOKo
rbij4SFKrscf2lrDb3j687SZO87rhUeuqH0w19GTP0EsNjuJkxjOWDdPu/Zhii85rUVDDq8Im3eE
XETvHibjilByH22ps6+y6uv8jgXvANTbc6OROkcJCuxCIEPuCfCkEBTZr6X/G3TxmI7prfJvgT6T
48Wdpgf2ZoezIqp00t0QngOm9elGZZGrrTgQjbjqDmnJ2lLBxwJdJazDOgV2vrzjAsfeS28Eu5Dn
mhjsgly9fCN+xeXTAa0rcdLdMKa7MIdgGRvt2aZN+v9xF+fEJgIt/ELj6c888uuh63xCOHoyz0Hb
gU+EVRzXOjLDnmavg6F5bB569EpAgJqHuPDBtwqhknCW8fp+pJhCaEblYXocIyUIK1Wbxp6ZfUS/
KjvoG6HEupZKZBM2exJC9g+8I6fVgexIe+Tk4SL9HHg+pXLQukrjmvrFl8EREko+v+uEbgwT2jgE
MepPGxYvD/kxYfRqjo6zTABeEHZnyn6OoYcDCPExZUjP33D5eoMYnIMVhUD2VsZQFAt9XqfZiO6y
a2wKbvTFLKAnKNT/4lrKWwVZUsUkZoFWprAaCutC+exojehG5IA3QEEcnJANXhxtbRBo3r3OALjh
Q4dPm30kjUCMdBQ0EpusNsFNpAI8gVR4KuosgPSGXWsu5mDDmG61WM/9aZ1hBMNbkt84omqOXQGO
uL3asgmR3qElGJtNr4+KFdqHQpYm1d5CTM2g+QI3YUAj5NqTew0pr+yvLXpc4HfbdZzQPCHuaeS6
dIlVmibzUdAW2peVOkuqHhY9tcLRbh4p6HwaMMbjhUYObvloAb/mzmHHtrUZbwPx8YVWt4LNtPRn
qcLIVxjJZx2h9Lj/NVdDWlVWLrCmPRVFH0/UTD57Mg3w22ovmbtihWpqWHAge67zomF5eor0BBnT
kw/avw0opgcqsgckwd5Iq7m2FmNvNT7rdK4vAMKt8KyKE4o9tOqkvKs6oDN4nRNi4gizEyLgDQyw
9aL2ZvOjUtUZTXDbSE5rnG5aBLJEbj0YGyup2jpj0F51Rm0CTcOHy5vuHxzBiiCDiGYMM4Bwt6mX
cquW7gUrjem+D8Q6z01jsBR86d5cTSPTHuM79zEskpuaFtFL4/zFX1OLlPs5ouiE/JEzZ5ZfmHWM
2XEt0KHYIqpjeeM65VlXNG141DkdhT2cbFk594L8dweB1D3jkn/f5m44GO7+i0YX1MSmd+79uHk5
vCPUt/uUnjRGoNu57WF0K7TXIlL5IORgSNJJBqfjfnRoEcT4bWSnUKJdBVNY1+ChYAWHm232QCO9
tTksr4OtBH0tEZsIJzJtomH2jpjFw19PU++0qN/WYEzrnvIHIpAI6N01IQg1t/e7lHXqk+VecQDf
fNX3pji+v6aojSRo8yqsktAqD6ZutmIf7pgiTu7YIM1aoP3f04t7ipRk/tRxiGZBJigoY8zmvwN7
iELJp+IxJOB9XcHKkSK0aA8NT4SjGhnG8VsH4t7WcghvUEJEfTtl7pc807xQ7ONz51j2v26Iqxsa
aY+ClF6F0thY2htNvNe1PIBS56oplWDboIEB2hQKij8TrubpRaxuuMI6w2KKGqY/JU2/kg+p/HdW
J1CcL7+mzhSSaq8DDbsN3UYnhyNx1EGxC9apv7u4xzKfcw5mUWP3KVgxTPY8sxUWMG3RrctXbgZX
EN9KppOaFl7TXWJ0NIxJrOja7gTt557qT7yyExp+Z+d9sPqrjpBkglZag5yFnNvqZjoSq68iLrDD
4J4TMGk5nl9P/OXjA+6AsNjPAqwVzBRn4a3uHFKFBxnsdewrwim/am8OU3C1Hr3jmJGWt0ejuBfl
Humdbqw6tiZtOaA/9szyD9kZvdKIXzWSdjujOZ1HQGUgfUiilE9b2ekHAvUsDGfW0P1gjz6CeUTt
47QhmY+Uymyz3DbB0HJOUwhdsCEpkUYNn0zbzyOfIlbFcUImpEHV3VnAYFTFeruSXv5VYH8mx5pC
kwzKAZutHHiV/53HJREQfC/cmORA8sW3cAkaGldswX0fv0JPlFQlML1m10cYdnb6NDIut7MTD20b
6pj6w0oxSlTCzr3ZodB+MqecnEKFxWToUXvBfljOoZPGmJsdjXbOYsoKVROgkvpPCPKyw/boxWtx
SJJHFL6YYpmoUJQi9rztE+6wLSiGAJWUsJ5bvM1I9vfg80BrH5YGGUNDKmmKo3VSzotKcmtX9RC9
Q6TbTQHh27UmNVF+63UWGWSce2LN/BExelEOh5bK5T1tEfJKVB+nkHKWcji7ZGcK/YNZ4aRAtsVh
NKFm45x9CIMa063wAK7hv+AhLoSBMObg2htUzPdUhe5aFI79eBYMxeUExdrwGPq3dYb6NWtCT7mw
GFa+r4O4fl//9yvN9wJRcEDBc9XxBxHb74VwGGSezrVmJ+MVeNx2auCdqzSexKywUvELoWTtqc4S
WdCv5En59le2v7FZ/6x1LRrZ7fY/z5kUCf/QCemqbst1UryOCIQ1Hbz2A/5hwvUTT0Y1hAQNJCjd
4S95ZYnbaOf5CZ1mbGP6lQf7tdlCm0Py7SoKc4pdVCgjazqyM7gFzHhoT4pfOVZmxtB5TaVQ/wDs
L23issjMPpb59FD3zBCTxixDCJZMiYOp8K4emzMc7B/FBw25+gGv8Niazi9vPqwXDFPvd5P3EwmV
uJOxwq5LclTOWU3YlZbSS2YXtUxrJwo7Hq4x+MXMzxZgmJdTKdD2CAe+7MSIMen++QCvZ7rlxbou
DW4gF+IZs07C9iJo9E1Tpv7AzQvn+JKpvJGAOQ9K73W2l6FabY1UW8o/vXMqc3DxT4B4haijhMOw
h+zRgOdYthFGV5LzJCO9nnKwIMg9KUwF+KgoNKUWRZnNNObQpuBz78gktddjbhnFL4q1nKxRd33+
z5Cevarcd+HmQotyGB98rCZChEyJBoJsFkrSOnDo9ulU0s4s1Gd4Ds4NkFGI5zmx7Dl+SGgegCKF
CUaWB/sc10XCgTe5GFXKJlGuns7AK5J9YPdOGgv+ambfVIyJZokaWd8a7+WBeN+VDXT14fBfKMGL
dfqSwRbS6rjOSKVhLFb5eGGOfW+je29zUUY1gfhdpAUbuS14sBLwsdMAIud7J2C2mi+B7oAw2sGE
/UER78xzpmFNQRvvewd+N/P3Q5ccuKFl71jBGVmPrdYglCWF5YcQA+Hv6EKYtbsMHY9KoUDdB9QP
6JZXgc4kWRfAQtrcRHlvv1Caxwvln5amuishGqj3VZA8wvVb2UKcXjwzEEFNiM8C44QA7z0r8N2q
QlSDHhRXVo8cKh0sD5ehZ7SASCcfeOqfxjrD0bAkO7QkqO6SMlbTdH7OgBumKK5mMQQJ61xMJn3h
CRevLxHgzVFVyLKhEoiAnzz91dHAAPf7IOwtZ1+cTfudJbp0oE2GjBVx6SI3MsZMkkcccfKcExEA
t33efC3EZGkG3BiW721aSJWXW4CJCTgclYL388tNmTDCK0x7E3a6pdmCnj24K67gfU/IxgjTB9Nh
bMaZWBYWO59lH+hd9/XKTaWRHV4dx5lSL6Ao9j0sSsZ3IfNUIFqsF3rOWUQy7MqMZMEh2pO8yUQv
veh4kmvFdJ8eEHWywujaghco0LUFa228gp8Phvde7HctGlpW07TVr/GYxvpXzBD1y9L60AhuAOKk
e9Z/EPUaac4N1IJHXxcLNiTJtLPKa3WIInqGRSzpRxfvT4WoF08c48NKl53FzPq/vP+Pyhar9kC8
KmBrJQK29ihuk1n4ciNhzzCJIiebAD1UtfWe7at7dD4Jtd90AWl/MNyZySUI2c7KxxdZV7wwyErB
FsOmSOic9lgIbpfqSgpCnjUfZJghYeQPWR1ayDMDaxxvyXINg/DBxlLINpj7B9SYN+8b8rOoMkxn
bIqG3/jwQR6cgbqAxT5dgGQfZMj9cmzUyxKbo56FKCIU/VcBWa10b09nP5ZkQO9AHY9MWQT4SG26
wxnti/Ql3+WHU1O5iREDEgZxT2WOb3HiKGraQkxsT16508xaTsDuedo68bnOdt7Dh5BetJUBY62s
H79D4CUr+N5875Y3pOlE0/v8OjcbIWjDgsyyn2wGV5afrti2WlTp1AgiOwvFm4xcD9pi5vdXhVii
1vaPYdEWc+WLpaAzz4rEFYbZ+f8/L4L1R0eRdR5oBcl7ZIQB/neoazOlduFW2Ne8ASoSB+d/8dt0
Gm8rbT85dswBQVBNMkDVDjW9UjSb6i2IXfpJrUXNWH8OwQVrLOGKR+YFSyD/rwT2bfkX9I7xJL3c
OEC9T/OFKyeTfpXPYd2lp7Z95DDMHS2VvUnJVGnoGzyoI2poLozkflMTQvpBcooXVZ2GtZqWe42t
gRUT604H2u6kn0T1wD+Ix+We+E0UgbULkgrMW1jcobncJoomNDTPrailb1fb1gXSRdmrp0UNLKFq
MuzQ/7JxpJIRDDLODVCW5tM4gieJ9d3GMro0qJE/aWESi1aX5Zv6CMISVxfivVk2dN/t9zsP/cyF
aeVFYZaziDsz34cYFBIMlgIUYnE3AZKfR7a66ZUGQWdRgx7byP4vVl/Z956JVD9KtxgH51Y7gMko
KeIvZktk9OLUPElw2jb6SraAXGIYhozSS6k+PmSc5CUXw6MVQrp1JkCYsJ+0VKf1TXcRouChO7QT
NlT1abrqv3c8eW78KE6mIoX2v/UA9n7clONgwe+JB95ll2347stT5N4VcCzNoci2I6KNdkn52bZN
J4KAqkvBqxOfcGhjZ4I7Iu+F/9xZAgrejA0DZXVuHMp6Vkb3GRVibOeIxuUp4A+M0T1owvAQ9emh
CuiOxu60uDPmi/ssJmiS/IIFs3qt+id3/Okc08MCPgW6SaJfFP4LO5thDj34ulOCgOdOYC/PTcOX
aGsfAZo2yaQGKjVmpydT7qf7Lp5wPQw1+6zekV1YgklknfV5Fuh6lMjUsyOSpSWAt14bFYCikFQA
/JqTC+ni7F/3qIuY41H++QF3xFMKengbHPfi4XMksL/dW5+N/bjLMnBSNbpKUA6hE98vA/jv3/rl
TdXTMePzzyx6U9PUHx94MJVAyfMORURnfTad5nNV441psC4xDgkwIR0Y+2mCCQiBPALkk3I1GA/3
vPwbwkUbJRso3+h9hdZHV/n+qbQJQzBnXCIuCraUeOSxu81u+xr9dzTX3b2UKo92HpblL99WmkdR
U6c1Ah0Orlv8liM23C6e0fQoMa3cqKju1fEdRXyiANXvpQuK4Bzabqq6oMCtX8doFzaOxOrOkGQj
IZiTXHge/0HXKMcgh+VEIsRxt1KX3VtygpI9wcY1/jHb2p3raQ5Nk7ORywItG4U7G3mTGnIqUCQ3
ZhJZHkAJ2fck5HkxvpWpil9jJRJcAK1dOC2Y9dwrfupPkyJGgzA8p4glqiJifF1QMd77Ip8yIq8V
5X1fR58KLtRs2llqbaV0dI5pBEtm50WhjzbsM50CPYH2BxvALavBpYfj8xpOmAw+cl5BQoj227Ql
mloyh5ogBvwQvIN/8cLMBMPq7GcBN/Oy1QqCBHE1lg67UMiD8gBahQizFhsDSNmYksHFA6gLpnMp
PLw02ZtruOgEbBb91bEoQJLtFi7WSk+tWhsiOOzFTxgx65QB8m0naOB7JvZey2umcJzO+SeKS7Zj
NJ9shXQHcQ7CHln4AmZR+QlMyhlUkpHBS4Z5j91U2Jjc7A/PqLonW76dJP01gVrOhxcTbYL0WvoJ
rOfUpQs4nI2ukP7z298T1N+5TABcUB92tP9DmIXG2h3HOR2U0zwKMReBFvTOIvSAOJi/Nx43zoWM
lOWp+b91z/jD28uzMICZOFR6hSGa29iciEcoB/L8lJBKnx2yo5rQPnFVCThckhro/3LCOAcXFao2
r32pILz8FVPNOLLj/4YFoI0q4u8yHzwqEFTizU3fn6CrgADR5pjjeT9DrMkAySrsFi7xSiTRuUbD
+2tylqkT97KWa2AAs9Epgwvw2ihzBUBpNbkYZQkTaXSM3CjwuXeJH0ihSdLzZsQvJtKVWJIeU+KG
vL88AhsV3UbrGGhp2gIMibTBPLqy591Aio8lurmyOKVCeyuPlLXHCRKHOM4DwdWU+LoWbk//JvtC
dE7Iik8RHqt/PATlEG+P5KyxMpFFwl1FuPrmNLb5uVzGbcV1lI7YyhXKMtMZWwruGSazaYcVKf75
laV9d42bt/Uz687fSfRP7QRLgUXtxeFYU8UdI5UQeS2G8qn8yM2kL5iBgOU0nQQZ4VUp+m8oO5Hm
jxaRbgld9bxIZZ7JgaxCt66Sh9xKZa+fJUWE6MkreMeZPBqBecIQt5+RXyD0XIh5tRjv9boZOYbY
U7vMjUkGb9cy3FpLyJevUOLi1S+ovvQMrD6uMseWTqjNqMxz08I6q+jsgFxqqJWmlgY5qVxeUtDt
6KJpdiSzBtJtBbo6NeTi2b3fCrPNu71DsczefurNnG5J93V8qnItA8ty9Z4YYL82f/2pCwjo+pPa
a51AyKOEXiRLoWaov+NvF8ZQILcDhhDqos5RMNckBLB6qlbjD5xFSiFcQJWEodFyyTXSvmc7jTnD
bvxUKr90OIhI/2MSTh5Nqzj7htlMwDhBwMA0JX5D1Cwy0DDkblIBbPVQcZFLVvGrtkizDd4EfevS
AdfHvCidiZ5FVyML9IaqgbdVpIshbaelAq41dYUNohDF8va9TEE58/QVsXhRABM+1khSQdBQD7H5
+Q4AKC5HHVfCyFWo6nBfL6hzuvr8H7wYH9rbQj+Imf0G4lLk/N0No8c55SxkeUcbPlwZyrZiLzCR
esV02z4vnPkhu3SaohVFDynUuSmIMqh1VjCBvSBeGPPvspSnQH4hqDBN2oRWTsZW/TFBZWT1cHft
eCHVh9nWBGpun/Bm8conQDOObouczOGS71MO6glLfhmqVf1WJUQN+o2dZZiVLWwxrRLBY4EmgMbx
oOFMGHcCn1l7nb9c76/yUls6vZxDe0koXXG5+fxELzh/eTXhyI8n8mziv9XT6t4BM6RK0NgIk6o6
6+dwKXLSksLNzIu1wYdZdDOxzVG3QB7VTsvKtdjTbZfADCBBrerqpcDM1RkA/V1UHMZJ/s11ydz2
50Hxy5zNeeDhGxwhuvo9sTcUMC3ibM6Vy0k26DD1Nm5KKTFapaK2fIVFFSLbx4DpntZ3SWLYsMYL
CqmNRtXv1kVhYgQemX8svD3y1v/YYW8Oe+pHbsJMqkgWla9AhtccAXN8T/Mt14xZ9+RUmjRzvCR/
gUMtfSLTrKvyiHcneeEgzoeXdVQQvYBFgHS08BUEuE2wq9cSgdMYpQGkA3a+o50h0fPJmZQQIWu5
vdhRZj2RHWw1UpBo8fa8iDpqhEHoZxaOAJYlIh75b/WxgpBUFXmxdKfvaEKbhSty2z7iotx8d3XN
kCgu1VrMn/C6u7+UBNqA/ldmHtRiKGnDg6ldDyVqCbvMB84IdwJk7HUqC+kcsfAfjeQyXYaRt5gO
9OMVLIzsJzaXyoYM5QdqIxJgP6KxX6MMvoao5V2hmmA7VvkbUuEEk7W7CjUIVxE0f38YI/CHSyBt
TVXTdFi9ZRJZfP3YBFLG/FR5KpYSr70IUlOfVwrwRJVnpwlrW5SBC8LfHQN8MapQJ8NYQsfT2u60
uHTcEkNLrDto2nv8UmrvBrnnt3ly2VZPQVG/NGh65TLNRPLrGwTf0KrHdYt89rbEwTcLr/NEqayW
KfOG0sdcfPYndkweUIoAU8/5FQh/jTs4/Re9LCbHTx0J0/MGL/79fqMiQoHt4VOWXsSmBAgH4Asu
oFzKBztqb7wnbCX/BUaoz2q3i5CUFZlooLXmgQIlI++N941eELMGcmNxLCY/xJhmhGKz8GjDdFAB
PVwywefx3bd8NqxPW1urupWCBLXvgmKLElvzmjY/+ShrDRafRncYQ+Y3gYrdP5c7laUpTRZtN6jg
vtyyqHkYr2Ly7j+HkxZkc8V8DvHxfglIIvnrQQq289XCGHlJ0pnh94pXi+P2EX/jeZdBSAsaUNDf
EUGXsMoBFlHrRspHBj4wS63te1iE9BXk8OkMv72hXqQrDBv0v96pvqKh9I5nMhNoIsPISNRmMPYF
YtPvPSh+JtGhNLM/WkeGIGARQ3kI+GfgolPBzmYqQkKZS8laWBpJhutOrjAIpUMdh7KJb1xIBINu
9Esz3b87yuF1ojBuGi/sm+2AAvPxkk3u3uDRWgYbck/Km3R4rZuK6BPHj5QOChc/5mKylCGecYdI
iSa0whT8NXTKJ+vC4hw7Ub+d5Xn4Z7mIetF2pkCSh+rEz7UgAr5zUAvFTOQwu705XZBmMWBqGYjq
izDdrgJOTjKOAm0pKvASnXBVw+n2nFRDIjjl/TosFDpWtT/FTffwUvw3JYulFRMTyk32O+KWfRQp
fY5Yep1y/ekZMz43RSCi1WIZ8MjEwlG0X9Iy0qZLV8/5X0Ntt/viw5sJFPHMsx0KICiUSXUU1fP1
Pmj+qCLUD9XKNf9cMgzdz6jU8TXlT+uu83Wzj36Oo+5JwAqv17ftgOhFIwhe4xb9OHlBIvutlbag
S2cWvd0DVbps5S0Br0cBSt+hxEabrwXs/AEFujBHZvFmhg0rJcouAxb+b6djWw5++zzSKp9AR21/
SPkaqLCQKUuzamg8MBQgjs0vYdJXxOI/x7OfewZMtUl+8ffziyP8tvypeCCGteDa1rf8WzlttTvg
v+OlVatGbtOyGlxxmXeCVSfG+4kflG0dC0Pi2nZw2Vieu7mEWXg/mwgkMnWvFSNuRzBahUQkx879
931iacHhjtlMtshDeHottkuBbcJhoMasDAFeckOXaI1slXGiCU5OIPXsVz+nMi4AsN+eOZoKFSPC
7P+o5JRYbWKlIbovSHQeD5ARaGvvgk+6MPle/g33khQIpvXDSgq3gNNrZO4b+2q8jak51YQW/A0P
DHw5Lu644WMPm+oTz+jmHNCqu7aukrFDbblM5cKI7OeX8vg8RN80sQY+cGsBpF0PrQZlT44F/Yk/
ydFgrm3ezHjUniSpkScyDtet4eBbfVTgFS66FFLPA3pLmnbuMTbwmxorvDEd6N+eKdSSCj8jcBUG
q3pVzT2CSTOCP+cxmucXCn+zWBLJWvC+yB5MaNMTrO9xBD43aT2pqi0HMnUwnD5E4DIaD3QDCwWH
sS2lbeH6HDZzDYPSb/xIYMakCO4PdBLiOSDIYA3N+eFTdCkyizCGYTQigH/amR8iHzU9egVJetiv
gO1GHff6hGDF21D5X1ovHQDwQhLmaatQnRk14J15RrDRXnZeaeM6/rWiEy4aibjaAKFz0VX4KZsb
TKjkbJz6T9eWduwXcLwFjSBLYDm8hBYXAK/McRCbzTUCFVKm5RBSD1kLNr+Yvg2EsYhYchG4w5d/
qMBlMcSBnEKLbZ3b9agsbgQTDz5KVDNSv7DJrG5Gjs06cwxINjG292LWaH920gbre4WhZYseZHLa
K5JEuLgYTGdMQ+2WRT4XFhOBOCacU/g8S5PWmuVtSSuWuGd7Vb/ikDJcLou48cdD54h6sm4xjoxF
/KLfwajzZXXhDHqwmq17Ilu5dW5Vzf7rrmjODtmpGM5TfYYu3y5//Q+bRH6RjdqmbOKNIZNUodJq
GMRsQqhWyYcJwlwz/Z0gMmyA2W+m1/lhVRH6ewiZva3/tfNkavqBHCYlg4fDXNPsfc3svZwM/71D
PzjsZaOysms+vrxCE9i4vvKxsZFUWcnzOyrMzDzSqhzAXl67dmgH45KdiXy9FMPphesouRsVvifw
jFBqJEtxG4BRrmAsABTjTNAlbLT9QznG25gLqFEb59+5V4+NQnRf9YW5bAikuhSwImzz3nYevKeB
BPSgXGpEp/o6sVoMJpS5QTWiZTuOWX27SdMFElUpuPyE9dvTU8BY5CkmfQwD+Rp53bfooXJjMFBM
95G4mqD8Ma0Ham2Sp6GLAVVVzmjDyIm+vgDRmJLXXrS7HoQAzlQQzsb375lnMXnT5o4ILDd82oBL
8nSgKeaWWsr96q7Rg8FflqhnlE9WpzYpi/ee1nuTq4qg0D8dw/kNPTg4himRHU224G72JblqA78O
TSm/NwlF7eKbMdDUqVLdyQ74B+9r8TmcmW9H6mvw1UgF4u5FlxgRvzV5r7mxTdQzVlCpfAMyzpnU
W0G2vgcoRlcUduNZzVWxWLtFtgykXeicBHBfYlqT158N3wgaiNHx77tqwlLpOb7Fj3vgl0BD2So6
IBAsQtMyFe4GZ4foqomZvxVA7jN7jni52SH0luJhBkIGyLkBRb96OzJnVos3tUITnyMsCIy63pvt
oJD2WzqYgjEQQKPjMWZXd/vdi4yLJXBSa8/Q5nS6nnKmCERl1unsrA1JsOgiB0IU3VccTAEhfHHU
M+6jc4XMRsuXBb62r7LbEB7xAM5fm4DJSc0lSVgt6Okc1nNvmO+9iDtkcO00pKbMSsUwIICnD7vi
BMH2ANAoZTJVNx8XBga2gHBBHi3ryTTJww9OHku4AiYifc9JTB1ZGfzWtD0PK9RK/Hy5uN5Fw0fQ
13vC3sgNSyFgA/g8roTQn4wKLSpvmZrzjLPI3rGrS5mjNNkrD3rIaE8wB8EJO15qd1w4EtjqCBNy
SVqERuzs4ENLwr0qU+ENZ+7x8CzdtCZXCPQk0ZmlRAf49WwlC1xYWcoizhCE98Q0W6yiDt95vmRB
6hublG+BHru98Zm5ogmrGfOvfY/fW5eBGYL2NVYaimJVtnQgz8wNgppA87hfuxUftTxCBHnAKyh6
2n3qrq22nPX2uX8GdEKeonUzLtWrYSz+OnIfivl5pXOP+xjDZ9LCBqMpJkMNFg0C0qBj5carXuud
Bpq0nFyD1n/2Y15FV70gdtdG1Y1w9IQhTBYeuecxbwzSGrUA/5rBKPGKJG7ihfIEjRn34AtTX8F4
VXNkdXFc5c3GaMlRrVkKSzdCtS8Gycq6yNiV83NaGK1C1fzg84MbhNpQWqAMDoYcIx4DUw/wFi30
aPmUQGMi8Fh2yaDF94v0D/pRtQn55kdzSAGsHt3dQRkk+LQhtVUyh8kn7JCiPJO/NcQRnniVxNHB
csgRE1MUvUJKjCdr65rM+vPrIBdqjMaLJxOLRkh1X3C6eWyQPW3tvtVXsd5eNCm5lRAFb/Hom3sl
hLROVRGEzseBS14SileiKqWy6S4uUbWKe7wh7yXy6zd/1kZxdcFoHvx34xVWM/LtRcbXn1VIMwwj
OFQ1kVt6LF2yuXDWA/5Ju8p0VoSt75acSpwWuF9hEl2J68Sj3OHtwV95lIoQFo5PnfqPCEZNTOV3
MdqwTZNU4hZalB/YCaXfX2g/O9D2Zz/xi40j4DkIV+1miTouzNzKNHASR3k/j+RakkbIx9ODnxPM
Ol9F/Bc10kChMd77PGgykBvE1+sHVTYp8SW3kqDwyvMwWsRCqRq7yCIXJ2HrloTPkNWxqRwJOScS
Kt2rnYbiv3R+il5EsIjwbZMQdzxyHDra70VmGVSL2LCt2Cf0k3rwYTmP7XQlYgR8ObAbycp9vSH4
9a3CQQr8jjm2XJ7HIvfyVSgtWCyf9Pz+zPK1mZh1I+i3wsdzkleUxEHpp8XYzx604YUp+6x4345Y
bKmP0cY/pnuGTFOiv8HtXGECHE7AYWNI+skyiX6zkW0fh/xZN2GXru7F5obeoaiIWqNFOkWKSK36
CtUdSrSaswns9jP1I7jIJGcrZ/a7OA/7PxWClgyGK/lAWdSAIzP1xcEcSpsTIS0SXWRqigkrNh+P
eVxgKO/mw4Yxik/hiag9qttxEYzPhRvvEZwWXjq9Jo7S7Zk+twwJ7X10qaCCh/s0E1lcM+A9DG1U
gmPjb7Mf5MfUMkDhItZEfH/H7bsVDeg8JMj2QE7nV02rD0jSdu2ch7n1vVYJpYFOAH9avYNzZmqJ
qAV5jOVw8M6gcygzqRSiLmLI1DXAJT7ovPTH5RYHEh9TMYMEcNpVtgUi0zi8DCq5234wt8bn9AGY
TzycUKwieJTfiAJZz8HOVwO4gNXFM9K/iUTxjY5j3CjEsCyKLNO4OpVl+F4nFns/qMr95N0zxwBL
430gWWK875iJpd0qmDB6lvvzERBUpiHvuWEhe5jhY3brS8qRQHFMr4XiA9AP/oTqtoHflCW9hP2P
MDRiP0wyQWnTvh2yixu6cJN+3oSMAXXp/ODt9S0C3dY2mBr6H2aeTPa5rDfRZAWvmMGfS/4gZhkI
hm4Awk/GLjgTQkSJNLgOqBFjYOt6fIbA5yNgamWb7rx01qB8DgonDo2QnMcuwtG43n0KXtAV+uAh
KCNZVx0qoB4zOPRpk0BdTo0CoIoyZI7uMyrULONrV/yrgmAmeRpTuSlfp5NOyuTUXl0BRcul9iT0
UMFRDp3KZ1xb0ydDfZ2Ue4WNPWpOuX7RFO+UfPaRcGfo7WNy9ZQjqAaNzhOf5+wRaZOtz0YB6L6r
THTlNhoJ3jQkCxWrafDqdEhwRuKAue3Z4ZfJtLk+7ROZQzhNBgKLjzGFnlbgad8L5ij4f8Le5Y8h
NCP2vq0Vz5ex0bh7kZkH5AMr9R0BJFPQ6mqko90EPevlwDIGTm2SnvU28y99auKRfPtd7nnOjoUK
7OHtfMV7bwAvII0z1aQqHD8jqLNZCtIWkG0O5SO08ESAXW5RePhh17lf/hzSLp41JTF98sQonfWe
XsSeubejiiHZZN6+rvZSj2L4XV910txy7S7mul27A6aBGaGxBJwC+xi/P4ObA6CifB6Wh2kKx1SL
EeN5rPlvicI8XXQG2ztak2/VO69ApP/bx2Gz9YWjoXpnXXpLIksvlUTJV6NaNVydHZ+fFip7/QCa
19bI8BOwClvXrBMFMlufnf6AnNeQLMNIxPLnsE4XV8pt5Hks1R/hbhlX1xkiGLtNcP1O/+j1qfXF
0/tHZoag1nCwWJN6HspsLDIT6VEj5BdbC3hL1poVc6ueJGTQ7WPfaSq6WBNqWz/FvGbtOG2OGS+C
yIpq+njGiPXdIHTys1hI8OaoZrcWRmgLIMZgD5EzgkpwccrqVjSeiK8sqCCWP9iejXWoPRpyi+Op
7amzr23omPiIZqalFLSsLgYcGNV9ht7GYQJvKEN+6nisa9LZX3/UGmu4ana0wD9sRxR0lmZwz4fv
EtDNgBIB4ak6A1rQNVuLd7sZp44CJFhw7hh4fj/wnLYdvYJMjh9bZr/QqKZ97w++kOoRl2q30rSz
BQ1HPXPaxDxlNkJLZ/Lnhic7mwgb8vwO/jaQo034CcMNPO7wMQ9S3Anb7MWUJ+xxJ3N+Y2FPeVwf
MuRvbMDrx6CoamDaFCpLLeVqkrglSG0ausgwWOiwLHSuiTezihJxRNm9UXO1+Jowvmg7B6q2NhVB
qPLWJ2hJaamqLo4YA/uxD9y87ROaC5UW+X4sYbpgaBSa+Hjg6XJyQcq5fFnR5wAPIRYn+P0VMB9j
sl3glr1GyFLufdI0pim4bxOlMc/4EvTZGdATPrI36cgU86ls6yQr3f3cyUNOoED8Ug2Y6a7xzCyn
Ag1dDinx/NOW1Fb4mXVL28Hpjp+lvF2jWy1eN7xsg8iKL1J71vcGo8uNiCwaGENKDhBgH3tjRFHJ
FrqrEJgf50HvIOvD3Q5rhzckbiGy6K2WXdvGqRoQ1OqrCJf4GWfQp913KOuRuaQZAzBNhkfjZKxD
R24jH2qg8mYz4kzfznMd23rDf6rmykWBIPgBLnmpu5jv4d4fV//MW7Du04JeqjDNIAW2VmSaU905
JkYJ7yv9EAa2iuFoZ3SB18A3MPHZeSzpw+0f0QFgIO549g5HB9rm/qpEaSO0IOYrrovnKFkDLTv8
MmOc77bIVj0tadePaXNRAlpgM8ywVLASE0iaptTThlbm1XYWgk2QjHYhkmo+LR3mHfbIlJ91u+I4
ntchnLulvFgXRKEUA074Oy/DFba3UFxW0UFWqT431fZPWUWuevKyPy917lGTUcHhEZupDHcbkHzx
k8jWBpGZDP59dLKCKiR3/7a05NY3ZKX3YinkxuiQ71qfy7CLQIpNOl93kphDCBOtYx5vC8HTh19r
hRpBi5hAftHZh5rzHNqAt2v3VYSQjXZotVEIGqd+NYrhSDbMOe2gBqX/g8KRlOEXf7ggym0JnOgw
xl6TZi59H/Q8Ocq4e6qxFe0TtfhoJJSHgvzIOmIE/Ethd26Vu841tLBinbkUUM8E8NsuHGMLv3HE
6c7g8uScCCY2UpCkNybYeXmfltIbcNRNW3YifcPpo2l8uH/QwVJdCTEbPKnjPlCotMiLbuWwuX3P
r+M/IVLBslMSzoprTdpucLJq9DITZ5WUe0HJY5tjWG/H381EKvxAvovOcLdlK/R4B9PTOsv2h55e
38I+jjkfIW566dz6RJM8NlzThOX1pBYP3oe7I1t4QYemCOQyar5iAyc1h/5d/M01jLULCHfh3sBl
N5z9kBEWlgCif9AJl9ejCFOQ7edvR6Q7Hiv0QsX6yX8tZqR+opRwBTeqmOH/7Ud+TMFReJcVgIp4
35UxabO7niTk2crz0cp+Osb1vpnbeVll9dBd50nOE11NxXfu8ieqlYoQ2ZMRhPoQyuxj1S86IAFk
K/LOVjs5wrqN1i+8Z5vx0FICBb/mnJK3+k83v16WvlEqH6Qb2uUUbb6v3iU/9cstPtqf6mUzTfAX
/TGvKOsCoYjilEdVTRy3OTTXCTcV1JWiD34M/zDoOIpy0fAvMPUyZRRBToSwljfiFNYMY1xdVQUV
fZjhcCuFcKAYsygvUYaw065KL2brutyi5Bec+/v1wWDd2g9qpoxRoq3bfW/Qo8vJX5/DCfSLRnec
wJFhfQ+SHCELQriyUosbozDO8Iw3mjKZjV4LF9ZtZGpcxltTA7/qLKjmvZYlHfaGS9Dxfu8IOsCq
wVqRwUdVVTioO7Jca3T6+tjmN8hlNA3UdA3BvAs7/6uHPz/FzHQVVHtBDiM378GE3vp6oXaAvyHO
djateQga8WyQKJDK13Q/asQobA6rJzpOi+u1olvK4umLc/umFgXU9XnFAj72ZZaOLX3xnTpQCSgm
HNbZ4H9r4ae7uzdxdkEKbxknoxipXfieK4MOMXwxj9DAxPcJUiu+a67sKI9lcyKH4gPVLSgh9q7V
Koz9bJ1Uo4rX4PSX6ceSk/xbAQ2Unn9w77Y+TXERYXLN6EtoihWcmhTSgCUwytz8fJlilm4cw2Sc
IrZD0XUjlc7T/LfeDnPyDdud73E3+gDI6zsns6cTa4zEUT2iaUUQH848Z1A3R0IUo0VzUgASz/We
iiKfRKSWamvExJHtLKB0WW5TTrgt9MZ/sbafGoznqLOJxFh8Vhbmkb2lsaeKnHb0cl7I6eOuRtWV
Jc3Ibun7MI6lc+D4KpwVZZ7WKAjvq1HDoggkXIu/EgnBwq3zQrLZaqL89EAbOehepwDuL382sLG1
m4S+1Q7OkO3rbU+XdWC9HZEb8mN9gCWMwEAgAUt41LrpJHKJUKK5BGyAGjksjRGIoh+fRohqh7n+
M1FcAGNTuu0zh13p2zBGBlNMB7k0m97glC5MBFWh2NrGOESu+RHFPTU3ughESlonRtGJHbhakdg3
ibMIMPoDrBUjGGbT9Ry6/yXD/yXEy4janKT3K0hDynDS+NVNRjldsiAwDIa/N5zXWZFDic1msNna
XEzK2sbaERvH+9G2m0+/w9NNV4aG8kjhO7xTqlpa4BxznLgX+D86KPEMbrSyn0hSaaNA6GwdBY+R
MKoSCXa/WCI7XmQHAUJeOJK2aN2bks3sjOHFjJYzJ2tvQyMtjlig+dei6bfoucNmgatEcyRyH3jr
CEEfMU+aU280CEAK1EMzdXXFxcHA1c83/H++HfYqvT7Lf/83eUwE4eMGwZ4RllurBtDrBoW2RShc
ykjEFnIi4y6adh+QEYJQ+sE8F5D5PL8tCRoWTBL9V6eErSJkHTH8f7RwyjjsGaN1EzmafJUPOzQS
4J4c+n/WvHs0vZixDVxA84ByI77iBmAk8EAOW0Lh7u7geWPAEdPD3kVmtxoypRYFJXA8IGF1EplV
Y4nOix4szT+u6zFA7LFBB8XxNS1zPu/IOEhaxQ3NUhbrudBP5nnsnq8RyfMvFB/akLp3+LcFTCge
UymPmE29lTMitzNHHviCU2Fw/nIwApRlfdtFCcmrRPtbEDHAsXSHTLG7IMR4/kPk7d3kBF0o2bbH
TL30ajZvuwRIOouL7NpR8kSUditcEd6MN+vrekCBCQnkD73KMRs6Ynj9moSwlHfn7JzKWTNS4KA8
evTZoI2/twa8fcUAXKRp4pDMmiYWhDSE6/B+BdKBOZkLrBrueG0f9XI84JyEsDB3RUl6sUQZq0HQ
/vyJeKdcuQHyLHadVo+vE/9Zh44pHH/RKka5C/bVHA1C7twqYFjR/qas8WHJIWWWQB5FI1dQR19w
LbyAK2sRPOoUctYfX2qk7hKqI+p54KTEmgQ96oL8GLMjxXs6GrKN4wxO8g==
`protect end_protected
