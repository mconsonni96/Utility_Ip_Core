`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
PFfrBlTYim0paCa2J3OlpWc9Acy79q2hOWA+FV+QjehGM4wcNCFX88yMHb/1BZRFSJ3248CeT94p
gr6E8rMPBKzi4hquWbR/LKv33CNYUckQESwt7VNDeNrGCGGZsg58OQTTGgOl5/JyQIGeEgrkBajJ
kGiMrFQYl+VmlYu+yK7C5mqoiAe1i1g0Bff7FlvVr2IHC+Y1DjaBoUQN5gmtqbTl9Q0awOXqoG4S
b+qaHTr7YRacdxUcmIQDum+nL913lyjRgf3erhoqTu1kdvqtNhck1V+27gmWYZX7zN2QFl8/khT2
W0EbPPiJQsTjBeQe3uc6N2GVcFYFeFf+YTVGmw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="tMND1DS181b6oiE4PzaYPwZo3fB76963D/A7lbBwg/E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17696)
`protect data_block
R47xKW742NKLvZn0wMeA7+Xt+7g9kkGolCh54JvJKF5H0RDjQgFh/qYc4YKqF/eR5elmxOGX9i3Q
hA/nSjhrb3XVrOJK5j3KTWA7DLa15tyZ9GKdow3TG0Gm1eBd0QewgK3ikDxhIp69rFnNaFk9FHtH
kakJL/H6CZ7g86m6zLm6NE3m+PseCCYO6U8VZzoT8fTYf8DnTKgLJCwKDEFzgd35D2Ro8hCK3jgK
LEcN0zY5ybqnrqfCC2FXy32q4+F17Y9vmZxEhGUFz1wMzoIoY48AP00fmqE7Ryeca/JjF7VzDU58
1TVKqRo8itmCq9Obrg38j5IPzGAyz6qE1LMWIxz+JFPeBAULAh2fA0emGMR15qFV8xgGMOZ5utd1
uaVnkv0KXmKdu1yzSa9z+FNue1BSqJdZ0T1ArXwAIgl27VeuPIrg5OgLZSwl7rPRhTTBJOgbVPhg
ZYfwL0m8kBcHstJiNKt2e5dMefwhITHIUBQzxSnNT7FOFP1BFB8pIs7HZcAkpUG7fXLrlQ6BjPNJ
rp32rJoD/yOASLNttfMotpyMZP3fgXJsoZqYRbELnQc9DRQSMffq57S+YtzjKsbadpn01oRId8Tu
Ij/mYVB7TVkKp7PPUXGC0Psmryltz9B+cHPko1szpQLcVqMtXjMjoqDdVrueb7YjUzmEY6ubA5Se
CVzBx9H25Ngsc6B7PoraFt0tlEYU02QSoLiVzh1T/4bxodcFPgO+zj60vIN301cLIqT1eHwvm7xa
xzeXNiGBVNEfMMY0+ZTV3/wT7HltNGECVbcV/Vi38nNnkESPiJANEPvk4QUp448DvXC6NmFdce53
qMqK/OjEmblfGqb6bP2o3Ck8jInYGSO6bN76fvxtVjrUmNiZiCskG5CpCV99ZSfI5ODh1IMhvvT1
qCSsmWUTac3KBxkP+ZJP8ubpg9yX/Se6XUr3iI5E80Aur/hd9HQM6d2+N2cC2PFYkj5BfiIwLNtz
CyQ4PgU07tnPUsv+GdkswYHQQKIhFbdy5MwuqKPYFWPpIaAFnXYVCZBXkIWJ3fQg9pfBgCYGJ810
ujEnssMt8r6RNA/jBuZCUY4hceSmr83Vo5NOLsmy1qn6+wrSJ24BY4rMCy84WchOtNpi/IvsvhRW
EVfsOKgCxQNVZN8wvC6naKYKjXS1exxsV+QApBfoGDFYI+iUNnYxx0zgf20fZTYu+Pa18v8A6DSA
dvUyYcF/MrH6EPt6IN68gmCKrq2Cz5dekzo3GmpV1aHMMtw2JsDT/0gVpc7wO5W+4t4I9AoRVIwn
Tdrsmp0kSCKw6C4Rp77XelDMywJn4kv1j5w+sDmYMsjOuaboOdk1qwODBQCg5MoIF90KLq7KBO+i
dOC70TdO4A2B3xMALpCyTBSAv55zhpmA5xGIh2Lrh0B+zEAK6vUSaejep5MjasVBsmud5BMRA1Rm
KeA69hbTSWZkw0UB8fAjwCukXFK9ia4vxRGr7SHFLTxb0poxwr85wGDvlRu3lkRGpyeVN6fX3yeX
kBKmpGDfR5qTDROOh1eTz/twEHr3yqLdKROPzWd8X8Zx6S7bgCiUJCNgFgPxviNHABgHaPOB4rb0
aUlBbEBvKiBnoJ6/coZO8fCI8cgETkkDCQZWWMU5V5+WN9/kJqFQvP+VKRm2dunAJ4UjM+DwssVL
SUFv36Ls3ulyRzaeBsXyVtzy3qxZ4MjOrK2wfEtMjvusIwfUw6xSev37suOCzlveStolM7KwSk0x
CFg7jcSRfIph3DzX55kmfTtEK64JyG6rC5Yk/49ngDaVo2n+zNyY/m7A3BpYe2Q4UVYVg1cWvFZf
Kosdg71nwXWE/J2qp4WJE6U/zZmmtxX4M+cftROpppDB+GvDWSoa8if1FgoSbgZ7qiuq7ytz2KyM
8jHIO9+y6fR+EKLYvd2j3XRKeeIkx0IphnH27B02Cmfr4H18tpDi2Sr5Gu1GX7SRGfOZ4erciDHK
1V/O7CJtoHVzKT8iH+4DfgcQNDt/PtgOtcjaaJbrJY1Pc3dx8DKWtgnXehBStcms48JF5bGSA7qg
5h9so8WL/4W8FXsypxUGNfren4nOGMlq7NFL7I52hzsMVrkcn0Avz9LnZuvkuqxj4YXN8RN1dfVX
3mi1PWeXuYxrghw3WtWSm8lJPqZ+VaeelBzDvjqN8sQx6yKyGFEjBc9QQ7KyIZMgMZjAuQ45Pxan
Gj5Pha1XRD+NH97t/mH4FmFHzke51GSITMAodHS+LZrQb4cZC/K/Ak4+IV4qz0rdgEFKrDDgriLf
gb3sxW49wg6WMLgoX6wr3+KkVwZ+jL977WBfFxGf9LKDEhr1shy2gP47pqSbdAORa/K+RVhkeGsP
RjZBA/muilP8s7Ejs9ocZJgvIkEB4QBxSiEfIubVmUC2AcylOu5H/lYsADV9ikyzSrCL0zs2IXfG
bFm2PIaEd5HZUZcq+MmqUwPfF+ebdInK+zfr60Ebr4w7Je8E1jq4jgGzokwOIzMvjYzT8E2VJfc5
HvCOXqiDqm0dQEmovQpzuab4BocmMOT8IyrQRRYZOUbqLFz0Lp5JbMpB2d/375pNUqkIW5QW3nLs
tca0kRfanYUUixBrlvHQvZKE4dVdbv4NN7wgjSMrfqYk3cd1yzBdwyJHmAtiBvfqP2LSGnXNd/Fx
doDIxnDWx+zyow8Z8Qx0hpZWcc+4VQt+HfrSwSHl1Yi1hIjk+TV/TGE5OX3xErvTffVNaKDf6D/U
sqCypF88m3TXYkh8ej3jCQ61SkKFU3IOI2G/94S0pGeTEgUYQsvyI1dKFui44DHke+Vx0L2K5tMa
LeQ6SApN2tcIVeeR4FPsS1q8kJCjrjFvGklZ9UYGY66mCkfCjm+hB/aSAPjE6tpAvnt7Dg8Yr2R5
lA2kEX2UOkV7VOFsMMLS861qevATMsLBK+ret0yBMqzN1WiH5B40MZAe9jSHixoiHri7mRjjMV2/
A+po6EUrM66hxhBZynZ2gqoXLtwcG39s4+VU/M5siFoh/v0lmdzuEE816CX7Fv0SNI6McbbwddKh
wH9kkGbZEmUCRsRaEmyjSYQ2M8v30TXb7n9isyrDZqT9qDasnfe78xQgdROYkTW9vl+YMTpIwZIz
pJiwzfO2qkMUqtNxQMcQ4Y3GIOqEY78tNoBBCJDdZU//BpMwlPrYoDb9ntkZi6AU6UK+B8XD9wC8
fSm2pL1+cicjpiX3w+Lk7gO2BPA7sCK+50NEQIxdk9NGFU5lmK8roqa70k+FEIKZW6GiHMdfvVBc
cHCXPuEyC+6+VHqNc28RtrQRWaLnKdmJDzJwSNM+3G42VvpbxSCd6cxqEeVlHnfSckcjzn5cpxWY
O0ZFatc5S6zr22JoCc3g96edeGhMp3TQSF/IzYfiNYqhJ6/fQ1vObWsFZd9XHq5epjroctiDBSDn
ex+L1MSzrX4VaQn5k/ll3vB2uMYfa1QkPmL6ZjzSshC+Uq+x0VM6mZISC3YzrXM0pk5E/73hDG+g
6irOyITzdN3IDF6R1f/fpZZXcXLoOYSUHFNZTqBlDS3Aquk+vacbc42aZrcrL8aGIzN7CygiPN0k
uBQogjLdO1Hl/vtOn+H9QnkAGBvWJyV9LZLg1knn9csNhNKy1oxzZ/dI8JrMjXOLJdnaB5+cuu6T
wzpVFhkVdBReOK9f++vY1g6GQnBQOJAPj9Y6lGRe/j9fb9+gseECiMf7NOFHFNMYvGb8pEXyUg5n
gJTZiIs2e5Bs1UPtRjLEsf0NHstmEA5VVD/JvpFBqBX2rC6bevwUyJpqm4A1jlaKFj64c1smvBT5
2t6KibzW2tZdx4yLxq4/CojkW9JQF5Ih/pfxS8F1vkZTvVESDCNYNjM7LSIXG/hE2FW2SC1jvu+o
010tJ17dlumef6wbtdO++ZKc8JSPRmYFgyz5XOtcEWsCUB4CTswPhuj9qQmYkmkpJOQY0Jh5Td1T
gWbX+ZCbbDD1afb1PhwJi9RNj6oCZtzCUg57PcptW7GUTnJT5w0Kg2ht/h5JQibSGjRMNV2t/O4l
FJxby/yWNl0DQeV45+wCRE4nskknEi2zv3NObNmw7BXM+fYx+TLuzbBDZPed5KQLB9WYXSqEqEwK
KXeLn+kx8jwcWxjosskB9ldg1IWdqkJI6834HaAqKGGWVgfx6lk6rJJMx+flNnXuzHltwLp52CkM
mKkI3rfPnGI+iLv6mWAcKacVu0KUzbuB0kDPu9GEJ7v0Jr4MDBWFl+a1ybJCENPIaA/nqOtg2XgP
YoXkhh8GbmID1s8eq2eK221EM9+RMa685sQ8h8IPu55oPz8VxRGixLBmZ3odWPgLCeo0VG0L01I2
6FOn9j9MAPIc4ihgU3uJ8HOSSHXDs4SLCHjdf6yjJNsKGUDbYocOC7iIff2431MNeEPj9piUeXUw
Ito4rAvqzKXMgcu/UJ76sAdA/Km99ojPTQ+575GTKN7fGNzc1IqgY215lK+qWCmTDntTa43/6Fv3
ZrYT/r/v6qctsvIjVHIfexP3F7DZrWKYF/SwZCAyNnLmKE70Rrl0uK1DDaejFzfN9sbCKljFGgMZ
NIzS6OrDTOtjO7fyU8dKTtTrQuiK0wX3eZ8qQ3Q1Gz0p9YZyTZsTxSRKL+an7sra7bcDzy8ea5OH
UWBkHvlEpGnowaV+B8KdzSJTshK9+p+UhcWqjdGfUb3EDK8HTaMOAoHcsDoYeqcHD4DG7hqQI/ec
NFFxKEKElcgA/j80PAQmfFd/wVZVefdqwDAsCMiMjTBf/52EbWN6CYkkcpU184/iTF3px057WnSG
LHHTSwOCWZG65ghjG5FkvDOJdTddQDLAzMTeoOZ/7hdsfs2QJyIGOJI3Gxd9SVP/ZZGggcRLat04
AljDoynV682NvoBbJwrkuGWPvbLVKf4J+ojk4BSTyTUnpvik0PFDJqUmoo/CTPdSE9fMmBAlj3IA
VnBr3dzrvN0S0+UV/PQe/YMNdPbcyaxvcOoXUASo56VdiWHiwakDg271L+SL/WZzrK4MoQV0d19l
RduMFD/5XXPSBUr2Au1gYG/d5ulvqp6kGgxh16aUXrkBd2vFPSAzcn0kQqBWSEglI2OloBHbCvO3
4qreY3EPtVkNEJhzB5q3BAHmtcCAsoSgXiWyVv0VeMZtKJGENoxK6eUNHgnvZWz93juRmzQHH0Yl
3nA87EkCTv9z2hF0DZVaPMKQSBGwmr2rAPSLbMI8oLTpn++HwW3s4OVQ1JTrrOt2oodLWUyRfDE0
NeEJvFi2ZNFTZ9Qr+dDQ+R+JZFBndTd9HOgAbSk+pAyuVjuG0+KCiIlYsaB7n8Ddi//PelEDgJMm
T3IZD0HlqmNjHG7utFC/uQu8u4u2+mTbqF0/cGoCI2ROiq6o5QGc8G7b0TdDYgVmHyu/6ghGFTSk
k4/8giHQD9eK/v92zuFhbv+hQCUZM21+vWtLhRAE7M1E9kW04CfRZDaJsTXATXWc8rtMC36TcQE/
7DFHPpig4tx8/jHCzRZsfSqMqd2ha0nW43N+7kjM+9nwVksRtLEpUiLsh+XM7MG1u8vwRwrrbTQe
NlVsSeMkC1GDulW30KbzrkDi4akNcCTo5OTbMdw9P+tASRH2YOEZ03B9rtjueY20PxQEKvcxj99U
x+CCeUsZIZ8q8d7Pn/ssrM+qU7D03+T7K+//bvkrBkfxtybLfoeNbaGZPNdwQSe516yv3FFV7mWv
BJKhPNZWlQONabLjh2939dXqwGEh9TVWb2t2bId3G2I79GuonuGKsO1oiWU5Pdx1j5Zvgy5XF3xx
4PmWmHrjj+0hkoXiDTcp1rjXX7Hc+NCue75zJXI/WNmNU3iSDdDKLDOyG2kaPXygLQl/WoP2lV22
ZAJBnxBUkcB0H+2zzORwEAPNnzMpJvVhNpQwhpH5Tl0BMfnJufL0ONuGClRgT4Pg3MiugiYXS3H8
XcWCpRi4BZlXEYTEOV4SyXxOb6dtneZglrFjGJzxx75B0IoiKa4VqZts1MIWoKhwmxCslnUQnk3w
mbR98xyDLpV9g25T9baadl+IjKurtjigTBdy/jABNgPE1hJpZevYv4BXcysj0hkaIwTikILty2eD
CfIyQ92lLB/7S3vqsO6B/ypJ88mG9NqTjziXMm/wgHGfFt2UgJcKM0QFvtQKxVsTEEmprCaac5If
oDg2D5JlhmueAfxFM9dxmypNfX0yV9ohZcsU4f4mNfhT78CK+9huLngGOPCV11oqwUdSOim3MglM
FW/voj5kBvKtWXiF1eEdp8Mj8XzdxOtvcMNXEoWxnOT84btmXbc8ycXxOdrKkrCeZ+w1DrvdpYwW
m+vRSy+GiwKBa2AHBW8qMiNotLbuGDglL01R5b+zItjtP6l7T+a0PRF+ejAuhR4fAysoxRgBLvHB
tF1eGdLbmQLieLuvodNs3HCuQubUcz9zmHBToWRQ8QUzkts1hBRSmh9DWew+gpfFUQ895pDN/3nK
nh9T1jatpCbZktVc7XfyqZVGmzfnpGnb9r8cO48HGs+5GWXr+epC/1IvlsNMUieuwOH7taYCMQ6u
cOEmIgTdf8mOOYkbEQmhunZGrWwT/MyHb++wVsk1IyZNsa1ENSm6Srre6p/HjH59mEaFB5DtNMnt
uci3eSN6jilkg5iWhutNOLoneqlQjiamzbMhBRzGA68bNiS7z4mpeFQRtupgXVQPOJDeKinCUIiS
DU5RqyGY1Q9SqYbUF8PKo63+TWdCNC8pGxkOaH3YCMDtBWSzWi4bAIJLSKt/AGp8qmuYovBor0xU
Rsc2n51tEmCMxQCthAoD3eqXL4CAaeYL2rupFpYO57V/Qw8hlTABWtfZjU79VuHKmKWMkzyqAvFL
D6Kj88fQ2ysTA5+h4Y6EjPA4ojPDwA1qWKM8cSdsWLLp+SGr/CHMspNBdzuN+z1hxuJQNuSu1IIk
bPxNtIfbl9LhAwBRBbaDVW1fHxsJ2zSvMVg/lfgV9q14Jv8AvXsswZzdsfTSPEHD07gkoao/WszL
3lDYsBBzkUGG+WowTkq7WMWKyXK64QeBD4TKwEDkFAvj3wMidk0CACW6RH8BP0jkHg56UUaEMvLd
2PJ+RvpaYRxYePAtYak7OC9UaorhUzZ+ELkkHgVAcMFLu83VtHhgnIDOcECacVFj73yqX0kpvXbw
E/lQRWrT55NT0vvBT8QE11l7FmJ1hQEvSvl57gTA2vE5QqyC0d6bm2natFUI1sbHiaoiNeEDSn+B
oP1OsTZWJElbWUPc+6ZMzrwhfW+nOjyKmHvM1aWyx+OhhThZTkQqYe0Vml0mMHwN5EL2e0/xO5x1
G9EtI28NS/gENTyrq+8aJk/HUoNRRN7FTFSaOeQvmtfrSuxOHCOE0XosXzeWxWh8hFeCtxiw/8B3
gc0gNghOdZmBxoCpQ5ZVpEOc9TY61r6Nm5lowZDfwuAKTFL/vhHwFqL220qo3SoOhe/Di2SUIMvr
WKJoKbbzzyMVRfFG7fbi3emLSTlWt8CuamB9sbabsnvIGihqVIovmbOdHS+aggRMvlxDdkoOcEZr
wi0XubXkyWyAlykLoMsbSn07Uk7UfUoaOSHEdfe5gbNCZ6VWQ0SFpiNP4+md6+2nl2ZZ/7CcL1Eh
99thczeM7ixodK1Qt9khAiszIHteriQnSwz+becRa6Qf+E1rU8Gi7zsptZZOjd9fLItwJzLtXXLU
lnnHhcFQsw6VjqmBnGmccUL4+mEgL/dvMH+hy4v4CqZwNjIJNZoBecfb+mLf0uGRnwfS526VQ1cD
XJ5Q8mirxVTQyQz6A1Cg+ybV2HXCF87ULEXOVJ+wK0hBAn8V4Rv/u3Ec0ag7CJHSu/Xv22y9k+Kh
dMDsPeCUZqM5dBMHMyvfASPgOVqOJsHos9NwyFqsD6mDg4dR9nxGzDlXj91Z+NOokI7w313lMs7d
roB9YNxgdceQdpsPFreJysJup/yJ3tTtIvqy/duvyLMrsxbyRFrkgJIq/qoLH788beBvut/JUtHU
wE4IX2LuAU7q/qrsHy2NusCVv6RqySeunthd2jgq1Y46msxLgOr+0Y3yJGGs+jN0Ql63DawIM76y
OKubXkjFG8cVQ2vgQ4rVU6pk7LnoeU43pDIesqzy4ATs9yRx/k5iJNkUApSGdBRS1TAeV1v0lkBS
qQSoiT3p6blj1RuM4AL0uX6BrOVBczPYy4cCfhdxMYzNam8kQg8wWc7ue0PZnleFtlODhg2PPKZi
FXZ6FqKlwfoLEqJttU8eERflcFvaYxLuiJnpBTMOeYzJkXNr0u/ZeVYFzUWzalQJzIfOZnQoNcD6
P56Xa7DRwdHYtiOvqRpBRxPIsGkLj2dJQh4iL2MhYVY0Y6Jl2khE3msghaKQf7fgbjnEKZs1/Rr/
kbvkMaDZL7/cW6mglW2rGAI165OFUGi/21CuaHqtuXF5aJqsTy7Y0DN/frrDaM1hEmDhG7Y0Z3I9
fuAsiMYywHmiBOONoLbXxhWzVZHbp7C96N3nruyZm4u/6Ri/RC3iF50CZlMKxG1Djh/HGIsuGNAD
C8vU+n9PJclzWqvbOSTwnoqq+Oxr0iGfT9z6sw4lMVruZKPfuXr3rUPH20gz8UKxo4iqDrx+mAQQ
OiWAGGmByVTDVBHAla9NZtZhVXcS8jO+bYDqSWq00bEpY6PPFkxYeSz66KLIcwiDtVxwh1EkzfHA
I40KKaf/Ib1rrPPiZdD8+5yPnftX3cJqjdITxf335mAdBkIjQMtrHxGw1VqrS2rsSe9Pqk9Z9VBt
wmgvb+Z7g37PdVqC28RqkoODF8EYLt+7FwyoQOk4hO5nDCW37rjK9ZnKgEcReyz0AjwzOtW86DiJ
iv3QdwUo4xbpxnYXjYgeL0I+FMf3rhdRjXtAZi9aMeaQcUtwo1BplmfjnYKFmr9SkvlKLMIe+UWn
7IhBtOZwVzCCEAeyR1+gEcYX9BoZmHZzZBX1GBCM+XNBK+Ci6Tp7FJr2wbjqCxxYrVGkv/GGEtl9
QponwcRWdB2ALF6xB7i8CbyhKRDIcfLQlj8LKUj81sVpXc4vDTLKRO7Hrq/qYbzeDnotgbWvJm5H
UXSLKTCM8NnWGsRcUYXBAWVPOMOx3L7SgnNFh0MCQ3X8UHnFQNXVQ0R032uWJmKYJ/tDOAs1LgLc
UiCIlWYv4sKDfVVtK4IIj4BvHaserwEnnxb6OAZyB3rqvi/7wc20mOii2qTarPHGjEX5nTtVic1J
zwzRIjla7rpO661cCklW/2CkiUC/EkwCwNszcPHZ1RW6SK+TnqjrYZomMrkVv748yE5yumnTvwN+
KNNL7Jk1V8t/smvLQ7mqXZW9jtS/mQbFoQKPdneNdxiEvLnM+/FwuFoLYVCN2D0Dz5MjVMy70nE7
afAXG6KEa/3UP5+sdh+Xbt5RruU5nYDfkMQKE4C85tFku8+PWxEy5bKIEBoTJww9wTKrEMdDDk0a
890o6WiJywm184x7wsIbRIwfRGJyD8jzFC51oWp2pkIhSQldCTNffXJ0Nkw1SVg68FqJt9D6tst0
sy29qqgb+7uLoaOMmlO3F9wGU2snYZGkDmXCc4yHh8GoMmBVXihrX2Xx3zNk8vf65s7/+8TlOGpm
IrMjGdIgFiyUdnBxGvCkLCzimf5GR17xWvHz/MoVCXYR0czJGaTTIp3zBZEZgVRXbDkmy9AD9KzB
Dtgts28KI8WN8oEDYkoj3Yj9GbOFOkdXGN5a/9hsYwG+tsRAdzoo+64vlYJL757Ah26Hre4dXGtu
5NDBoTJOijKtCZz0FZKPrCQvt/MWAeZnnUnPPC/XUaYL2zl4lWVt+rfRLiSbXoJIUhPiFWo2QM/J
Edl+FND8+NWjIP6cSd4reWoPkXujJ4HW2EcOHnx5SStXn8q4kh+UjooluTLY942Tp9xQ3AY1OqCd
3WoKFzUKfo03/qRx4SnS9HIXhEouXLiacnPZyK2YM74bZBjDvMTMpqL0+cmITersLu3z5S1GrRX1
Hpmv4S3GuX5IEirNzNN331R+3MZkxxD2FYL0WHsJFtryQ+8M/B/AU5mAB4O7sTecQl09dqtEIPSN
oEfegL8a23Z1CHofrK1AyOzGv9G8fyUW2p8HTwXlv1HmnDgbHJZuv+/7Mf06k7563yXxH6Bm87D8
GN1SCsfr0wvtbKATIS8YkIUN9yAEyL9MdT4abHOoWns6c8hvOlqUnYX/XK8hxzze1jdZGrxbtfWX
s6LHtNTSpbXKWHi737VSwLRgSSAE22wefaoecoOJl4nQg7OkuHuaGh2MRkiA6VVd26VLFjFZVcYO
GwzJpS4yEUpsAvHfO9Icp84kfCyrDVmEAAmxtGWdw3fjfeA7SVXNbixkA5gelxeb4GkwkjM88Tsj
Q7uy60KPD2bVxplqaPOqS7oMIXsXCqlHAttAiGsa5m8TjqV4VWPaUHxKCVgGsz9KKqVcZnxC1U/6
jwsI1Y+zz0nvjUfEtVKYb0pDy1yAEbtQXTazxyyKTRbO82t5cOAqVI2mbTtElJi4/oHpPdtm01IF
bPu3N8qOxSLIxic4Y+81bBXGSB6r3bBA+Z478RpK90uMU+N35r5YurWQOWKcH/97/xQ/spEWM1sV
/nVbcDJz8bQMhq3Wva8GSK1VdzUg+Z9OEKdu5eQB7PwFiSXiaY1Lpf+Q7e/L/rFxCDRWR8pQk/jA
HzUDHAIhilHsRssECx3rDV4zIZlSKGQDBnE8CI88E9Mj5HwRX/4RXiaWqYBDixVDN+Cb+qMFrr8+
PXZQpJVkbxtGKf1uXRxKDF5SK8YtPUQNjXGkiJtg5bhO+2V1+enLl4YabRRw3PTDIjlqfzzkbd6Z
oVExbxymySd7aH3r040mIonoGQBfIa5wYCeXRplDgF6JxQqQPTY58IXq7aBNX7+sOHDh9sRRt3aD
Noa6OsEhjNQ5slgKXJGr5DpwyLNYTzu5LZVTnW08hVdwwKtH0jlCIMv2Uw2OK+B/ijmaxEH2Nu1i
T0fAdOGqrepA+p+jDoxI6a2aFWqnruRSQZyz4anKjNLmS16Z80vCXBzaDS3F55x+dmccDgXS+3LS
cQrW/RP46a6AQdcccaP2aT2TDRDQonPUQRuP60L0MHQ8AEB9Xbl+c20pY6iYhBjM4ztPFc5BXod1
bVQvjMU1c87Bdzd0qzgjMAP4LYlRdlUBRzVwI66XcapvM+cUTghLC/9x88A2uc//rV/Ql4B1AVep
ASsBazA/kJN+edTYVHadUMzq5F/24P6aGA4c51Ez796zwdLtC6J7fS2zMmwHBBrklHissw/7nIk9
3AG8CqLwDQc0Vlec+GSx/U5EiLAvrwq97UqSVObSnQ1Dz/AZB7tC3qqW+4cAmw4djfkdgwG91Y5o
TTakSKLSAVlF0xF4VIk6i7e0O8n14xrpbksChQgeUUzp6fyDO26W+EPNOvBZ+bYGrjzwuUdV6Voe
0LIOQYCf363JvjIECOBin91pDFvaB6Ko73y4e/2gzvQDBFuXRyh2ehGYxTl3TCAWShd9FTS3ExNF
sa2aymMrDxGcgxlKpnjH4TuXsof7r0dMyRpfJEr+/Cwp6m0cDY5pOYENVCunlwwzXAZysosC6vjI
puJ1zFE4KQO0cs8zrlos1sMki4OLX5o6JliCZ66mdiRKG+r98V5h8Njz5FijdAFi8TPBy1vAKIw6
QHZFaH609gHjYp+WXnglbZaNSZSJcO+LERanaNg9I3X3OpfreId6zh+yP9b9QZR7hpiPBhcpa8zv
RW0fhijwHYabFGSLPzoQoqTprWh2VE2YtjolkRhG82PRjfU+tgeX1jKvJqt4l5+kB1s5B0Hgvcpt
AyYzFsjwb257v55+9CQkoGeaGNUdHO8v1aHRUHZC/s7+tF8dASrh4gR9eZYhj4MdcE4gi+EhC9xL
06XocmJ/xbxdeeO29R6tYhp4ms9M93E5KHwPx4fw8oGoBjmQFngbtSmcgV1GH3IsOm8uSB9ckx5I
dNhF/logYtC+FYPnk2LKPu1vYYKPjJTo78OlRoGL0ZYz182EbS0b5ofFKNMGbEwV+HGWJExRR+3X
Tw/U9RQ1zFXBJ75ehopMNdQz7n+iATY/SEwXM0+WTQp1KX6jEZg5B5PtCooY176Mfk4zgRABC+id
uTKcQ2nMIcFxFtfQQiarBZBytAtOSg45TtksPtcR77vacyS9tQO692+gPWVb6TowUuEks1fqJbQk
WKM8F1JWaqpjb0z5rJDw/6kAa+vozx3OwMrzGDkBfJ42pHnRC/9q+ixa7P7dra+90eRWJ8UF+oAC
OVYOlLNJ6TTXjLItX6K8T2yEuzeYYERUwwlJtZqa9jJAc9hBI3+XXTuNdBHs8uZdDFA6gKgYEmJQ
aT8pdtlhz/V2heympNC9ryv5w6arF0huRr7sYFpPsoYhkq95jCUMsQ5+8WZNt3Qah7mQD/jVd9Oi
D8+sTbwky+nwjZL67zbggcG9WQYeiyYj7sw4RtnWk06t73eLOGHaHwo9MLC4ms+AMmleF9VBSJYO
HITg8B21EOsaS2l8mXCUPNheCbtqLN0CJN9xyqYdjDXEkSgZwrgBmb49nKnIPUBYts7zRtn0epfu
qRjSuB3MTGdJiq4FdDW0jWp5j26FOpqvTmaRVn0x0dUtalt32LyzmhxsH+4yLSBFlJ1YDL5F3uvu
omdKnqjuIxb2FOkb77KQG28twIpL42h29wC0KU3/Ma+73Yklp+KLQR/zMwI9uYYfO7vJZ6KsEPyr
n2ntpNMaYstvMd7un2xyT3kNyAxs3stYU9x2ua3BEYA8C2O2BGhB9cniZ8AvRqqqpXehlpYhcpDC
dbzgDKXNP4f3Ksd+osu7szYy2+v8Ezhd3EDbhTLaWgIqybV9UP+1V9djcpa81o+AE8w12RBIQ8YV
+ZA/G8Qp2iyt8U1NxtGIi4e/tPG07nmsr+DM0JYyeHgfWqD+5MmuK3tf1OtP8LeWKUr8/GuPvEdT
ac4Cp8PMz/Fn/wCQ5Gv2N2OnSNzUDfqFhD62cnV/De/0J2aKjKccwKPLgvbREdUVxGX9BAjf0d1O
ohOA/NvZUe95jNfjTiJRBhn0usdbC6mPHGFefk8NTNeZlxNdHaoS2DX/187q943vIu/GebwdY1gQ
3kUNuPwnyHfjkEjbVZ59sBwC2G+fGNiuGgjkCf58GZPakiHu0P0dTF2vum/QUC5IuoFl9D5F2hDa
4ebyrKHbA6vdEyFRvcortIgiNyIfHM6OorefobZs/VHgpYMUaC7oxVZrkVzFoGXDqheFwnovLYRH
ptvFgOK3gtUmb+QIX9+ihdHyLk29ioubaznUnihhx1B1m7d8lR8wWBI7fhtAm4/jO12gBn4Drq72
49MdNuHqOUJK/EXsPvFTIYE+YZCVrX3pRFzMns6hcnq0LdbNNcNu68is6S21JO+ZVEAYF8aygR9Z
PYxOyInn0r8PGCSrKJTsAo+WgVg624uFsIz5+bOXolEbZCwh8r+LHMVijY4OaflqENdbPGgiRbCG
RlTaYXUpENtKT6xJJFpwJ5P9p19TwhjnB+7kRJtOnU1GLL4gKcgZ/pxGvo/q0iNIpSN19U1uXOp0
94yFoL3JEUiF8WXA40WDJR7p3tsxjJ6MaWvHe35psr/lk3c27Yy/+uiqYQraW0GCKUKPTyzkt/PU
v7jErlxWi+Biglq/uXpN7LAdKcWYlTSGHlaDzSkmiQK2CLjEOsBwXCTKv2Bl1hdnC3hHFtelLFLr
6/VTV0YnpUFIvo7AcJpEeiNahBUJgfwYChTgZBo87RdMCKp3FPdNoj++ACufZUk8c7i6pQnKFeUw
Ox6Nn1mZ7wqnkms9F7kEJIzShMu2JMp7uWrM1Z21UBsbJoaQojco6MMoTJxam6fh/Ck7hDbc8hUL
aMRI3hHVrcfqrOLX6sz6Z8SL+VrMPjrXJFFWFakCVVhFUThUYRwW/OgGu2OykN3I+yUYpJVSh7pH
duyMgzH77CC7JGcRuBeY/amym3WCMEwFJn3rw3YJtA/VFzJlvnWeLzczII+0UqUeQC+8GZ9f6IyY
MsVbn8yoEKfWuuD982+8xsHTKXaLbfXOw3+wd/XuSglcOmswHjS4s5hngmzRK45JwFicAZpRBHMu
NK8JlWY1rbfoO+QuCP0wa1XKoIlgpqzAk2GxRb7mTMds6ZC9XDJZyOuRGe1inLy20A0Q2JJ/r4uq
HwtwnUcJid1Sx5cHrgCi4U+9OaY2ZoGpraRRYhhwKPXS8+XLgKoTe4BaBukrR9CAKzm3nOBB3R9k
KPObx65zZzwJfoKdRkwRttphezVPEsO+zGteOj+94RRZQMufUSd9Nb1t5krLUCgXH5CYjK/p+O7w
VqdHNmx5lHjynu9pSsLisi0dySY1kN1B5nO3RY5YmUyhrHxg712a9cErfnqL+iOgqWP7ljW+aLmh
DtsVZHc+lT0Us/mmShFRqvFLw0g99kLxF5B4TilPYsIlujzcSUnxHm7fDue1KJUgIBDtYhdZh0mm
MoxQoCS/4QS4pzi1r+DG9+2ajU1iGkodqWxrqfDjr9m/9gXUZI9NSzw+nwZodUjDGUFKt5XZh90P
Fl0Oz2E53x58QjZo1H8XJFA600TV6FKPtWFNpHnachwBfV4U5zN/pLqXmFe6iXUSHnIG83dAhuyg
nBfTolHvtqg/jF1+JJ9641S06P+NNjonObjOJBlqSvDk/MRcuvO6rxaWx4oq710mdsQ0VZVXR3wW
TeZ5wztWd718jqAzMdTzN2He40RuJ8UvcVvxL+Xiqp7kJY70DjpRKOAOiJm4HCEVmjwyoxVxlSUy
Lmb5WEU6RGk6pw5MFScc1GwWhomkSqZ9dL0SwOwFxSD2RmeKmyPRSpLRTN9Uhd2gSEHRtQZ1HdAE
jaOvuyWJxJ7taPgfbEMfgRr5UoCxTy9xCbKHInWWV6Io7TrYuhb0ghWM3hsX0dzAY7QrAoBbyhLe
GA8nznNrRTf+oqxo6m5n0aOxisUo6bkmTJbcVk/s2Sfi/Ts1pwWOMxfZLFEBhfilqI4KnPKfKXfI
h7D0hpozl75hQg/Hd684VNAKP0Tf+rqrXPDPkAf/fwlN8YfWUCJwtsrYZ/3qlMDUE3rfJkapwTpp
yTotf2LNVwumy/rJKzsaClpTYp2FxlbbodUy7QsBFARXAI4uwuhCGhT5ELkzID8FNPIB6m5KBpo1
wo66KUK7Fu3eTjrd+U7gcifA8Tm4YJtah2SSglDfQ1TtxngC175coIMPaUtXcNoaVfYw2tblzLcC
oSKuIEIrmwz6cwSdbculDs+nZxaLtAeToJT+5nEs/W/DUAQuhjpfiuacMM7EZZfIj1B8fSIFYD5I
K2PrOO16DLVPpVqqa/6KQETvSo33Ff1FVDVuYhau2IA8JGJ0Y8o+miczQhbTnZEwBCJKjWOZTjND
XU4sRfeVkflqnqUcx/QskrNUZ1nKK8q0Xu5t7iOjZmDkEp35NMuClRz7QUF/ChGNrZDFIrQV5UZn
DsiUEWhjaQx31re42QxFwZ+QBKqvhzO8xqWE1bvAhdNkQ+nDRuNdXZryOp7l6ui2gnYAKdv+MAFU
avIF5kuh1KHVVGBuIAFFsqlm5SkmxCmIPmFXPma9epIStNpIsnmm4VO4Zb5tA/s2vZjQb7ygt8lD
VCGR6roOfuJro/UlWjXnZzB0022us25Ne3YPgr3jvs1Et7SVWg7O1riSwSIXovmL6YKRt066uIer
a0dBBlkR6Xy3EY541pLPwTwu/SddnQ44DN0WbEMai6S9y1BmR0vGFzBGlcc1RvWBkHSZ1b38Lpwl
mhwRMIi7EACxCbPCt7OxRvNa/uXnnH8M57QlI1YbV5f9yVk6kk9xtqu6GJI3538UjC/5w4qHhmHv
okLbMmgQLMmzpC9WUrx0JysO1fKiJCn+HdtjbVNxgX6DuqNDVNbQmR/gkDSBpvhTnoeluiUEdcp0
KR7VtpAxLV7yngqlKQ8MStwB9GkN0F+oFqkxVT6z/uKIE/IXhONTea6KQ5WU0llArnS7NLf0wQ7z
B+mbjJRh164s2NDLZ/waRNa4kxKfdQLUv5Se+HPamgHB0xR7kBezSxxXTxBYWswGEih1zvqc3yV7
UqmL14+JTDemshbxs/J9kKAeg/6bjMundt5yV/H6Xhb+ydWU01uyqu/CgWdgtCqmwuWMZ71AZQ0l
fhOP5DSll44qDsQk5cFJ2CjZ79811iWL2zNRtG+1bKE6hhV38lm7Ru/6EoWKn4TDBPICSVaxRjs9
TsBxIJlISEC9Ew8Ra1XX3zLlsAuOoL8vqT4m0nKJYFQAB7mZpX02BOGV3ImAfGrTf6RjLayTtJ3u
O19IQUiP+T02oouTWKHsFyuuC3bhIuxW0hjM3InFwxeom0oFyJ4VaqiClUJlZOzSTZ7hSUckjruR
Vcehym3hXeqvyY0CjIUgrU33p5UEDaBQDtpMBnyH5uxEB4/fcPvCnkXPTe2llkTN1zZEZToX8j9w
q4QwijG0QFaGPweir0QB8A2ioOBVomKdjfl+MJPNGrvon+GmBSpCYp8hpZWlhriiB3ISurBsWiZE
JvmAMddJaxMloSp0RfpA8A5uqPArWv/cKKNT9rARPWXN959DX6/lIhMLLJntxYxmr39uJ+yt1hjz
HfJVsXYk97yUtSai5gIIinfGP0JAGMxEGboDtd3RszrTicX/1blF9P4x6LoYUtgni5ZRC/k3mS92
QhAjztzcF3NJeqwaz1yQgjEb8wSXMMg0qK26ofi0nCjXm1wcdUE7AnW5uNmXhWIpT+CdK8Qu/+1k
iQQiUUyT+Din/IWwOIr+HNp4HgbxHyy3+mfTjHgSrFXHe9A8m6HWj8Jpf4AR1YT6RdF4jj7q9Qdk
te/I0hxHYuOgOzUEjZ/zIVOOK3WtK3/z5ZFZQxRxocuy+nsBKa4lW9X7AZ1pNV7HLtA7md7aZqBY
yTFkSYHh0T+oW7/UbBeJwIa9iLfGIwbZUKF7Nplq9fXNWlmL9um3Jf0rTATushJEgx71GPdxGObr
GA0anCTDtuaCnjYWT+KFwJzFCtJckgAiLGXx7RAXsGysMnYxAObvZMwmlL+cDHZgnKAp2Q5ZBfxR
JIU719PyzX3vaLfUZcn8jmvduQveRTLgUlffqTkj4j1lfUQuj0B4OBZmwASmDZhJBYRlvIYjasku
7qStX8LHm/qcKB2vRTJZaa1LZ5B9UjTZjccZ/QtlwxBSH9mCutCmZDORke4i8d/+oLlidtlpD7nb
x2wOtmqL6vePyBCOdSvyzQIlvv5GFdGaPyQ8N5E+fEDKiq2kNERnMwXYmEbDh0nNPFMlqw1aCszs
A8uzJnl9sZfO0VFQpEDGeeTv45M3JqlDjtVFJBDC7kmadsKuCFQb1v5ikhvDBI5rgwvB5FMCLEzx
/a2TzuSblWEwI4KPUV6xTp2PFGc0+Z+gYkWqUr5SdC8zxJcO8XIouSBm1TIYrM8n1BDjSZcUNsD3
UNa11JeS0FnFA2F2LZ7Ywewfamwkj/sScvNdf88s5LXt1qJv/wVnC6fjSBRYW6CNs3MeA3ksgf58
QmYBK/RfT0yKqqeL4TafOVzY3a/aiWMU6ti9Yztwlo+I1ZZ/g1JK0SvqLAmkUaNdmQYGjTerahzt
EoDbj/CYdQo6CCHdcnKxOuctmY0Zguneiew2XHZMD48nNTgZ5SrnUCg0ZTQE7XehX4tQVwMgNCpl
YJBhsCV7LkoRKsvjqhvQtdWRUKtr/gdAIkYVKJZRssxxfI0NH0zE+gqHFcGkXZWtQeLVtGW9lJln
D4Xr3sJsHckx5BvNSKn5yBAL1ThIUzQiQwKu19Q5fs7DoayhVKYNv5w0Kn/e4L00aaYJK8tlj+zh
ePOzDPF3g6H5oCIhXYGuUcSeNtHdtESRUH4iFbDfLPWFIyIPnssTTkTlUcgVHwVcU2f96365CPza
ExN2tzdtclXpTnewdQge3ogTsSzUdypaDNwCpF/mSNWaEsXvlGcA0Jx67H1cNFC6CGmPLjbMlWcU
YV4Vyy3Lw1XKPHfD9FvyGnVuZ/1V9+Pxe24gLLBWxSma5iA5Q37uRONHlqCjpaon4I/oj+UAuROB
BGa0FY9GoAWCBje6bJzpwzslI4p+ne9Y/JWccV64vCS0Y7YkBMP3gRUcax4OxIcGqpozQ73apNw8
ao71dS+0z4fxvMtjt2g7kwFJKumHVLeev1LmDcSZpQKhKZGXupeUM0ViSGJyglPS36CkG01+bHEN
K9L9EqxKg6jGes0oY76gaca6qC6YVQO9OSzQrzLMdXkN+MVUAzHZWHj5vKFc6QoEygvwavGFEo53
G3biAuio0u1QUKkpe/YEVl1lRC6yTtgS/UIWLOEigEfsl9Kep2HaN29LSKkms9+ch5ABnD8arAXh
2nsh55tUEuH3/uN8260Epv5Xhygu0jN0c/p5B+KxrmImfFtHV5ORzdI07s3Tce2Rjm284xegH1fx
D8OZjFZ1oye+lKHAIgxE6gD/7VdORJSL/9nyPHiToxJfmpJi8hPN3FzQN9v52CoyEoQ132gqKAMM
r1ga9Gj9kEehuoTCmK5TuyhAro3JwGD5N9lO7EcC59lJYmBU44nG35hXjYtmEzD2fsMKCOgYgmlW
RsDT+z/KMkiU026Y+Yth2KOwF/AwJhsDKXnsQsFVJ8uALtgTzu9GXR5TtdHB7KYlPws5Fb61C2e9
5zdicpp3E49+qX90LgpSBdUiyWpuR2PqpJlkE7MY4t9A7ceJYB+/2mtaGWpLBcb3+zHA+mGktngG
zeuC+Hcnj97+KaQ6u9t2shcfzKWQe5gYBLayvdFkNsozHKIWGlkZ21SOrKRxifMAlzj1lkM5AxZW
HViyMFdLMrxf1GZMhl6LPw12xk4iTGDea6OJXtOUFpb/QyG/PcdxTsSW+Oj8kUrOOhn8YmXKkB6S
du5JvaePb3FZX79xMAqZ5PhodJIZ3EvTfOqRstJGlgvcDOSnX/wULCIArRjShH7HmlufHW4pXha7
sR0htsYhxSl3KFEV5gnDHYWb2pI1DUXZ6UIj0YcjXBAZfmaOawNiVnLff/9fwcQL1/AZuaR95T0h
YMr3blylFBKpYBfM+imSUm7kDXODJlVQCfyl5D9lTVeavXGhL+bFllDdZRKxLAxKItkAwVR0FeFz
JSOtatMxEan3948uwYuwcVDHtbSNia7EyHl3JqD1m1c7UZ7I+Ko/7P7WxTUXNB6SM5evQLmBctqF
l7sIwPyiWXyrYz4JYOaabPZyYAoBTfBHeHr57z8hvRlT4/GQs39IfKlQE7YPGATtRtWbScX0dkhB
bhpfaJvvZZDf0BmQRIysXrapHClw50mweBHBVUZQNo8B4fxz+E3MP7BWhZ+3soOVf6814HQu9HWW
UQ8BjE9Q1VFRVM5tX6PgRI1aU/DTS+alqWxyyUrvn/L86dptwOjkLjwl9M3zYtZi/8K5df9jyGtg
uBJFZdm7m6xbBbmWUf9sQVZfigeSbPDoZOmPHwmUHfFdQq1KuJ+e83gvMZTpGZ8oEWzedCVTnzEn
H+UlOFzFIdhUflsMbL6ZjUajGZJYh9do1wr7y2RL45pWP9eXucAFPTJLdj972lAL2PmakBn5dNal
bKeLfQcRi3M2kSiDCgVxZrqdZFG/7v6uZ4VIU0NSiyhn/p7K43hXlzFIfOAr1siNWmrcjF/TfV0O
EZwE+KCS4JLa2wU0NCMIrpmnnFdoilE9p2AqKUOiTfGiq/VkB87V3NhaaQpczotGZgSxWPyAnuin
w/k2vp8FUk8Astm6rMp+zUd1whzIoB8pXe6bV3djYTBbevsQ1YzCoYf98ClkKjUhb2syIx1+DHxq
juA5gIKQQ2/qCj05mGNi6m9uRYbpoIO5LY+j7MjwIdd83piSOHyfXyiGONPXdahhrFnnKOXzEC7r
Da7Q6ZMSuwIKYlqEbjxIXZmn8VxtN27D6elc0+r4NoBMOWZDmCbR7gK0n44qZrjHQjHwV2dO9Jl5
1C0LIZwpBTgQZMFm9N85l+bthLKmyf8F6DoLMUcyOg+GfUwnVKfbEbd4Dw9leREW7nmsEY8gOqM5
oiunqRaDxDBZX0qnwDQK/8CsEeOoxHD2u5J9GRmknzjIXjXJ524GPS1JRp2d2kpD6mmns+UztcNJ
yXCw0Vu57WjKWElx6Vl1QRfLAasVwW9L4X/qyY0KCfIRY/9fyRvgDN4X6khmhyVcoQKE9sL+J1rY
0q0S0qUfDnf8/ch9LWhP/g+iGNWjwZDqT0op+Xsvih85X8bhJ+p1rGaiV4KlcM4IpCDJ43ygtx50
ELiVY4r5GdId+QKJeMBpAU8Lm90+NUvm7zStK4zPtjKTist7mpBNKixGtcNRsVhds/G3JokwLZYE
6fueSLT14o3xgGLGfg57rlgtwk6Ip2lqXx5sAq6w074FMgl0c7JS3tf+hYiav6Azy7ymzaddsZZr
Z65smU+PGh0B5SC0eomizE3Gz3dMpMYbCus+VJCCo81TE97Ir3QmfeXHAYtwRs+zcaUuOhuCmUfs
wMkxqOMw4JzN/VSc+yOt6ZtsXg3N0NLKY93OcB3KDlyC63YmHQebCm5J1Jr8AWuR0bMIgBxftdOq
LQgCykbI79AWc0s2cML9iYVipPV6ziEaDyC8fSkZ0I/azoFfjW70ZD/VnHkQwct0tMIPJqKqIGUw
IJdEH092UaILK66KE2ggjgltUvOMjmwNRtuiRjVCGmwFlbf0LH06OVnG8G9hes5bmYWb28IPqMLb
DS5W/4TYykWQ3GyGvlAMOtWu91DbKlqWqvliwtw+tmpWTfLyYNM1ky/0kj7gTyL5v0SuyisvcMKQ
7Qr/XhLf0hhpaZFHbVQM/tT1DP/AAF5gweq6/tfJnkfVjrJkuJhlN8OopYzuKDRDA1dtQQbyCIT7
OXYlZ/gXOe3tOj3aGGWCrv29W6Yog45tTM/YF/F3K+TKZYWrFmKleE3FFj+BsTQdEoOalksqnpRV
kHOfmceBfyzwTf28aexRz4/6AARQ4Vdf1cnz9snOR6uMNvGMywz4eERb4Nhd3uNb0dwe4LVVxrge
Wmt90CBlM5rIInARpATOF5a15y7LPqnRZQIMkGPjctw7ya+gBSfbI2ejx5D5FDU3LnlEi1P1Lhrb
afEhtetQbLz+rStfF2HZa9yqRgorh0/WKa0TIkosmTuEujcv8ow4hNCDpwRJLDW252wLaccwfvwi
ZFQ1cwt5Px9bXZGMhX/iGThu1K27PjGtugonkKpIdJo2CaLCVhVQTQfUJOPJQ9ROEMFxSquHC5L0
9gfOYzb3utLphOHA1XidnuwhGWQsXlENaozCBEgo7r89KgeSV0MtfJtYrhVs4KaHZ9+IKlZEJY4Z
LK6tehS6t8D7NweVNWmTWWX9+PSQ3bqYA0nJ1LgrNeIWcrFZ5Oji4Jq9okF0Z+VFohN7DOeGaZzs
g1kZtP6aOOgWfVj9c1cIoDEJ+B6db+1+5wGL1PlStWfJMfwtQ30qXt89YwuwIYxQ1uARThPzgEDr
1km4b+qMdBxEV+Iu5RCiXKOTB/k0T/BK2N88jGOb/OP377lrqTtde8W4tAiQgH9q5vmmuwUhrI3W
++3T7UpPSLMspupgXFqz6KdPX9y0pLm6XeJCfcHdK0IBRE1bKsfUs1z/KQGqR3j46vi4F6lEWcRk
UGS1XZQkq2I/TTmom614AOVMiSyGT9wDPoot+KtlD7yue2eguARmRTkuCPN++Sk7m0tkvb2TMcEH
XEfg/hQSLz+2s0z/odqqg7ce6qRVvBk0GPh2cDI3MxuTzkWGVb8MIKI6T3AYVENtMVJOSm09etL4
j5alsnpUoES1Aa0ygo3bplJinn4MMAkJF9IeQP20JbgyP9JfHkyK6YedSu9PeST9oChgz+vMHzRQ
l/Q+3D0lsH8D9gcGXEegyu7r4xFpJB1lvGXjRQt3z8iXemvjWuuJUjaUiG06eC0tTbNA9Ez10ssP
ZmoS+kyyisa+yYRn3gpp0xUMq0Yhw9MAqVVTzq6FKbINIzM2KURKU7/18yZFZ6V9Q3roR5/A3M2b
Ju1T5991/Xx3N+pD/+slTAKTAphWInt684+5gxb05Ti+pRdwoVecXl76oXSInvEZMZSXCMiDuqiH
y7l1nIhMcXaYgDy3ZOeZOICCkZBVonAfEXbMUvjbHNvAnTAd9V8Jyl0Z74lKhIg7GYLGsH1Q7mPI
THxz15Usn8mKyk4Zxlp1HEffXD7BMOEe3464D5FSnv4EWG8m8EyigRbIMf+mon4OOyGJOaKAEvmL
ZYgJrgY81gAfGYFA6WJyKJxETLkIYkdgYcs2sraAPmQWvwb1hJMXqSCNYUtdVCk1p1WKOodH/Lsb
zTlTsnj3mO5GJOLFBGdoAiN8H2i+a4PqZBhC2ePwPHOorp997yPBKK0kvj8H3Grsys3QOHizc5oj
aRlImhQqCsf5jzmslNGrfMBLESHYSrCRT4spWWM8v+qHi5BKNVuyCowadQYcc1u8WO+qYITXu8bz
TxaoMwVS1laxdChfLLepRcUko2RxGLo584nAfB4HJ1gz8hbbHu81iN2gauszgCixcOA6W+nE9keB
vXOy7hoGQrwLt0OBQ6yn4Z3Pi1G8plJnetZ5AORWWTwTAZAH9SX4Z/GcYxyxf5v+Vr/p9Nw/jkNQ
rtAs+gYyXLHUrqKkxpRIfUINS4oxNxVvw3j4FcrLHpi2u1rzY4e2B6AwEejtcPzk4dKunJfsmBF8
iI9baz1Djs8PAiDg0vkHwNVvkTGQyC9TznURuQUjXBAUMZJ91pmOr98P+TcVdpX7BwWIBK4a/3ph
ucyafki5XgeeVZNvCkoIgmTP4mgYif2NAokxQ396CAG03YHzV/VDXYs7Gz+G1cyl6gEtKG5nAaWL
vu3WWPyydRKfm+A58yBpceWPjYmUDr6Xo2t3IK2cYxW0SIEJVX4/tnJy/2PPoDPNFzrqg7adbmJs
UGykQ8gpTky+RaUUFQbdvJhAaf03bfqw1HBnPziF5aT4JyTrppysmMZW5rg5SMwdubcegyd/FrF5
rR++dXt7PBrCU0BVWx1Wd3CyRGSAX/SV3d9K10tk26N9M2ZkNkrzxmKJzUY14tuHYqaNXNMQaaJE
/lqb4CLdbb5jzx1SIVAR0fOCqWmddhJk9j0L6WV4UYfKBG5rRebxmQDLL90Rm0HGXtK2gBV3tmH7
lRdekW/wqoMubyBMe+fX+/wsWnRDowy99WxDcFzb/Mhqpo2VEnrVKTWHP3frpFmls/sKE6KwNBb8
L1VC3lNVmyllibecJXHdAl3bY23r6V+/q+90v1RYjNGqje6qkEzh8ebB6GKgPVPP4GXTjZ8AjFtD
DbalonIGrnPIa6Uh3/zy7uIDWNoLnGh5/BY/kbv27MkKzfRYnyqidQeplCvZrAxorjaYXvLnNzuy
2IkbjprONyKUVW+6jextdtWUzCoOrdrKNZPq8y7TTOfGEIBmnjFgwJE0dX24qxTF8413K11C88xD
EtLzWDeRQQNauByTTaPLKScrn6QyuECeJSQ4DBxMWYciA3LT19/+1sG8BGSFvEqt4XGRIybUs5I0
UvheXpddrn8f9xPKCRGz1NfZQC/zELH50bv1VqbPu8D9bC83+M0KK0SrvE+JS6DxbeEp1hZMNoJQ
vEglfLf9jfCq995E2SVzlUWBFnpJEk8TZNw=
`protect end_protected
