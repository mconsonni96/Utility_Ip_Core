`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
myyfT7v9Go4q7nQ8y+uF7/VRTsadURok4BIcFllS0F1zHL5/u4+/qYAAs09NA7fwS92esqYXyh3G
PJG386ygWtY4fqTpYI3xOVMQ8fBA3aZRVN/dkh9RF2ZxsFebsOfRPx6GKsJhhyH3h7JnHNnIwGzc
MLNNOsnEqrAMXmdJ7Q55BkSeSR8edMf4rxJ8g/ZIV6KDnxTrSNBV275iSP29IbqRYiCOKHacceTT
OPzquXDmmfx21yYs2WiYuKHNRUxhv5qNxs8IXjVJ0oayCyjicLcMd2rwcRCezrshYaVMFzMJU88j
k3a+yqwj7lFq6lraG7yBy3YNiVwIpY+vDW9FMw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="1vGf0auf1BjF/65BDoazcumZ2eLnd9mOP8OcBf0w5Go="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10048)
`protect data_block
VEUMOgxOMKXS/lFdZ4ouqgWQ1XuPCvJYMAkqcyIodmZrnTOGwzVobequvF9nwLZoXsFLzw+QOsE3
H3l3xLxhrT/5dIibF7Qvazro4x4wV7Y7VQbS7WQSkMvgp7jCH7FSoarKtTZHrMXzyk52X1pxbudh
IZ1M+hvxj0SmN7J0fWyx/wM4hASorGNO02l5929LFlAzLlxFjmWeE6KLZDQ7GXcEUtr7KUy0hejS
epo1cb+VrE5bCW9lUR7MRPPa8QRsWRCMrt2hXyxqlb0eDG+QYUWNbp6HRYu+A8lJX1/0z47nOfg0
9U7nARnaik0S3LqfqoXNBGnBpqOkdxwTEEEKn4SVPqRQxa09KoW/p1SlZuMF/H8WDbs9BntgOz5k
IrnV6m2zkWdnibuhPO8V0EBLvNk+8gWOqAGw4dDteW7jwq+xTEr7mfThVmzsnsSgmr75j+qNQObt
CfIh5CzWZLudHnYib60x/B4MymAavTmsosByMvdpvMzRg2K+1IKpvXwsOlpw1lxG2FzqGcuoM68Y
T40y7USWgOGj8iubLngMFsEl2AY7X0ENvvZYhUwHodybQxYMgTWapLGOutlJXNWFesU7PliPiimV
P9P5VrPS4DAVxwIIOtmY0caMAXjUagKV4IN2soywMr/m1HHcA7E0biGiHGDPOfaunaSIc/K7q3tJ
SHk1Tf/YVW8GKyF4tGE7yUzbCFngbpLx+cpCJtFQ3DG84BNAnao0qiBKkpcaeeIRzpyRerNJaBcI
gLlxW0VXRoahU1rkm79Dqz7acMWBoCLymFHoAhksxqvloEcjmNBVd/5OiSbE2GD9T0PlH1zbo0Yq
J1iCrWaKCUVapjRShY1K3TC2wVyAGrd7MlgJJESjQC0Wo0gSfci37agEI8+p8dsWPS4ymXcoEkUE
tgZfJJvVx2V0rDmq3ed0hCtEanS48CDKWO7KGNATrI+rYvt+pjmjXJ14J35Yn/689KfwJ4eRLQZo
4hKg0PfRgTHEo0dr9LdKmhWlhwhW2hYm69G+SfoxaIr+aFF3nt1hC/9bLp5y5DH5yuI4rohm4yNM
pzLnid89lAfQ8qKGfYMQnv9NZzctA57BxFG3j5MU7tulcEKRNSvScSW5KU7unBaNFFS2B3R6R3Uo
8gCJloEACM0bcZPL1vk2pzLeZgR2T4QOD/cTbO0PxffNdgIJnIy1Kc+fLAg91bBU3n2pQQ9FlHWG
HeyZbTlaerqix3+7oLCtf245EwJyYjof7Af3wuHVmBc6ezhzSMzPSsMsSWeIanhY5tsct5ypRl9m
/nN5HuJz1X+Q0WNIWlqLA3fvu9OquWVUvAHOGthVTy88gRdxTCXZKLd5UK8v/ilogMP6I8FpFFZX
OlIOJpyUTjSc0ChD9nJ+ICDUv6V+5fLh5VHzlpuEhOvff8i0niE8SXIksxUhZlCp5NMyVLhAcTMJ
XjpWDcKAkE1xOrluModbrssUjQeXKMZE1hRq/r/92keilH/NJjzwYP90SFr1xPXeu6lsG9vSwbpy
wCCQ9bd6lXWTOF04mETbzpOYvH2Y9xwg8CFmUWkhFykwFY1Xuk6J8F9orgYPunoGi0Ub3VvlOGRy
37QQlqBFtf5CraOrZNUGiKPAdtRX0AN0/lF/d/6ybO4GMud3iV3cz6jR/vQPVuYdOnoXTHlusS5J
u+hIoZFM+UkCSjJbk5MBViD2q762UDY457Y/OpBmjWeNwHIvuBvOrlMIYjg055qH+rutjTD9ooyh
ZDwJRk14frPVpNEVpphVXhWtk/wUAX6TCTV+/9gxFMXyMhjExp/VBTb5hazZdpgA8jgzOhtRYPgd
KpymjI5J+sTdSZjsM8aHIyYbmdlPlvp5G4RI5MAgzftxZa0PjtnDdRozxI9HkdQeH1wpjOUgGXLE
MjIJb6imNqqRCbmLIY+m5mH2t/wJPQk97CAWRFFCUNxMlX0wG3lmsduE+/3hVhud9I8cLlrGYyqQ
Q0I4Yk1PXCxjCEmCJCloXGFePvISCKzk3KO3ewAigTHtzPN/vD85cGap26hRpytGQuXrajVXap8T
g0Imm6n6ZAOK+dlSyQAp6/AWuFmE8QOCR7GKxBDHddyZHLuis2Bz42HKizqgar+IOf8LoxOAlaYQ
HGj1jx323Ythbszw3Gb0YpmyROk2YOG09xkkP0OE/7+t53s6UnF+Bbsd4KDlD4of0eceBMkwOwo4
I9/5dXOK5ljDyKl3IRPlCSfMX23jdK+kPZV3HJDmpdAfOVsUe7GN7ILitNxTZaX53hXo/waen1i4
cR3DApueb2XcNX1dATp0uYfxnNxXvS1M7kjkEpqokNKdJWUfvmvI1+lEanEpmam6hqe8F/T7ve7u
hy4Um7BhMX4A8NfQ+05+ICv+Vvq3OGYrW6bn9vRe5qjDBahtfxf0OFemLFv5KdaLebDnMaHMTSMs
LbcdZR2fza5HXsS59Q47Z1rwUZjPsmBVJoH33+p6DzckQbGe0tlvUxFoAW8sXo+aVlTCyn171kln
ETBcYCBo+xFdp4uotMVAn/hm2Z10bzw7YNz+FAnQVASOJBOdijP7n7+VpomENF/+475PAi46O1F0
ssuE/K9b99vK6P5sYYLQxpy2W/sEtEa61p3NyWhJgjBpFhSSO1JWozF+qZM8f5ft4Ka29WUckk7k
+cyjq8/t4lQJmguIM+s3LhOSIRYG4bkA1Wz+VINLPprq1kxaLtUnobTeHv7VzzlQmTMn1MgqXD+z
MzztTSehumOUL3DYaiYz77ISKcQOnVkU1tp2y+c1yD+G+/s9xz/V11TuimuzetWj91XmsxgPEQsF
VpC17s4ir5x1/RRx1w+hs3ZvggZRM9f3hOiG0fi1p/zA2i8wiJMydwwPrqKQCf8RhSr+URnJQdyN
DnHB0Tepv3P2xONKEvOvxQbsMbxbOP8F8nYG2pMIUhW6vwntKFdMU3GfZN66TzpabhRwYV8plKkD
iB/4mPOxR3OnztsQ6Py5mU1zQdb55zUltEYXx7ow36L9Nu5UVTrLh10V4S5TYZDfxyKWeM0Jx9+T
6ZAg/xkfVRmKiXfNjKP+vRgvzo/ScauWSlUtzSBhbzE6ANOImvUuHBbUtrIF1IMpGvGsznam47k6
a5HZ+5PPnB20kwIsFt01UIheh6tfW7an3E3Tyzr1mVil+l1M+oxpug9ahxOWSLyddgmdAW1eer3g
B94tKT0cm/hcDJV8aFaoB2qgmP0HSStPtQRR5htjE3Wd/L6hSvmNbttxtnCZuYfazk0otiFgvydZ
c2D1ojJkPPKmduAjF9STpitEF1Ga1PFoqIl7Dt9dLYzVExzSpLBKdzc9YkpAVqwunqEQKABIfHJb
O+1ukrQurFmYZM7LxUPYFVZollOdjJgBJPtLXW6a3+NSJZJhYQHxRDPLqmkKRErU9W+k9OFqspFj
2DiBcg2bQbYzy8PY2t8BgbZXN3DdJcGaFzdeh0nzjDSMigtvogzzdDnCtTxbfFc5LEcDM8xlyNvc
VPyOAKwZF65ba2XDNzDMe0XEMCn7sR3WNtSTes8ohmrIAeBZO0BYtxR/Ex7nPN2XR15+Iur4ZpWX
2vkZgi4gGwDSuixuT5DclQcPGa51qAQ5bnezCNzD8Az4OE615XimyXgN70B2Noy5MCVLHEsDYMBu
3mRz+Nja3nPuG7Rg1QOBDGmVTLQ8X1A4SAFaem22Z9uN+gumOsON55DZf2CtrnK4z7139lCxFRW5
KxaQEXeU8mM18DpPlB8uNuWrwNw6sJ9OfA7QV06ujYlXqDWafbR+aQUdmHAuxH6ew4JPUV+B9341
B7FtGy+09fzNKZUFZtcrSmN7O/92yM4AM4VuOgDdpaugnZKepCsVfP9ILhw1BrVqx8m0yMi9rdGj
Z+giQPnXxTbVfwPUcV4VvPrf83D/a+PvZlN2A9EKBG5sknHJiZZoukB1zu1EV8mS+YFNVme8kV/3
H+e76/dqVu5xfkxTMoqnwg8KXnSJn/9DXx5xr5C7d5/SRsIi2zdaXxa2qnSLN1D5hbHd5o1ge9gO
hOI8A+wC76+Kj6s7gRqApo6Jrc6376aJ4oqVgXO+xwYLAfTsuRgD1miaWOqmNVst5TyJyOBfwGdG
oXMzLVmmuvg0GgoF2PJK3z90v1aLdfzV/4D5iH3wddToaA1Sv9QtxFbNanvc7IB11A/6/aPcECn5
w3/pyWwGqL1+mto58n7O/3xRp2V7HyALsZ3BEy4VkaTa4I+sto0/m2WmyFBXxncJweEG4GspsWlR
yL1VQGBLwadGgjzxI2T2ZMc2Ww5XrV03JPV4CzEsGrOT+gYGDzKOHeC0nfyVTzGqynwQayAt7xMO
5P//w+2dwcMnyT5Akg362/vJfcqbSWcKNR/HPt15YhkG5mJw/kZI4aPisD3lf2ethGMnoDWA0A/p
uLBFiYtuCI380l0VOvpXKLzVDaRl8AMUlBwhA5LczS19Gn/luHlCPgnrdFpWerkVG5QUanrJuFhK
C1gorEy0qKLYBRZHhJnPqVv4t0Pnwja1zeybsu1NVQHYJU0sBHubE0TPdLdKqAnZbD7fe3x2ypxL
SpW6wxl5fsZT/N0bfVR8Ffmbe+kzhw7lH9BDo8uQb1mZiJviTXKNE3c7rekDigSmI55moZ7mXCdj
E3ndVERNNsSOg/RjsvYvqIifKai2EdE4ZAFfKfPkUnG4HlE9kazZ1SaWab2VFbR7+5lfuARLxr+/
MfNp5KcWV1dwREVAwRObtq4DllxrZJGk8hU2w6ut8b6AHrA9KV25OvfUphzZKiGIPGXaA8dkY9Qy
kajhzgcGbpSfpM84macpXLI+sK5PIIcEwiFZeNGCfnOONK4DKrDqPILC82U/URZn1nxGLfKOZs9p
LS+XbMNmhmNlEzOW5LCQVD+oyxSY6iRxIiRqDdCK9ax6btFMGrRIuddXnNZQmf8Y2nCE+Yb7RyhX
HEAAMipXUcU7FW+7dDfka5l0/0qZIApzi8geUIGBWnPG+ns7WS1XUCsgAWv59UZOdbKKR+lAhhFA
v4ttSy/ln2yWAwapC4rUQxcpT2naA/+0067qjpSEEcTeYnNOsLQJRiAYZbB83B3xjYt4/AzbURLd
idkniV0TVhiiNIHUKbVO0PWfPrePtLUibugIgVCFVvDfVNFzc+RAPLG/qfAc9olNXUACaNqSl3K0
ts4FOBIm1sZs8lOkw9IQKvsxgm6wGH/FZEszRCz+YORcL6zu6ZUgLBP77fheTKs3sd0m/sIC4iJq
6RafVwN4Z/C3e4L99+UMLm121L37fW5KVdvRTLMzCIpYfzX4KB2r83o61DAGUopRl62OaKXcOK/W
oB8M4hV/UBR/+D8mecaPbDMMzDB9upYTqGBlly+U7zBLb+1W5mKchfruX5/tu6B5RbRWiADbYQia
jLqeQj5kXdV00HDlVfzTo1kesWhVMjp01WZjtVsEiYJiux46VsSmR6zQCLgV9ZDFk/5eZ5UbIOHV
LSXZE0vRV/BHg8299coF1GN+rPlB8hVGMl1AGTZ8utyH53YEib8azwNDufl7cJ6fkYICUuNeNJu4
RRVUAKyP3yTZLWjEaDvc0W6fyao5VcpZKrSlM2uJ2ALPMP2AK1zasaoi3lZmAnBWcCphRioNdwxd
QsmPRjpa10eeE3Khbi6jkMwtecO0pBYx8UD8iU4w4uhDoNwQFJ07nbHgPrVEv7SGGhVDON57tdBa
VWEWWlZv2RZJCPHSY2wjTN4PX+hNvKiY/E6YxxzqRtNro3gtE00HLBDZYSSVzflCGXWAHCMC+4gF
f3OxJPsMkkxCL8kJKRd8zZgUVsft4sAU3Pqfne+2mvjo+BxurmduRZlX1shhzvdfAVWqxxtfIc27
4efSB1BbyPzeiqSuyWivv75zGOvNTE7HfWv0Wd/JlDf3c73AYO6b8YMHsZQnU+XnCkcigZqdZshk
E0ymjDBpYNSKG/fS8ViDThGacKpdhdXOYl64Twiy6gyeBvyW1fcGfIQLhSqrUZyutQqf4/ZBmg6x
66q1oD2bRDgjn7f1XUdjOsTnGGMlm98n/aVdJWUcjsuIapfvkqyeTpiJJ5MFUrfEy/O0eEV2B9JN
V9ZwP2Ewl1dwq8l/pgZgxZOG7LN3NKYjpC1MMHoOd/erZVNybmcBNpMkWAWldNqxfBa6Y60qa/bF
wSEwxUInUuE+Og1/76h/ngBdoE+t6ndlS/QZy6YZ5OG4MU1E7acopuajBd4Bu8u9pAqgWIxBg112
+fQsz1aFRzEm4FuLEcM9fbQK0UcM3KWvD8whHZIDDbL9OfitGjjbkOGmoQxXXqvR4hFp7db1BIuu
Sl98C505v9lYlkdY6fDqw9SvGxxfp9HEeJ+IFXcFBSFDTwo/A7s+hEc/0R++Mnv9jPYCfhi7ZFr3
q2ojCrToxsAvLJjiHq/jX6wCBtK+aEzOv61fKGGYCG82u2OMKmffkP6pX15dk/YQBQMp9O89VsOX
1Z5l4J3qi4xVCwoCpoBaeKfkSmILjh+WidGkejiXJUAvzLuozFAFYnfGkDQMTxpP2LRtPq2Ni/IU
OsDyTkrBPpmnv/TwstSkOhC64g85Bjz7OcrbSKJNfXTt/Yt7M0HpSvyHFbS9zwIUCJFT2vcLyBqA
s8tC+o+nzRHKfbpH95tqQnYNo+npSvZwRTnVocQ7PLos7cJl6V8monDGi3BMo2ltx5iGCJGFBZ/N
a4ct+rhvOmn83GmG0e3xN4CaZ+Li7F3Rr5SKrbYY5GjN8tS9wkm8QQcBrw6iBsvAsoRP99+IU00c
faSrm3+88M9JPHJqeA8/2lEM6tSv21psNgMCGJm6utCKq9PI/UTlDCwPkq8YE8DLGuOOLkE6ThdG
0DHo2U3tLMhfigdAUi2fUi46G/0TvMmXySlnjuRTXfEgXtnc4I6Cxhztr/PWseg8J1AluE0QaTz/
78iScUCvbty9PzV5Q9b+cUAe1pcXVS8TIOlESXiIbN5wTRwGLqyT7ellCQuHIUKDwkpOtJgSaYF4
vPKdoUJ0h0YYwG1hsbDMAl51rdwr2Gz+50W5RrJ9KTDw1RAbUBJ012BEPLpb1tFk8PvQXj5fqS6h
15Y4nCVNSfgz5AVPHCdv6+BQ+2M6d/VDFjcRwPBTqD3J1Hx9B4aHlSV4cX6ImUkn2sNRaz9EuE1C
MFAmmNus9BRMreG2AlTcy7b5mY58UAy7W9aRyuMem65jgzsWLg5s7eiVhc82/5lMmuSpdq/rupwN
XAQ6XvGrHCFEDNdmiMUk11MvowalaFQQqqkP5UQpaLs09FfDJNJkJ5QMtliWx9+47lCls6OSl6Dx
wWRT631odxh7hkwU6abiN8+1SHTOgD0DaKI7h+m+bDV3TOYhiPo19FOCqB5lKI0BP2xedLcwegsZ
v55SnCnaD8CpduhaX89yD6lq4How+rGxeqxd9Kat32MYtJVgWCfqV6ZWx7fWVCLhqQRLQn9MmfHR
eb2w0xfPdA+NvQEaWK/O1Z6U0RJNc20Y+ia0WeCPWPDarLLEbab22NQgaMkq6Qu1YslxHh11K4nD
mkfVQKy9irzQAJunC6cicZfPYzBArPsfIASpm1uY1u4cPMqdh6nMITlc9qpwsCGxHEHvpj9y4AV0
JMStMbG8XyP31HdlVEG+clexxbGNISL71hnfl7dJIb0wFM4hte24Sqt7xKX78AA7tnXuxwV3zBsO
ZQhR8uWp7n1MgIgmXqJhwUXKy/V+8Oh1veZ2aEvKuD/3KGAvbE4MTz8hxCQi0cFH6+EklC5RCNlD
kP8pL5EKK22aLfjpRtsCHeTaIHh9hRb7YFpMXBXWjxdQXvS1BUZR2LKpwlgiN/bj9lkMWa5SNdEr
n62g3U84lg9BGQ9XqJ1PtU+Tjke8RlVUhctYbOefKhHNXriU+0Z+KYZKkVgyz2QYGTBAenkp0Hvs
s4nBIh30SpFTL2Qca/zO4FUzfbmSLx3+4HxfC/6WRFTqj0OwqsDKeo+YlsxSFbOXrR+I/WBWHy7m
i8A8LAssUGKWkGnl2ndrNcimsstf5gwAlbMi2FQlPdqmCgoPBhdWiL+RGbCPoB+x13oB0dQvjrJI
y1FAfIvLV3XOpdTj8LEgdk8Cro2hS+lJWQi1cliQHMphEl/63SzjuUNP9wgWjtIq3VeZHBSjqZnI
usVCEuHidy4+FxtBY3mug/7PdjFsz0YkFg0mQKRqnamRx8LjZmzoueoGhipctJETB6AklpPUHlAz
st2ZqWC3sYFZ115hWSVMEuX9tIJwDWoTwfU3SajD8kkzaimRALZbLt+YGNgZDsTmuNmO7o6fFWQe
l4XmSp1nCzVjPv/+r/JEnAodIRzU6mMgZ38tzqpc+bu9cMOBLf3PAYbJ91LVcBU6v19U1CUFY+Q3
LWbz7lOiMd3HtSljluSZykMo0EwCH8WpQ+lmnDyiunfRgdhuKRJMaNjGR6ZQ3DkY0ac4bZdgmJAw
bQydfRkplh8EVV+YToCY1U93dyMbpjYuV4ADgF6sf6IZEUIhJ9EzzkedLjLf1IRNzZYf3O+RbwRl
7rplwcHo2bJP5r1fgS6aB3T4A1jBqyhojmVK8B1GvV+F9sUH6xlaY9fhJhO2u/teL9dvxZ03watN
pEbqkAfT9m7cLsfloQ6cCzLrbhGEXmHb5BVur1w7KPk9MA4C6VeX89QMumL/j0GyZIk11YdqoA3w
U+zEFAy636Ju07xKteTrnETgufiDa8KxQCx6rL/Y2loennoX8XJtyoLFQczAF+1b/C8OvdC+svUs
KdPlxM0+x/WybhaO4oaJpJwAZqvQiCNZwbEESGikeoAgaF6F7qVSeb1VAMgwX9rOJoddCntn1dpH
00FklabhX0/a894EXsLJ86XHtQG2OIVIm0Ys7VZZ+/oAfInEX15D6at1LFPv58Z2f23ORSW56/uZ
Sl76mDz4h/byHrf/aozk0Wv7X+N4zsvpKqI+1Isy64W/D62XBxQQzz8lRL88ygISV8z82BpGEw1A
zrmeu27rWll4eKwPtdYNU8hPNWzJ4jx9BiwQClJTvE0PBKGMo/yLEUJ2DYBH7K8JnMcNo/6zGheE
HvzYWB5L35fVUW9NlRwg7TG4QGobe+lyrJ1e7btR8E4HJChy5wSx0WVd1Ze8zk0Vv5+0PSRtm8Iw
1JFgkWOD9F1MaJzMdrZ6KXv/cG2ZnI1ZQrfcFQkrPwP+T/Jy7fp57q1Lcj557Ch85ExJw2tHsG3/
Aetp9dBDBj3di2Gl6X17vB4llnO8NveXaVj0fXjKd0QhepWVr7t2BwiK1yd/DoXXIXU8MBXMOd7d
Cy/YOAte1lMTpH9VjOyuMj1ppBp3qkxv0qwnR7YhxMYg8gcMNvAr8ESPsFL7jSIDZmYXonuqxRZX
G3ZxVOwNejL4qbUUVux6OMfRTYxzMS4UZen2y7DsNeN1Iui1xt9eNXJ4oQcD2Es5PW73KZp+95eA
ZI6X+S76jYGdRk1DHOo+AiqNOBh3094mPq7wOTYs6vOHSkKAschNFrAeuHHFZS58tUfiuy9ZwEyW
7X9mgBBIcEtzYA+ainmWEHEuL5zr+cuJJVS2/oZRzlMzx4QGzIxn8E2T+iCmcejrQQKB1LoQM9Rv
rWKLgEypDGKhwBprqkyN0wMNpR+ymXnm71q3WAZdNrpMSTWhHTgd6SJ7T6uZkVP4ntTc+NFFSS8w
KjheRcNdm3cBFpqEXO1eOFObJKKuSoxI5AtANBZY8l/91tjerckl6HWf4ZxcVc02bcmFe5mr7+Lc
puSIuYnJ8zDNRjIokNJAFtCTJHjJxjzKsfsGbSKHgXJWuF0k2sLCGuE0CeGb6Mfd3JYHeMSxIk3d
aLAewxfqUWU8sPm1NYVxVWijtFNMPTa1MTWjTaEHuPvfK4tlGFjRfTcR/6FOx7G/wA3rD3kKq9o9
iyuyCKYpRNrh+iQ2zkwJBZGAzUwhGnkY3Ih0Z2DSFYIVfhm8MGTMwVLVqY6vlOvMp6OWuLQFYg88
fy7/OHID2MV8wfxInfmDZBQBhm06qDBCus27fXtSF7QIEtd3J17wecsdtqQtEDCh3v8Op47FfdQK
szhhOd0P1kObfu/c4o9EFMr05Oli6W44mR6r6CKjVCKGSwJjtzID+R2lfOQvgXVlhjBA2u3gIayb
HomZc8MFBMzrWcV121Bru4gC4yj+sj9Q0yjLIXc2ATVswAfh3q9Kig2kHO5RNgqO/ToGm/xlXQD4
d2T+jLovbdlJhtYOFmqkuNSilQzXjPCEi7F4SwXohF4Ge/JwcF89X1Fug89Okfvf9JuSsXKdwEmH
UZ/rSvLPzyEaOLpyaCnTR7zRRPZeLU8iMHoTXP5TPiDTumHOeaLnXBr6z7VOEzmb+gMppa+cMCW8
ia0OODkk1picQFuDEMq4V1M4KwdDFx9zdjBv8tCRKORi2lRrQLzJPO2pfxcRcrUco0+YXjQn9kbi
gsp65n5DJzAGrisM5yU3grsm2fO5EKlY+fGmIv9Hv/wpkAl7ztdo9e9kXWDMqFvxfhMUOCeD+3bK
iCHtUQA6hQUUNkY5VVDjXSR+vLY/YTW3lp1BRVxpESRx8peWzXQLW0wjviNVri++LWOnDbKMBor0
iIpk3tAo8VlAyHw24bCENSm5eeZfwZfCy9gZQhEkSuOMJ7CiI2G7UkSc1jugZZpDi9dI8gU7O/q0
uvBavrAq18MkXDU/oFXo5+7yH9yXni0INomCLDokszbtCG59uYA2LAJvSifMOID3LdRUtpy+UNyf
1CKCmH+v+jrgOYkSm8FEzYM8lnp3QHoqX3TBqWMgzsKEQpyZz17V5URAx/2YIgNU0rNVUyYzyU3e
Gbiw0MFPqqdElohhJ+PO8dkpudndK9on9cbS2A0eIP3QtKr5jA3Atae1VYwDIhuoqztDEbGp0+QK
/BzO6ZC6TlmPhW/CX1+QAv/u7fzklWZCgtnGa2tSs2fEXErvq06F+32vLIpHJShWlmpwActqgvxu
LhLcoq0mAtznQLF9uYD548wjCa77uUsN2/y4L6Kq0z3bDaCJ9RqtpL3epfJkCc36i3x2ZpaYwA2A
oXIYyiPwjlvrfckOHszMevlFm+0GYhjs1+JeBRRq4LjFzUhyNZAlpvtrnBbsu/WoiF8HVGoDUinU
Z1AYGhA4r8nKg/m27OjUrDzxDzMVvHAX+bEV/O4b7C01AHbhf8DLf/N9Osp476581MMRmdgWJLpb
9huQBNZKOh5OVXOH5inzIansFPYA9k2o54q8cKegC+HdA8tax778NB0wQinC2kZgu5V4qFj4rknJ
3JlmCpk1AAsY5iDhiu1TMUi21y6C1UHe2/AhRViP62wLMiph10dkp1n6Mvb5m80Ey//NNR1UJ/nY
BzxvkRRpLeIM7Z+crp/E8Dd3aFr+isctVfjfNJE4O0PL1w6fZBA33+kiEDtIhGMjEM8hpJDdqbfB
OCdRkpO7TvsMvoho4S1I3F75ckKqAeaUayTtY+4umGVRdhqn7CHtp/fVSGEZSDHHY6OFEJz9pvrx
zN/S+6EyQByWx0mECx8gzl0RwqnTBB8jkU2YgvkMZhD/6N+faP8Uaqa/e1YVSi7na6KQUT21hG0c
hQcQbkPEKuwg9MLybIoTbOBFV1wGQPAfbNAixNKuA0X5jo5+ow7i+vSCgeBubnLzfjhfa/09Ea6D
i37hkH5vvFDkNBXpVqAaB1qum7mKc8TV5QSUm6DrHxylBtSOBxH9GEasYUqN8l0eZN+M4LJ9YL2R
7w0IgIP4EjUwMBOWvh6NOH1dHrf7mf2QmLzNePrZPDp41K3pLJAgG+8VjrXQzd9F8Za65YlF/L59
egWOCy0VbiVKPwQB/5ihtHqoTo5JjvIDy+BghEvxEht967rdc6Kmu5Zm6ytKKWsKGovLbeWYXiv+
k+xkW1cymhP+Hr3t3UOUpgAFM5tjML2b5HM8TFf/xpuW2DZqyRrr8I5pu9BIsqfMbV0EuwMStGym
+XhKTfuoJiTNcUX5Peu9hC5jjA3zZB6CYx4uQJutg/7HZTxW9wF4oqu5wfE8EjsWkAXpruvgtXE9
11eQ28PEB7jMeapFwq+s8kWfe5K27JWiWgRtyoG2G7g2Fb/Oh0mweV0feb/2DIMOocr8Z14jMBmo
dQexIU67Q+tLPTeXzSxjAYBZjhCuwDXt1YamEOIQUUJLJqqNET5rwPcGErTgleoiy+OSWIN/ddVM
1kSCmJq4bs4xTJG8IyfSWsC/lYUmmE7hvQ6B7DP6yKy3ia2+9abJq9gWnijIRjecVZT/d0mQwdkv
w//uvhrSHBn9/TteMmWvNUyvyQh0gNWYWBf2oXnjOlPrC2/azoNtpWy9+DJpyTcB+wpd9+LfyOUP
rBs3ytv3OeMSSY2ArHCMyX7KuHYkoTCU4yJ0yfcmcelcKXL7l8Q5v9LhHsDPxpvCxWRbn2pJat3d
1eoB9ry1LkM++1/Jl84IUMXMY1vT1yWCTIMoV1uV1vjWT5lnPklXpiLNhr7MPtmo1Nt1ySB7VN+y
S9B9JlsXTOiZkMo4JHxKuO72eF5t6EQx+rQorN0JVZt3CL6d7OFfDzwRfPdimc9lwOy1DYwhMhSA
RVsJfxRHQdwiLcQqKMgXPOuzv34ujTGNxQVTyRPV+B3FtpURHg9uTB8L5hQ5V7hiIiGYijVwj6DQ
UWE/1+XhgfuVuFp9gs8pfCOi2IiwY6xeTfIYlDtqyJi2cmw19Q0zpHKpWILcP02DwnvsfpQALz2a
U0M3VWFV9OhrdZ87sMIFf8g1AwG8Sp7dBn/E4drAnoOv1qj8ubI3+Zd1XCFerGjkka3LrTDeU1HT
VJTuA0OvYWGnOAyYtvJTsSG336T+SuglIS7tkD4gp+oDeeGRYt8GMHVx6I1WVIQMCoukxYUi9q9A
MVhUOiS5dc184UhWQk0AVazdfOqX33RqOc6Xbtq+GHm2eTbjAfuCDCfcMksz5PlPeU6wYqIAdNCN
b7z5J1wtITUo2VP6rZnGi8vuwjy1SUbncpn0+c0CAhY8GZdTiqJImise0FuNTcWySOuhr+dIg/y7
VUh3MO0IQYXs6hBnvE3HEz6eTG0EZBIsSsdADua9rttQtKiwSYzjMxin4PNPgug153qkze43y+5T
ZIutjuPPayAYt10bVVrNhhj7kAhGi78bNsJBsIcMCs/GobnwJ9fL2hvJdV9JlgBkK+nyH5jSvKqa
T93vxgSDz0TFvffau7zYi1UQ0CWuxNs7hxXCBGcitNK4rYm9ndKDcDj3Q++FQNrMSZ4bwq5Z61bS
pnm/cdO7XXcgNq9iKLzQuSSoswJDd/Aa/pkhySJR12yQAQoFV9YQF4P3dMpFuIp/tL4dh6sYCspw
IjsmGrn5U3uscT8UrRzFLLNvU0KjfZKOJb/9AieeDhbwDTOhvpFR9p5myySFUJITSeAZsC/NfE8i
dFYvHLD5FxXiNpd8GNGcBg==
`protect end_protected
