`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
SvP+SssjZngt/Mz22kM1uspCsH8CP77D8fJxBg9D03UIjiU5/6gVqtXPNS946PX3iuPS879tNUQ6
cLnoTEHcWiq8WddfiI6MPQhhTXKItCnr5MjWpu90LvrBVdfTye5e7AWXJOidR1iQQawp/+CCwr2p
1xJn9moJ7apaL0mxXFgFGR53Vq6L8m/BcyiqLlGo9TIeLBOJZc3U6VKF3z1FWPot5TwX3yQXEQ8S
7mTMAIgTzOaBIiF+Pw0yzcsaO8XCUJxXAv/Ov0sh9uqkZxTYqfV107Zgm8pYpfLpaxYDP7zqw3CP
NPRi3RMyrXeR9jB3DeBgs08dMzWM54JAKWIJ6w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="MOhOdr4DbGCGhVJUDVJOHbXl4UuUQldg8VxHUccpXFc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128096)
`protect data_block
Pi6CFhhYYkeE+KlJdi1nCeuPQdWDvTGQs9xC4efcLC/83iBcTqhXtyyoa2UVtSovCo7qgi+qMqvq
wdRzjVhLUqhOf1Yb64jp6BWAPOLKbk4eH1TnCJl16WboTN5CB6r7N7rn8ecrAOQgOHVAuLVCthSk
khQf/7MkNOvoHauPurVSu7VOEzOi+Fy5bA4sHYWv8XhEfDhZocv0Iiu9CgKcItlIYZHcwx0JEL1B
4XxHG2r/cYKW+Iq3REs9haigeSE+ORw540CX7ty+VvHdr8lT0L0jL4TcPY5bzBOFjhY2VGqIruyE
VeRi4/FoJHJY8JXhROxEh579HOSmP35b/tDRmUUTM+oCQHasbC9SfuIS9el+dXCZR164obsUeEWd
tB48VLYprbL+SpJfyhOHpKDiGgNAB7r38xb1tBPR517uU7a096ETThslv7VZAPI7PbSgN7UW6OW3
tcwqsoDZvdQYsA1+2PKljigmgfWzNgXurGYvm+dr/kCut0He+XJbEk+Kwz5pP+UdAMhiAr7jdyHQ
MsZEWCywgHkspmRs14osGJfiMhDSH3jLJXoR78itLufwS7ukO1OnBhuNh3g5GW41TXzYI9FO6WwQ
kjx8DFE04qLF855ekiSd+NYJVAnHV1lpnAq9iclxEJg+zbj6ydwuVHAp/OMsa5fJfZ9wr1sTaNS0
FrrKulwfqLGOLMCbjMzb6sWJY9rzoclDEulb+KpDVi5PVRZ9RCtBbQisJVahxMDEajYxAxHpcOo/
n+pjMt2/B+kd+DSrAquIMg2eXZJn01LiQgzunjvb3U4T0cGRQVTB0bE/D+JWq9MpTFQ8iGeJEBjl
SwBWrX7S+8IruxMiWDwRUtQKTh63mCNCOn/+luCxnopWbrrwARNa5T3++F41Vjh8kG2k0xR4460H
olboaYcHYboaHb5U+3+74DRA8LfSCRtNa69JL1AQmIYUz+IfRp8NooxiQpXm9ueUVi+VqruDGJJg
YdOgyNmIrhjsBVoLsvJiGo3Mtgggj9W178IrOYmFyyuPHfKYs6YJSdENZJE51JnOxh0EJJrlcayb
iWVeU6H7GmCqqrcS8a3yScQUF2Eof16/Vt7ApCzKcONqMw03RUvYFBF5siaF97Sndg8yZn5I6s21
wn1mnZjhzh8kjhlOenguXo4n9jzX1u7IZOJ7o91blpXqdju9wg2RVbUfcNHTWIux+lrZxfo/oKJC
Ak95S4h2Jav72usm90Ytxfpn77MjkJvni3bVNaC6c2iULQBZl9XjoFccHS0LYhuCGsHOaQ9tdatl
5Mm8lh38JRwbgKyoyycrhdmI9UFZpRAPmsT0YWF0C+Q4COpBLHe+nNNWv8+p5cdl/otW9Fq/gvPV
Nf+z65sL401CHFA0dgLyNf0DCWtAr3Vf88B4mYjsrSE3xqjsH4qx+uJjCP4mBp81nXJuDMJg0tsU
oofiVjuYAhmDn1UZUyjA3CEVNPbLfnzfWyhCwIaTm+/ridXyjQROleIkHCMzUm7A9y0KDruPgoxz
H4CSDXXW2g4scYpgOJs35WwaNFmz0D/62vtQCiSUE9wwZqr8lchWdLxQFe9nLHXb9JayHg2lWapC
vGKUhw8ovhQNsYusrSUa/XVEFP9C8dIwj2eCdaRBB4y++3ml0dT9066odxNPPFE5+19sfLYx33x3
NQrg7vAkdXCJWICk7eeRwy9/8m++1MRhO3T0fsNV3DXkpoqyqmxgWBA7RVic0qGiN9RgifFWOmCW
uz4U95kHHxM2+gmGGjGWJjLbjwsXtjon/te+WKm7b6vZ7MFyGoHN949aBLg2OLeSJADuiKlXXImA
JYptQpC44ZFwKbc7eybwhv2Zp0SKDaYpRCugrSJNipLWFVnh55ZWK+Qidqdayj73axk9FnpBEz9x
w5AA3mnrB0/4flVa35/1VGp3gmoQWMn1ONmM6hG4uyCiHcOBWb4nuhdgL5Pi7DlxXDos/8oZBauY
rMj/U1gZbeau4h+inTUkx+mr2FU5Ek0/KXhRHjD+yc9w9o+Bbh4RvMU7+VfOx4vVEDgW3rCDoWEX
XTDt/ejgYAVWm95nZRH7EVTMon9/mHgMPXzAH9cjlHpSafCVl5oaORk1eAEkf2z3M0Uftvr4JXnJ
y6QZFoxv8B/CJ7LtaBv92o+sjm59pb79te3UStlMi/tjysLVMrRzkRF6XfH6poLlv5PYoPoXGvN1
IlwW2kqBqfk28Hzt5mBS8EHPpvurHwNZKnlzJ/UZyCGZCs0zftfe8Rl7gWIzTcvLf9tvdDrDomTV
SCOhA0GA9XCUdCIqSt4E8sR5RSf2iU41L0bqHh3lbic5QdCiLEFgeWlTkeUaqm/CVVgiM43OPL7D
A1eB5BYOQZJdTQ6SYPA49OMu4NZbog5REUZzCzp5aQwnypDSJcYEakJz4QCQo6u6XH+kLMUm6wvQ
f8rWLg8aVfaFYehqCLREXDcYLngaloQTCQAW7vHVAZPxmofIqs0WBT5fjk2n2AdvEmlP6S04Hjgn
d9QWTZD9QtgFLzpKLE8ZUuqteNYIlxrxS9fsxWDJrW4laqLapuEOFtufO0bwNoJZUdlZ5IuYUw0e
wFues0ZZ1TPE/woRKOX4n355KmU6a7S4D/4aFvy8dWJoKHhI15twollKAHzoxhyvnS8fP5YSMFSN
a/Ssn4tQ18unZDAWtuFqM35SX21oyUMqQ8bLp6eRsTyVmxbnwum6DaN3QJBsRlf2hBcqzPkBpaFL
FdOxNi+um5nfKR1Awtr4OscLXjL5LVeSCWj3f8VfpX5hVOhgRbNNoFdQzvokGk0RAa66xyxf5Cdy
CzKglpcYO5djkgizjb6e5PFRPoa3sD+lzD6cwnIpwdzEZCkCU4ztA+1kLZlakDOsPzbvRLv+Echw
arzoT3w+Xoky+yNcNWAcsPept3NIqRsVO6D9AMkVe58/rtmjoNCqQDvK4SlUYfTfD3d2kVrvGzCH
s4z4saoPDr2aiVmbJSN4rlyIPqOMfMlX+D3EkHqstDSjHgvZCLYCtL2iqbynymkvJ7wJ55GC/sgJ
vinlptQDlAwVXcYdX4DAE1ZRZ1sakYED6ClNUl3QG2tZvCchR/NBnTU6Hf+Yc1IrlMOqMsxc0rnd
rGBERRSOPl9vr9OQ3sIEVC0zUBQ1OxueV9OoVAPu1EPOSqqIlvuwpaTrUCRnr+i6iqeusGvE6wDM
3VckLZftksQVzpryYwCBFlgKxa6xwASz8JvyhxWmrUdS9LBKzmMs3KclOKs93bhgnZB2pJwm6BF9
FKIX1IROgksR0At5b6Ol9C+AKboRBhOlcWgJ2MnkPg/Mo2juTEB6T9JRCe9t3/mtbD66pmpt9dsl
OKF7yDq7vdiCAY9UzTOlhFCOnSn6J/iUPQbpGVo7Gi6uN6G6Ck0JLoEkGra32nnDKFolisA5E2KD
EFGI2mroP9voZwMTBlNYcgQsv7RGXqC473LDleCDk4RgxuZUp2EMF4B9vCRl0DhQQ8EKzwGGC+fE
ST9YlAQGqUUymleUaBakTiS702CpcNrIgSXA7verWkjKMjZh60Sm2PrSuJc/bFAXRWtCq2h7fiLf
wZys5Lc17sRqzSvJXFKx9TIvrRnWsnpqgQWWhQOSLJ/jiu1fCdsZLvCdsqv/43ZVqu/25CqJ/Dqf
bp0kfgmLUWEMvWeizRyDu5SPsx9NAu6c8Oa9pNrrLDEpG6U0yMh4IVEUQpTvGKJMnPUul7DmUO1O
HhFMqm9oIrXIw0Jh0pbx4I+7NwcS3tywEIkVpvH9T2Nrs9F2evx4M31UgwxE1CVQs/eZsVOwc81U
+3fNWPo7P71y9ZBLX5DCM4YaTf8gOfCX2skDeSRK5gooOXcZvubYWdzp9dIr95vH5q7Js5zCHEBh
nnOouO1aIjo5/VCXSGpyGCUm60P1kQ2RuDqAAZY7qbEvL5VziUWl2wWyV12wqU21FXZCowuN8TXx
efmARamYU3HbIFwpMs/oeERYj7FWSgxeeCSobH6pA0NDrWH8TN97+JdUf1pUPKQ2f0OcG3p7JPj6
tHoBzMEioGePLkeRlfKgO6c3QdU/GCgE41iSpI747Z2YRU5jY1x9l9d9S2waMbG0TRIf9ABtYyMb
6Upnr/deN8AxU0SH8u6qm/nYBGezq21qGXvaVJQo3feG82CtyibkW3tbI3zlsOIoT+UxCCLosVsC
JcX8YIxbm9YpNfJCzguBHcXRqqFgaDjS7dt2dhWfJ1e5lDei4DvDPc5uTmL4MKJwo095Isl+gs+e
gaD0EqV96bKYUbtNCEZ3UDbnAhMRquwS6s158z8wpama9guN0HHeEZ25lSDc7fnHFdJ/vGGeiU1/
kSyPVqAL2jiQq777L1enNpc4/W9Avoy+rILZzDZj+fB28evyxFPiVMVoxb9oggs6hraR8smCv3Qq
JjQunZEZjYIlutb4tfLKh9BtnR+US8JQD1QcWII0eUcwQsbBhwj2e5W/EVUe+yMaYOu5AlwhELjN
YhavPKa6hb2UhvTDagnTW0aFTtf+TjYhLAzqCk4I3c/fZ22wNfdN46ZIkJgKcWTnG6MiBY/RXFbs
DTIH1DJ3DniJGB55kcLjAvxXgSq9VvG0xtAnDOhEBXBJc9ESp1BgOPUGmjZpnXMrg1NcozZiGybt
yZ8+DYpvehhrn577iDS9bw1fQ1+VujGUN8mhqHBWZ1xwlqrEDTb8gyjGIDqgz4sEEbiSITfz0fnh
xWiw7Ju80bSrZuwBaif0r75IQtSOTwiZQ9NPDKBhips4PjV17bLlQKGzZ7sq+DG4OOEDL4isjSqZ
6si642NJRrerkLEuWvGhgqG5QedNmTWMT9FkaGc94wTFJjP2OYpmdvuuiFX3gaW7oq4Vw467Aj30
1m8YwecHrGsx05tmUgpyFhkJ7e9xJGHcHTaNC6uiEDlvrMmTQInmRgoODJWs6gTJqu3YNGl7g3y1
fyeTmOpD6qXpySoGurDmnxRw3RqR7GnnELgOLd0yqxYrKb0qm7ZcBRW0WTiw1inhmKxqGmISfuEk
+E7GcG9MRPS4c+GUYUSVv24bTEqpcM5QGzz7u3IMxy6NAd2TKk2tfEXSEqfEKuw+V+lnrMUPO/1P
66h+FaZ9Xmko64xv72JY6sf0qF850NG2sBQtDtJuBHKXQOc7/cJGJTAvoahRQABxsiShraG3cRVW
qhYl+D3qqedVLIvv+SKlQAUycFppgdyORj6aJSHCbNISb5lXLIvdP+cIxV6l4SCIAGtsJsovKmNI
Bx9J1iZ+6UUUQTtsSqhikLcJF4t0hjpr8RYb1b9h7kXqWZvzYF6iVOYTgdftHe6DNO9ccrzlAb9g
WHAzqP7816iXOXkvn5vw1ZO3tAtuSdBOPl+n+bTuoufBgoE/4pV5Yw5XcxT1JpbUwwrZkDV7qCWj
ggKAo016TG4wkxrEV7Jmle1JYtiNGJdo8p237YthWVvdcfqsjsp9zcb6eWsLPOxUhqk6LJtvGu3f
KOl44A88DBju+KKm1rAxysA2Hj4CWpr7Xod56w1kdQCiqk0/UMGhT/Z6reZLDogjn/qx4ygshPL4
ScVOeLPukm7Vl3Uc+uniQN/WLO96x6LyGfBq6Ku4nGyFvTNqwegpAZm1+RQt/BANPYoMffvuz7mx
+VGn/aXLa0/sfKWkfQQ88cpAtziHdwiV5x0eaugoiSfK2uWTUVBV+qOIpODZUYUkJVjVw3aKuC87
cZdiOj4u0QI3AyWezgmwzwlKPCrqMOycbJQBycKJTiGXPxCMkI63K1uWwgasvARouXuweM0sqQk8
DvnFxnGJUHgoEmW57oq2azrBmaUKll3cXNmOiecMgUBJezvVaOryBwFaiqfdc04q7ocgzX4IKGra
g7039TxGNKz1ZnvFs7LFmp3WnG/rWeiVJparv2OP5iT1vXvvUmlX8VZCumEIQHkPsGysjFF9oK19
L3ZYz+z74929Fe73f7IwEWhHXhFLC3x1DDs4SqQE8+1UnQV+mVYLt054Xp7mmQ755W9XaAr7byH2
slZJ0x2wDss4Vzyumvk2BwZRM6OuRBBE6k9AziXwOFyLrILSXgJ6T3Nk9ujEVCxe6+xaTDd/uvJu
wJw05AexjZdfBVR9W8+p5EQgvlIu04MsROxmMEIoXNOM7H9jfZOnmPVVbriXVzkPjeJ+bnUYBZ4A
GDlxqDAJJaU7UpbkdAEKDtS6LwgMB5DgLId12R1y2gEVcL57BVxrjdKjCXgJ00O4/zuf+uZfcEmT
7MCCHgBA830tcVAlAS1S2OiUPY/tVhp2wqFq45YJmPlFdqm1ygSOyPk9iEfenGUVsJap9hcVsG1y
oIZ5T9CTiNiQJMu+qUBYRCrWG1cLlVZOpIFqtqRYeUuN0gAivyA2ywe1jDUShQh1dedDgPt1Ui/T
vj8je2ArFxZPdn/Kvjwfnzyb2K0CdxGRl59xdU+/PSUR0dc8AI29/ZcFEhTg0lOh8ZlfqfHKeWdP
qr5Ou3MMZ0ZZP8tMSCrxUe75tDWpLjhyAB4iai1sLHyojJF9nPVGGVbXWh4Uo9W6yE1PYQ/a1Lo2
GY4kNXcbJgDK/MZrioJCa7TaRmAvZBfhIXPBPm3PzFSslSU6s9dw+eGcDLBix91e53kIWn68fhsH
IGVq53e6rQxZ2HYOsLg4K/Ya2rkWKf5qK6cakq8rWRe1Gf+3qXEYHan5eVD7D8F0Rh9bphxEqVts
sp5Xl38DiZr6h4BIdqIrdjiRl+UXGa3gOYPmvBNtbdD9R+7FWiGzXeSWqz5O/RPaQDdJnwlWxF4U
V2RUkJswhEtuknX9FKkHrRYVGU4DiaQrVYjLuFhgKuBwyL9Qn+nRjkbdTyF8LTJvAvx+j1DkYPOL
SH7//iXcEjD6UreXxjCf/Jcu5duUPvq7KEg9lxgNiSZKNptCmw1s5WtHEERB1kNG8Mb7ZMsv2etB
FMvKzphR7zR5TyI+UB15qoVG6oguBi/HDzlD5MFtJP8/0/vwJ0HLAVAJJCx4t52m4mby0YSXn/QZ
Fc/qfvbLgneWy1mjzjPgiXS1WV5Lle6TXOGZ69VvKALCx2JsBn+MAu6JaLuLAa7SVj61S/zP9tBI
vC1oPGPJM5q2rfxOSo7iSmOAgN/XnNykpv4Rb3YnA6R91vg6QePrvvPJPmodGAj/FRWflXwd7k5m
resfDWS4Gf635pb4PwDwQwJPRl7ape2LLNX8HQgp4N+umT3cxjiN0GYVT8L1DAoY5YE0YzhTwoiG
dHvDUOGyayr8G7vvZAFbqgbgKkuvkjHT5vcrgnp1TTcOF6cu0GoDPxyDo8BQUr8KWHVyXX29NzeU
cQp9LbC4kaBse2ibJTfXGBcJVybtEZviWAsoGyb5DjrP1cekqVMEC5n1VnODDsFq6FwE/TzwmQ8t
FxFPeSPBKR2rfbPjNJgC91EZmS5bkw2gOj+nnWxiwGDbZqxWf5xuEwNm/n5rwv7y2kaa1CpaASli
WU0gZg1jrHFB+WfWHF7cGNxSBvHRw5xD4v9J4Gf5sBGrP8bQvVXx/foovo0tW7ulGrRlqWLexwMQ
LBG3C/PfrjtJfvFndrOoi1y96dFyyc0yXSrdC6jF8w0zGnV78NHe/HHKtm8ru5pqHbLQD9q/ae5r
7PjR7H/NGa+mhQWj1acFUzZTidQm8euS6SQYNOKwP9qSKE7E7jrnKqvZr8qZTpv+g7lpF7calyjo
s3eWqWhFDsxZNRPTfSXLudEaLLm6ufAiGU2SysMV/SDMTfhE2WjoqaVfdL5tF54WMp10Z6plVZUI
DfYqfHTsV84BdKtCZQfD58aKIBeP8ADZ2Vye3dQ3wtGtH8Synxz5XDbRAe2+XkI3Xpmm80FJMkPP
UVCaGxi1ZyKpH65nlhLlYLf7lI8k4Q2hNUHLMOIQbxebhanDpGvEl8v2XIsHCTZNlCN2fNHw7gRW
ky3PZCBzrFAm5hyHICgbYw1pc9gVgQdJMLqJFN8lszafLO3I6AB9HY9ukGRw/ZoLhasgSQBaZsSw
xG3Gb9dB5uLhYnaYxFul2RS3WvZCVQfD1lKMugPWtOHhZaDtZDzlEA3LZuEshsIul7xj0/GoCRYc
98cXlsgdk7b2Zfv4JIqhV6iu0VCZpHKIxWljQS0R03udXYtAUzVWuTFmiLUaoqXNwOc7hL+zqwO2
P82inn/U83bXylnxe08KVwUxsMjZU1YmL2ar0ilKJt3X2/My+8YgK/cW52mmZSNbGesh5uOc7bDL
PsThc71L6RcKtUpYx7ch/B7vNUGfOWGMWft0rU0TQes8MGgYlzMNmS6Xo6ZTi0e6yMuwOZ0cO+EK
un8oap9s8BT3cc/BZYW2jiHqmpDIn7lf4u6zrX5hhK/uJhjaEazfHX9VtOzq2/d4D/EFMRocS2E+
HmmanCZ+rpLTAynI0Au9Zu22OZSCdeiD0kHB6fOv+tCAMWhyvxhXRJstgi0yNQEWR6Ox9v+CJPo5
1ubl76h2IHWnhrwGYHyth53rO69xk4zXfofbOho5qYaNh+wkJT2AVzh66QPH7SNTBMfr9WHQlrxt
dYMaUAFtm/8qm59hQq3evwYEBKyxesiYuysPiTycGFdQ6ApF0anRANaK8q7oRD38kGqM1WVpqPeD
ZMlZJNsdCSJqM4P23R9RtxDYJVQ0sc+i++F4L+WM79n+Q0MlglVd34T/NwdgPpEMlBcv1nqq0/wO
FwWqVKcmMpsO/i/sZS6V+P0aRkb8IVH8jr5+hwCNvBbxzLEfto7ff/AmBgryxbWINT843fmO/zTG
qbrR48XNJXPL6+7ZRBK1Lj+2z6sTiAEO3exrWTQKCzywwcthOy351z/+AqEaOg3h6nUFf53TyjJ4
QFjFSqvda6rtA+O81JFyLyrOLwNTWyits9T9ZYFoK3a3yt6RK7XBXzJgSMsrKCDsbLrg8xThXwyG
C/hkvZVhkpqTLkpQcemGYUsF+TeGc/MoOD04EpMcAAAhB0vSnc+1fb0NxrxCkYQcfC21Q1gQwOMH
JzodF+6RYB+9j9lWPVU6/jmZ39Dm8bnRAxwuBy/OfSPtchCjgwj2PNBVWDrtRtztKzz00kkxy8xj
Im3r+CqTcV7ot8sc0kd4QImWbSmdNU+Xqa+BLKgSVycvQtQORl6/bGsGZ2dDSXplyLSS7WBqGrLP
lfKMpAp7Sh9JIziv+ZfsEsmhOHArW0V59h/nC3rVYtPzj8sGv0bj8aTfdM2ejo3PaSiAzrMAwiLX
k7XhTcGLmC5wXm+FZ8DTyc5mGeCWDav+RJk6JX+qC6qvjYzXfMCtaKmKyWPZXddJ2P6+GHiH01Rm
yyCLXSRqKHML4dYNJgZrxalYAOn77/I8U2LXPmKzTqsi2WIeuSYOF7MSigAy392g7X/pzEfhHCBp
nezT9dwSpjiPx54D5c7wuQ0/IklVHL8LYh5Pgzf4a6y3EKyLf2pyoNOdNRDHA7y4k24jZgHN5Api
38sV/tq4dZlFUeQHi8AUFnJfe1ycHLDZNlZDD7ZULEOrfMvQ91jvZRrjmwADyJOgEkXgXT/CDuBw
d71dRZ2PqHrWuEbjOiawXUkkF+easfpyy6KGEDTqy5ZMs3MVkAinPinrc9IM3VMcVEwNbfuJkufA
Ybn0EpYnKsFsM768HKQfWKAEUuBxF+f4qNiu4k8TJqEEFnnpsCqqKZSqQkHDqLa01UclgBK9Nqi5
1Y4z92FS78+wzZkZFMjyP3jWbHjIhBa5WnR1esZHWkvYbZG5450vjqfuwfGmkYbQYanBbgclNlLc
VhwBqNZZ+VEVyKr6qX9Bijfs0opO1s7EGf2FM2Z3foxDmD26C17Ac7qmzxDMJypyhQzDsS3VKr/I
0cbkzZULkbshL+LPpOD++K4ByAE7bzkUvOTl3B4yfTCXOEgFmerQGBP6jlIoLZlSGi9yRtyIUNFg
I1K70tlOtEOgpQYm//mIar37ymvwxphJugYgjWTjGKUA8NZUc9o4GRo27rpq9bJn6LlCJabct0CJ
5ud0sKM+QDI6OsG+IGUecs8qnWQfCDPijKgNGDu9Nsd/xfWqMLZLQes+7p+4gfw8mDfVog4z/TOl
PVcWKXbtrdLaudcUS3MCPyMgnNqwM9ys0vYOmJE018Ec6xmtkYbLbjQDqdRsgkC6tcj3SMf8I3Yu
1rl5KB8L7EdyZ8VvK+0oTpoast76bE6g5CgnFwZkqkrdaN8uxaCurHL9bEJJh3oCmA+TAcXYA/dC
QwTL0P5GJfFGJ//y6KTbDa7kFOfOE0mg1cvryivSd7EyPohymE2v0g2DtTT1Dx2A6pfmB81fFpl2
F3XdE7J/dgJq5QJ+Ui7cIfGvwt3NNkcgjDWw0NZIS6aqL55KLb4fb/EyTyld/r9/y6CU09yrtbrJ
MIpe+HJXlF/+kLBQqnBJgvlHc5csRC9+VYsOiWCbnypru+DmYp3kfGdkbEJ3ifO1z66+c3E+gLbr
8LFbRmzCj4C2daFw+eHY9harC+5yAYUcl2RCTkbXp8czUHdLmQmvYiXOaTLdkov28Z+vCKZF93xQ
GGwmFQxrtk2SAMIdlQE72ByBV+ZnzdUeSocsVwQTGgpPpp15UF6jUGqV0KsPIxQsJ7yJItGQqsR5
bsWPNsy+1eS94Rc0wJeWu9pX3NmzJ52B3DKI9QpbehygBaxNeju1eAN+Z+uHdwa+8O1oVIbgf50W
1h7WUHtF8H92ClM0h9TGPRMSa6EwHj6zBfqtZXkeFZoYXhz0zwJtKjKOErLkQrKOxFy7XD9EHG2n
vAEVlNqizj3lFUYEAR5SySbE3sJy3sEvij0nEl7uxJ+xFUlWOWMkxvBUuJZXB80/XYk7k0dD6OmS
/B7fFPG2PQxsr/ONg4BvbTxewaUVSFxdblszyzbUgXtilC/4PE1ChpBn5TMxjURjBaqqgG4LRyUV
5mIVuuzM/P3+tebtvPCwqY1ViDkEpBZGwcVAWc3G4QYBUXTrb+SFqvuE3n0OpEfZ2l/Gi4XdTZdw
2215Hrl2BqleuBmoWfhZBDWg89Plqt41v6Xyf7BOMF6AzQlukJH5Zes5qrSjxBZ3k/K9fiaE0XCq
EfDR30Z3xfZZyW5h2Ya/TGZ+dmzBrMK5DnEMUNn8LgvY1PcX5cIZruHDSYX+1VzFAdM6+st+inIC
50fsU+aN7YE/oud9cWYX91E5/JqI1pi8wQQrwYRqVK+j3N2DB/c6GAaPHEjQoInJ5QKL9UtR/5yt
Z2iCXdUiNl8GNsUDzBPq8KoFuB0muyQXpqj12iL27FMYhmQGY6xTOkpIODEq0NhAE0ysWVqMrZsu
P+Szr6eMjtJACL6GyU/0+GG4+DjJCsCG0QkE6t4z5kyxrh4TKeT9jBetuE+Ai6ulh5GLDivUXYlB
TMy4LXkdw1pdH16mOq2Zf/H87vmaubbQhCUomv1b0m1yBy1TSXfD/SiGpVTYYsSAIEqyCOLAJCUs
Af/29+DMZrMnxHiN7rdjVzWfBiavF4Y15kVUP3Kneq5dSTEMaSM99c0WRM8Re/uo07iB2+Xc3IUC
UD6VREhaLMf221NKK09mEcKuWeqaaGcMhz0JmQOJhqmC6/p4baU8ywHFCindqmHd2VCnY14UnhJc
Pve9UtWRz2Zpv4A+Xk13V2CBQlr3hmUH674loA2zxYLHfBApCgCtTF/hXmJh+SCKOdCSB2diUm0t
JUHE6Y7qiHlOZt4GT7N9XNGfJWwAG0Rj2v5SEyCQeot3MHVdKdP/R9Gr4mpi7rjFJR2JqRDGg2mY
5L1K3P7Ej+CJrLllUj/1OQYOysCQi8ARFGdeB2Lcd+RcEl93EKT7Cd6NRgp8A7RKCSCZP8To88Q2
r1XA5HyTVRSsF2h4BHfFh9wphA5cpQqyfPOx4o18mU7rAEU4wdGCPW/kyoCGq+LaN6nl39mQCzPy
eJljaRd3DKQ4erOJuQzKVs9DFMfHPXYSUJF9wUL41uSczmOLE1t39zBRfcgzedmQuwrN/nTXpv0x
frHoR4v4au0xe2jIznmFx6Z5/AJQkv8bfRRQNITbddg1x/exIvD/IVBzXqVVToNCejFXYa/bNlKs
X3QQ+Cb6t1RQDt+Ez/Ck7zJ9bxz922cTWWpHFZ8z5upwJOzrmtqj1b4W+oZf6ZQvgmuPb/Ss626G
JUNbp/jQP0DgM2oNs7DNvkn0ZMRWt72bGsv2by6eGXt/k2l/cawNMDXQXEoPsw7T6yk8dyakyvaW
iG6XxC2H/YufO/Y3EBVZJX3Zcckn341wInPosjGIQOH3ZrplNsoB6d7dFsQxQ66BiUavPbtNuLCh
i+mgzgj0fJZ3PRmys+6QsQvJG/3rPX4qogSBeQkJbgm2+JiMeEdu+9ptYeS64QsBIJXurI++fUPn
jS9NSRJag/Tx5FbJpLMG8cFTgaibyuCDHultSs742dqs65gcFX6j3XIlhI5WW4LrLSRnnKiiJc6G
BysO/ATYBBVhC8yZmQ4RshoSVb9lBwNWtlajkogmpRjw/gsSKK8nDctEafHfJSCBAgyB6UoflpIC
3po6NBQE4UyNAdy+Wa83/P0UP4fToHP0QBIFCD6f0REmiLAUwowuJbpyH01Wr9uqcBfNygZJQCP4
tGSn0u6tLy1zmBLr3ZISkp8FteSG+hB5ilAIdhDGLsib0G7lM//HWiSuZUYZiIviyH/xD7Tus/md
9fEIkQoQ1Wf4rSb/HEtI41qHF2WbSzcmlqNNEAGhsNhQVelXF/fJMSLkuhx92VnpVXHVEn6z6BB7
kDfbTFFErl2XOxhiPrI5SCag4azzJF4rA/mhYl5GjtbGQKoCNCfQX6SBWymFRm1satTqJUG/mUlL
rd9mcCGsa53rGktRKpoIDIfYTR2XPclUqJ1CneBZ/Nh3vdVzH8uc63wg4344tVT1C6poKOjJWRJl
oyrGJN4lKTN2RLjeBQbXpnDje4pE6yhRZ80Vs4hEd+pjNiKNRezxbDXJp9DSz3EiNE47gSbEqamR
9eUqUCxrHPDF6PkNU5B2Z76+OnABLHblB5j6p3gCsu1lNBe1wVSWnYHwFn31bKhsY/o4wyBZ6gYA
B9tfrOk1eKA7f0kItefHm61/lPXzhs1wDX+mjdlQgTFMRz5QNRSaptsrXVtXn216LdHSGh3SMQv+
0Dj/ZBGSjcx2pTduE30Oo96qPc1X0f/HFKY1R+pe2jq+2uwZZTojxhZX1Men9IyucNzUr1EqyFWY
ZfvMGMwGBjlO2h0L9RGLcRlMhDLEAtyPvY79JvGZsN2GX7gH7PJtzpWkKunG3Z2+bj5RaV2dUxBu
mRrkjNOTf8zX55S1woomTkkpmtU14hQruQCSokXxupl5Z00MHtjWPFEjkVjkU7Mrow4fdnaXoV47
a+dvuGz7RQFKmB4eaZunViBAd09zXZX3CIbyAbIngkRXi7rhKAG6+GyhVNB8wQI+/j8N3QiYOBrf
26Rym0RnWkN4lKa1I3SkBSDOxENoQKtvWMgtKjabIb1r9LVDU4lZLX7wokaTLFJ9l4He6BLq4Q3j
Y/w1u/O8tgLelvAz5rpr+0ZvgH6+Uvz6OpZWMVGu5ddWRbYi84sCLcvoJHwvAv2UsHKKnf3Uq4z/
DKOqr95Al/2GPirFvmQtU4cdE/KroiaLRZRm2PZGDHzXaQfDGyrjMpeGF/5yKLrqqsxsA2+soUzA
MvYZBOYgkJA0xrlHO4oMzmEYs/vmaSNuHMERL/VBNaHlYx2ALuJcVbyfYgK0l9q2jzhMd0VFZCAD
NjaUF105rM0RtGwynt+e4rGkgjAFRV5yrMr7KIWiXwUoNHq9QdBLiOrOHnDDfz0uy2bRjyTKp98T
AJSSikpl7VO7KK44vbeOOdSyjIYUHUA2yNRNUiTGKmEN1ciAYOoZyipsudia4UpYhLpsYn/WSEW5
fJY39CmVsFf16fwkuGBPIXXlN1zvRJhPMdmnlCMjfRswmDIjMSzcaKh2fZKORFJDwOu3yNKgtMPv
4cXys+IRhyyK0IMYEMB6OA9FR04mMSeh7DTmwOrQlONcA/aQsMOsrvQGesKbazBZ7fiJwqPdGmWn
EJ7jEpVjaB6lYg59Dg5xIlqn7paIiLzuQ/9avZr3i4XdN8BQSWnULEmSWo6VXIlhrvXQZgOtl1dd
+6u/niAR5qgXymoP1WK6Sbs5GyyOj8XyQVXT8DolU2Fzg5nwu6eHTmhQfA3fnYq/+UVwoFLb1iyb
kqN8I/XvvSNfS0Lpm6OJq1+jLI8j79KzT00CSbGqh0+5vfF0Pqc/vJFyTjaGoSspyQj73DGrgmcG
LPgJoFdap801c+BwEGwZpTzj/9j3LiEkJurEWjpKJ9jY0H6SiHfVQqwFHF+bvrwJ2aQlqJcvIePC
k8LcgrJ99fxz/6JNBJov2F6oYlmnHac9P/4G4GAVt/PSCkGLbjF+tP9KOKbPENsXTvB2no9D8OfR
yP7evIDTUIv/VkbXH4fBdnsGg6OM3hWUCfGLlbRcmUeEpqNgrWzPQIGMejSz0XyFiQAvsAp4fyYr
m+lI7L0XRSDZzbxv6AR+VLRNtDnSlsJhMpUcQRSf1ILtzarbYmWaQ7O8JzEd1erMuRk8n8NNHoJc
6sdvsNRrH4pntX3ElCcr2ENJVcI/5ZVZdS7NzpodpYIZ+kTdE0TlE6gMj7uaMLatzusiDI88J82O
TJ/DBzI/JJ/CJPYatO9AEOB78jdIn3v3wP+BTYIcVsywDTvhqhKcmCiulmGwrKdSBP7lJ69tE/Uq
ecwU/EYP/9aXuK3yJBLLLMWMjmnLjE2cirx0ZWZDqE7vajq54gv5hoXD9Kr85427zG0rLGwelYHf
1lwvTzW4aZvYQCwJUc4WCST9WAYeTFzO7/mYocD/7EJs/vrPSiASDz4UxgMRdS54SHTr5rL22WfN
M9WgW5Qi0XYyDYHAAhHcMdM2icchRnB+4JTx0jC0SCjloqnViJzYBXYticQSDQUpz+Y2IUNwqBpD
lGCWJDM/Sjjp52cRzh8vB+C3waEIaeQrwL/tZHxS3VeDlfmJ5yJrgNyw8+CiTW0uwsAIxbzZh8g9
lvaHzlS4n9X5Q4tYATpoqRbojcaEco8neIZkUCdYJHpJR96BvId1bsQ/RQCqEN+qepsRn1EK/jMO
fd+TmQaLvcO7lpQdVvw/3Uq6BU5yR+Ocb9dXxNOFJEE5snI7TRKdSBCZe5ZT/DHrhzXOV8x0DGm8
ROMSsLkqvqFPG44rxdiE571r4p7JUEhOSYnHM9y3LL98OYBPJB9KRMh1odwKo7NhdjQ1B5dykRLZ
q7YCDPgTjx+7aqLms/IuP7OaG743BbfKzcx8LdNfJ9MSwyQljiT9tsf0ad/DMqSUIosmhRe1+sgA
2O88/UaeJD9gj8cFTNSSsTIMYIBxczNXazoTuNh51rq2C8qRDQ6xR72vd7/OEMBihVA+UEwTJctV
giedbnvvzQt3OB+/d2wksFFB9br+UB1IcwjW8ImIOONL1hv8ktcRwK3+dZZigGUY4sjOK2j/NKnG
EuYkttfkUIvW1IUKzOX1nfM5uaP28QFuHXg6oQAkKDJdQ5BZUELlOY8lBpZ7Yrhal58y4MqsOShu
Iv5I4DFsE2+FEncvDPcRPv5fygzqfCqSszTZX66LcZrjauss031ew8QyjFyPDC4/zXaf58Jdr//g
tkq5jHhuVUjDcRuxJRKOhX6iQQGDwZY2RJer5BnzG2LcjB5nZ9l1YQQsfHOnvxbCpqWGD9yoSDXu
3vU5v7LFANDj4aDeZy+9V99iJ4uYfcu5Z1tndfM58bsxEc9vPusUVOyc1MVhbBnRdBMB3Tt1obsu
NCL5Tvj7Ib03lfxlABleXxKZ2OpvW9P8TBPH9RhmLFN/DdeZiRUiqGc58G26ynSj/EOCwmN3XFJK
1L/UATv/h+SEPvhJGh08N+55kszfGns9HtoFD6UGKHP96HkeKrmZGbvZv+7XId6yGnf2z9MNR1GY
EabPbN6yRGrze13InXBt4pvBfuYHiWNLAQ0LnDK63Oi9XvPpLPWdzJgsGU6ZsqpNhsmopBEvVgpA
DE85/3MWle14KmOGZ3P7cFbAUHQ8rR9sqm19oxDDecS5oVSBTVhsVo++edrlhnrh0UFI7WNLSJEm
c9yBo3vQ//9+4XzWxYIT9t3fAfX1YL3QjBNxXKZrqdnSOi0N+BJVXi34ZHtngyD3ycQn6Dwwzeqh
LBt384Vv+CuLtjV+ogVaElaDtwRcA44szNWbEDw38EjAqhxVup1k3g2Guv909BlKdPI6/GDXHs42
KfcN9TGVB77cA4UwUmgRYrZKQO0dK1YRk8DB0kNMU05CrygASwGj72PKDWnnaghu/R60ol+iB9ul
8UjEYgQi0NPIM1REVTnav1Wp/lrrmFtZpu8GrHT+/qWB8ow6CacB6OkhwPWsgGU0RJ5IctPzIY4C
4vqymRI/lUPOQXON1MmM6i9fDBFA27mDIOskF5b6bxkjsGs+uG6BqQScOLBHLJlx6Jmx5uftU79v
N1nqSxHlGFA/9pHCVAsh2GZBGH0Z+XOQnnS8w0t2pCO+1TAN8CRQYWeyn99PJjKo8x/9Mms8vHcN
2eS/WdOS+zMQPVaqxnKLwYiIRh2ewQfAh862z7ezBhm9rvYlEI99JQNyre04JC5F97sVvyxDDvgo
6X2YXbUAuYFVz9P0hL7bvlBszsYiE9KpUdYri9wtKBuaeDzZsyoK3BMYGdpUmVX0+z8VDY/8ZB76
akYveQxqJ+P1aD8bxdxxdvsrYMHJcaSUFeqitIKZiSM3TZis5EPiZPd3uuKPJ7XG7GUYlNyGOGS9
DKxIYlko5QQYbyDNhaIjUQXkBr5lr5ZZP6aov1L7ABtxtzeK8UfHzfiSQrLpEjpunSESZw7uckhm
q4+d+hVlcGvrzC5Fgjv5ymJB+S1CWs0jp2Hwiqs02oTk4fdcySh6hV89iXxdbuLnMa9uP7Kmvdej
y2uLgtBJu9Ti/RO3t7aDR3y8teTBCbgntiGkGB7sYrya/wA3wD4NZ2TXDHg9nWUF6pa2axi0/Gg1
u9VR1u/Iir5xWdUKEqjL11IyUeo5ap/36jwHGQWpwo5SLXqqV86NSyZMkCrB4KwOoFzeTcCq+CW/
1gBut6dMi/hyln6vAX8waccg90vgOcaJ7sQvgKfAxT+/lyB2b13k9q52iFFKammSl/0GWOdcUV0A
SKWeFh7uU89Uxqh5ih3gxVmlN39ftLVmYJiHTvUiRLfr7ZOpCbCuXsOfpA47MIvWUzJr2MolD5Rx
lmxWYIv9c2f9ZGv8/TQngzkXoERI+fulvGQY3k8x3rB+hOnPg01a0MXb7ZkeWwYU6C/sYeA0k7Vi
mBnK76UgHXBE8AhoUC4Mccxwa6nI2KO13booJZQfbJwe5ncEKNBpntjLNfL/4aO6jWiqK1PxLHvm
wBW0kq0tMlu8oPulBmcj8RzMUylEFIXIGP6It/lwfkuG6dr2g+TPR2Sw/AUBJQo7jVbyaRaTICyi
UEqRhwao5QbuK55MnfDDidywJPufKdvTj7QFtTm32/TGcfOH/pQK00ih7/ScnJhuOvNXMve2Y9sl
1rnIeEbNTaYzxUY3/+l4FE16Uk8VgUtBRXDNAUdKJlzCAPGI7VCa7t8BH3QMuGeo09agKpwZ5Ea2
1JD+A9RCWXWVLVK5LcDPBFcxNqGIw40LDbmfAQMQ2qHlloqF4PjIbfaqsDWGDqN67aieh8haTSTC
MqtTPfNwCGnpLiGhhMLVZXu7ZxHKxFEuFI1XX7dJ62Ug08Bs7yn92E7Ng8QBCKvZrbWL+dnTGpZV
AY/xTyv0BnzB2R34XbVPpp9uqJ6omWtvCRhSrIg39zVI8ZZ2kglll6Se6PQrtPe/TUxUqAuzoTer
yAc6pQeLkdAXrj6yvhUH9Ekg2QU4OiOPkPfZrShWhlwLo1LbufNPlBVkxMRCPqiLpadGeuL87OVz
54PijkccrgcB2joLluHhjtcd9fCSO8h/ZKQr5NlQvHsIh3mGzLbByT2uJgSA7QB66yy6Gw7PFdJ9
qeBT3rXJD4Wyh9KJjJzgJdgEmA1+OwntjjUaw0R/ZbSIfH+pvlxYUa/SVh9xhXXo4+GBMbXzr3VQ
zwmdjqN6nja5iA35W0pcYyFW5poU7GrvX9XTgnyMSTg+jSF8TewRhxMRr01Y5RnTt+LHlOyb2qM7
GsRRanSsyoJ0Qopw50KjxSnPx47en4I+vufHpqflZSWQMaOGY/p83Ybiiqhgcdn/ZuKMdBWbp6Jq
cJujdp4+DkXyRhKGyDrkKwF/eZEfOriYNrq/TUEjogwLfh8gY8kP3JTSL35TCBnXhyQfKI7ep0/f
2aGavwJJS7ro4c/HZvkIguRexjkR9Y8yOxgfS2ENgrLH+tuGT3UC2Pjb7K1PoVDydeDXIsgLhObY
zX0Ok2HYaYDhtWAZOcE4zwF51YFI6ToiICGRu9JiwERi1Bq74iqFgWhQND7iDyAxTx/iTwabJX34
koLPTiZ3P9nKfXjUovjl2+scsTR++keXl1HP9YhMtZRA1DTUYBDoumguTGslv4RWDhoWzkkQM0Xx
fmYMdrbR8wnBNAqZ5f8bvShFW+W5QC3eTJDwoL7jj0/M485x5Dgm3ajidWz5jGv/cTIwMK4nxei/
aUo6rOEcf8b4ik8bM0kE5ZpBsPgRCRwVhDqcP/CuWcwrwsoOL0mYEU2Q/wSWGBZF0mXbZV2687Kj
ezhgbaGX+REb7BVi/K+u2xIAKeC2FOWZ/pPs5SDhVOIfVPUxQwGFlnAtf4DNAB67KAgku9SbXUMR
Jsll6AiZDrmmSX+4qU0Bny5WC4eeD975JyKu1Gk9aEIRKQW7Ergnphm7EtlIXAvicczFjzY8KUjO
q0r+4m+cCiSy/5HYhKhQaoeREVEWBGLXJKwqraXUDnQiOYjnRhmi9CCahmwMeaIDiB5wBs1ib8Tw
iPHZ6jyn3g+jvUComQaPY+pvB0Np0rjc1OJCRmf7Bxb4aXdSfcBMB+GBWT2SKhz+kC9ppoNFlKbG
YGxCvRT2k2nzZCqZmWHf3fQGNS961tEL/8C+s8II/VqFKGPrd2gemfDFwzUskT8zu6WIJTWzX1AL
oKgqlPXdUtJosscXnX1eiK3QRPf3Er1LmxUaHowpI31Ymc9HmZzocUT0r9UKn3bEzDl7Z5tOoPsJ
OD/+kWjjMAB1Y0q/PwBeW3uSot2E2umCgAaTTwNZjxi1Hd2guJy1A9ct1grOVHkqX2oCP5dREs7z
eA5vhTRfk7m6H4x/DKWL9hnXfHngLgFH3aDy1tFI92O290764z0Ba/jhujeCNoY80PqQ4jWuqH3N
Ri0ZBTuTZTWQeX4cHFbsAkv6XQJ39O3kw8yFCnefz/g5zOHrWqaxYNJxbYU4UmeQpROdwuDXoP04
bXgnFcEUcLw7J2UOsLN7ePaQCVVIAyf9OSBSHu9qL5RPVhgAOZmjONAPJ+pGMfC5Hvf5ueGoBZJR
q9/PfikaGayfakBxPasE/aQele+N+XsfHenpEMJTmicc28Kaqc79qzLKqMNlCr+g9PFyyOKhjaWI
D8tiO3MMfuIHOc45PqhaUi9a1oivoIUheE6OBUHvRmlTZk+XkAwpCVV+L2SxxT8Obza4Lt689lTz
/5E1kMUuKW2LKLLhrmJwds+/ofshByUlaSDjybPr+AIUHX9TTyw2HJ2E4KAMuSks9PKcXS+WSR/G
o1cxhbSSMhZ5tZ9gLdVf7WVmcvFLh6+Ms/i6sFi8jMx9u+baZsQ0xDgK1WHoN1RMTvaOApsn8Ocd
jjVk+7/aiZbgLY7MnQCyK8b/Da+etRHdMzNxq2B7AZMFSrhk60j2nXBxMP3IZ22uRlwKBXFOKK1G
+hXTfRJpHW97aRRxz/WY0xQDTeU8BZePKIi/J24mrC9SMG/ueldIUM6FJ+rV72rn1YH2WJmMgeco
OxEBVlSGdxmiSVD2Js4xaCLHxm5aGeq8+eu9oK2/D4TBt7uzTSGqGNcSH8ZvyNK/ZYwK6IO5d1xv
2ssXa+yW0fSkd0758rXMEJ05Hs73e4bMeERiRahyI1mwAfsG4yqlM0vNa36MLfzcTY3EtYsXAqda
inDs3dQ1YyG41QqPtcvTtytX/K8k6y8Qy116XxxvpmGJT8oY6bFii/Hicm8HtuFt87tSm28xCd9X
xK2cTjPs3/4izmy5srX0e1/muCtFmLxAb5IhaTIJK70qjC1Ae698TN95ZJObfkSNigldWlIgHcuG
lL3IulWGIf62/d+R/KBcNr1XmEjKYF7nbBTo3giGjGRri0H7eHoWmbkbEbWnb1h115AUXtwDiiRf
97G2lDZM8nEnRIO1BIXq3YA7s3W5IVnUicSP1v7YHLwcARRI35LRt1+MSQtzWpn+SDv2dXqwA4iT
epb8WS8i+z7rPqDDrg1N5IIHpjlLviVp6jsOGwER9uUlXyJCyEI+JbxrQ0UIxVPAcaGY94i6FlTq
7PcdMMhNub+Qbi9oAd3cO67XajHC4IvurmrO/ckf5d3GFhcX8FJ6FSAMjjxrXceoh7pO0KvdYnKJ
cubT1FM41VtUyjciUVyHKXnkXxxzGvDeQDzpPIqXWRE3LV6KP6jJqutZQDEGIfVqDXqhwthY+kVs
fR2Rzetyet3tTOvvhH4MqadeA0VuknYV/aPGqlrQPO46TN/uIC4nQsbU0eSULr3i51OQwdk3MU0f
SQXipDgCxioYGiYNDS+sIfRCxCLpzGkaUHe/h/k/LUbR5bxHvysxusAqI6aVK6s0IMqeXujE9zQ9
KK/5F28HOQ5UQBnwKpcEo8D5WfHeIdE7Ya9SKJgKle58swP982TOuLh37h2SbVR2wkwo1NU3FAjm
pCw/ouPDY1TjVNtnD6j3ComBMdjKV4/f1oK22mMWfsBmMLSpgLTE+ZsRxVcYW3zCdkRw6TP88vS3
eEXszqoStgwJ/mmgWBRldpnlkDl1ZfJcRgU8SMKoe9Ucd/17uXOhJ7P14JuHbsHtw7fArpHDC2dy
2fY9UdvI7f9YYVuf9T9WCc+1O6c63XDa5ZEkIlhXR2GUz9f/qMy4PCzkGOy69d1b6MqxOtTD2I0D
yNNbHKi9rKvuYEO8VZyAEOx6IOmxfm2RfC3a8BEDJuMViRBHevWI3mzv9RkyhZ0MORHSnGOq/Gxd
lrUNlBUHtmWyzWtrVF/pjQJx96EfG2zO8eBfPQxoAswXW5lDmvjv5JUfdulF5c+O/2+a4h9pOEcS
Iq5Siqgt1UxSkCqUOyFpOCzBDBWippCfZ9+weiE+8rGtbYtgG8CtWhxN5Yx3kLPii9uqHV19RhOu
X6zSczCZDGvS1QzY+sVdNetr1KQJgWwEjzStY4BKBV53LJ4g1fUYZ0RVdEdGHopxN2oUrUH8Z9Qx
AkYV9tfe922Iadp/11kWpIfFtVE/8dCeqplWR8w54olICOqcfrRVozWRsQiY0YXsBcANyPfcS0Ej
BC6OJrTT7BpFCXUNAoQhfAZbgd61Vjs8+XcFPHuXS//vK1eGe5tQnNjJ7CRKeuZpbCA3pPWlTmzv
a2Qrj41eaxDNE7Ls8/p+RgkxC4bCfsap9SvcrtL5+YnbiOuOV3TjQwErQSsgdBTEkVOaa9YCUP9l
2B6S1ecta0A/P2U6f5UefKy+bJ/DgGBqTAcKzvUb16t1YNJuS+Ig0vUo88zwauuS1Dt5b3QDlpJ/
AeKFqN+LLsClw0Z8Lvh4YNpzzBNTDTgiCW815YqWipzhHFuOQIxHB4LE7OsjCw5xTRrBzllY4KrZ
eiBqyrNkBQhYjlMdUKZ85pV9XOV+dcuuB8U4j5BqYuRc45IYRVLt5EFDcTPnOZJWIPrbFEKFQOPb
/bkU/ACYi7M//E8VHPNqL4wVKD1owU2KHfvAih1f5WR0Fnn5X2bYLGTZmvv6pOeJcQSk79HuDMbK
Ujj4pEKCHB8lQlmFP5xSkchQoyz00alLTl4QaNU4t+0a+XvwEv3iTeCmSg3mda7UH1aadenj8GAT
IQNjlQ5kJcOkmUGmg79Emh/uic6JWyKZ5MuQriG4QOuUsTwLYOsWQD+3jYS5adix4+gE6TME5SIs
aP+KYGWEhH9QTK2RoHj+wxKUU+r1nmDo/LO3ydGrRDM0NrRkdrYuad51JQwU80yyWZXryjMM6C5b
voCkZMPKd5WyXaI//lboQOkKDXW5C/lK4Cbc7hq7QYCpanVDzgZJETecI6BMC/O+uofPR7WQy0+f
E0c0cw+R+Ehf/fabdKym8agQqX29A0qW/0sk9QhW7uoxcBou7K62fGTGWxU2scXhV8OoBKf6TAnt
CKU39NlxaKPpTyG5YIPpnABe5iD2s9RXuYa5Ik8tU/qkN3MV575btnGFrTb5tOQFUHmgFT45Xt5M
81aDAeNGDuowRapjeA9Quab6OzKxzmJDf9jVYBro7m2fGoliCj8I2Oe7mAYzv4ODtAnOyOdMr1cx
yTaoUD7R/BxEuff9yxG0bRIXEzqYOeoJUQ9ovVV2jEl6112CZK/Oc9DU+kdRGeTYxkX8iEhhfqrZ
Jv5Oeuv31uHlhSLwrI1NzsiDRt/St98u+1tTFeDrgTuroOfBcwyzF44LcZzsGG7U0B9xwJ6kwHg6
0KifISyAhptyePMgWNoi2dqZZ3uHcZH+F2Uyjf9zP+Q4S4BLGwcmL1MZukV/FV7TSdnuFjB2mK2i
jzCfgKIaOs7YcdfvqzuSSvgkxqXMys0ejG2DKuNAUb/oHtLZ9aVmGh19ArlifiHMbqRNIa/mCenJ
8CT/g/j7TidVzHojayw23TGckTWovtEWECYnSlcF+ZLTPGRg42nKo4YCAYhzJveISNVpRNAieIpF
aAN2c0pkk4aRNe3AqtbGYJoDj/E48S68kPo5z3iHJqkZNqaZ5i+f+oouLbL0+lbdFkfxVb6t7GDj
y1E9+B334U8fY7D0qz4vffnFkTqmyMIMnBPdYE3igdUYtVZvu32yXEteKKTdmnVS2tFJjjC9oYUd
70tWsFz2Lz5wU4BRxOEKQgv2KBj+2f+QECqFwBiYINVC0z5HrNPRHm8pd+L/JVy6VKBAB76Y9ETS
GAK3PLuoX3sVVSNCJKmGrVRi1/4nAuCPIEmaz+svwuzutuM+XT9Yir/2km8L4v6yadLeZIkTuGdQ
9L0LYOoMrwrPcDsIZwYkCebXoIu0RFbgGqmsgb4uXlx2edpdRNpB9/00I0dBZXXKIeBAUuLkP1de
DM8tEJ3pKB6ZTL95PhFoFzTy0CYoYPZpIzbc1f265P0o6v2eccYsEm1iBahflDVZ3kN2FBlcjT1j
IDnHGIyV5vOMGk7TRHxxrVmJg8PYsDZXvGaRDsi3DHooL9HXpNUftTg4DhdybWTp01RGHuprcosP
R+CGgbM27FY+ETJrjhA5+nnSty3FrYCjfkxEbkr5743TyPMABsRAT3xSleZ3NOs70H2j3Gpim1cz
rC5gMhiScjTZOV81n3QV2vqsZblyB2G/FVibEq0abALzhwYwOaSlQAh6PFrs82NNBV7fRP/Fo5bb
FawBTFQhGCBWA+oWHeX7pUSlmXHV6wFr+EHgWov0tBwaRxnLy4Aw+MmcnlvVusijVqYyKCsOKbc0
OyreuzkTlCDqsqkyixtm41MG9SZxem/fukGvIQZ48bUA1CtUQoRAgGRyFL34lBPdUzlcivhVLr0x
DzJfbYQxGF+ee9eesEOHib5MkYkYiibfuK6GYyx0+DJstnmTjSD68kwBiEWlcD/EvU0xFR9Slr+i
AFvZzk7ebV5mM/ndpRlepG7fAj69uBoE2GyrPRU8/FLNOv9b1NGkBDuO3pgso1ITRb6uwnPIl2vi
VznhJV/In7qSZcjXKJQQatGTdM+U0LG8cOJXe6DnzMa3/52Pk/c5jC9BEChd5gO3umdUBS+QrglL
EJvZd1w9Ms3cKQ1QpupmaZJ9iQ6eRfpqgYdbytySUzYfGIr3IiB+/wQRr1toIgNpANssx/aNJD3s
6JOlXdB8HH9ORiiPazlnT+2BKK8mFx7V/+NYxPXtZLZP3ETWOgf1GwYE9wf7nsq+8SYyUVpMOLcv
rgtIjWQ67dkEZYR1A6Yan7DNt9An5ctlgBDn9zEIWanaggVMG4rtb3fQfAg8R8p4+ud/rx+ZMcBD
2Q4cU79IbRjkpOwEbzyFKHqpxJw2QG6XQ6JPibcZQNtsn9rI5yDVKYgUK93dGFtqqW4g83XIQQtX
7Oe16Inz31SVLBhmdzzZ1s+enHKeogT4ECSuQYH/5R5LoWquJbazdlVv36WeYhow7npJSMKeXg1D
EVfmIfFqiXu+FDIBqkbK4gwwRbJhEExjzrwBbqaoXeqTHvTyMs0GRrAgRO3PPKwyhATm8vncr36U
ZNASzhr7EKJV6Ixpx6liHu8fFFuY6OOd00fiq9rYiYJqzsrfYr5E3TngS5VVI86Un1CdvmiFhRyb
9gRzyGh5BWbM+6Pwon58dfZTGk8WxYrdyWaVKsGLvnatFxF8TGzs7gPmxnOlFpIBFbgV5SPKDS3P
qE/1znzJLd43nLg+uB9+/rtgT/H/el3UtxKb9RbXZW80OnU1CcaMsjWyrUP3ybB6NEtzTCWPnEwT
ba2g4lkFwG5xcF0eJrc+44F3kDT8PDPJDIBwD1vrizpPqmi1Ol8zqzH/RkviqBGFRXBvXPEQEkKq
KqP5WCG7HP7EyhHwmXH7iU6obG/BPwUpx5fhI111wpd0v9EfB6xI/X++3z82eRNV6KZv589VyxXF
+OA7u8TThwo/Lkz5DoFQ64pjGfcBZWTJXtrIEbZPID3d7iHWGMsPT+mue+TrXpyteLsleHR+CsO1
JOLAnUzP70CzMffUSmwFbChx4nrjllQ76tSpRMZ7kAWqx0qHEi9wPtRENiz7syfZs4xdcrIBRcPK
3u6d4m+FmLjuayechQnYxdtvrbIA4MNnw+Y81x0da6EtBF3J0UlQz09PTwz3HU5J3jNJ1RAqcIht
vm+zZHz5wJ6Hr4LSi/XFLbRqKkX+lYX/g87YJAe2dC0EXVDVGQC+6iAij/hMlmaqYNvtLBDqwcDp
d/FxNu+cs16r5s7lzABC3Aw+pmyuB7VIjVJrgCxBSMtOroI0ul9HZpQzMlyCghctKf53mWUQTZag
JRHXKbiSFzBhwksUw1F9LJF3yS0TH6iYX3YLfX/+MLlzKzs6Bg2lsXcmw2L02m4cQHw1IKceyolW
MLzPl95hgYFuHmgIsQQtwWkxQIVDfjUd87GyIyzEU6/V09RhdsoLu68CvWZvv8OIsKwqJAbnhexT
ZZJb+iqWF8YuQUHD/8ZKaWexX/PPsmqDuHgOOxP1hpyuKjs8DTy+xeF4lOFX2TAc6gP6cDzpW/Y2
kOmDrss3tv9FwVj7iHf/tF0yJl2rWJ196acQGa72VYoGtq537dxrvjduy0ytGAtnU3Ff8JKyCYUi
7+3aCCx+H4ytBaV4ZI8BLnPLLfABKn/PUv8PUb9BSKjEeB3s3oq7bGgYCKXA4Jo+G9YXkhyiEXTY
s3K9lu2AERhmNkW2lAwD3pOj3OPDJGUKrBB4LQoSvYVEX1i0B4NqBA8qr3iJc2wEMkZJDiSOfR89
LUFmdby6+BK60+BuPudzongAjGSkUv4orn8gmRatApLJe4VPrEpqiWDXxMouXAN/xqaWi9Cjv58G
WEbUoVMZhAESKzy9l6k19+jMCO2RDhgEty5m3ZwTvBsDzLDsr5MXQ7MnMsfI7boHkZSGDXoZo4/M
pPTjuV+pc9g8OWeMO4GpKGJA5t53aBep8GnzKWn48OCJlBkbaonB+rKWrHlitKw8Vfy7Pud/5h6b
cvPBE0Q60eLRQrbDC5E2LPT6iUXz9vcmghg16FoWVFHy+yzTqCqaS0OUZmero7zr3QtgcS3lV4sz
WzmG53V9bAWvcmcq3qrQNHEFc45MluaH5F6fRo7j/tLT/FF5+6VEA9CtBrhSOJ/vzBQkjS2ijVyk
Rnmy6zf35da3P+ig6AhuTIctbK+PiIM7BeiT1oSpz0r1yTxcwLjx3NCAzgdwLxHucmPM+DfNrudO
OC6yXF3YkXj/uhEK8lPrv/l697+y1KnDB8n3o2QfZ1N55OojeVDVXr0pCOIkiiiQk6zyJWZN+nub
iy66kIq7pSzznvL6ShLAESYLoeShQL4V9FXGSh/QE3w+GdlMuIravl0no1CLd0OV/vsHcWJ+maZr
6+BUzHbovZfz5nUe14At4X0QAK1gkDQpdbweEIPql6FzNVlJfkiaBpF+uENlKh4OcnJGEA9MFIlr
WlJ9NjJWSAbQ2b734PJoyDkHrQdUJVoyptvACCv/YaZO7bwfNPze1/LJtWsV7dbf85G10ZueT+wI
zTUt4Em53QzJaQzp0zLKbJ4yrJ214NK6Yct4iQ0/TL6L/OuX0wudp0vUIM8QPIomEvvUBVfkAJmN
+FYb9upYqRCm1OvE0PO8CUfAZ93aj7oPJ4rwr7lG7f12ijkfR273TrjPVLiI+IMwe6Cp6FxE8EKh
p3KB9UqlHQ01Q9PvO0fmW7yR3AXnGGQ2AldIqHBR/IpXkUalvQPwC43gkj7qV5wBMF7vWHM74F8v
0in7mxONu9GUTP6o25+XlG22eLwRsvCtsD6rZmo0B8Xb50xQtbSqWgQmOUrBP5bRcyLqeZg+SQUq
hlXvT/P1fAl1O1fCD/YzbJsnWeCKwn2zGV4qEwGik+YzeQ6TuCWTJOxZ+/WuPmO62oLdpK62KEhx
bQftRIWYzwh7q+2Vde8Vn9U0E9jyCL5BDbt0R+1JWj1IksLvxqtXgZMkMRsdhfycMyB34WAvT9B/
XUwJ068o6rp2pOct+i7/Wvga8ukDQJVmK1Atc4GcP2563UkPUFtAlFJzBCG3gogMtuvO04UVO7DJ
JM9pNLx/qy8fBhfRgCV5n/XC+GWxJSPmx5YC9LhzmMxXn/Kf+IVWlfLdj+kFv20nLRNvVcatoK/0
E8uPyjgr/CUgO4/Kg3rYBGDlXcjLJwji9WAmkY6nz49t5X5nnf8BrbV8Zgx8YSU6utEHZOI6uTQX
izyWKDjEXNPnJ236ciGWdvObkWgYAmnV918pELzySL3WqYGGGG5g0fnp8HzcG8TrMt0CsC2E6GVp
f2o1eeRW8WhpDF/baiDe3hzxGJf7zNFv4Cg6dSAjXAJD5LyZ9u9w/SPT0SwCz3BM3jbRk9BCa/tl
y4RNTA3kxoJEUxvTM2wUYqL2Zzv7pj+kgM9AImreUZRmt9QjuPIj+SESwlX6bSqe0M0Q1zbozcOi
P5mzpGWb47ISqbGtmGrBPytAmqdIs3N0Pm424FEH+jSpvi+NSH9WVsr8geG6Nkm2fBsaqpOyCAT2
m+GCRy24leZXScACUIcgdRSMuTqwgPiLjcxqZBp0bbAnDVgubptJ8iWikTBtIenxzgr5zc23CAEg
0E6dcGch6xx65r923dd8cksz8lecYJgg0xHsE6ZDu41OqIO1wc/DLWu+VpHU1SNeMxi7sHmDPNXe
VZL9oIdjCJog1VCdsKINMalDuxLYoQd0dHPBz8pYBaQrsRZQRX6kdqFf4VzWybf2ryBJWLOYX/VW
rTAg2Fd+/+NTTl/tUeiKaYYj49373vooeUohl4fwSCEwczcJ6GtCgz1EBes2I/p46fqCcvSLO0/D
TYaPgro+OnOJyPGmCK94aYHB8ndjgVztiizlK0Mgsi1JqykeBeX/m7yQjLRmVFQuSLrEVG26C24a
37XN31Ne4Clomt1McsD/jBhks8o5MqsXigaEYHJqF/jq8JgYotwXMNo6xl/DQ+LeN//bc92yJqJ6
UGUhpGpQNwdRU/Eep/Zj7zCPyu/kNbUPCHf1qC4WQCBTj8EW6v+WGSUmXM5QqcdW3YiC0FI2ViB6
4UER5QEGKkBUEfKcGihB2hSNr+w+Fr5uHddu5JOsbdyGbOiD2w/xh8/OZETn5n+Kwc4VqlcMzW4/
q7jkwpBEl3+und3mshbKRBOBfTyb4J4vZZBr/gAc0vh06OsdGEhGtE0U/xlS9Ox5k9mATAX5i9NL
tKG1LvMmyvJHCcIALLOv5OrFRbMOiccTCg9NgFK+4S+WCf/i3m7VqsRCERHjtZmYYB1kJ6Gk7pNU
1BoxO1IHbp16bqGgv0Vpzh5KYOtkz4jgeQy4x1Sx/sGl8fAxh0kS974YKvjVIlxDGHAor/Y3mU9V
c2l+Y5xTIvx+CwYBd3MyCBo7O8lzCxg+xDLm5T2p22MNpq2FdO6vhzSRer7piywkp/18bpZbV1Es
MWgvifolMyOloeO1aNBQicQ+pGzJMF3faDA8DZHbHdFEOho7lR3RJuVnbeSvmR4Atkpsc0NDMx4h
XlUrnA1dA6IJ1E/WkSbZOsDPGyTMxWEOkTTccOvJvAAX6qEWBPeMVc8BgpyFqnjzLh5RrqaMdsZ9
nkexKYv/fPSBE7HdM+hEAB6yHh3/tyXi9FPq1VCJqNyI0Qiv08PyDO0JK+qo2NvdeRCyeiC93BcA
rRI+Ydnh6KngZwJycnaVQCaHIZne/d2ZM4RSjB4+djZrbV9gojClZ3x7nUaxdGyBxd3tu+RiufFg
qKEnDQOqWUFNe9rI/2ffTTSgmsIQPnz2yhzLTfC0mzH4qfnoWdMFT+eLf9X2O4k3s5WQlr39ZToo
YxsvyZTnZNwDnl5fsvMwoNF0+BsYNKPEwynJw+KlpwUhaXTJX1gzg8vV51ArVKHaHYf5PTIsEBoT
K65ka8duB6LhfyLigTVjs4YrJIwqXHyKpZVFgXfPoezQFHWgQDEjN0gQc482JSl+atVMQRx03TTX
lygb+6JMBJIskkHz7LAshqf4rGZTw3wRWWKDoAz3TzEXIluMOWKpA9DZT6u9GwLqfccnHd0LVRCX
WpnsKdpZHcV6JBZwmhxx2Dub4PPHZUujRsJb/HEEeyA3cqkRpo5sL6sab88V3N/uq+4CNnOgcdgQ
1t634BX/4+BHkC/2KYe3ZccyvtBHvR6PGigf+jEhIt5O4jIhqvOyBHex1DAEeW5soE5kvN53mZWN
88/uTXZZrosCBQPgvUBR58IVsXVunco4wudEaCbM5jpgWApY+8kPO4rpeEa68DKv9PksgsiFluMZ
CBAFpkFrHVE652Bznnij+AfIDFEp913Ui+vUcfgkBpPoDedsKUVHXgcLbvn7B6NzZk1jzwiC87x8
tx0+1zR4tf0drM1nBFnDfuF3TfrMecnehT71uv6y0iJ01JFi+RxOkS94BK6uuxpLxFydNkBv4zZj
0PXf0bilSHQt8PlHjceJZNUHh1KJajyIP9kcVk59Stj+G/7YTH2OdZi3q3AtzV2QbMWfFsowSzuB
Jw0OTBKKb9jRfCHKbaZZN0tPCIUFlAQLG35EhJWP/FBKLCfZ2OaZ17VQiqBQOYKZXBcT7Ef25fGe
7GqfspsGSfUS0QnZqtHCzwhIPcbRdNS0OFMRQEzx+StfpjxUkc16JV84xztYCm/QYpwLPcH0QUj1
xx9HhBnbOqe6DOi/PwVYJMHYajL/lbVtwGTgEDLAfsgn7U9nNhGpavBc7/npegxuRNj+XbhQWy6P
GTwLSwZ9lcwF6ZjzQL1ELd7PwXne2H4dmVPbwR0zHvbjFhPjcCm6gxqWRVAZa5lKsq9zGHx9eb6w
pnAPFijJeUErY8KWZwExv2SsdS/H/1AvSAZKkNkNQXHY49G9XqvtOGmekYX+9xc+RJfD2ebmp2lx
ngO5iGsaGcd9yOMT06IOmijZtDzzd7Cqy5W/nEpPEg36K26ohE4XdPa5yNQv1bPgRAAvIMvkkXf5
qDtYH/sYZoIwj6I8bmlgpaefi04nhpwQWNud+8m+CswOHCA8H3/se4ixe77xNaimzZuJ3Y+RZV44
t+H2RdB/BZ0C4VERrttSQ97KP9pUxrDGWmQ3dCMiPoDZFSxbSvo0NyNcovp0atwFZ5VomMAZLbPy
qoeuHS0iLQAHg47Fl8cNgcsPHXmqE8SXFIgqXN4ljrATZd7XCqfZ3usSSIbFnGd5aMwuNbWW7SXE
dx0u0pwzJMJnPNn3vFefl5greeU5QaVFQVVyKnc3jE6/afrZ6ZQFiS7GZX/NFJqbh+z88pr/BfaO
wdO2x8BhC78/muQOT6pNfM+z6jOoyHF8AS/c/7g1Nx/FsTqzjJOzwpY5KqUT07DVpjaVqWqVzUrD
ESdFZXSN0CYo3Bcw0ZxR6nHbB91azx3zOkjQ99hOmGbW+oSF8EDz6U9qSkl4LHdA+2a1ZVeBBu3t
13i+sz2lmJIir7PrjN2QKTRE2dOhVVklcQOwL2r7fTtOgZP792N1uv90WAx7xAs8j7c3ADmWiwp1
o+yRgx4ydi9hW/Btqs7QYf+cIRwx0jprqvvhv6xxoIT8ApueoLEs3Gw+HqqN9kJhF9ogyP30iA4e
4okSFUTbYbzNrc3JKvQ7LUL8oZXdPF5GxpMZqxwkYmDcItS7um0JGQ7DC1pi7OnuuF4aTtYJo2JL
R4Jh+yG1LWm7GT1OwSJ6yrDGaOeom/KZMuAwouMceL1JnxHh4zLFfXyLDng0nvA9gOX95/6e6WfN
fTTyxM3fPlI6RlC3eNlqlreWFRbnM0dPVd51sjwsjyOh4ah8KqLWcuUKaGvouaILuRQi7u5Vae9f
N06LDeCQ5n8gHbq0f4VFsbQg+wMWsI1KONSsDqWgzm4Chvi59xlWhf28qbjLbA4GrUFQHTxbGOjS
WrzUBjc5RkwvpRvwdBRsv5L/+F2kKQ7HKKWSva5+MCTsVKaRUvZZw2T0SCq7Xy/dVr7bcNjpA1Qw
LL741RUm1KNv2aq9FasbzhiV/BZSG86Q1+c5YEFd4RTKriOfB7pwNz4QIXcoYw5k1hzbFzw+ihdM
bon1ZmLj20GoAMrbQp3ido+N5M7pQM9bIIIRs5wYrm3HeiHQwW42YLhdMoR2FRqtdZy2TOOPGyjl
3MAlSj/q3NacvYxTPFbdPU2eoVEWC8GK2gDxX7ByiyYNBlHdta1pMJOXqZlX9DrO1440hc3lBOow
szoXMSHEo18bkVXzMA5wS2ClD9zrRGwtLcEDZcM+5Q4WVUv0woIaDR/SJgXWMKg5nSCknQUF8m0x
daxIkCCCQ131aaVooMyRYC1Ee+aB51Fj9E1+uULJdzxnGtJKPaL/ufqB8bHGAbEBxpluF6GhzYzo
qlh8rgDk7RGNMsUKUhFsuZSuZyWcklJwSG9GX3t/ppnKKPb4g4b989pMNEwJytwwNl5r36jKoey8
Ka8x5Eou7G4+1tnSjcSQP38WqdO++HM6wYBVHKC7azeuN7Y6Fejv+2Qqh1KpfRB0KslXQXBUmrEC
RG3t/2fl+phXTxw0Y+z9/10+ZLKs/nP9/gu6jPr2NdGDK+WkERPcEYqcLWzqVFFOHGw/kUcRXtQJ
Xg75hxMalTPUBN9ykxhaJ8UiVHhub7jd2mt7xBmvxQXw+bm8ZLo40F/Udmh4AEPog+DhunqzPk91
BEA3DKsyCaWLj59roFcaTBU0cTIYaEEjppocenHxf+nmYc6je8b4KGeHqhecvpt3gh4SYP0Z1ygG
WUZk9xFhOV4e07rG6ViMAFFFfqLrCnio9QltDA48Vii2doGafUU8BksQQrxLFIyh+daS2pnsC01o
MbBNe6RokeWjv6E5jhVrBUTRoiYhYz4dve64+PZ+PvKzVqczjap0vGl0pDoXT5KXTCjLb0bBq1JC
fHINI7xfuN5KHv1bUhIlpmpH9INF2je7931ItBevVhaaRueylu4VWchdHgvirmZgOfOV6PQ6KGg0
+Xhiikc1g8+hN6D5d1No5wQVagAPTaWgTD9hmk3c8haBrDJc/ciksYwaGuqy1HUO9R8Dv4pr+G79
oDXxzTS6/PzKCrHq/4LVolyamdMyWZEdmD2MeVNjxBDirjNvpNfraD6IFAdgse1QJ5oIn8uF26iz
jyNdQ3BQGdAEmHOzK774dJCDzc06LcXcLAWH2oH9wrbB7k5WbUodwpEXbsAwrq21v05z/P/OaTFb
xw+P6vjRa1o2NIaP+ENhCLUvdExArjAvSEg3lS2zq3aerhjucQjRLiatUcPwoScWErVxOyPjVtAo
mxtnVU7mmwhpSRM26ORuM96E9QDYXmjMfnWtUBT4sdJa7j766Ab+A4AH3ULmCkmHHV4+rNrtZ7hI
8NcVtRvoyK8tsuxg2pUT2hiGjXtPaTZT1LBRdpe05wo1Qoq8CP91bqxaN+QOC3eHNzJIz6HLPolX
OigtPKz0VvKuJ87g9d9O06hhGLSva6aY5rr6gBv9777J1PQBhqj0e95T2j+52ZNZ1utE7KlSzopz
fm+9QmejgfYRdp07LSmm5rUijbQbI5OSln7QuRadQmy5YpUwtgOYvyt6pA+GS5zfZ3snlE47Ciw2
BDF15yCaB5Jlf1Co7N6/ZtxOCMI+FSPr2e6Q03dqcw/vDv0Pfd07F6UATDevFyg5hXJS9oJPfx1Z
wzzjsS5uKwvre52DW+b3pIaR4XxFcxGWhWAfZjLqDYi0CWdZtKUjAfhNRq9/ZX89k0d86MoN+v72
A3ar6Z1WvggDIRIGlgdHN+szIJk1pLAnkGOmcs6wN/xe1k9JsgcUKO1MrXvGJxCUo1ufNxUlZz6f
bLQctwM4xhlhXdOnMd3XhRSYciK9Mj4oFK77tC43Vd78fKaFinEsRR6Bfrqw972aWEeEcXQ2N1jG
9Aksl4SkLTrQe8X93tZ1yRqgnNV+m6mSmnFE3LKqlqaqhiH1Q41MXv7OLN8Vq6XmSzrqr5u404K3
ZEspFsnuzCcdFSyQfRsQsn2uRGf8l32ULXu5SLHwrwpJ2ygDCVLEdXI12UpfW9SIpCRjAvdt/y4O
5XRw/zqKY50VNoZqwyNjBaiNJb8URuNhKzKUzeZi4lzVx99uSyH+334yzdSFo81kH/LrxYS930rN
CL67Qm0ts72Q6MNwH6h6Xer9YzYu2llLFHX87iKD4K61zWTz35b3/ZKQg0bSQYYXiM2f9hq77QgJ
ZZ9THG8S6PESojuSp8ogyI4SpgkaIXI0TXu1tbTtfaGZT7NcLacER+Ko4K8yI9gLg8P966m418dv
brx1jKY+mc4aXkFHUGOvatIOQv2tlf66GUqRJpsiWT6mT8JEl4PphHORGC9hgkyH87m4pBX31RQX
WgpCo1FAkIhJO3H8T33v2QqP5anTuy++UgICW/pL8EiIa236uU8I57D7NCcr1aDLC+pBR1fJXP45
Xk5LXqnjFgBLrTH4/Y5EoUj0v1D2yCWm3D1V2zJzEJXrwzwe8Fs+wGdWK7svrOCF3oc8MxIYYN9g
rxYYGv7dgPtZsk61hWNTRbFRYxASD9B12FvDgMSRrVpYB/09ZdGzkzmdi8UiHDkgkWJkkmmamaV8
lmzrCQIlBMYfmd/zdwz2w9FgYPP93FjwtTouzsgJDFPRekQH0IiFE/Vzo7Mt2QJeP5eYfatyu51c
WlInyLD7uMRLJm2GkIW4q0/E3Rkq45qULhgIwvZs3S3QugQE/jxY6BZLkJSj82LHPUKcFIURJn9q
T3S76MTeeEsX+ZQAVNxShW3wtxpcyD/4mxDyWMH4m+4m4fdLrFRVPEvRkp8RnM3ggEwgZGqLiuMn
L3OXM8Pi/BWzcS/Ljjy80t21Y6wbM0WztcB5osCYZNZP/1nxvdyHT2O9o5oFYq4INn7IUaKp6u05
wQs7kQGndDfO4CgPPmK6k6zivKKLDzy+m+EzjRRh0n/ljU4oIoJRVQvYAz1CZKTAd8LMfrfuo6hg
vX5TC6gKl9vKCgGs1rKD1F6WvaM3bcPOk3LOQeRIOfmkHm4CRfVuLbEEPcG40izuCvu0Vn11vw5g
7e55jeLh0Yty2pWJzWczI/Lf85LV/H6tGuVGV0o9UgiMwJf7OQ++jiLB112M//2EPDzXSMk5Q1Uk
CRYxVn2VbvOgBYhh/ZNclkk8NG6JzBsZ6fU3xK+xYgU3NPAxwmNzoAjMUbXe+MzlV4rq4LpKzy3V
3OJo/Q248x6acMQFzW8l0bvu3cTfRV6RQ57tsV8SFaALMGBBIRoPruxvXWsFVN8+1nOmuJYrSorj
BzM6haImSZrsoymsrCSanxM5DfKM5Z6PlQ7oV9SsrLCoC8r8krB0+U3tdfw6IsQ8WMTY4xR6ec/L
OiEb78cdHcerSfjdKRMP7P6cqymqsWZf0BxFspnHb0h1kGQ7aabT1VfGWQEDFiUzdt0ULz+tYPZT
dHcxQX0TpNW6VLmxTjIfSM4lhUiEJMU4F/VTqSDODQS6ayuLEXROWDy51BQBQaNg0C7bmUpQYW97
G/0BrBUbaGBEnLI/Y/yJKQ+N0iHoa9alUa1vkNAC6EIx3doWKaVo6TJ892jpUaz/Xglp/OWm3mXG
9+61Dqb8ehB1mwBfFPcMaraskFUHD+rveOyOpnywYxSpTaaE1djVJmEE8xguOMULm+Es1Mkch44Z
G1QMff3nABLd+XCYkM03O9FGarrpsKnCoGVbWsi4gjGckksGcOclCe1AAfz08GhyUGfKVAb56TdA
otSuC9FtbodFp6v4bg+npbYXVYUbKkCX7LRHfKO6vEp7qBi2r7xtJTD44ejR83fEiOvBaPeZ5RIb
S8cAndIgm3WK6m+Ippp6MbYLSAZOGbn1qXZzUXrswEB1snT37qWEgy/mwar91Xq9/NX8WeSqMyjW
dCrEv0Kb+xUJvzuAjSi8NmjLQFBDjnQOq+zrnGw673qyBnjQ48653VUrFvdjlVyD5lh3KA9HfLDW
fPc2vK6UFBDkiNOCHdPTbj/rF0B2IhenWStASdzu0imfJDdv4byFSbFKWvxM8KXRrKwXlywYrLqf
v04WlGC4ISE/9UTZ4MWjlmVOmjJEDUdJ2c+5Z4PeSuArDtoiTH/cFsuhTB69Yg731GKNEo7L1zgK
NuRiaT1/NDWUEFINq30zTbfVl1l4edAzOmFg0s+bp6KO1wlF6eTvUYLTOYP4sSCmaafpqfn/KlbF
kt0Z7s04HAbaj+yLN5kor5UqlHHQ8aQszi4vUUr/JcFpwGhuKubb05OKaoUOGHlkGdVwpgfu9P0q
i3/1JToRW/DL4Bk6ttxQfRjFX1d1MmZpLaju76YwaNEVA3A5h9PFxxnG6JWfCiBJ8dxtClB2p6qF
P2HfcweoLzmzGUvnkT5FdvE6tLfrRVF828LvdaYL7G4IQbzEQW0dl0Obn/n2ZAzYhTVn4uxeucAl
CWRIEgvoUZt/PKbpdVy0Esg8gHprintTU0Ze0PkvjF1n0Jh21f+XDmSy85DF35rxpduzQ7HqfEQ3
dhhqooqjZ/Yn6Gu05X33fyMhO1ktd8j8BBuvr7QReWD6FAjs5yQ0l3YwztZuK/zWSfDev92A5izp
yMKi0V9SjIc7I+TWhf4o4RNlCQ7rYMI9PFNiXRvhteOyDioQIXRV6CvdRGk8qENhKBEIiNrD5g5g
Yezyq6D/hqvDBevO+wi4MV+quuSQF/vSPFAiRAfjhnRmUTHu3uvsfEibxp08tfaatRnzGTAFD16M
IO+ubhy6YaEglMPZkkRq+ZbdZupksvlJwi9hnB5hpDYjc/J5+USlhubihZ0No2+aIp/dQdpFQHhF
XHdo7YpOJnwDS/Vbzu8KKXBEcUmwLQNxPA624zExfWUXN8OJKLVt+Pw4eva519rY4cIgIYCHCm3z
zrLPjYDNFT0kN3oQ+ID5QeT1JxAYaTq4MZVEvzY0qat2OX9J0v3LfRvyBvzGOLklQvEHbBwbPJDl
rL8I+dj0vjlN+x+6AZWDtjZ9vJgYVTnn12Wm/QR2BFUQhBkeyPvVn53WH5hkVqhFtmSSk1MZflZc
0BMlm3dGzmgD+WXhBlITRAWVBAJR4Urhu8QTeJJqcwDF6IsACmFZh68TzH63mU6fC0HHEx4wmNOU
+bwqfeMKIAFcB8indb4fyIxN2nOAs0sUBy8BBVlkQNtLLHlJMtrSMObw21SwrYPoxQsEPAmpqpL5
vDziZbshAJdvgi0SskHT2vFdLS19/trbKPTVjbX37byo81eiBJ1XzRlNxwO4AN1dPJyCSjpVN6Py
7iX1JY+M2FwpvROJHJERAK03wyaj1pRcOnQ6p9a2Akp2Rx8gqTk6mqdp+r9XOjUDZoBvuBIO8xZX
d8BebxiYjiXmvgSyWwTc8bhQonWbZIGWJPF3oZAcyqoFdn25nxAnazOHo7pxTnqIF3WXC3R4i14s
oKESsSWACsyYfPyKXNkv65JIPb58m4TKfozeep4PmVWdwulImwo8g+aZ22+DIH9W5cdpNQHKXj3J
1tvA+lo6C8QNWdLqhKlRdQ6l3WErf41xvzcek44MdJygXsfJk8ntpyUZ6p6E6dgHNsQAuMTyVXqj
bRXaRe/0LItmuKiA1RTB3ZxH70l4biLPJrz105Gs1cg7VsvgWQ394sFcQQ46uG6BAXFH6nGmGAnU
OIIWmEK2vgMNf9NsKpDEblPjvsXSbcUmEvPxRMc+8MU+CdfDmRON7EV2uCWggOD9suDqHq3lUuC6
LyxDZJ7WOwrM8UTpno97Tn90R0Jc5fC1/wsW5+uTBo8j0cEkHpxoo/DzdC2uxEF1ucJFA5aDd41+
lbvrBto8JHqdqCmNHJ5OdFfs+TMpZ5jBEQXOVPs/FWH8apTxCsnneJmw4C9EofZgZVZbUMdhYPY7
PeuWc0wxfkbpREWiNjwqv7SQ1+PI79y+tjYRfzeJYovbFiGVYXE8RawTay3HDXA+N/FFtmfNy2nE
lReiHsmg5yyZrY+BGjf4aNa0Onj3o1Ajd9vF0EYGuE0EGzzIvNxo6gZg4Oi/vt9rg4CJoIXoIBa+
+DijenZhULlR3qLJCi+NZQXkK2uWGTyzzP69BNo2n5ogduW0Ki4pV9xy8OcqEBeK2agv6hm5CneF
jWtEBdrjZK2lQK0HNG1P/yyU0tKDuYhYj8RGJ+5rMlrgK8MxmC6nsJxEZBCev2XS+uRc47TCo717
PJ1hKWyEgKZ3SwnuLf0wugS325HXjPQ/XTs9BEd/wOx/M851/1OpiO8QrVt7ho6s4n55pmkEbrwL
nhHjlZQGC0Gx3ui099AX5C2DLUDnnzKIvhSixTP5vYiiZ3SmNvyoIwaV/+d4sUqsPUH7go8SPc8g
5VzR9JZxsrDzc8nxIyPsHx/FOqADKyBWYF3cmZkh+3HIkcHi10ORjXx40y1S29oBR4gnXh9HYuKK
rO/3dB1Y8oaol68Fm4+JpRBIRmBRaBfZz0/hn4utDgJOcBVzaTx0sbXA5SXSHb0q/+J/ymi5GWdB
6DO3uUOcWzR/m0JW/G/FXzpC1LzdxVfYV3jbNUEJu1EOEDh6VRU/4HuCSD+gte0tdXfRF4uQpSmI
b+Y4Eysbrni/1e3fIrky1lgMAy53ygunOe1FRbZ3WFSadSvxwZTUU9/ixWX4XFxntLbaK1nj3UtN
Vv6R+PFXfhYD3Rhvv4DUCbLVz99uOBb7GuDRFR2V8yt3BbO9Cyv5Fs4FaRDQzMElnCjkxXcKssvX
87RLrQmUKMCd17vR8enZMYPuRm17s3XB7bf4AYgjbsr6FeqsU4aFsU2x1/KanK3Y40kNZMckVtl1
bx09J7qUSTCzfeKALJD4RMCXZMsMICIZrFNvXJj2vDXmST7/AjAvIXNr6wFabzU+/PNJGxCmr4xE
cddEP482p4IXfmvj+3aJ6uT2Dk1w5k8R/3HlPRJifW5QUNyGj5SWV+rD1TKTH5hBd5N8NMCQ6pZ2
4fHbdVk1BTfrsDUowHMDCH9gq6vzJNUoVRSnq5WsHRifV58wMI5wN3BNgw3YP1U1uJO9vcKjpEkN
tbRUSiya8LUe2wJHaZIIn9NrhjCpqMEkzydbnHJxvZ2OQRXhFnQ4UCQM4/dp7dQlXHtK1Z3TvK/M
Nx+SPQfEAdelrfocbaHH/Ub1QX8jhE8ayHY5COBfVRggcujjt9kVwnxCnhp08GYk5Xh447MZSvsF
Li9alnRHjevJDh2QUnzCbX33DdFbwCmT9A4cG9a2+OT44XKPVwdOwhApuBMdXpqlmzt9/LAELQbe
LVUQD1WjOHWeISVqFj8cjrutTb2tDXy0R3WGPNHYnSzS1YRHC/3vrIqQ/5S6vxAgGKFv+s3VQUH8
H+Iudv3b0cobHg+OzaT53GepZ84oaTZ3sRcLLF5Ke/q7XfmimusNitP9rdqBwNRUlHm1zKDzSdrZ
7UeAbZ+Cy8t/M1+/rh5INmeqxof2ezlXk6cd52suvWOFXGRShhLqXcLJYqjXGTgquvf82/h05pTu
5Apn+wx+AoOAfvCHjEUkEjyOfNelVar2EKvWT9cKEtkpRjkPH0fXE62rhJuLxd+fxeHpwoSFOtv0
FqjZQqnorL1YVFEXtlRxX6LsaV2BwEyT6uYAm8weFtsw5o4f/1UYwNwzwYIahSisVjKfG6ovify3
YK/TDwXhnoM03qV4dCy7B6vAmcipQcLd76rNCpNTMV5FBmClZKMOv/9fznXV39bN/KZIlRZzetw3
040miQw2UtxPXnYKzCFKz6F79IOZ/A6glS4I5j0IJwWz6LFOM8omcT7fOfM8hWXfbCSRWceyiMKr
bnOguWVZ6ZWttBUfTrcPSziIFOPogSza8KCmRSQywPLBvEfVcM1/NxSrieJEHgpjD1YketvITwy6
czVCL9sugBA75cOcg+twerZYus1WxJGpW0r1+fTuT/Xr9c7sevqNSppeGFVav666VXxeabP9h27I
X6pVMHmhYIG6f8aEnCtgQyaTKn8y4xOofP79uahDORYsQlFGH/Auqa+/qSD+w+i9sW2ubWABRCcA
RKnz8sIuQaX79i5Twx4EfH1P8cllfTWGDh8SeW6RqZJEyQX4+3ncGCLzOUWQ2OT/jJj0JNZlN33f
LJEeZGRR1jujvaiowztkoUBFV7kXw6XcPKTv6325G5OjBaNkMKyIhkY2AmyrB8ZdTcRaxgsIKZFb
MEP2bWiAtx00PW0behxBEZf5q1qMV+GHUJdohheYemFQcRQQa47bHeP7BK/flRs14yjLUH++CtE3
tKWGwXTZOJ5ThMjxIeydiBj+SQIUfgJtUmLCIjp/BRptBcT7STvUYj/pEAMTKEXqnvmcQZnMeWqo
BnkBaiud/nTypkafSNLzzc2iMjme7Ml74+ReaB436qfV4vAIn4V7vNHjVemsizKrZKFLAk58oC7F
R2FE25SjEaW5Ow9Fy9mUN3eHkUzCUm9nIJ1MemjY6GPlTqr0LYsvZjSzdcAEntmvx/udjuxvXFbB
GQwun03ZaYFmmbb8SXZ8/dyxRcdwseIUNHbrqlIRtagSybB9TlA93fTkjsjm4xBREtWacCocXJ57
xzODa06NTvdODhA9TmdF4uApEvwUaEdX+aQyjsA+fCRbNU2xZ9ycI8xaEpjEFhNNP8OVBiuAQ08C
+u/TSgZJekCwd6LbBGe84KuvuoVANXaOTvfJsrGPFBRKNvaGS7dfcCbxxNdzpxoskzi6lP/ersDv
y5ZOHQyx2YvL0Tofa7idIQz4t/j1nR83evrK4E26k2MS3drSP798GZYgY2cYUw0CgQJOC0Ohn5H9
I3ruw0ldY/X9bIccYACqoFs45HcfSlCSwcmTmUJhC2POetTbmAaPRMj+8jj51tBilzr3qZRxcOrk
Nf4v/IcYSKV1fmKFQpVtCc90I8fZHUbgOVKJZYD5wMdihvDCqrXI7jDk7DL6gdr618CXLOuL/uG4
a6LAABnoz8V6qBRAxxlSyDygEBERzCepw3IkizlIwdFQPDE7dcuBOWnlsmgCOeuwNojdIXuYoPdP
Z2OVJ31JOB9aPSiT3aEHcwP25BKFyXWAkhcEJLEhyH7zcWavyaKLPXWiq0CDCctctOBLsJAPEYZ7
OpBOvd87XP3QxtWDEYmKj6yGGfMSGG4vkOkN2n68/e6gRPlvS7U7XF4z9tWw1L3NGdp9lXOo8rgl
EVpFSEzGMiZEsvIEEog+3ShJViNrDrw0HREkgXuCEbVqUMPu0NV3ezyCQugzPwxOnkFZtEDWqeSZ
QXQxaykYnYb65P3jcisrPZKiyR4sroFp9BxNmrS0Hh36okEF3YemsY/wS1zdx2SlxRqkoGbBcIrP
XQgt/9zjiODRIxkDSUHAdANckAe6NRCagcTwZzKfNH4aktY/wGHD7tPpDtINfiRI+Qw8XB23f8Q2
cZGssMPTuTANeznaU2iJdNhCChwjm99uwNywD7RqUtHagScJy3hVFN6x/IT2pBFC4BhUcMUDFVYX
/BaeoF2UzZmGwReYxWuj9cvMohmerJ9MU3TTQW4YkFQSYE0syJtHL+GbTY6n7wUWw5V0sonOEeO+
rPp13CcaQuN8ELhOJJfAp/G29jadRwqxPH1MLIGt7AyRyIeGV12LOmBzrCCZlZ3dZTvhNVoPpCuk
so+1vgZQeUmh7KSddTq37DqJqrMeQlwNlbv7HDPXB7C3w6Zvg+uWmxbh/9kSWk8CAlyPqSNx8jwW
lN4QrzJC5uEpGVnW9eNY6CINSa398TLV3Zd6hg5hT8YxpLZcMTupuZZeDTuAm7ZtTjvlLdqaCpr1
9OzoONAOTPbcAmdOzu4cipPRTM7wh2NSjn5bWIDctSFg7ZBET+artwlDPV5/lohHqLl4xS/VVlfu
tmdjLriFVFkYyPWL6K3IvRd62hYIG05sCWeUenqxTWfSRO3xEVUyvqjAZ+AK9JyEyCNy3k5LScp6
D8XlK8Z1iJ1/esjjia/Q6E7TnLu08VBwKpOXwYSMqZwrM2QFw3e2CxEVwCeNt37BTfXEt+bUX1rC
S+OLFAZ4LI1yKm1h6dPU+k7VRB4On8fBRyAOfVnR/6rbMFhboJTCad1T3U0SqkjXgldK8x0FH9/C
/c6pgnFbuSH/fSUggNFOMs8N/3JVS4ssW91sonys2aqnan60S7DraRY5+GHjdKUQwT1a32GaoGyV
w472gVU7lG8zG1rbJxRjmHZBmKNhIk1yOZuEhEOsEPrDZHL14dod7c95nexRpYNM7Xg+762mqV9T
EI9yz4sAf5+JGJnHQyIbYOVWN31xizMC0o0AMnpu6yrMGAKqvl6lKn7TiX+dvXQ0M2b7dG6qNfwV
W5sdYyXfrYr+FIhdBqnfjV6gwUTFY8VLBPYlwdEebfC4ol8awRp3sDYdjrInuE5SQf6Bemu7W9oe
8ySyyx8+IQfjFN5pH8C7S9GUU0ji269GnbylUlcYGhtkdFwUpSpX5zs6XlURMk+SQTiS2w/455y3
ly/mKCL/4HsedfQZovddIRurS3GgWGyN0OpGInJR1m6E7ULcGSQ3jgBU6tleruitUZ/aRGtmAzwz
hUfaNs0k3AC/2IyWXwKrN7Ob/BM80VrrIPoxAbXCaLV3xKndplKFTkqBV10J6okfluvcwXBhbG8Y
nqNUTZtVIbJjEKbXvUH7y57lHLlts90mSTGYgjf9uaW76rGM8ybdn9gXq0yKjnw2fzSa+L/Em+KR
/5eZIKxT0fbUteAaiFNsT7rX0edtZ3kNfFlX4u1LBOoobEKpbq7RGpx+l6fpgcFpkdTRAuPO5L+R
ahhmz+sAnymjN4uUCpJIi/B7FaryTi7RUf9RuRjHDF3Dowqtzzxym8fmOYcSqrifGrVLcBGicduM
oG2DV9fbZaw21IkXDDsR83zAaC6R7xKXFYvwrl73zNmd8g21FdPrrsVWHo5uABXZxBtrRzJz1iKu
5QrPHymgvdl8WTINUXJMu/W0g9b26sjScjLsfZQ/rX+RG1n1RVbt6VqcIzgW4T6gQGo7Rcv0oI5I
Cs1dlAfeEahzFuP1EmNCTd5/kP+oQvq2EI5aS5u/SiK2zgOK+/g+rw7Jh81A3cCB5yYgQBR4SpAe
4DEEo9ZrZEFAB3O5RtLnvcUNfmAXZr3EBw54xLiFA/qfpJY4MoWBo2m8tFfDUFNiroCrL7LBDLaU
Lxul4Wxm15uQu9mJ/spA+fZ1pKTqhCwhke3X59TMID7xaJfSq6Cu40ph7/zomLnfhItr/xUASi4R
/hr5IUYPjp5NK2IKdgrYwQl/WMECmLaa9Rgp5s72OxMr1ap+D1cHybuITugXLz8XpmG9GlbitBTD
tRQtVhWD/OB7JNtWqM8xs+mL5BW9tpUF9BsuH9c5I52HSCuuq24bd7D/T33XCA5O93C7dgIqBcLp
t2F11zkx6e4GmquWcFq3rAP6YNN+jW/Bg1x8JHvd21AYd4V1roH3iVM++TlS8uYTy3MAB4ynzxK4
kvh5K4K5iJ49zPTCeFMHVid5t4VuF6Q68xtDuCvL24ooySYNHv2AC7JHy65HqboBwmUOdkMPn2SK
3hf4CtSOfYNdPeyxAf0gKXilTxVQXuKrWQpHfF7Xh87Vxvn6jbO/5YBijg+u6t5GyZ0LA8FJkAPQ
v/UmN/KuK5wHhZUMvYSzOEdwOv7gVjafnxUCWqUBIajfSfkk7euDy1I6jsftZKzcvCWP+GKkmvv5
JRtLpPWrbFIKAGYJcL+agVstHMFBqrUnJ1UCDIAkPuW9RaonKveW7/0zEU4jtv+kSeZJm3d1VeXt
D+8upxluSH86WSLyiNqK81FNRIjWdq4lbNqH6Et6dO7fssbRsrkFWMhYhzkVgmlAinZdUveebJqW
DgQxnug3Yam3VF5BiUbDcowGvyk36L4yJiZjMlHDfEcgf04m8Nt11WRRlUOQMmDzjZN++DFLg8Df
kzKPQ9fyZRwlfVHE4Q3yyY1hNQJBaaL8siZr+bakqPZBKj4Jwq1cUTaltLhtlXdsZUNGUz4YWLyb
+suUTF5M1aYr9Y6dX3YhuJyONFneBl0j1HTCxcy4ecFjnnJbEnT9eiEskhG6o0vQuEi9lDyYuRKN
EReJgugDAQ4H8HSwL5s8Hh0jtzs02ITX5xV6Vw5tzdSt3MfiF8svldn529844hf4aA9YyJUz46E6
MX4hQO+tZOL++hQaX5hGIuWFTEfTY2w5bwO5V+DZVsxOCH/LZJmnCh3FCeMisEER9b8ifZiek15P
eCTk/4k3GsKemYGi4UFiiMG2ej+biOtDWDgJXES/cpxQDtEy4zNOLYi/k2Zx3PtyBg/GZZS6jCMX
BKcmshjF0WZ2D63svKMCcnDZ5e3LE0H6yS/NnsKDscHOqYdHI6oSGNHyQYIcdc/itDHP9DSxemqa
AQoaIAdBf7qAc/h3TfoxxfxIqACZvTCqVoG/+WSf/WdRZxpAUPOwYYeY4I5KZFJw9lxF11n+BIQG
HaGTIWvv4ClfFriXPs1jxQ6jqf7iBX9op9zvoG49cm39p0qMa6uC+cEYkkK9/YKllabKDW/a27oG
MdDKYJLfcA9nht1IzhfF8mFwFTRx3boMIZ33QzwGA8Yf76yfSHdm6TVWjuTabWm5RYFo/J5GBYBQ
HqowQ68MkKn+Puiq3wSf/Lqy8sJVWJBEhZ3KPK6cQGPnAJdGqTkgMsauYYRvSUIbHmKZ2meri+7O
uHU2PvMTbEhUQN9TA6iwlJUf1/BwXNM+8/MSDE640rvZamgoTJdpGTWj+jSss/Lq/B5CXbsNtaYS
KvX0BZNnXl1WJginjMVfh0ZrwM0APKpMbsj1SNo/PWVCMIQKWf1MR6BvF9XexEyrmn/JluWlXyhh
n8d+XsFAbveoAI8z13d2iwMF5vIdUoHou/ESKjpA730wfQ70qpucBox3npaQqw5WrU4nBYYMWbJ+
UDAnGrzA6tHnIEFHgI/Wht6QTfjOMWV3/zfr7nB/aN1WhZ12zJ1+Bkx5nl0K5Gx5LU/7fxmtBW/i
sxCUW1xPjM+RuO20vsyaEvqZW4O5nrgeOZJSmyaHuiqQdQ+IY1WDfN0UnFtFpjBrmCzUUjQn4eI5
4SHWpAkyLd3iBn74784pcvzmPbQXhf5O+S3tD5b30H44nKdmfcyIdXlR1LExF76p7V09zKOZa9GN
fMTbFKbS+FHJtCgNZeJ1vMGxsZH9IMLEG4xv+K9Kzs0f7W2mMRmLQ9Y73DXIWnwY4SoPBwGK/nt0
Yf0HVENDA1vUwEoxQFjTB2Z6eNSPnKjlk8L/7LZ1QMczwXBvl6/sewlVud0g74F0i3Kwt6T5PolP
NYly12ZdLQyKQury8hPmLVZVKEQ77HOQbYZ6VR/L8izfR6nbfP5bRTfs5owgu+TSXHk2+bdx45hI
k14ndF8FALEnFhimv9VnJTfeO54aGZbl+A8H3mKn+R0fBsfX51H5RyoNb6GGkwA4hSQW/YPEzK3z
dAA9i1pSxQCPu+x1b48Cu5LYSj+cIYh8DyjJDBydCu5vYROngsDPHSxTj+FW3Zb5/TOnLjjS+TEd
rH4OmKsbPXgLOKUQFkMgZowmt0SCGLuimd6StcrOMbdhCtYmO2VodBMN20+LK9sMyQINMyNvjyX2
u5u60Mf2uB/kormXE6ZhsGBPdxlrGTbcfZWrCto+3XQwvhFld+ezlALJh7i6QQ0olPfhFjA9fRQ3
gs3DnF1g+GAJSZ8giX/zkX5ZBpiOnNFofF1ZnSE/peYGy8ZBqD71apfWhIIoSdZIcWGP+idfrA2E
Cntp0cqOR+aRs2yXuFY3YwVxMDxPeZClgyHU8wNPzChsf0Su8MrcpAqFpQ6/O710YMITCR0VoBTi
keq1qbSfadzGB2A+nHlA2Uf5lTf2w2PgTxSr8L3mS5llRDIHOC9acHrB51nKSs+QQlJzKP2FRAZy
QDeWrcUzS8zXrI7QvCIJ6N7PHDce/kXeeX0HrQei5p23xceyIC20lOuGC9UsO0V7rYXqBqolECIZ
HIphdel6opWMwy45P48RdcuvUTJJrqtV9ywOhZVMJcrrRHB79VKATVLMl8zGCuH8n8c83fBRnMzW
OeClBI31UYFDk8xaHIvp7/ANZGkyMU25xjy2R4Fo/HuLMYGTu+6XLyCrt+q/KUDv9sG1AfmqvVmd
3hS62MFGqfQG88d5mNQgZxCP/T1LcxNYbc3LxvTFTa7SjdpY8ljnfEcuMe5lP/hbngXzACq4gSf8
HFTsYpOtUzPZKD5zgcRwfE75KvlJ9M/OqQ4qdJtipTJ9c3NOJr0aBzMuccVnRQ1aE0Zjdbd+oQdF
zMkE1Cm322+4hNSFMYsKX2rvucm9D2DHUKUaqmjmVpWKsFyl/FqJVy334xWnm1tLYWy3H7IB3kxu
JawsDNvM06ywJjP0/QptV6jWzac2UBDYh3TzN0nfRXzh9wmex9v3XnmBlgydY3iiiNXavrZjWNje
N3psrEevbErxYfi2gJdkJmEVGiANgNScUmmp64LShCUg88rvr1Yp1wB0p0+e89iY/9Z8Iy/cM4qg
ntUPOD7mFc2O5OXMDYIDCgvnH2nzwcbZ+6d+YI0YuWJKN/aRz4QKJ30DTxBfCw1ISruk46nG4XWT
4joyLRWtxB9OkYo99KEn+aNQrYo1ILGzmGKyrPKceh4eSbmytpqatFKivp0WHs49fB9VyxYQrGLf
d/VQClxTEFyIhgV/GeHPX6rR52miToeyJBk6CDgAn0KBlzqYAw/YLN1Vh35xTYpaUbAiY3JPkRIY
H/BkVzEie/ocZnM5lCdC3pJAPHLbykHAkLHqYLyAlX7U9P3rHus42bwiFysyX+zz7+kKlPUYbTZF
0ObhqSL/pgBFhEyL3jFiopFy7QEjQkmCkz7fcXuy1CEtqKSOd+9R8UfDBZos82ofhgEe9BxNsIry
q7fV/V3N1EdPKVubpVhYJzvw4K5U+qCs9YJI+drxyyNNOErHWKp4F38sK9yGv+cyj2lW8J423n1h
kaeNLzwftVG/j08ZZzBV6TqsKH4W11tYQAu9CUaESaEcOVsZbkbKczJkp1nC7qNRCkeUyim5axky
l947G5iTBQWsXcJKAapt0gfpzVnSWiY6BWAWHheqXQrj9v61CgcjaHYrryu+glspBI7Ku53sAXNo
mssrBo+j6yEIFBsIJrqL3Vrz85O6QVmnI3AnoNZEnvyAD41eowGBNny6w8MFvtleaY3snKdKCVNa
m0MtkWcc7KNYcZ3UacIZ/m2IUZKFrc3Z3MBiQWg3RZxGrt3Rak4U49X++p/N5OKBlVI1aPmetluq
vzw7R+76/OsbB36ZHpii/SlaNQlqbaOWl9o7wz1lb4T9pQ/nnj2D9l6DxWZ56t0jF2DuAT8R7Gc3
gAKkdUIU222qrUG28ee8p0QAxxdk2qlmg0Jaog9xIRomXZg2Qnoj/1pAyY33hRkJeJjQdfPzeLi+
SpB1HiuO2Ua3fPa7Bg8fZDV/Cwg0FHksQhQYMl/llB9RuIfoUpxh4ZIr0YghNqg2q2Fh7t15SpiP
GCL/r8K1qKx9xuDpVP3ggc1T3mLkPuDSLV5O9gs2KpaQPtxcDunbr0G+5EYE8X79W87fglLmFLPO
2Y/06ogWwLTuXv4xEUtHCf6SZSzoCizlJsTjRqn+sxltTL/R1xfvNx0XJupVUVucs3HTv47rddTP
Dmt8/55de7gN7D/5wmvLKX45ol1x4xHMQJ3pSS+WqvCkNYjW/VsaxhbTEQekbQN56RK8ZkRNIWb3
IZxGOVT0PLys2d5JGjJQTuuyg03wejRCNeXE3dha4LP18rbAGFjt0mJjhia2vOzfxCXY9PJRjWv9
zFPXAmg3qMBFZcqrads5+twozO1tMWYK9YiMs6k56zJZ6SY/E7fZyjLoFPCMn9KrQLUDNeoiDQNU
WiGaO4VoTnXtDHm57AXqa8TL6/8J3l0PtoPvQSZC/wQUQtqtS6m6HGo/Rn2+cuXN+x+9rAmZmWSl
HOp72E9wQm0ZIQa4k6culGuowwHUE254Y+Yu8GpMnkCWYrsY4VHb+KQKiTmcK0XmFP9Gro5puFs1
IWZWdkfpXJ039hfA/vMR/vs7FBTPp1xJnRJbCgSVh+FfrWrzUMMEwMS+j+MatVImfPx1JWg/rhvU
mWPlh4BmvbJlNHrkqZFUAXDHLKB/x0Iu9hvVqjulHylKeCYgJyC1+lwc+Cbw+eEFXxtaMXUg/eo8
omK8TIVKNrJS2CA6GT9UjzN2fJAIMx4iOzSGrfzPqU3hD+KF5bYnSqt0P0W2VaLua1nj0fIRZ2Pq
k7D38rIX/7Rgs5moHUdAnsg6+b9itIn/360umOJUcssZPvoju0bERBWHHHFIrSgpMianRVzldf33
y3PmMW9ucGz3E/HLB3gX6SxFC8lY+2HRrOl6I7p7UdTANVfDgzXdm0lXcRHLacwMkejJjIrGXIjc
9CaSyixhZiFzHp7rA4K0v3V6fmmxyE3LmRkfMLcUdpsGII5KR+6XpcRDqk5eZSpEJ6+b9KlAebwM
meZJMFv2A2TmuJYHCVnrEB1xpCMF9OGDjEW9L4U1MxFIS31U1MpSRo09w07wMgVeP9a6HmVu2IIR
wmmONYCxRr5flRVT1F3qfC4VkjLBD45OLRyTXRDpdxYTVtBZVsSyWk1VwAR+E1qJbeyLCcVmjsWj
ZysTu3FxqznQCseziFVoFCKTJ7oKb5HfKagZxKSa2/G4Mde8ILbIYaQ979OLO3aTQci8HbOJaToj
nnnK5emob/PNC8eNNhiasboPvaJ/4dgT/jIwZpFdWRicXiRZwsD4cep2plarf3MVOBfDedyD9LDp
KiSKoyr+qgiNJEzKTWd5KzVVkYfExgVf1tVepUaCMghyplnFW+RFVJs8dBUdawWUl9pHyZ2ZGkFS
DqPMgaT3cE4ptvOyGnikM/PLjulqoQ5RHVJtgnj4Zk6hgUm9Bb/nF1Zyk6RTGfyXnSWwq3dVs5J4
UKnlTCtj+3u8NWKCJbbp/Q21On7F0W2N0RTM7Qn/by5RhpWA/uQ+81bmAqmnRsZVxt3l6MumoGYc
l6D8ZRFQ2oXQyl0MbHm5wQyBRvviXgw0zP07j3B/EcDCt8E+QCMgtF3bdbPNwwVcTqsfsBLvQOYa
DNcYprtFNEndUgD8ZiSUyVFuVYuDethM43ISrd8VCbTEhOMUK33ZjIkQwzjROtBSwtxx8PFUiUV2
gpQ3TQhZRL/HvTWk5QucpJv2heq0Wppq0kCBP0Zm6bbn9ggWr1a4Ce+IQOoGZ+bFsShVyPtwGC+J
81g4razg9P4c8C55q95wKO2nH865gq8st9QZa1m9LXhPURwIltIQcwVz33JX5CdAcRIj4Pgr6n7G
495FYgNWOH7AyDTzMhkIpp5A4I8RXWal1Zf2XwGLWhmcKqw0metvth/z6EfUCutjb0a3Nzgsmi0Q
PwdPDBy4Ic72R4DT8lvqDa9P4rBD/GuoIGk6Qf7084B9JMk/YiBXkZh2aPf3nV2xw1zLSfxP27yq
EP9/X+cKZq9L9hZCdtC3FCTzvk9WeJ5ULiA5C1JuoV0KT4bxdLX4IfZzzZTkmCh2f4Bivy/ZSncH
XOrINR24nyAm/e5lto/V7qggikJqv7qOCGI7pfTAQVLAqTJJpkTZ7zvs5kW4/McJDzP4EBCdeO3G
Z8PzN+zHblbcNGCSpl5ZT42DbCpItRNQMs7D1sxzOy5dBVsz18fKU3dQU18m29jrwr74UejAojUo
Iq6jvMqQZEOBjJhfZT01BtFHVk2UQwK6d8rVKZwLs7+49/piBoYmtI6STFP9JyAcXxnhXa11czep
/81q370aIHsySkc6Bj9srdaGMse/usv3ahrzHiflgJyLQjfhE6hz51vlF+nAHCiJG9HnQnpNxLXN
zrZpIZFToJvSUX+l5HtHPVaKwNlntUNgWMzR90hcTT2bSQioyPAXMFwbXztnTr4vRbGCnvZrcMrV
a/GALl8jnNIo/T+jWJdtJ2c7ulVRDb64F70Tm3XVisVIzQLBiu4ZKtQf4SJDbBFsadH6HjKp7mKq
Ny4qGC3STw5vLw5QbaPyEFK22RZYVQE6VEVX8nrMnCPAeqY0+K6B3Bvcb/+Ikyb5BgrfRU2HxkwG
cFi03URU7nJg+64+rcP6fgF4KDG2lpqEAPvlYyV4LOzovINrcaCjw3p2xkXMIkDge+INKkeOUHWW
MA4C1wejpGqz1BPkL+qvq4m6BHFS9uah2J/wa7A0/w0DgpBzBO7gXGJBceachpbTDjC4DiuEoBke
VZGFOylNSHyKlSFmi0x2WwHTNrBV5ue3oTc5zl2v336S/xUKislkUl5w2nEOqlsX+P2ra339ZnXR
n5aOMDi5ptt50eKfB0jN8NT+W/TKRGRx20JtSSg+3Nnxd9eRgNOWncp56B3ozP0vkCAsHGy5y8NW
neQHI+HIBmdC1KNn8YBSqBhB/jaVCM/Xz+RCyiiON5A+Hmchp8IEfmoFioFttLxHlwtSuDz4YX31
Y6dAsWSIilzTEoQnx6qColScbOd4zFEdeKqeaCRAX2CkG1Y+uDOSmEbfTgi3Qc0VSEaVfnbKbuB1
EXXMUiBNUbrfKEJUrxrKcZm/OM86+K/hNc+9luH7X3wMGfydvOuPoM/symis2ddAcCtlxk1QMKxS
jgqct18aJd/si0PmUEHxnC09xj8TvOpcbtb82lsjxRmozBJFOqHWzBZxoHoZRUn8a+AsN8JoyvZx
b6Il7Ap0BaPXd264Sm8yLeZwGo3kB8pEPWuW3GzVhgVo/g1gLS8pCVJzuHszoNQ72gVV3Mi+fd+V
l6ONId+sGv1l9AF2Hp7p2FdV7413hYSjW1gH0mfjgYho3WOgtNVWjrWYvBdaXx03hzpY20/rn4g3
plUjpeu/xX1DmWi+1lTJehTD2xiWX79lztRjuYYxYBEqpaS0ZBxndQt8b0Em/t1jjdVV3sl53yJm
bjFDcZoQCE8JLPH4AekSPDog7A46FCCD9ktOogonSKlk22J/jPeB8lohvz2QYfkL9+0JpoN5g76F
w5z8mv4PjFqCKNZUlZy0DkfaHYQcQYLJ/6dYioRrBskz4udiwokLt9F2IGRh1NezuA55bCOhLUGx
7tAsUOtMBXpZXa13tu6cq6DtuHBSdkEVqH/ms6gtVIz5m5V0aDcXp39aAstIRX/31HUSJXNXIqdF
Y+CiU3T+TnYbQy+4dd86AbIOaM26/BLcPPh8YZhF9gM1yHS2l8ChaXIEscGrB1cW3FJaM+dFtwuf
UsCRCO48MHkYaolvHD60Rhf6rgcR7WoL9BnA5gCkUQnRLei8hU2jVoXm38WjvAokGKGotl6EBVzu
Hgx5CVgXUX1jQIuONJJEgZsnJVrtY+HsHLCh7c34zFlLtpXh5gN43tdodoVRd+VxMqQqCKbLnv0V
IqUYVeciNrDu4agn/4OaxcOiYktgfkkZkjsXyOsWorbwUuyvK4LDKZ0scNNTwsUPuP4fJc3j8+2G
utnvnPrDJi+lChHwLjg7ae1C7DKaWbAJZ3FMFZMClISqBcLeXOnXFmiUdpeqUPu+qWWqcIwIDm9c
ydgNiCNHkUx1VqJXix+1qoxvZTZDlAJYpOnjYzXeTWG4vrvLupB+BF3oHP+l2MzeNJuQ0rrSma/J
RICRA4mNOd/OZC2rMAnbivnUXny/SQpYh+UsNYRFqe1dSe0R5qbp32cjtRQLRK2Y+QXGSTxKze+G
v3myQVGvTTszvI+35nC3llEibWr+acIU6i+oMFBk3xeiGvl8+RoTDX9uMEhpaQQsbcC3KYyB4hJI
M9wrISD9zIe7CDCWUXnaXu7iJr9nVRxfqoRui0pbSQVI+r7TYVnGmxkVS8o4ofATiEG6uSdGbiVx
GT9H71Y4a/RU8eaPWfvaN2jA2+fxrJkVcTtaqY8vOiQkb1eDlKKdAbqiW1XyjtFUN7badr9zIUW5
51jMmXyzIq8m8OFjbW3tS/SrYH5jWBJzux8XF0McVGgoDNgXZD2cgdqSh5lqFgwrSTjxvqZA+W4/
9knnlRJ3jgci+pnL944fUPOl3NscHUKaU6Q1E5MA2VnKmvPPTpjYq64JLlRf0KUEdhL9ItTI7v8a
rnNQtDGEQ7UG/B/KrZ9ecTM16GjoPh9e0Jr4293g7t4aC2wTiVfp6nzwUvq7nSjm80b9UL2e5IGd
W1ON2nCuQkdzgSib747QbEfHatgRvtV6TEoNPNmFlN2+a3EWh1q9orYwBfcIatxOKIcQEMbzgv16
ekcEqpYxD3YS7f+HTfnJX4tt7SVijfQVRaLlwczgn7ljos+IMjyj4HT3HpzEBq7qVH1mGLoYzVGe
IkOeKOY6Hrrwl2HJCRccP6/IHuyfbgEWZSR5L9EtIY0ZDMOYi7KJMAGIa+wjJYvHy6NOSWrTGYud
pUM/gr842FDV0R92VwdC6/cqBgn5tvVy50+9pfHBCq4wYK60wNYDmrcziMFRQJqF7u4/7CbwtmHU
TpXAWjNEalf0LLSfXRZgysBiSaIQwWD+2zRWsye2qhQqdm0zz4vDfAICfjbqBqnuZSA67BUEjXD6
vTH2WWOrRby+MI/RnwaRUklndmv8pr43Mr1J01g0WwIeD0xkUTvPJVBjE2BKfXSFR14O69N1WEz7
4xgtwR9VsbsDhplIjlfYHMEs6dZxpwrMKjhJCQC440rXtYOUs74FLnmUF6e/Je+3WbNVfQAXGlZD
ZnfTQuQNdbuGfoFQqldHG6Zia+StmSJJSmNbmEXvIt+NJxeS1U5QTyfpANNdJlRBeK3LtujlNt+T
QD2/Qew6ke2qQawIAw+pAEIezpK3l3MUibj5N2IMn7shb2DnIl8e4hFVQVpK9yOzx5P6FLH+ZyC/
gPb8/AlGIiWPUDYLj+n09PYyRtFZmOgf7Zc4D/D7pchRwFftaz0k5+cNwzmCL4JmmC0v2P7moFyD
kPEtHIqkuJ3AkW4MjFh+gxDv2CTPQ423WCUFoEYxmTKOI+ibJZ3KxBEWgnol2WqYmqGz33sEny/f
aPSvdrsU/edKp3r0bPPbREfRF9GVte1uKPjAlvg/BozESUqR34XeBhTWeN3H/AoD/Eh9MxakCcsZ
3dkI+2XZ+GkhRbU0SVcezLjWFnSFHThwFdVZHoaybl+zIQDNPhSFq/HIDCa0xvr7yGWU7RpXCb0M
R3pJHWMXmX9h6F74OX2InuFOD8iuc+RSqgxPLhMMgE5tNiBBZWfSEBaFpNCXZBtWyaPJs6RX3tVW
NPO25WbvPRxQBF5oRy0DaFy/tAwqo3OhGKEM544fQbFaFT1QuyU1qPx0KAf9CZWmTAjwEbal8k9m
pw16yjFHGmj+PG4MDWeaX7o3+fbcrJ0SquOjdCQ+48MyMeuL4IrfCVlQP6xS8xFGBDX27kEnLHfP
LvK2wXMqLONBYrReS/6zJBitPXiCpP5hm5azw0zyL1sOKRwSOEkl50xmNoOxmxJ/YZ+b7upGT3ua
15WeV5B6FXGYkd2Knyi28RzITrOdcpiJepuUuMSDXsVhzI7vlaIBOjP2cD9MamyxBr9+/KHerwFT
TFo6IXwCuDVJPvVaiKHFGLSq1Kzzl7aUY846f6S+opGEJnYy2zj0usC92GTjCUtEWannqYPO+CNF
1fjnJfVqMhH5iPWyOqsarohDAsj9GJ9Z9v52q/5Il/O/j/m0DXgm5GeCGo0Dl2GRAsp5IWOgyRwA
O+gUwbAVRWZve4v/K2lxGi39m5H3Xo9EVx/rfQmTrIOj0TfSYcZB/K+gf1yHEDiXupy7qQrAoz6S
7HjA2Aroy9CzBPSSKkVqDFxj55sKQ10lxk+2CtghuXjsSnVfOnU4TIppjT9R6+TwhXdKx61qL6lc
s2GtLF+SgNtnr2J3PMoSUwBP6HcCeN7eFsdmhAoar+I0wvYdVOKU9PK5qmwwC9WFSfHgYbMzKzVD
jXkiMYG5N5vWOEEX508WI748AHBg4OB/qlS7ZbHSC+eCEtbxR92+FzK6zGUp16tXQyY3tR4V0Jw4
lYscCnE8vrFIyEX588ljBVSyNa75gyynL87grCFmeAFgQIWKAM7x+J6KYbu9it0PabnusFnCJ23h
j9LNDzd7JkLdLXvrxMGFu6vhHvS48Raq582r6dORfeknCohA58kIj8W6TDM94jtoX49ck8Y1GigN
ULmSP5g57EUdGe/Ju1lvzTdEmqmgVPq5TOSWHHQHFLPLj399x3g/Fg3qesiy677dHgy5rma/fKex
lZASSFkgxPRcGFNhAAEwt9sSmVSt+KMp/WUYH2C86t2pO3lFhYlQsU4h4vpwP+YgOVaNPj1+iaqe
Ow0r/yCvAmEC51YEJaCUTA3gecE4lOnxwBWdmBkQnHHR+/PU4ACvO88au16aTyrk0cVJqYRLbYNr
JMLLpF3SEy4Rlf1Dz2EImEAJ7r0yVIcAoQwWACI2m59ZzDgcFF8Qu/b0n32mhjc24NeQ4OBGv6+C
uXVYAAiF3Y0c23lr7dhemHv54sCdB0HvX1umzbmSJCjMyR8rizS91HwNy8eXVvEG2M8CKIAyuvCv
sjaSRCFfhDJ1RcpRfmUZWNU2w+HBOa7wGcX4nSu3AJvCkMwseg5VSzWj5JX+A7QxTAnVfyruQVlJ
7GjkgytZ54UgeykYjIQ5n7Q8KvuWg3jscIByKaEn5GuqJ8ugA2KdE0nHa9dXzgnj/zjMbjG/wVJL
BdWUQQWKVWzdN963RyLIbG8qwSW0Ezg0iqcKWGN1ZeUYA52G9A53ljF6soA0p39Of0TiqRMYuBmA
giLcFvijT5t6tFzRuYuTJ0IHOLC0K7+cx9amFNy+2MVO6rt4UNuM29c5EEohA+zYmq1rDMNCy+64
UtdE8MEOD0DgYmneCssB6qoA7Dpsjhax8TGtsGieRdm2O47bJMD/2KcuTIa00orly84DmLyFPSYm
OzGmO8HFN8/xZod3DCsO1TMZ8v15F7AlliFolGzwVcThxwQmz0YcS0njRSv5c/PABGixAS2jYZU6
asvHGe9NKFEP7ahFbE60A4aD94kn6PMzZHX6x6Msz8/q9L+Zh3sF058L7WVS8AMAvIl5nzkgaQb5
D9nNJbfvOnL/A4xaUILqOlq11jV27/5G09wdiDf9NPeLxU5QqX5C9DyNWbZCNd/W/7MoXWOsMPhh
+Q90XL889eUPiQga21Yrnsmhugkom68rxaqDDYe/AIIR3fxI0gkrYlboO77hj0FrOWt5prFoOysl
NrGDIFOrMUALRO5G66+jJw2A3q5ZNkO0q/Sy859KNGPryvKKQpWgRQ7BZTOCBpqDXA+nmhZeMC14
/3OfjD/S6aww4yfmFvl6XQpfwlqBw3Bs1E1q2IjH/CAqxp8Ay46OJzGt71f/qMEHRm1cDrIo3Civ
Rwq8d/NYZYnj4v70bg1cAlmlstARfzL60uFlbxZ3aiF95LTOh1RXFCRiH9Sw8XNAQjgBBgojJlj3
6/cSHXP711mRcUq0jcEegcdLomgq4Ul3gu3wTL55cZCXU2KVB+KoaxQJ+lNv00BEAr19x9Thgvqh
z06B9gzjfT0BbxZSyjDJR4oIKovTWUuN94Y7NzqfS6dVh8AEsrWDsBJAgjRwj8cO2IIrTMdsmrXq
BRPeQPTFenbwc+MTABjItbbaVhaIRJ97h+LBoIMbvmmDFmfiyVun44DxQZhi1Nv66mDKbJ7tEsq8
A/sAbVI+HpbTCKOu/TY411moQ/sWwjklj1NMVSQ+L8ll2uZpxKeciGHHuGXmJO20TQJDa28dkJvZ
6kuJhOwVAUQCNbc17MhKWBEokRSHRdQ1bUuWIPm88X0ws3S1tZv9CPRrp6tMmBS3BgpPUvlmbbcK
03ty5FbXzjD4h2N0pTNsewFgkm7AO9g0ujbo/npfn1d40PWh0c3bVqUe/Zq9j6Lsky2C+RHQoMeL
TT00+wjQG4HAg36SpPl/L4XXUhsH8sbDb8yiWYktQQI71Ih7Mh/xxM7wMDoQFd0+87XfObVHj4F+
4pouQjatZVQpsIklhuBTJIzqyWFf04z4VgF+AXrya9t004A1G8OxUL1atipJs1nRJEdrw/tm4/Ut
a+aLvmChtpg5yqrEMsyCdxh2Iy4YSVdOWeoyzviJDxHZ/gn1MB02K9wi61bMuAxGlxkaLmuVmoWC
4sfAiPLlDXvvUU3ydZnCzTf4i26RdOp9C/KT+oBtD5V/cyRUwXm+V8jERRVIhUTEFUYta26emfTd
LOiVBP6zVkMJz5o8261XW4enEB1QX2tmrL1TBeMF+itkpWaq+zASQCvwf7HGfaIyFxouMp6Vq8T/
gBfd5OWGfXikrN3lJA1YnMbm5biAWNqa1B8QHrNJiAZ7cmRb3oa390AEl1Fq0RRz7wqA4pdes3v0
+TSrdBmd3KDZgDCnAqCgDxYJefbqUDl1hNykCxjvgwBkBtcpmZZnL8hBBXaCnsiMGYp2v0Wh48Vf
FlQwJ2Q2K00OEjBrpXyXWBe0R7V2wcT12BWVuF4fKtfJHKOiqtPc52pEP6q87Fy6dDn5jb9Wbl9O
1xnNua6cO1zQ/pLsUt9cM2dNoqtPFSVVJoXEcHpsW32wZnCZn9ePbDiFa3KMMFGu9KCsrNFp+D1G
s6hKJg2PkZ/BEI9grYbmNJ/0jv7GTNgeCvYX8HzRGcBNZ/OwgjA3pg6X+m79Ypv9+nBo1Nwz8+Hj
hwm91IXwyFHnwyHU5QTzN2C44Jwh1IfKfnBWsBL7sjLvw6wQp1IFSxKDzZu032h/vz743ZBl6BKx
EZ4G4PuHSzRvx0w0doCZuG9NBeG9PV0Bg62hzfuQbHGJaT4DG6bigG8hEVNr4z8jBzXLsYnUWD0X
uDpbJKz3ukwGcyZ208LUYpjhDVNKOM6KZ0teOKHvxVJfHDPnbWtfgOK1U87IqoGOcC2uOORsix3+
EgyJTJ00ARbpFQvCgC7PXcLWoBRckOddVdDF7RPo6zg9JTv7a1qCk99KSqQ5gNw0T8z+dg62t5v/
KVg7ChUV5nOBtAVze/20THgLAHM40Jw3ocNC+IKOhaIJ2XTMKPqW/kk9gFaHUzVSJDk87wh1g+/g
S9Mck0P1Yw/S/JYthQ08q7LZqjG5HAVjtvJHmVy/4tzhB8cBpDT+Af1guuKJq124zY8LNksHxL3B
5RzkEkYEEo/XjXuvOdaLyhePwHKRvy+vnFl/yB1zL290zHxLvIRWCl+gqSvM+pjCKp4QJ2UinA0J
Lzqct6MegiSjtYejxuZ05pX3YuAuaO2nyT/GE+rgaaRht3RIdAhFnDemdExzqPJLzZ0HbUdI8GMP
HGhggMXLNhEyXQUIPq+IgDoB2o9Blh9ict41+G3DtiNyLK19Yv5Xw/VA1Y8+lmVFsPtg78dKLt1R
p0nBJKr+U1ltbISKdAjTh/8iitI8k0EWvwE+Jr7qiAVjbcBeIZTwcYRqDV3IamR3v+fvM9Dr2tLa
Jyf8MUa5hFXQK27Tc+lTFaEtbR6Wh2DrXRDfXWbX6kkgqsevLolymIxwx1fX+9l7nlO5uagYi/ws
dJoBL8+YZRmEi+OvQspT+MkfVApn3AMJk9o2l3cCzhP09buzqwBQ/OBkWE07A8VxY++qkuGbzoQq
byXZ61VFDXq3/6ppjgDNKFV1+gxFsMc9NenuUjxr5B9HCvw8V+oJSDXqwZPa63OWVZ7XIzkPSBaB
ulPLuQziMoa5TeMWZoPkL80yC6Lpxw/nEZ8u0rOo0aMKhB8AZyDOrG5lsbeEaaObnaPtr+4p03e4
7W4Z7DLjYgjEtzsZSPO7Nl8npJhBmVNggUgv0OiG4k3Nve4fphnkiVNe+vkXgwXwVKWjTQyyEMwb
M9R0npqcKd6uBbrV1wA96Kul9gvE6mEbcwBT5/OMwRUAxhAxXTf22preSv4HlJquShzzGge7wDBH
qAYoaB72DK7R7NLGvfvZveC0uqJklpSYMpklbSi/lBk2u8/5WQ8d+2HrjQ7LRKvPat9GzdhdezOM
pBBujkAUdJlc+PkD67C5W2zxnUVfQv+sDOCq1Bd5b56xfOj9LcpBA4B+c2hhQsde8hgpHksCAsU9
y9criy1ku510BFqiw0RwHBOB7Y5PszulSy7Ju1rXk1WAHqTL21OODyHBesWu5txPX/QIsSM10/4A
avno0SkjyNKML5bYcqU97s8FOdG8JIg+b7nThf83g5boGv+p1zNABlAY0tV2iO4jbQ6GmYvS8rfs
uL4kWX3wKjLZCYgqO9n5K9RzB2tUwsdbIeECoSsTNHD9W8+lr8UHQzrcOsCOTLQj1V5nbq4DNXVd
Ke4KrnkDFxqd/U89X2yLuB3XRF5+fsKkR3/otEvho/ff6L7C6yseky/fID6ayeoKr+4xCK68ELrA
mIPDWkJx8zKK03Mjy84UWJGRvZnRU//O71HsWQbQIna/weWepBOUgLnM0BbKKCg7iMagDVulqACA
cmL4AwOyKIeEtqZigdos3An1BAxaUYN8elbbHGacWLoYG1ktqB7rJk/daCFVciRjnUHnw6ZivqZA
KyxuNDE1NiOCeEXHEtOP1XtOvKJJ61FS4QvGEZ5v/xkJer+NV6m0BP7OJueejQYL9QAob7v9HJDm
/23t+8nLFG4PujjxNwVlzW43p1xJbFsdLN2yjYyul9VpDdjUrx6Jk08nS1AovyariNCk5qXDfUvA
kJHnuu3UWadPIPQcMPYfVj50+cKfMFmkzKxqcTgkZQoDKrOfPSS7Zgg8orgh8f0Bw6vI7ckoFeWz
LZbGaCOJ2A61fSwCP+35XHdhUaMvdLgFJaolaEqhRvAcIjURhWHElMUsGnCzrHSy4r/kjA/blxXd
D/K7W+HmxXxX+lcsOrC4hval22zMQ6egMvaoE3VqPaEfxZ123jD+6sSBTvfcc8UFB0kMsWPnkUJy
c4EeYEDzUjOaxEgYvPQ8YY3Q2SKVs807lNVmoobCHk/FQFjBVVEuPjiO7R5EoJEfpgWwN+HjuGEG
3z28CFPH+ToSq+hOmNpg53N/fQRiXCaDS4tsZWoD7Lgb3iJElF+x+Kd8ffMHdA1Bjt8VKjs/IZyv
pB01jNX48JRqxBhkAEtJjuuB6MX0BFgsDEmMqT0m53evWnMfrvlRYtbRXqX3LjvEPVP06Cg1Ys0Q
8u2rPjOzGZhxgdMnXb1FMtXiuXfdK2Nm3JWWa9/BqK78OUZanQ9mQnDoQG9WGfpe/QWA+4WlEJhG
R026FhLLzUq/oW7xlKnBlvW8I7rYEhlM3PdxCK7GDuIB0YgAhwGyAQIyer1zKUZ8JZuYVyG/blX/
2T78z47gHhX++RvJB6iaO1EuoaXuzaJrYdvYsNfQywJGLLhwxwFn3cDiXnGuULtgpGPeQOtai/io
Cmd/dcgq5mO1mcJ6mAAUePwbmrwQh8e+/6VEKxBROxyglL12IVIKYJPrEecPR29t2LwbtADlFLYe
mPE8V92uvZBG7kx+GwEjj+1qEwh4PWp7WIMrNnFzkdxneY3w2fCxZSCkzJC7VywgPTEi18BPtAED
1XqyHM2dWEBBBSwJzzvK86HxunrEEfvoGVPKphwNYFKHN6tioNfo19zYi/QpmYSGTeOGN7ak3Tkc
GjAmg7BWZR2q1VPrtSo8waK7qQgb7SX9OZMxTjeFogICA4S+VKEGevYaH74Fq749dVFpNaRFBfsf
eIAC27hCLJeerbqPy08G2w7kCvAg1LSO6UmL2ZbpLYPyhMAtARXPdv4/3BgSZ+3zpeadH5ukEDRA
ez0FMbMaHP88gOxTMAuCYEdxbEq4qxdXC5uathaGDkxyubk817TMDNnNqwfye6eprnqadaFPmKQb
Zog2UZ1RRJS+f5K8SrRkC84I5mdH2TFEAtYxkCFcXQ+cgrXGLWDMiusbqAHkCp1umSg0RT+GtiTC
x94YOOUOcAQ7mMgsI4bwsSB8jUYL9sqW0V6hskYKvLNqsCvPuHdFEO4hSEfRjvU+MRT0cOf1mcYu
6PQnOHE4yalA+A4iwTwBj1jJPDOmw+PTril1SKpYIOMUngLkrsGi5I8075ijyIMEyFHdUUc+Yphj
JxrByriyUui1760TL38/YliXHhG561p9uJC/GQNRWv38IdDOxKdbmpkhinLBuqURaBuSTUUDWPLq
lP1LdUqkXD6RDzwhmTzw45G8Jm8puPZ9W6OnoC1EVS200UImtYExLmW/TNqbsE93/vN4E08HFSTD
1pxuGzR+TPCVW+LEqZ7X+3yZkmX32GsPLAvnEk4LrTB5oIdXgoCXJrmbRssQ3KbIWRtrjfuDBgvj
3EQ6XIMIhkNkvFJE8eDgK5AoHpIsET8czQ6irTg1OecY0EJPZ+0KrLt1uRdwQHOgevxd4nLoOfVV
X0uL0JzLHkibPmd8BoMNPs8vX0XnhT6cuZZz3wY2BHQj3Awyvk/Mev8BJ0DaMUFk4sG1rAbRO4fC
4d6hokQfDp6hDhI5qjjLAbYdCbY0QBhpIGLymTS4AAKjoOy0SKYd8vk0h/9ZyyI3u3XjtzrABAVy
HM6LFHcxfUGTL9k0GiMnxQjb3+Se0+wfsXgHnBsycd35VRvoJ2hY5Hie8Gp3spcq20ngOiRwhMQ5
bg0mXpX4YZSDlZuK0xqbI75doR98C2gRepKo0W7SaCq7bYZLwMItckWDW5KxkN1VLyWIDJ8Ih3EN
ZB3cM5Aog+NO1sLgo7hku9PL3UYq6V2nLutC8iJ1DFlMJhP0DX8/oqzWJd7WV/+WV6iL8XVtao30
LYab0uSloGGAQqffz8cEnh6+wtjvHIhFTfAFoYCF/FI6/pDWfXTCTFf9fYN9kF+HZN06g728P0Pb
ZBB+tqHYQBBLjFYFj4QxjxVrP4tMc5M2CDU2GhRgjVLa6EvqU5UZXDRN/irFi5p9uVHfrKUykant
16edgaWHR9LbtaG0LprpjdnpKSCWCyuFsXQicqJT0TFtgpXn3VmJoFgTaw4BwqXoK24yy7n93Gz3
4YY0wxtt6Z1OPhOji8TTDvp/2pcdzIf2fqKOAemZ5Eu0nvfcbPV85ZqZZ9zIKberekDlZ7keZ9Tk
K9Yqb4/2wnw3UPqPmAYllQSjwpG7wLd+4ddna+kl+G6CmoQrzAxe3lvRaslHz1iWbCi4Svu5I/oO
isRD3N6gn882/Y4lc70QdWNYAcbZ+xvwevqeVfGD5EkY/Ltw9JdtuIKLk2mbcvcPuBTMxif2ywxr
YWgtQZ3iSwBLKgkDmlSeqwlGGhWqAZ5UAq4PicR4rD5slWecy+a1iZs+PU3G43/5XcpvmFgIrZSf
FLVOeOyxFhmrGFH16OfBaxxI2cYjizrnxfQ8R4Aoe5RYpCgdvGVXvmpRwjcS0fhNcGaXwnSR8GYy
dyqwJxyJQ+2HEhvk8eIdHjWKznccNXCdk4O5qyXjDHIKV7zaYFd8we9rQQCtWPSHSycQR22JfhD/
h8iWnhCAAgNV15/GjGzJW3ZBJaKWbwm5fSdEvzqttI4OUMjFvrkMIHOVGKa4kr8lUADb7q6y/KaH
L4hMJDIiH2pFdjMpXIJTVnlQ/0O0Zj3fMR+ndO1744CM2q2GjR7EygxZUV74kaCd2hYnG4LipQIf
alcuKyu5Q0o8d/8KKkJ/3fe2SKJmpDy74x56SAL2wsQqMRtWA4lv6dniI+tB8SF4e6lJK/GgryZv
bRSjB0khbVMrBHF8mf9HkGOwGqFrljQGj49Y7QZm22kGj2/K34KaOSpFEJ0IkmfC78LtZGbBBMVP
6EIxNMeqj7Boo5dWQfQbCAxqnN6FCr/lSzBfUW1ZXJYSy49QmBtt789UiU6PnbqbNqyVDJTg7Zxh
DUwYCR3BeRjit4I2ixKDTqqHUsgQOWfnP7DaVeV+onXoynMR6ToVqdgB+LRfOCdeETKy1S0s9Lc1
XtQdjVLnYaRsgmney8+rYrRoaD+8/JHv7JpSrdCQJCZ0lUJ6quU+xd7kdNhfR8Eqfk4zhUC9/FfW
DpnxJv0/4FOvRynHSWrrG36rQVWxS8d8eGzAMqkzNUF8nTfsbTnI3KUftwir0rP/QHimcQC3C9e6
02VMo7kz8IfFqAajTBgS2zljUcVDQKosu8N2q2qzxTbC8ICpUNi/3Fb9u5YCaI4ksrATs7c/OgsE
P1AH7fdrgvRwICWfLa/NfeGPVDZq3tIS1lg7jhbNrVkngTcgWz/XC+BQIIqbE8mp9UtyCd0aHmuo
SOCJ0frptGJuPE4E3DHV4eM25eqFW1k1Mw5lJVfZyKWoRe6oicVeR2m0NTeg4/0AR73lxTOxhYWT
RGGnJDtHCsx1iMtjGhPraPyoqordCKiAheCLtqYbC33zdt9hdbZ7Bgwtvw9uybOu6Y5zo3q5NPky
o4GaUgU0EBIpm0N/BjMTbnsoiWvWSI1FLOs5ApD/emcCC8bsMazc+9BO6DQKWkqWl4MmE7rb/Otx
wt1E+Gzo9StkwTA85lbw/m7t4MQgH1gBP5dxFKTDseKk5HrkFqsdPSjt1gGNpJRjUHmLBB8EgCVC
/+cIHCG2GzLl6TIonbDHCQV1kdySChbYnYbrlnwOMigl7mpGa86pXt0UK7xqDewEJKIfGVtxYqCz
TInFZMJmLI4sR3mI5oweiqsyxnh+BNDC/OrY23filpd3eAENVWw1rWy8nOuQj6jZLN4GjGDq3tWZ
D0hIIk3pG5PVvtMaanS7f+4PD/vyJS4Zd1bHb8FjJJ1wpZ/qHmicBMR4TOnHATvG96v1LXl9zMaz
jeo4TM0pElSwFXJEnn8+zq9Pt88TPMOHummKEPvuVrpDWUfP02l5cpfVtF4TwqIbJWr7cVq2x0PM
FIypFF6uM84sFLJZaz0SACtWpBrqr7CFYSgORtVhM+155k1Cg0cb5Km337LdRdSDT+3vYh2zbOi1
C6Mdt8ac7SuKFUZbyVqJIhrrx/yMODAMpRzgW4fZwwqvLhaKC+dygoKX6+IS8dHA7hFwPf8tX70C
+B02K57eIZ8RnYsgwny5i0XiggbgXobyG5slyAwtgWZnsPT6z5zx4dJ03NyWDgwdkeFBnfjLApwp
jTYZ17B5Ra/U4CQKM7Rge1UmzYfX9+9fuqmd9gTcsEn9wPP4DHPDU86D/gF+b4T5iFVNc3UZmUFO
SIKtrgcKpmStx0KnmLjapc2gO5RB/YLa47AEw5+W1+ct0GabrNQi5wdDnurw2mWzii9+LO9kKp2e
zNPkbM0ntm5LJ6z6+sKG/z1t656keiPkPVpezVA+RCgx1PAXHsn90yjizvK8qfxM7H8zfO++ap6f
QfATWBHM+fszmHKHHdxle+cTwAPRC/b5vjVUiWMV5jsjucoM3AQ936/mhpSeAQjKfF1HSWaSi8v/
6O4dIoWLvPhAcHE+cO2m87nqRW68VRVK8QRoRFka+CInUwSCPB3A+1yUijGXpU6PJT30w+cCEjgh
DzAtSuu62eVXJuHHExq9+Ccd8TmIuf16Zmq0Gdd2dOWgLHCwxSXVk0Zm0RFqXFeEnH1PsO4tHjoS
c1PYLTw7zjXsdd0VmpfzxuNPgXzo+AL+DGtRSfXlvEjqQbIxEI91ij/gnJTV+/bxN8BP15EdldOg
bWzOpSpsFxxajLMhIaTY+kUYsb5vzM3XOitqziJvx0rUQjqFaVejz+3qTGXSFUsQLGdIun72CqHJ
OhlmzXab3bDhGpdQ2DtPspxLpR1+xWK+xhyn7LHWC3fmJe2gvIW2/ieHodaaaHTppjv/sAeizqTs
+to2RW1v6NO/yeE/hfE8j27cqCTXk2Dy7SkxRP5TSfv70Rx+Ny/yN9TUVCuczVdmdPst9oWQ9758
trniXf2g9/QIvBSl9Dz6/lFAoqRWaNdHmKggMYdfLr/+3C8BYJaVzYc7+x8dqDDZBPLRq86FUlEh
vg9/ZG1T6t26nL9Fm6lIjmTayMtHXq9N/B0VODVEhp3ByNY67r5dnXrCCN1PntS7gH3qqhdrFHIp
lEgZML2Y8AJJOqSBqPSGmXcukLIE4HiUhM2hHtR5T/xaqxyes3G+ZYroYmB4yji5TvLFLWgYhMK6
A8R/0mOviwcyn2yQ3GJGc9k+EDtZHxQ3AFlqGmzDR+hAtAkmVmjO4eu6UM6cJuXs6lx10GghjXkh
Y2hTrHjT/g9gEyw698E6mgDNCmecV07lR8aNJ3V+MkoX5w/Mk6Zfq8CWxSg8MMOiVykiM+UHAlny
ylA71KPOEEo0XjXo4KKZpVGo8SvELQDSgjGux5alN1bHZWfEPOtYohW0P+/JJXdqwlx5n4hE4bl9
wxcKIBSQoRWLSuRg22TXa0cYVLfxXkbP6kkgsHCdwLgreQMyGRTnPEG261Y+WSmx+VvqQH94pCe5
eh6RjrNvh2xuj4qHG4jQXTbQihhWQlhyUq532+aP8Qgsmf6bVv9aYZLmmSU6Z81bwDCcxbd0UtDu
QXiCtCjFnB80idlv7qZsL6VNhBm98Yktz0zHviHhSCxvUArD03i8hOaQgJXqXi4wIF2YnvgPWKev
Sd48PIOMAEe9GMU94pXxyae/TNDozifxae5jh6iYlYhPZP5JJi3cnmMvbW5KgnI1IqJmkUHiNOBp
UvPvvjKMDwmx4HOyUJDS9S9UWJjygBXaKRsuh05Sy9dYssQKzv32yj6muG/LMziQauYSbAUWcdPR
l7IBsoHXQHSX1tXhBva+nyl0cdF5czB5oAxVoMnRqBryVaFvdRl0avDhJYfetxLUWkthIDvDwKMI
e3YeXp7YfmjAHuK2QLAVYhMqPIOZs6ulW0x1MNUvYWb88mUUIvX9Qk3dEl9WI+ACnH/rLKcYLvQt
xnE57wl1xNIfyzJIi6klX3bIT9ricPwPv00cHsY10EOZm3yfp0pjFx8olYVQPaMraqUfAbyrigB2
2BGh5m9+kPVRrTuQKwH63GxrlqTqQ3h1oM0P5RsUPf255YpsutBrKBH04LO/5Xw9UWKiKX4v4tx9
cFueo1PNUcyAKON4+LJPA+mewYCshoGPZZqNaLyQuN6RVm7YTqFTIYoMqKJollkFQfIgqZTLR1cT
o0YWcWkPosfdzH1/xd4zx3/iaPaSRGNIKnuve/mniePKyKs9ILNmEaik7PD5tbZ+F+Gw7tkpMehK
hjEKuKD5PaGK34EyUhtO1cRL6NiIZOoTwQPx6i3f99kTKYFySd22BzdGZr1Wz9v6e/poDnYcqmRk
iOWZnuMrQjXb8+lT1VCw8rHDHWrkk28g89m1EsRmV0dlaTsPyGXrIny/HQ+4Sn/EBiunnCgM4OT/
F99gZxrAX71E0gnljDUqw/w9qC+TqbkUuMlJycjLa3E0yrTlu1QfvVJSNzQVAW6tFbuyawaflVU5
rsqZ/Y2IypbeLjzVy9DZo3S7QnoNnnhXgGLLLLGnmVXCuGo4GguaNTYepkMR4wUGz3yKeTgC5SKQ
h8V0SCaNfxAmY/1Ep1fq9XJ6geqxVprFxE7GY0+GwZly296X82GInnHyFtksupf77jgYQ3zl58F5
NDnL+L2zeESylLL24r5kd9CS0a0sdL+o2pQV4PIR0I/4e7RjxSbUp5P3sPnzcvsH4ZnxtSy5HRJq
668CfFSdmg9/DiWJbsZiIJTAyjhzCMq5PHYhmRITRBsr9JCo0mMRFZNV/IAkZWkZHQy2EivqvLwr
YA5GurjLVjfFy1fwVzuLcKjoK7g+sB6pukfnFgpgiVobdWQIFoYMkN70GctoPic/qxyCz62frZ7k
D8CaIIcEcwZ2nrPI3MO9jS5YkZN6UbqWHVX4EyWKAu6g5oQ7lYERHZfXhZdRwR6RKYZ71t4xUwJl
mxZjggHng3NP//ZEGl1rsEJRBZJZwrWvWWoVZBrXLAsZZ8T5jMDHeKNNj/zZfgQbs4cchIIviFrm
mcTRhyGDRRjgXwLYOUA1QRea7cpFMFioJaIJaaJB9Hllv7yWmCufiZVe1y3nj1mypUwsAI5r0OK0
cLpUGMhF4kiAtJSJpzL7eDafcIQO8r3M/v1Eh/ssAga+S2LiXUlHUll8ehDnK0SvJKf3L/8PC2h1
UcBu82UvMlaEbNeB26CXnbwsX56TIP/1D7/ldezT+mKT3pyHB2i8t2mYZXtxwhgCPnQ2QNTn69YL
7UXMl5v/lFgXXTLymEpK5Ctd+6UXaR2A8btNxJh6xLMOnQ0u6mgyZFJqmOcAKo8a2TSYou3bNe5P
BJnFUoSWRtWTn3a/Cj5PhnhNVO4ChomZ2ptPDZsH0FSIWRgJYztB0/EBw/V756v97o/mzon2HJ/W
V+Xdved+WSdZEjHZ4wew9ZQrlf4ZLs/SGLXRpSNA+5Mu2ubgupjGwTvdz1zf8k2ainlKEr6IC0le
AwgVntwCS1SwpqJjdHoBvvJoRCVx7tY2xLdyYC7qsNX7DWA5JElxSOu1Nhj9q65cBlZpC9v0vIzH
EAqAYosMODnmVmkJ1jxDH1+8K4+Shq6OqAeBEZnneqyaaTOEWxAQ3Rhg9tmoiEr5jsDvYbKfnox6
RJX+42eHpwoNXSWGehL0eJkPS00SAK/J82B5iPnqNPjCEQ8BRTPXONO6Dpy0mQfcL14RqkIzoabk
KCJU9l2KYHQ+hm1mp9AC7NoRO88bFSxdrp19K35LMfyq0/FXe7WmoTJ1+TUyrKQ94lr+PU63E8j6
y8QrUQb87TuzNqlV05n6sGBgyxpVjkyRSmr4wa9dPypL1DbrLYc4urasrlG/4Qc/w26hM9pFr7On
7FuqvWcmDpM7mt1Rz8RjgwL5cZNiUVnjCLylpeLlut9pX/skVpeoW1NnjMU709vaByfusRR9Aw8z
ujz+RT+xuJfF015ThHnVPWLebWRgMF2+QR32OhTQ7nvJbn43Y5nPvgtkT3D105/Txnq7EF3V7X/o
4BNdRl+zFQ3C/ZqkmnhXBAmNIdZ0hMRC21Ky6auzuT4+tzgME5fB1AiNuISznQHwBaova1dcWt3C
O7cQavJ2bnP7pCIYy5lRqmET+FlWflB7UYfk+jaVMsq4p2oKp3eNrzi6OyAU1RaNtiCaVO5XdNgY
/7Ew0cd4AmfMJFuR6E7eEeBR0TF59APILbrlnny0xOnYdwNmNBDWQsG6IZARJiMmc1EO3bumDo+d
f4F6kkheMiWpPjSOLS59O5ehprLKniZNmuIJXipqgkTt6JuULk/IsPXZLuuR/m3S9V700Skck6HA
1795lEONkdGNsRTDOQs+ALgq9ZyKmds5NPuF9ffDC4Lt0lWwXUwPkPyuXfJfa6IHdOCF+X10JGUr
CwQY5U4ctrxD/e86yDU2k3/Cx9gDQ/DrFnen+tEhxA7X2Dc5wkBbqGC8albfPbNxdeJoJQWT1EBw
+f8/zPAcPe87bK31lQm3H9BaNMHqRiDi1i8VCNp+GWEGBb74b4vYmNdkZ30LLdcu7l5cWa7ldxxe
jXrGuAp/zMGWm9euiihxm3ey/gKOULoc7t4capTs5MtcreO6MRtjN3hHfznSj9Lmvmj3yreEpZTD
gx0feNkSLpvf4Jx+IEiipDZfTDs2U9lAzo18zIVgEgkA+4DqZg+YIcRod4wOExEaqkQWLV/qX+4Z
zZj281zd92daNvbqLGkEZ4mb9bb+yz1DcB+QIyfnvaEgTqN8w0p/kZizYjiWhjyRuV87GfWpiRq3
DjUkKVwHYW7b4qc2eFJDWO/Ug58CtFKT6/gD7DlYknBHzwnbSe38LNbpgtLEazFDhweELZ/HFq4q
doOvXiWQJ+q0Gqxh1dG18oEUJAoID0D42nYvgsLJVjZm/JKl6V/rHJR9GrBokGTzuotzSF6nKSG7
3u06T2d7VGWTQAFRzrkEickIJKgLR4jUwJKO44FCSmE+Nak5JWH63ppYJ6yRVY+oasVmEgnHFroG
8PwxRUZKJm6p2MD38vQaYKCoxVF+eXph8y9shsfhspPb+0vOm027VZjFD9rppjD7aagtIgzeUQcf
2SIkLNn1eeZ+J9FQpw3WHftTtti4Sscg0qTU2YK4ai3z06VaFqinYtq3wLg9ExtOFFvPEfPFffMV
FhNydEBtCOlHJeyjcQE6wuwfFAtwKHDVLwasmrUcN3eRT7L6WeVUczx+40kQFphO80kjDvHzJQdj
2cWg3S9I/xuLJjmvSmEuZ6IRDZyOwelcMF+adeMin6ghcWVq+zM4Gez43fIZU5bQ3kENumZjYDMs
Tz0VR+JCLSRUz0yTxu7R8Rgoix6hcC5iZ7+1lqurr2KPsT2AFbKEoEfdpfvbvghVLFBhePop+q8q
tTtnVuqUt1UVpFmT7M6M6OlDYQ4x1a6r5Hjj/fYqdUIOpRPrFeak4bUJj++eAge65oVnqr83eRLn
fxrEa67S3kVBy4T5vin2Y2bOKJc+Jy5XNUZE6dTWlS6OKh6f+YE+SE9GekNugNlfTZD6V4G9OwoD
D5180GgMFeHhxxQeHe7Siz5vdXwYjlfElblNHrn/9pOxqK6uFNAzYEwg36rNHZ4I6BvF+0dTTgYj
g/TGsq8sTqldHDSOYY/06Aug70pQQj3rpakoMhTTasxS/ZQOpuEKRuTi9zA00XTP3Y/2jJst4nCq
2+2tddqfTvprkMYvfZa6erGPFq8kqgWP5WAvbjMKZrmkAR4bggsXUyZzRyv9f2YZ3Cu2o3AjXmPR
9XKo7UEuwSRc3uIAsfZLFSOLH18ACjwCK8mLwQkq//Yjp4aeoCYUQAIY3mHLKX5wy0ZXmgXcc1uK
JNS7IdIY9NJKyJ8Br5Yi9HQmqIyEuKNDlJhrWxX4rfwpW/cL7/x0+sFGhrAVQcBzc5S96sKCSg1K
rveoiqrHKm3BK3jaNGkWzDJfb+xQSBafhztwwgMLVEeUxB0RnIks20BG5OVZkIRAXloTfqblpfzu
j+b3uYtnx7NIo1UFNs1qyl0m98YrBQ6LpTUZRruiO3nkHJzleEdQ2oAgb3QHg+I/GFYfprRsqlRM
fxZoM2fB21i0Q+37YRNvf04rRWzT4ydELN50bxK0tphtqxuk4qp0/2OrUB0vfwJJZsYTGP2g9Wib
boyo7efYRHvzahwES3X0wWJGBbGUsqW34274TgkgCvHDtQML4R6lv6v2FFuQPKzW6U4iNadEBkLn
9kLzrlk5ofTnSSZIhGPJwgX5mtwbyOwB0QliRRRai1MYcWudTlu2gbx3ir2wHWQc+goMVc5thmcu
aOvX6dqBY9hK4hEMm508QUCGHLicGcMNRLo7vCf7n/7lxKugaQXGyvt0lcGgIfjZa22sW/fklYJg
XJqi8wRFefQOE7tvKpqR4zRqInNqMnPV+vbS76TOm1JUUNAOD+056U5tIG6JfIKyA1tfGgVRoinU
gZZHGE+inY4ZbUvbuQ7EdpB4kTXC6cQh59IAJAZMR07/pj/uN+9e75ol2SaNjhTCEiDNmH8X3+O3
YgnG5ZHLu6Jofd9/jiCepLP/Ue6yUDQq7Ys3vhvuPs9NK0kL7tm3FZi1g7y9d7qP2sYZqajKbnrX
Tc/MQWvOy2p6CuMWpwGuhA1P00lj3D6T2CzjJYjDV5gjS2oOEnPh6e+UNmA5hk/l9eNlLAc3yNfl
Y+K+Q93y/7APis+aMixCumBB8ivmz47T02eDFAJKftRrvBe6mhQk41f88R1YqhA867k0vsuUXq+M
0YoIRkLjpPXv+dnRaBi6+dRXSUkT1h3duRwWfcC2oYLN/pyYokpGmuvd8Qa1n1JTCZClbTWVFka8
AG1GKgDbi0QNQ25bqEDwqukZyTyGz+ZoSSEs+shvAV7VMKmi+fxMNTZz8Y/WXYqVl2hs2vxkaAQc
7aQF/Dq4k3pdtqRvJnSXD0jCjVjf9tm/SI+mVIxe2ig1LPYeo+ucr6W/WnymeK2Xp26Xxaz4LnIq
hDnftv1uTFRNXP4ly/dpBhUw0AQ6nUAqDBqZ+RR1ieYS0lRy5lSMpSk9Bt3wTWhL+hUxy2bAzPvx
pTB1eJVxg4jGjkOsvd2dPxIHKnNpEpvuc4s8Wo3zabWFY/d8sQhX0EdR5p+LDSwkHtMJadFYlunW
czt5DLcBdk+M00C0vAi5DFFI0K3ZBsj1pNJcLku9RrZ9qNMUSyCVREkFDNaTqlFj7DZm2btzi15p
9Ubka+PavCs0vHdaSGgAQioiRRzXixgjWqTXVvot7PefpUczwcmdFjaCojEzs1958Zoae5WMmyLi
0K0r6DAH3AMvRwhtnFnksfz+VWix3jRoU3DPOieNW2LVh1A/OX3SmAwhfpfLHX0SlVoe12CQNRKS
AJR9F85rhGWYwfGUjvmBqGkldnT311iVs//FlCAX8WGp04AHnYKsuw8mpbmgftbsjyxd9FClDXfs
FcYRh1nX316ewxtH/yCi05fcpsuT512p+spA6vUz3PSlSV0293mXztwxf+hY02/hIa2R9QGb7Tno
KqySzS1JT6tKk9MF6iAU1IgOJZTGhpDXguH+HmAlFE2PCvfd2TYHPe7Wi9GyCsB+FD9AiLfVv4Sx
r6ODl2M719NCV4Louhy5CRevwajeTFizlmTm02CvJsxZOyQbqhY4l8/cpusGt1AG3t4xC3wsbm7d
WF+xtq3/CBRRdgTh71LPLjOGTrxjh8etXPrbHOqCvx/j5JBzCzUnjeEvqSwTEy5m9SeE5F67NOOn
x/Crk/ijLN0DGgVqzUpx0gWdcBJ4LFVLukjHCqkJ9dkL95E3klMhwsnMI4ZEYEEwkzrATM8kyX7f
4XAmeOEbTLaGQXrP510nvcqykWg8BFO6ub28bdPNHtURGv6+T9SHv3guErQ7L9qeYPsaL28sZ6JT
q0/myTq1dRfcTxDT+x7Dxmyhqc997pgBMMnNU1NdJq34FYlYnURmtBjL7j6+HS2yeQ25HnxYX2j6
JOXAS/Rk60lJMBXtuP3RZ9bh+K17lpDarQuJqnZOLZZLJrckugDgIXUrOMMJ2PGi3CQ/QPNm16/Q
K0c5E74tjBWDsO04LX//yjE7gONDrVayGhvrIhOHyppcku/HlSPceV7G5EyH0WwnNQZXTHiGhU7N
2EfzIkhf7rVdj6CtSRUJ2gjE8byIM0uVESDMS4cm5+nNjjN5Rf91fywK0/4pSi4ufOvkbKSKf4oR
drN1Gou5+6En2tTOLAG+iGHBFvLdg1CcpH1Yzk8wo+AnvY/6I6GxA+qfe8J6nJox0RMastzq64It
UlSLlC3bhP8viqeW6wYqoV+K/Ml2JS5jH0DzsCY0uqnI3D0C9o1tK+MvSFFuuaB7kFfm+D/MIlDn
E5wrc2ev5RYqmTZcEFezRVvLhvxAsfWFa9g4soUFkNeqqys5PicYCNKj7tSQFQAhAoeiB1Ziv7Hv
kMaIRxDsL/YU7MHriT96wd9P+JUXMUGqCo5jquP/O1m7uFtdzrn3z5E3tQNVjXL4A8XrZY5beewj
nFNoq1g2B0okXjvuOv5zdpUgCW7GwV4UZnE6z6vHEAfqgVo8z8YIw6DaMZWfA9g4A7DvQmAc3dxl
FhEjH99CmdOsDGc7z5SX7ZRKFnr0Kik3HL3k2WtqDc5PlVeMK0wi19TKezR1LPnD3JMM4XreGRKU
9B/sF4IoE6lVyoarUyGlsV9jMc1qmdSzh2P4sSMtA/eQOPv4XeMa4WrL2jnIYD/qyZofB7nIEM42
JNXeT/AXIyBiYv/Xwv3auXwVO/EsXhwI6JW8uJmOeCkXKJg0ed2h9Oc9Ff1cIuOc2XrdcMgq2gRc
WLnAePzm0CtWDlsD8r60vEZpQMXa3xFzQYBMkIh8RIV+/jSJUM8Y7A2W6KWUub6t+e0ObLh47Y6V
GCVhhgqUnzHz67DoXWp3yE0km7R0o6l3YTmsgUr2WpK84o03mPoXW1icViUsQ8ZaYvi2DdgYcBlk
1twtgeKPNvYy9iCmIe4zw15mf8bofjYYIZG0VWCbcSvRvojlZVJ3/MkFwN3OhalygbhQfR+fU2BT
3PFbBsSHPxMzkM9LHUqW5z8Kq2QvLi1lhs4/LLptFjkGXyxPDJVJX931fv+N4+EhvkyFjOi9LYgS
rZGp9hleIk2yOPy38yjakUhD/nE74bpOjtsbmSRZMfH7Uupy+KbC4nNaqOjtNKOD3qLeSfxMPf/9
luzt1ahQMm0HCPSqkb5KnryC6M1vNBH6kM75K2q96uVSLo46gf9gnE2u5D3w6OOpoLdbxdStiQTr
MCMMSUPH9sIUUBon2yNj90gxb+ScN6XZrLvC8NBqVEGBFW9FQp8SsuF/s9bB4RSZe+lJQ0CouDgQ
n35DQRBnC1606ifKuCGAhhn6cUF55EPioaAisQ/oLW4rxWmoindVd3JoGBG1Zr9qfjgdczFlSMLN
MOQXaonVDuw61/4R+g+WQ5vpkYWgTho8x8zclrVvWDlDRQ65/pR2PAZ9u2+QJxUOj9lnU5eBWFLC
JjXp5qkyVYVVj41T96xSRrk8Ftu2QCqD/ka9UyVbIBPclMEDVodiegBrFFHy7nzbypSFfR2Ndb8B
vbvxTAdPdSA5scznLTflj07HC3Si1TWI7X8g4qyLPND2xjOgavCWngp4RJRLEQppEQZIrRP3En2q
g1Fr1iTRZiv4v7RLp/bvNrFlZrDGfA6OoYWMoragVO1SN7sMtHKR8rz/IPDqnkOqsSt5+TkOc6um
U0DqWMYLTSlinnXrFIiuhqA73XodEVXAz7IGp4rZQE32yTW5xBGscA+HfifpH/ufSt1oMWBdTrcA
WaiaaRSF5r4/3VAbNUf7/lPSROlIgq666ml8qZk/nM01eFUPGRTt8+QKGQo+0bSdtUQBHomYsKs/
9x9urB1bxgfpJY/yOzi3IrzjBzyGcbBQXfzzSVRdjlnLTnQinjNfgN15uRY9zliUo+GWTQ5k/pTJ
PvjTN267bDuFcqAAwTrViij4msAGCRfIz/fosRdLIb3trKQRQigVHRgbwEsWW0lCQ8MJS1t8Gmu2
1cXFrNTmFkayN9HsgLHsiDBcFHh2sx0tuF6tCysjscuvPwRZ2nTDn6hQVjtVEgRguT1ExAenM2zi
T3Aov6BXPTFMVRqj4vNsIudgY/hGpztKCA55s/twaCSy/6EiC2W2ZovZMjWQWnhQaIA3zLB2tuFQ
q5pYh1i90DUIJli7qVpVJmtkCFboCV8yFRJQasCri1Mv1pEy2DU9uLbz5lJOZKeSDGtLkRs9GIic
iefpciNcaXJxAhk/ml3e7TnxK2oDa9ZDypiW+o7zEdJfDPrPx/YuaYENkF/n/LSZixuk8ir1ABbY
M0YqjXQoiQXzvTv5r1ioEZ91wY9jIhsNOjby6egpBAzcMII1IYaeKN2sdqM+kbbEfYBAhghx8f/l
H/Z/EaKPzWO5EhZpMCuD4w4KD04Gw0IGr9a/Etsm6Wi/yyYIHN+aYICdxqo87MHmQJ20k2GAS3MZ
1ZmdWrEbTZtfmh5uHGl6FiPJO7WqOLtWxvolBaBxQdJ8YASlg3dhMWcOXLVktQ+2vaxNsnWczWXM
cEyY/pdB+C8ub1Y0U20kunSn4eZ5yrn01uYG0LiwM8xBQCZmlK6B7XQ/98oPJxzBJDj3wI9aoRB7
BaJmnHJc1QH9DWe9GH70/2qr+SWJwtVeO3BfOR94do/iBU23+9NQbeL9F2BK8zych0k9WvEF2x85
ydn39SRBQwRb1Ovxs6eP+gO+Vzsd4/fcBSPzIAOYonOlmkNoLCy9/KF4QL3W3rKcJKXAZQgVaYMU
b4vsM9jh72cYcTwK6KuxwOPL0iOoqSDL6GFxxNq200jDGBRh8zrg6jlINnRJgrcAZdDOhmILmVz/
oYRVIQhaunFFbunOeHOcX/9uY6+ZnyJ3M0yegAwWiNgZELHRzMOM6LEeLewIfc3GLp0s40P6LzSS
pqr8vC7nG+rxDqLnDXk6qgOOQySUFx59jvrV6FcAkeRqlM4+1Ocm57an3FyywDHDWBRjEF5wrLDz
BhZNCk5ugKqcluYRyQjubIK7nIacA9K064TwHbcXDZauuu0KndtHeiuXocZTZBsd1DtNyGeCCyzI
52OAs1hNSHeeqKRKtk4SsoXwD9tFDCsZMxCGSa7jFOTvQ4RLwBvqkvwctZRLi/5jXf8jaF8pJ8g5
sPL6zix2h0s5l7Gc2R90BXcCQeLalTuYftCeC7i6SLxdmQ0jIIbqC/uao1ZoFMOdRDX8V5J4MKKJ
yIN4muYeUMiuxhtwLSJhYFxW3w/s/eZuH3e8PWTv4ZkJ9YttrFBOUFPZWAFRcZ/OVbtvvUCSuMPB
OdbWYI5fxo2BkE7e9uOAc80XkJ2LeXfZ9tS6vR62W4biavhelBHpFWACYbokoCVdi4biOz3YdYmK
0NdPH2ySiv7o+wMV8CdwA2CHHH5DoPviYQqOkG99zEcBLvzx5u8E2P5cKcHa2s1f7fgQN5mJlCk6
zxlB6C43kTQbihABqj4Pbsx6CAPcFMdOZ7QXMSUptXx8JcwZizatoLGy8zqAGMkpJgDBkuduKQrb
B/YPC/hbqDqc11AupEQcSz2Oie9VsbxhDsGgD5hHvvkribyBUIt8VLSCVkq1Eg3TESS22yVTiYQI
yqGp4tTHsY+HtwsDmpUe026kBYMZaEw2scFiO3FdLvDJ5cq8tzlkYnH3Td/k2ExAie0RtZP+UuUx
gozRxi7c+AMD1jIP4XOgVcZwtC0goqEPYak16WE/dMZ9+N6Pq6khWyPbecoWnf1I90SYM74pe/qp
klk3gD77ZMRC5OnYr932YsvR/BGr7gABDCv9KaSIJ2TbLpOXrY//l/Ijxd3LiG01pNAamISEgLkt
/v75gmoOGrtAh70A1iMLJI/D2vlErA4VuFaxLDHwYgUsprbINhKnyztrM+oEqIyk7YEwkESm89Xp
HttBNBU0iSes//gfgnYgHxm3HnsD/e3RfPfVn2l77PQrRxN5V8oZ94VaaDYNu0n+C/5yl5KCYzSb
jxxHXg8EIs4Lk8PQUvK/4m3KdTO8/30CD/gssFq3hPu5datFnkbvUFaMzP9L1v9sZQnYZ5V8yA6f
NmKRwasUhSjEuDzQMmwgeqMaFIJac0yoEc7BewisLgUU+APIDHZEbuvkkXTWCOwcQaL2pIfheG27
MP9q13KwnVkdy4mMtmJYmg+md+dUnV+I2YOyyT5mpyTdpAXoxizZTwV9rZ6g4kN0ELK2Z0aGrW0N
EZpKPxuK0ENJalb+5IDZ4DzalmutlLYWgicbXRjZ9Di0LrKoQ1uUNWjxrKm1qPeavyKGnQMyFQQh
uyWOpdDrqkqKU1MdpxFnI0ZmDtA589saFi3bbBn1wK+hAkb9iRVoLFHqeywcac9Pgny/ajzfSSDV
5IWlmNMCOgO308OIdp70kOPTD1+nOMAOCsJIrNBMxYcyuCQzBhU4lemr09zh3pVH39BI7oLIns+k
hv1q86kRLj8nGukqKcTGV+8TBFQAyLiAbjWKCXdKIsMOFpwozzYX4lPGUCCgw49YDmnks/YN1u0Q
BCrFZ6LM9lSmtLunB6oUNyv70Z9aBZMF50mhJAqwcZc+qN3W12rd5pGLNUqmLrjLfopOL+CgFjHB
3T3GYYju9dGa2LposwTYXbBhOYvdFatTV6spI216SUiDxAOrj8DxsGRCwlq6ircNiB+2J+ziHR4k
E7/MJM+u5d/SEKZ2CZxX7/9lroLozty/We+ShK/17Txw0p9yxU1Oj0DcZqSr6lm7GwTff1ypFcoU
jenGHWDK6+yDItShBvjIexRoAKxBTXwP0yo4Iaz1a6HSxcN5KCTuSA8bEnzg4mMVLKgtJq2zPE99
/zxd330yFRCP+EaWKBEMBRd95n/cENQj6J+N1Vhh8RC7inKNOKYAknw2lYGvT53pJCPA3+Z2AVuJ
sfkgvwRvuqva/qWbsLVyu0MWqYiwXUVdh6dAO1j48pWPVPEOetKZACmvFQ+axb2zgRR4w81L+05/
oIPO/PiHBQbuuZkFa/PeKGuHJ2X4x9kP42kN00fMdmpj7P/he4wPGYM1pYs4tgzFSdy3hY5bR0J8
cNArYsnMPJqR2FYJZwfTpqUpQfH3pPHnsZuQ5DaFm7tiBhEhI24MKn60gqUiUUxIzqKWPB8WTJhd
K27m5tHHRSSLYyI2zDsF/7IynwbXGZCp9+3t0CU2vVTxYsZ9sDaGfCX80OEgpzjFtg+ORKCD3xyQ
ewf5+XNnCreMxf6sKtJ1rFsuut1/eVzT2zWm0dX60wdM32Ys7GxD/8pxoI1vjNS22R017Rz0yS3p
9DIgCOVd0YkBDUeepbMTVL6nxfmWikR5Gc8v99DC6sy+WT4rhhBxiTogMFdkJnnL0dXxg9JuaX5R
gCw10NZXwOcKWSUVt08sYgHzf3pCT1Uu975v6CRD02EooY9qKsx6ExXDn4GkilSEoLQ+hHgN1A3f
muYnk13D6UlPOvCJd72ZLhK3rkpfSVEToYCbGtNiDR0zqYyRw4jaI+OI7qEKTjlA0+0/ShNNhs3z
+NywjQUYAfqwdyae6m051wTHIDUVqXJ17av6bJFBXfuVsPZVBzgFoYAmiuf61fRvEbKJ4pDyMI2l
tfPsnPXyvV+dWewLwjS3hVPXMECoIS3lzu+YPZvySlxse200p+iH7K14hoRavIhiWF9UZxYWK++0
JOfbVbnFwNj9UOgPMAWwGKDBhRHOnracyj7p9DPSAMejZ8Td04Zr2xLNELn8R2uzyqyRgPgD+9PC
eII7hIQ95b5wSrnFURApYgLtf0g/Cnq06Dvqssccw4h87XhinrDqpkS9eGRoSOZddtfZUuZd240s
GY+7S1mg0lvAXuflL/BJWL1w++Z8py13yWAwt4Ew9b8RkYJURsPmmV+JIhotkLpGMx6UF7eovsXO
5QCPedTCWZC9kJrX8uMXMz/9M5Jq/SguUdjrvKZ7bmtkVhl3saNJ2eka2CGTY0e+GNtFtAWB40vE
ZSqiRsGhrTe2Q7e6XPNw84AU+zEtAWpNW4uLRz8Ugb06DEHOmvZnSvi79IACb3q7B0zLizaDNQQ/
4X27mnuUpQMRcV+JxI359xlFLfy4JThj8IlMXt8PPIuEJDd3IWcUzv7ZBfcbygY5K7tYt++zdQ7p
IyzEkXXJ6RZzTNk9LeS4ARfcZcAG6RJcUi3KVYGTfqj4QnLFXjNh5YxwFVJjgxffEsQkbd1re+wD
RksGbv332EErDmMNUghKl3Fyv0NZ56SP4Kathz6K/zcEyN3nJN2TByPz6YoEBOEmI7BYpPSNKzox
AsLl0qcKq5eCoBL3ApWwdpFIJST9ZMdGOKx+yuSAShkE3BMYjiCqFeEuqsLZec++k1tvSU2117+r
RJ1Db/etGitvQ+uNh/CxfVeQVOfxgu2SO0qB40W+B7ZqfriUmndj+iT/P0cGz4N+SiReiUQoJBH6
3TbJ6k4GnwQqrvGYwDcAdYUZDAGbxaqAgK5loBc23UO/+i488omGhzSTyWGTRhNdvOf8dc77rM38
bCt4SQ+qOeKjjolNVH5HUX/oUQm98j5C2m6MJqcv0Hg897t0YFrWPVponCiHqxViVfe76xOzJU/j
M6O1QqJOZu8H/abe0jtIkROjJKjo9YItkU2t3CtPbvBhY7aHUJDvEd6EbduhVSw7rsQy6huCVzbb
c0DcVv48E0OFwdjg5nKov0hUNSCgHQl7b8Q/s6m8O9gvUPOYUtoffMuDHLKY3hvtrDf2vE7SWCxv
kFpbiwdNa1bKcybsfYY1ooT2++mmInKh7q56QhcdT869sIdEFpB4vV5rvVUS48Kcp1iDgMkaMv62
WnjEXQYMNgsCU+dExxGu9RyR4sUXaWfGqNvKtfAdLyDZyIf/lEBfYfYjbgzcEhubfv3DWjSJNTWK
Kmvp3fbGUsZc6lnakpIpzUDVUYPhRnoQr+iwafsECNsLqKIiNVlUoS7XPn41ge6fDkiPkcbO4ZyT
xZXItjR9Y+eYZRmVVYx3RHGRj6xvHFiTJbdAvIhz8iJH4KGpvRs0h67zvQLcUWcF0nBOeN8RAMd+
ayQ1odMzN9CHZaulAW85aQs6D5JQTdyohOSqudqtcBCIsOd7z8bpSIJVOt5HEQjRg/7tC+w6CVoX
l/2hx8AT/Rgy9BBtdZLgPXrb/N2mI9QERGR49oCLCIAA1braKAVLoswQbWCK1EIbtN6Dr7rA/ZEk
adh1khtDHgj6oJXSvPezq5WomtJXvzl3rHg+6emjeMqwih9gHcPqJau/iJFC3RNB/8jzM2x+7Mgs
HUmFKP8zr+okGCrAZ8W3zG0vm+3nTQ9+ANfiL4BzQQ19JsWrLFm6P/QWwZEb2X7sVzjY46kBr7p7
ufs3G3I7Q1D68TuCqYvpvvifAjqaRXRwR3YhBidLkO3zfb4SOzgYX/KoH26R9c0/VYoAiRTS1kgB
bft54QqdnfGxlbShmwjf4f7FPbc1y1XxTbG/9DXzRnaNUDe1HalYfClHIfMPMPszn21IB4JoS2UH
OXnnbdtOezLd6xqJmAO6yD/B5LaVv3VrGqVGuncuvejkc28jdoj0WNhO4QhinNsrHnS4ej+gk1Kb
cgqBEnqW77pYLdBtgefwgjk5ukVrGwxZvIV2slLChPhWrYP7oT5FgeQ5+cb1XGICl9QWx6IEckI5
lWujgg5JD6bTYeGM0RHfOR7L3RR6K2Gk7kITYaNqOHr2dPlsBXfXm5T38IUloWWp3H7fORhncsQm
7pe9ATMg7STbCjBtE86SDMo9euJ5s8mKebVjHgcmTfPpN7foMzhW+XmivByXivI3z0HbKRrzuy2U
MtstMZTnOHMGWh47RiuCOj4lt7HP7GPtv4P2RP/eyAjTU0vvmhG8G2Ucja0+awBQPGiUjFVXPWAr
0SPW+74otA2SHUo1mTAIWhUYkfjQKTaNwzaU1C5/1LgEhoK7SNYGVL+5b/PFAM/d10KA8N7KpzWM
LiYOyiXrlFAdjBYirZigdGQS9XUXtBeMSQP26nl6gcNPOTyMJ2tB8dVnkjbwqAcQRYq9pmDTJ9Ze
T7HbLooFL4GJZb5zVE2YiJB89c4nLMl1I7kNbLhthJ5Vze9xJC5HZMxgW5gsYtxaW4ha06/3R9pb
XBAWKeBfNEBlq7dsfeR1cq86zBtRhm/OuLoJA1xMMCyR5WzDuvrb5rBcRswWe5TPzT8rxUxepaWU
Bkd1lgVHWhSepjrgCzohp/UIVbel1DEX3Av4hwQhxVXeqQDcCAARET7ex3Vj7WH3RqSC0/W06TMJ
Q/cxN/75ColPKP2rRhO0wU9xxdicBXZcj/iPgAtHT3T+zuiP0WF/siCWdURb4oylr259xM5BQvgu
V6gzPUL2/fs/6VPyBmuSEX5h5ebZh7JGacDHJc54UtgmvA6g7Cxe+2j73WfgQeuZ5a78kRjE8SGE
RwHHjZBqzPyz73/O7OwDp1a70QhuzLjWcUQcJZc8pZBpvl+Matrrujoy2yqE0hJ07EEmA36Uz1Ns
rWOhU+R/UDUWycBP5JMt2+ax9MbRchLh/euu7nECvFyOddVRTvM3Hh44cDeQDDNSA65WRJSrbOQE
6FxeAI4DE8kp/s/PtEXuc4KoeSaAACrb07nsTAaIh7qu5y/sH0stO/WPGZmnmGQDIh9ixYir5/XT
V9OpjcGXM9ZYe9iDPM1WZkyW85qkhW0UKNQ/JfHM00//UlMeNCx04Ijqfr4suT5qhT9+9w0E4GaB
nwgSJjjGR2n8Y1d7yTVxHaVs6gjZD3+PsC1OWaSV7DOIgw/yLezlhusbfQrxYwKSC+dFP5iujY6c
iNs2dgqMKirObUJw9aVwJM6xckZMm0EnGsHwblPOzUljQAm8GAqClS/RxBsyJS05LqYJgvlu903A
Ya9amPCe8bVEjJLCD8J3wfRJ1jvPn0q9ICfnDRR8wjAtkgXiqQREuUMiE+BTkbM5bQ7/O3aWpctY
WaPkDx6ir42ghVH8NyOkYCoMRKvvk/zsVlY50PQud8Tz8IIrQUw67DIdRTsVNvcGXvy7PUehI4sv
kONeAruVooye/fsjSRjCtdf/WZz4cF88fXyadog9sj9flxtxq6skF3BznzJhPRAYRNSd9nePAP+i
jEv+VU1xHi4nFg/IdjcpdCa7sWb6xutbDsnNro7CCWXVzx52+iMOpJRlgNzp0OT3zVU8krdf1Y9O
wYBpXja6U8oPj6AkWNZZVRDvSELAVcxpeyLFNpG/xSWi6VztwAT1GqEKz1tS3sFAB7APdtncG7/n
utR3wh8GfHWSsvrjeWKN9M7dBc6jr7JEz7NlsT3/47ugcBb6sh/mVHmOKlXMBGyfkVzQz3qukjq3
PYAxJwE0kwDmdBJpr2hHzuT54MQhxemVRwaWXJOOv4GcGlNG9kukJjM5YYdoJJFGYncBe0JLIwOn
2CSpvS194y4rbgx/3D0rl9BShVXall1euMes5+pR+qBAFFxdoY7UfP911vaNLYEUgeLpopOTy3Gl
7PPueriwpLNsbp+1qMR2eYHgGvAQznoN0Y1XuZFqWVgfCyCgeVK8Rb2yXo9NdrdXz+vP0Zg70PkA
bTN05q6L2x7/rL0o1lsWEmGFSNt1v8sPDxicLonCtpw/PEYjlYuJwzi0nEX+I/pBat+1YmP2VqzJ
hrAxgktXqUxLzWISczDhFF2O1WBbcJJn2JisarKK7M5GP0dv0W6uPbwu1zkxIWEELAHiqUYy3ell
k7lJzzfRWXTk6x1bR4/8vPHFTKoRnsY31Je76dPSineVv7QAjfYQHcSTSkeP5IfnQPp/mPCToVTn
mE5zbIZWeycrwOSlLmbNfQeq4ilcWvAClQlG14LLf5NtPaeAZ8ApYJwwlakZzCwYsJuvaECtpUB+
RvGUiM3fND6mzrLxVfM6wsQPF4MDIYG9eTuyAvNSmODh3D653gH0Pad9DzXr11vLxsw7YJ15Xrw0
in58CSEIw2QAStyQwaRb7AgUYnJFxSKbI3vy73nblHWXoD46VjwoV5HM1dvw8PyY2DHrPdh9j8Qi
BOFSlGx92ByWg/xIcLzoEbHBO5umK6P7JBJghp86ggK9L7VrS3Q41gWBKL9J7iUeNzo1D6IlY58O
GdYLULIqNceoc9wXde8OasS5ImR00C8zbX5S+wV8IqdNNYPqJU/Kh5/VXlV7F3B5PAmBAuzJjfBy
rYjYkeATE2HElJOQF6ckF4YdIF/Dnw8TVmfPbq3ZhPa7iQrwI5kRRGyp5B6mSStgxDL7nqMMOKwv
cXw/Gz5+DoNbwFc/sSDdSETX4PLQOUfYZOgEN8Swdh3Ju0Le920IBspicsqy/G9p70mEEbbrIQIo
b+9P8pcn5hTvRvGeYOCBRZo/yE+I4Nm0q4pjQTzpFqfZ6WX7rngTKSUq0OUKIaMch9ttSSCsk6Ck
RKNmOSwEvy1276gPMyRZMiHQJsFLfX17gawnHLBYsLP8g9usL86cb63GU5KBIgm3ddVa2TrOG6IF
aZ0Z8qf6I/Wct6JqITSD4l7lPOi2epV3DOx4D91Q3E7MZ4ngSJfRSrNang9Nogp1u0TZmTjdLNBs
3sIUIlZJdFAx4tf+ukR8LlXSDb9Z6UVNnDsbRxCBdBBVHqjw99MJV+xzqXL4AeNiXCp69P5r8iLW
GwXfG0oNHV8f6G9UFFp2rvTd0C5LFpQoDD/XdkPEgj2sI1kmBZ33XFWbg43a2XjbEB1rkv0kKFX5
vSklDuuKUqFtZv2vOuIyAQ9Ov0S28CX2bWoCYJCw6FmrEQ0jJizExYgTDPCrnpt5mpIoBp6bSZLx
Z60ogQXSDMTgp5lL6KiOP+wDrDeqqWaSPXWGZh+BAz3qT9FbiZLUto+VO21sMA5x3PcPMvT9+QTa
56xKKnujLvYT9hAurNK7QYz6Qe/ImfdvTfhr8gaxoKrWjX78ifquJrjdLnRYpKh1poRxKpBMnzIK
2B4R2/lilplyXxvg/tLLeRHv3i8t+Yh0cQCc/lXgr07sG2avZroqmtdDinuysWLi3DYgkB6eS5yk
nJh/jkh86udmmAxOdpk8S9+GnWygLQ+zm7DNUjBWacn/T4/ydIhUc7CJzzbMCxVzhUeQ/3wxvRlo
9nx0DhNQrlpN3ObCrfuTUNw/Fv/bRg+kMZz9+U69J0dnP/blNWOUAF3b3evG95jWCzHgARa/T/C+
tz9+7sEoUVh9jeeO0cPeZdfsRfco35q75aNzXN+F5uLYFzD/qFpDwIQjvEUfLCar8yWTus7uc8Bx
l27ewP+TvMQAcdhExmwGSpYWEwc6kHCR7zstv4PfkrlfsEx5y8K0/tMaQ+6fNAH+3cbtLT4vbL6R
Si3S2fKA9iE6yBntmtgOrzBYDOSgBsLBfVSNRI8D/LXeyq5oDSoo2L2kh9o/PWoPWa3wCo5bmDz2
CtGAR7yJl/s1IMUUk2P8UU0IWYEHLiyVQfkfrVsKtukxR1ftIAztLIHAdty23H5P8n52VGm4Aaef
YSAYw5/Gwa+fIBbmbZfgkKTYXIeFgLY+AN+a/lMZTCQy94TOCqKMHu/O87e9nn7TF5cUc0UGe3ih
oI28FsyjbrqygSgVDkOC3rCfsRZDBhF/kQem6Cr5MTi3MHt7q3VgMsT6YU73nlQnB3Q1pdWkGf3m
HV6FpoCf4grZrJdkOjg2e9oYZWGEJTaQuCTn659LcF4+HxsFijOYnxQMJBadUq1+vGv1N+t87rVz
FTMlAjNchSMHlHrHxV990sNJKRrBsQV5WSiHm8xACQyEuLcVPeFQPCksJYmE6UVRVdsw2TT5en7V
qITsOGC6prb9KL4A+hXFPB6mAMR82YcNYH6X5Hn8JD+crir470SsrzM1pRXPHbYzpdaaWVtM1VcH
0el1LbtKPuvSTqozvZK+TNe/9fR2UJFXvqUxuRfvTSilTuGuwOwc8GmAxr65UwdDYAMD94bDPdgZ
+qjf2qa0q+MvfWNrA1OXKS9ugVbEFJmcjpJP6XXYqj5Vbh9kg7PCWhz8e1T6urKtvf1UPk5DCRyE
H5mUj7pkRAWFC3CZ2ekee4qwhWEobzkSNW4wPiaQ8SvMt//JS8Ro1oBaNsC9SzW6x8Re+osIUhwT
LUtMuyyV9R5/Vxs2uOov/TUT2cVYMGrspwsA9jqScYUPOUX/fBN8vMSBf1y2JykCrtEx03LDYOeb
4LK7vPDcid/4XjIR6zLiA3b5UzJryjQsU1rjVdzhcPNG2fjoR8SsUjQz8ZrOpkYoRPUqoRuMbxj0
CvIcb3PDkwJq/2QE5wylaMd5lpXrwWUMSBgaAuiHwZq0RvMRf/+Y2DlXKQW8QZV8pETC7iVX+pnh
yBH1XZTM8DkS8uShYMgieMKCZzaChT5V4yhgETcqgza7vLmk5uhBI45Os5z0LhV/8HqPUj75DX1B
5xhHw1edvIc2tAXFDJJdi6vQ4rojispTZBftL6v/2PV9iPttrG4ZcPQnpbWWiQ3mMQqNR6tkHEO7
6szFXuvaZt6RJmcg9/zm/nAqwOAGtLoNrN7KmmsnVoyizV2CqKOa9/HbvOwWBN3DWdK1AaqTxonJ
5ZGzMUFu7oE5UA6U35S9rKjK6FppJS2mC+Jbdk6bNeasvCw0bgau7WVupgqi/pTUbRdU+KC85CRm
7onWmQd9m45+rpNIODnZGILACuCFgJt6A3IwkGXiOXPw87kBMV3W1zxDmomM2bVyGIUEsjKzi6Gp
aOwXLyQwL9tS0qVz3nIZRoc0kmlraFmi7JYSCas0RlEwjt6swEea0NOdou0tBYG/IrF3iwzWQ1KR
LO8RG4fn82TMZdLSPPNXCykkV2pbw9kAwSb+Fm+Qg4dRHat1Nk1yXVquTX3QNzp4kTx4TD2VYQtD
Nny+IMDjzb7r9vWBglR8/gxWPcuMoOtVps0eiSPuq4wezkoXV0rgTRYNWQNfV6lNtPWWdQLWxTyu
5LTBdl/Ofg1B0tK3k39CuBEdDCFpB/IIRfpSO3i+OX779FBtW21oXLp893lU1aZwVmlKd2YkRtkB
u3MC7wfmOouMs80/ptxUMvei5QKhVTzMaE0dBxfUgkRKZxHJbx/ATEwburGgx07jsj4Ctuxkb0u5
TLTm2yM3Cxb8Bq9rpyjBFvsgchNiaF+ZrEPuD7mU90HO9kBp1lqN+uRAdlm6Yx4pIYEWp0VyA5/L
okaS6ymdQOVIlCfHP25UaUb++jC9HvwWajDh5YlA9QRv+EySIiow79wgDZJkfA7LYCQkuiGK1zrW
zEFA39y8vuWa0m4v2Vz8inyxAeo1rnS0vxJ2gNvZupFMWTp55mAaEUHxyRWBj8w7+pUNcT3oBZJg
mindSw9SZJ4VZBoj4W6eeMtCPWREMilqZpDpU3XFATUCAFam+CQ7mZEV9VMYe5FnhNxX9Px5+mzF
XSon76FJi/qo8dQZvNP/Eg4t1TZEPyGGuPVstG7af0qrWb1SLbi0LQFys/+x3Xcv44X2zyRVp2uO
hvqcFj6XaTI/olS5idc8iVw76Sp4jOI3c0Lz6X/ETg6lbj2+gtqnz5fbisJ1KqW/mDQR+dDO+qYd
U5iOQtYj4dqq5sQ9yE10x/82dfXv38uPNgv8qY6gb+hO1SjFt0y1xExuwJs8/fKRjn6rPCuzvDD4
QWA5SMyyCJXpxfCa9XjKpUgnvTEORk16DRISoS2pGapu1j0TR6ptnF2Ykfc0n7kdjYCHlTM1LBto
5D4KaGd3qIsZNnsAbIroJQ1F6rw7cheW5Qb/gPdZK1sPOV8HeaU8PALdt2vinwXhVeS0O/vdjCIm
rYAbn2seZ97+IILsmXiaEqiXKyUzYe7HtIF+mbOSNiuhQ0RuCY6tCDU9OjYc8a4SWrEhj0FE945x
PtCMQT6yYG3Xy+tP4QXJ1K578D2txZ9x1a+Y1eIpCOQ8CeHzx0YlVZ4HbD18UqBTZkzxqm21d2Fn
eKCLYjYsac/+5CbTVUUEl2KaVBYuz5+agJ2iSyGpHznGw30EZLZa7PXD4vi+RR0ab5YDFdEP3V/L
x6ZUI85D+NjRVy1+rq3PxYIFcjWz9oAqAbw1F0zeyiq8+J2jx4xWVVfebzfbzcxcYMbShsUbcuer
JrfT+MLIKiuErMqcYFQel5fyg5uTgZtSGdZK2JLYcQrNgXYNvUPuxsEy926xUqwI7dVVsKliRWoc
N+eFBtZ4YDy6+2hBKxCTCtY8aQyUCPt8E5EM+SPt8pMEv9IAgSfAsa4NXhs/mBeEoJQd33KxqvNl
oWycXlh6Cm8yUDNuZz4+s1y0rBeVbO5+1HCJx1V6fHaiXyw7WNnxJzCKjEIFq2kMnllGA0ZYK0Zl
ghQe0JEZjDjRxUkQozJVSJiqTiK475SajmQ7JN2eMBIrshWZEbOLjobAD4cHUdmg6j3gbkdnX34T
F8eJmLn9MZ3l9oTpDyzWZycmtU2X21PuA9eeMrqZ4opB8vynbvQNK3L07yCOVa+Fr0mJiDzvvMGn
kaPMcjxH8bjWuKbrqJr2X/NGOvIGgaaeQ2O4VFgYtCGF5MV763ocDgrkV/aiiTnrbAPXK+VRJZTt
q0t7Gv31g5xliILcJm+PwiOU48PawBvg3956ZvbvDEca525l5o1uUns0/cyqE7bRreVHuMnTaPU+
U3nY5BtPlg4VU5jK+V5s2mYfUt8kuMQ5M8LC174cBszcb0lZIe6mOKLy4HNQLLiWWDpVEp6D3tKZ
u/EEJIDqj3rtcR3WF/+ZKSxia8xQvHYdlk2YAEJod7LCGbwk2eA/dgi8nTtov5x6bQO5vjofwArZ
Nb2uJYopHjRgEM0ewPeo6nsulFZwVrY+bTvE/9hgt6xrUZYpppJaA2Swkd4nWGIH0/b/u9Eiq3uI
N98twRHa5OXxf7uDgFTAMjx1L5Z/zR7KZZ4qprWOR5/ex5J/VHWEIq3DdYeDliLMpK3B9tQj9m+v
y/OX41g6/67/SvDqkXkuJejSwee+2NlJJSQ6QQrC16TnXtXW85M5u/r+WDJXMnt+blja+wnpOgCm
KzP2Xx9dkm30olQXh3fDG4PluAjF/cEG/bJDH8WLaxfZz2vOJ/mAXW+ZH0wuYyi+VURfRuMDSDtD
GhAQ3ExzbE2w3enOeSD0+uUJPvpeskRP0XcmgPeDQhZR9yRzuAspyCyisUa572EsqcqUCyk6jz7H
h4rwugXxvXSldL00HZK9yGgJJoB2wQLZvSseNJLgg/dm+oL/O2ao6NRzSEVdYhggcqlt8zaSl35s
MkETaPq1k8NqZY1l06g80hYkeWlYKKKN6vzDQpNvkC5DrsD8SteSV2hVuvjEzO4OTAFAcSm2s7DM
MHXc9ibFWRA96ri0VYzZTUlJcpK/9KMda34FlfT0/U1Zub4OLR85vPwvzxQwqTi+8URp6CBxOznj
vxH8JZuQY8HoN9s1cplCNY88uIvmsI9+KORjbKxl0gc/rrnAgADBZ1tY6KHIIcysmh1B/tu7bSEX
Py3/nJwGdXLOl8sByoefswxYVXBmCCb+4xI2l047VyjnDW1Ptbsf/7+LSihRC4KzMgT3PFlN9KpE
kx7HgGni5pbkSx0YkWj8mcdqXrK5YrW+oTnGQN8h74IYPLzkw2rnSwPnNab3piG0//VB0aO9cr6I
ZzSFhV7jG2nqBEKRX84q6s/JwjVGQyHC0pzfKtHgzplo35+uvmIU5sE7s4QYSNPebrLxNxn7jM2F
DKdLrez+1bXN+MHw20qsIXbI57M1pGdfU8ELJDRkMnOl4qTiVfYZQk+Y0GY4NosWyZG8yScJdByk
WQ75cfTHTF1oTi4IlTczFBpaBzZ1yoSWNF037igZ8P+JBhuELJneiB9BXwsctnmZOllEOGuPDlDA
KD8OO/nTq5pzUYMIh9Fz2h+Akq5oFml7OMjuHVHlO3YsePGqJTAviZVOAqBnfbNICIWg3NKu4Ohf
iO30RSuICJlRagL9YJVYjKU23ukbsFMkGAQaWe5vD2tPYt5J/PbPvnUrGBtdKKmmsxwK6WWzTFMs
3r9RU4FKQO9PEqLxN5vfE3S9dGm4RUrEBkmiAB56sesV4OE1k/H8GP0A7vX4di7ggODiLc3lD9s6
ecEN4Q/M/m9HF81hGXkwzi5nJf7SMDKHDkLpxK1WOa2l3xvsECwhM0v/sbKJqwf8FapnmqkF7S/l
GiAkkbVqMq5kCuIb7KbCcfW5LgdRXgf2jmv1ZzMn6ima6HKU3zphQOflU+Qt/cs1GJuj6vp5jG+W
jQoUdMeMIvVzdvli8ExkvoyfSnVRjP/gqi7NLbhSrFoV72UA97wGlVUeEzI8DHkmCu2ghghNWpPb
JsvE6PCbOXh7tdzP6kY6HHlyXUVdgW8CFNEQ0P3fx9CWyfkqMY7G5u9TdHYmihfBsPq9uSJydyS1
ce1FR2N+Q4/Z9D3rCv/9DRYptNt8HUcLaTGtecMdlX3exu3qDG//gqkSzjZQVlo4botbw0AnLK9R
C4DutSHXDVhSY48sDXjzIprO//Wd5Kj3lzKON8TSNPGFvF6SYgJuVL9RLlFk9W3E7uk5nMjChUsy
fWVwn2lOa3kPUEZ30Nn3XZIFLhT5x3o+Pyv/te+cJlU/eU0cNTZnA9sJ+NZGMJuZ9jndmRMaaZzF
vIqalqfKldYPAmvC6x9/4tThtNhWfghKC55jxGSTb7K1p3axTTuZ8GO3Ns0EP5mHEx6qE7pPRSm4
+YV7ZgVs7VTiZcmtb6rPvMLbh/wfPISQ5TedKLhuvKWxiBYUKNolZCRH2kUtJ3e+VzhUds093+uz
aoqB5oaOqQVYMZWVyvPQfQ9MeDfcAczkYnJ9lGac05vfbHUaE/VBoxXBK9bPaKCz8byY9qihwcvN
DCmt6OzExodMGFt5v4kBiXDltwTY8vm0v4+xLBu6HfTsYKNl5PUzQ84tXSC/2UgdeV3GImw2vfnH
5w+it006TzADpl6mIHQIju/u7HMaimdmkXS5Ip6e+rNmPgj0cr6FHVCCghV+a6C7955nnclnLkwl
3HaaMSaqaLSOXxPzVCUZ94o3jbrZc20axj7HezQW9CsMrjpfKx+FSSjkb33dOMrTmx7TKatJLXG5
GWUaCndCIJIUcCc56OaCohsG6PRonRLsFUGGOtd14OorqbaMDeEnPDEFjfwfwgG44RdAoiyIbsTg
GE2GQ46AYqsLpnwt26vDS/0EzcSM7EwQ0E2/PKVv/liMDq09uYrsU8nL8MdJ7iZccwWRD59AiZO/
aSyPwR6ZdLEa8pgIqi0A85AO2psxcED46qoZdhiC9PxWyFoOrs84rZ4q008BsrKzitWcOp1iCep4
4pEksy3cIeKaR/DOK5z9yWppJq6KocBMAxC1zeMFd02tmfDxHE0w5y9AnbDeLHPMG3DpNwqoTGyO
Qhg7EY2Ja0UZgKy5oFLOWFzpPNj7NihZrr2z+6oArg3nPf6d/57AiUlayXbxhMUtJlG7amVWUEb7
B7VJ3Gqu1MTPglX+xbKZmxUGDyvBlGbdqS1Y+0eSzua8OCBqltnUSAHSsxJ8gRdjTzLkx1E79wGG
QO8pYLLPnSpRltuLUQ16/alkQLk4XRraC91hrUAMFBYnVEGoW4NuIw2DvuqbxOKMQ9Hlpw5JwGdQ
NMXbPwa1sew37q6HF91BO+aRLf9WuTLBDv3u8p+1CyOOwkU2NdhWND4hRx9eSK2XMR2m6iK0N9eG
tff8W5VsLsVe0JzHBZjbJXejckjWfyXKVOJB4Mf8GjOVRDEEl674y/cOSIXprkRIG/E/vv4eXXzD
SgjLSrd6HdXXWSF6aaJofZ0GHY7/MxW3jGwHzAukkD7ren3dhBZxxDkuyFeEXcKUrD+BahzvY8Ks
IEBZOtJgJAVKz+0rJlXqRdQW9PopAgX6gGebeYo976eNMkbrZCXbGdyoGiibm4GtqLhozrBLO7xM
updJL5dt7fTdrJUMhOk8lAcrE6OGJgzJenJDsAKgx5tH9Q+hNHc+SkzAqzuO6BmZqLy18jU46v27
dLceJUwFh2ONQ4tfdM93vMOrTMeVx5MWj0ps5D9gJRPLVKv+YCOL4JBHPnf91pUJYwqYsbZCN1Ys
utK1i9OV1RBkcItot5e+md71pkJSXppSWKC4WQr2UZIM/KG/GRoQumg8SkqpWbMhJGODNsi3u7kb
V9YnHdOnZVweiNOiw9hvxd7c4vSQOuMEfN43Aw0J9J9lPdlvIEwss7Qx6Xv5kYQkEYgBZIPV4FUc
+RcEV3MhrDJgvMm25+GpjHvI7nl61otpRdSJh/Sf/AUg3QYAoXj4aXihTPPG1tmCjkADyCniE7bK
grG3+x3J5x8ZppuqmJvkTOd/rzef5GyePbZOovOsnG+blu1W+pvloa2RxMiOtyBgAcLoyVwtzs/Q
mtK7c0WZQUjXrlv0jCkP0E/DX9Gb/7mQXa/PB6O5s9ilOa23tQGFt3V2NdN7pzVRS7ePi5fukpEj
8eJbms+d8FF10cGZ/Wa/AJe42315DXbdSQP1O4+YpFiZVGa7CnGFc3x9yESdkthFD3qm5G1XLe9o
vGZyLnK0sHgcxr9s/6oLsRSyQrveGaTn1piJCmlTuccFof1ljF0EoZC4y67lzYgThjk+KMsLfeJe
nyeFAk2dpaKoy7d9FMAxDg2ZGW0C5P/fN31aQaSkm1L8bsVwQ80zsGSdgLZw8/uQ9j8mTJlP4tkE
MM6YVKopnkAPYJR1dqW3agePk2AiWLYGp/UZR0ituf6dNr7xLK4B4Szydp9cGR6EGhi4GmUeSm8C
OOFGkd7q8U98YB+7fMaSzFsGV26DBXZy1leIH9HrfQ4WS9TxyDntG6ksAnxGUwaoiMhfZgNJYlQh
dlwTYjltkJuSmLLfRUEgnBTVoNo5WgjaMgAPohHMvnCiGjkyMECM9+29R1HQhJPwc7Kqjsszymba
VNMWSwTr+7F9DIDBuzXRf8UiawIg0I4AFna5g0d3qwZldE5Rm5VPcPbQPSssZZjCQATNrNWeDxLW
+6YxahKD2ABOFilExxnRS0Y8CYDYJc672XwRszCsxSRmB0XPGaZgIqkfcDRGaB0+VLbe/sj3Al4e
Y0yxc66L7MmVKEWFYVUTMESTkf78C/FS/R905qAaacYdJ6HecdlHlEQO6YfFMZ70LPiApO3eliK9
skZWAQisd3RigeekADCcMyHSEhhuzRl8X2ZPtowcz3JHxyoYxzCHrePw7rHbz06Ia+ANKT0RkqE5
fN4zYuKk8RP+/v+gg4e9nf3B8ocqK/LfAxWZWcjKotZSO8xLrNdIfNDyOycP6+DGTn4ceFBKMBKf
tBlsYnK+RF/SK1p4HVMS3QVL8NwZmFb9uliFkDEio8h5vwCk50a9pJ7xtVDe7NVJxI+VWQjvEyGa
r63J+ulTzxw7I30uH9d2csZyI9Futn01e1fRvG2GiwSzkUnAVhxjiqTYGG1sX6rIk7+97Ak30tsg
ITviW0FCKsoY3RLqXFOW99tSSafrl/dMgdKHMVPOIeSWCLTimpW7rN/2j0s6Npc4etW3C2v2DxFj
IAZsOHUCzRFuVWNPCk8jO5NGCSIePrdGUztLTkwGjhPtP3aYjal5Hgw9Vsjg1bSFjRxvRScizm05
MxwljlKSBIbKTtx5cUqtk1jHIOQAyEKUrkMkuIQBJvFW52N9BIOWblR4YiNGXbv5MjIfwj9sS1Bx
2Wj1gMA2R+kq1Jn7/XGgmNkhbTq9OBm3vox8eEicuAPROlbTumzRZP9aWM6wx0IKZRLffLBfJquD
dv7toCzJI1JnbFGG7on3TXEdhekbyOnJm61mTC+Mg2vfVmNl3Ji5o9ZIi1TfmoXOSMBrefk5G7ul
1xYhDiM5byms81vlS6ArECHkXpArGCYMKA5L+Lu084qgQiITf4YTggLyoxsFU3F6iBsqlNn14RK3
pbW8zJi4CMwUXTW2Ddcnu+7jNTPgY5WxP5w/bjt6QUVgzoSrokx4xGmf4gGRv9vcwAx7L8OHbUN3
XBejDiRPW4R8agHwP7/LC9EPut4jJAN3SfQ0edQ/6304eBhugDAY+d4IpVuGNxelVE9DGswCeCYw
POsW0K+zz2MdLOMj4Nbwr+3qRi+vJWnbV+mchSJB1mi/ICp/vUz1ppSoItVzoqjvEaXon0GXMyFV
7W/H3yFOcwOXwiZzDJQl39p/ZG5cwWaGbfMucMecFLTLoMhQycWvOTQ7GudFXy9SRfBnhfK4w+jy
iIomhqxFp4auTcbe8QQwlF3lWZIJhOpvRZjjuwCN/6ztbfB0P3k51MJlj5FdeAa3HMkHuI/6Uz93
3heORyONcm2s3yW1svodNPlqeUyDFoLsB/Y6PIjOQIamUeQmShAs3Fg8+BkyQQhX6t7+KPemxr1M
jXgWJ6PPh6PU6ifcLWrO8EcLdciILIVKd12xf9Ppj/IDdKZvTFGg8DEdQEXzkCiTNv4anTvSL/n1
SGscs5pV+kn4E4dYnn03gmT3xfeDLdhyCgyv86b8n0KGKuKaWdIlU12CtGskc0Q1hYB30h+QKZR5
kb+3bfG7f+RtSSDqCT55fYXQ2AR8EMkZwChXu5RI7zGOKyhi541Mamn0Mym2Gco1IpFz/80KV2fm
Z8W5quU+0wK0ts8UIMGnWWqx3zgb+LZSnSz8XSTogLJ/cC5Uh5fr7P8noeZSr3EysRCMEZ8kHXoj
hYAKXWOfSRNOy+mAhGnSlQGsPiXPhxxD+5G75JenOMm4xo2y8JWIgG9xSxkhgO3AETzYxcKt5v6X
VnM4OdffSHXSrxCNc2EBfIuxE6NfHkEhPfe0oHcVKTpQ1FlAu2Xto81E1dFS6LiB4R9YderxesFA
7YqjLTzD+lwoKSgW0TUJaA0OxdLe7y/IkNW8DDioCjDQgqHe80Rx0IZQDcMjnpBJv/iUJs8v7b/i
N+v6+L/+cX74OHNud+W3lPqu/qI8TSOi/RSuYHRsbiisrRXqrvMP41BNMAaOfUSF4xMeIoblLApM
X7UH2j5zttG/dwk6YsT3JJQoJsOkw8nU1aLR4ink64SDqvPvo4zFyjg0MSVbcB5hA72M04G4yk49
4rz5DK5Rg3J2JtakqKvhaZu8YxChDr63XIWgSK1vjEWQIWUV6outdsf6QIjyfC+wbHGHNKJxymnD
Tui/t/QHNcuUx5bLbQjQG72vBzGa+NhvP17/7IgOIvT+IEBFQposebFZJGBPPd7yERhaSJkyLaTf
njhTmToUd38x3dkvQd+V+Q8XWsnuJNNdHQuPNs7wsSnGJmpbHkHUrsbERPPxYV3Fb01fvfwf6U2i
QfGXbB96/f4Pb2qkerxay1pZaovbJUQC7gFImlvQLGaxQaJvUSgPXdoHog0AHgGQHDxl+SAK3U5y
QBOYHn84iYSI9YbZKJgYW3JWkxl80RFsMYzZjIiQlDFwMJN5Wl6mqoey2b/t2cNfaqjyhMvvd4Cw
nvu5zlUDCt2I3VI8ExSoT5JTWKjo1kL/3FOQaD5BNVu4PT9Nza1kBle6keLjJlgpJBQiqlNtrCXK
+xOgaPzrOrR/xCsG3iZDc/6oYrLfzmdjVS0e2SNM1iSp+w/cHPz05D6TJwStYSl/GCf5Eos8EMaA
LdHXMV1VDmcV4a7jOyIxDsfgLsI1JTOTDb3BoPv5QSGgT2/Y2/ndxXJCWkUyueM/8OMZ5JRN95uM
RtkcD5z31HMuindWC8mPNL2Gq7I+zRLUIKmcnLAWkaVD9oXQTyxDGO4av0ayAQVq75joNLX0nR6Q
PiNlteDJjnNvPKVsa33YDt5iBUIriLvC4xIx8ZKRItQMvJGTH3fpQGi8ON1A3kdDPmlsBAMZJLz+
b7Ma+uWF40pl3E3WUFeuXLawjiDuoPEh6wWxkmb6Ftc9GLdDph/PjEAXtvTTLleRfinfyzU9ykQS
fl780xOqWAH0bni6O1Joy6fJovRgaob4z0ARLMZamHMFqGyvdbioAQsM8DVsII7r6rXaRxeBCqha
DJNUERRdl8tMQuQWRvyL0ZbnjQgYwyCBf+ve+yOvfE7SvaqDQF1tmTODlNnrU3iliB2D/MfNnLF2
bb/3e2Mfi6ll+iZS5mVH3CzdurcjJvc+0anUxLZi9s9d13XkTyxHMNl9JlmGouzwLJx28m6BvTFL
MnH424fdNnwgj932RcsIrD/cBy8AMQC0Bz3y0flbpxBTK+tLX0MitneGp0HBlo2cEkh7xZvbjqiH
aYAEMpatwBjc6tOxXkD5h9FuYduv/cP7p8/g5wykbA/JbggIn96GvFv7UZHdi2NpnIPItlXGTxbq
NBzVeQ5Z7c+wTmkQ1OurvBR6+H3ya+18TzdIBY0Hbz8MApkM8J6egzAR/OequbXKPTCEYR8aDlng
p/PjzlGEg0JBhUObA5v1KhYwBTUWz9xn/lv2ApOnpu4e0gtYBbFNfNhWF2Fgqb9JGAuLPqNNdAPt
9KLaoqqGYZn6kAhA1o+6z8EBPJRe8Ad2THU7H0CO6bj67vnZ8pLk1cFKNVAF7glCFWD2zO90tUN6
1zVNn4xpj/RxHtp1EOy6YfKKowYt58XOD7AtnBP25GdpahuEA7lK4WB6ngRbt3qb91Pl+zqQ5YfK
dkh8pZiHC3Q2N5oTZizWF1VF/I1+oeUR9A72YkqzTsX8ci8XwUmQ2oaSLdVgfcHnrTf0U3yb37G/
W34OLkk9w+07htXD+vEjxbMKwjUQrxx9+qL4vkOmOTtPyTL91ruU5JbWh6yHkumrmHgU+cHSPDAx
xlpqNWs8s3PM4MlkyCbwHeGjuY6yJRMznRGPPAUgx8/Jt26ALSJtkz0mw2qzub2mmvzGx/Uo0Z5s
UOp7f0XUfAw6SgwisLwCxwSL1Uj22XHFh9z+zooUl2cadqASCOQPkIpB+5ig+nvBaKamPSIQzf7b
g1KTouoakJx7Gl4zFCHeHHW2V0jEPI12rh1Kpq0rtK4XB/zO4jbSkW04yt9qoPWW0o/YXYida8bI
RjKKt0hDRDrlbjbbRV+gIpXOc0UNWR13mJenzGnaIVHXW7Ymr6o8L6OlwPAaxiuSET92YJeVwSQ4
rr0DQ+m24P7enBTiy4KE0TJYoh1/tIvO6eFO/95CRmKuUemLeGBkbit/10sQFVoH+H9xK9GrOQ4X
qw83zCy5Qg87xIgyJ8ZQDvMrDskyo+1pt3acL66Y+ICcXA/mMSCnt3I6dbN91e1MEz7IzeL9WxOm
BQ8Jw6k4X1y+gsf4nGYwRX+bBJL9zqWg1kl/5iXx1DrMyedwKuj+OSw0e6wAT2Jlomfze+eNPWZx
b9rcIGkZA8+pb/l+BsvEidQ+ZzjiK9kF/zLoLp6LiGPIdwsXErPAsbj/gI2V6cmXd+1cLyVJVxfF
Gi6QqrRkb+1nc/mvP7q04+erSBnloUWcG0/VBQzf/pDFMzsXwcH/Lg80aHMQOViChB5cPrGVbzRd
L6Cr1Wa0L/2NSzpKheJ8vJ/zuoQR29PUmYo0H3pLd1+3Aq05ke4IvAsR/b0fZk1OhzOvArh5uvYz
dX1LGycSFR3YlctJiixNFpTl3lXjkcla2N7SAsyauB8KsWO1M00BqPH5iC8KIw2bnrLOma1Zi1Wr
NB6uS/yKQJhBW+RUpFfVTfdWpNbs0E3WN379mkLHSDoGHPnXFrxiS5zz1fMWbmPZBTYkMgJBNJqH
+6VAS0qVHsLqWYRViZMfbBnB010YN3Kwmveul2j+qarKmj8mNQrmVIvQtiagh3cEb99WzNKdpjRs
FshU0U0GQvnJGWweFpuNo/JwC30z6JOE94cL55uVbo3peUtw9rnkjL5PsYWVaOTjUHLaFbVgnAzO
SQibI1PJDNPUYqVqlnqllD2pzatlf0xn4fpKBRE+LFKej3dfY2WrBD3qhq0zfWmHQp2eota8AUq8
IzgiqBU6V9x54uELQ/DDV8G6FcJ5Mttv+xQyZFDrhNMAFQCBCqZe63Q90DvYd6ZxjVyzeK1soc82
OL7SzA0JSL+83AsLG5IqQvtlyvpcOS4R5a5qSMRVP2ct/Wn8t/hvrRUpmWZYG5G8pKo0ZzKBVQOX
ckas1FZOSt1Spx3FUulTkeRqV2W9bc5ItFciOrG7AgqIOM8iBaY1outUnqwFCApiYT5rkpptq16p
yNdUB9sdKZQ/U/sMkRBNdf26pGaK8mmCBIEUi1D67y7DIlKSAaKkRVrkB240H1NUHqf5bIpcQOQ5
7n+tKZYlwh/g8Sl1R3nDEx/tU++ceiiRTtWFVIDXjgRhzuhe3k8ci3TlGyENffR4Y3e8NovyINUj
GEAG6b2fH9qZ8dsMzDNIYhyNlvrJ+Xo6J0Cx/UIq5Q/dqzY1rrLt1UuwK98v8yfLri2G4rvSll+T
Jkfpr+HqAXOcyNx8iZwgOpUk3eSV0vZ0/H20pvz0ywD4beyoGWkI+oB+tMNqLDEONc7GbHw5aEop
iiKDKlyVor/HL3cwq1iiVClvih0hF7ZbtNc6ulPS/4fcLxTOHnKDVMPkUH8joXuK/OpZ25bbKUUk
Jq3WlHeO+3KLllNpVnCu6NhdH0NnH5wmBxESI7wvy3KWNo1wXy23NHcdnvgfL6FSLWpTH1zBolkC
FymTx7BaIMKa4wd/ketd1w0UGC+58D3jhs6yO4ySy0osGvMfwb+1hhRWgpfM0zGjkUu24c/1Cr2O
NK/Kj59tRctTa00ZgF6p2MktNbul0fp65ThlP2GMIMtgfv73VvnXhrJeQWyJnskSQsJnuPYrYexm
VIe0xD2a3oq1imvHDB3i2V3ffx5uSZ+5zy+L25kqrOB7tGH0bZCZUBNRV2Nii2NOK4x2y2hc2bzv
JzkaNVCXVw3LkFR49IHmEd+vA+nuQfTnibmRIHM/I87yHTLtbNvh648rys1dSn+6gWv59lgp2Kld
kvoMqss1Rfg8XJ0buxEsaYkiz5MLm/TcDGlSLRyZtgCIJpgFEyUXur1uqIMYal9WlO9Hqip7BBJ9
EubJBKTjyejtqw8QISctEf3Z0PAt/GtgsK/Hn71mOgpaxTTbDc++lxeeXGVNryTP0c2PaCXWOl89
CIBb2vCi6mJVoCPLevSo++/muTDI3RPGlieBSf56PQtz9Qe5tP/qF5jXqt4mJrR7OoaOGeu8PEjD
oqPn5hDteuluzVDqsAqvSqde8KxclBqKunZidimjMVO6h9ry4vaQMjOkyVJKKKHVNOYayDDmsGh0
3uLWabAQFavz6yfDpuKCuTW0t3k87Xc2CCne+511AvA4zi+ANqYVvE4PSpE00GXA3P1xwxFB8anS
/hCd4OBLxozn0XftnuNn6HqYduGySpauFYHbThGPP+SrbkoBGQqT8i7pO0yPGgBDI7klUQKQu0Fr
1p2/WMBJ8OzKXtmB+BNThJ3MpeXkBjTcCPLxHQr+CTWTJvVJzzjY5bo0dmxlhKXfim1lzBw5DoEl
Ai+Ui6WZwZWbPCmYmHN8K0WCi8ZsoJELbyDgQujpjRvKKx58m61jlqLYy6hUb2gGtNo+MvG8GQlG
12b4PVlyzpTsFvVzSIO+nM55CeqZzUVxISJ9j1+Xq6p75FsKhb5X+AO5/v3vqJzDGDHATMslwnX7
n7RgoW5LyHJ4aT8I+l0mk7sjnrnuK/yFuKUCSnGja221wRmFxiPHSuh3Znn/WqgZ0wPgyuoXBtxz
iJXy/XuyiFCipo4kZU5i3mbt1/hh3EMgJ906YyowhaYnw8uKyFNC9KuvtiYcNLLdLEVBq0IFZqhe
3EgclxUR8qMZANopkArUDSjVhCvcazBiCPxoRYX3LwrSes1D0GQ91dD6Y9CgYMo3veDyrfPkVZV/
8sP8AyvCaVHTlJefLebbAan/pKD4pvOaLRTBgzB0L7mOU+HXwxTGRceS5M7zYGjePhCe3vRdg/PE
Uz1FXwzTZKaNxa7ki7RnHZUY3wDnlGCqrXTa0cmjV9PjPmzD1bTEQcAqAqnJKoSOiNd4ks+0agzl
d9PvsqVmsJ3qPYDF5bBH5SxWoy2NvkPWwOV4WFX90+D8R4s0DVPhsujSSMlu+LXVSd+Cn5mNH2/y
rXlN4Ez+qg3WsrWXhYd8hduilTkOh3C2WXohKex+6QSCSOHjCUWM1Qz4Rg3waMmWuPMBpcLGMKsJ
RitdXDYPfeQHWeZD02x0Bw7t2wVWZT9g/CL1pf9C9igHgW37KFntUBnLbmzCD6Ignhg1NpBcPGwX
4jdsvJxrYMweCVBcs+ogcB+GgwZDTyfVaysoof9JwJ8czck1ncUAcW25YQGitQLQnLj8Td5ZxzFj
hEJHUfAajeGX5iWPZPL40ut6NJVVJ8wvASPmcIm3HpYFGNLM4hCpEmOixWrDVKUcGVP/gW0kmp0B
erq9act+2RpTr81ifYUod4WsnasCtDcPjLEv5XfiK5smJIMLhHjcg4FlK9Wy9l/8psCmrgwPL82e
VjlvU6zoEgUGlbz5eEWplML/yRZn5A7jqXojp5poS0WDSiEkBHP8WuWC4XoQn08W3eO9kS4aprfD
s840r0+DcEQvXZE9EUYAaaezUxmCBlcYEA9sigUGBd1WP/+Ow29z2q3c0Rk2L4aWK3GlibFjS8Kq
ghd/R38TShdnrvch1XcjgZLK3gdbIwuf1m0gLMd6xfZoxxLxDNdXP4S6wODmjx6PAm7+LaAOMZcC
xiwUyxEfwXd9GPf2bUD5zIL1kGU4/ZmVbmqVkfuduE8zhlo2108Yxum4QsBGqwd780/x2ipmZLPB
Xx9SbuJ3v0OKzc+vjPOiH9oRGdIL30CWruEaT6BdPkKVS603P7rMNPjyTiR8VVpg9CN/5X9CUtbD
3t/JevkJ0k9ihSoV3kNFvFSP1IQOnG3oSf4r5QDEI6Jou68zfMMq+oRxQpm2LqRYBZPLqTdZZJuF
2e+QaHO0j6YvYcRqGNYiW5z9dP/QcT7zz8OLUnFcg9gdchGLMTVgH6tgZEv8mPfOQX93VoUHCW8s
P+M+cp07hrV1uyQFyPHGGkcsVzynfL2t4zEKKCuKFHP9XM18+ifQN+rgP9SnbTA5Lz60iEFCcE5e
/fBYmfMt8aAE0ojV/hm2zuxht3HSSTcIgoSAZi8t/YMw8lQWsKeKM6HTkmX2jcVZagmcMY8a5QnR
8qwGIcqZpQdG8/SXwX/HmzrtZ4vpohuXiGEl85+3Ibgk7YX54mmQVFQrjROQcGF6MCVMXqDA+SW7
3iZinbrjYx7UWfSLgdASnlKKNBI5ZkbKJPS0QPMUhUSYhPax+jUHAm+pYKFuGzes5Pj1TxXrmDOV
p9OKL3JecgbTB3EDnLVT8EjWbWlJSqMOKOr5EpiHDWILtrKDa+OOeSxpbz6x9kZc2Tu2qvKjYqyO
zQbAaKAtqquVkoXdl6sBRFj/cT+KQ7fPbafvYH66Qc2EYP8dqrultCDMKnvqEMNQBZLcsg3IJpBp
XBJFvKc5rSHoEiDIJ7OdFOatWkIQzEHxs8byTlarNd2QdR0NQwhJX9sgL6o/pkwTzcENQ7dB4KgD
doH++vOjOuahX2vKa6vXCc4Lu0yRyLWGfjOBH6snJIGMFnyyaOgB8LAnTbotwyuH/5p2GD6rHLWs
mt4tuP+CKG0Rng+vWF8/TcoFYxYixqEdvYX+BtsnhYP90bfaGXk2aoKu1RE3dx8NJa/IuQ9WBEqz
cJQg/ZeJjS+xcNp2mrtLM36QKblXqcXqmdtszPA921W7VJXz3TtvJ4EScIDDVt8bevUjYBQRQ2xq
FoXvoJO01GXGZMXyk/Kl4WXesT5r07Y8GzV72uG8CJR9Tqw7+wSiEi+o+Az6lGZ676wmhRrnMowh
5/iqnpiEIwYIXh2qKQ8jf+FlMUZ1vypQKypzg8g+jlzO6cwz6G12BcuBDTOj4FJy7zWpuMj6LHc+
AerJ+KEARzULgO2eRIXs+Hp0B0Rnn1B5esO73aR1miwblVSchCPoICyCqzMbSiBRM6IS9BRQazPW
VlrK8ERcrdpaUpxuYvO4b0009YTylnTp024gs/toJc8TKlbb8HzAXG6jq+XEa9/E1OTrFQ+etoez
sf4YQYoRIo6XRZ5gRKLPzA+5Pn63WHdZlh1wQMwbDZwCee/mXsvFLgvKtFdUwJbIfSQvWxJBLEFE
Y7Wlsthmv84yXi7qBi43k7o3nhCxuIM4shLbNXvQMXAYXQIE4jonE7j8qQXqXXQuUBDDEf/P+kMB
7kD2d8J+3aLWqD2BypkP10ETF9L85gY6S7gPbZIsTDyafqnGxDmrhr2HX745dqE4tBe31+XihBJK
PvqeBeWdqyJWHUP7Vm8llZDVYIZeRVF6JVsG9+vFI7dCPSUmiYFVgPVpg91F3pw1krgd/HHTZLO2
TFuEyFuOouK9JvaOgqfAiZ9J66y9FwGyxUp9GqLEfTf0CdquAXZC2rK2WGHV/65GNN/jE61GDF7o
MHEhH9DOvmDTyuOLlDdap7HV4+4yFuyl4Whe+u+7CVuaPZT37ftQjugSBQX1bP4ama+Gr2vdKEpy
6A2kwOqCaVM0zgHsmr6zvRxjmdZia9Yf+s6jPpHL4eiHhg+qhfSXES2AYDfCYo8xyn0vCF3mWiWe
dfPPlkV7+uP/rfI2g3N2uAnCZO9x0oub607/StBxXtJe5HRNkL+D2SWo0MpGqKHnfyj2n0GClc03
riypgEuUwz2jDjYqjcFkKDfeB3h2CM5qkB9UQY8lzJwDNcoFEMgo1Z4nxwpY+13YCUrwNxc91Clu
LOpPSGVQCOroIxWaDjYwmkLpz7I77pojFZgFrHs4Mi4zjkdu/DaDeM1gBSFOUUHyxFIFTogYiCQX
/VQ0P9PVXptJd02c7zV5PMjaVvCNCe+sfwmALXk0C+dfO1p9gNKS14dLcniQdAXxTleewGBQpI0l
g38ZLY5YxDqNaDZrF+dQwn5Urka0tw0oKz5i+iT5VMU2Q+09Nh481jnNnJbdw4JA/7nxFgUHksO8
vKu7YkzW0TEaewZD2nYfzBRoQgalkV6gw9rJumNrDILs8KO0nzD57mTdj3lx60SOlVI9ZXr/Vziw
n3MepoMCnUnE9s/aCUguzKcM9NfN1I1l5cntVs9IoDCrDE27wI7VsAnbrZ/qLd+Sy/PURQzVsgNA
icKijvHMr/FgVvOgGTXz4Sdl2nAEMnp0ERpaAwR5SAFFGvlJ9jAteZoV5v8XwJ6kmHgnm67bHxul
7kh+PLRbcBDVzbwOKMy6BvpdvNaZ2CaQOSfjvmdW9XOdhYXUB1G9zhJ2Akt5JzYoLxrsFqQ/Zb25
/TTbfZM+6IjekY3eI86TvhLgTNUJg+iucUQR/WKE56XD3LisPrcq94zwObs6WYhWZMtezTtXXvPw
fw88gEHApGAzS1U/z8C/UftzwW1dQUvLHD5YBC+vXB3fkKckN7/704z+Hx6L5mBYDWNJa7Vf1urq
hG2nlUU8KwikljlJDruZhr18RJ6fUVbAuYpu9YO4zQpz56UFsVqK5Fxt15xlKCGF/l2dn78ajp1W
O9c5KzN4S/avPuQBaioZEtLBXGGiKvwfB8nGHyxjzgNpr47INL/UStAAHBf5rx7qRpvyAx58xtdH
ozS1jDncKMKKYgOV77ZUxks8JCVbQnpIIqnHNgcK6WrA/TVxE7VVmDAM1xIPgeFNSBRGC4jaTFlj
/iAXh+RLDw5tNCzXl8yiexfTN5+vNb4lHFlnrzg4sscl3Cu6eoqKirDUpzBCBbeXQSaRJYGUJPvj
UkEGbBojRv1mnfRZLnwefZxsB4EHUg4mVeB2yk31UEt4xYnUT6D4RflKyG50GOQh/s21hnzz7L6p
3P/Ek7jpR2FW3uwpN0FIInIvNMEXP9GGPEXVnyALQSnFVA+b1GgA9uZK5FZUE97tyDaAJCIXKyrj
KY+8aandYRpcGmJ+XAdwYQUi3nS9SOiProQarpLy0//fv38VbAcNyhHMTR3UOhJn4Us+jg0h9Hdb
6sMSvQwCLa9/h5RbmotyiPVpzF7UYnrg6E95+iOrRSB5UkTELs5byX3xclDllkdheBHUQwaCplez
PBA8J8xHxez0oNntHd/7EPIzBtMmzi5RWgX2izTzZRmm/J3BoRzYhBsMgqP2nfBVMf5rkNhNfbBG
ghRetEme4hDtqpoJlkRjHdAHtkzgcBLxpH8kNHsa2mgqIacv7z9R1m8NJSI+VKaX16KgRJ+mlU8z
skRIqtSNk5jFrQVTfsC0JauWfjpSy/F3LbRY12cOMsgPiWDFKDgAuNXDvIQ0Z7fg0CmThZmPHXJ8
FOFvUhFM9RoUh+Sbkba9+Jo987Yfb676WZ+O2nB30gon1tmZc2k+0+Ui9cY6AAi8C/eCxvEi0FIR
5BbmTCT2cR7XP7xd37G9rlXuUaRInE9oRt0oweFzMtiZeSFybalR54LH+q2tzs+BGW3uTnka7C3Z
OFXA+PHAgwtpFxQLAo2seXHDGNjWUxksEhKXNa1M78HiHXE6Zmn9q6wqDRm9Un5ohvlE2YIeoKso
BmJB/+mRq49CYpZdW4ePmQLXjmW9+Jy/nCsbbI8inU7BBhlsqm/HZ2ihbG4dsEKjGoBrk4Bdshcz
GJN/QIKAqtCgnWgqhDTFG8wvGZd/vewtmNG40C7DqzgjTbIxV1gtZNglYaywdk2PsgrhQLMZ+zPy
qmHJFLXXctm3QkY58CUafeu3Guj7Gf3wMpmqZeB1stZMDYurcyy9Cq2w6+97XkJlaJJcjHcJk0gm
RtsYyCAmRq5Q8atynT7V0TTJ0vLEQ6h1UtJ4V78X8MaCLEXXWVnoySSGzXjcsBD6eTol+kZp1fdQ
sYaxzRe8xCwljYrZ7mbzvhR1yXg5mSKUgrDz5btpRO8z58lFcMwTDkJ8flkZaxtnozVeIVR5GJh8
g+9nvEDSZFRwVB15bsnvCVY6TJB2uEhFbdhqRbeobYhWT5v8+HN/PXiKNKt/C7i2sBmVtPVujCT/
qIXemOBB/dbbtD2Ghamstl61uJBmGQvN1aUWE8VZzj2v/m9tM+BdlIg3Mw6Gt+LjMvP+AmW4wN1t
LfJFQ5PV/BoPorhlpIntS9DDDT/HTujBeL9+SlsPTdR3cLnUvD0XCYpP/9yO1FwgCgBkNYR0aqiS
3D8HN3VcEj4W7NJ5z1RE5AoQ7HoNp/qe1FevZq0qPB0Laao7iVp9oZqkr2wbX7NKzGwMt8T9Ik0y
PudElMV+ILsCmPTiGb96nEJNa3wRUaYb4vgAw4g3Ww9yuw5C70djyxAa7lQkL39tZ6qYeK9dnoSy
mcxGnuUtf8orjUjONuNGLrqKg8rbi7iZyzdP6iW1srxEOJQNZRx/7PkgBgp7W9hDf8focNmIsEaR
/cu9lVme4mWeIaKPux3kqD8xxvCvEZhy8+OF5JhHsMBuqBUJTBPwYb6wbAzNNl8qEK5J/SouZcXt
Qhvm1ZghqN/eJbfYEcpKC4BwXfIphj0Y8p8XCfZkpQKtYOMoSQUUwPWk1wSYDYJs+xdBX3nv1E2I
yKzFPXAM+YOcl6iEu4ZrbOhF1HylF85f2XHqZ8cRe/xasfaJMAA0ZXJAWxz8PTK5jzfxT1aVlmvU
fbu8OnH6B0v+ypW7s88/ixSgalVLOUqc0p6OtNe6nvVDdkK4gkI5tNGgySS56q5A0jJzFpJ2WANA
nRu6jeif5XGugwZN7IzjdoDs8yzN2CKkWiBkMhQ3RFtpK6hDqoQ0Pus2/qctwnvU5HECoA6UAhne
/vrUI4xGlCSZi+F9CKmcdUyOcUG5i8bKx5YGVkYSblDzxp9StGa2gBCBQrs1rq33t4i14JQQGoSZ
ye5Vzkwn1zz96uscETD2ntXyDY/VI8f9pCLo/eQJL8EhJ5asaDKvDBTf0/PKRyLGmYZbov1hEDuf
Qyrc3vwitZONrV51asQxKNn2ykgPAP9iwO0DyPPZ9vHbacDmOfTn465TjO41+4/DUWZBAOiri6pv
MpHgD/C9Um8x3upscg/FuFjIDO6FB5Qnwx6WsflCBnoDn8J6PAMt65sPr/sVCv9yP7Tqox6JiYty
ywyT3Dnk6+5315aG5v+zgBHcspuyOhVVCQg8RAjO6njrxKIhSqGU2bZARmPyC1hgDa3TJjZ2xJ+P
CokqWlwbfGd8cGvB2DGow95RrvMBA/brNqk2SCoetFE/qPotgFCSV+NrlJhlHLDDEtsohHYzaJ5q
QMqf7kbD9A77LWLkkCgU7i308z5scMbzuhzQGvr04gtaL+nGda/j6HVwWWqH1ZqnbjQUwLsFGJrz
gt6V5FIixZda03WwGo4DpIKPukFuCkrxjTOYs+nSGo6zDx5IMa2UvAYmv2uDIOWEhylTGlMZ3C7C
jQOrmVoQ8me6x5HTPTqRd2cdktLKjFBURzxWqRhML9WXzY7DkJfy/dgUQtc/iJEXTASLRok27D1r
+RzwV6bbOihO9Rbscpq7FMXVu96mKU2IdIp8eXE7qqLsJlulGfKK48ZlcIgL+qtxqpEK8hIZi31I
Yt5qLCYiJMOpitb9C0hH3/OojgicKIzNxKI9+kf5K50w7edYkTh+rl8m9OErdP5U1XNGgRbkIyst
fto1NZ9jwvrVdPTdOv41hE090T3qOsvdnvEYR6PdE6IylVB/q89GyqbAvPGM1gqjyvCtJEOJgdo+
tEfXDcqpe5wdJiK5jfVBXPVqoswl8gaKqVBp5WoRBgWPKakhJsv9I74ZdC8q2hfXvd4BA/FJWP0J
StCg2aSxnX3QGvdlqj5S46dNb24bcE8x1owNqeGHfCPQ+BYk3ZCaN+r/cUlReakZhuZ0RfJtnPFu
hy06tJKzxdVU3+d7ShiCGuTMjGZP6atLZrpsDhZxYhc3ZHEkcVjiM7A8YecmKWlTMmV7LYYyGWhY
paET6iXitXZXifRoqadPpg4PBhaEwTybP4ZHVpAtMduvdkM1GuBcg7go8I6WMCyGI3zqUJVQ6RaW
G145+yFYSnuRIP+bpfYQGDjQacnK67gi8mgHwFxe/0dWVTa2VZoUQtd5no5Zns9/O2jCOThE6Mmb
UcIieojsHOVSN5mEo+K47K2wnu4FVu/BTTEFBE4lRC2NQ9tZA+pCOZj8h+71l2/jYhznYrnnL4K5
+GYnqhG5CgRbO4pqIXi9v3wLphQ/5l9fkRlCljfbpAxPHLb3wdSUfA/gI5/hjDRv8Qh4UgrwEbX/
FK25z2aTn2MYtK06s4jgzdf3ses0KJtLWfIFhRqUcJ0E1qvWAvFroD1ddlf+Nd28hhJRWyI6yncY
czAijkB2V+bohysdHBoXIHpE6NfSwh9+0oTIdLbdiv3oDsCHDzN389L6m+Punx8pS190yQ8BvUz+
j8ad3fgnbnwjLRHabqORJoeGSaLnAPl8g88EoJ4kBy582pIz0WYkBIbq1k0RRYtEYPXbAM63Z9tF
gt11mI3zZPU+ItNoGBlpnPcC48FUWuO214e6QhVqPEPPm8bMiEzpYnzd6iw4jMcet3hVyunUbGAq
KmF2cYOu5bdADk6H7Xj4p+x20qyqbihXcobNe/idRSR5/5GkYKBbjpRQAc3Da4meRtw70Onk4I7y
8VnaGY/ICB+X3idvsctowtnBuXBIPvHu5zDtJ3BE50t7BH1q/oNhgwN6vdtnJcB4ZLp/eBd4HuR4
uo6VfWjAyj+pZZ+JAfwrMyBXxzLYA/Sf0W0tuvHnHYyBuSQ/SpeulexE6EjnbAwNE9I7OezARn1n
KTKwGyGA78i7/k/qfjny+yI67ujtHOKCnVEun/44Icu8oCUT5CtIhDu2TV7+ndpWL2LS1PoILGbN
smtXTAROi/aPgk5mno1MDH4jl+p4EJg9DM2a91z3Xyy5eSRF7KPJpwcpbPdWidUh9ka/gIg9t+Uv
p/Yws2YA1SEQXUVILT2rtbGgIlUKkZswX4mMVvuIElN18ysBXbGOpHryP7kcTCYKJ9teBq6vk3Ky
nkDM6DskwJ2x750mvHmxL6CSz+gvmICuIvT/zZSdJqeJUUvYvpnab7PYcP/6z/olGkvn3kG7oQg2
nxVwk/FoUp98FVMO0cFPajbmQl2glofa4IesqwISe2ZZgph9pAl6Lal3WhVgw/RBitJjslKmrApD
4DdCUC3vjRdPxpzcfAp3+jxn3RP2NJmDJCnSfN3U67KtHxpibGTpQLCfKkJAGx2xeVGZCCx0dD/V
vyQ7LsYNq6g9gettsa3BH90GUdVlyupu5LdZekjOOs/81eeoTfraBklaYzsykhzUgiNDLHNGQ1fE
ON8lQN4lLCoJbj6NdmR/akUIyp/YHHSf6N56KqECAochjZPkwokQeVunjCFbNtkk4wZuSVwTiah+
kZlI8R6fUKqrJHatQ/3SQKtXx6jLJ1c5CtLrMtoaBWl9VqH8bWuTBevexkUTXNRgfd+ZeCjZd6F9
0lPy+AAaNUq/zFp9xQwOgb6Jas5Y2Mqin0ePDU4Kjih3yhWq2wA7/AcGvphcWEzbQWBi0q5tqrcb
hImw9kyoO9UwbsccCQWIlcwuwfALQTpuiKwSe04kLTp+Et5fgS+TY8rPTfj0IwMC5ZcWk/gOG9LV
A4vdZjFLM2Kd+7u4xytx2LiSafbqPKltEGqWWfD5sJ5ueLQ2m+hL5qrPwzkBpoLD0TlgnHHhNazl
s/pdw4Bve+xI7i65qN5ziEWrRtPVUCbDikLY9hxDg/137PmJvh3DPZfYoRy8xuebQRThqN1Jmvzn
fMoDtGAcjQiegFL0MLVtSU+yT55Bpbs5RTk954eyBwYu8ailB9cC76WMgZTXPoWBGnP2T7puKYgW
N60j8CMLuFyb4mgg5bpnSoCcXunKcAI9tCvSDdgHhfpSH1TcXISk53uD+nbSsSnVFnt6oL9sJUJI
GvBNcsgGyB6spUkuc2CAPXa+yF6yLzVC9SZa7VqbAemsHOeNoxGwrKr1xJkaqXq8IPfFUcTOF6oa
iY90fwj3kYBiGJb8boB7t41d6MV2EX5bS7gelJrPK8haOSstQUnxAXikRq36heXY5PZ4zOPtFOEC
6xkLyu5mgZ5sY37UZXDQ/IimSWiGDjeZBymVESh6dDVd479YnTBuiAT52Utr8sgFkgFqHB8thXA7
c7UCZH3+CxpFQ4psoJZDhWToV6F0Oh66lycJlAk027K8bCZkCPCdKfmF42a1coJT9w17MOdwcjNN
lf31KGFoPNaR7EuRhxx9D8hWSO4YI/XFU9AoxMowOvFNjVWfP1K0cHU09ZGCZsIeaSPmgd4a/fwH
0ROsQnq3gsCb7v6MKbw+AeHD2F5REozPMzBcJzCt8kAo/s7doTnFZGu2Ey4XBN+FYUq50cZ+uWjL
E29BUzpIdMd6vlrKzuCZdJ6RBLlgAXC4LmBorhi2YvTugNe6OKaLAzG0T1cRpfDVcFnsN0mSyRUm
XiohMC28xIXOLFw0xxr45pJmscny/j38nfHegplS1URwtb0IR+at9KjHP2gZVZWBL0N1hNLTD0TO
yW2ChjxLaeLqbJChv3DuGgNpLY5RgaezJQwuhgH5NGdGITvW2NZt8xYd1nBuiKZ6RMre6KKGaycX
bGFbEsyOvbK8ygmW6o1fugY2NKXGZKLf6n4S6eiMcF9NwYCequZoiONmywI2lLPy9n2DQzz5DHR9
8teqXWhAhFHiLROD4fHzKy18myYQRSBLItl6Frw4C9EIvVaPNvLweScrfCb4ws+KCdPKbIQfYOMu
r090hvCP34ybfvNTKUIjgEQzaiM7auLIzvMgut5AFIP8KZsDogZZi2upnk1AuxPrRdok/13au7iy
dJvpMJs7ycah/tzSmCZX8abgRZmYvzq4GSNvmEhQgPrgL8CVSVTf7VVN9bGcwi7HJ3ntAUFwF8zQ
fhimr7rr2fmfEM+c9DRlEorr5TDGJwBhsTFDad0cucX8v5++oLH4MLVQuJiTwwAMa3ZTHOBZOgqm
8ncKQZrJVo5mO8vgJ5ktQKQ24/XUZ5GpA30tM0oCZLyzCxDzVksyYxGliSc2/x6TEWLzLv4x0e23
VIpGxV+F63jWta4+AUKNLNwBcrFeLjskvCycleQ69veIthtJ5czEKEdqNoDzIqigK2IIsd8T38z0
YhGHIWFbqL1ho7iGil41U5aCWA/GucDvgNZ1Y5QwCauUl975XB+QtPh1bQ9Ja6jfH80rG4F7f7Aw
Pg1volDmlC0ycIWVayaqeQycFi9GTdVZK2/Okd0WEgomw6BOK1IIl6Dom7l9bAcY4Adcuz2XkSS4
pEEbLXS2fyAj+Oku7bZC554EQZByw568WS4qPy8sp1opUXZ4A9CvVGGXiY8IcV0IorKYQ3tl+Aeh
loSljzEjLofJHPN9Uz1FjZed2qmVdiq2d7OmuFEC/IydEyh93U3ER5YyUhAMr9NTD0U4/X7hrCBX
2QStJAm1GVdZ9sKMVuX6i8oVY9JC+9zvpVRk1TEqhXNxlarSiGkLB/6JpsUcNj/at8mwrTgNcEz1
BRGLQy0CuYPt3DNiTSgmkGKKeCjiwMLKTVPA1qQ01ag5qEMop4+C944h/F5LXrtEdbRHBPoB2r3n
A3QxcM52OFwnjQ3UfdIfuoHxKqVrR84m2Wi7u8E0r1AZ+V1sB/lFR1qeuNAApGy3EjP+iofFYCfX
1mtFYsFp2EVETjH9bSqbRwatPbTb9w7lj6RehMVTPSY/9G1CgIimKxOb+sXrqLPXeKnHOhcWtZub
7cOhmajgEcV/AeVfiYyCdTvQJk2XSu60pICCs8bU6Q7JISYp5z5zitYJtL7nc+B74NaXTwS5yjUp
vWy3/uyvDeX0x3oP8+YWdy/+vy64JNyl4drn1bPKF+1nO3SHcv/WKkgI81hJsalPgir5c9V83Q8i
cyjyT04HXTFnHnDQThw4D/4eEnFgvcSuef4LgZsSfnSdKfOO8B6aULxZfFXjiCd2gFtGRHONhQTG
dv7NsXPVR+02boyDKbn/MW4ANjhdHhCeRH8zYmY6i02/xapmbxzLhq/RVYFpnnjbMULNURF144G2
qGdDNx9kMTQ6qMi8PUWnyLm1Q0DBbmqwoO/Qy9zqWcP0cwnMY/kPTypTE7aZ0U5+ObwGkS0AM+4Y
j1w93pe6Y1wVlAVAgRNisgWDkR/kOJq1kiiIpHTpzslYf+u+78D8KAEEdGeEilkQgrzYq5FZjdbM
K9/xnMFi+8ho2JabyjmG8tU6S2uAoNC5qNiylM3sfPuhWQCuGZH5tzUKCqGKwWUMPuZAU9oE6dzc
N67PAsTbrbjoiBOi5B2LbEYHDEqhEuHGiwBHa7op6sFm7EifQ2UACNiFPaxX7k+6ajx3ORnDOH1w
1rSB4YMEUd1pnU6b8nVmiXx+GMwuQ6UUUeed8fiuCf3201VcLvL0S5bkZS/URQDeBhTuqDG7tEYR
g6I1pslNTrs53sqth49dqqkzT1C6UD2xGW+x+uMoGoGkm//FMFffUsx4K7uE+38R7JK7sTrs9Qmz
7ti7XFjujwyaDiDdqVmi1PzKFXVqMj0UBVD8m1OvuerlcMJ+k2J9DgHiITJh0Fo56iXI0JXL8Axl
kV2+9zWiX2/OAqLneNqUKAGHI4ny1WAd4EDt3ER5M9inVAac4+U0S/etDT5pLmf61rYmOvrtC9VK
Q6OX7yq8IpOeR6A1p+ed0cFaMGA2CVv6Z5sMM+krXyPXkQuBCuDq4xKRyuY3gGoEt5CDcE/DMLQ8
MHjGEtmDVfv2j8/mWmms/aw48x+Ct+UdM//GEYXmTWU3oXX3D8FUosfwWD67L6TxHFIijJzdhbro
BimoXXSAYULgfukc00pZNiczuL1ZKAXv+Qb+jvf8wdOUZwG1iVTMf2adAe5F7EohFRB2yeK4cTF6
kWTBFTlMxIKvuxrkX8EiCBJ/pYv6cmW+G/sRcL4ojdC6eieQHnUc9vEDc2TLytxHecZtSN/R5SUG
JsvFk9viH7TmeXqznqX26vtcOc054448DuTtdYFenfWLBPWLrxawO/I2kvlIQJVJ4ROi4qt/OGOI
e4W+5zNQ9+j/osA7dhX5It3z2d0szcejwsVQaZwJeZQT8+QQOYx3FImeNx+rutxoUCiB4Ra5T+nn
awpgfSTKX1vSE6YY3U+TBhOmVip0IBfyhijk029YlE/Y17oXMNsqj9setfZUwgo6V6+U2Fj5W0PM
NbePT1jX8ig3mZ7OSeyv3Oz9vqtysGZ2bEpiFbKUdCtEdIa6Ayd1XFaU8K98ZwWI3qhBkPcFYRjj
hVZBCT0aSNQfrbMYtv5LFoccXBeqSLnRpo3J2s9ZcEudAuzDN69nc+fdrliesH8VJ/8CclQt4JF0
zMoJCfZEHEwDsCgESMC9Nd/3WKA71FEZKKGQ4dvKdfWt0+SpkulVXM4YOry7HPoXM4XSjzKWO5UE
PPzJbnezZMpwvkr9rRd5xZqKNlVplKowMTurfCbxDPo4ADhBHZEzRiAnYGTk+d7qI1yxA0qOUyeE
jwfE3Rwe/Q8G6Ycz/Tkqm5hbbgWRxYr+5Y37mQZfj3ukej5t7dnID/eMB7AYEjgB2lMMql/30e8y
A9E5WKvnB7j5Z7KxuvDhHJVfGbK5t8F1EVzyr9BGru7gna9d4T2mbRymlPM/24jD1TfUh3xdm0YE
XOdGklHwJZ7svKqI7b5v/X14U3g6ZExMss1k8lEbC3sFikWLbn/gZxbJjXNEXthBv9ES2TJqKp4q
m4722PDcmNAOENM4lobFVlZiZGImoTpvUpCrqYQkof3oDXOQfDU2PBaO28UGqBIJ/sYcA3Ao5x87
/ZQ7XofcfxMdko1zVZvD3BD9rHX58JFJzt9ZhFYAcUwMNw2LLyMtNhIeHTvbXCVl1WgsWQsUqWx2
bAOUzIlM77N0CoC9iuPX41ZNcsgfIIYix4MJQ33Ccq9dH730zfGAJVw7882AaL2R2S266uNdNzX/
OFu47l5+X6X439fHLpKz1L/HNu/XN8i+QAQqFVU6x4unAWtq0Fcmm9ia7RY0FgytlqiI44pc0iVz
ZqRKW+R3qQaIIPkquRaMH9/Ua9qOi6+20MPsqgz7FFAzcaMY4kt1U5TqmLl5WztkTQ4qOMgKWH/7
AVww7w8BABWaYEBOtbSkri+d/KJzZsYMm15J88x9/nZxOllvn4eRwUemKrGb++DP5cy5K9QBpcEG
YEXRQX8kil44/t+FzZnV+J5SGeNbv65rX799TrKitCmsslCo4R+sRHpNgA3PfdRdd0RAHtMqeemT
oZOZQPTJ62wFNcdC9JqjaXhg957AACCq/qtRMMDcqnydEfpRoQ0LCSZepNkYswF5ASUtq/XxeZdz
gJ1TBkegnd5oLSQYVRYFFoSCrc/h0YRjIlAV7CRCAzpiouXpftZd+wFp0IHtv98yXAy4pQkrNmI8
1havtwJJZElhHPFv54pNBbGNJ12oMWlb00DV9Dj6WIQVT4kUcJjidwE9zlLD8ctgpqqK75ozbrn+
F7vThVNb1lqnp9EfXqx+DdFT/PzjH5JLzXuLLzCipWCht6UlS1NUcYxGTfRIZkuA7MYjUhEhLGyi
baU28KNZmag5bcdjCDBmidepYxCsmlX9iwjlXzW1EvL6LYmVcmJAufLVR3h04Ve2W8TdBzTPjRq5
6fWdIbYiNHU+i7OrtX3uUBeW4c0hm6ALEXSnqP5fh13SKOHliajLDgei9eIjpXUS74mkv3bBUoxc
FLBRER49+iPCCNfUA5bRH11VesA5ySW+djQjeufGY5FeIb+NfsbPTElKNJk1ik2rVoFaBDRcYJwq
G5OpS1I+l9jVnXGhsyjds8oI7GHhD0EbBithzMQ/tj1DLp1wbBKXGjztU5uAzOvsFSTcEb+2h92x
5doWyiMkxeUIFycRlfca/N3yQbS8EJKGG2j7RxBZPgb6M7GJzMr2IziwVqnjior4y19ogtjJEgUr
hNb1FdxpwVLQXS2MfJdKW6qYkcvixqu0gAUw9NQJskrkeAx5upOYNoYdoGfGfiPmR8Gy0bRGS64H
xCGiLTB23Tjbn09McMxL4tSv6fjyfT+/hNZBoAV1AHoD4wHPUYgvzn40qtJBzMYuZa9U/5YA9TP3
ZFpvZvv8rXU1B2bS5eU8uMva1fFHik53ggvapaY05kCkRXOKsr4B+KTM6kw4qd7rZ+w52eVmzZyM
pwmkR+z2rftsNABhsboGl5T9inc85683QBXgG3w6iQCmvl0NxXM9GiujhX4nnleAnfQdcUU8eCC5
+gazIqn8TCpslcOqFTDBRCbzn/MIbh7CyDm5Y5nzphq+QRcPE8vwFpnnO+O6Gwms4B3A5VnPthXm
2hXG3qP6yNWKqR7G8CMAXGrNIkIfYgcFH2B0r96MY8tMf9uPh31BscLsBo3bQenGXRfxbR0yMaNm
uV5bpIOKnAMfM57jUbQr+TY8sf84U2QB1oI18dwIw/+7Ap4/spG+72GoC1JfwIULfTK/Ri552oxu
JmYCpTDVDxI1o0CJRwzcSlic2yrKCfWUdLXdcU5TyiumRA3UFijJB08UelF2niuv37kKMCX+mjF8
9h5jEYvh+1WdZ0P9vdsxTXjTIuGgebXR35RINKVAfcqRyw0qy1NVZK4OAMshzbcM1YhmXrTzoDJO
71ylzI8K3XvzeX1wKdPXSXHf1fHXArbmVtyWXDWtTfwasrK3ENzMPHVPdVx4yC2HLuYUF4yRmIB9
gLE327BfcFspRQ4Czx3+TyLXce03FdAWheqWKOQ9LHYM0uGfjw9Wfktjd/7H4tXL1Ebpqv8uzRuq
BXGfX2XJiaaUYenXL4iH18AjCaJal+L8Q6d29pPbw6+IMMVnKkL9Ui6cBMsOZVDwrhZDSBg1nj0m
80YO+zz9/xJ4JVE1zCYwoHlXjRovorFxxd2ysJ4CoBKz3SZm7mQJVwLSTgyhqYynmb811QneN6WQ
qsAe+/ZqTuCjr9KUCR2K8KoKNtn+zeM0cgn/MSo0iDZ/ezn8lj/VA+N4OhtjGsD5YTScHx4xofQQ
IAGmQ28o1qNSxYwW9HpNFwi3wXDQ60f70BtQbw4pCFvt/YyUVaFcHZViSo6OwfJ5jz46h8WQoMak
vvVkAXtpC+8WuJH/sFqk9gZQeIaTly+0mTSWsY9alqx0Ix7xE4eYmmyRTwIAHxgkL9urgA7yGpRI
GkEsZrCzJGgRjpztswbQvDZDMlkvxDcCm1eJNW/SqPuGiX2aqaqBth/Y/p2OukX+3WqtBl5WEHLH
597I3eY1Gb4rRrYJb5c6OZ/RAtFpqOtkz+yCFcPT45NUwISjK4U94xXkQH00FOKzvIeyzAF26uVo
9X0pnKSsU+QYbxCjHu6qgjDpkBItB34i52G/dZhYLrkh++uN+B+Dlucw4ZH/y63jW4+5GmZfVn2u
l2cWddrOms3Qeb1XF1yN6bOspt/6uZsUx+Wq6bpaePhUAmVp9AltzxKPYbfp4on/r4RDkS4Q1Jvd
Cl7jX9Fzy3phcC7cro1W7H1O/Hy1tFizWQEGyHprebKaZRiqJb0tCCjL3sRMesvRlDg5wPTZ/ekB
pJ88yTC7yQxP94J4djFEyjvlujvc6bASIy/sp232SIj6qr76JLwnDyWKU/+fysLHC6/tyKPOYkcl
xePLrMdiTqEVHaD6BWLETjP7R28VwaPD++Vq6TEQHSWUASZwbb2mK1nqelirfWFOYtS1t3SAgUSG
zhdHH+pqmx3IJlS+LbLeOXE6xO3JnFBSISU+3YM9srSlyOrWP8hc1KENkotdVpTcmDHDIpPBjuMS
SNdfmbM0qz+c7HCTsq4Iqds8vTEup/KX9iRXO8BAvvzxZesVY0st8Smn0Q8zbNh6/i/qMD4O3PCw
BghogxcJ6XrZO6xi+CTcESBHY7+e/DjaGqkxzITA9QPIxLnUC0Gw7Z0hsunBNtSdG6JKUi7u6Vmm
dJRePimBPVX6kWwVwpY/DK25L+/0ygtJzwVD/m6gHQ21ToycOFarRaY5NKnFF4quHP1PUzHOXk83
Bo3S52qvzA5lSx//7mKDAhtBFlEEy1H/K9cfZVn4h8ngwRyLtCGPHGGN01ExnYdO4Tyu4eJye8Jr
d2IrI+v6grBwQNx518RINGzz0ddlQn0La9so9iPS6KQTaoEPntpjKBKb41H1aWWZClPGSIjQxZRY
jchdOxI4JdOntZqW2C5n/N5bdZBDSOQ3DAG8BuNtjnC0MoPESgy0jgbQkZRYCkhIhaOURi4bowh2
1sncCN4NPqbu6L3lNdwaeEFIsEvdLkjYW90qH5m0zq70p4IizH+WGwWjnKFFWw2AW9m12Q6VPfFq
wRjkKJvLrzH93QJiezssgmcVX+z/ogAR3Y6k0XQB3NxGtNzu4ATuGzumIl94EOzypCkzCzU/54m/
glwLH9rQU80MJ2IuTIx1EdfZkyyTui/nm4xChA2YOrDon9NTsVK2XTaOf4toIwUQiZhhy0TrJfF3
e9G4VdSo/gJ2RONd2Jsxsj83OIvCHjs9blK/E2ZnYk7iP4uEgfwLLGthMf+VMsD7+wuvCrewE8wt
MG7wXak/idgyaTPOgaloFebDJt7tHVZGvOUrwh91j2/ypi7LMyrVu2v9Qt3b3dgOY0G12oyTj+M8
E+opO0+6EeIRsQ6AyJiqehfNtR/JSqT9uI+kUZRAQKug3zvaXm47oKVxOLpO2eK41/rFyH9twrhb
qtWW5IpDFT249fHfbUvSwtytp38Zsb0F0pYlATyfBSjMFyPWnnNh7d8TGROhxj+KcXDQiZJbsTpR
///yp4yNP/6SQhPz0U7VZrpGwt70SSPelnJZGDMdSRdh287uuurtoKl4RETu88ud9JiWDGn1HgEN
g+kAmJQr8YlUgKYkt6cuEh+At+WH7gx2aXgxdDzzB6Slq+Uo6ea/HgVxT+UN9E3sygspuAO5/B1u
quB3BaiP4LJ0j76o55ZMrdPOaBT9bPjra/o5HW5t7WVhUPomJOXVuKsZ1ZK7/dDtQhr9ATdu0Ob5
87SH97FTxdi1FZfRURhc7fgvEqEZ83DqDmga0mnwB6NcSSnA7TxdCfHI253vNhhd8EQYwzPgq1dA
aRbyd2yOrdoOZGW4YFvtRzBcCt7DUbr8S7U4c3Ax9Vjpq0e+HQdYbiZr53RJI4yyPM1pM4KhDnib
YES4j3d2LGkE/JeYzzEPvzfncyVczXBVLBhN8X/bqlNPbcntRqLmAhHuoz+CXYrkyCLO+rpMrrnX
wp8qGjJnGDQoU8SFi0wlheuznhrwmdV7974LEXH01QoeKeUsi3crsYf0DGPzNndaZnbORqpJzaWh
q5TQS6XNdHua/Igm47tLcpOqHiDQALSqAGkjR0sXvPwXIIXDG4EDw8ejZHMpqUqQmND0zyVg3csW
7N9CDkbE00Cq7lc7D1luiik0KPY+KfC4FrTZo7HuU2/gRkVVNayXmn+2c+v/xh3fRukXJE0QcTuS
OZT8UWrqRjxHcBu4xG1L1Yys9StsptlOyX76RH4z99kCmbpc06URXoFXoiiEgKUiCrQ4soXbmYGS
IqIb22aFMlhsl42qm6tMR0eunP4raH3Fs7g4qQQ9A0Rqhe/4xt0mqGbxdFVFpyIB8fJ7XxFd8Vcz
K0L8kokUNrp3U0QJsyCu7LFkY525Zb3IVLmgzGdiGvRpbOFGOESEVmiuAfueyAoBXuKD6fW86nX0
7i/CbnssUsQg4oWMrxh1L4IoDQU3PxzCeFovmt+bpVVPb2gM2aVaB9k024BYmn6z5YpjjKyjfPH3
IsU5vqy5qetakVTLrgUBKIMjzf8e9Wr9nfMGu4srwKGGBmBphSt0cXsgpGf5/dJvIwW0ySA/G348
XtEy+rccwaASa45TRHwxaRxX9yS5RdURHVVTXraUCZvK4hPYy7tubcCaCfgACkKTtZ/EuMZ8JEJh
LEfZnDVkU989dKCo3vR62oPeR7B3BOAuju39rpztoZlTe/MdjLZmhAOUn1uOvj9pcEqy8CheuVcq
UblGXA96F8Gm2c9S+1nRLbv3An7xJKsHjCj+wlTmmkX/e306EuLsg2CI0eU2J76ZbPvFrJEIvFPx
nRyBkjj/ZKFmVcEjTKtAhbpsHKlfBs9/aL4hd4iBIiJ9ogfNeyMmVCLwTVxdwQhxvDDJbNsGy727
Q6xjYXz2mKAn/aDbNv+ESGZLUidyjoqoLAlu6SaETdvFBZEsJ7/wDFkQ1AFPyZ/FrY65R0oQjA5m
JSKOZuBjIsLHHjZzrLU37F/ESp79tXTCtNmz7pDot/1JV7nKnvKztJAwFFS2mjJy1L/esbvmAy59
CBI/U3Y0QmKPRWUY79NN/akox5SGRr2itW/S0odjsYJwxwnczVe3NwYuMiVBhYQI6UQjiSiBs/ET
uw7jQ+mmXS+miVozbZbgmqNTCWfnViCIh1CNIqRvu9/uA0Zn0DbxWntexloc/faxk1BXXQOedDbF
Znzad0GL2ls+pRNRW8VsDeIU+K6ePSCmvwjtA86zlNg/ldSnqodi46C4WnsyKbfjIpFg2O85Ny0r
37w0O2AjnQ43iKidF82VGyp/KWn+Xhm69v5RGODEg7Ff9f5J9H/tys/puLf5Fnag51PIkyKV4rFm
b7m+iBQI0f9QuvjhK81FoGbi+vbcb8lWGA5A8qvzcmazYkj+tV9RU9Y4eVOYhhJkJ2rVAnIoETi9
rnve9irYQpMLW5YNguLcpGT61CaIRQXmHrL8012EThvpoeab25Rk4981u7hjwctGF1uyJkpI9IfZ
4+KqEIF6hXm2911o3j7yrC4whWMHZXIVO0T4P63f72NE8spKn8WrDfx5qeSCwDarrMX2LfxmsnCk
HZjmV83lqgXxxXlHUS/zIBSdMfs2N+4WcvS+VFcBXgBxNGuG9jrTOuQMQxM3ijX82gShUpUVvayI
MsWh5i2BOuSWjT4vAMNa9duVoBnSg98UD495XOvuvaQ8sQFyGQuGY2sF1DeNBCfhrUqV8kpifhSp
fpbMQK4mhjPKyseb8Vn5PAQDB6WUQit9tqI78VgVI8BhOQOlTH0uLKAHxsBqVjmXEJgOqN9t9N5q
F9L1o1TIDabjrk/nSZiKNeIBpQiormwvT5m+WI2BS4ZaKSF/YdgHW4X4zrIEBtsAD5yTtEqkGP+x
nc692NDy++0LR54l9EBb03Robeed36z9je+bilvi834AIoe0iXTd9KN9dlOMV+QtaSQ9mQcaDizm
fkF87Svv17kAib+s90iazDWvPk766iXXcI5kgjuAjq0lkAV2m+QGDn5+4kjsryVq3O+Y4eqdf+Ci
VFS44Sl3UGOevESygY30hP8JVT1XDvE9bY3/Ot9aWSG/YAA3uDINIDEvZN/5SgBmrJtFPqqE1ia5
+WecQDYPuJTIZsxpfDYXgTN9RjRL8DuhFsOqR1enJCxPhkCJqilDrB29n9lQgBEo1nzm2Kns+h04
IKOh9iFRWkJUvkADqQpF4FTxTSNWyQxYrmPHofsDIcONvkudpdVygwG0MPf6QBVETNDMtQO40Xlg
gz5J9SQC70aaNVw4shDL4zjvvQGfpi0XEZF+okVZtAdL47L4z/P2z9dffusrNwjvDTCstD+CSFLt
TJvwJH5IVXs5JcWb+hMqULW2IZ/blHinGeHykLsTGXUJxwcDXqniZjLnplOKFm8BMOH6ZwnuuEj8
U0yX9qtvXXX1lEP+n1zxyfF9DNsmVgFZbEQuvlCdeSk4xAGd1HlAE1wc6u0zb8Oua6Ghw+9AbluZ
d29uLVy8nm0PrDwCNpvIozCVTkESI6oPcOaXGE/mIh1QPIOFbJ8oJz6puQourpzoRyCq5k8lL/kk
mPCztyyvVIL+ZBODiTmvK4XavsK8CoKMoWMfM9Fl7B0cgeQe0VBDJcPAZ+wGFs603EXbhy6zWnvL
gAcChOLB/mzWyoBvA0SPTqJJvLojrIy3wSia51RYKjLh7bvy0JUvZyoHzdkgS7wbak4fi6KTAb8T
bqvMIh4l2Np7EYCY1imBqe2/kN2ifYo913oSvzpygiHfNYZYthvErYzklqJpXVD/yEK+JsT5+mEV
NFLNxSHpfD2jliGvSpNJW/Og/clNw15H23cZyFCkvh8gcBK5A/gY1xri0IbtSUNqiHN73NJpVsdn
ABMCyzokhbNTVLxYav/Af7oDGJCm1gDrl1GmjVAgyp5jh/nDs9BSGBbgheZ2aNw8S2RAGpqlxaau
ancaLB9sO97YbYXEdSvRVHvRkXHXwEYOjHvG/VlZw48mNeQb+TuiAsAOkMlimlGmqNaxEu06TwHM
sY7ggemZGI4Qn05KC5XZsUTA1JdpKFvee2iE3AI/ORYqzeQX+C3tPwD+LatrMUpLuCEC0ASZnZO+
TiupZfTS2x9dEMOKj49Ienu/JJSW4pR6UdEnf4IYb0+BnxJfIjMJMXI2kGxWYmC1ZssmETLyAUGl
JIF9OMZBk7Z0J5/XYbSwGUaDo91mGlFjBXtU66Omvsp7zuz3u0NtaWthxtJiqg67WJhV56O55ws/
Pje+R4X0VZgSGBxl8dAC6QNpexo+/xQCS8XoEnmAvtNPiqigl0SC/C44h1yTsySLc4WowBKL2x53
SXVkmzwX+hoRoh6ElPCId3cryeQmyT+d/Vmdx4CR/0RbIYe79zK7dBA3LdAICsxtlM0CLQBAPCJQ
Pjw5DaXKYBWPzH8HDgwEL0cfVUkMqt4FgRiXLeLnuAug9ijBtpTTMwoUBJ4c1/R+sFiszHjzusg1
8QXYRFodulqwIQvgN49y7cFbdNZQgRHV8uNE7i5kiqIYTiY4VLVRTWhVrm0Rbntcvay9M2WqoAyv
3TH1DfWbIOt1TLMWdmxUr3M5kbx/4xoQW4Wu1ViiHO8nDyMWCqe/Qh9WIVBTORHIcRldBwVL81S3
+Q6mR+yScEf+7aizWsxpIpucej9OGVmoyfxrUQFIRF+MetYPtlkWyJJi4xi4MKzQYCuqcGfne8rN
FayEYsTF2g2PldtXsL4KLvCeL9tkzfQuHv3VFP5W/Z+rsWrhYm03vYFJeC73bxCKzAN9OSpKDry2
L5lTHtgrLeL2qFhwSC6tjqnnPvobBlkYcdjdWMYVeXWOOela+5mEeslBkxcXt9Yg4f7CkaBhvWwg
+x3l8+D2Dn7ExX31Z/ydkZNOHMbd29vWSvrP10WcjKu3o53wrJskty5GSKNdAJkEQ29KMK6rCC5s
l93qT0Abpo99wCXkf0aA4lS+aw/DG7UjU9xWq+zlgH+AT7MnL7mwKppMw+E/xicFfAr9948n6yzF
pv9AASgF/Xol+U3bQNa3R5VyMj5W6Uiv1xOFqo4f8+YUuvYF3LE7OuzSthxye8w71iqJNdLS+S+E
t5zFdSzbD7ffdc6YhaHTvinyQqZ6UrEK89Nm7iqEfIqDOq1XpC3XAnwOoQoVBVzU6/9qvhSejNam
/1V6B++3ODSz0q/R15C2CFW0AoOxtehYjrs3anXdr8Xv+bH5rpBipnG8+yE1Hy0Vj7/MHMebaa/p
NyZg926WVb67Pw2IONMdUAMk3bgdnZSrjX8FRJTzwTiO7p/uGnL0FSTNhFLH2/kE0OKDK4ILozs0
OG3qpHjrjxJCbyctWRlKmmK+qXa5lB8HA9ySxnNtC0+LkbfCcO4wMMvWjZwyWIBAvsTJfynl8rEg
3btrCrkPSQUDnvw4mSH70gfTcmcwhABJ2AXFwI28PZD5BWqMa6vd+b2oPd2zrU3l9ttn7spK2l29
xw1Vrjhzwdq0C95baIcl+Xh7hriE7+kf91/+faG9koxGxQRaxKQxSz7D4VyFMyET5Q9RPrnTyS4L
7IgZHEZbF/jhYYSeCZTIYKrWwPNd7MU4QyLz6ZHp7mJlTG21ar/G+gtDg8uFT2bDJiAxbWQtw883
gqLcf7ixM63luwx4AaHrl0qiH3lPMo1S1Tgfa4ObuoLGwVjavUH3y6AZezT1g33fox1TsqnhhXRc
25gE4b6OD47q40mfqrkRFppXFh7qyd30e948zuEz0JVBY+jVCA4NODbD0raKrf4gDU6tD4L1JV9j
ajwqP3t+uZhIQwwDK7477DkrltbncBK9iZMB6iErCSOVfPgc369vrLvbsG/67TQAvebI9/Dhj3gt
c8Jj5Ee72JUFUS4+FjlUy4rR39xzXPXujXi3JrBnmTkFXqebmJglTqr5vwtlVRwbr1RKQO4Pii2+
rOLXj9G9FW8HwLqf9pIcLHK10H6t/O+e7v/fpdF5VlDJpQUK+BQzXzVFXXTB//HthnLOadH6souM
QgYPZufiaqbQ+3Gvf6phKmdC/KIfWZ0+zk5D/KIwaFhLiSgvqbiHivIMrkaWD5mrtN/MT692uj5k
tfT/K3zCHKIdyCTG2TLTeF7z+yTl2agFzwcDNgAzsWWYwUo3vHwJfiS7/mCUqMgZiXpcjorEnr3G
/XAM9+yuSP1tJ4HVdtWoACFW3tMMG7HDdHJ4XQUffLxU8PISXA91Me+pg4/7LIUjFXLcMBSFzuTQ
aljhj38vq3EyWkMZHzoke3G14GO6hMsWimyBrrXkd22hIIHpyR+Ul4v4nVgRMSiZ8TRzunWU1vJn
9wHQKUWsz7C2eWL7gRGDRgZ9N/Qvwii2hkdXIdV5aFbRITvINzOfiOeGGmP/jXrpRxbJeMHG0aGW
WInjWUKvKxZRtqYrvgomXqFRpX4EFG36SyLG8n+S3nlo9OUswOLBt5bQHRVmSxV/S/6HsiDo/83A
A94ebvErC4jXu01RvJd/1YXlyZcVTwgpMeKtFkOViVDBewKXK/uPw0Y/OhXE9RCTKLYoHh1Dmar9
Z8ScFcBfXQHvb8pFMuzOu1+mb31HfzguFBHgT656IEdyGJzkRXwRq+6V6qC8kUfvrotUnnTey23m
El1sg7vSZvHr7liwhVhEOi/ORsGQsXPyWQxju+Mp+qaRzqQF6oQdZ17Rh8N471E0/DIngMcLNrCE
mLeBBPGpuQvPp6rPNy9HnjLlEbB+XHVNkgByMnovS1dRhTSDDwkdkplIRoyr7EKCfeCmvpym4hxA
kdPEvo57xbs1dJBNVXy5yt7bhrNjo4yVmtc7Uj/S4udjEOb++DMdj+nubOx3h5xobQfQPCFjN4pO
TsaeE8FkKa1M4dB5qhmn+VfjtoYtO6xxRSWFqmHAR25hTI8fNDHlHMSAFCUW+Sw8rC+UjQS//Rak
RGOWggWN6fkv0uaG3+blirlREG6/xL+JYi8Gsa+XWXl1xOqFvJ816QvYlEimTiulNrkIjpCFTLVL
wv9fpj/CNNTjdTAxruRl1U6HRgogY52SpCNPTC/j/jXEObClR1mXT10E452sGiZN+XeMm1CIW5FQ
9exK2oqWGbjQSLWXAww1wa6qCXHmQJ+Z/jie6OwiaEB8XLu5NNFRHvumzFlIS/HbIdEhfuG7OArE
56wkZwg7ecQvNOgLjd+DmSTjf8UHWCE9TEogbElWGppoXhMFLYhu05WGQs6UiC8szxyXgVYqEh69
paHl+8wP2piVuX2G9Wits4AQcAxYKaazQU7HQkZGu+sa5Q1Kdo0AN7GyMFfEqIPyVOzkv6RaN3v6
dthTX8YwwE3uEGMcU/9flbtL8gjhcJNlz/LZ9brpaUYO58vVzuAR43lxuf8s0Abt0b+ZWzt7Q6F4
o00x6soVp4p2yGBDAxsVltVvtB8x9zuHQKn8H3l2VusW2/mT4Ar6aqwRkaAp9cmVhd6qLTm0nYz1
mlHQ2i5yMUFBBjOsWJFigcRqn2mnYaOsaLVipFFVG9DER0Sg6W9RCxAkf4Y68b0zROtKosv72t5K
/eR0QtWWbb10VDfnjGRGOv27jMeddiW9w62nTKQ8jMgOk37Ts+5PbeCpYF5Szwc7i3eKRQqts4Ei
3p2OV6BT0jFJhNc7DXHUulsVoysHoEVJycLy6e0/aDUBIwZhXYICPNc65JYY5RYXpP2udT86U+7C
Sy2dvxoMCkI0xIhhhAy1856PPvDll5umJl6aqL8e7xSe6NG2N4LfuFXP51UrMG0CFcwID+tE3SNj
EPqgqyjriHRJ3WDb3SLz6J/hHm6DS0vgJDonRB5zpRG8s6he5gyDUkwfXrA4teEUOwN2Zq5oznrA
VSmQUrkf+7UNlme1gVCK+Jooy0s6IX8hYV9uKVx5YhjRIQTfY+05cwP1bQryqLyDmuYygm3slwIS
QCvJXpuxz7sddz8HbRCYpglS3HNAS4e7xYLf14+U2HqsKf6l8ZRJXBZ/2M7EnX1qt0sD+tSf57FV
vEHlPpFS2EuUovQX1d3eyXfpWJdpD44kXQYLMhO3O+B/hshbMrs9jfFQi1HBmHjCGe87pppvor6Q
A+FxGLcyyAiCqbFw7+A2qDyeSy2kb3Om4LKQdLOSv7XJL0RcUZY6lCd+N1HuntlBuRTk4UBtoLN9
aPAD10bWvJFz7AUOeyUasB++fXrU6SDuh08oZcGvLSWip+hV1oBUVkyQ2iusooMiGsz9ii4F1D+B
E/xZV4v+q1lS24eWmPgC2T22M2dP03ewROF5KT/gQYvVSrTmKaZ7tpM7k0DqX85dlw4cl/rB+i98
NbXr1kegMOmYCQ9Cp5dM3etxIaempqmlpbZf0kWn64xYMKra7RbmP1chssB2kh9hRCCb2V7h5KgH
/0UhjhY0NjQSK2hnJTWJVLzwhNbXaEvJE6NpP4v4uaJW/aWv3WKfYWRqcVvVs2SGEewQLx2juyKS
fn8WJitqVDr2tQ9Hk8gNsYT0i/Na+YUDezLf7PysYfKoeR71mCRHNglIBcm/0+zZWmW+F4goUDvJ
CLpC82AFesVA6nVUmZWCxHocHTQylXByIKwvChQ6lWCSd7oDEjPhU0jVmLlyuQ5zk14pUrSWYNCm
FRBp1EIjH9v4k0JklAzmBsmsky+DCpDjUDgA6CPj6S61d9m5z6u5B/+JN9K0Fkf+8sxXYX6DhVMg
VqBbhn+oycgGLYcG9d/c/XO/UXnxDsb77ni+q2YaiOdUZ/TnkKGV4kuk6+VxiOl1+1Ll9GpMoXm+
W2QbdPvDFUrmbTEPiOsPRAIpFqgmJSIIxq7vQ+f3RJJwiPcBtz8ntv5MOcydwqzBSpmnfemq+HeC
0lsFJ+jquUaObGf1PFtjPMNuUVucGYUv8pkgaGl+N2iy+q9YqER90Qr5BFZHFcjmCVeDFzh+ZoLD
Cyc099HwgK8fWy8Cc7rPoTyob/R2wUsLcX7Plrt54AGBx2aKXR6pBde8kR7vwZbQrsxGh6rylJyL
n6d4DFRrnACa66Tgue32f6zGdAlDJcJaFgUq9mtnK9GETFD0JTVWsWeVfr8jL8YUtM+K0jbouTAv
9YMStw/FHlypkP8HXrQxJd/ZzOUy5h6wERhAHUJ2d+jh/PGMHdcGb1M0dYlqANwVGvDMnkWF18P1
JEyUCBsPyXwZNpWCg5Y311hHcsD0ezWADekbBtE/Yv1vF21gVWBOcsdM2H23r4Ql3UaYTKICZC6W
DoPMWWmzGHy9y4JJe2yW4Ghft0lUa/zkYp9WBjPB8W0Bl2T7+80xeFq974vzZO9tMKmZVQl8vysM
Kx65/G0D1RqCPDADr2CU9ClsQfKZUNWsqX32O1UKS2u7abMF3kdbGwIf6Ofan2P3Y2m5+8EJb1o/
JmRtLB/bD5Hwzhgvqxqx0beLxnw7CCBRQjAiEoj2DO7hI2u1Jsye9Y/dQUF5AQ6MeRccZvpGplpB
FLcMHfJClQeRsKU6eZkJ6RvU5RwccG9Gybx0TP7vY0XpyduPs3/Nm0h5B1TxtSybIY3e0tNs2ZN3
GQ2LuGpndLGIqElmgslOoFbXQGYI2nlhiQW5lqL1RT8QNp/Z/j9wa2EdU+nsfqq31ETQMgitX8on
wmTKxm+nafPrgM/w8bgujGT759+hmSNGLaiLsedGL7ViDf/hxYE/U9gD4QSRDaGeK12sPCITxrjJ
8NrIJ+IO5yf/REStBnuFcspKdWIZF+faLW+yFxGi+Rn58UeLSlLZUr8v2mI5UH4NVofcOKMC3Lrk
7uXVzApOVDdPcysco0sqSxv6gnqnYVHwq2xN8Vg57LfPgRGxY1HrqmZRgpphhVUIQDQpqN1EAu0P
EQiqQqjj7R60UdTMgcAOv6Q/YK/dAlYQJ2v3L7wT8BIN91bjOE2GvxBaFwNpoCDqtnM3Gtbhmh0w
eBxni3SzD+6pAXmNWp9hF9QSkvYOG2pdS6AE1Ey/oZBznPs9GzB3ueFL2cZY2UYHnCiPdWXn3Let
3XVtem+FZCu37uC2p0/bPQWl7wd1TEiHyk7XTsNQ1UVI4Rtxgm7Ybjz+iOLjO7NR307xqSBalaJD
pzKCRIScAbz0TjUmxmzZ2/+VODsanfKACcakZ3mTXPGY2XkbH2FACSk3kVHu9A3I8kkON2FFnLAl
UZCMQf4bGfYiekMt6ROKiIm4AkMxb0sDhsu2tn2qOyz3/0fJEO/LksjFcidUY1ri6Gc1sFFbX/3a
HnKxtzl5GpGMouJegpBp3h7BlvljnXrHnR1jd21IUzAeTIIgbIiGwCPnc4I9p9e55gl3BVAxZJLA
Kc+77Bxt0XNog1ASWl3r1TgRRE8JJYQWxxI+uM1M60YvgDlTs0gwweMShtc40QtLciTtH3OYMkBM
pf3q3ejeZjwZqCGuFGA2EJt3Cvr1B4VHH/cEakYHzmrMYmYMvmGyTz6g7W9pN32q4uwsdyJ35X7k
OwVPjzL4uEpmk7apaC5ZMN0q2JkQBU3fMwXnOmmJdjQg4ahFHlow/cI3xVpVbNvB5oJILDiX51bd
HdFEeP85DjiDB/PyCRpeuBeu3FbaE+dg7GrQVacFbj3OAJIS99ioaTQL3nUARVwx6NJ/n4uJ4iSq
ezcGcCzaLd2JesgjOjpbdQyxPgG0/5KfE5ZUMOFuFGAkOThvnLsIFLpz3O4xNp75xMxWeTWhxkSp
2daH6Q7sgPriarvGJoKrbyfHP4hay4i30QK50IwP8LOJb9aJlgXUWDbCm4oLSzK+MK0gO8oc86bZ
i5nFCEAU/7T8eeNGSzVsSiJIqi0af6Buzf6t+oV384pQUD3PoHmdkx5B9Ym9OIJMNdOxzLMREPhd
tIbomaolEa69e+w+aCq0nH+LFYUF243CDN0KZHQl53sXdIzVGMqVcUK97UqYz8mI5IZXuMwV4yL4
XOOfHtBySeFuAK5PJVanyhVbgUodT/aKqU7D8VPXpv579zhh7VMqstB+oujhY86Mfryd4kYBmZ5D
R5cW8i+onKJbof+H4qxHRKN0PeTpalkBgOX6bF3oYp50mDp83nntAKj4FKZAqPUFv5LNSEHmkUX+
P6R1Uv6aDszNfWLCMZKXIWZH/W+t3inttba3W6r1Wo9Ks6FAmVUUi6EInWyF28Al6LcOXBIWEA/y
bUkrssdS0tUN7KoDXH7on7a4nSquba9bQVnYIIz8fB0EvoCAJuzJH5fUZosHb1s9t8XSreEqpT0z
hASRs37yWRjWtWJwPIOIsu0dhLmVEFVLoypOM3ynBxgrF/PYiXF4g369r3asklxzeCJCrRGVuBuq
bGOstSh6a6OIYGOuND9wfh007quJYEMfhpkx3a3Bvud2EqLuiVZYJ1z5p2sExsx0oewnr1I709U3
Uo5lsm4SWla7SyVlnisH9/c7a/0cC7F8ktpPL4RAzzsXHheZU3KT02SiSeKECkVEOpLNMDcISAhy
i655Wyk4IUbpiStH/SMc9TVZtajaBKyXD7Tu6SRI1o4gFzuLSE33Zev3ZOMUnkLO/Q0d/1bIU/oR
/PA1s8Z/q7kpoerLfIu7tds67Y3PKcl8O9b7mPQ7LWyKA4kp3yyZtc20dv4qlZvsWVnfAPvde7u6
TUhsRSSz23GiQMVROG5S7LJdjtep+rOYCrBA281OC3pHLVhuzqAm5JTGcmWyz6aE+7Z44Vt0iyBn
Ts0XJHM14hx+nhJarIGPq2p4u5uHnMXH02wp3J2K+8RBZOVCAMpyhQZy9TKGTM9ZGi+PsJFv9V68
bUrsxB2XHpG0foV9rRXZyp+nBVYJu8pQbQrs3/R+CoAcegfSERC1lqwIrzvghkj3iRYlehDcM7NN
3+r+5kbHvyi21ZSRZ9+tDJo4hOqpVWS/h+ybmmg47lZyVfAVzBWlL/JZEFv1vPs+bmyXgYme/z/6
hO2y9f3NODPoLJINO+x30qj0b6F9RZCJWZIvX3x8LOv5wf8DaV7GEoy3RsrmWu78lRwBUpbQXktV
tyLUxqt1RfpndjLCbn/v5igXCTpS6db86OZLK6GY+/Qw+USjEGrYU1ZDG3UEESw9zKSiGWOHsl+X
CC2JMuJaShqEJipPlTNZtpb+kJNSbZoGwaAd2EJnUPLBZSHRxOGSLDW7UJs41E8S1zUaB10AwW6X
4fYLInusGlXRh4k0dlEZf1ju54HAFULetWEbagiP8EFHvwUU2SIRGeMZ4QHf9n4vF2ibNeZxKm5y
vbDUm9TS9OZJUN/HV2hTSGU3zZjEYnd2nJ6xTYNkmCrqujOSvcizJqC0cyKICJy2Wbh0canpHI9o
Oq+OK6Kj16xjE/UF/7uPdlgIQHjxHG4k51pAI7Hz5UVUInnTqHZw8GvcSkjh45OLyIF9nap/w+UE
+e9y3J/hlCgXx0fhJco/Q3IISyDosGbJCDX341jvHSHL3BS78tYh4ECY0s6EuRW3BsSByVxxZnaJ
tyeSNagJFlr4mJzBKkekC0tH0yenrncVF2uwsvAdUwYi5LaQRi9wvF7+KIo3FrRdShg2pbNwGwez
u+n62XJ4MCIk41iwSJZ/Lu0vUk5J87B9x9ZPKbttlMIxP+uj7BdbT93gwhGqpcvTheLr7ZRTdWo2
6CqtS8iqCsASHl58V3sEFtQ41kNrqu2+JQALVaBIJnN5w3xKuwL0gX+LcJ6V356n8ZE082VCbvRT
BEdxz/TSv38AYa1QLK0Bw7ZobWuppb2R0wg6j5rsv9cr0DH8kMlg+7tXDdIpB6Na5jqiCPqAdmic
9qFjoDA8I7KivbbBSsHCVAodjMbtGEqMZ0a1bCjpRSw5ZvZeLUU+LMcbM8jp4D1TruVvOry+6Rbn
i47t3tLageGfT9odS2jrd7eqybD0B3mDgQRnvdfzr6tENhQ11p+dlIilqe/5Bav2tMrURue0etAO
+vvkJMQ1S2P1rsPtDUF5jwrwphrZGSfohJvRblwuIKC049dhgL5VKdaIsbV8bbDeYKg36aLTeDJl
U5M9GLCIVYLz+N3uxzzT7diQW7pdonlQixRyyd2Vs08ReA8+IsfiGyKKYOvYyybUGMs8BYfRm8Qe
CLDIAQWh/eP/QHVFWAO8dn8U9AL2Dd1dyupb2LnigeAoRcErL79vGqz768YFulUTnDBvW/IqBcLb
rC/vSIDJ8E3Q897y5LnOeiifNSecyf+CKtxpMj2ra/hOInupWoNQr3KZK8NwOx5dHTxhxbGuTgcb
bUJ2sL5865hhVA8qr3mDKQatmjY9JGEz9LvvWvikMvc9f+RZ2RcsOZhXzQpVGIms6U0yoNY5Trrj
mZyHg7m0irVRi0lxBFUO35/UhGeATyppkiUdebV5LRJmp8bebF2Z26JqTSaOPCFVIPc1WIckm2Rn
3yy3PI6OwkCuVz2C9VEtCtmErNuxLlGwYCJqD+FCKR9MhN+F9MIZG+H5O2hPlcvfx42thGszhCZG
m94r2PPSgIWIhJA0NguvZ57KOMpfPvWzncxitheevhuL6mGRATCCvZCwStgrChYoXTXFb8t1tDid
w5nIt29iDdqoBzCxqdKJqk3aCiWrNAVkfsNtWJ0WmUylXbW2ucLH5LsxkuIGeySJ1CdzfLMcFL97
OEohCWp5oZxCraLqjoYD8CRvpxW9xoSR5y5CYd2YlGaaRw0/fgO9/0MaaW8UfITYIwXApr5DuLWZ
p1MnHcT+GIM98xxP/qyjwLWW/PLX0I5RGTqqHjLKEQ3yCyUhd7+ZonlFk1qsY024McRySWvbLpN8
pBdT3MJ1q45ESrslv/WI4fWsLTLzx3jMVdrO050juzmsEQy7IQcbI9/xFPAowG3iymP3lK5BpuEv
BGC/+eLLJbyHIWzyeb0lvjLpiQk6w6P/GFPWyr4SmBJC77cE8SDUD8klc/ui2Ejimgy1eydAKf3a
qvUsmFgbNPoz62KnnftS7atvtLFoAe3/B50NLXfVvjLL2ni7/8huRvPO17lE8mS2Nxmln3R+zpmv
EKtx2c40Vo0jD0KhMB5GebSiCSGN0i2oS6JXpLfs4fveWfwcu/11tvKIDIwHnPuSuXeXUeNjbsBr
bnW3bAIwSvgzV0Y9L5o2iq+CKyBXUGWNUUulUDy8qP9BzaN2J4bdBP1iv7zLBLGLcmbrvzgWUkk0
eUJilTWOZo3dEvfwxxCg0vVnPo23GVsJbEU9D5El+hEs19debdRaqxexpZhYosCMr0DDYyUPeMUX
sVQT9wUppnUPMbuKYRcEihUOKZupwBj41zhlGrLr8MWcvOzfWTRRMcmBKwCZtfMU2eUn4rcV8xxe
BPliMjyP1g7aFI+eLy2FRACn7mH5aXBLW4TLkLnAW4IbnwQ335r/Wew+pUhFnqAl5GAa57F4VpwK
dw3DDcmwOawMMZ8TVaJk74+R/PWz5LruFE642XTn3wg9hBmMZL+wqIzyTrIfk3E8cVxkhh9E8AtP
SuVPEcgItsuKD5GXf2CmV90pN80jDCppZeQbSj9Q+wLaAOIugU0t6jYl01BTfmRF7NJgZQw9k14q
4JTllZnSe12Moo6t24hsIBNAWio+Pu244j4RlI0ID73fJZFH8+Fy9OWOhqyGcLaBJA1Ej64hoMKX
TekiudadCRfzkAXFn+CPBdwSz6b9bSx/udFoTBcyQ8a4KOQoWVJnMLUMCVvwSJkwH0QEjTW1N/s9
pS2zPv/x6ll3n/A2KaBvxnmL3GoymqvgCzNmSJj35Pw2VXj8JqdCZ1VKB+IrZWZcHBJXJ1sn5F2K
hMWifjxpYlgV7e97WOezYpP793jeCuaf5oF14HD4oykQtoXtGuh40mDhWbfnb25AuPX7plVWwHp2
5jdVmWVnhFJNLS2AXA9RJpzrkwBSS1nzUGJkCf4bobnQSI385kzow6lRerrrOj1eo6nOBTCmwI6i
RLgdGvps6F4tklmxVTgRtWWuLmOHi8If6F1TPnq1BOr+RFLPVzANGjdrPlu7E1GrAT0jus++jWVF
vssfOGcyVkOgwzq6+zy05vIcnkX9NeJi/DE4DDL5WqR1lIVxDv3wDTCnRSn6lAGziDJEBIbf0o3Y
TGjdlbUq8K2Xe7dOrKZow4JL2Car61JQsIDseAcNShKMSREufaiTgVMGlSQC1fhbhtvWAFtvcAAE
IUHnRW80aCvwXbJb3V54udsE0rJ4suNHmb2FYm7yek+oBlKJuXHyuXwUW0CmSaVRO5r9VfvScisY
c/fn+W1MMgkF37Cxt1RqHupK/Zm+wRM67YLddrcJ2bWGCicytRlnrf8de6tKu7mKrhLSSOTXD+fe
bjdrLT6SlsKMHSvmDl9VdeyH7kn5a6RAATCVNOStf9XUs4cGmMd2qan43F1iPBRL4mYN141wpjVJ
501vyG4dhI5+U/TymOy4K+ySx2+5ga0hzgMqiQUnZzgMxHBOVS3gd2sZjq6qNl3lzBkPQeHib9Hn
cdY8o7U9XyH4dpR34/GvOVTjC3st2b0zA30g9STz6HdZbOqvUMHqmwuw/yLi0mLMxKLh3iB+YNmm
iccV60F+gdYeXb1G1x7w+v+c6zTBwpnN1ExKg8q/q/+1GbBjhXEh6fEWRjDbpEvYPUqruyrzdcOW
C0NL97ftKBj8/mOlJyktLW588HD0bGxuB6pHbtJUXHUqfY9BlWlTYkeYQzahoOn4IjpXJB0Etf3L
h11O7D9wR4/+jR5T3b11nOpN5A7r14yZiqukHcP0BOz/b8nI9moPEF5TITym/gjLwcSOLBUfyVXq
u2jyxBf1Al5OJ+K76SPeduIInqSoFSxKtYiUG6Nwd32wp9+IWtzDNpxHwELrDpkm+twaGQOg8ndd
wHSYI+acVeEYU0+J9JnIWReYi9rC3qCsYmK7KzinKQnbgVhF2mjGjVPnPtnbzfXFgsdjyndmgLrR
kt7OM6pnum0Xfdd4EYDZnMd9ZgKQfEACSJDIpu1Dc0BSdOo3Z1dZO9Pd+aaAOFX+EjHtHVZCNFah
EeAVJWHudHnumYoJEtlw9szk9L2fFMr/gzpQGL/ShBAzQ8+dFdLO24BBZMwA2nQWm9DbLKUoR6Mo
xRqdQY8yUDpFeXdAaLeFW2gHMbSku45lzKxNQ/CxN7P1gJy3sKqoq3lT483RIyzSednBO8Z789GM
b3Y+i9Vrpu9DYQpVeHepfBWnFP5uTwMnkerJyYhquCzP9SRwuOWBzXNuJO2R0otMZwdvG87jHC/f
iR1hloFThCChnLCjFr8PuYE4zgE2ESjw116597ev3QVtKkSj1/Iz8vUSAOAutu2P9Y3npw/9gpU9
yanu2H8rRskTotfu7Lk+4tV+zOyUapKsnnkQl8dAFEMqsAfa/q8c3Ogg9hhJ88MhWqSVhCIoltPx
yelu+mRVuptemxMzTrbs3Cky+4jCfS9Fa/Dmf7BnM5jA87NdRlw1EapxGioUnt4971HyDz+jkzwO
/mDg78joszWiw/WpWxT0OgkYqEF22X4P436jFGc4KJff5kzXc1WRKGMd7vwRJiB2mSMc6fdR0Sop
yrsHPGEs3b3mPgL218AGVco0OCWAUnzIzdgkh/km5CwkTDB8INuZYnAP2pRI72qSL9ActJbHaK/H
a+FQS8OAzjkNNwtvb+qCuZSgseLrMzdyE4FosiUSLVD1ltaFAEB6RHgoo3j8xqTKonZl6nRYTM3q
IAzFSKwsT0DiNxAHr2r/S9Iyti7tGQIF5ADAcAOy6gieunLvTdmn+qMHto3DaX60gU1Lw93KOvG0
v9jUUmPs6sCYr809SyFC+Wn2v2FuCZghfcrYzhmD7aRB+4KOPRX/wW4gx2KP7uyiooo6GBb6VTUX
BHwEJCVUsE+7LBvmQ18Hjz/Lb7qzX//cEspMgiKwGlYs98UDtzaG7GQXI+CupOPJxs63yywrM6I/
Sv608U2tflrWf7rb7Wz5yMT69x5ZVIWynhe4SzI3Kke9DqqhFun6u2H6jzEz9N7ZfagojqomBmyu
afUYfP+7j41IOTTBTRC8AQbRB426T3IF8JHj0y8SChx9RatFa6e+s6geKeod0gUcX9J0L7NJMriY
OjeJ0PZ0d61orNU0ueMVdfSuk0JJiXidQfoQI735JKQS7/t+OHpVIIjUuVCrdiw4XO9iPUdKM21K
76vY00hc1gHm/rkowXU7RwhMY/SpmVBHHnATPhOoK1MkuwStuhohp2VYwtuH2x+zxeQKJUCqHuH1
IsYOkx8TsKvqyvtVjp8BlORpFnoYfsheNWCe6ac+EpDoltKIObh0z7P1fEf9b8iS4xQo3DQ47deR
k7uSQ7EqYH0oCjVqrNmf9Dm8Cvr8nwca/+IrgvcGFH/SGHOFzCZpUX5vh4SNxYaobOCXuPyGliyj
bA7pA96oPHVHILqDi1/ltoLxI7SurU4xizGhx0UFI3h0XtCNdIbEfIn7n0fTIAWC5h2y2GscJ4/r
FwJ6V6nHQdHXDyVrSL07TwESTN3by9JBTOlyF1RDa5HzTPiB0BVQqxGEUrFCimCZ2kbu6o5IMgBb
yr8qPcFv2rT94fGzecpYjjdwOoRY/Z6mAG3omPmDaOdPKgrV2uKbM7DPqdk/TwECo/Wd94qSt759
irZX2ApcTN2vQ/ITo7cwvdQORida15jsahWspqwuHwuH3kzW7jjLcHxa+6/8nQ3kNDn+IDXNbTeR
qj5Gdsqh6il5HsuNs82ME3eCS1NJZWpiyD92jeQAOiIXmhrqHQK9+3+DJAo5Kq2fR8tnutlHULHD
h5p0xCdTN2Y/ryMawKeEtpcK9fpENYh9aAkxvvzmCLyW9P6kvRK3aWjLSGFvprQDYmmwOEi7fvBZ
T+L7v3v4IMmmA+9He/08rwGMDKEjYlynyRN8kQ/1dSvrx7vZ5YN6oekVFfUziv6zAMYUaKovN5aj
WHfSi3kujNynK3WF0YGK3tm4/R7JzWo5Mz6NzEh2E/jGgU8yRYNXVrYaQSJsn6Cij5Cd6tfHbT0R
0VAjZ4w7xYiTZDSo4esuUojK3Qx5E6VzIbTVUW57IxnXoiCAABVTKXcvzY0RuiE9BJDAFn7o3uhH
msAkdjLYqI3naNz1ugPz7qQHLBs6Edl5aXw1I+ExE4TxHZirL84Gj5VOg8HIqYWbgIbDVLJmegjQ
PgxGRstKnksbju0rfqaYKqacFuGfD2wAh6isWbQuWPOc8mB44tucbHBfzpqL6QfTZt1z6ndgv4y5
px0dmy8ZPSX+6yLbBNZw9/cCsG4F1U5h7FYSpODjwikwUkUi0WazF8iy0LQBQzGV2pPARzwXfD5J
LfQu9DxSIe6EujJZD2mXGdNzmou03M9ZysUlXYaT5n+8oqQP6Vg1GJnX545id4S1tQo0Tq+njuIb
QJGACgm4BJ5Y+9jW7WHgboj6UrT3LTaeUfuLqSf7Nzw5AFQFNq0A/DXS/Zd9P7yx2vly2vopXUdd
YvmxCu1PrkeIa5gHQlO7wA39DesjRbTX5zEGLQgn9GSVlvAHEsEoHZGuiXEnk/bLTDOhnsfMgLG3
II0X9TQEhUDWEkVJai+h/DGpWurOoNQsK24pMoXCI8YmhYmSLkEnjdSqZX4NoypPDO53mfV12Hiq
aStrqjbq5KHGeUbeD31VW042jWZkkp9KgtHhinyjIwxZksAqCg+Ov1jjMJsKOlIIoZebEVM4nC2J
y8SQ7MbtMB4h3y+srJHrL5JrAVtbhuZPGtiim2t5vBfy+7xnJACrRsIgmN8T7sBSrZJPAd8vFERb
CDcQRWOwVRJS2rkg4vebW6khfzdKurC8hTLIfdXndWyWQqHQAPX/pa7Y8w9gTMUdclNm0I2eSsRz
u8k7DlOHWNsQ/qLuL/Cyxwr/SjyRnFAm3dX7X44LvALvzhYRxAe2tgJc97259eYctEJdlfBqtv7g
BGKKytcAT8vo9agwnPYool/tRTd8vTycvL5nJj5j4MmnTQb/r+q41/6rdAawxt7HkSdqh/WDmyx1
GClsQ6rq04o3l/IdgiNRTID+s0KEFQb5/n0qdL1VgKfrNv1SZgXVIynRuiTuhH6GaBpXWHq3xOGt
MIlJtLrWp28nsanWfBqPMl2In28zsxukHyCSYTVmcpU4zJmChJkxMFxu76y8mV8glBGwpP47LVh1
GV9QAjOjjS/lWRJDQn+pZRDFdoxGq8+NwXhfNhkAYrUGP/2JYb5PZOILSBzY5MrzFv3hlx1dk4Pw
i4SXr5BtevQRhjkbwfFp5qfa8QCzSIGK2IXkyvMuXXx7kDrQE/Fn8+iEF/zKJ2+KXO1HLqCDnqq6
yTynCmYlS/TTDe92hLcTuiFKjBN2Mt2O+9KyQIuipSqTIZco9z2UTYvKwXbhlsLvhTgJZPOkc/f4
QVRNteKhXZrfY/JG4LVmrCTv0Vt/ogEZvJQ+nx2pjkPkEkv7vBIAXEvQG/QX/Sp+BuQPqcGj1R4Z
DX5tFgDOY9UqIuhZ1WU9tud1uEnr0Y/wZIn7HC0ySsgbu/YmVbLtLI7tx2Y2WDWMht+dhxkehUjn
d5kRSMywdDsM1EB5oig3FGAp9Kv/sgHJndlVFP+Dslq+Q5kEL1PcuK66bSrdxRtd2B5ko9mngIyO
Yx/F+WYcYjFAzo1uUfLH+XsbgZHBogNNNcBLNQneLUJ++H0k/ByHb2VRHE8xJhRX0OWD7YA8aHD7
MTArvcJpHSHDExzd86xiYicl0oRQMAy3Om9RD+jAUYQ5fEU0rnYFqsqXkBS+9in7FooY3BFD3VLO
O5mzYWD6wZFpJRVDwq8hgiM0j1EgxOcBqqsXxjeM/GPe9ou2tnp+DEGgTVWJuc1vKbTQ6Mb0BHIs
2Yyz18+BbgpspxohozoR6Qeq0mJt6cGE3REiKCwUCtmE57817x87rFv4Cj7e7eZh1Gkxs0v7hrf+
xJLc0MxamjXXgxwexoOJHlBXjPy82cS3aZc/p0ZfnuO4BaDEZOVtbNBFy6cZHFHqKWXGMj2j84Ja
0sv0/CTP0k69N1iatOyG/LFYSUCYFGXvpmKX0ywyjGvyfVrQSFF4maPZWYcHnxX+OYMunhV4FHLT
2pjqrDq1Bo5jOurdfl6hyHgsiLvNp81nM4YHUfaoI9L346zyvZcbHx9heORhnmGyUd7mj0PDs/Ct
i24+x8Zo0MoPI5mLCWW8H88v6BWyZc12X/neCz7C7PQ2oL/JgeeD/c46YJmsrHTGfirTbHPFLf5S
GknLHSVniVJGZW+n1BIN7d1dozMlz/qj9Iz0xkTh9gsGHx5KKKQcsutG7A2ih+fi/c+BGqJaycRc
x599V/0bokKDdfoAHFM3THO53eXYJ3dLqF3GvX/Aa2fQP5FLd6ih3EIq+uIhDudaAHRR2E0KSFBt
jx3R9QXqcDcy0j8iF+Q7VWo9wANCNHz9KT6nTGSOs+nMpmBWdjczWqO1PYSu04inaA62Th5E4b9i
v4u9zP0E4T56w0Emsu4frksOomsQrdZGPYdvQPkPLwiRJaMI2gKCxokKkqsye0CiiEaqCwfh7KAN
lcMpCg6msqYt55hi/pmKrzRt+nFVE6sCxE2xb5O0Zw8N6yJqCXU7Koo4k+Z84NyFUcrnGUCSmGMz
IlPF4kvYP7jd6eHrTbWP3QVFzIOJMD1AP7z1ymrGtrwhPvEdOyNuWKkEmOM5JpWHKzbkhOKp6Y82
vHDTaPg5JssZwHyHoNV0ubqyow8OYJDJowfwodrPpAhslbM0XBuY8a8l80Ha+TKxPmBVK0UtkS1k
rRkwy7b4W3r1asafauoEs0VQKQ9f5jt3bMAaCuAuKmNtrx7prgX4DUWHEDGbmSLBDBe+Q/WDyqI+
/sqm9Q2nIax0SP+QVfn3EX7fjPx2e64pHUV4wSdUeyeX4pSaKevgQEmHnJy7PK0Sgu0JrVZnwfmk
X7ipV2D2wzNIW95NIDZ2tVYdK0xwu9pqeqSyhPOEPSo8ukJ3/cgVSnGtsduXi9vXvop3gXXEVw9G
CWgF2nQH4OTVbxZpOl8o8ROnrs8zWKygSTIeeruy5JFM/Pc1hQe+eGmzVA0Rji02jlHcTU7B12bz
yzvC3Fjbb1Stjr5PdZwBtBzpVgyjn/yep+rh9wHviJcVoJ/GdwyWnkHwQBa6IgMvSEB0mt9XgvP+
PLrIbb/XSuHOU6leJ8ooHOGZcVnq4zbvneg0IvU2T/DkYpy+6rCRe0CNFUZgyMyoJGTwK9VPPoSi
Os/G91q/i7cdBzMh0gzEi/yjHlk7aHHue28s5D+Ut/jx1Y6QBIX3GPN36di/hhBVZvanfKWGdsNa
N4tOmY5AQSt6qXDtAdEbgChy1nQxrEIgG7s8WC0ywNgi0VhJi1eClJj2RXoFLca2e8OO7Sz+/1+O
yVl+heasyynlQEIYA2haVWU+a9LKQJadxs4nBaMaxImaBEDcM/FsGg8HcLZJ1VCV8sBC/MXlVp/h
W9ugrE2lvv5T4pC/A+LI3fSQOUepCXtJQWBI7k9Ua/REmfL8B8FOuMFEXXDJ1aaI908e9tLQauYY
YRrGPkmI3kutongUR+mVy/EPj7EHj3Zg0dSfbsWssb2JYt8jhjqa/+Yjo91+wic56DNspJdAxitj
oWOD1BZVO2Ucqa4a+zU6grjHwOVPpWJT69ASHeIFoMHlsVv8UubaZ87SwjNLoRJA8/X5JP+xeAGo
tpY/ELV/RnxET5Z9pg3Nr6eK171AorCBAg+bc85cMnyRvGlBbXYhHfduuDGDVyRvBhqi3eWYQGuz
0m+lS3pOfAOvq2msjl8NjZ1UyVS5lYZ4Hl631pFBYJeK0hvun0Lp2Dc5bZXk/ghzfejS6PA2v8lG
t78Xqc7gJgDSJWpYRhpKcwA2gtCEJeE1/dVe1yxNeM949v2fIQusHXp44pPHOzFCJXyuWy1LSM1V
ps3p/sawycSeMsXTQxH23lq9tgzp93WLHT2ILAw8MpWTxRgXFyvJF1pYKbHt77183fEdHpCk+uvA
kIueBIyavqk50YCcntIFXfILoJ3XKixUcYd1FhQnZWFiv38YUigLxspgZgGkw/XsomqsD4L6QWYw
PE/P9Y0TA+qQS4I/fZJzDrQ7PDWd3dPlxeZehj/YsAvrNV7ytuDDS0II2mOBu/PNO1DXhspxllZn
6c5Q9X2UGYYxgv6rQDpNTT6sWg0ZZRbdCM96CGgv66CPxrOm924PKjPezYd+dhp0luYDL/XKxJHu
j1EyR7JbWstzLpQLpWcc8rH6hyShuLbq4rMqPd63adlzA1/baqQAmoTPT+DlMJzDTrB61cTF2OSS
CySPbpdqs186boiiEKfg0YZhgBjMsE6FEoeNzUbI5C3+zuwis1z+fI6LIV+IU2ulh7Bawziig5gy
Swne2GZ8wfet+4mctwMw1Vf18wUd75z6NPABcPp4j6yl7JypcF32OkKd+FUP3MFRGuggQ8MoGjIB
pAc5LuuPS5bGebo8PHHy/UJJcPFtKXOqLFwbero3nGWMrV9dx4VAd9q0wU6LMkVdmOujTM/pPVT7
81JiK+99Ckx+w/SDHCme0UP9QFewAoDUcwQI6mvcoA8ouIa6P2BzixHgFRXJAAW30xKbCgTrAD7L
elOAIj8Wpg3Gv9Ah8bCYmZ/ZB2x5pLxRFlFvOWuSTGfGvtlVcJsGTSQ1Gv9StyqnPOi/NibX3/Av
pw9OW9jEK8adwywAhcCq91Yaf01D4JUtzFtV2nFCf64xuB6oazfVzoyoCPzmFnEQb4YZCNxiJMNj
USwW/JHwyYA4leuxIlmhkIWgjl2OBLyTKlL2jbc8ORLX6FTCPewVTrwXnU0GTpduGZKZvM+T567p
4hk1cwf+NS1QgIe6C28rP1uMy9x2uGamh76eGsRxO14ZOataHQKO/V2rdMWx3aMms8BZy21gLdBr
hb2qR4ugAgd+QLTQUw0JXhp7giJ+ayoJgtpL77CIxJh9ZCwBExf7JJE9WZKHv8+geuIwZTxIYwPO
7bsuYDrSAkwRCmqX6tLInla7QxIvkhwKQWgMv21HJQBNop1Tn31y0sy9Ty2v7+oVF8P/6HZeUkGf
92at9gt/ftXkEg6H2aZkpv17bAH2PCYEbzXUAWUJoCP7N+KMEr//q/Z+AFSe9iFWOOSJc1GIGCPL
jWePlnHPN7u/X3sLaZJcxKKk3wpYAeCjXnmcuK+CmnBXV/w+DYdQpTIyZSPjJLhOq4WSttXclUc0
uvsah4eVgX1ZuozZJrln4WCuZRlgjbcMIFR27mIfGpQtbVX0RYIOA/7kedcQXlyX8rGj0y3c8A/6
AwElTFlOt4lUgV8bKb429qcgWkx5pys3euJZtOWDTdZe0vDOGnfEl0dwMfLbEnE2PoTT3bKoHDbg
ulS+yoduwPwbvdmoCDVuRnNQbPODd+tQsY4YsuXZvB8jYF+Z+8wileZz8GJJPXNhvYp82KfNOuBq
39BXUnd4inV0/w5C9SOrlhTMRB0dQAY5Xlx8q/pNx6gfErSl11WPSFj/glw5SalhJ8xcHWkK5bc+
YHPOsCgXTS0ekQlw2jzLe9Pa+zfw6z8KImkClEUzJQlk/jTEC7s4P1oSLhVex5vR4QIgCMXfODOM
V5px5IqOzPJSDKPZ+e23J4x3mXva0EPQ3prdXuO1O+IgW9OsXwyuz30427aVOpcOa+OMN8DPvtst
6WnthOht6COh6vBDJOxVlhv1PrABcJGBzEFr/mtybveg72WUil6lQkBEFBbWze2rV+sGB86bXjz2
CYxYBgSaqysUSONuVMx12KDDsX2AJ6qfkqYo1FY5kq5hZtDQdtj9lw7GlZm/fl8A4JhOyjHNvk2o
zfTDA8LaWuf706kVhmmrtKEWvw0eKXsOUB0gORp3L/eMLZmVwiLvttQUktbdehlnsxFM7M+jKnRJ
j3lUD0wMWezXTLcJPyb+rvgnJ4n0f+sayyWikkBSjUups266RxUUcfP/iU51E9CGqVQ1xXmfIp//
lytHVzZa5EXGpeq36aiA9h205Vy4yUaydH5Ik5w1R8dWjt9uvD4yy/e86G8a3RZi1JKdgfmXw+9W
WTV4+YJV//zKXr6asTpSvVPLG+loe2rBPdj7E7XTlVC1oT/0tzNMyR0r8Z/wVcOry0nsHzO1lDTn
lqLkEPoRlKsKVgypovtkDTpULQ5CRwiUucc0DwD0ozq11Y2SZsbFnA/5y2tNrPzrR6lHF+1J9GSA
2jBhcCiSRXKxxNnAsAS12JBVmOXQCh1P/WffJHvFV0w7nx2i1OozxN1qfQANfVUPD8bbcQ+/w4YF
2bJjQDYTtHyijmoSFi0fgUrQGefuhcFNztjEdNTeV60O7ejoqhmIX5vnIZfOgnNk8JfuhvF7lKbP
yoCwO/wjYOKQo66G6udU3BnFcP+ZqNvhQPySCgvknlyquNAjoECu4QrRn/7VqdH10B5WB7pw4B7t
X5nA8KiBC8SNO5IHo1lu6p9zHwtAOO1fIC76aPVzabrEiZy3FSk9QHVIpVZ0IZviW0vlkMha5Q25
m9KA8sfwe1rABQKzV/naH5tS9GxEucDpZe9UkSRTOSL9JqaOMfJLx07j/Z7ejScDRk5gcpWl+1P8
iP1eym5bplOVXCCN18frcybeK/8g9sxh4eacpJarSqnyUyoA+kzIjwCJRi82r9GpHv7AV+SM2dhk
yozvkacQGBXkgvlJp7ZtHaqznH/j9qpV1JhZ6l4hGTqgOpIRzjsFWcuKTcVS+v6raVYdpB7G/s4p
l+m3DvmRABZOs356+fz1YxNgL/kvAMt5ahfj7PD5sgHTs9Y7P6UN2NOGZZA/+KX8B64/49Aw3Bzg
2D/hiYIgovozNwcO104hZfbEcd4e+0G0t7xDOq3ySvRCx3XSNk2fF3zEpWDTp/2RDATHaTP2bdjX
JotfE9+7IkXGQjmu/CyzEloCbtnlONv8zjR+8wsCP1dEngXYy4DKPd9JkHNgrY+8spVnBjqYAvHn
vciUS19BkEIUHtq+l3bC9Mpg+xWVbKpa/Hxlx4xFoCBrK5B6W+eGjrXOY3yLGycEZethGMPiTgyT
Es/UlQVry+OTr7P3oEmkVcaXuM556XJx3zr+AwEnVLEPROZNb60tpKV913UeYWExyaYYWTLDZsUP
+C578d1ZMUpHksQYnwVk575iaiobPRlk1JcUjtFGZ0O1iXWOwDGxC8Ob5Ti6DggCIKdIhUI9kmxe
Cdh48QPp/PnyrKnZXNiSo+ncYzzHg7b0MBIS2/mpjm44PG7dMb5ABvlZovlka5YyXpZd0S52BrCI
HrihQFO+SCnLPmq0fQTKgC7KsY3X7zdH1nCN3F5AaVrZVhxgdPwDogIR9ERW76vcnRuaIg4pfye0
OVWLpLJ7fItYhcjCzdBHl0jENlGh0XhivEam+J+HIfqa2kz+sUnM7Ca9I+PIplZsL6FlNyg154B3
0/2G6iAbo167+489GiaPt+9t/V2A6VcAt4MUNWbWG64JB4LdN1XGSKRwGWk4LHx3EHB65N85S2MN
7BbQPQVcXFMOOfpGxY4cPuZqdGWjxfd4Bm3T6YfLL8OJEHkg5lfsBJKzpehpxkqZTUo5CQXk6Eji
39m5+d1DaEcjNpZ6kA8rrE36xeWzpAuedf0VKpzBGg19FNHDX7AYWzgXe5AlROVQOCepZKT9BBlo
ewb02jAKX1xPK4tXyNuYA0bmp5P+gaooEcIWpZGd0oBY4eBP6C4s10Uo9bhIjdx46+Ib1bx97Sph
vl7UCDcfyyMA3YW5n5i751IZThidE9kn6VrSRQl1e/eHMnMcS/acgLiS1YBjRxStS0CLBysxSLZL
OdDuCZZUEbgInc6GluyVrwe9sj/ybotUIttZH3jL21VkxItQ/rjaDJYKgbrVs3uIbOoIv+NlojM+
I/VHAObnvFCymhbytBcqFPMKW4zdIPCz+1Scalws0z+wu5ghBFeay5ymiIdjao7tWixCmVWVVB0q
DbONY5lkXwNNPTT8HTEUc6thyN7q53U27RRJFexnueAmqAqk9j2mkdXyhC7s64TUBDKQWohYZgr0
BjcE7+Y2GnLeE6aM1Ven/hv+oWpyQsaxyD9wnsmhNwXGKfmZTEhJRjLOiKa3VqKLN/bhs6EBDWSl
2XnQj6V84tZHQSOPMmmkV1io3xx6jZbgABEpeMfoIJkcfcpZsz0cNdU42z5W8/MojkfKZ6IVBCdh
YYWBmN+Ba0b3fHyb+GQ9o0IyLPLYWYFzChh+0k1xmIGy4LqJg59iF8CkBTcgIQvE4zS/tE8+GAf1
qPo8gPbQd/d+hz5ABA5uSdECvCwNfLID+rHDuzeF6GoQwlkxSGbYxwfKRDlWrmInQmRvohrpt6gS
wUhUPAaReJ1YFm2UqGsmku/8max241KBi8wz8CgVWklljiL77j/YZvDGh44pqAb2+ci6rKobfaxm
2Qm+gB4ASkgXzMHFa57qCnPt+NQPYzYGtvKnIGOiyuLVDosV1gN+jtwEYO6O/D5XKdK3SlkIIR5/
OzOfwrKfNoSkawsZaJPxSce2jE1HZcbp+KLSwin0+yGjc//rTFhJdAcQ7l/hn4fjotzxwrslEP2a
MZ8gczxSJZqfHQGinTPM+oLFr62E/AnE/k0d7dzQGsO1myaZ+HXPYrHKhpkL/VF/k550oufb9BS7
jjsWAFcLfVEo9iwsX9tCi6EFdII2JPYmI9bQlWLs4J8fTeBzYXmQOb05FIPyeK80AaqRgyNPXmVb
+wLgVR5phAX7/nMR1OaINFsrDPzJyCeLm8lEBwpgqFY1jiSvuGoH6YwciYR1jmUXzQiOEArdOXos
SoafEtfHZAPGMXAmabAPitVUHwEjS70aAhGx+yZeU1Qw6sOhv/TA1wH/9Ub/Nj4JM0N8qzOQEXws
Unc8a+QsNzIIrE343SYjlcZ9MoQMDXRDbq0Sr1EqspkQNd357VFvh6amYAlCqvWAc0aYVxRJAyET
VnHXmoFY80hYE1NTljoW5YT8AfOTtph9j+MQiTdouhyidU2zCUeek38MPMvBfwLK5XAkacipDIdH
AGNaqrJOi+cUd7qeLIUTsQQiD4QPKgwLEgWEFPNV4CVXLaNr9NnbrzYKeqI1B6KMzyTxpWauL/8Q
mExihSfUVkmhqA6lOsRXbPYGys5+AGEFHyctzEAD4hCSrbdD5aS85DmRugzr6kEO66JoEL1OXreJ
rttLN3/8yUWSVi4ANXxuQdTmyiXsDP6TElo9M3TEf12iwvnrkCN6XwamT63CD9GgHkobIezVG3An
3+s5ckq0oZpCJBdFnPZ1ZocWcGetx4ARmtc7qa3/O4WiPvbQPcJSN7S7TJxnFen7AMyRD58ha94K
0UJzV5WbKvJvRpBJaP6GXa/auRdFPWPmtN1XiRxMUvztWfHkE8kz4zHGfGWN1AzxfXqur0+UcYXz
qvdZk3VQoeuotsRgH4irUBPUEki0LTFjwdlnFOq02LQFJaDD/vIIvgq1vQ3IV+a88X0KXNpOi+kA
dP9iQS2JHNqiRoRCHrGGx0eCCFYXtjlJozQgUWt3g7K3d+R5WDrxcK1rLADcKtwGIMCD5e4wdrjd
5yhY7QR2pK7YrPXuFqr7yCYyapa4Q6X1Vayx6eh3QJJFTXaphaftWSYJgvqZLi35pstHG93Uqmax
5ecJBrJliRkt8Ce9Yt6dZEvmb5v7Qtv3IU9ZL/Jm8SbWRS49XJnGMef/xgTbpSwEU1ge0R/Bf2MX
3BR1/DT7ERemcmHmZibNKn1M0UTmzj/dnOksG1tQ7Ey3Wr93KQpqcGpaiMjWQJqsKb4O4lYtnGJT
lwHa/OSX7CqtgcIfgyV8q3kQE60GK3mQ/2aF5TtNSotjc5TyqBePisX/0pJLmOn95pAHr//9qnXb
/qSvbXlCAEa+kPFCIpRycAQFoDydjzD9F/kWtL9k9e6N3G1i6cAmDOfV5oXtRJ0YCEUaVj3ZdgTa
LRK1+HxyGduwcsx/LnC5Ue9z/DwP3YNU6klfYC99PmEsseN6Xwxv+9kMZcZmNq0aPwBSUxfMRwba
v428OQta9fabPvjPTk1E7zze+YkPyzxQNEQi6XuMP2UFRSJN/TjkxApNL3xhDJ9kGH/A3G/WFQlL
/47xw7H87O5/PN2dZoowjFZbDghvgC+DamTdKx/gt5QDId7NkUWmu1Egb5AMURpxAyfQ031dBaop
kS0TqcAQwuoxIYdz32Fhqv0FZrN/vSk0AMA4gOzoNG+GorZQ8+/4nNmhwkTzuPE8D2EZ7CLk+XiB
piSMM+I1N1PuOAxmayF/2vby/zB54Yu5HG52BurcbZRvaLMQYBdSfd4NesVoeImpBoMDRlRp0+Wr
KSScsM1N237GQ/9pyuvBUyf+RW4MOph4Y3FWb2Rqcs0m6EWEnArgLXv1ZmbI5oTdTbkOWQfRey4y
HL6raj6pcfQStuy85th9Vm+5EaAvkL/qSWV7dh2LQqZ/ieEMixSyVn0JbvwXEyGU5cDGg0mDxxYC
ANhNQaTXmE3aCYWAXIyXJenILZXpAnPE3o9z28PvqKPfhnCz46uU4/OwACyXGbLD7guxIg2LCfd7
t6XGgAmfX4uQGuRwo8YE8IzWVW83xoJTxS7SFa1ttLt2JCS5Oas/S4RdfAaKqHwqe07n5Cf5LMiq
ggV712AhJ1awWaPfZHBDjEZaDo+5tmZPsJWB9FNqZH21rQA27cs/Ttc6UIqLtVTQkVbPhpGtPKEf
YVHGlsxB0K68VL9WsMCQaqm9XwM4zQkz0VRL1wnhG/qTZYVqukFVbjmvqC8zOj9+sH/l/Xyk54bz
Hd//22wBIV+lrqdybsrM5AVag9B5Sr71pSGAjwGYghLf3b2rM/6WSWnDOZ8jLtxxmB76PM1Fj5kQ
bcCbrP8N7iryPihaPItgkBwybe3lf2TLZtdB12M0I2z5G4xbC6JMTqDtMD9KcZx0SfSP7YalpVrd
iswstqFEckb4XbtgWDxy7yJqLB8U3VjUDkYQ5WDaY30FOg4SjQOJeoeeGumjEtwo00zIee4hmECF
AzdpVuSEcw4ktNbQs0wUuoZrBeX6Hk1kck4ArjiH3NyDLFnlkgJI+prnfdd51uddHVqM06Ek5/y4
xSYuumVd6GHhT3Sg9p9OTaMZLp4ID3doEiX+zg7I6O9k1W3FLRWIZ4hwTvUfu819RE34TPX2Yuyl
SeVDQtAYSjztjR+59qOkcvdOo+u0j9hhriMfLfPpm4Ry4S1Oss8ZiLFstM8u4/F5YQeW9khptaIz
/U1SnH4052w0FlaokPXx0nq/sQMiZc+ZRSIcgoI7eWVAMS/O84TfHVB5d/moXM92T8iaSCRwTO2s
sDHfdW7M49xkQgWACo3efJlVibq5uTrkf4LUBrf0R7X3bVvo595ykre+M7FbQkYrhTniWQPZoGkw
BGM4VYG/rN4Qb9aLGCheDnZLjkYXr2D3is7TMmPMbaYk/pqiXRdxLuSJC4rOYD8SMculB+Y8K585
p21flsfDbYX/6kxu36vSNXesS/a3nFCR88VhXIN2VC6e6xbMYBjUP2xQDOzgQmGx4HIR4rBy05Jq
vGCWmYKjbGjAxnLQWtzEGCRMcF+EwxGOOjooWIrdj6DZMbfETB78Mz8K8meWamvqZXnkMeUXHDst
P1RJgQy/w6Prw1tmOtIRD/pEUs7irQQi8iDfEvDonEMGeZ+uR9j/NfsuAY7dlMUBpnQLJjBuHenN
Mv8JVg0J6qLCaS+wKgSksFe5XqN/NgTW3/psyOzCgIR9jtMaoadrHgC92hS7BDKR13t8q8G/Pnb/
JgGhtoIJmKQd07ju7UL0UB3oRcm7c+U959eWG7C5JcYyWdrwfmL4bcI5rvJqvl0yMryiHGJTCJ8T
lrOUqXQQtZL5ouW1VToFr4lx/ywUgXUd+sTmNPOspItTWg/e59r8hePNGjBaGHZvmMwzCYQIXzW+
87bDnJKSj7/ozqq+SkNj8Qwm78vsC95dqEWW1MVB4pkUGcKL051fizMwtBxNnCEMrTbZdAX78S0N
y+ofw6+hIIy6oXbxbWeEggOLImMzpVuS8FSJxZyUxjQLHktIvzmS+5RjDdgCtMYNxRSHkb/4Pqk7
UQXkn19tF/+TisgAFJvadI6kf4I2bJTvikvv21RqRK4LHVeh8flzZHnbO4qzSIjCcdRvVC+ALxyN
f1HOTIFSuB9kHkhMMKtBvvAeYDEOoSHnhXOKUz8dpgIHyI2o3jH0ILVk03zxkCINiOAZ+UYLOUTm
PTMgbonRYi6NqGRnh3hHyl5z+iAYzAifN0mpZWuw1OLShvWmtiIBAvegfjYoYqu5E7Jmb0ShgOiE
WF0Bcw/bmLG8dKBDfeOwjNDi1NIrPdGvMlqZyUVYbrVJoO6s6Ve5Qo7g5V61SX5BapC+Z+f3Rnn4
rlQHI+nG3lTdosm6N5IZqFTT1yxEeODe27E9TqmlXjCn7VfwpqDQodI77KoHoL0UpaiO+H5jp+SY
ipLkGZvRfIxJqCoXXKyx7/usX75BsODkSIxh8aTv7wT+cCRHlq9Ju/aqQp+FZO9uBcO7EBVpyJxc
Y2bmf7N8rLNrUXYCVUxlZhgV9Hm4euLeCL77+LMW9+6s0inhXfHfRBr+qjc0b418WakeJ7vDEa69
0faV35LWKyvSug2YiB3fglv/mY36bhyNa5rHOmZAJQendoxOljcWDs63/Xvo6FIwP7WcquyJP2DR
WNoZUTglQPuwnLMgGjJTAPe0AMI06DNRXKam18b34LOajBgsul4/aIEVkM7ZJ9bUuNx4LC5SHpAT
5Bn9IQELlx1h1y/vvgd0NQLIQX29rSj4iHwp4rNVOqwtjfDBoPCJt8fvqoenL5GUIA9dQ+tpg3JY
4topvQDH3IQACqhybruRyS/YYW7+PpW8gLoTeML5asjZtP5CctVroyvEEeqbZoFF0mf3mfCmig6o
N0Dr19R3oBIya4bxllqKHs18F0wKe6YyOFfr0MOFKMKQGRF42UDqOWRvTeDnL2LVXbMVZ+VKHrBI
6KvFhq6rEDbYePYSM6FV5/WeSqboM1RGtYOB8oxPwbFQlf1K7RUMoTLlZ2so6yf9IQ2cBMGy+oQH
D/4H4q/+fSQKbzcAaDXGdjmbmZRJwRnxJ05d6Y5VeSdAqa520wncieLGSkt5TdFVDJMIe6hvftS5
c/e8b8Ac/vqv+GnlR498xbvT4gDGd6fkWn+Y0OzOxnIrkleWSOCvLdRQ3dMtfF9dxii/XbND/bV9
BAAPVlm1Kx86OSoactV5ahrUwAqGXPassV652DmD+fYNZAI0TQAQdfox7EQmPs9r7hI2rHZsqgsO
R8vQJBo8SeUmXEa2n5BJSSy68rn+xggRqIWJlXiuABvESsZOci+pWslxIa68gJo5kDCaWkl98R1f
z303utNX883UziZ/wqf9eZolZHFiGqVtTpfT6sOgQEcxAW7RND7QfwrIkHpIj1UgRzKps+a6K4Ls
kgy42768hmwVNxxKapudFqAI7Vko6Blshp/qB1sFItyS+02kbC5Iry+cRdqLfcKTYFLpFsWACpnl
5p9z/DMTAovHbUfUoDYzmRcEPsMFwE6BtfiMFUDZcFVfDGG0q2f1lUGtQLmP082OT4d1pUXp8/t+
5JK+73cZ27WTaVAaiIMvJL4pgHDT2Uvq7AMfgXVCYJ9StdylYTXS72gfH5Ogu8s7CHciPqydVsWc
S8LT607L53YZHM20OHMAf01359MvvaCpBsXYEoXcTEq/C4ujfuObwMHOAvhSk/LCEofqC3RtBmYx
giQyGaLNLDBEDfFpty4UYPDliPZiF3sEydWBHr6aT1q5eD6W+/ZOCDTULg05qJPPjx0KD2+DfVVM
Eyk9O4EDIvoDa2yx1AjHu43mGVa34gwYL4XyGsNtVXrHxVB9Gv24xEurr8p1fnjoU317AK5K3FuQ
EQFMzQ29rX3t5VYFwtSP8T/CFVRQmysmBIpIIyxsTTuGt5XxtHwQCPnkh1M78rxA3D+EL1LUBvO7
dCTdzudYMa9X1AhZtMsJ33FBLdV4j3Qmdb9UlXgZJJBz8OzIog7QoWf3F+/RwkLpzXKbvYKCvTiq
lk2NlABELYB9/8UVSTaEuYV4r9atDUOrcxyQsNUhGWmrk0Tq7tZu0RPqWMMNufSyEiJ4eVA5S3HI
2c28pRN4Q+ubky+wNk/zvli3Qc3+XJFoLB44t4YpR/9Q2BJgGyOHsqNQsLgk5LeIogqA/WeUmf5o
xPGD+KD8HDvLYw0fWx7yXah3nSL4rocVdLQXf6a6e4KJ0lWzOo/Sy3I+ZGb15DoG1FEk8KwSFYk4
yVVJefDiQCKTmjJwPlKBt+lPfXKj9L+mpnCCq+Yx0uUqfbsjV31lnA87k2HZlF0II/4+HCMol4mm
owootXZRPmU9grTzH9ME/xTNL4NdjbdyUSY7jg7IMRy1OmjU/8Z2FmgQ22vBCKkPTVRbufwKwihL
X5U0C2O3io8JYPsjqCsTH2SRk9BoL9e2C4dBrJKmfcu92lh4hWKYPpKWIVsuN4BQlY+Q3wnZmCeQ
EIKib9b91da0524IsLLfOkQ3oWY22jR8if6S/V+PAkWby9+EpYRHz/bAgLfSNzXnfU2JrAeVfKY6
a+kD91SoIzEtaTKoTKbrq+61AHriIF7Mk5ZUD0Inxsj0X9VbmKshld5cUX6GPVSXcDBUkBEX5q4b
s+ExAG+qhn1Jjtsc0dlJVNHsrAmaYPSUyz3sdvKIACd0pUstB7d+L3LHTsvPLJ0VpSpQwTBriD8r
Cs4KzbechETHv422OZSN70FFzMi+MBOIfYKXppdPJA+dTFWsq9AdDpr9MOv87GuiXOWi/ez4N8DI
9OIKueSZaVxBhSynmJ+REn2dI/0B+NftqYDCVhc18SMgAVQWtob9LBMMg6VTsVNuuGZSLoZ5xmxR
O84BZhnFbv4qdN2g8s4pZFZIvCtz6Sj4xXKrXkNcLs37Ww+KRnEyGn1Djbi4vNM44P4I90xuCYce
m8Lo4fYPcIi1bAG3bcO7dZJrYSYmsmLjw5m1xSlkztazx8f3AQVb6KLnK/mVX/OBM2IEHiDnDkLZ
UuJuThd3PkHYe8E/n7rlw9ZZwHoYMMunfWTUJLGC5Uo9M9+rJVUAr+Rf5QSYwVpeM9qFOx0AUrn7
v1YgTbVda0dB/+coWeonpRTifKxzi0Bq0yIJDw1zyHu5gEYW9eu9Un0ztIiKkQ+wh/llMJTdJ/ub
tuF8xYGvkQSzh9LiwQCUZd+3tm25TDNTwGSMgOWwkEcuA6HPgT0ammc5H5vYj/JAAqJ5jMYpxHg5
bjU+2ENykH51C2p1qXcfLVJiYStgDbNzfRuBmqtoFFSmYYzOj2/MLTzon0JJ7ucU2eAaHPkuMi29
CWBbRRrw9G331/7+Rw9ftzYcgIMNjQQ3CPHolIOKCBiNHRnyG9Jgo6QSmexmZqfqu6ceZt97APOY
8SSu3NtOonaWyK+ZSXxfgXPJqRfJyaTPHfDDic+9uMTIAjNshNVB4yg/0rqlVwkZuU08SqeKqgMh
oXzfhrevmCSjoCZyFlGv8eMRo2xUXK2Yh4cvVoIIbYi1O0BO2zojhznqf0/pys/7mPCBM6kVQqJ5
4MH05fRSBjPq4C3HV1UvRkmvU7yxcFEAxLRviP1J5HoEtg+f+lDzt5QSahTancIWOUDKDTUj41OI
7vAmrH4kcV4uS9iovhNBRoEZHfI5tYXV/EV2uJKNyI9G9u1l0McgYiEpP5jKt6gv/gQQ8UAjLlL1
UXEuAc9CM59MVzOk3JIHxo57MzP9aMn+KpP/7PeMjKAdLAY6aMvdOm6hT6OgEwm/vYJ8ip4WhKvt
wAH0RsZkS/LFYigohZ8rogjugJcbxbcp/KI6A8zyZQp2RH/hHMvhS4UGuIGkT271HlDhn2q9FpIp
CXBp3+e0HFTpLA5WJD1SuWmF+W7Uc587MAjnndOXmBUIIKknDARrzPaK92GDCT3+NF+Y/+uYFpE8
Dz6U95ipjhkTG2xrE+0IMm9vOusHir6CQjUVPyZXG/ldF3Zse8SzFSRojmDn326xo4UXd5iIlKt2
YSOuaUGvkbUZYqm3ujuGBlnvWFrb2l2nngvSHZ4y8oaJmztwArz597vxppjrGvnituAIl/SAsS2G
isV+LV6dOGOroUI4z7oyKr/Afyj9y+Xs5p2vIVN74GC+PwzrkkxDWd3wf3TMzJrOvSV0qrH+aznW
eK/RepNgDm16ja9tzlOLrU7Krt69TrqUbGDHb6c/7wTVfwE2PRS1xWXnvbaOuto8mr1GY2KogC3b
hMm8hhOykmC4fkub2xJ4enu0IHzTfY1Gat2uWFVOLIL6av8TFgLumjP/lGgadubsanLDXlHF3JKs
vl1bNCtMFN8CYthjZiJ8hf74+jaenm9Nee2wqJNMb/zi4pU0GFlt7UKloiVcm6XdP8piBcVw4Fkd
YqBR9RycJczhPhAXmr+Qgb2Pac3UnInRHQiyOmpD4Rl4bHSpQYAjfS/gSX0oVRGxk2Mqt/zVERPi
ebStmowhYoLfNsgsyb/yyPh1IXaZnGBtaROrBKCdORXTFKNwOPXWYnjt2JTk1TMBLC1adQZTGiJe
LHuVfVhKmWIskaeRs00XzCBEAqM3tgKEfspVIqnasbjtTYGiHL7C+G5MdfjKD/FfOYlzz3LvegG3
o7v2dn0a7Nz2VFwiJNChganl+liM3EE6cpVoVJAGqqvGewP0yTj7eR+m8xdwvxXb85NB6Nr7Zirh
LIznqLFFkM5qEsT219xSweuJVeaez61qQ4FNodhtgFHYGxLMLD6kwe+OZh7I7H09+tctQXkoKsJE
ntRc49q5mbhgS+SndsAQk+/yNZj01rNe0TutF714y/aQ/zQygZ16wIYPl5GLy7GX2da3oOohfunA
IvkwTi7mEhp+yBHTjJ1fli/QNptXuUGyXPTN84FQ0lZh1pzaJQPgKJHUo3bVPaksQpIfu2KvieV+
TlWF46JEGnVndKE+z9AB8ND8cBKiocDAThxsUckyjIfu2RizUAlVnBMGk+1kV43xYevGHZY7hbjS
eTxHxJsmOR/l0V2J6rZWlTJW3TEeEINUgc70W8M5zKAshd1SPzJY+ZG9dMem4ZgR2xtp8LpR15Li
G4DZ8se3huKAMKqx0pLkUo78rZTg49R0XRrKPePme+bdHI0Ibc3n08XRS7qYz5n1/VCTmWiWz9De
zE10qoncT+E9S/PI+QB+X0rCbfEe8i06FZGLAEm1CDXHKJEOH9Ar+aS/oVtaPdIRaBnKNR776XMX
/dOSzg/Vg71Y0iEGmIv9VTYpVnD2Vui8XpnEHnM/vnC4kgS5yttrX8VXuzqctDGAiQh+cL6pTuvq
4efNhuKdS8hbMuyweQDsrkiiVN21AAVTlnck2OPGb5yjMli0H/Kk0MtLTJwqMnLQZhKvJXGn/nWm
u5F3oty7LmnaCqzFKc78cBQZlDNWIzflCNaLnpIrBLFRlr+IaiOEZagddOjsG58cl9k3I155jCDu
m/SecXh43ob8IuO9YiAR3V/yfSQaKTM/9i9QAtsUpQ0I9tXi6zl/aEReOJKQZTbUMpHQgWIp3wYu
vHPSivmQBKiFwv7OyfNNmcPiL/ndZts6revliZEt8LUGc8q93i3qzDUtE5B6KgoezSwxkqOEU8UN
KIEOMhRNi36kiEAdWFf84JG+2bqUQqSWTV1/UzZUKjiwxLyq1KAIpHqrAzsr71QqkCUKyXcjvBEu
H5mb4TuWgIE+4HXN8hBapW/HGcwPWYcCRDlSSm1AEBNxfktI3hK1LaDko8r6w0nWkNoVab01U+UV
RkeowePnmGPKle85ddiJY12WcVMgapNwv3IUs6YGaqtvPPbijBPjqgECIxXQUhh7k0uyNsP6EoPH
Vsj1yXRdjX+4Cr2OfRQ9hCZnGZg8seECC3PiHzDoYFWHrT+sI0IYEkNVIDy0RF4FMKxze7+a5FCa
po6DWYGiqZ865KfBNwEHBi34RownxOIBLKbTwGU6L17l2NuM0gEeoXQj9bQOLvYAvUhEfy6OeZak
BHER34N0z7ZnLxoJk6rE/o/ijzPxRFG1Hf+LOhKGJ7BBiZ6NcMpl7g9tUlsctSzBgGTrTJ6NRdWv
fs2I991Mc7T1M8XSyPPV4w9sNQCj2CoNEzR441J0T1XVfvaWUh0NyEJcvByZkDk6P3cr7pZ3zhQk
BPUhffluElK5OI7ztYcZ4P3aZ7WZ+foSlvhqI8GwWWfJIr0tYp+2X+ELIf4UtS5Ml4anpkAuBdNg
QOnjxXjLpb9gVNQ1j9MdbIIDOalUnaPrtxF+60tew/qGI7x2ymE3Q1LLwMYUx8c6LganWWEyNtRD
ISsD6eeSgMbpYB7omN8VdbDNPdjwy52XlSZMk2JgU/6IhY3Vrky85eMb4oKNbrBglf9wPlvKYld6
EyRjRebG5BqAjV8r05P/py4JZ00ecb/Fn9JnxlRig0TTUzCA7hdT6kqiqPLjf+k1OZ5ceybBaHVE
s7OLtOQCScmPZhqOffHtk/xoJvKWV9NvGcmOX0qF66gyUVuNXef7ImgjeiFeBbEchGN0m1aNFKlk
T6WC1z/H+dNvnOJLSnt+svg/PTSo6e3X8+0Ea2IDVdIT/PYZcm+KUGUFicyMIFdigWxp7V9MqrYB
oXKkF8/3SPY6AMX2HVE37y0OaMxtIq7j3mM5Rkfx4vYjT5EbUapbIhPPfw0iRWEIZ927EqDhNY5m
KA/vtFIw58FRUfhWVtT3FonnPeKijVpNo7DsBw17LMsCiAIVNmAJeDou/xoVsV5AFa0TtJTC/Pzq
VwwN9VHil980iUgLT8RK7nEG7V6lSG4Azibsr3rEqHAaOr+qapdv3k+a3N35R18DNpf/WijvqzDG
nRvC4IgtzGkN1Zjmk2uEaaaXhxXa0sbT+/W+dr+09KQSP+2IvGRnRpDZo2yCJHxBwsNdjzY0Kwni
WTrGuVmFE3gAcSytSTGCmQWbHbRrPZYrJiZe/Kz/QOeOd+hP+OZ9EgPj9exUDYYjph5inf8iQgfB
14M95z3LMmNr8XZaDWwhKRUg5fPBQLw1WiHflB8y9pcTXjTaMWNVs5rJLekOmp+Dp/zBjQDvV6Kn
i2yC4dKAnobhq6WLtnthn/czzm2pa8gKUZghBhn4xdSJvw/2V0UfZCK5dWDH3kOp56nh7+kg3EQ0
EmvkYwyg2QS1zmRDkRuujxfPIIlRNeZBoWvZYaCIoOQxaqRJMQpLidmKpNQVnoZ4sX9gTDSgc5aN
nHhx2vkLQWpzjSbxmMe6q/wLTCss95wr6CASVMs4uZrHt6RI3N8+I5YT4tr+CnSJOicBdUIVvkFr
iOFZ3grQZDrvJhPBBYPILwCmvSNQUuyU79gKPJ4iDGsXM07p1dXVfPEsqM7IhxW9VknSFS1KEl3n
9bVsrGtflDxSAyBnFDAl6vEc7wcD9E2UCvRKZyzFKEXTwuV0MMEEuWOeP/8pQFkDWAc8epieXMQW
B/uoAVCZonzR3PPvQcKCWJJP2U+FkFozeQ2NfITLcNLikRUJtvVs2wcoeG4Mo0JL71gDxeRUwI4E
0mXbRqfGkpGydn8OPj+b/KHaA7JgWPi/67qfeP6P+sPi+OGkrYzT0YdygKQo+aJjjNzmIIPtSmv7
p8cNwD3+m4OqeXckEHQvWryVYHZTF+StuIPWBpsIdI0ft7ZSaexa6m3goKb6KlUrQi0uN1ZHgIU2
qFAxGkUH2s+gJPRMGJy9FLX0F14t8KM7k5lN91hukv4Yy956Q6jHdwJrPt3lJ2HPbxFJXVsmTZO3
VhOiphdWNQFomRihjb8JsB0JdQod3cJvjhzgVJmSS13dZbMrxDhIZ9TRabMMSyOFOZsaTcLwB2GY
o7lPfBBg7NlE2bI4Q0pQEv/wUz7VKCMlU6NHvf56+oRE7me85MAPGRnwqtF1wGXYpb7YcUbDxrPG
ESXlNW89Rw2wyP9orlkI9uHDlSCZdzV6QNk+DTqYt+ZSB623TOgvXXIP0UGzl0ApTuXA1EpElqMR
je3VWHBAuAJ4f0zGD2Q6i2CE3br8smunqELsiBVtSstd0Z7sDxmtr8pkanGUsMTe1LZ45Autk6cw
SxjV6b/Q5bEr5+tmVNaU742BdgPc4HUwCB0L87cHhz07kwqQTQkXPLN3rscz8Nf442q0nYGVNOwg
CGDZ07l3rP7q6hZaho433qcnutQXajMsZrGUZ44nqIWvXt0f6uGmmxD4+HML6qzQ86L3YQZiXxZt
WnJ8MuKpSnL3ZQjPbO15QOr2shz6+DT/8by21rFAfXb/Zungo2NNtYwhfDKVOwNYu0gcZEOtDz+3
I1fzKip1ySXyY7eD07Iow4oraUYPCwdq0yP2j8ySfs77uJlaBx24uVOA1ZenYAmRqj1S37eG+GwQ
OwvILNpt211NrA/cIgEtSk2RR6d8aqIO1yr4JAikUWIzZtfv8Wpb50iONOIHif6b49iB7Arc2RdU
Xd03KXYlVuFDw3B0U+F3B3J2rNHsBcCUUp5cm4nxeIRZv047dv1CBcrnypcccNKWja6zaYABR7bJ
ItOHxRr+HPTizsirUrjNitadqnWvfaHmgfBIquW76J6OpIzYCDrW1izEymR5mUQ22rUCLNw/HK79
w9sFoL971X/tl2Mp1UXAVajmMatwTwOBnRXXxNphvTYsMO0HoOBtxncNWpRXwCj4xnoN0CAVpPoD
5XDYarwStDnpN7IfuLgNFo4N4STSrcy9fuepbQbY/PY4fPueNMetRqm9Z5qRI2TAHoV+hTkiXer9
T2bJDsJIh8OvYKRhEcg4NNiG1jGmplC2Xk3z5umIPDAqQ+UkwcXRdW7QhbvZdofqS575cF+dCYCl
o4BevmSg9Dy/41AOILHf6DoM/hcrdD8dB0objGZIRS3GjPEe1BPzWHK0ThRhPxFNtysxXCBwGxfW
4Vh0MiMAiiekO0kZ4gLGtiOEQimE/b3dv0nQOlNrJKjNB1ko+UoXCZasDosvEt4q0R/1vtksWvNg
Ffj+w4mQdwAbwDTR/q86HX3OP0YPAFSmctImXbBu2ygA4CFW/ogWZ5Z1O9b/aUcFStOavC07QxVM
Ty5EbHj09ByrnHHTcej04FaGmtCr5iMmsX3QBbfGTYEXM7g5DnZYNRQJHsYCHrwjPaAJIWa5Lu/G
AYW7ghVTqoMqFvnMo1H3VKxiYYFIVhZCk5j1PuWhMddIXa/GEWzUf0V9pJmL08/IMtj4rDjtwoG5
PV/810ctJodSVVsK9vsJQLEbRAFiUbIxas68MWidzQ5ZbQnL8SVhCr/a/W1tKehs3PPwkIxAk8Yi
I8x9DoDnSnW5WR89rxNdyqMqLFqRK/cX4z1MAm7qKqmOrKgmxFFb2vvkKF7+56u5QBJ/GaDyFSd1
NrKZvS9wcDVGLAAyTGGyY02fh5yGxoLB+ryjBW8djiTXu2WRLWHqLqPigr0z/lFLYQ71pG/SOYm9
Ljrn+JVkC+BwFVpo+qHLmamzKObUKg1rfPDrDJk2mzP2hABFqpDwQxY8vmeSL2IoTz6NA1Eg86iJ
JbTW1PQ2MX6L1C3oXt0FmsBFIFz+inH/ggsv5PWSCbqAqG+WHnPu1BR+WEBfqx8Rptc2NIs08xjd
nXMRjH99OI3Q0T8Q+gEQNX3eZdgcEJhHZxOiJxd1B2WMTDr1iZjTGyeFgOfHBupTojf3QhoWDePl
SUmynmj67gk3z7Ork5o1i453ZRVb2LXgzv7aDH+9PJvLH+/9kom/eVvLMkJfbtWxj5aPFQtlP7tz
s0Oh0pvOVQxX10l15HlyZkJKlL6VBPmZz8hONQp6c/Cgkr4hQp5Zg/QDDdIGy2n6skaPn31S/auf
3Yj9l9h2K3XyUJDskZGDHcj6WHY74c4ffMNJJzenDP129rsZ+Cy4KuN00b9LE8MyCoemMVOtsNK1
8+EpwMFD/hdZsfpjgozIkaVAeyv22mhcRpw0jie7FyyknD4du5Y4zwyVFu/66gch1droKMPY4Qw+
YCEmW/LmkagqImnsHbwqnnvSorh47wXf51r+WKGib/OYJrBRQG3syv8RZoMDMiuo1ZwwkMzeP7++
d8wnLEdVWbcqDa69n2hkyU0m9rbWfMeYvIwvNkkDDh7Gha/ft884pxp30LVrik2xNHbL6Er2OBVA
c/i+ETTulDmpRPHXxJyt12qc3lP8fDGh6sYnbVVRC0DfopzRyaeQbxECIWzAyQUsnMM81VMV0oLT
nKEVc/0RaaAsa+bNqah7wKgZevI+0moxmrFwTaVg+oeytvqBUJcwyAKZGfVFiBG9y1V2SfzIGFtE
xFypWdIiAZzY5acCXJCfsfWKeINIeGCL/WdCSHQcMSajiO/rZKbkgrw7HyUxhz48Q9qHB1ClFjSR
ZfBf3dfY1ewumiYVFmRWIbx8izdjZRGrXt6Utviv2VQqgh2Iz/fTFB+TGZ3nmX6686we/xk7PHXB
Tp+zn7lj3L13Xkyq7jCefnSHYk4cL665sFDlC9mS4Cc9CmH+8/NYaW9E1gUKi/0iRN3m2onAVSf4
JXdls+NmV3KBT+WVsF0E/oTxk1Rpre041OCWWjkCXr6zWNssItOgzOciqmFWhue4V9jUKXTXWELF
cDtnVe2JiqwAmse+annJ+UB4XJk1rGTnagPAlHBRh3HEK9ze8g+w5txRpAczNsZzrW/nCAwKV3u/
dsfOmwXoErIMGmvdeQLP/O6pcjOhq68KS78X3ySBrnzEEea9i8kjRoq51jLDT9XrPDlQrzU1/z00
STKp4K3ZerhjBomShEVV49onmmabpfAP/cwGeInx5Z160N38V1MmYWPHzkHBdWEAMSJMsce5u5h9
k8uuVm6fWiyU0PvKgptGI1ixJhRtD1atOXWd6YHnJmC+lYSypDvWGV9dAoBkNq3LrlqQuMNP6mO0
DuBhtKwBycr4jzdh3LIZA+dMMY1TNEAJTQyRmC9MCY8P6YuNPr3K30K85Qi9jQ2OpUlZk4KbAwp9
QQnOZa1iXP57SyfqsKO0DP9fA0LtlGcNna4SkeKS8tmTmmmN47NJAjChZNHiyH51NT/tug+4tZQq
MhrS/78N+q7ktuwyfex3zpMpnN+h3VvWUM2i5Y9+ihbOLDVQDcDgWAPNf9fGKXo2GcsJgwvk0D+U
hi7mZvF+A9iWRS2tTc51PDFoRmPKCiRGnUFo+3f8ku9AN6Txs+BuIHsWrCyh8ABGFmQj86yVO+Uh
InBfqjBvf5k4OiZRqydMY3JsxnkibKSEY9Wo4PiP9xd2Dl+RPOc8djIQ7Pto97QWze1S4woqqgyn
4p4ZC9l5ibX2VqQqE5UFIFBLrS6lv3aLKQ9cyISXyOUu2wptw3xlmWlI3dOooO2PpPow3DygXRYV
48+NrppK9G9RAm+zPqgX/gtNHeyjb1CSL2H3+CnbU6kBfF2U/3Ph97y8GbkjpszEe0wFuKA0Q42f
PIOAIsTGPYO+N6OW2GjjAh+kAKzUO9sFDWUWLgnCzrkDYunZFjRbUHTe3vXW4EHDb7VD+B54shDk
pbMuvF5/D42wGqzPyErpLSQ1TEkQ7Ib6rrW7PH3uzxeuGfkT9vBXNtqWg1CgIadK3KxuBZJp34Om
ZFRaDBQQ3RKNkZ+oE4bzWPlsYVJZOR/wjLxIt3Z9+OzgoiwmDZE7BNuCnfOBEItXLC8hb3tyr763
27QucQ0y5xJ+AV4nrAce/c4FROfcS30mdNFnMzi7DieRqI3Mwb59VvcRdQpmxCQ3C3TmpQfITg+/
JEWVhDtXLOHvz2ommb7pAMA4IRgK1hZ5I+K7zruBxNWf0TNJsP0npuIjwOpIKuLU/Efx73WzVR0j
gRAt+VjFaAdoqp2pOiMyra3xYFm05EPsEaQisyDr76EDpfQJoXOlGE9RrcFcSvBHaHnZeI3eqRW2
sVcTG0zrlBoDz3GK046pDKua+RTBt92cGEtyT6g9v+ZMGG0wlVV6rYdgFmraEPRnWcE+aHAYbVEM
4vJEbCL5RyxaFqlv/jSw3RXtgE0NztUdeoQweR59PKQsV4qC8B+0ZAELrW2jjeOrVYfyQ5N2q+sV
uXQSba0Pa04zKFf2ZNiFmBwYr4oSwKx9IHaKWLOvmKvRFs2ys5aNWEF4xUGvh91lng2MlLwbJXG1
oNOeYMgcd3y6X+evjJvh8LRKDR4FqHurRcHyeElRjYKE3ZLw7rUW2SDEixiY2bEJT2Ipcf+3QJBM
EhAV8PYe8tfeiHCKhDtJblT60CGt4RGNNymS4TC3gO8bei8IT6+tY5V/iEwgELxlivKtUq9TIfy8
m7S6uCsr1/kuGRxa5p8xEVr49rYSyGElRE+9/AdpH5SLu/EDU9qoHVYck/lb+S7SGDu0uEkdYN6w
Qgz2v0amiteI66iIe0qKrFLucEr3nHRJVLz17W34DzZlW944vnRPWVBR6tAq2MC3RHKSTvW9Wqed
ges/JeHenX+mJnuvcSi/386DfrpQWuRhnpnOl+CdEokpI6HkG1Ti0ji0D3GSEMQZvQoHxfb610ou
q1TC4OKrN8N/IXBFZpCIU57eDpjdhAkruhBI8qpk+lrD5hWIFJHsPDM5qlAP/0gjahHEn/s7L2sd
b4inCg/M73R1tf0IS+a2AawqIQvbtSsW3EaxIo4pQZIMMMqfC6TfF5WZbmD1W7Yb5X9uPyYT2CkN
bMKonGLmcasZ8o/cH1q8akhjSIHnuFS3TAI1/I+PaGBbWlINxOgvjiXLCNtMomH5AdOp/ICa3gvS
KYPjb8NGkpURPwrrPHDiNYmjThCdNWJiTibrMDVcXqxpZU9G+I801L+M1EIys+1quUZ6cVQMoDPf
dBCsE3/3zbm473UeL2AEGbCKLScS9ixVswxmPEwb7b5q4iaRSf7RE+JL1mWT0eZu4/vEseMHTsC9
+E6AvfpkPA6gFNAaCrPHQjxr2XdsGfL8RCPon4tYOKPJrVjHDjNZDLQM4WRoFxCDDHGroRoTylvW
cqrCwXX0/BjRZEPX2wub1QUC/hRy4xcFozXNLolPtHX8m1ORrzbHr/0dYtuFIC6sWK/I8yGSlrkt
uz1ET0wKElbLc+szXZNAhkVDXRldTqLSgHaX0Z9PtCHcd7CTR81TUwbI7owkfS9siUYbcpwh8xIj
ezfKDcVNO2/i/abABFkQ2TDr4xAw5Ycov/yDjH5dFoHvyEQxBxqBMcEhuzMZEkbSSH/eKvL+GLRs
reU34tUINGbsRPlc2I1ae9y/NTKSB9U5zuQrZgL4B10V+33UNn28Xopat3R8B6fCbcaUn73K14Zl
6UI3Ix1CyNU6HmczCAXfOqVMD4c3wx/Tg7xB7rJ3ILhLcbasBpICeVfxvQjDf3bsaClVJOJN6HLq
IMJppNXMvPir9/OGa76OrxCs1B6qqh1Fm/f3ZQiLD+9kFIfGhi4/lLyYJ//yCaFkdoJUjqb3gy0a
mbm0DeGWXPGLQc/1Bgw3SSOw11dOIyzV03euyIbUsZvpuvX/EAg0EJ933qhHdSQL9Qg7oWDwXMf2
NImL6chMrroG0iETAq3IvvVk3zXy0lXia7kOKCviltqgBVaWKOA61N5MpWz0vbon3XAT8DAWMO+g
AX+a2/OEFemH6w8Hq+5zaGPIbMHWrPu/5NZvfmKA0O9k2O4ODn6R2EC9fmClMygrWMnUzMO5Xmgs
ZKaiecikAKpeQAJc/NMJmMlbKQCZY1s7+jbKSi3ckQPQFDE9toYekOfOmhJLwwIUlgmj3Komgedo
o5nCfEGS1JF68Trp5NlPH6yiwVJJ8JrfVJsXaPwDu/SF3R5Q/d48n5lkgakaX7GwF8vcNAj5u5WS
fKKaYG9PTL2S/2ZjPH+vAA/Nb9+gsrV7ghdHsDdJLTL+g0xvBkF8h5Gq03qJAMNxuNaCNTDcUrkR
QaA0WMoazIpnOnE06Q9QdTrFafXo6d/SXHIF7BCTMF3XIAudIEPLbEGcfsQC8YuZXYVSuZyoeYsM
1bsJqXBIglLWW1vtZ5JQshmD+UKqASYkXZWcIwpcks7jXIMZiDLHXntccG5fMMfGGG1FqqbYFiDf
pt46u8q9Amr81qYAvyG75O3nNth2fuJLnpaLym7BYMoVceU6DDRXiCmH03OZ8oAXAyg2NTl7mFPB
GcAiKqMZdrtXWGT+E5KnUCb+4T8oDIeEFPAgde4gVHjdSjajFkCdvNv4v2nqnhTFemcLzNogYx7E
hkR/MzcLkXzveLiOUvDkvH1rSh8vV9ZJLN1KnLPLy4GPKbK52ZzafeecBu0ZauRldSXL9s+ukRXo
RCNMvvJM4onCYe9XibiNxEZllJ+J0brX3yRfKZnV2fvTuO5smvDjVovuNDkot4bhqJ5IgTJbcXwx
xjQpjv1kFE3xIBsCXqL9EVNHYn3oUh06LcOMF9+odnwpoISjpwrhYRViTdaeZXgzoQtocCb3RXI+
IMlsaAjuH/Sqs9f5BPLquskX2dD7V6goeowWAANdQGnMkZmx8BQRjvy2lXgPAKd8yGQqvuZOLlfI
nO73QXHt9XVdJOtL7mWhKoUk8RxAkBWCTvYZCka4SUPlSecisq2yUsKZ908Sn7fIN48uniQeBpkC
BPbzNT98Oc5LUHcAcEbFNd67fE/mDa9KtMcuHKf5RSQOw4DZbhuu0n0TxyuymZORShMKjr1h3iLl
/84oU7AApUMwsbPLm60g0RKyTnlwAQnNhdZrwRiuGnHzIJCZKg1qXsu5JZGQlwbLx121632nxd/h
FtF+goY7T/AE3nhBFV+Puk4EOplOfrpYSA8mJV7Wv6RhQiEmVp/U+T1qLTzcHNIH95tDtlOMOn5I
6HUOc7MP0FTdxWlqf6KuxDqouoKrgHlKGypAW7IScyuRMBw/GvLApJP49IG7k19JUSAzsj51ioX6
7u6UPfEWAEVVdgtIx7jCj1Hr/MZ9Xu3AU2O6nqCiTNDcRzDRrixEShAWhtvL2at2Qj9/Mo6S1Ees
596DReTwCd/iLkwUiCsBVJxCejJXffjWHOhsFUVaqHcRmldGhP693BVfrtaiq1SW5M5F9PSL1i5l
tz6ORHiNFdizMzVzkWz8uNBBdTID0v15oBs0jvIR292kBpdgKGeQozykSueIKkX2hgfzN5jKO4gi
5lg46Vm2aQ7gXomJcdujJUrN4DeddAanS9RYpFWLMNHHvV8l0xf3tA4cUwumndHfM2OQr9agdtQW
hxAPJfJ5YWOwmhL1WJuT1nRwL8tWrdEPI7meYi0omo/JjImCQgiyn385I7j10G+6jROTb/+xBye7
QB+BxAlSqHopJlLiqUqw11TiGUFD3p1rp0x1SCGCvHhLyWWFE7I6X3rK+g3M5c3wjZ7gPLxWaEEH
H0D5lkmSP7uqsdiTwD5Q+d+qXEjmFf/2Ia5UQn24XUHEyBGrzrwZEg/5miBNKdnAtUAm7MAwR3LD
bwtt7Mxn+SUTdsqUa0KP9tBgnO0y3JaclbKWni/zECfhBgofQzT+28iPUe374FzLbzDsWLRYDos/
Pte5v1V+wxy7BNbSdMJpiSI22p/ldnkXGmNt6Koq2oDJ9hMTaL+xjujIhdKgG76Nrb6sEnoJmAMt
kdsH4++EbSI5nS4zpyyyh/cxACx5z1uioPaJvGsDQeYEOmy1ua7rMz4ZlEPC8ZGAcmXK8/OIE+Dw
4vJ4oXk1Eh0Omy86qnx5EJlt3kNdl2MInxJpmXHLwXuiNCax+5x177Yq7cjoU6W3keRQ829d9WGy
9i4JhktJcuaN0pAQ4uDnd/yfXkDHyV5xM8lmR/dGT9BilUYQmPG+leRTx+TMDiwQQZh5hOtc0Pmv
begvq/AO5MPA7krBNUH0Ov/GgQmi6+PqlHgx/bVqC9RECqlb2Qt3dZrnPvGeYiJTEkqujg/egeFO
CA+yij4vq8ovrwvwLSzfFCzTPCPPZuVfxmgAMSf1LyhCDqTLLo8XseKj4ZUdT+WhMXm1xSb6lOEu
UQrjfHU7sDtrGn+peGJdyVbPoV2uZI+uwuZzrINBHgFllzOpTG54/yNwuVkTejPZTCe/iRk0imoV
gcbYwFEACGfzL+CJi4516xCiMeoHL81+gfa79fi+/FPtxE6llZyKgPI6IUaUMEBIcnMtEwwl5fwX
lf45oYXJgrwnw0Xqhoy/myNl3NOWCa9nbmnFYGoGlsDvytgWoLUN001tcintu2lWbOxUsje2zPkc
dkfwQX0IRk0N9OV/SFVJOFyFHCLDxuo/iiRBZWCsWIuW6e06/pkkB00pYQJTsEth7K0zDmdu1UQS
lSabIBJ18SutPhoi2bPG1QSaIJyOO3w+qNS3obpfl6nrSgU060krZSGcyGtHkbhS11rfR9Fmle5s
25FMwOL1Kd2PZLUkPQBhnwZEXRj3a/dBHhitP4tEKyTLaLhxos+d42jQYdOjv0zItnhYxd/dWFuy
DtKgd9+VrDKkIgaEJ6O7gb9oPIkQd3N1FIUeHfg+kXe3t8GBCezLciMjC9HNugf2O22E6zOz2x2k
FNF+KvaHRxq+45gKDxjXMKQoDNTPzI3/LBCoVysFOYl51PUz2gSuf+0BsXVc3gIY0fDQz/VSW9/L
rIeEiN5wsyYhbDeAANVFFhJIGtCptxptcaquRXBhv46jqLjFX2M++QVNU+KCZ55bADdE4ctSvJsX
I5q3vIyki98/A2DBxH2GbBk1/mEe4j9nM6WnNTZHSCrjlZlqjtU5LOKnb7eG+DAuU812kkuqmma9
LJGv6wJwELnwTk4Nk7vgmMr+IpiqGHZPTDZ1jvooV6Pr4C2DxNehcn9fMJ8nZnJNElg0ZDZNTJTK
t/70IfecCbYTUkJf7yxHc4GGltHlSRnqEVOFhyi7OzPOdEXmzuY4+HyeKcVjM8i75gn+8Dh4yN0I
pnuW592+GqyUbnOSpvsVlPmeqnY/d+DMvDkBxqN+RhG6qVVwIKFmirFJSjVxnjTKTN1dUxNfSbb1
Nz03BCC2EfmoGfhOa1Sx66VXe4TOChLhWoiIuO7QDRuhvXV0QyJFDqT8ot3ORtphYxdM/mQstexM
HwkwJxc8EYDjkG4Zrwofd0f2FZDGcTHcTPUCg9Bg43jCGYubPIp/YC1KpbjyqX5yUWUEcdQfpHO5
UvF7PBGBl7o07dInWuSt43yyWQs/1MeNn/3BQIbKDgR1BI/fBb0ArbGzOSQ18MvjX9ZVxZ+GdTMc
daJq71X3WPZgCNgwVO+y8lOPTMSUA4MGePrBRJozF4/XwXTn/To7mP2tjbSKqGZvUTEjif6NoghO
xscTju/uAZC+A2r/ylwOWLIEhcadMfy0Lgqq3Dz2JDdaShFg9ZkqIH3wGaZDiq+rc5aspKkK5Xvf
23ktXr9+qrshvnDrDwulDDRdHDeYbyDLMmRIMMKpNVH1jFH/bPbkbfsXIRVivDx3+m8e7HySVBVk
EIKW5ykHEZgfhFZPijx1YLbeYscsq1ARwmkWqLcFajVDTHP7IBUjRHcMcvNbux+XfpVlyBmVuZUj
WvUbEWpazADANC33Md8DqOblUaufFoOSlfHdpYM3gcUJUeLYOIUinoC9HZRP2QL88Y9+lLEw4x8w
QOrOfm9t4jLLvqWtbq2NX4AvC2Bp6xiLezwj2LZ/VIIUbszdxoYEoTwq7vn3hNyWdARN2S1640MG
RhfAL+ZhtyidtNCiqHNkV46lOFUqr0qmZHGtJNZHElG1eVwGqzH79p2rpZeb8L0D5nInA3MnZZVE
wYyt1rw4EIeSY2tqFDQZpZ+BA44yWtsF01mdtc1VrbTOINBg3oSVmj6KCCddY4sy/kfMBxPojQd5
NibyHooNIrXSlQ1BhaTBIYwI5Ro3bYYRP7pvvKZxlfV5PEvyTs3lbnPYW0QyH/qUttyq1OrkcVhJ
g5FxDUPWeFzDWwmOwhwc/MkCHSFzT4gWwdUKt5vktWb9YD/rNYd7NRj4m+Z7Y0hl+WNwPfPLtLhb
dI4NxG/zaatT7osdnMcbn5dJPAfc9PiI15DZ//1WKEOWUdVL/IKf7tfTOpNl4mM+Toflo6dDvxfQ
3u5sIO/Rrd9iVPaeHUgcN0bjmrVBfF7+9NwfgGUuLtceJOldk+HjQ+stICc33WM0d/fDnEszz69u
CgL87agZkyQMzqIWZjuNkypLXf3pSqheSPmkquz39PHp+8tBb5EUeAlcmPrQRr48C3ogRnbYbEKS
XNHJxY89gVfulgxGwyqDdYxLLiMl1CrcrZh64wzZnROpw9LG6DtDKgv7NbPlq/dZbLk2I2uh23Zj
SzhE3IqE0U08vpvUoEdp4ww955CTee/E5E0wdmSxXx45fH+kweWO700FLFogx5NtV7sLCmXFO3r1
6lp6CGLNU6DqrKUGQQMfJVepbt9vN6LR0Y7Ly3n00agsApL1EC8StJWYk4PTywZs1FjJ/dxUPPo+
igNxvK5zVOvpskg7PRXXoBEIaC6sOif3BZE/nrUwU6Mqsn1q8ONo0vpTG9qAraEomuZuQvfngAOy
HjzvYaWdxvC1mfn3w0bSBIu4bEBC/A7U1jZsLr5YzPpzLdIadh2ba2PhNRDTtlobsXiVwrFoGv8j
o/YgrYcoaQ5lXw92P9/kMdWQJetlkc7V0Lrkywtl0V00BVZFHdJ8O2cqG56ziCrUOc4E51+a6Kui
rv3EX9WNdsuEXqCs5WVZi+L2dMlDRz7a7oTyVOn2J9kHfYn/AWGiGoueZvI5NnDrtoY5N3KJuuWw
zO59XTqiv98a6/n1Too/behuFgcLby+eVYNasa9Nqn2igX5+MEPQzsjg5Pkwr6/mT2NMTw43yM51
tdy5JOWgGNHvXAOAwF0QAad014o/GgaVZtvbsGM+QUPn01RkTKv0ZMgN+oCVeiP3a46xG3W6eC2E
ZRU525dWbCDNL9RH/yWKafSZIyl8PDc8oPB0TXwI+XLzuwUKDw/Oy7aX9lTk3Ba0FMB2e/QmqquF
mcl/fOwUroo91ogL5LrgwqiJ89OZ7p0r2M6dR3d3WKPrWRFQwoBD5HBGYCtNA9LIdTZ1ooVTIZAY
OTgBgW+Fycabr+OkiCGUHUuzcb3TOvoyi8A4NrBERLneeonRdbVa3sxrefjaGsdKR2lOlvcHEy03
FzURr2ynEy7NUmw/RizImevMBox7iyo/VoXSQoUAlF3THCvmnDAAxyIxewC0nNN7V5v0FR89LiNX
OUSIOztDXxzlQqpbgq9N0ddbCPYPUwtr717Y384IoJx4vCmv35F0RTaESas1CnN18W/5mIJG56vU
bfjoySyeCScA1Ws5kqGx5xl+iQDMJYioG5jVTLTtdBu/BAjBEqvCvvkjsKny0a/j12GOEe5Rp/ud
ja+wqA8WZH+ukJ2NDy+Tml2OVQqW2jqlllG78koU+UyzG9mNpb/H1hyk3eDFOLJRrabViUakqULT
CUQHkMhxm0SEkxulV5cwmC/zm7bxTxqY8rdMEbE8RaqCUdxkqXh0U8gUsqARFiqt3klxwasJ+p5i
gdVyPWABDuDQJVmxLIDzBYyiTurjY/aCJbaEjXQObmxlMKvxQ1b4pm5uuCmIyxlSat7of7CHPTTm
2kikLVO6g/CzwZHKpgCLBNF5TOaReNN5bQsGWCyN+PRDNB222cDSH79FxXfrwVFhBNQYb/9yKaIu
J2+oEEDOf9vK4gcGCuzLPKhz2YomkTBk8qIW5BYat7lsdLCY3XnJxLFF1pp90Prx7VXSMMX/xvMc
6FsEmM4uRJQWGhNLeDItrQyasZ7M+lsIiTodewzLa9BfRqufzLfmRYK+OpPI+ZyK87nUTTvgsHBp
ysggDQo94aCnfCkl+qzCe7W2uWdlxnlafxvcpgq9rutDjqvG0L3twKvTl6YPz0HiQKEJiQy+2JN5
8p8LkHIEjRvbpRS6i2pPfg1giDErz/EiCac6EbDYi+kM3EE9tkXAMAdixY6nlpGFV/DeRLk4eK/d
yAauWX71F3PPM0xsivtMmEkVHcih3hIad9VYbcWPdVdV2+kxeTFduObLjkblQPJsZHvQdd8ezsHs
VxAh31r3dAMs1Cud9IdVgv1FqgTwUTiAk6Hjo6IAzv9pGS9fPDqIBP92HmS1AB4/a0rhyb3NDNhO
PWFHsErY/9hRh64WBQuVWK89kGKYn9kMwMtAa5gRTItr7Yl72piD5+FGfvrrf1bkLFWcui3ML1XM
YfiWw1sG3Dui4ZAlsMgcnnp4wMoSAkH6Fsdq4a2+cHyonZ7OMXnZ2w3zFuL48cSFzmcknUoVk0Wz
y15wjTZu7qOpHjf8QwHBvhilkkw2yU1ZawNlCruXh9sXHvw5095eVbqWgMCCpPfq0Vbu4ujTzHg6
B5BFo8STn7BU1z2mdiSGrOMIFjdDuidHbluGs/zM67vqxRF1i7LW35dzIUubxdSBqkpG/9ojgAKX
mIF50M19AGR8JvY+Fu1e4Bm0Ed5ICx9WlUNliTvhifksMGPT/bUzBZRTWDgtp4VQpY7oItjWhJhz
arpYdJJUEuGcXlvF584I8ypW5ZhVuBAIozck8asy2EHTkT140n0Wx7jqPLgsj1a2LzPgBCbMXu/T
gA6d3juC9+keuwTh7ri9nmkTszUrdXlT6LyxfOl4k/0E8IkrNdif2JsWV4EdVIY2RaucYTfJYS45
ucnpYnA+zr2achAIvfhGGuFeaWGlll1HEgSGOtytnhJffHx3ME0o8x+G4M1If0mIBBEW4sxejctW
EmHC7vXBHUu6RVyyJc5OtPoQ8JVfW+8kWfkIEsFnKaMVPl/YOlbHr6dOIB+2OyjAY1YhZoG4hFEC
BTZPqCjmE9fN424CYMMxD7A/dr2xBGf0aYT4TV1Wnt+YpqdoavCHP6Op1WXNMCm+lIR2XE9PNkEY
4cl9Q7rYvTwpZA5jXmwNlwKhj+IlY2anfv/TNybq7sGSJe6ovOQRbQPgyFH9jhh0piawLwiR2T3Z
VBvU6q2lOMZpP+aDKeaQ+EUcBME8n7mk3DifZHbxgMH4XciY583k8I88cZMt8L+EWKueFzIZ1qQH
BLPoFWf81bB6Gt8E35m5Ofs8+AO3zb13ey2OWanw8XIL4xYP18LatI78X/il54fwTFNW5PU+lV64
buOBeOMMe2WBCM8Equ/7emTHeQNjpn1w6h2apkiQQB/j3p7Rm/pL8G342mb5O6KNvbf99JzLCZO+
hYGkENdHxuggnb3qS7ZjuuwJI7/O7kMBF2cF4HSz7LnNKvPfHcN+UBqqbGt6wPEw5AXQ7moTHG02
bnr4RP6YZZeVEhkV4MIii2dpRH8VNhB1orQmyL1YmqvGqEyahGnka6kFExuzaeBHO+OEBSYQCmYM
86iwJsnfN4kj55oCbpayyda/j47yxXJI3CwV1GN4OP8jXmoFsU3ZAgclh9aG5zmuO4akIoR1dK+N
H6M19JD9cmyaoxiy6+7lIs674BPzIz2MhzvTovM5Z3Eow4JrQGFVPBAxcCPnvmQ8XaDj2Yt4Fale
6sc4Yqy39Sa2549jw61xIgcLWu1tN3R9pyE8oaowqavMohUVgWdv5Xf+73r1EUmudqiOH8z7KRZy
3xxawPPKk0/uJzJIUUE4sLlQO6xVgkN42M7unL2g9moEuZAJsBLxa9XmGt57YSmsrhh8Gl1/4DIF
2Ke6vr86cr3b3ZTziLq7RfsunsACTYNSVet/+bUnrkT0JS6tbuZW9TJp1VniDr9vB9MH4U3j+ZOg
NgmWb4L3XIlCmBKlU2LWNPF3dbK+qQY9fEmtlYMlrvKr3iEgsI6m2X3D6mb3CYf+gAlpAWwPiZj5
oiYlgYTk+kdiR4NJSbH+deirqImtQsiE+mll5+4eT7ZcaCeYUu3c1qseH2mfc7ghVItW5CF5M1Dr
UKFj8Bm8gUFu7nZXYCqEOAIxUQBXPep2ZVNHZU4l9cMFzKqYQljFmCA3XNsbkLY6f0PS3/T2NM+V
dr4uc4BYjE9dEE702jENx1C3H2lFHrAz2XBGBwF2JRRLytCQDJ2LMkrZJcOyRaOVzZJlRhkLT7cu
P2MM0m3OXeBXW6oD6xT+vFuY7SxuRRRQYPry5G/fx8QcnIVjxEB1Juxw2HaByiyaLDpGjQoYq4NA
p9qW2WK660imwmlKE0LHEIpA+LrkmPdKg8RRLPXYRbHQ240fxaOLd+YJowfp/kG24YT8FY0FObM+
0iscS5kNvwkeGxrw/HotWucCZU9fG6VknMY0HsoTfvuCvgB0K7bt0eAy4oJh9R/Hjee+fIz24BCk
c4SGfeaxZKda51H8qkx7HOnupYljmW9tA0IZnD8BNlDSX6o+2uiCywF3rxvNtUPyWuTUNA1LBEnX
0CJDgkU+UK2pf0rP/azfRe4SYLPtAgIn2ClhDWxskijYhxay+Q0xpui4G2o5sbPCQv3PVWl7sMgK
7TOQcm8/dkEr0K1IntMI62nZ1KaQrTJIGtz0mkGAIcEIYV+AVcfMl/uUBUDUN8W9PrpfT6b7+6sd
+a2pucKZh7JJQMRhFG8f5rknHjVLmNQ+b6uyy/OuDtog3KM14SH19BXbp2uQWIGRbGKx7++dGRWW
c/ZyY0L1OyUrzqmfGB2qSv1Efmri/b6h++8B4MdkotphlEK9Ee+KJfhjd5tz4+tEkONuDSUWGOjU
sEN5MB3oYOgGfJWWf2vjTQmuYdedTQNjzkw+CokyUEsa08xxDhvvcp1hW307h3rkCjLbBTcf6MJb
g6QEtNr6V/uqymx68ecTu71HqAMxYlxCS/Ke+q26C0DxOerM6kP1K36Sf+5y+mOhgtKEdi90jPCK
p1+BUcoyxlRcAVqQ117cWxoPkwmzovI1X0jtvXn9MmCHJwhS2KD00d6WvRYMBOgX+4wri4YXHhj7
UYlpUu3KSc6gQnlXz4g77wL9vuVDbn88Y4VWBOZCjbceec0iutuWEBB7neLfTgOnCG/8NTIfsy3N
4F82kotgPSePJYGbkIfPvFlIyKeXP51nQLVB+FGFn9xyBMA8oXPFWpQkSAxIBhq2/BuZq/HRXnmT
DzE32GsNFYyBTNVLp74Ag6z7JN3PgNqAs9uqf92F9F4udBIxVeKbJnXTXBgX6b9K7DeKI3vng/hU
7KE7tvQeMzo6/2bgC1iKq2hOvYS92zgMe4KpVVhRtfnNolDgslyda6jzmvFBsj1iRnbwo5MQ5vqK
vkwL9lQ6d5JTyxfPVOp2lF0Q9cUgo2xoWIahedKY+4oBh5wHGkmGpygQAw9wUIrU8/EPU598aGlG
9pfKYQv6arCbi+z0fOoQDpvycW6X7p+vkqfbJm7uGFk60aOQ90NrhzPLywvBXa4skXJvLKgJ345/
iLOVcuboB9EnmZ+ZE2hKuTv1Zcldso7PVUiM0/C2fyG51skUepXF9Bx/yPLNv9JypAlcYq6O9ZMP
r/FWklslplVOYr5DkAen96q9KGNpgHh+tPG4MwDfEaPZFoUa5p4xL17dhJn3smHdlyFDWTZVkaiP
dF9LAE33mpZjWJcOjMGAY6dEQEN236uVWaO49s9qXq1lXsRK7xnA0HMrv+aY9gbW3cpnFBFNIfqL
3t393BUvTURV1guG45u+CNMwio7cXUAfQL2dhYrwQf3aoVlgKzu9V/9CE3eLTBpAU/eORo4e/xeA
64NexCzD0mwoyBGtnMPw6xjm+sNWOFBahclkf20r2PqggSxgpx2kzMO2sXvIEuU711pE2I65oQ8B
fsYuDYqN9rGCMRWsHZHYxH+yviwZjJTCOanj0MhwQJSrcnZnnicS4OzVzP98bZpjc98YS6b5Zh65
6S8l5QVJS9a4DQ7WoLdw8ci9+JLVhAO69/Vere0s9kdDqMyOCB7ZY7wGTPLKTrXLpnuNPbv4wDpc
IBegka9O5pTBLxa2sislACkWhBa+a2MA1kCBY3euqXXXl+d989C07kuvCU2K26hLWRXp8cx9FILQ
OyQbKerxRn1s/KXhzJmnOYEk14HzhfzSRZ070UqqLsNpFvUVVmPUT8C/ez6r3OVt8b1J+eK5/5dc
089nXNK9OEPTlCUXbNweLzlIZljZXlSEbU5AQPaHwtZjQlqucx9OcqfU7HLnvpxW0tFgEzSlwx0D
xr2O+AXbvZ3XZYNqCkAHFURAUssyoD0hZv2v9Nz3J5oEBUOSpcqRVl43IxU6QAul5TiLeeOW06xR
ENXS9DX/gF6ge4ihcR4KrRk8nSfkD8WatbDrs9jQtO/P+QHe9Vh0TUrh8LXnNrO4Hiz8zP5EH8i7
3FUgRPhpVNIjW08pKsSj/+mrGFUAFNz/KB6PWwXtbFGljleXDjEgc34V9ENUI131omlGp+qXzA4q
HYnHg+2oAZl9r7BbUrPB3XY6W2B+48zW+Ia0owIU4vy5bkOv3+SPx3i/NsZgWX6kTk1Y2lGx4mPu
7O2yCBZ3aU26bmIt6lMqKQTNmpod2wYbXGtOa6S3/r2cnRi6eVwS+OWSaVNYQwXN8aBQUS95clgi
xPbZACE0rHK4Hq7pZk6AREeZVJftyboTuhYFNuzMYCjaFAv/GMJueLZQZ8kt+MHPQWImfD321Tc0
piiX905JlcOg6to5yT0yS1zBdLeJZWgJWar1OtP93voAVSkAoTcl1YySyntgFd6SV2XaAanIUQhZ
Di7lSupK0yAhO167bAWtvL38Xgn2RZY85jdLC2+BpnR/iIHRRMq8PG8TUNeQogPsl2d8799aw0zY
l30t6DFcdM73yqXoilQyauDU09T8RY2V8D+/iyQdDpQetA7SSYAE+ymzffBO801fL5o4UgWvuEyW
IX/uqxaO3gC8YLPROhC0RFXpdcPVClTPEN7mT/Vjrv7bGOj8x2gEAvLTkA/2Olvgdqk1KFAiQmf3
ohmTIfAGPjyaobVi5iZzrvytbQw1UkDn3kgSyiN7vKJXunnFLmxpQmJqufVjaXwTi6QzzOXiwDcs
xwyaVU10SWWm5UrdcD+h/rPcUWe7arziNxux41G/XqdakYm+zY9684aL09B8KWPunxY0Dr9e3IzT
o85VHLY1wtdnnS0osX0ofYs+1lg5SK3BYj3h7o1wZVQkGNb7AK0j4Dwz/0//1fok53eRjoPBBiUe
RU1TRyt1GFavhv/5eAK3zvLOzi46Yy6TbKmQ/wZcXx5C1kqjgfoJwGzHZKQn+Qvf1tY9sZ5mpqGa
8NKweWJ7jcA7Cwdm9fGTrKXWwzJoC2M8V44/cZpiF4kb82YFCY3aXmZdhB2uqnlnSEvWtLjn5fik
2gsb3pDNe8nak++IiS69YpRDp6tejmJVlaXBycCRDHsFzUhXLAOjiQs3V+rc/HHqHpCw4/TCkC16
cLEyT4md6uVXJrHpaxAIjkDEWhYzcrfBzN4nIrwGEnpZmM84rqSt49MExHD9rb2VmM+0F3b6V02y
ipK6Li+DBTBJ/Sq8+KvpuYPoO6kIOdaINi6fv+dk0G7iXRvksxwL+xExKsMSjngkzwH1c3nGtHzK
P62gTw3bJ7Eb1LTfNhsfA5ZlCSUtPgIFn6lL9uOFLC/QJ++RZu9DxEZT+7lB1f8DmTErVAOGjIFG
ASLTaJwgvND3ZkaUTFv41dC5dPWqroYnA5VaMK1ebaYpnN7RZydISKDCoXqOo3czBl+qiIuAJzYd
a0FSDsvvG1Q6BiwgEJ3kQGFUx+lM0X59Wep6s3dnP5JvTsagKZjQG1jvRg+EJrt8BLt8Pj7TTpRc
M0i8tcxgZah93BcI9FN2CDio3wguJ8pPhKTzHHfAK9wQ5wrgNjKXsJdag4MoS4uy2G9DMgFsJ0eW
QlK9o7EsMy0E9z2oqViugtVd+QORDsGMj9Pf3cJWyrXbHdPpKsCXW6dSld0TBCIJPGuRY4i/a2ES
GXmm8t4He+ZSY4Uj2WpoqNmxMimqyO8tbKKYjG3ZIdzPlHeyeSFn+rv86sTvzokN9/DtYXLeor/T
+mkaSFK6LZX07o7mgJIEvqroNT4tMO3nIdWEcrzbBeT7KKbi/kcNG6EQMdFVeK0BcFZa746K/8w7
4qLNGnuynbItsy4czvgby1y7YZKEfEnsKmLWuozbD+blIOUPnoQmFZ1m1TkG1z5ZQFZw7XSKSPEl
LaX61qQE2jNZY/qJnPqQtPLGrhkngwvYv2NSDer9NGlHjWCSF2piUc4wdcuCDwPS2zxYW6hhEBeF
rDa+N2dD/YHmZZVmk4FGDj1hKsd4GOwFHciiv+nQG5MTTLf6125pNGHzOYezcqOj72HS3NI6KA/d
Dy3LW50TduHW33AUPzbp9cE8WOI3oJDOGQ0Vp1MqPqji2O2l/kFpn0GlHvEF3xDtNSJWgUZyjEVW
yVCoFN4tcfiBLHQuMPei31Z0M36Y7wfXo4plAe3dAa1nVrOHXYBrK2eNmMDQRm1nl+0aomQbD8ea
Ed3fBpiMHjLzM5MnxZbd3RvCiSqyhay/xKfAUGNaFvBi6i904AX+T1VQk+PjOogTNr8rnN3X3sf0
7mvqooa9jKy1FCXrA/bFdQnBR4S5zm4yS6iAvvr4pbSYeFXbL28hnm4ztzVTksLAxS9vm175RqeY
Ze80+WCvT3YvyK6cmPu693rmPk18K0RmcyymX2FZhx29teWIPvPBNbmWUToP6ASTz0gAsfExGedh
x/c11oRIIwkune0shSHkQOi5dqvqvNLbDxvhJYZRrVh97mHKhLM5e324XWDyAjX3TE4H6huV8PMh
A/9wTjtayQ5pF63TYHS+N5OLQhOn7h2qQbppVGF9xKdv0wBOcho+aGlsdGLkCH68gsAWDuY8BoSD
td9yz1U62Sc25jUKQ0GUF7UqQRezBnZiwlUNHWlJulDQQksU69xWm1UwuIOEmeAX77LwuxPJo/ss
+roDhxcQVnlk4nkI63GwNPAyT8MZEe30kwM1x1y2VQaNnbHzC9/Dpo4GCW1ZQrYoDn2mMK3rE43O
H6OKR+1HbjgEgdSNBCEyxYXVq8GRkj4VlJigu20uAPFUYN2/rOvgcS4zljSJ1OXjWRmXIM+g2cPh
ptgqVp7mIjMRQHvwXUSIwhZsMMn+UjygiHIfx0RB1NdvZrOV6HsXpyH6EZ4NZUkJMiT2uGqvTdWx
r18iWaGUZ9hyBIqAOMA3ZuE/ZbEHQwv21GyMxrv7tt6zAjsMdlLX6YFHWgn1n+pkFevTyz9OETKD
6hw0zfRwYsNIb3JN7sE0PTnJnaLGYFsKcwRpM5AKrU8wDM6M0QGAFGF0MG+WMOfOo5pGo+6Y308M
sD46r8vna9nE5EZVInzc7+N/2kZUNUzuC5Y1BxxBpYE10zU5hunph4ZLnhgzfgMJefiOTcKMzGoU
1YDTJTERdb/ZJmS2n2QwrT9cn5uime3v2u/+gwurjOg9V0g0++YioU4hQmtuBxzDQ+LPE+478s0b
MthX5sWnvXf1xwG2wU5TFP0rqLMjamRNsqTqX5mxAuFXgAW3jAQJEPLCq7Gjsr6faIAvBu6yZlCv
8VZaj3ejhBggkxZiMYEvy4yDWNm9UVxkJtGwtZWpZWbPR2UTnCvptxqDbp2iDaxWMJhvpbudMjYi
49dt3KKViyp9QaC3Mj6QKJjS8zldjf32IypR/7JhMJbLZz5Q75Tpat0RqMRv49GCqwjWMFWSwFRX
0XoM9SiBeqiMJ8KWCyMU/RWaz8oXwBAhRK/iYvq0a64+X+P6gUkZ13iA0ATH4MJNET3Vwz6U4ld5
E8XyqcteOA9jB7unbHFjF6OEqcixBp4h9GGKgYPo3q4YphMqFXH2z/+k2XS2M7gaavRvRRF8Q2kU
YIYY5gucVibKf+9NXtNOHLwIkIiDxB/deYUhwZevmGqAgy4qcXDz2h6oXs+PGvaj91Yb+x3YKrLU
Zhig3z5DeCb7af0M26jqGVC1jZU9npg1Svl8aDaE90xzRspbBJ3PPJMwNblovMS+x8PJBXD17NY3
MVgKMCApJFsKCsrdCjTj4ek5Dtg0Z/PaOF6wfDmKH42gEGSWPshP6uhnWB2qeumW0xDoOEyg0gVs
JJIeD93Z1SD1PlBLAfsYDDXUCgdUsGeaXTm7pYzJexu7tkJY04NTlq+mWmq4+7JuRFbtH/fkl/XS
oiZ1mFX+5nE/4O/tuK4N1TZhAAMTEEaOEwCj6N8FW9gSkFQmULFO1uPWWQREQJtxdnCj4AJEYs0m
2sOGNUeztRf0a3n2xqO1Qk+qy1R4BDmophCWQffYGlDmGskX5VLSiU+vg9e/ZYC884iQ9zC3NYca
CwtsomAfyc0aks4+9CehAfzZlxrJVqc/iTwqtu0c4VOGxrEniY2mv2AtBK0g251HmAl09qOWSrZr
zX4Po8JTWoG15fS8kMsuuWMYTYM6PevCYtcA4hikQu81tHbFX4QHHq3KvfTQV9fexmg+UqVy99d+
Y2fPCpyFuO4R2/2gw1twI5tS++a6++ulqVNC8KSFYCmagRGt10DjtgWTQuiPb1ExIX+FV2+0DJla
PgJKPjKNOTD1XobKtEdIDSjaVRh+ea4a3ByottYSOGpA99zLQq6T9paGcAVxh+M4txU1Wf7yrwm4
mTpxYt7gfjFZcaApR8T/6KGXVsEbEZpTUQ7cFLabVMFNageH6MGtp1M0YmlItL/qxnvhAFc2zfHh
xdTcxQXxwMc5TfPHKfK/zIiF3sP7voANK2TuYcMcB1MwzzSAosBUn9fs/tK1caHOPlMmmIvZflJK
gp1raQlGpcV7tEO8RLj8HUNf95MK7leoOAVn7k2chqDx+m9+IEa0RM8JtmqzAuRnla1cA3KtmyhI
fu+oibvysj3b3kIlp/+J8pr2fR08I9Ht257KvYrgWYXYfJyXbodWLevIG60emltBIrX3KbpH3pUg
IP1+WUUdSbgEO2uGGc31Dw5pI8H5BJBch1N1Q7kMka/q/lU8bc5sm4YBxVEkFPw22oBcj3zipU3v
y2b5t0RVpDy1OpFBNwnKbkaorIF4R8rXhLnegZw2lIrJreyboLYv5E3Z8F/7wUxwUseuMXT4mdn9
OgFcWHrwdqrtWPbgjr0EB4Y3s8pVjowUci97qX0Dr4nLaUK5nMOEh0jEqOO2utnG56RpQj24wGQ3
LjCTRbmGNYUzEc7OvdRXlylLPVYL+id0rympOPgpYuvuvTCx6Sl889e87Uv6SxkM/hnQJu8s0XrD
e5tciCKAHbbBlgRZkTW00qSOsYQNeNS/Gx+J8tN3j8XRhSoUrW48xcd/hlPAmLridiMnbggYCBLO
WPtUFieET7kOwFmbKh4/7OSbCKjoH6DEh5/sjYvrJFOp8OsfszUFMHS+Ty/WWsiGAGl00g3/dDSX
BMP2BqiPEwIQoTmHkd6NgaC198ibW5cxK0Lb+8b724nMoju/MAQY8FM3+utTiSL63hQYxO9hjRyv
9hEC8SJCf1WJjNvwQIjQUr3lFhlEGJtIf7bQn7QA9GuZmb5Jvfg11doLXRxo1w+LecZbL8tLQn0w
gqPP0lCC5z7aAEfw+w4AM71ROWnIx/7RAyLcP6AVMaqz8B2FXIz5yPh9jeV/6OGz1cq7bE05E622
BQ1kycmKU8fzvD81oTar3ZfxBv56HSQgBSY5xkUIcX67S3qPFXv1zSN7qL78CVYJaQTLERG4GZCT
Xbn9cKzLNMgN+FeSbL5xXEG65hl8YCSP33VVDHrH3sFW7ElSZFFVYpuiQ4Ibq1VA/wsafo+60MB6
xvyRLNc3lx0m5aAcr5nwK+/Nj1EYhAgHN7dVxuUGRb/75GrIp0uRtzM9zgt6BVjpz/dXbGI+E5Yk
PD5KIyq5zdfSVFMqwg7EYW21bJtYoAK6V1NoCugl7KpjfioBdwtlptSOQM1W7C7bbjJyddDkAq/1
x2kJBntKNdr50V994i3+wxpNSfk7cr9cUo5l4/7BMW5aNVxdVRyqBreUqootMoNxk/h9PZ7dexlP
rUqpTlpWE08C/NRgaBvxhzNkiL8rLjbeDR8vWF8o2w5wxcvJY9VVDRJaVAalKWRsXwovn+FJ1BkL
3KwPDVYxaifhuN+akj+0SvM=
`protect end_protected
