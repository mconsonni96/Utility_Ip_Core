`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
sopS5OBTfEeovjOnsEhUVApgHmBomQDMid6/5nJjyM5DfKpYuOqSc9uHUkmFEQ6PtuIfw/qn4hGd
MZuMjZTPta9Ur+esgQPJxTjVg5nui3mr8KhGbMv7cav8oRGLq+edyj+vtgEVopZXKXbJjV0powfN
Fi9DKsZcLLauaT9RrY/mTuRk2LEUGOiC+1Vv2m1mP99kuxxlPszeI/nICpz5JWio07lY8631uLex
Y60dGmUmyxSX+AG0oYpVHvgxhdZXMxSiwBuqkfWCvnR+95KSSVIY3zcVAe3JzrycOAa08BisuWRG
45kI2s0jNAPbi8ld/1TojtApc8yrq8ECtsEO6A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="0p0GTpxOc+qoqosQLW7ayTgEtzx3+sxwMUyuMz3xExg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14720)
`protect data_block
rFJHlFYDJ7YAbX8natME47Kx9bRSIAMXKsTdF8udlnYy4/qfoWmy1Kq4AG7hBCRaPot5XIJq2/9Y
NxLk03qpQUXlpJmqfvPL4OHJaoJ+H+mmy/1mauQzkaHv7I7nbfuEh9A1XGMWmnp77GjC8zUP5OLs
aV0yIQCU+xiO1BkkZMlnbYqoA0ILA1RbyraL4M5Ae7YqzYYLavIfj2RO/FLJbCEeQ+NeDvwy/8Vb
2EPxDnI7G2KlHXkndN5rOnGETZDC03zQiVHK1BwUh9/xSWujAPajtsgIaU0P+3pUrKuZT1926B8N
QWmj+/ltlj6mQfb2tneM8aTol3tL6LkMqgOxqEefYwz9cmVplV7otGEz9Pmq3HKqdNCnuBt30+LW
F83f+eVDvm+GeqsXn9KXZ1XGGypzXHY4CePjcSyMU95G0SzM+uF4WfnHUwZ2/inDqHedjkst5F4Z
xsitg2Ko9nBqDkxz41HAWZAKgvpqwRRDFdCzR9dBI2/pbtSEwduMKHS/mkj+C06DVDkleQ7YZ22m
YeT6eG6DATCRWCnYy3NGwTDsvOj1wWFM9TQ1eGNl5PcQvdRieZ8fETECj+HzQTi+dyuWKmPGHSEo
zXJVoY9ssYCdE5rIBCsJtMf3vEO3Tzb2sLCjhdr4OjqjCkqVTAVxNcj3RlyhY5wAjnkH653HEciY
YWSHJmgjSwspM2S4Ggp9jqQjiCKLNjwB5yujn345ohjxGO1275qECbdL9NpnZ7OCulHglXNsxNSC
/wL/ckLbsE0nqgvYr+VTaJVYKt9Jpdg38W6MJwBwI7LSdQKTT/nqg3sQjWkVNdxVeXTGlBcB0b8a
ssuVtNPBvnSLHKEqfBuAz6uxtwaMrhO1uvA8QAd04qH5nzvHWFlEQZmQlvoykn3coK1cmpQ+xG2/
l2mDz6W5nyLaUCK41Sur/BEQWKz0EZXz0fCcOzMvOS+HgrhS76r2Q09x1D0Ei8nJ/0EIn5gn3F9d
yEeIIGCFmaoBSS9/09bgQQbY0sH4lrD3zE5nq7LFfwmIh4r7zO9KKKXm8w6CMCS8W4GRU9W3euxb
/w0vCnIqnh0JLLHxRh2fImDMoNySlU2JIzzcQhGgxK8lqPHmNualCnF0bwZhBBFcs8xPoWUNNuqm
48/yg5e2VqJXIeU67mUaomt41ap2ZF9HvKcZC2Zx5w8Fubr5WYRadaXuXFlN/rWYFSiINAVITgh5
zRAHYJshxkgCwhjYZBJuMYrOwhCIl8fUroVByKZ4hEGIL99kim0tRLs1f6Sb3LvzluhKTAHFa2CV
aEz4xJ1PTZE8rD3KlWKQndDCPyAa9LLQ3z+mo/XyQswseR9nMYXe/bZtA1gr5wNOuY3cEMRBnDwh
mxmnbFASUD/QiaBjHCPT0UAEv3rUVQZ/Gg88piTbcWUQnD8sgbpp6ocRU8L1UqcEhvElSOtVFTm1
Tukk6Bb3pUizE4/SXWKxi9NepoohrkjFI10ZFgUoLQ7MoVQUf0MsUhYwvOwrzkvw1dPG4RzZzdSW
sNEIoDpzFTxB3G1L8j5SztgxjR6SJJtPLk9wHyATF7IN6ELuP0X+NfeYBg2f8FC+y0fRFUMEzHCv
1V0NvMlTnW/4hiYaNjTsUNCcZFxH5veEb+QvSvlc+v8bAs/w3SIRgioDlr1VJ8dp+rjbxQBCtMIZ
94pcGeTxxkgRZNTWyZ6SPU4BR7+uXWEk4ZFVCtjt8wUbnMbWV589zdjIWnUhPytLBfhmDvNKGPAw
hCrTxWUKxd/f3mQTvxtDZSi8Jdgf9BHhBUEOI9o12z+DoO6G9nQpY6FuRgxCIoQ/phMTwaIiSpMV
aySMLclHm7aGLFOwueGDEuQjRRQejp2iFfP/TRSvpm2D7Uf/eykbBfnJUKJ+Mzw7mbgTlW7eCI5F
1dt1dhxFAfo/k/wx2ZXd5Ps4ug2JXPihCjvNfTE8tgXp5cVR4TqNZxoXdlzJ4ECHa2PSeETDuveX
xXESnoNojk6LmUiWTPHi1TTjb3yyT6QjjTblaJbXOpETkcLCaZndJxTQTp0GhaoWK1kz2swcHytQ
YKp2wnQ+bnnocuOAfLue2rTaOLJKC1IjFbCL6a28HniwdWqjGBsoOTkRNbkVaLDi4elX1ymNcWcG
s6QuQWZvxn+j+IEIDEd4X+q4S94bQ4IhFdvDFGpbwBu3xtgBlNlTRIq2g2m4PgouLYnASNhzTk4N
yjqswNBlWBkcbZac+Nd4PevKefQ8Wn/eferNdT+nbJsgApKG7pYrENbXt3sLj9uvMk4nBmwz+UVe
7SO6XfztQHWUX+mJIKIyk4hoXhX34NTjVlywurRZq7VNKqeG0deerfplXKMJz00JGffoBB9KOC7B
rJor+NqZeJtCngkanruZn0VSmVo2/8HHKIqEHelGmQkZh2CQuT/npIGsIV0MbrgHjU7TeTIYnU5n
3LSJxeZMLjbs4Vt2850XFACz0RB3OpXkjBBEkfEsbbGZ4xv5Cef0pXT/pQpfSWVdmjgo1aMEQpvL
RCzFcykpMPFnGsdl8m1BPWj1NKUoyfdarL4S11Ew81/Epn+WhvGFJ8GXvAXmbBDK8Z7jc4+/6chK
AneY2M6t6t+EkB2fXqhhVZ7cxUaQaxxkbeor5uPXGuimK+1QhbjL3XcEE95cV5+qM4EgLkklqjjm
gIobHhdXayZIrmcnOVeJJZHSRO6XNJa1mggYSWFn9gzBigjgfiiUb6wIweXGTg9/f2dzFgex0HFW
dxNhW0aYud22NQ3ZhjVdEQlmfrDgbOdusBwd/Ve8H2Nehs645ymNYrPpa2kFoeJ9Pi3P42wfdlDD
j5qDk5EOaQEgbNWXrdCLUJt/fkOOmf5EONLl4MzfsyRGR4JgEI1e8G1D7QWkdyVwODJdyb5HBSps
s+Mbrw4sQZT7mUqv+2Nk7L/vQilTMVpHlKi2+XK0j7p9Zmx/9LFWIX/hK5ai2dTh8zsxtyEETdhQ
yDi3ReFhYnqJXM7bHRBqoPvge+/ahv59yEXxcPPnrf+bnUuEXyDzGB+U+DVSo4eyL7I0gVTSF3xR
PG/08G1MUAbXAeZH3AGWcRue6f4raixyKATLlCYRTHv+uJPMf7mbT4sJbvLjMDpJHYYHudMWjg/S
EiIpY5T7i1CtfA97WtL+of86ZSkMYEsJHP28qWmdtUSRXniVeXDUGMK4fOABSvMH5Lcgjr8mF5Ba
ScLVsf+0X60XsWx3a9ZPFg2wKJGAZMYdhl+BIzKJ/tNFEPo1AxI7oDAwgVhNy+h54Pyp5amFAjvg
87yFGp1MQKcMYhTxkoFPJa/VaigaVsC/ZmRWmIIWSH3OjbG4KqSJ4Wt/76d2/x8Fdysdf6ncbmQ/
KVwynefgjI3UjOBsfUexdVKuqE1Y/+t+RwX0P54qz5ScZCyhFhJy/uiFrEvF5JR4VH2NFJAgK+b7
iYxKY4/r8HUVfUz+5seCaTSGRL8b3sXrEsDmdqJZd/r/iZ/Bhe4xy3LCRCwqrSAWn5JoJqlMN5xO
J2NsItugu/8MKz18EEqjX/FIq6Xcp/uhq0Lp3S4qkRDR64QG+yvxou3hShdMkZ5UBAC10llm1F2w
3i2ZGSktKCAIZP4bEHOsZusAfKz702OJkc5AIlnmEnoGWwW2tOS2fr1t6OQiFxVxcbnP4JkBZvw6
rla0t/iiJ5iY1V33NRblPhbbjmBS3oWRevBHLfhJlbkSEFkziugOUVl1CbkNTO0nIYHw+fh48og/
+MIheNoR1exmdAvkFCzQYIoBaIw1YzVWagZoMon8ans1eb8kgRm8Q22Ngcw5iM/fuBYIb19iQh0d
3L/IA5V2qcV9WRogAn/W+/dqLlQmBQRyh1VB8l2VDPK1kBwA8uucfTb6R2V5eQw0D1733EkiB+WA
JzqpWpmfodUkU6PXOf3pOBmzidkKSSkU/y0z80wunX/EFgjoRbpC0nphzBKzlsuHKzQqUTpWB3ru
tR9aKo0bNqoaRbf6x8Z32F74YvC4mdf0Iq0GXoiGnHCQve9+LZp8ztQ46ysbAgxQ3F/MNI45eDdI
X2mh14/GjCC7bfJG+IqkIb5/FzqlJNU1yd4BLpViyREiO+dm+9Zkousmnf91BR/jWKSvL31GFH3S
yj4rMKLKF/paY1IkOXuJM/V8VWx0Z09zK5Gbxl3lOWKQDYWl0yQddeEQ3Y8gzxjDiL3LIFs0CQK/
9NlFXvVWnkeUlmRgqJfvWfzRY+JZTgaUIbapVWufisZK19qh6jSAGE1fcC44sIJiYQ96DbCmneFb
kOkArBB3eNYx8TSMYBhr3Iwoah4MGY1Geev+VHKUaDMNCoFC+iPz2XKs+x+uTZ7lz4mGYRvhJ3vp
QBwDo7z/cEQ56Y0umHPn6jfHaMq/5SLq75ESEFx8TpqrMlPN0JaX5vdvKiP00v4nHXc/On3FE3+b
XcgXtO2P72ZXQn/2lxsD4Qi+BmSuZ1bvbXkGW2QPluM+p1kHKrO6kTotyqIG3mPgdVvPmRg6xTf4
ZebiQ0846fncQooqyihi6ufX49ikE5SYQ1bZBwUJBSgg4UlOrLBSYKSW3zcG0iBT6w2kevpf8d5g
dSH87bwr2EXnCLMy7R0rpvoVk1YkiXBkK711Kv4nKPYYPE5Umc8Pger9j5DYK6S911FXhm0wV5ZZ
IWJkJllrp0L6lsjBugD78SB6Mt1BfDZWDLnFSTwo4ghVGTCPG5I8zEFwTzfcE3O4/BpDBiF0Qtzt
HInuHxUzLxLnAZw/llFMcmDSETeVWYUzuK4+TClwEuhzM9PxqLiIQIp0W/B5jjm8apQ0G+vFSKRV
yaqDO82x5bjWv+rllkuR3aEoqyEfzMvx/1bITslpn7ozKUNZk1yByZHDHqKIU48UvZ8L6G4VZhXI
V3svRI8IwtFW8KSqR+PUemtwKvDWImWqr6770yVEm8HxzugpZuX8hLct3sNIkvKeMSdoCDkKys73
zf9KjFBIPtgdo0GL/kI7HpEPV6GRuBAg7dwDR3g2jm7+WKnOmvLZYJ2kjlSIGLwiV7T1k9ZqxHoS
xf0trS+aohgBRaZjBOhxi2kNwSt0O+xx+10SRxk68zwej1O9NpTReN91E8VORkGuvxsHOE3naTi8
b5cTq6qEMFxZzrdYSt/xacMC00XPaHejw14AQddDa1s4xVAwp/1vMv+c7Sy30m+daWtDY9AS2/ia
RCg0YzdX8lTN285Oo0xh4nzMsWleTwTbV8VfYPEqAf5DAGBMc4KYOG1cYSljAF6+X1ljul0+i2IJ
+ULkz0dlK5Dc1bRWzAbRlFTgVtCvrc2zI4twNcj/28n7YLE7XBmNhDnj1Ir1oU1ueUnqHpYAtsRO
AFllL28OYRhd59sAODvlOaUlo92so8Yiz04d0vCvQZoRNdrjjAxSk3Sv7tYU0yCYtpf8nTpX1cMT
dtqb4TRAFaMewj8aeYmeVFR59dXwUsAx1LWcT4AvX4a9H90hNnamnrZr9GteQRSdaiidBXYZ786n
aCUD9YX2Hki44Qazk9D7m943dYxbs8ohi+t+5rRkZD2vODT/j4dn/k/dAgrOk7wmOvFRMHRH6dCg
GDLvP90jNn5QWzuywWOnsTL0lCi5jYxMikpUBtbkNCHzCMsFnmqMFIfwAimO7+HaCahjVvwLL+KQ
RysN1EO0B/J0FhHq/Q5aDlDAJqUp4rsR3jKMrUvZn/7kR57aE6rLGk514Z4/v76B/Zc7ISVpqjKF
8Q39TOIt23ySEqG4oBd500HaObGICbxWYzBXUiL3PfylXkCL0WXniY7azhkSZppMwoUtGn1MOuxM
jzP9oqlZtxNCankc+58ieVpt0qhZL0msqPrWMxb7QmkjGMJGI76QgwcVSa8cpk/l2fg1+xPViWML
RjV+OKLFeSAlP7BRh38R2B/3vbVEJr99TKgHGqfstdfba+gPVCv2UvemLSxEiz8gHUS2QDRa/HUg
YojGAAdYBj6dONPOYUXzqTsx7faytaB5ohHCm67L4er020A6VwwVQBp4F0h9SxwfApRblCf1uUvn
KxCFza7mlrx28VRnmhw5zFdT52xVLEIGHs81QnfR5Xsy8Qp4LtycjA3cYDmUoHxug8m5sYaAFZpB
I74WeHeaB71x3ZRx8v4wBkoABbsnB3excbPvngNNO2n+30SrPQDzFu7Ihsi8Lu1SCFQeNBp0kvRY
hAQGjaeboJnmvE+4UsvXQZMhoZdANCY0NL54oJM3aG4z2VMFBHn7EUc9dMR6PdGfgwcZoOxlQVHv
qvigq7ZbBufVA1zhFwVZvMRZUb+zTgoMmU2bF5d5xunCV/VjWClBnu9Xo3uOVPK8u3hmqPhGPkdi
/Z2nVhm51OmNGbkZfFbCmG3V+DFwvTufSnJSExajyrJ4QoXdTStuEiyiLF0HQ/JZS9+gFzX2fU35
0pwZZzUZHFNpR7vKwfaFJcRyKcCMNnTb8I6XJmUHFt4s+seAYWa4Ed9wm48zNqZVaHY65JnzGPzu
Ak4QDBWHxGawbEK3ms1vUlopPD26SxNaNDTwQPkRLWR3GEefQWr/St47UopdS9/Rjsvi/7q6CR2B
O1MAWCWge5X+fDrvZgQG7rPR1Zg8OiLIpmiykGGkJtT9wfllZTbBvLlaW93xrX4aBBy3G/U8kR+c
g80vNhk7gZR8cI2Jlpf2TQh8hcB5JEH3EaX0FuuVl9RJk1BnfjveFFZzVUcx/94GRsfnDeZjXLBp
w4QBim19aqW6m9QkG7hkIi0WR91HmDQcOC28v7k6DS8LiENIS2oXOJBFJGeM91Y8uh+CFOjpVOY3
vwpd/VWIUMBzS4/JhJbdOyQPPzOh63fLirjdn0mFzFJtY8zTKzKR59BAnWY7wCPMiMOpcnxV42Td
WWmjPncfcaazC1asRxKscliiWEqjaBJs2u2oyr13+J3XNH+ABlZgVqgQ5c2RBle3x0nD53fFMKqt
xaHNwwuBnd4oLit3BOFOqRwBQsuMg6QhI/gi9yFjh88/XO7nKAvCTu3dpgYtxRFn8pkyM4qXnR+a
kMxafv+NaYFi8XH16wqr/U2s3Nhr/0BeNUzwjsaZAdsKc0yamGisTZHR8RY/eY5TTHpWOgot5c/S
+4BFombwQUx2JN2jSo1LtUtkrb9N1LfbxZ4G+O/R1uVTnqczrZxJOJ2eMOZj4OW/9d9UBGWQp3QL
ts7bMtMA15FrA/kV2l0EQlPGjxr0XBQ2CY11lXdIs1UBCeSIftdrTaLNHzHWstnRTE+lyU3nZnAs
GoVjCkqby58pWZMPrJ3OOcM5YoiUcYqx99PieRYHmNKgI4ZG8T2teBjoSPhDKvLShsnxUMKn0wh2
cgczznOa4/K8CCcl6NkjHj5EIGi2YP4CS0BZ0vI/gGbC7iQC+h5bhCmVwfVm2AvDhDFgCD9Ukm8T
Np+77JeEiwOPHMMShak0HSF/FCZnu1GOVZ/jjurA+AQsH+8p41DcCYpaashtkHXXsxxgM39U24Eg
IOjSZLdVhzijQ1Q4H505NigVmi79d44LkaQZIycDKnod7oP5YdtiiCyPlUCQpq6pwv/iWDIKnH6T
VT+WyKQxwLianc1dev5mIl5Bt/l5SFfXywaDDO2FeH/OkFXWBSTTLxyAVKBmO4oNNhH8oJvV41Y+
Msca+L4gn7Wld9sdpxfBSZI1oe/OmWoLehfUrlUhQJxlTqi1U43bokKcrZ9muFfVFJxNHJ/m9I6l
hN/fuLl0LYXLX+AYrOyx0ZdYXkAH0Mj+QE5x2bgzTNIzfHkFYO+g7Dnmbqkvl7XefOKQo5eMZCUm
Y3ppFOuXz5AWVJDSpdyDQxooKeZgxu8/zro2VC56saXJdSVG1MxBd9zsMlmOdd/NTqFBv7C5xIRY
Qt/Viy0hdumd1lKQ0l8VBWW48u7vFhDvOrjvk2A4+zEZ9oyfoiQURXWGjsUutV/fqoR6evbz6V6i
EONHq9ExcqPNPs3MFi4ImM29r0G6AYVO1dWeWw2HJftFDWIFn2sDIkdg0cT2276XwDUN8htvAmUM
TlROfLiv7qU7xZnWGkReYzhoR6DRCEh7+tHDBc6ewPrYm5uBaJIyKd7zDoY3UfuNulprrET7ig5J
HLAurn7aMViyDwwjlu95gsBwdmUnvFvqfBMjDdyYggPWbY7Dm7c8mcCF9VPkIUJsZM1na8d7PLG0
sqerdeez3K2drTXrbwqAWgNuDZXV8jHEksa/WEb/qQMm/9k3D0SO/f3ZwigdBvepNGRlmY5IK5tT
8yGkFSRKCa8BmiLZbsrPP2u0hFSWdISOrnYK4bQwozGySMcs7D26CltGZGOaBYzyPcoX8L+D1E7H
pyFPZ6rW4NhDFEUeDd9jqA/Z2VjXJQWhiSQw5QjPE+IPf7wD8gPfbDg/MCea9Sgs9HjiLk7pYzRh
WTw68GaNYZDf20nKaKDxdEfVuLmRFqR7O3p5//0ZN6c3yP6mCw2j5aYRBofKZMLFTVnT1Agx53qd
S9Cde7RcWWS5VVsAA+XJyI+UuNxMS4eUPnk5sze4TU3FXQuz+VvOfyCg/yrQmVBX8CFhZdu3RZxy
TKNB4YoNf3FsN/sbwvn3ev5l3bSaUxCBsZ2Fc0aDJoUN4a90FbUDa0Gno7AN7xV03POYrjrthM7p
+GosRXjkHYnf18/S+lL6PXHo21os6PKV4dBsU9r5FTLwyDKCK+AKvnkfBWjfF0qcW+CuLRrYyPFO
xC9iSCcYOVDNhfzsgq2ybdLHieH5nPbi5WGRhy1iuXAyktfLsB4hRyeWDQa9u6f07oJVddDQYgSc
41yY4OFQrP5YyjwJ0Wb6ds6QDVSQwyo0VDSKOXDYV/mqxGoKPN+vT3IORaHZCBllgUt6vr72r7GW
2ry7KNM7nqK7wQDFFjzVGFyHPVDXN5ld1x2uTTRg511scsz5by34vuWOJ/wUFi1ROMPF04tUt8W0
u6WdZs73DA/Fx7Cc2qrDJIpUucs1JXLaJKUgvy+tauVrbIp5z/81ZqiJC5PnBZxFlBvxNBkTxIYd
RmC0sntmJLcURMmDbbfJFktHZ22DEAaTYivVDXqMmRaUJC/e5yDxm6jrQIuZ+A/ZYosjvhO6AYcj
JEe9bXcMvg0hKkoJJEucOdQ4lkkw5QfXadNmPZZ6BfmkDH4hr1T4oaBmYDa7ABg+ISrRlNLZpVc+
I+ieTNsfQ5dlJNFtaE4/BnMYTZb1fMPTVkTRmUs4BJytYwzMbDQLRji638SD2IKhcUJ6Q+36lYDk
AO/udEyMAiKNaJDPpLwh9UehNNWrBPpbWYLPa2JhwXBP1j43vwo5dyRysdWKWZ7/LSXLLRhAc1q3
2ERaCQqbU7ZCtDV1Az5U7zGAvkc4cm0t8X3YL7HTMSCNwwpQ6C2BRbJ3kdQV7wMSMS8rDIo6rjje
rD5pWBHvBVBN8E7S95BlyVPZ8bsdTs4rDgdFaYtDLkT9a09f5UcnCWWURWOQga7gy+wTi/n7stBX
FKZA8MuafQY8ejdWVLO9JPndn/Y9+t17b3OSSMMWbSS8KlnzXGaCLeN4WUi/Hd+pZIGe+1KvD8nb
5JFCkpSeb46Gr0l4RgtQKgiAK9FjCuml0Fjzt966csxBeX6VJj65/ck6lE3l7GjHIO3r9hP9t0S7
hHQohzfRbLYogo+0G7eeQahtKSfvZcxj/XpHucI59yk3TsoJqTTfnyLUpx1cQekE7aPzFQSCmyLv
/fD69aoSCqYmtOoxiUzrNtVQT7nbvkGMuqoCmeYf3x69V2X31BM5GPXcYaTBzbDWQtGPkbi9TRfh
cBGvVYMJp72SefxPv8/FfpqkQBww97aHWOqGAmjNXewtnnBhVGDGBdfbcPmpaGUlyIMJFJYhb7xV
T4K3Khcj30mTVRthrQ7diq2v4xzJEASc2Kk2HOzzgitVhhcNoWJtdImTHUpbetqhOrLpaMG9PIvs
6jTCVdws3ue9XDt1NGdQbctWPVtzYTFkIx0fZXzzsPpJ3HMhmP1UPIl2/NwJ2MBCZLbz0hNjtmz4
RAURHe/kXXUwdjDIB1SYA0XcJcXDlXE1KLt8QZ6EG2+fgaZ8QadEqPet80goDvaRBZBqvSyWaugT
AOmPczuuFB8i06KaFNoPg8ne6RE0KoHMpIgP+4ynMBMEjktCh4IQTCNc7RZe684kkQeW1NL2h1F6
TP2X9yAeNTZhACt1gPUyRAo6XcDGv38fkaMfHjJ/99Y9VEnFWDWHIqWMus3HzBSESMEpLaOOqTZm
AvDqowleLL1droMxpyRxYcmou5gJ8bE+0gd+cgi1tOvTEGZvaJjFD5KTLgjYD+l9Br6CkWE+L+38
x4GHgt88YIpsPOJli/0Ycm6W7YOVIbjKqUW8c5YeuMySCgeuPWf7n4VIunwkX4pCI62/mfPbE8AY
eMTOA3CuEJFODFXizpBJvco5H7LVQclak9B0EfoN1mBaT0tp3exdXPUShtxO5CYG3mjHXumEf6Fc
Xg7/SuloHjigdpVMorvfCV1ixpG/S4GaHcm08h5XHNBpDp313F3/BWp85KkzJ9pWejrZ227LDa0h
lfvL1bh1cmIBov02xyg6BfFKu1v4dErQSVEeIZRZIO8rGPhp85Dop0KOye98s8Tigp4a5JtXrjAP
B+UrBYS6IwM2UU/7kES/FU0ebcpjtCfd0PyXycITEf1vju2UWakt3pplnJ77Pyz4zrCbv0YUr89N
4cSDK3qw2HhldQOBbrfgKEYtDj2idXjkAY/++FAf7YI209TVfriR46CFoz7vjWhir6lf3Tzkg0wl
Fpmg7ZgI5eOnfdKuLsgE1pYCs48JiaSswHTUtDej7dz6pnO3TmKCtQv1kvrThhugpnRmeP7TU/sN
xulvuFvuy1YgcvXdtGr7YwfQ0rikZoWxIJoegdk9g+AXAjDcjZH6KupsSy0SaC9OsJCQD6//nuEF
rTd3Io7xUuXvGrDJgrA5eEwi8IsBb2Uv0BKi495ZgOiib2VjwfyY3GgnR1gyshXCntZTX2lDceth
8E527qTUuT9O5os6Pw31LmSBbhwuCU0w2dQUhv9wgetz/dRbnYQY+IZxWJA4WYDLXp03++lof8rd
jjQ2QzXmQ06VKQN9x1CjGkzFTrMD7Gx0IIGruhmeIKZKKqMDzP6oPsKGsNurTXQMj2hhADrlXuiX
4dvFNlPQwNVP5v4fx53AEr7adgyqZvHu1JhMBb1jMN9dVnlNPB05oYnq8vCPvVogyQxabd0J0Egw
yAukwCnFjy/04ckn66Ms8vaV/k4410Se9coeLUy+OxUQhlNjFsjetPj1tO2i+NSdPWyv2xX5eU3+
X+SbSVckRFMVD4Amx2UWNihb3bsKRwQtk9dBx1Vc+0TEkPm0jEEz5CtyGOHzOs8KOG2wFFSZNlzE
9Fdy6xA3cBGE8olr9TfZObcnfsDk92WWb5MnaXkDJ9ODDDFZ2BozU7JbgIeNZycR3UVzWEBt2BKo
XsB+k7BtsiykXZBUwoeB4KV20qYWwvNsOWGp70NZNrvm3+4dQicpqtM2vkCZCwzfUHWdTpFN8lyj
UBC3PJ8gru2JeNSv6QAIQd+zN8OuncTxFwfXEg7mrgoy2nF8bqt86eqhEn9/gMwsoiE4yVlktIQI
cA+ErBYUWx7GBYH8sZ54xLf4dCY1zWzK5Fi/YYwrCrfP8q9KaNQeynYGnLfujvFWGEHyRKhyLaQM
kbmCvf7Ms7tRPHs9ooTL1yFODgvZBHNyDYZpNQHv3zUo8XXAx1zUwymUYd3rFFLVrPJ2VFVmgexd
c6KLvyTzOXWn8rdhwV5u9lX5V8BeOwU0gLq79Tp611d4LhlFkJQlMDqVb948dNNYDq0+n31PSixq
BnZmDEWjQ3aeRaMBmNYISbTVYwQt+upjCNjGANYdXKapmpX+6pJxTvZaL7Ge3NZ6k8HSQ2HcKN3g
TyCwdguKIwx406UnHcaEJikduxA3aNfaeWO0Wwp5f5YY+HUUHgLVifRk+u1z1x28MyoRTZqeYRfz
oGeQ/YwI/821ch/RPxfD73IdMKnAmvXdzRP9qMf3u1eu0t1yI80LdToWXL1w6W8occfIQDTQrHEB
jJk+xqySjb2DvTE+yhswBnoTjDfNCCAgdt43nn9FkpnbiSTnUkcmuxXtN8do9INlDxzZPgzDg/EZ
nCM4Hk1ea6K68YnIpmqqZln1LI5fhkjHtYg+LCQ4RvQIvHznmBRJuLaOZp/u7suIhRMr+/ZQhgVQ
8gzkRfn2lscCjY1uPWLOTxVugI0INPws4xOnsLuwfmriC5f1h4cE5FDGbDSCQTY/KyKzcbZsmCwS
MKzlCSZ4bTgnf9F910u7kiBzDghX8hst8eJosYTK3G88IIje2bQVSZinBjKEA+0P8MQ9uMex49Fu
n25CUvWF4XmulGL+3r6h9nbXWtBnoVGPxqhY1+DmlBZrtwyF3UjImTDWjxKzBnlOtk9Ih9XBY8x8
3UpZQtONqyq6XOBwU0eQiDUN1iFwbnJeLjyYhz2bu4urqCHQ8IVowu2Ys2heFMYejLNwX6m+E1L9
HFo2E3VhfMdUVqSbSKeztQU7RFGgsqrlGC3IQOZ7+M2gNwaHU3y5bFTdUm/fBrtWqk+ujtI99l1B
70a/DgKnheYwpcVl0Dp07zeR/cyOzuzhrAAN6u+nTal4T2mrRA9Pc8mzTNAUrpfn7wUPjRU9/Pll
qyXF5lCV8/A4AIjDO6qmmn5YO7EvKzAhUskqwXdlscy9g+ynF9LE55wHpfIVr/rcewIemo5yQaed
/S6NrL+CUoRZueoShrFebemQj10JdE0Ycz0nAkcY/Jcez6lvn7UKQ+uSMO7cKBtUsxU0pdCi3AtC
2TV6nsvh+MaFjAdfM2kM0APhrBV9D8ur1446oSYNFuVFhJkiaxBuVCmXlNLEtXRtO56iBrghByKE
h7vsQYzLHvvJrbq5xs13bJdCCalCi4uXuxLrzQCoGuJwVTzgzNPQa4Rnf5320omJRYq1krxFiCEy
7RhQnBWcIi2zBYAJFXYmNcRKZyQMVmtfxJZmzeKO/Z/XJm2sqrh28UK4hL23HhE4VsmpYWEMXJjn
eaZU1n36FWUxKXYckZwHnBFAWAShqh/WXlHlay3FK06v+G+73+YW52vaAIpyduyIbb5PRW3q4Bao
fbisEkX0kKrUblzpO+7iZoL7AD3WDmKstc1J/6NR8Z8vuKkmlzwX1jNi4mj/88KD2npLsqpyAqsy
V8qD9qOuD1rDDb7V4bLudB7ykn+23lJoucM22P5nBwdgGso7pa1Tb8xeKVjY7AqscT5uihH+pBOp
cbvSjNrPrlIDLB1+VF4TMMEruD5d0AnfzoTEmTVKOXdM3ywquItcpaR2ceo4NgiIAPR5pQFV6WbP
1CGtIU3Fu3mMl09enLFZg5TawQ1ocB2OFaXaMC2yB4mWqkxB7h1U7dMp+IStZPgD+ZpKir+6d+RS
NF7UvXmwr95Z38cJhSEfNJirxYrOHy6EXhyDMnJbnsJK7GQI7tRa9CEt9Ebna86CUYdQs0cKamps
guozc6AO1jlTHMw/eYJ+YIRGQ5USjYCkAsX6Ld3UbdciV5Pp0Fs+YDigmDxSOQxVg49LusXH+O+/
pYa0VWokX9m6mU4cwgkGysbt/RGdpSEfTEA1hnGi6UGCjHLYVGO7T1GWBFm887A5YRal/EAC8jVH
YBgRI4vvMJNpH8cuzTxnqJBMk/huo0C7Vh97dNOqhCq92u9432FZB53VdqI5x8EcDeDfztEVdRkJ
/fMyhsYYfXeLIdpS3l7ErxCMYmiO1D7dMF0M+lKn4sQ3m/40NAOieOCaQZPyxOmtK528Zn0L9INO
D1AXTwBtBy5iAZTFP49QfMCFQmjYLn/ld2LwJvKR7JjzC4S5DN2tMLqoypwKOv2ARDyU7gS5Sj2m
WZ0g5+tkdLUVFxy51u6EpToYnqKn2FekHw701KCMSVtd/Uv3UxBrTecevIr06btkjKyP7EwU8ixj
JypjRDdnIv24T8ruzX29XrE1ZIsyhEm0XzX4Fb8XYeuqnM77QiCDqNSA5UWk6cCQdG2kczWP7qmZ
t7cfxGsY6MGU73qqSwqAKbXbb3pw9FRPZcYK5ln7DnZqP3OKottPJkcvsUAd8o3v76kukNIAt9DH
mtGAocx+FNfiSTn0ZINiQTOgwhThoVjBYRW6i1OtTSGvS4QRIVsV/WQabHJPgU5JCOnVQtlXWje5
afSX7PBczOBrwzoJveDBgtDnOP5z0lf1nXZxjKfFyuTwjh1brUFtYytOyp1yDbgsNpXNvp0QONBR
w2IulcnN1vFISja+tG/a0L7uF/bIrAmdj6g/GU4NGZt5hrqpn9zbDxp7J30OzzMbpyfIuqSovuzf
m+2Ci3ZRmgY2qoQOGeOr2gnDeA1dvnlecstq5vY0ciOb1W0+wg5VyQLu3TeEm7usW1IInN4fRvgU
gz5ixRzTIP1RWtu6YqOKAZkZ5FZKO3UfQ0q2ql6ZHiQYMOGhhpGXEYARQvozGnlmpGsTf1Xc9ABw
Wo53gqG25EoYZTHNktTN2wOHKq36QATvjs9cPrrVI6Dg/iF6Rm1DjSRqk0X0Jt9E/o6OkRncZHca
M29HnEBbjZH+h76MqZAY5pgTxV1bsSD3YNJ1QkXqIV+PMthEHvIIk47HXSZssi32NjjcNTv9RpeG
2HGINMp1Du2E+iSc5UELVxFcnyp0ofq58UBo/Ul9K8qels8vTjTQ638qqGAYEsEEYLErpbHykEF6
KuYfm2Brm1La1huSJjYwCh7mXzSzhFF74ICXZeUqAtiUyZ3Vwyb1Cs/HMjOTrXXWn1CLK88UdBFX
htrGm6uqvX+XgssXpY+qSF1hwfEO/Az/KGBgon2frDkCHNdWelLJ1xCtcWa0PVNjHSqUgrUIIA6z
SDEDWAvuofSbmodoQx2uWrlD/KN+GWlsH3FBiiizmhDAaeQTK8HwA+Y+xk4mqgdwuxPybE4kEJgr
yQ4naiAhSR/p9Td3fyo0KPpj5FDF4wibOjS97yCgCVV7P0CKBtT4OcCzabEHC9Dc6cOxnogE/Ged
0gBa14Z3rSQu4Il3cN7JiNmQTXTED9bRP3ZwgylNxj6PgaVmPkvpv6wn3uJElrDttu2x1QJ3Orqq
l6dEq/uVTcJ6Q/eQJ2vMDiMMXBZ/kRl6GC250VtNz485sook0bvFn/ulLkyLm6ih4P3u9gL6losL
oQEQgeogrXD68Ouq7Nm9jW6FCVqRjtjYvRneAAu8JSdiwzN0C0c04tDstpqBq1MCWBgpBCHi9cno
b7M6R4v6ENGYGrum1dz2IRWDsXZuyhNPRGfULG6wecAfxfmwIv5n45+KcWNCdLuhDNZiPagtlSbW
l7mu6w4OkOjUWSMSF7Kd4vZ1KrEMOYfyfqjHtM9d9XYpTI5yu210l73Qyg5IIQIA1cbiBpRKBz8r
M7mfd+K4dR+2p2lue4jNNWoaTzi9OgZfakpO1vUkF7uYEASysY3SXOjamBbYqCyO5z/Z5RhYWnH5
UKnkk7HruxWnlF2l54j5SHO+p2sSWbMRWqhPF8RtnTO90iQ8ehPWsycUrSFeivBGDKxqKpWhcVHL
NgB0PiK6I36ZNKYpTQ8PKTS9AV5nNDdLNeNM9oZoEUKILvsFkfuhJA8W05sKE+M6cfHH4CnJQoN0
FW7/DoqQp8ycd5gT4YRYltUn0ISqmx70JYDwwegXSMYKuGQRu/8TdR4YCjQQHTF/+GmnaOB85Uml
RSAR9nGckRelGRWCRuMiDFVcE4mSnQnH44ppvkBTPXt4/idOb6vMSzCjQK2QrYXkIC/wRl04Qyia
HFriJRKSWzcVISFshODELLl1EVlDnL3/1DvkTx8OJ2cJf0iIFNPTiA0NCR4o7jmH+3TsClDRKDY9
UuZnkv1ds4F/kpD9Eiqr+EP4xzA551SYKlS7qShs11GbQV/2ty4q7vqB62enIHhbm41Ke1rrlnzP
oalwr/rqPr/YKj349BRVucquC9dw7dLLb1T2Tt9q6asXqlCLURIC+Af74GUjhTbagpcqlkG85rtg
lXC604EYgy+tfWJSRV3ugraAE8ukj+ImkIBWEf3ZHwQLR1fpuwYgzStxMY92zOga5gBtUNxF5M7X
Tz4j18TmCQnICPyyFR4B8tyhQ7CI1uLRUlot9+hrlXyRAbYwSfsXE8xMxNVa2b6O+o9W/n+KXgHS
+CCxoTvXWM+r/J5p9o2n9usUv+m7MhKRH7krzufLNuNdhs/iXqsPP48gCm2XugGxn+XVXnDdfN9S
SBUUKmrkkk2+u4vLjrO/pMo57KvFGLyVfbXnkyyNY94zD6e7WocIUYbsJ3XDsmohE5iSavDxz6I5
PHliN3VAJd7w9PeeIAkxsqGJtNPeLWBsmR9Nt6XZ8Djspe8GbUHabYVVP23izvLj3ldp7aTJ6rrz
NsmIfPmqEn1579kOkp1IcMCMk5L7isXVVi/9QRnR5RdI7n2Dhy/cw3T12u/K3z12rXWt2KvuWYDz
UcelgMYl1fIF1lCzL2GBqoNGPrpJZRAiV5PisauXZVmKX7HijqhbxPbYxZ4RBa0q5p4opKYEvYu3
3vaR/e5dyc3sCG5vz4QqB2V9IJhHT7knhMz1i94iTZyQWI/t4nK9wcvxWSN9s6tUlG7ps+vjiRyw
Uq1XNGlxJIOtaq4/FG9+4WYMbRm30+Vl9j89TsvI67FQLvXXireALsgZHm2fzAqdTqn4Aon+EhhC
0/aOEfAEHiZ4O3+gpjbBbJzfeJakDI9kA4TdmEeiRe9fO4fqKWc5hCVOqZ1gyYmaYdYbo6XK4eKk
Y6iGLWSGOXJFJVMBIsWKKyxxEvSEH7OQrIyDpA7XQBEzo7b85Z9eMY+feeqZwwFTOuki8A+gTUtI
Z7nMmcf4RH0zzdXNOcvbpi8LR3TOZT7t1x4iYHfGfbidee5GML4kNlRt+sJpy+G+r0Y5xeKRP5HE
7sWYgqVKIcePvnTkM6g0ZYLz3pJ1tQ+ov3siAo6cWsOMuSV+Ymmp9NGLq053gcxbZYgjNt8mY3J3
uhlR/UGYa+wAgUesfykl3s4EAhen3Re4cRbKG8uc8XsfTsSf1Lb8mJnYsAnvC2Jta6uIPMp9pQM3
XovnN5WFTyi4fprUMkn5s8aDLJWTLWuPQyAwBzSgP8eieA54Y5PL/LLt3UnKNMNDwbmx7XKkhccF
V/MKS2cKD5p4BcnYyQUh6FrpN+dXRzlpOQ+5WD72mZCh0y2spr+AwBAp2fqGppLkHI6PKMx5HUaK
WYh54Sde4PTHMTfGpsM5exPSkFMdc7NFl1ZjUPkX7UnG9KOZg0/SCLAf9JYclresMZjxO1w7F21o
rf+dvRC/5IMq0pFhMoS9woxE/lEBbS5N6Bb/gZr20XuIq1UVpwz4RLT+tx5AQG6oWzUdix6AZy2K
oa+5fuYqS92HPyHOjzLkHEh15TxEkr9BjxNVdzl2np+0cMDf3iFxhfRLAFIQ6HtmiQ7oB4xgDRwU
/PZwUNqfO3lCeTJedr2TmzG+MqzYID9nYZvB1bOGl7xrz8f3gTjl/FciBMvkoDU8UJO5RE4RzUe3
RP3xulplcHydcocvQv4BrjhULBFYnkqchYmS328AIeE6R3QTbieQUgPSoZbKDN++eh1znhbDkkJi
Lju3foW0eUCbUk2ehoNJKFPL8M9cfYt4MHu1/AcPMs7GrChY/S4Vt/ZPC5h1ySahQBCGXP7vLBFs
2Hq5iVh/KuSg7aO7ssJlrR+2Ob6JCjeurJeOJcOWn23Vz0Xsw+SreJNoLdG6TQ6yZNESnH6c8/ET
eU819DHlzyVZV65pLDFC1oHnBGVJLnVaC+GH+LilIK1lx9F1ksPpoKqCIvu+B+d2UlYiOcZtn72k
QGXalasmXAjm9ffhUDJrVRz4XDi2sNTo3Un2tDTlcAThCTWNc5NiC4+hq4sIYE2gydkefHuYP2yN
5RlWX0A8dbw/K/RmnLA0ASbUJJ4yFpnyCN2gJElktpSFxmvcuUkUZ9kANlL6kdhjiy2wGcNwrtkf
tmtbv+c6TpnLLp6KPSFNzUdIkg9n+itwh2Cj+xvwVCl93icmp4yLcYWvWKHWdusLVe6tj92Vkisc
cFoiobOqcUuX8+J7khQytdYDijB9Fyd/P+CIzNK2YgWXkVQP6P/0VpQYoXyJn8fDa/Cp2EebG1T1
yi5TrxsmO6hlKKsxRAD0O//1Zp6MWnwGpLtAFXyFzJgqDuwSaONxOdM0rmdJLJwU3n5+2G2v7EWN
5+3YSUKv/7eMsGRsfFsy3XTa97mIsRAFjHxEFMEbGaL9K9F7JpOmWMpc5DNfh87d21jFNG77o/pt
SFQeJyUivDy7Xr5XM5/saXwe/I5m05RA3XyptzzZmYJW/lVCcHIGEIZefH69I4d8ToKf9f/l4y/9
TuGSb1icrphgwC8iepQEqsMr5Ia9dU69P0TYpx+l6wI+4/GCacqmzm8F8Rz5AlbhPHQS7JkeObqC
Rru1uRIVv3VQxPxUoTvakOxJ0PJfBcgnIRQK+0iKTjzlVdU1WG0PM/ztrbgkoE/sg16NdwngRq/Y
6EGfwtIp7KZKUB0JLEubj19MS3kJUyJXp58C6z+EDUwOjn47Ib0X3C2jUZlkpau7cNUuYsuUpEoh
gflKnb425sNSN66ZPFcuXzqWLT5nIzwg/Or32yN1pnNFe+QG7vpLXBO9eiADIeE5pNEesRhRFOEq
hIY28qB3cepxP10EVzmqzUx/VAv90J+R4c/xKAcRfk2Xq5RRbnFr4JScQGSyrZf1ew30dI4020/S
d3elUdDgDHRW47ZCe7WhmkzkK7k6uzLIcHDBugEqEBHHO42uJjSHwDpe6iKkg2NeiXv0trmXY/85
ZVg5WkFkf5UYiTOrG8rs1gn3M/foyolL+0EAv+vmwwq34pGp/fde1jXVuxRK6UwSRzNRbnyY2DgN
3LIO4+M6hUPkDCsDAVsCvB/Yv/CpnFPgZM6uVoDTMWguFXUCmPUCaD48qEszcx/xavfR5UD9DM4Q
nIIqyX0vPgm/Xm8FnRQa70UXsw0voY9PEgZovPe3fPiGje+hB/SJG39LgTyxQE57r7nfREvLaHyV
47oDVHwIPcs5WKZymZhw2zK1K5FPzK4eYgBn244LGys/Ol6TX6Qc8aeQq2LAMumZNcyovSv2oiL3
HGiLKXCkxr3TwMgEhmmFW+y2EeQEXV4pN0P1mjxhddsHA7xg6XEfykdIJyXyRhnx0XIG4lttE64T
p06nQJvvU7KzYvIebO29XQbcpA//cIFz3WNH1AmwrttqkWnAmCdK8HOIkN33Rsp+GogSDg0frQRt
y8V5fErS5z5O/thLmUivirxRQPgDQTaykHeesPqB8uCgf93xTJUWs/Os4xA26IwoGDAHY4Nmkt2y
mLFqq0rEQnxj6f+H6jjfl9Pyv39BtIT8QzbM2szysOacAeBhkq5F0+/QozNEic2DWIgyDgzBRR6x
HbKh/+zK7U3pcfi88VaPIc/a4NmlQdW+xzR16+c7TAqusqANv770j6vUwO8rKqY2oF4AAOf8S7Yf
VZI96Qd0ChGiE4ScBNR4q2W1brq+bA87EyehkGHYCvXTf5HTC//Bf4JayeU1mhsnimB1tmt9Pkun
UB4Ypsyu7Djy7kywb0bHX4h72UTaTGBZ+5KoD9Du7mLlvLAduse8iMR0x4aAEdvARIRhjKZ5nlO0
yA8X/fwfAPQm4cjrvwA=
`protect end_protected
