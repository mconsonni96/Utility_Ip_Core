`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
MHxtFluiZ7Ff8DkU1jmG5e4uMz7MYE5/h2kniA/K5KICNZVWFPZYlWyvt1RCszOtdGxMkPqQc09p
zw4BidK+NW4iHWtK/eYYpBY1g88F8x/k5OKJl80QgfH2Zp7J8JSHhw2E6DVwhwtNf5ujN/dvy2hd
c5y33fArwwdEuVhK7mzjWFuNa+8E65VW59RvBO1JRsXZArisCWmIEuaFTyxa3ilQ5O/RG5EYQp33
8qRNqyQxOlsEHzxJjaWI5VgqzVRxDdoDMjt8YThQOeS4T5CZftjP10GwLm3zPZ2uuLMnHIKdUZjO
mOq7/SPSwo/CVFoyiW2N/FUgAjm1qWKJWt7m1A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="W96TBbj+lkxiTXTKzl/r50zV/Nic3DsZJp8iQTRi7Po="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12800)
`protect data_block
nWDpUGWJPxjrFE1xrb+RAylVSXf0Jylj9KXuwYL/LZQlUjg4dASYpTxqtc6P/sc9iECKA33JG15j
4jYnu6u8HyexLQigwJLmm94ayaoCqC2y+vIFsOmdnV4ZmHmxYvZ6qcHGaP420y/4jhjL9thT8WD0
yafOs86i5HhcRP5TvDXBJfbmStfGYMlgUPR5KNh+PKAq76O2JRVAS9WodOQ7g+obkRdQbgdgH+0e
uX7ZBNuKXlC3AlkGoOf12bpOUA8Bq6SjkH4pLShhuMF8I0lYw6VshjzPrBR8PTqfISw4B5jedk69
jDUWgYpn0C4l9dvG57QhxnrI3h8us9Fg6y0CUVmOFu9IUCkRLpnmXNwec2a5tGZwkJlXBVBiBtVm
06f8soTfnInYtumf1FFE0eAavPC5tKht9Rw7OJk5J+ikf5ZyOn1dL+yVKgfhYve+vBzYhNBe++En
nOFYssShvb201QMu/lmrp5OOjvUPsIvQYHQsn1SnzQrYdkyt4YO9cshF/yBEvP9qvOuKEXLz94M+
3F9g+qPI6fe7Np8qCaLS3mFIb3ev9aCrnXVneL5iXXJ/i0qPVWGiwuT49Zlt3PKdajLAmvGGWLOv
TlLpd/ojiszSxSJP4dt79lZ/f+Rb7fCmdoBnJmLvWpp92CJ/We9M2PD8p7jkBQ0PO9185Ckc20mn
HNKvTsahwGgb1pfk5IYwIktXgqD8MipwfPdr2kOAvKKsoLpK9PrVnHWY7WOXOV7PygYT7dwPdjr2
vi9+zjeaE0x4xy8n970lDZjOQTkRheJ9dH0fMgSa1+yCo4Ivrm3KywUD2lChwrz264fwmXjfYlqI
3gPbbWWGqGJnOi/ZQUC66n9MO5e3JfM9xVg5YPhk2T69uNBuVWI3CB2z5TuTYXLZnyV1B4EN2wdg
tu1m+qC+QOv/7dcuzKV6Si97w0Wtw7vD9X4MrYDqr3P164TKBQF8Pr/sYDInnZgxciTsAnbArexO
KdokqiIWcSTs0/ZoZg9sS/nvncrsDfuXaOT+2ZD3JKoq5UcqPgAOhJ1Rik4nmCeCnc+67bOvqVz/
emgG+M7obfyLddXuRO+3knYjkCQDBOPm+TjFSmyAdq9OZS0jum41V8UORxH7ZU3O9oBaA0F/PmNe
jSfy0/zo5445B4uh6zao06WCSJSnAvHFX74Je6/gMMkUSlOaGwt+n3S+FWyzmd4HBB6xLGrcZzSV
JWVVq+1M3VmYcTkcPexRV0jfa7fZbiPjRy+40yqir+TpRuhaWGG1ovu9lQy/0Op5r6y39FBmkNa4
Ly720BHMpiYlCj5hTLeJHzugjORt5GbvHm1r2z5BHghP9fQZDjHSErN4gAndiHMa++f1+t79nYwk
zFRTGS6efV/9Cy0xG+VLS+u/jPNB4T8h2po+Id9b6d5jE9zYM9eYhYU66Ud9YMjt63KVO+W0IjHT
aj+lAlYPXqF7hMp8xaB3Twt28prz54nQe73MlXOlzd6Mc/TUp3FSzcV9mjdgN/GIgaHMMGzqIb+u
WLeWZfcw1ofnfq+jMpUFdFl8imfHLS43oOYVmLheyDbqGAQDlo3U3x7C/N/MnoDDAH0F19c9CL+I
4DxnM9+PFBwZFx0E4Y0B7XTOtDBrVqj9imc0LTf/43I60Y54Wh+k/2iIvfNYVKisjy5MotfX8q8y
EP2IDURQQWjhfjGPj1szE5iLRilEzCsLVXWl+yC6CA0iSAirbvvvGN0hBhnpscaLJSTjtxI/1TLX
Uy7nW6WEUI3ypjtGCNQg2ZLXkEKojuTFuLuRg4VWwkg3bpU06SlxL628ipXx8AxfjC6MQTZRY9qn
8QWGw9OgcWtTs82SbKKs0XoEsKmXz0L1isla+Ohdfycw6KFhXke4o+n+Cr9wIYVz7AJaUhb/umF2
/d/MO6cxLSdRmG9/AbS/rfK2q0mKMFUGKplSY+qMqt6KhaZxVohPubUOAD2HNCmrCcuZTthfIWmM
VcrzhGd0XTg+67el2AaHkLCoQndCiRkCJ9wy1WQdaKm4/oMk9Sf3Sinuy2OzfVCtWztsJZmtJI4A
Q6KfwY3Wge6MmSo37k7gmFAM7kBUJwC4xYXL32CCTR3M1YRjkPAFXN8WT457zSXfuwRhMXk3swaC
gNuc4ULMmxZ0fyaLz29HRfML5JkWz0AqAYfYKhsHWd/kLlf0z+nkkFaZIcwB4aOzr2vSMlXPnnYZ
Ui1jds5EFf4+6fEGn8mCut5OKXjLz0J6/R0ls5+tqLMl8n99lX8TFvGBxegNJ5whaEWz73BbcwOd
UBNXBtu+y6dTc2b2TahydE3YNoEbegGnR64BvxtaowIbXSg20NZk8epzctqz8L5s6AJwrNBj3EnP
Dh2DAfxZEm2+Ge1QV5IE4dzGbvlPkab4UtuXVdUJ4YMOTqocfMT4VwgG/7nqE3LrRNFpGE6D9Ewc
qFgtbi/2BpTNhxEqcKyLMdNHHd2mDFYoUQWZUwmYs5llyoIOxeBRNFU8gUmhSfcR3paRd20eHbZB
u5M/V+kTol9s34lqf/dfBpRqw65O27K4MpPyJ1cvFCzKzMseiyBvl6MmEt3fX5OMD2o//ydRvW3+
C3UtbaQR9Zf6ee9PjNIOWanmGXBbog1UsXl/HLVeeB0xJTZUQan/LbqG9FMHYqZlxS3i4cs+sgid
VVXp5kt6nQUpIsbA7UBrljhHndaiAUYmdc+wgQuJnpiNGNQH6cxWQtrWYdjm76kHR/87Kt3m7OQ+
Hz8td5LKcp52DVCyqzcdFvx9nN7syXgWaqrNKZVRtLVEl4VgpJ+oJpX5Nu9MKvwMvEiFwmiRNdWv
h8nL8YmeCyH+8glYuo3D45uUwcJXrHgLKACpodJfJUYlIS/YcFDx+AlsU60aTSrW2VAfXQ1gSRob
uKtMGDtjuo8sNl3lzJ1LZDWqQwhhFm/T1Fnpp4QnqrWzlb+47DFwuMsjY9MtD3BMj0KEzAsMxjCk
i12wsPh7xQbznBHKZT1/J0sEotuEmv5QbTMC+KemedtE+CMF8i5ugLQyKlBzhP0VqriYKTFT1va+
nVKxKvklw/Q1cazjyU0QjTCNs5S4IT1+2ATyLedYveG6CwMp7QyMB9bHdKTKgG2AmgD8nAUTJooG
67oboYMWXPS7zVo0dbIswjZ1+PM6z4EktU+0gnKOb+4X6QyjmrgNoy2etCO0IO85fo76t5aihusZ
CVKSEcGRsO17L1QYi745BfvGmhNzxY/wYYusdcFOiXGyI2H33mGjviflFKEbsytpPacO0R/wfVaB
44MiCxoA8b3grpyTI1TAlT1QylCyusQeCHj7a2xMjo99oms2sYaXC1SK9XLrdHuhyBOVnFpNjNrr
aL3Ksh+3lQJa7SH3O9r0iNUhX+aAlTpibrTOoUBcO3gLC25fIoCEEPTUxBcyXWnIHSy9cxCztC36
CDO+IVXqFKa8a9IjdSKf303l4Qa8+dghgkLtNsZ3I9JZXeG0sAsx3hiN0TmKLUSz+EjFpeh3E2Fn
o/WMQ1mdXwIj8/AZiLnYole0WOhU04gkQphYh9mL9z5nt9ZCTv4R6q305ViZgs7mtoTd2qxjuD3Q
lnnhbRDEVV3MDVB3Y3CAnduj3V6CdAMlKxGDb/vewbq7sr6eU5n1oemG5YuvQkA5wB+a0tRa4X+Y
krqEZOIGX45nKNwQrMrKBsVqaxHV73AxItwVl7fdh7u+vfLOet7j8zUkymjT1Hv02hUp2OozGmDZ
knN3grlO9q4gCBwFFPe+zj2VKmU0J/u2m/Oi+AZQWLY2UwwVnGSnbCx/dfcuXdFASTBKt5uXMW1J
SLhey5hjoypEqPDIxpmF1PUdnU9mEQROGM+7PXglorILBWuMnFkzORfdX9ogILOoT3CTt0z1b1T1
7BVuc2IUqipJA8+N+SFS8Pp2Xa2bEl02HJG6XRwgKTVb1/4MApU5C21JnWKkpBemk/jY8hJ23tYh
Fyr7LV1RZY3UfgNczixthD/pdgIuVSQYD+YlM/BisI0cmWno07vD8TAWU4EYuInIHNf75arEqM2O
tudBklgS13Qe2T2BQfR1sTU/ZmWrnk2ur9HBACipqtn2/0k8JtIM/j0DbAV/EUXSb1ANX4HcmxN+
XLa2PZH994DkbM5eFkxfL0543KMTW6XkjXD0n3myeLplGCdc0AKTo1JYx1TKzL+jZcXNfHhIP2cn
so9xgqSC/TCTGDi3JK/a6u+PqR237zQ3yGnkqOuOZdSlhFYNIx26nhuQRqMsFrmo/eQosXGKIeVF
c0TLYLZR7ZwP6bEzBSP3iCGSx4oBy64Bnbvolx7EOnEWA04s+xr+qZ5U9ty2LSgK1XND1BUXP37t
1/1IcpjAeBN/DvMmMN+dHTksksSVjWRur0MzNEh+E8FaT4Zv+UFUytdzE5zIwgPr5TJwXnJ0MW5Z
SX3G3b4UqyovGDdVhvNC0Rcw+P18uwJ3OvKYVn6ETOMr4OzoynurL/LoO9WVZzlolTBNcPgF0kg9
+DZMsW9szTtZFm5Rwd/r9yCu9rNxwwtNxTJjbAE+bfkF76S2cvBwC02/JueQ+th1ktjp5ap6YLUh
29C1RZVUtTHkUix3KkLyyqsIKqTYuHWQ+Mu83ozrcJ8ZlcMRdp9XB6dGHMoHlGOqG6dKN+YnJrjj
QOI01bjGAWRTkLtVMD6yqJqLaaX4CAyXZ2Vx/MwhfDLhq5b3WTnZ4eyWOuazjlZtnh1+PI/2qe44
rOqzojvafnjMVX+VfNPnDxJ0nQ5wAjiwY/PSvaV4+qJojyB9OhHBZggjeUtoPvK8tVG/o6ylxUW9
xbTvYc3ebj1NAV0d2ZlZANkPo6gTJbwbsrKaSIdwLGXAhXnYhRlFXs0f8zIewf5F+GLJ8p9E5BSG
TMAiJmiLlMbBgXIGB9OvTzB2IIKMVoXLPIboW83SsUsbDntb3ug3All3mPvEzcxPZKmOwKCw/c3h
c7B+RPpmY3GYkUeWhmAmZ7Y82CmIaFKpieXKBriQKtI47bC/oQujB77/C6xYI9C074XdWGc7H4t2
JLw+ebhPASpKJH7TPD3fakIgodQ3uSCYOtOoKem7URLSZDJqx4XBUJoicBunfugroHO44uwbupzH
bRRwO09AVi/9190qPFfWXfaKmPE/48JrxqzPyAWT5cWYxGF+serq2LZhv6P1wwzsoK9DaIDZQ99N
DWkTF5st9eu6M6SqrkxfULR4fKnjPWlGJ1mRdFR32NGChbbZds4HIyp5/pgmW7OJAr5Ix6HipiLJ
tBNBvLlKEM5IT2S9dooHngvTzTJH1LOCci/P9v5X04k7JDuz+Y5vXeM4d/B2tDN9c6trup9ahZiV
YLdapyh1U4MCAc+1HGgRI0oIj6f03jQU3pGOz1zZgPkFuZML9fhsiv34818GU+OFO96W7qgIAYA0
ENSXjYMcEyAT4BVxq/3QlHMufUS8gm6R43Jwdq3z3v4M9nImrQBqFWxTUM0cbCWp43FtuM/y9SjB
leO/qeJBGpClaf6dXzoYkTMIKjBA8AqlCg7sonmQG/X69MKMFtSKVyFoxJuLTkVnhKEgOOS2ABG9
s1wgnQLj+s2dUonEUcnY3ZzzNjl5NHXpvOWzFBPTI4mcSIo8SGFCaP1IWqVKocrX+r/AvkdjnFnl
8of7Qy5Qg2YgK0LyoXknOIP2+rsiR4i7Rm3gjibSGal89xWR1x8Et0r1H6O8JC5LD9qpb+pwgd4v
g6dkaEG/rrMviEO5TsX2FsjwPqI5QKk9iWPcC194Bcn3x6qNFW/sIAnBgl1/oUvbg8FP3Gzi3tuR
9K+tVJaXAPU9bJg4wGBqJda2D79iSgfrIrS2oRX3U1Tse1AVaBIOdpI4aLAEBGdfMOOB7pA/thSv
DkxYs+Dg109eChiTSjFj5mVKDjsv0hSPsOZvvuNticHM4iJmkOl5D/jJsvAPeVvTUEmEi1ptSzPT
qz2E99/0Zrn/GOa4jNR0Kuhf+ZjsQXAyOVnLd7yX6mlkToLMbaES6s36aC2sWU4gBcldEOc2x9/y
gjC8gtYYz+21Hlkf6B3Mja+bXip1fAmXZwcqE3MV4s7mLuzd/R878Cil7zLcAX7OY52K8cg4UrMH
smM+hfFICewZzLoFn8KP9U19W+0rhu9T0cQFg339rnRhmC4Z/5SNVjCVkMK/dKHPUK3eiy+dZKdF
p0gwqCE4gKYR36kBqa63rvooI7QSeD1K6wXHrOG04Xh1mzXYVxc7JSmnqK/KXXto4gAvjTMgzhvL
+Drwxf76eDCY1ewBa13z0zrJVJrZV3PronGvNqOOnKG1WLRtb/L4ETTVXMctOADw8vpSkz3r9k6W
ujs1uX3s1TLBzxtCz6qaz/PgXMRdJkqebgcQvRJeKFeRl9clVDzwemCEHyMMzsW9FCfg/05PLw8q
ctdvNI8kfzmMrm18icMNfNujuYFd5FXQJUA5y393UZcDZNXojMM8V57kn2S2akAa1cVy95TmDI1G
osLoHus+ZA3iGTREl0yr3LcJt3Z088PIX39w2IPHQ6/KvkB2W7s4X3l36Hzo/YfVMekLCYX/KHzs
txxFR0tb8GeoTXRbX9uUTPSULtXuYIMLRzyLsE+g0jaVyKxnDFjEuNak1gsoLP97k70FnZO/JG9P
5tz+ojI+buxuwpX5Wd+WHMgHGcRD+weMAWFt3do1FSWApkSelCwjLkkj2tAwCo0Kx3AtV+ZNw9CK
Oen+0VhXl2DpOUx07P+YgolfrNKa3wjq8iF5hddVv8RChlNAGQwEysdQH/TFPvvy3uPjKkQEhevf
CUq7aPs0BTMcwslT12FP4KaizAGayaPJNhEkhoOD3uS8HNFq5FD8jTdt7WERWr8Ib0DD7/hvNL0W
VI6MiTZK4/qYtaBoDDsq7ahPbGQu9diZ3A2ehka5ptbS7ffvv0VwL2ASdMT/3cT43xd6mfbVpUZu
v9Eqr+FxlAbnsUMy5VJvtI4+qbVrcqmOfntn4k1AgNF2bFCX/AstnlAG0+l6RuwPfwRr4cmqvEjx
voQLlNzUVDCHnN7R+dYodcg3jhotRGB1J2MpNJIn7nkzhhP37+YBxQKjhLMtRiFzjAvW6vn3OjbB
anY6cKaFZeanRJOoxK2lg+/9bJYcVWthpPKzWn43lrnKvEYFhzHvnXBTntlBCToChgpW+F9DTZYY
fvA6EdkqHhToAoHQYxT4nwtHR4SCL0N44Gas3W7Omii4qVDeHkbkXMgq+TCbKCxutJ1pnQiVcD/1
7F67CUG2LLEwhWcZipg4olKQhUF8MUdWZ4nOareocb7uQGqn2g4e18NPKU3m9RXB1RkL62Naoybr
giDOquYGX6DcwmJge1scfqiwZ28tQ+TDmI1RbqFMzDYy7M8NohpbVv8oeyLZ3hYR0LKQNg6dWTuY
eU734bGnJdPjRgoPapoFL733sFfcda7OL93xSUCpLOZN9pO43towdTV6Pg+m9Vl8It6EoWHMou4Z
a0lAbH+S0O59eShi70G1d5IwqWUpVMQDTF8L+WlTN+SVjSYZtuksmBDxo7RpEeFiKbOxck2bjmZH
WODRyh/hlVc3rbgP+8EGeSt8DbXQVGH2rnw1jgtl3UdObMq1+2eTY0AxhREGnf5W9jqiAYCxlTr8
rFbQxydHPdeGuSNyHgBK9l7PUP8jIddpor6cJtSb8t8RqynxrUM+42QaWuOJ1DFjjyHMBPZk5evR
qj9F915hLXXsHgU6/6W94qWPJA+jHC5zGErpUE9KDAq68xAfyWj8Ro6yPxg4UbIKwsR6zVDzSZdj
BqaOvFE+5i0/BjwBc4KWhB/LxbBbvBuFNbQcyFt/lCHuYx6vL4yioCpxXZnc93LLntbHL39sikFs
k0xu5fcR5+aHRY7yPrhtviZUdLsd3kTJGkSnHloXbd4SqgigEaD+TUfA5lgsgfnolxwF398iE4bW
3GKgVR43kfUxbg7DWnYBmZ33Tp1RSxK2rxLWdmn4bCA3M70U0Yh/eu5GW7tPRzoCtR3cmzf9k3vC
eh4WFyd5FnCBItifngFWSjWys+h6PXj2GtsDLPchsdVhChYE/TZ2zpOT7lNisFC6/rb+bBic+Zv4
7zsL8KF5fCTVJwoBBvI4uj9FdskDswkUrDxbzGWx6dGiTaIMyJcKAF6wDXP2bQjEvL7aTwGMgmQr
u5Xm/0zmzESnlvPxrBLZ4lbTpwowxvZcGoXqZ4Zrgz6hcg7ZiUSYnobIB9nW2AwZV6yoOAPtyNK/
LDh7hMz2QLbAc/uCbY24QTpTQvJhSzkgOwWYxionF7iDTh5WOmlCtaXXrK+GHTUbaX1/26/Nt2d2
3b4aKIWTGpR46hDzpFAvdi0eiUH6iMaFuu0p14e0K/YyEQ9RP/bo46nbYjUOCrJVxUSQ841ub1do
j/qIkln+IYM6spo8AKdx9FJricK/DNisvkVwUnaZ+XcoxVSU81fCfMGOa7uIAg60K2Kqmxje1l7S
Z/Hx/zgyT6TIqHD4UgsWYUVpGxVYCynJ+trFiWKLYQnib0yMVS6/u07Op4jWWhTl0ovETbzSDo+f
htc8UOoDweZuZWE1YTzA9IwJFef3SreMeL53IIwANvSgWW54p6Db3NK0Xz6gnv8SMnQn6LRRykS5
hRocOxno7LOsFArZlr+5YrkrEAwz5ITk/nKNFLXC+SUBZd9gpRfqUjsoNA1QU2QJcrxOaN1afdih
6e2CbasxbW4MCN4pL03EsBM1eTyYyjN+OLgUpe82/zgIW1icimGee0nDppcPYV/yWbVzAimljOhl
f2/tOXKRiuyd7dRDDgSq/VDKUTrMZ+gR/ehSLcXM8iooiso8dfJI0OWXHyqojplvVcJXafVMFjQn
jWnfxFBtqXjPrS+mug4TDjO+8jgjXYOShV5AunSgfgJLMY/GJzb6TcrxJSCzOz19vKQvDatM8D4C
ijxhoiz5ptcXJqP+qyV5/7TKpZnXCg4gJPgeXrex8kR+AF+BPbxsO8LAqTpwYYZN0pjwHi94fa8A
UuuQ1MsrbRPfs2S1Pc+Khp42sDS18GMJpnhtQd0xIsqBZunQRb9CImorznAdUBPC/3NKCo6kJ+Y6
6cWMycASd8bnuYclY57AfalKpi+cE5QCGyddZwisjJK1RGU7v8eyYfMQE3HWMEJcAnWeu7bxusdE
Fnr0hzoTqMO6nuTAGzpHF2sIaBydnn19q++x553cdtjE0B3fAs7fT0dFbRHs92hpwmuCVenQK06X
9FCHQTey2BbHZ1BbxCm2FweqSBtZYL11At+jMm9qdDqr+qpUxBhCkACMTK5wyTRfJ4x0hT2fIoTR
ThPiBv0ZVfjeVBDsbJ8/U0lSmdbcm8BU0aoiIrGa7Sopopd0jHxjYIjWnNxxG3TQhokiDN1VXp9P
vFFfAfgCkzRWx4VBOmvbA+ZqDfoGsCU6gmrEKZcp23e7a4G/oLuqAUewrc+w6+88DOYFOV3jLL3Z
gh7qHZEqSxGGQhzH/l6F1TiKNy1KxeH0ZKv+8mvSnI23ZCQuA31XmZiTCdYtZlMVbSshnfpHinw4
r9YK6OAyTiehN0QqmQ3u/y1P41zIfugCnxCOErJqr0H2zwvIhy87whFHggOpvC8IF050WAAQXXlz
H4yHjSw4PD5Br1Pmp2QwocsGwIak8ymGFroVU0Oi+aRhm9ZbNde2RQC21yHNDucj8jozvx+94xOu
giueVZu3IipSylMnpL7Ludt43lu8g3GycUqyRqg6RFftGbRrbzO7QbuRpo2iFJDjNpn5ak3lfaDN
QomcVXdVzyScY/EpHNQjtu7zYijUeyOYkZiS2DGlny2KrVLn3WGFkM/vilYej53bw0GvIjNHTkrc
L8mpzx4DUTgz1aRylovznSDXJ18Jo7YPP4kYnBXFLGyEfsbHnBZPXo3gCVkU/4weHvDNX6rNzP5V
n4LVXPFuL++aswYb4/A/Nsm+Tg0alV/4a1aqvOlJYo+v1AmQEnT/hQTd4J44ma3TH1ni0s9vOphO
YQE8O1852ZN2Kd6LqVXDumbQYFP//eStBe51+W2+ySa3Jn5ydhX90MOnJota0fN0esOo06z8Lj/h
cvEIvGDM3F9ixU5u/o/i6uYaWHmE7Bluh/lp0Zxs2/X41S93XxFCW2Owo2KdZXsciXD3pXoxwS/c
FHLmA6G0im2xfw6R9lOCSGmmuWxEvT6mw1kGVOkrB5VtQaP927nwYbwvg8FO2Xeq9xLQZbp4/OSo
vBjy+prYr1rDciS7tdbtnH0J6NWV84UCxuol9RTRhkwiaeTHq+yl+icU6ET6RaCBo78O9/ABwXle
wEEF1FTHfrNzgYxQn3kVQl+T8WFWo9vzNLLbNdX2/m+l3ic1gh3ZYW7h0J674OrhKt4prgxdZm3d
f43WX3j+GJgHSqkN9tEulbHSs+KkEwXkzJJYnfNbDKQtWscg4ICDR1+PW3qQYFmjMSSUflvLVDph
EYRF60Un5vOzB6b7U96mzSCCYLOOfhj7ZhD6fSv0EUyBIoX8HsQIAAHvMKOTvk2qhl0DCDzR2qr4
OVN31wU6SCzna2kOWM5cYV8Coq+I90jXaoaBZyB4zEdYC38xUjBohX8B58fcseqGda5x5HtS7iVv
l2ooMWSEVTS9andYa/aIunaUbmFSEKOBlCc40I+yR4yma9NrOmFG1X8tCqTDEOLsE1Y3D8n+8Yx1
kF85Gh0ryylXLuouzTOE609SPuBNPhv7YwuvMBn+svqBKKdC0NSHrMWfwFnd6GfCLAb3Tb4XqyUF
O3hX3kSHj0rcvo4Nw7CymTBKwN3pY2VS4KCzY9XXCb3v4N0rmQJKeVT980lTI9255ZbpEagcBQeH
tD78qxLa2NVHV6sg/qepRm+8WbeZI+pP+zub/vBqs2aKhKSb7MXiN+N2E9nOAGQni8R2Ry1T9sSG
Asqp5uNdmoyqI1tQcX9vVB2dKRfz9GJEtUU1tEmsRLjycY7soSV0/lWyNc1zlDy0h0SQkT17zEj5
Ef1nTQRomLU5DFUI8n7K+XT2sZ0ixS4v6MPRql6Qo/daFcVp6ypZQ8CoPc9ZRQEqGb3p0Hq3S3w2
9X84aDTKTzfHcnum1K5nOVnfSyOtXupnrqRJO+1KeSdX3s/hTpvcvfPppI6kVyyXQ389fvqWhfiZ
FpX/mvX0GCUWPo3WSIzjqsgwBqVOiDTNAbYAM1c60tLkxN/Yxmx+NGDjfK5jmbkIzVwl4M+zfrgr
HzTJ9d/GwUby5R+AfSLCY5elx8+dH8RNBI8f+D39Jr9ZladTkBkQdsSmwxbakUZdwNU4xmGtcQuK
xI+Murq6icnreNmRmiCUFNc9IAtXtnqEWFZglK0JH+cQpueiwwin6+kSzldkY5SEjhl+gSgn/6zC
809JyO8aL/RUkpA6gTwrSm39qu9zZPMUGV2vdHg+6MkHIJZSD0/3ySiA39CiHV1AQ5MbsXnVC/pi
C++vdD7v4xDJM1mHW7GMhJULPCmuhcC119VByNCWijBwQkZk2o7F7eKWfxUSmXNAcK+Pd9FyF6ax
Xc1jt7G8sVtFz+/1PW8fRy5EZ6onf46TKe24zOQ1bgOdzK9rzZoJKkG21TddsOLnEndrPeCcDrdE
wOW5qEWDxWYJvy3qfO4b+/AJNPP6YTcVzSevyNiUEpZ7gX/zP25uwBiA/wF7P6oj1CyXmioShmGf
oMS97fvpHZ5jO3UQZ8dDbZzjx1TlVXK27cyIlud+eSstqe6cJjFpfBPeCrs3OWJsHH7kI69vaSWs
ADG9nALYd1mDJFirEgRySzlOWHoVgm9lqbBlx8zTaAtdz9GCY64v4pcVqn+SFygrguv42lcSEa1x
IeCykXwdd/2k303YU5prTYXjSjIt0Asfi7ODd/85E233Kshau9N3vjuoCWi0Mr/rPP9gPmcCoef1
YrWGHhB8VcD2ah548G6b7ASJb3i8JLSii9Zwp3asfe94HnJm6CGFe/Kj4hMAKp24eavy/h1YgpIv
YIAtGIkdiWilnxHHmeM/rhwIlgdJuSq/1C/iAxxZw8Q/bNy9rmqObI0F7oO0+Qg+tN+bBVUSVE8Q
4WEoXHb5PKBMb3ETzG9BhuEAABmV6rq3uVv+TN+pZ4KEOaJwJRf7Ng4Slwl6aLpwMguWl7lpLOST
tbBoUxzFG1id3NE1d0J6abSL28apq0kBCUX1Vd1hzyLD+azBXzoMfB6JAFhHkVn9BYzvMHM70rJ1
k3S2/VQYhPFnvZx+8ytWTVfhCWzq4hjdqk4VUzIdRIe96gfnHDLaGK8TXokkyFZkRI14p2J90Tni
nBy2SXEbBUCmedBIa6a4otuwgFWJg8cMq4Ohs0yoBIWWdggGqaeEbnqLIcvhk6dEAaia/ZzK1WJM
3dTnT3ZF9NVJVoywgYdHTmYszvWs9JaETKtiPnUKjJlwjYH7o09QlRsvjPqEYr2kQFruP5XpIo4s
SnhFqueBsCAWdLxUDYWyvxiTcMZY2rAc6CFDRJK+TPXnSVwiNkMn/Sj1CAVwqeiG9pmgbJ9ezhrq
ABEzXHGnlerB+UBYNHA1kxdMbgnxvH5PsueEn0/+6LAhT84F+vACshM28+6z057v0bSy9r/Med+w
AJT7zhLKWuewaI38JRMDFoKTzIByyHJxktrXfkBsbZjoWPAdaNgLrkqdR5frKaUIOWS3/9FaXX9E
BJOEoao0KG8So4cAgl5vlvZvqV5ZUJHT4wbKnMP2k2D9i8g8hBDlf3Je+SQLMYQ1KErewIQJ9r9M
e/0UNZKX4MmcwphaBrWmOCq4m+dxoGvNCGn2Nsv6PJWClVgjTJGHHifaKINwqaO3xBYb4JG19SXs
kM+3U5tx3DSbzmLYlsSSU0fx7JCeqV4Ke10ZYq8ELP9hOAT8nAMGWD2SvKAcDXLGZUDgXzKaO3ci
n++MVbIQTFpe1rq0P8XNZIonMaupg/ULF7onrBeM46YWLFkeoZ60NXPabiFLSKIKa0FuNHXEKT0n
J0tehwdzduwuPPmRsMIudGp6rARgb9tzQt3Ns2JMLZpCrSFkRGi7odwWd5+06m3HzAWS3NWPSpRt
bmQjq8cNCaqsoW2FsBQPEZK+E2RyncvAnZJFqJx3WIumXNAl/9nHc1QzueMQR7PPokAE8Vy+VYeM
7k2rl7zX7KKb3qQmLIAWe8+FJbD7SpFSoTg71MhbS7ImSZ0+bEPQTIenwCUVmooJ59hXQ8wWqOI8
dbdURjbnpt3wS7hUvp/3dxSiCK1FZsmD03tzpM3iedpJAwPZRrsNfUn9IXIgM13NjXWFFNkdxxk6
nn2QifG8U3om/4ZJX2u8dsGkh/AvygWzOchcLCrhJwHoBG6FEYOvibd+tjeKtzw+Ust4JiiUiOvq
FmM1DoXXl3VJKq49Kye+58Tit8SGpHSZzyz9mNLDnz6WKqgbetCmoQh8dv97r6TmAcLLXWnvQqO5
upMEbR/sGripo3i9fBvN2hJLz3Ln0TQoo/u5TGl4PdTuXK5kIWOssHfnnvRP7oHaYL2XTOycqT1S
cxY5oOxILfv7jau1cz3QGrPrlHR+v2X0HNfwNE0UzSU8RwhttwSpXftKKNWCGO1bBW2upG4ssS9k
rIFB2ARcmbC4kS65u6WU7YejesPFaLMcFlM+qIroZfboWueQDEqHyQt639RQobEjTalEaBfnq+PO
LH2LHuxX0mvG5xRa9UzMcduriVcF47rUnBnL4Zo24LE+3QYkMzWcNGmhsQQBzN4d2yJhWhZqLl2b
orzNnff4PixtvRrFzJPdEQNzrikWa5yVsthK8LtCjqBHvWxRqtB+j+98EVHSlrv3FV1hGLNuH8ml
1kZaabGVjXsc2g+4EPxcFtHxCTPchB2F32NdT5gdV2GigdogclhwI0O2RoSz5HQ/ALlKFl7f1Guj
JCn/HJ2SMDH/goctmaIgJMh9JgB4GGImqBV7lozOAPE3AHGjKPAYa8ST9nLT5QCNmQ0J7MyVEGeN
YYfkxA5GdqOhozRXtK9lBjJyNj5ZSAu/GmOdDbq6zxqkHyKiT8kOQQAtlIwsDYd/iy8vFhRy3X7B
rYO0ajMK4Pt8PggnSDkjrOGgDToxrAiu0Xyd7N3X5bmhAMm9/EIkSqJqJHcDfj1ONrCRKFa346ib
iSZXgNmzHlFvLxo8voLHBaXrEbmVEiBeMkwx9OA9i7B54rqotQr26a08hrtUrCv5DUweB6CRvIky
wsh9t8G80fUzIZ6Z2lJgQ49xEnajavyu9WNg6upwYSDX8p+gbp0h9h9Jbk60ls0HHXC6bFri6SCk
9GMa9IUOtfS/xnnFnJTaFFNlcdzL2deqH1ygEDBqiF36q1+ndQoQqiyv4d4dgL6WhL+GwxnWkX/b
SBXjKwi6Jf/SLxCKl7NZ1NoO1/QM6cd5h8fm+5qwiWH757sTzYOGihwaADMcOKI8K5PERJXRXAFq
HJU44x0M+Zbo+cYy3WhT4LKkUtEGaK9gtID2RWQW+4iS0o7mYQouWtotxmzoEaXgmwDAfcsbiDXb
b/Ph01jI1L5PfIw2FjNktyFSuHXXCLLhQw6MB7vwL+FWaTPty8WZmsxSC57maCBVajyp7kVDx6jq
l+JhcSoZSiqC9RCrp5c5sh3OO3cH9QPSXrboyc3FqyGZOw2sBVq+0jrlU1ODdewMdyoePIpMAF4g
6a1JKKUs210rjC9nXV1Z08UpFl+rspCFo7y45uqzHwDPkb4GmpKqRoqd5feobo/H/DbZFSiZtlg9
0hPScl5Zbtg0+k8D+gqDTIsu/YI804r51vOmHTtxGoqEZkS3GUZwwOkRGsOUAiJFrPiuaC4my8JR
hhKRPwpc+xKYG0WPvIMPbeoJIswS/544+VhBwXdzciVWG1xs8zAzk751Sravoc/8KooMspCE0k8d
80gKlzIhWM6OZleYezeDDM+ouP0MQ/NGfAFPaAPWOMWVR70Kj5Jv0GUVp08YfQe4aKkp9ff15IJ7
OxwhYROXc8Wqx384B8KxU8Ira+nn1AnbYULvYxIGFD/SY8JMqNDOse8qViGmYzwBRzSP2kw/RSI2
DoULBh7zaZPtyl4R4EKSa+do/Ir9j1zqgkwEiL4ymtIb9FCS1c2XavpDkl8mzXUSSbn/Mbk4EqQ3
gfFlV7dPZyxQ9eRdCcaZhM9PR6kwjtaA57hZgskiZZPq7qUUA4RWm+pgRHJDdB67NGFMpBme9mTw
Ffo0l69VyqVUjBUnEU/eKxY1jy2S5zElOq92IEnf6zaXsDulq+fGq9RIGt/XiKAw5E3YvkA7FHS8
XRV7KzXfk7M6N8ySfYDZNuXSBGaRjzkatW+Z8MwTN2aUb/goLzjIOEY0MI/1Q72MiPtTwIVZJ1Gb
PoEJcN0Zvmqb6FaJYRo1Z7v8fWwBsMhn8LxLDK0z/9GKS2eabaNKnlCPZ4k4wPJrIZAq6bPmscL5
u81FJMUclrD7stGegCHsGtUkSKkP3evlZtRchZ2ecRXyvqS194KeHcRa+w3P6kXc7lMegu2Lsjzl
KOs9EAKpYq1j7PXPDplsk+wHgL5MOceWOH7YAGYeFeXugy06J0umSEgS+vwssf7zmkA6P6mT8rIB
f1T3/UJlN67nEe3ZkpP2/AjHiJjLMtfdkRiZURNM6eoblJi7NOG99LGWLuNTwpPkgG6HtUUVGVHG
QK1rkRHYGBkEOpNrzf5Y1XLWIC5AoGll3tAa0HDbMM4Dkp02vVCfCty1yTsAK45Xqgrkiz6sfZjX
Xc7jBcgNwHpF/TjdlcVD11gLIS7n+fKF95ayRYZij0Is9rRFCs5JImMsUDD8+WsqbAdhD2BWrIPb
oHdhJOZ/GLroOZKB78JfZO2igIt2D1mRP2BV6GqrW0qOHJ5SXXcI6QP0IQXjBQ050VFZ7CE2X85R
nvMcPoZBOrgVdzXHqczOaZ1lt99dwtYhRa5rfZRJCwvUkLjypEffBNrZhBikh1r1uHl+L4Rmk9Tl
HOlGZpDBmxFsieWSR3JJIuHZxhjsYQi1krGAKlXl/ZH1bHZpME3oXNXG9x3fo7MoeRcTPi7y3saS
0Z1TLCMAQ7TC7cywSBJdC1yslFgi2fxxZaNR0ZWtjVqJ0VyoFdZEc3XNotgknIab7ZQ/SqAlCney
c9Ys97ydVoiY6miBXKGszbsLQUFrm+D/PvCX2Yc0fqOoKgqmmG54vT5v5XJul15VmRWjvQ5sr/l8
uIDhm7vH/6K8ILcV/0o6RXFoIjdNyVEya0+OKWbvkEJfX7FJfRtq2g3LEAkvd1gjGbMEq9W1Np6M
fML56WypdNqxGmfr+uLLq9nGvgp1RNDu8lWSxycUqneGhH2tn7BFkjz6STRIz2oqW3vMJKzk8pMm
B6srUd+ZD8Y/Jn6Dj/FyZzHJtl0kvuxfNMrRai+BurNqHHwetINC0hriZjVXf9+em7oKoMr1iDMQ
CCEl0rwJXa2ZKHbUieozpLCFXTlI8Huo3R+AR5cCQMG9JIZe9o+yswKaJa0GcM54WNlV/i5ETTEz
LPz4zfUhSlbU+WH93dLU3SlR+/uLj0GsTfnMaiAxE8E6nBfe4DccsWc6SMdNuJgKaEw08xZ067nc
GvEngDNXEUg1EoqLo/roaDIJ2AajpofoiNS2IEodcfRhqlfbXgnWJkzQKMkt4B01+loJmLBxKcBA
E1ytD9/19smGZymoTnyH6t+/6QtA51qpU7sudQb+57lHKOf/svP+HjcU87rAOJ5W1E3nzxYUUlds
hl+3XBOl/kSAbm5kxMCmWm4WDqwCPx+TongtZc+nzjY8LBQ2ZxCgZST6dRCuQT+hnOuGCJOc2QjP
Eu5O1f1V8fm1IDURdzzowufy+pyckCxvuTP2ULcJ8EUiinAjrkY7GBJh4YnsdUdvaSqf90EfxTTY
dlb2StrBRsvWoSICMOxoROmfhQhy7qFLtNRr8eipy0X1feUDNq11JzSLvBhus8BaPgjgVlJCt1ov
Zl6xmiHooVunIOO0JCNQ2y8WMaed55VLq/b1OfA3o4ApOK3x4V8PUWNG6jkYFFeBh5X6q3L5HIjb
ZgRuJ8ESyjUwmc/rVrZkcX/rSVzM7wjK4zc5sWwg9Y+vW5bT7PNExqARdXIKgWCBcgFom0Lb+e8L
4qx3svFpJkPW3enskostajW3tVJpTwnCmA4w4OZXkMM=
`protect end_protected
