`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
h7HqNKiqIEeXB5Xm2+jjy8Ol60BZlTMpaKcrYQxuaPMjAWTtXnDjR5YBxLDcwSUpbu4Iw1Y5ZZa5
NgVS+FhvfqrpD4S1L6xF3qRXhNDJGh77N9xLA+tjR/SKnHtbQZR6MNSDS3d8sk24ZGJX+XWid8zT
iTdq+Il0X+Di6gZ7M9VrEeEMnyVnCkTfsVDmgMU0nxC3rE2rRDrW3VQW0odHuGdDdvU2HM6jHVUS
TbolCwzA6O0Fq7eApq3w+vVr4OMxL8+Fz9TLRap4zzIUkYacNm6jR3/KOA6oM+xT+n3ZdHx2X+q8
HHxTRznVQqmWh/42gUdJFvTyxxPPaNePqiebxw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Qg3fSG3CNEBzjVmkFfiWYWtShaNq7pfLY0QRvq1XnbA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 139808)
`protect data_block
9TSGhGDVo6dTPM9ec6hDgqJGRySfsZtH7x1WRFIsPc4aDPTA0schk+3xmoNl9Ic3/NuSSAQQSxbn
k7QeV21ft4FzPW8UboZqFJYBoFYXipgszFKtVSCotDj5mUIihBz6hz2Evp7e7kc33qyJ6LT+sn/3
VZzG94jwzzzVROUxVKlZBmvSZBwPQZPNqAykaq2xudpetwCaawfz9+7P4ygUJUnslGnjhkKXfsCa
ecW4Is16BlDCwsjI5JxYNfVq98SywWY59TBsC53QiiRcP0XCSrPr7uWi3dnmACBUAnX/sIVakuyQ
BJTp3W0kfvmff3vo0+UW9euueTIl/0nLRd09f3JOunBHeTNMfeDhSC7cSLqdSw0T/r6zGyXwyZ2z
NwDmHfZsLoEhtR2SmZeYW813oVSVb/DCF2+LAAtM/OOOV8dDr7z+rBZ3xM5lXcX1zfLsUv6lOtjr
CqLw9RPU835xrrvKhPPHC46EOduZPsclUcAn5dELvW9eY1mR+bFelwno0vbWLaP0KoF1e4Kl34q4
y8EwgZKk0qx9eZEKqtIWEPz6PtiPwaNF63caj9LDttBNazWzqCW5dxiMHQeJciIqwSTmPRv38K52
bIgxnwhVk3W52kpENf7dKr+sIqPxtqewSMMxIxfwH31r5DFH1ZKzGqtPmLjU4yVpNrn6voFXPhgj
RpCqR+6D4EU7hKR4JTrsv6QHUxbWpAMAClnp3LfYn/QwIuxdFKOmK1KhZVejlOmnAHuoWM8heOKZ
8iT6mFofLeYmVfX5A74ufBHEJorwbkfJ0xwgaN0AptU4oCjT/49I7wvdeUuEGviH3WtOsORbjqiq
hCOtmr3gwZ2cro8Ez7ErRl4BSyvNGwV2JcMoCRs26p+EALqe7lo9OqbphtjjVU60Uhx99I9xedm/
KThsd751qoD4hF7MEX1KtsZC5uL7ST4Df2S0g8w5TwVzd57OXf12h9tbw7pVgjcTpr8HxTLymOUY
CwJZws4nIrAmTFsRSno84nWsmEzz1ZGyD2wcjQIBA8d1UU3VznZQccSz5CdNljIQtatinL+I5s0G
oFyX21V5ZTXsRJtwvIUOlsEA6eNiZfqrm3cykbzE6nRGmINRozB3GX9XkVUPYZ1eJSxeXQH3dAmu
AsYKzw0nXPAC04CAKwRrOmy3E9WL+rQ/mhHiQxgDuKNQZa450BNFLHmS5BDK7JPwzbaZumYy0UKc
UQkU7uuJfvo2ZDYINjeOqL4X6pVCD6kGVNf27mRA2MtMX8U3doPXfJxfL/fLG87rh5DdOWwi8eyr
b5AO9IFsFc7WJ/rNkFGSAzbKohwWeISorOQwGcsDwzzMJuzGfP4AmPcWl1Kg+0vbNfmbXi3cDRPl
Fp5ie9dhnwFzC8okji5KyYIB0ny+gzdtke5r2B3/+aYybXLRjKPjqRL+Ey01NPo25jYnySOKM8vv
FTc8c3uyIlhDbBtQ0PgHHmhajUTFA+bNyL24b16BSmRdwK8HA4H5FVFjD5fvaZCx3fJHBuEMtgJE
vaO7lSLtLYjS94dhygl24WXNhJWN0EDKDHbCVw2XcCpsEkQc9/syYkLT4MNoFVL4YXR/jOxQDOz8
GZKPxnvgsDsmOaY89LKfVebtzkqDDNuk+3c95EDeseeE5BJ6z2b6TExpGRUAzlANpegf2o0gE5In
zlGcce/6NDGh7xHKbJY1g/A/umI3sy5INTiazexVKeY1aEjVueBvg+ZnLWPd2FjDyXZaCxAjclE+
beTV5lp+jspEGnI8+iJxDcd0I+Lsm1RKvdKVCuNYSuQHtGTu7Dn2IEJt6AcEy9HN8PFm5hNuBFSW
hQCpprmvi1zOxPK+0hAxGrbP39+BaskO1JmPuC+mzuf4Pc/03uTadqQFMNScnq5M6fPey6KTWN5l
7WlBKkQ6RwIZIGi3ns41vQ7FiH+iz6t2rusL2aPJ/mPg0/oBN1wMBIaX2z/XC3u9x4sVjjwVEr8x
EqNi3ix1SAZMbQp8Zd3c0eFKxgg1bump+Tb0BT8WObJ/FCbt9K1KIXkHnar4c/POLEgxe00ctIW7
gNOgx6cpvn9jE9OwRUVUH0Hf92/oriPstmSb3xvR9BL6LBnY4vTFGx77bZ0VoDXGIgHpDZ/BZn1R
rhFev7jFOVsgjTeg7lVJXBDOdEtvj4tNKQrRPa41tQTLguIvkzlz6SZqUxq/61kn0bNj3Jx00AMh
t1e7/+FRtANuAZrg5JVSE1K4/Mupi1I/JTl+ZS6VZT6JOmXcLowX00Wmxm/Tpls9rRyzi17AHaDp
takiCVDGssddb5YWubeX5rCE9DoZx/vfaUTXAzDaPIoLosYfKfg7X5rel1EItm9p1DMdEJHmyQop
rjHw4+YewABOCnqglQjE7qG1Ac0h8uCF+N1st8B5Qn+U1Aww//p2iFDncPi4kLA93eKhlY/f0ASn
Owhlilul8MToyFnyEhE4L5DX35jeKH2YrcG4ygi0B6WNUWjyLwAcyPoU1/Dn+SBduxjtwbg3Wiwo
UX8c76qJdxOy0ocQFyqTwuK/IHZuF0xd5xB7X8mvBWmPx9f9NuqXT3fOXrpplxdZpYv+9ErH1fcc
OYbT6Ro4/fNpyPqxYxlgf2/aFEyFK1AdB+QxHtk9ITG0bOEC5Rug2r5fwrE7mTxygkxe+uNEeSgo
QEik/HZupM16focEYUT0t1zLAOCVXcVyoOrNw2KnQAwBULXyxxhlG6twvxfd86NuuzsVzQ5H5kSD
sZu7BFnzWy5EgdgTVfYu4yDScpZu7ZH+sf4KfWHSArD++ExA3LV+zKur0YXzXG/j7OwzED9Jt/xZ
pfaKERlg7tLfxDFAHZ2pCqypExCH8nCj5sayDIt1puFCgHWsSoob7UB8+iKbUb+NxwcLzOGTKIMI
ErkwMlV0MUaBRQGJhOvesVGhPDokNQPPhs1gD/IBmlVBkbCAYAaBog0Hu/oJwU9juROa0+DDDJsl
J3pxigClmBofbiz4xzIyS4m/YbqbLpLhUesVJQJyYIPXJANsJLX7Gt8BofYP5z2gOAtHBQamXp9k
qvx9RhsIuTxmApvX8QXtNFj99zXTIrbRAhyXjUlsiX8RqYPaACiH8iB8xWUAMY1tmnXj3o+4HzMj
tGn6AeGvLmLydvDkRctDVuv98ejqP9dcoSIGQ6oOgNQ1krJHQEN3NTVf02+F4YRUx3gC7gdyalZP
dxcP8u3jbhr2/RUxtmNVYlfnC8EdO0E1UZ9kHWpRTGNeCBL7oKSTdt3i5Cy6dl2Pfei8cfa1y84c
gb880MSuodkSobSYAjD5mKFB59FKPwwfMjV5483HhZA8+DsmtTMSTaWsPS2teV6gXU50pxyK9Qq5
9NeYhYUiUtgEL+PcyCjRSDZL3y0RNPwU6eT0YmFh85qM1WNlsggGM8fvR8z33GP0mmumG7LDqUwC
ZdJ5MI+CouY5zIT4gJxx7qWCm1ZEXXYH3FcJiK49l8YRo6SuNo0qVQ+NkHmBoZKB47WrEJz+0nDu
ygXhor9D92dCPAs9ixrcIy0OIDqzXUSYKbRjPXNQhe1RpO8hOrvVOvy6bAegYh18u3dFrrmqokD0
s2nWBJNwM/kzZyo9QgefiUUmH0ucnzBE4F2hbDKI7iec2ZmfJ33O3c60RQujRYsNxonDw6zjq85q
9VYg3as5aqzMmIwBbivZA1/VJiglYBsodMPbzlU3CFQ44yrb1186Q/qZSmjnJideXEx1vGOaEKuJ
58CRHDQtB6c5vyUiT0wmuGf3hx4Sw9C1nXS2rAtsWo4TaqboWCxlSTKYKAP0fDqhyxlHzTq4mHwh
SSgH9n+xD/QGxk4IzmfzNU/tIVOzanqpDUyS8COyFp3LQy7cg9zlpNjo1YbIA6t2KAMyd6TXcZgJ
t3kpLYkcBrIfuQTQdyCWGvbd0bCkESjClotCgASv5rCC4yEN3kKLRWSPGjQ9vndurBXeOku6woON
SkD5OGnUucKS7aca1IfSkqfIfR1JBDhVKgKWVd20bruz/bFM+L9VTjbk4oBiR6MCAh11aHtUjXMK
sa0lyInZ+0lH1/3sYmtiKAyxr0roLzhZPVyk4DTJtCl9y5GOSINh0+J4XzP2ajm0jjPKjBGDmc9C
Q75ClXG2ZhqIAIReNngLNFoxCT7RV7ljPjvjFKPj25tMHupTKbkJ97YW8A78ppEa+xTh7n0jOByo
Pj7RE7CuMCvUfvAOnayhAYk3bfqDb62cKT++JBXMyDJgOr8KJjUWS9CwPyupzTB0NMwgV64bM+Is
lhGouyHtpsAHhqa/JZfrftMfDQ/VLJypdC6FJQKYyLbs3kLy2HJnJrnLXkwTI4qiAPVUBbzD+2YG
aG0w/6Hc3R2vm5AXHQMG3Cy0u8zLHvbfZe/9xQTy1hOtNxijzTwjLgkmzX5oomjbK2ph+FZRfzf8
VcDmUCz2WGoiQ0+3hYDXb+5yh1V8o9PEJ3DCREmUawFnGqYleqSa6eh5KrRkbx+2Yj8qa5NonpIU
AYAldfDJsK0g44rP7pUKsVxiIAOj7E1JPGx8/cs5VwhRMLCXf1NIfV+YW7BqEAtHJDLuHz8TqtPG
0s67Qyy20n1alnuwD8LhSNTewUU21ybeUZJXT/KCRLAecS6ARwqaC5ckWCvkoBzA7aWAPtorL6e5
ZHdUmtLrNB88B0IzKSsZG5qh2BNkttXhTNodXKwr4+gK/0VlYlPXGnsQ0TJRYAHMTytW0bIg1UqJ
9uF9B9G1IYzTBIzYpTMV7wRxV9NPpd6164as7sRgp1XwB4aOTn/SIRJNUgdgTMpnUrWGlPNc8kSs
Bqzrm2h7loKInExN46ahbHc/0Lu2ZonsyUKz9tho84teKExZepuirCMlS8lYX9babKlEVOcyleH4
+5rYUQhtMC2mqR1vaW5Wgcbix+lJ6TPbClytXqWj+A0SXRl/RW36WOEjbiVrvC88HqvZ6ttQ7C3Q
UEKVI2OdkPGq2i6o/wxWjkj3TV+7J+LTsXgFFM4RKsX1FfEgWeZwddsWTGzczH2TTaMKzfezTCv4
9RyudkdppflbLkO1XjwKFYujMtt+JInFWM7hSJGlYWZiqVmOX+L4jp5HJXWLNE5kDxa2d2FVYuJY
YkNMJiojSj0eZtugaq1g2HmQ7ZhBFvHPcp21REK8dyDOciBE9d4wZBCUKyqTRWKZZKsr2+qu5eD9
oKAb3l64XxoqJhLBSpJvmACQoTN9OPM2xAD6qGf7iaSx1RqPGJhTwitrD/6RE3zYacu63fBjFBGr
G27xn3L4xSnyGBBpZHwYNhjbWxvvyXtWHuURmvgIIQcPviyE7cacSuJGV3Ig0pcyA1wAg06LTrqF
PDMwED3K3fBYqCcnn/aaly9uojLwIo+KlztvpulIN6As374N27p9a6hDlPc6pa91Xsj+zX5bxofl
TGCSn3oQ5zMwdSDCoAzNlJUVWdFAm9AzTDbxR4uuLbKLNLW/FKQOVk7/Zwl1R4Ne7FAGiTT2700Q
RBSVI0DiF59LaBnjmMgroo0q2aPAXNHTf3GtiGaP1Qj5KmGYI0DEtv3zpbk9ZP5RH4ztMHbH4RK8
ZW19jBK1lSDApDQCJi4BC9oJyY6VZiKeVh28zSt5eyVdvKUXj6jafXXhymGQsTw5efap/eov5S8P
42byFWF/SglTAWNTY8l5dPOIwX7XJf4/FRMzpRxdTePq5X5bDI9u3LZF1sa+qyrU4LwJIGa9sU3c
ow83SDFknqWQ6qTS/DRJMFFCQp/ltWG0HebwcItd4I+71MiMrgaMI2AIdXBhhH0B5EGAa2FKsmF6
9YcGAvY+j4ZHIO/9AlBPyNfaPRPTuaeiS/t1rGfk6jRTI3m/kY9p+bS3Glp+HTzeNJo7ocCn3wtJ
sty5ql5nzpNFJsnLubGOQRHkesnE1Jab07FtH97VCiMNDSM9M0OqJdbUPqbIdUl9Warp6vprNBxP
zZVvtJgvNJdKrQJS4zSzo8BRO1nTcaLnOmgSvrJTML3UaEU/xtFrUo+MHPdJdByaLqYYYatbMUSS
T06iyMC4MN2KIk8LQIRR3YMeENKi31oPX9THWVcXeLAZHKiEG7JJ5DyPQ4sbWoy6tVLfBlg/L/VQ
JaeSGysoIzwgpLtJ86AABBXQRnObqIfTUWpXa/KftQULxnya3g1L1qmyrjMgIuOazh6fDaoXCKIz
yPZe21oCU+e7I5tPG/z3VFKJyWf+laT7cIDT/aQ/yKr6FhqSv+dTdMnSImDrHdyiBr+B7hZo8fST
skvn0iLVmdzGyQ2NPDPDnfzpw8oMPkd7w1jyK2EMI0wSipl1j5YwhAVfQGyE6v5r/ZAj9Sh6q18Q
R43skeo3vZFBDHdASa887XCQ4bF+2ryhNDqph1ZCXdDXr5mndAdPYbNdpLBZLdiUbRS+w3/oPOMV
yNr10qUZb6fd1sGuZ9DW5mFpMVDKaqCXoJeoFTZjG54wWcFVkM2u9yIgUBa+UDKNwKX4q/wxZXPg
/VzK+ZHYcqgGFpRTkKg41RoWmhrxISchpUQbgs8vJwiTu/jLu4Lw88m2PT+1G0mp7vAQFT39xI+q
F1O5GeAiT4mEiVk7QnmPRMM9NcEYIveKyuxIXQE7C1EjRzWfETekBu3EDgVKa5+8proIvavuDEGP
P1qZvLtiU3+UcsOpwiTe5xxlvzM+mnKnpwL2F6gSFQqI8tHEne7MqM512c7TyurHAS77tTwD4W7i
OIyYylDVJzJDpThgQfA+51byGsj2wCvkoMk5tjRMyPmOL/uVWz+ftpGg0dGajqB9Ahigz6MxviWc
5sOhqJq1tRyyBeRZs2rMJwAIekRNnU3Rjg+xBEmS60twH22AM263XqWpJxv/nbDhf7pJ1PjOIkDj
xVkd9ehRPBMzZEGnAnnKUWJJT1jY3ewE0V86piYncghADw4pqpXwJCVkuUZFE9JZWfkbgNpmBy30
Mz5migG4hqzmKbcf6Z81HO8MxsjOiYQ7/KTPUiId5MIf5VZjsZuwNWVsm/jR/nKSxFxCkVno35Bu
mMbpp+fv+LWvc05aAANVnajYJbXtj2BL0RUMwCd2Xzmgc9e/UDSc1qOduILC8+S16HwH/toFgmua
SpYg1VA7Rl3OtXh9LIrPPvigSMj0HPzxqRmhbajRr1YvfB4yt9GCY0XPpfssaI81cMqQLvd+LsR8
YaU98YJtKhv1LjASDsBaNnxM7YlKCpTY4epRkYX2HNnAjjiyh4rzJ7ODgzUbu+sx+Q2A23C9AHXg
t6K5QUGu3gGml/TmoDKxfclI7UIOHuLFSKTOBUDIDs+YLQZGtqMko/hYeKvAfrPV6MIgeir8I4uk
v4tJ0pgezSE+/LrAGb73YFGVNEtvhtc7V8/FJJdNK1r6VS8lEp3D0oludUywPVDsHTRfkTPpFzPF
HsEd14iWkyK70tswifmQd895Ov6gakOoxXJWBvLi8ui5f/n6FYSu1jz1nvqt6CN+IQjmtLHXcmW4
Xn8aOxQoFkEqtN02KnGA5RBkX3mqwMYneZaB2x1tRUelVaEbKuRcbgM4HP3nYuEp1MwTtKeRrK4e
ajvkEs5nO8QYcK4d6MjW+OcwxKywBSjKMRNcuUgnmx84WHvv0z+OXx3FlC2A5n9qEGTLlBDTeAc4
aCkZ0b8+0aH9z7yAXtSueTlt/nzC0SOv+z3MmJeO4UmtqdW5DF4mK6LhnSenQ0DPo+7nH/tw2Eux
nM4MiFI5yqhqVVywB63Zm8fLoMMbqYsCcrDZHgvFl2YnPDE6CpmchTEB//+VUxVy6OKTaFRpa/g1
Jazi0T75Tveuaz43Ai5xycZP9hYFaheEuqe8TiOh7Li80lWkKF5jW44JwGouBONbPt8mVoFLd8E5
wOblx+daEiuncUZFqok4rCmXseO2eMuNC2yQDGqYO0jVzcK1tAPojBAWgPygoadjNsdxugstJ1jm
fG0sgVYMvX27v4sUYfFmCwruR/Y/7cNdtgrNVJPfTYh3uL98Lfa9OOUUwNUUvrRe45RpNsIPwQcQ
inhVUqNd0LgfevGQ1ZA2kvxb+856+ywpsmAw8ATVJjzVVmDtVU85inT/gIfqVbPxCoIJ63X2e6Mb
gbhchUmp3LzY6r2IOQit3kH3oioO8hhY5o4Yr/AMbwxAj6z1RYnQLT5WI7SrD6G2O1YYGiCPxH9o
QByBcWBiEyEGbt3EVzQmyo1xxE54V9q8JLo8l0NLHM3um0NWNcOrkLpwYOrqPSlxjhwkv2BRmca7
9krPJ2VjvK2abZH5VUSGXIs+JN+Ke1pEU1Hehiaqommj7lUi+pwdBg1pulJYOiH9q84lkXYftg/9
BejqsSwg/jUa+Dxu23dZNsj57pIMZ7c/3HMZkGXkT0yrNPT9vvrmrYGkn0UbRhZCRxNb8+CraPyS
U3vDuKBwSUNha2jJmDUr80u0aB4BZvYvBBlwePW6p02JI9yr/6mZwM8wk+RhpNxpCYTBa4vQCrAJ
LE7k8zYgGgxVliLL2BOT1SHeUygnfaNarGE/Vxf93w/589K9U2caA6dez8ZT3s/2a1aCOMhpRLdk
XbwyOUCE1bEcOIQg3iRHma3K3pdjFbcYoVmUM8BQiybK0X9vBG6biV5QlcUhgK4nQXUo0y5GdS9h
KjxVQmMWxTV4MzWi+2xRfF59h8zrej0pvlwC7HLBeqqhXJqPKIeyMFhUElduUEH3oRIrwsEQNBQJ
wQSoBG4lTDk8jNEZxe5b9FZrtg0zeBMa+7R4h2On8VSeBkRQT039RZ2/AEKaT/VdGgOYxFfLxzEk
N40xEumAAcSPg7FJW+QkdzAHlUO09EnkiTwNW70dudXHqUJLayhv42N+YRAXEb3c3KO2N+QpY7Fw
dZERwFoGrp/mt1Q9XHugm/3ijU+JIbkLMwxaSx9VsvmAW0rMXkf3P7FH57z8WUku2yeDa/RFKszo
tU+qyzAt3FJUwWg+wmytkKrkF4uSzEukWyUtTa4MFkqfTSy7P5+6gL2PV3WzDf9bSWVqAeirC79p
NQkzFpmfAEGLdoqiHbGSp0wST34bs4Y5CmozPae4mSwyZM/Xl19CSTMwkcCQceX3GkuWTOfThml1
8ZTsur4+oSo6XPYyQ2/yy+Igcj1DmwiMCTSPX10CEf7v+E2zFIysdo6Fe326zQHSDKztnpKJv8wl
yWubP+rdPWq4WIHGOZwfEPPHPqgGbn6XQrdUYcpT+2vzuGYP+JyPFsmgPkiWhI6tfVbPlwoCXdk3
G4dPniXVkbJkSFqtaCcP8zf71ifUSobG62b2fYaYCPDFcG+mGmbM0z8O8EXUW0qh8Ou0AggiI58a
FA8qESOKjCPe9aaWsgXMUmnFg6GrBuC6nELM98XyuM6MnJgVktZuxWF7mmVSlM9pvCyI3axY7bGz
hWSNStKPPAxHdueAiO1tPMGnKhIDeGQEzbd/pi/eRfBjMuwEpn1X8mMC7jc5Rw1Rmkmj7rpjv49s
/HpkvFe36+7C2nLz++QbYz6JnejEB2PI3bhqQ2Fc80IMlsNiJ1jcBJQXEwrv7hVpcjz18regw9Yh
xLjv8Lo+zT6KMQ3+RkHTcAc46bY7qdsDMRExBLbmv+fmKL4iGHSH3LdLYaM77kDaAlj9lzVwSTUu
RrWZ2TjPgdvNF+HFQkCDsWe4mlcu4hNf0GPQjJs9OomdTAtHL3kCoVmmGMCnSSwhfC4wuxX/VNJk
3akA5OXAQQ8UqpXG6utCvmsDtlohmnlaMwKjrNyAZLJBRAONTuVXdbS4suFLstGr7+lJIgDy3kT1
Jw4mv3ZeicTnFKt70sk7xbzHdL1AAoAzIWMwV7vc0bbJrwz8+TGHT9p1KUjbgEMIP/RMQfdKVJyr
AqZZx0fKVM0y2gLjuuBkH3i9a/9m3lyToEsT7qM0+zBJqZEGwy8NVJNOmBzCR8/a5s/KUIhnl0rC
MP6DBRfXgOS9eY83dJnKeCaBdUeSoBRpDgfdECHwt0UFNMrld3OoTP82XkBMWrQYMUlw99mM9Q4i
QhBNL7Sbns42z2tuKiXRkbltQnJDoEX7NaDeQRC+Suz8g4Xl8mPs4q8WbwgOjt8/WZbKN/NMquMk
ay63NVbaDfUj5cLghNTt5jdSHpjTizRlDSb6uoy6tgz2lrxA6MyhdXuOTZJeDcGgie3+nbDYqte6
5ERYLOtFiRjKSJH6g8UH1+R/yG474mABDO5Gz2X4UJ/HU57OPDjawhH1gXKLLoTT2513O4WHIpII
LRQBuh0STIM3YlrT5nTZakdlC/NG3b+5jYINT4Ic5mLff5d+67NYMvXUmoflvJHNMW79l3YUNFMi
k4MFJX+tbIykL+fQuuHA/YsSIzBKYwiFfk5Dnf85LTIx8obZCulLFiBIFH1VXJuuKDCxsxxOfPVK
Hc5IN1/n8dyCviMAK2PjDSe0eUmxuUgkK+A9VYRCL2c1cjZhkKk3uvE3VDupcumFRBqjItu84leC
ho+kWMNLOKvS54umm8TZnA0wr8W9FEsdgurWQHOPBIRvm1yOmmDaf6+oFPRb2N0QuUKE0dxeBDG6
B7LjMBwZVZnZWy1MttDolASFA+c6cjMXcievFKkaHImVyI66bSefKKDXvdp8ZzIaq/+uKMahePzZ
hqC8lYUCPQvyvG0/WwEkzi88KQpYp3vrN0xGNeOd7SJa51xVuzWOjDPnnrgkbPtcU3ggBvetlGAO
FwtRMCsRdGJO0Tya37a0NZJV8fz0bdrkkJQRKoAHeigyrlQ32giqCWIizPrpiH6VfjzjYA/+hGDt
V3k1ZIAhP/4vSSfAiPKSD4439tZG2GzjIYr4b7anynX0aTOWlrfG0zPdgIsKVQrF0hBESq3oS1R1
sxhVuKNNFEOYeYG5PvT3TlEu7FvkCoViATl4Re++/ZqsABTSpSnEZW9OpmTDjZZ8RYMbn5HDkFcj
JEgDeoZ960dhc7uGFZlJCU1bTu3rEVdZrSl2mA40gd14R8creAyfdQCIEw3AgvatvKW7EfdBZHlY
YqZlj/g0ewC3QYq1NWxjvhtOihdpQ+k13FlEeLNazGCEx+b6w57WkGCCtfNzKnJv51pxL1J9QFq0
DnMxypncGgV+GTXYdWRKq7DWcMILaHjxmDmLPgcgRqaQuMTpld/7T5iu3qaVHixCyQnhkXkv2xOx
t17MGBa1iYBIGN1RxpcuNaca2lwzFw9kIeuR9RanWZ5PVXhRe3zlbntAJ+MyPWd1Z85LlYRNLbE/
l/rVBmYpln456zffDoOnA5C0nMpQIlJN++NrmJl+wMuAEN+Ogh+/pf4OuFFIQZy70GHqDiK/Qgff
UOV6BfzJEJyw2KARckp4y6yk2a0lYnhkJsbqTaBwxuDi3fcAEOg8Vq8XiTqguEqL/qCYVCJrXiUA
lS/y2yXccn9ZC+2dO0oEiS7Ln4rOTXy+LRe40CbAKR2P2FJRhBZVEOuZupRorKdHMknE7tksG2BM
vaedn9VZjpLPztv9zn2OUy2Xr9Z4Yhz22a9nf05hMzr0gmU//5qMhwmxrRGDc6tY1PyTzcQQ3wm9
JN9wvU9rzBAUosSWUhOpa+EMdESLICAsUgil0OjkJFFXR6Hfpfh80SrK6RQReluMIOmB6qwq51M1
VoWWKulWnKXRqbKjxnn8h0DyVqThLCHfPW9pQ4RhVKy40A95Owd3zmJvT6AM/e0AYEe9UFYE+AsP
mW13o653kC/76d8q2zWAGWE0OQJY4UZJzdpuCkKdWc4/msBEqmsjYvrRie+ShHrzVS7AIzEF2Agx
Xu+udtc2u68jVeaabrZQdDX8mU+6JtDCuHCC1F4AiUBvAnTJ2YYh+9jMGWXUHXuLBjpXzILJqo0U
fRKVL+l9r5GO7ER1Bcw61JObCLzthsDmTmBCF7GqL3N4d2S/IxFl95Wz/QFtXT02XfYqYmSMxXDO
HsOd3cs2bVOGuMUcs1bCeIDV5vE+Ba+fA9TNMIJZfs3uC5YyslB2sdfpmxV7TE3dEYMrqkS91Qel
tUOJVbjpOrlPbQ+Pa8UxAolJgBHj2cNuakD0cNvorZQ+AgMQWVWcxxnOBn1gdJ2Xd5uWD/ppiBy7
MEfUdvfeo0xLJk4GsS/beNU3PxD27phhn87uG/VrkKWh70lYM2gAdcrYS62/fPjSjjQCibGhXIRp
h4JHeMOzrXmO7FS1nG5m2n+zR12XVRD0cITxmFdocZGAkhWTCgikWYnPbl+pr1GomWvG1OXIv0z3
I4ly+GWyouysTPngp++hzKTj9Akdng/T7HN4M06zJxMJ0lfYxS1z6v/58qemUUN09tPm6eRvPZr7
s+f4D02/ZVoVWIltMPYF6InwvWsiTcV7D5JUzi6L6VoOSF2laDrZEJ0K1TSihy2tPKZZOjZJ5Zhm
QCZhQ2IN0frMPird5z7f1aMYvCK0FRWqPr4oqOqGDwYS1EIbBmgEC87cati0JO1etM+WLybfJMMs
UEqNw2uQbebvDsZpDlg6UnLMyEI+1XJODzAP/NZgjvCCVd2IaL8AmunYSLKYWlUTgyw1qoEZEDWK
OeUcLTKfMfc9BJeUA2WnnPNehgIu6Sij9xaoBFpLYd2TBJSVdYM36E9dYd8QDAlv0gmIeUoBnogE
KI/L1/n7+kz+BCgSSe6GT/wt2z4ZVEHTg3Af23103NDpzgNxZO0OKP3+oYodUSpU/6skLPvIDgbP
7oNxtz22WhDKgXev+TDXTkMMEzC+saikl68XLxEav7UyakTYBD/UiaakV539HLgYqRPKoNEEz0rA
4oH595v5qnm7tVI9sRiMsa4UKhWEuUoQhpKARHuGF62f87FP9ocbvcdP8zt//oux0AvvO0x0dOaL
6qqmLePgY9lSRepyADb6l/+UTGw21l0TrIFbecV4rCwkkJB5Pe0aU0KGA3B7hXRanKkb1uK6Lkdx
IuAsmOSNKHKBuBB4UMhwlr71Hxdp5bnLx7rIlWJjdJEksJHNGIi6lpp/2v0ycJVyB3xygGXLSb73
LIBjzIyIw/oI2BX5l1ifSI+/YXSAtk9P14vpU1Epn2fGqJgREDNCz4MCCIMZYgrBkyPEZDCGzWmz
C5g2MPgpAb81P26Fkn9K9CJDDsiITl3PLqQ5B02Qe0QQ+1yvYAke9pkwLa0QvtcqNqQvo0SnOExi
h/yLg/ZNw6fygMyDhHlUvAGY6vv1GUF512Q6gsaBEnuYkWPTvnlh+yA4WihGFk8ix8zpzAt6t6tD
vfIqfDY14v/bcIVO3J3s6LiLQlGNXBb0hV4D0uQuqKUeoVYt4J5Bvamx5dofFjvppll9R08cc2IS
s99T7RlYKD7z9JXX4jgWtF9YgdIIqD3q/RO432xoOc2uYNvl+8h2Rk1FZm3SlR+kVS8s7v5TrnOB
ijfP7rONhWBeteG+D89PHwDLFPCwGV4vyJh8fRy/2Qck/a2Zp102GDyhpx9BS6dsX0unfXE6Fjxc
vbtLgvQony+agz9+/C4KBCPKPY+yW03ndoqo+YvsE+PGBFrbPt+YuppHM9Vo6cBjaU0tyIpTYpou
BUK56OAhClDUyM9uGNjVnRe7pA7Y/UFapXBOq2/4Zh52Pnl+EsTl99uFUgSK53j6TZ1XF8Lr37ha
jFFp8HSW3zgP/eCFX4fFC3GOwXm0SyO44kbjmc2mNo4Bsg9pyTnwgx1UiJtHJmjjGVXIXtxvWbax
jwjIU45VLUuZAx6i5S8eJBjRtfcyVL3WYLvun8bJwvNgpzUAgGDwIsib8rruoOmxSAkTCM8TILMg
gtMIczu2m8LTcN2OjOhzGuBBrUnDPf/g23Y1d0ocgIux2FO11gtqCSbVro3NCFpHXRGO7G5f4rEX
NsUOEGCG39Zb727aLUzZ0DXwSLrhm6YK/3PVwyYnQKoBewhzpc9eQ0ea2wrS08l5lyT7eowYetMT
8tAs6zxvUMr3u2L9suAGkAF8evkTi1JWBGCSCNxrP4peLV15EQV0DOB0X8hmWAh6tJK9kRj6oVTd
/7Cv80cnJUADoF6LdlSiaQi+rwKrGVIEypMZGOs++WIdHEqPhlFGK23fsZwYF+N+LCStWWdH0qn3
RSmptsTwL8F/H0HrpM1YKS4ci7He07isYsFeTBVieEiXxeA5x6igyk7M20uWSQyXcoIPW8Qp/57U
s7Nm+pFNdtpro3XRcWqBnnKg1S7ZXALaEg/tEdk1bMvyZhhdbMjaRlxVGlthPUDqL4NdIrg0flMy
Rei+gL7yWjmOncRWfGaRNnjCbanoy7XAVMX/FU29lVc78gfAKJUAirHxBitWlwXzBhPgH2e//alK
1AtU/jVcovjVsozw3CtbtVJLRARjG7sjBuB9v62soL/T16Ia5wlkFH0kn5eo7kJN09nxtaeWkaLp
Fe7XUKR7gvKDgOyidWgyxWyytTnMbU/cH40iVWXYHImPppLKY6o+BtZDLVJcMjGBL0rDEfdpf5nj
FBB1n6lIo7Gz+AAHYdDd7ZiN4piOO0MFrTvCeMdQ97uqiBo7IWsfiMxoYfj4+Y3p1vePyU4zgGiO
OSbLwLBx4ru+NgVDXqHFvqEnEtF3fr30V2GjEga37ToyGFYqvbVH7A2uzXGQFuGkvDQFXHGznivh
WwZ0wtidTLpPWhkQn8WJY08K/wMGtlRNB01KgRJ5b2e7Ip5m6GgpfmO5V1OTVHwGeTvNY56fCVyY
li770ohbUHNVRui9DF1vz2rVdbikjYI301i4sddDLVsFgpxKdQKFoMWdR0v476ovET+QSVMk48ak
0xNn/RqEqxnTSP7ugxSmnZEPGbmvJ17AEHfyubonY27QIJH/SxW+LaWJMWUTwWU6fcoa9WFfM59N
kTpFrPXbxtbUTpfe/jxxOIplpqt4Ktrbi7/O1LP4VFeXpr7AGGdlvoIGrDXwwtEzKZTiSCQDwMIg
4iTKmsuXUrWNLa2uN9JKg3GgWfldlZOrI0sYYw6WRg8pNWaqKFr2pf6WG/PpzlnX8N/FrAc1J1Gm
MdPGLuWT/lbIWMFB3IB649EAGCrOn96E3TZsQz1ijvF6mKoaKxs+2AmEYZnu09xEj+NqKfNEbNy8
y5D9KmVLFKEBDd2Uxawqs50Q9E7KoY1uXyGGxYuM8nXEIWwnez44BeESFG0yAKZTrgEdIIz5TsAh
m6SJOcGZEzatIrmGmDx9na74Qz9bl59IhAWKlx91glXGSc/EDwUTkWGdnqqEiA2YwdOkhcpLJIvU
jY7VkHfaG9N0Uc7wDJR/z/FNNUtyQ7e3Twyy9Qy/dxxtVk3VDfULvHFjIQtBv8gVUN0PynaZ08vF
StK3DKLzZhuhQK2XPX5EZcOc0vuFzJuqPSQHjI9Yi42Gik4vtjYF/scQZNBnKjF9OB6er4shYyGZ
VYD15cm8egiG2nS+3MAXmLJx5uxNBwL4vE0fSQ2ZJsOUBxd2+t3FLtHw1XwgF/o4JTseb8wBiXOc
NfEZLPOoErSX8eEkuJ45UbW+wca36cXPeiT5KvDLwhw8gQSGFc+7SkAimQVZP91oa/geDHSs6Q1w
OetTLodtOabuJxote5h/S1id7Y87WGVQKN/fl9CS6m+obPA55xw4flgrBrvz+EyYYLSIyLLMMNMr
l/TYD4JcakkvBPbgOk0h//vdbgJkZh+Mao3Vr9VX/pXSDI13F5IDBGrokUXV3B7ctsSb/7uBCm27
53aSkKsMI3DfXp0QrQCqMy74ECf7a3zMqE/AtBSOQR2FIKMc9y7MSQMngfgBr/Wd1pe32gmnapX/
c6nEgzvnXG3BjThszFTq+Tm7v/0uMwE17rxZb3H9PjGML5RQRCZpeWX3l/zeLfbpKhiBxn7lW0Ki
+W0dggxlyaNhxA7YARicnVOV6+tYxJEb4rI/a/Z0AIwPPciO3LsBkFzG7N9mWdLc5BrOO0/o6WGr
Y+Cjeqkubppx3HazRyV1l5Pi/8lE7NfN5ew+4AtC4NWyVNtT38hBwskYkaPCORk8f3f0gVJCwmfm
bKvmkQRxoA/takcVWM63V2okOLiGCGlwmc2/sWiMqSy2mEamj3pdzynDkTtQ+naWSTpTOeE0jV+S
8gvGjj3wt16iv0ysZczPmoz7GL9Cx+Kl8FwwSUV0vd5wJO4xdPhxhVinCRusr0UuK5V8XipGHiHY
HIm7PogC/Rce/woMM/HEHh/7Exx0t7ylFLC5XSPIz3/tJZltB0Tzv70GE2eyK+qRXRrDmzkpqSV+
DFEhD9vaiBytwlzt0pAzeyXsSWsZHi3lwH0Kt6sJ1MT0vs5HLXAgNMAOhSWiRLLCtits/ho8dnNV
KrH507E5f7CKhe5WV9e7+zYftAH1bKapVT02OUIzRcTnO9MxRiGfBm/f4RzQENHihIUTp1GgfzYb
mIWy88/9zNNwJizoYe/iuv+xTXr+Wg4GbvjL82tdqwMBraVka2S2jVKSMpbguzNWO/9xbYpWJfLL
heLazlO3yHQyh3OTPi9m20+zULmMbd/bcKeecegr4ujznRXe4Lp1saB7NpvZn8dLpHhZzt9ALzoc
qSo8CdQPT5eACNZ2BV9Jp2UrLjZaazBuA5GbUCtXa0oyn3KZkJemDa/1iduAI7O+D170n/sgwGEF
+kOqJeqg2CLSZxUEPv9toqNHSfbld/82xxmS+KOrHqZUmwUTuQvQubodzh0cESzbytu2yyuUA5sw
wLJ4sBte2HIGAwrRTXytcMwzHGFljQ6TpBrnbbfNX74eaEzw/GyrJ+x6Mpz/45ywkPZXABMWakyh
czx3fyBykaJFQkd83/UVF/JRWST+RlpFcimVyy6er4J2CtYcMNmwI/MAKiGtT+Kp9iDqdi8n/96/
p1uM4fZxZIOH+/+FhLfKn6LIYDAnIVFJZQkJEn5giq1B8LKt0xI0/4NLOuB17Iau1ZjYWL0XQhFY
Omm+eL/VNO5OrmBDHv5FjoVAyp1OOUtpZw+ovYJAtJqYjGQJWU7gDZrSbJ8IYvRhMFOKcyjJVwwd
tN3f4IJtOab59YTp6kljJmwbcLoda84h30fyX4T/na8d5R+VodJDKAD1maDLqngKg0NdzPGwm4tf
nrw9O5LOdAR+GQar73dVc0x0Zc2d+3DxRxq5nqoVk5yxjYyS1Z3T/vXUoAZWfGT7lQyPMCgb6DDr
iwcHXM581fnSaR7KplZutQ1leopYa0IGe/yO27aR76CWOwJ+yH0RTYeTZwtmtLCc5I9AKhFw0nBs
JgFeuFY5h1Y6ABKzRTJCSkHUsJGSvdUjKZ+rv9/U9oy09Cqq14NM50GBmyGa/+PJG+m4k8KN6LN8
ahwKS0F3Ihmlabn8fcg3A4PQ5/zq6McI3g/2G2XupEiBHolgl20/L9kTGuSYRDb10Q38zLx2hgKH
qjt3Bi1ntug7F0vfF2tSkHSP5ENNRHp2E962C570WdOWXrfKDV7AaQ+GJrtm1UY51hwMK8hbA1FO
F45iNatrijUfotZ78kzutsS3FdQcvvCNesrpzs+kE70Kqcsr2wEMUrx3cBkDegRwxVj7ggAoEqyn
w4XZB88JT3dVNneie6x7cr1cMnSY1IkCPpuOO1/0YygegbDdRj8ore0Gy/+b+CbvxTriqv03MHsj
uNE5ifdGUC4UGo0MMKVk5qOpwArIEDY2MxOcFVqeFeM5+2ImRNTb2grFzel3BYzD8mHLkKI9tHws
FvHXmWc/MD+50dV4SlG7NIHhkbjKQEdDieLwtzbFA1qy2gLae7Aec5i6OaNAolSFuid+2w+pb1aH
ZQQY8w2h8Gdc9+lCgntCnoYeignbMbINUCz2E28HSIRXn2EA9nzveappUYDKFMVIvUF0qxTXGeXy
qUTC/U4BrRY+/gboJb55ZETWGnzrNfNRDBlDjgR5+pRSDxevKyor9yBy2BojsyzzV6JErqQw7X7Q
EJZ4ktjPLGBrq9nE8RqaE0trFrHyQlG9ayeMRmVtD2jFI1shkf9rTaJvh7iozQU8bIcsG7yIyEPk
uYulT+8OFtqXHm4d/DEZYj3Y2pchOdMqijG2nkPrmj3VZ2xOtHOX8BdnliPIwsY6vHc4Ccu5pn/U
26tmO30h+DxNzsNhIilBthL9/uKFx5eyQguE3xsAAgr8ylp+pEDYvvSo2z7O/z7lQ1g0L8HqG33p
1rZfDDPA8gfGlF4/G7WMVhgn0gr4XTF3Za+vgbmX/rTrkGZWnEPIbrW4h4p54QHKftMSIy3lcP/c
UstxW8i6cE1tNkmmooieJ3+eJuaCuivSvxzyDDimaQ+B0dLl6wC8lPMWewx0ZuKaCQISUj3ZuBoO
auE7ZPajNDPdloz5jY+cxF9YLAf2+o03CJQfh4W4FPOtldTKbP3sQEz7pvU3Dou+jkgVOgK6MuYL
G3S6LuTks6FanIpPLiJGghBuebOWLxg7Kf6qTqJNcrEMCriNSKQzqrpZYL/M1hQRsfJQtsFO+04k
J4j9rimw2mfk8KrOR6NDMWaouEQEisstFDSz/KSxc+nM502mTfm+LvS4DD53Q/aMXSX7heCPBT0q
oxmHLZMeqee3X3ipomEFu4N7HeVwUAeD8PWnp0MkRn0XFps2Z6ZqHgxi3O2EOLZsWRngSqE7be3Y
IloRqoZBVW3rv7ZKB92DlY3j5BcKa6qiqJwcyfQjcnkJNTrDfBpg52xbI4Y5apUFpaJ/Quxlx3bq
evKQSHQVeovuetAPkqEnQP4Vrep+c1YhajjuoRpu6ZliShJy4TwI9x92UN58WbRjifogPYl+4hrb
Mg/UEgyaCInqMxbNJpemQLhFQ6P+gH0h43LoskfJOFdhrDgOdOyJtjfsEo/xuA5qkim6PTpHW9QY
ku644DeoKOej375aH6ryZAgY11lAX5BZpXguoUedM5GFrns+JC19jzcgzpZk6ikS1UXLoYsUy6sV
JLjLxXziVjFlxrpFXMtwVOIUBPkofOqo5zwtlMwsTwjmOeBfC0nKe69IB69WZZG8bWAU2312zbrT
CQOr12QTCZzGOvtEOdNvRkLTfByHeML18mXZtr4iObZy9iAaC8OkXeYKTHAx+kVZuj3QmyPiM8sY
Y7ztxi8O9nhk3d/m8v1lqCryzGkUT62KTjJ24he5G3w9KZ1nxL5mWSSS6DRvUd/IG0cLPT6jKB0N
Gmo1BUikVRTlKmoCHHM2Q09RsUpjTEaiNOUHhKnHzAwX5tuIbQ2yK7nu/Cc/ATCdBbtYfjObi+Ug
N13fRx6UIeQXg0LlvaShfVWQ9YZGE4+HnKfLF7QvkZjKgb3eG5K/3bS6X5e0nFxycGSwrp6Wq2PS
mOHM+0xj3lrQyFqvm34mh+qz5+olUiH9gqdvstusY1TIR59AeHTzJ6TKq5Li9WcjLgQ5YXsoDF24
173oDREd2/H80gi6MyDzlKoyLvXfkkHnLTwpC5Bg7hkMkCc0wf2v9WXVRcCByF5ddopbW5gdGbJ9
3NssGSWy5R1bE0Soy9jmNImsQZ6igjlgsLT30rcZy0sgNbndbmgf6BvdUrlSoxQr/n9QCj9nfcyC
ycdXK+mcis+UJNM6TXs2W0MfRVeNm2qqtHQZbRtJ28HI1+q7gZuT79+xEkfrqp1fGRMhYdCdNMIX
iyUO2bM+ieZlYEmH7aSmiJoS+hKkT2spZ7vA2TKIV1qVwexRVCjFurq4I/EqSsOUBZ/YD1Xa0Prt
bmWSEegXQl4pPmeQjIMZLWGY8c2SY61J5zMjDQ8U6DKbD/QPnHIHm6rrOUr8GDt0W+bLvT5nJ1ld
Q1XdxqGwJ+yMSy3nBkkK8NUSHdX9t17Q7VqlaB08v9Piozr/z7aSFoNAGlJapTDyCmHna1ECM+wT
tkQgEmltyGaT12TMvGfsf1IZe1LYJT2oUWKamtdD91Rmywyq8Z/F0ApwULCagqIBam+ZbQ6VTZJ6
OYWS4Ug8m0wvLbVLQ3TRUDVzgYNVVRWLFGYDxOuH8Rz3k4v0fJqm1zPF7ILDcnnTJTw7OVN0ktez
PAuo9FRUQYFdbEwcoWwyrCl8orKyAglJwluYArW0mn6e4LCfwZVu3IBEMI1A07WWevV9N8Wz8pW/
JBv5BRgzKdVYBRfCQAoRgtk8YzN/o3VOWmMieooFiMlHRb4LGKVkj3vCqgt6c0Zu83TFu3Vwl6bz
LX5TRXBKHes4Iq0tntt0nLT1OKmSLvDzqG9QEZexIAofJtPuBxqHbr65gQ4fom1m3KUL15RB/Bjz
uv7/wDES1yRg6mD0v9wDORKwDAAiXZOhN2bfNAqXn/g8ukwZLaacGSEFut+xKeQ3ap5oL02K24l+
BDjOPoX8+641xULPbcvNum7J9vhl5f62cdCyiXp2SDOqJiOY7cdQysNLqKGmp6i+S8cEoMdZyMxk
peCBIAZHhv5CaR8tOv65oZ/WMXHS4SlGq8VoecSWwVeUe7/dxEBbpGOeFOfmKRldAQIflIp9QcGf
uTnh2Y19XjwDn3B1KNu6zH/HU/mNaptq2Eo99lYrWj4HWgUgfAX5GICpWzpEBD6wyF/6DuEm1VKq
odGl4t+WhxL3XnCEYQH0KSgftTpazOEJAYu1OVW0vtgiOa94fJTGsTgssSwZDQUcvWOhULWEG2ar
MnASMeMYXC5jiD84mwLH88vU6GEuZ7W0g5meIgA4TiO/5mmSqKxCtvsuI7ogoTFNYnAnMoyvH08w
iWJAtC3dd4hOFzAy8ZtjscxUSINd7eQWyCUFWvYvdk7l2w9ssBwHegnmIo2vuteKUfuSFSPx4j/2
pMXczwULFqNJFtOwr/j7KK0vIWE9Ht5H1spcRaPvOKy6h/47AIiADZIZ3/BRNll4N8j89O+psA2P
9+1ZWRZzu8U0qdzXeWjoDz2MRR133Pxcl7dWfnaYmnk/IQi50Ftfkw72xTtNuMefQb1s1asSjAy8
f+76+z7hvZMVd6WRsEbiqjSVgRLGUJzytB9dZY8Z11A7vC6hsRwG4Mmkh25YtLXTTvM3xASB48Wi
gjS/SFX585MMa+5EnfNo/+ZK1A+QHAeH3GUUlHv2sQzK8U9M/+LTndGV/QslZlDHsPJoP+A1ClEq
ow/xW91SNwlatMmllKhcU8oYC4nPp8lcBrYh+a9Bqi5OOZVAAjqGbFR2KivQfTOBr15oHUHqRa8R
jjYJ9RChIeFWzOb1SuGjFtc7GWFy0M20XAbBJRjmMFLU/oAl9ffe7B4d9Z3iPVk7f5GbzHgCjc/G
HgFUWrNllxfXuyfGoyH1Ln8GVG/gS29OdDgpv5MHXmfDSZwwwaslU5z4EEBiT/c3CB+nfYZX/Luk
qfSx42hQh3sLk+hLF8TAlJ4A9OStupi93u9HyS/k6nOER+XgaPJeFt3pkiM0ndrEW4ymjKuKQo7R
4Y+hnk/jhph+/ihkdZ4YW1qm8nL/BQOXq/UrjCwMquXPuFHT3Ukv5jAf/rQ6MirB/uN2IFlPxbfL
9JdI3WbEyrZCiol2kdSHIm3cKIg0mjhH7DWIb+qWauwmnQoD7yKucVBH0huWQ2HHpDMhCNx9PFbf
mb8nusCtE4oUgBL5LuPJlmdIywhnOv9iYXr8V4p3zJOo+VcVWxjQG7XDCyUC5dQoEFtk6Y31EEzU
MKGC7DT+EKdcgaLRMuT3E9y+VxkS7b+Isw/9TyshIQHAgFJ2M1XuxNS5s4DdIXbDxPD0XWPZ5zwI
yIaclxxdTebkuCU5z+DR67P2Zi2gIJ5wp2khhPBBxGMraBPx0BxriKuFW+wYegdrg71boxSBHIqN
o2MylekkyMTMBa1+7ngOpKAEujbu2nyqOOKWBxQGwDOEkbE0ZuHe4NSiQli+h/6QKnJuBqoTFt3x
eaFKUXIcZoVyv3aSWX5PU3Ff+e8Cp+GsMpRNg9OQflbpyV23Mz0RWkbEh27CCUby1uQYgqwLnJAD
iuUbUU11K21pGj0Vs1kM03oIhQ+KNk8S/yxKJFZNL96oaAy8jEYI/DQebZZZKFQmGIef6S2/ZXGZ
8I50athapY7FG2aCSoiqg+FCL/I/Q38StbckEtm8hLpxEeE64emmEiYi+d46cUPoUq+/mkcyflnd
xTmC/6epV9R/+YQ8qNRZ8ed2FCphGy79v2n5JYPZjsMIUrlSIYMu5Mj7GK96RgTOig11A31jqsSH
lT7DVg3XE/2KuArEkUHov5dJXFtYYJIRae4Dcbr3kjpsI9u9Ud9kDj6wDWBoDaMcHLdzVkf6kHFR
FWcCSsVXf/ytw4j01poB9eKdS4s/Fw/jZp0FRWNIGFkCbVnm7Oi9fW6jSOJIegfbo7TdY3HZcnmq
rfdzLIyC0aaz7TdhCNDN771h2ocj0p6BiyroUzC7ZttuUJYuI1pROUOD38QBHJO/jo+AL7ih7+zS
KzNXSvKhD1TK6GK/KQevW//Hm8KUAQuCNuX7ETR4auH9Su8oFUPDofw2zX/UVkJngTepspqNalUE
g3JnBBPVFd59Cn6WD3N8KBax1/E8Q6rvI23nu7ySsbFOFpiCzB+ZGDo4FosnZzoJGqi5IO04wzo0
jAAEx2OYrtMJ0WsLh49RK+GGBPESnFFVD0+i/WxJ/egK3y1X4mpIBfQQ6YOviDy2CdtVKoDHyOQO
e16abHK6Qilpy+VXiFMS46qpZbuVF26dQOVKSZ+I4pciaGJNjGONSj4dm8FGJitVBgDkcZMKi1qy
jKdy9O4wUJeB/zjoR02l/PM6IlN0clCxDlwl3klzAme59BU9VXSwWxsItaKuQ4pJRLPreIhR6CdK
EFTJgPMPZu0nBnRwgkZ3d2xbiQYJn3xtbhAtRFYY4zrTPYGVBMaz//SPRqFpOk73qA3cuDA4C+Ay
EQcui0rJJPrOLtkMxGP0mtKsNFqxA1i2IYOWoJFvwrGUZYbVrKYecJYvI6pQ4DB2KucsjmOmG/2X
tILi6/KtP+pF4GPas77Xoz4BtW1htrp1V4GTbhmioMtWyAVpzWJnQi/S9wVSx4BEq3OXbPwyG2jt
pA2B/2FVrM5e5L5YGo8M3gLID6fWZgf+FdbeE4oT2I0zllbAhGGityB54AbKYcwIQeB+sF7kP+Ms
/f4b4gw8B0CQ/kyfrLUPyFWDPhgojJf9n/6ZlmCTKyLPyv4li+fNP21NNfIF1KNayQ5GxCaos1NR
lXdJ6VuDR4TduyyUIo3KwbMJDJUJxpxphAJkQl+uNqmFpHMxRx5PVAW0IEAsMpGt4rM8anrQQNwX
RAeXmttmozCjXlj5VzJrPqtaEdOPrU9u9oB+Whx//N1QqFR/CGk3mGaiOADPkI/wUeWIpIR3V1c/
WFSp7kjniKWBHFam8JWAEQbUBwonaaifchcyWv2CTweGYLqlCFNcjFg5Ffoo9J1VQL2HbEiIAnOh
VEL1l2/jP8e81SeN0oP2xxNTpRVLySdOkrkFM3mL2AEHp4gR8yYdroWsYdYOzanBpFgoWpUL+6qo
TctB2/4S3ImMIxfFPa6VRVitdM+5klUNsjnCOLBZme7Dlp59c4rFiHFqO/zamZufstZAiWprPlzv
6Xs/N/jpQgDOHPSxECO/bSk2zSPYwkz0mOD2VUxIJ/ga2o0b1hz1I/aKcbcWlw98GjZGtVz9RIWV
+WPQYKEDayxKI+CwRU5wLOgN0mKkyzstLYnZckOCtM13a5ZuJgjGCfZZ8oRR5UF/qKOHCg6BVpse
jOZP5pt3MDJwE/uCKW4lb06993EdjRVLnz1i7Q0VSHgfbvXazYhwCQWkzijAVzO0FGRiOg2fdSkz
r7VmPCZUq80zdk0gCxxtbp5X5yUHOPbq2xflvJTbMSgn337dcwJaTzbUfVmpl0hBLLKBM9WKU3qa
+h+GxKKG8+VdgUsjfalwSjx+QmALGy0j72nvHXvuteRGCDDBb35+5oqaZFcjRRjzamahfNzL5xTv
jTwVdLtS68AgAB8GuUY4YAwcxtL07UvVkldnXq7bI8cpUUpImjmUVCd6h1Qfm6F/tA6GKeYtvf/9
35p+lGbyPOrHDrOX7G4IapmazpvAcDWsgxNocRHicAsKEgnrjZfnX0AokW5Y6gnJvr13xyqcev0m
rO3sHpywjAAL8X0MqozbLsGMx2aOl9+61iZPtkz8OhrNCn8L5kG7kctfLFckAAUynldrTJctqn3+
nqgRTf8ptoFPZEIzuzTKJM+3HZ+HTy98k1Zan4hEN7Ms/G3p1vRqFYugRcT0LdShWwjj9g4GOWkj
LoB4usOMhPpvwK/pUEs/8PLgZUGhAFjVjQcVvNCTXA3odMub3ZyXA4ABOHREOgwh6BIjbytTLeqx
RnBiBGUqwo8LIaxMjR7mhbfNwHSMVM4iztvYBHPtQTRz7MixWKDBpHYNcKkIJzBPURjF1kU7XDlc
TiyIukmxOqYyAP5ewaJDVvGTpvIq5kasMDlo1gjAant60cvLj19YZ9R1NRcEAYdMg6TbPBMkGxig
UJh5kBQlvPqXP3k/3nDbsXMQ6AwMOSFw6eFWn4gnBuyVB8Q5nVMPTn1ndfMnJMni/DYp08RgxJay
7fvTYwQ2yVFlWU8PL8DrWq/SyUbGWL7KJoaO3E8CNHoTiGp4k6buJFtIeYM0+S9f04f5LjMeli30
ubUoh0Va7kWMtUBDN4+OcC53wjprrNaTWpdfdIIbORsUeuxDW47LD27hbc2he8ZF7iMDbVBgGdPF
taESamRHmk8dvlNyrWdRdbpWY+QFTwh4YdHi2ouis1MIjQDeqK4nAaniXY2j3GsQq5o0CStB+LGV
S4SzkQAqqNRMJI4UVqJ8c/TyJH5al172MR1WX932iHCNKo65qEgYS+g45CFUU5HqELJa4LE7ElFi
9AeMheqr6FAAbZANsmLH+nztpBQ8d0U2OyItRM5abBUo/k+mjImNykccp8sgAfwR6OFzSirukl6B
T0Wdmaw3N9hXlOvwVu6ciIsMwdhSaWKwjIMgoDIsYl52CeYRq9kpCWuFTd7h1csqt59FCsbrN7/6
WAiqzJm3ZiUoncdnxHGM5rEfFSemJeoY3bPWJCtG5ff1MM+cNtTyPtExZMb7xAYh7WZxZBBHo16x
qRfqNByNjDama62jWvMMgcOK3GYqXg9XIcvwYyESknCjScOuWMyqZvq/QniFQaAb4ZsHaRpZbGLu
LcGYVQu3n/N6yF/GA+3QhuhegE1WSHZatFdgjBagnIP6cBIKR/cXUjpJ1H8o0VuIDzdca5/SzYVD
KJ/RixnFajcGzk1zsm5Us6gk9ScOQ0oZxjAq5x5nTyVY3XZop5GosLeKcMWDMHhMXj70iSuUeRcc
FYsQ3iUvlpKDDo0KzXSlBuxhxxap31MkE6SI67u2G3UGaTuHQcg9fH2l1uLoduOFrKcjQf9BVmJ8
L522b0ph0vkemZShr6H3riGtd2zMYOMEdWIM+7qpc6X8xz2hTVqF/MqilkrEFK9dbrIa98C2CJ/Q
WKpqGkfQEZdNbP5AUE1JZqp90cWSaC46BBB49Y4wUuD8uQa9vaO8nrNTTVw+m1VDJLAAHWWfdcuG
h4+Ym5IDvbJVIWrDxozkb+nK30YXqobwNi99lk/hSAfDk/VxPaseDU3wCGVpYeBRuVM7WGbuTFUy
HNFirP52DhPcVprNBG7NNkAej6epdHIU4QNB2HHPQHO9zPSdWHMck3Xrvfj+LlyQwF3HGc2pa+RE
oI0XHTJ2YtZpoM6I3XEJ0lbk8RjriAy2EUsH/+dPouq3xbwwj0Y2TJSOThEMM9RQrFD82JWjyXDQ
OCq24gP8aznTeZxR1nT3wzl/bnwNj3PLoQT29e5vTXFLtMWJ5uCFpbbjBndHF4N/RLUJFBpUPDC/
SKxxH7vszhTjBfAqHkXwPqAh6vRlUExWokXH1ycmoMIOBneVzdu4VkcsZdqdcgSXoQTolTwpJCJg
Am0H28+IksODRn2+HHo+/Ak4MI03UPM7/6r0X9VP9M6UzyGQwYyfMMLJZU+jy8aykVn7y7kFOHlQ
tMWbpmrJST2vwphcFZJo+PX/YmvnrQ7c7GZdRLH5U7tMAyVzDfBqxsL6gZmaYWeoi5HloC7y4DTI
w0JB8QiF4+aRRP9hO/f9nLeSEhqZ2+6VVijY0rNqDjjLsCv186B69NeXYKVZMCZ8h7xgxIIsEDAS
rmNsiIkrw/PegXorD/QhzZGoYvQPgFBTN5lfqggw4Y0EUPK1S1wcORfSeZcUCFHElOUbxJuENt2y
jHy0PI2mNyBFAkuMgE6P+oZxnrvdHpxaD4lIOxTK4iEpNV4azJy6k5acfWipROe1vpaPZ4sGZHnS
QTfdBsx8fihfc+ckfwtU5F/WHBsY8K8ddM7+9/XNlrnTArcyDBylgDuzS1csM0MrqP53fB37IZRv
4yb/YVCZ6JbZJftFxSPm3eWZb4uZ1dxepcm2wKnqQcr9oVGo0S+A89uYSUnnyqD0r85MhhtKAzuz
b7mYB6wH6RNFlpe1zdBb/oq0mmXn+MtwG3BRrr5f+Se758UWipkE+/sccg2U6Ti2KgTF4ikzMBby
96kC/ohAf2R0uK1lnXC4nil8sBtTatXR/4Ln7O6Og+NkUghUqmr65OejgrUBDSFw6luqBWiYW6MD
5i1E/ucP1/ydcZoZUR9Dqnh/sMSd2AbKjvI+tyOlnVV+5tLTq5lghP6u37ofexzwEdufI4CB9hEj
1rlsR2/qsgs0keDD1Yy8okYloge3KoDHHpKGJ0j3hkiw0BCrzwk/5TdtOyT3MXgN0KoXuZUUqpYw
6a4h45h2Am3WQtyervpgMvp2DLaJy/kpmveY2AXs9a3TacJPPmrQimtzCoAVY3kvKu4lODE0RIub
vnCQvWxmnmRlTs1HUmnBt9/zo8BpIXcms/nkeNxZDnC1wbL7Y8ZNAbU4Fk5YDT+aCiHn4Nd0k2F4
NqV0uTdNU78pZaWUN8tWYA6s4i/3r4g/EQJCRY4FoV9twA1brt92pI/5KOPQwT5H9Ej8aY89DpXj
Gmgi5xfdaUSYQkDRNGuRJB8DCr0JGQSFP5YeoSIpNOUhAmyCdoM7aBHMymw1+Qq3mF2TE7TxQraQ
RsyZ5yNs8V2kv1/5xDobzd8tJMTv6mefPwH+mmwlbs41Jhz2GRhz1u3/gnLKMB6cyuuRLH39sgNz
ZkyVBc3sJ4Hy09gtbWJCUhOd1FBrSFzobbdmtAqV1d7p/PDE3FqgCu8vTKgKbfRstGF040fRMd/N
vKpnqAg0eWpa0X9l/6r0oWfpPWF81FnYlP2Lx43FUODZgpmpLnxhfzk89l6HAugQ98eWLcoufd30
60eNmVbCxqGrQKATJr9LsnR5gWCTpdmULFs28wbMP471/Duvexr973Rl6aQ3Q0LMgj5fAUu7/Iyt
Wpmv138dNN4C5CRFrWrdRAaKq/GIyfcuHeyavGPi45vkHNHObhlsrik48JpVbvubjkL2UBmO4MWi
rXkPIWP+R64jgsOhBNaKBjGrMi5b9bsmcD/BzwR/YK3GltUwonixeELdiZBMukLY06FOypSaG9c/
j5+gJTljqN+d7Q1L/uFpF6/sDf9OYFyEZvO1KDLJQ0hrdO6qTFaR0xWQiRFmWVhN1dwoDSKOzbNi
FPyY/wUrBIglmA2eA9iVslfTmu8vdNFdQZrKPMIMXsHMM6YkxAR0tZ5hm7YR0C6t4DjRiMW1KZVv
tYYVkTrfAapGizPG7scga98rFK6GEBf47yKPVFLQz0aNG9r+LQqr126Vda6+BKuJJ/f/vnSrcNn+
rTDvwSU7zOxsPUdHrTvfvvhEgsW6MkNdVLkF2FdsL2qmEgAsjIZpye+Q8ysn5/YWykL+TCOHrajY
p/vMERiNeWrboa81M9vaGEG7soDYqV5H6FG83ZVQO98JNNZLBAUCSYIQXTkKPwBDTokNLLwimde3
HZGQLFBHz6sj2XAikQ7MFHOJzPOlwkE6Pm8+Kxz9Ev5d/7qRcfi0SzX8aqNhZR3NI3SrI73XC664
7D7zl+a46EBjECBcFZtbPvobuf1POkRdi9ND7EO9uwPvAnrE9f51mZDDt+dtKVF8GaAjdd5aIM8i
YEeZPNn7RDzRrn7OIFB78C5dV2dsuyXT1XvzPTnOA5YaOzOKIlVqOuzphzh3pm0wU9HxHBL9l6fa
DUQSu+hUIJt21q3ZLq+upc+3kIgEfcOxe39VKn3JPW37qb0K9cxnQOq4Qv+Cgiy/LgbsPT3Kh1PV
c72nwUrzqbOrY8ngTh5ksgAF7DDnuJGNw/7dhpRQutBIAvjVVtCBXOLgGb1XC5M7gjp302Tz25Od
LpE+g5XabkSaPs+bpQwFL3k0DfI3Tl3kkqlE20S6fDfMtmrik2mRuwvvu83dSD7CL37QHVDa9V89
D8LRsXqka8uyGgWDuPsxT4Z6s0OudXxQvJukZeleRy4VGtuTpA0ZYXOqaNJiW1gFOE3KEYiONiXh
F3Bz5EzvKOxjseZHbSchs2lBhfgQzSl4/ejPDDDbUBgiW006O1MEalCLhvLHk+oJQjQ7CtsqNE9k
oicsCJkyJQZc0BO2s7iq2mg5zBDzlQ5BACMUDhUVuBEbFzXKuoZIbITtuxg5yTEN53gwP5+TjpyQ
6Lm/6vNZU/CbEKTmXKMHNomthNPxJuwdKox/UyJRCj9GZoz0pP6HnTDhva4HkERSDMCcRYCuFxiP
uyYMkmFHTALiErI20YDYKPPWNf/IGhLjs3iu0rPgMB6b+ZDq1QTkbmAQ/4eBRv5uf0YL/WxXrhkw
59OOg/FzZXlBHx81vemTt+I93PQd8i1tBAeS51Y52tt8rX/9EzXLlkfJcDWPFum0hWt0422HMG02
xWxhcldR8n5npH7Qdq7dCDrYEAVqPd7Nm5/hJkPY70R7D1W/DqvolHtKv58HyMtlAKQSfLfmfk8w
91oCUpXn9qlDKmvtNr8dt8epZWlHO2RBWm0vgtx7Lq/gmSoSrq/rWcL+ehb3ZQDRvDUAR2rhsrPf
AHxnQ43gS/L7FsA13ErdPkhuIwYB2Yvz53h4kwNIhyTJ44u43ZEl+fJxq62VaJ42n74VPCXGZ9Mr
39iVrnCTZBVO58Ql7uxhPj+6FQUK9qTYvo5JovjraWl0jMjUlZL00ygHWCfMsJ3LAumsBl31rS0l
WW3Iz9tCho7fITcdZMubdLu7qViynK5twlRJvx5bGbFFJMKPF3pfJsRLvZBXuNj6PRhtqSK7fsQz
FLY01+ZNAvGeg1hVAA3XbkWAopmbSQdivOWthFostd1SRp3RaznHDjocbgcFRiLhgEkZvEhZWxTZ
LBuFPAV8YINWjMImLMa6jl2KB0Bg4hThNAsaMiMC7wXj0XwFbJ8D1FsECyc1qzBOGZV0fHP87njC
WfQVkYJ2979zX5UxqlMROiF92TNnzrCCUqsaYqXoOEzjg/saUs3/MSOaYqanM14jxbnDe+4Zkzr8
8QDIhZJfW8T4nLNfN367BfdlQlRMtla0YsPsNg0XVKpw8ki/nkc5l7IcekMZA9l100iVQSebWNHZ
m+wCiP8gxdJ29CGc9EvrM94tdvYylv2It8kL+mMpuLmVevyJwJNY3FGW3ABx/dQBLbmNoSWJlvmm
/I5sSts4GfJMfVkasi39HDTxwwIE1LjFFlcaKrAEub8XswxDxVR2feJdcHjQejWOSf7KfGy35GVE
KNsWMsAtPEh+eyardEY3extZqT5vnEDVjouzZH1szKTTsyoGE65CIcwMmW+uUv18cm1i9sR6uDxv
3e74kfBuxF72FPtgTIO7uxC/Vf2IdQECDzyYaXWtpQdGq7z+usSbAj1brYE+vJ+SGBjxvhMPkUoH
jt023Xoa1UQX1sHFhbQmHPSrr92E7CfvEZGECntrWK6Lt0a29gRNilR2dnji7BH+y7oZEd/tzSLj
JpatMUclG+aj7wxh2j+McIlHxrmE9k13P41htB5pFTpDwmwiEtFP/FQ2IyvUKIG2mk1gqQ8Rsa6c
fvDo5e+wj5IKSggLLuKT57aQpqK5zga8tCOdRMw1QLaGno+5qcNKurB9E1v7lvCbi/9+yVtptU2I
qiCq6xnS/fs/10DhgjAG0tWB26YkkNzqchRDM24vXsW9ekWUXInfIKYtM0tylcFxdv7h34zrMsON
qeahuo/O1zpI+Vr1EK1eOTw7LFc5O73uk9VwioySiVXvUfFqLvaHBulRZ3MOEu4dS6WUdzBK69fJ
ZiPqslGt9slpob/FR3Dc269zaMY0nMRyGq5ua8D72HbPgBZMgqUriDoKkkX/thGnihhGtRp/exvx
LDLHISZWXkm0AHk8IrDoX+/MaKuR6Rs5PWi29deIKzJ3M0l7QlEaI0U20k3FVG241XMurIHRYzzt
+O9p84a8b+AI3SihhXFLgNkBAmZad3ZnhWvm7YWjAZdKpKSD3nb/5DOdfWy3XiCJm1vpu9OtPNAB
LdlGqyUPhndd2lw3vqtedRk58gQC6E+SaLltOurfICtOf29zC+a8ufuu91R+Tnymakey4z/qc0Jo
sl1IIKb9MURHv6KkjkuT6t96FkPe45pN7FxoNReaP6fiqrMJnRaWI36dRuknrtXzL4xK3RyhBAeO
u4BSAXVi4/YmnnUwRUjUVuKDnvKK6bLDaopXVi0UdGeTbO6+Yl7wphaWY62YJHp0COYcxr2m1CWX
DZz2EZW8tgzwjfivdNHNx+2hbtTMOzyBZ3H3JXV3CkEf6ODs07hOsQYypOxI8zhftJMgcL/8Gpyl
P7VW4fyVpvV0iESAZdd7pl/My8S8dTmeyU8DEUC2Gxz4weJNcZlBm1c/C91vqRhx4RPdoyijq7re
O40UUSrREimjAIuEPWCya5KudF6ngPBLkYQg6DwjLkl9Gn4UBZtJ70ZfCAwAcq0RPVk9DB6+j9wy
8xzrI6pWhfXb84wso1YPOkN6hXwShZqwZuS6kcVHPLNfdoYH5s5whgxYXkjt8g+EoPHJ7NwYHXER
wdlnygzeZOIE3dWl0M7CE0Z+UMdKetQMEH3rWNeZ5DZ/zt72/j7fdYyfaQmc16I26OL6z5aQJl/s
6VwCPn9rucqGLALfXKnoB9LuYAtHBo68ZMAXROTihgqL3f/LRTzLsR4nEMqEcKm9UIwGDkItTTFm
aUsvRI1tXd8igNjVX/ic+cVguYQVkwxi7N0ZgjDyJYhsYEckwnjyy+i2SdUQBOgSiO9h6CysUJ7v
3KrY1ZUqBraV/4xkNMUiQIMRRK2bXXPNmptMMakgKXbOUWKAupRaMMmw6BlMcq3OghutVC+i4zWZ
4Y2dmdBSXJggdyms6q84WK7DbqIidT21j7Qj5osutVY+B/x6CWDWOK/4egozrA9bBWz6lUu6Ckr3
TcH+ETagk1M6wJNyZrxpiP8nTdC/0Vk31OUQp9Nr/AqbKqVczHd8Dln1L0AK8KDbS2Y1TVCbR/jL
VNnXdL5nthq1bGNQvapTuEBce0xD/fgIePbbRiv4q9gB6cMOXbEC1lMjm1r9wf6TWetXz32EeWSA
fUMMXIupJKJq/XpE/eUW92CIyvuz6B5pGv8/eDEhANkRZYKgfGgKlU6Gd1W0T5TlsAf7Bh4vFre5
eN/Nu8J+4MHt+HVuX+/WqXsBx9lBIRf/Hkth3a6XX5m37jWANL6K9zF4mb9KG09QazQF8wbklCdd
0S8aLGgTWViyuI3WC+WsguWhclJ6Zp9iSl+pEnht5lHItZD3UUyCrtcAD+stcWsiVbK3oCJRo2eU
Crai2iWVcrhdrhaJTckAQqC7vmQlDBwUMnMPO8K6VUvPZnmLUk++cBos37UGifq/tHSTsT8mrwAK
aElHNiZFZZ18z69Y48rpENjHHChWP/87nXANy55QlzDitb+1IOTWzBo1NJYHN+JFssKGS50Bw8W9
wmG1gX5BfzoW3do5nvaW88WApcscPb1AlI8i6S1U8W9b2SVFY/J7d2+qD+yrR0J8N6rT1/Svjozq
PbEvtodCZsjRcmtQsiUJA4BdibukqbMocwhZYuHYDIEM5QXmSuLbu1UXLqjp1mHsIDrv2cohM+yS
+IW+GrZEhC206SA+zef+9O4BctDirN4oV5OKgXaaPZ5T7CAZaNREwOPgC6CBj/wJ9h2FWJ+XtfDr
QqppfMs2YNP71vnVAJqkrRJDUecX0Qn64l3e23ExTsWxf1/aPNHvhb1F78zKNQ9mVAyGnMUKEbJr
6wKBo53kSxiAZYwNJU2wlkQwSSx81obsInIAZ1y34Ka0DT+c+Rwz9PaKHntASVZ4rv0JoyI8f5cQ
ZXynnuMs/MQHRfF97R7s5WCFmZF70l3VTnQb/Qy/670nMWLXIvVZVp4gLON8lwM1m7k1kBgNhxm8
EDDzDIHuk6WzKS6CKvDsEJdIr4JAdOfiAsqZkVZvUNIJPJiAW9vZdUz6jTbgTYS40JIFugph96zv
uWL9LUY8T0Nmj9ABJ1XGPsO480mepS4p6U9R4cMr0HOPzolRfNPz4iKCIXT82bOQxw1pQiJnUlBL
WeSvsShzOqKfTeKlcTbKkw7r6iHdNPkjlL5JQT8ziZCrWMSfKR5KT2xxOea4BujuoO0YlHrVBgy/
TBPT4/OUZh/zfbKqHhoACEhQEqyphzGvgDO15yTGf6icn+X3PJOGBTIzSeN4Oxkl+KL7v+DyNLq3
4IS26mlfl8wMK5HFDJz4pBGW+YCr5rmY8W8b5v2IqmYIPJyajYQdNrJz6sta9EusHKizuFru0GKQ
XI008LlRzjJyLE2UqUHlu4fOVjCxyUHmYvcCpWdoPzlkEpMYW+MXhiFTyUjelsAqNtrlF1XdmEwd
PmL5l1Kce62ww7juo28llEX/CQ4T3haLORPVbeVCJb4xb2BBBSJ/mGB5a+dFRXA58INr9enoHYlI
72Y496fi1TlLO5/uplNqNx5EkCfGGVrQdWtTFVDC3cmZH13AA2Echylt8aXIIOCD/ZSoAcM2apWM
dXrPQpfDCyzqIkaRar8YaZuZMVY1SWNrjPe6ZpQ0qtMPz+UeGCTRk/tqCEtSHe9G06Fab5n+lnIg
tJE5ZKnsIsTgvXQ95jyG4cFjvQPQQVNuYWW4sXcSiK/Fos/fxvHTXAJUNGJvf8a6aza1gRfzh4BZ
B/D3FFt6W8J5PXUi86X0AP1ezLejI8u/J2Piqm7BXBUJG9i/ab3Gil7bF3250mGF93cqVfa1KeOz
GnXo/HCOmOQBGR+Xm4x408yHACyJ2raOswS6HCJ2tZtXLOMmxS7MddUWvdC2vyYqIb9lvc+hcY7B
FIzmYYKKtDLCVIR/6mHbgHliRv//xSxatsy6dE4xUvIgyLPET3djAOUsFMxVW34eWi71cS/2u+Vj
zAC8M0KtC98Z7YaOHJXycMjp0ct2KHGNjuNyqQ58yDkgsh03YF/CBpWmwu4jFrPVCjUekDrbQ16d
pBji1OcububDKRmvbI/vSZuu47zsvWnu7yuxr0CEMxeLaWlFbQxW9w61H6EDrU3f41Rl0Hmqti/P
i1HsThPLdHd1b5r39Z/kquk0yyubyGuJrNLAxilKvfO0xKVKIzt92QI3gN+PA7AcJZf12qou+lVG
GNNEdAK7wGL2KHLMcBGqGw6wBxzKIzPOeR8qoqFEiGfOoo7EzNVcsVtUBVpv85bUTABqp4uD1xWV
ciGzKRpoVAqkcbmpb9xdtttFahZFsDUT+J7vGgaIuUtfouSKaGKiiTmdWeVHJscf5c/nGlX424pQ
ZeSqrQdbsgGVvqhiRBslKWY0YWJn9t63qFkYJCfMoUT90sdra6zxuy72A6dotaxz+eON2s1vsSqW
NcwGwwrr0QDtxvC6OE33FGKRTeKg8l46fvtk+55rbLviedc4BefmwPp9pjcW1Rw2d1DQy03QHPaP
/lH61AhWVJpNAmaZhnC5bn4eAF31UJkJE6f/iMl4khfM4pO7GUzES7FH43/HxM+4m4yhga65zE/D
9aOhWLYZlgL7RAcEB3ycXF0pV6ZE+hFvNy54UGMFbjibMzwy3VuKDl3qA3QAqQiQuCbjKidvR3kx
JTgKMjG9rreA4nt3cFEij2nmhzejbV13DjRbc3XZz1RTFBrQEff96lIHWmYgh+RSRaaRAYNaui3d
WMle8uUMfEplsiefBP5Kgg1Y0hbNT2OdYZT/rGXwMAe/8le8MOECWK3hu9vunR+qatNxijjM9A/a
srlCm9HA7dXI/bIo87R2160RjOIgnVFk6Z/EIRwMSwFkfpiOnTau3n/hZKo5MDZA2mQoTKoHkREa
dn6G2AX1oTm4LSjLaZ1Gj3WGjHyFTnpcbU3UMuuDCOpjwOMK7jd240CWVp8nNr+LudYwoESCfnL2
Uu/dhfDLv/Jnf0yvT/GKypaSSHGeqkDznEm+5d2BzzbuZFEwmnatUddCF7rP6bmSKHrb9PL5L3YL
/XA1ACMjtSamkce0nJyhutpfshIsHpe/ORbmO2V4j8ua7NmHqxEZ/qZyjch5JJ+44GYjEpoGkCCl
IYpr3soyapIzBiLZQ5J0gGWQnwe/YXNuHW7i1I/Z0g7De3RwiVMKP1R8rgSr6MPcs3OCXSYE3SZV
NxzDIlR84ZQ2AX1e6/sWpXvoTxO1j+0oCGWS7mZrlGaehFGOv0QqqyxqkdEF7kT/we6F0MeoGz6e
EbsVk4C08QJwrobQae6CconPu5LDOfkI8446dJcrXhnqaMxtjPC0BSHZDN0amEa6dAUR2tbynAfs
sdOuOnB0ni+50tozBwOydJQWWnTOjPffFDcv8IicIVY7QKtnzHMePXwW/Y1FMqDvwx2lJScQmNyz
47qurq8XRlRxnXRzyHLHJVtACUS4li7JMn5hgI5/iWn/Fddq7AYE2FZSl92RFTeEkIw0ZMpAqm7o
btLL6kDBuBo6Xg2vteONCHlsFUEXZqTcWM4P6aaJFoyXw2GjFbAB8nN+9OUEolzvy9Hi5Qc5ePV1
k6BwbcvE8xQLYPk8iE9UJChW81D8oSo18hSgYHJ8LniDpxs8EKRPxmyxd7Ez+qu934kK5cD6Jo2I
T1ozdgx7awK8zKUWWXAi1s1nXJtHeqIFBjEpek+Fz2swS0zXf4dC45Qfdi0hlOIYQ+yW8VC+0itJ
49DJF7z6VEMvPggHzB+jsdxvyMe02k5PUopTfVUjwC36+4TJ5mkeyMUtpgdxPuN1IE35CDnia5Xy
mXWy26wp7NrBQdZN+gkWDOY98BxZUVRaQVYFnlRTqJN2XQg5ImTBD7KCNZlWFI5bw+ORHsopIMOD
r2BwGldysNjd9NCk/bBAe3ORVywdCP+M67N2IT4yLBsPXD89j+w3WSkYoU5KB29beLwNof6x++2o
zhP9/twX0HHsEdSs/tWWHhpWZdtQyUI81itjDxZEOj6kf0NpWKHjg9Z3J7WifcYeYQOsCsxGUlVt
lj8W37rUa9nJ9o4e7WKpYnjCpxqimQfpk1gQH6Fyr6TDjA1LOGO+5if0n4miaYXot4w1v8pN0BOz
G1LbiEDFi3kqCgwTWTGaMipvtQ65LDwTl8d3dSsaRHm7+hs28WKiL/Qbw6RR4ncsNCpovXVGaVJz
1sPkW560s0W9R47EvLjZuv7VpkmPLcm6rBjWSayKRBtKFcY01i17DGky0VYW5W2eGptHMp6wE/8f
ecL/igCuvB2146FfL5pBI2r98gdPV4F+YSqCn2ddMOBtm1C+58ngDOq0l8OpMElr8AyIi17q8Ddf
CpX4WCr4vjeT6WyCTk2XTrJL96fGz7O3TJ8lIW2iIumz/q3fpCVAEztBhkSDvMI96h7004PUiwpx
mCSjG00b4K/7tGbpuNnQ43FLpQSlvlX+PKIvNjJGNr4WhWXNOV3+JPA6bsUJFrhKQWymfmU7vrPI
o4ZkS0Rhtkgo36dtzlOoflZwV1or0jeULREchi6gF+UlP52op4IMLJjaSupnpiisrRBtUunpe+QX
oTUBMsvq0v5I97KAnaC761v9H8Ng4oqWAAPKf75wTtaWmWmzVfLyfH8WA0MVvbQVC2mPu7V8fEiq
3q9jiNwAHLtJI+wqXTujgCMKlB+G6DXxtXab8Fg/dCTtcESfKHS9vXhSw5X4vBU6FZwCqAVbegvd
67Ra7bQq6S7Wb1xGyEIyLn2khQRvkSOWfl6czYgIKRaoQqAZ+qurCayR8ppdGjPdNTgaX25g3fHO
9Zrbfb7dFWTUsKVPrN28+zbp+eeM4sfkYkWSXB0OKupcOXA8uXExU/3srtc/sfQS2PBEyccONNFL
ONEfkvU1pJbE9bj5DTzc+ErtdO4t4ojuPjD3VUWfh16gH788V+KxfjnUGcbFgnoHEjL49CvT/29R
4MRxK6eJlLcpfAKZJYiETDQWNIV/9DMCy4n8nLLp3mj1KVc4Wfujs/+HgObyaSNmnXDkHeLkUD91
ExszT351FRIitUaeEwHWxJDHoQEYltWABsO5e1vgG6on3DexHTRr0QitpSizWr69XcBzTZfUnTqN
E51ydbiO/EikJrM0qtlxc0KSbJCVJvc9byeoDfVUiONYQ0a350tN5PB3IXnKa4J2J/RPm2cd5/Vb
nsT+8L0wDijWeuGZPE2PYBybeDnGyLJ7XvO+dY8ZIWlXz7TViN2SWSjDBv7GD08oKBo8pcw6jPS5
+VZUeGR/uNGYEg+N6ILmXe1AYhEsq7pLb20wuWJQlSb8xY4iF3tlWw/2I4mCg8gxvhK9L4Wn0Syz
bEvUfom4HYzEUoABk77NtwXtmFIL+hv+svnAAPNAClceL2UhIiwRupBzFGauysmjEtik7iBwoAVY
XR/WFocezBhAS345SI4soAzwywB5jpAqgrOChr71hHcsQTjqeFeoSJQzVb7n7TZuWpuPizvX9Dc6
kFzmVulnvFNC6m7zdV22t9KiRkqffGsVLqDeuN6mrZmEw7oQOQrTIfxRD2RxTCtMjpqt2UKzjKxd
gUCByk3DPT3WRbMsuZIGl4AUIQZ6bXQ5r1y862h0N1Vp0dGB3rE0tKcDKLbLBoqvCciq1MpvKhMS
jralmrEfh9xMsUauVY/yXoO5wr7Bh3pDM4ovpS7T19C5z+ZZcvGG959IXCOjYxOkqgS/cIPxDPO/
xUc9eCnR/VrjMkSVSF82KPh6AB5IfB+OxLJfbDg/g0JmMvQFkpc0wpAGcl6KBlAaTGVH8QtIwe3C
0wuIumnkzyO0hWHuVt+qpgBlobv8CasACvEs6X2eSeE6lW7O21xqXeE1JucAyJqGwBnhrNWQEMes
JvU8fa+xuN7U/ghlIrJLShFIPv1C31CtsgD5/xIvy1oHwX+KOVvvSGzDOUu495B41qeyg8rsRfLu
mR7OTa5JGKpU5FdZMAe+Eb6Vc69EY4uyKhMnmQWVZ/m7RV2BbhMt7JT0CA40B0dr2AW0mzD3/coW
/NlzbEcHUifbRdCXIRcPs/lOuC6ToaG2Nkt9zMCGdzf0uJgrB9WjCVE1qZMOT1Ws99hfpAzdIrSp
OLdbS0yKWuMjFW1fPze+y3DTKG89yTDboHOekrHaRg/jUHWx6/xOai9WwUk30c1yCD/Lpc69LtBh
hAZjFj11ubgrQysg5pQnG96ZkQQIV+jdrdMUXoNwNZKtD45INcHjiT+UDvwceBd+HE2rtEMRwm7H
sMe5J5a5keB7fv+I+u8Gz8TbQ0rPzliH0SVFrqBZxqy0BxS/DniVakhvcWRjsRiA9D1PERHepkzP
9Duz70usymSXVV0ocHZcA7qNkmMg3foZgmmmNolFXbAiqFCzMR+RSMgItbe/aECm+9geYp+3zPT2
sHE0tX4+mMyQHxHUZ+dtkXUJZsef+w5uJKJKMu0r1oEgefx+bnoV1igKvN8p3Z5sVMbc0xvW1iTa
oys+G0I525QiIWKNjJ/nDuuQRE6P/UqA+2e9zYMuZszLAEze+fX/jAKtNQ2Y4n7javkquOKbt4pY
B3XwFwuMHf1Tlc00wa28gRytbLAp1vNLfNBjtO+zzG7qUJ7tljUTy3Q571s+VC8FeRHNklUfX5AH
shod313n23YGlhM6l05YM/XjeGdLsaen0JUeRXdiwmZ8B2f91TI88jBCHm/vf2KmkdOImgm3bPhA
4zTB1jiZbCIKA9aYrytaeqEnB4Qeqs6cQeuv73j1hiJuNUax6d6J3gV+ZFbEn+XuUR9HQTXJkcyi
zABJj2/96IdBiMSCN0+H1eBzaMnGoOHIwVcDF+KJXQ9t8+BfQXewiUMlmEj1mRtjA7o2fdeT4m52
7SyjuW+V5plDmVYZ+TAqChWq0Icxo9kxWSz2mCp5sucBXrTSM3YqXqi/0HejwdrgJWm0eEbJIv/m
33kbb6BH7E5Sl2pb3YjJKPckSSNPINUkw3BgyNDMl52iu3t2va14kjktToWWnv46Y2L0eeIqhseI
BStScelxBg421c1bxde3/kb5TUVjXkOIHGSR1Dh7LacAaj8NAwaFX/YGq4InMpsV4BEkbM4l7DSR
rHgwyvV/28P/rQWXX6jNJEOHm3WEGCdE29Nd1PxNF9n7lpm0qPkDajH52OoJadVYHnjtZmnVTdnr
F8crWrDxOnyz7teG069hXhlbjmIg3vu7MutHNjaXL15JahMAcaSLNEp23qTV8SJXPFfKZt0fqfpp
/sN+pzdEp2c5gw7RdgQecn/gKuHhkQ0f6is3Dhnxy3QRXdX1e8KAxDe/NcRzgd2CHP/M1dBAxk0S
UQA+775BKofIEoWfUU5HYJ6cj0li8GpT4zGwG6unx6SW/3OJOrBdgBhbTtlDq5JztDlCfutR3uWf
qDDPwvtpRIdyoZpSe6DCZuWFU+muuDvAnoFEH+rD51l9Qa1tlQh3HPJcmdLH5UHJrxGCRDl++Z7W
N7NEaCTAYbPc232w22pg2jf4SJEd0ejLSnRG35YQt5QuG+Lpo4YANfJ+5GrInYWm/2b1bqCoRSAj
3EAHp78EnM2rWwpmbW0MERxAFS65L+Z9MltRfzz3OXpDwBCkz7P6vurn4WRr7rfaHKmAk1GFuFPF
6aFXFB2W36ABsqDmCvHuuzPg7XQ6RW3sBuhoKzMrP7EHuYz3abAoYfliRlhljV0R61LGP4YNmWWk
bYn9JM+LljdyDjmPC2B+0m0nW3iHn1FN2B/IjArlWUW2OzlzUTgi5iumMF5s3qm16X/8AbdVEE6I
mkjnFebg/i+ZE9uCFmf6NwdmG+iSecmDrIk3/uE+dqFdqpBvvo5+JCb2vTe4kEjmFidtDCgMKAZf
7o71EgVr50vjq0hN2I00ExEj4LDpTbjhx1MT3sFuRTVNJtECdkfZBHQDcHBeuVTmVpLntjrP8ls+
6iNguJ7rQ+k1OdpkwKGSyLhq5SGWPR4WGjTWjLsyEOvSNsEZcempulKHz0QIS2PVjv4WMh2LabNk
a6GAiZjQuM5T5SbnYJYRrwGxBO33capsiJlTDb+FxtR1t6ATzCz0qKqfSD7E1/NMW6jOzdMDU9Hc
GIXKLfb2kA1Ne9ppJsd7cRONaljAYNa8mtT0Fntj2ryrV6+zYT5mO73YjEPbqR1KB7clAcukkEiN
HP31lfRgbgwuqqHjhsW2H70Q9grQTVqkKBU0GbJeE+dHM+AFQu+z7WyO/Ee0UPJT0was18HYaPdG
LAhXWPrWRx4GnLlCq+ap2AkJsTVkrOkR4d2uPtK1CwtFWGiSCxGWkmDb8OPgUaZ38IJaJbwXFjtV
/6YA0G6E20ZsBJa8QOAhEGdbc2KsC+McITpo9+/4of5ESkFHxpKpYDtAU6YoGgTh40lFtzHiNrw9
R4MLDXnb0oRnC/UxGNwJwSxggBlTpHdnVb8xOgsEHbhZHKRzn0Nl8Z2Fmtb3JwExEDrR9E8gQS9U
nZue1nU5rzcTanJjOrVmaMB57N70yUL50jzKw+9i7eMrcwwwdvqQaj1yp/NMRc2lnK5+jJevxeGb
8tdoCqeMl8Cw01e1/d3J6kEkt5Ryzxyj6lNSAcb5z4V8lfHJQJl6tf1MtZe22ZjMRVg4udKHZfW9
JBvz9KbZaZytbhrdsg4Cg78JQF0wC0Nwny4jVi83RkFJaHGmJf2g4cvgDpcfblAEFpuUJnQaXgUW
aftfQ+kn6hx1o+OdlnYYqq6L8b0zYmyTJIyrVO0IqFEwBzqxTe00gxGgaDSEVcHpnYU4BPrvIGgQ
Jg04cW9akVKYi7TTsbe4A3wjTq1BfpGluQqyj4AWZNoobFXWIanTvv5zGOoIeDT8c7OMKPNweqCy
mvkmd4WjXx+dE0YPWg9W0TbuJ0I1HsFlp6w83t/bGoLGwc+8qINYL55PboMaRgiDML/TOvVh+mGb
+hzFjP/hpAimugoACdeh2vQJ90rVMX1NuesAsFsLxsLsAxGg0HCTHUlQEEswp9EyTwT5inWmSKUy
lH+u0uIL5SWdWcgnDK/rApAcEcZzaYhQjA1q6YEZ2N6/o85/s2NrmXGptcbta2IJ7VBN/fxw0Qni
EDdX+EpoSd5vSMZbqo769j0LMsKjUv+C/GLGLLf+VWEj/d22zpAcX9UoAXnZmR/obma8TF2j+F/p
Olfm7r0uIzalYfYhYA51JjwB0V/j4X9LwhIJIc9CT8MtWEZpHH+5fz9+rq/3wANrZf3U1N36PYpd
kDaGa0XjqmX0p6Qk+oOqoaaglaX25Mg5SdpuWDEoxAM26M4YpMZlYb9SVBTrEhLzLddrf0jgo3wI
paLgscHV2f4sLcU0aO34ZhgRzTviAcVdBMwtPDNaqvAP2OAhyu5pm1VFCdc63SpZ529Ut+xNEkWw
R7dPUx2mJzOcI3zg6nDz24RdVZ94Td1ph0YedUZR/JmqO5Ht1sBiPkSpxFEG9N5FVkYKdAEiUYIG
QzF1nPdlJgrWkqQIGwW8L8iarhripeEbNPFqqqZ43vVBkAfbXS9/MDjp8ze3mIt4RV5i6HiKok6A
PnAJ4kyjXyEZlgnxYKrBvOamS3hjCFJnr1uEoiRCEXY9y8Iy49PIvycvMJnFvY7j+bg4Y39xxs+h
pYdCGf4rT+PpgW45/jyMw2FMLD6NEFHiWGq1ugkIkd+XHobdZsgBzKTHG9bKqOCbROBUEpzrZ+GH
v8AHKuzpObMoRqrDPUtFONpxepyhYkCrlXd1R+QP6noIJjwEBlZFE7wzYmKG//TVMtFrvkLfD2z+
1vXzArKCS5S49i4NRj5wPM1eix0hETWfpkSJnJ3lfcwvPqUlIYaPDPBGMMml+7alJ0cpvufq3Ku4
u0mKQKuuV2Dbce9Pveuvv7JPnCi5PB5CQTC8frhjMyduQ5T7u8QExKo3NDkKMGCnxaIyrFcQIAxb
A/P1Muano98M3iujy1iSSeQmWPFJNmvAvPz/LCkK2G0RcbaTg7qT5hMCOKm5cxJTn/jr+ygV+CCW
pL+tG+/l6LHYA1La9YWupt07SFlhUN5zixceOs9HZXGIznzGw/XeKZn7JBhMeDa5HhyTnJ0ubXn8
WumtbeOAke0aATQiwscBMsQxrRY69dKl8z8grdSRxIFjyu8uuNMj93FPzKLxSy8unb1Q8ukFYoWW
6T9DNHj3z7QlnyViCozYwpJsQX2K2d8lcRc25nUfXxNJ3rKvSoLMl0FlrGiACQ53c/79KvliPXkT
T92QiH5JcWCFBABsCOpbYhlLYYW5qW1t4hn7aoLn5bPmoeXb1ZieLggcCkNleRaQuQpxBiHCbA72
x4PyMC1CTDoqlR/FGJRvGN2WvX3bpGYb+sIcfLMEEyDpnBWdD4UtVPdHtrha2s/n9lMDyJtQ5z1I
iefqeQP2Ojt/zoyvbsSKMZiNiQWuIwmmSsEEQSoqvsokXngWnDhN3htuRZijr7cZoRHE+SBowBJ4
EPeSJVahx2VuCK439grBymaKhhNYCJDVsQm4DHa8+5osK77rrhAxJTu1VA35Zy606wCLaMrLS4Gy
88VbyGaihkW2n02KQUXvdjzE85jgcWpyun4soaxy8dd82laT7f2KE5LtaAuhJ/lA7WHeL1SRXDrg
X7Q4jH1NCGK/fXXymHWcaTLfj9lcZm7CbIK26ahkmBSFLgxm/Wd3XblLAMniGTqaqBiXrIwbqjae
jk0YJ6o3Uz1eHrOhsrP5Cc+cCxr3iCJLtYEGU7YE+pDMDpAQO1v7I6CAsIl4qwCWR6N2naGnKG4N
RXMiTuOVClNZihvy6VZBsCFr27Lbb64IWT2xdQLFBpDIWQfXwFp9Yj5uZl18S0VMEZMUfwnxXzgb
ga6UBWSD+sFVTb8aswulo7KsacqFf3glKepHy5jpIz+64Oq1wea/cb9gdzRRp4SjobaEuD6c+biM
pyef5znosHh4rWyni9Hp0USSjbRWF4HYw/MTnOyLWeScl7M0Is9T+LKfnpdmUnITikHUVkaBZciU
3cFuo44G2nG7Uh/ivNSerFObIKqKi/lJIq5/YhWAm4j9FO6UbMrfXl/pl6zJG5WMs7cDhwsgDsiz
zAK6gduqspBi1f5R5pJjSLz00Ibsnn7OdkScpx3yWDpNreiSg86YbB5roBIzI6buYlqzocs3v9lD
mD/O6kSQ2uFnta3T5my0wsf5Vzq0X7xlq8v27/3x7Gnmcr1zLh7oh0fNBv/q6m6g5Y6fVdJPm81m
9q4oHwbE/+9l+ewRKtKV/K4xdKQ5PqqStKFrP9bCdNHRJ438W7mIA42a6iWeYW5J1OteV8Hkn9lR
Z24n+mI90+RiWv+5ok6PcfBfhqCvJs5A0Q5StlYqubyXEnQ6vET2akHzWqO37O18sHeYu/tCJ+6b
apyOR0RlzqChDUqS30qcE/s5shYow7t9B+cf7g0ivw0qdznjW+HBYQGpiXRoXhrBnz9k/oH3ZWdm
ZENznKLLjlsy2OeaI9LBWnARadBOUgMz5if+43XQIVfeipzDZCMQS0GJfHpZDK5tLjjvJh9qDi+4
6WftJqRS9eNcLBCBPJfl8J3/Cxp4yGOdV26RCxWfglFRlmvoeT4NtmdPodYzGF2ZnnB3kYfbWmWU
r4n8Oq8baNF7BZoP2FHZ/8Xy9TQe9o4u5t0wbFNc9bZ/KG9ebDt7n2na2AbC/GQYz/V9VTRXTwJi
P207pNxN9kvBV3oL7R6Woa3NWC/31dt5gcByCK/kWrbO+gpaDlrhrnjpuNLJtvINwQXuSE6ZYRVd
1Efonf+0IWKOUwX+XpQQKYGLFXsy1cY7UdXvxMfuA7hsEe70nCnWTWoKR3xuHaRc6Ah75ToFv3Jk
n50dGlMvngv5t6szWSd875tSlVpkKYLzchdFKwROIqD2Usp+f7A6MCsYa57uR+uLEYEMcrKGA04C
D0hK1oU1aOxm6WbsvjeP2Ro9Q+afaoY2hHrTPR28yhHIFm6TbKNi7jJ/sfdMS/sMycJ3ZJbfC+l/
jjiYJGRd0DSGH+uiMcbCJW4K7FwePYSDnt4hS8BLm1FT+2ClO83ZviPoZ6Pq2g48fmF5HfgTterY
9O19tZJnYgbxXLDiUuDMwwaI/GDE7UrHcCBf8fhw8HyW4LG8sbJlDQnCp4s1uO2bmlUS2S4K48jk
lUtRnBUaJmb3W+rShTzU3lz1DyC5jQyi0mnoza9fCq9+KKqqWIez3RHU5h8aTuBqdAPk/PGMYpP9
8uNXZijQFN0qHGrsPNoVtVW1yimmG7oMcc+nDzJI7NvGkgTzZi4yy7WRNYdOR0Ljy4yRRO88dT98
67USdMEOhiw4Whn5XJtpv1lu9ySdEK/pujvjC2QVnuP6NCqCiDO0+ZGMdlQ1LiwCAFpJW2ykzWJs
W0JaXZIZCf+V2PK8HP0C5WTfD1C9u2lk+29vn/bNMMPDMXv+Xc9ANvy8sam3AJlUEw++kPdRAFyY
yO1ZQ1/a1g4rFkoZTSJet6yhpCq4bimUNKPIFRlwr04RWBsNcggbDAwGScGvtATZx337IrhUUEPz
zZNdXR3zAbF9D14ukgj/YPmf5xpc0OZXCfFYXEJGOefELlf/Ea9zM0CzobYnHJKacgY2e52KqBpv
2Ex9mthrvdu5rG4RQBGdPIBRBjjV55wqYO5DVT5UQfgl3KHkxq8jcTaBnpwNw8zRkDT7VPeDK9wa
PtcRyLH/o8kf8lofhqVdPeslL9nw7z9CpoUMOnFsIm85prlr1vN4LDDuSl0Wu+Z575s/cUycjZaW
wz9Q9dJsEgayZQ1kkL060FCuftHOX2ysunMxTZ3llvSpmcBkANhp4jS6JnmiYY3d2eJNsnhPwey7
Jy4x4gNHH9eidgkspZ8EN11c7HMA3768W4/s+XJ/HfdZbjMLPEftkcZ0LMv+QYudVKOUEmjCeMui
iyqdYl8fs8UwfgjQqS4TpSFtyx7sujq8a9OYYMXeqV9U5+aJeXHJKTauR4h+BC/k6vTt8+qwkWyy
8W/4bF311DriO8bIjZFzukZ1eEhSU2OOe3ObAkpS8JK5j/rSwfSRAUxu5Am6VRDGwIRMXLOw/AVr
ZXnb3JFUqMPGPd3GdP5eZ8Z9c/3rhjkjzEcCJRbv0cLuTM9Vp3Is2IoPZTy059lOSTGEROGjVk8C
yz4NgqdVHTKBMLtzj1owhGOa70aNT0Ir/3QY8wp2WFL8OXmnWiQN70DWET8ciuxOX5iar2iiSvBV
9UZRD0JiI9M1wUjXIEUlzlmZCsFDiG3IsUoBRx6xWkz1ArpPPaUH4oesDfIZ5EMe/fa4PaBecvB3
5ba9Yg7Fy1HL9z+6jd7GRpUFCUzB6+Ul5Uqp8HvRSK2XgOgXE03nNjShvBdN7dS7ge4NrdGqNDH/
F2up+6hG+ipu7duOtt7gNhLrebct6WKbKXQo/nWI0I32rTmsCkNz3bO+EB8VYpOmtGFIFo6TmGXI
ZkDnuXiVosN8hb0gSW/bNh5KVw/rWwWuuPJ4LHeZzbcelT3EJQjnGT4fx1aldD14Qg1xjgLkaQA7
HBlVeMgmah+J269QRxGVEopXZmlVqlF7FHofQDPjtW8peTDxhuLBkYVpFcMle4h5NsKvieHHNxxL
RynVKB2Sym4VvA8b9AYEVGmozcODKimnRj6vVu1H/3tgdt+hdZ8Cj8/TTsUqASvL2sF4Ghe0oLiz
DWxSFylm3odrdPOGYBNix0WXzF9uIf3h6CUvtwogKuyXhwparl/dNDIQaALPgtaQT4aQI9a7Sxn2
bCWb7yo+LoeoQ1oIBTJlkgqiniRLNFpaJ+/12/XvyU2FtlestUQscxUgATh9QyZ11q7YRjNPp8jX
g7c4vszb2bN9lB0jnWG6A9oGIWYHly59are2BsP5mKD5T+aVS2vGTW0uZJYx4GmwpUX4FTX7y300
D+jO3eUO9uoknAFM1/94mwEItkfTRrbm3u9Wo1RryYp7RQ9VhPgYTygJ/zmMBZn8ObcaP27jwiLg
M4DPRk6ndzaz94reiR8oJr7IgyOe0q8MiocKmPOSjGpinfXTqSR2SKTQ0IYXiyFzaZu/D6j7onDA
hqDG8ToGz/TswqTUn/6evQoOvApydA92qmdpdNrqvhQOhCdHqFYyB5oHDk3KsJQsK20l7nLv1FOG
m+pOBin4nCmprEHDtKVIe/NrkIkMEr8hUSTNhOodGyDc1YY5faAKVBK4p8XQDqoJ62/v9Egu8kka
u1xzW6WvojSQ/xnFJAZdd7L5zqIvzI5+XZ3yGUZAghSum5qBrWkVGIsYndni+OJ+43NhzlmdUv09
Mh98gKZKY8KjooH+OnkmgqDJ30rCoo/wwuHHnTqs5LO79mMBJGRGWPS0rbbrVuZU7SJxLwC6gdYa
j7i/A4yqpyk9YKjtnaerPTMVN6Uq82WNYxcAWdTE4C7ThQxFmIi+JZ+iD9ePLRb1EL25omgLHmmV
VWMpe2ykmthCuf5JL7udp8RVAvY/toId/HszNwhrz+iLcVR1lD02Pyq58Z/y10mek5eF45CArZOB
ZTXKbudbz6GhH6Fkn/OU1F7456ivtsPXYPFv5+GIZs4pW8Iv7VKtR+B/M5ULJOshq1TiVkIkV1fW
bQ9FLzmLLQ1MEvhoYmCcZ1kbpWaefxF3jVChrjKrEegM6TUZ2y/0BJ8uRJidqw/OBqFmvYPGi3f6
acm06YMZX5D2r+ixczWGNolmDmN1KpsmSN1V89KS7Zjk7D9Fmpl5DlBgT5eJlxNYU/ZaSw6xOVLk
gNyk9GiVRqzHEWPMg8saQz/j5RnjTt6SJRkzwBr0WWS748DojufuAXGgafIXgrtAdYSZ5GRelolX
fAhFM13i9NfVSfm1bSivLKTNRAX5szeY5OylbzP9et68KpEmD6e/WammDkhk2nGw0VAZpTjgHSY5
/m5UUn2MwKjmElhPMAssbsVid1nmS2MdjoJaIN9LWkN/16F9gE5NFnhcdGz4VpGyhfK7+hLzmJ6M
tPOEVNdAD624fLhYDJCZxHESEZCOSU8uks9yWNLe6KVBrY7pUc2hJ/Odsh7K45TVoahwVMSh7Q7V
sqSwBQYZTXDXzdxk6dWnlKEFPBKUlYiXN45DjADDhfQPfpnEbLytqtigzo7KYe8W5EM9x+mpWNy9
cvSdurArEkn1zbydse58H0OCakdKiNHhMsSIh7FR6Z4Zamgza8XIiLkhJSMG9eYgYXaKcSq7lIyV
Sk9Zg3uh4Z/nE8EjTPVYMRLDDitee+ZLHVgcU1Rywp0fhmgSpPhAMCqdBz8KfEHtPtx0RB+GUnpo
ThDe5iwIHwt41yfvcm3AroYyEpHnPYk1aNn4i7lZEZxlIrCsT8WWCCHrgmq6NLj4n6RLQZ15UvYs
ClcZudv644uF/HDXX2jAA379MPFZvfmGoSBX8E4RpG4bcnG8Ah/G/lfKyvAb7toAyThoZf08xNCu
L2vFEvU8R+Ue/A0mkXSudKdijahy/w4K7JtYJ9/QWxbT+hQVCywjWIZcGEM+7N6nfF8Lr63U98Sg
fL8/VR9w9X7fQZyYQ2HZjUyB/DxrZeSBmFG/DJaJo8JhTqE9F4/i5C9VyYHJCsxOHYLT1eDixt9s
kBTkENYcBM4Qy1aWk+vLhepzdjFsSkGhxGLRWphofuN5WJzfDUI6DP9rKZaA5w6lBhIIUlBe1Nhz
AHsRdoyQbdkywv5X1pw6/pN7Rm7phdRgtIWO7sCltEbCIDmdSHH9LA7DbPgN/SWET8Cz9SDY1O++
LrOe+0bNcmVDnGPZ7bvE7qYerVKyTwJkvlVOSQmq2UE7gY8FAz2qub4KyxqYe4GGRtxQWi9P0whi
Qy27GJNDz1Wl+K/GFxMtenx0dipzRv/dlBnN5w1vLMuTftax38glXa+9N9YoD0vDQ9iTL24VNwo+
I6uETb9kfcM27gIxMkJVlrW60B3mtGbRlvWh0iFBFGh/r3PJNBOgtAzKHDPyJbrDdGMHiMrE2sqS
0K54iP2NDY0gP7sjR1ROXGIuooEDc9alzjltUAAGs/Cb/R9Z+PBXKrxRDcXfKZsSIUv6CnIdtIs1
LYsy2rasJ3fPyMXSFyV/EA2puJMXaJSd3j2g6wF4pVsihwra9G5+/WD/c08SA0vJt8h9YUAc1Ibg
rN/sxw+vIHaY8soEVOfijbN8y7C7nz3CePNm5LXpzNwtn3ElEnCeb627zw6uqE/YylvMQFOzgUqw
WAYalOJ7sq2pab7N5T56szpGCgSMdnSEb5dEiSZhMgtCakv1aoJSZTc4d6gQw4KcHP9KqP9vE8Mz
Z10wLYjPc0tIRFOn26ccEyBFGH/c3Jrf3p9VdhFl4NZdHoSjykz+mKeYWSRhFnWcGyade3hzAiyJ
SY0Im6CoWp7QCCA7nTuwutcMwSQLa6Nvup7kbLxjppcPJzngl6UjmFp7fHMVLh7bYfOZqfyo5Eah
b+Kf8qPNiqM2Gt98QqzWGLwerLCyJWedBAcPYN4xNMXCrJevW5O023r9xW+HPyBoGRoy4xHVl24d
4A9qiMXw3l/FuvRbi6+eabfMLgW9vYumATKmLtLy05DPfs/rqFbAozMdF2oXYO2Qc0P7dMdu/LmB
lZIhHt+/v1qtIvs/8ET1HkLwqDLjISdaW4iXSrAwP5QuAA4137w2ETBiCiV5u7SJHKwvS2U3tO8j
oQ1MOePZg62SGqFJ9f/irUEslJ3QRg89ICSlBs0H/RQDRrpJSKySJLPtwX8Ah7cLEN7Caz57Xez5
e9V3o7H+sH6s0xOm79dSwl6zjEvcdT3OtRs1rx8ckaMu7sk1Wj6dcNFAZ1B/F0uupmZ4nmgn1hOo
bwbkvi9onhqtNu9nDLDqkoE72s4Eju4wXme6loZoOnsbF+GDMmyO48X1UfS72+ht2UdzI1Bci3gx
E6qX6z3IzIZfgH7EVC2oVgKnBZDwbZv8WBCGqp13x+2htltwrkFaRKIZWGu9QRPhTxwITi+aC82C
8nPg5Alg2kyPvf1DkhVycn4RBu/eNZnNtd25bB/c0nc9ElGzMRyl/qtccD1msCHxy37S59owi54u
6irj878FXM9ucfjrejCVYBsLN4lZjD3F4HdKkSJRQTRfDjINzWgKphpFq66iJ29LKR8wtggBbvby
ybGq80l20K1N6VStop2PMjiusrEsw4MlrHbLeqe5Tiksc3qBNKrRLmBdqUkq3nzJD+3ipw2c1PLJ
3wHl1IA/ejg7xtzx4rLocJ9kRwbAlfkFFn7K0pWO7EhqsMLoHpjbnPxvq/D/q5JBN0ZC4kqlZaa3
Gv0FNj5urjbpn+DF5b9GLdoEQK5aWnc3Xs+o2UoJhSEtIQ0y4SJzAIKJKVROf7ELhDI0iTS/lU9d
iTRju6sC50+knCTV+RnsU1B0Em5Vd82LEW/72+/fM3a6TZK5KxKQEt/S3tyfUS+GOXsmr6gg0ZGU
V1iTh5U87v4SZ8z/RccX38NVoB2Ku1Bpl9XLmXjqXa8xRNrBV2rpnqanWvLRGbyb6yMZkYHIKK0T
7uNjZa4UBff3eVKPqBDfHNoiLzPjw0wxeqWEZykDHOTjGC3F65DNxLsIgTh/DFpny3excPCwLrwT
4ZS4UJYOdbR1BdKYKEhWw9Xn4pDf3ysbbZiWuFJQj2pqvGU79Dt8c9PKjACHRUsz5mYpDj014oIF
QKeUyxiGNg4E1LKWqKdAySKXVO7P2PItiSu/HNpP/wFcFtEvOCY0GhGTMWjq1jx2VHZbFDMLuX92
cvs31QNH1qravarJn3KIb53maPRvAA7VNANvacW+Py01eMLk+5/Cz8e9trmmtmJyoMfru20egYmP
Ahye0W/hezc/cbut9F/UFkshaLJV9VTETluPNbopPGHSPuQyWeUORPWQ4upkoMOQ6iktVIgFV8dl
fMKr5Op+x+DDQcPALdJ//ZJYEkYFBmSeFq0y2eGa+xRODhyy1UrKgld1xjIB50Yin+E2HNeogFEK
Qra902dcQfnjd1eN1Qh+W6a5g2PcY0ZTdAHQUw1nsLY1u/K9J16yovfQwbPx15pjbVfd66c/gYUb
Q7Lw40ZdmhMrKrcKrZMhILAIGkKIkqKJHV4smO/em3hX2/4Bwl5txhK8T7/12H/I5T9e+RTwdI1s
Nc+3rKqd7pK5P0LTSYTHbNESptP+vit64fdDmAdBJ0oW8go8ccZoFyktDuLJA98adbAMV+WQJx/M
2VxelJt7qHyPYdVqoFBerNDLIH/FUnRMmW2/l1bqOI3ltsMjPk1DQ/7pubfbjp1Um8amKg0kHkIA
tfTxY5h6RvIdBcm3q16a9itgDdNv4YYN4n2Kh3vw4hZLqhspHUnGpkhd27/wexBecDJsKC/Q8K0f
oh1qDlnvfC0Udst6lKzfDNT/QtEM5y90UERpPfWjrB5RS4PgBHfhCuCFJKcdXLp63CwFyIEybyz8
t1uL9YZjC21gFyQ9CXcIATHp7H5J/vSXGShfqoa9UxtmitJx6OSaBNHP3M4AJHVinWUtarjr0Y9G
9IptRmkwhDYGX3QJwOx+j7/RQvX3ybEBkKH5jh1GIF7z5hmMT9xa1bWZi5BoUQL4YkNLLLcZft/N
9+qGs8bZ2MYHU6EhDdOr9q49EJRvcGnxomQgMTplbqsNRZlEAMZCMhyEcD1K9jVvTadBfvfaiDgn
EPoEqRK+Fjfo/QGrBKv5VifPCR8gJIEbLHxnnnvvlDR1epqnaOgTO7VkbVTRramp+TeR/kN2EKoB
S/DWYrHksbnlXEAXnfoV8AjJOMLCoGUKtuXi+8brJ2X5b7Ie7X9mwGw8ydgyjlwMu56vg0nfWf5a
788E0XIpy5bt6lGVW4P4TbCBdr7/TvN41sJkwpWc6hiZR20YmTftXTKbYBn8yhVoOM/6ij2Zz2v1
+J8mZ7XKmb50ZcnQXZPOsIJMzjjCV1kubiww10vDj7XJl7fiaq8VUk6cI/OLopsezpVw8DaS0mux
B0zLTIbkEFlOdQUg/eD7FBFTEkps67D0BHRXmZwsS+zL19ebl8GGrvxWbup70V6oma0V45cK7mBq
on9mvTZPXOIRbpydWbJJYeeyXrgclrUrzXbZHZfA/o74nTNDZCkA1D7uIyJeiYc7pTaVhkZaNZ9P
QerWMpuGTNMZ+qGHsD4PMgnfok8vH9FGZI/F7gFEeojQOd62jKg3b0Zel2rXRzbCseMsbVL7uoF8
jRH6wCpCdKEpFltbAOCWUITVomM8bc90N4YDL+O9EA1FGMc029mzPG1pdHEgpgqJXJp4a6KvROs+
Lcpy0wJh/AujfPKpTGo9/I8VcYQt6EnyULyZmW+/U8+6PROyCkGzfRMOjbqrCTnzHCkfWf07fIRD
CqyuBnuXLvfjSlhyLXywkG/ODwLO7CUrkcWgaxkON6Dbu6f2SdczVfYKmKZw8Gj9ySz2aKxztsI7
9DcLadFXrrmVKyWVEjBetDYlW1/POWv8eimeSs2/uk+U4wOdliEwCVRF9OK03Uot38gttltahbLG
XyHiZjTEd+IIeCoeabvc+dtPWlV+eWT+bgkAOGrHVbvKnjyWTYSTtzzBq5D9aXk7t7XtvbMzI3Nt
IfKiV5wnrvQTKlPD5cQK5P++KIPC9MNsgqr5aX2aEifi7ZmDYGALBweBv2UySF2UGzw4awnO2IXd
jPpb1TEQsNK+aMcyZUDph+42Nhl/SamhTqThePhpPwCtra8rNiEiEOVi4ers30HR+9vTJc16TNwA
QTu5+Hg2Y/+JVCiWqwfnVc0kvdKPKuvEumNjtQpK7RFYTgMMH/fQ3oGW8GsVH4u0pUd3dNdrrGud
W3VXFmvTuNT5c8HwtgAieaSL2Vx1UnnXRwOIGGFLOB78wgKn8RuGy1KIq0WeYWC/HKwFac3tVpcS
MMFF6AIUWizkMwSFHiXyqO0HVgPsIIRTTlgJ4r36IF6uu2XXJFY8sMZEuUKKmhqeg6f7d4yv0fVD
9t/PxcJfafxiDUGoSNXBhwuRUajVtCVeZKh1tEPh9E+FTdNQG+fiYWlbpk7D1SUH8k/vFANFm28g
fxqsbhVHfVCbyty6hn8eMaRFXGzCLModyvWu8s4mz8tl9NGhnr6KteHrPyvk39XNGefDS7usB+Zg
y/ol5/LBLheLadV4GFgVO5KbgRKDBRIHkDARM9Hi9We8uedHl6NXnT7HS94J/P+J2VfYcIHp086v
ffZ+ebh55+Ncz2kx1eu4XJk7OuNFvilObQ8cfnShJEuDhDxJJjkOJlAEn3z9OIXR6t8fpndUJyV9
oU1BcnCx6wqYUGF6f/UZ8Snin+H5YcNjEZk4oS3aybs4ZYkEkexBeId3Wp4ytz3DvYQR4P6Nu9zG
Y2srUWJy+MuIwdXAqbyYvGsOdixP7+qaK1O4XS4DQnN+YYPS4hAFBkX3IaadPdscomtPgbgtI5in
uNcVJ2n7QkkTeunNqi9LA0GS9du3RDRIZcpsG/C6J1G0o99ArbYC5X9k76EG7CcHTQX0jqerX3i+
OqEiKvnaAZSFbYNhh/zheW8rcucoo327MeiiZdIqFnici+iJPCl4VwVCjhhYWLlee+VbKH1qkeVL
beApNS335i3+ZIgRAZVMfbqhNYAUPbBegaPKBP4fPsUZooI5S1C6LKdRwN0xwT/lsv2dQQG1nsuW
vC8uh1PRCbYli3kK4dEH8yYJY3h19vhajU3M6WJyeWu5EeJekSM4dQIrBAtTFmgRwSMEhfCGsOgL
mV82+bGXiIY++Ls8vKMiN0HXN/7DdEcwJBozPr2IqPL0Lc2GT3nl2nd/QeTpcbHuzFp73cTQOTAi
fC0JRsmb41tSvv2vIlxFLM3+QeZcJTaKkakkrzqi/JHivbPtEawlcNHrflT/OF0MENqs/d3SPM1D
qdIDH1rHBZn6Z2haaRWlTNs7/jSvzKYWr3YtHMt4GlUzpkNTL1TmiBPk5RJmrmnQVTz/889Uh8dc
djFeh/DsCxZ6k2UHTOwOuD1DcIBsi/lGrEM3IYyXMfIqHFrLo3PYCLbwfP9/8e4g6NvYUoJpAILt
MMZFppRQB1Q42cOmcOnqvQWtwF3zZBwHyYW9T8NgQoUYnj6HG1rm5hAX/ThcTwMRQ4yhrQvNbvq4
FnmGKWP6lrWqQ6+FW/22/wQWk3ytSnF1BFgjb7/PZ3zDaoGCApZOGswx4KKVTfAIzRXWV/Lq3fxc
dz2Z21kca8U2YWjY3/hnZE+mozzN4dum7QEgMv/SgAN7I3XNeGxOLvfHTJRN4mh0vYqNePCn8Y58
b1teXOjWpHcvl6833mUcT6Pc6SeFjK5ZGnhLSmP+e4pxTCwPU13kvsSyPb2w9WKn+CknbQ4tPRXz
suhUyJnq0ywTgCthhDZvylq2h2LheJ37nujfNlTf2fCqSJOLAVMabDmUKRC/goWtDAyZbGYpmJFN
v6uRsq/qDZdtQPs/QRNOOLCvOBfqTII1h24sKGWtPElalzPSgZVxeJQM6UXjtOXwJsnwSgfOHDv5
QV428By9BatAWyaSqKlwMWuG+3MKSiZ3UCaGNWH43XxoSFYX8R2XahvPFCxamI+yFLF2MlKFal+j
Gxa8r0hVn0M4LUPEb32i4lSxor4n42VPU7y3dsXOdjJzIcEnjh4OaYf72oWA9m19pdbtaUf6LRm2
18b1+x0wJsIhP+GXVkLHw4DGpxZpadXy+4J99FebcoHWgOf+p44QINHNjHzIt7sD9EuBGm8CptSX
EpYBDCa5CBXSM05nxkznulTULQC3SavkX+sac4inCZ4Bk140Tzkeuq7goRMdzyo0VuaTxhFa1nRt
D45fggX8FxdSBzpujPKabtymXkLbeT0Qn1vn/FeMb59OpksdN7O7thwEVmCwHt/6zh9smnVw40Cx
NkAwNBgc1zbTbuS0DIWRblD28TJHgjvyhgX542ne56R6lGqz4BZb4Xdrb2OVDPMvjmIiSn9Zx8Ct
4pnYktvlJY1kcDzO9mTfhkYW9PMdkT6hgCbRpEYx7Id1a7ShWItTlf9aoJxWliVOanW3qDqJ4InY
lf8DL2PoF1s8HhE3t4ZcskqMW3buogUneBLhREfYncuy5vUQ0hIM7aLqG/Fav69+G00418ky1hQL
WHxeNY/0w+pZZuYdJnLHFE0fyAymeHpCJooi/JNt+r62Fm17v/rxwlhR628bGUJexoXyW2ToIPiN
6qnxeH77m9zpysGFgh3RTseB9f6Gbb0go+ICyfw/MUksEq+SEt+ezmHkQa9ZTBqFiSIUcVdP98EF
QUG843MRLd0H5XjRG643cZ9txzJssdUTCJevd5eMmtPXx/0Wi6Fox5elYbpg4sCOLQ+NHxyNw9U+
Z6AV3FJeHpBrqc1AdXY3DkTLC5tSqb5LwKIxyg1+fXl+1zs4dQdSwqWwogjhTkL/sjAs0rBTvn0T
4fyxTKNSsvtvn61xNM4XDOEJTiB9hOHpuQ/VJ2AzCfa3Ms+llDzniZ7m+/rZRYjWZPiUZzUBenyo
pcMaECkLK/4W7KH7ujYfzJURgH8kRRVc4W8HHtcAyP244MpuduzeI0do09Z0MpTNU/9AubDuKPEs
/k0I/0SPXDqTA16RbGQpzAOaSQGcn0ocM4/j6OEE1wG5iqb4bpxKapaVL3I9pmJ+lFPysXRHk6q3
5LRjAvfVkzw/QDpMVlRt68uQ2e8RHD0cTTGNKMIldj7kbTHrLrN9pFLUHY7uhF5ng1v+XyNhdEOY
aZcI80PAER16uS50jBJ1S07Puqfrc1Wlk9QCH23EL/GLL1LJ0Ojqn5cqnlVMkpSwtBQZIYImpsDq
xHy6a6n8XGinXt5Hlc96Mwvz57gHaJaF87dhmDQQRuSBFLbhXkI563uplFgHrNytE/XW8fwa3ekF
seEskdbiN6TL68I8E0jhKjufEq94IwE7VZXfS037afYMZ19Knpvg0nzLq4Y2rthiTBFBZqosHBEm
ZtAAI2BTvkIBOIPzYnfav6AqO8KMZCywBjjiOkjm3EhNwjGpNN8SxjGkhJcGT4hC+iAIm6Hz7b1X
lobeNzWxOaJILQ0UTLSZxubzUHhJM4DKiVH+iEKOKXMHzxqFm3AAPwMqNtAXZe2lBqg7+P/8bCr5
Y81Yj0/YHLvquWUFVxO+1175xRG112AyT6vN1kyw2m9d5V7PC7+fJ6wmATu34HbMbgD5LhI/oNyg
6keCtCmWWNjpkErsk+DgAp6jnW1dZS+VuSqCdazewy/NVYmq+iQ5CM3asPk/ZdexQQX4kf3NCLY2
pSvXgSDoKwtug0D9l3l10myhqt2cc7Ioh6hJzvtXonx1v3gEZ25LADYkzyud70DH6w8+MEUabGfk
CLubOTvdJnuxEgnpwZ5zvZuUW5JY0jj7lVJwy22NNLx4i4Kpf9wU63GKunuTcG3qI39AUrwVlG6/
ozCv0EPsed6KxjieMQ2N3MLHSCsQ98772RLs+Qc/3NOaUF8Rm8bsUx0BokvClEjaoFz2l6E2888N
vvaExhPi2r3qEMycLskJ/eXqDMLleR/42x/QJy91IR85swt/+iXQ+Lz90WA5JIyMzGvF/SE5pK9K
60506oghtaT30Cuzhv3Qe+9bDV7AfiBAtgnkBNyQIsmXw4zD2IfTx4FpALSOmMGH/WUhBtwF7p0H
mcRihf4zCYExlke7ZBFiHWc+FtIiJMubx3G8po/bQFNdVnbJySDby49Khqy5bUaPJKNP3GdgZU7l
7Fo1Z9H9IujALvxsOcp+i74GajLOsE+/9sE1cE0EmvL+RdkT2th8ilUG3AkyaLIf9lsh4EpMjBuk
OXhWtiS+0Pgw/6kohDaNCajfWebSnV6Rql3KnyhuvQ6KZoPtIiKwdwG9aqzjTGV/yNogEVZ8GYJZ
ykojMptko4eyE2PnLgjlL9Th4/uvbFDHoHlv+ZOCzv6daA7F3AmEBO2hCy/PRx6O4Rh4e4tbcS4Q
op0BOJXcoESWFW0im+Dx/oq6xFeH+TejVnRcyFH6GgPI+oZ2Z4cWgL75WDkFbgJSFVN9ngyguXI1
I4l0pgtZGJ9qvwFhHHkpcBFR1RJnKzaOy8o2Ql7IGt03u2RhHuh/zk95HPjbAghKcLRM1itO9AYE
/ZVDn7q7Wspoh1T0bzvcJwxuVMS4QZ4sMokEpcI9VDIhuTv4ax5c0udnUuwI1GvArpRUD1direhA
7e6FN4A7kgQasxTeTDPLQyPm5etc/rmm0hcaCJzGyz1x2UjtAawIpRk5Vf+T/O/gYnn5dNiN4+hW
ipziE7qtKfS8nabGnay3ceua5V8STQj+EQoVa4lB7GBixp4n/MkeszvQegG+ERxMNrW9+r0IYC0l
S0R3ySZWDJZNlvgoZaFWEDEFWUORfMBiexdHV8yGWJiDG+8eZbIhgV6c6W2d75k2JgF6BmeK8g4J
5V0U46TNqNVFN4ZksMTR3mTdWpjOdIX5sPSoAxsJaewB+2hF087tQZL6qGXVzYTcNuUSEGKaIpCG
3ydBSsB9qgZ5ENvcPItfhwD3BM758vvek3XH3aYjhTThN9OgwPLxPkt1b5pPV5cGrd9gt06Pp23T
IWRBLMkFjm2CrcgC+lqlrForFGh0NYFfq0n8yXlz5jtZCXkeUvPXODvMG6MU1M+GySdMt7GF/UJt
Z8k+Dw2s3y5ZvZvDDiEJMqJlfYiH617T/KBHtygs9on6UWxQAlPSMAsJCu10UIRGl2HH/YHM0VU8
nWoY+xdEXpEGr9awTTUT8R9oB0AbNnH94VKnKfK5PUp3gASDpVNo12aUoSit9AYQIlFwXIGTJ9GM
dp0gNDfFli77eW53fMJrltWRznkCC/rqV3FeiCmi1l6FAZ2Ks13n5lwO4W6Eo+ebDcdjitQxgU9/
vSAPbAv6eQUJnvdhtQ4GRk90waEHwN19K3zFjXwa7neUcyOPI9BjZk5IgrJ3tQT7ICBIoZ21RaQU
CgIUG5rVYwzhOqR8Pj/PJ8Wt1jNp2BaPuXwvRbACJKvxTWEdU8yciZWkQRys1XAqjxZu5FLpbEbP
V2oq9yxgbXQVLFb9RbVT6vhluCLVAqN8iUqGFYY8B3ymom3CvatT3Q6Yj39xPg/KzwpIPxY5Er4m
gx53UBAO98ExJzVTeI8gxN16yXalNCLx4NUclB/x8MOqX5VNqrTFLRG9PPg3SxpQlPHDMUDv2Et2
N26T2qrp7xTgVPCOszph6oPTU46eHUq8JEjptzCSH4I9IXzBBRG25bz6NEnkNO7wKi8hRE3cUN3R
PQcH3LQf6d/fU7vX0LSd4KaBoTChQHSn9SHzNog65EhkT+RTHxgJ7DcGuxJXpAEVzee4tzyy14JC
nNtKyg26Ld52QoQxFkoCmuf+jvPAMTuGCynkHMQ29VwBSLhfYA1Y9kX7RLX0tPvRbvC4wYoF/tzr
3ub7CObO1depMKIMzC8DiD66ZQUOjuC2rnQ0FZ/3suTP5NT0kDOAmW+cSxeDt9Tk+aQWF1cA0q5o
NOBR7FXDAb7yqfHDavSD3g73djj6anrxPGq+psWgIoTzYxUBpHiwovZZIVG0TXV0fY2gAujFKzBg
V1sGBZO515rwsi7ggk6mllEPWVPpUwIr/eIT5GHmjrXpw/1Cz6ijnOOuvaa04UhyyQusQkwDlDhv
SzS9XI+SLXJ4GYkyKVPQ5g3EVLDZYgCuDm+EfZbvPCKKRV1dJ6CzrNbSi5M+RUymRbFERUSm/Fj/
MbEALeYU3zOJHLYHeF3dTFksOweyy1+lsWxiKmmE/JoxHEU68eGGQ3har2SXyx7Is/A73KIA5k/V
3kDlLHyJ5Qy7zK190GsYz5Yx2pnebujs6Pnwjh2F+xwCRMIcppr7a1SZFMWr3BuXjed9ptIPHTDr
LPIDxfKQveKYqyR9bTsXNMLYyMC/Y79ExQ6rElcZoyFC9SKptJLuk8DzcsJMVyinW/DgMZ+8axkr
U6OvZb7SMZAoKrklJOP2D6v4QIy4vDMQb4NuzRZOUPK1RICJx/AYNAqybLH0szVYmw0agv1+gS7t
8EkCEjQ4usHY7JVofe3NquVbXt2i57LoYbL3ZjoS2QUAEivta/8TwA3i3pifUdsZOJk2K8nQ16vf
htwDhUL/H4xWqOed1YNjDUSq0L/V8D7tSx5IYOCPxxfg6jtv7aTmC+ZzkfuPR9ejqClxQDgCJvTu
uJEVMeUPz8uw+sGli7I33xDY5e1E4IY9u+vxj1UNmhdX0yJF9gQkx8JNh5Z25Rb90jml7YZK8atW
6EwtCJ6DdKr8ye7clQ3tQRAfYQDcQCQLUrLPF6d1a/LWlEEWZGohvo89KhMMs4OhLOAno8va7jNW
pxY2/PPo/1jW8rhUmydCEbWlqEiPgoDyUJs0qQpVoqnmlvu3WRSLezcJAd1CwBPgzJW89feqW14N
R4HEJ+aPBLaCcUPI08kVoUNqw9SsFnCAmddrSUjKru2lxryZ54/S2KnGJzliB7l6DwRaoCLtA3QU
K0LUKMsSQfNLoQ94GZ6Q9RSg4FNqKHuu6uit5goaDJlyS3a+ECHI6AoGuCOzwjeawRHzaye/PA3T
nHevj0KR3U8pqPdAETYQsC232XhawjfJZ3Bc9a4aJC3bMEY6744vOGqrkA2Oj8YdTwRCwTDVPbMB
SvCNvD+2N3pY/H9TYcpsmPxvb4yKhNxfLiGpJJs5nlljW+PVoRGJ44+g0lFdaYOz4Q82phwxDFsg
vuYRZ3nXmeCFVO9Y6Ch3k+faSVt5HiLNbljcZP38qKk2GpWBtFBe0YpCTrecNFi09ssX7eRd9O9N
iA+nqd/7OOE0ZVRXkWVDDXwTus1QlHCoImW27bOW98B6HzLo9Y5YJu0BV4PHxkSTkFLLRgrVgctk
pEWu8MFIP/GSE4i30+0SvB07UwJNm6+H2fO/OacxtPisTzyTiRvGxtVZtx+oPH+l/HBZalKsPLll
kWtorn9I+bvnn6wXOzC08kYCjcFVPixUtSHU5SaoB3dPESUvdLyJupqdwMhUyNn6EexBU8HxWVc1
LaGcSVSs97mnP7Kp6Tke+6aG63STdH7Ld1PqY1+UxTKpns19dScWkCUqpGoE6mnUdGKOSKM7tZOG
Hx2PXVY6mlIWe9VnnemaFE1lmVbwzgbPAjXq8zAiLkUNzZsvi1NluTvlOZpRPcXyJJVS13GiTcAl
z8Ji+aRLUhoUYjJyyuQE+9ko0yaRzaQqNoPWTuHw0XyGhsbWgbgxzdSAYK7TD631SYMNhYTSQyj7
Mf9n9gvpYVLZ8OAB02UbW+iCrW0TYRND/teikzmDeqNCSIvpAsla91FZOKafrUd3nmSNBPMqmS9r
ximc8fbZQG6P97mekk3A4WigZX5eSQqVbAvx3qURbbBVD+2TOIHgQeFjO9ymbIxOgv99OKWncCV2
xVu+o2uy6gUqDFDUOCiSRTcHSz8OdtoH8ey03K70YL3/YnaHr+se5VYICtAX7vhWkE/ZNVqaTbbL
n7QsxnBSFpK5b7CsvPmevqi3KH4E8255f2TkhIibTzqTCXEXBelFsPlVKbbP6+awe5VlP//09+cC
HJmvbWcRJaCZqzvaE/SnenyVIdMNkVwmOg1bJZYosT478eP/JCZSY00PqbY+x2Ii8zcetRdQNHYV
4F6o94TCJg5L8B8AKAdVbnl2a+NItM5v7gvdB3AoU7LB062TG9gl+bzpthRxRE89a4v9aShGIkWx
MQe4JFoIQpJTzNIw/cTK5J+R60STn6xSE6UbRhwkgYP9ASm5phEVR6EYQz7aWZ9qj9WSNX3rcikZ
CzuO5HN1I1J/tVp7O/8Rwk6sutmQ7s6LPfzM0fClMYP2sZqKUWXixcOtKJX2+WfIpD/ajNMiT9ZY
Y0FlbEKf9NWIMMjTuOwAnLl1NEXiO3mViXrYxvqUWvXgXXF4GR/NZ7l+lHhhMg43mk1gFbjIvtQM
yHUwARCTLkrEFQdi16UpORHROdzlIQW4ftC2Qre55ARaJgLxrRjLcg7flkzxxvPUo3tO4ggwjXuh
rc0XMMxkbWLM5yjT0EjuCtih+E3v/5lENyNLebsrYZSrfOzNYiGNuivC5jpWJ++ydpnlHyCfkNIR
CsqeF7KH8VRclxb799qajuYZDQV/LtOPdJPHHoJF8sv88TDD/oL5Jeu5ec5Q1Le60dMBtlYgm44y
bQ4flmaExrqbDpJuxjjMgH/W0yKs/+1kfgw4oSofeGiQx3T2lzURdel195rAYv7sU0zW4izcqx/A
KnUsPU1EKzvTe02cYJfZPNvrjaxJBdUsLJr6vjYxkMae0wHIa6aIOLHcpTg6sk4GDL0WIc9Eo40v
ESdlDLy2ekXK+jCIkrR3rHMMH+z1ErQyWqjiTgpxAfNlW0WLFX+BHduiKRKxP5nJfmkpCGbUrcCt
fPjC6ohJ1ycb71X4P5N1+1NSvGt7pWiGYieNFNXlAq5QT42VClHFfePPlAp0NaWfFUoBcCL+QaM5
lS1tNfolWoBWGEjSMozHb5jFXLCTHrKN3/lB6RthlIOpjqPELt4ZR4fhRt9+SfmsRe/vttCM9C7o
kbZq9M3VvOlqKBYgqubs44jNVNZo6JWjXQLjCdZIxksLg8yMXh5nfIxI9eboDcS3pTZS/HAucR8v
WRHOO7e4P9yPvGVX9BjelMbNRe14YTVbvVwfAtrY/iU/Jp1Cm10c9tSJE/fSMen6RY86sb6APQsd
HzVND/eTNue8dYAfPxG1YN0+LIs9/kDcs2Q5S08FYFnqfmdq/1OLl2tVC0Sy+CTq4xen0+OzQ+v1
iSeWHIfiHv+yE2F75msBV2heQmZc3X9EGPZKpn3niLyOlZP0Rgfn87dGffLTKwoHZulAbEdPNa/J
dB99U+IeVchkPpTFFT0PdlPyJE4EtESu5Hi1g30NRZ0TMOUhRZGRijtpPn2HjtJU7SWiLtMbLlk2
Fb2uCGj+bsa+P01896rmHPPGMAevWqgYelO0vEgBAWeG8mKop1LlJivu4Ax2opYgquXhpRmeovBj
TQaP6+9TJ+Q3iAxCdUkEP6RLoTas8fsCQx/xKqbctwQH0IJDp38NXTz1Cxj7sSoeqm99DYuGmNyq
ZUGfeEJ5vTspL4ifGOIxGTptwdBRNgovHk7/r5pLuIhpsmBxwKiNlM9T1+9caa7K7eoYLFrKPmtG
3iB4oLCEFKKamanbJK+c8xcF2wyvEnmPw/0Wl85taeUGDaDJve9ZmqURh7B6OpiUQYUS3CuKM03m
/errvwZqimYHulyMs/qQ7mUiFG3XWxnMwNFLwbu6rOEvytmcOXb65fnHEzwKy3cXOMKmKvIgo8Tt
Ucg5p0AENulHfq5RvK46x5Lf92UbmHcGaWVeIgQv7Ha4Yl/QO44w+ay8dqLi3x1tKmTQETU4TPw6
eeFeLgzHLbFKeUarh8HfZFPIop4ynogBtEUTQfR5r+G+1R9rthyRTNJF9VJoBnrb0p+tAjMXuvOg
igulT043PHtbnGN7olj7lEWaRG7Gvp1KIorpG5p8iTDHC16z9kdGmCdLoz/JuTwIIKO5AXZMSK7M
O0ghGL4P26hzdQ+N5lO9OM8AywmsilrIfcdPe2AMuwbpngF7b7l+vHEZAWi1oNH694ShP7eEV2yg
6lSyciciDUcwXJfddQ9F1uI5ZLHkZNOJUh5Qf9Ftmo3njwLsM9Obj9PvoG+n7WXKr3wBheDpwJ9W
QdF85wJh+FSM1kmqtATECv5S2IfCkAoufCm2vDn61dGryc10EHV8gjq/tImhOavbn7/CLJ2qT2kJ
MSqi5SBTmZj6DnaDQW0RheWJ1MD2KUVquUUN0OrtdnXmg0+yf1CVzFS09Kf9CopxGW4REEDThCV0
VxnmnlN7HxJT9dlcXsGN3OyTDmABVb1OKgcnZoGTMna9DfsJlhOvb9CTtkaixncP9oxvMt6k59Z2
fZ08+VNyj+ztRjsCDgKpGNQMSin1vYAGrSvkNLnH+yAImgjoNllQSd1Rwb8VhVbGJRiHDmYZvxJW
/ZoBD19/m0sx5dPP1Ztpgc0QZEVWZWHj/sDLcfoP6Mx3LHg1FjvDancd5qf7J+Sy0zucJ+pkD1JZ
dT3vQo7jHPMdfyvkFJE0xEed0R2qInWDsWVrLB+iXIE/fZuXk/1j5Qzw7xL/lh/YRJbh7XNNtTiV
bWztR/TiDetHE3/IXfYmtiIWgPU116L7dCKnPArOLq7+7LZR3B713AeP3HgufxPsRaMl7uYysCfn
i7ZJ6Q3p4IKp/oaitbjwjCWo6v0050OIBN+mkRQABWHBO3g0d4Lwn6Uwq+JSnhZHXyKMzN+ZBMDq
aE7mKXAH38oCaOfIOfFSglFvRuhZCBly+RLCfb1Ubl9uhciN35xsdqnEXMjTTAGJ+krb9JZAw+K4
IQrXg1KpmJUdDM3wSySWmEYMyA4uykSIrMKxGDoRmp1jZ9+3My9LhFcQabotztj3VSz7bWYFCJMv
djZUTKGiYhE1sOfEfOGqErKKXb6nQ3SqTy4Mfh6PJzPxF0yxbpl94IoH96ylEN1EJ+j20DpNS7TX
+M+538dg8A/+qJV0Z0ANLIgnE8FwuMT1z6UFWpNnYBa0sT1F5Utt6zm6huQ7Xhg9EGK/58t+9Gn/
Z3zG+zdkGAbUZnw1rGbEp1nhexGIhKa4lQlJi1+20MEjefYoC44uJDAccYbqkU4b6JNWfQoGrf+s
D1T87u8Roa0k7B88Yu6AUATlhchUAKUzJg3yTFP1Kz895o/grQSf7qzSG/WItBSVdE5KG5bIv/dN
DNrQnrwZXFOa3k2IVnz9o4EYy7iE3NxaWvsHC8u2cuZbjDJZ44CHrTDnigrQ55Y21w4KeQGQrwsS
Boqt12r9pNMPYbkJHG+S5TNXcvaCT++FVcY0BrU3RA74i+X8Lo7MG+kYbdC1J+MAvGNfZO+L2gyP
w3nfHe1Q54GhY4othY5YN8eDrYqo2bm/pv+v+YEvM7tpX00xxm5kPfWtUHzKEe9CmJBWNfg78VFu
QlqXJdFA2el1tlWY/HgZeTtcjXwXr8DShPrgSNh50kUoYcEu2wpkXdHpzKcettTfEaqgBUAnzeYy
Rpk4ytpvot515Y7zTDAIRfcZjQcam+cDBdl/wJDbrIjsImJ4s6IiM+4LrjaI/cuooFJA1kTeB7BH
c5/EOxmP6ooAiPVgTHvpSbCsN+ERvt2TpBTtmugo+qx7W28gBqnpKjBCPnyqyJYOB6yLXSb3MCmu
cmJ0RIlbQ6Oh/Wz99kGFeGFeikf88nfl3X5jpKMzaHl8nNClKL9boe73es/AKteNG3fPH1Wjn3ns
uK0OPNb3+WOzQlk+hoRilSY2AXPWvGqOGqSBJwOrHjN9J8+vJEA5kiCP/9V5vTvmLFg6KsVbMnqu
ZZosTk96tJMfYr7GACva0SRnZ2kupp8RrwBmYLvP5luxZrGjUNWesWbQz+sUajIAnWjbN15nKMns
sb9nvIat6/M/SnTBPzmHgzHlgUGC9Jbdoqe4MoPMQR2Td14hvo8TLaoXJCxJycV5m7O63FFog1xC
Eqeu6BMwzgnPvbwT9vPd8kizqo1gh2kpnvfhsrPnXEtiyBsxoIgMjDAklY3JgyYnHMN4MoFy9OlB
OBAFfXFFgbUvBYd8450eCq0Rfuw5sTjtiA1SSMI3s4GAErfK3gLKB2NbP1NyjBMYy4GRpBLccV9e
pi3RR/+oDFTkgD9tJ2YeRJdfEiKRjbmbjIubHFiFutOKQmCrTG9S6J1MoBT1xP7ziJnbQ2e7wTmS
/vsvrfhEva3yqkLFtXilpEyTjJRPdzFV07EKyqP621mgsMy+UoBHrnzc/Kh5wdat9mGR35zNiVkJ
omaLmemUHUOaPQ6dQLgS3334HbltyR1MxOF9DTg+Xs8vao4O9L3Gj6BX/EaFtqejaEBr25jVbbIh
pAV6xmex/T+kc/oQSr+WBFtnDoI/xSiMkqfTG0GfclgvebdTibhUHvOzazY1IfLm+zz3sm80gKJ7
B3FQwzS4cdg6kdGK1e8ufFGbI7vmpmee6ty366BuTSqwwFVtpvO8cdbvGQ+ZNcNavaqMXyxEzu/Y
FMbRjjbdf4Pnq/hFXk2zWiLP4eq8T/xpP0ff8I0rh4pVvuwBuyc5k7l1NGCWRfI2TQVgOvAnK8iM
9xVs6BhUL4HZWECaAwmj3UXo9C7fwVaTzPdjPC1TQO27qVjRSrqSrCL0OQStKeD5rzNBwbjpHRzY
Yc3M20dtN9vw6wxeGn1XK/g82az1j8LNtB1a38RzkcTxM8e/FKxL8eRfWjvraR5J+W6+yyM7LX7W
LipeCQa9ANBrSu/7PCm8qMWJWfw5WiwnQyM2oB4TiM6F57vaDKB/J7iHOho4krbGg2YB3wxSOG++
5RdA0CY2xKQhBgB7A4FCzFwUsakOmFx8IVFx4HWkzGkvdvVGSFT8EGs6mX5aZdbzMVcm0bMls5qD
VIslrJXyw5YkdI+EcwJFHBLOsWkYCf+Q+SNskGbN1jND99rYFeGMduZCdti9nqDseYgF5DlW6SMP
5gfVMEmZtQRBFTttq+oq4UwUc8v/m1YzyqtcUWqIkEPw4RkZyQoS2B1+J/GPKOzzlVzfVsyBOy+C
aKVimKrchNr6RhgaSnjtdajA89oNUlZwESabGeiMDM2ipWfpZaKqRmqjPYNjuvOkNoNyA+H9cc1q
p/prTF2ERP1QP9lUI3bz1CpdEez0oJM1IwpvD35ZZaze8DyBiIPr/eDUK5/wRD1pnT10FrDYxHJv
flWRkSIq1d8xX02a15BqPLln/UTGK7FkTHun7mxEOAR/uxa4gdU7EibPIYWBZ7DgETj97+qnYOfl
7Mvj40gpwmRJ4lWrcYmmeOzcHT1Jg/wBu988YsLzhZrakaEbDgJEVL1fGQ+WWVitHTY2TUg1Mc6U
+0LgwdhCT2RXcfzEWplGmzTDdrNxswGWCGJzfcpG8BTO9PCNuH6AxJl76gRLXD6cO8aki6CaLpHE
L+WTAIVnrg/r1PfgOF0aV6Hjlygxcfr8OSovMq7cg0XoOhSZvNXUmLUrbAERCTzKFAfIctytqvj3
l5M+jXLbHbaJVSFPKVit6sQGy1eehVoeUMFN518FTGk5k5oVI5Ekea/RcFmWa5dgXAZkiv3u+Jrz
KkTIQaAvSMp5vS+uXxnLEQpOmFIt6+K2pdHRKWTj9UFXZqyEwb+tUXj3tpDq2iU5jE/nZl9lRDvM
DqOTexEJ97BEH6mM5d3WqhJhAPytfJk8jG9iraaThKmSA2hTU8AEkAsazpQVhw6x5wQ2FL+RciPU
8eDDuLFef3o/ihlFHf51PoPz93RIwtF0vjA6vEjtkJkqOiuA/wAOrxDnVHpLorkd54YbCJS7ShOo
QGZb5zsV7Uqk3DJX7TW0IpuuHmj+04XiAhGIRN8Fg4pq2reDFBTLGd1Nm+MHnZgr2PQf0FpiN9J5
51AlBCmQlVi3oPPQdr/FiE1payaFzBNBnzb0u5vMidVxOth4kuXcwl1peBJ5aCc2m+4JBjoY4Rxf
ogKSE8mNWuOwsvijnuWohE2/lo77gbeqNvS8x+3wDNQagyautbsZjPibCdyrFmr1GatIcHhfllkK
ZJZ5YzYIE+o5ofH+Ja6I7kWDxKTzMYdV+kFaSUKm1muaLAIZuQcy1IouBbUx/W/lZsJQK2YsPMHM
eZ6PQmYjbd4ZD4cd4KYaVFVNPp61xTWhiVgbiU5du/HFV9dABGy0n3esBP3llsxK49v6AGcKlVsW
WxcTPLTwhlPo1gMVLA7++ba5imYckrkp/J2PXMBjfa18jNd5MIdyKRVVSx6nu/cCtTfnr8xkHtjx
nf4yhH5Mg4a7Qv6/vSKR2Q3+SECcsNk7Ef+oXauKCpRetZlZqAM7Fs1qiNgoyHV7ngG3b2cTf3Tc
tJeliqboLq7Bx51qz9QohD+7tR0GP8BsWfSmSXpgxfyEaJdNfOOvlKMBjUfeZC0rMccEm+wknPSR
xXCWg3P2mq+vruAnzjwLuG1j+W3ToY6OZMQae1XwPSp2iwHp4sTQuTk9VOKCHaaf6PFQTvPG++4Y
hajDNhBbyAdkaFiP90uf/0rEJ7NJuhhp1BWZN+zSASCIGLwuMWTbABUnryXOKXieB6CjduFk7X25
xfiG0Jk9Qhe3tFVstvNI/BDb3FPXEdDnYwSh/AEOvK6keaWTkmXvrwRXOYEzIskPv+2RngqBQhmA
ZC4/GTlkm2SHhw5YJs1zfgPozeNzsFy/l7Cq5PXt2OGG3P0y2kXBSopDzbJKJa59ttwW6kvzyp7z
gmAcbTlX78FpTK1ooZDK9L3QivO5ytMv8Z+Wh6IU1di8R83aLNMvH5oOKoW/ghv7KHdlUkJmCLZq
MD6MHwyOxQnEocmkKhc90Oh5MsjiGhSgUjJSx5TxQ9g/alwvTQNHwp2w/QVrhygwZYufIyOOoJQS
FvcKH7/YxyAl4gXyX94xdGomtxbqFHZ/JoH4CTethfIBNv4twsaX8trZJXKZoCGulHknalnePeDV
W6ALS2P3EYY9OYNMFbQtMj3bzu56JoVrVLd3hRiuYSOV1CqCKltdRIdVFKVNl7j8aLvSlP+SYzlk
Naw+CwrcbDGdSkghqyUfekVy6tq0a/niVAizHeVZTMjtJcxS5c2+R/cOSyM4ED8DuAOBn33gZuZw
L7RnwSWJN4xxMABC2vE5IVAWLOARefsxzkuZSvVGaQ9H20JWV0HnnNlB9SAUlt5Pxrf67eqJxyQX
tNfTx15mw3t+Nbr6HyK8o/w66FmIwKjoQESvjlVUMImL/D4dMG+g1Be7JXIZPJ8eoGpmnZ+SpaED
Nswpv/jOVCEqgkNfUPZ4tAEwbNL6s7QafmyUOATXODB4L4eTsqdIKXctJYV3QQ8qNAMHW5EqJM3F
NmoLs65QcgdpG6d+yisytSo2wOw6EERqX4Z+RjIS0bZVHo2swfnNqSQCsAG0SOgRUhCXaa9nptzE
d71ZmgfZgef4dWpOVVeq9JMmGGfbwi+B4jDDzevI1Ho1RnkBAuwEKiJdMwNigPWLrt8oUd4BnG4+
4ms4pJH95TnkTS/DwMAcksCbF37hbbOFax5RprYIY92A6IvsN3rr7+JCFPbYBl+dLWncEwkv4Bho
40gAUx48S1HmXbcusRcM5X5/PKE89PL/n+C+t7eO084QH2//Vx52adWNrmwJGKrhPPy8YDUc5cX2
VwO+MpXgQ7sN94JixU84BfS2ZKoZOIXMExF97P8XiXSN3NaXPYL02KB2ZK9LqkT5hZ8MQrMFrTcR
YRGm64xuWXB6zN6kVVRNCC13F6r/d2PjyQ1zJ4vzx3auMs2cD6ePOjgTHoxrvEDpWeyGqP1gnGMA
U4u/dwmEybuOhffN9vjF6d+th2miJltWuLCjsuLisGxsx6ZAHLK4H5er+por0kUy9eMYeU4wk9pp
4MnHO2X1LilZS4a0hGTJxAtnBzeKy+QeQN3BWRYOjFZWkY96OE/brnqj5abC7trhKZ9EScapsMUl
g/n8AgfoHZgGZ0dQal8WfsQ9cXTRTlhbAzOl6W1HJqy0H3R8O9QgD7C5Qt/fxj7Jxk3cJCrCVWLK
LcmManpDZsbyZWrzEsJV0mrZ/zOfXiN3OdFoDPVGsg4KbKEr/fkpNWe+1Z7QddE5tCT8Wsm9msmX
nmm2kB7MJW4FO/EAd6b2HNljfc7ulQcVaE9MBrOhOUiVNXwtvqF487ccUTF/fpn2M6Wdk70SLCiX
wF4YSdk6J5zXelSSBRltSH6jmgluFRUDSRwtCFEVSmqin1INr4hNm7Dpu0EJO/epn8nC9ewmrXNb
4noJiK7pPmkx68zMZsQ5yu6N3oj+gzTsj8332Nv7L54XFMKlU9dEbKPKx0BC/QnuHLflkmbURPq/
ohvwBPOuKOHP1Isuh5uH+/ehZA3ZRH9EXBdHhl91xgubHvA6hdIzoiZfnmmYOf7QGoq1jibyNbjH
0b7cD6sJeD5oV5oB+1ORKfX5i1yXMQv+sDP0vcM1Eaououh3rccZxCtlBUJkGj62VQuXUEixTonz
hy/op8zqIMUUhX2Q2dopqOO22daFrISIldy6LHSqYY22sv9LFOgqq+zH4isqDn9Gf4ubKyIZ8NnB
8cQyZJU9HfCJ+d4KCCWjnD+5JsCydlmRi63IOpqBZLISFy7D8KZh6C8H1HQ6pAVdP17mpOt1pbA6
M9/K/nANmNjx8PZIzd6qKlEvT++t2yPfJ4McWD9sjdvEH3dOMIDO8nJNeBG8tfRDe+89j5fgG5MQ
/OJ8RN7eZHatLCcWdXICzUvBloWWuT0OE+7kOE3FJxN/Q2T1DbA2qs9/GDgMwmHsZOBTsSeb3eFC
X3R4mmaoVfxS9BrPWAoBCeMoPDcShH0/7GBVVhCVxestmRMOLeqWHaJ64t/3XJtZX7AGP2SeNUsQ
raaPSU7Pf6+k6Qs9nWFUjw18rOnlLJ4nWnTnZ7KGfNTlOJN/Dwo8NZWkK1y2cP16FQd86WuQ4NcX
dGZbeXdgtQlVR3K+Wc/ty8g7hihJvpyhr913p2h/Okoun2oYAXhV0a9Uz4cPUo0SC58aSt2/P1dU
B7EUWM1iw0XXCHqvR2i2csfe/l86Z0me2GpfyAkpwy75zK4x98CWPwHwxlpCEqYPa6Zd1XSI97wk
1EtOHbDbIquaL8MYhFVp2KQS1DPkHWDHgXYsTHttTRpgsKL6JEiyvC58QsnTIBFHT3Hn61SLOmdB
mkMv6lcUq7NZcF7cwo5Gct2CJVheFaMuUoSlwXXLNQCGo2n5fMBRj8jxLGpZpqXaSQ/58CXWmMv8
vcLSN5oEKfQgtQBZYGk93E1n4M2VDaPc59c7aPW6ywKM2pHHIktW+WULG4YYWY4w+ozZ4LpINwop
D5+LuV2QbLTDsEilTs7GsvZV/jX477+ws2dz7S9OdqFeilasr+2nLKusSsp3LG/nIoLLU3FcgDZL
4BG95ErwEN6mzB/aROJgPR2CgwzxSkR2DGw1UPATHywsal5yj5AdAJSYLOS8zyiifPNFxnP9SytK
GQUkWTg6SSOCc4sT2inZiw8E+9ed+K1co/axuF1N6KvBD3BO6bhwEJAkO/tDJW2gQxawKagwZkWL
h1220mk1Vi+sRej48HbuMFPVAzXChebABWrEmiE/ydZN7fSFSHjO6/C7CgnYGT49ouH+cgK//ypY
R0PJAcZQEEkoYGO2q7QlhtM9HqMx7WHOhPZmKVHx+jxOPDoj88zp0S9zA7Q3qImZ6KzU/HpkQqIi
hTYrOVuP1lmwkv2yoHqP1dgJORloDQwoS+GjB0BBAz5K/0GvJRf7jxqQfBRpxTeNTIoAqY6e/5fn
J/c+PQPtTrcvIA2Ze75iVgs2Bo4ghwHFOHWnXpdatsZ48q29bmPmQ5XhTNo/epvFSIRadXuTPcAC
lH3Z6aHqKcuZ2LxETArftZNWBXfvu9KQgKHeECebZPPDDPDQXuZ4o16W6OtPcKmBexB7vF3SApyJ
0myiNPGOD1dZGKR1hrQHHFCif7vy3I2hZRtkZ4olLHZKApLnGcnqcHmWotl7M60Zw0UfFWzSHyEF
Xgn3IcWzqZX6GRurEOhJy6E5nODGKlw6Pn4qSbZqFQls5jHbFjJHv4wBivn06VkzsAGWu7k9YW0R
HOsERUHl9bu+A19gymb8Jl15DVdrwirONeCxXCB9jTcG/QhPeW202BCDrdv44X3z+Z8NuusYCoL/
JxVVo4aWyTqNiWwol9j0kgTp8Uutq7Lr6HYCUlrMFCNRhZE3n9Zz0NqgHNPcF7zYzg1HcyTULGcJ
10wSn84eq+yd7OxuinTk5j3+eDhrpK0QjBkNiwcPHpyhpPiDHe2+70XVgynZysbJWs3f7f/bpa66
VJVgKIyoKuLaTnTyKgEDkKIzdTjqbK86P4KsXCyXVNGoRnca9tJXvbt233RyPAlUbkFq6wCLOjWf
Hnmu5qYMiZwuWYrgseeq0H/fWA+ThELFuHXz9nDexusCB2ZvK9vNFMa0TjFDFNeQ6R8Rvpkg9iMH
Ut/Rg2UjFyv3hiCkmWXotixTZhldplhpGrUlxwbq40y70ej2LMzuE+8fmslGaxC6mNee3lQ8aQ20
57uNS+4BWO5riMY99BFt+gL0sRZwBtYWsbHDJvkb3+UOkdJPqxKwqczS0Sp3k0RNc88h+XRVtD8V
yzw4OOKWBNLxm967+9wQeaGkzIWWtJvgPVx8CpN2auyZBb0ZIrOoFrxlEWl0DyURzM8H4pk0H22f
0Ni8hUBYaEFEoBWePxMJlyLVHxu6zv7zfBR3/B5N7C+cXyTz0crCtP7XSMpWRwFNgaowprnzqZ5V
RDlGU9DmW3vjwDsBJh6hVPfO+SLhyTsbMycYc4DG8Wyuj57c4KGSLtG1l8lDy2yGEUyiaCaAgty3
L8HmKD1KSUbUSf5POoIeXh6dKslrqUWmMGeQlyh/R8BIov1PeqcODTukF8yiTpSd5dCFTcfljEcd
WRFn7OuopKBluBvQpLVYSHUPz0O6Dk2oO1MVtvJGKDi5oDyTspbBgp3U9z/SE/8geNZepUCooV4T
luzUoTyisuufb84Nncqe6tV9YHq701/bY66zgaEhfVNWLaWcQGTu+5Ij46kWdxw8NxckaRa3WfSY
Zgirl/Y6JUDOlnrtEKY8TdSWOceYS64LPZFZ5YfK0cRWNjdG9YVqPXsBt+GsSNXSCrY7NkVAGpek
W17wSshgFRdCHlr883MyM5Etojy3mXgNsZOpVsQsSn3CJDrHFDdoJHcSOHbahhU+jHv9Luv4mSih
rB+Z2ZHZYyYHKlQ7XMbnIt/wsbTaMrwh8D3OUub4eC2EWEazZLgFqtYgAxbOSAZ05MFJ91i5cC8P
DPntEP6BG9h6ZzIBHvo1kkmI5N4tHnYDpnTfLYrCNpMYYhmlsirODVzHHA2qzB9SsiBKvjLgp1Kw
DhL7vOGvgRf/UIcD3Lpo2DHX4hdYimPGPAP9joKZJ1+XtjaN6MmtHwWxjV51849cdoZ5AefutLBc
5fuuUWiKAC+a16VdWoz1XClxgNxooihSfTskoYVtbcGoIYlNiUOJjAI2/fb9bJimNGsLSFXwgRdC
s4Zf1Yhijf1TlYrfeacMrLansSwWeVAgE94byChkFEVx+8tcKQA7qwurZVr2/sQgZKRSOiVntnG5
7zYTWwS5IYbb4C+SPmzysDBdzQFckqD9yfvql5IFarEMYvqaDPJbiJuAUvBV2Td4cFXsLN4iyGZU
eVjmK5ILIN/MajqGqhoTrxXbIh41UBxdVI2RqU1HPJyb9cd8eClLtZShWhfniVDV+zW2noupQ0IX
0Dyeqt4DE+DHy458rejd7SxzMRUhQZYjC7ypdR/Y5QsksLyOJ2goymiEhyKM/2oVVkKqJMnPbk77
n7aN1bjiOnddGDCzyO4rFnZZK6PjlZUE2JOEjDohQk42epc//VdCWuyFvk3DSLd6trVmi8RkcWu4
S5Qhxlsa8RACAapajS4sIVSRQ1S4qlheZViH0biSSIjDGLjnUoTYL1pCICQPMuS0mH9zGONXJnFr
heviG3+PUWuKHYrWLBx5TSeByi4V2NXfRAa9t3rOjuyg0LOzoXi+n4l8vSQ8Y0NEV0w1APfc+Inf
Vmse70r5kjxyHyj6SehVl4EopEUqtrFB/SjN7raUNkbNeA5U/ALCb46jVTg+DaotlcS7pQN6ZZbP
noc3WAwmcYXV7s1NvA8qpJzXR/DvRIcz1IY44n7DCny4BglY2uw+K+eREhkS7C/KqRnYY1RiG0FT
//o0cz/GDuF643RLEEn6MlZm1IxTxB1Nu0+VbG4uTaOnlX7QANwfaU1/2Zu0cJPRrWLNa1ZNRr8W
kDbrEC3Q/rx9xD6SO4tGVO5vTlJF/dnurToYh2HLul2adsKL9Y++341pUPUj3aG8/96SFADOEBN0
UKwWxeIFM3aoFK1xH3IsCHyoRVcBwzxEOgrqHCNLXjjZpqv99cSeTAx9vPOPxw1zh7G19YrDtVyU
9gTFdxr0TCV3TBk8oRxmPUiH2YNwLKPU9nD4/AKmRD9XezohX7lplcOfjz99RTdCCatdnQl9MSQl
q911KLCM/NLSG2IjlFfqp34ikSEi107HJo3KR1S08LPK0MYrvEKavvqHaoDKNOEQfLStBC5TBYf4
ayeiQMsfiHPOHiSZaBFVdPRqoZMwLJvpGGK86q/T5C5BRF/Erj9ObASBX7/XMtekIIadK/0nkcF/
Gqi12ZNInluh74cfSX6fj4lMA+fMsA6Ej84P5LvZbE6pTImLEvAtQ8RN6qDqN6E1jHxslqn0+p3V
lIMogAtZDnWsRQwJ2cFO2AElXQWgM+dD7/VYceaUqIBHh2WnID+k5VWmwdgOsJJk0M+B/YP7rG8A
DUf242YMfVM19Rse4F1xvi4zHjYdIL1HPiKAU5L42V7yG47BlN42Zm0ZRUnPc42ontgsKuwh3pu6
jj4Ln2AhTp8aACXgB8iWpUOZPyWmiYYiAj2O88CVXhE3XfuLtRWuRK6q1ZzKLyMqI4AqDwPXurqp
dJlB+QdSeUDnOr5la9j4jNUCabyFytmPQ9QGGZfe7iNiIMqWEVsi+8f4RGNjE45/sOjpOEz2FoBp
VVmVsO5BLs4g0ZhSrrtMTr3N1YpTZpsRiQVzvBuK7LgdY+6ORgt+5fV9KaKuyWsbyzt14eHnHDug
fVuualFGh0Psa+tvjHgVYnw19Cu5/8IsV+H2ppAFfrNsQXEPARL3MHB0E9NSO3RpWJq2C4PUo6ga
I/kSyv9SEAZKn/aCaILxk6DxYyIyTcpK4Qp+bjB0H8pf6xWhZwnd+XRk8C1Iwp25P/sytqdYhOo2
br5zVKk9G56umGNsiznZE1Apz5tCY8rPZstFeKk8xIZNB46q5QnGr77s0aCV3SYGxVyEAJnrJ0jL
6qUoxOKn92VbxDOn4pT4G9EmLTVBJExfQlsLmP0pWPyc1Z05UqGVveNsX81tyxa5toEJEIwgWCLH
tj8/La1TeZMeovh+7cu7Dszpq4rnMp3edpnjswPLsUJ9iZycoaapl40Ksazb/TIvE5NVNh/CgXt3
e04Uq/c9jht2yYxG/sEZVfM+HKHaJjhzh+76tlyQg633tlhUITRkMCs46znhxKqnNyMkRHZEgiMD
yTQOEGkr3QioreHpiftjFt29F8aQan20utgZkZiiayA2xNPOlwaGuvc+DgHIRUlFpQb0K9UwYIMj
SHJbnIuWmvYbG8ct1h+Pec81ialJEXLyy/YQ0ZGVKE0rpw9qNiRG94ZR9Nof3ROb2BB2Vxakqmd4
mY6dalNX4YCV9AbB7JqdhfQupKBxmhNimpH9b0hIMbKSjf9qRmT7s9qpjzOY1B2LvN5zsQsJTjQN
XZp2K5r75cdgJh1RaNp6CatUEG4WIOKwluDlL5QwjD5U2Jt+8/bw7JZTXkfiYpl2BrBOVtErtVX8
P8ynfDri2bNXYJOUe6z1BGBRdlAtKgUXjbaULoec4hjXSlnV4ijRsEcGf4wau8qgE8nvWlOlpNdf
fH+i1Y6cQcJVM1o2WtXjZNSyX9ZxDj+scTrfzj+7BSmkF9dycBsaixEkaNfiRAvM9ID8TqPHzLpK
AXnplCyFxRtZrpB+Ma58ZahAnnXvgbUFJgaTMGyJ22xYCwBs1vpStQSjOUvYu0hAG7VYWon7/PHb
kMVx62eVVfTwZwShsRDTaSi4AzUkiOy2GTzJ6tFVQ7nEitYLseAr3mP3WWuwkYvHTsxBAE+l9DIj
4nnjWH66Gr++yVGHB86ZkY3+b+wyC9HTHi2F/vq2nUlgApbfXFOYmCtiagz87Pu1MTGmDnS4UG97
I0om2p+5pBF/buA/gNRza+YMBGaLI04+s/99o0ko9DQU1QVrriQxF3KoqhJeCUucVSerA8siT3fx
APiD7wtYf90GiakDHKDfUVMSyxPj1szjK40PrkY4KAbUjvWcwnLU+cIH6+gYsPHG4gF+l6gpE0vI
ma4gdnwRG3ANmnxY7Yyyvjrn8gSSjsTMpiUQ1l+ySx1bhHiNxjg7iNRI6SeHXvw98bFwTyGkNjPp
QDKoPNNaP7okWN2K5BLaSTPLwL7rC/Ay/WnrxPczZNEFBp1GfCboNqnnWRwUYKPM9yI8i1TF5ahG
wTWHDESanpK4gRJ6EVuD+fQmG09PgSFu6kW0xfUV1xG9crIDgXC18tkBemsetOBBO/GjZFW2WnG7
Px7r0UPFLSckHYYEXBJT+htaCPX3TiRTvX61UkLR/KMttOmET6vuyMG4KZJfvofuwwu3PX6bLNI9
lfeeyZ8AllMaHzSzUqbFis7Z15M9+pIN/brLBzMh9+BhQ6FWvTiTdp4Sgjl9mDaU0RjIqZfJV+uF
cFPIMzRQrBudwTzZUj252q8+t+DDsSjkTNAmke/84RqNYaxC/xOmo0kueywqvAwu6wfdldJeBiTS
uEUtMINXxVNTm+UlbpxEwNYU3U/lTqus3R1YjsSTXVfhC2owtBdLG8ZDEdv+/FJYsAY8rBdBB+z9
smcUNzQnaXrPpbNhyMGdnlR878mFD5F4zcgFwIFXClO/a6SsD7mIhYDsrlHv1h2InWwfPo8PgTwv
8W8iVnY+mcwsQihqmjQ3Zqnik/P94242peKqTlauxtAQ8UxjinDm9RUIh5rZiOOxTrVQ/t7NaHcp
03XyVxt2P5WAcKB9XVqoZKESVVDePos2hBVk1rlIRut/z5PPN/qa3jQp1sQVcHMxZhg6XWNIdgyh
azGpIh+zy/UaVtG16pTj1pC0XMWzeFXBMYDjTS9SL5qaNYi5pOvXH05cmBKh2AZZFAvqwdEGuG0g
dZhVsWWOs5umJNE2ha0tJ4+WiH5L8GsCWQwI5fwrYrXgwfWXYwZ8dauujKcfG4AgAO/FiveYlWZM
IdFT9rg1JEepF3j5pmqb4HkaHmAJ9rJr96712n6jIuwaYBxAi2DyJ7xRYDvO+HrpaWRBbdQ6iteE
hI7wLtYN6iM1aOVxuqqEKK8PkB1EHEIBl0f40eBtS+du200PQwPP0ngmPxL/YIGTcdzvjY9RjEUV
u92ha9ZJ6rg67jfdIy0JoxCfOPm3/cHcHZ4//TlLmKuOSkOx3gTy48+nOOWbxxzZtnzTm+fiezEP
//Py0nXEeQVAW/pt4p606NSE6lxr/BnCfCGzPK+sixtKEmE76TON/VgqlrB/xuf9bURUqa8KydzM
ooH81f9hIb1/Fs7qQaHguK47T5L+JfkqFQ6QW9nrVUzSEQrLZu7YHjVd/DhWuRGpBeP7yT9pSxfI
yqFW9EIlVNKhGHwq2yPCPYlzJ/roNYyjlOIoJjluHpArLelx4SM2/ACf2tAoLwL3P431Oi78A9js
lMJof5y70n2Hg9R4eV3jAeUrNSQIQVLVJzRMd6GiKE/I+UOsQKLy/vv3/9qhaGhczFns7OPSChQ1
nWaS0s7VXnkQ8psID89JkUl/AIuACfaSOkTHLqmXmp6tF8Sr8wDIFWq2nPkh5QnwkVIpU4TnX/Yn
9DkoE/uGF44adGKFp9KJbAxTKAxUuSR64WD+JvtJ5n+IvzsQOC1gViRhSOW0+YJSZ/G2MhwbDZfR
VzktjZW1eh6PWW8ai+LLCZrU0FLGj6x37+3VgXiupSSR6z21OtECLNh/LDqp28FV8fOSo3hN+CNJ
4U+u8rwdYItmJ3rUJcicGEUQhQnN+yIfmQsZmuqrdIYmgYwJmigDc8WJjFyPU2qw4vwkrB4AaHGb
pAvw8TD398oQdqkvZFXNbrMQAdQJMYhO8x26lq/viMssNxgmqUKhHlO1z0kTElrhFsvbCBAOHFz4
YDl4Vku72A/TSV5dI8gjnx2AvX1Z8QUT3AbeA63HIQ78N4dPpGOimHC80eVyzMpo/GVvclLplzGM
cCVBfEx/+VRSKKQcbStMv/K7IpiHP+ERLt5FgRmSzH5K5bcUnfzf908bkPtoLql0qn+2zNLqXAKL
Hx8bbAK8CN7A2laC92gdCZPQLPaPuw12apNZmG6gg2+SWdfiI9G6Mw5XxA6GOFpHdrZTcR2uaPdL
ybds8sELSc/6AMReWMEdLrNS7Agg2fyzBIO2FAZywQjy4RV76jPaGGuFY6MrQPXYTejzY9rxInHo
odfbXUTvQecQdmWBkPh4xgvu5IG/yQIYBVLUJ1Q3VcNITms+1q2892bKoy/KNhz/eV2FMXAgt8eE
yCWHpZwlgVpG1mS0Wt6Jl9f/PiG1JnX/1I0EvUy4/GKMvtaK2mmuJVNNlU0lZBk2aF9hPGSatEHA
o+8AD0KueLeajSJpihp2B2c/Qzsx4SwE9FUu6RP8BzQDgfd0oMYvGDA9UYF2zTYHY+5ruU44E06c
iFXb+WOc1hfAl8FbXUTBYTox79LbwO23X0P1dmNX0bCwzHWeouAEf2WEC7Khoiwz4dZKF522QO0F
QCyEVuhsKqHAEGwynsBSfV7upt8ZFraSglJlPjw5894axByq0aTaT04AVONQP82L17bFpnHn5QfP
GIJxvEDX44zEamufmCVHv8wRzqKTwDUNm3dZiqcK3mFERHM63ycUr3hrTGu4gAwWs/nPoWEjAIvU
5XhbBH7EZ1Xqe1HuVWTkXgaBuFfnsnYNxmQ4KOiad3Hb5fGDhS81djqG6EcsmrPBgzG9sKXd/YAn
sTMmsUq4GEXmL+V1mOopaL997nU/8samThMwPx+YY7S3NrGZRV00sTbxGFJvQSjNIkh6PBFDTv1j
wbE6/ep/gFAjmFq9DHStoGHyRStvyAjRcp5TyuRr1syoB3cJNuxOzU3NImQ0tfpWwSW0/8lCqFaY
vXcwRskRMqIP3Y3/+Bc68/lWKiTeEWEFCKirDQGZoTxAR7soxlUZVLTY2vc8kq2RseLxAYV8Inus
dm9NF2ETP8dntS71V2WVeD1ZRR1w9LHRpo3ku7zx5XYsC2bKqkIVMnsmMpCfY1J4pEo9e0zm3QOK
Mi8I5fg5zoC0l/I1tdAjAvY5jM+TwgXbIH77BgHOADNnQcH/TCNIVGNx0MrDOLeWWJG9zlCU6/1K
iEQ9MvFQi0M8JcDveSSL97j9HyDBYt2mfMuRFZG55FIaWc+Qt8UsOQC+Qy5IkYgOFsVHnCAOm+Q9
7AIyWX5DXwUOCuTlTXEsjKHxJeULnT9FVujxVG1rOkaWc4mycV5BnL7lIR3vOrmcFOcQc+Oo2PC4
H4r7Ad0ofbUWo1m7YaxAEB2Sa0DN4qiKAC25sMxeVpqGMJgkFjrPVZEioKdnq5X9Z5aj7grxCyn5
hJuNeMJnqUQpH0ojLylnWNOcUuwsGn/ORSfo04Iy+O8G2s/h5oqzuRYyTibZkZTXTdaiB/b1nnAA
VGWyDa+/nyQAvGP8weF6qUjyDw7GLSFJe1lRiE9HFV4XQkGzGwlcd1BdPvxWtKmg9Y87pazuokW+
9xnAZB7EZPG4QJ8buYyOrUtjyT17MsEZCdI4nFf6lJx5/4U1tUIa4GxLSi5ASk80SFPBVD5nOqCd
jPtkRtmMy7VAUjbrUuZrep7OpZrMbFP4TzsVciuUNtTdTV5MW+zfHamcve6xQzCmRIEFWO8C9TOh
lmBEk5c+/n1Ol5OaxyIcAd1lgtsoA6faIF+O2OgkepsjImttGpzGVwUcF3Srf67lytyMFTPltLby
F4Rpj66GPvIZoUp7DxcPPS+Ck7eWsrQEW0mM/uEJAc445OYZ5bKa0jUSNibac9W0FR+8U02NiEyW
Y9ft8TLoSF/basYiORubDfAweGOpI9DB1wfBL7SirkjnvJ3LscRshyA6QUO4LTczhobkVQTK0RVV
OCl1XtZdEzRF0oqsj4Og5IuubIC515Eg5qXZsQoWySXof0SAX2GCIyX6klmg+jtjzxsM2iMoc4YM
eXqW04fvNWufAVUIsLCjNUXABmrL1NPKIQNEBGG6VZIHRPkCIkim3ev9wPlrKdz/XXF81okL7MBH
eQlXMmg1pJXf0GetE3s8tQG6hV47lW8pFDKEX+BbOEpzVBEEC6YiThw1x641YRRdjAD1NinjZDdP
lFl3pf/0B8YIyMod2n394DPcRKEDTdJjy1tThzR9nB/LWJS7LDova4ShU5B+oEwE4Ctgy/aqH399
KmuSbD3BIbaPKCMVuCRF5c0/8x94VX20GxpRr+ipmZCiej2wWTrkct+I8TYzDPifywNgMV0vqXWM
q4kcPuBWGsdj6PqGwrGxCeA49+3CF4IlWZPD1lC8miV/Rt/hApICNEMQbUsknrJ1S3EDIAREpGKu
/gwUzcGQJZJPO7v+Yl4+7900BXgGK3gUWc6fa5ZOmSg+CXwFQkgGrf89iqaS9bO9GJEnmZajj3O0
w1ybj/dcNiS3w1x7yVT195YD1WcwymIQ6d/eLmnXjptfTAUDDBxwJuoHLGzt1OLPLGicYI6q3v6B
IRpsE+WTcgsGnaG4j1MidD0B/IvK66hbQb6RhoxxynXF323b3t1kVz8t7S66uIBbWqklw4X+JvHV
yaGiTUWExmekJ5Dyhi+opjKprBHIWygszA0oPQ4WvkNluifPNqls5vlbafcEEcjZQtAmjPmgzTRs
5/VAd0VtfAp/isTJyP/yONYEcRnx5vFaa/wuARtzBxLYdBEtwV/3Y69f3A0mzWTz9vB5ky8pPawI
4GxMYYrvCHlFewTX4IgP4L7d0P9rAQaUaHex6bxzH2xPV/v06lhuz3zPRcciYK5MIURV+Rgrn2IU
+L9KjNb6RLhSueZa857kiSoRhNRkHIQ7vbybvC/4jW+6gTSbELvUNnRF9prLEQu+dS5hAcVEqp8t
enw44A/HTMWxs6dv1woXr0eU052T18/g8OTdzq8C4uV7ehBME2wmnIrkvbPjutpyau5Y73SoaNky
nBMY3E+qI4xTEcX3r8coVPvW1LBpL9CaloBXh2q2blOtVytUMLIRoN9+tDKqWasz55yQK9kUZVOO
+r9EbxPbLUpmHiw8Fd83JnBAsvIxwqbptkUFvDg90DGnxJUuJdmGS3hv2rZ56oGV4vptgkGFc7av
gntTuVJpDVSR8EfGBtKYoK74vm4sfkOfjgpmgSdWK9nuiodcYIURd1XtZzvL1SuDl/R7/W0P0ECb
7gnLt8TXnwfU+W/+acJH1CFceWJQqMcdjNCJoEQ0Qr5qlXcgYqUT5Tv8hFSthHkUsQ0EtzbtLNFk
nI6qjtK09uOuLckViZkmQyejOZCsXqS0R9oLCRbjABacgK4IXIzWInstXUI1vbu78/1g7LyCABSD
k91OI8soVXR+/mhxtr0/zeIO4AkNap6iE2OBJVp1qaVEYzkNLLlaWpKAny1Yed81nB9+Ow2TKwgY
6jn5j59QVHfKs8Mw3Z2Bsbmj5aXxKFaY/cRAnbEXV5jor5cexNmuSRN5BiKnDuH6kaJVOBHkaPtO
QZIBKH3XkpXIQpe3mfVz2p1tovH+7tr915bsKh2b9dZg1dVrrOWqiL6UXqbCxlqZ7+gshFz7YKhT
Ha7t4KyaHIlsVrCrOxzN2Vi3vtiHRi+vAzMq38WZdgAqkkGMk78G1/U7ARctwPkbQi9updyh1zem
IV1fOyzpnAEfhIHENQ2S5qKfOy/wMslcGzDInfBgI1SstAPNOzPXvkuMZKm1R8oKlc+7wzMJqbE3
PKR2OU19eTQf5+yRM+f5BZ1xxX8yay0r3s+usmidxNWtfHTwbVl0B/xBCMpL0Z9UYEkdsCzd7+QO
x4pGdFMyQJW9bbdBe0lCiYTorvPSc3eCuWXfovImpHbkUM/hZl5/T6tFJ0fcqycBX31MQBrA0Crg
MzZ0CqGaMZCigXOW5Lqq13qId1+aIiFMcp5HYycfPVdfqTjyy4+0EtiwUwj9hqs8LuqkM8/q8bh4
X8x6zGZ7s71TKQ4MZaJEOE/0ZnRc0ewWMCeRZdHub80fOhBXZvJRtgF50C8T2JO+ljmmgPaTXlEf
1zu3sgfapmhRRilapXAA4Ztq7f7Df9YPxHTBWpdP1N0CJwt/JtWnQP2QcLHxeRkRok2Kd9cfPtiL
/MJHC0NIyIraC3A7udQlbRlkeoVLsBwt7f4bG17Fh1F9Ra/g45hrjZwrfTbCmJvaJ51VkX0MiDXE
m8JFMOfUkhzG9FTi+AMY8H/qw6PNjCI4yjWqt4yTN/o/X9IONjAkW8UdXRciQw6m4MZJrnehDjop
W1ayktnWWo2XoLpn8alWJ8yGWoFY41v9xpEAnQ8qxMYVVzXXaEQenXtmKyzgNOBv6KKuSF795gEa
QAbGrEn0marll4cCbpQIRPP4yWxEu76xo/jhhh+t2fI327zYyYRhC7NGsQopKNZmKIoDHFP8K3q8
DS2eybjyu9+h/AZm4QCzPhjSDXR4Ku6tu8EAc2B1ndhY6Fp75h53hAokNX9DaLq1kdPdHem+QBD/
VgVnwkGV2KPaIWoHdiaTgnUcGZf01YkQzb0HL+MbLdrO+XywAhOkko+HWWYhTLZdzlNNrPsD8h7n
K4W2OMpGIHd6xOCWC+v9iDZHr7RPqvR5JscyoNcrrRcQ2bwUfNXYt5FxU9zvyg8xIbZP7USXL+Qe
64BFmSEmbyoRNGyN6tiM6nXQDVBSpcckQuT/4nLtMZ1C90fn1VeugpyXKutbhxfzUpRneFAB2acy
fFSpVtY+TyD/7/an50YsfU/LqBN5WhwVOdYoTNbP7M/7FBqGxEYzvHpiVv8/Q4nfniM0e1bWk6Mq
9CCMOk8vwPWParJ3XaImHjN4sT509CSlt+zLHljTRljJJiJRtj5lWgIujzp9BoX7HsDfa+k3TSm4
Dexn9q4JT6aOnFKHLagZTKPSf8doLRLPdoMUGEb6rPsNbzC1+qqXbQ/NarC8Fz+jx4V24n1tn/4P
RsXn+42g23vEYtdhJ8D6d5Sd0zmQ9gWqeH2VF71j34QcaMU5wfst6I2Tk3V9dDvTCWl8YjfWa7d5
g7SYD0pY5UUZ6VqVt72YbvnjxT3tgJZzz/nwkvpktz/Olf7le0iYQ/qQXQFLivC/2h0oAbsHpas+
EOUIUpszVpoo4spUTdY8hJLJrI1qPHaVgkxHQUwtTjGROJePbp0TNoa8YV0YE8TjTJ4m2gJ6SiXb
8Vht5asBplBOgElZT0/jvgW07vL9AEU9QhdiUYbxC9SmFWXdQgxWvN1RfHe2CvBlUP23yZwxjTfy
yJRwE+rGF/pNRgD2aixZyKoMHmCaeNVaF/wbZW+9WQhAqwEfbdqeR71mI52F9lBkpswHcCK15H5s
Z2hI8EjVNgumRgE2+0VCHSa7k3zSf820WhGIwsks41gpboll/AatwNVvcBDCLtylnR3ES56NGIgM
DzJht3TNkikMSCsEHr4L8b94z0Y3Y4j7fio7xX/Gmv3H55U5V9QTMRw+uk/YKWG3oVzyZNR/51gB
WDCpiJI+5rjKfKM8oI/VQvkecKXbQYaDnLXR4UwZ1pW1jFFyrBxtlh56KmDl9vVJlH1t5yFlVcaZ
pZIl4LGUUqnSMSlbxB8Xx0nutGM+2gn0oNmjuTsjNjOzHhnzNdyYlVdnBgcROmR5zrQGguccXKey
yjovVbn7YhU1/48pgYlGGOI5+CIimhpkxc3Dm0RTlJYZopN0HcWGlhB9iqV4yl4LFj6OegOKvsGX
lwBNu5KaMxdW4k26uvEgcD66phXDvgSTRuGWR7Ahg2OQJNzaDuA+eaFGqztoy1fN47oEueeth8fb
9xtaaiG3zK5eOnTYTG1tPtE5PdnniQ/ydob0eLK+IRIF+Mn2gfnjLJWaFfrn29rmGTSlPQV5GTZ+
144Svkn1CECWK45q7o1zjugJFWEU/BQlCuFrMlXB4IA8nwavf7+JJKdsaiL+h6tUTl9ExaEas1wf
cVCuq8hQLiOhWYTYqNasV6kJCVy5VmlOZMR0tgPYxnikvOBn31h5L0CW/SeZpa/mWPTLMsIgxJTB
Pj6VlNaC/OCxmt5XOww5+RDIDamZBS9qIYpq0UAoNviZCwIInczaP0Hm9RUA2GttdKLkdYnCu9tW
Dt66SPHZblvD11Ln+JdjD7ebImxcc3ITu/VmGUGVdaD0xdsf0LjVcMoftWcO32dsnrB+5yzxyzQd
bc46tW8vRr6mKGVrHmHeAWbTsHgV17LlnX0KhH/2qpUC0clNLssNyfb3aGUtfrSGqppIB7bggc9I
X57sKCQOrW3zIZ8p3RElXOGZ2rpmFhyvu3EYdYP8VZ3tcpjdymdt9i80+T5J37CfIv8aTofrJHgM
VSLDvURwCovaevA0PJnMQIip7NBnCdG7BxC2lE7ySqSgDljECV5XRfpV3K5B9oV1QTeObVNZcFc3
9OR0vm1esjzeTj66d1DuN1n2z+kpkKWTDMo6bqIPwF1Sf1F0g2Y9uTS6G6p99eX4iAuG410Yxtmk
8U0lyQJYORwmE1e2RkE1fh1REqYPHi5qtX0EZYOSgdvxBhBLWPf/t+B570pzm5MA4xPRbz5Cifh3
ARX1qgo2yAyGxpLtmNmQJYD1lgKx0I25GWmg39hzkwKWYVgGO+0LgCvc4MNqTBdLJW6D7fBnd6By
8EWbn4SDV5e59NaJHiz46heRs9m0+qbWBfLsUrx7shK5o7Jn10nxpTXMQvXYvS7goZhMD+o2D/u+
4cWiYiEI3KKH0AD4nqq9EpdmQl4A9g3v2N0lR2xnPF+Em//6SpJ/MWoDeOtSa8EUli3PEJQSZrKg
U/BF1HrbpPUXlIMPGy3pt1wAss/Wq86A+r/po7rMgZdFsNN/GAZDO4uh5lhx5TbPqJtHguOoPRYW
19hTt1FRkhKSxJ7DLAj3gmYkr4mcuDnvgh3DqHXVn5eaC0W5tokwtJnNp74VJYbJcS16lRbg+b+P
VvrKK1sNbxfADC+35iamI0JwzUQR9BYNZPFLz2qNsupNIjDrdMOxFPAj2vHc8Y0evma7jau0UgJO
5Gtpk5sZUXm9XIl9OEF5OX0ZuwUChHc3XGwgQI+IMMvOUSRlRKu32OHMLU6lNwwBrEg6wCuVnjva
yQilw0KwKEoUccl9LWEXbpc6a7Chd3NX53ulqMu69iPjBJ4LpEwINKzCZs78bzL5PFZXoAdAoEIn
MXpc/cG1zxlsm0OypTnxmPrkVYDL6AY9OVLvw0Ok5XDs4btKTLzEqyEdC2R9YN0BAeCxzuLAzCBj
xKCzgXVEYNjeoBz3yS5S+ahv0ciKSR1Vb1QXqVDmorfulaBKSbO4i9Pym7K069kkrzMo/tE+/ke0
frTByTsloUn9avYBIcoa8W7kBMaVICFtgvbMaB/CATPId169niwrQEZCRvCgTyuQDGmHmhvcuH/l
wBsTRvA9V091vcKT9sJRhn9H+H9cBJWou89AIsdhkHDPQrx5ObnMJJ3SB72P95g9dmL5zd56zyON
xe97WZxCHL4CEIUebPAY9gnI45b3VFY9DROe8jt6XxlOkluLrUYeHVmuu8MkXpaUV1EUqnyGNnnP
XLaj/AujvUQJuT9qeNKhj66JNfSQN6nR4vc1DgzFC7fRH92qLaQbtx2TguZON6BgNStQfT7Qo9mu
PNFue5k6l9b1pYEq7RBu+UUsjjoNdvZAo3ZrvIyHNg3+rxp7D0Nm765CKyGr9jJVo7Qw2BxUicEy
gcTvhRtA1u9ZvMtuiAyJrQbCTkgFp/oVXC9og2r2cd8eRmtxO5WC42hC19MQYYxqzArY0b2cNXJL
omiPZOa+Uxu7apyeeHK8/Re3vu8KB2qwhvYHMSAtZIBteDN0XkFV/KYe1Pq/JWyRVoTzCCgR/ouv
sJVfNlddpZ7pEUWpVr29E9E8UDh0iYErQBLHIkLdL4rvpn0cY/sgmA25keRDKfO/UqojI42n6wqZ
ECcqP2XFgJo43COITGn1hi8pmr2FSGvL8hktvxFjraqPqx6LUk/VUkfrWOM/jfhgSHWcSA5AKjgW
S7FNKYOHEZrZRqg1u9NXORetocokNPV1xe3ZuJRXiTHJHg3uk3HP3oIamej+2uow54kNdVa5bm57
0N//b9xHMrrkoEMaADtFjCpS9Gz+fP3skBOgdYegcxeLEscPsPrSh35yk/mHUwYFPZmO7gBWx1xf
KQke/oaXM9IpZxebEyrekDZ+3bL/8NGLWDuAUqDMniT5QfXBC/nb4bnhOcQ89jkcm7LDx5OpmFWW
dG38C+bkQth+chVHTeA9FHjlhEjOIN/dca2gJ82LDr2q5tssZTw/kqzDaPjJVMAVRIfaiFhEePTG
w+gHV9ue575I7smagywjugvGhkElToBD/nvsbj8IHdY3rq+STTP33Rd59gHiRWZLCBmWWwOR79ky
5J82pwcXt6U82M0MhRJviV6j7xq3ibRrIRul+X2LS8pkcpyLemCe+lz5F/7kVMJmdjyqSJQDItsq
NWKgQnXQBwe053shMKvgJIeEz8lfg2GEn9vmvHsxs6HL5VROG98RGyVrwGQA9Uq7a/wje/6Im9d9
B0p5wrpCrGSUL6AQWooKbViySROVEAtQai05oRGHUVlljdhbMVYZG4WCIsXsGslpkGGMIkJ2lNbS
2mDqyIYh6lbNJXOvrAUZHGXe5oSl7fSAttDMB5OEaHH3b5o9+m5oZ422RJ+GpMAb9HfUwmMjLgnM
l5AmZcO2/d87Gs9maSUK9mG7tDIIrKT85VldeJAfSxvU/eLSjWXi81rUboXN5hQ3JPXnt7xof+iJ
f3JC+nezObYluGD9HTF+rZAe0X+dwB+g6tNSuj/wWjaiqUUc6hH9XgdmFIsko2WgmegdJTveVUXD
LEwVFke4M3w9UyKm9ZgRyu/+bitNWN504tX+aeWKdPhfvpqBafG/qjeUkROmoIU2oFISc95s7LPU
qAkPp8zCSCOgqaK1X3DXzEGTlXmFJ7lzBiETocDl7jO7nWnCNMIP1ypTadWkxHBhrGmxr0V07NOc
+5Q7Ug6cXBa0Qq92y/llo8ddaiJNBPUO+fZ+Ehk7a7sopBgv09RgYBfrL3MgbYeXL8a0OUM5k5D4
NpGOvDzcVImjcF4XsxAWUy0+qdfEb2nTzZd5CTef05ix05//MpBMj34QUo5qK5w0QACp6HQVpwDJ
IMmYQ3qi4Lo0ShZS123kWHt4LbFY3ochQXRXacWze78SA9bf7QSEFU8+o+cg0t72zmTDW/7s8MEm
dkc2+/lNqcsb4YwSawKP32hIP8YYAQfH9eUymIDYqzKdD5HY4rrasrUx8d49MilHAqGIBlNx0vKx
tXuH1Ho5+BumMiYR1qgON4mZ5DK2dNxU8K/T7bRjPNR0e/WqYz6OqAH42ViS4YMBGf1+RIArj1l1
/cyduIEfpV2zQHLN4jJoAQ5L0+zd9MYmb6INDoI6xqayTH1dG1OIq3eq/XR9aANJ28A1dEhesdCh
mux/G8hYooPPRxT8MMwLKRcwe9VymvMKH0ZjonBcE/aEucISpmBhY828xLFqjj16G1nERW4BON49
49yCauZJzegBF+q6ObtLlobL+N0f0mEgMvxMSSw48NMIovWduPEDRje/uW25phvIsw5EAVi4PEDP
yDtE8X8am38mjS8mhq3nhgiYCDhqQvH5vYr6tcTzmn7dYR8TAqgPTqiMLDbk5GBz1yyrZctXb9PS
TGmqztZozfFcudG2/l/klE7oCY5OhfliAF37Tb1wkKDWflllnS+A+/6UsafIz8wjN8gvV2ifE1ww
BMjLqWcrp3Z4Fqhf9GAmN88cmlBMUneKeE6JK67tNdUfjZOioaI3zqhSpPONws9IUcHfjEAuMP5l
s6z+C39qCR2/sCrTMuv8qtU3VXy/HoJn8NG2HzRrxpu2j/davb6oqxK1Rw9+CMwkAgy5E8RbvhXE
5Z5aYKePN49gR+jxwfRrQNoMJwi+Fpk+vE4jorB0RQvXkhiUjHX8l3fWF1pEaej2tgJIoWak/YmJ
h3LdMGzMwKDeHIdmweQW7plv/JOfdUoPS5NvD67ee1722CpaJYPINbfZWAm1CxpS7+n5bonKiZXD
rqJbwuTtDq8jASiWuKpBPaDKM6I6wOR5uTFhM3anvzKjzj8MVjJByKHM6amdDjwSfhmmXbQcTNGz
DwlPa+waxW1JJm5VnnGwcs9Su/oZXgT5tX0+zQAy0dY44bLHMN6Sc2ItAGtjkMhxfvrkR3zxAQ8x
jCUQHexa2pi6hOUaNq4u0tnGNU+GlJkT2Zvcas9JGVDsisr7rtKjMM/UmeFlyemznMlBoNS/FPHH
uOEXrcn+JX1dycRQTSjZ40A4hpHYI0nGxW6ubvfpQevUisjr5PSFDSOz7YsNSvKMubYoGuD9kT+y
StLXTsA8WwMRHbCOpQCQVr+FcEBmS9Vj0j9Yy7B/dtBLznWhvdqmStzlaw2+vM0l6bLx2tfc41DI
uwNJUNqfc9ifuYFT8PCb0CPEcpUyLRt+72PtS97z0RYoEFHaP4I/yhCHyxSGXe2d6VWM6skioTsz
Tig7q1/7Pt1wHVLYkDmDAg+CG9n7DMWk2Kk7+7zCIB0Z1SZm8JSe7e+mZ9o1LNm78V2zG7HbZsbN
x7+VnYL35d3XpX3gVuAFR3H2HFPt0WQeseMh4/B3GhUDQlzHSW0hAtAulZ1OQnlEH454hVmJC0Rt
OXla4eH4k3E3jJ5+qTNA5JLe5wcLP+JnANPT51UcNUElBVCLtVM0eyj51oAXKTVSHX/5f0XTEFNk
g6L/snZABuB3hOr0hC+klCXPVwxEJVodjE7BInrgCMbpp78xROF6wvNOT7FLOKILQYZB/xcJ3qPX
kxKmQN9fBeYYy8YMefTcdfJqVnhLhT4Qrv563wX+pOAZf5IDbxN7qB+bB4a1WzLc3xYviIzHUq4j
L/124kb/TuF5qA5sbAPDcF8ydWmMmli+sqoQCI5cKKYaZpMTYTLJhbnZ3MG3xWwI/1veMptm22mC
HUmDSRsFIc2WBatDraIrPYv3Ses9IiO0P1+ou2HUlS4PPgDTrpzSjKRZ7qC60BsYHJC+ZaDu0W+1
OEQUJ71giEmnORER7NVYnvc/+tQCrqVHF3mOLgZ8rnjxt5vBfJ2Eb7XVZQcGa7Un+wFw12Vqpldk
dtdNVnDmhdr9JvxD5/MezHFqfd5RpYhAr8pDnjj+ArzqaoPYFlMxOSjRHuyM7ITCh+/g6DXYXFhY
BAeUj89eCG0LEBX5v2mzoRsAtiqMsdRMiYfMu1kp6MxhcxK52urxB8NTOfnENQ+PaX7X/VH7erqT
9awUiRnwP8FcxT5l9nMP22rgLLtw8BxvjtrczAkd1u3ksVBsSp0hjX3IACdGOfEVp6WVtLU4WRVg
bUzZkLqBBVXVitSXbQ25cQ7NL4FWUFviEZQWNHMXWaIjVI+8OGuwtGKxxuBZY4qLTCOrqqkzeJX5
5sUzQUVgp+dZVve+1H62idQT4+K1S1RMJ3Plul3FG2Ew+LZht59FzFEPIe90QkcCNTo0aZtmfeHV
8njEYid3hCWY9F5w8uHziX1YPVuOkCyd3JP3UFod+D9k8lS10osyU0akbLLQQyY4ASN2khdNP5YC
Kjzyq6cTYV4DN7U62BCTzb7uCmexguLqYfFYUTArGpydlQWcuFp6FoUbIYvYzzJD0mOqH+DY9gBx
Ts0oG/tMCussdEK7OWwKgQae/sjk38onDOC8J5vYGc0w2nSph42c+68y8W3f8Z7ztzbSWK5Ckzk8
GyI2nUvwQCK+CoHsKh+I0yakZLA5GJ1IwrTtJ9Zloy9TrDCGFib4W3Tdxz4gOmCAS5H+2nBntHpn
DdaRgwy8VOdFo9ydXpzpgjBwmgrKRes85BqgcQ47tiSbjzJxhff65uWcqjy3r3r8w6AzFxr+CdlJ
xLO1PUcMEBV9drZ8VdwALgC2lbABfACfzrGYovPs7XBR2d2zQ/fmpBD+hu+IoZ4tf7DciiY+MUyJ
aXgxWT4fZTtt6+Q/6VSiH7A/cR5MBhVEyjXAIwRCX/aR7Y0csogj7jlz7Rs63dqarbp7Y8Aogss2
VA6WaboLSTD2xI8fk9PHVAJVq0S+oXHNybekfbv7Z36twwctIk9p/kc//knJjGcqWuacTteLhKS7
c2OTWheq84/kFJMniVDkLSnVZWiXt+ixlbIynmWare3foAfHgfO3p1+NfXlTXv6eZf+YfCYu8ReO
B/XbXHDP0ckhSqVP9CTgPVKSTXgFR55Un90GpafelIoea4YfWM96QjBcXNgDojvD55eIG852heTq
riVdod0gw/fI3ympOWHjUhB6toUPpo2AVxbnWP7dWnSpXYMN70GyfrZ6r0HEgWKimaxSw30TPPrH
2B7HaLGvw8ngDM7KzJP2pbMG2p1TfPmKiS/Jv+zQOTHi93I7VsK6P1IRAmy2N4M5EqwBXreFxYzI
0dEKTVug/NSThkYOHAeSJ223HoSkr3XpZdxhKyydKYD+PmI9T2hIGiaoYePkWa3TVWXIGX3G2yZ3
lyVK/gHUjdIFrUbjsSe62HvMKKliAGS/2LTvzxvHwQfh56lpoNuCm6f9zxhHKKEbNt8NHqzXQZ9l
fNLGJLT0RQZHRHP+yk3sOeVE46AiL9zHgbH++u+0s0fH9sXcp+P+fYjaRR6UOzeNP60ZpvJ9sHKe
0YzFqvvkRTj/1/1ysNQegylSNpHyRsTnMNT0xYz4CNRYLruhooCgBiXE4a86zFqXh6jXy+P3UkeE
wjajyk/LHcVqVnSPSa3mkSSCIzLj6Ks7FAb5OOdmoTtElRH3oOjHpPkMmfxFDwc0ad/hxs0Uc8Xz
o58KICT42QqHzCX521tZkaDqK2inTqovhiZXNVMSJQMPtVr4C8qtVvFMCi8A6DSXclq/phm59CZU
YcuCREg3xb4IovEqx8rKCD5LLlHOr7ObeDdNIwo7tdjI0Dv+R5YGfBww1ci4nne6BTUUSO9649rN
lAB9TylYKy9BYlrNAYy8zs/AOkqG1Wmz2oYfmdfg3p6259835YrFtt2k7DILSI0jAzdwqw3489zD
N1rhiHffi/RqgGIkwyQNK6NipxuJ9jLRX1JOSXH5CfkSquPfhA+xqLL6/OcpgML+93booYfnBxtm
3tUllkk5HUDggKctwX8Awoc49TQz101euXfNNM54f2ZF5J7jPmxSPzryGL5iNWaTHwt2M+Mjbsf9
DpiSyNdslIooEMspqf0x5dTH6Om13kcKNogyYIit3V1ysIL30r4jZ8ty3JuwVD+pUcPAF2zvIU+g
iWT2cGhWepJebo9fRuthK18wDvA2ocXwozvzdSPHa6gu+I2oXFSsQzgv2r0b6yzfldpX300YRH0f
wuyQJRKsHGsIn9Xhy7VQYk5zIc54C44QDF7m2KCn4nsRUcM0FHGYzW6F7j/kJZ4QuCHKUeqe52HC
k/kHhXne48F37bYHUVv+EovsgzMCN4V5bM56xFzc5sjc3iZ0decS0LYejOP/Nf6kGAmDCSvobQo5
bcPF43CGF2xcVxEkyGRo8GXSxxCGd9mI79dud7U/Z5bHmVmmEAUrnch/nFhzU86tPa51vqZmF0Ul
liOc5s1C8GpG6oMppkMgovsjaGoIpXETn8Iucemuoe7Hta0tfJruL3Wmhs9JZpkASufXUbU00dvr
RI9XHazyt85TnDmeGNleRzo6DXgtUSfr3DcYUCocjHwGEbU9pdt3reMof2X8Goqz3mKkKFnLc4NJ
73GdMneZCHOVJkmNWLdCak0nwOOABL/8LW0GBpggOLpfHVdCF3+UzusiASaNoGSbTUBNXNsK/LIr
nl+wuMV4jNldSdY4W7i78IgsxK6hzVReofj/RXgPYy9Nl66rZFyAYSmaq7LhKj+hvW3JHpE7ZLV8
xDYcZMLasilIQ2btQuoPuh0tuCC88XmBkSgVTqcm92/Nfl76gujtNJwlNPrLp2uVesqO0pv158JH
19rBB9pSFdSBMfXFMLLRBciEROkPXvvFEh09lm0fJJEcODCUlF6SvX9h/ECfP6N95vEm31GTKovy
JhVUPmCOaiI3PvR97yF6VhV+PC0+uiRxkUfDSPA2rUSaPWUT+V1/j8LRxaBYeqFmdgFq2pYSJpaa
40lL379ESzaBlOogi3/wJCnbFa2SY40f8lfWu57s7RQ+8SMtTUOvzIvuW15l3ntIK7PAggTCmhnX
dS59CXw7YImhNqOmcMw7Ca0Lh2RMHOgHXj8IyAhLm9ZJbFFigZx5XqcxRQBGLwFkMh5+gB6OYdcm
GlUyXs50xI0EVbE+A21GtgQw0qDy9CQj4o5aRlLAzgE5HCQlurwBho/VSby0fvVZyHjAjqpZPmQy
AgKs+WOH9M9b4y9vGesWpwC2BKOv3eTvoGYqxccFgB5xFiVIT9/X8rcRsF5A6z/TZlaW6JmCp4MD
i+n5zrROELqSlxkZkDiIHWNLDTRIsKt1Epgj4+edwy+F/TfEabf9rizyBabpezjYBlwhbjd+zDDN
3QsioCt1LE3MJ022IIkgTqB1+N3xDyh4lSmjK4ftpVQuMVNaMfAg6rSdOs/juF6+8rdBTDSM/MGG
xt6nR02Vp+IeLc1OB6BT8tMKmCEH573LttVidpiHu5eZDVRo1FFocs9IV/0bgLEviWND92lLEuEB
vjL+MqDzvMKua/wuWRqGcSvOY/M816SqhNlzyr76GJyv0g8pmVxSXPzLMadFVTI/o8JrS4vee+x9
JiilgVKNB0Chdd4R3l2rEueFrBE8wxnWDdWgCyJmvqHLmTqkrFWkBlTHWloUUV8MvvmRFqPvpj6d
2vE2e5Y6sPxUSoJjRgkRmGh5XXN6YKChKn1mhapJav29WypnRiNfHLkrF9EoAdLDZoF8bZdm2RWx
9UCwmEKBYnJN6bGk1KXGtioxsvpfqimo95+O0BcukcbZdrts6pO2D3AYGyeHZMhebV38EGxFL1Rj
PLCOoNmRfsqP2drqUdL8VuJ/9EUNJqoHBKQITuWRxMU/m1JkKqr6dK03w+UPErmkNmn+SURrkXLU
FO81eDi53X4AmHR4MKDfctR08sRh4Ji66EscMQ7iOWtiWMosjTNVCB4Kg9QXeeN22ZeRy/tR8UgQ
rfES356WSW6oMu+eXWq8GNbIBy1+9fBLF8QpxBzwn47mAw/M9/n88Wfi8KwKD8osYJbIzwdmaDGD
SVOtBS5Ne+PQu1aqMREPHtAPhPBKaHo5GsNlXwt4sqBdixdRHtVO9fSl+5U51s4MrPujh4qf5aIn
SswufYnP0WZkSOA1b6IBlxbxnm8JsJH+zy/DnHEdpvpRG9kWvQRZJZWXi8+f8drgnq19GHKYdxDd
UsFQn6XaVC2uS0xIuN+SU+E9AZrtG/nzOffHrRLefE5R7jUBA68Y5aKuB9DrUObBwR11u5qBTdKe
GloST4sxmSqdoGXpZ3YsQsFwbVPSh88yv6g+wfcEn14EI1RT/aH2GHY4jfxuPCXsbYDqJNAmStTd
LT8gKIOTkuGRUF0pARYzGKARmxa3kinTXai9d7ktthX4NBeLoLs0vHtuR1mduipa2nSATSe77RNK
sAv6s1t1db4sx90TkVtSmN/SCErVk7GhW5/X9Z+87ncO6HIUWh7zk1+EDaqNV3Qq8KlpiwRUh1DO
w2qvVaziVVbYTi+MKCdtohIKrmnXahEEst0iffsSJmomaaMVfdpSFhY9pc6ihA8M8eFMU/O6tKI3
XQ7ZRALkniDpmznDkG8mXiV6FldLio344uYkfkAtINYs20dPv7v6zgB0dgTAXOCV+gW5HCTIr+nr
efKyzOibdbiNqhXoWaSFw/LANtiUTd/FKRrVXE0Pex0HdJUKvDCnZDyRm9NdLq6fS93s8+p0Ebbq
mM8P4DP8jvOY6zXvpc0lYyN7vmbL6XAme5M2KRmD0FGxtFadR9VIm0gOYBKyZVNdvnFeNOJt/em3
EhhSPqHcIYEk6ePypPRh0PZC+Tcafx3Mtr+LmHEhGsBAg6DGf1kVGIWprwhIFAj/rK0x7nISI8Mm
aLzVVyFpUvs7I8LBVBUIT2a9CGwVP2d8KHKZynGN+jEIlOtA2dVhlAoLQ5RMIyV75q3iX6YMR2+6
TX/R0A5xYh5n48p2TScCVsrZ5BG0E6ecQmFf807OcCDx+ZTkFe0B/PIaVHDOBufHQ3qy7wA93QT7
diUK8/WQzqVhfndhBmtuluP3NHdK8rFZBaHU3OwVrgEZ+CsgwtFGBpviK2szByZ2kPbWoXYZDlod
nsnke0hsQJWg5E93prLbmePxfEj2rosO7pqUNI2UalDdnTkgaOsQurZuyEF37PE8aNuUk7Ub0JLS
JTckSe7AiMcFxSsT0MwTtMWTxxxVS9Lu9DmOlrLmRjOZWmKxZi/94S44nZKZV0h340q61zR9Ghbh
4rKxrpqYXO2t45ibk0fBFtfi4HfH4exvcFexF40IKIRFzkyB0DoB/nCGbNIUHCq7PFtCofSpvw/S
Q16v+vOlqyhaMurphEjW77qGMGbFCRqIXXjnuTmZjwzQ7B98oJUdd4CHtsM49RSjqjhIp1WQUYZF
RgnK2zti5W2qm+I+RWFqF6CUj5SjhRoSWZ+Qs/7VQPi7n5KWdouMAwTfBJ44klt8Zsp0TwlO4avT
f2HZmOvybxIgsOGu5fiBXeFdFLtt+hzWlD/oOtPFs+Jm/twegKWSzpfeLrAMOSQj+9L5mZajR4tN
nZDW1xButMk71R/wHG3kvPVcMB1liB7QvGkVi5uLPI//RPpqLNw0sHNp/FQoP99s+IuXI8t1dBoV
Mh6jIjNRimWkUAVQ73ftwgc0XPnFKLOymmsRrzVM01kPB/I0bUkcQ2hi2BDRIDnYfEu/68GnGRBj
F2FWbYa55wIlyp+WOSWyujcDNOpfzvuLm5kU0QE2baRxbRqjo/pReFLA31Vly3VXGb1awaFAUtGv
CehJgKiWNzEcmBuzmoywTCO6YRhdJwbz9KQeqyEqAtBtYAQJ40WKjazqu20mEnFv7gcr3cP3xtc3
zafrssqm56HOpa7py7YgOjawIceNv4e81QM4ClMgXuVPEgDvwfhIFoigcWHgvhCobUutFv1iugmE
1JdI6EG+uMHSIBgbQ1fVsBgEzEKj1RX5XEgu+gV8k8R8UxwhUTQtITuVs+loYtVq3USW0ilr52m5
WQQQ/vHXR6HZeI0qVV3rMMHF9P1O1XmhWgihTqjKG68difurz8mdq3edSCWYZtnKc7XKqGSHBcR8
TDl8Wb1OcIXAIxHm5l2beXsKBWHD1EMLfgSKCKVJzDCsQHAoYvKSvSxNUJ4HsBHg1Z645ymAcZeT
hDxxYee2R0sw3nLeOVVilgopnN5PZjPn7D5obNHHw5Ga0H/FxMWL4QcgUAunxesPn80MM+i/Di4j
QoEtifdoxuXvTK0n15Npb9GmLx5DIfk7Zt37LoOAmDaPThpQGngsNT/in+QigJ281PRcHfz6Qxfz
06Epk1U7gLxkQzfAaIAstxQCM/wvzReWUF6pXUJfb1fazKdDCkZopXuPjPn+Jdq/JnwKMIUsVEA2
Kg8TWgfw+HE6LQZLiGD6s11czSsVpVzTnesaS2KbVhzUDRA+jXgdtSmiA2B4mvi9oEzUeHlJQh7U
IY8lbLoQqP21akG6kVIcqmj4Yy5e38mnaoTCjpCvLGr/dwxZiEeAVcBwTPG3LoA+2efYHdUCvAm1
7u1f0kd43BbRiP1nAYTOyMqw+jTR3lenQeBQc26x9eam3BCZSwpMz7e7i2BDE8HRHpVFTacfLLKv
LSVOaOhu2+U1qJpBAmXUqYSEIzke8/8L9J+Nh29RmiyB8RXIpYzCwq1+GXph+zi0nHOnUZScd10P
gJDdzbLGMMiGNbujLL1n7cuEf2fy7gsT4ngwgQI6zTy5rRt0fGf/pTh5iROcfBqw8RiJ6jKmhHeC
0hgR0ndBtWK5+nAktqIioOhfjkcqw3t0DKQrH9GvRjQx11PrqDV8A2VxA0vMS/830/SbnlNpzOfH
XfJrM2HEnm8eiPBoW+KR2MAvzcp7TDET/UkT8He6goLIldEBuhAQ5iu/IPJlyRUUlBAYxP3VFZls
jAl7gdOojN8jaPTK7KymhR16kdh82GXjNjyR866XiDljq1f+tJX5ttYHPh+OvYvpSXqlFgFobanB
1MqcryX/pobhmMyfMl0WaekykIfFCj8aaKQI3+sn/GD8CqHqQdq2e8i2bLFuuGkQmlX3ln5Wuk+Q
jTPrWWPDt4ryMJH3jZJLvuDLDjXBCbm0tDDQQQ0/4jkh4GExYzf2z8r78evnRz3MrUiFT3iaQycJ
6/MJb8QczMYt19D+14ILZyjAYTT1L00kOZiSx78n/9RX+ZZZk5YOxf/bYGUjwgVt3UZHyIwX+t5S
6fkdB7OczAI1Yqsj1mdHiqI0zewEFL6X3VCZ3JbVIJMxEsoQyScJulymaUWEnCIWsK7W8o3/dD2y
qf7tB7g4oYpCU/xZ2LBv7r0EzXfE3Vzl6ik4DUSqHyDxOf2URThYJLyRnND8pXpZl/Ckb2w5Fywv
2A7e+iGFyQJKtNEhdS8xPV6BO554D/9B+soASNvcHJ0D7KyJrt29NHMHbL3rGEc3MrTkdaho/DSD
ExrUoLlVWXrGCPYxdbqIe+xNjnZZ22XrHKyR8GqbALN6KKM6zxPaWqB3+mPKTgEqt6r9Pms04m1j
MOf4v5fp2E/AVJ3ZsjsTjQjsAzZN+vzNlRbVPMQxnGNiZWYipxa+fSb4tA8SeLeYvhJpH+4gZa3Y
qFcbsfpEcHka+xkfcV6UmwSOQiDFPlKqAx0oD+4oujcEOAAl8i2MNauoU/WJ/tIieX3FxgbOKvI1
bnQaZ+meAF5CCd7BQxh45krMdePC1ftn9Le+6DtbO1lruSCiETzBzOMs1jfRa1Gr53ztXadXMJxG
zPeL3DJf9bspNwUHOVSm4hyrCnBQv8yLa2eO3m98QTmz6kQKsWT7Hk5GE6yqPR8m+6yyJhwcOx4j
ngaBDqT++EV62t8Ms5Q8dpqNQuEHqME2RR5ooUsW2kbaNASvk/O8VsN3cxzgHVIfdiWBDhQGIQWe
EJYe7KR8IJEuNfKhsJU+IULlLg1lAKZXEuGpaR6uLb/+JIM36b0/8WTfbMNPoCO9THh+O+8Rf9r5
vJwh9h8AJ+t4sEBMSSxAkBHb/d4QP32p1T9RFgdXvaTnq8j6JUaJ2EzMKzcOgjTwM7USj76RIlgD
hvkZcLiE4uV8PpxldSIP1rGCYmEOlZvjZmuATeQBJjyh6kwOgwX6T6yVxQgwsisBlseiM4hLzIRs
ZRz9qXCeOdb18TpCHhnEzc8SY1hjpsH44WR8Y0LUDw4ZG5QG6Ksn0y7nbohiMbgfUNdZMhBi5nLB
gB1gntUJFa8jTh1YIXuoRjiWb11OmMIf9n27AgKrZkJnZngSLU9xucHXpXmn3MoYiPsaMDW2s00D
4dCQLp5qZ2lZzPT9v1jnfZ1OjTYAPgRSa9U9j6CHXgsfi5ZB2G4MRienwJU8ldDV9yAJ6u2f8kC7
1IiCB74qRLDH1AadHFUzqGUz3J3ZV3MK529TSAP0+CuT7fSPABDEYGNf9dZKGwf66dMWeVenQild
RNYGbDwmXKGjXK813aZKGtu0GIyU0hT6t5kMjXJrqlhCdsk3I5ylt8m+GIr869xMH0NOUmzJm7S8
iv0q5R72kT9IU6MG3i+UlomDUA6/HGUHpc5+dT57awmNaSgwR2YLjFVFV18bA18P+b1s+quF75KU
YHEKnTU85UmesKWUX1i0j5olzQUGIkBAuNU+0LXtwmeTti1rdPeAESr0ldszZOSBru3CUVfSIVY1
ZRTzF9ZoTumVLI8gZkbR9KkpegJ8Pl6y683GL3vC3+1UYUSd7DNYfTbiv9oiJLTUvHp1NqkLs+ob
VSSl2UDsC54Q9UDu3XG4fmdz28pcSY1EmjbjO6sCPNVw7BZOUYpqkmvGINZacLxldaMQ/qik5ItY
6TbydEq/b9AnSaNMwAlq0GK2481HrzR17lGtLCDykx1w+5MTwkQc72TiHluS11O8N3B4b8T/9bVu
/v71IRyzisPw4Ve5qAOGRQaweWPyA5wawekDS0CRRjFkaVg9YiXARjIEDLqYOjoAq7Md+2A0O345
hV7poqOQMRbyccjIOThISwqCDfgRFt1grqnwmLUqBIgZJMkZGR/su7KKMMe4+FjiErwvebNB3M0S
ujesEeXB0f32o15jEspUxdWB0VIgYz3NLRANEXiJa5VufGaeBQ+uZw7tRNAlBr6bIBFIZIznPqZN
7sFpJPdJq/E4FSc9pyuDUk6W5cdZs2a6d09FWftuSeqrZpWRpKm+Ufu+LG9PPB+1yCvZ53Skbcm4
o6ZYRFhCJ/UNK5sIV5L8qGriJJCtP6Q5v6VisU7P6n9XfjfmXxED35IXqZsLlN0W3N23cij+pqBO
z9sld05ZrWNvabsOIoQlCHa9t6lHZ4ZPU6Tc2KvCNcuS1eO66IMembj5BUP8EO/N4C/pX0u6fIzX
p0EjTsLQDYTy6pjzW/6+PgOnHeXrLJX3xH/vvFx7zKYhwf035pWoSSLAkkEtLPGD2tb+T2zFQJQg
fjL/Kv/JqT/dA9f54dj2tMZA++sFtYoJNJ3JtPYKwdSyHw8UcQy3mMrg687NPhDN2Hyyw22IRQw5
G6umrEvLB7wgaQaweZOx3yRS044SgPTzePhldQwhPzS/wBKW4k9dpb2VNGXqzR2AzbxDQqiRULpo
HBcDsntpLxDRngmsMYgIW5AFdq6E4ZvMVkYnoUblgKk8oRuLy+C0+vayYpMH+P/NKbtSbKXjU2KK
Bnc62qgb0cfTCKZ1danadHoYZks7ToiBdLv4bC2YMhS1TDvoNxTLwpvHEu7ibCtTXf2OEb0sotre
7F2NYa4SEFgUDmA9q90l66oixKraDFJHCoHON8QWNwYe9FV5f9yp4F6p4urqfCo3/J5zHkq8gp3a
T9+LRp/DYK8tA2xVojEavIzJL2blcwG/PR+8HzIYlmd8BL0PX4TZf2qYWNtDHUYeVKzM7rFSYb8Z
/gvfbLIijCIuNe+24E4JxkEWN1QJTuhBrPeXKQQMAob78miDCOO/zT8V94CyPxLiPXQsNoEbaiFi
7BsOokxzN80NtTJpmShhbomrUYod2aeXdkbGsANgTFhKM9h6sC5tfglMvY2i+Olnm9N7Bv/+7zuo
k/EAndczjPKqAVs0TmPcdz3xoJuKgV76stBmph8sIYAZsSLheJDTOQzNEwVIGVf0UW5CwSs7ohV/
vXX5Q1lcjQTEyP3jc8JKUBikXzUhfKrxXwgjVkIMQ16lopTRBxqhcwclKCHYEFiMq1kgNF8iKJ4w
QVgDA2aOfeAjeLfUop0NlwxewS7+i2U99Xs7x3y7rbLuUsu/gi2PnvtrTKnE3P3uc734Vn8p/wfA
7FUKn4DrVLY1bLJyE6wGNr42hRF402BNc/SCBI4zj8fOiXJojGQzS1VEjcgaWJBEVKkviWXgNfUL
c4EWYMibbt9++4O9R1apWlrkVgI73YlPyauaMcP29n3Xk6MeIkZhrzr53QVv8myEfACY5YnLFfDP
iqQWtWofhbjyF9toPjtAm++CzUsdeC5XynBF1D2npMqXh/JYIfcT9wvSUyNGagwPshEtxE2751e1
NhQ82nh3Y2ayHbogMJMe3OCULq7dJDt1jo/Ej3mFt/G/tdL6aYLdd4gOvv1a67VZR9K6aJYdZsRm
S2TEB5CI5xJmqT/U/keYXKfUsrtn4w3NmRlQQX872c+MSNuqDSXVUvA7hOrbbnviqx7n8EU8LNRa
YZ/mSFOx7J/GMFLXWuZkekQBqGOd0BptGeWV9oG8hbJ6kq+vk9SMM+C1x9jz/nC1q9wjWCaMqV4A
U6GK7okLV2UomVruov4Nby3s50HvVqRcMWaCCHMroJm7+Ffr8VNveq7xliUCSzYRvtpYoEboNlnr
u7SBYwD4QdXmqJKUmpXkO95WIVO0M4aSCvXDBuz8CZ10lq8z4isx2jTiwiM+tpDCZWEkFq5NhL9s
jBQNHA9YHphpeGAbQco/9luuTNLh90qLelxgdRfCW8GyVyvFNyHObnPMxZX3erdKaEG1oKDb+sKJ
+XD5a1DGwUs8uFdCmsSQSmMw8ZPtsmo27P96l6u+s1y2l1QrZfCcUbMCEn9NSN3FX2+ZsxBHufGX
LPe+PaWTzJ7VAV5bPYZwCqLvc+4tkMDV9XJ8LPSUjO1YuCuGtlHWSNBXJTvFoRyowborNziU8NZU
ejaMsaNe8umGMCB+fZZ2uyO8LFWvqB2oaWs6AaoONwMFNlb45tijxiFtzrm/AWAWa92CMxabD5ME
Mqxqy8WPHKPTYiBGO3QNbfeiK+Eatf6hudsS1CVd1XN//0wfACwuq2sRar2vadzg15bGEg73kXiW
6l3MzdpqHjcVzQzZ4rKgBZVNcD5tuKBdKy3DZWokH/eFEyO6uRIUvW6MhB3Bz4JI8KUs4PFMgxlE
TfR8Q499aCCQ9vVa4Gb2wM5iHO/3MwNwIfp+oGJ7m69F63THQduPvmzH5mnsXr71p+3IXXnpJzBy
wqmNgK8maL8UWJ4DsLcUvnz/I5DovpklJ+1tFZUcLqyMo9ADOZKn8RJptnIL4TkwmsHkChuHowap
Mz3QH3wXC1Y2DMfm4wr7+7fxEy3dkB1K9ysCMznljFAhvWZAaV9HQAEJ/quQ9OukuzhjP9uDOIYT
siU3hDirs0Ch3OYHC5Z+fsWRbtm9F4GVGC1SFOiTnw/K+55/uuQRvk+wK7qKeUhpHdWbPmYj3/ab
9flZDJGFB6oiL3vw1n/MdNySaJs9XP+FyfnLfCz45mSZxvlxcK7EYXIHytEU65qnh95bd2jlHRVP
N3xQBRRaYfzK1UQaV5NrbjTRXHzSP4ZCbtuH0laTRaNt04eOM2uDV9lF3yUCnW4HzN1ME589dJtx
49fpLNoxPzwPFjo0KMt28nbT0d2Hdm+zCEK/Jxm0qyFlqIV4vydFshlaiG2IKpYz+znjilZGbOTc
hImE+acIlOnEAhZN1lPrtTjVAhYWlITAEylNRTT68/yIPEo4tFYCnOZpPoiDKl31EOq7God7yuK+
YcdHBzYRiETIOOYeui0B4AqOSFOUSDf8usptCufock6THRHujATuhEKdIQ+nEMmtu+ItOArOf78N
q/1zUDeCZHrJCiAf8Zn/oc2xAz8K6RqzZH3UBnzb4886QUBUlV7gKLSQrX6pKjGQ0QMUzyEVM13k
0FTishCGCdpD7I+xFsyf6LBFckQs1potZRiyRaRRh+/rL3DHTo5kKUHBY0rWfrUJ1HBDDcFiSYX/
f6JZrKbK9Wg/GxWGawcfDztndD59caA87JyoKTQ43NLPAteYFGC1nNQZF9MCQmhWcUIGGXmYagUU
fpx4ss7AQFiF48j9Cs/gmJtPNP1S734HqiC2OTbcRPpdnSpUJnmgKz7U6x0YamuuzaHmlFxMsJBR
LnTcz3VuxH7bY0pfe9XGuhVFv+g1s7jWuDuUrxrSt3Oc92rbMxqth1dVnp0MNaz58hYxK/Jei8Oi
FEPrBt9knoH6RMBo1S08y8Lk5/aBN1tp+uui5gCkeadR8GeoMOTq07clTic6QfOrSPgnB8zK/f6l
uDXlSmZ+gTHKAETvDXbQCFWhmkb8Rx01dvGfOyZJxa7MC9F43zjWLyQyXBIEYwEatLyDNgFIbvuS
9RM+Xyzjqm+mDH596BEVd9qpW2F+5KAhob4Xn7OyE/AKI1hRBna1Envg122wcuWbmES/Rnq+bidV
DVnlf9EOUTxBM4Mv3WjpqiZiQ42vnCan/tRtKtPmIIGo+RUoHKiKdvAxQSQmXpblSq+wwSKcpl7I
8NQm/hko2bQk2MHVanm1RFQDYMqYAgNXBurVnmU9m7Eh/qzMDphvY4ys+8ZiTOD/yQkcwEuo0i2x
jfxuaeV9QrBk9Zn2dZXzFb5B3Qpw9j2ZuUJ8ZQBJLSyhFJjlLegBVKeKEg77kxwDaaZS3U82E+Fz
d7kveaKtMngyem3d8WJqET5ruqKrzetlCnuF9TWTMufVd1/VHidCXdNal9do2ANja1FVxGO0huEd
F8b0jLLDxUhHvKf3qkpHokLnj/7OYQQczSPU5bmLX1woTI/eikjSPG7q/FgtupIB9mbRQ9mcME+y
APG2+AYE5fY3Owikylt9LeTObs+hzMy7NhAf4baVUhuVF9lrX/M0FwykrldoxXRBCqJA0y9PAJ1E
8OoBTzKdUUIYtaYiv3BWHdPbpNHPmgTvr8xz6F6bvOyxdBFE8kGTtp15APbyHw1UKmNrRnFXVBlw
SAFgtArMBpNpz0l97BigtYJhBFcPr39nJHYRKYdYaXiCwOK8PwmRyBVkDhh3wRzO/uOrXbq7LupP
SOSyxTemP1AiakGKP2kLH3xJDLkfZIBq5iuCWSm9XtIycoaDbphQKG4TxUyQVB8HykqlkfQct2MR
0tk5QXJp923TDH1Z14QqKoIBvhCLOTwEu+ZWHIUbxFQr3CMA7F+ycCxBHMg5ff5FUNniblM2XxTl
RNSj1n9Shu7pklLhtDSAluxSmvy9ntMuhajdG/fMZCx5YYuF4EnLbYxAT9D+s5MAfB6D5k1nZHNJ
14HeovS24JU81lVIv+Lbr/niakCA6yt8o/sqwaKiafUknl6RFGCYURNgycNrI5LqRwzRTyKmx339
NRHQ2tg9frlUQmR6Zzp3Yqq5NrhPc6soJH/8pA7FBmzj7wTAldoH9NryQL19wyJ65bS4oIscZ5jr
r6ya2pOA6CGIsjHg4YC862WniiY9zNGIeBbofqwzKcB1y6WH8jZ1F2aROgKDDFWj/JM/mBmoqUlM
Cx9VFod0SN+ME+Q9GnoGW5ozH61/j0iegboflk8r7kdKVMHLZ1JoxFkRB7QfhBi9qrBGMM8LQFz3
UcbcvTWOC3RPD1Oi54b9OsVfMgeMatNmgF4kIrWnmcKuYTBR2bgB6HVLaBoFi2pzWZoBIrDU9flu
1S6sZklB2aqN529gPaMcpVZAF4+Ss+DE+Qx8pvpS3DqEFBdCp+T4+cPPPYdfdHsgvhyMsQ+4BhFv
v50uhsMneMjRTs64aeNzMl6HSp33rpaQf2ZbDyf0mgv+pJ5B4v2JQoO41bBpIrJ3B/v7SjWJreHk
U1Zj/DADcohZjQmjnzITsRgLfief14RXruwLdqqOvskoZQr+IAXb6pHI6eyQMOW2v6QBnbNoP+BA
3dSzK4MCNA/Y4BDU8/uWYP7gqKMRbJaLdxEfUuiniInXEYGoGdqVpV9D/JMZuCYy9qzkWxfmC1AM
bXCFeOE1dv/6LL++eYTCHDDY5dwX8ISyk+YpGC0CwZqTumU/loS8u3M4oJmTMeZCpBuiBpUdKnXu
Ya1q74dBcWTp9kNTA6rIlmAe3We3jZsUIeqSA8NEDs9m7R/ORJWbCwy704Ezj9A79QWrZKqNggKz
AsG1+/SNbcy2PG8UoZNk6odDF2qDwxn1euTM8upUWRUGkEEX2PMnTUJbi4q7wQMTyTbdeoTOgdbS
0kZgMYGdPR41gX2bfFlXU4+wIOC8y2cd/rWaAhDSguFVzmmZy9bTVJ/JKI408hxD/6Vb4eiqYren
/zYtWGbdO/SRquBKLbMi98ziAPhMYULsq8Ab3t5sgJQGg371aWyw2WFzk9qgXIKjZ7VZMcdXmIUB
2/Ss62nADQA47bwfl0/5eC3T7m/JaBYJQx05N4QPWvy/RuNfHjE9Hz9zzeiTj6p1Du/Y53GdAiRz
xwK5EyjLVzmJF6JgVdaEoowf4xpM8YUq2NAvwUW23Lg1QrWkiINGC2r6qtFH1kP6ZrQjnaa6LPoW
qlY9cZQNauFd843lvRqHFITcow/Dz5wBFD0oyZoDipGeQj0XAAgBHb7ObEnhaMk2DLzR04YUqOgP
tJelgtV+8HVzPlJLkwJLtGFGS+ywIw0UQHeIYWlAgQK5I+wTyv0RPAuajPcDwr1ZtQSiq07BIt7b
7v66ItpJg32E/AN2+bCq69+HZeRIrjSjmjpRNz5Z6JlQ9PxKzyFFcgukQtxJrfZk2ecnvZxOE9SU
PfQUfivu53IeS6oYCgF4kxbiZmbf5aDqd8h5DQs44523nu2nhl8JxJbTpQBgRHHoG85tvY0/o3EC
NkR+v7OG/Qx/+RbmAr01J0oh+6i85vesIih5BYhgXNu8ZllutV+p67cNu8PEeAiDT7ZCX240VGpD
rJg17iyp8f2BRg2W4VRABX39a9n3oYMXtdZSlC1eTQ9BtUmU5dzqT6Zx4o1nsZ5wcU+IRSLy5iDH
JcCT8+iOCTZYMXtZfZwazTg2PbsSyKxJXKKqj2kRxtGgDFDrsg8iOKZbcGIWhiEs9wvv0PFlrkye
0N4EYDs4WrfWutXZSN1w0ohVh8ExjLCsc6fX5iaFB+4jadRjZ94f/tbS6mI4sF+KsZfUXMRxSjMK
/gkRYcDbjQEqAkw+U5w67yQiPrZWLk81VYZl6eUuxR2eYIL8ljbGxW3ac3szUZxz2+ZUhQfqySgJ
OUaIWPHIYP2cyjAx3QerJucHmu5fZVLGrbRcnKWu4ZAh95UKYru1XlJ2edH83rgKiKuVYdIqItsP
x0uBNn+V5yXoycUSvK0Lk9dl7rZLvplk9f0n9lMPmGQWEq3uEfLgGtSL1MX8kTgNPrR//rfKfqyh
UcqWZ4x/JEXMk5MLELhad0qgN+Vz14wpCcnwLF4bOXMjvKjuA5WDYzVxBS8qft/ketToJ0zgc+it
NO6oxcQ8LHxJWTHSlKo3jRR+HbyjUtG5+d/ua2NVjD/WXLB+U0dWGhWYTnby1VUMdrzeHottiq0Y
A9xeMYWfZY77AJt+Uy3DC8H3IZOXnZbk/7v1D5xAZg8EWANAfvcdYH0UHXxdLaIUurXFpEz7vO5t
KImGXhZpM+J2ljFGgiReGGKBOs7BHAHnlzFNnoziWRuWk1UL9YfC87GsC5YtG1KklbAMpa/cWzNF
YSfS4JYdKDeFGJe3+yODFXHQwolSIuPWpJpNNKPjgW7RslJZojh0Xlus6xQymYPZMMo6+FNZylyP
NLC0K9Aaj7ohXNpMzguHKX40Njytkuthq+207Z8382zS5yiufH98l54HMVxg22kJsdsIj0Mm2Owz
d7q8EVsXb5wPgub5nr06v5y//VLa0A7KvuaHwL9dNY4RSafuhaTVUF5GqwnVk8yEZt8R1xLRtGOn
3PKr3i72N/pn4x57WJhmYBUsl9nbZNZhPrHZKCdLhWFMEXZDSPfRVM3zwkwh+SCBljy6TcIlsKJR
wrMyKoNfZJFl602a0Yl9bXpNpJnyM3l3Moj8nWSFUtvYw3uy468S7hlLrYEuC9pQiM3QFGRRh++B
hNkPrmmL6EAzcTkSirMY5mVYn1bbZoQiTbPqtNOqx67PgGs8afqiMGdaSNKWotAEc44niThiN+ak
03i3ALYGpKHTtnPJEB/WY1IudfykYjEy1eJBGdLj4ZPM/vuziVTnuDiNO6Tdb7kRChw+/hprn+XO
PSobABSV0do5WWBVXaMG/86lBJb72YZe3vrugv7EnNTKXFPu030oFwQTxKO7G+hu16xUvMBVYWbc
F/SPBSzAgfUJGCNlPoE/Q/bMAJ8XP7iJyj2JZiI6M8cbJkWJxga1T1S3S32c0AOVcAt38M8VFBkP
jYm6BmtWCvu7+vc2GdZRP1vcmjrREeRz58NnDcFZwSzkhFw8HMMXvy3n5r+/uUvnQh97rtfZLP8v
Wo1e2H0FW4BTuiJhljWB0xylTypFl3tAj9IGkmS7wKIveDC9pzP4MYI52Cf3jeOzaYfjmLt2OvDM
I0fMT0RckVTPkwLC1A9mEvD9FiDVv/MHcstqc8XxD5o9a//HbNu+7eKOzQYTtp8NyFdyZT0143Gz
d+78ETJcUtPyhT9gHo/t6niU+mAFGcLoVN9RGXEeu2S4/LosLVRfgEM+fIG8poSSygzwQWN+0g5u
l4jDlolMqNrAxU0d73l/XYSpnQef1o5MZbgdcPSmKEcVRxKhmrPT9PtwMTZUVhL+NEjJiBd/Y3Rk
H9Idt9zN/PE96p5tX1z8s+b1ZfEEqTqVSxdbCmSF0ch70GVwYnKDZ7tSlUfDhwVVL1yO5bNQv5kD
E7odUlqooJdoS55U9HU9fQj/mZJYhtom3tk1oqKFD0vaXci9/TOK+9DC/JQewuVrlY42NeaqF3D3
gtV0CpDkGV8CYm9QFujvYofN5mogvgm61Mjvwj0FDWJbdbxlK2dXYUrUoG5Ya73wKpFVBx071wiM
X3lWc86zFFonpK5zQBkXMx2IHDI8yTEPnyQ/dYJv9OPB84+c7k2Zs5VgX5jLlWRKCQxiSatMkuZh
w5Eh/6MSVM2ZLKRdpI0LNMk+0o6SKzyRZn4fq1SQJrDshjW3GxoUv2I1k/2+/LOb/ON/iJRCUNf7
rvkYzJbADrXZ5NRPpDRUxsq2HsKoSYgRugGf+cb7R3Ysjz3JUHOb/QPNddNlniGTm5/ZbxvA2gUu
05yhEZqJCsyffF+OWJs3LCpmQ+m2o0Bf0reBeFwnKihhUOsdGme6PfzMStpNeRiUscA5qt3sLOlL
qwrbDc+zQeBN3r2w4Iupi4peRXqGIw1+0ga/rNj6TRU5u6vH3AHcIm3qs0r8jtI6RZmRSQDtWXpg
4LCNvwMvtzPSJLZH3D9F3wxuJUzQva1j9n/rAqmdHChwTvoNgFCLTW3jIx8upr9hmYosomGrminV
ja5bAj6nHcd62E+DjAOa4QqXyYuyhwNpMHFoIGpFxskofpEOErEBSUl/URHsyAjq5d5wUF6O/nlP
s+qfiXEN/H2H7pkqN08Pq9rQTODlSBizCNVAhs3C282JMIHiS7a3qNCshGGY6h+FHqA3Xq1PL7AM
rHUYahpjsMGFx+A2hywsJxXhDUhdRwaxy8WIF3G/NiOXY88rxXH4KEry7oFANdc572rwUE5l1y3g
PRGBZEs0rZeXA5vXperN2wc8+e3hlzfd0wkCVc4De8f6MXuGroQNfgft5rUdIRSNqko/sm7znPW8
rF14X3wBLF3Jl1AtZpY5eR59e8R7m9gBpHDpmCNSwLBi0aWbJM15iwLELl7/WRPwUMcopBT5rWjv
PnvqGQ6coTj+jGQwAAJcLR5hLk24rx0PZ8j7XRXclvdM6/5CzI972whcFnfTjed7F8O9+7UNPR1P
MF28KEV583WokeHk9vTzjg35xGGIJrnHMxQz/bUST9pvCavPxPMe82BM6Iypvo4JexR3o3KTtt1E
ed6H744bqnwPnNjAbbJtsBK8EhAkn1M3642pwSbnwZleC+yM6UJEBkIzA7/IfUuZXsBpIYHXiTFZ
txEKo8/ziM1JGDz7jOoFHHNZrXxqBB9RoXJlF7GPgojBPUl2RupwERMtw7/0ES9I3wRTUO/Uxdzb
S5BPHcN8osm5jNFi/VA2ybqrq6yGNSpEgMK/Fvhyo1VtfP4MovqddTmgBSMr5lpE8i2wIjwiTNqx
fHQfExs9JUTJLWslXf7owKJOc+XAl5bgu/Hqn5d8z3js+aKkT8XY0DNh1ZDVJnGonSPqtqqAXImv
aCsnlH764KTdp7zfLkr0avgSknX8kc+UfP443okBFaLoWyfWDKpbbLuC6X0x2uYuJEtWtruFEpo5
Cy9NhuqQ2QtpgR7/2Ihkx5R+WPmvxQWfkeYhA2wCAEmxSOC52vDacGw/OAVUeLAk+D2tuGL0+6MJ
BVUjmKUnIS6HxhjU3nnMnRT2OuAQgJnOzqzenlJ+a70UNFbE3bMEmm5fDECpVQXvoLf0T3MJRTJZ
hq0E1JFIS70fOTYQ9L8MbUoLCw/gv9T2WBE79N2qammuqMiFEaxuIc+tgh8XmlbSmt8m+6S+THxc
XDnSoMCB5z2+HBnR/7U83T02iis5uyCZ65vDIuJy73D0ON2441gDGk7HtuWogIaTXiGg8jImYa15
wC13+Dz90RN+QLehH9mtQ6clEuAMCVWfE0rzPeEJNmtW6APkDf8qlPI6Y8Cb5InJVl1wf/9XwzHK
u7Scqgfp6V5ES0bENhOE0HX8Vh6vastXKCoBxLPZ52iHHjZrd8u6XK1yUeOiQ/sLIIkYtGFy1pli
2lZ3A2fK43IA6UWcHKGA1oc5FKxBxnMQrp84A188l5A0mWerop5MyU3RDVj0A/+9wK7ymgaHo/Kd
vIFTuTFXRXSRWzIGlzuz/sGHOUO49E9pP8aqR0NxSTLaTJdi5AYQYyoxxDhFV0GGpf3HnxNRdWiw
kX49dyh3w01iTRCRVAFz+2AS4yTfbTiQ9wjKTFLGLLPlPOzwNyGPe81c25sU0SGqL6jUmHQ/Q8G0
1KNQLwvwth1RFVsTfxK1e9EOLxWInrOkp4kPsFakGeGRKGBo+m1y8PDB9lRaNnsPvDgXC+g6iKfZ
u9Sg3aoKsMjLlGaNDeoKpuNDTwRHRyHHRwmbxUUQw58gARwXQJ8/WFmX3QGSws6ewp90Esyy+PTM
p+ToKRwRqg00DJKbwYLj6cGp2rvBVpQnSyaIc7J4n4hFsmssElJpAqJ50dyoLcfddAi1lKbAHSoS
iyX7UhwA5H0SqlhumcoeMHtnyRbMOyjUJkX7ODgjQ9L3KIa97GmGAJwZSs0mgs7nUk36HL53/7Xq
oppROqFSGu9TX6KsE6AT9bIRVK77lyudpA7Fpivwv8WCMBS6QUURHn805DYN872dNastadJ6VPrS
E1Kl79Sd/277QltKM9U+BoVAH2fJJSFbwLy8rtZkJoY6HRPXUwbMX2yzq+i9rTTlac6blz+LpI8H
kzcFlu/FPZyXzC1aeXUulV+w6Ry8dFqgNtkqXA77aidxt4h9GCdoJudV3Q2SNbPn9FsbBdmu9IaL
VJ2HLTBf9h1P+bSXa3NMOHx/iNVuudcw2Z1D/BA1e11JJtFSQZHyWhneB8yin2fxKHlWIJWkP07e
e+B9BBPlr8hluW1cDkSWRxg8hPmhhRvabpZOBD9C+X7bW//c1Av3iaSfvNkHDqH0ftInQ+K0Xllx
BT/aw1Wko9HXqQY7BSsncSH2P+4/yWzXypt60K48Gz8BuK5N5OHosatS/NbOfLv5To/c4JsO7u5B
CvoUYlbbpMG3kBR2kyUH3/pDTK1jz3GSP4Ju9ljwHYgo5wTlwfk0EEQYz7Xp6AeXF4pnWu04YK+U
MvPzY1ugynAStWiheZSSP/HzXQyub1m1GodUh0FXdg9gYeuyrRK2MWU7fA6XVgSr31MwnoZu9i51
YIZjC4L6wwMw9cRPVG//y5v7DlKZqTQk/2nVyFu58b1GGtPV6M9tQnunLX7FT2pEMN6dtTKlbPPj
YQcyxeWVEPg9tjQFvSXWFBoL7e+y3zzsSSpl/DpKz+KnN12RsxiPSllVpDt4RTM2Ihk4eSx2SinV
VNowOjFj9xqulO/+WFCg3vFZcOFC+K06IeacLl8qxdXdKLp4zls9lbd+ladGKtDDirUX7Krn+mgs
sEMcysYCD+rWTRrgYV8eiecokDBe7RKUnxvGJRex0xwZgBRI4rWX9vFriSxg9LzZMZVMVP8AkioQ
Sm1q9vsJxpZ2m1QbdwBQ2IVvFnD2wVsxh7pldU8DmfFcRUw0IytBzOy4ndXlYOX+j3UuAFmvEelg
fpyxwwHPtW95U1zkzl831H4WjBOJTX4aQUweSa+X1Nt3tuN3gEGEdjfs07FrxA4V/AxJLBTqLzNO
6bW40OBEXR+hqwZGYt9RB0pQ3U7zJEiicKQ0vk8faPco4lGhIXMe4SJjddFN9B3iltFB85WIhxRZ
LOcA0U/8w/5juugvsNksX6a/4WO9RvNoMF3A/icpDJVZtongaHwdujLWv6DpST2sfVhX1dXipQtR
FUB6h15Iut3HeoCOqy7ZGhzYgjk8ORxOZ+TNVBv+ruO2sPvEMelVqBXlkzSvp4Klf446yBJWGydL
MVE6QN55RPfJ+/cODLUELayH7twV15Otuo00+z+4xozwe3IskyZfx8nct61ihHAVmjah0hPRdfex
kKjB+PgsTEGr4tm/+s8Sijx4SzVZWO1CvcUnR3lmVMFCkwq77+FMFfPnshN1zWs00IaLPNPMNnQu
a7H3W+LST2U0BzYCqkydnml8RP2A7BNLAXFp62GHpOyFomNyGlw20mBhRFN5Quj8d90jBARyGEYA
8M+CnHD5iXk3iutpphpGcaR9oXemCMBUKfG6by+e+QXi8Ej4i7vXnSJ3iMljCEVnm+q1lxEzi1ui
lG16INeBrYUd/WFdHEDp/4aF6F+l+XRaJL+96+6gvHj7/fTnQLgzlGb6FZL2ZMD5/xVZ+ZTmBZd0
vlIhHn3J92R/gqAp8V7QXsLmEOeufQ012dhAa3zxek1Bf08WSV9aoa4oDYfT3stqvEhgzzUUVIhE
0loeASEXqSCnfGtLK7gXVPSNU3oLRznYZ792hCDyHqWS+mlbtTWQFVQ7k2MXzZXXEEzV0CtRZfek
KvKpw/YrJHrC2LGSjOKDzxlL5X1E0iQR7JrhzCyXR5Oj/EIDHss4SD7nsUPlLBt1dvz3se/W+xdR
6RaTWT18vmRUtTdedk5J6WTOcNJfameafrGSiY7EV30xi0KHEPlQC4Y3jEFRn5wJWiuh/2ztvDi8
x8hGk5EjhU/hTLJ4pIpMyusSEsouFAADtR+1BZfCUNj7ISCyWsxQjvXABgpTcT9ZcBpTRlHtAyYQ
qeFcbclADUrswx6WwJ09xs0L/98m1MJSidHX5tQ/V7j1L/Y4x7hqlapoHLSwrg6U5HIfmlnNta6i
xmokS8cVo3AEpl7XgalQnrQx+1l3m69gGDQqkYC8g6T/O0ZWZYmcIb/4yJer4f5MoaQnJLTe5A9q
0LsicMIzmBb/sSQCiNnJ771NESe+OsH0uGB7mZWwbvtBnai7+8JGpTDbZsD3DYxr/leWbmgl8AIe
FJeYbX/HVS3+KxLun8lVWn6lEsqE5ng8ELmpqnLCV3oQVRdPXVqQJVC8Zxiy7e4vo601B13M+75D
n+Fsd557n2XWZaysteSj0TDb19AmfFpqugS/wtGbevjF8c9TdTdGmtcVEN3Capc/R/wGQd9jdF7j
xsc/dKFSBNziI3JSxMTvVimGOVTf2c5gVg+GOpeQz75KFTWCSaxCFFmTSZV153v0+/E9BOIAxtXQ
IMadoqPSAUoWoImY/8Xq8DpRiR2vkAKxQ/H/T9nDHELxTrBBs19ptR4F7f/MLXyXlI5acFtqtw+Z
tWqRSMK/wYSzY0T0xs5c7KN5kp8asY3l8Ce0zM9/NRIlaU0GCyOPS1/NAojY6ElwSr2zmA6Z8Tbq
+sQ2kXdawfHtnaWkWfU01+aSaaEW4ULMWD6nlwHnjSZLwrGUwOh57IJJt35b5OYe5fo6vNkabnS5
aFGBPidLg0mOiNYF5dRQyDyKq/zKSHvNr6+//3EQ0IrGBXmDa2OhtrtUWsrnemMb3TdP1bWQQkXs
CSrb0GoLf8237vjpzPaF7wzzHyA+v9RPHNgnq2ehqQPKSVV62PkG+vClM0NJQEIwF8diccF2VFAp
tyHu4/W3Rpnu295YrYZQkf5V63Ec9iChYEX9656VhNp9NoT6GW0WP1UeBeyNyaTGI23tZJ+lWQLT
Qes54sgCMQrg0wXz+tTsHWYgNBkKyJm7RdJM6+3h7lwqYxH7d9BL1/SyBUDKrC0zDrg3OUEHv2ls
6gFu641A65PEs7K7gRUCZB5oqNZ1HOCrXQEfUhEwN8AayAxvfJnVoF5E0rpTRvy9Vb+rlr6Pp7KW
qzZfSLYXvlYzOhjPC9AFUAmvrqj14Fue1gplQzlrCqRFyrDcuUCV7I4H9d6pXClOx0W+L88Rokwh
++TKjX3L+pxqh1Btq18fTrCFNxp5MnMQ6IfAWlcNZV1AUVf/5Ma+vW/OESJ0bcz1i94Z5PfzBQWi
cau4uK3alds7fxCvyu225KYKznPdRLPfZASfPDL0e42NnDFH81p/gZ20Oj6gra3ngGcy+VFZG14R
wuuEoDg1D8j4ESoLbGDDTH1Fi0likoLG4NRTQSAt+B4Z/3BQrLyqLazks9igpNP4PgUoAdC+RmXu
oNOxc8nwm5z0fONHIW0HQSKap2T7hRKDyghrfxLdg3wsvPeRZGuAOfwFa9IUTzXmlAVGa8NfasDI
utQUtoSU8hPYSeZ4YVB5xTSGZMW8bMx2EFloccOBmkawbZTFiJRprCGZr9p9eFhwW92Ils0AJcKt
Yz1mGxkdNq/hadXPdNgd8s2IbZRkNAHJW68CKPycWr5Ypnf4AyH3LbH9S/JlGjeOKnHS6Msy0QTi
asMyp2iOGHGL8z/xFpQXQ7KMcsfOQ142GY0s1tyvt2y0VJaSYFOo/brfTvs5qnUJQRLtT6fMWiQl
ivdOxi3c96UKFGbrIDguXr84/BXnN21F/xls+SQpNQB9zadaUmDbkRh/A89NMpcUPcqeP0nzUIQj
Y93+zBO+f74q2OPy5reC2fu/j46ImOimWjS4PlYITgqznhXVJXiuECcLPA1lSMoXp4m53XjtiuwG
mLYFF492Hm0eYA9apEYQ8rYCi2xUVaPGZ8ZHfpLWzOXaypGTXECGo6uzFOVixucPFlJx6DcXk6L2
AYmlmD2JndTC5QIrBF22mALZiT6YYa9BS0V5uX8zzOoYoqrflYuxTwHoKaMCVMsCDth3/rs+7h+w
lOp6ssA1dGgJkAn7VqeVkzg+1zGLvvo1NaDDGYXAbTW5JZ05cUqPwvdlfURDeuyyaVOdSu/4XfGd
jNQ7w6eE0oHGrmAjsp26wHYc0v/naAzpTL5KNI/zVhLnVL19OZ4VT78H35FdkUfd1IvqrwROdFtx
Y7o7E3ZUpskfUOtxiyqSK0AuTFNKe2tErv0wmTFKQI0JbPfVq+zjcOBl1IUHILofAELBYR780vMO
0+3RsLxOkXJzkrF4da4db+2ED7kyDDNqfjS6yF520erf/ayiIC2WjWsZQBvLgxrxkhjtRH1YyR5V
a0DwQyVoZIjTMklZW2THZ8i0LRl6fG4prnJ7hiLc/yp8NNGnzY4G8U8/BI9qq0QDbgkNIhPkHDrw
wXCfvZeIxjtkARAvjjH4DCz89646li5vdB3E/PW7H34U7nhigPhpbkJYQ2cIXgj3sW0GRDma2NR1
ZuOilZtzhYbaMGM9VXAarD106j12qzyJu7+VANaw2zw2Uj2PFK+u4gAdiNeTTLubuzo81Zt0yV4W
0u+KmlEYg7372aIHgZrkFlrPhSCALe6IyfOm1u0SPoTUcusl8wvjli4BWcm0NkeiaPlVoQrB03zR
UA3z8+buCEivsdqYGkW/QqZBFUK70oXM+npZqEAxXPBbI6P0fveCEezN72PgbBOtl9moO7FD37n8
ENB7H/FKG5MYJz6oX2j/uBCvdterQYQNwmyYaXtmQmSmFE5CUnsZfy9FXYkxtoATVTjR7J44eFRW
jnJAEKAJwyp861Ybj6iOFpSULDUjSIhv4SMfUGMqXevShOOOJxdDLFEw9nAGz9B+2KnbPA6vx2pe
hGvyNupr6DyBrQETuj8nYknyr08b8IPc85XAw9KEmzYHjI5VhtBHckV0LNeAI/WQgJofdixHC+LW
hu0E6a6/s2v7fvejBZuOlFh7hEIN1zG0QFZ6++W01SbO8hhRHy1Z7TepliVogSDeKaa9mFbPCT9k
hqxdcHpRdSaHsERtrTs4e5RNNSUQvSQ0vMlFMvSW8cTGiplzOtsbv7v0Z+eEPCfUvNerakq3c3Cl
xXWuhIzQs6dRfeZAW0DjB1TnAe3aJvHbLCuOaZEnyViaOpzhr4BUxYoviX8Y5/GPjIMvqhtEmKkg
29QnPPEpVkSpt01oG+beuivP5K1oNVqrHT5CKgBnit8bA6QJ7M1gQ77fNxgfnwLSCHyC0p4xf98n
nhpzIGo7fdm71NHBe0hb2v1+Ez2pIdaI4tiL++j095xdxhhGdU7e/aHhGgdy8fpL8+0jLJMYjz5v
EvI4u4Po/vwlmhX+s19TbtHD+PxLd6LFBu7M2M5t1VAa0bKyZhwGd+K2qbriKpozg89nTkEsY6x8
C+/VtH6r6UWc2a0bMHDa3P677Rh0mSnTBjDrQA88H/5fWbER/Y/KkRH5djHD2a4+jc/G6kExDovp
t2xXtBWwO1E55xGNlwg4IBxyf6461T6+8bGgfRvgvUNC6NqOfgHC7ufhPr1/6J+N1u4N6/RXkkcM
JGBDjFy2XWLVIohCMaVGxTcxETOEzJz2s1roMzUno9wbCxP2TyXtaWOCqlAddVK51sLFkwwPlTGK
Cc31628gKDIU0EEzmIO4LfDTX6VvX/dEiqLxugCp6f6rGmCa0pIh4wy5z1hWF9LeDn2KQ3qDJVNc
EYvItCG5Nt66y+zPcAAKMZfIYfOfHCbF0qwkGXcq5B4z1ZTaY0wPC9kNjhjhYtAcUQN2dxeNhTl/
/3tuR3SVVinycYFB0X78xn7SxX7sod8pDPl0dA8hqif8LoWilhxo657BTnSaF8KgBpvN0+2GXxmw
P5Czstu/SOkVAUHftp1iY+l4y2WCqRYkKEPYZI3orIdxjrT9VF1g5mFXeq333+9MnS56x5KnP69T
KQiqN9NdRUtuYQtCfD4xrAzoNmvD3IZYVyaVoBG18C8/Fhhbr4mnyrbA+0zvAWetBAlCRNgmnCwF
r1kHKML4sA50X72vzATMvNXrYyE5H/niFD7GpsURRNRFWHUA9I7p+9yM4kVGwWWrLW1+nOWM/6Sq
oyn8aSooQHiTgVzPszqHJN7bqerfz+9p2jbZrNkmiqMaXZwEgnRjLkuDdcRm1k8l8+wyuGZZ7yDt
oghDqedh++0O4oWIoaEE5clKCW0ERMZvMBlHy6MENmunYnv4soHGONlW6KexZ4DjiOm7h/wzrXBA
gTshg5b73apX4v8X4tgPedLMf4/80O3mKyp97rJFSu4xTeU0pkZLxYgP+pNEfNw4UhTJ6+Lcgk13
QgRWHOCkDIqNjG0gJ1QpoDMrOpSABfepEJIHTJFLl2nESYGizEK3YXsWXW14reqItASgrTQp8UFS
hgJQT07T1axSSmgWaafVfiksz3BtF1KGMixGiIX34NpWtEJApJqdrMrq04NV39tfJ0CoAYXAZ751
S24qf++jUukPRro5zwZdOqOd4qAiOe+HL7NyPym8bfvtqwTctQjgQgRK8hKHlASYjkGBuabIx+xh
xUlg3OnTMNjTar4vxGETKVduTJQB3mzRGy90zYgUqFfQAQ512UP5bulkDRUMVtCqW1G7SjXmvTMw
rsc58ya58PcSSJexAu4Nya7zoZ7zcJ4D8Nv9MQDoBgr99rvTrmAAZsrkqNv+BDWJYIjmaIAefxsL
0vJ2fLj4eo5tRA01DncoZfSlNt39uNMf+fCxApYXK6Q5flKn5tLjtksoJNeNadNOITcsoA2o+xqD
dSo+w9Kb6ynYuXz2117tA39QeQHoUwnyDPCNaUM7ILRedXqXsi2uaLp84yVw54dTewR4aBlrZxzw
8QNwmCBdLPMd4/MHV6kHKHVgHtfcDstem/bhlxH8MDW3+5jKC2UaP99PYR4+gPYUMAufQo/oUhkp
17ucRKHTZsdjYgKrrDkJ2yNV+gPulLXLrs9WDWgHRLDkB0pjV90Yh/qWfYebvXMzY/9hITty6/3Y
8cKxJkHp8xb49YERU698/wIzu3X53BmfBm6kqZZT0rjWyPlkd9zSbPj00b9IDnXpEQ4qsbMxM4AW
DYUuKW6zPLsQkpLVli0HAm+zjvCEzKwWq+O6x3Av6rXuukIgQBMsjYsrqASgNJbVjREe/HJo0a8N
a4GxBhiExCXxwGWKbO38wBWh4CIYF8I2zfEvO3WX9XxgQz3cvHjiw4RAWS1sXfDm+iCbL5gndyNv
423Uls8FaYzlGK7SOtCiyCSkiOcoJcZTtrgXdfv3Y7N6njDK1wmpubB3WMvwJDLZ6GDcR2oa1G6y
yN2UYQqGxcK+LW9f73whAfw3hpXf0XnntFTyl8AUd7fngMZZlzC+8su2ggBHhhGz8vZ/wC7SfcOt
T9JrNauJ0UuLpdgik/M3pZKaAnH6Mt0W12YbvbUQxYx5oOtwdC7slNwH286qmRv5znfCRf2ZME1b
mtnkge82zP2x+Pc4Nsu6b+Ii9PmYxC+//KwIjbbdMgTec7WyUIaVSLS811QP/YoVgv+WE7DjImkI
8/BWWDyKQK+OEVfKQa/up147PGtZ9OKqo95R98q7sH6A5KxcNXjbmx2vtB02+jrDW1c6aPoWjLGB
ZEsnvL44B+RFBGsxjXhjTJ+CMZ9Pcw2ZCWaP9rU/fV91lmguEou9/btXEUghcJzQYZ4C7AvmU/0N
tkMANCu52eB4hxQiQJKpQ7MDiJTZPKkxitF8DADx5xnnl4Zd3jt/XWQmkxJgtiBrNswyhKRDjYmG
gF9GxMlJODwSxWyQJgz+MJ/WTq1aYi61X4Wa9n4jS8YGre+Z2hA2USE5wZFmyx6zy50hjcWe5n4o
efSjGTFs4DtnAtHxLKsWC1u/0y1qmg4YuNgWTboEoC9AlY1AoRFfRm8keCMhC4b+GrwqQM+qRPK4
S3t4huusIyC9k+3CDTAvgEEd+ut9zg0PK/Vmbxv5VrVXbvwZjq+/Kue0Xjr0QqfHeaox3oBQ2xOC
iMM+iQV+VCENiK6DgniBQRse0TOthjeTbU4wpc4Aox8MD3L/Ib/5nu7LrJY4IoplrYPJzt2LNz6a
DIfAIC9kSVqYJAMbzwKBKQ9FSShpwo0Cc0aM7RJaRVK8jqIf1Qd/or7nA37mLfXS81hZ1BUUsl8M
DCiObQJrM86vhoer1N8v9u8Mna1PrDqzTUi55RiB9sss6ka4I2yTlqUb6+9rTjNxARQQBUD2nQv4
A5PihkYgr4YY0Lk/JFSoDVp4mG+VcaxBrnhnNwDRo4WXRTFTcg1IFbyfHDyRZSJa91Flr/2M0hWo
NKxGeiTRUbMCDzbp0UIXwuMMcvJZ89iYk0SxB2BblbfOQ82ZH2eUkuQPSrpKaim7la4QZALHuURZ
eNKADNTTEIwR0twMp9zwCa8YcKI/FqgwCG8bodkOwSBh+Kt8q8L9uac8wtAwkFN0MuoVI8VWDUy8
mjMxsNYZC6oPo3Yj0Lzj0TuRpeLFDNGLk0VLKwQ6KPqmRg34JSTrxXH7OeBFNxj56/OwIMF8mll/
zjGt5H4m0UXiEkgfnaPu9mv/Ockx9mWVt5vLdYN2YE6ZuRx5zrxdYaIDg1u/TaNKsYXhRBhFQ/jA
iGkIp3tSDJoln9cDllR4P8iV4eReNPV9vI7LWLzzZ13yuJVWBM3J2GUWQigzgjacRP+qSopbLsSX
P+hRoZ9JJ1IRyemm8evdUSzTVuHYda2iLqvwC0QQ+NkifuvhgBxr+alkI8VHZTGfIytv7nDPpxiv
rEzDMivbSD84PLgR5BRsIGASAri/a2hoFnLTr9Y8r44chT48fITXCW7ssCeGWqijitNBYOxHJL07
+maDCFpTHVYZ+c2Lf8uFljHvWbWU+NMH8AkvS45k5Rs6vE3/C0V4BlWyatkfL8+RdCtNuzOkHNKX
6z780E5ORr8Dzugnl7+mCkD3cYKu0NMxVSIPUc4flRrkWL0Uuv+RKHaHTgQe/rTrWzC7+slszgzC
vbjPP7J0I9Q+44XiB226HfRQImPaLudlmGA631Jf7jFHHQht0RhLE8qPS+oX2M6KULF27F9ASuuO
le/Kat5S6ppOEnSfi69c1GLcCJr2Xcj7mMbuTxJjyzfStS3wzuWFDxiHDfb5v86PIfzYsXPqMRqq
vsGxaMkfRdqtakHGK2uWD6ULhp0Jp5fOo5AesdgFZniAww6DNADkGRTRRx2dNu4ltRhQzgt24MDc
rla7LpjnRHHVO7e5D/1/5KF5JltN4kiM978cUpOTWb2CW502nzI2tGYYlBnNguJ092SHZ3drIx21
itpbSDhABE6zw66G32UJu2gHjbtxrx+zRnI8p24O1qeePMS6iGBn5ksOSg/QlUeKTf0FyfbNQ+PU
SJ7K2O8WCjLEClARcoAXeAKZqwdMJG7kQjvmIBqthrHuECpo20+JtCRo0F5z5i91SE4yPqW3bevx
WYa6/xbGChl4nB2BTS1D7H0h78XPuWKlAX/1Gy3eGLieanqXL/4JIEHSyXwBa1Ay9iQskE4Ae37U
G2YELkhQ4d8+SWV6qM2uThwUdQu/N/q/LQMrUp4E0rdTNzUJGa1yGO9LJiIF8jHrCnJXsoFbRIaF
ppnzSxC6s6KAVuWJtSBcA2MFfTDJ6PHKWOIe4WfJPRcRYUeHMJpHVBhOVIQnUEuWtGtJuU7tUWR4
K67D5dKBq2xjOgr+ugfhEDnygxQC5kgRSguniPy5ckGxqqUphibskF7BOL3jt2gJJwQ0UZtT1PAM
rIHm6ayP913U1sRB2laD0b486rNYQbCLKZkUV3iA1nC0jz0K8ibUhNJfqjyqktaaePEFFpzk5UyB
ZM0x24YaSBrWn9pkaNhmlyriuceZWJPJxFd2wuNysttCo3We5cKD1PRDDdVRvFcHtO2DZAVY+q8m
64Ox0wdCT3vLBttjSFgMuYMkkIcU/j7X1w/fk2Bc0gqlNtVQRfamYrULXtP01JIPqCGdbKzpC9F2
kk5YnSc55SXTej+FRXQulB9n8GwiiGX/EA30S/+syiai3I/WCzGS28WVyutSwvYpNGJ85cI22OcN
ApbQ9VqmHVct/XDDmsLTz+3jMUeEqlMu2VQHVs/ErHWeQWGhczyLNqxRU31P7GvK2xJjeETV7C9h
1zdhoE/OkfIBvrZpXgq3n4waIQLVakR5fZUSFizzRJyy3z4IRr3GxZp8+C4fMv0mdEas6OYJPPK9
azKeFYe6hFy+b6OBVW/iaWrKYn+Dsqc2hPVTllLN1oI8niED5h0KXxo87gl4036k1MLfKYHfJQO5
cnVpd+IpXZ5yJvTnAVVTwfH8YI7/5Zmwz8PinMyVwcoFBwwfLhzi/i7OCPnNpVQkAUZDcElJwXEm
rxpcUcJK/I3ybdfeb7E3Cuu2QJ4i9ena6jXQdJkYXNDY4cIE2p2J96kF0j1shrijQoHdDWEeS6RR
HSH9uNScBxHPULZ9K1D84ZIyYpcTvVpGs7hPWPArP7ylfGbG+BHJ6n1ba/p71agG6B49VWKRAGFg
eAUX6dUcSlrFszONlrBEeto4aNC5uDm5kruZeSuD7mxIxV9DGtdeVNQyPGSnK+Pz7QYV7Be6oWvI
dkGnbFUHWs1iDPAeHkUod/NjAPhSFTxXGoOHykM6ga36N5++bYMlf3rek/JC7C8IxSxDwHitCSuh
xXaHWnUq9WR4CT8KOmCdcgqKthHGDzqsN3ka31jBdA6TaVa6oaDJpBvfuz8QoMlpQmXfllSdzQj0
E9YCslmtMJ61cjYTqvk4YOv5JfCV9gdGwDcx7pNxHCGZI6LWdeOTtOeOae3PVwsKcO1VpsKWR4JB
h/hrM5D18py5o94ONEzXVJW6nSIiNquwS9a4+xzDiP66kHHrr/GzA7uAzcjMViRv7DeIy6haEQh6
mTASUf2nWoUHo4ZXIIYDkQbtDa11b4USzTDutVl62w+kPO1PrHHZbN7lWEWX36vz6BR0qIgcJS+A
XgUrNPzJGZB6jRYcjGPDmsRqHTFoXH/7ug4cS8veQCWlvPCOm87AanXLgubzY5VyID06GBcr3x6k
LHQSqZdpZ4ArtD/Z0O79XuwTb8O5v4bBQVgQzgbyY/KasB1Z9/uGaVrHR8+I/xAZumiWcsKNbLZy
hnnVmRRF4dCU6vaCGPyPZAcOmR7+dxGq4GGJcdyRsKKM3uOqQrQECWn+FDow3w6fR8D9+paxcMJU
T8ykGA+yH4QXelYp5UPRXmm3PohJnTXiQkorl7n4k/qnXcw1ge3TKBRRpFk3qea+HXzxGpmqvghq
h9azQZsb56bCAbG/lb6BByDUMVrB2im8EnDdbGDadSFfI5L8Y1GzeW6CwZTksX6qTovOn92RBXjw
mTkOZ8gOgXGBvzGMDmYEPtFskn85Nhe6syLyqPkeIax3ZtBYUehfxKRVbvY0BnmSLnUAZ9fUrj4b
Krt7DyiMmKAtCqCEnrBKQGLdW8rTyt90tCI3hgmS3hLXvYGy57x7QcIVpAXxSXfTl8fYlMqUlOBQ
5TinHcbrhcimCvO04y3Im4DwChUv7b0y5fFoZJPu3wZQ0bEf/jXvBB5j8RQr7unlmpgygWaZe5fP
x+uDO8J/H93Ti7BTgWCAGe+X/KlGYoWllFW3U7gIlLZgjIzhcKUvCpZpdawTHShBkA1sFW005mah
83viQ3rCEZ4uG5qVp1slnhVadE+vNbJ12KhbAYOiXw+dxDqJxeEUNJZdeKWMmSNoC4z6p8IWhvCL
/ey19/uTzNHtgeR03832YymBXOouDSiH96VjWie6wxVST41prSbQ2ta0bNrvHA2anUGOPYm1czOd
1MFE9c7YUbNpZoJz+TIOL+IiG4Ay/KsLtBANfxI8C58Bzxeynkv6xj5yJoUSfn6hwNENPN4mmsub
g/kSLFBkBTVIOm8G8OYdNJw/eBIBjp0PVl6sGHLP5WHAdX8hjyG9bzsOS2ngUC+8WJuTbmu2ICUs
tQe19SRnUjeQ7IKrZvxOwP2N/dI1BwwdM8g/KLZZFFBbwFEHzQw204WOZNNY1d3oy1Hc41GzH05o
f7OdxN46FUPYr06rVD6eyH0nHdsVykGDGfpiYhzNXwkrRN8hTYo1awW5r48L6+qQ2Rn02+ZesOWt
g6H4lGy04fxkKCJZQniB2g7mnON4F/vGIVCEBcRrTSC4XBVwzQM9LHDWzCWy/sYoHTLmIYI3+/S/
/vt/OZj4QzKola0w7m3czcMSCBBosgv/6AwLBS7eQmkCRhW5rnj20aKPxuAshTS/JtxHLZS5Vv7Q
6dY6sxCmLG5IiP9J4+adaAVazguhoIeEHIapn5AyIc7zFljxS+T3dvzyrgy9Y2oxyM/1s4id/PMR
4NoJhFb+2IKUrGVik/dhmVnbMLlw8ojMgtBMEpDmak8iz761/h/IurdcwN6WjgRMXEMsYUpuCTqF
5TTdUc7n8/W59KNOmbti/RVxeODMnvHL4FLoPnLDOQif9rBWZ4KeEU1wKortbbX2ta5vc7CjQFAo
9OAH+x4a5OvKlNRcIZz2SwZszioqN7KxC3VDlgqDm8OJlzkYFi/41ltc4ISVX0USDqNfu9N3kXw2
q/KoRSY0GaPeA9hzEYozunNzE19fkD03/CjU2EdNAqGpfwHC4Ihsg+NSPZEHib2xGOowpdP9hb2q
ZlKpRvbuTazfzt6Gi9y4rEGob3pt1ZW9T0/d0BpaBOj2Uf6IPg2lTfy+kioAzAN9qmAfqR3udm+h
cb10e/ViXGa675EgSuhiGduiT+2713JCnVbZXg8uEtGCBflOUjci701yziI80KXUTBI09L389IHb
w/tKE+Vkvr6zdK4nh4A70DWdUHzmbSwass3S/pa2sWtcIeR6vMBqnfL5WGNqecn6hBwn5wkMQ6tL
MOWKjgHkSxUPtFnxEQcOcFZwkmWB5JxjHk7wd4jfP9oZkBHkqycCABFpdVru2XPzAI8ygZOv+zcb
DJfxFeBfK9jjBujHjemXdjq61514571A9UTUiaCWPH9w0Y8W0O4fwaxCJCJqVIDxonOPd/72f2G2
OYGOhLKhyd7oXymceoAhX63/GbG6FDSiqAjZaEFYBlPDo9mkxSchx9TrdiTUtegqKEBe7sMQIbff
6ulqXjxRQpvDIgnQITC5OWyoPK293dwkHNz5u1u2Pz+hEqewhDdSa0zhSXS/G3pjDGatbpMGIxut
ThMtNlT919vbjnzyXXpCheTy5JzZox25z0dzeUb7rqfBYd89HuGppNss4iVoETKJBp7owrbyXtxo
c8qCIyFHnnh40H5VXvkbBftbK3ykmdZTfmEQMa8YxrTXoQ9DpUL0pLkNlkv4tdnQ4dInpbDu8Dfv
FewHpYsv4YfIWkdU/bkcLr1i6KA55cSUT7sWIIknf4sfVmFdW2ZoGzoGvAWxUtY2YacaWLXkjMqz
Va4Y/DoZ/eE65VQzh6RhIsBcILGButdWNQSYbyBlgpko/X82ONIM7qtdNIEZ5gqjt3+yZafAo9n+
Fa4+Z0P8f44GlG1RuwomfLW8ZkUJbwsPDu1ShuY1JqyRd73gwBqlr2EixIk3sOVdxROmMzwrXoxd
EEkxqzeq4rM69P1IknKHJhHQ6n4Kz6kw77e++n9rGg54Rcglv2TJn3DxrWSbIpmj7/KMU5VQwfiW
USbFi+jvu0gkur0hqoimp6wiCvcv4qNsgC/ZyQ7DC+ATl1UyKM0oAoEcFhbOrlQdwNLJFsZjb0q4
HLaKAR6cJHjq1gs4B6MKE2PKRQGGsHpCjAJtf5YaqYY2sdKm8ew/8xMmzZObSrLpsdzZjytGxTxt
cpQvAIBbI/M2XSL67pgC/xGx7M3gQieP8bGbqmIg+A+8a3YwxHzuXHTpp1TL5V/smAVdymUibYqu
5rxr6PDputmHnKUec/P3tWm7Vct5ylXMsVBs41xheups6QzmdvHWi1lvWqe9QdKF2vd0Ii8ufidT
w4AjhLd1LnJyS3+CFtyI1CyVbI1QsRT8WuRle+ezrtQQlDUMfdTYG5qxiVpmaA+LvwSP1TvvMAUu
VeF68DvAx33sD/E3JUp94QmIKmPSfOdHjgIm5oIJBQ7kGoLJD10436DPdjJ+BBhB3X1UkinDP9On
000TSOLvePU17BajheuCU1bybEnLp40EgnOthA4u7X8Vz3mVvKVpWmF0FznC85wyDTUe2oAJATaz
j7tvM3/EW8/dOsEbaaSIR6i5GG+njbcRdxetWXztBOoHqdQk6cqbvKOrN2D04X80b96uKAaK+a+e
UyWoi28WPTXieUwsUm4gmt2zCcKTy4MmKDCG6T/d7CCng/pSvWKCSgUzdMtSLndQmd7YV2YEcdK+
ASSUUqgmAe0EQv8PwPZobxEo+oYgZNlKwLGTTc49ZPX7ELY2JZPisSc+qlithoDYLbJKRbx8RQzK
uw4p1KWdU3GB5zM1AgqALdTjoKiaOynjJL6+ah6X1sR/7A201MwVkdlQaIEFLawjBAZJSJ+n94QN
xN729La3riKG45rrrEiEVA4SGPx7mIxXWiiJEYxOpi+5vAtYtYWiv+fevzHBm4LtUrHRefrMC/Ip
LEo3Q99XnDGAwFT1zwUxX8UqMQffTciiL3vqV+gQTc0E0BSNcxcVZWqMszl6Vl9pIyv63GttSM45
BqeOlIXCmPceI4UzW1MVVW5Wk4haO0KBaDfuMsI5didvCs9Pq6miMAkhaNEoBTs+EgUfr/P6Z5f8
b8Ql7g3neygB8MBCjoa7YNWxePzvUdQq82VTn7H4dKpzzlW7T8Z+GvjA88nZjIRb6a5dLjNiN3hI
6UOsccMmta2cQWslQ/OWrMvdJwi0sP+YDxmYMcJ7afSTAdTEJc+iVtatU6lscChpsaaB31ZlN/2I
XyfdhTinXeCWjTFf3IrmaiawVgX/6lXW5qIqjWmL5VeOCP7Y0XDM/hda80U7HKQmkoWjEghRtDQL
RsjYvjr7dkZwzb4XoRH5XvW5PY+vW91MMIDTdbJI+1D7PF9EoTHD2H3wtNJH6ZiMFXr6KTfsaoOP
ZuZ3AQF0AFAKY1CA32dLVdy2SnUn+uZl7VXJFliudyW5Y/ZoPaS+BYLZZx2Sa9ub/DeA3i4jQIOX
J0PnyDkV31MQRAfd1fBSK07l/FQy1vgSazs/vnlbqxQPZnP8dDzo9ze8xeE46DSORLgUApAGROIJ
ygy4CjUUeOx0950lk+9WrC3YnUNggVE3E1fAqKHrGbJO/PD0rtdkEtEci74zK33lUbF3ZFJA+sKO
lCjaEQlHKXoJfMxdwsLVO5i2OS1W3tM213Jmeq9N1tOnpEkiEzt89T5IyfWXumTVdyL9Jk9SVHKO
xgXjhqbJbLKanU6Mw1wmnma/5n5UzjiRCah9eMz4kL2GZVoRGaLnoxNE+mE/IO9h8ZXYAXri/MTa
S1Svc4CLvLcIskbX/qrTxsb74sVRXKNIoY+Zix1TzkjRXluUeKJoxDYaqnsqQPuxaXoZjta6/oX5
qv/S3MNR7RoCLR/hmC7GLfX6iwbmO1m9WhEsFOJ1CMCjwd4Ts3I8B2eKP8+qCld0ROph8eLjj9n2
mqqxSpHSzNOpNvKmdBXWWxrymENcZ2XDUosYF5wbv5N4sGH1YifaUCsYYpv16pAhQP3BmzkylNzV
cZYVlw8opl2I777r6gb+22NdhDprbdr5Xtv7P+KeFPOlOvb1hunhzs4CX2TTgX0Op7kDzAHAwDYt
cb3L9k8rokFipU8eeGwZlcRerc0SVkPw7Iklhz45G2J44loWnOdiAc6AKKfqGnG4Ph+0+vabsSnl
8k3dnvwLpL3qAIvS6NWQxlBZv+Pev0/KxM26vHE0EH7opAVxgfHqRQUWuwtqvOiND6FXO7OKSisj
uFEF/PWebN6/s9C7BxhcXbQCk4PFMBbmSuuHIhmqEgUT91vZeNWSRCLyE6JpsKGUQoC/+fAz8mdc
yIAct4HBnBTqSCoale3u4No7Gl1tEXGKEm5ro+7lXMcQG0erKMBNcI6UmOoUoeiJLu2HtSR56NnF
VXaHSD+jXCrUUOOhWXvyKhLc4J0BW79herS2Nhep+DRIBLnPImZn4ZrDqP99ZT6x7otpr+NBRzin
YfuN2o8JzuS5MUcd8VRAqnVxscvmLpxZODGqsvSxge06MGdtaGfkexmi9ktWEl/Jzh7qIyztSAcx
qfJ1ApioS9DEUirKGJKb6WjbClHkjJ34SU4qhbCOndWYD8m/PTgeux5bI95+YcH1j698vrBJfME5
aHOejCt7N2RZSSBYambcsItNY3ff29qJdrqclMpsMVpKItnBXsWYxpU1YDSIRf5/nwjr0AS1l21B
6f2JSWkU+Cwl1GsKlhlCMcJyR9p8le3RFPcRAUOTgp1asDrWFrFfYpFpsB1r61+YN9js9heOOwXJ
NJbvGfGKDrstUJdeGKhl3WxsMAXGC9Sl6g3Ov95PAPTaUKEFRp/LRxLPkCLYR9t4tM3POSE3BfGj
gdQRx8/M+zOgXkCPRLK+f90jixu5aBRgM3sDKXgPud22Qdkgi9huLDqi7IF7dD2EdOHhXiTyPb1i
WeEeN2+/dyg9ZxW5qlizf+9p8nTa2AcDnnCwcZr8befuXZi8UDR681140VlmZItsDhLlcazCgPhV
hRKh2sxXfZjyMXU+58y/Bb4gwfuwkC9kY3FpBkP3kAr0iPue2Rd8M8vRCJPpLjsbOMZKoY2a86Np
IhrzxIcU1jL1Wu4bFColN6RyLx3XhlowSQGChdepP1Qpg1+Hw4RzPjqQiZRpDpXt50lmvZunbEVi
0/vQ3JxYW7Oe5RRp77UVAiSyBTJP8pxCkJ2EHLuQ3LfALPtNCXZKhII16DxgHydHDhxugSXluYLA
ZgGv79F+IemBE8/kAqP8SUDU9f3VjDqHKop6jJsvPKCm6zbEQj2RMrQ+YKVPPOfz0044B4MNdar1
rI6z3U7gU8BwiO7kYDGHqZ6qpjtz+V1+PIh6DxGlTu39dUElxGbqcxeswypSMJSleVufdAwZjBIF
Z+5dxHfa3vsINiLba4qli+uxJ5PuOYvhyiNG10CmkHzXf7uA2chkrS+z/SQW0DyvxgjYSPIJYXBX
y/bB+eLrRHuPlBBDbRUe9HtuI676oPfJW/td8bB3e8/jEuytouN6zRoEEoKl4Oj47MJOIb+/Yhh/
bAArGFwnoJEWJEcW1qHFHFcBSuS7gmOVmnRgA/1rDDSawsgv58jW98Qd9qq2L93wFlTSLca0zKGj
FOJX1FdspxTX+ZCWlETBk+cBNggSK/JS0V7Ysi5XSxADTZUwVGEKWuUE3b/D/a3BAPiPt2AtGmVd
a3YqIwdG/TRXfHIqBjT13CAeGHLkpsvjzaMUYqWdVNRAyXLdsgcLM+qWX70+LkR1zmoh7mgfGtyk
7nIM1lzZoVC//bFtRVKY57NzLj34RyCCQznva+NKN6Uv9PMwGHpRT0qDTdEWn7LKuCWHp+K2ctCy
fBx6xiwigxWU0hpYHf/9UBaw15uE676LFjhIdqbOl1euA2CBtsuf+5g8pxHsQ5IWRuKOZJbnZrHP
WjHnrw45xOU19Rkw69PqJqknVIJSfbazw6QDpQBWhJPsz+36yjDLFPFirtGAxMgp1nnGvcEL8hHx
fAxoAjJ2fcjqTalFJAzgn3cNydLgOd07h0diLCiaL0NvxOqmT7f2H883Yf63J4pGuRVYbmTu2rRo
ZpqC2qURJlGWgbjVZz1izpTrUgoLYLtV3ywXrNofxFfP+DkmYN19GDLGuYbD1WbP0JegHOMpGxXD
uM/JUiF7YHuXxgqia8B8c/PFAU2VxFx/hKq19RtPMakifRr0DqLktX0/bVwLQAqFcWkzxzThp4Zq
GME51elqfW/LhrvJKSvBs+wTZ4+3lsnH140UgFnKTmyetYTs5sqcyOzjymGLm3QVTLHVBPTlfg8N
/3KtJPTAxmjNy1X4c6WTYvi2F+lxZRso8nkBv3+wt4zMOdbgaOZkHkBQI8EvDQoY2Ly7+1Pas7Gr
vtrpS42IPEE4vTuy3F+pzHMGuSECxrL32RotM6h1C71vl3VysK/5UBbwCxiTIQvAqF/OQPsWEs3r
wjcj52r2Etu0efmh7KvBdvmGq8KRx7/lfPbozPoE2yWuktpgunK4/hhhh+bFp/TpRtmTZr3UTT8j
u6djC35/h1J0p/hEtvK7w/6xnDa2EwlZ4GydVwAuExajjL6B1bkUIXk9/vQa8gAetXcrAsV/UZk3
2W1n4u1rQ7Bzssu3OveZqx6MiOuNCNjbM5KqmlWdtW2x+M+z2LbPbpTe9fWGyvDK6k4jZFou2HjS
v2dTv7KAv1AbIWNPZbA5E76PstiOGQ1pXHTSiugcvLcSrFF+9kzKGOcxjvmkSlf2OMw9xg8Rimkl
Ri3g6EPyc4qoQWTyjzSQ6iBGvwEUJYO9M/FrjDJI+wYPKCwoRe+fcKpUh5otkm/NKIw+aQLJXfzw
4QcW+QxbS9595dKLnPjdUjik3aquoVDvoViFWNJc4/vrB8JK6sgUXbndYgznuJjNBQTorzoorWtl
mgHJeyU6jnWrDomQWrNTQ1yzZIV2oGIrw7Yhgq5gt89Rb+vYVG7JWWD6KDymWk6JSN0hs4XflZSA
Vds8WaCZvhU3uGKjpqujKrgBWnJ6QYbcT8JXQztNuqgvlLj31+PM/N19bJ1OxUus33CR9agtTatZ
w290FkIZhws7o0lMmYXCUkuCqb7mkVEs9GKA1e7YEz9+WyZOPrqBSyz+cOYdyE7eiD1LjBuDvM3+
keiLyi0MiYjG1smO5SgR/bwiU4FcwkjSFfgZdae0ItYZakXo7KRtJ9tztm0EGwq4cyPIAzYQCpAe
FBqefte31lb9o45WIpA5ZQc4I6dkn0Y0b2Mqsuyekc00J2HbGNqD3GRvQkcMexswp2OQkKPJY/lG
pQ707ftGn4esxKcXgz4ejJnpoByPzqPO5twsO2+XryndqPXf9pR8OkxspMg7JSrmVbRgKgZ6j5X+
A2SkkR7L4wn/3AIypi2Iim9jxqMP4y6wOukJyeLOTe40FPax9w2NiVPEtxeVEEhij2hF9Lake23t
qnTW4aikE+b8Q6PIwpVtvGcTTm+mOj3ZB3fdOxD+zHjUpityOwAxrJzUFpab4gKJsipH0yT/bqQL
Ai3mBJGxdWIDH+qmhjBkxC5+U9luKHbxjCOG3Nte95fpk6luppHm/W+t8tV8yQfswLwDnysrswA6
5V+LBxTkJlp0LucYZRCM7av+rNePr6aOmIZ5/NdQKp0phdGAttD+vYF1n8d2l/9qN3c+xr/KgL/z
DlFa4e+LYtV6hUq7p64CVKpVPnttNDZBhw3sHtDV9LTf2Z8cHX2FIQS9vFAiJ04q7WdptIbOS4oo
ikUWHTd6P6gQt6haWrN2ZH7Laz9mkTTiNBqHcSj0GPh9Qc10ucY793ZR0VBsE62CzZIE0xSs/6Qd
jWhYsOklQcBc/pjEt7Rj/zEjpuk6tPL1jeYHeQGy9rXGYUiE4iWXSf0UN0riW1f9hKa/rnDEu0ZZ
qIl4MtNIRz/YqkpC9ST0VFnqXOs7fDaJdOOuXOTAx7tg051G7t8q1dKQP0oCPMnwLPNT17Ji0K6K
3BhaLTXORdwvNRztrzfG9cMI8MdbTLdTKIPJ+qRH43Pn6/930dozzzoN2Vw/PBe0gN8WXtf29dyk
AMLEVaXSmIoh3fiKEduykD6zMj3RZ/veoGDsh2IiuuprHuNoZmjuurHYnnyM5iWoCPPMDDR0FKPF
MFb1f/aBZkLiBdBUbl+lU9gIY0dKO67Zdg8g/I/vtqQzxLgmcFN4VZGXrjjjt9Xnl9lXerMqkMhP
IrFjz96q693PIvdA9U1WRI8jz1Oiggem5Bt1gAGhnzlTcMGDVdSiD8ZoPFlLSiqI6zFRSq5tAPFw
w0dvIccSsSPYCLr0EqXSdPug0OXeJOAc7aUgS1iPTqisA1t/k/xFfKaLWjwgq8iPpC94FH9JE4J8
UC9R7Gcvr9/epSCvwL1GldujlQMuhPuqKACO1NYP9/6EkUERTTpTjN40KriNJuyH+r9REK3C8ocO
GziAG0ORnNjJC7EyWpmYeEyT7umVLGgmbLqqysRUk5oQoWl4kyzaj1yrnPFdVlhX4hTA+ySMAWa2
HQS0WKi/RKBYP4Zal8tfmssZ2IN5bLdywR3qR2ibMjYi7LsrBfIx3XjjIpVngnuWgG3V3qIGgVZm
mOxcYc9R751GTIruf2rioWljxuc8hoeDErNuN8kRPiFvbDVBlzVQTGN8WXMy6H3XTeHl4CIoE1HK
uZKCph0p/qH7wClhOBLhP1nrb/kIoyoE/62jY48yl/RN6FoIW0D8vqbQ9cHL5BdsHn7T25ihFfAv
nqu5akOWoOjN45JBrSCgNZhbqWm662g7g/4kZjsLBAQ++Y2riicsYN0T74KL1fmp7X2feTG7EFxH
zppYxNtqc5M9lJp9tSCTwLKrS6up9S4DothwyF50EOU9OofB1zBsRDgB48HvAKwaElfghR7cwRbm
DcsXcqOESkd5k2so73dsa0W4AumeJMsiQ+ivBU6eP8vi5bdxQWUS8nzlQf3ydZsdGI6WLc/CAn8A
3P2XQ2DiiKWnNmpFF47/63zyVel11WOIsmTsi9O3FhGF2EmPgRkMBit2FoYhUkv90MPiGdqkSGav
LAEzsxoPZ5XRZApi5JJm9BXLhL59RoYZnup/R6N8jbvg0vcW8DtmeQ5/Gb/F14EOV2SGq/VVyL9S
cNVXh/gJH43HVqQKCgfp/u8IJ87BJvsNw4ePHC1cAgwgrIt3oM+D7qmKMA4jnYiKJ9R0B2rw4216
g5jD/akkEpZwVUU4xmR0hT/k/vYx2tX1SctQQ6E+qgeuQJCz006AtT5FWlPkddViBJ3RLLNagcsT
fgMC7AoP194tpK5q/n6t95YTaGRiLRaAEOUSK7/xx4zvGYFR9mI/0An/pGVbh7uvPGzwHQp0573A
NPwoNWNQ6dVZH05vEeoojBSp7/4x06HgqbCQqvdxK+bunbZqgT/5Jo/J18WBDzou/25Y3B1EprpD
/GVjALK+t1dAloH4aK78GlQqSuTqlpGhj9VJojWFHz/6TaSyN0nhKtelLzmjRbh3BHao1RIqeFkX
AmQ4ly/KdDQaCJqz3uiYOE0u7lKPWwz4qCO7/wcgktVLYA1ZUi923bMPER+SLzHO7/sWvGSDBn+x
fLcbwptiAztuj5yVm8hhqQxGw4MMn+gvjMn2J65LDXPc58V7w9/7Ci7pdxUGmV5BYuRA93+/mewG
kUmuiNiMQZdjrNWSEIzT9lBjrcC9J+aKaPpsRO4lzItjy9Dhbgi2IudzIvbw8WVMc6rwTUg1mJBc
IvfpSwjAbpD8cCYdMFrxXczTwXW8Kj0GE+xPXxrLkZp5hcK4qNgndzWCOPSpWcVaRdwyd0dKFXxF
cJ9IXiWZptTpyXUZgk9u5k9EPaKe0iN5dFuNiCMu2Oxe4owvD1ezV7zCI99sZMDWlpi6TawtB0h1
5LCBn/i7QGrdjZWj1NHSsxv10wxg/BI27qAFZ8hq2yu2SoIZ2z4J73IGsHQITmLIFp7q79iYP1vz
DbZlGDlSPNtahtSqQPCbHevVBZjZaRY6MmsKXgQCKgWJnQgVmD8wXiC1F5rLQEMiZSvSJ+kbVXE3
EJ3/H9h3iHndsbGeXjxyJ7webUzByW24142lrpdQVorYF7IpZtgS2LUqT1F945lOx7fFHY1ON1Fy
r9VQ5gmaz8CTg/n7rkpoYdMtkSHyVcCWye7BqShvV+EgrZCpeXKc1bw+1ZNstYLE1aOxYFu2MdgG
EZjl/5Ef0S50EsqkoIzCLezhGS+n7+IGdyz9w83L4qqWJB+ygm1YIvB80gRs6fgdeKxMnEKHNijZ
dOvyUXTiXfvLl/OpOhapmdmBwJ27BEu+VUXSgQoJEjWihg6/bI2KUKJOKFFShbOz8ExkT5Wm8Sel
0gh3gWRIeaU3I7iuRuOsWUgC7W/icXlYMqcfemXnmXx2m0HT4Xr40g+AOo7zhMwgbiGb/xcfK9tj
qWuKxfurmIwS2Cl8IZWouTXlgxxW4bLvae7zcuepc/Bla0mTw5XdlPUhjEjfTELJO3DOCjHTIFir
VW7wEhB2H3rhqKTMxkZrpLpbW2q67afyrSLQfUE8gjok7bC9nosTJ7Lb3BzRNb2QAvR/xEhaQOtO
+HCBRPK+xI7J6tckSIQga6uMdWETjWp+H2WdPV6Z3351/uGuzi0i1dZQsB/ksvgunBIpPrmEg7St
RvGN8Zyxd1LVRkgBEGBEk35PibynOeAg1QLYHNB4mTaPX3/dV77Czdbuk4iZkz99NPOIZEysAX6O
ep7G6Y7fngut44vJ2sOPqrFIUKcF4K/0Xt30cdWookxNROwsiRGmNOdz8HgXUs5RypIuuNjVX/6/
M0jbmpBGYvWs8ZWZyzXlKfnJ4MgwMtQdB46agBiR0OsNt0iT857AUbLKsrrKaCI+Yy/Zr0MqUYlc
1oxss/LJy1l+NXBXWpqITX8cFjuiO2reiMA0HoasaQZVp6wiJQ5L70WXVO2rpaWpCmndYYnURizS
lWp90s/C5+oYYy7WHA0NVHOYLm4+r5sJg6Evoh98Lubtyoxc4k20Qx9YrsYkTTPaM3OGV7qVGY4a
6+D8CwhjxbkYljn9bNzDvf1OueFc4U9Nnciu3ocGFfVfaDXPdb+Y4pMsjE5E0+mJcVwcLrnCJ7uF
xomj42z+SGC9VD3vOFtKktXnfbEP3OF5/wnXApKCF3rpOK/VsogcW0CeLyWJAgqucf1oUVspILu3
F19eDA2cmu56D23IKD1+zIZG+6K7Wwwr/+CQ4NJzDuo4og6dFKOmt/4fzPQhGChQogBI2xOYv5rk
WSIJz2JvQ3p5rVeLZBho4V/rbM6zfOLKPXfmq83zvBlSo0NJ+paTo6UVRhnhLlm+lbfqJkbGHu/d
N7jY5WR32ZOGfBHiC6NU/pHE/nmN4yMmrs9lbFmawpjRgH+gSZ3fFTazPqUah/yOX7kCD6cY//h1
Z9ulnppdySPgQvgXDuvjCqWWYcyuGQosYZBGHB0oOXdYc9vsAxMQrtBSacxcrwru63VZ7f1mk6Rf
bb9EzS4YrFz6SgK5zwVzm4bXz9g//TB+f8yO67GqMvdM8CjVWeLNDEvp2smVedkrF2TNcKF/arWx
gr3LRsrBYS9A2Ehmh+yCKx4wQEoA6DagDFfSwFX4hLiZx1kVIbTa0UR58jfYvAS+O9SXmnUi0mvK
/9yQ8e+wRES8lygf8l9XUM/ltzI+Z09tzY9SFzos8Cbud2UYMQa1Q0Q+Um/gjZRLCGAJZijoWJnv
TSpcozGk7ptI3g2gwoXrvrZNltEtra4xtFkiI9fypxGSEEGzDkdaSwENpk+W7aaNV5y2UV54W2lG
BxM5DaZYokSde2fz6pCZzGR5Ob/Uy3KbcoC4b7sLXm4XWo2gkkpDoZ2QkPqj2Sjxtrw51i/cPQIi
YPI8fEen/REEk6/YTY27eNGzdM98mLvThgmgwbXh3PQ3k4MCJHKFIfpo0no3k1qjMHx9+etQ9xAH
sItPGQG7hQPX02IxWYBcbB7/FeUmawPHUnKgCYGNgVwca9zGbkHDGya4TCVp4i3H6rwDvVmF/zRR
qLvDJGdm1ZdURFrZpE61rBISYw1GQjLrtVFvXwwv48Bhl1zEtHU3rhIGG85CqwWNpQRTlBRV4llu
+u6SC24vej72f07gAxWAAi6xFWA91WALlMKEtx3Fp1Hqbd2emH/A5hIyicBfoSGkrcPdTTj8BJOY
/ZjUqPzZYvGrOt2qlp2Ei++sn7tawooADn3i2Hjo4l/4AUd0aPKBKPHkyUgcwzPAC+fWLcREr9NF
u7H4/3S9gP6wTBceEVNFhXD8yxbECoBpXAd32bkRI8Wm1UqTb1gxlwYjxYIu5jHYhPq3UGYeVtVq
ObcaAyt5hpecVCF3UOMcCJaNbX3aLlhRAxzFHJphDF0D/eN/blmUcSR88EnFTQIVcpcbpUlveL3X
eW0C8WOFFPUIsXM5b8lC1BwScFE2VhvQLUfKEjW7O3UQi754JaSGkJQEywTUyEGKUnIpj+sprzI8
+ayuOv+s0IIjfBwSa8bo1xTKnR2zB62JZWubAr2jXfbb/79vK1XwcDtM61R/i1F9sdW8/B5FcBpO
XxYhn1Xp5TxuD9soMaciY7+dQuWEcyXr8Rx9IAU+NaAA2DtQI7amLwpUwmWN1OjQuf6g747+cOyk
oVmx7DP5wvRCPk9tdj19J5zlPlgeLTb9fhFSaNGlAN96hzhxcv+K82RHIYyWzF6wdGKAis1BuG1R
ttWAYohyxkZD9uBSMSxgqWy/1XjMs73llqcnyrwXEoXvvXDHNP2T6wcr4hLb9pAiMJw8zFrC8Cqt
1ry+EtWXvgpmao/haS+rmPQ4aEmbDc6g6ieGHI2YdTh7H7UbasVVZGPOiUmydXDhCPRcFVzNxYNd
hkkSFywOqTv23i0ZFmLL1CP35yIS7ErPxEkQmUIZIaNvzjSw/dZfyVwcbL1+lMK6Tq+MGZsvSprM
V5Rt48DJsj+dyfDks/eYhgnKcVZ/VOX37AxDYLtXlqf+y38hf043hYlCm96tQ2PVuRDIOP67T4ND
KFlMAWafuhaeyPROgpG1cGv/CuMW4GIsVHnw454WWVjwBKksToWV0BAD/Qbkmwglqz1SuzDajQKM
DBj0R/gE8Gdg9xq2St1jUezTJaB1zbNw28hFECc/tYJaht/tCE/ErlKOS9H+W/k6kETOtpN0VANH
3UHCtn4B0gynvWKQRQ5LHsYOssc0P5pAqa8yDhvDG2MJyreVl/LXvfDlNagH74xXWIfHmGp2sg0+
t94Kfr8LHFB3oV7qT0qeZJvXZU2T8QYZCHsnsidhp+J6UR+fIEQsuL6jhQ+ecoc6k6SibYvJhapp
4A6DAF+2Gr85kezna0RbU4XkSUNr9RprqfCB3SZl8E7LPQS2G2rs9uoshQVacMDlnihdV3Xg9hUg
ogAcWVxzaANrR495NGX33RXgyCW7RRgHOX/VVITGyDm8x5NkKXq0tC8BnhnGcyDy+CrT9mlLPGqZ
CH+KTN/CBRL6WgmYeUNEDOVMqM2PxneHy2p2/t+xNV2dGcAbk7l3ie8FoDp/y0ii0s6UlNnGapb2
0S2aJA7IlP0VdF6rqp+7fmNhECC2bjJ02samIcsiJyh7eCP9WyUPWrI7awAcPBHSypP0jkCY/N8n
8KjxS7SlALNUsJBcTKwxt/KmvnU7yvk0U2JKL31XFC8nQMQChW6Q7I9yaUMp50OmHBL9+k4YH+8s
yBR1RJKRWe3OwhH8XXwpH+6RZW0sEzXz5HFZeBJFabLURHoqIBO2ZTbWoIAg2sDh16O/HwIXWRpW
i5OB/ISeNe0394rWUyqM3oC05Ug+mrDOQB+sGwg/XloxBOkX8ngw+MEHDjeGwCa+CkM8ON0JnSyx
LcxwwPBrMUJIEKh+Noxxz/64RjDJeviuaEb13RHGAZFucv/1RMQcZymlQn2Lq/mrbozQLAYe5RWW
Ayo4hjQpQtwa2NSC7/v0ybiLv5eaRuY4/ay8WBXZw8wEt8RDu29918mgIZEPhgtI7Bvyu+wMyDTg
RD/uG5vWM8S15QXcsMcW6mIpmwUMLZFCEPKIFXt/r/PnHkEFPVrA74c/kN7yI7yommHtPbyUWjU2
JdD7dCoNU0SWgej2Ia63DLGPX2zBABiZSJZUvZOgeFDjQ/aDzlXoCv/4TmNcgSHgcsC393guAAOw
99NVxfJMVrnw5eF4TVXY7/R2l0IZpgaceNG+/69tylGd6gOxzNmazH5rV15ztMWPFPzjmzo0COK2
Q0VIn6dB6G8E7WMeAWyDoUwXT2+VwEnZ9bXYidl52fiepYLxcDJm+bxc2o8FBzr1Bs1QB84zxyL4
795SLE0LzyPxs/LyGiE5ibVs1LPsP6sjbWaavmR1J0pqcGnFULG/dHCIUzUfEtC4ThQjnMiBcaPS
rnLmtN0jL/HusdmmkMKx8jv3KR1yzRzodeN88rrkj/+H8203R/i15ipnkcNyWrQd2IJc+nNYYc6O
EUElmgpo30lXSy28QUxTwEQwQoA5+zzZCYnxCI5hZrkxqoRUD/I8rqSHVEVuAObI6XEXNFcJoW7A
zdvMpF3y2mmsMgRdtRrjTyvfq452dihTfWcuNg6rmhooAdVH4EmtHSpeYaP7tEodYqJYv/QFB2lc
etJBUmHvZnD3/67E5pwSjNmMI0aaTNJzhBIK6UYodPaBX7H+sVsKBa93qVhYZjDdGo+6eg0tJkV7
KFzKk/8YQ01WdNstgALd2Ioh1wbkQNrI9mEWYCilLqz8fQdEjD0fCZAQooQqOTL+E+5plRYMWLlh
GxwYmjG736hbWmifbWTI6JApv2b5k3IuVUmcznObC+fk4aVuoAHWQowPKUzTBCcSfkzXoCSu1te6
g/6UpMf68LYMtjnbmdfL9Z0IgmsvaXgPJH7l6ArwWyfXd2wEoWHNrFt6dInqv+7lyUCN4DVIkY31
vLGerksraqR3Rd8VWeVpVSjRR5NpJvRNQABHKh4VJZYyCl13wjLAhV1GH+oA20bqOyGDqBBMzAyD
ppeLMRovdmQ39R2ffhWXb3A/BmYIznJRrRJ87KRCVtCr/Ono2kXgHoJnm8JBwoXCK7YK4P4gV9pv
Bu+nmJd/BkUPK5f5DAuqOuawJkUeivgw80hj79E0AljVfxHDhXJ+1yztvkJHD6i0UNH6cisW2qou
r7UJYq+n+l2oDLYX8+Yh7BvB5aUBdJl6k7XmzgGpnRQx+2B4kpj1No1YPyMGcX2rg31XyxxuBice
sNz27xhYuRONjxh8O/punvZd/F5QNoGtY0n9QX9F2GTEwSh7UZIuQFe//p7UBd34uefb6VRbE3X2
Dg4LnxPGslS31MpAKaNE5hOlVPKSr/XqBGBAV920aMNt9pqXRI3TzJY39yzD+8fACV9lplkfRR4s
VKIP2YFGGjA6fBBmw34yXvbU3ya1ITKEQzfrV8lOFiQQRQJ/d2Da03ahvfpLBKQV/iJwa9MA5tqp
YHWHMC2bG+/m/fbqgW8r3Zc5pUWVRnjI78sSDhO6XT5XA9P/Dl0ljbQEtAGlP8NtD+qXbmo4h5zQ
GMfkeXiX3UoTjTT+ossYLBv483c8pR5T5aOMY5XUhArpryruL6prN5z9QZyvr9LDahhv5GgAit0o
lvW3w5zFsAVXivn7zfJKNM+MUHlEmzhWT0ojX1ulgh5uTYeoyuszLbJOQtems4XmtoWi1ryif2xp
rsOnH5dXHPX2RwVeUsQcP1/P8lITx/YrZdp7PtIkCdM/S2ZdZdduLlKyh2P9JOicX4+mzGk7oXvb
68o6vIndC+KtlGrIB/1f1DmAMOi87b76SxP3E3yU9CtjAU7WyQjsep9lni11Up09Z+XoYdSely49
PIMvSxyNWSk7+gvQcNemBb+7aIZMzP0cQi2DPnYhixZOoAoYoelVkTmCsWlb/UTy/668YzbgW44Y
TAA5WE0/BFo6eXa424n9ksnNQY4PEzTUrJLEzYxSL9KQ4VFUIN63lIXrKqHVqeeh7In8telJQr7A
feTuVzn0nxzSgkPOcUhCEWS09dCtFjEihygs4zPED9iCiUBMcDqQuYuEbkFNqAQtUfqIaqe2Gmkf
qV06CcYWGzXriRqz+CwNf+aTu8QfA6tdluwAwLxxaOF1cD/AN3jkxUpOx5g3o4sKqWmxslXgQ34d
fXONotuHeOyN9VR3LbFE+yQHTUCJMbcChpYwm9LThnGqr6dXF5NqzB87JuCYAoIHlb+AuQBH9Wr4
j1P6riSRMVCr/elRnaQC76PIAxaw/l1csqeAhdjLxKwlILcC3TTrLqrOsT2HN/ODRWD33FvJjiXS
H5X7i4KKKEk4BW8oeHC5k7bH1PUPN7CjsJla96Iyc7M/yshhF8YcA0XTjJ5s6ycnITM7thH2d3h/
vN6xtH4t+RfjNx7xcxdbBFU0HEYQkReziez1jojVNTGRLLtloNCu+IbjmcdMIu+CwhfGIgROZJRo
/UY1ubtFDCPFVfE/5CKQhvow+qXAYJ+q0zDEmrCm5HLQn05AWwgT/0wtBhjkQVI1d6bHyVcSjtXw
IQ3/nyeZXuwrUz7SU3oBgr0MdJyXk5ijovoxJCm5ea/v7HjHL5/hHnlBin0OfYgWa2m75lv/OXGU
dBgH+KrkZhEUscVOr2WdPPr9/rYcDuY5aWeq2GVWIoXM3w+ZQ7+ltseNraF5UF5CBqMM8buAtKiv
qnPVpKzPvrjqJOm2DdxYoAP81x/nX9NZ8pUoSQPWYTXvkH49EI/WnOSvLHoWy8MoV/WafXEUQr+l
2f3hGlapCoqtvBYfGjNxItEJDQOTkNEYaxq6TKyF/ds0iEYNbZNEVBR0AXKUvjiUCmgV91mJBVAi
YDFxiyqL1338UbrEvxEspaA+pKoHv7Sdo5OzFB8MTbYndQrkyxPDnnrhhIdbJG9wnfsdaY2LN5mg
HRQZ6PtTj+QjxCgKnqGIJBJhY8ajVfBxmDokyEKd+FUQ/tmfscnFzH7J1oEcXQvfQjBednwiozNo
goRdseRTkhuBF+mIw2orbP3kygzgqA2icTWEHORQZDt/6r80hKrzrTRa+6/oRKqf/Xe0gzs1qF3y
CDPms7qLENEz9NPCHLCRFuqSTCaBnZoLDulQgsj1y2RlbFfcr2kAxE2FuZg1AAV4KM4I86+RViBY
v90f/BPImhGr1AbssugAGgev4KavHIr98v757b9vsk94Xy9J0Edm5vEVH9Alu9BCjCvTk6KbRZi6
t3NjGkPeDcmjuMn8e/y1Xd6Tpy6rUWaMfFZkcgUmtc+JpUuIEopps3e4cUp6rswcuQt1isyFUwrD
ob6qGf5TPmUiZkflQQlsr7rEIKJL71B1ZLzFAimrHSE3kYGl4BEJ1W6PbWWv6MwqD4hvxanNvIgR
Bb9BbyBWwYHq10zi7W4RJnGjHUZcbbyymT9M7uTPmAyz+gyX5dsqdCCtU0ejvJNBHhsmpUxBzA9j
j5ItZivJV1q37vUlrqu5J1auY2lX8Fpl14EEUt/wmXHnxYBwo7u1xMXeLvd9EMFS1G+SyQ2JJMJs
0vkPX/SvrpQhPeTe0Yn2BMeJlqT9lGwEaj/o5Zo/9DdtLJjjSysCuTRhCkbH9siilhJ+PXuc7pFi
pSiNKGvvjezx2gVrOCEQJCv9NDGAW7q04NTy7UWYVGZfFjaqO4yxNv16ywNqjgVnRCVTMfPiM/tQ
DbN+edx5pDzaAbC2BJAsHNdbsW75oQRfkRkvJwvVw+19w91mD1Otk6t15O+wXyyVAzTf2pdEkJKo
xIOvVxHEXrwped78/bWgnhPNB8M1+eWF94CYVhlpg/A8Umzh2ArTCtsoK3mUtPDB3aKNVxcmJ0HW
Ypy0iRWlm5volujD1dLvfY78N8IgzKDyQssUPyaPzm5Z8HtXyM1u0XQLMUBg3f/jfFWQdtoLhJbm
QDQ53nRXG0Lm0y/vh1L/cr7bf7S8E8gzaAzTMBu7uScmsWv1j9S9kdEVvGJH80gqwBFaIYGqVZRn
BwaGVysMNtxr5FNUhDwXYTKQCZgFHnw+MYIJeUIZa5GI8VrySiYKK/JGgPXzt6ohZKp/3Oof8JQg
gavnJ3BfvltAGO8fZnrSgiAAaqk5e3mR6df+0lLxCzs82yuHFFob4gYetaTKkMhXnpdkxQ0QqB2g
K8dhhxM+u63qEJSOmLP0UcrLf7GHlJyz2fXZW0C+KgfSLd1vdg9/eDlSJH87pbzWa1dtEwOiBBVO
AdssV/oaZmhFrB7yIfluq/YcHYQ+WS5CqQoT26d+vnOYpk+fG2V12tbanywncmCQWJ/WxxEi44iL
sUWdoILoFtDWH9wJwa52bnSiE7SKyhfwq88jbrUGLMX1ixs4rdesElv9PFlmPlEvWwcsuUyW8PZS
RSddveUZ0DUyRCQ6FecokYd9p5gqRwrdESwq9dpob6Cbbb+xOwrNqzKvdYHNVcrFTGqFlOrBCu3m
3mDHwgkALmXl7GrjB0670Le4BoI7J67yCUI/bN/rZLi/8JktPLenu3bMu1eWaRInkWtF6r8ew9/u
T1chRbFtm3rXCWfp7r0UsHx4wpR3RhGeLQWr+922UXwcduwQU92D4ukl1eYWfCB9Nvu0W42mAxn9
MQ7mcmBmNNcAL0QSOMLLPXc33c9yOas5cm0ZuEcsCxIRd9pP1DCDumS+fgYIssXq0R9/mDoPyx8e
o8So8FdamS964f9eB1MW37PMZZCL4z4QjsXjCmBrqXescoZ283yqyZHMPKh413IvNK9yjE5uRfAn
wsXjSYUXy+TcizNZV+xLezoEBnvmaHdI5M+XJ2hTyxzyxEeLcrGL5N4/2PYT/pTpO/fZi3Bhbkox
MqdlaGL1yXDOPG3LVl7mBUEzuI3GCQGVMs0/110hFMF+x4/22ju/JWiVLzYdORzTykSnWygDVo8J
AirCW7oHBX2aThXnzMGHUdljlG2rSjF8dPs2wl1fVsQUhetIV1/PGrhsN3rWBX3txRGxhkj9zcPx
Xb7JFreEcj0sPJsc8XgPPBt4PJzPm99IEQ8GrpAOHNvRYC5b8h0zz2oc6PECgs8CxhgdsFCRps1y
h+jZd9tKIngWzTqZiCfkb6nQaOJ3MTKZXoVSH+v+A8jcNW1TzbH6uMqGImdZn9EZ1wHTNmkryiNf
CHTibqUh61JjrWVJmBrxK4vvAdcKnfuTeb5dcSuZ1rRuDAS7vz6Q8yfAajawt0KwFJsBiIwPLBdI
gKdCzsaBMX31c2NAoLoG8/S+N7/Sq9w/3/7bxEBQc8IJmkRfTrxyaumLLKhb0TzmhBmrPRtM16Uo
bLaAK8z7RiYw1kDUnWGA5nqr/zWVUtfR5CaijRgrbnX5R9VokvJSfMCvKBHF7sFJkhpPOLdr0u//
wCjHn35bl3Sha1l3kFmRmsPvOZOR5lEvgS+UaPAQ8Mp8szYRMmeaq0okvKjbGW0OZtK15ewWXkI3
hq39dQfjdRwq/PwrHZgcoANZ7aNX0d0BXMCL44/9hTJQg7bCSC/k8UeAHJ1U7gLlh7UezI+d8n+d
uf/r+tygbc5F8eD9oRrtxONUgnlx1c9RemEHV+p8RF3enZzeMdgC06SGmE3sdhlHzfqfdeyBNYPg
rm5mvO9otO1QemfYrc4gkQmvdXUeKI4q1GnHZWy7RK/DtGIPhKTurtSmZI9pqMlAHBhX6r6t1/1W
wdZXDlvWh+jYSqJJVX3BZ7kFCIkuXKZ0ZOIMzAtrShb4bXwrXKrnAG4N2GXR2h7x/sIY+ywLXZkc
C/uFk1+Wq93h83Y6q8+sB+NN4wCSQHblPHzjTJ+mS4a4IKZWzvh55Iu0w74OGkQu7qauNRIq8HEI
cht0QyTHokaKQZ+0nrS726udlyCXsceFtLTIDt9WTV0IHNES4AmrgDrrfovVVotsfzfZFPamKB/2
3srXVlRrCYD+eljZpAyeMQlG1sgagZhIxfPepEE57g3yTBQABz8RzQg7lHmR9GnAMblufyvmldbB
83nT3dDMSEKWXjWpgxYVqx3e8Bsr4viKA47QNkLZR7JeLnwFT+QJk1zE2h3BzDVPRAWOuDhHOeIz
ASWE2UU5htRsQO5JIBcNxaNISq/ZOPjUwOd+7F3Xe+vF4JEK+d53TxW7Hr0lSCDrwkNpZ7Ep4fPK
3e/41A64NbwGFfLQ2FTiccaB/N8zIzIMglm14Tld28tXhBftkzBrjxDEWGZIMBh6rIaJ7jUMWNRm
vqj8imFHpuBqV1elLnb4bgag0P3NyadivUE48yhwmxlmXPNn1JSy0x9crAnrnYMnT31XCxpfBVl4
JzptI5V3rmfuw9FmoL3tvF+PixQ4sGzxGZ3FUWVE1zxUOlMfEB0DDI6G6vgfxt7z2JME1ctzM6m8
FwMMOARQqC19KXMP5oghlSSFj/XW+6U7OFKST8VmcI6Hgc3sUQqLJFayZu+IXekmZzVnp3ANrUQq
i8wlq4ikUmNrnVPRJIOifG7nNqjOAwRhx7e9J4Igatg2mCv2RyFco+eoICdnYjbfNsP7jUcHp8bc
KFm26iibFZbYLvjReHTLjRsBL31jRh1nqHpTYh8uHDmEd3vrL58LQttNWWR02eSR1L+Bq42+/r0Y
3CaXC1J5zzNW3ish0bNBYZFQgxb8p2DoO0boc0b/HzWCp8vbYSYZJFbUKfw3IYStTtRRk3pOIxI9
ZjoVIEiYy5sueNXOVVY6UxyU6kNp9Uxcut9Z/6RReuxC7Bz0OILoxEBKtpXKzxepzNYeQzQ+aryY
I5Ja55oMQuJg6ZHv0n8HQjiz4eeghjRnR+jj3fgESg61I7YjI635Zz1EWqa4UsRxbLg3hS4AIIVo
0KvehChrd1WqNPzUa7kloYWnuId2mnhV+kjJIRPtjZwxbr+13RMbd0aHdvYg9jsaUy/GC2lSnTCh
gq1VJks5GQbHPFNJ0XTS+hE/k0VHnN2wmMfgiwaHxngdQORi0gYbzcbwSbe1pCGRCV+gw1HM1PG3
oPDVF1wjjve6WXycVxNVa2axpwtH4iVx6FVTDkvpLxz56NNjG3VXyTO2KjuVBAHBfqa9RDbFC4Jc
8TK8K9iXhSa3eBsWopoTrWB06GbUQAPsFGMC0SSV4GfqzA2Xg+eBWhv34P/MAAM34ok/kJUclEsP
nO9kqwwqBV03O35wjXQzEQMHqCR5GX39tojnlZz49I+keTMfqcun8e1ZnvnDYMMkgD0VtMI+tRn5
OQtY+UJUP729IpCWVwYj9EDc0o4RSyJ4Y0vI7Pp1PPZle1/XV68qYeDLwoAOeh+UzXtTQCZnMNSw
hYv53pE63t+iVyoJER3ZL+2124SbQzRDHZSyozE847q9FzWZ+dD0RpM0m5tcrB2Hx/u9u5g7VBuM
KY0tuvcr/ruEZe12mCwzWj/XxltXJYEnDVuDPxc+KiCZC4W9K5yqFcBgMDiE3AtEv+oSh2Jth5Z4
R9u+ueHELppjSSeTPiSbkdWPetMcn92xeqdOYW8WhPO2SNhSERyLL/j3DqdXmXcCoCqt71j86/St
30MM22Pe+kPanZu+SoZSM/sx+3jCth9Jip1x38zUBPxHvapBLHgqughSEFAIXXvIy4loG9iVr97d
oq9LeKR3HLHY3A39rrGF53odK0oFiYIWAKm5PAToTYuvlmGaoFc5VrS6q7SIcJ1/G1ReNqkN4Wo9
RqZrZuXJiQAAzj30z2HFR/grEAquxhOg5zbTPFK9u4Ict54ZYByIigX1kzCJDk2fZhC2pFKbdy9l
8Eja6JV0HCwp9bNQgwY7OYb7SSwnDkWL7V/zuvdfkvJFU9wEqnCIfivw/R5HGEFzbkxD8+/YdGKS
e5vlgCx4Obbq6eeqMLkpwT7sXvKf8feKsl4g2oggepuebRGBb6CN8DYHVINqO6Hn+N53ZDDqhr/5
t6cZz62gjaEIfY2wkMoY8gsofEVjX0caPCMI1x6fBxHecPghX2iVxKJjcMJPjVzoRkkUYc7wNu2X
/1oWuJ92IWpqhGEpLPhsdT2tDgcowN3+r3Ys7I62KcN2Zp3vvsO4aROyfLc7DuikPF7t+ZYkzgG6
MbX9+wmgcBDFZDP/DAumL32f8UyjTEP5kfzQeoy+agWF75GUZ2Es172+Y+kYIdfisdpRShNU3WUU
neM1MLC/TCnT+KeL2uO/DIryBtotClJfkV+bewsNWj/er/84amNmlqYcKdlw6WnI060rePInTeJz
d03PTIzqDkhWMQjgWJwMuHtcfv6f+eveC+hvAE4vtUqpuRXh251eQHkGr/1Ne/XVcrdCSWKFZmJN
LLpBMw543t6ilqc0IBjeiQpt36jMEKlWC0lMRNuhVbDffXzuLoDMG62wS5pMZNaooMBRy1gnFdgX
VsR9dHRDxfQITcXl+pFucC+XU7C6S8evWzWCYWKrLuDFhilF5n9BlLXJ8Tjs1iKMFYdLMOCdA5e+
8d+iME+zxcu0YZEemC8Vnwl+vMIXAi6FjAPxiYQPYt6QXC9B3fyZ6oBVf9DJe8PGHK8dDjgFtxNr
hD8no6H1TnKQhbIMDFfbFBXq4a4H8sprrOPsn+A9ecDXsLlps+7lhVO6pgeSfuAQmoJ8ndOYF6q8
v5ufdObKMXJGNP27i0+b1JryEcPMbwfgXTQKqnqxJL+Vx4r/SDdkkqFRZhI5tNNLj7tuOpS5wZXE
ySU7J3+LJlNolZ3IBYT3e7sBEI558rffQUqICj5tACNQTgGj5wTI4kCubCPgeKA9NTyTYqToMnCy
htwxduA+HignqzyH/YDGsChnuNignxS2s7OAWRePWB5OgMtCntDKokyHT5NnSa4fZ5znrln9CWtc
JQ5i6syrY9R36zKC4O2mwa3xUpHMPOv2XwCsCJeghmAIfC18W5RzSOFNY6f2RGd321HSLnRabNbi
svvMVri+n5djpciPJjHNLPBOg0PrgUVlGzi+aZkZy9fwuTO5nyP/NRgYKnBrpbDGRkZ2U/cNcndW
s7VsLpUM0jCEb6DF8GdHIdyqPe1hCVZdqn3WbyVnoxe1j6mYmr9w1t4T6TgeF9Nh5GKetY/nxHu+
fqMo5jadVJsGxjVK00mISx0Fpg5jBpLvMcHuR233lqhipnIrohrP0NF8hKvcn0vSLCknaWl4IS9U
cSVzQOBE/fvhExiwaKPFvdTIVeRBQhUPcJohanIqqFTesX8LJ+q8w45BfnZynZpWbihOC7TD8PrK
9RSlb219yeCP+CU3rRB1Bln4Clrl5JTF3g1FbUxH5WEYzAtyG9dLZ8ApzNZ2BAPOzaQVYp+aUahE
jhxg7j9ZqIAiHWf5z4l5l2CE8ghvByPUIF48aWQ5z0PlHDi3VfM1LbdbKvNXnJHiEO60kMDdSQLw
ai0x/JSeBN1Yy/tPAAUK29cvu04y3WaO5yyt740NeQ8NoOzY8fgcFFCEvNSoDRLVMDIsYnfxSJPx
nBpFpyrvAzI4qqjQrZqtlkM1McKziHxOHuAobDK+J2Kq79Knhxhtqd2oqUcz0/Z9E+4WarbhkIla
SZ+zwi3lS+EplNMQtI5mH7e1bfY8Zn9rrd9c8AhJoFumqtD0/GJ6N2smPTjYHpvkNobKhiXA0YHy
5mh82ymSVyrWHBqiTzxtAVjk7q1ur4qc1c45weMsOGkqkTiqkHWJElm8oKVcMep9GZMly1oWq4nH
FrzersFliG6M1qJPkRVLDGmNnqjCt8l1NP4YwvSUoSBr3+/yRTOFD0szkT5+jwJ8mtldyo4Cb6fi
N87ENXvHoUIrZVeW452QGGuEuFRV5sCAaeJeMswn22mHth47knkof0hi3fJoNWypaTcSd0Pu1yeC
gOijmJ1gwVYWVhpT/TKLIP07wMv6LnQD4fziJwA1wc7eqKHmnmzV1Z06k3TdBLqEEyn4qmCAxCbx
ZBI/0YfzQfDC/iero+BqhzLhbKZlKyYiqcxil0t2TyrCWdpUOT3dcb/kTimkFg7D61bCPI1odQmo
ql7a8ng76LCO3O49VaxypYV/cPzMX/LpRQTA67F2OkQCdMaZLhZGe/FKC6JHqKHYVxrmGc0CABE2
7ZJ1IJZbKGY6apWz73yUCnOJPy8vcsGK0z2gKJiNsMgPI6SV1yUHO9WnmmL5hiSQJd0/pdsnwHru
CHXa1m4KCPTfAvpdpADD4AH/wGYypZWQd0p9ndKiiM+QM2ZfX8U6Ffpd5ai1y/PWGRTU/8qK5d/r
FHqQXHjurIDYkf9o7NxlLINW8N7QwA+mvECoRxem1EhW9BnNkM7Oxsn1LgxEKwOlmgWbuOMz1pqZ
c3O/uaCK5dCFYn568q6IyXtEDKTRWQPbh7J3WNx1KbVfx/jjFV0mKhk4rXGE3apnq+4nDCBHwrhq
Wt1ryeZrOWdVM5wT0WLlcEx4pvC/ebOyMAsbXR0gxvpT12z+RjzTNtL50aMmlscMq6jjJQvfYxuq
iPT+MNKkvqgDGJj6NeRgUsVPKsIQinxorlOeknGoFcRgsh0paXm4fXskwzVvxqGoL3DwmD8zLjR1
DhXqy0DQ0V5M7eKtuoW9Z/n85ZcKm1U0tQt+X4aM6B3tZX0noVm7RYCRhxBb4gsHts100AViCHaJ
S7Bzjcq8QUWNSCgmhumMPHbBCVqmCuPK0noV8VVYT3yeYUyFYUmpZ7fI/Ksq7jLT8hb+mVJrK8A0
nlbSaaoImNAPMa/NE0ND1St8DRbRwHN9/o2XR+VZqDFUYczvnaO560iP5IhszsXkR8rYoIHMzWER
95MOSA3q4+bZV7BXl26HthlT95WIImF8fK2cWObv3ppXF+UBThUBzReZA+NrUbDxrA49EV5pBW8d
ysTMt0wqdFtZTZCLOia+W1UDIV6ad6c/TrS6KHzBioucIniN/52y7N+/2wNcpYBq3N/wJQfDRXCa
zWWpcRZcczWGseJ5f8E8jne8Vns1uXTT8hs3NPI2ilkSt7kOV309s5CMdOQVvGrbLshv6G5PY7Fh
quSM8VKHWutSDoqP1/qLKvUIDpb79E62Ex6OTSwqFx96JlrKioHkEjPopOfrULRbGU/34jlP1V0n
fHg1fSpRWR3EXezTVRgyWfy19AHmnVBRoFZD5Ptb/nbblYtGEFrA0Gn/fu3DzoAJ7av56nASI9tN
UDCu0txmCF8VOwYTYQsUUMxyYqVONKQV6f0hbL+NMLhWGWPjEmYukao6At8ri9KboMmXzOmVXKuN
OryXm9Mz1gC6oP6oGwb4sXtwVkZqoxBXKJKkF18eggWWw53GN75y9oWWGLpSodl/LljzngugLcz2
R3t96644zQ+28Ixm2KUd4Xm6vAYc4uSVcAXHGnKbAhTRAuHgBcnVFKbtQhhlia3/wtEiee+SHvaF
PakEcro758/wPKmxff8CzsuOnQiiuAux+sSJNh4hAol7/dpQdw2c+jUhbRZLPglZzqfJ9CkGNNEQ
lpc8iCS5sk1s7M6X3DTSYH0GiEBc4ZflOp6rpD0nxDJgulXWFXeMWoBzuOh3JbmisIfRoUHeSW8G
Hjyi/62zwDYKpAGZMXwoHMOlTSkvFJoNZ66QOTYewVE9/EblW/Em8k+niE2mhjtFWQ6IVd41WfFW
+71oBWFSdeIgUzj6MfzlLrgSomwxPHtUt2DQAkOeUKpDt52g1tIZ2lTX3ss1wi73mkaQfSS72lDK
CduzmWJhYPplzhU0t0xOM3aMKvzWsfrUCI/1xy56DNU9vuhAhx7Jwe3ARjFQU8lsH+VSpJ1/fcVo
lyTUdC0AccrE+boZEdTN9sH/mkL2P99E9Q8b/NOlfpgYEzxLU7OOWJUrv7YO+pWKCuWCE19CTP83
3PySH2SJSo7aW4RSTu4qSIIdc2MStXV7IajnnzjJotQv8h4+pIwKlbw0LJPTPupmMJ8GHpY6dtJt
Lm9FCoydyE+EJEpAflaWStLavI4WLb/nuTaH1gkE5EBCdE75c7/SNt6Nn0d1NEo1/k6kBLIJljB0
COr+zwyesjS1j4eNRcLtNkBEUwbOAx5jACzDgDVgHF4zentpcuYaG9ZA0mR0Mmjaq6LzSxvA1Pti
K+eUdAp6/6YvEjYb2HVgrJdWk7w1xMPuxA4sT5q4iAA1lLbNPCYoErCecYZEm/C2GvJxAvTn8THz
IKhEbs43BUn8Ws1nDdGh/TH/VQISFSytT+kMutKJa3vCdzhLBG7kTWJrHlG72aKv3k4XJ3YTMcC6
wSnZDnq2eWg755dKdo0P9Wn10S3XxveUkl5O0mlMffDJogmQeVg79IPWEcdmMhZ/IhUShLhuHX9T
MKRjEYQg/Fz5Bqq4UChqThN3GIrbDDizfpGO+v0EKJeWJR6fbLA78VaEKQe4newvkwU6XqFlXoVE
hjwWtvjqAaOGXSJAhok9zla315/SRgGUVUKFYhBGvDGONXhfp+A+EyGc+YrDdmIzo8PmtcxjvKWD
40Yx3y5DBwEgp8AU7NrDE6gSz7fM9+z4LulP0mddHY+P2ljqMdA5gIRVZIt/AZvSBaBb5Xe2W6s3
DJIbrO3TiEJJHb+iQc6eWin2byVwvmY3FjDFTvCciySSWhcCEK4NCuHB/ZLjIEdZrGuEj5dBiits
vHL/CscBDdE8m4Bp21AjDNe4sjugdV1FhQxgMZh16ZWu95y5KjdompJRW1KbFbTUg9s3l4+DjFl4
6yFSJWHUGpfojXlYn2PaGF7dF2u+y0pXrUX5AkSir5ptn54Qim0eh8oYkKMN4lQgewD9mg422Bc8
8/wdFGC6ipgniZAG5trqiiWnCZEcU16J2yFprnxRrOkEB3t4/3aClAWJyOHMKNE8AdfPv09VvY2S
HkfKYZdwzHv11hlA10TE7CeSRz3kFKjr1Pl5rras6/FctUtd8Z9P3KncryruSTUFZ0wnuV8tR7hF
GgpYP58CflRCv+AV71SZCAwQUWmdeGPWTkvIwXZtpuviZ9AxnHjohC+OhIZOm0ewIYizvCf+5tO9
/cNHunYGwkhLFDlCPSyKWwcNtYCveD/s2WtW+md4gIHt23Exex3UNa6IpMLtqzeuP8vhQsyY6duA
lV+7+eep6ONiRuzbkpesLvb7U9DqSGge7F8yWHIipoirJd4wfPyWiWBN3CM2H4yRmFzl0BbRoTiK
Wn7sY0NV5CkZ1CGVGBWJ2Ongp37laiTvdGVqlu6MlJeo9YnAa9bYIrkgY9NbZ5q1K5nfvsO97mzs
5NsHylZGzbQ0spJ2R14wSt2S5qJTgau8Lk9bN7BAlJ/WPuSqB9+tLDiOGFUmLtSxyQBjMLUixNYP
0Ylas2j5/fLalCc+1D09ngkoMHf9ytoJlYedk+kPUuOW8d1GZ+h+1mDp7YcsqFIQgkRaz8uVYaPn
w9t6D+XojmSL8Kz49i0IEIT2I5Awr+jXjIvSo6BdKkvmHXj1acklZbjH0O+iI8rboFIIKQJcD+LE
M3nZR3Tcr204XyoIZ4GIdKpyP4pf0q1xhj/TN2YY0Me6G/mLx1tehNXF851oKPvGM33eCwCGXQMI
69XaVfTOgwFyUGkV+Pry6+SP6nmgvmCCeN4kMsWXwGZWS4kSiZQXio3bKrgPi05SrSh3BrUxH5w+
BLpHTruGEsKwwOYFw+iwJWGauy8F/X79q+NrY78D51UZ0pxCi8QZi0OQdnab0A3U+3/EREFZCxJG
yPnJmFdkPsKgR1K7AxoWeRuY9pamvcnxc9j568nh3cfOxuU/nbVi++YjrUQAALFDG8c7LPLAPRfU
ygL60KPsdZVRjHWwkm7foYkMba03wBOPO4a5EzHlHrFMnBT8Cv0Y33in4P1lceSt8B2ql78wK2xr
jR7kQHxvD+VBCV+8u5JSoMgNTWDENClCJFGTJ+bmNi9aKtzAbaslW2xLS6DG9eQ85IsNvtKZ+QFY
i/NWc3ro2KjNpLmHS3h1in95omc2yGIHYyLZV1qAweUyUNkQrznlQXLPA4HwC0iBQOk/h7wD7/2C
NU8X/LIWwaCtQmtGKA4YyBLqK6CYTrMEfgvdQeTZjtgb+hb31FmePYTkoaOYVZF/lz/ck0icr1Tj
Ws7c7Szy4tR7L+Vw7zEFYgGY6TXoxqciectKcsprAOBpUtaCLTE75Z/uMJhO3vFAP3WUhnh5XDP5
yysDOGvQUrRxWyH0nmn+FjA8w9yBmojAXOMD7s/X4FysyE65i+6zwc6nbHb2T4nH8wkAd9M/L0JS
JI+r2ZoGoWilgwgM1NOVEnNu6avVWj6KVCCR81O2JLN1uqMQA88U7iyUwUjGfW0Cm9J24+tkGqun
mPSfZkf+xhkcQ+JlfS4uL/YUXlbSXtjFRmpfj+cZ15Ok5PfsW6N9tseiq0oRyc4tkFqaWi2z94JL
ZXzHYeITBqZGqfhg2ZI5SzX6cmB1bYuJpF35IOFR+kLLsjGYVwtLIQDcbICFptQF6WVJ4XhaVp5z
sgX+T8Kx2ZoEqMN74TVL2TkfzFH5vbsP7Mwi1zrEyOjh+TWkJcQs4Eu/UTef5Efs54FfcCfR4NMg
+MNxb4s467J0Cz5opPGDKi1K8WFI67Ds9yrlM72dm73sA+ITtC30Dlh+9qdma0ywzgmk+uf8J0YP
aaGwqs9Tsx/3Fz8z9Guzr5zqoY/r59zxeBR5tZ2kWyddqTNe5jNQ30RStU7k8u9nElnrdjSjMoPs
OFO9/9zxWIvxHqHhbzuwThlqqVpAZuUyo8GtxH7ClWYtzqyF4edDyILMJU91ll32Z+6jj97mDrEJ
9t4K8RtO6Ln2X8ie9qY5QN/hPe2eixp3o+IwE/Ls3NofrUI2IUvEAAsR/Sx5fGAMbARNIdzN50oa
N3UPdnOLOHm8MEFhhldeSPf/xR64yBY5M6fRRxlHJG81exxULoIccpgwg9o5l5JD0FLoeZ51FoBj
7WkxxTNIGto9HgBP5A3vbQgE3/CLfBg+d0R6rLwqf18LeinNBB93Or5mo64s2yfAiI8MfmGRyQ3l
jtNQZH5l1F7Q/z95bNNI1cGR91O61SPLyP5ib7PET8KBucl22dA/mk81J5RJvkL/+s8FbNT/uWaF
jEnBMMMX5F9fkeI1zw0O9CxVvbJzZH6LEgsrRgCZYGuY/+o7asd6lxtYYYnzSzSVpaOE+oP3OV3d
xvW4f0GTMh1Y82LcOde7xBtL+soU/FQVTiJiTtyYOvkKH/A0PlWgOAQOkgyYnJvCZDg1eMEZ6ukm
4BPwS4jNS2C7vvRmrG6k+WssCnO6SRrUfPO3l8B1fz0rp1emcJlsIiWDgKz0bpAao/Ep3CbJCKPS
aROcAZX5CdyVwrdNFO/uC1bodEDOg/n4WW2AbZlVmPVmgbdnEY1abxH/AoezjhEuxuADd8wEfTbu
s0K4Dzt3cJw9wTjKwglocFW8vLkyXdSOq51rlqfrtQ3LjJw502vHndmtfzDlc1L50KUaLtIeZ2YB
kDLLTs1dnYOMLkv1V/orkCMp+yVcCPxrGCBq/jcrSGViGv1iorbiyxfitX3W2tZoB92IZjhgRqUZ
M/708Dkq7AVVtS236FhUJn3KW7cxvXA2j3G5I9cW72+XfWmSsQ/bwuf//HuaHzAioSnKtWGCDVt8
KUbqDPVm0IPmSJUOV7dbaX7HSBlfA+XiVIQROSFAlNRz8VGr2WKZWFhxabKEw8MHqrC9Iv1qgZ+x
56lAXVc1vAnHOsfWfd2oB03HXabwFW8nVPomQ5xClmPTrskCVXoXZfxg3SmRnItGW4nkZ4ssJtRQ
9o5DJioNvy+hFdJVIqVxX5iAuNwjsxEhNSICb90AHBXmsoYorJwQlf5O4ZqFxFTuABl4MK5hLnKy
toE8tquGYgtBuAIBIQ9jFSPuh8KHz553He0KIIjavkYAmaMAs2sAAtI3Dq2CgVkcbEhA12mEBiP1
lifrcPMTa2DB4B8ZRy41NoloBKLVGQp+20o66h5qx5FIsnett8u72nCQK0NcTlMMGIiWPKu9+oJ4
8CWhGHGjHJ7ECqDikQrf6Er5UUl1BDezVEFDuxu22JicIfDF+dPkIE1EWJYn8ZR5NPSvzn/Oslpo
OJGgOTOcFFdCruNnV352bg0Xvuk4P1RK0kvwuY5zWWAMbbqgQSpZzJGvDERICz5tAxAFOBwWLKpV
vW5JC/Wk/HgRll20mxTuF3YWPm2Cdsm1bKw19r0xIff7OWBMC+Sgm0emKvPabZC+frI2mf6T1+nd
RLxojw+WJfpa44jX4g4H+BOfEcq0ywTZ34rFv/igVNZNPbCivuu1P347n5P3u/8MMywq/k8N4VRH
dWBk4KLzCxNU3qU7zU/oWMgHvH/ANNM/TGnAakXtXsFp0OGkgOQQ4a+H9kYdMZFZ6eyvDqKeyumg
P7+L+vcpetxy3w9zTYNOyTEGaomQtCeCuh8+p9WpQqJSlFFAb+u3av6in1TSlYven6XiVNzlxyfC
8b7pgWJ1DhqMYVKSQSB42+O3y/nPy5b0sg9mJBFCRpTYhjyrB7trjaB+wWid0//8s0y1Moj3SZyl
lDDwv6DIHRc77qagrXkjL/kVEP0QXdnSuStrFh8WjbR1VbhyvqM3BW7Of/r455YTC4byGWgjD+MV
WrWT+owpJhsgu2kOtUlDh9nPZJJ9+2bX9ri9yTYWr3+45ZomJoJULjbRVmWkCcSgRMNR43wrwwbH
z6kShzSPXMkunogU077qnNPlVTcQh3zyQKnaC4oo0w+Z9Vw0wh+TEZMgDGTYblOhLnv7ClW8EOA3
DFdsymDL529Ts9V4GTxRSsF/68wqUu4k3++QBrMfaqv4IiRQ3DdqejveQSEEiQ5hx2jGyJpJnECl
lbKFZ20UHblfdgVI1ZAsTU4CpKZWRlO4Y/iCHOHK+7OVoCvy2fgjRKephoNHRLRy4DyN0G0fPcns
Pv8LHYOO694d8X7K7mWUnGg+CJWJ846mWvVSIuvVz4eg/M+MTMlexDUvZFIALRfLl35HLd2ODjAd
CJhyLGq1V3WiBbXALpyjrVkaccZe7eS2ahOxHaLfb4TpijuXxUvR72FiQVxbdhM1GnGcswcbScyV
bV22ATlgyJgDvGbTlZGtlsi37SLBlw5MR5hPPYgkQMaow2BU6bY+j6sORy1pPZlZfEgB1UR+CWH+
GtT2VyeOAxbq6JiGGrGhc4ILj7i47OqYMP/0zDnGSAWTleNBGqsJv9QLrkIIua30t59oxoDa1363
h8Tzkz/0Nt+0uXjgQGkA4ocTBeZ7sTAuofU1up9qval67e/+Ok+KmxTxqCFuTO+uLx4aWdqBRowN
63X0QdLs806Y5mA45lXot9mKfe1n3L6dPy1ipIEOV9xRoE07/C5WWNFIKeCnJdTAiBDwZndH+H7O
CoB7VuG5OaXP+I2Um645JcU5QN+aFwn+J59r0TQeXim4p3O76x79sm7HuJn+KtOOcA1ZoZfNHHgg
rBhsd+sGxcDFYsVnAJnVrk7+RirQSbRFsQ9GoNg2JuqyC8pbrzXf07Ut4oXwBmlyCgSMbZaayr/B
N/XsRx6vS/gpUo6pUg5t2pWMtZDc7eqgzLBkHleeGKG8KvG+qBbZSqyBzf8DeYdJPo0oXmj31lFl
0jb+SrdIcmLBcnH3NFyiEJj0YjKTP5Wdijyl5f/EPLlvwYyAFUBN03tDgOwVOuARED0cuxgbAdyi
ygzzbKoLrt+I0tVQliykWVDoTpwOCca8qAcRs9voY5RGEgAFfo2F1U7duY4pGWFMM7W4M0MdSTGI
D0nGkxQ92I8O8cU77EN/FSYvLUTmcXhZ5iuPO+pIBCqn6LQM1re6CFuilz9QhgHF4gLfd4YQRl/O
/xipfesVA3ZB3APp06ou6woyg6e/w62xFVb+CezyqFt3gkgepDGRI3zNZ235ItONzt9xoXy9qKzl
KixUOc7VP+XA1iuuk/SrUuGa0yaBAv3sc2hiyt8BDQna2N2aRXUGQcFddOulMi8AxE9Z6cUs1r48
YtTwLBMislNT5roMlNh/k2JzzTXcjjO2iN7zXdIIrCBZH/pvqN6Qiz6eFaMGZ5KFwbZ6o028Tqqn
KduX/Q4G5EH5ODDKSVG+RM1L/NQiGcPBdnVU103lvniM73qUFimDcG5YfSYkCD+urHjknnBVenhg
iowXB6Jr52zbYXA6HaEx+9XabzJFQH8h+g30KXwQI7ESyRkw6y95jJYqaYKiyXZd/qOCuhd6dO14
d3WTv5AmhSMwnU5cDYJ6G1o8SOQ7r25PhVK9pbUO4wD301Zba5jZ+ggs0In8wL1trv28oOkCEpiZ
hJAO4ttyrI707YSP0d0V/wCSIwWJn6So8bzwRy9eGnk/CfZJeDXffvRQUL+SYQ5ErwrOaxwJI/S5
tpZJWLCVEQqhEAOlhlQM8Z6B8pj2NuE6AL5W1FzcnJ++C8LP+pHxI6VevXr5WVMbSrWJHU442wkJ
NIArJa08n+PNr6YrqVhSP4cXZvwWg1BOCczLtZ1MI9hgBqVbuTbzlemhzz/P/vJoXPxtnwQ5hWQ7
7Wbld/QPK9kukaVZQnU+2Z4FF/JqQbtYzJsGLgBBz+PJn9G/P69kHOxDFSIcGBZFYdWVi7i17vmg
iYLF5Md7ZPocaBw78kDBXxYBz320oUKi+Bj5UbIYGXGsqsl3irIa7ktz2biaSjrVIG8VEJAb5ZOZ
DMe5ZTfl4JWuisiRSHJ5jFi/iRc4bYZD0OUpf3GXWkYEv0uf/OgSVtyB/SDuYmu4T8Q1Bj88YXoR
JbR3srH2bW2JxNvPWhMxR86PERf7FDmOydN8siUVJ/1uUXwy3PHa5nQFahqSAN5R83tq9BRMN9BD
4x27sS3vh7QqNuFf3V5eCvW3/IgSCQUpqcr7KQgj/+nUPM6W1SuYQ3rF3a7qvM2wquzDBopSA79K
gU2xxCmiWqlw1GRYjEnhfCjUryOOSqOf5NPBsb09+c4arYwoRbqpburSIdQ/TbuPFJUFBUGixh4x
+5hT4z/aPpZwnaTXbNhcXEEnVpHihAV+dMLTabbo68VCxaR6KuK6ElW3CLiXek4vYMhtm9zKQ1rF
tUbwiSG2aQsXBQ923ll14lrn+gdSUr+a/rTIT37w+WhRRGKNNAV0YhA4djU0rFXxHmXzh4AZaYuk
gh4cn3aeNRo/x/sVrh4KIOMs4/cRQTarRzY5zyHoxVdxhOEaHFw+x5PU2kZYcYjr5vJn0MSj3LE+
QANIK+fQv3eyBUXjkQbANfwZMRYWoIJb9JOUh7o/PObUAAMECTaaigFzX+ruFv6GYv3BVqC2Dp6G
CNagJf64klpbVmeGVPb+5TW3edPK1x4AHlT9PVYuuC67gvuJ/F+qDzF4fyHqNLTTKbssdHXI0VVW
tWnccZpOOpnJP/xN8MmCY7ZHnanMrhXQ73r0b5xPoxW24JMERxIJGq7OFGw+e4oAtEj9YiwJXUny
b73q2L0r2n4IWT9mVq1IfyJ+T0Snd1Rn54qr4xuBz2/oAUOZ0bVDFUznbyvhGqiBqBjCQ5/R8do4
g0MFqaLHOagcD6BK+uqgIkew3TvGL8PAIfnE8FocwuZ/k4i5s7Q7pusC1HpCeO4AZO6KOGpfE/kW
aQLj6za+VsTA7QzZNR5OzE99bYxTsM0LAwARHVPp83h+s/tqqEkiTPUF4SKf5N7wpwxUm/Hwb8Wy
F3f+sHml1+ijFRbSK6tALPBAlPuho9tQlnGRuH2FFTTNfIblsmnq6ooNmpBYY3PlUhDILtxADuwI
SNqqXFsVHEgVhY9vgCsT6qZD5pfZtPMMfTdcfe2/kyZH4XBB3527LG+MhjfQH2ec557bh6YaVMTV
+1fBFBBdrcjvZxAgbptxETp8NAv0X8S3iYN5Uu6yLsZarDAl/RxQP99QjzU7JOXo4mp/qXohT1Kz
f90JSofox//lljnN/+jKi/EIO4n9B1Udb0PwUXTu8y+zURx7/9r3twObLp6dv2Oluh3kEfXSVVCU
CDj2b5ONRWZXcjWYr0QhosH6uI5QbWolcc4AYLu4S/9DfRFcMCJLsNPtw5aWA6Am8+E/GZgFF1Sk
SySVRYnpShQadb+4PCCJTib/q0lHvrnlNKlKQ5nDYZ3nPAUKsWUA0J6fGufNYQXmR+/Z/+Pd5+ub
YvxOB0WyqisSBvD9I1m2KJ3wAHDflMdZf7D6L3bIt6MGOqGkgrS5h4y/3esVk1Of+Xxtjd6/V+1m
dxTjM2zFrGsjVXcanjiYlInF0JjNL0h4up1ph6QLv2hqukpDJkP5z+6yFpJJ2OjZlspLvmUGNkNI
Oc8jFiatxgfoSveRPOOyfyjhip6HvNSWe8xwyKlNytGoCgqR4e927H1/Vd/DsQ/fv2qrGSkexoPB
jRYLW9ivnJF+inCHjHtkiXZ2ypbOWoPF+jJiV5OjiC+0lfwgfdj6RklP6/XbCOa5RZ6Tb6nsNo7w
Q01BSJZuNF2zWQQ6URVQHXQR8enIBRqpLALKaK4Ybb0UXPti/u8INsnQvG2Za2e9CGgB95IPzpmk
1j5pdtQscbD+cOr5abIpzoOf/W/DLVw/PqKejseJgAxFIc+1C8hKinqKN8A0cTolPgCT8vZoGKF7
kvUtwKcnygsFNC+yiRAc3CODB6SDxBWVtwOj4/S3vBTQuKifl/KpiAx9+10Pl2TLsRKsX7Y4n5qM
43/SEg3PKqnT/cwSamG4ey0TRkQECuMSOtfmIJDd7k/glG1e7lWUl7rAnRA6xn7Ql3bNf+WINYaf
IwKpU1khteXh3YZ0mSig6Bc0HldD9vRzRyFNIrtKglfv9CdR3Z4JuD8vmEq1t9nPhwjwsD4+4d0A
GXVnH8jyOsxEpOJYgbnuAW/Uy4BmCq4ynHjTBIF/giERlYn7h9SWJMPIvCId3z6Gog5cHHOLVfjq
s634xmq0MGUJm1ykbKwEkeJp0rtzBhaHRL8CHVmFmZo8FDULQ9s8GiuuPz16bLEOhGvwlsNIBQlJ
Tx17fUNlgXmwyZSZuyTLPTqdQd8+Q18ml2Br7nQtVuDuxV2fOZyk38tipS6svKtjzWQLIhSAAYhx
mYxGLizjkIeJPW1iroiSB8v3AcBLLyBk05tmOXKkQJR45OY3s/jHM4s1U3GMs/udey1l6cQSFWR4
tA7EnRAH03ymWTfnxXwM5ibZKRCQ8RP248DMDQVlMBuDlt5oK73820p8RpiYYWi8sMiDAWQJw89Z
5Q5iX1poC460Jflz6QKMvYG7dxpTvZ1OniC8qsvoDwXBHCPMrLBRSGKwNX78jb8gcJnLQ5p6Cq72
4e+gSzvLri3O4PmDBTPKwI5iaXVdRfruvkN+VH8HxaGoqjtWj76URjfcTlcnQLJRhat4mJJdNHHJ
Om4W8rxsyf5hpW4hqyBHstzQFT2gSahF6XAoPPVw30Wi+LrFhIA4dCKkrCFJPbx967rnmb9Z4O0p
e20RZwRJ79pWDIwTFeMEbqFiUtilXtNxQ9wGMApMKpA9Q0UciGgERqYbG3z9J/SwTUDZkeogYeeT
J//gx/sfpeT2FRsfKogTSdirCwhFjkhtjPRMnKgegbiLIydnsbXGcDdYCg3u6E/Hw8DLDExuGhd+
AZyEydAH6AVkHMtnhTXfGhSmccmC68nHN7xlCwAnWb/vbTQ25fkhxQDeCoabkTpY/eRatCoU1RWU
Fy3c+uKeOA86IbFMJpQ9gHTnv0ByyBr+f7zCOKnOADUp4Ofchg20XncfJmmdJrH99RGTdyv1mxSy
f4z9xr9ch5IR8ByXxaqLu1FROzHlOsDiEkFBulNIh+TZQwMMMungn43GVl+pYZW3I9CaanRZGW1L
rTnAZx44qvTkRCPSVeRfhvRuZpxvn31kPupTxNDxyPma+3VO3mlOdO5tZ9NoKYYx9BigpZ8qJ7SO
MUtDv+mUcjYhrw/saP4KNpfFkIB0eIZaj06zy7XgaGQvGJoHjjZ2vCKRfwDrFbd6BPL63Us6lX3w
S3fh5lg4wNavOi4cEy4pbfxZi4ll1PNAwC6qbyP9vKtILRPhrqwP58BkDXPC76y4eL910m+TAvRN
oFRFyBuPped1EFhhEY8IMXED3f3wXEJMmnazQIoWbEWtQ3pgkhPrRrnevrTC3hQ1XbAFleu8ZZQM
Ggy0OZG0wqUi1YguR7OJ7tsdVHcxJEdSR6HH5HO/lCedhuqMRiz7JQvq6/x4FiQBzP7t4c5wz0sy
qR/8CNpb+hJogq8r0IysQLL1Hp3PYp7F6Vm9mY8QNSQclLMVeAxpZ3BMG21My02mFNfmh4kLxxE5
OKXRL9kKsAa2U8JVlP3CNMrHBeaQeuvUEjYO/8fe522xLpmhXbpN4pSYniUZmjgjXoFnz6VbZQUG
pRN3N+HnTjs/SpLexd6IYV6jxW3QRI3wQClA13kw7adGBk2dSOckb+/eNRc4E8VyhMP5oKBDbrs/
RDJ2/YQxwgtBC9xw9l9D2qdT2I72LULilV3IZFWYUD6971q0Beukv+b4phvVx61PkS9cV5o4BHUx
NuaSOD1YYsW+FBmyxOA894zS7xOzRz1Tk7ZsWfmuJAfRv/46KYieTyOyLFXkawcpKJk1fBS93vXo
VJP3rk7GPVgvRQBZrnAzLAmqUo75PDed7o3EYlKdk3k0TyUOQORb3yAeiwyFXALmYB83ZptapnSA
k6Ah7//w9FX8ILwFGQelXNVQ1gWXTd7cJQwmcggvRrCIUrwxmcDpvrYfH4hLiSmvxPpt5DREuF0S
ChBA94TU2Cc7olYsemkpGKhbF6lcXDZHOP8UMmMwQHYk/pqY6sm2DsB1dPDDFJVrlSxmQVTVXj5X
K7wxOtHyFoP2bhx9aM52xSWi36OIN767A7bEoJrz1EDpnhId3YY4tcsIQU2nJzYupAJOD9XlZs5R
a6on4TohogNp+JZI7BHbXYkwSH/tzzS1iF4QmIhfBPDJhNTENDEaf/HVKBBjBRUhYzJ6r4nuvrNi
eD/CxC9/NTE0bs8HPS9IS6DUBXxJ6y/mvi9w68RzodnfflHlYdG1astcDBBUXm0pdrh1SLjlYR/s
uSGdEO5tp/kJKa1FFLOoKab1xtLs0r1fqjJxGCt4AeCJtn8lUZ/ruCifR0Hu7xyOJ4y6IJHwEyhy
0RksEIAu1XG5fG7Zw9Y8trN4tdw+JESfTIzschORZpbK41ttJqw72tr3DiiDJr1yr7NH+X25sY4u
uAQqnuj1eg5vNhZk0/X+mxpni9aLiJfba8MiJL6OtwVQrW6Tv1jESaXXiZIX2FxLBny5JRI+AUAo
90OEjorFdqR4L8R2ZdV9d8WnPBA53b23IFHHE4p8acAQCC6k5PZ+mmUEEdX2W1FWJZrPxtkUMqPz
miNPa07M7EoNYk48TqTmh4f/jNbIOoMIkFm7JAtDubaEhFn3KgpMMHRWO0egom3yDbWgGcB6FM6r
3VB28lqS+3+l2IIQktv1c7jR+DuVtc0UMsvtfhN0dPkT9VJKgbrOXUSiVTmR9TncCTsSNfwa4QWB
yEkycdbczki9zZ80v0Z/9TfpiNc8WSPe25PoKb+LHE3Fv9M+wOUM2UTF3axwbxkx4KTWwH6G3OYM
TWnQau7pxZioGV7nOEe+o8XTlsxEYY3kmFQIK5oPG3Zl+kXhYbHsJYpAfYAw8sZaNnJt1hTdeB2h
+NaO8O8+zTsSm7dOYC/eXBzC48SlgGRU15OvVZgjou7GDjw2c6XvE2/CyPlHnZUsb+eSTkJHVts7
qLfXA7ihzDCyap6CymlCr/cFNSp1pdbaZ2p/pYw5eFVdn88hUHSeAV/T0g4XUhLAYUrTV34IiBml
uXCYDXnRE4oKBbBdAsKaUULcTQH0TJV+xOZCaZ6AtihWM14ODRJZzOv6rjaw/pX3SHceujf8kMAe
5EgnK1UkCKSP1rVkOh9jR3oKWP5QU0WuLEhW0YupZf/156jSbh38LGqqbZDPoOMLDwWIyxNoPT81
m/e/gw+GSofFe3rteejQpZ0BQUBmmLjgcaPEPT2cK/iLWOO7xXXrjB0VbO+Uu/4rGsM7Np1txGL2
h3mTnWyn4SFj87mhowflXJN7ucYeFFj2WJp8KcKSupxfGIvHjNmelZVg9rmhj2APavVgrwNKssIV
nXp9BHrr1/gNFYXATn73IK1jFPwYXh8iaBPFyUqUDlI/RSiDX/jVUjVBd8PIlRA55ymQf8jLGeEP
zL+gkgZZLsaChAaZ/HzcptnIhIoPp/0mzoFtbAMv4g5x33Al2FK4efdEfrdzjJf+WB02JKQmAury
H6SrKh2cN6U8fdljhEsWNG/CJdi30bstYHR/xTuOERImHD+s059uWet5HYANKHDP58QaduAYQ8DZ
ss0Y26RqQHOH49P4rcOs+hjkEV4Ezq6Fzq3iCuXaAiq6BfXkg7X3JGysSIPrCHh8bbE3KHlKMPyo
xKiaagqTB3WSvzFQwXvH95Vh7t3MGGhrh4dzNm7Y0P0N3hu4dFio/UhV5nYcWnaYuolEFLmFHhpq
Ltzdx2aQxxfROE5lUsHRz/iF7gSi8L/I4M8Tx2W9hmu2pGuGLD+4ewcMUaZKc8rA7u/mCVlX7Fh1
j8eQUzlGFs4w/4l3sMh9BNIgMFBMehTLoR/OYscppLL/JwqZL4yPCd9iRxCmG+hNHALpRzQUpm0j
yTDXKhGhrsX8ReSFX0EwsU8VEZq98LnmD2CzS3+uzSW3oer+d8IUqTv/UqpusvXydpmAkgd2/tq4
j2tf7gk1J3P+2jwC9Pnp2m0ntkReybru2HTK3i94Qe8+Avr247y2H6QjEPvfav9T0sKTZi+in2az
MIkNobtyoA9kbd1TFTcOHkQQTDTpmU+f9Qq9bsiGft7+gj82rBGe1jSYbzneYyD7N5sqkCS26oNv
wgnyd1mrMMrkwmzou+OmPLzQqS50DwCqtEu9n7Kx9xiGxPjqCLcXlaQUCwdOqUhapXX+UJoJLaAO
PSL/dj4vAwaM29Np+aZrCXQfAC47TU40pely5IdHce5PxsQhDtzVPqIHsJSPXiGW311T0T13VFR2
Bq9s3MynfqL7D5AQjm7mg5VI4f0VPHd/WvK0/DvFM0gZj6Y8jE+GOn4e7yN8NyM18KNo56uReAgg
1qdeJvYsJDNNNWeP16RcwnO7dkoqJIci0tpeHsSkRpO/HbfS0BV9tig9P+RnB4LkMd52wjlDOBBC
UTsEku6O4hvNpYQUyFRefrldNwWqOZlS/nbKYAY4hQWXU2nJDaOg7F/ABmdR7fWq1XgIDBxWFI2m
LvDQEgorClLzFnk25qDA3e6eSvxvycxhwzZXDoQU/zBcAwkJZpdlhVbOGOJmp7fZl2PTw/Ccrj4s
z1jrqARegiBlbamAv6XInJD3BX4jkuOBNEH4AcRRXGlF6/iRIqRJwrm8D6d26kI1GoKVMdMBKaX3
TrhwbJJ8E1z1Zcy7qOFiSq3PnwwZd6DSn9t86VFFLfq46rtFQyet5w7qCrJWAm8qn19lHsmf6W8w
2A05lyPX78oBPfPBDZ9jlNWqaJoUt+KY9U/6fjlV/q8n5DGT4EHQlIB75PHNToZkBReFGdA+D46L
JyeBLHtys/lhIpfZI8vfHMSfrr5McCQ3pdN6UM5Q6wU9gC3ATsZHX6+HheJaFeIg2w7qHR5Yk5nQ
QftSpw1YLCHDRYi7JPp/TFCwEasxPxvciTZNyzTeWdWY7tq9I8Ro+CHlvey2dDtGWuoYStXFV0My
dgPON2KA9AaobQLv0UrjzbbK0GUhBkjcJHY8mex1p25mwhXdvclFnR47e2hJ8B50bRmiWf4Ze+Jg
YMvL84faNKRa5TSQszLlljcIueRH31xCAklpwXTCoQfs0MnspK5FHZxqwyM8iyN/9n0uKWaczM6m
1t4OVSYyIfpJVFJS1BOEAnGXWxTrWABoe52lDrQdgwGjKe0ORLh0ss/dI9OkaDHfjZlCELfxFVKj
1pco87X97FLfvUSJ4/4yzkfB5bLshTS22txfKkDMFbzQZalfU2wQMRQIrpVkDv+vwEW8HRovnShA
30REVFjImReXaOSjt75nwgSl7oR2S6NeJ+/KtBfHi9TKN+x1mvJkppVeUsZz4+vzXHrjdSl0nBGO
wSFzV7/QfLneB+U5wfmDGBYJamtAulAjtEF5H/QD/tFsIVESa6q/5M+piF8/xrDFs5ybVJLyZq1I
m35bdEB/RUqHjjItcEo73r/F1j2Zu2/Z2/jYBmUSWp1M5jJ8KLX6V7cmH2nqHUObiC16J6E4d0l+
is0Fc8ysYlK8RHLkpcGejFg1OW3ecPEnCSsRZGjAvuwm2BVoZJLsuhKNBBH9sbvIFSIdEL0mdxAl
+hL8TZeYT9xOCuJlbGRkXasTBKArZUF4ZgOWMtfmtT+MRIU5dyuHpazOls2EtTIPDyBMUOYZSvo5
VipXyT6It7sCX4xtIwzmcAcxtCkkgwh4HoXEcYv2z6IlpNRbC/rvtgBuhjloLKk/novkKkTcJ8Sh
/PB//cDQvwqTz9+xpepUfgr/RcjRz6El425xb/8GWYlGUK8/YxHqzZqxCiMWpNAoA7Tu3nkBK1Zp
1vO7ST8zoYrZa0WGVxA1/V6LTPiRA9obAp4jC+vX8aqdHVk3vpoF70IFYLQ7IB9L0DdCJTVZbcUm
/3JuX0KeMTgbOrDWr7+2DyYb/bawxIxpAjrNkNCoURcdx+H5MtaEAkpttiGZHGgli1dbROArC5ha
1hgTjk/tJx6r4Mcv8KVXP/5NN48Qv4bFSNG6MQOqA0dsI98mGyqbaKZrMBeurBhW+LpkEoKfHRGk
ZklOYIXMMKoTHusDi/aE8RzxLQdvZ4JilHwORTyU61n+n4+PlRIqEhlXYRPV5/I+s68wsanw9Rfn
ddoGXH3ir4z6GG6hBtnDGQkZXrPzoMnpwGiFuBXY0MEo49bvm8+KNryG4TY4Qr03dhmOf62UnG5Z
59j8puO9S7db2XfsVxwvL2BXQf6QJYxBnvHqxW2vE9SonUOzS/nfppSYG/4xB3j0zW5Ua4y77SGs
3n25Koaylm/bf9MrK1rkiX8d4pGVFQo6KSWwVr91zL0S2XizAr9m1VYiK1xn3f/Nev06HaSsRpou
0hXSdxyVpQs7fgkxOOXKoCA82spn9iZ4+wweS6sag2ipa73EYFtghEoJO9dXn3+K4AcWil3F0YNh
iTUzBofIyA2+N29JXfVGIwBZGY5Znd/6FnIrGbImOm0suqBWi0u0JfRHqaOaMGwlQiBBcUBOMFYF
8CDUENAzw2veGECws6M9EkYLdtb70KoP2QZxpNelKl8O4Zd5qkVXr9CePyPJhazEtR1z9mSKLABb
7iRjFRTBdY7wd3q0cVTNBJTmdPIcjD20BRwFdV4OFeN5hmfhvPytMdRrsvmWg4PqRa5TsuLgLciW
1DMJHD3pVm4EhEZdnNJuHikL/VDaXQb7xo1F2mLT9+j+jNHaGhlMAd5qO5poz5XskFfk6rq8UDiT
ao5gzOAXBqietFthcXEeEUDqiFIjYukF8U/wMVOoyZ2R8F4D3RpkDqIWheYdmDFWZEgGDDeM/z1V
dfCWbv/tIkYJzP6594vH9JtnScKm4ZEnVqvff4Kh47e4AZxSl7/hwPnqh8Z7RTpSj5kDVLTlyiRt
UrcVHvYP8kV85V6Z5FDCGnDnd9H8w11GWJTjOHR1xGS4Vn4UnjrSj8pQJfOGNd7iN5bQLACKunsK
+YjNTJ1pGl7SIt6j1cqj+2hgpW7wrMmry1dmBAp3VpXNZlM9c70be6eqkzC1mSWuZR37dQnIK34m
gJE7Cdyh351tAEvwPeM2Q3zQYVQT0f2BCfC6i8mM6dL/6DDv/e4pWY4EJlzu9vyLlpHOV0M7y8MI
aaVQU0s2A2KtMjNMsoLsjPGoBnq3410cRypeg2pGBaOwXAWDFygCerPVCaYHbZzGaVz2iX3WOzPB
T8q5zpXtI4y42R4zno4JKswDpqkGXpswgU3pe7sxrpsVzd5QFbIFS2niDaM4IDXXTNtKoiqzBj+G
nAA8rw/oTga66KnQBOvs3ju+LrYIiz8KlF30wwZjzfynEJ3CUw48k8sjMVhnQbcxOBBydrLiT2F2
nIKsYUThYfLNXZFNNkd/DlqoEIi2mbSG54fFzwBpIJzl/JTLXI1IETRCJjXkyv8XIlO4LWZzrgvu
UviTswTD+/aIFZrakcG3hvnGfMliVbTRtaYWNhDbfW/xr7nSTwaquSzFbFr5PkOpqTlXvTBKrXHo
D0oB+j0lGhwcuWVYs35WEXW1n0UmbX2nprrW1hJUTTS1y1qJQ6xbP7DwQZdR8xAHgG5HAPYlnczu
PYsdjFkwKScMvtxvcWZ9OreuyZq63ZwOrtiRKw3uI5c42DBY/1T++DzrtR2D1y2memHMaqP2p1jX
D/1rHOeTIrO+ty0lukTYMQBran2YagKofLOOCKYCEJeABS4IUoJtTDARqmF67GbgymPBLmWDzUkz
DZWKUORJtsA0qqQ8r0rPGAvWPb+SuzRoyvPu/F76tc1NKH4l4J6ScqqFo9UCCjXu3heA1Kfgx0Ww
dHrNe8biwG6dPA41LzVLcedcX9a8rF0+b4ECrJ0CAt11gjAj3isvFKw4uzAbKFLT+5b6NIctjkl3
0xDpGjZdEfo21i1ily0ecLd0XaR2xRQSeKVRkWgSxub8rwaWvN0ivGCm31mfphvc6E5L0Y6DaLXz
riqlU8woGsKdU1LwquVNahhz7yqk2vBEvtjkgbi0cQblZgpdwRWdqffsy8lQ4PSTnIQzpvFVIuM6
BP3L2A9ZaCOGIfriuSs6/BmDZS/UqkhBylKkajXXUO2XvkhjM2au+O2zReGJbtey22Xsw9Xn4+G6
/YgPDhQ12vHNcK8zzR/lFba1WBLvETfZyKu42rRLUSC7NXwazN8jSxy0pZmxRUG6Bpwq8Hk6HPvM
D72drwuv8xfJ19OPD41bgMHtvFAgrl2Dl5AgYvwLpHRY5Ej+N7aqkGEudvxO1obwwMU4S8lpRtS/
qcnJ/isa7W/hS83VvTSWzdtskXLat/CdOt+TeGxB41hFOur2S7a3GNdXukUguWUbFhRKZYZ8Tero
q28MYvFE6jow9mVGxwVq5JmgDDwKHZoZ749G8ICq1g4fYl2XWgRRl7hc7H7y/c8HdeD3pqidYEis
oe+uPjrIRnup5uND5GiD4tCELDSiZZ6XXj8mfpvspER2m4y7/penhvdxYRkjkZeRm2pDSs/ei/7s
v7u29QrDUXVTjwt4dOWlEBp7U0G/s7RKJ2F/48gk09sLUWuS2RmoAPzS0tevIlNHD6Pwogt14OeR
EyMnAO8SIZcUW+rdIfyP5moGig7JPtJywGDkCnPwbXWpdohrdCigsXP9NFrjlWSw8qYwQdiuLrQg
PzCCIyRMBKauhobm4iBi+HQKVigROqlICzjXJgwj1d1Wg3Y6BLpUfgQl4P6xkuM6gAIrbsqWfcf4
tDn8MXv/uUjXyqmlCmXM6m55MyhS85q96bOQh2oezQr67MTVSueH1qZpoZWS4+M1uImkHjlXOrN9
Ljj0qQNOHuhviXZodtZ032FPcO+Jm504wYaJ0hqfHLIRRcLYCGw5ZmbzF8u8h1qToG2cJuG0FasH
H0vTi+5kkAlekMzC09qNcyeLuJnfoAbKEofYWIfZ5r2d3VpuYNLvhsFZ0mi1qevH8kkbz40pIt7Z
SYI9ICX/Hum6IeunI3Mvp+Vxa4/6TNWV6+XQolO4bQrKyTbA5+ZjsLJNLCpSrRoeGC0VfsGSQmDI
8awWdh6r02dGPCrXRcJurMbwVZEcQKqMnzYFN12S9A8R713EY7HI25vWqAHGIMlUN/opL7MOq9Hq
nKrydptpOrtU1m5Mgc0G+8Hz6B4EHAkmqc13xlJybBPphjLWk/Ye3w+YncvaYiYY3qNyokGM1BwK
H5MyDXOo2f9b7BHJO486Q5wNGa0JkfESY8hoS5WGBdAAMliC9El/NR/CvOr5Dcyqvrux/pFvKdo8
pVaDbWWmzFp0cDn/U/7akErGuyZSBUP0Y5VfYyLtnIFW65+y6NCl+MSFfM3cfPg0uDmOz7W4RkFH
eX5Z7xmr6ONWC/pZ13+xdop6ghErd/WxZ+gGQz2ndtRpaCMRm1Z+hsPa29k5Q/sGXejAmvrb/uCF
BGdsJ633t/LThhPqJ0Ti/V6RGgUYavVgYvdsnmpsFpWB8Z/U1evfeEOdOm5BBEeBQQ+Ib1pVju1h
+e5J+vQ+EYSjMHA4B0n8MF2mBGtBYlK9ddqBpBsWp9qfjNo3LGd0XQ7fJFwAkod9PVOO4E1Ww2ZJ
R6BvZyd2kgtT/JW0NLNGAkFbRd1da+K8oauMMdvEfPahN+QSjU0KvvaQPhiIbMktkPzk3SJdlck3
NtGHCFLIr40hRU8jBpaUH//thahjY/yGnR7vz65PTxTM2hFNN117Zlh6oZqycpKdeGKJqANCBaOq
3MMNqDOMLvWJ8HpXA5/5X1jggq3qjVHxrDy193uOGNviT0kXGFxmjCpRYvc8uyUkjiNV2xIF4zAA
hq/I0XTKU9cM5Wd8cqLULCA2Yw8AK/zAA81vA14HIsGHK/PeVQtJKGsvK4uSAcVjEz+HkPFJTnXh
VZ62h4UMP/Dxhie0Aq0/eoGPoeScPUdYFUVaNtYG7V26rkDz0BsvLLCkEk74C9tb+9PFQNRaCeCR
Z9k1re9WWl7V5qLQ5+UvzEwlJsyJk1/N8PNU4swYcT5MNh2qyNqHApln7pMFVsUrJ0c2paMu8aSu
mqlfqYdN6j3VqqfI0Yu+s53dHCdI2WK4X2gwvc05xNE9fOoVUcG4Wiljey2+n1HcqLCI+XOtqdBD
BEt114FKdF6j93Fq767UaPy4aMYppChPKbqmkbmdREdYM9n1iJKFL/gnLn+yHV1E8/4/5/C6hUrd
qxN24iuDfmSeUP+cPCCfHZ5GWsU1bAeLb5M8pmjYwtfgr0biXK+H++lBRPo1O2TJfxRqEbicufVc
0pi4HTHdzFfPi6VF8b91LdZK577ALmqNDccTVUx0m+EI2B5pjFllE3rjMtIs9buy5EnMaMAIOgrA
d6u0nz6vYd+FpGbpoVsgHUqUUzd5XB6JPSaZvH4FUJDQphyYQzRqLFQeMwKAXkmJ2Avw8RzX9j+q
G26e3Yu1vEHlqrh3oyvw7Kl1QnvWOe9RkmSzOudovNuVCGKnkBCEdzLkdmetqi+A5r53BOxhQPBN
8UsigUDdvb05Sq9hUMrMu6ns1qK/botdsL22bQh7tt0wyQ7wA5HJ108Sex6Ovd/Z9cnmhpCw+McK
Vhyd6e6OJMBimm2hYIfJ86ARFeEFVkapTb65GT4siYjPWraGN87dfl2fOFO3Rk0De18r4mXIngUp
SKbbd8bU5mMPjACa7rPtRCU7Wp6jyNaR37WGvfI0v+cRQoIhNeLdz5yFMZMa7E+LGv6IdVVE0/oB
ly4372HAH9QF6DrrNxZBsolmj6ouKfpaWIKuuxtmXGdVSi5AJAhIL723Fnwtdfo6MO4nKUL8XFkq
9FMLsewUvXeEZgMDjKrLcjrqiJzUS3t6bVGwjTbvegWqEtbZ3A+TxnZMJq+JC0V/gDAj/WyqLwoM
e3ZGBGDTAY7A1JXg+kKiwvDMg9Oj8RbtEBbOLm69qGKg2uOh5+mIb+ZlclKchydE9e8THoHRVnru
iUeegpw1CJ1u36PeMGE+RWnTzAZMp40D61IlYRUObZHt1AAOHIpUbZ+Cbk+HyDLusquY/x8GzDJH
AzwhJnzuUJQQFESnvIEHVF0mOkOritNj7RcNdb/iG/y6jjaKNs4bZlwU8nTLg+LMEqWdV6WDvM3K
BhY9Ls/qdYlc4RsevmimDnvyKajNfgHnhAbXYGR3GHGA4sGBkbt1wOvG/8JWMzAbzZjnCa8BErdo
sXFx5H+IaMGhQtfi/qND7b5SZusH3IOMZtagcWqM2yDz2+b0TYLqV/LGbxtDRuGm80U9X2xramOH
5xNNOu7NbzrPoZTZLOruafbEIFVulgAAm8vVlmiGLRn2Do6JkzcWSCpP2sGY2wMWaULyQ5aqC+8Y
Tvva93UIFh4dcc4zUEEcEUfzQdfrNEArM+MwvYElKUhzxPQJoUGoRbOFs/A/6i5mvmc9yrETLTi0
g18L2sHw1ftx2bwZLJYrx0jjVzipacEh4NO0cAdt6Lgupdgrx5QF3gLEARNxD/tKBndelh0nSGS4
Edy0Narg7mz/my21yO0Bcjlo/kfVXYMVh6+pqGXKSd2VOuzSruftaYmGRqUtRHsidxXUhEStTz8O
yyyo980nSdvFuYjcPkvEUY4cmD86+/qHF3HJfTsAwq9QdkSOJSFIaQjiOuotb2NEdIL4kERtsf5x
XV3tFZU0Ls7iXZ1MqYAQRNAnGz7JYSkX+XnnVNLVIR/tCRPN/7iJXJAt8oVVRYl+pI9yz4WSVRKI
D5NGOtSYTUf2OQs3xt7yIhA2Nc1Tfs4/4mEyChk4R6oNllorlR64i4tyhjWTIFqWXnZRCz7BEp2Q
msdXHLcu6aInWeGxzovmR7p2UoCDlt08pKDVKzdwS34euPxvP6TSkCWrCNgzu2plxy/ZRsa3U14M
TC1kbVMKkQrnjOTTxzG0WoSRyPYpaLInerYVZ/PuwccbWjXv6GIWYqC1+yghaDv6tjG7doSDqLpm
s6RKg5xFAseTljizzoIQqffBp//cwNj+P5svWfq5Fpm9cT1HXn4nWwW3KGZmxq3QQDufH2jAP6Bj
Ngm46oRo5QsFBXYEmFgKm9hntAYPqAPkhOq+IwVV0LtZ/v5OH0HBEAUuR9Lpxsgylh24gB6MGOnn
hrtcADmhFXI40ofwQbbbxn/FATFrdK8GVcTF9pZ0RSJMgrfEpeJzaRTiRSeIlZUQKJWclFg8+rwI
BO9udIUgWwZtHkgF3gtkDjcM/PZGsjwzWRhqWJZekMQPkfi52IPXRJiNM4Mdi/ob6FxN/Qrpx7Ht
xz4jWsZfmWOHbZgh9elHU4ubDnDRLngziht2ehSRU4QtpfDoGH1VcMtT5wJZBHDRiKPn3y116xMB
xvbWOo5t0vFrF0yglMovHpTIPtvfsPbEeUYlobHhBHciqN/+zNyW8WF49hjwfnad2ErIEkwzFq9q
LxFT3ZDrLL4Aic4c6G40fcT22//CCE/JkdN1JOW0VeL1P5Pg9Xwl0RiuHlvIEo+uiefde2sBNzvS
mauq3UVYxnjFm7LrZ+S6ZcjRgWpW4IR59J4q7Heb0hvL/7w9dfw7XttLJ9ZpMyIcFiWre99vLplp
Rrs2asIf8a4rZfOOWR74mB3qpHtvphn0HYTjzEGAmYLXcEB7BxLFXXt/oiHV/lUwnOyYExXi9HT/
f44KlkGgFKaSslVW5m6xgDMICnDvZ0aOLoxu+lbziseh+XQ5XyrpqulcACJhorfcXYoD+i/uBrE/
fxHr+JIwAkiuyuNXSWT/iQWA/MqgxVrAMvTlAQj85RoGT14Ur0qiMYxapPOEhk5vin5gKaJXfC/C
Zltk1koId4G3qfL2JFUgBp17wpFS38xGMiR5hjfZ3CnxQ6qp5PveRGhbDS48DTkP//6xkbN+I9ag
U6A9tPqqgRKtaZEgkL6XpAd4FshQiROgmBCi2Kh2U8LOd9XhrR1znXypneg+ZXyyva3SuKlmYJEu
viNYNlN29hkUfnBe7SptyCKDRUA35s7XJnPCGcb4GqP/EhCXmGZvovPCOoYniJ+JSjICfmPS9YjB
ed4LO3MSwLVwjYhFukxOL4ZwfziyjhQZDwixQmMSbPdhJcww++4VISGgV2fxOXr9xPWl7i/VWw80
r7WSkteSSGtEdVVkc/10IOn0gFx1Y1DAhHejTWOycVPbla2SS6OCEOLpnxFI1dF08Oqaqf9AE7Ju
+Eu91eO/ndQ6QeFM9vf7JRv5au2c04kjGute6VKgrktQQfP0MOdsJKzDYlxQMQcQbH3lswFEhuM6
ReGEZJd4VFkjn4mh5RdfXXDWgiva1F/xeT44f4miSDV/yfhdj8M1MTTbNy49Bi+FxLIesTX7K8bi
s+2/Io8f/r31mzzTStuRmjGC2F9WQ4ly1SR/P3Woekj8TNO2L+XuLClQV3TYnCPsL5ktfIfIHUoM
qgiIA+VnLeiFHhL2G70K1EN4P04G7K823e6u7aa+Cv5mkvSviQ/qLHWZiexNol1SEraKBLnjW71T
sk5B+ysjb2Xg/aM5+QiFXsjwPh6hAQ+bK5819mm84Erewc6N7/xGMQU4zyqCWIwE5GLN/xx9jMUb
l5BK6LOYS1Qz+0f8SscYvZi7eek5c6x2IzWrihxsC3+7v23VXYfWE1JMjojuhB3mGYGTzopSbWAH
3WzWb2huiC1XCtytOELanRFi1qZFt8TrwYzUG/olvumo4Z6ExB2iSAzISUaM8GLbjnXiPXhH6krV
kHGxN8SJ25od0la/yzeHQDhuWSdVwrBRJuTuivsK9Fnsja5bMBgaOTQiqLKQR9yLyzro8AcQebVU
xHcNf8GyjzTSKoKanH1Sms/HMKkqWb4wAJFqh15hy/F4bmMJSWpl9HHtjcoHRhtPUf74NV+wHHZr
xeCxWCKReeWrcPeypOrnYDlnT2OV3Zw2SU8W+XKCUnQuAw8tf/8If+hM1hD8JcZwn5qpzcDiv/1h
+jKEXesw/49IuoBBeuYudjxL7jcU/q/ptJXGBx6dHU5jb4g4VEjb1S31iyG6aCWwplWmMsq520xK
8eBiT4PRBggTLIfWAa9fOLv66kXBMOdoqjdcCEwsK3yqgPqH0hcVBb656VSvwlscFKcCkc1zyQqf
5ydBTqlXrKLGeBQK2ZuL8sr9OFw+uP0uhGmF0kTFEF+VjT92Ob51PjGbLCA4DQTzn0llJNmUv3Uq
UjbnCCHe9KSiOTkbVk/Cq/rt7AbRytcrsCTRfc1skTpTu8UCL4+50QHPqAs4LXgEXO2t81fZqg2M
tWDntua327z5hRcNIxdkjuk+4zOxMoAiuC8n0RlOrpodYYLWK4fXQ9BqENvYUhrM8LsCIermkY1M
e13yvp8Z0kKT9S0KgPLQW0eGE+UG1kniSpT1FKQSz4S2sgBCXOP+b3pY2stDuOTu6Oib90+RGCfG
lErz8IhCN0/IQxE8t3eYHTOd34tyy8nXSA7MPRg2vy/1WmIiGR5nZgOBsPVSiEdXVh4Lakb4JSsa
Mq3vEUY6mSsehqjk8yJ/NSsfNQ1GPX/L5plIVa3XpAydTWMionf6ykRZXevLYLfKmRguBFTw39hC
Ny/Cd1EPBWJgAHx2lvBzJEnf1DW1qqVxtv0jfmwjaShV0ASNmfMsjNpI3/rLbl98w2BNopBZadFk
lwAydH+9VeYWjmHkBpJxjh8VgpO65PfcA+Hk410sbD+HUEQt4JziMUA+vhJGArF98asvb+/SqNDr
rSKE+Lku14FRT+VkipvSVvXPFkXAu5S5ajvvFw8BVLfo2CSWK2qu4muVTIePs8Yylyqe4k2R7EAK
kJBWSCvyK+EmXhmhJBeUMSQ9nLSxhJBQzmBqpei1nwV9xcKjZC9olyPtYkZM/dtVMhqgtDfCtcN5
SD9psWEcOzGnPxBaiDK7OuQsJ1fWuSr1WtTXRClxD3nUsGPucCQRm3shOGoM+Tdok34/Wl4nbce2
WvY02AwQZ7z1NlqrsV0jdBPPjew1EcYGoXP2EhEwp5u0ftEzr0egoA1ZD+SEKznxIQlh9oVZfK6s
mwyUv33o5YeF6V3/PesdHLsFd2HcxyhB0UrsRcJ4QPfW6Y+T1gbQNTxpCzgavts9UyFXUsz3gsyQ
vn/Bbvt3zC9SrBMOEBtq/EFBNksaa5aAEd2ofdIeR34DRYbLSM3BQj4jyGAP+3t2hU59iWNR+tcY
RurbMl4S+aVuvxZq5YTHRRnTFJqUYES/5R5bf2PFtrb6vwM5Y+E4LF6mqvTC35o2lMuJFB06ibVq
qZZ/rw3W7zp83XcbsW01fEniD6skKZYWMKKKfB0iqtYmJEGFBe82RHQS9IGlGGPTl3lAH1EL1d5o
iaa6LdIPLAu1cxmmQjWvhYMRnBsHapvdyWxmjO9rtu7duC5bz1JhGuCl+jdDGDoBNCcGSucWqZif
lyXQpUs5C8ilBSqfHGIx8bGxb5SXpf8jQcRJHHCf3qCRKTP5niwgLe3Lt4qFuNbpR+WOFF/2maSu
HcCtlX8H13FLtnKLFcPlb7O+9PPvgFi/Hgjv00Bk0BMrpYGY/BS3k2pHynuhIdQBB9Mf7GA3XL3w
v6w8bK+DXQi9bSqXYnuMyMhibmDoZx8nd39p6gxCCxZ+OJSWu9xwHpQSTpRod6E7IWLmUaT6PMjL
2NSxvy+3t4L/qJkBjpM5AlzbFmSG+5kURXRE01DyB5o7U+A0yuoRtM3Boan1Ro7IkL3T+y/NN9GX
++5n+YxcHTHVkixBvLwhBMsQUZVbjh5hBS03A2yvYlw8UjdA8LjIftk27YoFcxGmEf2W/oUgaG9i
dIGDk58Cllg0ka3JgqF+tCIVTBhaQkr10qqydg21T10gzi4LDL+lsJ7PIKZy8UEACnZ0Kv+780YZ
qBe0/haUuBOuiAe+bTf35GE63BMME+6OXKRqyC7XDibhjX/IZvaDyJaux/Fg48NvZOUIXU35WwLE
SxHOSS0qV1p4ZU3P9ZPMXDT8eLNwChoSO9oZ8e6nsKy7Q0ATpc3j+ZAO0hex25tEO58lrLxaFfx0
9VekP61Tk89un7J3n990mym1Dq7cOoqVR7vCUEHkcsQvrsG+CiLQnPKfy7uN7U6PVoInuvguU7XH
iijo+eLp/HWSnIr23ImqqdQ+Bb3+t+tORqBvVs0gAyyI89KNWhRCwA4uJVoX5AekivvZI+QLm67g
eLhTJA9AIsZEb6w1rDJB8rEJludCTYpsqKBf363Fi4+jAZpH29uFecQMHc+pRnsP+dfgjXg/rhQd
3GaWMCPUj1X1C0+cLj7rNRLBGV8ynTe0HhUeI49SVyQq28U8ZaC8AZ6IuLy2Ey6fRC7tMqOO4rXw
8QMeMU8ws2FzCqw/H35NFFfX4hC2fsnnZFJtwKQqBo6Yo8WpG4C7Q5fwdYQLEFNgaGwEwW/Gc9C9
+s8hnkKiJbJ1c9PkZA2AnmxL7AEJQKFylN6WTxs0XbELlqA1Pt5HVU/b8XErAPkotri4DiLgQJ7K
vtFFD/BPQY8/h6XNUjhiCXvandB1GrWRkwNay4XYhv5MgvIXU271umLJ1+QnNf+4xmJVqKtgv/TH
Sf0lnb10SS/10OeDXN6TMfH1Rnco9a+dkTJWWxPl4OoXXZsfVYf1DOUxMNdZytxCsxG5aE5OsfFc
ZSEOoPu0BDpWGk7PnxpKDmepTAUml3xAXdd1MBhsHlb2Ff+J7O0ZGb/I2cMTRql0DPhyvyvwcY7X
eAHZIvk4g2epaQ331EkEtyZ/8NhnpzyH6rkJxAUp40R3/nNOf94FCQPQpFYAnDombeU5hx2TMA44
63VnKQzWCqfu2jfyMQLyJv+rZtb9ER2P3Zoi+1kOWBqpkLHYq9p0mAV0/ARiO7+4DFXn9siWobty
VDwpPn5RiTALAJBE5hG9ncKWRVhV935ygltbmpRpT/j2/xBjhf90n+/D4bJBSuBSqz6NVBuYr+4A
s+XCjmRmj39e94Is2dwmWcZDcbjKaNXr7Q0r+hSNPc99QDQUezhFHEnCn+HYb045TI3MVQjAErsf
L/XwjZlNiueMQyQo+C3+5WiIChfAf19/QuEfu7IjJRMAnKyn25P3rP05gDPOGO07JmZ3dYYv9ukz
D1gRbWTe7zo5Mi25tw7HjR0ft8Y7IkLOT1PSxhtjFvytZvWmET9ZgA+qgrO66vy205NUaj1lxvN+
Tg18XC96d1eP5DfrcyyGjt17FFaBphUORbS9nibWI83Rwk42FvLM5+8blu82w03vXJV4J0c59ybN
2Q2dogIaVMr3oqm0tFHejN87JBtM/jKZuRRNsY3S2q3JSdILV1UqpbjQVIsWFLlHmeUHqOyTzXTe
buMfuvccU71YU9ZC6mP0C9rKO4htowBsXDYzfz6cdM37QLCUmmuOvFyRhd1gStXASP7zPOCF9Uqf
DAnMaFM0vwlaLw1hZF2yDkBdtrVdMLAVlZm68OJBDnX4vZjn/XaeGfy4qPxLitqXEh0LBFEAVuwm
Lar74QR3jdhexDmgAgSM2pBTL8upkKBsmIHU8lZaFm37Ve2md6/6kiN1UM1SOujS0ms31d1XEBzQ
fDd+gN+zjxupEBlobXUOrl+RRBzKqW7fVySN7VSMbHDbmbwv467CPiZ3ZJmOzc8FOmQquOJRYhgS
86peoW6aL8vJ8D3WFm4XRRk8VT2217Q674OYXsHxl1UA3wux6Am9RhDctuhLh9mZIzS/5nXX0qZG
UomeCvoUcGrl3snDu51x7eMBLgeR3gfN4SaM22E37O8WBfBMXmUpvWMqUrWhgtOOz5xjQ5PGLfi1
PHGvmwGtGttvoszPWPS/8EkqB4IygK8urvglIu86y9DBRgT1/RBN/0w+k0Qps3z+IAydxph6ezFH
S+iGze+hO6825KBSbs/E5t1WF9WDFUiKjQ1XF6mTUKcBXZCdTed8asw8uTcz++6+D0biaqHjNCn+
RuT8TghXYxRt2C7h6EL622G86Vzuz9AAGR+D8KVxCF/OujakOzQs4n2s3bfe5rbi5+7Gn0ZP2rMK
6Us8LcF1YPyuFj9H53dN84PR41yjlBkKLv17dr5ZQ0BghfXXB11WVXsZAyLE811gonUZ4SKWGYnb
NvbPxIwzfZLZFZg8U4QOsuy4500C/wRVi0Az7nCyl5nzlqtZocYPkj47eaeW9Q/J88m84pScZ10R
rjlGClGXyVsPJj4wGLvt0k1/JJW2cEJwuKDHybPUAZvdwAC88G9og4+Ow7nWnKHpWxSbJ/WUdCMX
vOp119bzFYwHLfZDpJ0O3sUe0OJL1UznNs4CM1tu5cOMeycQY9Ay3BGRp+mJN8dBliWivzcpfvgV
Z7hqz1cNQkA8iBH5DH7bcabSE2+Ykma43M/Sm5sj3fPRf9SyETN4mdgAtIT8Rhni6Zi8sS/MX9rL
gacWfvMQKUbOR1qjaxHA/cqg7LRH/rqoLp59pGL6vj3+NpNhK201iBKemP05/qYEOsdrEmdP4ZAD
ZV9uX1+2Hom5HQbnda1Ar1ZToe3OdYnmi3bgTKlyhFbtdvnLhyqsWvwQAZBc6u9TP6caO3dVLQwJ
6rQ/Zf4YUgXM09jdHXT+ENbhQwBSmQ1W6iYmlEJ+ijIOvZQYxXYqHQl3tZIJ3WjzPaDh7FFX+iqS
ofHC02V1VGvLsscDsblC5Atu2/ctySHxH7mmJWDUjy5pUNCxcaaJUTnqIiSqwsqsDL/AIBBQHaKj
rY9DaKlT/rbUKYM//WrtEFjp4NHsBwQ6tl8Z2pnD44UjhC2lCV0L0OZUQYbEhlkvuBOdKb5qM/03
LelzMDQmEeTP+Y/mrcqTKdJ5ES3mJ1x2ohQdQpZKIU3CCMS9WyoGREyZJrBmayUK2xEEFnUox5je
Nh3bzsoRIRSAyrsymoBS3oqu4SU2kwB5/hkPtXnOAjFEuBvBSHzNFZJFQ0I5Mx95HmYj276aJUlw
dN48kDhhRq3EarPOqW4c1PosB1z75t1pmK59sJY+hI3T6FiPxH9J0kDUJnx6z3biPww8U67FwdKx
gHfcbAsIJ/CYp6EAI8WyzVKwr8zhVMVXLOvbVoGnya78wElljFn5a9eXPmb9Ww8T4IovJnkFMkk2
/8pi8eqzu1z5W1Fo0ltYlCT8ys27vaXEaSYWfEMWnoR+nvINqFplfxz0opczSZNiyrp1SGBOkGZ1
h30bVzDIe2qHCb6304PSxKvUZMPTxf72yhRIJTdrBEwzixqDW9mYnfiT4M98T9wOpHkgnxo937QA
9NNmGQYv/qtOBJT44MHqZ1mMyhhaF6kSo4SExFxGx+7FKaTsptbSGqv+iRBMLXu379Iot5W3fqM3
kVtSH0L+GMYXk9BLsqYlKz0dqScQOx0CgW5ia3HpoQbpC8S6HD4xBKYYpePlWareIVmxZmZjtxvZ
fdemqY0zTcWTy8qyLcUR5RHlCH0npEVxAi/wg75e6m7x6zXQa5F94za0lAJvOFbtQNxR3PsDGFff
IDiIHOYRtBdvSWsEyO1hxj+vx3Vu4GSLFvAcmVM0D0EiPTFERE9Jzt4NnhrfpoQzRytGWBzBmT58
TelLQ+YDRdvSWrn4S2emdyjbvRQnVDGd3Tu5FsewXwFKL02D7x22jXC62O7odIOwkDsmEAlAZtwr
i3Aa+Xst8vOxg3tCI7dcEBmucawLffxwe+cY/TFyPO3ehaMgIJZ9DQiSTJz1W4gNJ7Rb7a93Og+U
LYP9ygdeM3WhS7eyLr9WmU7iX5shOjP0kJdRLJArAH0ceIzXhZFJszJOCZ2RXcJnBV6kM4ifBB8g
sDoWfIKpGSEV7MAaEKE6OBxmWke4NUi4/yLtI99AnhDY94ABS7QQrv+dw0W0KQZlwlYfbc1jtJQ2
v/ImlejMED7rmtgAcej+XT90S7zm77ahBpi0qkxuFwIe8YqNX9/dKtDLj29OmiKyStcFQ/a6drQS
aKdaEQznefghalBsj2fUt53wrPp+nqnL/R8QYCQYDgUG4qkezvrWE2kjeBLxrdRK/4nSPGxQWnaJ
VmZN6XK140a7cXyZDNmMVDIrHx41lOSRtn5Fq7/qGIiNtBQCh0qzGSbOoGB6vn56ekbhMQwZKre/
Br2v/KXTdncxn6CUThTtxcO2jUVhCdihgxCyrFEMyfjREUpsHnZMR8LEI3g07J+o7YZduseZAlX5
jZAcX9/Vw2WMF0oOcw+SciEbuZtEASyz5Z2JsXTh99c1mXhUoMBuvRI1bf9xLrzk3pyIG8h/bf0L
B0u6O7U/szzLSNBhh/t4+ZeI5diKacq4GItwhewzPtYfQzmb1gCXeGVmg2w78VfKEzdlHY0Fu7oe
1wMnFcwkKdpJVwhrkQhPH//KfpbyusPX5RitfaBaWoNlg6HbMj1zM5c9TM5Hu3bv9XjbVCkfZzim
wpxyvxGNwT5JAitl8TVo4cUBufqJh8ykkd+cGOxBWAQAFxihS287HU+JWTJgh7X9YCnm0rmiDClj
Fvt4lKoaCw/A5sHB8F544HcXKH4XTMbWooZ1fC/cvjTXFrRe3gEWr5UlU3fUArKT1XDdJYukYheU
65P2foSjRnMcPdB5bsfAOOXJlC3pCHXehX1hNAwIOIYPvkSc5pUsteR9nbG3/o1M9W/Bm2LvsRaM
NAyASD/bRZ8AD8672oL+x9XkUI1aOMp3WijXJqoV4sWQJCXHuGVaXv7ZUoQa590YbXYErqv4Gzvt
PWky228433zOCG2GnA1zN5anZN2oF32HH9T1uAwAlr8alMGa/NztB05tmYAsZgCqjMzhpaS6s5Xv
iyQKukV1WOY7oxL0doZ6rhE/sFu+dyMou2h8SB2gFjofju2DSEDI4CHgjUAr6sqeVGHnmBbgZhzb
+9pItaRJXSJo8ggE0Y+EQfnwtF+2iuRcham0S86S0Nioi1w+8+0r9s7vAoinKwyt3A0elE9ik67f
4e+hsD5+P5OWFkhARxJ48WxbbwsWIDk8sXWBF5wNI3bwm4au10nsicd5F92ss9cQsn43YeSWF7Cn
SHl0u/+mauVzWFczUUgvpVa7QNZ2Xyi8HhrHyhYwDZaEiDWZvrGgxWKava5emgodj8BsSCDK6fp/
n1v123tphZJAseBTFDZXjOHbm5zkKFTwAhjmEDBugZxgSc/A31dmflDYlwVoyRX80+B6ZQy9uyae
yD4TIlpNZ8mm8hmt83Hqyq755YJbVxwcoCRCxPDbUl4EY+/GWXqxcFcaprO2ERWXEbT8WJW9D8r/
TnrpGdoV60S06pdyXqniQ7ucMcw9piEvqduMY1KIrZcnexrFTU7ug7l/a433gFwKgqvjWvip1Spd
tcJuZpcRaL6r5rOhDETJCqbwkAqnvE4vXpTAtu55K7kG/N9XPRNkDkxBIrOJD2yuQvHl1UGu3dvg
KEcZlBZgxaOpJjQHXz8nP9hMyViqgrv+9Xa1ooiqWI46kYsDIM0zSFbeqqxf0wPdhNDbgISDgLkO
1dZUrLcfvSBJ+/XOC2OXl4tW61IgI2qby145nNX/tja65ise8MjksazZKdtZwb2BU+behJ69g0XU
b4HQ607xTll+/x3bKCwEpCMNmUrxic+KTEdkaqQ6/tmZduJ4LdCmpJYK9ePYr6tzplCVEQvNBkjv
4Jy1RXPiqRvX8D4rg3RvmuWxERsyec01jFXUpfud7IwlN4qO/ZinWaeS9AoISHnc0+eErEEElvut
bM5u0JhtXiPwHHQZJYMRza/SXl+iiQ+brO+doUnmnejlXYXVeVVqObzfr03tB73xPtJDp8fT1YRE
9g3Me1OcS1/ofWBPEhhSDlGdCpXAS2GoUwc1529yUbcJ9KWwMcIkzhiUB+mtWBnX+aj33x51xuZm
GIkw8kBx4J1nfUNLDQr0XQPmZcy+wxMTxbFNFBJoAezqegpVk17ZTEKfTzbk3uxaHFIvpI/Q0QLq
t2uweGEZshfDmU+qhT8SkADh82LAzcOCFRkxPd1pGKWXwf2bPhpuMLknWVkSirYLo8ZEeLg+wnlG
HFf4idIb3H9Vngkd9mnLtXlffuuRmh/ip63qUsBxzSp4pk5AlxvjyAJY7xS0/3fVHWEWPlRUwEcE
jZaNlqj51hko34/3hx3DzDX3+hKKn8zZO+GNyGoJ9Uq9CRTN1yYj7LadU8LcJ4Juy5CUVGWfW/hf
Dy0mKalxuw45nI68VayDtFb2+/Zs58yvCzcdNrBoMghMM/MawIaZ+6sB4w3Tyln8xVFyt06FtMUA
PknzYQEJTYsZoM0WpfdRtmKWUjF/qv7N+C6gQOXLiogR4beWmzs464qK3N7Elh40kaIJWDfxarWk
G62lpacB/b9fLsxmqgQyqi1iDQUMM0dI7I404qnz3K4iSr97TKEhQlRQgWVA4Y0rv5BPbOVsaMMF
pcbgqmO+tSVe41UA4MJMR5gbiq2BvPbboSlZpnNa4FnjIs/Y7FhtinLJfVEU0XaFsj2Pq/DtLZ3h
DO7vyvIT3XtYqrRnUch5Z6bRmBEVPULSpu6rI2JZ0DyGi0Bl9JWvN9w/aK8eaX8eHh5YqDTuifWA
i6m15N50w4IVotUoQP2mhxEBmFfFkVmbg8eUh1ra8dBiUh2JkjkEPDrERd6CJcJVVbj3R80Ct8Nl
8fBBRyk2QJGnpH/aOJV8BXv88cw3IuQSWqbdSFi7q7KuOcRV6cMsXPzE3cR05F3szwQahTxQW320
wr6mcRee3/raYLEnY9ujD5nPayo6Gcq/EYtKYlwFgvVrn0o3uiSwyLSgFxSDHHD+4BSZKfwcgQie
atBl3Y0R8WGDVcO4grWOptlBaTvV+W0/OvIZE+GqzbYM3W9WKEh7r2SWI214GhUk7S94ucUwFJ1r
R8mms7XnPYS+vwrZzLmE39b8s+55jQ3echyMPS/K1Y6rfKgmEf9WCKwOpU/zKlx40ciPfhYw6CPs
RcLC8kMge4NNLaWgAbG1DijonGpIwQJHwsxipEuUj9Q/IjdSbCaoiwO+rJ8isZkHePcKiufntWvM
HM9cwOkh83tUfXre9TyU0rHFZZM9NwyWZrv6g6bYzVqbO8I037I8HKU2r2CR7m+AdootEGowPmuE
Ecivk/T6uKTa0adABIo6vuT4yfJYCPz5xply+mcZY7jjjQ+gjjbMZPlBTc3tUtYYKcvjLC5e13G2
2nc/OLs+2GVexy0+VouAH3FVDTOLiWbSuPgmt3VBZtueJc2/YUt024fL2qtSiMW3/2mdiBC1EEAH
qn9/8m0wqHNJr/4tQIWtfGY40kLSejPzf2sbDp91b5gOGkYAQQxP1hBvf3pN0YbWhnOlShlkuGAY
LOYXyr+ZopWifoOGnNZbnWtkMHvxHaV7yFrdPB2n7wPBoRUDDyo7Cp5HKRc7V/rsOU/bYfa7I4Zy
5SuXpcXm9nxLSjyg1XlR+RLyjeb6ZqUOBs1O3UNLArhzi0CpiNKnh73xUL3hdfL8P1QDTbFmyMha
TL7Z2W2YnAL5r8QuZbmJIeDDAWfG5p/7W4P2CaLq1ejhxSK+D6dDB18y/45/rB4yRaitz8IVl2eP
cRex1MUdQYXXyDcbXXZxy1sY9nTGV+uhPv8oBORQynu1mXeKw+WnQtfIbab764Ub4m+7d6aLn+3I
vYLVayuLECuI67OZ6Kpc6UgZq3HdGOV0aV4uQ002TlSnWDBDSYPVPGMGWWk1sI2zALvRlcumGqcj
bKla2V7kI6IoE69GBTLITV6PRqUdgfVOJe2HHcaDHX04bk/tRd/wAmgKKssq5wcPF6RsfNDGBn64
dohF1bmqR0ut33pbj84ZAf3bNFXonaw3D0MVnLQ5Fq9V75+lQUp4dBKb2H4dRZa7m0WqJM47XNA6
9uxH1Ma9AKz8+ErF1RInAo0w0ZKHroggTGqZtLgP5R671Q+avtbyffelJF3Jf5du/zbmjH/09oCU
MYQRue2PBPym3OrTKDlUSVda00fwMhX4RGiMUB6Gzk782IwYKUhCnxw7/pMlT4G+YGFIeNS0kDqJ
O6eYRFrwmKPoyMzHDP+7iOKkxL2ZnLlTkfMucQcuqUVNvH5X/WjObds9Z5myFU2V8q3ivtdVGC6U
SPQAzK6G0w3AQwI6MXflw5rRT/rzYA07iAFyyfroQeDjf1K85308H6RnppqJojXc4shvtWbBKIs1
qPLO2VPHDjAaDaEDsZfzP02hF/1VDbG92DebCN2pkipJNUzEWhuyl1LFeKLfL8b6aaqQVEr08uCQ
0YPMrQtXSbhvBaq46UGUbpn/eWd1G4K7/G5lZkOcIQhf2Cn9EhK162orzgEAHKRQSfzI/TYRjOiV
0oqWJOyD/54fxoFryiZQ5f5e2uWECTIUDhQclMN0nKR4WyphVojseaG1bqRguqf4QCJbsdlXSvbz
IanqPAZlT4UU1cSJzHQ2vhxxE302dNj3VvW0OwLL4EMqrpE7Nf+duD1HNJZ0xERw9x9hdblok4fn
OiQ3gxuBV5tk9GMqWePxi3DlmjF1Olf1XvifPLcmXg5TM4a4nNlPFqxOlCRZ3MzFU7GXdynHAa07
C8nacGLeTQ2sAoLsFI1zKvKN3mfxV5nJ5E9d83qMe22QSQzTMwnVy/nBmlEDacWJLO9s8bLSEnzo
7b66OwKMky3SWqVq3eYWLTJOgl2glEqYoJvb1UlTKYLnnqWHdiiHRCHIvmmVDoJpJ3zcPgQ1ZH9J
Ng9xeg2Z9602f8ef65orJmvk+uVziscEY+zGHz2ZocEXLUnn0o0ecDwClAwFCkyWxntNqMZqku/X
htqjJHsQrMZUEXL6N6lZRK5IZ3Chy5ecPZsW27XWJ/AbFkBS8od7+qiqMETnJaFdQJKqps/nmXGK
v6t3YY63/HzG1+0DfgMMBsbfeWFz8capYuCksv7gkn5JPe2QhE7VbJuydqr84UxeFRSCezxoZgsx
kz9v8E57MU2s9fSjjvUzqa0hlki2cKj6D7hRs/B74RhHdM1UHmubwG3xooH5icsxPdWPIDvg6BUe
nl0kBeUBROBeMH3NBbJqfmItmmw4LF9yLT5twB8AoO5S3xQWbhZoUTfJQG8gZCFhB4qSvdHmJErX
QkNbpCPzIPfGYGXVa5AyJePksCt1dsmtN8KJKsm9yOBFJXlSZ1IIRkmTKDTbGNNV//6UwZshKM1f
etBKLilIe4MBVg3gVdY9pPtikdoG843XoNS4TZh6TDWsvCIyWYUiDPiG3a4RTuVGO9JQHF+jzEW6
iiHX5p37JqQPRH/ED7r+VzL/YiniiJjYWENc+xdL/yuU9ANPPoBdy4Mtb6vTvpcpAX420QxwWI27
K8b2xqFtb+UsJBslcFzQbyBxt2k9n+uCKHQQsBEyrdfL6bAgAxgOqrntIXF7RrLnlcfPG0onu6cF
oDVC7UZysmJC8rjz6fzrYLGoTMeywJ4Ytt97G1eZWfi032s3R0JLXNBIMui3W+B5d6UWspCkT5hD
wpou4kxfbWo8TxdqIlmNJ1AIXpwc6n6au8caWLVyI0d3iylH4YccDWctpR6f1ivABxY8Wczpmmmj
8hqIpAGB4HyVAQ8FISEXDngE4/gmuDkYX8/19qCnAP70cacAz57TR3yiwcgwNCZ01OdBXb2WFEyY
hNHH6DN0i9uUjPtUgJM8h5qZuG26Ja5121uBPjVVEB/a23vo/+jF2K5nP8YxyJaa9StqSlyJj7q+
sZYj3N2axJp6PfXZAQ/YLTPbBjjBp92YK+AkH5yca9XEi95sZcBoS3HTyqzEjU9U38c6E0q+yE9g
hd23acBUT9WdzQjtEcXSoMbbY34AglVzpCT37fKG1OgoOcLbe1LAifXu9tO//XRAq3KNIaRZQ1T1
2k9zcNGpz5skJruRN1LJqN+TvzAMzhKD7xrfFRTYttC8Gk/yFDVKrqUWCzklBJqW5cqGX1+ARtnC
SCXTEmFMpDdtio6SqAjerkacWyF2hdJV0FSBnq5WaO/v97cbFlavW6kWzwAsEITBj87W2W08ihNU
M/ieeS9z4reqcbJmqIU4V9MCJpvixKLVL+5aHbCuWJe74UP+O7hkP6pWG+NeU/B6Pk1rzeaFGvt/
xUEw09t7CENMm530ps13txtBsmFIV7G2zBc7OvJXcTpbc/1m2764v0g/wFCBXdWLqngOzNu1eUsM
kQzpUt8K3d/dIuJ9/wXpPrxDfx90NJtvXQTFZyre/5seFiwt/pJZQQ1abnOoOTfq3+dxaYNuyyC4
jsyGwUo1z0vQprONd6cnWTxsXxuUT/9vMKwhK0mqKTB6ZG690BOgS2Fy9lRe4H2wJzog/WGvXwgQ
ftMxWNr86956o0EUVUbJJJLdrNjgIKG0b8IxD00SNezYadwOIxB0aKZyYcp40NXVvoDsJdURKpdp
h2F19JZCjWoSrGxrxZ31Gc3gobwBWmG8xaLHAbEckKzZ9DLQy0Dqxy/7W7AOm68BaJ6tRb1+DC2z
OlxL+L39laSRSrlz7sLcrvRKmMfazDhqGXSQPUI85U+zt4J2nd3/eQ0qC5ULwLIJH7TZP6QUAbjj
UMrbPfHkwMdLu4evHxyLxf+TRrTMH48c4BjvWup/wT/90AT25l3pzGstPorgLq9w3dJ/aKZ8cu0m
ZsIIH3QeLl5u+tSr8Hf/zFvMDTZ5Y8eyo88HjH4H10P8FadNv5xWqUKzrAryb0yB5bG231d85FSA
Xc1Kqgl8C680Jc39lg0fr3PW9xFdCYXp7S2Dae3MuXF/S2YZUgzncYX9zNMrbNu2AamOw2OqptmD
bsY4qC1i4RO28mWET+y9eUuCxdU6QbvfO7BAEpZHUIuccpAkOyv+UrTObNgumUQWtlaKLQBw3wYO
KnYEXF9bp/ZSGv90cox7MJIIuCPHNyLPNCGkaNQYZDXWOIDvQmBOPrULWXwE74v+Ih8kp6MtCL0c
K+7hzVqrG8gARw9OOvm19bHJPEfQXSMX0ClX+6Xx7foiiSD8bLiyMITHh8Zj4awAJenG1+bLIHw0
Ww0JpJ6xE3OwsIv2OyQHvcMNHxZw0i9eZ3ISqdNW7gY9owYDLRJEvj90MXpbkubXGTyfKb5xk/kr
4xUjwpbggugYK7qHMW/BC/++IuwEPwEe+BmR4vEHHqrNF2EbAhNmdtfXXylKSz/dIg+ZRk5tU9Ao
8YY9ZuOF6eiHgBVYy4NXlzjDXgswdfKAl1Mb7dubjZu1HMpfQx4agxEHUGB79pwls5YFsF5LvkiD
B32Pt100jmp+2UC2BzI/GtmoAN2WWmjaCt3MqZmlQrKFFnBkA3+mPBs7UaOFkKrLLvV+LSwDfCKS
jTpiDzhddBT80gXGWZuNHdWB/f4I6bedSZ7FA7zio4YcJnn191cwAp7yGo4bApIa68GngO4i16qg
z09NW4z+26SozfYh4/TPg6O0nT9OnCcNVHI7jzPCGIR2qHxcC9FYUUVKnTrl9fU6bqAQDqZ2SpDB
wsHd6dc1j/TwRDgEmiNV9EgrIolXEnR95wD3Xah7/+JGPxMzAT/tSxrdpZ5uArrVNrYQVApjYyeS
HLcbTF1MwtLk3L0d1XF4tKk/ZQUnzVLyfQSLbibyfCRQEw69MMnICp62BPp1mDcoNHrd/YM/O9yF
wHDz6DMlmtsjk7SrERaRY/1pvxpDkbyKQy0HdFR8FKvbpPwcpHyT9Ind1RL1D+wmIGjuUD/7OlDN
8n0HhZDbaG1VbyPBKsQTRc29KCGyfEsvbpbgKmMzFoFY9OC2NWDI0tlsmMXGubGLAo5Gg/pRIMkn
2CPw2D8ZlZ9ljUQEf49ExnNsvL8PXQyWu12t6Z8o3swQPQYA58FGFHNHs44TlWBAkyiMv8A8Mat6
ERqd+Inrhgx2ekA5vW8w7CjD4QTx9KWys4d+0pWieVFX+/7SioTTZoxN0W+0ZCRb+CHvA2f4px4N
BG5meBzE5v2t6Ewv2QiYpOLp7N5e2vlEY2z0VyFSi/v8YbkKk2HRFL2HuN0wILy4BCH11j0lX/wR
NLoYO09fyifpUQGsa+Tkvk4V/6EnwnRDevwrcvQGMQ5PrOQdc2tBER5uv+pMxR4gx+VyFx/D3Duc
nnEs6WPCOTfjnGjwIIRc5MLbMcurZZI1OLSmZOam+AP/cOIBtS1TLo/LCgXEAIhEP+TL8dLra5/Z
WbjlW9poURaHc3OCjRYN0BOWbH8Np5F3twjd2luR1qqX0vNP6WlimallSjBlz9pRwcGD1vXpI32S
CZC8cvpTVHliz30B9IopgT6hluZAHhsfHV7bnd1k8ACcW0q6KMqEADwoecNoaDla5weBGN44v3rC
pOVG8H4m+e3hRpqna2tHPsbThLEF13lur2lFZnrEfWK/iJCcJ+YLcLEHLPKIKsfCBtJY796+Dq5B
cQIj1+WWGvQNliWSTjR8Ix78Pwe37uQsYJNriOorHxeRfyIFjHYpr8PmEWC2/R4iUXQTF7TywyJQ
OpDdhuN/IN2tlLx0iH3aeRcrZ7dFSYoebudNQe7YhjQ7NyBsfOa4l7jWtxZAlErTY653xNIRqRLc
zuuInFEug4hKEhUZKi60hDvvtSaWTEOEGYDL/kKLUyhU4dDdwl/d3kutZbsjFn8ZD+MQFG5sTkhb
3bYKHxUm5IqQNM5eFMzgaEVapXL1/5v0ZEkUAkDgWoGVIyU1WOtgPgA32bs467HrIHP/1PkBWv59
DB47D5fIy21BFj893mtPx9e9WTzcjx95M92RKDxEc+CzMqPNvlvbS534q16XovHNusvXHUFYJeA7
dnMmcgc6hNn9uxjxa13qQn3LD85JqJ1sYuQshCTNchkQsl4PpGzxNwgUwdvUn1iBpuBcBnPS8+3T
Nve+bStF4e64e5bsgcfldRRArWeYObhQbsUoOvvh9YnAgTNwcCUtp5FrS6fsaPw2d/puf7K/CnwF
GeIUjTeQUUZ9lP/Y+L9cnChlFWWWLtANh9yXITkxa5CJKqmhxnrZFPTntxmnRwshdfLJ/0rUjRY1
5xFWxYhFbSWGaItxQ1DiZeXn80uR3u6kPnK+FpBxzNPovckGeGedeXjaP63TzU4AdSUwTPQwveMX
nt/5Xyc15SW2lSU5F/wrm7nAcVHVeolYtLXz3xLJeSWvrkLAVzY5vN7kfRn38C/Ef330LOvDdyLJ
61K/hA+/thAXF8lMZTL8Xz7Abpud8rkAqfUTnUrkoyOsKeNJddevId4OnuBUc7/Inb8u8Q2oUOHX
fZlI+FwVMQ8EolK7432Y7Fh9KW+QXR+Lm7jHw9eT+vLz4OqEcJ/Gwlqn/W1nwMlGeed4Po5HapFX
AGZ4+p/wNap3v3deH0p7rUnTtedlAOcyq8W44t/QJhp1LcQU+jCU6dNc/Q3q1MpB1G8YA8iLUE3X
1oKJiOx7kkEs+recZe7BYd0xU/NNO0vZbzbYFoJ9myWxEGSyeZBZXHp7RK8Rn31wDi+LvQBRCn1w
nBkvVdZ488m4Q4PKUQDn8fp1ck8uMLLK+GehTmgufb3A5C/UyLWREWgjeF0fiGfq9y5ImOSWqs5C
CQ7uAaI4n8I0Vh1XXDUQjC0BniP5eTFnX4/JPvrdLSnb27x/hjIH7662CcCLP0QJE8aPriA3uiS0
ddK19OKTRzX1QqYBGhvXiFjqbRoygSwD8IPMRo3lCaZ+xhSbmWL9RGhMkI6zAs9hdSemg3k3Gcpn
SKbsuo8Y1r6CX7bPQ5odvN4k+VcnppGz9EaUve49Gvq7QvW1qWRx/orjMuwWHa1SEed3Uqx83CoA
5K8kRnsBikFg8IqZi2Zwb6Pxc1vfqZl47V8RX56toDbsMaCQRLUaMTlw7O0fhckpcpCkiwt21k5X
GTIwZ4IyVlPlDPZYMmziXWQDPmk6Tw/uO8NCJFxowGubtAQ91Chf1IJuu4ng2/GAm0dXJYH7ftHj
A84gszCqnD75D/WloVagnPWuOIjJ69TbnW/xAKZVgV7Yim631VjAe1SAxLPdgYDd01EPjV1wvGGo
WDIabWVzGefP+psfFGLDSXLxDfNkTirLftJ4zFLdqeh0BoZy2YWm824BHkrTehXJtukBeKO/N8x5
5KfbEyU9MPRW2TgiRpUfp5JTtQ94IydzoVOEuyDMwSkTAKm4rNUD4KAksC60HFKg9Vj5S9wE75Nn
d1N1/VIH/s2avNdO7ZfO5lQynhdAhFbx8TP4TMW0Pd8mbYvjWx49qp7diah5AX+/IIACLwydJBll
sbGoncW0/lZk7kllkbg/cKZU+0kG1NE14TqX0BTQujcTBjVZCKgToQPIlDBsBrfj0oI54hmQMIbM
Nl42sTXhhbB3Rg7KyjWsGzRb/SZHjZ1mbW6zZWxVpb6Pm51RQAOJD2nswS/z4MwkJSK8EAZV2yDN
B+FkhCtT7WlD7u6wBDVPaYlmHnQCmErZul82Y4nYZ66jW05BYbKz8SpeX0ft2CAJYUG+FETEwdHL
sU6AfArAPMGroDfYEK+bqofBHvKYS5D64ULXHuWWX9UoA4VzzLwLDIbw1MzCQiwkHLcqSNVtVeBy
WTVbi489J4KELHRCjV7cEqWAu//GJKoMjbyDUofKST8T4tQkZaboUOIMjEAuOqARHEwk69Mf6ZTz
5LWfU765d6yAXZ3DJQfFgkPBUuv/cUmbyhVcSBXdltyJw615YKJOJ9yT9WAQszuWxp8JWkjEa+DR
hIV//WjKDbHkt1JMppO0RTH4T7N0hD8NUx5/FSVDHfiXIKRGlNYsKSslIA27+4DV7S71oZPKJvrE
ktdHpZLgGEEi5bTdmjRr9vND0t9Q+dAZFut6UFxezrUFuS4kjo934VjsJIzEu78MuVAHSuUhU8yk
XMlcxCNtGOkUQmNZ+4zYPL8YPUH8so1FRYT/tMzYL8E5cjw+p+roQfvKiZY00MMCCJ/UI6nwsbWA
qy2FmKKLrtTxQoiT6UT6kapewvbX8vFdwNK26Mz6RajMsvv2MiJ9QwVd82Nt9kN4W+6M2uJeFA4x
TOECcYindbYYEJ62Qem52CBKWg78ADhkcjIeA85Vi5Xk/XYye0sWn1QiZC2MIJCqgeeX5HyTECFV
k0TzLKpbRKktLdLhanXuZJE2Ma9jz+zTppbn6QhotytMSiMv8472SQeE66W0pRi3pSftAui0U+w3
Ssr/OPYsmJ5+7rDOX0QJpSTGjq8o7mtXW4z9481SnWDE56iixrhkbOic/r2D9URDaU+36/YD8/y/
b6dKsnLODLLjFlqtLL/7dP3zld5zbQZeQ1W7i4bVxLxyrl9F7j5OfNurcjHLSA6Dh57cMcHE4JlE
32LbUaCVy95Wy39QJwGR2SIn2jmo+PSIMbonA4BDtG2UBhETDpLO8dz7NVpPOHB3CgfEFUFgtE3Z
tBsFHv4+sw/sX+uyxFUoJwSFsRDYj541mOcbgx2CERa5jgL0CWSWFWH4gtSDJJDophbiE9TixKsa
FXdcr8qiyaywunfJQxJWtcfmsstE20pN29aGbl7waCG4U3ffRDmQgGamuYWxam4kuxNcKnKQM54s
/2cuZD84Wg3eWmkmVu0xN9wzUkGqWxVPb0X5KfRf7/ih6nB0fSA8YZOy0TfSgkRMPDdtuCGAudy+
oxU1pM+F6d98bFJVUgFs7NWoTRwSVA9lpRL8DZVJg6r21R1AmVt28rbybZZBmSAJAkCw9T1E4amz
mWAKja1l3+tRhSYvcD+J7iF5USKNHyZ9y98jqo9tGTBE1MsNaxokAbIZeSqkazb1CV0gUkOxOdYu
l3rAV0Z6O2+tjq2DdG+c0ttTKPiinDatjT50DUUlmauXWu/1XrC2/VGNxwDPsD7EQkPLnyk0Gm6a
cdVbUkCSBSHzqtSkuvRfA4KJR9dTVTX3sOy+iQQLtu7mC9J5orPdiGOZxXyLG+GF5yY9GzRM5d0+
pVZG2KIDHUnoLtrLH10itWEsEiwvy9PVekAgPSUyyPfFK4C/OZrXzvVEPzqICERJEKFDg13Kb/yd
FRiszQY2UsyQN8vD9c8UnguIIgI4OvH6iEIDLv9gRg9Dklpkt0tfAgc7IKdTm/UwuJykrmNwxe65
Jg96TFY0RBcaWgNoJCo0TSahX6xaw8icW6k136lJmaGaAjt+8Ihjwib0cuMW3bLfvTeC1ECsj+f7
KtK3iyuSEpdRUC1GlUsdyLVeY4FTeOylQch8pd+A1NxMQH9RmuE80vycqGLKnjFadlsp1p0dxCO3
alsH2ovTahwhrHvV7hJ3IqBBlZ9ABKcOEbVbc4/UbqhMibiBIPzGHMZeOXjx8vowROudipfuuWnl
/bAxC4fp1Lk43IZ/8+0FKibl3Lnbw0xl5R//dnkgojMt6p61WNm1N/UGfkrUFGXqT9Dswc4fKtK0
bg8PFRXTu04zkiU5RKntRGdGVh5jaFxze8jgfkN/u6A7RvW5PrXZzR0bMhV17ehbfg4+XbOtzYkO
8BUqIJ764b28IQYAvETMefNMdrWe+ep4N+xTF1w5ODlvfoDnOl1uQytTWlBrVCsiJF8nHwmiZbLV
jtKA9uf5gwXn0XH7+aw+lkkp+QOgGambBdG+/veSTMQyGHsSGLqxWESkUZcKoSSCy6m92ezKqxkR
2855jItoRah8Gswpigu9yv4cyGMQsQRAhGgMxzuy6Q6hJbtO0rCLjqnkg4aS+dHT4oPE7FRgVOoh
HEIdYb40ScK1ea8MbGtG1C3gNF71aruzWWdrYgx7B5mWSzWUwyMuQTBlvCeSbM4OdfScqwtUYRMd
UhabMUovbdYmrSn2XHGuIHM65eVxEN4nxNd3SZ0ifvuMwJJ4xgZGTGSg1IFzbUA8dEPXtDBoJp2r
XnMZlOT1aihZmDD9LEBAk92u1SJpQqcRnH92qBFjbqsnKbv4eZwzpsjqjyOhmDmP2pRZSjaOb3pW
Ng7koFn4XBu6a4+NLVQaCMH6Nbm0Bppvnn8qVGijrivSzd2nENdacyKo66dJL3J5yzuF+yp8mYf4
ps8l84cwgLaoXPFGa1Ji91eME1B6NaQmPCckSxoiXUpcVg/f5ggzIrHQ0utZCnIvZCUR7qPsu3Rp
n9Us0/dTSJaQ0AH5tK8OS6n9fZBZ3+SEX4GPoEtfneMV0cRbobc+NkOuYiVxPxoXzJn+m5DUurDj
FUoaDqNbeRqFjLis+FMCo919oIC08N9xpdjbtWYXQGMJtvI1hQYd9/iHF6HqGr24UHhuMf3Xv+OE
7EhXG3YcRUZjc2HIRyr2L1CP8CBijYKzuyiCKknakzSJH+8G7rLJNaQQbUjCwl40sQiyJ3TdgapW
UmkED2+m36ZuDik53zXM58BvHhEI3KdXyDsGCvp+Ce3ndZ6Fy4z/NgDLCbhDbgTzYxeUkt4GTCTh
+58gJP755Rgjd1i0tVDejWIQCPi9T6y5SU5bTwI8NI1SMzbxhUfpFRv/xX7MDUoHYlcTEfdWFobI
uea/TucxuGeH39PL7YI+zN4Y0g+w8GoYKDfnzf2J7Qgh60jXAVT6iE0avMsxeoLFFM12yv7BJ836
ZNDaBPafbd0hkePQzB3nYFFRTNiZZKQLit8UjlQnJ38dAI6EfpXlhjpjqAB3KzdByMcnOUnF1fdQ
JuENhv4GmtUlS68I+/IESVQnxGuShsydGvv/LKAPgcdeXmHFZcta1tToRJSuPJVGTexVHdgbpKDd
9/YqbHZ8UodGLJ5h7538uv4Cb6FuB8woLRd88t0pPCpYjEfBtnqJAU/S9SxP3SX1WiWcE31bB05Y
w5JI0toH2eoywc3dIQhH3SPKdJCozTJ7J/kXOy8vX7j2/Sn4HSG/4q9W//acI0oV5xLaslQ+PTFQ
gEh22WLOTjvpfuR2lf46KFgwI7v5l6jA9T9QlSd+J4ZaA46FWSWrwbZ36elWEcAkOrpm6CBglrgq
AqydI0yG7SKebPCtTLCkDRdXE0N8QyZNrWnlhvH7AbjAcwyTmOIQTwWlVCjFq22OW/Q6Vc3lFlIz
TPFpCXgYBJznt8eOqwXpTT1qZaCTru3Fwby1N8+NAASry5oZwDiuJnrtgfiyR8Y6tWotSlB7+s/I
13bV5c8xdvRetNKReu9cvy5Y08oglHACbWQDIbgfvKr56ObpwDuRlEn5hSQaK41RDlwcBcWi77Yp
FWVOMjOxRZHtDRFZM/3ASLV5cK3kIahem9dCBCe9sze0+1YMCVANsGJA/Pc7nKUoYjH/KnEhkh3t
b8UZTVdBAPhOQRdqrIYqbEYk/UXga9hpbDNXPaD9FduCQjwdyGAtbTc8jj5AZazGlYwSyQ3l3C+H
KApF5IDO/WM/SYznUXU7heKFBjKDCHEY0fOntctujextV1sjQcUbkKPDv8FisrwhKy1A4oTOotNY
52U8ekVMC8fZCteDV14xaS3/0jfQJBQ7A6ed/aSPOC2zEdua4CWFbyKHHv1Jmg7qTy9mp8TClm3a
pX7PtkR8SfUXkx6RoB0Vli2bKVmDrFo+bXctVspniK+1BEOzhCgl98y2wMfxJzsXRN4A2uEaPw0h
FzADUa+Y5T3x8sNgq6yBUiv74S9wBPSBYIwqFbrnpUBY1jSLXRCTBYajpcbMk1+rFx6ssgbZrepJ
1zmuCU8ed0nTaaCPGddffs82ljZ8AYlwnse1JtJrrwUxQPXpsd8F1uAlOSXpcnFi62Eyr7ZJdIvj
cHfIPIWmWEzNNfVrOql9YFXSQd4UaowTvvajuSft+hzBpWb6oe7sPRZQz0m0iwq/3Sfms3GE0HCw
m4dnFPbmBE6CIrDo3Vta9OK6qW3aJ1FHMKkTSqz/odA5t3VrmO/bMYX3m+79/xuWmPqQ59ixgxpW
ZkrHxjgmfz11c74bo8sSWNlSfTGhV0HBEFZDN0VAuyQEQL2TCd6KDWdUSY2t6NeR7U37GleWU1yY
9UW5Hwx8zXFp2GGOtOGoCuDMPHc8SRnznEmZHGwGFc4gY6NAd0dTbnu2D0Rxdox/l6XDEZTrQKCq
L9hyBUUV/XaECnTzBVAP90GlY5cJQP5Bu9HGU3Kyb8EGyvcF7qjfds6HTKbeLlDRq7XR+WGyr760
MjAVZtykRDQaPFVan0xh6k1Ys0u3KLl1NrGDTwFy8TrDJkqXgZGDEpyd/sWrldn0X18MoTQs8wO5
NIJHXNxW2K65SxsL0D1qx2PAibxuAOwcsr2NbKhqZ4DVDk1+kZYJai/Q7sHuu4BdP8VyyfGk8H8S
kLSRTC2vhJaKksHz6WOi8xH9yJYunqNIljq6t1pO+QV6Ia1R+ODTkyklk5jkm46ck+Cpwsqo5v5i
fCokyOFgWDXPGLsYBX6PJ+haYI5iYlTI/prvRb9RwzPHdCi/LeXifQIVB4tIU2mEdIi5WGDvUpdf
eCpPTlY26EFXGUhIYE2ZHUAo/TzetTpEkXykrN3hRpsSmUNV5SfMNTkyRW8=
`protect end_protected
