`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
l5kxVQHg3bYJL88bXYQFJlQjk7kH3h5rGItYbhTKcXRQsdxiB3c52a0/5Iwbc2QuYFOaDTt8YbIU
RE10J8E0u7ez/ZzoNXvXKxx8ggqRMs8QyEj1NNFeAMoY5/mcfgdZ52mz55uQ3RpE5GSYkjF6u1tm
xGzdkljDivGlq2sqDpoV9+15TKS1QE7YQf0v1DvUtP7S5HXRJXFvGbhTW6NNfwPPRDHZbLtnSIYZ
elG+42+Nl2186ScS1IwxqZ/86NlRTJiXCLoSJyjx8wnDnuJERxodWvoOnK1NNU7eV3ubZ4GfUyGe
Lc7uaW+2Bo3dOSXjbnQjxHWAxpf+rXjHDZLJrQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="mimOHq2mvicWh4a2EkTLKtDN8IvHSZb2mDbu5Qqgg7E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9104)
`protect data_block
TCunvpoaiCevMLa7IgQ2Nsg+4mwFoMcV30J04Bw12OcVf8jgXSEId8tnSyEpf+IEJ3vF8pav7z86
CDGsU1LL2qvaXTHTvnZf53WSC/EEvg2WfWXRxsBjUYP715tToTJOPq7SGnXBNZxw4o4HJsHZrcOY
vfDE4OQD1DW4DYUFSRy8Pdfi5QMenhjK2yujdpVhd/wrX0X4mWoIFDB7S19bXj5yRxg1vmn4pjLx
iog/Zl3cFMk/8dC60zAk+xx6Tk4Jh/dZpHhKPsqS2h2t7267o3JESQ/zvxLL7UofGSSZavk9Wr+G
7bt2dflLAJsWLg+WFOJGG3KNCPujU81CMpXj5Cw/lcpktAY6/77bVyxKLKiKjo3OGX3uzHCkyQkf
uAR0jaBXnyQC3ckhb6cboMMpKUokL9ZHwflfsWmuhfACAx43p9VPrsG1OisSkkvx5mSdgnzuVRd2
aKWzE8QoTFVFqb91EubH3dFB04eU8/77LmPrzmSxBYlc4bZHdOzB38wFm8fx6upefYOPgPO8ipzX
GATnRb6uSPD/Gu1F7KgeZf3ZFUq+G0Majte6DFeZrGc6OMs35Xx5+le2q5N6dLdVcZNEoAUuxl56
GpZrTx8HD1z7FqHXulM4jIbVIw10jdyDTZA0sWbiOV8b7bSkWVeTHOcgKKOQwm2HRAcJB6rj533y
lpD4aE7S9Q3hxluXKhotpZ54D5EXT/LS6hhDVfs9CN2MUgmzRPeB0mt34pwxOp52l6JMb6dntoSs
YKh/Ko5RV7QLxVufwJRhYyPAV22kzwWxxUzbma16TRwfgjK2VCWFawOt+3AQ8GCozEqEX7y2y7gg
ypMZOFquAz6ykuPkOrTf9XnynRPWHSw+3fyrxrLZvcJFZRHOd1mIIY5t1lo3ZpeqipJcqRnEYNT8
pvjCUM8biibMzinfpJqatwczB5s69IQbt9sncbM86vqQANghd4HdgGF59uIT8fsdmAHHUBGLisYI
kQVIlQqq34p/2dNJeum6WBLgwtel3YK7APlhKhLRpryUW+brK++E06PdOvJ7WqXvbsf4lRubP0E2
IZfFEQkV0fC9bki11qg9CDY9vcGX5HbADGMOB/d114g13yg47ILmfOKwc6YhLbDJ5/Sx/8o23lZh
vfsHYsCd0XWBTgzlYW1RXK/hiORPfqTW5pBhOuC3Q7Jr1/ML8aTdN1vW3s1MTRuozYB15hwzW43q
fHKI2OjPqEt/8sPpttiTJ6JglBGQHPIbXWg7dtnKzbd7MFpLgYVQqidarh0TdQ0oKcAGBIsh+h37
jmGseunvp5cvjZ+3pXlUFdnd858D7ICU2Fl4LBIAabaXSRXvRKog+hbnS2FzAYwXk2UKxMmIWSuS
9PF3ZjPOrTM9MqhVeNJouq0DTG91ZaZjQ/1tiQGpx6QGpkjcDP7DCpAST+gaRo2ei+z74gmFAA/p
xIh0MMtc5bFCVEWABZk4/LlHGVkZ8RuzRS38qz/+dHl+zcINibfE9j3PZMirha54EZx+FQGBoJl5
q4hqimohya9xGa/qVYzz64NoBWR14PGD+q7QZh2BydJ4JChCUXyPm9qwYqxquKvOr8740rEHPWh6
9Zn/3+ObZQE4qndDWTl80f7ehyVIvdmO3V51jHIUBSdaKobNY/bq3r1VN2j10rPT0rIpy86qjwhv
OxwHEU5gy1CA0NONwQcPULlqp2pI6I+MvD26gB18tLW6aw21+JNNsIRGFcfn0r5aEsY2Qh+exQIx
5APoVgAR6pkXH54z3NDS3d7hH2jXl4cDB6yKVA6xSpg0RqsthLjmZF9PmuQSzNBOkWB8hNPe0NZh
9sP4FWdQQRWukJCVAGbrq5QjPx5mrAJmL4OSQNjNd4kt2POAEkFGFUtJihWJY9ZlQTMgj20bxb6K
RPOMsAxAfJceU/fWRI/OCHykRdRFo760An+Ms2jtzO0IN7CMOm+i7gBGoxBk7UScgaXTW9iy5buS
EbTaZAZbX9KszXNN0viLVQxxkbQK0P3aeF2VZAQIQcha73D3jacoC72HmkBO+qtkVQGcoJ1ISStV
DkJ+UAxiXUCoN16XLCYK938dJxgXk/52iXCsxhhqq4H2uVZ0xWKn0FArqQFDd2QAMe2Nb1l6h7W8
YVUnUy8cZUnRLw7Occ5lZ632BgwnoNvwdyAeFonNEKjZq+QA+ZlBH/b3JklN0JY9/27DkncvmKPA
c0Hl0yes1311pd2EcUoY+BWRgLGYCnsjfKkt7mfNZ3uQw1hUuBFA8g8Sv5c2YaL3O75bq9alvbc/
w8m3LwDcK5Ufap5U3LcdCEI8S9O1RdzVe1bPeRRB0aoiMVlOSublrxoTBuVbL0ZlzIPMEwLXherM
ptwAMZM+dNvmo+5lrn7I5h4ToDLB/I2qpHouPN9tumIj83c1M8TPTBz4QvcFmANPx3Yz9IurEm1A
XDf9WO+PkfNSSN/365R8akO05/LtxpgQAMykpv+pc2kqYf6n5e6pDSJZDAiglrbwbn1K3x9qdU24
o9bVNPElV7qB+Rs3TmtZ23Jz+SCgkm75cvLXvkoLWVtYy/KWDYLrthsoYiCZgT3BekIou+oGnk7j
inoWgUuRU/glgohGCUcNn/MpVtEbJsA29/MefdEVglvl9mpuBsAwth4ObHgbLz3nN/oY0KKeDaO4
XBdnJSHGysruQ2STrf75Iuj6qI/mBOIc2/ixTNyxWqFrhkAXr8qqqz03qmpaS2wXCqbzj5nqJ4XX
KJrKStqCQ44LNTe97aQSvasjny6gCSborZEnMYINaypeOjsq+xyVJMrt7CUTxqoUc95nj1Hml1OY
PPdc0Os4MnmzXTgSGfl94ra5rqr8ZmOtf/XqTn8O9Fkv2FXMICRDgJacWGmGc9xaZuIswYtAeZEO
sT96mGM294UCh2y7iQBL6vWY2Nfp/xiUJZRR1kksX8NwmNnXKC+mLxan/3Z+gQocFN//CIDtERry
nwfnOSyc5v7yd/3lubGLfxc0Ze1OPA79ePEaDkED7xATVfjDB9wLn6tNEjAIZl3w/GPdjg0CM9wz
k7yj1HzT8HzT+1yiGR8vjSbUWwTiZgBPa24sM8tBYxz50kqoinUgMjQqkCIxfQ5PGFJ+xYItFOCN
YSHwWIjs0xgAD12H6z400vtWoCUUn7PqZGFtS4VJCa1vJNZudhjkEw5EvN20SHqoclFI6pXYure+
6de4UPaF+eB7XXn+YfKgTO86SnMKlPbNwWHNcsXitoRlaJwI9vg2yTmlNk+1Q61r2Kljdrwk9hs3
8ePzHc7CA1fC5m3ULa6GrN3q8C/jzKDE0BrfiU6GvX8FAbRA29pWIvh87pUwb2TguqKCdTor9zSb
RtInF/CXozvkOjFS6qugy6lXAWnYeLPGTHal49qewi4Ac7mlIkIHsCbafxjRuOIl3rLTAZm9ZvS1
o1hHCMq4jhktuJDm1eLkSOiWaAGEGRltxPcpEMg8Izs04rQiJdfHScX2GsLFkoHq7qbtpGYgu5bN
dcjU1gUDMZ0amhNYjTV5GYY86Ja3tIGhZCs+GtUpctHJKUcgVNAYDg+4vB3Suo2uJlkZENNmAUx3
6cl2pfOpch+f9fuwJywV52Xtnk5/HD8kZLfcsva6pbXCuD76Rqyas8h04dTMOMeVFntXLj6rT3MH
0KTBGoFvhQu9Ox1BNqG9EZaM4YPN/JnJCs4+KO+f1XY3PIRI8s99dTDE7PWOJ64T4j1LC5QpcxZx
rtTdS1L7y2/AVKHa4591LJSzBCLp/keyiG4bTIlPoCT2qzkbZ6zBvYHVil+z1N8X08JxwB0iLfit
czT/RfwHMdJ5MP0oznsuhlAx75TWPMjumyQ7rBxZ+CKNY3hUsKvOGcC+EMLIVYLBP1Ev8RIniDX3
IQRHDJ4IQNOwVfa8uvTgfysnsEb/cWCof8uyiwuUoZd6QkQL1S54m/EHDdxsdsR0GGZlsL+SVQPf
wyCAdTgMa4VRy+sw3Oo/vzCnck+eQsj94Vfk1p37sAh5lOzYFaTw0Yd2qqjKnO589ZZYqsDhmcWV
jHPUlU5vvFEXPY+LZequoC4t1ycswx2lmj1tkyFlA9xWDhdd6BGeM+Wvz+iPOVnurqLJejRxwf2i
cSSxz5QL1WyWwq61WVxmLuSj79jh+DMXw4L+hisJqr55eemP3Ufdm3ui9A42fumyQxnlUBAIzcS1
UBvWsW9gN4zytHH/qtOhCEbE0PkmC66r8u+TnJ5cf03j5IbMkcyFQ/rH7xrqpfBgFtzy0z88fyFH
NjrfUn+KrSiP4ju0NTHhodxipYfpxTQOf2lFB47ZZvtvpoxjiaSPXSz9VtUAX/EeCQrWtmW+egEj
QgakkasrVW5CbpcwEToMp3xOKt6GelU1W3qds4jssaH37C41voU2CSi4vCJ17yVM+CC23SpPZQA+
9WEZH0p8iVgGuBNvCQPgtdw2XO8QlPNVH8UbawPfusC0Rbv/TH4qw6g0fVLw1sDGEmvS9XeWInGa
UbSgjbYg275GPaFx8XEygs7cZ/rxOLvdd5Vfbxt/A5eyCtmzMXXmFOdzO0xouMaHY2T5pDKEx0BX
oVbeVOyY21Pk8DdXRgyyqiGau+vxvgwP0PjNDKxp2xGlwB0Vb8IWgYa2jPKjuBIn6ohxT4+ptCEO
yosStvFRlaZKBSdZ4UrSt2Ljq/IEZzOvUxmPhkzRnNUljJwGv9qClS6um1gV6BfQ4ixEqq0YMOzJ
c6cxpabeK+f5ieehiJBzjiA9I6AiEi7GqV9Sz8ZRsOKnQmRup4YRwYXx1yIn0uTEBM0kk8wmuCQp
uLsAyGH5wMSxMxRTIFO9RmD44WX+n2leSOs+TobWJhQ/QSggCShqiHOprgmc+tUgbp+zA3NBCLnU
m75wYux5qD8Ipq+Wr+Hjt4lq3VRTAIYVrPJUWqA/t/vbbA6Arc9C5ay5kX731IIwLWqcknQHmNbj
SOY8BEKhu5G17ot0QxKRXwcqbRmrCEnbC77e5+A/8P2R6ikuyBo79ZyPkAMcbVOJRWYW4CcLIv0G
UlahJbxKXHo9G1tq0LxZQ8oBkXRCMPB86DNmbPkUNHf3udMJS6V4Qyo/L0IigZCwGnj8cxm3ld4o
oYimNRlYaRKeprq005ja5RWMY/MDtpz6BThkKR8mAxg7Gk/PeNtnE9BBUcHopoD+wbDmylsC+fCQ
EZ1iuqEKeMgkJ22/iDn8Pki5sL1v1q3Yfmw+LPSLwRMdh0UFyygvDlY73m6Z77v0DAI3eZEffcq5
Ma776oo0Vh7fLWz2ThigRKhQGRDntj6wAtRvKrdwQRb4CTswMMIWJA31fKxi+VtONjVChs8RoEuZ
en8vsX90MrQgVQrlAIort0tGk+5hhjWCU6yyy7lPnO5Z4d5pHTXDcKRnJDpH+EeGhs+h3A4s8Mrm
MMJtPH/Ob3AwubADC06VAZb6JsoTmMO3bFBFywW1dchL0em03ZzxWxro63RYoy8be+KygYbxhlv5
z+UouboGRiMuyLEaTmyXiJIdrRs1lOlVSbUEve/7KvfQWshOiHBM62UfxpLvU3nxIqqZzCRF4rGB
a0Z1UOiZ9h6eyNWm/elUJgMg2n9fiotH1VUTsVSn+W3bcJBtHZiPVbvn1cpwmTfr2FbJ4lddiCY+
6YnhJd211cN7P8dCimLs0be0kOjqXs/fxFPEA+kyHaQTIztNGGsAgHDfmYiPdFFE6l9A+TBRDwJa
EHwGnK6CYzJm+/OcQmLQpC6SYbZo/FV8v0LgxFdhezbPaoUU7vhyiEx7tNBf8TlElv5RsTU8V+vz
jbN+JqKmSsckkYHteHARJrPDiiEvK6kXyrKEX073j/CI8P55M3XSHPG5cS4SX5Z+8d1wjMo18vq3
gQ8uE8WRRK+qeuNk5jKzKqIuwjAlVHKA9Xc9NG9gabAV0RR9yWlLHHUcLvQiNWtvYzh23wdVr5sE
au2TAiqi2mszVEDkfBovo7gd5u8FeSMCLc7TDY3Xbz3DKxkWiDPFSe+87ITX0mTNHb//aUud3xAe
zn7Nf8toIeTTIT/dUVVmu916W4EvHpUbbaIRrVDTMhkYtcrw+Mp12C1qBiGYGP29qT+oQCX4ds+d
r3I0OaGM+dL0C5/5/Cg+kNB1VOmNvBFyUecPT+qaEotrgFcx3oumd6qYa7GzN/2R7z3Tk1cVao5u
hVrv18as1ZLSnJwwDVch4WB5ClbdaiGSbOQoRYq1FiLLiGhk+9B+023xaotaqC6mxN1xD4bQA8fi
NSxzHl0gKK/dtCeD+h8Q3fSTqkiWWkI7OuRS/BtLD63xzPpo/PSicWbq0JVTKGmW6vAbvJHoScZX
tTOuRfQLXqyhd4hqeEE2Oc4ilKRvNxEGsVa9XCHNLTSDXQ8G/NWBl+uW0S6ZNTu7zTkb/+Z7Y4Gg
3Gvkc/r6e4lwAC5i+mL5bp+GUgjg9CmiSEVC1IlHwtL/S5DHhBng+oXy4cPiO8KC+QFED+E1RriR
e3U8r6QFjyqNUs2tKWNO+LR0T1tXxI+rb3taKpVLS5ivSX+AvfaI9YUtFXX7E7ACeTxbWRLJaI++
X4FcFea4Yd+43EWl1krKTt2aA75PvNvTf8/ItXIjg6MQDt7U88QsmP1YqBB41LCDWAYBiZ+s0MSd
a/+Czp+bqSSyC4pJHljnDI8SHLf+/YJa+Ie2tnm735OagALsHVWSoPCKAu7xoudvGTrAdqf8SjcD
M2Ei9UPl/3i3g48pzu13DqcxOzMfi3z0tVAaP5w+ri3XnssH/x/CLJO34F0eId2zTqYsJubo2STn
ZZE4kilxjR8j2XPqjxbsEgUN5kQXSGE2GAgtVrFSu29XgALpbnODnrqTGx2WDGUMy/0runs00SZd
HlNx4xRvnnnwker5Tc7q5Md3vBCnYprAFRRxZDJA3V21Sy77iCfAc2ZKpGPYrXulEY4Jv+qaipLV
jYoK+6dCusPVIaOkrC3E+ePA7LMPAcqibj5rMWkHpxR48ZifCUAn+2cqbZdPU+YfJobToeV3q7us
YUR81nM8rqnTjRR3A10bDj1EEBaD11xhkk/upJpPF+m1hm1JCPRTVOd6tEVGZ12ptgczhuwzAfXe
lrgqeOc24XY50HHDPm5u4P/gYgpKm3kNdau5c/+Bds2OpBL7brLwsiXtt7xXETOuAmo7Hd7jCpDj
0WeqjUk3ssux+hM7srTzznTASgUmbBwPnz1aWJbLROxNeAiftEbd9/mXqV/yhahkdxqi9VPGbjzt
kkFPISfqXmlUkEwgi+8ShyDZoxH+DuwIs5Evuh9RbI+EM+3LezyQY1+cXMx1bgsbzxdNa55vxmi4
vTLKpodylslLfm0BEsVFIwohesSk2M9/t7cjEYKvHalMQr2nHoiUOJZPRyIY2jARRcdmSY81yRQf
L1QXc/xhl9vKOWTVjFcribfr9T5bCMXPEFNWVM7EoN7Jkh1u1N+UgEPD8ZZol7M+nkda8pxiCx0S
4UrGYbxqGW/dDmxj0zHi8GM78dN5qcpmPjdO2yBjL4K2u3ylJqhbqB5Vvd4i8Yrcy/FTHn4B5X4C
UpGfOjWQRy61jGMGzgNEpEWfwGJCUIofYzh+SJxhWhV1TP/r19serdBqx2nLislNZcSWO5aiqaPq
ycU6fJvwxUidlLeqeBzD2DlkjTNotY0CbYEcRALHNrgGgJULOe1EX6Ie4y5R6ZSZyOpdHWESojxs
H6fLpmCHffnfr8E11dairjSP1RX/XqnF8AsSXY9wC5dmZACcX++HoxOhIHyj4AGljmgYri6T0v8c
2dGlEd/CR5a1arybdBpN0LOnNoffkPX428L54hDjx74r68RBvJ9uFRJ1JWVjwClhRqxSyXU5vvzE
QheLbwDpB3bkSsjrw2PPMic3ecCBx34xjxZGtjTV1PLh02hBotSFUFWHFQXzIWS8vq5EP6d+o9/c
6YEinbkmBbHG850fNm0YpvQVk+CSuKFs9f9pfHJ7Ij/o1lK91XoGtODCdUq9t6pNKEFs26gL/67G
HRKjbKqPUNoQ03q67u2joY9D2jMWpNSk+sSYhwCL2OKOMezjnYIkXEhGV+bF0EeknLm/wlLBWBkx
AMnMd7P08mewRPgTfzIM4AaMvIVwQVRnEkAbqXmG/L2BSiv1uvythLbqgEiA4LhQoZy7M6JfJ685
lY5vmjZDf9A3n4mUytuvfPjlVBt11eLIPhgalAlhz0P0/vUJ6bLFsSkSnUpr/o1u6q2Mp6rtczPC
WnnRLsHRjoVvHITviwiosd5no2O6gSf8XzDLNqPSyNdp8Kv7KRD91LPGUiu9t708JH8yrBeJrLWZ
NAvRNPGsTLjqO2qlnEjNIudg0U6g15vNTxZNLP3xmwKM6lOEIf5/kqC/EYcIL1LVTAdcT8rCMBTL
W11Z7Tb/c6xuNzQzTZZULtq7j67Awnek83Vv2RQ0ENvA1n5ITEp+TOeCOc0h888/fe4qKnY+trXW
CXiPmOau68+lFD9hSIVHweZJl9/Xwb0rwOlkvTnRAFtr6Ttv6PWkcc/ydyf56QoOVyiY7jQE1+CV
O8WSNGE3gCZIAd1V0Z4SFLu3wG99IplvY5GxtJEQfMJy5uBbrRSA0ThEGJeYW9Oz383+2TkWkTqz
yXzlN36EuOgLo+yZ+LX8/+2WBbjFLN9/cfsn+EdpHodk86qca7nj7hCT4Rq7jCTvqk8OeEcm4TTT
NSp4HwujdNCiKqClOLZPSbkYhr9UVjjVmuCdeU/WfyHbsomokSzhoLFSn86YV5YC9NnlEdu4ZFjC
7gu9mMhniCjlZ4AUKPMGZ0S34bZno7aP0EM1dmW1kib9KCcbHCSAvU7JqQBa8v2sPD01ZRS6dEoq
mtzjLq+qC1MGRVHLOPpyKqyt5HqzAKv2ZFjoXjkE2Y3NXo2nNcsQU66ypg+CNZtdkaE8HEH5v/tq
1pso3BlNChQvllopOlH3bJ3QwJ6TN0+QIgd8rlTIgRaXg4uF4Wyw3meJGBdtxifl/Eerh59n5o7a
1DOAcoxO9zWJlK7Cw0J8izmlB+ZeYTp5dx3uSmJMsKMbZ5FuKv7HsAvA7X1Jhk0PAhpB6MtDVhif
Nl+L+imiV3+/gX3UCom3R1Psa97r07yNckxIhyOuVJIJZJDjWDUFHIRt2Wiz/T9SjevFHXS5IPJe
biGVgYnAeYm6STnbDa3o2L5VfXTW/XfZWgYyqjsK39/1KUnlncTxVPCoq8mYTmQSazFDlGGvRNc0
IJvt2nA++pw60NFKyaVQmie0Y+CvW9GW+54bPJj27hTgiOrHftLlR/CWvNC0M1EaGgyEDrjDbt3v
PVHyoBGth8aoh/n+ud3cIoAB40GNYfhn+4TxHA7nta8QQvr21KED2bLwtxdqKc5G8Ur4nT83Md6L
IPfXXcr+X1ZSfvq3kONSzZwylABFpjqmZi79nPn3Bt/ax3UzMbh9ZehPVsO2ZEUhtCtV49cK/gFM
+zqnN8c7nL5A9N8GW+gBevjG0QGcU+7OQFeg3iCDzySNjPuxw8kTDHhbnSFNvlw0YrA4CVl2jyfE
X0IUNJvW4xpw+O3MU4ZRsxeEsh3UyS9UbT89H0pmXi836/jlubCb5ubxwbBG9GVsmiCGhkDAfBaJ
57CTTmzbEtnq18i35f1zxMtOsSud2chvJjXtTymVW+i/d5rySSlhRgHnVAhTxW8Ex+bizrUBoEtF
DuLFpYxTLbRA0abhsKTHkWaBHmZyDOROntooL92gOgoCLRWqmWtvgyhVEc4+UzTVujOYLb8f8Qjn
bDcCerZ3QmzMvg2YLvMGxri9wJhAB5WTvSCDB5PTsCWGLk+JjLEP9hPJS+La+LEGLnedj2pVR/zt
qbP590qKWSl9y0AzguEYXO7NKQer5DiSHBHANuFRyMJcFVAWyS42waFEodOiugBt1iR2vfTgGWpo
BL54q7CiEp29o8aXpC3snaQqF2jpdMAP0aFYyIMSnxhUPxgPoBLwOvuGmiGb/a286DosCLxAoCUy
m2y7s4t5oLEZqz+o0fT9ExZ7qavcO8BiIGEyBMAKI+7Quq0GHUkxn0hk2DyH/5nOgU7Ld/uVIZtl
1mnG4Y2+z9dozNhOypZ6WJ1G1Vuir/Xq5Dqo1iPuv4sJ2N41wFBqyAZP+BfNgzD6Oi+nPmERazIb
N/s6OljlrQh3YwzQ2f5W5+pjIYZcRSpKH7/Rn0gWEYgAKiiqqZ3Xg31h7d+sd6SD0UUkjMFyvQTc
zNPCD3+4G1a/CVu4VsLPFYOboYBmla8Yq4grx/wOJgguHaozfmORhvyTcb7ea6OtlQDyRb+otWWX
IKcfHh0K3VJ4nsaF6sYGGiTdB5Nmv3o2NZE4dr8Qp3hldZyoUboXD9nW+QXlpdJCa/U4QzSZxErO
jkDJCrl7e8J4qRtuz35ug0XQ8hWbC+q+AqnvnEJ1lDrQbnVmhz5wCRux6ucUmQbS1tpYEIxjIOw7
yAIc2nO8GBkHvvVOcdO0FB4mKga9QsuKI0hAg0kwdpBwZvL7PX7HInvBmxZaz5qpDWdNBZbr7sz4
7ZVVehEYGPL0iU9rfjCCf0i4ljxjlbcrWM3cuvGH2IVU4wv04SaPWeQQVUWmaXMB1i/f5bVV8/iY
DrZFtE9IBvX6AqYcn3kd7sDEPS26abYUXnDebkJ9yYozfry+uPlFOcfPHVG/ihA2VL0HlRk4Aj59
CjTISUzyXOaag6UmCnvEBUYopouXx1wJk2GPd5inK2Z7PZ387OKYs1XCAnFEDSvm/3w3n1fRZ4kZ
GReF57F6YyxaIsIYx4irvvE853KmGm3EhdeZs2AiPGd4n6Bfo+RaMBeLNKke9dd4jvzq0NiavSvh
1R6waYy2Z+IPXt8yXCCUeyxxnGIgSdhSVC8MGOmtGhcBgxALOxt+Et1QmWRElNNGf4ZdjpP4r632
7PITHIQ520dKFiLBqZaCO0mdT3ciSW/nr/YaO//KgljRJU+f2nHad2LCbz0KoN0TXM2y9vOOKZwH
Cx7ble78/xuuiETM8FnUdeORcBtL+5W4Uq4PGUWeQnjB1wys0Cf3+Goh5xS2GXSwhQ0IBriHSm0H
+EfVn71HEwv3r4k6fqOcfW8cNyiMogRhs45z8dOSGt4kQr/hrfk24LqDGs1K4VCMQlKJHT6DuXDa
LbXZSdI0R2aDVQ7TAUFLxd71uaKFGAenVeS+B29KZTKCzYspAk4W+69UFlhUHtn10Qu9XLG7XqR6
mDqchQUa7LOBhd/kyEd0iIcxN90mcNgFgUiGwltUmqmY6zU0srKFJ8FPH6Z8RjMM/0+4meCRk98r
0gi/uqU+PK197S2YpxX+5IA4lKVCslzy8MS4izP0LGX7sXmCAsesDVQxhABEmoAvLDUnhwmpzg1l
CsRkf3UB0N5gCuZJdVfKRZ8MlniuW60PqHdMWbNM8IYdgzCg0m8EL0ZkvwwBEX6fjAM64/CG0k9u
TRVWJRljvtPxAGvaQjNZZhwHlr87F/qDwtvuFIbnAcuRr9gOMPm+gonKg0NjubsNVmpOQTuwua97
vchV8BtHiguHsAgFVTmgBft7blmEf6+HRw2e7rFn73+nZKGNqruWAUPldMQNqh624v50FmeQJd6G
Vpo5NHcteiYJVobeRe3z98nUAEQKhcI26P2SxlyuC2BoSqlZNhMuxpNIs07gcHXI8xR7Xyw9Rijl
nbChbkNOH8K0y+smxyfCrGjQHRhACiAkBErhygAsmPti4kkLK6QFqJEYV2B3GT2ACtaT9K+Amf0p
w6Eu7AaeQJ8DSF4p6IJ0VFV10/1pDuk1jblip34LiomEYQ1D+uxBMmd/mQuUysi/ldN/VZ8LXpQT
a20GoCfwW/XFk79nmS42gSIc2En5GRh6EUW1HudBnTQGfA4ty53WLST2QJbqXWlBAloKUe53na42
+xdSwoCqJoHsaR36eQd7V6dftWtm1qstzlRG1t4krh8sTxygU7jpFuRGCsKdtcwLS0TOG6h79B/f
MEdV5pP+LZphR7om1Ybqq657OuqicPG5uRrkHtPMn1TqhFEDTffOPRxsl086DPrg3FLzeTYDbERl
zydADyrCZiNk8VVaXDhnTyv1a3PiaHv4tjmQv1a4tC29DgOU2HHgkwZzClvensKSoBhuMp7J532R
qRM0obE0rSp6Oih5jOY6efKdkqmfKNqBJlAwD08KzyN9jFMvd327OeE=
`protect end_protected
