`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
XaWKJhoeEYCuQe2H4A0E7yqZd+sogr8YhtrT2qXnKMyHKK0U0ubToey1fJGHw7P+9lKnhIfZTyw/
czrZZ6SGfZKsXlrAxiz310EKaXvWMGKYK8J3CrkULT/MrqkRUDXmy0Zaanki4VRWXJQQp+nnFcqs
wTqTCaBwTFbzhCi+rF8vx0mLvxNpOiH/TfTqtF+1aK4cdS1toOwDk6Hmo6x1vv2hnPfXp0QB7ugY
BSBPtM7XV7aaswq9yVTPiVOkG6oo7tcm3CY2lU+m2ng2osGjo3YFvMS/B6TpOA3tynSuZLXmVgoE
kPLx7taE+V4RqNhzQBEkVKVToYFfLXIzi6j5iA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ZfYE42WY/Dl560FM210lJTk+uIjrRqhAcCmUHVtd5Aw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9872)
`protect data_block
DNwmgsOqwR62PFZn6YmmkGHGTrMd230O1Hsf35UTgqXDhaKX/e7WWeWwLAdrLLwer4ijAMbCgAzN
7+Kl7Zx36gBhvGnnUHbDF7C13VAeeo130p4mb7Y6ismnxTeZekjB5SZxfQ/TIrt4CjSnwwdDftUQ
I5x6WzwV9mkye+hi7zi6Zb5Zxvdl0XiQ1ezXz9H1nvzBIaBwnA3UwKkcx3UowQZaY/xlEethtmLr
U8oQsB1JrLIL1JSigF+msA0ROYV6M+jrppp6vQ+BEvoSKt/Tlt0x0IWlMl2SLQN8Gn8phhcL7ObH
Nk25vFpVort/2Fn0UTK9ok4l3EWvnFoS6vvgjPdqEmnIZ8ZdSQ85X+srrGBAnWqcyp+k0kM8D9bw
YldIKLutzsSmxvvpdA5KsbhiYvqrGDDKLP8so6w7SvXJ+X8rX/jeUMOqth+hpdeiNhTUuAPPVtZT
5JXBNdd6tH/MTzzChIelCOBylGLBWhZiQ/CkoH/9TPubYa61DqOqErlah26AVsygTxEyIXi9n7en
ExTmkOve0/9k9wlCSeE4t7F59TcesJ/Wjfkm3VBHq8D50nLEDcbO6oEJieFag7iia7BUHP0ST3lQ
Z3mlEhrm1yk3So6yl9qVUdEYlDS0kOTUFHJS8F+45+R5FKBkrUIK45MtDWX31xO770a2+Psw4vq9
CzDqQqtpNMPHoqjEtA1Us+rrzp6H68SHs44z7uigvHr5Ho79+t5gS+wk2+YMc7pcHnVLDbyifyZF
XTA1C4WLIsxK8W0eSNf4De4qcjBn03jR0I8oBf3ek7Ujxr2GpyblARrY24V/GnQnObVnbUQlY7Iq
pHbxEVh/fRSbvQFhYcEutlPxVMJo5azD/RTL2z4L1bzGGFJTm6jWC5Kttmm3DBfh6V3PB96eOoYA
NbSiJMwJ9h7hJ6Ib7l41vJGhlg1nyyJpcnFH7Zu6w9rYWqKNm3JLgUDVMRJVJ36CPAM7BYeOKk4n
RJvuYgkbPtDYhFTWL5OUJqJPicDwZA/B7ycEwvsFOmbJfwL+sQ/fWdaRp/n0RNjIAJlEkwxzZZ+L
Z0OrP+6HFeceNo7OKfKP5PMrvReX4OcDVhibxlbgC+RTFUDNMNIS1kBZflUrlD2zbwC7K4fZtK+0
nLwsMBbwJhoSgh58mgqf36b4tKPHcChXxi4v9gz8StWK+ana4kRCDoIpowHQsDJgfqqRnAgYfvxT
s3ztC9KSmr9eLabEzqKU+cFtn2AgHofGaBJPrpxUV6XQfcxHS6WS11LUHoe7SPVH/fPJ2xoRJbHB
2cOcbrmiqAf6qkw/2LiKtP0Pz/G/KCut8ghK9f8YtQRseIe+OVrmpuhfcNFNxBLRxszmC6DNDTqM
lfk1mKr/b05fQFJPWSxcVb+hmU5li2NRpj2Bc4NzY3TgwL4bDss8sT8uoMTTO2UusoiloukOX26S
QTBka95mWWP96d36bKe2AyeFtFfzDbNzFhPeJbFGqflPU4IXiuWm6eOC6PV3RSMPr1j3srdhwIse
/NNZI7QH/4IptMLe10e1kNQEvve2gcQUDkh2vb7DtoKnjYPjObpXHY/IVQCb1NyTx1/t8IR33340
XmFLMRjslVvGdV6Yd61evTZjEPj8vi1GVb5ziFM/ZnEpsmVwh/2Js3Q9w0OmfSLwIjasjchaatkl
o9jUALYiGP6geLgd+l84uzrMHtTaYNVDsBqtM6GC3BbMeMFfoFq+N+0ybc8Sc7LMwtGZ0t404A6O
YiCe4iKtnWP+auedJmVLq6I0D+uHI8ExnM7xqqfL4vw12EGEqZh2WIpwVf/A/5gH3YvonNyJyWQR
smi20j2w/erBnmP14jL0aI5hNY/Yp3bFeK+phWEvy8xEtl4sRbXBUQDFgjiJV5BZGttJX8NeSJDF
8Zgt9MVn3N0pRMJUl7hopGUzct2zhrcmhDOHr+5oMEaxxXmMf04NnruDgi+ato8Sq6MEIc6IJEx6
9CPsYOadm6GskncyuRjY+OVc7L/qOCqS5Px4jxuEyW9MVQvP+kBCUoITHrMd7aIFUaOsLVTmfHMv
vd5sTQh2xrnW4sRld/wcdWXMqq5Z7ZOWrVfyR4ASsHcYG9by4G20iXi3p9ONRGmx4CTKp589osxo
5qc4+iFPr059O0l4zgSBtw5pdZVRzjEeaOLIFYa/Y2aZAE7w4Yx8INNq0d6MJXf3fTWJ4KDBCxkr
B8bFHdLYn9LuDNVPGs1HJLMqPkaNhpA/+z8cYhnjnITT1L/E2P03bETmN4M2zPMXFbvYhC95AlQS
p+37vTPznWG3JWHzECDoz4zeZI0+QwgnrEsPyDudDXOA2j4bns9mguPAKJvunJIR5KKFiTwGBmVB
jhY0QnVGnwdC/ZerzBJEsUtJik/18jj5XyEGJU6XbdTgGm2XO///XJV0B6Q0Dk0sN0zjybyZ1vof
SsrhNvf88QHcNaP1Oga0rd/kAvkMSbShzTaijwI89hpZaQHGyE20Hova9ycIXh3RTuD9IztxLEDB
2Oe+VRBsisayWZceno29gv2X3K9vm2EzkALWAnrl8rysZn0EhLxILRXq6iWQMODzIfOXj/5IPWHa
gFCyogzTKaWHBPqij6drzIfShqN0GbgQ5VUGc97/ifFV68DD4P33SJgtJIpEFv5KZAEY28bWOehX
yvI3CqYWQAbTp+BQhosBR+kB5rsvnpA9jFdzKqci+L0X9IU6YgGZJdOqBC1w0W2SaC7Eq3fU1JcK
V6Pv0t/ethmILQg+u+/2NtBeRZ+SODnOS7QW8SKl+u7/H0TsVt0pfenD0zF9B6T0sPLpnYZD0K3g
2CtxY40vx8n5cPW95qfpxMOjYjYeLwT7r7H2A1Moz0JbrDK6YiGy5YsHDe33QE4i7NMXIFA8bUl7
WoPBTy+potHklxW8Df1Zfr4hWx54Md0mucUBOp9N2wBc3KmRSn0KVu6Ryk+UHhbsFqnRQd6/z4yq
WqTQyxVscRj3eVxQpinh2JPmvs2O8NxPYTMMRJSM7wlf7Muqt2FUnfg/dfogKauBiZ4XTbiarLym
ap3ybg0udJR+3vJANxvi9GMUp18hcC8yKUhDFwrVITmiipcpBDa99qtMRXtdZNSSVAB4nkbAGdlx
0dWc3mRT2KjorHfOXJPAKUs7ABel95WZu1WFeUSenIN03dXk0g9FHz0VCX8Bbbtx+c9B/7x86G/x
h7nk0e66OEaevh6LkizJdkEITQytumxln5ef3fWIw401sC+td/wpBsNyhyExX1dx1SqjHH/VFipg
R/yAx5re+GlJFbDRPTWqtX9U2sCYyN6k9ilqgWM4b2pJJQp5b7BIlxiY+0VLmuyqLFo3mgUvI8pP
29nbTiDCeb8gFOatzp6e5OvqMP8Ce6F67V4l1VKpLEW6xkduoGR1X7k+FfCD17V/36B3vMQ9fdgB
7W/FB6asfNGVhJYw8ftbawMGJk0SwNcJcVfm/AN0TpEdZzNUYisStneCh4jxl+083oPklZ21VKI3
WXyuyKirsNWTlzgro6T2yL2spHbX/a1LGzbpop+kNwdag6iGnl/osn8I0nCDDIZFCoTxoJOFTGis
/TS4mYyG3dyQiVhkzj/0Ju53MGJr5p8k/jPYWpEigrKkPHTA2cgSqK64YsOpZk6pKwpdsWV5mbhB
HVtDwkat4Gk+FPzmsjSp2lHlKpWVge+CcV5vfO03nBzmG5WQFMc3VDj/lRb1s1F0s/DcXllzfgWy
G9p4OTEBTrNDHp2Wn7WRLiOBIibYRongF72WNLTGaq1OsT4weozMi61gP51XWwbwWP16g+ZIOpB6
lp4Z2WjWGs2wKFC1uIkfew1mBJachrivoZ3mhXSRTAyUWVwriwu0yHubS7YSAX9MAn/kWOmxojiD
rQtD+b/m7lSlq4VG15GKHR0AhkTfHxSYY5BwbxwjZENvpw41f7YgfQ5ZOemVNxB0eUapz5kH+rw3
Fg1lnjJKkgc0+0vPqfdPGyeKOrpe/2ePFAI1l4sVPdqMgIWNd/RxfOW0fzWXn+w5tKqavl1J/Gby
BvFwIGLvdSICaatCYUpqrlx5P2/YgYUDpP6ErdbY56ps4Ko3MxCKlntQtvi+iUcSrUtrJE83VFCY
A+ytyxshFWQI+wnFiolXNiXMkW9KR0L51jPuf3tDY3MhjSZ6fu53Sfs9KdxujkjtFHcoExm3rNdc
0uuBhRjrOKE43SZx2cIySCYd3z1QweXbvkU6LvBfaSjY8VlBQqokbdQPtczlCYv2pC2vF1i2Bkfb
qKIfQ7Y0SYRWULBwy6FNicP5wOdIC1obHSIULz3a6I1AS8q3Z2mH3p7gfiF5qpf01P7v8D9S9rRk
9WBy6ZaOOrDSYJKm7sQihStzT2IDrNrFef/wqWZYf1V3Y9zSrrL5vxCN6dmcR+Pm9pA9X3uAl456
AAzk0cOYDCDgzeBhQzIRdqi+qIA++r92cT6Fpi2aUjS7dBaOhtgIUnZaV4DnBZH2F21QMfCGUmRm
wc75yAyi4goWAEhrjo4dkqE5UT8VSl/b6tOtSEiV8PpHHan3tbHiA21er+o3YymlNJ86C6xqFJB9
QKUqWS2kxHzqx2rpPE7RqRKnLf14jwvKy915u94Q23WyVj2OoZJkslnnC9qid0cTG5avKHHSVvSM
zHOJp1lFGFOhqls9zWrgqCk/tOxIbPhTRpmkLvbxA5RmOXgCxuAQSqiVyxUMTu4avMhvY/UZx2Tx
YxPW7JuOjZSv2XDMtTFAC1v8/3VhBZUzQCXpl1kpJby9a/5p7ZLAea7RTTIiHOqglGQYIwLVikJP
0+0vHoRfTg05L1kAYH2ushBitYWktQJOcbUrCLcO/Og3WAcdLFlueDgb4qOf6qvdy0WYgCm8tsjb
eiLCHhWJvfxU9MgnlhKRR+U+1GzJ24pYxbAU3+JI4Cn0a9IYOccdw0YO90Bz2WkvdIdfHmhHREOD
7581EfsGzSU7J9yGM27IqlufDUCrWBUu13k1payT8VWSjROfbGDJa8z8Tz+M4M0gKnM6nAgWWrWi
mypCgcrOnh2J4iKdMV+3JnDYQDl6qAyl3bfYCTmC0mgv94C+eBHqmd+Bvsq/0p5BjgMKUl/f30ol
ZCun8idlpxe3C5qKWp0jlKHlQzA2xOqp6/cIvD3PCrkF2LLJ0dL+/iPfFZVfwxJ/vEZSVA62T/ad
d9w9SDVZxJX0W4sGF2YoTH6PJKtKi0R576VM1jU2LAO+5YgtM65+NAUtiV30PjNy/k3PKepD25zm
ZtxBc2Lkmzeju+xKSYOPM/+++V2tBL7yOyYrTrM2Hsd6GZH2XCzzbFiA5Ri1cW0WQh++dtPrCVZr
qpAm3ei+YkZeqn623W29/uh5i39weX5DdCOAcx3K2iEcJ+eYfbdUIWoXpgRqLwrftwJC7qlxgpCD
0uVXHLhpOmAITvULOiCW5UcL1svpfNXukgYmrMP04PpjxrqHQgopEjfBeMe+ZxmQpkRTEqlavwKt
croMlh3FNfX5dWZGe0Rs2vLB4YdFvc6GD4Fp5QD9q9NT3XkUZCZfIlkmFZccBs6aQs6QEuG10bK/
Tdg+ytlE6zf1M9sKRarumDApV6nE0qe8PcF9hdU8fCJQTiLl3XVM8iVdtwZunomoV9pOtjp1kcgj
CC3r/v+8U7/Zpn4HmpYEuOxlm/tFzCtf6ijo8RIUYd42M5safaMuFVqOHwF53O/aDinx0wiR00fj
4yYA9UdWRGoVuPYVHwbqKV7cZA/P2E0oLwJC1hjCwd2RiUkd8x4uliSEEHAAN9Y3DJ3T4Cwr4iyx
OmquHdzcMrJS5wE0U4M90zUeNBJk4gn4/oNFhouBCoGh8iLOg9VeiIlghhCQdyoBxNEekJqxGk5J
3ZnDPY3P/FWXacmCSEbchuOKilypv7iawYlX2Mg7drZoa3AmbtLenV6Lu/2VyiuLPOriJGzsZA8M
rsMJSeqaTqQMLu/sPotbIetlIn01ACc3U8PDaqvIFPCdA22eBVeVg79nj0rbq1eLqNBE9KNQGP9Q
8iSWLdarIOuUPDi5wr8GSHdjKZNmAsSKWxgYBT+0Igtq4db8/u5BYwzm+zhgYxovaPh82CIrYP4x
ce+HDp4N/qcpUxokwrKWrhrgYUhCvDfGI+CwVS2BExQm8jT8Z/Jgq0gqv09vGM4YunwsseegIwai
3NHtGAwSgnwde2uZBRXCcTfdqi7krpZiPxc17VKbAnK6h6ZyEaV2VCDXMbobOfNVK5Lgnd8aWflk
xPKh4znV4vIrx3NyvW4rsgPzqdPZLl3Jgmd2XYR0lJLyjrl0EgziGDJa7FiH2uGHMiNocxNB6V7z
q8JDpgfxH09vpmmCrjR4mLAnwdbfem56/SodtunELKS44UmJMsFiVYecKXwo7AG7WQoZbNW+HNj9
vPJ+bmd622tllKvbUBLETr9WFszIhPOTZm3D/AhFOJ7bGw9dxWgaS3N/YTTM14EZbpCi+C254A6j
pHRLJn4NXsRbMxDpsbClqrHCbnMQHtFb1gMzgRJr7FmSZuHHnbGG/U5+UmfuYvVkFD0Hak+o9N5f
3eydG1CVmV15kEmw6IXH6pvqWZlrPqJ1sSrv5gdk2WWquhSEghiZSK3f3GmDr/uau4nPcO6XszC7
oiWp40LVb1JyfAU+0b1Du+YK39QdsqOTHkqnkDBWxvc+hK9OOTdcz6NaWQbWoOI1ncJrxPwTmm4g
mtGUF8Qtg03PvqPbqqhYqYFsgaBe5qp77QF4v789B3SYTvdlnsz4a2Vf5qoZHgWrWFdFWDrDmMIR
LeEwP0q/Wfc5Dhzs+zGFMY2J5rnMVfkgX/6b69GlV8pKGtzG4/H5vQGlEoq4BnWWqqetTS50Bxyd
BWwdkGJfOXnxx3o1aTWdsSujQmE1ILYqzbcbknpo6PsvkqWcb/QEzEr8iSXBmpEqrTyOdlogs8/8
r3UYv4GFmt88bc621LySjMrEwTt2b6HVHz3LxITnvPU9gfn7myGZh7VPyqSqJa17wkxQ2Bs6HYYd
OAqzei2hn9j6dgrzqHzRIbTtW5y67+nUNPoEUexGulQIonLVdL/VvQZsKsLsuKQ+Yso079WsrGEv
pfRs5uHhcurfU46gjHVAYnI0qaFjGJyA0NXoNRiu1tEsgetNm7JEibl2wSwH+wkkDr2oH1nOTypY
qJE07Y1zFjnh6EvEHwZNGFItEo2pfKRebUg9sdvc8DepV4hu2LA+pkSbe1CRaOb7qGk6ESlt/c13
oZMLG3oCKCio2BzbUevFLWSeR9SZaLBd7mtUn8TIZ2C/7l28tUqUFPnWVa7D4uOy2tyeZjTLmrYp
VX3V2WXq+tmr+/umjTO8Jy1o9TDABFhFZWYud3vdrDu8vBGATxp6FkebCxYI7H2QP0BkSh0Ns1hQ
0H2s+oZgxCOLnVIxzgNVjqR7RRFUYzHKFIzLt2DjtPrUrl5xygpMGvwqJ8hkuAg3R9BzY34lhSmY
QeVWNufS4ey/h124Lf3UizpZv16u42YlHXuCgLUd2t18fSWVdoAxTELpO0eUkTZ1i2jaxByNaHAU
GwF70RyEloCDfshr3flLncFyvw6W5oNInnJbMEQ3YQ+hoc+z6US/9XIrkEbVOpxGYWkF0XjR1Txw
+cy5M6sxRRZ0XveImkI2Ts+BCo/qIZEieOjf0dl1Ukf16QB1WFr/ccUhonlAMx/vIcxbfKZkXPcH
pQqLPvUFEej5hAAo8uwqmu7ZHf0SUJn8/73LnfsydgOM3TQt/N7k5f1UKYAT9QQNPuWqetLnBzf6
Mj63NPG0JL8LZXDLjyS0a++p5yZRT+GsdCx+6PJ+48jkfquuY+B3+3NAh6+zFbhK4unQb+Ddlw6o
w3c8UmwegkpGbe0lTxe33LuiT5ZrZ2yqzuguaOc3109fiNqScyn6p7ZBek4L3bKnBKDVRtRuKo1k
Ka3do/hvT73Taw1mmLmXPDNN1/0cQdGrayeUt92u4ua0uehSea6ywgXV+gyDdg+LT0XnoVVqW7lm
wgP7R/rEsiSPwHrOzkh+iNTzMwUiMknbqp/RXhMY0B8sWcaC+gCM/3HZ8qq3QnhGvNMSwz+KO/u9
YgjPYcl4r92Thsui2z006pKEyWv1ztzv40IVy8N2CNC5t8EjXNVIAZHihtuzm7mg5ZaeOW6MTUwe
mC5zeNtEgG3pw2Bv3r5OW8wgAGGWH1KOVM6Lkd22gIutjLrlXP8QsuJgd3o9jEkwvwc0sbS+/Jno
HnNggEaSa0DIWN9q/3xUm54e9Rm5wpuFz9c4D+pODlLgDgMdcA38A4YnkZLjsW6EJKEUUQ5zru3t
gpNsbu15ghXYbFZU5U6td59m9j4qVHq9ROWAA5YHcmd3JKV7Rh7MngRG+eRxXrmZ2YvdarqHiYNc
2WfVnd/CzGIcsfPYBgpFfsljOUIrVRfVGEUjfAcXbampeJe4X011MTXnYWKniRx6DOoHE7kuCXW4
GsGAVqVqb10M9qYJORwFEcqEClHqL0iSfReKTKuq1C7KgA7JYsro+DWAKx+kWVGYCzNDiXwIov0u
e53XoruhQg7O+PLlg73ZLig0dqCPLBB0No/dXKQhsrnAEv4ZPSrsGxAPhKtV+zXFu7ZPP9lqtj7P
3PnR49ROzB5bEcq1kAy5fpEb+WrFy+08XKKlsR0sAVk7AUpqERiysoDs05qQE08o+23Yx0OQjiQx
5JddsIhzh9mO9k6hi8j9TGLkiPglDSDa6xYM+O9eaKmgwB+Ecub56vtxQBl7YZ/vEeNX5zamFNm9
QYBmmZvaum+iMPxlBY1rcoYyWYnLaBo35DKpDkNF0twMf/XXxsQCUD3zbpNvj5YEiBqJluu1P4oK
VGZOFWTO7Lv9qVswAwCudBWMNF7ZerIXE/iMY/la5wPlmami6VZ1APQBmIwgNF/xI9+QRfy9sFR3
PG69WzU9uZjJMOUbsFT7NbwU79kfSNCHNB3x7N7U1bAXnn1wMjMEELpsm/cle3v53ssutJqxjuUh
mJvl0mm3tJYz0DG1O/NvbxNY48a6V7qAO+QLTvzNDRHN0u1UEpgwpBhfxGf6YDQ6adB3Ojg+UH4v
gTIHr9e3FCfVRF9AjBovqFs0z4QG3gCdGZTp+KPAv4CERbW4m3o3S/kiwN9lamikLRGwAI6+Qxj3
IkGyMh8X2zZpbABw1eDApl9IS2YSUNizfLNe0egkychFqbyK3UM+eZZdo+/b9V3t4abBSpEpl01v
jwJDRtPsgXFpxn49Nr6zMT0VewQq59mYV3pEQLxs17708d+4k9AtXUsiI2rtBK0Ad3LqGzIlQziU
WUTFNb5JuNK9SUtmvTDdGEoczMk9o4W+sjF3eZlRXgXvyZvyXOO1z4ikSVedI1OxPLVPMAabowj0
wVyruQiv+2m9HxNc7La6zqyy3durb8gG55dLnT5+sWtM9tNolw3VfBfG2aBlG0ouBt/4s8mmZYOC
PC17XrdbmEVDU99vReKeSb8OujxDCvXbzJ1leHAdKwW3SaS16Wfd1YvlqPHodw3MQ2fB72d9mpAC
AicLt1mxpXS2o10NcgEMjH8g/vhcJ9HY0e28V6IplblhhQ5BMPS+XPlcNqXmqQIcqU1tv75xowjl
NlZ+uxfvt/jshiRgTPqcs28TZci7/nrRszhz3PcTD37Y7GcdkD9AA5vY7XrVi68iLWPAyhpivtZY
Ty6uNx2B3WpAXZt0teENMcevQMeMnfLw9+YyEP24j867GnQ2kguRDCj1SnfS4YyZnoHc8kkPcth6
ejzx5kAU8EhvNbyYfDXqJG5qy2fKgId2EKI8qdSI8lG/+eu7O2EjcneirV6DXdbI4glNFtQDaHu3
5tXFiOsByQgrFb+fRYhhaX0hVTCJpgN6Dcqsba+kzmcqNrdVO848T3Js0fEGLV9ChwnMn3SjCXGJ
7fWVfRnPrNw8Wla1FBeU3AjOLmz2p0nlTSrGK6YxmctQhZnvK99bgJ5OLyskLy1DK0chYxQNMLoC
o5SP9sHX4FN5aQ1cohN4TRsz8kXmdfozZaa/tM2LkbuPfklCXytxeuVgh4i88ri6r1ruG1Ii14fc
rP+Ip/InlEgBI4FLWT2kDz6bNmT1Y+kO1vMhIocms+NlqTbaDmWWdt4C/SoUSk7m+FBl2ZOMcTwj
2khk5KXOjRNClKxpO7jt2VfQOuDHRd0l4NJccrIf+rnyNfL6HMZ6IdfgrVcVu22SISSMdeOkx/si
PFDJc2WjxX/kXH64jmjlr8QAhC2uBFNWmE1WUlaKRo6sxgpPdSgcr6PhzWJqQ7XLNV2Khc3gVEku
Yo8X5zbTk2nxc25VZLivtccMeIPVgMpfmU7NYft5QAiBQJKEkPfv4RSK9Kb1anni4iws94Zbpoih
cI3MsQRpGP2DfcA7/g3inDk4EmOmJRKV2BNEmXXdzjuKsGq4eRcWEfgj+BcdZxaOqKQ92uXqOkSp
x6fSx9tz5LGFEXRG9i9bZWZp7qJUKT9O0GvzkGUottcw0TVWBE5443rX+Sq4dekewH4zqsw75tnP
YvQQD9cTnVX87EuFhKggCpfQHtUi7ag6boib78IF2oODx17kr/ZlHdAymP21RyvHpEDJcmBJa8tM
W9d9J8X7JcFjMmB9ip05vRufR5QvG5KKN6qRUVOWIjoItVPbgcO4eEYz5PAL8CNFA1ysSgXwtkLl
TROGYFhmXqkXc2RhzXnmBhETDnIpRMWpW2/NHOapYPNyq1NAi+bNwqYfs5TP0FwHlsTzdLf9foL2
3aU4jlNf9JgqcpeK+7xJB70YrNGZfB4AgKzmEXvT7k01PF+FMQZrRLiIz/zh+frVbbxLdckh9v0s
tRwRGl/L0z0QmElo+MfQm7c3BVpL7R5TILQ2FhCwmt2zBV4GfToBNukL3tgdelN2uvZfrgZ4hCF7
gsK0iFCcKGBbZpLMM6DjC1V61YuItlBGlG8rz3q9Hbn6jYuV2IQ8JKNqH5HM5s1mHX2kMJ+bCTq+
dRkuCLgqfvSi2HQe06gAwcFENb0vODrKslQREGG3uHamst/VMM+i9VdoTbOIU/mR/bcqv4tFM2NV
B1z+27E3BSsgkXMGyRc3ntgd2hyrXWDz3XyV/YE3I0mQ7ewpJ1lipYlaGNJUre5oZDreril/TEg5
MT8Y5ds8VqRQdhxyQF1pTzDLrmcO1N4hcLPy0Z3IVUibHvAfBS8iEdYhu56OWAFfcyT6aVvNhcF8
VAmzFX+KZ7Am9cTjC+9gupUOoH3qdmBy6YiE/r5uZxj4SyX7dYTdXXr+Ptv8/tsFrtH6kg+ysD1j
RrpOzghjiQUK1awsWBY4p7lJdBQevVcVvPZUpQv6nOAKHOkt8FmQQY3xDACPlSqKwW/VQSPwCcv/
t38H95d8flTr5F1I6HpQGQXf9Wk/3tE9+EWVRpfQcvNHRtj2AC4wNlhHKMtYPbX+jsiptXuJtyEM
ptUSFL++bTbJ6Ptq+W3g8h9F40tjN8LZZBqhQwS1csu3k1mJ1aGmJSQ2ggoM4Z7vk13hNlvyU9tX
OQiej9ko8aFCVrcrASDkPw3MuBLw5I7NgGYV+W35yqK6+1fa98lc8tEtSerb0aUYpR+7CoQ5wnx2
YqaG6hb5eDF3sCEpSBiQ+pWXwmxDGO0BaDEvbHfD5nSGrJoVWjLrp3XMNKJItcgiwPeStthWfw1C
KTmwrdMxoXo3xt1jEsX1JsiNlSHpfqCV4z1JIsOdUloK3QY6bzlh7e+XfTF8izaqhJNaUPH5p4fh
rUindxWzxkFyS5w8Crp2yitjeiXctsQz6NTE8OICFhn5VTajvXRIjBFI5V8Ou0C0k5TihMQ9o80J
lzP01ssN1sineAwGqdZtkxLDf1OzZmLkYCQjHJTrThv+Vcq0bH68RSzqbxrSiNQZHRou+dvShQRR
LJFJ6OpZsqBA/qRRg2q4NcgizOhwJnDghhBIjtuBaikKSbxlYOb1VvPU4goqo7GEV7KbVSnfLGD2
fUMJoHQGC/0/OsNbM5/YpkO/Ena15gIk6A+cc7EPVKDiQDJ1TXQgy57fRZhWFQlilHUXZoKsrljx
saIEZ9zkVFsCiW6LxmS/yl4XFe6QV+W/XbEsYt151qFhEgGqt62WnhqpHWxvGNtyOvGkMATm4VmT
WUjlauca3iMRgO1zm8pigXQ9YihLgRZEk10vD3nydaUJtFdO6xwxLFLC4lws/3K4hNh/fAa8j1Fc
3BqOBcwtXUcBR1zOeQFy89r3uksy21N9QCLoMANZbT6rvpHrmnMq7d0rEyTlRRAUVi0US/R8vCQn
ygMj13/4DHJ/ZndGHV3XugQ7tUdFLCnaBe7Jol8qzEWtgZ37pNoFiMNmm0EFnCdcDrdBAGep3ffT
odVkU4M+Afq8gdrQhb6kq38UZimTjBv+4m99gcKHKXXia0lDlfF92h9R/O34s+7iXmiD7JWFpMnY
Qr5hyrcrrwSX559MsqnSrD87+XHnD/9fsOZMTUxWbkgSUiCZZYOycDhOeFaxjlKDiaUeP255Jf38
YHigg6/4HQJaSZ7wnoWt1lnnrGY+/Lwy6ncm3KsvXD80ox8xRxEp/qj6gBfnEbfGkh8kwTWDMG3+
7eBMNGVur8Q3o8SaI8ChATtZghQ3kPJLm9spf3ZLZre7wAePo2tncXOSbV2U/wKtSM5fbR7GcLl5
8IU7fU6JXWdfxWXVLMC6nVu3TNVPTSQY8MUIrJb4luROvqOm9NUDcmZtLGD8JHpqatr0Gxkf0FOk
rsqjML3Qw5envvQNv4dR95ysskqF24wFoBKuaLAu8q39PWqWRH+KFZWe1osv7PfwH5J8iz42YGtj
4FdjVbkHD7Hn5Y28hnfwDM1zSbhEKUL5AhEuB9KdrOBQPeCMBUuM1zRIh6JGpRVTnO4oFgbDwKhs
7PH3boyqk4Zb5wIae0my/I9ZovimuXCt5v/CvLUEcKHwTzPtb17QHxTMqpKXRGZ/My93Nf08xebR
QPRurJ6bQNp7y8lusa0XcCVq46nMycCXEba+QqstIdFWZhM+PdtmWktj0R6+5U79gtrbDzggBYpa
iqtREpSOXLioEuTX9tJeSjGPPBvk0HCRimrcG5botFsrZqyGOkFXh7H+iKPZTsRyY8roGU+EQZbO
B/lUAyff2ZNNCuZFgZbJkdNPCloQr9bHcH+51cohhi9HX9vF5y7M5vVCdMXfKFu1JYpfnaR69qu3
RhK8szGuwIhfOs0=
`protect end_protected
