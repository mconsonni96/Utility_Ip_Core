`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
JIrfVvigpE9WaADoJfKb6VynW5O0HMcZ46NLWQUM49Z3veps6VPEeRiJCU2Vqvd8hB/CMUgtWXvi
4bb7wBr1Wj3IstPeO7FiQqaKh2pmYsPBCeJn+zp6/DbA7+/A7fjRFPSS2OcuOyY3HQe1MFcftny5
ZdIyleOSkrc9mZ9X5aybXJAfBDQask8u+c0MJ855h1fpKxw0aKYXqgZ4h1QBJF94KZwEDcyr0xTl
ZN+etvkGqFYs8ZOM3Z0Yizb0rZzNpL/rp36Wnn/qyX+wjoFRS4AJqSUbEoDsYEIkSo9c06IjaOVA
gDTWinEq4IeSGEYv+OZOJq28RWXaNEdzb/CMiA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="nbn94IeGBnvD9WwLuRoNw7w78haTndn3VhChtn6hjsE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19344)
`protect data_block
XlWbTtHciM3qsJRaRI0i0AphQI4T78LXpAnf/v2cA/r73aqd/aq3fRf7scILlYgeAfQ8Vr7DJlcq
Mtnz9ZpR2Xed+yGyPNSR5tAZSljA/Tiir8GW+oC6MhVKn543QFj3anIX8r42kLGq6hoPC7zXz8Cg
xtY2prRt25Ch7mni9b2T7mZg/KrLLIYRmBS/niDXWJnAJpd6sK2m6OO0sR2N27H9A1DavYGYi9nt
GhrBRUugdsOjDKXC2WPp3TJKsC3R4ial7o8l70HSJzzGrWT6sujmW0divqsM/qQ70PrA5PjbAEk8
VY8BuDON+V1hjKLCYfuyrwopqVHweISkOjDpBFG/ibol00CJW4zRChAaq28lGrRvcG3ZE058ba1w
zaEZdwoOj8CaoJQWLrl+wvI/4uMBrqoFSLCIJqxDf+agQfRNgO6hAdfLas1O8+QTKISZFHqgho8M
M03dpqL+3aynnZiH2jxsgJW+ExknlaSIv1Y4Gr0D13Yw15t0gAns3yWbrU+jWWnwokGLp2ShizSE
cjlLW6H5OGv+UvUiKRFHDIl0JnLi+V7hORUh62oLnvu+RsARCJGi4OXACpsx81d5nOkc7Si05erE
EJbRSta3h4bOOhS5epYjeA7BWWTZN9pn6KaHN/O+D6lILfT0K7JaoLWmd2Hysipd6egEo3pAM+T+
G4BVEWYrdReIbfd7PXxup9AYx8qi2bVr9jhpM70VT51ie7ORg4ljkO4e2z4nCJTCDmd/Ctb7/wzz
d7X/Jt74Jndbu+Q/EmCnRXIZFLVd33AAeSD59Kc81USQq9ie0Y+zK4jVMyX94Jj+rwcdglzzoODj
cpe4Rz4yNnQL53T/wFN3DCyLQOwJ7imGo6kczuDRnqHpyda9VT+zmi33LezOd5XCBnSeW/av5/NV
SK0m7DNXig+nB9lmcl66xrzSvpI2owcdEMKvMQVtqx/0Qq4F6JBe6jYIASaca8MvlSBfX5FqDYT6
16lFDcJbcH3SkjePb0CPX3eNHHM6VNTBlcZeIbvXuU+VIP9r97rtbEsu4FMhPmUcvJy04Tfj9HLr
fqtGB15GUcdM2wxW7ShJHxIG/uTmfMkZ18ma9ZHWjMlTdE7LE61gesPYtbc9r17yJJ+mRowaNeWp
WnYCYaPyOgJ7pOS4uKuWBwUxVzpHudBkJBu9QmkOjIHEO6riK8ZKFxSnOdUy3KAWXPT2kIbo57zR
xRe6fve6UUHOxIeSKuaH36H6urgOAXgNp6kr8KNr3TD+Q2x0Xa+oHe8qUfe3w/qAuOgvJL5nFmM7
DJ01mQOnY13Yh5T9+zos1UOFYQgg6v8pj/cAqj4VVOgUPFlUeIXHmJTfPbZFm/B1J1u9NcQc6D4p
DbWoEpQbo0TPYNlf6vGreyN5yHyMkecRR4WK4+/+/YNEtG28qG4HbLIVaOk0CkuBLTWxAePRXEKt
iiT9E2QeHxuoGzNRnuH1KMoQHzBgUXX0yyZwFvDAMDWQT6YR6TWGxhUABDh+nY5Dvs1qew4Xhd3h
8VF2XLWFZsA+FT7+Tk1/51W6XpaZMi/zD6PGa7M+P4kF5ha8GdmYKmwC/lfQ8GtjvxTg93jrPjFb
I9c5sGkxSd8xDDmDqESKi8/Q7mhxJuARiUr+vWYlL8tep6ry7+ltQ6rq1mFNPsmAuuhaVxE2ZtDH
wHTF8dEaqV+rK0lvJ8pUGx6jnwrtPpohpBRLEAxJHC+GmwPWpyjeeL6glQzETqpySdvbC1IhIpYf
EKNCX9pAmsJo4cmKaEx4P3/CxAPOauv4F7tk/tHthIRsyitRpZQLArJLI6RHS4uUii+D8XCRcy1G
HFCUKVK3oriwzcRVT0LqbyTNs66WvKl5AuIO+YzbJF8CmSlQRWeoR7UOsP5MB1qRzPAKAnCbfye1
zt7HpP912xjcgS5gNKLvkTr6r1XWInvVKR1W8zmHQA8eERsoUWapOpUO5ucJ5tc5YAUEbptu/MLV
4rubVvLy//7We6KEVoB+3lvzGHJ1orKcq5jR4K08Gh0nzBCzCOdZ/qCx3S1qm6PgGsmU3d7WSx1c
SbtrhK+VXqBar59EOTBZ1Rdrh34r63hsQByp0eMOG11JLmKkQPJFAclqWBh9uXzumX3e4PQj2yXz
SztqO7ZBrklRul6tiMzt36FFaWb8x314gldxz0mSIE1gJVObsNirFFMQROwlOB8ZL0f15nv9QUsG
CDDARdyZcyGbuvE8BercPk4islGuT3j4EXczt/752Kz6vNqTWsbcXYS8/2qW/QVJ8Mloojy1yNhP
rzSk9nb3mlyvUz0ghZmfBrMfv8lWdjERKssoX7AhiaM0k6zZ8y8HFb0q36Q9+MCn+28XiT9YciAJ
otlMTG5OoAlcixCAh+vRs1G9UjaPl9Hpld7KqQ5o2Fw6sP9qmX2aFSsLJmRzfMnvFwjK5la25luV
Z7BnfecUestvRyoAVQ/kE9pb4y/Qm9pYn20mDv9W9yDIdzCjnzAzx2rKI0FczYqS/2TqGIO3azmm
V4SSTRC490yYLzx5aC+WXttEgAPU2p0qrglZuAkTyGAoU1hrpqIZUciFCA9zG1SLxctCsJ99hMOg
o5ABkH/exRKa0CcSCEddQ5McpbAaFE7bAYfUDUVIhvWdc+8YgpgATR/8iFWbJ+Hl2WAbkUviRpIV
HTrLnqfZsVBxRHPiq7gqeXVGHiMfawNTIB++27XtA9rF9cMnNKcxHIcMSossAAcJSgUa8iy6EHhC
Ow78XhYKacr7ybP7UfZhMZBggJrFK4UouuO39oyylZVlJUXeJhkc1elHkaYbwHQUv7+WBEelJf8o
nuXu80HS3J9bFKkh7i2DtQmh1UEoBpnalp9vWaBSglCEAri2DHLZ4tSKU6bfuknBSZ4sMSfmTiu7
Cab4v4Ik4Q6OTtoTzZCyyc18C17jysUjolu8qt3lYvO4hlPXWqsfcCKZcR0+FrFQvm3tpyr3IWhe
i+2WoQsTVRdDnrBEB0YrS3o9anj+/sd/9qXu/jwrd+O36FFo/WlsGN4VMCUwTz2a0F+TUo07N36v
v9yttTe5zCnSvyFlfIgisX3SfZB9ir/BlMA/xOhWmQt6NbcDCmWXXvxGms976SqZ/vO8mzTp0/df
gaWOqPmPdJ/3kwcv5oRlmN7rNmUUBeNT0CQwzyo10e/Qb/3iwF9GGIjkJsPfIlMJ6+Jpj1FzGYuQ
qQwMQWNUy2mycpTPx838qYB38hbOEw0z4KnUFcqhUVaBLoTh2UjjfKnLpYhWjqYvXM/Yv836i0Ql
jkUkKqgN8HC8N+5l51MrdyE+QVsiho5ZaIdy+nW72ZItkam+C5Mwi2VwQbXnYZIKH1DjhINvS1VK
sDGsJnJk9Xg6qrdcAnQPAiiK4pf/pYpkg+cDJvfCTstfHiLGIQu4s7RR/KcxpQBfBinqL+Mt1pUj
9DGw1P85cMO1LCmKthQaomRdzjp1zUS/e8EZRLileKKqXKLUPFp/J4YXGJ7AVX+383jzNx73nYrp
jONAvXnqhAiFMs5m1dovnNr1oYxcG5jS4Sk7hsYt81pb/IsQBETK2j2z7Yo3jik45EhW7V8nvUGP
tLuECuKuyIbR2JlcjE8lnbb3PBxg9yWhM+FQnYZl7LYXhkxO+hUAewfo7J1CVMRnguxHmH0O5iD5
N7SeIn+oYy0CTvK2fSms4K2pDugs+XGtSMj5bnZZnps3P0ksolVMhWQbHJhw37ncpiAeKdY00AM1
aPs8+vz9e/hdwpjEbUhoPtmAfc6Ge3D3/CtB/J4YTPP8kFM4IEURnKBPUaZoAg+kFxo4vvIRXm1J
ddMxMGybznb6tIbzdos1md0r+3/BmqGhB6PjjBK4iylGJa25hOLMG+Syldcu5NVleMoYh77iTPX9
AV7HtjNHh4UlI3zbznIXI95bgv3IyFowk1ddVkBtnVYYPdfsB3nXGijO1XEmtau8BGqVmklBXMiV
NVNgFUwljHM3RA4Teh+UnsM19J5VnuDXq1Pi/+TzeKIOLb/xQ8lF/u+fuohTfLalW/LIa1posKtr
uh3hUf1qG8V4eBYkhn3H+A5erxhZN68W7V3rTyLel/9cq8IZt4MPwTpIeZvuKTacYtA+q09b0eK5
zt2B8B44KSWqFxvHAlZpxOft0KjlLcxYeg6pRx5pAAA52grTogCLiUhu2mK2hYqSocR2JMtYGam4
0sUhY92bKYLfhO1ZoAYV872pGZcIn0Y0MOiiwftA/lb6KzJzerPo2K2S+HcMvA/El5Mvrv4xKCH2
dHQp0AbXlQs3HWQwjjanhw1IbNuKUAe9n8QFgHn3gbEL5riRn7mzT+HnutOt09tmTS/sbPWmHtGy
o/897mxYRGyH4iPdoyHGVjegK79djRP915UOBlkgP5JTp1SKFaey9YFPj+cLKqKk2dwVmEQdTCd1
T0BiXrN8l1igN9H3CBBt6S3ESE1gdISfds+ycsj1r44JlTfrpn4nF8kgcthU5CrsT5lYNRAICMnd
B/DHeQPRbTOgw0AdnvAfWCojbXM9ObguEoP82puRQakNuXyCRySlYNt5qtgvan84n4dJhU9aWTtd
wNEbeiJmy9woKcEG1GCH/8tX/Fwxf48CNsPPLaFCXPGFZrar55VHfBtL2UUPd6GiecwiAZ518wXy
4lvHr8NLlybe6Y0702yXLsUpRLqfLZojMxXzSL6HkSt+ijp98PwTls9knP6SqcXE+F7MJarxzAKX
+/aQsvM5QoeyYe9TYiQbL9MJX7TIm6LreWpYTMAtuNFE6rq1ymluO+hA/SWLuxBBKBDYL4lIdSP0
mWINQ600hr9yIIr4uq9uu6pyB+fe5m/1e3qqKewPQ/Du66X2bcqHnJiCgluxeLpdF4ByqbH1IlFg
rHWgqoT2mB00WaOcR0lA2TYEEooXeLdcoGOGXxFrRi+hgDKZtniHN288H2fRORNLm4ET2hW+3GTX
JZObH3GehsbvAr1RM5ZxUuo+X5xvw9233xbyoMMjQT42NMoZE+4y6W0xKM5a6vua5KNJssHHjkYh
0bPb4miLQ492dMrweA9vC0THFq2rdvWesSzAUwFpAKjwUgA75AgvRrHY3Fqf/tcNv7xalwTrLXqD
KrYQIXPCvWPM/Xz37G7etbL9JA5cUGsbnJR5ZF7bJ6SS69F6VXC5B7m89FlmUcrgXfxv4L/hyMWd
i0xsi5yjecf20DvxpY8aLWjwy9tT5FERw/8e4Ae9WEzUOZEf0ZBTfyq9ORo5tiK+hn6dVjyJ8yZQ
525fQFAe4lA4Hpy7ygE4pZct1Ar1daMhx4j9T4WKONYYEg7Ib8SIADbsaHrj9+iC5BZe7fJ1N5I9
CsIpmsoMvQyEv4G3mbnu0tyZv1tRxlocidg3m2aE2qzb7gklRyzonHIaz/Dh8U6g8kcPRK2T4y/n
fLDh/o8WM/u+A/eyilXxL2env0URxlIWjlfxBzs5GkuOlxz0CDr8qC+moJfJ8Lj8gYPCnXxf1QPn
XugcS8zujV+O12Wwkhs6NSQJrE9hL5SoKp3x2tdP4XAhX4M0sfAOKPYV9GOj4nuKgOnDovq/L++Y
c5cBhZis9VZ+DxDHHF1lXnOEJKySV+0q+hRjIA6Ef2VKnS4H17d9mZlRpmZx2/H4+8oGcs4TS9J3
l7jdX1R593sYTO5xvQi4Uzl3qtOtT4HdpfG3UvG08ZGrFj4kvG+AfFAv3WYCzSzu9ixllZs8j/Kk
kCJNh2QVoWLUVLeLV7lhQdErM6cc3zPkXR/m7Z/VOzIzIYpEcrk+bABVNPq2MtFMUq/kLv/5Wdh6
mioRkGbLQpselTGgQ+qE8BTKkMaS74Y4gjYbaCOuyYPIIOFE+GfSD7nZSLFTObh2bzTMUhdEnuZ+
Xx59SsMZ5jWXLoJPYS0rMORolNKXKhszAqaheZMiZbQgtefuQsFTkyzJutz5fmCuyf5rqzthhaRi
ALFpU06TRQw9Z8+BHYD8xubYKDFIkLd7m6z/XCLQvvMO1KdkQisqJRfmzymUBfVWm/aGY4Jesjn+
q4kdEEUKRRsBV3RvKRoMKCctcbC8kQxiFqdY3Z2c+CpSgrcHQ8OjvtC+fr65C03YiHHfzR093J+9
o5oS9zyu3tYeMK/GPTXRijterVklrLyyRB5QuyUkfO/HtptooLqSvzltVaMApCvEsN3UoRWC9YYQ
HRXrQ9CknoGgO36qcVYFkuiLdWaaoD+hOLktTJ6lNL3ww6gq9Vtw/X0Tmz5WoYw6EbnMqHQt0AjI
lpvrQenbJTCQ7ZZpDai3px07qeonewTLk6OAfB72HlivlzEcWqLrYogE4xZMzvxVBqFu73n7AVMN
b6hsPYMAadnjOYV4xLLGwiR34HQ029I4NFpTXdp8Qfs9ah9UlROCDG40tBcXsB4LQAJyP1y6sclo
XJA6E13AvTIfK6NkbZuE0TcrCpwwZRLGI1SDO3Qk8C/GSGluUckspFLWCsLkBnZOjawVr8DKIMkJ
pkMmXJePm0QMCQ1QUaoLTCH4OpZVYb/2Shei1jwo3kJtN4mwse8469TBysWkygHlD7dFJnjqFuIC
2tejTtqPf5LK7ziI4umeOgrByg2o+hgk6FBvfCUjM5pl0wFac6GMCVRoyBr4Tr7tvA9Qb+xt17TQ
K75Jj1KA56RHN+YCf0B3usIttr4WOBqGGKQM3HcPmr0dsOnQlaUobcH3P9BVvZlkfbTbEPRVyb3x
9H9tZm6qdufCB/Job3wYeJy/dPox0wlSHJoz01V98U69DaGCRJzMCjCbJusj9OzAjrGZ9aMEjYCk
CXYbJOjxEhJeduIqONWuF4WcySbDp0HVtiRUYzpZAW+B1/K7y1+oJu+orq/gy8JYzG8RD0Nk4pp8
b6+al62bp1y/trh6kTcmVGXEaF2nhLIIRdyNAN9DB+vWSX5s/xY7u2KmPsgJ/meWdT4ZeYD+unWs
JIOJVvYDIxS7tfe9N8njBx/sxW1d6yij0mGMTuJTG91q3rXE0Bo1vH8vAgOyrLyS/M/Jb5YcdHXE
jod98gVbK1HJOCkbCceeozdY9NwLLBSkEqem4iYcDmixXSyPVYwYizGBKMCCQ/uvkVvQEzWx6yYb
ZdGPIhreiltkIdLZPT+4gD5CD6XfoIhEfH80XvqghdzxzdPeQbgjt+Kdm0cP0vKjYBfwu6NInsGV
Fir6U/2jGTN2TNpCigvgB1jO9kwrWsmFOvo75t/Uh6lW8ixQ0F1GTeryDJz+vcNk9NbX4nUV2sXv
mWIcJdFLWGUg6Dysd4/mni7UFy8WjlpuNM4lABkTwatZ7qDAJ0ByzH4ZSsj1OIpu8hr6v1PS1ziU
j9ylpYuTYKTPpaF8zPZGPN6KPEP7t5QGHG5mCn0+QksxayKlgaLboV6/syaBWxFmfVJoaMp+862T
6xympmMxbPXNX4PRTTv8ja4vLZpF5ywDIejTNEi/TXbg3HWgVGKgtZh26MmNmtfY4E5NbFMJpOnT
v0Fl37xWwgHnz2iG58UfQCmCE5CDSubZ8gbEDP7V9F0SJVtc+kWaY3TvrMJa5RTdcmsNFluT7H59
p7Yy+LrwG1qzFUwgEUjw7g6FZIJDaYGmKTIQbn1Y6Wsggt6Z1khh99C0gaknU0pCKb3zwPYMpBaA
jDJqfQPHOUOdUIVZD9r+9X9NqdSL0AajcwgN3tj06PeBFdTK3CYIYGRl+chpu1brx3AhoausQs+s
fe9Cj9LXdAN58BrviEnZ8Y4+u/olWeX9LzSJ1szir6+Q3q5YiLdB84h5R8U2qtvQyTEXLamPgf9X
VpJr6bUHDR02B0tp3cPbb1PplMRQsdpzRpgfaGSaZ4eJKMTigWPQi2nZjgWpsHsoLXXM7Zp6Pa0w
HW+fiFHz6jV0LolGl5ZyYu72/5rV60XZs7/+KUujUi8tVj1C6rVGUl6shuLJRRzOH83+vzm99DV5
dLnWpNlRaGkVasmpqsMicxyp8cfcwxbUQdK0kIjItvtP2anICal36utuyM3w7hheC96eDzw1gAoB
wJIhOJKlJ9uV4fqHZw1uNauRvB1su2k51xiCQqaTf3iU/IX2AqGAbVxlEqDzwA09iYo+hBewVPVG
NE6cSvJVKCujnPSduKR2omMgPCsJJI+w/mspplECW+tjZHHcvsN1sy1LAExZ7W5/K0iGgX4GvZaS
guGFySphQpw4C5ZeoIOJDQrRrratMxHf6KEPK/xPFtqlM0ncCAuMelcW5GejdVAr+UvvqVBF/x/F
+OtYqUobNch+GDU1nrYBYsLOZspYL/mr4G3ppJ79tyANV0XEaAC3VVHxnIiXcLPPEZOQygt2bIvA
ZIBcEjUtU+fA+FB6Xnd800GEdjfW9TutujZysgA1ctPzrqjCqFEwKjQEYnU3Lkkm1XHs7LfMfw1X
fOitVE081RASOc59gLiV4/q7Aom0X0jtPjTp1VrtMWl7L32bYdJj8hJ3Xi4JeG2fKR/xtzkaT1aS
fd8YaO6wPwUrKfdOp42od/HrU/izXc8W6d6jZHl6GtwRQFDDj9sf6j1L5L+x3XphNtD+nQpCHInu
D7PxVhi7cS7cOV8nOjBdjkUJ2SiOrVQIQk/Q1G4HHADoTfWOgVEFqRNqVZPNdEZzBsgJDev6GxAy
OskUdw6dUCpkNCKEXcQ3EDDTQV6WWrckOlaPq0dO65YFqMz20V+aF1dw031kleG+a45j/P9oMv7D
lmBAxtLfzsqsRHPJ4XqyHRkCRhEWdMlKnAlupCgJF+65154vEJ+nr/ONYwitcoEBz3/8WeFWAUwa
+4wr8I8JX3f8WhxmIGxLl6jGYkKr2UzILABIWzRV4HcSFc1Bwb9lFjcu6zgcDC3pcqRp7/AgKtjI
zfskPLCJKTBTrUhohn+Sodn4QtEAavPMoF95rFm9gV0CmE4NN2UbuB1vDJFNSEJHMTGmUmg7FuYt
Mvm6mCKoKg9/vbc+WjvJTFX/9Z3yhFffsM+FaKGK59I8rA9m3bf8PSuNK2QFe05z7F7VaiiwOk7m
sQLgx+jYvXNrCXBhHDFtDghfGEyMqOmjcmyZK4lsCII+nqwFqfTpk9wPaUiJrNiQsbaPWhrpkHdZ
aBnuR7w0D18at9lhLPcOcLX5vkU1Le3Y+BIbwHOTB2d6FA3mTEPg6qc+Yhe/N7gZNGyIHepakRAD
BAcWPJx2ebKOzyLe8r+3w1hnpAPq6UrVzv6Q/PUy+YpUmnxMd8A5m/bjxkMKZOuNQwrwb9i7WQFs
DprOQVsQGzXcwrawf32xnwvqWCcwOej1s4qfBOXxWp91Biya4yLocjCoh6xo6pbHpdFD7MrbCZlQ
2KvPxce7LDLonTzf//qIDaBuChAbLF+4rLSSUq/N4PZR8xYhSjPFIeE6lh8rHjKxWHS7XWNu+8x3
ovb3Dk5tAWAETvcekxlgAJwzFSXEGedN1XITMj3IBYyhzwXm/FbJe87CSNKQLREMQuJDHMu0VKnX
xF/g7Z+oqERx+lqKUgVAYRUjVsGXDRJcUlQ7o16ACkMN+WFSsiB/B+1evWz6A1Y+gjsN2XAxZNwF
Hr17BoID55Vw1uC0MoGF77Q046OUXRnqbbYEC36NP5SMXyugM4PLpa/EKZiJgnU533uOO4zZW0qz
mbJtG+8E/7ygpxJMygy7Gss0pXYWZOdgbgXVwc8Z5fgBiPNo6VnSfUzUpzgb0690ybB85VAgzg2m
kkeBBzd767FZg+4RsX4baS03XRUGRa7VH7Rh4u92ncpktg8TMMLW8mI8LK7Tb5ERSnMl1qc6bg+Z
7wkwC2tXR0LKnZA+EECNSLF5shIEsQWvlSBwEs8T47Hkw+lyGILNrLIgZq/ULD3SzC16LUnwhQoS
LNjS02UuXzK/awi7Lr78YWTPiGb3T8/gsUEdA6vZzpKP845ho11pglTIctSgHvdRodcwb9A88aiU
za7xjf55pZC6a1j/LJHwKe75b0/RL538WGyGWePCAYMtIitTOXLAOpEJUeWdeOA9wECP1QJlHhmB
lS5YXto6CMxdNkPGPf4JuBxvu8BLVPc7yE3KCLFoC+hEUpDJTHN6NpCGsbH05C+Oscg1zJHEZwhV
QXJNeLHXr4Yw0D5TF7QLiuhcr+7GWcOzlzJDC2yg6caj9S+TJjqLftIp70qcr1o+p00l67zqGIFj
wPkF05isdUQFOuIa1s0+1bukI7HGTzhszsO7Ms4qg+TmBvLBU/15kf38tTbthfafIm2ElFBaz/qY
pDmUVBxp9pGQZaOx58cferSVObs0XbBGWN7uS2CDDsALkpza8XzujahYkmgmBv4Bwae8qp/YTm53
oVREN9PR+793HfdmpNtYPaoqEaNsDCDCaS8igWb4RHkpTenqOAzB+LKRZsImaYAjEoea+eACpsPk
1L4IX0qcgs/cyHLnTWy1BYBspigPBv8kU8B95uD5xve9FLliIVUw0bWdYXjbFm37LjJkOLNVJj4Y
GUUxYrmkXQHHcCQ1bjNC2LEY1wR1heQBXHn4LPNyzY42RN0fHa+ePbX1PV0u4PbQ8MKjyRUm0QyD
Pk9ZrH1if+ESPGT7MswTfd+iacaXaM4Y+xp/GdA6zwjFHD5bNHZ/RlDXnO3DzYKMCg0KW//oKEzI
VxEdC590dGb+dbegEdMjkN2/q/VTtxaUsEtA/x7zS2Xcz+JbGgi+Qsgjg4BxMkS+pofXXx8OsPwT
j2rCTFz0U5ucHQ4u0hiBNWt9Dc1vYfT7ywN4R2i1EGmcl+1cswfbKFS2nDPdPIBSdOT/zSUgTN9Z
AYfHsgSbTfgLulVljFaFgheeeVnXCXN9deLN1IS9xaVRxPpOdA4MIbR8Fzf42WcnoqjEw7tKAuec
8Fco129JUUAI5jmY4nNPPFWBgengVWI8+WNmzH9aTmt0Tr8ECFgCoUMUbtxFCiJmLPGqQZSwFTbM
lLBUfP6mDchW++87abSlRNLbbIyzSlMVx8FNW6cIiW7Sqqt65QiIEngVSf/g56WghimoQ1ZYPfKz
WA/g9jKDySNj9ocrq2kEJry4zeYMl/wFhEd1xE8AvntOdhia6IM0/K7ddXEYmqIG0ZfiIv4pk6IJ
udKYnCt7w2b/YAhSEhEdKRgENDAOBbyQu9FXoE6P2JF1JmZqX6LnLlHdRP5e/MNGM8GmEAk82PD8
leryuH4B9Lqz/XoYlVNcUH3FwBKZNcZ53JzHeMfDBJabUily9WgRH0YQC1uDhaLVIEvurQSGElQl
SAOQZq61+l7PJqaGU01IU5+S2ZVrUo/2KNIiWZRXtYQRdtBTwlk+PY3DeDS71ANSJqftiLXxm044
oC4lYKbrRwONuu9n/wQdPNnWbhlxWLTe8dTMEX/i9+hKvZIuO0LWuaYqiswF1+LqCvwq6+e5KObf
HjgtSjgLWEF41HB1QNGXty7G9wgB/VxMGUByY1dgqRU9wrpYPzNoBjKtekMIJz6cPehLHocDX0v0
ICSqH4A859ck5SMnWKARAiKOfuf0ISaIv/H227TTuSPm8Su/+qHaSSBvYDY3Z1SBcE1HBiKPmMrS
Z0mTX89MZXCacDcOiUfxdbO9mDdXGullBhF/6pUi/KWL1Suw+BaIt7Q2WJf4gupTasmRzZGjgXnQ
VY9BwyTpl1MC9oZmIlaOP0iZ61YBtzZ0Vfbvla0QTPe7/R72Kk0nuPrp9Imw2tUULlCbLnGwaJr6
mgquKcLQxAVrVJHq8DBAHCVZAXRI2aBuC2shADZVfMXcfCxZJ1PlttZovxdsVBJYWi4ytus27kVW
UFUiELnciH8N3d9ozb62jpR3fDobHme1N7125hFfKhjTb7DliF0noF1mJ+EfV/fk7A4Ncceyof8f
pNwV5U8AznLYHATlJhfCpolTcOCFeMnJuzrNPAY41PVNdm7RFWv1p3jzusKx9Crvw03kZn3zfxrf
/aG0EodgELD5KcWhw9W6oLbbPEci6hxiXMBLpLcMTG4l0nW5eOe7i4M4lKQw92irS0Nos49uMast
uWgQYJNSV9r5fUCZWlukM/bkwUDRjpGqfXJNa8TrHUB/FWAVuOrgX/y138qtpvZnqmNsaWJ/wB2+
fIExbHcYQv8zJRu1rqO7WIqvDzI0BKYaSEDQojUYrx4iCoQyA/VQMxBn5RwiWksnqWgWFQsQErEI
A/St5XqP69XhULsuacLGP/u5cwpPIT4EBsEh9Qiwm1PgFY5ycBP2y8FcIdcXZe+NKqG4jDMqMvHA
GVpEdKfKuNrLgXtYZsrgXB4Qczf+t61FgFtoOFzQCvqRMuou742xsmHMW9GY6C/cn3Etr5N1DmuW
prNpe3OztDRviT2EN1u7cEIXDK6keWk+Wo2efEjLHPQ55KfqrjSshI96qZg3tLxgv7NsYHRhf5w9
/SoG9uXbXUVTxq32WkrUSb4YMieY9CS/A9SdzlKYPi6UMyElt2aH/WoxyTT0mjC5NEVdaZxz4S6u
bybU6QYYrrkBasF8vidPejzZFuAUejjyVLBuHTz68Q4tzkQQPG1fUCKjIe6GuQYwbzI5FaQxYNfc
eE1Bm5hjeExwLrpm4xnD5PxwOrkDCumsIJaUSD4sqVCNdOHCSsUjyKrBfRobPshCQr8H4fDw0Qij
VeY4PJ7WZTr5HGnAw3m8oPkcxrj/SERJuAaRynk51xiDvQJ7bX7WR0FhOPgs/EQJ9/wG9HHYmmJi
POF+ETmAe4uUaceLq1AWho4/EMPb23w2o7mkHvIVd5vMNnJutnSu69mASMcneoXYVIP9y9YiPp9M
8u3DKEtZO7VpCtt5LeeIvunZdcxYduetkEIWNA83VH5W29Iqz7CZyI3rNVbtBx6VbFaIbHS4B48n
LutmrkSeauqHXtYVuHg2hA1FyOysgxt/+BMNSbNpI5manBPG9+Dl52k4/OsVKZQxdAHiwgowtSXi
luet2p5cqeIpSmy0H6Jk3YCeRRwyefdW9QuOgKUwQo5X+iEYv7Tr8cnd5j7WVCm9IlXkVvw2qZiJ
mRYYd4joXSLY+rLGGLNOYHYvRXycEn8aCBbJjAN9Ki79sMO1mDxxX+X4OFvo7pTJcJGGp7sRUoT4
ZzeXy4YeKujWSQS2yZ0eO69o3EDttuX/7zLgXEVizU1jKYNVf3UvUHiPk/Q8JlSInNLHw/Arj86W
Hhz4BFtUKPp9+bYlpSn0kJZRTSRuoTiwZhSFTgT2mrDFvHZNT43MguV9UNosXmzufikqNDHhHl+J
Sf3xvXShIRyt7lYZj9NfDu0ib2kx14yxFA4pkWl0BuviVyn7VdDevDMhynqoEsk8emXKNZ14rZB+
+LePeN9z7qaywnyX8fGHjNfq60NfT4mTGXVehJfTX/NdhAWXQ2SzQOkYc1Semaor5sWyaebHmJY4
1OB/V71eJFBJgQbzGi8yzULCtdzW5W87p7KD4bpG7698MmXm6K49jrj3gZMylVi5A7mImNWj5GVb
wGFFS5M0Q/6l+IFNKtix8qFYESknunNaswPtrdrDFPLzwGnwL3wC3N1JP3mXf9ED+lQ89/MjCiVn
D8J6TEbvig2sCfOBHqcz7+2MY3emGx3fKzT1I6TOe9Zv9h4kNphmZPB5yIIrI7KQxlqBzvyDRS6s
8z7sU9ba9PY8Yp+jFKToEYs2gzsBPKeGjlrl6UufqPkk04cd1xYkSE5VpsLdyRKlNkJUiA3AEHmG
V84L2O9aPYsGZIiWDzKwe8MZtXo/AlrJeOjzV7WWsyeFeW8lMIDpaXHJ7nR40YULoHxdKMivQVGU
x8S8XXys0HRkLfd3zxt6Jc+eKkulMbCEoUfM9mjfAUZh9mntfKj0rBBddjGOXQdsRh3imR9aH0Xx
SiAWIAiKFbUoBkVb6uWIIRRNYTm4jfJV09BmfzznmN/D+S/owdylfn3U0slTYQR5TOybDzNMrJT8
/bSWyXGk7d7bnY7AZahggn8pYUjX2M+0QwT7430zPkoVl+QtQQi0TojH7LMVcb57x11KYnh+zfMc
3kDDjlnMkOtf9BqtJrMvAeaCSiu8byWfM52y5tB5426S60EiXFYgMmjIOiK9cvrl3oK89+jaIXDA
8NUPU+JSXrVC2VL6yYexC6bXE9jf72NXrpTMuwycOZQDYioIoa1eI3FvEeJmklLvzv4kzZw0j0IT
Jr6OIBcB4jBvjuvwQzeHifCCZWjPt+2Wu+0olIjoYrN1H62KZJcwzwnHDytJOzvg6FXrMcQQ4m2U
3QzKvNspRJNeVK8EK0wfIXtAuiybLO6UhlEBW0VuSYk4nbO6L02h6E5FoSB5BU1A/+nys4qtG7XB
nkZYGtKJJ+L/Wpm1ytjiAgfq6VNJ96mfHrBN/7oCPd0v93v7yweGvoCQNFrNtFNojMmxC9rsEoQT
nDVBYwv55F8q+WqaO0XWndXVVtr5fg5eQC+V9Za7UhG9Vfqxbxn6wNpTw9sM5Va9elc9yelFDQeE
xbzp9Oy6hOPR8oP1rHPoSc9qR8wfal+XNFVaGTgnbV/1fMB4A0SpeCOM0aqi7dtSY6Fx6LNdQHDv
frA4rN96Ee8zWq66lTgkxq2mMiYP3+9wEYSWiZzwFWf3LP0mnOLIU3eOtv2OpRtqUZF+9vESdQvR
JNYlmHR2Uc568AuwlvAxB92Sywn5tQXoKQ0h0+4+K+paCi1jsczlTNRDMV64oaPEjsvaDHb5B2dm
J/DI/HZdotZuWPIUtHEdoiX5G6h8OLds68x4ZpgTF55sDx6EgJNvyKaR6RKSLnn5nod7OEz6gE5D
NsfqoumACMKfHKtabOmaZUBEQ80AUT9fS62Kq9EBrTOqyapkqTZG2rf57ohSbclV2XXCeHtwooKQ
X9jwHX2zvAEgICM19B4izOD2ywGxjwgVZSoYLxYanSmSOfgOc4xlvjX1wa5DB4wWFIwoXSDJYbLd
+KvY3dNp8gKso5dlcpxIvUuYNg/kH6uOs4vG/m/XoDgvaOYkLs+Ws+uSAp+XSdLF+BEvb6PLY43B
GJMCdizC/fbMP40BG+ZmP5IkAB/z3VeieXAmdDPzHxPeKnYBmbX/m6j0A95Ehso379lm3Y04y48g
Qj44s4kCP9KTz7hnBjYmOJFpW17IaiKed9iZ315CGXP0DG6jycY7AsIBtqFMAYDl3rUzmUzXz34N
faMrxtBkNkBum26gJljm5bRnUFauEp0fPtw012oInXb544e7UBFerHoXAkwFIFekjk2nuU5eIEIa
KZMhnkEzFuOpr83Nu8dNJuaBX7QZ4k6UOm+mprVKDoGmLHFS1eXNQlO6//E3WXZ9dwHEIB6s1vQM
hVSA215DqCVNdSyeoA78vlF+gHHOHmYkbtCSs0m68KEFsnc9qWHFVSd2UO7sAJR7t2smviuz7D34
cEogTJWnrf5SAL5UxCSlWQUZZHM9T6WTOvYoYq1JIuEFrkitXsocHeMXtjyjjQVUuO5TurbVOldE
8/8RaD9yTYvOJc0PpNqb2UEURAH3DHsRB4mRXSrvlRZ8E8LNG61tkdoBkBTHbapnQ0mKmeh+rpAS
CSuvcpyFzbfTAlk562IMBiiFoNNWWy2eQp1spcWyQ+jQPEm2tph/LPmlVSErw6/Sp1gNspt3GfoW
lZAH8Si5Q8p4SyomS3SQpaI6h4s4AB1vD/ahNctGXSgN1ZI9ZPunOOVe4BhpSfBILaUQJm1tpZQV
5JhWwDcNe8+H8UgA09iqah95V6wD228mgfi9hLaRG8Rej6PAvUhjGfw+9eky2CMqXCuM/v6KqE7E
7RxgSnfEnyT2NFvq6T8LkmtoZBOul5mD/YORj19WhLYrbaP6TRm/uZndhtlOGnNpvRNebZjMMwO3
QLJPZgaU7ztcXM1S7edLSyW/mVmiRgcLLCwR24BUN2dyMtR9zleL1dmAWGd8XrM98QxBASQ+kT1X
ZScMcEN4ICZX2PAEST+0n2KqBS1wLtRzSf1wu9mxeurEgqorcWYIFLwZvzct4Wn/MMJtNOL573k4
l7eDj9P9Mm+t8PoLnp+6hKErjZNxkA9wSuUnMYblUmOuJpiRTtGsMY2yKHtXyd2H4VYvKVwjhmKx
PIU6cvsLfbSc7UlHaooX5FH2ViYg/Fhwde5OfPwjnKvBE3dY4jKLr1u5TYlfT6Lz1nliGGYSX2e0
ac8MGiE/rZDcUHeFY3+r22vVNLhsun1UVTbcB5UKf7C/gN1Ok09hiMn8g1MQGY0TIqLc05ip/ucR
d/oFjyWxs4xalXdmf838vm7a+jg6nZjAmFd8meLN7cDC/KySQxUmXcdxB2QLAcfxUTAmm2AnNZK6
NzI6vf/jjGVGnepMeVN7Zeql+kXtl9ogLRcJjE09NQoTAfyrs7+ybhN97jyEEypyqq4nzKNFn82I
RpOrbMmRvygzsGLbFDUbGZu7joDleFxMSIWgil8f+JGNof21Vb6rq52B3V/lM1Hm2W3Q1VFWPIy+
MiZvYs25IZ6ltVZwuzlhwhGPuwDp/SHx647CJw6bw2Oaz7SkVg0gBS0qTsuFx0y+GEYaQgUIoAh/
LQTjTOvwPXu4YFR2qkV6iFiik7tYFDZDt96bmDNuzwNZ1jeVUC/DsKX4ouMz5iQ94woKDG/41aa+
7a9k7qYOcEFRAY0DNt45CX0KC/MgfhPxoVefrYBqr6FRZUwpY4hbB2khwH5ObTTiyTH0WdQIetqV
uQUi/9j9e2FaAZORcjwoEyLKVZX5jxq/5gGvy/pL2bnt+6fHK3BaslfBzrzprJ3AHrDzQFA8UbhW
3RpNsenUrAr8e8U8XpMXbGGW76ipOuh0PH/dOLVf313MJSf23dfqhsJmnJ6wTg1wVEmZVmGXHpy3
80DLpUdSLCmlTMjBJxyrvSNZbtBuXFnT7e9y/1dpdVRAn7RyvTIhAyaPtX6Q/sUzd8sCK8W5H8ak
UNWUOpl7yenwdeh8EtdTxyU5Y2PR9XRFyfnSOY4LOn+6C02D7wDR2U+RDEM+aPcuO1bBSq2dtraM
/vbjmwh2TFt7VBdmxy7OROTc3m6bkTT34/KREagRTuqkGyhkAw2Y/J6S5sr7YrnVAqZrl81FOugT
/buJEBfEtgwwfazgb4YBvlzei+/B69BTjrTpTo88OTCgA9c1qpf+S7uhZaInpHRnLD5vbsi1y7BJ
CI5Hy/5cE2Ikzy327hRBhERgIPcAq/aclQnf8JHRKfPVl3hmml/dQE3ckqyMygRONIZeWwvgRTtV
vSEpVU6v1D3ypHsGdjKt2bnYHCPNfWcqFX7L9PzLTecV4wI4RFO9osCo3dNm3QyttsCn2szQnxYw
UHdFYpq/g6kWw1gcBglcLSq2OCtS2x20ZPOGn22K1rXXLaibFAM0URdXxZwp0MRAv6X8qtv3Y5lE
Vgmz3RNn7vyilm75ssyrEBzMtvrZW2Kvc/opE+vdKOmaXtBPKIoB3Ute9ukJ3Jz6kibSEwZ/o9L4
0jg3Mty88yr5YmM0TK/z6P4WZ+p9uTE1MsBjk+bGXdUb0YCt11CtJMWmCvxVvlheRRcpOqEELB64
hPcbx7zCB2bjKDG7nxsvce5zB8cvdz2Crq+ypzQi/5PJVl2GTp+xKdPmSxwh1bOjZU/BGrMJpSYi
oVFyTMLZuWgcTki5+nCASS+HDUFxdOrAqfDSifXIFPTXpaVqVnT/gJKXr69ORlTeOais5H5qUCk2
Nt45dXN8vEhU0cBIYNLjSPloZNpIbd7dsJEMrEA0m6hdR6AdrdpX+3POxWiWB4OYNdl/HQvf91n0
Ju2rGOTduoKMFZRhYVFJQ3VglHaS8lzRGBLLlZvbF+TE92Rp01uasJAfY26a3NEActgzEDNPpTEJ
9AIpPRIis0oCgaO50nmKc/CNNrpf8IFO2hVs0DgC7QtA77oG8UwPsffd/4KSWUhkvWoD4EiYwAZS
uM575WvWACdv4hgb/op7lhzAG7vHLWTIndWKZqBomQfY0wiLJBmyaEx9KkEg5N7PXdeJo815frlx
3tph9Ik7t/qlu9FbbwmymNofZQDFZAThQJ1zfEj3Doj4u7tf5bGxKUHaBd5oIrT0jzx3ct41bQvt
gAl+XbnUMG9vR+GnkwMYx1Wu0EwqTy7/Euqxkx8BTwIE4gZWkDAEZikBcYvarDxPwjD1VPoxMQ6p
dWv4ij6V1+X7uNXAZw5k3SSyInrLpRyABXk67ZKCtHwH4jDbechPcr3sVPFxKR2PZMWgEUEREW+o
b1BuKFPlg2S2EiGnFLfnINyTlqsbh2Pz0/Kdz5j4q6JlYyhEC83LLo9ExedjfDOYUxbMtxLqc0lj
QVr9ChLFP7XSUnDczYUOfkQZFSDt+8THMyMbta0kADSZ4A/WTyl9PxPdyHkfO34v1i2p65ZZfc9y
m7U6qwa7Djvm37oDD6wkbN67SRAJgS/PNmFFH+HriuDLxUw0dXNBVZf5GiuRd3Jh9x2p0B63GV/K
OjjpEUGCMem1VodwSGw7+0gH4DcVLz0yOtsBoqftBcKhWumQUHTQS1rqsmMJ0oxmdEf3WOJAhzdX
me0nquOuTsq/GYOOKqIzYgQf60FR1dnIOwT237NmOCfIHRenlREJgYjHeK6EZExAkFHNTrADwo+u
/383vYQyyI6MEP9JNJ0+4rYzc9wpS6w35vEosGFD4BBVY1t/Lp1szWawbB9UyjBwpIg4InNCjqRQ
ULAt+uNE4zZ2FB8dM92mRv0FwaEQDsy4jHwSIKuTm84H4aKBIhwUyD3DZw6m25sR+yByibjzhLoc
5JLEe6WkVqOGcGdpEfZM4qKL1d03KZvzh1uv5Paj/yVUKPiCDoI+Z4UWmNo7H+alPe9ReIsMDYwm
q2hAt17w1oWUpWIlHRztMvR51RWfzKJbIBL3f9hgEKVL2HLxOFfU50lRshvLXDQBoGtRAmIK1nCv
v17apyd7EOp8xi6zKXa4hdX/TcuNdnZdgcOmKYCaLw84qYQierW83/cyXc6ajtiHvYP0tFpn3COK
vTXIA9KefF8xiRQMR/l0Hrk+jpFhJfYyAiBwrxzkD8pSPuzaCoJV03cJM+ibnfL8H+kJQOxw25aY
d8pYB8O+ME1tc938yLv2c/jmARBOv+MrSdZbwx+7hdTJEpcteXLtdKsD4MYtf3kTqQN7oJodMXFM
zoUIm7lyOfWKr9TAvbaUUP4U74qSB+lfDStuwJDPmAQVsC9jc6lRt6yf2Ec8mGheVQx7idqJblTt
BzxznjPGI+M5aRRojN9ZzD8coSe8UTdiqTtmDkt/2xKf7J4ijz4mvNoF+FKqZ38kNHXlfZNNoiOU
Ks2uAoM2SGxZD1cuWHORDiFpa12/JZON6od2eyKSaR/FoXeMjZaaFycXGd6/4rPWOk+fT0MgMKU4
r8KW71T36Ihe/iMdFGaBthkony9VEjaXlVY53TzRmJ8OzGmptwktEujbTblHc5M2A77F+Mtl8nTj
AXLwv66yET34MN7VrW8t94C9fO/VBThBkSDc8wicV83PgEqoeLQd1EKk5yfSLlc3GwH6O78OM8QK
cOJO/lKEuj9GI3n4cIw77OLe+ZMV366NflSuJaZ3zEfFreVLJ2bDUtoqtDQmblabfbyMbThO/HVF
uF1cdZHHopAo/L96gtAQrPaXMjT7Y6+1hZRyz08s91E0y6d3Mbx2PusXbUHeMFlsT/xqfj20+bje
4utWlsr7hyybxRRbuUzth1vJxpd7bskxAXbKtoxkon5fdakfv91SyIAaijw1KxFD8DLNGVsR2P5T
4u3sssRgRWb6Kn8ReDuxLOaqD/kp0zRCGodVKyxNnKptOgE0Sx1x910lqnIHSMgBRFO0CbRJE5y1
Z7PV4dQpuGJ3mGDqpos90bgdnw0EJWTEbR/E1jNeG/gwxf4NakqG5d8bdqRuZ4dMMn0s7i6qLdUA
EemMGgHg70yGD50pQqUHRnchXzn5Tv0f6DmVx3oz2DJCyGyQyuCcmeosQZk1yRVUA5JCS85KO8wR
Lxtmxhx2YeRpsE2outVe+tDethRCvZ46OPvf5+qPknBz53Yj5rUt5KvduZXRxWlDpq7GsDQeu2Be
J3RT7RIe9mBfzTtLaEocTp3kuksAQXuOyQNVhWS7YjJgGz9L5OLhPmVKOI8rKFu6OBNjEdaxbUdJ
LLi9sRxrLATAiSziqY0wCmXNu4dJVzZ75HvsSLCkcxEBO384r0qpBY3NvP2TNBBNE3pavKiEuiPF
ox7Iq3it9ngC+pNMf809qFzz2xW5AyXU7ZFym8gB2cQkkMZeGRQYyzXoJB2BjXLSv3IsThWYPOAZ
YfPf/ZnTC7X1UeLX1w+UBuSv+EoQHHDKIiZcT+ZSPj03Bz10qM8FHiqxfDOM99IulvBKpXSr2umI
5BUVC4aYboexpegcr4y+Z6n2Q00anJ4L8dXNw2b0SebYcGLn59rEN7xOfuTkUtp0AtlUAJWPZDG/
BXD+HFFYZ6xvlItHAGJznvSDa2a7WRsX0+O7gD5aJUrizvwlGlzyMeebUaQSgEYivrMrCO0VvwLK
/yiy5+6uwHqBV2JMQKUnQfTp7TayRJ27B92fuCXnWxm7CHg2Gru3zJuXfhdThUz1qliJDzYj1Y1Z
JbQgBExPrRpFLad+lE1XXgbq1b5J0K28VzLnlRi2c9+ssU2ZcJtt3C1VUN7rLso3pDD9DeHCUcio
qtxJvfRm9O4gGfjxOwN6aGTN3RwWuOOaEU+T8rdFKFzIjQ69hJZFJut4E1hfBjDZHmeTfQyTTovs
qahp1NgL7bxMY/EIdDrHHou+f64e4GGKqUqu8WoK6jbBZ2QsyWFDAzB0W/lXo7BIHirTyiZqwjtb
lZMExJKOYCQTy8gQ84JSkZstbwkFHWQR9eoEuRrCAtcvAvRYhTfkGyfciXxGg4dGI+mU9/tdbo8U
XhATuMpQzhzgCSjeihTdp0iKovV6jnX9pAldgxdEnWWUdjP2yIKcE3pMcX+lfX9ozKWUZxYXvMlO
CyVuGQdYuff2mAzHqq0z2JfJtoXXphB7eSfVVRFigNlZbZyTYZZwdwN4I1DJE3lXIGjbQw93Gwcs
3LH3Bkkk4XkPPFD8Lq8ewz7MbWkxietUKl5Kd/g6XLpKchRa1uoBhiTt4rGVFURC6QZsgkoocs4a
3ivEKm/ZvA0Ln1MoOlGSYiJBVi7E7BlR19bXm2xWns+Mu3QL1Un0DMyxhgaAWX5YZcwLOUL2ZvyZ
QPIN5+DF5RzuQ6hbnUhOPWBsVK0iLbnq5xyqCgJjTVH3m7Z0Yz0H9U8q5FjdGY+azjl3G1YxMwv2
fawoTSfHJ+hN6KR6mf8cszM4b8AZvdHNyx0rJnF4cKq3tQUlZOU4wl0sY6gnj8NiWUltJt9JQnAP
rtwpwgmZmdajD2396/v+8sS02J5LL+9iZg3MSe75ArlGRPon6EEWVRqBzklmL8l4TGpSQNVltsoi
YNPWbOZgcEF3fxxGB8iasVUoxlJK6c0bJJSY6iRuGrS9t4YincINAzvXM95DsLT8leCS18RVuKNL
31JXpZ327vpmtyNgU1mRvGEv7RBJdQB0/bDlGC41kIjR82+Q8VhNcizsHdGS3wzSSOv19hGL4Yiq
CxEivLzh+t0B/VRWxYuRPfmV15Hhqs1hNdve9Oa9xOp7ZifZvn79vVcwt8mEfibjrq/gjRLOwoXs
BSfMXoZOaFQz6Lu9GCp1efA8kztNr6FctbX6cuD0Q+tY1qarvVyYQjdQnCyjmQITWigHEAjXXlj6
kUn855YrOJVpYS/70VysDA362Y3ut5L4zqGlsMKqZdEXSbdkYTq0sEZYNZay85GqirZppr6/m3Rj
DOGN6Xw0zobD0pGIPT5gbToyGsrP3fczD62n9Tkww8FGZLXZuReqNqUdzVeePd7/ZgW15MUc1Lrv
YuNFjhp8cULX62+ZA3GhGOWHy69P6h/f34l4iFLISCWfHpU8oD5V8JENQ7v6ZCEfr+TrV3/MwyP9
3oC9fUNXRbs80Sb9xDLDMynRhnkxQBdNng18Ern2eFnuLhP0tZzVn6obK/W+X7uS5869OWVydHMz
iB5Lpy55YQmfFkiIpi1jqD2BDjLNTiZNw9QQHbyig/eSAbYpFP7IPLMS6MZP8VA4e/3PhtXI/hut
pmvyaI59mI3nhRSqGwBSO65qv+od2r3fhZ1wyfuUnVyI+vVN6VUeXXpqy7lKfECJTdllsUPPRSkw
8EZ1h6BcwAtxyNPj62mFEO+fAZU7xo4mTFrEIS8hdk8B8wJsYJhsyy39m1SoDUCvGIg5Y5dhkUIP
PWuomEUwJNAu34tlI6OmBICp0lATqlbtg3KzAnsp2WUkWMun4Wx69ol/WXmHW/n2DX/TXxJ1p8C1
CLcw52gxudKzAdFUsVOGL63CUvDcp4k15fxk+x35MyEQp8L1L0m946Zb5y1TXXhLUJJkBSnAxkaL
YmqPQKI6qkqcZTdYdATzF5FORaSvLdso3Ll9YvwbrZZ19pElnJXubuwWNflZpOxarSvVsD9/LXs5
s4JYVtmld8Nxv5j4e/7zsNUmiZ0qVJP29z940+X+VOxHXDTMUhKWE5T75mGhLUUqxd6MASI7R/hc
+58V2Q/pcOMRyQ6B8lXbhhzin8AnFreu+9MJFkUpqyKlRTRyZJ5QWV1sESHpbB9Cv85p1nsos3Bg
r8ut8A8QUfS0yp/ak5vjyCb0p2s+rjoO9SadoaJmMa70xlLUnovcOI/cQcy9awwnd7RiyyiZQ+tX
/2I4GOxdoRlCRQg6RbF/600k51UoZH474BIxt/xdzMSXX36kxtX8f4K+sISDuSQ5usvnyE6OHwwo
lr6ay7w+xtPF4rnxpfeolvlGHm55Qd2DxthO/wi3voRRNvLLEjG/Ht6tS1eVcGpgdP9x48m6EGrt
W365jf9fuGcY32Y7F/4QXLFOb2NP1AYRSBQFGTaU50FJLQjt7QuWkXFynoRxPlX3oPJbLr0NJInm
rBkXcnoEiGhilraC10faZBgPOUZ2cscZilstNkp+vh0xUGj2nXydwSLMWvYPKGvEnJm6AAvWGAMr
S7iaqzoyJS1FmNMH97x6MAp0Mp8fctAOI/2K7x4EhclGRwzZJDkzks/Gs4NWOtwSmUSSdnv+ufG3
zKLwEj4yD/k1njVsY64miiT5US/UroT4H9WJDtr/qFvXB4wofvxBSQMbsEqj6JrVHtpLEfhACj5G
qCRKfRsyQztFgvlrzOmOqWd1U4oRDErQALq+k4WhRBBEpu6Qsqa/2Afa7wiplRbfvb0QxEXrmLKL
HJKF62h/EhiStBb+Y0zAB3Q3JFCtD12h4f6HHsQuTwakeBP6+6NY+hzfF8+Kv+9jToKOCmSo+0cy
01J6zy+eIGJ0bQk+SUUOHpgZ7AjIzjRaYUiZknDJvqjNQoUW8ldQqRz9Mu6Re9a/QFHLZXqi9dhp
eCsivJRC1+X5GW8By65jj7Tw03TP6TeFSOKW0B0Ys3FFCE/DlquzZiuYUoLNjsdBfkFN/oC83Qyu
0SoYTuANhvazrh/O58psw5oesv51x4FxAnnVKWOOgT5Bp+qMV7rrZpRxUaQfKz2yKlNxxbn7vl6G
6TOf+BWdgTcU6wMyhlhEB49Glru6yZkUwPmkQ+1sFNZgMBOuzewwUiG4I1VKAVaKfUC5LPK+xwQq
sxlIfJc8tUrAKMPzrhOZFBzhPy0ccVyC/+Y156X6fchI0j9DehJG/97fouNdFfnSCdKnKmy77AqM
4b5YGPJqhkcLa0sq7LYVeJqQrTBPQDcbkjIqotxf62Qrkupp97dFl6JpWNSS1/xZwmJ5ckTh68/a
5cHUuXAeX+qpH+TgaBxXSEpTKnOiA90s7ApSTdjD+gpS8GJCnYYSFFvQECgZKbjwUc6Ap5GDNSJt
4OJxN5xN3Pi44grEhCuN8RSYrUQIUgaC6jlKWCbAIOw6d3OB65VWBeMYyMTc+WpPP0dnUd5vQPLz
nQRmQcKMrbP24flq5qAcUnuHwx1OR1e52D1ZmgL/gqOfyyAd5SM+bFWkjd+3rCVdeCB5pvuvmF7g
mb6r+Gb5n7mb7NoaMtuw0/vkkE5SrEmbhZyxRGCYGP9D0Iq96wudOWocJNaSvwXPDRyUOx+cxEWn
eOyO9bl4GYTCHPH0zVH2OpDbyE0ePliIjtSvQSgAW8EG2aP48iL03WqBE4UiBjk3T+3VYXdG5f4U
3t/r2PlwM0X3ktPwJXPNKYvqtKZ+P6jS227K0DmTIgpy8xbkbux/kh4vS5x9p6eWnLFg4TPzzbwr
UIWls8vTmqaeGf199nhKy1nMxrfFfDugK8hoq8HTNYtXVvLHuk6ZAxVQDolE3bbGpjXt+XhDn2uf
4UPDRDFggTWe34VYv3FaNGAkHmoKd+bCIkPuwWP3n2IeYPuXD+mO56nLov1Gj2GmTyAkCBrC4cCs
TvomLEUxy1VgUksiGe0aaOqk73MuoDQwfWiGLqP5b9Wbssnw028zbby8cp3hOToDHrxjND5bQD+Y
9n6k7hABhrnGj/IAywH9Q+/ODDYuGACKdEQsCBmXQdYrxfghlu2W3fFMxl6NuXrl1A/BrJCWl/th
Cnkrhwce1Kt3VdBVO2zK4rT3QBvMRi9XaCeC6qDwQiKIDqlW6BGO8XBRtl66sLiVCVOedUBWI8rp
2kU8JVGOnVhSvgyaCNKNcR6x8ySkJc70EUpCAyOi7B3EmFRD7RKm1IjpKs7dxr1j2DvAfs5kLA9X
z62Nn/SRKya90PHIFSuFnuLaqjXIY8RjmSIRI0b5m904BOxVSkcUSMoGtMpPu2W3rEUnJcb/GP8y
cjPipQzbB1UHZ2WIhWUrLAm68efVrSM2E4gTuEOB6seg/ShkNJWwuiUkO5PpE01QU+NI36fov4/M
VK4JwMnc7/f41g3NH9UOL03UO2DUgGFXnLSCsx8QXFWqEU7Ta1jetTcbQVlW+x+/YFZ3zE+42ldT
Ve16bcEMPWRiPbWzQ6t7y2G+HN7FHY5+POH7eaRi2y3otgPDN9hNVSoN+C96DGhxpUdhQR+0qJX3
Y5KZdKaGbkXT5zeqba1AntMQOk6IA6IyGvBdnzrOKmnw9NcwJRYvtGl/MMTXlmOPXffn6yJGdXtM
jhlnnO94WLnglPdEcOiBd6VD5cIeQyEVFg82sO7KBntQsCD7+VALvX8ICRL2tX1oCkOtwmsxse0E
3wos2hXqUxROvXIHRy1nncgtsuVlA3CitYWbM901OFQvVesnOJ9xY/C8oT/PzuqPGY52z2UAgmc7
2mgScNVNTSXvpMeFIw7LDtSYMxiXABiPCD8A/+ECHWEhEZy/xRGh0KfZJrGmrDakYqVBnYLfzmkp
6I1WQm/cJfYReiURMXu++sjblBq16Z8F1enQwTBid5tebLLDlwIqcHHYVSUBh3vgS9hxQwa9ULqz
R9FoyFfBo2wWQKHxoYG6ppNVcN9LsXUyPmc3/6uiOySp/eHv/TSChMGNozh9hLt5htzG46jaC/rV
PT2VeYZPizj2dxPMfEqbETRdWqH4eUSqaPxfMUEnoxNKiUBELBueQnkBf/QBd82Y+jBNTgZ4fM8n
IQSxu0LkkfLwt1lKfRbuwgFsJHnLL3SII5tG/TcK+/wF7bMt3fvIEUGdOYd094xxiKrIkZSSVONp
eUPlBtZwU3vRQh/vVsaGiZqQAGCt9mO6I9f2T0+jtrisV7D62RfCtE5inZeQPjEU9gs1gr/l29FO
qpVlvmFVkRjWOcj7wfNmfm8maaYBfSba4LATh0oYCClWe8KJYebh3g/dORC0uc7FKMFjqEjMutVi
Vj8NJFNU5hI5VBRh9QLT8wW6ZFypy7yPzEC/mbFK6H8sk66hKbZcFkQjCBVi+EbLCACal013093Z
tNcTI8xQ9tg13d1JtFg4hIsxyWNDnim47UOstGijVU02cGf9AQ1iGyITJCpz/GtMCKS+lkJIXk3S
3O18lRHt1uxeXtL8r07nzE8GHAg6
`protect end_protected
