`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
S0Z5K+NBYWAdvRysItZc8oqkqICKRRUYpiXa+0/cK10j66PXzUB2Ka5ZZwtCmVF2r6koVA1j+NWG
zTGfRVXEvIaES5DGRcwvPycGte91SaMkzZNvrxSOU509xWx2YXZWqvHhzmUp/X8CaRyRmZ9DjHab
BJevvEifeTpPCjQiSXiMxQFQV+RN7wp8fzNRTkOWOLGf8EFXbXBkGGO+Y67HUK6jOY2i8Dp2kOKE
Eu6sWszS21WkKLftsqYPWjrdL/OlJrEDt6J2eP2uUyWb7SbWpUeQpwTOPiSnqQXytsXwqj64nSGw
RPyXDyUymScmBRH39e8akHiWAAOMkTWp0HBwpQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="0kH3KSVm9sQHjARPhtl2SGQD+lu4EP8vrLfnb7fCPqU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11648)
`protect data_block
8TS/1+F3WckJuOUN6nn/dLDG/ikBXK45C/17KzwGaercKkbViFahBHFaOWuQ7n1hd05s5/FvkpDH
8VuXxWLmyvQ1vSRSwCFHz7+jHYGxgDvix36d+i9zE5a+CttxyRT0rTEYphrIuu5qB+8+CHc2zcUP
Nnshb9GaNnnxJ0jPMTJEhyaIKlUeZ+TFPAdbw1v1L2ZYoFH/2rVNd4jxihkHN45M9FV8Ny2juJVO
JEdZkiyVkHLAaTC8uGzBWMAUXfS5RPt9J2Sa5BivNWk/UuDqSJKe8dNRul2fnQdCKOTuV0AQ9Jqm
noechgKmurIRNiE533KFLoBUw9mO5t7nDnhYKxqGM53cFA4cy8Q+15lJ3H2ebiXdOWP1uqPZpR4d
VEZLFJFkA7lC9HoJFtYqJdCC4OhB7tEBhW5gYooJnTeImedO/oYAr1sc52ni5TReTYqT4VcKpAow
2tA4p9Ucx06Q9n1ypl+2GtocrFniOR+mR1jKP/rnijO8wFfdpCRGJh0UiKJQMOSW9+kE8CKEn/g8
Y/TL3RUOtwbFh0EeObmXnptnUFNA5qQzryGTpf+tav6YF4xhgi3YCOfHKaeZhYg8bvFb+c4M9RkU
zGlQQprwtF845qXxTFXQI53t83op3dnh+eGhCUbGs8HiICYWYFPELCukYCU26CIiEMfZN/i0Pbuu
hw88J1zYxOExG1aiR6czt1QxHn2DsxF3dEV+sP3YxJFAc49LTvJBMATRNUGeZ8pqIR891dYNuXMa
hkd0noknqHZydh9ZiarNGsRN2zORGcn68DDjrz4bC4dl+3+pDveYgJIedSywJiWI99D3AYX2yQ7T
5gwMJ0XWKUy7deWWOPKP+RQZFWWJj4IFuumlVJ3sUKSWHlVD7Xt5GuEksnPnitKCff7ICFeT0JXj
ikpGeFRYHryJu9WyEZtV7nr3e+ey4UYtlQ1R5MehKcLmuF9e1G6gHabJg077c6I6N3XtWubMn9cm
yNNH0wy9mtNqJ3WBa1WYXesDG/knv6OLHSG0cHOcxVxZXxuZH1eNwdcO0uQM0/h8pGvvg2ug3vO3
RaLyu64veJDEG+cXURNqz9N5VTlyBwUb/wvf461YBNs1/5G16pCkBDb0UnLhd+byvLEfxkWTHhHB
vptBVgQR6tMzHJNop2EG7Tnt0lhSfP1lRZAHI+16DRo5X/QYq45jKujVgNCLzbtu7m0npbA4XWVZ
kVDm2p8uQDdrPXGw5+MhTxixCt5XkIOIb6W8NO+gDBa2/fHELbakZLmICF9q0ff+9faiHSJiPgo+
iQ5a9BVrEK6bP7AJtlDaXFLBi73tAkVX3sLZX2IfF+GsTI9KnW5VGmjgvRNrBjA0fFz35EIdjulI
6qj/HmGsdDw8DT3sQZsOxMsYy7h2OOqFtllGXUJ44Iij/oQIU/6Om2zpHtt7yMYR6S/KPtr3uNlM
4vFun7rvl3iHlGAkn2F5ySXERhoA4N1k+cKm6gMLaKnX2xlDkLIQMyNFoNIypvedAnWwnn/wiiZr
HxFGofUikdBF/rqXryl4pkn4hYRQAaGaKdxqsIjsltk6IjW9ouk1xttGQNLHlgHUWR6RNMEqz1dd
7x7L1esP5e9s5+/qGP49Nv9FVuGbFgQIr3xfFAPFA/WYAALkt7kKw6QZ2i5iWZTIKR7uEY4TDNAd
VOPZ+vmmic7pColOSi4ytCepDwAC5AdAFMwCiz1r6z24Pons0KMxFj6pJHzZIvAeeGiGeQOUIQHE
pA5X1uxDsSRdm4oQRXR2ZvyJL30HmQs4fXXv78IYh42q5/zoC6bNONHwPcMkKZamATjzKNv5T8F8
xaswuKB1FNuEwJB25oLHzbnsZmewIVqXEnRMG+TosTL04tMmgFkX9kXpgQqmQqaM6s9BMsWL36Fs
3vriOapts+3veqmOa7MRD2O1Lti7J3qSWXYHh6EULGoaOrUNbH+GcjCaKCvcprpqK2PfcKhFc8xl
Wv7k+NsBsWL5kMtJYWJ7W+hBLZ7cjG4Vh3vP4D2ZfcPFPnXQLIeYXt0lySbGCrxnDS5P7E7hAsos
2rNi9/XUXgA3dDLNSAJSQTbAlsRdE82V9v8Uf/lXtlFQl26RLPVLd8okFMy1cVBk5pgH1nl1rs6z
fSozgurzBkUKv22VXHsGGCEorgQWae/LntdJ0FMdpTSd4LUE2zSvET1WgzpvKfU2nX2XluQY/Wb0
S0Y9UVM7Nd009wcc8UIRtipbHV0oouCXpWWx1fXBjqXg0PiQ1hPJytngkCnEx8NQBl9a9N8OAmn8
VfafcjMy4oyR9PTGzwxu9tjF1M/UKbzlSL2L03cW92gfazq2SYTzgnHeMg9tvJIsXVeGrzumDoUY
NsAc0GuS5WDd97+NaLjpjKQqq7f0JWn3sLEvICllW2FImz+VhBqOr3Cb+zZsnEDNSxW81pBYMbYL
+O8uKAZoCQwlXjG995URpuffWuMaJvFMlbS26sJwZrdbYxa2OqthGZjoFS2v0f4is+yW0c/mfzIf
Btxw3I58y5ZGFRLEqtShtxXpfazEVHQT4j83baQYDBy5xX7RbMcRDqaJjeD1w9LbCNs2sebbGIRk
35oXrkW9/nNjvD4Lf3KD0KCpVyNT9dvNo5tQAaibxKUE/RdXB18q1s9FSP19RnnHBX+BzPUFKL+q
lDk/nVtnAlY1pVIRdFewYSfkOb7ALU+OoShg5uEdu+Xzfg+dUkgiZVT1QyEf4MyT7QryLzuSPtmd
MtyTIBcXZLwBb0W6MSMjd5qJ/EvLOxfXTYaLsXq0mdwO3ezMBm7ilcJdmeazumQ6Kfe9B2WWETnG
I+o1g0IyciYVff6MNvuazpcsDvBxx5XamnhJDAHXFGpdp4Vp0+K0bCtCg4Wee8ANxNyVaotSSk86
DL2mfpUA1qahT2q6pJf9lH0nxHk/amoY5h/PO6vdBwhS6GqPGo2ZOAoN2eshoKHH6ET/W/ONpp0u
cCNEtU8XuXElwm3uBxBpxqvnQGEbfYQKD97qobCJ8ZW8N6P4+tiv69p1KXP+r+IQE1Jz5ahdIVC5
lz39sCIF/x5ZqKZ6xCyYovBUuHTbdFFfsv5jnKuuROzKIdmN9b3GSGEn+qFHfwDmK++1eF0F+2V3
csDwFlfhOREhl+tVE7oEXMalYyV1Y2p+8LZOO1YAyP8czuKdRl6Pz76+rfbkWK22aVuak79x283v
7yZ4AFFBVCHfkClkIWmk0Z0jrrkZzdqNvh0OE0elhPmUMYtHwh6LBsvC8El5raHKZsUSCK14ZCG9
ybpjASSrV17UoGVIwp45RZsRzxeeW6fdilXwQiDptr2FETfyIh8TeJi/3aOEYr5wqcS8oa6id+YI
nEOze+5IU17ceoqMlUG8wkI0fL/swhpAAHpKJMhdsMwHOj2Z4P7qGQ5ndo8/rHa3Ev+OhRBJz2/w
GGrwmkFpkGP0P43b9RAhcgYoRGEJu19aGG+PuoXGUYjI1L0gL8rjCk9Y5yOdHong2zQ6gEKi2GPJ
2/71LUVKBM19c4GleVR+0LJKf7X4J/04bOkahrPeJ8EV6hEfyIFeZJ2GjgW56lpDTIkvlY0dXjyB
GLw14cMVyPdCrxkW4iIe0SKg/QGRKKLVkdVW3DnpwKU1mJR1Z3Oh6Q60EdoJ6VWA1kp19Tv5QXE/
nBdaXdaUAiiGrStS1JhX7ncUfWoXE3plXWNYqCei3WBZkhBwpYfsnqdQ9mAAfPtG7C899mjt2B9P
hxxnh5a49ua3YeufDu3U+/PNV7Ie2DSbdf7T6036tmd8aabxr57QEhSjVZcL/Hiy7Nxr67x1rB+N
bPI/pe7ZEhZ/m4FgJqd5Q8f/WZ8EkKRcXUsqBNCcmBVyIhEBwYxlTX50Lo8BfEelW2KNl4S9VfwM
ZhT3v3CKD6Vx/ghb0S0VuADbufpEiDh+O4AlJmfqQk3o8q7tx4VB4YK0wROIW2Tjqhch58KsA//E
6MCaXgx6fKfLfnrxMU5gyCtiHK7o2yFJywVrg5c+oTgNGBPGVE//hCXbXeXSEpKRF1YK0FrtuZZP
Zlgu3I7mIYLVwB3ijINHI8CYWGwswXoUg1yXgLgvxzes2iJr1dD/6JTK6+o3s3PpdIcD6BgnXXJI
HEBEh8JYfIZ2FMp3kJ7fuUgQ6FRfGfU5/iK7BT+qwksgIFAsB/tyt6dxsPdETDp7ZSsp7fVFsaav
bcu3R775FzIOQNCUo1IUZQmUNZ83/8GLxQxNt3Me5D0NqBWNu0ar9gZFcqLydc0mV1Z11NX/ymYy
RQcwnUGeCidvuief/fd7G6OZ04N4bNChN8FbEPUdz9wgaI7Q/Y7U0XvPg0Q6uxNk2tB6e69yJX6E
TAoY48qAZucTec0zIbpizBjpgJE6rDaVeKanBHOiTXCagYvFjTiolNPREyzAaQr+N8+RMz8gg1Js
/C/Oh7jrl48jPzPOhUFZ8wyzsTl/qPEaah75Ncoa4XViLMLs/1Tdq7thfQOl1CyFncmTu3LQ8lEo
u2cLIMv7OR47xDL/BGPu21FHfOhR14SDov1qd8T0dtlzn0Se0lS5T5VJgE4BGpIqLMB9jzAS8nGc
RZDn6Q3May6qgLXirqY03xfRg0DmBwADRv78BK1jkMD4I/zbci6Jzyi7WMJboFW/gE6IBxYhgJUP
HOu27CaekyeXZGJ21kR+TEMsGgKBibhuNYoSHs5HiqVr6dtZSE8YFtNzwht4lo9CTI5lAoD+TfIp
XQiTKEcmpUstHAW68rnz4T4YLeYbF9RnbiZSKFXisTJfD0SzoOfAse8wTkG+HIDPS8NzyBs8xdeW
17woPD9dMftC0WW74gQ66Nc/7Y8vtHweT20I4lfJSz+96MH6MgT5cdhIYZJUoI7NqqPWiAFvNNql
JtgyUlzHyCRBuMtGNF8Xc3ewMUI2WA/O3smjPsTq4VGW3TGpkvDsmP3cnnWpFq8j0e3DeHDcgnr0
NSjamwxE3ylXxz25ott153REOspFAklqqSnc28SVQOO+hKNgQs3ONYBO7KJ91nGGqCGEPPbL/suH
tuIkZnVXRqcclgJJri97N+xHuMXWqrG52FO9V9wzjWFDBaQr+GwzdyAWhacG6MI56zey06albmdS
FLiUdRufl8IQOBmwVRGXLFb/4+0HsdEb89duqzjzNZmLK+V/VQvzJrD9KoPpl8UeoPflbq6e42pC
GtVH8mmkC8OKQ3qkndtm0k7TsjptQgBkSRthrwxk2pk+BILerWGkk+887w544TPN32ahF3gGH52W
1mEsQnbYAsl898ojoPRvkccH5aj6d84n9Rr8To3uOus0h1G7Sv5PCxI6w9SDe3M7VDIBOP3W0MTh
EVJL+HktHEsh8Ves1c+F6nBnJnABCmvtFQCnyRqj5ZOcgrqR5CXhlh6Yu82pywtDsRGprtmvXDS3
4R7QEtBEGni5hnrtoxthYkUb5JUqC5Z0sMltCHypFgoSyiLwkGwD20GhuLf/btyr+sXMsSX5EeJ2
FzkPIq8L6S3KWqPhwra2NfptPJJBq2m0bjKKFaeTLOm8IhjYSkHpt0Cygw/a3Bh7uabNJmESpGPK
ELsuJI2WKLDyBOVFfwFydshkgxaQxBAsxtpsCWlQ3SiFG0luqOBAce3ByJUaBkgfNaUuipoyFhmC
c1Y5SIXFMokaiyWm0DgJJX2joMgnD8ArI/hFD+Nt+dmKHvvReBZKpKJ4sCFOjtjv7UiFk+F6F2aG
oiHZ93Q+zzVgckEecqvicijfNIG7ojSBmlKt5+siU3NFRFYrbwpVTvZo33nm/AhypwhKGqeVN0JA
7U5nJdviIJ5b+ZvsM7na0Q82NvxXEavKrM4k700FBSBs4fdhi120C6TldlDrYxSQ+tvl0kQISFN/
5uRsjM7+YvzV/5hG6mfWI134prc+8XUiPlzdGU6K/EJOo0WJIxmpLBukSo1/ZX341n27WYF4pkJN
M5Zd4HGdq7LypLQbmYeSqCW9Sf2d9BcT5tyJuY80ROxsJfLTEbnFB0Mv4EsvGZNIhmruXE4mejxN
dsecmzRO62kiIGGNLNZHhwX22SmFv4VOkxvDYMOR+A7exUI/4LFLu+sPHovT3pEdGGrjToVq428C
eLhTPOH95DQVg3JA/YEo+GH0HhrVZCg7k8IiyKWbzzuR3XOtCY671KNWHGjpe1PtBy5mSxbgQypI
5BMg1RgHHuSS4c063suRCm/DV5h2+zOwUBSDAGteBUC4XFUSJdiVFMStVMwzrJ/mN0uUFmtcwV6e
f2kU12gfZ1zvOpTrmM16VTcW5Hmw5kkEPqTKXzlHL1octeXPDGzCiZrbHcCQZc93CRVDYvcStXbj
+xcx+QH1EM4Q/myjP5z5C8Mt9dzssuAtxcWsfYdDtzLBYi+2SP31tp+SfLKLFiYX3glkKeDAUn09
V5325iMO9vUOXFDCIpWFBmehPoFSEr6/yzv5xVXjUAjxHJvHiU3IRNlIwWFOoeHoigDm0SN9srF/
dprO2sH6vxEB5mq/HGn7TCdImOkXokrJRELVyYTbsNJ5TDGWYJ3jLJ+w8yxN4Mu26/3jGR2PL973
U3Huin6Ka1sMLicg3wu16Bqaf5+yr+3YtpIIKeOgFBVFS3QELIfVQl+FAW/oZZIUjOH5+GAdPEFb
RgzJEVhf5H2a8sikVitmu88QoiFeschjEAiis3ADo022LxmJnu4X4YxxNDVvblxTwY/JPdo1M6Z+
wJlFDds9UZ5TFmUsV6J3ALWCiNA/m47zMT25OFYWYzSLm7/J+xK/8C1dAWY+qjUK20vFZIm0lqyj
HyLe0TWp0CAd2cd8miQNrJmebEkdHHBUdaXbBmsl3qS/bz6Cx6PwppHLCgMMUjvdzDoKcW+IIfiH
dRiWUTSv/o4fBKvCgVd6ByUu6CkPbbv95Y557BQVEMPyN8S5FQTYmVJ1aLjjwC/Vxo8xjgDQF00J
pCqHkMXQ4GSQf2put6eEGgzx/q7tL5DM9EfY4zFll9v8z0ezLK0oa8TsE8LVRv5M7ZOljg01N+0T
wNZ+ESczM8ULpb2RAeY1KbbGjWxgpVwoTJ8gLNUJ86mBipVVNMJ9itVcdt0hlvf4bY6UHOR82IgR
PEpGUQmrKOQ/rvE/MgmKMMI/uY9rQ58+P3+p3/4sj/yB0TU/UxH8EF/sIEQ+9tZoVFTUE2ml3ydq
1f4auCMQMwACMlcrl0qQ23UHZV9wy1SK5WGCc6rTslCxbbMtxfltr9CbbWk5m0KJpRBIEAC/86yb
l0wFAb/U+CNaVa9P0QvMeaCNXA8WDld2BHsTIls/87OrArdkkO7wRW6/DuORWa3Na4PKaYnndtf+
G0BftvEgoyScZEd4gap/DRQ6XRxvb9kZTBDKkpXDZOZCudXjkvzCndsPqgkmf81s38V/ept5r87m
AEVyWyJYpw89s1lYl0V5dfLZSjrKKZdMpuQy5u3gRLsF6mkCbklPNJj1b3w7H2INB5sMclaSWo/f
xI4aYEp7lIUqZ9MsXfXHGRGMmnR2eMHVP826fTaS4h+0+8bTDGmKkgzka7sWMKx9zvnA/RCw/KAA
uAGQnk59AH06q/ejHV814khNZThOxScoFbrqr2Bf+keBHzf65HS0+ODW0iHdoneyH/sncrV1NUyx
ebgIX0Vklstik417c2e09YbMnpk5H6YNmhRGvs0jT8Xcjfl5bFvz53hnSQLk+qGl3LqgSSnJ0Ufp
47JeS+lgQHDhFaq6h2JY9vqK2mQHOwTHIMygD8U/uthx1qADQB0BoHXoIjfTMJat1Dfjgo4HfnEZ
9lQR+dLQszCZiggmw1KjwpbkaewgvEgv0U0Si0l2OEutmKTXOQzKgbKmBYcG18/4RtUgcFO+kQ/B
0CqF4MhPMXzSib4OiImUbf10NO6/5sK8tTdDBWV8OufvUQtqsUD4f7UQk2uJKKLbm59cf3+qq1PY
DcVsw+pw6dZVJ47844fDxgm/FOjQDhimnU9Z9Ws4uVug0bgOU2ATeZup9p7W4wZ1NlZ0CZ0vsgFM
kqBuWU3ecID5gYKwnD5NRa7nE4+INaAjI5sM8XiinS16LcSL+j1kXmMQ7eQnq7dEZE80wUcLatZ9
AlbVFWwWgfGCneu01GMGJquWT5DQEyUB1bOL9JtLoToax8d08Z3mSA9uNX7qq4y25mta93n88W2w
705ld/6ei/He0uuncWN3l/vSJGmTzZgV17FzMsJxi0lE7JZbMB56O+JlYGWR6qAoGWuTEdmzCFZN
jdNoJgzRGgy+8kXCm4HiQwDPhqLPvJDyqTVuvWPkMR0vHFG5sf/a7js7ZgNhPXuh3/idGHUD4+jo
8gJye67eHV693sGACyy7x1b9zWxBqe6kniCKXImy1+RMA5IIOHkCEpBXeBT9iWp257iSJk9KJf3M
JgwAvS1ZNxg2HeshglnNYTqrZO/mPdm9Kme3q5XFV0NEBOTZkd2pFNtGABnM26Ak6G0qMgVyv73T
XUCsAmt0jFRdjMwMannpq8MyToxUT3tyJ5EvMOsVo15nAQhSn5rKKpt2/8pj4qtiPD3WP5lvO7GN
2raL/lgq0/dlhkQHQtRIaJVYV5VDShK7BOVWognb+xD4QTjeeUvBbJOEJbFiHtjzQwneGl7If3+G
MFhL7q/U926jl+xaFs+vO9RyrxJUjH3O6haufrt6oDMkH7eW5KxLKsLTQFadrcDgv5mzsyZki9jQ
/M01UcXUEPBd+X2HGH3hR5n8Riej4ygpZE8rc3Pm+dWnAruqNoLSA53wWJrU01au2jlb1uTyYq34
hLLCoA1b80lBPJ9O4J/CCdL5hWA13FkMD4NR6YQU677SKPIXELPq9TMoyNpWKPVMh7CXBA1oY/Au
KHwntRzc8wg4xIL0LhYZJCiEvUjSnMo9uKqVcqPkGd01gTXnF5UkroGvWSSkU6QvYjFAiAucGAk3
XuAJ2pHIRB7wfu0Zu01EYKTkWkaKI3vYPlNFqPBTZ7D9upvotB5f8fRFc9YRtr+MG1mMkt8oh8bi
wrOFL6JDibvWmBRNgQ6aofAdkH+9Ex5aWMKQy3hrjio9ikP0FBKtdOP/Wj3ncjSbgWWNdzChAvje
N55nyxYldJutT95k+qJKB0CvP/njsGC4fjr03k3TDI+ZJcOp2datUWGFBymY222NwhvaRV2NQGwE
4OVxLdpRLiJ7K0TYaLKIRBB2PR3pymfG4YlpDLlgSfVOOod/7BMlDHSOmneem1csr2ObiioQ8Ecw
C59oGgGFjl8L6LknMo3B0V6+6VrrYasWNKPJJTCa0OJ7B0otLeyoHt35DjmgaoBx9kvNoDu80nVw
0uuPGVjEssJJAR84WoDSRYe13bJAD20FKp4XFgwMmNM8xSA0Ev9jRv9gii5rESfTVd9fIHCvGLlx
kdStaNb0o4wk3gi3Rvy0UCHhiKop20gJqFhcDk3NdjY94vNfQ9TKSZ6AfaKph+9v3oWnDCMBlzw7
YedzIqERBXOGzg/4nxE0EFLDhaQaAOb+TKlP5aSf5IgqaB1yyp3WEYN3SDwZqCnDUTJtVoT4HvEF
1HDfAaFOZ3XlrjtPZarfqe0ZvjUXTgOysk5OGb7FvdGZqIJsIkvWrgchCro/nuCESFUmj2XvCc/Y
x9uMJ0DOEF6FeMa/3NG7EkemO2RUt6dCsl8n6p7j8POKKGF7TMgn0+ekKtAdvZtNVzwGkb20QExr
j2FKAX32wmV9MCA+eMtOMn/U8qFo2C8Mv2O8dFgxADA6XJwkY2FRdIr22reqtfhRwfJv6IxxnLOH
O3ITPeNZsqy7WJym/seXgH7I/lLabwQOBLi6cg7gM6NLysx1VX38Zrxw7ZKKlSZPEULuxyH6me8k
o9lteFM9FBoIgVrDYVV7FrxwOE0A/4K0Su4CgC+IdDiYW4gneakTdZuIEnz5j4SKFrcylhyB9stC
Tmhqs608vS4rcnbwu7+cWTw76e7ixpChxgI32EdT4xP2IAMrWkYrBGzsd+Q0puSJz8i1pmRJ7sIL
2hF0u+/+mmqtf9jUt9HcGR67Jl9j+RFtwxyxCP5ck/PoG3W25eNZRvAGj0eiOnGU+RsdBDU8c/SY
gmbbHPAVeXE1Hbq0Jw0ZGWH/aJeOsJM3rK7XgxTg4cYioN5ps5CTK62X2Q+e++DJEgWgKNOFDnPr
G7r2i5kRLmEDsNfM5UhmNBK65Nu7D3LastFYfqxvA+DtXItoPJUkqoxnzbzW3PmhC55dBt5bcGsx
rqqFYYrqUEIbDD0LczXLhUws8C374Fow6um6hjdB/lAekATR8OPEnYFVYl44I2rnDrTWoDdjdM/R
zV6MwOTJbQ0Jw/1fCpWt4vmlk0qlW4BZqezGaFIjcTZNl/IoFjKRy1aQ7MtDolEEmXC2Ti5iNaKd
Q7k9aKWZ61o/v2Mo1JH51OmtPFsdIoN9ikcSaeP8NL8w62F+b6GwlUa0DSPKrsajvLK1hSLjSm11
6wyQV2FZM8y3PMdUIKjEAeKx/kaaVoqI09R30Ovg+4KvoSzMnSOzicU69ZeTT9h7AoSkJ1r+UrD9
2rk36LFrDQtLnO7MbGZskzxk9ysbHEZBbbXd7O5GDBjiEtD1k/YEQ5LsvRfH4bHydUx8/YDA784j
YPMzw4vBZFfh03BvZ7kfse+oY6VkKZcP9/9kN4cjx6et5jgKLHrf8ZGMcqIKYqD53bcHqTmIIvtC
6FIkZttWoRIXa2WfCmFnHhsJJmm5QLLM8t7YoJ6DvG5seS8AYpDu+Btactu6Ycbm2kWt3aXWEM7V
bGo48fnz1LG0YWzu2FcWZBNapModWaO9X6V3HM7Ws1h5xSHjomayJ/nJT87I6iIX2JYQDMzsKOOn
kRYi7QG27AgjUMrGlLaQSD+hIhkG9IjPZzJZSFMrYiWPR524vEq5IQoIZVix6i6YoKD50V8lRwK2
AygZ+XSSIPLBLQoMmVnSzfLhiILgtajiwTE5x7iGt9W1Ku2E0eATnVQn0lJ4gZnd/mO34eY1H72f
erw9BT2Wo3EI0cX1yHSFwe9JADtfBxd9ZRDIYUtNL9WpevikEI+jjMKuNSIzJut4dD/Zw6qE0Kgl
yRiIZcnqNqsTaIwogs6aQ7ZFCLZ1xZQInsr6W63ngyxogfdwGffyEWhhORW9Z+cOwoGktFH+gKJf
YQ0eMxMsEKSEK89B0sV0eJUGmEpeyibenKdyGUWjvf2UrW+UZ6p/m0fXIFqhGleTYrtiK9wno2zh
nIm44/lOCtQXTAGBhqXXf2BjWpfdigRQ8fZDakC9bxJ68acEfBE3OiOR6EtxDvupdsSJ8npUfbX+
T+HKc1PzjTXAPW48kWdIgNg6q6DRqtMK/ggZEBiKldInnx9l2w4kYFiN/iMG+N6cYpohc0QsK1ZG
omk7qbDQvIvPo/C16Xv3V9Ckq7HxduYEHTkXd6jhSJf6hS5rWtrNv11KRdgXk5sj66LGWnC3GARv
F1K7in5l24mnk8ZTsk0A4cvs+E92bYGaPgiLWSQWypxzgY68mKbF8q5gqJb3o1tnyZ21FlPmGn/d
7Uh3GT7YbPs1OM0kzljD3ee96Msfk31V0r38PoHKQ5vrwzpMTZqaw+LmfKW8h2654HztIgBOAKKH
CX+HgARCAwO3ewH36LUDb9p4FyqxxRvG+t/mDiCu1Jp1EDzTS/Xo+FXPMIbmu6kww1Dse9vUBHNa
YeDQqdnrZkENZqtOGJFCV7iPYf4PlNL/2S7zbVUSUusLc34bthsVsVopTXwXzA9ogim9H5E5eg3p
nBD4DXKHrT0XyfXyMLTcOUnHMki5lftIKzvmcBUTI1MzY6R3JkH21dFgLK7OinnF9uvhyf0c7g3I
z+jqhzVCbZ5U07Q5KrAeQODwklm7GPpYmuEirwRj/Mgi0Lgpjln34YT1YvokXyXzM8PKyFkJqq1w
kZvEbjERll/NMo/pocOu74Ze9KXNwYyJrbAV54vqlqDRHCLQg+30vYgDSGkANUD+znegKvxBzfT0
zAN0J460PXIb7PW9s0XPnDKXE9oQ6kWnMb2Jw1+9ZiT0sy+IQ3KKD23POLO6vV2HZdgs5VSWJZv4
JnOxsFrZyyjQy4pRKZvN+0LLyZa+jX6qUxwvVVBHqoHgUtIi/J2nRxw5UlXGcAYkv0AvDZQr04Fv
ezChRhajDTu0B3JYeinZ82Yx/xVXbIhO1E/YcTiMBGvAUd8BkmUXDyb73tniCKnP49is67miRyu1
TeCb2CltGWMx1vBhRRH5/8bVn7FPb4XOx1lKlhJXlgPzWTmpajQJfQUsJ0jj420qdIZDvDJcbI+b
x9hS4l9qsIxCc4vKm/VqhXpMAsNWjLpjnUeSFhkPgapYw0x86swD8R26z9y4zDiL4lGxW61Fxndh
LP2O2TM0kaylSD6zafa0ba1MoiZ7RAIikmhnnmm1euIRto3/vKggJxFQk34GTpbtt+Tn+tDBNpYg
4NE5GTqcGyFZrJSPFfzh/Qkw/7HnjsauyhU7kiAcdI9j4WLw2yfE5Yt1fX+AIMIc43qHo2X4n+Ml
WvwUJJlE6q76L9TipaxkFAZ1nRnQIPOfN0k7DGQjwSl8cHkP/nFN+0W++KcmzN2wpQ3HTr1+izXP
S2rutQvxnkg6H7rRgNeifuV9nNc5HowfZXn1yq4lnlDWzwzOnjTYAqGlmWxrKo76aovQGSSu2y2D
SmPFCAJ30KOSAU/bSc+aqNdjwI7G4LnhMS5Tt3q+TBfGK8CK4/PUpD+TgttFehBa/Mk8rlHQG5qa
ptvC9HB1xJM1AnyRMkx7ZXFSwsM6RTVDqbxxbKhQJC6Q3UzRE+U+22Zd5RoZMSxlTiBOnJnA9y/u
Zz7NEzy/gRgQOlq2oCjS4NJl81H7lrS9UBLV60k2RP2n35b3M2dWWI/MU8fEg7QPy1K6j4p2tA1e
PZbjz6kUIhe1dl/4N5mYKMqzY7PkZ+G5QLJfEYqI4nEellsT2it8N2dv5zNnjE5TtFJQEnj9QhfD
cFJ7SeR53sdpgS2WofJ3NmPF4S4/bvfIvbD7FvBfY2V1dhToY2szCQdrbbmwf4rnCPTyARGFBgeS
yj7uTvm44bNMlPorPkC/hABQMnl0dUI7WvIIu5Nlp8NjuA0hfi7q20G05hRoaP/5YLaE7zqMzK0R
XP8z6k60CZ+jA2vOsv2qEYNpGjaCIwD2IznJj2iYmSgSgP1bgs+BtUIkEYrqwbPGyuD+VE90HAdt
N49BaNocUDtJYsobqu82P9UX3KlxUblQ3+dbAm+3anKUHc4KN4tVkDOueMT9ls4vN1Tv6waHSE0i
CRGZ3miNsrjeoiF70ekEyJ+kus4BSaj1m95CdILPZBqU9t+f1YdCxfut6WSae9Y0Z9LIoAf9rPAO
AWabJwxpQ7m3I9vO8fW5tBO+jgy5FK24w2FDAp6/Ygs6TkstRlAX70m+RJgnWHwqgFICTCZYXn20
mxbdIBVmmKtKeAGURyNq2be+Ve5ciq3316wZb2grkVoN6ixPvRWEUY7qw4V8zKJqujWR39jcUHd/
ZiCh8e9B/mz6gXNwUdFIqpsQ4RShraK1RZyN3ntZfHTNkiK8r/0ooKSUgIZOTAg0+c2HbzdSTCap
+gvmCH1ExTQNs8BcnpVST/V3BhvGAQTbdS3x9xOXahnoJaMyFa4hZcBzzZSj46krrYmKfbJwg/0Y
5lFvxCvd86BQTfQzqcMgPx/i5X/Ow64C5bkts8QOYg2sMxeHeQZZyoXpT3Y5j+taz0kabYNt5f0A
ZzVi2DkcO2GmPCreePHzmTvm/06UYoS2/qoQLgPpjYKBQffWOz3Ub04D/rGKH+BuOF/JKO20M02H
aNtaesLLuMd2xMPMfFxzp8LmYEEzB4UttZTLxsScbi1PtvM2EiZ2LtgiDRDYEvGa+j/ISkAJzEYs
7WXBwE0/eu/D0YnVpQ6+ofSmRbodEaZIRWSA8pXLierXpPIx1qwYYJSWJl0FOlGQFtCTAYZNdFOa
ZwC2MW7SLiT3GEN8OcKUa2n0rV30ibucvGz4pLHIN6mLdTD8g7/+0FC4tCMnkKMa13/8aCVhQFXA
gtSBaebAHFbIAbzNL3G88QnOPejFFRQysCMo45u5v/+A1o4G6IADBTSmvbUWAr0CY2LsrzrGt5ju
vcVyN/O6S7vtksRnHA1Tu6ZOo3qslNbseS4hnXp358E+6qaVVL0muD5owK67tDmvXD/SykjkmovR
6G8VaIU7bj0U/p23E4j/gGG+2w5EhBAsj3sBaA+yBgKrHoMI9qVeq9WaG0UIV5wnAiC8LZ/TsH5u
EC1opG7pwiy4vWiBl8Wwrx79xq9grd6PE8S+03vSQtFh6+aacMXDDQpZHWclRivviRvPyH1J1YD6
ULzmouJh2Cmah0mvlTaAU7zspImBU7o4HIZA21fYyo1orLBgvXs2E5iARctSw10rhg1KyqKGThI8
fDUsJwyj6phY1QzhV4s1EPR/R4CsM0DYqCQkNaQCa1ud2O2sLjgULo3GmmPrQ9Vlj4gW3JIbaKtB
UOpMpshAx/pxNp9URzGlBdTCiMf8BonodxrnxwazbNm+19kvBopiiE8RacGVaKSP9S1p7qlr91lo
Cl09VmcVarvg9y1yM51JhLj3ivmXCWoSOM18UUG9ogldlzGS3FsTppiQdh0jZqYh1W8TRcA9uxro
peqS3Megf1qFzm5gg91+hskRp/hSA2UAKfCuGGkVK38ZWTy0/GhE0ghLusq0hd1wnKj9bxcGdlf1
BjgRObNJsXlnnj01ERZodoWy7soxN35OVkBRNO6xIhQKqoGC91X8Llr5kBxPe1nItDbdHPHX9jR3
2k8KD8JiD0QeMvfUIlk0lFzOPnsIACgoKEJCpPgxapMbnwvrOX70X4c2C/gOI42ZNs8Ej8dgVCOy
0olNLRp60Wh/e+8cSDQylBbRMAAxzFZEfYRYyecgp4CA/9IutBlfp+uwGIQXulZ+390pxP7Tuhbk
PPzx07MjahR5oozpMHs582p2dMS95UAisALo9ik8Il3iCU44UY1yoQHVVGwxk5SxA06du4s79wXn
TreGSrH+47nrG3wJxVMrnGjwm9p2BgoDM1smAxkYrB6NNu8vdXV7Hn47bCchx/XoM85+h9nauXyW
iDm3qyK20nH7r61y9av1KrHRwAV1PIpyKQxMk229KcSSkv4nd/9S2E4IS9uSJUuKyEzSVqT6rBx9
hEg3ybLUJxjCzk6HPNheLihOPmGNAk2rIkcRlS+2MO2YriUVFNOd7EiZwpFSFZeT0pjsTTgHAmUl
XxRGfQpxpL1qe3Lm95nFm+uWwwsuD4KWlHjtnSVxw/C1lnf9cvaca6lqGme2Gv2Ol85UVv476YTf
azC9oB3On7tTUP5wVCyPyhFZ5Rmm3FD38u19uw2eG9km8f7M0uzxKwPIK3LnXoE50FlSDuCibW3g
Tc95wYe25GPZ7VGjMiWEoS6W7SeMCxHyr6pL+A+0SLpeyweflGDppNhP1qKhBxoCvg4qEj0EPXzP
uWHISwDBXiWGfs95t0NtQch89kS5S+NbZTvuGMGHrj7AMqwvvBeT9/1dJMTvcwjs72W7nuSH7qVM
K/3UjlXHALowl5D97kNfDJuElFM=
`protect end_protected
