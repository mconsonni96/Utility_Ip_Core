`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dF7T9FS7E1CalkRA7L2RyjA9JxraYk7pI/Khdknzw8pwX64E0XdD89N3uhh1+sRWcPOxai103mZd
1Tu/QHvRP975JTq1wVaeOFwy0mxtPhmcC0vyCMJV4oW838oL29heq9bF4YvOrN5QWUsyViraDfoK
LuNMycEv1Gb10/nFpx3KUegEZV7Ew4BlhM6+K12m2rndCaxFfXr1LbsCs5KqvqI5og7lmAQZDkHL
DmqOawPXBhBD3N+T4T0/AETfeY8xLE/WJkPTQA8w/sRP5QeRXwMSOnaDcYd4Xe3nYh4bjM0CqUJN
/bUc/lzStNx6mLytcsYPO9SE9A4+043jwGDiyw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="WBaExLfB/8igPd9nzCCNPltsadRp2L1/ZO3Y/hVCrEY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25088)
`protect data_block
8gyWBkkRzmA2ur0vihw1NZR5uP4p5K6ptpkli+wqP4TW5896vVEnhmqAxL7bQdctsFd3zwfwmd66
hgbG6V2AvRGIPBsodiy0APJX6BH3PH5d7wkq1/YDxlSbtj4ZCSqOVgg2kY24za9sNfm0UNV3faXh
nxioMv68qdRkN+AGPOqcgwC0p/1IqO7kPtzI4Ab7oSW3G0vmzyhSZaj8htKwoucJTtvtCXJlk4eK
iF0J3o6TZYJw0aE8s4G1dyRT2YN7BHQBv9UMnmCeSDVnajj2MWL8nmgS7IRAzpGlfnniTgqTm46q
x+NqDgaG12ZZ1wnIKrO+PehSHW5IA5kWbEifPuf5/Bio96bZEapJ/AAv9KbW7ATRAKy/Fizo0K4w
5kQzVkkk0MOFem+77h1bZj6+HeAdIYhvMbuM4si1b+GEXic/IkeApyyH/q1zrJrSrySeRldN1fck
o8mQyIGZxeQO3rZS6QSnjbhZrfRNwchA0z8didZYh+QREh9StjlEFP2b1OIk+mUqbKAM+6oHLG6K
LqXEZmh07L0Qs1SRdRjQLKADuYqQ7uyMG3W0UF+h8Cp1rBfzaOE7H97e71N5xM4IMPJvWnFIp9aZ
j/P5cwH6EyzBG3xZLpy9T6siJee7A6dguEJ9G8PI10TlLG2BkWOtHlWwcb/30nbPi2abC+nNnsVO
xpJMod+hXK2R9dmH3f8dMbKplCCmzHkEoFNqcyQUE6SFUKs8eQApwfV881/XyCY5Z3NazRuMjxX2
qVSu2qNRHMKFTMNYJhLdZFKQLHydjH+Qwq32dJ8GC07loBgpnm1MfZ9dVUao2O9hj9cPWB2QSWCB
Ixp6VOXSU21zWxMoSlLTdZT9g/p4iD089SeDlC3jWJTir3B7MqBWQXhoWHsRnTpUQnB96XFMdaOb
JHrRXmnnOdU9PuyraaX1JirdMvAM3wzwp9w3nK0dlZa8xoXxs2hwFGu8EAqLdzrYpBm9pctCfSZO
0DbqD7dosBnxpICmVvfxqS8XyMYxcX4NEjx/qNH2R1SZPqozTVE6Kgbzd6D2wWZklM8XkjhfJqwE
v1wYjfWiA7WjfuDkmpc6uBWnxoJ4BWwioGUtXjKeGVK0haU2uZAgnmZ24YmS0s8WkOomVIaRGBz5
bBlkQwk4S4tdMnOUMwKJ9AuTBjykO7cpGXMq6/8qmegt6IMpMMkY29JTBAyN3jTCBpkhlfc6eWEM
Ul4j/7rflsGuN4m1zNksDUDnyRUY46MgoEmhrBiRrSpp1pCileE05P4AgkPTGy+4jJjhvmELGbUV
YFdMK14F1W41SETkYcMR0qU998w7VqJ3Z07u1HRzRg9ENMmC6BBmXI8iTRwea5GNFZl7ROZdUXMu
F+CV29SQtEys1yZZi+f2IhhGsIvLTS1DQIu/6lT1MnzLyOjvPKvTcKCnZceXSrppkUbENFl6d83u
qtuzST1ZleQKXfWxjJwHxd/GzhrBZm0bmYY7OKOrxxushZB5JIo5AsGyWwlAhLW/jZyKrUZUMnML
9uFlxo7WVF3HBbwmketDmM3DeNhSN6Bej8QeN7IIjeR+xKcZY9UkaEcY88FrqA1a+7Y4xkAwRy7N
OABYqmIRY/Yt/G41ViMUNuhSArWdBU72IDVOLlyrs7FZN3QGCajnIhX4HkJim1f8/VTxLtdDdNOZ
2C0348TB7hJ7PuFMhKaM4s8656ASwADD0aZ3sT4etuqPah1qUQ1zKK5WWHGzFOhfA3r7A7ZyHVr0
39loKNe+9Br8bYqfh4DDvqrCBMphu9SkLRez2g9hGWvjiyspQ6pIHfnfGK/EkJLfP7p3ziayw+N7
h26zBwRhCfg7Qdi/kYXfRvzRf6I3k4RzfHYp8waLakL8xjjA8PAlp59EsDvnWPX0iL6aaEBLT55l
SKU1kV562pqArvfdqtZrfqiXOlLcjHZCK7kkQcbN+zfs1ICph6aOS0C4eyK7Gtna/DinlyyjU+Ll
bQC0Ja5CqMIcSmpGeavQpF9LifqQ77GA/ByAGnZc2IRpPNs0J8SIfZj8R5gW7G0b/JTUvRC17Mnt
J1gol7oDcjJNOFENhxcMEyMH8RoY61CaFIx4KjOXrFG5cvYfF0jfuRFQu02yTUEChD7u/g1t+dnn
0rKMDOt9QpyVGZth7tC2KNl7A8U6/tItZBpdSDqX+4WzfGSElMJ/jjetH36PPrxEsa5B88VdCldF
nFUjlDuc/oTPmXwqo9Ryl00jQnsIkAoBpzPyGEL5Arl5qIJ3qC09FbS/NyjFltJvlmrJ2NlRsu5p
dm/MctZHcllod3+MHx30ZQ+6wUNVx9s5uY0KWjpf7GvMWvIRHf5lfyRShpQsHqeDo3hwVa8ZGFjR
Rdwc0yhEheplV+cbdR9/zct2PqrbBnBcjybGzWtjzv+G+4nAE9BqG+p9fHbaOdZo3pG61THPSNY0
MmAQ3xdPsvVXjYeYCVuMNIBeWqqQyWHdqnatrdrBOy5Ut2wbSLZmJgUZ+TEFud/Oc29N+LM+a1gV
vC41Pf2P2eyfwbo46Jpxi4W5w5XTyvtbZFjarne7/OHQBIISssVAmN9wKGQ1rtHUiAAJtNr3/H8i
O2LmxLpurBfAdALB00r1qxnCyvkZifeOQtL+qUNC6YS+wImcExZErDovos6yFG+cj/sbewsbqImj
9H2CvPwa0Dr2bu6BcjWhmOsmPPT/R75+4zrX7H2LGqXiYNxlyi0IonI5yGuTBPKhMuLrDhal192W
HygGFrWYjYNHUSX0EN4/KtAtHMQW93eGsFj3mYu3JN7PpyA7LG161SruT3pjd0gh7wHVPW6v0D9c
Fw0HnGI8kCTcJ9DTIUPioiWL2HvTuA2bMaupVst+bMO08o833Bxr6z7zvxtpzzkk9bLeGRvVZ/Nz
fZyGG2t1O63Iwl9Z713PyasPK6VYK2i8jXokLjxTBkHWC1txJevrAnubnB0V6ufLlrUFV/JdyYkB
9+Nw1EWWEuaLwu4qdZUGULoK2UD0c8nf3fuNoY7vhYSGFkk0C7vm3cWh5Jz0hF/H2omnWH/3e3k4
JglP6KtpCuqjELZtgVGge79zkk0hRfTxIT7P6/hjeG++Pnmmx38gkLyfgWzObTEm7E4jW8sG6/4h
supjL158g5LrGo2H4IfMBCX4nmHAEuq2W+SzF1xFCJaL4EqmV34QVlo1Zc6AKuiLqVfAHU+6fmX9
0XE0mp68ZeO0CALklBV+8WXhwqATIgxDSsN8eV/Q3lrFdBGtG9vONpmt/bhdKYsrkggYNAKcZrE9
k0NYmWskcCXhCePcB6E7QaYrEvnxtt+lxOVlVn1QZtF21CaFcGrPgQHnfA1moY8oLVFV3EJ/M3Qw
TeOmV8xTTFtBtRus0I6h6s1lip5LlfMaU7RFbBMmF5YzAIWXmtrD4pjJpZicVM1cxBpqgyTRCYCZ
UJFiidrCJGnxXjbXKq9Fuo/fetZmCHw0quUxt1dQ2ydkmjcq2H6gPNgVMVjzRn+AFpCYs0//5VVl
UWRRvkQz6brEBec/z7F88QYjTuworu4pY5sUHLa2WCRz2FHN+0H57kxRHl3cE/ZOOXrqn1K8CKk+
p6opBKm9NlcrXhvHNNj//rUKMQb4v6rEXVKPbTCYIQqFYLzWqOyaB6PKxjd7888bLiI+g7oGZ7FH
dYBdrZIKB8b8bH9MIBk+6FYUM/qLBCR/rp5IbJdN1N2Q3fEaM7SgdSXNPG66X3jnAv+tMegB4i7i
nptowiu8v9fU/Gy+3U1I1XoY7gD5yrRi0jfkVyR8WZnAyGGe1Lmk9ugcVCnbch5H7z8puUW6So10
+6cTyVnR8ug9JOVSuGhEDuiHyKaYYP0OZ28GcacBHlkBHoXGTuTfxhaIZ/7nz1OjDJRSPkA+CH6S
TC/SQWT0aqlBdZUT+I+cd5xmyug6Mq9dFT75SVMbezRhLMvhrdWgo4LEYZIR0Yt8k30L5BT1XzaH
SCY6bel4aTH1ZcGUMosp81vtxmlUTzEKAG8MsfBHRYiT+OxuLl9zOzbHGUr3U7RLVJx6etv1+WEK
VlGJVCzEB6IrRrnV7bIBETwSO34ysI2VR0OGjFKP+om5LVVvoUM1nTAKKDadPBBRVEIPpaRHgHpi
jcSainN7q/rH67hTFwRsVVGF5Ab6+oohygO85dOLsT39J14LHthiR8gweTxp0Ru69aIRFymKWALG
S4mOIHgBQ0CEsRYcFXjOCm/DyRJlkWPa6FV0Ko94jtJWxYYt8JIVUBGCcykh9e7v6W0EUHBdp5Wv
KThsFswD1nmWt9H2FtjXlZzFyhoFPbdvNOMGwiIAyHuhRD+fOrPW3mkwKjg5gOkW2T2gmKInGTEw
2qPp1XSVvh52qBVbkGEr18xv6JeGhnhZLTvba4gbhTwTXS6Fun2l9fo4Jqx9gEwMaYh3QqEI9+4L
xqZgeVGe2GQsF1P1u3PWECah7PPoGsrvYhvMfrj/ODjEN0BEQ6pbWqsrhTiSXiQLXOiQIEsLDJCM
4+td5GusQFVZGq0kAF3kFHxYyERzPvuL6OzMl+c1uhFKVG1AXdmhFtjl8xOaUf8CIVgCZ3tEhyXt
763ZkAQW2Fw6EB0IkJ/a47uSkIjtTBzbarhRG+dwu8nraxmYWDnJuK8ZxNfHcUqmiXKfnVRudbAO
AosHlf9AxjKxw5I6RdvTM+jVGGijU4N38VQKuyRq08FMB9N52N3oJJNrp/OakcIP4GHvPciC4MZv
768+8gjlTRuvuJm+S6j8n9iSI6e7aoq4PdiQvYRZoX6uuOKdr0j5HTk9GCAwOsV2N6n3R5s5UB1B
noK0uM8j98KMhq2slH89nxgaR8bxWjBz30TQmEde5skguDrYdm/UUnPuNptWGbgegR7LJ8TKz+/v
AXgL7xqm72psP2V6grpA/kuc8gjdTYU43LBXEXoizUCY/JJluyPjrWOHSZFzOI8GnFQgxWwff0qd
9B+I76W0bLS9fQyZYw8Mr0uwBIz4fnWJLYORKtaFjW87kdz5Q7AfYK3o6OfNkJVI2nc05hNvOv83
JkhhrZC9hDtUEs3oJiHrZcbs+nga6yfP3MFLsVSiBS/XcvJobv+flV/ZSNzVEVr62PEb2U+N+K8R
HmHqcPig4ED+ZgHuZboNIqDq/9f+Nc8T72PI7tBbjBPF0Np4HzbNRa0Bpp5S9ip86VgkTaxuKnc7
+ZNkjO5ptHpaAthtejbdn2IvYjNYYTlWr7RVrccQY4EYODo9T8zT/VTpr9jSJAdRKP+84/7Xi9j0
kOLCa+3lM5j0/aJqhaKUoO+tmeD6BGberX4Wyep7t7eN4ZW6+v8KyjaLhS9Wv6AqLSh2RdWrPkVj
NVi3t7RiIxKEwzyJ7qV7/gL7wA2+8//z0GgS1lFcrMgoKfIYWyjtV561gDHQDUxxC0EWpTp+Bnfe
5p+URBMFdxmdit/0B7To0IxP801PzGjrz+N2nlktfKhN55W+qK6E54O0eO0aVRhQJNztluV7i8Rf
IV8bUs9oVsuZygQtJy8gELQHoIkmATVZQeTcRlI8RjbUXL6xPqJoN9yxN2HEsCg+HYZw5jgGyg6D
dfwrKgMxQ2tuudUKDm0nV60bPlUDJ4Vw/ZRlA6xiIZOua5gNJpMPxXuaw4YOTLF1RdSP89hLB59O
pcSvnl2T0V4D1uLSwEPuYSmFGIUoiAw+g8OgfNJBO6KgtjCIYRWB4smN+1XrpXByvx81sKDlDGW2
Wao5AjxU6GA4hOhw8HoSebuf8GeKh8UryNt/pL2KVbe3lo9jGIHg+/CsFfdM8xi6xluB7Hue1fjC
dXI/tUSlqvjbz1oQmaZ8DlVHDzbYaDphpb3Twgt6z7Ns5zZ45EqbMOvis+oUIuH3RM4BQwbePXFj
RE/aqZ5vFVBQKm0nkqOqx6ZDfccJnTuuVKX3DLxrmQ52BSA5PwNZbS8kMgl0wYfk3b7mLBPkg3/7
B1tWDnmtV9SqCvjB7uq9+PgWC3XcRgfe2del1golRg3cR/P47RRl/2EOHh0OehPucBsuSaNxE6vC
DTtuVU7GSkUivHMBvgdJC8twwGI62+vbYy6TZ2E558W/BX3KGlcrXCB1kMl+jUdOTLeHHt6BeLxF
i2R/qrz+hFuS+OFHFP88OetJ5gAnW/2T3ok89dRNK7wpYYDLLyHbmA7IW0LAKuER/78UIK92Nyzh
EQLG7W7g+JmU8kF0bj+3B0ijGKcaMpNBKkaOnmbQraAM842f8PFsDsUwKe5I/mZFu4IWBnupFosS
RIlv7F3lhD/ODWVlrWJG+YqqAoJnTlKai6zaEREKkwLDxDfJA0UCunv/fJZ2H5+PQCZ5+V0DcpRe
LLGBGbKB/AF0KKcljrgty+lm2VDNGtiosCvjFfjxgkNIRs1dITEskZ0fBW3ElTiv+FaDBm3uO6Y2
0qXAHXmPSoh5CSYfx5frZNWnwHWsywMyjtjq+mZRaxL32C7dx8MUOed3jglflMddVGQFLNeiCVQn
VWXasnn9LACu6chwmMHJC2NhbHE9WWu9jT7dlYtsZsx2v2JTcy+QRcP3owkmdqRRA7m4F3M4zFBs
Z/8+OBIhFmvb1+a/dD50HHVcCmMoiFMup+Qn81rXm+W4zfrdRt7CFmAq9VqJDDP6jEOLp1Kwh1Ic
+gwd6PN4ytPGAkSFu2CdD/a8co0Z6daPmAz2K4fIX3ZAcYMfqEd8Kb4h+KxKBm8Wzj4EXYggcvsn
55qYiSyvihHYjpBBUMmqUVMngIcy3nJWM46elfFkWbfjjWQ0bS5LNCM+5QAnFKlkBaWP3Vl4iRTE
V7lalLlrisudcOQnj+Mq3RtBEvVlDNnr5mqkCvL1hA0zCdu0NSz7JpM6Wr7u9qfwT3zMeLSvkuFj
8EDmm+D84neCI/t/O1xy+yKVRGav1BipLb9cVdJhL5tq2nDUiSqm09z793vnLeumFkfjT5X2WQK5
NLjb423bhZF9pHUbhC9ekbtS6yYehadEoPjHxXV+HHk/WWyBomqmU/pnahDHcZFJfIxsazBd7BHc
szzis1aAVnurhdCBp23CP0hcm77WvWO6/wzlBy5jGZIgyJIa2dcv9eJcSy27eU/lMimtiapm0yNC
/bVNSOoqLR7LX0+2l9kpmfYMBTvHgX529bt1+udNjKM3UlyitABBCZnLjOuJJrRTXZfdDMyTMIFT
2u8Xaui/twJKC5pF/4G09Y5OJxhgt4VaOKzD0IclgZxrkOZT6wE0ttWrhy308ecCQ0b8Uvhvqycy
oadVPzbqrjs7B83N6/yIYzRLWEvy5UUkE0OBWRBSztUh9FS2AcpCJ9FxGl6YDwI5VlTXka9g2aIo
TeKkhVAAKaG7ITp0VxdCoYFe2yL816+yvCc8t9tpuwuDIyMwvql04mcrdlnn1996Is97x1ewFhxF
j3s330LwrRteLeV7L4ccn9xO5AWsuajO5dUjiCQUf610JEYYd9esDc5wd3PhL8CD0Oi7N7VbtUHo
cEudpF8EF1RNDFlCen7OyWBUlZ/kbObZMX8Ek27mSwdtxjh8xTU12SBvzC4l7FvZ8fWs70USRnwD
5+qqypKOp5AFm5+SEekk+Wnu2BijVyfsbGk5NZ/thoasXR/NUxjtGkA0PVUfmpuAlDept9yZX78c
va5uDDYj+MEATlFZeQCXQy26ZAuNkXAlAiXLpbNvNF2Yob41r3gCp0CsRjarA8QTBK4vOL2j91Cx
beuDUnLq6rGyWSWmZ657SHlttvJlGO803UfoL4IZ5zSk4f4A5U9nY7ilCrkH7JJl4QeIJ+SQoivz
S+xob5fjSCoZuaz/MqjPKedXXYJBA8yMNOMpGu+EkBrnsQEsjpxDDyIG+s7opDh0lzBBNX5Kvg/D
/fbnCnV46cBdxTS21HAtfStF7aZC8T2XMx0VbrPq20MPGDuvBv/mPwzBIWtueyGvSPgIvQP76nVZ
pp//oOaCWKXIsCurrnlhsZLAGrtvuaFLFNKg+Fz0aOE3mOuTmrftEICCE0Ipg8yeAhD4ymRlLu42
A6L8TK79sciXuhT0PWrcufK9YFsuam7CHz4XgnNJ3BYfBz8VXHscDNWwQrlgnuqgFlxLTAamINsZ
mjjEpcR5BmVB+1cYIKupvu/Ag2BWZAB6izE8T4pWdsfwCuyMo2iVcApztHgnm6EkGQO4c+rmhGhI
rSFjDAboMzNYeuEV57CFrkvdWxz2q3t/yU3WGmOvwBigZh0UZrGcSV7k8enLBObY8i6BYj43TaHr
PWNsXJv0zQ6Sk9c2OxAXhMumg8IcB8EGhpFUhD5iLbgvvbw4CbD+AOH9ZZkCH5hgsIqVeTbTs2uc
+eBYxbRps8O2sWr+GkNCO3LUqpurUqhtzheYdNK3yXDFIyIEm3VtfCHzxYnTuUiZUTFULEUjSKS1
KszrZuvT+ISDF/i+wI6BDmOONLMHSMB4tpcC2S7ue+NW/c3F1XDCf6ORD4q4QFohGU1o3yhVge5L
qgtZcJhei9AKiNG/RrG0H8F6ZeYc1O00X1F0CGVBWyDiXWiFYoZagEZ9QZj8TTQSIcXzUYJKY6x2
UpwWtvPUVqmxJf0IS1vkgR7YLWyl9tjL1eXuYTCAV0xVJVMOj5cK1Pqe5fPF3XjrwHycRntyVRlL
RKXQ9UqWGeQvGZ4G01bdVza4fFSOdYk62gvAHZ4hsz5PLFQd1lgOcVQ6Y0jorhmHyrAnLcSVQFzn
rqfkNx2+2WVZIMVmgW0OGeUrjHGcdp3jXhJBxcGMGzWYkfv5+YTfMv3xokvo0uVdEARisLs/zPdF
w7XdCB6IPZX9XnxHKiGAahubuAiMhlbdWPZ42Z0IAtdCjbjKn0jwOMl0VkPK4PcQpxmRLSTp0Hr4
WZz9c5Jve1SvWledKseSZtOHx3L78va5FjWNJKuCGOqvEP9GIcAucd7DuXX56cYKtP1+FYW/d83n
Edo4oCmz9/95mNoxdmLBEKwexI44jWkLT0wpJX8ATtA9tn5JXF5hlz3jASGezHZgB6XWpWDRdnNr
3a/rKSjhFS26nA/4NTANBqZS8wqqNqsYVXBlWxaOWsf25r3AL5oD/f3PTqoY3hUogfSUibBs8vjm
dwwPs/otFMz5ZIk3qR2Z7TkV8PDwUZflyd8JV/FgxXJgLincUUnnS7+Zk0CHIN3bFqfT0Xy1eqBQ
nA7S+1cfbMP/ijEumtRAJjTfjwb1UVkCZFdHNpSDpWHBJz8++y4cjaonTvZNyRxe0Cace0X3m9On
tjQZkp7yITVniHsZDNEb8TwvmaoSCCniDnMzjd4TemqACkASyK8EHUwKeE6TnEWUgl0himbNvTuS
4iSyVuvm8dpbvLiI8VVewhgcEcgELA4/i5pblHmOKhOgTF30UkvbgQS0aPapX6ZPFrZlssWCrM8U
Uo848F1LEnuSPyf8yUAQhy9CIiN60m9BMgQZMc5rDyz+YOmpd4+NrHjIKRTtUcNiLFOLJkJJqBVH
OnxCgPTWg8vSsVNOyS0q03Tkqp75UNNfPO3Cl2frG+Sg//5gtQqyzj9jkxoF8N9PPnC2nNSRdrNr
11oEAgQFawEO4+ju8l+gcXYJ/evDD+obYagoC8CDyRNaZidUKYLcqb5di3j6yu77Wz04n6vAIjp2
+9d0dWwZ3W8GUVwNdh/OSpFELAGPbuacg7Lz6Y8qiCJRNQKhDd7SlPX1Z1OLVu/uHILXS3GKO5WS
76wIxCIJu/sskwLPeZ1ZC01u15FOpA2SjZbdKszcU/rS3VZ+/4jULct5lC/Hfw97TvdiqZOZ4hKp
D6BJ3ud2wciFzFscRTLJp5u4ezhc8k9/RHsFCGbq/ov73Uh94tTAckyv/im100zu4xdipYJt8NLw
5/jjpcu1FO0QdvkC5NmBVPGOdWAjLLGNnpn+LdAXRt11L0oe2NwosRXLkGhWKwtBVlF0ZRdGFqfa
1e0yxBbRPygbUxBVD6tnPDxvh/d9Cr0a8PEVc3CsoXNnEBvYD7rUw5Nk07y0aKK8dCjj2T9RbdG6
qo/FOld+pVFTAyVs2DzApLRXUUa2n/QP9eUDY1VC3MaZkt6hvbE8zKw4446Cm33Eu3rQgSw618Ju
RHwlqaMudkbGiKYh6cqahbzB5up19b6LMJvc8HaPiriXA99Ptpoy01aIms0LZcpskfs2rzbc7bXb
fk2SAEu/BgS73oFBUYqPI+oDPOte0m+RcNmyhu9wjwUr0Ft+NddSlDiFuxdH5Z3/bG0umXWJ+Bgh
KyNeretY/kV8fMahB3haJYMJqJAIQrdKiOUJSqKT62QRfD0hs8dO1X1coIDEq8762w3OTIuhUTFk
JcfdYrxQJ0/dQKqU1941eYLgs4eTcv4bJqRuh1CJgYA/3uClC2yKZt+yWdVpbSIBqarcRfg9lMFn
S95yUxqVDe/VoIQobcouBGWnKuqhDiFN+V4NwS9xXPfVwjLUBmVkRpSsGfwkkjmppgaeYGrLz5Jx
52hxMJJ6nzGc+4hxLFW9HwCW5Er6xhfIWEJAnZQaN0a6WdX6BeteAJgMiib/UUiWOE9m8d7fPTNv
RN76la5mpfjP33R2/k7FxwzSEN/e6IIWkcyYXFxWizXfoqNWX999Bxyaru3u3CeMxJLQJWP9/S91
BwBqRadKPZVuF96l6Z5VPiNeKfGX7zt20RApmEP1M9Rm+rDrdIUBnuL02/GeZJYSqY2OWzOR1mXn
YRQYstRYChMnmstmJ4fMnP3sZU67nzf9mtn2Mdq/F1fXw7KcL7yQqfeqJskymst9Zrs8hhT4lnOy
LbN0aWTmtMEH0hGQROc3rI0E1GBy1nkXR+Qd7hX/ySk1+j/q3ud3GmvOPG1l8QzYyJDZkXEuGZo4
1i9r6EIRIU1MJSsRlNrEFw2SKSDLktBqbDB6WbwNzr9ZDyzwdXjyxGBg6ztcQeHI9Uf7nkmKu5Md
ISrNpH7kLVjh2g0BILfQZ5e9G7XVag8bqyVI2rXdhS8p2QAsJJHjFgJfl7dllW5pN75ozq8pmOFq
GIqxIyY4kgvkYSIBKhkj0e5RdMzzNTa6dn7wZ5JPmo0zDVsVd+3yqXRhhiBk4r89Vba5Jc/epWjv
E3sn2kpAxkybNKDkByz6M/Eulw2cHX8E7fL/Xc/ACByi9ZGLawjT47Jk0NydQGEzEhNJ/Q5F21XP
UaNhfpDJV4PY3sQY6Tcgjcfw5640/dZG23OfIROJ40eXixAgV85xDvW/u3PK9U4AM4RIGbgI1m+D
eKTur9AOL0XH7ENhngbtIoyo4EVebOPMG6gK/ZC4lu7246mrshOtUH1TG4Saj1Mbs/i876XkbRFk
S56OD61PTxLSmoz5+dCCXH5Lfa+LKiJoOfs5NdEHg8I7YfMkSFALn4jmgLzxjMBLOl1x2TOxkfkk
vtZ8gB/Fmy6cZmebv2k1MrHWM7dFWYmp5fqtaHIfM1clwops9hKa33GcdRSQYVrg5//qC1f4QZV2
jz6lvWEqBeXeLcIIqWYCS6FTU4aD2pV+epOF6mu8zC4QQ99ftfJ3GCJYND1NKJ5s7BIwlVFZNtga
g3Azcj+e68lADh07RcE0JfQcp53MI6P4FHxdQ6rscPa6llfHfchgECxDIHv+dnvRbxJ/lqa/oZkB
PEPaySktbpiP5SfgxKcL+BGiO49/anvf4tpkdWhBX5O6tEnOcMC1sEhtz4ZPNHtGgAdEL+vBP0bF
Of3hc+2vQkfKwDjHD7ds7dQpZ1caMa1dzrs2mhGFt3NYF49JwcpoLfWlcfcvoNBiGnMrIakYaDlT
Hs2tWEbDqJVuzcF9lf5G92VVWT4EvJGeYtR0ghh32N6CgBQKcMs9RA6eZtSUxyxTSk9uK3zOi/By
H4PcVhPBwHqYuh+hF1stIxi7feOw1sczeeu1CR2Bn18yzlwFMRssoyhm5U/xa0tUZS8eUoR8AVWX
AoIvnCmFNRStvykOpyfj2jYRxy9jyzXbExUQGSGJBbKALRWUQvZxFW/AOtFE6IBj8x8QgCGsSCEK
wUQjD7aCWtsXeXMgKUM1H5MuYzQs6jcCompL5Xecj1osSB1oGZtkPAKDZwO3IwhkKvxT3BhSF86b
5eSSUf1Q6LiiZIDTmKXTpxIehoJC00ngy3ZULGUyzCRW9Vqwn3wD/HcnD8v+bYKHUevldhGrfmY3
noa642J4Ed15Q1oc2nZycb0vC2aT7qnqZgccJfi7refSK7i1psGrFX4ibzFasaXZ9PeTvXenqXWN
umkfe1RkhNS3BH8LJeJF9De5+7PO0XExEHlSYsF/x9jfl1wpP9qnE49VwDTYYr7qCF0JgDrhzb7W
FVTE26YZ3/jNcUIOr44ljSZVe319VM/ynh5M9lMPkLS3J165XHa5Eu0of2TSLN0rqGUsk7wsMBEr
Z+6Qwd1/HAXAcjlZO9/fXLy8VVOI3wR3TezZMWxLSptuAuwyxmunMdjuv0QVor9s3N+AfRUedJFF
1kULYb8760zAHKnIjfLKGiaUapwZNJCpQX3nZHdS+vFbJhEQLBX9RYSJbs1UeNInlLIRON4fOd9F
CdTrb5qtqMQ13uoOS1zWBIvfcefEYUL5LkXXaczodZz7msYQ04gozxhv4RKjoJnWclqkICjLRo5N
zznhhiKW9WU5tbN15chmymZmcyW+O2Gz6xr83Cd03DeyryLwscMUX92ilo9PdUzkCCGmsyGJRLDs
3MwyeFGzh2q9AfxTvFjVNluO3mSlF5PmP+tcdA+oV3eK8S/Vn4F0TGuNzGrtPRDjqe2gsR6rq52/
iQUd6ES/4Y+Ej8rVFIVQ+6oJOh+gfXO/FnFuBkkee4HjmHUmbvil32HSDTu4TxsZGORAod/DJwrc
iQyRKvvbSheS2qznnXkS0sgwLxpqQ5ro1AK14PMDB5NLoZlcvIQ+XD7G/M/9BFV+3tyi6jEihdau
V5FntPJWzgoEoESaClBZWxS0TkCgEWbNtrgxclNBNfdJeAE5ExwVrBgL8rFI9Zn3YWiNrpMtM/oE
hhMZOEK7l9JUeiaptMdwUqOH3uAY+F6g5o7wVCxYsaKTiVeH21kZyLZX86TzUND5pqPGpXz+Gi3b
vhlzpPZ06YxIth0l6awuqEltSweDw4+3fZXcAXe4a+/wBqH39orourEh+Le5hAahG7JC1vcifTkK
5cyGL8SRYAECFgA14V6srekZFkoMZA36xzwUNHk/6Nf6tVB53KZhpJgrenk24vockIdOjWcw4YyL
ezqfrgTW1fcaJDuyyX/elRLALZ9J2Llxu7x0swOAkhgJpUz2ndJmcvHOu7zKnGTMLWXFmxUHUMjW
vTG+lfJrLkyNlsuZPRrwGR4SMoanfvpZXj/03WEoVrP6O6XB2myG8iuVz+PGkFRB9t61YKZ1zaKw
ewwRn+zNbVva2XPD1YcHKEc3kNSYk8wRrNHnNgeKr3plUZAxUxzD5/XKSXKIsuhHdn6D4AQ8J6ti
Y2jSAhf3D3RDalHMnaN2VbgxqGuLMj5+Z5yHbvCsArAfyxenumU8B6qVWOBqrdpEePqmzC8D094B
Pg6UEuEZhQX3fqQhyNfUhFkdkTFf6LrFtQRzrGGU2xrGB8H9uJl7tdRDSsS3DFrf0J9kA9SH+aXZ
qeaVSiFDFO5tGQKtSmcst9Nn29Fd0QXtzidHQkR5Axcbxb8oJaJZqD3fFYH7RR4/sJjgpUTBAEXx
0DH2lLhiRHAKSwXS8fFMHvwvbmFm2CwdMy3eXP2r5b9IOK3alY3/DDt2Payj8PS6vTKv+p33dvq/
tSR1TX5yaX+xBCj7hboC/zrTzemx4wMaqIDbIfrrE0k5O6DvzKnP2HVhqasNU1JnwEpTkC0nz817
0nPuiobTYy6I872bwlVWUhixHPWJnBqxveaLNSNK47ysLox3FZ9H9rDhg/M3azXPBeWhaopUfXr1
5kkRLXy18EoK+t69rLltjxv7muud1VVEuVqMxjx7wUiG/IfVtCPlQKxtexSMws2hdyQuBiYO/UNy
8RL54FpWNnDe303CVliYEn70Jm6Q7AQvr9ouqQY2RpJ94cQFl0RbL2tWKQPGG7e6oH2MMAeimGEj
X72OGc/YV+IuHlXlWP6O4B1xieeeFYoC/VDBX173KG+u+9IVaSeWcBaXDMtSnso7AYbCAj8jbJ8W
EIAlZnh/L9zltc/3h5TXhA/p0oeSv6ZJsY+uNRzjerHZJ8nF9gG5loxTXOUcn6hs1whPqpE5disG
GSfr82i7pHUyt846tASHm7v6T+mZitsEx9BNLkHjmog3pQYOdazXZtv2pPkP/43CiB2I0EkM66FP
xwH9VBPzuO15HdRNrz+uK8PUa/Py3EltxYcb06D6qAe0sZ05LNBA3JlZPQeLDqosfetZTsnup3MY
IVjgjVpJ9rh9Pyv8SRClAyaRBfw16u5H3wyc9blbdvYdRYy0zGKF5pXrF1rhkrWKu8/FGyZssuoe
XoCsbIoNBmLeefa9DD7dW48/R1lIOP6Z3gnczjRbIEmK0bNiwIsBoYICWt/SgL6oyHs696fhzMlF
ldCVAui5cFz4bd4DBuaOpnI1EzaLBAdIVa2nCEGEW8Dk6knOVMHR/6PWZZcVj4zVMwfD79vp1S7K
1dHAE1a0k5xWfNTHH7omgc2GSb6aErjKbFQZwMybaH0qMtnvKLMxmBrlXFVgVuurGfSWDF9i/krs
9I0uHbGZVskWpyxCyV/lN7/VFmFbQx5MB9cxHAIFhw4ij9aYeQepAA6wgba5RyiPUEId+18ikURN
wxyZyM58BQV4kNq3Zf+UI8pZxIW9rMlGcFhQ2nYne57g+1UJf0UdTtX/Idyhnh7B32sZC/EYYowd
Foo8PvmT/o0doJYOBXcMkh6wHWqdtpoLxaeGQ5esVTJ7Tci0fw45UgrEB+cokXQ4zDnliayDy/Vw
StYYRpuBZZU7TlxTzu1TCRRXcP08jsM6ByAN5N7Irduy+tQcs11Z2/6+v8UKowrmjEUhaN5mPBF4
MGNhSqfyS7cEKLtchCwUqNI5DmzM7ikD2j4nWmSagsEV66RXe8hxiGOyyh9Hizh0gRt/F/Wic37V
tFx02EqtKn60y7FbnzEGlnfxQSkFc2vKX7HgMik27AmE+n7ohgFgIXICF/VKcab5b7UfsxZPLDRi
gVYZX+oUn86nYiB9AJg09MrhfH+fdwkzhyKb4OgBRzoaMipFP6YsILNeg3TY4SyBQTeRPayy9Pe2
5H/RrV5zrkSraDtDGyhLdBCtF+GW+LmDcMDv6CVT7Hin1AgcD+23mYR+/WgWtTOEi9g1Cha8SEUw
2QE1M6IwhTZZEkG4AzY9fiaEZ8zhyHCHe/QiaFNpSgJDUW007yk/YIyt+6MQKf2Ng0I6oTSRpa00
+jN+QJtk7TLJ7vIftg3BgoQGpoD3auyhitQuD2elL0W0Lwci44nJ/Cq0PfDGYAcO8njVHJ32rEyO
Fa7o/WNBMldcG4QqvQu5iCncvvUi+vZoba9S4j2bLBhNV8UNy/CFaHYcNnka9B1i0ervyn49plOO
KM4RGnZatPtezqexa+li/ap8y3iO/3JJ3J4gd6PA4nHticqgwF/Ozeu9Q8TFL1XYQ3CyQVYeRTLv
67V1Uih+v155z5BnL5QfDlipPbEnlwksRDpHGJnavq3Vo+Ku6wYfEGZCLlsYBRvCLUbmfcoZ8fdQ
itGtZmR28IsjHvqYTbQvBWzIzNH41X9qCSMKJfEsOuy0ISv8ZQgX5jdOwXC9ZObZx8336sZdhPVC
wXluqyZraz+L0HkNMQGU1RGEBi9+FPVonMTm5A2Ls0zZetRdxSjbMD0rdsLwkHtPdUD0unL5qqmi
gtci+2ofnzX/fUAWHFAdw87lyRN1IR9uvtZ6cG48JHIAUpGvHcuCrbf3XkzQiFL82IgVc/cacu5j
r0PGjnF9MtW0+RTNm4Ka0kZmmDiJ1/GxarcyTXKAgWhLKrVzmr+or4zDmgocolopbMW3F9o2in9R
JjXCr7SbrpayPftmCr+PnD8FB+/aa+FGj0DlzCcK3650nH5yFHO31+IUGM1jP4/UbGU4s6O66SZj
hLkBhE/bcEVb4h+8Cmdzkdl+vhpF25lD+SV3ykCriCgm5lFBMna8RF2mqKwfaADWaBirBpytN/+D
lafhxCS+xUJqWWe6RThfPFae6Qroys4gBAXeohq7hDht5/lI04t0QGTbMahExLG9MnQHTct6WLS5
gbpt6UZf8kKWznCODgDMnXCR7PVFTles550akX4J4lIpuqmtNSvxpoVqJUYhpJmOnYp/yHSe8wI4
ruqQSvFiXPfT8T2q4eqAiMTfXU/1I8BCEpyG+ZcnXjdXkMQh0m2bIih5bcGy7HB09khq6JZKYQKC
dinyOdPIfZoo5g979Lll9i1SpSrcG1pRGzTBPXwxUKVYKsxD9N0zPdBH2kqN9mmRpUC5Vv7oF+uq
EkvjVda/8TX7BrNe3Tm9qloE3rNk2wX5FY7R6TVud6xactA77IDQp8AIooRIZ42+4ywjb6mWPrju
RY4KtrEWkp3Zok5HxvhfmoKqLHv4cbIvB5Z8ZtRRRfqeSh5QGywzTepR7AWhf+czOt9ISlv/WaEG
BvGqBMGzCXedm+ZaLQyVp6iY4olfpQPJJipDfizcoCbG4KQmZEnaq+Vigr5vsUFYApT7L7wsKazJ
KdarAz0s0eaSBPf8avOTBI/PRvUSgX4V37B+Bwr4ADDzP73Nd/n7NTWXs9poDZekBqwlu4USeVzQ
mHpCRzKL8tN56lb9z7SIwhLCrWNJQcZuyzV+vDFqAD2q2jLPIipG5gE4ywcRlV1K8C1zASTObZdI
X7bozDcKa0esmUVdAj0KKRxjcFAMG7y415QRDClO05YAnTWd4DtF3RrQ8w1Iff4H76C4qVD7PLyl
YYPiFGAXMi7euWB5PlpspK+SYN0zYVU2Gbcoe6r4PbeID6dRgPpUr8h+cowAoAsODWlHNq68tKQ0
jcCk27/9Sbjgk4HKQXLQbcWVMvypE3HUbBtmOs4m8Z/NsjuCLrUK1j+W9SY8/2/LZMyesmU6XQ2i
x3t+G5bsIWzO1qOBAAuCm8KxOfuXxfz42aA4r5fUG7wJx3wxXe8Lj2WmFlyKY2nWL84jNFUD4YUI
QLKaDye3o7PBto0TQaTTXRmre5BIoGAP9MuCMqymUujtf+cVRE1OVffecfcrt2uGQ8Q7LA/0feOi
8ljdBR4XArMDmqy9oimxpe9TCrYOI1Gz1x7+T6O/G3GKcHoiAeng1KY36sIGR2YHWdhpcIKXiVF/
hb4v9Obq6dkjaNh++kt55wNkEjCDYAZyRaXt5gjkgYXVVhIGZiKPbUBQDasCDdE1eOkETloNSof/
MvgYKptsYzrzeUl5SShsftbXvhzEfdOZKdxNE+trvHIj4gu4204GfA7Bwwe5h2XIK+uAdlL+OQZy
51UGxH9lZoOYytPb12CAZEuQpwFMnnX49ZoUDp+YZydCDptuKZuQBmh3wy0TnWWhcTsh4KoxpE5P
gUdNKybmdqQD7WH9mmxKvNNIIGaKQMV7SjgxYWWcN2Ur4t6FcItPx11cY5H8maCT9u35wGXtinWy
iZVguZAgTb3/F0FRW3T5v2NBximFsLxRG99YB+prI6x5+i+sDQUIh83auZVFh1a5rKQB3em+TtUD
iWJgUheVwfnpERIJ0KUWU0Nbh6D9tM6WUOE7Bg8G/1/1JCQlfGXZ2RuIkEOZi8BAs8PsgKYFOeo6
79TI+hyuoiB17d/3rByczhq/14149CcAaVHrqSUDaRm6HXtTwhmSe+H64uUryqqJOJunOIidOglK
vf0RnzPzREN86LsjKMa1FngXhaCTBJISo9EdeJ1aIvJOb5Z/dXMBmZibHirQysb7BK8IdkUymfRX
M+XriJSbs9mfCwAH18lAhA5JJLnFryhV45OWZsrzWjeyqTDb3Kqty8qiusX4zCGnWHI35TMMQqT9
wXodu++9cdbikk/0Z6yC93Qs7GxRnAwyv1ZM5t9cgkNR5jZW9bWjs7FfHbifC+u/HlH6SRxfwj/C
hxMYm3KWswt09dYcRuCyB+G/Q+0ORcQuFvv32PSb3WSsKq09IEIpYuMDAxxCYueTBhkwQqVCd8eG
0YLszSvxLphYpGw++BJObcOZr1/Dzg9huzr5IlN2zg3NOD31k79RM9YE9FQYTaU3iJgaJ5Gz+87h
J69Uy1uAsVUPlodsnSEEHueKAOffnh8wUO4A1FJuj0SQDqoJAsWC3vsnxqR0FVnV7hiOOxn2LXXU
0o4aKcoDXw7yiRVXmB0boWVZ+eHNqcfm7CJUXwzzBmwT6Wh+7EnFrkRYi9YCpO0/6GLYkJDZd/Kq
ZsC1sc41Cy1EM8ZJHfyhaXOFO8ADHWfm9x2jNKdlXwfd/qr/dFv4NRJW1kJ9SflkzrpJm5lMHRfv
dj7e/N5I66Z8oaPtlRmiqeNTvX1tFKd7Bas3sV0mN6CtYyU3Y/7PZUUC2f3jKbQdqj7x9NTkX9Ux
gpxSitSSToYzdi0Nf7ERmt/rQj3l4FShD6qUwztA81frgxhsiJP7ZtFVdruNFIE2vvPFOC6hE2ig
zbrBV5+1WZc3m5yBGyjehS7vPb7sSvIVOed5kX/2gsZHJ6RFB9KJkX7xleiSOAIm8dYp84gy8Z/Y
4KI1mZIB14a3hAHRaUp8Rm6Xoxc0d9iDs5xiw5r1frHH2ghXUv+ZucmmgEAtVicbM4ZsYqo8XTDc
mMwifGsIjbjb2Qtg5iuXbk7C1EcqwMKpkD/oJkmRdKce34pgQY9HcZNVBVVPGXf58NaW0fpHV8nd
IaEsAICDytT5jhuA4dc8mgjRHKSUhyaUI915Z/70LECRtM05xUMopm8hyWheC/Gm/gA/ucm4/meX
r+cFRdy8aeal5okeAUY3EWXxmbHAn/lOFMMfoq+QUm63b0PGuHevs0XxqBCB+LI8tQD9R6EAFIGa
Q/+5ct94giA1uo04L4Je0XXuCtvD90tdUPOSmVX/Gb214Ojay7lBKyVru+Qv0l+Z+lD3MUwpKW5b
j6kpxnmIt0dvQPkhhKMdyluPPMmJ68/bSR20cd7fcShWvyorFQzHHoDkJj03qiZj9oOy/a4Iex+f
HexnjAAwqObwQQVbOn4sI5Odl2ET+7KIRfw/MQA/eCRWOJif3s08PXKIj91K36mBFf3FkuYxGwXF
xHlH4JkQHhm4/5hf0023H+krabUryutLpL/nO6iQ/z2GA3bR9pcGMQwRizNLtc69awfLUoUjXn1w
yUluUTp4WH3Q+oreF67eYFkxHMXPb8BpuAdlYL83+65jddHUqdbbY8s+X7xeYdhrOxq43hKkMvxs
fYQ+RUAfu7BPyfsGUtel2Vs1DMWcJpGT61cdxLWSn3f5oMrtM9fLHis8IWPKy+EUh4G+9wZRdyNr
Z+kKQFr6NK+WEzRo1gLUpVCepUAQPBRv5wi/BQJ49qjxapyJ1u1aTO+L5kt8+t5v38XA2ZDTUZU1
uAsUwK5c3W37kKY1zs58HnTSYmUCy5NV9tmsplFK+jZ+t2fr1ZeNPofs4jn06F6bPW8Sa4pDTqjm
VvGqq7qCAEm7BTx89fB1PN9RPhoBOWsZL91sFTDm2NmveEKW1gPanOh6Dm6JIPOSB59Y+mmLb1rt
Ht7n3+9KwXLMv+UvT3lmGgXOY45CWLzz6OUS8T17iBZDmYOzm217linA2qMXRXtMq3GrS/tQ/hK0
4OeVOoN+ACgUeCOt1lmgy0IwrvjEx4hAqVT6R7wgHW6vTuCIB7iASpUhzU9gCnj+T5axeq8x53YA
w5GIavvDRZ03uRB7HNWbvKAm9Dzf4AWis3bCUyOALRaH85MruU51on3KYB9GM+gnWRPB1k+Su2Co
n9KGJRJLvpr3npRKxYXExe3Ux19mZwuM0GAzceZA9OZ5kXcvdQXMxWJqGXId5T87ouziB9Kkh42t
sZoBPnP6Cp8sll6p15dRzHiUE2/JSW1D37vBvWyfNAd+lAnSb32BVm0sfhZPHqk+faaQ3hfoaxLU
aRNqGhVWQ6khjoGeON+NeKGaN8NOXZ+DpQSCSBT0y8xqtGFRK2L/4Nrcv0emhV+lC5kPQJxcPuwx
4cvVcxumpnWbGOscvpeP5d37cKHqb+YjiFFQSQ+shsSHJUTgGOF00TEkvEUCL+rLvvksG1cEkyLL
hD0WKvLrywBfjupjE78VYLnIgztXGo4SFT0uA6Nw7/2pMck0iuP0aYv9iYzHisZus5k3/Gi4Sezi
WF4FYdtz2x/VhIuLXl7gn50dJKakksN5Tq2TSRyVH9TpRPyresisNnDk1stR+EGkjp6duuVAG5ah
VDfboXTUOMAK3iwMAvjNVp2Iiz+yH197iGRTRY39zE8g5LLViK4KY+oeRAtYvy2kpD4Mq1aNsw1s
XWsE/xRB0NCUiHV9LpKjXGB4gqtpzEiNP9d/dBz7HlUNFukNjxjWEN223T9NGYuSqt00OVLvojQy
sEyMpvN9x3NE70FjDDTER7hAVCmJbO3cLZGf5itFgs1aKNf+NKjetoGZre/2kHGp1kHszaJDFpa5
yuwlpHsGtDjw/WvwIsPtB9KD5rngTe8F9rwW4NjQHLXnpESDXiYA0o926D6lHrHouJSL/0C+G16L
SdGBAUIWWsdy9M6bvmJGDybqyQPfOGN+LV2F8KkW0qg1BwMVxEWrYMjrfKpOSXSxYkA21hwJkBD3
pkoG5iyTWlwWLRgzMEt6ql7KgMYpXAIinKnGAGbRW7jcNf3sGcbUVAmTMzMvJn+9gSNZNmBVjsvE
A/6zWSwsJtyie1YSKhK6YrGlmCFMLBwfL6OVlPdsX4vMGlHz8FJz4c6HD7jC1+p6wzO+6+xr+Ukv
XQJPaqWHwGJ1+phsnYV/mrs0veIaNMfRZ3ggyFVopypqINfqKzA1OtpHBQHg2elJbv6Xlf5thX/6
0ygD0FPI/ITCF9f3GJ6a6M5R441Bbv2UHPPepebBP3quxGfmEIufcFZdl4PSmQ9GVbpTPmUzcxW7
htWhrEI5bB0q1gRikXjbitaiDC2qsT0RcSWpzVe+AzY2XO/6CIjc3KnFzATQc97JZ430hRYgTgZq
iLSv/VCEyrtDXgk6xhW0Gn9CquhOUS1vzxT7F5hxycSQwJGnU8r7yZWMItnzazf89a/Qdfql9Y2Z
F9b275N6qbe27ZrR3cs20frSJnVrAnKHdzkTOsq0QeaKOfY7YOuUTf2XFbhgsUA/QXb9TBxYU/Xg
LBeTzQiUEKUv8VPnVGjoeAGfKT9G3I7xksloQJMfR3TPtPAGRDl9Lpp8oX93uktHVLGraXMB1QdG
XTh0QD3RZLbWrejHsDYrPyCno1MXSf5MadDbaYKi49nJMQ17qgzefFtvPndg7TGfunNbxXQ0texC
5CTDTAHvKkF78udFboxmnCqtzrPMKLC9fk7PEZPobknFBVOvPLpkO+D6nqlMHB+sXt//pC3Hpr6X
/mbLix8ISd4axWi9F6vFfB194oTDusQbUOe5hTnx6od3Vz+tXS8EhJWQLU5AyVXBs+YTglzpA/3y
GCpathNtrq3O39G+Zf4fI1g2V/tLZiR9vvVujNU7+uIsWaERcjU6EtkbGlt490xygTF1gtANMX6I
wgvenVZODCWrlqO5VyjEBwO2c9Nr3N1rlJsuZgY4Qr2hUtUS5BOoASqDKtXK7Lzl+OHOlfep3l9L
qcko461XmOkJdrjRhTlJVQcer2jaJq5bXPVQII5GKkD7Mgw3tfNKxCzNMGFOvHK2UrL8QuOVi301
mg2V8J5PUzXg56dwYHXk7v8VdU/HSQsZRZpyGuZjgIS4/3Lln6fvBVmmEE3kxKjT3S4DdVWQjcRT
5OvopFbspHpXl/cUDKOknbMwMXkhy/xxAr6srZdsqXMlHdceEiSdD555gObZJy7VC5nwxIYZzHb1
seXUh0VP3P4utdt745aNgNTTv56/toitwn1TE4pB/erLwYwpmu+Gihu+ebulDSGjtmYLHZoVBlwJ
Yud5RVA5C5fEvdMRw93c1QumE2axyMkKGODsgjRvCbTzR3p4SKe9Ivf3h/vII76IGG9hFaZTt6Hp
qEb+Sd2Uifron7t4gh5D/lMV09udZGT7L6UtBXgHznxBIa7VALspyfPxMEq7O4FHFWEU4ossQtS2
Lc3hPpP4DZHWNuQqmNUnWLdiDPPxntx+gKVM1z5J8J1zGVp9Gz8YGtpA+EHd71owsEdsya/Ck3Fo
MWlWT7rryqMF8gGICH64uLwG5JeET+e3mMWVnFGFv74bbO9P6KvL932/GyLFe8jrMmYeLQ7Z5k9g
CUMmSIAoROUkc76QCbypfqpv61cHaQgs3K8hHs6fgYFa5qF2bPYgpneS2wZMqkVMBNCo1CEzpSfB
KxB0e7rKni+r3CF9h6GQ+IfHkONY+p0mE1CO5Y/DjcGuUQSNZfdocRqhVcxkJeX7khJzta1HCp4N
t8HW4GjfJEkzRO30q25xIHQ9RFo/5MPpZYMzZUSZS8XnL0EgD5N2lVXpJvoAWFJSgWy0T/PRmKSl
v9xzV8kypZekL8mXVCpcP7etuGFQlXptwTmUjPirJjAioF8pVtj0+hTmJHBPSpsJaWiMdlV9gjrJ
ljG4GcxuRIr1X2W4NA+7iNGvChJiCB/RVJCYZbQpi80VC5MKA9MAoEXo5hIReAI6s/pTA0SrDiAv
/D5OkfELKOw+vOukwYT/lw4SwI1iVWfsZ3Bl1JHAOYOpYRABq3Oz5WaUocYBJg+QR53NxtI9hIyo
TV+OayFB6JclBV+YpqpchrOWO2c5Tp91TYhu1SzTVfe6cXymXLEWMznA49L6N+2+VcY0ycSL4E2j
3KAsX5Ee/LlBdyud9oBNHIXjbRXrK4zEw3dSXMBSGHeGKcu2v1nkbIrK46DITZk4/gJ3kG5pLtny
iurf2u+eWMrs3PdJMrYDG80/LGZFsHWju4+bpceP2ynaZNLtakkeuAoPb8Auy/L0MmixzSWzi6KR
oS2/poATJfEcd91vfN9pGs5NSy1YlXB0NfiQMUcr2v+4v+GCVGYm0jst4rJ/Gt+MZg7KiN8q0A1R
zOiQLVl5oeleXwFYDUC7tVccVpJ9bJobDd/O3Z0yOUnIstJVxMDKEt9c6dhkWcZK4/poE6jpFcNH
GthugAf89MazF7UX2VpZYxpd+9gVTlidgtIGt1zVti7ugxa1YKmn6prY0Ht3P/OXB3oYJWB6Abaq
9+hAlaqLBGV1CY5tOdQn9jgw3u2Sb/UQjxglG7c2Ed8YEeOV7Ub748jV+i45z/S2OUE302c515EB
tRXT3uC4d2JNvdIsxiyFKTHiILbCUTXSisuafY2e7cXV6UWzlAAl0tiLmbFu+Ac6mrCyCjbPQSPD
Psm6Ym20dMiAua6jE1js6VZKOstoqSxR3HIzDJKQWNa8cf38jt5N6ZiUaExPwIhkVl3fjkN3oPJO
RqsXEwkZdrCY7q3j9/IXj3ZHPQkhnUOdwGE2L8Mq7x21Wqy1aX+I48p+701IVZXw9M6AF74RK9FC
0kGUyxTZUA045724ZNSY8d899UAmu42BmQhLXR3S4yAk9v5wPpaUuTXvVEJPBW+VWrA9h7ZWHtDh
fFe03VuC6w4Qc+aGGgNVN9E/CcAmfee69WwfSOHreHRFfdMMktTcJM27PJi3cpVIAZCKT2TZwU00
nVqJwb1bo0vByTyT8+B8WYVZoaB9BfD0pufcbXvQ4KxwOehkJCFaGaYS/dL8A72y7Wh8jWavboWu
RLF2+w1ugMvFrfSIsNypCn3sUFa0zRjO7otig07ARHdhQyOj3cURBtJIMfsj0eedZ2clcGkPTOfK
3AUrIlm/dBqOwGWNUCwbkazMq2ds6Ct0RNLavzcg0IgteeUJeZNF/5SpD/FOBgCyDMHlK1gly87Y
mP5r+ZUFaFeDI0w8w+dlZb1SZPv4vAfVw1INCYAb/dFbN/By/cSFh/Yy3FSySJED4YKIcz8Q/Fe9
ek1GX4ykPDJpRcDrFNtI3fGFmel+AmeOC1Y7nreY1lPurF6HgSCVGZkopA/FtufW3/pAzbcgdtfw
Q/LzYfADYjV0cwwpfeG+5orZCDH04dAUpzM9HjOQIJSAceXqIzmaKLNY+NYBgMlUhgti3NWeAKqJ
1lOplM/+nHvGzxlPpzBhcQHnQYYEeQR5OROjlcYy8+G1aE6NHA6zQej5SpcLpkNj+qcpmfjk0k2A
DpHxi6L0NxnvRRKqs+p4Au5UIgruITBvT1Ljxe79eJ864huBe+GzP8htAiqfS8Rig8E4lPym7qjT
fVjpLVEZlf/ZKAWn69/hgWNs9qHhFCDZb5EcJ59SeIAGO+9D5CqRwrBdrRkNYbmiwfWsn6uhO7ZQ
T/XyslpQ5xQXSwGcXTea3hP6sDtnH/oKOyGdFBTiZqqEcbzsqrZoYe5eYsctv7TSPiIsb2HfeFaW
yqh4/60BT4IGXAMA/5BuJyHd3RTd/SGivLcER11Qp+svhX8LEDv6Kk0n07f9pGTWlYO1bJlie9M7
MMYaew+X7ZHhV6GKg14YK7kyRxJwy6NWR6XI0SXKcyP4Q7IKz7saAYjdIlPq4nx0h0zh7ArsxPoq
W6ZkX17MawmwGxT1exuHfOGJOhp6tGQPers5YJEq9K/yH3yR858tCLC6UrUQSFNQM99guH4xgoRQ
j09VOit74lZNvuEfvM5XcIyVc1vylRmJFKNav3vgnpWfyrcOX3DYexbyMRkTQxMz4J8WYFxaYeMQ
+1BHefEzCqu/b7mWFmkTtR3hnMJtkKqj1FJYZuHci7Yy+WOBU7rU3CdtSGatGF+SSOPDBuo1ytBf
aWkJOb6DW+/ZhGNIYnT1uqx1p43VAhyLQk244gMxW847pIyHpLejSfQyADsFthbSEUxK7XLaP3EB
0aNxTOmBeArBLWuXBEnHzTqFfOKu9wyIQuERbIidcXAh9A1lUATzG0AvubSEWpT0JhvtauHkag9U
dR/Jcsr/imX6PcuHoKAKJQkigXYHuuChDoXHJ4AfCIdYcGD97Yqd+n9Jf3JH9zUy4pK/2eEQK16Y
/55ThdeHByr2P9MqRLHDwFmffGzwwld16+sz2N9UJNiedU37kXeq9LU4NWp6n7dNQ0edF8prsyNq
wYb5qBO8xWJw8bgUowfW2EyXCdWnemOUJjynzerlFDnhwSkRAC4KvWQbydg+RnSoYiHc/aCcsQBa
7PXB6H0TBsKz98ihvuyBq+NArLaRGJolE0xTmFU9xBZAI1QzLyYSH1VprX8ZxkTR0eEDq0uUOblM
yaaxFFiTLyZTNFZUGYaM4puRZyIDpS613rNe+J62JXwWP7tQT7BLBA6iEwpFNmMGxKadja5x3iqL
oYa0dQlU8BOU3eCCWrX/HVy2snm7Ys9OPwovvPYUrWslgPvSXbR5275QBcJpdmwmBoThkeBZ4WOm
Y5qEbTfIpT4aVoWinrqIrMa6wbrYns54cZ4AStymUOtAHRELzq6d9kYdVcZSXZlLeLXuxtp7apML
YUjz+v/9y6NFCuCr0R5ufwEFiIlOfRxlIzJk9AZn4dUrR6FbAkKJxtaVhgrv5+gRAbICVDqsp4zo
Xn3QIBzgUvZwHi77yJ/8nTYaDiEprZlMFKXHHYDgkm9JkRn6eNlvIlEEjKT18LvHAnUuz65AMG1Y
GaheULwSdIqZChxlITm/oW2ZYjOXssMCOH/75POfFBBcPJWOEHqIVJfLljVr8VYBgjfZaR1IKeD/
GKEurx3M6E5PxmkoGAgKxBZ3e5EJMOZeLHfhij3rsjDegCdKFxVJh4qCr12OZSgXOrNhg/gpG52n
zRVzIcYjlzzFY7PujTb+xqnUfWU5wwSgNKtq/XjRoGs4etkY36O650XH3Y5tm/yzyuA4kYOH8tut
2Mc/0b+cl1WS4Q8/PdR2nXNnO+fls8CR6jiRjO/epMVjvwnx67cx6XF9pC+AH+bfBljtM10nvVVh
WcDMO+xUnGnDwsrdJM5i+8IS41+cY8OJk+GrRMLNyVYlAQdKANXBEOpvfDHzKgxzjitS/88g+98H
/fThXSy4UMuwM+uIcisGjbYGIF5sB/UCNQo6rX46eqZSlhFdtMMPmftcF1bzc17v7k5rsSN7DPhB
H+IxNg7ao5JuoIoVEIiY98sGl3ezoC/1f+CiJYIUyAiCPzw2PmpOxCyQcAKTQOSPTz7lAGdMx8Kd
6mswRPo7Pl4E7at1KTrSxuxi4RsALqrCMZ9XsMDhRjGw7mg35RgS27sNdStzao2qzOEXJweAtI6h
cA9kJKoZAEAB19keFGaKvYESanJbiG06iafaQwgYZ9S0j7bplq8z0TkEqNk52qTs9dgWsYPrqgom
AkqWIUr0KNkW4eEbDd+2putHqVhvFLezaGuWXvt/NDmCkretVc2HSmenW+OWonvwX2gzH8qeatqv
pyONzUSfiOQbREZs40NBSXB0G8b5EKKl+MiLsWQ3OLYgU8NtikGFKkfbO0vXEv7Y+C4zW8WJ/LPY
VyXRhDfIdL7iBG+F5q5KOvk5usLy3iSNqPI0ZGLreMZHMbP0wuOA+qzZf1AKSoL3JOCNIuH55hy1
L4ME1wlY/7d99mQFbt5Itaw2E5PvuRtwdPzsI/SfGemrdAusB0vu4UTvEaMsluDRiPGKH1VJkQDW
H4Lmkh0hxDjmpqDG/0VYK02T1jqHA7oeGDrg2zlzfMTfA52VXYWWZDdvsJzjyvgQ/cNo6C/AjT31
+C/h/GafX6vsVwej8v/2k0FPHkYGY7NSAlbF0+tOa4jw/PSNdvlhHmDepxg09e1pRWmBQXLcbpwj
YhHB4E1fm/MapkG8Ss/U5MmiO1kNL9O7NipWb0AXM6c/RsDitjjBE/bCKOrIe4Qv9vCMmHg+D2pn
7vxdxmi1RISPr6v15/QR1SvkJvQXzdsshITFOhs7ZH5tGPRCDMCCPVHFDHb62lDwcw2Rb2nLkAcp
sfzIG5lzutepmktP5M9r7NI4fYCPfCWbzWVVuZeAS8cgnmGRf4sJ6QVN3SPemtq8FkEXrR2/bOH+
qaBUvheL4+IoFx1TtA2kugTwyCTtJ0zG1jXvOLK+yeOm4KFJ7Gm1aTKMVDpsYDrEfCVVcYvS6AU8
cfM9ZBnBFkE5F4dCfKigltaRXjHV1HjZSJDm5LdE7/uaCoaQD89FrvMBpdlRzfFq/arAkYHWimg3
RruTPDqqnYJaHe1X1ckcLD56GtCxCThZ4Gnaxqbz06pbnYprVUeccyL2+xQZyjqO+U8DUlGBmTa6
zwTFSjZpDrJvuAXb7oCRQaZkQ5/6Gj4D+hZSaZl9sAXgda2xYVkbAOPhttr1bEhpEviX1n5BU4md
H7OHFQhdNVC0ir4ks+5SUlVojCIEEYmTg1neNHUKKgLYqddSvKCJ9EyVb8c+LRd8bHfKTvJeVJi2
0xOcRuG+eMSA7WHhADHboxNMZcCTWek8eqskhSkxVZ83NAFx0WjbTJrpW7ViCjh0ybB/mdwwKWt4
tPzZA61xL7BSNcgPXbd0aUVB3h+adHiydHcszCC/O7ztDcIKmngCSb1bdh3NwDCNUFL6ENC9SJ1W
Sh/a1dG0VjH73m9mE9z4HnP46rTa77WknmOHoSVPz9oYOc3foooOgvmFDvel1VvtcmrmFK+uOa3I
SPWsChUl2zgrZvRJuC7jJYmWYtpbBLvHzixCEYHuwZnaVWh9xekDHd95XpqgtVETYJ8EBdyRSKux
ERO7PiRwGZSEIcMCREwg8hh8lLuSq1+IJIefaoHNmGB9AZWY00zMjVRYUB0foo0vQN5Pxtb9soQD
/aFi3rh4pElJ1dNv/CEr5weEdoLag3pEp1GUFsOE/pUZNGqRkX+7zMU/feIgzrWOjgfVJVv58+Fh
AXAK0OfdAnIpMLvs11brV0WQRZU8K/8SEnFag9cz5MULv2p5HHmr/G4zZ4FTMidp6xDjWbhVkN9U
zDr1zCqWm/fmdSksLCP2IIkKAVLDAvH5CpnY00qSQF1wxwrNMCfwljdNt3ktGlGYJRNVqsPIazG0
eiz/cJonyDgXSzyvgxCgYiDG/eQTduQW+f8VlSj8iphgHDgHYU8NWDue7VGEOYIXH1JGq2WfWb1m
UrDPLkctFR2PJVEmOfdJ2N656GhsyY8hH8RL+Wtci/qQWB6p7ICjA9s/iIzGklR9Vs+CLinant72
dX3LQxEDU9c7NP4xpVZZ4RiLXSli4TvqIQKycsmFvkgvatqegiX3pHhDeK2tSx/GkMcdreNlVhYG
pctEQaUizDg+79AbNyGJdHXIKeSyYQMJtwuIkDHHZg1827Y7YVtT6GKoi9DbUiR3fR6GIAYCpq4F
pCXNTHbbVVk4EuarwbUKPT99JXK5JfW5U8HsrIveqqBNgabZuSDmcwq1Km25yTW7jaPaO8nH6WMK
QCkvat+oNhS8ryvVl7AWm9taD6X1zqV4pK+bWhcedXDbaE9U4Ze5LcDZ1bQMd79jIA5Kqto5zkPt
2LPfbq7ArU851g1zoMXDi++CCgvWYEx3Hr0mtYSXlcdtYDbf75nJFLFOaRQ5NMz358YVAT0APgnB
RTYm9l4+r56yEogl10QUm/OP69aTTNdkot73slTO3yK+8tQAg+iDbdM2dTZpmR3PfVMMcSe5/o7Y
4QkH5Payl7gw+0pvk9xB2nGZvMN9AWjuAo2pEZJrD4mRFB5Ufa+PTEg3HHqIVa0LJvw5xqZzuneF
ff/PbJyE/cCVNDvP39CCyUNKI4qvEFAGbKPz8Gff7Qvr9mrDuMQg67cpkTBKsL9jr+OjMSv2tfVu
8SkFlfmDLi/Zk2qVlvd+Zv2RNk/9I1hCglMJsxEZaKDlLxC1qRmJXoeQtDbhPwo0B6v3V//vQrbP
RcPQ+VFahTHoFtZ3ViF5Xu2FyfDQNkgMleJmCNckhEt5mLvVvZs3ITj/QMIm5rEGZX3pwhnd4vxO
VeZ8hza2Rb7seWUeCi1UoMMeMSjl/8vZyYe+7ItHZE22GPLEqwK/KfI8OWi/53y3Lj+N0V6h5HKi
0/c/vNBA+HKbmyZmKA2O6lYMHuwGBfHzLTGpC41l6CbiLm1HIVN3P/dJV4jsGS9bK69f8n2TrPSE
z8Khb/3IygnhJN4QfpWvN51baa4KvMDdtrmOmqfNK+w8jqtVIdLn607l5rkq1ikJC5S9FkGU03ua
c4ccY/vYZny6ZedsczexN2wOfWIgPeXRHhQcRtMrkh3uoIrERxF0Q2SsLYtyfEBgL9QbKJrOFwSS
rC/8TADNqJoVA9SXF56GHRUT3B2J3ecfWAquXoNjALKKMIrKVwL+yNYGMWeXqe9D5X2T0M6zP9X6
/xQma0ADtuJHQ5r1/UvU5xmKMEgNftafKNySCl5C6/i/1WjEzKpnAmnMhN8JAKU1NKISZzR3JbqX
RcXMaApZaHZiBY410+PZQf54jRjCtZy7U6CLgVtnyXu8IBzYYHGrjrO2JUBKtIlY3/t8sZfpdts8
eE5En94PPk+qbGvRmiHoBrzJduDKLoCkenXXhfHss9TIqOqb1FUtvFrGiNtUA7Effsa3NxE9em02
x6GDc7NmFDEEVfOCm7sjh1l563ZqHhLSxnghmwR79bExclYLLqzrlKI704KwfAW/neB22NUNa6ao
so7WMyUkUs+TT5gi7rXAgYbUOdQCZG7/1D7aLMPGmX2B1D49EBCp4GONOtAsHuIfqkvXiAnzvORy
ABYUYQlMneX7WFo8PFePELdUJPyKo14Kd3gyWbKEuc1C3SvsnmJsIK8/MB45ZMa7jPcex+ysrTRg
Bon0RTnx10qGetBM+BmQFKSQtcll6BMYjImNG1Vpx1GW/Ibs+dSSL1PoDGDoQ4VDx86f7YVSkfzq
FnILHfGbRF1NKDKs5AmtEchUEz+QmZSHsvgd/L/i+wwIpY5nMCzIF9ZH/K/FlqDHXBnOgCMT2x42
NpviCC6N5T1GWcOpvv/CWm5B/sjESQvBHdiiX76Mz0ZJilmJ5VdMJX+H82KOtHoEoZErPVJb5l8A
v1gHV1+r0t0+ftHiMShBbtNw+zBZ1WMe9VuiCQ4RehP7Kwv+hp9JL6gtB4xKY2ZsmpncWnmxlZ3H
bdwfFz79fN5f7gZK6dqPjws/nxZSRWSWP95l8NWJdsnyULJuBwo5XTDd8cei7JV4noJsECuMGt1X
KEzap9ZzkN7fZe6YhWWRwpJ8LmDMoGPPU6or716VTHhYhXEUJ5+RZNjSey+TAc9sxd2L+YjNtpSX
Q3RcnRq7oYI+0i+sx1Hi5p6IBgouB47OAtbdAv03RFs+8H52quo0y/h2RtmWkPFkip4c/Yd4F9JK
uOTNb5dbfU0csn+FimP3gVcRaXkn/ANKq2JTPt1DGMuxg02dlpHB+ZAB1i+iRcQyMCLiLOXLz6MI
mwnQ+5WxOxkS/o1hutZbhgIZxolyNN5Zh3dKH5RJ6EOSkpOPvXJDlAvUIlUUCcsDWdYZpnATafpJ
m6DOfWYWaj6JL/KAVDXwSU6oXCJxFnHZkF1WVWoDW8XQSNBd4OA07RbTqUm9kFLGcA4DEXwFs7pv
bBayggvVgOFCuK5gXdQsOP3fhewbJ5+9NDGYF9zz6ZiCWg5m8YU9UKtyeTUIIQLX48OKOvMxABWO
EC79mj/XhhYfiXICU5rRDN8kPBKCJJK16wZeIuM+Wu6XLSDHPuIfRlg4ciEyJ2blzTX7ppwkTFqN
SP5vLZ5tF9jw5BbFb64sMslMdxCUzetNnt0V4GuBpEciiZST3sKqIGFVZTGYwOMyhDAHoF4d+H5n
AW63U+FYmbbWam8t0nOx51LsFW5CDa+He78Q71BdHn4qzYZNDwEMIm1DVJ0EpnAozseUK0S1MRwr
boC5C5NvfFuX5Rypelc7pU9PZLzo23+4y98CnHh90hT9gfcEtc9ePyH2v8b8Nl125JlKIZX0z9mB
1LOUfQQNGR7BOFzGsdFtq8L1FSg63uvBskkAl4epThS08IMwkwzNPBcB1dJ9wIomz/TxgtegZjJf
X8HU6oz3ELYcSrpIwMVku4xt8cYG/dW9yh5xoWirXZkol1WANCKk0t8JjhJB7Ai7e0mRPoFZLmfT
D1KvmQUQt2attzW0OBPY9Ka0QUpAwNy1pw5xvZUHQ7SeDKZXasrOrczp/XOT6Up+WwJKK5hIxsPp
Kn4u+Q5Vw/wfkFL/83DyB0/1MrSdfxC1otDdYKmtjNIp40lkY1wSKDi05T1jBL/h1A9IYgaA2z0P
dcrOa2mx7ayvVr97A10HLGZ0G+9wxe9mvACf5O8JyaKiHXiQcthEKFA6Rd9iZWbmi+lFHv57H2yF
eQYgIjr/Z2Tdw6uwTjpMuyyxadJhs33LJbReTPw8Zii/XjGpocz0INhTo133pOWMim2bSsFsjFBq
evUpt01GGg0xWbjUUygj0rzbnvIFXwbYY1qFxBuhbsps3/zHvPMfCf9UP7H6Jv5IKEfYViNg4Y2W
V0Nx2C9kc44lHS+hbl2F3kydb3Pq32UHCJKe0D8TKkuCC4I988ppYVxaZwUsZ5zByiUCTRM4zqvv
0wIgYv6bBmuUOEjTSoTRrn4EPZzg/qDyP69sr9YHxgVT9+gLn664QV19b2Z9pBqW+PrMJL/jqm1s
PGHcKr1XFLi8XN3ts5SQD7pBnE6YYE564bHaeO+kGuyiiZYxWJAr+nGPhvQPtnNZjoqnwOOJFLlZ
ehzYaJgW6UHWdSc0IqjCZoChWRXZlgv3BM+JiaStcaT9IBP2q5gpnqzW1RjKb2kCcOoa9iDrgd7i
QuGqjuhx74gSBRLgzyZwraQEYJV8XAYrjmu/7UV0HSLwSZszwSBtnRVRNnKJUoCDtGDZNvs/rfzJ
0zAZ773XpWsBJ78ATxagV45g2xHw1PjYX7x/Pyjt8iQDhPqLpwwGkzTPOa+uxHYCHWc48MYxBF7P
kBaeS10q9nED1GoGtjXmTyySVRBmXtD7M3QW6jeHfOQGJKcwlp3fQbQcAGUG8HnDqkRFGal5qY0z
KF9Fpmm8hFxJfA+qwHnNnwwQCgexO0kgCvUIcjOxJ+37T4Qhtc1Cfnzo0YukQNzuntIbYrCWbCMV
MB7XbT2JUteGRrxg/VWpGIO1qi32Mxz2ECwDNStJp9Fq52XXFN3XZ2liMKTNb/MbNioDTM8L6rZ/
ZK5NeiH2ZjE5IzkffVhzl9oBQZzA+Wpj9fM5brdVtQb16bdQ/kW3hXNwO1hJPPRvWvrWPpu5uxg2
wtTDMv4sZ5kuEZDuQzaiPif4z+eiUGUXaYc5ia281yHWvOf9+yB44JG2EwiaZx1NOBo0LsY3gMR1
xmZNGofnuPmh4I1KAurnDu1cczDfD1+1T+jtVa01YDBwYrNOi7emVFh5aqNK3vzSf1xnqe83kWSz
udKAmbR/cw3IFA//fhXPsQdu9pdW+cYtUY8cay9E5g8rSlUBaufkXfEhQWwLbT5acI4vr09Tgsdp
PITiWFzBgz7HFRVCCJwVtb3uzNHUB2btCwgp+lepsChjVh5L+uwRylWLxyZ7UOpvroue5q4TGtTd
EBPWj5j0p32KhXLafZiJYb7szOuez8Iunu1G5AuG4CSqHjrcHRNmZD4McSTzsjWboVJT9JApXDm/
LL0UkdsuxkDZDHkyHY+FZliF3en5Mn8Sp2Fhw6IWm68jk0KgYzaTso0xm59EtfVBcdqEJI8jFTuZ
3fgKrtDUOG+QLcThHd8VY3vECJUYK5vjlBTnZDfe9JCt0x7y5UZRsxkMJT8FUcoo0Y2hU9qQ/BM5
KG4OR17NDnF2oPGPiqI8A387IkEiI4c1+z3c5BOHol8l+bP1Ow0ARZB0+hYVOgdzgsaPou8LuT3R
TRkcyb2grjVJt7TEgEaIEjI2gxJFXjZjrNN5HN9xPYnpKTT5DmjA3GDWByeox3sRmQvuy8mvBLCr
fHWWaajmHX80i2JLPeA+nKY3IHqN1uKgjllYrUizBTHV3o/fzz3HXxEwPYXU9dQ001Gi28RvadIe
rrrHM3cmeyJTaDKet04vZ1AaiX+NIxrc3rHgRqmeHYH33ZchWK0Kla0lVG99orF2Cf4ZX4tX17kx
BuDiXZkutuzveSBE2NROTCcqe1EmLdygze6qYY04tuAUoU399fbidzL6yB0icFvHK01hPW33Iba3
L4Ne1J8LCFcQ0dO7+EYdWKrhLrLq4zzMoyTgphsC/4ZC+yx724JTj4Bn727OBkpTHfdWd9b+kgQ8
Pm+oZGMbl47rEmisP2dHh8DCxaGLfUTFO38EbMeThNGJmgbxTdkFDuTfbC5hbq3ObnyCWMHrMKrj
u6MAKhz1/SbLk1cncapp2DlvjJ6XPE9mUHI9irIZnc3riaSfSCjauD4LurPknX5z4WmcI/N/PKMr
rROtA6MD8TqTUHmt3/V+f94hJcLUnHTc+OXABABrnkVZcexfOR4oXzIq8Ca6gATTsFAK6EkV21Kv
gEnKUYbay2vEGA9WYzvQ7rMgM51s+GY18W/c1Q0hWDA3d39QzBxUuVnzMI+zjkUTsaEj+Yl5WiuH
sYBuKFgIZv0o4giABiZBIU6cq62BtHb5SIyB2aQzoRhvE1OQoyoUdAHiUH+FWG41FJmzxj+AdroL
yk63Zcui18U=
`protect end_protected
