`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Hjp61rcFB+kjWpWLOV2qx4U1CK0zNOAWId8pzU+G7Cv8VLLL0+1k2N2GrTKa93DIZTpAOXCtZWWJ
m693RxSGAf10Yiz8cX4k98pNrHmAFit7OzEBAmEqThf3eatohv+w50ofV+bc1PYPIxCjJKGwgSNc
dUifZC+gt2toWDyisiyNWl6ky13xG60a7xprFvCuzKBQTiqCBsC2M4sBSso1Wi9GHZzxjdLeyF1m
UaBDUZ0OWpeHqp23icyFmWQAbFOewAKbsyxbEhkM5OBRKAFA+fvVmTNxmFctNeyZ7VI2VMkZ3Go4
xijVIvziVVWn8J98ifGf1+bnacSrhn3E/D7JTw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="JP8hBI7DIGMGgaWS9g5oQhT/44BH4RYbHDcHzlu2xpg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37552)
`protect data_block
mzK2dPELsf9m4DYXjR6+qKbsrG/UMVZ0pD1WSZuTjjShwkWbsHc3I5ASB9ha1iWp3k6ZymRC6BQ4
zeYwktR28u0UtmyvWHp6BVAm3uYuJSBM/BrEUdBYA/tM8tQ2FswQzEW+TEGSLYPivivMbybEgyVm
zXxRrdgpZcLKYz8D5Hwr5owxLysl9SDLZnAo0R+/SshGBbCW1W3iFVWAbcXSRivI1/3+pw1ZDfj4
fQMLpvRiIAYgO0C7ezg9AaVBvvCNomEh8hbA4lTZr89D+iftw45ttoM5hcIkwtVnsXfNdLBA6sb0
aet51UQWC2vkj8XI+ZbsBdUeNrw+ARdEv15CAsmV9C/6XaXWuKxS9aSWQBezf1pPVOCtOLy9wnc0
T+7X/BbfIg5kvJtTKiG9tJMF9tvFHXHVkYnzdX8SSvd+erPZVoGCZgdfp5hBddeN/6o17mgvUsTq
7Ccv6rs3hzg0cuDp2W3I8D+Nd0Mm4znY1HgCgt2mxgORt3TpsgB6YDhMlRDNIZjkMBilmuAyAPxy
5XISpdwhkMpGU2ItNunmFGGpqlPTSE1h300P+mPCigxKUXUFsqwRJZ2Coi3P+OzHpXtd2TiiU89z
u94/GijDTrkDPYGAP34Qd51d/DkcZGpYSvEf40HBIrYzRKxTn4IURQ+q8jLGZo6wEmiWCLvDMlCp
YePky6QFqLv8lpXYhjIXcnuT2+r4y5uopUsMS1dfvavMrU+Gu2OxivLllH6bWR2oQ7ThvXAjEVf1
nMMRjZ6J4OI7GwQee+vRDacWHz1sTfcy6wGqheD70r78jROwsDlSxMpiu4dPJjrdKXVK4XNTMHrN
3vArRA60x8TVosUT6fban/DIlAPhzWSfhkKuO+LIAL4PvWwd2wDqo+whQpFZQYmuCO+T5AHxr7Kj
Z88hvNVGwweME7f9t9NCZWusTu/1PEHrnoLUhS1xNfcqdMnMALe/+p9YEE4Gd5xa1RNu8nCCUzvY
F7VzuI/jXXcPQo7UJO7ZN/K8lCrLT0rkm0up3I1LjF9/RxJhBsZcK3ozKKZDw7crcPrjmrIM1N57
urZbKG/TcKYvs521Z2jSxSkh5/gKsY17trjqcG6JR/2kq6OlSzn2/8fMQXWsHt4Z5PPS1PEifPG3
QLzm/nvbXPQ4R8B+gfmvb/In7bD5PkxuRnClkZPgC9lEWHEy81vweV01oh03CbMvcXL6T6YAlopB
7+z/c+RvFZ3r0u8z6apK395QA01RQdL5llA0t9ZDQzfPI4JqhHM6iOyjFHc6iH499ttJ+AwNfhRA
bx1gHY2uQKlBCtD0hGnwOZ4RBwSjEZwFhLECiWN/BEOlrRVMKMrqfpaulqzdrnCF+KwQl+XMqrIY
yroDIHdaPwD5jKpLzZoEiUdrhACrbKq/8rb1+nt0kbmvgbmvCRsFCxecNI6oUUd6mVM9J3IQBseM
27POtbfLPs1VVqdRXepZKCHoC9xsQpFcZg4JZZ3UMI+XSQ5kQjWsMChcnmHP64+BUKLPDAs9azSy
pf7fPoIEq9JenOxvNbNCy5Z+ne72foOP9ybP4+5P9PIsYXrYRivRHpnRryGmTL5ihDC3NyZTip1n
HkQt37iCupSHfN9xrw2Du4Q6Isc3chkZs0McPaYB7lJeZoqyHYLJnkYic02WuyIGkdbwq8iTgYw1
f6ui2yyT5ATnx+oSbx/Hn7LOOfoWmpogoaEvNT2bX7awW6mueH8b/VKPpnP8AcuWmR55gaAN8x39
wttxA/HB8RoslaapoNVrqO+c1mJh9YutxK3usf2xNCUXBfBDXaEylRk0ScB93fomfq8u5aCF8djr
+ExERU6sHuu/puV7Mbd+/p/omv9YlMufh5dXBBm9joqtBQjfr0zxbzNGLBA6xye0VQRrOcNkiBtb
KzP7ogqQXuFs3y52t5FgPGHKJKBUkOTOtOlOK0KztFmSER2Mwb0M3JvyQqCbgL6x1AcdbBPmZvQ8
oAB2GYm8hv8Qg+fZ7Njowu0EKyVdsvkafGs0tBSblaqCQAyJ6j0qzPOQ5Pj0SppwmCST29m2hq+4
ZTqjr9hC7uaE3t4lplFgIojWGiPIoUFd7sBeKIiYZlB9WvLV85eae4iW+O2yKZDe8JqGundXSloE
SQNdox55Fhu9Zpfu48c/cJgLY0UpwXttWadPEn7MX0P3FZcGI1ve8Mtp3f9t7M/An6Tjz9pgxpkQ
16BiOBV3VD9TMbuTtqnyxZe9QrSQRTgkZrK7CC4L/ZRr3RxtauiI0wrtfqH6RY+DHKelJ6xOKdhj
v2eYKpf7b+8FnwgmnD3dk91q2osC60go95zFgHRDIfVd00K8Jv1Ilyo0/C+OgNeYd1jbfrR7yftV
W9w4vhGGxFakct6GrFbHv/iWFHcdhcIe/xDd6j7/dxdxs9rGiLx8xFV5hxwO+z/ImNnT+wzdOm+y
zkrkkpdTiTwCtYy2/40nxUcFAR9ZSY8ONV9+QpxbsF+GpOVi9Olkajq+3XQJMzXmXKfhzubZL0G6
b39aOyWpRoJNOz7wpRiZxeoXkFPmC5pco3ZLFbmdrOSerbM+Y390P2Mmb74Qvuj1b6fNgJADa0Fw
OeRfxoGgvSkJJCdwZjU24Ew7ho7CyglprNa/XpKFcewhx6211/txvEHdwBKCVnEo6pftEHggU2cP
lS0eW4J7wwDt8GfcF1Kw5MfPTTCfA9vFasGOoy7IeLXQjICRKlmgTXyFk0X6HIVoqiEmo1PvXUfH
br7Y7btU+O7VHOv6vutZYxTUJt77u/1CQSiCSW1fL7qagf3bDI9zLtBgCyiwqalrgGEiKek02trH
+xj1eOg5m+0w16LV1OyXb61fCXEkbX0vcN9mh+n7KAeYOZsMCrsWFSC+dSIyiJgL40pghgLjurvO
1oD4CJsWNExp1RKaYM83aNtxoorlqZS9dX4td3Bgvkc3zbFPW15zqQ36Dl8LlNAHrxg1G3kbu/4m
fGTmq5+LDkF5+gJJkFlKoMxc0N8SSOXBI28hUrFHV4gr+5JolNEcjU0VyuPCIBEqzqwwGM8VKFIV
Yh6jDe8UqyXdWAj6M+yVqedCmHVc5KgMFxNhHtdh7cTv2C6z19kh/RhrZdlu3lJsloA6HM5NCd+4
6OUgUi/00AbZzrfYjgs3cPAaHJ7hQ5ju6LyffXTNNvYkvpx/ZngxeoKuy/Myy2kiKK6nRKt7qz2o
wTQbL5m80jMHLBMo/AegbnHJF6xg//k5i6FSWP4VXsJmiBB8Ab4whyG6rBPhVuJ2QbSDnYlhGGaP
NytAhDZifGhjevvkch+4BIkGg3N+UoruGi77QVVUDSU1uTrKU1y3SXKVEQi4Ha5T9+9aIUicQDaa
syFugTpYTwu8zY+YRSgL6JuYfTUlV2NYrGyOjfzKLSn8b5MF0sb8D3Fr9B3O8t6xfxUYD4sT9ksS
V+Rd4KLwh38EZMVY4XzSRo3Ga3LHFpgZYn+WemTn9WI6yIeAnKviAQEuGoKVOwsRfC4nVd/YwK3t
wkDFB6g60GDt4k7ZJCH1NJlrnlyyEkV5KlH5Fhi1jg1T9FmH558l+ePkOWARjWxmuHF/lKQ8Hdel
ngVruZUyjM7pA1tTlbteFE2sbmoPdM5xI8FMelNntK8akiqXJLSTlnUy1ecDLVFxvkDTceUlRwbH
ql4a5ZL14UZjR5edYTXOxsjXH8O+n7h58+UDNzF9i13NbL8MUSpsLArKPeBqMnm801PsKqXrSbiG
Qn2ABKalKc27PuC63LNRvhYkZ6wPCA/e7UtlySm/kS6k4qe53+EMS3YR7JEeubO7Uc7goACg0OGw
Ajj7/g/FgjkMpuCReoY9U5CDhFO1ejCzdCXkHPfx9rAouY6EH4eCpozPTNXurRcuChZwhgCURs8a
Vn5/IltS1OilVBSiY7dYtvTEgxkHujcHitKEAjl8/JirC0f9o+LV5AM6z920tpU2tsKiUVxZj4h+
4BA/e4vHE5BY8jgxjlOHcweTneD3vjuy2tefIuvDaYDI+REM7LVoW0EQeUI4W4Y/GyyAkGCZMzSv
nfzX39erS7/i3nasBRYPdISpL6OyHrEkDg6UFnyU7pMH2uM9MxeudDFp4son4udP9Hk0QAKfJ85h
oxcufvEGIOmjX0EdFiFau/lgAwASfOAfvvXfGDQf1eHPNqfTKG2dnL/BHBPNrFy9+HYhHVEQIIwV
IGJ99wYrJ6WNRah2+vDL0M17s4/Tfu63HCK1ehM6UUqo+3Su7HhY4CgvyGnMEm7GOv1ZoRCNQrtX
EZvcP2X+tRnrmxqECF7uNG3Ovls0U9/t4GSxbYw3W/Q4p93dqobMaShf4hasVPWUCyUOATKxICyF
PRrCcrwIgg9cP6f9Tdfh3XEBJ4NS4M7oSsSXUT7I5u1YYUwh5nhyOmKyosvxu0Ko7AuQbCbMFZZF
PYv5D6Ys8UzOY+Th0pO+jwzmsUs8zJJoqmMABk2YCrw1M4OMMjDS5HvCQR8zAJvC7YdjghLX6+4s
vhXBjflASbVzKnGsB0C+E5nrXzbnAeKJUv87W6mu+v4nGCfAKqzOxaPvjNXQweyUqFMbzpCiV9xy
aZHkBTBVOAiSEGDy2fJkMww4tSKWQK3TF/yuaW+jQaRJyXszQR3uAXM9bT3qTeUR7S3FjiWJp8pW
vaN4JvEEGyA9dLqCozFp0qxjM9DdC5qZtig1RKsPN9MSjHjSQLu1iIebWVCoNarXQwAYyXxxvBLa
t8NjWPgwycZxGWCQ724pF1QNfwidgcyYGlAakNNcG7Kqe8v0xmswzC/2qoRZjQDBnhMk2CmqFVc6
oakbbyodP4M+MzjjuLZdcl1wsHlzZipr/qrRMmaGEbKRHmWdzxiCVy2ukxZTTnRyqUSDZPDMjoYg
uqe12QYQLAK75WvlfnkkOW4qmwza9cZ/NgN7eoY3aaluKDmkML+eVKf4OuGrBMncEHYNGvm9K7jB
h+LNtNW4qjiek/aHTkJTdJcIDpIJgMmnM32TcGUx5DkJzxXOCavrpg39MU9SWqKXsHRxuIBkuOsy
pI9DORzKVoyB9QTLnrSCIaBb4ZIM2EqdCCHjtGOF9KN+XU/2KHe3qM7TsSZ+5+Yit0CBFYXRthCr
JVPiSiyoWGdQdUvMpgaplDbwJ400JvgyObFnSpsiA1mtBMLn4V6RtnVcodC1XcvccNz2Yats2Frq
Oi/uALg6K/cyeNlM6mirHqlJnEW7mN06kRcbQjc63LnSkUApCI7NWrQ2uXjFtq0Eg7/WBV8w3Tqv
fcZj0gbefQ/39gDXVV2kge+oARoSCsLmM+Z4b/rx5tNDXgiXKSRduZWVjgKdc0Wdh0WR7xZVsIFU
IApt2rVcE0TxwhMCXNrcARZpmffDHiGLeRLsI5eexffQmPWFlIYhyskCC1Y+81NAbGsv412+PxAK
Z5Z1CVOJU0K1FDDchmQeFlO7IiiJOIzymRrwfQHiyrOFW1c+QYUzlTOdmjN0lav2h/SpbYUalUeC
RhRr+o0Yu6/UnC5cKlN2qB7jfE4lxn8SJ2mOBMjevbPMtZRGl+rDZ2Mc8jyi5notQqdgUmxujwvj
6Kq4f8kJZzE0WVfr99xqVURJxQWc8MRmzNn17VLkysdnniDe5gj3y2g5sYbcZeEzx1b4gS/0aDHs
ZBbyUGG2ixVv+5yuhRImS/ADc1g9EZj+VPKK6AGCRkk0MbqQAAop0vPsQr9VRvVtjWlV/5IEYDVU
AIMVyPLU+9Vf8+9x1rnuK7t8xQikyVLtwhzMSbtIQxrnVtmDz0jar8AOqRXZS/ikAYAk9b6JbqGu
BdvpgXm2xzGsGQZ0hLaTs2xhvSgNncgkNeQXlSqedsCqsR62t7K5U2fBqQaWzcVacAfhauqH5idU
25wNsQf8DcFU5XzFnrFolVwZQcLfotTYxAREm3JHKWAHkxajM3qvwii9zOlDydjUOZ2vaxoUbhr9
Ao5P14npLuwNcjme7tygCOIZt46hmUIdiSHUM8AhFLl4G6grJSE3glSV2nvLMKoIGKcpCQy34y5g
S8nAZ43YiAQ7DtUx/RmAof98gy2RxDHrXAsfQiXVtXxMBe1jDmv3CyVxBpCVkD3EJk+BbTYUAPhB
SwpaUgEcCCXvFceYXJRTan0PqewGefrRfGCSQGyYroOVQofeJ9FZoEH4TZYW4uXAzBJbzVGuMmZW
eQsJoQg5I7wgPByWWDFAsY2e2+e9aqtLHhyztMrc6TwOYgkZX6x/BgG4kVn0LvwrV6n2Wiw2XvjD
TN+JXU4y8PewF2GtJ4pIORpMO5H1MSoWKY9MdZT0OzYa57F4FcTFunkcJhgmwo/XT037fDEY7yaF
8iPS7wi4+/jlRO2mbZh9H3uXb1O92743WcPoXmQX//y9YUnCUme5f6zEldmaqq5e1dZKJj352EtR
QCe6Pg2p/RR5GoGPgFO/ECBpBH7YELYJsCJKan6ga5gyDtQLDEj0SeFNRrUYzhKGzchWLDoOuAyh
6Omvvypxp6tWBI/nuJ7TXYZJSE8ysMvoEvRwiD9Pu/QLNchWy8XVpQ6+NrtNgpz50IcU7FAEyvF4
C+hKJRr50AL9PTv2ROkxP2ab1x4mDtvFf5N4u+ZQkY7zdcAtqJx39thAFxUSAoKs22KmFB7LlMpO
d5vNlXUgDcMqaz+9r83SFGiNXbU3cdg8dZsUYS4kXy3l9ZIaYqlogG0ED1CTCVrx8yJrNvF1bmsp
dLKagHGNF1ZCSh7h+IZZhc7toUVTYgRr2U021+qdKN8pi81NGSM72NbAypZtICEswu9tYSfrVYYF
qzc8F4uaYAf7htPpZLKodOocU3On4IstrJTCOiy4NaChGVIJMGSGS6RntWLepx0SXw+sS2Fkpw5S
8eK38RzFLqCW1LhliR3Vzh81uczisAUNZidgECrsVCrhhlsbAr1ZQOaPQ+zJj9IGG4UDwUpPp+xz
F9werUoCz6QEUyT7rxCvT1Z1nm0ZNgx8bNeFGVIr1Tg9kc+YXf41/A6dyqYVcHzhIDo3wnRsDBzK
8BImdBOoaRxbuLLuwHiUmhuQT6AWOh+X4kzhyPd6E47CZsDPZDaYe9PkeI41JrBreNSdKfn+qAWg
3yItCkt89Pq2BoKzByF4XmVWGKzS/xx0jhv3heX2cmPoo0pnZIw+bRZ53HxuNMch5LGHU71u1uFs
FcUM/QXKJ0hyY2DKeDxnHFi9tRpMe1sfJ3guT2y3sXhfAv7/QenqMjn2o//kccXiZITRRkndeo2E
XJBOlUbk8gL2XHdlnNQcrme4qL+M14oirab6rlOzx2y+h/92i0M05e5QHQbo9TfExVh+WgdfcWLu
vgoCLNt+DLPtGLuXtAtJ/HN4oLK3xRsOlMvfCHrIYSpm6xXb7HySrKxNPK8zjpfjTbcOM9iFjciX
BMSQ4gCGooir9U4UJ5DRcinL3NCARBUjWeTWttdR5KpdnkFmniUWoaE3eRBcEmahglipvlxe43DH
sJqVok4JmSnAGfXIr0eWAEHHRuiY/sf9Q/65wNTmOp16n97KysiWoUoJrw2HqxXHltGkQxD/ujgn
86hWecLCExCYZaUMPNDMw7sItJbckteuhlSWqYYqoj/6+BCRcvJ29T/bjXAcv3Lyma7cDGCNhAnt
VkhGLoCp5jXpKP4+uMKqhnl5pq3/sy04D+MlL4Uszu+WnGQRqWMYGDwrbbmLgspEK17NA9nkzHcf
oRbBTcPk24nqUt5ySkz/v8PP31weowTw4dMIdBG1dtseltcMZ4HNA9LZZnhQgoikGacCT6NG174g
iibuAWDm43/F3jPUVNhbKp+Z57Icc1cdkq2ikk1T0xir69VMN0iB9WZ8UjJ0XMXNQ5RAV0l3M0gW
rEzbwXx/la0YuJ6/a3w7YndHq8BkF3fMV7XMPWPVvQny8rXY0WP6IopW7WM/rdAAXCHNoKcdlnOB
cKztmtfCJ75i7Sj0coyFg3pWeQW12NkIyT2Kmt9aibQOLN92CCWrJRQc+Qs4YMRXNvPyUye2Ntby
an8gCQGK4qB3DQwaE+In7DNsoBCLmRo9BBBHFDCZ5jojg/2CXvUIRPuW9gvqji5ihckK4hvgHSiR
UcNuO1Yn/xyrmKk2dI3YUPQfM+lI5zOzNJlEK7wPZjLf8kydGo7XmRUp7goFM6mNgGYobY/4WWHN
1TTtWB/2TfCxjTHlLjkL2miPCd8teJ9qnjICAKyRwmPOjO0Hs9upOZlILO6h+/6sGAijMMjkeImG
YxEbSeJqDf4wQ94J9xLG8wQY74tojWa9HQIqTW5F7GmpAACsiOUjRmYuI0v5wmKYuPF7p5QdKuMh
aGQ2LsHT4Z3SJacBQl2VPfdBPS86e2JVXCLxN6hZ+Lr0D6NGHtJLTYjJkScpU8r6UGXPK3Rbz5o6
PUVAfPPMYHgN1OxsRMlM4y7CQH9ScM+GPLSVLAmrMds299hqdGJHZL9+FYMfeAkhrp5ebzAeGUwH
FtNbXzH70TKvM4jCewxiih19Mg+dzIG39x5P+95YmNQv2E3XW8y0YdXUoJpFh2nGiM41nZYm7NMM
BTMvi5d4xqVPgF2CUcMAKg26Wx27qgZn58RN/XFl0RtwaCDE2c58EFwj1YBrgEF1+GzIJGqEdLT7
/NeVJSyvr4JvZH8C6OLDhfFa4llUdwogoKZDo22YGQa3aZkU6S9tLUfZgMryuMhEl0MCqEMUL59r
xdfofRLqXyKe3GG+hTTAattWVRCmn8XiMJRCbtEdwCymWHOqQNYxX5asDAMKPTR023Sr0Q7KA2X6
QIhXMDruf4UiB7BC4F1pGvp2lOfbNkA+lDoqr8MwFvxVAxiY2us1ZCfHLekdIgEbjf5123JYizRA
UE2S00p8Gk2Nz67H0OPwFL4DwRrQt2XG2g8W9vFovySuwokbadSjDL/o75vWUvRAjVHMqimkNm56
ejPc3rAWA4L9M4bfDvt9xreCzloGBf60gBrMl9Gnv0NpAUz+37TyIkf4MkXzajXn08CunY1gaz00
ceVA2VBpC/u3xI6YPOWZ/jCrcCwl62SRn7OpvOoIREyt+71qIbZOVd3TKaPW1PMqedajr1oLjGcN
QHrHR4FTL8cscHgonTeuFnumeLvAzHUq3O7+ZEQokYR7SLQFAXESEvRKP4szNd1EqJ6zLOSx/Dzu
MPtiEzaNzJqRkT0FYVQKzRU+zFumim1ngG36sIzq71jdxmcoO22khJ/cDTcOvtujgJOv/DJI6DPX
vBNzHG/rGoBJbGmyjOQQNn/ht3x2YRrqAdhhjJpCJJ+QeEBrHDB20prQsAUj3DSQrQmFNkQ6USZs
TsPDLotUxzWtO92gN12wkOIJGbfa4skMxuVuJX/MgZtiJBayOeCAP/UvUn+dewTGJHcM5CvYrfCe
lw8sHYkCOPrrce4ERRJJv305ctOrSTQoXg9sPwbIa/u4Iv6VuAeMu6fx1uRzD4A6JCGSua101O0T
Aq++Nt553JHPwx9hUPhsGEb5Q+yphnvqqpDoRb9qEkoPanWZrOMUM6GBIUBwxgEntAJB/QY3fZb2
2714pjn1kq/GnwbWctCG4czhx3b9VZtvFyfkK60gZGOZLHusupETVNlR1B9IMdDhkBjY/lX5gRmm
xECIm3L9bAcP1osG5ec2siAMA0vfkhIKMVEM3ZeWTMCS+Biv9kfgt+1/H2L7c9aGP4HVmM9vPqgf
kX9HFUf5G7Le47cXlBjix8HSdtHTxMCfC/k6NanmYQcOJKeMu5FpwnoFv/AQpwYiZcVhRHorW8r9
FC4MTEmcGDlHQlo65I08T55S7UYseO57ys2XZpo6XdE2lMDUNfMKLm+POfYWSonAmTa0LJ8JajTm
zX9OVZVVzy80ZKHir42RZ+LZbTBDx9+8EmrRqnRqn2YC8snrDVepL+S3TDlbczxRZcQky6Kc9D/P
cI6MNhe1OI7ADNyLlRcnKcqgLm0d6NT4CUkHJsuUHAIOfnNyTzOuKpI3K5P+JxuaXMrVhaHXI02E
iiXqzzM4BQpAc9/c/2gRsfhdeL57h0vU5ijvdWfm5uHsnVkXOkmR/0Fb6h1by7eR/YqqfnCeaEBw
fdLdRSBscpaD6Q64SnkCb/bqooPWxN0cxdStq7/6TM90SwI6GXXzIRWyLSW5ay6we2WGJDomjby8
kVZpy0UdMQxdBwsPPJy74hR+HffvNDLNBpK+FdePvsQHqM61UjDA5mAAzruNHLX9xYqkeMQiUju4
3wiy/85f6znXZv6xw+tB/skkg4FXy4rg5305xiJ+vdojKyxlw9vGKDxn++6En0l8OHeDeh9ox7y9
Zr2msL93+4jmoniMy3NEnbFcHUakV+Be0eciwradf2K8009IX3o4jFGQRM4P2qmOvue1Ay2C9Uyv
nRem3Fz86h7YdgZZEjqdUrwrgjjdERYvpTwbk5rhsVQ8M2FMAZRKP9mrr0WHhXaY4i0jbpcgiwxS
b1GElOWXefzAeRELJTIT+6zRDc3YFlcjJtBYRqa0UCisnl9woMchMA9Sh8tvoyLkdATdXq6MXtd2
p80/i6RD8AaaCyJwnIP65P7lryynhG9vQ91OLxaeRBsdUrjdXwUcw66BK5b1phDohg5kskFX/MI9
nSR8HEOthT21FQQIbrGpjK8ar2TbmbcxgRUjZeCPZsD0DpJSvkYNl/fsveVp9x1NKYrPMe36g+78
bgI8MbDOIPrvb/Y7U7K6sqYh2Kj2jmKS6t1NAgRmjOI3mU3CXC4V24Kg/C2GOKy511PiKUHXexwf
m6FluEDyFfbqUh9eMbGOfgJNeoejjdDwT4fGWZYHwFDLOSn+GcdfYCbuue0Wh5uNUqhKCnJw01o8
9aO1GSqpd9CTNzpRoDcTEZ780TimaLjZfHORIicHbaB8Yn9z5F5ZULtOfWOIuMw68VCs8QjIU1O5
tPNqylw4NttsyGw7QKWkIrDzJqrH5V//euJS+KZOrVLejk73Lquhf+KQ9pBWaleyqUPBAG6Q5bNJ
/kriJpW3Fq79jmSkosafkPJIbozhyCtt0PS+E3w5RzL91epGEt72TzTwg/pDGcam7uh5RAMYa/W9
HV4YaCqcHkFAWFwMPqrjyyqEtNxEcH0iiL+qe5y2zbYvvFxel+Bive9Db9gNSWNPHbyyd3HISo17
2bJYdHi/XwUb/pSbsCuJf/sPhlFJe8IskG/WWF5A3W8rsBj3fJFbPnIDe3+4oNOUuw3n9CAO60lc
0Gtr+tEoi882ILUODyDr0Q+x4QJqsylBFnuZ/Q273fTD3mTwoeqfA0ImVzOafTeRx72Pq00XSfqP
db0V8hXWZr/fvzQT3FrDgSqFNPkDOrWX5oN33tX4BpHnuNaOL2WVkxXYUIQVIfzVYIlBpNvc2cfO
9HNDcRxgfbJI54aZTFP2Vs6MTIhBfjRvf6R5EGnCU6ScFHsbCmMaZuJmVYok34eit6wPWFAYpNGW
X/169+xxQBJTEjZP7epLsULEXrSAxTUGJ5HYiVdqjdLDpW65WOw/VnaN3jx3fKqMZckydDdD2RBH
PH67UXmjJcMytV8dbVkQ1Nn8NS0aT9WHHLoWAfHWBIdUp+uWSnemubJyaWaDBH2yL/mLxS3BOryQ
YRwWEyZy7s2fz4Eb6PdCpe2ZQkxC0RIUBfLWTU5yzlnvdbovEhzB8O8uxH4u1heYUYwVKkqBujog
cEsqnBJRd8dvAi9JtsCZ1SKQefCFRFoTM5oHOaS518EEcz7rxrJsJqUCmZvTy1yP9y90SwCNPmqS
MAIusc2jt77J2+1HQTbm1aoaoZWtrDeqc4UPOT2KtrOQea64yh8pip6KurU7Z2uQWH8sX7wfoD5R
Q4au0RW4vx2uGlDHnBBSpjIr8uNNdzQrnZ74Y3v6/i4bQWiQ2wwP0TppyoM0d3uj2k/XvoBQZwUa
TbtajQo6IuX2iqdi0OwxeiPE13zAFygMrO5TwUDinQtdtC2gQy8jwjpzS6291GFXLO40wuyJPX/B
p8kl06CXLNvho8qNwDLtXuDQ4EAd0lSUjkSzDMZm3yoPzd2NNeRdY1cXOW+Y5m6t3NFnEPQbmRzk
SJWvJTZ7Qax8ut3ekGgmukWXXT8DAPAKVVtmmf3wkceQVcJIWAEw73vz5srl5lVfeUgNGDJ+UutU
M10NqjLko8Co33A5yvWl+sXNvXt8HJe//qHdjHRjgTe4sTHd0T/y2Pvr3EDyIoYWkObwH+iDzadw
bIryfTr4WJsGVSJHcWzkMayjJ+WwlO+Pe9qwJ8BFCZjmty3qRmpyNilXc++GlYab+8dnosJ/84mh
CPOpDS/zn85BzvvzGQ3rNznRq+IvxWfhIBn2l++GitFWNFVohj5G96xTnyExUzQXu6VvE9OXUi/u
/ppmicz5Uw1vZPsCTjfbXYomEvqRyHkLhjfLDgjGAc5EQ/i/dUp3R9mxHJq4t46OrR8XobEd56IG
RiGWGcuGeKaXf7sh1onlwKHALQrm/zXObDlwnYnoHuqLe6+js8a7sEkCp8EczPjyQ1zWugUSGU6s
RJAvA+UxoL+5fTmOQrwfUgMdSbjS9PNvjAXpUhHnk+MoydeFD4FP2Ebbdf9p+qS2qtBpMWmjeXp3
SEHt9bSjbbcfA6ADe7JohlbxxxD7t/Cc45OVaCMCaOgbNRyuY7lAf/dhNI4pe66qTSfLGEbTS2Up
9ZaudrmAs9KFtf0R3jdNs8FLIkRwawCn9BxR7fLh5V1IBssy2HWHCnayqmsFL59hEJ8QUbWdhjHH
mOJSDS//zx6WWVGuzWCcl9hXL91k55FpQp1D0DxVBk5Gf8YRJC8pOWOL3QH1+BHaG1O+eokrVS4c
dV9GhtrBZtHMKKSv/ueJKl4Qf5s8t1DgT053nUJJKIJ3AMBpkGIqQR+sq9YCH2DV/YRm8bWOGoLM
M25XhMzSd9gV0nltNeGCs3jybMej0spo59pkkiq54Wj/UYADGtPJue4M1bLhpDmwY89CDqNJAPBz
419Ry8ghoqO9jfKElIElpdAPwoRnai93x75gQwlzP7Ri1rbtLNau0A+nRS3J9eEMxH0dA0bSN8H8
ocABhqAxVSu+NZitSuGYtfOFakSyHHdYrVdfQb5UcYrsQ/8ziJPacXr9ch2aGTBPgGkWl42gurco
MKOFREDiIid19V8aw54ccKBw/CXRmH4nsvF+XD1US9ZJBfs7U92Kgj2pUDyjav9HuzESBXnSvK0s
u/3DbsQGFEroqVjXevwq5k5lcJlJEPzvt0W240YvNwda8shkZrKbQ57ilMAOpWgXKceGYbuvnN4L
KlEzPsfIr3sGUkV1JIfPgMgv/H9CEnw792VKw4zdzY+eqCW0TssDXW+0kFalE+BW0CZ0tuWl0fh7
TN3a/YV6WoRHZBpU8HpYeAL2mUdSg8hHFczIRr8rtojoto1LrH73ctM1iDgt4cWIg3xRSO4/aCLU
Fx97sx2xTU4CwqDzKMqCcTYg1M1AeaIFWOSqlafmrOr/jc4/YtnzWaqeg4c55ZM6VlAyD9ylS+hO
RlTerep+ERXsWkQxDoRHXoyxDBm7fUI0zQJR8weAe+oAaZdq7bgWwTMW0MRFxsCqTubdg5HQ9FgX
jpbLGQsHyQ2zxKWp+Wo8ijMupDJDRDrEAWnCtEdc3uysBC4fBftcj+Lnb4PpMigqjX6XUL/6t/Oz
8l6rPWR3bZkvVLPiYbqrT0L0b3nCRxEk+y65HW/s2XICHHUyZiqSxfI6DHUGsUMG4HC92FB4C5L/
s5bufUneYAJcVEZY4bl7mj+B2nSYOKfNjgq8f4pNrgYwMbstbGFYqIrfBBLf0nYeM9OBaibzqCQZ
5Nvdv/KHAYMGNQ0oaseBNGhh06wwoduPqnqmZWoKDtrhyUR9Ubb4KtJVZTdvLFunxdH9I4gepUw8
YNi8JZHQYCTyFiKdfo4LebtETanNpTQvS5THsBQbATPLjl4gdptl3wE0JYo7hc0YxUQES4vRigFG
QW00t4NdqD7Fe3FhDNQRXWiWdti9pb0Gvd7CiYBWoQygZw02H7EK/DxAngMaNUxNcdpoPTRnw3lG
n4LnudYr5cR8WRTgHkBmRv/F7OOl8ADBz5rGqCgW3wkyoazSfCo03yrhUyjpl6v25B4AVgMqdasa
GDCx+GUfpXdz0UdKAr7YXMzsHijaoHksmMzR639HMFtZ+mlQft6HLtu90WwutvvDTHyJ4oawxFHH
5hjy+Gl5xDnEeWwK+qa10iYXrqCLQM2HNkuunZZeUX6mtQWdfJBVkfiCQKj+Q2A/BCY777s5dNqX
joXov2AXy487tcfTZhpmhUUeZQL/AB0BoHJE6pw+4fYKsiE9iEH2odm0ly0kZsYl12aRiexBmz+g
5U6pDoBNzSz8jzynbR/nA7OLNVJFwa6cNx9IrsfZ33n/ph6Rz/82ijByoxTbTQpM8KndM0aRmAx7
2FOZlj1/biQZXjDblooxfxFRXUgqhK41d+1HNhc29VudWftSUbZSshMGwppzkeuIXnWeIDtxSa0k
9/Aw9etjLVrAznJW9fuVpsLoJIYAZxlGwEEVItbFxiGOejgz5P7P5QP5gUdYM+6Vc0IsmGRCGp1O
3LilrDmnS3k95FsFTjFn+r+v7twsGECNPyMc6EQqQ2pasaMiay1G40OnbTMJ++ewmDwv3z+37Wsl
O1sJ5P7PiRQW6QxRYNSJhf22ncYoFgcF+aHrK7nnDapWCycV9XqAMNIk64iUz1vh3BFfqOrWtjUQ
hjqcQUWIFWMoxUL5r9S86Nsqt2AQ/xTydDvRVzHuahaVqLZTRzN725ovUlZjRCB52F2uCVgPV2fK
ZNRjyvaVLH9mJ566YLbkY6A8mHsCS2uY4CMfMycBgVa9uxQbG6TdznsiZBU5cgJPRfGxck8FjtCr
0tv8+72Up7qNhJjSyvX8jw3flYbuXdDRpylWQ5qxcoF8veDoIse1FUCgS+sB3RGX9W9aVB1uo4IZ
AkQCr1MEqtTTn1fo9LBj6zUpl/iMz2sA6xm5aX+DA9EaxlyyVlV5DF0Lq77MwSAjOAGf2S+FjPqm
1RDfuibLJorpeRoZZmoBlW9n7n3Q5fxu2eGWZtadnO/7Ajd9Vdre5sd0D93EQrgxPC1RpxpLZOpY
D/8dxt3WB2xqUcXjz+svC32wI2O9er/W89BLpDlpr7pVsEWPu+i9Yn/xz3apjQz9+5exVFecrLsM
DZRZl0dNucvFJQUUdAio54pL+cMzwohKmhsbaTuITF/WAnQMgzL4cx9Ro540sahOdJ10klQRuj4a
AWFpudnWErWLuM2VbYwtuHVMFrxF2nmOyXeZBieCEG7nMXzffZDal4DqbhtDhuyICkE8eZmZQR+g
j1Xgzvz8pD8GRhE5Aylz26b+MCfDOVDP4JUxk0C+Vn1rZNSQsxHeR1Ml+jS0rXidbBa0s1bkaJiJ
rME2SxVjcSH8+P9FB2BqICAVgpGLmU2cJvsKUMPrqeacKHZUDyGMWv4LPNotNLCfmRH6c7dUawQ4
MHd1jnVUTU9ZSSR+NlIWIa+9+LVg0s1HWY7v1kT4DkHDSzmezxbqeaREUwiFRUFVAJD//vqJIoqM
s4Duzs1AwdRs2bpfC4mlx4WIVIrqAc908BQNOeUNyXzI5126nBEFUk1WS2vXnYzpMtdsxQQ80yOC
wvTsNN1HkeeHMw4inohkDWtVyUbCYpM8Km/LKhvzd40jGqFEjMHPsayVW5qvn+oIJQWWSz7h3zUJ
hLxaFiuC1zKA0u/ZFYyNJCA5k/HWKKZ0to3yGkbIAIZ5VAX3AlyIZe0mA9CQf1vwPCpq5HfE1xGC
rJdELil3pjX7iXB+gWjqqLNcdXidh9FTssOIhn7CUWQZl9uNqD2Eaa7KcVykXo2rtN3k46M9VdFx
iL7/JQdsULj71QrhZ9xeaziUn0SOv/0ZBcPnlq6i/UcsbZ/eX/5Zv3tCYLgwQPyyIqIQOwCWUk2y
8KNz0TctgZd2poMATZP0bo3OC8fMIVbtMYzU0ipvsHGRzLRufu9nOyVKCm2hxMPhTJ2SM5EWqWyW
cTNHdkGKALYzf2Tz/lu4o+NiErakZOIW+9DoeFUR/JoKyug1HL+yS8Eph7QwlTqXWO5LrJYydWw3
wb1JZLGRJCuAkA02tth072Qrys+UqqDQMSvMqd72jDbRFMk6h+h2PsOI26X/W8f02cC2HyDJ9joR
zbLM9UU9oxAA6/O4a8kL17wgc5y6swlUNeTGe9LQN4K+XSO3pibeqTWvSLBDUoBiYrr9ljz9CygY
Jeaxxs5fc5D7HaUdd+xvMK91xvPKv4DnIfUajEObNn910qrNw0W17XPWngAp75D3DXwlJU/Nt2J7
q049NL+YQrcGsM/tluYYzq13ybRuILEHJENGR/XMTaCU0I0bZqXRxi8RRFUXMsw7aDQ/AckviCE5
eNWqzih2Kwqm+m7ghshYnGU2BOMAN2L3NV2Rtm8+lKs5NTS2oLU2Z2qAWLueWc+HiryiYAlhINat
TVxtEL/PQmP96yIsFJLgbWdV738HaxtVR23lgc36Yf75/uUJjRqyWa1x03F0KKgSDwjazmG+FGxa
80KTOkkM9odxCTK5a2Jpg5GJ8P4/gu4e3+6FE079TATTmssGs++pBqkas6QkkHEEKiKKbQEzE6To
2Ur8hZihAIQOeLEEDuIXkC3y4k07+EqZCVG5jqgSD7VC3ICa+0TJD0mA9DdYPOvfnZkugG8fN+5T
C80FXnmGyFSYVy5E1TaI3bMyGC3ZXWkN60w34bYBab3P+cBi1I6clF+Vh769ek7EXa3RA65IU+8q
Tb1ZYHYTbQZMeIqgyqJms1g+xjMAXK7o8h5bryUR3dIdORw7fajuegVQSLZf9NpEJMPU1+1b7gcr
G+gB3y6LZ0AMhW+Ej2d+G5ClPsXTqXTTShI3zsSqZ2TzIOWsrFjeTnFUNiea2GqH64LtnB6sq9mT
OJenA+NCOIU0jfxtzygG/Pu35rIzyo7MHOcs320jXoKf3KIjL7D6BkCD9aZJWeIjuU8rHWhed7NZ
6jDekIu5CLrge812zaCmPMQ/t399aaFDJvFJDI95WFXsSxKCTobFzyK9qto+6JdXTlME16KBrde6
albPfCfS3wKN30HFtC11mxQ6HO+UHMSYsrvNkGXzVikXLkph+lrM7OHQ1/6vyRbb+BIXqqbBjR/F
1HLxOYKpdoVind/wDg1z+ODTtRpdQHduixHtGjLyQg2dZM7jrunBSnU/PwJLX7c2+fmYbHeOA2nE
6XzAB5StXL9ydgmaNbOfO0bBsql7SnE6mOcFn1rmvL4K98mRJmmsVUFdZjR63VUIM/t31Joo9uJ4
BT0l1xw8DdBlyDK1qcbEhzSFjqYMlLIoHu2uJVHO+VvvbuYrFw1uSKlEGkuGu3F8tVNas/qm3aaZ
F6vj13Bj8uEhGo41jP2V+xMH7CF0e56fpxHpNnGpBMuXMLvlhBXaZuXKqHIULyHN+PcEdG+eAuoI
s5gLIPhC6hjFb7/KUTnAApA/Th978O4aesojZQdKFcCzxcAt3cvMva2dXWln5KTu9jWKYxxS3rjl
bMh/6/luXpgBK69EqgMalXty8NSXLTVzzr+JOcxzFtTWMV6ouLHoSv9McMfCRxjXTtKLd4qvcyc0
J4046SoPOP04EStBYRIfIpEPDPVnqx+0oj696+5L6GsA+J1/0HRAduedDzdZ2PuDIwmJgKkMNQMW
nWtJCKgQNqfYwjonbiXfb1eRGHujigTZha0zQt24AvrU4mlU54WIYMNhV568Tucg+dRwu/KzRisd
z9BucHWln9fPYxoJ6Lj4zGd8BTw/YuFn1C3fkGZ/z8dZw52SRTzeqKoy87sqimESj7LamPGie5PS
2AYeDXxmmfI9jviYIW/9HJo592YqzpCT0mVrOEPStYctVBGeAxwCF2Cj/yZ+qAi6jTME7CNzznGt
lrmJ3Vl9WAH1uQq49AiID4cCwjCz0TqhCORsse5ZJVrn9W/FRAuxOVe+m2jrAmoZVL3ZlrJI9ZQb
axk7eTsGksRpAYJPkl/Mj5aXu71uelL0EBE9ZER5MAZq1X+8MBZw49jpdjNvlYfCN52diHRMdQfC
CBi7ORzxg+oka2ikQUIMhr8QzJMYOGtMiqnV0H3WUlMcJtHD54wPZOfkYikIiry7Ju6OMhexgPH6
HMU2HoXQN7Y7F8FoZbsYA9rYUgq1xCIVvReXLOJ8mZDSvKHeY2uOYti0KJuXhdJxOYoSVw+H2H4y
H1d1S5lwlgUam48pNHc4gqQLkttTxx0lHSaPFerwiJkBjEpXw+kzyU0+9jY35wWj11hHf/3bKsdj
W2h5CI3g2Umv429nznx+hdNJf3jlzFsrYQ4OauNy92aiOJldU/b0SQOsq2bfa0F+OqM1V+p3IpOX
3AzEU/v7HJOP/8BbfSYbbQmh90Y3jvqatn5fMObP7S8sG7PsS1DlvIZ5LWzndcGk7ov24A7wwopZ
MDY/+//fs/ViCq7eCWc7kSnsiN4zEmkigdF1FFBd91qS/SeZGxOKfb1aK8W5IRw9V4OnF9WkTjMl
czFuOx++AlWv5zjj0Dcnhzll7NASePwPnV65a7UAGrhaUXTHXsDLVJ1NG11Soh7mGN6P369rvwxI
k/A5TlmHcpibKBXxcOvUK5pYKPgcJGtcWG8ol9S/kMVrRZZpc4XH1COfv1cs4eg/TaZzcuaLOSV/
qz+uK+4kLORyb/Nj6NpsFhoTD2fxFTSW/Y+ro6xpEDLPXV3YEIlWfAwdWiNir5nPk9sG6CDbvNp/
10R4v0HgVKRCFz/YbkNMoUtZaflImKdokrnwmJuVD8ysNIAEiA8Bc7n68R8aBbLfrz3GRxRFzkOJ
r1niEHSjOIN17x/x4S85PtLnyIlNyBuWUkyO8IDBUkyXn1jwHVvIRjdlkPRAZm7K1otNxIELYvVf
GzaqvG8pT9WFUgt42UuGa3eTnDylhkzWpcC6kbzTxckwOU+zTZEihysk81Zhbz5brDDRYvlMSNlD
8sAw9mJxz/rih5dtFIvnfvZcj6wr6jTuFXT+wIxtZ9IZ1eU8vulvY/h/n5vXilSldJ0WbJk1Glh7
VAmHF3/YGILO2Al2GDZxK0KivNbvVxlrDF1L46QTlHWqGK0gA9k5atl8UYa9KjdARQVFHshM33Vr
iCaX15caPS9oUkf1D0dOx+92elZGOf1P2Bfu7xBR9bOJUQSruGCLRAUkVBDiiKLjgGemZXNSckEO
k3qyqsw5Qj+OcLGsnd6zNrmUdKhgoqqw+moyEcoWn/6BQHMvTL9grDqVar/CioHIm7suAa0X9Xkm
XrTBFhygaK0Y6D5FW7lP6WUDSShqCSKb6BwtteuFT+hqD2TDuPs5Npq/DEHKi01xKD/DyH0XofVa
DYfv1e3TVJnC36rmi1u657vOH3DZ+zUzDB6UtrNyAN+TYMTEJJtbZVB7sJ5Rpy+jheo5ujOYN1gm
w1Ppwd66IBNT9pGjyxSMWKcH2Ze25Omi9tEKi7g5DaZh0BHEm7yj9OY2sBFbx57LZFdBNLQ4gbms
8Cbx5gQowo9e+26aoue9RI7Gy5gZeC6Q+ubgPqtsJIovMssRitxhAsJyd25sxfNkvXTMxKyGU8sv
vfFBVWhP9yk0QPEWoK7maSWvqx470Nl4KKs6MYTC9+g/J8iB62fJV/dnSlQ004WNmOsWkztIhqN5
ptk0cRo4gq7WKJnkRP2cr+bK+Ih8t/IgqLLwOU5DO74+cXu/7hvLRcnxbglIkM6KTInIigY4cQna
pHnQ8IvLxEVpe7Bytax9J7/Twp+WlGfzVueJv/Oa3mG+PK5j3vRBa+37KqhOPhejt1meKOgXClxS
OQLWUyj2Sgm8YiDmPgaC/zCxQrrzAdTU7kh/ZpaIFSBTaohvy7Fo1gElwk5n2FY10Lp3fgYwPwjl
akT9w1j14aaMFB915TdXPmXZgLUChlah+opOuoCToWm+Cv7Vcn8pxWpm5EHWBuRgrxnMLw8OTZJj
z1bzrBMDl1X6gyQ11nFgMkKftACZk+oS9yhKJ3oqgMkY7LSLhkiWJF+5BEzgNCrb6BXLFknMUMNr
6+AASoyV6t7qe+BHguSmrToTQk9emD7sI7Sv13XyQVUAAGWPWLiL6SLnie4UU3TJr2mcZr6Gstuq
MhpQ0twwPEaUszYp1tHmqMcAwi0V5mO38LaV9FKGob7VasNlJldNTzgpXhLutnYZo30OV4MnNE+i
CzGNKpPZ1oUE582eVY9OAyPMWuQj/Et+iZz+ZoMVxXubamFknBwMP4NbyuJlopO0qCOGBQEp16RX
GiW28UC4K7WGKSHy8cAStpBUmri754lcaw5VRDbcm/+uFf+LjwKNLUrf25wNlkXvq4V1rxGFkQUh
7P0t2f8Bgp5qrvaOrImqEhAjvfUXpRwS3iDat4YUo9h52wKtCTnmDOhkwBK1NKqr6cyZqDC7nea8
y31hgmsUFEQJ2bWw2B72BM/Al88DWfrujL3pqIcp3HkjtGnWZoQtdcB1iajl8FcEP0V0VyWBFoAb
nHxmEX0JyLT9QlDy7sICiVdz49PDnBTZGvQi6IANxvDV5KpNiRQ5JEEqbf1dL6NaOD6wGMuKYQta
OaNB9aywCwi+sBjh09IOiSQMAEV7Ew1sCtsyoNVhpriWn5KXGG1vGDkeBxw27Ybp2QWZszzvQp58
vKjQWlAcZYeTU4EvsI7VQfshp+Xj4vc3CHvWgXZpBtHfjcwh9Z8ev9EyOT2S1p7JdkU5HdLHb093
TchGMNsPBs1CQz9RFtUezcQ0G1ZIcDnWLHrd5ywTbS9Q6ZfHcf8lB5Lvlx8ZSDILFHOECCW2Osa2
5stZtSS52pel94myqEYI5y+sWUqWnS9vWS1nodypX6kSXaUIEu2rfOizbqPcMujPVG67l9EQNDhU
H0raT4KXqvBnRU8lmJjkwXrcrqM2UkRCbul2KCIjMUgD+2tp5AXjHVuVoGOiTm4JkGwvz7LNEcVf
rfr5BAoCRLB8GD1CMbgx1vwrqih3D1vXoeVg9eQ2qKJew/8uYAZ6kwVpW8BQ1eysyg9ryzw2k5+r
ZJ+v6iADKkpV6V+mvtGE1nduVGkHivgygfGtmd+S3qrcnsbL2mNJq56j1YoSN1toX1Gg1rI33t/h
N3dFOxnkmbFDo2pHecjAn6caO8Nxvij7cN1Q0POzdaAdtUFJhtIzn7GrHw+kK7aMUyGAgVMRjJgZ
bZiulOxkeJyOww9co/DWDkoaQ1s3L3BMnWzzGzZsjzjTo+ztn7iazOz69alzvtCX8+HIHniMQ6PL
FVB/LSKSEQeZnJ5NSuz6UpIL4nVp6D+Tv/VyhTyqP2x7w48S3Ya4AB71q6EaPEjCqRCHf3qDiKng
d87/RHK2mtDhS8269hZHePSEVW5Aw1moJ0QemsgJQjhU7+QUMpExYUAbOV0Fkl7cq1e/E3d3+dX7
/rQ94YHVMbdVYL/cZptY/7rmk0dpCC5lFS/ARJXYcGsFDdOI4NYfrgQXr87mH4y4kkjewZaZ+4DK
BaRaEp4TAgXWQVc37+48IC0NmPgK8Fi2XXaRUYzTiDyP13WuCBMeDap5zNMgWIX/FniyuaDWU896
DOCcf7bK7CVp4ZtMWJei/UuXmwHz3bMnL2a/OE2/UjNX9ogHPkVmVQysnomrZAP/7AEWa+C85jjJ
bugsNV0GYZOvr0iWa0fMQxcNLcwu+3OyjVwlTMuKGi3vvWwYunCigtj2kMSn9GIxo5JvESqA7m37
ESTM0yK4+zioAPgqIWqumsT1mp5RGiCQObk+iJnrLqPm2HA0BiDm5XofJV0xIGTA7jUbtay7L7ly
wBfkVWFIbO9wSq37HYpjUnO3MARVA16e4/Fix8XEQ8sG7YuS2a0+6GGwkYh6STwthNiiyMPc2dYX
8HR0enZIk+MESvM1qh3xgSE7ACFwPqsezai32AiWRebsXtKfOXAMPryvCwOrTDh8WFnuuPUk+S7D
D9TqkKncUPOeXdt9VwM2PUP7Vwj+YgdlgOT4+AURByENIfz8pkWTyCA4TTCpfGgNKdV0s52bFMKr
yPt1peJDyqbWnN+/38NJq0yIBYvQiqcsTfHyqQsBNKvyZstkNoSBv95moOa53Cv47XjTEyINkuWO
Ijq6oyIgYWmxNVVw0XxmJuO1HgGimJstTHlqbaZDHg/t0Qz2AvodJIbhkXnYYRsXzZX4z2tFuJdp
uE2KGK8uxpCdQaUIVGHSxLhukrIJG6BCWrtZt7LgH4qgYANnfHwCkfys+FuvcyGsxEPmnS2Zr7Yx
NXpoka3hhCK6h+NGCZU66wecYCp/ZXE7xlzN6scpuxHKIcawnzMgei22TxJmMuiQMYvl1tw985EP
kG1wMvPr2SyhnSqvlWGg6sNv/gD7a/Qhh85PXRlf8JmzBVXf2eg7ipcuCsqvpBjtnqMVpIjGgTnF
KAX0cOPKy0QvLSPtt9GBJDhGqM6lhU7FsxS+10t7xehRs9Qvng0t3xfs/nP/Uh43BrpbJM416jja
yRyUDdkG2/nz+FbA8d7DpwQs2QqWaWiVSQBAryguHtNlt9TvC660xzJ16+IBr5VeyCtR0YTr91Sf
2nT3HPkuX/amcZBccL3aXjjxZNEiFOq1rG0cHpcQK/3s7lcBLmN1mvM0Lb9Ih6RyDTBC8qHHShsm
SpIr9PlxuvMjtg2de2+sZipb2j80Z27v0NMWlLns1eDeV4we1LD7DCKUwGZOaXCmCpDkYV5SA4mW
0VUd7zp8m5KslQDFDv+NTBHDBlSMP9Ensc2Kjb5IUc4+WePI0OcoPMBTtT8zWNHqZvaL+Sd05jba
1UqQv2ShFmXPr7k13BKt9bZnqSedToPf9/K+jI9Hnlu8ocn7aSEPu/zjeAIMYKKipa2OoxLnH3A9
Yz7+o1NBAgcK/pj3jFWXCljjAPXWzoJO5DjGhIFd5ZLJtLdKNR1EuIR0KXBmVqhK0nRBwX55nAVj
qZo8IU0BY7+wVnVnE8PuNb0LYthwjnliIgR0mYGPT7rIm02ypKZPP3t0o1eiWXTKltrksuundAFE
VypV8Klh8mGiE3jzt2C13ZM9pwfvDdzuTdx5qohxu6q+su91v2pjb5/ouUcw6zpVRTijM/+wttl2
26ld/YAAHd0AaYaK1uD+lY9g9tQQO4tB/7W/RDY5rSgzHm4ZNzD0WTWOGUvsXmvyW0KAahTiMcO8
16eV2nCHuqmefQiqvkZLJ1itcJEmTxbzSUlQniRu3V37Flzhh7WgkSDpsyu+ijj5laVz6aad9DeK
rk+Ng2CkzTWGZpWPABlz6C6lkf27Gzz/AvPdmGlxqcL/QcaODUSqmyQTwoYaRjLq9vFJBy9ttCSE
q+qy6R0NSec73M3a54ehgb9Y7BdOavoHr+D25Llg3e+L4/leA5MHG4ZWkFCrn3ohz+U2+ngjdwqx
Xd6TCgxFb2WCrmJvUZt3BZkJ9hqpQSzf+VrlUNZG/IpSJ7683ODSGpFAhPD7K0akbX+pX4zVkh7s
zup4TgIeX0udjrz/I3OW5gYbhCl8zwvOpVEg7P1zoSFs09uqp3B563nPmxIdg5EqSWIs2DfXsPmz
1+JToODZQAFJwyVTCvpVRW0wofG7dSL9fzfXhNiUSjwCT8TsUMVYcPGO84lmPQCY51M/ZfrQz5jm
x7aXgPFeSDt73+x1A4uauDfM7R83FKfcm06HrcxKxVMEEArKgRJa3jDLkCT+ahS2lAWN4lXJ/Aig
beoO3mNvfpWLeN8CmGMVU3dV5q5JtkRyDgzAbIcZlk9XYVbh/4lEdIb5gvEhxb1nkEcprIWI4Z61
oRPV7f79Zly0A3wLuxgmfBBGATgNv/+XIf56A8LNxUkqPfm7Ow1xzbC3Q9q/qHKOew4jy2ikXjY/
1Nqw/kuV26MrUj2Ww2gemeKdgEtatQrPsfTph3KXHmTXvW3vZf2jLEU8SDf5mGEOugidJggxJX8Y
zKDfn7BBIbisfpTTfGXCRkpAqXzudMktnLkIGtYFJ6+MG7sbnZdePsRhOX8yqIe2cBv33qncFwCN
oWb6d2KHpqZu12V+uJhoj0OiwzyFy9BiqMzSpcpSCvjEZQEfDNF/XztPvUNKjaW5igqbTCzydwKf
tiq3pWU4V6jjhF0dqB1J7pzUNfaYluKoh/naxvELU8f9y9kS8P+p3+Kcn18BKNwq4wUuIVjB1Ki5
qHoWqdwlETgRlF1yBsARzRO2c9WgdphLFSip/aApJ/BDkeRDAb9ebwhD3mrPynmH1lqrr99B520l
P/s08NcGAiBrgECiNcg/5hrBFpr6zlZUiG6U8kWTrD+M6ZQ0uK70G8WBPBb4virSj01/WtV0STev
3gp55KpeZfCa/BbqkI1kRXQWrYvApCAg1Zk1k8k5/LZKIEsmQLYQXDPqKVJwAF28kX3CL+2OFxcK
mEKewRLtVePYt8otcmB2JYGivpabxP5xBZ9M+5cEqG3/d5hkIIGvpo7Gj0Rg256wyHi3BCmRpmDF
+u9OW4N4otBHiZBmbK5u7RJUVQQxUpKUfz2ndOeQmy54dScpIBgB+eX+38649AvJt0hwuCMXv2f8
4NgLmrGE+mSo/DEemxwWcGa6azV6TP9KTuPE9furHN2PQt2c4XkHE2pewFojAbfaQiyG7CjV2R76
OHc8jwOJ1j7u53r28MrlhQ8k1tWob7ARYLGd1s9nwByThfP2xeYGxfhpiUwpPgyq9CK6BhBTKE10
W4pPYyv8c2TwHgvf9QS6BHey2RRZ4ZwbGCc0kElnyVyqizz4Y55GudK64DJ3VIOz/7LBU43dg5La
3K6Q0AQAkg+5Kme/bIsnQ/YLGyBUNo8wJ3zH5weK/X/MRpnhMReTB249ZqHqPuoJnCnNF9fi4f/z
kbGCDhc4jOR7Ngd2t7N4606YnDHgOxEvuPDglOyY/LBDBBUUiCIj650Z3rHoO5XNdwCrPV+0OGO+
e3cnWdQxSh+iG8kvSlw5i995fePigNEk28Jnl5+AKV0ssZfSpZgpCNXJaPI9tszNspNGIjlgGy0v
qRuZ0IcFzDibq0SVVbd+KkLkCCftzp7pfKp5dZKZ9LPwI/iW/jGxT153OpgfmVod1d1y+/TKGzPf
ixiHtX04JpVppAUwjvPvvIZTRNLCd8gTA9CU8TL6rWyTHIT+FlydnWwGWJemZo6tR92k1sWKtovq
d0EtTLQg/Xxfg3OZHTncporCTjDlIg0ShOfMdkE5uHTmE/ao/mwr9zgd2d7pU+bHjN+p+c2/vC4+
hBB2TVTyKmUrDC/bWAZ2VN2nb6Cd0mmAcA7MaPr//lUSkqWJboA0YSWEGZT3X/sRF42jxki4aoQj
LBhr8fLF3GkuR6zBoT/mUaAtcbD+1mujoxfkCjYymWxiz7LpqYazkRP2xKwP28GZy9gyODRlP8Cm
aXB+He7jYgFR/f/IMpJT+Rr30fPuDAa917RaIamdMBjgd/Qlo+onXdPDmyQViS7PxLFTJjNdp9Zu
W4HEDOKN/Ig6DtW4nJxhEEChH3Y96BdnAqk++WgIrq+ad/GKHREd+Wbe1wAblAw3EQ04Lf0cnhzB
wWJhriGqfhXpV67fq7aK+o1CBRDJNrWdis2qdO2qZvBEz59ve4FFrCLMgjFXD1/RD79rbz1dcCUC
i3tx4cth/vnhCsPbr3WDkAbAfBsspa+9q029S2A/qpsUOZllOA6fXTvRuvdEKeb4HUSt7EySoVMU
G4PjU613ZvbeUUSbENQcLjzWdyaz44MYYxbBzE9gf6TvX1zMHyeItzjYpi2z8QYfgcJ1MHCmNPmR
GUAZK2AyJgLanN4AOfuimTXsOABr05pFETJQJL35XB6JvureMq76ub92zkZwJ3+9ULh1lN7DH67B
lpAb1lCEqdokQGu9oZ6j879bdfj27beJU4VR1Uw4SawDpsDZhFifDJHMIEASJqmzSODxMGzeKscP
nFZh5ysKd4sxbxum9ih6hurLAkb5X+g6ZzBv2iFYoRMkiBjBHoFyfrbECq1R2awRmUW8i3CIV4Fr
iAZ47k616Asu4U4MZPefa2YLu1EZURbkXFWfN12HYELokr47jSbl6e9S5gWsS9ms6ZuExToe6rT7
eZCmk7v7lr9cAx2d7P+PE/jFj4pP7KZEYnjCJ0OcRBUNeGcnaPahbrhC3SeOvadwg1QYxDYSQwhs
ccL+C5afILfzNxEtgtiZP+DLmW516HdnXjHU0BpbGQRn+bpMTYFwrpgKsp/EXYMYQ1TQGpSPy1AZ
yEo7p2GdZd5C69vsrMb6TJV+BpmgqrsspLpoUQnvEw4+LRRj9oOgOEYjkGL2DDHJNcCNElP+T45G
/cwt9LKsQ/Ytb0d4EIWiiZrEMb6LjXSIURFPVL6P466E5URIT1vxmsWOP7BUD+yQd3yD5oapFukH
WMi3coUCr5tgjdDAVmdvRWHS4PaW0Je7AN0E3Gm7NvK3DTfNEbRIwbxaGj0PP/NmRXlZwFY6Df5n
nIrZU7eFKKkHkmraAHP6O5pJEO1mIqo8HILFl0DQFIn9wZKqxy7bcPIj4DUjRX15eoWAdwF8KR9X
7Z48qSGFu+lZ8clWPKD6cezQrA1tmJiuIx0XnZRzCXlw7WszFVc/jI24gF4GzjNAtEmlt9xX2fc5
KoM/36uevTONs5PwRDzlHPYU/eBbKMVSA9GZyCfxZl+NM5C+40+gnylJEYlo1Hxb6EVsUjlM7SRS
w+trFU/YbvR/B0qNAaAWajoRAuZmlai0FDwWYsUSM9zdRdoP5ihSJMuv4VRng4/2Oo6fztB/3QLv
VmwjniOB/iVPBzvCZ/s1ax7eCwgoAKLYtkavbIW9D59hYwc2k7ia8Pi4DTlBzdpPZZ/ZXHQ/ffMF
4jm+ebLhieF1fUih2L4KstqjG5pR3uy5u/FFarBDvHNQq5mqXBJnjn3xjEMmZoF86CHYDBnWPhUZ
/dGYF8O+mPLL5//sjx5EaITX4TSOywKxrT6R2Hu+pnlRqVkYVIzuvUWDu0u2TepEiz4/ukkN7jTN
M3XKxYsr4HB+9IaR90WKSsmI3jeYkpUjWbFY+/+fTbT01NikGow67FKm0vQyL47TPtbIcTrc5HFI
lEa/Bx6YpzMipV4eE1WHOY3YcE7JZ8zgr9NKKZQ2BJI56dN6Ib6ypr+t//m37VYnjlC7az0mOUOQ
PZHc8wVoBvwuat4ZmSwrBBW5hw5zInvxU2fo1A3UoMRzADuXy6jBJkQn6ISNzrt1QiJdnKj/WOFf
6zHVFpYIVswML80S+MTY6wFho4J2nJBjrZXZ5yI3y/0+HyJmzY6PMfxqFZxQwfOhVEkLhQuIi+f3
9lrie6+kBsXhAwtAQj2Y+bJSPQtzmzGVNHpAkPBC0vUYb43dTBAMVVMmtXOM+54MdBPlfpgH0Yq1
1pTiq+4E0JJXO/6XVKfDZniv2rIjWRWPplDeiRCwSgjLR2JR2kPqz8RmBKm6Sef2QwyTDNMHT/GB
JwQvBKCqwoK5osxe5j97T+1MlPQvLs1r/foeRDwjBtaqcDf3qXR6pEmweVnTU7o5RAm9Uc1okdE+
VFd6HvzzgJnWFN7j60YI8HZ/KLHSOnJWlI3vjt9YqmBy0O9yAMrxgRsfgTr1qdURC/ZQ889fFpUT
OPJDHRbPk34IaNNJFDd6kU/GS6S7xfVhtimpncnqpFh4lmk65gU2mYQVARvdDu33RK0Wbv/x++Xz
QoYNDHED2DufiPaSLyNaEadT80gGPehvGkpDr82rz+sTsmi06rmXS6MXyKZN9KKN2HDhpxAtAGjv
5gB4Gzcfa/E7YyU+9gkxIJMvlcFRTWyaWx6xAurNGABW55vSIM2tJOuRBmgxSC0EbHvwsWDPKx2T
BUun3+tf1sm3Jn5NjRflA0vZEXA3X/TaYLJT5n7QjUmEXVsJo617ODMGdcZO+41YzlcObgX2tZkl
QV+7KFctveFDfqppzDjEqheiVejiS77/PP5f1XQfTqL2ZQi4nHWsgMwscXTW//yjfTFVp/X3GB+i
3+0ALVtuZWqxKWNiPqu15KOXJBk93uyQfOVByES1Z5G0JJs0G0dFTx6+zPTL1PFD5Qhe5IfCkpdy
Q3rvabYS6M3KRqSV4y0lEAIOm41le3ZeAFBrHFSulRmg8NyMLgfUP69Pn+jihTF+zjOlTA+dRKzw
EMCuNl8WR9hrNoeNf3pvED081K5jAGWo5D5B5yPX2xgImKaM+z40xAGPGFICSxVRP7EfNF9YpJCp
WwjiktS9KZ/+DYBqk6ohkjyx71o0R1pkPLoQ8TZ8pb+5VU8x3Q2C1l+xaJHL1CszmhElIqqROeiv
ImeN2PaOU4IlOsQ9fIB4Sj5JBhTkM/pg3/K7plfbXd+Vwq+8Lwc7QZgKebf7rVXZDbRGnZb2YGn/
Cx2dCJ8IiWIY23MOk3m6C1zL90KyPYeD0gAEe6mJEraWHkDH2Hk9xOLy+8smjqbnRJIflcj1qCS1
NUMxQUC5Am8EtVvoUPcfnMqc4DVubNpLp4jgVtW/E+3Ows6xgPI6vVMS/mUDNiuJu6dt3y2AtOG5
f/QZeTeAVYMBIUL1yE7wLIQPL4eXLCrYo5FZzgcXAxWfZR4HJHnfrp3qXmrxMGaUyUZOrlPBiX4g
y6v6BPKNaXnI+tJBscM8pqCrZ8AbJk/fTI9WqYdJfO1AtPpwr1ufTrdvWhEz1QUt3uQpFN/U0Z6z
riPM61De02eyCRvfIn02KF2Xdjxw6MiaAUtJwbjIrUbbXOoL8HCn2Dfm7vh8pkySM4muK8AMUWm5
HmrN/o4ErD3qLyHPjr2u3g0rhvsZUk3XTTlEmCf7HDdebKGhPN9D2Elv9ZD3Qrg5PGwOdheH7To2
FSWppH7CiCGLDqPFzelfhyIhLQHV3wsQ6SlwNaUkuEpZKm/wxSE3PCg8XJ497ny415rD0L5uXwQY
yEFfnVoXMI876NjLeWhtg8lZG0QeUCP37QhQDjqY9rB2OovP7vklzb1z73NXsTSe3yVWyLTDcet6
1WzdEss7BFf52WKuYNKonYuOhk1WW7voZiqWzMTSgej0hxeuvh5iJmz7jW8df6U1zWGpC0hhbEhL
9XFq+7vJYmjCnaGV0yt8Qt6Qk1f1u+hh00aga+N3C8BybCMa6oYJWNWXzBg5GW5clXleBQIENY1c
OB8Rf5wVyyXwnk7XNXYS/JDvGc07tQEr4l0xpuu+tcyOhk2U7NlNd7/8iZUM+7o+ZjYaXDoxfGp+
lb5SeLJ/d8iQx2Da6T+6U7E+4WBuqfeIqRXHvQINOYMJNU0uc1szK/g4KhqTX/2eyOn9fFTf4kNx
rayEFD469pIouA+c2cLcGhJxAI8yS/UhKbg3drhcb/TeJMzhfV/zklPRfkDAx/BsQtYiy7niZJfr
mshUUnptawtBT5AQxx0hmkjZewTdBgE/rJPjLl3FLTqZjjDcENn12zwbBX8FYOtRhyiZ9iiO0v9d
KKCT1cwcD0KFKxvFNUsXgke9WMemPK5bQYskquL59Q3hLkgsrhQjoHVN6UtnjundRoRMLj8xDaeh
F4XTgbRkH3GjrqDeqEckugik6Jx8yNlMbXWiNrA4YY7LyvYMBHoRZnd8y4qvUVkSSM6gOR7B+iG6
Hoxw/JcTo05z7srp87NRHozS5GON82FvLZHCJPAVPboaVRNmVJ3e9bnjYm0OCWQajDLGatoRqJ7y
QPNQDoceEmJ2iMfdVI6JbTAsTRMh5oXcxL8tt89l4P8Rcrlb4KV0+pfHqvD9RL3QK3ZsaG/dkUft
i1nw2y5+GO1zakEBXn8iTUbfXjSn71gxNuMHuKiVmcbjA6kOguuvE772fZmtLaXNjBM4fHv45DFt
W/LEp1UYMpVixF3G9AGEeLwrtUBiZn/eY8l6ZxajeSlJCQ9oZjhBdnVXoLE4bBRA1eYhSIBIZ0Ew
k6ZC/7MatNsJ/VQT8aUXuxOPUhSBe3MHf2MPCadDzZVqmOXcsUrFVQQZUNmdUPpe0ynJ3yjSxDLS
1WiOuo4WTkvyXUj5M2wqdG21/9AV0MUgOpY+Yb7iyCdQokcYMwoV5UreK28o2V8p/U+NUR5m//2A
8DomsOrkbk2ZbgDvT5e7DubWazFfdPzNU/eCIiKPFFtYAG++B7r2Jl0C5soyIb3MbBusGOEHg2F0
ht1sGxedExkDNWflj/yIiSocZZXsV4pmrmU99ANsvFjJUIH/mSxX9GVvPpy6otHge04yB/0wGxzC
KXGtl+/l/s7zvqvRWehW60bpmY4HM3LaTRhRg/aZbvOfDpHXi/f/r++jDdox4OENqQYILaHgrtp3
w8SuXHiEuQA+LtKlCiZY6P+IIbAp3BO5VNjRw6/VX5HJym+/PDnLq1BQAMfRzrbmWeWVTEao1rxD
NTpWVo35iViICpI8xwzqCT1aA6FbNsWNyqiaXxBTBIY5ww8tD8q6gakfru2gxCzjb2tZKmDS9H2W
Z4M4v8pnyopsP4O5pSpbBsxHE4SVrunY67YDddJcVicX+mnb5GZhKAJezR9abNmNL8iuNBVtCJdo
1R5/pWZUKrrfLsD4WFjyLsZqcLtGOMW09I8DdzqIxjXDQmRJGEV/p3cJ2QCAhKVYr6e7WYU9MZds
keo2ziCuoUwD1LiarSCsjfwa53f7hdmhc5Fn+kqPU9KeXK85cEOI3WhPxK0NF9jX/s3H7jZrTW5j
Pknwr6oJw2mMBwRJ2kJeLu9YrAjgY9GsmvKInX/fourXOrOIlpW+wz9pVLaDJSjUS+DqfuDJsTQo
TYKuTvYsOId8JEE29pkK0cSJuan/Lx02o43yAZAy7o2eoIRvaMfNmBH0/bNOyZ/EJF7VqpOgo9Pd
SK1AqMnXBzz1T6LhAZF4G/6ut/+2GSWY8vMph/wlyrHTzaJYgtJ5Ina6qllRdo3n0fRFbDbSwVwa
8NA10m9u8/N0RDmZh3UH79K7wEccz+xq0xVltgfO3Tr1AvV9X5YNIOX8p5wR4wE9uYCpL0TMwUjC
1kwD2KM8yPJ3Gw8BY0KmzL0yMx2LgeWiaIamHagTLYmEwPceXWFCZV7rN5T6AX8aX4786HUV68IW
U8viFJrtj6kUClzfjxQ9JkKciZC16A56cYzZJIijbgbt4/7I5AtF1NOXIZ2ZoP7jWhxatT+KplGW
eAuu+qI5RXNrGs5dvc23GXrACrzofL9cV1VXztNg9qPsAnTYBdLdIkBwT6bYGR83i8c8DFHCDv5N
S67KeMIf5KdhUVuURKOt1ZyXwz3CkciAk8zpoZ+svud/g3VCD3zVjc/qjpMcdfYdxJESvUgvwR7r
SxGqLPEUuRRdUdg5dqxgLIEnfHXguhFxfd5pRgTe4oGYP8RIA0eoHVnER5wibf8lSvBus/nZXBl9
kc0TTdqTlHGhR+VUQuUGYHZKCVds4vpHq0Te99PRehtljp1CyhS1I3iDB3FLNK610nkREBHBagXt
ZvFBN3vKmT6OPX+sybd/eqXtIXsTeZl6k5Ysyy6nhbgNky/nY20a2Kws5/dcL+vm7X1fD+KXHWzW
zxNNUUaRfzyNI7vQKM2gp3PcZIA1HmyueP1zcAefQFD7vsQUPcbn4iPt83l5/i8tJJT6DRW3wAHR
9KEXkQKfVJHarGkTHOq6V1mYYly7CEiBqxhrgeaxSPPpYji7YSa3G8yBjlgSJlsOkv+6VfiygrPv
e0VPp+tSKJ2+pNocMJbGLTGmHmTvd54rjXjLHkf31Lkzj+//hKrdEOMc3j7sr1+mBnPpim+hSy8l
Hl0GWE/PrBPH2/9R+lZCftlimU5QQpJ7aozf3mKbqA9lNVzt6dOJbmswEUIhgEFE0ZLBOAjlsiru
bQGD0NHfNc6Cmkbo2e3Px1rri8SU6C6ZzfL4UNRwRwtwqpPqcEiS4Y2YRZyZXToB/fvpzuOdn9ww
HyQSnIwrnLajqd4N878E6W4oXHQJjjn+axD0J1hkNw+3zkgUuPmgb4d339C9dnaDNVArdM3rkGmY
xm7r/9moDUFcZej4qoA6PNbLyJW/6n9YPlERS4dV0hOHQBWGJjWC60i+nN6ZCxbY8MU/CDzpIjJS
fXxo4osIceBDHq5MBsZHNwyH0latcYvuMnSYSoVmJF5UMmYhxf/b989ZrpeV/mpVmsLLHj/T8OzC
2jtorWBGHi97oPztJP4ry/OssFtUJcj51dmtVtqFMGUPL0TQ4bVlQmOHI7R0ABY8idsliNxQhQuB
lfaydDstibodU/osuUJZeiJEPRl9XdZC8u7fvJUiUeluNvvwN1ZS6RoWgKwZjxNRvgGfztx20QQW
MxKaFwLYVI/K4wt/sP+2x7Y1nsyHAKtRlcvPfQ+iJyhxIZS3qcWujjOilNpE25Xvy9CfGKFw94wd
F6aL88xzmJ+yiJG3+KvoQBAXdmRHHdIDNkZOyzGjlzfWi1c9FrlH5qTb9mfHpOxm5sL+M3Cfy2Dg
uwnV5pG3Qoq11vYvxPrKFlubshb68hbJevIjF0nYdXxP8xEWRRk8TkQlVbzhgEZCPebBLX53g53m
jwpiku6Q0zIWY0ZmGM7lLLC/TNORGMmK5ilHqPa5JVx6iUYi9tRleD7/tt6nl0celkhqClD42Z9q
wJomBpNt1x3/s8FipQ4qPfp7jSPGeTzIQT2jif3EJyxOQKG9P9b0HLiDMtyPtYODLdCiP3jBi8mi
DD/t1+wrY8GgRri0u2PhZQY6HkBfSB4AKoNGDDK0u8L5cgl6H3zdXKQi2B/6qwnFVbkdptwlkfSd
GqGJpi1lWXTa4ObBVE3PYjga08+5INBjeaC/RxXvJMxbnJBqtvR6tMhxJhVoB/5fxKqZ5dQRv+DE
uQLwvXbGFFCjyiuvMn2/4j/nT8XG/2f82i28b4e+nPXTk5I817akuriMQQoDtyCS0uMEZ1ivnKvm
Hdw3MkTJrF0gEkB34UR6jVyGzTKsBDetFLwn3hK5xnt965gwHaQXyoYOogFOAQvL8WZTT700wkIK
GZ+oUhh0b0Fi+mgw4nkbOVyAJ1AOYVhSMhEmfV2qr5CkgebWPf/xBGZtzAG9cHvda0GZbGRZihTE
X62UUZWxxoxOCY/Iv8hkITlFa3NUTxSQ3vsqzHwazF6NL+j3V7OwKsF7Tr9+kNqeA3g/YYEili/C
SCSGY9MjxR5aOC2jXL7ADPlrVjsDj2WuU+8BN9u7cgIGRQygTUryRyRXURuAvhz1L90etezy8Qa2
xA0lQCX1npuAre+33s6dFICvrRb3e/+KWfg5Gx1+qBUaciu5RWKV2RIwPrnwKQd0bt9B7LX9te8D
XjdcmkgYP7IOJs5oZKOIFgw2H0rb6f7BRq8wap3DwcN32wQmSuM+WCvXxh8R5qlXrpDduiWQsaEj
RY404/+8+UrF97asmzs7wSVZHx5Q2UV4HCfMM8+NRqWK2I3UaGMYtdYRhrwmTCbLQ6vEufhfWarW
nsq2020BTtXb3+c1Y2NidM1HYKyPobjZjmumDJsBbIpNMdOALKCdOAvU24ETVke2Ib5g7IxdW3gE
6jx0b9bNzSZQz9oXyjMFpHCC8TdKj7UlJb8ak7crwh5HApY/UnyKNr5BYzMKgnctiBGLikDPpP1d
4oQ6gY981kYPR5W4xz3eChyMlWIOEMNy9x5IBxqv1wf4lPexWHof2/rNwNiHkQegmvgg4bSK0U9y
Pqkarc2Y8dRtdnaR3A3SsGXI3QcNlim5A3S8zpkgHhVYCX1ZmZEdItRUODrW8oHBlmYzmVeVbdS8
KR9P/MtZO204xCqRjj3A9Ma9bfEVaO3hxybwlh3rNNmfFqDXHsPI9A9mv+WDOb7nmdfUkYngO56o
/8nEL7B8MEX8fq2Afr7ygtXwPJJYR5quKOWRXQYYGZdkRDNi71ifwzvcAYvNhlXZ8LfR1XH0j1sX
wlaq8YzVWXtCqF2OxvuqDI52+2X78Ile00zoEJ5bRI3fje+wSldFk7jWTnoMcB3YGoYK6QIGptYT
I2SS6EeNLmnTzV78Y66k05ZKQypTfIncSVRiYNl0h0/rsiEaNxc6EF6IR1tnAzW+UrSO99t/i0Qm
SE1of8ETnmdxXzhNRvig8HPK7sHTsSb5Cauc9kqx9xB50N14zQhLOMF17EsglVc49a0+0CN3PZAx
B7SxoS6eGNOjMNK5ePwE6Z+Ywtf2liw/9h9oauTZ7dlmPU8xf4cIpWoM2oc4G4inRA+LLbr5d2UK
pymvgpGEEqEpBLeIaZCnlxBKRa7YvpeYBzENn1+GpUdrok0y9/o3vmA/5wJgBC2M31P+n2p95fMq
EBg4Slc74pyViywvZ6utL97a3PUF/B9ABbPLyERLxmMu6hOhg0iDtIZo+OHFEChSy5qK4o/rqMwk
GQAsugZBoyHBntoisJmSOwHpzF4UhjB7gV0leC8CCgpt6Hp2O/32mmmv8uiV8vndo7GYEX8RjH2y
RtzQMyLHwcjLcLlSXS6zGdrZu0+XiSTRUKIuSuVoS6tlwjlUGPQcLn+TWeemhiMqp8oOjfMcBE1B
sp1+LZMDTmdM88Bpi9IqCY+K077Umye70drqRvrZ9itF6O8J4jN24pbf2luxMuXkiShhkSa2jrgl
mU6vRPkQo4f+1byLmQs73ltKcIGLjFXXMacQkohOpbdS5TCv+L6GVF8EMLvlmyXZhaEEJ6YBd9C0
wjFjfCX3G/z3tS3WrFs3h9oHp6+F0L+FYmyO3gs5z5KcLrdUwC7+ZLzw7izwHLkkqeOeljL34uPm
1fDZjnOkQyA4BjCDRcyGSGxNrggHHoYIxkevxu9KfzuEVChciPgveb0QPG1Y62PQpqQ0xo/ktbI5
+fZrGyK2VnhaC5284TC0oLHllF7qUPb+n9MuCqhrMrdhm2XKlXi5KnQPENjTQkEim774t+fRGQVo
ASDP0vdaRrr7pDkVS2MHuUP4UcbwKlcGvMk6T8iyCWnkup3p23mPXE23Qy5PYJ9TJtqmA3AmskpT
/73ykt2uWO1NCYd5Dvdi7OaVph3F65wBMEE0Kh48RK49pTr4b/2vj9foG/nbgwy8hR9R/XW9RICi
b/Wr9BPKfkNOCRyAfcSlC6uMzmKSvIwhZz4LXrJG+hpqSgF4gPvJXGq1Vmbd0hZRdfwjHHfGSb9p
B0rg4mXRXMihNtKT0xuyfzkZ0cZ2469/ticl3Y5t/HrQwnQWYcTw6ihNPnfcBcQLNlJGoqBl78yp
w4x9hNUZ1YZldSy74LU2uJ/jFCkb2ZwgtdA3JJ4vur5fF0BvWOHqZ6CCs53nd2WvRAq+t4zni4Vc
JY7q1VEReXWf7x7ipjLI/zVOPpY/9NB4q2sEmKJejpzrQCqySS0OdaOElTrXaOdrldMkL2xiRZhW
ALF54gHZFG4b6q8WTNhe2uXcdtLoATgXe4lSw88xDBAzlWcvQFY2OHvYspF78g+P6AOZGgW0Fjbn
k5Wjt4gTWNUsVhAiYXTrwXjX/0Fkna4aj8vZCJf2dN5/0tQz1YStlRhjtIFTD6OvBz75aWV8BXiF
pxczNzD25DjUpSbvbWX7Q7pFn/XSj75IBdJexdPdo4F7POEufGA7g7MtDwjjLX0UJQI7uCKR2hem
aOFVJN2FSV84fbYIZPhVo7FD2vyz3BUqfrqh+IPbtBjHPcjgUv1BazDLwi8mpXWJM5m9rrjf/pZQ
bzX+ZTPQ+qe/PzE6qYNO8bpXapz/RmOrmus1DozVBe3orcVit4AMBReqE+V9GbWmglXg27No/Bq/
kHpv58CBkwvGwIBAtXAHhgPKroZYUIplA/jrjDiDRPr9zSmZBS4RGZp2jz7E2wW5NzNM3SFp82I5
E9Xl25h3+Qx5XlbsRolquQKJU/2GxDnxutxdcg7s4rfHapKrWInj8OhVrw4r+Iqa1icsSzMY5AYk
GkQFHOHkLsKYgvoldeKCWb0y8VD51/I6aRJbFdYn35B+z2RVaS52daCs1DKs7qsb08xTCaWqxKpt
G+4xA7UKp9ksTbYzZvdGSRyFtAMVPstTB//vAijNBuUAkk3cFcAoQRvZ+sBhQK01Po5oxFCwFmc+
0enTmdnb62QXGWGuRBZTz6PxR7UhwltdV5QnY0oGmYjl1iotpflciq14lg/nyKPu1Y1AHdZnZFyG
InxqSjdwJr1P/w5WiRB3PPqZObXtdnMRcc2mlYorjJHGNPEFc6HlKmTl11QAGDJ+VYPp0urAVdWE
A1A8mE5lwaZ34sWEbWCG7bbz4yRSaQWSvPz/yH16sEjOdIcyOL3ciJkc9MMEjWLknYDcHrLepLr8
EneqdirHEHItBo4BFu4olBaarfRQtaKkHYaGogpIDUVbKrMhPZfqGEzxud09eMIByRtYT6fE6//n
YoBtie2y/0D3F6ZxUBSzzzty0z4GB8P1HqyGRFiFZpUKolC3q8+mGbvnDKrGH3bsdyLfbtLStdFM
AEZ0eoBteYWg45fw0mIp/zcshim/Aab95+0LRDnka6RxZZNv87BrGvfSmOGbUTOOlOInMgeexmR3
2lABbnFuQRCr8/5jtdDlv9yamtxW2SZWS1UrcxsCJXduuDfbYRK5/e/0ocpoMkCME8zDQA/L6f5r
H+hXsl6euB+e/z6l+uKQoPcbWYUesJ1o0ATjKxllqGvcyWkO87wpqaRcQRC3/96QNT6Aoi4bhaHy
GW6Nehptoc8XXeEc4NP4uhdk9aemi7dhKpUHRrVOC/iSBBe33ditfPV5FfakdgDshZEY67/2x2OE
+w2FFjyEihBCAouvyR/SuSZjmSBOmeQh3FbXgk0zBXWab3SevI4Heu0flC3R3sIjibJ1hBZrMEDk
dpvfk9zgamtT7lebZbs/Oe8CsD++hNVy7O9OSccFqGfRcMnWqGBWlA35810rN1SsfBjN653s1152
AXeSk8cfqTMMpGGHX2g1V0lotLM0OrkbGOeH6iNlous4i+juCJMWJk0i2XO0PopKE9HrmLjGXsmT
+eMqqZnbnJ7oiLCdzUDS1VZS3PDrcVh57JleKd7g8FBq9VMIzzsvp0DICbYES9YehfdpZJwxJEHO
OiAV3F3dlj0JzKetka+vtDHXMC7sco6iy2d0p41KbTQxbwO7MbCvlKMD+q90D8/TWmLTTMuH/8uT
m5P/SFik/0aMjGh6s9ZUqHSZzpCtQD1voZNfV7xydXZAb8aVEhOI4sX7g0oeGyT0codjJd+aL1uA
4nfxuBGNUHIpMhbfDyZq1LRl5sXsgHzaae+Ka3lkpxkmX3LdHnf5U4147JFrxHvrAubpaUA3OWDo
zoBVDRSqcZfMa1ImAxMYDU81YFVCAS0TVS6B2IIvxooOKxF2fE/DG9t0+5DQiS1YsZaIROJ4yLoJ
Usjw4aCac/RwukIZW3Zrq/IpAok+9wdWMolHGvnWkur3hfkg+RlH6ZoG20WS8gXFmCQlIFO+1P4V
tTa+I1gnFH5COBQHKt6V9nEmumMIW9d7quyyG4Nm/+VepYsxpQEXw9BTk2V1neS/eKt1Fj1Az6RK
A+W18IjZJZHLiTGO8KVM1p2NtHiz9SwcNdriOwilWaxkIz6jGAMLWDuKc3qdj1TYxp1U32tHbVks
FhQkZD9DNd2zqnobila/oAqYfW4i5tk7rTAmg9iBC1ngIqKXoZBGs1tPM8x6H0ufoxBbcGQZe323
B/hbCts/Pw1KmkGSwvHqkoDRBED3hORX04JSu9r7pUMCWcKfh8riYnpnpxF9o3PwjN+5mIQNJH5C
qq1ber9gvuLXUoLmk/LSGNB3l+PfCsL0WBzBkgHCZftkio9886+muKSbQAis0BGi5Q6mKAMTi8Xz
/M73X204ceZf8+fT8eIfG1FAE9ZvsIrCmmPhSOf7OO/GGVprShCWDeSzIcTTMuDzAsk2/HbGur/a
hwG4N2xEFpt5PsvMFpiFtBNoFTVZB9BbsGkLBGLRXALLg1zw9L4sF50KOZgPmKRnl+koYIkoQsJc
U15yMQm06cz58lV1mrun4D5AmgGEd+DId+t0EgxfaZSXaUeEMDBpn1RxvxJ4ogvF+UorryD+z2/c
CgwrYdKI75n4MU1RAT2yV3Gn6U6UB6e276sluHX1Iw6FhwMOaVGihp30p5XSG6hdgCVzI2RY+Sx6
uONUW+5D7IFoI/LJhJViikRRNL7dm6ggDcV/qI3n78p9LD1SDthoDX16O8f3k4ZYUWij6YSJkB1o
EMtRzC4udglRbolJeiOgFueuiGSBluFmxrLcxur1kgTa5LgTm6b8kPeAC8O0+zjYqiNe6eFtTBD2
KyTWX2hCXkV/frC+nfGIcGPqegpRVt1olOY2n9P2ifjhiN6Ji9XEdU6G6ytfkfINZHQHsA+WjWQV
4UJuJmQY7XTt8j2VGvtp8LUUyAP/QvVsn+x8H460b4ImlDecsCiZF5WxZbWzptzH7K8oOtlMQyKD
sYJPALm2FOvlfaplcZHDODvtJJfRg+1kcpfq6/XB/9N1JSKyYXn0YW/qK+oouys9bRlltVfks5E8
egE7qpBtVDEu4YDKeksdMSoY/OImKUUs0SoiCO/ahtibYpIvq589ZU6yD355NkqqYR95hFOsBhU9
43nSNDSGqnIhRvpMfG1Ibe7JczwxVRu3e9O6nYQvN+7RDoDLcNH3Y3hXCQPHdAjXuDazBhSX563n
0xdcaJ4uLZ+GoEdYwS3ZMB/kBvnb+O1yRoPfnJwujkPinGB1d9PSpGgQqSjhQsyc43H9rhIOPLJz
vZ9uHVF0lcyZqSkr5q5wyCA7CdDEUqubGMy4NK3q3lpH0aarI6AU7yraHX+2stZqs+AK+xseNdIM
kO5/KLY/5kn3q5u7xSbx4JJXbamgMj5AWDx1qesqVj4jWOiDRcK7rX9UgEgn+/z16uoQYDbi3rWN
H/gpPkPwdOxtb1vsFEfBJzeIoCZjBYdyJkH3NFqSpfIrMCfSObbbIjNPT2/4jEuVO8Hlw8MEjhus
XnxxtbYDCoiMNF+hmTghs/zX7R+4zrNIxlJljK+4grpn4PMAre/XM/tH5fIvMTtExBEewBYXoJbG
W/t85rpV8uE1M000iRD6QYBOHEGGpqg9NQmcPaxJQSy4QFJDGjEpgI1CtvboVVZQwcd2p/w57nsI
x2P7Dniu6520L7CnidkzLSw534l92bWyEqP2hJshDIO2oXgeu4vrz7dR8YdLU5/SEFA4hx5MpzN7
0DmKAPx5af6D0V0w5a0YIpaZdHCLqtj2ph4GQ+krUxdQ2N7VFW6gEw+gNy0D6TV5ZUTzR/+PGCt1
8k7Jbp1SHVenwuES71aRAdYXc63GQhautKzoDCjuJmv7tBSqMBNvygXT+GINnjdoz47kaWgZAWvW
z594j5/J6MJUVtoNPTXEs5SzRfVOTJIAAViuKT+JW/NuJuvAvQwAR9yt0rPGYQf92KyHJXCKufd1
fgZFfRBh08w3Im8VZBT1F6xHW/d6P6Tbh9C0s4yr0b0p//j9PfA9obuM5nR3MEgBlwONeiKvSEQW
1OmChvry3R7WAiyUMx2Rih5hE/P8a5vOGQjhUrJBq/EDGbLX4e+WgCRN8mIq+KjlxhbRr1F/Vgnx
RN7gZYMrUtJ2TwFwQTZa0mH8SKlNuaoB+EWSAksNDkgwk5kEbJL53lkI1S65aB0K5AuOSpB62Npm
iUFYep2C2NE5NXj24YKlilKJmR9Elnr0G39ZXdliJvxaLFxNLtv20k/l81FM0dXNC6BI50Bk1fZZ
oLaukU4dhUUqT0gHuq+XyzG+OLeWk3s0BA8Fhlo9Wdvsl4qiC+eZRFwxuBqO3vIrGKy6BaMbZOQU
KDG2RV4YrYFBFemx/e8Jn10jD9cJVzzqJBk2MKRzCus4l9WRoRqF8bGItIps6aT9doA+SCegzXOB
J2we/+MAVXeqq4g7v2uvexgtApLPlaeJOdWLbwgs2VM93YB2n2sE0UXu/Tjp7Gh8lerVgUeS0LpT
lgJPxQOGyniY3F+O39crIWewV2g1mIvazkdjAiLnRzUvGTO00f+3PbAYZrfhW6X+2XQK2SaE/s7V
mNq7O7aPTXp/VHL/6nmAdgXYABnDKkPD4E16/598yGZhfqkcJxnrRx0Dgg7vzSwClPqiHZhCN043
jlx0b2f4jGCakJTiqKRGN1yIYPGe9uolxUBelgLpycoAR+F/6t8BUzhMaA5+0GdYzr7xe9ir6ug1
nkp811xCphaMEhciABy8DZOysC2PiMWOsvX6byCr3BWq9O9oky3RoV0MJvcWNQ4481NghOR7vheF
FCfKyYFB7T+N7ynrzWoSgBwOBfh6DLAl8SkSRfG65/zLjiHCB3ZGq4jqoRyv5NTOO+ZwUppW5q/0
s3TU/g590fIC1e3/dm+oB2GBzgU08GFxTMLVBv6HbECa+ThMZlWSxHKF8/EtGxX/n5/7C1Pg5Vgf
VMHAxTTwm5hK314QE0tJipwP/+uzTaDeG87zIbtGiO5jsqQl4TqbReoADnX7x5D8+dowaplPPzkR
OH8Tb/8LiYn5VDyHXo0Qo6azhzHA1I5mrnPpAYHhLmvsP9XVEburCRvJQXmbjwOCQnobE0N51OxI
hngHb1QtifuY7ZCnhg663B5zb0NrH8sBp73nOycCM9s8dUkLFCI6KHamFs2yCleC/xV5ttkNoy2A
0REb9TIlWeAoN1Xa+8+X1g8ZnihIVX0HK++AFTpRczc6UjCNBqJAonMCrwQbZVdW2UlPbdtMcOMt
+Wm/DTNX8ec7TiZn332NWRWxK36RhCvf8PrkHd/OjVaKgT9Dab8jv2Ux8WkT9QJhQKQxQr7lCMAh
hIUg2jHW1nFsu4CH6mjhAotEdrm+CMhjfLqbtgj8V9h/6N4R0vMfGOktWGSjSj/stsWjGRVLjMMa
egEXBwhsv+8KYdzGEfb54DxoUVp4nJtQrfVXAEx2vf5zWDX2SR2ToMbWfgWBQcbZ9FYH2/UNu20o
xsdx9U51sMxPA1VSfq0/DxYeS5S+hF8gRSLMbeSQzSWp+WbZaw1ThCRJO8jcl9Rf3sw4F7CkI+0z
oGe4TUZFlKI7/nl2I5F9+/fVAqV2tj5pMYEfckTbzPR8+2GyJ/OfTqUpy/Yh6MFjyTeH8ty8lLs3
0cqR1MQpyEb/7B+eOzd4LlsWYvU5qR8i+CW7gm5L3Pk9HpFXIDX+qN4zTGCRw2wvdTZu5LHPyIM8
m3+xcmYbgOZL7iLlOVfvruWt2/ojQGeZV3xMU2wPA25f6kVnx7wdC04Dpy2jCbDaxC1UmhGDAcmx
BcMwux+Qx4TZXO8MdDt/GFLzeRLZk+JQ40pwMDUBe/QbvXi6t+T+qzLDVWWEmY+eMFEN+CS67Jxv
xR4bWb+3Bl886SQjW4IMeH7WsLJe0A2uuFfP7qgv8Q64hebOcm4kQxW00xMu+qUTbdhOQRdhMlam
/h137eQ8UBarZLFCyF2eenspoKRs8Vh14CL/IBDLdvPGXEa4BMZlgW9N1u19/hFfITJI7LvKr4i2
plKp3mWm7LrlPjOFBrYYPySrQN8GyS/gi7pH2HiJfLpXFSa/p1J8kuxjp6MCD8XX2irQbWyURqgn
UN1UGom6vYpxqjOiwdcyGVvnDLY2Sqkn2TgcCm5uU6OgH91Ltfj0HPLAzjfeKMxBPqBizRlJVqTG
s+blT6UTFBCUKpPWXkyn8sXN1fhqcw6CqNbT73svRZlRXqhn5AqQilZSjJXwJ38bL4F8LvnjdFzf
AiO8xpsisFDtWlKvgrIJGZFLVa3uuiG39bcJkVYu0nF2vkK9eCZg7gbS9tYkCMFmLk5oZhw0OUDe
pvHAy/1xdaYpOZNYQRRCu/GS3pqvEYL++6zrS5K8kCYJswFSmjiKOpMjOS7naDKNp5wxGFph8VJy
0vx9zlpqZYwQnlzwfm0f/MGlZIdxRSHag2ItY7OTZ6FJOoFYpvs58+Al0LzRfh2ZWlLbmes7nc52
+WpZV/5vsbv3JADSSE4bV6JOnwIA8vpgdrYUpFM/36peNrHdOpZRTPYyleS6PntdOorGuCML0/ae
yp7FFCDyquyfmFzLsW2KsB1lrmcNdA6uZs3YdilUgR8OxN/t32eQqZkFfijHbx7UsndEfqcqqiAG
2Yu0oSbxs8VaMXMhxrKHGV13Gfw6EwxqRpL1U/meQK7cSmtU3OFurKXcSr1lDwWLcZCGNWZ4W3Na
PfFM29EwP4c/Itbpj+NjH40VfWdXV0CD+cwvVEVvzWyIzSXxqHTLCcM4BH3Texb9WcH/EFUne4Gj
dbwF9SW6XLxWIoGwmenHBfoE8eBQHgqpYTEjLi9LyNq3/vAh/hBCeCWF2gwPN0LxT8MzQgLROXaE
Be+O6X8BxI4u53sduqoXWZpd8H9q7krNaF86tQsqBOaKEYIVfTURSBuDqmrNW6oNYLoN1U7MkdUl
qFxMhlNCrbnfFZwJ/g43DWfMva9sanmDvP4fsMRF92h2D3W5C4xJLspknyXFVvGDJXtR017hDFFL
8skG1p9pwroubXxl2EkzOZUNm6jb3pWjHYS39tlHUeZZJC4vuFJd0zNt+ks/Ntdd1BGBy7cZ8mb8
Jdk8vxqwPjpWNcAKjK/g4tk9GK+AFkb/teXlq2gcsVxsMv46TKhokh/wdke6YtIGqKdVD0FOvVxb
JySx0nUGjBGLUZ1hCMzvvUVwTr0pC5TNSVo41b7KbCOX9EQ/Ji7VNmbRglPY/haA+jbIsd+0M2Aa
unaxOMU/D3p+gh7xu2Cm70/5SRy/jbuqT6HqG1aLI4Qd+WJFiGKWYyARUTy7/uPCe9+RGP0V6NBJ
JRZEvRvkuaNJw+YbJXhkUmmfM765DE+AMXWsmn+GmNgKQOcTmIEczuOLh+qgPYeD8URMQOJbHKN1
TvGP8RdWCknHreLGLsoUusliWOnyk4rs3Lw7x04j5cyJW0tj7BySYPp72DWn8gx0DAMoekV7ILFC
jk9Vlfr165NuOGqcixAk0JrB1vHCAU9ngj+JB8VJVrjeBwIyFdTkZys9h/aD18PBzAbCaeHgHrEo
aC8hx6WQlNQS8cdzL5wHTJOd0o+r4g0rQLRQ7UAfnEWHE2UPdpaWkpa6rPRAiAUMWVfmyG2Gql2q
EsRBcoohT0GK251XPD5hFHM5aoL6jh4OEkpbwtjKXe6UFjsV9GbaYtLteZZJ98kuWKotit/6MIVh
/Ny4qR6Ekr8mgLjBrMjGX2F7NArnRVyM1UX3QrHPFXpzLi+SKpT97h8B3wV5FIRlCXrR0YtDhVtA
dYGw59h+i0N7FfJ787BJZD06yoxew62J9UTrbD/ONLGrR05QyMwxkFWeROewPg6Hb2OnNo+f6Q2s
pGuLzgcP14rpefUlUiEVMrce1VbHHpV1Sa8OqzCXvqUMsXsGl1wsBe6nhWLfVXJUwmyFrvHjGTq7
zjpYyn77oStOGAlKo/xP0KBuHz0RKULUG9mD14wquD+b/j17ofjRRAHeSIV+90L1Q9PNKN6rekp7
teOcA4qRhA3SxJYw91c0YvJiPRK2FFN3315DxMEqPCLodTj/TDjaSxdh7IULIOUZ+eleTQme6bfD
XpZSkpl2bKPZG2Iza1kG4XY5VJzBfP5sNHyG/PGBXoVjvDlesL3cPQeflv7e0wr/k8nulJZ2wJHc
qO3qQZFkmfl9k3KADBMuqpwVZicvuqBThI0l3cIgSBb4BXgoOgHnUOiSgB5FVViXs9cYeJSUxz3X
Q0FKo+mlqMTCcffSubuqSOS7FR0iFdWuUyUSrb514kRddXzAfabnoyNcNJtrc+AKeVBxqfgpRqQs
lgwRumgJdeeV/dDHvOgqwVxE3tv7da1bSw7Jjoxwg+QP1TyJEkrINIbBh6zm8y7052u0JmUZvTeZ
w3qEv156ocf6wglAv5HB4OtasC1V4wJefITduKbkQcWcIX7Uq8PbRz30fDdsXfq0hkI2sKWgHhO4
ZpUDDawEBtf9R4w41tUNCCUvBOvrgvIppwXGPkLdXzmNDi03+x32j1gAbl7qFNvKffsmS8zcKlNr
J2kKjAo0VxCHnkFg3kXmQSmkxZ7zaQOKb70IJugnJRTaY8rkLdaUuXuR/MRbOVNGk8v7xWI9TbTY
5Py3luOWMnm0ahzMVgZBDMLs//kohmTe3jkiS+v7a3k5URSe6a3aC/toWqCD2gom8GihHrSm+wfe
tdXfSQhHNEHKBHUIBRlj8mmTS5jlv7TeCMv2yhqYNfq0kJvYfpSWrtkogvohVIx+Na/AAkNug456
Jy3mXAzk61PZAkHTERDbyh/Yfe0Hsgen3zxTv0+NFj8BPPl0d891Yb6ZljChIUU3cg2qZfzhbMbC
w1ek4dcBsiTgqPrha0QQDNnh9S7OW4iQ938Gj7qHjEDuEKjXxNFiB2ZEkpVx3xXsfPIdKYHkNXKn
2qyD55W2vWXzKoKfq977TY6ExHNHWSSPfApYFAO76yTZv40WhX9g0qkFLlTvZsJGpd7j4Wj2lUrX
lxGNsQJhyrd8QckyMgxK6mT3AgIRBlvk1/+en28yV8DKw5KTs3ngDD7eErAGfS9/ODr+H/jMBkXS
NTs+JQwjU2mokmdwGSoIKy0JCh0Qp6cPeSRulSDhhczQAyvXD30+HzqPbiMzjGOA62U4HvOjWU4t
6ICWnVY0AI5WwW+v1aW0hb0RQ4RLfGO+QSLmZuxAamyHdjtDRljYgrNaTUo5ba2lvl9dtsfqFM7X
z1B/LFaiEEKpOhTyqv7gB8Cx8P3/IN/FDBXYuyPGuhOSKFbRi70+wSyDX7vhcXksS0bgRjGSnJOw
GOKrX13FVFZ3YMG1wCBq7NwOrjiAYUyMcbB0ZJQ4ao4QdbKQUmH18MXlnbKw3zZ9gq1ehIvtZRPx
+Q06Ox2TXMxQfjr0UJKyUZ8wwc3emBs3yKnlMgi8X98FOCprCq+bA2jPFiSQNwLb+nUGZbL4vVXJ
iI92mxHO8Ajy02grlgujsrwGHXB+0dDixIknAfiRukfqS7Y97hdikRUxolS18CFTvDhyAyHSyZwZ
f0qobm0iRIKgQ1d5a2Y5IoqcIIFvfZaiUTGILKo/tpYrejyRHSvS1FZLqAcRojuwzY9tvczpf4id
2/Lk9nUE846UWPm2ga9WtMc4WNVypa1ReU4pA99mFgH95WnaOvyFAVj0wR4kQar8t9l9umGzYin1
06u7ePKC12zPvmTOwpBgsFc38CDhtifxuHeK71ilT0kG12QmCH5AGQc3uC+7MAiHEgUNB94Kok0N
OzDLrLlQBKfaRQRqbMLKHr/iwTm+p/v272uhcuOEmEdA/fTQb/+ICBZDUBsrRD3KdxTsfoYjgY30
bDgu+3RdusHq+7QSWJXVAeyAeCD/No8eyj6YAb+N6lApCN2xKEEndxnYPxffLcIly3FBu76WUD9F
Qb3/F+3p1Ur5NKvzPNp+Inzz0RBQJKbO/8iTDb7e/TS8+yuzoMoRwUvvmHau0aI77ei380LPtG3B
ZHF+vI4YukxcMbQoVqxFyNLXJyA6C1jul2gRPue6S2ANPOdiv39Jbn3IDdBa4J1YJzZO7j4GExi2
sDe1DZyMOoxsrepKBFBfAoxcKUcyfYIod/198Zued16rL6RPF9Cu7XAjtVFvm7zFRQOkfQzPXue5
XlOg4suEfz+ZDGm19kACjq/ugzzh5iS6Kp1KxmXrpstsCLi/u5NoDvb7HNG4ohI+zLNJjBq20NKc
VRaxpPMvW6ES37om8L0YP/kyqQVdXsfhbZHdWfNOuvj08aXdv+kjEfGNLb0RVGDeZQAXTuBO/bVG
lVpix/2pfAPHKP7lyHVLnJuvKq1XCQNouQwVcsyr04KSG3CyKCm+YkBmIi1t1p8KKHr+5obZKNhr
asHPvOMvN2X0RIj3zn3lXxtgiYRoQdO+u/9sfNTFY22ndgzQEY1TthnrNY2JKlh4rwbN6biwfDld
FoS62C8JNOImg5Z7781kaTT3XeDRtVrLin1Av/uyIQntBSLTOU1FA/oFuzUGnfHkw/Tm77xRlRwt
elUSxAY9PhcBVva4Af9pBSJVCTaAcJQ0nfhU3QZyM8Et4vTNPWkASn262Ex4DToOVGEgUjBVSmk6
slKELvbO1EDAB7phJIR2yvWGOoecqAJKmI709RtPFIfgU4ZaL2I1ZryKofQPqDYrpeePFX/c86wZ
nD0a0iHXTJwNSpvkZvMYwYsByv0el/antmDxrAKnW+DUEDBR/NTbKxGTIZhkTXK2cm08RhkLXQQD
FKeRpR9FYeOhOavblHgxGD0cAeuMIiZI0wnPRClR7KddlHcpiXTSJdCZUeBZ5vzWqO1SqgIECYY7
1K2mKgh0vzNj16a6AOrfRAr2Twyx0ZxMIiIJqdzK/p7Zc/wb2fNTSfivp4rwbv8Z2fhPYlvEnsQf
Qt5zRMVJ1bAaOmr6bNE+1zQlO4+eTIYi/suRVdGcPV0GO6Ymq0LNsP3sGrRvIFtrg/+VLDBy0QZU
rHH+eW7hs31M9wl4l0mW6Pu7yiKjPSebyjhiaRrak2RCUnjboWcg59wxexp1nopA7YoB4RbXjdol
wXdUmNr5/AQqR3BpahnXo0t7e5JYBQuGrcdRXzuNZknHXa1Wdj8xayG3TvjuPk/fKpGHBQkLHMHE
2YQkXyBvU6+LaltWj9pYhWYPbqLzYsKt7V33j+QKwxdmi5f2pRSuYPbzwmbz0OFYelf1X4YRZswQ
QU7dae9ksgCogt9yvz1MxAmhTQt1MPFcwCo9o4KKEbHdMpBRUhCbet9M3uAs5DtIiX/4ZLf3SrmZ
u2uicrfVde0iF5l5uXVRX0/mfpg/1zgX79Aid98DYp4MmLuOvarXXAi9WW6MVMGG1A4Q33v3G8WP
lCAcNQTd3S6FnY2DbVmuodYH1cMF54YT9cyqM3RTcpFv9mUXmjjMEn+ZQpgKgsyrDN4uMylqNTBb
SU2mtNT50/qnVJV7q/C+VNkpTnSUnj3Ic/1QvBuVMn/rZHLMWFmEWs7wnVhEfnNct2bO/nGj3g3B
984ugeMfukOVRQALKgQMDf2ctGNWwwOfJbrAbAQcQaXin/zJ6hV/MWCBxqX0OFB2Pk1TF53Thh4Z
686uHfxeZuldIlsIyn+J6YkeytQC56fWF5sJoO1gAAf7hHmcTJ8WoXa472VF6Bxalj9wKbA5rELc
CplFk0sHxlyp4yZEHShMR73OoTnEM0fqe+H3qE3kEZastGrZVhXuIbyu6ELb0q35KvY/tFNlO8OP
DO/riHlFe33AO1C+xsSCAqGUR2QSTabJ5IDF56sdhidiVhxlT+b3Fq61NXfrZxdJw7j38wp+M5JD
uojUu3iRtW6sdvPkvySxQ6AgXWOtfQcoLXcVO5Ed0MT1k5JwZualAoAgXOlPsSyQn1gRzILVqRDs
BkEBu854KoOW3z/kgHZhxwMedR/JUZ5WpFzFsYwH1L/ViATEAv/t6hUZJoYNlEOxFazVxVQmqkux
bMYfRVrimHipIU/Se0OvZeVi1VHVrTvLRpAAtwzN0Nowhf0UsKJbHT74dLyskNEvf0EJoxiojNUx
MfLg4Sev41qHhR9NhiXYp0hRUW111lq7NtODCBjAdDGWltVv7WIw9TKxiUZ2WbLWKhRPA6J+QzkS
Uv/uXPjEG4C6ZjwIOpt6csAO2nQgEsQO0iWiBVWozsnOVyxTZLhCjg0ZlLIOi3wODolbhA6r9JRU
v3ShMFFLmm3n+1GP6PG9emlfGxPxOkG8God7bIu8BY4WbogtAmEJdNQ0u4ZTSuvxEA6gu7qwhtDA
GdHPIg6yL2TE84ycHHsyum5YBUT8xrhJLipvds2gW0QMgiPUdVSzEAHkfOLTRmV4nwUdPM5Cya24
yGouEmXcYhgqbfIVQq8WF4gl0r4xWmUdxSNz45MBj9SQWpkqmivRT9eXnnSfxBzrHAzQyruynIuZ
NFaBflejrEC1mRjfqTEHH9TWYAM1bndMHFiUJqlieDC2vF03O5L89hZHFbwtxl9M6bSKF9zBEXJ8
HYXsZ7+9+6jAKJcj6bHK5Jowhg3YzVsfbmnWDUVlRlJsaFiTj1d/tyAzcxVsagF1TbilhRNhQmOw
kX0cUxDp10gVFuAqG7W4Sm9h3OMM59IEnlhqQu0JrMyT3zK2bFsXiyJBieUC0wlcX4sicfBghsvb
NkrIwDvUAubhJNCUklsI1k6iO3wHcRmALyuyYKwiZrqvNWaU6/KNyx7a+4ozLohf/YnmBqAs6KMS
BFoFWvosrVHJXYCPEsBbw3ZjJbjRReNnDXQMRikZ5UcU2otkq7r5gCNJ/MCeSjJL19cdxKtququd
S3x3M1JZB14SumFQwg3R2SXbSeaOyTfE/WVlqj5dEZgNSlZ476sFxYalKY0UEAXa59ErmlbD9Ct5
Awqvbef/78yh0TF4nLM2eCFjq8MRvW+JR5BTw2GankhCRxjTV+Lhp7lYHiPkDZwd/vL73TzXsp2+
4zUTZ6EQEl/NWsJJcmRZoDnhckCLHFEUcIkBZ9wD7tLvz7PpY5dV85eNvXht52rBlsHNZ3DTVam0
sAzQQqsS40x2V43w8ZEEXYDQ30n+cSarYM8n4nkJppqS74QfvkiFGOvjNSSeZqQmSvt+L7V50JAl
MEhN2osrwVPJOKNkT4lqvEIbKdgT5itGsYG4w0jLfh6zrVhrrbsWs5E8aS2j7DZoz4OQ9XXSkSX1
fcRod5ONoloBEhAq3KGgWm9ONzbxhBHsch73KMaGXqvrSJMSUOxyWLnxhMTPTxst6q2QAhXKwDlv
2j9sw6S6yyJ1YKJrSguAfHMLvPA1dWYYl5x/F5kVJ9xEa6VirmjHepbPdXXTSUcLT9sBmmNJ34Q0
1sS1zkQ2nAdp9z1gMpzFvgkaKYQLixmyaBrAS7yC2mQBCECc4L8U2JP9h/7ccj9trcggasdgsLSA
G8c5AC3EDe/psMB5RU1Vv6OwTokgppgxApAqHRfRJouyGsObsO2Ye1dHKwJ1XaSBqJBF026znjKl
ijuBc8pbjUAFpE36nih/ITUGFWJ1dPzSbOy7xZ8yEvQOH778x+kvTCI07fVK7SM6dxxXuSbUyp0g
8P3h2WmovxTIU2O9Ky8IFBxuQ8wiANdG7qrEy/RqX5oA8ozHtX3DALYmu7po6qPowKnl9KtHrRST
h8AIS+jDSOpJ1MCoTBqpvJmsHkogG+nIhx0g/fdtAvlnvGVKmmNSZPKj52FCxatyHXiTHXVKJ2nt
5nbylX6z+Vqxr5RY+VFj21+AgXeiNkiyidaUxrnyQkwDcrLmU7V0cWTvx/qkljKPhs22d2Gx7xRU
hTz1UrICXDrXXX3PZCroGDIgDPUW9LDIuQYRDAID1bVJrhj34Yy5i9+RzIV7/YlpdBr2BNlaWYF+
Kx/gf0ufQjFI1UE2e6h7K7O5SuAsoesEcGsiknwHMFWcq+p98iMBDYlOzHPWOlFGnajjoanKyETi
UNKuAT+LjFLkyQTl9lKWxyKMgJa70VDDvSVrhUNakFTBIl+jgbVu4l62TWVBLlLOEIAOMKaWbFCJ
Dp3upScz5qE+h8p7OGDY2Ln/53B1QZJSlhPq5TN7qDUnlCP2ecIodkMWU2Yo666Kjzjeltyr1aEh
LRjzbzwSWlNpdpQ3N8ghDIbtMGozxKa1WCWz2xEb9tpeQ9PubqU7AtrBlkyY0BuItCZhQdHAD04p
6N9qCXRBNrtXE3PSpIc5V0vROCo9ZcmbRpHg0EX0PDJscQ9wUFPnMlynhZKxAKrEHtUBDsNa/VDG
y0AIaSr5XQVF2lXf9c44X9athTyMuEB+H1S2m09gjJIbmgQVy0AfkZaWWeefSCrljwQSOk35CLG5
2JTMY5srVNrx/l8WMrUsgHA+eJ5DYhp8RDoNK2OLkXTBRK0HC7Sem+MKu6VUBvl7Cx7sKmvOwcxY
VnrUiQqoFoljsVWvbmju5Sf9ich5cYG/fVpGgzWwCnmx4LkoPPcz+UKMuZdC6oqhFNtilvkHW5eo
8GqgVe6LqDIEk5rxMau9oNd8YvxjiUDlKPaH3B14g/y9dCFq5wLf56QYFI0N5RM1DgGV3N+1qFQO
Rh6kyVU1YVrrJ6qMWqCTas80+YvG8hi4Q5pwGNMu8PPEjLXZkoEPU6Pwze9cibLNF4csh0JWU2M8
lRlYJ+BIIKGlcWFPd650Ytuw+GOmMfSvPaCI1nmkuIHsjchK8DMEB8/XQt6M7t93kXa4m1FIfgGn
nJaMQoH5s5g+p5OH/CL4GUhjT3/FA0mVj1ZyqDJhjN9tmYvKOh0FV8CWkS9zg8cecZci9MT8d+K4
83xa3IrVcWgPZDKZPzmm1SZ+iR7r1/1qWLlwQ/7wNISPk78uJznrZ1WS0oz9Zg==
`protect end_protected
