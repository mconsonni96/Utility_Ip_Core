`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
mshY2eieYaWuiesW+im1bu54eUJ6jMfynVhiLateu8Fg4e6zPzDyUlT4BjQMvPcQW2lJyckfEdnF
hB9K2w2AH6fm+cU4cBCfuiB0pCzNnE/H0QxxPZZ441fm/8wxf+SQOWaj8CVm6IkDJm4gjftYmUMz
Z2HY54ecnmLR0/Czwxsdf6iIlGn15AWqLDr7UKnHUt80P4okgmOC9+kI1esc4IT22CZPlFNjk3Lu
Ja5o0SQOsu59DDmjjYwHa/hI+wsXeP83wi7cK8Txi/qu+wC5MTXjhN2lVbjXcC04zEyBp4ItnWx5
QVPixaR3qnQrTdjGM5HX8pATAh5Y6eUOzFfL4g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="9aQcpHWvTVU8qSZsfz4fMCg8qDrnuyI18ArpPIY70sg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16912)
`protect data_block
BcA99RvGqNbDuVGfq12KZnyvPX700EwPTXAzRpvjtGQG1wMeoKHl4NkKWPgJT6ZQxTiiTJEgy9d8
8I8xdfzYGGx3JVK89j/C9nkXnlb6LbEmyyfHHPr5ZSDNAup0g3xZ6rMPYcny2CIQX71tEwCJD56z
gseuw8E/Uv0wlt2nWeXXVcrrIqaRyWHhW710yTlKJ1zrhHR7eWlvSo5/+46GqqPbtQ5y6UZnVuWB
HenIwNkyUXw/aW3afkAPWfNFWcrYZ8IcWQDclETVM0jKFyuU28J+GJHOcCgsLgyvuG8Z1neyjLL1
mAyjUqwziC/NbUpXilMp/LbsB7W0J7rB1CGIN3AKN0c5UOznk+Kk+d/IaT0Gg7qA3XdJ9KNZLOKU
AAc2DpPuA6ZmFPBDXXW7k3pM6V5uh4qCLSbJRYlrHJUF9H2VKHSNWxyw9rCOgG4nmH3w+jsFq9Dx
KqFA/znudEHw9Cq1EpA2P4/ENmeq7Yhm8oAq75yRwPenrsEtmWlvTafGzLse2hr2VK/dBirgzSji
wLuDbrFGjjlTB7smdwslsLQipbQFNsRBbDT0C54bj0GXVuRyF+3wfDT018Cs2rsBJN+EiEjHaYLV
fJ46lPr02Si+xX3PpV/S/Bhe4UL0R7EMfqIDkQqDIjNvwJwxSV8lTgJU04rc4YEB997Cdvznk6H3
4KA+JJd/6pPFVTiEkSYtfRdDHVu2mTXTHsq5yZbp6mHSMIZ80VYfdSvCjktZpsbBFoKNodD2xpYg
XTCMeKXedZVHvQrV+NYdpHEBcV2JsnWCjjUKJQ2jp8RqU67EkFIDkh2lkWgCnOa/ePSjhiRMEFxD
RWlM9n11e2OI/Zh6adCTLtUjH5DW2yWloczyccpcxp+yknl4G1w8KEodwxliVhAgDJkUiuiuespa
a9oIjws/gTdEZ7f/KCxj9u497nb84f0QmuFeV1MiRGw+6QW7VA+jv9iiPU93QckhBBy5hAgbkgjK
AWd3TYPCH0rqdo1m6NNKKzQvOkOdVR5sqtU53Oas4w7Rfhdrgc4wT2IfFAeflFO4aiXVQ3dTQnQn
kvvAtzgLweDEHOmMtZfaUwtdzxRmqLuARPFtI3JQwG6jTjs2MeziCPvVS2ABXnkK0Xgnyk47BaSr
yxfRiGvdPgsLWtxqE/P/QPqHYC4zZyqyotv8nyePRzBYEr5WdeKd+L1LAHhO9Z15x6U9idop4c5k
OyreQJfytuyWh3Wrpi33FFgs9XgGDJoKVY9UkgZLWkB1+RZW4q4NRjOdokSQz/AFk1vr6t0vqygq
QVr6Mc21pDbBS83AvsUbqtdu2BZHIESCEoH3yJoi2Rexa9W3pNtCg+p72RGWQ+jynU2CYBbf9erZ
BDCnbPeDTjK9iA5JQct3o4XoCuTsgsq/jKLz5EkadP7+sU1Si1bIG8YkAsjlpU8RGVpKY/iVU8HZ
cQsuhAufo+U+m5jqCUC2v6X/klXNoryAKP2/knkJr6ORiQ0ZflvZHGkYurydZ4UFq0dIigdkfpIw
Kr5K/9K+VGxC5ozXON4xE4PR0d6xqkSLk5hRzM81gR75+kMe2yttXFG4LANbXjOzHa3T43MmIS0h
OT39iii0CXuAxXJuGda3p9alB6nbDKN0Ps42EUyeX7Bty+c02aLR6FxXMrPpqrFLAnp3EIuUJZV1
PHTs/8Grdt/8Oxy189im5io1XqJgYNIlAku5L0TTgZNOosNAESABATWZk3438RU6/FLs7HETHLf6
XCFnT+oeixroVjzcRNTiSU+3J8vFjcsMTJhdv+r0AuvHRST/uyw1o26M6n4lw+VEwRdvfqj5XP1P
gCaFdC2Wq6mNQFHi/VpQIwSqV3YpY6mn5MhH8VA7CfDcpEWfAOIlDYp/9RUBaZmOd6lceNOxMq8T
6sVkgQsLEtcrKZawSsa0U2gVE30HjD9x8HYcLgdQFeXjN6iBPVaLhGQwtbi+m+el2bOR8eBrtAkh
pD1Ej2T5P81OUGIVqK689YK4+3pFPrwooVLSrp8GwF6BeLRw03Y8E5Kp+roC4V22r4X4GwK+WFfw
7ZMtpJ22FmrLiDxE0M6i3uS86Vdt11plIXcalBPJDWDs6bnJdjAKc+MSM0SrLNXz18nuKQDn6Gto
bDIX5CgBC25/Ers4D2UBFoJ4/OvpY5lfBzLbmLs1AFtT0lWZTF8Lq/bgEhpAkO15p8oW1S9baJUD
EKQ+E49QnB0hoExSxzoRcuHbUDUbK1HHR9cvaindiCS2v+OuImQSqjnFAJzMoCLz+/7YsGvwkwdu
i7Ryuwj/fL4A+B/sfmQh2KJZXJTj/TI7FOJ7dpNJpDEhCRPL7OtaPtBv1pyfwhIOvG39ObG/vuEY
R9UUPkt7N2vo+g1EanX7UZDWyKH9oSqW+mvZ8p+jalKIRfdSxEszxBhvuUVtCxivIJZT7QxbvO1+
y5WS1gkfVYlVjEPeI6m7kwHIzpCSAahDNBrMBYGl1spud8JH9p4HxBaj6ohyrVxaE6KxRiArlUNT
W8RJ/L5BImraKne7zjmJnU04tV7DEIOGrFjcNnoGITiW+2BCiabKYC+6BM9tDBziJVinmQDZlbct
djtIcasNpPfxH135eE/KkUK3wqs1s3t3R0JJurFDVVa9rDrMDnzaf6Jym8eEsAmmiQiedw+vEwud
xDr1YVq9fb2Jokdp577ogmY6HEgng/y2a8+BvQwJ+pnucsbbLc2WjRJhLEvSxw/mnlMt72ZAktGW
tSis+zJc2m3VxOyF4dT2lpab4srAgDjMnBqie2nzt4IrOuA748hwxFv8FA0GQhOLzFJWgbztywfK
SI3yd4AHFSEhj3/FvcHUhsxipXmkQ7ONtuHJgA6v46N4RL9HL+v/1pC4ohewQFVvG2/boen8tsd1
+3D3NvFHW+cykeYUrzKgz0nFjeezNvDIQcCsQmKjNDgMVXWz4A/QbS119I8wUJAngj68Utogf26f
RxyA0ZxcjpEhFh58i88b9GrrIw5TcB4Gj9rpNnnFJ2OJ+IzstSr2ZmEi5zA0t0SNjymIh+dOfwM1
yCcFg6pvFrguiOLK0IsVuZP2Gxd9ZHCVHJGm+jkmK71rBQdarte8fDQv6cpiK5CQEOesQAnOgLps
pysEGRCenWE23zx+h2B1tKpbo0cdGuZ6SNkluQSLf2SzAAjnir5uvHqjl9pGK9BajnvEB3L1+biK
P5iLPzD2ozopfER78cRB//jUOMIvTa1HIFKGDNJLC3qxShW7bSW98KC3rXO9n21ualBcCz30+MCr
c2wMEQ5/tenhLOBqJuyIQ17vq9lIFq4OSiM/vWZHcS+vhAYr0/aoceOJ8vRt5HEAnmrMBdlDDKRt
F+5wWtlAjICyJ4twyasFMNXGMbuf8G/GSwpp8cxEcvC7bMX9qzHkOXsx478vwxPUPM6hIGgKTfOD
HK/kEF3JHRMbzf1hxSb9Q41RnpSUOf9k6NF5/ZZufNmKcCOzEPRvHlkq2yd7I/HO7xTeU+V7Apk9
+Tbv75VBx0QbtAd18J6TA13HAwpTyWErlqj2UHRzuNEEZB6L7obuT1kFIM3CmgQjNGZ2aMjCPSFE
D9tmec+RbEMIdEyx0EtmPEM0x6IbIYbKFzxa2hXa2zjZX+DFje0uRYIfH7s3ibyytuYKgrXOFZYU
AeiMFYNd1OK3OJ1JjdXRkSO64PPiLntDIuYLDl1fEMXkBbMtLTWIehRgnNOo36bxare0+vZRv82S
EVzp15aoYkdCNj3m86n58AxDC4A7k/l/PHqR6la8JuV/NYEeEwc6jt9me8vSforB69CfsZzQ2rVK
tGMzOzqVxHlukTn9dxp6NVimoWGDIXKp8+n3ymAV86fOkhT059y9FCslKS4rvraLuLmc5MAC63Zf
+KW0G7P65eU0r7+7wm+CW04lR3z6n0tgsStWjIlJEo6hsgEFi9I9kuGbgV2giBOVKwODWzqUZqjc
iXbZerHusC7PYhxDm5Wl5NwBW28s72/lj4NfJ/NJ9AToAWEXyh2mKgAUdOAzBzv9okn+oUxiW93k
0mQSsFyYBjy7w97lM9wBf5ZPIAOeJ5d625fTUUmW+CDagB96Zk5cLBe5WKIiSlHW5JqBegvnem9l
3F/GLjARZNkuY3oJQsJahz8O7jHsCYgVum49whHKB5B/VRvIQz346lBd+0vGxAYkHZCHRzr5CAvJ
wPi49lZBIpY+eDsCdi4GR5vNDkqhRpndficbxwyKAan3CeSnz+ZCpV9DeFCxDSC04Hyr2dinTxlz
C+XDADLFALZRLr4M/ZdtyaH6buUuhKcA81G64RHgXiybW9CrvG0KLI32BMZLmw799u342dQdWykS
db7/xEx/U4Zu8k5E1WSEIy/k7JYfewuxXgV6tK8nIEOJaBJ7oe5RYJJYv9CdPFOge+BFgmTi+5sR
IKH67Nd7SpvUFThwA4/HbQoNhiqI8Ugf/f/16ZuZrvPUo2FnHX3bDTkru00/MpvNkLssULScG4K+
KlxsdKXPMKPrb13jvDivwRP72Q7sfJcabif3CxoNwXt0KOVfQodzGWgti/5qMYaBolfl5jWiiZW2
glyAoFiSVzKGchzuDL0AyMmZ+FqnT4/T/s+kke5PuBUVgRw3EsifhGhgV3GWBPj767UdMMfaD0SW
ADaBgDWRyTtRDTsZs4cdVejoJBmbRQuoOJF0GvW8VkvqPMIKh7dXv/2G3VBhl2TKxEsuMNEQwmzH
i3nqU5MlzqwroKZ2zlf6SB6drtN3i2v3zC88FH97J1yd5+mbM8DclH3s+RW1VWaz998WUla31iPT
DdfXNonZChkJnV6JFsq5/8Bav/lPrVJy40+Jk6a+qGyHBKhn4ZOBGCuoomAta9QjcgVyp8g4lhLy
1DcpKoDasP+rPNKNfMFiDKnK8ShugsKjk49AvQ2cx6Gh7oI6geScCVu6udntg9PcKptDOP9IBwFi
llRjirrAhquTYjXl0ehw7hJfYwS5DvNv8UJwsdA+qIHvRs9/QD36+VQHIDgBmZsX3/oZX5zGL0H4
n1BHkqWoTRRBBKbZ3I5RoxU4odyxkpcyIE1g8uImXd/59M/hbSL0ZZCDFmUcTDJv0CcAsjByv5yd
/tFQoaA3QpbNRu+TnnRWDkceTtErh3QBuaTyAWGxG2GBq0n8lF3cmaGKgQHiQJATSd/Bs/nR1obX
15RWYBhcTLfrDJlMCp1O4vvykFX438lf/mY2LIuhBujVw5V80ahYXyAZRhOmjXC4fwhOh7jQR8aN
HeVEPiQhc6yGkJlasjKrvYonX4w7rH1RU1kNEJmQWi1lTLI4ANaG4CmrKIFBK4uA5jm1lFV27nNG
CPnWEjfIJz5dSSx0BUCDXk+u4it6EveVkNXuE+75iPgSsOfC045JIVNsnWHCdcndNX9tEr4kcWVb
1OAMZWrVLchV8vygqz7lX94G0jdTaE8gDQJFIsLZaNY3kMR4VfWC5LzULXU1kMe8/k/Hb8T2cF6q
9BYAPxDGa0Z0iY0y6gKlFORVP5ypTdPfjcquAJskgGyLbrorFy/7W4lJt8ujxyJne5uK8RxvhfG8
dKX013vCNi0TE1yT8dr2EwxdHANC3IQlLzyRGXUXXZju1YuStXJrou3F+8fRAm3zBce5S5jkj57B
hvObTvPWzRCmGjpbOv6KmKJJwICq3wcNvEs/NEv5Hqu16sRlIBOr9fpufvDedPQU3tUoyFIEspNM
GQrzNMMpjcfquSEOXK7YEFGXPFJdc3sjfUgNDd1MJO+CROT0GndkLaTiAoN+QY1+nxz/R1hnn1zd
J+vkJsb+nZOXcvsUErKQ0J+AZv9kV5NeK/JdkwY/1e4sUMeUqhcsllSOswjoTB7ZKjSOUDYNbpcE
BIdEvRTdSOk0uda+mrakYQNJ1x/TNbvfw3QBqocO1/aJOXh93DzUEyAPjFxxohEGQs8yCHtH8agf
UUicC/nRWIKLH1n7R/9fWlINdEimuRzE32cRbFfRjGgZHne4pm+l/8P8vvemAiDnmHpSyzCDekd7
ei24dUo0ImLmnTnWQYtVLH3Nx7kwOlRfKrE/LXX5y8hQzz23nwWki/JUTMqx6g1nmtKb5mmHeuN/
EXyNx/1OwlMYZZqj8BNNFgotzVKbmALXY4hUWXZW0xCSH6oIfZ6GNXTqZXaw4QMO9s8gtVM+zWdf
xTlfqwfqOpLB6SI5kUIo2CiAk863sjguHFr5LRaCrvmTRkkUa0AjNQMD3UVr+w+fvl7KvA/VZ9RR
rj4iu2aSfqCCGqngqKYro6/3a3/S1mAIpBH0m29QWoOhGYe4PiYHqp5HUIySxO4vg2cWUiHoHyaI
ava4ZoU3lqly7rb6TjViGipFV9VE1YEgKtAShDvcBS9Cat9U5SGtbBjDrNH1e2uyBTZ+hdV164g6
biTUrigZ9Ay6WVNhy/73OFCYX8zMvYmmCciO/tQaA+ynjnuHyVPele5JH0VM4eBiol9KBrVPM9/z
hmzlXBKqr2GdPkUMzUqHLY2VOegClBGSoCheB9LNYxoqtwn1Ex8pi2S/xh8Dz/GVlEx2WfZYRyjt
edvRI1rLMTucw68V3IF2VLg6rqpcIgoeCf5UAA/Rz0rnN0rUEqLpWPnnhuKa47KIIHQLZ5kklgd7
2XKJn65n7XoqgGIjwZaM5tVLb6mS2zaaNupn4M8Np/8mqqLnIu8vjHGHy+DQF3tFA/XBxYivtACx
g81I3SnLi/6lXsETqxAK3/b6xwbB/YYVT6CdQ8cW3HEdWHlZh9TVBYYgCPExRtASw+sXttmh5tN0
8sYU1JiBMLO9r5Gl3F2x6IdlkJrJ56NeKIIsoaEurdaoZxcBDuBMhntx+H6okdacs5Nfc+nNqWJi
gxHUa+ixq+mpWoPWa/kj9orhtAGEnh+sDc6jzr0o9ELlBM74UGRwZ7mNQdiQqGfpAKjBzSFHoyR1
KqYIWJv8XBteqM1izFa3NL4U0RtApCrCeDH7XeTGyo4399oSMi+gTD/YEOpSCbkqFhTTqrnpTBSF
cNhI0fy7Ci2uYwUQ4imbhiLymnu8jHidAX4tZybBkUSPNej4P7sgOJNQOjVysksusoGZs6Lta68w
gCmlN+N4HzeyDTu+AHg6lAix/6sL6ORNIt36zs6U7BarBXqnDzUG9DgdAVoOmI7cln/Ox/bPqZXx
WCBO5HSevCdpV6vcH/ZB6qlm13Yd5bZHM+lFNfGmgNwFAmSsjJ1mBBqFi6GWU61MI+YR34st3AKM
YLwEGuRuuUpngqzrHNl5VElBEgAKP91dBtFwDAaZU4LL8W2SWlGJLgxCyyDnZmDG9oKAIloBgyOM
804zvuxZgu+/4YrFIFqPihONAY52UstwOaf775H4t/ZVcJigPGUOaS3um4Ge09hE4Todc1Qtw4Bm
7AS5wgJw02REovPf4OoSeZYqgG4IClAbe0ie0dFBgCxjtq8+ymWoiwsYP55NJfN40xAZCXb8B2i9
+s+vsMfckM0Av2yO2s7So3f4MLpefhHoQz/spVrjppBIDP59L8kwJpDRzF1cHVTzxcULLdWaM5TK
GchybNQluq+E2H4wEFdw1P2yl3ARGoZII8qZs7PACHmCpmhi/IOSH70qyuVMurS0CdwV2YviBo8H
bi6pCdzrlWqzJJ6gbwxUslcNfUa6iSUXUV1RHyQUIIGhd/l2T/Fns/YReEBFkJZhOuqGFMQtKmZh
pXBV4qEIBDZDZgvr7XdrpAWaS5Tqs57cl+7Te8L2ujH9Nrwn//Bz6DOMBR6YP4LV7UT2z1rb9ysh
Woc9+z3Ztf6Lf5eD012YA5RnuVhz8PqF5nODLDoMOpJUN1fZv3zHBCnNnBiacAM6p3u+TukAqbTe
kGYaO8SP5g3u6urCX9suzGf1U11cTQeu8zslVg69uCTc28lIh6Hum9mQ854xxSD3ULioV4cdVYRE
J6VQ01RISPQG6kJPcs1CUH9oc5nZU7hHIbnBwzP6ycF/SedmVUKQe+6/1H0AQdXpKvXCSU4QOBLm
bt6Wj7yx9VWQqxI/EBINgfXJ26GWNuAovjroOB3QdXKjlxYAf2w06oqv0lk+e/xkKre2m4dO8O2f
/mjLUSUd29WnjVzDgT1AhcMEoiUfrwzl09iwPCvoNSJtLfTvctM+f25AovQNbh3Yt99PS2Dm+ePF
cmbbKk/1S5q21Z4iFk6OHFraeEvHOvVy2vUBdD6azd2jnsRRwVh/rv6tB78dh/0p2lLuXkLKbFxK
DIevuSCFJw5pYNdq/iIHzt50Ow15bYVK77Xt9etQl8xIzLYi+P8mKm7c3+/sAQ4nxdu9LumdE7iA
+cQngpO8Zy88XUW6XLGRM8wp1p5VYZo55XMOcAaUXqyK5ZAOvdAiGvSzMslFsjFu9JFfoEKYN55W
VHXz6w5k2Ky/s8Bkd/CkDFNYtpXP8reFjOM3bKeY+X7/FXcJXJyp3SMCfuVoN2Ab//EYVPtWhH12
8U1wrqRCXh7YhtMVuMI2ihzayB0GCXRH4nJhIsMiRgPrW9t0PYC2V279IjB9fBnlsMn1Hqp6dXZy
2AgqANJTGeSkDe72ak56cUkOB7RSaG6aFoD7cX6vdwybm7SggefmwXSIjlk9uszq468cJl77hTgI
HYBTDVvVpASaj7jlYqfoJDYa4utN7ccoVC1K5EkQ7jTdSRZYkn7dq3KZTebD7KZzu3xddfMYv/TU
YHagZQY/ZbaZSi2lj3OPxmvno7Dhp/sAXEovnfNN4HeYJ1gMJlrH+o0Gwj2b569lWPBX32cgGUYd
gA1gFmoRBXh29gwjA6W/zND++qLicCkGEAtobcHo8yjd6qcyPAjAho6MwpHIhZ7lotDSC/5W+EgP
W/2cEFGElwZVOg21HUC9f1MN7b8RrLeABocxE0N/ZqYc4tfZbtK8Gm/WqvCqBpx5CWV8VADUBt6x
oXatM3gVrMA3iV1lYcfyQK4BeSwQYRZ3w9SfrDZTw0obpcjn1xMDah/XjqQ1ieZ1Earc4/voWbp9
d0pmp83WKevDTC/Wz35HwIjHUookx+DX+aOhlH+CbR3M+gL3PF0C1f22IyLdDHX8HFwBRFP+JlBz
BuESwFFR9vm+xYZ2kE78Lfvd8i7rUCgUFQcImAqeQTmA2c9EoF+248+TFjOkLGpedyqBUVGAqZiL
UL3U+G5uWoszbq32LnYRSEDCBkj9k/vFurR73gD0UoH54z6qXQP2nR/czIxkFT+GRSCE+o9T/NlG
hVNCbT92yH19TT/ebMuhVGexe+njS9mHIqnvbTCYUDozCtaY3Djagb1PP+IlltJpql7O52GZGtmy
k4sYgRw1cflpbzKQD+wg98gP/pq7/s7vLbH9n6QkvonYJqM4RLUSAiJWUFTLoSO+V068ei8/f6CG
1Uq5q0azSlyRk7P+HzDQxL+D1oTbWvYwi5kEWFQgZJo4o7WHUv6ylRXk3M8Ef3U76KtijheRoFch
7JyO8hGxDocDD7iAFKMragiWPMef0rQKr2G0hQW+4tH8Z9IyYUoR+rzm5+Cw0KrVPBcME7q5TtbW
2B6gjkgohFQsaoR6OODFeD2igL8m3yARQms4IA9pXQ3xSrCiLxPSxLX12jrwjHVc5Gmxgg+BYqzj
6+joFVJvf6bWJuRERAlUNl6zMBx642BR9l10NEdHCwpc84MClDyQZCfbgG1gii26ui2CEEzUHFWP
YR/sZU7OWLrCTPOXWANdrCQFo3RTAdqWD9HtpsPlT0aLzhi9aHYy2UawuygdPaN+1XeuQbbqz4zB
X9sZr1wT/Q8V1I44n3XsORHeRHUNX4S/vSqldWFeuYuHVigiG5uxNRBTtKxFN/lYny1r0baapCb1
7Hz5NIaS6hxZb6on5X766otoj7+C5Pzd5EZ3BPdorxqM3lE9Gp47PJ59rW9c66pBZytsNn8u7l6f
AeZa3nDHUZpXFZB3Lbn1jhI8Y4qy6Lg8TwFrGme/LOiZYIWqrgbO8JcI4vzsuKVo3cx8+IahRMMl
MqRBI8r7ZsCBwTDUjYugIS4neEY6+AgFAjwt++TZaZP4bekf73LdqjAG+aJeOGoJBIzQYAB9B6Q8
ntzYKOT2OUZC+Y60xxQi1aa4hlaKxuDI28f0LKICu7HUaMLZdPOhaucBVA+9P62PqyYzRLfjTreu
QSkkFKsLJq9yXK583TK5VxYT23ncfnJmXD7H4JBEfhin7FEg4a9lhXp+1SJM9NNneAMQQ337SRIl
i9uPKfzd9p5gCf+LbHw5EhgnopWvs2n+K+9ndXvqfdUCixosMrSpX2wF/GHQCZdKGkN4/ko6gp0o
xqzH4aoDR44pW0hdZEOQY62fV2+otSgDPvcJazK3CBzwISDTaIv+Xd/IKJJBdplUwud0gqh6SRd1
mS7AqDrbH5tIWXkynePAgURKkswCpWZAFHCIC9brV/XSb+OXuDgiuPFZu6IRusScW1zuvoYqUuto
HI3VJ1ioXdKtBP56A82LFhiume0jBfbLubhJYjXKZfp4UlSgSh+Xa4R2fVWJSTD/8kMrgV/FoUzO
SO1GSRDO0938Vic3LAR76jyRmZcaI84+5YH+HyDWnQOli5cHKOuXFtIYysSFk9qZ7VdQlL9GvdUC
i5U4sDin8nOuFOohjiOwcuB6ZK/kShRfc6SQJY2I5HNsbDnrqpFmIa3oGpBMX1BdAdGI7+vFTAAf
ZixFTNPsa6EOnJMJySbjpsRadw9MpuExBJIzVqEgxLBPJVi5MKvIU82QQO63M8+J7hKXbeDzrjTa
BkNPwK5yxTz3pr8rMbkRWVO0AibJNQ7bie/sofixUFhtwp1O5EHAj1Dc4LDB7dszw0NyOjuOFYh4
4ZK9XDH8F4jfBuv0B8VA562iJKkT1OJxp4iIaPbtUpYep2ALHecBqagX1G0jOErJI0uZPXfyOgEw
U0kyeyBeuWK0carL0Gb60pOQp6K83i9yfc7twOJ0KbuwGfEhO0cfB3qqPJFB7wkkzetAMqC6jGmb
9lF2KM3hOoxjDdWnXYdzkRbTAC9DFH18GkR1AsA2xgl68t+UfjAg/jXYIyybB3ZzvXpy0qhr5Yap
1z8sAC046Q7ugQz9qdyYkpyw0s5S1+ofdHlPjx+16ao9UPor86vagGPkORDXmwzyY6cKMd6QybdN
XBt8lbOE+xDF8HNmHaduxVdzcDqaxoNSmso6Dfw0/Ph4rmf7X/fP3FLQVVyZxehKrEqCDxoS98rl
gAbXa/dR2mYA1Rx/EU45JHVVDlqwXcgNE8omnHMyfty5E/UwK4LjG+4ekwH/OUsjxtbKvWNl65Pw
JFlOjq5S2p1ao46gd3x0W9P+fQZD157G57zq1Z5n/i7bG+rngpVIz2A5ti7U9ilmb0qdDuy35jFh
M2QMCBlFer9SKMbRp/e7jBtB39AHgWcvVsMfvUA9WdHmcr6hiJ8usrh00CWdkBIox7jKravfMyZf
LYilTh7KAlrwasogOJ47kbxBPeqZpL3CYwHpBrDF8WFXxdCO58uxwIwX84vBjuCKl/JGvQjpM9Qa
K2iqWT6+Tpluqhb2UsJHJLeG3Z9CueVORcwvz/cD9KdMP1ufSwyg9UlZulI5mvPYYbYdm64rrqpE
H67LG2w9v7QPz9sdsZQn3SStd5bIRaTAVlJlFSNNfUVgvDF8QXkuk/NJaAAyxTGZJ0CZnvjODPcp
4uqgbKG+QWuOv8O0Op/8ECO6GaAa43Zz8WgWJywBMYabQAMk5qwXs8zuQWdCOm0hbnNEKH69LYnP
i0lQ3H7yWEa6jiildhn0XNmT3LZ/WcZlgJsQwW7MrHvLeZZ1ugWFNmyMA1VlKeDZvZgU/1NsCyhy
6XMHWfgKi39wN3bWxBeil91q/4UUFi2phXDYWjOM87vrJqvyo1r+YRQa7urNHwIDvlELNVVmkOL8
Kg0xWdRWH5EuryfAHoj2Shy4SgdC8JrZPPkAIPmvbL99T/U9i5OnGy53Dq7MQBAlLi7i4hjyqxb7
1nm3gEAJyY7IRs7uh266qdV2smZbzVIaGuCl2tqIMXjUcAU2gIYj8hIZYPUYDj0g+O+817iO3EKT
pbVTIA0LNAUR980Rv/Id3lrCL30nNmNhpWQPX6wqn+zDRLnIXGC6hZDNXSNeq6FhHDnWq+ce2eL9
NpysQ5dHRHEwfeIMR/KXZ71kw8KOmUJrl3hEk3f90csQOCo1LtL12Tp8aasXdflo6LPQZMUaKAUr
P4lqDqgBUB2G9TPEL31smcV2h5sjhxA4eqfbT/KB263D8sVp7JMa8HoEftJ8SAuceqgjvf8Un/Tm
u7G1e6dnApDPkcu1X9f9kNG7dc41rlRbl5cHqVf3bVW8bts211FZNM0BE35PHqTXoTASEnJfC/NK
8C/4uAP/wBQ9pLyJHhl+2hyPTDQkdO4UtmNcWDWG0wvZGKgXuhMUpYltyGl3XR/mpyRGvj3bIjx9
mvpiLiZGbdPpqzh92s53PCFaH6MDToD4cWmmpuKqz4OuC3XyJq1wnzPXoj3x+rtSxI5C/xK14kWo
j1qxSrSnJzQJP+aZ7pyXbDLipg1A4u7S0lgXZY/3iXLZXD6Wak7Py9qNHojKyxj/EncwPheRlrZk
84pmkt+sKZGL0ZlZUlEs3IgKw1Pr2AcrvLBKBXOVL9FrFOmUsfCpruFIYFgE2hxiKcaSYTpiTg8d
g3NAD/LvM5Yx/mpJG8az1c5RnSiWeYVEhfjUYklIOdf7baOxaYW23JF/cMD/7hqw50A9/prcra77
3R69x5iFNo3Y8lDhiV8JajcR2fu/3EwffsCpopg/uiz6NxF5cMxdjdozMn795g8JkQZgcnE++WfU
AFdI39UHBzaECDEq56BwciPwMR9JoRju8GwEAdL8FZX6CCMKWuB8hcDKrkEgt5R1oCHfntF1EoEk
t3BWWKtaD3iHl5lQvq0t6DzAnBSLg0d4JHHpNcb1MHZJHBUSVQNnyLksvgmNL4paKUZK5hZo2o7W
bfalNk5/DlPKSGnUwAqO5WvkORRtnTQ4YKTiMdjtTHuN7uImYV2JUjpdbcvHOkiqgnQTbKBi0HR7
vx1pXfDURqHW1tST4N7rnRI88i9EVCsA9A63AgDV3esippnotWiLksLJqRbqsyf9OhMzh7QqXwHX
biwwZlzptLjAn0Qc963CmnKR/XW1rA/nFVgXwE3UudmcfHFCF0n45/jzrRtW5SgDya5Dz/1qnesJ
mi4tSOrPNLee6tXnjw6LOhfWt1G4Ld5gjN5IFoSdzbbUpcWKhxkdRLsFpvg8XdQYHo6DR7SjmXHq
r4jj8PKDhoSulo2XzhKr3biub24U1KBHirZRIqF53mf15jVE9N9hFc7KvEK0ve8EhlZmbogmW9ei
fvPCwIXlrlL6drL0+gFbV8ts37i+oGo0NTlBvkSrnGb8eb8VxSgPTxcM+gEoLA3U++JM15qnuJ7+
tvQ+jy0AlOOYy3Tj6gZF4GI7rTp6j1SWW7msKVo3B9lsNH7/hp4W1j9IiSMgkRNNZttNivNRoEta
q2BjwMWQgLAEoWtft5fjQCoAlhe3u6KQxiUF6BU00sYGREm+YSMZ3ScdWr9eo7eAHMPGQXF0BhVp
seynXwl89iVfeL4vWz0cDBlrtZw0H/QkvNRVmQMDUi0dK+ZvuOsHFOxAMzYQonVayR8F7AY53i7T
/jw1GR7cthFw04HR3caOl0mNIZnRUJVIq5GDCq4LTUruzDtHHoHhGN9DEQCAEE0XYEFqLEpOlcGa
QXnVjImGCgoAw1d3qDHCiSeoZKxcQ50FzbGHOqFqy9i/dLk30dVkPRjmC2u3dp3iNQHkRSAc2VxK
6jvp56U6bpQ6KybbF3PJJjaBdq3yFH9vTgNdeM6c7q/Vwzyl0AWJnnkVGIT+S6xScnRiChGL3Z4Q
nC4OPXNbWUXzELHEY3CATU4MWs3ExWlVvv0O5ai4mMWaWuPSrDsxAsk5I2/ErOY85TZ2s1Nj1rIM
f3fbYXR8BpupT4BIcRc3Ggb4eCMA1SLWvCdqb49KTcyTq5IFHT9IQ3ffHLqEz2h4PI16h/c2ajHm
xKP5erwFVgbHcXO9R2VKi5cBly81fVgF30kXGFRyHMF7XbWgZV2FjT89pOIeKLO/XU0stMWvopxX
F6UUWMhrKrPCsdEqA2vOd2qCiKBN77xOdK/4OsBlR1d3BKZXPSwBik7yuBHL7Ge0zXkgrqMlkeXJ
Fyp6tesrFjT14KXOs66IUkomjgzxa4JdBAM+e2rP0zPNzwHFty4dOovXXzlLIb3WwJEM5CE9jST8
4TdHYz/mVAP13kEREUU6TAeH0MosL03nzhRRYVvBInd48AFnXSqi5vB0rdZConsaoyop/MXM1YjL
AJPAHsiV7mVppWHZkmor8xYcg5ylWLNjdH37B9e0pO5f7vSrCxSZ+F3ASxChqhQrpK2GT/RAkojM
8g6MTVaxM15AatzdDBdKS4MY5bxIqbc5f8OmgtXS8FhoNLicV/P63pYdboLJQjoqrBeALe8OFsVS
CXyaPIWh7MnEsl6e4yWWqHn9hwkd+wN7IJwJcaVl19NENnlT1Inxjy1HjA1fJ7H67PNyKti+MjF3
eJM3cN7PdgeoMMI09qy1TTz0NG+ErbYPKWnJVwLA7U9Kb0feT2oLTzaMpvcohqGfNnAkcV+7d1MO
Y2rabJt9ZIeb9s3jPTp+ugrepUfiCBwdzICOmhX6eWeDSQzPJHaOkLeVljOf9q+6w7RxgaSyoK6s
KfVNB8N18SP5GMjHldwtLpYMqkE+xoVWg4ow1C25lgHLlBxr17q8s4VSZGXcM3cj+qMf+GLvZuB1
l1lb4M4g5RIWhiJ2hhbGxmqmIXHiuQwsSCFlgkHOraiN+p4hxf44cpez7kca1N/FcDBy//nuuk1k
dOSRo2HSbp+8W4WWI9zNv/XqeS2jePum9mmaOtzrL+PsbpSYZOJVlPEcxJuavMUhyn1d5VRGQb4X
0fDvN/PwioVOvW3DFACsxW/sxbKBFjce5jYX48t0vLdhTTPzp4wsNTC6OtbhK+rXLT2RJObX3M0P
lAi2zkbI1eEQZocoRwxSSbYb7GHIY8675yJ7JIEwst4p7hWKoMrbdRsCawXKJOsYTSuMFbgW1OFH
hLrnt3BgzuxW+hjbgD15HVwNUh54WqGoba4cN5Okrd21DcoJgEJmqz9KR5nJA9mVtPJZxqPiNqg1
iOS2hXQuDjQsDJa7M8LZM7HyUmQeRXONa8J2fMnK/1/E4318tkQnk6JH+Cylqh7tCWB0STQO3WtC
U4xQdTpXWwUFWooC2Cs1tlQuZd9IQSTANKr8WfviIT219k066p+BmpwfdrSzXTZFrDdQW2hT6ZP8
gnKged1zDEomisYRg+Km7ldo+JpkkDH3DnpqOMX93u8dfSKwIfw7X3s7TXRYAQGx36d4KsxTclNw
k68AnlPj4bb9YgXWGn7WDR0+8pGMcDA24Hno456BpJTVnhSlWhoPxpncurc4ShBNhRcsTseitXHn
2kLTdcj9mexKsjlDFjy1ZavMcCY5zzhFuZcz++WQ3xWHSjSTWYYe2MzraTz3MaZKrSQjw7amTuBc
37OxHstwWsRCa+/0z+MG1mcy7FBxpdE4jhXJYPSVmR2bI3SI93hkW6EKxm0Krr9lumqu0mPzmdyT
WupM2t3qGeBGZ0ASQ8Qp5noRdD/4tRJHYdHPfXqsUzvJyPxUNzGlX6pHdN60a5poQuwtkB2Vr8np
N6Lxvgbfs1P0BzRKjDuaYp2376xBnXf4rWQ5dYF90RHcC35b5axTfTChrBkm8js3UyPC22MARXgF
BG1E4xDRyzRD8M4HLcecmLvADJkW/dJIF84rhRZnu6i0QICJfTLUsBC3UOrhPZuP714g4ZiDQlgm
7BFCNI0WxbfAHpgnbW2lWVy9CJ5Tg+GVhoRo8sFWDXa8x/vmJHF3WKc0rbITA4CHX5YpNlxCm+uw
h8U1DFQoKL+mJITVnfurHSBIRLME2iFuyseHI1HHM2Onx+1ujpWJDQG2DZUgMSuzWOSNUeAn1M0w
OYq+kr4gcIYRhoLGTPDX+exuEd0EI4KNkP9nx1gXko+x5JdUPx/3OBWgpjdVWx/yKyq1rZ8CELgb
pjclsjWC5Xtna/yNrzXyolx+g2ikpLjhxINbcQt9RPDqdHfR9937Adj5ovz8drRlhFl+qM8ydXAz
MKhtG25yIA81wnIhtTxc4EqJuL1UeR4J0MefKehjkj0eZLrOdQUMqWi3VV9FuUWxkT9TryMNnG7J
lanC1aFv191etSu5FBgFFsdYcqKmgVo/OAXeNnxbwvJfunOrvvJilPRHQBC0QSiW+KHuzrBYWzYN
9i01MnYXUPhIG2hXwnF04GGpkSrWyxpYIfuuLNQ2gsnMzbzA3/qU3bVFrBMRnUBVdJo9pZKHTLJF
U5vwlhVIG7PtOSRIN5J9jawSL0YXDY4JGsEZ8FVQVD60p44TUJmbkTIB5IFoC3NpMV5tZeNNKBL3
MR9xq9Dm1P6aTxoJD3YYiDjedbKTqCMxZdZ5VAxWmn0hZArtUUyUfsKFjuWMSsSBV7nVEeJu1CDz
YqTVLyK/X5u3YPacXe8KIQv9Bon3iEHw2rlAc4Yik987VVIBx3Xj9DYYtTWhPKNTnnXQ/efO+p53
5lgUPJqHY/+B35r7V0BBwuXYOCyNsDy706GFnU2la/JuVi6odLjPsO4VPNP9VqdRhRYp5PKSjFad
89O3gkSO6QO/9dtM14D3VlEiQLbX2B5mVArHgFY0+/HSxcNcDnrPsqh1HnZGmIY682d/bQGIApD0
43mAvgt5E7k0PN3Uq6yqC/jMTwL/6tEQSpHxD2lkAf/l2Eo11RdBUiQTpEyQAQS1es53VTf2vrtF
sBS9e2sWmLk7ZMFPvT6r7gRMKOFYWRCaoOxIF142ZUFB5BPTK7xFg2sACOWIa/vA3qv6IizirYgQ
yZwAV9u97ZATwTXGAI8DvLIGQtp8Gq/y2wpEgBDEpDY4a9Et5SdePAWE3um2qSSxFHaX5B1b6Prf
YsIwJS1yESNvul8eBl7h8mCMyTN2hM5s/oCu7xrBkzIVGadIikuYPLjsj2rmg6oujMmUi6faHznP
X6VkYJ4bozFnKGcZTAqASxU0XzuoYxqq6eKEv3uGmvUauVIoLcgLCHZyRwTVVNi328hu+BIuIa3O
M1aXChiOxLmaPySZDpyxQ/3jn3RSBUlt4MlbJJok+bDeop4OFmZ2Qk0hgVgDZSzK9fynUmQiB0va
PKRy0oZCQMsdZLMMBlX1d/teXqxjBeBBiw66PsPgcz1YOYydc79XUrJmiFUwxpV5s43eJEX+lKTP
QO/lYpl2ZdeI981OR4C1ULV35bUeNk7pTdzjth6G/C9jwkHLry+POe9Qb1V/wDtvMy+nIaM5FHly
+w0ISKkhfHN/dthw1yZS7kLLJKaN9z2my1X+wy1vDqwRHxTOTVZz0qF2vTiAtHncp0JGn83NMpRB
cemMNYq3Y0pqkHHjSd6T4u+5lFNGKUIbHrN5jmrcK0YYoGWPpmcDOdhOiGBdXrRLxcAJo1G22JZj
bC8VKgBRqvNTvpfYWyiIqEmSitfraTInaQzbbv3KgbYt3QgEYSFX0Pej5C+GEKpjnLYm1OoqGeG0
LRFMDhdtA5dGk5KZDLPYtSAnYXZ7W9amId5sIq9v3t9YHs09tF5mh1wS/vhRN58m+lriKZ0Wsslx
8LEdc8ilMQKtx5MF66Lkoz7ar9zXYg7dYz6hyWjcIkgYg+AFGltLpiIpUTrEFFYjDnCQAvqNrEVG
jW4nYjXWAUnHRQB3owsMoP8pv7aqeNkxgvN6rbnZqBnzWq0pOzvp8NXnqKdoZ2Lq1n8lqLfmd8EG
ymahaI103C5LoJFQVsOVwkW/2u1bMfBp9FYmdf+6+6k3s818P2tvZ394T/5rbhH6FeD1L+sSadiV
4qujF7ZEMo/wh9eBqye9cFMJ9gz35fIj8qG1fix2jXod1xU+fkTkEhP0cbuPLtTsr1F4jH2M3ZHr
BWP9qRZizqVz6qmdatFGQkrCGs9WRo+5qIRSxX/GkIvQ1SlLYCHxeGwW8SNC7pEodEi/64BLUYMo
8DG/CvfVwEmzqrKFJTwGArSheLf2m3L0g8t7MyoZlb9ykHPexlcpL3xfAnD90oX2EBA5YnKQJz9N
jZP3+qKfdyjHRq6PZjrlRY6KNqpjUtBYN1xA5lHqHKTl//vTY51+BztlXV11x3ez2sdn74lNTC8h
Mtp4Nn/1LOKLvNQdmjormjKFazFmRUqGPtVRoElXimDyr2rafFDCyaeQHmiG6lMv3B9QzDtUxyqc
/Q+kn7aMTZi5r0fKX/Q7urlP5BE3AShUjvFYQlzeibzOIgRQXNy/vcCj7XlDNdnKlBlzmKLLhzQv
yN9UDUEgaTnUYHsAuWbD0ep1/xtXiZaWhI/5pexTsM9BMMsOxpvGbT7IQfnYiBqyFMNhMMeN4C51
CbKzoDHkhYvCbaYTXgQUjM9Bywsfsu4wSaCY/JKhPENAKB87AP/GvJ97tn+uNuLw+JsmFaflHc/S
WgvNfZfbIEfNMqkbKiMAIRPD9WwBwvyCPKWtSOGylEasR/Xh6EFRYATZw251BaX+Y9lN8XZwn027
KH52Bv9Pfv02GYyN6D5BTLmhsaJjKxrD7dOv58gHe1CJjVvay60Iud+9cjX14Yhgjz3ZEECILA83
+FNf5kL4fIYm2JOfSPemaRK/Cw6NhU7yl71TDb/wTjo7nYjImcsGtF6UZjc20IhBPrr6R4E09bJl
8/3G65PnMrjkHshTX5tmyIEAFB5kSBvzvaBlJPOooIVKNV6aLzqTKqbVUY3kEY+tZW7hWHpj6Bge
UFv5qT83R01GAj0yhciDSEMG1P/VWYi1y6FAlCx34Sn0S6a/wS66NJxoJoMOG0auZ36MuKUjHkaU
TopdciAIQVKifymoxjw1bD6NCLO0GRaO8NNdATEXzdDVSEXtbdmcJXsl7s/xeh55dCqjGrl6Mq9D
Puo3ad875CHUdLWC9Kc2xk8kZrRVJguoVpYC1dN235aq3wzkjhihswjc+OFS4zlY20znYZRqrWn4
pexWM5zuCVyQnljy77d5oadBmuss84V009fmK+kuV18z/fMEDeqlYy6bPixuVCBjOvIEQnyjWbyM
vPh53RVu5EyeMDoo+KP2ATwraw1TMdBF4RcQf3AEcleMl8ecYdeLFNejvC21XqXg9ul48C4K00Ji
SU0jzCJPu81sTLCegdG6277qMU7tZasFTxyRcXFqz6ogchVKo6+nlSS6X1odEYFA1tn766tw8AZB
zEiqk0gH18m3rbsa5UaqRuElKaSjKjDEdYfjDNRi70g0Ta4d80U34o4Qi+GASTJ7I+FzvcYEHyBy
CCGreunR6TXGPeGfJ2e8wkEojbhPZsDUljnl7tLxKVrvfK7YuVQ2A9ZtZQzWYwJaMK69RTbkmn8K
1aoRmZ7kE21BAQfaXKHsihCSpUMmK3ZVbDWddd2obwLrTSvG8YwJ8y74H+Tcp3qtZJvVMKP2Dcob
zYYo5j4ABT0hF8TUQi6Wi1lccQt+KMulYDlzRI8d6PiFeoVFc6XnZwovrj6Dg8DOQVwUD9YWAgsJ
x3ieyTnBJHfECK4fOPKuMVBibctlSw/vn7apLnYxFbp0Qe1FLBha8RjvL0i5poZ7VmFHcTy8Y92R
TtjY4aCWFvbO0ajcfXS9JhY2GaAyoMZWl5mgHrHUJWpJEkIg+pUQmkfWf1lJ3f7h9dvuSKOG4BYX
8aDxpX4WRLoGItSNkT8loRdR/+ht8ttPkyOJTqTcjEAwd+SgImEIn94iEPeK7nUFXmKtr30OAFRA
MfnrPDGqpbYuKvnsM6ZrDdktyAFcztWe6fW1gyxjWjTHFjF0yv6mvUuBQXXejkfPS0ygWldkKjwm
KUV6ZNLVy9JUIccG8tTuxgbvxK8rDVBOoF/fNobpq4f8g91SyEcoCUgX/xtds8vqos0qOuzGNs4U
FVkPFOAPjMsr/dHGmsCLCAKpIzc4QhYB+xaw3fqK3krMDLHf4fIF9TL/EpBTa/qWZdvqHQq+Y0OZ
u7JsEiMd0kWKin20GVFeq02QoN08v1v0bWc4TPLbS6SKGRRDNdOFSAG6UxS8AV44NlHgR2+j+Yn0
jgBTY7hByDz5Pe5Fp8WmkWoV/gzgrp2jx2nDTMQ/XjT3vSwgP6rD+OCwnJk1YoR23USUb1QdtRB8
ExUhftZxsqKWYV8hPEhz3R0kmWA3Xb+ByXs1zQdDiDgRLmZwOm9TPgkqqPPTGIUaEz3rSUvMvPDX
DkVAkxpyv4pVdAB2270sbPlzR7/m6OxkWKB5NN9NPYyf9fSpEen1jGjNujTlCk9x2B37ARBc4S7q
02DmaE8uvXix1kgNlNNf9Cut60haTMip3eOk1yT3xavCE35S4wmi09LbphIRNoNKBpDqC1Uwa0Ji
aG9Ql1bt1f5pVoHcsw6AmO8q9reLUUtSY8eX8v/mn9GAEylHHHlt1mD7fF5vlFf0i6csExJh26qS
uMt0tF2r7hoVZVo1/ays3q/nCkdqM0k6uK4a/fY6tbISwy016cO7dm9qPVJjid4gHTBc0I6qcrEx
axkbllhFcuekzkr2hC1QX8WnHsL/jyGWMvyU1T+xVqYzeL7Ok+HZof5xlyz4HZjwJh8mpS2G9dul
umDizBXGI0kOycoyNWZZSusMGxNc5EqR98Ww2SE3yzwyotheErUNWrJlWh/hx7R1gUPYBhDrt5X5
W7gTcg8ghHrcLsSlYMazB0XFDJeNI84oCIqGCATiUK8aEYrgoSRbw/43I6B51wG3OqT1QiER5XwV
TSraFtBMU/+44m86FsYPEHqjWBTZuWff4qI540o0fc6nIKuaLUICiHMyEjc613J0PcPx9+C0Vm4j
XZKfzOze0UqXEh2m0cCOFXexzPScj4FRwQlbP0K9xP7/KVJX3ZiYeivYyELPVpYOAIHUlT2wHONC
wKOP7AQpJ8FlGTLYPz6hNk865fKb0Ld4IY8wm/eytcQblAxQgqaOf1I0qVNT3EAgX9vv1cVsdq18
ANfeWDhKOC/ggOsV5yS+a2DjOfh+4JzNTvUza29AfrrKQm9ty+5UFvMp6G+/z02qtiZ+Qd1Bqdg1
i1k+DUmzAisy0ojtiCp++J/jfqljPgI7zQRgABQRHYArl7rkpRiN8D89VeAmNZ/fRa2C4vNcSIIf
JbdOEpiDmc2ghkFceQ6BU6pOi3kOTJGqMwGh+zn3iXv/KoXQI4/iv1kBPGD9N38Ie6YVlORjyPPT
bK7RVnoTpcwCBGL3go5ZRDdbFI1yPiw++CNA7Bnq2LAH8LuG+J5XtnPrF2Ag6AF6Ru1kiqYNvcpY
ntRf9ZQUZCpJH9vHat8kmHI09xaPWgK7xqh+ck7m3a0ysY2FAa3ZPpH1w9S3bhQdRQV/TpxzlXUQ
dfPpghUGxAQeHpE0nTlr6NTqPFoCrG02RjKdDGazXVGuHGK4oVR9Ud/ZLzuC7+gFfmifXOiY/x84
thJXaBqtoIactJsfJ3G5B1R+UPss2sEZZ0PEz2LAj6gGo13kJM71xpfol8x6FR8kooGDv6emrhjB
fDwNEfbO9pUaikdL4EmZ5JXSY2Kv4Tou6j2yBEZasmoxDOBe3U4gvNNyi2OMePOoMjWOriTBTCXg
eGfzmnl8OUK1TE7cpdZK2YNbwgEmEZa0Rlhsl26gWTlp3o5IIzJUlsEg+OgOuLb5pTYB5b1NVYJk
KqSsWshpcWrqmyj90Fs7XDeyHEz4xdPs47wouz8PDU/b7a4yR+kUpZCBvVA/L+zutdzVcxvGR8T9
zaKk10A65kkbklLr2xZd2aC9EO58CiMTg+kMMgFiaaEuCERaEu/G2FnBz0KQtccljDcgTZmwVtaf
1TQLehbAGIIo+AzfDysJN4GoeKkX+HNL28uY9u8s/LAlx4exFGd7niloU1q8ysM3K3p3x4jYEGX0
iNY1MuKlz5ieWU92KMwW8d7zkY3C+337nFkrbLPZrvQDe0tDjy65J4b8IeezhOY+ZVhXrTiklBI7
0Rk8rLDVFzxZc+6/vbr5KNPOF4T3HgjVJx5Usbxkt2acojj+BWuQ68xaEPFmG4ngS46oNtK6+PRj
4txB3Z9zQhwmANf3sbuXUowCE0aGKmXTYBFklMmEB9XXWvCJaKJAiHaxKrSD2QdeoIJrOtoBQYNT
dU+ehSrcMDsNuyufo6HfeNKgNqtLsB6QkbeyGjbUjuyLiX7OAXW4R7L4DVeSZG0vLwmjbNJH5Pub
axT8V8OD5Ptt4HfAm/ljcz7zpcxIVr59LWDZgcpUUQFhnAxYe2e7xv7Vb0DgDyYt9X9h3VJZknb3
cEbf8eutnyxjGqdjW5jMZDj7DlTbm6flwT3VIvjhuAEqapA1pDHl5siwE/TNLZmxf7W4Ck5OC/fx
S86L7kgNQawG9g6aSFPESUjMkbDljCTGF9ryErFCdBkcMuKPLvFsAr+g56jeYZQfpBwfoBFX2G/4
cF9h2ogtNFCtJ1w3JG59NhmwvHwma2IM8T5ydIqU26FhYY8agFLjHp2/3DRvU4Otz6Ti3JbKsfw7
HyB1REhGs8xP2c8PxPbsRGszVPEeT6h+mWwGkP/F7N5y4oiI76ZtzQ==
`protect end_protected
