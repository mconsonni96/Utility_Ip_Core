`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
I6d4/hC9ccSPk05vR6Di8h5boixTHtVXnc7OK6aijVR1KdD4JSh0W4xLlwuu+i9FPv79ocd24ObQ
uYNigh6xWrOcOyTimdRkVi1W3m5smu1SdXtD9gnLBftbLpRtkF+xWHmrkc9fQSSWp9qDJfKxdCE4
U3cn8nMwO4eLgPIpOyue04fxFFO6af8jYgoMzmoc47XfenNMIBUB66slfdfbR6OjAMlVoAMjv4co
C6YE0QE7XL+ZYhL5WsR1m9aaUHQcg5nnSCNdBE9kuS1iKOgb32LnO06jxxCjIjvhxVXkNdC/EO4H
/rbcjpoZEGzph/B4nbBXDMyThOMI9zpdvefQuQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="QDfvNPS5lTlCjHUtf7g/dLT3cCcLPesLeC3/V8ndiWU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9232)
`protect data_block
23Ov2fcLODdpc6BwxVItEvQrv+EkkjPj2r3THGiSAN9ipR+k5FrjULRnDC0E0Al1DzVi6tPn+R9h
YMcglTOoL84fv5irBUt26jXxv+b+X98NEvmTNUbKRA0OC5RGbvQrY0Bnq7boA3JlAYHP+ND963gI
T7+5YXJgOxk9bd1WDbcFaZN9qGLLvob5OsgK1Q139BT/6IVVJJXK2voqOSmrRCam2oCxXqu6s1Qf
ReLLoWDcFFg2YYn2yUfB/ktRdorm7jgJMEB2Z7geVlpkv+9M6fmLnDWNOU/qNNmDO8Cx2vkip6Pm
l7HqDRDTbt/cSX4QFM5mLhPdnhg9uxetn9ah4MJiVNETiL2YPnXZIj8UE/rzRmu9KMQJgjHOjZ9q
OhZ3kLdiNSHhkkw8sMTAHcrmi0LjSgn3YKHxn/qmhF1Ck5O9BqJHJjRwSYV2ZN6Zg2FnBa9vWzYB
qtosO8RzqzLhiHut6Jk9pro+aQbMgzjQWQ3P/N1Wk/wATJflokHJW6S8p/JfZm/G8nbktNIUKWet
IrNXsn31kpegTg62KeujOLauQIBBJRzBrJpMW49nXDGNjH12MV6JZXWJ01tFzS0ZF885KHXn7Mgi
iy/qIma/piDCRGS0o+F2QzCkdne8uBMY+K+GoJ2ofWoX15ua3cDkHkUGj95f8vPGhdX7pvCsxbqS
9MxeIFp9JYjneBFgx79DzSHqJJIo+ZW2Dd6GxClb92dACWUcdNN3gHAJ1tju9u9CR8dq3WaM0bQh
0fzAi93nWbE+MQFj8+fn8QTaVbIvGd90OOqHWkPKWBUfnt3rsPCDubpMXe0xgWQv43JwCNGvYr81
fhRqi/S0SrSHjVpurOdtJGCnbnKO754wQx2U0BmcqgqSEUoyhkNTo3pHSFQeyLP2T5I3bT3TfKQa
oARCqZpw5IWTl3MyxyAdQ/maLoZmQhxr6JqYUEDXvtKtZUHRezpqTC44e0tCQjQaYY/5HtN/oLtg
KwWacJY8wN3fnHPIAQ59JLTS7NmLTSV5BF5cDgDSJ68liIPzvNCzZJTnAaGuSLcri5GPHoyaEk2M
BNCTGPspBySZIzY8CHR4cc6zYH/OLZU6/svAsm541d5FE/bbgYq9N3z4p6ymyBOsGgjikNzoEQNU
WgIezkp2KDBgh5F72uwvemrnGVogRGN95etXLxYUiNcWsMy0FPzft49ID74m4tzKOzbP9h7EB5cf
aI+icvpx4n24FRnj3ffDjkqHWb/t4tamBEV0tJvKGzydIyvecrF7aldjrPTvRm5LhevCZOBaH1sG
3US2dzk27IBj+4MqRBMOaYpd1hGE18Dl3WcOWXRTctRI84q8OCxbzskaAuGjqHOjny/nMbGs8i5p
lbrVs7tV0ke0FfeFsgxVRwgkPY9YX6n4ibVogV/sibMM948s0wqVwdGUzg5Ng0Br7sg52mmBA+O7
fFwirpc41d4x+5yqReQkKgckbYWeMOVyFnNIGGRXhWjW6XOf7hK5oabLeGRPbHWQnsfqMPLFqehN
p2nYbmWaBAzV3NYWCyaktQwve9xpyym9FaQoxI83OtJSLxaFpz+S3LUhaNBYagGGeJFg/kO3N0lQ
eNugXxaZbzFEtYp37ovra+On5FOmPv6lj7ij3jVtZttZPNqU9jscrnM0Gk1HKsSs4kM4es/sTUor
wMGwi/eAK5A0PAk2+PliXzeTtLefrfHhifgwZqxcvnusuNl5jD5ELJN4jyj1e7OaDyptUbNpMS+f
xgrL7Y78YvGqksMuTVLYplQ7XzBU3gntAtLYb9wFOZwdGb0oywRkPWpy6H1hn3wt1a3FaNT/NM/A
Z4xkGXO9XG2KMJVQ22pEDmcM0ftFIIRFYU/5FyoWOsh6h3PsAbYhlIKXJ5cWkTMVboZtc0VnAA3K
2vbLHTcbLkqXH4qWmMVpwt9hwaCBBHlhfA4+O/0PZ7fQd6f+p3e7U5zd7L1bxkteyL+8g++eCVT4
4tw6SgbLi4qnK9KJYBRinf7gSPy3/6fXxJXTqjYJ/PwhBIbKNQTdbK11NMHPc3ywJ0en5+Trf0nL
6NEGh/0x77Exkk1bYVrNm3mXlYFrvZMjXXffCRklXxYu+IuudH4mHWrChv8xM1dkHgEoLCl8jLrU
LaOgvbFKxbB3JUjTUYu8OPSyvor5Pdd1WGhwnc0ervJFks4j+auXRQgb7DyCNL1NP7+jkIEZhjKB
tP1GEwh1EyvfOKJ2FrWPfxtyCXNdgzs1Wj13P8DKT0HOURARHNsbniQxChDPJeRB2n5r/CV+DPq4
3tV8NktAHRyk9mlg5C4oEJ7HhCt1E0LmEqwYk0iIUeh2anWWOT7xG/5SZlbr76ZjSNb/7AG603r/
IVuVn5Tndj1jx0bGTuLduW82S36rtA+5zM15V+UGWQ4uU7krSMIM/s3ETad7lF2IutP+uk0EoVpi
ywro0VP9v9ks7u9IcrLGCiJIRq/swHZWod7en25ZBqjRYS6H7BSVgQaRNLAsGsoJqPjrwI0Pl+EF
a61SGRUtVGATtVb51soz230zaUnLJHPqhY9W/aoi1YH3OrV3Y1bJqZOsj5hPtKY/y0bw3FWvNtuk
zT11zI1Ij4qq0w/Fng98FXYfZTYed9rDquedJFnGVrYgcZAmcwB9F+JJ/H19WS9SvV/tlYOCaxcQ
JKoPw099RuS5Kl03gCaOY2x0ZVkbWZwYFVmE/JHq2y1ystKQjBG9kD/QpP/qkfJ79qaMbXZxHZfC
digoo1Q9jFAfNifuSjGwOtSK6thi99hSPJw9uGAc+0IqehKI60Ps8F0VWilo2XEahWBQrsKjqX8g
FbFrvVrElHxBQMnnC4m8QkEhe3x4MT15uak94eFxoz7sp1K5bhLStTZRG5JryrCDZGHROjRWSW4V
zsShBgioDCu0O/5jqkTMlaChDviiPMXFR0LORu/F8TcH0eCZgi001oAgdPDEJanhYYoiu+rA7fLf
7fq2uxVlhSAc2AGCEwLJeKf/TvFCNfoDYap/6sGiXNa+/zVk4V6zIUWnLnitZ2beE3M/tGT+13VV
18TBqThzTt46D9BuD0fezWnS9UKfrz65sNvOA1B9VEUephFQfVOCcHf67dHjncS+RxOoUYDMdm2I
inuDtGrenrQM2y8hZrzlLzTrkUldjSPqRpuhdnvIGiBsflHe966Wdf+EjV3/FZsY5QyypMnUvi/U
Z6d5SklXTp1RFKdCnkNtYmfbC7B/Pfpasj2mmmQAX4EAT8aOrJnNqJgmoyrUQU0N8mu5VnY992vb
lUf6XcO5yTe2bwgiEMucG8o5IR7/8IM3EznS88B7Ykm/if7sbVZ/0mSQt9dNNqOJf/TN6eExOahz
d84hRIGrSwZtjLutkQxkueXdEFQd3nLlLRF+d0FsWGObcCROUKRzTLZ0CKMD9GX0uuReHmD/qBF5
qTnCagL+uUQZcP0VR2Ti5+XuCYB5FW00PXi4gcvw+SwPM8JoydH39cntRHGoLC1TImlL+JomxbnX
Gbp3SSqS5HtjkeM8cCoXOqKLH+7gyukDr2ZLsKILul5pGDSsmQ53kcGzLRs3EZ8qSZ2Wb1GOHkMX
Vs7hFOl1S7Evp/zAf76YnkIcAnYzQLJBJP7k9B/uFNO5fTcvs+51pFtQDpTdJOghzztHfiEGZd5k
uT6UdrU6hzN5M3IzSsEfuwTKYi4fj7Kl9kQ/wFE1vlq5R5QzR3q9/c3Hs1A+/PXvclS65aJGcBah
LdFrPbN04UZFvI50XrU4VShvl1nrAAStExlgLIHNmsphOEnA6OaGc5M/D+dg7p1ZqDWLoM/0ZlWh
3/W173OP5Aa8o37B9XS3pFqs7nPn7q92IJHvIhk7+scDG5Se05B49uphTKKeyFHQfegWPuvXdhhI
Qg9BSo7dmOOCbMyhmo3P8bRWVKJjTTR7OEt/3i4t1Mk+m36oHqQ58+QX+KmZD95AMN4XCryAqOPT
+UKfPVrTRQrI31MfIUuD7tIlESw+i1YNXACrPoanyVvnUWZ1SDekfwKqTdOfCWpnOgq2Bx4U1pur
S47k4h8BBJtwaovixUqQUIU9zRD5O6ChXLB8gXHwj6hmE/krU5XQLcTSb17Kiye8uDOsEW40ge4S
VZbNmeJPH2JG6i7hYCIwzp0g7cYLRta/jevHIecS9hXTSx0gv4slnFrGCMq+xpmVHpGaKrLp/xmz
bQNQB/Mmr6YZrmZnBdQVMFPSMtPA1l0tXcNQUI0DqrllgLVizf8icgeQZ4eB3MccxFb8p+zzMfzb
4HR0WDXkp+yMe1ibtk0vVKxJlu17AcYVAPhg2x62BUj91uzoHq3kxYmQRrUjhu7Wlqw8HQ4zAhhJ
pEU1OmNtr7jqgrDQlkQV42nuXlNKbcUDFqZu6SiAEmYe1dnaD+HQBP9XM9apeEVePMYEsVXpWjGD
4+QrDNNCoOmCKVAxI8fVNCEMZJpFDSzbD3m8JlEwS0pcBSXJTH2ivOUaqndaZdsGw9gHguCa9jbG
OjRRG6utOYvmv2kzaYEb0LPD3UiZ8Nx+LADW2Vy9EDka6dbo4E6KWWupNz9W8tbEJImAANil5L6g
xjjOu8zlDPQyLhQbhkQ49Ktct/XdouFjUd764TOEAstvedclXbFqT11OkQq6WGx3jvAwgiCisHiZ
9fIxc38V2OD/amSVD3AqyVTG4C9lu2Nptn3exzvpJkCL9rhMLXo96+z243Zt2FO3vAOwogDLjZ5B
5MS7vOi1iT4H8PwnNzGdMW8lcv7fkC1s10NuDwB3uy1digovAyO0js8AopkbAqfeEW9iqo5XW8Yx
dz5zcRJagY+8ByVEK8/5RpsLIA4iTeot4gIRfH/tNDhdNA/NvjnqlWyOIgPsfFtarRi+wc6ZDRqk
YGtsAcwyehNjuFfjg8oTa3HSAGRRg4tQwtxS4zfSDgBbteYbQqdnOOvuENf4tbQ5qhvG/IHUckHu
RoeZGt58DPU4jAIc5XaKitoQgqPsJCkR47du+4HHeTMicgLzIhEQjEggLm34jURYaHr4FxiUGbeG
U+kiZ4ginnaLicqd3jZUC30MyY6/9tDrko8H7IwdDk/Fqyo+y1ZKhmHatH6jjXTG90R/oq50zICs
RM3pAA9R8d4zUIf8v6/PEnq2jGczv/guEcxCdiIjbxoLyX+5vKj7cjWZr3SSaS3HchB3X0V+U1SF
ekdP/8fepLQzmGuIZsgS+7gDw6ZsBYpme1Qg5KYvzSacCjBYbfRDaRfmU85Pq2hNIk7wkFLIyarz
MGrlO10wWx+M4yBQ9GjBkbG7fYIjYoRBxFIIIUwCLm83/a45ayXmZW8z9e7pCxzmENEyBKKd+EzW
YKNzKDerWm78zhBrHbfDUaUKpA0y1qdz9zbfgSEbvy6nkBiDItrLPM844BODR9S5q+/PbCh3EhdD
FpyT5/s8EzI6/r+ttFdTEahneQ1WrRgLjyx+R+no2/YbbNViPZDYVkzuGolQPscKXSJ4RovNyn0S
FhvhXuW3HxbztKSePkWVFsvALhu07peywVJkPIYrb6gaKtSrNw63uCIDE8mbpA7p8yBcuXg5gKHF
b26Vo7TaAhlEY77GeX7PesrC0AtGCo6VfA7oE4t81S7wxHdTire47JPSCQS0E6xPPAEjeeWKr4DY
oCunZKd7Cc+g7byBgXrfZNmpC70hTQcwmlWUfu4mRp3qV8FPnt4lm0cqFd5c5UmNUmNcX3rT5i8K
rGPnhsMAoRGfRui2pd4zpuhARz9hFLMxJOJGUb97YiK9uDV/ZE/PWppBkKUOgxGthA2+E2CYiFIi
QfdIJ7vAhOIsBKGp0PJlPTeIeZAiJVdfyzTZlQRz2TRb0MEAMAG4ZZ0/UeizdXPoSmnsW9cW0ggu
nG8AXHD2dHjwPHTCExWUedqraWEhnWS6InaBNaBnt1aJpnBE1L8mSBxZrzCeXzM4V21br7WupKYm
Gw1gxUEPOejKljn6bMx+CxmW/fzFaOEcmC4OlSS2dCnt4jzlkjzFo22+UDe7CxFfZqOx2LP5Zcuz
SEoFr0G6mOdVZijm6p0scKXsj/uHv3HQ98705zRePncBnMhdczJMm9flvLBjwQWln+ruAGKgciDr
Poccq+NaaSaZYTH3P2dgvk65cPbzE0ylkJqNvZEef1jplvgD0Ulkx776hV3SAzAZl3SqijOC/SLK
h7xpq0A4He88xAwztERUthh/MGvyo+eWCJa4wl7NMfgPPZRg3m1bhwlju1vhtUdw6vRKp6sZjDST
VNaVehgIbXqcMWxLC1eRykq/1PGlFVqb8bKpRS4HawNWXtuu6FuybsT+z+Qv8FMSM85vWgovAKxg
YU9Q0y+z2iUXc+0+TmD++2CQtrMiYGLh9KPc/ccHb4pQw0poyHYSxjyx8v3afg0SYTyAMuyntFPG
FVtDTsY7KaU4XW5dVhDFNrJCY1xx6MxXdU5wNiqbELlL96XAsSbhc7F9eV4AEZ0K4Ueq3nbjuU03
/KOSFQ/a8vT+in86+y6/PHtD3qrO7x8RoFM4C/4S54zO4N7GbX1E4P04L7NoNyEeYDds79VJj+sK
9TdgTAmg4bECZn2cPwpc7LMrGibY1axTqu3zHyo01x+ZZwuUCj0sMzSsHZU7RlBcp3ugJnNeWd+H
dRXeKJiyVKvgGCTWQnmd2+yexc7tSVf1HWgObyjEeT2LRcTBaePyAeVoDr+lXLxPCO+AATwcRofW
gls0zrhoO3TbP+bn+g0QhF29WNpN3u8EZt2rty2pSytuuhE+fZVXmxTcNqPiXmQagivZnFQkBsDD
Co/j9cjfaPb0Qg1E9WrQ5wBssnWTY8c5L4cni7JhVx4Vq4Yua/FvyRAUKeMFimflypqX0JqYfuoa
knBzt/qwCqihJnzdkOz3fikZKQ6xzyI3h++POJ6z+9Chx557A9rlOMMVimNlOX1wgVh6FnQlGP2l
ov/336pCpZIy5mZJqVeqL9IUtAGeJJ/puKysFd+FVme4bCQwS2DCcmvmSLOPzMmic9GTpQbB09g4
vR0ACnkzilJEq57dfSgyhPKXgD9zbqbh50RnnQQJDoAbY780PzrhNW0kVmIZnypbe1QyoomjYVEn
UQiuMUgPHIknegjEGggMQrWHh+8wrghPpWKQ6RDJl8XuPY8zheJAC9mKDxggxbOmp8XGJzWkSjbv
WGwRAfu3D1WqxBm/wdPabbYduYVE2cshc6vo6oNNHXUN6dOK7jxfxaNYxn7BfoORTN8rTfEikwfo
55wEG8ee0EbIcal+ZgRv2COajrpj9+3zqVCwqy3Pqga5NuU1LPxrkQ4hKJzKHfVJW53QC5xxowUw
0usIgNfv+iPtSWqWd5cL7PQsDfrIj6DdHq0SpyBGpLS1Qfjtcmk7jk6hqQFzezsF/4axvJQl4rXv
VTwC9niob4EDbzJWYk8qRLhX0eybfMNVRgl5kT4yeikwhcCHoALbJPHGZtO5J5c1yZxzDTeEdFv6
jXepyPZKSD5OqxKbcTWQAz312J8mJqNxRcU6uTi3Dht96Uy9xTpkPPd9ZGx21AiFCNNmscz0r3PO
4gc0ZhNOOCc+AiWhGCYaFjkxlDCwiGviyKzkAaLcy0rCZNXQxhdiMO29BskFuDmlLXxiwSn804mX
Xq3wGVUHndbsgQlNH0waqORnVZsoev5PhnjkJxwNAYZ0SB+kt5LAZFXGacJPaTmZWjHDfPoSna0d
Wm+wFth661KlKtoxWOWL62vbV8xpCn8hfNaVYFSvG/rWCtkSqzM1/MrqS9XkkdySS9kD8GgnMyE4
TSzzjpvKEfxLg/P7vDEhJjg6i5UUsrYSTzMDJ9DAL6Yj9M9VKaHXxDvmQoFvO46IoJd43it4wsao
hAybKUde0h9mDly6Bc6mPHoTjHU0jhfuat4LnGOxAV47y6pa/74wy1xUmPNaQZMmPq/V60AN7H+x
pLzc83g8SN/H8wZTfgcezpKTjBdrkPYd6rspk2Qe3micXiyX5EhO9qB78a5xXNoMNrjHy3useg3a
lxpcP78/uGhTtVRFwT/rJrDQPKBHDn7Nau+ZiJJXA0dbs9UFXvjDJS5j9h/Nay5fXiuE7eVzXZ4d
tFRw552AGnm65fvbSENTXLAbvUjFj1wJYe5wsWqYhuuhgsCU1NvblGlbUNMV6C5Yl9p5C9ZlpcFo
6ctopCdFKtMJw46UrZv9V1A9j751orP2VfeVMW2Hll0UZyEOMcWWpWigjlEL12A8fgdJnKtlHaB9
6pydHUdnLMmB+VUTK5U0x57uBCmMGbG/HsFF8+mk7eYHWKmSyCMqoh1Y0CqaVCONrCPjZ+tBPhb+
xUDY4n2Fc6xP6uRzTiPJtWLfInPuPDwtfDCLe8aheIB2r0Yi4WRTiZyUC/sGGDQW68jsLAI2hRpS
ZDf9QNPyuYEuwg7cdktHlt1PsI5YTRpa8pBdiL9/Cb4bkI5lklM320ZibX4I+FRWLSskn4NtxKxR
0cgOwQ+zRtt5OkkT1EQ4g7Xn5Wdj2z19fYTfsCXN9UAMi5F3NupXsePkj8yOWnm77LxdHWpgsBwc
STDWTVWA81fZ5w5HvyhtABDVm9mLBvx1xebIITjkMsTzruSqLXm633TQ4sjlfm3LtypuGxi6vhjp
fJNpmoclcl3h5tAachGznu63yrNNYOn+tnJHWMO2sS4fdLO+6JlzwakuyVJ1rUR6NYdP5iU8Y656
2rr4q56NEvie1SdP7XaUJD0C/wk0Hb9r9S4QvTh2qmA2aTQE9D5nWFmopIIwN2JgXG9mvmRaXrt9
r9x3Fw9CscmJ88AG3f73Y6cD8auSNqAUhAj4+3/LBqQRFlmTAzSlCEoz7wJh2grMOPpCExscvn9w
RDDC4IACv9DgZWg4yhD0c4AiLRC40REL+Cs/sI+kUwZdrJYKKNMbsJj209Z347AFiBd9w/VXBzQ7
dteiBMqPrMrKWl8jsYTfyqG+SDPPq29VXGhovy29k1AivWai50A6ySn121wXkinZ+WnXZH5qpCo+
VGEWN22HQ31keQiqIfwfjXQtj8ACytX2oWyWFnMbjbmLDlawoJRl9T9Bb2fMIGGvf9LMjI3/CdCl
AxLAotd6gW79YkZs9n2jfjkPgKQ0mKk/BRNgUk8z1z4iLhSpY+t+dPWg+YeFgdyGv44GMXCg+Y5+
WQNZG+Gma/Y3eIGgC8RiMJONU+JokAtvoKPI9fbfeD/zEv1a4enfAiT1AyiNCy/Jj/dDuUpntX/o
gKeTRcPLm54MiA/ANWmdLOsRhWxZFwW87Mb6WXLALdm3+RbVSPZXyUrSnttwhLm7PHqkeaAvF0K0
rGLOgjy+x71/7HeV/10eCPzCR3Fc/r72lmm+q/kbJsrrpjsBRFZd01HM4qY73Bx5KTWVQIFOx/iw
t1NJz3XCmbU8hEKBCo7/qPA5zu1xNjbvw6kdJcP4wxUThuYxKVUDNK5vGUxPHvuomZ44v6PG4yRL
g7NvGRh6LhxxgHMMzCfa7jFcvjb88E8H1bzGNDyQDSUTbfVHUkQcDDPp84dnHeoZkZozOusabku2
dPKuydlcFzD39hjfIlUX1/61g4W3npCwGE3zQlZLl5Vu6zwVGIZf0m0b1jkFI0qz1bzjDfTviFOR
WvXdW/n1C9DXo8gnHln3FjUBw6Oclgm2fx20oLPBE2zUEJWGXmtDl4pbDwHkvWxcoYkKNb0MRrsP
Pn00CB+JBzR+fD9QzJNVf5jt2nYMkAJRzfdZSE53FP3PHL1Wu5zHl/pq4XJxD9pmj1iKoH1RTCys
cgCbn7jv9vb8ISWVa3oPabYL7AIMAQFYvcPvvqmHqT/8hTQB060SmscYsatB5HRT7tBhwZf0btZQ
lBmq6tBOMkWdw7M01h2oIvPhxaJUxwAuCJYD9DT/W3ppjZhLf7lb+EmWFKBbg1k5zvurMZlfxwS/
2bohKMaa9Ld6Wz2nmEhN1uWWVDVs+hwGPulbNqo3XbuoMN1uDLrxTXX7Q8RD/b+hh9zpxJG0OrJr
rN+sivw/Tq7cWrct3HdNoSGZVFD42pCpVrfKHV6vqwnjG7HeuaSqF1GNiVsBdic/YNkwNwXEM/D6
dEZR8jGqzpylKKYuzR9qqnpuqMSfi2X3EQLJxEemUot92bxUjQ1BUjOAP0JNo+BtvCafqH8SKLWd
tolURFUAAgbtTvUo9E+8Yasv7CfC+U6FP7S2JtiEiApLgVTTpzH+xsnc8wBxMdRoapsCAiMhoyts
OLboAcWIv8ahdiMEqSfks+5wKO3Y/XWlaSxJiCWJfkfnyRUc7J0fyFAIXmMWrk5SyAjnCNxQDiau
gYdR1z/ZCEO+/pTQXxwxv0RfrX+gJel1aXV9M1wLhFTQ4R4RQuUo9T8EcZlEzLgWSICfeFjR/Qtm
r2jLvPxjiyxDqd1gTJ4CBENALUsxKOGfHbRcIPRTW9hYDa1nzQhAOAlnWP4LrQaJxKMP12eItypb
DYMx4jVg/He0nMz9dHOxr6nOlKb+cpp9QaL6rA//JQPSSh/7nTKWig3RNNQdmM1wVwyLgNl20TIa
4iP72Tax9cXJJtf5LBCJAd8BdbDdwqPA4QE88Zhgl5mnnWrcgjictD5xfr3cX3Cii43xOp8d44ji
CvpSPb5SvPNeDi/dnoqNyfIVcGl+BGQQVxDky3cqClBgc/idCgHdQ83XW+WWbWgrOXDCh9fQ2+OH
ChNyZL97mnmXGmNwsK6phip/2dhsIPFsDglCEXE+LxVFyfzIN88Ofl6GgUX4gGlVWq3Fp6q/onKt
F6ZmUaeJluo1sVHhUtO93FRSTwO0lgvZiS05QSjaiZIgBiPRgZvsgdiHWcmg2IYo9FlNOkzU7X58
bCR83nBjOwjGcxvdEo6hvG8Qiy4LeEodk3XOTLY3MPMfrY+lx7W7GSRXDTCaHce/iumh+61ocCdG
4ynhAVcdd89gmgSzl+IxWk+G4AKr3DXZBfjJQX/2zLqxqA/IhzatTj+j6mPwy04LI0S0ITFxjEes
k+c3Hnz/VQr19WOZXyFc7I0iypLS7zddnyvqRn33KgHX/0mVyevVR2QTCwgl8ahN/6xcMUmF7qx5
8B7t7+C5ojSYgeKn1yRwYOuZQ5joG/NOHJ6+y8LXpIsEm8F1hemrvwnxbKv/4DGU2TwR3uwu65tI
mG+7F2UqnFfSEci6JhdfcLuGL5GQ0bJePe0ZH0pp5KP6fJ1WTmfKNy7zz0Gp8rhhDjfLPIgLMis8
kAu6tLD/WoLoBKlF28bD3TjhP+DWtaAxKyGe6srT6wIomlNv5/uonMC7wmpCwvQuoKudcmK2y30c
+Br6gFXgqcntYmJvBqDHTwolntOWT3sngbGW66cJFzEYZNkU4PCmQWACPWHw32IyvnA0LlX//vlt
96UCfStNM4KXGdIqaciFjbTo6/Jl4hK5JF/+/To7atwRR3OmfknNee0O469q14jd+3mZ+gr/eW7y
/72uxBYqfeS46SkEy3o3T+fIpBPpsyI/SsLP3/QWN3vNFWZlzPUlAqVh1/u3HahrgDVuc3+6Sp8e
Auq7TJnItWVSlP2hWiinet1XItFT/F6QSdZORF2jUiYOpp6y4wgpADdZq1MvETHWAN1G48u/Sn3I
JRwHdBa4rFu2e8x2ZbJevvPRPU7dJrf84nVztDtYmKQkKcvzL38YwNXVZO19bS2ghfIR+7XB6TRp
eRg1dqSoJRFEme9aIzwEFNUZNQVMCEJUWaeCx5fLmF998Ok00fTs3zY8EQ407phjDTexxTVbuJ+k
bzFbexi8c67C+OHqADRjHtKAV5KZ7F/S51tZqvRvAHNfLq0AMnR8K0FTILkS0tBzA8Wzc+YJCoA1
VRS5W0d/8nsEY3fpA4QpbAxaWIs+6isyvkp80VxSe0/eyIkGZ5feLo7smufJmKKQnnB9dCYfUX5q
A5axkRkkOHPndrwWrhm8ClPsQvEMX9iNTJIAZsgwO5Oh0Qc8G4dWCvjEtLmJFrvetBlSU/CZ/cav
7Rhf9ReF+iP2qjq/YAMhYA2jH7snin6T3/EHEBjh+uyAQJ/gV37OqO/IppoGHKXFOv3IYTCyFLQo
qKgFLX6XpO6ngRYsyyKHI2pWbcPeI3BVR7dWtYmciWs631zDOIVW8I1d7RhoxZvMmqKQa+pMfymy
zFWgteY4k9Pw9D1I7NqtQO149BkkBU4v++HaOcoLBiwburObL2/kqBCGQMTBk+SWt6R1xAdaZ725
e5oeFnx09x/xLQO/xdke9lGHeI0HPS6lLbJevqGZy9A9hPlRjlMtp6XGU7oLfozncDWw9/LAteHJ
Zx7dGwn24UWKXtKtVFezm2m/y9WNhHMFNCbu/wB5CGxuuxfOOyfJCI8cwx1QsEXzf34gWKfzSg==
`protect end_protected
