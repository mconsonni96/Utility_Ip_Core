`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
abEiIGJNhzS7llaaYKhPrUeEWliUJXbXRMu9YJ8aJJPqDVkFNGVRpRuOAS/KM9zAg9BPOuvxY0EH
gofdsj0DHdka/v7H/Phd/9PNP91NmzCAWre4NNLochxdiSR0eWY+C+37slWJm88VnHECRxZ0Zk11
aMI+pu5CP68U1Dsgr8SyfCUdjuVu5EGkW+md3NKRaUPrHsy6qRbjkOmS4mZLf7g6yJ3BAdVxQx2c
X2OsqMkj7WQQwEysNPl/TPlDq7IN8DzOyWiHXKFnLxpPLHDXsMtEuunO6yJ0AeySw9WjzoUE+vwF
Oqrjco6sbEz+99DoYN960+1e2Ba8jLfUTipl0Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="k9zR12EVyFcWhvJnn5m423oo/0t3LSQxmB8JT/LKvuE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16320)
`protect data_block
rvM7y7tdy5nKuC7riHhUZuxBHsCQ2FsRfoONJj8n/nPkUl4OPKPXBC/MutNnRTe0k99HIqwwitKT
o0TPD3hi2slL7U5JsJhmeOu335EptB9mY8pGVuqTpyDV2derXUK6RhHEXQOVHH5Jqba5DCaHn15O
bgg2QtALxjLujnadSHQiu7eilkCjZiIf9AfRGcY8RCWfAVcAtzHZ/Cw+ufJsMkWBsg2MjktEwn9i
CQmvS6BjmwgqmFIbp1iboJCRUE3qcichOHS3W0oqsl/QPfM2yYSZSdKgajliqjxDaxghWjCXbkIP
DcQ108dfbcnqSd8Av3iiCe2EZQqIi9kioiyE1O1J5uGjn0pO5/QU93MZ3i+rrEtTYqL0hCM7YBYK
97eax7V1c3Eg+SxezC/g2abctcns5BUFczU/vaE9dp8ZW2ECM+vJua/igdT/zmzab+RSFFjHWbyw
IflGNgKaGnOF1k1r751lASAT4XFAc0L8qUoTg/3/rSIe4m2BbcmPq3mphD4E6oYDeg1fr+6mqWsi
uvKHBh+C+zipWBxZcwBUcjwZBSpPsBBJMURFtL9AnsXxye6MH/JtnjaiWHThCIDedge+aFMBUozH
e8v+3CkKMW/k6EDGXvK8xtzFu6Nnf8fwr7Bne1lEEluBA8BG1+sxB7dav0qR76MH9O3KIj1ioxqF
stQeGwraH1MOQKvpIMvYbYCsPgAPShqEcTPJ7dyAZlI+5x8yH0/CdNoxXsARbvHH+uQGOxeVo7lo
chlf6Iec0SEG3eRv1Jy2/jnoJ9JyqYTP+VPvdjrbpN8Ix03nqfMFkgt5XZbiCI0iWkoWia16MJf2
F0pyHPGIe5M/Hhdl6pMCwn2RPp56QOlv5l233XZxTLEKHhoO70GHTysdPeWtsFcHqMXO+GJwK2tk
aOgdZ4Ac+gv9duAWQx7Y2cegI6n5NbqpLvDP7VELBPIKPysu/z7cFoCX/uHygUvxQxlgC7JWg2Pg
ls1Rz9kACTrDfPVzJNg5ezEZbABSzTIZkT9yfAH4vgA1A2TkcwYU1WgkFNFhcuuIezkBz5QNyRB5
IFl7iawBOCY2cO6EnZqR8XR6hoSkpIK4suyWg36sCKm06CjCvJAUDnjDjwThUrmWP2gR5H+/Yc2i
3J6M82LSM26UjkAxmzHp62Bgxt1DRZg2/PEXTjGLyF15N85FYaZM7UmWGBLiVxqsPXfpcOCnnbrV
Icmb/vJ30X61Q1tK2srxRTpY+AcAEwRx0cffZIvOl8JZ5znY2urJfzowB1ybrQ3ww5eB5Npb7tcO
TAjqC4br3SBk0MxfxXV/4YfT6GmxeoBiLEqudZ1tiMA6PQ/T74capW/HrMFXzFbMinRnyq+hfHTC
MdQ4sKfz4l6Xqs4oC67MGy4GkYyS++ykcpGGSe2LolkwyacPH/s2xVZI6nlCFoD62uhEdFfoyV/P
rRtJAwFHejyg0dQHDnDwogMZiLa8OzLXA/y+iCPmZ8PBdf9upFH8MGd+YVFkzi/J/qPxE4BYqk84
KplkP7smvh5m7aYbF/VF00KMHCHWV2fCK6YO9z8WJpb/Gj7JsvlAXIBMTIloyw5tp0PDGJIis/kU
JwWxOuppq0+D+gkQHi7iXhquvfhOm1zEETNTO8t42xhtI3tTNqNBVy4EIv8Eo/nmNLwRPCOIqiJd
DseLTB/4Ykh3IHUjnAQ/4KIVjDtK5QPsyj+zi5+FSyK31R+gsQ2eOEZEq6V5kNt1mKYRh0RLQ2Rg
3BiIZ1BEAM/huAa3yann/YpBHaw3f1RlNmhOhxToz+deC9KgiYkHj6sg9tM2wfq83ZM0I+nmYaes
SQsmSATZ9hKs6R6+P8ADs1319L7t+XgY5haGUgOS/USx27hG26jI9PItLafIYSgRD1bWuSQm1Hcf
zc+bZxOFw/x9Qt8OajGr2Wg7WwRRIQ+JuCVSlZB9BKZ/sFBjuJKXv97plJZs5WDfbnxSxOF/l4hQ
Hmcxanc63IAafhbSEPPMS5K6wNK2xGS328ylLhYy4hD/+kPWnLrPHWfzOyTN5D6HtzAPR0BXzj7j
zMp7dCTKlJOxAuIO1r9qCLtzhK/P7ryrnGaGHVWfmOuoxNJMNnaaEAz7EAIqbeqYPqNz+qD9UDyX
umjCks/Ecy0HxKLytdSju+e05FhrDo/5rxfwAClSGf5zocei8D7QoqEUyXy0K6N18BGWIWi3F4vc
jIDbQdodafohpn85ORqot27qOExxXElSeGGFN2iblQeauB+0xm67bgIfMv4RcvUcyL94FLQIW/7A
B7vn0QSx7r6vWyBdWU/vZawjbjZhaeW55E9SS+9SmjB+/a71yjjhzkbBRqOKYIpnv1bkWn55gyIV
F74Tp8a765A0nNrAb9OnGbnjBYMXc6jTsckc1EgMZ2pIcgXkPfyTWnVO/mRgh5s6LCsoRyhbObfo
G83o+dZ+iSJWjgPiR7GZExs6zeAxRJ9zNskdWAkvumhZPBHaeV3XWWesvKol+viNM7lKbVnZj/rU
PbVwiFkrb9t64DikqXwmv6VHymTxwSY03OtjcUGYhCkNkvNmUtxZibAXsNzlQIu8QdN3NZVLx+5V
TqANVSSeysiX/vun2Inlbq0jSsxECAltV/f5z9ek1v5i/UQczSXV85VPDqLqu7rDXOboJ7u++HMG
RpJCRh7EcsRjn3PBcQcr0g0tfMEBU2s6MmxkW+o1qfs5x0+2jemWTUq0/zhw22HtUM6fgM0TVOZr
XTQ6SeMz5UzY5rvAYYKQEiFZK8JsY2qgC1clOpbi9FYrFRNZ5w4Scn0J/szGXb+XPmJpr3C4GGp7
nSW/B5BXJPXxcX7+Nw2aYHSGEimbpY+jhx/xKHQuIHjsoho9rszvVxDKzBzoKqSHu1GrL+v3kZl9
dOY+WapZ4koZPuS022ATsMv4v5zoQD2I6hHcAQJWijnLT2Wvl6vfrcrxTrcvpCZyKLndW/QmZ7rK
Xz72DW3ZKfzWlOY5SbG+iJeYUiX2xXWa2puLKVFDJQ2blUFnA/RnWU2LfsD0KgcXCpQYo8F0rTFf
POG6AWD5tTAggOKGyWOrgeevD9F3i6nN2/EpqCzfmB3etehAMjLm82zztQLOH5sabD9OOMJ7jbXn
p64FCcF6j0oKs/H3uQWCo1uIdX/ege9qSjl0Qq4htI+xTT/JFQ3Yt9WhvseRPXoEyUJX9tIlGjre
St5U3Eu/dXGqugJUxl1L0Dc8CdCYD2u4+WJQmG/mVoBIaaXmCt13Tv7oT9kmlbunewpUMAz3tWB/
h/2Y3vOkJGamnjl4X3USjID6olNeCTIrfpPGNvBjlQEXLcEPpS96GFnBMjQTXz7tv/M55wIv88on
YaxN6ze6SG0J5YRisuAEyAMjqUG6NuD1Q2DsHFX6bcd0zmp+k5V50OiU2V2fBljs5KOYzztkbady
4kJLVZuWILEEuTwmmgXvioj5+p1wOK1Snsy59orW4X8rHXqd9QuyeaAUEY2rev03ZRTGlJN0QchS
LwOv8xkJNy6GudorMndN2PrM6HBqkgjsjSYiFcqkodf4cVH3nEg91Hiif4CSB+KxYxGmBoN+eKoF
iU5rYIlZZcBwMYRHAWZZQfeXmrjwA2dMd4bF9edx0ouo9ll//hYD4e/rCgqsQ6eK/Mz/peeBcNfp
l8tBAwXgpdV1/YCKVqdfIjofMSD7BgqctBF/aT+p4qodavzKhM/i30Bg7Umlx2DyyVu/Sul2JiPA
J3iDnGvWW//ZEmxbNTSNha1/oHMuFFQWmI30WK7CNVB0t5hJ9PWbZexqbZCTqZcQGDhTPe0Saj48
N3uMEKs8NLZfIfKjZEmHolsAxkbiJUxCI3Ajfh/QfLX6pqwdS2DPbZj099+jU1k8ljOEiwZri3uA
c5tpdph0tYAlvMs00ZQ/hNz7j5k5ExTVuk+U3MhsGDiKUpZkUUZiWmPTrwmdT9ePaa4qoi6xLxoe
RhTl4hhQ9Do2tLR83U7GpAL5Yqkykm80SY12JQN6ETHZrPXVPLyIkbxRLaaMUkOTrKc4aW/EzuQ7
9Lg9POolbfZTmXyS6X9WoUNTKb+ClQR7v7a6Xu0KV86mscDQkPeX2apVEpH5xjiUwTcOd9xE6+2Z
6dCcLsCF89nhvpMcRJvPH86BTwHuWIe8TMcdbN5I8+hhx+8wY17jW9IyC2rtCJjFr+58knwJtbz3
F+uviaU9OxniV6QJU9pQADZAQ75z1aTP4fERrTGqzfAbVi5kfXqXx92j8Pkt+YcoQ35AwnfLA/mR
BFKNeGo94JYcV8hsHoJeXwkqlcg0UthuKnP7JZCkIyXgHG/sToVdYVLAvdcpp4WhPh2joT5vkJVq
iaPXltCu8qp4WTLdNY/dW4A60d1LyGS5Ge4NjAEKy7z3Qexuii9utcoLxR03QdNUOkI8JxVRFcdU
JG7dRdHOVz5NspQLApkeUt3R+86L1/IauBGSPn5PW/BjkmtXGqPfuyEWPRmiQOWNCQWAVaynDa3H
rmAaBYKrTKh3vAPXvY19RGy61mAENhYs3A3LjDzzoYVOMA4+UJgPibjaImaI4SnuXgZxU/Xpv8OM
Qv5RV3Dm9asF95ZaWeCUWgKsdW37m4BJnGDchv3eYL7q9rvA0enIxwAKdG9dHnXrKg/AITkB1Bxd
Kia8l4fBcPtTN4nZ/+ilqyF5AWyKo1MeGMgdatCanGV/TAGiKu6tx5cVaQ8JlQ3zIpx089LO/iDC
iF+7CWEEwaUBoeEyZYNWWhO3QI1cSoNZrG239zJhs892poqeai1nXfHohFcKZGhZL/4NXLxf7Aea
jecHe5xIP3/Pk342KVgQhv/19SlW12qp4VywvBBg4KXgJbPWBcyhfMSpvrLyzbN7TL1W57SHQfDC
xJkLeX+/0w06bvgCy6uFk4g+7ykl0J8jA4xP0Lkj0ofuf0iy47LhQY5Ar13JYLSqqYkDslx3vH/B
iwfZ82z1mxhzLOAsRiZe1iu91VL9LpmXWTOXz5FOEAQfOmVlhaTH0wUJiHKNTboghAZEcKgs71iP
jO300uGkeTe03IuDcqs3YRLI94Ed9mBKzEN1TyLZBOt7hF/aQFxTPpwBFq0CNub327W4McDtT/iO
/2+NZT6L+hifmaUT9YToRS2pLpI8afIOsP5urU2rqCWcv/jLAfxdkJ1+LAEU8EoHOJ1tfgh2rUw0
a0mhiGblwMbh5Aa75chdScUPRmLrtKqtk8aQa6emZUMSyZrxMZzZwsWBX1qvBa4KVOFx1zRV6eKJ
ECfiv82WIm2+HsWdj45LeID2GizzkoJ1fmaTxS8iB2rQJRv8W/foqD8lZbHesOrGtNjYHZ4Yx56Y
CsgjciiGlXNbN5hbwZxLwI0h9zk4zrSIP+QdwYLqHHKfD8JxJGsZbRPGUjgUa9H7B1uKRE+C5zwY
qwvwEbC7/Rs6JYbqvlKHI9O0jl1UZnBhqq7wlJwiat7fIId9gmOgtUGcTHOtZ4UdFchLwCYhsg1C
Xy6Ghep/k8Ou+W3PO7tHwjxbx8iR59RYXuCTz8sqelNTo9xM80LB56FOl1qtpM64ol2sbP2IrI94
gmciSUNwSlv6kRXtGcfcAfSYZv/5yQ2TCxSVZt+l3LcQknBxf0yioTPRK+qlyPgpRjdWoJZ3Nuhz
9mF1PbTNZJUOUJhWkdVPbjfktbFNkgu1cylzUEgRPTHTuHheLXpsIwIQYK31IQ/bREi4V9eXB2Je
tE6ttqNRqAUmoKUJA0fazM9oUnO1wkfWO47HsVC+3zZLFcBjdEv+v9eC9QcmUWQ8Qet47M6iPRCW
ew3lQyNwJfcN26+pGOzOMnrkaTI0henk8GxnDFFpg8jGBiC/MZ5eB+nhhxNNrVNWajk8P2iYiL2T
lVdlnOa9vuriHKy+TrmuJn4e9mWYMW+9vN5aVh8vFe0ojnooBMKgPb9Y41jI8QfZNPZNOG+03pVz
kePAs+sDe4OvgdL+wPQJIv5ECiF6SCy3/06FjKXHY9CNA8gJKSjeDvU72FAUCLm8NGV7DAcAYDQa
a/hkRbW8GOPJhEa6vrBPkV7OihlA75EXO87l9d4Znd0qWuZkew8UxydAEqGy0Nmduw+ne2ACQzDD
VqZjCB/sUOJhG/m8JU5YMTCG8q2W+UWH+VPOybWUAW6lbVOZrPm5hbckV3w9l8SBpLCkQPpVEEKi
apJlApe5qtrA82y3UrvOIb8xnKgGwcAaAKNWWSSdY4C1bN2f0uvH6rAB6ugHQ/VbhTw8vmvJHVc0
wTToKP7cWAzw6wEmu7bkfThM0Ku3D1P3LJNqg+IWtG5QBa1MISnXNp4wsu5sBCoO9zAWQaFwoQTH
P7mMYv6lOaIS5fM5jqJRyx1zDGlKq1OiTXmtaUsh1SKGzS6BXz77nNEqDZ1GOAhqvbue4CSEq4uE
TU1eik68gFivhhGbY/hx5Lv04Vyn/XH2wzVdXZQ+XAhgNT6U6Vu8zk/zYPitvGmdh0fahLgB0j3p
vlln5PxIussvqrIwAJ81GoLd9ld/LO0qb+5Vw2RVLQi3mLfzSpV+4fHNEtXoHrfWgJRp5UMGvbX4
z1D0eY9ZVtfcsCFqnI2ayrq478SdG675pIu5ebUIM6XJhfK0pyhJr1Xe1N29Cr4uSIC+tC4MFvq0
jUSPZGIGBFPXREE6Cx/9wPJxxpgwAwWS6ljntTQsU+J0ldM3DINjDhRr0+CqvCcYRhUKnDPmNICM
sFtgeLILHM+eY/Vg5KcLKElNu+y+T8NAm9hb9s+ir9OUPwY+ZuhUPTcPoCkIIxtvGo6hePD4XfyX
BzlHU0thizn7OXd7qH5xnF8X0v2SEjrSgwH2DcGjSpICc2F/kiMs9R17X+Otx67X9LZUFS96rshX
fiXlUMiijO01Il5fU2puobzgN+sDoqgGGLSzaIuwstZzddUFIxckIx/xgHh+VwMPhXRojWMo5FF0
QmxAE7+Bb+G15yKvhHuDRXQV3R0PobHWEGcNhG1LJs/DhaDek6YvGJZsrzv7u51Fy3GiuSkh6cWU
r4l8sqysA+syI096BSXOCN/Fa8eYVFrTQ/5RfZdnQTZphTVLSO5inGVfIaAc8d6nnsCpRTFb5NSf
ONzVnrnuhoVZZTQGRUMN2gEoDwy4r8YKx8aKL+gUj/dn6AfE/3GmFlXR7PRFSanmqzt2gPY0lhmz
lQNl7FyLBjXOpmnbY496zK5EbX0FSbwR1keJT5fe9UDrBUMf36BmPUDVZYIwHdP05qG/kPrPOVUG
iarOD6GMH3cyLO0KhOBjMsRlc6pGqXIxDaSnk9u3oTcYIEOa3L/rl4Y8c3wxun6utxDkdZUWd4uY
u7GnJP4xor72Rf25m7v8sQEsHWHmYSL1ctQ1l+QFDH7f0xJOcbCpuI5eHFOxoQoGLqqDHLYimlA8
T1ZGISQAqXUSAfgqXFKlHMmRKguxxrER3xAsf06TJDT5KvGh44Sm3TigJl+gKkefLfXETZ37V78b
vf4/MQWHbzVyjursu2Q2fbnRER9AG5mRPuVCPGFGGvyPw0UJPyGNUIRbC/xxw5DVmwWYPPXiMyN9
yll01JKpeUAbl6oyus7+P51q2Ea/ou1BJxayd9tm2pp5M1AnJkDZri3gFlG7vyN9uLUCCDHlgoim
0GDm1vksFxB4VWweAsk4bayVz5U1oIPADEibn3mQDnfZNmIu7fGpLLHannkmdclkPqKrYDvF8I20
fwlEo4yciq/WjfnPpV/ckRInTo2tGxennfU/HZugGMa/Hjqn/2fkQV/g5TgeSCuUlYpRe+K++bdl
uaj8WzdQgm1wjqDEmQ8sRklQcKqOEkEvHZCdbk7jwMbwf3rTSD2fTsYlJoYnIbIfIBbcXGYd0FrL
PpnDr5nU6tZLUqT5NL8Y1dyh7uH4ALKp6nRKMw67wz5tiqhPaexE+zW0l3vGYqMdsPf88OUzgEvk
kSBQBGgPYvjJ07e8uRLGQ19yvj7kKxCebz79kiE2Zjwf7aez1TSxm9jw7Z6XZaFgRTG8stIZbEOL
ew75PC9jXw69JDTx71g1Ti7KzOFE4oYaH5zfVjYBQTZYJWjVt2uySJx41VGeda6nAjU6+K1//ni9
ggrG0dHr2JdEAjEOaQ2KllLDidIhu0xRVDhvI7VK7Zjt+aG6PbQ6TAzyCTP6l1KjwyYIo6hE2DKE
i20HH8FkQwh86MQarVYThGh4GuWHqjehxHyM1pwk54PJ75fQGXvsuGkWyx+Jcr8yhC5VmLslPsB3
typhXs+78bvJANPZa9ZJviDOfreso2a/B2P5IVXFdpEY1iKq7dkqguziiNtl9tusBrcwHHod3sYA
0YjU8eNVPvMmuf4NFsexGK8bazkIzQc5xrHmTYwJizb2n6RTLF5MlBKeSR/Fo4XmIX3q1UVzRlno
vT/Br5TY04idx9cjrCh9hLLgJUKaXT12ye/isRlnxWmLy/68NzFomgqSoHi2pTlzapcxlE51XNS8
eJNlx9ALLPyF6xwvi/i0k4K2aTMXuPyO/FwtnOPNY8UJmteOK36gBownLiOVYkpWykzIsiXTXEEr
gcZg/t5oEeEpQYNQaG0S+gcMHYrQYFzIMBh/xv0f4Wp5K5VDfXjwtfjG9k9FHV51Cy4n0qV9prQs
jv+ykhnJol2qmvpvTnAb2dcp1NWp6OOEUlY9yhlNtOd4BF3Hh/CNfoi/zRnzcdjBCxH9Q+GThyY+
pE4ATYIkFj7vY1c7TxSJIuLVhKXsBVJcNQ78AttOTS+nx9IhtQEngb+5C+H+cbkRAxb4Vwqi6zlN
lK+VZ7bML+omzSZnW+asxstcvZ1LM8ydIEeMg+BAy2Oz+nIWPOJSkklrdPlCff7QQ9op9v3xXKip
UaaazxUuo3F4jnCgwAMQWmK6u7XCzcZFE0XPir+H7+VUZEmNPzC3lpIq/Hnkm8AZ/jBPuXHF9qVA
m1IfLVlmbZs29mLEz/kEME9JhnUuXndvIWJTjof2/O9663K1aKYZG3/zB8eQfkyJ2VqKmC9sdW2p
z9L8unpLEeS3M5yjdnaYum4Ln9oIMYSenFiLypiTAuH5mC3DTjDBWZlcAvCTsVW3X5vk3l+CqSlG
Wq4aU5/R/oRuKhShh+SWMmpeOJf+MT6VnsFX226xWSIThlpRsBjoqNGgcJJsrv0k2N8vbD8eEf5c
Sl8b37xPvI8YNnlOF+Yikvpfh/45kZbKZhieOjoyNEYXxOCwFqBX6zwkkhCBAW8P1woHtPixajAC
wDY69zym1ptbdZERwPACKlMlsfs+ywNQz8S7V/JRtfwblIcTL0IQ6nPemVc0KjzPqvAIIktmsGI3
X9ALq2EQtOZoGDLu23uOhY6F7OHseLytAsWw+CzqDLG20NbwWdmLQX+JxOi8QoaTEox4M4ksZoVR
oVWn2kw9wMuQ2Q91IG+iOjmEAXNiI84nIbZob8H8Q2DtBtr9mwGg1n584zxfC+2T6D2wLcWn6yPC
vduizr6DmX8QcNqg1ak05WGF3qFpprDXqZmM5LUdgF5wqJNv8L1lwm6sBeDWJ5oSWKSwxrXv/qqS
e5j+cSGBaxV8G+k+VgCf54NYgKAWjYHdoE7gG2jWzOKhKTGNk1lbg2iZlxzQOSF8R+sF8D9g2q9E
rnevCaFjkwk1hwK3m4OjHk6Z8r97eCZ4Y0hXIicyzCxmbVmlWPHFqpNU08NQV0ZJxIHJfPXhXC3m
0vrmnNGPaI6UHIGXNm0qep7y6xX3JgQHSKFMvqKEn3IPJ3gaS8YMAzExA7WhfZwGcrqwIeBAUBGn
TLU/+8EvAjm4G1/x3tgFcndoFDLgKUeemSZjZc4FaAsssJqRTKmWGQS6CL/2lMBGPvmVPgrLKnJE
z1BFBPMCb2qVYlO/psrvsCl/pJPrqU1Cc8HiHzceOx+whTifs7scl6OyqtW46ROMv2WSEh0VN60b
Ps8QJTG33mmsJ3RHdTyoGpYSPP63krP+0XTB1WdBkAE1uTUj+v6Ul+a1Qh4pkrImQV9YHobsqbIE
LR+n5K9LfQOV67vX2t+RS3MjzjZeSRuh85iwWW9PznPF4aUvJeB3XILIwKfBzvHf1lLID82uljQT
pgoZ8ay3SOL1Y1NcM+4UDcQPKCa+4+gDmdKle1Rnj27rLS62JGnrijhkhcpuoRAluQGa+A4DOvLI
X+ntaGdfDRLPZ+r1hpZY2hOiGQpp9Nde/m3WYrU/g+FOSnZtD9cvL84CC/E687d/KjAZeM10VYwF
k19Sst+LEN1mZv2z/3IOX4Klosv5wJ5ChDS+bkD3l8vnpZMN6PGR1LodRdK0vwI12Jo0LZk6By5T
d34PzbQq4DpOORbFCj1AD+fSxpov4dYexY6HMJsA09OE1IWvLC0E32qRTgRoeRNMzOlhoiHyVUyg
oZFGwtI9JpMdX9dpVHrVF9/8VHfqZo+cpuETVilp92yUA1zhRN4Z7dWUCRRXW8oVhY9w+6Kgn4Zo
lOGVMW18pLAenq2KIAX209M9OcHJaCJBSJI7VGKBgmkbOlveyJyMnXD9+66Uc7ililR8etyPfLEM
Y5PdFd+F8J1SO8B7f8gQ/NnKrARTozV7QCmGZLvRBlPI85eO1TEtrRVuIO7H0dgt9P6Lw2ZrCxpw
p9y7HEJH1Hd/QJVMysgt9Otq+Re3TXAO9ipF1M5yoNQsZ3yuMtDVmZ3OcHtUl+ngZ8Tnug+ZrOtc
th6DHicr1rZgU/uZlpRP+9dF0rZMrxWBW0SINgbAJ1Xn0WiuwXB68J/eUWKBWP8JGdWzwujSB3vO
Vrq8wDlRY/mVdKt/OahenerQSAMrrcPoPbz7sbkMB8jRgEndJ1K5g7gfCEGo+4i7F/G2wXSn88d4
K1bo7Xgv6b0fVdS69tpBFGe9cBW+Wd4crZQBdZQpLRIBxPqC1eNnkScltHfxCvVDcaY72ZGfAFGb
sNWQrosTX8quU3soCznBpBXcn5xe10chOoeQvyK1SdcnbL/LM6zz64+OouxPmuouINMffChDJ3ao
vGtCCiKKFQWCE77gbD281bwvzGQ2WDfvIeyO2S8nFCeH16L60LeRbE0HWGc+eYNn2Xmuu4Lk9e9l
8NxKvqKhh7BeZkg+8KE0GsQQlBWFum8TNY62mHrcu83c2cprSn0fLFsgpsGNfD8pzZtVXkc4zJvg
NSWs7GSwbV3B//XC5unfui7WCEW7ClxSwapxwxT9Rg4IndWgHsv18hnfxtoIYIqsvkj3NyedHQfn
wTorhkL8HB8tKhQeuNUZZn1QrTOxtEzxbLXegO6+D/Cofwmqj88TlTtvrr2f3vxtgYsdQtgtITSZ
Pf3AcE3b77lO5kLj/XIe476oMI41iWjxhKwotLHipFc9XiwRn/Urw68AvLGsextbSOPnzz4H7El7
jyoH9551baO+zQB0hJLNWeK/gEECo6D+p21gKIuHQjrTJSZt+HpZZKvoF2r+G/uokKSNMg1qzHJe
s+3uREI9/f7zhrpvIMRXEMHlyhS20z+jzSfdDqRlSU5hFGKLoljdYoqR1x+QURoFGt+KPpWP70//
b2bV5/zGSZQDb9yl9erCcGktdiNYLYKn3tK0K5bOEmDWpN75hqmwh7m+Oxal75C6uGVoyX1lbsgQ
JVvhkx4czweauKO9T1+GfaHAuulP49xXcNF/eepVkStXtWeCOZ4kOcznt+piCGV9J3ttRbk6wPoW
bO0o+Tof5YE1JsohtnoGTcqFeneKujTsrmwp0ZJsnL9UsyrAbneQn5zv0RD8KEIaBlm9fkEEechu
zkpp6jcuUBFJkI6GXLt7FcYKGYMbvcgGwCYRze8LSgh9sy7zpcqYFrVE062dasPp5QdpG6xYzUmf
msqinfhTGGv8qgJg8WCyNLoMKLweKuroj7T4X6I/2SQB4HDuoeUYLGPKLy3oDXVvvVX7TbKNy4MA
9x07Ea1tmfPUKuZs9x/HWR6DsDNuwWFmLy1I9Ethfw1KeED0RFilKabUFQ7iLVkCOKA76BUYOuPk
4ChFWp1UZlcnlMxHIr08t6AID8qGXX9qTO9iYTrBZ3JTtXouX5Oh2iiKrLSyVOlBWHMvuwCcs+XT
PuOBwuy7Pj/ref6DjqUU/91REABsq6GMirM8OPM84UffMHgAsECIQCIQ6f5i6q7Vdfqk17Di/Wk2
FMY3yPjvoGekgBuz6SR7WfhKKRkJ9w2wSDpv4xwkmnc/gPAT9SSNxI3/Uve3/MzYGrRMN5xyraBr
+LFmzKMNs0/SEwAi39yAD/AtmFnzXekpG9l94dP6iSiot0EgKuDac+JxQZaz4LJnhaf0vVaBKVZ6
6bBvbdJpYhy6jWXVz/InPqgDjTteMqr0CkXNwGXxTLzKVDMBkJQsRWwC8feE7HQ2LwPL2Qpp4Upq
WOA3GkL3/nkWd5mvM27fEuHJZAQPgpErqvkMnz6cY9Dj8d5ppIu16uJ5TorXx1R8S2mFUrbzPwzb
ZhkD1sNu/P/7S3J0G3MsQVvCRYriR87hilVytqEZ8AWSTYahA3swyeqz222tnHCKmGhbUFS5OPsK
r2qLKxLqrLCr/cj8M7y17syzjrNm8bHQz6NpbmRgA4uSogABtRI2JhLXhSEdDVI2s19curZNPHFm
q5A5O7h693J5Yza6b2Zftts1j9zBNcSaJhOhMCYNwSwMGsAwoXQC7YA1Fcr2ui++41N2bLzdtPEk
JNjYHGj8x/SMFOsO9Cmv/c3k6jvVpmROloyPI0sfWQ48abUh4rpYmsx6DTcMV7RPM7fWk7V2VGLW
J+OHMLiuF1DocowcsNaQnXqLxLhktagZdyG9uQYyEu1q00zFoWl2USW7LCxICHfyO5Vv8Oj8LANQ
op3YbjvoUk6GjlhbI75HYbj1f6i+bcwo//ddwY4jvMFwD+9OSNXbytstpArGtHyYR1WyTKra6ZgV
X8Qj6WEwzYhqNNQxjj9oIOS5Jh5PVFoeLiruysRxdsNoj56ye/ZQ10vQZ6ytq0twJ/g+GzSshBnP
yeYxu+iKed8ewY2GymyodSvbM8BECeViYw/YQtFdE1qFSMETYFnl4BKPKJRz8QbjdWxM3VbC0paA
9/JIsfzn7BSW/ozRMZmKhxt0/kVXMs/wx4OrumXk1VEjYvh4/mZ576WHiCswmwDivQoYXHS47WcH
zK88VKpB12H5zsyxC0PTMZkRXq6ZDyF4qO7rmFRK8msCah5Uk8TNliKQH8c5a/KeG/fW7c31FqD4
TN3qnDBYNRdcgsN5q3yVMoIT+5brL8XNHcNqEjqU1YXJeeog+pbdqKzavz08uuXHQDX8VKylvly1
Tn+s7SmDmWInVJg6bQB8Qu6jT071nPNhbmHXUSnv3NVPUh2c+5uxGFXllH1DpwIWdxGglrgOoaR7
RUBfMGl9/TfNW3dCvoHTs1vOq4HGB2FBnSS2dVJw666MDCeq7spA3xMGjH/+0fRQwzu+gFdSu6Oz
EFTz4LB5foUkvYGl7GPbF5AYqjXTz2VMbviY3qkG5u/ohF0Bi+sW3tq9uujre2Esln9PT+EjRTUB
F40hb+sW4/ejXzoOpGcDRIvmzith48OeC73/qQULyOa9a19SwzoHKojjZNMaA+UGucBcH55W6qBC
NL3jDtZ8QOQQ/8TX3/7OqHybjnlZ1iO+u+KayuH3xYghzQEyc+H06nvIsaNhIzmpnpJmXVawyWA8
apsCJ353n1aAu3rXt5GVngEA2ocAxd9E0BcZ/2UjQgQtq/Gw+H/NGHae34MyoKFoC/EIeprYOOZr
9r+ZUn3xIdXvk1H7jTVKneQGJJE4w1sBmW1yoKiKCi+Soqvg8sLCj6e4cCuf3VpIDs4ivkLtoyav
ulgrdwt7KN4ycYU50MmG4bTijIz6qJAFutFR9HdANKxWoVmmdr33UO2jDD3bzBHNVwv5BYOIAC02
ajF1s03LyPWVN0ARJehT/DNWizAESmN1U4BdebcXg40Jyf2gaFUWyz3H2H3qPBT4ol/8Ew3RXb9Q
rKt2nPCC/zdQQzISAjCnbhLRD86Xik8Nmmdb05opP5cfgJ0RifJfi8if1H/O4tbiLO3S9ri16RE1
KI2MWxX0uLY4suY5F0HuOUbjyOf1NLQvm/5G2cl69PHFhCYKjPzskfUQNoUZwsjHn7J9K0H5VHr/
GfSO55YT4p1DnGKDICKHood+D6EK6I2IwYsVOZMzYosy9IX72FNpT6tx4qh0G7t34JNiU3ofnhxH
VAu6obBTFBuwCtIiEz4yeLN+Y/rvBLnqfM1bfCdGotPoRKrzNtS5WnSkvmhqN0lOrAhKQAdJ4V3G
Cf3t1h4JhwgMR1nMCRpYatoGicXAmfCsICdLGIkB6dcI6o4l5c2J3NF6p9ovKK8NyQEm8NJ8jSFV
03wgvyUOPdZdEJsH30BIRiy3aSQg5jgkkYH/OliDOBTHWGICSNBIosUN/GbHqm05/avoBjhO/ahS
TbMZ7V3l+FtqczF7HI1SdIt73Nov0IPbhJ7d299x1jjY1BeO/S4C2wCoegb4gZzgeD7AvDibDLII
MEdBKKIlsTLSy1Vi0QHH/zTX+i9StJYZgQhpFijDggkz46LjSYMvBDKzG6Bei1EpTsxPVPJg5vBN
u9WI8V/idgHQEZdeAqvavDIdfLBC+NLWvrPqxV2o3DC8/+Xp66FsBm0r/cDnAmXNKeSuIQ5UR31m
XiRXsJe4W2VPsUAcKeXEyTs9g8k1GT+GYzi4otAmZRsaiCWXmnKciAr0ugYUL1hV5Wf66GYcE/LC
ikBH4wC+ztek6khewd0zc5UsuC2uLubzY0hI8EPYJYKWbrx/yaOewtne0Qk9KD26hnThuXEtwGd0
Kk+IlqgUZZ0Z/lg72Tz/gasFU5DOpcAdaDNgn2VcQtbbH5OyOUmrcJwcEjFWQpIPqy4sfFWMnlFI
EtfNNBBYkmIVrQKHHAesfureCwJY+ugoGUpL9zKXbBQ6n2KPLUR3jjkvCrbA7W9UMmHYdI944OgK
Ybgl4w5yZ0uv6zVevppMcgVSd+kpeaVwo2ClmHTrRm+S32UVzJ0kM0PF5ukreGZ24R8goyhCeYaG
mfsn9ZZsg5pkBov2l691zCmOO0ksZF/8KCzwzedm64uTiQZVP5ZgHoylXKvzp2HN9C/K3IrqbU0D
J0I+ZP84+tXtUrfBgCPRsQrkH3xFZ7dPUCyZ89qSRyBXsJMdR402aXAPXWMjr12+mPvsqI53+KIU
wUE9K4MiOKQLce0dpryq+3SiTfxSk6rgzpMTRj7bwcJHF8oyqIw3/Jk6iP2hnyy53C/b0AoeYRsI
t+FwDod4G9U9uKi8YMx+dTCdAZhj03kOaFUkZMtqMEVdwM3+78u8dTuvrdfG0xxOseij4Y2y5Sys
hKrdLhXZHu7w4qYtc1VZDLaZ4R1elGMOvnVYdv5MSrz4/ADHMDZAGY/MG7sEhT9ETwY2iBvzwDOW
VqKKrDCTNAEr3t4xLALTTLiFhnwRwAEombma6AjAkFpSCGSghV9KdB8IVwVrNsdKg4xRJXGc9UOo
OdWUzn53nrvDNYLoSumdi96W3KuxVx/ZZp8/AtZuiqCtWHq1biwoxIOjf+wg2HZIssU3zKntN5Tk
1p85sp+zmS812jGrf9S+yfoTQ6VmoHc14OedddgoTwEaRrcElKLCl6nRChKnvTD39oitx5EApJvw
50znc7od0tFf3E5vf+SZSUmMBBgiXxstUlnCiCO8+Si+Ob4xV4A68SYH59qhlS/8zUizfSsojApm
XShq6xHj3hjBbvTUcu/KKpiIgEA6kXa6922grwohCE3FroW3pSBUPvrxOkmlJM/D782NXyCbxFwN
j6ek1XY1fp46SD0oLc616/IqxUSjFxl6celRGkvCbofbTWPoI/kmvJ0Phe0blz4QuNHRqsO3K9zw
vNm84df9C2RqbwbOwmW9LV82Rx/LLjmv7Z/f/RIV0v3a3ZKxX64OEIseRSBGFxEkYyOaWl4uLKtY
2d9rxr2Jt8CmAdznLUYz0rKmHbKA2LqMoKCZcAOBHK8QjKcsovFkK5c6X5wu2SGwYxM0Ah8/tgAh
nk0dymmSkt5bpqQymkoWNRkEomJItyhR+jFKteejHesuKTgKQlmkDAhDHxIIrnMrCRA7y1i/zADy
dmcuv5RMBoLtJvCCnV/sJFP2PvbA0zypA0J3dVeDIStr6B9F9khs2dCmwc4wPKkIFy7Wo5ofTwpO
WYU41xeLqM/B2twR3/whbxMgwchfVW3XT8eJu9rfhzWXqoVwj6UdGwXpfarAnLa4iYQJPh3G6AAK
MQvP2u1bMDvprBwbs869RHYg0sQiRWP0/YAjQqgWeIU6cGrmjIM5sEZDq9ME0KHP7pQhA0ZwA+mz
X4SyH9F2tK4XLx3TGUsSAyQZtwBQtOY9ZUYJRt3ZDxoqXg8gijvMlpTdCIXBfd2Wp+5oyjvqup4b
itPZLZxAggpluFS3mL+RfhqyJBBdrh+aynvhbgSxR3a3X14LheVfqQtymK5OpQIyZFkOKsaEZX/B
YhRQhxXEO+YvAoNcIulz1vpSzFHx64O1K8Sl+sDRo21IpkGVzzsspImF2phwc755UeTyWfNkN1Mc
RZofMn+oYkfZXPrG9j3pfGKQ58zKMU7S+De1J1Kb6WvjmWFU14O7kxpugneSGj7o9jyjO2vF8zNO
ArXvx6lCczeBxIJhfDZKe8UDEz9XS6vtib1YrwJWdKyA/X2s5GvLKfnjjH+KkfxAHNTn1vE8uKJg
UTxiU9o7KjFuiYMMwod3ao2e+Islip+CZ+FioiFzwhTxamtXzqz+dwCzLWnoDxCsgWAaZUJXuqEG
If22HWl2zutDYYIAWrZSz7rC7Y5svWVFqmk8nk0TSCcQcixpSFnCZLJ5Ni2kEsjt4en4y2P+yrd7
xdhNqk1tGUsVE2DA6B4KI35iRU6waaJaMzjrcZOQV4R1nipdXUxiOwVOmzDPScYsQPe+/CLbHjQ7
RS10tEuDz0aQBbq+htbgkG6o2v92t5N+rpkF/8rLbdB0GHPLmKBWSNubtMKm583LGAUBJeWz8SwW
gGRFEQ3mHF+zwxGSR1xmdNKETLXMt2E+mHsrH1s18IuDdOTyxTQN8MBVsg6rGohvG0Tey2gXV0uj
SFcpXapm2JpAALOHJr0ZPgLLk7z1lK3tW7EvehRCcq9ZAdLY7C8UCXEU8SObNgySXxlunx5gS7BH
4HevMHkR9NdNi3wncuUZ7+EAwYh941e8voFgYtE6DTV6YX54C3uXN58PL5WsRyY8Fdz/4DN2nfT7
jWF3wI4DN7pAzTWgWgMKAV3HtAk6+2sMgBX+BLBVfcLldN4jyK+mYjqWHPQEMiJaka36ZOpMVD8t
pDMlSpXaQWlZmT/ubimPLDJgGb1vHypll+TOSc8ALMsf8/6URIzRHCHTrDDTl8Lzp3oLvjYi17Dd
lQL1MwmEOr6c5vxAeV48KD3SJZbyq/8rPrsb1R0pdXoRYuvyageUSiEVUorNbESUf7EriSWOmaUN
pgjcDfajSCnFR/A3YXAS0vFPggEmU2e2cJ3ahwuJVEOOA9xcDXKAcHOhykMO6+AmEtkuCa/64rO0
+YIjl5NOXtw0+lfvciSfJ1oXPsKO6VzoCPPMbYcnWTu04eW56abXLqIkeIjA64qC9UZcOjMJLc0D
UJfbkJHptefvzrijW56shBOAqBt/DcE+V17E4s00g+6UBwwedenaNoHr2a5YCqaVpHZQe8shJQSZ
ehlOCIJVuJ2BkFt+tCAiRf+wlzIyoHPsGT1hRW1OVGLbKFTRteIJ83Lt1+R1+2rWlZReN1Litwnl
9MEshwT2p4ylGJn2oJpv7NtsC4Aw8IhZFeR8J3MeF4U4cFPC4y27NfcpZUD/sZ3RnY/Ugs+AXEjM
7bLfekn53jbxxW0Muco9glbBpg0reKKVHUa/OqNfMZTTC9PUUrD2vQlr1o2/LnQvM6eP/8lCWItO
fxdKCsS7IU4WhXKKFTjlelLTpUP9djTQJ6yW5D2Zdi/wI68AloCRh3DPPw/th84P8wzaqCA/zQ7M
4m9NY8NdU9kadpMFr30u7fGcIhN5pRajl5Kh/NVKVQzfD595DOvtNn7m4WWerHEbpAAk6FO8wS9y
tAveh9kYPPA1tHi8iM9jO4ohlkGwsdvn1uMflJy69SBUPeDuYmqSne+7iKql4lz1umUNFMpljZea
WJlMMTnfZUSvTnjV0JVNiOpDcxZ0pTRl+EhK5tuHc3IOs+NXnI2QcKZLY+j2J/FQCNH0TIBZoyJi
rqsKg040f6g8Y10TrUgd3UNfvvwNrTmMAxbBR76OZqPsFF5oEW8N+UtquZ2/hbr3BmgPJNj90fWG
nGYEjG+y1+qcKz+jyxSwbQ7xKijl0xBWwB024E1GHkeKZ/Q4IcoCH54DuZrvC68GyRFkVB05/SDn
OMvCjHNXi8w4qMk3suJhnYNydGYTlGpin4Gbe3/JeOpBFrxcMKlZc0z46kdHr0Loe5UsXUz6/mi6
3nvaIDIK7Wh6QXgzE4CH/aA17GDyM0MXPBY1/bTNTNBvQOfkj535kiwvmHc1BLBXqhJXQmLz7ouF
fQqBF3564AcH+yXmVfSh274/ARY22E/Vprlh4FhxYzWYn/u2t5++q/KQm2AlMBfDUuo0yZyrb1WG
Ugm47dYM9xiLE3s7i1uMq8ymmS6yUSsVUsBbNdZqzTPEPonDu9AHK2gNUjio5bsT6ELN0zr1Thq1
WrUTCFTNKgZOLC3vw08NpS2qP9PGZjak6GyRSVfBxWpkfalD8Rme4V1ytWJNZG9wsV1hgOHyjBS4
/JvK1xVCOwraH8OMaaYxRsvmkk8TXmdUV5pG+RbTXGzYzRw5/0FpKFO1KNKSLMuAcDU7TChOk5Ff
hWe5kzPEnJe0bHTIVpvXW/DwM16WPvTw8y2OsuTg41BsYxwdmOyLIS2dJns4XHV45Ue0590q8DLi
RQcYOBO4uOBDm3vhD/VBjjq8QXPfsmBHVTN9KW8XYAThFWCWULA1lh1zFIYarTt8UnHNJvs4jMmG
bpYqwgq0BxytfFx0WqKr78FFa/oeB6LUxSW++uDXHiN7wcBZZ4QXyncHQRjRuJCYAa75GaBMUBnh
vG5taVf6Ooyv1IpZb3Am9npycg9sCoHsUexmrWFP1Np2pxar+JwbliknEWhkcOfi1sIUBijb+MOc
U4UYB+F8IRM+V5bVzn5l3Suw7C3Exw6I/1y68vYC/77TvFSu9KfmxcOOvTY3HyD/bg2WCY/dLAHy
NOyIYVjFT6liwaIyfyY49l12HfgHbNuhBD+W2YujyV25Pta6D1U4gM7azNIeCtrvqyVrPC73lwLe
B84suWK/ivRegRauFGPV+GaUdPp2/k0lt4bRN3aqf3ELOWgcJOmQBjbVMPB4cLxYnWcvBNWZDim4
HYEXyasc7hv4hZhls/TaWCJhp4La1Mm68Zdp8T9EsljjkXLEwGNErItDZll46afO7vdRTV4WwxQr
SIqmUXQJJv0drAyazEUshE1AbhvrV/rmrcq7Gbd3czOJhCvbPFCwZ8O4FVKwe5T9fP9DPDT+rOPL
aCDvY5mEqf80b+oNLtAONNuYf3wOxNLOaAFyTprXc6Vyai1450xnSo5lZOrSNA5p1yNoXaxZcfqg
7YnLddLTCq/fFTKQd7NAki0SNsCupwN3YKCdDBszOXws84wWaCp/sgbB6aj/M0WHxR1XqXAIuPwu
SOA0IXu8KxoM1SBThmMOtp615sqO+qlZoIn5grN1yVdCESGBsrf7s6Hv4TAyCiPHKAkBgMYXWZX/
ZoZcdJxX1pvOKV9OVckFmstk7GXt9/DJECbor6gez9HzxG08AbxY+TzIdbVQPUPMQ2ItONqjEv+i
pQC5WkB+OojUmXLKiauKEPw68lZQN0bFq+FC/9H8E8Zuh8Ow0JTXcsCSoUq+7Walya24KgouVwT4
mWWL83MYwATY1jR8fdSSWrcLcdnu5aL5wDaQ2DV47jHmvL1Il3vsg+RfqHSmoDx72CTm/KPX1ICT
R2kNwG4RAnD74Fy0LA8I/rj8ozyBdpXxHuALRgNH6UT5pCfGbqrSjkoKTym3JJBqN5fjs3ybdxZX
LB9neygOXIiMEXd6xnC/IXS9yLUYS0MkDCpt/ATAvwvRFcLLkrxqviV/XPBxDJLmlrDffackUnz4
bUkWBY/dyNNpbss2JNnAw2KzkveSKYZl8bp7zH2VenrBWygCSAv6WZSsRF/hT1MMJofCaS2VsyxZ
V2nCyMf9efqy27Rq3Vio7NwoKhr1xtPETaEQmQPq71mkZ2PnlRNhsVHYqbVsxlT6SxgHL4NdwgOX
L0TITrJ+JcLgQVHGVO/nsTL20Z9HrtrF2FBYqtB3WfsWh0dd+3uLSKOQzQ1eukAf1iarXrigVu4h
adyZYA+us5ZrxrmtXJWXVZDrVGxEElnFTOre6fW8Y4agCTMgPpMJOQYAKHwv/99OciEZmYG2kd8f
hfq2P+QmB085u2RIaTDsh3rQCMFFm9NELMONpeQUEBxwtpZKYbe7osTgpeUdRY92dAreok+K9/Bt
GJwNl9MzUrEiSasBuiP6wSAqFBQlK5Vi1nFwBRmvzYCHcak7zGVj0O9zHgobyYdZL9SP0wP4bV8G
vd68B3hWm6s1ODIAx1l7wtRF7KQ6bUL7oJLF1M6Q4Je/lLyPAoIJoTt2jzAl/SbtItZSy4Iwj3WY
DAQpjjWrGsk4gF7gYRplKEIuRYa7y7s9400uXElc0Ahty+BexsXAt8GbYL/1C45LBjDMg6VX1PqK
NgHbI7U6KOtYtgaoUWY0KY8i0HCiWyczVVKAcy8INQjg4ffO/Oj3yb+oVZXX75m9ykn+23l1LCyJ
lNb3igjd989MBudNSMV5+UOfxs2VwUE/oprGjeMQdlWozGgxSW1iU8/zsDfm5NWb6o+8mjVdYz5Q
F/ncNedxPwR3nPLLXCtTU9TYsN49630/8Wv73Jb55lgFssDw+Gt+W5F3c2i7ZO0M1et76c1EkR94
TkaxLrWzjXjay7rJpysRA9Bck2v3NmmHR/nNAblm0lQGlsGLxIOvRb8enLLvIL+gNv71/S9nt1aC
8uP/lkcRqedUziqsidhngPpNx4BOvzzRvUijmy+ZLMznkaPVergk7kjgqiLCfRdn3PdL5IGTvmz7
ilVifEkcR0KtEuoiWj4V+ubuYVXQuQRP+A+VgrYpxvk19/RzC9PWUoBbNvySR3qpLsbkzi8CdYf8
wQD+V/LbbP04X8csPFBDd1KlKfYXZPaLxwKIVItzgd0tGFA88GHc5u66gRxRY2Dt3gyubTb7InfJ
GhTM3m52XI7t4q7xWe9yDTNwJg9m3RP/uoVW8Bk2XlHcCTSlr4Pkr8Y7spxdj0NrmafCgMbtoHyX
d/s40nOgwe8p2EdevOMvXt7nWUyABi2VIa0Rgc+n2z+a10rb7tHPf/2JjonNZpdOuwyJ3c1A0vGv
WMltCy7AWqhfCMYEo9UYVN2EfSz2ecuvfD7NtY43Rqn5SXvnByofq1f+ctkBqyVqiwuFuOVSFp/z
JInDuxxY+ergDFN5n8MmKu1Mi0MdIgqcKxpWeGBIo49AfZIj042Q9BtG+urZ1x8hiN1fX8erRoPC
YouZLwMzuQz+JFj7V1ChPUdgeUOo/mf0G8GJWg0I9D6gQVLzqxskaSo0aFTLykhce9zX41J1nhY7
s2h0QD+0AtWF0RHvIqEztoazpomZ7t1HlbsOYeZUSGZ52zsgxLKbm9p0Kj3zJ1yWUfVEYbnX6hAC
lbUD7NpxGGysrQqiDkfDSCUuXDLwwZXaPSJB/oRsPGXBCLiq293nHhp7MlbagWANISzttSaI7uQz
XSP08r59y3OmJzP9xQYK7UQ6
`protect end_protected
