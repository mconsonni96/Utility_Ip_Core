`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
fwvRoMsY5esf1wJuMwFS2xPWMScL8i17FMykIuzli/NRtRd7wT4An8AkqeMg2FYGSXPJw3j0mwd8
5fhLCJnPaLd5UWhQyIPQB25p9MDYm2vbYaVWaJsM3km6ZhTNnDUkGIcHnWuE8+ghO0XviWNgUUqq
kXv8PwOYig4wQM5opuJTIXJingVejjX6/zrcHDjK/gvLOCyjdkfNtlX1HuFALl2phIGtOTktjjxM
9yGOh39LFaqIjahmq611HVeYHAixyqmXeygMPF3bmfozXIEYuafa0BTM3SsSbp+jHLhDBGgsVGZf
I3SYoFq221q+mDYSonv4RGscFjp94dv9rhT4gw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="3aFqaunnO7XHzFIx099ayqJcP4icTlWRalHaG9JENDE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11264)
`protect data_block
/H3APbJq4cLK/Va9PFU/+8NaqdJi471yxDhrntJnFuec4FNvYN//2tbMMvtcbCLBe7snn+3E9Ftz
ZqIZ+XY137b85Q65vciWB5SD+LG0XZc7OJhqVGcrQUkTOvh03sxujeYg4gwMa+P6HvR0ZpqC/BVs
YDQHHqwRhCrOtNPUqEdxWChNv6P7wTIXpi5V2a7L1j6zgrnuKS1iW94jfAWYEJTkYMQAzQvGqfeS
PwvOJnbuv79lsvUdCfJo0LSgZRhRBT32W++wRsRJRGtojbuzc/p8PCRjR0zz3vQ0/61d0Si5QDc/
Yuipl0ZPcZgDj5ywMdtg5SNkMd56c3fV9BMEoAKL9GvGsDR8hp0zBCFJHNCIPfxYRPQnfiHuXxSa
TJcESqitESUhPDRq666SKNcWszUiWLzXrKeVi2N49xvU0ZoPBqKVLMJvGv0/BwxM6l0pkbwcbjyY
qBtapcIQmViaENpyXCO0ASQ3gMDE6hSql+8N10FEzbe1QlV+Mm5VgAI12hCFF9dxwVr5P+m+bWyB
68ANCHiB5TJVz8hesqVX4ez6Mi4Taqv2NauNH036gVWTReHYBdIyb1qP9k75EYcxeX63YPvSNY7K
qkjC8mXob9i4L7bWDZQ5V8ZbuTw2dUgoAhtXijQYaanGtoaA0fpkiu5on5eMIYgpl5SF9/IJyeCg
VUWMrrEtjEpsL4kJ7+u5qfD8LH86eOCRtRY6XDjEzsy2DNKXuS96hh+g9mb5QppuSfFJUCy8pJak
0q44tFML+uTJOOt8sdNtiZne0zW4StPNBIv/bG/Lvox7c6jNYVBcL22VlwyUMZx21weOB/mrMT5t
OG70keEpey74Sq5cY6FmaoUKk5H5f8Hro1lbpFLYK6G9+dF5jAPeQEK+bT7+zs44FBf2DqYcIigH
bgdlwBuo95I+GjLwVpPHRwwiAIKyVa/aOfCW5Z2rwJooCzv6JNk/MSaqa/snZ0Mk04uDJejRIKcF
ixWI40m761ahw3o+qBHAyKvDmpw28r0nyVAjZFJPY7LZLSPFj7iWR3cVWWIGhMoBh3QlfuPaxlPG
cllij7BrSqdjKxCVRSO2YolutplGPiQdWp7w9P9tpcNSri3Y1n6x2hdW2qAFfLjgtWY+eoLhyjJ3
VebIu3rrFPcj/tooZpq7K7zaQasnqA/BIMRk/DskfPLBpDp2uYmCwJZBLNdS5GmtTVw613MzkWN4
YQqpHUSGyUcV6K/B5LoRpgutniYL6mkDgc5xv/f0KH7+yGgGhImDvmY7z/T1HCbT8cGxPB12eX2B
uVt97SZlgdee87o9vFVuhaV9t0Fap+f3qHP4TyFPKc4vjbssjzBfixEPEFOfPjmAc5rlSC2C9ij8
rI3f4weN6Vf5HBUuxwTBQYNicrxbbxgkt8hJoTorQB+aM9TeNzmsx4+LhEgda/s9qdzQidiuHiga
37PGgN2B7HUsL3jneyMihP17VjFnzbIVR1sj/czVa0idfFsNITbosMjPIXg9nLf4DRChdvArE5kD
r5I28AT9Km1Fuk+Z/N8HbM3uEaOQ0YpVpiUFMVtke0luO+91ngbYM70SQA2Khy9/GCr6eAe7h2/H
XeNpCz4OzHeuz1X6HHSm5iCgMW0SaPrXxhyDVqHLumjf3UhN5w26tUwPS3+Gz3zx7eNp5ixju9tn
Raly08mnes9chsausGTzQfH/99d7H6imtqiJWKHBEUjM5KtEQx+gLYLw6OGaRJ7+4BfAQORZL0NS
KM2im+GR8O3ynzaj/yL+dMfRZMnoofXtN446L3iI8Y3O1n09iI72YyOmi/MXRj7NZhHKn13UXa0f
ngzrxVM+GcUNCLL8Nqo1uwsVcPc8Cmmz2ZEGUVFjEmbPuHW28PkFdxOzY2gO51fHQLnIEiu4aEaY
Fs1NnkXQ2xDGYwPqaXdPElUBJ/d2TOqLXy+TkWx0geg70oVk8ZEjLeRgRjOF/lE7MEyK+bu14kuj
tyyD1D6nzKXynvb1VbbHlzmut+t8A5EpDFI5mOVOs4D5r6BDkjUwy+2RwB9LKxjQZ/uYbNJSJe+d
s87MmZ9WR37e8j8LJCqAL+FPuhxktAJGThcEQCVqy6a9J/iC6wY7kkGd6MLPiE23LixCBfywUgjq
dRVPx6TLt1vxkOlyvnBZ9Zuy2zE7rMU1UsHcW7wlI4w3L8xy/92bDQ6hxXFLrXdXI+ql6cNQPwV7
Si/2eYRX5IPjL3bp+IM7ygeCaA2b7PS+4Wtwg8NVXxHlssL9hutBw0sROH6dZ9c1BsBrViqDevlQ
ab8lyVxUQ7VTyUuXD5b4lZ6ARhi+wxjJXJHR2DjPFs9BhrWk9gR0kW82wn4Jk+RloYXMDidVgHRX
Ssg6GoM9o4NpSAGOBbLWMKXPAEC7WxXRFxD/ii7ml6iMu9WdmEx2UNC5/GK7zLDzG1P9Ola7oDKF
mAaUAjeTxXgZDylETDFM6fdaOH0BZBPVcIp/Zrs6o1zIT3NEgq9BhVtTqdz8gP+xAdgPwmKMijUP
Gsku4M06WmGdaZAiJLzbQ82E85llvJGQiwehWtfXw58bOsj8dtwaD6ZM8Wu/glI8FC3Ze6HPR1h+
0eDxtmMJb+e0q0WwtbSjiYzF7vUoUzvo+h4j/2Sx1d6Fzso87/zslh2YUWaRdoS3G9tB0QMEWCpm
MT2YXLJcGfrDIJpfdXxefCXBeYYoGvQsF5DgE6vFcgWtfMEGznvDotv0MWTT7U2Or/AxHgf4gNgG
GDI/X3dPccBCumeGE/8qeILN4SCMl+I5/uwpeEZEVMP5HVVCGJ5JwKaIsnEYEMNQkbW428qSWoIn
x9xsG5WT50xRlS32p/QoPTZk3LKrb+UMZnRw/iWYhCusuJz7vGqExlvHZsuHKiEsTdacd/2c32HG
yqbQc+HIpzViOiDJr5AOOMVnzc7ahSVxcH39Mg6LTB9tHlkWOGAnIO4SSBGBhYHjX9QdDoxU8AIt
qwTzrxNNAeAoWDSJDExV/vHEx2PjW1skUyRE3tLx8mMH03DMAvbR58j/fSPlFKFdr3E3ec3KGoyJ
FciKHlVObdV8t+evvocz4XgSWpFwgkfQvcnPqX6lFpvEXBGvn1LLejOxTtMhNGE/QHWq4rnL7p1D
1xq8e6IVjjGXRESIjDaxqJOLZhKMMUvkepIfrGbw6SEIsq0n9cVf+DCILpKb+vyTC4k3nQvh6KS5
+AC8f01vtaHefZx1CwhwAm4FuDkrz480yaMGQCZ9MizajWuXIq06/k0maIaq/uMc2AQadJ35v4VR
hb2W3THFUM3RdWBuLIC+ul5bLUbECRmQbOTY8fyYEZ/ypYxCMVN2rlfuqT0czFEedztJMBAbG6X7
82zi9V00ItRVJUFuOhejNP2bHuLxy+VNfFsrxNPrODxkW3WPm6xylEHW3sOI0O6c015KuRx7/2Wa
Nr5Hb+Nga7IU3QDhAfDFtCUJO6gvkRjHgxpsBBq55eDee4rmS7lQMr88A9/CKnt/PEvJ0Y0LJKV2
nnqSCUDQ43USgwIA+6NMSPxwG5yeOrcSObybaytGI1blKHNETczPjYALNoDwdI+PRUuc7K1CZcsO
dKQ2S3aXC81u8ofihOhGSjjFi5zRXD8yZ1MBWH3Dmf+t4pvw5vJ3kRHN0eCFcuugVPQhbUpgbjSv
KTFd9b3mMlr7kU5i3zLa/jc0DQEZROa+7s0W0iHz2OxWjJNbHH1/o8p87b4aZ3DLPQz7FhZD2P3U
33J+DUONdtQK0Iwaoevjxf97xDKyyCs8CM6osnlgeVgUURvpbD9qxOC6jSXwiPHcNq9rRFlQwIxY
1/Wz1S1muhz/yX3UeLK69dKMdaHuNT7UG/G4xkQxPVSNAqaU9urqXscCHDkfD4FXlG3vf7z8b6xT
CkVaFolpDtkPxA07YibpPT0lS2Mw9OqIi0qYtOWswG5qTYO4dA9u/VBivS6E/rIx3EvSrE1DeiH0
Zizy2n3hLkhR8QLE0WwpjF02Iq4swYpxim0bwP9TckWvSe76pYNQTukXN8jy8no1TaWLGkSBRY1q
pGGrdRkRsyFxyr6W/R3BW3OebmwfuTZUxy4BC5FjmAgSvxVCaCVoKMiL/xeXXdwxZLH0f1f27MOL
lqULYywZwZNc6F4nroyYMZBpjv1ds1S1ZLeLR90xBJutQb+rplE6sWAmmBptD+GE4V7Tsauthnhd
JPUs9oRziw4ARCTv28YPxu1zlyGYFxf0oVWXHV72R8QBJ4aq6ZdXWUmIIeUfvrD4x7/w+1vKZwnP
KyOqetnbpBgHCRgPA4nSX76LbAVW+M3d+va6PWpqo3HLnUgJti0C+GkwJ5n+6sX8eUe4lcsnEuEb
XzYPkRF+xAw4XSJoAdAYgYzHWCeIGRqfVMU5QL04PFaf/DZmCnmv8oekx2gl6f1j66vIbln6ktnl
2+iVsokk2voJ5ksGT4OPBgwO5uDHwWOI6N/xmoDWoOxGy5kJMWSZ9i0C3ilmn+QCndHglSNB/cFX
xW2LYAvCnQd8jDo0dRZfdIhyTSaJ7ncasGV6ldBkkI8aAYjaewiRLCkEowW1EYGojI7kzxQVq6O4
qpawGQwqOreiEWN6MXGPudLBsEXbboX2b4LhCb50DI91ON82MLEMWkBYcPJY3dd32jS0x9expDUx
J3PgnrwkZnuaSh0MLdEGengoVurNA3ZRwH3+m6NVxFauEhIEo0C/aNb4V3r8W3+1QAYV3/zqYVI1
mKUxOzqvxYdPKO4LbDEIsnziYfzPWowZ7lDPpKI+FeMtvxsu5Q8coziYoTFmoKvXVU9nA/U52igO
RHHl7cinHek8mpv1uqMcLF6g2kngUOSl4mGElLZmlEACeY1CGg2lanoYyjCs5Kzg514nRnfcobja
3cwA10SO4enDBaqgys0u2M54fe24nPLQ72jcJbsSyyoa4gMxPM2b2hhz1P8eBuZmP5p2KTEOJNIB
yOtwvfXktriTgoAnYBDOgO+T2uthoIEAkIKBwX8UqnR+QqzNo4IkGR3IJfpX3vXjBYpjuEcWUtsY
/UHMvpcKGUHQ+i+AhnRmrSfFkxNkPKnEGWgXyU6bi9ewtEMwXFV3y1Eip10fA2os+A/N2PRGLEFt
+jk3CE73ZAmNI4XlcOBqv43bcLbSVNEEEqn32TOC/YXAHUHs2KseKV7haYhgvW8eabANwexk3bnT
c9TCdLgarslfEpagtgW0I/cws9eb93qasaN3jI+xoyfhkMik6Z+N2UzZclYapuSQeoMswg9Z5TUL
l8Fa9KP0jlyg3POn5rthSttvllB729kAxXX/JLMyVmGyJrxKRjzIRsQ36QuQSYRne3QJDh+H2tID
FNjgf1lBaEt4cDdsbsx/fR/hw2Gst5R901ppo8DZaz56jlO7b3FSRXRfqhDxV5wrcuTTOndFBYCU
ya7+VRtVG5gAR9TGuus/7IMuXBoVRVjdqB7nevd8TvM+9NEIdKjjTkAphRiCatBBSGEMIVhXkWnZ
BgoScGSh8JDjD7jqJyD0WVtiw5BrXa3ZsmxV+Rf73U74ZVCZ9godMPOW5SagG+HQi84QX4o209Ts
YrKXQ5xmvYRiHDEDNMrUH9+J/VmHJ4KUy5Tv+IGx1KGFkNdIuD3PJU6ASU3QNNck/wA+J9JIlEEQ
3ev8oEOnsfoXCbuAxsENdl561nuF+pfx3GR2qXnjAFIa5ZbossT8llF0wJcZhpOUOs/VnbtFqVL/
aB7Gu+exFQ/NVHvvFpvmmJn1PpyIU9ihwRROlPeQw1BQBCV73U8wa2Uneibm5BSsctTOE72t6FqL
WGOJ/PvWKwPqxvTxXDrQ06bOtAIGsfmorVFeiHsD8XgTsbd/8cx8EeqiGifmiy24UVZn2cGbSjej
yJAxagTklVJBgNfgo29ta7JxV69n9VjP8RoEy+n6VA4KdhzfBJLdPmhBS4HwB6hFhLsU0BTp9Pyz
YkWDCOuDKxEV4FhqrazF713D5GDD5L3SB90erBWd5NMsuD3o/I7G07blSvV4W5a6g9b8voSWHkgD
rRRdz0c8WjT5zdkB7oMpj9/LZ8NDYiRz/Kc+9U8Mm4DGuqbM5blqsD/9gM290W6iJvN+3Rk6O/o8
YRIWdfQpcjV25/2dcUzDc2sf9cqWNxe6qic4uNalAnqk/vVamv50uMt95Lpwrk0qxIZeEOo4QtSy
qpOQGSTQV53IBdujNGOYNf11yAzgTPiPNLWIpPZN74a8zr18Pdd90O/v13k/75594acfzt25bakA
My+Yh0oBtNZcYIbOJ0ZNZJMivvjxem4NBGuixtjKEn9rkdq6oDTrKaiz+qxnnCWV/FN0cKqRzdzG
Gmu6iKRIjwfPBnpXvoWybkz4R7pVF3W473YovU/m2/pJWJZF8EagfsEFMcXxMyXGBhJvSv0frG92
y1WgGzCHY5Y55c5871AoNI7jPrXkN+EWvjejgKM1lPxlkbbF6xOIh4/WJQfJB7naRNiol3ndTT2C
3Ftp8ywkWuJu/G69DsgjJs95Vtm7YXXNXtePZ1DbNQdqPtmQv+5Hmw1l0UehCirmiXgnARE/yoig
ypfm/EpzM7M8BS891o6MQK1ekle7jKiDuHmTBUOd38qcfQulBvE9KqhZahgW/ZhjQKbAyaIm8k3H
HIEBR6ri/+ErDSss8cpAjsWJ3J4tPRMrjmVV8zNAEPRBj6cugtCe4X4AYyPXTegJCyDGjj+KCD/m
ZUd29Z3/H8qPye+wxOKS1fI/lmEZC6KwXPhQSmn9JvT21L6BIda5iCk9g4Tmmmw0GDL+6Q9YZNsi
B4jim7lFgmaD6VMuiqv11nIhihKqDrTY7dKkUQwBqOvonoJG6d/v5YsLYaBZpOxDimhXTdzO1HnH
KlTDp7Q10zksc72vZB5JVONZBsMxBFjTTRbliR42tunl/XJvve9MDdlXVNHi7zgTH6EzP/wR6wzJ
YV3vs+cy3W7Zm+cLgnu+9iyWgzjzU+dLu1PCoe2R3S4hPU6GOYAmfeMe9f2RKjRnlttVntBrpCI9
/61Z/tpRyxFzMvS1XcGyHinPh/RVJXPzQsFNsZi0Dx9j3nOo3251onKTUrM/K7KfTTwtmf7ilai8
sdwpYK89WPc9vom0dcwozBCDqvwjqiFGzMH/ZdvaQbM6GWlYb06T5+Uml0PWEndmvw2kHeucGIQ0
tBlchZN+uczv6YnhBg+TVVJ15DODUaAzcoz5pRwcqdDdYpEt7f8Ww/huTlkauS7NMrik+3sLZTVd
rl3EuF4+YicFGMoKf4utL6Q19amKeo4VMYgZ2k3mw2UOR8Djmp2inhFBPEBkvbaDWBvEe9MxXe2s
T1SetTcpQ5Q1Nld+zTjiyyjEQT2z3y2AVt4NHEtTQ3bss3Se32R36Ymc265W/hTEOTRhfwnQFhoX
6Tcdi3CBkhgaeboC/zmSevGbGde0pBitOzzQkSXkGIysDtsdBEbPUqlEAGWtwC/tpm1yaDmNObgH
sLNYlpCKIfiH+MeKg9tjH5F6Zzb3R1t08hLrtXDnQKimYcHBO51CLeNulyySzGPrWN41RYC3rlY8
ggmD7JMZMCgcyLCYRqZQPycFUP9pyQjseZ0EiioxIXNa8sPLYM+9B7RAbfYdVYuNcqlA60k6C4w1
B+5QMIsB8tjVMbyk3pARY7fqxaMrZTx94GcfIeEQJW+m5MlKYbFTj/sObLwLhCxGBXO1ubpmwDc9
QnfZPmdOGiTWP63XUFUJJPHPmZIn7tPf5gVcK4gcDj9s/Xsqm+QtrTkp+632CIzdHrgqjnKqm3Fn
sne/kMSefKw38v8QwcqQtwMPcBGe38woe9F/C8QqX6CVDS7ZUnGP3oh+o7s3vXoKul+fIAFDDC/e
Be86I6Lm6TKn4WZy2n947hoe5U05+tZJoXnHPr+k17m1OYbvEuy4DeFIXLZwCC6m767VE4vGpuSQ
cjIa6MnzYJGKkFpSuckesjeyY8yB1tbUgGNwEaObY3eeyEBMC+wqIWU/AFRY3XD7BpBL1QY5xZ0z
uwN8L+TciGtsxR/HYGaK4R8DBALTguFaLjvsHd6BNEw/gTpzqxsy0PCSYHalBwZG3ottKjS95P66
oPSdYv34QiosWhvGp/fQVa5MJ4PfH/xZ975MaTKWX6JarZeEggcAnWQvPRRfgR1aJ1RzSERI4eim
gJ7l+RaRzrUEcxVONhypj1ZMgG/72nRHA8QHqKj13tDiQnaVN2tSV8ZoRMb5EnqU4cS1ble3cxrx
9wn1PIJ7PmsTKo1oGJ5MhZm2XY1HPY+hAwxcHqYdlqPDkfqqvwKTdc/WYVXx+U0pgUaBCik00vYI
0CiKMVuSWuVD5Ehkjc6ZkRPO4bzmlPfRQw8I342OaldMKK0UAey1m6feEm7qKGtdyxRMXzn36JNf
u3l+J3CFEdZCE+bqCGJCdIL545P1cIGXXNhBmva1Ns46C2xk2uWYLjIs8ofrRFpAByCuoS/pN72b
Fz8EUmM8esfjLGtIlN/inDyAh15ubihnoA26SaansCuoSAAVpNEZO6tCepkNVf7XyujxVBGBUSUT
si07SpOBZ0prr8iXOmDeFBWaViIlnX/4dhL+HQtvM0DxxYFuNUgFU1P78q03+1Eyr4j7ogEcg7+f
jIjUKiZxUV12757Zwer+X0cdI44RNNkHgQ8GkfXhXjJMeGrcwz7UFaCNiVVmXudZ90TGP/oysesY
Y9ddS8rZAjrjeLaC0JHYesKM3JyF2BDb759Tq+X5sFSKVYIWWpzVPL9ZicAh9C6kFchykpuoINbA
oaGsBc+x0oIf2nmS5zPLxwMnHyw9ccJGgT/Aolbfr6cutKaeD3oWo33BKEuwdyfjo07WRawYWRLc
T4Bs7JJCqBiE27Ng8JDVpfNUXkGVTI8GgT4AB8BOmD+Jef/Q2zVHVNx6TjS0VE/AqwA5HSGs65hr
p2htLfkj84n3uMsacDCOcGQa/NLZrBpN+eW7RKXWQj5xlVdZnIlOWhn7fDzhYgwm7KnNWQsnJ/4r
StWYpchhU279uDhtOdUadomrfBIrzoawwAGU0HEzHGTBeq2VuYZdP5YrVNFiJQhvyUVHJdMmNvUe
16djnxgLY9dOTJDqx7i48VNO9LwuES4juJWWEp6RNdlMh9oNkPlrbvmg8cIrapSv8xuAUW6LOEDF
yMiixlkA6ymUmNmhBs1nhmcEe8XEaDzSScbjyguTn4mAtZeq8NC4d12/JJsiTL3IM+JAPbhZjQ4n
iaAGi98+ALI7SPmeHdZue9NZ7im2m7f542PDCsBNZshD3LPlXcIrBETTe159F3QUKQp9Calj7bfR
lA6xsVxLQCdwEg2bpsgZVsXjOS82PuR8LXDup5qAsTPI/qEJT4yDVG8dRkXm1ixch1FezYSuETHC
5kXAYz3ylcGCjB2doFByqSgEPAQKijq+KsAjeM50kLhRRh+Ww4k0VuU9I18Mjwqd+3nEXyfrHls0
lBoU99tRWp5mahdFQEJUZUEyfEsnE14VcepjwIuB07deNlbqAnJrbg6ZyAV8i3a05EdCu8v5+vhh
CaodkhL99Q5QmFKALCWFISiIKDPE+kUC88OI/ozCPSMA9hrev2i5uTECHuVaOejmYTdPItghRcPm
BI4iNO9eqO0JYtTCFOT4dw3qAAc97kXVH6Dk4gk9S8nQE7WZETgCeh7xqmYd45SRDnidyAZx3GJ0
NcWuT1m5VQ9al5zL2SIr1UHrVRfhYSSAfD3fSJ0pwI5lowcdcoOJi0Unyx7dR11xft3Y0xfiaKaX
1C9PJtqE3L5y/otTvR9o3UYVzMfIN+C5qEhLVRwECB1/6xJ0HGIYbMnWZZ/bLusJbvl1hUSMCYkt
2P+YV9lF/aImUyoZVMcmmITXqsGDp5iBe9cvZRi3OtftCATpCV+4ESpHL40Pkzj1mw9qsd8/maQb
ro8+y04NSp39BuhxxgCQ3oJxHyPq0dL9pMg0qxDihzx7bjU+MkS7q08BAd9IO32X/vxiGfRVe7Tm
MagysmZ+omLUqM9nxvTv+fs0y3irW8wDxcIzvzKtw1084pRwEr6415mqCsfNskdfjV9yp0XTRcwr
Av5buXFGSPD1Yz8gL8IKFhtQTnTP/gD1dPvGzEJoLkmbwIFH8Z+9s0T3v88XwAH2cG+jGt9lAjlk
HU+t2YDmL6UHyxTiMBBGEDoazmedea0iJELbhwp5brzWR7Zn/MLvoq1DiEelbmOz4fnWYFzUVU6k
yjT4cB4qMA+PjLt/6RO6RyTeh8GrqobdExq4JcYCfYqDppIlpYVrklrBm6Js99ColGcEoHvAaFaB
3/bA0rkPxT8uOFlCipFXfAM5pfR81+yWJleclXsHlNU/J9IO0+3NJXfudlgoueEjy7wu/k7SUa6k
vNAP1VZClr21yCEZ4Vpb2k33VoLrNF9RZsVauszC9H7ORqGsGOCpI9l+LwoGTG1JnDVPv8yzRHW6
L0mBuMhDl/J8e19t51CuDYAmDstsTEi4H6wB5Za7fVjJkff0OxBKZaEUpsanG/WoV9bvTI5ohtEL
QSIiIvdI9RY/fKrk9Q4Bri6+5E+H8RPuGkwthxGjxzDn+daeEdLeSmatmW+YiktaYTI7ecZXXcMn
bgijFhkIqKR7mrTQA2xCDgWHiOXvn6LXZYN6FQ0m4LxLgaK77VPRdpws4QYio3Nn1pGsunoH6QmJ
iIFOZGalgwCFRRYw5aq3L+BoW4DeZpbpLSNRuuswQCBgQFpfUNpq/xJcrSHtsvju42NeyqUdHB56
O51wIzo85mS6B4Mt+LiB233W9azFYs6STSwRvKEHHauJQ+INhTI22Ibf7A8ogVH7TUJeN+wXf9LO
sFN6wx/Vo5B6Ptb+g6mwrJ2pG8VSb0KgqAOA16uQ63qoHdKrg/kUMGZ3B47bO3NDt2QkP8pXFecu
w7Ia5/zcVJzakn8HPHeIi5n2Ev0UP4AswVxV2wDO9VHX7L4/4vlpkvXFLC9CdX+Pz0e9g+dtFw9E
MDaiQrBWRWRaZqCK+z2iZvxKb87El5bvHRRTCRSU4KmcIDqmrLrcLKoARtf1cVew0uRTPl0atQSJ
B65Q5OYX8m6k1Shnw6sTNuqOnuVD3JD6+4HY5q683MmSIEaBCyWgpRN6ly0JpnAMrtVpQKRb7uRk
LLLixtM2XgIguOxfZLwJqj/DKfb7milgNP3zeQKX6mU8GtJKu0XfNNyLL3X5WbHCNbUJM+IEAJoC
rWgy5wE1ibxrT8r2T4KcG1RSk3Rc4bMBZ8vT95ZmVyirjKIuQi86Wc4Ao4weC9WKc/VKlBbeqjb7
EVTcQWue4qUDwXzP4wtlDWurkc2FGwRV8qthyHMSjrXVY2hTqBKBcQ79vyHYDjU+2hedLKMXnIFG
9E+oXxekSDMiQY5jeVGh5LEU9eQ71J1lUDDQtjypXUczsfRb80cjWkl+aQ3gbRTdNb73qlUAsvEo
0MOPGr1gsEGg88hhvHVna6Tb2W11FIE93vZl4CG13sXkqYE92oGYdiJ3FXF6gW8xKYMTpiB6+Efp
T5i1rUFWtC4OxBJ3bwEvvYPKM+J+tzPfhih2pbvEhDHV6YFVQs5t3qlp1lgwdUk9n02i/oCr9Pda
vL0aT3ZOjipmgapShO7DT/Az+vmr80mLFVov0oZBl5OYTRESaFYuHMfbFmlHJPAWYgBlgf24WAhM
g0aRBqnXwwIlwRnVi4hM9asR++piMfeJVmAKMe7oO57iEVAJYhMr0f7GZBVOpRNXhPgah4VR07vQ
LIUXyQyUKTyD34Mh8bcuWtZEOG2pAmFXPnyEetNV+8Ob6xpMJaziKL0M4hOuhvmD4Ofo6fTWn877
zMISeOwWtA2GuPSslxPN1xhRGFwVIHqZPcQIYcZQHAxTfZ/uQJkrTS2f11Y0dSqA6NgfL2F8uSPO
2W5wgvMoUcwlpZgMJ9n4Bi280ZtB65/h+Jew1bF0IAPcTIFjdmeKWx5syLzTDxwZm2+kwElaAGE2
wACsKF+tU/KAQ2TgbVtbLIzCVP7RD7fmRoqFwtwLXqA3Bz031wyYSSJJS/VYQPLekE9jkz4YhXb8
jmbkPw/8pJXhXIwkuMM/1KAboJeI3/a/1qDnJASHWIfxYALoOg0ii+DzQsYxyOLCVPbkK0zTHWl+
+YiMe93xZYyXPjPgxoWNIqO2/lxy5JCoHe0AZZU9MAByfcGBC83qzew6Ikw1V6uMx9B1wobaH/yH
OLksWoeJfRnUaMgMMtrRnfcHsK0LbrSo55T4m8ZeAT7XujtfaY/FzoxdZj9NkV3GwRnaHnKrx27N
ttH3dKGNIyGnUW2AyLO8cBEsyjsOCP0Ys3Z85vz44kpYZrG0mslmmRV5WS0t9MJVRRLWzsotRTL1
re6pyUeOVv7W+aIRqUMAVE9sisJCS8swVpxq0e5/JEXSECjjdt9TJoI0B0jNElToRKMYN8KS8Di9
Yyv3fm3BTi+SQzYSuQ8/K5lN20ADAb6I+0uLO5t8bcDIu4dRT9bMXH5hdb/wSaefkfxoIuWZHn5r
lqziMuyBiSiQC2zXtad1s6uj1dVnnz2amUQrag4IrICnxN8lt+BrVeUimYY6QKF5fAlgvWzG8lUT
SfybVW/nSCZreDknEu02IN5JTJfjOPXjFj6E2VbMZcmCq+zPqpIrrYG+VN6l2Z2om2hQEQ8wBhfD
2XdpNM+wJQkp2RQPR+Ppyg/oI15DAtKVrOtQ+l0KZ75BYDgsRHccxwrIGvkoJEJ5jYkRmN0rSNKB
pbfcXkzpbnh5YYfh9/I0zTOevPXOfShSXzOC404GQOvRPrfuZJyb8rI2bmka4ic6NULONhu6uQYp
LLIhN3hWpZ41ZBC45HP/fNQ+24E20w5qyxa6S4B2xkdqXiuxAuqt1mkpuy7PlzLAq5asBm+yo/bM
R77GUErZxc2Sbc/CsYgqBUzNd+MM4xkpV0Ea2kOteWrgmUZRrIGaPY4bxGBH52AQi+xMhjlGqIDu
vKq5QLfxGV7LDjrK8wDVnoRed3duQU0Yze1a0kfB/oqxjANdvKDFQT9aZmAk+QxJJP9cuKkXVWat
xSQ7ugWAuDrzy39lUDX/ad1z0yjuu9lc1ZJRpwB+pvDRdc6DPM94OE5oZ0il9qYbfq2n8pXf4KI0
+0LyL4uTTHJbNKKti1giKU6zOv9HrY+Ks/bbVq+qANNMBE0u1f9f6VUAzdnY8yzn3sZAtwrNZvK+
VGvLZz1+wLra2F25MHFvZQep9VF0xJpSpvRm6t7qZiJR7tKkg0YR5f9BrIUqFkQhg0ltlAbnYkil
H+fg7idhxNYpY5Pfxai+3ZKaeI9mTCAQYeVXat4oxaFhZ5Y9z38NyVMACe1spBxIMOjxXXN/Ujbd
Aytd0xTft6XrFf85ag6scbKn7OZ+HXJff/YCzyzlunMXXeVnz7568KmI/1GcdJEpCdKCnCUf1xQ3
fq3CynmFmSS88BrVFL2tm8lyGbfben9ZtqYtbBMzSBji0HE0w4o/CvJCifPOZkH0mxWzHKuzSJiD
Y6T9WRA5ZXZD7ymuUT7ldwm9+S7VfRzfiJVQkL3eZee9K44MwRlCZ468hxfu+pRKheAptUetH+RQ
YkivoPSqMCU/P8zZEMCLhuEutFKBSMqoc7ZS2VbbADPgJCENROEHQugVc1qcb3K9HoqjaFD/P+jp
8BhDg01fRgVUqybubRBu61khAWoT0Pkogss9ciGccx/2IchHPSdsTwoe/jC8sLcbnbboOMfogrD5
XWpuWM60glSLFdewloY8sfhsfZsnI66tfsN5wdTdbTdSlmkUZxEbdZ2ofxGrJy7mG4iQUwQb/I+w
ogBoq+8OeCTGTDgS+56i3sA2Vk/xQuRhgUYs8tNRStN6d+gkVzQ5QMf1joA2p3jnsw4De3PQ4ses
gmfyvJ84IcSYZacRr3eSIuNGFWS4bPPYVbSwEm2YLeEah58pFRoJpids8KpK+kPII95Ci4b8cmEC
rCbVZQmWE7yfXkqTHiM8oQn0yswrqgWPAe+mCdrSGNo/1vp2BzuKbRcISnqvI5gDETjMni5BRCAd
USVBrOB7FDZmgRG1WvKjkWEGcOAUy5IulwmeRLZ2s8uxKapc5Ht2q+zLZvTCxbjOeXKlR7iTowMn
QVQcCLPVIznrcIZ8IF5rGEl7ZDWayny+Ole1AFnsDFdisFrDYNcH+rFlp3X0EBxY+B54YR0F3D/v
Yh14W/CdraP+iwQmfmvg2ER+SDjsryefxdB1rfxhD5yhzNXoBrChUfNui3c4uidvuT05m/OhNZjW
Rp6c2mVp5J/04eA//Ql9TNC4K2kr+SkOP34YbA7cmFlE4PB/GAWNIGIOusmn8KYYgIrEfBi2evQk
yi4/1MtkT5cWwEP/QlI22zoZztoWvmjnTB8LhP9662DbmW2Nh51mmCEOrI9F6gZjXgPtwJKs0io2
KS2ZEgIA646S9e3rjXsKVm7apX5V0to7QyIwZVrAN3zJSSpupZpngPAQK0FykcaE8D2x8z0J7YYz
K2WB8097DI4Xe55o/GD3tcqJS26cUFyGXs5+n3W4tMPXbiOORxqmdKtqWPyuWSLQeJ/Ntj2NjpA4
bHvK44SBLxJiesYLV4MCe0TapCdkkkH45wcHRbLmupCrtFIZNQm26eYQjn2g31VAjNa5KbLPxfuU
tSyt8pc3GfgrV+o9YlvpxqqU85biqf4zJXZaaVglteSVe/wk0HyBzmWJDCs+v2xWBOIpMvxg9cNM
juGXO7dzH0xpLa4CMMkhyOxblbE81KxBDd3KAuwSNPdIDe7qVonEEyri0Kc4JcHqt46DbYhUfqzb
R0AOg7YgKHSGpO5B0h0Gi8VWTWkeKa1TpaYDLw4ntUT7DPSgQK6ZOprrrTFlkg6eJT0s/RcV150y
y6r3C0EuCF77Ps4gmQeR64RnAkzkko9wk3zig5Uign4+NulPkenOrO4fyqu9Zwq4s9p3SCt+guqR
ue1lrZcgc4O8DmYmfE11DAQKwLU6UCE1eFnQgFhylbrNneqL0pjVYDzlaSn6AhaXUn0IoFa2y9ZF
ypiPlG0VUjnbitJeY/vuP1WkgiovbwGrONC9lAfOZ6G2N1U=
`protect end_protected
