`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
SuCYZDjXbCwBqdL1vAOG3qslFas0K4dFvgPZbrJAecEne0gvgu7DcL7RWU2R9hQK7ZzR65AV91YY
a0N6Qh6O8ZT2uWmE24ZtaRmc/K5dujRjVWXszLy7UvDIWfRUX6gYEdK89t21hUvH8sXnSFm3ujvS
yywdIpJimPiKH0CGS99Lr6RvpzQKD1zD9fuNMglCzyKOd40A3eu/aBigFTmjPkqoNSogJmLcLtGl
svLaElPDKk4N5eF+GzXeDkFC+9EEL+j6W64ugSWWwOeGAp+2XvxwSRwmlk5GvjqQKPy1wJYrAX2A
V7FhHlBedAWP61YX+UkElrOyYs2i7RhPCBKzCw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="9uuZk5Xcsve8Juo4r4YO3PwntZ2ZNj53IXzYU626/Do="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30112)
`protect data_block
XwAN9LZY1q2/NpEyIJcBdxzOgb4sTYiDJwurJohZVE5yAKDMVCznWOn7ZYIcd16/Ct5Z7ogJ0PGa
xxb3VlchMqWwz37KJGI6ws42oJkwIhOM4IP7O3vUi+5o3Ug9Asf4YsNKm+sTAgzBVU4F2okLMVtZ
5qFCRyJpiK1NaLQvEh5FrfNDWVRa48yCH9WVEs//HYXqYyCk13ZK+mGYtuE3K4tRakhgGvun0XYs
rOON2Ma3TECwrG3MLiFZXOxR+bKQNLMEp/8XgHY1BFuonEhIt5L79Q1M90rfFfow4B9CODn1lJ26
14+wICGlTGjKxNHIiGoReLoCBWGzffsvS6gQN0Twm182TMcZYsTFULaG8Cxc8uH3K7akJA3LEOan
QN9hlkzhZQxFnOiNTsrDkkjAHKwnx/0LZXkZeo/56MJKiTQLpZxsq1ouKpTbymubij+FNLDaY4zt
0HMvCrRIgmUPPWci6/PmJO51M99DZkgAXZFFS/KRiRvQFt3nGQQaRiKxw8rdB41h66rrtmHeoRE7
mnRPkfWnxm3yUIwPFf0J8fwFe4X/xnSWu5c7cqR2xJTkdNLMa8GZjGfRWRDypezcr780AjOsr25I
9IUScm0O7vyM6habRZZmm2iuygZwkyPrLCdeqjtVQ5JkeplXTNtUY/OYIEYdun0FuwvKr3IdFiw3
xZqs93d4TNr5TernRKGF2UniLLHzUoAb7uEUNhAj7qvzNgfLoW849hDN20y55TeAyvXq+eYUMSM+
H3SA8qIqM//BP3AosMnKeqLbXP3ffBgy4DuamhmWMUJ8y8qyrS6HemU4Qm6XSl4MjHYM3UDx6bcj
tDeG0w7Zi73WCZ2BjCarTLPCjIqahSztlBcn20rfZJfBETiMDLhQHP93SZgb9OLDUov2WR231hvq
PJq9zLMi4xmN93vi2IoGOnenqULbN/WSM2/ynYO6knje5dpO7/UprZQRbLRA9lMGWTYxd1uCOzgv
KbQbAMbjoDyXqF+C4qJbMvX2sVpVvXfSE4tK7UXx/RYh3+GfVKD38yxFoIPG80kPlaafWzroJBjj
WRMoKG/XmvPjtWUZr8IbyLRFFOjCg9vpkJkQwTtHncBEu1zSBrpN87XRsCD96PIlJa5Xh/tnVegJ
jGuSyYC7cOVEOR/brEcnogzcLaCAEWX1y8A1vnx6oIIbLkIeMpJ3QdcUvy/0ihqtUukf/RfZKzG0
iGrnAq82H/6W5KdSdQfvAnl5mEgIM/xv2Gv8X1JBlozCe2I83WLel+zyjUWGAD2uqjMs6a0RWhZs
pa8H+LXuNyDHsRIz9pga9G/zJzjz5LbzR6mWpcC6sGlyQX0hANOGZtnbSQ/tJN78fg2bV1b/wj05
bEMmsI6d/upUCvLAN2SMEcyNJhnOXv+MHFR1+mrYCZglWX/CrC9emvrliVvtWrk93SLfsvA72jiL
p/+rDctXMFsQnLXCWMPJBeLnM1OCHSfZb0N8nfFdpEtUDDHRIrWOvfslvjUR4igejgq9mapOP3RK
qvil1I1k418x3/oY2mmyWl7dsvYQPYnHHu+faVBXH4vVYa1D8ZsZynyEmoqQGYQwyOwhrrOh8rOV
/rTG8rU5oAnLsMx+5q+gp78SdvDVUfWUzo4389gE2dgiREbnnSJmC8Oy0rDrfFoH1KgcqVY1sqNY
v7dmeOw39RBUwdTtHe3P7dMVSvOcUB5MiNOGRIwJtYrBgLpIg+woVH2s9qObIs9yV97tNGnZBJNI
I4iMgWaskgOfUf7iHJ5D3J+DWtY76dfuKA+KhVgXc/eF+lu8/xg6s4dnEYtuIYFJR90Q/vG+MY3X
DG5Wf8C5miPJGVJQtRIn6496AI0rKQzl1sAB9CT1U0gXuuaVpxBumff76dypODE8wsmD9Nzxa/6C
ApjVyArQwmCAgRzRuqkrD8Znm8pAZD1Z1ioRMouCYNb0YA5w7tH2lqTt9Xi2VAMosrAPBXl4rTO3
Gk+XTNgITJnf6zqaSw04/Jz+7KIAxmPZ7Ma/mhClkpn2sWN1I+cjMIo6tR0pdwVWhPnFMGsMZihh
PCJMqrReTVIVlF03gRgyVa+thOLfLgLsfSvziXkN8PtBtY8TO6WqunpkroqPR+3bbIaszoEsXWMt
1+XZn+iaV4D+vjS6CVLR48okxLDf+II0cfmF+wayx6h0h1O9FOBZAjXc/rICHrUY9kbGUsWrFbIs
upo6mUQsVEILyKltOrSE4urD/7XqsjhmvcKOJKIPtMcjGRL7Vyy/mZjbb6AcP7+PDDobnrumnpuX
v9vTHHtr7C9TLUmxgKezy5jwHe9V+7kkZNHs7NsZuu5zW+gh4YaJVb6go7FL6+YAhx69MMteSdOF
EvA3ZtAUZfWITxo7dwMm+pdAzsqsqLWhMyHzIKkOMo5xcKXjoClgCaK1/OuZBBSIB/qbxiKqRKls
xC/wtNTbKUuoENmy4G0OvXDaMWyHJpDAHY1CE9ihrWi3O3MobtEdxDfBOjlDi7tlDboLHqAMdyGt
WQFY+k6zxUkMKHk8vt/8Dc0//zdqzdVoddbiHjtjD3FN14pdOKNMnatQ72IVo6232uuUeEU/luVs
R99TuuQlVdVh4ywgK41cOFnn2O/PTOoGLciCodJAabu6KFvidMhJ6nqCXcOLAMQ7HxeGwWwzft5Z
DaGtZAJ7VLQBpJYNGho4iwHpeLzmR2wFksfgLch7m54cjOFJmcI8JgmiIDOGIuwZSG57SufP4Ayl
mjvEZi9Xd3oDyDMIw+5i0aAYyGaBpOMbY0dd2uUKqPFtYOZE8LQWhpM0u7PVmqRj7O/4SO+xGnXU
kmyMt+dVWCywe1fpOCgyd2+Vx4/QpgTFo6+6ecIS0rWuwVt+RSnmp9rOri1TjnD68HJv73Y0rUN5
jpglmvxsvclglWIJyYN8rg1mJg4Mzi9O0447QVGmyvboANt2YwXlGiWENXcgrVE3Ab7L0i3j1zmM
20Dqx8njPXctsstcfZEew+YCShFVuJdWUnAMnYv/GUnBYh46fq6Qi91CmyH4YZcbagHc4VNY6d4w
xlPuHrv7DD92qSaZ65E5FyCT9enphF8l134BOdVbl3AHxy6o6XbxujxsepFiG+BEu7gzPnjlgb53
Y2hiFeVmk8CKvO8qLLcCX+NmU2HWTr1eALFpjd9LQMqjIzs9jv3qhdBFRhLiPzlcmoRx/wlLXgym
LFGWiqrpBaJLNnURyvpnCzhWbKI5cX5xGYll6zHg7XpqejNCu8Xa5KGZo93XN184UhMnIq2SmQ0b
UVlPA0+2CX/fuXJn0WjYASf2ncLv3drges0ai2DADVUH9zql60Rw5mUbXs9myzpo8pr5cOBZ156d
r5beCeDgM3keg16Hvh3iETO5upQ4C4Bebxf/3yQeLKE1PSp6P1IGCrmPwPYbEuGDNoOWlcW2tF1J
ZxfRTAZWw+Wc1E/7VxUGURXIxW76YAohYmEfxrzru8hsYS7WF8d21KL4MnE7Ah4ngq27ovjfHd9h
Qp0q0QqdOWX5pNnlPF/ErT2O05UniCcuZqftBO44pwe75qow5kWf7T1A/BpzAvGV8tjHhGYEB0VW
0V3QO6vrqGDmIxiUn7bL+h/HCNyByY4Gfiv3ooAeM3nZxvkL0tMwpGJTaLCrN12xRordtZCWWXcM
jhp2wp6Ml9EWslrDzsBFRmv1k615YbChQKnriNZwFE/3WhODZJ1sBnlF2ZJ7NHWgQ9S/qlxp/jVJ
BAmoWcFy5MWbGA0zC/dzQSJNtldyOH3mkgW2EQVHWJ/zz8ZGmG6vfPDHF47CncoKTibnAFTv11pE
S28RowRnQ97a9GFz8L2Nf3WQBryPXsCG9uiSmFNI7F9qsROtgHOvGdRXwLHwJ2sSNx5I6WgmGs4u
JyoVciwFWnky72Ft8IZd/k5BQ9LoD61HbF70GYg316Mfz9EIYdzeAuF6quWBkOXMdZY8CxfH0Zu1
yZFg+sGaHWFcFwXAr/sSZbHqMluX3pXiOsfkvMGte9gdhNTGnCHTP6b1BMYKsj1uFRVuBJqw4Nxd
e78RrdVZYHQDVryeJvdT+mnclICNpJaXs9hWkeVrt23WC+cFx42N9Z/q75i+pqaIfVpJQMMu8JT2
nPChsyigVfoUzc9Bc+6J9EhMBYus4rZUXzTektd2odR5Bk+jaag/kPtrALyh3jJoHcUfn1w043uJ
5nj/1gTdyPNkNlB1qBenDWK4PmxkxtCuv7hUA36PGZHzLtsRcmAJl9yPIbY3jpa+AtjkzxeuzZVj
Ye5RkyXpNXTDOSvIZXpRPNoKuyW3hbPWWjS+sWxnTBvSBJokxhkx6Dkz+SBr4Wl2reYvIegmg38I
IpRgXE7Qm6I/GwZd8i61MWtMj6i7+PEmLnlwW/8UngwHvcNXw8L0umra7Gf1N5UU+qGeteRkp+Ot
Kertaf2abJkKfcd6TLSMmIGj9P8Mtry/RF/M8n9UxpOrgougkgysMpp+WNVZdX2eKqFpF2ZSR4W7
96abD9oJvibygqnNld+LN747m0J3cHi/+lDaNtPwbwQbxqd+qQu4gRa+kImnACbfVBTWs0bVnwcn
VbBjjSPPUYLJt+6UpvT4w+TRq/3D+mdS8o3go6409JI3XImXbpkmY8CN6pxem+KYVAgFcJu0kVYw
JIJQna2NjUEWtkCrImMIa49iAcuh5FBuU92iQswm6FTFwQsk0nRNLJzPDRNAillAURu22T7ifKvW
zN3bOMlm15O3ldhB02pKa0Tz5dVUUk5pto/T5b/Bt712P3mtLNSrQwsvq70MM6pyGd8mL8G5YJwA
UqI0WQfK4721cnp6lYcRzpv1TFJgty4ShQyNhOK0Gooy72mGnHF/8HRl4Cm0osKk6PGztz8Km5Pu
1GPDDxAhd1VZ7qYWyr4msCT472qsCvT8iEg1IFSpzWf14pGHJ5MbK00oSdnbbv5lJGn30ZmjaTZ8
pPqewjlyqlFwqgjdynZG18GiIZgAUy3GwJKZwj7kBXdQd57RlquVGhrilNTpeW/Qef65Y0lKqu8f
PPcmQ+e7YKS5l9j1Rc86fEAy3mweNzCnrmEm/rP6Ud9nQ7zryEPvBdmfdviZr7zWIa/X+L+VDb1E
YF2b/im7kSiFOsiI83F/4uriA6bkS++89Avkpg8on2zdWgx9V1Yu3h77jgmYvaTMJivkamvBEhYb
Zztrej348U/w205piRmUw4NMmyscNQQm0usUi/oIHYQbV+WxbFE1z5s9qGMmPohOPOBRJghtmUTo
7+sEW1yNJQlw2HMjRQs5pEigHWF2PEodsC1mQw2SZ80+8kzRWo8R1BhhmEGVKX4yX72MNKgs7i5V
wSoqg2pGKKopW0DO7q8fxKt/LC7djdPMQuR0TkpXWpcKJitidSXfuGzgMvPPS+TZ2s2Vn0N0+KK9
BPsVGhBS7dQye/xX43sPgmBmU55s1pNqP/6ct9ofoBBEApZKMcJlBU52Jbos8VGKFOx8bYd4YwNF
r8igSRRqJF/FyIYMupeusocnG+B5EPP66RC29e8jn9X3Xz9XqbXLmL7rirX7hAVoQ5Iswcb1ijRo
Ao0/fdZZT2+Ztu61s4k5qqUhLazGtOCsxBg1UCxNnUiNtrMM84dAEPQ1/hJ75Xd1ggon8q5b2POT
k99DoafwSgS63CHblTlXTlqwIpgST7XpMudGUyyrSd4mseL/GkErMRcOwCIOd4RIqelZ/v+L+AfF
Ar8kYALdEJkd+vnvKymNB7o7erWy4We9M8OKtLMJEwTAzI9x948IKlXcJLMqh1dok8xmMtGx+AWp
GsRaOe8akm7nvowowvDNa9xKL6LoFBv13j+8JEXki0x653l5IQqb8zzZDUES71OsoOAaJaUkj3lr
ErOrlxofhBbrHA9MvCBF2CHT1MN+ImxG0sV+sKXLEM3W1zZHyQs829sLt2Bkp8KPRvbb2OmOlcta
M6KXVjTLjKeEZhI/BOtm0efsrN82Z9fwPraEY3zT2WixgTf6nQgTW0AOGZG+s+iqDqzvghW3F6fx
9iyAQu6OhItuKq6VMV+chaEAohy/QHIY7awml4bFxkYgTU99ZHdoexSamEnooqBI1AqrwLbZDhAx
ObUe+U0ortsCaSGa5NLJzg0MpQawqKGAZS+xmsD5yImPS90F6q9AYOT/XwtDR3RhEkRim8t4COS4
D8JfD+kT28nLmHMDoQLLRHeGBMUki+7EgdksSlkutaR4MgA/ZFKAllzJm7ORmUJj2LV5vKqs1+zc
cGRI8lvKK4UpVF8cZtzyPV/p5DW9hLAAmUNuWL2mb+hc4dqmu4R0o1Jnhh5nKRdD3f5+ZsmH+m3w
368uEKd/qAMmIsYl+FCC/kN8M2sOIHgeGFcRHvwrycZCit2f+Mk5690HOJBc/Hn3AXb9Px7rTfq+
vJQP9ACHxPzZ9YiPMsyOT3CQkLfsqnvx12GD7uKWIwj2anV0+OKy6cMsQ90R5y+Simoh1KIZmG2s
0puLf7vi9FN97YWoFnql3EAAd/b0j7On2nI2NdoMQgC5wwpu1Xd5YL4kSCIvdrEce0T9cybiciUu
0rhpQNgcdBD8Xm7c3+iI+IIQiX8e73NrcmH1o6v/wktcoJKoPcYozWykOJn7+5XwXdT0mrzHIm3y
B3PcxjAlZHIGiiaruT1SflW1b/O4PsDCCZggb2ytZoT5JFWzspwNhQpc6/qmhCCT/UvLnSjlwWC3
HHkOGaL+icniR/FoclNGKMwoJZ57jCCNX+aEkkSQch/Q8sq+9zuPCiFqVYy7sxwTWDIMQLz7nm4F
X0Uw7hGrxo6KRVQYxUVRYv3tkqeI+X6bFWlZkqDxr8tx6ECZS5B5TrPa2cFEVTQMuKANHnpD1M9r
BDOl7yUYYFuqMkmODbvk2Ul3hmn4emfTqijIk76iJY+EcVG9LlXlzyJBKrpXTp3i++HMmm7mz/ax
HJvzPCEOTkLC6Hun4a2Oz3zKib7SXUXmNpPjblPU0U64rqphmcGEV/8Iy5AnZNuDrpi9KUg9FXA7
/52jdJ/MhwbaIzcwln9dx4VgF8Zfq9P6+kwxRfz8SwQjl7+pWSiseNNnbMLG2W1ZHwMUahmBnOpf
VKW+ysiTdvY0sfvAMmuvHgwAHNdkv8Vmbg/ovIx8FJ7Dhp2vLzGNZewKFu26mxxMQJ8W5Zu7yuX3
kMBTGFacbO1hAj2CXZOI5EcdoOmgo8lBzgURGgLYC8gThxI7fherk3bCH6QNsk6ghj4cHUl5foAP
rAV1Hs0AvtqvOz58r4JPsgp5mHmn7bkN5EllE2twsUc9k0IQPruB1EZAKILxHLWC56xpn3PIWEeT
xN/92C2knjvaFb1lnkmhzuiYsn/3Sr8DTz0+/h1nUofo2DcK9Xj9QwE1lQ+panV35lX79NZB2wG9
H4TR+pfHyIJuq0CNCakGPWqcbcrnwp24Q84USYG+QXZOT8npY+0x9BlG14NXu11u4JCKA4Qn8ell
6L+DPy7A0h2sQj6J5vw/fDlzmeuBiiYUIHn9Xhv+ZA1CqrF/guhRd0mtBZWWTJekq4ryoXq5wfxX
SpsgkO9/ChjWX/lfQY4p0VT2orrxk48lX7/c+dRsY1mGKvJw55jMJZhtYRn5Oggd5APWI7czZ1Vz
eHuJNZUzfDPFuhLR8Vt8e/ZRSgUbND5dkwveB8nnrUqcdaZSpIHgoUhGpi/MOxh4jMjmzqa5/CYJ
xIsJ1dT2JSvEk4u/NvR5ZsnspXerOGcsYw9s3QL5JhYJ6JlDib/hcIJmwVrro8lKg01rqMQqXLci
+V2CnwRkeKAoSUW47iwpr8FlnRZ+TcqD7rmPYo3NGjuZ4UEoW5k8lcyruCk6ALIR0OTcU546lMdZ
QRhfGjkwHZk8hdOVF+z1RqCd+cLrrpoWaL+37VDRZHKbbSpmW+jJTrevJK2UE1JMlo2pL/j88qJN
1ygUr+tL05zN54VEBmaEWhakqTOLAcWDGP89jFNwifp72F1lT03H1aPZ3s8mpwOVoG0UKE4vrb0Z
KwD8LDsofnHvk88eKTi/qfRNKfRYjwwQA4z4AsGiKRJIm0jWYpuA4VoC4+Tv/xl9mxKWj2BiCVbK
qi0JwulnJKIXg9vSlT9TMXJXtUOZFg6EhxdbZ2SClD1zzrOUxfB28t+6wqooqK4dA4oGnAhkedal
hsnMggi6+MIfnSrc7R0YqDqacE+JiR3dYJMU55lMWrYZAN15YT9yvMRLu3ggGo4WhOiZXdwF6q5b
vpuNynal0oPxIovfk05qLR01ZbpjmxPRYL0ZACZpGIzAYNtpqs/9qlwErLlEAObrPvPlCvHfbeb3
qvKTCu0VUBMkS1mJX/gmzaQhiJ3WcvDtH+xkxtXFBUVkoVaiQf2GAthzU1t5DKQFnuHEm+fUWvRF
AD+JDNJ0S1N13BUil/u2/Yl+0/sZj2X2AcBlkkWBwf17a4b1zTQqsYZOkL2JgKsQHxajEzK+/fje
EO8s73vM2r7xPjCakUhq3iwtIJ+d3/g7AtWzXk9irK9hF1ROmpne5hgD4Cd6xKIdTzKsuM8mllnd
akLCvJk4PpjVVFCRgMdEaYogbXP5Acd0ppdw5qfbRyFOxUpZNT0oQKTsCqXrlfwGUem+M8RvUZgI
VlSz5Fx7P0knnHCLtRqRn9BgBxvD7+EgPT8aGgWxCDpJ6vEgBcJSQZQkq9CC5ciKnUHF1sFkSs93
rEyo3eIdGL6z1Zc9rorSjBO4cFH8+Bgvb9HqU//iaqPYIS8ll2L1TJ9+SkQ3sMVZsc0WIIGfWYbq
XrEgn47fwaFpT+mNdDQOQOTm6Dy2Xndk0uKXFZNMRlCTtI8lm5td6Y39++3c2INi51y7XUUmQwqm
h02R/i/cf+ez3V2ZtFZnb9TfW9JlBOU7dc2aRf8ld0Y0mx0lMA/J9TrzffH7ASGe/tKRoT7HsaEQ
1rWV+9f+64zgKIyPosjaBhRtIzT+EU5stYHL19dIe5v8U4tNCAuQjvDGx8Qp65ZqDhIammbGy3h2
l2QUYwwkLPgl+UfA7kJvsUo6Nza+cDE+DVA6Q+gxStqYyLSa91+5r23O0dtNYOkFHIBBfgNEXCF0
caO8ZKESlgtMFeLEJo79/Eb2VfTxsRCVwMrnpk9zbTMHqsR9S/13ESr3RP1Zg/P9b9n8JdrZ0uJt
GrOB+c1D6eImc7bFWzfkgTPw1gAOyDOZJ8ICMOMc7D2y5JWWfpGUCQtjtNqjLkpcU5X4c6WpF1rB
ceE3Trs7GFasUqeczS/Upu1VR+vKeQ2IIpkndCMD2n6hebGVJtymRjK2n/Rjp7IJWdZQ0ZLHYoPl
O+cNXIBgfiTAVxHt0WK3ikggWg7BEDqDbkZkDHVjF83aE67WE5XI/lffwap9Xn/lYWicr/GIddI1
UwSg5jWwrk+y1YqCUcqQF9vReLIzO9J8rvHTu940lxuRNhiasZuXRhCWSSHW5G2rA0UuV2G7Mgdu
n3NXs8h8Bcl35XKigQRCit0zOXMDHb0p86vMF3QzRVsZQef4sGx9lTLeNi9kzrU0SSu/ppq/5qS0
o0CSnHJ1LLLiNYv0uLkMakrcAaZMihr3FyibMol5Dx5nc4y17/lolqPbEuvpzJJ79B4cgIscrS27
D8mIwVzMLx81tggek8OLJQg6bXtQktSzcJFnn0lws6M70g1tvTA2euBHlN/z09Gu1kDz8cPW4gNQ
EwTF3/y10KphdAm73R4KFl5uDFicc6wJveuiWLwPVV74Z0LEHEZxAI6ctExAdNcWo36NNAZaQiHV
vGvx1sCgYy3izu5hTZkWThuRKr2k6Em/Nt0l99gEcdEwpQBUg/8HWdAwYmOp0dudkVyCK6B8S8jr
Jly/6U71dv6X0MATEdd+JyCZ5gACH3C4W/34YcU859vyvsV+CkqTZ44wAwAyVkn5EZNrgZh6SoUl
WiGJCUX+S4xza9e2OTbU9SISIdHL7bxTU3OKhRsfEXeQuhHwfsT7HO9btV2+EbkZaOCpLf5tlVwN
XCY75rKlDmjrmOy13am7Vo92cAYD+YmU/sfmHLIZDuvKu9rSp+3dnKZ4gK6JxhCx5dLzui1L2B/L
ybhGIvvHYghiiHv3KQht6iiibnOOVlNsIO3CyV0wvBf9BLEVzFp6hLv5HoBsvhNcpXpeqmGiimuk
W4JgZJD8BlfSVHyxnoR90uPUtAWY0zB3/w9Qg6yB1Pi77qFYpApzbamoY1yuosveu2XEL0aY9VoD
tGkMaFBpxHYyjIuX58z27Yrn4sNsXhJlGr4TKpAe3HVeQyvmtwPJe6CY4Fktq1R5pedpa01CbLfk
9xvdMBx4dRYPvEeIN4aqvfdLs0Y4ttNR8zCIo+Dg7PDd6zxCtpXJJmL8MdgoVnbUDTIXpKgdf6Q2
Y6kZUMiJNgQ3G9fxNotfRRNgs9IoT5xhunf6BhkpaOSgUs3Wc8VOTpoI0x9xmpC2XbhEzLCAtaze
t3QZ3fGnpqe4rKTzAguYdgFVM9EEnbVVF4y/1yhWZtAgt5UO63wT/vvunpuMIKteMnd5sf6uM53l
BReLyLznuSjpucfCzKnEI38BRjhMTkFhuCn6oFNB42xrI6oIwCw+jJBOzvmnAeOZgVJtopdzuWtA
qV8NKxLtNoO1iUOIGi/Xs7OA+cy1UnsZxqGiFO4fTkFJDMv94BWyfv2JDOlLbB1IT4u7bGk8sRhn
cT2IgdJM8LfHvLnCKHX21zC9VLZImXb2HM5IvxO+8ilc8GsUj2aqrnlbtemmVvPW9u1aMPA0R7J5
ZHaDDjFvV93p1k6nWrKuzmMSVRjulC2yuSDG//xkmkADxUH96LOwJYZS4hRgV42QUWqKNNqaKCHQ
rFZ96id3INBZvwamwQQI5c2JviMdBLobTJrniybJ7NAzKIKeciX3iyxq9i3p4iYj43Cdtq3JC0AQ
xtHRHg+bRzjZ32C4kIJriAJm7H5GbcivtlGbhGs3Xx5MzVmfovBfjzGkMZ5fWoRTdnP6Q4KZZk+G
06mTUmUEEXsSBOOE9QqP2gP8BNQqCLyTwYH8DNqCwtV2IzjByhMVOy8EVEQgmIaa83eyhmgIZkP+
lacfV9cHNJjDtIosq0z2X1O2m5yVihORAq90jSgo0N64AI9PrZ6gf/4IZVURTeEzfe/w6nDXLihZ
Mw5MHAHZzIlP+uwrlcZFy4NWbhZtbE9J+/h6Es4Ouj/0z+TAeS5hrjBG3I0PbxwXspENbwh4VJWT
jq+9IbWKIXdrj/wH945S33eShGh0IjcuMBUX3o+kzPevo7OzgQKPKymxcaeEWVXxc+MGsN7AYmOo
ucvu9vu0QbJtA1tTkpLL93ny5gcjVkzQnk23m+pTM4gATcldSeURsdUhTd0507zBcuKFy0PV8lpd
8hi4g7u0BcmY0gByhZAuIoNVylt6YO4Ke2KLB13vDuwk9/kjJTu3Wwqv2fRv8hRuT5YuhcB/2aeL
xKnpKIXQHx9nBf2Efdmgj/kJQAdROgQxcMvfyjknQxQ1voU/I+h42VEW3jI1I7whwOzx07FZcGCc
eiGhRsaWSspRJtYCzBF4TOWJtW7BlZj/NI9oW8wpvnrfZ71pKLzDfu3kxIffJI5udHBqBBLUbhwT
FEDQBiCeiLvq7O8/eYdEqn4nGJmTewvQrRmlMPyqkfN3ijQ9DOxRIcTIYZiKI+G0h1gLNZdbbzPj
R/U9ZaYhxug8ffqPsOg8sw4vroM3NBms4VGY5PtwS1pftgAo19fyIajw01hF5SMpiD96RzUkpjEl
AQVcJl4bedK2+tiExrR6IKXG5p3RnygOoEoUP+4Wn18rSF0rgiOnHdlbBud0PRBmU2+tQI3p6FYs
1nrRwXbby7ecSZdv4kXCvnjP+M3J9cUJEfKj4LcJDjX5OuQX2Ptul1UDizdZI/XktydaO9Rsd48D
5zk/jDiMom+Oj/Bo9U0z/BJTrBBXExHk071UvEiODC7x/sh+GHsUSeX+A8JYPNDXQ/CZwrsycHzT
ndc30K77Do8a8AUYAcsfzmx9SgkDQFETsD9ZxufnPwz3Yu+AZZW3vldn7rRCCubroq0cm1XzYBs8
BBsTZrPBIND59/mX/+/QVSb8LpoHIL2wQNEvm9ym6S4wV12UxRJEpI+U/rzr2R0xJUXe+jbSeeU0
3qItrXpZR12NEz57bZVtBIch3u1PrT929MOeRMu5C5iOM4AgITU0luJilZFNpBNHvkGldhrzlIUS
0WSPNMCPaigolQPbs4tZQz1wInHyxjol0h4wPtg5TnUIuKRsfLaRmUyao/pipJ7VBxIfX52qwi+j
/mstKZXhJSzmbOieP62UB0Ho7HHQebHpQXTpdXzuZZO4Es0bqy1ZJK841/8rFpEj2Ae0LulzM9fP
TwY8p7e+/0WP3mRTgjCq3i4N92igFoQVqne5SYySYA3JopUYYg0Zg9FsllZ/Pt9e5Qtaz0VcoVL9
aae1Ihr54IJJMFFyZWe1i98/oqGtrOUsodTJ7yJQb2KRsxm+FJmQB06c55j2GeGqzoHUaXVm2RVz
QTsjcq6D+4IDeeEYmi3ytyr4Sdf+7jKE2xzAj99elK6o0JU9b4/g+CO+KiJDP7xD2od/VxChBPI3
qJ3TlLOSZLLpXfX1t5wpC8AYhAiRjeCS5ZkkYP1bM55WpHwWRFpLynrHtJrPTAYX5VqCKs2Un7/W
3DHcCDGSHIX+LAJVGweRbtEntbo7Id0zzeWc/xKIC/ha7mPR8vmSL966+uUVjLDTK3kAFDd4sN+e
b3XupJyQuzZy5yobojxHZlcvHI33RFUg/LmTtbxc+wpqA+gu71m14gPpRSpJHH49dh0msX0HIb7q
Cr8eZ96enz+dLdH/r/A4y3pyVmWkOjzEqnbTE78uKS8hQol3IbqBpwsPxKQfzBimNnEcXF0JIfWn
lBqnX48ZuVBfiUMgQzNjS2XRSaApjXlQVBduqucYrjUMnK8On6msGZgW2/mtXS4xCGYB/kjON0CM
XN83Z90pmIjWXXJyYIRYLczz3SZy2OgymeyVE4xE3M7RFZhfNdqj0OcgL/nQYmYC4ub5sWz3yBhn
fkAL6L/HOizAh7jiSW1xzTxv8JtwmWT4no8WyfRaxCeIXKpvm6N95g9Hr2HouAUGEEYwHlizSdnO
5FMmATtI7LzbJ6Kov7FVogmegoHim41OzGzqZjMPOT0VqPsnje/QYx75Nhl+h2M16fsnBobGIxo1
G+Mduoiwt2Popie8HyV4VDxNejYJSEikmKQCx8u+UIHD9u8Pjm97dWmCgs/PaAKLvUi4rLEVbCP7
665pC6wNdi7+Et411ZQoFpdDsrJKhOzIAxm8KVJngtGjesbYRvToUUj8bscjEad8PN9H3XCJvTI1
eapTb1wyWvk3j4gHwbm4tNwUXFvGxf2kqMqBtQ5SDgutzNysdi66eW9qGj0W9V9AXx1NQNI1bgxP
uVDP5XUlHRF8OE13yOV+976Np6Hpf+jAQnb6G7upjXQoWiT8wRtL3H2GqHodw/DOlQWTm2mCqOzg
21cCHxlBNSyiHDlLuEPmWsGLCya7TEpFZVo1s1uL13Yz42aANjrysfB633DN6d+J1zB+nWIh6nCb
FAf7J4sSmpUyfwf39qrS6sQ9rHpCz+T4vlGLFYBh4mZKaNCFuPQBD4NofpOCURtMTmBCACy9oZa1
JWS5ySf74eE7HUmbSm5iQKa2ROTAB4uR2DCQA1twtLlymSbmPyaVluYuB3zeTEET5UqTnk9VL0Nx
CP0dZZSN1EFamyHKs48QfxZlsRGs1CRRHMqozSqGnAkkGs5aAZtGCbUnJEjaJrN+x+DUerRV+tQl
RzwUTtbSJlk1h7SNw4hZgnMQMVG1rTJVjiTBnW/ocjtmEKWTHRzZALtrfCDQxu2jSZM9kewpMqKG
ZXwavzZMoW35nYG2to+3nyApcMR+NNN0acp7pSzSLO3LiWWTh20zNgHAZ3C3JrCTn1+if+1V4n8g
MD8UhHTwn2KqgJcuFCBEwrn8DP+iKmcnNn0FoKdgrr/sp6MUKb5AuLvtFGi3pkmLw5+rUk3vVA+2
UKffYUwGEm2b0JxXm86W7dYbpiRgK2lWzX7A6M1Bm1vWmI7US6lnZbuSyRLa/AQppyi/0m1ARdl8
zD9XZQo0JWY8M3q+pojh3AP1r44HvthhaCk23ru1SCggwLc72pTf4Tagfp8I/ZYqLYzUvpeoVCQs
kqZbYK7X2h0y88AlL6WvjE3ZcsAnkdJ0rNLuBQH2r05+2FIm6PELld/4xYfImg2FINARucDpmQ3e
RGJpQXcT8oUGD+C9FaYLWZCGyT8rROCjIXMnEPmDbYo9js5V+tWqSDCmboOgiRAeYWcdcSwISJfA
0QZIehul3JDc8SWfNR9g339CJ1fQkiJmdp/3pbeVGmTF81WhNkwkzIH9OARQcSZVipmfuYILDXGp
zpMjTtnlsaVVqujNfudBFkLQWCSJodqgLNuYrvHaKIbPbV+T48Z2inhj84VY3SOjRL4N0IiYqWnf
6urkhq1cUNJQAXw6vZu4TUqav7aQO7bhDskAehpedPIh7AhvcjaP29x7FZFLgn7o9NHEF7yPA+sq
vlVyiKpiHGPWVBq12/GbbjrW+TamoTi/6wVE10yGugIk9qS3h0XrIlA72qtEwZHytR50TRGJ6Psj
l+d7XmBe/j4AjlT43GXuZaSlOtSqiM8bx918ZQpMocNvKn4/oPL9soskdZHOE32YkIHzvQ7om0P8
mRp1Uh31/bgkTIeuDUeRYA1/J1FujMgKWsGM8HfKIiWjLfn6gfjBv4GZ4sifItFe5y4DXiaS0afv
f6rpdT3TjMLsBCsMF/iR7NbXKhIg4YI5KZUiI7bYT8+pWISSJQJLqFNZJCe76izWXbbDpix0I7Y/
lqrT6kdCFpxykyl+SJ6buuqJ8WDWrbLGBa8CMTyLt/Sj3TjDga0n0X+8wVYBUl7ZDbZJE8BeS8q4
dm/6FlBUNwPW19u507Kk1g3Y5wazsxdKyEofRtE2jilupE+/25Ui35eaRV5R4n7pFHBABHqQgZ0H
Sq8sAks3fpyk1w8FG3okV2APXlg7O4OXMUnoZReUgh77KoW2bi3HUQ6XpmStiHAaAJBEUda9WXaX
GmHqktCy8kaTCOioW2ERNRXlf0Ol7HHYUU6pIDBQ2gySMEv0CzEBjMx0vgcQuF/Qhzmy/jdwqeVR
1LCN5wVYX84Qta6deaDtuTDBsUU1S/G2lwg4nXGKNGbWPskO02b7u2uAXfFJddx87qVflxq/FcFa
24GsvzgzshCRPrAB5Uo3jSDCH8C57uU+H8/3Fvi4zqYcyJNPYbtH2e62GxirVnZDk5D/hcTj3jGa
FDCQRbXB9hKSojsPMM5Uw8gd4x76O8hV05rK9rKTnxHxkJmdJJvPL5Q1tBSrZiOTzYziL2v5EQky
PEgmtOMTRgWnYaVBRZXjv9T2VuGnmLuzVA5pv7ZrikzWjJkXbXc+vIyjJWhIJWB1ECdCC1wKGMRv
AyfO/16Kdb39ti6yg0lNt96Rk2QnWh/y2a6B2t+nsmalJ09kVZ2fvcWomi5PxBfFOoEVgJ7Bj6oN
/jl87RVtNarBdtI6Efr5mskpqjUF22SJ5FuLuZfMD79bL5QW7K6rJzMK9TSU9ZwFraVGdHKTM9Lh
mCHWQtdoPHeZL40DJZHOgb7jqWYIdsp0C3JPvmeyPov6Q+zZm7HRbs63oHkHxknAMe0/wZ60+3Ks
yJpRW3D9wl2dTe2VVYABPIuAjX3fENPeGjqN6pO6caBoPfGwIYHdhJJxCrf42+IwymFyhx47/KNP
QxwMcqQ2pFvXDs3Bi0Inq8nJxh5rKjQw6GxkzYjx7U+64jAzrJ00ZyhvXCCgECwChFGbe75L6F8G
2x3I4dYUWIlb00tHnl4tP5Hay8e3y7UjBT8bn3yKDIwNhg/PCU9vvyGWeLcYvhiKG1RWXcBmlJd6
5VFWD1vYEgL2ElWFb2M4zhzx+1Tez3Hd6M+bbcWQsEbROo1fw6dzZvuTK/KNyDVueV22RKZ6HCNg
KP6HFjGd/k9K/4p7WzRPBgCIDHydM8hLWwbi6Zr52B3hILxgPVzNyV2TU5+80moxzNQrOa+A87lO
MhdWxBpkgu04Rl5rAqaRQoKUdYVTOg8Ck5PWr6mF70Xt97uskW9dXABgYv+D9tHsd3cXNAORGo3J
i2OaHq8PDo1MlbHNuA+cx6aOL+y+ws2GDWcx08e7sQ1N0EZsf0qF1DiZN55rZhl/B8SmrPHHYLXg
nJdChYD8QBZccxY4ct4hGRGtk0wCULFJ81lHltX2ZDB+gJkss1OtBDfxYakFN5Haam61KJOK1FNB
+coWjawtLUz4EOEBeeVlRwwEiPQXbWlue2nCMAaGKUYSlqpGTd/Z/FkAUl+f+SyiUZ04REuu7zms
I7rj0Varp0thneMuDuhpo8hwQ4VZjfdwTz4SkhltMpXYw8g+i8KIMkF5UHKwHMwfFXii223fO0U6
RPsPN2rSg8tJTQxtAswPwpzVpRfSfKfo0ZqqKi6IqDk7PnDipC8RCvOG9TI/tfui1rkF8mCfJJoY
BLvoMNvKmBoiuFVwv10ODQpy/Er9vSY0Mjgd+rwO9/418UDUfZpp+OVYnI1it9YQ/rxRcGfC08zs
E6+xcpGnRCzjglwuhmc1vK77QIeKUM1spHJ9XwWDG7ODogu9wIIBmlDKY1jXhuxZLe4YJ6ToM44D
X+XnjpHDdU1wfqV9ywgZlPxCI4E9TFkm/5zNUnr346xpwdEx9t/iKFR7TCSd9uIqY46sDl5fYOXP
7JnLtMA+uiB+03xTGzrGycCqaQ/pS2m0Xa/5FLAucVTTMBh7z/ioVyK5tprKOlhqfMp4FM9Y10Te
nlhQNMBuj9dajLpp1t+gh5XqCFSX0xT3PBYrtZ1gMygsjMSOfU4TAB8mhorctlceD1dR7SRJov1W
E0gkRroF07ldS7dbq1DUNnp8hKI7aAKNqJYvxW5TXNNMtW/fdzST9afOJaenGByENazUWUKwzNwE
gsODYyjsCDi9MKFsGFOO0i7bnGxSr96eWIZh7IzWcL+OIuj70Cc+g4scOYIL+v+y8f5WLeYU+JQp
Q2sSPV1YBAq3WObuI9ZdVUO+ZMLsysNYg20g/P4DAGKD1jLHJ5JYx2Wnp8vfJO3b82PrEZJd/9jD
/AVZvmbno3kZX+vRqJNqlF2dOuUaSqr1xmu/9YksaDQ1+H1W21KDQ4QKzv1IrfDO+/GT/oGZKqT0
Bl7z+ya00pk80UYP3iLqZpVScL2IR2Jqlp2nPd1BNzP07J8zOBDMA7tv4CnFsDryiCwF0KJAxdI9
AZnW3/tEY6eGxxdfGhgxnt7AZWoS3B0d/qkrrqgd4J8ITdtjqYdz01MfoQggttec15bL412HMDIX
kCxOj7XncJq6nAS+kMCD6/6ALywQcXq/9hCCFn4pGQKyxSgI7eRNsLZ2kiiwbf33K4xBngUY5qlB
3UfblAxSkne7KJqArajwRX6QI5uuPL2rkxpPhxPeZXw1X3vtuiql4UhtHX93Y6jUgov5porYoHoW
whwSfgzfxNPO4LQD1ytGPNHT8ewelHIyNAQMBkWGQ1SN2ZlloXWTJN0X8llAzzCkTc+gjU8AWH91
Q/YV/0ZXnn5ln3TeNtAfn7xTu1kKOg9YqcUBVFZ/A53kgQEK/WG+QQH+jma9SgYcLlKAmC9uaExu
wLP35IJRkNp3vKJOY3gG378IfjGooxj0BpA+virZFVVuiUa2RWP+sITu7+exWjAEfx9vvJjspWbC
KqXYyO1pyuELYwkhokPQdYDzoNGsRastPzL1bqwJMBLOqbLsDKwJB4eQ2mMMVQl7LgfuLOaodrOQ
IAiUz6S2ZwD+SSF3ThiyTVjxBPKowBQlpngwKbhZkMjhYkNSbiM4v0QA9ZQwaC1DUXzgHQs248B/
dzeW7T2TtMmTRiramWWz4o2dhH9EDpRZZEY/WUqxeEF8JSz06YSiyq5P+deGLHq+1cf8/pGt/B3n
GZzqZvqVe5Ao8F5WFWN8q1ll+JRglTUvrvQYs4QUwqbZMexUdFRqYATg1QCZPxGkzFGwB8kP+KBb
ietFtaBhoOZDKvtg/6Wy4ZWrhy8CnvkHnd36+bTFCoTJSuA2kEyuswjnkuX896nZ0npgqinv+jBC
v9SPY4iB8bwBBWq8XavNZQgRJw2mkuRlNlRoloGpD9FqBOK2RotHm2dFUwmFclG1Rdkp66JwhbDp
7tkx1nYwwGChBtBVUjGWX0ekMnk4vrWHHJCyTfmq1O8LR+g3hMB/sEvBcCLSyGgYRo3sbnP4tcXz
QXKT84feUj+RHs2/wQu2Ky0/a+FlOOLhNVYhJvsw7To7/xu/vYxUMupy3TwqwmaMbWzPIh+smoX9
oLAEBmqq/7aEr8JY32gOETd3ZsSpFdodMgWQRbi5UOkrjHumDwQA0Q19jEO1kSBO046OZFnoVuee
G+HL1ihDzho4NDbr3r/fmnMJWijO2mLEifm/VEYjOFOQCpo7EGevRZs/4KX1C+L0CiV2x0ps5dSd
CZ/1S4yV/Hi1AGlhOU5A1g+Qyl7j4+DQf9aOrR/NI4qKIiTWNdplo+T5vm3k694kdkPBC+21nNkU
YQpOWdYT+r9FmLTYpkTMm3ldKEGfMi4UJn9Kt2vA/NEm6H59xBnJD284StEbMaSFRWF5X0V0hgtA
vyrX8XG0/3N1SozBHpGwCn7Pg0ool8iCY4yWTdi5wJUqQdqR2fQx2WPVl4IREgxCKIkL/DFDldWT
DW01HPiy9+/fjDeSHJQvcSxUc8LDlybUaRgsab3/JU/nfEHaD0qX62o4ICMftJ+s25no/YeCz5V+
6j5jiZ845fnwyEhyrdPrqq7WuV4v60ZgYdVMUANTAVThZ2lKbH8V2fU6rmgQZUmg9iaJzmSuVRGL
i9DIWB1y6SVkSsdSGgu8NgkRxHbOWzlXmyTu9CQg+ohP/2P/niSzXKHDpLeQMlQcpP8weVCqooYJ
7renX5300au5hA4/VLttkRkkQGYKt2/luoXfP1yRM3cPsOaGFvanu236ty7Mce+mFBZDDsFrKE8C
OdToSIJmymj1/dPTlE0aEHDRBYbRF8Zk+MiUt4Y+gObS04Vnj484aWpZ0yTZomDifYLb/hqoRP/a
48ox1YCAWlLvsWa2CMMdAhSONoBl1VvHyUqyO6puw+z19CDLSKYX9mMtJ8i2yu9bBiyOBGz91CDJ
1oVHNICyLrRpcH5IQh6yXg9R4W/qkThP4pBj/CWmZFaKQjWg/F7vjuygi1xbRVex+S7tSqX5kwVd
MdE3Z6mRPsVmUOJ0UZrwk5j3+B9iWuvOW5JKYmFf1Il6AxGSSJO5Vu/vB7ZzV2gd4Nw5H+/VHDef
fMKzNlXN82YgCMieUhNvm2oTqHgs/34bkpfS9LgfYrPRg+6gyeRYmEXpX3xkls9WuYXYSishX+1j
OG/6Ukvyy1pGKBGnzIj3UA67Jh1vvVy1RwA0CXrRLAoDcdjASHs4jP3yeEG29u01Ms1ucROPYh9F
9rZVAAez4Z0CKO6rNeO5Zz8tF1k/kGgeXIOB3wLTf+8ZNTc2JxiAdMuiINxJ159en3kQZX2b2Tt6
MtNpTndQ0gkpSFvYAUjCDrS75UaNcXPNd2NfGEw5DwnSLqamdvuRwWGCMsFemj5MMggvdeiGZEBZ
UpLpwII9DTnw4RgW6y0Wu36sgr8B7+1VG7BkF9qROLTjBGtKQtaYUycBq6pVkJDupmWCZu2rQl/U
xHmXkMq9BIUOoDFERusuDLxJ4rJSM4S8al6w6F9oGTMy8bzGuQ1pf0Gzxs1x7kkbGIuri7Nt2siA
GrI4BqTvcBGxZsbGLEPxFKuPBnSto2FIrEKX8XzInUVCJES6cJ/ixtklHy2wOdh36h3gmxa+noWK
SpHBy0JMPd6lgw5qybwKw8IbDQdZD5DRAdF1mlsFyPQFBLgt6udkzffiJq1zxaw1CO+1cEk7k6PK
sC9RprZjq1+QA58vr4jLcioF6L4swWAXzlQYX4L9eeM8KtoF2X39oxM7bNlpMCBqCp/oFKrt7QfM
jZ9zcC+U1FDr+6ZKgb5G7xxWTx8VW0BzAQvZgiMKnRz37Gfg2hamopYLlfoOlQBrpDDvRhlQtZVM
sqr1Qt7/6ndBUyHYXw+Rnq6PAcPFQ5T66s2m48z1rfMicx8dpES4UscYn1FT7U6b4+lrhlMR+ge2
As/FeLgduTrNL+CGOPwUi3kQbSGIW/TmCJAGqwo7VhveLm0NeZ8GQNE4XLVDYupr9M0GZL35SYmV
IcxRoj0DSGAm2UGK6H0UmcEgbSKJ25aZsr36xf8XDnOPekgf/OeZO/7RWpUtpJf+m8aSDOYJuHWI
HTYrjgXgusrSaUDB8AZi7vAaFI2tzv+ufTSFwPDkaQrrLMXIoExfTo2D3th/RxOrsgkuxQ3hZvKx
aqKMlAjI6WzIPIXq0Asn7234FTTe16PyWjLQfQhnVNju80OfFIIqzGFBWdLjcYea25Nz1S/LELSj
W+tAnj3ort47zvn8atg6hWd5KUSvFLmgLL5GQhL+xKiVCQrj3NUFDRcvfqaO+Fr4ygBXGJzv88D3
VIjQiRgXR3c4Ze3mKWJZDKSdsFwvxoCXcDAaarU3sDi61DkYnXNQk6zbRHZMTHm9TXEMdpGpW0mH
wp+VpfMo0u9dJvn86HbaN3XQJhn7a+tX/tk2s0ZOO2hYd8A0rcIIjl55q8N8F1UNdnHDm9wmrrTb
a7XMDcr/TfjQ/zWCc9p1oRWqKLbencmGuwXgUJ5HsWkA1KvLNsCDdmkwjmXdUKvlw225dzOjLOun
lvMXHvwwN1TLKdyok4A9mP0X4Iv/Iw9fzoLa+N5zxqdekz+WsO6xFU8okgUvm1+9ORHnFgy7YKWd
/r2uIqTkYnbLKupTXfTUjsabzLM4I+FCAMF4Ok5k6TSJwDolPx3IV4LjsOYUI72GG3E4k76kYDBU
snCZJby55XX/DOwIvW5gLVBx6ljgLqg9kjZbJ9AsHm0Lnc5MmLb5Q+yix+WXnHY2VkHtUzbPQRyL
Zwc2SQ4rNJ9+PKvwQH53E8xKli6DQ19fPVlen8ALSdaIwzaYp5GWkD4B9w01XZe9Sp7tmPNcESF5
/+yzaGGyvEUnPX1NgvlUkGeyZTzmYaDrOci60sqGHGIYAiyU616QwrsfHwRkgJ5zCIKr6n2ulYnb
fBPTmmXPj9I4EHq9OYysGDMDnPV4k4jNV5XBgi9cFdJUWkXk7ADBnzjpyNohzFxzbFDnYXu5vq7Y
aF6DAkCChuN3QXX5/lFGdHEyuh9Y+2TQE5hzBAVhnKyg+BY0RcofGblLKY1v6XDSruBqS9ikmsyF
YnL9Xn79hTI0K+7HnjEVc++Fs7deY/TTnDA3op3bDSC3h+fWO857lGocVQ7V9vIvDKHejvhSr1Aa
zHZC552gwH2ED00/roqmExGA2scxWf8DxowAMd/vvnuoZxoRCViL5ODVwZ0m1RjoBDRvZyQ/RmGn
b4ayT+vTiNkrft4zEvLdhwZX6PpuONTc/c5lqmuFcS2bOpEWV0WydNcsI5nHs0aweltT3DeNgJ8m
WzFJNajPh6+Ib7hqIKWzancvvF5fNoKEZfkQb9el8tjFcCYAjRz9vwXl90tCKi3wbArJv7AIfD6A
KdSAiGFaFXonoqeBmpIJuTDKKM0EaLhcjN0pk0Fwkzn4TrDynNUfKuI3NiUN33ApkIzOAmQB8AB2
8Za3IkDXFGAyq6K6qqqPSuD7nCcNEv2kwgYRyY7mZmvtpV/J1X5Z6541M9E0p6IQzgDLNtA4NabX
sBXl9kR+zood0P0s3A6nTRbSWU8rzxQDz2PpF2imuzmU1UurfIa2VPrYdu/KE190moa+uoOqhoMR
rzZvR3b7eLean5F9G4DeZmjsyfIuQxJyLXAq6J4LbiUxll2B3E8qDzjH9CtJgz+leUuOvfKdd4Gy
M+ApKZDSrOMXxPvpiqgJptv1cSaASpyH6zT2XJY+1paFflBgbI0VC2nmum3u/sAM90CksEzU4Z5L
qnOuMaJe816miRrPNdqGtDnw7u3GGScQyvucldF1WpyXWiWepvl2i8QILoe2nXMYfvNpJ5TvAkRx
FPOYC3TwB+MgFLmAJH13Uuhu82s4Xk9p/r8Py8ek9KQDE1ldyfjBGDaLrVlbaY8nYp2A6zNbbJ2l
lFg6AZTw4MgdOwY/5OGTyBSGUtANacSAw/6EH/e1LCx0mQE3FgM5wnTutFIgAzZXyeqDiczxLlET
DscaPDFXcqF0Y96WTz55mxbAGzVarT0a9yeKJxpxLWope3q3X6Ss1YdbQgOGvuN18wJmAcw6VOpS
6CVqOKrK+IlF3Fvy8jqcrXQyPk+aahzDtf3egiGV7RKjTsR2w/S3HGd0mGrmjqP3LD2C1LuPu07Q
RLlV+KHnltbP0PBTMT/pVm/ti7Gbm/WOntq1ZvN0TCdSk4att3A2IMB1LPQVZIA7+ojCBavYyw/T
FJUbgBNRogCuFk/AbfWX2zjsdjMFiiKV44qRCJj4b7hiLf5W9fAGpFTC5TXo8bV3o+riibVh7fCR
pgUyTWkIaxv6HZLQfz90czZIpOJxlOKtelG1e9y9/SAk/EWaT/p5klOaw/y4uu+ft7wrDlv4bOr9
6Ukk33H3lR3weBsxxvDrMFPWaR+VObPmbKq1Yc2qSNgIKZ0l9IO8TwmmTIu0+8v78IIk5tymfhch
VCWI+SVkQFHPQ2eodL23uRHrJgt9EJBDx0Trj7+0k1Y9pzxoYXMCoZC83wKyrJD+3LuOncv+2D+U
QluOlsqNl2pyJ9+x03JLirH7xqonfppERmgRefV7APZx3buj5cyJ5k1ERAufGIS/6GLtyv2fue2J
uPOsINOAKl3uwp/D13GgS0lMnSiSLoSxqTbM8UH+uDAS3TCID143/JfQkOPDwGZolo8P2mjBuZoG
5oypw8CKHuiUBCPaktZIUHm0oQVybn6Xho3uLbt801v/ZqeOLqQkvf0yFJQpSkwmxa5QbWb40Qgr
GGt1Qv3UkxJxENjLlV8VMY4M9w2tfepsiPhP2fcuExvH3AthnxdXEwg2upm7QotLrKLd/4O3ClT6
t0DtlM3iHjCwHzTbJxOk6oX3fEIxwvAuBPu0h1SoOoU5Pm1xT9AWQwJu2vzCy9VGtQS7814IiNp1
24HRmCfhoJ2XCYvaana+FK5j+OZKfYWC4V/Gh6UJq3/OraT7kybZvCWvcduodKMQRD2UjHbU4dHQ
C6YTBBanSdaVy/GstjPOr1rVOLhz+QgTqqo5faR6hhu5H+NUXV1psaYPkJfb7sLVxdzE//PYVGhy
famCBn0TQMzAMnWC5xIjP1WN96UcCn6JCRohVO6jzTs483kkuZCSTfZAAqQIyfi47CMIsqc7d/wJ
ygaJpI2z0SRiVp9McEd2Lamapg45QM5qRWhDShtBNPcLpnY9kqFffrq/MxSpBt7Dt2B7u1ZHaeap
p/BLtZvkhGf//uioPeIdTd2wuCAYqlS6U2CYgYMDajLzYcdZQ0HtGYcox8yMi8inyrZidN4kWvmN
o4Jdg3SNFwREKltDXH6MuKkqZmJOMpwbe+29Rw++fG44grG9X8S6+zm6AiTUXXomWaqGkBMa6vNG
ev05CE6JlgWHa0XxR6EpkZpf6+cBXjJZqncFeYAjuKzykjo149ws0JnW87mLQxcwpe+Rr31Ub4IK
3dDGSg0EA7/Kmh/tlqnzMBGADu1ztIDCWSdF3y/l0RFwYSMk0xl0Og1GbI2hy/hJY7pafcnAv9qd
gxOijRvHENa77UpobnQ7oNNADjDUhBS6fxchn58V45sR6XVYQaljegWevGgWn8EW6aUmqAPEH81n
9inw/Ch5uz7nvrr6yh+Vbm9IlF/XqlhWJiMNM+3z4F0KWtIpT2X5nXcBxCOyM+iwqoQ9B5cPZzIf
Q7OVM4LIh7SCjWjmpZvSY3bQ5WImH6dYZ9fUciJjQ0bxLoP5XLRCH38ceROR+FHq8U+sy0xSH8Yf
VCtnxQinYanYFKPK00ePlTrUMO00jmbGwTPESmTjCdrT0Huo4EghT7un4Q3xcOqhBbPDnqj6ygQP
2sbyKjHv8NjQ+IdP8kfinXqj7YkGgYYI2eXjJSY2k0Dst7JFM7pBuiKCLuip5eYwiSu0pLHn7k/q
7pHCmbKUnTIe7vnPh/16Zgn7W4uGcPI61+P45ffb2ZobhSM8cyELDt/QUj/B+x9bIZI8QLu0hZn9
S0pEPlQYAd06TRDJzGs6HUOT+69JhcoEkosxnTj8JDx8qyH6wggKZ7oYhZTaU9v7xEQ2mPBlGps6
KG3y96Vrl+FatcG3DoA0Ma2np0jES/Y9MBqcnLXo6vJ24Z+XYaXbgZMMP7d/XTUm4Bpuqzq9HFhU
YHpa/zlrhZCG+G+Bew/lDxxv4sTrtFQ1p/RRSjtV0qlfGPhIA71VHVboA1aaMzf6+lvwjLrf2KFA
Fm0m6MtJevwDTcv7hE7pyC5ulhSnGPBiSHiu9iekgUVN0KwgFNdoYj3PGgMduNCVu13ulvXBAjtp
SpndpJiG8yDfpjrmnRp2aKkZKdQElYMmHnPqUqmYfhyrekveWykB1rs676CzrHGd4liU8j9VeJ0s
J08gk5vdIfywFDTyZ7cLWPPgwTnT2iKA0zqRTxxiBpIGBnwDJsHnwIz/8M7iohEZw6TAQ5nokYLQ
8VysNJevkUQwPfhJrBZs6UzSoNg3csxGjnpnGwtq+FVuvRAex8opCLfJCvIDbPerB0qHNtTXyWqV
VpmzSHxuVx06p+ZrrQW/rVgRLQajmh037AsXC4OrEEY8S9b+/ZWenvnAtxYPvoq/SrAivtFdUaBQ
rlHASpZooBra3eJuOxDNtv8/gFFKzV7OqATxp30UJKFvz9nORIP7Pl1wCZxcJs2v4vxAP9WH5+bP
S21WONjUvcP0iaCJmdVYPHa3fA6H18PWdrjyoLSyCjLs/SxQH5PTuxZ7nS5ZjoTBwenc9ux39Rjy
RaeTIp8IL0AX/MH5IUTtvkinqg+vcj3KCAon8fccED8vEk01OyUMNGsGoRLgb2oIuqpl4C2wbbfZ
msYsj3yhpf+gHPA4e4OMNDxD4XnOBKmw5BPefZGNjVbcOUNsOS+1y69i5L1g23C3+n0rNHYhRObi
09RxvwYWkbukmgr3lisWW8ykGAM5QkPvAV4XRXEVJ+NHKdGlJ0nxgOcetWgwn89ZS3+siPxRETRB
D1ZXYuvJATiucR5sNf0zpnEoLCSqGy+HOCZCZ2FzazX7gtL0od0c2QTrmIM0mjr391VEozRaOxYP
Z6vyuJbkBniadoFiE/qpMbVLwVCfhUmHKJx14ZUz4raGHYF/URU9XVW7rSrRdtqlt/8R5zHdf4et
0gSXXIHeQlnLrbZtUeRnOxN211XgvI4AscK6coceE/mkFiYTk5UNujnxOOA8QQvFFhIAmQ2rB/f1
vFmQZG/9RpJH9E4+lLC1nsgsQdYBubmfTFsNiFOnNnD0Pb6Auc+n62xUVSOvjcT6NOIj2w/k8dee
UMheTDFrQ1rOSPrd8MYQR9eQWJ1EOjs90u3GUX3lUUIRuoKV/zWx+eDCrOH05ni7G94Oqb9RGRHE
L6PsM1/qYQBd9649mwMx44aTHQPWVSrdaTMy4d8iQ5b83uBgRao7w1iitXZcjQweBtOCp2kk6sND
b2Uwe9Z5gC/cyv8ybbx4dJI6C448f771M8T9KCuxBG4ZGZYFz7ltKlCQTwkM1Mn4B+BsqKWl7NAX
iHUOZ0u9V+eCRM3E8a4Vm/HZCN+gq19iOyRjBN878ZCwQNvcOB+mm8Edaw6KkqHJfHmGtSdP09Gn
SIKsfPXoou0grnjuwO5O2P5j6O1m/tHOJytzz9J5me5Ji3asdcCndB90TsVkXTh1znZqaNQ3fC5M
QRZmCmQ3Tqr9UaEdT62KVOjj8eA/GwfwG3XeaIzdrS3w9ZBhDHyIcPwhW0vZzNjH5efO/Tau3WnQ
yfAjk9IfXK4hb0LnRre511whyHTEJHVSdTn0V3vMpqxlVIjbWEheK3O3Fb0893VtBPFxHO8oJosz
+txRmLcGT/MocKolZlmBcjut/WMzM5KEnxX6nP8y0KO1jkKUfPYCRVKugmy899mWC2jq9SUz9192
GflIcMM2jYXnEaOY4inUWTZVI6gX51DFTIyR2JEzm8qFcI2pTWKftSVRqix5vCdSruXglub9vLfc
F8qW5lz5lBXVxp+/dq5fdF6eM9KYTaezwZX7l2y8ysj2hZv3KtDcT1EISR/9sXcxfZD9LSPLUcsk
9hUznv5OU+TFGG2Ys7CC0BKdbD+c6qPajtBImvb2DhVMK5BmRvMOSI8S84oWkZ+n03iZPfqSZX6u
ud8+Lgep2VA6Icx4Su2ORD5HZGkRcboQ7TCIE9CCVPrM0+m9BZEtMcP0yyz5XyvsPmjDBJnrsm+e
h2Uf3lh2tAGlV+pvwKUw/J4aOw3qv3xTJJQGqWekL37Z7UE/3lxv8oHzmwUQV/UObd7eaq3k/Xtj
ZmUV7Wok5sAsGZz2Yfm/fioPF69mBcaEBIbPxdw9ObYPBQw+IKmO20t2a17lqfCqG2gGHtmf+nxk
iphJ7xtowffWCyOgdPxcT81MmxcdpqhRoOqV4uu8eoDGjpNEgB0GtlJBgNxoVET55gpQ3+1U9bBn
Z+8dqpKpKCFbqNQdwjvVwTHsUUTNIMVUwXJHCKYCwsr2tfTnLPEA7g+0bZ6CGJvcToFUU+qaB7Uo
GtS6bJn5BUrc0YJUxWOEpjxHr+nQ1pBItoom7NrVRK4DXSViTxFoA3ADD4JAcBkdEMpI7J7tHNlN
rltJrbE1XjbyU1WD+jZ7qRqSOEusRsQCPaI1gYGnm+UqAU+rR2PEciV9+gSsF2Mc7/ZsteDyAhS1
o2vOp0T+4pPEuYKgr2de2V87sTSKs9NLFiX332WG8JSSYOELkbpGsQnRvvzYvsUxW2SrM54uDNV0
dcmfPD6y23oagmh5qolnnLMLflnFl/v3WSMUNDkPJ/utbnbqBsXZuO4GcHXOXR7nXXcfejqAJqU9
AvhjD5yAHx4kVFZoORJKogxyGgZZrZE9iu92yn+3z3PjK/vhlstOO8r+CwGlyt8IlR1K0rGfXt0a
gGbFHNNfqS2DVROjZm8AoALZzuUC26F8ptGGEVE4flw5JozCP40lpdH7I06DStiGKDvrVmuoQfP4
gRB2QYCudRupLytmw0bLwxa5SdOR93sLe7B4o0JhXl1Kkq+OjmxuGeqyEpq7uCjRndMD9FdCuAKX
IKD3IvehfOgomUbax2wRQ2mKNIKu841RpZqEc0d8BsCakUcLJlA6ITKZhtgj6Zi45qfKS+OllgQP
Y9DckT6UhLHKYyRGL5VRWm0d0/HsJRk4n8/VAhAouFWNgdsPSk76i7yuJvSel5hqLwrxelTHb0xU
yh9mnMGOY+LY9m9M4XoCHs5mzkn0DRJo3POWSeSbwqvLCKSY4a6ePdy+t9150SbQS20Jrd1uFYFY
hi9Ky264GxwhtZKNSNnfP6TXJlhxYDCH8e4Vrh0TZQUrX/H0rf4Gp+Z/NrM5x0cBU4cynpSdV2z2
3CwDoPM5zcKMYhFCzB+eXUuxtaHUL6OoESfOUEBGUtnJvV8USV+7qeffjq6gC8DeY1M3oVLy4gOP
aMIAI15CwIGSwCron05oARZABRiRMJWtNeXsVXDKymRKfCeM6254TwqC6ow0zSdBbLrHM2aF8ZfD
OG9tgn+Vnr9CCbN1uf2UQ6QZ9C2fPKhhJVzVAI7ajRG6GOSAw783qFlAMISLAno620bPmup1iwqr
+RHT1S6lznTmpSbGl/a2/QoHZXQ7/TzJNSm2/12Pm4pM3RrRuf3aN5ZbyZh/gYJ11vy70COm2AJq
AkfHrsHMsMZQaATJV+YyeMQckb41QGFHgsZAfg0keTdm85zriIM+Z0/XUu9RvrnOc0P7HOupWW/0
KqxHdcHRaWg0qTewgoWYkdrgIzcxil641aiDERIa6b9oHrwR9DyT54W3VZHhNqtVcBYr78S9nvwv
ISoCVHDmo5C+sRvcm4ikf48kPVlXH+0CGz2TuSow9RA5X3TfiaLlLGwelL0jz5k7y3IkgKoHDVGJ
rltOdOIAyomS0SVTmS5Tf/ipf03uEURf5DcvmXPJMh9IkCkOs2j6Ckd8oqXQFn3Fe0zhd5DPBHPy
ZTxg9dGzzPgRGJ7EB9JbSmKtq5OE9vlh+It/WyZA+6fo0wPavevYCUe1R0aeZMqPRL6cswG7de3o
boigwAHx87gLUgpWjrDuXb+BY5N4zjG8E9WHfFv4xiLjiJGsKCmAbZ7eLusv/t1mWwYxmQIrcg0F
qvDGlymqh0gJWnUcHJ076/EHHrYjQOc7/pp6K3MUBNWFt9M1YWPRf3W4FjfiCFSOfR0X3VkHk2ze
ylo/Axo4XRwIOANDbUcyUFOI3A0S4clCnsPpAZY+h0I1s2EXpNg+KnoeGBphwR7wsRWZCr2o0S7U
/Wju1wAHx4k+4wtLp76xUzSoMWWAQtMeSZ60zqdJkS3OAXIvAz7kU4C55tt26MR9q3buBh3suw6a
98PvN/gyeM9aNAPUtrT8qNn+MJD/Q4BF5w+pXEMxThCa554hdVqQ3zMgpO3KWvXTbryjDKIC/IQT
720VCQfOW8Sw15dFw67oTbU1Rmmhge5YUZVNB4nr8ol8/0rAsjebqwqhUaPa0HLoG3z4wuOZQK91
iWE0+BsDC0RAT6Oi1dRnD1ITF+DkBsyuLcUud+0I6LgHKDq86fsIKmCoGeigGB/J0gk6XbMkEfjY
/Ko1Nu5UiG43ibLsu3xAVl/3TM8o+uWcRYEOGNgGT5Wo4zNz+ARP5QYZMcRv2fQn+6dfSE6/oDWZ
u3QE5CuZmvJkGNhRrniTbcMUgwetPqSSXCKZ5HYKNdswvZlmlTuPpRxFKaa6lX9KvrtVwrtQV7Za
ILCAalmpLdb1ipLdcgGTLr92jkIMJbtFZFu9ogl1aUEwQCox68eHswPsxGabe/hjQaRjwT3OAEoM
5VYx+p0RzUAHMp5bnGlkHOroO2IfyfYbt60BdMVzjsrZPNW4wXV9A1Qi0UZksYdssG/opnT7GfUh
eBg6bYnpkixYjJ9U3kkoTnO3tGCPc5o30iExAUVQPKTuHjzHi62EKg19/c/rRwwFLLw/a0lgmE7i
1PknaezVg5g+Mw5+q/jg8McUE17T74Y4Rr1atF822xsDQ6bqbk58DaRpPGLkM4p/YgHLOswwJaT5
ZwhXn7OjvBPcMuM9y4RfSPRtwenyDh4cSNf9kX0oxwWatCzFjyPf2QFE17BWlQcmYKEFdr47J2IV
8fxKrkA1XnJOVE9hsqE+NmwRmhNa/EDu4AjNqEynVi5C+9vhINHnCfHiXGXZ319rox1fo0AsHkmi
jzWgivPRVVrh/oFRQN7E8lGLir+yy7+31LF5xuA9Elvzp6IHdiy4ebPrTQSJl2AfIksNaZ8QoSEc
Jt2MMr1x4wKPvFgEqjRrE/ySvGX43vvgcWdnb+9ftMeND6weDZjUCy1qQhPO6H3fVpPbrhrff582
j6O2FiAtsf3WuWmsAno+82iO05ncrGdNt5hmR71J7YSQLSsfFgC5yMj73DkOIklmhRRGu0m/MjUY
NzHjo8f/ZtySYqae0P+fpLld2y2/A2sJY3dBNQJe+e7TC6V3m6eqsBtB528jEXqQnl+ZyDU+KSob
DGfDt+2x754P3XFtkIpchuutSSC/zyhgagiBH13txSyLwognP0+IFkikSNEXB4HMgzZTeHAtbQjd
Ku4agvirhpMiRY2TnxWh5sz28PiJGsAiojAhtvvqC3fS9o7mEPO/pwnQDdcBBORnXVcpR+Jrge/Y
Qv+hNmWq+DaoFPJFrbkzKfVwHqWouauhkrmdq0tZv1o+/nXvQ6BSYQm5PPTKKkeYfHkulRZEY5ql
H7bHroIK9oENb+++7cbSxgaiaIChaBuqNl6GMum5NePYWiXTCx1R67wsAr+KMK5LiUumUjh+RHas
uV5MiOi8g1+fUwGjLA5D2YYUoUoWTsikyWx6Ld0nzUOJMB6DgzSQtcrtA2RoLwHd4whvuBnXTNYc
iQiVoLCnZvneknlDl5tF3gUjyQSlpragl2wWMiQ34ahToWLbaJcJAgrOEA/p65kCCXncqOM4ksUD
b5O/GTeQV1GqPun06R0xVytHlAxPEWBcHQA+b58X76H0MQACLHd787xT2+FFXLezztwhjukLrQM5
v+IEXKH1e7yKBtZkrlQMACw16s3Z23ZPV/B4+H8AC73UmL5QugkaoLozeWmZLNXfCodaQ1hKwMhD
NKwLHvBhAF7qXKlCctlPAlIm7Fm6J3GxFi2KjgJ8CpvFtqdjrdjCL6Dj5/Pq+KiE6P+O12MB19Om
x4tUfMBhUE7PJGYljQKfMXPtuvbYEwYCZS4s7DWBislSoHAyHsl5m4orWlKlB0uC9euELjt5mp7J
/kV1FwcgPOU3gW8USEtoIhSSv2s8y9Xf3UdZQ9oG7Jcc1MoV8yCecaDLrEdQXTZCv3k0YbIAyiBb
cEywnBxBseWJEQuwgdoDZbJGQuxkPkN9fwCx++PNiAFhk+g620s43VFzxPnhjzyrPAn1OpFv+2Y8
zRyrlf44b39fN77nwyj/5ONkyug+Bjin67BTOI+g1YUSBfKgnAoEasWIaj6k5ZVytXGg241Ph9/W
GIlmTT+GJEsXmNUM1pChFgEHgqVdCMU7qdenJEErYeTVS9BAXvgnZX7Hak/D3BvVRAPYWdyuDDda
BLcayHvv9sf/G7MIe/eQYoDAyXnWo0w+LrXEOJT1sNFW+NF0pcj0BqcHKdKUPHOmO7AucOF9jpb0
VL2s5M5MvVuDH1pBs9iedw8K6h85E+fktQxyitEzGaepjXW43EPJClXlbgJcnYLUCY/1wMmi7AcJ
pvPTpS+yDs7BHDpPMY02NjYDVyZRw+I1vHSDMFD1Kpzt5J6JUNKuwZf6VC8hbVV5yFQUJzDrjy39
gnfZ95MxL372I4IF5pSpt39dqKD/Pa+mHvpRiC8UJ/K/QS6ekDZJmxSFEkfk7VVs59OQe/Xo0Txa
XoRtC+12LlNqEx/Qku1zg24vj5k6d89nipPnqBFVpefF1qVt0LCqjMQ24cfQ8o0rjv1fQG97BQ4p
9y/ckg4Twyy17yrhXxQ2nA9LUrHWSHupZcrF4l9cPJLV7sKZ3OvNoPepk8Wp3smHYxXekTGOO+hb
WdceK5ADwvIW0EtvXSuCf+TB7IegSD9hrQwWtkfir3cEt7OLUIk3eV1m03sGHdXbtOZxcawiYV6x
2N1qyjpJO5JghZiRc745WXciexdkXj2li8irebwI93ad4UDcxf2VtxCwTcNiqPP9Nh+aE3JPYf/u
0uKVXWmdmB5B9MWM9p/4+XovbWkGabz2wsojaC4aM4AqKOLeHCnu2OKrCbaStzsvw74XB2rABBeD
LCSQ62v3zWNj9ci9HuIEpEKz8JkOpFBOtjh4CqWB0u8Ixo4CXwztxkkM4Gjx1ZIn/umJma9P8Gxm
knzMSOBvDu/9wKv6UmfRGmyAp3C+g3NiGWt20Ktb3kBuOco79CdOvp3roiwPGHg8UtF1NKPrjnam
xkQY3JCckL+qe+H3X+UgLdEHhzDJ/o0hJstKqjB+C0l36KFVkCQPOy3Fus/bcxovLD4ClfUZF1Fr
PUWheUvIlyd/9xS3Ad0II2kiu2q3mH0e9c+j4JmvewCrGtHIok0tZ4/umpCz+VYiMqN4EIgtfarQ
NIosdL0m4WAESn4xZM40RxUm+Gx4l8jHHbf4B1Od3jNJ8gkDiNOIZCx3WLFaOWNNe6PnAAKLV4ax
P2KsfP88dc81mj+Vy53YHyRPPUSyTsuGL0fmMeuY3GBQhsSe7Cor2/fe26Jm6AAv7uWk+B05kSIM
UV1grL0/c/ADMRyaKlHo0bugHhTTQl94cPAb7L+p0u31tli3e5WMS/7Ju/UA2ZJxqeH16aeGzID6
32jwvglzUOgPqhQFsPPNL/jnidYDrC8OAf1g4On5bk50jMPHIWxW2vyQjnkpVH6TI1Qo0dNAvaiW
K+6oqwJxRNepMu2ndoq+C0KIYk1fPY49rMIXURZ0kx388bSDc7uUtDgx4MLfytupKA6CR7x4rsTc
vYIQ0cNdZdKLPwvFsptyUwilWyG9sc2iHKshWwKYL0s+4SFfkdRYcgu2G2D4YtXDEJj2llJdnDR0
g70HWHuzbytJJhtae8T7ceNaCmTHEwUNeQTU1RO0XZEVhT/hvPsNzyqfwu1f41qst9pZuw7DkV0v
V52o4N15A4skoQyM5ZtSz7rgQLiMt1tYCr0Vge7qiRJolNUa37e1XgNguBT70DCAdgwsUVwwBX7u
3AFRBQZSSXgWXHx4rRmEYgIlzaT+S6KdpUyOoGMSTepJQbZiwz0xUT0DzODHS6XXs5HonZ5SY6Xu
7acmE9U/C82FiSGU98Q3xSjXgLFLMiSCrskoju5RKv6noH65waWuftUVglAPtOFJlIftNbYXN1bg
P77QVCowgJj8Lquz4qYhgHzf8C+EVjb1pHt8lDvSTLqJzXBirIJNbYPJ5FNgG8cM/Iqt9pBfhle8
CaOEXbGWuOSDTN5Y/fZ8r1jCQ5gFnehOm0DKMUf6ObOQC/xQBPjS1YGf2JbZVPRZn98gl7SL4vJs
WnPveAPJvAymWLR3AuzMYgogtJBRBa+Fs/Hcjgon0JJKblwOu/1loKnnQxNO+7/CrAkNsj3wM4GV
AYB+sMO6RufZn4t2WUooVrLI3faO4dmGWseuGQq9hg9qk4kLNrRaq30Nm5aShlBJGtNVTzyelOAf
wDeIJZCo9e++rNRi6bnJadZaRvfZMzcgi/tuc7I26UMufUKuJrpjY46klVFs3m4oZJ5641Z/NwSC
hv4Du6P6LKB566SYYMbe15dPlqs+4Z7dhL0ErBSjEfBVnEE320NeKdTKmsMdsX+Qg5x1vfNQhluB
NhLPtMAq0Edp5AbPgPH++HocqW9ITFwFvmaKY8no98DuLvE/CeGKthynaPEXZwV2lS0xCDYkMSDY
VHD5bN61uARr/2fu8AXRqfVjWGsNgRvTAzMf8QCTpYmV1oBqyfmpjTDGieSIX5xIel/YBrEwheXd
ppXEvVxqlCTNiSssVfDl9mQVQPsM0zlzhDGqg9zvGoC2Unm+GTxi1qIPGmp9145c7z3QuaPbpcoD
5n0THrNdhcbTRlriVQ/Kk7MQFQPK72pAIE0j8pxBzIcxaCcWeGaN71tFqmqkdrxWfc8j8eRxmw++
5AHVTRa7jO+Vdkzd2UDzZHtrVnOGsGfE7sUzRlCLBL/C4xRAWYkT91YdXPy5FdEoX7ZywGYs5/0a
Z+29aeR5DhjlvPkNJ6GLbVe4pcEIR73M38yGy9wKYwL2pVk+8obyqfTiDhHdS1AG2LmziN2O7lSV
8ks7AB15onuFnIfS4WwvNbbdDjuuLXTgZkqq0advCylDt9SbFQQptdV9c9/H5c5QyF5Xlyo7QkVC
4em3H8PIEkrF6x3r6WVTG/SdIE8ou+U6YT9/Z488Outg4RpCIOXoMutTH86CxFLytKRR/0asBmDK
C9Q4mwU7qMYBavX0Geykqc4NZqqEtIl7+7+3wUfr+Andv79JBLyG9qdLb/zQLO/aE3HhBMVQSNbe
sTrmJ3a0QOh6Lm95vAigTFCzraG2ymL66xGXoZKga8kCteXeHdwlqfFr2W97Yp1nm2lRXQ8h7l0U
G4olX5W907dbLh90GrVu7OGAFKXa/X/IvxHRooNuOjP8zjJT2yyfJF3lnKYxEHafqJAvY/lN/Tb0
kAkwtSwUGxiOFh3rEj1jWkhsPgM3I74YfM/Esw79pxHDEhnacwpatmbQ4mb7RbFuG0ACw6EMBaDq
XxdE+9S4L6C6wMUmqjkJbNk+Fq0u6O5lNawCPT9pZm/b7674B+105iDWHqIEZbbJJBQI5skiAWAa
5Cp3v39ATgm3EAZH7G8UoBHeJaAB+Soyc5LbjGeN70pjwaZn/z05DO2haD8cs5Y3nz2O/pV0n8dn
WRr5SAgxC+yTSoB73+8J/bQ7fvnmLqiCFbUNmBajRGHF0qyUI9SrO1Y+piz/IzdohZD2pgb0552I
kO0OVEbqWiPzagowDv1XfbdWsZ0m2VAd1GDTBqO9oifd2qsqgnP/esSetuEuCrMxp9PhxBn7wTwH
t0PxvB6q2fXzgJDyG7jrxf/ITRL3F8PnFqTG4Ly/YtR+DsY5//iIXLKE+Dj/iFVzzKlqC5uGbyA0
jwtXCq8toC/yewQOHAqhO/8gYb4wHNoM+rsi7IOVrrCtld+5M/990/a/E+Hc4FuZNM3DCsn+K5jw
AFqrEaYF1P8phc9S6V2oxqexCbVEkmyNfrXmEZecleolKFlQ5dKsBaqkwI9Fe+VfnLJ2cQY8/qRA
nB/l4Cp2nsfdjSpI3kh9pNU9vD7mriqWJTu8mk2ydkQ5VMmTlPBs9ar+Df+Vszq6cLTBE93TdPxT
WHpTh6/wzwi6jJbCA3+lhkOmaObATQGvxKAxY0fC/UBaKlYdTuUTfSePftEsAL1I6J1TqxXNdVpc
g4S0rWWa5raRlzIJ/2hsCQA0WsheCx3uXhc5tekTddkK5LSikdsfYphVtGpRy2FTPC/+5tawLgy7
C4DCSDXS8oJweo3wv+024Oae5YVQqxyM3a/OSXf6GGIpJ0np4kYhRkpwjUYUFXeH0Pi4P9I/fDU0
bQN4l6PF2mC+BHj4b2VxBEMyWfpQH0JdKN3iZsYzGiTaLG+/qKFcFOqrJtoNex5XX9fDZPQmS44L
rF2sOH8OTDE/Kl7vcYtllrI5KRuVhGPilZdsq/YqRLFwrnyTsATeQGgtnqYm4mT6hnyT/jXdfQoO
oMy1JAd5ZVCJEjrlgRk71DMgXdZZnTAs9o4Py2D5nDpLzUZsPQNL6ULdSToB31eCNrVFQ38Ta5Q/
xf466WUUltaWMLlFt/UntFM4M69JdUc30gPHtqg17koLYkUZzSu8n2VPV6hiCw+7zQ6o00jW/WTx
C82OaZKdvy/NIdyOsr6KGzvxC6by9VczjM+N777DjD5xSralEI8SHwe1tGTupMCl4YEUGwN94VPq
o0OPb01A/2eNalU+MWNqIzVGZXQ1aOLOYe2Pp3phGZiIzmT5x+ix8zWHsWh6jCOzg5kOgyI4zgw5
I5rOeSx1xymJTMfNABC60DfeSVWJua2HKIpc2vIwzhFhUslAFBzpD1oUeyfFCGQ0qYXQD5PXm0im
naHdaIf/+nQN4/DRp8VpHTvcRYNLbk9ZDNulSlhU6x8Q5U1XTG39drj/IeSRJECm/yeJpmAi0iKU
mf+jkSesM8GUDFGwt5o5dv3QwiCmk/iELlJrJu7tWT0mZGP0VSw55dW7i/zWxK7WtW1HTLbIf1bY
OWHmShzVIHvIlvnZ2+M6HmOZUoAZ+n2uvyxEJJCBUeqpTWJiE4TwjeYwQWcykdUzklaGUvyDOKr6
aAoepFjSeOm03s5b01YKhz9X+1PPU8LqYz47NjzJO221ZJ3z+U+QQ00bVFaFosJdaadVKUDM5klX
RB8wlvOyWT0hSNqZYsSJfvMYTAV1FqB8utOdFTY/XL7VkPtNxB9MULr2oP7QkfByk/zkrilDmpeU
8FMP4FfgTW0nK2RXmdPLTy77AlVUHcOmPIPwoo4KijJ0p/KHgKEcvBjZ0xJ6dOs6iNIS5I3KsxNL
U+quiHFJvoi9J9ZVEtv9vtZuhM0yqs27zx0FmSu4KKJS4mZUaQqVTJQFNbJQ/5R79FEIAzMYUw6Y
PsGzMcpJVctCtO8lsRC+kD6TrMuq4j1zhjxed9MWHbIYa3yzD3917qpP64WITUIoKgHpL2j2HUpa
hbt+GlVlutkKJgmSbLtGSlfKgmH5xLh9AkhGUomd4m0R+qlT/9gnVWXGE1MMtfvEK3pZAJHoClQH
Iz0v4Ypp3e/GK19aY2qlLSGLo/gzoOZTCU5hoYHLrdLMHklW/owM3XsVXPcxdzdaAmxelhXJHIgU
8clPjzjjCpMorIKEnFFbwJ3A3mMhygdVK7nDT7C7akPLQKheroA+4ImkXUHNu69IQ9sC87oJZfhv
k5ZMDOjKAiT/MfW69POWpeJS5ELKzCc/TzXtuzDMFZAcZdW+fFdh7+lJ3dG9DGTR1AimLFO+kr4E
zInPw8BVnd58+OUHbjWXR+q7zbd/Wt8CSVTKFku+wzmzi4TgMHCZFlViioV22EHY7p3qa9OCOdN/
EhM2tSV4Mm+KX6XcHyPg19YdkEub9ZYs1xFIX09G1C+f7DkH5wJLCoyVIXAs+NQ8TsgzH/ceAWjG
ze/XAyvowjcuyWKnRxC/tcREM0ygRCKeWXCLMT0LNQtGSM7koKyH8tmGC72J5Pwmn+Sj0+aMHCXY
tIXsDvOKz/Y1BgshrK8UVpOd8HN//c2Wv8EOM22dcD2dJfexhmxGGClDSF353bXQN/WIEYAmk04J
qeJkeJ2kIYyG+mjJOGe0IwbbI6I1+QglGH2GvgyXXw3MbeiUnKL1w1rEDxfBWqphCSaorCqhM7W3
Sp9eYQaGpfjkpRO3xcew/hf/tTUkCXEJ9Ui8S1fLa5TUQXWUBsLJFGwS0s+WqnuT5D3+UxWtOZgK
0+yt4EUj5dpT7We0gRo8ddF4WpZKyg4uSH42F3UvIjHShZUGlH/0ADYOw8YyAfF0aElccuKT9tPx
KJ6WznlzCbl/QA8L9Ec0W7OAEhGjk0J6CxKFdr+ofSmqTnj8PKjoArvzq8FLNJebhxIK6TZ/cYzW
fwz+Ucvp9sE+ORw840QQNth/6nGu03aexSKnHyEs081B6eXgiKWUj3MlRG8W7uaI52SnfVho27ss
qQLT9nX1jS5wxGyUSSewzQDdBNGvp7eeeeut/CMhLcIKYGu9VRVNL4oGRTR5Vu8G/E/gsLIQk8ES
ZNqZfd1F89boQD7oo8dy/At5hHgPH4WaAjMsUUMNOwxhx1RK9Z9JgnlLf/OHz1pFT2C1vuARI9mF
R4tZW+0Mv9UfSLCUkyJNbz1BqPhwm021ZM/hy6oirXsQLSWNcbQY1z7qe3UBvV1HD9rCLkKk61Fj
Wqa72ZXel0I8NoC81zR2+e8JZ3myDckTyy4sbs6/ycFaglDiBZ5L7WvgNhu6PpdBwvFyrei2q1Aq
5Z2c32JDiOE/L0teD0NFDdhHw3vQc9yly5+kNPuUegBExts7EsCqRgzID62gb/oJyF5jgS/XaAvh
q0ZbNr0AAyOiFsUNNUGZ9ef56LLIG/EaZKFACRCbMqLNvc6PDq70M+l6ZSIavwjv6DSAEDXOr54q
4q+bVNzgckOzXSgWR+aeGT63FWu/VVDFDHEKd08Yj+SQyYSJ8UyFntH0AAbUpiElULrSYADMMfSi
34ufRjnd7jxP/MwaKi1zcvPOh7t+a+WH586kqd45rjE4neK8B8lyk0Zsw+MxUTF3B3mW8eS7W9tW
0u+jV567SM/+JmYo5khwTwpsu0BezqRk73aRv+TJb6SkxWfEciMNH0eAM0ncp1bFUnD1UM/imgD4
itY/s+M4gbvmyGgQduzPFUuw35lIe8nCMidmrVbM9KInkX+cT4GgVg1+Gt+pNOkAtWNsSlSKTVuH
CSaC6gvps/iDjvdYsYnaA5JLC9oNk9WPCqK4OlCZX6sNBKABH8xQc0hnWJIblNaqTaqgZiZBomMs
f2wX8AuSRSw1ZAIqoyxXz1e+nEjNGE+N1qcFA2oV4+wj66AsTOyLn1gM9yMQHSql0QNwpdqpbrYk
49a/Ztcjc0Pym3fEd2qmiJAio6cdNJjS+RWgTpQZio4GC8QwfYOLuBFvyuOgFQMRvOvERgNp3jb7
SgUdhhhpmeU7AlTalJ+jkwXBB6r8bYGLBvdZwFPAGF2enVkMWRsadoRbFEJVWrXuKnSPgIrT26Wz
5zCCnE+2HwtBM6cAGo1zp2toex8WepIdpFjzla0fMCIGA+hLsUmq2ct7g3KR7YgEla1wwt51moMn
YYFQIoiHwLsCzDdCgNUl+0WowQE+ERDobA7QAeW4iP0w9DRnok/owkvrhNpSzoeiFuujnyBVchzX
PiK3huGlHbmXD5TnUW8FYrBDYbPS6z9HfxLLz/SoxjlNcEIIqTVS1kYaWDTJ5ZJEKNftOkQMzXBg
/LjkKtFQWFUOGAB8JdC337sOtx49WfUtg93OfCF1Nz5MQsydp/dcNrZOqpHTNslEpaxWGXgAhBoQ
BAas/C2k7G5iJzwRHWO6coWJHFnZ9u8/RvyiR9y7cAOMFxU83Qyjzd2Octui88DZvlXlJEmcHViK
oZWDrindBnpnqsjne+qMYfWnMVgdfHco2CqLr31Qb/yM7qeGDZ6EfSGXWh2xHpVT9fQnsru6Uv4c
FUUxLQYy4fgKnz5IdmI50nUDrN7v4l0BZ5+OUhdN8l0F5u/aGld7A7oVVq67sBoOBGFQlBQTTzgL
4aVW+KhN155ELA0NvwW2pQpsjhzXdrRCVGgAmGKTkbL9n/RTAmrmBmr24wZFf2W7h/GAkAlghVQp
f2apugtDNAzVljQzetF/Eqmx3iaJSpZNisPKveLf8LeWt6laO02qfaWcXGrdAKEB0wl9JbEgchw8
Ahn/75LOrLCUnZzwh5flN7RQ75W8kukN70DIFRwDtX9LvDODBhuOC5QVa3Tc/nKLfCuv2+7fjLhF
V4fSAoJ5yvByceherKVRYhOO+lchKpgmO/xU5SVyRffFwq/S2kki0aK6FhYz5qdyd7sO7GGHVDwO
ENp3t9BHIg06PV5W8ycWjYgVURlNWUBMjj23QIrMuJTyJCwXtAMnQCTDU7Uh75wZfQdvp5MaEGAS
XGvZCX5YQBsUB/DoEEkXIonmxuhOnRowh70p009MmF58xpUBDSjIRXIXqjkfGf5dIESlxyEoak7v
bcwUTFJUp/XMianttzEe8O6jFT2GPnMndWZlNU7OVlQ6GsfvcnfSNXrVyT9bo05ugAQvPJzbya06
p1k1aFpU8LIORX5oNeU1C8jHeegUlW5h1sAu+lcoX6aADmmYEykOU6V+2LCThILZNKPqoxyroM+g
zFGsEGiNtlfqK6866ekcutXR9eVNdLoR6oj3VxOLGFQgStleF3c42u+jP1zOXnOYzuS37SrAF8yc
ZvtgNXQKAFuiA5l69zsPS9u2gWWOCXSYOiIkZsKKoILLh9DDU0B2c3IJaN1/h/RqrdiCYuRm1kIW
1XaiEVHS46Z8VWtUPBxujEDPYgarixmr4z+4mjni0ZEvyGr7Q2JO+nZLNT+6Dc4ldEBuLGgIrnwW
G6lIG72pJJBw++c4y5zO41JRf2q6dWSQjkK+2kckf1iqqGI0gF7sc/q10G3Ubg39Mzf/CIuMwL2M
LK1Ke7NrMBPuAou9LiawUGFU4oyHHPILR//yeyiBRAs3f+zwUI+AUj9VWuk84oklMV7fJwxe6AdY
fHfTLUtArKqiqtaEuY9zM+u28Vr+Zu/g19ySD31tfMG5f37TXDsS2MLpTVx9B656OflzVJucNF04
K1Ae7GYNE3QSHG/FXuzdSz/znl+bcgE0vaHPKYxc/t0ysPT4yVn9MXlv+hLcJ3Ymt3IZ0exs5g6x
9xy3u9stc1d3sw5Jl4vHLXF0+Pg+kRCSKnoUUrwXIfng2btpi39GwFg7+eiwbweFClDEN+tDLexZ
VplwmuGaDLqc+XGWPx4Yn/8S3GsPIdhqEbaWbO+cTPhpqUZzatyFm0LyunCnhSptNeSDoZU1uhJ2
Wsbv6j2jDHvJxB9lMl4Er01YB3/1bRLzOYjSGJ43hbU7o58B9erHQPJzSqO27mgGiE+n6Xl4mIw4
KuZCuRmARnXjhC/Vn3pJVGaDIOo0p/fUFRkX9Udj73NxhEaz4XJVa3JVpyDnTECEVsqwl8vVB4yQ
zC6G89bLs1PaR/syz0ManLniiFJ0UDCNox33D5NoAw4VkXZnNdDac/Uw66Vz3tY4tA+lQnIM6eRh
PZ0SRsi7EGcQur4CpE2r2FFwK8AqEwFe6Un5cv581ozu+SY3HrrJsuTWFKh9yA7lBo+DAIPmrGxg
XFTklPG3lyUMDq9r3zi/Po+DmUTHlCXoaSWlSSTiDp84/opxkKOkHir5zQzTkRliQC5aRsJRWxSV
yZj6TOoXP43cqarNTDjfgZ5wlk8FagvXwotfGNcy1+ZBvZCKq+x7DDeTzqnQOecioTI/yiX3lY5l
fxpEwNdNFNR5f9k73lWpRQ==
`protect end_protected
