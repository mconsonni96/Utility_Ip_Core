`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
tzIDlW6WhZZ3OLQ4BkKDiK9Ilec8Y+QeJ6Oi7TXWQflF/xTt5QDsowifi3CXWqDfPCbLAZl22mUq
/DDrLioQ3o0ZP1aZnpo7Zr2RYLjf26K1hkgdBcxEseBlGE1oYQw9Mx9wHk4rYA8SfegYrApkB1Ev
9k+PPXMNjMW6wRxjGkVkyrHCF7+kjXGmj5lUegjN5rcvBgP4iOW0/TlXZZgMkxPxSuPzrfLRWXLE
Gr8Qlw/nBXHaumFoir3OKXqstEZ1ytx1a5HnzZjvrDKfUVkTC5Mv6vyDFDhzYuH6QvMpcE9dK3Td
pJzbdQWhT2NtDQ3hWHFQV4UeVNx6SyZ65jlGCQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="RL3Hpo8TRSJ5/YJWu+BfWkn6r0HjwK88PfP2RqS/Rt0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17168)
`protect data_block
8cwrOenX5zZ8hjOF0WZQSvL/FO3gIT9gyIQvZl0I6UnKB2R3FUnOIi4N50m7wnOHnRHfdhg8JuRR
RWFGogIE9BaTmQUdeK0Iaw696Vphit+fvVa/LqNbYEjUBsx1VEcyKsFaNmpPyh6grw6hatdLnUT0
mAYd8Y3uBQxUb7l9dMUzMr5SxAKs4MALNS0beAbf/RPl9czWIJEPD71eDm/KWULBAxxpvHuFpsiM
znvZPkNZAE/1fYxaU7nDkc1LQEI119rCWZBTB4+Uvq01tqp2gTvHPcs+S8N/EUm+qhlIAwx14+vD
4HufoRDpZCCTr2DVmOh9lmm7hV1FRFZB9NykLaFYahES+5358lZrC+rdlDN5f9IRHZ1sR0praE2y
ZNBhI8D9yV89N9aETFK/wZ27BET2inO18ceuL8a2Ddga1T3J3HfQbxH8i7euPgWAnF5eR8Jp/V9k
BWIt/XibpeAeGOvPt0zXgfn3TSGlB1UQp2AaCEnwxZXhKTZ4mDyn2m22H4dO5x76NRxwem0/JgM2
WwEzWoKVhglRhpR6kGE1qZOFsdbR2VtZB/NPDC986wRtCt6XZRDBraKlNElWKkYnh3F5Ibia+pYj
MZ/ZaUFz255G6gn+v3O3wVymLzp6L0Hbwm08HBMgY43IHLLU6Dl+LI9+MTYuhxAl2zMqWmOsamnJ
qu8XuaKlOB9CSYKUw46wDbx9U2QEen+JEPiYRrHDh0Qfwx7t66aItXyJZeraajGX8Ol24z1n8YNw
+td7c64RbdnOzFvHM5NJOdwQhJDorjyb5ycRxLIm9AQIn9odfvXpLkgXwTJZjgycW91w7FPSLrTp
cd3ef9FslZw3NB8l9imAjPE3xS1hqHImhJBgrUvsZv231s1m6PAOsadDZdJ+J1FKfNrvMWUHG7+a
lTsAqXyMQ0ZI+sK93ghmTzor0PBzCy/XWPrJtd3TlQqxblLjz7A91FsaD3U7Ai0HM4TilFyVh+Mn
E4nP7ZyGXf2rzXvPT868rVcHMaUEl4x0YLLwfzlpMuKhJEF1wUijHMNWa2REuMzSvtS+bE+OJleN
4Ga9v1RSFxD8mL4AQjCcNj06in75lhb93XAde4QE7YcrNFUBtqV1Sfy8Rskaj8eE2p7unz/oa/7N
VDwL13vTsGQnqZtahw50aJ4eAWLMiA0vQ5U9cIzzYphEUH9mevqAjVXTVFOuV+k0IeA3N3v1Wl6q
rwi2ffsi6fvP++8WwSUZPCmh1e66a19lCvhDzXABxfNwrm/5DDSBTLAK4tbxhZ8BliW+zXIyjW4K
5ap+C8JvCStWqHwgU1gzkXoAG0/QomjTllxIYbDBSsPcLI95XFfngEkrQijiY007ho3ZJmfKut4A
b1/AknPZ7ByOW9laxwDvfLSXXyAiiiq1SKynm9TPSRiEIJ28+hKmOvHSG/ZxuzlNstSpbJZs5v3r
fQQHLor3WRjE8jNCrNG7+wSmTx9VhGuxvrD5uPTEbNyPfcylJhvmt4cCoQor/tWRKw22N5nzLE5i
WZp1cr85CtDKSF5jVOCT6LVmqzG02cy9GNyIcG6ydbAGeYlKeZZJuaYnRNS8P6FUV5cJZETge2/Y
+pjRQEK8dYZHRLj+YWdKjJvKCd67UjZ9NQxYGnEP4Y5aFX/egGF7o96/jbw/AtIZ1zhOyT+F4jEU
S4w+Nvjb96H0VHHE8kseejAmZqGw4PM8qffgNoMoed8qm7t+0BKz2lbDPfajHjq5h2w6EVSnL+18
jQP3QwHGJMUG++EGAbSSFAnuvf6kxmr3SEckurlI8vsiq52Velv/yJ1AxNrLfKCuImTkMftUoWon
d7LNh6PfC0CpsBcAz1fVVnZNQHd+m0pJOqeHrK2Fs09Ceq/HyMNnm8Ygz1WT83njmLtLBuuzlFQB
4EGATp87wlT1kTNdMLsx+ama/uq/6BNO6UTLEiGLLVqcbSykfyvrFNno67CdBEYZTBpi9UP1NrC+
Icy3eyS653Sqz8cQuifbefqKwLZvrV3OZ0fcNnRNAPTsPW2/Sry3Dvq66bbM43fDsPzGo7T0FEjH
x9IkdYtV1Rw5JWn5RC/ju6nLKvKnw2zh548mmKrTNh8oZJ5IK1tNYjF9OsRQTITi1BLsQLXLLu0O
fKpsWRR+wpz+IZNhjpmCslNk/74RsKo9O6MTNdcE5ZhzOV+0SlwLZBPB/HF4LdYdWcdlDrN6lSUu
lJXK4WD8y3t0kiyOm953vKYHRDPkE/5zA2Nb58vlpP3ClJS24J3SPgm+7tQA0ecL6/Arjck1VzIo
Utr3PL7iW165ip8tO0ufOCaO3AlPF+ADFUIEkp+jiYd+1xFa89aQset4f206+pf+NIPlF/ORfndk
OTYYAxUv7OXsP5Kf4oZ6+0rPXHPtMbYh0DgiDR0ajYOfmv1qtASdwiR4IcvbGuR68j+tT1a6j41X
I+Vs64MbvyWEYMS8F4fsLBjgYz+Ewd6nWSpj7/jGZ54ivSs4EZSmnqg3ycj9nfKd2URBfCTlYjte
RSbvVJ4NmSl427/v2f0AFGdM9rYbhWCjkFIlWk2a4tXi9097kd0+q+M1cRzvlSAy1+f9rzUfF7sj
ViktH467Lo6fn5GrnrHplrmEJMdQ6RYxBhbl3s5BuTO0BcBQmIY0v5MZ1L4y746ars8DhDCiD1f3
08R+ApVoZLVGE54JU5bxOl38HNx29NsHiebqKcpzpajJj4OTzSWKrjHkQe8L6Hgd8OtyNhyymFKI
Kwti45dSbAwWADMr9cUIAXBSYwbcYZoavjcixZa3sOzI5bmnABjf5YzJgS0ke0psJVtqfqWTZwA1
HD9tjiIOIhmZ1uyvsnBKkCtm7+tpGRxG0LTEPic+AOZAkVR3/RRm2AM9+BmXTKLk9+jURgwK8R/W
VaPjxZHJDbN9LypKV9s8RbRhIx/vruUcJr2u+Pk4a40gVa3xEfvjizPsdiq1jkEPepEBjRQ+LjBD
8lHegFA9fuzy/vck9bkWDCRt84u7BWU1T9lL4VZfoUsQFr3qmBF3LsR/Q73D5OL0uWRV7Yr2AmSO
atGktqN7uKDNuAuOHdvmdln9O/C0J1rZ+ohjcJVOFqdDDcJ7FHkDXMf5NcvEUzlRAHIPe1DZLXFW
RB26ZkdfFWRAK9DLQFPOcDUP5tvTUZHrMtF1MH8v10dMZDRcK1jn6Gk+o6YPHteHYW7HNy/qKgr7
yr112KKQ8hmP1DNj1Ge/+we+aVxe0QvYCW3aZUsOcVyGb5TXZ7IOfaly/3hbcI0lln92p25hRHy1
l9wz2pHZVNh3fD3JogaUbB2ScKpjaZgLZzgnrYGsK4uslBVKHRb4UA1eyTnvykhycM7TQpGWL1OD
cIsN+sP01O+XRlzY2sQx+oL1ZiDhZ0rUsXUWlCbWOvpDQk6T8Bt5izvn6MJgYgFPL9y42ue6MgvX
q+TCZpknoZ+vTDxcBBJmrIat5qZluk8fpxFUbgkzKepjnvIKwaKNegIuksDIWSqTlmJaahHIQa/m
MR4ZFleKbnjFUv0kqVQVA2AGxvRd/I0gmzLwFALSxVepAgs6NaICoQlIBelCWCWwH9lXDi+pZNol
9lL4Co5JHASe5uVWVyfaYbDvknVQWPXvi2eLiqxaCvaX6BjvmvNQBA2BAgROm9K2Mj89NkVLXiuj
vqP94EUv+ahIm+gPBrodcaQlEtKw4AzA3179bYRxdchyzkVrDDm96xdGc9FJtiREzFX6Z2yQRei+
4E7WpzK+oWtY2hbwuZWQ51LCBr/DSjww8Xz90v5TijzaUz7c7fPBVpHrbpz5bHZUh9Py0eBLWqLr
tDrBZzGzPjB02fP3RxaKFUysf07col00Tx5f7jfUzXdnMgMjvmASgvmjr8JihjFclTImn0dzg0IO
5PUoQQH+4opK3PFKufPwV6P8vW76B/g7nJwv2xiU8H6gsonTztUrjZs12ij3S2tByE9jRQZK9RyS
5x2LqDb2KQdUVF2jkcQmpebvxWmUZO/7H1mPIOagvIed2qE5ZXdeC04RCVGvadOM/b5khbo/rY9P
FyxRJUUknMsvh4SWri0oQz7JQAMVRXkBt9F6FwO1kifXf/ZPxxKmJ/yO1/FDN2GJX3DNlicJeWBX
sycqlhNpIHbP5xrC0QYzESZ13XiKFk+VFC//OFgFsrZrvRW3uN//4TDuJfFouH6qwXH7RxDX2laj
4ii4kfEzPvVdBOFqHx3odlZJ424Xp0o3X5YSQZrG0D3UXtNtNU7Dj2g2A33XRVhjTGtkEHD5luoR
KEByi51B7mgn1BQSEZnpIiza7Q9H0+bzQ74NZEMABP3RpmZ74NSXEgapqDplhyMdu7azYOXed62Z
VHVKcWeAzHNl1Az+zQLGc2vnhv6EWH02R9wlh45hHYIb1grKY/OvvX74DkKNGDo30f6OZl+g/B1k
65cgQAh+Xd2lElvolGBieQMHD3ltDWc2PUZOkYLu3ivx0VFVI+/EVCeVC+3R9U+VNbTxtPvHq+EP
dx7BbDt7chV3Q1/S2tiYI7OPYnMf+ffx8VNg6Mg3ilowuQDDQbEbTua7hLb72k6+bsQfq7BxAx+H
xdCASWfX3rwOpLUt9LVry1ce+vAqrljnHC0B72n53nAST0vvwlAVEtQUr3F4tSXj1dDgUqjM+vrg
+C9ZGykGVKS9OQargLtZmz+mgDO20REUea2/4kZ4gEZaZrb9X3RpdeUHbXaZoLtM7xy1VvJojznB
9Zv4KWz6QrzmR5nBiVL0HZhXm2dUriipePenkWGqhqn7Tm8VQ71xSKelP+X2nsr/puKv8Cvob8+C
X8WsdQhooSMqOGfHcvdtt85/ERUT31Hr6Bibi0i1l/0w1BDYdKaruwzyG124LocbJcAojkmvDA2B
Rwy70OGMcVa2opHyzlttXTyPM0ioMeK+IWV5DOTVvmO9J2QxE/TifC1Al3seFN+VFl/vxqam6ccX
xQ+tr0uYaF12vLGg6p6O9ihiFuH9bg0Y8worPzDnyAFNB8I9dG13iAG7D6pfwy77tWRQwWDfjD/0
cAAsTuQIbur+PFFePR3Pw1mQASjyYi1fh115SqCb9oTPQtFhyk0NDSqpiN8debCLmywDnlh+NZ3e
D43nL3WwsooZvZh7wzkXwcGd8Bt2AE5RIxVku52F1ZObNicYDdosL/EL2au7+NsdqPu3+GDQf3qg
tqTNZgFrTNv7faKLCYTqrLH1fL02W33XD+H06Ss9y4oOhvEFzv0BV78RTiVfjdb/NIlbDvwl76PD
oDA0kXN9sE244amC4bIhyGKop+u48/CmaIkMX57AhlpN7WAJyinKYUku31jn3L0hrQ8pCvxzCCOf
ahQ0SpUtlN5T6EbAZRUbdmMD/QVqH5V78NztOksYVc8YdfIeXfXY5RJ5mmaAfLL7oMAqctep7RvS
mKa2c0UakSarkByTyRlsjHNno/Re0Dqo8isWZGLHXIT/3QBQZtMbbGed1QEPCFJL3kJGhlBRnqpA
3ZIlAU4HH549imRig8+h/YeCESt010tJQKlEMurWdYcnrs/kBGGZjjZOoxrT11vnl2Nk1vXPzuRs
OfZaNMIPwFHqrvFJjVjg269ytWf3ezbiBToFCGCHd2RWcSpzR6wgOvmy3nJi6HUTDmB+ECmXPmA9
9juGwaVI+o7S4tuOiYcNEogiinmoHPF3e0KxwMycT/mK/E9vb0LuW4U/+ohkE6G2HFMtYy3qCwrF
TX8qaTjgmSKSAJGCqzJ/8hq5/4/tFpRL6N/vG0NQUyt4Juargn5hsbn2L9ZTWR9EJQ2Uw9P1iDpP
kme9+5WAPGO9OR3rZYA0MccGSHZHp1WcGSOczHsnkCxKtgqN6jG5R6Fb0qWSAu9BEQ4fleHeL4hc
6WLHiodZKRBLfd9DAvKyYqGhbVDTZPQ2tJIDa27Lex7dT2gfhEFfbPCaHlFkdUD51rpfnALFyLN4
yShY5Nr1VNtG3IBgdxCPxhHMx7IMKcqL3uVQe8h1m4yvLB3WwT+hmS0760UBAC262j7Bi3ISwXCe
tJGsJqQMFNEyQVJVakrizhOPoFgchRGPoYTFTkz+cCM5USHXJ9wmSKq507tCJj+Dl27F9kd1UJ2d
t2n7SEpn+1+NdGcHUhm95c84dYF5eb3gKFDOrSKLv5hgrI3u6+wucq2QrRvTlTIFDctFbXOzrwS5
yopHF7RzNOa3xHV9fNe969ME2d7VvEf+uIPvOcH1IZyWT7y4Fx3dizMGrYUaJ8Tj8sK15up24uz7
ahP7gEr45CEntS9L6jme6H4jlElux7k9/oCpQyHut47DLJCkfPz6qfWn1Zj1YIJyLlRaNOh7y11/
4c7qUeyoUBEf0Xk0XthNodwBg00v5qPcql9l4xkuGuU/hXNKaP9NsGBMICtgdRiBWPh7Bj7xV5bv
J8pmkHR6zAeMFBvcya8YoleqW4npyyYObqT2xZwPiWWDaePIl/EtkQHMbG0jJMC3LAPmEU5sGUpI
ALwKKdGKLT7l7qYzd1ZHzt2gHxnPoTCUfWMK7YII1gWudko3GQwo1UMS+I8tIem605JHqFRAkIDq
reD5goHxoUe1fPlgTuQx7gsj6GmpX8CL7EzgBWXQcEmX2oLCms5cAX+wVxA8UEv0Nw0+IXe7jjeA
FL2erB7IDMBxm4s2PTIqh84oYS4EasztCMoYuMh8AA/zBx4fPHYjbt027pNQEJeRGRxquJbo8sgI
iGu4Q60HGHW4y6IMOMUhQ7ldPta83HnosSsQf4sw3YqhEyK6IA+UAz/P/yFv7ryrFeTXmtlz4p6y
fdYPTSnJisbuhZsd+8o3XvxCoBj1JCMf1jBwD6AFNRj9bN7j5lfTwhqm3Eu8/hSmCVTbSeH5jRuZ
9N6EMr9kDmjOgfYfq4ydrDYsuvXfDlPYnzDa3pP1vx5px3Dc/haZXbAdM+C8g7b4L1RC1BcB+wSA
1iI2bHigdlJDq1ZqefPQ6Osa2Xi7eKM+I0kodmqpkcwaKxw7uAUiHKDp6B2q8o8zB9QKH8ABXq6L
aoDAR3TFcEMEjJZq1DqgQpEvEOwUlGol2kx62uyH/2/kyiyvNy991vTDc7Tat/5UxrmKHkjE0c/N
JssL/fm2WNONHMtW7r7zmENbHiKwWsfJxl8ozuUfeSdgG9dAP5IzHvdw/NWcuRPaI1ceWMfe6RkI
YTiSAVRldUX9IvDPXlF5mBownNclOtKGNwMaS8KHzecB2ENjxzitv1eihCw0OCVEf4pVpDntLk9P
kdkexJHkRJVsrkxKVVxhAI/qq9dGYiC10sksIpfy0fmnof805uJOPoCxP4eP4feQJifcyauoiuea
65DzKhCKq+VNjsm/3lpVF1vU58yYq9sFA0RoMRTVN3iTepf5VpeFTAqQZJYX32S3iclfZ5jAIvue
uN73Xla0U7dd9TBoLbEKmZhctRbs+Qxgvnfg5W+Zjj64/LnzO1TxVX+7oQU3itJip8WVzczf7HIi
O1l0kWWFyLyJJ55wix7bWs9MV296+stJU5pFqM38HYINlfPO/qzxBj37ix4s+kRgxw1Uww3cRg3J
ws7EvdShDweFCYmgDoLhHg7fhYGekLLd7XucRSdW4QbKuEnfU8SsRV/Vy6FlQ+ZMk9yBEBaKcQHw
52/MvZDSQzgruRr6OgqmUnClPrLnH2toVJP1mCpCmLAlOC7K+E31uhCypb3fv52quBSlUdXEzUOp
h5HMbcZBeWTSRE07x0oEoEVTZ8DHMnXWaRg4E5DAzTcy9dEjrBkCTzeEkAcmpTmLK3kP6m+mQ7se
JElpJP9/i8tGmt2RPx2dZPHsctjL360ixgdrae2sSqeqNZLvVQ8mJggiTUj+ZD/z3u4UcrP76RCg
1j023AQtcVVQURDycChvRsQpIkPhx6RCOoF6r5joARnSBmK5QGKxeNBpHJZJJoA2ypnohELwrVRH
Yo7y01MF6Ihzvngnlz5URzWAFTiiVSt1v3xv4eIHmrhSe50wddPF0Mb9SiL+IHei+O3rYpGn8ucc
AzuxSuaa20Fts8ZaebI2OfGnrub7gFLP3xHsGIrCr1LklcsSN+UMlFgb95y1MmYbWEPFjqdFQ0zG
IgAQsMcHlfnKXeVukCfUPF2QqPeU1ls26WP+x8ovmg3h/c3Zw916vOLA/7mMgEceFFwDv9gkZ53E
Zn8M8/5b+nEDOiqmLq5rMwKLl2VVq3ShiofeD1RZdX6LkrFqNK3a8wx93BW0cGSjJ1ElNTUXl3T1
fm4bIM6VueE7hOXHNJk66K+i3MBV6YtwksENQudCNExTtvueFndJouLm8aRP+WDlKKsOXn2rrVm3
C+QiegTl/4x1gDu9rcLsne1ifQz6AM+9T+ES9GRH8VMsAeh9gKuO9L/nn1cFS957yzhwIl0J20H4
EnrzeloA3VoCkdsz/rtxj43ubj5Um9YN2TUluDgUKltUhsiFjgu8NCuyxujUpjMHD05rzimepMnK
h6fzsRbBq+UJXyh9CPBKjFPFzefipNjs+nuGQtyTwVZPu/jhxZDXj0TkY7ynF4Dn9U/ucrAqfYwC
5EzNbVrRH/TL71n4yLbl/3FvLK0ghJe4y/qp75j7W+jSq7DX8V0lxMnu3GzR/fmH8gzpPWv7PjHM
iGTUbtswbvJFdracv+yqElFKWvbjXIXDAXFOC0Ca3PeCiD741rJ4r0fE0PGyz/3YBJiPL8NP8C5F
IJqKQ/RgnP5iqOy/2dGpRbfha7oo/QIIfk2H//2/4D/wN5O9bwQoAdJQW8b70TTm6ItLBBGox1TM
yAFAYm7R6vFZ5DfC7fEqxQRRovQWY0miR3KeGVVyVb0t1d4WTsgBSDJdfyHsHWjynfFr5/MHN9y5
AwNWuUtf1Q6bOCavQiORvnyWhWB00OOIrXORg6d1p1WMmk++w2pbe8hBi21TV4jOfvYp4hHmC4t6
3MI/NRGa/JHmnQqKw0aBSVnXlwtwI7ilRRVBtrgp3QFkFzdaX9s9u3nlQEk0FqiwJKeYp3IvWXr/
aBYCYi7+rDZJKIKGJwn+Wn2qLqV8VNhx/7z/jG4G5b9RsRi6wgrFONjJg2ktjbfxL4TYKgSA1XvV
y8kr+4hczYe8bdK9fwECHOzJ7Y8q0mBr+4Gyr/gt82i/KGMptn8U30WBV4b6B97wDzm9NEhxQnOu
ti+RomgB404QFLEDTFHfVYdbRf7XGFdZY4EMvgSgL46j8ZV2PjwRbNCfRS/DdjHNzvb2epJi89bi
nR/xDtSPR5CPl2lLMTybVlRz76FOW1qlfYX0A5wqBxFDV2lQ+cOmiC1XRSTu8Ax/M/tNdckUnc2R
z/IhTm+OSXN1SRhPeNI4ciQMjIyDOMKw7Ww4wA1sqtjWUQXTLP6Vz6F+k+oK259bKcLVOL/8YreW
SD05+0SRQQqFSJdxhglukRISypIn8v3jOlJUD0EQxMyZorCnyz61n1mJaQsMNrCZPyMnNq+wMinl
31fUvtsDDyUrQK5GX0V98wKmN3pyavgQ/XeIXP+Oj0tReO9aJRaRiZ5YHUyDst5xFLR5C4cGuvYJ
ocRx/IlggzZY5JxI0ZDi8QkplJ/VL/y00VS6OT5boO8qD1P22/u6U2ApkGvupCUWoPluEn2YvYWp
ZQzG/cwxdEopsEpU4i5ittkyhxbDPckRgYVqykMsZWLM/rUXFrIlCHAzcG/X377Ig7qQ1zfInWIr
3tgOjQdyUQOZWrxsv0xGOk6xqaxAD9hVcHmo5ySSOzMhrfAv+FA8Ond1kciDcyYhPKJ35nXO7y38
E6uvMKmSaCLgZkhgckrILzJXAlT2JBUqtcP059jiDVGxS4I00XdztY5vtltwE4pAXVmyki0z3EcR
uA9+v4gb38J0sqiCcxVQehhMyTO8O+7vp94HpkLjeQVvLRLnm46u41z74mC8Sn+NZzR4YDZl6+cZ
p9ESE1tc946DA/zECnCJ+xUYtey9JzJPpI8hvTkFS1+U5V40bsS6krrMZNFhGstNv5VT8cRRxoy+
F9wqPqQS+vAQw8bB+ZBaHp+BDsfNEsszizEBm2zhi8NRKz1xyIIDpSMJgxrsoACZpDVrfJs/hOHB
37QsQ9cBPpwI+ijee02z0xqPSMCdlD8CnpkauweGJkq4VH//ZyWifti4D+bfZJdIpagYl9m1My9+
wohOeWWiyXd8mO6YMMnpP/n8qK35/N1B0trlSnM+BdHwCF4jzoe5BgTyk3G5H4S9nR07+VoJSgxP
wHl59V1ZK+e8vyCo+2yK814Ko5GYNEolMO/dTv5IFynr/Ifrb8I3HtgzGt0Sf3p24nsLFGI1aBkG
AyS9PbAgSJfHhiUPsQRRtEpSuzXOu80jEehQ8T8ZjWl6endYxCBF0iI6GEflVOmc3TXljzLTTcQH
rviSm8jtH0LbE/tTxNHvNjNTfMtJH2VJP4VuvD4TkMzoK0hht8CeqcoT9T4vo3GmxK6nC77TryU5
bNeJBjJwnJgxfJLY6HJOmxH9a9PoJoBOTsGpI/K051m2RfyMLIuIAv95QJ2+qIqfoO/Vya9t+Rt7
P5Ztvr5QJYqqU/zRkEY1JEva2bdATitDTCKB0FnLVNJsWYGhkhZDzQUiLurqmFci2BRhUOQrBjMV
ZYky7z8K5SMi3zu4HIjw+wJA1If1E/Yo32cbtpyP0nZA5rN8gGhiwZwcaM0XcgHnJXf9yylKxQqb
peIkTutQyOe8bOSqG4EmNu/NHOBWGxCvdoyXueJ36jUL1XoTlESopuekqXch5/qBUO/oa0o7agVE
IiX+i7gnRibpBFqbcIrFU0ST3oxgW8Mgcx7szIUCFft4x5KGejbkAT55w58gyCZc7S7fhVYTqF/I
KowRfy9pajvw+cFvCi1z+PBGp3W8LWZway19Du8PzM3KIBlU93ZWMponHfZqDG0ebS1EObmDHW/b
IMupTpZAR6mcS9NM1gHix9/5zXLzhzIfh0IVoHWLW01T8Tb4T9HwhubvxtNhkTShl6Xt7RY0TPiu
jRuxhTpGzREBmzsbQB2aWFg6xHmvVHGbg6oc0mGTbqMO/WaemwC0MN4zQZOXMmAdkWj4UAMorRaq
m2sVzFOyIebupC0LxhcwCTOTsJIIVZolMsHc90l1/sGTT/hToBIqJ5ph8YacFX1BnNkIFL+Fxg3z
Cvpn25QARm1zvrBoi831quYHhWEVkV121JtErbqndPWHXQkU9AoyUdJ6xXOOqBtoIuytHJJT613y
rscCitbOF+s9/5Hjaklnzy99m3Ar7yCaWFCzlH4+Kh1ufmlrkFpxn5haGVFShMvprVGiStQ4SkjQ
POz7UM3WGv+tyZ6BxjCFzzIxIg97AxHdyFGBeDhn6QDGjLWnQ61ahIToJLjZ4QnOuhfcRgv2lDcA
GGzYv0Y4nibqLv9uw8In8NfTJwlYmxQsBw5hZSfvj1mKqu5zG7PnHvxVc/UoEr9oswPU1dPoShhp
N6nxIohP624E7CS5E1VPfGZ9OPUIzpmjPNOMQwv5+Sc4CR3h1z0ZjxcYeghUtw503Se54Eb/x537
3FNL0Cd0UUdGxn/Iwve9T9Hu2dMnChkf30Wdb9klUQq4ICu/rFBBBmHM1P7JEvtcd353QEwRqsZb
psgAtCkgV0UeI0H5WMhP3aeDAm2RHZGWpiA7h1QaV1nEG98OSyR4hzL5v2jbSFZPClAipIT2keJJ
3NLbL0e6iF9Bm73MnaCcbII682CvoV3sK8qSdcEf40JkjmpqpOrSZeST4u/76/uMwZsrk4LMP8I8
/hZEnL0Ss7yKilyqodY78V4AzKc+aNpXADGiqouhM4RMDqeTBdX6R9XdNfe0MtX1XujFGDdXHm1/
VQnVO3moMhY5r48GIPFRZ9nmnad21yRo5kCZpYJgOJZ5jINqrp8zkux+DAN9HoZ2L1fKV7i4v8OX
qVf1d38SewOwHbg7orEhL/IsnnvORobSdaPXqJb0Pl/QFr7DkXVVTAf9GqS2Zx1bwu/ieel6tmsW
TEyJf+fFGC6OI/yBIWbWqX4r8RNjKG0Cae5wJRkwlmcMpozbdWRBXQkF2SQy4cnbWdwXifQ/Tz0G
V9XCzcbiqJtAzOwh7I/60ENRXIgs+LP8Yh+3McolVeZ9rx+7gCfmkshHgVv4yqefJcu6Q6wPFt6D
PCBoDx/fGv9jf0XTGya7/X8lkJi3trhu7Essy8N/yz1IenBtxZpa1ONqwl+ThG1s5RxDkv1o+u3d
J1Pq2rZJfytcPHLhCRKpdSlmp3iXt+L18qPBeE6Cn+gtQ3sB0uA1etpd98hkgRyR5BYgHJM3vTCt
zKQMD/6eyNZDdBN9e7KzoArG2ThTg4KumcQ0rN0SCRZDq6t40U+9IkwRIb1xy3itD9s3sYCsYlKY
1yGfsBELeFGGJVN+0BooGDeDaCQ+BEWR6XxMrRtu+luA4OBi3WxirQgPOt/xejl/39qjgxZNp/6L
YrdmtEglHT2s9Tqr8s58jQLpYbIJhFAebuQLtmuDtUZJG06IHjeG9oHWIe8L4Z0Ui6IOEBKlYwH4
FEmyWbe0lYz+v6UnpJWu96PSEx4yOA3bHKPKONcKwbQRsLSb1UNuVjcJOEfjZFqX7UsgaCAx8QGz
0z6x8TGRyUB7FXio85/7ZnnZMTcW0yuMQmGXlWwHvXeoxcrm2V271elail4ryFzTVCUEgK8gDXBb
eA3V7ycGl6ykpCKgtzGirp2qoRFJTxn6E8+ql+0W74J5XrYGy/ChUr5YtBhNQ1ORcJI9DOaMsKS4
IfhZ5zYM/qur4XdQThA0ygKK9OVzpp+sV7RGg4gfpO7ET72M4W/Z2So4q3m3+asAyFE+B7zWQnYY
fCyjWAsTsgVOjBiysHvYXkoQ/a3jcGlZzFTREF84PAuFHYBCe8iru/QA0Qbq/A1lZ+tipmVZIhVt
wbXILPB5njbI+4a6tOxJBX75o/6eN23zzVJZWy3mljquvtluwpFnQDB/nU8ZO5DWkIVMWaAW/WAa
JriI/M1GnXd/7OLnVcVkTCRx/6l4NonfapcIv6Go7a0b6MRAIIbNFNfdZfeHtgbesuTrv/6dt0BG
FKflIIt+nypvByvzRlaGymNwsHINQibRJVle2rZ1PIsh/fX+c0+6jqYr06oEkock4ALcT8d1qEX+
DfNp6R4fLk8OoEUhWCwV8Y2WKAxfyyDJF0V0ZxExoYyRJ1d+Dj6rHajWpj2fJnRPCmTlfki6Swss
fsitoxfkOrNk5oL5y91tB287WT09BbliESuZWmQzJjhki0UJiWQCrJzUwHLLndRulQwXe2lDK3rr
/9+FKzeYoOKKD8ry0S0XQr5qiOqW6fAy6T1nDBStxecLXWNujpdPnqMqt13fRVmdbfZZuGBDsK8w
CE62pFeu1QxCEachKHx180oP/UnLoDS+AVNJpZ03GMd0D+rgNud9DkffoR13S6LCLryyS2jOepHk
dgp5T6a64DxBtMg9B17xkPQQZol8T4aI0EzQgxymY72RUkLE4IlGxkAA3oXeFgXtP+YgJYrYiItj
RwELJsQxTmqAnEu+tseBjus8un2acMxbErvpnNBW9uZrrOkEHeaKCtfhHwu9wCTs2cP37cfqAV6I
CDO9m9ipXP0f1+voFMINtiUO7mGVrEK0CRoNhkwrluT1Jpcb1SQUM0Qo7JBp9IZ2YJEgLn5yd2Bm
U8jJ+hftNW0HRyGqcbfxTONw+qh7DJbol5s56YAq+7dabF2Ij1vZAWKgqllZ0UTdPBN7QXL3rBc3
7Zd/I0dDnKQnMU6kp6/awbfwVhq9hjwhxrUJkr3d/LZK6J7mLltuI3EKJ7InzgHTsaKZCgtLUo9l
HeeKK96Wkux5f1Fwi0PrQdcBfKgfRUamZXfTG0enA0eJI/mfRlOqLiKdL+g2xSO/rdCEz2MvKo2V
44k8jZOghjnP8tTJzzPJw27zk4jVEhKve38yO/3ziZtApbymnipNORgmYUvmviQWoMZVXz0CTpH+
zqrNmQ/YEBESkKgwwIn+M/jEmdKuWr+E7Cxkb0Edzpz800B311NQXQBVPqZO62Pyzyi6xZnVO90u
g6XXa0CascJnziWCHJOiWZe3eAa8AxZ4835QdZDZzQCCv2LCNuu/wPo5+FWwEdC8puq8QKk2OKm2
tym3+x4vebt6V+LB0AnptzYGOj1wPRkNJwEi24C9ZqLjudObI4P9chpazvWhFC6Z1mEf40iZK8Rw
gGuDqg9ZlPKdXZWxYkB6y8VmEhCz6bgGePqj14orG2imgmgrROp6nyfWATNTGTTBVzSPL+fwooJz
Xu/nj/MZRU6KuHMZNEg6VqvXeGitcN3Yq/VG8sQ8tJejFfK9RkWJEiNbTvgtPJN0zg52IVFestku
M+DT+GbcBD/3yIjdG+G5vYUrqCK7I7JT/6wgRal+C3k7EML8Z/EWn+/BKVefVFvMYP/lTpUYw/ms
qbnWI9gKU0VzhhRmnv/DAKGUAbGbhc6ewJMY6SI5EjoVCyRA+5t3EywUWa1YQgd4FImj1LTFm+V3
Ot1SgYZjqFmC4hcDfRSpbnYiSVKC//gxNmld7juP1z0fXOt16mp3LKB8EOd8m20Q1PJewSJMCZv5
lf4xPWo5bVbPyi4VCEy/e+CZv1Wa/hx/XAWIw0mzV71OqhBj1mc3zIU9xGVpdvRJvTZU22GNn+1T
T318pL90AGFX0DM/udinhTz5cA4neV5IGS8E9ovcGIrmXDGS6GwXIGzNdx7nratAyrxYkH5iOSAh
J66xwcdFBP0/Quuu0ELMPU9Lh90fE9DE7kDzKp/SzGUUuJ56dax5EB3jNpIk8G9xpVMNB5r6K4Aa
qGZeYZTmSYXiWqZRZTiljI4tuRtnjd7xfl5BWHqQEnxRgGJs+wg9DAOYsXPTSffsfGnhvNyf60v9
LFEryVM6GySD0HFX6o2BR/P7pVQN1M43GERGl6LSnETVticJ86ofPsecFxdr7sr0n5VzzSn01G+J
zPg2PXbtAsshZE2VgKMN9NZu5HQbTIytEHpsQhSNuD3ADW27OLj/Jw9seTRt1IKE+A7O5h+pICNX
TkcA/iJRDzIFy2InttUK5KkM5VSjP/Pw30xW61cMN75qSfiViSMxI1w86HzC7deop+agAIydN8Ae
phNJ5n7rzUM8yFxRhH4q6J6ty5yO1mvlKqpvTkvhKGEaUoN1+Jo851/HEr9WamNxUEg/BxJayR8F
E9OPXQhjzCXLLPN0mQbO/WKdRDmedJuPpPg9F1/xOuyyfEZ+ZV6hqjd8onBbtyU2wMzY1ZYqwUUF
41r0soPWkTt618jmEaHVVO/tYqq/3ZH0MbsVR/A36rPsfzv/Utlnw/ZC/CMdRI/FNdhJ1IXT8rNj
Cfa3vPMU6rstPATJh1PD8TKfCxi3EnRO39oFWH24fDAVdVW6louE7y2T9fJANfUciD1dyIStFF1R
+ITX1P91yLchgvU/rrls6Wj8J1RjfSQ6gFw9+O7x/iVi6ocAy3C/4QGTrQagZ6Ct/cWROZnkWCdd
DfebJenaP4thdTX+mkZHmSAVimcbiKyiV2lHSWSvdtxDMJB84Z6cTmH7zMWBbGMynhyigIDok7/p
ANCBF+pbd9Gnl2+fFv85pbFfuuYQCfGYFJzbOKNO1UE1ORugpCBao2rccqaMC69qYm0YTG6wq21g
pBZaCfHFwC7kWSpMEJpHDj6RdZHuwQBEFpeqPXepPVo4Qo2piGCOjnG47Ak/hTJDnlM5+uCl7rBl
ThrgnsiJs2zDasOP6Pq2CUpI/3EmZCtEHH8kaBK1Tg4HSeXB/KWIKdTCbhLW9v/WTuq2lkVIjc86
3r4WhbDgz8plGUphkTLV2nLF+dLWlV3U5sLW519vc3EDOOBuklsqDCXNupCKQW8l4HtjUIu3ZFgp
vWuOHUVoKrTuSSFoiTptGsrTjDx0if5Nx8SYn+tdnkANUecl6ov1hG4sYO/t53zKtoF+CCpijvCe
GCiDHBIeivCGy2EEvW9lEdUj7WqcelEcCMIZba2/ZAdZdyKs/VsNu/vr1cnFptN+fH0blLhLxVW0
JgFtL5JXcm01Znlpb1UTZLwb6D5tQltvTWRMF1Vj4jTW0jjajvoGGSQWU09Z+l/6efrjF01MsJnP
+HYzfFn25Uh8UBZP4YF+jowKWyVhAwvy9Z24wqZC3Bl2Z6scsQdfwmgvbTsoqf5kfGq0lG5zWsrc
U2EcUErigaIuFrq4nPB5XLwpTu8nuv3yjHXQK5VRVWbGfB9CCDw5M2eAwH1jpcqaXUlfGiJ+1TCu
U8Ygr8jqinsYCQQ/JK2dwBD1/HLHMO0Cy2EU6E2cpQDICuAdr76+QruLYoKcou7cT4Lp/OjuZlNI
c0CF1V8R5O1Xh6zyelZcL7pXq8owmiweTT57Xlo30klqThw9U3UejHw8gjE2WLtBOTDgKveZBYbL
1kbsL0UsXrZCP3SiE1q/MozGj2iyWQIVrUyJigWJQaPYNu659ARnch5Jk0ke7pFYhP2i0K7ZkgZG
vZZElUC5VYbTasqiIBXZD+IOhd9L8Vvs5dvekJWDosOfSIQwVZ+4l2RR7HGiytgAGwYuoFw9ip5l
3Xo1vgNvvfp8pbP7UauCQXABszOrqVPYJsI3gApKzPgTAPu5qsOChaFE7Vl9681+HxHJKAk56h+B
vxZam1OZtL61Jp2S/UpiHUqffXhhlXgSmLLUXEf6FqQf/5MBH8rU5cDkh+xkKl+iH8tjpwtoeT37
1sUTQb8oldVDEy+S96czVz6C6ZXqsZ7jfOc7MlxoMHUg2VxQZk1393TauzhlBi0MOSigZGbNFEfD
wSDyn00nPu3zaWxNWhJ7eHzPDPAldrTPLWBozWagtv/V5/7pz6l9kmS8N4yrNcGu+g8YMvyLHAQG
7lV30S+HIDZddqIQGyzCwMqXbWbPO2/LFZiiziHcTuCvoPyP/2kqzG6ooTgF/vqVvT4S/gCq619c
wemkrkWwQwmSndMan1DsN/8IGTKYQiCoMraTZ6Oo/onrrePHtO3yk+Q132XuCVV72kNmSyNPZvTo
HIsLolilUKexudasb0LZxmlJtOqd4dYyn14bew67Y4Jgf+tye9i+lbdPbCEvHiTQmXPPGo+8fRmV
qi3JTrzAMKx2XgLEsnNZ85S/xxqTCjvlgs9yg20doTyqDONo1R9X+5r2K+RiWH6Isu2rGeKoHrX7
CJdyEze/HLqmDAyXEz5N4xUIBPWaGizpPBpJpM0UOZnF4X/8bp3tmVWlxeHPxNa2QEZgxPiuAPbr
cgLDRb5Zg9UYoKTj/ENLZN4nQnm49x2l5o8SG59oIwUe/MwJS414m0XQX55H3mT8XCQmyBCp3emr
Kvc+ShSYtTi1nQp6oAighN+JgLiYg2I2eZBQPL74B/jwckjOjhl+PCSt5gZulc2Iv8CLvnnOLoba
tyhvG1Pmzf+fuB2G8VTt6itsNrIra/etIcK/1+Tay/NDaqtfTI9n0ct1s2MBKpAlbsiYc4Qkuz4v
4kAAxpb9lHC4UF5uFWhi04noG/IelU5dAZD6x4VCb4vSHkLqeJuvqMZSr++SYGlZDOxmZLOERY3U
2sm3ulZGywygAriEGiLyQqw8S7lUFuJJO9wBm1juSEXr6Z8Qf7c3D4fAeAmr7fZ8sYjp+7tNAZVO
TlSFFaruq3OeeK9fJf4m7gIcIr5RpCbmQy2iquTlcMlw05BZoo2M1tRl2o6hW9q1R3qb8xuZKejw
yRe7Sd7/Ggj9DQMYZxDGA0depO0YSjsPQySK+7S79aVkQhM3f+2ygrSirSi+R7M3o0LmXrpFLrzN
MY2DEAvWJqvxTSQDBGotKRix3dcmOBvVdvjTD9bfRbVwDEy+en9UxVRnYPWpNydvDhtju+70RGw3
rEAEPRsiwqpwQTY5QbvcscI5hJofGHQi1M8VbOyEdYBrsKRurql+Q+F5YU+9XFe8AKYAa0w6JQdb
AJQcuelWTe4MF1hvvYqSFecoSXEEIApMhqJjssehVg6Tw5Pfos/2LYiiCSquI2CRhkMMqjpUw83a
i3ESriJfgJGWJdrfnNR6EDIg4nL/b6kOcOebVzSxGJaR1RQUIZdm+s6ls66W/j+6CsW54txnzBWA
f03ysf0JdfgYS5vFBhi40XMUPZUTrVJl0SzT7j6y++gfF7y4G2LVlENHjImsogTxBf3i6FzQHrrD
VpDh4Pag2H+Dz8fVH0Av/v83ALjO1r80y8YyC9ZFN8kVNl23n2+lhlyfnEqkDBlLkuyYx9BXjh26
3RL5saQlztRpA8EZ9iYZIUuwCLlB46nFxVsCtIsNrwTjLHBi6CRqJj92WUw26k5hlNTg5sCpYRMM
gnxYd1JRge+9xLdVRt1T+Ds/4Kie9if3VCtoXdp6t35JMuca0yKX9ihz/hOWZLzQ8BYS6Y4meit+
uKRvkLvnMBZZ+KLI8LOG7PxAJQ3ferC8B55DXICW4Qsi7ZIrBy5T0V38C2ACbcwyuUXjnUwOBRiL
JtIVm4fyX/Ayne/AgD8yUYxjfX5kXPhSRjV65it1TmbDlqOZ5/NMJWTH6gXtHKQVoBtJMPdUMK52
I3j2RkjdlQpXho2oGRPJBhpWUWVDh32qEXXVdSc3Pf/jzJ0rLY9qz82Qra5BaQl+mmtlXnIrAiy5
7UAScRunwhlcJs8tvOOw025/9MC6OlKQFX8NI1y9XLY+CmO/7VOBEc0oCnWBW/eCYb6kRtIiaPRG
wX78dWt1GEhZmMtrbyEYe5i6op/ZF2b+Fyg0aeOJsLkIzAA+qjac0gxbzlciU7QsdchRE65svoJn
voSF1Gbv0czpjPK/AODw/mlh05fexzj9gHb4tFqe5qKi0yjHGTXarU9jNUIMvIbJEgJqhJLkJQCQ
tkYpjgkAI7rDme7uyz9G8OgYkWuEhaPUAanN6yugoLpjURiAwUvSoeRZBVHjT+x0I2mDs7TcqSNv
uROovsQSeNVlkITB9ioLmnxw3/13QzFWg/CdB8m0Ymv7bhX/Rd32j9o8sy4DS+HD9Y1EVYijQvD+
yqCqrtp+TSVLVBC/UwbM+EVCdXGv1+04QJN3nj9pw1PMIgMtF8xu48quOsTrkmmZIDEtUEi6klF7
Ftfd5p1ZYLg0WNIILXYbVASjCzefMmr89Fb0tBMuNQvIQbQd1fXnBitd0ZFtEWWgmbu7adlPNzdY
F3DyIlkKJvV1vxemRgls8PtOA0hi7m/siGUj4HKE11Y0jrr6a87pqNXfw7lFoG33LettRbQnEafv
ZI/S3WulBEd3745GPy9d4E28S0tCPE+Uvzw5092DJeq6kpB8N0JPhDJgQrYYOXoBOA+LlwY2AJp1
Kfw0pz+i7/FZkiOIhd6LatcKdrBUBa2bDzjaN6XgQQbEs5DlzCGCIXNcfo7L+KM1R5GAftvklFk4
sPOONexIb0o5j9b2N1UKOR5/IqaNKwUceauRIkvIpJ3YsYQd24yY1dxxT1x7scqCN+jOqjleZTn3
1v/f2nDCLu5MEbhetgIS91NqHY9ZVFNE3oIbmRv2452vdjqhhC2B3iDWs3ciw7cItiLQBsUu+keF
SpZ8YOYrtxUf5wA/vqnM5Tc+k0Dmvx9hp5YZqHdgNuoecN+fBO9+rEKIS7gJe6gBlhKVtS+O/yjG
0xpROEp6da/EFBg3mk/GEuH2kCKXz/B+EJnFOxGTvGp6WK72EuU+SzPLxaoqJPSeRFyP8IlCuLlD
Sx+QIOMoCMjmHTtY52DfJGKKUh92qQ2S4pTgxCPb2wC+IRbrvftaa6cXj+a7WQmOGuyUKc7qrhsl
XCZsW7yumaA0siLevKsCWEnvZvyqLqqST5+dOQiVpy1QFLbUihqID1EDK7N+utVtA05bDUDDPlpg
rBcfV50TekGBN/j1O0X/BH/C8an1qxeGIU1skRkrzrPTKkzkVuKSEPfNC0WO2swYa/nOdUaZeuv7
znjDRXmXVrkUJzRgsbgLxQQ5GCzfZe/aK+FfGW4XZsPgF7CaqStA+dfwTMuO83CTogkACvkyoI0u
sigVZwojXI0ovbktO9PpCsOFSlRQd1U4LyAPFdOOLgU3clVbTNE8C/nHRJb5ptm9Sr3fMk6DKGKA
e5W/g9FWmyPiVWWQcDVuyVer6EQJMPXtgXatKm7NeirqvhnjG4VlptxQUwayvavqzldIQ4kQ6lXH
ghk4rRRMRFr/DQrChnrA/xa6l9DDbXW7g2DLmDcba4F78XVBCwSdljAX/UmzJPznLLRqZQro7mPK
nDEH7ORyIvLGzVg9i3X5SbEA1dE1OosX/Iqg6j2rhhh1a2UvTFs7kWWkhSKuIju0nff1ulREvqOB
ytv4quvf95SdIfHSgKI9aVBTKISaV8NvZHUVnRad+m9elyLiZiRruRicz0faU0o0LrqkDvLsdZGX
yS+F52qLv8QW+Amvb9pBqelLrNuI5NKnp0UYMuJ5w4YKceHAdIpXlIuCbliQI7kvYZ9ytCU8+1kF
92CuUCLmIKQQ33YmA/bOchkWEGUMJXv8atrq61NBQyI5Yn+hTLJWPPRPeDTOX+FJTMONPDfKvqat
fhiWD2V9tm/VLzc6C0yko9iD1MT56PonwU4qz3omToT3S2fes+UgpBeSzRipeJA+Y6PFsgVmMbHp
pSH77Kj00qppbvGbKTCtkPrV9OwGE7F7BGpKfHQpOzO8BVrC6sBiNU+Rm7WlE5SXzm+rZRCnobBt
b3Fq91L5Ogp+3jawOQJ5zNppt/U2QcZ75M2+ZHd5GfsytkOT8/oS5clrkaJal4vS+dNrcXv7140I
P63DmCcXGw1EgUHpFNjqeVVo5W0qPfNp3DhOzabLj/60d7sARGzw5SDQoVOLRf/3E1R9bz49mnIm
9hYMu+QdCH9PLwdavkVP7q6N+39XrKJFNOwOJwEbwDNxBrkVtVUYAfWqLRourgrd3Xae/2+C8Tbt
YZnuYbmvGzLYJD4FX8boER9uYMxlPkbU3vX8f9bUUQ7B1IPXUeojb7jvujnPYMt7IR+VMhXEKVEC
VBg1ugDkJsEQ00R+hH5faEHScmkgzYhcAOadDs2uAV52PdUBJpzrGOijLW7vFUczvPd98/f1pj3E
Wd1VJWTloOLSGrFjtLksAFDWRrdXsaJ+IbxdRTgGQUgqP0MufXZhB4V4F0xPG3WcJY5mHu1c+Ruu
YvbTiKokwsmYE6/+PGrvZ2+qxabJMXTtdMf0eSDoLYdHZruyoMIUPVBZekqoLTGG2TnMCtBX0NZ3
Us3kqwiXjct7F/9+qLY4zpXMXYYnacpW4lycxWMYxnE2+2dtZYoeHXhKqnx3/2jNTvkk4+R73LXq
POFAhcTu2Fw+Ooun1o810ved021IwWPInE2aYZEdG975Y/+fKoONqnti1iPsP8bZUouxuw8hb9yI
+9DngTQ0t3iZS1G3QmR+73RAEXX2Y6TYQJxSA/z1y5C3klIq9GwwSS2e4xbzAB1otCv3z2iCwsc0
yYDouf0YDi5uK9nsuo8bH0OomW+z7yLnG3AXEspLj4iXpfBW8+3ejVKgLfB5zQ2cBlZ9RjO6FEdy
GReDp6RSRSyxIRywRUcJgPDxPUKzjXFLtiD1cXwTUMji1Zwhu2Nx6M1ee5HdzxHxZ0Ql8tSYXhB3
8ODHk5UJHqua5quuX5v4Jlktx0zXk/cvL3Ssj2BcmTnl7Ld0lJkf3bOKGRM1OXClAFY2Uwd81Dnb
99QgQIV7jPgQ6O+UjaylWNemYrnuuooLasjhr5rXxadDVdmyYoNqPqH5kLcANTGP2anpo5LZtCZ6
HHYYcnic/v7ndu/xSc1bY0gwPKWWmPN4uhjLl9xL5axrrKJ4JyknE+qRklDCjMqt0Yltwi8iAxFl
ged19J2J2UvbYkdiEF6MWqbIAuUw7j6bjo2VXO/33ttXKYK6lc8zbYEK0lyhxsRlXV2MqrKm4YO+
1tbLo8UBQyyb79u3sTTTwV8zWlkaHVuwBRWMTyBGjMfB2jRitRRdu7o/9SKt1ZltNtR8AU1mO9TX
C1gEkKdWM2hMzPG24O3wdjGsJdOlKzhEahrP8ydclimGoJADrKIzEGY6ZnqfWO0eNE1BGf9jUqf1
dMvq9tIdMINme3vNfeglkxVQp3B74avUx1BikxKIsjA99RSK8T4WxP4wYs4N48QSWY+lYJ7XCp1Y
AmliHjzgtCyUGQVoymGGQf7DOrqGCRPFohdZnyBJ1kQPxRcWdk5Qs7qsQuxfa0C6IQIKVcleQJ8Y
wgIoE9g+O2fq8ieYAYzx1txsTI+cycK75i+JxOfjH3jBAVgeyH4+dNj366TSOon2MWvItjlxWZWE
yEOAxUYo0O25bqqQW4u/VLvDx+NmfTvxD5oLvbbL5tv6QmxtQqB8aeY57CeZWC83AXBA7BRBz5vF
otz2xFx3a8TgGmicAOpW2TaMEH8Jp6ZBID07PcTPZZEh7BAO8P2f4Cyo/eNNPcQvmUG1tR8FJymO
2uusumM3o3ib3Knn6J1sJIRb6Mc/VglxkPWuPJNSlFE0hbp+Tz/mp8z9AW+aruWFkzCC+k8mT4Zw
BV9TkcBqpXP9h7k+fZxvaoO8PzCz5tC2E01oU6Gwi8AY+6N1SE14Yw/rIzAhjIlrDX2d9IJ8zs4I
59mIjH29TNkZRNhej9y5nX3/FtDXXagR33QB2k4gDSvqJxuFfOAIwO+EtuzoDNiddsGs2LSY5pjk
GOlL5Keon9lWlAm3mJ9UMY8Dpz2MigLdWdYkSNLGvF4x1AWcQfya7a75nDkSQkeT8ek6RAzFN7Bu
Gx1RbVqZ4EbGRUtyCOaPjWLKev1Naancnf4TgnNEHmFv6X5bXEJA4MhmWb/mhx8uX3d6KM9iZC37
VS/28e25H8Bwf4cyvAkfuHqUvTITEpy3axPIHrkseJfg04uzzZs/ci13Chs+fdpmWHgtaGy/n710
KMMOw/hc47mrwHGvzYIYKfKQdRpVg+qfDnSfdPwM2X8jh1ahgARZJdOgDsZqqR2gLg76EIg55yot
C9O5U0KJNizZGJI=
`protect end_protected
