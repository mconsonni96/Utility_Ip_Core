`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ZbH2Jz1i38wJgNaxNfV+nhm7Xyv574OMqnMpp3q0rTGiHPpEV6M7OoKsHbIWUI/tJvW0molPTRMf
ORfarQAlepHERGKXpZ8H+XNJkLh7z1OP9uP4+RT2OnYMsqqVf97BSZzNIt8P27gK+eQm3PXkS+XQ
8Rm/iW2SGrwGTrbIulUDmLo/SrVVWy7CESmmHfymYhI66xLDgURg1KLScYRku5GIaZnwDaXky6+F
BR2IElIaE9ZyxaHxR9nxR7YUllhejvxYPLWwIbX6leXagliEJVpmMVslCkm1/hqJhyY8H2D7dY3H
keHi4BKRpJJ5l2d6ptDWs14gY4akVpeBx0agjA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="sCVeH4sZk+y+b/3aNn3TCyh5NDORSipwnUl2lG8bccY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11056)
`protect data_block
306kLAEa54M7kQiTqV8SGsyuaj5HvVLfYyKChRja7p9jf7t7/WUciuDWIF3ULy9J7C9YoeIKXV+X
hcWqhD2K5YeDjZ9wmEswTVWqN64TJV5LzTgAwhZj29oYJWc6i6NrS9szKxLwjGSn39xeocbq3kBY
rE5wJbsfP+uhdJcom8rclX/UGQx/lYLA9gr55tjKwo2PLsT1vtN/o+qOKpBJTcKB9g+lm3lfU3bF
wH69pity1eddejvO9/JCdFW313i+3DlO3N9qnWtNCJ74RwBmGhsAFvnsgTCDo6KQisgXAOgHECkW
EIzpsPQubK1Yy2/8zVIecpoHqzt9Rwr4paNsILSJKFasmkZMNQKKCi13Hi5yOiYyajmY2Gkn9528
Brc6rfpi5eA3KiJHFC2VcaNGDXjNYKuStzh/yskBFhQWNSJbdevNKNobfhxnHfwLeYbfZMqmAQOb
d5+wXyXf0VfK+6pcOJnqkb6oXIA+KkvRkOHkLSKAf3AdBcTF/o5m1O2QHa2m/GJNW3ewrVbKtLLB
DebLVSndxM3pIIaxiQb2UzbA3s9uGRCRiW+EX5aqHMRDlqrqTsxZMZrLrA2DVg6VWMDnqxLQj+re
lgMeIXnTeINf5jEVpkh2PxLj12zu6XQYgG5piIjXh1bbSVdrtIKCuV64VqNfNeMAxs13n/ULGSG3
8QwW1cGhKQVZdaV0Wa8/yk4VJuaL/rZaVT0tO5SK0LSLrbmgsi8qKOdghKESAnuuw3WBcWEkDvAh
X3Ueu54gpGkJnb8UbbwioLC7ooDLLp7ErNTmHy0Jov2dnuRb7subCrV0KmizPtrflJXRwYkKu7gO
q3A1joCihKI3bI2HxOveq54/j3sr09UuKHYrk9f7MDQ2ECfhGxpOhKoOiHX7drEkddb1V2gamrM8
8lDhDwUhDiUf2flKDODrgeD9/qkNIRREx8zYsV5R3Pev19FVss6JkCG45qmgc51kDRiQiKk6vxv3
ETHl543Pv0gOnR8TXTuAYA/DZsslsdvctFcNwW9GrL5uEzs5MhFIOeH1W2EW9EE/NQEFiGTeuH3d
SUvcALFjgIMv/MDytMd5lX3ZOKBYVUBXKoOW6aM6GYvPufho3t2h2PpEDQ2FoRuEvQHRa33RNcjO
REcv+PqUgZptCZFf//3pybGuqsjRxwqwkmRN8lLApC7VIMz5lrt7UgFHq0EwvYbJiSzUbQm+gXfi
XHRpNeZuJ2poMlieHDLLzoWUnK9hL0Lc1SMhxq8E2NUVx1N3N6SQmIw86l0EV4Ud4Nxg9BflFDjC
CQXdTJyhqHikzDUJBlfyQh0lO/jINIxI0uwboe/Q2Yr030g5JNRAdar1wLg5nEJtA18If5kUcO6J
nKe7/t3QFs+NdlFcmS5+x425aQSg4XWSquXy7zg45fY0YDumM6ErhLydAHkj6a/6kiifNINe4LDp
dCmiKnsYxjXYD0k9E1aO3a/SeMP7xNkH5YW4VSq/zxxNzEXpJ9EBleEX1tWh1JIL380bhkKwnrY0
VJbJqfHw5k8ZwBq63InUIwRo60MSgtzIDg/y1v3K51QKdVPjWiVw0krrflnRjljUABk/E5umhexU
Z2BLr5fnHfvmr2KycZ31QRfh1XmL2aFFVU26394/G9oDUT2kyrf370RRwbAdTx3bD61ZuAoZkflU
jSrFHXfyfumdRC7PrAJQRETyiosmd41z+OC6On0xfviZKxIvcvofr7FCk1j58qaSEvV02HNVys/B
mAylq5iUXZlDNTMC2K1ccarD9SirKzJrlZCbIKARwPB63k8xSp4namg/fh0grf+sEM51iuAbMX84
MpkF/0BWHH4lVei1PesBOp/akjK+moSMhTa0i7+aYKf3UQdmjOaRXZzcxfI5GWQIz349A6hW8K2E
V7nKMvUAKM/xCY4R/p227fjuIRPVXUDXheC0ivFsbfG4p4kAYGQCwVnPy1/nn/4NnGpn/XqLy37r
FAxYZJGsz7yJ98enYlU/7/ld/itkI0voT70XCOi51jpNfLiuVtP7zrct7eaxVAaakvf9dZLNGPrs
DZHLzw1+Kl5miXh++OJxESpbs3OPLC3xy27R9YVRug7QM7Tntt78Zz0Cb5b4P9akGPt0Pw/dk6FH
WqzO/1TY5TaP2eNdz83jq1iH8ol932ANeLzE0WOy1z3hJndwc+ntI+BaOH/+3PLjoDNjmzyZlinC
7CgNsnNw6zQDDFjuqPWf5gkiuZxFpTjidvvQ6I5vti/fQmgqaRPbI9ygDFwQe+4gZA7kNtw5t16m
aqZuWRPIs3+xlJ7k8etVIsbPyHuiBpZHNczTYyqvmqZVdVXQlD8h3tmNAaKqYiS9alVZVw/05pWr
3JyabymDHVPB8qA+o3wWvfWHs1SDfOcZIl5mjwx+4g2JoDksJFN+tyF7Q0oMsh0IzQgae6pFw9Mq
VwHY8oTEFfsyTqwvQadYxSPgo4HcXFf115a51EJpK9R8bM/n7bjKhEESxX6JbuHQh43kXTLCTxEq
2ffWWCBUqfqoAFW1WmU4aYNPNZayOZxOE0y7kEcY1LYloc7hpKUALTNBHg1VEspcVcbuqdlsD72o
HsL9e8kmDxvbIYVZOY5SGalqgdtSd8EAjxZVwFNRneduxshzLWnoIcV5oSDcaOD6pGEg/B4Hf8gb
IJixtR/OjYQPt8I4Jd+zNqrcaSNnc630HYZ+mHv0wmbcE3kVlOEa283E+wrenxhoOq80UhFTF1/c
NvTWprKSkFWYzjWPpT6IYEUS6/nu5jXyJ39jctSJrbAW5w+2g8CgHCQX7SMMXG7wokL8Ia/q5l2i
Ibt/l3Uu0bfNh/D6XuLcn+7RKaLWiyC1hea7MFdGgp9TH9UjoLMHd9FogpJP7wFEmZ3kNaXRl5oa
nQ1AJ2AFSb3fVi2KnCy4qoUvTsHkdlNx244jVyEuqvbzewon/o2w5CRVHPPtft4yEVWkSPo6/vXY
4lpWBw18ZZpqxzdpCHu6+1uF1WvQIuskqUtVq/m3tmC66SNB081fb0TjvpY1Ot7c81pCBr53qlNW
43x30Ya8ZSpRQPknsRJXDqrHGaK3oyznJocR2RyVvK3I5WpfNhSVjfUR9UaDlDz5exZ4ZKS08KwY
ju4soIO7xVI4OL8RsCpq6UoFqOKmw4UszFc7r8qphhYanwGyf7WNRRC5WtrpLjbqrvfLNnxhqTAr
VGpXVEmKiHjfivrUnvZLcCVoqR1PhZkD84F++KgCbD63Ovr77eoCyTshEnROrT+4FAmLXysiTw8k
258OtpmTgienz6UmReyB+p8Xzw+C+X0d209vgGPSTvz0ePD8rUqpSg1K5gvL1hFWemwkCm1tbiUc
rFhImkus3n5poVyNhF55aqpPEHMyePDp7+ZTOuor7dDP8BFrQPmD9e8NoaYf5N0wu7u/NkroulNj
P62wUlNCDWgbDqW1Nw/H/+lILzCKbtcu4XGbPL4r9IUt4Pt+b5IB2gtAe8aetnVNZ60Vw2EVRwWl
6TymqlTc1soUqETybcRHPpjjY/UchEBppfrruHYMpjZxLAlnwFmbKiuIzSV6wL1pwl9Q8MOOF+y8
Ox1TnRi7FnrQTRrGvCeK/2OccoDd5PXWvou0NlseKe71Lq2WjUT6avCm/FbFyaPTnW7MCJRWRslY
5vQG8WVkE1T26SueQWaKIjIuUSCTJqDDNkVY4ijmfserx2c4aPBVkwcH6lE2JemmTnRg9dhD6P5I
PGnsNdpEoi8EfxzU3HJByiNFLyULfRPOcIiGuRfsj+zFcogaMK8yHU5kO4ptXCtK+BmY/T9OhVS+
n9wVDt9bx5+V8OTb+QFXb93JMTPUYST6i4zTC0MNDzM9VDfAwmG2pGqvW7TlfwBy19fxi2MA67hz
fU+KQakXrbO7qnLSOLmCEynIYsna9HCZakuk1Ol6Oqpz4xX/KnI0KD5Ogme922QYNcd2BO6hBNs1
GIfQpcDMslQVKnbTdiuAtIQvRZTmOUO/5I7sGVXN6l3OZYxTxivxu4TJk5DeM++jTQvP3/CtLgIJ
hMY4zTbOfQtO8sGTFyBUAwftcQb4d9nYgLDSaAtvBsnE94dBF/B3df+rEaN/CF0lPR5lp+RpQcym
NtkP4nNas1u5geWVl89FJUhqoA1Ok/JqCKuwHra8PT0aNax9AC7pR5zytrKN8+WMzR87hHlS6y7j
W2hmg1FOFIk2FKVnP/Mru3XVvZogW8eYnK0ORudOMA7Wbz4ctgmiMGvGFlw9pj+IocYSif7ZrCG8
e2ZAUlxxeEtlKvpYAkT+B9U8BCyYst4kd9zuzq5ccNALDBJXCfeTfiR8ssHjls07PyBSWRM+6OWX
ARglmYHM7nPqQ+v/YSavPPY82M1Jo9F/+QVCpuCBlt0udS+CR/oCGczFak4ApEaFynW164hTPMxo
XfKTxPvfDCTNPU8iBwYR1kt/+TqAd6XraOAuQa1sGfImFlMe7ZU6kNh5vuwxNkmoMvjg8C9+diNx
IRtsxw4OKYZ/caGV0LvOKar0WNREmXqg3t+B06hWImw92lerOMgOMrZP/W6g+IG9ZyUxOCNjyqKu
DHEWJwBdjDaJZ9jcq4VTpTsXs48FRZbrgH968HYjyuSwHEc0xJOkEqcbw40iM/sATd+Le1QhZrfK
dnXAqxq+HeKtAFyg0M1SVSVKGdVEr5cZwKoLS74ZELHj67DrCgvIRyxZz3E2U88StRoYOd3RGJCb
0l18tJoMulEuFPscGMsJx80I+x/OyGveDFZZsyK48+A4QGIjovBWVklVqNEhElqAfQCLUVFJE1ki
a+t+pm9zVerEjFSn/IbwK70dw7WlDktFc2xdAVV/Jhm1gdfwdE0IHLb+i5C+AVaJD17nT/EvUvLQ
tBIB2TQFxEuyKjATaoedrd9sb4TfTex5rUVko0785imDiJtuIUvzNvc+O+UsLBpnsid3+a7G4hTO
6P5gujGlINrNvX9Vh+viXJJkNt/LtiRJtE5uMdvZyVdDliBYmPL0ckhl3t52fcU0FPd2/OFGO+u9
sgy6T75LYC4K4jw/rYDLiu/ldgqdhZlGvwxNJ0HD4fr35IlPUlddEBzmV5tSh2kE/OLP/Pigw4HE
YPzJ40kLfcxYFoqnyeWg96vGwBxbpy4VpDfN8/WW0QuKY+AwxR3E4N5tNOBgA/kBDY4Q22jqFe1w
nbCkI7EnO2RG7NCXJC6vOdvG46PGztLH7Y4oaugC7mo5txyXipPUieBWCO7ugCSQ105iH4fd6YNm
LCgfpuhGk/ME9GKi60UnzyebiwTyesdFvSGXAZyevtuXhbyj6d994jlux7e0SER39ApEZhJcivDg
fvyzlnbsuagUkOTDjTROG+DCr8q/oOpvET7Kax3VdCGFBCY2WRiKG1TfW9+qLLkhs3sX/IhiAVHX
84DvSgzr1rVnYY79ZhCUIH0tJIMqeiMs0isx2hPbZ1x2HMvapwF5Wy70CzvBwk2K+ibFubEqu6E4
6allJ/8ybkp+VXr5xxJSNoFtVHBWmB9XfyTCUY8HQFvYTP5XVkAKAw55aOTkf1sC6YgznzXydrtR
HTmHvNgRQkRM51QsZj+SSxtFDTRJptDoNktdVJIEnCl2EZ+mfAw1SEXwuKjGzc2dVgPOov5+CP5f
46kHdjOiAe+D0i1Pm23gLa7n4XsJfQPdpq9KV/ANtjd7vMW49tsTSl4+lQYmQbD8pVNc2KrfeOoT
pvSIW3LMwDGFoWuBktUCROZr1jhr6YxK+9QaH+T99EgKlQi7KJ7o1q7JQp9+in0Rr1NO/3TerLyL
ANUUfTyj6dq2fisqyCgwf+8T5SFbCNajRCfaX28ympVpLX9FNeBoLWegizAw1Ob+6BIdr6bOGP5i
BDteE/zqsqdOwGVMQv5ZCbZs7FSE0zUdhisKqMMQwbYT6siSsgBn9dDVCpZ/QsdYDGvfj2iPXAnn
UvAb54tUvZdfQaN4rgHKvaJn8u4KkTbkHMAXW6creGNg7JbQkAkhS+lHcR8gWTO6s8MH6ayT24S7
q0CatjXfn3YUPvhqxaKF6VwumovYTNOBUrMcpOhM7Ys5r7rTO44i/WsSXk9Zd62LuAKkmJd3Eltm
R3gfBPrJnHnABOQd4DmoXvSGLKEVZ/7jx4MKxgbI+AnbvhaR+ecWgNrc4ffvQ2Pjh56rNExYgmrX
BpkgCmCLu1K/rMwGK+FbyajpVA3LEChF6aO0yQOCdNEc2dwYjkeKUw0wxU9nP1XMK9IVAKp56+ds
H/r8wNYiq8sO43KepBB4WbTdoPbgRehhk1oykmqXZ3jOhYyvlbmW9q4y78hc01mI6oaXnAtue+bm
oVapiUcGmeuX6W0prDWndpAfHVc/5UHtjda1PAbKuibIzZTeGRzCxI0IqaD2F6K5AFI3Q/j8Z/6m
ORxk9FALjVxKAuSfdxFiEeeVd4LnXtz8cdBKl/1kGmYSlx9D7IteL/sSovtDGaB8NkVn8+YX8xOS
GL/zSc+PGDeBjcRlO5RUzIbOXelVQASfu6D+33r7zO5bYtzCzGGQJ2ePmrokgjYXa2AOkKRgU1V5
9o3b6oNDtn90dTn+RblAjLFmpQfVpPAHoAiudchkSLZi0+zTEbpAfj1Ta1YaeMcuwFMMGDU0Sb3e
3w5GC+cHafYV8Q3T5rBNYPbmD1v0cMvY7MzdpGSYMczH3ZvIuNUkLcfRGcOyMFmaLTaauWLF13vk
dMD7BMuXbZufzWli6tAXA5hWuoF2zvLv7+c2g7T7aVP6biwh6tjjqrVQTY9z2bQit6gUV+ucrkpm
yVeeU6+jt7JcBZYKrdWljf3eM2ftItcXU5jIak9dUfmrnVP5A0Y/j6p+kGNLrbMT9lbdY36trwi5
gFVvgocHw57vB4CvN97o6nii67QeKxYfU2B4YtEqkX1iA7NPgubqfRPuoqbvdv4bcXRQRpObzfPN
YJaQC8aVpk0iuJJYS39vMUIjnUF8AcQzgO5KE6W3h9rHw/r2QQILTcqNEdnm654e0Oe2nVzlZ752
4WCBvK8vKEUmAmXasDMFGOja0XXwUjY84YEXlHQN6dt7X7cOPe1g2kRNopxB/uz5VAjlMwYjdqJB
q4N9fzBajtof6DoiTVntwyQtZHIctOhk2GlI6S1sYf8iPR5haMQIET1LzUCuVeTkTdMatuKIxRGK
b2kGKZ8rI/EVdEBtlDUbWhRD/GTFQ4FQQdCIZzj+5iUeIFtBd4tr9nRon/xjuVybnVMCDJbDfUtA
TbuEWVsmXrgVkl+U6DPzG2cFDRpTx+R+RK2SM/i0O/tNtKlflazm3xGyBfRzN3yrW49pknKGNrx6
i7LKnigoOWE6gDzJCJnjwLZfWFnJdilT8XPMjx9QSQ27+BdjRd5Mhd3JkgIubMzbR59r5WIItUaP
MKjf3nxQT5nIDY1JQM0VrSaD/30cF11ptRkt25AOzLD6mHJHQSaEkksacNHBr3lTf33davZsHSOT
Zp/l0GEoYX0DmATM5OrxYqfFDFPQjcKYSYXAKYhj/vc58pd6hKdlXSfxV6kTG1R8BNw5HsLm/UWZ
ZzVaHSZS1y98Sj4RYnEQEIFTNF/wbOy+tUVIV3DIOvuwpx4GFGob34+3rOZN9RU7vGL5V+S1pOki
8UOCbdaKw40pzD9p3hxW+vZzrWFIgeLEOsN6ARs/vQQnlcqZ3Us+Ns6KhdddSfhtGPULCS02HArC
PE0M6MmW7ExrT5JjD1fY025YPfZgI3RVZs0YzmFG5lKlR7XOCP5LM+ZZvmLHdPxvlRHWtTayr/f2
+PlWLVJsu/WvgrMPe3ALrZGyQfKwpIOw5OFOFI11HNCCqTHCpeB5ilTiid/TgxIluw/Vh/i2vBWs
2CZGKHwdyQ4qEfagWu68M569MJeNADnBVxIAnixe2u+BHo70WIm2mDMPb46ZKGFo1lw0iZo3eAUe
w+yNkTeSsJ8OzYioQ8PU5Rjxjv2zHtJl/OzKg0noZ6rJXSMFrHKlcgyqunTXZmOdt6tXUgJuzb61
EFFV3tExmy8tlAk777/lAfT9+m3sH2jd7/4Ha4ksR3EDIxzQP9wcuHcuYlqm1sD5dZGoQbPH2OPc
b2ffq1OsMM+fTdoPYdWtJmG1Z8roTywUtihi37x9VBV8tzYJEN6DsxyBjweZ0oCr+c98ZPAeE/2j
gFFKeMYy/fFJ9Fb7KgX52R++Pwe6HJN4p8lRE04jN2G/CgNHUQlo7/QPtCTFyR8qkABPVR4I3GVR
Obih0QJbGhfG+WEu3x7fGRCO+vsejIcd2e1J0SuiC3TOEL/0p9m065w6M4jw1J2VWvmpUQnIeael
qaJfREEPZPHAkyBWyRxZzv5XE7vtxtHIqDxHMmLIArUJhmcZy7ZUI3alSNV9qeFK6nSx5v1Qhm3d
jNcmr2SozsRTbO8ec+ORzPZS8198BpBEl6H00eicyWyOLiVXMuefA60BM6KClPKwqAqdcqT6P552
hIaeKRietC50V37asce21gZxxnOVHb6e76fVWYBm72/E9safQWVHqY6+8XSG52JuZl6OyRwqQ911
sBvUmCG3+FjJVhazzTvms0pLVQJDFEwY63DqElqTdvBaA9l+0/YhjnSeieEFp5Ma00OupOzPDvQg
P/mmA7aIM1yOiMoCOGSHttSfrr5I5G7yPuejYx71HeExVDuYMF8lAe26Hw82jevw4AvHWvqCzClw
1emXUwQZmau11kwgn2K93QeKAV3U6FETNazdxO5IKf+GD9WqVeNjRoD8PWEA+vjqxfxB6Ex/v6Qy
34a/m+oo0u0sGxjXJErhin7rDJMAXWpoWbE5qHQtqxTdGwco1pVn6FBNMPs7AtkXrmQzfmVZW2+L
d3zUzq7dKv6xeUxjVzARQoI29c14is7EkhrnKv1gEEdYpKq8qsTV2aT3ena+02X0MB+n5elnYWqI
+7tce6dOcd0vcRMiecHlf1HNywLs1uZYwi+DadwqmB2LYqDC3TA6U3adrT/OU6Nme3rRMC9LknGc
QjsBsZoGpZcmiekyYyyDTgSnmKmvf6SlsmudIhtO+iqDlMLFeXksW1qzCUnwwCCZ/G87+hSigcJD
zF2+EJp7U7ZRT/VUbdSLvRHxzEUnFmJpsZXGpJeUHMaflcFM34pTDlXxs/K25NkHqP0dGvvgygzA
H/ih1B0Frix++13V6kBu2P5IELGJube4p7D+L1r0CTwB6Y77gGUhfbGnWVMD9fTHk4gOqH+Ai2Ki
E0xfEpy3ccTI8qfpQxHzARWeM0njpzQtY3yfNxONYBkpvi33nhSbcalkRn3uP1YY4mSiG58m3VKC
PXtbArynXU/BEkNwtpWIO3x3PRIS8iBUvEcZGLUe6EKgH6stI9AHzf8+oWrj/fOkPqjOGENDvOL7
bY/4P2I0pTrMBuewbpUAvYqc3QWEyM5f/dmdQiwFZLKl/ELlB76e9xVhw3GARO5hdtmIfiS9jCoj
kc20tEjZbOZctJNCujuymq8xi3yKIZ/7wJmUN0SRBZ4+w2kAvLll9VBuIgJtTMKitca1B1/eVlrL
KXiaLBjoPcO994geNvVKLbX0S0wZaWZn4hpCWYk78AZZFSYaP4/p0earSi1HBEM7l8d0TappJLei
94zXiFRJNp+7V2Kj/6twegyQzAd2uWhxQgf/0aqiw/MNvQJZMHRttbyyoHGUXTOkiTjQiCC+taeA
KW5X8aIuMOnIm/rIiJXAoEXoWbrA/9J9KFriJ9AvtGCmpa2cJWhkNU4JzOXDDDIOsEAAfyj50Kkd
BZilnzUTOdcZSIhhlXattPG+uwDuh+NRDDIOBhL5aj/iCtDFc4htdL9yyExSPDslWxIlG5g0GMq/
i3CxppGoLUSGS57zW6LPNUefkZMb0zFTrlTACXs3XXAX47UuTOzkdjwEzxDX1lY+8psc5Amg4uKm
YB29CTC/++2V2r6cT5PtJ7uYK+7jiLqcRo2NClYd91ruBeEELdPVUAx9CeTcCFEW5KyaP4rcSER1
T43oLfwcYILXzf6/rJ2VmVOC9lWUBKbOcmopccpnJTRLvEWp+qGf0N17tz/rbr9RZXr/pgzu1Ba2
zGRAa/+q7iCR0hd4OkkitamqkHzQht/NMR1AVAYdi8AOL3Kyllgu30nDTLr0N2Xxk6flV2A64Edt
LXLfBhWq+bmjj0evoDsff6kF9MN0oNfBQI9YKEGe0WGl4kDG/ytLbjD7VzFfFMurkEDdF/bWjs6Y
510egwYXPaWtC5YBsJgz08Gb+ihcPe6VLFkW4Gru/i1Y0j7pcoW8wpYr/exJ2nIDEARG0/rgZ4RH
2HTkBmAaBUcLdy7d3G15/HaHppszBwTjRd9f+gatfTxwqwJpx2SM8b8SJqH8qwGoOoLUdHTb35Bu
+sV7/FBHZEUTn0ebSOBrfZsb3/o/H7BT1XcfivdvBUW5FYaSh+aZu4Wl86V1qba3Vkd+LU6Je93d
V1I72fK1xKbLd7Sw2ofL54JPIFKshN9p6SPqwXGivWe9J5WKc4Yjfm9F+E0aB21Q9ulbgtfqzIoq
N+0fWmBPIGelQYLLqqpF0DQi4WjcgY6ZXLQQzMXqH8CN/5FStACJBRgSJcsrw06cZeMSBudJq6H1
0GS6ss5tSgyJh6mf9e1dI23EGn7deSJHqxC3jVcenS5F4SwFiNOYTDFGEBiK5Mu2xjWSwYwcWYgR
2PgLSSkFV0s0iYhZ+fZtgacexzTSeGDpHeAXl/GiUkY3kYShlkjIrmQBCLnWAIqUGK1dtywX7u+Q
ZuqYV8SfBeTo+uoMcnytrNqz1M01VYsLqs9TMgbVD593QhY7gFt9l1M9TcLXI4S+YXBHPjHMvBqQ
PEGnA4fJDTBLlFWj3uJl484FlqNFR29HozK30SXdLalCoS+hXeC95Qzk1IXf5YGRZhe1tPUUIvpK
thz2Oop5VAZJ/sUkY1hWVDalipCy2H64rB9hFDKn0lgMTKECAr1Ko8te/SoYZaf3DdxjlQ8c+4V0
7gNQB36hO7MQaNWIuTr6kGNe75W4KmGQ4XOh772PMov/vxeJbusvgITbXxNzkXQu6aPSWM96klI2
9gTL8GkEZ/TtGI9FKrTgedvksnt54Kfori20o8gE0iO7237Hdka/9sjpqHlnuLPQhLufitKbY63Q
tydc5XxIVx1w/BnWCEX1XVjv8/nRny77E5OykB89P+il8kQ16AFTwNDX6PZg7d3V5x9HFKNLyzuM
gb8xVM3zW8MOojw+zFiI7cAkQUzFvGZE3YJMN6JI0Ai8vpcH78PjspZtXmjyEXjRC6uIY38J/9n2
B+6RehJ+nWIoQwsp98PUOZvk5pReXpg0Yj6k762i0a2DCJJgqTBRiYh2r3+VCGiB79vAiY9W148x
czM3Y7d995ciZlRdyHwPCedC2kJDSRXCLXEWE7+Gj3p2VE+sq7sLA/5E2H0Khda2NHpOqgWCIizr
zr98hkdrrG6/WovvPUpJV+Ymbs63PV2Qvk/IsSxZuPgQRo/D7awb2GAhgEHAAPg0zYj4z6ipEVzg
F9ZMZM/nivQFt7q9k1VEcwE6+HSw+yq7JUTYP22JIYn0v9nBxJzLK06FHAS8h1PiaXYakfVfiFRs
FMWUmV07lu+/Hnq3ixPoM4/4VU2K9gDyPm2D6WibBVAOGwMxCwEgCXeCi8FrqTFdwahu+qFSH26H
QN3Chh6n63a4zWRrpxcuQD0sz40GhNDZIYsMt1LKcQTqhQMhp2ybKRDCdhD+Qm7IV0iFFYHY+Bfy
X24ICwkQUcTt5AbAzgicusIPnMXm9X58MgSsEo3Ehm7dkpO54jIY009EU9aLUnwfANcyLquAzaYF
8d+Wzc8IMIesjtre52ejPlHW14XwuWH7/rFPXWbDZ2d9Q6q2qakvaxGOAqNqLpraNU+0V59KHRji
tKPCRRRWg2tVSmoPWVviLj1MpM/iLYgSNNgNAHKKpiusiWMZGv7CbPFVLnoVw/Aj/aBLZrvzXUH1
TIUuXwBeREesHSfSYQRYjF4YCkCLz+kRRxK5gZYwEHpHLXZnRw4EYTgHXdEBuSGv6qpgydYb6U4q
85TB6Iop2IVPLQpI/wtHiCOYohR7Xn9f2qBWbYPTFxDVaZP9BOVL/Vb+G4LS37PADi5JHQ44YO84
eDw9SOYY5d0RyXqzN2opyCOYl3Ts2HlYloBX+o1k4Sod83V4ultbiva+INFCSSP5oiyDYA3jZX3o
1W9eMsK9v+ZdFFVSkkrLs6RZE80PzllhDt49vym8xvDJBVQz/yYdkSLaNqUBxBp78fa1kTS2+8CL
onoKdp41LyCIR+LBx34uB9rCi0M3k6+tEfaI4xM5/yZokJpwgmTJM7tDiGzFt5Esiv0cRvFsPMEe
c2VF+hc65AHfqZF/TuXklA8aOUNMHTwjIe9qO3ekWnLhbuNsfokE1EK5b/zJJR7hb4gIj7+UoetR
XenYLw0aWnP2x6+rkgZFg8xL6vmkK5KrOip6LaXR9JeRBj7XPHtN0yfzCwSsOT1S81bGkDvVzUDp
m5PgSObKc9dbIuvGLOK6ekDTV5LgANEgDR1VbnMthoVPCcWFBAXVDH5qQd27IBNGhZcH0CDOi5xH
mlXrY8F8keQQDJH+HE4wl35OIDVWBrQa1YKWyQFEiDEy8KkTS0UxoxY76bWzPNVYKfv6wLZCLCIb
0T7vh8AMDz+8y+wfOGeyRMM/ZzBnzuebr8TBZeD3xOA8071paq4fg+KeSgxRBQ8rEOBpuMBgZ1wP
XrGErn7ULMe0u+iU3vxIAn5LRVhvUNcoeRGlepakVTyyZe4p9ifK0FswYiCAmiMU935bEor3NjMd
ZbRcCTkcNygjFOK4oJ4Q26j203JHsSkRHNoTnL3wfkDXI0LGTx8GkUlhXq77bED+2tkR791cC8hs
5ZWvXkx1yTZmij0dViEOJfLiXcvNorkvR6agMQHIv7wBCJFejbrEITGfYXYAhDUNhvSvLpptquui
1ZRZkYqZnAktnplML3hWkOsK6I/FVnRwAHf22yyEaJZ9lX+GweIBdhzDonz7jiunHELyEWB6J8yv
HBwnMZRK+Bupo+pyGd+DhpoDsKic18ROsugJqN/yxbHcHxDd/yC1qXGnzgFpqvKDwjghN0koJ1zA
gf4uFngoNNBDQbxmD75gsASebDopUa6xIFbIPqnC1/rMbYPLloDEuTGb9y8knn8swcQFo5GEd4Sp
G+9cJU8UX0xn98amiOboSUs9XMkQCpuqtQURV3h6N3kxQy4rt35UWEgQZ3U3aUcJt4JEJ6o5z/9V
loY7FZd3snqNqHvsU80rm3MDvH+tGE0tWrNu/H2ijRjfOTXJHFoBRcqXzOKyXFVAKcMgNFV/qQ90
vLSoEv/8ooipKirAwcce02Lq7OOQN/baUdbTocKFGgfyJO/tFB8I7q56u1MM+eiV7Y6eLDLWhFiR
9b6UOz480d4Kz7zcOxonT+szLUATKzyxp8Vdo5AeR3RvchdlMqAIC9fI52TaMk+3TT0IndSk0iFE
Ui9++EdW58m95pBmh7OtCxlOhr/SBjpggrFpinkaW08KcunwhTxqR0Pujr4pUXcuF+EXTJhwiWfx
4ecxsSgqHNMlPvY2zTzsaa22eduO7NHF/nKS7LvHtB/cK2oKqI9NiGZw9+4ET0wkzI0OVYczuoMy
7XdzJjzwfO4cxuQLoziTU3/vENuwr/4/To67dn2A7qXzDwFd74u4YXdPm1hqT63b2gqF8+JyFn5W
GSNvjysVNiSWgy0u5tUHFIHoygLNCO+HjKtUW7c4ZGedot1+WmVISWOvM0a1j1A9VaOh+wHqTZXl
7DtxaRz55FCYQNvlz3iVI309BCJ7WfVvYvqTezsFLuYngGatzD1n4/g9sPbN+szAamz9WokgKu4G
l7pTGR/ZAy8aml4fgRZTpcQHSvdgTSLJRfrsaPTMb1PtMSufOcCUPsXH+Fzwh0jEyTvuxnBtDncl
pix4EOrzrL243ZnThKBu341GOXhu6eOrhzK9Hs1Tmgq1jCsagobHFrXWGkq53/utv3U33mlGnrYK
tiv5APM9f3bx2Q8LHB2l6OFscUS1DCC6b7ARl1qTMkwCEgm7EyKww6MY7I7uxFxLOvrQzubxaCC0
DNSH/KuxD4aTcJpAlsHWU/SHxltEONX2kKZrbnGX4PcXecTuMmzAFgo/tNtbf3wJvMHCMwPEyg2L
Ekq01gzS3Y00yqBvAKAQfqO1QNmG5vK/D2XF604b8L3aCrSUX88W+Mv4Hq6GAx+RgHexJPRSkJNc
elwmJ1kAId3e48zBbWbXlnlSW9CfY+0C8K0UI1bGooAwm6IGeQSLtV9pHZx+4L0zYvIwc+xyMoe8
0H5Nmio3kK4WrP8G1rJupMuH7zPrj0C3Om0k0vJKfXqHvJJO60R+sBhxp1zrD0WOeZfpDydly1zn
00KGX8218tSaMxyJCkfc/myb4deDhRAVCIKKDYQfXDihXQsT9hIsNlxQEXsXeYLWnnFzKJWtaxLj
WOtF3dqNwV+VDjFC2b2YJPQMonkpdl0ubDOp9QG2K/U0uhiTx6dnq6ghLXK6VrcMhOkk1bWpv7ip
T0MDOOzVDvLp+7XqE2xiacYQ//BhsReYebS0XCc3PEUC4j2jd4wXGw9eLV7PHFvyIDVgBKYo0IQb
m18IxJATo/YZwNaW7WV2DYxx7UZsM2MOVA+mTLuPC7Q10v4ByAWL83Agcx7l2jT9LoCrQHmbXkAA
jdn1nlIPJvKf9rKp2ELWLI5FfydTEFFt8WmAZ8j3GERQ2By6z2/NGXM9RTvWyNqIE93Fr5ncEw==
`protect end_protected
