`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
cvytd1gcLOv16HshKQiqVCShB/35NuAOImJqqpECS4P8vof2idrYbxa+Nr/dYBCjLV2mDM2bb8v/
I8DfdKEJ0d4IxrUJGw4NJ4803Q+VGAAkHfLiZvPDNScunpWV7ND1vdtTal990wEhFyB4PMyHQOir
5v6lK0zWpanauVYxD4tdWZOzvGrvagOTN5zrtuKdw2XX+g1GJe6P7APO2jWbEOicDMqhnIYVcyP5
QZPr7s9NfqJIxZL8Yt5ZqbSy226fCrMxan3vw9G4Hxv/BuS/Vhak0Wyx2TYbzPyOpeGUXjJaEcBI
g1HJVVlhjpgP1NMSfLX8v1usLyXqKQZHUjvGMw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="64GJQcUNnQZXrys3MbaLd6MaHSdccL8iNc866EyUIo0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37216)
`protect data_block
sPdqLmKOxwf/ezdEeDVCPbjQWdsUcOcO2ArXZPpoyEuqQrNww+h5vhRaU5TImMx6cbotBwdPc7Zq
ByZL7Ud47jyRGYd9KwW31RVKX7KVzm7FYI6v80xeB2AHUv6Xsro5h//mHoQdoRihUHbtc0oBm4qN
XFxorMfCuowGITmQM3S8nAqHVgOaY4Al5sr9TAcFGBjTHXmBnD/zR8GFBdbRpPqyJIVRN4prblVl
tyR8RHKKmpFn/3Ux9Drk8JN+wlU6aFKPual5UHY6wx1n2gxI6dE/nYvCWr/1/5Xfa6h8mZnROnKE
9zeyomJLmdjlhQIXwAwvpiHjB9s/BSiXzbkidJQU2ynMcPtZf5mDOeL+twhuHhIdXfNME2DtJDFo
1JP/T2AEczK8Q7uLVx5MoBoAIp+Kp+NpyoIQU8vYww41s8NxWtPa+RXy4NiE5pSUiVqZvNSMfEYd
Du1VB+Bsg/gpBdGaXoMAKzq+PeA7Hwh6pLZF15wvSoz+HvcbVNHLXqQKt3GrMik0TQ5GOyvNqVuz
L5FUe67d9C6hsJyUwGmBgZ1+rC2Kp8Nvz7LULHK39XHdfPnkFLGBRTUJSQRBG1S9b7dzVUZPsGS5
eZ3aRMoUlgYRTSkASRONMSLFA8VlZ0r8T5cRYTv3uPr/niWN8YIzgGbA6FTplY0bvK4oEqHM6jTj
4roiItwFGQcWQtXYwBfXjLxgfbMsIxlg42om1tpNR1wMGZYiga2dnOhsCMDiPOpdV4BEkts/bJd9
HLeGMzbK5o90QjQQ0Prn3lswuFbN4CKsrwjGOXwgJRhBanJg9CARlsqs+4mvWaQpp73vuboS5VIH
ggpGW70PtTw7oam9Xzb+ZnC0tzQt5EWIrwNDmpTOlnP4Lt3G4ZCZDptX8CLqADRTWTgYXLdzSpqM
DYDUK3i80zXUWSz2XBusamjj1znhAk/+gV/jg4+gasjc05k9o4h5JTRz92QxHThjj+wLTtmwMYB3
IUjkS0IO5iJXhEEPOqwiPWORNw+OK/tEUMBSh2ITzMyRJwsrwyhKgVtosGLwKE715EqB9b8LzIGe
rBO09/qQvmPoDVxPorXa8Gm2eHRIywXqXfuZBcOZcM9KghxEZTpsFeYCY+T11TkObDQZ0rTAuY6y
V8JkVlttowR+rxVsT9cQ3bhaqA7Omeuq8rLXnxD//KopNfXv7uten2OFwvUukmh9iPaS9g3L15Yi
yizsv1rzkELsOvFxFquB7ICxHv3i74P6HoUHwWAmnEtLgzfaf8UXTJO9i8l011lInuOhDVRCihXH
CyTHUB8bocXJTKvvJH3tMYrenXgbyMOW9xOxxiqaSTJyV4qcdPf2qm7/eT0t8Gw3FX0Q7pi1cJfL
F439VcWkdZPiQvlUPrj7/odSH8Rfvm+cf82QjEf+Nl8lRqaL1R5kq/pE+2QKZIcyUMPYsrYRokRz
T74WwOGjgW1M1owFnSvy4K6VVCrb4zObnDFG7n33316v0U4tbMOTyxLSsE0fez2uDYhbhUOe+ekY
UD1XNqLAUvWYYJBh5I6K+YiZ/zovn35aD22JgyxSUbiGPWBSqN/TOnAJivTqQ8hOaDmHqOdwyNt1
OYnBOfd8p+a+pG870ZxNykJK6NREQoez0d1U6Qino2R+Ww6iYyY+ro/d16Gn89ulcIQjczrmJqMk
5zOg9AEpAnDaR6JT4dwTX8Kik3eGjJLTETyc4IEBMeLMTapWIr6sx2BzTyztOqHcyk6MnnN9hCHT
J/8WL2XIgKruZnw7mIMmBqlpoQEwPqvERQLhpTBy/NmxU/oKo9OIGVUcZaEkElTZl7w2Q7NTRgVm
zDakPPndcbhnFIvt2AXorfrDCGisRVj9y6lpGF0WH2eBD71LktCBRZddnM8nyhXxGx+9vv9mhM2d
AVUnwx0uxqk+a4oIVBhPwfKAYVsuh8PuJTk0JQK/Onk9h37A2CAKXrkdxc20rC5vC1sHuPWVUvvG
2NXFJ74dlEaYNkfr7IhsLJ/kxiGWtI1VG/GgmS8GxIAjGpcNOy727J1Xu2F/Mf+HUs4GauAn0AA+
pPqjaAI2O4KB96lhXPnotKwttCdnsebv13MuvJ9fojdjGoD1MgO4stQskGgy8C4nMGgQBL/7Z89t
y2IaEIqtYfk54ggG6EF4cWymgcyogHCpXlyNBCWZ0Pdxf5//lPY1a3t1Jg7AiGImmF8eNuzgwj/D
GpCew840i5NYcRHVtQ4AjsUn9E+jzynZ69H6Ac/Z3hJTQoxQ47ZYxS6iZzQz5mdQu8cG+dVUv5X2
6HbV8vWOXh9blRDeFstCbLpGGLUWJbFvMPEpjg+QIQXzc1KqHE/c2+X/kne1j/PmsHM9TaR5s7/X
eObtvy9/MbNy0BkUYMVHu2qGWqEaCPbiruSOH5C9DdAEwN1nU2WsNyCp0UfgNSBNkhliQ/fFN9Li
o17V5QJnocru2Nz1/dCc3z0ccDRVEAkZFYz3ja5xmOhKzoMSX3e7EPkzOBB1nyrSXSo1rV5xxMIr
GJvj0Nora7KlUA/PZ6bFe/Bb65t/acKeJ9T0EEYcShTvqrMwrmmuGROrjNtN+kDguYJPiRNG6H/T
xU7JLvYKUWg7K/SeCzJA+xoN7ZGw25CQ3wg5tl13PRgxJL01Dhj9khm9m4kSZmYI0VoqsUiRErzX
7HriGWDJyUYIwf+WU0LRbuKFLRTwdhoNN4Uh8RLGOH0FhyNJtcQhcy+3etJ8OZwyxyzbHwToodeR
exX84PWiP22p17D3B7y3NLPHjkrQf6B+ZhYnTX3KxttRIjBoiMbBmUY8cLQ0w8x2OWt33Vag3bAR
C9xmBe3q4g97nSHQG3+4qGrIiJItQJSis77h9vOKhNrNENNLIJsbbkxSUvbESelFEYhMUHLN9Fi5
7b5twfafoyKLozSFF6Hp7VLrpn4HNHBBzJ1pEqyT3GvEABkC3hycFLIt/Fp+fJH+VIDpiCIatwfV
Y2fKKxZVWEcKAuUJbvR9JQY29flUrRe/p7QRl2CWwt+LS2MORQJgVVoAvYvKiQ/2KoJk7okDJVq6
oRUwcdpwkzUK8rHbYiD9RsYPEABf8nZEv3DYrzXI13z1j2bwSAd0VrWkXVdJXm/Xk6H3ecAVQddv
twUfIx6xHBAcGwaaSistSZKIY+o4l2XssNd7+VFQZ1NQ+Twxq9fUcDhxfbG/wxovLwXdHLkkNg5J
qIrI9fH+b1X+9DRSG6IX4BH/TOwh5HN5dhg30EoRk6XCdFx8+9OmXPp7a9AlZz4q1ZpPIAupYTxp
2JoJcbgJQJ67YtZ3+p/NcVDfAqsCHECjhuEBJrZvGyp7xHa7tupq5aK3JtZUtD+gSBAcCj70g14O
BANmqtEjrpa/frktjCK+ZfrsQz3+8UlCytyz2cE3Njhh6tAyDKiYh7kMT+DtV+bzaWEm0M1hN12I
/w3gxjIrciBi6zMAJPDQVCJJH/lRl3Wy7vyImoFzz9OJUmWjvzBpBi0DP+mqUOphOYQoFZLyXwDY
ZVFirY8CVoIltIQ/5vTSqv3+tLsssmdqkDqsCFt+kgUO2aQQ25nwBl40+iZwop+raVhKRo0jgkKp
6ZtQzn8tJlLSTUZFXA11h62czLj0Y0RV7PXcpKcgd67VM8Qb6TeBxkLhXjQWkXDHfk8UXVCZvuRv
LPhvk4UA8IVJu2pfKkxA7qdMt0ondTIR5o6lS6fz5rAHfgjXyW60OKgfVYovMdILuhbjxJC/X8Qc
Qpu0D+tLm76yN2MFTwbA8hd3RDaIVClIAJ2gdn5aE8AsojllYblIso2/8mN76EAD608FvnMJ80vK
b5KqREnc9AAUuh2dhj4v6sEnP6Qvpx66rJrOa3gxBWzd6Eb6FGO05QR3yrNmjVR2iEUv6TJwKRg1
G+D4MeETmVMSw36nh+QklBL2FCvdoa8WuUji41wMpsL/4oQBaa8nlJEV9KNSDN8foEydhKbp3xNb
JfsVCuVo4Zax3SxPcbwhMSeG4y8aXf8zKMEKOZ9nmzFxuAzAdMuwal3aPcNblUJ6QUlhQXc2r+5X
uzS1ElSX4qMhX243TF6/uEC0ZqpgODH6aNb4tAq+IUqiWPcY5Cmc35jTVk+90rrXTABzIhamSxy4
FvomHqMvU6ebkVrm0OWhcdCePKDcsRSJ20VsrJRxvfsx0U2f5r297TNDELgvmSFZuc2I2RKBTjHO
HgP0mofga6c35Ws6ROl8VsUprr8a6E4bbZORZyHfp3vp+GGSAIMKdeilIvl0yBBaBpHZ7jbVcc0Y
IRLU1taYosj1hDWdVXBuax86Ldaxc8BhK89q73SuXl/hIz1s/QuNbttOVfhSTiAG6l84PivfwgT+
Vj0N1BYH6PrTKfA/h7KhE0AV8PJvgnIasGAKEgslX74PkZ2JD6pxfM4V5dC9CWkyT2XHCZBi2EZs
BmumwfJz7glPGTdytJJsDxR1aJRKTQNWOJ6PIsWg6Y2cYh0llj+GZHmBFzp3tqWTf79WA3IlbLjt
sAH/Y3OL9EVv4Dw741Kp/vFzW+rTqp3YThu0h9ME5S4Zl2ALRbXqYeCyMu9Rd4ZzHmMszFCX9Cse
lm8tClr/Ez+PJ2bHubHlpPX6s3YY5DDVWGT72asJDE4TOWVhR28UahmNJ7eANt9Fj2FtJCFSKpc0
U8wcTmrwS7FWFhvgR66XQHPKksgu88igmYdQaYLdyfUvRsjLX2BjmAB4Mcv8s7NBhfpv7k6oPWvw
hW0IVPup6TmZKNQotpve/bmagPZfuSey1KXVChU74//k7GA42FP7e78vNGVC5EEA7knHqMZRDF9t
g+91y4fYHToeLwt7iv6Y7722/sLybgJUY647o+tREHPSqYpiiJMxuzq7ZfrUnUAtDBxqULjfjs9z
d1ALTNTP92owghZU1EgiMk0Sr0BjtFp4liH5f2sGvDfrLxWGJqT8OCDw2bL8KIleHyHiF2pqGGxD
/119BRJPAqC1wzgIYAPzMtFpADQVpVtF1bQciX6pxAf7pSps/cSpUV9aPmflX7hoLhIxR/5qmnI/
xLujN7XSJ9W6OY797xfd6tyODyJaFfBuneXR+ENWkiX3qvrVXGcQZuycuerKXFaE3xQM04YBKGNh
N5BepiR6z7OWbI1tNYo9FLr7bd8RNVZLBi6qpGl5dfiCT2Cu6ryt1ISoaIZ6SxXGKGQufRHT2gG7
3p8+D4Lvkb9BLJsNN5SH9/w1VzsIr4Ue5jT7fD9y2/XorEruoimR1tScb9KJLCEO/5uQi24EVbPW
kJ+qrWCYA6Zz/PpSIDJ35Cd7sdy074V3GMYK4PaJxSj+a+6FAvyP/yhOvM2OlFD4maA/RFxhGHVu
zU16tVUK1/ii3p1JmeKuZQ+vi0sKTvWEHm30Rb/sXWfK1Pys03UwUOPLc+9aw1u1q8uzk2theUh2
hT8m73c9kIQPPh4PGtJa+rqEC89nYbmOApiLfrvlqIpv+ay/K/9N8jvqy2eTIQBcimCw2/xVjqm1
dhYSjdzY21iLws2P4ZdZ1u0wkontMoFKNxfbbbjOVNbxogSUdTKgoAqAmxZo+iynFmim0CEFTlu6
BmQS4OZsUEAQqO5/OFZfpNh1EYFjGe0jUGSN/VxihZ8i8JLgyboCUXI4uQZKAjCRqVHh9UdxCQWC
7Arw878fHOwa+q4wUIrulr2cq9bk0qLkUdIHCpKMgbtoHkayARmbDbbPpatmHCIzValZvazXnwSJ
eYHe3PqWLBIFCbHazKibNwcpw/X9aIogY61t2vDysiLGmXvEWNDWYGYuzQQnPCDMAL0oh453wzwV
4ky2sYn/6Dj0BN1Pggx0u4G2ApoX+G3iEpi4Y2rP+ZYsBd65V3LwSOVVD9b/DvXEa90CxZchf1AN
TzjrjbJH1+/Z0LMYkEZAt1+tZ9JqLRL3Jq4yJKeiYfPuydXrVfKdgqEY7moUFwoxtESpaN/ODD+O
yPvn6DpncuKTiESoqjvlkB9NgA/SfUjlfR65lRMT4iMc6w34KTqLc0yoXuKSBbna2DL/2uZAtVjU
Rwz3T2Eprx4xacjYScaOJRypdYZAwqE//7I2xJ27rZuM1h+hStH1KFsIe/vVOPqzQlj7CiBDxIvX
99hd6E1arp1h7i66qaslOAx4QJ73CIPNCQ+fQWzaPujt89oLz2I2Q1XEufjru7EMihjqV4XTMIB3
jAnTFqH7Nx862gwyOlR2C0C2/ASUhOhjvNEzxylgb+2s4dTV275c4c9DO0XlYiGoCTFj56JUZOaQ
mJ85z/vk7vNhEhSeS+2elhvYLvrsZrp34alZrwwgxHMFu022PUW3qXHJRUJrSr4PWTd6yKzxr0d5
p36ZOhj9CnweWOMbe1UgDB/nU9CGVMzbL2ZKTYQowZc1dzM0KWcKy9Zp6fKAAC7E93srhX17Dl2Y
2BXfxMd0xW5sfoUvu83TjzFwcONIv8uRqspvuwbgdHGe/f4ELsFJNk/eXop7/WXDRzo3r32vwF17
K9/en1P7HcvyI/ox4kI7nqcuFKMnvIVDeg9OrcVRmlf09PowZPM+884HrY0FbJM6KI7UITamC8BQ
pQwq1HtkZaKAWW8XxymrpXKjhyO9aybgibFCmpql0ZnVq9R+6XO4pZgr81a34v+C1Cij6FLqtHmU
CobM+l8IjLuqRpZnHMN2izfP3xevkZVFFmDwdJSK2XyWS5E0CYszzTkrVX6+DwOgSdPINZDutP+7
/ivrM7dw03hu+2ZdPLBGbVYMGCdhBGMug0Bdh96iXi0N5jZKRzB/68hik0UvYp696vmu6ECsgrl2
Zv6/TMF85wgrB2RY+ZEqn6mkFwiExnwEEzwd0pTvB0IvByofLVP2mhOuP63T1cp9y7nj+JSyMCq+
cYfZpYSxh13KJo+e8jx+ztD3LSlYSOpyDs19XsfyzGDHxNx05unEiM/MEHfIZItiVhPPVkLItlKm
zuDkdW7AXFp8QAtu9i9pon0X+buObHDnOkrr1x7/gUmF9Bxm8tbtx29pkGY90/8uDMogLHH1OQ89
06KOd8E0bQYFH5/JH6kkdkFfCktXIYFC6IryD7dq9qto5yjbF8V+3274d96RgpV4IhzjAUXqwalg
cXZTI7t4hqxiH3UEHNKM6TPUbp11YRPCI6ioY8ailqyjskpUXg040DuFLD/J5anXwMySDyVgq4eo
oJbPxU1YvRxT8BB0bKsuhI/cvDjq+5UVmB03S7jIPcG6jS34i06mPGAAoX8MIF5U35WTgvZo/iN5
6OknN5OqSOK9/PTEVmyPgSuBvBCzYlzrUYp0Onh/XDeZxeydC1Wr/yFuQXKRZjNxV5YMizfI3Xhp
/nzdNtoQVEfBu500khjAgCL7kg1bAtlk+3jMnfGIPhbA9iD8jbow85RHxN/OfqOzgrDU3Ap3dP/J
+nIozlWaHpWj8OwBOJVyF2yVMSv5TLjHfZRH9/ohlRc8/TRU6ZIfLw2jKc3k+W8b3240XyV8cnjT
f21GMZ06Q2FdEww6INUOseNm4CeGDOXvBfGeIMK3Z6ukdoIkKLgAnJgEokPv7Jg+zH3MLELAufP4
SteCUG8/hU9ULj2AX8Hyhov2YquUruAkuqb5RTTKU3NA2ty72Q7TE+hQxRpfbP3BicNWLv0SfUaW
FJ0hv8k3Xrn21XEPbBcSwmePcUpM9S2dRW1z73cGYdgztrwtwAtFyUw46Muek3B9g33sxAkJnoPf
bSjm3eB+z3UJ+BHYo9e9yd+gMX8KOXa82/KWvgzfdDshjnO2zlEuJdDFfdCGVJilfuyTx9NtO6CE
QT51IZzkgDW17Hnq7XWicuB+MwKIl9aYf1y//aeRX6ItqL6SlXXR33aQiGZJUzBrs6lbJ+6OT2CS
AkG6/QhTirHLmm41p9uY2heWP7W6VOGhYMldOU0uxYiOtBwqbF/Yr63p4E+eR08f/GP2LzQWs+tE
CHv/fZtryPtxmc1TaLpS4ihTnMSKNQSrbrDGw/SdcAMfjQBV1WerI6mR3fEn/qIfRxFRjnWnueuk
AaV1uGHRCT+yBuu0mSXfnzmuZJQpMR7uVLcwD0N7Aw7ZJEwd7zkgbgxdq+b6owENS3MU92yuMSMm
I4qNll/NUWPsz0KcR1DZ6Xn7yBxtnJjjIgntcirH7FS2Y2HcvZNV5mSzANSlXVnPODiKiNlZQV6Z
FP+768kpOosZaobDYF1qsORwk7PyXHTco0AJI8pQdu6C/eWfmXrlDpweTSlg5/jvwnYeJhEIVa5B
MUc1KrCRY3KyMwvT8fB6gvDXRoh0nRnIUx5WtdV45q4kSgPSg6ezAeFH72dFU/N4Se0xfhA5TNGk
rX5q+j/FXPO5Wd9yAX9psBnQk9X2UHzhHZybKjk1yM4SbxpieoJGP9ETuUV7NEJiQu6tRtcx6Ddw
Tq4/LahwpJosB0G2vZzRIgSo0yTkbXdkdKiUgsqos6bXUQ3haE1EkBkQh4GzxmQwxFPO686lsObO
hY+pQoT5FUSGEz5WKTUHRnhVATWwVSNwQDu/o930nE6dO/QDUhwzvSpegCKR6Tr7cYxFlYvXsYWD
nN4NhwXpT3kxhqBpXFDbwh7vMCHdc3pasRCMIDxJso7dc9khALmolIYZ6SZf2Se9hqqT3O94wbRk
O8xOoCdcPrDBYQKOh7r+QdpIW8tr+DWlt1iBdYzWyFLAk/H91B0tZc0b1nbNc4y8K2mt8v1FrHwS
Ri9NJXhXxRdIKqZTcmlDkB00NDvJSM2OattqZHCVp96elvZqWBV3KbFE+EBh/8ZgMD95EdO7bb9U
MVgngpNsuz/CJTDIT4lqqKUz2m5/whlSTrEB1MWnxH3LpdjYhIe6Oh6V+SVpa3Qq3kDkuC64sdkb
jsMqbMi8hkZ1nEFz8UvjXhOxRNm6v40HxP53n2FqbhUFMT55oGssR9ppFVdnoPLJohWtnwj/ci0d
WgVsJIbHpexxqBr1/WtSUvar6s5uoljolv9ry/nyH9NsT5V0hkM+3rLBjZlQQ8V6bYYyNX3+0HWQ
dVSLZCrefVZXyLC9tVx4Gsj066GmSrESCObc6wDbFU9u1eWy9odqul5eLMf3lXaMmND2hlnp6PpA
woXCH7Q+k9jwCabswqsH4UnG+s0fblvktBtjf7iskNwMD5eX32CW314hBfJHIS+eoups2eKxmqpr
v3NdBAMS5ZB/hpfNEbO9tdoDCerMyi9TkqPGNjkNKj6XxKpGfjkeBEkHk3lGHXmEvJC7ooPgxJzj
Khi2wzdn/5JEWIwd0sIeq2aANsU5ZeS5Sx7UOxhczRp8qKgWaCSSsSREFqJk5mn7UwX0+I5zpaVO
co9uZ2S9PZBT4/ACRp30wRNuSN0fHe/bsMdn4AN4bbgsSeNKMmuwRbrJlWDLCxkEP7+xo8m088NO
GWPP59rLKhUBR4frTez724coIhocnbqnIjMclh6qgdrAThlwbo7b5/HJZ3B07p4TKmnwG5Od/NmZ
ssJZX2wk7RZwMslDojdAc+AzWlFtyHF8gfQRgsjJDaOHfT9yNgWPV/Vsc6KQhQ+DuHZw0XAPdM4P
SX9IB/sTfcxquLNkDTdP8A8eFAcVhWPPjBd8/pAh0ty4f8+xLORzzmS3wtmuqW8YDPrftPnJbWK3
1KuCK0QsN7KFQehYmCIhy3w/kYsak6j2MaZwjHXISBHiVv1XfxSgjKI4tbB9P7IHBqUEueVcUWgN
+Oc10CIqAxgceiyb/P/5zgi5gNN4aYG59Hlq7GdjLYWiJP127O/UXNhVW+61h6gABjWTIZBLrLUc
ocehrTBVNwij2m8Hmx2e9PmLmwI3gbinFZD5q/RrTFRvlnMOLXVwn5xlmOzUBliZWQrDwkjFi5Ly
Nhfcm0IZc5Q5GHOMZv34qwYWc5TIpPoC55k2CnHw/zc3MnSwhC+NcEkzSFwLWJ2TxlsDBYJkXLrO
5Stl/ICZ2u/QCyCgCN18qgz1dmgZEvXCWqPp3pBfZMIwBaYPl8HtVHGUuekz85PI8iqlsCBy3Nk+
UsgJrUw0MQw7uLMc0ItOBYjvND0IyIJYhggTyOoqLOHrL8qfy27I43xT+sGxfoKocwVcck3tymAO
G57GBtg53xdYoPqyIpIwPWpvQ/TsT2Vd6d9GsoSxBHQzfyj3iX0N2tWIOHX38e2eLvhp3Bqp2v8o
doOtgpQWx5YIM0KauLQEikCU3JGo84JZUjoEF5CSAfLz4NmZROTyKhXDCrDNSEmscawqH9RVSVEc
L0uPvQmVOJMLV1WW7hKVErhICQejabd7Nj3QhNhfIP+BUR8dNhd4Tq13y+wNPxS3huZPOyYSLtEx
Vz1pthwYGnEYT1OnoT1WdIx6dTnFt1oCk49d1rhvbfnwNs99i2reD7CGyp8eFqQ70cJQkicz3B06
82zzOARpoEgroHnM6e5Gu6tHuIq9K4XcL4KBClGd5rrzbX1sFPMy//yZDKQu4a8NYkIFkj6GMMWx
PI+Auans4HX6jN4vFdWRc4+8dz2uXAv3hlN5ozYACO02mJEibuEvJqwylyr6nQwa6dzpwjI8dl/L
Z1b877D4ZfwnYLAyoyvGIAE1oJSxJ3Q2PFPyG8bP8jnpJFxNFP6+oE5jciBOBysi2cwKVukd+pFJ
STSNSZ8DgDU0CNMObVfJalrcvHG5n5pvSjAJ0Z8EVlV+NpfoDZBg82A2L920z2fGrpZPiFav+oLQ
niuSWSev4gR9WRXAtwmah0gkRmV6Kr7mp41G23fNIHsUUBz57KX9UK5mhvRkfRl4CI7w+USLZ/O5
IWWYAVcxSkiYBJVm0DHC3hm7DCGISeqOb5xKVtTbzE9yyTa/zR3IZUouP6yMuulHYj13WgWlAuhm
8CO2Fyiz/HzOf/l2LOWpbGb26MIyG02hihDpYCRLvmOPJYOq89Kd/cYiJxwPu3yUefDXxxdI4mjw
EDm7Pdlr2SQ4NW+woIj8286jAt8RmozfTN4xOKHSSwMLuazFo+DSo6c9XnwR2TCmsNaEeD7ORpQg
isNQkCDsfioTHFE+oDLAj/2f8k/XklGge32sy62jvPrfCWAdig+9Zz9PIO8tf8B7yu0h9SUCf1zS
HxWeKUavWqb7GE93RU7vBz9CukoQRxYLMcdCJFQpFHu+0NM4ugdpxI9fFHk5mW/LUdw5DXd8486V
/KgQTaAnV7FedbalGKywig4eiwevpY5M2vf241k3nJ96DdQB8Zn4mDHAQGRez1QvWawNlrWaWIPz
HYh0/6RlknpLQDQQv0c4FSgOn0LxzriPbZiJk9CJfeSFNnmFJ2NMMO75l9f8qC+vCXK9RN7QPpYc
TC73xjJASuoUuemKDC+MQHLh7BbwIq8by1BD0InPv9QSjwgFwAoViAuWZnhSECHeEoV968ueJyOQ
6cvPoJRO+GWn+2b/cd+il+dYC3PbsdPLhYl+fC02sbkpyArylF8sAXnEmP1XR5d8sGJ0dg0mDLA6
jAWDiKhxkLP+H6olrPJLed4y4n+u2R+b8S/EnrHX9ktqdDVHSoasrP+4wz+HSfuyl4vg2mlC3W//
y5/6Lz/OTM+9LihCyOq4rqGH7EGtsB92U5bRnvWgKESy+UROfeYe2al/Z43v1ZXYhMVJNXgVmVT4
HIVmk5rMDcsYyf86CwTPQVVx4xIwUAwNYzRC+C3iSIIF8jlxjhb/bbJdkgzMmCIUKAz27oiDhKu1
9wR+eWxjY9qeLulabkaHezO/FVq7Gyvt4mEhxt+O/NN51ahk/asm3rUIStGjWCdEpxH3Iqxu2E8x
mHLJsUtuxNYVdQaAPUZVAVpSGCjqqu9zhNbEeO/WhCG00Z7EpB1sylQuVri/x9vf9MbVRSFU0hdD
RK33M5hYfd1PC3oAxzCLTHEtHJHICRCEwOc975DWSDFBHUi95ep3rmaba1g3E35n6f1WmG+r06oW
/ogos5Aq72Rjz4AO3x+QqPe+mWAN4fvhWhlXeY5uQQ53A4G+Rrna9kFUyvfGsNB784RUje6yqXXB
NhcW0kHtw87o1Dy+/6xsNCH4z48G0/GS6yAhHaHku0TfpZvtuHaSHQMeqX2QtAb4FryXLZz3pH9g
9a2OAC6BkYdajJibQbedv2KrNKk0Jx8TmTFucsD8lLxowkHIgPnTwuzp8twI+pYmaTsG8+d429xz
LcLip1jAwqoEv6H0qCeQWG8pjH/mNfGuDtq34VOaPggwc6eNjUFGStoEnIo+ZNPuZQmFevJCq8vr
C6aOBUbd2BIzUtOShpLsvGF+O2sTHzMK3IAKtvzA4Rw791i5GHdzcsbPZ22WZbxEjJtz8z/BozoM
diMRWxxlPN38tHivVorOa7CZKGCWBMdlSOpVBxPZjH257Ihha4u3ZVHIqulUWNVLXbC9LAd6shoQ
8FDnRFHQmDNI9+JrlxZ/J69+pptOrWVOS3X0mxKJLi7nbudhCieK7CeLoWnvpyvITaAOJD0lbw1e
ofuxomst9BgSnyfiCKPtUXv2bR7ufReBkwv2sU70LCWuMYdrp0lOo3Z83cGYUDtv9Urag3jxTX/M
BpPvpT10LG1ys7sJmg5OSlK8irTQ0ZiMxbeT8ySFMO6iHtt+VhHxqst8qAMXxm/W9d1nr8dZ3n9u
6A1dSrg6O/TAnk6YFTwAv7qdRgFNoxD8H5cYtuSkzV3fds2y7J4COPKUMq7Cbec0nedidfXGVCSM
jI++EKKF42TxWmpswZixC1oNxNOi4vZz2dGaV85D4GpAEQ8bJPsCZsxlPn/mLNU6kWQZIQKoYyFU
lSbyjlVTd8B0A1Ze0R3LoV9rmFNfg5HBLEWcOoCf1Omp5Lat0fqCUfo97u4sekmi2TwztccFZF+S
4/JmUfVsaRZ1N7GbYDtoo6WtraB4icBHdEwrSRqVY0B59bT5ehUKPFkLbUUS4KmeZo08ZadDihYY
2zaS5VJk2zLsY76vTtaYblKZ0F3Z8u62qVs9COtxtgScLQOXQ2z9cD/YUblWpvgYzwEvszItihbL
xUVOThJ9j20P5jMpIIQ34OEhlEAWOvaV0CczT5SBkTBHOR2Bs3Xz56rYpFgiHfKugmwe9zDzjlSS
pPfRTK2Fh/raRWkFdlxPKVMw+UtVffdx6ZmkG3ivF9kajhSOZLV4Onr/DatVtMMZy3Pqy9L76i2G
9kNg4AdkxsbWI1XYpCqOSjEQWefm3yBii7Tf6SnbBhTkTKU9pipcg+BevjflseFs2t4zS8ubbb8i
EILYocFA9vQ3x2tADztMuvTAjh5KOT3sSdoxzUFVPA/Jivj34CIVEDg1ClQpSRlfwCGs5OdLjiS3
BvZvOjY8Z3ntkUnUgQbml1HE7iUpAUfQJkAZ0hRzo/XKEyPKH0U5WtJFslBHcp4aWBQ78bZ6+LOh
ZwlarqWlbeQ0Aacw/np/rMoSAbqWKOqQcU64tKXlS0xsorvwEalloJjBRIpfgEc0FHRyO4FRd5nH
5SizAqeq2m6EuI61RPjY8pO8fsWI4cmmo2myouwV9JpAtVYSF/koDs0g5StEtguqIF9mD9vtepNm
lzVSaKRGpCXO/YwXq7tgnmOKDK8KaZVgc0etG6ABOwF4Rw5BuleJSX6It+uDgcB3OaUUDT1DNu+S
97qHffhaJxizVb+b5GfT4/dBBzRXO4vdQYxkyiuf5Jjt+kOSMthLCJkR7QoWozU3ixY5Grtlsp4A
3YIIPxlnPKORQ9Fsfm1itTR25qzU7tD3VulE/9hjymjOsXefk+PhJ5R1NCRy7T002iv6CqLBH3Yg
wcFOw+KeQcikoVrNhHBzG3KjnJUNZ2RhiFCbI8Zq8iPVVBkyPW3+ClBjauRPkGmmodHJq3a4uTEU
AT8YKwhRjQ82TQ03T6tN600XmI+JLPklR922Z4B7rO4aLOQJ7Y0fTL9MVSylIoPLPeMzlUkkK93o
/UZP+qjLVTscCAk/ISJ59sje1roBwydr5Y+91sf7qXrt7KUcFy8CV82DHKO9OucFR9dI6izxr2pF
cVTVU8zFX9xQ5/v7adK0h2UMqgW7kPVuz6Ri9BpYzQfsjno48slo7OmGvET5zACJgoZioVGrvQG8
A0YQv/DLZwGeDlluXlZVV1U9AK/K2yohB3GeX4ERhgKmsrK7dSaKRJCeeyFK0PGtPGQoVR3D5G38
03OB349kvYRKGKn8oR2juVBkUdkwqQrriiKp5kbAuenzUSwE41Oash1DYY4qUnBL7c53qeV0jlB1
6ADYldHoZQLidN5TCOenToqbusr8SqHRdES0G0kxtMnKQEJFG6xsa+qN0bvdFCCp02733nw/rZo0
7guKy73feAYEbDWxJ+Q1AYnMXuGcda/1beCtGJFa23cQy8iTXC2ol4hg5GkB3b0WyjiT+HpyipAb
Q8ihx3YpQI797goPkNKco/awbkyT3/Ba/0rj0iYUXuAXI5hA7mAoLvVG9jFdJtORRMF3Cm/OyYQM
rwj22qr04OXF7mKF9XOLOYZvTRlAZRAgHy+zNNy7grkO9BT6yXrMHgK8ZVKcAuxPAY1J39AQWCe9
ZF1BQ/BXNvaDJ6U0X5XAdsdtUQE3qKFKhcsmhpuFdtWN8cFrE+NfAKdtro3bkf4ckU5hYSv9Sf4n
mWEG6wSxMqdkGc8g8OdXtWJTXCGYMr3iWNUhGagEGRXEbxOMwm9Cnj+9w/sBeRzrBGz4TIlrAwie
4fuRl+y8SCE8Dqn0dGX0DDMlC53whz59274dqlY+o8RTPo2PR1l7YMBUS6kjBYARkSjnbmyA8GcL
Oc4viJ9yCzbyotAO0KSzH95bBHKak08Z60L8kBRVJh6e62M9xxMk1XsTPTDLuZ2hscY8SluYuLik
dkl59vvxps2Zpz7GBbXgwYPqY2h5Mxqx/WFCTYvCMLbKSmiUa47heN5TkpBUyrnmK5CLuuxvpVKc
ppiKjOq0PiNzG7kywi0ySV5Umho0c3wulh+F8DxS41WGUnrzJVjbVjLoFZoR8SKblrB6FHQZNvP5
N28Iw1eEYN3VPh69Jg5wcNavl6XQRn1MfJmtF6tkKwHUb5in3R/+7Y+K+D9/3uNZFMufwVIVZBAD
j3npihfAf59D1v0UAaBDIurC1mGGsNywZglih+83PIPuSZC/PT02k+/1FR52nlv35Mx6i6lvX1NG
Rq7GV/KjLIRXSiWKr27MQtuJTfzxQ2ILOxr4LXp9tGhxfk4yrmN0uXV996YXm8r6XuuZ/sg95PoN
bz/d/TN5mnC1yO1NKE4yBkwrYOVznyTl5uiaysgQV+tSyIC6PXi4nFCq4xC0fNORQPOxg6HeTTD/
e0ihoT+ycb2p48KoDqksxeoLUfBddubxIbGGtrlT4L/40vFqcVId7eqIXEuHVZLtsLqQgz9l9aWZ
CIFyjMhS5gj/uCItP56rFauu81YUHjsGsIhufz/vpd9ElieVkqP40BUSofjrUnE81EbYlx6Nx5ws
YCVfgwtSujW8/lYHl7Fnb2GfJoM1xrrnlefhEmWvCs+4/QbOQAshJKOmFHuhwnkIRe7gIRkSFhkI
koRGC801dMd5XcfFHTl6PVRuNdqV+yZ4URywpfityBsWl3msiThHW9exa5OoeGWsuHBWxNa2kIk3
3ZfuZUO8R5mGZlBwBM8EuszSeCV5IF6b3zxugwsBoulQ+35X6260MgeXfvJKI32YBEYpD1DqvTcs
UoMq+TRcFXALMzIXLEG1goLu1gZyxWF1f6oiQ+1hbWBdJfYRgKw6Pkq+d8Xb6CBY8w7ZCUV7JgZs
7DC7eRVtlF1OED4x+wK/JW5ji8Y+GSMzeoLEii+sKsyJCAiUrOIjhVhedYPSv1XQTDslfPhNE05u
M1JXZ4iX+2W3Z/SzRodNLm4s+VjRrj9sV2Jh9RrvZBHTaabdbzW/v4AH64QuU1+z/90ey8GRwNYe
RkTR0sHVhSyKFJOUhHSWBtT7LkjcXdSCN74IPz/gCCeBMn9xDvHAsjueIb1nmx4Hg9ZtaUjNu63+
40YG4lDxeB3TMd3iM4EaBNdIuFAGHGlPwRGi3dlU36tkLggD7EoZwsVgWIqnqw43tdkwp9cdnvly
q/jFw0vJzlbC4VCMmdbYOF2gQr0qBfkqLqhc2pusX/BtBcYWls8clhJ/TdICNuto590s+4f52A/C
SmeC2dt4qjhg0vQxJJl+7h1eM5ofpq8c/6DDK/v9aKzQeZq29KOtsVr1NQ7TXcamC4PcZmJZGuD3
TuKAEcLG/YBp0IPZ8Fb6M4+kZaPqcTC8zvsrKaPWNp2TLlLaYxMJzhj6+8c5PI8gTDENrHmxVm/6
TQevLhmU3BNEK8iSHRYWMSbmCnEulTQxK6RjWGHbMZF4BkzvOvdRXWrbwfxxxUhi3uf5ypsUmYy+
vhbfwVDlZTYJWKFgTdrjANmEa+RzzuIDJnHGjh32QOVPl5K9ICc+SWgsourOCoV5AAGLEU5t3sPs
odko7oFP+rccPp8IpQt+W5Eo0DlHLwmbQevc9dJc3nLzgtgEH4DDlHBvr0PAZsBzMOyRxUE0f0OG
RMI30hkIs6AJYcWRB8UxAjs1AWZ/GNmRckbDGBQfafdYydM4tHXYnmPNFHuFEqisr3zaGGdryXu8
65licjh0wV9eEjsvhu4Jbbpoae9P/7L20RYKWzp9pEt6lWUACCFCKdzKi39H3sryOzbWfceisJxR
7bdYKz6MUj+imCtKqq/ydtFyC8+9p1hjAXL72ARLLBssAcvuqgwRs/cmqdrkZLTDNDSH1lbtMpW4
UDUh9St6SloUCKoP2dQm/pIE028on8OITDd6NC8ryBCJslvJqRdJNNb5lLu9J7JhDWTzJ5SsCo95
jbe3EykGnUWHaW/Oj0JQo405XjLOfC7lhSSdMcQybFi/s16/DrdbXWwA/F+VpMKOnnQwRe7d3+qb
0OXIVbFZB+Png8UhS9a3LTrCfEb2vUQUvsArtVMI4XqO5OTa36/lhc7aEPAYuG7b+htvcbR8C5MK
BgW2mTwtOnGIk1KrA98/AOTqqS64feVvBJJSgSy0feMN864ib4ztkfXWS1w8qjDWgb+tJb3bnGrD
tsPYkPY9Tu+GqlhpLyPtRmcxu9vp9WXMNrJ5GOAKOSrHVq5WEkDoJ2Q0hUT2ws1AkL9lJ+yxhcp2
QJRbIoma0aKA5KyIbM0lzjSYGjXqY3lpXUEro81qxqSBDAgtxZjztFRY5FwIvHMgMKrc4/38aDXv
dYAuUBeEy95tRYiFuzjcDZCgCulBdPchsxUJ03MKL1EOqeM72bypWrOi7ThQhHOjS40QbZvlhOyG
wKNX/4K6cWkoUntOlvEmd87mEdQOi33Jrc0E3xjIA67cw+xh4FNZJFhEmOVq0tWArifPwNojOwcx
UQvCQJNU6wZJtNRkQu3hqSNg5z9A7b4egw+JlqCdFfVd8SM37wXsHsk8xbCyl5vqkQ6a5ijcWocv
TS/69DQ+1app1znSIaIYhqar5sRgYVcCPPAqt7UzxE20vD8iCyPosabQB5LpqbKbajCkDg9NGjbD
id9mY2bakqJgpzCHO+NlnZGUy2oSLKCf2BNrPcm9IdLb7bLKjfEEdYjgfC2PvDDkC60hd3MfSbM+
9SNULiPrRtqeTmG2/klnylcsd0xI1Umxd/sb8oaVfXpAH62P9ipe1zn7awHa6fjMZvjwO168aFlp
Rcr5ZbV0b37lJQE7JcSnTPzAShjf08cywBVTU37+6sFQL/+EtOO+X3gPbohjg9Jlg4KKc6Qczwrn
aH96JLsoGajphkop/T7JsIr+FL8jiAuI2rA5GE/Vb0DUpsqRpnJiN5ZzhMPwS1tYXM/cCrLznwUO
lnWh5PRljFaTA0ea1Byad7wNmrTxaagnAzSbzULHutCE1YLowwH+EN7kGSPqad1TFTl7VSOrMRUm
o9W5akEYY3sATe7yVHXxLEZp/UHdxz1Hdc7B+8Pwkna4PkFIBV8hXs4IG3YpvwGrYKtFCc/rid/8
vd2GrGEvVKiGyjakvWafozoQjDgTzSE1xLWzd1efmCyg8AaeWO4AJsNPlNnQcIZRUKJfZ07swfoq
HkpjHAf//gGvQ8qX+qkqxFOyine/lzp0jNQixXP2NA2pjhLQITbvySP5IickAn7gmfaLULAeHL1V
Bq8a57hJ4gr0K3nv0fR3TNxbOr3Z5Qwdf5Irba/xaUpUBaF6Mv5ZNzExdKvRBDW9r98dT+T9qNO4
DM7E7NTZXPoaudEP+D0Pcni79CpdtDxjWBMKcWcE95K1F83O+n/sSi+NcK1VTVR+cxMsVFZwmUYj
ilNn6rOqmnQ7jgAtgcJ7DfFjq+FmdvxWkbZ3zQM/uA5HVkN8PwiI08gYD/kwVgYwG1qPCtEjZ/Nb
YX4nm3drBim5ljWdIo9nqV0QY7WuagqQpfivLBL9MAjo9FN6FjrclMCipX7/bGoaY61gbMFlvmkg
1WJ+Ab/Omp4NSCCpF+MWCWO9NEqS6W/SxwDYeboseihT556B9xzuw46lf5XI3J/Mwz2dpryPt/7X
7bWZAGt45gr8apUMi/A9vpR91ASTxKzrBN9ivxEL+TGVScrWNREo1DVC6Nkpk7G99VAjvXvhEZEr
C7dsgWZls3WxRT5wsKxM/A5otpplsmBU6koZkMFfaPBUaFnVg7/Ve0td9FqJLzbGN7iee1UdVHn3
wjxKxzh+JqmVSvQmACAIo1ZiGwOjD9Zim5H4h0no+GlVAquWwixMN8c/XN/ZXprKTnIEvCSYVyAI
tpm+0gV6fumNeMvFuctbZpN4TEukQVWUBj7sESyVB9c/DXqGryfdFvf9wSua7Mxpaciy19wPcipb
5e64kHAFfM4vHCDg5efW05vr2N71iKCgPDAeeD6Vdab2fDjvTLAV1HKLeiRYteHR63YCmHpMZG0n
ZQi/WlkO0wEl75QapcaWm0HGIOdXMNuIaCBUKyPiamQ/qGx6Ahlfauc3VwGc/kHMHPU3ZMNdRXUP
qWgGEdNHQJ+P62Mr/t/DoPbCM4T1uOACodx4EDAUEQF5FHVKqjLv5oKrqOguxTD5ctwakbhKwpch
WCWUUx1bJ3VV+e1qJh9M/e9gCy01Pemr6qq9tDki4MPvUUn70nv2LvOhJUXWc/wIhkmBU2mGk7kP
SPGnNkCcKoHOtIF8AFL9A96VaHLsF2oR3dXmJ1WVFeG0u95XSeEzd+Rxj1djc9rMKYCZSamhUWxn
R/cNAJ5Qd3pnDIbU0Zh6coHvXOLWo83fRMKd2T3xvsPVhmS29VyN56SRN8hJXaA6xcYxlo+FHkiT
TrIkgnDnh/66frdLp5dubFq4tzAOqsDHxWbRY8aU6h/5xrfshjhjLxgsqDruwQTgT7QtmBLmzY1o
mQnqXsgn8upqJduHGn2wcXXHEkwzYw1w1Lieowg9Y1SzFbq24ufxYGEeqr74Vym3kA8pk9ipo97K
o/C4E30N74908IP+ZVhwpsKKlVfmJg2I5X0CUBKqHpAw2+koqaxsB6f2zFbFsuKuMMUT4wMDNu53
DJnVoCyQWiLPgA+i1lTL+SZZlCC9p/wO+kqrS9NujixSHB/f3Fut7a3x38e3mMx7+/QwrPJyNzle
TFV80iK90yUrKkko0ZNcvObDREebDadzjV6xnXtSZoSdyfYYNqqM72eJHNHevn0jkCHp7xxQ8Tqr
H2IGEgts1BdqTjUdQOxrcMSOwFcIBQgUEdZz38r6g0cJ+Wtbpg2Rxh8xNh/I9UaHVsJv+xuxH+wm
bBJdrY/+YxKm2Jalp7RD/aa1Sx98Q6nvnmdwvic77DkAhyMDbXO59VoGUg60ZJ5B06I9nDXpJfTb
Lnnu3NcURykkChPcng1bFEecZDGY0xQOnMNHKyYlDrLGiSihr4cioP/0Fc1IJdAK7BjQYttVD6Qw
eeFFuo/lDyfFNeEF76YxaGi4h5SxsrMYkAHJ8coEXHW2dhVq1aJhDwXKXpSpMskZAEawEVouFPgq
V1CJ/IG9MBA6o5logH0vw/k7dKp5EBAE60E/xgU79c9Bnv8E2VidU6nQgq6I6Tuq/K6/xzpNR4Ir
gXL4uQ3cWezAyj8KyON1+5JQJtA1iWdQOlH/tDgZMxBb3fkPfneVZdsJdh6LJQvfNRV0q9VTGWLa
b0MoliHyhMIXL32V10vWb8ejTZNASArf7FBv3YAWB6SqD91X9pKorV/kFumnqt14Qp2zI/CjJG0U
Ztu/eSse+QsTIlq/kTiziGDMDw8uGR+87M3XwKrmrv/Y2rlNNzEh+3afsf7GRu0QMU8XTIVXLqRp
YtU1X+jlZXQl66xuVQNC3kRYNzWfCCjVh8mMce8ZEm/gwJ2Yz0qVX9+HLMktj9tafAfbB2+e/9UD
V9Jpcdx5UM/h9EYE0kOG53TkQ+Q0bm9w01BPbALHpxIrZBlI4GlrvK2FJx2Nl1vI/mKagx4UOhiy
iPrBzyYyxiBSgD7SK7pRxL2SttXdNjzQW56Thh3TAZmSrsK9vpTHsh8ZTk+1rxikKzV8JG4KmyOP
nc/TAALYwL+mvvmmqjm07RxEQU6OXAOGzeUKK8i434nnVsgcifulx4sYomDNqxQb3xGZZFDyBBjT
BfepkcG7sFKKnvyhh+vjFML2ZYQySXfygb9272cH3iuh4x8gdbjf044/YsIU636UuHBnOCNb/JMu
8rTpVw2bWJAJO9u9VtSduQhsfKgMsRL7W/VV+zXvYoUyknhsei8mLz6dbCI5WgLGNvc31rnly+PO
pd999pKfunGFdo2AVYsO3zaviwRgacJ2tDw0Wjn267ZCA+umo7I5OIPa1KcMZ+aOFnAXHKSw2PJM
6L5DpN5xKbpv6nUiIMH/PNu8KSQ+I+bra/ogclOh12iUpTlEGQw5Trg+rXLvE++2QFg/ClGcGyog
vCPzHKtNpHAT5dLcNWt0tPPmDvPt1PZ3niFLtkOlIK0W3q9iN6Yix4abggAwx3xQ5BeZUv/sw0GT
9vZ76ODxhzxr7mbrU7mUZg2p20WuMY4ECWscsvKCeOC8goI4/EPFtqNP4HvjkC4k/3sf9DaMa8ci
1qP7V/IUQHNmMHDdGiZHVotqs91Jw/X0bMI8eolU7Hpa1XF0gT2ZVESOopFpE9sols1w/FEwtjrb
7kyrySxBaFsabwW81XVrWX8oPn3FWDY6KBGk6a8Aaq1NfDjkzJq9TTf7NP8nB37tMpKNxRoaCpft
ScjuMvJAlzfRolknq5qdtOfd3XtkcvsC+5gWGvf92KquluAmYp3ejBfBB0AkRfzjIc8kst+M4CZT
e5vl4LUZJxcdSc0eVzt+2JHRNpAeXSz70HGRtW70I2DQudhNYx+NdhnidDO6RPzUUMavBS12yqnh
OORIbBt/AlpopgqWrHKdvToV6ytfZvhZgfc6pZ7V2LnlZZTeWr2a6MWNdxaamYUnrwU4mW+8a8Pg
mNGQjWzW+cg/40bvKQPRK2BEXWot/093OOXRkl8nRdohJ0cO8l+ht0FkFC6tMCV09mXhZxNOmO3S
g4/Ix5r1pUKFX4Iu9HanPQV0rGLFAF6KIM4rGhjhQbURNcUT09HaJW/SN4nLLSOgOc/1jjoVdlJK
BCsY9COslm3GZm2DD4MenMPWuViqlHgjMUeoQ8fdzqTQCLjgqOISVBTpFk6IMXDPp4JkJwU7fM81
Edw3Ul/FnRM/PJApKLIMgYozvtDYAoZ12kG3T/jOnAhBVDJS/1yu/OIAojwCIKtsaVgSk73cfI9z
aOkn+zKPbIkV/RmjhpuyhJSNEsjgx9+64Nd4PRLIXLPfna/ShVr71dRGuWB70vHI9dsaR3Djgwzh
2qnGMsb31AMNK44nX7OSDAtIPYaiK48vq5SpXR9SyxwqGm9CwyodFtx3q4ez7ynobyFbJVexwhMs
skraKZYCTXCaZS0wf170s1i8IaPSp7INTBjG3Be/4AfQwThx9IpnnTSVMZOVNoCOSlMvRxdegroG
BV8iDVbKcDR415wGsrHIFC3WYREhpp5TsLZuVRivOUtnyOuYIsp5GxCxGnwzRV+HOVngw2ECnL2s
QxM4CVkzmaVvEIPGfQQX6YurNTYc/+lhUnIJyCazXX46yTjihTdbHXkBCQN//yDCnyvw1dAjhQCQ
xTUocinCl5nAZypl34b+KbBotcAtecfl6FgBpALQtMGh4+rDWOS10EfzLwQ6cD7x+gLJ6G/FW9yW
iWLlbgPqSlxVZjn7+p0flWxERf4iwJQiRwGpKgR3nzzEu4obRWxMSmZ466LsAX6I8dDHZQEc64mr
BMNXyExgvXHLvrtBVRQd8t227vOhs3K/iBdKIBrG0fX3LdvdmEdoW2B3IEt9vyE2F7KftmLf80/8
CErI0yUdikU1t3vLUYXQMhmS7U9FghXex5uL7vz2HpH7kpmzbmxUon3E209yyn3D1yPqia4aq5Fz
hGOM/pQKd1ad+O68FOTJTxc2OH0fPonsVlRju02BFnwqQEhaLuievT8Kwyx90dDOLganXCk+/a97
j5hfJBSUqH9BdIY3KnLLBxel/4C2qTB0tpzMFLcrDDZTFErQoiRAp5dI9eDyl6WpRR8jT7PmhehS
/fUpdbm/yj2vYClKUaNVDep8+Nspi2N3yEr3p3t2lkN9Hn8LA6hBeWRz0lHkH14InVTPkdF6WQoG
DNhZxV1m9DgxVdD7VpD5T1rrbYMSyXlRcL1CvY06IbQHZ9Y4dWU5gjb38vfYNpaODB2qXiu5vjKo
C8ekh1gq2pldoLMmmbFyvHsh4yX2E8MZ4diE26cXERwvdE0kBFg3A8H4VKwnk/HTRnopC8JTWqny
aP98zsmXdXRbLZ0Iivk63UEnKl7CNzeX4grViZMU51NPoSpkyzHQ4w5xQi/nLC+DEKPVPY/Z2GvB
GOix/vXi7R0nosYpglKmARSCXPwnRXzLsxr6rcMDTXCnF+N0XZ2TY852y+4Lk1UaNt9XSAULT3TJ
wHAYbf3xundln8cbcPUjmkS4NFRoiR9xa+XUXcv7Cr77jOM4ob+9heRThdvZOCoJOmpxLvM/TDQZ
APls80zbriiKCFRTXDCIlER1UqkfHR1CHMuDCNlm5oJcPclQCEQSqyzevCGrn3AMRKuDGKv5HBtZ
Ed6Z/jo0AcKYzDN5w7GDKRsIQFkgTZ80+EPQV+vAzIaMCTPWYdWWffnET4zBQdrms+aItuNGLDWz
0uCub3OOeBe6zEVwQefa9BQi/SZnDKfxMJYfrKOlEILZ6kG/lsp+FdedHihr8l1kwUH7oUJqMUaG
9OSidEU2pQ2feK7sUiypWjakCrcPcpoZiOmpRY35HY5rcpKtL/4fu6mQ8mzaRi8DNsiEgs2bfwP/
69RaheEVFvaPXHTveaLe2P8FZYmPRS2Jgg0KDa3sDeafVDH0LWr2CYpvmhJk7ZUDfIhyMDmZIeog
srUMb8PV/oekhg678TdeUQ2/Mj4wcTucHc8/IXazuAXITA83U7BRfYylActS9LrLqUJjcB1YleIO
6DhW0WK41s2k/HMnRzc3vw+qDbq6seuzxwCyvBd7oY1nWZSNu2UIdw4D+WNTH1LVSvf25EvvjcHc
QeZkypA0krrk9Px9zK6zyp/Dxnps+zYrDRBgj/qRyjqtNrcq7njLo0vdRjN1NWd7DXXd80ONiW7e
7WmjW7SzGsfWjcdUonE6R+vlx4AUTzdWL1bVscQFi4/0GTqMKzA/vjowpd/1m1y+BlnxHjA4EM32
zpGSsNJM+Fx3WNBcNWe4VLBb3l2+LbI0OgygZENmgWRkhFFrAvGxy5DPwrlNZYI1npaTDykR/xZ/
Rgb8jZG+4NSnSlE1CCa8gP/7uVEpeTGlSjG6CF4JJ6RGv7SMQAtPRMtvOngGkVoxG1mFOSKFd6jY
r+anq0I9kAbluOTjkwZ2wO8C02zz8gDR7oZ7VNKd9sFLZyUgSB9z3RtnB6zzbDvXy8+HTEjltvJ2
9YjDjPsxmSqJzfwLerBzYp6a8kwdKiR4ts4sIpHzbDKe5U1KH7+FzllaeJJ7aCqmyALAaoLHEp6Q
jT0eWxIk/6EhEbZISRSuJiyX8bnxMdUPA2hvWJANo82E2EnqHcF0ZoS7aUCwZn1Ls5uT0JUfqDhQ
AKu5NX6VH03dsbve4t1xgt5/mP6UxJ5cIFTWYdYHYWBr4vLvNXLf64BMhEPywh3IChh9z7XPN0qX
d3k2CugVzwG/yDG5yfjYLrgvsvoc+/mBUI8xrukO8C1m6t3I/RYyQ1/tHIAu72t39OGP9cOkHfEa
F7P6nxyPZXLIQ0D3anaxiN4uxMr1Y+QSBdsD13PTCizHEanUHP2GWk31lkZESmugPKmXZrbp2P6Y
Ak37C9pHeo1fSdQ2OKV2SYuXnHy08Krp77owgP3aMfYsZqw8gDtTapzqFLc1rtzRfa9qrg7nAk0d
qfUCvAKyEnjK4Mc57CR+YziPn3qCJHr7ssWxBNSa3d7r+LEo7Vmb8M6zS7YEmckbAfQeVxUVxNjE
4R4Y0uC+aUwXRct1t66BPTCJ5v5H1RvBknnONKSnVcL/rknp2+3OslP1CTLVwgzCZ21kBWzAHocP
mc3hCui3pY8KWierBcy8IwPMpKerb4ja04jjn9VXk1olMq+gi8ZmhNP/T+rMZYPj5+FKTPBrb9cB
/EebjxdTVy0K1H7LjR9wirH9V8KHNO6bzB1Xxf5CJIkZVi3C8g2L67DoF3MZx6XPKqxMjCWSBxPT
FVfY097kXOT9/YfEChnYKFgVHBAxU8U3zgSzexad+Dc30KAM1HCPAeeAxJgeT5Izxkha/ONUmfrR
A6+IvSnXJCxdTCpVub3/6n+PX7PqZGpfppOtNcLRExhdee3mxH/NEzC+LxpeE4a/z/G1RJSNFR4O
CsSwYFAuK8a5Ynggxaldgt2cA6tpLuGkI5wQf0n3nWGwYA1UHqbxkZVllAWJZaNFcTiM/oJx2XoQ
epeUof/1plI7U4DUnEpT+/9ZJCw0ty/IHn+9wcCkRdXM/7Jc1cmheQOIqX8deLDMbOB0UjomGszP
KrpNneekA2rP4HfwALJQxlwVrBc98B3zaGG3otVopaetJi/Wvw4qNfpb2qbUq8DfN1RM7DA7qLQz
qCuZsPqcm3auD9ZjZIJ/lesg4hBNAonJ5qPh2b9K9Zc1YuPEobfT1ZUdPf0bFlHbQdxb4Mi1AxRu
0/hmQPQZ6lfMVcc/iFGnGAxkCoqYVG4IUvnyaUMXUf5y1dhlHC5bg89qa5o2sEGWoScyJeAbmPuO
T6nzblfpzOo4kbGCXQdcjnDSp0VqR91Wv4iTOIKrWLLHQkObTIiivMbNcgXV3Sbx2AZUF704AFB5
mgHX/Jcln6YUeo2hzTRKUHnRSk+2tHMpXAzOb+kfJXiMFnrCyOhg0N8GFED1/PxT1zG0S+m1TWqf
7AWpcj+p399sxsxGNrb/cYhP/RupLn6EUjPAnBmxuRqY+hj6rmoYmnLLJJ+/iPElT6RNiDZQz8gb
b6I7D8vWqI7WiZ60W8qkuyn7Q7Nnz4G6apGe5CtKjNoIjYj85zRlwvQlQUhSUq++lJ0pjv/o8RxR
Lwbvzpx+1BN1asCcbIFp3kZVZbW5Yl9EMazO7OtNF4v7Vzk51074DX968KoSZX7XGx3QtaUORb1o
xmx2F/j52uKfRnX2JZxucGaMYhm740JiumOry3ogB2A+m9NEE2YlXszNIaZBJQC/Cm/eJ6izTY5u
lK9gyaYHfvKpYb49fjBpgYLRJmmfxSw2KJ91S0gdDVzeOp6IntOI+E0BM9Olp2MQRLI6Gvs9nWcb
Ud4DW5E+Nlm80YUpx2hbUbOzulG1BVsHhtXT6u8Bp6GNU/BR1H+rYbYHhz+7VwatuUdmbDuFZ4VC
YYMExyYtE8EDUqeekZdwaFl00ejQDsohIhvrNvT+ltx1V4a9KrsxrL8Jd2B0VeLHH2dFbBnMAq2s
IHBh26JJjV+peIYJBzN+ehtPa2SuCCieTddhz2z9IkKxrZAxWqyPAmewEa+nvMVynPI5+0yxqzn7
H/bICKdHKHfh5zlNCWhiSEtseXbCPQpX3fKjT+hCUPAbcVeEOkQq9GRVUHZWfhkT92AblLcmOXdB
Oq+qyG3FC65h8WEaOwhfzewBraOWgSA4+BtsginApZ/9nZ42SEHrcIvv8SjDPTFsBN87aki5i/e8
KTGHlQret1kNvyiP/wL4Ev7ELruNjcKUn1uBUgndDULb5w8Erez8heDwKy5w1vOGI1hBSo2yrDqG
3mANNInQnUZ7AIDN4YZ297hcygmp3z7sRAlML7CtXQKmg/UOemd6U3RMq1cKx3PIXk2B3r55EJaP
8/DM7xMkXKJk6Dt8kg2C43gxyhX0+4hn4T4Xf227CPsefpTkx5m1lkU2lCO4QIg+49mXXfn3SYQt
Vp+G3lFJdyzxpnOT5MXi7/gRYhkLhOQ5VYvcxL0nbdHr2iY2YNmh4CTT2r/s5RCrHuz8vSI1rEMb
APmSQDzSj3wcFCACClVXxLz7fLs77+LjSofIlMAivXSWk0NF+F/irS/ESukuVcithj0NxjcfTplm
DX2lMb7Ww6/bzgsi3b/D/wcYDGwAR/POKaaSSBZUHJNvZWuneL/oHjHHAooInqwtkKmETDhuSIwK
e1gwEcdFIM4zUIiPW2UGq+4mXtJDTCKQ4lqvcg46/bt25sk6hTY5KI3bi397GtUIoKMLvBQXLRUi
df7+DK1EZ54E3iJuJaDJItwu+DoMDjbKHcn8hRUP7rmaQOUsjxmGf75eLCIeD5NEbNyEZDyY6PqW
KGvWGjxG4RRlLhSDu4OsTdWCqDgr7DW9gEGKI+FlwNUP6BlRLl/6QQLVq1/V03ySBrfXFq0OATlF
igNkjM5iXPAxazeksChN+cXczPPzr2chru1Lj6iiHMZKovFNYE5YbLCJJSHE0Wu/Q52BsZvFCmEW
fGkRUSkFykWJySJ025KdzgmYZMJqmdPY7wrnlmTuhFeelWJwReezeq7eYbNjSvcQpMKzE+HAAoSx
qjcL+QkJIZgOCQ45BtB7MKrpntnIAJmO32md2VJkfMKK4yC6jjPcEOMmirbebSViQFDtkbuwFgoJ
+WnH8LCl16PTCCuGqZ2xVa1iDQhVTkTuviSNHWBPZVYjgKZDyXOmr/PKp3RpsOZZin5QaIuTZp/p
nrVsQ7MiDl1QmZS5KziiDyjPIdViiN/9atDnx86rZLmmGaQ2Ue3OeyYket+UWVg/+sSHrEqVxOLE
4moijwaTigR96xPQT9vxK59x6H5EeLUVY7HM2ZRLuPwlOUDLS1KSitEj0d3Zg6Wm2Rr8D82qFKFQ
1iA4y7sELePtQiQjsNiEDamVs4XT/MBGrnBopZJTPyVOBK4BhVYtCT098p7DFK+IHwgVgSV0UIro
CXDirzLQTGwu5v2PKPqVrMlq7mOUw22DU14NW0hzDsq9SVLR0x+b3qQr9ICV7USvVgH2dG+d4uUO
17uI17NxjJfchIjAzX7Ya1E0NlG29baexlG4dKOjTZM2MNivo439n1BJR1mLjTSNCFgmWfe1MZK/
Zil1cOt/71vuGeJ06IT0c8b3jTlW/dEy60kpzvAflOL616C5m/sup/wWTaw7U2a8iE1i2kuz88yB
w3mxIIOkV77NOUR1mSDYikNtpItEh4TeG54P/NPksUK9tEqy4eAE/r2lu7GCnEiJHQEW1CT1J1YA
gE8D71ygB59klaYyeaRgjy1deoH3Jm/cuelDP7g+RfUEe3NiGzpy97eiKWzC9g4idhroaFdytVIl
K91t0BbiDl7Glq8vdVWk2RpJZ8PvY4leKfcXlTyvQkY7bGKdvvJDbF19VeZOiNq+tGV7vVUVteGD
cqIr2WLVyEQR4962yK/2EtVVT5iDosI48Oyq2400dnHtXObVl4Q0/s0aVtA++Q6NKAIZtms2ImLG
8mnf2iCY/MJ/ebb0vElIGazMpK/70ug4fyq/OLwxWk72RSXzJCOccPu0x5+OJ3PI7QupXP1uPC0Y
3AuT7LVVFxRbV0Rms3vOq/lrnCBBtMbvXWQ5FdI1qFIZc1oRvdVp/V+lBcaSynhz8Vw6/mOROlLP
7qvlBeR5sA3vm9Yhkl/zqel0QIKnLtwIchspw354EuhLcb8fj9Cvlxzy6i+ITvCzbtwf7EKlEVKe
6YK11pzaq8KbN66Tc0RrJntuTFeg+tUtZ4D9JrmnFcfuSi/5rQrgnGGHaBDfvxGrYotqiSZD2Tkj
9G1TSDd1LIUZ6/6mo4yp+jtW8xyHDJVkY+5BsvDsOLi86WjSBjvFaT+yGwZpo/UdCTceoqT7zpx0
06WqJm5HtEyCS3FjtfcLpq9JV9KRmWqfh/J1djVaCIdxHNhNQvWq2w05hU3785vsrh412sEtkosb
Fu9LECbKa8ED11olg3l7gY89dkiTbwFuO6fFyO0zw73uhkvmWaEvxZsLwPvzYlgqZP8FTe1YQjOg
/ou0UrQk89JNZ9p8PQ3/udBz9sli52737zvuerUCeYmZ4ZLukK6aoLmZ2w62Nrvmtao8kPp/lsA7
l7Jpl0RssyrOHIFEWcmE2g5iCiVLb6Qq0lcHdCl5/Zsrr3daWE+djPSIEm5clriqK4Ek9W5762GU
+pFUinEzVrrQM5W3UidWjIsaET8AaYJ0TMgiBGncNI+h6c+PmnLh+ankBW/UkjRIP8yiPPY51ebe
jfb4ahjprGcFK6RuDjBsUW4y6Hceolq7X0x3B+WKRm6HejmLCcUz9rw2xQMY5kJSTOfCz0ZyY3uT
0UmigzUq+wuXuYI44F7GCNWL8ml0EhMDtATrfg2fsVvnJK9dSCeSfEa9tUDzQmgpU2fFwopXRYjo
gt5u1gDvgzXPTdyRE+5X/fG+whO3CI2lliMKSwg2xMo3WV05t4Neh2U2K1Vfep27YxRXmGSKRn5g
HR14yMwJ8mVwKiEK6ocGtKgv5zCxlTsRaFjunq4gSvugugVZALzKuECxUBn/3Iyyxr25Vqa5Tmnj
f5+SVbJ15kCrU7fxDIb6rb0l+Tsb9POXzfJnU/sSQUWHMaVfQgJhYnlG9oCfpKJ+45zXOe5oo5wk
XVEa6Y0L8rgYcP6aeQCHrCI0+7p/2cDa+TVP3sUFWQsoJ2TJF03qWJQncOJL6QJ84k2BBckl5JXY
11UqBeycBxSWb7Bvwu7WN18eyPL04FbFhhR/7Iu2tjC+aIdZ+rao/U/B/+Ip/d7o5dIDYx8oG1hZ
1CiGrDKUUL1eVtPCrM7j/rjz/XhXIeb2iSc47fsJ+keOnDMIud8YEd6PNdVAieFN/kdvLifXx7qi
L92r5TF7K9cMGw9457hTLX0aAJOlFP+lBpJ76v/of3HBX4neVi5wjtbRT9GVX5uJQgq4LPjtndCG
3FsSEkRuVSylYa7znYISwXoy79S0CXf2JcK7A4eim3YKMVNjC2Jb+kmrFG7b503X8+FD05H82nRE
YClFTY7vujJoBaAZkyup1SujklW6D7TM7rDab9YHtBMj4N7j5IMoadVgrMZW5fF0NboPWAQNwP7O
5KA5N5KeKx/8z2zCFBKZOhFI7A6uSwEJqaR+GMPLq3fjOnOppCioYSeOkEkNYvfqrX/eCI814LqQ
D9AotVYWP8NTYSC6ihjgpgZv/PWVlrLD3U3V7AGq/mpSZMgm/9AliL027wAH1rHsHY0euAqrYXnx
cKrpR3Qsom8SRKtSOM9IZKj50SYD/+IWYQAKmVgUjf8tNZDpZSViEK5WST5ZT6nUgnJty2vBX/gx
kB1XDAzdebeAilbJdSwwzqzKXZ+c1QPBAT4/CiQp72CEyin71vkT/+4++m5umAQgL7cKkTz21gHf
M3nQcfHGFIunveAlv2MKK2qBP4NF6YSKPRNBaPnFo0cQBVwd+O6R1nyR+Qhabe4OwtLjlQsf3v3v
fBYLtVSGhkHWkUMPizjWcKjbqj2jQQ5uX4J93MZ798zCL3xTwpU1zVXol5d9FGqJDHGRNMlCh/Zd
OI7Vz7riHtGwmYr3VzagRvD69S57P3+RWdcTiCx69LgQCYa6DUnL+rPYu/M2cx0PZT5UzK3Z0iA5
XZdcC0Pl3bsGAifLuatmv8N715QCTtlAQH1p/RFKe+mPDnR45lMeTLvQs80/m1gDHxSmI0DHqG0s
Yx2eYTK41Rgb8C8jbjJUvYwc3/kynb9pxNRFaH5k8pYHCOjpCn2j8daYewTyViW6YyYAaaxJjbPI
PsN67hjdvwr94dy2uEn1GOvPPWCJ28mb+as2m13zIYWDfLuHV1ve1rN3HYIpRjgUc8zHxfN3INV/
om7hcRkXpdJtu+0CzHPrFw0FIMC6fJ21iYFyyq/TqVAG0YYQeoUof2GQdXVT2m39X0MAY+IOUcAA
e2S1mkrU/AtFlwJbX8DHzYmkzxUHD36X6Eqq3wKvPdE6ZDO0PVOK6slOXl3F7asje6POxzA4bIiT
lTOldx4xMcULD/FXRWccWLfczE6BBMI05wcnO3hGGHt+YLkYQzPrAAVcwiSxTVQx0Vpo5mK2iWZP
wZP7FWXN3+nDFct23ZmdTogl4eSzzrW1aMSN39VDR5J4HTijon0P2DjyMcSPyYHMhswOFb5J1d1P
svrVq6qpzw7jxSYYHSNvaTEFW0lxOKYZpinUPHOcPk/aEm3lczDZ0SWp3yFOLqZJ4Cf3l6M7aO9x
5zs9AuIJ4fIY9nONxx+8w0HyTGWWxa73q5+RKXJtItac7P0M0RVTsSZnNDKG4FgtzMcGecAtAPea
nBaEWxGjOm2nhs0cL+Z0kvGakPFLra7vLlhlMsiVCVsX4Vbzzmb4cXe03CpjBz1mLQoTlH2dfCB5
yyM2fgWxPu+BCmhvZKE7tBgZzV/p3AhitGyzmX31Ol1kH60cAu43BMaNPQsZDzJt8efUSJNhWxp9
s+RHyG/Z/WRZJ9n+QxL4xYsNA1GYMxUsd0S0u/8ZhBGUWtTr7R5D+3km/W+13/Hqyji3oASrlBcL
qfbglshCptUaLAjiOUxXVUs/0VWuBlH7VLSqigBZhnuvTWmFvWPgtKbeQPnol5ThQ70y5qrajb/f
WCLlh8gwNy1xzbmGjG+qUScuvVb3k+ZiX6mgTGJ4028/7jVFTODYwh7IIgPnxZuy7yXCQLsczl/V
TQ6VBgdL/uqbPdDSyJ8z/DImQ0zrFdoqvvrPdIhOeLtobr0wRHhHMKOseOzcEnwyDQcEMGh2BUcB
Q8i+34lmDnVa5zqIuILc+2e3P6Jj0zuSHVOkdx14nj6b+S6WVHjI5epoTkj0k61MvykUeGnGtfR1
wDIFyXGzpHA5u6pZaHppe9ntgo5Ugw9Op97ojCXgXSvXfl7neX5l2RYxznDY8isSc1tFsFbmmKTU
DLlHnbhL7l4oPkQJTrZkBaBhZ0O4wqdjRnavDS93PpyhUIVcq35zc+dQudcnaZL/4qgsI5kyZlMI
xWyYFs/T4TO9DuAWcZfZThz4QQerH0laEMX2F2gj83yfkWfZUoBW6WjXryRT+Sz/+Hziz7XQII/2
W8RH9ULRnw+7ZZ8fF4miS8IwgoJLwC4ifDzHaQUtbt5bUmWY66kLXihMVoV6CrAdcv1WYoFg/5qc
4TDWKYSXUNJTwUBDh/InM811w2DjuNFuBklqtFWf9lX4E9ZnrUMTEobz5ct+x5QQEKOhbxnLMaGG
gKm1JCeQSDknPuzfBZpLi2UZseWBWekfC18j3sKXZmNxODICFfaHbbxnJLCJl/MQ6KCEkM8XwU0c
9cqnrwco0M6AsimfXBis0oW37mM+jocFaBZ6RkICZXjNnecD8b0LF8v49Hc4zWittSw6KwTy3MPb
5e6L6TH5kmyBRB0x/rNuznMa7u8yDRSOLKUQ7Wa3HY32wZqGgKg/Z1PpEhiePwcDedn7H3nDju+a
mboQxPNaq0/gAVbT7+G5IdmRSTWAaqM7Y20n/MhxVT5Kqi/I7EaYB4cJSuBntn/AW+BvzW8hbqaz
hUwqxvwtgH4sCvtj9bVZ7vQY0+buMegG3FI4j6om8XtD8o1VPLKiAHJyFxmAlLe0BFjyCg9dxsgX
XUqbgI2k4+rC5DEpuFTt3W2GDExGGF7oWEgZp55m00Yh4gsQwRi1WuZbAMoX751bROM0bgEvDlBL
ucxQWtLkT8MxrOYKc/kcNQ+GMV9hdFN9kwfSc7FDwbtWmXbfdZ8YnC9dcCYWX3GhBcwejocWVOWX
IFoKfWuR6ijzb85WOXNQ1UEoinXJOtC/NUrIXMjobpJcvJfM7OFBGaGEY1pnyxcf5kFrzrnZrGBY
G6ePAcgFRQzYwdH5AMyOo7nOFrjVY3sbUd26Vj8Sj43uLHDc0a0ednA8US2fnZ4QOn8aorH2/MuZ
6LiHSgc+S3W8xjds57WgTqjOlCY4/y381PtcNtiXLgfArH1LmZTfCQT6rsWrqSjNT5YQEYRA61q2
TgOEAZxlbEkccwQAIv9w9pkRJTiIWW7bznt8b5Ci7Ck/WpzcDzoQ9MXiLUrKqJjEKuf87tMArGVn
JVuHg5EzXm/pIr9XhGoWtasSh7PYwyLaxgdzOpsM+PRAQps78CPrYMB9guwbwmH+Hrarn1Xu1dxi
7TWMCn0CLeFBorys3M9sBx4wt5lXvwISmI/wScylgX1EcgHX5IJ/Fy1jM9cRbk9D2KJoWhc/Fye3
XSGzPX8Gc8iyMK4cr+U9+vfFcbB4bR2MDpwU2OzGr9DGjPpJ7QbJMsAxH7d+y6dbEg/WGq3j5Vq5
aBI8Md9royc+HNCfB0HVbwLmt/fKOHwCXO+Ca44V4RVL88yqycPh+EVmx3hthspV+5iZVwCw3lBJ
+TKKSbXloHHS8+Nhgt+abmg5ETP7QuFtaOinM+H8EC/x/M/6fJNmaPDH2epooTOCmOepRYaY/y+A
IS+DAS0exLfbWZmZbUHziFTerHgBSLLZsBm7258UzI0fO92IQlgHJt5o3hn+4VL77Rk3urdDzsvm
RYsokbmFsgvog7PqACYeHlTU8yml0Fz0KT2UXFJgAweUNzBg/HGIbEYJK0xKYFHyv0a2kRcXYv07
tQf9qZC0Cs1uuCNs9LPJP5bk2s3xFI0emZlKvYKAVGmsIoQKYYWnYJIy5CB1Tn/zPLwAYSMXRmus
TXG03rETzxY7cTrz663pa8ko9xRIDYUnkHCBnvIue3rQL+sVsfK8Smq74xK66ltQJgzi6Rd/HSd/
TRYLkdvtpk3g6OzVCZ1eY7R4Dx1QWPP2wu981GX3q9zEZV/jOAv6RrGJsKaYhdTLFf4KxIKRTuXw
XUV4Lx5kKsCdIrgK4AYyRcqXceVtqfuszthGrYrMBT57MtloZwc8f57EQehdDbO2juaiKrNxl3b7
8eDffK5dcNPJHICXjllKMFWi9HnppQTk9fTOYGgPJ59D3VMIl/37plNgHNqoBOS1GNh0uKNkoznZ
gG4nfh8nePlCs4ku4X15t27SHWampsBikFMDb7psUlrSi4u7ZzYCp7Fhhm4XI3heOwV0Co72DbyW
mNMSEUPzhtpeHeg1oUzpL+irMQVZizMOtHlreNq4ZvWXw0jljQnKfIOnVnAj7RlJKmQN3VqplOkQ
EpcfwKPCjzaebs0aTPhNMk1MwuN/eXyYTCiTmFpZtJ0s3vK8LEkbEUUiMXmVJVFa3xlMjLpzcRVt
njeU0euPHFt7FgF492iZAr1yD94BUKsdIgMZPC2BuIOt726nMpc+PwVgX7hA2EQAtukQt9OPLhYn
nz+NymGdC6LikQ0qlXdQCsdE88ZHNeWnOnAiUSYfFK8l6STbZMHPY7YwYcqbhdCymMvhpxYJrImc
NCZ7E6POHyhpZsOCqvnnhuDI7bCTvC0wBpFg+mO9eBWMMXrGFXhqaH9UcwuopdNz3rcmlcTZUX3H
zzNvAHgZ1u3mTb+fARw693jL6F9fev8sQMbVwfp1EWYV2WvXANYHwQ5OxWEMz8yNWPzapn4oAEQ0
nuBBgepypszyVnNs7pkeoWxhDPATj7zDeu3gmkExq/tzQIhnlKhEfnNJ4klhZrBt7pThBQjOMByx
r6hQH2onQFgHbl+ZPZUuLr/8M9FQe331PgqJLnL1Fe4RxzSM+6P8AKgacfoUIG8hS9NI8cMiPeMy
j2H63YeqZ3DqcaAXLy/e7SI28U9CaYdcIUBJD4ea1hxIa8nT+IIoPhUiZ5+1jBIZOp+Jh7Xts5P5
bohhubEF4xPo/wLMh6Pus3773EZSvxib0eVAbt4VaNvKhdr2qgXNvCzlxjbOxsLm/Ld+oNEw8SzC
Oz7LXPswV8nu46GhtqMbrnfCn0qhE4apjX8/8nD6M0gOXgtko8wbhRUXHclSuTmIiK2wKzn5Mopy
8/PQ/lo9lXG+cG/zBljIYlDyuPB1glK/MPNZFHr4QyeaRULTO6hy93SwkV6W0kuFRGFOG50HCFrN
NnDbAcGYjAOOcPHhmRoN7MXm6hB892oWxCkBJwp5Xl1UKDJMVZZpVYEHDctzYAXN3a2i+M8PNqRU
vu2XmAkkS66pOyGvOkTRaNyzDrSecHUT8UBr3DEqsxhVgxhQ54f3/eyiEPYtS3AwdM0kcYJ2YETc
UM9uaSWxkqY+UPS4nHvJ11M6BechnbLNMzB9pkwA1zAPrYKlm3laHd7DeRsUTL26DLM9XsKqHYV7
DtdMUVCd3iBZrIInK5KZLd+NcqHLA72Zy7X/1RfFqjNVLx+QxFuhyR0Yga5yDuBhZbTSDMJ77VCQ
JpGVt9jHXKDWrUN/XfcW+kgk9MB5D5vUEUdnwWTL34SNy25bgcI9v464cfa0/yrbEjOGCF8kK/Nh
Mqi7S2tDO6afPeVvZKfgsdLKgFCTs22/uX3Kor29CAf5cnVMYvy4lVsAubf13Mw+WOd1vddxU5is
3crsQkdASWuchFcSv3uVI07urBVxnmTAyC2zdKHmYVCth4B3ktLHT1C6+UDZyt6O1NscI1ZxfJeu
uswwmBfnFjB9aDp1F542x64yowhnUkvY2A2UT/jKxyr2J/2s6fEah6SEwG/HVPliXxCfk+PJkAF3
q2zzpY78aNuZix4WjH6pENjM0SOgXF1YubyIisongx4dLelldUBrTlQmHBB77OZtKyByX2Y0M6ZD
iDmGya8Bon27Ca0/seHe2cGerdVQinKGPLilKsTt/kLAcVlxDBXUcopoz/37LymPzN11/JrLkiFN
zZ9H/UKtHJ0L+DMJcXhSQiGsZpruYIZGivg8sX5uTWfmuj/CBPmTRcafMq1Z4EMy8DO/E3HNGfs7
bsrt6Z2kxJenqhjq//hGcYD9mStSmo+fOq1z4E7ofZ6ExZ0AbCa2F9aqjFzf1JP3Y+dDcUtfPD2L
16HPAmxmPLEVVW6K0LeeH+3blT8kQ2V64l4+FzAkxaP4ljK5OmM/nMteqC02E8yfqWYkMJsvivy0
WiOJJjkCGzMKASsJwEqtCAq1OWDXEtqXMpywTN4WHeUpNJcVUvtdjR7cXyWJ8jdQedhgoDjoDfzV
7FrY09Qi5t++5oS7vBW0wc9qR3xQ8MKzOGa7vAGjFg+DqdwXDau+SXLhh8CjoOoBJaxTz3ssLXv2
xz1OMlUKcvorhaW7YeLR6uKxpbWT33fgmjtNas5+NlDhhm09gV6xbncKD7IF9Xxcor+o9yoF17I3
my4VhNOwVV0/pQ/wvzP9Yb1BSwJoDvNscRDH3QH2YweEMFW9lg0UHLb3aQ3TVz6Yhmw/Bgaolu0S
TNtL0JtdIuGxloKlJVLsoW9plArRLCPOJyQQ9eM4xWR7Xy9wmmGPRc0uLhwv7uqPhip0N0zwMEca
/v0Hdy7OjqZ98gqJjl/hqydWaGdxGpQprxC1jZni0MeaCM7hqMLHseZfFRaldmVT4n/sGPiJnJ7N
3fmC+MPz5G/xdgMR1Dd9iVyjCZJJ29znFElz6Zicq7TfE5FUl+kaHgEyIzn4ILEBPMucZ335hFr4
bcHDZphG9vMnzXkJZLERcSMZvTi34fQiBRFTV8yuE00hzI4J6vqDrXQ5FWfMxUY1SQhy6jm3e20C
UBKPljaphZr782Qf8xAcVPtUYUxLdPH4Tyw4ZEMB5+ZFQfJ15P0k9F/emKWA1LNH7YxTJUt/VhXH
50chIfLwi/PUJcrf3mvEyEASC1pJItzM/N51NQkT7mq+bY6goRZiwUFfhp8hVpKkjmGQ12UibfA4
gzfCC7dQWalbLxg59dmlAAk6/iRSinwzHIyNaVGo52OYk78N7abXAwOUa8N1j7QaGRtUK9ipvwWB
BSqpcVdEThRU7/beQgpBVnTsOdlBbEzhJ4+BD9QxahXXXJtd69M/vpVNnoY6bE43kbj/8jMMTARl
wGv0IWUQs9Lr1bgAevK/43by0Oj2Ma8EiPEr4Oc2L3GDajjh5a8gYjRAMwRmTPw9QcVCgkirQXHL
s1800wioRxeN34EQZmIZjr0+TjcQ8TpIOts4ISe03HU5Jb0XeqwfekRWCBU2HoAC/geFkHFJx3Sn
0MjLNp5hlbskMpXgQeJHBfi1GHXRDe1g1eJqHZrtIQL4eST5fFQrhsx0vOaMavWUvgOorSO/TEm8
aId5xMLgF8H9cKzE8mEJoA6f8qde5oypv0K4YEPEAqHJO6Oq3rJBugNFNV+PepViDj8yU9Vs8HHE
IWTjC/2CzW9oVIY/lkwbbwcke5jH1m/GPn3HaDW7NoVI9bk/PpRvE8VBcH95+SyqN8YBBP3Iy1gA
hzzhNgzS01zCvoL3XbrkRe/uRykIW8UaqflBnaN5U4rg0YikGhcK62dahkp+bar9yf3iGgQCOLAd
VfdVoz3IGqLrsFU5xw7N8Ta8eoFoKDwOFV7CmCgittWAwJFotsDoLazOehfeIHDKa6hw1P2eQTKn
pte+e0iyD8+BLrQvFjJez0oGUrHgYi/PDw0RXd7bd5+gXdB0lvTFzeUlzifxBVyAzkagefUEnDeo
yiPb4i0it+1G0uJvpLRXpB26ux7GGbqXVi1VdLqAAS5XtpfVQqhoBdDQJjJsTbEzov6AH15+Lj6d
W1HhtgEARWn41/DiOM+z71tzHGy0D2S0Tp+e3xVkPeXMj5SHMpx8ZpJhJSkCJkOOCTTE21UrWiy4
a2POYkxwblJHYI59basc+ws552u2gVxG6omRexTdNQ4BJRwD/9vZrSgRpcMcJwl2byc7AW72+YnH
wvY5EA1grg8Yu+p/xbEr1cA+hNwNbQD3pI+rvI9j317ctso7qt3bSjBWtRPvOKUadTHqeEE6Aze5
feC6qKjmIETzHugi9RENmjlUBEEVhvJ5O8Lipqo4Co0rhyFQwXJAQ8qj+ajKsxJ2YS+LvQonIuzu
LZiLaQ5I2tWqkbnPalRAQLpkiRtpZRKmwvwU2lXhE1svCapd4inxExU1xosgp5YzzFCz9nU+IW1I
/aJtiN9qb4H1zrkZcFxIPcSqVdZ2DwU0cFA4sfmQdqmODzAAUFczn2FarIfv/I0IqYiAXQy8KM90
8bLZaOHRui/x14m+s69Jy6Nfw24zQHUzqQpnMOabI0LoWk4mvIlLO/H6FPBqfehTn6swgZ83iRJs
MOsM+5CdjES0fJRQZqZ0DLbABXd9DTsXhcdspuW6+V+wv1CsPLjHHYkUT86lPDIFqlUVMiN5Y9eg
Kq+1CFmwv9ZcI6HncsH8v4mD3rwf8LGzKU7MHheW4qUHQ71JWnSr80Hy3uV35s1vuFckcRujwQ2W
A9rZwbsxpBTvULi4aV3L4RpX81P/3yiifAgF8f8UtJ79ridSuFUFMrGAK6I2mCZwpmke9NZ5zWC4
a5rZfezdeiw6CU25PBAZ18Y25sLS71bnmEfZXczo1+oIhtu0fYGo/sNsOE2txbI62RRHrbq98LLh
+QtYv4ATlgR9jRkGQ9uTr3rxAYWSq8PmA9+6oCCwoxZbV6aiUaDCTW06JT8hJ+BsrITKG3vVadb8
i7sZYsmTT41vCEztK+Qaz0x63c3AaK/vwm82Z5sMg2SXJS2+B4qblHUseAfqa1qXQrahQLnhIWdX
l1gO8vfZmLuzaW71SbbotOm91MOMRgzloZsId2z9MM0PBBDIDJ+3JKr+bkhGRctvMBz/bcsoVDE4
3Ax3jldIk2w6OWz6kcs+c0H0Tsk3yARjFAzYiGDH8RPk9qFKLMqmCPULE+q3F+OkJT0TXHyXD9I6
i0q6Lr8gTe2uVsSFkYG/uOspM4i+2sIJ3VMTzNqRUf8rOqwIYdZmyBEauuso3hZH+s31uSzJSzBU
gECFHmUW90Xu4RS2ZJNxZMIvIYLC+DMyibRuCfWYjsYcZLCF+0GeXZLKCh+GGzuDNltMA+7d7c94
kywjkHeW6XyuvGfrnh9lsLUg0KqdogWBorsGzM1Km+8Ktxj337/3lNTHHE8Lnbxwqql/f0Y9615n
Dvj/RvyRD7eQKz15fPRDNc+2qJzcpw7Bt1FkwK4vyhZNfMSYic/fRz7tDaz0xUvNAfJkBk1Y7UKK
y9Abo07k4HiT6UxrqaANLgRwK7agSd01p7fw1At2Ljbh2JjlQt/lvoINV5aEXyw58dRNOYgtZ5or
wMdl1c3GXycWNbzCIYP/gxapqjxktD8WDM/2tNeHOYlRK7TDa+k3QVtUFmZnniy4lXojNU6AdP4/
NeDPPPUQhDCpsB5Gyk9YX7Qjkrj4is6WTgr0QOXAt8QPznhASKuSOSGbNhSqJerEnTbyJcee3IW1
Ta5KXjxl8Itep+uWb4829uzCv45mmZ7l2PkrzgBaps52MLnqr/LZre7OM2TItT8WRwiQPBLpv5/I
MxDHy39/fqyf2liqleOPvFqg8k0LXI2asVBAEZzEct/ABJ0v3/a8Nj2ns8bB0AlBpixYZcOPU6Bd
0+iyYqRfEvkomwDGJy7FlKVOLWsrS6dOesCaI+0dz5fFk7XEXRSGsVRKW2uznA+vp9MxaF/Y1OHk
tuMwooQLIUvHzSVyqC2g3XGJdi5c2RUNLxuZX5Ivysx17bfNXTPykrMwPv5K3xTNW7Q1VMxms5KU
i9bkTv7VR7FzNeZ0NvEY/mCr5WkFfLzBXTiVmNInEDBL9QCMpsXOctzxOUUALu+mEYgA733zbmP2
v1/r96lSstdvE91gqus2iaW+N1iTnYQcRzyi+6TLbnw2pA4DXsyPK5j+NLYEZc0/Loqyjt8v5VfX
nEBCvnbtAhNF3YKGhrKKpmDqrnvJiwkdwNfA0pZEGwGv+y6k2EV1lKZU41vFbvTLpYHZ4Jsh2jj5
t/X0YZcRcNTBo/3Rf0ubk9eW8ULB/uQikJ3mdXBrfm/Ns3j1OxUYznZg3k80AwtBx8kvsgjNGDfn
zdjlRI6JITf3YbdVoLhmZEocQ622RAx2YsGgg5YAiU7as7q4CH7CcY2AgOzoD3uQEhJB9m0Gvg+O
kNLqcuv4IcA6g1psdRCm2VDz5WCk7STDIuH/ZFR8jL2+nxagZDCCrfVBsm8jJGI7odyfezgszEYB
Uu92yXUw4O/9Or7msYFPtEH4VgboPEdpFDo0fUXOUPqD3LzHL40oPNSE59emPhmD/rePP5wT77ui
GAZhDoWGeAMG+UJ8yXijs8ajBjM3jAHunRwTpNMs7CJ4STgpmSLd36mN5BPJL6/fI03y1iSXxAtM
PZ+rjynq3zIIO70p2e2TsShGTGdC/l8nbgRL0CTThtbAW7cOs/ZlxW8CeHTnhwIHmSYCiFwB5icg
90y/8ARmwmXABnD/yhGM1OQ2WZwtX/WVlepEUdJciGCiRk7GiyaJUDYozP0FXp+DbfBjmvexql2i
Ev/Or/dbYTfj5S4+eHRVSMIXii4fnzBbHQOaV8zvdYg5SdIAE7Sm4H7vYgtHi5epldQBNTvfvNa7
TtH7KO0sTH/Q83Lnncs/tMPVpBk2keGK7TnDn9/+esAn5j7M9iiUTdUx3AmS2The2Coh0dNZbiVI
GepQxF/FlTdGjFvvmY/wH6XH6GYUbWXZf9zyPFDdFV8gttTPDhJnEfIRymQ2e9ZHRaT99hMuhYa7
6gspqrmt4x8oJEypoTkrsc2MV4jYNIN8QUDNMHSKaGyKq+J/7ifL3phkAUSlNqC0pdDzO9DCTRUv
5ry6W+EDMQS5EVdGESR2Svqyrl9A+qM8TuBTa0/oR9kQYSMFKshalqQWA4GZcHwmOgq68isG8KvW
VZkuGwSxqk5QTUEyNRloW8oCg5oSwjat//RdXEQHGmvwiqnLpSOHSDhSq1+1HoFz1KIiJAMxdv8V
ZcW+9LczyOwDsMKEy2jXE5vQIa1Mbof5N2dL9cQ2f49gdMbW+1kQyAi/e3kFf6n4MJg6vmeIpHjn
7bQ11pG3axYsJoMaHCji24e8iHFbsfswe+94R9aIQhEq0yxmGDWSvJ5sloaNRSySDsrOXVMGWBXO
/UN1yI71xr1B8TnHh5ecRv3FaWJjZmXsNMqvXo/4Op89ItoZ0nt1E/9ScOSZZ1FkxM9jhZbOckBS
yLkzv2+Y/I8aoLJYhBMeCQA1hDeGNLJQVodRonPf51r/e85GEw5a80REdrVl7be32KXaXoTReQAU
eBhCbbozh6cEBf/nWOJip9YZm0i+NxhvdzUJfrDYXDNOw9SSVHWhpoMEGz8rdYJJcgYPCaijextF
cGUaJwwzuh83lB04qQGFSwZ5QPtzo1LdvO7JVK4w7nd19VhnRoX+uZuCpT0/r9EqB611RRC6WwMC
53r6ufKvZp/M/Gfsx29BuKR1Z9piYF96/7eK+dz+BXX7q7CttaSFqah98TAybFgvJkwnfq5U3YuE
PBUZN/zq2Q1t/qxtn4nKrh+Zt4a4YOoCCOfCDXpuMVQMWjK/Iw9IS2T+zc2hBiYCR+u4Wuykb0Tx
IADz+yA5FG7FcFG1L89f2GN3pC90RS3CkX1QKegXXLX7Spm2vpO/8GGmFkgRunvpCGJkbtI8DxNp
WxWEmR69c7K7s9z8SJiLwznJsljbWYWJFBRtsi5P0i/gW2jVD0nn4zUdMoZeNp4ibOnWNlRib4hq
4DutCAWigIu3BUhSl0oQcQYE5F+eMLJT/d24/DpGusbiUY+ZSxSqnkb9jEGHpryTOV7QHl27sFzE
gEiJqyOM7HI0ODvpb+P7uNSTCVTx0n1jWFih7q3JW30PXZ08bK6F4vQPijshn9BcISqOGUYdeZiD
EblirrLlJL55Ijxbel9xvxCC+fvXwMPvM4MZ8vbbSSd3Sw3I+c6G46BRPRpax8Y1oHInVwT/l1OW
vHCozWjjKu9sBYX5/JD21F10HczJd0qW9UKfrt2fD/Q85IYTxhl3uKCuxz+k0BOfE0Gpz6SGXsJd
zCoBM60EEC6SLwWHSDYPHJglftHHfsmLHE1U1zLKl4G+4KRvetq7vLb4PX01MNkYdvy2AQw9aeuD
uY0CQhAPl7ysV8Fc0fxRNT/wT/VV304q8tx0w32SuwbqxtKde8upPN/9+cOnV6sHpKlwL9lCHPWC
9xHRnh9zsWTDsXNwheecOQArUPgvxU/Vz4uTDgs/jhxxALTve7EPeRHE+h9Srn/ofcmmWcmKeoCU
2QLVt2MQo5E9/kgCtV5oXTwgEv0qdPHKJde4EeaSGkCyRvl01yqkHMINH1LvVF4+3Np99/nvRDKm
cUz9lbn6pMEZ5gN/8wIjZchXQrcoIYm3rUp8GivuifhsbqutfjoBA0dP+e+NdU0ccIw3YBfsmExL
DY4e+5b17GcRL51Rj5o93rmufOAYW/l1Tgc9b8YQa5kqRC2E4cYcb4HCmPNFlk9mFnYjRMCDaQUY
ztFu9TpTWSp7TI2Hf2AFKebWeiDnW0+WzKdPEL9NLpL6hS2SbpH6Ou06NLxhIu8sWR6CZth9ojBD
LLwLq6tle33fqxMJkGIWekZR63uLVh/7Z4pTho/xEoLHUrZkhSIc/KITkBa949+8WA/rrSbMNzWs
KeqBKule5+NYn926rFIpViGoIfA6AtDZVj6v1WvRFe14ci4tuYKlu3CaHJfZrj0hZWAA6an/pjMz
uEVwPkl9rNHcAuHiUBHQcJ3U1rJ6OjxFxOcGrzP/tx9awdJJmKi/gRc9GfzucWPWDO2h3GJMBqg9
hJ3JXwtoPOyRysGlMZImznTXR1RPVJ7Zyrikp3J3l7m80W25827gulu8CpEuj+bcsHhnusxMH5l/
3fDMbqcyE6JOSLm+mis0U0VOv2Xbf55QBgjKN+AkyXNAuG0JDNv1+3rtCIEM4twr/qPDZH8eVKzH
1qhQmkbyafkUzadBFleGOpPfF4mMcAd6iR8sHcbQErapIYi9NuVPzHQJ0rNubFoulZU+LCkfMjGc
wW/Y0WoaklCyv40KA0gIULZFqMWVqCvJ5a+Brgd2f39/DBeQ5xNWRgfo6d/25Jtl1gpmz4GBUmRd
vS8+Z3WZmnEHeJJ2+EQSeOSNTPWmeDU0WChAz5orUEL5cYruyAufMAAHGUOJ2WnfCarrkqMk8rnO
0vwP/rb3MBhb/fF096jiQhLA/MRekm8jgOzaDCVIZ2+L+68dAAt+0QAvcQPiYOC+k0LMvz7IxpSx
QKhwKdGBEVL8SzBs1hKPRHUVh+afbMIFPY5Gzaep4QnSVRsYVp6Z23LWHtYY7MvI/7mezm7nW/x3
0hThT8RcqDNBaZfaRikuUaai9/+jgmHXM9tVxKeGpu9pKRNK/V0kJGdMzew1o0cq/TwGjHeeRFF1
qVWNxvaQIaWlDI8teHwypSp6T6Fu/qWjs9N55I4FG5U4c66+56ZswJnfJ3cxBX2wlPXiVoL5N8Nk
9exn2bEpaL/9mXYxvvRzgORaGD/CnPAK3O8T3LAqYH0BBPGU2q8DnQkbb0+HUremyRpk7+/bRVno
f5U3b4dEZggFy2KdXZ40UlX/JWMIPGyfcqjYXdYK1hZNxaArNEowMPMpStuvlQ+hV/uXnKpCBQ6c
p3H7gLKQupXfd8+8sa6SJ5Qm/qA9TZUC8C47aJesYtFGHE0huzD/Yq+99Z43kIfJLT1T6dMd9E87
WUnYGB+Asjg3ho+yaHwtnpIF/B1O8eCHlBCPf5apB8n5DKyEDWDIPSxKCLtUuJ8gas1bUqd5l1Q1
h1DkVDOzTfDo7VymyMUhlhzQtqY0b9nipJV0w6eNDn+fnsNrJp6WMLoFnOkC6N7c22aa0M0cMVDB
nVv05WTQyMjns+0dqNPZ/bF422y4XkLHkUpJssJiCB+AORHJnTC48BU20arJznspqsOvM8ZSzwmx
gzd+zpLtjuQgKsremx3W5BFflP5wPnLnrlsDCCJHt80OfeBkuHNvxuAqg1agC9C0MfvlC9RPLsME
nV2hObaJoF/fXksuLf+kDx4aNhjTFw+PkgqcPaZj6DMgVy/q1Tgqb1+FQbPRJka3Z0BH3oOXNt99
1Z9xrgc2HKgdMY7bNON//epesQ+vlAi2OVuJrGpDdOX9I8xMWEv5ZB+g94MTTlhl6Yauop9Wmuv6
ulV0xiSqZul7zaYMUfmgbNuITyQRqKq0s8usNCyOzf4tPnXxHRpnig9E5WDzNFM+PbRBl7/zDxc1
RFFmWXE/z7MohC92PZfW4KIW1lFZ9rOlGHr0gojEWu6HhquUo1d3be+C+TexSIGbnD6Bhv3XZDXU
fSnhf6xS+En/fY4QXFyGbpWEesPEJgo8kOr0HZL4kxD8jSWdNUdhPagcF0/oPwEL+dlSUjt/j6PJ
yv9XG6fIl3hgVuN+1mGytkw9HkqKdrApyG6CILLl0iVe4PDHLpo0kni9wLPJleQiIO8ds7E72edr
bmJbfA4bsyFkHxxJHI35Yx033C7agOIlXuT1wO/ks7rCHpSRgNUuDYs2DvJv3EUUOIUS73B6D35B
18WaFuPwmk4fwQgBNzDDkGhvuat2ITEJfTOGcPbBdSh9rUqJ6hQ0bMN2NYlV40TlV/SzxnHv1KZ4
4X5L5DkZ0iifLCB4W4IkpA7GDr/PQHTQ7ZAR2E7vVNsVEF6IWpcvrxVkxVii9dJvCuE+zZeavBnV
aknnon9qgvf6vwNMRCZnFWoCMCZBzbaS8u+21S6W9zHBUrxnTpCIQk5u6d0mk7HHWQM+nIN13u95
wa7oYv2K1lZ2gB0PqHuGdc68t1QlxawIa3tDVPDmNriFHLQdwUFqDQzx2we6f1CmfZIVwJQ1sh8v
O0elAegdnJxul3HUrg0nNc6u2iS3i3AJ7jjU6bzMhyd5AvsgFlzolTaS3Z9wIIXbHrLe7jUkNe58
2NC8NZbHS/I7XQUiOWdtB8zvCXgWlPH/v7qflpQ3bkyLrJKcplCsrfGkuMOUoPsxuyZY6WnMZeB5
GVSxLmJ9oB84mDphModtD+CdB2ZrhKKZ7pd7GCVzypmebI6WzgHglXLXN5d0jmkPBsI0Y2zqkrSX
tFydYykmvjCcUjNcih+kwRGPvX8SK2XtkYW3np3sTdbMJb4Rgpx00NcyC18nny9LTNjfsM2jmipM
ywEHKIrVsuiC4ML5xoWcrWLJOYwtSGbki9PanES1RtjnfDa60oWGkvREAjHhDpLQ48m+S/r3zy2X
Ti6hSfOW28d3YF70XuWv1vqovbWOhE5ZttqW+mpn1l7ucGsyBK4ztjCiid8qRJcO8ICnvv8GxoK0
XieN0hYfoxEvtDEsaGuYhy+IkSBfn5t1JeEvvFipFwMU0hypMly0bX6gPyVXwM3OBTP3WAI0yWY9
J7XNBLX6LKtj95euv9/H4XCV09BSO78Pgg8fTE2IhvGdx7s6hrMy3BXep35YpBC337Xn5g5Tdspb
VrtoyPBHQCGKeF4GhAbpkKSAAOsOJTQ3OMDDEzbAvJMtV9y157LXzkoWNujVzlCWXduaahFK4GXX
VWhQHAuDxcU1RaIQAGSCUj8CuPgqgKJ/FCpe63YDYOohvP3CHiAHz0pAxNSQmHC2oNGc3B1eVL4s
pNamIasRXC4EGs0itBuOcnrDUGCzY3L46haD126XbQR9m7ju0m4YtRlhMMU5md1TM05F5eCoU54U
Pk5HOh/XfOw/+/bq0DX0ZkhlKP8fIdoDKWGeelMpUGvIRx0RSgQieBLiM1V+9PTpTs2anPXWHQ0H
Ibow+tryZzzZYm4DCk8y50CNvTwzOHNAUIhMBSAT5QJeqW63S0o8weqR35/e/VZw/5tV/E1Mu591
kFLsjZFhAV7BwXKak/CSM03Vn2ilxkkOvVlPOcgwHDr20thNYuyVUCmMQbckMOVV6SmvkaW/YjOs
ViHHUsfSTymmZSExahAaLZxHgNb4R/VzZ745MemHIv3gA2dm0B+eucMKqK+3oeEu/gp0WOOc9/8C
4mD9TY0T3t337G2l7WeVb133kfNKlNIZs7hUGYiIORLMpH8VzkuQKxiQajYZQFWboH9oWf+nfJZF
x81lilONbi/ae2NAVyspQIPeYKUVehMJpCMlvVBCDdqTVvHbMxiijxW/nLhT6S3K9zm+tx5qoqYH
XJv9EBZdk5+B+eA/a5FvoEHljR+2WIRwPc+n1FhZgCi0dqDWlE7CT0oX/AkATL1XCfrbu4mo3e3U
kS7eMm1AQyqUll1Pwl0Jee6tf4S7VL/8j53UpcdG79aP3N2FsyqTQn7dgU3qzdFk/uoMFpnkMpwx
vtETPbPB2MIY3kEzLxpcTOVuDkfDyGzrDwWQfF5iwkHDEG+ZogxqpQxqml8kHH1m1smdbDAwdUXo
RpSsvG2idwQ+P5gXlELMqYnuNs39uxHh8ME5Q4/Yulj0p8FgUqJGQnfwxm/nV6pd7ihiy1uo97YY
euEQATHYMnbJQnyrFV5Jm2JUAF7zpqQBsGR9WuXkNl45e4rqriES64BlGWzOUthAKgcaSiVG1dNC
SKcEN+PERhLqypc7qnV0bOwHygBemuP1iCHXluk6Mq4kRcHpkngGwG0/ES9RzUZGXJs1ipLUe1sg
tm1Ha3Y6SuSIW2FueHsDBq2uZes1de7gpcOsQE0mwOpBX/Gw69/4Jv6rQ95oy2SC5dC5ifWdaelG
LW10MAsjqAgtxPihymrFT/SlmEYsTDwc3dIPzEoxSmERLw9mpBSaIk0Wxoi16g4D3DqMjz8VwHyI
MMA+bg4tJPYep9iN0/51mhRzkbre3U1i7hkuMa0jpnGLNbebZRTrOYYww8MrbiSn3rSFebtwxK31
A/DOJfYPQopNHdYuqWQTCxFfL//Z30rZ84f+p4f7qJvGbziRtyDAZ9RWW0ezaCAd+PMLNUxfmSS1
M8TPhdbKmCuAxAjCWggAiOuoshQDboutYAkWmJItgF65P5vgxb+HjhptD6mL6pfiV/z8oFVVqR6W
k96x6ioUqxoEMaywdhqy3KHcp6kSQqstQNzghr9KEKB+5iFmhk+vhz9juXsI6PXP3mA4KOrJvhac
tiHcrp3Q4O4KS2k+PH5WGrlWzhI2YEzywYBOjCGW/aVYavkRTm0SexyKi24RJNY9+hFAf8+HKMse
vDNCKOa/d5Vz3vnorGoZxkt6fy/NsLXu7dJCXG+V5JXEgJsKY8588G0ZP9vuG4aqzZlXeirXT+RZ
DX/J+v/nY3hLjJjOprApYTZtN+/h28JCS0Chm0EyN5DfD5a5PnjwEUmFVkG9WPR86MwiJ2aVt6f1
MHY6hCZiVI4EPBL+De/Qk4Hva//LkYlCnMhuk9/RyYfv+Q3Jb3+wjQuL90AJr8y2HDy4P5wDyl/t
3fhqHcyYDZ/9MLany6SWD3JEtN6HZ9dQ70U8yGKUwitw4KZAry03eTr+uQlITgsqnRtmAf4G8BrG
cykrSQePKVkiys7M03xH64dcXr6aeuIYc+OM4FAlpQ49QFlXmD2JvkdOFEp5qwyUG0kHjPBhUxHL
OtebqU0TOYZeRWQUqiNP9sPaSLZK+/wuTyryQemv1I9k6hnFEVHEGT/tM3TXUhT0yAZ7iF5OKUfm
58UOVRCOjrQVfXCpcxuVC7zFpTLXpnS8w2OmSLYrzjA6ji8grRtGOP3Y4slVUduPxmIO/3VaRFIV
kfwn75YbaZixxPC0D1AKOAdXjrgJ8MzlCj/DcrcmaF2FTx3HQMtfjlHcg7vwuR0rwH7rGDZD9VUz
BKCyIWlZMftPXyo6JB9y+2rL/AOwAvjByo40xDiLv4kfbn5ir1no8r/Nm50MXPI22JZLqPVaxZ4Z
ezL6pHSx7mqQ6flf3IlgfriY8GGq0jibBAMuST+6sHJA6dGtand0iLpNHuIO8grmyU8RsClQdNiu
hrj0ZxshSE3NaN22xAV1KhagbW9vc2o2s47hx1rCHGiarVwro5I4AKndGz+Wsuc35KFjZOBQsNOm
IKuuQ0u2Ig94Bgm6GzD6bEgVqnMnxV6reyNp4pi/nNXxlWFud+A88X+93DGfbUCUHDB6oBhA5eG3
HhGzGX6V0StFBvuxg4D7lwIpGXyv2V1+NJTiFLW69UHQhUZBznk6x+EsFwILl5EU9rUQ4cs9sh2t
Jps01P/vXFjVqx1XxHjruYJ0YWNlUi01BitkqD6QxOR+Hg5NdUcR4RAB/SmrkfXC85xvj8nGseR/
g4/NELIhKUXNDn3BBYptkGgPICS6UG1aF8nCkVYRmDDmkVcZ8LSejCqcirPGfiNtLjSTFC/9YOCQ
xMWNVbHunZ4oieDx0q5DXmKhPur51OlzuV/a9Tn8319rdoayVAjkyGrfMzO/G2HW0N6jfTXO7hF1
ecLgYdDfA8dO5RGQbMk1REPOWpEwCl5dX/ne7ZIbV0GpTooMBye8WAWPp5nM0lIYLIy4EHnh8dAI
Hseho939I1O2xkTXli9iZkX+ZiDF46U4aluGMkatwMjHi8rwhbVgVy6JZAGO9mSVmjNd/1TVorp0
LVwor7BVYsNWKPOHvvrOZfTysWklHPebme0wxCP8gopJRscUl2FdR0iG2lV0hwtSLnW8+4N4GlBr
KQcjVzVNzqgSCIpuXDE9VEe00w8eTPzQCehX+TCLQ5fsTgb+QSjve0AFNitUFYAPRk5Vp9ThBKfW
tvUzEbOk6m5e30ouyyKCbuHMD0v5AJGBALek5y6C8KnBZgvCKv9I7sKDjqY9RQbX2af3vLRboi7f
1tjqZ2VjASpFrltTxrZcDw0mPlqUtJpJtBRvpk5cBH1le0Os0eLd46PJIBJZNfwGFljfWZIgAwYf
whJg3XuXh9hUymwBx1TO/fQUzOrpT34Ci69UCBW3TsvsOWZdFyF18sdJCsvKOMHx5nc/4ycSM5Ql
CeBaK9tQtgMMCBtSHsbf+XVYBShopvI7tS8DTBbB//n2E7OTQcnLCPHSaNz6SixrnVLzK8xk593H
YA1ErveAckvSc6PvL7GkHU7MFTW5PipBhNIPeqEWAUUgYOhCql8k7CWY/ON4STENOP2DzmEEA+h8
zu+R8846qJEbP8A9y6fJ74Lc0yERdtEQDv7phJwFJi534BrH91BuLytqrckd+e0wHuv79oOP8JF9
BwA6XHUxAUrGs3nXmzKNeG/fku94fITz7LiA+de5G3+OOg08yqnXTSgsVvBOHt344fu5KiDnu+dE
TCNruYvQno/lXMTGJySgI+SCeZbKBsWu85+1OofHDNwPUImx8Gz5wHzRlEZlmncANppD2N8/ohTp
lNbV4bHSo5s8Vo9cg16LMPn4Qi8K4qD55E25wdcdYNZCRP4IbBXkCHXKAw6Qycflbek/9hvJK2TU
foK7kxQC8ntgiKsP0HQCw3lbB/HOMg3pHMiwV7m5vALRqdGZZc31ESJ1h52//Az5JnqhgNCaG9/0
1HPB1nFhXf8AuZ4Ya1/3dhkZShiZ5yUT4SlzIvWgRpqUNQks8wjE23T1pDcmCV2/bT6kEPsXUZU9
BWLetveT8/4SpdVs1RU02Zn+XfOP0bB5KUhHrTkos76r98/gGdSuVQIvH06M0fCml8U1Ee9yjmzS
o1MxULCsLFHhKcCJFA6V/PlSjaTtED6dBCj4Jt+m4ltZI4u16dZppQ8NR+Bl5urcmvUVMSxXBa8N
HU37+ZABEw9EPhWmT9iVYrI0R31831fZGTrEsPs3otNPyxrLQ56KyulGw36gfzLtAIWRn5L7haTD
ZUO+saVTeWEIi85YK2yH//Ik1T8wMYFz9BJPDdPXrZENk+VJ4PcGfPlxeB8Mv5JzG0je6VlFl3l3
J3VDChbkv2VZX+2864RDuchm0lwawWHN5AihJ3P/IGnqzYBJF6J6jUlNIYKahvBqsXuxt4pV6VE8
Sg+wiqycyxS945oKFh+efmHzLscb+a8zMsKnGupgq5aSzHu9wIxSJPtwNLk3yVsyqgtL3/DX9eH5
iYUSClvOaGrAyYnfK0dI0Gj9v1BX0enGQ2+1jTNQFBcLdZO9pEad6BqAqaGLkbkOgvORD3EVMwWy
xX/APgfGcZXAhTU+15qXSiRu9UvBh08IFGqTShYC9b51p+h/14W0cDs1rtYXRjZDI5ySwyTww82o
ElqDtv2kgnhvsbz9KikPWRwDMWYn6xDNoiyjzo6kAFfc0vpxPZtQO/bJUeGGaWrVx/6j35FneNTj
A9U6eT0EL/mLAkM/Hf9iBu8J7DK6CIzsdwPvg0mnV7Xfs7ArypS5DTLHEDb/taZ1e9pG3pEi6CKy
i6m9QS4ZeCMzUfX3+B+/34g+WKuudkpw+exKqZiQA2kV5qCoZAyNZwXVfXPLrKPfwigsod3K9eU0
TYw+PlcZQplOKD1JszR5POP7ZbwLZ6fXu/jXs3WhvNNd5Gs++HwFjRdR3gnwAF//9SicXygivgmQ
Jc1rdW2ciDIM7UvsuBdx2cDrARz8whJcDsYCf+65+bsQw7w2rRSJv0qv2MryngxMMIysqO2tuvoR
NX8S4W/fbKbBetExno45ybgiaByu7Bs9KwuDfZfm4G6ehtMPXTdivRsplxYutCy2gxDcn3jg1Zc6
54JaQryVvfukKOKtlG1qfYh4OUHp9lypy5V6xCUEQSctuesVisYpAW0ilodnUopxwDgN1g==
`protect end_protected
