`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
S3c2Fp6L4+SHN/7T/I97dSAu0iq4i/nrJjJxWv5pq+q1JExi8JOTLdPmGPeIBbD/UxX8JpIuS4vL
tjtRNCHi/xyM1VzwCIW6vAJyVmnuCoI5Pk448T4iIhbAmc0i2O8/LjkurNW3wEK6kfv+CaMmwzUH
LBEEWtb2SNnV1pzOsORT4ocM61duO4OsZN24x4bpfR7aL5iXCZwJBCuIt4Hynq72U6BCzxc94mhh
Heh8RUPKqMrZCWaI2cHDkVpNbi5r3WwgqRzWnb5kkkSXncYO4JqMLBnDR1kuBj6/WtW38AdrrzkA
hNvRyaaD9D4N8DAK8zRu+vMv6Rdln7ePB+b5eQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="sY7Uobb6tD0LasDxmDkX4h/uBxNFfDbHuXOXqfooCJ8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8624)
`protect data_block
5pF5MV30OYZpJKn7BLZpzHzgOiVfdqh0rIEb+YW+ICPToTwnPkTvqg+szxyTeVdoUkuYov5XsDT5
/nl+rCSKyFb9r1nesWwEjYcH60I4LXyX0Z/0XS/x0B7xZXBGZQlD+HwLGLzTJfcOe1MQwXgrBeoQ
BfjYj5Z9Ltr3g+j8teYTf4L6CyTW1hjWYtE23KBvAjkz6yOj1b+mc9Xy2sBJirP/J663hAbRleKp
yobvTwhg5wVqM6yKDZ0NzhanL9gk/8C8wPNRWRUkomLbiaj3AGFy0tXAPe6oJFsLHpdWJPWoPuol
MCwwm0uhhGo5dBlethTvSl2wMVr1fAQ1AVP245AwTI4J0vFWx++xKYrPajy7jj6xyWZJEbXBxDkN
IzULFhNU2vl5H3JdyWNvPDlRmvOsMlt6kSVu5lSbWRIL+FoRfGCRXoBjBQmSD0zFZwKL7DHD/n7c
UwhCCWjI57WoAz2D66jvWjtBNf2fySZ2yFTSEAz4XpDfTuatPqqUAYVIVcAyY0d9YfLHZNWtpPz4
zGrvyIXk3fcFLCyiRMyGYZWn+6ukuj3Js0Qx7XMPXqzLcbYn25dX1SgmZIKUjcMBbHfx6QXphiES
9PHGmIj+j84j9jOVsl5Rx/umjCwlMt4AYua8c4CqDHyAbXDXH69TjFoKzwd8G0Aq1sprzCwarkoA
vhs0EAUzZYleXRepo3N3a2HO/gZUBjAPMnTfEmFXX+RyGoFnK9aTStqLXYpWmUU/aYWhXm94f5iC
ko61eI696Z5M/WjOliKgjvr0qgP7Kv0xyaTjmBPEp8/nfn4vNy9jmfPJ89hnVmv9XV6+vuwTeQJH
98l2lJGKR3f8jjUO+99bO4v2yaqHQ/njM4ESRN+7ks4SqdaCFOTXzXXtRm+49PomvP7PluIVonG+
rnmem678PyZ7HZyz8zIhEmh529YDFKSP51+XK8CpikpOP9tsR48RpQ1akvoIsl1l8UIkLWP/MxYQ
JFUsONmkUL/isRU60gk+XCdJzzKMI+D3nk8XQFl8iF35b8vmnuu5HmIAqZoJBCNh9XYYbxbayyEc
MEmn90RIORQECWy/HjakIWYzfJWqOOAk667Xgdq2sSiFO5HcFdXk70LjHBzVDsq/wKpmCIw9BZfN
nBYf7/8Sv5bdFEfYt9+H0pMfcrIBG473QO8aKcBsWsbHEJPvtpF2KsMDtgL4fb72t/o2yIjHk6te
R0HAT0hVWw1DdKoZdcxCJ+IVejHif7yLHPybswRcO/tv1N/SieuTQOvVEgmNc+xmxG2Jib13oJvN
gkC04xXhs9Gx2ylrnTLSQ9iukjk1heLNDoLHyanXYesQxyPd0Ooz1h7ZfEP7k/MMv4SnAVVBteoo
ijxRGgA2E/nILRgf4KzSzUIYV4ydCMSCFrNLNVJ6PGGbVjebnt6/rN/0gKUzH0EhP7TzmB6MF2Ve
RzKqVGzJU9zgEFT+wXrQAvEwKOodG35rDJUlK/8328Dlr/vkwy3YvFoashS/UGKVpB4rFHyvt48X
qpekop1hZKV1pLlrwKlX1fLT+2BQ4oFN2jRxnL6RBPNP8GdSo0SrdAiKoA9LOWwrYWr/GCq3c6Em
AI8UNbQLAjypjlC24fQjgRiyoJPmPeXZxU7H6Q+ekxVUI7jvUxVq4m/kY74qTvHA0O8xPrJ7Ueye
UD3O5Vr2NuxpW55dwGv5iPB+i2JGM8M18ScJ4YdXtryv2yzCIMM+DscCZi5AqffrPDWAsHD1bAqg
9VeLP6cxZddk8n1IEAK68XRY95THh7NySoGBfO6kWfW+USRitgrV+N8XuZS0Wg5NjNogUQJE/d1C
MHzcGMww80oCYd2HMzux/Nc49/vEA3AwdsN92C5YO00z5FBTMvc809QaY3XroYgi+Q3SHE7frSmu
kOBWjJ6dyPF5RaDwMwkqG3PdBGq441Yf0cEHW4ei9mRBdynB8i+nyXBGGwABO5FzRun5MPitJ3mf
/O0VnIIvOC83R7gl6D4xqN7tbbMiJNzKKzqu8NdXze36vX7bd/xXQA4BREaQbLguwLHWsefugESS
+vRaV5o2aNn6kWmPiVJP95DbO1xXQa2LxrwNuOCpMzdM2IfJKIG3Hx9C7f7dZbkgejs+2cCvcMRR
BZHOHC4K8euYA+DetNCkcioPm3kKCg2L0JByFmmfna1N+J/GBTpgV3ZJUzP1mZFvoLjLO1jN1ZKy
th77mMiMpz+GT0k19+jVwwdnLBg2BjTKlqZKYHGkBEqLKIqdjz+2dF8xJ4ad8JqSV4zktPnkltzy
KYW7ogrIrNGmJq4TGYi4cw9GuiDVcwMoLZ6QUPagluEykcAA03YOzTfClf0TJ2BU4lgakSk7ASMU
RJmvjIGTqASUtj+/WFXnrr+Nnjxt0KRXoAOpJUZKVVQa/XTaMDM+csM+5qycb9SW43HV28li1aQS
UAil2h9IjRNyR2X+rezEjj9J060AAinfzodcZiOLUO7QC0OmOqReymhc7XHegJhVJFMWja2yab4i
OlRI/R6pXF5q3Nq+CGIddpwh/KPVzrVhttgXedJRlTohUUNpj9PaRyBRM7VExfQnZ6cn8+eaeWMH
xOxYMeE1+QRwltJ8SgPx9tsEqWy72lcha58yzpVP+6b8y+k/JSTzDDpDSinqh+57BCpBkcSd6nol
pS1HZPWu7CMRML9Be+3NXReu50cqdfFMCFme7W6QXCcE9/xtuAcFqTkqgJC9pvNL8eItHBOKCuTg
e0gWRkh7Ua4NYSFOoIQgZveQKywdkX7/CSzv6vq287jznfKMsyU6Ja6QpAaXMRIh8URmKz6Dtz1f
+c/0tHSmEkqKiK5oWyzanSvFuLYDW7Tf/mzbMgNdnmrF35Eh4DifelM6SAznP/FJZ1ivIMEPYnUK
PnsADp3qYXBRTss+A2EL63Oe9h1dBnjmMG2dks/lpojy/nkYx4FCDKWlA0ma5cmPe5mgRANpUId0
LG7fDf9dVg0vJfy90RQdqb7mzVuqpk/Z3crknT6bnIz5yIN/2MsKQWrEB9zqTixJ51+M7aCupTZs
Zdz8br78qYYuuVwNU5LRDNz4wT/kRSln4/L/QncgeiRsB8OwDa0M9qavDjqTUzm2S1UkhjCdL1uv
oy0LspF/9u2Itgtw7unoJfekFtyDbGFyc0UjP0IQLPtEyiv3Be93NF6gcfA1/N6WZb2fpgDiPkCq
F1hjyObUDVBKJmH3bFiczwR+yfoGmOzT1wYfnarssg4x5+yhRKrM/4FdWwBXnezhpNK6rCFBBRE4
JNpqrV7b5d0re+DlJPnptJUFtYKPjhHDgMuekEfAWqTQgDrkxjEGM9hiTftzHKrxTA22vkc2YcMt
zvQNVXxf1waGtNtU1sKT19WMe8DySXQa8Z43rbRdgIf8cO2DTP3gzqLNflrqceGC0M47hjALR9xr
NvQv61Fsega2zpLRAwr0zvusYecGFRj1VRUKaUu/qb33GlXrWZWvg2J+LO1rwJ9twkO/On0cJrVr
14ZKcUeB667wJv8mhURtIfBjnEg0iPRzx81BMiAXWNUpYQLSgu9c+K9Q2Q1ELhaW41kgOLEiXoaD
ABfhScyJUyW7Uc8HpBjGhJ7WQt38S1B7gFKG/2ACbc9ZaCGxOsxNgd0a660dmw0JyMWr5pfBZamc
zJb+kJJC4gMv5GyFe2DyBQLA/hxdv0w+Oz5b3rvSRnvxbLbdgYk3cDYcN5ZqlQthgedtIehVn0uZ
0kS+fjVRxMak97rHLe4EtmSiQM0CEpqVdjBHskgfaw2L9DD5wYofhWKbFLL8m0sXrvchbw1eCO+Y
IlfYyGyLQHgQ8rx2RAajouSC/PCIGBa5tH2Cel24NIAhvVeBBRGvneUvWlaGxt3TQy+jMFjtMio/
3SCFZFzbiyYZEFTOe0NT5H14EtBsaAF0uUnpS86FQr5P3tkgUrzrA5PbuDq7gT+ImMhS06h324jQ
0ie9rym0suHibxLgMQ5YQE2xYEcorAsWKLy2oQmG6jd65TljnNHXYRoKpSjrW8K3cLUHkIOnH/Er
5LjqSBDxSNJJgLisDGiRw7YA4kBr8Q01qcfoNaSs/oHqPRhbnpmeY469qpjPaV3bxAHSSVYDEhMY
9V07cXWIiupaSXpzbpcQmwuezP3Z9Kb2qrQVrw8LAreUgIVb2XsSz3uBCjhaN8afNyLh59IRUJNk
iWZ9ReIY3oNxr8+eVw0BxFEgLnaXGv1E1FLf+ZhGo1Hr9ofkppocgH7g/sXA94ZTBPmkx69cUkQ6
3bZyObCWMpozoaGpR5k54c8drspaGF+PNkkmKvlFG2tg94GKocz8In1zFQqBIaK/qXhYmJoe5bXw
cH2PSGH1IUExggltOKZYDc1mFcJZ+P2DIQ5XXlIMbYSIcctHg8wYLecQOq+tfnJTwbQcz93Id0q6
ebaPFMD3Pb9/Txt+QIQG0BJqrEEzUYq4CW4VhDFUjmL4erBh4eYIeS0T40oSwqmvWxAyXADSyC7x
G+TwOGiY/1NE/sBudCBSsG5SP1Bhzsa/2/lZu400ORCSZfS2gP1BjaCA+U6fvYISGhmEcr3JGgDS
ai+vpyy4s25eE4D82CXJO+exU+5dSOIKlmsMFX4ipf6CRgUAfsLndL+fDaRBzLtxiuBnbG0E/6hR
NJ1+iIge4yqkKACLdRgPdOZIcOc40SGNS7M0tBhww6drYV+N/sV7F8DHWuf12on+r/8e5L5sHXu/
c5tGjD6O2R3U2T856MELPboRs8pH+RPC21HiahZ98tvlGfYr8i/I6oUA8HNTQ6eMrnQrOkubTY4w
invV96iJyel3fJPBmcBlclSLvZp6CQSJJ2GjSynLcotBNaf36scsvetcOl4IQa/s/WGg6p27GITy
8qQL5k8BuNaedpPCSXSsWYw+hy2HvQx3JLN+IyJIJgQhKUI2et52hR8OhWjWLaLhmD0eH1FW8UW1
fiMnukyHn/631Oiy9ATrKFDxABtn58Wc3GIab1lGOEwoIrHPoHd9p7A0Tt6yvJoslQN6PnpCFRC2
XaOhOXMi/hBTcGt9my1NHJ+KtnL61TWEj5hTVSO2DXMKIMdBH/iHsK/Hy7/VkaOCyH6+d4B+dsKk
XToK3t5scdBsOIvoqaZx7Vekku2Ef5HuZPbVmvc8rWXWN/5VMzUtzYk04OW5tPBob3v30+SeHo8+
vEBBDcLGjAVelPLvB+PFp7Et8Jt/lAxg7eHQ2Po9vUqRJRQY1N0OYrN1ifHdRezMnc7ZvBa/gWkp
j3T1hHJCcUa75GTCjZXQkkjlLZfZlPAV3HvFXyPSdb0qD8dhzJzLWcfxQJQOyYsc+4F29dWQYw9R
ph3LNPUnPZO/CNEm9ZIT7xRIrduCx2/Jmn3v/JGfC/7sjaVUO0p52pjfnW8mO1hf11A8yMFb+Fni
hTHFihEFvMWdHmK3JowUfI32m6DfdPjeQzoiRw5174PG5e+QR1XTRwMQdaGI4wFbZ+0DNd0rZst0
iHvBwCl6Dn/x+IJ5VaBgXV/o4Eou1ppPO8/i5u7cHHCdvBZchnO8Hm39fe8wjoJ9lFDmrwZXDFAu
hklvSouvUHd7HhI8X/ARk2x+QGFrs6gkMz1JlbrBdER1rsk+rmBtALGIX095+oCfsphxwHQJOHQS
vQrxe4mMLg9po8b3O8aL9VEQ+1HM+9AA4Wz8jCmTjL3BUfoMrDiU5VtZfX2JdiqXVCO1/tGcIUIo
2EW/1glTrFXdhGit7ALaaHk3Ip2J0s5J0PvfJVS04lViLWqztRP24h6g6bofKKJacXIfxjmob1Mr
kbX768Gm4JK3EePYlwbX5c/a+hlTzsXZRqGzrRJJwKjkg7hKBceD4BQXE9zuf3hFSeXIWosHk2BQ
AXtUCF3VJhCovCRnP9xadt+j1P44DUGAm0bx/425btmOd8jiC6fPKt1ke6WEYiy8u2/ICK21+56Z
K1QnE3mU7jKucl3z0JgcYdcN6ql/AbxosSw6PRuAaelGaTudO09sr7vKFQx1AQEale/vtXywQb8z
VgLbYhZDJCj8SPIZo9Kazt5YE4zgCAqKURjU4GKeWc+TbJQf2f0S5oL+z6ujwz0wdL2b19Y/8GSe
+q7gLzyyDjepXzte2P5lvGvtPCjLpiCjJJHfdTawY3yzRuzRFtOn9goztTz6PuxEhVDST8zuOerz
OxD0P8SEjpKdDerz8ZdUpZ82hx2v78lANKc4bUF9A9r53TNVX0gyIPalV4YHEP3fsRTXYUwM53M2
i3simWAJS5XNJSPniNIOwMnQr2sxcSKInfvoLxyEsjDqvdia6MwTSFSu/tQO298G3KFZKa1U3QhT
l5APCN4jIVtSGkK4nj/QeapnWW8qbqOBbkdCwB6RVY5YaYZvl5dj2EFMdkDaS6BKoti70azXi2kC
Zo2DIz83ZzN23QVxHtcLUtKplycnborHoq7+TaE6cYkxnnzCNUG7vc/YXCzD/XSKgxb/Qa6DZCCv
io5MYtHboPdni0J+YabNrn31gX8K8P/PjYCDalXVqQc8AA1anwgYf2BmpN4qUEp+T+wcK07MNDmy
rfz4smBbLHoJuSibRJhiLzfV6dCUwpqI70tAAJbi2WTuuxBc8SnG6l7N49+HJefAjOx/CBbn3Xv0
ECRF0QsBLIWImAdnY1LCIls1tSpGQzw7LMsf4dQzsrFWDXoG8fnVRae3b03YFaVZsVZZABM8U3L0
cMjyuZmqYSfW8hHXwiaQHdTjwh2qE4qyycBFEKQFYey56QysGibrCU6ldbpqQRQ3vs23KXToZXya
xGyDvniyp/xeK4vV30RjF2Af8Kmr5rMvwirEJq6+CctKMuNnYRAF1YJD/zWJ5JF0T3V/9dw2AcBP
CD5VZA+ZymDAPSvB6hf6E8+YCm6VjnExWynhTwjOBXOR+m3IpEaO6YQFZNcQuqqZWGMM15+HJFih
LfFeau2Ra4HjzjeqBS/9cBnY7lQWkelGtP0MZqUBSL/UOaXl7W7xVSPa/XoFay6o0XZ/e12q9fpS
GAV2rbATWdKHFt2IfQa/yGdkpfYmUHQOvF950d89vOqRoMQSCEySJJCHf8u9ywxTgxljSXCi/HXr
P5+u0p1XjSXf1u+5gJ0RppVU9fVJBF9nEG7qvb6gCd8pPpKXvtt6xhBdqckb6EtLDVhxHYajnWgG
P5Fh1XI1LxQB9bCRhCLVjUynigWbMxxbm9f7dQAoHRPgfWNajrBAyycF+pwfX78i455EHQQaTFvB
0oVo3dZwo6DzYSssJyUZNXeVU7F148RJocb6bR86jU7I8GIaajp6JakgBP7dqXF4ysgYq2bpE3D5
TRw6/DcI3Yh6Dl6WVhTDKPh1A4WgV41iGwJRdyLHThHDGwm31/LGymec/jwD7h7/zMcxjQEGhwce
ygB8CUvBnr0SB9Vu1P4SNjdMIqC3Sd5rgRe0LJQZwSVLolSo0ee/STgZZsfre+IT28q7tMYoY4Z9
H/1ILYNXtiGvz8VbB4IsbHbGXdAQrvbBCkC/D6z/52AMbW6BP4je6tEcmEjfVyx/VATikNM8U3bP
L9S/Vwet1G+gy1X76B3u0BVzZepHvyaJHZ2G0qTa1FXZ6D7bkacbVyWkcRow2fcQx5GV9DsGy06U
p8HZwR+V1Lne+vae/RK7DiUc+7HnHjh6wJbP68GiNXI4OPvmUOsYuCBfZoUVLYxDMk9k6oj0K8eP
C7uwgndvooYG6kdqn+iVRD/LZ5Upj4yQYaaPEy2Wtu15v8SctvWaoLlmj9ABJ3iTXF0ItLV6klNX
p42ilnbI7ZKqsX3qSS4y9EuHiaj5h8WrdbLOo0KsXi+zyObp8Kdb0vyWKU0ipqn59RP+aVN4M2q5
9P50dpg2R3dK04aJraIawvtkvm4G89Sf0GDA0OvZLpwIflGHdv9h70WdGIxZBJDmqtT/QM0LH7DZ
u1Wa5xX8Y4oXnjB20Hs1DNMX7zxbqKJnZWdMXSTTRMCpBQS/noOkQAOzZevRpUQ+RDf8NHVVaFA8
TXHa7IpVsasgQ1gQcjSxF/2xP7fgXhOud4YsIFwDdsOYNZjA3BeA6Owq2LKZUsMQ3JSGzU0XfvOM
Eka/ZZyevTrU6LaT4FGjc10F7PjjS4oYqOSEZ6oqvjTengkIqHgYF2stv7QBNmC3nHtA2iMCsXrW
ocjZE0Hr5z/i75/ue6x2eZPajIdFpRdv1qAxO5G8VVjxtXxIBdNiIrr4RQfo8CH56gzyhWvFEDQ9
hKsvswMYKBpML1i/WqtESUPE5m1yIxRFCe1PvzlxVD8nKHw3SQAmykO3v1jFC9zJ/+O0xPtsTUUK
dikG5UzOXEB/bKB50AL5V93LWZuEMtChmsIUd6KZKG9WKhn3CDZbjTZNDo08nkJb9BcY8MuwuiWf
auROFU/7kSMkVa/47J/jY4ZfHN5DywGnr4MDNIO3RGJJYa+AoLl3/gLwLUhSzlGZcq8zf+pslHsx
p/o8/4U2SaMhn+fb+EHVw5z0BrAcNfCAQXrQExazfaqLz2JLj4lKqKRZ2z1KAzW3XSVb4lDPqoh0
mwoAl7lzckFf5BLqkDc95Pycs4PqYS5C3tq/+m1a1tIa4JaWRVoLxA1zeUhlYTMaMRlYyAUjpJCT
4THldtjmud4gXE8D7GDCBVxMJExm5yB+nWtS8JZ4NG3qLCYJ5nq0avmusO5GbRXP2PTJ4JO2W5i0
yr6+F334ELuczvtKVyUrRh3bSPQsWGqVXIhCaKdWsuBAsBkx7U9UUYMYlFd3QhRWW6/aLs7tf4Sx
xK0bwlzAo41GmALF9P/lW7YA3fyHevs6R1QV9mskygqq7dyXJCOpxFNxscakVxDm9yJj7JOLemEP
RdzPzRtYaY5wSEIGCL+Y6zHsrZ83W3BQXlmG8MKfmCr+Yjjoji8w8+/R/b5EKhKdnQAxZQpy9Njr
VyafMbyr3TQ4o8aYG9dt8vZRR60Xy7zT3mNyOnGeSiCnQz1PwXQAVZl8di/RhSbo8DteONgE/sZx
R2N2C2mpYyIxXPdH44FRchWMNkqCIYP+tfvEhqq5tC641QrCvtplFC7JFQPxW1/jP4R8CfLiZ3Kq
QlLJDb0EKCucDijDl10/7BTuYuiAZoP/6KI4P2BAtF+4GZo8c6ls+cJhBVXaTlOZLNP55Os5Ooga
B4SN75/L+Re5xucARg470A8IQ1ow+Qr/M327Zu4FJEdj8ohBkIjd/A3y9w81Z5b/SicoO2qGPkhA
QX5s2sBMvZCHeK18Qk7nnkVXWgYeLa65jX50xbp99fZjLocbEl5y8VNw5djGC01LJLbzgH9Lf6im
/7o/R2Ll4lU7xlWnxKbIX6ltxLUYF5epfM1WZFx+mFqWSczLC3txAMQTJ5GtNwVyGyUenhVjZ9/g
uNB/XGqnt+HkgpaSlfPA1n+hNMjAEAhTIlkVmLEAbVYheB7lg5Z3w9nBZnOV7It6jeZFZKzoZivA
mHLD21zyrIMSyP5b/7jkJMMLjvUppnlN7q9EhDIQF8d8b6tklDJ5rVYVgMA37BK5GWDfKTpoJf7e
p+Y3IwW3XMiUMnqJ8IByJ4UL29MwORfktCMXjIkN5x5duYif+TgSvpQtkA7stY1NTx32dZcWk9lX
Z8/zyVPSxQovnnqF51WejL7Tp+f2s4RlNwjI0dLYhBznXFDMCFaftPwDW9MUA4AYsnp9ob6kY6z/
sHoCTtOfjcZUWaFnl/HHowV2I9ij2D80CbHXqK7JFMBfmZYqwwG5CLojWgiDz/ePkWyezA8Z+sXT
6ZMLVpVEfcLPA/cqJ/Zni3GZqArUzb4bslLo2cIaoJGwFgk715wLhffG8jv46LVsLzILUq/IdLxP
vSQnLmpGbdwugsFmAZCccJb462kTKU4cuF/m/Ko1dNIStZGjWUjdT9M2fGRVV4jglm4fU9NYeyQ8
dVv2Y0d12C77zuYg/55Ho4MoA1gF6YaVtGBVm307gfXvrc2laskDADJxXtlQO5dwxhrnuiuYvvVa
jM2bM2lzDSRWPN6CxxZguOOC3pSiOb3jO8okWMFDUK1E0LfSleSFvV6/GgjD/ei3u1buqIp9KrP6
zy/jwNwqkxHS6HVL0uhxdjw5EERF+P05M64uwNyk+td4Aw+7Cd4lcAhDKFkFaKGvsoWgcnjWyKbQ
LDSoHCWIFSZ0jMFsXuXi+KjxzbZUooLeQpMbt/lXwgbDhpGZXZUa77x0TgcoCGMKEVDQw8KU8dRv
GShZ0XiLjWiRI6sTaM61jR60CLMwoS9s2x2xXp063sEhYm/yJ/fOZwf8Hp5LT5FKXwEFvSL/oPlq
1Su8d2wXhZ8oUfpz0J8pgXbsohHfw22xyb/rovW0ewrA+wryEqVDfPLPFt2BH+fa/fWOkK3T/gD/
T3a1+AhboHPPJ2tFYZ9rgyn268iBqcnk33ydGe8LZCSKlP8cDxY/TYT6qqBgkAOc0ToAV36aBrWd
IsYoSIBI5qSaJf6esAc6Abi05+bwYmnJkful1Ap7Yt0zIcePF8EtTQD+Gd7i8iVxdvgbyf4zPmd4
WpgfuOXsW6K6+lwTM/VGUhuyUIZ8UnIsut7R5X5D/CrspBI11P0yixGK+natSFmgvv3Tyt8hQg0d
OQfxd3T5hodbtbgub0x/VddPf0fcHhJFxcL4tsm49KbaDX8dix6PP58wn/G+KM8P0xv7dp/c5nrS
l1QmN9wB2vgk/NefIJ9yDtu8Kvi6Ov1Xqry3Gr8L8k9ve1ECZCZdYdX4l7d95BKpFRKgRkY42KIZ
nKqURrIhkyeZmcy01D0JLNGzV31F3cCQ8rtNV25oH1hO9ELlefKTKGGutE4B4Tly3PTvL/P3EgE0
6j4pLi6qjtWA5L+Y5ELIJFzXEQU3mcNpOj1PsvIawXJIdaEaCfF8vDZPyfJEd9Enk/1u2KKt0urN
Sp03hKUXVmjKT9Es4ZTag8llcLV8STmpJMMiztZR/KsFEV/kos7fAOmQKydAwfF7JDh/Ue0QOiz3
uJPfZrZG3oUfKvzVH7f1DOzlZj7jJFNWYknaV9N0Qaa4MCXLSQ5ZhDme/ZWpu0wZFhgvtMI76Y5j
/h28maa8Cj+lAIUbzOjKriCdiNP5UYUkopvOzWQ6PbSyPW6ogAoD1dmO/E4Mf7i2Y30jZ48JySwI
qhKqf9wmIuYPKaKWKj0mktA6pL7LJ3H5eJjU+BMck6iAFFwSAMkPhvaqIidxy9jLYvL2GMu+rHqB
6t7fTxW5LMMuKPytQCrpwgPw+4ZRW1qcdlqMasMjbYpvRFCy7SMnMkkr36ikDw/Vqo+diZ5/j/yR
4NvpDf0+fd25TkHIbqTGHy7+xLpOYSFwVJjnecnMicTEhPfJ67FNJBGJcv+7PDmQSD9Cm++HkbSk
37XJln9m8HU9pBAENXVkw3gGBTGzslsV4Mki8KeydVkRiq3pINyZilcN2B2JA5zBvqNbzXt1J5Lr
Js1VgrEYyJzqPJVwjFdI7CHavuq8I3bbVTxevpBpy4nA/S58LDkQFfQOEPwdqkrPJDU7aunKYUoS
eXOKlbQleTMgyzCOG58WeDI=
`protect end_protected
