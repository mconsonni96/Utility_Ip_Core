`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
U8oS4GRZfU5faE/Ha+jK/4Vr3yHG+o7sMwNNHyKAZyR6FQ9tEhROR8qguVxm2TgJ8YRN46qkDAuy
paKiTatQMjma4pncmjE+eGoT14Pihe9E/ekTgtrEy/8gxaoG3gu3zt3yenPdo+ESDtNVK8sETlh6
lvk9xDy7b0IAkG9cTe+h1RWa1KPI5qBZhU9belY0FGTdhBC2iT+6ImncbML81Br0TcaVyB0pdUT8
/yQxZjLZRByljaDMLz7Zb5xHtfskUwir7et1H1zDWiXbDRvvC71vgPp7/+25fWFXMBrIQbHh7H5M
KGEwMZRgVnHcRm+DboXm2E8WnW9xRNHf+TazlA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="FiiuI3A0QT1jx4clPQxBXnHe8r0NnpXYaWK1unlpHRo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54560)
`protect data_block
GiqW2lOH+GXdm7Nq3Y2NNAIh+SRPRX3XUtXUtgjdw67mfQZRfS4/TYpEs/LjoFF+UsOsBE8dULHr
AFkokeYm+uuhMVm718KRIjkO6WWZF0JGO2dZ5a1J3a07E0w50uYvMROnIhFCXTCeXGT9h2/pLROX
gQWiXa28R7y9xuuVoEYJ9lZxzNOqbGI8nZ06Z2PyOVadS7u30MrPiLkb3YasyYHY06BuHGMisdNS
FK2uGzx5KTI0eNLtuAIPYqw1b1GrQ2uo+4uK90mvsNQCeTa2MS1zVlY0JIqjZw1gsOMrXufcawRn
HIgfAdu1kgq7lu8i/D0dsuN6vfClimRxrFXch243wBrRsoFC6oRy2btPIqErS0xdmA4gnBnlIX4P
e4dp/YBkS47JgAsCvhBbOYZPWpydUgAPnv0Oa9PLgg1oWhbF7fiQtB371/7CsNNqcxhKNpwWV2XD
NDDevT8Ag8fluK9ET3HBPlqsyPle0shBF1m/XtQ1vHqM/3bWFcqelgp04yQ1xuda4oqn5kNlVaM/
25KBx0OKQwGuH093fQroW5YGC3V5KtVWgLmt5D5K5ZfOAw1zY2hjnu64mVhZ+oDgnHccyE06A3iY
PZXyFuK2qETFsyqssYcxBczXq+V4WZOD+xv/NpK7ekLdsKdV5pVXauWheD0vKRqZ1npseNXPHDPV
DY8avRHGDWpMxEd1uSAKmg+dLoyAN5IUnvDZBwsjYRwAhhBNTX3P0KNeX56o4SpKfGoI7m2TKYUw
Wp3H+Ms4bOFZ8qnNvSaLW99Qsu5/jfjfotdQSRVvplAM1BTxttfRAnOwzQbwBrJS8JLscQ0ZYOxC
CFnTRMj5mxIRga/MVI/wka8SNyN3OtGLmOWjLxK3aHNl3RSGkP9GDnPsWGTZ3dVmuCAxncoQF2zJ
5UDJAbmHvwwWJU4UJu386Emu4jLQGDJE3Dvq1i1XKp/0jPhjVCiSXZwiTNsRJrxyEgs9zqLYKBL6
L7Ld7HiYAy0GbZafZ3OJ5OZaaEmc6+qqlYosOgr8n+ai21JO60kkof2gdEqlsRCV6FMMmIzO+BdQ
l/qkFvl2LsPdC5rnSLIKYVIbdZhScFvLWDWQ2Ls/NtHs4PN44Drd5nqZrr+O8FZmvQpFpnC7etio
vtpDErfZ6zktLdcRqC4mxgOezQGQ+IBkNq1KYWbWaEXzunUPVLoOAsTe+9JKXcbeJVSz9vDXNc0G
JMXUBVno4Hiw56tWxPTLwevtCivpZn7FWr0JNh6lwLCU8Vo1j/NL1llBXmpXm2gSlpTUjV1hYzAB
BG2E6HKaaCoG6GK0tnR4v1KlSvUZb3kT33XI0Vh4Hl2qFDTtszTcpGj2ICJffR+Ag4xs4WgaTMU9
xxUyba24O+gCWjJ/Dlv6eLRGTruzlRl2YR8xhmTolrrECy5Lbcgw1D9dNerH1Ki0rIrLtHfuscSJ
SJ5ttXs8XMq0WPtOcF6uzPQyJ29GDbAHjPFz/Gvz/SM8Lm8GhQ+Gwv473KKWSdbBH9lmt0LILzRe
5EJmQB7+tX5Fw94X2eRIV99dj7Y8BV1KZGCt6QOkb5tsF8VSglf1N16d9ZqVSL6grltstW5r8gbn
xCeAZBulBFiGCWxz4TuMfby8W3d+cZEVcnoOAo3XgEDmbuIi8o1Alq6e75f7vsOhMSXv+FLx18V7
vz+XJSP+LbYUHRbm0qg96OhZL3V5x7gREkUabk0O4hEtWK50Y9XoGp53NY2w+Mv2C5zcW2R5AbLF
k5b5TVjguevVsVf7wKS8x4jGhvdw3Lsuv/EIyQ81jH1CcegPyqhLGGXNoMMuLRamdB5oULLpXCQN
dQIlGD0csN5B+Vn7p9W65bgT0wzrZjaKQP3BohhqlOj+YPaVWvggkxpQ6zhyXQym77zRC8mE1Nir
QFqWBCBrHz9Js8EZJsoPUJujN5C9N2UsWmary0LoX2OjpJ3K25+/2Lr+l/84XLppkXy8PeQT9QZ9
c6ZQ3BO+lEippu089qWzQuUq0I0Cnjta0X56mMJ2cQnjFc/e55XhxsXJfFBGOYJErlHt3wgWytB2
8NU9QyLnal4+ceHIpQwGjELnU4E8ctUlZEV6ntMnr+o3Ij1aOQup0vg34mUFxhLr3VEi7x41exx9
MVNjiW+t/i+N0UsXBARlojjf3HaINYR3crJ/qPdG6dFLZ04GV61V06GCbPNlG4HV33Y1wsTh2huo
02RRc5PgQ9kZxrXrAA1K3M4z9UlNp6vbkNGbqopAt7OBN0BHb7U4X9kQ4F8qwSdSLgR2oJdJy8t2
lhEJzew0DukVhbFcSEfvaQbP3lu7wsE4GExXfu08byxCbVOmQMVuejfQ9WQKktQJIZfYVM36w7hy
2Az6g4ZHTzcjDa8HA/IcQkwSdksl/CjsqptOUycbAMJiiNLsv7b9uRRdiQuQbFHkEBEsZEkxyPG2
LZO57lSnfcCuAzv4JTS9Nec6dAHdSfO6fjpJhH08OgsysZSAVRHp8h6D/YqdlTXAhcUOH+kGbgap
WmeW3aOTON7G/9WKQQG2EHhPY5x/4+s3qkkCY9xfw8p7vRN+f0b8Ja1CboqoCXwODRiRmwFo56e7
RrP8EW1kGi4qNKE5wm5/eRhGR3BtOm6w8WHqDRUaS79ma0Wn4Rn6po27rv37AbITYK0fqSmkvs63
Dxn8hyaw9n5phhgf+JRAfxxfaSHVCpUC4BmXkWoDFFL0LGXdtZjasFECZFls40RAX9bkM5rHYtI0
DlQ0O49K9KMY3Jk68YCSrdO8y+nbMfX5UbEQf8BLzktSj/AL5xF5+cz6W3Vki5E4+6Toybm28/fj
a18IU1qbs9B/nDSAnhgFQj1r/qOtqlTow7I1cOCSuu7eAaYhzcm8Uzgb9zK7KtBmtpuWKUs8OJxz
0c1guNTZDd0n/GNUaXubomgMNnTiGYsqvzNQ25nWdaCQijO3hklbyNh/UjfiP4U8viGySA+8f3Po
ZTNihPxXszUMsFlQFgMQGdz5lVObJ2yGgDbwgHGHtdBGTmq3NPnMIn59Quh55Xcv/kUPSNTZMWmA
N5NDk+dEOneZkyjIUs6Zd9itQNULrcI5V6fZAN+wCCTYwMyl5YceGmLv+b14fMS/lMGc7tGPSGJE
EL9/PjnfAyzk9IxA2vsfhInB8d9bW37pvteueSa+YTy6/EXC+f4O45eJ6xBUxFkspT6wfDU1Cy7B
cTsndWDHCLPaQrNhp38Gik/Rmn1bKxyUMpV9yAtDC1ZW3/uAiJNMgrbbJuJjHhHZcPVbu9d4TRn4
O2HxygIJQAntFX+UY/43Eu+DS/b0uW/VB2IKhKY1zPGd6rEF1TSOOSZDeatz73yPzJKXc7d/JM/3
igG8V7Xss1p+mCbGsBD8QjMOJurrwqDov7dn9oHnwOp9bPJuRygqrVH38vMWqatlcEsK6mALEtbV
roHJ5pYtge44pb7gG5ENQxZ9mee5BaHofGhVsdWA/f6y22iSkp5E0pBMFzvjHM3m6L2u7+AsAqrF
oI/kAxH3btERRk9zOXIkuOPnYIqo19OiZUlMAC8guAhkNvm/vC2Awha4vFvMIti5qW1C5ZQUCSJo
+IJlR1PEe9Y+YTJDVHuaDiErQb5HQWWH1jDfq8V9MroB520YhjecaOaJWPECTnnkwjlClv2Ml+G9
YUb2essUMjMv5eJEA14ZIlOvF0sp6Vniz9ljj4oZPrRPCJRd1d6IcnJj10+6cxHSO6NFgJrNbmkn
qblxbOYbA9MclaWaBTJJyM7B2EZ61ugQ4YhYByysdYnjiBI0WNnoSnEWEBrf70OU+IV+poJ0/JFw
xmsqFmjYWiZF6woPfBmhauSzoeW0mXqhtXvwyVPcZJIlkqo+lW12klYfuaijnTD9C5M3S7HDSGL2
SOVx/x1Pvjx019osmklXxUMHwVpFRioNfnWV/h0v6m3qCQC91qSMAd2j+hG+2devg/6oejy5yZYP
yHSkDIeW1NtcgRa/TNUg6o6RCBP+pOI2sy5KuC56fnSZBd3LAZFLx848OazCnipSEfWl8Rindvj9
HZhixG4nLKiTXwYNx0wr11jnWWg3NuVXR5YvNsU2V50N++WWVQYs3N9gIcBxaIV8X4hWnKG4Zj8K
31mj7cFecyO9pGv9863RRiUnfXDxQsJWYukv+Bir2jjpoLnBQqVZ6XLnav8EGH/2ljSXVpFekNAR
G2/2yRlzhHih8fetBkZr4aDurHdqD3Dm7ZETop1doCdP5w6IEBtRT4SdI91FWrJnCW0csKO5d4TY
mbingZPk8Nz2gSwXzneiswUnQSRXM1TteOioF3n1Kk0g6dPkoKVmKuQtURkttAvQb9+ipGUSDkJe
svkP9wwqT6jkfcPO/XLMWrQDPp5CwpD66YyNbtPWhPQRrzWYNCVWjmzGG24QpS+TthArciKx623Q
FHhxyOwvVyPHDtaAb1heJ+Vc7+TUF18XfH014CDlrhN9XOFXXKk+oqyVuVSYvQU9J/Cce3+8fbGL
BrfTP/Lazyucu3CpEeHq98mZ1qP/4r61lO85WqFt439LIZj2w45RVoQZ2j2VICUoZRKNuoTl2Ktz
Og95K2vsLZ9hmD55uTWRRFEIXVpBFFrFRjY4ZmEgyuj1gDWnjVEnGAnwjbLOSIxA66wmOlt5IvJ3
hx42WN3H3o7SXsTjIllokrYwJI9okZBqAtSrkVvYgWZlUEBTeAXTYlpph7xAOjsac7wVBCWAQVv/
IMiN0djS3kxTJ/+XRhTD5Fb6ZA5OPfvC14Y3sEXUlrU9bpXn5OBSlaUdc/TTKUExkR/Ums+rtEmM
wP88vNwOvh++71yOwlmHOrI9Rlx/6zRqzht+O9bBf7ahibvxQwBehEdMzv6/rzvNCwNY/g0CyOKB
U4Ka95BltAEJFrm8IVmT9ptI637k+rSedJ4D1buXI/Z4bdG8LIJ2+CpiK0sCPrMf5279FDRplZGg
OFhCe+CCnOKeoK6CtJ7CV3KWoqdd9GDKU3A/LDkZbjwHPkIHHPwRC03IxPkpMK1/7PAfW7u4IcNC
j3xXWsmprsoauLNyh815XdllmDGSvIJhK7MYZ9PknB4eTkFGChyZM5Smu8wAtQBHBMvpuy7TryyM
UtvH7UNkfv49LY6vNPUFqzmb/NMWeygd9VtiqQ9/N8yZhXh0BFUAgTXurjVaoxOvJBu3ftfYqu4O
cqCHZJXLSGQ9c4c1SRKwHS9fWavBU7Jlq6LLJS/MYHox5n3nMeVwgntw+jRTm6hsvn+aIRVn6suZ
p1x5KXNDOLqrSIoVK9w/Yb8kXMBK7stRlh+qPU6o30vwB7ftS8MxvXb0vNBZsHOPaedY29bbOYsd
REs+hwriuHj5eSlNbRwhRY4E3XsUazKSnfXY11vRkSsHpaMhjBz+M14JSe4qW7W9C4wXKz3p6N8h
Ypdhch1nNew/C3NYnYnNX3Tle9xWWh88IpebkNqQKTRQGirZjIAy8Iq4tyMl4/SDVih+4+X12ekT
u6nM87cHg4u/1/QggjQLZcfaA+BL6/eJX1BJZ78APil0E2ifdJV3u0vwKMxjMf+5n5S3V2fg4oYI
M3hriy+KRvaE5jAJt5U0VMSNYDJKKif9EaqF7m3A+5Ikb60OTvHw/EVePsDOkew4A53yyHF2DL/D
W9G6IkdF4FbnpcDddGIOx5AJNDkp6Ctqd10KaVbGvBVXgsrw4bUiAEaevKctQE0nqaZWqnofiAE5
rUQhi3IfbPaDy8A/scDetho9+nm+Rh69qUZ1UK3DdwJxEzMv8GaiMiTTi9AUmaHIUVnMGo44NHk9
XZlH5L7h9wxjZIlGYzQUT2J505KijKggPC2XJlRj2X46Aq5DxUjF9yfYTYaHwgEpwKxPnYHBSNNO
ss5wbeRkFpO0whl6dFVzRGPVQE5R4Cq5qljlnLO9URt8ZqXM+swnNwmbozElfFuel/b72opyO6ow
c4jqciImkvKXT/xxh06t1RU+46Newu1GKz0AZYNsvWkAo4ZPSu3QGldOVAvnyyf+WkvlsERYdbfs
qqg9nfh8hX5ItHFO8IVBo0e30BYWal4gVcj5BtbllQ5KpvotY3rpZLUV4NBXrpwTSn5/bt/oGfj7
tMFekGRxRSaWm8VW+bIkA7ZEMT/TZ8yEzITQhY4zpPOs138jKLRuhYN563nu3qRfSkHyccgKdnE0
PWxHsTpkQSCjphWK8tCJcBGypuuycjcHLfA9STZLP6BS/2g/unyL/DLSxtDos8x8BuvAB2gHQ0gF
NXgYlGFlwk7Rv0e0x2Pc8HwFtatn/TwsHZRfvNhkITkG9lcCP8b9bAfj7m+qkgc0kWNNDJHiTr0u
NANG54spHxxLWtqBMiPg1lBPSh/K5iPW4ZPXx02n9fGOLYADD54LIV3xVupQnurB85TLe76YhDDG
U3eF5+0kfAu8fHVxrUCDvtdNiPKhxi0iZ9bf+kz2+x1pXU30gK+PcfSP0lnSE7sH8433pBwjRE6t
8Cnuo1Sqb+sUv63VkdLwTRQ9Y3ER5XUd77wdR5ALWmPFgDKHsTv9oOdjL7sMy6GnorJSt5VidNov
H+9hEyRLYE+XEGplZJPBzMn+hT01CDFnAX+BlFnEr4lNRAu39a7h0sG7iUBDCh99FduVST4UjZLL
FtnDz8lz5Pphhn1TOIInSwU4e4oms808Sk/cU4XN7vz7vTT4WFi8LpWlisUn7EowRcY2Xak5fsDz
Cdk6e8vjJ1jgAKwKQkrnDFToIVGAbmvWfilfn/VvfYdIhLC3svtOl7t1ztWuAp/XIUbfuXdWokEo
zwJWQ4UuaHXs3xGqAZPa7WJWvlNxw4i7/YjxjsrjbCMuS2ii8rBGtQyjMfTTKgfx6KiwdLAxCkPC
FSFC3RgwTpXur/QpeilbVWFN4GXzk6yv/nLykXHqWHyIZ+31adsAZBP8OQtJcq4cKxF5z6JZqvOP
NVNYNY+NdWiyUcbSy8bs4bqxutK6k4gJsJ+WOi29eArMz+Sv98Lpu0E6JoMx6/BM0g+quSfle0Yd
tGU/ZdOs5Lfykzc/xUBt/6gsjx3GyBtOURaFvytILaeq1WYXlpiR8jdtGQADERNKlJbuh0OV7iar
gW3/SHKpT9Jae6JNbsDqfems20LCaBkaKNgPCnX404StGkEHKa4+1OrWJwzJxZkYk3eUEjlciYdL
hMwyGU8tk82uM41W9cVF7HWYetOZzADCyip+IOvQN1Mbdap//csRx2JryXr6va3E7XTvKStwm0IK
Yk4hrAxW8ru4SSroiLBxmCSDzTcaL/OHksYnScTpja6GC1jvfNWICCiYPdeuziLdVTCGPTsS+yZV
gZMPynJV+RbRtoE8gg6dFdppa0C91IlgJCAguEG8lbkVOxWX4tewjw1gDnDPKs4esku1JqaXHkts
P4btsNBWSXsyFMtRLcSRfcMvfsWkNe1ya3AQJlxZpZ+EGWIkrsLYf2Y4k3IuLDUsI/Sz9i9DG2Yp
IAA4Xf4vb/QBLsQvNf1eLfqX5KkmfnED8P6wx21cH1Fj4Y80AtFkrJAq8yTwAbQA+4RkUX7zM8KV
zelgRI418vgKIxb+bAYwuEbRwEjtsoXAjh1RKvvweJvzz+FZn3AiHQoNsJR/uurLjU3i/M65gd/K
4pe39eY/2bjJedrFxpW2u60mq+6nI1+j7oBBR6MhJuonZC72ERv9zY3K9jFvViH46B6+6SgNZX1R
5WjVCHOJcMK0W7It0PVV27Tn0DTLkZuOCHpdRfgcUhIfHoiw/YR8mkE1nrWtUuDdhIm40VmyKNvT
Fe28CtaTZN257UUlt3HVPOL84atvn/3Xnth6MxXztvqMmmVWTec+95xvAjwNBUBoA8UsFJI/0Jho
oAlUJyCsMG6FWWfy2OddWSGs7vlxBaevNzVWbYJmykHkW6KnoFvmFZ1LwUHRAjNFX7ZJqzttJPGS
pPN4VvvP5EYSsv8a7m/07fhuiBbht472a72tB1AQFUc5KdMKXUjX2BisPSd8FXrJwYoa6BRksHk4
M52f0olkqKjRXGhrtBA7cxLgVsmZ7xLspfj/0eNwxjy69A+5bNsT4TKgivPQCPrAv9E9fKl5jt5X
phLWwZwfelPXBfiX3K886FplOa5zS/w472qPO/njHsclCIm0fW8CVVg0EVkUU4z9bIuoy4rhX633
ntbOYvgzNsSmuaEl4OB8DUNTp20l+loc691V1xSSm6nYoMYoyw6q0UvoU1Lb082Oo2VvEali9U/8
m4VQBiO7x8gPv/T67pRiKw4jvSrEokp/XPFoJ5CPLSTFXYZp2n2HwPUd8njgzkmu24mC+3rp8tS9
6Nb4+rpuD5HU7p1Vdeed96nErXm4o3yJfsgBbD7bcpurwf93W498LX2CKVkfLgjEt+xSc1CkhjD0
qdL4lyIik338WthubZLCT3nnSCXL2hI0rRZS7C7c8ECh9bf7+p0WdjD/OIqwd4ykpnE6Ppjlyagh
y1ayGfd/SWtRpESuDJ10uarFVNQ7OvwDO3Q/wTFjgHTC9VOYPVkgklVSIqi97qTmg9xJYsCIRgkL
t0Git3ZpKtAolTxy2ycLIj9Tun9DDgP1f46dzDkJZqs+aKCsfgYVE5yTtpYsAI6YjV2GT/wf+N0q
Is2ObPdHr88W1AnS3UydUrh8FZWqkOUbP44248wh+dUoVdedEpS1GnrZW0QwzqrWV/rP+WnSL6p3
JfIt0gRwVcIY8cyEAS5yeq/ZhcduM3u01SLqSyEKq5i87C07zZNRr3TcrJnfae2AyXNvuOpUBcGo
S4LCYWSfx32BACKaclOp9IiJ3B7GudAOpJ9oQda+PA2pLeWxnd387vIWs0Gh6fYciRFJrJm3y4L8
QpPCHLRol16ecmUOfErPVqGkBalN6/eJxiNw0BITJ+IsGle9Lcxr0nlfoqsiQ7y7sbP6TmWSgC1l
N4lSLTHtkzzD2MUx4alB7f1jYIEy6tfTtS2HmdAvnKIbf1MfRsA9dPtZc1Wv+Cq5LegMTRlXwujR
spzQvqI5kubpl4u4vzwXNkhIP84nEow5gtmWz4iy6TH6L1caqKQ9sUXPTKOtS+yI/PUVpacnxpQP
cGSwVvXLKu9Y0J0oq2vupbVbAdRmaXToRYQwZTSEaac/+6rzhIG9EcelzeoI6+BVJ8MwRdO/VUcR
kmCH+AYqsnY1hELMEzFB0I4MFSKzV9TcRnKEFPUDMb2Zawk3nA9MZWNyGOzyLGMI/ppAJNvBF5Lc
1xa381nfRWdvf9PSuMOMSK/5JcJAkSRaPGU3nkbeOxlhlglHF49yA+7IQrySPVbduZFAwT33Qovy
UaQ8V5DBId5vRQjPptyx96QQGyuvzEUHsxeiEUNoH6a22ZEV0FcJcPWIg0qAFOxo1LU5xC9klYNd
yeTqLOH/FkgQJ88nvA/wiLdGy53VJDIZn6yzzgGBGU3Qr7pKXMNAR1PO740UUz40jWISTK+qIKVH
3I7SYQCQ4+bWsbezbIUuKAIA3eRZb5XuDJYdL2iM0VniVRRc0WHx/MUUcz41vqzOfY4L5Kjhrqly
bnfC9xYRfCtNE6hLKeEu0SLk/GpXszVHbtljUqGNiP6h8Kbti2GEiaoO5ijX1yHlLrJ0IpYmmXZF
6ARty8wXET8qpduQNlZfFN8whLvktCOFSMJ3yOiNkOAl/521BNUUz1qZksa/295cCG9Y5aPVS8gK
MMisKzqib4i9dz3/cU/aT95esyAgovIfctMbPgCd/gYmHisS9q555M+6ztECwWnc267BVdavIK21
2+ZrA2JHzFs4y4qIU79w+hjz4MfL6IDiJD2pdshQ3CDHexRQs21/6XB9X3HqOKH3cv44Pq2QxUj7
EiZywWJv6PwlJgN7A4xY3BZpeJKl9sy18Z7MYYqSQZN9QYViFQJ7OJNpaphMmumyE2A340lHPOYa
+YvQ4dAqx8+LIE23co+1diQlqgRcrNApzx+XbYpWkVUzvfPALOW6buWSzvOEo+ZaTlyQFd2/Kgv2
5UUcdi4oL1EmNqJMTo0pXqMzMOVQ+8LUD3gpLPPc3ZLnmwgGnQPGop7ZMhrE3sFqNJ29QTJVPrp3
ORY5H5L2fMNXIjDhtec9SZ3gqE34iaKfX/BCeSYRXOZOnAbcayJFf31iWDLFO1EW+GrWAcRUVdq4
CRwsMWip5zqSfcs6YVd6/2TgxuHI0U6RgCxLJ+oGgH1avErLJtphoKBjNgFKaxrHJCJYsFph3UnB
K9gToVuhLH5ODgrMpAS+2SXJBM2RBuuLQh/u3WYPHh4BSz6Xu2m+xvAiMfErbmpku8VXhUZiBApk
XzX//WeqMLyxYnahOPL1JCy7z3mY2YgRMREEe3k763aR77MEm9hhaa13R1EWNeIfWeNzlxzz2CHz
gIW36SKbKnQRAyjxWvOM2RQ/WlMONcibB32JpJ27YCGdsUvRvbiaeaKN73Mjfq8Nx7KO7H5dgx4Z
I8VaoYWTV6Q0xD99xxD4d5ivo01y/daNeZV3GJoqCPDDehoyO9cOhymTBEMlgWQZ0v5oDzJpMUp6
rghxugbU8Z7oK/x7vRU/6dfpy9ORCJ5EYghF7+MJ3y3LQV5JcOsZqTbV7UdAwVcmAzbJyf5JY+Jt
S7jOlIsS2+dPFL22LT9xOhAx2MuH8HLm39Go9f0+FdoaKAwLDDixbrB9yUO26R9a66RNspwohXyz
/mJ9ZnbKWaKQcQYawVevxvUbGFVI7DYxK4D2wtAybDq1CGbj2SgGvKNCqHgq6OrAOG6X7bW/FVm3
Xn7lR2JjB7skfV9W+1ws1d5nLeRjGnfHhwxhwhWiaZbYilYX8ROdJ2KY4yuT5gm/Nf8JMZdIbGmG
KdqfRTl+KEOgUAF/p86HgTxvFtOn4Wlc+0Ix4ifNGmn9sqA03qqAS5f96Rs+d4cW2blzgJ+iP/ap
LyVfa/LQMURV+N9ZTMgd0WwQBKw+uWSNGPjsHdE0VdTyrkLbaxNDuG4MZQGamgmS7zDEUihkm/AZ
+IgMN5zz3yQOu3CjU3j7P2yB56Axgkd39K6ccBfrC3hyBHwJrWxObWT53ic5vtOyixj467+hoqjK
CwlZkXdWzgOKTjAdmnK6i7MaiJcLgMpzDlRZtWr6ucy41Hj0KJHvXyy4W0B1CUBPxbGQ8OaY/Mr2
auyN1KIU/eGmDpV6DuRl78FvdNYSoOFs6S5jFJ/9WMJ9LPGEIQhfwlVLrZtcTmlEVn1PpwGUaZFK
uhoXB60fZcEtr0aU2ijS913tj0LGtERi65uF5yKPFE9Xu+1oSz5ioFJopb3zUAxM6BWWbMs0awwG
Q3neMUtpcYHMdFE/EaJZmf/6dZCJrRih+nvGQOLbbk8wXtYaaHSV0Upc+D3u2msBTgLpzKmR4me4
MTHF2xJj1v/CRi8jANIlNE56AMrjUnSuoGgEgbT3NTwdwaxysiM2GgQTGPu1yXjUGsS7cbZmnF9d
V7BJ2mMOzMkPxGmXDPPRcxQuPDwxwFA1hhTsPqla3WNXfdfc0VQQOYtT3BeLEroq6wy/xceIDHzh
WH4tmeqVwO+0A8w8wIG0ObqH+DWNq6/yOMyjlDc4be36Auvr5P/zY8VybIF7CGAoAPPjBUxVXQf7
vk4Ypp3fjSL9+1i03DgIykAEF7IjI1JPDUYDSspXZfcWUyFVeynFMPzY9yAE3L/VnuDjFnCii03Z
wpGzYwCt6AnBxvgX09wqY1FoQsJQAUMqrp27J490KgDdx9xwE7uYdAbpx68xCAFY+m+RhnR4ExHR
d5elY7FAhrqMmYx/5v8bjxqO5KJQLKxhhHfJey/WDDXeYHLcHch9yIQj9ZlVVuX4uh9bEp07KwK9
numFTmm5GUX/jsfHXVfQjzZJE4UHxY4YGDxjBd5YX8Qj3y7KUtPrySojshfvPpdNd+qytV0ry7jt
6yo8NljKE0hESIMpRtMUPVqa47oX6zrh1WRUPX9cdDCvUKMi58TGtkY9zUMrvfD3sUhVqQXJHoEL
NhTkkztfuWawbN0qAxoTsUq1UmmuE13ulq43HQZpeetnOuBwDV+JPahi4M/zYIrVUuna6lJFvT3l
S8s8MgGBvkpaW5svNwUdzReEFeYXRaf80zmI9d561hMP0q+LsPbBwp2tFGb6/qXcCp1tkTeJHZBn
+pDWix7uWd8kP0nj+iPVBOycQI6Ldmal7O7DVZVH+fJBbAlxDNZYRipM4LjDKSTARYUk49GTEngR
gztwVyyxvFANBVEJU0hTi0H3vqczr7IRVHAPc1sh+hJcqBSFrP98o6Q0ox0iejFVddTsCknh9B91
LTFHu8n1z4RqDNeIKInRDsfjgbEQAq8MNc4Q5POcaHF+Zra3I+MRigOP9SGUEv8lc4yle7u/1Fmr
WGniIWtj91QgUcTajeIHXhPoWipsqCp+7mmn5N3MgPeXQd04qtYD/V/rsl66z/Xesw1Yya4bCxTb
16PUbGn6qkH3/1b23OK9NZQZ4XLGbf8+oMBWcrxuWSl35nnJfcmUP+6OITuAyBy9XHQighVQb9mw
hPy+nCrac7aOJ8qMvXnrsyEp1RvNAbruxkXUThQDUkUYtzWyCj26stkLgkk49tM/021ZFgTMXhFG
dSBhzWXeo5pR47fxT6Dqrv8KPIFdH7hRmfWs5aLtcnYLpXz11mJb6YmTJOipgdoBanM+mK1/wyEb
ot+GYhl04Exi02P+ANrPmiYixf9y7TMDV0ceyNN2D9YdJGUg3/2Q1aOWcRlJ/n9VrxtDEAVqBIjE
isg/h1eSdZVLidIaJ3aounY2t7ecgd0DW0IdYyN5JR2fTmjcZpplwHhb6tyI/sK6Nbt+7Xx1R9ly
AhEi5qRu8TGUNYSqX1BYDUyoCuJFy6ai71z4CCAjmzPVqktCwqYFRgShioG1H4yq3zYuaGbd5c7m
Fjo8m/sO+9lKudj/7F20Zw50q3Vi6AJMz/tKsCHlMFSgm08707jFQZsSnS+MTYgJNrpsqKyF8KZl
Nq0kVJQDIr/wF59NxBJG+u2SXIR1YV4Z8W1FLqcpwUCIq0IpvQFggr09bKF7/jnfXW+xnnGv3kgu
sjyWz/eBPW8MovQHYa8ameJIe3YWfsO8CGt0j88vpwyh5K7zP7h/La/lrkUPv0C3NKBHQZ4eAIgE
i04XgFcxBAet68FDktLAl6r6WPcO6TeaJ8F6x7NS1tL8j5z5x+PD1J+yNcUpayRpOAbzG7DajqSw
FFr7mRvT17tj6eedMtfQvyzsGs0KU6uv63s5UxstJUdQvXAFEAj93TXoNm+tDMYs0QjWOIkRD4O4
pIQ5c5X2QkwMC008guHlQZoB3HJ7+jR0iL3E5qHZO1elZ0aV9dedvAQ+fsGUiOJSHISqQZ+I0IpC
I211UlEo0Qx54ZBdaxJTwxfarF0uWl0/jVBgIfYl1/NZswxTnTSw7bWZ4USHzXG4M8DZKXrU7Ymm
kbZvwXL0kqn/tg8Ij3Da8HBmfsqPTLazm7kyr4qlqWr0hK8FbTPRAUzKUlrMHasQwOCxub1tzwWL
CPtXLll0uG/ZaE668hKJAvlYr+AjI/D0PsafPHGj/aQ+GVVtJJgMqzAAycRoZIVl4GACo7tmTe1q
/mbp3qMK3XcI5YwUXGwSNQ9krWjPy6JjzLAZCWTLfiYZ7afXo0N90QrlBQkQTvAVUrPi9No4A6wD
ZRSn5V/wJbWvrYtfU6/rzr0Ikqd/x8jE/m4K6wdRJqGkUP92j+DAtNeoSdaRd6yYBjBHoA7wn3vx
FV5QDyyVZImQvTClfrTXd2kpkguPZ9xXgcLgBwwAqZtJzDbcm8YcZoF/9YNgC/IvZS/m3IT1wiPm
ck/Inzr32G6bJokWHeLQCoew/QHtjuIZ0lZ9VrUY7wxJLTBfcz40k6xjV8sCk5lW1x6wFnEpyGjE
3Lvat+DCzL5VKEZFb4ZnC7+QsrSM/zYVZAnZfLjI5uDLgBFQnSWfMD9jwmTU7yR2yNf/jQ7hODDS
hutXcJ/Xz97Pwd/AjoV3oyYJSRayCiqOa3b2M+J6gwTpi237YHQM6DFKKlP+JYeb3owcxLrfxClN
cSKa1aYiPPKSmz6wXb9kxpA+2297yMRk818h22oy6TDkNMJCg0ScDob0YtT+Msulpuug8reYD4f0
RoH9t4fFPg8HMmp6KOcyTMWk0QhHt70fk3vhY7NbEHcBktAZhCWc09AV+I4ariE5BH7HIAfcMxYn
qbEsOfmvA9g50XuACuNMAkGVn8zkuAO6KtXtmMoh22oERrZZbFio5V6anO8R9FR8GVZXtksdqPEv
YBfJuOX6qCJkQPehKpSA6ZGr3MuAG3BBQG1tw0X8t0ejLlXLYkAqMg7VbYFnphGoyLeU28YDCCyU
McidH6qtlhgJ+tOhEW7VNEn/ouZG4HSCUMSJyYtGbpDyO2dG6G4Wd5TWFANUkyTsy7wyl6oW8yn0
WHpQAJSyvjgk3q3mWP4FsnBcmh9uh/n9S7mpLUH3HDM88AAB+rqgGyDNeiijOzh2wA6HjhAM6kxC
g1tXSqV6CQ83P86Madvh2cBGFCp11ifl++C2XHnJFifZgk4UOzmsTgkfGAD5uD5XTNLF7LNhyRdZ
NetMLEwqJcYr4BHgvon1mw0H+5q7N31toMk1w/ripAeQfS4ulFEIQHtRs1QgPZtuoqn268g2AQb2
datVdoPDIHk41UhN9k1oVJbUTEoA0jzRiUnIATbeP/WAx5VQNrKwccqBI6Jho8OXugAweKKb0k14
TC2KHi3+R5p9uMC1EWAx4Ezx2xLdyjZkjkybDeFvYzonbExzrJRD8L46uyHuICZOxFJB5qwL6N5i
5wLlXBlc521R7OY8nxrmIH+jNFjsijAYFSIMxHQ0+QIKiYtJrYSEuUx7gZIfWDaoRYXUr4GWxcpV
Fr7MvvpDzmj6LPs0uEaa57uSZ6ziTdsBa9uDmfcUKpZqoHIOO/Ehpu5K0A6qmw/Lh/gU9TskwPEv
qI0WfbW1hOI5PhqNXZjBGyVrtMuBV5pAilgyIja/+Qsgn2uy6szvDUJHKnZ/MiCWxYhh2AuWoXlN
1YJYSTdRrwZvLHnPnAMzHJ8KBul+dwFa1aHwT4PJMFGfKqAK88cb4I271Taw48ZTmZEXENZeqMt1
ma0fgz6RE7eKsmTHc0jNM3bA8FeGodMADUGbOH7c/y3O3QtpCQZ67valgS8a+PFo68sYhXTkmXf7
jQQob+nV/QmEn3d1zBEXB1K+guzFf5eda/+7jrmEzqiiPubEq1dzNs6kAsuSJvP+z6//FHwqfPrq
+kD0sRZ3hksC8i+XSxZ9/7qN7vIClN+xZ5mDxnV/QEqj6J9DSPSX10fM0sCvB9dVdZPAlZUDKjkN
RuPvf75X5nHS1UlE/G6yu7M0KKg07imnQM9tNZP6gd9EGq2UVuNwmZp4Sm8aoR9QtXIe03B3Kf9H
WgSUVRq3bpXchpnigWo4vVNShp0fh2/NiCVwHR86TgtdeNKXtn62u9J9omxYtOHzaEFN012ormU6
qRoknwVvhvGXsgTPaEMBLe5mGwehimV5t4a9RTO0PRubRJak9lskrhDQWpRugiLWxLVgMmJakPP0
fB2bvHFkfZtM1rW8Lyc4aIa1/CFqj6dNqSPNuBk35SktinIVH1DbllDquYTUsGCukA/OJtZxDzrV
OSe9V8FZrD1EZEzHYff/Cp5XaudeyBAdusvY0wZIpsGlh8u2iTrTzkOIHIlBGv8b6yLjZ8Zr7vkW
POElktVduJMowo4+xVIEUFdBOxTMSsO7IJAz6TIjbbJlI9ZyIRd8MvXLn5gXB4l+PyVD7LEMwYbt
8Qsl3hpPyS6miJjpJbkWw0seyf2ii7Eh4d2S+PHcrgW8OiHLeppw3GJARhcu3JbDMQrQYwpoZEjB
esiZyuHImzjH1a3KakHny6kQdSbTil34QRDh0EbG1QU9I0kZHS87jxppbU+GVPzZVwdGaCZfWVFv
Tki6uN0DhyX+bLRF4pty6elLYVqQrJuI+21guPhNIGVtIFjLGpfUNQDyJd+PE2Fl7xhlBBrO3D/t
1xVOHSk9LaPHSE5oJ36QSmgrRflZAheDQZmfFTF2HCHJRFhEtzknYppc3RzYT0BEv20KuYPZmtHp
caHA8MPGLfhhKm+U8PUTwjf3yoRMRf7lNPFI2E5kF6A4bOEyi+6OgG7JShEJszkF0JPSAytlWz8F
LA4g7PHEIbfkhYvfQX1n4VGoegtjbUrdrZAZk0jD58txEaMdwlVi2Yut1NYmjITh7BymtwWd0LE8
ce+S+k8NdtltCiGMxiwcJipIWbyaKI+Nc0ybtsmnymngJMBbECt402npVL29R2bFpKb/BhP0B7SU
t/wcDp/O8wcj25akhOhQvmnSjLiBbpE/j5nqqHeFN5ZV64YZlOfcXNqfWO3iab+niGNit7U9JpqH
kXLdEikT/4fLJBWbXrLi+4ijVtzQKe+2QukJO65kpzyRXqrQ9Hs20Z/ctpyg7LLyNIDFDAjADVAp
FZaJETwE22hp8FpVv57nnTdsfxY+2E3Y/sqFHNtFEikP09YvQayW6H+pmyjxQy4Kulm2SFa5+e3w
oqaFr2e8zE0XCzxJ8oGo8B2DNg53MtVVh12hpDhWGnGLyzfuUG8dQCR+CIHwX9Jfi7BO5VsPYoBY
BJwkslm2PVz1HRXIzKCnrzP6Fq83JcTTQWuR9gxPGJ5+6MKUyysE9jViHwD4Cpy/zQDuD3+4zk3O
8MS1CQ/qoBxUvB7KCHXxodmVsmrnD+ZgAu/E67Lz8iP8mIPjAgQfnN8VRi0Yz+49MsERVl73+pyy
a/Nvs7NvpSQfuEx3iSmAm4Hu8W+CKleRqNanprkALFTOaVQtf5/qIRvuwhj7uIE/McexVHhrbhFu
7fUE5rUjbANsxYdO5IyJDbPCpArBXec0fBCYPDPEz2Ab/F8w/goVZvYjgjoFv2ouS7r6cdpBF5vw
NZY7sUEnSsJoFCuXizsqE0TuGsNxiGpGy/DGHemnbRjfqIuGOnDhOEhJFZca012T2Utk3L9ncXqJ
jTaAZ7lWV9ytFh16LoY9bQ5dvYe9v0XEL9d5R66rltuoF8qxfStXnn2WAQHCzcjan+hJjUmxFzMe
8KcN5J7q/3ibOggaNUqNAcjiuNJrTfDQs+l/3Vqo/RWA8uLko1aXVVdkDqgrVXDg6GUYUtKen+/F
Pn78N8I/6hVba2POuDTnQbzVE99va2eVFLwBrTEq2orXZuqU6OpvGVI5rmFImt6pGkL5u1wpgH1r
zyqq8SCfQuv576GrQ1TzFadEWabR/os9TCDlkPyyq6o0U4JCIqaO4dRWfusjJbgNA/+iDP/5hx6f
luCL6SDM98RD7xXt2oYV8mBqMp+M9xHV1s0MxHAMglDkvvMqq86CcYXlMshKLHoj5MOM8XW1t69t
hhqxeUc0/6UHC41mPjftDvw2NNgMxm3i3vSrBkLq2N3PRNXLrthdui9MlrGsNB42LAtizi04UxBn
+AUh4sQHfkilod4kwdpCBIp/3+dh67TE8Hysl2qGtSy6Qxcf5mMz8/SF7JeBfxGmULKNI4cJU36P
gjxqXjWO3ATNrqD4R5ATQn7kbs5ePydkEG6hRau8HJDAVsM+BzGh5yJ+fYWJ65d6KuPK9BcnLm4i
K2uJmNhdaLQwJ3SVmifrS7fEN3oymLm4kRDt3L6A7bykaKVFHYjLP16FTgaVlu4jxTYzCGO7JoRI
c/XNgcjAuJ/mZ/ADtgjYNkeGUAdf0jEJajPvi8+iXUF7t5pWjphh4rNvmqRE41fMPjHZ8q3jlILn
zHJTvBU/d/T5M0pYwJto5LoGjfWFtE2+almiZbl4Q+HE1MPqSQnzJcJ4PZD9dcUhkE0xepv1gLNh
f56eg+02tZeMmFfUGPZZHFkFB+qdTPdRwWUnR+7dXcif//QThuoom6aGgd37Zwr7D9J3uWXy7eFi
Y6j/Ub0yxKgtbOgGCe4BEOfnThKHDiRR/oDvd5W0MDDhcSwPHKSxMVBYKWWu153BwR+n3E9V5Pzd
/MIXXrSZTZB/e98mLqEulKJzFUwhNvvsmARAq3JFrjyZwWOUdPnuoIhRGk37dK5bd+HvYAiqbK6M
mAkSrqhTjzawbDh4SuCG0JJll6CBgMetar4zgU6KYtPjqYRzELSIBW/kOafda1fWWAsdL8RCRute
ChNeFwM/upyyfyU7XtGlGUjlr7szFvfKC9e77S68V5yCAVVR5T59eUfbI4WWZVhWfb3ykxp+7CgU
xsV2v84fVgyRN33k1sGUF/CUegdRO6f6eJXKXNnxD/OlnjUwRS4zt5erX9vHQdNqy+SMGtBh7t/J
8L5BJmpF44RpHh88RinJIp7fIPrSq5J/sJrBFUxQCM0IBgcsjy7JODRhb+jJ8S1lhSM71TYC/P78
YAs5/FH5daNBIIKfkssFwxSmf/r5xbbZs0z9KSmy1hiPW2sUPx3tTJwaMaxTD9lD5K8MbGdFlxUN
0akUC+CwT1RssHFGIKLn3R+hy0/L13PsrtsnoSIRuFGe2XFOqI3KIGGIKMxZZ0PW1cG0cr9mDI0j
7Ufn/WhS9UQqUIBgBx9CXH0TGPnsPnRVPCtWMtK/RbX5dEWSHYi0NN0u874ORDOzA+/bzRiydzG3
Vx/47BpCUmIp117ynipMVUtHVD5zGtmcjUFZhdhLkV2KSQHt7Xoo8zSKqF10bOdIKBZQVIIF5YVx
EmrmymYvvZFlYnIkD+0CfDkyu/oyHceRm8PX7A3K9Cx4Ntz188pJzbqz4S2YP5vLr0mHExAKg3C1
zgeumCm7WdvtvR0oYb2YeE36zJSOSNa7TCcMpK7n2x1mlDwOaWqoRjATXmF4KCFoJzxxtrs+N7vO
mmEUQms08ipbo9VtOHJyl6q/InKhZ2AuHa+7Q2Y8InBOb4j3t3IDW55ztd6wZvaVvepclM3PkuJ1
JAIYj8ELOA/2EOFKI08BnpIWHWsdiSzqMONJhTD3aatA8IZHcuPFI/vgJoB+7VTE+mXL8oRD8OlP
dzIDHg62+HktKmavxE2QsWEcgmYePsk1B+2Kiz3ZHoSqKkGIeoumXLYexJSDKXqgg9jO8EqjC3a3
CApg07Npwelg1EUJFDZ1PDYFRAf0NCYx/wiuUqRpkvZzJMMMH6Okj0apSqqtv8N/PFylTXZCL2wG
dhWIjXvC+wG2T2bBaPcWjsD5TdVSPN4ZfgRKzY1TROV1SIGK5VY9WIsACwIOHl7O6eXht6HqV80i
tN5UaOI4tciQrHKe8LUU/pcoPov20+Dkxt8nnN+yrPI9apuJ5u1mOOTiCrah8qFITVv+SyxuWziH
yO7s2GDeZmd1quJ8nQ7DS8vLHflnI0NK3ufZxF2KdDRJ/5V3i768LyiRxMXrsCUt9HIpM5UKNCli
qyEo/puFw+XoJWsTEh4ZDwOu2/x4vS6UqXAcrj2Bqw9MxPeNFUk8z2A1/aIr3Ss7ckoxCNunQP8N
8g6D9m7fPyfYZSYZ7qJ7J8Aqwi50Sy/WN3usM/S9MZJLtc/+ku8ysSupbQIk0L54d+n+6cRJpDUA
EM5m47nlCsDl6Jjob0qbfQHIyD/emWOdeWJznTmSmqyeH3M8w34FiLyciIxk5pK8x+gCsNgkQ4bv
7bosLXYTs5IDd72IlC4Z831ja/j6oPu0/Aa+MBB85NFlridkLMif8xpFWTJE/uprmsF1XaPQpFda
66/WZKysFi1tTIhjlst07ymzh13nXNxM0LtJfKnsQTmftU6NmzGEb0oTIz58dr1ileRL9y18WLOu
ezK8ynonir9Aosw/DVTqgCkl0tN1RP+q4e11VGC29E3pN9MF1Bl1sE8uf+BU3QZWr/hU6U5+Ehv1
Zh3wgNtaNMfskfOv7ysNLqbDkoQE3cdoQ6Oyx8ociSM0dvacLkZxh+NudAD8XZ4ELNKunL1qeJo0
m8wKhZzZrAl9LKufRpUr9mu9AItQqYi2oDoXrCmgIC4a1ZYI1PSzkNVtMiRCrgeOCqD0L9Zc1Kpr
Bp53bEuGnrP+erDByGYOGoL1LXxEOBCfGo73f6TKtWAuRAeTp3afq8ERMNa8Ctyjogcu2Gq4gZJf
2VbpW1mEiJ6bQ+niKUWYZVdO6jViztergC4KoD3LIe/Jed+QW36Lt2AwIiOMCXcJNLE+PUx+DBdN
w+4urd3R3Nr1n5+dJrbS98PqiQobXAef8eYQ5hO1IBWYBcF2lzDvqBXWhmSTfke7SSxCxZmLoaDo
7Up+p3oLKdYaPFPnI+tlS/Tu8Ro8svk/3kSK2R6EXUnCb0+8dj0DUhR0BSqJ3feVI7bcrfGzIt9a
e6sav3VguniXAKpTTQWv4t+djqzHf73F7l1rHDPFZTJV3CEiAP3hP8uKcjeBi518cniTu83ap+D/
q1jJyc3RPq+bD3SmDhPo1dEsQ6BmWOAc/EP06RlNed+zVOMlrXQ80oKrczl3GFOrXJVHcPAVsIn0
9CPYT+0tcWbkGlRu04up9BfZAJI/slyQHA+BUEJ//Lh2tzz+FVTLUPVw3Ga+fE8DCBJRj8yad0tx
ZO/9CB7kMhDfHR/4/z62ytLWjF3LGubRtr1DoCxJSPU9z7Qq4+sTL1mbD3hXZ8sCiNuO9+ikghCP
rJLhm6qHZqJIARAkBIFnqyiY9lOY7UqZ1mDHVSnIrtLzDKL0+nEDjBK6u0pg/GgP3rETEV5rwF/C
KDPv96eDtTJG9vNcFjYhlW4wzQew1L7+fdN6clYkoHksRlXjvV1ITI4GiKnTdZvncwx8YmDRqJNE
0DtREPkgFgU7MvVDzRsX4ZqtysBg7iwBWu3qoT87ytZxDPNV2tylzMnC+6gPp3bOT8FZ5L0fmV3p
FbDqmL8Yh9guBn6oaBVRVKunijgFhktG0R6whC6o8dc/IoMIyO/bf0OyTeePkTc/UiPU1gFe8SDz
j4OyM+CjsxXpxGPW7a77V/MJ+I4TK2zP/1yfJS1/bHRF2+qHjNABjfgFD9AimKhLz1yCjF1kVtXX
/Hqa6IdfWuRvZ8BNFBkVNiUIgSaZLjc7B9z80QZ1qbzhtd76ojh++NUc9p67991QCKuR8w/61ukQ
d8IF2emZY3k79NNiYnBghA2FmD642O2KjqFxeqKqgzVBHkffyucMn5WZ2p85Uz8GlAQqKlblHZLM
eQU9FlCyR9eKm4X9QGWipUn5nprNeXU85B00dg6Qs/EIkRTO+Yd+xEnOScLNeB9phoeL0m6ie6fz
zkPVMchLnMWGCj7FVPhFNPEDC/6gmGDIPANH3k981qz74IG6CifmjA/DcSVR0IpsvGz7Z4S9mMOB
C44nlXX5oje6nTI+Ln/TzLDaNpbT7czYp/dNVDVDocfPLNwA4wLiZYv8YM8zuo5SjcPvaYajM6Z7
NYG+jnSlUSSGx7dLf2ixg5A5D70yPNUtSbBZRyxXiHF7xS1uVsZu7JuR6K6p6ywNd5ctKjXiYlsE
2YBaU0mU/CbO1UX3hV1lk084C19+bFcHmBt9RSJ/VrrKqaedJhhWNQJXWSaQHQN3fMjZkU/V20Vn
EwG8CpVLBvvzyL971KaloDd89C8Xe5psy+kq+UhzK07sNjOYJWcW7j49fMBFyL56Z6fLcgmjN0co
FZYhpFelJ9C0m+zRH6IOm3upRlNlVzP9PQSeW4RUZQgqIAkEhRFQQsnEXeCOrutffeSnbyZuPe4w
5kp0zFN7yckOvlsID+QI7fBOOnhkzY6AyeL3l5pdnL3NSfP6/LuEhzDOKwK+JcOqWbOBl5ddsHLE
SExOP3AAm+Hf252SMTwmzhY1Ynd+4rhFzjj02wiDTI+NW2cFXt9N5KRjTL+pNS+9tJk+m2vgxaFf
i31i6UHwXI3kd0eJXoHLWldIMu1ovzTeEVCfS1ubBeCFDeHI0FSlqxKECJZEr+JKfcbqlGiZK66V
x3tGobAhoD+NgyEPLyIVZe4poh8KIiEBmMY6/VxNdmclL95MGRoihYduW4Tq9vkEkFQEZZq1fou3
qtU02oY8TqCWYn7dfiaj7vhmH1mQUKXe/qp5RP0npdfcrsfPveYNKjTKlDXTNLW9xFVsUcn5dQ3N
P3w9XgE/zFuUCtctURDXUCnG9XdmtcRUCmIvxiFXElhbpx5+xBvwiqHvN4iAhBDbsRS4TgcAxGmy
T0GZ0pqsw/gbQrzhDIy59dcsZzwIzZB0E56qpdRjwt4zAJ8E+82wZpvXleQuWhKoilJTJWYmavxR
ipK4a8dUUM1AC7945Tg3UyN5uY4KcmHDS58X6BCNOLjlFnIBXwDEIUXLIUvSmDRUAEI7PomXeVzQ
6qe3PmWHjbJ9kJvaQLvM82btAPDzImhIJjd9pk4VzFmhA+j6E3z0NIvjxkGq4twC19EsfT+OPBd7
0nEDSh4kakjlZFrLc8Lrg1H2kcxlvvHaA2MaGfjfXWXTTL35qi8VpgHUX7pWYxOxvVfJ+bAGmPc+
omWtNdGQai9FpSOz/yHQNeVhc7O26ZnJ0XqaxZmFbtPvrQuxeKHB0nKkqqcnQKQN/+41zv5C5lnx
Ak3K7XLazET+Uq7GYqauWjK2c9EvLufU8mZcsEIPH5uR0HfBisECZaas1WhrO3B8xYEed6E95mha
Q2cmkZnkWUABPE3ye4P6wf8SpE6Y2KfMoFSmBu+X2Gq08whm2fwpo0iQtPX9E8HMH6hOr5KrRToy
HGSLujpZFwfZHajKsxVS3/VF7eQ38/w7QsqjUCjCczId5iNxETqvG5tMlQlxk61/e2PpW36jOy69
9W1wIlrvE85VtKYHsmcoSQpQOOPzMl+fWv7Re6a+dSgAAQpxRMfHy3bL43Vn12Prk0Bf+9pr1ZrZ
DpUL+JmIK37deHVsIzgSqy1PkCnF3+e2LHAgbelRRkTvZmakvCAk3HieJhG9pxXJIxZdnDXh5oGf
NMz+R7csyaYfFwXrSx9dctSduwJoikGr2psLDE/NXUSkPmubeU7/l+sg2fIzsCYTJYEmu5b8vr36
1ucJk2eczrm/AVvNl5CynjJVH5ZfWkfQgB85UKUTpZt74YiLv8nlNyN81q2gHV+iRLgVOYI5mXbG
ZtXOxFCM0ETPsSDrbpLuuqFw/KEyBzJRj9uIrzZ6q+KE7F2s1mx5cGDzfu0Eu2pM64olTBjCeIQU
v1OItJjdwAWog/NS9aWmR9UwUYm1J6AkcNbZju4exGyo5wSIqYScmROB4VT1uTEvlvIKDCxZDEY5
esouXFJFLc+bu7IlRXNGSyvsnYG9ThwOup1+3WmEs2Ee0blx9qc5RV5v7rck56npM51KK1NBqwPl
Bozlonw1jyMmhGCgIm2hNtYSTgALnvfjqviVsxyQwLmj9MQ0kHFj3LQ6xdUX1Ycwl7rfWr94rgqz
wFo96gbel5+8zY67kojViqYcPqhduAsACdzDxt+Sgn++8dHDCQXMAxz2yoMUfocZr9rBVlxurjXS
kLr1LO28m2WuJX/bIkS+si+0u8jmCe3Qjf1cLjudvaY3uS4ps8/RejgW+zQceqzsS8BI2T/8Zkq9
sEvNE1OxRuCNAQatgZSQ/cbHqkaHk2TXEERKUDWI50bgGr8/h68WyCFiOzkSCpT3wvkFyGwJDiRC
vkGVxYE04hmG3Bol61+ZjERDEWzRiiWSPj18+RCFhQhdlawQ8OHYIAhITh4arYMMcLUOW2Rn0Qct
beT2uZVF6plL0YWQY3SL5XBCqETe3uaMxePKDXJd8/QUvEEnc47mWzx3nFLrYemIt5vcA3RFiFKS
AD1MMO1ABWcM7OUhzAZ3vAX3mh+hpvZHpinSnpq2aTaw20Fm/jc2lHhADZH4aDURQTFxR7zIbvrG
Hz1nKp7gVsGsHb9X0L7rQDQ68u80yDvf72SwvwnsLY1NXwRzMyYXD7/nYzWH6SnyapCOFgS0+p0Y
u3aH4/4Co1ZxJUGMr9ZsMUIY3Y3l+kCroSMN1Jtj0WrNJDxLWwkQAXVLCwEbFGx7A0wudtqjKo0p
bbr04juZYE10phQ/T23bDG6IVIMISks3C5Ze0CJfEQr4s0Eg9LyErrm/5O+ryPUa19UPFLJK6aQo
Ed0MLkgxT3ArSYVpH9a88Eew1cTVSq78BmGqe3jBl6kGahDcoNLJIOmGLcrWIw/+Q+Tabj9q83y4
Xa20BpsHi8vk5N80OBQUsNtIh7p4cWJJyz2PqvnnAO/w/A4iKydccRKQAP5jg1lMIUnHYNxBZ3Tr
IV7ZZ3IbWIZVfa0mzAgfMuq0IHtNPdqqa83vP4FUrPRrTEh7WpF2gt6J3piQhwqasyKwa5n867Ty
pDapKx0EX6rKcVVVa4LoNL8ahnRwIDIPenPK701DOGpWiq4f9Z0tpdQg2zZSTrGmnc9qKAP12MDw
x0i79VgCXbCU1VWbqVf405F+sJPR4Dw6xhn6bQFhdv/3JtlCHI3mnaJL+PvaD5Qb0sA8YQ9K4GWp
uV00PuzPthg+hFx7/fvYUekj2innWDajKJe9qQqJKBIVRP9spusHeVImLi0cjdDFzc51ElWK9R1b
WPeZba0nALQIuiWqD9EdvZPCfWDNfECRLFrBIsGkwH0KY9l97avzS4bObFnbrkZxEf3MF6AxC54J
JhVH7q2GP9C3WzbsPQtpTswRVEVbkCjXdwfqc8evMlwmEDWHA4ajrxKZ8UGpJR6IxD+Vxt3JmYlE
MLE4++1F5+momlXFhwnBy+jdC/3T9PVYB5ESosAdHTxh3Bhzu1+pnbraheCI+tGh0uP7LUb5TDWT
GCSpX1ouCYm2iJoObEEk+ofSh/NYp3Ngt2JmbVdZiZHJRp6fWKRqiXhW2bS3xaC5dhA8PoiwYuqs
y3bb01LrAG3m4q0QX26jbI0KX0BO036jZIkn+r36xOsrvolJ5S4FshCRuYsDQmQP6qCp91rjPCxF
KsyMe30/LpDDqM4K6uFZmCMsQdQVvRDQStxGd08LIlAFC5Q6i2DsHSJCvHXSP/Ol3gSDtYjd0GCa
k5x4uutlKWQ+ec003OdYCHQvZtMVl+MB6B1aP9bRTvL7db9kgb5ybUSpbUtYOHGLti17cVaV1euC
P2pOY8DtaFRcMk9+qmuJ0Hp4aVY6e6RmOx69mD8ZHIz+v403oJqT5c9DC5w79XpKFrd9LBOtLIUW
8uGMzMTZMnKJ7zzRdIIDEr26c4FLeHs080UhN9lLMzM9kBY+sgX179QMdl2y7FtbHRTSkqGDlzEK
t2iWERaGJu29ounnWFa3n3YdyXsqdEc4gmNu6lGiSxYj+tqL1tVwRD4eDyP6qi8wIrOkUOMO6WDt
d0yq6oeWUonPrAQuZsullWyXjkBmx7xvvdCLFtpD4mbAGJL0Kmimr/9zrvoBIU7zc01/7TF2Cg8I
lz00EPNvHzYdDoT6+Z38e56U3qDxmAroY6p5cweu3ZV6L99GNFGjximsJHNwN+3t46/m+nPxn3as
pndfOLXFgVVWyw7PjDZ6/HCchjCHMc8eF7AdoZHumkP5B+vTKEPJUtnV1pRqnZPG8va6E5lmdGib
e4ENAE1GkUv11JiYwvSfxRhzqTMq1lIoyw0Z6JIgsTZOt+CzJ5uuQDLDF2BW+ggqeGIzVJwCjF9C
IxEdktVjZu3RDkVqde7qGmz4Gea/wZMEYNxDK//73VmZvCMQyblSVFdWzFXkagAMjN8xglfRCVTB
5CVRo3uM2qolTMdwxB5JdxuOCSi5AaKUKEUEQWfGiHDp/mk1m9tsJqnsG8PHXh8blevwddNlivbM
upN75VsCQiitGabMoQZBS+rcEtWGFEnE5Oh0blhJuxaotepsl0AEHSaviDXiz2Tu24Jn2u6VD3aK
403UhY08jtbYUDaNa7sMA/ZedHA8g/hVa7igAehcZRrgh4jnoXutjTyHLKJjt5DA0KCSpXMBErZ2
MqI8sZNYMMVjL5ZQ7327KdpTn56fN9f79HxX1/nuuKWXNxyH22FSz+V5DM70LUii44Wn8YrA4IAe
llDHUKtY/GfMGuiAOOvygl00/w2BZjoHxLwdCis4N+YXUk+ekjdkByZoCv1e7ye4FAJymMesudO/
LApQHT8u/OLdNcSKvxnKi2+oBeimqNJsrrwg/xor4U+HLdJ4ydo3FWPSkdWd/twxlRldviMwcVWG
RvfDwqsEXYgL6DNb10FfX6TwuletF0uiQLfpiuY82JlIc98aOrsszFS/2af7xOZ4/LD+0mJvEsPX
CircaumJiVCkvyEldTk9b5RTNT4weqklWTsrO8sSR/bOKeE/48BdW3p+dp7yThhmDWY6iASphowS
YmfhFyQrXV70jRlKumrdKjSK1ka+WtQzQeR3A3cJey1wBSEHF1kVzaAudMoBYeh5pk/uMr84jZU2
80qz4KfI0QpXYC1//hA09PCetfyCAsCUMgfdO595GgiVECuPczF3dDgF0/wLpAbGXNQPwlsykrfI
rzgHyg31fz+mVgU2wuDKz3hhGf62eR19So2kp9Yj00ejrdQR6sFJDV4LgisvA9p3BemiZ+VG0/qU
7im2G0LTIdk0Dv6AvK2wOTWM2fUFFKPY+WQBTGQj6yFLbp1f7qhJFoFstUn6q1r42JPDu6J1R1y8
rLccrDcYbjles9PR1gHu7V4VS3sqEkOt1u9360i53bdkAlXQZaEdK7PE+A8/hpoldb4AAhXPOr6J
lA0hijGZFI82X8jsj+rOlqgXU0J8CPXRrUjVf5kzS7mIE8FnJDlX+ScKwJpur3k+PuhK/TXwB2mQ
WIuaRdivY+TcuedpPQ+ewgWH4XKyGyAn+o8OvLUhOWA4rv1uf238UJZqK/TWtoADamrjn/otvra2
tAKVKh/eawzmqwcdHo1mroOcHT3djrseA+31kW3zoqOCOwgNlW5ll94JyhPv3ITX2JpklRYQxDgo
F7ZqHYN8Xm8JW0CXW4WCP7rKh0JihEulKPWjIQtgLHcxVikJBSD/FlyO7Dsu6AyHSIcT0J/BQCLx
dmSA2WiUWp8cn+X+zBOEd20E45127CV3TdcRH8o51ZdYQqXBi7vXzrQvw6mY5uPjCAdwst8xDCMW
1XB6Fq9iBlzB+cxYJFZtwueekysQBC5Glp+zCyLDqH30/6032u/YD2pekQTj0OBzgKVf8r56mpu1
sJZOh5+xZxyW/qIHqS90Fik9uYJjaSWOH5S8hiMPHRGtV8rYpiP72OA4l+BbSbNEhUYE3yulKfmF
9W09D3q0DWmEB/3xWbcG7LkU4evaDwD7i3U1yexKcu88cml8sKL0sV+VBSredyLslpgL3X9cDYBG
CS2MTccOsVVgEQoZ/RGG2tzfX959eIAfjgAyfKMIraVwrCS5oTUvCWwKFFxG9Dblt18Ed30xNbTJ
Ge9HyohfK/0BSBPE0qF8f7H63RBs3dH2aWAL383ZxxDPHwvjVaVXhlKiiJqD3bAeBq9G9fRyNm3w
Ayz+LV5q9lU0QupOVz5oujSvKo6fPFQo7sJlA/Y9pNkg3SGu7gfrGbNuQT6coq/YlRhJ/7h+VNlu
+GBQ0a8M4tLkSBlswxIMUaLvHOZluoo6yctejpaVz8P1TdlpFX7mzgfWhfvD/wl8Ixq33qLpV3Re
7nb2Vg04DFKUjqiskPWaKg0yzBcfkKdaoLU4daFLARMvqr2ee114k30BmFzUfVmAlwwsk1wOBmne
v1UWD6i0YvpANqvZVUFy6ufwBZ1pvHe0os050nhDqSQ3HZqg15knAseE9vfPe8dUWuQkwC4dVWs7
fVS4VAZ5TkUkg4YWdirza76B/FmmwUco/hMzh36tWQFfGyfE2jhLNg/cnZnN1cdmR8hiPrIDJByi
lJcmQJgqmdzrTMWXDbbOoRDnxHDkkRxic2L/yYU69TOlFoBUcJfDrwKq2fTWJQYmYPsXF6XnTVrd
nA4/upam/2lTcfmF2MnaReYyhrcQROzf9+jfWp7mlTWZzacwaWITrRjBj0Tc2PjsPQBziRGNiwOS
wtltfEh60YCimZsvq8fWdKIVJGMi5egnM2y2/nvhDZjGMtO2B1WMfKz9i/DRAZomsTAMcIxz7Ygo
BGfUHN1G0qrq/6/M/3ge0qBegCiW6eaLGl/8d1OgtbN1K3hynkrs4w3ZRTvSJmEAj7ClPhfvtpmu
IunxtYvl4eInIQPH3VCOEaIvFGY2HKG2Vf9UOP6En1rvawn/YuOdBFPmF75eh7WXl7JV0xQRbyQA
Jrojh4c2bHfYZ7sGFr+mxMPF4wcN5Th9IwKXk3Lm+v/zIo45nZv/pf2+ZL5A01PojK+YAFpK7SsT
UTuBt/0K2gpyPCnQIspvXRWsTByUU6gotfxn9dKPGNFGjTG7kBr13Rt4LzlPyWk9oZHAfh6lJphM
2GWZ20/a5PMJDja3NkvPXO39igJBg0VpO7hLDzQaxbNbhwAnOY2PMBdOVNxWoSCLs6l9Lw4CwH8o
BUkv8kfbFxq7avH3U0n5zfo44bOZ0DliKAvVP76jjGuMAV0SKXUGKozXNyvla84j2IGjaeLzVvOu
i8bOWWaXG38wKlrXAplBMruIi5v3/UjbUn8VRKPngYSPp/2AMGACYUkIs7WlDEz0AONknmICWiyz
gBrFn4nCr6i5lBsHfqgJlHaami4vfOMhVRsAlzZTECiKQ3I1uJO44unlGWz/YK0DlrB7FWKuwZZN
EANdQKikHUjafkHuyiGZtEK3cdT7HvP07tRqOsSkGDCMQwB/85B3pYHgTncftEmNcbNJHZ0VSpnp
jRZu9+unO4xRpFSPSO1mymxFQ5WPqH5CbzB5tToOJn4earUzSh5aBsFV+0TOa1olkSuxS9WsIs0e
ENuZsonAGZeYH1N98nZTsFwSFaWsNX1ID+NwM7zz+Getlpf4bID7HjyYGN+V7AR8eb53emPkmRa9
ND7qdioy2vIs7t47xRp2hYZiaW1VF93kKFs7QCx9mdJZ/B/Bwm43j8GkwHhfQcTHvqxZ4pvG2E7v
RwRhyHLlyixjMebJz/nPxfKorKcHDXmBa8johtSW1jJYNvq75h44SiU7oJ1uJxEQr8EquCu53VgA
LWo2C9EOqnYCJaLzhUJ6uTRkO70b0kOpLxHB25rViSFpBqcZfOKju5qV5cFc9dTmmU+bSGEoPPRa
2wZqf7o/pDZpSdqxXlp9rm+3wug6G3JCvdLUmBeaWm+rlnzLWcHLm024+ZJbpIRF0Pdlhr/AqG+E
5bimoEnYdDKuMjJ7P/O/0zQ9FyxZYx225p59W1DwO+wzOQc7dPkDe0k5x0/Q+b9r2do06XJRVnbJ
bqp0EWNVeBd9T1SbM4TMOjCVI84r+ufsStj27KGThwNXuSjuZK0fusZaog43WV6c/Oq6/q2LJmL0
qxld64vJIvXxehq4THcb5J4+dv2XOuZfHaOdPlwL5Zb/vIZ7aDwaqlauHBJTNC1OhQk4yIWjC1op
5a4rJp1IQ9H4JFaS0TERh9t5MP+MI3VRu37c5A5fOI/TT+M3y2ZnUGqJsumlhPGZokRb7QjDl+57
t02f7TM9WIeo0dRaLoISqaI+VOmuAsgpmrfElYR7nehdM52aXUOAeY1Bwj7lp7wkha+mg8HRs5Z8
hqJNgME/FKp4I+lt47Sfjb2BUJFpqiyhG9rd7wfvVir+vQMMMnv6VvSJ73QdLhztQVUoO579E4aD
Jo+uyGQ2Bfp1gquE1JNRwJc5V5+hvsl5RjoFsPiFM9UF4UPCSVlW6MPwVM42MNnQueGs7KlFFDPw
QHHVq/8EmNgtVU0ZVB5SYI4k2SOdSIyQeWiMypZLMxlWP0fxXM0d04a4SvvJfNx01l8QlfLJ3Zt2
wnL9FhX6eHAHEY+6+8QMljBEpqllYJDVgOBYElFsO0utQ/38eZoGnNmiL7PpEY+qGEujDAFhNjdH
e4yxHKnVNSmVhREtWcQReOa+ikYlaoIXwof3W3c5t+ZlAA0D1eQIgjLMxv2F9VgjZOU5QaeFzImm
mC9rGUomjtcuFKPuXMfngz7GgJItKUGKD0MUrgqmxxOYb1RPTZgWB4HWgFsOGZoPZCF2CkT0elTO
RsPowClh5UYOTZkBNg3mnv4VXWzDnl0WaKj+PUYvlJ+fqcct2nuVzyt9MlyR9pdfuMMn+dafHz5Q
hHj1hFmadtTPNiBJbyJ0vvuXo36mj7JM/C4MmafOL7cmsrgDuU9U+42gp6lM83LPs2xPFec6PmCE
b5Q9P53cEt7h6hTRVA5TnsYrz8AluVUDs/K0/fQScwsPbVYeIVY5WR17uTbfvJYVL5pCGdA1n4HQ
biVFUOTnMtKdizwhfdZoctm8UaTyzIeWskXrm+9r4Z7eD0RogSatEZiupEP7zseJP9Z47sQi+gva
IJtfgSHvDj7I4HDTDGaoCBO0Z4Op9cJZuKvq6rSqUgzf0mIC4yMXPAcDkjDB4sc4/uVuLu8P3+W6
RUqLtP57mBw+nqovNLPG5M+mON6TsCbd8iObcCEjBe8z9nKvEpxLbnxI49umq8ApvAr/kqtTAEoM
XxjrnF4zGoKV3TYGFEsY4tukGBW7o3pZNTPNCok6VgseXKNRq4Z3urHAnMJyjtSOUmqNL2oWvx7Q
Tgkt0jDMwtOjExLQ8dbx4o/iCWP+QhY/TP4/Szrb6rOmUd8nWKlRBNrhfobW9NNs3zpKLezTJDrI
iKMFH9itmlahd+rivvmLT0pGjLt1hBGDmZcnNOQKYgXh4XMQLCpInrwdNxGsfl4YPA1PqiGZsKJr
7FWkOH7EdSMnlHbMp3IT/MsnYvCY8Rbtjuwu0i2+RQAR1WOdPr4tP4+dQtgNHz+bYo0bBQKF+s/z
ipmc/yaBPyCVJVVOdtLp6eH0Rehl26rsdpxM9N7+ALzihnZ/p+3Ab18UIn3RRBltdAE9xR0EUuMY
tTOf7NWCnASjNzGJSj3hlJKbh4WFWsTmPOSkTs25G/z32MtszMWcrwZ+yycSkSjyrgU7t6r6QZOn
DxYezba1UHNGYN56ut1liDR/Tb6BzC+KrLg7DEGqV2zU8MrKBZ+vFSp2qjdUHGlKidMLFhWRy+lL
Mxbk5iiTJMjEnyjivg7fcNXIs8xn/CPHZPtqUxj7Yctnpynlkv/6m21d9k83hIvBBQOaY85HdB6E
3DetjlQVb2x0s5qPZ/TmbQe/6/LWOClNScaDMOwcDWXc3aTIwQWQJFFi7uLytio2Ou9Fn+ORtwDB
Bih+Qmt6hV6YcmnQa+IT/0XZyChNuhXr4JO0I9n+Am9sSYi9k0ZknNXujJDDTDmSe9iy84065Nhg
q6Vohn/G60HxYOHb9rrnO+zW3H5JLomPMEkSpXiYdMwO1mAZs5nUTRPgdRoCAAzrEFrUOBRNQZ3v
AWbqRyDXWS05U0gQrMgnv188H1h9ASOeDohWOUyiwh7B7l85S9aURWJcx6XoJKRWtoyUbydmeJnm
CwqAoVPxyMhNOeUJPSMAUrKHIZo+w/mTJrDD7hPPUl1GikORod2jzmRSEzen91dnbHHEQewi3qgj
h/554iDeFBcZcF7XMhzhLEbcy138oXGFFTZmwQKmrezJPvzZ3k2TWY58JiDQLgtur/jShKmjPsO6
C7yT47aNlq7nBCkTvo+PC76Q8CCgTiTzBJ3g9K4/liOdGSK1SXfQlKXWQJApZjqMKFRwYGC8TW/B
7Y6UvNFm4vgUy/pVGfwX2oJTvPpveGf1w2glMmHBbPJyhIc/zVQiZKNvDKeV6JFO8UmFPd9+w3tY
TSVl1V95G9MUwmsR/DdUiPjuLNoe1zIg1vUr8y6M+OjaFI6GbZd9n1Xoh37SpYrEhD6N2oYrCCI3
bhLz0HTlnoCbB8ulWLwc/gaVIAYFaR8d9vdA3rMBNho5rsSXSS0FGLzP0APOdh1l+nFK5Uo/plaX
B9el18OGtW+ugygW9bx87qApiKItm3+Ab6J8iLhpbKPdL1qXecJZMDti0XyVKHGlb7nRrSehW1Hq
qKJns4gHzpxWUE5TqCM+L+tpM+ekTkooAiIpzImuTGLvpEdpv7evg/xpYyxFFig2YMNJSlXV/TLm
7NfNXEkMK7T+JoZdNuB23mw6BaDvk++iDzIkhDkVWgu0CkwfQ9JFRGsLpbJKK10vv4e78YST6m/9
MFjUTo2wsS4qlCHvZ5Y4OVJZA4JG4dE7y3L37I+cZkJlmEkJM+lF8w4cHCf0QNtWLD30TYmgUA4W
yf0dH0swOuzP23x9WI0nLdiHBvivoVl96GK+KV9MAssUWEeW1YPsjwHdbreuWuIQkykRM2sPCgQ6
5sI9x7fALXKDbCFb2GShPQigcyRhlR+8gatHq2So2kYzxDHqKvyVV39Qzt1C7IgtSMAdTJFyUiUg
0bGeZDrgFJCD+Zj2fYYbRTdFmPIwNUZKTl1Gv6cKQ44rfKXrHJYaal5wALEGMLjdi/uyUa/l6SPa
FgZssfLuBQKiPQFXwPvoAAGkklxD1Hu0CKdqfTK3RNEl6eo/HpPncOSMpomm1SqYmeV3Bt4J6QFJ
tg7WRXWBe4euLc2wjiFPTXopBbimzqk3NOw6fHyjzbaOn2OYJsCCMa+Cswjape+Dr1omCFNkLwB3
hWRgoXiyiRQeboH/3lCzXYZ+i+kqQN2+uHyY1JjZ8NWGlMM5ay1QxLHn/P/FfP8EUkIOQn61ioV7
nX5p7gcTcra+pDxSaHLnbwYbd4OvhHYZpqc+sjPTkCa+qv2Vlo6PSaTrwS6rjBKs0FcRGJmjBt9t
7c5hxmKq3uHN44AW1A2AfG0GwEdNB5PEkJrHCW7XGvlkTicIncGrZMT8ljt200u90w4My0ALg0bl
QBQC0O9IvTyiJZGYyGYW28MQ34gNNjtXPCGhmouFuC0Xj6dJYOKXcjwl7M0MtoEK0wDuUguSzWzh
1VSbta97vjZi8NnfhK/ILCUpYk+jSWTxkX3n79Pivev5DNPdRyJn8mQT7j1fFL0JhtPjQt1sdhLI
AjWpAIdgbd6IpbUsyO6jLV6neLOKrdNt06xd5oFEnwjKYZDx4dWT+w2WZu9u3Hs4DMlmEv+V2bKo
8/nQBc9H8XOEIo5OhR5271zIU/OVHr1NkToivJvTGTCdS2bBq0qWmlq+hgVnMJdVRv0K7TUgVpMQ
m92aDvOanNXHtfGXRF0Arpk6I9+SSrA3G2mqqr2n6v0O9GDzBXNxPKgjyICtOzq9CDEFdnPAwZ6e
fcC4HREz0Y57Uyze5FpgnUuD5l5WNEYtAvI+cy1V/LXi5qYXksmoSJNo3HA/3X77SDUKZIVKK+R2
9tQaA8QSoXpYGB3ruAbxWPpjaLbyiQWpN/fmxEOq10mDBFBogs+O4EGwRTBSwZXZNAwWrspBl7g/
U3Gu30IRA0YqqcutAlvoNX04NyJ5KMMG0lohsKv3JQUS3Gf+C0gzZoqQK2IhuKsiluiOtCMeo3pj
s1ovMrkqrQsvDB0jQNC5Kuc320NAXYa1aPXKAAIELyArMYagw2pOOGQGhpvTpbBUspEZXQPT3kLd
6bjWqgG3kQ4ZYgAhqf8kK1HRN/P8yvPGCpPDaKhCAJ9mO52L56n7I70GLn4Q/Mi20SiYXY4dYdex
2jbUGVFahypkdLXzVxJ7zJ4y1DC4dQxoWO8WAy9MVCNCcl7ir1eTl4kj4fe7O03crZc0wKI3KWfs
5AqaAaVY9ipYdqjUc8Fz6jHIcVIJ+Tq7OUx1Uk1s1eMz+CIQq93gGZtnqJVhNbN3A5jobRGoPVzn
K6l9b8qtMjSwDxMorLE4pF83RSg5/nNO6mfzdWofLVAb/x6LtfZwZiS8GJBRjm5ODL7cSgw+1W58
ZVrq3aId/i94JcZpnUOrvCPRmwSkXEWN2YMjx282cqnZ7Y2OxEBrvNiUdzON6dS6smCSIweB9eeI
UuUTSgt1qp/6NnoSGuInmCNN04VXs92GnSnZdpc6Fr+21OQQf7IAW8VrOhmP1KA64XSM6FZBjrAL
OoyEY5gn7TkF2a6LmroHfMKbszjYkcaN7YskC0EJVnRwzlTIYymBAJFk963D14C168Zn1nLT0vO6
f60SVMxqino3j2Es3vAklICyFp9PjEkKrLV32KnDgIaQy9WvuZh/DEiEVWZ7nbD5omev65R58iZS
8uHotPqy3qeryxwj2uc75tB13+5nk1VUlYpvg2usMHfFOVH6MLAVGq4KAQ6iQiUJb1LbKDcM3uXV
tQsIdU7VKT3hGEJWOO0jjer21MEzkHjdUC+jW1CaWZjpgwKQWOik95t2Fk71h2ut9BWvhscygeT0
IrigwUvLuXM4QiDRPyntUjzl9oYeGabjNTs/8MTxLxguJw8kR9W9j2TBKNfrV7i3N7htXnY/xUZe
ZS/8AkNfgPOur+cyiXABxOfpKB3aXIwCK68v9T+bSgF7yimEKj0YMQB0WnoNuMKqHFO9iJg/E0uS
L/c73EUvTqL3V5yiGxf7kwtsAdEARZ102hRebMaGElDUdV7HZ1/ykQHEE+9i9j46gw/OFwfDK3V6
4GDpUeBIGsG3R8R6qzDpyBW63RBIyUfcERCXIKko4rOQDsr5Ya9LdtLzdqIoV7CzbVdPoyzBuWbY
hP/nct5zNSHBQFC+hMyCdGfJK7GsPY3KPxZyUd6nhWWCwgUI6EfXAVVADQfvbubwlkk/Yq+zx7Lr
SSQaiKZcSBPvuIeoU4qXWt9/MxbciC/BHdUy/2W3xXTpafVt+dR1RCWOvwfF9NUdBzfshfDKAMsw
q3K1Qm+shbibCZgUwHo8unC9sDRd50Owi5nZ+6eQ3F4KUnsRAU49eiFSiqAXs17ilVY4bN5P4ZYD
U70dHoq0wHutG+yv8cq+M64KE00zXCN5Pw7bU2Q8KRy9ohPxFXb17/k3jPoLozOA53uUjrVEh5Dw
yErq443ztKv6ke1lX932dDM5YFS4WXE0zNsPgvcBnir6asd47PdoDkYejvyCZxJx1Xck3MOXK1H8
CGjkp68eYuTpyRLAH2aN8vwjWUVlMzyBIE+QTLYr68pwLSc7Pkhk1WHPsujEYGluInfDtGLD/kRp
MSh7CWSW7CM39s+XEhCNNcwYs7aUhq7IJ5Y307iufP7ipFtRimywmhyNq6qJHL3+g6XOt05cn1u6
pPgPa08UUZCYEP9akmF5KQo+c/gu+2p1VmD8jKVCPGHSChSTuqMDxunknYA3htnsfAEN2D45HLjm
AaOzjXxlKiPsI6HsRUdm+Zm3Yoz50y/XRNJMiPt9lVzFBKa6Vd+oHAmucLtyv9AROjLzmEfzaqcu
KR6qrhmgs5bZu6pHRLkzhLhmoF8PVixfb8je/Wx8AQbwNsPlR/YySVxuIgptu8srV0adwJ5hwiJu
RCofAUdbYs6MOorKtCxNKyYM5zCC0wavXSH//FF91oX3U9QAV5VADV9Hx9Xq25UhAHNlH7FqSHZm
GBb7WTyn1+RhMgQKpeJKiXcJuwcnJHV+PT0W4aLirsek+12Bm4i8Umbolhw5bPR3LoGwNDemQmKc
OXxFb+VvskWNaITMM5SyjYEEW5TfynO/QBn5fBeRgv2Y76mzqEqIl3+k2+r2HkeuLNewX+jJEhO8
DwOa7/zQFZaYNCdmBWOzHF5+gRVgwtnVW/vtUq2nHKOESz0S/tgfem1exStHT7taD8lKlbaHm398
WWbbZBetMvYm2QPY1mhg/A60aZxMWHIbu4ewfygCgZQAEYFCFJebp+/scS6xh5UbPxtjWyl2aS/k
0bqsAvnyj3JN2J2Xs1UaxvIYRojBcj/uVuerWftG4SVbHfBIDnvp9YoUlQ7+jEftNen9vJK2eZVG
A1l4XMg+DOeWHIcLugHjh2hn/YXgareRt+LaWh8LL86RnhomIKti7ncKlautB67m9cpuvile4AGs
lkCVjPfzJlnrHJhN3T4ZIjlfVWLrtocdmcd1vJIb8f4QlzJnwAzvHFiZuAAKKbRInYMpAycXMnpA
r+XuLoK35b7uI4JiCDlLsrXJ1HrIQklPrQc/oPjtfbUfGkyzZfvBWcxD08vH0RwmhJEjKbB8mAVz
kOaDAZ5WKBcAyQ16AADn9ZAXWkp0Dpo6K9EcO3j+z1n5v3RFWkwch5CmDy7Jh4ey4dN3fBjJtkuB
TwqU/o0dK2pKBgMgfdYj6KJxwmGWxjg+13Rz4rJmStA5uNe65n/yGQElouvHj+n9xHmwT21OEFxW
982XAPwyFi8pQ0Aol38+BzXCbWoSPTiQJLLLvfTdEdbMChF6fxnC26TiZMbnCr4M07XrotVbj2HC
+wEYyVO/x/p+k4ouDXJ1u7BL55EwiqlLCgWhY+R7EoXPIsmY1KCLnvRcbCpdxwMok/BJWpNIdN9m
TWgfI/HSbAO9R2wI0Lkshzp3HZjr5vTDE9MGEdjtYkd9682y1k0tm7xHUclxj/4olcpAGVk6ahpG
ZFqxg8tzqeAVgxpxgtN/N3KwYC8JEY+i1EAi6s5sBrVZ47WgeRVYk49q1Cf6XxPGiJaEzOJR9Z0M
6rvI8P3xExveyBydPyFd3P9UY/QlT0gDqxF3AUoBIMtQD2HbZZpSIngwTJ8w8L4R/yulBQzsbzLQ
6alCDN7qSspwvEO/j9kcbI6MyZI0Kt91UhyraaNT3tyPHlBfe7lecWlv9xgbgunTHvTFFNPHRIx2
QKPIEvYDPz+g72bD2SCO3yddveydjEw1NhwBmkFc7IIS4a787LOmeFH3iZHU+QPthewTLwcDDeDy
/sJ9QC2q/RliKCTOdU2U6j57r9dJn5Iwmk2pZUD6H6noDdfovK8EmN8M+b5+AyxNfS4pZ6NNJoSd
aIiJzkhbAYmbaTkoUjjavzFFF3miBsfWkNPsbYeEkQDhicrmi6mMQyMSutzTC3DCFw5YapJVftei
GUGOjcTdP6AzKVPA1N6EgS4Un1UwaSKBqgqX1XDyZmOs/vKHxOr/taoGyBzzZVmOmMLzHM/8F8R0
2RBJHZBQ1XamJQDVMcVsnMwlQBFHFBgunkYDtPPjBoeIcq3e1MtxT8f8EB/I23A8ZRLElz2RbMCM
NiW/NEttNBzIcR2UUv7i0cUE9gnd3XNpWevAg7Oc/KpnLWsJcfHA/rQvCaYi7yDVOPvzRqjTHbdG
N/1YeEnmci/C1Zi5LvZYM/PshImQbz4NHb4gdWaHgWaXIHdEMP++fTf8rg3vgS3m0wOpb3+i2tul
7SsrJIPxI73Vz+nEjVCmO404Fe9WbMa2/qk62eBPOmWxG7TpuUDlHT2VKTBNGMXUSARSWVhEXzCJ
5ymHHNARGD8CxDqhBU/aQZdJ2MC8m0l9LQeZ1kxGI7Dhc+alk/cWw2eiNDHmx8Y1qU6E+EbZZ3HU
EWBuXAUwgAyEqONx085YrsrJGWcPjRqmszNZxFJSjUwEfqd0cGNLRmsJc6ACHeRDyDgTEtbWhlpD
xdCuu4ncDMj2DlS85OrB26fgVf8SBwlwNxz4gT/wRuqWQJcbHl1CMbB4TC8VPcCDzD0d4kmpsoqY
lST23D4UCMz3Hpblm/R6nQ8DgQzgA6A5vhsHH7O6lhR8QaWoxf1CLCga/7GQ53jIxQkg4bUmp5mm
DSgNmW3D7HFeKtBOpBPF74K5GeqvE3xKUaBjHKw21QVsvrxusXlyRNt/w/qEYOt02gFQ/uxVsPsP
RpVd1VUVdyshkLnKNdyEtyNdnf7IlhxFh7SxT2wD2xJWxYzh1CsxClMiDdImfFrUx5UTpqx5kVm9
rRSF5x6K+xjSF+BERSyGro5pYw0OUdzwIVlRnR3saVcHK96gm1edecKtJzmkgrfYDqgvbxUGx0sh
yJrV4At5L+awJ+Bs/Nj4WnQEXaDfHdu47JOEygMeaD46yq27wbj84ZpusvmTNdAbC+V7CBplZw9F
NJGm7E1Ds9cxK1hUuHwg45ytd8Eb6uidLJCPkycn8SBrDJwIGhcGSpqAOBa7/RFm6zCgZI8KMPwv
rmwXlaFD3U95Uk92eh3AxnyPTGVuKrLRXWNa4MPXz61z0NJas5uX7kxBT+ZJJVblu7JmVsEKXGBq
h8YJUiCOEIBgTb/D9q/7JlB6+QJ9BQi0Th3hcMCOCrWcgvEbFrDhqHefe712Gl/+jaOU93N/t9Hh
SBh2Uf8Xd18pQmxAbTdJV5jRGQvmB0a3y3MWjZpEATCvry6lu2K3O+J+LhN/z67x9O1aLNrUVW01
NdJ68yoaHjJU0iG75hjVXfoSZbHfZpjZTIeAUKrBzV7D7I6WHgYgXe1GfCbKFgb0cxwzQyQen3Ht
B54yJ8yNR57kk19quv5ZBzucaVJS3TaBQwhCYLrFmEUAL6yHMYYbkf4eoyw2SbpL7OG2RpZWpZxr
kksl2GBb2miWFxDLl9LEifu3ipjT7SiuLzdqNu6Vir1QdzaUzEBH3n9DzPn+S1QzVC+mYvle8FAN
gXXovnOwIE2MjN/1iRXB/8WORZl7sKS/+q6WU/D4gjDN7SUg2VyMwKe9rzYwM9snabT6iw0Zd6Pv
XQZsxXPHLwDDo8bOO6RQE6NjKKORv2JZh3iQcAQak5oMUul0olJC6cEzVWUiPsMryDWVujERozMA
roSHwr2CTEOCgpdMu/dtZ6E8+8S8TBzjH2Yuem+9lgG2y2rT5Ygg68jZFnZwX5zH4hC5yqB66J1g
ZWUgjUy6NS6S6Pmz+7IvVSV23weQtlhuUshoy5QqQ7eckK4fg/BjvvttiRdF/pvAVVE09qi8HfGd
WxzI2Jcr12JepwIGxGr+7xkDIyfSjiv8P7hGvVq4QflGDC9nTEycnHKiCgRsVzyY2uGWl65CexQv
cQTctRWzu/gralbc2tRBIO/p8qtMuk96GHnttruu1q3CBfVZYfFauugb2N2CCtR6yPTu0fDHLY3m
QDYAPxEreuZO8l5jW7seXLyZlu8VfgO3ecPvXUI6tQdTcqtvRvvyyfIqc4tS9FRuHqq3FmqGobB7
O5Vxk7XCg8TGC45wIJiGHj7ciCfxiG1Kqy6XTzuH8OsWkeEKEAvoROT9HfDVCTauHfw3Y059/2kb
vEEUenZ6l2u8W0TsaUwh8EU3eMFzLcSnxc99fm4WrNWAiC+hd2WwKw/BpG77dsfbn6O4n12YwCB1
cuVXEiJmq0vOgtEPuemDrTjAcabzLHk6I0BR+xlTjkcD6Q2/cWK+w23duTLTPfdXQ8AantWoI8Kf
z7bNvZEXeUFesWKoT3F45zhaOJ2XZ6t4uG7GJtaGuziqXc78kYo//IDFFU9P91ryBf6+kfwzPLBM
tE1Hevdv4TwVQIPblQGiH93gggH2SRoAEBtDQJugtcj/DeaKDT9BOHGIs03hUphMwkcpy5Qgq3L+
SMMZJVZA1eQvQIG4b70svlXUoe6BDv+dYyaI07pCP4eQJTiSj85ZJ0rQVwHZg2q1NGlgD7yPNEe8
AZLqjzarPywbtvtz56rWqWjWVYwJ7Em4f4G+WA78WCE4BBIM+41fJd8SdLCKGeyYKfb1PwGtvqzD
th9UvisFPnnYOkcsg7OS2gGYSrl9rt/leX+Mq1N8OOrO7+7Eiq4+6mUomhTolcPY0A79SWAi1aBe
Aq41z9TPVmBlM4SQbI2jr8j0yxLbe4ZHAx7nhb6kEQmtbbhIALk40AXlpCO1TB4l8dFrv8Ab0/Fr
hmFQw8YlmtJhYi5Cjm+b5fvbgbV1PSwCz63J0RupmkG48RkY9lOhVhGrx9x3blcVf0C/zrSG8P7o
pv/YTdl2DE/BBXwKMZR9Lkr9Oxl+3pSzlIAGkr248br4XY+RKyJqaOt9fafpsWvvZnByysEjbtIj
o1HPxE1yoh28y+dZniLHf+yFNR5ILj0CLa9Tmw8dLHdtnMxxiFdGqBeJoLCoGpAsYtJNsM6cDD/A
EPhB3gqdUcCsa5sNVRN7sx9/+HZ0d2jt8jJFxLmMUu2RqhDumx/bhcVOpDPnfLTYwt478elFftNw
sDseXdRl6Y7gW8ILR6hvPuFN8qupJvrZT1iT7HgIpErbk72YGcRJpJCEhibMV24nuYtD/bfRGPMY
jA2Gppv2ev9HOvPZWuN9ifm0oGI7ItHD6ily0CATtf0lxI+2qzFAYQjQ9xG/ITEfOUfgf4ZW0Oq6
Ch7FFFcxXrEDP+6Akxug9m1/c/ozFikfyX5m82eIJQpi41Qm46998hO1UlUejl/eAsc85MdMrxFl
i6qYxLWRr6ThHE5T3zQLuCckTnJM12MweMXguhKndi1aTY52SSMbwJAlmpLhyyAdQTHj5tHIBjuw
i4iCvMDdvFFl/xXQsX55VpbzHbPXPonUyaPVsu31Qm8Z2p0ZIKTDm6omGf/1J4nS3BditRH1nOhX
9q3UtFQ8kSDftzAs08v7xj6SqAfCyy/hSxv05NMuVsBHfec4seccZrRnB7QlyQWdVpnU/FK94kXb
zJ5J9bsuoAzWRXkIZ0gZnJP3q3X86/Fohjl2Pm4SzNoxfyWIWi0FwyJYFSZJDbjawEPkxR0epuvC
cxCyeB1UwTlkbwV9mjph6KYFEbBM9jHqLdL2U9GBN7FUgH/U1d3hnvFT/k/VCBqm2s9ElLvEU/hp
Wwm52mGd5JoZBxCROAXjJzBIOJkamczw96diqPmZVrPsPqgA3ZEpG2GgYYPwHUbqYBnctfddiRmX
bHabyE1Xi0v/FR8X22qstNKmcWJVQTtgO2sbtzcjC+ku4fuanqLV/a/Xgl1rP6EPiHaa/tRZoLOz
O1na6WI3R3qj14Q7Yk0ovnB8We5osm9bisLC5HlLREQZd2LlY3WKjJpP8rah6Udx3pZGtl7rBhrz
lANOFibgi8ku+1VlLL2PjthouyuAfTjIgGhlS1JUet5vONKP8iH2+SLmbY9uHTWLto0HvuhKpLzY
A36GFNUbIPp6AK2G/b55ylPvJ55vjPyVUjzRKCkqKn2Bbd/DoHUVs/naEtjUohzPHEhUDkeEdxZH
GODp8rVoKI2mydJGfs1SChWG7Iv7DfpWu1oCFrFWTmBd5mUgN8159QdABxQZErZe8Dc+xbPHAQd3
vApn3dufZ6/ugA9w8qpgzJ/pJPLGFcCw0h91XpN4ypbA5zRIR4br1Onl3Mdxp1wQ9022/keLJddW
jymLPLBq1OGrP32vDyQjXKJbTDO9HIqvxD2Cr6yUUswMhFAmwnUi8d9riGSB7c64CLlANOq6ExpA
2H236tuHGnAWci3QtGKkVEoSWauGxUMmUqaURRO/gZfbbUZRJ/ZXvMJMy5Bo171avW3qj5GGfh0y
RXIPD7WZgLpJ+Mt9Vc+B33UFZF1claN4YwUZ+qrcNghVrZfV2enJig14YSXH9mGBdLm+qd+YSYhE
Cq06akLQR0z+6J/L57ti6dWMxCdm8Q/YdVE7MY1h+a55n3sv57NfedbHRdGPCMgNnmVfApSQFy+r
q21Vr9kBdVWyUw/t3fCXoXro6UCtIsuww0jSx3RWp5ZMe1H7WxPFiTuP0MoW4Naz11cguoApJlAn
iOawOJtV5y6Qn57x/hDqPjXO2+dCioRQwDNeoDMc+SuEuXhdHEWO32AtXFWSMGG0DaTIr1/cgtMF
OgO60wrtud3z4QudPKO8p8cghvPGN+I0mRcotPOWqQDHJzjdb/vs+KCfz0GJOKzIAg8+uXA5FSdt
HxgANivkKzNz8SNtUpQCLhmXA+nvhUW8hiVE2Ksx0ZIo9g5nLb7bVHcMo6nqRVbIhAX279i+OxUb
1peCS/+/kLgyglRqGh1gU3YnPB+NDJC1+ktzQCeDtWBf5fPmdUn2/uC6WoNCIA2CieJTKmtA4XDn
ejIqDK1BNrHpxFPfarwm7emiFiASABpr71gx+3xiPRD68EfbWXwfBVd+HXBej1AEEHFSJnHnKzsT
JR0437g29I+FYoD/NLHJOpUlpgfeCojYi9BaIT2fs8IZ/DD8L5Td0Ud1D/btBbIwpb4CSfpNTGAs
CmGLQI2wiaF4NlOx3E1iR3lPwtskhGPq2sjTgrB13wU8NDLjcqpfD52Y60LkU/k9749CDkdUVtqC
n+MKDLmrxuF7QKXp0SElsl6U6SXZfenESPsj7DA4us3SMNO0z2H2dMFiMYD0bDwtVPJgPyLmvHvk
gHTxELzBDav0kPVvAfzYbt8y9n3Kx9WXNGK35pfT70SrSaAN93lx56iLDl6O/XaViMY4gkmjRipT
beHhJ2YG2vPK+RolSDQUexB2aJdkUlt1tMnOr5YWCcqd0ehiov3rmfXohE/E0bIPD8aBxjs656Do
GVH3dFc9nY0jW+LOjDy05ZXcbmcq8KK6PdkQEcnkCcjeKSQSEaOZqHK+moUKRuKBpmUOd50+6U3n
JONgxAnSxgCQu1gUsURLhm4FjhTciTtbjepfAYFNNCNiiLVt+c/Th0i9MejnbUNNevnRXVn8myoh
WgP8Zy8vkwE+NapUHFdGkn/HXpjilt9FJ3OYKc2IMHyIQ+FydwaElGhDU3+hXQtpK1AipjI24Ggj
/955tHx38Jp09PDJ1T7b8VxTrRBvVa/HC4WpaYmoY+Sl5rawCRgG7vcUVTfLFZosbLu7FWHyW28n
SaTPayZrdYvIiJdeNvZl6EsHWm/Uq2hB9GSU/niXoqT/smMATA0bATzjxF16RQLDl5qtaojwz2sQ
o6p466DJSKISVbcg1MszUsRy1AGsqp/rCXELAzCYp/zkk5D7uQ0V8KSDlwvY/xu2QlGJNrNrkp0h
UwdjSZoD3jbYyiJ+itWZ0nDfKpG2m5FRIGU389j6n6M3pDxvW+gu5LTYFVEqip3CKVTsJ90I5g2v
s7kTIDKemWkN2pUZnN2T9m9CqTPp+s0kygdrYuZEWeNrRqZ9X3IREmrRcg3uhZxTlEr4Qut/pMGy
mftE4aPbHZqlI6wH8d9pkotfXSInXza2vtn6/2LAVqyM//UAaycVjF+dPe+Du/UyW5o95f76gUuv
ofTHCgwxeVYYt7IGMt5kw9Hdbadl+mJwxfB2aU7Y+ahpbk7oRBPQNNN7V4NLNpszr7pIL+q0H/fy
BXHFDq0qQsecPImrOphQM6+HR/x7Gt8VmOzwEksR3MsGW+pcAmpCb+EDunqMkINLHIbe60GU2Szb
zy0EbWODEMF7jSfkXgUTD9fx90vpw/ZoLwpB/52YepBuGr+xP8+M8vQXMRwrZkxjJO66cL6xUr10
dTbnjZ1EcyvnyxJvNMrr4dgjy8r6seUzQ1eILjwhliRNr96m4x8Qzfd7e0jCsiFbzdM5NHnp6tP/
WNg4JUAWiULAsN9Q6I5g4k+U47hzmzox/SUgEmQfW9GuOT9djI1Y/Qss44Nne3EHoVwDHx3tlxnN
qQgNfF4nH1j5Vd1oJNfBpf448GmrA7rUR1qzUbYvBXjqBSMEye6c3O4nGxpPEGydoSpexReV6Tdl
BWpQeDsRMPq9+c74fY1/5QjKLk3xRP0VAY4Q0mmvEFoE9osaynYqhmKzx0HpykKwvspPqvk99szg
Fx5joukZJV9m8myPC+B7jlLqB7uIvV5Wp8S0FZIqJ2RvZhX4skz73hRDBNxhHsG3X3H+qcyvEtvU
/PWBpHHgTzLT/1uirKeQvtM3bO3Cadd8qKBrZxHjKez3FYvKIkcqxDRK2sxB+F40NSnDl+nPt1Cs
c+y0BIcpvYWf9mjaIoTD26PCAmU87fk+5CijR3nAPv5NLf3eYZF65cFM2R3WEUFUL9I+vWWKqNtc
xuuj7fkM8lPY8/YwExCgHc45i/x863dCzsyb4DCDRO7iL53q7EDQ/5iG8SkCrAPRVthAqJXSku1W
4zufxOzVTDC1xYWxWRp6nIV7IUXysIVz82gHFdL+W3Od2aFIL4GAATaa2Jwgfhb1d4g2/uINI+d4
Nd2qjn/j1ZXUbwQTTad3GOOTT2GbGavDR7pJUdIm1VowecKbL0Mru/QoVB0y5ytxdKHjiTKjAt9M
c0XSBtW3pvC+VTUPjCh+5p/iXm+F3xJFVMdPCPmQBo/A6rZFRjPg1IY5+tbZVzCkaPDSbe+cJgJZ
FU6+onymTQYxEAMeMLaYIX7xHstcyEaP7t+0BkOzH7xKOwo1fqkgk4cImBIq3CaROUFxb+wQuvVv
GvG9ISqSZRAtBvCfevHE6cVf6SqJRtaYnLtcwW4nRagU16zqRT1XNGnX7utT8grVNMdVaUiYPMsE
P2NgOFynDD9lqdxYpuZlWEM1Maltcr9LG+vaF/DYtkki3/4fIMuEmwKDq6OvFEnDehh4W2zWTs+a
OMw0TuHZ92lxR7kHOxnylpP2So50DltlGT3h3yXO5SnuNSJK1WgIHrnjdWMi9VjTCywyBsulbWXx
L141M1YqwEInK5vNU2a06tkjmWCmtyDuek5OJihh17U+t2Vzq5lMhGOyEtl7ZVCwwo59w1sIvoM9
V20ah1rXlCDEH+SCkoPYxtu976937bSASKgER8H+dJcujGNZs0JEq8Aza1LZZuOt6FGS49tU9fdn
YpICquMMTTpZljF5Go9ezIUOo7ccJTWjkRdQ02A4sEjxTeGmy3Ko6/CbVwaRxJpIsTSrh2aB6Swz
xXW7oJZ5uQuxVnXmdfROBnNzcaYvRSaD20I79sBBuV6CYAMYbWqaZNAT6tIOjdkgmR3vhg1UR/eB
9kMWcwSB/naGoHfC6s0yGHkN6PSxTJfzOfftoi44Xymkx/lPUy9KLGMQkrahrsr13rFl0ouzW/Il
h9d6FbH0DqJBBk8xiO98BlAt9wJv/QZb3nR05ZmRKGbrg2AebXcF8bKL8HAiL+M3OB6Fuo/6AZK7
PeUsicjm8PbIyMGR/ZSON8uPDmmEhNHVaGOAngHM7SMhtj7pIMlbcrSvXgXo44AZ6el2kdw3F0jO
q9l+d4Qyi1wufM9lLWdbQiUt6y0bFdjg0IdC98qXDQYtjVRU3IAOGeIsM4wzej9loxRC/ZfCJqMa
uawhfni8zLSgTH0Kjyfi8EzbKSzhTb8xIX74XeZwuD2GjKArA0g/ewf3vtp7JH5sczFy/lhrBjrE
iDb5ff9JKBGVf7B4iPEaMgdJEnCG5X/fClrdPjx6mAD8rwk1aJsO7wuzMF3lHNHSX7775ZsxdYfa
7PlgYzeHsz0g9k6tRRmt4+ZqS407vlKX2OafHC87b2t/kmmY2xL5ExMJdYPUnaXo97m5J0H058bQ
6xGs/fRL8RCqClezeeOczlvH904Yjhtvx91vm+4dl1cKVEf8iobCTbaUJgZqsfUoMTdTDj/IYxVn
6YVpBfxwkVw+Ppdm7Q7JXlZCLASHuxJVws1gEzYg/SoPgPHJqfihVwpLAMMgmKspgxGTo/Pi2E1y
ocWXH7lXupm2cfySXxBvEGkjhUyM1fOqxG44LnB5IuPAzDFx2lJNKZGYz3KvcKuEv6RHNNWhHp39
nAi75bmqbCsR8og0Y1T0OU+ODUV3XbhOmYWHz9U42A+RKm+yOzGh1izH5ZV0Dl1unAR5cqQnsuNN
6IL+/Mv2SsF0Viqy52nhW9JLKp835pqmH7sb+OtiqrnyJFaZyjR5e9hCm+eHOcfkmxjPiWv2kvZS
RImAyMSabwC7kbmDS1MUK6m57mrdeB/SPelzipa0NP0CEopHDwFntvCYTALx1ryTF4wClwZKvo53
aSOBHaAnwKCJrXtNlIbXuizn+SNwVM2N1CCwdSft4ciNZeAs/P2+y4Ol8maonlytuj9XcNdrtDHU
qvkZgxx6XxDdrMKfTnvk9IvsCfxUGxWWI/4FuQCZD4LMXVbXavEP2ZezSeg3k9vpJtSOQgWugORp
kY7R/SkbNQRd3LdbyMOd1R3dG3Ck7hUZa02HAf/tZr8PJ8s0UOgUv3ij+XcKuekHs6gwKmGvHuyP
aiqWjkGuSq0I82eWWWPpTluR/BAnQR6hzHYx+Dbq69uOnvexxAXMHF7DK3ZUT9ut/dZr2PTBli5x
HWiCwxTwMb+UT2dUTjzC2Jw5RC9KIP70vJiWy5mmj1picznw2sUpFAMa/pOVTUGJAjA2GJahW9bk
KWqC2MDcVR3v0r5OHHGO5w+pCrkPJ/sxBNdUQtzM9PCzikf5Db9/m2bTIcik/LUNN1xJRF7S7DX1
j0ADyn7ktWmFTtSVYVLbB36xdvZceNQwnRW9UqTp99cnRQibR7/GUgcFFtk7PumWiA0vF6Mi1/DU
X2/pZEK/JPpgjO7Gxlcbzgf2LEFaj/XsvxMZr5QEX0c7EKmFtTRDHvLsYbbTXA/jWo/BfRAmVJJP
0zM4lpWe9NSiE4zlaIStGFyqDC9GaCk3lr4rDci7nDhUR26MDG2n2SEN5hf7s6AyMcK04l7AJJJC
n0pXpq348bVivRLITy+EoVwXp2fY/ayimRGGTWZ6gVtLcggOretkFKOO03bqvZL+k9INYiRJQC5k
smJzjqUxasEnLihWa4Yw5glRAYskzr6X+D2hsRqPuDx04iPPke/OiS0gg2RHfart5lotXKp+Dq68
jnB1ydep+Uq64hKfrdAr9gblNrUq2rBCFO5NONjEHb74VwaGoukFgdrk68LJUpgwUDgpFKKgfcsM
ULMbTrkufoINPEJc4lyNZykNxiG54S3NIF2pRggTXsIBVHsPUyxXLMRNKgDiEVWnhk2VqX+vso0N
ubYG+eNGco7IcIYTBkuzA5aihSIzw6qsabgVgVeyEZILqcHAHrglGIArSxEAIb6vfAlLsoty+dqt
Xu1Q3NVDx9Gjf9KvVRWwiI0HWNj5NvaDlZsOPL+2Ji0MwXR79kKWL10KWBQWBlcQWkyOb07s9ee5
6UZfKjbrZodpeS0/W34lwhaXKNldxvLEjxCCfMr23WRO14ZDYggmRIRX3TvgPFijQ+aOYb8OZgHN
kfcI+6+wuT2W1S0n97w+y7+N5Sz/AQpRCjOQFXvSIGoxz0Hz3S8nsM6HllElcVRIElOGOEs0LzHG
9kn422FIaCyvuJhQLkY8v9cP39u7AKBIspzQrxr8478CupziTgU3pqEOZxDP1BXl6T2Wm26sL7ie
AIFdQa2AMSxtEMLR9pqXdupKdYlvqUUAedk66l3z12YPuUmzuxhdNF67fJsEt+zI8QXI9/rqj76N
pfkHZCUG5N+OtqejpR6ZbPH/f2KnFrBsyeXZHwEN7CBlCAFb0aN6VX0NeEVzD3zKKY8n1xhj7GtN
w21RNkLP0JUoT+92H0ko88w1ZP5q7cq0EumYbsWs/FRM2ayqNhjv+Zoo7mUQpTBxuxcj3RBsQZER
4mmsiM5eO04I9UNBIJJb/NoyllUc0ePMjOutlIqnQOP+tH2soGGdba/LCUBLm1LxPXpNo27CFrvb
TC+lqmspfPSqQQXN4FvEnaaNW3p3BIVgNArf7kfdJppDNgJNd9p4MDQ3+9DU9rUGBapQu2G6Q10M
rTu8ki1icOJUwktq666hZFJiwKAwOvwicc9uDGwsnzUy4OJq7BRws1NJhaz8+pot4Arbqbx6yvH8
VMTM91gC8ly9L9IVAvcrpHwaOZR+lKjb2ulBH42c8MFm2XBiTJO5NDegR0wjkQqne9jjoIBxOcRf
hlqAAb9NEd0j7g3vNzRCmJMIc4NTBmQiLPGGRucjkelFNt+G31RKjiLgoLtm3H3XsLLSzLw7/41G
D0qy9V2p+uwyqEFJxkb8Qyk9Tiuxm4UUOfC/H/Wxx5n20Z1LZP09AYNSe0rmcwq3kK+MHbAwKNQN
21UDY4WSqiWxqGbm4syU7xmbhfm2nUss2Eielt6/p0jS4mQVVABR05UAlcBQDKUEor1+raKhc9UX
V0IASB/7Nkg45wLAYZX4RH0C/JjMs8d+V46lBKZn0pSrlI8c9ZS7VKIorMmceA7CAKKi8XE91oFA
LgCO8IbFrc0HuZgUj3HxUT2TfUrPHFRaycad788bb2Bqyhc/NXhuvqTsLf8LJMT91q35r9V4O+fT
Ergh/upp2kyLVxHi0fNZTmgx6IZDc9cld4keVWLeVvTdOkjnsAq4bHe0qTwru7JixVuNFwrvZNvI
z2ThezLet/KkKlbw7xGCVsdC/iXjkVK4Tj5RT27O8D/av4KpSUDtigVo7FWSLeuKUhypU/wVgHGg
5Gb4RlKzSPWi8j374bQSPwRGbmCV8hzWaHX6ceNjLtC82YYwZTEG9+ZQuBjXarhohqZQTTqh0t3U
mVWUKDelvQeuLwdJd0jRudo3GViMnSMZWSLKYw1s9CTU0Lic6ZtJRImgjyM5VGo7XzT+5kYtM1p5
fpsQk7Jf0NQWJovqdjteI0JT9oNKaxYqIolNHgQNEYixx+jxkZz17tTBVDnInkI65j5i4tqjAUf3
DryIUcDuTOF/Wwbx0NdIhFQdo6c/AcRFDBsMUMI8BoXcgjV6zhWf+JjAEkDi0LkViNLFVZb3T/br
F0Zlm6XiI76mZcZsuCFBG716cdq0SCjyX2PYkbWuyuWDsGHh7B+DN9nBxRyWMY7SnPYh0yUqy+GF
6y9YXnUeSsr+g5KJaduVXfZxCJJxG6avGm8/+EMn8LuOrDWNfDd8Xu1kO+F9n8Fap+yl4/E40ibR
nnRYCHkqElvJLkTP3Sj3ryJMNi29pyb2iQWbwE8T6kTBb8kdH0+xO4bkhuc6HgsZF4959xkTgpM8
qS+pO0I08DCq9W1bXbr/WFnQlKCP8FPlhaq8V1BDD7RDvdf/Vz/Q9J0fu5AYES/ps6i+ejjxsMHW
hZYygE7ST0loq2a1Z3awfJrNrVvlloNjA1IlSGyLZCfu6JmIGUBpCY9dKOTgwnhfu4KINBp0GYpM
PKxgpkjIV0phwDf+ICGGA/F7rLxDOOsavHitQCTJS0o7VG9zhnwrdeoWWq9T0v/W3tBl4IvY8G4v
e1XVejipy4rxYl58V2tyiYTDwqxPMDroxtKGH4JeL3qhjElQf0zGxE572XUD+TYFbW6Pf18YPQlX
EUkdYKtFrTB+v76CR1BKGlN5ndSmr4qGpbzse4g084Inf8XlbV4p74S1SHDYLxTlh60K1+dDLAsw
EqWRKxqdYRlzxKCjeGjAYscqQ+5Oe2528PvFj7ZQbPLhrjHe7Nm1yogDBMDucD4oI/FRl4n9HAm8
vLPMsLl7Dzk5U1pjelHbb32rugXwVAmX6dGC6JLHyY5L4EHjDoB4v5+rlGJhrpgBBTlwQNeTJ2vH
Ql2LVIJBUarWVbMz6YwwmbOp1KpnpbJmpuWQJpwKqt7rEkFdgkhiQr3wpAEDxze6ds3IRK1elwlg
3ZbA3Of7OX+TxDmjpDM53XeZAUFzAbueQ548A7IRzOczQJAuvY1IeWxYHxzawGed7rujw7RVypH+
A+eTztjj5ZR7bTUV+VHoz9S156P/5hJUjH2MlTKT2WMPHgFVEsLXAlnP8yyYEfWEyA7ZBVRFoA7B
UMzNw+dmH0FYeZxuDA+GET+YOwa3agkmqflfi4Zd+qhwBAuXkczea3wXuf+BKuCQQcCD/YmAmc4M
xXQGmVzEn/17k7kQqcXwptI3nSA9/Ibhe4bsO1ln1iSyeV2jghujGwmMgG5oQ/NvglY42nVxrL7/
yWXWwNsiGrJKFaYi0B2KCo6WJXlvjYTsCixecNIHsy+MBgu4AzUVWWrDwofS7GUpEaSb8cHJvkcN
60T+udBsAQLQkAtEkU+Qj7JnBPUt3zNtnt25fqV+6QXG94MZgAelezpzHMn0V0L4L5WaqeU2t7hR
AYfzeh93HCK6k0MVtmqtkYW/DYX+brhWLHh3pOCD94ASYy6G/eOYpJHtINVM11Rg++Hwb+GlR6Jv
uOjI3YXXdfeH+DVWkeANVq2pxjjoHZX0JyAlzDh3k/hb7ku2EAST58qqvHMXEB97WU8OFCTtMiAM
n43KcybeFnelIwS5PqOWlTAL268rbzrTJNU6FqBOvm43orHaX9Z4B/BrfZkmZdFZWwBwLXo79Brd
5m3U3986U28hu39tzVUcE28DV/kXTZDqB8fEpfGSRX7q5eyXhV5Fo/VUS23aAY+tysLjhc6El538
FNLEHuGqMC5bKcQ6WeTH+kXlGf9NIwnerQwTwjrvjI7yiCnzW5A4Vq91KsP7t9nEIQTHp8MdiIld
PqevhisLwisojrJg0LyqqK07jGxBFQuWrtuOh2uvKi1Owy/0DGKrjC5YnA/xlLgy+VXrg/67FNVs
W2MqOLAq0CsEVJsqlz5Z/TbXu7CHoz/sTZ0Mcbf9nReqXR6kBRfOW/ZKT80z/73y3NULDvyzuIZJ
K8vx6DXQJ5mDRo9WnViZT+qPffAS+DHYTrxJJ/0zWFgPxloHhg2BFiGuC2oxP8jHyAWFbvxqFiou
Bmk1votOX1gxhLlNfMGceaGTx/oIUOkGoQnJQ4orQ4wbk+Udgv3jxI0rYIivZpvCbjDlzw1VrDkk
Oq+M6Sc9pD85Ifu2mtrIbyY92rhdhVc6hhBVaOoCRA39tsr1UM/HZosY4JT5tjnkvWQ2FHTDibxj
RnBCHkYotPk3k1I4c2vCatHd5MtEPDziZ/MTBDzhtNVLvMh7kC5BK8+LleZpJu4YXCWwe/bqT0RD
NPcpeAEseKWX1SLxlo248mI29rcpUIepRBvbXC4i2Ty/uln1r+DRzu4Z/adKbN5M7cCANQHTtvpM
3lm0WjCYHpBqR9Ar7H8Q2SqX3kQLf2DzR8yTO93ZFl5CX3J5X3INCFX2aWR+97EcqRWNJVsbJErv
2lPK4OjDM0Bmmb9CA1aIZ7mi1l0989W7LOrFSIG66/WjJFvQJj+nsG0cs77lILb9U400YM1Smw6b
05xk111Hvjdl1OCAPdRz446qIa7Uu+th4++gDK9tkwDBvQJcdbiE1uertEqVLDuexLK3BpSL8Edb
2ObyY/8f3QmglUeSIjhYlGba/h6KLcuxNc2ahQZhxpJQVOU8XGvODFbBL/0qJikckDRV6M31sl1G
PiUOPb9lY79vxSZ5HiSs38TnGkm/5r9lzSX7fhj3XpgG9rgFx8Bj+Mw1Ge7cTGsRl/JH57TQ2vDg
YUg44ovSlGk5V1y61jKibUnn4OTdL+RgWSpb8yazAivegpG6isPwLRvnNiuewlzm0jTVTa8cc79C
b95TBGyJM6cSbvyHQXgltYt0rJfyQhCjXn3fitoYHyP00MNLhoSBYDlcZGy6/1rtqB/eWJDjmkeK
mE3KnSF8ROVXvGSHcgtFzvYY/VCht53Pzzw9mjGO+7zxlf2NuaFI9gChtgtEmMZHFhio0YRJlwLr
AgvHGniyGqtFTl7OSYpXiYDsayWa0vnLooonaSxLGFbFYgQZmKk8WSdm5lPFwA5B31TueOl6GP4c
HHm20iLQQx0JY1p3khLMgjQSQs8F/lvtA2cCjRILirmgFNYlZ9Z7DpDrnNCSqDndO+T5J+o6a1KP
X1UM7LXqnjbDbSUrjhJUfJCc+RE75AmB/A/9pIEySH/VJDKafscHAZIWk/u8P8hJE10aqtuKGlA4
xzlby/UFTD38nK89NZ5Mc49ydxFrNKCJO6jHggel2sG9PQUkWY8xdKtCBpxIf4KVu2U9zBmcexCV
ZNzzT4tc4TprBWCTWurA+CADqLi0f4v1nbvN+474hnNs+DgTVLjV4sKSAFf7rDIZrKpJeXurcZkR
ivuq/BPlGbg/a5QvT+Dd0nQ8GYrA2WiOX6QrmvK53brkzhteHMDB0oRBrsCXNYcwBU+d0k6tE3/Y
BF2yBYExGHL32rWOdh0NaSQtaca96jdc08zL2ZL42RQq8jY+s69gC8R55S3MdjWd/pFdyLeWs6Lk
LoDQCkMzcRMHcseWRAVqcE+MBTdBR2OAKc1Z64V30SdiMIOv2bkvjezkx2VtAj6zVnHOqQ3heNLc
r21Y6N1mz4WAgd83ok/xwvcJ/G01a2RSMKrjYXKc5XGhrW3wIoS9pYn0BbWg3+6kiXw1E9f1+rjs
fXnAuHQpXesI4ztg+IPXYDThZSwRY0CR9hvRz6R8H5jYgDPm6/8VQESKEZr4NfO2lmV/UGJO7F5o
ed6kjDQw/EyphlqF4D6C0eiA6EwTGWpbm2eHZqytcUufGSpPzNBJGFG5Ugm5t7yqmhg7zk76RtEi
YQ0qWk04+PWPwVv9gguh/HdR/UiPhgU9fMwHvHkmd2ntcudnB6+topfNZeLTWkoWDNW2nV1TdIFz
a4flQfzcquQEs9H+vBIhRqgTS3QijuE4orVL6ddtZUGoq8mt/gKv3AJ1wO3ARqd/FhCZEpqqaTCU
9Mx3HRFycoO//7xx31W+kJI3zjx9pk32NU3Z8dkYFTH6F77Rb2eF5CoQWRq97zau7laOhqT/eP61
Ariz0o7jFRiTIcrGu+aA3nQ16eEGzMA24TFMwPxyL0BOgYcO+I8VAaeLoMeE5+SesJEW/vhFTeyi
yv4MfOkLi8O9futqdfnhmw2L9f4MtrAAEK9cI+CfixF2RbVwF5upIqwysR3c3DF549i8jFLtdPLN
dvNeUfBPNGAz9qzyYq9N4keGcO5XDDbhQjXPqiG7Bx+OlSDQ8IzKCqKoPFOAwBj3wHai4UhZIwq+
R0l1ABgXpfHZbTqj8ln6BLUtv6lcPpaLLiBCeF1LY5IeZdwZ1kE+1FUBeep2662uSfZtpCIVPqCV
DvFpjb7HJBaU1479wl/JEwqHWyybgWLF5jl6HvcGNaE+Cd5sORTFRj/jXQz5tMQyRAs5kjQ6tKp2
a0+sX/iHJxd4kRsmE51AD5utfnc6Q4CA0IeaG2j3xHT9r3gXJ/4Y98dXg/UPnHu/17OiU2KJ/t01
t/Cg/CWWeb1uj1NuvhEj8WlhH1+BdkmgcO8+ZOfkWWWg+8vpABX6QybiJ2BGkGb4Omz4Ep3wVKLu
jjvVsxxl4ojfu7G7m/qEZJs9szJI6NaiNRMqtRO72c69/QQNhtvnML5CY920IGVEzMzhAX7luzkn
6YfI2InGsg3/lR5R7hFY85EuNBCkvSyXhBYCavqcKcomv+/RSC37O7KdzvB4PJTuBZ2tr5b2ARKD
1VHQxN5goIImsFZwyg6Yuih1T43CI99gNwXEou1ZU4UuSX+ZIcrcXRrda/aDpjtNXEFxTYxTZBCa
aChcp/7eJtQH5x7JohoCsDS3mh0wWtckMW8ClmnE1rqZWn/MgSe3nJRxAj/Vt3Q44QzKJh4d9FSd
qCumeftBlTUJ6DLYrq/pmrHzmoLH5cJz9wbTH0CdmTEbQ8iHfJPMXv9LPxzhKbQyJaI2hD1q00Iy
YVTsDrCRN6b2S1uRkGZUFsIr61uKlGlpxPGTpX4lac6jevNzqLKL0hg0azwA9+NfXdRADVhwGEKM
js1mHgmtiu+rt+y32WaSTmAqGLLQdjNCSUBlZwfnEvYuQInzUED84976/qEthfep63wZDW+ZmAzk
LO62724/h6UOTUIiBrkD824IhV5xzXs1lWDa2R0VMT40rOQeZDY2tqX7Q9mdIAQvAaOKzIu2BUKL
f6csGEleqUC7zOaMVgvELuWLbmgWFAbQnghBf2yfp9KfOO3BIXsM6EydbKXfhluGYdZVOfOImbdF
cNJ4HAKeaTKfzJWkLA3NVMFiJpunrREC72CYLIUOXTmf8tOc7wrHzfL8MI89ISoyQUKfJAfUSVL4
ZRdCSbn1TN/dJsfNof4C0sbBIjVNy0HxZhC7bIMo/fL3lCFsXihBwtRtQxjZg9eLDi6nbcPkKMNr
wXDxKjzXN6R7P9ZjLtm8PYpmjmVFLqEkch/V7W4sfJVhVYqX1rECd8s+sPOxTofPdN+e5ImZan0e
bgIK+aSkL3uLW8qZdSsA4jIlFy5MEQs82Jx4+adnYHkdGymVVdX588ufofKlOndYa5yo+u86htZQ
CV4DFUGDBex+R0yBsweS5W74V4nQkRTlPkihupXQNFeThgVg6LjpzMfII2/DH+ovPA++v/lMCqw/
39mnRySfGxcghbRnj42LFT+r8ToNYUW8GnnBNQmHTq6aTEnjLUq2Q4UO+pUIVFNmaBeXjiIU6nIY
BGLZDHL0mmubaQsvGMH/ADuybk49NCif6b+2ubuLJ2HwZ4ECpJp+6mLLg0rKE6tusJpVGDpRzG8L
ZnyrEyQcNiDHRxPA/GUeuorExWb7WR4YaaMb+qN4EAtA590EEei1VZz96noWndLvP02wCFJ0NeCt
Bb7ER0kwyI9tReD94aTIWGy0vJikKFD5TT23C1UHM/qpMcXLLDptWV/yiR/eKR+UOf9ibkEfCc41
jlWk2MOLnCAOSkAk+f0FXkwINa6LA09PUJ9xmNrYPEMPd0H9qBqyJo5v/T6cl8Gqgvm8uz7s1y0R
M21lvvdefQh//6p8e9Cb/p8papT/Zr+oeHx5rTqNo1xGTJvZqYoLUSh8Ws7YRuY88qHB7MwFUydU
PBGdwLM/COMerNtIKSG8ngukhvx3RVJY3b4TaKCaWxmgM0jRFoviygkhPvqpjkqvTZBycP5ufbel
ZgfG5fpFMwUBYrJMaBLc9tzBTboR3UW0dk+OmfmQPj1MMqRmtaSH3PHiQAcruxsV9ozH1oTTvRuD
zYjXgJlKvBy7AWMmGvqaFXo8BMynVZ2w9s093QiqK6ku/LTXDzwhENjXMD5muPE5TDmyw9fw7CGT
KL83rTsmjVLSbEv7f9quKM6ubi9CD5uhr2ihK2HaIqiUZ5F6b1YsxJFq3ALm/XBicRh7iHB0rMbG
6sT1tp0ktkLPceJGUG1SLzZtOC7Li7KpSV3//xJP5R38z5k3reL9HFhWpplEWqCYS1KCImmA8SFZ
sytU2btuz10NRG+BO6dkUWeOebSd0vV+375I5/2j4wWbpUYX4jKxZSkOXPdyBfwNVqE4w9Dzgc76
Vjddi/U9TsTDyhSIuDYH9/f09HCP6pMthhLKeNAiGNBaSKPNJ9h8GhzmNEopHHrBUmBa2jyCBVzh
B10keGFtiaNSFrDsybe503Zf+WF8eWV0i9U0iB9RQ1IIno/BiIvymGkcxQ+Fv+bmTEi577hO+amA
2TCHM6R95wIZHguHpsmTEy2Q3k7RFoGrmi6G3QxXgdduMjty+FevOy02dSDDWSCtVILM5jJCCo+c
DavskG6VwEvrqHfiK4jzyiYPl/VV9Z/7MDGc6nT3HGUWPx3T2mtXioS3tHRoJIoVvSn9UGiqJ52X
JZCPpU4+VSBiL16yNYa/VHJ/LNAbqiroEWi4qdrsIxl9+o7GHOg1thzz8i8z9PwnSyDe1Gr2sm/8
Kyd80LWIGqYyIx93rgkofT6FnkU7ZEk4O1uagKdwn+ttn3eOMYR+zds3gwFouZKh3mGFoLrF6y4y
KCkUgBVlXxYWrBejmJdU7n813iCEU56jj72vxLxokio3aOWvW0baqQ07tTXsJvWDBcbLeCdr6usl
H+GCWNEhAUOuYCItODCSqad3huv33AF9+Ls+Fkyjs6nY9Asb00LQtqG7HPd6WcTBNk0Gm94ufrqN
hPVFIi/B0RtZdbJIwazNDPx1yLyAeJ1zV34Z4ASFja/WhL8qnzZ3LHwHhhnwO+c+vgldaYQXAfZF
rjRJXu4/BPsdFiCifhYjAtnm1zeo7qgJQvu03etTbeDyWInh9JmqAZGH7m/1Flby4C/F38ApYZXl
a+wCZyu7nFGGVkWVexxaHXQHT0phw9pVnmDuNwnUBW3QyzYflndE9+NTolJaXvXj99p1bYG+SNTY
UC6tFtyO5Xyldahf+BD3ejxXyuA1j/6b8vU+LAMkoYLJmo540LT+XXnn/Rs+B1jP6rqKMhwWNRzi
IO2AXLx0LxrsN94QgwsxoqhNRmSVj+7ONrA1zQUILk3+/pmBwvDfYSQz8BD7ETouHhFfVe1NJq0H
l/YaeTXihtyvFY9JyzhKv2QZZxOAV45sUfidVEaHUNdUesIoX8IagvUh8RUeFEGqS8DudMOEJIu/
ip41oLAa0DHEmkrrEGPBHJo/WK5BGW3LFq4n0jlWCf+OAKsAxxxTnJ0U6KKtvrpr3U44QTE91WOh
YG+aTqQCfji0KMowLDLCNr9/imbP0yKlhXOV+mUgoY6DRbr0kHu7pmC7iTTTXuRe65bL5ejWjDbA
CrhcwQ4n8FHwEZbzOGCygjTgPMzv2BWh1FDVGOaMpMfHR17g/Bgv+ukF6NEENGk7eXqay7wOFFmb
AcNs1uqtm0unjGwG/gZ9oskYV/di4GFIQe5uA3eFS+5X1ujlvNwTmvwPV4rB6/bZIrxvjysMBuSz
fqh6B/hHgujuYV4KpG3hTOdGmoQHZu9AG3QueelxyxldQvs1queZNaIm5vH/lT0g4+W1U0h+R5nP
XyLcCrZHbgT3tNxasp6PRxgfkaY82ewMzEx1Uw5kOk32Fo2wQXpsFhoiPjqpNpapIGy/od/sfuG6
ppqkyGUu7pBPD2+1lvc3QpGFx+zLYypOV4VNZ+HJULp9CNlhFZHN6Wnfhe4BDNrWkGtRskfD7tJc
SXQR2eCvgb3dXuzif0pKwDDLw3Pf5+3DZFq7kg/egNXs1Q/qQnLxsoZTNQE6CSEmmDZdkFPXlRPc
CwqkCJju/T7vDiRl4E+irF4cD8hZpKDQmTVvo3G/JDTPV8zFDyFaZ7g04VdIEzXVg5KgNeYHtfhX
RfZWUrnErbdPZ/TBsGdfs8QpjlqspuaqG3uCPM8AohI8X+kNDJt2aBGMHSrghBTtkTH/BnhVkJtu
A/EyS8ENeCYW3Qd4TqYwhhFl1YrNTq263047R6pq2xep3X6MkOUOLy+n3Gl9hK7P+MDmAGBzezyU
QN8hxGpO60EyqvDQ+ZLMN/ahmMxd1mhQRohsJlUl/bZVMUwEQOgIJg3tilDRs5VdIooujVj4iMdQ
H1fcpezo69dvf/aSPKtVzDZHRXoDQwgtyej0u4xcRyFQ4EsgpF4VVxkO6wP8NLba3HGDpXVCyrxX
Xn+SYC1IF4xUGDFJo4FnILD+bpgTSh0QKPx3if1RxqgysL7cBBrNdgWf58CfGg4zinjUfLQMJJxE
s9RPj9uwGmJ0vBWo3aNqBAywLOUzsM1bYywWNa9eRxiIz19cRr5wzpLMwwf5p8L+t95z+38Cd0cI
8Zv7Edsi6BU6eJXCBrpkxW8QQAFcdjY2ebinqiF4EtxCMC/xyxHitju6+gI0pRiHb3qL49Wt8cg4
P/sbUzvoY1/Y0cBLptJMQdyZuCtfCM8rd3olzYFJW4rDSKu4x1vl7FZG+rf38hX4szdwiOly4+KZ
t3/qum/yKlQK2Uu2cqjmyhEXvyACQW1bLi8YE+nZ6RhGxplH6EKHKeGXUYMKrX6+UEzmi/FQiudt
M0IUVDx7SIpm1waj/LKB6EDaQbkFPZCK790ntgTlticspCL91NEzgjVn6kFqATn9MPnrNuAazmAH
setMSzFvRVMYVq2dwVd4ATvANkZxoDZULXdJuamgjBoo5PruC4tN8KOV8jhrzKHspHWC+xsW7/Qv
aKKz4Xbt84xfO7yyFGl905umhZQoSx6LlK1DSOX9feIu3pDXLDmFWgnVbpJhiX57Nv8UxhFoH7Po
bjnS6fE/VCkkjT7/7p0Rp4k37N5IeGEB9QGSkcGuODadSnRHeohIql5kmDQfGT9m09Zwm/m3A5Hk
k1drqcyQehW07V4V6lwmbHrcP/9mYB1+VEQ0Iqyeg96IB1QwXsYEMUyMUJl1xuLTyPyCSLG2xpbH
Rdx7oyh4LZ/y+UrFeUrGTMyu4xX+7q5nCIrUMvVacAle+Zj/r/4MPDmJL2zO3uflKYmEH8gmHMC+
6TThHafOmsuM4j94yVZY0A5KZbSTno+gABbpKcHXRZeOwjHftKakuWPlzS6IP9pgwuY6u1eMOOXB
tok9H5skBMVvgI9RLrXi6g9FAdjgd1b65QEelt00GO1uo0gjsUMYUeHgVGKh6ccM2RN3S3sMcSfq
+xfszyc9ByQfNV/nHshMu9rE6mzOT/lJJwCeN7YKiEXSAZ4XN/H4lpop+1G83CYIfDBCYTe7TX8N
6hOmk/uSRHPhvhTqm4gMpFtA0ATIduLRYefAqVwG5sQoXuJfiSSQsgI4LX4mh1OYD6rYkbJcq1ml
+WkVGXZAecn5TlcMCWfc1wKeDNH7Mc0kb0/5WO33PJ5vu7s20ZsZ9ZAVEtfw2PgLe8++ybEoBYMs
fu/RrE8so13dDqmnzmWIIaeOjXytkjvV9vLCSYEOTXPVZHfTt/SuDWw/VJ3EpspVdTZutLxZTwSJ
NF1lcl8iBV2Bwt1SuD0stVjrcVBPHa7cXBCQysjheT/qgDwIHXU0Ox1ItNdEd71V++AgktafYAfn
duyVr+eHAJDcVVMSHSYEuCjOZglndzcnoTstH6PuEEPZOaqbYPc3DmcW7wX339JDGfITFc2E+j38
LqJYzPu8nwIkGuAkPSkO3k/OscP/f+qUkl3G/ebZV+cPsFdjM1Lh9AVJFc3I9Bvhlrm1UPcZywUW
z8z5bSEkdm+FRRZ8le/T9z2qjQCam8cO/Q8L0II8M4M2GlU2f0JP78J0iMieg8VRStNaheNsBTDq
7/BpLKATlNvYnIgLTV/F408s7pIKVe/s1j8hrUacK4PaPogk1EJl2sRaMapewdZSx6nxnCrUh9Ay
wAibnSKdIDW8EQ0oNvWEvA0Y+89LmTJ5vBAGTv3XP7Qh/OXu6a/jWmu6GWM6dIrjluHymXeW3Z5D
fZ3l80Crw2HSFWNjI+yrpNgi7mZya/3lFCHPG2GTeJV8hLHUxpa4A7PG9VThZ4UhdWrBzFonqSbs
QGqbPdJbcW0JH8KNtmgS6DIOSqP3Y61apeRWuNNzxX+HD66dm5rXmlwe8OiAhkGAUfPhHDZkzxml
UDB/RQyYhwDzpDNXSDvtzNIO6pjzIVyt9+Ye9kWjPC5JO7rz6mK4zc+jUzY+UOcoPHt027CQm1S1
cGn+P72iFTouFp+0IBSsZHwVX/Wcfjrpy/DqkGS7DiB7JzN6PNpQwGaHLlwMiFQAuCOMjUN97jvi
9Y7goWrs7cKR+zwSa/opzpKfYv/vbyQx9dfIdKElR9xuvLgTJBUCqhyVarJaLJ+xx2fJe2N9PzlO
igIAMo40wD/LA/rz3d481ILWJkxINGpbcAv2UcEEsXsKwB8EfCK7Y/IRFonPBqkv+Cw8Mn4w8/dv
48fvD9CIfCSh8SlVF4BrJyvVpcsKh/FTbA+YX4osltRACcSMdXhxEsRdzaX/8u2ECSHuZImTiaJy
F2VKroQQlVLUcxMlGw2kHFr7Lbo17d2wIrSKUOW2jIMQMz6vahoOM/nUR+o7BH4VP12OpqNgtIR/
OiwL0WlB3020c3Jse3hnPTqjhvpVTH5BpoCCMh2Z28/JLbAmQWVqsGNkAV9ySRUvvGWp+q7jVJYH
i6xACU0dLqo4s+uVjp+qRzQKOdzrBhtIH0qQ6gyKG0QZr5JK943JEyZkmw5Q5j5JLNmuuLIBCyLR
4bE4MbeCoIAxo1VmSUZf80XD4yFf8y90wBMolqeqelynlcngkyziFbl3TZOy2WWj35r3k15pJQLl
9Bnv6YHAUDtvFe8bpV9P0Cyeeqf6CZQKlcLrhIDHvExTkr/p34QaNeqqfx4APVn3JrFAE1o0VxGL
VrCRXsZKzyZiYVwXQYqHOq+zEeFbdImul+uKYvcdFOAh8/VxBIHqOlZcupztzqpC+xJtGn46TB2y
5v0zsplkdM/5CAQJXgc5SWVYYLuIqxgK5rPcUH/OBlMeD57slwiiBWNOdJi8gAI7pvzRW3gVdrAL
6g6Yj2QRxa3mLzhCKahfMlHIiE/rNk1obSAoq6uQ4YI9ZIT2cJAel0UHPVmR+fA1z/n6Xx0U3xsF
MKPtVobx9QSLXxjhdLEJxdHSz80gSC+oqOT/87nb63VJrB8PNDGkOwXcDp3zyelBN/PTUVq6RxRN
mMsHZhltg9NMvNPTQFihdOIfv9MeEHteZf+aj2NLsFqLWEUSptRNIIY14fZgF6InYEHSyjViFH1W
PYbgi79M4098UMe46XxqVBxgduRTXCXWBt5B/ms2/yOUTEUjMCsl1wwq8+cf5XUf2Ah7+GOOR6Nz
swOW7It9IpcxYoo/WZi1N02GkVI5x4g8PeTrrTaIoI4LD95L4xYymAeL6nygFPE3MqSVjWPboKZA
doNFbfABgPEiY6AkQsPEBfBHJV/huQ2KF4Drh9xjvwD3RhzH3qeICsxsl7JBLIKJRi3z7Iiho4ww
CSj3LvRl8TkXcGE7Xh/E120wQPL1tvr8Z0OAsXNskj6XvpXHdPEUEvfCx5rJj9gqonp73rg9XBsB
bml2eC82RDy95IAlgIiyxzj9CGc57wyjo0WFUuORiCDpOtVevkBcjyotSFX5XICjRmSeWAhO3KIY
PRRIMYA9DIV/RbRBLJBz0jYtzgMAGOE7Xi4Z/5WfSGsM7fAGq/7x3dMnQfA7VK05TY7Y+hj4bUaK
sRJjilj+Ke9hOqr24Mn24SaS2eW7VD7AFTibcg4XhjCjZIUj408ITwtqM59mP7Ngg1Vx0S2C3UA3
3JaTsspMETB4Dyt9fXQjjWEhtabWrzDQ7zxyIA0RQ0WdJWKoSuPsXlYimBu6c4qtkJFgJr1tV6Er
xo8CWuB0jm4eA/bxzydBosLQ2PWop/ZevQm/VwbivS24PwWSr+Cf36hj8ctnogWR7A71QiEKGT4w
CHuwV3NIUHBuFV2Fi+Ux/uzAe/0hDLHlnIrjD52KAwIIz9TnOdBq9laJB2CarZ+H0pG0btl1jQaL
/bil05Ib0tj0rxZd3RjmNsOBmm6YKCdbMcbskUh1Bu7PyMHHJzgtMB6AM/1kgbgpd21MJnWdXY6Z
PWaVXWNZua8hcZNo55BS9hG8LtUUV07jjbY+iDEnII/auLlMCwlaaRdI3XBcPCOBRWjExbcvhOBh
EEIJOJNXeFfmfamawjddflJAaH9IQLgAlczs3zHNYCBilqeZ29lMUNJXXy6GqmCCFHtwonhXWgra
6DAiUCqJ8Jmca5KQmyLUlm8yOCiL8bHjR7AICylkgxREuw1br5p0VAl0SJHiYQvF4aXfz1Ubf4JH
EFA7LwqyTVBjE3BfNaEME2dogyjODrr6v4mEot5jWyMQ3OMNbQPeYBzANuVJX+xn/l+Dik23lEaA
HUoXmx6Kn/4nxXFtySMM255qD2mrHOfECRiWI8aSJAyih8z+fzWGjxO8uwSKPQ+01ZDsJnBa3UmC
2ygXQfwhbj0WK0FAAuQPajXZyWOLlS0UoQakxcr677rZyO9K+duL0RevHLJGJbBmx+11N08YYoNc
VfQXlQeDMCVP200lAquaAn8x516afLyWyeGKxnFij7xhAdsuHF8whpJeczUs2OF8DyZAiA4m9JAd
+p8gHsUxXOgpxDw24y71/cQw6q3+I/WxMZgxgCGpI3wel4GfsqHsQZMm+fo7mT1CSYBlKibsRXPZ
VWML8KX2adqivX69x6zuo0Ez38o3vmjruTHcDiZ9fnZtb8Mg01s+27fb7anvXdKDnJtaBoG781AG
M2WGoEKkDwPbU4I5THJhbejxPCxUEVH6CyORLTz1JfVndJijn4uCn6T8hYnFIBArCy16qBqF6PA+
hwwrs9ANdgVkg589gzE0iP19RTUxm2VPN9Xe6EjEMWjvv3xSar/A2bM9g5ggPUsvRix1tEnWtvIy
9PwIJ4n4R0gx7Uw13u954qNEmY4mBwR/COItXuXpPSQm01+7aMC2hwPh9BvVsrvhKzDpOaS1mYLs
Mibmjp9sZe3DNM1fDjPtqN5Jg706Jx9STiQS+GLuEdZMN7cu5iwSjw6dZYVipXWCK3Nk6hQeE/0N
0f7NYF7HnCi7e6zd4Yu7Mq4et/WUH14nz70vEqBnyv3uLn5ZChx0t8xHSLyKXOqn7LKkNuH6bMYV
8W4uc8QNA4WRaIuDNGDbrl4sTcvT7aZ0Jjl41tUU7kcGDkmlxesbHLJwz96bLzTB790NjlCk/JZd
VqNe6FJ4Fo+H0M3A85RzEBb8+0aA0iN97Do0ngFtI/PpYa6dT2KPaqrt7NyrIHUxhinmUYVQdGHo
aFfuINUA5fvzdKslVBzxZg0wYSSguMtVG5MCrRF5QMLq5pRN4Ai/xT2S9I4iLgyb3P+vGnuNblhF
bfogDAYQiKLoXA/WCOz9jcMByGxdsmTsGjcw+p7zelSChphSMiVrtKZ1Tt6NHTTOCVkAbe+kl9jH
PlIR1jDoA5SxxoqCH9VuPtuqNAFZjrfA3WfSUHvscYONuYcvxwfS9V03AypSb/6BXHHqAVtn7xk5
V4LUtsV5jhNOSgzFjwHjsfYe6kOawDxGc69hOdXX7mi+HSGBBRAZC0iMKrfcpCxmtcfLThiSTvmh
WykLL0WVs76Yxu0QlMlK41gmho7B46/btDY3z2rnRxTU4/GiPkEcbqxNBC6lEfbIZFJQYIvA39wi
Cr2a5rNIsHqUuunVFJjU40hewb3HpeCCRcpRn9h7+QMvsOkqvnvHgUxB9ehksDnhr5MRtuwUEbgn
2T5F/XgE0L42gM7QxmpFHKNvOh3OdMavnIa3CS4J1U46f+SHoyW5L5u18BGxu9cbZSMZ6JCne/cz
HitdPiDvq5xAzORKb6+xqNTi/N5AQAGRSoLuknDg/wyg6gQs640N05QRCi3xUJFMyg96PcB8j/fY
nL99Zwf+mJfQERIYAK9kflCjE8KwqTIu+zxETFnuOIk0JGvdHiRlkuPOUyf2ntEdCMOeP6ReHhpZ
Gum/l2TLU90w4Uhgv4azGHoDc0WMKo+fEozH6WZU4KzMXGjNXXZjQqPSrT5U4o1Yx1rG9Cr5uY7V
GcccFCkDFMR1WHeWhRSAc1Mu8zzWw6Zumm0Y6oTnW+Q4Xue2EipT5wabAfFUAVvaTKX+5SCN47lZ
ii6JbkjDggllwcINbxexvKp50Q4VsSeGy7JUmXi6PIEjM0CXFj7cW/pIrCGD1ya4R4PU7Huj0NMX
vvikop843GJ2KOG3i00k3muhDx4TUkpKbOOs2bC3yZ42Sprjz4xU6jewT8q3DCLAAnKuQK6qfuQN
goAbfOz4rV0Lv0DqF+k/pPchABQjklY/K4Q2nT0yD6IuJOj0PKjUlTdZVQzw+hGms91hxcGEDQjA
N4t3A6xdsHdDEpkO21pgBqtAI5Ml1yG3qsXJasVIADSpyp3PhQEvxRTxk2u2UGUET9BPhJCWEDdX
sUPPkT2rVqoOceRnstRrv0JitsGRjQ6zC4lYAl0WxqS+FZtqv5VwFnaRvUMptp2ihst8rCx9BfGK
NF822ja4VkKoOFg19sSOOnSVZ2KU5eFfpud8xDk/SkRNT5CIeuwkPB4tn4aA7wL+xszNUuhlRKJX
1zQk/ksCfPNlJZDz92qFC4P1pnkls++/XIeN1XhatxvYq+WWJmC3W51+nIjii9aYX/Bs3+o1+l0u
mxjVZc7F7vw/Lgxc6VrQg6urIbX0P3ZyJVJufRfEHVJAYzMHK5QxLtxZgX2Yi8oYUzpwgumUvudP
Dc1tMA0RPCJ90GrB+zAw6F+JvuqFaH4lWWnODYlunavi42rxrd/YN8OUigvw+owocR+JTdfGY/UE
sR0PCIBxpNgxThzv/c9P2ESEws+Fd9MOqltWUnvE4+I13201l/o0Hj4XvbNJZLRpGEJbfCug1b+l
dIMLinM89wC+Zs5Jjoy1JU3N8ei/bj17+BJzj50vNxgsiTJ85z/ZoEE8zLCPNqJzRrO2vdJgzuJx
dMeMkzGPyZwdXDbsN1iSFpHHK2Czy9ufxPqA0tl34Pfc5FJkXascid3pq3xXDSa+zEl3k3BC+VCt
6qMcKLnMuCiOfSOQT/4tqybDyfUtjnIwhfLJtXNB0yeet/F2N9qIywrM/zrvqic1oY2RxUlxfDEb
tDCfzV3ZmIQB5VKLELIG344wB2kHbs1QTJ1P/Hn1+X3OW7yiESFZ4fodGuNAfnqyBzf5vrOr+GoF
xYqa/sHbwiGLq61pUTC/g0qE73mf/eGJbppOS5VahGwTZmc8JGc5aQHeiFbZXddQ+MFpLDWfY34e
Aukv2tQYzSidXpQ6BD+WiNZzEM5U4wiWcx5Un5r9pI5bOaVMt4qK6AaOC2fu/X+4NiaMI+eaUENp
oz9wxyLpg1/zxd0aXulwFF638RY93kQZ0TeElLXrkCAmkfP5jVYAhO5wkLWSvjM50OYK4r7qUTxC
kGHuHa77j/pYHIwAvLks/axoKqdIB4IB5JASrtvc9aqxoW3kSya9o33zrzzAXDUhVYixLPs9mvef
71rni16KlSWZ7dNhn62rdallK88UbbibtQLWOGIpitUpCu6hm8i0TZK6xqg3+J2lnGmu32czMCZ7
6JvPrpYHmiUbpytU6A/Ia2bF2h9/Z6MNK9GLN1r1qPh/Xc/3dbhMYlBat93ZPK92hU9Rbtx9aDVB
NVd3a6lvTv1ODaBkIJ7OkcK9zljCZW1IX56LFssbhI17eU+NJQ7iWTjOgNyZOSrXNjQeOh0d+TNp
j1ZDeZBtDu3t/LIQ5ioab9+rKKa3zalwDylh4Utq8C3kE9edq4SyA/A7kYreXuedLDE7A9LqbWmB
jopgll1jGXxwxAYZVYHhB96z0YXzZ4eTBEiSK/ax7fOeovUbHZP4XLjmqPV5OW2kZrdESnQ3ChcT
IenfQbeLG3ozbDp1fuT7tqMt+jAbr2AFxui5PCd73lLLLBvQPtZx2y1JQmhKCEPMaSjzagWVA9dV
Cm0kFBYd7z9uZReFJMG+iSdPU+6iRtub4ScGLSIFc+PqMirbmOEaS3HsWFgo54A0/iC6kk838P5O
ZZPqDRAWqgPjN9k0rrBl7B2kz7ULCZyZnQnH0VnmepC49HOHuvNxUcHUOxhzM+GbVDPgZlOy04pb
rfCpW8TuqLUK/RKmcFJzQgU8dpJSL8MkOI+liPrvIucfIooCJR+5mS3lfbgRBfVNUeoRPFJ/ost6
kqEGpYHZDBDU9GvPJW8w+4rmC+5kEraJu2rKSa36JUrmTCeH/h6apjzM8xw3NZNELWX/e3ZkHx0P
qQqXeSrTR6xNXGnIKY2yA3wm6qfv9QNYBaxAe0b2DwA+hGAIXxlbj+UN7wCoDvmDASCr6bGjJ5zu
PX1vQcTr7WyTPyBLd6gAnaGofzUuF4YP44BCqQDwLk9wFN1+zaIWC7cuzrOMzVec+BFcGyTLg6lC
TV5raBgIdLsXRiHkmdXMhEq2aaYFagebN1Lmo2kNwCwRg3zQQafPY1GUMOkkJ2gWJlDSk3ws5kMc
TFk6zSZhE2f0jL8un/lldxAzn45dV495c5obektYUgxAC8KmewBZ+i0ruJazRyzKKIaGzXJNgUs4
FFto+RquhjrM+nBF3bRP/dkovva4uBufnjefsbNGnz/+ALHol1a93c1j2rmF6EU1ZCU+jqDYt5ET
r/gK1/5GSS0VUjYt3bdb7zzGwhND9PFhsAQufs3ZFm1r5tivGBM4OZTnKDyrHVMa5iL7JwR9VSkA
HTGdYCQgu+cvCkSwM94/DQm6klA95d1oguDHpMWscQbdIGgN1OTrqAGhx6Vk/FUVEnKr2vZLcZkX
dWXZiIQ3q7sfgWuoIOLIzJR+/CdxIwBo8KkXHatqWkrkKBZf8LTBsm30/dFk0+vaURYcVJCECWcD
//SSlA52TtpNOr7jjYl415MY2mnnMo1aPqdE28n+bKvK2mC0Tg3CZ9p1tl12xqLBnYpq4z55xF8y
YDrbuRkWIW4wIpnJRhykMy0Z54pwVYXiHdf5XA8NsA5JizJev5O9JMWKtucuRMRfi/+U0j7ZdyRT
rbvSY3x8G8xFETCp846jHFKwkic748yIAnRmbGyv8813JBnHUKVWQG/35Q5+ccCJOutHXRuayIpn
DS3AWnO04m0Ltnh34Mrs/ePq4sr7NUVJHgZ5PlUbpwGvpQ3xt99+23AeCy6W52QMS03bBcs9dtuN
3QiO8WIbiT2Lc3Fv91HoRAyEnWXDY+6XSpNQ0LeLVUOGPG3/qsf0JkpBnyFSJCuBr6tKf4wV8cI0
hCT2V4ZRyBQ1fzQaZJDUXzSylrCwyMW35Myl4CAc1uUfdtd3mTQNckQpZpLv8eCRFLYRPvoqrN8Z
cvBxMTFj7bf3hIekeGwitrg7TcJXI3W2DeqoMft08GqD6k7/4GYwIAyXfnKmdNJ0W7813hjN03wU
hShEMMWW1luh00n8xcw7fpII9s4A06pTE4zgPf4vfVkXki6XBWmCqISlmt000sW57gADumy25+qo
fec1gkf/AE3+1cGDLZqMTOStQo9pRFgftcnG9srQrTxc2QC/yvYaDPEI9ZNYfInJ8ZdFaYSlFBxM
BJH15Jfw5cwI6/GQYEqqo7cszoH2h9h6X0aEoVYcUh6pUOxzMuSpzi1ZGdOIwXb5fVWj5BnKYmWH
0ZC+wrCIkO0CH9gcKzQ9OhZARSxEE2xa1LVaEhvtzwtHEfKv4XGN9/QloDWhpo55VEb9AOS/RkUx
GSFmi8buK5bqaOwRUdOPdVEPAVgOytDL8o/lLpmMhP/FvzcXNTcj22dR/DHVGw2mlaHBbmeP1BFM
RuoVqkxaEE5IBq3Qiynle+SP/rXoLzdFkQQiN0wBlorqudp31dK/VEVogmFQ2K6/lHBJfSO70vka
XwjN2WkXeuAyICDMGVRAcf6kTdL6prDeqV1Zv2ecEAlfaO7XCPLKxY+0UUtJqE0RW+xFjb3Hm/Nw
dI+vC7yfnS5zAIOIKDADuYh51do0FwfpINRAk2lbT8SZmNZhCHKZXfRNogqNMP2u21zjSLoVFzwo
4rkzDJr4sGjdYD58EqKCLPh93rcY9Yvmn+5gr6C6a+SQ09ohm04Hz0uc/TeKIDLK36SkSY2K8hbD
n5J7YP4ozDHNNOv9Me3GhzMVjM6V1GWKZTzEJiB4FH2cGl0Is6D+S1lrqMu64N/2oipAy/PcsuX9
r7Kft3Sj3gIMP/0cwKl91FKQvVx28XASAsk9+NXiRD9m01bK+1f/m8KAc1w4rzqrtY7nnGEFTvOj
7UHIoOoLMtmxhtJ43pRDK9TaQzeXGSsCxa4HJ4TVZM+mFv8lhKirqpb+jI3OWCWPWgRdOZkl3Rrv
P+nG/DlKHIPLIbIJd+pV5h9k1Mr315ngbyG/TtN5W2K+ZF65KKP2jj+g/peYy+eCyT5FRRtw6JiE
ae3stMoeBktqGSaBVaQ0ckhEs70M1yOfC3z9n7VfBdw5tcP9OHhhy4J28unZuP1VTeXEelms9pAH
cl9t89ixpGZPOZT4pNEV7dmXxDfKNw8kCowPsOwu04ksJTFAAHJrz7FoNltqmRRKTBIPpGRHfln3
hKkjC6qm2HGRKh4CfgdQOumciOOCLn6g5kqMLeYew0HScn/d/8yaTg1tM7C3x5d+ATngqCLMwkCK
RAPr5FJpdMIHpTiPNFM0nNJlgibwlOt+c73I8KOkiTUCe7fn3Y6l0ZFxc1sTy9zbLO+wfcMan89e
Eec7kn4LDSh5sPvDr88zzi2h/nilEtfqde+R/au0/5FIUEDxNJzbDlpOylioRRMaHCqSGLv9dJd3
aInIxUYTepU2aoXpGLHrVikd1shi5kOsAzvV/p0SA4Wmqh/UUvYf2ZnDxAdRmemI7mH1YsNZ5CLe
mBXePQQPWsxT8+cjtZxcne50U49JUtVikD/1e9jifHj/QadFUmDPISM7Gld2T7XdCVVrgmV1nfGo
+E+nZirjJMGpOU9VaSJEbS0Hx6x0z0qTL3lwKJUN/GlWvYhQtDj2TnLLVhKS8GewyLP9GhrsEVa5
XcHuBHO58mqOZvU9XJ9M2esxexM8rWNFjs+piQOUpuKnOWU9+Q8B1whB/qew1l/TAp18NagptnUX
gAq/vcRUuQw2jI6rIAeXzewq2XecH5p/LK39XX0xweDdnvI3LUqrg38bwzOAaH8ey0UiaXP9ZOZc
CPTsvwkqLyZuiHolsRzmJ+9jXbZR2DhxK6QOFbgnBKghOKSwuhswvpeiApvmQ34VE0sBoUJyrtwQ
JDgcYnJEEf35QVx5lpA4Y7CsxYkm3oO5NeOlB2FrjdWzDf3LeM1MwLF88wELcnRiHexJLqekZBQZ
U9luwbJ6qZ4RE8G1BUhAWXSJYdA8lrvjVvt4CsKE5DIal9jD+GX17x9p33JfZhL2ZytUuGDN3kvt
Mv5oyUDKQ9eNpX3C+Y6nh3MslF+mOEop1m3lTchyk8O+IhTIwKFzZNCgntvPs/jNPyB2FcPpsL2b
fkme4tGf9o2v8klkj/HHQHFA90+MGv2NPT0QErkJ0Ai2e4c85j5sIjPZvd5np5lgXmRtKfOunyzG
qL9nmlFzepd6U+u9SMbtC0WkQ4aNjR6OZpQCkeo/AQDlUo+wdZNSdBq2Reao13iYgBOEjGYm9gjw
0hkytl3Ct6mJv591M1wewL+qqVHmneRwxlzUJnWXLVMG6FE2C4R24TsWbwnJPWTO/7Btk8TWC/oA
hGB48GkSpcCpFGtIJ1snakxLwFhsZAm6HQgYcwbSrarsY/97cfdnFFtpNxk1v96Xz+hGKHjwYJHU
Eg39c1sepSb4RhIokQ0CATC1KR0kTAe27W0+KjWQTz2/Ck6S0LY79BCwwF2BIulfjOI2q/8nbrJI
NkBkSS4XgkTtOqcqI0yH1N1mzh4kUWOv7MXkDH0xC0up6JQZorEPHpVNsMRx/+OCS5OebMamolkb
qxV/gVD/BGd9JsHQO9Ovk8vb0/8LIIf90VucPA8/0lwSzWdMHS5CHVpznmP9tht2GpOTAO6iOOZO
cgPH8vI2dTdbVPtZan4bDbd2ADHBIQW6WBEExR72+LJCSnxfD2Zve42j7drsSFagUDZgMFQSnn6W
zq5f87dRpYQ4z/+OL5XRybLsIsADqQ9Sr2YJH7Dyb4toXAGB3z86/4Kk3pvoCsP2HAYmy+m/t9Bn
cYB6uwOfMveHuiIVdie7FCYr90Ai+1/iYldVn2pHbZ/6nmIIrj2iS8CQvDGD2Y7ytwptvVWLWgrC
tkbagacfhM32cOfqbifEMt2ZqYDsJ38Q7jJppL+OFl1ikCue0VD+fBPndGJNWQ4bnzOlsWxh4gQE
x/PqB4ssWm5o+BESY5oi4dlNz+VWGEKzgy1R0l2ubA3GmaDePloTszfSD4NOnfFg3ulaJ9pGElJa
2JS31c7sxKKi1vFW7O8BqeSsVB5iGsDSd8OT3vm0UYKt8F1hVwxes6MOquCbeuE/S+nwsqjNurwb
6HdAqygMUWRw8AoUA6T0r5Xn//+xLKvjl6yATVpa9KZHXWYdfpaJS7eOaZSu97oCdSUdLuEuqLrE
2doJyI4+H6Pw7dDQBysIH4zu2VrACcWBcXqF2JRWhHEqoF6A3VrGjIYaF0ftC5CBIAW0cfk11mNW
fXm/aSzY21uwSzwxfQR6zPe9yt9WVJX1cHUwJt72iK8Q/HVsO83Og2l1aaCY0wkZkH9Rnm5exiAO
1yq9ngHxMZcD9X8iOXgXDf9lkJyS5ypTjpALxhTBozzxFybky+ZXG8+18l9OjGNHs+wD5s/rY3m8
CfuJm/yyL6tARjZBjO9PeBIMVleuRquGPaRWv184/MxrowkbPl+0uN/DVBn/S6wSUaogmcMVMkz3
5nWEEcNPkBi5sQUDCmOeidJIRB7oQAkemYqFBfSzSRZeu7rCZUatHiE+1FtDGo+tCNOO1fD0cV9H
oMyYZgeV2Kg8n5qQd5e6SE3l21ZtSvwMmteHRUOxEy/KYJHX8ecPg2JIicVZ9CjiVH52gTPHJCit
Z7Q2fKNv8XpfaJ3nAIswgEeWaBnF8mCoQ7z1YCTh7wF/2HunmJzBltZkSsJNn1KbGqa4bdMZCwpr
wGXB7N77dlhDX/T1MDH83vLmrIbD7BEvFig5BJEtoSzMnxBIB4azjlD/zhxD30jwegNfXSmiUOX1
n6bauWu6WeBxlxg7mpOX3lIoP6QWUsdX5ep5OUr3Zgmcz4uKWtRXfdGUTcDtuuR52lR8Ue/Mc03t
IICqIR3eJsy2x3GfZDCLUCI/lHEhIrPpevGi/Eh5ODmxdCll9y2v8brGSpDQ1zpPLgR0aBiF5BhD
LQyuxO6GzfGcoAw9wSqRt7ZijS367lu99uCUBtQdt6sAvYOzhmVJGbp3ducwO+EidEgpurAixGUe
5Kl42imC6ppL4YPZL6UAa5LSSgvX2Zu1FfWu+a4ozfki8f9X385I7LTED2laCTGX93NgZX5FCPQ9
6wA/R0SqGp14u4fPpOSrlqRRrgu7NMZwFiGtTsZcoJJ7/APEB14DXtwcuj0/yEtoXY+SJ8zOPHF4
7tLztedzZS8IH+XwBgLTKoyIVlIdI0axaCyHQB27SttEJh/3ZDmC907BmX5BbbZw3alXJFNp5FRp
BwwcFi4919+LnpftinoKfdy65lhW1buZrD+orL7kNG8vnRHCK6LkU0yKutrKslL0bOcUvMFeAbl/
ukstrCL/IXqYNSmlhmtR9U+JRsJbHUyNSAMbi6oPw5odOI6i7RKreYvni24OPP2y3GHeg63LGVD6
pLlaoJb3QqtHRP30sH73IHyNxKIR4Q/9an80MzxGIR0ByezbuJdZscrzdxutPHWyMx1fdZ5xsNxX
3ZN3MO04TQNJ/gbVXm51rfF/jypAgF/LHkk4bS329u1y7hszCHtwRGG/uUHcfRu2zLaADz+90zRT
kLzrCBuw9cqe2Zav0w6jK8XIb0vIpZQJ/teTBvlF81pnDDkpmlMvQW4af/CjSzBGmVvHP2vl9DPK
0w+feOjfd08HNN+3uJLDMDceX0FKXdQGTWavGBZ80yC0iTiFndFQPDMcWcuYCCXLYNLos0AK5JL1
ruMyZTBTChONEl9VRbkV4Z8Gn2thX0xrr7vgtX+tl12difiPxTO/JaPWf5LxRbSgPiPhmdekyw3j
3kmqlAh3bRfoy2EK8LKJk6w4p5bc0A83Q8Uqn2GVHrzc91sRh9Q0jhMAycvb0xh8GS2UHb7bS8wO
U+UH4Exo6XdcG5+d7CJWsI6UyggewlG19LFA6zIisBd6zVhwhW66sszR/9V0EfqPLyvwdqJrNUGv
TOU7kcoDIe7BSQHofzOlM3qRwDc5U0hAx2cVKd60WRn6t8LVSkEFgCKfck419Ok70a1N5k4zMjIp
RBTQqHLJRjxjxhoyUQmGwCZ0dYz8OAYslX/IBi61XbpS+i6mitr7cPMXZgVP7y1HL51g76EFsvAy
bXWPEAuzQG8EnMIpH7+E6OAl7FoMynDNWuJY0sC73iltpddBqS2E77GJmTa3GjSmOc1KLdI4E8v8
tjl7A0Ec6x1QL1c2bbja5/BjRhzLeAAOWoa3tmkXgXG0ChmNHtnkYSriMGy8UFMtht8hAp3KRItE
+N6FYr8xCh4Jg/Uo7IGSERjMsjZeomQLfwesyMcwG6V5L4OhB93PH1l6NjKlw4TOesS6pW0KmI8u
lys0VRg4kM2PGAJKv5q1HVUtyGapZGOeYHag5y0dTdaAoteF2W+Mqu58qTh9uwzEzbgAj1+REEfe
i3z6CFeZsaUOkHnfjVCGbseFP43YrV287nsKKHfaiBh90MMDAHNJQXwElbPVffglKb+/IDyEftVX
ho5Gtd12hg8l1hfnxHAqJp9LXAlxwbuf9RvrBI43rmyluay1gAKwfXERZQQ0pZ8EbvKrQzmdteSs
2R4XproC9afnyi45bAZNUvin/tqsBH96juiWMIMqulnBDC1nvYuxQxZS+uLs8Oi447lLu+sv95A0
/mMkf11YlMJMVmdEAT/OTyHK5WgQZwnSqJH4LfuBbNB41MfC2hrpEZQdlaP0KtIQVBvqzsXLjhN3
GxoISqoQOfkuYXkfE9/xuhhMJs4xHLp7RqzMsl4n6H669Z+KCFX08EyvD/+6LuoGmgq4Z9IneFSA
GDrtxr0FJwNnPXJ7WekSsnXyvMclmHdbaPaTeFCmAooAFQskB7hHggXFXClHNcBsrDR7QdxVkdkB
N5cUWEXbjP7uY0VawVkrrUVA/pP7VOxk+I+DmqtInXNpjMDHrbt/ouoOoLEkIqDVR2xRbHVY58Lc
IbULA+MCjkKkATZn+mT7AsRgIpOIdbUx2ZCTSa7ndjPr+reMhmxDiyv4ExA0t4Tb6zPzMpG2bPRZ
EZhQWnb6raf5J/x1z21MbTCAugQYNx/zDtmxF7CSk4bUpb7nYorON/37paxmCdYcYABf/CFELuwB
HY1FXpLW57z87lyIhoBclQQ7MqmAZdJa/8Sj73WtR/9pEOQQ08ln0iRwJKrwhAFPToPgAf4li6KX
KqcUgB1Z/ouwMEIYJkomvaoBY7LfZe9ryxvTrlPFaKqtM2rcP4A+8VdV738vizEzrhkYt2PEzq8R
lMG4MiG39pLvl+goJK38W6j7eZsFvq+1pMPi+b4Sw5RJEaYNJtlaxuBvDMDJgqig+ZsxrysHO/12
2mItmGFlxrCcPECm0/W/tQIRvC3zRU/sxNQIdjEspz5dRIrs2g+614wEVdK8ijbpVrhYJnUvuSg+
vhot5i3BDDwsZVQ8DOYFzmlPUOIwAWjE9KM1ubLI1z/hnUeYHHrsncGHQzA1BxUTpkddMcQKO4wx
iEgW8Pk5/aR8RXHdxW9CPB/0/OCF/e/yLVkdVcDHNsGt+3DxhF7cEEZz5cKKyC5nI+rMEXRsze1j
2VLFzPYEFrWdqFp+WsFnWbBM9SfPMHCmSsbuRRiZ+v+KzGdGv1OHJpkuXHXKit55WBxofKI3dVXK
3f3oqH/MuWAyc0IRbSGcVPxPj1P+WpshD1FxqgZl0PpzTdOswwRKNld/lEG8N5vi3Qkr0JkxN/xw
ZlLGVL0KVUyBJVmoE8N49MaHk+ulK+hy5fqiTare06DEtBmaqqCVV5DR23IsjNjhni+qdC46saks
Xtr08TyiLxo+SsRlDhHfTKv9Qb4eMdW2u/nA96AWAY9qsqB1dEUwEfZLZHUqTu8t+mQ04HzNbi4z
K4yNUSr13PBEGjmBH0LGU5vVOnG8th5kvKyjdq8wmtgpFheMH267J+O4z3q5v/TkWjRG+TUdgBsS
cteUxIrUyBP8Z8jD3FKc0zzFVMewJs2BNzaQqFnxyTA3q8fkUGuL8zUJwnf2ljnMdv0zaESWT/he
yQ1q81VkwD1jQMxEytaiJg1nwkFcbMcXyK8JvfPXp07YdR397kB64czKFQepJdOG3Be2YkGHXOyA
0hQBPebNmnOWthxCAL3BrjHlAbp66qQWT+qlqcdJWqB22yOCe5EnQav8NA2qzG8GUj2lLVVOs0gO
qMqKxw87Cturfu0=
`protect end_protected
