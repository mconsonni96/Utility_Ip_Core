`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
sGzgGk5inMbWvFYa1CTgigoQViVmopvUFLOOCmRncKkvzz48Lpudh1jvyswJKq2Dwakqyz2lu6JP
SGQXC0pXm42txHxJl9JAml0MgSNM/ynmDmqBCkhjG6GliFUgKf+n97EKDi1nDeYPtiFs1FeCAcAQ
JA+/MBze1ZtXdX+E5Zc0Ifg4fsxncoTJGf/cM3GBTN24kbZU8hFM3KPv/wBbn5H0dZOXrsTWArr5
LLSWn3Dz0R4dnm15xu4EuJxDw3GFxDEoW1kGQNHy83pwVeHuwOZkoOdFeahieMyapN54JWjQlBcs
NV/cZQw5gxJXvArVgDTXjOYad3sPZOwGW8eRaA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="qBZ0GuGfhEAgM5gjj+qy4rZK20JRwx3dV88ge30GW6I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21040)
`protect data_block
xWBQEHYWwTxIjQ5Ln2XPI3izdvKfZ+WFFX4SeJpO5kqkZaTn0C4CdpN1WSvHQ39XT3Ce467rWvVv
iUVHVbWA2ALYTM/R1IJMVi9/V3YqPcKaV51wkYhzhnbacLSYcnDJfgkaKX1tXKSxKndWuN2lFeqT
3O2qWD+FRlrVyc9ChXdJ3X46Ldmpvc452Rcx1bvuGl63E3mwyhUf0IZKNLFc8wh4mKWCmLF9qYqV
pBVqnyae+A3a7bZq5EmjUK0+g2eIatkES15wNTV1UDDX4pX4fB/IlY8LruPvzRZD2xSCRAPR8mXS
4+K/iANGs+sj90yx2hEf+LWnW7j0KuXJgezT5V/A+i8mhu1tJY4QaHaJh2ShvyftrMO0rr0T0+Cm
c/xFCuHqKBSl4ekLhjkiFq9rQlAfd/oAD94j4QLB0q5r6NPaWMXUedzTBeDUeG3SahxJAVrJ5JmN
93Stj/WbUpTd2+7ZEs5iO+D3YLwMbzfRmSjkgxYJr2409U+Pi2UtmGgZZMMyV+hbNBDqjmyDpnfS
5fK0AXDlOccO/CfRLobn0+Xt693ZkAk0FGy2cnDpNTxF2EpahKmI0oe242//bN8jp0S2hWsKjeL6
Pcr1iSmmsDUK/DIb0CIIaYuLQNIqK4L1n8NtBRUAIwLQ9x3IepKVDAhWps4KhKEtPlNmjtNkCY7c
EKaIHI59mtJPgijtOUvggMtBxzYn7c0R33fdAQAHqoXZ0gzVIIFTunzjtnjxSidko5Gd7dV7SmcZ
47Kd/xTBSs7ZTla6K7rQ/tU3jpzWWBdEnoW1rxodFsHsomQQhIreC+XubK6d0qcUWoWBrbYldS/P
1FTG/WvApM+J2t7raAgLVJaLthQ2IKWotdPoIOwtzpdMVmyxIjnQcKJa1n4HhlOs+7/tn7v7YLWT
CbkbgUYk+IJ3vis9/9qLMQbQVj7C/zjIWU0c34EYkJIpL1I27AVGDFvK3r6Nfe/f/bNfJuZAeIED
D60CF7O2ysLbc8VIsEdBXZ1k+CF/8RxxImkPk8VfSAR6zIWVQJWMYeclEqZJdBQ8PlhDyblkYHWQ
Z/GEKKKo87/PrqwwlU6y+t23XZKbcjLSWLw7wLZH/FZcKCtAkKWCUAC6jXPNzxKk5J2owUbOdaK3
gdjjUJ+IaMyOoenkksfSUwX0vujXu6ieaAbcj5C5sy9NZVsPZDObdxIX8XR+g/ZIvqLwn7BKoWCk
xqzRh06FFhVuqPo8XgpUkVeYr2pFYqTWGZS92yWW7Y8kJ8LjtS1lAyDs6N4UImncMdcUfSwV5SnU
nccqD5fd4vWcIWI7jlL1F5+7D7iqvIjtsBPHOmnPzWUMwHshlKg1+f4KxwWC0sMP8vLDtBApS/no
bMUWUMLo5XG5cGPfTHwSPMB30HDBGTH5h+BdBu0A3951Q3PeTf8sythAAfOpCQPyFCc/8OxJPNFZ
8X6qhewL0/oB04U52JN+f4Jn4AJBcxEuCIhjbfm7LEKSIEDfxRoq2hTFtbqveihJxIOcm3dPywvj
/bUU/6/qpQan5ElOvzqfu1XrCswS1l1PSfvzYSRNcCuo/Wr9bu+9nB0/PrLBXJuW2qBGZKy58tKi
/hhjmXvdu8qnyftZ5unxjK2twbPkU21/hobyi5occNyKbODpm3oz+SxQ/b39ZoDf1nh54kG0dGUx
SE6cxNdYtaWzP+eQT868liT14TnQD8ZU7X5s571ahLEiUFf5un9vVciwjxiQKO7MtHmw/ASVz4JP
6T0ZTE61ViU9wmXb4QU2imBur6Kh7OP2iq6Kfy8hU0CApwUud2CpkC6UtG+cl4jimvZXt2AeTIlH
/P6M5fVqsKzRQaG7tn2s6fq12hHMdd6HMIxFTyBd/nTybgBugVpnRcPkNVzrg/LBukD5zFkTeulZ
Q2jICtkALZ99O6csEdkDPD9nJ6S9nFKtjYGYVJdRPIJC4oH6r/Jw6WvsxwXbhkCbzPOK1jDxe1Lg
23PoV41bykLsDwP9g2apmDEpH/6h3KFodBcTsoguTozcI/I4L8lcIH9/sDoxgreXrBuEDPhBkmc7
yq5G454DHleVULvvZq6JahdbtSIDXO+WRHNUJHs6fMZwf4vXHdc2AHXlUEhd+QqbAVmY64duVn92
cgBXl7VROZrS4rgDa8PQr+JDDBRZDe9YFrerFIw//x71gILI2hjVKEbyC+epRo9Fa+OTpSOh9AwC
C0LzreeYnNAX9sMq0PiYEI2/neY2HKCC7NR+khSVB1iepCf8q9LMPLW37Ol9ozsMTfkJ1LxTdJKD
pFbI7IvF3uLBQAQCuYM+23/QOAQ/5PygKH7OCFk7Q9WdNroav+2hvrIz4Xjn45J7LCJnASEpd5Tb
i/YP4sO2YFGgBhitb576BhItRvQ1l+gHFdHUOYGS2g44D0ZynbXfWNMgmIaEDNyMd5YhOmifpp7I
UmOFnAERvv5VBEaILgnI/bejfEDzxQ/FmCRlNHomGr+xaFbSNKK31r2VrNS8UWpNUNP/7K0d3JIe
wEfAhoU4o8XKMbkmZlsPVX9HgXc6FljVg81dOBGVZT7UyQPkb3/9FkYDnuZPUtytUjS7fk9MOspb
3QX7XA/LT8vudv0GAZuEgbuUTpvDYG7glP6FpBZkHQMJ6gk3lY6VUopcTfxCpWWHLyc8JjJNUJbU
xbD77tw9wZ7aZGpMdek/inU2k2tlMEJxYyY+u2E8e2dJScjAwebysp/VRXjnFYX5SoiuwpKKwuvj
gZYNaqBw9rnHJKa5vaLKY0DU00JtY79LNsK2QyPXd8BeoP02XcSvPTo10nW8NggCm8SpOjAuqzYx
5uFAwkEk6nSJIqBAj2Mp+qKeoqQCMLbLA76AZBzqybflCJkd5Azc7U6MAE8DrdnYe4qn5bOoHb57
qOI6MzipDrh0j1wAXvJzCGO7nSIyY3T+AX1W82WjHrjMz4/Fv3GxdgLO+zJLxkv2xnYn8oEnsuMK
DCY2UxrA6lUhrD6ZSG7hLSxMjrPoVZJnAOlysyVPC4TcuaSw6w0SJBFK7AQvXEXn+4fC9BGv4ET4
De69H2q3U4BtJz9ohlntYtntL5zUsrPIaj7bbubmjTB+4fyoBXRSHNMPqwl8OtLuLnCFckd80Jdb
yJ26w3Y5I88Xgbrh66klSvOpMv//xMuek5d3DWyDPjyOzyMWtIO8+1V+1wmS/rzi2YvqCrJ+Jq2L
1HX0MHF4LH8fXGc4ppFOHIKQAXwUish2JxVq1tuOhUrJ9BPfuSC9s7VCwchndwG8a/bQHz0oeU4i
lPQMAR32oii7Z2vZ92Txzvu/MgRUcfUORjoMnHLBMy67hBWTPcIF7PDA4BcQSx77DWao9DqYPtN6
x8OknrPrjrqgzTCNMXuEMwJS15u1lEsfW5e+lopqCPfzET21BmCiDDRDrb4OApyp+KgoEeF8bHwf
FlWoyohjHHN2ALyrGjCfN1FaY8+Ce9X0Itbi3cfkl6NXHSeYp2I1F1OhAF9NMhRF1TIyvLMgYt9Y
pHnWjr8PZdIvWc7dUEGNW6m6o7CHv6S3ICOcCc+IJSt9B2n8tHPITaLp+pF06j3/0e48unF4H5iD
+Ufs+sJ+00cPf4FCfQBfdDLSP0a7PXBtAcvIa6/JSw12qtAHQAYZb203cBEudoHuPeGWB+WuxkuZ
qqqrYVZRghy8XU3rKj9EpC+UYPH4CB9ob63BJY8k6LN4pDZIk+Zaa6jxvD5QLr91wfwwNu+ZeeqL
y8Avxmoa88Ga0BOwa8lodr/ObQD4ijTA4bOahOw7iQJSe73Tj3IUy/euyH+RU9q4JzZ61UbzveH7
ip7jn2xV0r63DVoss+syO0Yi1ejHlpbuXiQOasZRapPfPgkTnV3Mq0mFcXwdswNZanh+IcQcqKk2
Q7YqMNr/4/nQeolEFEZhCR5KFfzRferRuBqxZ6iCrmGIinfxmi6YDGTR4au38EJhF5npzvXVp9+F
w5egDLOyrP5Xb0uxVvOOtq+GkIDPEQUn5B59yeQJtk78Cd4Jwylu12g1NWnqak4MW3uX2qh3tqI3
M0qAEq8Su/tK9bDargOZoJUMPWpDVYta59Y31vcY4tqB6flMHahng+EZ5Ye+nhel8og2Cd+pKHrS
N6/mHLK0F1pixcz/lyF2JpCmg6VNqRD86/LX9ulpzJ3dMF2WV1mdyxQ1BtV7hJQDqM6aBbYOsphQ
vAhFE0DojqeAr9crRwcYOqCSmMPbcX4osxgBV17LQ+vds/Ev/x20VVR+oYdZRWN62MOqFrAA5KUe
z08vsBQUe+oMNej4xLPCnMJeRudn1PyHXt9Ua/5tZfuswh1ZqE00O1xUvhlKli8gqJV+HS6c0++j
Y+MzwhTqsqclPQWCZsjuskR7ejwE3YkbSyvbcnRucGE8GDgyweUNg2lFkFMpeG8y4WqPdpIGEjc3
3lhCIRQ0NOLm7WPmtNlVZTH5W6PnfzNLTmKSKifiiTDir4AeSDIEo+MF1BLnzPjsyGlfE9cCT04J
0SNkrlFqs5POKroSzqE5BwmHIGzw/cxafyD33sfYNpoDxJ+TzF3KGQ3P6nSzt/NeUSMGM9xD5cgH
9vo0aFexjgk4XmVmmsvgdGs8w7pZKYHNIhJ17+VxQ3/xbYa82/TtCp6FS0/an2cxMktXYeQqCAcj
YLy3VlnUIOu7PBaK7z0Hb/LWC7oy3uwu/rqvgbbOUQC4ycxPhsfYkLU7B98qP77TGnQ4rpxDT2B8
7ZSY1k2ylXVHDsHph5OxOqpa7KqUzlMzUV9Z1Gcrxm21oqAO/teuT914zrqdT/6E4NPJXCyjusLr
iWZOFNKSOvTtJgRT1M/feUuLJT4ieOhKLCP8YywG0bH4JZyEm0b1f0uRyHqUgwHlJof3+By089ld
ZaSQ9IpHEETKllFCYxJ/4kiinEKLlpPz7+JHMX7evwWXlrnr142trVIFkl76yFVwTheNGKS5dmRx
8qxkrgdHhBVnZizUjYRkYIiw4Fc+xoUv2h5kZ+W5hfR6E8k94ylxDKUs6m2Bduwtc2+byUPCJmTM
YXemLII7OWPIoponIAyGixV5QwXMbu08Z6rCn9DZptHlqph20njYB4SWj6SqFvIOCncl0wLQ05ka
FS0BYKhh6t47wGt0EHNxsf4ZFuGWBjAD5P+HGbwNpXtzdkVQ46l/7mNaBF8JZNDCZfYzsjppzOn6
1vOExnODKIo8KWE9/YjxGXJ+s9S5yCIGksamRGbcqc2WOd23MzGpI1zJ5hOWHC6bZwqx4wk5YYEK
WuF6lIPbpMMyftAkX0nIA2D8uixHNZ5UEyd5rfJFrXUJk+5SQ8KMNUYOPPAHNh48za4wutN28z1l
fQPvcSy5to39DAfjJnZVtc2FYe28fPlOYTldL8fTp+8yDrVae/myeScyDBSisfoDHCF/Pr54+/rK
5ZGwKBL5ISeVS1Dhtb2ZFHhwT+VkAyyCjZsMyseNUDGl802Cyd6Er1e1PLQEK2N0ZNrsDvjmCAf3
X26HqUFAs6Bg1Qgks+B3dYXrd1mrlHL4l5QiibhRagHEiGUpP7Y1b/2f6CFenNO3s9EiPP7Njluz
u+xzhXLkPQ+j324f5rFxD8A6fc0JfhjFqewcfoRz8yZrKYxG3S2dx70xU7RXq2PA8xHoiXg96DrJ
MDEWQ1qcqyVmFHj+hePNqNTdLPpbLbzoqBFo1XgJE821ha2ngjL/y+XtRwQGIO0O8WbTRDTybX8e
XQ3kN10Z44vIhjqUf3+jAjCaQE1pOdLjFNu7mxpxJOK5OGZssfk9JkxGg+ggLzFmoYOiZ5I7QqtZ
JQY90ZQeauRBrFbCfCz1YwM+H82saleRT+hkT3XSaNixoy+9I0IAs7Y4UfSfzVk9zN3tIaNl9Y/o
oC1PjFCD0OXCayTCqubMh5I9qNm7VXYF7yYjPWQI0ujoocicCPugV8Fe6zAEseIAwBV5zEWQn663
KnuHDnHH2gqMLO3vQzfe8H6k00wyo6Jn24y5Ces2FmXpyMTK6YHxbaepJPjIjxT/+pybv9u1blge
ex8QfADDuArINY3/01WzlovaNjEPRulhCWbrmpk4SSLZLWTQP1RrnbANXa5+Yp5ZzwZzZj7l5wyh
Pw3xbXD51ya5IAApGqtnpxbsoHvVt/thjPWgeuWXWRQ2lRVTprDx9pxszbLoMMLRtdahHX1Sex0D
rIX74bDHI/NtvrlmL7ng0P001HOAoXy2e97utRHON6MMpC/qNwWLTyxcCRnPwx7vveuZcpw0krM6
LZf85VusiinqejzDjnrNclr6btMiHB43ZbBf153QyapkeSy67HolNH2X2b4jPU2KQTdLt507Ib7j
nJKcJy33VQo48pjFeSaSHIAWMzOYfv5wJl7kPdHQ4rS1OHdOLKWmUhwP6YBwXW6E1rPWkTf6nA7A
S9xhhoX6jl+0LLfnGXCuFch4MHbnLcvgVugaSmHVzr5wBJic7ghxEP2BE/uthb/CLstiYmSwA0Jz
JgKawe66xTkn56vXYEpRBeW3RDe0c08UO+qwPPOA3zwCesDSvvi7XhN5nrq8XHd0FvoAwwOFByrL
CDzll7EEU9q93zLKQKt2K7rBN0sSfhzmHkEM/LqEidpQ5eghkdjNoSahWJmnyQWRakjGpYVOWbZT
LtI7EqwQLMA0F56BfayWndX7hkWWW5BNXOx6cs0q+HnY7GrgAaIaENt8aE3tdh/tsER2rxxoIGZy
k+nNpSC3cY/1hglrqOFx7ie+zWvQveZGRe21ETB5OXwZMYPoN3p3ErLFLe7QwsSLRkNGzWd6JV9J
l9VIAlVeCVWD9JB2upDMq3CWvk14jLPUOqC3P9fMjiElXebuO19y1D6xVruWh/3v4cUnlHdhDW6M
OXJ5ktrystq4REDkkGRyJmg4WHoBptezfeRGSWKBUVkAmk4FIJl+aMP/UQnBV5WCsSs8K1QwtK/b
Nqm4/ihV98nZicbxIkCSPJxJ9lhbolSNvcAz6vF1mH4pgn0KtjvaE2saNAJ56XHiBBwiwvtt1NNL
pdLJRQ9DYk3zi+W3kPYuztinhT3nSVTOR4eZdk+Qz5EVkmiutj3uB2PoGa0F/j4J0rQHqBgR5HWG
svkOZ8gH7AzTWhEQqP2sWwWmzLYJ4QPszjoarzWei/2v2BrFz8FtG6+bVNuMj96L7dVGU80G7ugn
01Zk5LkjLcBd0fl431fH2t79Vl6uQB1YF6njD98eMHO4DpBdYhcJVU8UDEapR79t/2wvWX+jd4EK
txeJutRJYv1m+k9fwoTXtucfoCz58E0+9CJsz9ZOWl8D0swKg2PgStPXVvgH2PVptXj35EhlieWG
UcfEQT5GFGwLBIzFDr92KFIyHUxTPj7L8vuQgq9iDmfC40YtRefj1DqbtHN/dUyWSRBIffAykBwa
7uSLhpWmaYY9Ml60112cjgDMqHXXEx+69W6gO9jXYcSkwweVGRvlg4ae9BROGFGdxKDXooKuDfp2
8x5VMY3+bNLRDfIMY+itO3R+VeUX6s7kmB/Y+uehVTYiBi/WiqakhpjGxBQor8Y/kAwJiF9JOnEK
0c04MP5M1lldfQqeJIjEN1+4G4HKRjZHvZktnnSHEn7AdaDRcAPPympJiLzzFqqg+lThOXICfC3X
124yxw0Eh0kJNDHa1Xbpx9tKfr7QQDcrPfqJI5xk6LnysQB9S+pNrm1i7LLsIvqjSit9fqa09aoo
KkKwyi+W9koypN2c511ljsjA0q+F6ZI3+F02YqR8ERRiU4r4bN+18eYbTZdtaQcYxBeK1+6UTHXr
dYxamSsC7a/2Y4q3psWAaOR8VtpAgYpscicxUggKXVhzriFxkTXv5J8l+GmopD1YqylO09zktP0q
BFrbjogcwkPu/brRxx9I55YuWg6VfdQ9YNxGNTrhEg616DDgzh+v4NFlNCO9u1IvGQW7cAMpuXL0
DCFI1M1/LdWp02zrBtsUavB1dKm5z3iHQ0FBmlQ2Fvw1qfq8seyRj2YgGqUVM/sHpSMHUngLZEoH
hemOhoUpoBIMm+MvHLXAe+j/fQCkMEL+/cHwSEGf32A4DTnrUJCx/OIKJmMNtHeqD2Q2P+rStsJf
TSy9pt2eK62O3qBrY92XBIR0DUUx8h9v29n5Ii/V01gmZexhh2168XYnFc5pp1WCVKP0z/LLoyu9
qxIHRwlpT3S4myPg/HS8113k/5uiy4BaX0epnKPNHBmroSrahKK/VrlRIeV2LAo4lX6lF7S30wtk
ovchu9f3vaBqhUPb4BkpAR7TVp1q6BeIFuFdTe/IxmmRQYk7dg+m4qCK3SIIa7nlzyS/FGpe9HFW
bIS5/nYEEE910G3R0fnX/p5YCKDVITNnZ6Pm+3LaCixAZTG68hbNOdPWk7+OtB5FGb0Us1FDFHr2
/jLEagkfFOPuhEEgCdybnQSdjR+QOpJPh+wkMD75jlA/FEPqc3/GFN7N7fAA1jT/loiKxTFWArmi
QkO5PNccAsUGxUWi532RdyZmdZabf98mbm1MXxV9XcZaXBU9JdU8TzvoemUPH0xv+cqFyctNkQWw
v5hmVVJnueCe5UARXC966KCevc2QKL1QVjNMRIBLybqOllnOPZvJvkTZliZCOo6hwyYkShj2ZN/3
XO8Om9qlQAfw7E8aI3VHK4nnGKFchAV6hvi9V8v0YKyr96XgEZEt+7SxZUREXWttNv6BYjotD5Hk
el/9YJx//M+1sscmWtuGyeQZoUMtQF5vyyvdohwbj+gOrf1aKCATjlLFVJKbiHukxAQMThkyISNj
50RFKX0LoziAVlEsPtkd3UONznTqf9HOhttP9QrCnKG9AEdP260V6Dj2ZiKsg5xzWrqqUfekSHms
/qIHyxyBApEdN96eSUSP7isaClXRyg4FWRnwMI8bo9Vjg+HVrIl8nybdqZ2IV4jR8U2sPc7HOL5n
CQqGuCOv4YYbOifJDuz9Pbe7msfLECHbNlYxKkFimXuW+3EcMH68Wrsl6CCtC5y/hcPpQIm5U7r3
ABgCgK2nRU+ymvNyhEUJNZWU4e8S2c8dCcAp1a1SDK2PZb06aqm6Z3vT73o6KTB3ppZNPuXrMpJW
vPnLqkA8t1C+9ygw5ClXiF+ySSuJWIP819XAWuKC1tpBtQQ7EygIBGNxsCGD+ZoLO/xHDwkdVtd7
+oHxLG0gS1q17BrjleVvPF9vXzw7oHowlN1wpsWTEtwKYQqdJBU4FnTKKhZ2qzrxIKPMfVQkM/HP
kvXBYgbB3wTwnsYGs1X3miRRQis3GQqXVFx5JUTmUnTIJO7cNDYBZGGQYqS9DDX9Y5WerfqiXm5h
ueABhA4vFsmOnbLGY5CHtBzu30wgeC4MeXvcXP3kXxmWnUeyIOpryvNi/gFBlrUWwd5O8cag8sM4
0kxPvlBFFyXiuZAcZIH4AXEGI7QsS0kjYLSt2S8k1nm5/81K0Zk4Y3MZ8zORjACMJOzVzTnhagQ3
/35cMqtVS7bXBXHjgPlnxGxyJ013OcgczsLw4yLIfYpL2pR1Yzr5JfgGtNLgqKgnbP3k41tGfcZ2
PNEtauIdqV4rMTsofYNkhFxQex762a2lTPzKc1bJHDLAu9vsTH50ASQuznG1uhooa8O6VkQIGiQZ
pTBYHdSPFf4tLHLsewzNHr4nNXxityK0RzjoSA3NGpXBLSa842YLYPwktGQ8sXnbT+ic4FxbZeN9
mjQcWmddJuYGA9GLD3/pfJ9QAFNnkSZmTC078Noh6NMTOoQp4pAxdevYsejVrVVR4czrLxDmaWYF
29s3ubS3cw1QIHhARgQvovW3QLpeP1F/fwKdjsQhLP8CINOTfYslN/L+ncOg+Qh5xCHrMUgEgt72
XQ1IqJA6QgsJhxd+cfyQxI7tSf1tYRfXVhBo3MKMAgeV1aMUEDXNEi9b1f+k6o6oyU8LuN6uebfS
KaCgC8zmYTr+5DNe2RU696zDaohwSqkP9Zm63sNIiBV7ymUOhTdZ63CWn1Mjxj1KdQ552oD88yfK
Mj/uPJibUvpHO9XG/UPR+1YvTRss64XL4FbjCwcr76K9z0PDVwkdv4QjapiAxoHHUcVE1Y1bmHOl
9gtz6Iib34tqgKVu0Byki4SUrteQ4SlbhHNYVYzHmWsTlZCGRZc6qJVjpvPsNBDLzwS5AfF9xjvT
AzIl4ENUZaCu/vfU+1x/JAKJOruiwzNu5X2+hvUpFMB2zYcDhOkFpSFEmvjKHfVT5bAljmfc64QR
kpGygxC6U2qg9snaL0fxJfnbVdBAXvq5tCl5Az4v4Pf2oTUs8FgC7aTX9ZKFU4aSaVaM6QHUQ5UG
EwjKhY26qQmk0vX9T0p1ZcOjlIqzYdUfIMrPN5OTQ5EF8vhb1Wtw7OCl5DuTFpWtbTVfvhSReLJR
B4m2INb4tVZc57/EIZ3CZrAccCZ1cg9+c4Ig7gkLiKQvR/givYs4IF/XlWcM9gBu5CK4EFy2IVNb
sg34yA1PiYxByFiVVPaAU1GuQHScqGBKdlf9MbOp84fV14J9EtFVBJfqmcPUxsM3KyOyKMWDJ1Qr
USMqvSMfpItj+6ri/iy96UitiE8W7eKBHRqPtYLTg6xDSybbDsHjDXR9QzSRpQh+f/lHfMkHTkZ9
UBJ0OcXvVsYJQ+wq1VhaHFD0xFpf72BV8dxP2dux5daKB6xB1Lsi0rcXw/rhWwU77r4umKaSnbV1
xLMu2E5tFLcIIlV/WRm48PJ/kDle6vffWAcIfpLfcVUGqV/5fhNyfwiSkaRS+vC1oj9ElFRu0V34
5g3Ywz/4vb5uEF9Avq9uuvagM+br6ipIfSVcjVsusl5FfGaPfaotvCywm6WPOFQQUqwSJKxhE84w
cnrSIPVNANukq6T34gLWxsc2tG44Yi8w5qNVvEHm+qoxyv5iJaXF+M9QtaojLNiA22lj09ZgQYkL
HXuZCOgPuMgQWQrk/Xlz+/9rOYLdo2xZY0bArBL4Uo/WMQwVNfDeIIPgqNmMWGajG52Gqs9xzWbX
Jw+ajWpB2KtAIgz/Iq7QTmmDfddWzZHkcis5iTO7STK8Qn8GGTZQRiKGMImSSRBNkEZ73gF6kyjX
PD2dwBWhz10N4l1Sp6vlhou3he5Uu5wpyR3GmNuwI57cUM6wrT1XSW9nYUxGed4I06QgOj9M8wbv
/o5DdP0+iYWQX3bqqI25EPgB+XcHx+DBMen3NrTd0LNhrycmmQQW+wjPE1sBZntDqbdbkLgfhxPr
tvqqnVqeBB9U+U5+z+RBVNUaIVLXlMQ+rOsfI5xBCoPUfRM/rsB0TclyEkGPA7BdjNLpuslC8feM
aLciNzeQlL91Fd/DQPfVAmic+W8oHqesq45ISuRV6eZo+++3PPROIgXALmSskkDfDFHLPYDLJhRV
sKH7UDqHQ0gHXA3FqblEJsBXvDSd8vF8pc5O7g383i3Qfh7RDimIrGx5rpFilFsH4y3QRH2suXQO
1G68zPzYdKkOjSf8pcYCa9EZoDqReDJnGtZqLUjqkXO0GhZkCtCtW+6Z2czbYSjnMTTqFbf5Nj7W
SR1PTDzm39ZHh2HTvVqtXMjnZvQ4i887csRsFdzgy6LkBZRUGfthORVN6FMQWZ97iMKS0GknndIz
A4xniAts0GjpVK+ShFdjyx28glnva3rn+AHP9IfojfN/QFEXAD9NRO2QIIDPalMKd6Vqvq3gVWeF
iXRKmnKnBEBkz8zxZqPoTI7T+QHGe+YAij4Bs45ts8Ygtgsj4+9tJ8a8R/L/ylNpOx5Mc/Os2eOm
XLAyCksTN+3GCIa9f7t9aGxTAD5+PuAFWEgUFzQkpArHtfjUuhqbT167VdHXi+x0cqgRpgVs0VuB
wMB+xcxBsQ32mUebMX49lIn/iFWCPjmPVrl5kOKLMX4yfEdW/5jcuPmA0dk4P7t1+5GACkjSrLRX
X+llqnuQPclhBWRuCwXo5EH1GSCTdnWDYIWgCQLgkY+7zzWruQXNzvXZDL1yDITyoTxIwwsxSEgJ
p24XwbflFMmfuM8j/OHoFLV/1hNFdC55QfmBSqDG+q0KF4Fa9+2oGVeQUDofhIHG/HDTIFLtMClq
A1+NBoiRFdhKTsJ+K6tp/CFG1wnZXXxmYJejC6HNdJyvjN9zVExUyVbw4FHB5/Dxiv/lXkgO4Lc7
UNce/HSHHjmDTjNDR2d2rXR40szxzd5xk0xQPhL8w2wPwuqOHrj+e0SZzZtImuw5kQUzf3Dg6C8J
S0vbANqVXEGIeJcZ27KMrGqpUfTDF+BkhNL9cgi0XO4Zj5M9TpFZus1FuZPAdlCzWWv4YU60uqnE
7mTP7eDccsZ3nEhnHh8ARTmSOhfLpr1XCYgbrgeJzOwpzoeWCggXdwBFQOQpK/Z6PyXEeBdh0EEk
0YtN8kq8finX6Iqixu2LhGmSwNldoCe2uQl/bJzFlfqU40yeziZZpPwu3QciNjg4I/tAwONtoim1
agtYdRB6H1c5Q/BHbqFb+qLEBMl5myEdE2+5ARzN0YYSvO0NXKYwCP4Tqcx97tUZ6B6i6YkjAas8
OcpyzIbt+yjhZSjq4hUqAyzHxkJy/EtsCQUQpXWzEKSJmPOQgtR+GtU0+nFdo81JFfye15B3MBNL
tcJtmGzKJXiIa9nz4tnkZzCqRTeA7RlffntZ8gxcDdQ+dGkr2w/G7ZJ3WsT+hi+b1+bCx128Ws58
6ZbbZu3y/j4wnXHzCInhOIuz62noBSWZEFfSkmYJYHWjE8MPH38OS03Uy/qcuPOD/Y+S1t5mcsqP
HZ6IOH3qrZ4vGy3ExDgwEs2bEl4ULEGfQjfqSartEKkYTtTC6uapV8fBKn2RcMQErRqJ2DELIuEl
xYTBWk7H61vfg6j+EawGTbDXG2KHYgEZUEgVgEJuDKw3rc4RP9dvzhNNMRgcGqPzWirCqxPvxdUe
GyRIgdHbuIAeMszW/8C9+VM9VuSCKmRYkIrDqQe7xmXw3gFF9B8hHA8RGPL7HRSPDNj5ibpfAeiR
C4fVQUgz4rV6RqNlel/pkyJw6XwJB0iSwMygKbbIrnzVaQeAy/QyZGVsQga61p7bCxNWCvg0PGHh
Bc4eKsoQWqpkk8AmnnOWtK4S7tglBFjPV8ig0NHgX7XswxjQT4yYtwbGZZu3+Beh7G0Bc/uQI0k/
6G+IwLZlktnLXCAPhZ3z5g3WAUJcjLEdHOXiGG+FbeoPU0ttBJDkTa/+qKOr0gLO2+dV9lRaGsDC
gB4k78YNIEAVACmlEA+OUq69OSD9QPalDLLZqKejH0EyQYbIMkCA4MBGigr4oQBvgtQ6Q9bYyEaF
fnX7As/pI2ERUIkpLp7C6HG1xXN15mzVwGQF0zbMt//sIomG9GWC8WIyWWDIfTa5QoFZnleq/Ic4
z3QG0tSq5Hvae6LGlV5Ck/TdtYM9GEo5f9YhGe9nznLx1E7SPdXnb1UC98p7QkZnObsWEC19a0oL
C5DDPFZCAcV+hJA0rwZO7G1XGbXlR18SWY4SrJy2njV/FER2acf2m0t5zlEC1ZCEzi4gYPlFwK8s
zb55YwkXCfJpovcauLqUOlh4cA9VFxB2SZgg2SISpKqGvIFkYDrCu5vzbCz/khJKi51zhM+onX42
5/VHv3q04wBKQ0YzENqEXtz6BzhS1PfYxuSvs/uX6vANvpZbPJM4bOLVSEVw05rMEKUopXNm5r6A
kuVfK2O/oeh4qNeuu2PXFS9omWAfkh+EyUurT6NAx/2gruAORVa5NKMAVmYhLbBLLmH41LAD+aAD
mdsHr4x6ph0/getLPxtKP0T8ke8G4ETQqgA/lUvrPZ6tt3FwvvrRxug02uzoU0+Rs6qCfBCvaMNH
xjAxQ3Z1bTYlt4HgOQhFVqbPTG7PK4Hzr/dqLhZi9MJWgXq1yeTXRyd7RhpnlReHOCDvjFFKbpy9
TzqSivYH9K3NIExnr+bLJOZ1pSpM9ByimzDbQ3BNK4gVoqelGqvepUDmREuEFmnhhInPVaFIltZu
ODVP7V7CtZeFBEt5I02fyQQRPv4RApWyfOu1hKhXEwlRFAP7wedzy7mU9QnROWYIeqjAtcpnQKic
+ULOoHenoxJh0lHTCwA4faXwOygmv70BNL/IKhw8JxMp+vxLNCuptzCahb2ql9XjH3zpElJBqRC+
R5FYxYDaNJRK6hwIApxlG+VRaWsSPpAHXl+MuJCqlUBvWXGzB5Um//Fm0ounBWLYfgTMUtcij96w
0aX/rZjiA04xkooXO48nfxZfNkIj4lZD+rTvwD714S/K8L45jvN66TJjLwL9QCwC7iuXWISsTO4+
bgyzewR1LOE3M5J5jtxvmruxarkx1dqWb92gSh8ZlKj82GPUFhgur1WYlqzl/+2EM5BeUUlyMrAO
4yICLqhrddyaPHCSAA0WeZNwHC0ZhKmbkhk92u4Vr45cF0+jr44VGiM0hVbKWrA7+3AgMyfbghWB
mKdeeoXSv+mSNAiObW+/7XmN6/lH77ad489TrxxSgjb3Dx4h34+LR1nAdN6zwhr+S4QvxL/w9as+
s0ZerwayX7daweGgmwNGkOT5+RfN79tgTXkQgekz60p8F4L40F6xwWIykbLU7/xTZHLeyIbdVucm
nbZpisgwT9/ImtEQSd6MyXX6L1t8wlchcvblhhk6zo2OVUBCVQClX08hcgkJRfeC3mGkn+fs99QH
tqV0f6WO4FTY3g4b02iDJaPBRuesViWUleIk+YczsTwWDGM3m4RQsvag80XXcVFb4KfHyQgEz4ly
4RddmRq7t4zzW9PU3hbh+HaMevWb1utFQNjwSoH0gUKLDUd7AUJ47GluVraUdZUWBGMp4Dp61gEM
DsjZUE6loiLdzKOnMywy/x6M85RZI5hAuE4dKFjbPG4/S0/1DSY5wu3rGDL6Y5kC38n9KfcSv6uy
HPa22/dNkH5zDq+PLEsbpTlOIvUDEdWOSQWhbaZTfn+RwtB8ovDLKiNlQHgwMntgPoraSE+2a9NH
0jXUPnUTZMzYerMbqlUGKUxiFDDVfnkDSibzrIwaSoHTfHmfkKESykByEGpHiy4I+XPhGaVB3VLj
AQhc/j3ZpvSw6XOv9gsDDee1zRaEYbzQr0aNtMnwOvEKSk73ttVDljKrEUBxA74wcn+glaica/FP
i/Vh0c8SrFzSDrQsqwcqIm7xJlHdSdVECoF/amfYE/Uinr6766VSZcVl9bL5sO5J5glqnZgc/OMw
A/uVPgeAGNARkEvEkqp27DzxSy0cVnFqp6xQor0iJSD1t/aA8dckyOXdBOA/u6ZYFrJ2Hbh6oTwG
IzXFfLH34E0OPbnZ27SRSCf9Vaifp1QvSabylnuwyVqLCUIRKYcuJYtXqNlE39LBO3MQpjr/y+P3
Rw/e2y+VNBu3M91BqLn66dYADEMmozbty8tFCItZ9gm6KqPOS9npCE4B6StCi0m/I2DY3TP91Gso
clfsX+VpdGGepI5kAUthk81JvUqCNODe/SFFkeQ7MPsSbOta3760BXFwRypbG015NJU6TG9AlNOM
Mi19j3ng65lM6hxJP8k/rzdizuni4XrIsdDNbxLNVdvgPwOM0J2OqErj6lGV/EJcFt3nJAaNe/TM
wvw61HoWAzCiV74aGbskoiXVSXuRVjWmD6Bz80R17YDSDPttLLcoGzI2q+QhzVj6kOCPF60ymMO/
ycnd4cgd8lX/mK6+gnfcYNqhs5q+rEDqG0sVkLdWDMiOSVI3toSIMgKRJmhMS0I5gi0rSKP7ExwX
i0CHF0yO8HhltDRz/zyAlUknQwphBebBtHTBh68Ch/Mx5MUG34OYE9NAFIiIRW1icS4/+fdEX91Q
+QA+SHciMwZVhNnloY1ZNt2TE3fNn4Nd8Npsh+588T92qm/sFfGgYTIKx4J4LT5qvjP7L1jSdUfv
bEEP/1hFHPbNGhzO8KvqiFnYvcXuGCB4jAmmzNSLC6Y4EFPkgzFz8DJ9D/BHeiYSbrOqJojj5yL5
mvIjuVTIJSxEnocGJyTcCvxMJUgWU7o3t+b13wtiCAjJf+NmQBRv+xVzR6wSP1qJMuz/wyRI+lYG
vv4+Zkud4Q0tzNjH3/1ywJ28G73p46Kyr0b48rPhCvcRkF9OZ+lCo8h70CxEG1bdC9sgyA33oB+X
F4qumxIY6QgHEj812lsgTzQIcXplAYQlVgnRF2je3bdNKkwZVSkbAroOEWtwJpdArMh5JnxDGGAn
hmv/K3WCSIzGecMJuOxB5daEAI65dxRNMyOZPEUs48wQx2LqeyUZET1FcjLfqo3/aStQo8oTI6Bo
ydpdJP1qabH8wNsCHRBhEbdskh2O7fZgYeV9/2wmXjnULPY5uuwNYSVm7pmlHfjsD8hyrkWQTwS2
iLmMicO8PnIZ07Mw/yMsT4PIXqELS0CzN6+Ayeg5VosjhNXoYOSPW9KxUn49Ib6t1k5w1WoSxgxy
MFRnIA2RBBA4RbmbvRjm7yATjuW6X+1EpMtKaIjz52HV9skxrfjYbUhRAw6USUfIp6jVL2QBCeRm
1swn9HLk59cTZW6mpMx5iNK+3WXMqcMGEIPBfGWO+uH78fdALrCfn23d6YhmcpClWCY/jAa905uy
YQVk97u3syg0qBJ1jW5Q8rIcASqmxYOsTvPtXpGY5OGAj1Ydw/+rl2P5qLf9WDorRs79O3wEJzNu
S//0soH2msqOcZglRwI3L1xU0JAoatuI/INn/ecCNHu9CHSSMdIVFU7nyFBzonLgp5v7RXPz68+I
owzipQbj0geZ7ulVxjKCAissxHJcyv6iaIYDE3zR3JpcL7NNPKCU2OePmXG5+J0NAkM1hiVlB77o
tgg+C3KWVv2g0e3C36WEODg2IhpSREH1rPcj7rRqzzHB536d94ethv/ahAOPpM1JEO7yo9xw7AZL
ml+3UXtkxcCD1+n0IEvOYTxbsqJLIHUsuqdJDWYqR+SVyjhJQ9nDyIEeckBbITjUXaStRIvGJ6VR
j20TXJBX7NWE1pmTgJyIMk0qw6bxbsn1ND4bzPdn7HqdYv+TdyOQiNmWdidK/lSL0OQxBasGfCU3
+eaAWeYrBgAXStJylIvd1V3WvKzuh5uZC2iH9gIQcFklHjS6QxRvc/+DaQa4OOtrz/lMTdIWdPqd
wC+jpqZAyFMXzoFMT6lUGKj49Eih3ZFWtVs58dW2g02g9Oh6eZS9Kivk6KFRg4H86oiONtv4357a
xOpQK1Qq2qKPfl2YOoHqbLiIcol0Xey2Oa5379m/cIkCwENndccZi84+iPCt8EY1tApAbaQMhymd
PLC9wWUBMKN9DzrYptSAFvQUuH8in6CZeshb14a9/kNqtFJF8qOx8sXH7uOnhp9OFramZ2FlAaGz
NrP6XjcbnlRUUHnoVQb/KMzRlv3B0zNfcmfcc1Fl5j+AEk9QM0xAf2HM2SQVvAlmuu4CrzU14dNo
4uDSfUwH0iTx+8gnxYi9lt7F2ftOuYvCrC5CaXLrk98l18m10skiHexSzRI3jqORegIWE0oFE6JR
JoinNmNnCTtSvhuzDo2KYGBnkcE/KQI8ERxeVMnuG4YEy50BsGIbugeiOgJNjFKAZvp3LQK3kiDr
t2jIcREBL9cwh7wM/FKDX+lSfW40ojngRhfgUBU/dhnd94Www+LgCuKdjlZZC10u2zWvUtV8roMh
4CAF5zkmGEDP+Wo4UEawzbA4I3Wdhq2G1VwHbURprfnju+vD2JIY9sbxt6Hzchu+iy7/YWPdPPc3
gWI0IdOLrnR/vTT2iK3yhulJ6Fx2qoCH8sx6BCwCOnZ+4+8BODFQPOwN9p02OGCgka5bZ8Fdn0Ca
rXus0uEHOk48JOI8Hu3MYCOAUn8pDLnnfX/0d9AoPjRv0xOTgDidZ0YNoAKj57OiF4mWrE8YHnPZ
yKqbz3IF47beGWe1LqYYfDy1Q5M1jB/YEaqe9ry8caEmz2WykHBjVKTypP5OkyToe2HRc+9nORxV
52zhbOQcT/LDsfBeAC16wPSQd+094gzcxwbkH+584PjBOAPSLMivXpfEqHceFd+5OcuHokHIFLc8
wBh7+UOaikJ3HpwHYGMPNj8Aw8fXgmE7h4SC++b8mKy1TYY+BEwMGGyvylMqwCk4yph/6IJvNKXj
l7CHd5N7+N8jpr6Cp40Az/PFAN/cusXkSZ76ALjK9EOcBg6BGcS7dEGJuvg8mZ5nHVnYfi6FnBaO
hKHxZBshxHVbXbx8jhG6G/ZAKsCLyAsp06I0dAIfA9Ps74jIJqx+77n5wnM3Fg+76EaiT2jJWUBK
cjtPkOnSM+HAoQ1LV2rLaw+lfrOALldmf1Q9Gr0xK9s07eBylRZG54rBrBWN4F00fEL7EGN8DQf9
jr1u7OAZz51UgynYhcr76fRyaiqn7xTFGQetdvDKL1mL/dHcmQu+dGzEz6z2b/sjvUjIxqxkxGSS
7v9fiL7b8Sxob1H9QQMtgIUVWXfsMED2j0tZpDvwD7A4bZFSvssLgePqzhYPZYkx0DW0vPfQ+3MP
wqhfwJgGkbgPUwe92v3kEQA4R1+X0Gqn2sswTPLkOsnh6m02hfKoj9Z7UQlWXMIYbhR1PkVe30FU
wCs3MZSR7oBnlSpxV0x3XhrdLPFzSMcVNCi+HBZyFXNj9WdS/jOgU+Dze+Pfbpxn+oISzW2MXopp
67qfo+7b/puyUyzbg9s2MbKhIC6ML/hd2Z6mBb3ABn36H0wQ2xsOHNoqzEZlGi+aYYu0D271LmCj
r1M8G4W78J+i86IdzK4kKa9flP8GBBefKwimTtcbI/yqGpRQguVnZSX0KBMwD48w0hxpx5W3ffcv
dB87n47neIKmx2OZGkohE7cYj4LUXjDBLxErE5UqAUYzmF9KGnOOFzuHqhpWLZlqC8dD9boHWKSS
AvTSdNib9kM2q//sL/YqOpVIrJElYUQUy84r1gx3hDNn1TCnvyE880RcLZ1VxK7DXNdoXSD1dUoB
dWEv/qwhWHhWieO5ue6DdCo5aGRvzZGTqqboIlafwatrU7AMtThdFe+/B4Bby6/Fve3SQrzYMHBL
9nzJSuMgilaShC1OBVF0VpoBfr4x60eYtd4vpUnXEYP2efmbT1YDtRUsKvTuZm+lZAHGxhTQohzo
SVgYr50Qx4nkqiNVnn+dqhFQ6UYx86L7Q56yuLBrcoOQ/Di8rqyXS8u7sZFRYSoe0MfrU+viIcHf
ozYlzG+RQARexLHc4qTbZ+p5gjB+VefeXny31fdONih1Ib9aYR4Zr0gy6YXThDyyNlV5WKjE0MGb
bbfDU6lFKhvNbVPL0kl2otzFdji/8Yw25m5br1UlKnHQjQ+H2DQ+A76uJ1myWTxNAN7xWWkTsULR
SezAsWuEwJayRV4QSu8yKAUOCTR1+5H/nGRCjhjpYzblIps22WM3MHkIkKTWpwS2bzC27Zb0tVNV
F5cCqzyACcpzAzPPwI+0TrQBGDwzGvWqPbtcoV7YkuSeUW0cDnDE46kszALoWnkgu0wZIiOv4duN
kPkqWcthnENqiKHOnJZIMo6pZxSDL3IEFgCLaQ+osxZs6Hnon24zKj5UX4EJL4eTUIkk4wZqfGP4
mBqpVhA4mlp9GpoTFsrzkw1IlU+BaUjLCk1MPdoAX39yMFMAL1d+Y+QE0x9b7cRkq6NUux0oS7sa
2HPTLU9sYjf0Co2kwucDpON6QmJ7I1RWuIpi20iBK2bYhimUHyioceL8eincicBxjULuuLXoPc2W
SFLvXMXyekM+eOjKcWxymwnc8FWL1zOqiSUBjDrtC2M5o14qdN1NEwhdnRWLknEJHzzTvHsuhINl
KPCtUs9Y0Ji+b4FTgdfoODLpexu7xnM0KsDYwrLR3GR5mvKNCgMaJ1JUZmOkwV9ve1kqaNUsGr7a
/YWC0bHPOKClcwh4/L9wNz34wyUv80WiE3Neb7BvQgugCOVMy8WApp/TA0+WX6Wb3QG7A6BwBDuk
5DPgDxL5Nb8+1jtMtKDIuljWlevzNyYiL1YlRWEoFCfhkyq0Xb+V9QpQikRd1pi7Zx+jCrhOh0pA
HwMBGWVjPGz8NQL6ztT3UdGZrvXJRzLA4JotAcps6okyDhiHhZ6FJRIj7vsH+UmxqFpSzXgfR75Z
NlyaXTm1NanKtjBNOzEKh3ENLPiYcoEW4ShJ5RcIEZp4wuKpeUxiIPnAegtFgjfuIMlknaATKdrv
XOavPqGj+L+RDYmSsiN1DDaMDcy5BaN8aEooRsVSi08m1HQI4U7JPjfb+Z2O/fRF7tSrSsEUWL+f
HmBd4M1yZPYZAcKFim7vjrbFvCi3E9okbJbmPfXZl2cUTU53ROEPmSf7i0yOdC3g60XMbIpEwHqw
Vc+Uj3y+cG26G6QVvlnq+esK4CYhxTvgOzaMBJHkHeL/8/mBvKLr/u11iWw1OoKoZ/Z8j1rpt2n5
nJNLxEKdnRcZEcOp91FA2VmnzktLbebpJpDApysMOppVmy8CdoHjCRu/Gwrj42LcINPmc+vJV2cB
FBOjwzxwcLlCHFDymuxZiSXCvteuSIFLULSQ2WBWXn42benJcxiQpEyG+VrohJBMsYgFp6x6Doai
AO5t+NcV1rKePt1/RMTXdAO0JZ5Ts1Vn2fSJHP+KPOP4chKo5UBe7KOxCrncj7qjnSaenIOS3Pur
GNL60NlgXDPTxLdV3JjyhXY/ZahiNyMPBWhLZoi/ukqfIDE8EpPVcQ7oIlEnVkB+EPwK+X/seL1e
pX/Y93JtCz7xvJEW6c0CIXNgHfk4jae//KIELhX6L9JUkJm7p1wdj54XySn4lzAa2ZUUcXdsoQ/U
1tobSbYPKRZcd43eWfegEFOhsOPGcbdSDJXbeW+yhmKrv25s1uNb/jjAWfySy+j5TR0NUWbbTJxu
uwJCb12r2mf0jKPBkqQN6MUhl96GWqp5cr4vn2wH+ELg1muBszW5P8T7SvSfzTztfVDKARPRK4KA
DoQ6a0GsrEedRAYdmNJHf8stVPb2vdRMbNrbu5eC1L3lO6jDRWcNdhK5peJOv3XSNbWXEZFJujoE
E2ZE7i7HKaNTAutdPVskprR0zD/ucPj0gsg/VSLqBGVbuFXIBgECbwcvpLGlcDhqEwiB3xxcJebO
h0ck5kC4d59n64eykPkMfKv8k25QijxjgzVCrlgbQNiS/whBggUWTH93zeskXiBwUoqXvOsHtWp6
MzP2A3ep/dl1qYSPZxnxT23peXEBkfHt1HbTK+l2SmHlBtLiH/tesOWnQkV29e+02p2wdKP4vwIN
pVbvEeb5+PsPDqO4LRpqaLeH9tTfDip7cS7r7v3XUFsS33Ib8IHl9yhjbm8KOD2cR2e6MLViXuTE
ag65IZe4DrHwfuvslS7Xn0PA8Ux4AL4YWXG+YTOD4yFUDQ3walDpNhm7aB+bXtDPthSPDVIyXnNz
AgoBXKq8Z+KUO6gn9v99/XEmmaT1u3vGzwcjpbaUr1Ph1ZCf8yvxVJ/XTrTGOlOEKVS5Q3cwKZRt
4WEQYgeUzkOSW/OngEeQD43jFTzBsH2XeSH9dUX9UwrJd3ZzBJj0D5O3e8M+3yGHC5wfy51wiPnx
D/3PDX9MzbnAApFtUMEhjb4EgSqe/UYch8FD1zoBe6U0J0uYI+QZK7ZFXAOcjxHh0nKOALx/PbP5
ugDaxX/X+FAUgw/RWi0H18syXk7pNMNIL3vGwJhllizBzEJjbI2yE6ANBh28Ox3wIJdpkfMaLdFx
Rt41sRz9fs3tY1pQ7qM8zICZ5iIHsp1U7iVt3qrLLpqhTF0BghMI87jMXeIyjt60jQsYrs/RPEiH
mzNWE0Sl6NeA6iCBkqKYYTAXCf3X2qq1YmJnoTF0lh28YivAKDcaHaNz+781RIp4ahYdcPz6u0Av
Mx2Wd36JOwyDFm8vLXFFLAnUatC8GSwXZPQjgHaoOQzWg0hG+49M1Vr1AA/W/IPD7irIpLbYO6I8
CRnSWzQ+3Ufwxy1jk+Z3zpsvxwahrSE3z6szUl+pesqiB4nDp2XPtfUI3RZPNYgzllZL6dhzH7JG
0dk+DAM6Rijncnn0g2+leEDPFDfyT21xvgM/jVj+ZHr2KeBzF0Am19byI3SJSTDnbeBekzRaofAF
pvNSbXGPDYOYYILHAOL+xxu4gpwJtVFl8Jp0bJxvHPrf888lHALbCJIJDQpMTBmB/c48t8YYkdnp
7Q8JNgNWwwLxyzluXkmu8xHLks2rPeXlls4PY2yF1w1bmjhcvC9QT4IKKR+bRXjfkjtlHPOlieeV
RiBgGKdGKREV0DuXbQ/OUHe9qFFCxqJ1iCftkb5jTP+KG9XexP75mtWS7O3AV8UcPEm/s9vKd2Hz
y8m7ewE5YLGxqZThxtrO8br8uWSuCkvy8TxWHngZmQ8yVBwX0l3B8NU18E1lQwy7KPhFzElDjaDp
0Oqw2taIQqIWiFvMmBiLavU5qDGrb3h8vIUuqqdvT2ZkKfSKK6L5VQB1SBUI8RAYQML0+LjB2BuP
VPUlG80fx8bBYgFX0zPQirTlRA19bRivs3H1yoqGZPUBlY7lq89xav5Ge2Cy1DQN1E7kYfqTrCqq
+uzt22f0mDhCzILMWlzbeCLSiOJby3ZYa0jqykHsbUT0YFL0pXnuNn/MPUyJMl7NpTrJ7qN+VGKy
/L9tSE0GytW7fmtclhKg8/8K0uvXFq8Q/I8dFElhElIcaSgkC/R95O3kDUFsEmhLGFisBSADOh5u
KreFrpHQwRaTwW8sRsrZGLVLfhFjqSABsiNFDBhQ11GQyhv7naeEgBib29MOuETuWMz79XFRd+En
Vqx+J6uMseo+J4kkN8M+HMTIc1eiV6fC60p7TPDGbtoglL/EIf4SQo/7/KJ1k5QU/OJDWUhiF4Ea
WH6uK+uccFpiwZJ1n2cHfTrZwEOD2tc33w0Vgm9UWtkJ46krdU84KM6Bk4/KweEuo3od94QVCZjF
1lS0R8/5QkZfmLEGYku3y+/fspJQ4FZhyKTSzJ2FuBZszAMISxga7UO4YM8MZPIh397uIJ9hcnzz
Eh8tlir2UJEsztdiQCIlhHNgqz6aFb8OWWk14dcAqNxWNjUN114Ov4jgOK9psVoDxUPygygeckQt
2f4cAACktI2jiWejpzjiUv9tzNATb4Dbaorg99Vjxrk/pLBqZMSI4cE8x8DzzOA7a5Ww+f1e8x/w
VNORE1JFrlLYXFFxixpzTaNQ9N2o2FDxubiD0V580liShkElG+aRV9xX3k+LduXbgT5pyhWlfFkh
wMdM1wS3oDPVrFCygdr2frPmcRBD1IwEhTWutk18sj1GFsIvAA8XNpgcmIvzAkdRtRQNJx8ht4Jp
eNOq7aM9Ln89XeA+b2AIEwF7dDfieFRvFY0zHOoEJVsua+kXjMxo3a3s6Z5eNk35jwux9ra6mraP
Elil/SIc9ZE5zt347XuU4LQtxBSWpf2g8V3LhGUr6kwKlG6gAZzgfL6iREJPLEdNTbSbQfwnfVmd
VfwOdu/GtTLW33cZ6rgpCYmJ2JrZKMgoYQ0o9JlOfAqPV5xYQidoTQPEmY6v2yFRKIx1ZMfr3E4C
PTHuLkaHcTpxV4rZgxhhQYd5BDSq23QhYEoHUSJJmRCPXOmRrRqG/7OJa1+VzzGkMLObQtBll59E
oWnTGE5wKGT+bNU+aQuQAVALhnW1KYMd8y+5aS6sq4EbOZDXg6x47R5jkge6IPqzdgfrpmHPpYWV
xjLNe2JIsS2DENgo2BxSaHPT5q3NDDC9ZUiLDKLkOOF3ebT3drxjFD0TOpX2DLq7CE+am3IwrHZ6
DHkkZ/tE2JoJJj1/M19jkunmQy4jLGUr5cf1HCbJILxNwb5jHechuYXJYfdIpc9wyyKD9+AcRX4M
U5+dZ0Pgm7BIux+U3+7AWu6l0qEdgjg2PZ4WbsZZPczGcl+rgTjELGY4NktVzwVTxZOmE8gDZNcS
tHiKtUMq5V/JeFdILXE0STdk1owIf44MFqerI+iavdVd7FeKHqXDaYB2x042tAIpV5jSsWdLU6C5
DbHVNZCtTOwk4lNsctD1vkGx9bDthxexIX2tc2NZfqMN9fW7Vo/m611ns0ki+iqgsabIC9brPHpW
EuMA/UoJWh1t87Mk+ekUo6Yk6U7/UL/eJjWql5E8ozL3rB1oyyvGjcfSEEQTR58N6Obh7+ZEQvI1
wc/KDs8OBPPR2ub44f5KAA1iiclzDISr1Q6TNDe9fcKGevZdS/P1DfSAXR1ixNncDn3BxX13Gwiv
jLPMjZG5Y0IhHd3FSRxXNF78tfg0cDpap2d8Ot5rgAlsz11ldKv3rIr/FsVma8EshQ8lWqE1ZX5c
FV1JrFOinW9OiaOYfTtOBs8hYugsSZiSIeFV4/uD/Ez3r0/mkmZ5ZurSdx1Cuy4ZFdGdhi41Xvod
A2XQJDDT6z1SgFHf1yl3w8OZbzrardpphO7A2rdQcmV08VN4AmzFaxsRP3kr7wyobQHoiSlDsZu0
dCVfTfehpFbe7VEbY/nS1LwWFsJIkHutdmOBAoPV38sQcCaD1SJsggdS3ovgb1E0Wn7W7qbwcnB2
WIjYc/JUD8Qz6IVcdo0r+vWG0wdpBxidia4YrBx7dpe/F04ZXj3l6jKYOpOSKlbTZdp/WCY6Ge3R
VxIJlZUeiLTG/0ckjOaw+kxTit6ZtKOx9qpUD9TIgja77k9oJvL56e8fpQvfjf3irY8Z8SUiPXpT
t51EL/6Vl3GAoxHX//LCBK7LBgDTzd+MrotO1FYtFLq7NtZUHHfgW3/n56vZhosWf2cljrAAhaka
f63gpj8XjcS91g2vgLw8teVST+AMtgrE9hFAuDFmCxXw7JuHFLEixSLWcRBZGj7a+ZIgq9m9jOAc
cd/UDl1t6SHYtxQPIsshdzmCOKdMYLsdOIfNtmsLZH4T/pPAeqd5IXdXlLTq9C+gMDAIC2cOiEff
ZrMwydq2yhmojvstRYyB6Lx9nYuM+YTm4wdYG/UUgQrJAs/vkJtSO2KKAxguVd/oKggVjx2JuSpk
fet59MDwhassK6jmNqKZyGV0ioGGNydmdk5wGsHa9y2BSGMK3SRmb4jTl6L/9qOJUIdodPKd0lC4
dK8qMCYDxsFi4FBSZEhHEziLnrDmA9oWRYEbl3Yrb0qBigbzpUaQ0aWvNPnQxIprXgOKASrcPLti
FR9dNns3CN43k9U38aGDiBAyUaiOni5PCgtG8zHAeA3TC6AIdD+YVRqWjqdR9c+gjC04bQPdkIdV
vLRf1r24gX0TC9x1XSVo32dEFXC4E5Km+reW0eRZSvgHeGoRoOlWhMQNPhP5kV/BX1PI5RK0EYBp
ElEPLQflhE48nDO9PRdah31Liab7KLV/Xa3QQyy2danVtsLlwBBnJB8qJxUn7kz4m1xQ7WG32C4s
BF2a3wBXdBCY7xRSUhBqRaDmMtWzfkEBLRXUvBBEYhlNtgHtclG7E53eK1AyKZgZb6/ae05BAHtb
EkRdyiM1L/qgY4fwpSDl9rgIlsoTzqWFACrqgsRkFkTph1GN9tyc7+wpDh+m6sE1HlFONgMw6elF
ht67JRYUsef1+lzisDA1cO2k1awDGy+CYFRhCwWAJL2a7QXlse9qqk4NJMKdH7880/XbWodA9E3r
IIAa2M1TiOuJBZN2ghROAqzs6TXRK2rw2Kvp3d/0eX67S9vB5pl+3aFHPDU3CM8bGV/hCW2NMK4X
fZfuVqtdg47orQsKgkZtwqRPxCzR9glgvGpEu3v9KQXCymDM1be+k7xDbPQwwfdjsTIJI+d0pR+z
BOi2tT6s653SWSRuzx3ahGRhisyhsClSqWgPI4OkMLX1kNYtLQnLLI1SoyifA3RB8mHIo5HLyDKv
C5bqY/d9aFMQTL6pa8ptweJJowncQ4Zx65Gyu9b5t7eZchygrqq6wPrz867WE5ScIOZ6NYQQ2oOO
yYnUbJdFVOU6zomTBlgmFLh4UgDwvq52WyCwczTQlLFuKKwQv7b1oXu777l2rMHhCGJt1Ah9MzRG
VimnsT8VcT8qwsGgtV9SBl3ekMQVD9qmtZgYEwineO5qSyQLD8S+XU9ArH9KnvHDH6QUK/d//w3Q
hKuSSYaSkc5DcQAhWtPB3QP7ARvgJsN5kpK4dydmtJUeQ+QQcJ3cOnuBkqlhq24AWU0ijjdqX5aQ
yYKoAf/5fsLIG+Yf3AHkJCrx6If3YdJHtZh0qv2efw4yef4mYtJ7hOWfS5okbSDS0cU+ndsCFwsm
vpjAUNSENDYqEbpjxXpq27ELhGxVcsKNp4Pqb26f9oL2ELHKd+hSTqQjVX7Swb/uTXJP5ISh1jlb
9ErdprEtxPwaHX0iDalMCMCPFfLL5/MAOj1eqkwiY3mQlWICxKKpJD0dDR/OaeF3UjXjDGpSB5ea
oKsxWDyUaDoRWckZlo/Cchex9FxrZBz6mWkq4WzBXUKXk6kHuz0IWeVNTZMtIiXKIV+RavVUXDxe
ohDRynjaLgQ7ALNwEmPAFf1e+LPSLN8GX5nrHpufbDE8v1WQjnGif5CEvSwRwna+0RX9R/cZ1+pz
2AAXlVG7quut36EhpJgj6+bfObdbW1QMYsOR8aaG67XJXWhE9MDgZSLq7wkEy6aJcgWiAjmBhl+1
PmVcTdAYZrAMxf0JhE2NWcsfmzM2/vyjywtwqT/uY7OLnTvftZS/5c08BJFPukpCv6YcbE7WhhXY
qLfHvKRyGxjDGAXILhFPKhmsRYcjVDM5/NgKVMLx7/pxpNY83iZhBSOtWV+j7n6j1GEJruoAxgff
0VWtO4WYI21vhHTNoTLtDHp77DTyUJ67YiJgmWb17PuU0ghRVScyic33u7eNpg4T1DIJCXrv9NII
u5fZioMH7JPTAMtlaNCjpb6LR1FxvXnQR8iing4jbCNpLiOCagwL+FgbnIfJhD/i2ekASPFDTxHv
wY3d4MxlbSZTwcj0LEd3LQZNRUDqBOO7Wn58j62WZUJJGkj1UdZBmCD0/aCirhQzjIFPceCyBSDC
El7XkCE/hw5tdW275Sg79nOG546Zl1hpDNZMC5o1OXX/JOz2BI5Y6f+eANhR5fCVVCEDa+rf3eoL
/YFvMRawHtyzg9IidVLh5vZBY52Z3m3QRGZOO+p9VoQUlaOVBGezPuVaQfnLHm/wvqUQ1z/SgXpy
kxZkeg9M2T7A2BxB6IUDDE21V8RFuxpJdACLXjwqQijSNdvR3cFTq2DO2x63dgEPMokT+IsEv4FP
q43d+7lNIrPN2y1EOAbHZQKk6JEAHT2/r1UNHwBa0WKxEOiNhgmQvnGJZDbs8rd64uaXio68X5yS
4DKZLlcuy53LREQ1IYIdJ3revB65XGFKGwvT6t13smXPSKJpzNNUNeLYZzDi1K+AMjsgU0yIDtOI
CqBmIGhrkJTTMthmYhqxqHXKrmhHXoNw/OXRJEn/IlxxIan/cflG490xDqMe4nKRT3h53idjrncK
AlBquEwot4HReU//w33O/oTtNFWk4D9OIte9xUzbFV7g/ZLNeZ1v8OIg2VahNdMvwYT2Cdxx6SDv
pNHDSp/hbAJHLivgdklYLNwb4uZCqe23TF8GmIThxThS8g/4yAgthOnt8ebf8xwLvo+FOGCd+Rsl
Y5ejNvNVK2W6IjZQEab1M+umagJxsMaAFHs5n3Vwlre9H20rAL3xcZgKGfS1IluySqEHJ99mOlIx
xc4oMkO5s9Tybpq6JU5MzoreWZoacZbLhKpbKrn7HMJHlEjDuGmXb0WJBmLpOK3t1h4AQ88M9Fy8
YoKFXWDKLsZXD1/rvriFk47IkykngV7XD5gOG56TCtddF8Ab1Wiu7l4nGeDKm3/+JlTi8jttOCDA
3BvtPsMFHBFt++6fkz/x4gzdQXIZW49VdL5oYclTdFD159+J/2X9iUaYTUkNN2MtFisZz5YLFGNF
xq8n4+y/E7OeQOB+3AK9wwDklOe2eVnmmcA8ae6ASQr4a1DO+TkCzmcD9s/+fHuyqHYIbKIFGilB
7USDkgfqdPnpJ+ZV/17UCv7JAYlrevbft5uckXMGeixMywOQS3Xfy95TufaGkCPKP8RQYi5cDQVM
O6a1RWJ4aankoQwIeWPq+xQ94f7ulJLKLS3GPf140zTgswwdBeHj47+FCOamvrFFemHX0VJ0KJ+O
u3N49jsHEI9cuclbVvCx7JUedOgVv9Zc2TFn4LkIcJ/qcp3abr3Ws881t2xsE25MFg3GB8trub+u
VZrgdF7dWQ==
`protect end_protected
