`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
c4yY4Ds/ih80H8ktO4iwEXZ0p45iFFfJQDh/vhCoP7scl3iebmuZ4f8SbRIKJldlNRp4/zYMURt2
czPF03tDLqURfpMHoQfLfhBCgwI1nQt8YMqMTUptrZz+UeoSuHwAS/+5vVIyvoWtMuD38blTgOhS
mcbfkdC6G5sbSq26vmtKP2K9hOUa+DOjnWbYHjUWRZTF/jK4cKM02y3fRYJsVYig/Kkx/mXcjgE8
BIwablZV0XK5gEft8fg1d8aV68W6a39vNn5sYe40BLrztweYQBiwW9Br37WL4QZzTMN54Ptr1G2B
Xu1JKOFgfv44h1tZjoii0Pza+zKYb0/5+nGvog==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Cc2wXRaxGIcvv03oC7spxwtdENfwKd/asT2rhpOyI/4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15712)
`protect data_block
dmXEAn1Bxk5gkwy28NApf6ZWl6WNx8Cvl12yEj79RHJFQHI9SViDTS8enTKtNSIF6zQwVADff7X9
0jzhrr65zJdAFKhD5TK6RvsblNK1t1zbqyx7AUuJFRiHSWVE7a/kNh9hBM3FvhS9gz8/Iejo8L8Y
odlDOona+RFnBIgoTjuS5TSz8G/riSC2P8zdkvvdWUh+C6VyfQ/6LTYPTbpE4Hmq5pNQF4IKh+tz
if9BtPWgjCqYiZ0eG3EGKIzyr1r/UpFlImrvlnAOp7AZM5DLYQmRJYvlopKzDlBB3s//43lL6eOp
L7d8Zib/UjK6TwKynua5JSY71w115bKx/64oR7x6OHXPY41s/yQvHRZD2QjPTR9Ya0Ju0mQZlsDQ
ffkKnabOXpbDz5z9evVmWwKBMkbLIKTttdtAIJ0yobqjRJJ1Wc0Z5WMQKHFrJlf7ORthC3j+S03e
+ljA+5eEuhUlONcz/zjUZbkwLBpR7fPnxnVR6IvNefuYneiHjmiauYyxoeVKl3J+aVi3kXKq4AMA
SC2jXdfgmen0R2MYKLT+dba9GKkpNpmPg6J/1xQ3FdQaokjDThGbuwMxHSlugDx34EsQdDn8F4mn
8q67At389r6M30qXUcOOfnFg0KzAJ81Ri48EACElnbaPQaOoH+w/ZJPBWHr2W5X4/+uCDAAhErZB
obgPeoqZO5F0h5+qxPSSIieefZJrgsNQH8RMqqsgiBEornx1XyjjHMY6k0Xlr/N15gqbnSnNGvpF
ZM4m7rfQRjEaQ+8pmcLT6ZfKWr6pIdT4PwJ13QAsG2RrXLn+7CAZKglPustk+J8XvECDRcnCKH4T
88BjImwN43PhhDZ7seW0bkya58ThELG9L/1MHdiJ6e+OtNQpgNnsaWRnWBvu2oCu2ZL3+d1DwBRG
BrsKpjzNnDJ4TF5WleEochYl7B+dFhSUKCL//5G0Ya/bObnCSXyA+oeJFgf5/OVE2LzDezInrGxx
b4OSOVaftzAiYZJ3D/ejaK8i62cfyh4/ZhrpflMEJ+sXJ4Lhaq3SEVJGjJfy+u1rWSYZ/7pooKjR
1oxkyqRhvoGB2J9BVkyoh5A0mCjXnVwDYViJ+jFq1cXsENMeudq51Yst+cCBFgP8oHGX0aiGvu/s
sfXjjBMJ26W8iIGyTb1N7/OD5puJZOQXfCklWQYikTsTaW1LNa0lY1fBQTK7d7lpj8EUGnCx30Q0
CElYY1ahkKdV/UnNi+cCHTVqdNSN5eWKsw0EzQ2UaHsL8VULtL5JqHtpIPe2DZWZ4Cq5ORPaP0xq
NIL/ScSfgjNVybSFj85OlYLs2mGFKCVmAYN4L1ruw6OyP/7/08oDmLBOPVBNo0slWrdx7bWUnqqJ
/dVVBo+8peGcMDUhjAG+54UV1rMvBL3eEoRXUqlkDxdUbmv6VDGjkkjj3fGHx7e6QT6auoIR2Pti
LZqvUkP8na5PPYJxtTqaPB/9IBkE9kW2uMDOkRXKUlpvzcbRNIqFddYqw5NxvZcqGnF7GpVAskc8
4ceIFKrNWbVo5rqnBgR1G/axBzoPxc2vx/8sy4C7bx0t0pNx1ahMUTAOGGsuPUHcYRp15PL+aBso
HzlaM9+sfBXwk7nQ8z0Uubj9h22HhCKQMHHNj4D4EY+obvWuLbWYVJ/Oj14pgNtO21Kff/B29TRL
e5jQiC/baoWHWnie8VR3xVX9QzwB9pjUvt92FFgOD4lqQqaj376kEFqTj4ZVG34ksHKDRNmpxbLD
4mjCcSXDjimpsuKrXa4N3pIdiIUWsDCVVWYYckbbZhGvlYkIlSvqQS7QAp/9w6juyA8zQ9ZSyHn2
txj/w+ruNval11axeeMPhXl/BMEObSGbtf6RrDVI5dLGYVTrF6DtaTEUed9zsz2jKz+XMdPX3i7N
L77c8Zru23taI27SBSS1iQLN5paJRvTA4VYpM2ohKlvEYI2N+yrsJwoK3HcZ2LzQDYbM5HxecVjR
eBm7MDOyaiiUvTq8ehpOYLGzhrO9v59gbtymCp9fcCsnrHMeFFeHV2MsRfYWuE3xwBhHLc0lksRu
x6H/M7LU8fwG+/I7rljTGXlmHBOKP+EEsT7IV9LwIhbFXXdCchyWMAgaZ0256Sk8WD9wyfxN3jGh
pyjSctYPUFHVQ4VEk/F63GSdUXczk5NBPaz2CWXYhlwG6XSYeTnlQnhMMcRyMjR3VSaeRF3Z7ZIx
BBRGtIDOqfmT9A3OvCfzNdxIt4ClznDQ64nE/ctd9PU12+eJ+h4dc6zbHOe22ym6pN3c9P1dIsdC
vXN7E43berr5F7H6snL+2PooE217yiFvKVLGv3c0GG74hjR6jcSYg2a7nw0204h0hKd/hYiqxYkr
qSL6OpZlmYsZRkmLWyVbyzNlxw435ydSTNRZZG8p9Lh0EIdJslfGzSUOSuXymLt4HIV9mTSFL2rF
aZ3L+Fpvx7upBrMRfajcVKIMqXxtACKVOpf2w1Qpt6xmEqT2vF5I7bKgcdW91QSy3S0ZQtZDlWuS
mGpsAWYrMLwmY5WCMxsEw7VdLKtP5os64pvPRamdmU1dyFC4wa0gDmNYew9OrT+eFADHQAuJ+D5P
gURu97QaeMoiwqva8msGwQZ4c2Fy6csG8VTCz8SA3F0/3rRjNuAs+5/ilNXIGXOV9xyza+6sqnH/
Rz4n8b/eHEMnEbayjUEzBxnvfYGkoPL+gw3kQQiTNrNCs9vDWsSwgxOYe8Lq/hqQLK/8hBiovPal
caQhZ82ixF0u3+473xJhe5F9/qSV1vyIBV3caIecUH1aLAwUfu3F7+NhQpWuT8gEvmOo+soCKQCT
egY7F/OHfUygNzFfTy/ihn/MrAsuwN5T0eb90N+/8lHY2SeifG8O5eO3N5BxFVf9pyyvnon8G9Wl
lPvRuDWI3f7uCw6GyU4IhfCWmpW16MSyVRx2qLtalbTU+S34dk+F5YPfAOfTOzXr1ljnfwuIU98U
sbedohO6ygxrqF8Cm5V+e3TzIBtSaDgVjbDoO3LAEjSfHvey+d5AHyHNPfW80Qsag3BfA3Q/xzye
FDc/JqSmyU0cz63EcdiWvJW5dvR1C4Rg1PxikpEnFNUn6+YAbi7bB+h6ILdZMoGQqINGJukqsHJY
OEA7PcoN/jV99dUXJmscPZPG2rar2ZImYFafErKJIc4Qu636LoSqbLTNC8Y+qBdOcshj6crArd40
lg+seiiX14ii7x3KwqyihW6IWe0c/5wJn83r23Y6BPqr4DarFH4/6p8Cx2QRHd6qpud3RlS025we
YL0YTihv/nw3HN4taKrwWIwZSWBuVpmyOtNteZ2GQLax4y5iOLHrz17KX+J4/i4VFox8+YBFwM34
obaKadJY1X25eiSXN7cf15SeIlv0dx5AaKHQL5di1SpFU2aMtltbbEEuYl4z5IZV7pLVK3Q4bODE
8hQT0X7qIOWsv88EPVhAOiLHZtlAo4I+1zfxdW5/vXiiSb1i3lDVtjp6JhA4IJCK2P/369So4Dkr
D/grcG0v3SWVc8eMruAlRkLbp/sNG8Pwbgi2Ik+FMa9cz2fGWtruBQiTrl+nmrdzonDtiun/2BCR
mE8+PrPfrPdyRzV85nJcbutMZCYg+aVqQQSbzo0pi7RA8EbfYk0IC6tGes8KfYWppqbT8cixZINI
FwozKM5H05k9CrMsZlgiUisyCDZszgOHpzBDffs17Xhwd6tOLTv2kJ1p08YmcmDwBfAp1Htn/uRj
BT78vHvaaOLsMWjckwrHXFvFLENo6+bGmPWDdJgNosPAHh4JGBHkVLR9uUNxPlF3GUBEt4JW3OTS
rqIoXwgMoRfuQ4yfMvfJwtzHoKRPMlT4+30+ukw4EtaxyqV40kDeO1tBvjjazSM14K/hPDYXJyk4
iDQNEy+OjPte8kYYw9vztUPcR1Kwcy44/1z9BYbrHFNTanXFBeIhczUa035rOXHm7mTSWIyG9Q4T
7K3Hv9TTHP0AS1RKG2P2dXmCCq1Mm/x24m/dcIjI+4WpOkhWHku6um2SNohFx/lGAffnPGSvytGC
MNzALdF/osljfOV1B97RpIplIQDJQr7aHQsqJz5Ve+1g2l9b274l+3/tc7+cFxfZcDBdSf3jFT2M
KvgYtqsdx3MsV75JzA+/My61w5CbVU2LF+r4Is1wpqT/A2ZK8asXfDXhrW0Rb+mBRMHuCUlSycd2
ponSR8H0G8sooL4QX6cNEqqEiFq+IGHDUPFn8YxybIHCRyldb8BsrGKzGGA66cZ02aBDKewwN43A
Ft9Tp1y4Z73CcZfAq+5hQ7hVYDaJ4s0GqsJLLfS3HCsKwxJHla0zkaXBjkXLP2fYsSkkffrsrsjA
3nRdjYUkvqEUiltnkTbDCFVXD6vzv9s1CfOKZKiYh8dxSYG4ds+16AAeS+sgLn4uAigZTwY3TeP6
6/QJbh14gKLM746XmRPm6DoCv4nE9mvf4TQKTOFRgordS3K+oGC6FUokXVTNHDX7rmXU3e2RYKh/
R2AgnKxMD/H3Ay7oaKPFade+l1N8dWvXS+rT/GvaDplW/hoM7UgGklV/e1fN/8T+Uy06FU++kftF
aKe9xuak7FB6h3Ylj587Z9m8CxyfElBNxoLbrTGpfwpXbZpKyGwSdhaVIxMrq0yapz9dXDMGjx4z
lh6mpnSl2e65jJATf/Rx+GapEaV+4TUxXbIaOckOC4lLW5moQVmPK2Fjjl3Bw5+flGFk3Sg+INoG
y6Hw3JG0Cc/MdgeTq7RBFYPprzu0MkBom6NfXYce49M/QetKTG4aS31KgTJs4Vhw4/mJsXrYL0x2
eDUCpdMkX9C8x/i98zFgaSRbWcKKI/mo+lJI7fnkKvD7kOXqCpnHxO46rG0X5TOMV9RfrFIEIDZD
JnY2OBhMz7FpuwoVYuZKK43Cg+1knymSdnJ25eemlr5hfzSVsE443104io3m0P5/YLOvHomhTY0D
mXVS4yL+eXAqCocoEVrBYdIlJc/NjIqDJpLxK8kVKNBjoYR1kT0ml+LKWw6gQ/jTwNHTuyAzN2Rx
p78RggnuwHzrn44STxaPl06f62f+FdI7S/QyLijL3wqgrK6nw8zWT1Kc3l12FHwKLI5h/qTqscFE
b12tGbEsGb+s8PQ+6J3XqFWeWpGtSVl0cq6Q9sQr5ZHoY2xBE2RS2CVkRvnHH0/y7pZ38za5jWbj
e7AZ6ij0raPv7TsjFymt3UkGyfnHGy6YK+lhVoCuaA4QzNKzLqV8pUL2XxVFtCyMVsNAYc9EnrXB
D4GqRZlS/dWAp0MgJCbUVhNd6/smBc/GTN/4BtyPiYAsnknfEokD3jUK0E0k3pW4chVn23+ywegI
aDO1Ze3W0iNnP+BV1nVya+hv/J53zlDrktE6vRe1iNuzir3H0rIiltLDCPYm7Nr5mTawo0Abhyy0
NfqLGJCwWbAbUYxp1+xwFw6lNXQHYyR+hqwgTWC/xF27Nmf9ujdTfpFsviHfIjudF4OIlw0U1Rn3
nNP938FECihp4OWB9e2MeQQmZ57fvosgUvaB8EK+XY7UYp3Jnnsu5PoNuFb8xUC9pL2M+xp+7mkV
RmjgIBXsxk+BJVDTEczmY6ojUpZZGhcL/clkjT8nJGP/KqUJpY+FF4fMt7LnzBBchsK8IN4xIF73
G7p4gWg8pOlBPcAd7qJd1vViYIkxv/5n5aRbYRTvQCNFkc1oKthIck24RNCdKdGICABTxDxIOequ
oNLuDmPHsLDH84DENBa4sIuERxE710SEt55ZggghdMFPoDpkYYCr+G8rH2Jb684WNDqfninNJ3rY
jYR8Q7BKPsQHPVMP+Og0OmhWEuWLXizgeAYVNqM0/q7yzA8Yx4KEQ+j1e88/QTNwRb/H/xDVhPLS
OYUii+3VsuJeCQly7M6vRYEnG80Y/BxN+9/SJK/C2kMb+BXK+WlJkhLilA18WfptvujVYzmpH+84
Tbsu4QI7bMBKgiU5GN74mvAxp7lwXQWItN0oE3wFYyD7l8+5oyMsspuk6k2qWkGWIUWM2Ykxh1UV
cy5lCzEn3OLB77WPQl0+Z2vQwUPtyfTRm7sCujFChRYjW9YJLcYNb42kDat+TXFb00fR8FW00r5V
i7cbEEbEHPZY3jeF6wHuiHO65EI3r+2Z8nfvjHqyKIUxLCZBPhb3X1pfFD/X/BPXoAfzOHpZwIKN
AYAqVuz1Rtg8AzBcKpDLh3NE89rOX/KPdImiqDelCak5+UN4gQpbUIWsUWrgcD/fbUPki6822I0F
ptmX9aTuqkBf8LJCSPtopzqF33Qr61FgzuAF3KD2Kd4xbuijHk6yDW35EL+HqQ8rmvLCdAEIaWp8
6vqkVBMLx4IxPSf3tRsdd66Syrs3tpBAvmgeNbmvnzCXV5Gb5IamsHbXOCx67V2dGBUA5c0U68yA
LyymGM5n6DrdKkZxGX4fxYqD2gbSyH5fXIsG81rRXF2APxCFvM5zOos3gLN5EqIy36U59gopMqWR
A9Pvh3kDcERKVxRCAMEPrrPcLoEzabr9GSe4QszF+dhBoITupNSfh3FXaxn8QEoagXCvGhZ9u/TL
/EXTJEOaBP5fQLMVJUN8XcS7n/PZ84AObj1e2epHVYhWnYP1ILjZM3mL1i36d5rbil+EBVzKgEXS
Gjdj02PMLN8mOd/cA1mXcLYtuDtuSMO1Jd74Z8Pu1xiOcN2OxSAC43RcDL0ji9ZzRNLmUQRUU3Uf
BAH0x1jLcgtAs21b850kuiZTBacem//pbMBkQ4IwH4QgbcViW7JrENcLwiPV57Lrj0+ufu6X2w/n
z5vxrr9LK06pcTj5u28tVP/bDT1JJj+fi6QU7Abml2XzgHUYcwAuibq3mYu9fgfnkE1z+3eECHGB
Siz86tupClFim6wtu2ne3n+fpf/OcvMSZBJWKl9uRd3L6qUlJI0SrAnJyNuP+S4nPy2te8TO9Liw
S0VUPsMkoDCyWuow19j7osU3aU4kmlVsbrrefyWv8Gl9oTUSc/fBoy5Ob+c7Fg0WIQOBnjcikrFo
rR63Zfoo4nhfg9bcEwBZs0Y1a6DDuZrZVL9XM5dy5Zs7nT98HqqqpX6KluPC9OnUcScBUDDtBUFj
ngrZ1uTNSVJ67IXqgQLRC0jY87IA04f7EZ8AdZHamUhq7+SuRY+qLgKxZpFMPkJiUIuXsZBwF7T5
usZYz81J2vZeABQnbP5ueG762zLI24ISky6jZymC93Hn9o/PlyLlcn8m6QNeB5ALAC9Cnj56RhME
Jmx/47ZN5BMbP+62cm3qMKirns+iBfazNjx6s60SLwnLcXSbEFrlY5uOypUkwFSCEXk42U2xiCve
VkhVikXHTHs9zyndwCFj+zmTBIiNjugrGnp1Tip3R3MlwogCgPqwEuIq+dG1VHLNSIYXfrMejj9x
wy8ayaxIUKzGf8rimxqZLYpLFTzmcTWBU04BafiHCN+3bhAKS1lP5KdlS+ewqxLb8+lbMiBjaewI
2fZHp/IbqNEi65KaY14ZgX6Sv5B3YwdXM934l7XMd2MkReO4UFGohiCK7wT3SM4dou58D+Q/aWBD
c0GUcXzzdLoaxhQU07bq+tffXNDAM/xpSIl/ySjGJz48BBw81LI2e2dyc/zQsLvy3K4sDJxuLayj
VfxraWw6zy7kH7HLlLFC1V0oIT6ND54zHN3RiZS0Fj/1m6sffvym5QDB61+hNC5NgtXtp5uZfK74
MOycjXdvKZy5mR5hTCxkkdrUXamOpmvvU2W3ypwQLjRQp/BKxSOKTI12+nZ5tSYTGOMYvdCJ5IXy
cbFDBqzzjuWrA04lYDUVXd8JLEpIBDP4dwDRTev71WBM/KoXZNBdXMTG8KQiXD97MveY4tC6pWFV
vpg6+pA9prc/lK0tzHAdw3Cy7sNR6XpTdeJ5sa1hoW2W3gy1Kl72tlRHJN81WhPGx2BQq7i07ZR/
cme45T5JdFby/mUK07Z/9cyzvr56LwHFfcLLpjoM24B8aCo7/XEoY3I9V994hl3GJa/E1Y7+mqDM
GDa6OHYoL23Jfx4AuT/8nst8W6jHob2T4ztgce0//G7jvx4tWKttj0lseX1nYqZZLAFAf2PLBqNF
24DWsinwKspaqvIEvWgHS4VvpmGfYh3wjyQvR2oyV/QY3Eoxf3xvR4CHxvtv0jPHMTOa3/q+Aglb
GNIqZhfYOy1eqvc4L9leOUDSZszi52NtqWZYQ49om5pWl72bTdjZ38eX1zpB6RmOTYnhWMRV+XVs
s18TSUkvF0aDHJ4/r0xXkapzM0o128ckhXJr5CWOKTfQj93NcmXXvEfxoX8QFI0eR5qi+VTOn8wB
o9FXeULGB74bZm4ltU4x3R7a9GzSg5ubrjPKg5b7V0y1W35+z9fXIF9fpi3xKoxtEoqFBRYaQcec
r32qLhvZ3Lq5zumwInzoasXMDt7Zzq4/aSFgCv21rl8icoFtOFIlKdlrA0L4wYzXAHvfGaUjpaHx
sSuYs719hwHBjS4zCjCYTgp+F8O8gAd0AtedPubrNq6QQTWY5PLxzC+Aw61LaksgwC4ajLQw2uO9
dLL9jAXfgo+10KhGmvmt78ytMgcX9ce3Q8sSQS3n4+PrdVZ9GJ4pD0glsrtqsb3IPMM3nxuFCx7B
ecK4Rg/hKH7uq+/chmMiXj1SLDMOTRBkTFZmnaa4FE28oqAvuGHa25gBpKFQcGazdkDWvlQptBBW
lxN8YLO/ysx7hhzpTUdczs4rY/VlkzPAMKYGVBzvs+6C3H7JwTEyh9pYMYVccxFYIWE55c6vUOpQ
6zbCLcTcGNWliGcgLHpvUAf5p388S2LJqr8losFSuMuvYsLTCYbn1cqUNQ4xyCq6lSzU5LxndHK3
RURQpDbaCCjXF0SCAh5QwvBdCHPAAxOGOZMVzciy42iAa4CyO1ohwErYIjL9pBRnZEo7D/eXL6NJ
wmr7A2BNBHpM5NpHyHwVPz64sAKZIZMcbNHkxDMNAuRCJrQidCiZGrAtQqqsZk7vokDe7yejsXxe
H1amK4CVnDJIPsGkpmEIoNiuvV2wRcsmrhokom8dZg3QZ6GQ6EX8In40b9zOFWaSfw8XNHSuzdu3
StoEcMBEElFzMZG8PkKJfUVHlRx03mpDagvQAcwewxEFpwkcnmWTrPHRG0z5YB6JzL4DNv0cqjbO
DacdVvNDCW4WKNgBV2aLAFCJNvfdB807BkzSvDLqfDuBphLf7kF0zVNIVi8JwkBQH6nh1Q4oOZvp
K+pgjZ2YnNbl2GHUraQUQTMOwUWMloa8S683QNhvdzeUUPByjtVCnXYOoiQxen/IgNYZBafsbH0L
NqOFbU8rNad32iN/IVIbNC9xSypjf+0qpQRBr3T35C52I6P3w0d+Mmdffui+pI3hWF3nSPuyvS5v
UsVgA4xB8j2TMKRaYWHMGzokCes2xk9hN+wx9QFbAKhu/y1+zPoVFHtFIICiAIYJcpEybo4xJSDU
kKYGsMW6qkIsesSvqX5Wu5/geydFOHMmKSHZU9thrk4t738V5H4BbdeGE2XA5x+U/L+/cLBwp22r
oU6qPKKwR3YYBagpb62K17R6TY8GsRae2Lf7Ue71eqnqWlWJtGjGmJF0bt7buveUZhpc74Y1gt3y
1Rqkr5ZBVQ69TZ6hJAn9YWcD9/23ocaVdSkew/g0TjLVZdJPAhfjgXAm2cRPdwSOQl7tSTkzYhW4
3sCjtOw/jzagI/mUfLE19pCnQI0F6Tm3+KDfAz8EKhkjIPYegAm4qdxvrcaT2d3k0U1rru7J2fIe
9rLVKRRgzFy3di+iCPyp+zXj+F/sWf7BuXZZH+/sgNyb9LZPPJbJTfhbwB4BsatWRZTwg+zkZ5Qb
C02ePVHx+6H6nXFfTKFS/no65dVJ/EiasLOKQAuVNG4E1hGDkfxHMVfE6JwnLYPHLyTBwCz/JixL
1Pz1taVEKogCDKSRgjTSGvczJGqGSD0Loxc5xEykfPCQaF9kWykqLmP9aQOGKYmi5FYPc0SXE1ol
71UX8ES+5LKda0hRs5UKzfaChz13/JXv5WoyUf+e3GeLK526K38MiRqki3LmxEN1/OxrF6uXDaZM
sK59Zm6U+Q3Kolh8jtPiKnuTj5zg9YjbK/i8IfZQI+wXsbD7iNGzFxc8cM49hY4z5Rno6fFh06qP
K+OihDTx6aTma1VOq/Bl5IxY8CiIt63cDgk268dMqjZklCSpqhNWdUDnX8swKCFk748ezhu4htSW
/n02SLW0BgZung9+kyeQc9uYE4GNV76CqaiZGrzGRvd8fIoYOlNN1KKATOehOHNYKkBgjk2lVTgQ
oWMPjTF08p8QzFhRwFO1LNIpcRFBEP4sbfRgbZEUWs8sL+DcyMWVCQa+SSll/Fn7O7Mik9gEa+wP
+MT/1OmK7ort8kJH6R7uUHL+icNAH4tSFhlOkVQThXCLdvK0HO0i+SU6Zq7Zz3+5ozZZgqp01wiO
/YQX6zmKX0jpMMlNDrXMruPf3QcZjeySAPNaJWfHb9WeofeqdhrOr+6zBbpbuCaJmIajISxRcqCc
k8993wblssxhIhi19NNd6Qi/dq951FisMce4P5fANkEJ5Saw2mx7if3C+X41G9V4o+mr9O42UMD3
t7SaTyECG5use9Nbeb1nIlKf3FVl/rp9XkBzAh912cVdGEwHneXf1rC5SyOGnIyujrUK690rqwHu
lgmt1yEpPMBbqwoZEYL1FysiaeuEvTtSD8GM30XaSwKlG95T4WFgixIvTibhMIKF9zU0tT1somx+
jt+p9N/1qDyQoBD5XJyS3Pu4TI4i+lCFzQjRQXCXx/mixYOeRHgGR+rgYA4FPtyS3Y07A5AbEKT8
W3bzjqvKM3loDxnZWDZNvhhnHUsiONrLvT6ry1iD8V8FPtOV/XMuQT+0j83DSi5zEDoOV8tkLlPQ
b2fD40fq8KkxYdGMJ04afVjcGHXbr+rf+p8KWcuhgaXedhE1nbGcQvHaHhDVV3/wqTgt/7FyWrPk
6tdK9YzfqfTwRPOBBWq/h/jIX8p+t3ipqBctYRJPG+H+eBxeyYBtOh40ACP7eH9ibXJItH9bI8VY
7ieVrjAsfU8E9kccqxhnXrNYJFxJAbbD/o3NTTd+invCCiU5IrU2TEujyWCK/0h1XjBWDpAI+uqY
2k/Idh6VNTcGEeVq7YePcvO8mRhHhVO0Abk4MyPCqGaEYqJhMfUXEx2AyfekAW6Axjtvdv0PTCkl
orb5RDrxAv8UrE+O2ed7kPFqaGrT7CTA6XCJ9uHRkBa9nTbk0sfKLdqoBvgTOH7AANKLTzVGdRg1
bCcXWc9gDsNcOmczhL4OFv9DvoIWIK2v/a5FlEmrftdoZRIiLG5n4So26abdnR91zifEQYkBFiU7
lRaQaw8zKyIFeQaam8nv2jnB0IzI2h6dcoBsetZNIiGqSxMrmpb37JTUOfK8nAEULNdR8YQShBc7
8bZ4CybK9CfAlbEgyewIhciwi/Rneria9X5heh4huSCl/96JSJSC3Eq31SG5IG2QRlLpQmbma5eA
32J0C080RWFpSVzgoAipRa9HbZzksYJGtjDi3TgCxGOKH05BH9VilFezCvocllt1YMbOyP9kgT6o
JFhn0aL9P43DEuCss19890az3ee05zN9WwYd2LzgdpztmTVTW5AcX/R3JQL5eCEWuIIrJqO5QEYN
CCbL5JKqYNxBDuYh+m8kSGbM9rG2LYLowmzCQx9kIT7sobAnb3I73V8/mEwKNE4L5r82tyHPUnAI
FVlMTlSScQf1+SbAoEl6nsYipQcCJKDeYBtZV8GTbrskIYd9MNNy9P5qWkIc/zGWvRL+sZyO6K6G
BnpVUl7au0Y4OXeF+DB7XJ8ekiAI8MwP26PjDpKIxduLS1sDCEEdnu5xNGxxITobOidlnFtHAgx7
oi8gusye1WTsnhrJgHmKrYZU8DARydkU7BtrPKs+ZbNGMn05je49BQL8M+UBgUzJwUIpmswVEDD3
4H5KFayagik1ehWBIBfswKQQNgpedUoTZT8bIBDdjKGW+Iwardd1hvsmA1dpeFo1h/fELvD6rz+q
Hm0PEQutffwuyoCt/xrS/xsHYLkRASrAKx956wSVeO0z5POqCb7Q751Mhhl9+2xDhIXHTC7eFFUV
+XJsvmTxj70jQMDgiNvicnsMj7EeAafF7MGn4GAu1AGJxnSiMT1q8HBCFtANtjHK41o/CiUP4fWi
T+IA0yWgcIbVzOdA2TRTVmmZRU0vw7joHYNJhtsAXfej9ULgwEYlGh9n+0BoaSGhLv1TMWn7WKZ0
OswitTVcTnqn0mc5WhXezLQuf8XtYom4N4+xwgmUf9cy7WW2eVUQEvScUZ1Pm5GJjXt2MDOjw22X
WPtSGXfoduJ5p7N5bVq37Ddv16MX5DJ1Z0d6kBuUWMs/28NXPbd90PQBFMY1yi0GO3jNd0Uq9REE
NXFOLEZTflsyUdCOFaPHPeMDX7qnOzMvimLaD0LKLqyw6QHMDT/P/PKlw9IDPiJXz8WKUN10DL12
oD21ctHRcW4k3Ez/nzWlqmFL1nXo1ods681mngS/k0zOqcPzZJN7f3bwr0gUvtXKF76y11dwadW/
CTRi8XsvY0Ly11GWqDaM0mTSa3MsYkUR176OKXo0LpnO8V4hTyyqirIe7bBQoC5AWTR9doScSMEz
yYLB3iBHb3x3R6TXKq4IcGMbsacCtcSbYdjPCaeJS0W1Ja42rgfnK/HLRFpDXdf/4ia7JffSczYo
ziYYzLZJVEDLXti4gvnnDxKqrOR8pVTY572f9mNN120c7iHflT3dd2YTUM3uYKDYCNjHtHiu/XDq
Zjh+aP9x3HYsCLGkwCmgRc3nbwgHae25sH3Wr2R7ucDYIaRoCLvq0pQeWRRqPef6FK5zI9Hx9Hdx
Bg/7/RfowIwVbuWaJWADG38X75EXrqhgxQXc+TJyRX4qoSK+VOFvXXzY7OJc/Df5/e0uMRWhfrsH
yJK7Chv2M+eN5jMSqyHwAiPP9Gzr6uhrzSXprQFU520IhJqNHTgIQE+kaVsiWwAWfcqDvhVN3WgJ
oA/ZI+fe7+r4HxfFC9u3Na6sgef9yfhKOJjyb9jon2gLwZ6odAKLJiXkUiix0AVcMnhZkqpuMCaa
RU4Jsx7s+UEaBS/5jp4CKXlk7QmKsQHXiV2WhZRkIyxMJHsfzROQwK69VVv391skMYYfgENBSzcy
sUrKcIHbVotAoySfjfDlJpWF72CuyUYFWgZW6B119lzZA8P2uSTzDHy4tS/4Yj3KQKFuareKrhT6
blfuLPLIpeDKoSCzmzqYtkgPLYEeBZzsQPzQGw5yC7E+97onUpzOtowuXn5Tp3s41Yuie70JBvJp
eBsDOJFxeDXtWjAZEMjxintGVO9ihV8W4ILm64N74CyLFzV668BrXfi1LejgBDuDQVynLBWhMGYF
gNg1Qc2p1U/hpFW0LdnAkEjTbUoJaOmgpnKQypRCml0NcGLg+diI+ZQGljaIpzgHFuecimwgSCjU
10HHNl8wQx/Y5Rar895VELG9J/f6o2XPCQlezXSUuvX6z6O7kMPZUTziXDObDFuw/nXnlwSIJsv8
0wqMinhbzpJVDhow2gzZB/4msJ8/DN4lPkC6Ch6Hn8byezh74gqww/14rgvbAxhqBcoXiDAD17b4
3qZlMy6+o0qHGNzMoqsVkFRm7ZrLCUbsz46PfaIvRJB04vXKjvfVF50aqXE82qh2ICC5neu0UbyD
5QhuLnGiZGtkPxFkPnfNO5Dl9bbUBc6yGa22gIjtvK/pDk3AEtXBu8UlGlsVI3NPdQxJSdEyIa9S
BeLz0l/p+GQg0CZeoj0Q4wAV4HmC+KGUekPZRAA8Lp9dgHHqpgJVXuCKAsCxrozzgbjMQ02VA1XV
fUixCZyJyGB4/RMh54zUvmF5sE47L6OofcWKEkPySsJVlC9k7QyGcqA8BdMHkwQi7Et1CJh0idea
sVOqeRMiolrPradEUE6dMRpRfSYvUhdMkGlsU85hlVHGeT+7+KX7yQHNhzgi1ZskiNnnMTMHb5VB
Hgb1wEYTsc+N+CNJByCHFFUnYclYCY2aafDUgwkgnIOY1lyKq1224C7nMqnrOrW+f7LRhaxPtjn5
QIeOLuEct9omvd8Z+uk0aLmTbNlodo1LU80c5hy+glsxcNj1/H5KKierkTtJbTzlnsof5J/otjy3
7RLN9hG7RqVmQsWg3iBaBwOVYKrpF8O7m8VjvCSpKYeSEoqYbfdc/IHu6JWoOvtF3fMb/HFICgwc
HnW3a3fOYRA964ZjT2N2HeUDzsd2Md519fbDDJAaUS0oSBVxPdGJNvAXgGj7MmekA/NuAWiOdbAC
iR/H/o3c48Jw09G3wTMTo3brtgzQJ2QAnVrRFBm8Wac7NB4DcM3VE+IrEfwq7T+XK4RiZdAUouiN
TQyNrfdWdc9pqsZHrxib86TtVPphOnUVYdAQRANvbREVGzZGwPuQpGa2u+3s1RdNQ6xSc+CK7P9X
vx0Z/Aqatbuh2vd+lxYTlMJ9vJWe7OvY+1avdxvXRvhBBp1znanYeRdpazgWyAs+s6we9lqcGO1G
YApZYLYt2/pvCuaOIlOkrBcq+8tmORY2KNALpudCVNEKFcj/OMhPWnbNe9c9MPYKMYJ7+gKN8K5R
QQfKhrxkqly0b/V6b5YNHugQKu3ecDuIdZHPxNxYabteblTmHOQfwAoy5y6dVriCss6+a71MrnV9
LThTGsulaWmgx1J7lxBIjIwFzwUyUpRqKWdxMT+glUqqPl/U1UibhLLFmLNSSGxq4PQX/KLwa9nG
qlXFVRF5GaScpQiPx4e+5b68/44GIYNsoAwKdZGZbSFSxPM0HS3uQWgEkG504VSXQUOX5UPjnurg
bkWmKFlxJSYPxc9DsOlr7prw3a9eXGKMaiSOV6GFmIVavJpAfChksU2LQSWH2Voq+mLkaBHnRXR+
X1MW0aZuE7kqwiKtvhdUpQT8ILGyElHpo2MVwiAoBJha5kH3auB5tmiCSwmYkiFyZm1i9rbo/+wV
UILt7chPhBpUewTF23rPRBbNUmSDotkILfLh5rsGa8GEqlph4f5lHWw+u9NlVwDKfLO4bq/9vT7E
o+rMYQ01tBgmLmtrBxGgd+JxlFf+zYq/vh/y3Ie8jASOmnNxNSISQn1ZsSFxeGD+lS3egwwiqvxK
SiYQVPKyBIcR/+a7dSrc9gh4zvcoWZYd+/cCKfhW/NWUSIGYRxm0G6z6ZEkoECfZJKX3gr4lUEDc
Jxl17angbYMiaQC0FR23Ko2BGffPtSfLWKczAo6Q1+s8tswztRy79H3T+SXOBlse98h0yF39eoMn
3rRDIt8HzFA21iqC2M+Ml0qW/z52fIJhf5++lzXxvxxhxFFLQfaCeO2yvQInkqAzqFI2JqNhHwYV
wxo+Ld/wnPjk3L+UThTmQdbxEa695ciVzzPwuj7q3sM3V9yk+25mRLJrJmmKYP3KtWUFE+MQFYLz
BzWksyYzGolrHpYqbxqT2XDij1bXxk9l80k5ncX7rseEAMIXLCDkFey+tIUbu2xSpm/gxbzQ9Vg9
vbM2+gAq5db2r7gFG/5VZmiQWtcEx7pDvikxZkzgKqdcCgpMB8cjxftz613zrp6xuiTiZTtBdTvT
3QRsWpNINsyQHAyjHf/28C3ukSGTJPVePI5le+8tCUWYSkTG5xOrpxYsLs8C9PcgJPaNOMsReaE/
nqjWpw++LA/WwEvDkYynJ189ioq3F6CCUIV/R01ENQ1VXyq63OHaOhTcdcM12rm56QBUzq1J66lh
F0RK+axJzhF7AGoMc+TE3V1FvYXvAm9cPlbJBCg3sWMO8YbF+b8xaDTMEFpVRsWZaTpn3XXry03G
i9fjpiojha3DaL6rUO5YF2NpE/ZOeqDQg2k0U2CK+0nGYZZ1hO/Cvu/M2lVa9kdcaoe829zD1EPC
tPCYV6gPaWLitE8IVqe5S2pegcjULJ9U/nfhVhGsWB72wgmsMLJRq5Fp1Yo+vENzSxX73t9Wpt00
vfZ5CuBovXNWQEga1i32Il3ub+rdLhtGVJSdCXdHbsbBL+F9dNWHsXc0J7Mw9E5nOcoP2hlRuFuv
K/TRgum8vKSYewgY0cO22DWNzMXOEqOZO12LUrppx4OteADltbQ7wWVBQMpAsRgp1rqiWXH/8P36
xrHrWiWXKFhLlZr/Dn9GDRpXm2VSWnS+2aGY0p9+Ee7o1PJyGhPSkrd1iowzHjyXrknADey6O5Zy
uTxA6p5Q/HQDwNfFJNzZoeU0kNMXX/fuliL3GfLp6Wpd2ghoe/1WQiE9p1skGGoI4kSSTqcQl14q
mZa3ocCU3GP+Yags41v7z4D+2looief2Btfx1GZHmdT3HsayheiK4Sfjkfk5EGR1tqCYQpzAAOki
jIGItTkhYOT2u2c6olkOMOQgtG455M/NHTVzuJ4YCjCSgxeYke8W3kvLm4dPOw0w2d67hW4vZv0Y
lEhlRghXtpjEjsaBm3eqbl/YG7EBODZEnHCCJeM4J4amBOeGnawZMcfRy5nOu2o2fvrf9Q1rli/v
y61VPq6qvErfgCTUq7Lc72BVQ9pRuEKp6cjmgsDLqPTt7o+A6Tl+427Jf+SyjVufWyifyWksQUTv
O1peq4E5Lx9GJS9geYQgYUWQkuV4tDzo88KPgfil9Ak26JFDia68FtefelUALWqLEah7sm/ADd7p
zcwC80Y7qkfNEDuaI6vMm0zr/YEYMYzrZsaDOQVJEVhZEtn835AVsyM3k42MzdO4CK7GgL9C9fiF
S+ZernBWLDN+xSZT//YgjDTYO7LTsbJpFcCRwa4eeCFpnVbdqP4/s0RRntIAdRATPjvezHZS6Yya
zOsGnZbJlh4I4ZnKyVOBq3n34S8JDFVP713w5BT5Q+60IqgPowNKt1HXntro0y2HJJnmnA7vDuGo
hPL08/tJtEoWcqfuO9hl6RurSYXQ3PANqnoWDFvIVdq5kKyLmmqU8mu5l6UeTd9Wc+ttvSoRhcHi
nwMDbazwfIjoXjauPJIGIZcZgeG/2Dup0snFy1n3vNJdcNnEU3LFq0J0C7RzwwS0hh1r94JRP3J2
h0F6RcU3EMGVly/o/d+gRkxx+hOKL/OlOQXcRsOvEYa6Z2xthc8u5yZjz62SLE8GBIlFPTnOMU/r
X2twyiId7RsjjidtTRTvA9NCmzFAZPVONpqF59rlWZB2ovBlwu1U2dLIgesAnOjE9NStVzS4A5Ya
0SU49FWL/tbwohMIsW/enBCt/1gmQETVQLuC5b5Pc07yKi2gW2COfIdyVXi/4vCnxAErm9ZktMqB
ydAGW45h+RPGufT7ul1M/Y7SnC/bMMKPdkUGBvft32KYykWIMRT5czH5dYTXrbR5acHQi7zPii3s
hLukSheNJoyI2obV+HmWliIDvb8AAicdPQx3lSXX1FmXGX8hR9I3AMskUtMDVV+qxrGF9WPD2VcG
creTAKHE0+4YLAUjFAdmWP6yz8WdCEUO4HliZSWkW2jPzmP/FNjoW4sgsWIMy4Xou37pXZa4OfRU
WcXjdhC2tLruQBZUDPnHXf0lNqWMJHwEl2FohEVzNhVgVbjqTOQs5J6zZmrxZIcsXdVnSQmreig/
Q1dqrZnDsdn+HV7CROi8g8A8t/bWsjbZN2LWS47EXJHRH/yDSBpa2MO5M2vFK+g+zc1WtrtnSItN
G9hLEfGuowYS1vIQM7px55jgMxzgjZnxmJf5M3tk0ACxNgoJqLL8kf9XuWy0e7/HZUkKcSdgwzK0
QcAd84cnO6mP1VsbYaqvs4ozJ5Ya9dwDAhMmJr71feO2bBGBGO3pXfZJDMj2Kqtctus4sb0NfIkt
q3/F7IfzHG4SEYFUYtzY9EBNte9NNNdZN9Dyya2D/ReTemz3ggdcgyWEWNdGlsS1c7vR4hfyZsa5
h61Dws/ctebN9DYbrU5J2nHtscWhxbj+LVxF1jVqrZDtjz22BF7tHsXh4VqnHiJ6SJVmqnLt1gwY
wpGoE05YYVRBso2xxKrznWWZM1gMvYuy5fEEbN1neFblu+kIp/lTJCMjXdACBNDSQ3+0qZjtjGB0
nmuAsIn41edGHd1mQ4dhRB7KTKfHWKbxjYTF5xk6wr3tHRI9ARpWWazTGa8QBsaAS0P+Mbz4UhDq
5tcfx9aP4614xpBrzsVW3tAq+RP/IsdglEOwknxEAAah0vTg41jMgKaNBxfzZeyQq5b72R63vAyB
3Th5izCnR+PdYdoKmdpKLzOpjzCZL3mTylaSsKuyVzT5FPRkuFLY4Ey0muOH8Z41fJ0k/1Yk9HEv
3ClaB40nc3jCOvUvQL54ZXMpegZp+fvQ2Ns6yRp9uIihuPWnMPzrj5fMsVqNGTL4zVnuK2fxOxhp
OaYZ2ZlyeV8tkPX4qeZ7/ZxRXSqIjcJ9qZYWNoCiPw5W5Ywo/2tTMWdB2ngl1iiGnXr5zK98MCYT
G+8aeI5mMfhCluZvws8sdPWZQ+/Om5puzfggwFi3QrDS1B77WjaZ1md2AER5oLkxK8Mo0oggdCEF
KG1vGxso3g8tZj/GMXUbQdvPZ1BcRe8PGZqcxtMM6/yPyFlyxTqQa4he6sL0+uml7mFytMvx0EgY
aX76m7T2iDEtkIb43yEFRxDSL+W/355pnjCM1g/i9ypJ28OTMTQv4K5NzJsabJjH0sORFVsPSsyG
OQ0TB4hFPXa2Jp3m5qXcmBcAoA71x5I/7/IrJHDa0z2A3PLdsN6OkBMpfTPR+TewGi+FcnsW1+hd
fzBAOCk3uBk0I/aTN5+jRZB69/dNUXHQSpVCl5MTTS5142VjUhhcO+g5a+oHbWT8kEzyE2j6fRCH
0ucsYJ2WJD7hgzfoAA0RRznQk4sP8pK682xjm6DuKgSLEBGSp0SCev9W8PYBgb+tM49pTwi05s9z
03pK2qAnVLnIUpWji+cASgzaaza/n64B27gZSn7DdZne10E4VhXlbcVBiNB/3G0BXh+jKgRv39vG
o1cCVKQi+c/ETxq6MCzW41+TI4yHDvbVIR+ELCz2UyT8rZQnEDM72iLsrHg3ZNu28f+AjemG4RyC
/rpS2ezsJpjtF7gBpNkbNXAN5oAwSTjfirj+PhzQlMdou7HfKjeY+UXhwQax0wSrsSGTJR21JZ/i
OrywDLy+5m+EdIRLzKPyEk6myHKxGeVncuVGQDpQnl51gYOLN+EgbhP0k6S0pw4AOtg1okOj1CAE
lV77HzROs6LuYKojDFtYHwu9qgJV+zoKpbNTcVUTK5cBBjBU0TSjo7NoANOaJDquyTA2AqbcwAEd
5ZzlbIxkjXihqVfqN2v2Befctq9aAJ1Q1NqMnjiuM3a5Kex8gSd/y6CH9Xc546v8x9U+KfnvZ04j
fF+pkdu8YbBnMIJ5BATZDkeaBXxs2IVFySdkh3n58bdnBz+CixASA9xVEnigwtrpYncQc8P3yIM5
cb+kR9uZiqazYI58KJuCOHYtq787tC64soiNUD1Ue/lAbBA+knf5vtP+8YjT8x2fj9ALdlt6Gt5f
FQ+ZhZ8rXmcZrgWFp69gpYFtUrj6SqWlgWKtnpEhIFmzHNyR1Yhk42voZRosf6OHtfCcsRzUY/Yr
hwMz84cQ/zMfqQHi12o6XeqlI8RYPlrA5TmY/HZF4al307r9y0anSNyUDI/uYk20uPK9noPcMUzb
qESJ5MLEUZisvY3poVO9OBEEAjR2Ke2NnpqBDhRvNNIla19FIbv4oWEcLUdigu+BXTHEFRcopCo8
vrQcBax1eJUYqYdPSx57jby5vIRaN1pwDPLGa5fFR/3zSEDPczHeDYQjDNVN56ILhhXx5tuUTmyD
Q0X3COVRXJFSbvEQ7Vhx43u0buWfpYfJDtzdT93Eeu9FlzfXtlJ7BK5yw6o0MUWmrtbwNz4V0T8V
7XBkyYT6FpHNTUyO7HCqKSuH0Wcn32LOVuKNCLdcxlRg12U/3dX1t6HTUA9Iw+cs/5c3YiNuVU6i
MUMpeztMvBaGTKTGE51LMMd51NjY3o4riU/uEDk32LZalI5Pn0f871o8USC5CCn/+NJgMLw+Mvt7
UF+xGbqf8JjwYF1Nb0id8VT+W5rtSGEb+jUPQVzCy8sWpbAEsfiJMBjXiXo11yOWcCpJfIjKSqcP
fdKKRb7Z/8QU6UEEXg9L6sqCXgvXiQPQ7e2AgfQ8YOnhqDwXtKbKjUKEKdiBJIsRdylyOzmvKDv8
oaW0LbNFE6EMUkpjjP1xXcLaN2y4jswaA1VW2VNyuyVsLgb/jFAkkTx8q82NbE1g6fiOb+b+dikN
M9Rv9mblTg6B7FPXXZEYa83nlD9XnujRMBWvYF+q5REVkTWTCjXPToQ2TqVWLy8TQxIwWrmCAVqv
+27Bj2HN8WG9kkA8v26vZhQG5diRng/FZNcEaI+2YVEJWBpQOWkxxE9DdP1JjQA0XRp2vX88KVRu
wywD/1oY3Fn7WLau5hIuxbdTWijgC0OMhIfs/kU6KzFvz+pScmiqw6wb30DzS5Dus3UhoGQgu0Ey
FGq1gZJ12yZT8enGfQqhLTNaTGa/Mc7b71ppaUn7zovpFfXACevzEOBWsej6hdO2DSXVGinVfi1P
4FCRodLOBaKzX71UJuXyya2xPqzedAnxocZjndDvC9RKDRqF0PZoTDwtHi9R8fiZBspGzWO2n9fC
m6O6fR5IIE5tR6cJrzqs6K+35rlFtp2liQr7C5KodgtRUoRSHS/rZHeapZqezsSYHKV9Yd6++PJH
ZLpHzoauzmILH8W1+vJ8C0/ugh76Pr/KMuLYI4jkhzb2VqL7wYZ3RpuXJHLVAjuEu0DydGPtiMRI
TCGlQoJAsbD4UFGredHq5790helWUOFjOLHVHLbuOsVElX4cZ5RX/jDkScjphXXfIhm91gSiw60E
uD4IwQ+3JGwaklmLMCozDpQgASENAV3zyNjQn1zajp/IflvKj8T4oTkFzsAeBOSfTnEstCP4CvoH
jj61K+Fd+iY300Uo4H66TlsB+95ScLsoBhzf/4lB3HogC2h7rQ==
`protect end_protected
