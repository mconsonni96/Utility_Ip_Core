`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Q3pj4Ia0otxsd0gXZkt5syd9NiDLgRxapedfdV5qoTIkdsvgbBryOOflmVNhnkJ/hbIg2rqeqK2v
hKtUlm6U7PhmSTlz/EFt7z8W3zMHekHNsDGwnah1jn3ODNeo3NPEIHczGACFqBfaci97etMFXCSV
GMILyjij4n5K3BD9mAGpS073LcEoKe24OpyuLlFYB8pVF1z6bqmrQNwufs2WgjOy8gOV2k4sdpGM
d0NgJ5RRqqCADu7AxjNzsfpXPtWCEPP5I1A6S6+YrAi+SMotBvOmGdF8m7Uc2oQdSjKOBrrTTh8X
cU+aw6LieRXBJNgyh1tmxen7JuP/GdWS9aIGiw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="CEs0CxkmuEoLtryMeMOVJl54/WXTWvqaQ7sHoP3tWEk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10160)
`protect data_block
WorbMdZLYtYvtW3J/YyZZOyiyKG+6Em2TGtr0mBXuRo68982jGhiuhXE5FpkotDKhD9XP1o/WyPc
ND+RlLkATlPC5Cg3/jD2cSxa3s7IW8ONBhRauQJwcOV8KxmZrG6Lne+VCIQsEZQFGhpIw0rCrr7D
9WilENh8E7bPONptGzS9iERbvMkVXudZIgMVJKMtg6CLM3YH6dYLAVPSDg/+PbcIUJv331G3Lle1
AyG7beViZtYRs4xMR3o1CG7vuPqmmSdVgV/Qy55pNZSKW72QzqfJTD9PkafLZd7HEM26nEMmMDPr
vUmStN3jJRPRPu5Y5aW605/qR0fnMMZ4Abpvk2lFxPhg8T8qD1k3ADtadQOb2lduKlqLrDtJU/uL
I5cBQuAaQF56FH4D+GjC/hgh7DyXM3jgYymfFOAs1vePlNgs+4h7pe5v5C0+9hvDhs6eks7S2Aur
HZMPBz7fiGNCATgCdM9641LdPyl37TCczOoUDs2teGJPLF8H66FvWySXGwWuWNjCZWJ3CccG7b4y
fIYNmvA3H8yuS93RaBvqr29k0LouTLUi8y76JcReWWEvaQUFAQK48FV7R/JRcnPC5mfERcCdfvQ/
4rOIcP7+2NbqyyfC9DbqWevwMESIRe+Xxyipa+5Az309+VWu2DPT/1yW4TWE0xMertzF1QeGjol6
VPEiSPlTq53tnQww6g1EjPqcf0V0rf1kEjX0C4A4k31ERzcHjKMZNzfSdWbOi3+2yVPu01fUVa6U
LcKAgciB6d4XUeirkx+gp0mFXE/ksNrGavZMZgJIj7dLK8mAN+nt6SZTkPb/bq1MTqC5zVZY7N1f
w9+sF7WhqkTba1UhSU1DeHGe60OpVlVLrsNAlUI6iBsWu/rZ5C6G2c3QMw176fUYr7Q4C1acweOf
ZrKUOEAW/KftIoBuV0ItOdImluW1hUEVestWDdhKw781kTqs75SOaKVRTEzeskXc5j3Nin1fVS4W
V3flr5Elc+xfqROG4FGqqpSAIJdH0tzlaci5YiKOU+xae9W2W9CmSQM9PBaPepV16Rg2kw2BGp9x
vG5iXK23N2HBn4gNB5EJLlR1T59UNa7Bq7lunQhyCwglbU0jZcwd/19+GIgDKB83WHh7qEZPIzDs
DIJU0XMyuvg2zWZGmRfax5IzJ/uDqmvyvrhswyw5yAeL6cV2hc+P4jgx8xPnr1aEhe3Atxo8mNPl
IPyRNSKYg4H8XSLS0kKcWDseWizHX21UW0p/r09ksKg3VuU8cuoDHQDP3V3vKoRHGq0cY0N8PbFS
5QX9+UG9vcI05nT5wLh5yA8AxKoe5CdzNsVXNyA9W6TsYRGkPmT+y+OvQDcpVGXrZmw0eeH8Nzo7
J+xQEI5zQXRAwGG+AYQIQXTCUb4XqYlqa5NMPISmfsNMx2FMEjrUN2+xAxBsHRQw74VV1Gf6bsdh
+gMFCYZDUmd4FCi9+E4VoCyZ2wI7N+Aex2nWqA+XhoZZ4rPrpg2/iD7FoZ5qH83lCe4B0MTltNDQ
xJlCWORAmAxTzDpxMdoGtYD5KGBWSgq5hKBytlIEFdnuzbov9Aqr5LQs9GdIMsJbJ+Y+F27Oiad5
vWAFRm18NrXDQCClZYkBAOP6vegz1p+qPfPOteHLTMqHDKqpDXQIPmeK64x5FvgkWU/CTbkboPIo
ksCkRIt5H6HXfdZrknNGfaDWNritYbixfsHjXhqa4pzCFtb16DHoYdZ6AdIRMO22fLcaQ6CsHOhl
mnBcXpX86yNnKefSOIW6nHEjFsg6YHkhmYw42m48QdBVlcP8/WiZOQRsPpllN5TLB0ZTQOAygIej
qoQ0bL8tKVwlMxuF52dnwOEnmZfZ5fBcLbRr7gIJy1jiu4oDFbeg5JwHodtXKwkli6fCZ5rz6XMq
Vf3ezV4/U0/tJ6PK2V9BJwix2OGeOnjCK677/ChYr8vW6vUgZOB8v4g0qxmJRFw9+oUBNAKGmVX5
F/X4hO7NQOPnnNGo8dU+fg9tH1QHPUen83gJdFgr0YQ1GHua5Wb3DtlmbTZZD4FG4fwXkzGc1mQg
vJLfljg938uiMtE0HztZiitxD2OUd3D226pqbqZY+Y8HMucXhAJkOLOHqwSuGTt3XK+fR+RPaPCP
AYk4jKuDq0tRXAL4Uv4JtJ5FZf0jOX5RwvQ+aywIIQClCcPs09EcEyIlmagATdAFZmKy2RULjwGA
R8495vaHKMEmcoQT/C6pEOeHHuM9N3yMkt+iaqUzVWPcWWALkdCn62gRSZ9EvMUrILN7IYU2SsPB
CIqbKexjB5OKcMLrnAmXAi0dg62jc58MUyx5a6WJDgU7XFJcLJm36Pt+4vRTX9XoHoYsDoHxut7F
LQwCU0ds5gTxoRuoJ0eh0sXWy/xZFffjrpXD37sNZ9k4vzzgVqB7JcykjkxmPR9eoHegy36t5qmO
g90LSr8VGzKclhwaA0HmxmPYpkJNThyNWgL85s843bDK4oxFQBYFGbnuPnTjC691gSDJ4ofoaZi3
0DbnTut0nFFr2gKS+QOIUiJJTUgjyWNv10dXknG/SH1I74hz2t8a/X3oAVpJDvBKmThKsJzweMYP
9xpirhCuwr7lrq7PZuB+ArCCjPeam7BGVJ0tLQ3PmPCmCqYdX5EQjwlDHE/TVT62WMbR1YkuMqQB
XjJxgNBsrT4qTp3ius8f1pNwq+FBk4AsECn3dK65BqNHG2a4EaUri3x4bOrmZPg/xIeigS9yFmbz
4qQATSh9Dyt1iOMhUXcDtYuk/55EPzqYLWUG8MVwbeg7HKvhue78PmtBVZi/e/AY0TM3kXi20rfp
NMUiTuRrcnOQ3ic9CBt+tr6fljG90Da3qiOio7OTySSN9+7ASfud/auH7are6pYXoDOOrQPpwb4C
OmQv6IqCgemeSTpJHDIGL2/vsddf//KRqXm6GS3Wj30VyZvu3LfeSLhw+RmuS5U8LsOtegrRuE4X
a68HHkDAxq2j7BVaX7uNshFUB5fKbgvAIa9v9oNNZCYx4/dN1NGLVi6CzSZIiv7hJM1KXXCWjdtB
zxQpSRjIMCd5uqnjS5gNDIdLxLDmyiZlfMi1qiK5e+HrLIqJb447UJuWDKCEmj3fSbvtmKqkIPLO
sn2RnVyRmnl6XTqQUhJvTs8moMNGHl1MMgpIyORd7swaTrtRpfgRguLgWI+jpjIxsPpiV4pA+/pa
mAQZhEgOG48xnZA52KwQV9GQ4/GiuYqCSQ0LR3BxI50q7MbNhDPEdALBaiiW89VcOx4wWkYbEznq
PusOghXKRxqZt2mUlroFzOCXr0tspBqiRDanNfZrFhMd5HBB7d3uJTR6Vhl94Pk/gz6iNqHzMp+/
toBEWnwWzfwG1Wdpq9+MEyWP6q5d7vSp3oORKFScc7JmaNJfurJcTk5E1idGHs6CU8Vc8z92d06s
mzXYJAakznPkj7s+esKTsUvBt9J6kpAdNq7SZE34n95L+Dxmov7mxeb6Zmgs0VR/X+a3ZHmOHWkG
1lBO1CV6KaYehXOjg2rByJCB1sQ6zHMI8C+f2h3JNCAAyMsVeXwiR/FajJ06RpxmGp/X5fvQxNxP
i+IcdEEtdtV61BW0dELSZBEvSD1f4WESwTp5doeVl4/MD0TtK4FMT5dJxDQr33Lq9wN4ZgDr3NY1
CirBMhyxSb38SCRSbVhGQfjI2lly68lkfMyWRS0dFoE2xBjTsX6y0mwohGyvB9NZkJjLLgQZklfD
l+s10GF2wBPucO7EM1LH8hTSfpf+xwg7W2aPjRibK0S2oGZK3kEtOD6xAA8sSAK8Dj/go3aObaRm
2jTp8kO32tU3l2KY2duIrpJgNFjEokk0IKQIrjEaH6a7JBG4DBobT5xa7KngQgrG+aI4g9Q7ITh5
HMU99K72C1cmgasYHpS/d9PfVhzbIc5nCNdtTZpJwPjK+J7MRWkb6zXgkDCPk99zecwyeFaLD3Kv
KxHF/P6M1ADMKLRx/SKEiY3uEoLrtQ5Kt0qwVvtFhuxQ8NARJ7gXN3BVJLv4VI3dHH0zG+SOc+KZ
7w1nuAp+qf36/dl+6XWCILvlzmNKs9+RvHWId7Nee4feMaICwPROL/cf6USfQGDrxYvSxt+zH84l
oxqujbsxDJu3MBcWS9HinlG26jS+2a19i5lRgYNH1jphrqxTu+zsy9EM93M3gxJm3OIMSEuYdGQ8
seTVUi8pkjOgL9Oi3Ub5bYCCWxcb9FErbGgb0dQOrHmse0RCrKxzVtFBqsZXK1luhq2cl4GrVBvG
i2QRZkK2RzR7YuqmnqHHPOSLRnqyFU6flDbLPvVv/mVBHSNAUEb8ugcUtmnmK557gcAbVczaNAQw
ZR2X0X7TqunIhhTwVpRDQAHsOE70QkLg24QU/2bVDscEUqls6cj8PiGmOV8a9+iTeK6rBGeMgCRQ
qemPvvMyt1HbboO4KYImHUCU4qf2Wjd4twBZvoEQHLuSsW+vfBBkgStsartZpC15QQ0iz00s+WNg
3izGgGIa63G9vOI6WnoGYfwK4uJC5iVkARLcFcG4yxR3j8lImx+uAQiPE7fYbXYHj0j3BPFldYsN
6A5PcgUE15YZJt0l922KVLp4ZtkdIhjjTnZDqQI5eL5NUUN5mnuzzKjsWF45yg4xKrwWK13bjHm2
pX77bgve72pZ4w93MILN8ypIjNSYDWWbdl+dgD4S2EzVFk+r8Exnpr43AIAMAhcgQbCK30m7D8q3
Ya8kZmFHTxFScj2RcTSnMFXHuD8e0YbST+IM33kXKHfxzHkS8swbzsMb1Q9ZZR62bNWjAyutg4u3
AN28RwrAetcDPxD8JecrhxnquFe61g6NmTgUMNbv22CnFS5t9FFK2kaOiexvyWQPsJdjDWLMvTVN
59B/uSTu9lgW+7/C+zD6COcu86wZ0MXGBuWzOIUSzfZCeRNOlyT+AfpKtfHYokpCHx+GksJfOJw6
rF1TOfAe8/h/EJzP5IpM3YSRYzqq7sYGZvTdJYtKQoVYrkGQxRHmcaAvJw1gzl/3/I4jLJJZcPqV
zcfaDVIzDfgxrbAtZ31M6rO1hpcby6+at4jv+y+y3RvIwyuRBToRfnxLFHONVmMG4oN4LdjqnpKE
eOgOVOg8v7ThWnlJG9BIV8BWWulr0AzWWuNRkaO2VrlU136sszR/QmDOWQlIcWJOmcF6Nnq83Jrx
c7VzXW6RklmbHTZTJBXOJpTMpQHpgXIFBhJjKJG1/AIYTk6YBfyCv7490ifk7ofoAdYNIEJTokcS
ZfNUMeTxGsKMI86s8RQSurGQmxK91ZdfXCoImBLluGJu1lEdoK7GkN7u3RrgRTF2mQRJPqFq7tK0
IpZg1sjDvz3iWf/FOqNC50rXXGl8beSNzkUhd8ZO9lrwO/2Amda7x8Z6eEwaaJD9h3MbQy5qyjdE
1lBZ03HkxnA5aqxmnLDPC1cIL59eSbZzGTdQ35SvQo6P/+dfuJ2UIdfajyUhPQOakbIACYb80Unt
HzdRTlGPwc3rP4sEtprWaZfqV2rMM57ccizDyxgD9Ek6egPW4awNxz+Rgbv4AyESB2nArA5IA2jS
Vpz9EKPfTY/iLDJkN/qOOHPY4Pm2omE+hFU5xP99NelDw/t6fCQAgrZzhfG5zdS79b1sqLHoVnV9
TfwnXtktvGjBsHId3/7w5R+k2amsoLBYvyJtV2h/tDwgAmOZMgEbMxPyjyN5rX9LT05gc4opdcZq
z7Rn0lEw3tUlZAYYy2yzCjw8/aeA3JDqOkEAv2iXZmuGtQoLMVcJzTWeTLJbkB+SAO3l8mjzw/oo
ZT5I8vf/biqHL8465s4YYSDnYzmDhtad3vAHfPa+hsdzpUeFrlqFvxTMbuSExiRPg2wUxheRikJ7
zc2vpTHuQdfzYecsWCi+9X/dzu13yd2pl3xRzIJMpqwHwvp6Owik1FMzdVEQDv9NKlmNyRLI/tZY
HOxGgRmbWQ/0fMJvVkOOJtyBz90hfu0tZWpyraaE8WZndIkI+gY/h6UM0dlxW+xS1g1X3FQ5zabI
yEiwSD6KvVcNG1q8qQq9LGzRVvTp7jGbeX3EmLsSVjypqB+GRD0/PuPp8Z5Jx6JO8FeTA57KptuU
S04x3omI5Qp3/mQZ2zVaVcynV2daRZ0sKyqU7Vhy5pwslVk3/rGwvL8PRvdJnVDTkN/ukdFfq22+
/efj6b/n5rIcuywp8xXsyCozuEM+PtyvMhQdMSLqt2yAVJ/BDTfHF9duJhPMvOIQndLlnvo8OnNf
+zP8X4nwYm1WZ0YEcNB75nPe2U+4/GpmZCjdWVuSVdMjC6LAExDD1AqmEAt2tKhMl2fAQxqCoB2O
TZDBUiMF8qUd9OclhPHN5aPT98qkUuxYsMtgwX22MBeMU/uyblaWeYO8Sy4cKq/VWHWpjpYkIL3w
SlfEu9quRVtVgZ/9t/t/0TsBhJ2TanipAMplZtVdOg7V3CKczg/+mjHBLdO61Rh7axOEs3rBqAeO
dWGvvu+vmIWVQZqiLerOBlASgYXUuLv4QxECEA65faDr2KmH6g3qk97n/Ff/OXPgj8RAlY4RvNlQ
fnMaENqEZczVJOPZ1F6BmaufxtZij3figTQPQfSwdpmc/Q2Y3ASxonClvyldZty3i1E+CL1oRLco
qsgh6VrOdPhG6YQ2aviZqFlsK2U+ThwzhTyuO398z9GkQ48OCzVlUj2PtKChmubcK0a/Af5U8Bf8
LzK/VzKwvLuMyRYwjeWtrP6KneO2D5c6t71jPHBK159uB51kQcl4yvds/xTpq6douVZrW9r6YV6w
+a1SmvjNN0bxWbZwqUmsFzdWwx2xA0nrtckW4BLLsvyxbP7sU3yyWyJqYl7uKOdmTZjaeH+mCkXn
niqv6Bikq9CzxSS59Bg7Yw56yDrb9zeGlj7buLKBWlNJ993LmYU4VUeOwLlniID6Z7eeGI2TQ3cy
N3iuy4n2FiKUyPTJkx2bQ1Z13yieZx7Pe0IRnLFAm9MslmfQz79yZFDjA0F9VhP7okq52zl32MUm
NpjE42RhXSoH3tNCI99KKT1ctTXduZ4DbEoNFPUSFqraA8074hb6B4I9+ssU6d3AeQq9P8aXihef
zJzjyJFAHbYNstTVhzeJQKZd2/Vjd6Gq94fEtlaDLAYu0ktOUSB77aOjLj3qwzs9Jc2cV+tgAmBp
qJnlbNZAcZonVcCLRjxXI7mpucqs/WmKu5zA4xs7oAYXTCuqfv4pUTn3djtHsZLbF4OugJ+1P77b
5A704q0qIKCB6pwk+NVlqX+1pXOUqjqoneWyCmR+aGDIySvsJBil5IOdH5sMjN9ioGqTe+sryTNr
GJnZzgTexbDqHjfyvMBRKBfv4IuicN35wabjSt5Nn/POPvmu/k6lOdinF/413gnZa8q1HzihnFmi
8U0JeU2qan9Lr3aruaHVD3vrWnXFd+h/k4Ydy/P2OxNCtsgRNcRb8YGoxwz2ZNBdUJzqa8CqNxJg
HC3RLDbZ69jco0ckGpbrXd7Z2PoHmuZ333U+OPFb1xSaGdQOiMkJMC81C4qyPcY5N0TXN9BKcMLq
E9bv4C+DeNVBCpM0OgNceBQUBXwjby7shVoxredav6NNoShBt2puqDZVP3ka67BEjmKL/F8f9Sy7
ElnLiAMV3VKKwOOZrn2JuscLVwNGQDx1DOurKXBZmAmx7Av9gcvHRUTIZ7rYM67fO85nFVbtkPZV
C9G6deCay1Tfd3R6MVdV27dnPALphedxXITrvLYTf1QrVarO9gMuBbow+vVh5UIzYK4IG7pD9/Pw
DAtpOJq9YPj/Wx964AsL3a7fFoHrQYT3D2kHWQ5qoV/ig9bOigw1/yjwRJQIUhUhbfrxqWtw48Go
zPsrFb19KDrrai/TvFQ4eYoW8XRWlvS0bQ9HxWo3/tPo1W0Q4UOcbV9PXUKOW6oApjDFBtYnbBjY
8EbixFgjuS6mDLOpydEwgPUN0OGYeMRrsQ4o4+3E7H60eXanyURRbTjQxPl2Y5DZQW91OwqaAvyl
oYVNrQqjfLk+rqgs4arx7ukDI3SEkAZWf17sF5SBxA+FEnt7K0kdlsIxqSjk1mIsxg+fdcB+RbfT
nwLYPEtZlbJR5ZZybIrG3v2MJaoEIhahW6+xWBvZKSpTZEUZ8GyGTi63NjLF+Kzep3npVADz0x3z
ez2MIuumiKXZTbCju/GhsoQbxSkQFrtbXyTYC8cPn1fS/auujLQlBGs3sIUWIXYrW4/ww4a8L2f6
k1seMCKdKRWdWUBkfIWOacEVSs0cyMvi1azMxiDUbtUyrzFS8MPibwvc3OXwh8V7Z8aNwvXn8/IT
UmvHaoAa/+vs87mu7THA5PAE3yEh0F8A7FEKo55f2eXWHUngRZg4XQWwY9mz5ZBFUmXYVzZxnCh4
Jr4rRWTO8g+CEF5SByN0SMLyHArEs3ApGO8h7bWR0UuJMy9cSgZlxsjFJFUz2csuamLkbtjALJkb
EBqou3tXEYpxcmm+q3tTAsjhXp/e0pl7SwbeXEMZusi68jpW8inhy1U3V9aW5EmT6Ed5Xj/2EmnV
bWc/zbSXLXdtuS9p1Em+fyAhQUDeK7x4BN8sEHONmzOEiZx/9ycp4PkTZtJpkP33Dm1r3hM0wj+a
vtXaJfiaTIKts5aUk/aU/QvTITd1BjvPPH4/8RIKtJjKAmQNohQfvVks6uyH+SZsCoe4K8onKKmc
BPOvaxKBNvgepSKgqFP9Th+as3ve58UI/zbgtERROl0WfVtjoq9Zw6m1zIjKl9vmNrNSx2JvZ901
2EqpYl2xL5iPu27SLbB5wYNhK0nKysV5+h1hNmwpsCh64Wacz0JYn8Ao4wRfAQvFMf9yOhQq+Ex/
nSHJUPS7QAhGZ0BMBmxUISvdC/r3bP5IZ+dQ+hh2RRI89lLjsl/Cn0eI/+2BLOk/wsWPprAJx27S
VxDdfGzeZ9cLNaSBc7VSTaNizi+JI7/285U9sn0yutrroauKo/Mc3FQ5GA05UM0E5kUnsXDSplSE
7N4Z3GxERVzV2NmfLBSQJY0WDIZsCald2bN4jaY4XSHBcHrp2MQfOKkpHe5YaFYCXfXab0DkTPlm
/vX2FgZ27uvIyO5dTil/sxEQtq3+hzA7/8tguo5LbwtH9QGv8pL1Ny+G1Fw5HPbbec24Bqq42dL9
Usp1bo6pYArnP2CKKgi/E+mr4lrPJfw8blbJSZFbbALBKgyTx34r9L1IbqDV85dh2xvUg0/i1u76
BiAbm8W2o8gDQou4TbttP8rVFQpNktLUK1ITxn0Rjm/8xx5msnwJ3waTBXZj2d0JiQCL44IktXOZ
haydiCccjfFKlpWA3ZHgqXJ4+CDKJzzrMzDW5f19yexIApdi8OU88yPhwn+1PZzlJMwJ9cDttPXH
dde00u24q+T8NEG7eoPcwNEcePk7G33ojz2Sr5shQHm8bGHhpsVSJOllg4sp+fqMX9B1S/PrV1Ed
WBbF6gso/EyDHur4xQPkpXruxRQXHOUsIacwCuOc9BS7KmFcdRnNyiLmdqmoMaajLlrRieThn5pT
3eeNvZuKJ2997VC6j+qNwKh7x37UQuAtd2Xk4VsOzNQvz7awM3g7qKVDyilKqmwJdunoPHsUCu5l
KkUT1KSxFVSTCBfPr72rJ62qILlbkv8fJRqOef9+U3CAoS44LZ6U72mI33p/NyAShksi/+559vRq
SEYnhXCkSUnXR8pPrkhKMGoHR88FMt14FPDasOh6p2ywQO1pWF0wC36hic1WSFeIYAVaAcHb07jM
BfNktVBEpdVIuI0UcU2CdBfyxwy0I5tL3bDSCFjUgAu+IMct4tlGPAwGRY9mQj2N0iUlC90SP0wK
NE7XmTotM7vm3g/nKFTxKI7+tppIyXFjJqDlPcmKyBtgWXDaTwsyEKsee2B1DuJtnYWZjpfxbg5V
kzSD89zIPUZn239zSmygi/DyuzHeLgmS0WKzkC3ep4gwNwBMdKQds/uwgU1yFnu3OBANZbjkMlM/
Bu87ujzzRtT7cZRzCsISw6+KduZi/FzE0KTZNhjeXeHoU296LTP07SkSGB9ggjtA1tSVJu8d8CRc
7E9szM2LFkqq0z98NmFEPEnSug2sKDYVRAzAmwbHsotw45sirFDOBSj2pb53L3PwJMH8A7SWeYj8
n68YjKiTNfdkL0xOhA4TW6JY2zE/sYSycM9DLtldaABC1EihUdR9dPxgIFsuBWhAaryelxS4995Z
4XgjkLitL35y4kBbYi1gS+GIyMvZsEXenPp2AXF0hPP7+72ha2L5arhuXKcdpUnYdYapS9eVAWkT
IQRmtGQcLcWve5QUzNaSSY5W4+MNIp+IqXPJMBBf+px6BtqDFqXOkDYURxvqsTfiddquaZsiX+ZH
zoigdz0aSm0f2Ku6zU8Xt03NENR8dwN2A9zYR1WQ0aQjj8EYOWVj6qF8Y67X7l18eB1jtE8LTZk7
PU3nCEoxz38vpiJZm6rxpRefgxoWAQYnNZObvA6CXTK2vOCQ7urMGnicb5HDLBz0jbqRdBrUP6rf
xVc53H5KGPKgwDcxzRLS+iDN3I39a2LNEwDCRwaYRw7oeC5TDoJzLDHJzdCboUb/ok0BulznzQ+f
ljHt8VDKe8+fba5RrEjhxE4mvKy1R3p2ICSYoa9ns4EyOtAz7wzogDDQoL8LqxIo83OI6JShMONS
GLQYhJ++HFzsO4L0CL5PkLbtDOonuWmOdnGCAksnZgvzGQAMXxlmta2ik2jC+BLC42kLgiZqpUk8
K1wJ/GIPilFqcjnvIjtYOb7CHDI0Xo4Rp8mzO5r5ra9IezEmq8g5G9lRQ+Mz/pZnMmOX3d+XtLOK
ShT4C6710nVU5O7mTASmLEKsR8ZVgWSM+MlymdQ9ZmyEzhfSrZxGmN5H4zH9USNsWEVDgI62HHzp
H6vqDaDlMl+rZ1SBvElhyS0xbqnzmQjWVymk0GGHovRzRUHFWpV+7KepcLxuVnWPg8FsX0z3ovk4
/GtpjR1hCZ3+W851Q0EqEkSHHbe0qNgotIq+MBWeqSkeoLyzQqrQKkpe28dK8TUzmW5WnrShlyt0
mVF8IyyEULimshXtmWpVoyX1ALCCQ80UnVTN45phq5nRkFB8GQcUpdM2h4CjmgWTQ01LA2frF0Vk
G+qRm2F1r2AmKTml1H9xwm6S2dvzphGR+RsPI2oXljaLhyQpWsK1xzorwnm9Q/O/12NuKmr0ta0w
V5lmtngkV2eJOiycXCzRNaEG8tVYFTKP1Z2NJSW4rOxJUwnkUcyStqIpCEYMPeCX92ef+uUI84Ow
Gj0NgxNJqXabmWGk39zv0WzrqoHVideS5ObPIs1XOFuefgzk0G5HqRduJRlQFHnlQds+eCRcdisn
sHkLPI81xcoqTBUBw+iJVOF4qX/zcQNeGia34ro6A+sgu/ehimcqae89isoMmTwlCAo2qPkCWGV9
0LQpPNnvgAwEr4gFizKJtH8VVowl6m2cocGqMmHWajJS2jsWTs3JzfKX65B1u+4wrSCW/ahpfy3Q
6MnsOTp2i1cFWng1qpTxpiOiz6mabYEMq/C1w4C4qOO0d4gh6jHaEJSgYyBKM39hvljNQvxIzvW4
26LhxxJ5IwvQTwXozN/7qGCTuekDaUq470jB4cb/V1SisFJbCEG1bFu5SQTJZo70RGRRdYEB+PkL
Y61wTvSBI1KzL09O5nOPnwf51l6RgKvOY/ySSYgMREBYX5vM+1edMQ4NoIeo1Vi5CZgGLkEFgN8v
Ym82pqsOx1kxBJnIBPidMckXGL2tRwa9yGswHPR/E1XMFU2+1rKcRx7yPhEkY6tHJzlPYoRh1Oem
4RV5/X29o2I6AJUnGHVboeA8av+dbEup4Q2Cu9okW241zcEFUobdLHDY7aZggXYFQCKaKMy9mf5M
NBHTTVWpl/RYBPSXWqh+DF1+59N9c8Ltbg8feEhfb7s56t3rawyoCTYLxfrkXZ28NSGEtZCLobz9
zHku0KO6PtmMZq8gPX9YWaSaPrKB+ywt6bjbWDS9njlO0nNNXkHQv9MpeOMebj97cph+nCYBY0oV
KEZE7T+S1G2r7HX1me84HOE3Jndi/6P0sFS4YkFGIksTrVl8f98LXVurHJbytIzQPqxC/lM25dGE
JJf2EX1cpb5OY8zDUugCmxcH/xcMI5RjiOW4f3LxQLhm44XZNnbRQRFkZIgZahxTHAUrY5Kzn+vB
lR8dPwKYaRbqhRg5HGFm0AdUqRevRbsE/cciANZs455M3cD0w6T6cSyR5a+dBpqfWwcOqqgkpVED
N66p3EVG53/s0wW5aUJnEpctdO2M9JWjUcgGQTx0TvNkupwvQ4ixkP4ZsFSaSXht8zoHJcFe+h5M
fNuA1I8F40frJcmW+8OSoZC0n+PPgK5Vv1JPG2wQhRit64ZxIHzPtwe/8mX4r8TBUzH1T/RX62DA
uB2BSM2oi1pGhHhE6ZFfjKmYs8bVgMQxtmjqTwG6vj2j6DCqm5k2Vs0l1l30j5xKZvDm7D8PXGM/
TgPdhSgaCatsZciSnOax6BCMadLYQfmO9+5DM+IEv8yFDd18s9/U91j6JZT3QhjA3BgUluajehQo
10epHkxSc/B1UoBx7gWx/OzHtV0rk+iH2ztxlGadkKViRXzse4YUXVueKzZ8fmkFThyYBaur5xAJ
1GOUpeaQfswgKc7Ooy/KXndmFmlU2K1nHF5nZ25A91PCTt5Ne56qX855ZG7JKMtn/s3cx5wshANR
Blu5kLM7EI5SnF1vOAKaXYb1fjC4uddLyawqAgBNh74wvak1eL6oEdr5EI0owY0b63D8gGDco7ps
mcUIQJkxjsda0AGrB1Aq7sT57Z//2gIdKWZrGnGgt32un3/zgA4O0AEtv4ZZxHiWtv1Lm/siG+aF
1EqU9ahGgT8jP63aE7otw5px1cxD+JCSmKTHxPehgK3hznks8pb9S4mZtYU9WKJphTmuT1+rKpDp
P4AQ0vePiXCVyzLur04oU/vtDOOEb3K58dQuLoFbcGVKVPhwi6i9LoQJgs+6pqFNQVGvlL1zHkJD
42yCMHQhaChpAtNjlhY3bIWNH4mH2KEQxdkfqS1nQZM+XGBdtFgTnBIbqtpEISwtKxuMc0cNYPwT
EimKQkb1E6aAjc1Huiss7zUHLx7+Rjha5kQARizGwORhhePYv2fUrwlufc6uem4RAw9lS9ePfgb4
1Ul2t44x1XnI+UvaCS3HYXS09KnHUzE/daisDJAu/EM/L3nyzugSVtJfikp8P7wztT4c//Kmzxok
K39pmYUWF/SQ5TnIFmag8rGd0nYoh3oSE1oUpNyoDCV3aRnJ6JALy1+pSoeXpY/rqVkW2gP7tg9M
GkIqAu6aMNchw2hlDZQwy76ZlqCRLG/dZ6abgyIk+atr2jU76asjk6FRDGbYsAE79boOLCaQ7fEZ
4ZzbcvhXU+8Cl1Il0JquhtljaBHYum9ES3HCWWK7S2/uGG+37+yUGyrJI50yvhCKEX79sK5DlzS2
d9yCJELwgj3vw6xBEQXjv3Vw8rxkINMpBdWqZgpCuDRojMdqnKtNw4+tMNrU2ISUjVDstsIoGNnM
nQiH1VVWzIK46Aoouds=
`protect end_protected
