`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
mZKCjVKZ/OqvnR17vn3ZI2yfTBRXnqZvkUG5MgAVxnKxOsRNswO2kWeRHMnLzPFxlLzzY+ydnoJZ
H+LWE/VNrs28Mx3JsHlhL+3lvFSsTXF16YRgJfq0Bpd/7nFzHzX9KpYzWauHW4dPitlv9M1goQye
A++VkwTYD3sdumAr8cG/tycXhuh4MMguqq8WBLZ1xmRJyv0Es4g+PUJVumpqBVlX6jiEeSuY13/O
QPiFa9n8xZqbN6hO+k3dQ3n6fDomY28hx983BMvLaDQsyQjH2CLAt8dDMg1iy9iEhosysS+976z6
R0d7cHGP7G77c28TQBb3J6m41dfqDPywE4XUlg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="urdjMkJ3rDDszpJsCIbJmOq7NX2JUw0L9yutSIIeGp0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 205840)
`protect data_block
jmYC76ga9uSw/f1hk0JzcQBP4v/C9n5j1/XMOw8ARyrImJJXRtipoShhjuXfo3b8gT1av2qq7Wyx
kRFsFuePptk/QyjTajgHfVnuDJpjPIbgSsxmvSub5rFAWijke/xfaxSpuvcXDjaOWsXP3GIRVvQK
HHjRoqPEWSc6fod3tlsAwAA69a7cLc4YoBJz01oiZB1ZNJbprZZDj4X6U4qmdSM279/vrr0tvEOo
bblVq+m78W+PgUrFbllu8yJv+lRbT9F1tkSWKhcjS27Af9ais0HYMZjVoyh2PUY1zG3W4pEgfm68
GCAf4FA7DMKajM2upUkJ3sL12IpMN8wwfLQiw7776os+eaXyecPRkATdzMXKZGBZcgcXzXTl/MXh
TU+eCF8MO6ZuglO+i2DHk66yUbmAt8UKFJKNXIbtgY4voapqU4DvMIo0SlfLOcMIP5vB5O3s2W8h
Ce1/gNtgBj9r1qdf8xq14beddW1oZ9rGqeczYI2h7OV/FK7sk2/SzRDwqSAIGO6APhymwjuPphw7
otRRESPhoEPq/7JK74JGBU09QPWnCRtMozwALPMk3pV7e4jcB6rTGFWnfzJHTaEITYE0MCiytGy9
Qq4pji2f/FT7lqOTTCOk5uqNXdOXmfA4VQBjh2MnzXtQ8z8OFSfMHIVoGUaJcirvHZdqV6W+gm8P
/V/0HUmRhZdhxNiz6gTcnVVSuCKLdwuSRZRyNFmpeVo7AHzwbn75TJTSETllIT051syba7H4++lp
krIA8e38jYMd36jO9wpYIw5PSVpf8gcADWpXkJSuxckM8Pt+qW9gI39wh5yVjLKVo7t7kU2U8uHF
YT3zItmRlN0VY8WiVLtY6lG0HEI7+BMduya21ShBb7kczANOJmfy4RUGvJqNeQNlkpQoSD//te6F
6OchjumVED+Zm4DO2KjNtA3ZMlGWHMC0VnLCPg2Kx7T9CqWdj3tgtmQ45r+T61MPKMYmHgVBhE6v
MyEWQnooJ2glGauNEw30d3dDipbyFbiOx57/KdnukBC/21+J5J9mvS9nG+5H08k8XPJ/DrtZvso/
n4PaGPO4JvvdE0xOFnGpEhx5lrk4LsoDpGPQqAu3nY9o44xff8Z+UmcniICOhyxaAOecuWppERd3
sPAaBPKZr6uM1Q0zcU/8uy1zXbfP4PNmHnA4AnanZ9DaSgEBQ9T5KoKLYIK/o9CMk97010MNj4LF
yTFMQzy4iPSoFVJBymP+7dY2Be0mKm/Rp+V8cRnQEcW2qzAPzcIRlcT7yofbL0WzuYt/CgJqC/BM
PFAkbtbElFazNhyaFOQkUG40KgNeggD0ydbIjVLlcsVDDZe/mntrDIeR+aOIsYKDK9o38AiXNJmc
DkAGkJODqknCaQOtCdQpu2oG/dvQ2HS5rAcTHysUComXB2zFJIEIdgKBOYGxP4sjCA3ugSwTwwsf
rfuVjexPPrCvlGMn6szqelNo2cfwLy1v+3W/6WRRd04vKjQPrubIMFIZLrMpE//z22PUJAALzdX6
lLF8hceuoemEScYO85qnKCDyWFiv7jstuDcGHBVUo/8rH6zbDryfkmYYPjct88B1G+urI7VxE8JG
9wy/LTp3AGhnJNvPw9BvpCAilPokFM0PG9104F46GONhnWw0An144msDrnoSQQL3pzEyQ+LTvRcR
7XTsHZvQ+vAsI3TtMgXT3VMC5C7tIeSa3DBwb6wg2OT9fhlRMnMOrUM77AVHwG7Ybd90EhztgQ9d
u6Ci2pfLSeLnBk1saMDMquvJtuVtWImL4zG1ggvFb0FiUXZHq6kXa/fu8/y0qgSa6aUNJbBNVB3/
2BnsEXc2gHjSogZ/PsGH1uREOFrJl0R93IsD4pVX43E3NL0L+IihzUTocJRysUnCR3aP05EQmtlU
hC1YGb7r2SvIRUbLAgvwX+5L3PNnVvlNzM/Y6I7P8NcFcm8V40MosohZX9iNV81C/fv64x5NOZwC
WSO6dGmvkqWQEycOnfDDi4d7vAIR2f80mBKzDLiD/gsuFUuPDsjEEIRjN3pGik23qXzcQa9n+bve
2jnguWavPa+uwb5E8nMpZ7Oyk5LcrsTBj9qUd8LmhF+PCHyC8DQoL1BXZu4H6RgcuNZXvfmdQsqr
jwYjF7YcH+64IjOi+H60qml3bhv44ad8cJIEKb8JlDW/6cqfpe1QvOjd6q+BibsY5tPPSpPWl8mr
IWFoozeRlcZbopUnVybEhgqTi37dxdA1o+J34pUj0vEvuRHdj1nG2CqKM4wp70tF9+ZrgOWTuj6U
ewye+VgYPUBXcZJuEVMoa6Rz3r4ALA5mSAJhRGC4d1YgXqBa5vAPV++vNh3TFrOJnIDHfykpDuVB
CXwR/yYRBt8xV23u7QExZ2ggw1zeFB7v78gyJh0x3PSOgTj5smRYq7fcx3DsH2KfjM4V9XgUseta
GQl1fqt5L9iXdRSeQGlOd3tOQU49vksbaX9Y0SiMShjtNI1Jkbp8jzmztZl5Rl5ENvjUgi/8Jltx
LnocankRGzNKinUS9e70CZAVwlQPWVqIKimBTh8CGBl4YEiuxHzkzrymL0IB3u/l74LyqSDwmUQV
EiVW38ND3rvelts+QkFWY01hGAx6Ke/zbMHXzqwqNN+JSbihFq1KQZG5D72PgSl+o9XZ8mUEwNtO
YvtSK8HYN5DMvpE/Wbmfkchfc4+st0PDqg1WsoOeDfLugn9C1UuXTJR3zyJvHgSKntFc0I8sNYRS
CuAAuLTRW1APu3S2xViGwzHSB8rY3HRsrnn7Ul6VTy/W/ziwHwvJAiAhWsc+azzzDg3iv+zXlIro
WPJkjqBO7kp2KaTIhMZFEa8RlFB8tFTzQhz5w9bKkutAxbOt317bv7c7e4XeF/biSfOBZygPMiZ3
rZ039g7AUd/zWk2MKXFQHxs8ZsVC5Qd7BinFPA6SSHgEUIU7hzCZQ/bdlzDQyTsAt7rPn3D/q7bk
cxKgJKae+NCbjl/SPqxiYlJ1lnx4DVPsRlgRMZ+eXSHR51v14p9mUw7hXLbgfZlRkDE7wTgGDOxq
py/ie3RcM0akyrc2Sa4QAjuan+6cFPicYQXMTo3Vvna3D6d+X3UkF/e17uKHIlIIYF2LDarWmg+6
MF2PSJJ1r03JS7H3H/6F1PMJ16tEdI+e37a1ldhPrnixWF09FA9ZYg3VDnvYGsCz7UnIdEQYeiVe
sG27Io+1JX/89dAZIh5wfDp/OkkWXeYf56PEtKJOgYoZxfF5H6kgj2NGRkhvRKRKQDxPZzebvm4j
6/T3KS+e1LA8naOP9odZ3veacBf930KM3dX1e8rMBvqdinE90YLz1f3x18DqXLrpvg0atuLetsIb
pyh6E6+uo5MYrltmCYPbOdG3E5XaZ2s9l5EKyLE2JOR6yFFzUqTW7XDiVNhp+zS79yxmLHam3D5O
WuRUEOlpno+HV4EuCG/ebqhPksC2fzvHgm4udSnFXHjttbwfGrqsvfkparTffJBsVwpfbe6CEpWc
DVTy1P3M7+icJVyqs57ydIrgDoLWwmfbdvyVJ+YQRlgY5SX6R0ryiihqRazcktyqnvleTmqe8pco
z+SK1d7Xitsy7yBPxnYTNPr2QMLkKlsWQLjDyGSstImGqvg1qQ4MNNKR9MlycwiK3vYjaaEeq+yx
CE7gdiOKKY5TIORY8hkU8mlOrY89QEpgVqq0IG4FGdXjqxSyGAxpAQPD52HhO0vopUHjKDbbllK8
q3rRHuTAA3QhaTV0qXXsGafZU6wCGP7PX5I6IGJCzkXhSOFO+Es7f/sSl8v/Cbu0/dQU3nN01UDJ
6chcpVPEfk8TY/NXHxAp7HCpvGG83vRpxDqf2G8Ia/y2S9ixOSIDH0rvsq2VuJCptsbJ/WgqiIQn
pjWtMBnkRPK9oIochuCuVwmj1ypPvSxihMIR4gPtpFWXmgTN4ONF7RYRdzORV9F1CJVrpPdgFKRh
U4wziLfj0fCOv/vhOO5/Zzc2DevO0ybGCBuhgUqCT92ew3W4trLDPIYC5CM6+b5qTDeQhB9dAORN
dPmcPABwHlzHZ67b6J0twtXRQDsESSk4gr9HJMeZI0i5dcaiekr8nv1o6X8vHJsunETywK963RPp
PZN9x4YXXT6uW/pIt3ltE1CkLpw6FPwnegQtBP+GXbOzBXARPhQRLDr9BFo3LWog6i5IbhU+VqpQ
BEUvl0IsHs2KDeNtlvyK9qVBKbDRlybisvcKJh1DUGkfuWzw8KwmV0Yo7XGwZZG0I4FRi7AV+zHI
pdm9BCqqVmdxcsFKqg8rnNcH5zmCs8WDV0dCJ4U7RDN34Y1IlYS8FVGXfs2Cs3IKmvDOntWe3Wqt
vmkbH5vlgRXhke3tAJAHh5qmQzQMbQ8UXrFKIfDy7RV3uPejdDuiGPBzhKH8fg416r1t4LPga9KK
FkMxmafaerfx6AazuXF0HWXT0g6EvM9zeyVdE2x8mLcVHYn6gF5Jh7cZmGk0wgy51EmoqQo8ZtTt
RKHA6GshrAaEn2bBgKuabl0IQ+C6Vi1nCOTeqUe5Mlb3TgdkYXGnva3aT61FqMZtc03BXIwsEBax
2gXfKlg++OCRUeLgbrt132Sld/POX1LSsv+5GJBAY532nPFwLMEBsuw3W0LKL9oWLHLCRlb7pFqj
SQjUndHUXg1nxXtzxCmozy1laNgkT3wGYDgZyIeE0X7HW8cl0NSIfdzVzm8cL5TT6OBauXljTHsi
b8TG/A5xM+YAL1VATEMJK9SqkuP8Hf34Ui41KV35oBLEaucOd/+cms6fiy/C43DnwUHgYBBz2ur1
DUQDsvxQ1aAYUc430QsGgxEOFIFkYdJ++JQfhKlONy2OJUrGgo9BXvZ4ZaB2Pv+d3g+FsVlGBNJ0
mLYSH7DiGtZcD4xL4TFquoIpXANLIRgNObq5PQdS7ZZTy/Z1f+IMRJQp69c8RMF76y+NMA0Mwadi
jxUwrzXdUKOtHOgIKTSm9ATGHruMt1lMJ+q/8UDB3fNmLLvNiE9mq2e94SXb2YznFCEkUChKXoxZ
EV6vDDhRJGAJ8QW2tqa8sh1Jz3p7zosHxCqm9Umpyw/Pn7654ctuvz9MiiSH9VWDJQ6UmryByYTV
ARxCOic4PX37mx0KSLRrlGTxxkI7YuLkU8Qf89w5QJ7qmCLP2IU4VWYiLw8PN95jIDn97ZXxqfDa
hEFi4rQzjoI4LpBDEvqnT2V0foYD+jnlUvy1OKaEZxkiD7w4d59iViQsBcEgl+9WqnAMo9vUXdWE
sZXlYbYm4fS4rM+Yhoz0W1K9TV3nK94brREgHPl0HIK4pZy5rb05gPpG3L/vBOmn8u00cmmXcKqr
05FIZHdiU7fvcwNbH1qEbNx3IX+QIhyQ2Xkxg23OIbnStaAOjWuMGGBiZfvlRrBQGzjse/+H59qI
q744VwkRaa+tkVfSgvNy4USDvs/XMPEMRngZmhuv70uGT7lvUd2HXentQLHx8AuDQhRhYkF3lm1E
Yqq/3YgSpTDKXQn2BJE39bflADsKyCjhhqbVqISfvef06E5kqAQM7VYiMatwnUMc8C7eU2pICYvB
JvygekyXEgzxSvv6HnpDd6hOmZ+CH/RP6XbLN9/QJxKAM27E58/gKHUsTG4IWVnjMZP2SWGjGbha
U/5Lyyb9zsF5GLhI9bjTdSOLfWt/9I3uxcJuYxzTL0Ppl/ysfyj3haET/kxrNeiErAJF/nRtfd1P
qPXaqamnPp/S2Lk/SNdhxTrpbOvZlrEABcXIWKg7aAHp3tdgvPfiiCSbvl6+MuK8eefTlx9Blusa
rqNwd7pHz04TIdvxSINkqsvtTxnaGD45+vaNteHafItrv1fC9a2ukIi8LiCfmFME9lNgmGRDKeud
vxxPlg4g0waTMjZoCLrquBSWaCRHAlGFdxqGI/z9qWl3Sn99A6cbZ/pvYYWbZ6DKJyQh6TvAg8NE
cSUjs9zUusd7os3tgm+BSnp+l5MGk+cE1eh2x8DlF0yTOu7GBksRkHQBbPYg2mzQdhXgq1UCcA87
shdKOXG1/so2v7u61ut1g5kRt3lL6e2EQoRWZhhAo9C2e7IOrAwCTz3jkgW8KGBYDKxVL+SAZJS9
6kSGAvd0bboI0eIZNv2FIWwTeNdMfOJ2QbM12/Jagt2A0BeAlDGRwJDL+aTkqAuA/pdvjbIz67Qo
6jiQPmttAqS2IWBuuXXccWKN/Mu5P00Dx1O2Nsy6sPMDSyWVlAkgwnjh/34AI/LwXSrhkIfrA3QZ
qd4ajTVA4u4pcJivjdoR97Bbuen4zXFfX53L/0G1SpsdlYq6e7g6kcVTP2dLepweCEOW3VW/rZLm
Zop0U11bSAW24Dk9i7bF1B1SJFOusuucHjhgLwSz/Dw7M5dhXMYIQh5fiSMIsqFIwu1baR52JC68
+zXtcrSmPCV8bNTAZ8t+/OJz2d0NMFtOTUd/kULc/DpQQ/Wj/pY4u/U11Crscj9R16xIWCOujRSq
LY4IBeEFzmnZd1t2EElAtmo8uvZtKVHOMGdu0OZ3cBGxlYCoO0TWq93gGW+vCzOfx/KUU4tN5S1D
U5MWuMgz2gDi09VF5pNspBl7FF+h9rDIfJ4U32T/IfAlDg0LHGTWexBVvTBtD6balw6GJUJPdlXp
LCTFE+uYtVJIjhjMhA4V7GzUqlRGpWasiQ2YXMg8mvesKKmDf57HkBFPCKNvo8BHSGkr5xla9k1M
VU9xWQ75zN/vFfEkJ0bQXe43TwDm36MSRNI3s07T9Vpd/qDjHSh6A3jZr/eEnJkDtXaEk2N9mV2I
ku9l9b/VQrsKTDr94yuyXLrY1IqOEjLW3A4EvKwHdmGHXHoISsLXzzqbwX5snkcxPF/kT4alg6Rx
8ESFcLJKR6tudm9GedPky1N0P1NAOe+THdg11tMWYM+2JANp04lKCRAajaTAC8/PY8wYJyu+PDXZ
t0CyyoAldLoqomiy2gZxqn1OdfQwHypr9v888PxTb3XQoskhW/gxXv+bzxNFx/ehIHuKc2szL8GK
Xs2duP1fayZKiYsJH5lsPLfuJ4UMEcm5RS8uNWqH3rWriZpSN8axyUWxL4SyKor3K1ZFbM37he9u
ZmfRuvpE0CK7sTQGsQ0kWURUDBLVyJRoS0m/2hNtEyVdIi2oF/9S97hjRxrOAZ5gxXV9ZWUI4hnr
GpJjIBbfaX0AVS7b1mu3zj4Awjzdavd1t0fcj2UxO8BDmVb0ebP5B1IEEx5KNHXNrh0velbRybbg
5O5wAx2XSe0KnPavsjY3C1ULXsMWB8jw1BEk/n+Fzks0pgLz3SGq9fzfl/EIs6eVN3Jm+vpQBlA3
1GcjcQxgFgp47K34uBjyTkU9xVyDLGQDQnFhdmPxdPQF7rEZldAYo2yAQj6390XBPhcX4XhLcF51
SWfr4BVf3os6UAqMNBIx1/it+MWSpiz0yfThFzZ3zNMM1C2yffZ4SY2jLiEfWuZ7bdIo3zK5olgc
7z5+8QYBwU1a8dkRIL0WKDxrYuQoHoORw8ao627tty4vxM8io+WezhUZAziI20Egb0WM6fphMDy6
Yo6KWRth6/N5xD7pddoSwTKCg69pov+IEyhhwjt/p4ymaljZ9bifywKiLYeW2f9jkpvEbz9TchfI
YUfn4wXtTx5DWtQ+QDEYROpG0vWOZzIjuppTjjqXY4D6Q14i1GiiL9qWQ6i8i2L73zefLMeAj6SQ
5vUbYBLIkLYkBLWC8TXL7HS/i9u6d9EBzgMC4k34ZWP8/UcQt6F38TicuQXQsrb+qqEORi1N79qW
7WFJ0IPv18PqNJAol0vw2Dlh5YWSuKfWCmaNxDD7FmIyvgA1M0VgPJ0dgV5iRhuSF5S0loQUqHUY
KJzNoun10Q2U5a9OloW5eRegqLMo7zzM58PVdxJ05WjeK3XbUF8DgSdETv96CY8rL3rnVU8bm24Y
03gRxxmXO88NsOngSuOmQAgGmAYFYaGu2rHAReKammjge+mmQVzA8V56AtYZv5cWRmnd1qEycMJU
1SLiPsELq/iXyjbDukbT9tpGucI34dy3oNyGB2y0ZeZ3Og8Z1wk7WSS3vpDYCCAA12fF5LmgMJ0m
MTv8j5xdA9oy4xaQOcQ89HebQjT6Sow56pHuoXMBL5Aik0mPJzwV/K0LSJjBtlpkQR7HBNARPycl
eqxP+AayYfT3Z+U1v//xy6Or7y3rbqLzcgFIaTZGOI3G6zhLzXiTne0RhMevcwQHYyJPNxe6vvCN
2PV/SwfMAFInU6VcdynMOtu5yzG3mZ4nMC2NElWvz4vp1UG0EFkq0r0T0XE4pyDtXBcP8hWUnXGS
iqduUWflF7RBe9uluFL8iTAdgqcReJNAafpRtBR3lSQnt1Th+7y5lpQNDoLzlW6m8VPz/B3j9sZW
tvHu/97HZjjnWeMY49Qsdu7D/LXj+mpJI0IJQ59NXO0VtQYoA8JHv7F3V1vNq3FkAJGhRQyyd5Hv
53XocwQVJhNfKpbEfOwtCS8mBY6mkjDGBLCRsyA4HmqZTZhXCm61T6RF84soWmNDNYghu+Y9Co1R
6csS7pz6vwu6wG7idpKs27afPdQSTvBRGJwHQxoRVOsfncNMcY8FbgsMRQqx7UfD2W9UXtn0/MtX
tcLswB3gsNyKoVNQik3bmr32vnkAaEPXBzzyeqtE9iBZ5oNJFj3weY6gVemwULpn+8nm1Bccw5kf
1vM+Erb3dQkEt2JO4U9pjIDpkdURrrC9/opzhRaanM+cK0WN3eiBkjaUxqOAGArNpTFzaV/6sjVU
rMZPVHVxBFqcRdxZ5sCo64F+dMOVFtKi5v1rVE+LSjp9ZpfGr0gBVoiH9pxQeAyVi4gi/nqSoj2R
Kxe5UYRz//tN6ec87wOhOFfm8NuZ/6MTBE6u0smfT/mdh3GkuJXoWikDly1OUjJSu+/10OVJxnqA
o1wGUBReD5Yqdoz3bBZtimRs11A0X2xTBTnCAHjMRg5OOIzqTlW9RsZA+gMSJdmFahf/nL0UIvBx
4yxuSccSnXpeZBqHoBGiyaoCnzOz3OqQ/r/8XxzJ+7pgJuDGNZI7BZ/hJ0QsQ/VW/p1a5GMkOsgR
IOGpsIjJW5syrgLvcjrSY623F3T1EZBw/tmgCsKPFpUlMHyonz+sLR0umFDFjoO/8thCrLjeCEJl
Hm6mh/eFv4x3oPDa0sW3Cj/Jq6nLC6+pAC3dCagey7Q9pYIHnpcZc4sbWJhUfTsGfcZPWc+4dv2c
FzBaxI/TGnNoJc5C2E0wzWIe1EkabImpwWxtSWUbruJ0asvHEzWYT4d7jnq8p+ATQoX7TubjUUSy
NvS1j+umdQuVNP4kY33aKsXOJSSQEKLbS548+mUPn+aRbMm2zIHchQgSew13Yi6/cPZ3aa68ixNU
u6uJKW3Q5ASWEmcfKjaS7APyeoCQqvHeFpg3IpJpSWc3nC85DiQShzAXsRRphgvt01waJssxHVz+
pRPhSiQkYSGVO2a7IFCPFThbyL42YC4i1ZhEuClM8BeOOHgm/X8F8zV0kDPFCOi9sjRJByOVCXwJ
1tP17s6BG6yV9HQYkZdXjiCQr3fLK9U47gOYiEXueOyCkW/qZqlh7AULiukhpOLk3UgfMFZNfXi1
7FHHHkL+uEYxyag5qrGbYcxXh8i5df/0u9QWyr9lI7jXI3v2Fms2jO/n6G5vlKIVt4gSzWiJlblx
QY138cv60WBIwE7MiOsqGcVrs+507GijIdlwfPFUiluAuiDeGtlKlMB6Aqdyf2rBlz5G/kC1loEb
OZ59hbx6utd+5avpOmJu7z6wPrhjgU7Cs0WlOzNztKpADsdRYfkSxqAURg4LgcheO88rv83d9UIN
VVzu1HGygoes9TzT4TsahpijT4gR/FUZlNlvZNeWtrBpRk0IlwqwXnThMAll6F/J6S7mhq3SBo1d
zimWC0lUoBCi1oXB+7ifo1ntw2RX6G7fCDdwAUA3s4YCeIPlgRl9FMSYBZ3bK4Qd0esviLalI5RJ
bELPTSAOSZ6sPKv34EnA8lVoyNV7tzCH9fGDuFZbYIJFv+z17cgfKrd4U6ci1pe3Ebh5rE364Dzx
xO+YXvZvlY1cp8FMBYPFbIZuAOrwbq+5dN48yXC7mVGrCzYYUF4vqkzJffYyBaVYW4WsiWZ0+ySO
zfs2TSYFc3iKmfzn8p6jnIDggjtOw+8qB/TM2v55BKgNnOM0TDOYQhueTzfxuHOKJLo5VBuDNPXQ
KwlBeqOoYTr4jSBnTNzeq4iSzDiLSoTtAKLWbBG56HKZpnX1fvciwDzlKhTlSIjkBECwi9UAD0dQ
mgTBKw8Zoa/82PG3RsEEenQGFwKg2815Yg8U6wXVW/S7cJcIGx/mxcafWVhmIZllr+RnG/PoQvfn
7Af6sxN3iMXXo3zZz343S5ZeVTW4rF2uVmrPBMFXBvVhQIFG+SPR9S5QOMwUwZynPbCCLY9pRmUY
Thx/MaX2dPF6l/76geiwFCnNpLpjjkFBaYQUC7ln3kcRvZzaw+iGA/MnLzGbzt8GVF0x77c51+RS
gSG8KPNS29aCY8jiYlrfeW7UZ0Pcp+aoK47zGp6lwdCYTjUOjFTPdp3k+OBp0ZzIJD2I9Rwn8mId
OxRZyD6lQs7EAcjrzaqobo3kNJVNsjlfRLxN6LM0v/qhrji3IFeH2FwVFuallJTV5zc34O9k3a2I
eNhuu6ra3GNqZh8QgnsTZbn8boKeUTjzlzyO/qWs9ZGM7MFEwH1MHPOmkS6jpwOg5qFhyhl03hai
wmRqhXLCqGLGrQ9EtJjoqKFeKWmBw9SB9XgEv66eozkx/LP5laKynze8RBZpJZkWuz3Uq5P0Nh/L
u3ridzjcI4xNfY+orQYXLY45qFWWhGK02YZWHUfL2RguHti2kc2hPylpEOlDhvJGqS2jZF4PpBbQ
mScrW/+GLRiAosGvDxt2L7kPM+NFPyLKEcrK1RjgJplyJUOSZYNA+J7Ow5wDykuTBfFXXryMv3k/
9CMLCIZ5EWZdheD2SyybMCvSKYYNHI2f07zDubUT3R/ckk89phBS0GySn1orqJzp6PWzFF5IkOw8
3jwI7+Cc0qGKGwaVgohj8kkOS3VHq4HV0Xfl9fBZ83Rx/GqiTMX7eldKtIScQndJI8TX6YZwvCFk
2obIR+hSFNnrBlO3GNUplJu6MB0LmgBQ8Jsi5qtCSs/xpCADO/ps8dEP3qZh/C8eVRP9VKPOhtMW
7DkSj6y2EgPUwM0IOEMQ5tmJL9aexwZD3Or6lpyWAEQyiB7aT8zs+1mMB3tRoZxT3ZIIUBNWcQ+x
W78pyH8up6JTgl3b6mV4C2vX6eLxXuuRQgPRyG0Iv5DjnJ/C9HAIsb+U8BUWray3kFLuTMKMQ05L
3n3VVChCLdueDBawYzBblbzvpQpcMsAF0e/WYUfZQ3sAZGbkwJL68X8BpP2c1da94EPtDpJpe83B
ZxmkxbWnMcncp4LhItNlRdmPYPLDAtFs4OMC0Ml4r/COKVL83J8AfxWnwFqFnA92GbFFEnn6/7ps
Hyw90BEmGJDA8Q8C2opd4L8WxxEtvYR559kFhV2QKshtPq4O6RaFxFU4sbSlo0OteQd8bk6aaGP8
6ViefD2m876IiMJHvlTTo1Z76WQ1ealot9dUiMVlIKteyhZXY5q5OR/JwjXFiyo3t37KEiqJLNM0
qw0qsjaMmw9shEgm1JZZuWN/c9be5f4u7thYDRuUsyW+OZXF1pOlKVNAAAtNlySCT7xSoXi6ol9U
L0wt6DNVft2IPHiwlGi9lsuA0aqyB84ORJfW00NK84osPoQ4pqVEP6ey4s9s1UMd8J98U4/NI3iM
hzqk5OI1P5BgOpB+Tak/hsfBNMMB1Jr6pLmADlS0AhQdg1hEc34iqFXalN1TlAo5RUiuMQ80fbfU
SbsXzyAZ9d1dIqkVVFDkFoTgIGemoIwXjHMZXza70BWKqv1lCZzkuk3P+HfRKVAIIdnt/5IOlPTz
J1Kx4BJ1Fzcohre48UpGM8ZnxAMcEMREQ3CSoRMwW0ETsc8ke6OcXC3ywWEwUxEOW2yOHeOEdGsp
gXBZvUhqgOPktv2sWVNvgwiC5LhNP/m9mJsjF7dqeop2ZfTR+yfufp14h1MiH4O8QD8kz6DIU0ik
LQ3FmIZyt1rPikQLK13obFatcwCcWs+u2tP/hPr07RCHzHcAXKnli8b7s2ImTV0y81G/+g18Gh8t
GRs0rhsHHQj1H1SsVxv52LlxJ4Lt0KZSwN9nL7sbGtauo/sYeLitWunz1/Jlgy7TnNTmzxz38cFf
D0zGQmxawAtY07I9sxRHlRfqRr9LtoMwbEBgotO0rBWn/PUGbyBXfidJqtCergT9bG5xdW9bI48V
+cKWXmo4qVdvM8acCjDGHIdTiFOTv6HPoH0Nca+odRayjl6VJ1vTMGstyTlds1+6eOIsjl9DvLSM
tj/LBTjHQYzdnMrGSjJhH8Z8DoPKjDDPnjvp0IhqQr4XgYfxDo2nC+6HlvUbGBF/SKh6XVer2hbg
KyOALhEDtnTQ+UD7DsGAFAvBpmVLB2B8UROZPedM5W32kivmYalA9X+EtSyjZyZ9G6zBZKxVGBzI
e7jtCwS081gmF76rUxF/Z9V8gWixWKHO9ZQ2sAdR8EAnIOaBXm56XIR4Z3s/S0htauAOcL/jPzHY
0xLurLz6Ekkt952Qug/PwzQJ38ZkLW+O27oWzVG3koMzVP3PzjCUqFNfQMsDeJXRu+7xvNBosj5z
r6/Km7Yf5Jjff/EsB+pExacwCYZc7evPQgKGxwsS0EmnK+EWy4k4RCJNaoOT5Dm07V+2fNAccPtH
oDpxvqudkJNoLG5YWyO9D2ZJPj6pEzp7WqMXQ3U7or/D9674581pVdG7/8OwsLDQQ1EzHb8v1c2C
shx1kOsgleeWFIqny14wno9ipsMYbpD3zR0CE/w6HMLIApml0rxmLscjoe9N9+o2XZfsxeBVua6o
uFQpDJidFTGA29RZyPU7lOpjLrakkwer2qDg5lY2dHUdX+mndjxj3UM7s4lYem8Od7pEAagFWUsd
XV25QFrDgH0ceuuWi+8k1P6zqu2m4OdZgOZnpqWfAQGcbPHRFqREb28GAgMr1RFvzi1wf3pkqpT1
5o1zk/N8QhAZ8TbWXWhJQUCrGaxLho5X6xesXD0EOoClEndNhDN4r1QJOUk/Oyrndkd4o8ETBVSA
HQYT0SbgcQShf+385Rx+R7MMbBX+Wp/Rq6hSa3Wk85UCuimtG6TdlsRQKXUT0dda5ouexx8XxfpM
1nLq9VirAguE7UYm3UAwh22nh4gNAQYQNJgidMiJZ4TJVwxLeV3uP5xO8TAb7Sk/7vmt7UoPn9RZ
4dBVRKrD7hwm4f/ITM5yF2icWumljzimztrMleGFpOmtZC4lfcCd7I8L5/FsJbcxZwpOlaFY5tsH
1h5UMpMx/vbf9PU/Pk2w+/YRqrnzLMPqEKU8mwfB9SIE5UA5bQiFnE7yZ0w4X9/MyCWA/cbUpfDA
a6QHSQXFtmNiyQ/Mn4qoEiHAij3zUZ3fV2NIBPbad8ClQ6YcvpaMIedakNUSL/3Vob1BKyS+Rsn2
wiWh21MNyH1m6cUtkcHiTGd/XqubXAd4USSi/7Fa159umwzJPMxscxBe6Ql1ifNL5zuc4pjwHOSs
NfAFTwkwjkPkDAdT7t560ZJcmwy/YgBHdUrgyqbnr3L7d5L86dQZzgRhxPD953gzQ/jw8r20PmLu
/rI1cxd4wZed+S4DMrHP02mMI2MrDyecZn1asn+AH5sQyD4lp8sOaY8NZfsAvukakGDVUKTwneNk
DfmIBqw79/rChtOloUDR/hybRlq3OQKTeJisVBzI0DmCiKC89kmcjas7aVtIhS24vOpDUVj4jm9l
kuqmmj86FJks8uZTmOIJgkBfGYKjv5fFOABuC0mD0xwPzwplTQWbpRkZ+zU6MbTt915rkygO5vae
+3qZfPuLRxzhktzYvfJMgmiazAz46ot/bSPBkxunlgc6F3E8a9XegO7NGQ49uw4hKjY/rVIekabO
wJX8UabIbeoEWf4e1IKrdThru0xbZRO98CS0wvzveeBr0r2+69f9VtLK9qXM3Ya37XtiDxq/Zc50
wxyqK1ffpk0fffUXeW/Eg/SeS2n7Pqb7GLYwhIzM4mmgAmYVPb9lfcJUBbbM1+KqyGyBYDzEn+Vl
rGH7zlM3pebS1IIy9q/+2FxIYaF0ulqb7aqBZxwsuAAXXQYq4zxNaxdvK5zwj2V7CIMNdbaSva+p
mt/bnI7ZEP+W9kSc8Sr7KMlUMLKALYfGJvraZgFPDfnKBpKiqt2LpyPKycGaWdhu7lXxt+rhpr88
odMsu/Pkxjxn278KW+G0TtC4MtA16wqjrgdMJQOuIhr94kgWoY4w8LfM7g0XvQcHQ2gESs7h3yiV
EZTq8L2m6dmtsOt1ZsUOumNZ1Pl5V0mdlc04UjeIsw0+Vp0L5Ju3DmnfK5NwK01Dg8WE+MBCBidq
7P7husnyDMuZDi1OQvKPEMhsfMFqsE4mWZm1iVPDsy8zLghtAtSK419/7fK/uHrC87AMZJkNdykY
WsYDMCdfrOUnuylIDM/ndAJ4XSJRo2/hTbGdRD6xkUU3f0PArw6orgSoSgNOuC8aN/ghRaOwUXH4
vB9P00178ApbdyojCGIAADCM4ch/50buDoRdcrX3UMgn1q2CQktkIkaAO4kqV4Y2X2FbBDIp7J0P
s+1FDACxfyr38Za8GxaJM48/xkPvdRDDY8fQ/JFnvlUb+3mSzCd0J6CEZuZA7DKzX1cbij19bNlL
4IBLGHRJKCUpJyp4WCdJhrimhwsu4EdPOCnbjfs+g1exq1nPs9DkRDTP0xIei/mG79Jf2zM0ycH/
MT7HrAkfP+NaL/1FD+iGm9kajfSt3RMASA/eIkcTNgNm53VaIC5SvLkEYhXnVF/7qWfpsgginvas
XZaehHCK69DJnLLQ3Uv8DBdIkQtXk6/CfB1hkkMm1MCHVZe4pbxKWxzsE1WYIYmOg0sthPtF/xdW
b1bkIsfyYA8W9X4tiXYS0I47VHuVuP7q9DH/B/kGEaRR6QYR2BZVXGGhrKcalGDcVIoiC99sJ0+a
g0yVH8Jiz3gq5Irxr2zKHJ1EqUhWSpoV0HD9n51d9IdqUbOGpdndsA0Y43rCjA7bllddNEnRrXSc
95Sd1WyhPXnj+txHfkpIcxYxk+l2N2djIAf6Qn8glMBy6cyPPnd03taMFJ6thPgkaVop/XSja6u+
dFkks3kcQu1qW09eCuDcsw2FNFUY/WUKLutr5DvJ1lU62lZ5mIxD4w9iWC2CTnUSr+2lAska/oO8
zBgX9BRfxR2j2hDrnzbANVpyIt4CZ+ruZJ+TpKfX/X4AhYAzf3QEo05X3QxOCJIsodDnXB/EXIJs
+UISFb3cJdS9BXLR4ESQ2ShNLo1fP3le5eH5jDEZbatmnv79+QxfdaVsDJzXqgZWO5aHqFDacgVz
c8ZjZm7fhYl/V96QCNpAthVFEsoK/TKD2kByuTQtm5AG5FRb+lZX3U5ZgdU2EYwneRh4BjYuunOS
Om0FC32DsKlZCB8+F3yNA0NwrwmCkgm1NhFDCU+B00sC+LMc2BCfbPOlMJnkG0vFT33qZWbsGhF8
wCv8ARwfzxfvoIrhZl4ZgciqlRahVNGpUFA2E+YkZdQjihr8r1M8blIlKzKLJYrw68DN7febGdZK
J8a3uJ+o+2qMzNsuueVLolipYrsPzivngRyjzUuy6rruxSAmUXkHj/cbfpD9Ccqx07c/+u40Ivhk
wt7+I8PRxH8FbUnV3CPWzZHzVxwqoxk6DHYjPi9INWDQkRZ/dbhjyqYvs+hNBKiGSH5daC8FvB+H
eXDqhHZCEJtvApV7B9m/duddJ+izD2Wneq/PxT7/b0EYgUz+G3ExWbJohBPJw7FRIiw68PNpqO3N
iIsNacZkhxOKcwNKkes6k3xrK12iXOP9NpBubDvVTH0vCxklTy/3/Jmd1u8W9gV5Ep7mPBhvdV8k
ju8vrkLjahHXmNSV5TrswmF9vzduYD8iNyYYtlEYYVWx4l1zk+DmeiC0aQ7ClSx+ifvv1Gi9LQ2Z
mlr6HSHpOsRg7QxNzIEOPM4rcTgIhUvtjeHukYNlEncOMD/dVGNE//0u6lJstLanb0rSauTKo2cc
x6cD9Gq1JMgOzupqICfKKVmf4XTiv3Zt6BiYSL+oodomjMSyincrfpZ3HOebfXZneFATPPspurwX
T5BlaMsQCpwy6oYL3ObvG+QbXfdiDu6EXSpECM8bFWn/2MYlNmiXSmi7nhYqLpHvV0kY7GA6p9jl
eBPKLOk9ap3cROry7snHFlC1sAA+smkoJwy94eoQe2Q7ns29olq4pBSIhoVx0ZgdfCd0oAhmFPro
q0ZSxy/ovjFPTmu0B6xSFkoItJiUjYlsblEezSqa61JWgTEvEG7qvK/31TRfK4jMGoIynl1SzWRS
/72EwHwc/5T4lHX+2i2PsPxHE8kinr/utyEipsZM+lu/T2E7B2Pd+P93/6oXOusEBFrxSIF4wxIS
bR022TIX8N5/5WrW5ABB/cSWpyHI8eBGe7+hhNh1JmzBEHY3xtrFim5N2E4CdXUWNfs/IrR7w160
oIPauMGNX4MSZGRGsdP9UlEUWePAS5dwdNbBrt0IRii9YiLy3ZMzyeB0er0fPfTWJddLb5V7FHo5
NFyN8Tu/mUNImwB4Kg3++qx6fZWvxYUpeyTBBl3qrxkuw88babJHs0GopaNck7s/eXfHQfNOxdjj
TVDHalPDYa0r7JyY98Za6dJ3UtCmbelACo/uOs3j3Eqe6TzIOiS5puN+61FekpmiV5NjstF2AzPG
7D21rfUJ+nNST6R9amzMTJo0oBf5diMbrRPMOohrHwjhQvMtMgdVoIFy/J1yOODSfvhFJdAlsy9C
YgFF/yd2aHkgpTLR1Caz8tAuRaQhW8Wv+hsPtlGxQ5gqeJwZyJHQtxOfcA/yXWbD6vORp3heiZLq
SpheYqm5ElW48iVvVAXYBQJpDz3qZojwVfp+13Sgif9LDUdzF1HZ+CRl4ZCz6NR3hCF3S/pWksXp
jiUgNabN4UE6tKKedDlRiipq5QKFmlLON7X9pIJUimOdZz7N6iNzydqvRzyNbM2E2f26mlxDAkM4
eS1QoWhwF8knVbg4/auteLYcCDHMs7vam8RJsuqBV++TjCA20PAUbwi2ISPALbVAuilMLxU24SNs
TVVgMFp++lzbobOYTlgyyepbRloBxH2cz7K6nuPdp8XH6GciPYulluEug4+14F9MCvl5WR6vgFN/
InlBMFxSeQQQMr3fQBScLPLuNu7ow50d+28OhEvGieRC69gx8kCwpc0NM8eXN/h8VKw0QjmIHw8g
pHO1F2ql0KJvt8Y3Y2LVDv1ofuEmB92+Un8O9EGrKES3LIT84yUJoQlVuOU0JjkOWqHLQoLD/HO5
ZQBo+cV7dNB797tedSkTnmeUNNhlDyr3YDDXYnBRyvaxQOT2HuCtgXdBM4E/FLOPG+PNnB0uDAe/
8pS84omdUU63VeiOL5fJtZmS5z/q+axtxeKCl4LedMXbVohYqeTJGCyL/xIbxkZ7yFjH2ooEIvCB
6OIkE66d1eMzW+FRDzWohbJIIeHafsrGsuT/PEvrmrXF0JpSO/rnsiJw9hTKOIWcQi1wH5BgWj19
y0Dv/nuofO7+F3BZGt8INWG+jQ2pAHF2UVTD7OUYwmtwFTRPxZRDcZ6JBemDKjoHByHqQnPqnBCE
+ZOTMRZRkHQAgDqUa3lULTqLkyNULbhFuVcsSAfBjA51Y1mH9Z/sxfnvfoENvTFjBcWJtwmAQP5F
Z0xQndDBPK+7n0bdhBnHm0etO3Fop65Eu+RVipHwHrqkDNPYQ2r+difKaxrb4/ioA8b4DGJDdxzT
Z8lMVNl/4PfT6msttxEtA1UzdNt0YjZmFAcvVPXWvnziT5PQ1agNUqmn4/tw4FSQyT4dLEs/O0ze
0ot/Zj/zoVuo7ztpThhrRG06J6neItovJQgX3VuGI0ns3A1XpCYWCTbM6YoCihVw0ygyEXnT/GjO
rAMbCOKPWLlZZueclOXCFxZ7YecAuuL1SeNZDek1xBJPOjznG2UBvrlMN5yRmH+cSv2AwgN3OEem
Bn9AeSjfKiNuZt34QFOES7XIheCUEfgsgI7448sV9qm9DbWfAo5ADaB1k/nKak705ObO9EQh72qd
V524Ak8uitCPh5TdzcSnVYX/NqU6rU4eSPxX0QSi396Cn9qT9s7B1aE6dz0HZfLJE1g5FWO1q4YB
gILSqeqYhBReI4O42zkw1ms2CrICy11bIwLFM2/zkOchyOBUIE43H7yhQiwKQ4hDhavPYKWy+9Ue
T9t6effd2Mgai2ebggnaAqUgYVNDFUjrtlLvnnKWrx67SRw/n6mZugWeCuILfsPQG/8fIC3OUczs
b58hFR+j7dxCuOsWloROPThpUI0MoqnUNs24gGBwdItz9FXa+yet2bveRsA/jDIjmRWjsFvl5/2A
UMwoYs1TKY1jwBNo1cxTb/620MZEYkxhOCnyREzqo/a/BYfLafxKobirvMpdHGuVBPPMRn2Q09wp
iDliEKdLqQcZuM+cTFiVIdBjUm1lOilplyqR4aXxlg3BHlwZwYLlV8ABBxCqiL6Bh0OOaDuazwYm
edbvUenhscacJVRlZS6n+L6zpePbCazLgHDuJn5pQBgnIdofU9C4OzXIXTVrttcle4d7wFsczRkp
6ZjpaEpJJ05Onlgkn7CNfnNyQL4IvB7qPqNS/TOwBCyCLe/WnOiICX61S3QGr9B+/Vm4oTmy8Tgh
lGXs/ydpbVijW/hpnzp/tJ3ACDwLLqARelcnzlRDiDT2toJ6CmZTwe8kHSCw5OTSgwyPibDs+e+T
PgWzKJ5LG30a6WaZj6ziRUok4NXQk9Qre+AAiO/0BHfbFlBH9Aqw/TJibO4aWlda9re6UnQtVGEo
FbyhXOgheSUjsmWsdCCJVZ7j4r9sTpVP3ohZMoXZn2etmrbwoHxyts5f3PR5/NEZAyrd2cPl5rqk
OPrDrgtzjWgbSesM6mefmQjpSKfP4n8HFUvAD3R7BXt4fmeRzeU7lI7jkT1UNujyylIv2A5S2XHE
PHlql2CjcHjDykGE5Bovoa/LKzKKMdtLgf62xAQ5FG2PYSjYm7rtTwy70wgfzA6J0Vw+relcnWtL
F7jdCjc14u53+nLfqcfZm6RgvJYgbx1S80HBROeCbl7VIYSLUywKsl2PnzUyE+ptdNvybcihtAm8
2akoEqtigmxwHv201K65xTYizUZLaLMzyj8QU81NPC/cMSCmIfXBkixVK2zmRsTB5+cw04+oC6Bw
Qpr8U8hsxP3Avz4/VcBhZdnqk3ytgRcVcbbE8fwxHvoCickj/c9Mz60fekiW1caw1LBlpkrk3X4M
o+aT50ZhyriUd4NBKQorD4P2KvkYDoWMsMGJlPPJOzs+GtJPg0BjigTC05UlTyFS0ZKiWU3lI1aJ
XlzdRP6B6vHXWSJ0UVBCz9RLPue+piRhG47yvO2NSMX9ykjiVeaVtlEnd/C+s8coaZ48mPrmT++/
ABWwANJ41v0LyCvU1KN+crTPUQUDThY8kwZN2QywW2rmOlLU3rw2bJxHFukbK/A9bJIWzYI8G2P2
RQZhxLKMg17vcoEZ2bMedw6nVyXUlU28L1wDxFN/bm06l0Ug9awDFnoF08v6MxPUulbyJex+UG4l
PshlcR5IAR8D0bKdcmPqCEoR7I79+FXOF5jXAJKK6eo35jCkCciWATuQC61PF77098m5W7L/HJHb
8sHc8n1+HAhW9ywq8mazduyDnO88NH+aww8g3O79GmqSFCQqAZnn5uOGOWaUrQ2ObhplcrR539JY
tkadPEJm9Q8OItqH9Tt5lwSa5/nWqMhGPhVCqyAI4IOVg7Ds9i62TSha/32iMtNeJWihFfXgHW+A
fCSqYjWswVzN/o/jz5s4V60FI9Lr7R/dOKVUJBx/Jhl6CTzcaGcUyWFXMLB4Rnbrv2ioVMiFKuO5
8miXT/cCRYwg//wV/1p0yzT/QeGxjkwZbi6eyU04PLzeb0v8Iya9xG+zS73oPBvFKlO7wlWaCTRQ
wBEy2v38qU0m75BtqWYZQYD64r6V+sVjus04x5vyKQiymgJShYsQGBaU7Ti3J56iDIKn0uUGJ4oO
CJIsJfR38naxVJr/IIQMBCJDW2+p51luvJpV5piToimlWkvLO1lOmXavfbRzIv6CTQKcLb295Zh0
lwRsO0ykJGr+Acq16SH7JuaaqjGA0SbXlaphW+Y7eKF5Ihx37QBX2dmQpkATlxHjUnjfvv/7UQQ3
r3B3jqdRt3Ax+UZmZXCVxyJZ29PCbJ9/idy6xfz9HTFom46bAzBpoJii/eIx7H2mpPg1+5TYwhe6
V1ED/Fv56gqXU1BsCce4tlB+ngjK09wQxZtcJs9dNGuCtNxfpCJgpwbjZ5vevjoRWhY/qOYkBDqZ
hVUpWEsjgYIlGNRqyaUvmiO73Ls9GKoy0DN/s5urYJ9V6QEMe1mIDIDmcJ+DDKc7FE8hqUruacjP
NoRUG4qVUkrFcd8G+cOGVQB1rqzGXsM7E5SM1PCSVpmr3N5rCjOBwochs1LyBwVFui7W/bucYfKi
/5VW4z5Rm1IPnGTm0fM9+GgexJ89drmyW1c7WwztlHDNxRijjSuiYhXuO1rKlT6Yo/cagxXbnfYr
r1B4wXKT/txonETnEO+m0tBnF+TMWA8AdMimnWHnPm+nJ8wmJ7Vzptgp8aMokCNqpyCy1D7AD3/+
CwnAmuQdaaQ2Z/j7KV2B59mnmPVdAs4bEArZHYynxt+Gmrr9qeY+js7eNAeqwY4Ltn6dlKnAbqeN
wFL0p5vukw+5t0gjSPLI7uQL1fbo4Y7+R3Scg2vrgfdqHqfMc711mZ3F4I9nLTLpZ0Ug0JU7n1EF
GAuGs+lSB44+7ZRlaY582kXDyb9Am9OfJHtMMTnFnrxiCB1Toe/Ihc8uSNV4qlanGe24+IrQFo+u
G8LWmI4yYlcGTGyESw5NKaRrwwJ+eFtuW36eJzuk72cf1PHs6cWbOQvMza08zvPetJIkhDng5M6M
6RIFeGCvkhv7eYamY/QPh/Aa2gN7FH5j0oH0xUD2d2idF/tZpqCdRmOH0O6j7yMyAQDltlCVe45m
0zmYk9Sv07nxFYJ2oZ/qHjDzViFU+2NZN1j787xE9uqXOeHq8/IFWiiy6f7WF8HGa9RFFlBLxP8e
gPKjeluasqPLBGILDD4ejILIfdpyyN1z6/hyi2qeqE88CYLwjpCVgZ8MChBUN+dl7qqWfm6EzcJm
vEi+n04m4FtPsuRW+oJJCY+iBuTx01Z9U9GinUAQQ2BoOizH7hJEOSWJcdtNwt++7s2FLidy6sNB
SYvIw43L6IanPbW4+hcyplaNlBSGsZ8L9c/o37gnS++pjQEc2z/aOrumlphepYgzk8KK07A4eENq
OGDzGzA8cOXsr8mkYLpp5tFJfOWR9D56LBwdJ/Mn6uvxcJTFsPmtCKquv04Uc8F4hlvf/Pv03mpa
XpfM8r/ItxUC8dH7sB5zLOAm8qauouvdTnBqAilQ/Lwb7hqOZgfS2R3la7zEBH+rgPRwC5+ex1nY
6Vc+qp8Wk4H6JWewAHGq0ST3JFPBhIAi9ZXA3D1FxvGSFbx3wDoPn/AMx8Ih2576DDasdQTLENEu
lv4ZHlfg8xRQ3KrYxsXOULS9Tvv1V72yjPPfVjYha9ZrTZq6wyPYXJYAqFOJimzUqpncZYvVmfpr
YRhdqS7pfzDVz6xbulxMgp9xJ+z7fWHaEoRWYoVuY7l9FJkliskDWswjEJiH8yvgdXszGJOxmQ1t
WPXYFo7jO371M7rZdauU/zrK0P1D+3QDFbBxCaBoguSowiaCkKUs5Ux74aw6Cf+QzYL4/l7iK63D
WVp1JVEw30rE8JybTGfwE+sj+eGSJNPMquCvFIhpWXQ9od68Sg1V8771ihqnVwMBDkPYTEfhDo1m
thmYwtY+vuIOcbjxwug1Xdo98aJHy0n0mqKBq/ytlp0Jv20UxPHefztHeMunHzy0QDGKiO8mlb6K
kIUsA7N06xy2zkfGS/HQ0+Iw4gq8ndY7Gc+A/8Tjv2EDnVXEecBEEZfR4JoXw1v4K0p5UlokwALu
Xreu4MDHVSCSANdzQKdjGCVueoLcOSVyJTkpxRGAc1y89glRiPPoszfItL/R/7OPUJtufkT3Sh3+
ICogidCfhRMdW7IDOOb/QY9l7ZSCGTGd5jrAtwFC1tOty0emyEY9kIpbuxkrdREalMd6re5Nn2gV
qJYa6hK95jQMTv3XyW9vABRUuLfJq88UpaGdVk6Z05JD4koJ8Ht25xi2RHDaBjjmWL1iju7tBDV0
9w+3xZ5Y3lwR+GQcJTiQPKFJGvKAvQemCLLuQD2M3ONBM/7xUUT6YqTmkg41fr1T7x2BQxq0wblY
Nx4H1M4ObnbW1HO5Cn1gGsSNDOr4A/PEh1khf0IG7e7ItXglApENUURw2mSq8SkljzVduPDqnzfH
Ow5Bi1L69BGdNIrEYU0/llK8/MaR4UA2TtAI1peEd1tzNmnLgF37OVYO2hAgNa0lWB6ax5DZB0Nx
YwHe6gjPPAq6F7GSHEhkyTrBDyqMu6WsQgJpPpkbsLCe6gkv0nN25E4D1yskzmUwMT1/2lvuc+H/
sDeaERWFefZ2EEfD3t3hGP+CUhZKUSPT+pC6yFyBFMCeXG4cN84exgmii6zkOLfHRlmLUSIPu6am
MJv51UWM90zL06AiOo4N3cHuJOF0YWySDpXKbadKcY+dHgzt8wdLYXFBwZnVLl8J0yia/stGLXQp
/Iicv2gtZERe4lVHv/Couqnuats6QLPwB63YpgeBfj0tjckpv96qO2R1b3DnpIkcZJvYRv+av1qL
+3Cz95U0WNWMywWNyQa0C8BTIjn1Onpvl1eWoWn4OaEhjeW98dUZ2VwcMII5JUXLSnjTM6wFiQQi
S4a1KnKbcsDCdMu8EDz6oDQrKjeBY5hiWxa4RG7qyzviTf0fbB5HBZzt0t1TZoBaNckaBTF8sd8Q
Kr/K7kEfDTTwGUlf/sJZEV9SQaZ9gnl4qWpsUSp5jVgUI0I4cDWoz5dp9y7XmvPfvWCkSY11fEQz
s0yE9nyE9vt/R59qdK8pRWwf2H6NANO7Nnp8pXqVWWAvuTNZTW8J6JL+aR8QwHAdJg6UlV69iBYV
MF454WldbLU9zgjNRKHtWixLptnFw90x3s2uKVQ5XVKxKOblv7vkM226bACW+1SHxEepexZbZ4zO
umXN0+vIl/sDEgMXYvJz0LB2mJawA0LZ+M3MwSf6U/vEqQwfoB9SPHj0rx3cpxle+OocDu/FDp0F
ZLkiC+VzdtjKpzZ7993ksgW66ZOnc+RfwX/EKW+FGgAN7DMYHe8ZM39orZ1lFl97ANSBqYg6M3sn
1oRd22yw1wUSvkY4G5w0q9UEsOImrm+64XfjB5mJOylwFOuwhjjIZJDrhIOkwHT8kNalXf0TvapA
siHgdp95l/eMAqD6Dvm9GEob7E6CV0RmJ7LykNkwO1U4CAaZbDpnT7E0j8UTiyy23s9Bax9GeTy1
Qgo09MosPXzv/fPzhKn+PSaq4mlOJkLlsjmkCW/7pEr0Fn0P8EIaAfOlqOjPCG0hKSKZUgjmvR5S
ULhCe7NhJ4IqfpOuNxr6C6zAfhcJQ2b2DJqFtcpGS6jiZVzd9yPDvLadomzOAZlH2NZ+Zu/HfbVt
BhUs6wp4Y589uX0bXi6sTSKwiIP1WTGeavxj/fTD/DeS0mrL1h3cJafzjLm+5IbZZZ1cL6qT/HBT
lhHbOP6JHmBEBtmCNc+J02rJ3F0TKQ9U6RjLNAh0NgTZlbjC2/pe4VMCuja6ll4N8WVgvIO9GtUv
QjJ8kZdMQjicAL9CJxHrqiZLsZzLBDNLdF32dv1+w7Wapf2P1h+xxn6UQpdfSzP+U+onz83RMm8y
o7yyycbpbjjkZ2jeXsBhMWQhCC7ODFjVsZzJjycVQ9CkXYUUN3NXRtwMIgtfwP7hPdMbI8i58l6l
aHqk2PR/rKT6o0K63G15OJZpWy755uLfDjOmV1N3eRbMRvTOS7i6VFqimEmQj90v2/UWfAbBQM10
xPwOhuOup4ufWKWdWCHiRv29Jpm7yHJpOG8g3dnY5E6S/Vz+3p0O5JhaNhAET/lWEQrqedi3NwTK
pQW+hjPcjBD5zgsckIApH25Alc6iacz1KvRUwgGD7byaXFsxLDWdCH4PzHwdWy/+E0AwJEH2lk1A
I4UVXyrIyI3qtOiaX9WyUN8E3Joy8EcoACdLITN1ZA4VQqYBb03TvpfLgJwi7ikYAGlF/5PkKVlH
ZJh4d/Mw99FkKSeBZIzdBZE7kmFBS9Dr5ST1p+1Eg7kVjLSwh4kzwJSxklyrut1Gg3FcngRsOgnB
JVmp4gAacyON8RUfHuErCFqJbliyww+7jEUwecyTt964cTRjlYwZm+gdwK7XWf0PAMSiS09res+C
IxpCToicMrpcO9Aersgkfhv3s9Rw+ALqvko1cfG/9yiaEpqkYHwEjaASvhXvzBqK+HOsO4twt2hQ
SBp47P0PFG0gp8v+fIrnNJFSygGlBePSSRGotAdPcHA8daO5v9nNXSb/x92gKh41991egscrfu9j
vS3pu76AMRba8P//G9Se9FIhxcEkX+E0SFSp/NeH6/UhKTguP4cfRT4HEA1yc8hETJuWKOQRE1lh
rVozZWAtq0Srvinx2o3w1cb4zv8vnPEhaWRyMxbVtmUHg8zQssNURXoszZgbMCclDzdw5vSd1ShW
ZKz4GtdyXWPCXeGnHzbb3GXE8rTfZLhOlvtedMnpLA0/05zirLnbn0NjI0ILFKmSBig5/0nX8EHl
nCpBLgE08CeZ8AIpDYoID4Cd0uely3xhzOUKuhgUeV7azD6C1fAbFTbWTKdJnF5k0h+Id4N4f2Hi
1mMY3zDJ8RCHSsRz8TomGKniBjJwqb3RqgWHqyiYMCeti4grd22ibODTCkJmsOWItGBiPGXn7ZAO
jc7bEaiYF8Zj6Tl0VbJ62gzqRo1N7l0LCwIXpl7b7SqYhjBCj10+GzGm4sytvF/8n44zXjJ/X+na
YyWq0hHgUmlABfFF24+x0QpMRCMIxJ+0RZmkhcWtiNv690m/p5mm4GnuA8fY35k3kkI2cwY5PbRV
vqgObMOWfysKFuq+RcSe6liH7KV1DPuS3aGDqQ9/5d3bRG6BuUxEXAMvdv6vlBPK1EyhAZc73Ewq
r8+2OJkN7Hldq2ttZOjpn8ak63OnoNARJWOKNUqxYpd5RKlCDoupJxdlSWeNuHo59ykO14d45ZrB
vmVKJuOtL6I+vWmsGOZdXD/zIh6Wfz7bqP2KZIRuldr9NJBVTuRdN28tGCcvpjqkLZZtI4qwZbLZ
fihUSqNEU5LYhnINk4aXir/MReHvwwgQoVzqk9tuF6FQYupXh8vHownPbmcRsUuq89gq6zGm25MP
eHG5X+CDRnxwOOtBbR+2F6k/1pv0DPteoWo9thMGWneTpviX7zDxTU/XqaOc49zJTmSXfH9+l+uP
2hRAIcCKsDSLbYmCYqK4zJPUzOELd9TIiWKJNGx3pn9WRPFsspxM7oy7VKHVFcPs4EvfSgwr+l5D
WG4ObYVfw2QqGxFA3B/+AIZ5EhXQ9RVuUuYskoRZFvEVwUuYfMyQERo5Karw7iRZKuzCKQnAS6N0
oYg63B0WjwG/MAD4rlUBo7NtjLrNaMz7O3VYb7tdKZlmUJ3SBdz89F+U6DFMcjjcnTE0Amk2tXWX
OPsH7TRKE4u5KjV4WpVOdW3A56fczkvNWixecrpri2qnuhiHhYBOm9lXG2iBrOHHwGMBNNDPvR98
NOEn328NmwC0fuZSAJh9a3c0P1VpAdH2I4mVCYW/1FKq4gsT5bXvgAfOZ/Z2EcbZ0gOBfd/+JjIg
Tse3oqjxGrfUFlR8JvHcOmNTzeOoWxJaxksuCKwweuvpbYldv2a0+3asqPeUjtBCI9j7yreRfF/k
vfdBfoij+mHR0fQkk/nnIXtJDeX3JWj/1bw0sIRGljljsmuoWXoRZibrDX2XnmSTY1Z+X3a1gL1N
eWBE9EUxqePgrpbnYx+aOzsJ4jiSOFqttut+2emgY3YpqAvBYBCT7/gjvWVudqfrqN2JbF8t9gys
G+JdzWITj3vSqH8xRk/mUmdl7qws7bh3pjQMcI7fyILQoOtMWhkbW+2/9BNKlSt+mYj7fFbdIv1s
FMaVHowNhsf+J4k9AW0grFVGxd0tu7gmBtt2qzZmMYwM3urhCWE2e54uVsVR+oYjSKKiga9Xf981
i773jNCd4+jhL11WpJ3h7Trkz+NrajAh7fa+lpYnAMh9vQocnLYVN6jkuFwHnjqwKiM57etby7k7
WzsFSJJ3VLo7LKLgUzSuN/s/+71cwHuiWN6+/9JARkTrzdnGJ4GSzWsicapJFS4tBVIgYpRvZYam
ijbuPaxX+hnyeWwJTx9Oz1fAZpDBXiUVqFdilTDxKGmC66Uanklxb0Nner1L6C/ApSfmT9aFjwoi
3YKJs9pUB0urQoISVTgGnIpClR++eN+Yeex0KThYR4ItruxfsCbCTepezR7LEPAV2XExESe18qZt
Tes3mOga5YRckdizzEUb0ncWS171Mq1cGT0Jwk19+buXcq86z5sRpX8EhVJolD466nviONEtOwQZ
JvpbRwbwwMuLKkHA/sXGDW4S0i01wFtvk/d12zFkCwomTEz3z+MANUER5fbIrhf4BCEIzCz0NEhM
haZX/OFXL2NATPvbQV/IeuqwskAMZyyH/Ss/c4O3Qx2c362ZFpHuLXZb9CRcmh5pwbfesxmUDQ5x
A9ZQ87VI51dEvqlsmdc+jhDjv7pMkJYxXcoaoGR1n+rqdnqgGBIvMmW3qxG7/cpx+76/6ISghKxu
IUbr54IpTQV+YrB6uy6Lo2A8TctWq5UYQdTpF9DY6s1u6bN7BsotbXAHBwHYNHYycq7gX7Rswcrm
cIWyRThRJpx+O51A+IkursIir/Q4n9AyVD3yigWme1Pr/p5/JQmkn1tR/sTHTCVU0Phkz4qXt4Fa
SR2p18FR+H8TiWqgL2GqB0Pt/ZkV75+cRgkk29/EQprtr37LgnNjcdO44F410MuRXRtuJ6ElBD6Z
F+hii9+cdhFpouNGIrNyC2rfp+ay1DDJtS2K5ClZOOT6SONd5JqLguA3Hy87duLgiHI14n3VProD
MNql+YcPru9f9YsOCst65KPVrOqEzbnwmzihWalFyRERuUwtvSu4Nq1K6Y+4uF7q7qTT79KWJqmN
BfDxHW4gEJoCHTgQxT+OhVgjBYAMdfFKLZj9wyh9Heh3YzB4648BO09qWq5HQT9a6sNP8gE2STRP
lfBjRrpjXemFOhrXCUd64NgAYN5QlKe35klG1lLhvpkKvhwiFR92hD2IV6+GepuEbUOIKi/xHtDU
lH+xi+sx2anShacXMj7c5oZISzd3Xpe/8/pRt7j0wtlZz+OyEpG/bnjPSUqsm/Iz5yaq5s+kCRHm
sMh2fgAiv/+O4531iROxX0EkOHz7EaMjmZzb+u89Ig8n3TcUW4nmbWNHSwWjJYT12ZmAJw9bsgKY
rQ/0h4KstBJwus0D8VdBomcRZZ+TuLYXH3wVPR+QJ9jLPGenrHgw9iwLYn+OCOsKSI6XGflCtSst
m3EcrJ4yTy14yVbQ1EhjCOM8mmtlnltbUTVfAQ0g6XZOKB1kai0HM3pVWjTnrQSc6zzkId2iDmXt
T2iwHliYaA7fLPsIeeSrm2ZwwCYeIqPmDzVwYp03kCILzQYU9if9L/k35y5FCeCQGyLJ6GfabUar
seUBas7TLJMmNFgImvNnzXVEl8FX66krfy8ZTtyXo1O8xDoYQ2GeZKG5TmztRoh8ARJDggfgG4dc
fs9CJ56khKou33B7aIcag0IHGldZADNR8/ejaadZpyDdx36N/SBdDOXGlT4/RFIyYp/n2mLBuusl
LkSqTn3v3czK4jZ4smTNl6IyPLpxZNrSrFSRF2fniuLYf6qljBGgqvC277mYqZhnI9s84kaWhsyV
6EOemii0Qd04wWzaiPRdoY1jojL3dqd3NoV9agrtHvGy9aUL3gzw0MFlf2S5l0mbkWCwLhWbLI9u
ZgZhghHq+Z0bfqqeqfWMFT8I/kpZcV1Z6qL8pxMlcjm2An/OtqB9F3sXMrxq+ucQ5Q3VYOww4hNl
jNrAmLQzspzE7e4+YXJuydOySiMfnRqv8fFvM3UMLY8844fN6TJeOyDUKbZlRmGVn1tYaPTt2QuF
AkxHOEQtw5eMoh96raiwX6lzMLJb0sAA1UG8+GlHZOhsohArk+0Jy0QeL6G5MvxNH7P5MMEfluUm
AXvSxer3kmhO2BnORJEdSdIcS/RHzR0gomuuxRX7CnQQ3K5ZiB9Ox4MxLknWMTEg5WJOR4cDMHoz
y60Mlk+4cwqWHktv2P4uhL9qmNIW9/gvq34GOPTvo96fmQr1U+JYn4R8ufu70/tdtsYV4hzXoFg3
3sUsiUGRg/c6iGEnnMDRNPxe3RvWKn4xkRElyEEGVp7mDRr0uhuWOwBkkxvRCiI6RnChpI57mXw3
EFEwzSF+InsTR9+pw7lyrkPhcUagPnhUZWKrxFAbQ0YAO6ms8WUYl+7CIB/dIfC7Xu3deAOdn2PF
y376p4EqN1cXpO67Oy2GJlb65iDVXpmRRWHvN9tVEyv9Pk6rkc2kRr0dX6d0wgMQODkv13hW/nuz
C/2iVQ+dmeYKyXkE5cHninQ4D0CKSUNpMSTk28Sd3yeSerlVAgYg7IfV8KJlKLQ+3aU4/Q3MBKqt
h3UYQkMP9LFtmHzPp5HMJstOMzLl1b/7AW1Fi/IfHr9S+AuEs8Ya/3cys8B/ufIXxK/ovGFmpucX
IcARQ9wxJjF7Ph3N8nJAbMTaLyup0yclN6QUW/GwtboTmrCJbHCoRARXcuBIdM4P/2BwP2qYKWI1
kXqdfx25OxvomjsNapv4LFNYJTkZJsqxLkg/L27uu3QKK5n5H44CT85yuR0ez22yA1RjdPsHjLnq
EHmHlJx53KuaSkNEvw2hYhShibD30SO9+2SmZeV6Njw2gCboQldZ2swFe3kcm78dqkXzXgHQmwID
oN3VeitKg98c12oaIwVFxwqyrHSWJjQmJmKFG51pVCj/cb3b+KeypCNqD4AePBRROS0wKMmCOTcI
JR/NoM+J9bFBsWl0xZ4DjdiP+UguE2jtMHCHEt/QGfFhtD9YRJ6Jc7HyyXIj/EftEAVi5rDFFQ2V
NCGbCnla933AebH85i1TfEA6vBnWXjHAw96xVk3qkuFhkV+RLC41bMlgH5oP2EnH65q9Vriio94+
aObEBSQ5jI6lvDw6kfb9hm/gNJJtlswZ6M/nnRjpln9fHpVuJQ0izIl+oake8udyfwJPV9gzLU7T
D9oqpIz+4xv4weD5aDSJVbycbG/S9yOC0B16XXbgGiufCE2Ijxg38+uLRHrXYmsVcTfSUQHIpQXY
HzbangaelZMM0+mjyNs2k2WDm+Se+cyE9Fzkq012zwCbwfkFv4pXxf/NJHtzl6t/9CjgGHCEtEgF
9i9uGWk8C9CWkTbJRhdPS3T9M4qhDcKs/a1rSfS2DiUkxF640jv/JzUsUegUx/aZ5iG4YHps4bfh
wV/m9cKJTtqcIoYH1MxTfuzoI0p9fB6G+uCPOPmcZTHr5xFIv7O5B39X09++o3zjs+U/dyAwZ5Jg
areMhSsmtLDOq4Czwt31ruwToF5wrKjTGijPcewH9L544n7/t5ng9TUYCOM/3wwDIMfTVufwb9MF
piHF6b/DB/uOzYcds7ZrO5pPsNoRkwvr8VvdPjxVTL4F3M/ne/8du0CuVq4wZh8Yhn3CuzE7uWEZ
MmM5xbIbcUcVTAhSHHKAp+4P2ZZzeeHF+qFpfHTlLVSiTcDb8hCxG9c+cB4ZWNwVmCoh+j26iku3
HAPQoSD5TUWj37j/geU+/DtDwSpen+EQK/BzQP7ghpv/QEUKxLi8tofu6geDfaYS3Y0LB/s+IKat
I+ELP/MCWXO/N3WttOB/PdleCY2mqw9RtJQwk2Ch8mZ10xbXM8j8F3wrogu0qNbC9hoBOAF7Fa0j
VcR4ISZ6cZRSwwiMQ2gW+yWw5vLpNZv7VX0X1EycSh0iqMHq0hfo7en/fMcguF5WXjdYiOSRZNgm
LiINAAEYMh5zPgE4FmbOE3Qa0R+3PtQKLNtnfU9pvqJPRtwOFcxdWIgMA+Md9GM9PEhBTEOJwbJ5
obb5wC7mh4DQMdrIHrpjfnmEhD8js5DqpjQkButYOQsALceUtgcEnasQdB93bBvdsk9xVLeeNBRB
c6RHj7DJppcc0949D0LmcdxLwcQxFyj6icHTlmm7E7C7thhkYZjr0m27yas6y/OkGbduRKvAXg0R
cgmNueNUMG3553t0JtIkA4TF5JDV64BS+4wNt2BWKWESdfzZzw5HAdHK+uH9ANwWql3EnwSUnLaC
JxQAkgzuKoGoEj2z/cWhTMofmdZBiV5lx8nuPZZOenWmOmdvF8o8XZgokiPubk5usIKe5RPFdUWQ
onCJzQ8S2SodK/APjKucBnoJRXmiwc2CNaJtZ3zgA9BJRGyUmsFhEqtBcVT8kETFms96rCy37gKV
4woMEPxNPfxOuQEPDagMByztfhDKWoytEMq0OSyDhJCpvYmm5zgicdMYcccLegqS8QTHF7uKc1e7
MhLluKVCg74fdgpXVORg+guLUuT/7MPk9KhmNv5ClMUblr8T+p5pTTkEWu08551cvoPpY53rN5dX
feza6SvGa1EvmCJbRYI6RauOmt4ilAODhrtt9S02t1WLbTa1E8MWAmgTEvkSZP0mvTbPt36XLU5k
1RwZGHEMeG1pv/xyaX8pjx4DjEf6yqqGqjY/9LXh17FNSQP6kmhQ1FZGMHtXfnBazZyG7L+Cy/7K
zn9m6cJf/+Rb0ooLRIUWlI/2rRcRWxmYD4uVlmsHEQZJkUvlI7JR/NZQsf0JggzAQ6hVfb1cNvC7
m5EcOJk1QykdqpOhQgUtrN6uCiMID9T7ijpIT+gQwEYGCmrDeNHhm9PdwnegZ7ccGU+YI0VdC6Eb
QU3B8NQpEbpbO9t3jU8ab9r3CB7sT5FFO/PsaHKTUT8PQMqo8sI5hc6Mset+FwNGqEQrXcw0gEXU
7r98+FoWyclQLHazjaIOkbPY3SM/4ntxSAVzO7KzI5ifnDDYX8Jm6AFMtYRwdPi6S1WXWnV+Y9BV
iz4ymNaobvtTqVNXMm23ds6JF099zIEaB0hli5dihaU+h5FVsQ8+dEHgXznz61IG7SpUzQz56aY5
Qk8a8s+q4ayx14Twz93vUQImY71CbrHRKnRU4co9jbr2lbfUkxsY5Aq/D+ztaluVjefMLrY2t89O
6HRu/KR2Blo0odWg/BccWuxR44MCI6ODpOR9W2SxCpccBttoHEP0NqZBOYroL+FUsraOALwASe1B
PqgpX2IFH112oQdg51ExwiRA6Q9rX+pFdNja39arNz1GOhMeAQ6Wc0shejFs/pnWv1v9ESwVlP+4
uZ1hYudBBaObsPWXynQY83MsK1Wf0tXn18+xLGFSju5yYzR/TrVpSiytJn04ieD4Dj3v7DnCXaj5
W3xxuNe0/yvHxGyrg4yhjlKyEDaFU9SKRljusJi8B+xZ/P0JLTiW7FLDVbYoa1iDQw7WBf2eo8xE
QEHEPa+Afb/VRGEfPCmhdxQpFUwM9ghtvYlvuTdj/CnzBh4QLd3LNJb9x0gn4CsLlSkND+GLfQ+E
ziiVHrkXu7+X3s8WyseyviAnjM0oIT6rcZslFswTfsopkWsEvRZc5As+WJcULQbLshTU3EX9xPJy
MTyWUXwmBkr2L5jf8yPWk5nEqpks9mnyGfvILnRBTRHZQUhgGZTP7mL5+h2ax4Ar230GeooHgDxT
pOvFTOzZBrDBZPPciZFaHXPlg5bJGZrH+Ks1qJFN+TptdPggU/GkuHZN0BusiQvSO3tZ+h8FjOJA
1XGFNi2ClNWx89OXhth8b4kBi1K2XRR1p8dbUmYFQikkbekvnhjcuBW0nwDJ/bNI0taVspuxsN0F
29t6r0PBIcV6uWPR9NPRfGYO950n8jrHZU96iLfrSJJohKTsYLiVtwoXhlRE6EBNeKwvrFLu9zae
nJDVequ94YxzelYtQgK1QC0t0JlmO1YDDYMnieK+N4gokG1W9KGxikK0EQCunIMYdC0YTgkfudH5
7Ph1KqEQkZS5mdMo40gtnVVANa0XA9sDFbM8/doHlLFFYZOQ0iPfFcVgyFTUout4ktN6uB+rIBGc
NVJzvkuKrwVYivToHPe/ORwZjrDkO1xttGiqb283SeM7K4GONHLNI1DaEUUFYZXlgU+/fdMqyWja
3vvy+L9jir4veit8qXJIUyriKvMvMxAEUF5SS8vPvn5lutt2fM7/GNS73jczznetyLgesYKQiGBF
v+IeeTYnsaOqe8IetQNLJ58y/Bu3qe2SAsT2FcBRlcAp+H0oxmOZcpS2Yv38mxN7Jwu3g07a9nwV
Yf+LJfGTiRQlp/75SZLvmMLjVRkTCTWwvpWHufzPY+XMLNQcJUyfvApvFztMwErMgaPbGCLn2jsV
EFuR+pcAaJ+0L40EjqjsBc2HHFK4g0zXLGhKRDIVAqS9Lt71cnJ/LzH7PnOiURuM6mOSgyA3o6Pw
MH0CqMDAklk3G8Tz691BrZetcIHK+qlSwbCUbqrOtbyBNLnev0YeTCS3weqYZecTfCE79iT+NWTc
mbltFcoOQEuYF+YsSfjTCm48lI5J3+ORzXPkYECdK3gl0oTpJv+PEj1IsffddQcGn7jJ7UeNE9/H
6yvsdrFfzHqAf6UrBTPtU0KNNJ27zIH5+MRwZ4fAWbewF4DBXJp3LTaC9JcWk/bWKsqNxZrKVlfx
l8WLjwxAPRjqYdq7MjnS2U+Rraz1HOFPGjwEXRdCnoMUcUBpE9zib07Kc26ytvzFKBteoe5PkaXc
nqXvuvW4ua4yIfgvGAQ2W8Qnecid8oVL/6tfH4hlbYLDDUSZJUWKmJL8Dp99wXF28+Ia3ggjvXxN
7k9DWwhp4e9k+F/Bsa3Gp55A+dTASg/vpbGYTAUWPef3f/hBQhkfZIcYHE8HtmlxiYu5arBtq5D7
lTt4Guqqz76Zlin2C8RnNV5IrOaWknuv7Hjakv2GD/1gpWHIMEKZVQgVuCQaclghWD0bVduhCGgg
eywPuB/1LU0KrLgZVNXGjnI3jyaU2CZmvOWGfik57e5A+k8DIThttJFB3+u94lxpomeKauI5jxF0
DTo4iI8e1FJlwQc0r2opRHeP872Zhmv8Pj/Z9xxv7gwkfBgyvipBU3HEp7C154eL7QREG2+H9lvL
/sj6+qVTBxjYv9cX7EbtTlnfzz/IV3cqf+CbdbkYF9wGUc9GWfxRNh/4oTMFHyc/m0oIeNz9gza4
onqHpjnLe3CkM4t/85Lc9MIkNoko8BuNqG85SSNjsqNtBGM7Dnx6YHqo7H3mzsAW7HC8rbHn+QhM
gjkX7kZ6qMgfRA7Ke9pWsxRrJgolIV2sytotamsk9OqTkJ7jRJ25Zm36tjG35cex13TTd9SH3wnk
DSoXbIwo2IjuyGrZULygXf14LQaY75LVQGMuxTli6KUkpGTZMmzBiGnOu13Ayx82sp1Uo4R6Ej87
8u+kufxjR5+yqU/RipAt3xTY8+w2sWY0kAfw8oPyp7AoecTMv8fbShlPZr9sOoEW9N37dGYCyU6u
CtVLV6rRvsfjFaRbKXJjxNSfN1mjUFw1sTLI2m8SK5WJZ7SGV8SpChvDpGUlddQ1UQpA+mX1vtLo
AYu8CES8HTytrm2t97Fe4+KHHGMSRc0O0SDBxOjptX/pdZ56Wa44+MTZNtGJraEEUOEJ614vloJi
my3EUhk8K0jmC+9er11eJQB8Fc6wUtTGeISC0lpIWf4JMH6NZPwMt96iGaVcGwBTMySl5Z87CLf+
iNACft9K0QYKpBsQdvc9AppjWtBC5toC7g2j5z0sPoPmn98yCLSc+weaNS24Acme9wmpN2aJgcG9
e978lTzilkKjjN5KNyyw76uzvMZAxQT1apFNNiH+oVGrBRlvTGvbYjvrYsDmlwsL6fY4iG1n87EZ
LcDFzQrCtm9hnFjtqy00VRnt5iLHtztGpEq5JXDQ/CrmgoKdDpbqEKLbXlwaNTWEk2bbrtzCtKhE
BP08PrrfMFGet9jX6PDoPASYaFfq8tg0xE+d3mKRhCGoetOOrH4Kwvd3JCYWUMhJuPnjtavRbwbk
+2uKIIAPIslx+7mojwuNv3xMppd39Lb354xAwIoo0PnbS0IDY9DG3ww9W8++NaKzr4x3A1+Sg5Xi
/+j5JXVMS+D3g7XziH+8IvW06ML8Eg5IxT+bRoYWkpfO1fl54OVC71qG4ZyeuaK/i6DvP0QO0HgJ
Ot38LZuaudzdEcp4xXas6ZWYDkjCpmq9e5lSeulRISQwkOVmoeq204VnmY9TPpCRmmzUKMP+xTN+
0Y7gTK5hbef6bzKHOsbsNFzPJw4vcEQ1YaiTvxZGrrXfFCR7uDS+tUB1e//QIY/obEyNyOro9n3F
r/V64ANvkgMd+dzDION5RQtaTOgOBCvFtkyqFJ0KnhERhdRnd/NQFpvj5iXMip2D8iTyZ8Z9QowJ
Hvt/bN5sj+4h1gQ8K3XiRuE8knLv+jc+T3Pc0OhiWLYQ9zM2dPwIP44rBwcv1BNA6cHv8ZuvhGs0
7T8eawcS+Z7fTD+023P16v9igY57WpTzaYhXktrKMFFjgaLTCr5x7Xo0LNGtayCLQwhUVwiE68ZE
aggEhuCe5qHirkMekjyRkpXj149tI0u/hyixUkkjzmZV1unEVC1yXsuB5hcrIxQdDvo2ZSEh4fC0
OmtdA2wT0lTt+NMV3d/NcNQwzzMhlIN4iOctkzX+fEtD7Swj34xHRw+HA93nDvbrcSutS08RV93c
hOCMoSGuAJNHqH53W83ivPwChmtpgFTdEI9zOpIO5lRJkJSEF92nbYPm621S4Wi9BfWJKFLUQ35k
L9kqwLWRz6XmH3EN3xNl7PnQ5erfg71nt8MrI55ARNoPGfEFIlJ2KNYj1twvI+oJs3/gtqegN/rh
ogr6kdlIEyhA9NCllNWrZdKoFCy1QetsIqGII8s6iTsASOEaixAVObX2AVpY3TTn3N2ULlmD6lms
74rQe+VOWySRqreqmGJl79PjAtvW8Y/l53g0JfyWhdWkhriZhtQNIJNk2/a+ZhcFvv9ESowNTCgP
oJxs0AWq/XZjQlqVOwCDEY7g+a4/r6rsZ8OYI27iEDdKQv7aUncePE/l9cF+Mm+37BNKwLh8rc0Y
O/KutnSEYMKtj4DGwrLMpavgXtEaRG1zRKLvDRJUseiC032c+h+6LhHl4f6MJWxFtd485ytsIwJH
LTfUC1tty/+KceYk+2DcDtGTZkxSE07q3VykTWCuu9KVU6wxbwRGJX5JCglA/Y4FvFbAv7ajZ9Wp
5FpctyYAiAvXt3IK6g9bMp+ThrVKpBMOGbPHGzHNTns9/P5VukzwMFsYNljXXHqog+sl82d90qln
23ep2JIdDRvkB0v72dg1eEdbkAUy1+IB1Z2e9VGtGzyvS+wIXh58abB4v5jdP7BdHcnM2jIUb2Z4
Q23DPxTUj7TWBi/9zACcXTbkDUhsaxoODR+IM92VQfcPV+c3RBgMhwoVJqPVBhEb3qedWUFbd+Ug
oQj56N1UeddXTvcZXxAjN7h8eGkuHm3CAv6cmbJgLFFc8jcHEMCkIdxEajTrCghTr8YDyyLC9p88
ieG6t3Nhyl9tIbD6VmVigg+cJdY9wSyih4aN04qWJpVB3Qgo3+mAJ/WGefiY1yFxvD52qDSiPAzZ
TO0LvAp5rEGb+la0ARIrk+vMwgtWKMpYLQj+Mu96wzGLk2oo/s1dqK39udiqNLQgC+giV8ss1okN
FghQP45r3Nr/OGO8/t/r9nJCtjQ4cEqg+7Q3TUO0cjq91SPhEQAeaAg04CSmfOmnrONuzZf1IG7l
FaOfkE/WC6Ti5+3VeFbkv/RKP+rvJa0BPVvxZxJ9G1kqjaY+W4RCniIh52xwe3LqGsvchOsUl4B9
Zo7hiwQ0s2QG8lHUkLOayNA2c+431vkoJ7BRUTsGd+gdoE6PeQMxBbf5HObS6BHjm2GsWUpcd8qC
Sc88oZINFlYw1B7N57KkrXv7u1b5ZCAtfeh7EO1AMJNHIrOMMk0v9mAIAR3IGJFKFXzEEcvvhw6N
2LpfNEA6Yug3osWm6Iummar5kW8hq4KUvHpKEpMoIPWtMEFYugmRGt8qovIinmwUnu3I+ybT3/SD
sziNHeGBNihihcTieOnzgJOgIPxK1+2NXjlGTS7OZLPuDHpmwXg7AnBjbR8sPhcGw1mOXCFms6IH
h4CkudTLmWM5PyfK7KPZoZ8bZSd0y+bVOGDrslSxpgZ7D1COC3pTQlw2OyJWT0e44wZBYX/5e4Sb
qlRPpfr4goBCN8QBSjWLauiw/jRO1FPqBDi7+SI/Y7Jz7Tw8HqDV36DRWLx9mpKs/Jc9g6AP5q1w
ESXncgvZ3XWVEk25QTguiOVMAydVL9Ka8m0wSExNZoFFntDnmJagisrEj3GO8Tx0j6UoAoYcrnFX
bB6Q9ZXtGim9NzPvzPGgTBBV8pa/KlNqnT+wz9TNWeL8Ca+a95OuC3MIin4v5JN7743g4BVFMnb8
nQ4fNLhZE8LMr+eBOrAUd241+qcYG72jlnfT//ufIalNg/I0tG4HGwhEkwpM3BlH7INYhvtZBuvz
aITXGCTq1zQQSk4wpr6px/NiWM4BP6l63nHqcOwlvjBbXuuTXBixaQ8/COkOoROHgbiQ0enOWV76
+UP1/4S8eii6iCG6bf68UZfoyCS9Re3FBqjAcFDp2nuq8U3PW9enC1gohQ+X+rnvL8RKV3nwGIFQ
SCdvfg2Z4xAHGTwYsEeRDlmh/Hb2KmQOUNTmOso8hxebXBxjtcPX4UFpV1XVmRcvQAfjVWlF++zy
L9OCOddHhP4d0Xx07+of0YLcj8m1ADEu12OPiKLJdLp5l0Bx6Hx+4ZSzPobjRJLSTPH9HiKOcSjf
mNshrVdaNvfVbm5DQQI8WScxkMmz2nV8g1niJg+as0FnG/1y1BeJyIKDfgJM3cwkk55Dl6v0DcA+
hDWJJO7R31ISC5GrnJZy2d2q+wVX5IGBW3WF1Qplqys22yz1FXiUyFlak33VuDd1EmB6yU6Ne3ln
PqEAX0Pj9e6iz70tgue/MCoaK4tzcCSaWUsRPGIs+fPlKJsXXcQqKJsLxmmhmZ0O80sgH5Hrp14O
HEUvl10mdfOCY8hndkRxzJFmxghXA2JKPn1qG0JybZyBNuK+LDoRyVnyExzLfTzh11EitgRURBDj
Q7m8UB2U7dEpol+kyOleFqfzotHiywwEvTxQx9quDjyRo2iJSL9XjTTa2vk+MXmcGfU7YO+rtw+y
J3kDzDDiQeNKA2nVlrldfpofUqjQDjGvJkZjH7ljzAgG41cQtP7v59/KrxoylthuaZM6cT4HSsUX
AMfaujG4mKjgIpP0SWlN8oBKSiwTL3I/gB32i5mFZhrTUhpc/iNFOBCCfxMdx28rDBp5fbLKCLa9
OfbSwgzPiNJc7CN6r2fs8BSFSxe4B0T7pBofnkAjgf/shSYQYJ4aPjfNEsncDlLWNe2ailDIv4L0
30iBk2c7HUxSeKE9RJf9xbubci9Un5Wp/qL+mcAORH/P49wKQ7k0tV+YG8vy5o+l+ApV88x7R4+K
3dnOls9A7m5kSH5ta45c+iAIZ9r7Y2Q5+B0lMa7dmHcclSzBcxqoPlUa5Fx1t8OEuwlgTmzu7jya
qHL+l4rBD4CxM+IyGe8NnwmjQr9XdZTHCfmrFvkCxisqPOhA3qQlohf298ZcyXD+Z6yMg3kRfIC9
E3H+5gwFwqZA27wMKBiy0mB8/FgxjhgFVdUs4QvM6KLctHZVaBCOij9QCq22A6WuWQT2YveTXWGL
MHBQpA8Qx/9fi5JekIkDUed5/8zjQOCB+OlRMhTrzpFU1s+UxXmjpJXXigR4V5Ac2FeCHWe6zRW8
HKzkeXNCCrK6lzguo/2XlOlmhDd8l6Y1penOzEA9S9zcQoJPW8UIAM7gaHQO89FsJNJ0E/xHiH5M
mnUpIMvjrqN/oky06mH/1+mM3DyCQ+sH43AwOO3vd2si1wg2QB3LCFSyKak3Uay5ltf/ygto0Oov
P+p7fP5brHQ8f+Vy9+4bJd/vTQMBTN+SjGZDdEsVdMsKxWmJ3+CxXHnxwr1I3H+qYYhYlAxngYM5
h8fhDqL2Sav9n0GpBx/ZB3ARskn5XfdzzNPv3A9NX5QeOnR8D/mwn6t9HlDBIkR//4H6lJJw/d7L
x2mHykl9qeztx+ishf6Ndl2mfvz0flzyPI+UQjHHCoSIonlI2rqv5uRLcf9RV+vltbRmOnrTAVQv
CUpoozzitoNPvUHWs8CVPTFzMY0tJ1M1pIN3hQ8ClNrNIzCl5n4G5e3a04E2Isd+RrD/i/X24gnP
7EY4S0kBBjcUlZzMM8GJlI0JWQNy/SC5vfsKP125yeciQjnkD5TW71O1C/R5wntckO6flrvpLW7f
lDUyQY9TBFKeHZeVRrohiXfPXUAHu4P1DvkE7jhULSlhek+R4itOueSC3nWOAOOlBYmdfm5wWn1M
Vg9w/UQKavZqSSROqwRFJCCyDxAjCihCb/mjm7i75JL6WUe9HYlrilQmJarXGVBCJMKIUIpaW5/U
4nwFLJ9M+tlUdmm5YNgLtdHBAWEW4mFbtxJnT7jFfI3UHjiBovssQyfE6/Ml7nCXL4Qty+tWfOrQ
vyDBtbw/u50Q3Kczy4yFFmZle6bFcKuXMh232DPEHV63wY3CqR/my2Uf1Hau++/g2IM9iPrLSCwr
LrXqapfJGhuvPNLg7y+gFExnP6A3qwwIayBKe7ZeGhCwYnKvOvxIyqdviv3qpiast0+mjca4P9tP
ybbqOFVIqYpTRTDqfYg+hq4rTu0ns/0b9f/+HMr3B4DZl8CpcWNPMuVbSCQ0jw/9lsu167yynCkw
uYtj5Xt4IB7QWYHy1prOzNXyNrWHcRcmeMI6SVGoqo67gaCqSKmE0R+vcTczU3qiKlEIUSc2+P+q
v5Cz33NFm8LRqH6od0nFNgIKw1iIQijNqCnvOYwoK3rlH/ETukBOgTSxR5UPK6LTTc0Fzs4aG3t2
HatJxQVPLCS7C8ayo1DfKA1iCEidyinmozLINIWyUE0prjxlZH92TDnbWEs/iyEH6XQ1507l9NnG
cRiEs1pfEjGvngTDHoXtJSPXUVy45BJHmmxdNUlr7Q2vwHH9pxyFsprPi01tN0wZ6XqHq9Qpq+7S
YPyk126hKBBmhK87l8Rt1WVGoJd//5bmOUAPMS0Q/YXHhwABBwFnBIADx6mCxpix3MsERbl3VTHh
YFXdXaT+StLjkYkIJZeT88Vnuavf+VRqzhbWbQYqdOjLK0WhAFnlICxQwx0oe+Bit5J65smDGt+d
OYtyeD3Na5ddOevTJE+1LOXhi1NQ+bX07tWAEAOx1EGctkbDrnPJpTOC2hKBmO/HBwSkUU9zfdl3
UeLvyHfBuKBLePwhKCEUO8D7SS3kcK8ZooviT8G3mwOs578TVu7+L8IfQu1lyJ1mrelg6goChtKD
ftYuaPk8j1w0dTAfMxnrZCQcUqWVaZQkLHQZGx0mdACAvb94fCoa35W9+Burc5pTyYjqOEWpkPxl
UJTKP++Qtzr7V/+/Dmo93kHAND6BWJSd39YYsZyTvd4tg3z4MAbw7rE8Cs52TO0WcvfihWJ8oK8f
gn1JJhCnN6tRbrAaD2d5d5CgEmurh0J+oTjlpJfH4bRKjUbLKNgHVL2wDHS2CMepAYZQWVsqso4t
94M8Oy44e0uBJ51BchiCA+bLhy5HfyE19MwF10Zt5xz/gTj1avaVvw+XtnlDxzTOHIFB9mOlA5g9
sm6En4yAPg7oQeqN7/zZPtpU0DqVqQSHjIKtpek7b3wmmJ788Do2aydv7RtJ4Z7ri6HhFpIkVNb2
2bHsJ2mGLGe45VC+859wxRzELgrjnykzfS0K04qmynQu6Z72RcLLewuBA3RUAo9fLznJY89H1EkU
LpH3OLbYsSW/8ypE+3cQ94KjjDjbJ12UP+4l/zRSvgNnUfIdnismu/8XMBCY0y431uTw+TqQI548
nq4L+2q7gGX7zSIwX2g2G2FvrbPf2QJPVkaf6YOF/om2XaESHoT0lJ7DteJAIymx/hFY8utFQG4Z
M5w2FKiZoN//Q4bKfkKl/9kUH2+uuMjXc2xpg5ammTCRvDUaSa3dxFtkLVQVs80ETIxlOfqokEWS
G6NE4zAAdhjLyQK1x51prUsK7+wZYnzExqoEZ3MMGSVSh1PFk2vSbYX9JDska9JlgX7WN1X3HFLo
DklrHo0FV03wUETboQd1YB8A2t+dc43imm0IGuOedwt6sgfXcNN7V4ntW/3MOe1J822WGuqi7LKe
nt6YdAaMO422D1f+u84DmL4EGe+DXM/1dBAwIRD0VAqst8Mc7XuUb+AgiwOd0WVpY5pgIWA1hdk3
OJz7+R6O1NkuvVx0bq0p9b5gMJ196lVlfVH91WaAg9EtxYfWHcPvbVNz0QDmE+upCf3tzQ/el809
kQ1FvbkPm76wPlStfdzQMsITAlUVt76vLfd+PG/HsZGfj7SdEL+xsQsMJI/s8/hEm6xQWhlE/CtP
ovMRbaNPol412cuSuAHvcdU36KM9OVDCDFvsKzK6RtRXyBmFsC26nkYRj9+MPRMK/osfG8pjtcuM
al6sThvCuzek6X+Z6ZBmEHXRgisI5Hkbat0qsC4uVBVSsBD7rNUqZSM9vWIEkQZsLhQSso13fwvF
rHTHLKmX61uV46l6dEeRtpe9P0nny7oauakoq3+SNSEN9Hi5GgakUT8kgiy25H73p+CG8oC69UIY
pEOhm/oKhuNSilT0FBW7HKfiQYWHD6DTmG/K9QoFrxJjH+nr7EYJtM1RJ3wGiNxo6X7bSz2zNfCy
l2cn9fc5TauBc1U+XAr8QR4Vun0IRcRg1hjKhMjo6Sfyug1DQ0jKXWqkOB71KA0EsQr0RfvBn2uU
dMc0nhjr9VsM3+WIGtRwrARq0faPPO6xMpY7HqqU6bQNPVKKFhRvxh0Rnsro9kg9xI4jYgkJexyF
8d95ZRTQawBHJ6u5ux4v/vY/g+mXV/yyi4Q6kb2bP9AVKfjqBDJs9GCWl8lfvpyoXp7LIsubTKF6
neEAt98AKQsKTd9qrRseM3xMnep4m2peC3xPgLuyK08ziyDC3JEnS7cbS0YHFFDey1659fKF2xNO
BMT3gJfvtaXHIlQLsl/cHeEjFKfiWmMKej2mtzV53jTjd08zrryxtRBsKrH3AQ9kNz3G4kp9Z5lT
MfugXVNOGBoB/xhkatkW7B7vFMD50jyYoda9VMhPzqkfs1CFetLEbdNgM6TXW1eGLWP6tmmygIA2
rxNI7A3NQXBa3Uk3H5EzDQYD4vjHCxAMz0JSFasPcu8v4XBSv5XfceIq1+3uoLiAfNEXNlghdrj8
YqmGJbzcPC+6oz+xbCqangxS2vllrqYSUpX3zOg976FrFB2jV2XuaRVuIF1TBblaDNUi6Y5OqG6L
hFnjVUjyN7P09EkDrKOBR+3xwN+PoVitaR/XBzFx1YppSWKpkCmp/stTn1glhskFT0JigMpgh8IA
Msq5aib5nAh6vGdRf7hKN7be6iuynvJjM0U4TcackIemEdQukZwdiiZ+jFAFqTCu3smvm+cB/iLG
0pfG9RcKDTV2wOCWBiDPWutyWoOz9FjN52Qhq/HZ/JNLqdjbKpN1PHyOesRHtZA+JIIsVBzF6Oxk
I8GgGdYKBYZrh6+gbj4mmSmzfLhTxksO/tcAAHxY86iTCHM4X8Twnni4DQaIvxpR3wAu99HqM1NQ
L++Vg1bGj2gcR+9hbFwIfKtNijgKLMuQGlhGWdvhaaTnMm9LrFxhoPF/kSo2+wDwgYpAphZ795ZY
I0EfFcAoIceoibLoCMWBrXLW0jQV5KHAz/iIQpzL3S2Fx7F1qK2TahBuciiSref7I5ZE2esCUAYU
P7rso9z3+Kk/iyYc4JiSGJyTNG9qU4qwtoMHuBckjxe3w64lkhQq0FlYX2H6Ek8P+Ug16RQHNw7I
Xa3XQ/6QixTJzwo8nEmTSTH6hoJM5tl75YmGBu0sAkGsClrEpZzDzaeWv0svtEQI2FM2mhzAdDLx
cA/wrXYxZmfJvNk40r1ylp/6HoAuuRkf4APKg7n+S1tJHRWiW9HUAhOPO4n52apGcNK3CYcpoP+9
cLF6QKuoIB2xNwWxduTCmFB9lxBMRiwF3hRiVE7AfhpUL5eRR4+rRfifSaGWo1/5yBOKpR+eNLRL
shmR+fGFHII2RaEmS+4WDe00dufG+FQF7SbApaq8lpdp3XYCZhVyHF2Ix8B2ROkmd3IPy/bsZ+Sr
fnrMdO4dnD8Y+UpPAzYDIAEyj1YQITEikz0zSMYih85eXz1o7Dx52K9NuG5tFuW6uc+14YAWF5dl
BGkmJcxYG+EtoAgmF2RlucU+LVPO93S7zqXxosyKczkevAQpO/n5f/k6bod7mcRKbvuMzkSH2WY7
njW59Ujg5DKki8RWJZd1bH2faOkvhsxfboIi+4VvIcu+jZw+sOjMbcGRIh0/PHakr03odwU+z+RZ
cHeu+aegvgYhpBlU/9Cu9ZLB0wSnrQYBGc4g3EYl2+1wTdzPQjs7nIpX8h4n+q/uYe192ZsAtj6f
tqLgonQ65Iqxzxg+RF8ttE33tI3nEAu+yRBT/+B1Nn1ZzQiyXWWqVX1/dOsyG85X8SCUmlY39hcg
LnyukHdMOODkXI+M+4/N8yjJdllXG/vHzn306QPU2EbDB2/yCQmvvmEnQVc8QQuf/6gMxXFPnvbQ
OodeTq0h8aImhO8Biyy9QzTIZD/TWj49/fET2rlivhW/ra3id5AqAov+VsU4THLShss8jkgahyUA
Kc4OBJt1IASTiFJAiJ5dUmKkCLlgJOIbbVf2Bt0CDDICfxKrrpI6KeuXR8OS+3E7TehUU2iA4cdb
Cb7ITYNiS5TXgMt0chaCdvA8TcoI3uExeDzdbIJA0W1/G/M1+LkOjTmz30/vh5//sIWyVN0peYN/
jMocLLTg6L8QygO065O0o+Idc8LAPN+Kr0qMW97S3Pwca/56eka1owfVo1+Ej9xDElGalhiKXMBY
1kcXk6Ooj7dIiLb8DvGqvAKg4+9fAj+x5FeuTVeKXm6NdsrJ9vUbna7Yp9v2iHDkAplOa9fQ8UST
Z4YYAyXAdu5k+T8MWfa7If2dV90bD69cqsRkIAcw0lHYjDPdsGxd7nkbpbUc7DdGX8pVZSL+tsYz
MwyMVHo8hIh72hUAyNHDxa8hQARJZ2ygaEiX21rM1O4BhQkGvg4ecxVf2iZJUplbjbqgZxOpNkvB
pKTe9J3bxVqKfIyjtqAknfrFm6s21HoqhGbdqHC//CYCDVTV2saF3QjmlK5we0RENe5A7xJSZjBc
UxxAvfAkztKWvU3+I2bvWhtZvXkOoBOSVOHm/if8vswgn7Aqusl+pB4j5Y0t8ZjWc/HhRg7c8o10
KJvndXpx1DiGTVqqpHMCHU3nTlGmyBpKgilIdvdzLq79ySvjqW92SYQbXgN/ZtQ6ZqFxuhrRXeKi
YCgb+eqeVIn8nEoULN3cL6nQAV6/oRm34I1NxJp66v2x8tTMeu5t41GzUa9jkK0r9hT9MMJScgO6
/THRRIpBKU2fvnBj/uvOkC2Gz2+kpCK8N7h9uyCzOjwzuqVXgR6YMnhEWzNyaXWku6dPgDRSfidp
agJwW0wYka/oz/KSDkvD9/uO3Q1XBLPNHilThkAb5MhK6rRgPdGWH9mWdyE+BHwU2qGKQk4pecZo
5mzwlmpPJ1Z+vn3nM6f+hQMp4ve8NDUaopG02hV3YdGk/uOZbxrjVajbplAlGJLFNNudp4CFbNRj
ZmuviX+KEuuCFqoMg7EnipQCwuUdW5yUgG3qWubllL5iG4TCgrOxg/92qin+vToHdYR64s0hXJ9d
OdiWEBDD6iXcB68g+QFvvS3qD/ga4sU9IJzhQeSifSfNuITtFgKsotqjBatV7DLg4hvjp/cMnaq8
xSVztJTcirKglFdGsRhhXivSAJ4RYuA263jN8CjyaDX5uFQWG1BVJMOeQ/KG3pBTSgdqI+OqgvI8
R2UeDJA7EOsENOhrcWx48MU2kBCzDI9jtrsETZs+uydQyYTOADLeg5lrOSpSgFWzihK9/ewjX6tC
EXKiFinxOMqNtzmmBT/ovNu3Ss22MgP0gVKaD6mGjZ7tzWlTf5G4gzKpsYEcZxfU7yeRjaXi2gev
Q5XLltqgX3CB5vOmLz0RIdZzLlhH4L7nha/VdN2dU6FJuZk6+I5NIIEMK+HsPsiwMiMaoFYVhgIs
9O5vjQCHSl/Rp2Z/96o3lLuU7yY84/+uNXotRt7KpIyefnLhkcD7n0cvxFCisqlJCWycnw2Y/ouC
FExUK4hxRwEZhnx2dWxXIyqrhC3xtn3m7jnoL6aUWRT4A51yOcwdQ8B4gs2FTe8S6gsLZli/4D4I
1LgV3LjsNfAvq04R/jfdqY94TMJUxOMihYyqm8lV84WWRGgSre1wcxZXpMnV4lt4VDwmwug9P+8Y
Bk1PguRLYml0cBG1jSwZZTqlD7zQKFX+OBSXGrnT4nNKCXMwYfdhZasKR/fybtSDJNM9+jhnxPrt
Df2rU0HgKFQJPp/Rby4UfzYdhv5j9XXFoSkfEgp7E8puqIgzsac6hV6gpN0XRX0HvxqkR1So4d4w
aVXSg6iOhz8RmHPV5Uc/dP64R5li6sTTxZ5l2D5eX4Kua10y0tdUFUfPae/0JXt84v2UdVz9Pvzn
o9cFLQkqJH2w0dM3PeGRreg3lou6pmMoRaGGuHbs1QWcBL5m07EoMgXuSmSCiJet1oPCr61tOKBQ
fYcjxsR/Byp5m/MtKDyIJdSOEPnyzKk8H/9hL47rFAtlo7WuxlfdUxML7VDUdZ8iKnrgYO+ytZhX
tn36UoTBvqIXS38Nw0W5LafwKCPbHubx3/KugR6euOnFenosa3Os4eJAMzmgpDVSiuElxmVQzNuo
qabKeVHeycrDFxk56YIIelc6N+1bjD3CbQbxl/tnGZqXEyunrf2kvdeAxiygOKC3l4PQQdnQkhbE
a+8Xee9e15zr+SbzkP2joXA3tXfw7paUisPjsZMwfOpZCAsYir30eFy6w10bpkeuv3bGIwQTgPLV
XEIRb/o4EyJxDYjnzrfpboYIRH92YifSEDk4WcWJLLyELIPfDxw/wNPDBEps5ZeWKCwhKd1UreFA
SERfDdVWVUBqaUcisKAevoloX6BiCu0vC06MA0gfnkI26Iqi7gKj0Gu8vYCkMVUEEOeCicoOjclW
/hiplJuupkCf3TEgwya0qHV3KJsjaODrXYvat/TF5rzk+COUJI3CnBXbd/l96pBgj2m4ezkev4vY
XdMR9DjJuTHkXv5Ps38TBWB0oJebM0cedDO5a9qxyyn//t5axDkjkYGBTVsY/eoIAfDopHnO8DZs
g4f1AhTwWs+gLx2SKvdHhmCMlMRbedsMFPs/X7IhCKvY4ySf2sZ4u7QdjKTw1q9PwrF1rIuJVjbV
fsJRClnP6S9kNYOiqVQoSDhlWOzKl0H1byhGfwIU3g6h/qPuwTen/1D+Cq6kkRoRGXj48irnfv1Z
KYCe5oImmDB5iH9GDmKryDM+VliDIeYQVDyED3S4w0rwu8BXFMOi234FBt+3u8enJWVq13FqZ0ZM
szwHt2ZOpn467FOvYhyFHmbYuQyiifWl4HbzHTpCHWBLsLKk3S8tXtXN6l2IRZ2GBb71Pj8rtqIs
XPwvThoiR2zfFcGIntp7p2XAiZg0zkRQF+oilsxiQQDbRXidca+ZvMeXApu9KslyAgOHUFvU9H6/
1i8MW0w56Rhazvw3hrufM1wBqCPCddJChsWuXnoL2cZCS+N+qOPAGn1tElCZPgrnFsypCpwubyrS
mxRLilVcze5MFST0UD57i1FZPwra1iRzSXAmm+3q7mV/cJalREBANpqHqcSdvtnnwlUvrXkmH6UK
oislWzu7u76h1xu+AMad1DtvfSJVy5BEN3HoBBil+nDfIHrKD21MxWnFjbplDmPJryBHyw79rfzw
jIqfTEMhdT+yNpw095GYo/oPFCSNAFe5Ybrk5DCS7oBIHRv3/r/q1PvKUGIz01rrjHUGNskeK5Nt
4E/WkrdcSoii67QXhSflrXpwuoAPaUAz3ef4C/lt9oTQ06z6bcj3AzFBfkplCfTF5WHBYyFW8Xkl
OncC4o3Ck74nrBUd6+vkFI0JHmDiw6Pp2zxU7ILtilxwosamATugY7Lan22dzw/BbxD5XawFx70R
dRZgN3NEOMrzeuIJpAVxA/wmSfhicqx0WVkUp90k05kAvajky9rJ0CoPVPWwgQyaEVF3DZi8XNkh
stLwZwQO+KyLnEHF1nC39rTws6nZEm9/5+T0MNvTw2JV13GsKa6fBIZNMo4kYgO/basXxrahnwf2
dh6xH2eU62TN0hXEj0jSeTqHz+pXZ9MVrneLfpyU8SR40uO6KQBZksfEA7ExtxAdVVSb7ICvMOi3
lO+4An+z/Ziw+VsHR0/gJ4a/jiTIXPC2IisicJVhQK4B5jo/oiPXERloVyOgxUh6kmE7WiLivwxX
MWahkodlHQARVckGH0h9G53ZZKl+Th26aPK1zSlwKpJCndUCeN0kyFKPAmRHzu6YLxetGe0fRpMh
8dgSihCvNDZezryw8JuFE8A3LEfO8Vovj7ciUxEa5A8GqXotMjIFDwop0Hu0nSy+QfY0/6RpJk5h
K/gWO+W76QjYmGTCpqKJNrA3fTpaBFyX+UwDfszrBjt4TQ3YNUN3CuE0ispxiISfB/hWlsgzBRcQ
Du1RfXxgy3vZNFIk+k6h8wtGiMWEz7PaArH0at9bBveDeIHAZEZbOYN8TK6Xcq6UrLk7yB3+VzeI
RwIKlR0ccpM1ecoK/hMRj3vywiN0rkxfwJJ5f9BgS6IUgifATpBeCgNme/tN3ytlDuyrKVA6KiAX
1Ns+LPnyOIj7pN6milK6hJbwznST0osrbhvN5vaz5YElHOe7931CWdU2piTs7/fDhDqlKW4upTNY
YhpN7yrRWz/PM74+tPM8+0wRDX23p1FmIyOdLVxKUuZegCQ1hz3TAJ5IF0gQQBgwO8sjIubP5VHQ
FYVHJV44n/NtY5BA16jNKk+VwZmQBEvZpg1hP/qjKbYAFlYS3255/Dl2mlg4EK1E0BiOWaVG/PYT
e30g6lUHin9Zt2g7hW7bS7IW+i+LNjqYIyUp22xKnC2o3HqDWc7ZKI19LCCd5ada5mPcuulj1M5L
nh+thkTQQf9cJcmSBLXcCif9ZyhYPJ1OzBeuO641fWdGT381t0jOus3lGUvjTjhZD/sZ5Ddagtyr
tJga1WxGX4BfuuW40IvzUVfV9f6KK5OL+4MBmzwdV91pQajsZbDe2QZNgQVFeAMKudLfwV6Qzog6
P3bKTAuD1kWJinCHFG0zfBda9VsHWeiItWihn9x++nf/ad2DaIsj9sTmzZB7EfH/EohhLHgCSl6w
4m+NRwEKx0Tt4eGQlyrwR9x6Tgtlnl/3nyoBUaptN6s9yt2RSWSp4z7fAfkA2iZBYdCr1JyqjRmr
iFCqWIHz6atujCgHNAMqJXM2Cjqqovm9mQJiitoOcuqcZL+YFJVi+EhR6l5YDy5TF448V9Ofvaoo
5smwDdeYraJ6MH12doGlgFZfrOA15iUICyDY7b4Zy+KQ8QSCTdeKo7Atv9SMOaqaoweI6p3rAWwZ
5MjKbz1qJj/qLAxx6450uxYHAkr4uMw4FzW5dtR4cAGo6xgJWQL7rUuqckeQtIoOGPTvEYkZIXw0
b/KetnyZjf35z/gVwCXxPTB8oYPI/QGxL6uoRXFg0e4r5ek5MS4igrwKkNFCzBATlD3wn41g03uB
aEa+TLgC/r6w37QiVStU2ng8tObtMnCg4tXOoUnkK99pniil8xdedZe+jRsmoqmxCSlgUmZQkTw/
2Ln5LVldU2ixs5onuuP8Fdc4dgUDiq7qj6e3DffexZtehwXo00G4TJsXttysozOTfQnDdjulppYu
1cX8+QnfFFxgf3GE8NBBCU6D1/Bgi/I9JRt6TENrezeTXCL6erIl3laQRYWI2hzZAUfGeje3+q+7
6cunN6+hsN7yjqNJCJKB8eLg3lGXTl2oisGZPBN0nRtWNgAFagxHw9JuPdReqzkqzeq3nE1G0Jkw
zFJ3oTbChRI1vZ4m/Q11A9TnyiWwmzqvLmQgiDyyRYkqWSEBsQ8IneMdPAVcUXNJuEtN/MM8+c/L
XHEneywgsw06FTwJJS7/ctaxDLu8C8i+6+P33DU08apA3aAMcPZpO+yOIDyaurlgOgJNz6m0f9mi
69iSHkal2MemSli7riO1qN+hf8d6V+nV+AzqD6jTYYnGrpuUzjz/KfCkS6Pi2cHsq5eXyTnM9opA
PIpXVxmRqYwC8j1tAzCg7/9DMQKaN59HlN5/jpgZPbIZs0PXLQRraA3uoShbTiZb7jcfKHixsdr2
gb2T8iNLgc7vRMhTtEEjY7XRNwpwEEV3cTTxP+ClMVktN2PrZWuMsWneanDbG3yXd+sPFpymN30m
BKCUYzssHWEC6gB+e2srV7Ju9WPvJEToG6/3j6cfwOl74bXNnxIADN/KfL4i76+Om3WGtgIbZ4XX
9YsCqDRPjA8uTW7o5iWOdtG8NAm/2ld2c2H/5tLtAPxJjTQIldIhSOcIBXPb6CendH56ibDGb/zU
Dg3518zCLr/1TfNlGLiZdCvSRczGD+fWeF+3Cu49jjXVUwbd6wJHHp0JBXYGRJ0+LdkZxpnm4FLg
wPCxkwAWtK3ptmu+JNwVJ+MH5K1PeRziFW8rRuqqQGiMWIVF7lYPT/rwq6fkx+Guo/pvoVkYh3R6
B6OngTQ6T/6a+tO/iz17hBq/tTaf3dQjO31hpoHzQ6sNIV9YxwnNkHJiX8F6pZCWmtsB0CUVhsTw
3zxutrNV6y27fD6cEPR+BRYJzb3P4Oe4eLZrYVA2El7YJc2wcSEtOJa7SVsqGUsy/EfygrJMLTWm
HojhQJJz4tAjypbIzoDrF/08NwVGbXCoRwG2obifgKaQ6I+fmeu67b6jM+IZ+8wEvy/G8u5SGteQ
1K5sOhVfc2JrfD08uj/Frn4bigOSYOByP4pdRTAlDKjtkmycMN1gfy54M9dmCCPraeNptTiNViOp
LQF7ev1mNFbKiaZFCUusU0FP0swe2xmQEwd5bUyhHOpdUQTQ3Hb4HYxnp7VC3u+49wC38YSHlq+4
wM8Vha/dDjHbKsKZ0b3CuIpwO/cLv4hJorIv0pSTgWxe4qcH7Vthn7/8Ty4jM/2dUXzux+F5HaWQ
gjGRFAkkTABe0UGKJqvwDdTFp2lDTR4UXInMsrZK8CmXkhAGJ8X5/RJbVyoBjDgvpBPB5LQdx2uR
Kn8vsonBoGF7Vk8xaUGOTtnXsdKS972YOhCzgl2p+hNJgulQZ6M5/9837nNe/RssxL5CXcStKOvG
ThhHImXD038EEFfPWQzdwBdlryZINrIg14UbUL2Tr3OPqYOhKJczqvKzh3MjfWA/XRJCyf0AhxYS
DMfiUvYQq6z9beuLvlUvZ3pjx0Cj/P4kc9ng57hsMLraeb2DcOHQjZvuJ6D23UDOyGgtS+dcmUag
vBOzhLV3/D3uRccXBrOc6YXF8TrMMEd52gZBX+R3cnNhgQ7tycoDiySmocxYvs+0FPHPwu6Vb7vE
hGCkY1NxclSAd8EjuYCZM3PbJwfomMHgCxx3lY6zH6bMWw1cY13RLD1dehO24UJ4PqdJR1UyXJ0x
DGCdjDR+BRXsU572yzgLYc/8f+GfEXL4SslIEQik7ZZ2GEuv8xE1goTymUxZhHDuCSjaf0NXTUR0
SgWEaGfVOC4kohPWkdcP6giiojEILsxBDuglt7yNMW7zqaY5o5xeQu/kv3SBYfMrVJIWwvdoiDie
siQ15o+ubGz0QdMWiUjDKg8I+MmvaDxIe6HRCyWiw6bPWA8dpFoHf6rN5h3BckY8SYsN840AaFEH
j2NcuoTiAY8XWU4ujd1yWi87mRBVgrILSv/LuLY4r2xgAN/gNDtCEsscuQs5ooUoYNVx71tVRKVC
GJBo47a5hcj45L/nvzzRQLe4X7MldBgNWw2iMhfDQrmEsPFSeqz5f7DgLJ+sJyBHc5SskSSCcgw/
JBDgMqwGkhFR6Li3NRQ1fmPbjXdgXFvb3JPV9mPy4+RsT7y0L7TQIC/vruPUvAOFGd8dmve/PCqV
8T63nbO4VzAStxQ2T9ZJzI/2dVrvvBgG8xm9kWaQkcDv3CU3ZdOAJMT5U1PjVvR6Ii2x0xv44KR5
mbKE7dmRN4XlwWcZpgdhnmxDPbpQzLhhk/9ICgEBC6W+1L4+/mtZtI2o151fwv7O5QLzQqpCA8sR
b1SjAn9A0ULBP98olFQFkOUCsfTxzLlY2oM47YZTYdVDDGYjSDxU7DIANjePyEgqgs7IuH/zqOxf
s4rcRkMVVF522BisJKMwKZNm1qsPrEuKgGOJZOupcT3rouNp6/KCUK07hnhp1mUa6X3u8LKx22Hf
G/9AzjJ929wdAM4RXR9xb3pGrNXpykL7MgRapeZ2m5pjHJ5dAHSLhU0e1ADXw3PsREnLzYrmmrYD
ogJcnKK6cvGkK54CQb2w0lFMz9f/lCkQhtKfOqHqRbT2HQ93w+HGdfLLIIiaLsrVQ/Q+MbURH5pW
YSN5QM4BiHsfDtF9YHFnbPg13zn7O3yKiRk4OaZLACb9DBLKXJvL0D7tshdb81UTfoueVYx0cydm
LZE/8ApuLr5/sAeN0YDBLcGeDwLoK5aXrFc/30W0Hq7qb8iczAF+S2dd7MDzQXSNxLY2Tz5m3SR7
oAeoftH781LFalfwQLygnj1kDS6AiK57Oevo57V4hc78AgD9T3kkIEASiAR9frUNXOGs58xMq0tl
3kNkaArPdeTtCRl4SUxnfkwf6SiNkuqOqFoytVPl+XorOArDF+hmxL5baOOxTOIK6MWtW9JDt2MP
lMu7oru/LgL2QBQ2PFK3R2GDoIj1/HbvAjXaLw/AKAOPrxK1TpnbVd7t2kvFBuIQIBhT0g5j/v1+
ZslBZ1yJesHiA1HSxcxZO4QFTmYlVTcSkWvYij9Bbqg+L7UcmJ/+XkQN3jVaG25fpxO5eD57CJ64
ZyyHFLmn+Fx8aa4naPk+QOP5r1/sDz3/1ntuBBuLythSovLXwBLSa/+2WwUudUHmc9HBw+U4zaaF
cH4G9arZG8y4WCaF0IE/jEuvoJNLubEz44730hU+dzbrv6IQiGOjhJSmfyUtZhEIgSAp5jl/ONnd
zdtBjwwuZkesbofbmSw3X+HyAXJnuT+FhUwQyTyxbvVyt2H/QiEdB2swLZPHTyo/0tUA3GsNTr2s
41QYIWCy1PxXF0fVAHGjqlgeTW1u+ORybLcHHrGIcD9m+wE1usn3s6gWftYuRgbuI7WcPA/B1TR3
dRsx7Waiq5uzKdt+Oo+h2rTV6OcMWek6ndhQmP4Fo71qyyIbA2o4TXEs/eg8Ey9sbmvoC5pUOU2U
Zvukmkpwn+lrsmwZPfoiNfByBEBVuLruCd/o3pZMlZQXQUgLuJNRIwUXszJiRIaaLLJQZhN91+LT
ZI6wWg3cWdGpNmleVnfeX6yT3BmmpVKTJOu6oO7+ZYt0s8X1pB83YNv95cU14bTUJuQqQ/N8q0Dd
Jj2C3OIFaORmebF+DOaZwHAIrK+rZtXcC39OarSixIcMDZ20DRwJe3p0HgYH2rz7Z4KyyMLjSxV9
vPQjovKjKSbTv824oGF5DvfSRRGsfD/tivpt4UkNgeDyrzrg7VAklbajPoJQBfLWaO61dXezGhAa
/fU5PxUiM5sNk9A7Gc03MqtkBUpkJPifC/yWixAe4lbP4A74XXBBRsFaAtf/5J5LF2eYFl2cYlBO
l9rrfR4VaBFKBm8FD8tZ8I19RUMdPtQZTz4XPV/vtMz8n0ZL5xTLQuyL3ojruzLjJkJNJMG7G2UW
DG1A+IufXuo7kWc5YhThTQ9FG/U8UtqFqiUI5xzi3MUUG+t8y/epfuMgR7RPwvZGb+3+0e17Zz74
JGdf2uHFtQG/J1WE5amooMwhR51VAtsZrtCsRNujTY+kbQhof5NpFgZe7sn/KiyVWUOHt7qmtDQO
SJToK1TcMesTxi44hNiBjGXqCjhuFTOlNoDE+tnIZXgOt/38P5kkEuwbX1kSFHKSNZJoQp4OUmTJ
Ir3KlqIroL0Oo3bz21lzc10Fhs0jd/QpsiyLfNXlFfLAIW/Fj9L5jvlSGpEHzbks6WqJFB3Z7SpY
oyC3Xgzhr0Srl8ldkBu/ziOSaDGKRdhk6OhSE/gURghQYuXvW9bdtdlx4ft68Vd1Z1y2dYiIAfGj
xxssiuXQ0BzMcOGmfmQtaXyV5NMZQRb4/W7ichgjRGrC3w6HrFl2Mu7ONUfZoaIgdLOlIdbgZnxi
Cn1EQiYoedW9v40W31UeAm1PJYvizN9y/P8hWON7jCYw4QCIItg5MEUpUw44spUfNxkOlvs3g4N3
kJUP5plG1zSg0kTju7ns7i+ghgSbKyehi4GtKTLVqR70sMHHoko7TIQaDgudGJISU21hicDJs1RA
ctk0cjw48V3BEOuLUncKmsYRquwoBtDlimILHdW3WuFfuMSYFiUF8CjOO4Ls/36u5RGdplM+F0th
WfR1ECf/K7b+5Su6U1OkAaT+fMjkBCxkSm4VkMrO2rDx+ghm6PsS1NkvB5II8JXLITWmwYjTo056
gpCKv8xj7dyWbuWMQyCMKttNJk9Ai7sgUk3OPQ9epgC8ewcbuTA+Q7CSOu8QRIvJ6A1XIfWMdB4A
RQtWkrrZ8QwVFbejxRCuJlxC+yiOdXzC8+n0oB2jIjAxWbVT+DG/cYN0wH6QnNvWF6pPbSR4NFUy
1TNUrFbZVmj5Q3w069NjN3Qad6H0be7XbflDWUR5hSUylrmKT4dvoOzp5H1KCbQUiEnedZXX/r2d
Rx1dl4iw6rClOJy3HNIQ/XTSf3vAfFmhAaILCiOQsqa/Lvx9d1kgEEoV9vyrGtP3CSixXaLMfexv
09elHPnPLzD7636ITAauZGSPzOo4unprsonXnGmvV9wRXpqT7sEVzJnbzVtQhg70Pw47Gn03ckjY
5QcCCf5nYqnq1yhQ/R1x9KTp2e+5OjzAsZrZlrO2OYi/mVa9mNN85pHqAs6gP686JwQb6yz86Cke
hRuwYiJjTPIDqWmaZBt5YpMqu5uKUyBWVN9iGwkHnMWZBIR87dZj48ZheQr5z0lWktaTqGbmDvw7
kRdPf4/JmJKBnXnKfD0JM/dRi16HIq0wZU7NSPfa9LK0U7jeW5va0YRO98C/cO/5/LTMkHnjXTGG
D+HwPb4MFH2B9dY5hubwD55YX0txOXIddBiFJ3zo+9l+YByut1/BzVnNDU3t/oGujQf364GrF/QW
VVv8/qRJ8R0uuWVJLv/t3U24tb3IcOTMw5ohd8Ms7iKgJCIO0SzpjeNnOtPgh7bUFFiZGoviKQyM
hsy0cXQMdtIWKrbKNTuLJYZvfxTgqltnJhfIBq6lOgtV/VrSlSfFsPDpKDAcJQ80GyEG0UpInI2e
WWzKkjZDmlK8U9SZSzXTJrcfH/fHZsYuXFQSpU3NCqFI8XkrNUXlV/X/TjCPVPa96ScwR+sS1qk7
q06WiZnzOwkWN9XpxkgaW8e78Yj3ziM+O5/ik9lo24k00iEEZ3u4+hF8Rpg6uYz7gwIugvUGG677
eekcSbM9jUJrZB9dr6bRmYYRBQnDcQphk4hpf3TI0YrC1SOxOGztRX5RZ89G/ifkGyrpx8b618oi
DvLmWpzeibUP8SDcUr3zAnbjuytHNKa6G1rY1zaAB/uyklj/gI4Td7s1WGgyY2uCFdgokQE1d7Go
uvOfmsrIaaOL4AN19Q8LU6AQTEjg7a21meZo/IP7jyh8G71ZlW8d7XDY3de2cjpH22vZ4DGfM2er
VnNQfMuXQnJdwAjiBNRYkkJFqhtczS9a/BCo89Jsqao87X09smHpOcQH3R0d2fSoGeWzBO5EhWD0
B/ZoTYVuxUkEi4IjuI3HPz4N7xbCK+Il5KlkVocHlDyS0KpbxiEyJEgsNLQUSzFYOiR2Nrq+B9qP
YStu6mBfzH6Jbb4/7vAyNwxTks/k1JHdF/mN9CumjHauygQFunH1DuZLk1UH7mkW4xZI4Tn0GGej
S6noFT+6F/ywvvpbXtTaOr26wPeEuTcnYg760QHXZvD/EJaopSmUeXKV+3lF5eqywDZn3Y6MGuZh
Usn3vWDPfZDj3zLbyS4m+aG4S7tqKhpWyUnD9CP0Uu2Gd73b13NZXFwi+H06M/+ahMgxcZNGDe2A
4MeW9YGnaCXorJPAhn/Tu3gB4fTnQzMAdkWb3bsrDm8Gi0TDCz+zxoa/toVNr0tvWP5pXx4ZQVFQ
ZanZ9UenBULX468U8x2Z1wZSMd08SHlh5oQ9ebu98rVjqNxEpcvtAiaqZaA+qrztliE93eQAGhDH
xB88dQy0jE3mIrgKtw/GH0pe35UtffLFvMHhrI0bPKr63hA8aya50iB2dItKEK4s6yErTgi8goSL
K1ZtgFbwJcYpFJ2inykGFDz9EyxGffT0THIrNrbEfT2Sa8TZD0XsFA4CIRpSbzl021zJcsqSky8p
XEPTns6JWiaCeV4jNMpBe2+nFZl++jRhzOY+/ZeD2MBaZa6hc4vT7e6eS2JBe8cUKKbEH437UoRc
LPu466OZ0lpppDeSTqVtRbWQqKoQnq2uTXid1GiRBRe7GFdEGX1bQ2K3DlWgmafv+RkxExtHIKbb
pMqiPJaWAtoD3NNEwGc+HgKKrT6SyjwpOHuakmUvy1ztPcd/niKhBkHZMPrmI50lrdvchMti43VB
4vjL9buBOEc4R0/DO53jQ7J7eUtMqdnEgDfnQWxDuxcZnY46OtnxlZT2kRjRVCyCsGC+xM4MnHN5
c2TeJEe4fpTMnS5ctjSGFCcsHTisK0/fefBr+H+bQJEjmN7F4gR4y+U/9ZEvw76orIG7u37i7Nbh
wBEUNMALYBXfbjHK5OPDw7ci8hU7EOm3/NotBhfNwUB6Z1/96nc2NEs1UblRLJPhn9mj0I7wDR3r
5wmKzS+uw+9y1Ac/sOzg3MlMKxr6qXt3kWzWmaPSMtetUpnwIdrUafnzUuJMJmBpaOp/HdOEFosL
ISwWicsSZCZUXLbTnmJM/pSQ/OycZawAYbqavETSpBpE7627coNjEI/DWSrJ7le2db7KL2EkeAga
18HIEzBU+C20VQFbWqOnht3Mxheu8PjQRCbE6+aKjP576XDe8K4H3ld0DLo7LyKcsRu+rKMtULuy
O+tou05DV03ujdqT/yD2ozmFaCXhr/+U6jGDuaroxQn/K+Gd1k8VwUGP4TcZlwmZlDwjjlR+ImSx
/3S03ApDcz1KmAHyE3Lwv/zrBcwDXm8wKQu8D3k8KTZCRrwBmmYuh2oOmj6ETXE6Z6wjywpMJAEU
F0/toravS370Hew5i7gg442VBllNPLYJexLV5DtsRTNlVpQLbFkzJrL5FPZ+LEjl3gxOWKcCZvb+
DaO5NSUbEBpawpflZLj4aPaCCi/RPl6lYMtMxSm2C7pE/SBF25A/slmpx69PjNke9762gWjsdZ+o
3tG1dskXEE4811a0g0h9+F8zijHTfob88HUl05Yo+3JbVUEQc7GBHLOOFNUO666hG03q3McWnf8w
NrXVtUsgWT51wot4h76PqAq9iUA7UsNoSS0XgbBmpLULSt2GFdhM/yrZMZRDJG8Yy5C31AYtAGhs
uRRUsvaOuNTCtR5tRrjAiLlql60a3SQJJ29aIoOkzj/urDLji5oG2oXoG8sbNZd8cX2h3P5cljDG
+PsMzBk1VrCb7K1F8ven2vLsnsjkuK+3I2TVdlZcBFHox8dzulowoiYF9B/LxndGpxVuyYj/iOIq
3fhw7cJDsDg+vapODg1srPi8nGwYWNjKgQBX4e/ihGmT9HpQfHd3uBHHJ8Eoea+gRr0C1Nh3cF3i
9S8pEyKDdU5X1/wSrG29zxF4dNQdWUyyHXtiDV1zSbQYM2zzYPc1BlFPoBUzKEL68KSLPvmKQk3v
BgNKghtN/uvz1jNRqBvxlB52LWwW/qfpYWCiez4WETZXhEeP+pQHv/TTj7MQGEkIZH7KkUBTA4eU
6nNf1O2iCNRC5Sy3VOyD0xmSuu2Sm5Ik0l7h/T9lsaj2RwOOq91TpxPTzJ7z6OltF1Wa2SpxAFHi
e9qCMZfxpVQOpS7ZGC4P2XWovFx3qOYo0oViXG+eNwX03ezr5EDMEr0En3JBWbtsQaA4nu+SaqAD
K6K3IbghTlcldv6GOemkuTsMOBY9z6AcGEPYVQfj++xTLyVBfJX/PZ52laECkDw8bMYItmHmnK17
6FWysLvq9HmcXlu+NyZVUlQsIO0Ke29n4evbrtF0fieQwQR4VKEbRkrE1jWyNwb8jQJ7mPAe/eCa
Z6UwlmXuY/xqmcpsQPGGjzX7HgujiAGwLnozb0/Mf/1hyEWkd2qIvYw+ag26b/+AgZo164CW97OW
QtNknkY/a67Z1PuTjxvdIvSsTXrbJ8pvGaxtlRLN+pqdnVlB1dxkyUo1dfq40YFt4FfKLZQwmLYS
cYEfP92k3CsTxC1kRwvb2DBjDlrWtvLfErePSYlfw4jdelntyjCPQErf0G9TNH15uniuYKqO1Jzz
1paO/qD/LoCajXhHS5hUXoJEdhmhDajFZjZOrpB8lR4V/NO4GJOI3UxoCTvkb+D7KgChAnkt2GSe
OT2Nc6ZPqNTmv09lI4x/5JjxnLD5lrD5DO/qWgt8Z4sEciN0/DIl4Hjg2EHJZg4qnLVnwquHCQRj
/lGYAORImS4y6odDxE1itGOLMVXDOhbBesqcF6Ya1/08JyTRefJyPKV4oaEafMkDLBlCWmZIVrXq
ANsCACGYKfr0yPvMHcRQ0N55iez/wmhAJIwx2zQ2cOT9LdEBh22UILKIzlA5gsUCX/qpFSMUB61V
+YSv0aARcmFUA32kgU9M4Bau46wLNdN+xnxa4LMt+7/Eg2abyS6V1wkSbUFcJkoB/J108rBZQQJO
dSRAo1tDUZadqHEJnSHywLKDAgyXlZrixvmcJh9g0N+NsZ9Nl7+3V9I1u8x9UG9man8E9vAjcIvP
WQEZiwNFXb0g0EBQ9romGoii+PJzHhCXhdZSdewRGkhx5H3TDKQxfQnrd1h+nerAlAKcsP9kt5D5
bOy8RmMfPRtwiwKvsNvtk4U4oYEkX6RlGsNRT2Vnj3vv0S/lqJSkFP9jYoKdGQFydGZrDuvzMdTp
crfA8+Huri2qFNbB+P2nnS+6/uDsMRbg6LCaC5pq+/8RndWZNlH47obZq2nAA4Xe7bo1n1RyR4tF
DYmZkwiCOCEDKm7Xdfa+/6iCNOJ2iIR/hl+uIglmVMA815c5pGPN1knXVf/LvHco/blsLLYOih7j
+qIYpJlMRhNUm9gm8diXNSEQFw9Bsb65GeWYxXrKbyUYVqX8rWPm2ujK3B1FoeVuV0qOI4ke2KOS
Fuy0TqM3I/XKEt68/qXtQnMB+jUrNXmR1xOpGGyIR8g5+IsfX6Y9oS4s5yXssK1rJOsdhBhWMSMF
kbffsxmCrOALjbmRidToGmFnTyJb+s9roiFBUSw+MpDEm88bzZtW0BYYi/fQ2uBwifrPJw995qcX
UGU3PFetcUWvBdeX3KndsNdOF3dNUHqKUd/xSQQ167JKZWkuB33PWCWb2b3N159Fwgy5MDK8R8PU
v1Lla6tr46X0phLeX9L1LlskBZDHxTjQZG+tXTdH1oyJ7x0AcdjVsKte4usvR4XqmfGK5Pm7ILXM
IkntWoUFDI6p2yGmkjqR+Xg0RYkoJVrd/kYK0m8+R47p6iwyLyPEiPJWDmE+k32lDaVzd9RXX6rw
ne/znpdMQ5EnxCKMPRkGUZpXF3SHKokq/BMWjmWLmj8G959M1M+RfjSGBYps212XG6ynMlVIIfq+
w/J9Gkt+Dcu1mjnpPa9qYfIFP4smHQbOBJQfejuV4f12lociG9+BGz6fs2S16gSn3625EvIJnxdC
frEST3xAhWJRb0g2FD5h0wJjkxW7OaaGvxRceiudGANNmflxg5y1+seZ2vK+uhHsnX50Ad/tN3G0
EIoMgwtjWR+iI7g4vxApEhQqjgpgpg6c/oc36ptn6s3mMJKlYJSpC2otNk7+DTOlNVH0JLkJDgP5
WRzBUeay+q9NzYpiFBYr3+RPF9VZMlzmx+boj0zPLRiWiX0IyN4Ndc1QkNIS7NnPrZLZD7gNMSJ9
gz/D59j2StQCeA4enVELzCKvgL0zylyjv+elLUEokjxW8wqeRb1UhA90FGE3EaVx6tHFQZRQ0nQx
AQM6RRrISFR2pt1he+SXYGzoJHDYbVuEhzHKPWsQmh1xfNcGFIb0VFOjO34C4bIuFUH8TrKtNJq/
5at3uLfFDbXY8aJh37JBBBYWYMXIwf6EuQZC1l0xJUY4wFOPlX1lO760XPwLfxd1azO/X+zD+jZP
UXk28/6UOe6pUqTbg1S+BTzcPZCf30k645CqtuVKZE6Ta21LN9BlkCK8jHH9XIbI7Mt7lD7kMr3o
4S7Dxt6vBRvnRHx+m1N7MNC/Pqu7ztu4i2BCoaGplakV23DhdsTAHNCusR4kxBOkmQw3N6WB33st
+x0/URKdFzfw9Qkk8PR62wBobood1jAZurT+Zczq/OkRzxFc56EQU6DPRh++4lMs/goclMpgxiYD
fjD06F8H+Fye/anTifINSRrXS35FtDhPKjVastnGH1cxdhkQBxzG3JUI0cT4r4596CLz0VqSuGld
++LBju1Z5sKChwMbH8wWk5QefXjlpM6FBLIHtycSXKqhC0Pw9ppnMZhv58KGeyORXkAEPOAvOYRU
4Oh/7KxwWfmbOdwTBTeiwoFTfqwki5ItxXOeEXSni8Hi4leIte7Zn2+Bc9ThnjpjH3SpfpMuqUYi
zN/GQer8oD/y+eVqi4/H3aixwfSzg/67z7pjWijkNTVLTJK+BzLgRoOBgJqxobgFATfjsOPz0qW2
am03Ditw1b+B8krvg77h8+iFkChodF6VBMGTR4R0LHVURSmfnnzeJgMulHbZsPvZWuLLCR6Czeyn
PVL9FI5uhfJiO9s1PFED1asq819I3ZGbH9iDvLOtwxzYOlYD+LPiHDMB/j0sR/j+G/cHS3waXlJX
Rn4agqt3C9xsloRF4htJHHZ1OCxzxJODBaAT2qEy+H+VClcKGFSKRoBxPxOw53tN1cACc0W9Jo+I
xhTsdjLYknYz5anR9a8IxVJQqVGR4qTJzJUAI0959wWv3zWADrtwK30b+z6aSbQWh4NCKoO77lp0
CGZcWs4RLt9nCeqaVGqqntdQbgINywgXlozA8DFJwWjjLZYCvjHvB4ZL+FXjOCzAeWGx4rpB7DgO
k2jnhhYlk+kzDT2qAYUN+W0+k6eJnHC66814Qp21QaTDM4KZ00ZpWlyHe0hVPNreFDiE4U4F7kiX
WMeaEg5X1OcR2N8YEOBQtW9iBgitJplo69F5iwvn3BTtVXJEMDXaWhQPrB0EPuRsKUENO8JvpjUY
EqUf5nBqnWI/l9HVipX/4syuNC19qLTgasrF/5AyLQ8Y73kqEndWJpB0G70oKfKcGWjcJhjOS+UK
lUs+z70h1NYLDSVaXOFyOFUblWMA7cRTPFY++ZoVz0fBROBr2PniNMh3BJ+KTljC2ruFZH/hwuW0
PvO6YZGsKrsYAYaL7mNYRh0jGta+LThgh+hGhS3flstCJ8JZfC/eLvhLsCn/L+4M+/6r4SvU2HAK
4XupTIEF3ZSliqSMjQVu18LTo1oq2fV7MDCLRhxrXM+CM5wiVyyZKUPLeWYQNEn+k2WGiM5YdYu1
CW/GwHt5mTcMX6DxDMD3ZWUMTkTdqvbykOYZVxxEmPSCj99NspyjSMdF4zLlpwhpC6umxMB/alhz
qPO99WmJ8EsLz0fIotIkr01R0OZQidAYW7BHqBnRLGY0Vwx9aw10hLlc6R+ObAYmE9/+og+J3PNd
Xp4XqKE4hsaNLDbRx6v1ebn98/1o6rpxeheDnPnNlTr8M0s6TRVUWkFwaFOTNAnYl6IPwNaCPJ6y
OgdAOEm+S1moePe5UCxKFfz+4iBQ1f0lEWl9La9rBEt2wIULD4ukizqP89tr6FEjleXGvkqBxdjN
TFW7oT5ajSxihDWo8FS51Jp1ApVXkSfwcuAhIQ8xmCCYS7pSzrqOkvDPyuJ+1anFS5bRFAtm9ev2
NogQe9H8QnWayOjniiUYF3ii7Ac1YxXyAO4KyZje6VyFYJKQBIKV4A0ckizvXYPQriz9J7HDU4vr
il8bLfyzfqdKZ6A1wViEwOQ7kZY8jTFO7CK7mUzrudvhnqo95m6f39RRMvq86WvaVYviVz+TKqmi
aH0qX8iNyIUCfvgb42jaXV4ebx2/Vtn5Z9KcQvEXq/HPUQWOC71OD+smOjGvY62+gXkB+Myjrsxj
hxLh8p45wyN1TOpD/QA1ysteIUXlEty/j+vS6s0ku/+VW1laivCyKpVCJl1Bc00aZaGUbXqr2dK+
+Zqv7CfAiBETiWdata8vha625dJBnydneKGwpTM8/ygmqKOxakCmOjBfrXu5wUH6VqUIeDB8XYtu
GDjjG+HMWyIsG1+JkwY+c8pC6MttEJuHonLPuozIF4WrkRAeBoCjx6wWN5eUYtRMRhLsLh8saZfB
6qOAQM/YON26ofz5AxOrQW0gCuhIWMTrH9pBQOxaPL1zrwb3mfv0NM4mzDJ+HpRd5f7u/5yHqsJo
5BC2Ri2dVeCJ2Mbl2Jxg6HWORhzGwUMHFlbI7ZZYyIgVvZkVv08A6WkdIwlkCAMY5eeBhhhzw7ks
vWvQBw3rNYS18zOr9OlT43z1WAziFoCMUzaZ205OWKnFZGcoFSbCizpo0MBcTO5TOlNoX3C1iCd6
vqjjtKJ3UGrPEc51j+7FiWF5ulw7FxZJaKutrVO6TZB7EH684rb57K3+SWmnD9l7I+lJ5qK96N9o
pnY7Cv0CVNru2b8E8+kybjxRu+EfS/k3No2oq1kRKk0n+ZztxtDkD5pGSenrzA3jwy+SJ69XPWSk
Tq2x7Ulcs6UT+nRFpwx/Pe6YmN5yTY2s6RLefN+taU4k3UupXfY9lTklvAJTU25DjDV6En/h6zcs
yRzel0jhsE7ef+aq7NGnS5xlWXQlB3mEyhJDk343Dos6WH8VM70odEhbuFczl35xGf+mhEyCsHtA
1TZq/ICmBDHXAZKsL/R1iUnNE0v6eFOcUFNbkxjwDXrMH/NsteOvfww2JAWdPRlIFFQg5QGlX7y+
2rPRqd3RpBqv/6cq/uptM3EK3vfKnExpElKNMH0MzUIWYxPKNVUsx52XVkElJZz9oQW6lcL5XOOP
PKFCQTYUNZZfEkMZXRVYo5WYPv5wfDAnUjJD+DVDg9S2rHTPl3RFyhHn87XLYvH4+gGlGZrbF7vl
HrFS885+P/CSSYZbIlRc65AWXoShzfMs4ypD4Xkdl+VGeJTsAKIdVljc0XNjQnWDh9VXC5ZXw0uK
MdwJa1qZVEp1JtcstZQPMM1JwABmgwJyF3E77brgq6TRmuvGkf4cQBB/L/q7ndac7TYQ/zQh3kU3
0mh+jC96XgdxkiJmV96Bq9pHSOY3EJNuaBHhEhP4Axdf01FcKOVl3/5xgvrlR4QdW10FYk2b0xlL
GgIE2lb3ZR+PMcjvj41UYDOInbWmSLvHVoZXmN3w/6a/FStZVmvIC1074CDC0fAPljrcAuwiudIp
WrA8+yOWRdLO1k2XCl7nWfQ4bQaTJ9NzFjifb5dN4LYdHCKQwDwKynThKSJ2+H3+wxc9hGvr2PO2
SHc8+df8ZMGFrXjyYBbJtcUemvyNulGRsgiPnAYINywW07/1kTKTuzvy4Do1Ntu4PodSzi2MKhBs
kDleFlm2pdr7gt6B7wVp4FzxFvgYYc0sGV6aOXw6FDBeaYp5Qdjm5qiHJ7A0a44631X4ild3k/EI
VAAP9V4ZAenEkWRwJCl5Dt2X41/LN7lYwKFKGY3uz5jc6o2Ws11l1B7PGnG9bbNkXwDzYKUwQ47B
X+unjbmZKpB8qFirittZ07DNNQ/1THnktcEik1i106aT34aqGbdwkBqcjFtUeM4g0pIDBWb4tvGA
OiLnq9HmE2oMfIHGjLoxQ9JzSLK3QPIEYO+4i0zali6jIkReFBC6+5wanAG0bjNubdo/f4cYYrlk
ZGlTN8NW2SZ7r4gnvRqajwy32tAmkRB9pLDovnk+xRDXyIkkQZ2ijo3rtFJ/zcO4vn++iLuHnGp6
DxiPEXRD7E9X0xHEspc0IrDL2yqVaXsX4P6fVuVJiYiVLPelNdMW/CleCuKBNLhdDOgjT48ol88+
Ec6oxyv82Q0WQu6/oEwVJzDw/jDESyrphE7N+MFZdAjt4Fysm6eroY8lgJXAK2e0wmCC5BNMjpTo
YTqv5ZMUWMI2pWfKbOcHfS41B06/GsDfOJ5+hA+yHA6oaovXoHoG+EWvoZSLodmBCxAq/+vniJlY
mTZuw16dxcGY/68e4ZOwQ/tdbUertFn713y/YScCjAVWcBTjnw97mfG8fkVRZFaoDLjOdseofTyG
BcVw2gVPuct9qi3m0pu7Yi8TU0VyNs8kOtXoQF2rABFRnaPjEXIencjNw1KsHwRvQYsDZR2LkpBg
uhQlg6+YAQCvy7ZNWQt4sw/QW14NrgRrCEw8EmprpZUeL+bi1eHoXmXfK2UUf6NybnscLEp5LPvI
iej0BR0gXYJNbq1sDdnxKlVvSBUdtJIAMbIogUFPIXh5JpjeAbHJ2pR9z4Z720SM5EBSHvOUA0Bf
zjCZXaS9+DW9lznzj0M/QtkyRS7A5ltiLpAmJUunEmWwFwzzaFCP379FQLiC8q3oUmc22GMSR9Vx
yNKgzUNHT8eyLYeWm1B1SntjMezJMsZ7nJQghSXD05otlNtNsIbm5R26DFOXW/HRzaU+ZdJLkaCI
5Cx4UQBpzS+DZn7bxp13FIbW/p95HEIm+T6ENcQjJ3qoyXp7NYdxqnsHKsngdoLPPqazo7sjbvQr
MFBl2+noC5jPELj/Xm1MIBr+Eo11ezpjn7y4DDVyuWIh3aUyDRAqb4I3mzf5z5XoDdcozAgaYDCQ
dsnSr6XwT+EEH7IsaTeEShaM4637H8d41UVpW/ieVgqSK8zaSsaa6eB4yXzvBtjE58jdegLcPLAu
518/mTK+NcxmFe3uS6rIm7KW1GzKKzAWqBz7/GEHYmX7TpXWuzWztDnnMsQeJOJrrKjAUUjG8twl
Tmu/5s2m9FDgUo8qqCMX2f+wGx7yDYy3Fd/Fr83RYtrfKc4ndGrDW0ac0+HSEWXZxPdX0TCtbhVG
ONZ//CiGOn2sVBqeIUaT4tp/8mzjRuMGJh6QDExYMJAHFjVoJNWsMb1UOyfUsPJIHcoJfKI53x13
OFIQGcxrwjHIZGS/Dgf3e/23m3bh12kSgucl5PvVG3h1W+LruvZR6Ws/xm+UyAo+KlakVJuqSr2M
LHgwUzMyvRb8d0p6fhSE5nzuRMsQicMa5WVZU39nVK5ug13Jep0aXcRVZCO76jsP/1fj0eYw9p5i
xWtfFq4aexy9ySkNdHzf4F386Xvc6RJEJj+bQ2oR2CDkDGz+xA25z+MLyMy0fzbXweI8YgbHwWUF
tY4F3hotzjLPz9bgZH+MLWnySLz9sCoheAd0QpP8QaErKYmLnOBgK7jAruvu9iNU6AXUaeTjN6m3
j+dh7r+dS1OpWgsrQM3tFKuWCwNHo9KRBmRIxVRGHHPReTrnAztGxZE6Q4nq+C0/gyA/e5nNy5BX
ndhu9ylvrxLMn3gChlOgzWe0BIQtxUqI2t28zgJKE/YleoSI3XiMaRNFdXp7axGJKxl3EHvCts+K
/P0gh4e+DnKaWOtnhSM3AAMafJSbaKPrqRlWJhevI9T1dKDYa6gOF2kXJiJUCPGZqW9zxr9hYC/S
jg5WmB8U/LT8sMXBeezO8eYSNES2su4fuLIyXnCFsQkvAMVHXQewAFXLFmFZ3aAyzQjWplmCWLVF
2z2SqFm5aPkccKt62FeCjxWv1CIbstoxK0r0Ts4fSRfjGRj8H2/yGBJdlEfawEU4byCh1C/O1OIx
9HAL1jjLXe6udoVmWbaIg2MNdPu2DRR1kLwwQ4tEadI55RNHf20GRW6H+lvXrSJuKEn997VxVxxu
RBK6rXxSc9u5M4qRhOilntca0aDG+g4yeOjlb8qvwpa1HECxfo6hbE7bL8k4xJaEgtahAa6VNIQD
kRJvrHqLhZwOb12qX1Gk+Co2pdMrHeVAVGjmFDbcyo7BxECnRrkGFrMq68e9nwxkqzgC5WFYUES5
7+zO8W//U2Jqgv8YhFtDYirXBt++P4Djz2LcfoB4DJrpgW1y0zcNSiazznO9Wh30jLYmXCye8rYf
97oWcbrz3tJWTTkUeajGWbGDDD3rLXXjN9gWLg02V/EcdzjoQnPq/V8hIGLS8yyJ1DHlOuK/zpOY
R/C9iuUOt6g33pOZvksPlSi+RIoCv8G60kGFWkdBMwVpS3zYmgJF0HMeqtvYrnKID7t7ZuqYIapQ
oz2Mwbq4hPkJwSX9tk2zAZMKfQBJX8N3VKTtgs7XvMl9udfR9GCg9XGGvySXsCOvQxGO9wY3xLxu
mF9NdxCN8b2HOF799LDBnhw+QCnRX779axUEVGX3FkviF8L9V7LlI7tpCi4j0CRf1bvaMmpteLkf
rICdj15/sxBnRaURuhlG83u2L+LR892xy20zB/2eWcZJRwoRkeSgBE5XojeDmq5g4tF5CILj251a
XoFa6Aw/HhXQHeRel/3KiwacDEkviUUcx7GypxbrF6IfKy4PT982kh0MI4E4r3mOxHj2ORD0RBt8
k0WJsRbhYzZWu/vVRisrbzvGcVMuFrat3HkupG22vz0zIpJ0/u7IS65f67mhlkJ1hE+V+i7TwzHh
87VmPZ2qL2mbNnkFToMipRRbcosx2VvVuNvrdGqlUuPlArR3/MvuXOXn/DOzZY6J1L5VkFT2zx+G
6oqlnupT36y7JUMu9eRvs7+PjB1T2v9ytTgeoWdjhGa/wvl+dQb9rd50N6VLugdWYF38WXBjQ6Ft
FntEsTbgpjSB7c/dyYx8DsBUM0nfxnz7EaUmvF1bM2hvV/xV6H03jBAphdi3Frvy54z5cNhsJGU9
pre+C4OpDGlBJHMnqh24MyP/tG4lpz5NkJ8XN9jwbDHd33JA2AphIV+oT5NhyoNcazI0MAYvybja
ztO+rfoS8cnZ6vqhT334DDEcmQWEIFXKhoRh3ZxaolHzO4/osS9Hh6a2An4hl5CWNcaXE+lYPFGH
hzTMdD2ueIKZaF/B15CT/slqNtsipHOgL7CvjdyAwfDR5OcncIDiCE5+2RlWNBPdYU+wM+womvE5
RVcwJPnwZWt4wVXjBCq3GpmyfNreZ4xo9xVCsj2ntocpjLfh/UsoVyC+pC3EDrpIbIXoP6XIc/Lb
K9rhX2XwYAi7IWSCqWAkX/AzvD3UdOOoeDBcaLI9CDwPcZbX105tviTFIw+Rz+A90uZAttsjG/5q
v/PApvBZYgcb2+GKFru5uv5MUSESDIfY1Av03AdRa0LK/SuBFVmbTdsia5/PNQYGFJRQC/vZzrKz
OANRkoqf/6d/ED18fi+Y/JuGsKFVfpTMI32g1CwHMa+zYj1cwru79y5CH3nbwrr5/cs7KiIb5VW+
PFi8jF7UGz3RV+rwOkw2YndRAeREtY6wIowVqGyT/ZWDTbF5XZoyfCRDCjGkCSGzLcc7BbdP1800
n9ChGwYQmcehLci2UUTsryE2ZtsrWEGoS50dqAO5SoS2GSFB5sEkHCC8neHVJpSKTAcTmL214Lll
bCu6XdwhBOx36ckw/Wx0Rs4QAKAam+gn6pw2Ul+K9Oksg8EcFfjEoIya0TX8Beq3u5mAVjc0xasr
j+LUnMuyYR3XG3jlos//PqG2obSP8VQ9miJ31LJIR3YsZ4M4aTslqZEJY3WrDrIs5OPnYuPS2uCd
lv/WuZM9bR4VVmVOAxNRxbr1q8PRolbHl4fJ+0i43CNX735no6VtFWAviJY9q5ay1MCQXd6pJRQw
5d40CQvTN+Kwp1TmYaf46K8vzoaCY9UOUYyuXvLzxqYBQ479Yr6SCuxNn7hur3k7xWHwq6diaVqW
Dc+V9BArdKMDJQdoxpC/XmW1NpgUui7nNByVWiMOBjgMMYPdnilqxWjV2T2mKb+MqedYBEd3hELm
8Uh3dfi19NDrp5gYVbSo51Fg+IFqN7xsGwyaSpTDQ/I9ni4yFmiWec32I1aQ5NnXAy5TEZcCwUin
yjpT/r0BcJkeHSIMsLo/xudmmIRNqRFWSKoD2/rQiGRFPEGI3T+Xi+fX1P9Fyc92Ck9FmRK6Iujf
f6VaWIb1rGhZf4VKd8q85xqhcIbM/Zu5WOxoHbsXqGe8lmhZhjrVtiL5DHW6rTcqL+u/RLuvur9n
1hoBB/+Y7RBBIzBuEQ59+It241Q5rLqx7kYZApeQIqn07sFKNgVZ/YS62TYnpbuo/GVo8466fKnW
1MtMTvs1+N8YKGfERJg27hnhkIzrNzbJ+CjeYPIm7jfWNV7mqwdH2bd2YlYuv3shYjiVCG3rGp8I
PQuFLoo2eSTF5tWQVM+udRBySAA3xYF6CKR0Kk84XOb8LekaCkaCWxNCPrlW+iUeHrxNe305Bhm1
Hcg6bGO/ILiPxUzWC/SyrWKfimEOJpr7/Oc8mEZ0UVOVXM963guTgOkhmdEGLXizmgU33cvajtN4
IPZ/eukAbWSUJvi9YKubrtrc3iHnOBqUBzpZkiWlj8YKRYqTqRt1idW6XVU+Ir70/ib5A7GD5Ohk
hM57qrbLmj8SzpfdIq6Bjjfo32gNqsKbzMGZgfhkbu5fHyihug7YslSmFg7/eZymM687SDW2SIdU
yXvt04giMHFpfrDcIdbGXHOCaxFxP15IneOHEXrSwJpehC7lObH1X9zmW1rGG+SAq+HokZJ8fMPH
JfyGCwBzMVzL38cPlIJP4p9ptyA5lp25H8r/P34N6Lnt7wRsBl9boyEFC7Ls52tBkow37r3Q8Q3c
clJIjZqzj74n00uOmXrg5bLXrfHrEu90Y9smRiC4CPTIpUXerqv6qHqc6sHRdTIIkDTEr26CIiV9
E87chnE0GsU8sNgqK+z32wVKK15HzHdQ3qPumLCxVPFnz+8PB2HNV/wrM5MKekuyr41jksDJgLyG
6iPu/VQipCRVXNcFAvl8t4PRiAbBkBEh8RMpyaFTr6hSZtJWlZRigxkXlNVvae1VF+RrYBNMRs4Z
8YQPriRPTJNqxTQwBJjsNW6jwPD5JbRpbh1At/hHPkSziRa6ZwtjpVPijAoCvaCCbJeLR8fwd4LN
/8sjndjEdKdF0irLkq+Z27T0Aivg+mNSK3Ma+F1Gr0VRtMSoirKMgrJdSaf0SEKbsu9iVIJt82bv
vvynsIkTEKlhKr1Z0c5FOKgTWngkxbn7L2rrC7WGIwZGww9jiCDiLl8ZEqYIOyeuBTIMlTAMWZ0K
V7WzFqQsThk7JGnb1PhHLIcmo/fOmMTPyoNmDIgQU8c4LyaBUuIJjPuhLVJGmA7WETBw4TN/GHRc
zGoKxdYx0aBnBcvhycUeZECrJjG++miJNhqdPMOVBLDJ0yrW54S6SDOiO4EIoTrPwa7HHzRolDh1
XYw/QCxeG0C5/FEXdDLgQGV61w8DGGbzS21GlJAVuIf/xjtPo2z/4ruT2Itvxj6dloBbBODtU/va
CT/FDdnhRYWJrmKVFrfdFUtTl3LrhX3t2Ws4Xg+fli1PyDZXlI3Cu1by6EwgEC0Q5KvOERU0lNht
eLaqQWuNq3QqlSI7YAAt1cfG5tDVgPkHuSrfwvBENUAUz/gFux/mzx+2TzW8YuwLVRHT0OFd0hMW
ini95UXLwFUdkBWVzlNgi/ogCVQ8u3e0j9SLWSJXlz62dBvalLZAFHrW9WCcKZuaEhtTl6UelCCf
Nya79zw5Y9icjXfj0YRknH7p0+YHj2L7YefT5a+zb+kpy0PevtAXJbclXgkrJRT4gb20C9PFpJqK
e5nCmlBLyREgjWCtdnmcTj8u3w8mNMTABmvW4ROdIBUna/QSIDI3wYPZXvJRYt9n5hOaleT5lSXe
A7JJT8gXuKyJtJ0Nz3A08KSaoEE1w5Jt7pn3nstyROGL54OUKOsHVj/+gIfaCBVCVNqhIyk2E3H5
V59gbmhFrrI00kEx6YbDAXOHn6QCcLUbShbkb5yphtOO47HuWqV0t8D/pgIPooxEa9JucBq7YTeI
yBYu+f6EoMpa4ocKcxKSRR3VwLe7mbqVd8y/BpjUtncqHfiyyxV9MdeyMdOs/oGihAgRNwQgV4dB
7wspNyI5g7qFSD5TUFuSuH9TfRdFmllX2EMdhV0+m1gDqTvZp4DfcAsoH45jh9A1PDfPIsZeGUf6
7ZjBE90HCQKBgVS9jUqPcARpwbJR64rGhDrvFTjrR6ERGuOS9U1vWrFX8cC/C3LyUfZVS4TQmTox
87IeS1YBWKtzDWW7cT8U9It8/MiOjM6wlOHogEBL9897nYbRWuOLVdoYK/mthdqnF3wXhpRYqJuZ
BTuYCbdiaPm5EGuvT8gqnGWTLlg6IEIDil4XL+6SK4EHqV+39VBz/+ulTrZVP2vGFSmiPHX/xYOy
sWuRUQEYoVTOqQCV8lmPc8rdEaVafrDTmS5xnH0wuQKsicx6tJU8yUksiXYXnng25gPjd5qPqsd1
LWb7bFCUmIEWWKL5fH8X+dbc94LqN6Qwq+x1mxeMbeHvuSK07a+gwkuJjxm4qRx+4gF62FTFfNut
AXSWVA7XlYUqFW6Byt0tWMCGxKErVAGKV5gv89DkYWDOYmtWL4sUDD084LNN81mRUN8OTBf40LUM
C7KPT6p/vBDNKtPNrllfZxT8UelYD/dZClZ/Mk8M16TtxrONxAFmb2ovO3SE9qnrxyek8UnUqz/e
kgZ9l0ppV9YuPshafAd7gT9UpbZr8evj0WEwBWSNRZo+E+lb+5G5URQtTbHS6YHU5/Gd4jeqXIiC
rNcIFnWtqKYpOMEteVOMkGF7DnVUlHYmttBkarGhSIR7ivT1FpeC20/BXObzigLr+muBuzpasM6o
JLi7AQLPVQgre6VhApjAkeRb1Tl1bQk4BdZuwL0u3J3YS6ahXTLj6Gyq+VZCAFlGhLry+GOWnJj1
nJVVjkNXW20eNnP7j5OZElDRYU3C6tW8aX5X3RxX3K3DXB5dtC4uWSsK6WhYfYMpx5MBPajkh9p+
2X3C5EChSP4ACWDM2Y4Rgf61SLTAWvBdG4OqfkTvwYV7Bk9U7hjEOtlSQEX28z5cWzpMGocQv/DT
wh37z7bEt6QoeB3cnKxr2/0m9HACOdylcjZ96BJ4b0uhIQmaEDf/uEMt+xTCdIFiGZyQ7T/omww9
J33Tc3chGUrofW508xA97WHVqtibB1mQbKqk3Kzp5KtjHQXn/WJT1jdR7LakxeIYC3DqNEHlEX9y
dXRZJoLBuDdDzhy8Mdhvj1cdFCTdNCww55azsuTD+CFESZOTRCpiVdu6vnUsYGmHNf5eX11GovbF
PIrKal1ZVeAyr9te6pbk657KmNhbozUy6c0ZcoLqKEx353SiVQqJVeaHRpmITCw+1WilPNRT5KQo
3W8fcAXYAgd0JvPxyyrnPebM9supfcxCNnq9tkYBa2u5fZKqY0w8O01oJoCWPo1nZz1mnRh/jgF4
gqg8b46mdrbl2Xcj/zoY2OGvaLkSx12KbffCzhFoTIy3QqCIC0g1NbV9NMvSrO37PM+UOH/J+brj
PX/IGD2Cams6FgknKJdGMqGWOh94qApi4B9PqOJP38bb7JJIPgL4waWYbMfE1Q5/keqb3lDwlJaQ
3tKK0BTLIrzrxEOAWeHblyTj6MLgH8yXGA0ylAe1tacUeJK1f0ouGU5sUz6ZyhZ48nZTk/A9VhOT
GxDVdabtGVkQSvbFutNmB69N7HzzulycH+YHQqXNHLQW8NEjhlaXP+HGrMiwAp/H883oeSespbCL
kTDsoAqFKn45PFwsgdaOJ+c1EO4lSN3WMvGjyhtYJ71Po0YhOHbKveAhR6FB2ZjXfIhbezTnDln1
nBR5I01/r/eN5K7rSwhin2RRE+ZB7KXsqKsTMRLBzrjOvN4DUSL+bBpxQ7BNLOYXg0Ch0JB49kKn
OdfCq7KznNRclqMVJZDbCb2PXqc2fc5gWgNPZdlz5/rubej0tr+anqGBtNaVX5wzbuopVlXA6uD4
whQPK9VZuOxOlksQ4AME/j+DmMM7oS4ls9xz8hZatOu753c/2AL+2Qi1hKoUjcmgntyUnKhmuYSg
lR3G7YD4eli4lN2/7VCKNkPTKb9w6jPRWDBXl45WK+EvQtak1acRFft5KH05W6XfPLuYtJ52LMo8
wUD6yRWViHZNau0pzw4wQ/ZE2+OE3Vw3zs2qs5QyBTU6H7PVZkFqiyzEuIYrvrtUg5NhFPffwrsG
Hy6iMJPMjOEim/FD3MolJEv90LGYRCY+HCtveUF1W4I4DjBLjc0/HMfU0PDya5OCiHdOxbdL9WXS
DKZyZDVu8Y+NzeuXnE/4rnExOjCG7jhQkajcjwAfXM+C9J3rfFpPne2cIGwKYtqT84YV9DbQQjfz
v4QuRUcdTg3jFLc1hCheZN59gTT2WyX0/y+kQUrtWnaNaokeB968b5F6cu9u76BE9N9H0AEw7mg0
iM47nw8AwLy2xYq0Ziv9U8p+AlnAd+j/QYXDumIkDOQ7TvBtzScDDB4nq4AV23iV+MSmzYYnDhHE
aurs1EY74PFvFDb5t6F0TXNb5wxzB2gM84i0hIBe6YQObV8Ge7EP0dzyJJy/SDnV2k3eyhqq0MZh
qDT2xJkzh1aawLQ5lpOfNyisxhRvQMRH7r/u1nCjci64aaKJTHHsi7fBja6n6d6Nc+m1jOLV5HAp
tqRcNWl9yqbaMyJCir7HXfVjBQneKHj4smgP1Qs86/qqgEKHF1wGtVTympfWgKIE2m5FGctc0Wow
B/2ddDChdgJzWIt8gHPurctsKK0cc+IWpuOAy1OpFr0sg1Mc4sE/BQOgMXeTNg3JkWTJy7nipaCP
lO1pqQ4R4rZ7fYTRcnFEoH9y3cV8J5p7DK2u+XFozOb9XTq0aVNBgU4/J1prQeaTAiHu6YArPOsv
y14w2bOItb6Q8Xq/XGQpYebHK80jFC/rHpdtbAQlcQShX+cTKdHmvO4s1ugCMF8HLIuJnbB7A+/w
+Tlq//uAQE7aErOhB5V7EViDc7pYwDZkHr3hPsrKRHjdGzSxSq0IISw0JUaHexjttx8nPNBlQ409
Z89pSvJMwezlw88tY8aUQJYiaDhcr7iflZKqB5yy8cDqPeNsb3TdtCLBvZUqKD56WtJ7+Udk3cKn
9VnuXkVy1iIgYn/DQhCwVTuO17O/faAwtfk58+jTGqvG/Izd55fL6shkCUy5N7Z7A0DV88Y1rkoI
FQ6W2ZiT3khtt2I/Y6kqKvw67lgEodjhWbrNwcoh5c01+NAStpPttws5WfqNTPOLbVOCxh6GUzNe
q03CmjHTttEvMQ//CJlfSeRO0fk+QnF8GRZIQYkTtN9nbLLh+F34nott/sTVpOEL27bVEIVPP+sP
R4mRV/Z5Z3utRDrL75A6hZfW6J+MfO+DeXcZ7vLuLImySpqRSuPqDLaamDNVMw5LoSVXYFCCG3Ys
0wATDrcYMNlAVGyvkO2yo5LF2P2pFov/kDar8q4ValgnHROBPu1MiRtfnUK5vlA246kldkosntrd
KUrNBET4QRzFWksXK2RB2UlRki6/y3fA6oNz61M5oBmhNY59koGd9eMtW41Pr6qmn0Z0K7KZpHsw
jcmkLN8Nc4Vx5/xGgTht0fWxuMxFPSxgNa08/Rq60G5IyTTP4M+XDZBrYLg/pTcXzHSPKHa2yWZI
OrG2mYaOS+7oCQxH6j9Fk6LTriwyJQaOCgoLXduEDh88fEMyo2aA5J9/PkpiAtGKh8zydPYE+u08
gfvFgdJGVZV2r1ENRfeW5E1GlHpKzJOLdKGKAQ1NqxGmVt6xvQad6fISRukjB/371h2UC6tHgXE5
cZdFHW+PKGJDS3qhLZDymq4XWSYvJcM0qyKYLFc2zatLNOpyzqeUigXsNKVntkhqYxDZTWqLmpdu
N02LxJ1CDBCd/V3doY+pI6EKDHnxzdW0qRJ709R9FANBQ4IniwquTdjTIzSsDEvJp4xCprAvZRLk
O8uizLH0ppOxcWfrGbmSgtBSHNBDFrd3zwIdfXTyhlzxJ4m4vMYZA/tw7/6KFZVcf3LXl8d+rLfe
QYQqUvwYlMvgEQuqktZBnw+oMxH0HH3LdbSW3VdzxIRvKd9c5cy7ou20LA5bNFM7PcpVOuzyd4o7
NLoWO83vMME0dNzwTxgvuq1vQd4SvQq6v0Ga7eincb6TJ2CjyD+iU0LTzlodVjj9DrrX0d+DD26w
1QhXKGwFD5VID2LSKyB1RMEb0+MOoJGtlAEtyD2a4leJ/se06UMk+MXHF7xcNKoNNZHBC4p7ZJBi
wzVl4+aC5Jkj8v7rYYgO3drI9KU5qYt0BA8/pI+eYoVWpGgDNCMgmNRj4jm25O861PlyrXmCl/n4
A7FnNIyg/brvGOJHCYvQnP1+RRhdl3nqUuFxDitSNcKQOnL5fAXILYXQXmg3iMth+AsMDIzKUqMd
3/Bi85rUpvCB/lopdumFl6yil8zvNRo1Om9VdO9WriM+9NB/Y4xgTABa5UAQ8zWlhwoL96PRq2+b
94NAD53b4Ii0RBO8LsiQ2MFUJYoZoqJsAgBH8y3YSTA+3cILV5oSxKNXCiUu6J29VwvjNlcILWv+
7PU//9D89x2t40H5RcGYWPT7ZgYE0IGagThT7QgbI5mj78e2DRoVJas0Al+oPeuH1p5RnaOgi1Gv
nRawVMVMaQplDvHADHq02bVZ2iQh5pvSDd9ZKL19Io/ZHTh++OaX6N6baeE7sTO+Bxmv4dwP1wL/
PLbp0juHTCDkF5dqrzQOL5IymVqHItTMZ5RLZ2F7WHGsxkEtL3UfeXsoUBqozubuOPCyK9yiv86K
sCelz96+YJuvHG448PvQKpvuWbpWAVuO0Fw1WxIDN3IfR4AhcKYgTSrYsBBSvkhK4xEjW4iOkUIh
NgQkVs+hvntHukw6El87HJy9ReLCugO8/oPSqG0bKGxnZ+14NIivMxunmiEMmX8+iS7MUGncOhg1
UiDx1CIhdTUgg7T/sEAglgeGpbOr4GHxmNQB8xL5ceNNS5RkpDph4E9zciBRwLu1OJNrgdkT840j
84lQTcfBUwf/MBchk7pKUCx2574f7QH99AOtZU5hmlWwJ9QW+fyNqPmzeS8nd8FyFMcSfYMEMcnT
E3SNuCkIOLEJIoSUqH6WABJxo2JP8KZK8XgAWOsw2XEjAd7haQaJRRidDE+c7kOQg6qppa4M3yxc
ucnWmCU/JIULE3ynExfd/SO3flP6toCSOIOF/pzndQoTLBYlUj9Ipt29sb+r4gCtlXmFB38qg3up
BiRFY/DqkzJmTMEqeks0OyM2uVjheV8ltYGGz87vGqkh0YzrKn/5xJ+BGS+FdI8MtMMCTrre9SZP
HZPgGyorxkp9v37G7HXVh6u9ueo9lJVhnS80/5kZPtF+kfd6zMdR0asBS09u32ll/h8bFVSFvXMh
Mq6VGCVP9Vh5JPf6shRH6VIru8OvfY9r9tHETGN3+694CAj2tEJLJ98c2EIZkQ/rltTCb1qv2+fU
msTf51oQ4jAyqK9kwNKz6bEsIR7QOmaeUQjHsVKeh/ptVPtGf7M/1cYHS0aryh8jCO3UZqcOybF/
uLNM6hhwFHn/7DU9IGLy0F782Vtmb/Xi0Y2WBh49JnV7++D+rMau5+3XMf5a7wTJt7mgCRWYxUyY
MwTIU+DwVBCWaPdwXMEt74LSdIGg76ci9u22UDoRlpmM//lnkaG3/AnzpCBpb/3Tx7wia8l5VkTQ
eimmGqU4e7qNrqjk5Q3jhHtoLvgg2IvsiEOuf7zgzLffalALWTpRTssop29EfJyfcAYMCqsz5mGo
WngIYDzFptFHev9ROcMPR+gj8ekMJeDkeIIQDIJNH1BkUGViqPkkZnpcPJhJoT83J4YP9PZ/bOE/
TOPBVdoH/KtgcQh4qLFKaJRnhYed1Iy40Wl2qchz2+V/rU+408/MEfY4RTbwHnLsiWhd8wL/da6n
Sb5R4jUReMLdzEhkS0AoSYBscSPV/wrOQjpHl42OkmueEmb8X1URQFBPPLekV9iZ4WjUMqjdqU/4
vpgDFBfiqlZm/MziHr6Mjsk9jo32N7ogXrLCieHgV2Ff43S1vxD7uxmkHAvzdT+NaqbmsqSdoxgi
C7yvBqNrMOHgR+D19DpldUhepnQE3kO5XKy/j2xh5+RaO+XkTHV6kRRCxi1v8KTxwLA0aR7dnK7t
XPvIQSbPW8Fnp+JIH+0Z6782053MKgzg8XEGZm+r7H4uZnYFa/VM7zalutDfFRcE3sWzpRmkx8H4
sfAQKzYvVPHYAJeWqoLEhX9pt7tqV0CDgbUBtzWdB8o50/IK1L3+MbysvwxZMcOCX7WXWJeAKxUt
IxHwrho8wY27Uek5jBnjdrDyKMeKP/hl0pTeQx2Fm/PTNaFKE9mR0QcB39DRrDsR2UEnZGsz+q1c
me5vcTg2K1sFWp6J5ACwkHDsD3A7H6gudQxBE2kEwVtD9grEm+10mWF7salgT5e5jX2173kXqcNE
Xloag1zCNjR0ht2MX4zruUVILBMstFjeHpgKaMbV0/50A9XYb8ZGqVRAqvy9WqUfSFY6BdqdHGG6
NsjiUYpIh/LKUXax0++dvYp6WZvwP1rN7SPHsmEht3zxhx4lKMilwbowi6E/2JKuY7ikXR9K2x7E
PcqfR5yhmC07fOuEwWgPtjH3rv6gYEVMnCy8Muk19OewinlGUSH4O+ix327vXJ+OqrVzBc5Nu4HS
DiPDUTujYH7xepXDWrx9ySeFG6BaDt9MDFgc663HN5BOD3yc3LAHMubawZtTy5nwdaeMt54FRjzB
LphA2rfIx4vRkYGYImgRFDJbG995dSj+tdUVfskZF74dg/YGWPj9QXDocJ7FYXnpwM5k7mRZUwje
8c3sUOqLX1GMsX0lm7Ma4WeihWjRYoPNIunanzWb8GOFnyBUJJkE2YDfrqLmAq17srcIRaKiTcsf
7WTkLDnBvKStGT+yWbnvQOreKqxfOYOCpmyt6Ct6CT53ffePtCTrCqjyCzbt211GAlgS0wCIDycc
Dzz/fQi26ahgiPqnw+pQaOIlteNFo2xfBfjLwECjq6/tV+R1+9+O3/8nYyR3Y1TF7KAcYt/2s4SM
DsidQySqUPMIn+E9TbvG0UHnhTldpQGFdNnWnyBfXDlCnOJ95ZC3MHQGErvFfuovCV7L4COdLtX1
JoIMHBhhYzi+NZRwkqVo0mttB8osqXaAaZLEsk5MjMEAAh+txBghs794Je3hNiTEfD9FvHli4KAS
/jZ9JVD4wnwL3VQRRSSCKor95vsq5WkH5c3HU76U7X6+pqvuzYvbiu4oMX8sJDGLOoreNNNQ2EBd
I3OGHAhSgsVRDIwl0z7jlKelRX1G1no0b0mgjPrgXDYJnE2VoiChSEDkFuHlEewZzx626jLPj+xE
ZG2E1b428YBooclQ8YjmeJ/3kX31EIBqKjEl1HEIUOLmGqtA35IPwgINPXX0y3naKhGtkIadTAWN
jwZCQxMDWrp+M4U9bB0u+TSLslE9xNaT2ThdyEt13hmS4MOPSdayaCbFhpZRupHGWydwn8fuRF0O
CofeBioTN+J1hFYfioeaJ9Cil1RlC8DoRCO8H+G7HXQO/GSs0Dz219L0i/ETusY9+F+2ZUqghXhr
nHxSkN1BtXSJrQ197EWEuuRDnSebInSZupar8O1H8+nfkesVJ19aaJ4254TeE40n55w0xc4XMRf6
t81mt+JgC+5ULEVYGKjtVNwAEtofZVDW4dnLcWuMFYs96Z3wa4mpeFdvwOA/Ma7/6n1g6tyiracR
n2jOfzr6r/UlqEUYuBhJmkTi65LQp3k1+s/QWOPYJ/xD9DxAtIVkNb/WDU0kHes7Qggh/AIsHk9g
W9kfjXii+jiQnERxIWsW9nsY37MncE4tLjxa7Nt6+Ij4RlN88/ov3Q81q3phszW2cTg2hLzBiDNg
GLcBPryK3yavueRZr5ioVYQbDEYjuQThbO/wvXg5QbOgyojNIYeABu6y+MIuoOfMX1693O6cnDh7
ChlG6mEmiIqBpfCKAz97xQPMxhCPmSKnJZ8Ei+CP/Moj7NsSMVQQxQIp0dKRMteYRDJvH4b0cwWP
gkVUYm4zNJm754Vm4q5eumAMwZkv+ZL4oFRTP6TpegdQpyTszLgiLpZpjdXO5+Y9VgwaP0QAE1r/
KbkfixsjSRNVHk58e/qZnshWjS74Wd2EAIOxJBzZYRoTcz8csLzi4lwjevVKssQp+tLo10zDgBmo
3jo7400C+1+bss8+4h9KpHhxdyeJEkGfPnoMwoHN89mf7PB7NnZw+FgKG6dusx+oR5+7yr9KLJZ1
MUKzNDuMbgMew0QU0przOKTVElf4cOKcT1LYYQ0EWy/MG8snyxmCdx74ICyp0TybG9ZSN7ZTh6kR
tWwo5b89uO6wB+0qTgH0w5gXrT85Xe5BU21P8ywGqH53gyWMCwactJMT1WVDMpP7wzRBzVfhNzDZ
mRL6vYBAdJSjNYbXzCnIqrugqvdOFN8y8XJOgV3O4tZXHbVgHe8Q/9e48yEGGk45FaI5wK4Kyrf4
pL7JxwqdciX3td+HjJiPHrkKglsdwApKLbRT6HeRGqXHBkl7BnMcZSdtc5UUiMmvv9BCcJw36ATR
hp0qbAaFvpVtTdBQpmBqtG0hnuK5Htte+7NVBwvWnTSkiav+36PRvc/U+KqUEZiFDazLDlrUiIs9
hDXPgnMTI/NevTTS11UdS71StlCYctHyf4NPxreU/TYKmeLJwuOlBU4xB/j5iz/G8qYZOHCeyaRh
HD7pQUEJp2cEX9H28Q215NSZKDKzHyTGR+xIX3fJ2Z2sjWBX7HCNLy7WkKd5jnvqEFCDxfvki/VN
Gje2rPUqoVIk0c0xN9cFeXdTV3Hql86UDOkaKZn2riHi5v25wEA7YqCx8tWeLwum4a3oZ5xPERIq
xKlTIKv4cYYoKMfIUxKw0FyoYhuZ5rZd1xMGGiJ9HCqcThh22L5gtmHJk8S6IcLniA42ef/ucdzd
HQlYbXwmP6WBX8FlorrKhRyWJmwOihjLx83c7weu3wW+0cvUHXb7serth4FQix+lDcOmAE788PM2
5Lj7m0J4BgP5jxEYq8IZYkVOJ5S8Cz2HMwo6gkPkeemarp1TJrZUXxbeFB84lc+5+C1hn6r/BoGI
T3rTRRemkKmEbJv/zH0Apr7NWi5iibp3I34/I3MKSju4QxFSACaKxeu8VrXWHnrCqm5e+LFrerbz
GOk0hIiGIYYvbgHcO/qMk6d+BLvGuwj2XXr3nTcnNTtAzzpU9vRscr5HvC4c2ydHb21I/2rVyyOQ
Fd76jAZKdPCBdT91XpnDOVfyF0U9JyEw6fWF/jnxp0SMiFsNMDO+GIpcb/r+x3fPJCNaqvfthWph
UpOo1yNNcdkbyR7chELXFWgQ53AeHr2R0YTcm7ZlugzWkYenPBWHxLZpwv0PAYnmRweAwcFBhBkf
9pTI0V3LlTWvGZO8/YAb8MEQEBJQj87ZT1SvpjYa3DaBHdXlIdb2jDJiLoyv7HoEKTMC60ubPRbv
7ogtyKxcwWhif58VkwPQIFl1ZxOtPor1dVa0uopUbaahFpYkIWFcohDv1tu9nNVXcCrPJLnj7QLg
pdrJ/fxT7NJ7plfITNN3je18K0OLfLPCMKH/0s7Lj6kN7IUTZtRrSXfD0n+Ul36+se0LMBdHamx9
RDWGtshO9fy7AmLJlwB/kZc+74uR1tnv+Mkyw7zo61qWQw+77Yz/o3q2Nei2A1dKm+AqUtXIeiQH
0G/0sb6w9oMt7OBTZa2jjjk/9rVilM90++2+ExSfMhqvTig2Qf8cTKAxMWkHPevdq0FgU0FaePFG
NyNKbq1L0LKUx1/rjdk9bHNJ3/sLHNjRWHTTZvJfn9+2azYaicFaTA3UfesAzAarI5QbfzzvtzxG
hYzFTCi4n/U7W6VJNJ6rbhXUbklEGlqa7mZdigXSxta9rwRpU5/jcWAw9zjacrGSFaIIYEs4FOYD
BEd7LzUdXvgbAz81Eh5/muAiJn2CfacykQByvTqast6A3t6VpPM9ovDJd3yqAt8QQPJya/TCtHv8
z/4tLWV6NlWvUUMNECawXKOGxiVzaamnRifpI7qGgKNQbCi5ajTZjOHs/tvslqhQoHZGysKH/FB2
gHORj1iN6NyfkNaKOWtOp7MFVcI0MMAxf2RaNnl2iP0meIWEylwvDf8iR6/xlOA8nvWpdUHS4mRf
npv1TYOKWIuWkAg4z97aIsCsqudISF45EJR7mNHvzneCJdhjUwDET4GtgepJJ2K0HL8MU5sOD8/m
SoMaK6E9jt/Zlj0MidC0ZLD8gRjgqGRSFQo1QNj2cOzLUXzxPE3wRqxEYQcWT9YtiP4i958CqEB2
ir0i/W+mh6renaDfpYV90OcE4YdnNelCMoIyiKnFf3IiUAMGK/GgMHWbMZnlzqc8UdTVqdLAq5xp
Pndi6TP6XFIcV98ICynVHwnh4n7tRdP0m+WMZSwYDdGgKXM9NB7msDn9JEFXjd/kfMPNNcMOYo/+
VURHQrhqGzDNl6UWC8WoR1NgOkZ/YE8SLiiIygO7CdbiHlCN0uVomurxbltEk07Eiev1pQoCUaUz
N/oLbwT5rvBFxYajlzClHBAoj5lHcsstHRASWbXQDpSuP+o3XmMeAbdUsHyLenh3p0ZPXbOE0gcD
NRRrwLc7nrdB15MozOGbdi2PUJFiP1lm7HNdv5lqWYSqyqva7tJDElWFzyvSxkoZGHD4Vh/YtgrA
uYOpepirFR5huJ3aFHCptGj/Z9+PLEf64+WVy7AF5ZfPpzNMdqhZYjFszItAS2fDmrdo3AJ4Xmtb
pT4xtzayLI8HttLAYZNY27P3k+BX8jXmwTA1na4vCwudK1VnBejfr6b67GyHEPE3xp7XZxHjmFww
/E4qbSgrjAg/kZuCrCUsD6HIQFn2Z9TOEDivIWOdxv5ouboY9YtpadcZlg5SdljE5nB7o5Lq0Bqn
qj7RwyhABc4MyIb3OC2KicnoCYeFRjn8xW5mP9ThFrM0nexMqX2ObHhcfUVEwA79nC0fhpLDZNez
fD7YHiAoSeirpp54pJqRz+A9ltfmQwKaWTaU8raYfY8TYSrzstihNN/dTeaKZzOzmBjSpICwGmcH
D1uIdYnfceafiWqn+d/pOowrEWCJ9MTWdYi7M0dJ3uIBlhTKyVU+hHerjxHVocdogBdBa5syVuMd
rsNHauJwHT59uDDHddOeG+uw7r1xXT75v21V9zHpohig6K/8at4P9aSMzzFi8NvtD3c5kTXh6p6M
hnwcq8Jbtq2PZeNOfYPllAu03eJhZGBISl/oSLp/j74QSZWLRz2UNrbAOrCdaF6NnjnSxN2e/j78
tONlJzM1A5A8hZ2K4hZnx/FW1XicoZtHDuqD5DeWIWK7+ZdrYxxfqTmCrB+19pEOJEnQr7ql5QXt
vicVmHoDvv8Ffmv3IXPmlYx7or4kliOY5I4BI0N7/JKYa9l7ZiY0aBrqUZtnOIFB5Cmyyx8rZbR0
kEV9XmSD+3MiZBfbx1vICkpJOHu6af2BfgS+LjRclHi1KSlU7DZ6LbkWKZjbGN6Kj7ZyfUpysSUv
qyRg0Us+A99B0ksGJHQjueINCmjUgXypxIvi3iX+3wQ993/GsCJCFGx2nDcRWfY/EcHKOnqanMJn
hAO/XQ1wvnglxLk5h0yn46bDvMjnajp2ZoS1obvGwN+TZpV2rNVEgYDeF1A25mmt1bVVM3Ekv5N+
nxoZ+JyjpamHMDS5Rrn7zMJA3WvJm4WXsr7pWP+aGT/qJWmjkuJOBbLzwSJOlOlvr8lxIjx3lIds
CuxdTI9GRpjVc7B8wbGy0+Pgyn/uZoXw6nfvBX8fyWHjqaU6u4W05530p9jMVZXabvdeYki+jb5t
24tK6H23YBR5GVy5pE4Ah5UmVMiiHrKpi04cn1aj6YMs4yRGxJReAbMHs/sMhc/pJ+QICE8FCRIh
cGpgOBAHabX5mQT6tv2gnNqCCTDV3uo3xw7qo6msyzIlO4yux4f0sAbpQDGp7hLeSY+dbwLbPXWm
5bJyWWV8o9EKAI8G+Owmb6nAEz54E4sZcWA2D7Oo2V3wKKm1z9h/Jyosu2zcFMngDJPrXcz1u9ai
P0vC+9BSZvBNNHvHOqdsFFrCHq3ph3RPgB/Qhf60lCgNjzIH2nIc/Lal6mQonLv1ieUaqh7IGPjh
X9L21PsrC+pbt6kDorkdT2cksVVB2zeBrKLPVog+mTmBl6TLXQVX5O9yx0+yZLAuFTRgDCC0nkqp
oDgIyxaBPMTaFqr/xNeb7Fhngf8pjxPD2y1iygCX5E5P0s4K6XggNsjfHNL21Od4REP86rrf+JwV
wr3Bm7TbzI9WayibJJcV/XjIMlNS0LN7bnHdKCtdQPFL824nU5B7ygt+xbt/xRK0oTg/3lyrcgC0
DVFbB5VAdkNXOVgDtHl5o1ltjBQsHsB922T62TUurWV0FAj87QQL1Jlkr4wy7PG1VpzVmCNY9jpT
j8DOwZ+J+rKDeDJBxV4UTm43Rv8fiseFdYYZRfsCyYHhp6jcTHU8LH+7hI9XdtfEUn6qTbQeL1l3
iJ9geXLC1ELz5BWKAPettgXAKiZeir4xE7onbHAVSF8mwbjS3dzO4heBgJA0roNbuBQn+6XihShv
ANiSrGh/0Ud4trDEQZKvrQLXB/GVd9ETGQez+lyZRFgxcz9gK4eK2IFiwKEqxjrQdtj7c5/YNK/a
cMZSH2pE1NUQMCAl20WLq26Xyn4hEUzpeI1afMk7ZMD5iud4wGoJ0AVCrndQ57mVqsFGu3PD/fyY
RQ0TbvlxmOQGQLMSwABBSvCP2JN7RfZx7XU57pdJPa9I1JkEhuoeWRX7DbtmmCl3Z9zmCfPh0RBh
VsLx9E75/oaRr68CdcJgwUSoM0qkAyJSJ6mCKASMltVZfGm+JYg+TLJd3AZUpA5wtfVcT9uFZrN1
gqLjH81YaR5MIIpYTJ+R6egzb354XCrA2f6tHP4wFKxuFHhsZj+wCr/+XS52Et1bvdyBqxQ5ASPq
zzO7JFjDsyrY8EDgWWx2rokDxcpHNhlxnAxxxrATN0wXKuk+S7x8usiCPhnffLln5/WWxcQ0F84t
PIfvWK243XWJ2SbLxOCHTorA9Ch5Y9g90kiO2L00AqHCPmvEWTXJ3KKdgZqXnFjhm1cC3VbZ8ykh
+nZ7r1b9zE9yUrzTu4v9uYZGyfv3vUt8VXtokT4JawLEeCsri5OMUrgBxQBGjI0zOtCcwday8ZjQ
+AHBoUCjw+a6TWJns387D48ynbETkAY1lixYJo2M9Qzp71SHN8VeiHR+cdgzAZJ9uDcy56NgTL3u
FVXDs9XFswqfSsVJM6AW1c4sHiHU1hFFoxa2HkB3OsXym7RNEiqB0utXD2bm7gQvKIFU0KXbm1qo
KIAaGSP+mkds32M/LuCIauJFdP+OCxLbhUKrrfMpPYwKYVJeEWRN1lkT4nVzk8y6UOjUCB+4msMd
Ih1MmCApNIq6U2r80XOeyzLOCa2rM2QBzMm0bONN289tocN5fG/sNEJOnz0cBj8giv82CEyDQEb/
WZmscvu/rdMv6d3nKJq0Uh/Pyz2WaGgZ5Okuve15nlKjT1Ndsn4/c66lPU5ngtps4Nrl0fpQZiH1
chOcipC/qUOcO+RW8i65e5q0IKAWsZ0F/YTue8TbOzSQX70VKCsLLyX4h8olqi2vAN1kJonx8GV7
HZg8PPTCN4n2vTwPb30Jt58fusi9AvgiCuYy9/BiE8v28VXcU5cLEXkIIADiLdP+5rtyF1fCjMqz
Lt1zeBWtQmqo2YwLFAuR9XxggkntBC9s1XTbsa/1bQ2saJENyFUAC2Tan6Brbo67c041+Gz/vG7P
hZeZ2EdOm5La6BY19eH+M2Knwh9ygxJjQMIOAljHdLBVDUv76/00TfFbyjE/7wTwmCygdzSUfZff
dG27go7TPS12aQ7SWoK6NoYeHl2agtgeEYHpqzSCXoCzpzNfMUH+AKaLfe2z614Ij9TZe4LmrWVN
0HkgwW+mSM+PFt6BsYKRL2mfgLz5cz13gcxcTcZs5Njaqel+D302XO+zv0F19iiU4dxoKfyHEPvj
azv+nHd8JI5UQ105XLCyMiNbK7NMbHO8MQl96ijP6CKrd3CZ9ey0iSmVK5BD8ZtbFVhIuRuxah6j
xiNHt3FkZ+Frv2iTZoIGRNvQILbL+xbFsbjfdupPfQf/BOLbvGm8aG3Owff3swEHzAjl+NKV2ss6
60BbQDkWnWkxrlNLv6knMgFbCnHKRcokKGqSNaym2V5BFwA7vEDKDibUFeZH3MSTh8iKhj+gBmaV
eqIpi4VZgakGK8MnJ9tynoAR2fPZ9pu5v64DG8NwlxAgXmrup22v7jCcXLyt7mpbb8YkEUzUIHSy
yiGKacuxCwOm/SatxwQCWiif2d3heD68XtakjgFxNe/05c2JaJqfqJ/wm3BvhREoRbFZauORwpf1
V++wD1Y/plHlgMW4NH5MdSyilv44g/2MA+Ym/hyaGPz+X17tWGcDaeKYfdKTq1udzGHBarnRTl7D
vFmIFnqRr1aTXuHC+Nn5+UzDA1s/rLWWuiZLdISL+kfCyhMLnrSmhKTEtKgDFI0tzKxwYupl8NXf
/4mwt5UMaWf02rRSlwxun0QWgrxdC5iHH8Pu2UuPZ//PPVdRwBLA5aJZrUveDJaRl+yxUC1FwDtV
B4hqz7zgtNaKgdlPG/DNdnpTsBVKDTehUzuUoYiAWtQaE/lKT6zi+IjPfhU4Hh4RgUZCxEWmo4H5
Z6MbMyPz+YXZxobCzGRbgjStW9Hba0Zvt0v7SxsUvHzgilMKu0UYlaSdyjq6GSl4b6f5PszG0l8C
0UJwSsoH622Wz9TDmBxgu4AGEkIqbzgbtL+ZIihYoF5RKnMGzrt9BZfBH/vduanODE/v6UzT4S4J
ChElI0bPp0+TX+nVR2BD4b7p8xfGJBEcsKt/YbugDxFpZ3JOJO++uEECmoh+dDNYnKuZQClv1bOB
BAnX+1dmJ/epn/xeSaavJpUGSNAOQaT6V4DyneXJkKzAk8wRLTh88yvHIkp6XRbZr/N9GCLCSSvD
ddzqLNjIhJ2M5KSx7uWMxoZ9wlJUVUXTH6L9MllfnvhSYwygsZKjFN8cB7rSZwIL+n3WkRjNQu4O
0zA1X1snZKkOp2F3J8FPDzoynvxWUWbfzkvyDrkK1E2g4Qm9gCDVW5hQb6O2/JXt0Jwk4sYWA6fE
lkwaKrSoGcoqQAHNkHovzLowszlwBdh6tg7St22EFU0GabMucUjuvBTma7H4JYbek3XnDeC5Sln0
RJQD3r2mGvLkYZFAQx5azVcWpay6yxgulmW3oIMUk1yem2KlR9kBChcGjl0WF5ef1p8VJnMXXSL2
dysEecOK9SCepRpaQtzcIOU9j3K5LahIaMS0pvT0IG4QSYRvgJ4JpnSZrIrdgaNyuvoBgXWzGDRB
uJkvfc03kMCffNvvC5U6ASZSBhdWCFiIILWLuVObUeiiMpjepy7Dmwx16Gsg3+0uGUGmE/2tPevl
KEifi8Tm9nXCLw7qyAGpvCEJwsDXQZ4SO6cc+h4rWisZzt7Gtg/I6RXjZXUqYXKPj3Q36PSw7y1m
XZssjb2+BH7LY5+uDP9pkDUbD2cy9qeAWzn6CJuU50UvOiUDI8QBXWMJ9V43wrpl2t9b88h2xFtM
Jtpku6NweJSu0zOUiRUS8LfO15n1JqB6ROuw1R2iDCZaZsVXnRMs9Kz7VxD8jenJU+p0Y4wbLzLS
3Qe1Nc9J000wgItWjmjOoNojqevtyFg6BVx9jtEqsdx72KHdGDjCogyB7jJ+hJg4TNBwjzgcSRvY
Rj8fqeBeRYc1qcls8u9KFxLJTU7smgVIEALR6R7X6UqIPNeQ6mvQwgkaqUZeBFjXG3Z7iJeoky7N
WxYtBl6401NftILrWX5L3k4fkP4YpLky6jiYbJIRKVMG0C1sGpFTtBD3gDfDJpH/B+KiYkxEbhjK
o/PiXOpUiOSzWlBuRCYy1PyLrq+g+w6J/AZfBIJ4Jdutg9Te7AY2jpJPG5YrZHMhYG84lqE5zBve
ZhcDPbQQ91WZ36atOEyuEm1tVwuqfSb3nBHwtyXK3jVTknwoOQ8SGMVvQRqnGOO9YcfAt9xkMfBy
NaIPncmkDXg905iRKQfAkgZ360YwMWjrY+whZLJSi4L+Na9MKTNu1lKhMR9Q98TRyFBryHzCLW57
AkPCj/fQzf7oMplJmPsrGvRLI0gzroMOMuVK0c7MIFNEvjZS5KX8OcrnAqbZ/M7ge71D8CEAf4Vz
RI7RH8pSJkpc3iZ2p2U1ivIw309jnNxSl7uawpfdB6Kdzkmcly2syjOeDRAjhs0LyF8a2MAYq8Dl
0qhOjA92NvOmQXk9TRE0rA5vpYf1BOf7PPKxJngl9JellZOgnLd6IzZD33dnH7TLT/grBegAeTbF
ZviEy/CIAwQ25Y9Iqqbpi3/w8t7XfKiEs5Hx0xXYOqqfcSSPeZ9i5jqgDYIaXdJTyCc+5HLswzit
DVl0Ol5OcGg1agv4RRv7SCb23oE2gbVSQ/RItDUXK2jB/AnmSyRxACTycA5Mz+SiA7TBDL8G7Few
xYZ0xOZWkIMzeP4Cn2PuvLk6qbMnDhFUybz4kJioXuJeGM6V114LZIrsOd++M9Pmhr2hWJE4wSkB
2Sms9KLA9r3ETIiwtB0wF5a7z2GroHMMNwtrRHK3H8M5c3EbywSqwPnA43EcA875M/f97CBjcyzy
qmS4HdODN2W+CB8/hEs2z+oOj1Q4CrAy+eD4Y6ksmBMgX6sMfwMx3RP7km/IUFvJOKT0yo1acLQf
o9eSbgrNF2Fk11tazPUzcgSODGV4+FSGi8iGA9m+Cp3EYmJV7Uha7oLr6srbwE8yyfQMIr203nZm
/i2Xn/5fSPnbuBDf6cykJnXyTzFwHJG1jDwR7CocYT9xcqXIOENV8iH5bTJ2L87l51qfYSZJvQhC
frW3uKc4QOtaaVBZke0eIKSBRsDSzNfkzQbg4kCUnGmOihopMiNAeUwwOFgAKhrgQtvXWZC0H4ou
GCLTv3QP9axyNnfnNIOp7tcykwwuIC6m3HlFPcxfqqYnbvD2nLtkddFyEt5IM9KATtEhxg4sin70
o8BCxttIF72c6FGJnCvj4edc6+5IgYYY4wWay0mpggOei1gbVdvGtZVV9Rrt7CNpWum/TjLBzfYw
WJQ9NcD4pQfaSKult/z1k68lXLd1YJRfVM1GUnyio8K8OkZKzwMwbCW+S/m2n4VnnvinDZ5hYppD
4YVOJ/S7YifqhiZaMKN722Ns8hTcef8ex4kTzug5TL3evHAi46pdPma+7MWqRUPHMlqqIBOegFtn
Lz1CUi/8UdvInhqJoT6pOMLQzlQ76uuxagRVUhXihJOm6rTy0bUkpb07xITkZDV1BJarqtnywlal
KG/CuHU8AwW/yRJo50kaHwsHvIjwowaIcbwpNoG3btDgczFVOKvFUf+Aw6KcDibQ/hjhKkdizYlJ
l7l8Vu4aQpiewpyOhK75l4gyOaYUUIoULALuy2XcNiO0YxfbbNBA3IiWb4E2c7qYFAwzR6gCwnh+
63t02VfDs9ERoO7Wu7D24Qtu2hMOOnbwwRxp+vUSp0xEtw6GHQZMCFehKBm6gqrzUG7oyAN+Mzg0
n//ktbssHls6jzUYcBqGgOMAJXUvkYojWPXPhz0046B5HB+NtlFqMXzoTXmVsYG6AQoVCAmB7Rrz
b4lRqPlJ3RgBHSHqfPRRH/Umi5oJuf4pFL2Ltk01vr4hxfe33u4e7WsKYmRVwT80QTHwmVmn3Otr
SXVcJvtpzMksAq8g2/YnR02jWaZVf/gkU9gN4evQQzNEaVcHvmd0XImlpNppwrLkXsJhePbj/ZSJ
l7LfLIgOTzzw/nkSqxERHRj50GNl9OLYeUpZiyTpcYQFAfnZjSaw7m1aysE0wlcuLFGPBGlEyLCu
IX0FXG6c3K9qCYkkp2X0tH0v0s2rwD0SNIKfsTx8uU62MN3fASVYcLsbUYpWAxlA8aGknEvXGH8U
NDQMNq8RbrYZEY8AkY8mMTuvhLmKoQdgIdsDUw122cigG4XNho3TaNeFf34KJaxjtpXTprAbEY3+
arUtvLxRc3MZzjnqCHi/OBxo0hxaERkpyCAPjzDiKOsEpFZRD/mOYbA2OWS0nGuAfsEqW/40wJcV
1ol9vN1eBRdV63j9CXUcZiq/jiQByTpHGfBq0NhaYWKcUgTVv6RJ+lpwm6TxuiGn2Ro12pWq9jFq
ho4xiBhRkB6u8iAiXLI3k1YLzPYPtOouy+TsPCno4YTDkS3pNk/Lrvmhh9+q7650y4jF6nZuvjMK
y31OCSOhQZEPCOBaX6xNIXoXp0Tr4uCSm0tSrqk5Rd83O6pgIg507zL3xn5CNZNBHFjDLDO+m5fG
KgEFPJV2rbV7xCa0MsEORfcuZ6fJo4AJ09bJbSiZmtWtnmKqahjuy+HC2J/ZAE5unYqoI774/xCj
Uj2KyJKu9AAfh5MRwkt0BfolOXvHVIjVXHy5cBFYWMHgCHLqB536t8U8+xoe/g3GcaAIZR7/esF/
XNK874GfZKEbaRwDxy/7IgCCnImnOEVzjOQsvkmtbRML+Md7acDUbOfW6NY3q8QNTfhsFzkLeLrh
/SMoqCWbwkZnOd6riWocm7u5xMG6qWbkzT6f0I8/MqhHYmHoQR4lu6UqTJuBPBNl2LRB8ql9O3Rc
MmqRYfynN3scMI84hSlFNc1D+tpcjyzzxh34e3WKg8m2CHf6kkwkGDl90SPZyjXK5Fr55g8ZuHf7
oeLIlNOU9Z3mkrZXU/9yZAH4oYTjO7F8I/YUY2ydYGErMbqBvqfurRjU9RQC5/24lg8zsrnoK3gU
T260Gw7Ua2dgouKh7RS9E6AKw1Q2k0m3mCJFLcKoxLG98i5ZBC8dsyoLg2eGNPPv1uqA5wkRsZtZ
SXxa895xF5HMCM1KtwJCGVSeZR/57Luva0gSInWwUr17H410dlUZ8NdCzA4Kz6PbdPbVf5FRDRZm
ereLurQfEZBzSe/WtSlvt0AuGe/QmSXlhp635Gn1l6ATRffMOs8ZndbMTXRZFyyFfabCYgfVLcWN
tlJU3aj6ds3UY311b4ADYF/khJnC3QNfbXkAv9RBSlBAa8SThAbx3+wfMta6Tr2IrGCVw3ciwzvf
JNkMN0Kft9suwBV4nCjTMnjod3/T3zTr2oa1Db7xpItILmzVAr+3L8ltNzPbc54APV6KQtAW8GMW
HGh17FSeskLkZiAEYKdIxLE/JvnyuWfwfEddhcYqP5DNdUbpoi4tvoN6XBAVeiKoMxlGDhN2izlR
/wappTF9e/fcFbIZjppaqKxd2TOvFFsP6ROJaWOs7z5H+8NDotUhulSFt4QVf/fgHcjzETFg+5Ud
UjXgrapMxZgrnMMJobnwDZlvFJWgRJwQatMerpajD+r9AYxmlLzKP80q5ZotjJmGjGsQ7w1+qnaJ
7wcB/3JaasfBniA67CUxrmrD7r/ym1EvKWeXRLfvrHnO7tJiRSHGyP5RLRCirUaGP+K6Vnstu52C
qkwVdpo0mf1LAcyPt5iy/2DaratjIlofik6fqcVGBW2/e9uukhgec8qW8S4Yb0LVhdb3nUNhF5Yc
f5jwmcJgjqatewYBmoAfSZO8Ok043bMJW1fJXcgnfy78f8DVF8F4MRvPSB/ZbyD/emmFp+avozoY
W7pcxTVeOD7jpG1RtyYjqYDZeCSn/uGb2Xe41E78mfDw3GTirqoTL0F77RYh0EMmrfC2qsv4Ptcs
2H7EK3oMyPU8YvgeIIzfu7EzG9N563UTncojoUBiCRTp6KFT/fu2rVa181CSszSKREBVpM9IRbG3
16UaoVWRm00UAoGjdM6ZygtL8k/9EBqRuk61J0cFfb+XRCaYVfxi/5pORjIOWo9euV+2saJXZCzr
l+PM6n7E5D3BHxnhQT0vsUb8DTkwy86Ms3iECR+ZOr4g9u4okMa0b0cKGiE7WZXelJ3V40Ag99kA
D07ycbAI+1CbtCum8PGYiAYVl4sofNl/Vlq/nfQR7jyc8OgwtMjml2f6ykvXpOcb/+L4eFnBLdN8
v1GkfNBqEYLxAGKDJQO4ekfgkTLtmAy6IvxNHXz1c4flfdFQmVrQoQ0aTBc2IumEHXLAMY6rUBAx
PGwbbMrgbTb2MVZ1ArMXF7M/jt4yBpeMex3kZ7F5DBhw8agBsurdp+YbFMSs37v6FxLsMLfN+TU8
+P+TByZJ6n6e0S99rpf/rElCjw6GqUK1VeU/gey2GV2+usfoz0yBt2d5FmzIW70g30iFzyr+3yqC
lrQxVzggsKNbo/ZNihI+tpQwXQky8gXdJxUZarYBZTVhGMdxLu1LTLDNFcdIx2TLh6AnGl8B/90Z
TBJNosqmeYAt+EJyuvHsz15HBgjfOQTvAwfAbgLcpRPlnGGf3/2941P5UtuFqGKpec3puzwXRXwD
jZ076kwe4uPv7EYt7V91e4rW9GgUwXUOKz3qajEjGNdbIQ4GpFJjheqWDM2xWpqY9REr8c3HZ+7d
sYKsc910iOK45elqAFHETHwsoxrjKmI6ZjcIG5txdRZAg+qZetZ0pHXStZIs/dBs+jwCmrpQSBWI
ZCmGp/JxKoy6rfemveJGXj7lKK1vfO2wUxmJpDiprvzRmG0VyiM+JaS77tFldemG8IREZMVDa19n
8e4tG9v0dJBohsk+e1/SqkBPdlKjRUBDJxduxGLEBHdZliBf2rUSJzyMbyMaeXjOeguDJ3KyRyvv
GKELRMCVTSWBz+efUhnYdrYsBqmVylojULrq20mCsv2/VYUtEjFVr6ngYOstYvNYLCUzUS7HE/o6
HplOmpW8leeHroaulVyiaZoaPuWWvEk65UMDdrTSnBb/50NKb4mllTdhutk84hbui6hDTU9Pl+wy
L9sDk0jjsWbsAGloKVPt08AMA17ncLuYgCiXR3tpOdl+JpxeDW4r5SeFP6A1uUxtXD46KF+xccPq
9Pop83rb6V9cYr9AVsoUnx/wOA5wV9SWrYRv6gbZryJQTjApktMQse/FT4UsN1HFt1lKb03WQXaW
H6312elrCckqLgCZ8jo/8+ZhJLhuoZWDiDypSpp3Uc+MdmoUrCbvWD/i2Tn+qQYWa5Glwak3S6n3
zHL+xVP6ecj3wTlmi35ojkgxvkhoRUpEunLOghFWUKYJL4bS1tkcMaSDZFkwOpDgs/zxf2KjhWDm
hDg9305Z9jWodgmZ+dNAWmfOq/qgZtsbPAd6HDyYR2MWIefHo/s1ieZJ1sSaZyrKod6WpkCrB7ka
S1rzY1YCJOi1gdJQYE3IPqtYppJXtjo0F90XjBY/EcELPjS0WLhQnBeJMlrQnYFNDJPx6weWPuqh
MbdfZcQlADVot5Xu3GwpghKDQSyOj1H4h9xNpJp3QbylHrb9U0nDei8wdXWg2LcV2cl1enS1v036
F8gTYamQ4QghLAWQR6Jrpkn3nzYltf9Tv6yOXGvHMP5Odae0H0QRjOLrLlMdG7pU/+e8AVhkUR7H
hnxaGb4g0NogxZlDvMFXMwuJVRSiQ2Uoe8+vEAePz8EERWCKyrFl31pqT157YRv13uUymzFPMM3d
egfpXOxT0MYUOFzB8KsFIdMD9tKvCPfjpIHibkLOREHZeYtPu11clMyj5jULGxvjM8C007N/qHbs
Ux6E2fLUZ0sppxxk5ADE0Rpwqe5yH8DQljwrnlnQ4NZfzlF6mm8BnpVvCuVtOs6unQh+RXW7nAs1
PIv8WQ8BDUtmq+UOsLy7nuV4MQj4mABgxeC/lND4dm+kgA7le6stA1fTQSSdAESsMtwTrkoIGGWf
DUUI9iyUPUuBn8E7GMFwICh3a65vMHcnee7X04ukEBSc6NEIAQZmhs/JhMH4fmldq1cduGLuOngM
2JcHjDlk0UjlBLA8ytlFih/F2pdnu587lX7PHgflMhuNAHr6Y6rmB/oQoBj5ZnkFo2wf5ADCXG7p
+VaA42YspaJuihMhXledb/HXhLeVqVZcI5+ZfjCQGEGSGGn2NvTy2czoc306FfacIZAef8Abl7o9
wDnGvhbRD2spFqbjxDJ4bhLrTsB3dg+UD9FbJuIdRe40F6GOdde5jSvCLMb2FuZsUa1G5YTMV6tL
Bzqd8PTIYf4uuX9g+F+sJJ7gZcLGcs0p5GVJ4KdduoAokFXV3+l03TwBpBURWDu/sIslVuWe04Na
ntgCnEsIDsQpQYoW+vhJBp/rFqVcj0n03sLTyvifRxAewKybs9uy57oRABr+wU4XO+d4LBwQugfJ
b9AxV7GW0T6nML/L6uVXzr3me2bZUTQnO9oC4i0OZDiguZ3vzJApADWSYW+AKQjWDkGvzTnndju4
atkDxrxT67bxEzN31H5+txYT2WI5CmjIwm+LV8Ry7v6rv3B/63jEtYJRd+VFyuR/VZZRhLKz5e6u
79/ktBEjccyqz5ceIQJF08y2F6qYup1FPMViToar4cjAD5570spHf/MAEOGlcNWgufM8ewlpFmMN
0Kh43n47bf4k9QswPoOMP1sMQ9Z6m+0c3dILivvYC9tpND79WoeQnodDZrFCsykweGcxKCziQl/y
6ISFD6y7ptHjbS1k0gBatCnnbPgCjQ5e/Kk4aaH8UG9mUBwj8j0L792KcvgCUctCs/sUQ2gQ+Z7G
OUmiS/QNb/CryEhV0nu47NqXy35gFBVYkIz/6I0Ni+jZ2iffytB19SD/URCfJ2EB5DBL4cFG9A/p
8V2rzKgBQo7QNHZDejYvj4MohZOqkqIt7LedEnmJXoZjHQSytAyXWwl3fbminUdGozTJUzVW60Ts
R79L+3ZGWUTS9+r83+RBSIhuHRKM9AdcYPPdFhRftvPTllGjBL7MK/mjVlRjEwNF2BnAtXXE7F3f
f0vxPptaFklHI+EZQE8k7/XRDQXps5APrRrQYHQBiqKtGKt4luEM5MzjPA2KuxdUfQSNiA5Cgm8E
ePU3X9eETgBakaRfRdjy0PebkXH6jjSRgptOR0Z6Z/gxr6aBP/nehA9HPaJ5WnENwZY9jhgXbpjQ
LERQRYzDNbes/9kEkhAHvlVEnGj4S/1Wv0VNC42Rzd1clHKzWpw1DYwIR0SLOTwYe6H+3we80SCI
IFF5bfj3o3+uhN7r7/ptEOs2Q8rWgWxZDPNK5RqH4UlvOyZekMHDpjknz4rSWnm1XJPlDzqbpSmx
FY/CXYEprZop1W7FEZxL/V2MuSro6pgsYW7DvuFSpdxN4VLIA5bDibP6c63u3S2d/h9oQ/LMPOjh
A8leb030qo7l04Onea5TkF7uEg2nLNTtOiO9VSRlf8YhkD4+6JJQa16AO2WqOK1mC8NEZj+Bfg70
Jumvnzmic035+kjd/5bVxv38DZI9G1BtgamWRDjeCiGFEkHsVqIhR3J7+swtF6Zn0SM6wwVZZT7/
MGjJ4cup6DPcNKJiUf85sVr3AYRRN0yjQGGwVU9uC9hs5hqOW/Af2nTKm1GXmco5IFPg6mDeWDyZ
uYu2M50GHgY5VWF4f0wb7FEsm+MwWCEjMTpX9r1tL1eMtVNFdwDkhquH778a26A7igRA9yXT+FeH
DqJFAOks0vZHITeQFh8nhjmuThfIN8oACAzAD7NYmOOt4nb5pPTbN3x5h64EEgAR7luCGXQ1d/NB
tp1I4zZDKwY8fSNTKAWNQVoTQMfImGLzA032OhgLU+DoI2kZLGuItNDoxkqIEZUlKAav1R3A9csm
PkuvTgafBdYAWXHCM75TmosQ8OOU4JU0dVsy+/J+bKO8fl/Apuq2m/aYnXadRu++ZDxdF/fFepz7
/iQzTNIIn3OIl3pQHKjiQixlYS8b96Wyfsfe74wYoZNp3p6S5D20IbxDX6e3KteYjNG9p2Jd2aae
eBzC+1CihkdqQIHSuCpKzUocuqS7zG5F8M+YNmxx9hZpJhzMcKv/63YPty/tDlUgx/FPAErKecrG
XQIdDp1U8Hu3tHx9O4i0k5kMEog19DHACwwLE152YIrgCvM+CctzX30jtZKOcSIpMJ2Twrgvh+RK
Lq9Vez/88QImIP3k2HtC8VI4ycmETHEkIWmoa8y2ba7scJphLasOMn5pCs/yP2wlSGARSkRg1oMw
TL83TAKjWf3LmVP92gjb9agJQt1zMnfVdHLTelrDp60y6PP8J/k8c8z+cAMl/gD5Ms+8K+BrSbkg
BLyj99qy2IhC5MVBUApKZyFT9b2PeGH7Y4wnFsfDQc8Ne3ExaaAc9KzZWrMAkWpNk/JPMopNkK27
0XTDT1M2vQ1ErUFZV7RT0F521ejnmBYWKLzkY7AQuRM6GGRTeXFruPhYnurwPesmLOYnDyoeGt8o
n3fzyW5yhsIEYJAciBH7aeIgXW74AP3Vhqd+pdSTaciuIydoNr5/RrSuNafOV/LnHFfleYhO0WUg
3kWdWeHG+JvdGzW8TEXrFkKcdE6Xpjrc4TDxJEXjtX27i1RVMK0cF4b7Js/Yp1YnRXNZsCyqVjD8
iuQCRMnaW9VXsldomSnDiW4vHxpzXvkH4SONnYk2Zk3IIUtxDZ481LjB5SaPBnXJeX4gbJdR0qeU
cOEuYsRleqU72JzNn6hqePQgdmgme1gmUAJ9RAF1SbCpBiKHlvTGNr/w66fy2Ka9JUtXziaKY8DG
lixBUG3CmvV5HLIuBPxmiiRYWFwi5P8jCoAksdtbgZYIUq5AcvNqgWF1ka+naSz5UxxXRWB7R2+7
GpzxTI8MGfai/QMVJ4B/yUUzI1EnExDg7IR160XlBzxPYLCmJMxxr+sy2G5DhFPpI7YG2fWdPiAX
2ZhqCDSo3zlJ584Mb9fjVO2tSAhYpvLKewIXAj0govYkrp15tD7bmsCBhj2cy59TPd56pH6r7rrH
e55M+qqvnPUA/z90ajDEXLiyes33u/L6iKzq8H+SmRtXFZPp5a4AQFVtKQws/sCuL3hrHVPUJ6ch
aq0FuBa/Hm2CMPSKk8O3sEVn5Rhu9YXUxuQxLxU3gK9mYviS4wYAya1XA1EnJGbs7VItu4Cb06xf
r6iC9TtYo9Q8ORU0iafnGtMc/T8RHeK9FO7Nn4vjLM7Ba2TzmY9qmikMJgphsG8oixfJXgldMl3k
qtyq94N3kxTJ3c1Askzw6wk7vGNgsw+zrXlQmecTByrzomD6e4Nggk2q19jwEgSEVVFq1mT27AD9
rNMWEIvQ64z6N9dfPjvwT90ku16r/D2eDcqM69dNaekKgp7qUr++O3Y13LI8Qp+We7ru5ju+3NaZ
KkqWfHOJztLR/6ww9nhP24t/akHEg/HodLqyZ5RCm2KYQjqGO0nWLrLnRXe+r5Uty1HO4tCFbD9x
98JPxkDSRrXuD5hiQnDKAmQ81ApxzUU89B+MIXZX2DvyBi0oU1z+pIqM9rQtCRrwHJzvQaLH3NTr
eESgWB5zrIWB4skdsO/lHTuY9OYSE1/O5pgvtlhbWKmID7pgz4wZBazKGmPlpljgNG0Q9Cd1qJQ1
TvFdmQMZsQvcS4FG+VhDnlRrhmhN6b9c9t3lUg2pydDmVX72T2Tz7gvppQFruzbvUhGAV+z7Mbe6
BfwQH2itALLdNYKhIipvnc11YEos5qknEoIcwuwLPVOhsXIICwu9hhCjiA/pPMz4W2cw8FMIW/Zn
onY41+WJAEkmgWiVtWnpuwuBAClL0kMV406QjJSnCYNXOg3CN3ZwkorKDdV1/pnTa+fI5VZ1AFEb
oNVxttgY5Rc6+V5uOvmxL4egpafux2w2XOl9Kh8fuaxqU8PBSvoM2cP7OElNyncvS5mqFPSyWc/j
jFxbDRDAahseyrNGS392DxQZDvqDi6u1AgxGH2WvN3oBwAgvfb65vRQ5Z/3s4Dj5s2hxPbga23sN
8eq0Yhzoz7/yr1DyQEIQJwnRXjiSBfgJUx1IFx7twK121Kmyj5YyeH1mYAJqHv5YqYQfdvh7cbcv
ZwD6uR2Mvj/U7tbY9gC3EYS4f4XXxbFDxi+zeA8AKvBKjexA3YpTeuPYfWKhnZGolKyvxq5Wjn9h
SG4r4oJrrynz8QFezfMjzUpfU/rwNQfstdpfknvdLHdfnvSyE+ffP0J9Hnp/tJg8PSDR/VHgayU2
oomB9HJ2lnsOGvo1ist9K596vNIMjvqDuJ1xS1noTneb7u2qcDmqQlQtV/RWO4FL6rkefXFLmE1u
1LRH0uQ7q5f53z6DQXzj69c3gm44rxh/3ROt8r2ty7hdq88EdSjFVPL1tyqmI6//7pZURDAwv3tQ
7Nn7dqybwfzFktTZjTnV1i0XQ1cYCL/KkyFUHLu8s3/azWQyimjGF27EgDGepOKGdnXh/PMeg1z7
DGhDMk7HaHAYAeq3w9mb3B2fbMmcA2WqlSfLIQfiWj5ROAGjtidBVzMVzO+SJjB5kVDUoD2/StYd
Mjo6TUG3iSfKPz+yV0zmXLRnN9+mImmgYvo2phtycjp1EaWYyI3uKFLdeLg0ucwWV969zPRyodBt
qMqJdK8Vzr6qVdMdiBvmvwocwuraHY2fZQX1rTzwoZH7gm38LKMPeEoF3U/o9eK4jLFA86jLvjT5
7g3R62dIH9VIld4mOzU11PcMdMk16LL4Wsu9NKSHDFSWNX9eMjhSMo7E505xgfpqL17HqBVdTa0x
S9h8hi5uxq9X9u8wNyLSmJTPNcCR1J6TJfm4j/7ev7rsxBYBDJxCD3ygISki9l6W/4SkOGzo0n18
+KMyMGpuwPtdAajGIgZLf0pzr+zGFguMbl+yo0gBlXJO3xDloKrix3BCnjLxq+CwJojsut6D9gII
QEjS2K/Iqyh5x5VBsyfTtmNZwepq0J07C5MHzfiov+v7N85M3DjokBYYp8ZYAoOjxL1gSUb0lKK3
MWkd2ltLelbAJL+iDgV54ZQeslm9+f/UG0vCN8HhABemTV4zhftrVhbEogav1p4h+R/9SyHejpOM
QaiCCg2Gw6G9M8Hwmdsg8g4YpU/wM3wXfH2ojtGu/AUbtr6WqQ3l3uwXXY6aHur/g2b6KujPiVG0
K6b72xK2NOqBQAEjVgcDY1YPm+9XLt3okw7UgC55iI7IR42RMIyBYof/eDrtgH9np/tATZErEvUb
vpfpKt/Q56PgbvXf+SFVvYR+kXwfqzeBiIONn5thtSkYTRHuwco8j76zC8cLUigpa4qKYw8140XL
AA7wh9jCwkOf8NTHvAH3CddM4iYChtv0K1rJNc+uqTi4GKqudd4AZw20OqSqsITY3+5dzMdANS7y
WyUTS4iDCQ05WfT1iPTrocObKgdx3dBelrhn7+GrCwdd83ASEuyDOD21cx0adM3OF5+MSXxw+ziH
n/4gJ6zRRXToFIGBpcSz6RcwrYHbdayCci3rUhjTy+Zqz8mniAPqnvBf0lDaIl/yvBjyx2SB42zo
v3VZ0LMCNX8kKw8wBr4tBhO5PVnNsQyhglSoC8tqwTw1D2YFyOO4I/gU4Ew0i8ClrPbvJqrZYE5j
V+fc4gSpxgXOqdNYiLVhUklPz8EFTefY/+eZPdwc/xE6KbZxrUP2U0Ev+3UOMr2gssgKnJwwNttj
lpPQAIDxBAQvr1sBzGgP/Dc7zgOnTq+0RIs/zUn4+hy2pt3wA1YgNgYvwd12c+5FKhpZjxkMvnCl
/xd2z1JluSwrxFbml2eQ8JElYwo5/96b/J87r65u09q6yW706NVUFv6MHjug35t1uroOaM7+e5vZ
pVe604RdNccp731ajKlhXYUSTAu7TbZg2xI3L1HhMrzQp2MQcwpLa5Vjw/fuWPspJlBEcjbw5mb2
k0VelvltFsQZD/AIaYSTFVqu8HtYuziLeAGEly9QbBs6Y98aQHWf0OMPoWmcPkIDZ8zfwDACOeWP
AoJkThKLMuGwUX5k+rJrZ+78k5bqLhp+VwotXeyj1ci8kZBtPpXwq5uEa4L+KtQk12upuNggEQLN
rW/qu1BbeCAbK+zC4qAJ1MY+qL8KUkTnVh8sHf7GwV/jfevyb82lbr8URqueXuUN4Up+v/m0b+T9
TlLrd0dxLKv89Bu+uxf1zzTzuQTZobSuourfftziOGeSgAuwZ9Z+qInRXimpwp7ZS9nXzED9719h
MgCsmDKFDfWluibOscEfEVRgajpeoFBv7vpmAZRSt+M4tkIPlJkwO2r7ABLF3Qvcb1eSF/mTS6/1
gja1E/WuS7slDwSREiANBGsfQjRWRIh5vz9KMZ74svdh/F/cTiufXd5j86SrKwE8MxoCYoCyU/5T
l4h/8bcTCKwZsL/CFNc7N4ogezfqEwSyFS2MeiX3qIPmBzEqerv4qxkMRBgbm+3kmYIdj2gsTghv
J4WhgNRZ4i4y7FqoDp14mTjtotXjMeoiBsoMeA5Tz9mZTEIrqtn4aFq0avy/06LD348/WjOcynoP
PVkf1gCle0ljR+0/1sDCnmIx1DtkxnmTHcSIt2FeQYioyGFUKIaajCVjF7gerZ2X1C28XoX9vcj7
ToYycmfxbBQ0plo0DZrruWSDOK+AW3s5nr/tUMVlUSgIU+Ipb3u8ZiQWATHb7sf0TH/JgHlWxQc3
PZWQbQDgueNp5lxTTPWek/YR87ep3GQX9zg50Yj2sV0Xl+cofhnry1gd4l63j2gsmkrwyc0U754O
62/LLToAvkBg3JVa4aZ6OkCLzRo1db6JVFpDxXleAJ0aRAy0k3Hj2qW/9QOMC4zwXs3GdPVqVGxp
vzxvTUTviH09RlLH8Fml6pSPv/XIY/fMdOMQ5D0ukIFYFmsmrfu1/PqaTe16saMwylnJLlgotB4o
2dthX8p7XiF6yAv6g1vjb8p+lg78aOrKD7TYdOe/IH7sas3sl4TI4IzZ7iC/j462CnOn8/drMuEK
KvwrNpMPTMMa9u4Cl9jfnWy3mCt63kneH6L3u59MellecDZ6+q176+aa13LsBL4ST6OXpqzDDSh8
/X1hFO0XUpNDnOKX6mzfMViJzoDXILOkL3zaTEUZZtAawUS+lvEW3bb8C1ip3Q4ras7Za6XYul4T
BUMA7V5wdOjy+gjy04cHp0rDxadNinnom6qVbKyAL26NX628iIaco5NT9/n76pBCjBwh70M8wiVz
wjjLbMB/+t7Ds2Rzw378eX4Id2qgLomyJnl20xkBCRxoI4hJ4/kd8yZe7U8ywpJA+EoeMZfp6nwo
dD2T/DuVdcLBkSq4jHmRgQNP4/Ww7q+Hpu0XdgjDZsVs+1DGWAaTW4MextSc1tHe7x7lE9w+aA9x
aT9JDMvZ0ImCOmNnnH6LR/MGNZtXOStuNkuALuac/jc98UtRyjguqzcyUme4m44LwJG+OT2eB3Xd
fQ8kiQ6nEHw1eYfpvFGfDA4KTWuz8XgwvunB3aYz6UNL/TP5/qiWBSxY1yavB9PWVVOscu6gFuY3
mNaSJO0E2/F6aYYIFqPaSS9XLZdG1QAxfdpQFQtDPkHS3R9DwRbf0PyFEN5tEFLw9lzkL6NCMkfm
Og9S2Trp90Gr3ddemgH6g1mNT0VlxOGTqhNeC7iKwak8/i65mRwimsZS6clAgox0fSXaJr4GDwYo
Chy81eOTjwpcsQM8Coz6Ridq8N3v4TnsLZWfq1KuC7g+D48TxoQogtU9cyb0R3gSPK/48qRkVApK
ZJ2YdNsh6VZKJsu63bFYDS04eRveQMInzQQ0DcTNgtFJkLteC7xfj+XfSLQ83eo/f+adtPm8mM+R
j7qDnKalEEmGLYC91mDfAXDk7Vlye7bPpll20agz7mVv4c6uFL3gEqzJ0ZxY3BKG0q0tMReDU61p
5FYgEizJugkqut5hBxFO0LEGEApt5duDfwLV64vd8wYeM+MAE+75WpC2yGFbkA1jHaHxldr4NLD7
GiDvd+uOU1PlhFVpKLycwGDWvGnuqiXpoTpG/Oc8r6TYTBfRBUOjLIK5Mk9TNGYC+XdFwELxZ+zS
SpVoRq/xUqXF+g1v1aj34r6O8uSr7ssyyBmUeD97Zzbmh4/PiGDrwT+sjPOcdG0OHyrssw6geSuB
Dbu9pl1J5GyLU2NytnDCZFsq8i9UVpBLlfwV3k9YGprYmraBtV8CNB2bxSEjg1Pv6ZQIUklldEB3
hXlMh6dk1RO4plWvepcc+a0OacWSbwyi81Bxi/foIub0n0W9apIYBYSKSYmJCnKmxomReztUrnzF
oclageyudiAlMDrZA3NcHJFS5Zys6Ys6PTd5goPpzUfyoFLWdbyJiWJUvHeLt2HAzsv8P0B2kusR
SzxdpChTmMe47zxtyaWh3dbImeTL+eIWIzNE8/Z9j9jSGfo7/OrFMfXb9PiwoZ5UHkBzQszebMX7
971fHXonFlQLufpSFR1OQHI6WaHgdVAzS60vIH8O7stR8reSUxzNlHCrktot6/MS+SHiRe6LCBbW
/q1cjFnQuplFQo/MJAfeyyMotxh3M0WvmIenpl/pWeOIEkTsxpJJdFV9SHKN/NXhdIRAh2Hd0Dgs
uM1dfhDTJyfl7sxFd7+ou+r5E1vZaWAnyCPL634s4+67LuqWYY5g4j73WGmHg1OuyoQGBQ98gOVe
HQhBx/hzXtqejaX4w2b3efrfWuww+k8qOz2ogpl3Y4gugJWdqg/0ddEuvj2rdMP+7+4YccyJbMns
OiWcYtGgzi6/DbX7F/8CqOF8dYtz4dO/KsK1zcl2S4GH67EsI0eUZvo71AoZE2PwiYYk7zixdrtP
8DzVuJkaVxxGB8HvhPu3/oIpi/pmlWzxzKNtrIJyTUQQ1ZtBeKoeZeiPSqx2Zqs6MH1jxrBP8nX4
/bsVMfst+yjlPXYK7fcaPxZgSj8Yu/8xD1Lb0OrbF6lGn18pE4SQJdRzclb9LMDqHQGdJvDU3M4J
lkVWKlOT7geX5u150JyO3X8gEstpe1f9lvWcI/SEJSHgHcjqm8ahd+fyfqlBNKQHl6Gyzms2JT4E
4w5MD4+w1lVn53hFxJLJpJXrAsYx+i0+A4SYa6GHKbmGDbxjMChb8St/55clHEMfuoGIQg+D9SBj
j5eArW2wM6cD2KO8//mv2apDzR4R5dE7w+mExEYA264sJ/kTQL9SStyasKd0PUVXz6DJRdpMnrV3
r26RRcLNM89MNj9Ou0b9DiLN9kZD6oA/DKwXGbk6aII4sx01ceipoA2ZXADA6jYu621g3SD8nld+
JJ4jJNuy8C0Qsw8xMxu6PCS3jUOYSzshPbJcNuGIus0fbW+w+gxwYFw38mYXhqoWdn1qDModsGyQ
BPAMz63MD5Ksgisxm+uDVpUJTLLCHyEQy4KdZ8U9iVxNiu9vxXu1WpXU00fmMiMLN+k6rFxjzSI8
tv2Y3fS1BrN34e6BtT/zimvmei1hNp2olU6OAYVRjuCaO9zH+9njNhcyW7+ty6QiEzbZR1m63jYm
RSIS48iZPeE+fu1LCvoD8p3fBVeaJbOErYfYeZWZrMokTbbr37Et18eXXmbkDkjwZtB4ZUGZ57XT
4zBgdUClEbEPgisCEm4EEz5nexTafJTfHu0c3QIkevXlcdOnouLKUjQGJHIx4LOpQniL+dTu49oE
bbeb6NIYM38eaMWleJQqtL9ARUCCbLSUUTb3vVhxYheH9evTMbloT3zWxTtQgXdL79/AkiozY8R0
hKYW2Nueqj1vUI6xieQ60HeTfK2SDghfEluT6vP5D8zFgSkCx851N2XuuFSSdMN9JjHSFB6ZURKY
OSgz3YHXhQIRnnaD+5afSJ6Ocwu0iNH1pOo975xfOX9VLjhzbfAaca6Yq0impAyzaqn02Y9OpY+z
tZN7CUcMBah/Tz0oKl02yb8OB93CMZMYOdCzy5D97K9B0IoqIH4Jj9nuyHL/byLAU37RDKAi2Ik5
RRpSRCR1T6w5aztJQhkE/sOjZixYRoF2aKQcq8F1IUbnA/wsyajoSV23dGiztSqDcVhv5HtZZiHQ
RwNU78SEdKfkyo+Wa2RNoOU+77ArqiPuBjCFlxsY3vIPLWmz+y4CpXdI+MxCugYJEHkxlaA8X3to
PTzyNHOhobdWXV7eBRxgISbgh03deBppShnoweP6I076P3j7YJkOD0LaIB89OPwvfmM22efZqJxg
uY1ZTvscJ8SUQOg5bWRKNer+kYF/zY8e54EjYW07Z46SE2bYsJzgfHSq6FrYLnFzkzLrlTqGJ+lr
HOsAyWchFGz9Ya9UF8O2ZYWtflDbwSGYq+YH8uUt6QEKBzjM1Uppuv0tE/yioWyZPX2BMGI31xoy
0q+NVILzYbxbbdmDIyRCBfKgrTP8bezy4OnX/m9zMg6eMB0bOPXazwHgkCsxHJeqgNwwAgiO3le5
qhVQRNTzIFEbR3Z2F6XQfTcR03bH48Mcwesp/SF9OyFXJ9iQxFfeoCS80ttUpL/y39m2iehsEJNb
XBTlB8UeMYlW4b2IK2N6POtjYbtVSeHfPQIWiU+nd58y2aCRwwNAsUz9OhvH5Uw1Hmz3sVhDBPQQ
ER1H5xc10gWFRCBtgKHi/BxA9PxSJiFbA2T6A+l2U3L+KWmDAFChZHmNcSZbxqVhgO4C7j4O6Isl
OmXWP1Pv/hDoHPGfj38BRyaerOI71iyYqFQr+IRxaeMNHP+32GVBzIGVsQTrWq5M4VVw7IKIhPls
CMFjW/E+KU44XluKWWGbOE4WR5E71PcMY+w6vmry3K5duO83PVVUP3YavWmW2rjqDL2++M2qQRcx
BvqiMpbkxkMvR81Kp8aVuIpMGe2m/CfTFrMFy2KvcDhdiw3iG0KzfxF5Big9feOJIwGaU4a63Vmj
FfH+KnUoHR9wa32t9eXik4f9bbHvyHhn3aKlQhBmIZiVjWeEZ+BD47xXKB1nBYQmeM+OupQQeGD5
2tidwmhMNld6QmL0gFxvqcfhOB/CNPZpP0PWruU1kdch5GTkE9JSTdFVOaUi+usH+g3ZS9Exoh8o
mtdEOfXdU+JOfTNm2fXNVR9ElModCmo7jlEORqj4GAuXn32XAFzAse58bN00g4VnxSwwqavHptSh
LrPC2lIBEJF/b8VrpsS6JGB+3E8PiuEg9XllnQSu2GtFyJVQS/o8+duQuybHUvgvWvIH5UVS/3Cm
UpPLcWCLCLlqNE2Zi8/BhZWh4MQcJWFFyNbm+j56SLSLv8ixYZCKit2CdPgQMI4nM2hUcxrDLQMf
w28XESnKK0x5iGO8OTWY44ogIIzxpbGw+evf+yzko+HPwyJNPyaDgZ/CHE/60cK32Pzl6rND2/Jv
Rug0oDi7vdfSEaU6aU1HtSzkJhLOKAdpj1tyVc2823ZjCU96wm7zUVj2LYKHZgTQoV0IQraRb0Dy
C9BzQ15gdFn7ADWtCR52JLK0fJDmpAknbSHOCArBindYQAufyyLAmxuCxoThEt8RcAoewbMJyQH+
SdsYkk7KysjJvjN2OXOLkYAlFdWTDGddcKU+ZBWhVaA54VYeCJZ+rKolciB3QLs9uk6pdMUbBFOG
Ma+Gnm1+GSnnI/L2xPP4mS7hIVNqujnYKeJ2TlNUV/tSPM+CNyt0VQ+7LWAxLxXLAv0TbqE7Tkvc
AZejumkBmn5Dd/ww7zFAt0Rf8oc1nB3cM3QP2T7IfeTi0W8LZUt5dBWMPnEirhffzThxFdnm8RFg
HutjSKqktsXGGwYpkbKRey8/Di9qXkBMl+sXX/XodRvVwcorNytcPVCd0bWClaBVTZBzsAx7/u0P
8uxbskpie+haAEOK7NiIXrxQpmmC3A4mpTkhb51M8MNZaPMX/MfHNvx3SRvylJ4mS4CwsW/daM1o
ZStUhjchOEQzvN1Ej/LCD0IrO6Ffsh4ZOUPuBdNfzpX/rBMYhkbyFMMSTqFdqYXHjplsi/2Fgv8I
RB962MUAYI5oslGUSuUN4mQ0FGx/1kCLJnQ7FZT92IjznDTlS5Tf07SYNT8u6uyQ01GMq5I4crsl
Oa3RVdaB2kXn7hmOStLGzqr1SccifmOpVuHd46M4NZVI++fPSy7Ap6pmxl6PfT+5UdeT+wz/TtgN
ZSEftsTOKxBu5BNAbR+d/C75yNeKjkSI3R9WuBrdL1cxBJE5lpxz6xqQuEB+yr8sG68zl2QhT/AY
I5plY+vJ5K52taBP/ele3siimQU2vIokKre232R0qjXF7W1g17/HLWyzpi9ITX0Wiks1COe9z7fL
5i2zUgxl645CI8JelZfX+jWeaMWBKz90c+esctCmBD5aOAwgvP6xHJVTOBvoUFS0oa13kG5OGEQx
dF35pA2B6Lm7tgRpr6Wct75gMM0A81BVHT2yZcQ5KD7h8PhE5tMo9EEaQ876UzK2lJGQWaCnPwO9
y+FHaaf9P/5xmDQ72khgXO+v7fIUqPKZKNSGuyLY303qsPS5aH9fc/MBLkfRCvaSvRGLq5eLDunw
j/7WnuPSt1SdDTEPRchuoxzo2kBNzQEluAXtDOTDmZZScJ0V8HioXhzsxT6DDayxerSWQQaCNNxZ
bxPWRkSl5kaqs2+YNhjWRS12OHOryRVRKNkuLZ9tIIlO0E41TVD31yijy8C+CunhhyASmyK6kC0L
fMXEGElMbzmBkzMwQ45VoCtezA30qenKIJvCn75SJqDLL1alzFK6cV6XYHE+OF3YOeqhN2dLz7S8
EAfQUZwQd76ucX97XYIUciwaaTGPvlgkCybknzI74sMDukJqErTpbAgTkWvAEjEPIhYFO4CA2QvU
1puiivQG+oQjQrcUQzwIWSc2XZ1ygL7UDTEdWS7GrEmqS5d8hpKxYsFWX7/QZgXDOcxmnFqk64Uc
Qsn4xjwb+U2X6kC7tMIhlkcQCZJ7X6/XwBS9LNVOOk/svQsC0TYvjvvCSohSquc8wwOMV57ySrZl
zO5uIg4tRdnrv/Ksy+tYNu3i5zYYuT/F+MbuowFh7p9OnNLfXfpBOR6IZQQe8Mux+ZObfrhGs75V
MocCo548X25Mt8yOA82/jwjZipYBmPt6tXN3AEFWQ8CM+mamOiGqftrN/u8c7SKF7QU3xkM280i1
bJfdkpDhXWLpsNHwuzqFC+zgEUWgtCUPMGZjtBzNgLBehMjnavlFX4JFvk15FXY2soRFkxGA/L+B
wmQyO/k8rVLK6NcZ+rN+IscE5JwtJ9r1CUVZOXhpsO1HUHrpDLY8fUgl6qrMbujdJeHhh22S0vZL
NVBNRh0wXSCM0GnEry8rkSU/Dqg1wEir7eXOjuVbhyWFcJjSeeR8iAygGpZZHJqEdrOgMTWc7klb
HOyCCoopVLYze8r0Rio6X309m7V8WnNE/yfUPuKRhZ2srH6957pgpAu8wZ6CD/WMTCcCeE10d+e6
dlw3HGwsKfUxxkhIKv9YTAGiCr8NFHNd/70+qgPqxIEsJzvqngaJVipvqc56wYygPZJNxhcEgCu6
ghu5K1Y+m8HiPpo+JVuqbc2DOHGa9uoI//pA5MTWqBGcEFEeKMwlEslp3FM9fMoLSFiH43VzIDuw
bFnF5rOSvm/Pn31iRX7UlYo0qc1UY7RyFNqcB3Xe9iwTim1ADqM3Bb7qgzRzum7lDcXNbtSRWeKk
paKIF8xyjneLJx94Gc6c5pyHCeUt9Cw1pISibMApkl7P9cHyRrumFzQTSLPHftwJoQB4KuqR7a65
Kw7/AOD2Moxm5pun4SH59IGUB8UY7fCnzzUjDRTX5VcCyfmP3zByfll5vfJkzaXJEWZQ8xDZ6CHb
OM7BUg2yTBMkFGfGJLUcJkqTpihCoWeMf0kcFGMpKCzmj3zpFn84HNbjfqG/Y2p/4vb1ohMg9QOY
KNHNUrN68AXOZLgMVeQ8ZUgiUqgt7QxtQvcw9e/tcecCkZ6W7I69VpCZLbFJSQ1x76/suM3foRHV
asALdaoLIieOIIRD07UfTCjwB0NSes3RGIPqrbRIRB4ZMAaUwUOs4W52RTdtuwik3+m10yCJQv/i
o7SvGBErUZp3bQmsGzdId97tFVOqC6bue+LmN9thFBj+J2A+pRmQNydHP3qkUyKczT8UAUQVaDAr
E9R2zcPQd90+i+Jr+8ySfyfoUM4/w9WgMvXWrCoYOZS5ToWAx9+va0POB68dtAAUwzGsbWKx1GFS
v5WFp3WJvYV5hIqHy/pat1Vxp9zNmk7hFMhYxxD+4T/u4Vwhk9wrxjNmsuObCqsFUuVsXfPGISfw
XhcD0NW5iZBlGmRi8Z+XpPlL+PjX3xwAt3G4C+kO83Ku/0kgzX5Zukv1FKHrS4UqMZbiYALl1yYl
9/ByMNki/nhxvTjbjoEQw4YnpAURjRgiZvgrx5iwu5QUC5EfZ5ZsYc4Oixqmv2FPjdT03tGrRQCP
MlNf56iRvfBcZT1AI1fUQiEYDhzUdpZ3sbGuP0OWc3j/VbUXNGxd/8z6kXLWCgBcMzUZ0ZZGj/rG
n8LuyuwtyrxpfkkaOJz5UGyJ8K8mx+96xE4eTIoud/JEWt3fV3ZdeYiYNpWBRqz4Am3WxtKlh+ai
mExl/qdyzf53266xy50YCF4hYlQSigRxUqAzeeN7CBKvqaoWl+Kiwb82A01XJ/a8pUjhpS4uXbfY
lAxHiBO/smPktFemOKZKYL0+p8foSsbtwVTapWcGSSTu9odJafuUE/udGLUwd5tnyG6+hsxi4aft
gGFEEmuzYvMU9X1k8VG5v5OE5j6fTq5Z3JuI4ZfINcPbdCJMJelV20kV3Pz8qS9+UzPLrEOf7+Tl
VFS9/V92Xai9vjeacLZOWU0TYaekKcRZjPDZyzsVB0WxtwlECBfo3AkMvik0a4XITme2jlIC9WGt
3gGFEFyAkgRRb3soe/AFaJ3XCmqiZn8V20ygzMkQn+j9ZiT6iE1C57tAE+gJ6xCfxVPRBhPgmOnB
gb78COyia+W35k8920cbMohJ+Ge/Wr/tA9UqWJfnYhpQZqwVAviSliupaSJLjNpzbtrKeeB1dkQg
i/+/jSR53nYNSYeIN7oAFZ8YcXMpZP0ZlNvlCTTlRVnpGTCBqkEU97XHV4Bx/v8LAs2Db4HC7a22
R8VbG5RKnjgh7IvyJBgHk+M6ZlercZdWZXrTQKk/u+DHMd0jFk5tFcU4vLi3hxspfTOfsIFJBgwv
h+/51EjLu+0zz/2g+lqkZJi9VsyLAufmbY9HL+AQpJS6LenpzWqvMb5Vgkt6+6FgUhE4x+9LrLyT
tnkDiteaMXcXoinmLOWV6sEXolW+wekXDcSkTonjRf8oSu42+vlfZu389PKUBWgiiLvugzQV2RJM
kSmCRx2qboU2Wc4FaB9yY/k1UUybnSzFunOrm/7389dNMmPCoFpx6nDZoB+fLJQy3rOXf4y8sxZR
3BtKgXSNhRwt3ikOuOFXjUJm5PWpLQyf2WuBFWw1Vy38zpJITzNt/d9jZub/X3eh/rnlJ3SBZdjg
lIspo8zX6CsiNAdvGSepuGWL6QXj2v0lTywIJ6vw3CfHNb8B2iWx0q0W9JKtNO2lRl9Zh1hv/Wsh
xHBLf4FZEKvohWVcSleM081L/Mu/n+5/naHfT+lDylHl3YjP+FX1PM9L27f+qIXo5dIqB0kPHZPJ
eQ5LhN32HKnPzrg9yO4/ukgj38C/dYbNsWHPiNz5gm+mLhPC7ih2GgiF/lVQT/nZIXsDEuHyaN0r
GS/APn9hD6CrNqpdZl8vgavSRGP1lGAgOI3RqZNryDaJlLFvO+ScaZ3Q6QbelaMUqozVUfGXQHFi
QF58QOhJMVUcgbWPLheXVjIjYr6+brU14HRRUm51W6QVlYiulqJ4APNFae/b5iRuYBFoehvNNx6+
mEMoFUQm1ahmuCVW3WQmw4i1jHWORCSnQhFr+eOPPDP55cv9bLiraZ4vOQK5UN5ce+pgUx0Bdi9C
ronOGZzFR+JXkemceaNxfCaBiUFKx1HfJA1EVGMHTsudw/2zln4Z7fVtI4AR27BJRnjJ5fiagcez
Q8noc5/uZAu+Ez1zvVdaipGPqdo8s5jgAH0eTkpVfnwZHL7Ny25huD7j3vicVjtuSzsjN5yoA8iQ
5v93C37MfveZWInfmWVbB7MBaqUO5GaFEmYChhwcznE+n9eqc6jjgKEIV7w9qy5bOh6CDZmf+vej
6NCL8MPDIB52g4iE16vrdNML+9mCkqh46qC7cr5coSl9QLx/YeEQSnKxHoJOnrDg0mX8vcCtlIrw
WOTHrcqYciS4QwKST1/Lly6ezN+zUeYrABoXsbLY1CoUsK604KjTWqytdH7jaSULi/cGffoT1HcE
HF1nkRC6ukhuASzxO+mdUdTvl/B3s5ISGSQv8r9Q6reda+1K4z73PgpucJooQWLx3YEEPL38wldW
6Ytg77/eE9m6+T4YSC7NoG6KjR2yIGGuWWuqXbivJEYYevz535Z16GRzVOLTg4U3WtXEtAHUBWOJ
WL9+TWEDvxjsdX7gfsGMtfFXlC8yl7guYUumXfnBpXkpPaPUR6Z9TgksXDgpvLqtRcyywIFBA9Uc
cEfepmSBOsA1kYLMoX72TAiKZrn0KqKqfBXnQRDWgLh4Ch4SgKSCMnl/HnY0wonRKLwBuSzle5QL
rc4ATr2Nlj9rnwRKIUr1QbZfQcyjE9xqxLw6tuGjXhL32K3JAaoPhLj0Awr1vJOJaO3u8Rcdyvgo
+NqHC5qkbhbw19jJyS0zG3mGXfVkVID/McBziLFIU2s+IizovG04MyaZk6d31HhgNNbbWBKg8/l3
e+jsSkY+I8p0e16zaEtOV3YFZlI9B6DsUZlYvJ271n3U6osOOytUgSm9ZK0BMKapU9qw/uE5EMmp
lzdbqLTlZNfxVDz7qJd2Fteiii/dNUNFGIMkXFEvcBZgAxcrmH1ux38O+dcDxn9KJ7zlp/AvEM5q
DG91Rjy2PWrMGSA7OIwiAzYXxuK98HRDynwbcdk213LTu3l4uutPCIp6fA1PLgZqYKuLyj+3type
kLvpNRkUNsyN/E4bN5fNmEDKFmzJfl3YZYB+JS2zOmZ6vairZhoEOkPBth4zFOSHHfUfiUOqfbaU
W+T1VvOzLOhrObsl4U0xVtBtP2+N3yHZ+Dnb3b78or0OJVQXJeWdscxsZK2r8NLf/i66XV7z2eEC
B75Bk68kaE/THyq6bbTsB7lpCCX1v54X14vZVJsrJD5lJf1dU0Yv4JLoxYnkQF1pP10Q+WnA/3ru
72TBs/WhUoHKlooh0H0O9cGndmrBX1RYxvPTEXiWNF2FVfi6yLGrmLClEmDKYYiL58R5Rme94b6s
w4pK+EbmhzQJtOtet8OWZWTtko0q/kNos4q1ItpnnBXFxtaPBRfBu683+zOP2moP+Tk4ipXBkPUc
5tfaYi+SsGAlzK6kKdvt/qpPcm/9ab/PORTwbus9OmsAa7QC3l0tVRb2NRUujFjAL5+1SfpDJH1X
1Wc5S+YmHHsn+L9FgGHli2Ws4z4qxHADpOW1GDBxkHkWNMb0azHQzW1X+ZUzAbvdNrekaOOax13S
hrcUrGXN4D5qxL3SDx2vjr59631T3NP+brNBEFbnRUB5HaZtzT62V3msKdFAYY6pvOQCLcLLOUBy
Hh/bM0Rvodug4+BZAvnsRILh/WSxJUWacFLpOHpsQhr0nf735w6dMxfX3U/znmJw4vsVwcGmRZv1
Y0ovjEWTzPwjAg9y3aGb6HJiGJJoE+05RGeQ8NFwCkm/ehzHPEml/Q23uvyfpYOgZyf8TPEUOiEG
5SnO2lQ2/L4j8mM9VA6CdZrtEwOicWQLKLh81rdnQZqvRDebk9H43i3Ja41x+qJcaVUud08D04fw
8ZZHqkqNBwRVfUNy6WzOayzkD2xA+Ov1Qa/xzvGXs5yknl5pN/LVDilCq5jsMvfTOGYIuyRbdW3l
LSktVc2jR69/ZwIVTczW6l0K62eoFQsxAQvGkFxmqw4UCOer66y7WEr/K6I6xGS/vFv5CAcdbQF2
4R/SIexlu9ZhBYsrwFgJA0nxtPzSt0KhDE3k0OF9tIofaOeuSJlyifLoId9wYJWNFh0z3E1fq+Ga
1IVEGeE8WzaEvDqH820VKruMEOycOUzBcYgAZPMDAd9CecrQHy/mlQrNc8YhAmrhNF2T9pXK1ZvP
2L38dzEfDDefdwYP93IAcHCXkHLdd8givLvnGVP9+KHSIlibe1w8wCXGlRKFrDsFdbYCJ6U07+rk
WJoGHaAgc+dA6PnfaVkPKmddmXcpWvJ40ArKSfMNQ1X1874ucTYHQH9a5+uCcaLxTMTmtX0qb3jG
15OAnBBNpyOP2gIcNt80OkuXFkT8FbHr3ez3Ux923AgNSe0cstSg21/ifwezvtMUf9EUJ6BSuKCg
Evxm9+YetIPaye9m6mLfDv1aE2979giURPk8Le8ruByIAdldFgq1grKlPto89xAcKAt5VF5VPGK9
hdkNcl2F+fc53hH13OQ5wGwOKx6nexNP3hkYbSHHLEsCMOCyqlpJgLYSZjc7f9vKKV3EvGt6VDqM
dd5OS8noMGMQ04RuYk5DeWhFA/JijQ21oIOogHIOR2qepSKiPVUN9DTHsZ8bNFwS2quVpdiskiFO
kWdQHNUvjtxpIOCf5PjDoGRiSmGaYVI9w63S8m9ki5JXp6/EKbQCGYFdFPWIl9B2SB3K0vR0yHdT
WL3WsBHiYAb7AblewrMNh0+l1pCtMbL9Hx5zzdzZiW6x1sE1boTLqDLTSF1RZjPFa32zqp0jiuQo
m+qpPQxDIC21Z9bUL7psjLc6q0beC8Zm9/5ZcuyoTyHdO/ayryXBk5ww4XFa7E1jAOLVMjoESUVZ
+Xj4BKmU16zDBwcdIsWsd6u7Xn518TdOMyaRsHYMnRWQbjonnpvVPWcIhNXGH+BY5LXUdHyKMsdX
L5blxv085CCuPx/4FF9Gc5nCnVYGcLbzH88OTc+3GTUr3GlDPvW2VECwcr2TGSfZ6pz88Imiqz6S
YgsgCr6fEn7o35A1hrNA25OTo8MkgyAg8vF1UTZutYAOKV5nGS1TBdCsolRl/q/9XKIRO0a+IcA2
KVd6XFTkN9cSp2PjqFQl3ULyYNPiCbnAgwFzRGrrDvaKZqQKPXyID1nLR0ItJFvX3MiYoFkzwlm4
0t5Uwx6aG4lG6/21q3G1d73/UqzkdpPbP+8n7XeOZc0DfBZSIsQgaVtKbZz/bedSif/SO7kRv/M6
8rPGvUJdqLgFhbvU228TaRbjFYXk8aPaiUUXvH1g8U3sRmGXuyE0tLo27pglquQ5ViC1SaR0nmzY
qB84+09wYNCt5AlcN8CSSf9twORLoJ2TAnsihLxIaoYawygs+5zQlDT/WkwBsUMMe21vviJaecwc
y4CNchJ+fyeez+Fc4O/uzWMZxb6uBOomyo4WOJAMmkXL0NnjweR1ZI31BlCm/8pgDnSNq2G66Z1k
lbeXv6SgSdlMUiRd3grqY5iktYvblXWIkkGOFpF6unzx5AGrISDASTZNGwMnJKDtoFh4hGZeK5t7
nKLj/fLMwOQdHvP1nl/tA8XiS56zCZcW9pY0a76e8xLZM7LCHOy4TDuddDTw3PXmp8l5e7xzOyXJ
4wQEcUxFJLY09b+2XyvxXgYGP2MPFJ+cZG4cml71/D74CiVBN7Tx/pATTEzcKVDwIy1jKS/E0zf+
995OjK58aMuJiPzsmo9RNBIpFqGlocNMwQDxrIs8hmyBZvOlv0OdXpA4cXCRRIsl1X1ZjNcmA66C
ubMR8eNnDHs8cpc4gJ/Z4yX9kj35BpbqsnUZOR/aQHwEcXcX1yNzt17WvZWi4G92rF40ek7nMGPr
pGYffFs1IeGLCj+IF2uhUJqulNzsDlhSOMZzMreEPxivEZX94dfaL1Ehs5RocktvfSJoNGX8VSG7
HscLq5oTze5TD3pjEVFRIjGz5tzFvihUojbizVxPWovIPej0DMlyK9hptS7dUOzYXaZQdQXZ2txS
7EvofxQ/650f2nNfC3XMttVFXKIxEZvIuqoGvnAI6yFy0342kInSP27u8xXwsbclKkdMXQAxvh9C
Zv+05UlyzjQAQZgEFDDKFXzHpKTVgD65UQVSRO2HN6izVbOMmqkufCfVUa8vQ0qudsD0fBin9zVB
zgr6qj2951Kli6N/u4wukGx0tdhdbKAlTvd3PW0VkACizscHlWuj51MS4/TydLzuWTDxRCx2/Yfj
LMCUMNQjnOcrltsh7xHttI8FUT5dqAzgwXTl5LOV0kYPVt6J92soZtX8q7BmCi5hpnVxCZWk1WZF
NjFcz4ASmwsbnluTrAQC+WzrRZnuD354X0ClhT5TjJGAdtShykwfjCx7uyZoPrdaJwVtxVmxOSed
Xh9unHu9DgGTshvNR/z9e6RxN+kWnhp7wlEmhpkmLwzpQa+yZ/FwTMqZsfGMxcAuPzq/FYK8Oc73
9ML8tNYQn2z4SPyc6YoTpQUqJUf2vvV3Ivf+NgfHK8D8yx+LSiPRojJ2WkRmypnM9S3QvnomQGjm
zIDhkVYCyQCUdfDIgP/nZizToCIW7GPFDSWM/bUVlgDeKnLVcF4xrJyY9gX2gmx8vlSYpOqcpbDD
Zy/AA07RR6uQ9EIOaUgb8A6Bw88ObGPnZpUuMhDUEwwyblp3BQjy51D0VWHAsxBqQnr2vHoJoQI9
2sTc3XMtFdCrblc+oxkfq+T+aqYNvjIgenQsHzKQG4tC/MoOKdGabePK6vVrEiiksJGjTDPClFj/
XIAcVxlQ1NuEWV/FoUu4+wQSCGgIZ4/l3688RIQhlMRHqZwvDZVnrf4woJoqoaT7TlMI0rFvIw1+
FnWyJlgjYh6a290fTpO7RT7sHgu1sDmjKPjzNCmeAXW1raPlGnMhwcBaYlDhTu/sb0CM583axHBq
vGdkdw8Rmr1UxMGigNPZ6B6/kOPvNH6TZ+l61Bp3LTMoF5qapBlLXf9WcLNYwyNHM/D+/vNIhezL
tYn0aGJNOidooGLCrinN3XfB/8W4YZz8bNexwzjWCXSi5d5mcfGqwHZP1mnz78ZFJuvm1Gox5ixo
Qp6HRljMISRmwMLBojB5hru0qNTHSS4S4e7I8hQqx35tHPnD3vGqTih1/o1w8f05nyGIffgndudO
OQzA6sbw5x/nQKUkAbbybdHVjrrg5T8oiKpqPib0/DDbEI33dbK0zmCbjsTPivW17MWYJBs1SaLC
9Jwq1V8CZrzx37nKolnrqnvQwPKfbwQoCUhCxRJkquMckQbRIXG09cN0CTNSC/lQ95QYGNCqztbw
GDOLOrA9rOinI3lcvjnpmSS04LdUrcszvQge0ZaH5iXCpMIXcq91bQ8Zs9B+U7FI3jyMy8M1vg4q
BZfGh+ZJS6BndLPxzc/hA1/q83lBitTO5u1xEFDyLTQ240h1NqoskIs93QKJnLBJGx9WdCqyaq3z
wl69thYc6iS0KDcQziVMywWhC39cP3OQ7gA2hSim5LKx4nyD2Nk/4Avt/EURJ97ac0GT7683fSo9
uzzzt/nzL2GaMoLApBgAhxSkKhSML1cCjEDPsGAv6e9DJVMG1CavK/v5wXHcg8wYrWg2LOtHyanY
bOG3j08THUWub8prVX4OgYLFK3CceaY1YY5Y0PsVpqAcVfa9x3s9E3dyCIIJGgpvGEQRWDMTxwzW
gLa7GsDrlLT84nX7ARkLWy6g8sdniZkrjtsjF14kV0bshCdDQqLaUpl8A7HutAtvBNA2tS8A71xq
e8Miw0iU5k57I6aE1ftM9hZMmNfgiQHEirezIQyGZAXBckbCJAINf15PfujdeQdfm0sjJwANDH+z
o/+6oLVjxzE3KveGuMOeGmuPFLM8EbuQMjdaFntF/RwIDyBd74MXV5iCIL0/7cNnYnjgCgJQeQee
Zi3l/tFM3fqqtzRqsrpF038wkCj3vUcUvVDCwQfD8g1JYe9geeW8UUAvjYH/mCT6VwGz658Dn7vy
B2wOuW+GP0hteFlpTad/l8d44duy3I097vVJvLuEKtF4aK1S4NaVycRhvGz1Gn5k10n+70841RTu
Qt7j7bf83T6BCf6NdKSHFDpsw3C6SnV9VqwunWinzCM5nczmoDSx5O7sCyTmfBoNqJD90js9ejpS
TI90zYuXdfIoqzyyPa8yOQOVRAs48KOfraOXbKGMENlfmEi1PEwWCpodkCQ7NXIvQpa/ESzOSTjT
a15KL6Nh59An1gL3ia0Lgb9ld4scW1wTR0W4iY74Drt+b1Kwl+vN30AcoAnV2R6SvzhqxNwU4Kz/
vyfRotqY9OfUpI0hzte5dCEUV7OE0ZgC8gjfzmKXaxvE1lL8tCI6VVlHPNhoKUobsP+R4emZBUTn
cxbxPQS0biyZvplvz2r/1Nj+vU11k4XTMumHNud3WoxtsVqLP0zuA3wQxtAmORIjMbqqDWeFn74Y
e+P97ALbNX61OnGadpljcCFqhlYbG2js7Nt+ZWXZd8WhgsqpfvJh9EqJ1kVTt0uA8LbMJfHmwb4K
xY3d0X32KBgLaePkZTGgu4YF/wAOzddOj7jd7qJG4tjDnJkmcL5WgnsFc6o9b1juCzLsu8iQP/vF
mbE+j2nkhmiO1KpHPrlfb6pBmgDqK3pZN4OWEKBpCS9rHzYCMZTxS4YD4hlydoUlL+WpOlTsdmi0
LJhTz4zf360GWbIIa50Dt9d3k1fgp6jzFCsU8ZEXIWMqvIrA5HZ9XW/d66fga0Ee4yHAuD1qgVY0
50WUaia9IfbOnuyj/LajNhudCEwPLSzjThV0Q/yKXcTvtJ7jK/Bshh5gfZ6GPe7GZSkTk3uAxouM
AXNZN72GOXcqKTY6UgY8ixzec9z45nfIOdVOFlu5gizBHmWHTPL7hEUxjQUz7PXcm0nCNNX46ifV
+AujUuDHn4xKtwyPKRWnxM7J9DZSS12zCdDLBpVkN7Q248iRjhL6jwYooC6U9BV6p/ccVfgw5KaY
ga5NOjLbT+5R9vBWbEkxkaIglI0v27TzXKklBsX1JqnaGo5qnE/B591zcDv/S9wt7dTQxaLSNysO
IUHX5BLTnAUVJUJzkMLR2vj8W1P+MBUppIgGWWyr4v3BpHIy3XBKvHLqytYimwCwtwMHiWEp+FTe
aDgXAWdijRhIGaC4/zszw6lMgAhJXNuCDAOzKwmRi+VbXI+A4wlVZQycpT6vupWVcsJJe8ZWC5B7
a6Ymkld5Ym2BZ28vU475/hiea2O/6/P9aXfUl2ZphRa1oXP4ys0lWmDWCk95kmpSAXjfXk5ApnLf
HnImcbxMhSq+K6aPQPkUT2j36fS+vKc/XVQo9imUoZjaupV42vf+snA4CPbqaTgc40tnhmdjLVCi
Emdfzj485JX0slMJ/QTSP9ihtw1UYN0lCasdma8NTX4JOJcnCYRqsoj27sd91fzpIe0gcMDrLuwh
00LdRhRxJbW2dIY/jJ39c3tFyiRxxaQQTwKsrvxxrY7RGL/twM9OeXeh9Vt1RDG/T9OiNzhz5OlX
rkCTCyaigjjHJ/Ew2UWwxRYUkv3fj0CxdURBBJWRiVkUap4g3B/PBj37SCEumJ7MlhWZ5peeuPu1
jcdtNOLfG8foCaQI+F5c+h8qv7vyMlsZ67Xiazns3WoCfLJYpc4Ne0ErJ9netKsT8qOSJStaHpBX
UET0xHPrZqEOeVlTOGoQNgEqfdjm0iXsoG9+7SmBDuJ7tPLQIVRmlITssbivn+B1oUvraB2ydCvg
84LhG5Cv7FWJkXVKsBarwmbP0eFacQVHdPso1oDYmofOpYbJEBv2i7eS1y/Kq/rM4j2qY0sLpk3R
e1kintmPMANWJi/KWWT8yiZCM/E5e2jSAdA+HlP4CpMSNL1pmnTXOLt+Pwsx2fy/OXXkI57HrVLY
DeljFeT2uvlAyeXj2S1i8o2VHmgj4td3o0GfbaT0qJifgrP1LzmOMzelOnZ9Y160V7jvw1cHY29F
BIAOAEjNGS+4SKj/xHAPie4AzY2Y1n26sBgMYgo8Ftw1dyAA2dtVWPnPVXZ0eKOZFB+1yCHCLdcO
mT6aa1vTsOQSeSboxmPie0dGSmSSBZ5pnjgGYouqVEQ+ykaSUtH/hImyQFSlbGDKlddyfaK+/0qk
KoYyF0O/uD1VddGMQF+98dSw5oromUDDuoU+VnUvL+Wjgx9hcdAGR7E1NKvhNOd2zwZPEFvzskOd
DkCpY4lV0wiuWJFuehshOJ9lnqeLe07pywnM0wzlctQ9Qbfj4frBAj8TZadxdMDdY/wMVadqwMeS
AQ9nEOxopLSWRnBmqWacQ5/Yo7yOyL5ubg/Adh6UyEbx6JpopEZ3Viea5OY1pCKDOrY1NghlLRt/
TKBWbUDyu2Soa6FBdjf6NNowlAq8HokfKpiXtZZ7A7xXpckIshCmujZCa3xHOCaVlIi2+xMqHuIf
1qSO+LixL02AH9bxjysssXhe4FxsiU2sMGJPF9K3MKjTDeLM98Z+81A6lbObz2mmTm/hvfn3ryII
jw2Cqfjz/hpBIgE/5dGL1MmEOenOZtbelYGnQ3+Ix8PJCAZmxHOrQ/bm3mECnXHj0hhC5tFvKKL7
y7wQdiCk6fd554v+LvdTNEGRD+Cm0111qCweoBCLqajqiR6rt31dyRk8B/I93Mpmxysr+lCof5UN
l8YQQiJy9z8OfPJ+AEel5XX4EW2B+3hFEiwRynZ4G2sPD5irREEDLHumwvT8U/N7grbtyhm1nGm3
nS/n8+a1jbJsR5F0Dn8Bvipol/ZPMLcV5wThGy2KUwQmbDPIeZRqBF8kkjtRSb80ipQf3cDj5QQM
Yg0LSY4kdi8s0WIN/BxJKxOmKfZVWx6SAy57P5R0XY9QuUhy356I7hyN5VA/ImMuV9vW6jSxHyT9
Om9V3QlH++voRXehIOvnP/n9/m84FKCtBJejav9YM1HUjynlYjztAmsCPS4wCkLgC7Q3vR9wbUnr
hf+zFjrZbEJLZVUkhzBb/oyRHANiIkSdXoZBjybm3rL6ocLrZf4/94yF+8MH34BPaDVP8aA3w5mD
uPkveHidcxRRvJ+Jiw5abBnfwPuqSpKhUUu88OSuk0n/elsxP08uuhPxUN7bdRSSK9rB98FNYPOQ
LHuB/Ch+DyH4tS+ppDA13nEgwAIWB9Di9bw8MKfyf3Ziq6jpip6JfX3bSXsGRPZ9ZY9im8HpMwqQ
SHglyu+tanrWAl+snIjt19haKhHg//CosOgOyPao7ygTrXwI9NImuaSi0L/nGnswXSGXDI+S0joX
1EIr7A/YGTvXwlUA7WnjEHGIJD9ZBUeeZEFvXhvrSc98HxGAXhIrHyzoUHk0pQBlC+my8fhzJLMd
gOERlIKQJrQRMGYeOVVDaenVrWISh7YrDNPGy21Z1KVO1eDBr2XpJJpXkJBj4piHFMQBJAQaA8tx
ruxz6ILUpr8HXX+Qnb505OU4PqfwWKpadAi7tMvwM/yF+GJknTUveQVpenRR0ONrPA/+3AWniuV3
FGdbZPrOLFMA7OKf1JAITu3R8fAOuX4eRhtB7k2ysBV+2tHJanIhP/l1Ht71q1P5p5a7HFfLSwcu
HYX1jJLpM1uYYIh4rlkl+snud619GXnnqR20GVg9GQLXkPci2lgF0epjvaBAXMgjKViqN18C2Jvm
TQSDoEsKpnGs1DKyRXI+042y0vocYHres5hB8dO4tBWaPL70WGZGawiqMFXU5Ac+swKMAlRJqiaj
p3XpiwsjU+ufHyN77jpsteyZGynnjePiwc8zhue8qSbL853qx1kmj72506hzXYB/UIzvsVafkiJb
5BTNVCQLJcZttOGOHhuodW3RS8tcLfXrg7+UXZo4pWxAMLLbJdXN702zSn8UMNa3Ikx5RAuTZl8i
PELbUJ8xZlgCs2NPo5lKuwk4Sbmzz4J2sT+VOjUlM9JWrhuQzCxNXfbHM4c08Pj4RfS0s3WKm3a4
DblDk0g3k2Fwa6D0mUgH5PQpXm5AcC5L7K6bSJqTSRJOGyOmtSc3w7WiU5flARQI26UynHs8M9Bq
ZuTtUHEMat9BdGIH7LTy3Hpy2KBPwaKhz0chN4SauEQ1eXqkNOWdvHNsHu9syJcspVO3xHrDzula
PIdn+lbPjNSRRCNNh8l28l+UqkwsmdJl4yqOWGqsjr5H+OxJD6C4zXNiyU3TFwtCH8pdzU/nomuR
u/+iEzxm7xz0qt1CO8drwRbAz4zcaUp/3/DduvO0QtlDfQRQJ9q4OLSQZU2LN4uHhr6gH3WPS66k
MFkzX4G6nVfnduX9rt++LbacgbUis33axPgVcDIoptHe+r7axMjQM5GRsxc4Aeowat4e/VfOnBrn
lUn+lj4RNzax9MuOOEl88ZHZbtR1CQpd3dRHN5IbZH6oKf+j/G1Su5S+QxZUGRCryaagIzxN4h17
TQNMFEXL0RVsezbRwJAexqB7aGxQBbXrsEhye82bSXIuDFaLlRoeHBEiY1EImC+eGi0USZHqHDO0
uWcln9bVPmu/CHr4O5/tr3O4ZgvUh6p9hrVugLYcMmFn9nv00Dl4Z8q8h1M2RE25zQx4xzL2ShFT
0WSNA5X1nWa9DSTh4d1h9TLtkE1W3IctSjygREe+gPOARnzKGTf7X80+WTbWANzb5LgmyE8rV2xL
pq68L/40O4eNGSX4J04AhXP9/lkpHHGvnY41GGw/R2K5+YUqWexpVW8I4qjZEWu37nV96eQ48b53
E9R6yuwb0B5E7LHLpVuLT5eNQ2vrlgf8mDAD7ywuxyFGvXFziGzo2G5qADkRb8gLvDgVQ0YsvESw
DtyAGGFS321Va4qW7ZfnokSeo2UTAwxFGNk0BWdiYDPg/QR8gz1x0Y/pCnodFD6eyZf3hA98PuGu
XWCeiKhiq2vIUV+N5tFD5LSRxY/Klwrlse8eTfB77jxUeyM786GnlxkqqPqxfmntNMB4YbeLOPjg
itlGLlQUUEdwPHlkF8o+BxxQb6UD3QcEm+huB4Rci2rKyrv1FU+0lz1x9vPuLfCIcGlpqZds/NMd
5OUNww7E1BUmNFeD2isO4DCEahUaJcE/143RKJnw7SG62u3tFdZOAw1N0QZaeNadDGYIGaEvRZia
aXJfhnTY2XsCr8ad9GBLVTJvU4Vk6MKJoMIonKQcg4TMlaSRJLJnyZju8dTsyYzDu1IG4PoNCJje
7etkud1VrMLoqSSrozZhCpa9vdbZ8lzJLn2Eb3W4MyRSZvKIQXMgxCNCUw5hcjKkHhJ1xGqgP6Wz
8bTf6wqJnEwTr7GxZPA5J1Vdso6tsMZuiQJrvvQYiXpN8t/sdrbdpmZP6vuDIG8k72NZmHgBydbs
lUYiBVz1mUS4mz4BW64b6ezYdESuj8Xk+u58v27u4atIG5G5M9tniQDuN4cpH9Oj6VG7eQzOhdy0
mNN2RYFCpMPs8dEybaZmjwCGYoRvTZXPzF6o+LeB7mO7M4l13B1Ts2nMHxcGFp+BVp5lpoDWEqRS
3XJrrQBpOUnKDFDTmM93jPdrrdOBKS27zfZINC2reJKDiVNrNu4eyDf+x14XeaVer6bn1fbcyDKl
SY/zxFmNn+hGrd/IQj6lpw+7XE2LyAS3G+tl5hfCKBoYSWkRnOEnwy7P2cC7AmJWx+fu7L7+bHTA
AK3pg0Mf4UkErofjrK+X9BxP9qBWBTI03+14S7IFPU6vyY+gz+Mjj18czjSmHpe5QS8JNf1XTZzY
FneFeK5AKSXOctPdgDVGsiOxKlG1pAPM1CI2B/nBPKrhlPVcF+PnSlHhpK1mIM92jm8LPZT1mPfY
rUX9B4Qpbdjdir2j6GLDEBODf71wt3zpcraZo5loNb8IFo0a1kyY9A3qBzLGWj+DwBASisNGZRZW
OZkTaSl7zLCO8pMVnnnXltbQZhfzNbbDMB/8uYnbaWrclaxdNZ5ww//N0BU61eQ/F7A9Oc3SMuqa
TwoEwBkjpG3L+MNELxVjnl1hqv608grswZzXiAGDOCGvPBABS0eptTYWGy/SDrffVcOLTTyg6BnF
drQdSjd5yqhi1TmGihY3TaVOZEqFnQAjH3xIixU/kZ5S9O00Q5V/f3gejRBw2xm0E9o7/dyWnCxh
W1AyVQYULNuSsLDXzZ3bPN5xhilXNJU+QUFh5nwzrcx92jVKIQO0AP6bpxqyWVuy/FR1l1kPteyg
5170/lWYd6V0LpIyl6osw1ju8C/SUoMZdbw6F7AL4TaEHSHLGzpcqaR1zP5+ATyQX6aa6tMcrTaI
DAU7Pgi2aUQ3agqmFzSEA5KJR7sHvN290gYHtCgDjBXRcMyMaklhfcs4Fes2DnHT6vgve83gIAoI
KwLntpOiQit4nzkHF3/WJjWsHO+mWOBrOsWpiTITdy7oq/c/hyfTRhoP0Y7OYgb3/j76AnaJWU/V
TKe6odEerd2mrQsWDK5WpYxM7LHu21YisnE3Cr7+usfdGzRvQWW9JOtI7HMG4tvyoeA0nETbsZWi
tyZxu8vfsU4cA6zeC5spabqtDJ7DZzoJPDoWNoUYw1Q+poJiwJUQvinWuEu3Tot6qhA8A9UhruLP
kmWrJZkTAon2pq1IF5sEr3rfvPX3drdhZNmNxxXU9YjbI0jYkzGxZUps8L1SFcsSo+myQip2TLFT
WfTzpe0IecUFiCXb+jAt3SDMWliXKMkg+SvPJ75A/ZqpRjfYwpV4PhZDyiN5mMP/vQ9bD8UMtpVz
5XcunGWWZphY1+kcOB72lReqUcbL+U+Kzlmo1w/gnMUt/QyGNACQYDnoX3Bj+WA9alFCscdxbk3V
AxAlPYsgVslrFseCO1VmuMFHkKD8dRgxWBD7MDJ90pXcgeXTm/xMfJo5sd7XeLm/+uNQHRBvAalf
hZhiweMVHwkfH8gOmW+4YhyuxScNWEVAQk/9o0Jm8h2YU9uUC/s6sb7zFZ8Rnn4KvFoTz4JpFNCX
XYL6vP2RtZMvp1/2ncADGirShtwuKL6nmjieL7lwTWoLiQTokBdIPO/fv91IH3CPQGRI1Red1U1w
F32SRJ/m559cJfAHmeGf81dRpVaUJb/DOGAwJ/ycdh/BQHazL1l3xe/wOrx+WSmULowwHolw5Lbp
5WvCIqbNSjXKCDzJG9bR5AzostPL34oXTf0m0UmfwYh0ztQuKWi3fgUMLRlih1WBEve0Gm8hv8Mk
NFADIcMzrAJiSHs2cDjsMUkQjzBqH+hP04uqB/uq1FOa8Y3K0cLtmn1aCf/MorEI4f2rnk0Ybt7i
oGLsDZVJbvsesPWdMrxTOZeQkcZHbhyPwpVoKBf6pbL1FG15s9lVChVvat/EQFWvEHRKpoV0KgA4
C1Gj0eKq8TTLxNq80NCtLJrSupjUowbvnjsuKbES03zO2G2TiI1xNed7LcYtnKgXJGntvcWPPmrW
BYOZaeHvI5x1gplodAyXj8/OibCDFmb5l1DfMzQR5ykOpXQCWWwE2rIZHJhTlf6kVuQcXOibG/lW
8vCiCC3BX90r2ktw6KaleAOvz+tz2WRL4F4NNho4UPa7+1Wv/LUfymY7RbRrRcSQ6Wm1kHSuMhmk
k7cq2lRZ46De/Vef7BeYZI2MzB8KSbIFM/jMUvta66C3ZONDSdu2GzU8hcX/cXhhNGK4taIM3acM
vuCbqEFQgCEEfMGJJm90QSgM00Ja5HhraueBTM2TZtWqwTEqNvuDPdymO7ZQwF3oBCyInd+lsukm
edl0qc0uuktw2kB2ZYp6e1qGE6LR4W7U/Sq4fxrgGWoWDQkwNU+dumr/ozPDzoygCjPssE+nu1I/
DWqUQwP8Ucz6srjRrNPZNu7RxJIgVUuHcc6+MDbGFc3xDCll1/H6b3cUYyjorBe8ARMnCEM2CL4Z
StadlYjVNTZleZLE/tHPRi5/D8Ik7lEDxKiVojM5eVfXb7Z6rfIIxs6gsgy7JQXCXDgyVdDwefh9
bZ6uIln2dx7pyZFDZl98KnU3o0n9g7wx0wjTrVJQ6dny5Q/wuRD8FXW+1mbT3gRp67MI6f7ehwn5
/GArmBQDr7T5LjnaH7Fx3p2fvG26ZwjV5OTdwFfJrapedYMNaeR5SfWP66edkjFXV1F9grZqUA5v
vU2knoKHQtT7/g9ienPbwWuvxXX4hqmADEdaUnEeZctpfG2CbvRP2dxr3O/Hoy3R9BKc9ftE0NaG
wmMZzJpRu6EnSuJsd0LxSZPPcf3VzqW/PiDwXG8ErJzK6YYDDFdmhikBGxMTt1KEXOUSBSbEgbh1
1ZMiYmkxrpClB8nhO7JrM1dPp/N1hcrBKVNDfj0Eb4KCBNSyb4vegS0tTu2hl3nESJM4bDo9OdkS
KZBqs93NKIcYtSTMzGaDxnQnXIbvVL3RmxNw6raAEzOeIW5ztySI9kvpIekkZPvc8gY9uVI2Hazj
mYIehBShY+wVM5gZfK3Bcb/j7RsuIueaoT8Z7v8S0EoEZ7N0/dhGrYqxhmqED7lPdeLzZ4FBqfgK
5jzKiNQN2HmdhthgKMA+XSGWWpXbtRGSeL7rvWFhcJJx9c9dlic92U+Tz+WwIRsVznmAjSa7lSg0
yoOu/QSWDLmWN+5ek/jip8hGm/annZDQ9pQEpbqTdvNJ0Zcdk0WtfZ8etou0QllQ48fPpIuhGPVh
b3Kwttz5CtxlWv6Po5aHtA6NKnbyOc4fV7T8P9wL0e5mok/hZxbcVNTR170OO4W0P2s0CK2wE6o1
ODBWvIz4DJTRjXbztsTVJYu+HoWVkC9v8FRzIGt2Oo7whZLmjSZOt9EqatVx0zV4pZMEAzuYmVX+
JRcKMFOemDg1saBzlP8wl8cToBKzb9ABORhIW5t+woCZFOPGtmUk3FpA8iCts1V3qqo7fpyzZcyJ
lssZupUZxZikyNy15JMklTii3wcAWqUBgg1HD45Gur866PYAA9YchRrJB+UC73+avJ05WUhHQYhM
77nG04uRf/DTzrGqFMTZXK9ebod/WfyexxVFQ7blfMQ6NJQglHKfdkGbO25JteJl6GkDJ9o6im+A
BqWgSbW09S0oCHCeez804k6e1pABk6rrkgy1RnRfe7ru5UKQ2AXxhsq8hXBi87w4u0VOlPm6vxZL
WkW+U/s/Iclo0z7lfStay0BwgK4Y9YPjQrrJVGL8cMfEDq4WVjsdhHTE9TvcfNP3Y0yHou/TtCQq
u+Izi8L7jlICpQQm0iMIv5KdgpmWeETLCE8ofh8PK6pm0pPxuX76ZSYJzMn7igAxIyDbRmo0m8sK
1YE6JpscSjh4rYkVEV/BTy/1Si1YbwhsV5URYEGtbvWAbSy6Bj3QPo8QInf0Bq35aOBzRNW4iiaA
adSuhBgVt8/kZ5EgmN7HrHaeB6kC12gNsXNBZXilMnzjwIzt6A/5QgsaxJcrl+wuLFYJDwJMSkD2
RXXUH1MrLEdhm66NExypXkHp+vAGDdILslLmtj19eBctVbanz2k3m02dvq3wa1yy3bqatNIpJiRf
fH/TuI+8GDV7HkKlB3dH/345Lfk1IxWDTp95WpPQJsVv0b/qBKewucabMJXZL9PrIjQ54KEEybiD
wUp7ALAZXFToEuvbAd/Qe9mHkH/jmG6rrEAw8WB8pOwl+a+C9DpD/7MQ4Bve9EEQWkGgHNgKLfqf
Pt3DsiZbF+AmgUOykhAvSIy5jQCliC4WgtJPzsKscp3vcjy+YY+PCbhLMG+vjwwVp8tG9xCQZE0y
x6Jxx5Z0Wljus0XNe2Z/+pyEC6x3+3bEMq10uQBtsWwoKPnwu4FOLrM9ttC1zYct330SsYtPMSs9
m1rFWPsOeF1wUInnRvYyHNTDy4pUGg/tc+f4ygUqOEra3Oqv7ME/ngulRi5YRvyB+FHoVTe2pf7Q
wurgdMVzWWEX5UbhCG0X/kE3LijNMZwZSNLrDwDa6MDM+LQaUf/Xan8+durDxcE+q36poWDT/uSa
zlMdyxUj1uuUrjRoXRM766SmfcTAyjXNfLbd9mkCstytvT/qZEW/yFlWz2DPevpOJ8RLdmljlaAF
UyvP52/3SV3u7b0xYTCLTgt3ln+nLFt8l+XWHir6qJHXLyS5K6npUKkW22aMqS4vFoWhneSahSCo
8bcsb9zMD7fydKFgpPGmEUg2lQZzK/J75K5AuC1HDSCVe3GdWZEsNtVbUAidDTT4IMTz/oFqjlc2
BXw5j/cDEzgnfF0p2vXadG75fASRRlXIXsZi319AJt9MchOEbMd8I1bPRrM3lKIVfvAcHLKeP3wi
vW9ThqIlsra5o6VlBaFGHzjvL5xJLOt5Cj/G72lgiT0E08TvjhlR36zW8aRNpDvxZTqrJgRPAk0N
CurJJs826/4AC0Bapo+IlZxp85tBFMxBG8TBqJXJXSUp5VN+lpWDPs6RY+4dRm2UjZU+GHTBANYK
/YzBQDYGzx15fc9OK4fhpoKFjgJxVNVuI9Oo2jsFUMRypXhcMUHzGkuQqm0HfTiNtK31C8Ex6b8K
2pubLC/5Zeikc1Dk0WVbSr2flJhGSKrHZ5PvbkYraS+Zv4bS+32QXBvpzpIZYD+mVG5t8HoqDJX1
fxeXC31JZ2DLoeb8bNzM/g7ediZovURafM7tTZ2mEC/KXzyqXCnHI15hHVWrWG5CvA65cGqk3rAp
nA2BD+H5Si/02OiFthAkrwmMPxH4nRHwpqlVzw2yQys8+KPGN9Q4VRPt4BzgNGjgUDLmmY4l52V6
vO016c9+754XAiQS38ZtCDB2A5kWwPlodNTFvnw7wKPgsGqph4zaw75VADlB2Y4b26DJaUFPk6sV
bcG4MkoVsXsRnTgAB/XKNtt6swzjwAMAdP7hDMpCVhioHMLdc+h0b6pwkVv8VBN9KytuxC8Kuhir
qWYuEcP9/Ektx5ysXuJlZI83N7LV9sxGueVFuD3rOOFku0/o3kzM1g5s0VUbQA6N3Au3wOJyFJIA
vQzBMwKa6P9JbREEHmBOv046BLvHkAJAuSUWRWcSz/b0Ou/MHDrO+gSFrMcP1iT2ECGdhytVcoSX
xCi9o5H2Ew2BQJ9iRkk/eTvB8rQdfyHcweAt6YJ/ElRFbWJMH2EBvVv040MAkdjcOlZ/GQTRIRy3
gkuTjTa0QSxE0CjZ1rFM+LVm3nyda5urZwfFlifntdY8ASGhWg3nfUJxBbngZ9JGKCG7RK36+uYv
Ua5oZfzQMPFCLPo5jRDwMHd/4sVrDa2oZJZmPGQ1kaZPDtW5uLh2bOkx+fs3UVOpyu9bmWJxxYQI
THZYIpbBkSQkzHGcjsuy6FzeNJ1hiKhEtr8ffwP24XYAnttTDmv89hLKSR/HNcwJFMZ3t3YLuCDK
psqdYomj6+ZzQxA9pluYqdFly2qauG2YnWSW+DC/W8qxI5GhvQTgck9J0baTTWrtLvJoINPfz+mZ
r3End799RrKXMY610jYY5y4buX83Tdbne4JlnIEgULzeg/nhDrgXg4dbsKjW2D1+5K6XC4HWrsYI
fqwxSGUoIsErUVWQtP4KLDr4ras8sOD9LXmBVSpgh7b9jhNtrxq14YNKSGcPK6FO7siinit6MTw8
zWAYth1tUlb5GCzX50h02Dwk9mUwDJ1C5xpLtqkSjFXLWLC4vZRZ4RND6S4OS4smSaHx5KRj1PsV
4c6BbPoOO/d6Cwxd9/MXVju6VZkTVxQlVpyX9aO8AT4N1El8PiIPt4AMxvI87DpKtHTDADYNdCMx
l/Pj65qiWs8c1rXONwT6/hTYBxfSHIuzsX3nxFQ7/tkI7DPW6zGqlPhrn9nq52Mrs+dVRNAH8hAV
hdNbo54MPm8cmznJeAhfAe2S9biwGgFaruxojkekvR8nExx+qBxR4xl8KEwMT/tbW8GYPRhs1KqC
KDY8szGN1HXVZXzkP1Gs/iWA+7xED+deNoD5w1EJgvwNeM4FsCDcW7buaD59VuVLPLURiy9ZryX+
Zfcza2IXWWF8luoK5ZJEWtXFOK0YDTYW6LrF3BPXy6UMrwftWYEYVhF9pU+hj8xsMNJsFGEdza13
HiN4ejRW8iLMfz1Hyv3OX3W1UpoE/FBU5VKhq30Uu2IiR2HgnD6bK1S9d/RSdVsIvNMA35sWbRwM
FDP5FjAw0HW5HQkN+J9fqiiNnd6b6r2vavHscEfIQypkVrxvYULRfJSBXDyhnYUJBri/Qaq1xO9+
Eti9uIGRfHPXFSI2j1FGb3WsfDcM83aQBrDpi2Ra8pKmPF3S5S97T3Jp/D8D0LX9K2lv9EP6fhfA
Dtk2QmtUzm6PQJO0nHAam/2qjgoYhSyltLA0kaCPV+s/902Z+H2KMBebU8qlvzb/Pp9SL4GzF3lb
01f0b/+0jn9teeenIs3cZPLozkwfvzqefWBnSDZ9ALMKMYNLzq0uXZT/ST7V4weK2/OHwdZUqDlE
DbDCeg4qBP7L2zfppQIkdZq0lJRnVmFDqtIH2RohpyFgHK3pb9klwmMCaTx0gU2oH1BmwVslyBIZ
sle122eNZLi/wS3bPgtZh3dLrwG1ynS0rLUMMVdPPZVAn+XmH8ba4ioXJdVKOTM97ER7DtgFuour
YK6GhmegOSe8UXJ2ZnC9ddTxOAd4OXU5Mfj1vqbKpV3fLtRB3BUSA8vkiFxfAi0NT+hkv0cSbnpr
ttenaJNht3KHSHiwJ6AULa2a6cv5L8swXIq2cbLJEPSuFE7KFrlGv/o/amFg1RLvTd1EiPTWt5tg
iGvaF7/xwyramldvZjOPfPOdc76+OevUNnIFrRpACut8DcXF1kmbX2bbcZjjJBtcoccooDdgROnb
M5XwbkKzl+GJR1DAGQ5Ok9bBUcxEGCk9Oe5d5DP/47MFvt1lPEKQRb13yT82/YnSu+6wlUiY1CVI
hDuwKwWwkPQE2QKo5KWJigzWPPNq1JJak87EFdcAyqxhzG+u3TdudL2v4GmyP1Wnz0lGpWFlH40i
3ApIDAiCQaqy0uvB7cIGbMObAt8+i0WYDUWYLgLvA95Bix1weoyv4qTsC608xbtZhht9066YMVv2
l3whVUHRH24OCkOU2ffqVRT/QfXxkeBlq8hznxsM85zzXgHYCPIhHyBNprihBO77gc0z8YX5EX7j
HsQUfDMsXYfB6bLzouIuA6UeBxRvqhoADUVTRORwN3+Uzqb6m8O7hp34BVKcITC15zdnTH1Voh2c
jP/PYCYkjmtgbwhVqZwMDfj5XCG9s6Jaa+wzk0b6L8pAr4datS9Sz9Cdhx9v8euFohUPpOSCz/gE
Rxx/s5YaSE39oXLYwEGPFdbZ8W7iLH170t6QWAaQiyRa0ILYyEwa/66pc0eq4a8FV2SgY/P5WgbV
TweUqTuraxmAYjnrYZzcW/ih8qpMKKRq+ZKiWFSO3qoKBuS7j+JfgXFhR3tO9kABxOkZ4ftNtm1H
A48IX7TYMM9kgL+fQsqg3QJbhJIj91YujKWZxiGZfZh2SqqVUd69tN4rObR+rr2pTyh58FJS/ihP
4nD0Z12fQySuPzDAbt+XTjkC+SlqdYyQgkYWp03T2M8Et2EsAgfL0ZhWGNuHZefoawpDINgrZ6rr
bsANTlBGyZDBlC8tRITdgJqEl1mjnXCe7KhLED71gASJ/hRGFM9gpoY5KnWOuxDLqSb2zJ675enM
XZJ1f9dvoyuhhVJj+fsapczuSBY9jet8P59FDkORvGlsYNmjqhIbffZmzuJk0K0SxAAJDdLYxZCA
5ulMkDG1MLzG38frWrxZKCIypLJu2dcZ2dUyPn1/KYI3sfRyw/ucLy9xM7DC3/BXiUCg3JpFs8pd
+S/tZ4h852h2BvvRLcMumtpNvGsA8fzFtiO4Y45QW3hhWb8iYxxC+Qfon2ywTNRe6aYBFAzWkMzq
EbA3+6jjxZBuNFzI4aAQUjbhlMx+1sOW7+vNnOWzmPLrF8qjHX6ZAzQK3QrKka6FqrXn4jePf7AZ
XaWUk9gBBbTmAiRWr1jTd0O/kKN4skNMnZAZ+WkMIhjZrPD+67k4L9KDiB8+chfGWcgeS6pH/kd4
X53aNSrhAR2y0WT5YMR7caRVA67ixMOaxAoMQEbLbJLEO2N0MBAy4mh8LU6/9KhB+yyPnnjcIZpI
CoGufLZ/C39Z8GjnhqQ1SrF46rL/vONZR2QC9ah68lXBQTkW8xlyL/SoH5uBV2OsKm8jLDif4+E1
QsB63Wxm61Kr4PpvPMdoI59AfG7jINBy+uWELMZPC1+ncuf+LKU1MPbC27xj0Xw+qd66Hkv3tlUH
yuK+/Ioy3Uk0ObUZgUC5Yw4VDT2s8J1+0IbO+MDz6WwOy37j8SX7hfguIb0JlJd2dfiaf7d4xv6q
nj9wOImlZpYhfa7YClgBLbkb7MYAvalRipmGRZnTv/1G4AJp8+VVCCtEQfsjazChH/vwQRVdRId9
UsfvXjyWbiEU063mv32xIPWXADo0DAu5C/pykgxOzjlFBHO7q+g86b+cqr/QXgHrNMPnjwWeEZbq
04PDSKetEcJexfbWo5R89NlKlrsvF0ffCXvowMuow5zyv9jOSo4sQt0tHufuUJymajkrq8SnkjFJ
7bJ/Eino5st4+9eIAlVvGg4phVp7YrCIbgp0RxtbYuAFoU1UyHJQOEP9NUpgv2aR1MgIsrjrq4bJ
jObior5cQ4lAvQW6GuBRmhPW/OXxUVwLriGYZsL4+gslnEAJd3OTusjc2on+cVl1wowq3M3AKgPz
GJqYEAksZeOs1iGWnZ+Nh0mXfam/L/zV4KEz8QxPrNz0N5X6yFzG7LhsljZfdJ5/uqqJ6+9A9aaU
Si7lq7zjjODTrV3GxXpAjY7xemKL+0ToY6vqdgQNg9X1Cl2JH03zCL6oeJU/EFicJoLMmtmqYr93
2SILv20WwgAIG1zUZAP0M9mmtIhS/bOH4CEJckfBueCv5XlG6IpLP1UgSuDzBVroYqi7eH50+q9O
8J8Et2qSl8Gmm8J7WYixDHR00w8ec+N0Zze9pUawIF0l27xmo7F+iKQiqjEPSpO43a5iNegc7g3c
w2MzwEE1aaCEnkbXDJo+5WYFKrrmLdys5BzsEFEQLtQHpFr4Ic1yBwMgh/q+eeMDdYjF0RQKMXu0
Lpg1X5pYmHOBd9ZcGofUyp3t1RN81hURKTVl/itezArlWvk2osq5SWMxsUYjEW2ZF+x8/+i4ABlS
WvtgcMJTLaFBm12TpDbnYH989KUzl5Wp/hCGzQcuxLLGKj8eceMuD201Zl7ZIcVjBAanfJLS4DJ5
a43sTAdpmPK1ZZDxn/1o7luvUjEqJAiNN+qBzYUwQ8WEndrBdKR1uQUNIPWCWu6W8gIFLWfNOH5i
JEId8K3h9t4gnVOJeQbjgNbfCMfpkLMfipUFIYYbYojM5s+PX70ZuhPcBMV04YdYxkTu93FVGi3K
c1E8zqlfVCe82bTgf5fYeScVt++HHNM5ifbjbCApQ0LFLD17XLwfP9MfzUwhkepqL9/Ud/OqOV8g
Lx5cpPja7KSbg9mTHccr2057bg+ND8lArvgJkFqFOM6xQHMCFLhc2KfUQM7iyzosapetXPMoikxx
VDYusvuUknCoVFHG2jJDhlLFUkULM+p1YEc852k7JebLUwdYAJHKdfA8oVqSuTGuMLuS2jVEoSDM
ZOHFERiNdNy7iqkxQ3T9a8cRo9ZYvcnLsJNYWiV67VMujnvihN1fK6hIDCkTfkPDdnKOUiIqZd7x
f3skBTzg+KNYk3qm8i+D48vjJZE2GBypJJ2IajuUcw2nK13gl7sMRO/sQBhPnYCKSF4R0Ccqgxwv
maHHhpnm+SZn5w1+W6FikJ51ExjTGWIyFkjX8AUUQb9uTfCoctOnguUJ1vYEXndupZBPMXE4sHQS
3SoSwGi/vmznBu4MK900L/qT+ruHMFmDSJz8d3kc8aF+ywiebtodda577bg0V90y3JIelh7medMq
Y1zqxqWBy/46e7pa9ZWn27J2ejy+ADWdMR7ONkCrUhtt8VNczbzCxkucnYeJuL1Y7AwW9vuTVhBI
CiZmZq4vqfVHecGSjwQWRgxAkXC8Wghd31maTrHvD8VQRt4m2waX36jX3UxeWS2O4zBPaJXz8mDD
r1MrjZ0HuqVGquQRoUgsfwbEipVHbnQF1dRsiGIo4PEQ9q6Y1fk66eZjFATZU5RyiMnwzf/ZuMdp
krc4CZclBtNxwlgQLp4MYmHkgQSLpkziZCKb8NO1D+FiLi0ESrIzDqQHdUCkVSFV2GWpB9CC3QXA
MVCjDIfFPbTZnL4DzBM372qWtNEupPtHm+UW2sh9wsjv76FthWr5MUflr9hP6VtvwGr696I6/oFa
d1YVDzZvpYCKyrbXazxdD1UFH+ETfZYbi2CDTck2jDUaVYvCaJBPWyMh6n7Ti/CHH4LdDUQCIhWa
Tq79wVQpvaZSHkNlolQcBAhH9HMjjby1iKbGTO4LtTLfLly0iHuZcSDnDXIoxxu4BlHlcKITJYAh
1RGzqYvzm3Je6QCB4oLVbwfV9Z4HWF/tEJndro27vG44lOLmAIJXHQBzEYJFb6KeWGlwcMTzT+zw
HySSNGW7k9q4fy8y2FKWna76/9BdUI4TWy3mBcYdoASxy812C3UTZLjaZRLitcSerpsZl8eGWOKs
bZCB4XMBknzpQPi+cA4UAQrSKJLW7xjvr/zUb2qPq869f7fygLwSmzDYRkcvlIrWea60FXvOMPWk
AIr//F0piIE1TkyRFo8OEs1AEeRBU9xYEsnzdWaY8U5AKJydZwHG+pdmuwMeP6pEqtmBNuYs7BKd
2rz9Yr/FbAWB8x2kcxoE9JTmFQ9reYNccUYJaqRZNMT/K3PVIhqZLjYKVFmaN9Eec+tM0s1q9b7X
JlF6WZOCnj5/tHHYb7guvsuY9jGFB0X/fnR6S6PYn5SO0/A23cSm1NE/9Ag3HGXSLHlELsP8tgKD
NNzSMhdHjTZ21ufVjo2G4t/klkHUlKP79J9iTqRofzN7zrIpp3MuMzwrG5LXrwW/jPQKsNqFxiH5
sP6+kUYguldVk3RKUKkFnb0A+IhrfXJaCe0RtgFLVhetH0W+l/Ba5ZoFaOV2V2hEh2LIYcGJvOol
zjU+2+2qXgafQTrYrI8qJ0iy3nxDo+W5wVPIQql0buyZS2fWFxV77GJK2VYcz9kQHPkIcmFg3Ii9
zW2+UO/2hmPZZTxF11tg0DfjGAtcNXn4/vmjrrhDgq65AQMp9sqYWYN9GCPa2kavL/dg6Ktb+Aop
W2OEgIoogAmuqJQ1PLM91sjPJpRabkWYFl1MVXRar8U0AJ9P9kHm/0P7DNC3RkWQvZplPVVydDkA
kB4cpbPPq+CwSlwxnS/wcrX5O/H7sBajHLs70t3BMM/r2CMYKLuha4CsMnwKMfKe94zd9+A+nMRf
gnLf0o+8hnnspYSRmIKbpKzzbgxsIChP7q26crCGyC0DyJRgls/wGK7u9igacTQ1uXEGEBI3vBYh
b4TyV18HhlffkqhXQnYcVTv00Jyj9Qw1dhdQ+y+ZRgaKas9gPkWYp3DIS63Iqnb9pbq6ej466DBF
bsC4K1ufLUFf/CYzTAZ2e/lGKOHTIamMQdrJtuK6ZLX346np+TJevsSLhC7LFf7Xm0bl+VIMT1WT
+qsvm+Q58wGb924f/abEQrwkLpoBmyGvCgloXTspKgZ9QVrmSZG7peELYMwd4qKH3xyCk87dM5E/
lB8UTPs7+YcgJZr+LD/g+XP/9SHQQmmNlzgcFRSMwuywfD0LX4/mf5b4wr/bDzz7y8ZgEjN4e2c8
VTBm2NTonHL5mPcT1XbfkS8aEPBPQRLx79Lzf9A9bvau6W4WwOv6Sr+VxMPDg/sLOMuGIaEnJi1a
y7FAexo7uGem3ThegtMWRCu2qrFI0i95RcIHzop9buqo0sEKSvfnWmBG8nm7Ud+afsn1nxmUJXbl
4O3jMjmYiN0Ub0/6XH+goLQlyNFg9ViRYSX0JoTwU1m7FOw6d8q6OHdNBC18kndP53kulpvIAPpG
3R1i7ZRsMEDjgL/Pq991ajNQA0/wVqc/WUh9lhvqYX24E2brpVPaAZnnsLizyUOjsnR2qPCUSX/c
+bKhnEJf0wGRbRydSKXfQfi4CqO8oxKWHQriI8scjtY9mw7FjxtMqNNyoTJZG4KH8vs36Ceo4ux5
6BbnkkDrjuq2BBLmQ3TRM6bKc3+EXwgnQInNw5NL2Bvap7u/bJ3hzJRb7bCobLT9mf/9yc+Rpa7n
CJQzOey8BKBKcOyTBY5H5CeGfJ+42fx/Km+8rV4uXtPO7NIQof1f/pyM4VU4gDH6ErIqYUYCfsIK
6mVkfbaWkIGnidVhrhrykWF+CBDDqfMmgkZsbTje8eB/8bCZ14UpIDYT+5U4rd/1ymgKCu5DpzNx
8r2UYkL13+WCozfmaPdWjl8UnFj++DBREsdQUkwnDbgt6aEf6IApSyc6DOsD2TEujnN3Uel59cZX
ibso8Is2AMlEmxvtmhW5Bm91UTxzuut+gBo2TKY7/toQuoVm2HG9YxI+AS+x+jeMtVGNrNiyXxO1
jXfqlVXh/LVThK/PUS+qf/9yzMCBDV5L3hDhlUs5LHq634LMA3wK+vzFPBj7Q4IlvcN+FOihhCzv
JYkXkvqOcf+CFhLDiMFmwpMKAmfNMRHDbZLv2mWYMjhMan4K7vzvamBWmfMvpRwks1varFvGPOpp
qxS+giFUE8nQPykFICS5RXNbQtz34iOsM2CIbrJfqUGN1zC4WGQhC3lXwyjXcwkejeKlxWZeL0sX
kiwL7zzZ7yu7WFfHGnJ3uWQHlWobhxJpTYZwDdQq9hwjnzgw6CY0++OlPhno3TdJv9l6eJFiI5SE
zzEe8d/5nZKJ66TFUQk8HnBE0T08SqvRuLz4NM3umMA/2qsLcpPO1Y8LjcNRwAwZJPPr6Jn3aHWw
ZyBvKNu8qIWcsMsKk7JGJSZtprlmZSWmT1XoAWaCBgetv4wDx+CaWSqQ/lgFPLRE7SXU0schJ5vt
Q0SBHkI/E+IGNJ5yqgNrYgxl0g6biTPstlv9pwDnBYFU41Pr2oeC93aeisLpr3POkwy38qgsvLBy
dET9BfaxjSFjFf9N9QEx01/JqTtUcLFgO/0mkEHwb3hiMyS33B+3wS7yvZTHXtM2dUSONVOl/wO3
gxdS+e9R5hfSlTY1fiFnKXE/ig0DajwSPsKimEr0vXXK6vN7OfC1r9PeKuYZdq/2iYJxXKqz04Sb
Aq0ROg1Tn3yn4U8iG+qANE1I3rvTcXdxkmdlOxqj4KDs6ygTvpPW37L8HgoraKBOH3w7OP1h8g7b
7OGyEMCoAXUGwchR7RJhvOkDFpBfcCZJ1gpBs6uzjBOxD+/nLx3diOt0giyNUSAmSG8Yo/awGb1S
kd26HCLYRxlbHifBFYCLxkrr5cwiZ754ctYqumEW8uQ4+nAZvvHdlAbYigEn9046qpeE81LkPU8I
Ob+vlBKWPWOF428/6inp06FWP/15ZIsra0it0Yq8M3DZXuwndpPfTv/7TzrqRwKUx3SNk0COO6Qt
U1U67VRuj+TZFkm3puCjprwpsJpB2tqnTfn8Oc3auM9+PL4DeZ5PqwQbKjDreGbaE6EXFAbdi36q
d2xEPUojiPpvJHP2leqIdj2fU5pQLJT+G4T24BvQB37izIbC//PKoYXA/rUaCzQG4zyxuQbSRUZM
HMXQUZqcDHEbxFr67G2da+jPqKxzArU7RKehv+P5ZoGpNwuFWgz9esD8lieDZSvbs5yorGZLbJ07
ALfUjkWXgMThW9quj0IsL71fGqXGaOAnNkVx/27MBdEWbz4oYOvQ3mn2GoiT8okzX8339iinLIzG
pgpvVX7aq2l0/uLNsbNFX4M1iq5N8UgZBEtvOm8UG5Fdfq8GfCpUIHMQIhkj5vmRB0ASMnK+7oVH
M2ECA0O1WP61Ko1O4/NCHWSnOPEBaqQl3nxv0JnSxH2Sg2NMemVNYUUwPlTy5/q+daQiYSaDvi/A
Yg11EJNlN+expPK5NQUFGyYMkL8hobdDngFNtVqp+behMmt+JQ/teo1sP2AH2C46TvsukubayXPE
WxWRwS/4bgDikXLFKyM7VCTrhhNORdDN0/z9olsxl8uhs8VK85XoJOleIGJnGGBH9bMFoyuPc5zi
a3PAnqZWzXY5u8N/J/HQW/ksQyC4QiLtBN5XjGvhIWDmHimyyrXNHlPZacJcmM0RZHdOEAAiPxTc
wsjStlDwMk150dQA/javD+gt9VkcNvP+g1hThItXtiXS9MiaZvU7YfjibA5MmPBNtd0b0alFNFoJ
SPWap8M/DyywGi6Qg0cJdpkh7batngGEMoz5NeHUK8GX+aYweAgWJ2boPYfRbGhnZQeFvnUkY1We
scQYHgdXQHz6eFh/mylfjHT899UmsOX9VbIFtMWRpQipMNNqyUtAZKiFK+hbYMlWcX/0R2/IJOo7
5j8vNQeLu8ucFPldgXoeasx7bnzp/jZRRGugUdPiUZX7ikq0QRWE/rOAEHM47QXlL5zzwozc708U
lf47NIZiPlS/aucZeNTG01MJbSc4vqrKeEwbOLPepNhOBusPQRmks7ciNgY+J1QicoQmLqUEc58E
gZRy5w3VgiBQzUM87d7lmE6Qzhozzmj9+RV6yZNqprac8ZdWP8PGesPYZFCeOyNsZ3Sr+UVy7OFx
e5EQoBCFp/TjvLLxMNESmFB0s+zhaWBNT/UIj07EKPo0QgHqYikJbtIUfRtqFXVldiqu24PePz6C
780akn1ICTT2tghZ72reilxLNrpjcASjbGrULH3zVgq/z3KJQaUggtlRiQYXPj5ChVjFDeyS05+x
VjawImxFTboSlLBMb00PfhXSe8Pe1PR0WzbwydQhkYtCKQsWM34iRfLqL2ZkM6nXYIIKAM44a8av
weUF7nc/2kXmRtVN0UBRdoD3UBAdY2l4rnqTa2RctnzacHk94YbT3pY15jyVyI+DrXx4E69DeCIP
+YUzPjZuITWj1uql+zpdKWglzEo1S3M6n/9Tf9RZt2ltiEKl+PXvxy9ap4RyIkfO/3TOHxxZnHot
rL3yEPaStYGJbPZBQNdbj/cuoMvDoWZAKsh2/N5GMMI3nr/97/g1lo9K/6n9LNXYbRND0Xxf7+eX
3yIZikCQO9jkAEbSvF5FwS6yXabmlKTL6DaqKxL2gr0EiJAmLqy5Zx1eq8iYtVmD6WHPRNhivmcZ
VdYh56wVfcs/matn8FfEkVMSPpY6NfXB96wUmQUEx8iVnZLSvx+XlAM//sg5o1hCtRRj/oJPMOPE
hxchx4OPy6QDP3Gq8SXZRpiL+0DONPNyc1hY3TmvyyeMsl3NT/f9GTjYG/KgGO7mvHRxXQZFzoPt
Zh3bu8jnqVVWljdlwA6Y8PDHonJuW0yLLtcMTfUdgJVY9eiZa3pEvpqdxM3BHXvX8qZReDtYSbEX
peDOnxZoYb1W5fAjSgTfzbLWDKWB+EWYIzQJGVNW3oi04TRrORQVmECx6c3DX/jP4ka9N8CdvXnZ
GXlkrTcbQoobyzjoi8Qj36Xl8dquCk/DbTiE08+Zhfl/3fX2dC+9OVVo/9F/llwlHHc60HJD1pam
01xe7ux9nDhcNUUt8XUDV1GKtzdRqtn28oG9M7zhofasGCFQvg8z1en/rrvN/Er4rLZVT9yb/7T3
Ah03pdetfLQSdKWMoRgvfGKYchRfpWYSEyV64Zc0p4jae0NzlC9SpjEWJKFUX9kk0HrnIYep8R8J
sG83l941HpEF58S0z8tkUgJPZFkQt56pLDTAZVZqI29fc0d9lrbzOkw7ftH6VtWzG7ya8Xq1EOvN
/i7gFm5AdU8Ab/ykJbFhszGpyqgSIoLQCqnasZkoy0wuYYQG0Xpri/d5wE0cG8xlks51CAbIa7bQ
eLAsZGbKiyvbN7+2zb5AaAtLi/y6i+RopWGDfnLEbXSO1g/ArJpKN4lFS3vOwoBebthUK4FBSTM5
OTyeQ0pY2vXI1UxCko9WoBAlbhrATh6ZlVbycDffSinph8Uhn33GEvlxWFkZT89NrGL2z+a7e928
Mf74wPMeVHc4/Tf6MpR2ubhIjfaMQNkgYMuDuOY3qPYOA3CQBfdbkDLuA7Xbv9Zjzw09asdx+G0+
jBAQqniboUb2UGVtDlk76ygKccgcW2fEA0dmANKjqlfCmQFt7ozYu0hgb0MPIZ185Hb5td9fhzhP
G5430QwERlsottUsLrFkefribeO/KkcGNoKh4dy/BVJPy0YWI4kDkONjL6Qh2R0odUTo5TehQYtz
hYkVUtU+uDufJPU1bf6ZPF4kz5EkaymJdVkl2XSDxlfZBq5pG04bdQnyHjXox06b6R70eF1x89TM
I2RDxCWJap9sJaNXkPjHei5b2PwqEbO+eOICTLByA9xDbucdZcGkGVbITOjHHt4YvUHq/C+Yjigq
ya1t8jX+grYZjOUN1+zJGZ4IwsoYUkXkBG+Bn2noU86XV6Acu9kdDGyDrV2rQNQJJREfqsHt085g
0EtmxCn8tW5wjC4my0Vyxyk7jCDoU3n/rjCTqEltmVhtvJ+NaMJSFq7hqOKlUgkeloG4y1gSU7FX
kUGJsqPV4aS+iR5nbutcErqHxsBM0PKU1wmGcFWJcq+MzwjKoUJMH7iNfijupOXrSK2l9LltcQC7
JrJ6pJc9Kztye0iJUdPcwobe+RiPMfkewUd8zGg4unBPavXR/YfSoTo74c3OxQQUsixP0KIcBNYM
0m/gKOz5eQYef8Oh1SID7w5ePKqg+IMub4dyQhth5JEACp3m+mps3l94Ixij6hhvHA2HoT4mNb0S
WgzcXYxdcjMGM2oFODpfI4RqLFlfLz7KkE81Yo/nxujM3guywvEj5vizsYxLfZ985ikvfnw9YvVK
Ldk5Nj8jzivt82KaYh25l4y+JdBKfctGJA8qZpDUfUyzE+gjq8+DactHRrdILrY0hFMx5JBDNtEn
K4AnqEafH/b7jrIaNAo1SW5P0+l9EgzkSzPUsycGXGmqF9Tuov71I/vmsjEnfI7H9zDT+GjiBLwr
MPc0gV9MH2kb4atE68gplmaP/wdQpyoEqtMBQ9i1Ak0eu+kqZ/5uef5ovp36sPELxe+q9x3Zjxa8
nqi2RbiUp6zREs5cSagVj8krEELMI9Mw5f1lHugh9Fjx+X5KcKUkzWb591F2qCPxVvH3s/ZNfeGV
CdKQgU9rO8BOanaNpOWv82r93p74LrIjP4klk7EgDQ3wVevqX4wPwVqxPJp+ldh/gEkBKbc/hLQI
8capP88azYe/uRESvyXKMbjjfn7v2bmHz91WzgFqR91yUfIAi0rQuVFeJ2rSSzBUAf31rCupLOWh
T14DsiysledIYGDV8sdORYNIeDhtpvFnT/e6BPHLn7kfu8ilVjmvYtbiiDWAS2mhSXk70ixa0Z9p
1ygnJxqmzyVVPzVSKcVL/W7e+vZhUrXJrrulXHQ2DFVVwUHiPqZ1sYg6PCnM1/sOFzAP5/3KSff/
XCpJvG2gdfXxzxwGietAp+0ygd3vkbCx5dgJx8JNGpxXgCF4oQbwKDWnSRmS7RkFK5oEDiTkeqPS
/zXNm2OYqSMkkh2yv8edhn0dB4axltpaGfegD/KX2MGzaF38rVnXPrBLxf8mqi8KHcWaZxWDupbU
umrbmH5cBR7zxiJf0jf1HoJ23X2XKJjiRYn1gGkbtZiopFgciz3oQPv4rumn1ZlB5X4ooAsevZ/f
G+kE7hg5RbGS50i38PZxR+Ja9iYUGClvyZW+X1vqkH1gRfuwyxsD9EgB4t66jd1YUw9Y7ZfP59wX
DulOZPKEtrdsrl/Ah28Q851AFTiVJeaWqrM7+iO235QvZrB0CFqip2ZXWaP5OWQ1qmrgu0AL0oLF
DEiRymFj96KEcuQJGOhneMtyRohATS6apIkX70K9Wh91OsmdA3fgvdRGS3W/oBx9u+m0zMa7zg/t
BM001F/ewnLSoSYisVdsC8mroQEGTqftLPcYDgEUnWmBcqO/37z/EkmgW3ApMmS5nK8N7aJMRla9
KVw6GWZucPFlLFiY0HT113dE25XnFPibQPozjH1MZDixFkYEc3PMf6f5F/kqBZQ4GWYuEB/JQaXd
mjyCYrt1xDjPQilJbnQSbkT2LxTVTSS0YH73RB71he45CfwedMSh4R4VhDM1d51Duqtujnfzg3ja
+2XHixEWBmarOFpINiP9s7636cgz3OhS66OSc9ZYrnOW7kUgzwomY5oxEMGklDm9fY3jHSZVix1E
+W67Agt8i8KZTp417rPKazVnBvvf5bUpXcjfwkMfuLRk1ECdddxFFxJ+uot1DooIBCk8kUW+fd9k
wk72hHaV+QhuYUNSP9fycvYNYQ7mPBNrvy8wDAXGpwq0ufjz65ViTHNvsamt4mfFSvpZrHnBuh4h
RF9rplf8eTa8HBfYA2BcwWz0HCYPsXkLD55hfeVB8oBeHhuuxr0MErQARsutS3HOtWeMqZmi6QHZ
Ui+GrhZq7Ah6RrGZA2Jm1kWzUBsRpcQiCm2fEIDcPvEXIMk/RPveVg0Cg3NxLPsE5FNHoer4c4eq
qdFKNHiwoCPt3NxvKnkm1w9Yi63dbp7BFSNVkEf+nNTxsRNeODFokd020r9msPFykUHAKJFYyRHG
Do4MZBtPdbXBQ62HeliooBT9L8IpdsvTEmrP8ZGAkkXvm9m7xR4bvJHWU+kQaKtzmm9cEaJjUzKm
a075v306fjzewMVao5BIKfm0mjhpVo4yTR5C5lYrW6ri5ovqCsqT0O2Pon+UGnpKjXqKDioMLVQa
0zzwFtNNC78Ux/9ddlzji78F/QyKHTeo7gwlnbXqC+KrDQI2pK0vIIMBx57Ys8pdwMbba4aAWBxd
npdWUupBWA9iSZyydM+4TtQQFgm8D2znCP1yrYLW1OAgQwW3fVvk3WUdpC6bRh5t8drsTtmagqH9
Bw7QfYGgSzvWUgpsK+sHXOsTm/oeDmaw2ggbp/tuyOxWgOCC3qD9GCnaSY+f4u+Gg3dSSJvK9oEQ
ZSNxw/dzg+QIJzYNVkxARAp95eYlvONn5yeUOsjdWXUFFF90nrWlpo15UYstj1BYWxRl4K63yrM0
XqveUxUusl6IwEGx0LaT+N+uEmvpwUbjQ2a6Hr/Iq6SuhGugPXor6AVWpxscoo1J7DSl2WU7Bl1g
1KWJv+qWV+1o4u81QxggDHgHstHblJVswlDUEYszfBuYZUE/Z9Y+nfNLS+igeSookmm6TKn/hYr4
cTYjOWaQDo3oEfvTlGxchV7M/yLG677TgP7PCUQQpwMHgMSU5Bu94CnNpLAC+5mQw6rzRyU7iy5g
aFAkkwq0BV7Fwx4u/659FBU/7xzQI21sS4guiBCqQctFYktJZ48A08TwuIKWy4RQbfDsa/Ze/+0d
JQMYhH1rEEtPCfii8BVyFGStUaf7KZ6P9IWCV2ZBaJ+fTKYgWBBnbsRcAOvPMG5LSjRIdw/PMlc0
8XDJeuaHY4QfZrntAkI6UOfdCIN1CdEDpp+GcXV//DtaF+JO1RzrA2mvS2HeX2F5TivUSKEGehG5
TW5DViSxfjzanGZTHVZFF5JqE8qC3rdLYSKDwXN2knrh1p8heUlsLS6lDroU5XJoJJ/fRev1sQwd
jngBvbxpG0aLkrlsDCsilq+wrnseAg/2i9SMDN4hWTCquBBYOZeSJ5DmxQFL6HeTmQxObGdL4NA8
J8maLR8dxXMaNNSxrIIzYOBCfUSlJIlBAnN01d/3ut7VHrUeBmB/Pwd9FC7HBG2JdQRAgtoMXDje
4mxg4s6HjExw8F8bflXAR7qioUG8kjmNtcQ3+lV+ygbjeO/B7i/fUwYTKrepk0kd3wr11zfAwIyb
dpRMcw/w6iEmJ2nc77dz0uqWqgFvoXU+uKI2z2oYmYb07cZd9idg4EXQuWJIcaokIbVl3rurR6/m
0BpjF5oHdL9CtNrrNCfUGFz9x2DZiAkvJ34aH32jIIyrGGBa7C9WSM+At4LuzZfgrjjtIH+8POnm
CinW3Sr/MWlLKBtWMZGCMawPUAuF1SA0N+OBQq0pXMgZ/gXTfEimztRMlDSXZotnvIcyFjUKh4T6
jonZVX0yaK/3wOAwSstGPhj7dwPGMsEdJYODz/IfqnxoQZmDQFYkqq5UiPZC1qrTgERJUHIoBqzs
EylHicIT0Ri2Qfs965cPFHZ/fsz/6Y4w+tpwgRqf0VRTZuziVBUc66Qzmj+rIcoadAihfu1MH1M4
6HCD4Whzto1UD0bcBrR4GwxBs2wzdnU1SPnn+k30wTJN98NjGE8VBLeJTKJ/W/SJC6au72uMbuoo
gL/YOzKUftCq8n/6kvNV1r4DojR1TFFnncK8rltiKW9TQ35gYjr7ABmloHrdA5D9i0suFXdwCEc/
1Llixyd7uuQ0Db+jsjo664rhFE+n6sOnKb3+s69Tdait2VkSRBnL9WL8Z0fsnPZ83t4ZF3+8yMfl
ONBD6MayDdosVggunfbz0Qxy8XGk/CzsaIIWTg+162ciH6B2wv/hSXVmF08+5j2ozwkurnWdNPem
DW7zD3LM8ePjyCw+DZjDKzKloakamsKx894JTZwgkSzdyt0R2SkF/Q4f4CIXjpVBuwKJMc9b5RGZ
e+jKVQabspUcwOgFT81OukAdYLOpbxBxji4BdoGW2O+05RAB4kp3I9ANgJAJiJxcxHYmjlD0ERtY
HdSRkNMQEleN1Uwhrz43Jkr3LFva9WqqyqVrLOlx1v/OColb5Bj2Iqj3wJ7iSEemXv24t/BeVeoy
DTs0dP2dnj7AA3Og5iLfBgMWxsgZcA4lsT/oiDeWLcvfiXbogk19ib96Nk29oDIsIAENseQc2IJ0
Vzn6MdfJ5Uk7+DqLMI1Y6cNKLYTEmVUtlIzjExSv1jhDTU3BeR0rVANQJxq7zzAXU+T4zZ8pf0yi
p5bsxsmAxuKhDXDqshvQva3eDe1rlkY7R8+qfoTkNNskpHeGHs521EjLy8YVw2q2biPw/nA/Ek0g
DpMFdbZHU6Bt+Sp7y40S+lJQxQr9/PoT2DpgPSeGdvbqsj/v10wjzxtiZgCKqcUHGGL3AZ1qkJzp
r4wKcpqrrSFRzrvdNfBjO74ENVyyJoQIjfj/ehb43BTes9pG9hCp8ltA+OCyVbKSUA0ecSBD38/W
GIdMX5agpiArig0QXYXC3z5glHsSfx+34yh3B1wz/HyxxOSG7Hm5sSNSH0BBuFpa9LH4NzrCGksQ
aNBWMm4SC0IMdozB47DK5H1wF6RDk521ffmVQK4bB3cl6/zMxUKyFXJ006iMhQRfB8RCITF+050p
L3HVesGrW78UmKxHo2LsJOl8kMAsqSlLa44ni0WEONpw+vpOiL+7UErzb0wfUoJVVidNXbo4JpWT
G8LWYmWWmKRnu26sZr5Lgp5N8pMHSZh0E8mFxa9k70k6mD1KtfJyJxr+aOZQNMxGBfplfFz1hIfq
JyLz7bJ3U99xuBy70s2SyHauvuerliQEbBri7ZdOhIwEU1xdvwl3axwligRdTNOcwLp8Mwf7HIS1
dFw+5V1jxpvh9VgYFDzo/0gUpsDGYaMgC1nhm5lW3SIfL1HBtwbCbejevYYPIzSWFqKJ0XT4iUqN
awDHF++lrspCuOFMad3O7tX+/cux/4jnIejHVFfQfbfT40MpYOlNH+BHBXU0q++Tj29FR2zd++A1
L5/SF84e30tAlyCyXnNwvDdEB8PHltQGuqmRb0N0xHRn0As5g2iYOO6Zgy5nwukxW7TU8pTYMWKG
vhyXCoa/nKoP5jOdqzTwbssvyvEGy0ihw7w8eLpKm9aHPomUnHrGsdmVlaHlOdU45wYcqshYOpG/
scN5VBHn4Kht/NhfRTSz1+naro9GyQuGXBmVab8X5YHHLWMr+nX1qzMJJekksCpnEMrOioAXTmXM
lMEsmH3hVmFyl6Xa5CTlsOuGsIs4mOjYhOd4/tP4HrDpobmnvw2LErp8XMD4HsGwjqVFd86vao3U
qXDuyhozKimoVIQYtsKANsiox1QU0iTssCt1Y4uGURUeMhRcHCOFxLQIuvjQTp3223jP0dI9+bKS
OCsh3UBDjq9GltCGq/QDsih809iY0D0UGh+IpbbdQdUUeJcjjCplhhbzeLtK8I/xz4cWanDF5u5Q
TKoHXS6VEMc1sbNa1TckSn8TmNaFpon9HwBWa2fkPrlqmYhA4Dv7C9gikbZxNy/QF5sva6v4KpPz
XAzKwYpCgRsErsJSxArH/jvt/s9Cf5qMu5NPC0GeO9YPDSHf6Nh3GG+Lb4SZiHvHPjP1fhEWikvS
No7pglpm3x4jd7IFCp51AVdCQ5rYseWMtLUtBHUXgoyQ6yOVUTRBQ9ES+iPmlHiKGZsoMNSmG1O5
XS3CFHoxd1m1iduB20fF3t5RFDViFI8r5hlvCKgg3Uq+yptYDRx0W+1TYdMXIWfJh/wp/U3bu6wC
USCWO2KLGifmiMERFIbmx+dGM9C4d4Qgm2l7T9wKSdAKa7OeQdy4auWsx5Ytt1msDtVwftj++s23
x/a5lpw2NkfktczFdZon8cMXCAw/YjjZTyhkmrmOO57qskeS9WU+dDue1p5Sfml1a77gSKRyg/Oc
RBKSHxCwOIZ3eYQZIIpk19SI6OqIwUKjSMDAKdZSCZdA4Jk9bQMWRf9mHt3Cegp90qqbpuaQBRXh
XCQnXntL7sIVqXhsXF69o49FE/kGkkbhKPb0Scp8jCOfEEVctInoUhkwtY1Bg+h51lmpZy2UaCVK
o70upuSQFDG7U2vUC07NEVmoAl2PKVleVaA6lrzhcWAr/IJm7msHWMQSEQAUmohaXSZEotiZS4Bd
KV6bYx/vDo9yr8T1aslTrvlrXKf8GPl5p9LdpbnuF3lN5lcEVD03V4Lh4VjKSmqOWbOZMcYMU1k7
YVjwGhz+rATj7702OAI0+hr7qlavi3fD++6H1eoPiSgZ9Cghk1047AAT/mO0xjt9YX+DuweSBYeE
liVVS8ScTGT2ci+lhrCFQrYXc1l0QC13cxpv3VGPQKLzcVzZjp2TmshteYx+Fnul+xMjDpUgL/gr
ZtW4Yu5nXY+fcKhALJLkFFl1BsYLxpOl61AdZPRBx57BWmdNCZ2EC11xBscDOVja4ooiIzQXlyVN
FKVOfiXqiviTASM1UA+PpHT1thNOWDDsA8X+2EEfAkHEROr+qSv6RZnCSaHTzT1GRK/vPmYfYAPb
hRVqV8Gz6NsoC96z6tUJnsvaz3p1Zkp+wiZyKn660ZEvUfqgjva90nIy43uY+S7hJdEHtywh9XnV
NmKw5AbCS1EpvMIblAMtGGACpRt43jIuM6/UwGmaSnNqE5tYZGbHrj+aAWRMm8icUwcz2nOCQszr
tg2aF81s1auAUC676bWrT/yBFmJfIplDquW/yw7f7ad3KYhjAVD+wzFgPosJRjGIjpaf0yT1PwSl
bzADT1Uap7lBuMXBcx0/+ZWd/GWjXGC247lo7kAVnMFx3YowWf1wafzALJPgTFftEPAzUUKnzfEb
hQIHIcfJNxsOxiZqwhI+kkaVmBmgdgsycrwsyYGjBwhL0DY0L77cTAJ0FY5KSO0hgN6jr9eRGDp0
APy5Gc4xUSQOAFtHDro3dpI8bLeaj/ar9mSrGvNwv59dJrdRSqhTKeTsJBsUM6v2wOZybBo3tXzl
cTFmq9+dhRyEcgoMRaz8khPSSrdznUULz5pConCiznGpqtQnN+o06SIwkejfxU9AAPzWe9jGA2so
2pHn6ReRPowoGu6ZIdqw4MhYS/14tmFzhTKSJlfDPNyNz6PVLI7v0Lhps55NIERz0catmxKF7jZp
SM9/uUF1JTv88To5Z1596TWGnetMEwJD+MZmGIOWcrI6NaVm0rmF0SOeSwkyb/JnLf2/Xw9jhRMN
hZ2uaYnREUKePtiNGQbwxpX4AUi64aNmqZeaUYAvb8oaHl2Zv8E2Zo+88Fo4oOs4HWz4RxmO7lvl
83Uxzw/toMe/8c2wvJgmyhDL902sflQJf8AyOYEUWHgY+k+aHW6eVs/Q35/huLhxX+2xhwCLA8fq
MBefD1LyBz+ndkbti7avtgnymXbGuk24bufT9LdK19or7s/kY9DbJKFu3r9vbUaGbGnrTL4iYMsQ
1N6fscxY0Rux6WSXY8XeCf8FfFFyhf3NC8ZdYOyLMCwXZOdWatfglRJqGt7J8MqZa0kJDqVlRPWC
bREs6P5pT3A657xzyGMzoD+juAAg5RCqedp5EKiFq5U7ojnO0lX/xGfy6rCGwf+ic1+mWARttRAB
+uvWBqHyL60eX7QA37drPH65KtPrwMClOkk70EcZ02UOO2aJ+79czTpmBwZleOoe79OiM6qJMdpt
qdxAP1Lw0bDo3KK+7x8SU6CH8FM8Omw154Rcr08i45x9dXAMKVj6LAlfCdfxCGZdJ44+GPwTmKn5
YWQRhRaF1VmHyz4XyLZdQXzHzSWDHZJ9sjenNNKlkTDihITCq6GPRb0YSpP2KwdFfEOs77fiZenh
4KGIiyamtYCA4leK11pBv8ImxeuLt61e+oZggx5HmoHUkdO5VrB7VfFVh9vnbA0m9LTdM3MVKfgq
OOpMN0gc374gZ+6TjDZmGofNWtPMKIVG/+5/rFhXRQYDEU7Tplx1C9sg0kLB8ZhEVHYVfVe1AKI8
XvY4Qfs3Lh+li1lBLnIWzRraE9RcYoRBAfKZggXlHHLmcR6RM9KzH+/sXAkSW6XsBKjJ04tPEje3
g4lsFGDPDDeo5vGS7erx/cnrDQQqCBsMTdjm30enEjBmjBMODb3ahYtWY9p+upvSadJTcqBCdjH1
sxmpljkcBOU14Zc8uaOauhKq6wOZgUy6rCd2wlwIbI3aq/yvK6eg/TRCBYVuZduicK1miXuVdP6X
yH19cMWYwYF9CjxjS8DogfO9WR029FJaG2JtkObOHghIWHbuY/rK4gKZD2TtEEhJj+b2IqUj0TUF
w+xg56pg15gdwntWaLaguTf1a+JwMAz20SWgdjnlxnyGdGZCC5nDQhLdubiJSzNlTqbV2jeMiN6B
bDFC8NVpbNG6EtQBoWENjIq2bFvdOZDpr6D2X+KSbTjz6HoJLIKQ7l8BoJTqo1R9AwZcxxxVPb2M
R+LfSDU1Sh1T04PEWnjbSMaa5y2G/5MMCzNuGWWAjJuMKK9Rlr1sTonnPvhia8MVBuUa1Gmx2rSy
VGmwyAatgLTcAGUZiyadqazuG10gkpwxcETnQ7ic9VLBG+smbxZ1SQLirQAJL6/T5Z1nfhGbXB82
g8ftv7SgHENFD1wnEyZw1EBakWXbQavb+E97kcOQ/JOppxvj3wQdma+BL8yj4yOSHQseXsHTi4se
+WG/RBprBzXuaR2FxMifuXRd9r4w90CKtedUdTlRYGAkdMjYVreevqRIDQhtIgj1jQZNr8I4yGtX
EwJfVwDCrZraQM/UWUMWjh6ujPHZWCDn/LsVDCbvfJBFo1HzWsvRrq8OlZ+tLtTs94n10yEpLDDg
jHCyp00ljxiZFjce6qI4eKR2mOQvOPcV+9P9M76TAWH0tM1fFVmh8/aQJF23ZhD7108lUXGacdgF
loGOq0LBlwYpMtQE7w4K8VflfDZUF94TwIO33NOVMsLu3eXwqAwNZ67Sl35XOv3ie7xphV0VTC0k
bUQ4cFM1APlx8AFAsNnHW0od+2kD9CpQFAQQ0ukiZqXZLCYRWfAtJ7yBRKXI/49FrN9Z8oihw1v9
YlWWtOoHwvQ9hhdKtTi5Wt/xbOxmMPBP4IF88VRMbmcFhO+lW9psZoXX23lFP8RqCDwjG7DcfKRp
IOjjvZE02v/4Q90mvdy09A9eiQChXweX8mjPecYZjhq5q5NNQTdNRbSiYVmCPczjnXsT8q7bDOX4
FjtpX+zqqmYnjllPNLThD6a4WpOVZjxUUURPkKbEaz6/N38XhXbEQlUITcAbj6W/sVaJJVWyTavI
muMKCRXsZlbj73geryVPXD6kuCo4RNRvfYU9fIXGOmVsnS09Zrec5nO8iGdtfsWRgDc/DF+xTBnh
Lryl0gCXgwrwFRgEh0Qy7O523YQCAtS1cjDI62Bwsyys9+WwL+0UuIGPl+XtSCDRNe5AAwWRZOYb
Hw8wtuQ5SqWvzsbLuRWB3E1bhF0k5LOg/uyMET9idprBqvmS4gkVJDCnU074/nxjNPUUkqNBuJa+
MjwOyiS1oyGO6XHIz9m/nePsNmxWPwGhRbZbl4ZcOB941spKjy04dszo7V1DN+qDe+mujs3I0tHh
Ek3QR2jDPKqtbRsmYhWrHrFWVBwIntWuMN7LWzvyRLf5jjolEXQo3G+JJcnwJU3RdZyQYu4x20pC
5TDBxogC3wKgZh5n5qUIm7GkyEGnxyIs5IvLO2xUj+2k2J90KepS8y9VVOENjUWnmHFfh5KDQzUQ
tSg7Ft8PiAku0C1m9ZzldH0C8ODQUrDxRC9lF94IpNZKAKAM/KidUlBW2o6fsvWlK0gs423EcUyK
VZIs6H2HnuKicsqoeHfIW/3Ze1jNu4EwQ9uuBfY2Vqgpn48/0g+u5ktkFOBwQGPkNyNeU8kXYlbM
zVhLt0nM589A4cSwbC2KBqXUfPW00KLi8ULRqvjiRXwLdg0eARiuW8vFQv5aSfjU+Fiboifaeor9
fWmhB6xKIosK9GwrfVd2DGx7GZLpsZEAbFhiEAkAM153qM+LVT1dyC38EfUdvsGZ13e3Z8STBZV8
7T1bPtMY3pf5KMlR5Oije0emttwhzplSbCoLZPcrcVPQrt6rOeefYpS6sqTFZnlZoT3Zf4axS/HC
iKwjXXz/5RvHGmePmw8RvXOY/Pn1F0CDv8bKQbJb95hg/O/NZTQW7TcI9E+Q6K4JIyHpN5jgoIcV
WfwqH4XPtgvPumA4xPdhOykNZHbUkFlS+Tek11XtJi5khMYdi9pjIqTssXOwDRUKTIWJ/L4VwIFp
urU2LCl3lxlv3EA7vFcgWdKowzBR1zfk6G/kM70KOWU+WJZkB4iPPS7Qm3myD6T+iMECEbzcKfq5
FCV5zJtDvq1/d11ne5DpgtRsSWvJk2Bn6K+jtIoF5z/d5/vFBPE4TKdUseZELe+8eQDHGnxcirU1
Oq0+omL6hhrHQaRv0Yl5gJY08Vrm8YFu9jpZHeHlU0oepFHKRjCtXrcpbRwrUqftP5DPKRtoiY4K
3JsSep12+6jbyQHqEKWB3IRoo77MFPJI06lck7VbvXkFjMBltIWQMAJ4qmexSVHg/PpO+dTAOerq
6OkMVFpvoW5yc5Sc6z8EiVXuQBS9w66TRoW2Bznahe/Xk9546/EtBwe54FS7iZxALVhbFciN5koO
V2MkFPrqOMQI3MEDOVMcfEEptDHVVV/NBiKDHYoOw2w4WChV7WMhN0rsVLEYOsH+Aj4ZSMzxTFs+
q3MCnWE9cmqisr4RglJxChnoCYiLD2nxvK9FBtgLBUe9P/uGuVEeago0KCTRm6LdzwoFg00Dopr0
A11bzB987Sbf0yOgZZKzsYOJcpSeroKYZZJAPVOaCNOw6gmtv9irZfumkDaeF3EltVAHmMOxju9o
PKd3C+c53e0tFtkqn3gyr0OZMBV6P+Ni3Oo0zjZ18vtvxWkUGOq63qGHBkAKHXY48ee4UWWZ+M0O
eRa1JjnoWZiMsOxF5K4NGrAd7DVI5OAEQ/TdouOFARn+Fukd40Wc2i4DspvToot3inp8lWsxUvjM
Pb9QqquPAhsot14tI4moyWBxITWKZMYhbMRaw8IcOZ6WCBQVnRPE3CR+w591UbC/k+n3n+5AdD7+
Zl6js0jnK9KcCh872nPL5StmcGPGigJjv0XKkquNObVdDK7YWglAAwNzOd9s3X7ID2lNI2kaVe45
tpOsH9bns72IaTEn+m5j2IOInUg6SWs3uA4wFrCwwd5jhuX5RfF0Y2mUnGVa/uP6MnFBN+aMbsU5
BM9bQemUEwp3jLDNEtNj33pRv72fM0ULbF3p2ffjxoUilqDp9lfmI/2e37hpTQTtNnlhD3js6m7j
t9qAkQhoUwoR6M163hdixL/7kN6ThlqRCuqELL6Sc/AqrBbmPlRCOaqzc1hsTN5J1KYrDm2TKLxg
4CBYFNWCyPoUv9/qpF45Gagrkg7VHLAQDoewbmYhg1gbGRq3WYJf01ITNErNLnpW+PJv/hnqJKFO
8L9lTHjfoBYzrDzIIwoVy6/msFqzkz/AW+OnY39d0RXodXfmFS3dN4jRa8ESkpoQSmXVPWnJtHq8
MCGZ6zIAXSVYqbPT0SHJJ26/3IhZIs5hzpLSsfgZH6w+Y1kbnex9qVYuhX8pgb8ysDWomvYlfYCA
eGwBJfSFQyEfHzFKFT/SgugzxRBSsYr+pgSY6BoFWTNJTGiozU8+0OLjdHi60CnK3c2+oG+cc11L
K3AtaMhD3Z9dlClB8arixTUP/jnTz3YmgEi1lwtvzHyS7JNVn51eMLFrl59zEGaX0geOZ3Zcwn0R
c/pfP02e7WgAxwuuT/xVfE7dPNbgS4vKVL1cI/uZZpuoIYWujfdDEkLctvifEAfg3vTwgUjsDtjx
PuyQGpfbOL0yPuQizuLGDJ3IMW/1TwInM+cbpnQnfTRULzHrv2lh/gRx0+ei9e/pp7h7GBGyaarq
wSgC3GOlr8g3e9RAnIu5B4VAljH6ZxdtZsjXGhMzLQkLuyYZvxdyV2xQnouUtCKOa4MzfEtwBLZH
BHTMJX9a48MRZLL9P5jSQXphywUbklCmrwfVJul54CXvkPi3zZ7l4wrSQCWxHbgJpVjOanRok8ss
CIul+SObNnsnCTXJ5sM+nD58eKQtTm5KM/JObnkNBu8uqnNfRMZO6RIv3W+qNeRUZ1n2+AmCFvNg
0NgcYW6P6rHOthsxwdo4OCQDI5Ar1mOW8Oqvyjjd366Z69qjPiNk6FrIezA9bp3U87+efvVsvM2p
IZAmuK/m9lyMCR+qX+ox/43tZeNsWpOc/d1i67YEtap93L9fHhJHGpSL0OJuEW3lvoirXVp+RRSi
HO/S2TgUlKx4zdYlDJsP//OAk/Fg4JiW0D8M2aZU7u40wE3fXykl1Hj/j/33CqOLHrun7wYjwuRR
SZ8Zdp9I/DDYHP2yaSzU4E3cpYLBwckzw+DNvHEkq88A3vUSLnvXWqblqZp+ppRUtuKD1Yh3bj2f
o6ih0eu4exb6x8q2z8oKuvk1QBO/4fMZ3StTm2mli55IVjCS9+xWENHCWA6ymz/8cbf58xLHNdGt
RE5LslTdjH3thmO8PdJ1qbwlmGkOcgpReTzIF+xkHpseYfew3VcxROCSju88cQgY+VjtdL5+ZHzp
vG30+r562uIRO9xUbKe+pUdSfhHmPPD7l3zjTWYzVjHrM2Ja4sR+z1GQiDjY20gjKvyXg2EJh5+t
zn4/3wOabs2YzqhwA6Bwr6eEEVkEi8TM3V9Ff5hkrAD9/cVUstxV0no+GMPEHBh9zsprkwZWf8AL
AQsPLedAOLucu1+pJNuzqxtVG94+IRTc48XEVotZv+Fb9rB8wsOB//z0kdpBBejjNam/pxlO86EQ
UTvwdqL28XWdnDTesWaVIBBBteiDbcjoDeaqncdxhIqdyhSf5jyWl3inC0lGjA/iv+ATvQEemULs
TdjD0p5m+OdfvDGnIV2IHI2dy4/X+F9x0S92lR4j9DhMOVzO9/3Ep/vqrEMhxtbwApD5S84Yw2CG
1eyGeMYFH4mKP998HM8QgiCdmVvb+bGIgMmS41oNaF380zzczr9akxXN+hOxf7zqFU0mNQY1dInM
/vYUE7Yk2Evyb6e5P5i2AuCz13QHhjagmeHI2hFa/FSYVf/RqxGYIWFfR7uQSRVEeSGdAHshneGF
f+DZwTLt1T5zDXqAfjxsUD6HTOrI6rVsbw9iwuJMhLyHEN6g98db4RqR3BB9Fo36LGKlkMa9tm/g
FH+1xs6q7S49UYbEXNLVLXTrXtoFHS9sh13QzsWJCbkLYQIxhACHj8vRmcZKgtcAlw+A/3hbUO/4
UmU78AakvYmqJHVJp0Wrx4S0bfO/GaSTMpdsq3BZJulTFCLQ8c66InC/yTWLHgZSVsUmjqxwpo2h
nWHf4aABxwKQKxDsF/xIfwwEGtm1bFo4li0BLjH//4R+cEhjTf0G8Vno1vb2aozwmeRUsUtrAUpM
YAVv03RJW748FcSKwcnzZfuqLiBrQuEbqEtT/XdrB+iFdhpCXYLdeMWyT+SC+BrB5/ft5K14UDJz
7Sn4Tintla2yaO10K0Vjj8qNBiwHOBs7joKypgckC+8u42yVQ6poyIaI0S+x1uJr7gDnawMUG6DR
RppcdcHiNfbOo+sCgO8/sGZeTDgMxf7uZzwJBBbhbTAnkl58/wHHvcKCJgCj7Wg5rzxbXzpBpwbs
XihlXAaf4DvQeKjWzTk9TPULVBNjNCDhEwoGKYcyNavFIaujNw2y6WK1Rg+hxmaZ7kPFXrDISEfK
dJId5bnQaNJcICG5x9S+DZYEWFxjjtjsUr9tFnWqJTVPYLT0/6ZmidCc0c/C6ba/BI+hgQQj83rI
K7v6ZZEFaaInc5kVHFiOsaeSSF6JoA8evArN9A65XfRu3h76IClZlqvCEB/NA7J8me5LAWy/AVf+
1m8ylIYFPBqrAQIbq3K/hJ0lGys9g4qCcLZOERfAALdF2CgdhZhfStBTxvPWWuCsxfFTAkI69zyk
4GU5aSiq6BDDU6oTAmxH7EkcbgcwdDKKQ8KohVL944rOFRrRHD/unLjVoa92kYoo40i9C7Et1dvX
KjCOrnLkKSa3+9j047bmoRGLGIJvFQZGBc1iPl3Y1gjbY0A0YPFFvlUJYwsj09VToBJcUqocKgw+
Hj2M61QpRb5JJHbcfHKqhpRx2CZZxTBgzMSgU75+amg1NJYm5B15JFECURwzEOMwRovo05rqgus7
n3URob+Zo0AXw4pz9RRy690+h83vFmMBqT4yIIsUJFkMqMbz/0r0PBkCC7F2qJsQH0pwPbhEIjnq
FRC8WCA4uYaP5jqzrzaCxcEXgK9KjEFk647cWToxnQCksgrXDnopvsjltm9vGvWUQoaUPDXwbgOn
okXQyQSoV8eT/SdBu4UY+Xdh6JPQMGCyoQyHAzHSYJrSwGPjGnNmzVFyASBAsLq+aZegIpDfCnnJ
jr/rAA5eecJaGOJJbEyrfn97w8UhvqSltFJuF7hAh3hZABVQQlVdAFbi2+1XkvOr7o99PmwqHKwn
C4W+m8f/XeKLTqN/O4Gf4JEJWVQamDsdvhwfauLZ8WhXq0f7AVGIDVdVSQckk6QPFOoppX+oGX1V
caL0E97+Du0nypvZVmPBl9E0XOgbDd6JI1RogTiXWuy0xiPeLoAlimEkbZU8/0LluOKT2HqFPIKL
7kSCr+mMGlh3lMrMZ3+o+3tYqgRdYLpRtc2eiFNfXWp6HrXgpG5HATwKg1bAHXgSFIECl96chr3p
GAdi46C26lX6Y7bld8d30sQQSA8LkTIz1MeHIqA+ljJn9eypluaCvDg5oFRPLZUbuO2QugOR/uiT
Dyi12g3r/plBAQY/wHqyv2dzfJ7tyOuMvxqy+/w/vMVfwX59cyHTYPVLVS6Hsa+0XSSaaHKQRcFp
cT24xyBTpqzJu01VwOgWVpeWbM4R5B7w+PPbwXCKhY08Czq2eFuOv3JIYrawzjR0XuBa5Rh2zLzC
w8Sm38yaKkOyPdNrW1xnSdz9Nb+pXyJ/7jo3g4Dw1r6N0/AMazxSzh3o69GLXnpgDiDe6sQ+v1BZ
3zSJ3ds9vdqeqYvIDjaIcSyGnZSfOcL1mm470tBtn14AUXLADe/7bTAv6BXAZntuWZNloUUV4gcE
M8TTIse0AqDQkk+laciJp/0m4BVcAjzUw4D/s/PCkmrA85kp2bB2DY2tqtmBM4e2F7MM6GkxvQuy
0byfrFD1uJDSN4W6g5jDdl93JSVBrkE3gQn/9DZ9jZHA8x3AH9lPFId8fiehT+7gVyBeSar3gWRC
usJSptC9wNQQ0g1ehNuRucjZJqISU86LSGZlkkqydF0sV6xHFGSJw9sYD+pu895UaU/R1CbxeEsd
C3fmv+j+qNjeZVAXAHnnqHyYSBu4h+9zahuQ+OLi4i+pcMN9doUOdsDfPoKeyU3Dulc6A6Wcvi0q
3Cj4ZRElrig88qGL3WgJoHMB2BuAXgqpOMTIzePQsKZz7RDe+gAnlCDwaupq+xr0SJEzG6YtFG+H
Oxzgv2HEjfbIi0358kSMVVW9BlEwJClfGRPlALq63fDc7V80K7hbHE3c4D0+nZ844gTRxiSrj5zL
tTUYL9bpbCSr+OiEkxk9yNcsey7DTZXwAOJbHOD63awAkA1Afi73q4f6Hf/459zYAC964no6XC6H
e8O/XaqMUffgWk5OITZVsKEYJSeMUJF1fb2vkrjlg97G5xSFPAasPcmBHEcdPcvt1QWpy/KCpDiq
eKqgjJ3vKQzjpOvn8HHt7MxZ2ztEN9nDJd2zq5qqkUrIZzox7x3BjBIfawhIk+6LXcyLarhjVJDv
qnpVazVFmEHgdQIdEoWGSkxShpmTWwaqgfPmxDaBbCUK238x04FAkg3exvHHyFXQoNnOPS3sCZ8A
hxNJMRAOklED0SBgdvxX9Ud4K8PcfJKsnyDzaxOUOJ/HG/F//jQ1lehaPC7/QUqOHyT+07LJ4wXS
JH2K/Mf13nXHOtN28z59cjfu1oznnaDipoG1ufyoS9YAP/AZSFH5abSYN6W0xrKKKP1MsIlAlnun
NDhpkdQ5jlsotutoxIn9wCp2ZjX00g/3lc5hTZ+iX0QqoKgbr/JRBrtklT1evnijW/OwW5r8senR
Z6Z8LiyeUUL+ml+JF3exnCTgckW0VXB1/vksXCv+YRUqb64zhm5PxIrAQ1VqlYy/3hgPj71Bp7/0
Jpn1hgfGnFKKlgW9WW+6/4ryfbFIdmJKCxsZ/HI5cB+HBXXY7eCPYqIopmKwWgIOyR2ZCdTNknRC
TO6ZVG0V2/w5HfGZkIaT8QlQcHxHxnDR6/xknJpqeTUl/FQGE6+7ariEvKrK5qoT349mJgfPwrKk
V9uPEe+KaKXlQ9OmiwIHBPJKj6rxJCB6Zxqq2iDMK3kbYSCM9VtcJUhc+kSYsqD4pXzZ5aLpVbiT
SDhU/8MTEYLdS8aCtZySi/257Q2NRoGxBOT8TyzCupFmHl/BzJ7vbDSeEPXp8mQiUFbRBB3ZjhPQ
PWL+htLKNKcSSkjY/SWSfFhx788FrcJt4axg+1VYb+6qhcZVNnWgA4G1IxGJK67NHC+HPXcv1xwW
mJSrcFguzjavcvj2naqY8I2Hxvoruue/lu30JrDdvd63fmq35auEpljlw2pECQV49prfbPaze+3w
TBrU3+OYT5yEfP5mmolL/zYewrWyl8ADNtnG3Vqml1/VYPcOERXg5RxUBnjT9PbVOfopMXv8OrLZ
ekow5Y/hcIBHVQ4EsRjErOx+htd235mAWuqitf5EDnj8Npja8OzxgKYsNNp4OK1A0DfgYI2TGPsE
N6KODVL7u2TAs9JtPM0u9SwCDf/8Ny7mog6izhL+RwTwMMaplFIwDoERHqBapYBa9XXaJP1ZnhoP
VFI40POrbbR/vlPRL6Xj4jBmcb7PcFQr7BPZslmLqvSwHCadQod2XjFndHO86yQ5fN1AAViBu5Uh
QMPgYOMiIpzRrBoKGUx05IjkTn41cyF9ooW3FVQkHU6jdZKXingoNZiEdbs/AfKlSNDCPLwWVDb5
4V9WV408N0C3idlYWF6ovIE6rZ3zN5AgEd5sh5e+PVQCyOaRk2av5qAoXP6RoB/FgiXrD1lVjkrH
65NP6YQBslqvLkOcnidHNqbK6adHTf/FbCQdUHBupfqZumFVqIgiOg0hvu51IP5cG3oRcOtM7IaA
fQyIoN6ad9WwB0eZX2YjikHLlnlzHqBnnlJh2eVpq2RkmeUgO8CVFoFj00/otTjoOdenZjLtKzbO
rMF334eZP3BZTsdpeOnuv0s5pdZGE8OInsvZXBlnsVEo1k9YdRv8V7ZKaBtb1f0LaP2RBXlCEix3
sls4WMTLjpHxZoC6SYn0hsur8HmfOnNIEZx/7QQX3dKVJ5hKQbZZy8K6aVXVnAQ20jbA+xpj10wA
SkE85E+cA+PDvxjpr4j7UFK7qnmEH1uBC5x3S+zI7fi8WRnOYVi0JcZGHijzbRlWvHHhPBgbY0Y1
C1AoAdFG7LxOrkmKJO+DS+lZ5lHQbwyn+WFcUp5emPNe/TmsYH8H4RgWlucYuBmg+xndAiA85glK
VKz47FDzBUasVTV2Hb9CFdgzMyJG9A4/SH3DzDGIsB9U53um1EsXo0TJD6N42inOhIo7lDwtfQAM
Y4iY3v7pKIHVIEH6bo9O6+J2VtH4fjbLclBJ7BQkrhNeKNPoAV/L0AP+3vL01SccJ4V0Tr8gwviZ
a4xXZYpxIAQ2vQaMrOco6KcTV5NP80T3ujgZhbGRIPLe7viik+f/VhMWF/3gi1tCd2rfU8BoV/W3
ZwJiV8CoFlLFvmHAZLMbJbifbeY39wp488ggvvDzInOnNPqvSA3oOOtzaO4kGM/FpqdXYoP1R/Nv
cx0yY2VNNc2wz2E5any9VwR6mgaE/JolHK1QR9R8pK8H4NfomxMgDXvKABVs3ljCKyLMJEu4kRyV
x/G1qzamv058cnWVwkLkrI5st63k8CNrBr36MY61GZwiknOrW8CtvJcuyeK7eCqvMNx1fnB8uQW5
44ENQB6KsWUkQylp2DxqDM2jFhbEUmnNtl9VZk6lqLgzlXqSg2K0CCZjAhkf8rk57M4xxxAdi9I1
5b6eFt8cK1cl1jKonn8EeU36AMqCpLchVvu+hTLUdj9Ws8OHC68vKun2Uimp6pdDNUTlzEiOpct5
ltyWYKy5I4i77yVvTFuBpGBYnmI8HxY05/lNTxhbIvHzcr+CWvCqFdeWJFbpnU4ovFG1jzNbVcVL
utEMN+mCeK96w4yLmaF1pQCoMLCugJLo7HfGN76J+AeRe01lXMvd4uHq0JXmFcgJYIw+GSfQzcMX
NGMd8ynlX61cjfrowh2tZJ1lEO+aAdxXfpCEDA91rimQ5P+UAP7gbxJ9wkB4s97BmdlxZFNgfnei
SFtc/EXbp5EzX9Zfg7Q0J2p9rLfRYMXVhBQIvhYp3k+RWdRfroPGK2x2Tgn0Cj7OwbybPeHWJ4WT
DWoD2MdMByC8iysL1QryVHXwfYv4OWPku9GABIL1QYJy6PAczqCudCNWbqFxlfeVTDqw0fnfJHwu
R1ZvXvBBt/cUKSpmXLo+De8EyPBD41nUQgRdc5/NlwR9VhDHzjRMO0CpIg2yTdflYcsI1jKS6rfQ
NOxrYB7FdsdDKYk81F240Z/HwcLLk6xGvspl+qN2/fwtX8LT31hTzDOK8m1x/fEI7xkHLhOkto9e
a2g9/FBvDx2zLP49k0fQmisFWJ1FKbAkwhvH9OjowhktoNjxuzTjSqWMQsNRceYQZ/avfo4VOe4t
f5f5HqNVoLiewTml15Q7K0CmGEn4mh7ssbN9Kg6tQHnSpmyGDHzCzZL8MiSHr9DaSCHrIofXzlvJ
2Da8LNhIrXKzQbTGiAGlQljA4yD0dmhQVy+/FuSirhvxaLm151uOzDOgAdBJTRSsFJGare8qVPgI
PRiCViY59+l88M35mPcdoychhIDpgtjSN9ba1FZjOtGbo7vSZ3qaWPohSkBQbfRGjmZgqeni6O4+
QEu+n52oADBzgl4PtkjbDyCiN7R3MhljkSjZ/7p1ZqVHi67qVnY7jU1KVs7Dl1rmUbvZ8wk/h1Bu
2gr3RDhzWOLCYRXX28xeWxYCeYnLXcreOyb5tqA6k53EtCjgPuA67/PeSOIjRxUkIBIIL9pR+d+s
KVwKDiknWG6AsRPMaU+AO54cSz7tkIMwD9cZng0lyae2NQpwFNVH+7wetsI4hUly3Yiaub+2eAfR
1epWRolu9JA5IbRIYCmvF71Kuoii3rcf6ie/hYHSbzlHVvDR6Y1kBzm/KO52/+vGn6vGEP0IhCzf
xVm9rkybdM53zF/o8lSMH3Slr7e8blNJK7/UzSpOxZ7LKTY7YtGDDyAlrqnTS94D008oMYCCHH1n
Atna5zYCWNNkBjQiTNlkeX6VjRKNrpIfKxY0W6CqOfRS6aTfKn8h0zwA0VNJuaB7MR1l8Idzf0QS
LNokfpLBhswomm+kKgsUGMdCXjvckZJrYe573UlD1+ZhIn0GjaDqjUkpJxvDK4ILx/GXgMZBBxYk
4m3pwuC60RhYjXjs6ihFWXVJzrI66tX0mZTtciTrXxJ1eQ/uehZuRF4sSxI76lk493ajv+paI7RV
Vd6HmUOdcZzBc/+adF+UwVNq8Fog6iNtKyMlLjE+Xq/u2EOtgnjfzyZvq6BKImrLRCc9R1h7KdcH
F87NqDFLXqvVad/vd4t02vjkKtBMYl8nDek4t540Yfq9bUev+bTAI4YOMweNti60Z5pUBAfLgwk7
UVhmPL2/EbRHFRUvx0t1T8LMFRGxgbmE4qKl1iQOGYud1pEjV6/qkPENxcd+EqyolT/X20ty+XJb
Z5GjX5uYwVtVEM6Api4sV6W1LmCGk6ZL2WpHwZ0bbycDaQzbHdGsiFzL1qSZMlaN0mvSLbjgJytN
fkyNuxQplNgOX3FZln67xI0fonQbsBKepLCpCz5rX64cmL8ePdVd/WMQPivgm6ZGdeCW17W9p9mo
/vAs19du4LHMQwuaZ2nJ7NXoWcB1FzE/4wq8S0hpU/jrnzQyTrFP0hVEf5Ej4XVtEjhqkdpOpoLI
pcHLuyeA9SyO2bpy5hKWrL4TYdDL8mXZzK3sZK3n4oIzG+dXyEeyIasyw/q9MJAFwxXu2pK8dlLd
UTVScqzCroorIMGvGTF9Fc0929zOPnSr+5bQtAmkQQO2JnbzcJLN6iLt1eL5EWowOvc29l4rJDQW
+u7mXNRnEkQDBW9A/1M0YGb3BInPb5CGw1/bahJ5qfvbFZNKPYor7a7mLth46dSbb50erCkUOv2V
9qeDG6NPOFDt656eFoO8m+Q/q72XKE2UIeEGiKOnqa7Y0Sw98SFWcEHzjUGTEiUvgjxWqMFwQv8C
Yr0hXkhpdvSjaIwwoAvqID1d19GVkbE/UvSDE4Nxo5z5+QknMSWV+lhy30f6dM6A+2QGtSUTP+wF
vzBQlEnLZDl/2iGatSPFJ51WUIhTcxBFulHuFqVs+zP/vFo5HGtqpYCNNXPFmnNZiTgha1dRlQq+
m9sXeREu4EzA9yiF/zt9WezDm8Hn015N2umBzwCzaqFhirf6rUp42XWU1w2zVY6J53xFi3MQeJ1s
MOjRALUSMv2imVVUF6D41KszXh543WbPkhPqtzmWvPzYkHf2OjbZZu61eP1Fa1raAPFA+Tdlp8d5
PpZvKSPPC3wcQv+sbF6hNdbbJJfdHQFHgeQhNQaYohMqv+PThZhwFzsmFrBl5/7LG8i4ENklAKFC
PdQX4su8wItwXQatElPjxTjGROmIS1OgvJd5f6lILPdA03DJpfGP+xfUAvcd1jY0S+0mByp3Jo6E
+rqbznByyhlOoajKhE6+E9LNr7xenxnC9L3gxtThoGaV8HQG5QCM+0/uIvSAfzuI9Fr4+hD1bv7o
MCQ+FJrLLPsUKvwbMmjWfUfJv4HYuUK5ctJw9/g4Amy6ATTUz/n4kWSi9tzStt4J0YOpw199jsfn
IO+zvJsYpOWyDvZSnpuie1UatYPKtFI8kHWIjdULErtu+QZZAnQqCeO/F5jJN+CD8pEH/WqZ35+Y
g07mNh7paDHGfYHcBYowd2K/83V8A76zGJXik+P/fY8z2D+NPBtvxMVNHiXeqB08j4rvaPgUJCJz
BKUuSEZ5A2flGS9kAFoScksTytPOPeyV3WPCl7jBDxsdeoiO9USwBFO7q0XNJ3oKXgziah/32VlJ
gxV28DOUvAjtpqivc4kJtVe9tx7fN4IGtqtxTcxw+y4UTEmrpePDB6UWU43HHwJnkmeNTRuG4ygD
OIrJX2leT5cvVEpSyyZdSwGKPBet+vkzP6kZYDG7veA4OKvCOvRJImLTn/LrQsTRWaqs7ajbRKSQ
ZMzl1db7WPUq2QSZPeYBjzii1F4dAem18Nzsc6sYljnm7KJnO+VdLm6xUoUIVIZKVLDsCKUHsTo5
dxlwyH+QbBAEcq3uWGV7sDNe4O/TgA/I31n7ex3lofzwpe8wEUfyXIjoOnNwlw0lvP3LDFqwq3Ed
Gict2r29EQiDwuPK0ltkSMjsWmN1X9uJ0CXKfIqPiG9J79mPgdCYv0XpJEUkjsPSclUEhbl6u9ti
aevg3aBK8IRA/WStmVv314gxm7Rt12lqHwPEJoBxZv3aZ4fxxiEb60RRN6FRrGUbGFSPZFGdIHJ5
TjgzZ6vtnK32s/Cm0RsbaIFHPN4NKFVb1D6PDSCw/5BswWGtiWp+RX/rFc2GP7f1KIStgTZBfaaO
1FiD4LeamuMuxE2vP4XggIQ4dc1GnuXXxR/6fbcNnuhRJot8xkg/uM2B5pjM6TYXvAPv7KR13s7D
iUl8xk7l+jkWa1zmQPEq6iXt6P7fj9m9beyFRcfPnlpueeEStMIAwGXrNiJerRsHxoK7/uGOQd8x
po6357yv3Wtw3leBxJJ3t9x1RK1CJE5KFQPd7Chm6qFY57Rmg14dNurhubN0Q2a/Zf7swDoB0ZF0
hYKLjQKv37dwftox6Px3idzMj0spqM8K3rzv3OE4sSlCnirVM6y0DiAoYfGkCwxRFDUFYBReZgBd
8Z0iob8NR8ZCSfL1TbIV3/p2QyzK0OzMdp93VqJL4BgCgNqMg56jCLb0LeJjWZv8K/ah7eMt838e
h9BR2qvqF3cGu03a00Imgz+X8AwidcHxN3+NQq89I844hzgPliYxqbN74fGSJCbBi2i2jt/rtn4S
cHX6DVTxaloN78uBmQYtB8z8gC1Wcf0RDMnX1ivwS/Yzas10uKa76YhrZBSvLQb04e/Knhn7PdHB
6CdAwd/K4lr9p1HqK3g/RP9h7C3PyQMJdrmVe8KyA7LOjQuq12IvkScdwg6nrPp1fG1n9gzvnHiq
HVKYfOyc05Nh8EXI53q+fNZ+jVcG+pyWcAB/AyXyxmQe4YOzNdKYWzsxGiViAkAEImoNra1EVDTM
p6KqNEtui3CibxKWIu5tOw1bmTzCUhfZ/t2cBUBsLMBLxP1wTnZd37gs5bgmHWcAUKXBS9cPEoar
9hKwPxvhOATasmZJVxyuTpF6ybT3tt80RBv8NZC4VnQrPxhLQWoFmD1BnqIxva8ilI7RW6aw10qE
1g2B8zMAAti7+lq4x2JObg3iFNpeArLAdd9nivQ1vQEEV5pUmor/jZqP10ZPq8x8e8Kg80kXbKXl
btQvTm9zlsluM69gl0mKjidZjatd35VnyAMBFg0Qrqg6Ub+RVRZ+N7SVbjHteANzN9iEjis3/7G4
xIYLm5fdxttoPVNwwbxBJ9uCtb6Fnh0mgYAnfMxCZ3MbIFKCVYX6+hdvxtXI84qP+FfzB7uPJzkX
e/Ku+P303lCiEu3N/GmdHTSRxbOwEOBdoGaBbWn1vvsZSzDM93/OSoqKMiiMWCy4zbh5yJjRCK1Q
1vizCcQd5gCBw7cm1YO1leDgpamhWGISvXb9iiPLr6Two1H+2YZQMI/vm9wgYk5OsaK35+fxvLk+
GT220aq0i/4zYFk/OiPGUVYqc4miXkPJGrL56nkw4MGaKsku0CAKmeuVRgZ8XumLONyfc+tAgrJy
ea99ku9URBp4rawSOENOBY6zg1QyEMH4kEDrYoqlgw27Q6JFSEC3QgK8pq7TYzOAQLa/kIxu7Q8/
uGOmPY8QQrSsDOsGLE1TjLZTP/JEUhpD6CW2Z/HPPlL3DtobH1i/MO5JGL9DB1mUPMEPd8cF4eut
xJBDSsY8J6NcAE9wRQ+LFMocLFILHT2UyTjWLSAMVyqlW1XujbVfEYZuLSR0c/B8FytDynMcEULW
j6LnHMim3a55yzcGe5P9fKQ2xMDnky12yuyp7u9QFr3ATwMPBnsZrIcpuPtmEkKXbfh7lko7Gwkz
AhJ2DobzAONFMwkA0BvBznf1lZbV6Eg+CMuvM4jcEGCS93vxP/+M83ZivkFNM7U7g0vlWm91FQVN
yMWuf7hnBbn6xBu7SUdmbGJbmEC8sKplKrNSz9xy6SxWwczguO3I6asLozTb1x6BnKD9cgFFIaXS
GD09fZuM8KEyGB/J9932PlgxskUG/9+1lUnyFaCmfrVTGKVYsXXYqqhngbunYTWVKEwaUuI4k1Rq
zN/64WALVWw9ESgYPIvGPfKBpNRBmEvMCVhZreXIJfmlpmi0GFBENfCi9gZpG0qVdj29yf9ryzsT
Jj9VSvWGHnYnDpdOQSjJA6HMatezAW/iPF1eo0BjkVrtbUvbCpwpsRJjYR0tmi5o5fdcM3bwC9ZQ
/88V8f58UnPjaJcC4qDTJdZNt9u8CLO6tnOR3VCqr0WPKdtQqbl4ilqEmiUg5F1b0sKZGDGRZxJj
ALF2XcIhzjZsPU0lqqtCRG3I1M7xHCyQpmfKKQvaK/WMJmj9wwJVOEwBD8fTZOpK6sH2DNubTsuZ
ExMkhhkq1sBhqScdDCvzhoD8qQkqtWOTiIzY1XevRR3PSSCaoWeOYTfErIqPn3l1c/qqNpZt2w2T
7m80cZ8WxLJYKLaKqyElbFcuQBQ0MPMcZGWKtbL3HZTHRSdNAFyUSU9FSTNemgfnX/B9sjKhvg/z
//DCr+tp3B9fx21D4IHDBIQfNvU17cnW9CZLpzZ3SdwGUC3AU4kyh9LcYdKPGHEGZJ0i7S1eKCVZ
M04hByaoIu7jLdbzs7ZKiHXjWDJ59mAzARr00P5oAkzpNoZqBH1jlX935GYO/1T5EtncMhvZJp3B
P62nAPUfr2I5+exwqZzUEL1ejyQhXoRF05SPSeLLaBCNrDVTmM4e76yYy5RwHEzD/IqBwgNbdJDZ
IL9YJFlBaXy8nbAvjWof7JpfwEmZi+xf31lTc5hT30Soukt5i+FMUSqE/pGf9RWlHbQ1b/6hRtzh
1xjLzD05SGyXLrhBB5TknQcSzg44JwzBSUVIt28erZI9X8Dx5Ra4j89SEVx2KZam/FAfqx6Xxsnp
nX4pt3IVazlSSiCeL4tQLlynfhbftU/g7ncBYFmoDjOvjt8bLaXkgROaB9AKM8GKYiN/kNQtDzZU
7ImUQO9Gkcu1Gi27CNhaeLS4+SA4RLK2oxuPSnjHT7/ajBxe3JXxYY6O8yvwGJcqaY6XsUs9/YHK
As0U3KnmLVPLuiRCCx4rET8CwzMaZZqNHdrz6O4nqRF9MFF2zd3Ux85fQ2tUrNGHQInqrm9vfOo9
/BtNXwz/TQgHm0uuWU7R4AYHc54/lTMxgNC6UnJ/ZmVsCFKskvkE2chf/+DPxSVR2+r3LsPQuDh8
Ts371tV16wtnPjRiJP6BVImsN6HITHN5K4GqtJF3Mp01t3xnndtvlnJbwGTyF9zzRtNaVbBMMkQU
wH9g4I/kGV37SzlH9pB6+WpkcdhL9CDLAXT//t5KFiTOxZHk3Gj9COSSBdamId3BPiAgu6lVT24g
QALU9Fm3s0WA/d5zrAwbVfVjAKh1eq3uNPJfIG4JyfKoMrtgHLXESFyqJmpgPRmRKmOHhMuq3Sdz
RvOHJoU6NDJLh0dKbddHd++zqyyxl0GMNOpn14OefvST1fD8IAFyQkuQDTRBLK2ySLOhNHL83kRP
d+RFQ7DnCkXH+LAfaUK3S9v13dMC2I9ESmGOtHxhX1XfWHkns/jwWGEr0diMbbQhk5zRM/KcSBQ6
heuzK+kvJ7Sp5TkRdwKc14LDeR1fY75udGhmHmHPBl7rc5upMt2P4xKDdNzAARtF1Uw60zEeCabr
L/Js8TyDG6L53d1QavJ20d+fsofpp0RyNlekcXvJh8oeGTvUUKSXb1PhG5vDmWZcQPSFzGevUTof
0DckPEhRXiMq39k2zW4QY579/xInlBUx/4t1gWUwD8/nQi3eSQSiySj8UpGbe7YPaGUEnVobhocn
S/HE9RpuKA7gc/+VP/afVu/bZ50HT+yfVsIkvzDP4aLthbTp3r5IDL2RuvNCAuo35ysIcpiZKA+I
IcPXBOVRXMVJSBeHSXdmkdlM5iFSCsivsrDxzL8x1p4UJz1qN6g+dgzJyetoytvOtjKukyP/bt45
u86jeIwQBKiMXMs5HIPjtY89YNIqI1vSeOkCVUg9uTb7I5YHaUd59JuUoHFqekX4BEhwhzo9n+3J
YKCmb4Zvv2ta/KfQ90mzFQ+eeqAgmSAEiR7AO0a9Ssq+VNYHIZrq41RuPivWWQuVxcgb0LjL69J2
WgqwKuC/M4Fhq8padlpG4v1/33hh4IDV13KOTZ8aWH/tLyKiF1PLkN6X/8eSI4skritpHZj3Gheu
9atkd56k1xc1hUqgREm1Su7PJSIw1TgtI6Q2J82ebIv+ig9Q0gsmCO+52KYS8zGENPJbb2IE6ajD
HlZwtVx9mYwKvHv5UYU8XI6920cNoSuuhd8SCMAa/Snl5Lf2ditIluBpibriPkm4uJxV5xvAGq73
nTftt9RMge6D5n5ZuwFK0cbB8nqI5e/V601qNn7hCtRH+a3wAMtwEYoLupcUPs/MmwktqXNMoLMc
cgo9jOeCeldNjeHZE9CDkEwxrFrjP0N7jWnbsg//DkzG0LRtd+pz6StH12d5VsCqLDKWJdHbhLNi
cpx+9gnT2fxTGutXuS8QUPKAFvbGPVWIZUA6spk22fR5ITEv5i1Yrj67XBbfP2l54+p52VyFQ4zw
M4Mzox8lzgfO69MQZkf6GfNveDKKY+WmX/c8IEuLOqk1vUEnZBsGRKK6iQ3+FJWhAfmw/Cg3nVV6
tOeIUJ+jkF6w98u6kqflyDMT98tVvTYY7zSyHlMeuCqfwQK1TAGhLd+b2TSa5IbazWdruQs8KMzc
dpRuU/V1cqD5/ZDLIVOG8KvQnPgbNShM7exo+LYteNWlLs3NN9ZlBV7noq9ql5/GG/fzA/KNLAU0
MdjonXVheukXRf6QmHyYF2gIcP5jkd64n4w2Gzwq7wLzt0wBorVrYeaHN5fWiV4uoQ0o0XPoROCp
8U6IY95zT6SJWaCZcdpvXCFSUUDriaovb2tcxtz7YQ6OkRqVxGC6uDO5DH7k6P3o3eK7hhj7bIQ0
eEoirvYEaQ3i1/UTnmyb/suSI/G+ZVI14CR6FvnOaz/QL/63spna4dWf97hql0EoDBvytVO0pnAW
Ejz31SNXZ+Jga+Rz4/KGYfY0zl27EtJt/lK/XNN6lWxp/jxX72an+4kd9h2Os+AUOJ+Dgi/eU9da
KciwqACkhVwV9BeQKSUrbwE//hcaEGQnVSft9uVAimixhg3QG68Ko08s0aAAsfKYyUIwtwCNoz92
+MVxFFJbSyCVpnbcH+FrXNfOOP8xnSC+Mj7RHxbTOjvuijpkzooWHGoHWSHi86VPx/2ZBrZronrw
E5l+1+MvskhYut3mpu8oBlChqjgmk4QXAhaF+cZC3nbdn0BIskdOMkMJ3PAmOEZGaECiXw/yvWmR
iZuQK1EmB6Vb8tKIZcsLx06vYKJpWJNZwj5ca4DispfQxKi8A6utbgXU6FFA1wyP6RBh17c3bXJK
WuMHCY76OFh2wVvgVRiH/A36ws9G0Iw4abuU6M+gcNg3u8Kmi3bkqywctuJ6l3Lu9kWJvvqBPBo6
SvSB7QQpFVUfNr5fTJscCrRPF2d0CdsbfHMQYEod2UR/f5ZlPWFbZuFwSnKTFbRAvct6oeVR+sX9
xgMlRsZHg6FDf06cEj93gsjZDkkzTxjqJrtXYd1q3JBnvKq1fo8uz1JZjfDLEIOusVZNp7HRTt2y
lpSsv++3ls53l5SFd4BOg6PKSyExNgYo8r974kPZEFyn0i97jv2LEsmpw31GRFb6QLYuPxFRRDNo
u+eIKbtl81FJr/zoDHYDOsXs+DX7spARXccCecvyhuOSuTSYGxLf/lzOvbjhKjDaNOiHJa1sqHMC
Ebc64YIIbz7qZ9tZQ/Tu7EAPxtVDGKee4OJHV2F0IDg6Edo4guu2VtWcQIeq9Bps1nzWUwyq230g
/M4db8UG1p+8hzVfFyiiI8121gf+kRfSHNrpe9+lpA1Vxg1ih4jorX+yUMVINlglqz++cz8dRSf4
ISApslaCJ0xUaKhfv4l9xTS3VkYcRSvUjARm4AfAbdsyyisfdkfMjfaeFnKZOlUpq/K9FsZex+sz
2KLDu4spJpoERyBgSmEVPHhEM9pRfxoDrpRzK7L2eJzLXlEQ3ElUTc0y9n78w7d5957KT8z1nHiS
qC78iBp0/AIeYiU20/Nzp1xQyPHp10V6IMw1LAZ/Qy4Z9/ksgUL2xe8NTm6kxCuNOwdtGMr26GMT
O/NX8qAv4d07nF4OriPRaaGaiwY2yqxc/yEIQAWnm+XKKJ+r+kL3o8q6rT5sMtqwReYxrCWF5OOk
ycI+UF2M9hluQuor3k3yOrh1MiP1xtg4Jmvvy4Ma59RbKJa0BLAfBPxZyShdYgc3Fqppdqq9FAmf
qQqu4IecvZO4+bePQP96Na/Z5X0KCbmkT3xjB5Mv+RZmQ8MDd9WfZQEdavTPFVW7P1sJf0opjQWX
iYHGi35Vvr0j96Nn0/xSrft68wQU5phPZtyib/CWntjk5y+WQPc2TKUjJhn8IU6i/BxGPYrYfr6d
6qZNuSFWJD8wGroMLkTGcJAWf6oIXIfofT76Ir5y4QL2PUfAQcrM/x6Heern22YkuoVWBWek1OW8
eOZPdexlJA5PHgbNoX/vRVE5bXHLuJ+rK1vnkrtVT1sk12AiN+CXGPkCI+Z3a4PEYf7fy51SqEc1
NrSkJBtOGT1dYITnewxYa5UnoTf2SkaG3+/LsHThq7/wCMt2oGWU9rjk6687k25pX3GdVYtUS6kZ
50NH2s+gebtGhtm4fdf4Esqk0YsUtMd93JQsq6NG1H/d1Cy3lpJyHzLWb9UHHrbJ/ziq98FfRteq
SEWaDwTnw2WI8gISb4y9CqHQmninAnlNT5TBTeKImYdjTbaw/588I+y+g2h7yw6DmoZPgGwY4Jip
GQ6IDDTXDlQ+j54utUDWOGgf7+7ka4JmJ43C4I4AM+UJsHmphf1gMh2WV3fKb9q+tajCpsSa5YKN
fRThpNqEIOzmxzVvtKlYUNguK6boqDmNbQL/1UI3u76vRfoFzveQ6OfieQPpPgPHGUrIiVqpFGXp
L9752x8dBxMZHzBgReZWH/Ndk4k/+MlkuN0eKC6+EtF++3u+PLflP144hm3zmeUq3bzrbToim06n
mgnINBegJxX6WEb9pZZFBGaCTfJ8e/ab/ZrbE/oxSvTrgNzqpMJHqczt3WWgD+Px6QKcxOck7jKQ
MV6bUsPXfgbfdr4eOTAjjxe6IpFHNeVVsz5gL50vLDSze58HNd/hNLoCd47CCMnpl843EtgM9a0c
16T4KkSmtlZsFENf1X2+EYHEfZFJNHscZy0jGScQL0zCsC33ixdFQyFyZSwUAtpY9PEWoH52vjRX
CdJcs9hauX9w9NPtFRG7dF1AwpcsdFkKzH+WK+U+v+ztD9B6Fo7sBOYOCaiyeI+T5vzLJY+ONm8w
XrEuaFbJiZcMKIW/M9B3tjdL9wkjZTuwP/otnVpmJwgqs0nhGLmP8eEuqsjcmgmDS9A9tcXNMd7S
KEp1UGdOdNDXJukhuTFes8y/OqHee+QuJ6RLlT9K8l0wTvK+dURdC+vnneQUe79cKRvE7C7Z3Xh5
p0HdU7nRm2ybRUALoFaN7RiPl+YwNursNUPUwmP09uDmCjjC096FL5FWvUqsbuHli/P1zozr7Gg2
/WOVs/WBaHKJpuERIV8Gp0p4mUxUUng6s3Vb/osKVL6hkQmVDxxforkIKAOZL72fprngnHHs3oVa
5S4Ucf0ITeF5ck/h7UlW6TEyJ4q0VG/gJXE2XlBHMQFen47C8+28mOnLefFMx2+hT98rQ83urtvv
EpYTUs+grlulfWwN9H1CyfEfN9yeVGYPZtmyu623I+wynODFaJhpKG925tvDGI9S4CLTVJePLdpN
dtORUSsLTb4FbxqXdTxisjp/KTwRjEFqjgiv4qXahssnAhNMe/rbgvFufjzo6IuswUuPqdC+6oxq
7YWXDoln6mH1od+XQ2DVjAbse0l2ZQQ90Yhb39r6gkDPyRn1aTvtonjfSzA7H5KBwyhTChBGMk/y
TTrZ23Fvja4AmJ9KTcs/rEWlerpXieTvlhCs6vLjNKcwhRheILKoCfVsURogf8Vz/rjYQtn8vXWD
iYga/LMqr/sA7AIyN1TQf/OZnS/fuEXWOQJ3R/6cKN/KD3BhJ07B7lnyzEJlKek6hvBdoGqP6tKe
QB+UqJYp14yJ9Da9CGBwfUfS2dfkf/3dBw89ABK6rlE1AUqh6Kh8RCuKEnGVlXGUGbkF6FObHMuG
XR1+31AZRpibYxUjJ+OiYI/lLvCPCFE4ucrysUJldguA44D7BWq1WBzBKo3NO95AzUx5zC6/YegU
i/S4JZvyuhiXI1BLbBseU1yB3RBhmyR/K4r/4urUznigrzk/CB9Rwcbb/Dh7QgseE94fIPXl5NGh
cgJ2kZfXjYZSamhw2w+HVtKFt3WyX47oVAaVAZnCd19W9G/6fYOMsP8CKU41QoFv/22jGlKQ29bA
wx7lXgytTMjX8aQ1AlSyZI/6sL4LYPxBmfqT4w+HuLM4qplgjFcJJTVYlngX2uDrRdIU7JJKm7Hu
Ind0yThGAXM2mbAS38DEen+XG36sALQaCgeKpKCn97tFAmi8bT3IXXzjqoqnWh2fqv2zGkuJw5i1
ylZ26w7cIikxPe3xLNaJ9yvWCLVZIetYtmEqgOO4o68HQMaMx8hzcoDskXK1XBeZn1nw3L9FZay4
qHf20PWwHsqnWxuUeh0Aws2T7zfcKFAdTPIZw6g086smp6Ysg9dOmpfzzlBhSq6TUK2ZLRf06unX
PhoF0xZYJtY5McAQl8avaFREJs12y8wADJ8V6s9KbGBh4XgXl1xpzyINHDD567fg8kTR7siq+bMj
LRpQMH1HjvgKwNfcv6OSfKrQjnyhPx8ZXVk8kGlOI9jmq0tN0JRPzlnUQYgPj9b0515gyZ3ugZsG
AW37owL9W83u0QQwcZ9asNNHZnbI6+2XyqcrqJNrldL2xpTxCGBjQeHIz1JkVeo2ifnuTS8Dcedk
z3FZVpO9ylFRBSQThEJSoyN/xwHMQ+I24SCRu26lDrRugdNnLmY3HYPvBjJ2YiBcjeCIiMjxoL+T
aR1ZxdZvr7+cxXHdVy48JegZkPLlMUO8FOz6mI5uf88+IWdGSTWHpcH9d5bjVqtZXZC3FD6ykv5O
MzYi32ffgLNPKqvS+/xzqKKrOPm/i/EiPofW7ZmxRcfgOQymYnbOuguIFs/yXpyQse6voEdiQ3az
U8lBjCKVSIUqvqKUZxKQ82D3mfrvvPfphKjCKc2TmQx6Xa4BvkhgEB5pWkru95kYBICbkgwnt438
XKwhYVnOeIZ0irCmGWCRVdWOGiBgkOgJ5Gq76dRtdh5kf3QJw6wvf8bZSfBvaEFz3xq2QACMFQZz
PboaKDl6xibvyUAxFkhBIdqnIsNz0icEOXolP5mWg853VFjSU+iKI1HjOXy5sttBLFsX2jMAuBn8
9VS/EnK6G44e9EhvK9wYnpJbpVjzWp2JdXpVf18qM9+qZofp3mynGDF4Kjb3Bpu8AcxoKyk8geCv
pbzXnMmxeysm9qd9slo9cZdrD8v0uUzfxHLZirx/4oDsfj5ca/0zImO9mS5P0wnzVxyy13+vTw4q
38FrPymY97VmqXrbws86B0AEVOElPszo3I88omho91081zvR7WJ3y7dVHWum2FS08aAS3V7NMS11
IpXXWzfbHRzgaNKElt1K6FltYzYj4kXcVllmOUY6kkk6jTE0jhd6j09yuS+yA7q68j6+xBH/UxKH
s25tU/xnG8sAgxyXRzzDT182zPBnozh2r5HIqifO6l9SOfyx/yujO+kgH3yw07q/7lmvKYDkU8qq
aI9doP4mT2Zym0HXXy4wry90La3vWxyBbS2ok2DoUlHqzrDt4hUrsc0s9Dp/GAkvz4WU1IIEINzU
85pfU8nDMGwtYhcX/YuJQyRFtua/kbcts0mpLjg/fd4GaLNuUgRrKKIYbrlIe3KyiJ3Kn29701zx
tfIIHP0ODQthKb0WyBQTv/GLMzI904LUR+bCl37b3uQLqkP18dv2QmMuNFQk6Mhdx5NdMXT88evU
deKY1dMbYTQHYyIBXE9xntzNLcJg7IygaA5PxDmLMhpeK4eatqoXOFe+sT80JZWJ0mQ91nQlKKq9
N/xd7Ews27r34TnAOk0og6PQZHhDea1mDHw4B+KdndJqhlZInX/H6FqxztReBsCss3WPULyzVCas
gE1GMiDZSQxxkZSuzwM6r0/7uXKNRDKZXxX7m/x0vSjA7s7RGuLa/tGS/k7+PKrKr6Dbej9fVmKm
SSvPfgnUaTt0p/NZDraieTp4S4Dc6xzTBO5Co5lg9fZ8zHlaWl9Z1RKob+7mGhqJGgnGXi1VZzWf
2U5lyYtrid14h1JReCKl2En/ZUw7tv+6Os3ecLdhM3sG1c3/RA+knHA8pb/y0zKDM3HDDfzW74sh
HMZqRQm8UNY+u0SRnE58Xt1KTs4FKPYrxa2rjEpMtUnsvojLvlRQaem7gqxMa5IuojWqU/4g9nNP
TRb5eD9E5YxRFyR0Mt5JHCwiSCDXVYwdaOX4XbWBz3cPanNwUzM1cYK3Ijmhh9+wtkFiXmjnQJX0
xg52ggdvbsI8ovGqMDN2M3iM6CbXyXntwMS0Zh1gMehrUvDo7xRojbbT1ev2P1u190a7H93SRwcs
phiGJVnBV/CYJitAhpQ2+avuYstFtPQqCy3ktpUnmac/bJos1dis2OaIcx4zWtvxvYrU3ypv01dF
ybcdF4Hc0/sEW+PTXUln9w6m+HQKc/yxVDu6svOIOpuMxCUmjT3ZfxIoLmTrOunZNGkW66Zaclp7
c3oz0yhhAZvZPxxgP0YkOy/3ZRZi1rhV4p3E3n9peH9eABX0cTh9gEJU0yixn83kEVjJROvJNW6+
j4YTkXJUryAEPj51XWomMFh379LB6XNpIIDwDoxRHpTrqtp92K/BYLQ7R+XB6J05hIhnFcB+TWOx
4LE37XVgqqM7xluOTSRMjkGgx/w/QggJ0X5qTAzNfp23TB+RcuSoUmFQ+UDCpcjW+gdnA1lRDEeU
nWRWyGYlYSm521VsKs2pbmCKiLzAtLwyHnCayipd4exuSmjg2APB7UJt4tKs4/rT90PSbyV5/YBx
Pf9zt9zgx0v/sAC/dZGjWwrRhWW2Xj6raisLdJJ7Wvz2MH5TUfD38lSSwuTe7bm8gBBrOsf/g61G
U5zSjFgy677EbhXeieusJPbVRuzF0qLqdeS/bGhzdZMR2clfWO5r7xruHyx9STH7KaXI44KsQVku
3wWhakuk9XhF4RiarFg8YJw66DMxqJjfuUYsJsZKEy4sydYUTCv2aIvUTxIvHrjX1Ppco3lkDsGF
gjty4GCM9SnFNSLKCIY8wmm4RNT/K+K9s53zJDXvGFgVj0etXm5hJdihbW4eDzcA2nEvu1raYzrf
2ChCLa4rIw0aM6q9ZuP+raUSPbuhZD8FwAYB4uOMh+CgItAQsy9P/Hn9qyLeKYgQ/Fh5lLikGQm6
54eyvGmbQMmDcN1nNj9vNsF2njBS1c1ZOE/F1aTVp0JAHiYqAbS190pw+YA0uuuOI/xgo0X1SlAv
Cqt7DVmZWtNvC+AcUXRR47p0n8lkBDifi5uzmqWjs2dRrDBt2iRKbyywhlzzlHK/J0WUEmEoB5hT
htVlWQrkGlSUjd8LZnkJcIHyzej5+KJThB0BCHQ6bLdX7PnUlMp8AqMa3a+ZobnUXIrcv/XtMKjs
mFONQeVcQdCevdbG3TEk2Y5BRAF+uW1ub1eTi0LPRlPkGzfQp2dFhS4kIi39hpwDd4kEWQKVB+R2
qd0kGfYV017rlFy9dmFg1DskIRYJa9bVlW1/xQcdRtQwuyNyP0BcUDjNok/xOWUoJJ80OKhZtaOS
Wy+N0NRd+i6bSuH1zoQcHOhXMq71Z1oUwVjnmJ1q2b3V0QcFGwrvtzwe43Gd2d6XB1nNjmkhUhwu
ZQs4s56Bwzde4QwumHLxmIO1dDOsmrN9oUZqccIghseIfrKNq3cshXVFqqM+Ly0Sq84gTd1ki0RF
FaQ9m+0zwaqpU/9DJKfNs3cio747lrY0Oyp7v11mjJvm9BJbYTmvTHmiv9VbXDImJEiRnRg4Ow9n
+PkZgJVmUynCasTLwiszgjm+xQvHQAKEmUY5GYB0VbBFElWP2N16HGyq6teUG/hOoV34EU7+Io9C
g99yPkB7iHIiM/eU3I7g5j+kyG2juUKgjkzwKCdIZvmMVbYllWsAWIi0RhxpmYY6BI9w+GJeDRXV
CVRnrK3mUHbXgDjSoXBxMnJv0Z0F3ZJJRJUqvCl4x/yHIEkUvBIhevu95wbSQWDxCVN2WWIHFgOg
FoGqRrlhoTQDC+w8euQnH/hkQBeqv/4Zt6J9jatdFN1Q073O8zNVJcsg5E9mP+1hRcnDw9Ac9Iv3
ejHZ+3+6+sXDmsOIDd1ph7Use+29bx14/aB7dw3Ek3B6WeCpsPOmVRWOvLliZtKncSdi7CMx26Cv
GDguYeaPsy48qrgr/ZFq2N2SaiQFaEXYEUa0yz7nOgZy6YusuI1TDuhVAVcU5tnH9U04h+48CPdF
dA5yiMtWyZBYtRNJu8q6iCHkYI4G9K8CRlCdY/2OUxyZdulhyv+nWrlKqPlOKORRLXjHjlCyz7oY
+1NTc1v8lNirIeYAV0pjrLc+Ye17QFUf//fpsITxYXCMcDeef89gTSA02lAnBihx3+1D1Zeoxur1
BZHjCDodPOH0v5xxWMVPgQaL8iW+Pofit2R8Oo2fJsP768tBDqeODP8ixBIv+cQZkPdSaRrqVQ+0
lwtI6C4yBDBdrilVtYzKMzUukXH2oxL4Uunx3XVCyWxNnbAPmDbZek/XCfsg+jk/wlsQ2GToKmwH
n6J1YQ2kSJl6K64pGXnaEnX69tCaWj4lu1Yc2+euU9VVFZBbb2hrcdWqEufRBDa1/ExU8higTsas
pP3XHIeTqQ4EENPX0AQBTrZ3PfA76MS7UOPwsjDADu0JwdxNgI3pfdpF9BNCEbs9eSDUFkYUvOJI
Wd2psACeJv8D7BSslGWi0qgANJPnDtHoL/Wo7iRx6R50+Nu9syhKImRLqEB7hrVw7C2KGjgpNFcD
FjDsivaE7uacC2X2Vf0KUi/mFMzylE6D+JgHooIPB+4vQqMqkJHG29Vv9T/57/3BgawGJV5izlni
IIqNTKYdXM31/1HR5zKx2eehiSUawdFk6+0+RA2+bVH9Z2KN/vFq7OzrDwqpP7Id0CS3vpkL2yf0
5071Tu3geEqCVbJpmEOnBbnAY9/A3KdkcPPw7cA35GppYaiTTaYNOyjjgUZSc5nLX4AFAhjFol3K
2gyVcQrsN2H/6k8RvIPQOzsNarxVWq5IVGOJbB1l+8qOutTDe7KRZOlKe6sOCgRliyrYrRZzL1DD
uzjr9iqWz1nCwKmtWtTBg8k5OSPf9/ibv7zstFh3Nfwyz3piIIFrri8oSr63klCu8ObwidpYYmhU
eJ7fKPFsVGSdXPQA8w4GxlMBr74H3LPKvTZH3XwXkI8oi4fQoRF+/PIOiRbsEyqWB1Vg61pBzhez
1Ec/AlbkrUVCsmL8tBGgUZwYocpH1WrxZEC09FlJPAPaQMwJDHx0fnE3uHlBjyQtxCKUMZ9Vx2dr
5g8ZmcV8NQNZwbRd7AP32gzNedvPi+KkSK6KZr23GwfkUsJNb0jHBYZfmH7FVQ269bi0BwZGHE4F
sm3io/QxqtfjynrwzcB/qfUKtSuyj3D88hemStFuRdAMoKiEMJ2IA+/nUZ1VRBNYpt8fGRQ3HIKy
EMKf/SPgtZpxGwIUjFiz2pOk34ST9LoOcwOuEWTZQVODLOCRBw0DkTLrpHhda/VSy9L3B/+tUrOs
j7raMu+4nOJHoVznLbDKSw6SQS+IpUuoyLYTkS3gWXJVzJ88/IwmzUzk/Wu/xf5FYtndoJJESMzt
NeIF29DkDSH1kdCMC3BpHZdqNBE3+mOZA1985ZnIIrlM3Mil/o3wI42tnvcV44tVr4cHCwDrbdLf
aHE0tOclBTagzVurNwxfDBtgYnUqdA0cuJcmIdkz3djJb0ixipPNq9Ujw0IoqQYdxO43rmO3dSY4
/BjvFQBWyaVsIBzHBINX8oY5EjEkgQGR8JViV1nL/pWgNk5VRa9k2p7e0lnnlqToDUaUSL2s33vf
WxaAlgv+/wdcKx9SxHAsI385n5x0wdqrA2FUDyzo+hmluvijbu1NJnVD+JnAlhsJOKHWTus5tJDT
wZbjz0r/V2kVpP7m/XmfQ+wV+twdvea7C+Q0uQCLF19hxr+W6pUC/ncMHIkJLSe76KydBKRF3yJ+
i49+8T1qg2WrljBiBUJr+/AJh19mhyCcJLoYDPipXUkNo7eRF8yEyLj3gWDIk8bSiU1/26eaEa6V
n+5TctH2PjCp4xP+I7J/097bsaDxUdl1WQTd6CpKfkjhorz9BKd5iQOzaZpc1ivCa+dVXyj7jKJ6
HxUIUw/245YKWefCW0fTXqLK4Ad0FnUxJHRNwprEQjx5sR89PCt5uGq35D4VQUTydSyen9ghDgl6
k1mSaw5mYFAhAjMPjYWa1I7ktgOaaTFaEjCCeqKKnXQtFbrnirsrSa3J0CmwgbQhKby2+ZdpY8nY
KyMwXbVZyhHH17iclKn49V9gjF2mrYWgU/uHKzUkOBppY4pGHE3cCl9lurIIjLxk4W8bLuvQUveX
9IwsvEZvogzwB4MK/7jP+xIYJJUypD0H3LMHUvk9Lprzb7kQZFy0Urfs4bjlTceUWkXneIVeTC07
ux/2o3yHJtb68lIaaM2iuR52dz4RnL/j0deOliSMZqiPD7qLUrHiYKUDhzQe3KbEDOPHp9QFzndd
5reJSt6pcoUpbGSdF/n0UqJHVNF87WznR9fRSZxffadzD70gFK4CWrwPRwrnLGpj/roWFe6Cfdct
7TMEEDAsT1bSl0uL1OY8iB/Whz+XJzS7fD18K8y/NVcS7xoBa5/FG+M0vE8d2qBKWb9hl1W0JinP
sZF5dVie25ONIYevPglOG4rG1X2HXeM9bqORLXsPDqS6pFWZ1xT+Vkbmmff/llYu+QZgALAtgr7Y
cibbpJFIJc/GQwF2qdsDVBMWCrAl9FY+6T0P/icBrZft+Q+wGeNtrGStTcgT3wLvdFGbFn5LsYE9
EhdYJOAG5odaI/xGJVvR2tzjKmBT23QP1lTQvZhGQg+6/bTO3q1PJ2l2WJXocgC1gxR7SXQl4F70
J6Ww55lo21JYx70K9WFAAc8hnmon3+YzcRlMA2bR4bMqZP3k1ZnkZzIRFIGYpgN1BmRVA+MfO1/1
50iSIGqeVD/Bo+y8WgIodaO3n2qL8ceVgTxrvtseqleDfICs0uZr9bHHJoEsJVFfZ4wxGrPRB8uB
ltJCpUOACz3W3EkynIAqLUP7T01f1QnYI9xW6Wxk0Je81QVLRe/BvElDBJmFPk5abnkbq4tF7wMd
OO2iBbl5Cfc6TRomYazxhie1O1Wec94r3tmm+9tcGC/69FZuie9mBbS+LoRtMGpJMVP1bJM8yuIH
RNxtRdRYuLR6N8UJPx4q87yfyxTcNbceeuBarmT9NbalHvcrdNsWjv/2HbSifE8mlFpBDBMWk7u1
Sj11Xc0oyPrL0d2nl+BOmCa8qPkGgSSYpeCI2HHY83uphVCbpUyhHEohXytVMpZ12SVkzZet0fa5
Yxp/xi1Z/pniFDsZ2t0LDlkNOddbFGPkVCz041lA9BJgb8o77X6rWucF7RSQhp6pVqsJUEi+JwcR
nLkjBgnI2tC9rH1Lcqw0oERZTvcfbGtJUfY5aNP30UQqk4J+zvGWSbawjVaRLb2l72NP0fc4m0Eu
c3qRlzW34ZxKUbx5sWB1SY377vtpkLx+iYqd650fB4f1sZSDThO7CPhWHDfZ7Le5H0+sULA2cE93
P2mipLMscNLxZJ+xb35QFH//IejUb1LjIQUoeOUH8R9Sk2ojsAGyQX+OiDLtNdF5OTfQWZvfsHWh
xwV4eV/m8RTxdd4P+WRVuTyYCysdSI/FOf26apkLKOCVbBlC8rGra/+Gh6+HVWutzv944qEwphnX
rqZxiY3ZZmfvQ7d6HZ64wIZfbSfohFdpVax8XaGe3s4CYH1a4WRqrBI+F0ArRBN4nOR9pS/jNlrR
jWwLkZIdmpIjRoZnNAVNUVOSTcjxuvHyPxIhrDywVLBtX4CXk27Beo5hqzeSvo38glqUxMD11z+U
4VPtBpwM1I3jvV87MVGoHdzzuFz51HlocRehT2zkBbOEP5gD6s6jl0wctNiI+pawb4J3HM7NfwXu
su5MJu5YCI3/211TrHQK47Ari4sOpULrKJejMDO0YqUwbR0zs7GZ6iQN5QsOtdv4f1n7Cq7lWjNB
fO08smSJHu1+MteZGSBIxoNtFPP2sppDme0ul9mYlyvgcNCvNI60NwsWBOxjF/mJJNcE7DOXrnpN
UuuN4L43Bm8sjYUnzLVm35kV5TP47GtdZb2BP/ItmOi/ZG8wB/No2ZCoGovzDswKUei9KPs/CJa5
+2dNA2UK1SXXSa6MdKqPfNxXZL5Npg5izNObcDM6RUIMlmhnHjpZrByZG9yxb0I6kEr9pXXewunT
YYEfUz5TfznU6oFJiqiiAWOLfWTLMNfRWKkgxw8SmGldOoGJpESmQZyJgYnKSdO4GBD7VggGcXsL
vToHokm5mMkTs6CHVy2WBRpGHVpr7HmJ6frx+Yy4yzbG5fkr4I/vbyuafLUkh/KdDjJHtT9KnwHB
vW5CPEUk1Z1saxcbBPfU7QcISUkAKKXXlOFIn52iojVGTcX0P85VTz9JQ9aelXDxhzYBCXJchNcu
0eri1zfgVjdEh5ZikwcSR5QxnKV2LJ7/6jof4nXZ5O3hbhfcrFXxoEEqknXBvVAt0zEdcPsjKwQ3
HnGUw0AuPqSctg0ScNpOK3uavNltfpbKjyT4N0/93c7BuD1zpPYVawsuWYevwrobPR0kr6ubcQLN
JQw3OC25+iIfLiGrQVbR77imIYEPbyJB+OcZrw7X518UuP+HtUJl45rEkw6b2UUjGu8y/C7GfQ5e
kVZGwpCz9Ag3Iz2pQGy+OBKA7iYLTGfauBAPE/zK2eBnYxoUOHA9L5bEQcDmaC/WVfqMl6YA8kbi
VxXbyfEa9xkL4VaH6usumb6ltKbkOYq/9aQ/KI1u1QW+ip3shNZETcntEuoIB2G8Exh3wWjKPNqb
epqWV/Nq0wdeDg7jhtF50s3yAq0c8lGruQM8jWAIrqdZQqEAfhwSFOUrziMmzN26qusbZ0pnccF/
jXjuatspDvNvaLKlerels67wYRUIxyjdXSRtPMOzbBAzvd+dFQSIbpOnGM1h5uU7/yPFLpO6/+kf
qvI9FRaaWCX0KNI8NzoijE71Qjeu0kRr6FnajjUl89dLJ64qIyMNBTgmuT3I0ulI+hmmUXJtxFNy
UfcyYWIoeqGBK+mZx+HfJ9atwXe3L3shr+IOJIVa27rJUTLONErdotxruV2ePhO38qPr0VqW1x4Z
ogYuYynI2JywqcIuM9YkaQeP4Gtmo/wFGbcVM/QR0/N0qdrqTu+8ntSnjFLVldXOak9cPV3eDd0L
EBuRozYdDOtwkSuMGm5m6tlMCnoY1KS2yjOLOniBqe2mfGNGNaTRbcEYzDtlZEBEAfyI+O7qUK9X
YOCcrF3ylQtpSc3CggH3ITKkdKwFwqzkwLWMXNXPi45UCGYAbVWuIU3uVnzyM6PRPOQi/3UosdmU
thyg8PzzmOiwda3GKxM9B1f1r4PRzkplZ0LtgJ8ILfnrXLcvxGY3PMW+C1IL7Dyazpc0gGsC3Vnn
zGYGSgrXDtmnxU8z3CTii2bhb2qCxop7xV9buI296UbA/OeZ4esy6AEB2xeIit0JD2kQiKAaNiZL
t+aXo2H5GoCzdN1pSCXoWn9+NxCro0ijjeZyVs1yEeju283JTuSQlg8y7iF55imZnRlXBRqmrr8n
I/MtBoI2kcxew5lVU3jqSLeMHr5ps8VzzhUe1KXeUJGIh9df/4K/cjcNi6lbixQho9WVr+EXN0Fl
tt/orkz74vBdQhooJicf4B4vnAEuZJ40sIhWfRN+ayU195UnnmM1/XgG/YC/DWWDUSBBOf3dqr0u
lY+7nUq23XUdoBa46kxMopzxp3kLgfirMuC16qzQQedoqikvXVcF/UiYzidsSGE04C1p5/ZF5xKn
5aJAntGhCTVkAk9mhVFNqBdLQISn9tiyEZ4ZFqx249H405swOydMgZ9SH4carZxBHmT3p+eKVT0s
zLfwT8lEieKpX4zOk/mjhluXYJHB8qBH0Kb+AP34QTwhOZ/I6/2j1uHm6wGUBFPflqpYS5dG/+4e
HtBW+It1TRGVASWIKDivPjiM1/OuJotCqSF7edwde9y+OxsbNNij4IA0RLUb01ltY8b8ICrH288V
hxXxL50y7SWKFs7BpL8TsvyvU+JLOnbNRn7+nf2lhuP+c13KaNjrsZ+KGXVMPd5L4k1VGsl4lZFi
9rgN/JaTZFscCrB2ppm8ZSWXxlGglpcjL10aVZ2sEQe5l8ux+YkBJCkAxWR4GqwJfXTLgURQss8H
yo32ecDfyV9oAL8ANFlMAdPn7qcXjhRMujswF2JxK6/9Axrq1G8kTGu6AVN1vKEBdi1z+bh8LgVA
IOHHJY4KSTZ0Q9y5MLLfgOMmTQO+/BnyTC2c4+LqnYxI06Gd83xiS9a/8aODMnz2TyVUFm2prJ1D
DL5hABRyck+jLCmF4KYyNGLG7vgfIPOu4kmJ/h3YSdC8+ycl8Tp+hcoIpSAcvkpg2+XO8feksSVY
29QweHeR3L+XepT09YJC1ZpfeyneiznSUJQrL3KoWb9s8HlYVez8gZng7Z6SFT07AmyJkKjomuEj
GrgwJaon2zKi0kF2XBvz2QyDyh4P7W5MyomRl0GcMX5TV/2Y4vNCG6l7AwBJz/YKmEpPrD6C7/yK
EWTmW8jAwNeDTCXu53Zd0Wp4DTAYEY4MuXvW1FBPfC+MmvZDW39TGMwn3DlSrX0ONLQ3qXfzgYOW
sIuy58tRdMQh9AtUAOAkLlSU/1uZGO+iePqjjuYeDbw/rFuCj+UBL2DhX+DDREIBBad309wtMmG3
wLHTzNdik0dP/h5fXAbnfF8RCfMbsSFl8mwu7GtqiYEjiSMk4+tdkm3dVUBZX+gH9g+DNktCaYHs
6w3Ax2pgUWZG6Kxjb8Y+ldrafE9t0iosjhxg/BH2GaKiGGZFrL1CEl04FPAvLQW/0J19MwskVwNj
k8X5G9rKeulai2gvFBtTSKnIpt24bCGCV0P1+s8v4jYcw56BD7Je7AKCUa+X/FEedE46hflTKRMD
CPsDNBRn/8R2fTyRUs/lmjtXC9fUkKi2OZ7A+ICVgXY3brpo0FcbXSBZsCezCO2GQ604cFu3KPZb
YCNz1lMLt/3ZElIz1w1Cy48pR4vVFbn6kP5YhCs1PMa9YI+nb45VvXt7NDFdaMsKk1cV+AaHv5+A
eb9A5P/hUPRiX9Ky232/JPqLJbyPvUa2nKpABFTIxAWA4Hgm6n7fr0gMp0SJWEbZK3smP2MDuYEW
bJiv1DArb2UJsBvSrpU/ovDCNPyf2tfn29Lzlh2gDQgrKLYJoPNyS1O1zCtQqg6GIAeUT1EtqrJV
23A+lVYellFye1PwMR+HhaUo+Nn7NEgkAAPvkMdO2gPac+c61IC38T2S8qErpZXvjoUhkhcJdG5i
mjcDOBH7feL5joCsnk55sYi/1pkv23RDlEWwKUPx8DMJL8YtLKwfPFHlFpYQu6kCOR4BNMepRPd5
J8n8rU19FknRO5vFgsHeJLpT4IlLqM6naAXSA2eVXvLwRdZ7QJP00VdVP7rhuKwIdZWCwjyYW6+e
NklIvRsrZqRaKwEVvOwuoprSd1MRlvZ1XILAvCee9WBZnXPPkjwtR9I5yZApvdXRGsupxXeOv8bP
NdtX1psJ8P6HtKBXnvfKQzNnfCmyI+2xZmC4oVDsf2gAbw+ejSg7kTW2z+1vazCDsHmUCZjNbcsh
pMYqhXzhjGu1ALAjoLfHJnBNDfdrFnn3XUx/fiPuOb3Znmz2RlJ9EZ+vxkUOh6HWsAZ/g5dlP3Pl
TWHB3WkMD+IjfXsvk1iU5/3U2x/kim/UzeXvBmZ9dBa4lz+TFgEUAZi1hdJvugHu/1yxMYKd4lTQ
SkMhbAdirbXKSrk9lygsIW5fGkEh8f9ONHFl7FRvsr81SXGJ0MIpwMAnWa8cpOLwM3IiJ3FEskV0
OMDWM3WHWDm7u2M+yuZ2Wtq0QEWJ5+E4yMH2d3zhopwMwFQAznMfvJGWzpgcpQJ0K1IdoDtk/kxr
hBYKTLO4oO0aAcrTATMsO36Ynh43hfJtO72rFAD/D9uvU4k3iYfxIGxIcHPlP7pKlCxTQ/9KwkX+
qSe54TcWgdShsyGkxrppTxXDddQnyc9uUH8we3bFuCt0xQUR+KOkrH3hdVba57f/QoJH3lB0HNX1
vyw4uM5iq7VcAwt535GYMpZBCba2JTfjvult/8CZOLQ6E5aW3Iy5+AL2aosMhpqA589+wUB7f5Sn
L5HilNNGW6P/eTllZFgaZeQCLm+nt9vLCtQqn/Amoxl6c45haYYW7iVlyyEDh5mYbqNpxOyDLddQ
Ws4F8F9hUXRNdzkGVKbJf+HXjs/X9bTb8+SuRggqsC/MnUy4C0x5M06CEaunSBlhs3qO3+7NAgsS
Jmpdpl+73cgN9XpKCiFc6mKNTdbpbo6ruwWXg4B0nblRLhFh1EDfWmd9yYn5rbjPJmfg76zoFxlT
ZY4X76JdgEXCr3O/7A3qnOGYXic7tHLcGBUOhIobv4jRvMDaxuIzcN2pAPUMtBmuX1Jdp2RFAOOg
w0BpEt2E4qV6bgnp8fv1qbWLnybFHHSQCaP8U0bSuI0hj/KD8aJkhinU6ZfYKfS1OQmJjEYWS4Z7
e7AMeMkrYOtwWqtO8gUnXBxtjPCB3PEkRb3+M5x8kATOd5L6oetrk+ZUf3V+telJVnkAZFD5zyRk
aMTkY2neesmIZpjRiXj7Z4BpWEiIoOrAX8gaGkYkZIYp/mxHxJh7MNGnRzN4tFZkOxrcCn/JcRzb
fQ8M7q1zwzjPgCfVSJTKa5RxWrY9AV2PPOGfxoJVxBiw3SzGQYI+PZ6qC4biBVUaEyUpanEceh0y
Cr58DbX95thc0DKludQERa4y2NVDGSS+dTmYvrfRLLxjkwu50kTLr2+WUWJUFJMNcn7KpgAsNtQN
F6hJZLuyAK0zM90y5dWlP9U1UZKEFEbevx642QUGuN8QsAsdC8J5TJYN5PHKL+YvcwB2vl6cKlsm
92K2h85IVj3uUaPD7p+31RwVhMOWuPRlMww56trTeznWinb06pIcpQqMmrhKVz8jE/mVu5BuPmr7
/u6OnMuNDhnI8bDJQBX1XFMJ/keRja6zUVOupCDx9vC4j+2wcxbQJ24I0sUjlBL+ET6hsd1Q1+fx
is3ugDaaDILbbYQE2g+u41i9PWI/mkWTgX4aPV+Ylt7PlEdONtpC6kU/gLA/bYKBCTyRn3oqonFs
M5NnN6qfycV/zcbleb72bBtjaZB1HF3MhVS2tOYaBD4W97b9RDWBEsbDO56bBVT0InW7CN4zmb7V
YUYO1G1bC58H4kLUmf9SbKbjgrRbrEuOU5lZwBNTqP5jQFd3cVV2uM5+tZBaBSOz5ltjeFIVYiPU
tNzzokXOShGekQq4OWhsEtujLYiqMzgcE7JV3+3V2A6otZ1ciJjtmrVO18J9I839W5TdYpjIWRih
ijGxwIe8yiD+Go6k4Ipit9Lv8a/BFTxIwTTMJ/zUKGY9rzR8yjZnqY7quXSuucGL5NrgTFcqu/1A
PF/coyiXo4nKFOhOASi6mJuo/d7uhIiWw32SxL6eD6Eq30Rmm6Rt02n+VzTcQ+yi6f3MgVnCcb0R
uhwyii4/+LUWDA02RqUnCPgmRzblc/MWCfvCZ8vn45sPLjamZj2YzfZiclbdUKcRKMOF7BCFSfJe
FONGWMb4PmqWezin+TOo1G97a8FZsaVgXCdrFYo9v2qsAEyHR2eF2mKhfxoM3qsC5X8zrykS6n1c
UYSHGWoA303LLCUzFiXThF2LV7sPAuNYSk4P70QRpy1BVajTA1PW828hTGwHbFx2ZMpG4qG14rYP
9pe80S/WK5hX21OFODvfU9dwuZMOHbn7hxMdtEztbfv4Mjf8epMok/hTncvAwadaKTGYzmBiXkDW
FBGYPbQ+dwfIbD69XfRZ17M60d6ijJJMIuhCdMsnRmk99paIHQMLR4TbWoVoySI2wrbYlvKFVL3z
XsHLvUynobQQ3zDru94kKK+B3iG0/S5h20IIG1OilgiUpihdGAopWjbtVLVwPk6ZaTeMYnX7Wkjv
DKpJnNny+p+9toEtZPt7qLHB9tu2akWAOGgeLwxaZoXWLtoNbZWAZ2NOvSvu8DOFfQtr6RVfrak1
H2KLYfl3U8pQuEYcTnBqK75DG3rbL08C8Rqv432huMqG5YxyVHExSs6tGmFjWSPp/oriAyYKEvZB
fSdEwmvRLY0Ylhq1ErJuRvlEGUf5AWmz1nL6fO+O7Ea/8G5AejS/rTOMcxaPw02h8rlF16GQkDQi
bKA0GxgoDNu7xjK/yxU8lZnydJRHWCbB1NUi2bGEUN+ICZsw6DCsulfspJ66YrduITrlhBwRZ0a1
MSVPH7EJQ7BliRRjorUSKM11q4fY/YDl0GaPnxWT+XDXVARU/aiWK0fAfKZ5BTwU0r7JmfaAEdGI
lopglEiiPdVk3Znjh+W0PoHEYAVLxrJEBSJJWAwMW/6DLtJWdScQn3jjQ3Fx1EEVco0M7GBj00nI
0sybS2FUqoFPCQw8th9D/gpJhDJo4xdnFkke5wyTFfNgba0qy9hg1AT0xypUabpZQjIHYSyXBdoj
cE8gagfouwiwATEjovg8MdaLUQi+162gsZz3jAWgw/FaiWA11Bjc7Mny8sEEIAdZSK+6Fyfk3d/m
DGbeRvG1A0blj2EbMRw0yi1GXqxFYKFRBRcG5yD5L9YtWP6cHHlvJK+FB4GaG+1o0N+ylagJAeX7
0ZzeU3cJuIwifi1jP4nLWut1u9QtRsghuBQ0WG7vdkUk9vI7YT702DqrCiLjyMLtjaJkg620xrkL
V1Ke5yshMe28tyFruKgTBPGzILYtGsdQl0UQ9xR2cFEs4m80FruAqkehGK6YZC+q3ie4JhfG+Qiu
cwdNutNwdOF5WwSq3RACXcpW8Fxp5pOisTViwbksOUX/i16q5tKwakzJLr6Vz44ov8w3sQ9HiviU
aJOMACGMi8dMM8h4ArB2Hoc1zPYf+RpZHnR7a1tggocjLAUWx2+zz0HOMx7YJJE30Q8Kpt3EAu4L
GR/ge2+imaFmqcadhk040BwRJno4ze2uVVtJBP3r7bhLusfwxrTUNaze80HISGHVQWMJdkcES+H/
dOYieJMEGwT1VmW0S8a9A8ZsWcpYmiGocWcyyPwmxHYIyKFBYZ+nTahdeoHoakvKFPxV/cndvytE
IFwD8qNx+ZZDn2gcJYeMCzSd8QZJHAjMzWzboVTidrHbqgvREzv13C/tnZcXVHcJN4BxZ/w7dFFN
fzJBllbwTm/B3XnkiBsCOkzTI2F89bNXXAoQHRPtf/YczkRafvgDre/iGMvalbOprSN6h/ADgAqs
tlFXKUuSvMQbQfN/PLY9QflgVNAl2y4Qc6sietO0TdTQMzJFgqPPa52u9h5JAqvEk+iq81hEER1P
r09/4tyYxwqOy6J708UH01Cp5wKCFdrxJJl9t6RraY8KrsFaBMeRsNhNNps1rGlQ6HHHbf5h2M/i
FxWJOsuwRPhchR79Oa+K8vkE+6PR50Eo3hUl/7eNvPwhe+Y1SAEAANOmksLGdNTL3Gebh8Rcwgne
U6BO9Y1pv2bH94t5/mB23ZwvoHPrSEY25JJGWB7oTbedB0tVKKhalB89od9MK+CAzl/gsb46viHk
WoXx272tncReI5Bcy9cj/DG2EFMySBEqFMHHJu6jX58IUD+DkJbmvtZJoIVnPIVCAnRpV2ghhHRp
8xGbSxLhwaLoiECzlgvUI6rHxjWckiSwO775tYVXJsVx9SmDJ68dd6LYTg54CIAulBcB0a8mNhS6
8crc0G1T2tC2dWHUUftT0tIs7FWmHD47Y3KNawigsfshseX7E/pTOqWHlsdvmMalBCSlG2li3853
+PwvrH3aVb/OtB0QVDJx4TNmahbV4WJVIjVGxgVYmKVOfrwEhr68DG5volow2M2Mxyxq6E6rAL6D
OtxGXGgc0I42V5fwZOvQ/tPcLJTkkwEiGwc2YbJ6tJBJCWHuchI/SwqHUvnhvmyyjD3bLs28941J
UGPf8ZZGjY/C6dNk9poqag+VpU8SEOLx4MGinUH7Skq32OgIZoT2lw3TwllqeYPJZcVQjU1aty84
YHHpvqhr4KfnFijYOU+asoM78R7iWQgcot71ET/Zlsr/pVGATX1agz+Eek8Bxbsl+qoO6d2NVst/
rRZ2WX/tDgnjrUAGZxwxtgzWXbomaX74o1F+O8vSN/uXeUiJBOrbR4PB1LqtZIdjFdxUs18aeSnb
Rq3+4iOT7oEfPM44HRT6EBqYyglmWMjbgRusv28vh99Of8Ah9C/on+YdaK2GmUBAu7PMmRB2wI7K
TasggVEDkJvC6C52865qjitZQQWb7J3XW5uu0+87PfVMPYWwYe8HumA8bkijQjhK0FqWhYEQgcPX
odAr5Tm25+lRm2Vx+CmG+TjRpI/HiQSBb9t07urLEYIkvKc+8qfIqrtrmBfevZefSBxYbJAN7SxU
+2ubiRy95ZdK78wr5vD/A1BNJ/vt2GXNCFhHZKYLzYcH/dYTnYvCf+ZYv2AGMP31VGzVhx9b/27L
o+eWj2q8AIkrSj6BMmjIVFL5ZnaRSZKDwaypgJ/cW0NecweOPfLYMmGZ11ho+V6nndSbbxUjSVpn
SW32ZrrLQtbdk1EjAqUsTaXGOFw66bPr4yfUsIm/NkybosYyHA4LbtweMdNUFMQuaYrT6dbpAuJp
Y7IUkWu34ZgaoU6BSq0Rz5U6sYON87gTh+Yaewpm59wphSC2R7m10yozHd41CMxvZtKoTY1OENuO
J99kP7737s+fsPUHxOOSO6pF53aBR6ptrpxZFd6SPxZzv9llaQPHc4lmRmuf6AJCRmXXzekQJVbF
Uacf4748khSkFdV1HWt/Je0jnKcJfUZ5s91uyznntBUVmg3l9zUGrETuipqnmLUcuEHwqhSq6Ys5
yIt7Fv9yai2l7eD5fSaj6DGp4FsiFFK1W0OCnHTY5b4CYorPKOkD6mNesXo9TamNEqguCVBGS4mN
qE6EdIlbBlF5rWXd2Bj+oIvuaPv5kppbyChuPcK+OkLPwmLJwZc2nS2wKsKeFSvJ+rz2vp/5hA8M
D0ExwKWDuuPw3PPx8XkzELtNh8z8Og5al4AYasWGXLs/lNYsxtzZbGYQiJOqb1cqnZFt9U4NXp26
9bVoeFPs3PWVJSa2CXK7A8RhcTE0E+UB7TDVuIEMDAv541r4p/zd2yubnBwyhX8dO7wC+4D2YoNn
F2jxWDyUfEsJderzwpB1gLk5vQARNLrvr4m8hUymub5816hVLXPLPQbQN/RHgWuFB/ILz+4qzxsN
7reCKAkp5zwX+7JnstRpcAa9PXcUv3c2tubAUDQxPnSJoh3486nuY3QkkgaoELsoLlii1JbQy7pc
S+cgX12ZY8ChweVLTpK7PRTrApPJBT9Ym1CKF8kgu8N5MVgciW+OBnsl9QEclA5h+AiG7TzjuB+N
m7h3DmEysEpu1cxhtWCpkyBGE6jzScK9EmKHIP3wbh0hbXFtJlCDJdHqWG9Opkcj4kfIVJFY9lsc
pgXQUpvraD6SIH8n1AqUrd79kNY5+ndPdPmzgYpsytcbtmlwHiTuMxxv9gvFti0e/tY8MjD+TvYX
pgMJsooZpIq1uw/ubzz+3CkCVqBx2gstiOQ5TSbOOXK8OxlGP1TyCb0hIOiHjXRM/buBD3Sf+Dvl
SI04YP58us7L+deHVWjqYqT01q+y11IzqPAaj5NYb/1MFenVMUum4M/bD6BSCfgJpIsjiK813oUk
DBCJ2K92pl/nzpTGZTHd8o56Kjn5bVlTtLevTe9ntjgdvXe1QwCZjTJVXfikKY/mFItJDEn88lrL
D9D3a1tploczpQDlSC3D+1U+H0vEtz2Oj/+KVRUPNN5cPbMMXYceqCWjxMmFTJY5HLdYVvt1TkLm
OqlsX/XGJCSDuFGWDEZzQ5MWAaF2w60zF1Dr78CtfaNtyFfxM0CP/evqpO4BW2ZDi63v5y5s5i4/
gdy5pCJOhbG6mR9pHmhAvukdKj/NAzQX2cL1r9IUMziNQ8tuMLJcAdqeE8vzemBFB6LNJKA+yiOZ
moolTy/CnBl6IpMCmr/vQjpZjRv3WZc/3l8/TdzHwRm/lv+gIyNcDnuNJB9S2WX3ni//Shrlh+Pv
ukc6TVlT5lJ2WVJZlbqMcPhlfgYD+2wRihwg4+3YMxLfTO9I2goBJWBJJATfXqvlZx7a1sRmge+4
bj8/0XzTajo2ApUopU5+Dn2lZNijwuFOiJBvyhnhF8OYJXcffNPcI/YoiAc2PU0wda8d+GXEAa6i
ttyriP0hZNXG8eClnuK08A93aFkbSQIZGtrdPa+Wv/gRaDJv5P5dhi3Ds6YczrDdwYpcZIqxCyY6
BkcQU+dxIF7V7uCBULYJhcXNxd3zLPlp2xbEWjRLLOM4T8QxKNDpW89hbJG9t7SRK10i2X+pFFyW
XbY62tST5Bf4+7w2azV7sXalkKGFGmS1FbqzaaqhPuE+2zQofAh3ccglW0tCbpsKhPScdKGP+cwS
gnK86BpT74TczPm0Om+LLQY+n1Aozbw7PtPw0LoJpDeGn7s9vPEGgYAF+RAgCgZlC8i9c+UUEQjP
6Hbn/3eocXWpKhhe+QLDZPspsQHhFh2tbYlU5OKVpknmx540L2twyZ0TIFFukWXQSJKHub1fL0cd
2sfwZPM2k+740GgJ8OWCrP58ZN2eQ3KvYVN80QlDLTR6OdixvTNuIaxqyNtDxvIauiUWMUB3m0jE
ECeWfm8aThGPdG/D1ljj4tEXLtNVBjHm3Lxk9C2gGTVIpcYSixwfvBLvDPG57JeB+Tq22kJ1/8Vb
/ajpoCe1USwbohWIxexeX4rwGq7ZanhjUFapXR+sN0iJPXPqSskGK8v8Zn7xJylAuB5kdmExG4cv
wXZ03gqsnMb+YTPh0GACHQLlibphoXsEjwfCeMfZYxlxThLPbUlT1KOH5esM/pPNALUzJtYoZ27S
IN4zm2NWdF3YOGFC4qcqnpt5ZjjWxWUR9JENaELhFyJTQFMncpuONHeiRLrkRhcgkx9IcfGvdQ3d
tARMWFbgq/nCVRM99GInIwokCAYh5oLhJC+sNZpUsHwOw/dj+TRK+/Szj1Swlxaqed07OQJia/ma
I1rimq3KLtY2LKhI/m89OzjyXG08Bm4ZVULoYq3C5CjLkP4CIxaOC+wRjXzxu8IGfKym18IszQ7L
EHfLAGZGYL3gAJRL6fHY+dVrLlCzS7AiO+rbGVD7ckvdRmA6w1axs5Dq7Bjza6MDwKBP1jq/rrqM
AYKIFZ516yGo8ReUiv9AgbqBbjymIKPbDULBV9+ZTq6uIZaXuOnvfgXSD5Vwp1n8acfC1HnO6Txb
SpU000iGT/NMo0lHNsIKW4oBTC868b3XASLby5PPARJv7AROjmhu0dm7ET4ht2ZyjTYERYaxfnVF
nygxzgmhmZvFmKt0hJgWYW6yttEDacMEkWpco1aTW793vBZc7pIxIKG5lRT1uKCh51QxSokHZSJT
C02Y9mEfmgGFbQ1X71YCmBWlhFivdDX+8g9jqxyAXluJRHK6db+Qu9VNQjMI9n7HI4NqjDStidlx
ZD4x0t09XmY+R74iwGnvh9DfmaM87DkE39XLdC1JVW3hmNrll7jOy/XAW/d2hg7DeuDOZtwJW8ua
PDzlXLqm1IBZ6hkQmCjV90l5OcKpdBnbtK/cnSn4tSA6ypKR0dfp+NSuhNcRCzDyoSp8s9NyW9qV
Xhb7oISrn3JqrVJmkIHcNuh73Hwl+uuYySaS4rWosLGcMHiY+jAckLweS3uchgBCfOTl2Hrm0Q1k
pJsJ8B/GCi0q0zvGyMpFmIXW2guS8XFTgiYYK2+pe0UfzeWoHXSM+pxqIYJIoTQKIkdkcje2oaG0
/5EStKW7+S7q5QCdzMmJrHZLtmpBPCnvTlrsVGslAlszb4bo51kPJ9LiZ0gecVtKCQ2RTwMiqrr3
OEU0FQWanjSBVR458vw/9BAtwCi1MbeiTNxvKRUfbfS475HJ22A4bMSFSdPiBeJOq36yONn4e1lB
4/4MA/DdHNPZiX3ut7rpiGQg0sGdlL+HOcIeOP1lKG9CB/cOmyVnI1Su8vUAMHs1X20kfOedgPET
PUWxJaYdLUrtkZ4Avd4LO8LTYRJ2rkRiEgNOHm7w3Po1xYKx3eA3UYvdRcQjL1+3MTfvlgF1/lvB
7IFhJ35tqk24CCWaBPOnYNw2yP5p5IPvp1wBb68t00iKHVkqUvobDYcSyZDbQ/3j+tVaF/ewj2La
Bah5r68K1Y8uj01C6aG/pi9FYfq1aizNe0aLJO6F0ek/on/dE9EhyJcl+cdLpcrL3Zn2DylUkLdU
iJepfzqmzGZtNOcDPuAuhGEwdex1JDsG4+FZCw2hu0koF3mXtg4mT8JbyvsSXyZbap2/3Br9pKh9
JPhu/nIwhsmq+Jmv/8LQFyi70pLH+NGSLTZAaT+Jfi0z3cd6PvUI5sJboYLxy/sOPiPRgD7g27Bu
pq9W85kDr15+LPAbg3HhQRetxjRgMYDcdAU68UmMnA4W26BMu5JUh7/U6GHASWPt8WGNV4gFghdV
IIiWhuYBpLxJF6Yo923w4w8t96AFAbFNl4PL11qyqQUOtofN8eqHGya1e/rZUqSzioYOBnUv0THu
iSnLnvsGP2S+60hbIZSai+FNIZCmn+H6lodZ9RJVh5iAedvIAbEmSCklxDZE8OIpX1pVDR126Dla
2a40y1XsY8YC1ffpo53jzNGwN6rFgG6fAbybiBUTsBcXWaq9WXUMzbJBXhn7vQVK9apijHStm+XZ
S+UMD/kpAaAcb19yVMRGDSwl8ZRbgT+cDD9KT//Tc6Ezi5vAOku5x/SHXGSwhUDlQGLaVoztEXMn
4tGmCUdAtcDifXnWhb5nD8kmHQSnaM37yFJGGUfKgaBJWlWvb2Pd3/++H3qDTt5HuTt2MMgoXgjn
31EEQ3Q1fiXJ9jVhB5DsXIQ27xO182R3yKmtCiBcu9kUE6jIQlLE9O5qUI/VhoI6VicPEpADjEB1
w50IxsAvqb5jMc3Xe/iNQw+mYsgKLPYQcpQ9F1DM+SJlFVH4dh7vLS+ZMTtduzuzk6wI+uTLO91W
30v0qCxEiGlacgzvxBRLnTHNRXxQJQSLeNtPzLUGPQGw9iPXgDNAJ28yJQnv2e0+hEMmRcrKq+Cf
YU9Cjz6l8RD5/U1ylVsigVCey4oGL158iVUxqJLVlRQ260epz5MVNbhwUYlkOdjPJL7W4qZ0tdGm
zwDZyaKnom5x3LfzC190GIdHHj6i3n9Cc8ItbcnTXrgDMpihcpNEG1bKKHflZsK/O0uvmV6ZVbVl
OGXkeJX+bH7w96GRLnDy+OwUAkGZ74hUNcX1Z+dIK7p0hJ+YxmGeTBrh5nJvaQrhAZImUNxtvpvE
1jr+KdFItspKnitakTkvfJGZ8mCyFQHsmGdyHbrOiP6+2MNHzsPYcaW0mCMFUlXq1HvpBYSW8iQ1
4q8VyfAhMwXAxHRGTq2VchL8zVOTnPVdtM0jDL6QYZEm+Nn7mZOs1cMEVNtN1KJpVOS8yL5msF+9
4DCNCpsmt4C+W+yHtCUH13rEp3iwxN+Bo5q7th5wkhZJXDgom+nLiVAFTlk2966qkza5JeNlrrKP
eBTp2WzW3Bb4DtZ8DD8xqbxG1HpkjUZJorksCkkTaUhjBbf0nmujdoB2pWLGzdpt5s4Ee6FvYZOj
9eBXBSKvtkZmvKDdIoLcoLXjtOmIIWHCVwnyUgG6tOJ4nNHwYxxWMXPRowasFRuL+BctOULWeYqP
TL7igdxxx4HX2e6Lm1JyR2SWVjkffVSGWje3klOxb8Oj6LaxkdRmrV299Yhoniu9eTs176l5AQMj
6lTm5OUXzOp0A64FRjFb9E9xHyZflltHhimDViFKiY+H0W2NC2NaTS08LNtYi2jacrhLcdq+a1xk
3qDQAoLo3g1T/juJkABhKwmPUx+F/y5D1Rmx4AXdJnDnCvUeYqt8hudr+2qqe1TWchDjGUBcmzIT
wlCsKU6TrkhUVxeZRx9dC+5c4Fqy5iFk8PXkw8FMZ+Yt1v41fY+OO2ZnlTnLnMurHydDEFW7sq4e
9/g+ECv6tJFm+EmqRnXVl6mo0FG8artcvAifWiEQ3Nx9ZisFgEi10C0ebjLg8ljdV0FGB05kulZy
Cr5T2S1ZbzauMPhM7dF0reVPsq1kcjHWLlQNCKVnd9puGYIeyKmBmdOSfxuUpbHpYJxITa9nfnVj
Ub3y3+0AbP40n0a1XAzQTWCzVy7wc/EWl1KgFOvndrFW9l6D8o8E6fZFw7XpfUEoUt0Q3+qeB4Lf
+Cr8dGrPWVJGqILY4a6dLedN8C4UVxPTrEefPMASoQNk8iicPWuAJfzfh46X+BCAwWbYp1FWRWZr
kidYX9enTrsUDt+nfYR5CRy3L7FrQhseJBL+ytaJBYLAy6njuI6JxrhMf9ZZs6GXn/slqt7y3G5s
dwhxxh0+/IcgD9c5zlVaB5YjgLNPHvMozV8FRdyjDrVCec73dtvKUO/gFls8CPPkL0ugHtywcu2w
QyR6++1h23CVaowkIXvG9bv25Q9JJFq0q0lMjFziC+nhpKVnOXxzJoI3Fwe14kcCo8Pqot1mS4he
XL8b4YZ0O3gWYH27Qr8vPVqYf6VGM+3hwZqhEbvoochCuuff4Aca9YBmKizsilm4uuhr4Aj777Mg
OkI9/KsGW7fi0bukbB4O57GATp1QZ84EDGJaRhWMwBpURn695wkZ9zznEmOL7i3LA+jl6m7iKsSZ
GOz8QEI2sKI9ayRJ9rvxyvH1rgvB6Yj9igq57Fz9HoBTpAELtTx/v+wKLqBga+LmRos3abYRHwhc
Ux8S7k77X43xf8q1OKK/uQX56jDti5JyChfj4ZUPcskpyDvoXb/0o42OyxSX/IcdiFBPgLIBHqaq
1GibyIzWc73jxac7B3EngWJxsnImsa/dS4oGU5HXpGX0HXwpXm4Xbph1fsYb8gZmcCRMG2LAzLeH
/lGuTqg97+AOg7qM+eorw55DMQD+M+/1f23x8V7BusmMET9KBA5OM2OarG3NAsGu7Ypv48ljimIl
QVXPJrr9DdBvgOluVuiiOzrHIi6Qr7qoUG8TBflku5P+xUW1o2Do1wlCaZZ/PNR8zkdEaVEjBimx
G0EWI7iJ98A0YAUZt/NMCd8vfLujNAcPqNieST6w6rOwBxbh8RQgXptyBt43heiWhZ3tljXBfmfX
lZTWUmUzLf3VaapRkai68cPQ8p7XCLChULwAw5B0W/wcGS8CrSFwm8sdC0FmP9EtFjcLx6GWMgyv
KGHcu2Vwc+vpp/n2/yQO3wh+HTtnz99r6LZAT/b6jmTSjQVD67uMK+zVVScyWlGgJXVE9dv3kkUD
kBJtn5O1NebBxkg8GFP7xD+wECen3Pi9+1Z7u/J+Pd6O4p80JtmrsXpTn7IYHv9gUc5nV6S9UCuD
nnhhvVmAOPxZYhJGZJ2RfB71fVIS6TdSIC1NCqyL8UOdvX5xSrIez0In9puOXb1qnjoMCxAvXpMF
8cYsuMLKwP5kHHOAr7nbpTeB5hf8Fn4v1XqexveF0j8Xj7D3PvGkKaUOuHEMHuB/vVxUrGSdv80+
3mDU/1+SxPvFYkMcg93bmibHTEhZyqRanlQJ/aqt/O7toj692v1HvlgEAEZxGLP+5WcLUXanRR8D
WARLTDn+DPNz+/d1ys+R75KpWN0AgsZvipKe2DLzbZeHrQZBsUJbyM027CuJWx+czGvu8yk1Dp/P
moJJTssJ4cp7mHJnju2QiWne3w3Ac7VtUmfn7qC/x6erI8+gKko5IqGPkER2CXvPO85lKceAD310
3wunSyj3PZF2Kyyi6hdd+vGkHVjhcEtMw+xHJGKb2v92H+jRt+4shVthsD4XUw/xdiJ+gszPZjKA
Uvrh8Y6W4V4siTozVeEdl+YWQ6DcxVsPXG569J6ZC1yFKnWpKWUJOByaTH7nSwr6dHpQk34M7YLs
2t3xdghfiBeQ94WR3ckUCO4dOLCikOua4/5zj4Nrcfr1qUyojj9ug6EAw6C4P+OI4S91W2fAXoyl
EyebPSGh757hQkfmkE0GebQntKogE/1Xk41G3Pk+7FNho1A3Ha7h8sZVhepukV+gXlcf8uCpQTRN
2DIxQ8YdXK66h7A9h9S1eiM7XB3i7WNUyzG6cAdIy+vINgfRxmj/34gmmLMCoS5BGZS7Olqx849G
pT9bKZFd5SVB24WQgmvmeffbyU3neXlLCykUiS1qJyKGWPYun8o8+viCJ0pDghxT5Y0sJKWRje6D
PEprwxIeh8+zCXlWwksDBNLIVKREqAectEbvqCLYFdFkUJRvtYOk5EvCaancTzl2y7+vLtlE6s3R
AlIW4YpHkw/bTlJOEiW3ZgbURcNBUHg1IPCg3jYKoSYb96cDw1YnjQ07ATG7/sMhnxQeDDjVjtqc
XTpJm5KWN+h4GkgTwygU6wjq0jM/Ji6+VrUS4JpwPgouvRlgYXmSJUDt8ufOHPmCpTTYSE9i8zhn
Vug9V03x6dgVsOXGr0BB2ucCV2lZt60SvFTU16pi4j54/sXreo+1LpDmUcB/bhaLN8DHmvZWTbK6
SchQjpBMk03nusDhEinOr1XFk9aTKeySXzwppZxMxwY3S8BFAXz99JJveys4ctk5WwP9HVCksxIh
204tWLuz9dIpuAmdGawT6nWwmVMJ8FME5DoJBB7oP+7e3ptksK9pwZouz1l7xh5IsekHK5E3nCOH
RBT9ZMzKVHt0XjyP5BoTpGsD7wFYx2Z3rqIJuryA9/tjeJUNG0tsz40+N9HpuV16CNsr5ZJIT9Ze
rIaT8PWNyQata3F0239DZu3rthMygL076YAzTaq9PuHTf129ScMRj/TM3jxHoDu4oT/urTIAlvMW
PNKkKXOuPrMjBAHYxT8W0QYdHdfas3WQsgi5/bZt3CaKMeqdvfjFdi+HUjiU7nEoWwBHR8CijfAR
hGsRklgP0Js7pucVE5sSTQD4e6fgboQH/lZRLEaPEPnMTZyf+gxeLiAY/9VF2+SwF7NjhyXvxb4Y
S3P4po7E/Omh84d6ow7rPiCuAPcJsywes1atVKYZrt449bzM+0hdXeoFRADsFC7eDkHVD6e5ufaU
xWJu54oA1xuywk5+NxY54HLQuOeCuyAjRa+V5LwV6pUTHZp+psoAr2dMvLA43PdTjh/YFVf89ZIR
CZeRhfW5ycIW9V5+RpsXPkgbA1VAXFi4F3sJOBpW3hURpu+hivH65+G3YK+52XX8SjedzarLO4Ex
UwhPUNVt59lHjkqzcEKJYlo6CReGKMF8CyRBMR1W6DdtRig9TmP2DCuUcfrEWO03iQ60Lvdqc/RO
4hL821ZQd+lpEfj0eDTC3+3Dl/SQ/7oE0LV9WbCtvbtMoF5HdoeksN3/XX/fLaXLaOhEyKFbjK5B
MtEGq6jL5F1bcneueSe8yl25UEytqKfJYcmBnU+eKur9yJguCW+/PYm6PGKAXFKLp6iGKOnyIC9m
HBEinTiBBLC6GSDiYvEzB9hdlKOfogs1nxgYPN8Kpc4Mj/kpCOLDheyl6ucO9eWdz+3it0K9CZcJ
O1hyOsOtevfUuAt+b6b88CjzcD+DuLZZQPb/9lrGrFdTj7VXW3675DslTa/XWdgZ3ybSCq+f4dUm
rIQtZJSkElji0S2NJw7N0w3gdqCUf0QKIzRkdNy0pwFAQUFcYcwVHeY0zsmPJxhJy1l8hjanLDnk
2Oms2LlAFh0XG5+GvszAW+plH9CnRbsJLtTngF68wSbjr2e+glxN52r3OY/73xYAeir+c7NLrZ6X
Hci1xe0IiZf0sczQQJPwZeqiExQ6ExHh8tLEaRomSWcc5O25WG5lRkMhwIvULxaWSa5U+8eL7+Id
LHkHyeCH2hKE2XWLMyS7TZkz7sBOwisAg+4ntRhiDP0MHH2+vCn5fdG5iH6uHuekUbo5aqx56WOr
hHAntp+eCoyxMESuvxmD31WyZqoalzhvIMtXRR9uDiU1nqRmpQ9zXwnNi7llSmBtG/ePAkqO6sCe
+uX8KPymjYcoSE9JROWKLxJwDBg55fdweqVlOmCG5MVMV6IKp6J2fAPiVKBFkRz/R/Ei4IYHkZ4K
tcmmmyimME0x3PtEI1/Rryxm0/I+NAarIvHUuVMlVbixcQSIJQc3k1Wj/d+w5zhM8UWAL61p6J4v
T3gol6zPGIDWQ5PNXq3XBni13nxPeG9mt9XPYaiZYCvfGJ9PGga94WzCG0rajA/YNlIkgjbXelnv
lOnv6I+ITnJJ1YQj1i32RYZKZiYzekedIu6tFg3xlVwbIwRMadx+QxDdYrbuElM244YccbjY76gL
yHfmtb+gD0FwFZcEHdVpNTfMvrMLLTl/ncDYDylKDktLFt4+dmnrWv5lk7FBRdpHzXHTmF0/JrC3
dl5p82DRwJZxdYbisyLuyWi07IT8Zu6F1D+sZR/PFXLbGNIAHgGsLyeBKfgtL1wb+C/rS70+MBNB
YHLOafcVXLapwh+z3AkmpsF0Ok3M6PAz/aGA0+zWJTnlGkBJ2Kt9xQnXfo2tgcPhKFdH8rpFwBZg
eljE+HLN4Z6T9a5/ku0us8xJYPMueokfA9ATcmMHAoWvOxrfBXinyxv46Huh6ZVVslRpilXLxaxj
03uIrNTS/GsczaDjpq5NHE8kIR3PDuwAKNnAXRJ9fAjvqjDTeiOfLuFg/cmugBQyEOefz5huKEuh
OheJO3Ap2IaX1N1HQpiHWJ9ZaJhm0Nk7Q7CdDBZDChzU3b2BVNPHhwPJQ7xYPr2BUyaOeTB31Qf1
DYYcKzZ0RrSMUzgYFBBOZHA2SxCEKYPScKvyQZu8z17SD+YtBUgPVRz7rLB/WaAy/SEzy6zt9RX8
kzRYSwips3B1qjwj7NDYnucoqQTN9T4jmlOI9RUDYQEhXD7Hd7lPd5PrFEJvJn91gnR5lFlQ3Or8
yUG54Kc3Va+1vrFhBbzKXr1YAjF0AXBojm6fDRffpeFoEsREPGZh9xaQvxZ9d0UqymXnGPURWDpc
yL+sx5gbpchWfgBwLrTlFGM6JAao1udkMcGuUX6GG9856vEuU8uwBwt/ArK/d5P4UN4je9OGRsd3
SKixq9ejdJJIVwuEUU9ky2BXuAyJGzj8abrn0rYU8GyaDr50fibtMWfYocS/FJvBYZpQ731QU8iE
KPeWLy2hKPO3cYzODvRPYAsAuzXdd969o+02bk7ctiiHPPIkv8e0iEBMBIZqI9S3lSpJxwOQsFrK
c5IJlv1xXw6ASTuYiic7+NdBDi2/9XyF67WWEioz8sZ9uAAZ0Xq08MLyL4YLD7p2bp2iL7qJF34j
+jJpLAv/ulFAZLxQhc/s1eMeVgcyiIBPi7B6zEtKDLGjXmAqX6rtbgiw+jWWYAmeLxKl9VcOPr/8
wX1vKqee9pkeDt8R1MhdTX6IduAiaDM+fXyE5P6+InWgySmuozHCnkV/I3fpJfTV7daV46WTNZbD
EzLZwjleLbEfB1jQyvFFbT+Zlht4jgD3wKS+naBcwkNfvbkFGxZZmvI1YVP6CsRf0Vdqj029a/H2
1wyoppcqqU1HW268otcgHxy4RGDBgDA05T+zvy0jvRhQKcEDogghWvpMcmThjsybSEPJNAJed96Y
eHLJ0ml9mbHmKbYerAERkSaK0JN0FBxp4jFC09tD/VIJBWtwWFZNxSSlBoaxH0r12VjBR6ce+R1F
4iyYE9d5M0p23kCdXE28P4oaqK1stGv8Mx1NKEYbFI7xSw610dllNPFrYuWVlxuR457qRsNl5yLi
j0da3z0aOFKc54bn2/dafcbk36W3jSctaKHrmLlJxY9VmC7uK6DvDtr03IxL9B+Qb9MB7hqlHh35
GjQ5fAsYR2nBW/D4CjG5potxBBAZnOcUgLyhk5UnQf9xt5SZe/m0oDFJIyPTa+A53chBGVSrl7gV
KfZwgZpRIIyf02q5/tNKLtDIHn3cgknIxmQSQE0ev3gOT935dfK5WSCAhigaS5F+MWTaO01NXEx6
CLWm6PKyHqp1yojkZn7ELDft/4UeBwaub21UOY7ZBLdY7kH/Ut45TIVMeqekremsARqDRjpoS8d6
s3trO7UflHPpZVH+EBprcFk2MjVjLkaey8l5GI5/JaJuPyxcc7UlB0RtCkpwBDigCiCCWAR8+/4x
nWSn5YZDlzdgjZ2EkDLzc/gxsYOuIzxAuLzxgycidBF7z3pnfNVIAsN3GVPA1BFUTMMsWJ+bKE5W
21scXoumJwgu002zGjstU43Ha/5SQHetDnfxYhgN0U/gYd4+KDhgqC2ecH9izmWKnWfr2/wvdvjG
y6YYpvqgHR/Crdr0gkmFpb+Q+9cn8gtHFJHMXmwoYoOfepkx0RMMGbCXHwXi8P2iqafoQegbTA+G
Ma6bXLnnkWBxn/E7UX7blwz+90LeJSwoxB/j/c0/JNHnID98dX2nBooe2S2jB6kN634QT7Dxqvzk
D0tIitavoME1mLRfYuA4YCUn5410/NhhkkZ/AS77JZFPUFTrJGuoVDVy7YTszEwGZC12wKAEjN3c
elmmNMdP8hHSuvgQxDfZ62b9TxIBtJLKp/jyCW/ZwPWrlxdABDYTIuyRefRvWpqQUIn7fi3vz2Ft
+xRsJ0VPnxWtkUeCFHh87ySPq/EZsaBG9DcWJ63yByT+4wcwS9DUu/ZmafzNHeKXpec25pmPDgIW
YGwD9Mali/uvK0s/gqyQa8IpLFsvhNNxzyzfMMMaB+ugYlmm293ePIlsGvE+4n3An79HtboND+ag
Xg0Ic/kTVNn8dlnGfEZ1Mo5HsdIZf3KE6lFqVQlOEM48a47YhWjtJEgcyJBjtNVOmor2C1hbMA1S
e/3era8GDh9kuM/U+qOetoCvPXkwJHylNEbs2SaOKWNpYqTi52XdBpObxEKYLAWFPJEpb+HyTk5v
dIWPWyU+QvRaMzXDsfIA4vuX28NWNsKWQhrQRw7tR2ik949SuCdinsUvN5MSaG+F085B6Q+nd6gd
lXumJ3i31c1/aby31azmrGIACn9v7v7WmYltSvkneSg3yIOE+81FQkjHXdMe3w7PWkuHOTUEwI2N
Bwh+HtdOTscrsqxsABixb85bAFNG57up7ODY73DJ9abXn/+b9cXTOb0py1fJL2Fb8o1tf2UPQbMJ
52iYJwS0I6f/w5IiB9PDLp4kjKRR0moWHVyohBaM92+VZuPaYElfNlUcNwipdZmOUmig0e+BWU36
hdblTViVpkRsoqX/rc7kQI894U+Lctn09uHokpJeVQLNcUGRi9s4HlXQXhjQ+JSMyWOwHsLQP0Fb
qbQsQQVNF51cEpkcs5sMKZmqc6tULeLa2k/NX0am4w5rFuk+/kJCs8+94b/H/iUb45Nlo9xCNubT
6FhNFXsRCWQEWDp3cJR8Oe7UeEBG16uPUKzS9wfUxpW7VzaObgoYAk8uc6qmEqMoWZZiD/9Kdlcd
DtSJdCAXA0uBDupTYs0Mqp+yMpNfREowKyOxWuAeTtFv1BCqNRmKyQnNE5iXWpWkF/K9x3xZBiZO
iZYYEA+8qLSXiTPPzoOzRRtL+ctfOKARllyiJtTHN7Wxhuln5R7kODGsmEhqtsRKnCoAXvrLarVy
Q1AvczlcbPiDHSp8T9X8TAX4zz9Tv/E+kD6RHK45MRl7hXJdgZ8TGmgmOsgWfB3ddWhc/MAwIG3t
YJAVxJQzAcqjfXPiVVlmkr6yKsvh1gNJmmn2HjpftKhvdiadTMgl5H8PszN8ns4mSNDqIRJL58gH
fkuYkTCQle1Xl8X0nAfrASo1FZ6AvKzUMcHSTVUd8mRXfjek6xTDa1C1/CQ0HZUtwpE+a0S3PfGP
KZ5ad/fqN+DVBU1C23DuRnZ+rR14/XVZ4q5hHr6TZ/h05JuOaQP4GhBTFZuboe/zBWMsEiwoY0q5
chVofXVvVQivEHe1sy97OwmXtLQJm7GyTlcu40XXfIdOpfWJQqgcon8jcl/LSVxng5fX5+48HHAe
zggPtYVyn2bVK27jTNhF/SAL7yYpX+BHswZLf75mZ+sxMPLyGSG9puXkiLYQrhHJxgGkmr6AYAN5
aS+xwus9032e7HwD/mbzXxx5BTbRNoFwhXk9/71T930XqFViHULgZBcd1185CqjbNcyAK8/ljett
AGSIZ4e1LC89fpeWSUFVs96uEZ6V1zR+NWVUsP1xj4BPCQRYPq4bi720oybbjx4Ac6/Qm5pehedU
5DP1LpLppl1m0PqS6xSRHbWuXowgzW2f1x9UoV1L0mvu3Vbi8abhH5lBzH3ILUP70OFwJoR1m1wT
7Ljs9bCNwiWH5NAch3gzKv/SkpRJM9zyt4YoM8XpRCsWr2C/gDoITg2BwV0AqBTTDvdKm8WkXM3e
crYaq1hr/X0YzScdh1mEqILo9f496YikGhlYlNzshnbPKhIHkg3n5fU7k2EN009ct3evR/JUHQYg
mXgDH3pSuuMon5uBwaWWUPI0vy5MIT/pJaCwdVoSW2n8XJSxHzNatU5Ch6BrgNMlmLUvZcJv3ix8
HDcTMEzqzxvwlh1sGO+ceY1msrX0Ka8QzmeacU1ONL2dAVoG3wQkCz3C8Ce+PyR09rqjWnn3zoit
rV9sxbpWqRQbw7vpDu0hOTPjQ/u6AmAh+OWPZ8G5d8qeNZGJdjDwSsaNHGpdz8MZIUJo59U4lsK6
MgW8dXlA6iINKJmRr3998gleP0vwVt7Cl1ovrdoQwoux1IfbOTyyLwXIy9kiPx8oVpoYmg1VKzpx
S6LFpKkigkjr+mQy4tqJHrS51mbW0GkxKlLTSws5bHU9PgAOn+Ur3MieCSMFInWwU+AuS4l3XB0h
5dk3Rn64hPb0Q87dyJ0XgdeY9Zs/HLSjunpX5eIDegBzU1ay+wymcy0wITRLSfmUJmPK255+jmJ+
luH90HncAOSlUddTiwlxpu+qNjhEtaErZ6W0bc+/Nr8EbLAgnqaIIP6E0o4hyTk4ygdhe/ReQGbB
1e4rmWFIyaSTnD9UNW1Scv/FRb36clXm499+XQJLfnKwz/m9M8EQbQdcMhcYBB1/lJQ/4dBATyDP
6XFeoua8EmiNr+avitt7vTg8+LSc1kf7tBh3ZQhqkSXrq4mH0pAThQnh3ezAuLiFRi3mdSYZqAWO
J1mIfv1JScfZHLLOkr2x1AP1sj5oZ925IrpP6mcj5/Nlz5zieXRyX+wypcthgudii7addvu1sFEd
hAk1jPzKAZgzN4Lpt7olxUBRKXhxwqLWaHOT76oPqEK3DBs6prhi3YnErViYl+RIA79zA+I4SVcE
EasqUvM51bRWHIAwCt7kuXX9Sxkxa4xja1x5rZNWWjn3dgOBY8J1PgFBWp3BUNWM+DfDtH0wcvLV
7y3NLLERJwvL4RcLpvnpnrV3qMeukwOXh40uLon+WwiXCri2F88bQ94NNvie+KGgc3uvY23n4X4B
LXbp0M/PrfMEWvclV8x1lZskEznUwnoDXnJr5z6y0wrpDeKPXEyNpHd7CxIbWo/rLH4QjJEicQ6U
GyJwFZkQo6PxavBnY2sl4BUxEUi37AE2AzD7riJd40BXky5uXHn2inicvhb5r0Z84Z4EXkR7XCZL
9IuDEFbTBf5xC2zQSHhzMjQGy0niq3OUczSdaRoEOpkhOJR0lrC2E7UIBDiEoHER61w4LH0g0vER
KyMSSgrpx9QBygEs/RWawcczLCJ+PFvL7KrtJW6Qp+95FGra/BBCE9cfnnD2+eaqEVQG/yV3p4M2
r/vMSnrKdu5ELV18LzYXyHGex3Cax9iE/9kLVFVtvzDV+5QKVD0TbojLRHVgDGdcdSAi2sWmtmm3
VJOmEgTvc2Rcj1JpAS5LcoZ9Yl5oJpnA1jVvZAP1P55oOnJPxRyHkW7WuzNxNvuMYUpbt2zaovbK
PuOEeRVjEhXEgbxNEMXr8uszw5/JzFtgSc+YKW1pUgai7rEtVGZSHudDe24WYFWxGt+OUWDSlgyq
cqK6Feq5gkQudm26pGALhTJqIGH6v/SaT7/HJOTEJWoUAZ+dSuCGs+6UaEnHEFeWhHQJAiY2J452
ReqJFr8OsKubtF/To/4mZYPymudcXjle7L72uD8EFZs2CGUwLQhL2L70QqOErVwRe+YIkvfITlkc
Nr3J4EkmYCN9fVIvMXSdggk7kixL/+8iWPeVIoxyatERz/LMIDYA4Amj1uhXdVefyCHlzzA2S7P1
UDWHPorQBaka+kewqUh48d+St6GPJRK7+J9EM6w6TGk6ndNfNncjSL4FXhIdJrpvnV7BKaeTckf8
iELfymikxV8pIid2b33RX6UI+3g+MvktF2D3zD1FEVnDYv/AAR2Ual624lV7Qf1vjlog/loDtL3g
rK4Zg9I4lE6VpqZIjxeGksTcf7CYiZaZGd1npM5McSPn5dOGiSAKUkr3R7RZMOy6KcJ/pS9f7/UA
ryolPNG/6Rk5+NKdEa+yGgOCeij/knDZw0R5G2vekFKkvC+s/t3EXd96MWlkilKR9uKUsnaiyxKp
+fW4U0JumtQ+roI8zzY+i76+igLDGosU4Dd7SZvXY2gFpSgGD16RUEi0Mn3eMR/v4pvR7F2ogwS5
xx9PL4srwZE4yMDPn1wEoddo0vrfYt8S/1a+Bx6Ibt35dT/pvGSxfpgBx27JHXWQGRYKTESpCSk6
OwmrGRvuZ2eOEf8NB1xOb4T/4ARANz7AJrl92K7GisZC3jdtFpKE6kQlkULDk2jaEG6ek3SC24U7
xaUdDf/9/INBoQEea+y8GSziNygwnI8Y/qEFC+sQwFuQqIZcjXKJ8MsnYbVNP7gYgEu3UQYhk6uM
Fj2JUm/YMcwC/QNWw/D+UAe7wKloHz38LHy4Mt97skn99GbmAUNgOVjGJD5IZqjt/EvYQfVRUzVQ
JoN7pUDRh7mTETI5/lKdN3TaOX2lS7OubDakn8djHdyOdeoxu3DFGm+0pWzWYQjuITqYLoRHuGmW
bOIYvXNgAsm7tRrcpZd+XuMT5b2JapO17s5l1o4I3A5Z3z6gFlZ4MhMiI0fD7RHLtoKueXtKQSRL
tScoZ0bQHlzXGs4hI/uIuXLoPgoyGg5T2eWx9Fc2kXR6yQ+wcIOzwt1UY1tq3w0biwIqZQxSR+2a
avltpCZBLYpmBKjVC4tKclv1me3fGrWr6Y2aBmq51HkSckSIkvk4F4izD93g0RWvRLnJv66CFdi0
ra7X2tjlXlCFCbzkdO4fK0MStCkus0S/oMgGzq2Uxi+NaIX4tT94/B2WDcfEneYexgHr8nr+rngC
AOksD1WH833zXYNTWmNAy0L+vDKK4UQOjQkr9YHBBnmnZT9y9oQswbru0IrDub8HnR1hjPH68sXV
ljv0dbvOm/zLMJ3c0fER6mlMMVGtytuLb9j/NO0f5W4os0wDwRwfxQGxnH9VP5gl5K+dOBIlfHQH
Bvv4+XKa0gr6tGRBk1TLT0gL1yV/aRh2x2b0CaUjClWevuLY32AIUtK3s6nxqXT3kum5IsZCkxfv
Xs19o9BWZ7lMZ2bejovmmRD/meGu8eDofbI1rho7RBIJ+c1danqDlhzPurto04CTBhBlpIKwaLtY
c7Q3by3yo2CO9ZbugweDh7auIIIFhDtSwdwudyV9of2GqLTHWNh7olecxjkCLoO4oB4S12FABwoH
a1IksjW2ska8CGul+AQq4uW6WpJCg4AFo4rtDdILTS2fdELXaQa500L6APowjjXePT78JnxerCOn
6lx85oyxiNtbVJYj+ApOGH0E7tQ1Uf+aSATwlV+K5GmW+0pC/9JEJ1D/IrgGewEh0u+VaJuOtIuX
xUnWsUCH2X4io/lzre/7HFmtCZqohm+4K7Xokj3yWkdmguGA+FmO9Wipp64j43w6zrfwNJQXPnUf
3cDh9S3gu2FO8p4TPCV+/JY+pjk/uAUceqRSpYeDvkbCT1USyY5cqvoMTpDtKz4lJHNUF8jsBLnR
++GyB8UH+NtXV9WvaJgmkOWTszjSsrD8bjo6Srff2xj9lzhriFR+0uPAYE/6FdSQRo3WEQ7BOZaj
LwkoFPkbS07ZOIVoJyMVdQBZPNzqXtCuwIrMBp6e28m/Y8bIQxMQ7kxOPTQAYuEqkt3UV0ZxWYCB
cnsx5SVAOhob7HSneFLTBLEJmmYG5v725POCD8b1qH9v3ZCi2dEysrtl6jvuFORjy75KoeoZx7rf
1ruTUZgy+p8+9U32auV4ctvNQkqrobQD59qGkZBaaC/hToxfL3lqytk0UjjC+GXSXnPc4tjVrHbO
YY9/3pHAKC1JtuNXoyBIz6/xcerUSta02+ExFz0dBqAX3YBgKXdsaooZSMltvPUvLeNDgW6bc5Xe
STw2o8yX4Xza0F0ltytM3XORAHE7tp6bPGOFZnc5mrYPYM5J2Z8wcQ+9ZydmGZqiDGSl33J4XLrb
wO/e7WdEK9sF1A5wmJUwtbKooSoD1wtidUJXMfnrKAkw1c/9UocT1YJdEetUL5xGYpcICCbkO/e6
hKSV8p7ZcHFa+BKYBFDA38m+hxLVTdgGvsZXTNNjPuqTZb0Ld4XDHIsiBL9vJYJGy6vb9kVMxVsZ
Xv6h6s+KQU/+I6ObKlL5CWCajbcin52RUhDY84Fn6+pGsyWg2hd05Egmf05oVsuZBrTRGBf9CpQb
dJBC7BXzrPKo+8Kg18rLvBOHWNi+Ax8BbTDUlIttroAmfqcU/PXJFhZMi9F/IBCJBKc8aDbDpToB
6i2hgVZU0MRA6Xp4PEUTZa/XPbFHu5fpJ9mGqGfHcnda3EqH36BUWP/bwZQ2kMYvit6+S0SBTovp
oOXTaE+PmMZgEbVME3nMvOsN4u5loAWR7gaOA6n0iB0KrO7uSy8oQRsyhm7ZBgaDWONJY6TcPQYu
MZ1g9Wyuj665SKMI6dPRwda1hGmTSjzr1VszlDJixBU6aUDfOtTGBB4aME1yl+PqC9NXFTlfi5am
KgHPrFqq8iXP+ItSAXhHLXE+Fo/zt+MhJMT4pu48rrusdaoH0SmYBE80NI3YJFngf/mg6CrOFAn2
nw68gm0TxXX7SFrPx7IDWAcO34PvfJKLH5mY/IUe/uOTGSX0WG4reG3K095zKV3PlDgBOhs2eNeP
I9FPRmYFvtyYwe7zT13Xr+/K3g664MP7bkFOXp8VD4YsxXLEm8sA1bHCOHc9NP4qJFBCpBiVb0sP
qBmzZ1SpzWTK4cTs8EN8JsT3at2YLPJboDg781/FY/Fufg+EusRUWgtYqfWfpHUJyFvsia7ih1K+
+dZinKHe4UdfjzNkwVfJtleGA+hZLAiChAkSUU5SBlRZCv9+fM662v2+LoXDk4K8HUkt6UcR8gLc
2VoBgNEwWDaKVvY/gsg5NsBZlDqPkv1pfj5CvIbFadIFMTenVfLLsCevN9jNXugFH7kDHr4H8HbT
fyWasSQHYRqphX06CAMYNIrg7vkjZaT/EgnrDrA+S440Bd/zIgEgMZWC5LEQGwmlkVys7AeT78zQ
DWOpVupPk0cQEtufqvUon4Wg8cmegYfeOJmumA9qSPZdI6r+9S/91AOYu62o99DpZynWHKrlJ9Ed
IKrTF0Ak0ywe2a2ON0ffGWJIDPeDnNVWXsM1yRu2FZsb8rx/A83AESPEj0/a8S1MHNcfgnMtWDWf
TgcTamm3qyy1MsFOnu6Q+Y3E3Nj06bdbRI3X04/SE4T76MQKx9J0RF9vGCbguZV8oG/x8sxkmYxl
XAe0ydvD81iQf7C2ABSC/N+5FgJK9HKK+b3sgAkGiW6FqD/ovvGMEkxe/r8XWICko90S2aeM+xYt
gGO//Hvc/7ADSNgx8e8hyooDIyFZKNScwrI06neIrslCyNUcodMF4lRP9CQE6EA5c5lAi7ECZhPy
PMfXeQUizCsbKTv0f1CX9aZ15BS92kxv33jgx/Rv6EBCf3gXOmKbRwRdf3MqaYNYdCLiE5xCxkvK
aXBT9vL4DIgCPWqG6x0ci0Qwr/zdI9sqDB1DxwyCAv7vNVTyuo2zv+0QKo3/8ul1dK2t9TI9f3b+
ca3OxQhgJ2213agS7O5+szusxvFOlIdcxQvMpn/AdKD9W6nVh9WPm8F0atZwdSC9UMPFHFPfTtdc
5jBJFdnW4VjL2dlciUWUy+fH+CNUozc80jM/W8LxM6UiTVu7aDPd0Xv4mgyCkH6PzmvotgP1atwc
avRSreI3/3Sdh2Svl07p0MJCuCg4p6uLzlwYbuO4xbthcCrxTJvjiBDnfu07H1Mw7virhTwUhwie
Kox69bvhsT39RKr+vfEZIc5qldPwnEUlLC090FaRP22xrQudwJf2UOy+1xm3y/tziwZPPj38JAMC
KxHmVBWl9yzOeytvnZxwbbqQfNg76fziI8GE1u80JE/hb41XiV/AEOFKhjMFr9sGCmFdHEh6WciC
/xroLOHiqVbnatzHOcjuOCaKgROw4G4V5dYu64x6BcqAooUaNxexfZGZBIUgsg+L2t33kxMKfGZz
lPVXMeNEAs196WWgnh5kxE+NhTLRZ/CNQ3v/lfMnTDvVcYBUqAk8TF2SGYpGBQrhCmrOJ8bOKnp8
OHVsubqwmVaT3s2OjB8A8cvFzHD2VLUR/iqnmrcDxD+tLAXAmNeKjScrPYtJbMgwE4Mx8LFOtwYo
DBD9cK+D6ok1OgLfFwkNrrw092XgR/e/yeGwFtm/VD/0jDWoh8sVMu6EMoOKIkdToQzl0FTqP6to
tMxeQb6/5WpWLiokL+eZb6zLelXCZwMshonpiXPU4Tb7KdvGgIZT9pSYzDrvEgh8ZAKuBCHyvgx4
uiUZ3UMIuv+e6E5Mn6vgKm2BslEplUHTDF9QMsLGuwleT57HfOSzAeb1iytcg3Fx2v5LMgO5u2Wm
Z9ca6fmVzWgoTv5/yadQqzqYDzJgYMwKUhSPWQETbELNX+qVby98ADB0kyv3toxN7tubm8HhC29f
dTX0zYHOThLkqWFLDwZogu7JdgNyVf979gumtxfQTHhWmkBh8lZfFm/hveX+ytsMkZHtpXbrfzre
YOV7TvUGDBC4Mup1fnS82E9cqLIJs1j2BZYkDblUDOTZOHOZCViJERKpqCrd1uXZQjXlLZLIzkfi
QCkDJHO1nj+Fhd/yskMZRi4kdLxX2IHa8Nu+V1Otb+65PK8EZwKc3nbi3BVEbLXQa4o38kCTv6Uf
bZ1T+AEM2yDm2VVZ0Q9C+gXVBS2aWznbg3MN6E4aYvT67LPzdg2gQII27+kKaQNq+uXXqTTbjZBy
Rzr/QVCRfIQ7e70g2vUUG+K2+/dUvGtRGvlQUM+PCUTOUILncU58QuEF2wUwZ2cvzM4eUpcJ273K
UELp1xSbULZoaPAmVPfrfbS1yTv5O+RrJNzDSLtiHODr+7xbsjYSYmyZxnGhmTJjUp6yLiwKHPwM
6eUBRgV3qMDc/UmXacomIAxNqowDWaUbSPdmGxJmVCJc/BE5SO9IwNGPfv84F1JUyL9N8ZlQT+jM
vne7zsmf7A1CMkTOrqPJ54LbkaOCAEE3mD5sUS6pbj506Yiz8UngCZ7XFTRvZG5yZbtwiUMz9RFp
5F/K5WyooTD/0pDMlEzfd4iQQ3Te6fX5G0H8aqC5adP9BxH3qeHDxecI8xx4oXzXQvUw4c2smlCj
RqKsJfPpM8tP2KT5vryzmVTJYQYXTl3Iz82Gpuq7efxfCVDAkmi4hOzVUm2TTdPQJmTJXBVJg4pI
fbiSUnpz19lWlnEnvMUU6gFIAnT1MdbFQgp2N38/1rRTNglMBR5FaouGJDdxSPVRHXkGUUwGC1se
moQBLdYDb3TFDDfH9m+7tQjObjDACdF3LlEI8pzP3Z+fYuqcTK/rKp8Tp8P/SxB7wWVH7Mp8UEW4
DRFbSggXmlVLUEFypwy5O9ezAUBsn4hQY3aZSNvg9ZoFHpABcy8sjAmJb4QqZ5QHuhi3mpEMj9dk
sXZy8/UQQ4ENg6QEISZ8I39d6VWgrdIsoYzZ1XsyteSi30ThHzK8ALIL2QrJQph7Tz+/40QVJtWp
rQ7ABiQxLeg96CKOSbvQAu0IMa+q+xIMvXTRfJNhejaJ2q+iwdXakX7KNMQL7mbJY1KtPTlCKbbC
E7uTl+UogbBemrdEKiLgkAHZgKjDv0CFRbvCDJi2LyGppxYeX4/PIvU+g+2vWWCyOgkvwTtiaT9g
HB1/BSKYA0qFNIVsJaLpGtpqlqRk6z6VXJs2f4pF8Us+LIvF3KD5fHCpvk7wNA0Xvrudulxbdw76
3vFYyk3wsunArV5tSkK8opmKfkSLSeTU+pX1PNTG9He4xVZr86JcanNObLTFsmglAQRLPAnpNWdU
TloH9FghT2Km2q0hl5PIAUuxtV4M0sgFf0W/2TVuy31QvwmQ3tJRZPDZobW601JmoRKlIeRUsL5u
IRN4w/1oWttPUSpdqFNkRGPDkPgRxz7kg0JRY+eyEnLovvX5aQ8mkjd1xBniJT4TB9MnB47zUHMG
MgU2nxfaYJOzR93DkhGAX4dLYH4c3MsAN/KzdAvY3WrRtUH3+RAcBBc3CZlFnhfgjkiGL8s3+O7Y
GvbtOvrEG8uy4ScILIxR1pO3F0ddqBGps4V8NFfSeypRR4Lpp7WrPikm/DK13x3XFbR3nuUZOep5
I5egI+U63u7mx6pyGz3Y3Ke2jY2kME6vxi3h0e/r7fybsNCtALF02Gx/uYlDlluu2cBPuRYtnZVx
ubMXXpmBbwDWwrGzOPXknzyCH+VkGRPp2lHTxA7zsvu1288X474zqJg3vzxlqmldsP/15d8i3Tgp
IpUil7r1H80fWrSDysU8MjJ6RRzexNCy854QDgx6w99bThw/9XYiOrR6YMRyr4coyqkKC/2uR9mJ
UoKM55fAQ47Vyn10CzFVyFL9MwYlq+g3663lH8DxsdOpp0RfpANuIZmzhd/R0ZekNmKaJi1BHWX4
jv0q0ZHDC84fv2gxevbntZbyAsbkb3ncBPwtMUbxJ7IMHqsSmmobHc7MrpsCOLpJeNjQcWV0qshK
xKYyg6xguwSGE7ZUyL6Lfn58Db/fyahDwT7TKc2079tKmoO4LIU9Gich9sYlK6YBat2TEgjGe7SH
GNkOuluOYh87cHvO9MYIL+x3T9GNS7QsjmP5avMKrtmMZW2jt5wmVXbD3S64q43MtMSkUFlTwZGL
YTecpNe7iVQwP1eDUvmluVo5BEgM7OJ5IeoyBDIgqW4njzcEUHHHEryHUI6jncUKCnVPoBgfxRpM
XFG1mjiML/+uDSJSjaEE0n9BnYOSsBAOCk+1HdP2BJEHkAVn0wknBsE7Wf7JrlmHCpAzWbtad/4h
M4RSIGmMSzDvAiDZQWiqoKi2Td18GcvL0ns2fO6mmJlj95h4WhCsb8tYfTxTNSSMiABDA8qXLzXK
yTV//NuhbhLLYEfyiN/RjuEFYvW+4wNgV3Bho/vLA0/RikmQ3oSwX5QxOcIipKV6sNiHnTBpJ3Lj
81+YIvNk9YkSJ2UAsiSsxQSmNeBKwlAp8yNvs263mSdQN/+hLmWlm98XKaU+CPiB6CP49AF5BnI6
ub8eApwEaZXldDmua1Fr/raDKGYw3t0ItAzpewpr0S9sqPhFgJqTmiBrZBmQCIkJtHAHNFsnaox+
mPanheERVGOTi+W9swQZflKLFZ6Azop3pBstsCZU0ni4UM1M7QW5mYAt6YNZEFSoCnsVobzez1J6
cHktHnKJpHSRsS6NihDBKhhhdbOvaeZAvVRM1lpp4CzXDyaCQn0oBT6n9qnGRB53lhSvvOlM4iCn
vFbJkAFpnvNpfGuxUfAg3/BNVS7FJh4D2DOpiDIkIOPpK9C1OIfOFBALM0X5FWMNRw6nmA6SybHl
4eIgI22o3Xnw1PVqkXg+XU+KKaZWBy87XVEVSqHfn2HLXv/Qi+MJ64vUQEfFmpqsSZGPKlf+H2YN
QSCm608I4ocnZvs+0TLU+5S/Obug8tdBsrUbtb/P+DmHDx17iHt7egL13lZtR918o0iTaAeON+0C
VZEF9/D0e43VRUQHzMovAxd7L22j6XR2+jKTNOuDj+myvMTepmfz9s+OhIN+LwYH4jWWglMpM3BD
On+dtNyJUSTZrAvvEC6FPH22TX2MKQcqfl7yVjcWSmylrSQZe434R2LwGIoBk6iD9+a+Baaaeebr
hVDvXNoPl4pxvpn+iM5t7HZ8KG3uEGdg/RXD3Z+MwawnZ0mDk9XLrYxa4/8jjuySfRzT2h4jvPj3
yQUs1EKpu2ArLkRYmHmud2gmsuLwXZdvbJUR57W/PDY9uJkepfgDxQd5K7rD2Ie60/PDSlN7u9Hj
07z/INwBTMyOrwa6+6ikcWiOl32ZKQna+AmnrZP25nZEi6c/8uULPDUCWatIb0eA/gdRqgrTVu2K
AVo5zMDBsE0uOo7za0FcaEVJfqFaipy9dnYUgEblWbxgqytMj7kXozGSGy8QOpXYAr1AX+RSFXHm
+fdXALA0ijL/+qglkTZpDehPfl9S+n8RgDoQI1eYCx6i10Elam1IiN620U9DBcVo2xPXHGAtM1Yi
A35Tf2SEcgHEq7+Mv8+PQ7eUCl5rlChEc5TMkjCa6ZsLU1Hb0pyXwPf/2D90vrCIhjFc/oXAyKtC
mDu6/2vd3ulmcFioxyHlOcB5VWilZ+ujFA4F6R5LBb2xDhRlR2lEHgyTRgti+z9W0PlKMJk35i3x
q4TcdZM6RXYlNC0La11WBTjKDlHiNekJyGzRrNZxzV5Pn5GZQOjcM7ggFsq/wljIUZdtlClYl+qx
cjQiA2w1qr9pyqzTkuF/XkHh/B8xFsgFEL6q+RndYOPOtxg94xf0ZIemzqcXWqKS4UIwVI5uqKR5
MdW0UD/8B4M8TM3Nlda3fz4RU5qJqPv5+ZuirhMI/lHZgBpiqUd5kizKDadBuS2xdL0X0b56hAjI
msgdY81ecNutTX1mDPmo6FX+dK26YyxDqso23+N709fxGwNhxXoGV8Mw/P3QB5SFb0JtICCsPrFQ
HuGer9tw/d3ijO06nwTsvT/gOmswS0xPzA1JP9vBIZ8QsN1z5tOIyrXWFKSFkiaz2v2G8WcRAfbh
HJbl12MQCVdINtMgnlCyEJUeEvcGo9p0vcA6h5b6x62vgwPaM+dnsmMPkNUtNRjvJpjwGiTCyTU7
sxDgEjgIZNVOsvQn45yxBOpn1NJSK/lz+Un7MVeFoHiGINb1jcS7eIkPxh3GM/QAew0w4kJ0FH0U
yQ7yzYH2H7MMYxXsRIXwqFx9rfESWPwYX6zQQLVONO/fGmJzNNfSTG/+EMCKhaHzK7Z6AHjSi98/
DmKP0ghQgnk81prZXclqtpY1LY2eCSvIAJN1zlXb9H4rY2CxygTx3FE/1fN3kE23HeShpdwk0ayy
49RdBcqT1lORpA5fmojhMdz2/15ift3furR3KWbfHaK3jaB9lcySfKUjmVMoFriQ1pFjlnESgGJ+
j3zywUSpZDQO6ADhI2P/yjbTmV7LEBv7GR4wziWwsxNH25xBNB2CWceaMKfSmo/HrjVFu5h9CEoB
7BnUWI/IGDMmRlxXotCDcbQv4WwWjPRVz2vLS2CW5wU2ecnr2DQhiUiGtxjeVacpZmgh9mUgzVsj
rjHai36dVZcM71FuZmZrMzo85I/k6+qPqA6MCzKY8pjBvHllM5E4eqwpMUVT78Weuaqvt89jRWkJ
OJVxrqqsO/w/xMDI4wQ4Goc/DL6A8339jr0axtxbc0ZyMMrCU4B1ukvYPgCszgi6zU4VZ6kjuG/S
jTDdPFcl9snqG36VJeDhHYX2M11t94zoGWDW3jEHd584lyRd8WkWkV6i69PTlNB0stLlYKzVIGQ1
mKQodtnbQo9BNoQXhtfOYNXpq5wMy92NoqzGelW+stSMdxVWcQwbzhXB+YUmkcHsZpzQ9kIIUnHX
2l/+1a56gEbMS364BShYA56VROPfq6XUI2TlPuUZA8a1dIhYzE7rGqD0fMIS++c8jMVo7W0omjeF
khuvr+SCg8DnTDIXthVzFgHcEP3ex2OiC97APX/R8ePWVJa6LrkKQ8m2CoI5CscgZ5C4b4GUrUOA
itI7RbYTzOAZlKqXJx/QgVhXW+bIs5/nCOUVgn4BjSMp/MLJhgROJ+DvDglceT+aVxAV8D1ejcdt
D/4FGb/HVO8JENLCLru5Mz/dcZ/IUKYf4fu8Mki1/RosrL0PVbxhDRqonpgrbImskvZP9STa2Ojg
9mcZyXWDfGyYzUSpdMTDS6zuqZZ/grdTeQEYSX9dNuFcyKttTSqMEYmtArmraP+A+dMdHIPzCg/+
2ZePq194eyYKBjoit28WEq/WicF995Ua6n5N47oRROflwIldMYFfVp/LMPw2+ikp/to30gaBNI24
+1l+JOYVHD2jtWbg0Dwfvzc+TXh+aR5vnRx14DiiXWhO1zo4eB/xiEfNIBjqicrRG38+T1Z8U+FH
2KHXTaCYVLnAI5ezPbDBdpmoiBK9uEPM57T1gQVfR2iNpjaCZmLGqNpzO8Z9hJNPl+/aaHLaeOoP
6kchH/f2DmdLpwkWjiL32I95ah5fkK6OYkdDIkuxinws1ltu/tQi7iOSY0zXpyP6PLDXSfQaWQO2
4axbbU7NQWI0OBj+9ReZHbkApTPJruH54g9IystltptXk2E/+YUIQi/7L0y/l6r1a54x9IpuLNvv
KvbMx+wvBlnmEwUGDGUUxRryKOBtwXdXtmgaWJgOggqD+J//LoFVncz45oaaOpYgqgVGTwN0TlkK
kihHxT22yC2wOBQjoV8x8E9D6JGmBeKw71H21jbXfAqtLpGwbMpU+sS4LqsxkQLc5X0GqRXzZ5y5
ii/4CkYCeoNUcmed7nBbD9AiuNMxJPuPyruw3pNBXpMB3l4n1SKd7+AFr7knfqyCQwb3vyT8dUG6
CPpkoMeIIBZCAc0oRZzMv/v+MozEIMrMoBv4DuDJ0UxGYvmSn8Cy5sYpVMy0brwf89Gy0SkWKE06
ww4xuh5yHwoaoXsNaHK4vjkMO/RNxnLgICk+x8Jh47YkwZaZyOSWQ0gZwN9XCnE84Ak/tnhoQtw7
PWSzD8L2tnl59XpxrCT8luIZBnkxq5w1YxWifRbsVwb8e7jzc8E5k663XIZ2dO1x4qshTGeTG1Oo
ncCpXeEQVsZQNlfFpSX5Fnx4Z1DbgDGHttHfl1aKPjt82nSJbM5ygV/cRXTHzR+bzZB6NlwQjkpi
cAuEIx9Jc9YANE7Rx19+e1HFnMeWhFzQcMIxKwarrHooaJYv9tmijZ6XvdWUCiGyNU1tNcnzwyAD
8Bl0NknvOK0D/jM2ziXehYqHo/doStxEowITCRztloG6OVVnsSwjUXoV8xmOFs9+mNgH9SDTOV24
QImfTirIkDZcHYbWUG88gzZtXuFBDLM3Ne7wVDt37ZIXx3LzxJx3/JOvKRUYMPqZ46bdM7lm44pe
v1qqs4OZEDFkVJyb2YX7ejue1vQwuBTnwnmZ5nWKd8NX6NoJhZn/Kh7D+wb2eA6lbHUnN2WroPiF
IK4khlnM8d9rkwUX7QE15PosFxM7tg3EIqFOU2b5ez14NX3JSv4HiuIHPLhacHWC0l4AdVQzKtqO
GOZwJwNftFSrieyd6NlfavpAROqHDacCShGWAqKOmY1CVl39fYjEr2+21kvlFbwiSLw0q9XC8rRa
TM2gd2EOMS74SIxiu0ZnfhBOODKk8EVzDpQhgsm7Thq79PmSJ6UC7IRJujOs6cf/NVZcw5msylIE
QGK7+jNw6IPBxgAlABTUjrq5+sXQ6kwT9y0xrvaKwmMHdFtvlKoFK59IyZzeyfh12AGKwXw89fF3
X6v1ZobZzHtJA3iU0xhIhs/SKRKFPmMjckvJNPRLefldLGfVcqRT0Paldk5wnZAsGKj/K1YWrJdW
um5Ja8Yz+MWn8brh/5yK36b4I1KPPGKZEWldWMBNGa86reM3HStCDl4pKIx1QLHG+xOS79WvnByz
x1G8gBhTGfS+GxgCEXQf4IKLM5z8YsRfmVYtITsel1pVYdl5KJNBAQNHwRCCnEnmp2ImBUm1GBGu
iama19/yWiLE0QxYwmIxzzAZZO8W6j5ptmEHizqIkb5yUexyhghXze7DPEmOS/vOEZI1wkKYacwT
OJerBiuyxf9aII5RLreimXRrTQH3kUkuovQ9oVIUFUsIkVPDXiDyArSMpjjrpLAuoJbjfMbeAc4G
khGMjuIniYjEdIqMG9q7UhmksP6rgsKKbz8UWnwN+I94SoEWQcKtTtDe49byUVhIDcWQ2bvaN7wU
UPx68Tit0PbbcOLBXeho4heYSDcPEh2NT/3EJDQbhSOM1Q7ax8V1qDCjHoewJQ1heMMLWrPtejir
aZ/SsLRhRISvoHQ6tm64ORrD2Q2SQBMiY4/aZg93FwGtXixW5WLN68eBj4Lk271H1sSoletr4jKJ
2yX7SqEP6dY6oyhEB1he02sgaTEmyqEA20ljG5XTsJSYpLOs9PoTj72UXrOq66E/y8Mk3afY418Q
HeVzscm1L63v6cIBkMPHdOOXK5macvK6XGTSgR+SL/wds5/IKwHuP5iEQZJTbsCi5S5u1SxNpwKT
OinePzGKv+D9zPbPn8/OpnLJKA/NZDoVoL7vq+YpqeJt4iBrnF+rP3nTTDW5PF2wjUbDtLZQT8ZI
Vk/yYbTU0Gjo4Pn7K8qWUiqj1ZpljkrZQPUpoP9kujzd2fnDfSm77qLvQxwT16ibe4YvyZGOcl3g
Po+4+TNbjoA+JlWSrqf4d6T8821m+NN4rM7+ZaSlCWkbf91TO6uhpKpsk5V++39IMYwjS6IVVTWW
EW4K6XXoUFjASqYfqvvPUasJyKlQQTxsHcB9SJ9krEq2yv3f2P1uHuPUOu4T2kay0JC5SqgMKmGu
PLi7UKT45A30MBp3Vk5ETqhcg+wh+DGbXSPs/Kl0U3bWGkGO38X6fooqcAuVtfMXo8NGnlvlhK4c
qs3L68PEGqUONtqZ3NTnqlCE4KIHqu0Cj62XOWX57APBQ+SovG/3lqjjAACgC8XSwHgp4ZN3TYtH
vRD3C6DBNeZGoWBVJgcOUMwvaqK2tjQLJIKb3gaBUy69pV3ay/RXLKxo+4CtqLR1Wgn+HX1dX26j
GHwhZNOWG7xuEJK1n6n75RqIzH3yNt2etZo0jRwbRM4pZfb9hxlEHtD0IasYFi2v3EUTwxJH8ILP
ZnOeAgMiICvo4lPVD0qTwCLN4EoHgq3jcDeRD6IJtW3EmKsK7Tw2aS9lDxyxLY2crXGeYryJVakU
YTHM6emb9v21PWCzg75hX9RMoSMPWatrJXxAJFVkYWN5zDcmOWAXA7CNqwY8eW374rvNMsxDEBrz
gL+qSA5YrxR5OYAZTsttz0KE+wu6HQhe6uBAKbBkmkEqcfUhJyf4Za32uixq/XITNhVb1K3UFmAq
BLUGqgu7VbZu77WuId4QQNvF7hpOQA+mD+egehpE/N8B1cwONVByKPA2mH5ZtGJGiegSMhhICMQw
HnuHi0s7fZHpz5OZH0CPVtnhYmyiprBfVqbsYUCHFgHimGKjbSx++vw24kRAlsM4FR74yENTFTgH
2U8D3sr+5qooxAfDemXW2EBOU5Ik6Aetrv9VFjtONRG8/FGtpANvUmIKU5yG8FgM8jriolS0kkPu
9W/XioCAg683LZI4ahgr3Xuwc33q3b9cR+JJzbk11ovaOJlflJ16S2qUXDA/DjzaLcY/DFsnvB3l
idMiffM5IrucnoB8DAacUv/pQPgN6J4txZE6s+M71iepQbMxiE0svl3o5eG3ndpknd0ATcGgvJPl
rFQH9ZTntXHBHU2yGpdNapPJ2j81a7IjHQyU+CUIiKjciFR7M5KycE/mKQHj3OGzKMbxfSzo2zDN
Oik+OdzO7N1qBjvPdsLwVqpKkgK/a6yZA/uz3mpjhNG62EcTAl9BgwIbG9HEvajHNGNPf/bpCP9i
ysTMa0GgcvdCRxw7W/7rG3241lw/Do5Jo64kvfE0EttV5vHJy+TyQtrX4Gg5n6ewD6eWCh0vCTS4
ktVxpua7lu5J74Z0JLD57l8K6KwAdjqmXAQzfRwZug4ILBDfdvjtaA0NMC3HCfHSFSkFsSv3ldsG
E+07txKB3lP/Apz0Y9+i4WXNkWS7YfJv4N9uci3/RjWccw7e1dBWTHNh6H6JKo1vn5N7pt1CkIp0
EnTNp5aSwjo1RO7hrFqjmys9PAwTuwRzWbKQQBXa96KSstdQZ3SpiYVSNoAAmY63IKPw9QhKUIUY
nia4fzfzWLZeN9orNROAkOl1wUsxcWHQ2bfyntIMRAOsej005EclV7jqjyxeHOAx4sBiNR2lVwL0
6FfcPlL89Ghz10P8HlyF8wL9ogf61basuxPv/eytnTA23r/JZh5I6SpVVfOhactYSX4wC5nmDmGq
FHeS20/ozsWWzye9+Tj9POckyo1myGM9uQs4TLX6qABotOkB4I794dYQlbmWhpoISlnQWn4Uj7hm
rEJhQBqKiiSgE2qEwTrssrsU/tQTbLLDk6tt4celI5NjqKrhOVFXCZjGmBpIdjX+L6IRxQ73Iy2t
ccDneTadN3R3kk3FXJl9nLTRgQWBwBeYuVlKizVKh/+ue/TV3826n3ek1t5vvCZNO0xw0R5yhSeh
GT7S+adFx/Pf1z0ayJtXQnFImU4d9tWaoHAcqD09SrO3gEpiALhJE1wGIUMVh5R/SQC44FD9t9fn
nT92XFI4XZbZr5U0lExcerhtUtX1sTZZDFiV/GGEQnXkULCUNLxAYf0auGXSJ/o+IyAlIerwo64v
78Jdq0IDCGMO0I8X1YcSghSmU2mTcj6nfqYC3SrWwL6THLxJks/f0owOd/hYYDkt904eRSOBxOb2
pPm3hVgR6072YnXpz9CDFi3IYm+JeId2FeXbDC7OiNv/IxKjoalwxWMmymy7jJUMsrnh2rvDjURr
+kzkJ47uJsXTqQJTbE+EKTMvA6qNYphT/Sy9rr55WQu5vUyZnC6XCbblGz3mVy8jTtN6dgADWz8B
c3dd7ysIAraKxtxEFXCrDAuHuAQNelVut32BC1Jdo67p9epVlGKBoecuDzwkP//QSLGDLdEInTtB
9kEB+DOaGlc+I1yb3lbXUenOjcHz0M0MkDT/IRrEYgsfeWIFL81ebGe7qxCeVJXqV1rAbploPJZr
dAHR+HJWP/hug+Yy0coCN8Q5ZI6wKRegCgdFUinGE8lpWOtPePJ9RQ5NUnXzvw5a9DHoCynkyGkh
EesEFrrr0qqYkhMRgYOlFPW377OOylz+rQ9CpmjfRrul3ENrxBbuG8ISO0Qkg7PlhIH1jnKIstV3
Pr00Gr98/RptcMoY2ffLrRMl/QxS44UC0ij8E5RzHeY6m3gkf38XWDBtYoZGqfJ0vUfa+KELmBbI
ehOojX7VfLAsfS6Xysbni7gdVfDhuV4yyT2amw+JOustqiMvOEAorkU5PIN5czeuBPHqfrv28V/e
h75ioQbO95mqqeN+FPtJuuTOqFes+7WRx6WmmrzSgpN1rS4zBIJmD42iCf8ba8SST/aCTJm/P/Jp
VvF/H51DSWsYpujzUYd2L1uKCiau//E1yA7CBYQDhzcHKCeudpiKSxeJqmtCH8ZOd6uOtu3ztQWk
2K5ozixi3I8z558rmfs4OD2lO0JeL/qOw1RzNowizfg8d7UQhqWBMeqK7BkBzNW2qegLBp75oE4d
QZh4TNxfvlbHgGuC+z6qOBXHz61dL/5vYFzJ9loj9I7WAa86yMDiK3nyHgrqcZU/aL7lO7cRTwhH
7+GEYhID68sNO19pr/aPGSpCRnskOK6ljGpDV3y/KdrFgNf+W4NsreoRoclvGwYJOBCCWR6ou9jO
5If1Ri0RhWQtJsdcoKFrXMxqBs2nlwJkDqxbk4KwSTqy+qnaxyLiwCma/rCsqRxbFMXlfGXcNwWH
WfDZWZKZ5FgiDrYc5zNVuQoOQyNaZV6xTEHsh6IPLugSIOzowmTjxUmubUYP+28F44MtFw0eVoOC
93cjdBhFuTV8Vkfmcq/MmlgvsvWYTT47xXF+T7d9shhKbsijIIfoKGY+bUssNVYWYQx3C8IcBWHB
8ZZsmVexsbaw6U7IYSECEtPXi4BZdTLlX2s2ejWwD2r8tf3gINEZadTAWKGZ52NgXVQUvgr65wBF
F/TVktfXobXOwcrOIB1+8VwvZQSua/U4SQZgGRwJV0x9RmfZtCVOzVLUtJqKYzWLOR25xATAhkll
SGVZ8nJ1BPja7jC/dsI+dua8Phao+XTh8HTYy5Fe574JRqtJLE0sYpjUrJY0qQILd8mZAygxFBbJ
jFhiMZNejWou/FVVZ9O12uYStZXHhF3LFkMjc/bGK0JU0STtmIxDU/ddOY9fgtCDbs6EQ3/pMlJs
VSATl6HpCfV5A/okOYbwYo7GntXEQUrsmXhj6KpUoEs41HxStBNPbUWWxYlblsSmh2PViYMFE4+6
2cNklsgZ9NPmXyFOANC0OthAZ17zT44leVPVtLO4jvsoXE4LPIYbUAnSniMhpkC+n2jMMvR/KKKv
giI5anWkbBS96ola6akhQURczLXGXSunFf2ks997o/j00DA95LLIpEB86g4//akk5eZSLUccn2lp
07KY3okU1m1dL5zXAReNJF0D5t5ofP5z0sLX4mINw9KRtBNEqypFS3L7J0iQqTDPiDRD3hQj6BfR
1R3ZR5jOHvNRQRTZpXqiaQxfCsCPlDRAPbQD9vr1NxJyj82PoprkCjZ8v5LA6l/eeton4NWSdRU8
lD6ya7yYJaE/b4mVkrqf6HzTJjLKFZNvsR249I5+t1+UuDK/9DZnd8bwQ//ALsY3kdiXDFS9TmoM
HnBDUt0w1JZordXUVqZIRuz/AIQk1e4HIGzaa7X5oavLUwn0YEV4WMrmPKvI5FLPMrovZcu6pk1u
Vjl2sMYoJiUbp/tK8eQM/bL/ldCMRwDi6Xuae1lWsg42bFQMf6HJhfFgIn+HnlVADWTDle1TkjyN
Vv464wlMVV3ORXZClZAgDJdxLZE9L5J9+dbcpUkjrojuHSRfvU7h3atNYHzeyicoIKEIZAlWxj1m
rRxYBXK/RYRS98qw8w75orQIN7gIGvyc6o6JVAimsrMsk0fy0xKQ31v8/OOPugAJQygxMcdcTHDB
04JWJ8P026Gyq8lXQvO1ISuJ47N9rVoy1tam5KSmC/AF5NJkeOXBh8oRMbCgvHWQOLkGamu8H3TN
YGysu+Q5yY9jRV66T/VE2cbkixNxGtkbG8ZoW/2k1CjtoYQEj19ByFrLro8p15BJjeTM9hzJFd/D
V3ztCyzGjOU2zMu+ZhXDi3gK6ItRfDHXioI7sd+yyjIIBFqPwr4ieV8xt7kRTk5iSTwLcsUd4Ho9
yR8nA1Ou15EyPMqSLss5K+PtU9WuifUMZup7NBvHEaVtkwx9fjlHvtha/En3+xSlOBxpvu5OosuF
zlPTx0q33vhmFUr3C/6Ak5IUDKciWjD3ikY+hx+3RqtmhvJsecXdhmeshgmDVK1B5C9zMX0hgMAC
vOWsY+MmE6QW39l7dpwOBFNweP1BIZK9Th2ocLcr7l1/Uwf5gjtzEN9bJPTmbinFxwaT/X3PHsWb
xQWG7eiiqKOf65T+eT+ZoJZQ4EDEPkIjosDIRkXBZED1yHj4uxs7BMzmJ65M+jmHyn37oBasI5gR
ED+zXQvRSpfY612cPxpEg6Uz+yrJ7fsoq0h2luq45royKAViy27e2arwHjk9KAPcETeWhrllD1ya
hcg/+QDAC9jNJuySq3l6cPJPrR3iqB5EtSgq0meb0x9UXaTBJflCNf56Pd42cxWqYeZAu3f1K7mw
QhvQl/JcERFCN4/IwZNFsx3P98S2XoeqwAP9+xHCB6uQ92/OBNKK7NIDLDjTaU+UYjBWSxl9aLCq
SOS3B+tZ+AkvG3tzcx12VHGlcWd4SBMhhPPUOgb+jPx3Pmt3L1Wwph+qSLhvfZq/jcRnm0tAhtEL
OgYF5Opr7NvXmXqvxwRo4VLqi8Vyo/v6gbySyppVdN8YCFwFb8LwSVxxR9wmkK1n3goBx6qdgOJp
ZsJZwY6wVdIR1e9knkf7WWVjzd2jCb1Bo9gbrgUpyPtBktjFRkwz1RjYRhiz2HBouT8g/atmuMzy
wM2xWuDOkmaYy4MtQctPABDR5+Uh5GohiWirY+9l7DkNNfIl+XiDpB8iO3YiIAChOR8QxpXAn4Ga
NBiUrPyhzSkyDPRQ0t0nyMp0sIE6A/Jcxgg7YsOL3EzKsRXWeyI7g2LqLsfLS6avkVh1Td9t/3kk
A5aiC3Or1I7ND86LaDyXJvdzu1RlPQfsjZnjw+a5va0rPBkH+0Z/kJX/mPr7taN3wMaWa4N6PZsd
eEcstcYe9Ci3/oaj7srnL9dm67zkqf7w0lnANRtEbr7wgHkgLEONsOwk6zm3XuyVfLC9w0/75oTE
fS/CAIajeIc2cCi7mGP3BBxfhX5etKlNRcnSP95tiQXQ5djaJCjFUIRuu7FbOTkCjwe0ftGXr//2
YLzCaNqqnQ2T5suJtQFumhbYF4muw99Cpo9Po2tA5r0DwBmOvTtuIuopgkXj2D4l8sThoDvKwlEO
yAK+D7KE/iR9i06KNaaSjNfQfk+Vrueu6NGQzsjl0Q+k60eWBP7iR+nQ6bMalPBiqMkW5LbDU790
gnxC1INeyNSinVQEdh6FRa3S2DWxAP5gtJU9vK0Uz+ZCFYWErbqkoG5hDDZ3r7XqIPEqnopN1vPG
us2AeQD5oMc2+obEEcyEJX/4XX1W7vqP2xlBnmJnYEmY7YHm8aUIcWS4VVC5PcovlN83bfvFDr1b
KgnGKgPmx1x6EHPgYOofcBN/hduRl5W/ZZdoqCLBR+90NmhuNpyXwbYAtaBpsgS7GJBowA5cJ+ef
1tLg6O0PgvdxtEG9qqw7TXstgIL2KpANnmuZBNeBbrcUnANyOrABe/36AMI+HH8vFosfzPAtCyLM
tgAq6nb/HT8vr45Aw+qF4WNUZlSdmIf71gqGMcchEhRTQCBFsvojKjMfd0/QfnZnVrKqQ40NeOYk
wQPwhkb/bPxqQiKPRQQyIXXOjQWSpAAlTTDOuOEYUA4hoRpCMFiOfcnnFIJuOxn8NYQtKLv3ANZn
x3baLCnxSMZTQKQsuhamLrnfCK9ixCdx/Pb7zBC2D1qS3KZivhNj22wu0VoYxOcW7WvBriDCL+iD
/aCl5xl/2XCJL3YdT6/gB+uFSZJtGrfVau03EIXkN0X5UPJe0VZnNyE4JjtOciEH3CksKzy6k+zP
qTojscW9F5sT3TVTxT7QhPRRk0BKsceFkw/PrLu/ZdIqiM3QKDESynxkDs/RRejLva0hkeysS5zU
KQXdCGJKMtBPeDt7watB+JR644dCLw0gYP8SRwpPpn0I7kxYXI4Nj83bSLNHHpGWzOPQApGtcM55
DHZhScqmvVRErOM85jTxxn3ZkXe/GDZeE+1DnxgfQWiXCd3oqNU1s5vMmiMO/YbW9gdjPShmBANc
4LUzodipqRZTbhNqggE2xkfsTjG5RC1M4oS6LjozQ2qGU+cI2/K5Qnig/fnV5oFxd04GMq2uBvhe
Mk9LYXIozs4rRxi7uxMZ8NV+YvgyieeA0VYBzkhKklqADQNYoA81fWTJqWNKIonsF1fnXJMNTDlQ
F1sgCTTp3f/WpSAKqNPk6ojpgfVJi5rhlZrl2z7m0OudgyE73ROB+c9RnQnJOT0251SaCEk7IqtF
nQt5SH+8EpozQvY1Vw51Sy7G6boL9WJg9iUfR+BCe0ZhHKMbo0UqKrFlHZ++cLX+G08Zipt4dZ89
vXBWs1jI/CiZLjh6JdhN3fH87ROVXdLpVGZNQHqziTZhpMuLTAXIIvJQYZ4tMZSHzk1cLeEWGDgi
XkqRf2cNAELOUnZQysiXSFHJJevs9pFrhscskhmujD/9CYI2MtAac/3+UwvXWJZcHrWUGn5Hkasf
uwqgxt4S5oLbfOcq+RbSNJglIzzxYwSB85eg9tkDtq3sEIARgMa4fba08TI/TBIyGwmcq7Fk46Cy
hUiuEXuAIW1EfFnnFh7KMidf8wTvQtokJmXjqXLbmjxysgCl+e6Ub5tPFUtzxhGnRYPFODZqnxV+
6+VK1ovYEF3i+ESDN6lyowb3R0+hHrfVebKTSO99VObbzpr8kwqQ+F26DW+43off86PD9FTnYZg/
zFBNsqu6d+cl9fGIcJIp9hzr3tMezbIhfjMR+AJw1L8qGZWb4bbvoVNh7pDaszPFNaoK8LxJKgHc
trdlaovmBIOpc1Oj4y7CBmNzB3mHU6lE3ldiJPFQfP3c4RJNv/vxxDF5sXDkvF//6CYzuCKgQOK3
6ULX5tO1zutWauZ0yX3Wqq3xJQpJvHzBeCos/69UQUFujMQjVb2yYluWNkeQtWFwwX+JD1Nlw2ai
q+LIYxKj8WRbkoL8BAUbv9hd36isn4DgZEHviIyOaJ0iCztyZahEvDM8YzwfuL1OLFMdAbwzbyqJ
R0G/Yjb0Mi8/mSafB0Cj7HyFG4O88Wdi7Ls5LnMUUR1aSSUV1R7Q42w411SY9RWefq5uZdK+YRhI
5ZmQUAP4PWnz0G+as1c+UiB5QnhpK6zfwT1L1yL8VOXs8zUc3TEURib9QDPGgiGhjCkBpJfBtQFF
hRPY94JrQeA/BOEjecMOVb3Y7863pSK/2w1oir4C1x7XIlRhJkpkjNxJuQsfpeWRvAqmZgjlcAxe
Vd6tgZdPUIDlCLYTgXKYr99jzFUcTKf+ySQ9NlytNESqL645pCFzxxmx8PKDlEPhV4fVZmi1UbzU
WgGAvv2rZ+PSycsNFbn04IcKB550l7YH925PblsdIYlKY6rd8Gy/WDUcgDoKdqMuEXRD3z+BDcOf
UbENB3c5++anz+m+B7D2jXkwvC5ustiiQfoVwyyA5Erh3+B65z1D31kUXn9zekCCtCrunt7X4hD5
HRZHJduKrsRNv8YolIPPEOvo9PVMkBho2gEyiTaW0Y8V9EXnTUcyJgcY1XcCQNAIZXX6SsQLgWwv
RGoFnb6EUuTf/rEssa5/Gvd4NeP1HvkYs54Cp2We8bEUaIFHZCdaF5ACUUvOxww5sLUs2jNWwq7f
jF4aWnKOcRo2Yt0SL0KaIqtjy6FNac7DgaRO4DH7yZK2cC1a4DWp+nJ0pYjFquIL3nWDjJkpvJlh
3f785yBBh6nzIDYggYWXD1PuFZC5KyKJYDQnUJn6I3cSOn5/y5BHtrut27RDP+EHf9n0mTGEqoo3
BG0/x/jR1ISBkdgBSFaUn6D3dlBGBxeQNcfsSBsSdUO7RaULcf9SWU6obyXfiYrb8dwkwx2qVnbZ
TBE5NwlxHm/uthty9mDSKbLJnDtM/Zuc1vIdBwt7N8fWS7BYqhGXZTBnGzrshcCiKL2UfvuxtxIC
zWEBFkx19FEdUHC1K7NgDdias+uh3lR8Q8UQ/2PJrctb+EOrqRD8xaUZypql34fHjEJUaUJcES2A
CWIzIzUJSXzFfdlMyhBgUWjT59MJ3Q6ym4BWWDJa6vid5a+GZUBFoOlFNDmcAiYTxgpWmBOy4IG9
1tXn1vnWgEzZjanX4+PamXvx3L81Cn81F/+HGKEPsVGQskl5k7Jz6bZq4SM6Le39tLohY4HvYhsA
Y/6WUKTTtr1m/4Fq6tRp/5xQ3WgVRdxT42eKerzxC2SINnNYe6OZ9EyL7NdGd3XPBlZuczQE99zn
4+BnHp73sQ94hMCWfDUv92zSYEihYQfruUBhCMMK0//001mtLCTAQaqEkLkba4yBMTzTHdG58arF
PqeiX5wjSVUneIP2jrm+4pEHM4orNhdTBWkT4+GuZawxc2V5HvHtN8pI24BA/sqtFco6NEaG8sok
Vsl1A0WsZQIUi6W6Or4diH+a8P63k7rpVoJKc6NRps110Zu37f7IYBDMzetxg5IVxzKzQxQOrzPs
AZm6/TdZ9y3vtGWbHimidNXkkLCy8iKWOLQYIl2deaeUrKMU7egtew1+vFqkc+cP2CNdBFiaHyHx
96C5I2Uwz3oeCMlu6qIojSK3jx2ZcMxZ6pHj9U9kyYC+jmfya7Rjsy3YC2HMtmKmzoX/ZBnzr0jH
vKG4dxdITF7JdHYxfiDrMa6uE9KDUue3U32DH5V9OY1eCXc6thXAG64JPlKl6wVWBpf4ICGN58H9
pS2dnsOBhMopIhXxYxiESr3RHMoH7W/fcTsw/me83Tut99xigAMWm0vaYN4bZ2PG9HIDvpbExcL3
XRjLHOBkT97mHE2E0nhFiaMqXDjuxqMxcFkZPTPtU7CVD7NeJl/WjFMQTIy37fyyL4fSEIZGAHfn
6VvPjHdG32mnMlm7HdyH0qOpb0f2WuSNdSiNrcUQTUrr77lxI2lsSxwAsmDKK4TAhakntJuJBSsg
vrHMmUfoJdHEeo6/bAofE6ttLwcxRihhDgLZcdvmWTCfCyYmoKCTgc4+UlgZQd4pPJAVrucWQyB8
zWmMNy1sWRtur7Xrd29sIxvBeKjHeL+9y5U0d5FZ2q7YqqTesXeRjx6Szl8fj1eSYZlLmN8RHn7n
ci94jdcVP4r1r3rptDWWkdVDmZCaa37ZwYl/W+ytbXPfiralou2RAxuGMLiUPtPwnRWxDGNVEJHB
UHcGnJARL/VT6kZJlOJ23TOY8A/6MXpWuL+JL7fY84lEup4r6cYZSF9HHGd4jiH/fLkFf40yxr0I
i/C/5dHAn9leiS7UfNl04KTazaU8PxD96GitS+se/e3yz4zhwseWVaWsGgKcTnSvwrdBC1rJZggn
mIvc+6f+8U2suicqQBQmrphPnJWZ8Q0i1hHZtXuEeFl186YyPXgJk+zcQfmkxiGNkOmedNh9/uMr
osErl4UlAV5kp2iA/+Fx8hvsd/2L3W09dyY5zwPY4id1O8DJlyXKm2dmXCSCfiLl0BFMynRciLfl
Cp0O35qecFzlrlt1uRPOAVdoVSsoxT+9GWgcNtojbU7Nv6Qa4JUDMcFioPAS2wETe/+Km6SvxDTO
Mehja7kXW+X0XWJTYmIDT9UURBx0wd28TxDpKNo041rpI1gSW7KDWR8RU7ppVAvJ0gScGV7DTtoK
2/3o3hoEIP5rfv3F/UbHXsgYM57Pp6rcOWyggbo1r1ziC4aOq3fcsa8pPOPxoF9slGU9Q1ReS1gK
X4EtPmunnp/c7QTw5WS+f3sdZYQzaksLwBFdAWLg6th6fTpKCpLVmuyxwjh6h44H3xjN88DrWAOY
znmV+MmGJqM+GvD8PWF5KxqWhmsfa/LbC2Mloc9CFtMU0bbzJrV1NRJWmxXu+I182Z1St5iTIeIx
qnQ/sun2taHI5TvanpXfg7/LX6eOMYllqKG/j6+ewUKaIrUigY5ok3RKE0JqNZqyR4QNqzkjONBd
6KOPfVsKV2RwrunCd+jNSdrUziL72IdqpdehXFOUjqScW1tcK3C5G78eWzU41mZxyKCr1ndJw65+
Ikd7Y+SLrD2kati7LkWyZ29JvY9tKXn1jRl36M9M44klnu/VqA0W7Bqooj6VlBOIs8X9IjT/pgcC
GqtvfmRL5bf98S/WoZ0DmZMow83HXW7o26cp9ejbe5aewtql44vY688A63gQ5waiYaMvMO+25UgJ
1PXijCJfG76EwveIMbddDkIN40//ym9r6HyC8QN1V+J+zvE2baQFbvVXF7zgqQKsMoyULVZE9Xnl
K/rj9txbhkwK7Ckox9b69WYOiuzoNPza5cuOCNjOaltUjS97eUCPipPKHP8T+lQlPQtIPIMhz4iF
NdYOA0mv39Bc3RUiez0U0OEp/l4swfX2w/ZQjL9FVKMLyKJXAhSFKXEYPRBeaVP0fe0CY9uhQCrr
9N6njddAZNXZQFxJvqVA9sJumdMN0fuebt9Zg/vvkFf9Lvd4ERbx0kdso9x3Y5i+4rf/lsNrQe9Y
cUnaHNbzG7pEBsE2Pu951Dhp/qm4q2DKdiMpnYs/YrectXX5bqf+e9o0KonXsFq65OO12tyqaA4g
1UcgNXnTD3wBl384sCcwLNWJgDKFDF08fFw3t9k8uDlSWI88+5jP8X9Z3CdSBqCp4YBVfLrdRZv6
KC4dL1L5kzpKVx/T3IYwilLUsw5vgofHwRzAsrjEaIPkK373xWj38grkH+6Sfx0ytTE4yi/RTBq8
vBEjyGfkpKyJ8Q21AmOqXKIwp41UqhxIbo67OAKiYUdttd0CZrs2tuAlkJXSUyCCZQ0xGLDdgxrX
gt8+zaLrzqUMSm++Z+8NYewXYYxdLmI90TQntxjqnUXEesQ7IOZz7eqmYAmHi5yOAeNYBDPLC4XQ
yhX1cUcLR5HKh4gbuCXPzoTpAVG/SEnnInNDC759s/neMdpFA8sz83n4qdkzGSSU+Bzft0istomO
1uH0HY1ucyUFzczIbAC6Gai0kYo54+xtd/uUwio5iQFvATiCEbIiJorMAiRne/lQc192vpInBwEH
3YcS+NFS0pBcnwM9ZyNfwsl1ssi8AueuWj6m4vc9xJbCycdxetmB5UnnG6fDXfIk8BfG9tAksOza
iX1B/M6pcNFwnmFW3Sw2uoZFW5MDlCX1HKlFjgvqFU8+CRTDlVTCTWkS02Su2B1doSe+AZMyo3sS
IbJgPTT9xEnu9n7xs/auwyX/ZseLPpAx/eTo7FhY2bP1Pdqdi7IDl17TkUGdZlstI5N1+0weEeAa
8z5z6AoKPAvaxtGE3bZM4eOt9ruXFwK6Cz1vG2YgCfUO65to8JexfSdX3o3Lo3ap4Vg/5nfjSaST
tespS5diZNbKa6Ss+IdhA8dBo5z+2F+Mhqnmpdh0ePG+zOzY3wycKY9odNbF7Oyyt4Hq/iYOnXbc
82vjXxc7g5erBI/HC1ihSaCn0fLskemCclF0EqxGCFJqO7nhJQkwh3QGCumprRWV1ohBqJOH44Wj
W9JvC/aIsYoRaE7BE9ydf/PD1/HVdi9jeMFcZg70y8xuUJRPp9hZpbD3UR9afmRDojsZd+NacMH5
MLRvT6ufPYrKvqU0h8F8D3+Ug0uTZLSO+jtj4ZA1vnaVJwSP4tgEMgBHz8PCXgPCX1VJ7VqVPHTt
z2LMmbMccIYtV7OnyR7pBRmA2UmTVf9EruYFf3lUixjVjp1DmMClXpicPAOay13YsCFImGj2x8M5
fs7w0GemGBEC0Y3aVe3l2GSMxoJxaP7GvmmAMHbukhXxd8EZ77DgpFZpoN3Fb3/Iqbm8c9b5baCs
KjUztQQ31/pqJA7eRjsNYmCkZ1tX/jvsEv6voA8hMZf+TE5hlGzdM7ZlWOD7MRIJmB5e20o3qgP/
55BbsNm9YyG5YeAGJnuWI0BiFiJZ4aBfb7nQhbK8zBf+tHGad4GHaDkdt8UTfbnZAZrxf0BExvfc
Xubb3tUy21Ugv91K1ZY5HC8zAsCckovvflkOLOuAhP7MY/gaAG9QcIS2sNELC+KFlhW0Sc+Sd7O2
WWmwt5lWMN8faiSN/kkHdE4NhB1rdEwbGvGUvljCrELmcd7B66d3Sw0H7XMt/DvsKcJjPFpd8Jeu
R2Qu7o7hqX64bQVgzatg1hnATJVYar7rTImGiq81vWZjK/29rIQ6p4nExxh3KA3Nk6fXA2cU7Ho0
sLn+XJYs5/VvwkPNMkUGClwBJZcYHnQqccZV2ss1re/kOeoKgl08+05KhiDK/3mxNGSI9M+2FGpu
4lrNUIQ/neGeglbCzc7Qc917OQ+toe7M6emElHQXYEyUjDIlQkxEfvikTHWFlfu/3JG1h6P/rC9s
k6SSKs4bSuQyE97XOir+7jsYdP2+IOWZ2KboRMwMKUCZTKQTNlpv19MizNEStoqqBQfdjhVMjm3A
RoyEpHxQIcPaDkb4PCW8idhFi7M2Aj6ZdBYViTOfEKrsJdKG3igMOJH4twLupijMN13t2J9gFN35
QZc4OjRYH99BwY7yfSblfqNlidrU8cyWFIT+xB6NfqE5yU+i3CckEp7QAIDAfA/M9RugGQXDOMS1
qLHEfVyUfHP/9sCQxW5nUaLVWuNa6WYMZUo3E4qy2KtT8czEAGw6L5xtvzUUejldZ6J8jIPrOG0v
113YyfgaRilFELjcaWVeripC8N835pT6qsvT3HKYD5XXnXX6INwvg0zNwqkaIGbg3Ye0PHzaET/a
8LPPG2p0mq4A4FXgCCvtJSAQMJNdozP4UhXkXapeDu4zFS8rFd5NP9iV0VuQ267CUD2igagTISLY
SZIG5/8227B23axXSnV5IFZN6iPKkczodhAS4tOgPDtRgxHKRXX2UaNHbMGdgi6Q7gCWubWQd5UQ
Es0NA3I3ExfYQaNRy5SUyns9avfhRZV9YA2ymkUGVa7+TRwwM/FMhc73Odjw+oFh4ZnEC84+mMRa
lkh3mOA2lQ/fe7iafUEOIwRcdyOqORbAbzPXC8wrWYqvq5g0j/wycSWmLTZxwqo4bdq84Aq8ajdJ
DKOPvBlFsPLvPy4Nwypa22+1xFqUVCWY1agY+udGR4qyVKmZqSyp1pFf0p2+5wyXbOMOW25cXnD8
TbxkhR2aJw6AtMSl3Spx4FznoFb+i+purR4bTIYlj2ScMejI76ubndY4MCmoJ8fjoaxq2kOc2QRh
Z3rlfxglIVoEPyiZ+l+E3Vcdi8hsU5HlPVsEG/HWGsN+pFHq7lvOJNygQH2lVg0wrRbSpUgGZRel
NYl24YjhwFFAqxAP+HTstBVe6W2s0UUDcOjrYeFiCpLEk4sX3rQkgnxEGg4o1HzdJKoZv5lQ6GCJ
3iI/YziBhVI089+ITZhtm6xqpgiwUQA6fZ6FOOf+PCgQbnPTPrWe3lxVLSu8T9r8upBi+HBMw13+
vNbxvSjCzya4d+KkHfqUWLYJrtwDVme/QxScnZARRUhng4evQHUjFoOfcb/Rkj2cjLLHAtZVs56L
Ahh7oJQtAnOnoqSeDnUfRBImYUYM7FkeKgSAuFMFUh1/VCzJpcYX7ZRQkMdZXWUQQsa+xtYmeLA7
Y0FQzGz/EPqz1ecK9etS+d7EJEn+ofpH7plWZv3gsWEXHrbbw3MsleNK/SvjnOlg5xhM5+h9q+52
e71QI5my2O+qveKHOE90pzzgdZxUXbPprSUcaCmM3Z3P9ZL7VMD+51CSa/Ww71fpzKhaRqAgcc/C
CCW6HIrc9JJRHKe7ccABBbEn2SRb2oDbFo8LUO9KFSEUhwWX7ZlT1PfnOtKvx37abtFoSZsn3IXs
vR2V8Di0ykcdKBHud+sIZ2gWSKQAa3OsREzfBoS+YXjwwd1jzn97ILHUgQxrVMqCsx1yLgW3DlIJ
P8p6IgeekOaWNOpIs1MmegDCui977yQiUJVXoqh7jrRFPB5AGT2Q0NH094ELM8EtzEqLh/GGEeud
4wErTK5G0fD88FSF4bHi9sLLrS/YhHSuwPfMONhY4UvGA7cT+sHq7D+9lUWe+unVHUQcDGtOmZ4y
PK8J/cGjlMSKWyF5YFnDWs+Mo3I6wc0ha4PDcya4F/PE7qlCnTN52/ih+ePYl/EP7QtQZ7oBmGVv
Jh+qXLWqf2pNmWMrxjOACKZV4r0vodCRJBtoHnEBCG5o54+lPd91WyDUZ1rKXmVkVCs2YZZdlLtB
pmSiynTLmiT/lEj3Ouu4GPHkifgKdC2G2XrzKg4D7QAoyv9t6nKkKwwTYO8vXFCNbS5s0pBT29cJ
h48XJ6gIPkPywlVjNGHpnPsCOqBZdSUoxh5zhIH12i9p6UFRwV8AJe8Lp1gT21oLfm8FUSQxlBdq
+yFfcdILXEsp6T5RzxDdgTkWq8feBJ3WDCJd0eyTElHKT7iib8wDk0AQJd3dYLC/6Sng3fXI4T/W
KrVF4MzHp6z7jB+ccId0cXY9GQ+YcIzddLbDwDD1qzXEEj8iR/CQyEgg+27NM9HKiHBUbN9Et6SZ
D65PeicRdDrT9EQxLKRsUcF5kBQ+h8lvgeLxK2dRQ/pZ9/TLLpys4CkY/zGSTzYddHBaUozaePe9
SlEQYmdr32Rl+UgNVmkZdYEzKrGPNTObJDL+tOLAO+08ZKWmHDvmuX2oAM7NCPt+QvXRRDdvsoIs
BzZKAeMXvGbB7rIGHEsZ/yXs61lJ9hqDfHKAS8UE4GN0tnO5gg7xltJS87c+aLa0lr+6L5QiJywu
0dGDvgwnjPV2z/2fsLB2jna8xBCsWzXc/ztbh7r2oBHMgyTb8Fgxu2G1Dku3WvlChfdDzomf4PMY
i6e2SjMSzFxCNBIlsV+mWZbAxqwhGcehKqDQrE2l7H8tTktIEStqT8OHMQ78YGW997zja5DbCRIR
ZthjAsbSgKb8NYOHPI8vOmbDTY+wxvGtW22o4BD/xeDaXSxgRXND3ZPNWAYhO229R4RG93OjTgIm
K25t6Bg2i/nOPiAmMKxwhQ3A0VPId8Dq43HgYQ1PzAzTcJRtvJf4LMIdzCIx2od/sbslbaKwrEJ4
SX3fMBKrsrp2gBVnuoONlDe9VJ1or1quUd6otxz8Cb07O1VuPQZDgSY045sBkcpuKYGiUsa4O+sJ
0P5PWup9JokFzny+bKrdjm6Ewwi5p3LeQ5H6/LDluGMALS0hzj9z2B5+mpKaFdAgZ8BH2oaPHN8z
V+3PD27JhSSf+HuyQ5wHfKKPbsXEg3I/q8vK6XaQ6GpXL6LJVVcDV7xNwflwZOtHJE43QB8OlwwW
8FQ5CchDQCF2pqz9jaqRQIclEIPoP/KT04rrDtF0ynCAosEtABjRv9SYT5WOLmWNVpLKQxmw4NyE
qJ86EJP7lkpdKqSBmOaU/8dugrtRgUd7q9WSTz8do0d+z8l20AxJyt1Zv0tprcMavAKBw20jsq1r
lE3SBmjOU55o5o+cdcJY1n7awprwqgJnfow9qKorDzEpwlbQFd4HxjF5ZIOApOvnmv87CbcW4UKm
KInTzQ+rpAVA/JzrwD73SQ0vPF5BINP8SxATPvIqYhTND/YYrcUkk5Hf8JPnQ/XXbjGF8u5f1UYF
qDDvzeAfRnIYvK6E1cD37RV1jVS+XgVz/2xK4hL6PCRKEwKenE61XQb1jVP/zH+M1YgTN+fZfnYL
FXAAwW8JE9knnQAbEXw7Tmj7gDZM+HrN+88NfmJGwwjuwtztyaQk75fv4c27IjfcjEN6Jcaclu/S
vu8b8LU0OvL2g9kU3+e00tcTz2YG196QFPe0v34mVTcfUNImR6c5YWOet+qzcP3jFjbCoTh7iVMG
kGq9by9mcTeBLpeLhGuUBUcmgWkzl0agpaDlbyLDzlcUU7cO6llVdAoYEto9C4NRb9IvNPSCcsIR
PESG1WjzsGyvdz9rbZhFhCFw2JMh790fYCbhynKH0BYSkp9uk7mLD8uD9XYkE3kPi5s7OPDcTT9Q
bvynQAxWXDzSsRr/RQ4MUU6SV8uqfMabmH6pQLSBRqvAxQ5Jh7UN9JI2WRoczSpSO1GCcVynEvR8
JSRqE9Z/R+6vEcArcBZjqi3LwzzzA16UHOt609g2H+edETw0pUMrTNB17eqkGVbFYtKl5N4inFQ4
Jn2T/3iUhVk/OWJ0f+sORPjjLcbLhQGnv1HoCDis+0Fhsxi/sjxsyl+dH3YJNnismtcCXTwcTwCt
55M21trAJUmwAYWZL4tL4h5VH1JnYY2xOSQVhXOBEvQ59TqpyVnNeofAlyibnhPRh+MFikAEd+iG
hfoX6eAYnrzgFNj8E4uJadsm83K+gYJqhpJzNM+2FtiOcstRtFPk8kBrUafYkz/PCmC6gRMDWTRA
bEIcNIZWqRKWLl/ox7F5lj1Q5bIQPnsxCPJQRAHAiAX5Z1HMMnAPBZOAy06iy7wijcW+HJ7Yeooj
hpCucyNHzNRjraQ/xNfGHSlwzCrcXvtDceeiTNOQGtcoJACdSrr+pmKnA02Hvl+mmXqGb9hFr1R9
Tw20qiCdFBOQN6zAsA+YOKuvRTdBCdvIy0zeq1XE/BndJqR6YmlHukT7AdPbKHaUrptcQQeVUj3j
xC0F++fOzwe18ZGQ2HGv1x35oiICIEGjp+35P4OiIG3TUUBBeNcaroA02y+IBVFE9/uWKVXklmEg
Jo9V5325upHMtyH5LXepov+AFftbEb3BBX63SKAB4nkWpLwV/LOC3slOA2EXwXH9bwRH0yD5aghA
i6IQk8S/Lcyf2rf78x4RrPTeErgs6+XmpiwS7H4bzTDhPVxM5ce0DSQ685SH6WgIp5+QkqiUBfJ9
Wp+Wn2GWgW5r92gQ3Zal6rOyTLbO/7SAgj9LXqp3vA1cHybNgav+pcOYNdgDw0M1cVL0GyaStsZL
wuZa/ZhcEPi5o/rO/8pmj+k7TKJUySQ03uez5r1xpcgSqtO25RHSoo6GdLA0NRSYCWMzl7UayPU0
tJVNV+AG12V1O0PDrNCSsgkzEnFfHQJD2nwaCYMYtGsxTA6KTIl8xNzrqxgkUjwgGV41By+x3ArH
BMIBjCJTbIuQcvP9S566EJdhvBBRQwimFIdeulVDZ6WCcT9GA5RqknsM4iXCC4tySO8SVWpJyXgm
kpYce5TSxPfh/zfIsNQD1DKe0kHx3fAD286wpXuPp3jb7zSoRTX5lJAPS4FfIoltLKwj/qNwVbz0
TOG+OZ5GqU5LuknTdWcqvscqR8rxkNcxR5DsZ1QqRBI13y02WkmmtGbAXVA+R9CtYw+KZcbczLNg
uCjhGQcnK4bUPMdxn43yiQn3i/bLTmDBK0t4vsmfgYxHqYsPDGog0eW4aDFlTnPbin5Q9OLOWjSY
fP/lK1mX2R3gihDo2P01SvSc0/Lr9Sbkjz39GI4K5EfEtWVLXEAi4TaZff940AWz+VjNdhsoJJii
OT5WlysYsk1Wh+Kv7MMEzN1iYhLWSYU/hsTfXVD69CxXirN+8BwXvug4o56oXoR+qAhUJy/7lRtC
k/mUGPrWb1DwRq9pTwcc6lAhRtpRzpfyFa7fdKyxv4pv4y1TiAND29RuE1FOC6nw0XI/N68ujvJl
UdQek3vtlH8+5MGTpJbfluj64zVVKfeeeeq7OkCqoQpW0fMJ4E7fK2Nt1QPQu8IHqNRKzPdx36Fz
eyn2rPm1FiwGDjzD4JMTMT5huRqQ9Q+HD8t/FZfu19qjaoodk5U7qpOVBhcnSlF+TiUy0GXHfqKt
rJB89I1h3Gl79uy4wZHWkEKLjNHr5vGdft80jNoee46GE/d+D8arJvOqYISbujhJ2YylfXGmo2l2
qAM3BPwwAK26dns2lP9M3ez652GV//Uf7N62SENVmixNUjXlwFQF8S2LJZ/wk5fx9pNgmvQ3ymOI
IR2nx69o+ZQZ8LY+mUtIWOCzj9V9ptsWydge66rLs94dGUhYYzZgn6eKL/Bwn0XU2Obpd4isTqOO
p7E9hIQztTlb0jhN/Qx0Zh0xPh1IjJV8sNNcifWhnJcU3zbgXVAHiaRyNnbFxDpJ2wZ1+TfbbkAU
2ZG5WduI6mp6bB1NXvIES19Ejr+RW8aihDyWfYdGbtNkEi8n4PlEZuM+JBf7EdopVggYdHc5B7H3
tKN/nHPvH9J7A7KM/CvB+C5Lm95xGNhf3v1DGjzI1iCRloTw7rBRc3mYBeJ/0gu9/HiU90UfILCo
8fvHh1lSnNjG/bPKCqaxtRaGHyH6FNtCc+Zmw+ZgW27+P4wU+QDI+fIFBA8u3qMUQdp538DYrgWU
FLysfmVYThh7jTPDn7LSVF3fCNuS9ylkJoycR0E1IubEEo3nzd+KeQYn9Q1uT1rlWu/LruT6NVkX
u/BMxS5BkVXqtZCnVo/ux6gV1rC9ynkUu7Wm7FKxTIZebWZ1KNhUCToavS31u2Gb25Hxma6T+xin
ZZFfQD0WHogXMSpCDiCE8RWvdPpUR6l3MedQFjV/EPIMSilkyMZXz9LQvDg+nTg95No7/NBf85o3
Mg/Ag4q9dQgU1Zwp3rUnb+7ry5PIcaxhFlVxMFzGQiDZDk09cjmcUhObJkRicr2PdxGEl9g7/OWO
UYXAOn2FtMsNa0mqSE4+EiizBxLEiPr2NIjcpNgf0HWwNVUj9ZdC6EfSVzprv1llQmC+B8xZgdWC
fWnssmWk36OuayW6euQjDmty3Ccrik4cxrM8UsNYtIhhzDXyG5s5Fe1DUuR6dAbMNXdv1tgbsK/c
nS6Ne1ne9jETSya/B8YOvv8WjLFpO1zdJvU2PqmvlxVsIUrFWVM0J2VfCpf0kaW2kw0SnKZRLd3Y
BrFo18oYvEOge3wQ9dhUc9nS0wsLitV1V9MYN+XceDrhzpC0qa/ytmB35gmjRJ2783cGJPfA73yx
shd5hEVRFFhu7yr58pNQTntx7G7Lh/dcTDfKCNEOXx6Th04bX7OlFVFkin+WjiExqzjMA965/G8B
9SSxjChlyBijt9OpmaZytsdx1sdyPio2G3Ba0Fk56mG2UOJDYEKxHPzDimIjs4SiVri6OTDtzS24
7rVbauUufV2HyMbdXIHsS2OLAzZB18oIpK7Utv6vzhG1/7Eeww91GDy++mrxVP/kE84qT2Q874Ik
WqfFGuk1/ZWhe+tR1MnGO0TZzDgKKPyejZ147DGNruhn28jSaeakGsVj5rkZDm+wnBz9Hrudffgy
dQp7PYytIS5geznpdwArl3lW5wgwa162sgY3ucRW6QxHrhy1oQ8s1XwaJy8LZ7PxvvC3vt51csqs
v1rP6JfO9/+Ovbe4A0/WN3pzHPjra1vBW8zNmRAyAoXanJ03qbmrDzg6H3QCSL/SlZYENU6lD0l/
r0vQFCK73pnZMXOCBd2UEKcxrr+sRQZFgsTjtKZmNmhSe9mHdglj46HU8Mcxy1SBF1J/DK8kUChR
0oLmBya5f7jcfDjAaia3o6gCvrgmJS3Hdv5yhN1r8urV5/0xQ0P+wlwAFQSe56DC6DlrT/WvpOPk
mGwpviteH4064QdELbauhdl610l7iYiCnj0G8NYpX0h/3hq1vY0DEdUHIvaLuFrYpxKB+OLXTrUS
0j038SCay82fT4NBxR+TyTA+G5saAe8nNBUf1qY7LfDoGc6/EW3TMCssL+2P2FUfXuJGQGSZq3cW
YfTeYW5qLax3ASl4TDxjfMPVf/2MZ+cI7lt+ZWK6scgLJwfTw9v2oelvZbgBGlg/GIfhEVwBmeyo
zTI9EL49lhg8Xi2BGJv+1mU6vDqt3A7nFGBDL3k9j/vFsSpVAOAT4CEVxw7ecAJ88KFFBH0v+JCJ
dz692Rb09VZaWlWndHjnvN7P65xdWrN2he/8L4k7Yel1xoncTBwcogPhxc/oiKN8vX7Hck/YX+cU
nYGIV7wwABZbMfttvSjSdpl27va0KOLNSrPCtn0kZGPn/rZmZGqtqfFpONZVOakGfofJVdrRozw4
nVUYG4VwiYr+u9tQNDcz8Wr+uxgcaoSw24jFZGLozGM/B76YvNbGQoqq6eG69GUy/C6d8trHS77z
jz8j58513UtRIF1pjHvTjK4veT0cb0rpKAu98Lsie7+qn21l2EZ00DInUwMOASqD4q+A0RGZycEL
TRstKsAuR1EMcGviwVfMC3wKV5TdiYIkPwc0A8PBDObfWEJFWplqFJb1b/ByfXQTG23Tonwtfd/n
uqjSC9OeDfNU9YHgtA7PcWcjI3/ov7OSKxFqP09iFN2xQ31SMX+oIt8pxdMLnXsQIgrsGeGymmkd
bNlxMEYIKdLNG7ouxjNccqQtAi6XFw9Er9DAzSBuNwhJ9SzA0RWj9t4/kEYbNXQK11w3qhIOteRN
VekHCZlyMcka266IkFgFPEe5W+C9TSdWgYJ0X5qOkAutUZ5KVA7GZnFZcqXPNbRO8WDL9sWz28R/
h30G0KssXeJciv/JNT1Hnxm6UeXueu5fHPmIs/xpqeooZxFMlgV+rX3ElNjftYLF0KKRLqUmQW2L
O/3uBcSc1yUi3yNkM7aWX4HBT40KpZ9x9+TF3T3uRONrt758qtn2x9XbSL8lYBS3kEuvN7/QdCaq
OTzmyTITql/tdZD5mfkyuQ4A33Uk4YItRqQ7hXjiVMEwi5/SwKKt5E4n3FyVIMnGUfZh7CFVlqPw
3SqPf7GP5vtjh8WTBxp1ClFPPrqp/X8Isud4fVEncGkaFUuvoatu6ixaLt2fRmCq+95Y9QkXdIxk
5BCQAUBp7EP6j8YoLXnIfQ3hlHM+9MMEIn744QhR4L27Ujt5faNWS+JzUFJUkVsgFYaXD2zKS6te
XrF/USsccz6CQYzBQsKtyafsPp6j1fz3/TdzhkolEOoff5wXS+98v09PGkw5Oem488AOEM/9+/yv
4WU/CvOxglXKIrIMNK3qVYKShKQEIK0UGpd+Ft90prKMHJ8sEHvMnhh4ux238oKgH52uWaGBALc+
mK3CctY1CPJCbMzc5NfvT7fXQkt438Fw89Xjuh0T9Tu0VnhoBHN5zlo63hXE7mb2IedFEJLboXXO
rS6pHnHwswX7XFxd+Sb++n17cZbilxAimdPs32aujEW2UjeOgDMK1+nTMe6FELoDINwl88+Gben9
dIi3mNlgTH+zm8YiIoVuKUcshgDeNjmJZ5ZIXQr4ZiUdqOGTc20xp1WWMeMY8N5A2kG3Z2W+8hgS
mzprfxI/et+xog1RJmwIWEbuKOhE2LPplzHfFKopZUUjM/NSQTetXCl6XEJBxp5y/Qen/GpKA3t+
lSkLRA6HVbH0FMLDMfFc1/wlgXXbZVYzuIuyiun6S8ErXUtRdiCsJ7zIN5Phk+3xQOQ9vUfvILFO
ne7CLiq2n402ed4MxdqLjcHAs7GvJpWvzLU9akraau/MJs9rL+/IpPFuTvl+K0nNz4noxeWWi2kb
Vzk+CB3AI2c5PmAg3QaiwpJ0JIR3DzcIG5D+ROM9igA2dcgxit2MRAEyK6BqWJzLEshcyakQloVx
mfIRBtvtpMAajJgHq4oUHajSuwbiqSI5PCb5BC+4oDV+EOMsHHL7UKE7UJawV0WQXlm+/ThbGbcQ
Zvg38pn5WK51Os8ZK5qb2Gqi2bTkUr1j3bLS8mk5SvINdGWqFAI3/Jt/khEVLAcjU1Md/mUVk/9h
6A5PmcAwPX5PHNNyV9Z1mHDlWVzFKeB6squ2yFuIGpKj5N8cIPSODiy3bYcD6e3T1GQ3wkWEwrzW
tTrWlohmFItUeC4nTmWxzZB3q9NqTDgFmA9ieV8Q1FSj5LxuGofANS9O6VrKn1zZA6GlIAJyEX3i
bsAHr6lZThr+qFJGCjPtvnV5+hkPrSrHN6AmUmlTuQjEIm0YXF44BigfPFE9wviPuMFQKOE7MNaI
B5F6CKdij06Gvth93CagzVIbbNP2Wis17XmmxDjEC9krF+bLXFr9zRK660Uj7k5/+oZ7gaxLs4t/
ojez8qlA7SfRhuUWS6f4MfRnB7xxXw5Aei/5meznwaGmIu9/XnUtgyMQiM1tQ0XsaUAAu/oXM3GG
5lwBUJLLd2RSeo/VUdJXke6n/XB5c/tS9FVNLmiT7BTVctJYXETmumEJync5UxGoyfPvsewspJBF
FdFRU/Jz04IM9tEtZMZ919SkWTGvZsViMNFsIb2LgtN2YgtgYhDxRARac8VBBuAB72l1OYwjMnB3
aTQNy3dKDOFalmNaeSczceVWCBpXycuK2Tx5kR+7Krb5zSkR2Kx2CyqTSAznqp9WX8FGnPvSYzjx
Sacyv5kcRtOi9IF3qQmdUPJseKN1XpMqIScrdfnmu2Ds1+eWzjTZx6hjDY1iN06N69ViUfgr2tD/
CJyORh6a7GT2YUbbXO1KfhT2cDdbytD1QktBlLipVeQNqpWY6+5JWY6bmKidYW1UPj3kgEmnK9Bu
Q25sFBEK1jjztLrhatWtys2UTjp9xcsV3feqrzSoycuHTU6RmnYfYWqcTOMerpdvCthtm/jKpjWU
cjTQ2s/9K1c/QS3U06EHcfRhvBNcujupT70/qGjgvYGV/iGxsuwUaO7hQS2ieMLBuxcVt6VnUSIt
RAq9w6s01ntaV1K15aIxQfOBCPae3xPqCa32YVpMiT9VFCCLI2EcRWf3DN/1jN0vDY4VSMTameU/
8PSUPryLTJvOU4a7fWU2VCFln5scCniymjQXfxxqMF5aDDdEiWxghlr9rrJtIxe1wuC+ukkzvBvW
nMVF9Aj689ofQ3e5nx9JviAZVWNaH/3tk7+2+ZJvew5qeg9IR/9Ti8nysgYU6LRUMtTI9AM1kJDS
PAJl3AsRbOKL+cJCBW/EUZCDVCQtWIypwSyLVt4pFDcfGG/RH863aoScYc+OyWyaa9nge2A4/PqD
2HF6En5ZGUOB8/99fYnUzA7xGMFoFBs/RTeJO7SCCkrL1XhMa+rVBJfhvS2+RQp3G5YGBwPvYeOB
Yaety2HzhRCsqznCin4kJn3BVXUAH8QhEf1pYmZSPPZtvWJLLEPs1Md6QyPKoi2r8neQQdYda6/i
AlvvbHv5mAcddIHotvBtWCd1mGS5UFxcTMJkBrb5Vgupglj3zwhAsB5mdADGmARmQv8bJwO6HKYV
SgqOjGAJiiHMM0/a5cjryRecIxiycEEcbyB7WF6mzAxEBKRXyELQRbs2ov1mU3yj5NeeyELDScJ/
f3+9zsJmt6xv5y4BptcUk2hYTYQiYsi80kPB1/Tkp/lWQwk9XE6lvyEXZrjNzPVXk9MLLLDxTrfF
OU013fXzSBZ/2GeDYtGv886DbTRPVrTDvGlU+73/yaELfrl6N2q8bQNNrNuKuxPo6YPAvIzsI4jZ
a9d4cA+T4B+vWRvNEGthLTrAPy3jttx1MtIRStEPGOHZpJYQOxtY5YrKBFYuP1K+8jh2E32oi1xk
GiKcZCFqLA4g7ZtU4eNe7PZCbxoGC/TpYyLapr5uR0qJwitLbrfWFnn7AsSMGnCgifoT6Th94IP0
FniRmvfpmYSM09JQD8LEc3vYfNtixBXUdr3vn3f79CefkyMozHYPRCDJLfLAVkdr7mxQlx/Dw4ca
vfxbWH8tFwMlqCN0irpKeeurxfyHTWR0V8gheyVjvte+xVIw15fCmCgJ6RJHtuaLZQU0ce30Z9o9
/3gIzTZQBK8lpGQQ/5/i4Ip+MDlU4yePDQjYvlXhxMLMw5+1NU5oIbSGEkZx8idKaRae8iQbNxc7
2iBgaTMN3GKJfwyiuj5+BzbZpWXEoCN3MKVMbcpZZVfTK8+OpiYQnF6DRWTZRRaCcEcpOcydUl9N
xAOK9wqSvYJOeblZ1tsOy6XTiWoaxcrgtXpcL2dA0L74gd2J3UyQAjaQ47EfmQP/uZXhFn1ufILA
OVaF7tf9r5Xmpfzk1SsnOEJD4qwitc0ZAtBB0FhbnmkbkZFx4HKTA1PjPw/a0Vqpjf1V3nOYcK5Z
SCWHKoXkhik/QVg1X6oH/lXgrjG33wJfTZTtU4vnQgbi2Iu9hXPBy1xeNp6uQgPvSduG/2VQIgPt
kxm+rYUyu91C06jCcYIWOJ7isbDgFmx7t6MFc323jcl6VvmbzGh4WCBPT5BN0Az8UYv44R8Bwh+G
ZsiY84Vnoy9asJMytnqCKKdDjGLC0Aa0cspCKpNmWiUbE9CASPtwFFdj5dljRl52+EjZCjhqxmvg
yZviN11b9NsMETpd+ZZlzgHNc4Gzvqukw6smQ/2B29qFblMg53R36J3vcDyMAN8yx1ismCcZAJci
Hkv5LNpZvqRbKpYvs/K0PnYGksHLXrqsZc3ByJVHemIZn547j38LUyKrN0DZiWh/NJPPUOutcDgY
MBpPQESHFTCaEJv+plHxSkVKMW80TcOuQczeYvIptkcAf/usUwx1Spmqjqzn2GU+ucE4vgtfDOJY
ACddPaJE2/Zu8nmMGMuUAQpd5u4VLKDGJh4hh0MHrtaV88VHEMqgPH75t0w7IGowXuAwCdWTgBFB
AqQL8OijYb9xrR0rWxT84bECS7qTH+PCjW7dViaKacgEw+hOq+labdlT5GtpDFQXxmGSEmqEoSiG
vidupsYhn8QdSfnn//GZeMbSBguP77Ed6xWfUlJAk5sNrnp2HQHyxAd4NdTxtpRHrRlCZfyWdojH
JNxD/T6AgCppjO/owVKJ1Gwj8cbt6cPshIdF03Cp3onBEbDyW8GDAVsDcBqfzqlTL3Cy1M7riLI0
Cf14CK8M0sdLjtqiJZrzeS8C6rJZChtEzx/TTSCntGs5W21kMbvshjhpbe/KHYE+uI4xVLFsJo88
WsbRk4jmjn5prHKRicRujelS3NVjdRyIZWLLZ7yZ1UryU4vR+WAKzZ+HoD4jrylEEWguvZAhmhQ+
7L1C6Pc95w9jcg6LjoEe8pbBAOIttoxzuypHv43YajDId4j7YQeF0ACMIz1D1Oe0QNi3ZDcf1YDt
B2jO5OihWRFqJiSlPfNGS2nGZDl/5EQ42HruIZUcjiRmOPrLd+qylE5NMAiSlvnMiE/jc1kXt9SS
KVKCk53SOJP9SeZbchgrqEdwDVLxoJ2e/EZbSFFFVbWILv2+LZCpYRAbOY7FAKa8enwWlJm6wOa8
ToMM9bZ6eil3QpjLvIzrOB45sZV0w4PGBFkD8xkqmgexYlDNJNP4fJMlBXc4mM0x7cTXfBIWiGnU
3O1F3ERt1T7CdTVmRrQyjFaeCKXZUzd/ezB+QZGfWIZsoJEu7QLj99wU9HR7SZqu34RuZaW8EOxP
dF5O2zKoFxlCnTFdNjh0y8lR+xwvynpMDD8Gh8CwfhQ4yGkdpjzZyJ/HrBkMAC6HTS1DqI8wrZnY
z0bqSa+pEzXD5aXyc8EQgVj/Aen5UUiORMOH2/+rK5Dcg9FYDr2T7VL0x6hJtIgHeTejqL4W33vv
1+k4a7qUlw/Y8034eg4k8cx4+/qqiV79dDkWAOZtR3bmxqZ6L7GPpL6mBhMxzcOVlIitw9UNyEzN
ZOi85u2D92TI9oUVHZ6h4d/YIvsZFYBLumBSIOmbKQVfNZ4HaJf5D7YfZ4uD5rOLj3Y34/Z5tIKZ
a36Tav0IJaMBf6dUWaWb1ggpHX7hkgJZX7fg4oHogRDDhMZGrJDKlr0A8Uv3WFTrMSea9/QPsKAc
rtw0RbUo+4yeKB8ym9ZOzwn2fYiXWLt/JOZC5ARkLPCujOKM4qS6nTXMb0S601hvYjnX4Wu6y3va
8trErcKPeTRsszzde4/UDDpZlNlCrqcqqiiw+JqJXdBBDAIsXbA2OinYETOVjveqphKDfMr3aJnG
jQm/Q/4usOEFWpGbdionC3vlfXORQxIo/WCrAdgQWwpNeybukgsJxx5iWFhSM3BapXt22WJRDraQ
NXG3Fn0kim6xmvenmgfx+F5daNIRHEMyDEPnXUrv+Khwc+W95YFWtgFXPrp6DR5FZfL+jjj5G1qE
HN1Vka3AGUCTQiSHwbhNZFcyWbh1qe5D4ffGISirPabGEiqpyU6vJ8XMQv0X2a5zsqByLp+b2z0p
F1Ek5pdTwy+/c1c+vgx3G4Qgqvc269WQRhJDY4m2SfUvOi7FfQUao5pPVPkoYVXDGfrdK4q5imkj
aov+NX7+4kTeBQD3EdJ5cn0PnL1mga9kpotLMF9hSR68tIt740vH3PxnjGJGRDTowyv1128wc6E8
2jPBaHGB95uppNqqfIX0TuXXDd9bA7qYNpfdbuT4yiP0W+NLAlmIcmI+Z6nyM3lpZTf2OIcrUpHy
hMLL7/R6xYGqqfa5vqoZshtu0PAo5mZEteFhNimZR5ORTTYUhIaLaYQ1bIxMQAteNeQ4jPOjUf6M
ajhKaY3mGIXLGart7OWS7c+71NNIwV/yXxlE0E+MiQU2aiBXKu/PVrENjiHZbPrpnTg2Xo58MZOl
6/0LPhul1aCUrpJbLSf+SJGqDYO2BO1JSBfyA8qtRrkw31gt1hYUHmV8TtwP/QCDgdTcgrLfXv0J
tuTs3SYJDlgx5EsyUYdSdbM3drXDAamm3DIJZMYGAYxyunsfabpD3reg7ijMO9f3gO02PflfjSku
JWtFS724rVIsMX9ju9gt30ZqBXp6rFWeFdiwje+O0FhJjjU8r8tWRc2vjFT05jrIonXC/U8yUKxl
QPQQ7RP9k7VGrOXwCKjWSjhPJMqjVCwQ1ElCZPJLJxB1W4dMgXqu4s3LB2RHDKbMLhBUq4gerSlo
mOOgxx9HpCnSbnYihLIlEhsR2vbFn5W6g5lSlGt/zZxL+V4POH15zg8VDd5AjeA7e+oMXoageg/U
ETE8w6BNOuYxLa7sb2+bYenjNdMIz2+AI+J3MU8uZGfk/YilMGbBt9/bvYfvwIV0Xj3jD9yT7vvj
dLpFPu1B7Smff8iLjr666Tr1LlkzgZcqAFsgv3b4Ed7jlgcky1aA7+9ZfE4+lfZvNkX66Z4cR6/d
iFg3d1s3GQW2q1MMhXIFI5RJNWkO/l1AhtkDKMNO96Ilg5fPUVeh8bWPYbMRXReZuA76TWdFjivo
hMYcua4DJgIChTeH+XrRnRA6hnMCHPBNCEWkWJagMsB1R/XyE3YNKiZVsxb0cmU4gFrjmEoAASbX
r1vBdSKFd+gQLMxSO1+TddG+G5qMKBbAG9X9snTeWU6CJSCjK8si/Y3sgbxtPpCpDcMlQt0DkZWu
+gQYcv/mUKrmmCq7VRDLahgxuBFjrWcUj+itkhdFiPcuq0EohkC8IaVZVdaDlYt5qQQ8nVpxCWMv
iHZGJUXLNGCTLa8BlLhFUtVP6aT0geF8cf+HK4ZdHfXoORb1StCTll2Ub+k+IIVLTCHRSrQentfv
bbLEt3eRmAzar+e+gaal1m8obxr1xC3S3i0qgNfAHoSEoldadIb/Isnx0s8Qn7SFmDhF9c9EsoW1
ykOWxAkPolTpvdiIOH86SqcrnE//ulbIiGDiIhygfIoYV20Y+cWlsn21lNU3n+E0XswJcFUXTYPp
emkRo0mHQ1uXGuTwdP33SmVL4Az18VrxAV/JgtTsQGHmwuAMoPHiMlOjmOO8Ffmp6YBGbL+SbaYP
z8OGMlTjcHJ3ZEJx6JLiHABcVXX9c1Apr9k5OrGs3VkvUP1FaJSmKuWAadLixQxfvH2Nxp1pFbb2
kcdroVsUsnUlKbisYLJFWXgXIic9UgJecXH8ZSY13CgxdbaFF1OGG+hzjZQLFidV+jGF+PjFv1Jy
PJjfS0gVittByFyLEoP0nB0v6AUlEKO5PEvYqun158RLFLm0D9DfmjQaO+u5KhRR5Krc5F/1HCiP
Z5y9DnPp3Pxs1pKydjlC/79a8CMpz/tlgnudyE/g540ogCOf4rhQ5DhGCDO8j0Tn7WQWXndRx7FH
Wp/limMB5iHbc1kuniRnEc1IpU6fpvQByz2qb0LHQPe4tVSfjrnn4UCWEdcTyevxyxargsXNw5o6
yYpX2eQysL3M++4b38mZVCHkzQgCU3cp7LkGCnzQb5mC/5SFq4hEbdcEsF4f7kLXDvPDoJ1hU7vt
fSYBGHve/kjVTbrdj5aMBvv3rZJOuZZgYf4WZ1rRN4OfbAcOzCuPpZ5V6MGk/MwcAsdJ33S7taHZ
Q8TF43OpUSi4kiRP59OMoW2K8egqXeyuar+nlozY/4wdmTmrdCumm99lFg9T0lwOZZ/ubPl4/1NP
H9ICO+E/kJvi3Ie6JcLY2HNqV0HB86niI9UOu0NvpbPMReRoh2mCUq3B/44fx2aFnErQqicBzUgk
FnRkIuVp3Iu+eRhLXTRTVd8SjvIeTSPzDcPlZK0YdIBIpWdwCrqY/CXFMXKfDWIwhp89Uyb4nIXR
fpBvTSB2seUa+wjJbgc6w7HI4x1RZyZQbepUntI0y+4wWRgJIoe0j+oO8bXMyp/z5+M5NZg32fLz
KPc3ZJsS2cuKio4x29ZZP+l1UgWAZFYsudqWSvBRLchGf6wKaNfBGvU8spM1V1NVr9d/4yjsbQAS
nGgHEnucCmaXTb8Fn0oZq/WDaSBvjbjv2w2j34wtKUv9/5uJF2JRjpO5LcalUio7MZddCCHOScZb
SgVDbHp0KCf7f6fieOkQ2TlIWImcqitaW/kirJXNoDdGIM8uko/KW6a4dLBDH/lCUpC/IzUxTB+X
VElSyFk9qD/lttafnygI2UKuLuCRiRhzM0UTLp1U6sFcx/WdIGi8chJDFuIwhOmAGMklB4iGSd8U
bnTQ/JwGaFkFjdJC33lT5pfppxi84oo1NybTdvmP35LoDLVxTvcESYIewWI5ewBkRNfsRexr1VV7
YqccH1/oAkTUCmD2wyE9LnYl6SPi/G2/xVW8xrlrVO/ffGxLWwsOAb8XDJH2cLSoVtcKUJstzRl8
wEukVEKZxxuoEXgC2Uxt2dA2LDXvNVjripdRt14/QW7YHx59u+eXUM3PjDFQ4ykxmXtC8ECJNAjl
V1+ZmwcY9v6UzrERNfVlCFfozBd5w9LmIVE+Rc3fHaYN67MmNTH9B4lMh5aKTKLr3PAL/Y7wHldW
MjPQuipcuaO4IUIRvBN1Eff9AZOBcX812byeAs1AEjv6stTV3KzMs+4Jr3tR+Ps70QYI/Wamfk3o
QDsIJ0hdQ3LQ59KG4nz1grW9MiSU4eRRDHLgGPjS0Fl/quPVQf1aC6p5pNgRWUf9DhD7dHWSceNt
4voziQv8daY1HRFQJKK0kQ76cg8Q6YCWlbdh9I/n5cHgS4PTtd9nO13+8nH8wo4qE3fuuowdisYc
ICTezn2hO2Sl7XrYeg4bhv0RadCzkzub/jeXWKru3YaHPJTS49AggYW4Ocl5OxCQh3EsxN0deDN3
XHc+JRZqBEZYUz0Gz3ovoiCYJfzAeztfmevlkJS3bHLH/4cuVnkueY7PSBdiLobjJitAe+acnXs/
1jR+DHjEn0GVyLZGZSNQUqDqfVgI1RWS5qFd8MigdrPqXK2z95g76y++f8lqHdW4CViZ0lf3rnQP
uuqRxgBuNEw0Mu2fxDjlF4IqRbr+7oxMO6SSsW7BPAF/7Wkohc8ZIER1rCFSHgTODFxAaozXViQE
XdOiaGyoeY7M9crYZNKdVSfrkYIWXSkSWCtHJVJJVi4StGCO7EfrtQ6YRbL9fU+j3j5uxLPmzw90
cwNzYrQ4PCkHJcsHAQt+FK1GeEdNuoNInQg9xtzWs6A+V/2gE9TmghrMh5qONEDxDKYm+ONX5SCV
+NXTZaaqFlsj7VglgTRULvgbl5ts91Uhsr7/Kvt7bCtCGmUkY6T56qlgoCUnNn4u9ryAU1d5Ibkn
vuh9BYByaaTwAt+GTc8VdcKqcdgz0rX6ISU+VCpWa06RNOi13SRKsvTj4IbZNdcIT6VTm+T59/7Y
bliNyajBDXNB3OnOs48YtqTuLB5BCq+FJnSRxLJZh+K9w26s642dsGd3l8EpoPqYnmjVxRyTJX4g
6bHoi/L4K5kph2XnrnlfLxJSSqVYqoDu10/yZJNitf0Bc1jZInuhmFpgMJJbLQiX1VYDMGP1Y8If
hPOzLjlYGqnKYikMFsrCa26VoiUty3+b3u5DdXG97Nhb7nmF2o1dhxkXJwbCYl7a7utcPGjKjn6Q
SNAtyvAhW8DQ+YAGBN2dOsM5ROhM1VRiusRcISkYbVKP9uMA8/Wo3aaEqkdskqDrU6wk/HyrcC46
ILCXHPsEryXIa8MYWX84nPCuL/pkQ/IIdtKEflJRIE/V3ml4BmvZIe4kn/ZUQc9RkO5eqwV7m5lh
PeiVRz5kucscboEw9oDXyOjRJfC5X/lQgKpLp2dYa90gGRyujE9aITVUB4vit5XpuD2+EjJm8u10
WLHxAyg6Ab1wu4yJJJNOKGBOyqAqVxQS7ncuQEp+QZEYjHmjM1BMSaqzAF4LtQwuC1i4KO9Z11CC
pPJpVKZYu3BNoEO7RmBEBLX3ECo4/RDTE0js1jk3/5/TW2ykP1qT2C/9kdIjmQDxoVnuBDhpwCHk
m+KtIViq0Nu5/BhPWvyUCABtzAy5hwXEtMYva5rE21JH6yFa4eqB8dTEFl4GBXL7DiJNv7YR73u5
Yd0zns3EEAfPCuZP3enNGrhAo3jAKmF/xhP9DZ4Dfj1DxrpdxpcTgYmktUZAbb9OPZy/EBBWpXQv
l60BJkB19JKFJJrgJI93dKpCqGFTciebWTcvYdpkvCmzyS1l7rGsEGXyvNi9WZIE941KoraIu/xY
iLL0wO3rtqzmPuiopGwvqXU06FtJoF6qyh2z3BbwbKIu5w/JGYRS6a5l/q76H7ismyZNOrtbFOvE
XYG4WKTaPOYaFzjVdLB9tR+Nd44u9V8DnycnvhIR60d/A4sf8URKGHOA2+yWfhjTeD9YXNd8zKPE
qPupqz9328HTDrFK/ZITod1e8zMvbPuAfX/hownedWO+jVGuZcukkofctYseXgPxG8ZwvLIEe1J9
Ij2pSHntauaLIYsRdIq1X0INNmvfjGewDdHXXvIOdDAud8xYGVMsUNBDWVkLLiLcR38tvOFnrceQ
0nlxH1PEDt1fh3VxmIyblyfGuav2n5IC6/tn2WtSk6SJyf26xsT7qSBV2eNCqN3stUnGf3p21LJ2
XEplSae4QzCX1BxA7W1uXzScO8rMrwQ6r14vQtuSfgOsm/a6hj47am3rpsTV4XV6curVtda1/rG7
tZftUq3bWeC+u3oFUMSTyHvmtWVqsc/5T8WtBt2uj1ShN2/jwH6QKWGYT+4CYroPqeZ4S8x5+Vjd
hl1e/DHmT3bkur11GZCeO01Spn20fR/xhs+c3yNi/QEm8NonYaLOyWR4Syb0yh8ptm0snOsQnjLK
c0YmaWMqUl5MJ+xHaO+fEBmOfgeLnnO/ANBSv+G2hpOtL9XNC5frn0y7zu7I0+nx932vJv1n6LQR
wlm6v/SwC4MehVC8YJ5PzBGpCWLPg82kRm+Bm7TRbi3Jx+ubdaG8D9TqRrE7snWub6KmNpOw1//P
5rGWGJMCWzUPcnKsUF2CJ+vopMVDxldjFphD6QwxIJ2NWlBRgRtsxGC2StLGuZNsSwlkMfGyR6aw
HHycX/EiS2upCSl4uTdCquNgocxpPhOjVHdyaAeu9humI8czZsK9fEsNf/vgBXPJr4HirWEw0eAp
KtoYVDEDsYTgJ86k4+0FqsqBRYNiK+gWIzfcd2b8+BFsJb+Uaqq6hGSyEjB0q1XhSt/FK9Ui46Qv
dZvBg9WhC/b7eFK9+xCMujdhG5E4wusroP1zjmyhoiVX6eqYXwGQjSHzj0EzpGknH68vjQcGtPU0
3H7oyoXqHMZYZpKAZYalJNLTI078GpCDCNw9fx1OfQZH4kdq5K+zMw71kNCxoc3gfQ4rZw/LaRDV
0qwfz+NRcuYZXoqrsAsSs0Qgu3+f0K6XL+mVJFCKVKcJhZKNLxcgrfr1Db/ascujfiAzGxntbKZv
9eL7+l+xwS/UcngjSbi+f/quTgTPi6A9YBNfbjH+cg79iqueNcqLt96mfMLHF1vu37nqs/8lsZKF
nxcZ00VFN2iH4ITJnTvD/h/XaVw9MlXFN3WC6LXErsQvWKvrIFD0FjU81l7aqaluINrRFyLvrbAb
vmp9ZG8Z7knECFB9x+GKvuae0dYA8m7kaiY0AirLRZIMN4yx8eGB7pJIbVDPFrjyNbyjwmCcHq4M
zGqCknjaT1nu6A3KIwYIeaJ2MTR42yV2NIVxlGFUY6Pv12fK1EIHbvIjlHnJNY3yfRNn19VzLWlF
aViNWgcYm3On43ku8lweF7oIrbkpOyZ3Ae6jx2PsxniEPL1YrgunExLGyYtw0Jby7tCyACECngf3
c9UBpULOcnxj6MVvJuyK0VSmf+5cEiV6O81gViqvHNDzSebk/eWAguZryR8nG933sj5NrfU/WY+j
RuB9cJikk9YkRApw72aApP3NsmkDOlPg42ZkoI5cWV5pkF6qcf793Xf+YF3ac7n8DzcX8U3D1Fcy
wU+OQxr1xT/gZ5RwYgg1ce8nBpmGy4AuiqNAf6eotzCkVdcXNPHhfYFjl8LPZKQQCUe2X/l3dTLF
lBYR5QmxXhnbl3Xz7iuMpmllYpiR5UPU7XVNXkrN4QlEYunlDD2+Wg/QrKT2GUo6WhHvS/iCH2HH
IIV0FFG1gXUd6BXGUeeYcmuoibT39AYAFDihtxJgFSmRO0cHIdjUG80anAnNFX8BRWkJVFzd5vV+
ulwMeijFExZ4+q9Hblj78s4N/TUJqSV2GXhHsZc7XbNkduNrbvqHFb9QVcQMoYIyGGvd/M3Pa5Im
8rWUI4S4RjTRA0r7TX9EqqozCo/QCkkoMYFmqdLcjD81uEpDk5hTxPmd04SSTyXe2+ZOrFFdtvYN
AvPJAyNofNZpuMyrY88NJt9jyQb4sbkKu0n2q01UFtsHbtarV5wMgrJaSHqfiApETif/6gmc9KZR
3e13YF2SFWvdP7z4447QV+AEJJyPxu2CfDolZcnBRlLFtzqSq1J7VQZgQk3o6pS3HJ27ZRilv4AU
z2gESGqtkq+HjDSDyAuxwyF8J2bjK4HZxpgPN0VwY77LetI+5SDPiFJDmUBGDBp9kWdfgnqGSB7X
6Bphu1D3aSW1UEpH892xNK1yfq19E3yCc4R2XjKbcoljALKTRnxVyVxHR2egK29u0+sZgoRhzojM
48J2RDXCSwSzHQuKcbMalQ/iV8RkZ38lw9FNIsUE8H12E/QcPTn35shotDglBm7AiHYVCzfLKCer
jaSQC3yQzHI6MezdyX0Ey68rQ/ST+p5KT8O6anJVUpaXOsQzlmIAlQkIMbg6/wxxBdQumV47x2Nr
yxaXsMjHA6XiyaUAiVKIqP8IEYZYTdj5a9dRDKh5qO3YeKag6xoELcydQz0BqhFZVkbtL5Ft/Gh3
KzqkmjX1A58HkfwF2CF0tbW9fgpF0jpq1C9gVq0bxYrOk5yJ04+qdxHm9RmW6E9TsRmUpxRlEOIE
LBalwMjv1u361e1WP5TNfNIM70PGLx11xd8vwF7aux+DkvEwbTvLgqBXRoGZukOBzrYO1M+Poypx
bXYi4VICYaf/sjYLK+yB6nFQ/Fazku6NBerWPla8VsjWryZQC6RNEGVRchT7O3uMd43RszEjrojh
7JZxH4pQT0EAbAOTgJhnvYKgHkcaKxhCy30h6lMPhB2cDmK+kS0dNyZ+GQIw0MpPMU3khQBXwIzE
aP6BkUTIHTR0v2K5IrbXBqOcExi8Z81PZtZ/8o1SsSVJ0UsD6zgULTJpUjuXfVhFv1BQFGHzO5uq
ht2kTr6P1WqJxYJAJMGrz0qcqffp9rm4uqpJuFRoDS92eenffJoUXQLqSaZgxb8o2JOg73gVOalL
XzqbUCbzGlg8JJKP1dKvYiwSUXDMSJG3Xb5eiJoj/o7cxwFLvcDPqRqKSbrZi8ctfTehmUTLbISs
Hx/udmBqJaWRAnzilILxykE5CViVGFH46EKGmj+HoEEKJ0if37aowxnvjbDliSaUUvK89kO3FHbq
CGnCvokLMIXwapZmeOCh5JcBepAhFFRJiQBBMki+MLkMEGJQx+dJg9GD+/9XImjNqS03MRTB1zz5
A/mSWb6j/4rEjM3x46gzuCvZjmISe73rq8PnJbhLs7kfEzC9YvbYbB09GAHirD24hgUAFbltK+qt
7SiuI20bYWRJfh4zm8rIudSdTdpde5XnS3HRL3OlylUXLSjGAnTfzYyVOIEuKk62Xp2unJvRDL/6
4CIAeje1fXdC4l/zDVCKSwirXKN2ifsviZ9ffDZT9dvmWo9MkhH/r7vuGzNtKomYso5Z9L/MsZX9
swIbEFbc/wfl/crgeEFc2CDvtvxw8Z0zPPTSgOLcxj19E6njp5yfAQLI2JU/p6FXXgDkDwvxVJAD
w00fNQugLll9XNYrkzrK3FnMtRrUYSU/o98i5+5cqczmBThA90vAbtu+RXeX4ENGbPCcQv9CNkSq
eDjAkSFR2vtEI1eAqbPBw84nRF3vB0YR67szlVBWjaHzKXmM5HvA4EqoXqjGGdCsGk/roBSdDtEH
gKy/OFnNASo2sLG4mL3julU0vUx1WlrE8VQkIg7smc4PMyR7hB4vFpx9r9HlronVPs9t8ggum6Iz
nAkwJyrN1tm0xIUCOxHl+pQYxwwS1ccF30qcz6x09TAvmqdp+40PWB87EfNxe2mhEuq40SPDP7Qs
KT8HsiPJqTa68SCYfFfLhHuY+A8h+ZMOoM4GRl9+ffgcXBQbup0LvsgqNKKqClV2xJYR3G5dXHqT
lLvOEUNyMgvIIrD8btbM/TXR8Z12aMktWZS2NXba99euQf3RhyT2TDr641N9faqD3ccSBL8eS3f9
rPaLfHFPfgSQDINjQ5uxC8j8uyjMPRtIztbeUZce7/l4HOt7Kt6u+tkhcXVSY6D9Or2XqO2SNQSe
cMDchGqPR6WUmK6mdh6m9nGYhljGeiOamRfGY2615l78D6XR8oooDLeiR/jgZpsuKpIu4vcSrwYW
lI2uQSqSKeZQE1/1EpyiAfIX1ooF3BaIQvscr0q/tum99UR+/UTXhkWkP3IPQh7tbrQKVMI0KSqM
n1qeOVT2lCS/wgsCaHNf2BLM44PegY5kyzi4/ylHSdQumVs7SLy9AXjxIz5JEKXyqPGv8WiSzQis
DZyPOhPkjwjri+tT1k6dQmjBI1Zha8aN8tUSluem52NvrYyayO1yt3VJH49TYhrwjubJ078swKP3
1+3NSyI8toTgPUT9S78ZKBpbwu4caF8YyUUBiU50hPvwzlAGWMGMf3Lf3e7vlwo4ksiFGT5S5Swl
X3dmc8+iZz/DMPZ0Cwc4mL6dOFm5DI/Ta7zFSTX3AKTgk6YqI2CX7ujxli6YO/LDV7avjaBj6UBJ
Cq341OdbVcDviyZ8HZt3BFIAiOMjK1h/G9GYQcN7m2K3UdfVtB3RuyYA/qDXSl0TqGUNuNIHu2Ay
DKBxteNHvt0dsviLdhtrmXFu5+/igEF2fT+blaykBmNyplYZh1tIDgYteu5D1KXvloWFbKmjLbHh
eupBMBSBM/Mfu/XehHeBu5XUtfnBdWJRTSmVyUtZskjJLOtned8B3vlXnu1f/gMGBz1F/EPoKrGw
kswtk09RIujpARO4aS8srnMwhGJPXtRIY3AceH7++DwckjlaNTKCnDfO6da3+J5yoKMR2Tg7BT/6
ZTSg1M70Kuv0qiTf5rraFjJc1tHYHUroGIMRvblRd/1o6OaFLtACrCMy+tDEa11WXfWH56h7bixA
psNr+ibDX+exEYch+/1nzWlE+nhBAtvjf/p4KoLKDGctRNz0sULpWFn2R4AZPhhQ7oJcIDpvM2j0
phPGKHUo2NdR1nLX2yAIil9qxMTkrOAxd7niNL3qdzRG7QUoM7PZh3bl2EMqbNXWXvgIoHeW25Pd
vPyzlcd/Y+Vq8PmXirEI1xY/EDeIMnkYP4EgxXjN4Gn3HS4KldEGnNZNkIFIfGffDYEiK4u5JaRV
dAE3K2Fi6Qm5c9brg4ksdJX6TR2OYJBuLyqmqf+VsdXq9aPUOo+LpXGo3c5ZzTJqua6ej/xCc+Sz
glmR+niH0OmeK0dVTGb5EycBZ0OL4pNdubegcHcPyGw2mYyCRD2VmA3RPNMVoWsFsiMHZcqoJMzB
kNlXzCSF/eGHTd9vcUb8TS2in8PlrL7Oo+JeNvW0yLM4JCkPm69YlMMuwBWJfAYTUWdHAhpdQd1F
p5JFrXUvtZkjfRuuvnuSVdyIu74OSjgOol4KeWF/ok3DCj/CzkGY7CwZf0Z/Zx+Vg7aHpVQBWXr6
c8wogtJGkYADaR1BwmrvpPsMGTFvrAZrxEnz241vmUz8nV0/FjqytimIZf3Na9cEOElh9A0WPOH/
yLX06zkzlStU2FIWjF0rkVujO5yS4GT3nqAza+RDmsgUW0k5MWuuq1LwGhoA0Z0M0a9thZijEnuv
hSdIMhdcauKJgeAC5TwFYEdmUy4CCSOzQvRbqm6j/uq7nvbUfwswmyabmJVrEnJGlB/RK2yHI3Fl
ep25QZMriuagiNnezStvI0KleixSVSvNVGboWflKXLwSbX65RgGWHQq1B2wc5Nv3Y0LAttZZlaiF
KjyQNUcWWFeysvh/wCdWPTbwDuG5+2/VEYdM9cxhkK/NFUpyHpG7G5JgaSv1NARAj/U/m6wM9e1k
c9Pr1YEGGgF9e4ezgB8acKvQ9CjmaLpFWooWqBRhqS6UyCOG+l3NyL6Lczr+xQgFWzEArDVfjJ1t
M9eSRcdGR2KmiHKKmzJ6/dA89p1FpHAim+SyvhU9VhXkD3TD4ojN/3POqbIVWP8T2vJUT9KbTKGO
hicQfuucWEYhPirVmY2pHVHD7LTBFLNaeABM9Uq66OkB96/xd3F0d50RrZR4d3Na2nBiR96qoT4/
/r3UfRZbQ2g8dQFYmpFA7XyZe2fOnafLg5pK67ldlU/FTzePsDG4Fu2B97kRCYhWbV76csDshnDP
B2CjRSG8BXGsua96HLZyEjMF6tdIQ9wbd+n+w+/H7Bwivh8Ig4Yfx7we3cijlPFvZja1Xh6flq+t
Jr22zW1Syk2I699PR8RwirAFJBKeGLsGla+SatoAJ5iuqwhD4k143hB4CLtseltNiZ+SZM1F8R9d
z/kTaeMiCLeSgfi/hKSRdh/Y13NJBWgttELW0vaRrDAqa+R6KdDBIqJuHXd45dZmgaMhKiBO0u/h
KUoPiZ1Ifxrfrrp3Mj4k9csNgor6+ePSFzWU8ctCCSDL3C8oWNSpYFWOy2BF6TC9xgO9GZjyBqgl
bFfP2q2yMhba1rqTpkfqnymPuKA7NRCI6C+QejodLBHXqnHzVBsv5Rs0o4wmhWH3Ix+EMcKqMukO
L+xVomxRSUZdREvsF7HNMZQauPv+4pHlz4ePqWHiCJwTOljje6scuDAFDExOWXMBuGylW35uDkJB
lFc+nT1oqn0xCDpPJPQwDvqPvjESXH4vz82Ph03iXHng0XE75I0UhoCKMBMd1kR7wXhToxJ0OY9o
uCCacDmxEsG0AMI2leds0fbvv4rF7i/bH2C74U/3y7JYwCFA2NCqaVIBBgdZrwz0sHoeh0HHGJeI
kM/V/3lWfuigxe912jkWU1DGktOO652Hvs+wkjlCOc3f5GnuT7Vgr32X+llQ/+TuYieVxISP4kEW
E1KciZrm24mAELV4trsNpRIQa8bGv+EOwEw6nhJZOSATKRc120G1TJO3GwvFWFwGDWMhf0CeioJ4
9lUiAayu2rRammcbMFqSb7Grzfa5wjMXCJP6dKJySLAc90jrdExLAaEk3ZBbhYU/hwlRfkEl5Kj/
R9BNId5UzHAFfcbmL4mMYsasFSThVOOFgGgYeopIcqAR3q++xyWLrkImPF1Gy2Z62M/y4DrBixKO
pwpCp3uKuoWvoKEA1+Q1DvZ3XpiLN7K1M4jokWJpAgKj+33Xl5XtXkGVGBse1rIcSIGGcimTPSwQ
6h3k9SqSn0HtJigNiDkNcU9GXkjgxYOa5Vj6CnVe/54NTn5jMNKv6MdrNiqBinxRM0vn46Ctzp+E
B2PA75/ql6caEuqQLpkAmraviOeFgV41MhVJSejYq5QGjQ3OZEAaiyLw7CqjykAOMefhc5m4Mhpl
G6LJ7oHc361FnZn+0XcZM6DZecU5QWcQc5ECuW7Q8E9SpHSI4GtAdqQbQowOOQQ+cIkjZIFo0Ul3
hhbA4iLmpsLjpZAB+02UTezyr0W9e/n/SCLaXdetz0uIygDbVVRxkIiyPM8puctqhpLX8iRGLZxx
0OYqACtp5tHLiwFlEIj5Whm/s3eSztiVrtGyHACyH7FthF8cv8+sZpoXbv/9qT9qMnPWPy+SL0cc
q4JY6p3ek+iAD4m3Htv3bkr8lB+Oklq2gWSDG32ZZJ2vOj2Y4ApDjnPtHgpHlSIVOWpmdDe1caAM
XYIQ26kh6QyI/v/usgvSxwF5CxdYqhc5BbLKA1GdLSGNCYWQjTVEfWiRDcdAuzoOyMV124J0bVhz
dOnck+j958y40e2urGv/jzfCc1inJE5miWoPHSkeJuwl1Tvaaw8ZpgzvlVF4dH4VOFHLlSI/JT/J
FW4szTIYz1niK/v8+iuA1Nkt78wZNG+qmpchUCFfsTcVXJ9zq915cCW6Q9nGyzIMSk7XHe27SkxG
g5smLUMErMO+dnF+eWK/zFT7oo6fksrUiPMh2C42Odi3JO66MY+HJM7c/gLODOT7bZ8d73kUR3CT
2l1KDOXGNHYoZ1NSX9g2uLhUJB1RNQmVJXWzeKFsK9Emsgj1oYmaa+s2HRCpM/Gph9GXNq1s0Qyb
Wmbf1W4MRtL7vuIq6/ev5tpS8lRW8S0pPS784gB0llx5qtWnrK752Wc03MDLfcyb+8he417p3ILF
32A8mnLpSH1sZNQ3/i6+iWV51jTwWHuaiTyC4mXU3Zedn5WoT1lyzxuRQhiXRgr3m88dJV3NtWzn
UV+8Zbed1ASVSTB/whDA3+wS73By5lWG+FIR5xskjdGfqswlNicP0Ju6lLplokFbHiWGrQtQIKeC
WD1aNNdYYwrGCe/ozkz2mEObalzTWw6QGvWl3uqSStVmJ7k/pvuf4CibPGpfGBXtye6UMhezSCSv
mvrYkZs+DNJQCt6VyX/KVtOzbvSbqemsQDjF0uZkRm0xtd5caZMFlSS2DJv0gqi4GwK54E7LvG2t
tWCzhwQBYf/l3H5llQO4dVSlNvCHgxRp4HVfwpv2kdF9xrM06pw36NjnEGtfhAmCQzWHwWRavbGe
zzFx7G38BwS4JzLAjtQXwk0UxtE2bw5Kiuno//j28+2AQaeKOdKD2076ZS43HVqUz78orEN4Sw4u
jCFRoKZyFpQfQMLzU6UulHdQ+IHM1ikcNutTKqTbU//zErN53Z6HX+WO9Vpa2pp9UG6fSXYybkUZ
EMPt8CmPx/lw0R/n9Gse9Nb9e9KTEc3vimcL4/bKnQTbXQwaTALjBTBYc9SVECzRrIwSPs9hVida
ZJqJHdkm5aUinAm5Y0PUpMHBbBjjR0pJp39vS6VRLTmrliXpJXqU/zHKMpu/rTohgeInY7j1bDTk
hWt4i+TASl/A1SGug9gyEGZ5AZUv3R+vL9eDR9TLHDyZ+QqCF9BEXaxDNHSUfEF6PpQz47fFGUzh
TFSP5oDZx11Nepvr3pCoBhFJ+3cEkG04mai+CklM7gWFkyBBtk9I1etFwuvHmvEZmJgW+e5CtkMm
Q2PI12hx3UDEVOMDehJ78Foou2ykmJkufQpjZUv8N424IR5ya+RCEMp06S5WfXilYxYCjxBFdYpT
bJCi5Wq/SiMdMcs2FYhfHqH1bQxmgBDfTtbX4XwrskXYoOnFNvgD5bL9NYvCACUzfzGgRjlZlddP
3t9dxGimlnRIU6EJiZhMhl0crK5uqzJfWve4R4SIgYF1nyfC1O8kknN0bd7JR+6I5IbodNODs9dm
m7+rLuZ2i0hjzhEh6v3G8twxiRHzJCVhK9Fjqtwl74hXIXhNYWB0lervj0+RevweZUvU2xp8fozd
F/LunMOW5zmb20iijGdKfrbk8SA0AlosWt1QBYiDPiqFQN4LxuBdNxaSLFj3oNkrOsilI1FzPxlH
rBWgPjSBvMURmZSCP3uhWYE/KHVBs3mRPvtcamymsFjdYl1J4O2Auwd8BB9x633LLvfB15Ddp8G+
xumLZ0PG5oxSL5TmFh0x8AZweF7VAH7pxvzmGge8JhoFBvnWMyDsXfwAV9FVHgh5FlDtXxztkbs6
xPZSKIylc+hmkAgpVHsUccFE2oZremtEAtHBpEVIWDdNx3FB05ltV/cby2/ybeT6lNi7XVyOLzp/
eKn89kz7u3nkRFgzjKdINLkrG//UmqdrNnF6/TET+Av9NM9S63LUIXVrM115DpvViih4irS9fqp/
R9gANxf1+/yZ+eEIkCsqJxliDhNtoBAe7chI9ECj22JCCk6JKRt8scOXfEyOeroGS8R905VJoI27
6vsT/JfQ5T8Lo2lbEl6bCzrLfxl7vI2GBurt9t2vCwHhrhzc7LxIf/ksXjjlOU18yokj9kPeHhfJ
FdXcMRNZEqVb3+RHK0uUQRIUCJCtAmNDIT2sqd9ib95/CtgPytXUBHhXn1ItKxE8a45OEpdjAmMb
wNINvSpl6Hb/PAhfZgaVvkaF9RG/m7HTcogEjK3DIDtJe5n916UduTM7RvMkwmRrPAHcThuV2QyU
EWcS/Vb68BDqPl+0n1ipI/v+4fIDJEv+ubg9r5nA+WS1yQUgIz8E0P6nncSXlW2W3R3isuI34Otb
wXj5mudRQFLDZ9OWSlqzXTgpr4TZIS2duolGfOQ0DnrVJH/uk4tkk3S1cxZUzaUeupeTXEy1dyEf
jyAnjcxY/KX56s4cESI5h1buCY1QRUHzNsx9c1xM/1JvW4mJg0pmOz6j1SqUQx2BMo5pC4iTY/Sz
N9ejB1B0+Kub1DSZx6jGwka3xacDlmLRViqBLjBYLvvePoi/V9aVo63A272nGcBtcb6v5YDlQmBa
Sp8NBwzjDfwuxbUmWZB11Xr7r5joQVEqUY+qkn+f2gb63BIsNQox29lU+79uyqglGlEbmVPVnqDB
J/JP4MHn1LcfGlndAxppfdPgQtFP11wuJCBrqGN1IO7sF15AIqZuEYiyIXM7fsRSkIRwgbHeFc+W
wnPLBpVKmxm/m5Tl/czJ66R2VXOFBUjqGxUk6cFTfRSiqJQuoFNkVv+URk+x58ghMCb6/nKw/F9a
+Iroe6Wllk284iDResYV0g7DJj/h80rVLEXa/2hFKXhrVwv0s4cpr0HiqabcYfg0BGcMESHedKmi
IL/1mI3namAzPWTXHuRZABT1vLiAFl8+zE3zW0vvxWE0bKowl48peKnG31vCbL/msJ62PNAYBxza
a7X9IHChjpbPwkxeAtaAEr77alf1/xX4p5rzXs/7BjYQUSDTLkjQXgV6iPjbf4CF7jRftw1X8GaF
/NjJ3LqXHnF3fLNCuMwDikvNnHgq7XzATbfCnG2xI0Dfwd1/Go+FGUKNicD4G45vptxZrahVSrq7
H2QNM5JbqM1I6S1dbhfjhxy/uH8XXUqFXkhlgVn/NQEllridY7Ii9nsChrXO6H+++o6Zj8eX12Ue
3oqheW/cFZ8FnksZ5MVUGYxmzd8rU0JMRaxddYxEOF9sXZoV16eJrmoUKE6RzoAgufrhebE12lUj
HcCfYipiEZtW2qciXXt5oRjKwbLYN59JGgLMPXlQIt4lAEyKzohwdtNMGpZVBVsfK9RJQ8W70Ur1
MZz22iItuc55hyIgik+CYCdpg93ARCqRDfszdSLLZnbgetHkttvPfDVvo9Hir9/X4p4UP1aJDNoz
usgWipt5+/1W5ABWSJwIzjtrkbyL/tRgAx9PYo4zCnea0MgzBSYwcDe7stmPR+fn2z1U6pH/5ohK
t40HELxRS9V/63XO/lHa0ed8Ggb5+ftBF3IYIQgXxu8SYA97dhepuDVfuyClBPXxcQtz37M/W4eZ
vuL0dYTxVL1h52eyRqI99HyB9WJfWc4sQ5txQ2CFVtc3gTLN9ZOJY/AmeR0Oc3cKYSlaIBrYLrTD
VWPwIgy6I6k5RSGgWvKJjrnSG2JXBTZHmXaDeJcPRoLcv4JYglJT9ilaNuBY7+pFBtCj/S+h2KAD
Gu9YmTDmC1Zh2rMR2ca+36B/9VZ9e0A74hW32Kt1w/J8RQWWuT2e9EPmfE23iMwxp/rYTrJdNiJ3
QbDloDGhxaCuVQt6H3ZHHHNWIX2O0PCLCxeFkrkQ+sm8aGCGaZV45isROBUIjvtwcmw0u7Q9tZAC
+7PtFwsQUlwdZnm/iAbIzuNLGD+3I/zG5TmulusFiccKElMaIndjegLshxgJcMy+QE2OofvOTQ6L
GdXb1b1Z/QKaJ2CvR8Fb1yxFTQUhrR/XmpdO3pmShQqK7yWnPUjouF1tODKH9mBYmxVosPpRVQGr
2JJu1zpz/mcYGrBJDIidScUXANGTHacm0uBVQjlqQGpvjT51TahPrl40YpZKImGeZJ8Z0iy/HO5O
abJDe2UiGSbN+VTZLn8ryvmivwtm9zq7uMuDY35i2PFa7GpF73hDq/9cxHsVm4T22d9qXeSjf68u
vGWS8lNUqHncOAMNDpXWqt2kgKrN5KR61x2J1xLARWSXNdNUBf7iHYT2AnGfLpAmHubzZmes2fJy
afD48QNmzLCCauFaePWvV7aFkV78KNqnEuddvY5zcrz/tvnatpp8KDWNrXE/bwbx6dEhFPph0mzT
u+Aehp0oRSmeYM77hu45COnz5DEzpUZJxI8tGQerk99DM6h2IlVv+3tSuOcP12ZC/6ZXIj+WMKiR
VdM5/4cO8iQsjCyddc3hO8i6l139ULvBqJtXsy9SutzHGErca1rZeAeK/yctt3JBu/kAeBjJkM5N
gu/tqO9QiOaEydaIOP7RXyJaZ8tVFLlI5YRYFgXbtHM76h7l16JK6k15+fUOpsgHum8TJkIukY8M
lDlrb/V9ZdYmC7yBEtG4IBiZhS7+kCTXyTjMZba65dlo433Tt3J2jjXQ6KMDRM8DCFgwjQ6FW6RC
NXv2Ba/iHP0/HTe9TEJ3QZ3c3UwSqEgghO+UvUVdPOjV5f0lqxji7Bn4osO6TkaaqRXGMnyN2blh
PvJs8zjaGnwMyxyyDi95K1D7Pw9k409ZUDT2wENn8tmyGGjrG3VVULESM0u9g94FKMHzuqJPGN82
Uzg9WK+aRXeR0FRhgXRhNZtkhWOlmxehaiMnsA70Mkt5hDTZgCIsm71P5kWGDWA5KxZp99omgTRQ
BeDqp2t377QtSIY7nNsUc7plXedOF5IgxvpVkjYsY4zAHVIE58nb5UTa/O/HhbipO/5WyZXEvthQ
0R+tfuo59o48dJ0ulqZWITiGlH8NooYiovCodiWBtpSJ8ZN12Eq85/LtPPVRPZREUfVA1aGeDkDd
tN378QAYzzfmWNcqaZ8ri341jpBYRF9a5KvmJEPStJs5Eh0zQ+ivClGA+qaKRWBr6zC23gB011eY
aohN6WIHPb1wD4mfu5mNuOCq7/uWHbb7nWcbt3FwZlRgcfNK3AfwYosOYs6833HWKTNHq48RrN+y
hswr4rHSyGzUSwvDQe02Bk+PVfT64KbdHnOHDrJcxeXW90gopPzDrEYsAbP1hgeCP9XbkqErbuW2
XUxymbhOEpNC/z8UkR213vlA9ThpyOwh8kmexhiq2QwU+oXigIQKT92oJmSbIAUcLlluMJDHTGsU
FbUeG73ZhgSVwlOvh1yqgeGe63wwHWyIs6ha6Xx/T9KeMJklwQkCghOCpofCFD2agWQsty3EiJfp
bwWI9Hqj4UI29DgWfQF+qxdszvkzYDd/SCHt/8F0eqEOHrNDewOHfzvDh7pyMUWkmSzgfXyTrWIP
7UW7m5VAHTTQo2F/hWsGUS+tEBprTz2lknkW5puTsGwjdSRgpvLA4od6GhB12CAP7WIYb7pvEgfR
+VX/AFYDm4iOr8Q4aH9YjSGyPWpiIsOwAPKMTJxtD1ecULZoiTmAsQELya1RoIV2nPiCx59AjcBC
RzGkMqtxun084QFZGxxdF//LSElp1kFBlcfyT85IYEy4PzU5cTWVqcmlvzXHsvEWzZXvm5BVJokd
noUA9H7f8SWT5FlJeSZJba4vZ0BwYBzeQhkLhp2lpu7u+tZLl/r6eJ9QtEd/A7xzx2ntbeBniqEd
08UzZpTIfDtleTYqjzLBy5LJYaH+6KUNuCYh0Kdxz6vtMlJKMahGDkaoj8WEIMkFxexKOnOVn9w3
qhjUGgCRNOXMlg2EAhfEbTLcG01cAKH7+/teqCmTuY2Vx8ueK9EOwr55p/C7zY2UAVjLlAythSjQ
4N2xMiP+kuK+hiAYRaTSu5n7961nac5FJ71yOlUEoc6lR2wJUf0ruYgtsqSf96rwJ2ObBJeXNMZu
ITufQJ13tmxLMSg1fUoe0cHf/0UeYWM3fG415v7DPLdbEXXNyZWrrUZo1B//kKIAhpITQUMbNWu+
D5IJFOiURBHRYFWrnMXJh8BSglJVW7wyoz2BT5t2hWp8yWFvJIZn+4Gq0eboEN69x7JeqdbS/dMX
HM2TKxEL/AUO5L6hDWYbwIcObA1WaEtdRd8OC/8pMVEyQ6dGxyh2dg9QKm+1aQy7jIg5/W7uU/5u
Oq46IUqzfreQxISdda1bgg5NuvIaMpxpgZnfa7sNQXBgkIIo6XlT18iCv3BSISHSnv3g/R+MKmkG
tdBy+OoXVuI6OmzLoRL5a8vh2Tu1Nh1Et5YaZN5sfS0qmGEP5ngMPyZopuq2lUaeJoG5+EXFZpt0
9lv7yGgefO7XWWZtLIvCc1BYbgmiMkbJIl+AHfswbTQYaLAUjGO/PZ4f2h7OfjiEJPZ7yH2hUdF6
pjE5SoFs/Mux6xl9FNNSgzTFbVxvL12LqMofIrljSMw6xLtgKE2kUC0nZLHo/MyU4jSDNEfRvNuB
6gXJHUQnvFjgGaIEr11/6JwMpGs6CGk3oqjxeGBPFNKna0Fu9hYREauNCzcqYiU3bCcm7V3sAOyZ
tBylDV3iCPhG3/ALIF2l3U/3Gd893oR9ESMGAk4NH1XehEOjXZ9zoV5RfkvN5spoUpvJfSaRhH1+
vidQrq/0lyNuPlORtpj4MEiWdi7G3QhFVTKpgYavC35cvJkBR6lz0I//9AqCJhmDf0i2t5h2GWEu
AP23/BVpOSaiqa6vwmXFPm1NOwHAvgB6aGQN+dQCgbWozaUbejxgnw4FNGS3ZMm2OjJz489U2Hce
9oC72zUK/mcb4E1dTYdhhFVWsgsmWH6u1yQHXphBQeWeAinPQiUN1ODdDv0SUMnNXyB5IwkxCmJL
CBDM4O2KNgWdSDkVbDorO/lSn7QYHadajd5rzDIaq6XeCACJrpn01TsKV6hWj+q46D9FgvHzNxch
Z1JnI2t8jCYsZGzjLh+1kgaS5JTbMHSqZDaeQGgThOpCBz04TOSBm7ybTh1qD3MvB5qGRI2eoPZn
3IrHhY/Eewgej3+xn8MOW5P3F30FJ1Bpe873LoZXidWDcY5Rfg22NXNiR2go+/YRMlCRh4TcTePR
FQZrO3RhQhOGSSLV6ParUt9uPAqYmOmx0lXnb8LxUF7vgcOY/gDCUPrGMou+lxImF5DYXQskSl85
qXdidf7BeDvEXRK6orc5h9xJiJjxkVdtlJUFumG4PPFIj728kSkbetvo75+9SsdOLgz3OdjU/EQI
PbY33JnRT0wecLugY7WvvN52v8JokCMfE75jq4Pjilomc/cWnE4WAfYu0lxH1w4Cokky4UczpISj
ydoGtdUs2Vud1ZZaaxRYXKHrMyoD0cqgOSUP+etSX9XY1cyU78q1rThoEq4jlLg2s82Jco1MNPQI
3ME/VnnsO1t3YoSFnBV+79ShDy73A9yVU6x6v1eSpELatoLS0/BFZHcOQ2wmgFkmV5JhEtv2A12G
Di7juleEsZ5S773QDSO2KxOrNrGof01m6UuuN939JC5z0lp7mvxiFhFE24rmadi/DB/OoJ8lPivC
3iSEidXFR1tvhB9vQqHsTwOJrN676s4TNv91U+2+v+ko6a/SnnXot9+RsZQVbk6R8l2otWroM5OT
3eTw77ux4tKmVXCeXnaKFvpmE72QdCdVgMFmFTKpBs5hEOENMT9t9xOJJuir7ncb5e+is0N0tO5T
3901Nt2laKtYwf0bNk7p1c29/8sJ8HtCaQBlE9sgfi2bSgTVgzxPTr0TNmzA8E3DO5SS7/3nqXx7
3lrV2/k4MshigJTp5ylT9gSBJioPA5l7wA7cb3aecoYVloCFdKyZSMh2n/3gk9Tv1G/450ChYUkC
6YG5tUXpzKiroe2+WpNPC/+nlyRUWKt1ou8v8SIKmNmx/5l0e8FO62A54sBaJYQ3TRfgNkj7O38H
AvtfoLYXhXo1ZrYeImP1IAs2WOFXu8AJLxVwWVKFv/RaxoK/ldOSdJ3nbiUmwj03zBbtXoWzZrbG
62l5A2QYpSDFesvsb3MX2gvCjgzhbG5YwHjGxlI0S9UMda+FWQWG9rgJDfg9jP1VyAxERiwQvK0V
Wfz5dnn/9lgvWSzVamHqmhQZ97x6IeOEV70PMcYFpCewiObZYwWtz+QU2t5Gut0O5qGGEg8lCWhY
IHbW2IiBPO8QGcmyeLRW2g72h9owKIYRwdRr+q4ncC4jvz2T/B4VKQix5kzI1BNV3EV1tDeIBigv
zkBDsd3Q6gFOBKBWbKOVctUHSTxtMwNM5XIxnT2xTQHQSsmx0Mu2rrSy53LYT7ZpNoG/YJHdgrAy
928z9N38S0E+iaWCQrwEArJiwbwCThKU1roLdf0aXpXYjLcwqXl2bo89HvubG3MSxEDdIVhUuHRd
m2SmvVpNk+cg5s8ua6b6HHHkKGMWs5Y/QrBVZirXiZPQqX1ka6hMeIv81kp6SrJoenZj8AH7sLam
HaIq/KQ/77jQWMvURruiSFgwXbcgY9wIuedZ6A9A/s6DTRRYlvES7jgRuaCWCBQ62BpTIAUiLXc1
5JHJyxyfkymgJbEeJfJkeLL/Kg7yvxdidfwHhHCVePyXED2YF+wTAZhlkXMcgtu9kVHvxaFDQU+b
V1LFHcHPjwegFdcu6RLQEoHwMfQk+Sov5qzzLi9DdQsIq6JmJEYiemr4VT5kSpqW9zmf5qc7FJpO
52drVRD4b4v5zHm2PCoUqGNtHbK/K9UkA5LMmP4WBFQB2GkO3AaC4NbqdACcEhSXAHXeNKUjYgfq
G/Hb3AwpT1E3p/Ss4sYNdrrR2fSRPrLZ46ENNVLI+LGa39wBeXOwVVMyK2fZW49jl9djzMhzvQbw
lAmTetTjezCIk8WRL72hMU+SmHwkfz8n1+Q0iglqbyNa9gIw9R8FX63fy4GFG8B2gCg47cfHj72V
7qk60LYyzVb5VWz1YkNFv2FXU3SFJuSoqOyKwaMByYt+hHssdtRglGjli/yjWa9WTVjIzmxAOHBq
EjHgYd5EkGtx6N04bjkTm5hVFBtfzUrPCj17EIsst2hKGdFRFTfuBJFnJU0vpBiXqnhj/n4qwS4J
jyIo2C9wwz3V4Xud4wOAPsncVERGEh/twSaQ8SFvO14JJEPkME8zIuSrobtANvka1xnoSfIQLaZo
1ON3VG70KvcLlzK0vssyl8vK3rn6xvvqIP/tskNEZJ7ZNmzOM947D7vKZ0km5qp0w9DVKMQx02YQ
lljVLZ0xbwgBpcn9H6Xe9N8+PCVG5c5Qe8/n/Q5sg1PBf1XmPikEFS8s9qfbOh7WfKygzcf+0Czs
CVH6XvQHRWmFYpBU+epROsmtmYwsIZT155/VYmeEVC+PjR4AF5c58bIFCffwCtUFtUxzJJL+rRdG
aGSGIpchEcNIs7jzkKCddqNocU2ML/d4itg3R9DzxhAwjfvpJ9JCCh5om4MB01srbufoRxHB8vsz
jAI7ctw4cDaLLj23u9whTrrgLhIrJz0f6UOhoZRbgO0vm8g9qulCOGKwzUJyA6wAT+ZN3KywyXfS
NAo8sxkqFdU+F6t1ssvSBou6WkmoQBK5z6ivlpADaTScmIfdWVaIfXZJL7lvUfwMtrOIB+NhqJ6N
xpa5yj/WhtQ9Bly/qErVDCX+Do2VEEIbzNjF47M8nY3xE+Yc+vjEUeY1GrCvJDk90BNjpS/qxzAs
D3iurj3sTdEbHSFpjncL1HTW4Xbz3q4TP3RnLMcG7BpfkqJf4c/8T0GvehJFYB6i0/qqvlgJO4gU
z7whTd+WTfz4WdQgZYrBdwFs6r6T8eatbxhDIvzElnJrbGfYGIeqtjg04MUuk8K6zFHuyCEUnPTs
fDsyYCtHGhwWHFZKinq772sO3UU5jzabT/mZeyKY+azVQpwyU3QXlAvmOsIrmsF9wWQwbzf8i8xm
L2qnm5WHs7jVZ+xKDx1zg2coHUI0NZLyTHVsG4AL3ndRGi6jca0yaBBoXBc/nLOalY7Kb44xuoh4
2qBNmY9XSt2WNkg2U1gOjKt4KyTgUlr2F0QuxbL2o8OOYzvQ7JJ6XiPTHDEavafY1MVHoA2Rgw6j
Ip7CZplIvhtV8yNdyIWzE4CjHc+r3vAuLdY1n+GCyC49jYsw0/DUrqCwG8lMuAL1BAOwFPF/X9w1
MpEba98E8mzBpGkMsqwf9NJP5dOIWe5oHf9bx0VKM2JhL3DX3kETIL+nPFiaOQAFOdRD0pGaPdVM
AyoLOD8ouA3X/A6xslwQjp3aJOc5PJYniOQtB6G5hftfenrx1OnCXj+b9IsIHxkkMgcQ2HpWWMnU
rp9SZtD8AWo9Sj1a3/RzQGFjknX+Tse5W01fpqzVsKXjDWkB4sE+1kJeBs6MmOxhOvv0aqOfZFtk
pJRXqirOGqsVHM9e0ONG3VaB43vbZaGucnm/mPrdo/uhrBWkhlK0N2afpaXIFZGSoLauoYicQFeT
wAw55t1OiI9WomdJDeZ02NfytVunNBtwD8dAPbsI8Se14Y1S+1xxIqFdFZNPrhS0PeDYUnt2xoeR
/hX8Fw11fop9nyhzatfQzNwrr5/awqIy1nB5F2w5xQbFV4v4rXCKggHC+CSdl41eko6plOPUL2lj
iZs5haIiIT08ZAdQ7RtGLW50I+ERabK/4o2FbUZyKrooO/2YU1pE6YBv0qyYkHvCr/APM/ZFAlZy
RQ+pI3roAAYKeBA9zR9H+E+rkwAlzDXeEaWxvexVig7h/Y4BEpYpmyopgHrVXRAke5V0RHCyMmMa
ce4w7m70Q2fmHBQ6PzrIZSXBYeQl1RZ3EYE6biwX9Agtap91IT+if2SfRDcaOHHaQsW4O6/3sQO+
0orvQ6zwSomdNWhRj0RY+/hGvDwK1TX3olHdkEfBBfOfAH/DNZGwSb2E41YH5yi11d1irNns4ZV7
2jNqrRAAMTygApUvzWmoPiLKEHG9+57ucuCRJvJJliZLswopFh9hKiYBD2/SB+CULZakh+1j10FV
cR8d3gYAlXXbUpDsXRsKDAvxDYqTSGTqtQ/TLXASP1F6iQst3qBiSwruPLvZ2pTTK146S/Y9l5Rj
+fvaOlP+VTvU8JzO5728+9Kq6CIjSGxgztSJ5Una+6CbKn8Et98CS4qwULlnswYY+V2z5Ul1CWKs
vcoxDn+gEWQt9gNVClYgvUMituKgw7mWD0dLuI/UWgxXAUMUvSGi3P+CatWR1bprn2YtAlMCMY+L
zs66NVwtwkCRtozsnN/hNxxF1rVC9/N7UMGkwlP++eL78WPOtYNE5qpDclGHrL8CzPb4fScI7ASu
1SSMhg3LPdGPMbDXDkUdqhliycp/g5VFjho1N3ZY/jnKE5ACvboBNPH0aiihHvDcSBFjswadmqUL
hCa1KCKWu2tov2OLz0ndvOa9/o4N9YAxhlCA+Xg7Gm48dw4Wc0ajtpHlzwHKTECIQvP0e/HpEKjs
VLmYKPANUDSA9iNVwTk4BPfznHvcbhipH6C/zCr0sVH0EVqz5seZMuOowVWO/xGyPnAfQ6tSSdiQ
wPIN9cHDJ6U2fym7QhCDfhFvGqAOZAF0aoNxeZUuAspCOXDByJRi58wFLHGskVx5dYlsi7assi9T
aq6u09I51J59ddDdHxhfAbFnwD7Uv8Ibq7GqwXxgtwFZd7nt8K4agSdHzgOhk6dC69yu8bRNCegr
JXQ2yEBhTPnVC0Ai54C16zACmenkd3LYvZ51ZioYLugLtR5G5Sc8Vp9ptcLG6/V8n83Qov26nJX1
wuO7tWpVhlNhyxOoFDGta9vw93f5//IuJLHlG5HZ2rQJjLloH2jGTuM1Ddqy/gDLtb3aizQUHWTL
AuViAl1dV6anyz6PmlKobTupuj9ywKdYM4/hjP2OgunyS2Vjh+6sPKfwooH/2KEgmGhs29duoTco
6oU1yNSTuukdJ3YFbbWdm+v4JNFRSp8FtVBS9C/k2G/bLx5pQcCZ8xIYDetvypHz3tIMcs89NlPf
uXy6jw1qH1MOwibktmk1DIwakLKw8rxUdb+VfNJLC+gHs5jugR8SeY2UGYdSaZzDMlCyKPSsMkUz
WYR53L3nM1E2lJfB4J6UE3BBh8ZENhiLA50Kh92Zgsk1mTWXBdM2akUwRPW30dJL8L6lFuLCUN6w
THDFOlM1HJolSGEx+yqlJ0rcX3kdR/yS1cjHTN4TBEQ7wg8DK5jP2Lp19qkcsCKc7x1FFMTBQIt8
WhjwPoEvNgbOwwsxAPkupACc4oe6G3VreIPpocT7MLQ8Eq5mjndC5vtmv4f//mTl8dAhhm+CTU97
5+l1l6VVwRYxolXy/SFFAvw9U1ehiV/4KNNdTQeqepiM7UiuprZYAuW5pq5L9FK5C6SrX3tFGFbt
GuHqdXbngGxHWzqurT66iIdzoiJXf5X3ut1VE4wFYT116IS49JE2qDjlIhbSTBQd+e5I5VW28aA2
tGskvcYxsV4GK6vDFQk1FUVB/M7ZkqMpxirBH5E2sP+Fox1D9lAt1yWS0TSY+JKwOfGCbnM6lDAW
Mi073cm7TeRseX7O+E5Znr0qLujdQ4eqm7vbC9H0ERvuITrij6I5cK9R2KEQor5ySLtiRb5/cEuL
edoDTbDafTcI38U6fynKxLgGhX9Jz1Tg2NN9D67qGjTjmBYHm7kapAPoE+KDuhBdcB092uOL2PjH
qxG9VZpdJmB3RAky0XUvo06JGFtTZaCWrSvzSBbgmaVxQ+Wuktfpr581MY+GWbPn+0fE/pNMKoks
e+zo3+vBZxIQTJV1hJjqdsc6x7n93CGpEX8/htGa7pqHUs6Uocyx00Fm7xSkZ8mIYUd6EMM+MKGj
srhpBiHu7/IILO2UVdm70Iy1/JPeCka2aAJDk3UJkd58PWmtOuXFIPQqPe82Bp6ZZNNMQNpd/bHG
BOrr4bmqttpvWGlf1CjCpgAj0TLWOOOXa3RsR1oWShx97kN5Z9Qe8lwYF1L3w9Ahzzu8tPhR0cxN
Gma0hnZWcZvBM5k7LQlnDIz99bP+CMJp1wun0Qr+ubLklgRl8Yws9cqGgXi96/gTICVpU1XfXIez
LoaKU1cVC2cyIXmtMwUk9c0XJZy8oiVgr4ZmhmjCF0neVkysGxscf5hqinppiibWBDK8z87jE9ke
xREsq8YfXk/jxQGMJIADqnMKyyOsr3wxJ59BdU5Aci5IZEujZBJtj9BVji1viw40OKAPUH63JgJ9
ysc6TCg+M+K9slbOr1xzv9IJSrUSJSRyPEPDrZWVK3/3b4G15tmG5Ast5uT7q/ZadpwYiPQ5xuP6
aohPBCmFfwmF+uxnnSPQMoitcmq90H7CntTMU+m6kVySBVaBjz4mchWcW+fnBBqaa7cfGRgABV5k
8dTBv0yjF8fJm97JpizWCTRb20lQ45Rxelpe1VBtL5Q5nH/sgZCsazw7nz/yoCfrSsGmp9T5peVV
CEQSayezwUMkg3rTBY0XNAGKvCS+vDJ+1ziGcMGDv+3EbnwrKcD8Jb3XrZD9AMeFv6WuNlkKOSoC
CfsIe5B8G+VYVFtP4zO6/PjCvjXOiWs/V6ynsjqxHIYBCuIC6imGGqqGoSVr6OtaxMVYp+VheSun
i5ES1NtNx6cmS5MkYslF7H033KlHS564LMNxztz1VhIRnTQ5p32yEN/sc8qCRm6qsnoMmRk0kfUL
7HAiExt608bkmvO/4Q2Py+K/z52oiWhhdAyNUhkAceLKxWuwh8wRtKwRyN8fbpSLETsvTvYdQLKc
ym6B9oNCmbACJaGHCRYUgfkvdW1eIaIIsDgvSM/WTgfiXcFBYSpi0p7+Ilk+EoY9bnEvF+RmKIs9
1P9MmMdpI6szNkZTNcGmFKQf1kSUi4OeEA2wGP3iRPq6MeSrAd+xgyr4ocZc2kn/IKHFbdE6tu99
Klff65ZbplcDI82iaFDCOP3gbuw8jHy8gY0cxcHoX2HDLbtJ6H+pW1fUx/KigveXEpOGnlublDbH
HkqRH8yfxjH60bmv7LxsPDSBYDofnjA1a5z/MmD4+YBAZecurO+ozie3lJAtsFbMPy9DGS76cQjQ
Gison5vySxoJCC9b6fqwh+9UZYopuUYVxRC4bHNZ3njt5v3M4UQymMX1nKxk95103TdKHW+wR/EV
5NWOIoY++sdcF8C8Ral6HoXhYRD7q6rnx5c9YTGrQfpRi+CqifB6TDAqZHc+EoJ+lCwHY1X9zO+Z
AZb7jnpMGDOPltfp8zdHe8CMv4BZu8RTpWs1qG/NX3LK3PSQzI+Znw0LHRQL81rSkb5ZX1Qad+7e
+/CpByJNtbbYsHLrDM5Tiu25hqBiU2TJTy4PHaZpkJTZdB+s9q7ODJWbdBCaxOzPNbZpUgaQ0A5J
D9t0gqIkykSvfF0kM84HnP27Nc8z7JskH3BvonfIzJ/yZSpdcDL3XMf4esD9U5lFWzH8+aDLoxbq
d3RTLlRw0Yf7rOmmciC1d3AuIyZ2QVZH1TE9jpmYI9jDVoLv95g4smTPZ3n5rvIJidi4goXXGCgZ
ZJB/zhR44V9aG6s8Vh5HXR7b0UNMP78NsARWViEMG2FYDoj2TlK+OkSd6iscjQdQ1ttWnsepTjfU
ulnEDq2ylbGHV8PXVOr1J1IoeXf5+TZ8K5ssSQscBRkzVLEH44u1rikB1jmmkZZio6YEdk7gg5ea
DWtEBuOXrorIdv0XdkXigJhEvmT9bXiTo5XsTK+evwR9gQS/ZB1jcr8bvQQeFWK05Z82M0eiEC8Z
oCTfBAlNpAXjLb25DvJ295Jv21Hw+oWxPKDinz4GPtFermY1sEQ3POAGXOuoCGsEShLQqjwEo1CM
geUDP7n4NpMZOyZyYTwpuyPJ4KAXDW96XlpdCd1OmEFOCOY9S+a9RgSfJXmENhBYW/ecObaF80Mi
PkfKlktOkxmBQo85BMvYa0B2JjLPpaOueTuLcyph3xIdpqz1EVBfjfKnGogKbMCKU6DEyszxIcCN
A/Lyy9ssh6vRSFqCnvwSCDJYEbjyy06R/QjyDSI9sZjlTqDHx6H+CL3Z50HtBxHTFz9t/Vnw2uUg
D6/IRao7UJN8k9Bm6eehIpo8c/UP1xz0SINVzERVgvhxEFEMcyso3/s3LCXYk1Q9ME0sLThhGb9r
Vwlr7sK6Uz7Q2yZMB2qUMCYgLnCNKiwjKMmfYlf6W46ylQfjn29KPdNH9bpptFqyTRlKsXhDFlgq
eGA/expqWpMtbhkbDM8A0lfmbWFqa3g8jHjrRIwkHCsLXYZzXPmZXYEYYCuoQwD+gy/2i0kG7cHu
xl+WQwcPnGOdS1FIt83sp94Ill4vVxUjYhoLc2a3VZ3rmclszOYvHOy5GZ7PlLNUkbXooEQrGjGp
btPGyxy03quQ8yPXq98V+tam6FdzAnmBtdJsicT/1LAdGJ/She8MhsMjtWA4I7VUF/09q7GrARRp
JUEbsweMQNMO7i2RLAfHWRBSOWvmZErGp4Pab7H3qwitQVkFVAPwIpJZ+Ah8wHY48NkO2IUCv7cu
BJG5zWQhmk9dTffptokKD+NToYW5SRdqKJExjUwTVNJb8MLm7f6UWv/S/85MOSlBlz9FenFy2NAH
CEUU2JK/Nq+vfKhp9xI/wkHy+QppVUe9ATUnaK9+5CYYWiJS1i9ISeXxjXZmgenYNKB8vatoIDc8
zHgdpOGxOZCYuII8ftwDVJw1snSG4VPQ0C9mr4947FERSV/PFlCMCJ1ICYoEgcxbiEqcIXD3V3aN
uasTPou9GDHo5kh9L8RKGghaxGwqcYcK6WBqZKtm8c03vhDt1wGDTguI9NPqTHX7mvIqvV3YlEBy
fKvunEAvlIV5OdrKeeeqALsu3xqS+jw3YQvccJiJPSLJDCj150TUn9RYweXezNTMyw/Axswsor81
+T6Y5w1VIdQRjvPpAeTYGvjPZs5tMnGzyaCPJj4HtdY7g4XmvzLgts4Z+hILyHz4baAp9iN9onuK
vYfaMX4DR22dbiLFaweNAqzg4ys/+yQpDeOgrtd4/vyk7AZuHEmzkft0aHB7YQepvc63cOXPMuH/
6+ZjWFQODvHach/tSc8rkTQIqiC10C2tgC9OTY1nxMqsnFCjWXSRHaJrygj8OI+Lo/QSdWidug66
f6dG/iu2g18zP9WE/aAw7SKFpdBfgC+OrtwRAB99aYKrYmPOsNMUu4kKqfEMesUoIybfh2hShd+i
/BMl3tbeYp4ToKcH8TpMGZElM+llVdSMkm1K7ipzYWQA5AT5yJRUYoD3vBS3xFd1T5f7PvmZkhV1
XpWyp1dNhZ1FbDSJlyC20kbBtgK6SRb0oPpYwbM5lJHwoZxLBEB0i2pDQM4+KfQ8UjcJQKaktymr
1fM/0ChWMdrBY24IXs26/fMrc1WH/EmcXlhiMWPTgKkr3VIZg0BRqdGqhtDH8uA8C80GXCfYUVVU
4ctEUFK2mkA2WnBNYgZOb3E3hCDJfZq2ZHU2bJu/vX5v1qUSfLqsq2Ud1Z/+rFA/ZNRAGO2FH5pl
X3WRAxcQgtSjvllMkwbP+A/RjWaPIE9y0OVeFfzC1heCsVR//aKsiS3UCdUU9L/MxSl7RKqZX5xe
2+fH7uzl7kS7DhLMPlVtQf1mQwIhiQreirLr8NwN0nMhSqh4GC/C04raSECMXZokegjtT5NjlrXW
6YZHj3UTcHfLYb/cJ7y8vkrFzwMDac5xv6vzxokd9w3c2ZXOVOEa8NwmeIcV1DGWVLlpZrj+BDab
RypgyNLVIE+wiLeIKAPcgj2Vn/rlee6GckRhw3zmuLXjR1H9ykgyVQkajiX/XEEdJc3vENUin+El
xZejxp+7jxjKlynSapOHg6m+H6T04YUMysdnNfeG/oycepHG12+3py1dyIGpreGxJQRTiOd5kBy3
ESUUJZnKdOtn2XC54en/tENcImDJ/cDYHekGAKj7gVbqtcp8GEPllVEGexfkqzvQuf4nBL1jJoJS
2kQwqG1thXc1H8KikqZZpHEyLI8MXel6D4epVEd8Rpgp2Yx571MwHHARdjQHHkHpbXqSu9botllS
Y2VBIvskqXi68IlvZbwOb3X4cgR6+d6U5bLf2n8SImALE/IpvW0JjqdCfDhJ8G0sP0bAzyh+afEU
qUD8D3c3bDK9wDhFX8pqDumpWt+fys3FmMqYJoAlhuQ0fzjhVZVaPuLy04SRlzPis/Sp09kkOwpy
lNNVpwAs1v46BNHTOquigd7lrF5eyb07IHBZSEMrLqlVj4JUXYl3XS6AwqD28UyNH77iSuLgDfMa
x6Zs2xzSZ34N9LTVWtIyVAUgffUbqTUs1bcD3PE9BU/oO6LlKZ62plJrNvcaM9TYsbNxaVztESi/
pHUIjWox22/zzgw2+hkzfF+Y6mqZqMLf8nJgI4j7SF0E6pY5V0yQhQp1Z7lMF6farBZzHdKSX+h3
oVXWDsDV9Xsn0r8rpZaxmwS9n7pE8I3BYPVR5WTOLhF/sBoTbGK0udzrA/EPY5NUKTCIlBTqAvFl
WxVDZH79K6knNFOMJ3NxFdSMrUYWEoiedl1pOc6vRCpwOFL5KNEMufHBFBsMVtaAC4FzhZ0hj8vh
w1HVMXbhaFx4b0WyA9/pgPANjPqlWPXUdKqoQrS0zRH8dt9Mh9rnuFFY5xNAZjYUalzyMCSu2JCY
vI4jcgLIXeJInBFRzOTpc9jfMiwOyHVC40gKo27aYXIS7kQLr3CFxIsSuKEKJSDnR/+TL44kJkzJ
RvinVsOrn7xQDtaDEPYU7yiae6eROykK0+BKhqvdIsz3E6LyAYh4kyTeb74SDufGNw1+ny5UbZQ0
xZVKEHUQXvRENojN6SHV5Nb7kNm66VzQovUio66b6uVOy90brT/8QN7Q8PpTVCX2Mm/xogN117p0
PZoYkkWmMGKycrTXDBv/tb3lAeYqlYViVrTm/hiiWT5uH9aUF4Zt5nfkUbwJd1XdjLkfZq2IjZaB
oYx4dzhLoTEeDKg4dD7wNhQr6uU84D+dGpuEaEa87fkX4m3hXDARID0AIo8T2hcgPFZeav9V3eEY
J9GAv1XnjdjOkLw3ZutVDk+xAqvJY61tb+pURiSEVp7m7SMLrCm4ribE0PIDauc1M4rQsYVwmIoV
rxBHQWoA/5ZK8KmsJUT3i9k5fXdzNLJk/wCgVPLuJhuWrkiBVaymYfRqrHdglYEV4+vlw9igs7pV
hGPfP3BdN5G8cPOdNhhA8A19FSCRhcH+0SgbITJIKpnAUwXtViWHn4yesH57UdfOhdRKUlXV0C8N
f/Bzx6qbw6GoQa7M7EOdZkk3SJw6uQEzEGIewoihvFS/8kcFCW6LvVT3SUz1ReUFQhK9ezZY/Ixl
tomLTCHkZas8VuLMhagfoTJqNmgVTP+9x4JNJrJjJzQNtrgXqg2dsKVJy/IJHddEPh8Nc4r5nAS/
rNdXI+iF+x+tLS05midac4+bHkNebVEihMiWPMBzrG0zSOZVMmmFfIc3KUmx2frMB7nzU/KL/uVr
DPmvOCQWGrRIK/OKorxmBHlDl7Dd5wKbcVA0bcLhzeV7BPJuzXpHVZiPjVxZPjEw9B1L17fRn/iv
g5sorKvNftvkRmxAdHwtjte2duK6at1mThHNA2U5pIFJ1rHw3e69EFnbnroBScFUcoXdSVZQinPK
iSEHFHvHiyEkf2uWXDc9jJf3G9joHCKQlekw3x1yZCGyp5UlkyQY1jTTCXxxv1Nvp1wRriTOYhph
XE0C5397hT+huq/KQUFmOnZm+uW5aytreZPrKDZOPIwPIrhG7iEzU/3WZZF3TDz6tkp8Ijn8HLsb
wclpV0AOt89XBAWCipM5i+3O0JJ1GQd58kp9q7lGE973IDXOjx2T+CMhzK3wfJ0qX3LJv5qCmk2o
5OutLzOHaruaqtP5Uk7QDQlVK2TJzzfMZmB9cpQ0JGOh969K2PQfHhV6G9BZNKCZ++iHjBUVrOL6
4j3IAGgoWC2gANY74TgwlC5uWY/NPkMtwtpTnSkYbtPiFgl+M6mtJBEAb58zWyUjZM5pl7jKy6jO
dSiBhGkGwbCqtCZ20IdKuYmZQwP+iLksXpbd0uRvsHGVhHKJOo3qq1IkKf62YuXk0ZqUxfSycd1L
WCBklnt4m7f9/vAt+cNpio5HHLukAfENIHKUig4iqsjgXAAKlBTW//NEY9n4vI3J6ax13vsEyVn/
cEmxiImdH2NvIFifHYhxJoKXpcKLWXl8KQzv8S74HXQZmnHXl0FgRHXFtJ6Nz3K+oVqQPBx6XJgT
kK6mJV0EvOkMouRr3oYuK3VUeQFf2rW+oKTYN/byeeZ/NrG+JnT/DJxQFaA0TcfqQZXBjDq0b9o/
o7V5/3owkUw3CWUPW1jrrVlT3e3P90azxQYkNguUoq4BGm0//JTAn2xLJJyrmEd/u0XCu44Suu6s
oCbpuy8Yqr0PffAXLH3GOoK3NdxunO/my9WPAk2WGVdnk0UKWjIraycVr4VljdqVhmp34NmgmM0R
Het+Y/xn75MXEIzNFvtFqQq2JB9mCwbKD+GSyuYD3KsUhQUoBTikNatW93QE9oJbK8a6DG8hSiIl
/6rWzI1RYT9n+nU1XWUFoQGzeFRB5O3JuBIuqZlRA+5Oj34kmaRXgpMI9kqtYyEpd+iAc/R8GpeW
Ca/IMDoCX0xX/zzMkRToFr0mAKrcvWGiEyTWcH7yXgUyXz9+w7C96UYq2nrJI6F40nS6KOrpIzQz
Bk4Xg+ZqXHmcnr9Sr8ynyWv2A6yQ/iAMdQnCPbPNKwYAi8XJPuTUmPvXSwz8i9h9LIjfdlJ23sM8
HAKw2EmG2UnSxMbMZmdVqvVdqzg9rZFFwdnH27wHD02U1AaJsMkFK9s5bw16k9SghIMsqI2uhOWL
C+P+coRizylAfgATGy++ZJHXmf4wbZ8P/o9bG5DmZbpEBph1uef6EpLO584wjT+dN541w1NbxCyN
6NJSgju/iHHOXcyK1OWKUm759AB6XxYz56ktzz96ejDOj3/egyoJqGSl+Jo9VjvBzuvj8riH8szj
zVDjNbVW7XduJ/NgbfAO0+i/sxqR1Q3LRh6RLLDPzIiowEnRaRaNLycGwVTAAq5Hi0GpBjhQlbrC
AbG60SnHeTIe9HrKBxT+hIm0Hjs9c7vy0JVon+7R9KjuUTUci9cLyLYZrP+Mw0xRkxhXrvNLCCRE
CoRanuuPCEXGouG1iRqf75+yiQm/iokL8qEKJTbMpWvD0cVLWbAGC/7J53j+gjIaX9v6EVXENaSt
iw0Llq58wZPLDuB5SFxe6emFTEe/yNVHtdGcTuioigfHFiYNjfkYPArhZkKWLWGVfyJd3v5A33SW
f46gKfnr3bKtWqK8utIOF/QlT5g08Kmu8iMurzV3bUQIj5O7roRC7YwUJVJ4OH8uasplyOofB/RF
opUpc7owOYMC0yyt1JATI0U7j/y/h9f1dXl+JcSsW/qKwpVN213fGYnHHtHl8EAuzN1iruvN6kV8
s28gn4KS04C2S6BEtVZ6T8kWmtv8m/TyJ7oDhTFoJClXSAsHIPNGD3hAN9ljTMxrVKVS4lrsCBu8
Flzs2o7ZZ4WkMHGV5WnRSc36Bx8UzMNRcssiFiiRQZFztrOyW0je0V88sGThDMknBGeTVpF41+wi
t1vxC+jXpgkBimqZXYSiJ5KP1VQNiXvW8X8qakXznnAAjzoovYdccbz3Dgf1T2KxiB5n+62P61mr
g0By7zXVimEy3r80WClg6U4QxF35GFFTgFCV3oJAKZf76TR1oFSqmEporzG3Xc0dVNPyUfXxK0q4
v4dzgNjisd7/xOsYJPawsiwuHmAUXsxuda821AuRuQgxHuns7QB7iZc4Ks/CuIN1I4HPRjNF8y/g
VH+el/m/tVNP7jMTV4YW01yJ36NqeJ+ho6E+96d1GrGmmoGDkd7qFCh6M+J9WgmbrWUc173SNGgh
oHIXhCK0jQjB1PBDn86EeUIMk2H+P4Qf3RlMHqqdhUTzVNtIAGZGY0gwyRsQYLGaKZbF0Npb9DAu
zL8Yc9CkSZ1tz9DkC3Zbxp7wkYaaJUdL9mNP7txpIZU/Qv5XAmiRup3rErx0yFucE05sQJpF1C9U
pUGfV2Vt83TML14TlPDpCfVSU4zhHCSIZeBPXPxaQMjGxmuGuNNs1/3bdZRcI1T9rVYwiGTuD0KV
CaDBNAiK6sTDNNdzMohgzjvup0mfNEwMdPP5CwamRsnpncBuccVvDLh+hKbFnmZK3bFLRZN0FYo9
L9eu7D/VxQ1BI5naDcw3MCzfPdQ/xkcsP2trdRumllthK/DtzBEIH+xSHxASk9uAb8VZXji5fwII
XPbwXk8dv3XGTMOEnFdGXNek+FqGI9106xK+9oO2+t6+0/Pu33OC7dszW5RYI64Zutk8MbWtVAvn
1xYQLFGTMyvJBciPT6kdDGMksB2EIGTVMxXv7P/SYVa/yFPnyHzT7y1Tjaz7ykBkU9h7NsgOlRdm
0yB0aPNQfq7wK9wp6KNSuhgoO6dgnMpJ4Wx5cMQBC7Bwolu3hGsxYsZTIG8Bb5Saa7x68TmBljWy
nE4eCGcdznPsrprcyG1Vs15C8w4FtUGrCRPVHtcO4faJdVX7e6Oo49jP/f5uelPn/ApJoiMKzCYC
Y9kDwdgVTcfYVlx8iRP5ta1K7FUYkPPRCsiBEvODoO6YYCYBdoZxD49WJBAK3jhrqYomaKGB4+pA
bocMvNe3SrF9yuuiKMUR4zzcVj4WPRVqUQVxZX+KXkW3YWQnMyfu8YFkmA/ejXVk6CDLI0UqKAVt
xCdVr5GyddFx6uBK1NHvc2VTrTx5CVj8G+M+UR8jHDSPsJI7rjrUaEt8uJLIcqetWRHnVENTgDJz
nP/DiJZkEb2KvYAUE6eozVQyCSrLNStf8SgFv5S/935CNXRWY6DFqi2mbbqY4t+BJ/qwRGoAiCrX
ZLepyDlput+NLh7CXVeIz1QqnbqVU21ZuRO/xzLOPpHGknBPsiubYM+8Gd/Wb7QVhtEUVb+VX6oo
jBh+cjYW75wmcoQuQqorFo20lgIeyL6YG22UFfpIIGepgn+mFQp5HCFv4SpXa25JQCB73heYHY/D
tHDGThY5pIUUZfhvslQhzR+tiyt4ALvwTwZwSFbW6fwT6yZvNJdTd+6mQVdfpCGzm0tKIE7EIDSh
tYxDryg57+iohBxFISDiiHhxL0k2uC66pYmma9WHhhB+E7g/oN4gaIJhSWyqEu8VVAc5Nzqj9hZE
zKw7SnBZNlSPalNP5ZX/zzxyQjOF2bRGx85US9o8uO4lPH2L8KoFtHm4/shHfnP45sbE+mb3xFNL
I8jLjL4Y3L+pve7T1XUvdQxiZFJgqUXjMubqqwfbcRzbrBeuOjoTK25ZIia0OpUNZnMNsC6W7CT1
kqlGtxNSByQboXXA9O1xaKN2qvmYWJtQlrTfKicreOINnhpBjgovQLX+spL00FthKep9H+PpqHfZ
DxJKm1onBIw83g35EaBu9JLk8YeHCKhXgZ20va5x7yc4su/tcJxvg6J2PlRsqv5ms72VHvoeosD+
EX6T63jVKNiRb14PDBMYkgfLG3UjGGmECZPfLTd80CqipVNPajMW9hDoGEhNyF7NUwqrpVSxuQnd
CrxSzIUYqC4WQRgw9z8966fFxioDVyxHY8qlRC2TFT45Wtn713AUQzgm/JE7jIwi6rf6F5Zr6Bhz
2uMWoeIM/j6bjOaGIEzMsYdZyaUSENfbFxHkqc9Nz6AK18PwtJ+xa1lnCPflzTcdzxHglojDu8Do
LL07a9Ish7LvQLbSHriwXJnIpkGfSUaLVDAZhEPrBiIW36mmGDgK6hsyJAECsMMeQMRYfcJhFnum
6eWS/kuC3K8rksAeKZuBpWmTM8pQhXmhN9CSOJXyGDfwdUTwWcWlHyfsnl9uz986EesYNrtACTKL
fu0fMiFtCyh2SLDkFg8xWPprfTQ3g3RrduVpT4n9A8A8vnAf8eTR8j0Z9UJ+CouXQgHe/9fLiR1c
gMZ23JuE5+9+VJTYQNOy1QWIOjX3XoJaJGZa06Pz6AE5z2GyFPv8QhWCv+831f8FOlksvpfVzbTg
jUqowTaqMrutoaEByiKqRgcgSeYVGNW6lx/8s3g1cOzOLyt18kOyf9vU43FWCIohtCOh/32ddPbm
IMRE3W0B4rgK5Ri12jj10E9g0nUX4UW7Yie4wEO99699OqF7kdhRsI4G5Da8M8Ts+ppLxwy/1Zdr
q5RuuD9U+HHsQN3I3DKPnXv8I1OGn+zf+VW5g8S0ThFS3Q7UoUucHNwsFXNJQqpwUDYzVOc6UzyT
aiLzridhNXRoQZgKxQbVvMLYDh1dHueRuCRtQmag4HXGeR1oreAvkCUyOIrqp1wjsul3rwXqY4fw
K2Ey9U24K1t8m0gY7XUT5s5iF4VPaWbCfALo6RGzniuCVLmckUEr4522lc4yNLvAxkygM/kLftcA
dKiiyT2Mk4s1Zy7mC4CS5DzVB7+8Dx1b+T07RumqlcuL5z4ICxWUtMnTA//T0YJaZphLChUg1asI
8KhxS+doHvsju9uvRg5xuy8/cWaK2Jci3+KIK0Fo+bgHSZF3PyjwzqPmtX5EogkTrW86dOrdKi+H
HDSlzG2rbFq5ZieWmpJIGeW0mlmWY03bM1qE7KSIKvdiEaeFv9tyY/0hFdgSQ9WW2cxO8j+ayFVl
lH7E3T0qSbsKao+v1yb88EuvfJFfRCOLh5MQ9ffftadhM3qLrDXvhKHxgdDEvA7AQ00TVATotUuo
0AevTT3kJINNoHK/ULEpB9GoM5eh2EVqNMquSufK9lFa0m9sqfiiFDYPYlHBSYOFSrk5+iimjZDi
EcOjWgjVpO8mt7mDIJrOzb2bETypYJesM0ZhaLNSHsXo66m8DMer5hg3IA0SXyAFboLnWEGF9dB5
dycU9ZvmyKIp3hNwrHaxmWi3uTO5GhldyQ1fNi66Fgo7oJ3fvO9e37OAd2/oax8GsvSy5iZSa/rO
g9Iu3EJW4+eahP7JkTB/6AtSjZsd1l303oq0DrImZXDfEwk4g2pE4ueRxi1isXVeAcUNVcbBszky
xvzdF9xT++534PPqLf/i0mBopTUMa4BXhn0fEdB5IZrLj0RVMg0w58uP6uzPuW1RhIMcJXrqSMBC
amkObiMy628FxDZ5ijHGMV4NE7bdbIPz8Ij2M7aQd4IQfvF2Z7/ENLLAkhiT4AIqxKVfgLNW2hjc
bf8qE1YA/pZnF9xzq/ptJY3JUOvdmoIkYib9HCwbntNoJKK4Sl4zN4oW3ccPrrd6qve7xEXvHWbj
pntbzrCG3X05WuqiD6c1sUbVdjwHR7uC1ozt58SWnBzhGpcwIg0cwwHv1uSaJQDbFnesqg+MwXmK
xjCKH0FAxktXzfy2yanbR6KW0kIqFiLsJJ4H5brsMn7l2Go1HxfcJqFi/ix7MB3Nc2HREfu83HN4
wXH1MIL8739Z/jBrYN9Vs5gb/kIAmtr1k4tHaOEbLrC7cmwZeMEJmZ5080HPaaOMKVhM3K8Z9lTo
o7XylLfA8qkwOf9k1OkqXZvatkNCJZsebrdKx89mW5fuRpB6VLaYl3uq0TMhLy1XPGfSUF5gq6qY
I1jeI4zpTr0/I2BCeg0RMqc1c6ijG4gYk+d3Q1NIbtK7uSxgRyQIFSY9JNkE+uIw0gWE5cnOYbVf
6qZev6gt47wdGQVItdQadJg3PCwn0jU3K74U/rBFGnpwQM8blpdGwDiJU4Wj8eD4gyYeIwDuqPhr
bjSE/rx0HXSaQ53G+GyIETSJ3WdC2eZuCqqt3Gp6VMPLJy8+IFqUo92rnGAy4TNFxdrLjJ1FmMza
CoQc8N2nnXPI4FnWlrePwpMEDt+mriWz/zZqwokK9SIwmXS4uQD2d+9ERqybkXa2aMSk1N7VHD2t
Yhp+DbplNUxYmKjo6mGdczwYX/RqpVPjErrdEZhrlkL5XHF6nwpXj5+Jj7zNPWX7YnAFDCErISa6
b8slA8s1wylbznV1hAOse6AFKVGNkYsjKFEaUAWMxNX4XmcqLMMh/ovuCP/HV9w9aUrUtwJVKPmY
UC87xIw+4h7HCliUISc+NIK9yp5XMmGteyMubOsZDiFvw0bAeAnmP3Wu7idGxSe0hp0x0ljW9yzM
NJx/32AUCjSYoyjnZlCK4E781G3AMUmT+D5/FpZ+AFD16w98x0S3iQQbKkfpCHuTt0wpv2dw+P0s
5UjUi7lWzsgzEJiUMODj5voexqEdcRnL8ZwOeZqlK5AOQG1aprbORmOySKls2RUwNtsnmvwXM2yP
u7SSGMzZxcHT1KwqYCuArPxR/KEAZqKqvYlNOJpVYtwnV+EKdtqLNuk10HiFfwvndD3RH+Myx7iD
2KtrnSiwe+H0l+Wi4o3lipRKwQlp2F2Onn+bUeaBr+qB1oL2hIAvO+7gZjC6ScIDhByt66/GrSHV
AYZVb6VlkpUovzE/4b8u5SS4p/INJvgA3ZQaIZd3V+h+WnRMyBQGsa3+RVPcOJAKmO05S+0GDsDF
YORY9B8alfqwd0dADbzyPXncXPeuQ81IRHdb8haQU+NeOeIgMl8cdN20lhqbaF0yZ3DrWcNryyUi
VVmPQUaK341KoUwcqYLgX7cS34UEv1S5neSm0UfkNt6jmDoOv4uuwzaGB1F/mn2A0QWzKvoCNaxU
ItMZNaO3tL8Zj70DyDnXvRUNiICOcUrEbrac2JFtfdIvR3i+cYx7qdV4iSqbZytpbnNcLAo4jaIZ
7kHVrIOWb/avzpYUW8IR5yWfFbdrE4SboHco4yntSPqGXiavA2ciHORHfMXv1q5ohKwJmhxVq5vf
h+U2alGgMf7vtHbkKlWCrlEvDlnkV+VUWvvETxH3VBDcWg9Cvo5oTFhhOed0zrep7FDgWp6MDMHb
JWhILhc5uX57erre8edLM5V474WcUtyagt7Qz0dWeRugdE/AdZvhS8xf6zwMgT+JUXSy8NMVLXkz
BGOp8hJYagz9BEN2s+W9aufYIzxXOZwUKlSCljrW/Ui7eZbpC+h8KEhKKJCTaLuistPZYUmCUqa6
i4W3+AE65GSaxNZZXpZu2ZOEOLsv6wt2JVkcONAdLJMv4YC9/W3uBTSORzeZq+u7rvUQs5eF3bvg
6nnMDoHA24iIfqEabT+KP6e5poG0Ut/5DpRszG920wLh4E+iHvUDBZWuM5BUr14p0+0bz7iwtxFn
CDbdzMRWg7W0lT1+14uqoc/DE2oPN7j6+htKR24B/+elNGt3H/QXM75uA9Jj641SwIM3u3D00/F6
xgXvkim6Ri2I6xo0FKcfVekhqR2Zxix8XcMCKrhINIOKrYZ+ECasXVzenG/naWg8/nJfhmozOPfM
fxzo4TCwi4h3mr90yPqoekkUacuNbxNyitUJp70bkVBEBP9euQZX1RaCZ6c5pz7EMTe+rxxK+AGh
v26WvM4jOupGONXqGaPQiTSE73Fo2w+uY781HMfpcQNQoWszJ401dn1keS9C9/Gc/0HoJLNchn5O
befbhj5TgyxpdvaHHA==
`protect end_protected
