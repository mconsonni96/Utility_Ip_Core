`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Wfi9WPOwvbcW2FDDEzxoBYiwDZii2t/LcF5z8CG/Ba29xxD2XXHbiZ+dh9I3wUYmAPQoQ73mQNjz
v66USymVJJiwXv1pLZCUPIkWVZWJo9Ju8y4hH3FY6j8FT9bZYmpmbu3dB9NbXvN11OVrC2gboH8N
TGHMWZkK/zmiFrrv/cssqzuuJHpz8Wk5lPVav2aNkTEWE5HArXEPH7JT2yJvqKtzIG8Wrc6wuDGu
5dX7BrTuozrK/Oc5KIKw+dZOXjNAWJptcU2nAeLKUPnj0QQYAn2rc2M4YvPHS7PtMzwBnq8+ePqk
awuFBVdTg6fu2TxwBmlMzsSrpflAKRXIJUzPqA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="er+pffphlR+arktANYhHKpFXvn+WBGLWDWEJxDD9Nms="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5472)
`protect data_block
7H/th/UQA9X70Iv//gQslCt76OD6MKPQvveGAKzGFkmvQL7559kmfPgKERhb6vH2n1/R2oTg/xFv
U4knbCCDp1NIVvUoswn0gcayM0s2Ql/+FyEUPnsQ17GUrG4oe9c105D5gVxMJTxxyFk9w63HO1/G
36BKCgJiGJgecaw1AQDOU/iORFKDPNXSVMZt30zVM9Iif3+wJ3MPEQoBqr6EqvkuZk5mQVzULM8L
uqQ519aeZaD8gqWMtDsCp4jCGpBzO4h+dfW6687ndcEV14NEZPVlmYDJ383oG+QfUvwl/mDmfKVu
+/guDqUSo1qzALryS4SW+xtNBjqj6x1QIpI7Cy+TID68iQSYx5MwMUYt9RNwoWhywt0VNKlvpwwt
HQycKagcXbH+e00wmcxSt2SWxb9eICPDfPabumxLM4RWZA48lxdBVL0izIMubIH9PUWHowNILBf9
TmiBbHcXMNwSNwsgLag2AzLWXHj3aIpTMBcdy/kjeKkc8PpFLKwt2COfQXejV/jO5M4uaDKK+f4f
YPrk7wtvI4uuBpnctgrHjysiNjRn40K/mJWGZxFSMDEYFVQPeMu3jsk/Wet3HcWmv5eQAkn4ZVQy
Nfp8i2H/aMsPtg7Gu+knr53p5BdXcpHn9gfP63IIRM+6QoRktxke363jBVvWiSQiDTi7hfryU8mI
J553I7xqay8HCe5AWnfQH/cVmhxj/UeheqcXK6rDdXacYRbMJJQOwkarmnmWNTySo7GtqFpEVIRT
AjWv+WdhvSwOl6lB+T61YYXIVNn/2e3ybZQEZqaRpkQ/cQSesvlDOBfHN7IwwsBrTv4BCn6XhUzy
8GDY9zQsgJiBsZ5564WVjTQdAxF1BhVMtjfr4kC/Lrlg1LWFN3VpR0mT27deM8sspjBOer4Q83WC
gnfn2djAJxYGUeSOfgr8Kd6i27wfRTF6cWuvjMHmU9gYBmVT3wHZBcXKtrRun/vWODSHkkNwQprO
TjTJdAVF3qYPorVfeheOmOaAEnWRjtk5Z95Jmiy1HzddF99vcRCehp4NPE7erPXscL4WGe1DTZUZ
BbVOnm3PAZfleubIUsAmDYfpukCoLS+/PvDhqlvc+qmSYO/E2CfdGT/MSvz7JRjNK34ANd9WMEdl
v1n9nER8gj2xrAAhQ4Ha3qXecU7u+k3oye07VB9UNlXTbEDMvifP6CEqcsxKD6yJSZc1WVCZVisa
/P7Bj65/28V06TkOcK+XcpBrsSMpsppecJTdvZn3mmXQWTo8DtoqKotjIA6UMPvhE5W9QG2MJZF4
WCxZSNpSWatno+m0QBY3H+6/69lEZYNupzBpuCggjCnLls5cguF+HbbcM3efc3Uif4iunw64k4ZJ
m97MiIcDVaAXrNtqXhXRRyO5Rnm/vt8EgpWWDu9/sYnVP+XrEdcXOfmmuhZyJVQC7skTzI3ok6VI
TKylF8hiQ5pFI1NtDy0Y/1Xgx1NxoVS9GvdkqS+Jnfv7gMHgygkfnl5jSjcOzi9FCb5ISZgc5F3g
OiyESCrT5a4XHYnx+XvHkndww+Lpv157/E2ubWEyPsmIKnSkUEf1yh1JCx/BKVmdMI29p9tnJyZI
hVer90ftdsGoa8ihLcJEotQJVCjQSpbB6E1kGaQXUvqM0D4osqRYkI5aiKJgfyqKvp53nsoM3x84
S/dSlWGzoPWxmRT1b51yWk9anfckccd6BBDY/1wXPeEsIqzx9ElykQIp1C9+pcQKQh74mQqXUPxq
nzWq2OhcV/Yc5z4E/l+Aa4ngtEuhdv9/Uaw0c+EPedIlysISRVqpeXQMYbNSJGVqzPGZQxiKVH8m
A9rZj6sXDYodq7euTVOzoxtKXrhlf08xXt0inH0Ql+o79halC/jHFDUpUu0iXXKS29UVOf/OSPI1
jkkdj79rtv4ReBa0Drl/LHDRm4CWC3oyk2SLQSRtY4y2OSWt2gbpN/iIrymKT14tbrSaKkuQnPtB
st3IB9qJwMif8jwZxBqseKg7petNwyrYgLYX4HgyhR79FK7JmUkxqOopqGMlxXBQgjxO2xAfpeVQ
lUk+U1nXJVdCMN5/PakP1Hni1xjQfjaT3gVXOcrA9aujPWd84yZbrpkYNzVfPfhXpaqC6I/w2jAX
gNOy8AsaSadTAPdr+QvZdVMzEivkz0vPa4KneVAGY/uR5hwC6U0Vh2FfPsk69aZxA3AaOZAWdKI9
PRpd7HmrJopamLioIM6fM22eqpoS6M7WiVpaZUfu2CwsLNXHx6r+NvsIqz2kQpuIIpGK0L6OpgAm
2GDpR85PXKudC1kUM3pjiJeq5W8R+vGeHzlL5QbFWefMc2wACWDnvlI3XjiqDXIUGkZN1vtU8EVS
bgbHqBsHO2gcC2XNrXihVOtZit+lX+d5+WaD129Z5X2TD8KAD6MXzWtonWkkIYftwzEw5vy588np
hZS9Yl7iD2MiHv4OeWUI2m4Huj+x0wXlmKwEkKrSIl0Wq8y6WweJeGb8WHlSmg5qmV99tZQ6amhL
jtW2Q2zfDe0yQbdXJ4n1/AnbFG6iCDMnRLh0m7ha1Rz/Oyg17Ky1qSbN/1aopuFzsXF/z2Syy0J0
usKQx/lks7lbLwqMxUmLHKNG4xcAvP2+jw9IhYq8rX6iZLqIw4vqmyVkPhmnE4W5aBmol0+zlUkZ
fkFRR3E7mPw3J33R6/Ju4TnKJdTsly30mrJq7X9yCVD9SR0p1lkfQ9BJNyYgeFLFMPjwVKY3ICVl
3HCmN5WGqCoKWfvoh9xFNTDRyRkK73RTvzyziCveOFBka0gs1bw1euQf5hj4LKILrkWHdRW+5YkP
AqV5rg8XfWtEEdoFd7kWYBnj+0p3FYTqinAqiHZbBr0YSRScASe+1omREbqvTackxi1vtmkWWqOy
WCp04Ev+nD2MPMAGINZpBF2gEh/SlHSmFlYYAImLG2nICOy9wVJ/G8HLTs82/RoWAornrBJ/VLHq
hi+ZoxRryF8pdgplnz7NNR6ZkdQjQhAOV/gnIU9q5i4YEiPnQ2Cg2+QLATDJutUW0bp0Y93K/a8o
5pMpBFsEa3PDDHaShgrdto3NQ9LFht9NcCUGVf+wVHo7ZnVxT0OboKbW4bkybLM/BnjksZbwNAPD
687Zr2e+7jffhjhzHfAKcjPXoXDpzs0re7YS+I8geyvfHoLIEfzENN1dIzRXEcD6gnufBeDYCeD0
DNc9HiGBA7rNzFPiuAxsLWokqIxIY2xoEUrOoYb2/467pEtM47YMPWM/PkGsGCkL/udQEM39UI2J
UrlHnrzw5EN1pVpMjgvP8s6GZvqbadkjVfIhb/UViBPFji/2egdMyoDEyFxlHEncFsNcF4Km/n7q
dl8C65M03LD3GQMdrlw8FtpZW/qKvtNH55qAEzDyIa7Q+w572HHdG6jwWLOKHhdav3wVtMsbzEG6
cWlF7VG7k/xj1/3XoZDE7NlnyW5GuoxskvLtlUB2VI7BL+Ud4edT9ZQ3X9sVz5oJueyKWwXcXABb
dFfjJMpTQwz3TpWeI3W3l5sGDua1ghq0FGKIth6PwDpFUzYq1zLsqNhEECMEq9NLF5GVb3uDHJk2
dXVmKKPsJEeInMON25HVttzSbxVO/d6mFZ1+VB/fcd7IIFHzDK+LHT7q6CcMeO0JyoSYk6Xpp2mW
h8T1HBOY6+B0GbCqZg844KkvK5afYW6uYpfXTdJji+8MZEOcy1NXCkJpwPgqO7dQeqcZfwz5DwZS
WbWKJC6buIeo1riA4QlFXkj5oM13w4VpQqmlW/Q0Vz5opfmse7TTY2nEAOrKVeK3rirIkdcVu6aq
X5UEPm90LS0Dxe3Z/yHAUstmP/GD4uvm9MWwo/KC/YeIj35dn+QwVkpFZbZ8AmpBobHpySP2Wzo9
3rva6NJUmVC8vex6Z3Y9Nhw7LxfIKSuavIt+urkOxQQ0lomws2mvIOMKIaoEltgsfVB46ro1cdnD
REBme8BviV4SFFx7QSuV3p6ypYECRZS8LVrjL4xymBmSVGt1o16A2biO8USWpHE0OJoOjjN0txb8
GdG5PsgnS4NMiab+T3y/9/2GqlZ/aDR+Ef/Ig1Dd0+yUTz0FQzVQINW/B5+kRHwPNn4XDi7GSavv
HemATKX3wSovKbkAgQfKDaM6C3O2e1C+efCcg1JOZevO+/WuPQn5dSlXizkLGqqD0a9hVOuMiwUo
IUZXWHFAEXl44E1jI9T5Xyzg/tDDOMQMgN1rYfr6Fio+WmocgOUo11/ner5JIWlNSDlDtwNRIb+Y
hKYCP+EREqogPOZPGf+0XE1GPvO99exbU4g9nczWugRZrbGh7KCNC1ZebgS2SqAraMo5lKlyjIAl
+7NBGEULssXbLubCjkLwo2/3q4lvJkYSry8EcG/LBBS7H6d0+KIpa5OJB1fit9W9R+Yrkk6WKRer
4m6uml/aTQeuwaLsz6BoS/SyskoSHc1r+K/mZl/LEm1hO17QeSwGuIAxgJQn7qX0PJPU/1RPeOZf
lIfFblruwG9RUEQgEPWo/pSJc8Yx3+QB0ElvCQGnmH4aIE/u4hI/wJHRs9siK0NKbyEYVf703rEn
xzzypGdUXo40EpkdtAIsOvs7gGRa54lm6NUqAU3uOZ0W9HieykeMJBybXRM6yyeesXJwaX4FU6ej
qWShNLAiFWqG1arrEbu758xkQT9dcRtCBdIVd78525NAW8zYXEIe+fBD1hC6ZhdZBhchEekg5o0Y
SOBfxm+lxvfgvo2P6RSbZyfRQcER0TKyyusXmgPwTsGFeX5vP6zLohvQWdqWP+TpfJ1kriIaU2GQ
nOOSHJGM1ptXGlToCtxpRzJZlLwuqXas/xMuDiosNmyrotXvIpKsYIjnSA/87DS2tomUb85Jc5ys
I+pDG+umW8njxfdj7CtHGHlHzpMlhjpxXM+hZ/v0mTUDNSRqagTAT2XMJFXshnx1X2JSOSkijceT
I1lRMVGLV51kNHuFYw+o7/Z+LjRbu6FUf11sSU+iaaz3o21RYZ3/m7Y+OnZkH3AaQkd1s5Y3jp/k
tc+TYjFNibdACBgTjwpbi66BJyqQ4RzRKAXg+m07dez/PgmbIsRrJLyfW0spUYtaVPar80+/ctG1
Grx1mga4wa2YbOX9xYzzrbhIvpoZp9MlqBaaBcelc73xhVgmf42j+kpwAWZBw+V48ie/PyJMfETp
PZnhK+EfuDRbOQULN009wuLQ2jEU6aOCiP8C8cbQgkBHbyHn3grnRw5JU3hcSroquduvVp/IbxGr
OtXqAshc1RNoi2UIQfFrvxpbADMDRoH5qLflanLD2J0xyOiqG2SJHlwPtgsNPSMkk174GX5Xdj6D
iCMr9qVB0WPU8S7DoGn/0mzSlE8cCuvNqu3RUD59uwoLUA4usbx7S27l8Cg8kseWtiYqbRLzFwlT
kssF+9fMdXXwCTU43igJ8XLPXJwScnmtRkPglibY3ZiHHYYusBSVdBxSNqaA9SSbUmS9A2RGEXvh
NtE8BxfZjaXYwcQud6eRunTDEG8htxFmHV9SmR50/UGBKGGrfqMqlydJ5NeMnIO9Orry5hgmJL1D
1KB4Wylst/Ezalg/H7T8cOyH1SYneRZ0Quf+FGB38Sp9Mk/gxFdE/ohb2xOc5rd+xOSRxTHqPkUu
Kk2lmq4+kQMHcsbsW4PkXksmWzQIgUFaBzLoGUAivGpyaHtoiQGZwzxOF8Wa20GeOus9C8zWydQM
/w0d4ja3FTh9GZO7UkhI4ErGCQ7b2y1K6aan20otKjNBBPH+bcZqB7teeBLcHeSDl2xvHHuWb1b6
eEo0Mf9ef4NPdsBIEMhUJnSoPBlTvWEUZJ1uZwYd5uPFkrMuVt04ZDPb2PtY0UCBZEpp/YSjLs6r
v43X+Mvb/NR2T1LMIn40Vo6thHXHUohG/xQO2HYVdTjHda7SOGqI8HkaKuXWvfGLNCnE5pby+2t2
HSa6gUQ8U87V4iiqdfQTXsbOArAkAvcz4hyI/1bMxPFpRvQWYUPjftmNctI07nemd6UBowB783vn
xWN/+R8gzy06ExzYzWUn4Jz+RK9L3HH4Cb//bAfgXMs7SCFY8xh+KZ4l0LNYWhTVVPNKM/sjtNWZ
Sk0ZLlzFvvbOvoNgl4AEPpB1iCLI3XafhvKhhMc20Z6Vcq3zQT98hVB1+XYeqNx9oGEw1KFAj0ce
8W1ooCWA0o3w3PXWDWnEVB9ltuezcr3CKhWtYkYoDSBRuZnU+t6iU1cHYokJCsCUYQB9fvVIImJU
Ftai61Xv0xpPZhzMXeCz3CGIWvCN6vaiAxk14pJqXcXSKED/uHqYWxM3MNKaTIKiarDDLcHRkSDb
efURDqizCKnNruco7Q56L2aTWEdgObeT+iLZJttCbKMBowGsIleNtdI/H8/LKk/WL+rp7TDxE4qa
Qn7buBR/sr1jm21/QkDzr85Pg7O14zBnIP9EmkxzhKw+1JC4Kh0jQqdnyYgDr9WG5DdXy+hgEcax
TDdFGntQT1RPXsYPh0xAhLnDwMhc4eHHqzpWBJ4sK0WaOQmspk4Q/4cQPTeR2ZokrjP2c6hdJ2Hd
SS0DVN6hKfFokLDTGsQ4D+85dzdiqNfP4Cjdea/lKXJ5m9RGVKIvc1lHgrTU1plTIi7hkcoULU+x
5Sd+XVoUox3jl1QfHV0HT+n0n9IKTeRfoJDBdUdDdBKjNF5Yo64jUfJ6SfHtTn+khztf6V9GcB2q
3VCHvS2JOPngBwJ3MLURgh6G+xeSIFQxXlRB9XvUWBooMTQXipTBCnjsHquqoH8SJqTbORDKFzW6
vca4OrYOeglz+lS8oUdWkvEHaaNqfEjuioqD+0JM6GHB00Bq+tguHJKxrvtkdhbSkaRCRLqwd0eN
zKVXRRhFEYFoK0aWBaVTV5s65pnLptMOgIsKNXtEE1IANEX+qREZW+DtFE7Ewr9yGpRK9aANzkEi
UKvs0U9BskbCuqYih1CBWHjwtHD2pgDF/BlsjpV3ZkwOk7c8Zfg22XFZpkO4rxwJe0AXzE3pdiVn
NrY6y0EEfVmlrwdfP0klAc89rbTgbxH7Ln4b3A9PYEJdD098MzAyt8L7XuL0hrq9Ueuq1YoXiZ7M
o1vAgDzCtzPgvHiuQab+xZL5piR4DuZ5sgV40NdblzCVK3e4vn7dNOmR3nAY9sH1XA83EU3qPUOo
HwmFRnym/DgWSiJabl2NEkxafEAFNvDAem9mDjh3Fryjy23uy1PrPx6FRh3WOqE04V/xxoky8pK7
RcuRUPfVVylc6+Z7qR86CWO1DP6i//aEf390xUPQ64QNp2PO3cddLZNBte78mFFhck/2vWALSRYb
`protect end_protected
