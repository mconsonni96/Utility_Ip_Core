`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ii8Qj79CzQXvE05qMjNVaIJjLwvbigLfay5X+83LE3vZio+OU4QZhag5i00vzdQbL9p0G6Clz3DX
iZSLefLLa3rvMbmpD12+c/GdXTLUs2InZ5CawkiU4fO6s0u8vG8cS10/yElSZ2cbCUVTQvCU1+hv
Lr+cTdfoR4BDC8gipjQQD8SWZFFoeLxaljKv0le5zSDbwk99Jsjuk59SBZCykyesbpGqbhuWdVU0
mDUM/isvk/cwch9aNfQBgyB2BM92INkZGqdogIakBNaII6q06OxDtiSHrjmyzG1zepUhfUgYR/qH
pyI06+YQdJ4Km1xE3awTLAY7glU8jV6h3sYqzw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="CN5Fv7r42iWO/eQmzfDXjtGg94vWIeZ0lZRbWbOUcdw="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73872)
`protect data_block
gN2BbFqkan2wXW/ZM5UEQxyP/SFEVO3hgeoc6xhZGBaR+NHn4o4nkZnw15gdK9L7ki4F273pc5Yl
B1edKy8pRL6F9tRBnkjX76xRUEX6jI4oYSywi2VqqKJD7yONGkLMzTyvi223m++ZVwD5toaI3w3j
Uj7HRkIqkbXXU24grKvKSB91fjCeKXuAX1BkZ3WVnAdv0vFnGbUkr3fTcApVnhFF/k5ruXLdlJSI
YXUvtJn2MJPWsrzE9lhRM2msVVO32Q6ClstyadOyy/LVanxCla5FjrIYquj3K3yZJrQwD9BfP0YY
RrSbZXj6c8i+JCanuLpUWb0XfasUHfRecNoi1y8w22LAUMYGzSBLAaCynEU+nrQ9UPqby/58AK8T
+F1wWeYfl0NvyqUJtyQoCxI8mYoKM35ZUZ8yTUkQ+zxRaP5Rc2ATrLOc6VJzRPVVBWo96vYyLZZR
aKSPkZdMFuAQaJ7kzfxFmW6OwmyifVz6ryPPVVcVRvPEDJLfyPJ3SNefJYuf1RwatVAETH/axZ0u
GGmFnsElYLmCu79IsJuJiPqWz/+g7wPPwtDCLgPrcNhXmWfb8dQKRZmc2e3DMT7XwY9tV5dXGb0X
yh07r8bxGvt/C8Dl27zoQzW+JkKx52sEv/2PKULCRa5FzaXUsI2xAa/60O658/xOMORWJWeMS5W7
u56mG9LNgLGxcx5NEDHOht1Lzvl7Cefmy+OXt48spOXjpbYl1lT2QAb8zKwdBpKYmn2qIX3/gZqI
VEgtNHQawjZaffLwDFoMi85a4+b95BZtKIXZn+XMNb3m1wCt4mnlHVuhXs6zBHT24qikYkc2fssg
bCauE6K0H+RhEtClSVKJwr6VgbXkR+HErW1qNJL+HJioVFcxGavElr/jVwO9KHut1dPFe5pq2dvx
XnEuQZ64DbqFqRtRCXeGtg2jN0SqOv3lCE4lqKVTNQFH6iNcm6891ZUo41PH5n0fmDWvjfzLalF3
TNKv4A5Ja9PGOtS3f45i5CQR9TnFVmHtQW1XTj3xytvBpH278mffW8H9nXp45mh6wNwsXEwDsQ9y
0KmsPQ0iWIiV33e4+85BUM56ecDsGAvzFcWRUTdy4pmYdYXBazioeon7l49u2egP5z2dYmS3AJm2
ARPDow1yGZvT1oiAdhvQV2pYifGPWjgwUDAEBT4iq8VNdhT1lsPeUd5BtGLFsr4JXRTNeIdBxFmp
sMV2WXw7RB5wFond/K5794nxVbwmJ1ZhwKR7+tnU00huBDwBzLng5VOwaVUAA7KnqzNuAxqZNugY
GXB8Cq0A3HVcSGne+xvyr1IGEW8vWyogcW+7UipsNBTvw5iRZxFzOo0oAXFziw7Og+HE7qVYicjU
xFHUMYoFi9LZSqtgWSC8r5xO8G6q8LXTgetL3w0/w9c4/kTlyWsl/Ci664aqKf4HwXjUdCs7O4Hf
TwbkfF2qpyRTLkukp+l2YgKs5S46kaAewjwcWy1z38JIK6xOMbKpp6lKmz1G+SJ2eTNzd1t5S/Xx
hfgVzfXOXYH6su75nMw28ay0XRAQHM5IlLKtbKjNRoJUoiFmmBZh45NdM8XRKt5rFrci6k/10Lvt
/h5HK9q0XDAdbj6oqW+ThS91aWsR6rg3fHncZSiZxFUyKLs99IrymMaHvpKO3KoBpcGjngEDY88s
XbJxhai+wIqRKXPAb6AYomvCFKqZR4VtVxv4Y3IzPdRjwJulNVReEJjbD4JCbMuE8XC/qZuQNdCV
E8hofWrE90DdpQHIm2tpE2zJG3k52qNRDRQiX4d1tcvL6Z75JAcaclHaeuF6I8pJmcWF5hXdgUr/
uz7+1q0diZ4AKTUZAPRj7XKxEN4bMB2VBRkiT3tw1b098Z594kcTzR4aZ42ImDkijqhLmKm/rPD7
RfEA+u7N2eEATP/OHez2E+5nGTV+KXg8a0LMvAMLsoZuOjaD/yIYABFl8zsJjMyvlw1Hco06Z8Um
wUd3d1W1GLc6GhkjAdQfCEtnRFrvK+z11DZBHCdWkXr90Qttcu43Ndpr7z42gqPfyMiUbaacp0us
MW5JMSMgObgzjAERm3lkOVz3VrKF8l2ZWCpzhySRGAv52lhJB20roXsek3K9V56l9a7928YKSxEW
5BNGn8A687/QGGlGYriQpMmN0Ru+76uixhCTn1YOLO3R45FnBfezhckT4ZB/Eoggkn0BZp5cK482
VFjVibr+G6wTDAo0ypGeQYHegJTdswMk/h+PPKb8w+iRvMCysqN5tu6f3sV1Qhh/vn6pO1bD3knI
GMxIBYZ8OHGPdErz4T3ClIv5vsMpUDotdubOCg5YX5YvZ66AxwEvbfA5VyB7VDVVPpaLq0J+fC4z
HrwQfTm7/d8exBTNW8FSY8DzTnXs+XQnjF1OJ0s+qeLDu7FNjUHE8G3xQRpL6GAgqTMvmNu2MynR
DlabMgwnXerQAjsxqAd6hlgai439lU5Uo8XDNm+4WZ4PD/ArsUQitAUmpjsveKXRyTCKFuKcxeT0
UAwj3Z9dzh9lqRIkfaahredmXOYK/k/tec9MSi8kSERRXba8E1WOIb2jDlGBJPSoOE1cOLZwq+Hs
cqFbN/p9Epbq1RsyXocd6hZy0AKpYIwRF0AhAuvbvd+rNwr6C6yV3egQbz0seIIi+mb94gZIT0Em
pHyVKzrzKmqmu4WdvVt0KT4cu2rD/7esfbw2wbIHN/vN4VcZQUOJsigA5SeIJXo/TQFF+2iCTLEW
ECs9ak89NQwmtdNYIUoFpnJg/rmUiWX2VzS8X2CDEqxpy5UNirN4OmzoRSpMtXtvbjfGfjmds6Mc
lM7xVP1c6qloZe4TT4/6UX6tKMjNV0OIOX1Rg4ssfgGhgpwcK5ygDEDnyM6oQ5+dYkwMS1S6xAjt
3Lxy8n+oPvJVIkp448ceYfX3s5Jrpcs+aERbp7owNIYmRgZ6fhQu2pb6d34sIoapI+m9c1aK7LuA
HQeBfqA88YXMwLy8g5Wgw8K02imR4nmDqFald8aNq+k/yf9BbmSji5BEyD0v8efEUEsLVPxej45r
uQFTBgsrxrVhIEvqizpYOAxbO6DE7tPXciPhVhFEVH/sjasNPRVEqMRhqLaVq1tE67vMDW3TfEd5
GfR/r0AWDcqeQvQ1RgWJFX6XnXcOXZFjQ3U9SL2VOwBunuq5Q4U1wuhcW5p8/zJhsEJboeqgGPDF
jBbqZaD+IMFdTv1cPR3VN5/KDmMm+/NKQRQBCrFh2dDNMAaAUwmpIQObhI3y7tWCipdbBCQVfUsc
9/ALMtlYYtXZg6pFgoImeO+nRwxKHqIJ5UTQN8b5tv1mFplZWct8xFYrgpAMbvFSxaXo3Z3MDNGt
pUXvZnZKGwWVXV1bLK1Y3NgSccrtCdUCYCQoagw4obcwkv6ADL0LST/dA1H1TPB/TAceNlJsUs5f
ROA2qQBQg6mwVE8BBTlsLqk+RgMFvKCs84+Qsi6gcE4q/+GWp1opxhzuLLbUxEP9Raiazj4OIzRW
yoCMrXqV2SHel12J6R1HVRTaejyz/z79z5nb9WPXy5BtYhDFtI9TLcU/IfcfZa9Zch1U6wJOxiDB
6ZmhW9QqRfGLsG/JRaYKbCeuTt1K0fZ11gLxCHYydoTKWB5v8I2d2IXiK9PKme5Jnp64GAJEvIDv
msxJjhPR3FJX7g3MW+c96PvbSb6iAd/low+/ZPoFdUhlk2DsKOMm51Qc0++jn1pSlAx33CHYBYjf
bgTVs1+tcxjY79H6sqW5vlZphDA2dnChPOzF5xZpJYAB6b6Ofd3S7AOfQxSXv6yrIb8kifDI2KJY
xPI4jz7w1ebd+necNSIEdM1lGRLc189QxkN87oXGGVicTMGtghpATj8g0DG4yA7vtkA9wXf1ZYK0
UsY1SjU5ubzdt8Yebve2Z8Cl1dfugfIu34gbRF+Cd6th2Pilgrtnigx6doPjJsRtawy4UEJP0xHT
jiJbeDCeOUf4OPdFd6rRMHv1MiXplOxMu6U0laC8hrq718rP4o+h5wMV7ln10lRFC7W+1srE7qbJ
cnduvkhA4TiISn0IiBgAxvkVpNlHFNedirO35GPPNRad1RmOeXoa/gjlE0KmjnqZepwxcWruNyg/
Reeqo0ofL9cTcR7+OGxExQKgFgw9wfClXv9JsIi7XzLQn/BQILHgJIWkVRDEGudT7jNzk4guHlO3
jJEpa5N3d5qGZFei+JF3oBbrv2bE3aeU4qm6/GUPQhMRwjMqd93bXivn27WvUvc5IceJrGMUsjSB
yGtvMlwDLzip7E7kyznQYzTyxigkA8UrXrqc3c/mnWU4Lj5/hXHXGHfwBZA58I0Zo86L5UsIn0BO
bf5VHu2YWNQ8N9e5h96wZGtsOlVwKjd5h3v4q+vk3rNO+SmwZdtbGKljcnroPkCp1c+IbGYXRoiz
LzJPKEGlb4GKrNGHPGb9VDJl5h6z4784JL727ErcQTk+n5g8OBYhOxRz6LfDcJZFVsXlwg+lsc8y
XTdc/EXBSfMou2q+vFKfLL/YRg82tLC3JCj/zDj7nKU/LT7U5Dk/cnA8YbUoL99Bz3J1JPlFeotQ
9claK5+VDFKkvKiHSZB/paT3GtijryGyD+21HmP+U2xAdv5IhqEcL1jaQpo3cmJcoa/2HdO3gNGo
wBEymi0s6xR3nw+1EDLz/ZGGjfMQeV+P6y+EojMQKMcfjJdECgPhNhsFC7Vf+6qoByEXz7JoHpBe
sot8bZz9PzcvMMv4TOBCyRWtihZyIRRVFI4M2H+iKaA9Lbc5Hb7XMUveZkpwp5oVG0bI5mCmD6XW
GyJzjJegR+nsl5ybXBd8pWaWA5e4O3O87reK5uj/ibrhE7LJX1PT3NsadvOHXK23o3q5bevt/pE2
tLV0jPdMwu0oXhr0dpcBtuIDIeAQhmik7qJiS6C5qHYr/LvNFwRNDaaGmy1PBMWjNmuJxkXN38lh
3wXY4i95TH2aWk7Mv1qFtlDuk/3QiKy2aAKPQ9O2JxK5Yqb5Vkq89YObEgBHSmQAuedVgqWrjJhO
qebk+gDQk4Y0ROnhf9gFoK51J+7mH8uC6SEzy9Qh0Sn7B8KqTrOEzhT1drlifjS2JjzequolITDl
vAcSHUyRF3KlB3SmmvyNveGzmXOc0wGsKo/zS6eQBdlU5iPHHhBGehu6kp4thUKFCadf67OvCOyT
crd8cbfFGl70un0jGxrOS18ypr/RH23olXdqwBZ5GRSTc+WwnLicr+XnAUJvz4LrjPUKNxrTZ2ln
LitGQnfzCv6ESqSItJ5FY11iHr1h2/kcjE3uRRQ9LnxSfJmflyIcB4kp1Tw6U1hFBgxpRiyt8rOa
IuA+W9Qms/i0GaVBZjN6NGsuDPR7lmKr+eSHYmiyd0IYDWp2JEzPThf4Maq0rDdo/1v98JudvTLt
HAnmqiBmqk8dxnYypHj0gxCD8/m4sZl0xNo7Sb8kror+LURBgKq/Fsko/3CuJjCFsnMPy37vRnUG
cRrYhYmB4iDu5y7YYq8cR/iOk76HGrbJSC0MVdG1qHpFBGGIbn3n15ZP+D0gj7Vcc1BkgGQ8/ldn
UARxBYdeX1sL+eQS+axbkByWSS88l8KNixudLfZc/2KeM6OPDV/YqawXaSiPOC/UkhjntSjgPY/I
KaYtY9tV+fwLHMDbpME7UE4vipxZHNNAvxpvj/ViQIQIPhPGfiIQhLQigt7rLU7JWCvr+CjRtj3u
iPnll0RurkvLawlqrio1qFEBXM8++j4VPdhb7rU3YhBiDfrDQq2jKTBF7dZPfJZO4mi23Db1u1xa
0W5WM3Ejp60Yy+mRLJy1hhuAsvKdRD5gh5R/1EPojGs1cJhKBERunUSq/9K3wKRfvG0hG5d0hS7W
NgFGBSzBjhz8KvWTOsbg6rHaI2waN+8wVqdnHO7j143yV126VRxIkdNalEqOKx6dJAw7Z62nwiy5
S/lX3AaNeNmfaLPM993+fkfYjez+TuaZn6dfxxcTN9DgjhX/vfADvfnm8a8nBqqMo0DgwhUrZEsn
bsBS1aZoyWUhumXQjP0bYeqvuuKPUiUO6K+/w01zcgT+D/rmT69U9Tb/7Ezgrztm27Lv62gdZpqQ
tQSAuHm1+7MhoNzt/LD6X1nXNKjQUWO5wDDiXLIITlJDyBtsO9GtHJAtWCwzcf/alnKv+u7ZRTYH
jhWX+pZRQBWzNH+L1R28MKVZiBPYYi/fwrAvCxneWxPS4J9yPdnVNQWTM4Ce8Qr8bHL+MjC5boYa
9wQ3Hm5X9qe3B2oApwhqVS9kG8XxLLivMQuw37ojqUfCwl5npD5TZOrvsPjmOIEcRtBlWIf6VdIk
R/ZVaUJNyh/srrlTD/t4MnPGPwxrBZFb73YM7rJ9Hx67j0UFuyPxO2mJ17xUptmwyNxb56yXHCuZ
RwPVsovbR9Bh+CicsWfs/IMcWWwzBRpfyCuOmx+D2p7DHHzGIjVnAHIXdQZpJSKLUDXeVB7stZW0
gy4nLHDN3XeoylhKLyndTZ6oFnvqG2YSQ+Jv28NybGFic6JELrXJHFkN8IW6MRcfZ3v80UgwJyI/
rFtx47NA6Ey2LDt0SPqXtd3Nx+Hdf1fYHfxTZ0sEL6vnWZPW7Ode02LU254YcDvGT5J5QweLk0yA
fZjhfQrqVBkZquMzXMzn9Fq97rj43jv7mft0RXjJFcuyccbDNTpkk9th0w+OJl0Dm5iiJ7Uqc8/w
J9CRxkEEDL1i52FFBpm4NQtt5Cpijn/+eOENxUpCkwYXI3TUEardmi7GSCFyjI3N5YQ7x0+at6gY
i4TiFBcvD3DstCU1xUIJQayum1OZ7ug6SRCujQsze1sA0wbYVWahCBX5ZDcx/jST4wlGlZJDqegz
ao3m1HjO1+Lw48Oq/Z9Pok1izy06zmig3eOjqUnDwBL4M0P8K6gdh9LSwRf3Mldon5xmi3jgAjVc
3KEW8UDRE/2rqG+qP2OOeko+pSSg1sAxvIQQkstMDG9wEbq1hnsNiN8k9MIoq2QNkUUelBdM9pO5
ltdR1fg2G9z5AXo1lkgW4sux07viE+cuz+oIMiQgerNogTIiQbGOlnoNBF+mOM3pG4mRR84XegLt
K3muT+/I8xZD7qCxlFy9d4qPvZDLDj1ql1KK5yQEnna5yeIfo52PA9oKfIsC9is45pP0p3cFtBYY
x7CgL6huuXQxw5PxVtyHKixw1PWJSvsja3D3pU7PvwgKGKK0dAJQuMtcJ7DI+R3rtBm74eQkeV12
mcmuxWTf5yV9PI/94hKY9uWSV/1rAmrD8zlikG5sP892BZKbzl3+NsGj3QF54NSJao/4T5hRGbFj
v2GsEO7TUo90VX13ElncE4xvgxPvfNpc77JW7e5A6RTqWG8OA9pwnvZkbotRkTnyMbPMGH0ABy4d
2mUdAWYf3AfvseqRGz8A08/FSuNUctktCoStZJy+DXDCa68chGjvUagfhYET89pUxMnXNwO9uQNv
APxYds93NuCHUo/Uf81qYO+nWbRdfW+rLuDxVsAybHUFqYbg/p2sSO0c84UnligLRMHE0rdPKcyc
tc0jIEuTR+f/2JW9SusRBxWtNYCxNGyH2qQCq9lyP3Tsp94RW+neOKrBXZYbWbkfkg/WgDGQIG7j
hsonVglRUIybFL/Bi2qDy8HcrQ5pmwBsfk53gUFp1ewTka2HrD7OVjlZ/4xjxEOXbjz283SinjCV
FR/WCyaCMu2UWvuZ6aQzpkqtfjkrGyG0tkndKlYdFUxmMLAoDS/2Zpahw3zuDUFO18W/99urOxcC
OH0CbtfRjUui6caOFIDG06Taw+WavJLaJGXLI+pxWo7fFktR3fkRuIIpHmyYAKc5KGyYFgTAwJOv
asqs+KcNeNvIwsJw/A53V7hnGPAoUFdxLkiuLSaR4MDzjDAjD//pv/MDPH5uNAMOigIw8SF5TBb5
8xeMgs+AfeIkMpatlQ1pMKok8DSkDGb/gROK/w9ldJX1gHvwFBwnX/SXS0JP1/KwlBWg0Z56q96d
+i2vtJdjZLNc1w7c71IguNVOd2+tyvT9UjZRC9wb895H+z2tCD4/ziZwIC0W2pI6qMAZBclLfLSD
F+KruttMhn8J8WE5EbhkHWhcA5wfASDvBNw4aB2ugPW/m0Rx4QAai7rkt4WEaFvp+0Whmvg16Fkx
lZSpHhi3HUbssuAhwIV/5ra37Ts0K2B/+FJCzLKw2vX9eGsbiYquYr4KHI8hMbSmv570Zq43HwIy
o9B5tl7R+LGrb1JPfIVFocp4OxcEa/JXa2dQs0V/D2HxhcVaHWa0FRVuihxo5GIXZsLFJlE/gozg
Z2tlh5WpnFl9/goUow+vdLVnKdv6qathGSMSCBCFf1Sgpd1O1oAJ4Ezs8w8kSK2OXJwA7K8zNvuo
NrhCldHeHqzKGL2RbF6PVEjbMPM3DP79bLyqzNWcNpCC6OQ0QDbnar1xwxFjolKtd/nvqd7ljLF3
+c/3HJ+0M1KIylXxtYAhXkbSpqVzj/1OPb01NPcthtxAAxk3otiNEn3wd4o273+H13ELM3WzD2kJ
2SS8FIkCJZ31JsHoPw6c7wu9CE3osgS1g7a++uZAvKyIRB0i9idzdCYsiopPH0DmZbBchR8+kiQ3
le1YXq2wAOohK4lWsLpHNfaVYv/QEdSbUQN2AFA+kl4axFc9RUkwwIKVJ0eGykAOEH1hcmssIXRm
s5hQE993PSQlfJBQUkjPlFbmhtZq7G6AxAkGBVEhzFmtoGDt/hFwyiNEn+R51ce2dhU45zukTTgK
s/kUStJ2mNMi7OkjyVuj29pmmS1KoWOLJCzlWT0n+ZS8mQRyLry5caPgmaOpvoUiqpZtTgtXLcBL
6LkJwn3Y+80S4A/6kLeqXcyKNRRJI91Kub/nM+RA4t+IwwIJGQVPU1JRdyomWqby5l13RLMQd5SI
alzk0TF/Qkg0YrAQZZGOvuW6tklVotYmQ7FkGc8H4AMbesEnDVqm8NqVPnwsrRaBWbGq+66RGMFm
IX7hXmNgHWwRHL/xD253IYZJF+q9hCEMHyjELUTWDT52gBvfkjTrbATpKGcyzyzhSRQQUxeaLwVC
jv4rHNEK5g4YGyDQy12dDRc5t/osVddLkNHqnBWi4jX13KrmDgF/IVQF+olSVXCxO06FoEjpOSKn
ZO9N/HWMPqTFnkbsu1m9iYFl8pDAPubXsM13buR+9X+CWEg6N9V3ITBvJtSrtaVjjx9m9juWLifI
5HXmcNxpVYuyXwby5hNn+Us2iJLK03ccn396V/P8YCHy0JPV2/u4W8Yaf/DQrLfbqbxxSloyFabc
etK+7RaywZEJAbCH5doEFFPGEj1HW5Nrf35mVuq5gSsW2JS68Ga+fxGSVvsUgdrniLbBOA0lhvxU
g9kzRwQhYGJQRz/weVynPTSVgLQ11yGfznn6jCwLPMSaf/cAnQy1eJelLH+30IdUtxYE/zhOEovO
pfLWCdAcHgfROyHpKxdjdrvWEtEMwG8BS9CAmuGw+mGpuGI6zZAa6ZhPAttAyzR/QNqtBMUG5lSo
Em1NvVNSfMpgE+dQqtMZk3+8sX+qC1hA40P7HZlcuiOUZaCcnptJNM9OjpM95KtdjVGXPZy4FhSb
Y3eN6dQVef68WlTVOntR+xxlLYXVjgLr9qfNLlAh2ywUTExI9ehaOlhiAZM0N6mZNV7t0Cw0NNmh
tadTeM2Ppi2riPi7dH1p4o8ng4pt7K3tIQLiABWyKPCS3KzDpSbsE0iWhiEPKbvFS6Ct71j2tz+Q
BJlZp2lYEv76eqNg7Klnurkqopzp/Cs96JRujB/9RIiAF7DhtU4q85tbZO7pElKxgXpxwqKjB5iC
mLgQQKfQsHq8wMSrwP6yrPuUkLKb96UIvgNiATA75u2wYPQ4mSvo2CgigLsLGpEUUIc1tFr7Ukk8
tuwg4Lg6g3+gt30DPaKmrEwEHPm+rLVc1+UjHjQMY1FJh3zcYCGYh1qlP8aVgn9JiglIKsM7cVpt
/i0U5efI8RVZLuR3rOGx/bKL5INp1ZJvRojv2dAV+JB49S2kJmb+GNAA327CjS1De7zJUKNj8M4e
IQgYeZUKzOOTMTAKDh9uOSxW+DScDQSFELU2hwGBV+8jbFLYbddbsDQc/8aLFVaZaTEhZck46s7e
EfyFJEBTETQ113R6u4McQS5h1jpLK3DE+GQU9donGthwqIjE4CK+oVe5cQjxy9p7+uPpMx/u7q2K
oXmuYT6JVDWJtKjmm26NSsYbVdmy3KkqgvPPK5n/cAg3QqyTJ2mTFyLcmJFltNDIe+nGuffOlxqE
BShy9MY4mkdoDWGIaYw0oswFl7N6VLIQMMeOUwcHmbsnDFMyspCavU/vTma82pe+aXr2y+878jT/
Q2GSgI4+yEu6cZrWSNuAIGEHp2T+yL+DPCgkWkHoKvGa7MYhWhSqB5IqabuQPK1PUcQ3CTeT5KqE
sS1XksostTiQ8AXj6ln1wv7yxqRBnvt8qUt+LmWSRvTqBLXveDBlR+q+yd7TbQJ9aON/2OD9o3Eh
FHRSjQyySdJB04uwK6K8XSDIMP/heCxxPHwi4+Hc8Iqo7u4Tc+Z47cepWgxF2IUBpgnIsx+EZXy+
AZEMfdeS2JXcJIOELkTz1gxEnlAKdd3Had/oaMCG1eYTy0rMGcXM33+523fZm52K/9X8Z4XcVq17
fhAIOIDaeXcONBypMGhhJdpr/LjzxPQrGyKUgm3IM3yshmrm9WTx9hPMG0x+3ZRnJheY6sDGSCkG
0OHdtnLmO9ok9VYykMK5IXsyF9LaSpruQ2zWHWWgDrY+qaGJPiXCnU/ez6sv7q6WYMpikreQNNYX
BAlAO6O7c6BWsvdgWqQpqqSUgJT597jymqQuNcTzfR5ZqgaV88Hy3vCPv0AcVdl/2nq48Iiczn2E
TAuG0oZTO8XTCC/opEZA0Rk43VBt2eoPJCPcSSM8lYK0R47uC3X0k3dcN1KdKjop7N9jcgcS/sFr
jREkX717ZA+eb0Osi9DN7u2jE6uvKjuLQiPfh5zIoGbeZcVsulNNZCSy4sbViNABYXmI5yeVkzam
9ZSmky2/crKb6ud9xCvloaRkkzDnUfPFtnmBUkQhVX3F85u2qfhq8li4EBhPUk6ciBwoiZK6ICV+
lLmWdOJUxnJMH5nnv+bfJk7hH9F9roKeU4X+B8KRVQ0lQQlVtYV0jkVQXrNgVGfRhQg26MLac8Sn
4DlNs2gEmDyxePlBoBNOJ0TamPn1XLfJg32DaNuS9VMwyyCtJ7RwuNXTie/XS4EHo3iYDgDbFB4y
Xet0A9A9xGjqJDHvSib1zPlJB4rDa5+ET0xRsvsEAP0i7Jt/MB8E/m9ie6F9Q5iNqg5LFSJdF7Va
PXEjMQi0tOKSAJr/X7DdyyYTREkOLFM7Ri2KpgdzEMyLrKd6t9J0KFWbvEynD5RtoA+ag8oFbDw7
sedxo4uJGdVO7pEZ/+1JQrL/OHsdvlZNIXv8gla7o9n5oD4BLb02hftNGDDgXMqepvPPgYzKM6yu
ZMLFJGJTd/n/zVvm3niV9u91ory8KWf4cdZFpPtncV2otl5GwfpT6zBUBW9WxnEDkCO1nhgPrys/
vW7UEF43b09ilPv5K3LCxWGbs1r01jFTXnKmkkQ6faw09flpztaCV6NLMUcxGyy85ELP+02fQtgi
RubY1cuqpAUTIxN0DMY+wUzqceIrvXnMryGX/hxbFs4LSUK20q72tOd7XB2Dr0BOY6DO0TigwKWI
zz8E1ai/696xKooKh2PxRT8FBo3eqfK2aYgpwYmqhQUzGBxCSIFbp/CvYrB+SqXNiCrmNLQaLNFo
EirT0zGQ1rwljGs0VPP4zEHuz38twlFjcT7Urru3r1FanaLYWonMAMH9/PkCF3XFxtdeStpNwSr1
LoN1BvDU55WnalvflBC7Zzjsayg5OHjNum54DQ0GczFw+oF1zqwbDwCHDjNvwyGfqSGsnVvfVeLV
1lMM0dVb4ft2UnaJXYf9Lqnum39En7szb8kVxzzrGKYtQY99k/cN8N3tgBQYDUJRAbHUwYHPwnZm
P6jdLW6IjFNKiz90Kv9ayfMQWzh7sRKpW5S5VYHuXyQgO4F69xHooEtCih9BNyi4ytJfdva3uMch
dpup7I36tAgNKUUBMvjXwrmw3AnPkXiars+ydOKJizcUKnvAYlfU2g75BQfJkMabbDow1x9WWhLh
bWPSelIiLPSCCgx7AW7Gn27c0JnTOQXXXFbF+1+GIFcUoNqEKEfkUmS//E8iDt5+/NiL/nqpPUGk
mx0rsOBvSmxGvHZpFh26suCaaBTi/ygCPtb5GWg5hr1G81iwAm3zlJRkfsJp+mZ2FRrUzlRRb4xU
jkugawgXTwURItckz/eT0oSoKpFp+XIECt0r6sNbVDxFBwbGaiszA6atlOVhlzmpbUkfxQk9+/FN
sEhObLHAy78ZXLCbDism8P0QX+xe0yuA2x6Bm9MA0N0i47ijLVk2BCR8UgI0t61efAHWRs3ZLvBM
fbbL96cgVOIh+U9BfYl5A1yFqZJUl3hhReJ8pVurRFXD+DzotrHvuTdV1SiASky/9uKu3OfLAMzb
4tWLQ5vAQF9JfZUEpLXPkO4mQwLYu3pA7JHwImhtPXkAfvZRHMLVQRVciueGwnk5F7PuQ3uV3axV
vwfbtcl80j1UD8QWLJZ67d6Go5abOPy1/PeaIuYWtYZKjNnKj7fSKm7+9TsxIWnyOrZTa4uk06ak
lOOLUhf1O+7XkIk8S+s4ipgUX+bSdfMubbEelSuyxQq2wEN//9FrlgAvBnS/GnFUCvSJMN+6bfQs
TmnZqgcEdN3nAiROE7VPp/F9pHQF85SHe5fNTrtpII5hffev02huNx4oFoZNM35gQ3m3LpYK0YIB
HT11BHVDjApPYNIIRSQinL6Pgv69Hy5H6o9Fm2zoZIwuLprhw39f69nGE5LLAYtLPbTXuYnbsl3s
xLLNBFy+Tc9jJdN9qvyInqlDgLJjKhOv9S1rZxJbbvylCU6PttjYBMd++CcGzM9Zt/QZq3HTQRA/
4isbcdXYw3S/3K8aLFVWZYjY3XnuFzhNHuHOFFryHCdZ7DLIQMulsPbPjScYRGLGTKaF018pRqON
ggebFz3uGPP+XFpqS++kwalLk1hCmZDNT+WPOOXFaW+MUDTBU/fTgyotKr+JESaw13SX8t9p9puu
rBVQgx5lFiNx8bxK0Qj/eaB3pX9LqLX3lzPTGu1tpg1YTlEeL8SmrPXng23Pj9YfdMadKeTt/cRB
As2My2Aa/sCtA6Qf9P/rZoRFRc2Mh4zN3t9uFczl/y3BIasXBVNS4UfxmRjRS3eKcc8mq/w1DSVt
Vgdxl3TiigK0rPO/eppR1q9qAB3zQVDhTHpnVE5hL0bHfIvZx4jGH15J+LOQXETDR/8EpgfE12Th
Jsi0vdBgz2/at3FbRIv5z4E4GXpBq9M3w/PDkBVetZ+pvlxCE3tYzxIj2DbkzJ3GjiEWh3EBbFyK
cihrq+hYZo0vBWWfFeilsZaOCTk3hzxb4dSprRQN2ZzlRfENyhTamPDaIapEPRg9J/wACcXYoXwD
TlcbHtKrkG8f795ehw7S+yfE4fjE6ZZfBRIsBUc6MfZFjqh97AYPK+Euj1ToqbVzLbyEi/CkUeGD
4Q12s7NfURKI+s7qIhXrZNCzTcZ/6T/7dZqYouYihjOzQ5hnmbjRZo0LsabwL+DyveIdgTQ2KvEi
PJ61e5s9Ad0Z1xE+pbl59qbL4+qX0Lubs22UNDA695W8WmLZ3OQqE9FX/zoGT3sazHCfEaimWiqJ
5DXZ1XkRN9c7yAwSR6szicwRxkbUPDZv6s9SN6atTvK0XI1Y08iC2Q38C6rC32qnzlxQFannFInO
dRuUR67tl49ioovla7D3ESORHHhu6HJIvTbEYu0071iRuVfcytEe6HaqQVf5kFfxWUj2OvXDbPuE
XxK2fX2cM9DuOH/ksZLDcXvHvLerAd3f6azMPDdRAPB9QlhlJbryH5Hnyqsol/dIXg5TplRppVmT
jCpiZl2eRpwF7tSLtSb+bCV7RZdzOgfafxa96FY5pRwlwaoKb8eiPq2DzmygoWsJDDhzoKLQwK/l
5moIv+I9RkoRT2k+xGg/pH58vHIDg8FvOxHC+pV5uhsphQhQmozjpFl86jrL0qTAYSRqVjKB7ohi
IEpGZ/ETxOdF9bKTmxrPY2zf5tEroNiYQfGGNhRMKE+1NsCKFbBrJ5mLiFHqf1sD5Db7GLoMpdHg
rRgaH3E+FVAzzx6IOMgLdRXPA7XPXIWB6MoYfRq2i6wCPCmmwoATQwGgBWKvPqjJkL5Td8P5sPt7
5qkd4b389/s8SlLYNjkenlkx5tv59ifx8Q1aY33e+XzMRG6cSTDgQyQE6yTdlwPgC1F2+ietZkF0
mCPMqleUIDH4zY5W3NYko5K3hGTbGkIRLFnIlhtt0zJG1d3ZbnTGRk9UBhN9OnaSImRuMOHD6a4n
Cdaufw+Ui+Dj8pZBHAiW5U/9eAQL1pPm4EzcUZspAl8FwdigeyqnH6k51aUEmP+PHcNufWvkiiZA
+xGj+6w7N0wI8LXAJjD5F2psE3VKSbInZhjpWos7fHZ/KP8s72YWo9R03P9lM9/ivecl+fpI7ijs
+Yoicf//TX5CZOMPO2Dpr+3t1bHPkROU0y8lGcKe/fE8ugWwgm5rQQY9R3iEUle1uigWD4fgeE/q
dLU94Ug5DrL6K279Wejq3LQv1gx5B3Cp+fjK33eOjuGi7chHjvsPwMnBSznbbfDxD8IfQ9qd+tZT
G+WXI52dfHtAJN8PCwt2UKqXkfe+Hwd71+y+idcwJaA92PWjJ/salx1s4Rt5/lKWLKS0iFxAtJey
SDzYIuNth2THjby7rIafvb5RefnJ9IcDdPV1iDexI6IOkx4mPe2Zeli7gul8gHij9rIBIYiAVHcy
apllusQCB2udX7cTOTNyDjbMJSZF3cBSt6o9ZtG8bLBAh+2VZ5LUkpSpIFEHAJoWOmms05MJvZKQ
mAP85GSJp6dQn2km2vqa7gt1Ekg50QH3AMjbgFs4tD21EbHl9SyyJXEff8l5uYkddevxoM4nL7kr
KPMGTw88D67AfSK/Xz2g6r55llTS8xCZ2NHFLI3RfV4rJxjeznrgglC/OeGWuSD8AY4CH4bmHR/+
bVzdXKJuG51dQkHxHQgZcRuS7dVdHq0JcRVrU6NnydYCMOdIgoTINkb1EuzWWt6laIs40syfzn8A
l2O9i9OsDaXOL9iURFOs7UANweOc/0JMK57S3UpI31gSHWNW5oOSEn1MRA2l8b9Y7mEkcGBo9ddh
XXFIuFmCPy2jWuEoASSm0dVowx+DFkzWIpiAsIPwoLzC8zC//dSTtBoT/bviOzSI9tLj1YIiAWO9
ikezpe+ySqYwOf2Mxmc6R3rSicBylycUPLGfjWNAuKiwG3Yqn13xF/MdY0OEe/0/ucOW3Ek5GLWa
mCOMtnRiYqmhDSeuvcGtqW3egEW5MM/zDRZQWs+bC8E6lpj16+adtVzCstnlvwUpOMi3QOUIN0gf
liYgMHxWHuQSt9bsdSRQ7NPezMdVhd+29pHguzdGVv5rvf86/dEOu/UN+7Hvv+4uZJm2jpYNMaEN
rPuPd0mCwuV6YdERb432mq/zU+as6S8y+b2Pwk2I/iEiMU3eaIzTKYrMahXf0G1GTQRt8sofZIoj
HtDCrltfyYFu1u/HDfOWlZ0Dirlffvj2VMP92+Y8ROTzbGyCemULBi/77wJk42sTH0bu2wLY4py6
bitEPFqO6KlD1oYeQjTXNwbnrTa0OJwf9HT79szRp0fWM6d4vi4u36F5TYCCtxhvKvSvAOUv+61n
d/HOvTiDwaWZRooI0EjDkjx4oLK0IRby2MutCe/li8Yr2LX9Xdv29ZQJ65CQGjgQmDZV7JKq+y5L
qjrn24pfADzHgIWFxOPJ5aPO5kPNN+pfahz6YzYN0PMESft4HMfSHp7Q5MeppPI/D7dJGYoAjjCo
4HlT5SuuH1puDK4gGly/lzU6KeHwDvSr2OYKF9rM106Rv2WGvzSnaIoGzjZUNfuZDVZMi/lr2dEA
oy2/I6F703u/ZL1JbJaybkKowj5mm0UDxNiisXsrWuWP3OuiULy4/qg90m6LodOi41waB2ZqXsgk
dJ4/3kO4ihW0dRhjVbmnMDj2vqxGA6XielrPaI7I24qNN23iP45CipbzgNfl/NcMk9OOR4xix6gt
ky68YeW8JFtb1gSLMAz3tcV3ePyRYjDLyFylpLEOsPd4zwYTPN73ALdUMyQU69KKJszHiuoVFDEr
vQ7hWt4P5jP4Pca9jYdFS65tB8CWi1C5UQaTjAR3AzKZZlnWEeZCseEIGDeaPb6ixnlmePGJBKjn
G7Z5lu/K4EV8LkFj3fXMJADbS+rfffc3boMx1er5Mfd/QAp6Rg+Hm+IDFnC1r1MlZi5VcC8Zh3U1
4zfDFPOnthFawDKPmjCFae7BZhWNHi3UcT0BMsGZY5kX/Vc1+VmCdLqcLdmddzupeyi+TNfH2T/+
BvVW7wo81f981mhl91caovGONOWX/O1kFh1sbTEkt+0iGx+5FgLlgUk3V/vv89NXLMtziHuj8okj
hbCRXyTW0GU9ORsmJhLgc1IASqgJgjulIYUpVBRhR5N3+qQIh9nzD3QUvGamzsYPPSj79BE2tu0c
XIJyWKBDK4R9amRBY+sjjR/vTjmTAofOUoUdcWs2NDrOXOZxt94OM7BkVKX9fHzy7VyBG8CSVNrT
keeFeTdHPDC07ySWfi03SMbJrdFAiP8+f41BALUv5BNyTAbCVkoK70G/CVtPTlXCqwfdDsABG9Mr
iPAOWE1mCooqzCJVNIa9ExJX/xDaE000UdeMTTRxqN1nIWAUv1YjUkmZqGOh+4IY7Np0yU2LQyoW
wTY5Alf7+jV27JjAGqY1egKsVfVtFaGEiaPr31z9rXBii7uqP1qSbxkYjZGt8AOwSjjx6xAFPNZZ
udUuP0c6ve9Sofy6kVTjuiHi37smn1qk7yfPR4S0Ex4VjuhhufI0sw3pD4hhSdJRw5v5JosvphkX
Wl/g+7Dj4lMMtgcDnF8jaVbuRIYhmUSim85WqRnmA7dTWyEr3ozj9mQFgsfZaVh01zlMkvGs6kPZ
uvl729CZxl1TzQVLuNl8TGJ3e5kUSOBVeJRRx8fTuCcH0DgXAt+bfBVkJJ2176tW4z8Mbtm0NBqh
3dope2Eb1cpeboaAw9baxwH6WReHr+Yxg+wSBV4XxjV1LVGwpLGgHuzyvIH8t88VHZxPzw+u2PqT
8h6Bg7oJ1QwUsVDl6lPXzRa0pkRnO0IkV8HNpi6hXpZJns8g41uOReO/wEbvakf0VFnymMEGRKCE
QG+sJUoCmhtrbURe6K2Ksoe3CyXJ0SCF2fcwNi0Mhh4BMWI0wZGQ7Hxq9oyBbQ3PZTsDXK9QMQLc
ZJnMqKao/1FTuB19LizxO6VCSMM+v5zQUDHV7+/tBtELnPS6UdhEZI7Fh8Zq2NH40tmjfbSo2eRd
rZMblF2dmI1qHiTRyrsaCIVdIsyzvNi9uneo84iUPJe9nz4gvpBEe3KASbvfx0Hq7zsJZ9vdDN3A
B25rP4fC/FGDN0VMtkV4PkMWyPhWxZmAEzJVER4v6jQdICwQbaKzfKCMIbbte3CSGTINdUXkU1KF
ZUP/gGj4IMBdsvX0EhNPngB7291TOQQGSfcjdv8ao5LKTtRfRA0Kx/dL7wpTVU0ub8NflGDiHUcJ
T1CE+qP6ODvHoaHQkaQSI1WPK0EOH6b5Bce3FdKs05Wk/+0Kh7FV0UmAgImgFFwuyB9YZYoT17Y0
y0nms9fh612qlQgR96aL8mkXwEaQqRwl5iAXBjXrXiDxVU9wePhGqLw8cLp8lzMTUkTFQtsk281U
b+Luuwq1gtvBRR3bAKrXixoaHPiLFwNJCQOg3DUSgfxPtlPx5OpNxSsZX5fvg45pXDzjIjiMlEff
PknsWP1ZPEEcLmd3ZQQrb8mziWgx6HvgcCf+EmMgbXP1rvKIvEXy3Agwx6jiAIYe0Zyi23NA997+
iPNEbBLGLp9alMxWBUPCxULBW40UsOzOFgSldx37yansBUfe2KKrRVdocqO0Ed3wAzooXiq7fwhI
M+4rfXsquTDM7vK0FPFE4ikCE/sRWBwPLH8UrkdjmrwBVP/w+ZRoep8274p4ILyj4C/hK5GQxVJo
5P9p9OOAmjLJoEF3RuW4wOFosYD1XgxdQ22VW00hIdVkEBZ0gNdgyTR48i8wYm2eOYILz7HFmDvw
3uMQdZE7zxkR+Q53Uwtkavi95PXTS9MCguJDhZQzxLFTtJn2qjScClIm0wA15wGZFwsY/HT1dbyS
zZdHXu1Xk9psEIvJlt0WYOvsfoF2Lgknsb+tcAqJCtxiUJYpyzXxYS7HflpWP/hhx45pL7hIMUFX
gsM89kdtckVtooWDD36Vqoza/eBNcq+JWKXfZLSYFn2typanzZbseQYM7y4lTSxieZdGAke9Tycn
EuvlJaDlmkNypXsg9RME69HIWO4Ursra6StXybl7plVpeoiWAv/N3/7evnS9MBgU54yuIWefjwL8
5+6rKWkUKSDm4Osg2fhcXCf90ClhB15lfgOnf7ND80Gjp65vQ/YhKrN5mEhGqtOdWUg/nH4kZDAp
7C0GSh7AczOYo1oyaQAiQ75gGzZ9NCcJRhjvvAEaiTN1gfR4x1xWgOUlfJiwjLNuWFwjhfAptkwq
zSpOrGj6358ksIJvV4/D3mouvM3s1lOHXXgLyTBVUczz/QPIPVJSEzF5QDnRPVKn5ZSTLvuWa7y8
1ISjtrLfU34+wayMAPn1lLoc23mChlyxr6NV9+pcyIkcWz4XOdIoni2UHBbdYeQwOJP1I7ZYL+BE
U4eC3mVjExJ6w0PdPY/a0qQKIAY5hfJy4MY2qT1jap77iNXdql6CDOKBkxqtN1fPW+IS4CH3636U
hpwX41u4/a1LnDEUsR1zpw+0GOnKPuwuyc2+5sUKauUo6HqFy3pqF9gwOX/VAQGKm628M0+rPsUL
PviIY4PKIteyVB8VGjyAdnw2DzFGA4jdHKEg+7n0BFVGcbWWB1EE9apVVDo7jaBHyzyXuzCIGh3b
cH3McaFP78gZLowKwqbl6KUBg3JwyDJxbnvoA5UowJu5il9f/LDmYIL8hfMGNd4xFxptPIIGsyLi
6WVaXHSQQe/yTILbxhWoHRN34clc0JY2L5x+1v4pX3788Xe/buyIZ6X4eBd2bzcfBo9pqa7JWf1+
uyHHu8W4cRvGEBFPuuF2ao8kD01cs1da7evVQ/DjEZZsu0S21NnPiuJwrRYjdAmRG8P7CeYjglDX
3JuBAPMQ3Jo5CM2IlGR+RDsFS4Z0wcMqH+RK61TUBdxuihi5EO0o1S/U9dH8iUveyPJBWJLjdb8k
oClfYPzaPVOw0aY4D+KdwX5L1fO4XeZGjKYeCGuPqaIlWh/0ufnriTVvJecU74PBvYDZRd7d0Rqm
UKgC5h9Uo8pJx5WC/06O43st+i+6V9FyWBiV80CzMCCA0sssZqni6MEYy/ZmOkZmPwadtf+dEeJc
R6zr50AN8ocVBedCiWXiAv1P2O1R5LOrf1nI7dyAlc2vzfhYoigy3iutiKrNuaAwYPxRYNT8JNvY
+aQbIEFWjaEp7tL3vRnDJBD7bWD6ZnBA0YbAM8l98Ii1ztgsR98imfkjxYRC3NyoTGOjiM3yHF/u
hgUuCxf0NBOYYd3Rh0p8P8xT+FPl2KuED6DzL/DG0i43YW/wWlyOLjzpUm0Z6cwlo74FT1XG9507
IzcRvrZqlMjx8T3QOb/pLlR+PUDS4xgR/8VumWO6xR7k3imsXSSEsKczT5zwsh+DyMxWXE+EgjFi
PD62mrx3cx1OSNIXpQe2uOTXeEQMKPIbh7KGlsZRhsdvq4CoLEFL3+tom8YrT9IKNx1E3/YFtO26
gwMkVoQzInfjtuFLdTij0t3JlP18SOPHAPj2mdYTn2sHie8r1oRktJy0JBz/g0XbxEWrWfIaFbfM
x4Ev+P1ZFiZWD9MlTGHGFH+ssi0ENX/W5qLxiokAfG4c5ceujbmPyeWQWny18fKdo13MMXD7367m
BCSxbkNbEmaouoUIfPnM8i3igNU/1lSZ4SBvwc9DfOOlsif0nYNyTsrcIJOBdhZtn9yNEzjZVqGn
hj1FF+W0yByXUL8pAv3H1QHQMULr98gRF8EHqK+nbOezju/n7vKJPtaP0nG+vPcRGgIC4PKD/D9M
mU8ovIl7PKkIA9dXNa8TP2neKaZm8dA0Ts1JaN4RcEjq53G4SLqVVj7ADSU7gPByn/MxSqD2mD7c
eD+pNQp+XW+ldg1qpCRtFzhdS212klpNo5Nxs05nmJSloO68wAhxlYDMSfp+38DIdbcdUK/Yqlm+
bwPst+0CUnTjO+dFhdpFSunl9WzlgtQXPqQc1M1mwoVsIosGTLJ/tvO7axWqR8lBr1C2lYLgzIYN
6GPDVUTusdnFhutFAS9e2BV/YUmiiz5cL/PX5aq/Ioena1Ap13tXD/TNvIIElqA16UW7lC8kocGn
5Umw2FdW2S0o9lrDUD6uJPjeXBlRdUX7mVkGFXCShvbmWJiNvXThU8yYUS2A8f6HEe+PVBGJWeas
5sLO5e2iMncY/WOzI93VzS/yUIoVikbbamfifSyU0nLnWQHfmN520DN/1Z8H7/wuCCZiRRcUVExz
puJxA4ZCQ+f+yq6h7BbzeBcutbnGz/mG8yBFIADHc0ybd4ulR8OXjvk+hqd02z3tRVWYzI37dGAA
iYDLZtddDJ+DNCdHVUFKDvJIyvnlplmQ5wwETnhTHta38sH/VlSRvEYIuiQA669xXKtT7p5Adqz8
IQ4tN1nq8ZIVmtdck2i0ZQVjQI/+50Zjlfuas+SGN58RophWP27TLvoiqMTSPtwnu5+xbrW+0g2u
5rGlrAbSW/Sp2QNdOQ3OVVdu1oTcYlnQsDgNpqjaq9RzFiK7ai5554pRWyGiLoFYhRB7XgeJRCMq
evBiZftfa+vJCXXDUV+tZ7cZRmaZ0iKWnHVR6Haactv/K623xpH+OSqzPEAnexU6MFwkE4KgSgT3
DYX8tacx/Rz1yQd1XaOJrMTK4f/XzI++TAYW7Z1XbcRwSfDEUebmVSo8MIzp3EpSK7+yhsRh1F+v
f4RBdJh5O9X9YDOXm2K8XrMyFJUN2Kd9qPGYoXjrQ/nMeN47aeZAjJEHA1zUbEFtNC5yo3vy9hpV
wR9td77NSWWdJ5DVLlj4We+M/YX4t1Kbzpq0ozPcYsjC5+3mrwITULfulO1pWsx4Weq7gR3K6xj+
HRcG4qjY9OZzoP6h0LgV6NFnvgHhJfELy7/GxA4XCmWK2FG0ElVDjO44S+Z8dMzyK4RDKmx5Dq7n
3j+Tcy1ToDk1jBsDnfVQHBbnVaNLoBKd70FrkwrFRs9dmss1qEhAgB/0JJJkO81dqh8Nbyer/cWn
7O9v+Pp/UU8YKQG9Q4L8YzekG1X8YlJghPq4uRMNXtMt1OOyPQ2OxoT441yeJhC7eO7GldTnEPwv
NloOrDb4XuzYOPkFU9SlAa0IhCVndlMi521EMtR9IfZWrVN/me5G7MSDmep+meMr1ywfVs+GZ7gQ
h70JmrMs3/YE62lbMIPPnElV0zZWnXEmizCzSjHmcUy6WwZlbD52O5mzsVGxNjmS9kCy750HL5X9
ol1ESSshlGCplP09x9e02u+yeJIo4WgCS364nX1pVdMSVe9VPws6QeWlRL5I6R6jPsqZFUH6A4P6
6qrd6aDIqxH+9LyirgHtEJC1ibUVt6IUErb+M9a5JqUOS1amG/KGfbscMF/Rlhyz68LasWOAvodB
cNAvIeWSurJkV0CcknX7zjeAbkLouslnoWvEVpAv+bcdy3KzYjIFuJmf4sCeX3lWPkM4Mp7CDx87
qlLIa7pqGeyFdYoQWYMSwwgXCpt6X1l/D6FB2abDkk4t0PmDyRQj0YGuZ4zshuytNekjUvNasUat
GmEjpCLx3KZAe8emPEiWloTVTV/R5hmyzSr2ALu3JT4TB2kp7JwgLqA6Vo97gwIPFVeOyTUc4qv8
n8jfx0kI+EElHDoqGSE322QT4mCeRFPVRDma6Svf/eFdULub5X7vL98Uu336ZxrK6UMQqdjrP014
UhkmuzA0glYVIkH6GnNmlos61i4C6Ufj0O3wt6RF3+LWq+CaFhITKNWiWIEUsUe0c+ZkgH8ihEzD
+B3AoX2aSPZQVHTwFEIR9am2dYo2aXlKeA/DM48M1ijvInL67LLe/ERPj1MNs6UJ0yu5AWXcl4G1
NvT9B9jwHnWqo4gIehL8Nptv8zQpGpDW/WAFwRcZO9JKum7S6vVVpeuJ3PDP46MgRzqKbw5fkpd9
BuECEFBUFNQ2JWUO3C9bqC7e8Au0uTBuFLhhgr9RbsTOrDioSz+j5/eqw1JyDLJdf9edK7pcx3IN
5NIOq3Lkt7pdN1l6OGtpmAzqqK1GJ1+NCef57lZ9CBadpKkSCcT6jTKnoO8YIP8IjQCLeTomqTED
gmTJOkYsNbzXOR1rJvwNyCtBsn9r6SB1x9QvHYmOYsZ8XmnyGeJ6wW2JSkfO+2OIiHue+7laXziG
kHGz19bmrPuvM8fJcwpwKaXlvH++nJ4W0MHXMpWWLTCYcryhIn62HOOiHVnc5ZIaaXdFlIan7U85
l/7V/EfAe2NCxh+pj5GeoP1i41u/VqOBe7sM3MpVtNyA90vgeKv6FKlHJ6n4R4dWcgrWvSDpdo1s
AtInD2He6Gsg7fwFP5wkdJ8IE6fJAr7Nv8FiGBUizIhlxeh4bRk1gIzqrEHSY1CYQcy60NaXLpx0
QIqkc6yH+v6Mc7Ph5MTeIbKg/MW7EUaCsz4ztNVxnhUKs3ye0lCARK9vbH5KT+0Yz9OjgVLZbfnE
sPngJ3yJYP7kYvdJlQoTwNYYZGWV+mUblGfQN8qLmM3QCNz+rr90+OL1eI21uGK99Z9/VYe+g9v8
qrhnXiaxr4tmqFTpP58uLQWUF2GKl7dtIwRJQ8hY3ObPT2onAhjVkR+4+IyqKeU9hbmAJNOusw11
iwU06LuNwszXesBq20DTY/OCcDc9iLoNC0pCVtiVWT4OD1ZnXrkDGBerRww9dOG/POHBkjgNPm53
J8SqUX65pHWqJphNAJWyW5Jgoby7YYVurDPZVwnMB1Ds6CH9qQGo30dC4kXSRcrBnXR7BuAdy3vH
laNwZTB/LwKx+sSf7lyjNxquTmYWzban5yyMJLt4wQ96Cyl79dNgBq/V6d79GNphl6NsGtai81ws
QlXpQvNbR0QkSAyO3rXUFFFX1jDCSB/F+Yi7pd5ITbfpoz3lF6B3IdhO0JfkGRahyFjUO3ENDw1n
46o67iKi0pxF9B2sl8YDp7CTiz6ozwbwncTCLelaUoxY1OwIAqo/6moGdD7fm94wDD8a8jXuCQ7b
1aWc0mn/tbKCVHzbWR8tYd2einclRQMjDsT1NyBFbCqrZXPzR4zEmR9e51U63dsWvaetLgzIIypu
GvqF/n/4B7OL+Dt3MwvtNEB0TGqWvOJCpiURaxkCurvQpsOf5oqFQBym1TJSlBoQo8tDQhLg5X0B
hMPJ1PUbY/LOffZDmYm84EtDHxHHH/NahiuJzq0juOnyLC6O1/aAzEhbh3+oOAxSmFEW+/MxKhno
JZFpRwoyNsUBDEqH0H3gEdaqz9sjkHT31rGXO9CWd5X+z7+QfjXOp52WP7SvbHxiDM3+wkHsdr74
sbQ2PwLtL90Qh28kXH/QB9PbJJYN+k04tD4pjmAU2NoQN4cwwvgkZ9S05/pHZ3y5gIBJ9sdftWOG
e281bTt4dyOYnZjZQoKVTYw6przHmIPaYGUT9BW9N3s491DlzmQROBZAQzmJEAK8bDvzmwS+7EiF
NIKBM+lX5z2Tf/FPnmD72yAajBiBMvsta6dbllBJeeJG7/EHrO77IdjkdCC4nfTVtnZxi09O5G4s
d4KrDbSCdQqVnwDyn4AHHyH55t25fXnJrmoxDMIsMeuswaFCDK0FSGDMo01QmAEoxLV/Qq5tuvfR
agp6pWt+8jUXNzk/WOMURfVPzzhjytdWEFJXO1WeHxOaepsM05TUOjypJXf1PDttoiCOQ6eo6la8
Mszb2pdxXbkgazC3PBQKDlQ2oynfNCkgOLsuxtGl1wNhsEB5A0TF2JQEx9XFRpODKp8sJIdZXsSK
M40f6fEYGon3E4hP4QUBo8MI5Aac3ez6lxvqkq2tgz/56HMlHDXpv3mdMRQ47ivzjIYV1Rg5xWXK
7Y4FWw8Xih0l1PH4sDG9tz/JlCGG31XkUSll34Y7P9G2ru/6uulctiYnjHN8xcvpsuAQOo4OxUuv
M8FP6fZfkPMzlKNk6MHgmykSBKoh4Bn9nEQHKsSgLm7V9qY1ge3ip2Hha4xRlLgdU818DW6oQNR7
P3MbeVcCpuvJS1S74dz6DfbFP3BZyFRvf2pgXcGqwtxcQkgzztm+34TGem4gTDudzAKSPDLJaQGj
U/UvwtQqz7sTXlOJRa5jhQqQgxf8pdGCrO5w+2jvkHC0oZAbAkz1uP+jIg3Jl8adSDEF/g5czcTS
K6Vu8cZ3U7oAHdMwXBTXqNJ7n6FABjDySy0kLuuDKDsN7+DVLWEkaCRHsnT83Dd4rFKOrDCCR2T9
00q0xmCeeEUMGLu0dsm/unTNYQPo+qnGfEvApDqHB7Kvv94z1lPd0DrvO0Zl5+exEr+KDD9HjJUR
9Flpceb8fK4VqLpnyF08nkPGyb/2+OyStIwE3eV8LjDQ93mw5KWzCAc80JBhDvMIHHk0xDLAk1VS
oVmKanUpLw/FMIqts7JgBizSoMwQn91NY/7ZNpM9vTwEO5XtDTCLhKRhhPA42F1b06PK5Vfh6j0D
dzW4zhYFVWnjtohGcBXOPQHlK3R8WZMh3/EvUmRPRlVTU80fgwWvsZDJxq68GaoGuaoyAgQiFUQi
wtBHn1IXE12IZnUUKW7XKHif46WGul/iylLlJKf163l7mvYUdKaLuPcGDodMJQ3L8kxR76urAIyc
swcaW7Wd1pv0LP3eWb0WuozJEO25Tghlq6QuYK7Zm1J4N5u2giRJ1ga2LPjNRfLusSBoRJON1ZUn
w8B7/OYTd6Z4lEu6zIhNUhuqisArxSYJBy/bvTItd5prTlD/iTGSbFBD9ULa3NugQS+z+C9N6OjJ
uQR5P1AiXJuooWrWDoGjItJbQUiFBUuMXUB4s8P/nOERIM48Q4mb3BLm4OKzIEmob/3jj7tBx76L
/pLVqOuxIEMnDlG1JzCMlClgHfe6TdHwKHVJGG/zOV4zW7BxWrAp24xyvj15ELsBRwI5QehBBaHQ
TPKKM7mAajnA41ta71WK+Ybe7/DwG3+4zTP4VOJnfXZmr+TsVTEkBUh5ZQzEpB45oWA3POQ10n5+
d6q2DTNlHujUViB9ONtM+dF2umsdw2CA9q71SMaBPkgN/AIbQgXpC5mzh1XHDwa/6g9Gk/XoN2RN
z+R/j5TfgB3GLdtPErOiI7XjADxNmWOmP1pHEPft5m+yJIA2GjdrKkBhKDSDLM4lFMeYTeWeXf9Y
/o43iu//z0QhtsKNZTBlaBoIbo2P1Y+zGaLe3UFbNY0OsC7Jqr1Dr2AMu0nUirQo8ZEGdsUYMfDQ
gj0e3NCCjw895LPCjAzm9YSQv+HSawCqUj/f5fWizp2Ie+/MYxS6yZ06Zi3z1EdzQGs34RcjqIgP
24F8iKu7LF0C5j+o7YII5DCiENkQLbl3Njpy0w7Ozs4hp9d0a0bh7XIqk/ybvxeGSym/CSJ4r31n
R65tq+NJ02LU5U/pjljfnfb00YPCNRB/wz6NHDMk38PqDQRytPK1kRInDY7rueIkfoySeXWzPj8t
2dZFCPSOQ/d7nb+GbDXH2Lkp3t4x0ksoBtacfJbxd+LEPCHSa6/iXOYa6fOZKmMcLZbzMgjWYtG6
d/H8NMZ65dn6WVZiSedREV0SSUu9fPw2UF6j769PrqB1pWAJrltjTsnt0OhxHWptEr3JZ5KdCWaw
NcPV/NaNtNgSKRU7Uc/wxEANk815Zc6z5VRwtXK7oMPvo95ziKtuIgjZ1UJI0I3Fbwa1S0TQsDRS
iJWIVoJhw7YP3AZ3hNDQdpwUs2f1HFKrG5Z8y95y6VLk3NBniOIJA2MD6O/EiwpKG/RPLmZ6w22c
MCU6jrWFbxgJSADhC9BvVrU5S1Bj8esrqrJZkuQsUVcOUr9GF2n1gIprSC6hWuzeD8IgVaAM6nFF
V7emyS0U4pADL2lGHU1TpDRJ+vbYcSM1Qdoss31k8IfnW6Fwb7OHrLa8+SqPEqLw699PoZfP3Xts
l/Ui39YfxJ9IAJNuoGe4srpF5qtYj3sTq+gsWIkPXus3Tv1gG+uz+NuIdrX4tDVaw3iAwbV50ykp
xDDB8+9Qn8JIIF+EKbSObxxdHyl/mhteicC6PyFd4iOJnh3s7dPgggsCKV93Bns4U8cFD+2fwy9L
miviSgA1EkNdSu30/xFz/lejFsFq+kC1BtkC6fmnLKIJipk+GB6EfXiF6fx/9/ghuWPrZYNG5FuY
n6oZxOiuPo3/08n5ExLWKUV8C3/1Nv6iY2XiiPWumMUeG9ihwushqTsF6t8oh1TWB2Z20/bvyo09
V5uW1VDyRlQ6An9WKm/gEQsQJh1EiClTs/HMNJAEqyufee7TfJuhC16aJCTmKnGlfS7VFmv7Fc00
5RN5rPd0rDBx3fs5KD0iLXVfEOCsC39qZgp6+06NgaWLXTeA29wjDFj2zCHlPGYbScykxeBjX4gj
tEsT2l3l9yD4GG3SGIldHtGq3KmW/HieCRFNkVNfJN0pikFo9az4XPw5ur+XFI4uw2csA2ibaFFL
USWWUPENVIfZ+piYXWB/IHDtkv1/2UvTwVMFEphWzocCptiaxAyKrdmtQhhim0shbB9U6CcnIlqE
dJ5/bIx29d+iphzm8SPEV8a7f5lGOaP6rGUZKT8Lw83xak7UM239qW+Wr0URChy47F51IdDB3lBG
l5d5t10YGQnh1FilNZECZCFEbo3X2PI7MG4J4XmLD/vVK3mu3qJ6hngdla/XoeerIpPkPxsPi64e
84Kw17oAbSvqiVqL/+cqF6lfBv/SjNbbvqBMUgwhFETu/3uqqTlzr9Rn+IjEQcsSNIBGmIu0fOVF
kD3K9D4cZknr3eA2jcEHQ5oBIoWY1qrAGXuXL9VISUbyCP02uts06ZbeGg6pU0duf1KbWE0k3Dza
BBFsKx5gD/BwRwQk0l4PsUnepHuZHee7pQcmVpx8nQWnZsFufLg12i9s5XGU46rFFspp8H31oC6l
JwmQX9JyUmmU5WyZ55L7yobhZ53RIJ0iy2ojZMf2XmXmOo55+jiWDUYOKNR+jX00xNQlHhObhlfF
42jGKJPKX0XMjVLVucZmgRYu7szaZj1P84cg1139nqYC6jaBTlCS5hdr3raqeTOAVxKg7MMXirPM
/IIh6FdW5PXpL4OHcApLHBs+TJQ4oPT/hhemygTtim/r0WPRM9raKYh5EAqm3FC2Lp1xoGgzXsGH
b23Kbm/xkQ2chEc+0IHO/VxMRvZTP3o5lVObdwsfivF0em57puErbbUnIpa9aNNTqWvQlO5561pJ
yghTYh44y53Uc90kgpuT5oCqFVq4UIshjHeS8D2Wr2WsN3pvNtViAW22a/lNB2MJB4SH3ZA7VX8J
XgXxQFbLC9g40u4a2JF0TLD3gCe4PuR1MRVmGdgn4drlU5bFBkzmfiG7V5uAdihpCD8XhQ8qxL4K
3Jg0U5pVi+WV+aOBxg2aMFzq4h+oLXq5j97qgSRlbJ/9tneQq4ikWcpXxgZYYz7lb5Bc4P+vFuof
1f0VlCYpkD3Hr2Z+dlA9B4WNt8d0LFko3JPqHMBviKagKOnG22YBOMSK/QoaYq22sBYMBuUAO6ZS
8T+BTsgrw04aIg/IIyyLcH8pqGTnz7rKbZNLSGQAUcl6pWR18SDjJr5nfMaCoNKxg4suM9DWxaoC
Rcxile2iy5qr5d7R9ECMfG3cCspPrxrHhxYh4DnBtfeCQMwcnR1yh6APnyCmF+QC/IR+/rSe5Tow
0rTRBfqkShwuqmEGifpIJalMjsPXdpe+0iAOczoVaac2JkW4nX+MT0kkD3kNtK2Q+9bbxkfH/weI
9uKMP9Pxscxpric6NpextudTjYzP2I72swQypi6zMcUtxMiqunnmoQrIqWd6PEaC3r06fRJwqn9J
rxM2IEXbCuzMIsdBbs2qyeHzVkT4aQ6OMFhpHcFVhCKZkUy+VAynvtFkgQ/pO1XB/MleHHkgbSeU
HLaiLnwID1Yrn352zLBdEb2jTO/OcchEAR8G0EG+70EjAd2kJQlwXFpswfkvKYj9FYBXp/Zo4xhH
Ax3pKBRZ4g2BotANV5KnaZJfsfb/xzPeu79X7JmJ5mkhU3raWhujJt9nPlUU1XivS/cWCYyV18lu
CHualCH36nV+DwaplP5h618Dm3OW2ZZFbI9b+HOu4R/gybhnx3Se+SgCILDyUd86tdyNBE2g/urU
EMdlRWHjJ/rfR+j65kahGWDgRwwfa6ELqNo0XdcVCt0qlaUfCYmE7ejrNekfToZRSP7EF+DI2jL8
uM1yV2JogPsrjQRLPdzL9m9HeurtpR0OP8phlls8Ms3o2IWHrTUFnKyb8uWdA0xrMJNKvOem+YDV
OPsDrn3Xetlie9ZK5Q4lwe0xTJ+7g4bqGSCRoOpnCvDc6vicWGGOkYnLrleYrQhDhqNixnIi+IP0
+2b/ZK9jJvp2Wais8hOlVHg+IXmHBdlqs0wzuas8H1W5ug8CLVWCC6zaiHWRqLyPaMH2ni+xbn43
sf8T+LIMPwnacvT9QMGLk6nDNOckLr1ZinhSYyEcXRLNodx/fcIaModjTbQ/uhu14Lq9x0FnFs/d
9wnPYp8aLuOz4mCGd0zQ++/rJpMMRIcrmmoy2SKGB6+piYzRiLCebRxMB3KFf/y8PdGvD2nCSqsU
BwY7Dx1LjVSdl7HGGb9f5yIdmJcQinYEEeYuPNE26al571C47jHvLyc70/EhWBtMgRaAcmRgjpmG
1J1m/BDv9QBvJMU1tSC5SPNX0PhEsm/BSNHEOjf8o47pa2Dmn0FexvISBY6B/EAD8G28/Ypa2zvi
nfxNI52fzkr60oCfo5YTDrpPl5H6Fo8SKGsectzzHgOPd2zDDcf0Mpd1ZAEijAPZ5yw3EqOiCYq+
srvqxn49GQeWcadwYEOafENIYctsdWwGWZCaoEI8NSsraf5YQ4TilDnE1wa4BNpjzPHVlLJlQQ+b
rJ+TeJuQsLsnqETbioMH//2Wlvs+FMg9S+RpoTb+iiE/J8p1XvDNCr3SMV/N6C8cQjDm4jZPuiJE
WsgAaukS9jkw2D9sZhMHbpLwbMqnuGHwul9GtMM4zAyIZRcNmvSZXg8V7CgDWEi4vPQvn6ZDQlnI
vMxBL9pGWChpkMMG1Nz1ZWipxT+x2H+bc9f6udUaRMOm+STsJgiA9KMt1RWC3Arx3xPhuABpg5QR
W/ldAoaSSoqZb08UkYNPXT9hVGo+30gJIkNWRIlr0Xd9+VoNZCl+w6xMf2jcqThB6fLJFYIVoJTn
kp/ROZXaW9V1Kr6XLWTE++Y9hbNKWQCmhwVNRt/GtKVPhNEqi2T+f7HwK3lxu0H8U27xbtYU4zrZ
WzLuli9GzkoCeGHLw2H/hyQvICGTM9Xg8NXGzHkBZBd+uKdJZO+SmBSOz++biJQ1qI4uo7bzx800
ShG8/suUiD67c3O0o5TQENdnL09/eUqXOqCMGudUuema8FbCTVbgxMFX7ne2tlNlK9mpxSGWGg1q
APA5Q7X6nAQViY1j+y9RyUniVMWFlcuMxS7wxK2je1EON9bAGYdlHthRiTxEanSXmSstRJLA7woU
7M4wrJRpSN9zA4XeN9Y7aQTTBEHUdZdRAehjHcYb92AwoEaCgf2HQwsFmfmraVFRsuVp5bpSrL/9
yvZwb7L5+L7alJMaj+j+WagM2EQaR7yWqm8grtcKJMtrcnfFGLxlCavtu7THXVrQEqt5PSOOqxce
T9kParLOz1m0uO5eWjO0T6NcGwKMl+9ymRv8quiJsiJzGiNyH8XeKbi55VzsG0uYIa3CFnumizSc
xqUtCXXWXRTQY9I2hgzlbiKnopf4vGMvFL1fMU9d/zSZO+Ot+5OBE+kGH2nyEyLtCOd5oaiF15G2
guvyZU089yQO8O/e5wcw6loyfDlA1zNJRq4CLLir5cTvPIVC6vf4xQ+eJl05z22g4bU0NgSRvT7g
8OQUSAYBtNht4k5xKXf7cIGTMBxybAgJKxgI7KMTs59Tp+EtJlu3VU8Wx/R/zoaow/qiWJQRCqRY
X836Sgf5Bx1qChZULY4Sw4KpX0J4t39v1plL/NQVVJVkz0R+BsqbKpLqq8pY7ZlsgIwsJh0X9yv8
6v1MC8i9QnZpTGnqMOW2ujXhyqvctwCIOpTy3kiJMP4qldqei/bTiADu5uNvtsLp8ihAr+a+WCm7
woa2UtObMCCspshhk8UZ3q+lLWnOlLs1y8GLWT2WN/BgDhG7I1ut2oVg9kt4XmfuIL5UKEZJAgPt
0WRTpbUzSEMoahVciK3aYOnxdShwGrW7KaDvRilXisIjc5u4bU7QrkRD9dPJ+Hquy4fd9CXJ37y4
2lShK/pOWsyUMO1k5aFsX4rCrR2bh5e8D6ACWGLPhpj9wtz36bagyhslUhg2Mj2ZluwLkermx4VP
QHhpTClFNPXOTGd1gRCS8oj3zkVo6+1Bzj8NqU/aZkhOWG2k7Z/Wsx5uokY33/7Lc1rUG9fGtQ12
EP8AAIxn/HEvvXfvN/BdPnmd36NrULXjM0YmAR6HVUDnSRUOAeC15XQKhbw891+Dk6R02Bvu6p3G
WAHyHNWho22iDXJPJ8qGtko1CQ1wkyiZ2dQZA2kpTqTsZIgIQE2V+XXSuvuQfvGZIcMev5wKvi9W
Qur3/ERR42J0qWNEU9Ay8wGf8WGUppgUBO4LC9pFpD/Lr8P9DyGcR/yjpfnT3i7IBZrb0mhWuy+h
HyKTc7i2b9AjS4x4hP3uAGXJ7mcyjPS2+tVM0iysDVU5qjpr7SGO0sU4D+/GOtR3nJAgZV3a/DaP
q/vRwCOfQlykv1mWBgaKml9welCYod6WL96/bgeQmGUtuWZLGIeBBFYNvpGiGtbQZ/U+tTKIk/Cj
djiGzw1NQsq6K3Fjbf28yV8r+lzQ+tyaaBiMvcxxZyAMZGogwgfu6tTUIEKpoR4NxrOYG+AO0kqU
8Fe03k4lB/zyaOnGSjY3feyDAbzkwOaUROeMeJGC4LZdunlYv1Q7/CanRcCl7Bv0RrXfMLm7MmCL
0X47TFbMdoLk5HSMOoQ4W6/gLJQ/P0ezL2cKtEqkkZ+LldThMgKnC0bj1aHKiZedL9+jFqrw1fKA
JCBgBAoTXr2hifnEn8L5JMLmW+sdYoxvz7seQ6FZdBGxuFDo7uTNowFrqudiPKO9g9Sje46VGRn2
tKG8hg3Y42pBWjg9o4+/s5uOAhuD46+vI25HufdLYVsXpv/l/h05ptwPsJM737oOvOK/jOcUOxGx
ckR//3iIz0zSL4rHQ632SXc23prxp/eNAA7Ruw4Kx5hVnHTQjUVhUFDc3JvD3vKuZh3dkwG5eIes
MonXe0ufCwx/4bSXT7Y/SMcZgD3XdiiIyXBDXhTVKL28Hdb7i/RADBkAozqXonaNZI/jzvYkxI0G
cGGt585gJvoHEJIaSekJsSfmqsqyKobmnfkNn/Wwl6xPoTtPwMBLk1rL/WuJQUjd3v9BSqtYsIWk
Rk/N4c4jHr7R/a2cV2b44hHYTYjMCnP2r5IUlG/I5VYGJYgvUmyq/uViAiXDM9FdMHDuL/lUgb3Y
XOgS1QMP1eooIl2P3yg062yZwF+jlR/TtF9y2IhU8WTrLp/XWDskBOCBHkzYpwK+mBkGbTwIGM0H
E0O7iMCHdIz1hqbsg15NK45yhAx0fLjly3SNz3zT/jghYai2m8PC3QLXVcWgCQaRUcxTB35pXYD6
EEmJyigSBa4QHOh9AQ2CcrvzU7zWhQaWOMzJvLbZbtMs23ugIZlXkm4FpS4B09tQ7/T/VIkYCbKy
fnLIFi8QJQRYBfNPFV4Y2kFBKTy/VY3+JhNcdwjeEhwM8UGZEMKblG0Hb5Ub+DG2apOWsFhnJLqT
DALPTdiGnJ3mIoWstNxPr4Ap4drP0TCi+xvp9I2Eoz3ttNaTHs1EzxZg8NMf7ZrNoLFbIc2uq6uh
BJbD2othaN4qbnlsCLHK4qqYOs75pY3gG3lX7loMuQ3O2IaCVrQwYmweB4nJS4yyqAWvS5g/izSz
ViFcEVskFOXrSQVvI2KhKaxBHSXYqDBCujUTrRh9ug5KKSQVD/R07GLkhr9SphIyo6KTcMSNynJ0
98+snKCwxB5+k3pQqosW0+2mQx8Wa1voxv8yQOpf8ySXB6sDyNJl29DsbX9l8Q8SIwgccQcIMV5K
I/sSN54qauOD+IG4fokzzhkkfx/Mz2PTztG5Duw7ib5jfUGwM0H8q8MI+df/ljDKVRzXIIb6TuiQ
b1Wawotiz4q+ISJbDXRXtlBduWneFdp3b7GNuxS2wEez1lMesnZfG3NVkoW8EkjOLFWNO+6JDYZD
IQO56iQ8c8urK92hM3KxJg+yx92c4z9UVIVgXmjhfUI58Xj1TQ/RgeCVz1GcUChyELKXfTVm8C4s
RuoLSex7uqxvAjWvYcrc1qHDRLJ698nHZlH9RwkLDm3X2cG63Dc+6GVRyHz90NV0gQE0lYD6VNcV
TB4XiqaEIVKAbXC2T1A5mESAFqSjz75CyPWb2HqssEA5VkshTY3z1BZTIn0fLnffz8oGMdB2YXQt
bCwIACs5JUrMmlHEe5zyOBze+2cnTnGk2xswLmIUlB5OoLhtsqPaCf/n3gYjT1ys9msn6JGEcDSn
5OE51+Un+HrU5CmRmfd5+bt51clNY09ulBOe/Al/DMyZIAsbhYaolzePFocq24mZb8ZKxj6DiWpX
jKiTn/OgIQpjWULA3xRad6NW9D0lw4eJEOc3w/0PkbTPRkWMdrw7z2QiNWhAALlU5iufDOhqWIMG
t9aVDtz8qcpgFPz1xucTz/vPnrtEYnPC8dKrlNl34TKp87pocVGR0lOBbk+sP3uJxHJUc+1eLxGw
1WKbMvqseUuj6Sp+ghovkBYMATifSo1sr4MpEgmKXrrid6RjgklNszfQioI4vfPeUXApNa/g2qUR
DBpVnosXKlV5D0ZeG25Z8r+Vwace8w98tfs7uqU+JD02ffY1gcQwitUSj8K9tQbxHc12EJvjBvEL
faO/s+C2aaoDcMhWcIibONwOf9xauaCenvJ5ikC9RhVXHtpoFT+qe0AJbCoIfHT0ImjGI2yWivqg
SCxT5KAZl+f9JhuEvRya6GcGvYr0Dw8Mo0ZuvL/8Qqqn4rGQ5KYlFzWWlCb3ez/roEb5yPncO6+C
WHgINvEqeNODLlgxGRpR0ToIcs7wYkQBNozNTOMg74qi4DfeBd3gBAEGJBI/sR/fOp4H+wyULqki
kp79bh/dS9+zvXnFZJ+hA6FoukFRWdQdEpDfDh6YO+jlTUv8BQHJxrsT9ArQMDGBl8BjSy+pacgP
3CBJSujLcyC/0N7GT4AISpvRUJHmwAGDw2RTpt8CSUlFJxBBj+3jz9J7YxnyVwUt86JxDdWTnJg1
Ro+l+dTDTgRXoMGFt07654cvvHs9K8DD7IRWAA63U3sMUVTZZXYpoJIMMQsvRich9ftgEx2hFazY
QR35PE3qofM7WFi27b8jobMRsGyGwI8fAt8MlOF7zi/Dv75zQg/eFp6uXKch2MZRgASJI5edAPY7
Wt+EU4fuNqEdYDEIaxQvxmMlWFfKYvDwqMek7+sR5eCdSpasuREdqK5W6NQ0niSA5ya7CNeK82u3
D45RDLGX3gcwnxHAZrpI5hncJUf2kCgf6C8JRj7Fu1H9fyIbPwlK3qAeKbdjddGK6HDT4gQd869U
qZY96YabpKa6qK3eCsVS2BbQ1WNfxB9hR03w6/mc7L0DviO3146aOqwqn0ehUsouwq19Yk/ZzXhS
jrmrtqfPnDQqdO6kYXezW5WZ2NLemqUT7WdAa7KiHhJbwNYDmShoDEvs+aojXN4XOG1uFguP6QPe
vtFCHiD3S+r9mENZUwEo75PFEXOFgcMrDxbQ1Eqj/2wPMPVShcE72sMB73NsaCnzenL6S7G/hdM9
I0X8PqzjtQwwyELoEYisXBWfO6bDWir+M2/N8TT+W04LiWlUob8BylEYR8ddPa8RX1Djj0NL8JAN
20yyn4afrdRlJ6JT59HgMSln/UpPR2hevk8IdnH8kNsdS0BFn8mdzwsFekcKy3hJ387VKOUO0Mf8
tZHp+hVJdsPqo3JRblOt/SLNBfRc2AUPNR1yCUsSkB+EZ43dQShQ3oIibVGhLjT98T8kzBVmSat8
cVfpyq7yITrxbPAm5Yel9JLDos/2x89t3j2l+NNVvu0Xj7tJ5qAo3uTlYw9Zcx/ZLP+7EMPCWRCr
FURKyDTUfFQR8aPhK2DhnX036qtnfttglmLNbJCvvZeCuxpjk9ojdE1VObshh8ESigq82a6Coc91
L/3lX4qsBiASs2kgQrCqoUDyDMvh9/9KAR7UT4QmNuTnnHYIBucxbBa0+JMzriJLPBRP7oYXmpas
sdY0SCoH8O3eK0Y+NCy7OKfffLY9dnL135ojWtZAp0GR5Ok8V1tJ3kgqwFWtnfq9DueLjsnjSlSE
QZnoKvYh9lSFHMyYx51W29R7HkhRpiVf6/+BfxzZ94nGwD01xNUkLOTDKSKS4McGUPLIAEoDO7IC
HlISLzuLEDCdRrlYO6vBJ+fJ0NVHtRymClszcfTtFHyCL6No6yWPC2iol+vMLca7fRMaXWSKVn/z
vrhFgsxy1c0yoA4cC9cfvELpaJfT4Mi0FNJt6UrJseSReLbgVVhWcVNCuM7rfqy8tQn1tFDAKqjG
7isOFlBiqw4K2N8W+mrrtuOrww1l6Mr6akMeCZ0EGS0pecvufj2YLMCP74ht7jBqJNHNikrFUakn
zo6j/ujTB++0/e/nKg1D8iKKbYxkGEEAB2J1gipw0q5f52BZ7hE0qjWhLLULSDiBTkAbneOuGnX4
v3XYRnGU4XsTQ+ZUGScexe8cx0IQ9/GSRgMjLmzv+reYwvgPBEAnIVkCqbQQ4mvq9IE0hmu+zpnj
RoOWcfv4nzpbBdPW8UVEqDqPeD4AXbaa79Ck7FcrN8Bu7gz//HTQvvk+HOrzdh9FqOr7vKoqMyqG
ZIl6hOOEe9t+PxrJNmXgchaKKLbfr/LN1DzsGYBbMdy74WvCcTr5el7hIt799rAprGJpQpHwRo12
zipikK6ipB3jPayNj3N7XikbkJuWK6b/oP2AB9ayu02dH/S1vH6Xa5iwA4OAyVdZIhjN3/VXN6me
6YBy0ASJ+xi1m9mH4uVeFMSzPIQZO3CvCZdn6fELA6Rp4nj9+py+tnO92zbhbSeHBs7CxfsGqrnR
zXee4b8Q059RAvB1h7dcf8vUh+Zln87t2rzHqEt6TOhx+Q8htvoCO9qByt02LLHWVH94HNLvFzMG
PbDPh7zlgu7EvOOf4ghWyqdiXpW8fTYF28iAxgV0qK1YXWS/SRSbSlzXR5dwvHyJhG9flEzgfbqW
N/cDpmSm5ECdauTagwi/YG8AYOYftXKIh75MBwq8UVgm9hD1Vj6XArp6jfaj53+kc4qpgLSwPZ2A
7Sb4ojfkn3AXlBt8CRkEpp0iGNQ8RiAOGxV1ez2VvLphAW7OVsV+HPJSCKaK8bSvWQEblcPdkuzG
7dbegTEBV9xSI7eYXNcty9mVECthalHw0eGLbASAeOlErRxzlHuk6tNVKt2mcERn0YW3EBT5Tsh8
qNkVCW97qYldsCBVW2naaltdflJd02q5Gzd8oS5BCFuXoNdUn/PGkbqD9EQoxMQEiBs37ClCyFHU
WODJMWaWvBwTV7EnmsNT4u+AtpVcg8VSPuI9QFr1ndR+p5Ruvy2vCvfGk7j4Zv8HUbuLodZUW+TR
+9YcpcjzHt58AB2feP25EZwBTlN6T+yqbYlGRmd7uzWZbIUvEOfJHibQq5GPb1F68IKhTPBGnLKy
Fh5C3TUCWg1WaCNoNir2gb3dpzWaKg2McaLl+aB3FvRZdKOSYkoIlBsalzOL/md3rsECKMUzCQ6h
GmKIEJR0iMhH+P/ZftOp1mQFicrpIGKYlTR51G69w3VThcAceUihW8DmYGgE97TCsGiVQbF5ukuC
06qYgVjTCiQbNfAf54PehEn7BL8YJ7GgCKJvBOi63gOE9TDydXXRxFHTzn7C6ryBiPq0Ee5id9s9
xWkAiuCOAytiPszUUifUgidEr9Ryhw7DICv06K+iGCJeRzRs9Pi/r4p6MPKzotudBYpl2oRYty+r
Vb+RdtD+StyMCXywJBhvij21Ap4kp/s5VIAKXUXgkyCjF0LWuj2CgRiXtb1Q02Z37CoHhl3KaQqt
No9j+QS2yU/7b0LAf+l64SoYgSfqkq13Npjus7qsZU7v/ozWqzyVrxg93ODzMcQu0ZaaaZ8r3tSV
hzhxdlzwtwc5jFmeuIwNZyCVyYgJ4SOOPH/TYMilKDqYwjk2Ce1uaZhp9gHXofp7ymQFltccHVXp
ygh4s9vdT4Cr+y/1zkqOAFyY6jTp5Lw972n7nEyD2RJz6/ms+RaVZ3XKCBgBslBpkTmyPk+z7UNy
ctlCYM1Ey8ipKg8ByZu5d4w+Y6pmAf5JlqqBqxv9eXnIek4IOulOpauPU6qg8ttnuLqjLlt+DJ1m
eVQGGCYmJeoh7UWZnY8yKKe0x6l7mf1PzKdLEpuUJndh2NWqr+QGyv81XRpmCcw0Z7uczW8BAHMg
fXdI+2aCJ6OZdRplaWYrlR+nmLcwks/BLIBIlgd91FF07byhV0VziOJAts8b3w7gYNv2DAeg46L/
qHEqup8am556+UjSfOD2Jpv14DFUrUOJojKA3/nbBuKKS3RVpudos6GazTF7kGO7rJX9fCV1DGfi
T9dJAb7KecO99B4DLmZjRaIKo5nWO93AEYjVumw7p63RdgFeurho3emUjg37vDsI/Prl5LRU1DoF
s8TEj1upXBPef3Ze3ZMtLJTX/OqB7EMIzcGh9KYH6z4OUclFIOawUkh7eiPp5m4sH4pL32NAHbuw
BMSFhalYl/1zrOcgUXM+cErNtmvQ6v27xvRG4K0MxZyGdmEZ0zpucF2wjz/XRHZapzbvlKMNIEiy
tY3TOLKXq0cVCLvpgJwTKj3s/8jFr7kcXAe1rbkTH2/pW71zqFLKTTzn/cX3PQXOhNEplOAQo7UF
Jb1DpWbXJnbn5C8eaj72l3qteIOqTX6a15eP4ZL7CvFKI1vAy4XAn50w4pBGUpiXG+uRHhNVP2GI
Isw6MTFZ3Q+2zD6T31DHdR4/TJoLW6gHc0WbeJkn9trlhKZrZpST0u10AGSauGgEc9u2qY0+Ilki
C0YeG5xc6nKbyZ8wsJOjoiKjHmedpViWfCKrBfPzjHPKZzn3NdKk8EoBUBAmiBsi3n8+TZauBfNF
jKtove1FlF3dKOwQbfrXJBfgtFejnF61Bz5nj5zrP2KFgjM0WFeXGDjvIuln47GaNrANlONxrXlX
oU1sj46vrSxf/bORpdj3PIm9c6MT+mfbnO7ybT4J6CitKHo+XyMzoWJRSbY2iNJ5L3gmF4HA4cBd
ATvj0PY0DXVu3mzRa37IDBAKbB675NNI7qpZfV+7kh4PRp3WzXnAj5Hd5xQoJ3TR9oeAHhalUcMw
wto1y9NZGT105E3RQy4X/ahJXQxuF2qPB4Wo6YNyvNZcPz55Ka0mZqfN0p3JXNfdHbQeikD7/z05
pe8embCc5Oe91letBfB7XC6WaW9QHvxOqqaPRQNOWvIFZ1tf953Qs9XgIR7+GwB5zS49tnYcM3oF
/+b7D7J7T5s3XQNDIYIm2xbbHt1hf+rPG/KAkVgTb0Vo+K9QiV6E53GMVnyECcUq54ElyRvecA6h
KOGrHYCZD0pPMp13kmtDP/f/oWHYQiqbDlBXzQootha4KcSZNBCYGK7yRRcgvcZj67c62PBxLMCe
TUoVIgJ0Zz5FsNoi2adOnz+/KAvC4BDmDUwV8gzo4ZminWVsD+5UpFCdo1FCGfN2BzFBktIgdp+i
lZsRLeNyibqGTqKuDLVuCqv/8FqPILsC6Ljt9NwJqDZDdS8HPtiRQ66XfI2SCEcMEVWVlw5n/zvH
SoxtbA2phH9eFtW4hkjt8fF2QSgIIsY2pXflmFZL4PKZTGM1mx4nIPLhSebgckiUzO1EogeJlNfm
1ptg9X7nK582CljSFnB4RoG85ZMTDCZ5CHvHLfq7kG7xaduti5cNSdSzt2SZBbMp3Hfag+Q27qhq
+HcrLP/DphyYH55WfV6gvo+5VMgDoAn6XBEInknpEjWy2/aBwf+boD7xGS7uDEqfrHPOz2VA/FGK
JpRmkn1+vx/CnL9GGZzK+ZyMspRiej2MA6HmASA/9LGESWoMjpWLZiSOQt9TkjgJfWm85MlCfl+u
TK9OXblw5SYUnx+HTvl6nRw/0M+udFQZYBarMoi7X52aCgwlf0Akb9r5tXdJ/i/grF33nyCeRWxa
3crInsXLV0SYE5MS6MWwvcO7YdOBgOr99yqt2x7OIzAns4cZ5aUk4PcVxXSxRW9BJSy3D1AMuGxA
D2mBrH8tQHS3r17qEuESsLMifB7pc3/Td54VN6DpPFzR3ad8dUZJA+fRLdbxFWfJuIusZWxT97k+
v8m9MOv2oYpcvZEzwPfRswA/tOdYIbVrCMX4ljvsuyRk4x2w0bIwqb6Mwz1PZ653xNJuTZnfP+t8
6L4F1qWCp5JHROFeRiUk+78JrC4+MTE58rOXGvkbz7LMrcyYMXt4yRJAXq8ydq4vsFhtmYdJeP3o
K6VrT9CaL/wte5BsYvcZhFzY7VuWxaZqaEKNjkhEBGcG3GLyM9TKw26aa2g/qOl+jiE7BPbRNohj
0zfiH+kXvhEF3IVZOwdm/NBOPoEpJMJxRVGb50NCrT93nbWEsxRSfYFNdQSitEeCCS+c9wegIMDo
e/j3JOiks51fDCi0L9I/ZLyZWIPDNEluMLHuv3HG0FTpIR4a5vFnzPXd4wOJam9aI6mG0XfMW6di
9rEf2p8oFS3nU56B320O4HZjg+slWXTPnS1Ep6a2q8x/BOjOMVOC4oQpu2VYvBU1vzphyMU7UtvT
TMCQcwaLhJ/gcDiI46vh0Q5L2IavHrRS2BcyAluofDBYiFbn/stZZ5Q1wUVuR8SoFcDKjfeUnqmT
wDl4mAwFIouVv/L+d6ozZm4wDoHBNfehUY9AvS+3lXvy1W24u5w4K0RyMeUATRs0ce/Pwgx/sDHG
pIWB2NJHJTte51gJYQ7oHlrDexniB7gS9sSKkhaMW0Kw5ODTOQhzyWuh6AbzRLPUTj9FO10KDC1O
d/R1OfkEr9Jjo7GXXF5CrEY0XNo2MgRj50cwYQM9O4Gr27D0ImhNJDJhk0M3+bcIdATv42Pmim0u
wZfZ4szagCd1l4KdZngfpap+LRQvHshUIfCh4DnMsr12RQxDXK5uWy5qIFGjU/CP9lA6oJYV4ezf
bsXXyTYwLomqV5EEyFyav1F7vBl2G/0g+SvlqWddi5TYDYQ/145CEVpknSLNgG/l2W3A+uMw02QF
8BBb4ZwGwnIehWX346SDt+aOCqFcxcNa9OVvuPER+CdmEvWKer+4B3tmDpX/+7iFhD6A6gpRGjoB
dMldn6nC+gkAEiYgfaxcaDtLznIN2cVu6pVzWy/rIzFmW/fLQsK2QhJud7WVcN8l7LvKsRId/N5p
vzQ5q4YhGV/2Oo6lv/8PTb9u1Kc0Ru/DdVs1mMIj7GXcVb6cuUnEj8cbF0CXczPP8bE02bgxC8x5
SqdAFmn6Nxp2rlQclnWZR2VLP0ZG6/yaB0iMnp+eF5OAFR4I0hpStevp2T5bGJBA3pM+id/9QIgM
8qG56JLyu9Z3wWvkKiTX8AMeKPISGVgnk25onkAD3lG94BM9d8YoqLzXcQVyHuhKQDYMya+PCZdi
i5iE2x//1gE3o64/zsPycYfR+/+8n+Zb2Ez3IW2uzuewMe7NQgdl/Xa+w6RIYr/qsgpzkf8vLIPg
0CPH/7JTYDtK0hTMxQh3/8ZxM8F89GU73HiQ9Jv4rmn5JwVtEQT/dk9h9WzxyvervkoAS1c1E+yI
DILdtZEuwB3gPGKCFaZHZFJ4vQNK7nLoPNuuEu5mW6DBd5yoM0M12AB9t5lDOI4vG1/jKiuSsjS7
SEdKiOpgyc49EDjg6RY5aCC/52Uddhh1TT2gMTQ7tP0KS5I/FhjA09cBFMr3Igs8vDNUDSvArdAc
yTORlcmertVMU36oyz8OOZGDIlBwUhvncw72bcDWxXgKO873q+hQElQr8wwj30Lye+S9uL/vlUvd
WnRR6cG3n+TBBetx0z+0vSpEhQB2tqPNBDReDu+f19D2YOy8OqTKx7v08S+prB6Hqhttl6/Foa7t
dEWp+lWO2tN7zh6LalV2opR9ToxO2vjsMxAEBQmrdk39rhF4WldaXbar51AnVKCrAKlXHAgxPEBE
l11J3YCtnaxL6gmzVVe0xz9+MvERsVcP9ti2PljRNukk4TQQAwDe9i8GiIn2b0+UO9HWpghQDmX0
KoklsHnDRAmK8+gzre5ceDuLaLdkZg4WuCt0ac9oaRlIiN/UK0HyInW4YOtEAj0/C1uYRocm7hI4
PPNCeOr95PWHu+A/wICl00Ul2MldRDEeWt4CfjRaNuJT55hoDSF3jwGxEYxJ9mE9dG1tT4ZJ9Q5c
ScBrAEFCVMxPcTEAA9lgAQERB/Dqe//uGYQD5pABL+K3eHjJ50onTQqnprVU865+ZgQ1CIsy66zf
YftaRogDoGsujKs8QSVRvEfZQebfhz55GPGvjz0IW6SMJibd4X+BvjjT8n5Hi8K9XtKx/Nir++At
1ZOfMH4oFKUlNI6hFJZucdmviyHt40IS1/vK8goQzRsGvsPWBsekpvvgLsHW7omCgCmAZeXbYux6
rtMY9Xq2svoiMIlAb98FOQbCeRJSDbor1RY3Ou8CRJlI4clm5CeQUiY6Yey2jJvTpQFUzqfI8gm+
uCHs154ECK7Kx7izWCC7g9JiEur3OaReRMZVKOsPuvMX2AFIigWTX78Cdymj8xacrsIzQWFNiTy7
LsoTb7sxapdBr2pskPua8cY39LZEFxBint5mptQ7DETjyJpJGCWe3rq9er/la8wKgh7kKmy4LCIs
q7vJcu4i3B4kgcbdGyhyS2GCL0e8lCrrYQGljHod1jOIMBvCkz6YXUJTMFTbIOKJuhyWyOq4siBQ
tztMZseGrvfWPXCWkC/0FNyPJER/xTkTPHtE66BHFOjn1YVQ70ZcC+5OvBU+7US9nJl8ZECGMw7b
5LZIa6XTE3jX4o/rI9fluPBtN3zz9nsJ81azgys7IxcYxnkey7JqV3AGFBRDybKEuPY/F3HN1Ty9
tvI0zNw6Kn/b6PgBSPqbzkEzJQ1zOveslXgkelFQzhV5Hy66ooSWfH/0Y9Zd1DBCtbS+LxdHh/Ei
P4TTrpDmHAxWX0PG3gV3B0TTlnm0MN1oVoafiwU7a66f2iMbzCn+Ti3WbhjxAGoEx3kHGJHpPlXl
LZxv2AteZF/0OOHaQ6jlK00pl58NmyaiqjO/AEVPkFSfI2XricwAK2/LfpqC/P1VuGhkG77C9ByZ
DsyOoMywcjB43Le947fT9QpFjmK7gqCC7TdwHxvL0NoNUa4to4USA2RY0YDb3KHUzz+jSux4AQ3B
aThNUiafcVuvmETl28rtv0h20N2PIyWmkpr6ijn1bIGK9SvXA+wD/O8weJjTTs7ULneLSfXyU6f4
+KKSf4brtXKk7djpMrqptqTyn3XMAF1NRT9LtL06lafaUZ2MdSVXiG+MIU4ooqv6wVGxvN1HiZBm
jqeKzvOfz5ctWZju2xM1FpvjaLPGCzYoYnJtSih6CPrFwUTj4qvAeQ9ncvne+xUdQ1uD3W01ud7I
38EAyfRCw3h6fHks8zaTz1VlKAL8IteqrKI0H2tpvwTUKURgmzdJZBCiyCDTCcB00U2992wAYtnj
1xMwFrX4pDkYuCOzJAd48E/iQj8fR0wa0kUkYe5z/XzfvJLSqI2kBsATK/bESx6NCMpERDsuh+FG
ct7NFNwmDpbzZjTqPr+GbGosbTsBp8KWJy5PEghoU+GjDplceWZZr7SWtBIM65DMKuMi4FbU2oUP
c8eOtF1GDCNnd9Gma4YGauJsdU8Dh3gD+YrD38TJJ9y1Fv1G1dRNZpZMkGEpMQaUyTyu5kTqWhtJ
cLJilIqdZk8fKRWipgE1MmA1gE7v2qTYEAxGuL9Q9BgfwvK0KlNAcgkZhKQaAkpUfyifUGiAd3s4
VskinNwLcbOUcarAfkDvu3K0m56tza0xXtJBrdIjo3xde8cpbNM3Sv/W7N5f8d/xxka01saXhrUu
i7JduzdTSnWUDNadpOO32LbxwgMM+qQREc8vsREci2zKKdQf1Fn2nKcK+vtmjkpNWbXtloFHE7Ic
aFgXuNpzF3kiVC3h0BLt8dxSJ6vr9ACy5izt9MPEeRuHdvmEcup6w4E61bYpcyvHrsxa8EnOsLiV
0/SmCkPbqUo7HaM4+UdqhqVoBIbABZm/benpRQ3L9z7QmOQ1zutzD5Z7u6uiVnUG/XStT8eOhJDd
0JXXZ6r6KSjLngWp8jGcq7bddgXUgIPsqaxmBNIWhG4tegvJPfLJ/8qCk7yCYvb1NYTXh4pTO38V
6YFSqPQfAjNeByjIX689x+oRFGi/cGO5reqzQ/u8Ox0b/TiYM0mCK1wmQDwfTJy0KaPiNNhvIbUn
i0DfUPG0VERJMwH52egOGF8GNch5mFmdcFztexKPt4HqzANfq8eEIIROb08gGXNzBkVxVdW+bO3v
82cd10WIVY3aNo8LHMBXYs2DudXn1PQemPPuUm37toeiWwOfOKYNbiu6s8NLeZAcTRJxUREEd6Nj
kwGmuU09f53Ggr/tjYJMNPYd7mWP0JPOQzNpsQe8eTQOJhNcUaFvHI/2t8nTXuCORrjFI+qOQTrB
f+GZ2w+XBs9LB/vOGSJGB5BHd3Syb2AArtE6ytViqWSZe5EBsESXodSzRARwIiiSIviYoaWCLczd
bzBac4eRFOsPco7x6X1HQ8S/84FBqDoAuYUW35t3Tf+r6220SW9i0YrhxTD2f2ET7OU57LM3ynlu
WmAedk6yxhA0Bp5a4cRINJs8ZJI+4SE/0jS2ZG5n94/y+lDhAdcULpX0LmTGybldrQ62JBLjello
+TjObxmA2ue4SyQ6H6gq7KBgZQNCZi/Mq4KBkl4SOuAGNofovzRzU6jeCzonnDMyCGbT5P2P9yxD
mYAPDhj7pzuJ6dB1kjug79Rg2tC/h3mSLRXd1OBmr9SKczdvZl46Sj3QuW9VR2GbOhZ3g0/WKpPa
3qLQYyWY1dgY9jsimlhRJ2Qn0q8gcI3KrygMP/rGjzGicNpBpAcJ0zxDqcbXlfyvNLkYeie5FPFA
lKg3GjgnKiD/yvWWYR/kQSVZVhPieFPrMEFL8sAMP1saN/KAvfzjgGotwwF18Z87kNxp7ZNNW76k
YyzsCY6xVyfatg8cVHkTnuc1PkAURTEmWFUcJ3xHGqUhv+DVLCku240xDoQh5jhzsylzPQYgswwS
7pwvaHGRnMGJeYe0kZy56nLFx3ZqRfZ0Wx9i+hyNiSAOBgqGjbBPlCJa8XjUEDJsXAOfvwPHBdwC
8giGepxunG0RRmALaVtMcaYjT6lhKE1Hr9JjyGKA96w/68mACiioUIfTIEmvSbxZ/cWbtuOpbWeZ
Ay+X76aW+Qntd7twepgDwq/gc5YR21V0qak+u7HzYzt+MDXhlbyKV06ditJMdS4rNLrkpm/hSYrX
XHvsaKjAj70R4x37VuT6dIpJEH5RYxFisCrUKWaI2u0yLwDQS8I1TZm1SogWd5Kz3ALZFtRs70Ih
dldZMaDovzB7KxVvRTMqdJtfN2RDbc/OQNUJPabKUCODBk7Cu1idx05marxAus///4209sBkMP37
23GfusUAmc/n/gAD/a2uaVCOW71ioakmuB9s9ckRnoaGf0A6qYtgRfKWw+zWl9M2XItg4vJh+sGl
g24ITOWvkcsRT9/zKuEI4KlN+J0roA/coCwzMrLsMnoiyYOlyOYjGLm5vpR3KMwUQzfxSiv8tuCa
Gfwpx7xGeOVA0OuHvUhZxILyOTOdQJr8A7mYn+KyOP83KaCWjVOZydqaTd5wrvxB51aPhOjbXf1L
vnE+o4srWzywyhIXQpNaCr4HyZfefld3u5DPtwtfIDtaHYKsqzuURIUyTVaLICbGk4MYkMNuwmpv
q0q5pWuQrUuVO6dyzOoNQYilEEQY0DmqSI/QNvasI19f2Bl6Auc7X/ZCtCV5HS/O9Jnimr/VwUAK
3EKJ1LL3annAL1ZbEAKMNjlbEmqun0WcpHe0U6XUjjhju940kTsCZ9oCQVySlRiZT/eIm6GvqXVf
9rmf7/Q+wU3JlHQPXWnEs781Kk8GLG+algnSA9bGeHZIy6CJtQA7sDGQsppd+KuNt5W06GDU96rV
scH/KxCLh9qvWt2Puu2VjHgUTDktFuyFVIQ2bHYSDbz5PW+t+EXShAc+DmqcbBbqROku7ApBbq12
3mykFO26Q5QTXZkQxr4t5wu/xe6Ov/8YUVoMh+/ulfAnUvMEfh2DQIYm2Yfn/eKolRnbBIz3natm
oypjD/fYMCpi9wpMmleYLxsvGV80JRXkn02nHX3sqUjD7bKshAhtURKgDcwjP3NsWIbcYCEBioWQ
/67//Rc3RXwXZr0pmus2PkFTgNi7dFdSIkQrpo3Vzjg5vv6kWp4M5TuFmVbSHDsA5+H5qrvLj/yi
PO+PLegwkg+Wy/lZ5IEMQzMeFbk8oNuUzwFbN/RxD19zXlCVZtQbMCukkxuzy+jKZYko4DzSHtRE
e7AMbtuzJaPgesKctetpKrWFoWU9d7ySCUZYzOPyR8ukdyzPemi4yR72oOvoOe140zW3UaPA4tEZ
Ug/b4FZL33uDKJveYWUstrhxvM2ylaWrN/i+psESdXQN6aU/h63fF+nuMERjd+2EJm7EeGzuBVnE
kRbUuB7DypRF+OGkli5nshTsf2XpRSYuffUPysbcRUdYkMmE7h2kGACxw2jjj6U50Tw3Yq4ye85i
X8s42RdiavxSw0eNJKdXf0iMgJ3sKZoShQu3v6oP6Sn4KAiZt1dqAy4oHY64YAiu7AuoIWxi0XA2
UQjuygVJueD9Xi7Kz4C+uBwgWFDfq7fB60cwsa016Ouv2Lv3Jb9fFiGhzD7MRF2iyvuZblK2atEK
oTIwV3QdViCneYnj7P91dEbyZuQmXV9W9IYJ/Kn5P04tCwExFbvLYd556k0wl/FNFn4FAdHMHHfp
AtlLVr/izMOhNymdR7OE77VWP5iPOiaovaisZgRRieywUhjMSpHeRzHhQIYBQsEzl6AvRgSEe7BO
gZq8U1tur5gs4lmQenw3vZ/MjRq/qN2vGT0slDz0yV9GAK/GYRGC7dscs7+hkaO/AUrciOJ484Iy
fVi9c8s7Zb39ZNBs3okuxLxy4PXrCZOEhHhriWXtswW7G0QAsv55s2vNHEiEceYcyCYDgltVXe+g
bXh33sxyAgjtX59F7mFLB0mA2FtxvxF00UW+fLJ6xjqgOoRBNb2ai0gk+oxTN8VAjuHa5vh9EMu5
4LmLg3xLaFvDxE3GMvGkYc/vg/hRbmQgKDMy/4UIx+DfBr8tVHfTh2nQaHiYEqQq5E3wgO/dugk5
FLI6LjoOw1I3hfNxB/elUhi3s+IJAAmxoHZfZrfK/PoO14KY0OHlnx6ucprkoqg1Hf8ogRCwx+eJ
RtSxGSldxOzf0qVZGtghVNn2Quv7F2WDSYJeop4EeBiEiSNL2cfWrqNJKnpjxQZ0ifELl8llKod+
rQSFBXShMkRRekZf2tK9UWWQ7voCZvYWF4abQRiBtadikByp9Q0pWQtxNCsP2bgJNhlYdz+qfJwX
i4VhSLbgF+XSeFug12l1feMtiukEeAkD+5GUaWxoxUgvsbtYDHnaMKyNV2f7k7c8L+wf/Fgwz2rn
4cyPO6mORwoLzIkJeaznGzSk0PIOrg+CMFFx6Mt8NEWMuv4RpJvmGA4Io7UQl7rPrsRFzg84nt8G
pAMKkV5BxGdmCSj7DhaB+GKUPff9EWzQUxXIDwyhUrPRfWCj/T6ITlapBDobPeiofKijmPDzy8Xi
pjMq/AX0wOL9sJwtrHI2R3nZAxINHFO3iifp2g30sLayf5tC5sEA7vuyYKFl+RE3dL0Fu/qA71Uz
0/kmEtGkHx+LqhBqwIRzroCo0eFcyoKRJ2LnmpXKPr7yhNfGQ+M+R8rXEMmT11K0sisW50DalsUF
FBzUo3HUi18h+k+3J69tzzQGcMXDYNgIv0W95sk9oMvOaKa2+Dlap1hXwXjxWpXDy6PyhYS6wGn7
uWKNBgr5rzT6Nnm/4nFpY8JfKtUlbXTUEBZXLj+MiziQNcENl7uuu2h+/hTJ7SrmfJ5zVs4Q+tnZ
bf7Zx8OiAqfhLl1T3W7KL0RSSQgVDjNvBnaLsdK+wMvURH3z2q58BYt511SL6j+HnvXtiTI/GIAB
tNu/lDGzCyrG3Yw7hH635s7BledZSP3gJqpshNO43ZhH2akeacHzkwZuXp+GhHljbGHzTo3wam91
uV5hpBDcKxCH+42Wp8G7oUKLUXwyY15cO450EpHG+lxkZUaQ5N7KyLD9XHmnD+L6xqVHHDri1FzJ
mF3lp26x+9tYXRrGuUjJb+qoUeXKAUEWK9nZR+GrvsNdJbivDFow/IaTVPQiH8X6HXEpg5MuwQf2
IEpzyp+Hzv3c8m8QtOCIqQmY+OLMe15R74vNBLKbbCxG11IRHh8aJIMkBI8r1TzBJ/1qi7lJSn+6
7D8o3WVCaCE9Fi6quW2Fk4lxd63CTnjnCnrNk9g9mCzgifvWsrbrK+LSSuKh3yy+8Ea5KjxH8cOm
f0VBBZuqz13i6Mf6LkjzZrfeAoY+iO+ATjPFqqBmia+n+1r73ywVPidVvxwIds3mtR2H0HxuJ9/u
ghwBX64YDz7Ez7NycihHWH2npuV2BZSjU+EpZlzhKb7OTCDtutpbYYk+ffWa8fuvR9x8fpnkepdA
V/paa9vTUh73fGo8yoPFUOGLl6QrSKjDeRyJ68bIhuGYoT+VoBCffGw7CYifr0uMR3wROVheO5yn
+fKibrhpBPVHHivTvk6N3hWb6cwlODaVNrh0LeANh4wJQdZgtS8VRjb1CrVQ8ptw69ZkJEtFRfnL
VY74XfpKVl4RGApbP0t1u7RtxWOQLWnBzvrGp3iJgCrTLcBCS8D8+781IIZvSJNnzicLmbxoKiI4
7V7a5QWG+bWYICfZXDLxgQD4FNMUKbqD2rddlMN+1JYgujQ46Lz0hh1y93hUPsSo73suK9zKYdRl
B+qlgEbG7T94xojm2M/1XPtbyycqw7oTJsSMYEJqFmGw6hjO5SnEkKOnIgx5oVEk+Ikt69L1cM8V
AIMMZ2B23bwBA9u4pzrfGobxy6oz1IJs0ujLXc/l2aIj9NW5UXHLc+Su7157b3MfggXTuf18x9zE
8YH52X6KnhGjQQGWpmMgeL5ZtUbHcGfHm01sa8j4cY+rkXSUYcP79QlBSQP0wgme5wXACNFBVs/7
tPO5sXhC9Rt1xU6+6HNsV068SSq+60oVwfhRrlopurCuhu07iY1QsBCQ+qmoEgG3BfEMdlPRENVQ
9tG/9uTewr922ae1G/FKxfuAgxqAN0wkbjPCUGXsVTRtHQBXBN5VtAyh94Q0hhNiM+X8K4gT4TeG
QIfagC1Zy9NIamZNofoDxkAEg1pehKMmV3t8+aBU5JdKiXlXkeyEGCEAga1XFXbNeNp/V/p0aqAG
arFyPElfkTk0iTSrjbjtunsFEZJYAXo3PZN3i6bg2sZszzEbvN08rkE9ofse/hWlurY6f5V55nam
axjnaVDglLxu0bfJEdiwnBhkY5PNuMWCZjJk25+Kv7ATNasFf92tRe7sSwWs/lQVdDjbzyD5ldMZ
Rlezi2mA9nQlLKGXFz75cLUtJWeLpvjG2GDbUDeIbScpzyf2S5c+a6gVjcOoWlnacn62lOyB5z/V
OMIOtRFvqkqfJj6pju2sI49NizcFj/ysDYjqujvYClLmj8f154KhAxmek7SmpSk/bHzJYhQzJ8G2
057fSYRBu+Ylhm5jD3bntMd3K0jZKom9Nh/E35p4VIri2fQy0PhH+3jOROoaaG5H8WLq2l8CvMBb
lfm4U0HCOMO4BhV9hSBjiQ13MnQVLLQ92NVdPJnHQ1/XIDf+mhiIk7TexKsEjuVwuuPSlwhQoPbY
iMdku0fKih6kVKQlYP8fP6GBfa4ECouv6Oj8Z6JLclo6ZuHnTqX0RvXxuS+hI5TcqL5HXK+ZM0EO
vZKpIfJsRNrNJXqNrnJilaV0olbICvg1ixmrEddOzbGOyjpg18UtGy9mguAZdAObX/n+uXwU38p9
NwVEU2mSyV9guXtmpC72dR7nGMCfaBKzD9mue6BGveZ1MDd1xlIRe1Qbe4aLSC1n8QjTjNd+3ACC
9youvOvdzSHrduxepNPhFK02qi6IkGJYF3BFY90vX2T8DJSuvBDMko9NANRQ0+7wHaAYEDk/4/TT
uqcUxkTesE86KHz3uW09pv98EiV0B549BePgBDmRPO6SSNygJj6AOjRiOkVxTztZzel4a9K4gELC
6RHdGHsGZe9h/c2vvNfoTSr6kMJkIuIOscL5PUF0huJsdkvIJcLIswh8yNVrtOlkRzRhE7Y1LMl8
37j1u42pEYP2IRiM+ohK5v99olv9y3SXJ1hCbd4XMOyqKiHELnHFUzjqSsF4aITwueSCcsjmRFLS
VIs3a7YUspu8C1F/saNGJU5w/0Ixq4YszXlflX7btnoyMqhmSITwjxMru8DeKmKDddn9z0WZdLn2
NxQIyO8iXpHVVAhPn2k9NhQ91FmiKKU5Rri/56xjr0DpMkRR2iEeC92sgIItHHkeqA+eT5YMqVUy
mxMqwfRAuxR8y+Zq21dpiYfDs08KraGbAI9OA45K0l1p/K+KD20bCSiPb9yhOnfbtcLv2oianK3r
3WZmcwr11Ohs7NDIRacC8kL8OoMOIGvK9Ed+Gwze+YAFhe3pBObUXryhlKyw9NnkBYQZjmPnjNZ5
h55lamurmMggSn+25Q2T+bjgEqoS3orp5Q82PUWyVK4D9b8iiLej2w2RA970pypp8sxu9zGNJWAK
XhSHvjvXwFR6N9B9aXN/ZZC8KMsiwt8vfu5f2NMCNtqnm2IMNguZEUU9IoF/z5qQR7zzNiVSHl5C
XWpLvFSZgfOyDmMXCYJL/d4ljLaJmxw26wujbIFYKXWmsNEzVn+95lDDtyP4KURuxo7WqV5Tih1J
WWWJeUjq4HwxEAp/yk10o92D828+lrIZ/BwgxQ49BKGHhz77JU9Ih8BkO6T4K0bL6POeByIiS5Eb
VeJlun7QXu+afHbhjPxWKnDRk0F4SdU6c3ZW11nwjsxdfVJ3XrCFhMggkJiXh4Ck0EBBB5cQvMBv
F6oGIxezr5dJpO+0YfRE4CsU4TgP+3q/0DLiGfWsLuvSWY3dKlLT1+Dk+pM/hO0wxrpZTrViC12P
JWG0m0YZBUTtBsbRGH2QYjmsqBrfi5KfmN3o56/wMYyQ1QLg1t5mTs9MJyjP5bY5RP50lM2jaKDx
snpEP4GHbvXpFXimW2rRZ7kM6R3OocQTjtI4f3U8YgDH+h78jBQFgXzaGIHSMxhT3XXaZV2jfARq
SLlmA7FU00wWbB4wYfPRYNmVWG+7WdHu/qU8GQ2azUje0HUxvf442EJYSutLBvy99lFaT2d2eqYL
Y6n9a3c+T3TnWXxXZsAr9CmMSSBNhGcx3Zo65z0r6f4JVzIR2q5VgOyXpWrNR5X4iHjAukpsrp3t
xxt/PZC7nno86aAgR7qgpN1dB7JTk+2yPkQWA4o5LiQ+QUVqvC032fmoJS1azYnKdGNZ6f11Hn1E
+45csa0SZrzMylMWol570FPqtcpF8TtEsYwHf8rwa+5Z9lXGo/M6We1VjlEdSnrJ+mbr92iQ+dVL
TefWDPBRhusGB4vcu2E9CHu+eq4EqJU81Z+C1S9ShiqyX/+rtCxfAz+050uSn5gKMlRP8kQPtGie
AnaL7WSQynRe6TnywQeDj8sIPo9kXhFLn5yQaGSX86qoT6EsAu4Vh5M7xYrKoVWIyZdG+nd+3m//
LzqMzG/IsX1O42LHJgrMViBsVHnv7VCV8GYSG5PSz0womxO3osNHr80EKcwrbErJ6pKtlMyv4Km4
9a/TBTlmRphjTpwNLGRDjiSec9Pp5EMWKV/5bGth+6IPLYzXq6JlZKeM9gB4DZMLO6VcboAOp/5g
GgOkW6MEqAGqbwaqIzgiLGj+ofB6b6p+ivfToBcbfZhHtlNGlCag3+eKhhQtKDrijg/vViEA6pAE
uLPjl2NPt1wyby1Oz1ormamuUJvCrQHwPDdHp9llFEoHwuoOpzUpcxo/7DfLh1X0sbLozVrmU2IU
8qOYYQRmt9cOXzvJycq+zf3VAD8t01pobK/QgLPAqiiZpNZc2JsK8YXnSsgUbgkE/MjDQKSXnvkn
SqMm/Ni2CukFIFlhZ8xO2R2vRQHeTY072CzLul5M8PhfJNXLnWw4LH8ofMs7Qw+q6+hv8VJKuf0/
wJjNQ8Qu1c1hU/I2lkwtJ5gXGx2lPTbYQMTb6PDhlrUSv0XFvJkVqmSPBqITmcG8TFbOLkVSHSoz
CpK8XTnATtkZJa/0jzCG4RtWdL5+fF4Jl8/Mx6hzz/n0ZZE2QCpDnUGiit4vMEcIFwvU3IosT75C
m+zTkiZyBH6EDUmcXrPsVlvm1NCXRZMMW7h5xzUz0WpprK+WweZVXTpi7EjQvDN0lMDsPlj8tPA5
wACyvlkLeypWS2OrHTywy0auoL+MHayOqAXpCmX0G3a200UESwnQDEZ/Laj7uV9v62ICKDo+8Biv
aeTk5ccc8nhDfVDtnWd68d12zlSOi+WKrLKpblWDxSUFSvZXOjDFxu4gcf9V0IofSo5kEiIqqi+L
Mw9rmWVj6RtkXIcJMVU/ubYVHSZXUtAYIzu1TWtoNR2CmWDFA0cHMDtxOH6wyjhMSj32HaqcDjFJ
YoTypt7pYFosa6dLaYUl+j3H8E8W+iFK7YqPl/rnQ4CGT5reH0t85PR+4jmKa/4LYWm973U8ui3N
J/6OV3MlqqE17+yT2ItbjwlYx9ulpGP3qZhHGAETIsd+nH+4xBKeqQFqWT0GiB0j0TOxIecBFcQW
miBUPYhYm+4GvXHLUDdM/V+A/v0hEo35ewjD9Y6IEfRYdJyhJVgfBp1cp8cbagasm8xlqwq5Ky2a
7DFHlNvrVSRCXKgvU/gGOOMc8zfBnez2I+fiIA/nleZgrW9scn/GahX3eykLg/jmajvxsoDP82nZ
VfyNLOPZfK0cTl2QZIkl47OSoM3FteH73wlBhrhm7ScnpvWoP1pagi0EFYIuGWVxGf6zxOjB9Knj
3eE2thcukOdp8GiDu7f548eZZXzv3nnOo94piwM4suj5Ftn49w4BeN/iir7mTzgne8xxZV300mwN
J+XWUxJfHcozQSuItg37Kht+EpqTciI8RaGds+kLaW7hgeNL6JUZjz01jw9nzhzOS5MjMUE9rDwM
HmoDt/dAXRFGOnfkjzJtBfdrKCRsi+RAHPXDnWLcNBa0cuENsMQ5/3CGDBb140/Fqq4kRSHmIyZe
WcHZHQhBLdNBHb2PgiXl+laIRJWZj9CyYUaxAkllCFLo1Xzuk1mOKiPW07dcdcGLZ1e3z0SP5xP5
NmDuueYxkbqYy6PInoyP30Dh5x6NV513C+JhE3rLz4jlH+WAZU607jjEkJMDStFwmrTdVsj2N8Y9
b2C/yBJY+UgMyIDPGwMptlAzUJOL93Dnq9DZ4ZfHQWUJhfziq1O1JmS5ZAQlDYhCZGI7kq6ps2tw
jj61bJ/VSKXWO6Y1IydCME+NuPVQHkxY5bRWuI8SP4KnpnTRGdby/PmvqCUdyz5mxGTRCsXkjjke
CG6H4U53BjMSniVbdUw2dyjgV/EmgvwZAECFnXf4uxCKv2jlVAeIQAJcd9pkNp66fM/JVyVF76BE
hqY3IH27HffbMRXXZZpa8GnmrSRigBSIbt1+Pzq1zWL0+QS5iUfyGxksv7gv3yfUV0N7C5V7ul+d
uEvFuzeHVhR68VhTyIeqtUyRdJtZplkDibwBJERaYMTjq2nA3/4DKVErhY3XqH18LhO5qF5WIoN0
43pP9HG7qcs75gcfzyHUNndR52offrU+PLcJhy/KBK4z9l5k0ZZZ5tSLYqdMt2eD4dSr7QpjnJ+3
4YuVq3Zdy41UN13iKI3/JQSIYUGUDjsOjM2ICgMZvqkC0ulLRE3IIvBE0XFWSbTNKXPWl4YzEQfF
SeR4Eg/pRaTM95sgCL0Crev9Q1bBCOUwJqtcyUlWAc+0eQD93Yp2P7nVrL9lTKKLktwMpKDP4LCn
aL0iEB6fDOplVFKkzfmU/aurQF2jhna8tAd/EJSHVsHq8gBhGDIoRL+Km0B2WJSziI9J+6hrW/bs
chrM4WNeowOwj2W9mfL09Ws7W6Z7DBKD22R4JobZcuESFdHJMRAy2MBse+35TVpKExygX3wcYz1A
3x7N88PAuyXG8ux+SKs7wQ2K3Im2jYUr0q5chNBPaVP/26NduCMEfAC+YhFhCIKFmN/f1SRooWWm
f16uZKS+HNNl4UD0YlM3Xs6pDFAENm4nyhtmmuhlx/9xV6gH+MTP3HLaOIiurYIhKY97KH/2BqMo
D8O1WWbbcRPyiP/ON9qqFXx+6kX2FCgdjhR2Q3EAdQCGtxFwo439QbXMh8PEAaF88UD48UyGq9LH
5ciwnQa4z+REbmR1oDn5QBg35C2UpCYeSY7AaJe4aIpt12jFiatnYNOLoiuF7xnUfiuu/bwqYFx1
HyLt/ZiX6o7Lax3VCYU5/eK0f9HUmH/joqIiiFsQju6B26qLB8Ig/GSTAE7OSq0M/ABt0MDj05hQ
dlbcdmsGpVD1wTo3TO6E+Pftr6AXR20akhVmgrpfJFgGIkI6aI363+mWLyTyE9tZ9SC46u1Cwl2/
LTJ5BzXFuB3uH7cSFgMN9UHNHwLSHHOjD0XYeq2+6G+hNZ/ry6gge/cuVkmpJHYyH4O/KvuygMZV
xXmBSkgBP2hwjVccuFjOAlPLXkh81Ww4p3exAjMigIj5oLXvmXeuJ62BhwZ6gYiI4W8hQufgamJu
+etagMjzvu4U9RJ/bBQMZEqEKlpLn+zx3HQ9twzWjQsf08iPyJCOO7eCVA9nsQnI5WOVOFVAFyHm
Q/XDz7teNNc1mqIaUA6m4TA3BvjpoRg/dLnl4BEQXsuJfrxTaiAHc1lS3EJMzCbrpiIHiYjXLzB7
idTUJ2IU9Uu4ZmXipa6LEGiT4Z2tJfvxFFe4LENZxAKvbmyHPGX9OIql5JAGcmsSPVn7ylN3214b
rHFwMXyGdLhW7yCzkYIzHaBxzLZ/Lamfv/UhdOZS4Ar2UENusEKMLvE/IKrZJ+M1mFIVse74fi7r
VAi034L+zXP0PUiE1j1oIH+2xv9+Yc+Yu93XKYsqXrQT1WMGYGQ+N+XyQ5PSGjtzDeNyjOrs+qgO
GPmxswuwMLWdVrxQOXBUGEwXeFnJ950bvqqt1RBjjNywC+RxCp6y6RdKwt1VHpMNmhm1udcu5QEP
x+sDOy5w9EtxCchz8gtVxmXW19Mk3KpT25PiQSP+T3bLRWXb14tnWSV9PCsvrxBnNeMyKogWA32m
xW3m+3C1dy9o4GLjSwexFWq/VMv3RCj4iX95SXNU3cizLQz1OagTu6Ajym4riXUSlkocaVfsN+lW
N3SGw+wD2v6++ib4GBbKKScIAsIfkimoNhx5UZt+SL/GzDEkwAjTXPyRgW2L2keAMxGC25F1ISz+
Sr7t2nXIErUPXl4JrR2s2X7BQvOFhHkgzl4TUT35sqA9O773HGnl3DPMU8QR1ulG1snBTA3rMlI1
x2oi2ykWJF/+fxz+qHsOF24A/Hln/B/MCzvbj4fRzM/NUEtG5X2zmpH657/JVH2HD0bPW2QADV9X
lAmIwTUR/U7if0mRyNkOuUSHrixIM0gOiR8H9ikjxJ81WKIcqBWlYA8ZvtRhDsWZYwl+JJyCxU0x
XULwJcS/wuTLT+cMMzosnQk0yEGCk/0vjLPsNRbI4dNvZAlnxnHy56fXecKbcTtwbgzcLWFQ5YDp
knPFGX/N+Y0tbyOU9CFQme/AkQgVPpAb5McVncDiiJGjNlyP79FBBa9Eo0ABOk7WsKpYWUTsXm9Z
WKFg5TIbVfoI42p4ffcPQqJmAjx4/y/JFpDxf1epBFh9sxPcbWlML+HP1e2r9t5GVlLbbdROjXmL
hiTkI1nM8chy4gfACp4+7hpT0fwN4LybLRe/GeZPHRWLVq5VXg1ppqjiW38M8Ed4QX5rr7JqRXcB
yfr2b50rfIskzXCqHfxHU2eddlVJDNU3k8IsoxASNjkrrkikuIruF1k1CHMg6Rblu5U3Vxg7atU7
Zsym4DU6fBMxcefrD2S8P1Rw7BWGFebuSCdPTVwt5dZOo4GUgUjBn8JgVWgPsC2ogNLM0KHiwTbj
TmiJNKtRHG7yaSy+CXhJt4VnOW+99H7K1gVUVgaS4nEcBDS84Z4EsFXvNhXWDhFvUv7cZH4Sqfzo
IjVMtjiDZebz2VBczQmVbkAgIpMHet7EPQpOHIO4q3mpIN4ypNxNQaQXhVwkBGO/Zv7jVgz2gvNA
oZs/F9AWhNUGVFV36wTOyYa8WcSF8VJocYeNJyPf7wWx7LEMZGBptlpeQr4qcbtquvia4ImakRxT
d9OVMG9zZ0cQvzuuUBQFEpUnoiT2kdkrcYnX/oshQXrkCA6Aqr4hLtku0KjHfAARg6wZhs0ASHw0
3rx9IJtCGAtLkMFEY1fkcOLC4OR9UOi3t/c+/U5Sxr2Li3KVXKopOx0qpXi9NI5qriMyl8kdr8tW
Nzuu774BQYvpv4ln2IiBKLdIsPnOHp8JS5Zg7phLaaHZUJrO5nHz+ND29j9utr1ETIpJaXsdczNb
qQ8BBIy3g17AgDUcywwYKrd0lkd9v696Dc47RcWDP4qG/24AichHEOcSWMDrxAxSnzOxrfkxCPP9
Ao2i+EAZ5UPt+Se1bCQyo6kTRT2ry9v5UOj6qKrrF68k/T9S6Sw+5tLsbih/8XwsqDm1mgVtGGrO
eiAchkiDhqlYzK6TPmWOwz1eWvy23fxYm0JpC/Kp4VQabfdXlhXVdH68ffIaEPUfzYVgyCxssGcq
dWbjNHVKnfDRxu1V1U23/imGBwEBR21Kj1Kw0eIkQWo9SNTkfQXwj66qYrc9rpV+E0N6AlhvJj73
KOliXzpJBN1VDLfKAvGXHe9SqXPH3CxIDI77Xx1j4fwm2B2+4EnloBgNYLDXa060HZ9alSjSMD9H
mLvNpHLoxtgZ1nbFbCRiWcPs0Cc1bqQGIBbdoJd87hVIpoPaNGQf3AJxuMd654f7S1r3bKPQ4kyn
PnQTfpsO0OoFoQU+beRJM7GzZ1oePkZpOceLA7ekpEDM0LfdqUWNDQpSkShQjl9xojKttKnQOdkT
DTAoKeaHFHSVnfmUsdi6dR7WJ9iTWz0cogIejh45o2Wi+hM2gvPLMJqOOkZ4z2fEd6d0Qto9oBzN
7NYo1CYmqwuPc6CwaQZ5p91untl0SNAn4zjaqM8zxMvnKJPrsPMy8EoeXjKLzsRdfD+8xuJMlz3Y
/OW4pC84AS0c/dLIKT1F9vmFVX5fTsMnPcO6GbpyX7sOal7o7doDzUjwke16EQ6ouhR6MDGD3qvb
V87//XqBJFcMsvCrLzcfsB0mqvdDw+iOPp2nbj3b3EwlQAOz2oCzl5tc4tjuIXcBR+LoMlhnHV2G
ipg9HuxxyGS0EGmrLc2fopqqLK0+ITXTUbH6VUy8v/lmEIsPo+Z255NhCzf/hAGLd7pzOI/v7mPj
yyDGUUiKcziBEUhh26XNSZDU3FIt2pd+EWlO+xu7x/T9IepoJ9fwGSRL7ErD3lTdrUn/4r1hJHNL
AqkP3LIu+UxQMg9GrTMz6mBnwpkouqE39bKUdOch4nCRVPyn2OlLUg0vcD3vrLMNRYOFTGuniC/2
Qpm+mU4AyuPqf5CqqEn/6vRbJTMbnywqCxdriLyXsfDUXNkZP1PZNXZifANKxZoOwzryfyOcs8XP
f0jC1XMeIcuZCb/6nAMOG7HiSQMwBLGcAxQYDXBnmdEgzVtRJ9hCz0iKb1D2UOnKoS1V3p2LsvAJ
haOGvxwsP7lhqL7D7ugb/qkCfTOlKY+CxtqOCSvJXyVt2xKgpSxMCRhiTYddEV/1hIIs1DkjHNER
QLWYizSPIUEhpqvoACPeQk0b4v0qJvU2hc8y/1dL19RbDkDZOwYu42BuicmYTnZCsbsFUhxZ+2Qu
vs00/DQyvGfhNwmDxbgiInLx8reZMabgziSMKkohj5F5V2tTrvwfn0gp3Rexe/tSy/0Id6G4ZuJe
aV0+x0SpiObG2qaFFO/0kdcTxHwrRg0gN59Jy4b5uwLvVYPsHymrnUseEDatwjpb1rV2cgDd9HZ6
1tdKXKj+YNoFpk1PckcV1JUDUkbYoRX1fTffKtljEdPo89VYFnaaOU4rDNriFysATxk9l/SdXHPC
6TDoNlC1KaXAeWU4l4fSJ/IWMJnU9SkQI3bMuVpmusBn43aQKnf+ecyun7KtQmMQQWeGOd2my+LU
UOgf8Jk3SWpDdJ9WDGxJGoMIQRramMTbFbDFsXyYhyejTrEHbrJy1otPqCZPMCyOOMYe7PeOyl1v
WIZqSqYkb5CaY4uIjgevaT3FnIfzHsLGFB6ae32MJ/NGc4D9hcT5uVVjldQB95170YhMsrD/hEed
8O4f0BHhIheHdjwO/CwbNLrSprlP88CjKZI76ltLUtHRSvh0Cg0hWfqUFh21e/9a7KmwXKuJgrZG
TJ/Ktr/iIq70uI1DGtY1DPFpG91KJ90j4XA08x+t34MbDFK/tPb4fT9LM2UociKWhL9vRCJy6vSf
+/p+UpxzM+dOYetpDDQiR5ynr6QRwRMM/YGBmzUBup3OUFanL1e69837jiqeTsjVRqPrkBXOqSkU
wWOK1LSpTC3a+G8917yyVTyMvMENRdipWScQHLASTXDQS/gcba8jbTJnF34Foiu4CwtFUHTeFxL3
qFfyYnVQywu1QU66dL4qdufMSFVcw6JSEaOwBvmERVkWHkH4TtaaNgbaHOZtzkyqGouXkO/BdblN
t49ZElAlIBYEGz0Ln1pbcRCQCM9q2+xDfGxKgbFW12JGAmHsqmGdrMiq3kmxfmulLpBtnnEquqcX
zWEI3AATO+7F0g5QsuEHfBlrTOZGugSEwyEQ+qQN0Gc8AN+439o4VJC06vGKmoj9PMW0Ly3k1+ka
k2ZGvZX95XFG6X6BuIGC9eZpPLIlwdO3gkYkTSdRNW0b8UWnNfcYIqCd9ZoF7WUAmjvgtTLb1UKy
J2/sb4Si4z2Arg+7bWCNEMsgLp25fKsyb+ZPzgdWIR4TLOCxY3IscK9ocFHbxHx2b2LUL2niAsMt
kK21048aFCSGSsQjpPJg71BSBO9pWWRoyZEr6TQeiChURpTm+aPDdQ5zp5YO5cFskL0Nh5eebC9x
0eq8phs010RqGcqW/9g5ezal+ipBvFgn5E+tJ5q6t2QINSBZCMMkVidyWVrS484qgwmZEBlFZqsg
IZo+fxkXTy+EhMk7mOp/9pREDhd58+Cl1tPhvPZTU5i4rGffHvuYxcp3wllcWbc4iTqvTIlUzhAn
TnvaKfehBTHX3J3XFUVRyBLh5/odLHQ1cah7EPWoRVD/MHKyNVxVR3E8DdslMIytcuuH/ud7KzZ9
G8YAf0Wpt5HddWt911qPGO8ZZgGFydIlI7HZRZ3zEMHakdESth2KefdIYQR/+Z2bIGuGSz9FOpxO
kre9wwcN47ieC3ukdqv9A2ZHN0ch+AsJ5D7Vd1YnZcavkqoEPcwiMMEOKeNl6qgUTtLHOLQ6HVeM
S6nfWWzp2FW16KU3JyCzF/5lgDqGb7b2MKRL6zLMXUcl+MUI+easiNxdMEWRVEXedX8p+rcjuszw
YG8GqRYJYCLbdu7+tp+3n2MbmgezWV1V8loJ70IanqHL4w/uvcwM8dp3ZQSqqDSVwxKYIL0E9H0o
6mxcrXAcKOgl7zfqzH6x1jdxRzckhB8QzvSA19Mp6UojW5wJcdPRzwgi/FeW/QJsFK8XluxqUlZb
4uhcjJKEQDqbUbhtiD5fT0s+5Aj7032Hr9k/sRGbxoD001dImIPeeqCooOZAB93MaWD6QhFe9cdv
3BHr7DK+AVElH2b90809O46STL/++1vSctShfoMi73Ei/werYdSaQHcRPl7DYvU7U7AkKJIRhX6s
/In7PJWb5eU93mCSNSXuWdJgOMy+fGah8PKv5mWlqYnv4ue2m6jjJsPpZI1uFWsqWStqM0XSb+1P
6geR3OAah8LyQbx3EGgwr54CUm27LC47OGtrrS8ZWnMMYm7DLaC8hoN0ns+k+ScFgWLcq05fYAFx
rUhbi9PDx8wh2JTtn2iQJFTDHQCrVENYyd3YPsS0yMI8Zfl6FvD3424YqaH0CQH3oX55V4F6/rOj
KksFoqgKNoo9wr29FEuyKbtoerEEpqEMsBjWOUdSuYsoF4b0msEzMvC7LD2+6+Ee/MAF0WcjOQRd
bqbCQf4YzaAjQhxR8MlAKYozxMRcw3k7Y269i1kUwYSVg0gi3+d/Kx9qYTgUcZMIMl+Is/0RwD1E
20SVp3C3BZioC9qNF05On+vxCmaSc6rCeePRqANhUcXOaL9V7VcJhFI/vW8G1XWcA7iin3GLDF0w
EllOgD5loUsAbLsWpSfmBSVQzyFgSRWZmKGjRVUBZRcOkGzZr6Dg9+NTbeIJQLPRW4MHY8q1MEdL
qa0hglheFLAiV4kckt+o9W+empAES8CL/yAMKnKZatb04xRec4wldGcVFHrUS7s2LoVNkkR7PRmH
oa5jOqZmIYIk8Xhe/oJOrpjq0Ts9XYbeNEWfV7zjoBdWFRktRuP+0qgmLxMT8CA7CUUY5XvMxHPh
CAaZOForbAtmQl2RAFfl4bQkJ3mqnL6ibQ+RRAqzOuFcE7y8wkEP//2+VZTVaeHhtTJWBBILfbtf
aPZ0C3KZMv9fr8nIAXou/55/ksNQXJbLbxeXGnVEW50/9fdjZpVGOAoitrzIrpnhw0o1Cs4VPCDl
kkUEzUasGN1uCjCStgY2esGBn3xG9VeU3nCNxCgeux+nWj6gL4cjupjFMC3g7rECWNNf8BA+fyvU
91TjWrQ69wLR17FTGjIEsbaUMQIJKYVNp5B31P+71sKvjLeDq1NYlmdYkgIILJfSJYhJUcOwYaau
kH2IE4zFpTw2ceRkMolCd2F8qgePy2vtqVpxiXAgLNWZ+Jn42cDR96sS6Arl5VILDL3c1KJkGZVx
qW4/tnLuvC00H6odpQxtmOQtCGuyt+E5hXAJ4LRtU6DNCiUdWKblGyS0uszR+FjbJLTbcLEzD8KV
xlk3oAoEF6C/H5YtqO2JpdyCB8HDtOu+fcsYF9eQdytGdVbnGjhTyowewVQmBPx2m/vXVcKBiOnj
WtNI5RyYfDrVGTNqkG4/CTyS7dew9zkSoxX0Kh3zhS7QVlCZJ2FW2ydCwHOWTLowP3BNsN0pxrlI
/BG/r1HAUOV4h8N15s2vmeFcfVU7cqU3o40UeQ8cZYGj65YyDUYgtuZhBJxu3Tqlglm2WIOFURCp
GfggowtScu59vCUJXCzaDRyg+OtQBGH6mibw++B1TvGyF8zsVDUXWGvBO88Cn36dTIf2VaGzF+qc
IgvlZWFqEIZksL2FVz3JHoLrcXU7RTXU8QhMYbbyHUdIsaeYgmg7od+Hm8ZdlkTJjW1RQqQKhNA4
xVtIfyCeScS5M08nO020AQKgc4f1uIKcMUw0+LeX3DIheIXFLb6WnTg8WRyOKyxWHwUy5fk8AxSx
q9wFysxpGSPetceONXoBmmLFhN+CaRFQeuMj2ZyUsAV/fTpqL61o8vc6vuaPxEuGpvaXH8VAvXKv
PgYIUNUJwKLoXgVBYhyiYII0/4tf2zsDICXma2RlYTP2yUGyZN2rmIOO1vY6SnKLL+2/AmnG7a2m
BNYG3kkM3kPZi2kdj2V+AmKv3Lsda/bhHi7eChU0y96t0IczCAIxCoO7Bp8QDGBU+xqxU2H8OkJ0
+9RW9ck9v1Iub61qaJZVO5OyYKO3KIANmNimmdLWaFmUMh+PgkXKi5pKJWgUMCUdDCrpV6a/7nPN
jzvaRX3H7hrW+JwRf4bJp+y+QX+r2HKEOtYig9yJRdMSLudhtSM7QU8veKPBXS3vq7lpw95nCelb
5P3eQ05PWcjXlRyVqSKGpKV4k01K+pBvdgzIguUWT3IJM6yu/zi+QymY5bq5s8J+9nRCGmCxnuYN
jTXMPHhlUk2/wHawtjpRPVeXsQEVdOVL2YiAiXRdlJvJZDbvxdUbo2o15VHnhy0P+UktF7FSaRIL
MH/2XRAbJK182wf+IwDTtHkz8eci+OLEtfeVUroRTdWCpXibZmxSVkF27/SiDyMz/H7V5aGY3IFV
0TYc0dGA/+E8i0xcdFceTH7UBeQ8rUd/2quBa5HIYqz717CQtC3wyaPZflul19a5YNYldS25EBY7
ZSnskXPJQeOXiEOHY58/88imkhdDNz+0SHvmu6S9B8jGgijK5lor07V29m2ppkqVDaWmPEH+H8jE
ZuPDo3wFmKEeaQcuTt5BJ6rxkFVcrL+rjbVn4s2ukWiJiD1BAfCtBJZmL9EZjbv0C2vUu5+kZxlE
mrMN9gC7p7EFBtBfEr24Gl1QgsZCBWOK/TbQz90sI5PCtFGrxE4ClXrzn+ybbgVZHvVfjfKPImpB
HS/ldUqUIF3If3iV+DuihjXvMNGQpajS4gNGhGOSLC1/avns8a18pxieFOtOirb8Vx1DKvrmdngc
u7WfUaNHiir7ahqTJbdpWXd1cVr/lAz+gScr/VgQh4cn4YyElmzjcohMOZv48KWeMVDz7sEj0U07
I0YMEFy5pA42KJAKYSxQS1Hq7p8A0d7M6kcqCkf+nZ9UalHwQnthj11Fl/W60hlSaOBJaq/vuK81
O5TfkghuB+uq2xkNvjRhEw8uuoa862dAkJMCCG/RigWjT4KYfRzaoWR2pybR8J4At2JZwmHqxaRp
n+4MPVLah6f03o+7K0paaEs+I1ChZVjAOArDudnQTpaBC7pRym8mKRNEZ2Exg1vMmMRKLCcDBQ4n
L0vSvbYQoK19JMIGS5SRfnS/kXDN9kGFTv8ZnMclgrYGFF6s5axKP+qgyqFQi9nVSxCtSesPvXx3
Z4STvIRpJ1GbH4/VAHLf99tBRHzqXOKnIJLEePlTqrr96xWPDLdcxYRWgoq4Eg7+AjhaTxTsLQgg
La0mRtNU1Z2ZiK3DV4W7mkRyk3SqcMV14a9PW2xIN5h6YGJUYf4MoxXY1uwGk8tsCMLDAdzPHiqy
QypAWqqjGDi9u+ULT508M9uVTkb3fNRZz2AtP5JNczQpd14ZtIq1DOqOpDi3rH4jLAZWpvftfYRw
WoSi3vhkj4xZ2MaPpy8nZ1Z1BkQmXjsWMro5GiAJNkrpkNGsy1Ce8RCmAQgeKaolAAaZMV/d755P
jjcu5GnG17JDNeIGy9nb3jymTIviORk/VlDAei7ZO/3JCl925pLNxxGovMGfcXocYLUej+3BZM0i
hQONlNAYpv2PBO9MMuHttHaaBId49GDHXzwN+e9by+5/QnduYHA5v5ePTXkek+wZll92EQ9Fuhi1
o6ZiQyRuyDZgtd5CmSY1FpGMtI88ommk0vfTxnGYtSjbu2SroMaHjRdGSqQEejBrJbTuSdr0Kpf3
YX2/YvsjHAThduhlz+qhDNW0AUaQm7qoRXwZYL6tkzObnUllCJt0U6jRVdNh2bvnSbo2ntFwzhEJ
R0s4qwUrnp9L1wA7USj8dGVaNGR3pRylI32mS1RaLe0dyCukhuhro0e6bZLiTQ+e6B/YBsXxIC9L
ZQ7QVIfGK03y2os1sbacHuCSntSmRSpU3rp9Vek81bsc2ahM2hKGhwdQK5kitrmlp2iWzF9uU9rR
QOfH4KccA9aGo8ENu2mX7PW3hf7EMPgpttljlUmjPPN+Ym0PjEpUD3DWuWFhKWnAAVdEuYsGzF0x
e6KZPLjoKdYiXswYLh0eo4VA3kOYnVJdtoaRwYyl3mn4T9msIV+YAbUXqDCRljaoWNULZ386oVQM
AHfWkkJ1xK3XHcU9urZwesXW0KZFh3kA0bIXUBXGh9gjPQ69e29KXE0fk1kruTdzhKQfQMEVEHkS
hsC8OOXNFKR7JnkUWSJIw8EwwM8PJdZYqURZnigWSUX23hDcgQSY5bvSRTH9I7SMJ19mdAY2y+Iw
3Uhhdpx7dMCwhuQFe/qS0r9rDJzVE6y5eqf762D6d0/iFVNE/57aQIe97B1I++ujiyoy91z/sx3h
oJkJ98crbkHir4YJ08gLDcpzY9XbmcC4r1tIZ/aU5fdkDDiqIWpefUdTMZ8fiktvQQIylPdY0vcP
m52ij0IsfXvLP62bmdtNMMO+pi59mxJ8ZR2L+KT54UE5wMkN6a/LtG+OVhx5/ttoa40tirGTGM2M
RNNdzxthlrJokWMBgZbKhvCpAkqBmKWpvDNVNQwuVvuvvmRBPRRXCIUywrJR2mrxrKE+ikii2iME
Tnl/BTimjmrMB0A4CJxZWHxpw2wrsD++43Gxa1hx++vJ5Nex8mCVotfG6uoXNMk5TaQL/60Kw7e7
roefw+w3YXKQVEYKHVxAj7a3OXMAzbUpl7FQ5XwVqsNlQ90YDq7d5CaIVFZ6HFDYshG0j85XVUkk
rVINLFwWIQDtx0EnnUqQ6yrHCGN5GjXw/RRel6kmxaW1mnEmG6Llld4S8/eTmsvNB66iRJ/XW2oa
ck+T329UzABnruDsGfV/dzmE/uN1Uo9dhHAVAk8rr/x5HtkWcpyI1O0LDzZpSnNDF4Laub19Toft
AbZgB+S0hTw9Y3k19CTHVdYTAG/xJcLlJCBNXDcpvaPLX4wOID4el3ij/xg8wnZ4vh5u8ylBGoYQ
PdJHEy+zm0T1IjzZXMOMa4zdcA+Qo+zwtudKLcYxsJGgL6htcKIn0QubS6/1zJYd5dwS5XQXY4NT
32JB+Dao6TqBt8n/CxQNoLDcIsKZ4AljPK53eUhFr2T5OsGa3grCVI7rFK/D++6tdhZQ5LWpeIhO
eMd9c52ZAtTciqpV5gKVPh2QqBlmaH9BB+pBCTuSb/mOTv4Ut3lDNGQyFgew1locdAxDCXQQRfiA
BZZgj6gV1HKAox1lQQTSRqv26UekYUHkTgJqs1mlOvzj8yGBxzV5mibryETltwriQ47ZQx0buO3o
cj65oEXq++yB/oFIfOE2tvXbpPxkYb/X4ikWrsPgdsaupOxLQSrUSYfcEbnUfik3M5hIypqJI7Iw
d0lpsCf4gYB7hopENX6RX0+yhIaAveEWvYwWRAVPK3cQYLsGEqg1JRbPADEi7yXN7BsNIWF8nDZV
zdjt5lqcZfXjKkXLCaryOU11A6Mk07StlW8a696Ez7hKuWfOqKC7jcAYFnbwKLi82m47mlUTQmVU
e9INEQ5qcyTHetONDD8ljaQZxE1aHJFcdPWdBqDcoNNYNrWL20Dsd/XNErc8sjxn5Mp4DB9SxI8C
sFDjQrdNTw9cREqAQRHhcDNhqz9gP8P/PFQPFLpB2lrbVyoKAS0+wRdgAFDdgrRWg3aysy7V80fQ
zUpitRVV4xbucIxC2uWLQiEqRoSgaKcwFcdGIXFCSv8bASNGkchAs3+WLmpdZjUMfKiBtYBPp60I
HgQm0ynMC/L7Ty0q534L5tW2ZJaNL8VGLQ310HKPkZRvbP5oHOSu/ZE6OdC3WbxI60Fb91dhqm8X
RrfMtxXCI3UTphWkpn957iJcBTZHsbtFT7P+uwXKu195EAWnojLXqIOywIku0hPE1ty3XGw3jE2R
uJ0GJAAe4B4qKyABcZyU5PWvmt6DaZ8dLk9hmue8XdvAMjWPlSSnQ6PPwJM4Pv6GT3Fip5iUh6pv
ANf03sPngGE4TJfKptjFo2nSdf+zC1p+20ATTa+zVWdFg2FApmIegrF0qqztJu9IeCQG+pz+y9vA
YKUPvKBV3qtGNv7aeCIbDBBlFizSg/LQ24bfq0nz1Z5zoooRVP24Myf/UEdqqibEkugQwbytKn6y
jFkt/o78hm92xNxw9ldT2ZcqDLNUuc++hFqn6i0OSSlZzD/kBAxHthnETBOzK/xMFR9CbN4SanOw
z4YZ5kIY0yoV6G+zqHMKQ79vQX1PCKBYDnuvpFis7FC7UcyIFApq0RDXKdCgp21R4tVJBhK5faOJ
6l2OJ+afjgSjeUbblLo71dKd2GKi/a8tXCMtJESBxYy+ru7mzHO+YakbPLZz4jQS+KmR5LuK1HPN
LtB0IoUWPQ2iDxetAGCMTAuD2RdlRlUtCUk5pXSmHVn2cTGrneWEQrIgwyLANGShqcAtiH+17cUs
SXdWWJEVFaoECxizRg0flCOEKYHenhmQjFbJxk3/Up+xt4aaYyMGCWHVE2btnBpZxGkOxW6w/1TS
nJCmjA/i8puoTy+O8VVGQlLBbfLD0M3hU0UlDEzhb9Hs8+2sd1TU2qZ4jhABQJJbngEveFsd4nZM
mD3pvtLv+WgkylWO5FC7as743xGwIwTIaGD3UpERmKtkdOxxE/WBs+46SaTTICf4/VmQG1WUZ4ML
zBRs+wATZ7GaoCBDJuUhiBsKx0jTrSIuGm3R7VSMm4iNnWWvcaIgppWSO5JvLbtsnQASSkSs+ELn
KYcdKVlTd8bBJ4xenAiGBi8bx27b8+m2WSECkhOYl9hBOEHxqhP7d9+4RPBPYSS0fh1cFzqMgV2l
dmtiQlkgKmruzGtW6tGRT42PohfN6tp/0QYmRF+qrwgacH8sgTvGgyLyAIVHxCws5UCBCL7zwwY8
iYHl7308EEYCt7Rfbv0j7JU+S8HJMm1szA3wtc2iWdzE+s5vd7RawasFk1jmFy7s2vB4zLX3ftmd
NWOLzmHQHveQ2pg4Tn/Od9Wc5C1I9dYBBoBJFfrHfsoHS4O2O1fq1rEHzM3gbe+eH+Tu34ljHhiI
ZOdpWiwtzje7ylyjPhOmouNrXBQq3d85eSg8OToPMG3D8OvV8onZP/R6QlUdPNkDwJFv5+MYIPrX
N7Ud673LEK8bTH0kjhYWDNm63dPr6v8DxqR8cerGrl+44JFTxUCe+9yQZCU5MmQR49LA5Fu+/ec8
tgQMSKlYtSPtVpEzU76olRmKx1SZixxi2f9r/8p2rKjSf9lY7Z2q0g7aJetAUlkra/rACWFkhepw
cl8WE50yddjMw0pVFHSQSuTXhqH81qGz/iwu6xWS9xPZh7GJvetz/MS29LS0w23ia840YIp3TD+f
kwl3G0pj34ANpdr78Hpo8uzr0RQJVzQ3KNxONotNUQbdGDYW7io523OZWata1AbLi+tcYG3eeOA9
AnZ+Vh9r+Z6+g14UGtADLXKh3/kJEyAMmR6/GVgEMMqR5YZ9JwTK/ia66iZDNxhayicOjBffmZBI
OOUN0Wm5ry9C1QeGeCgRNkAS9eQ7Ben9IYH99Icu5sqDWOoXOYzk+x1FTm/VQvdiujJWpi20p3Fz
SD7R09V8gU9G2SqNfxqVY5rH7AARd4gtqsAdZXUBsxWAJZED4my2qEf4ISSUQtMne4hlfkFLlCgi
BzY8DHZhhi2RWoAkEwmkuWDuBfiMF/Y4sNvYjqNbfX4+hfWTVOWTStomngnpTlw9TZiMPlucMYU2
QSTOBtckw4g54VS3/h8wf/bj1AvoBK+rZ6qKypIzCA8VcMVhFa+fvsAe2N+to2AwhjwA+jFJLhnc
3KHoNFodZkU/KB+kPzE9v5LRwJaRbmOWsxazBgv+F/jeXnf8khkyZnwceYUO4Tn6GAQsmtEaytiv
/UYSGcmdD5f3E0B9xAuEybcWgM/UOdUhOHu4aESMCg0zv/COr66t1bhwcZcU+ASHVYd7HI2JYkvw
/r1KCNyquW8FbTz326UoEsXU313Wt1FKEnkr4qD5impHFUGUt7ShiSo+6lgH8Uxa0fC14aKDA0nt
zj4gMibrF24b7X6OTilFE+juatopwa32JreUR2628OmxiHEKyxNVEyPHGF2oF1xfatwq0SZqWZma
U8R9+Xo6FXiA5EpZQYJFat1W5uTKsQbbMAqw3Pl+Sfo7cgrR6U1B726TB9erXD2v3wT2wBJURY4N
eSZ04or9WOPmIVFphtvNRfXITzBy57LrkfkLimwM6qVT5jsT1gIYBMk1dJfhC4NFLaqmSFGqQ43m
9hdzaFgPyHQ5M/rfwLdFJFzF0LnBZd9XvHNThi+pqhdRqnL7+t3uJN9XDqsAUqyGLiV47MXdPzSm
BxVtivxSAimC6rrzg/NkD5Xaxqg6bFiWmuZ0iJQteNEyW8iznSnyTHrEmYjCcQ8TXNFXpM78lqVu
oEnqcoPAPboRbf4nMH7eZxNy8O4K5Gs/2vZqvxVc7hiI9nR/eTlAyML390GG42834g3BhReZMAwh
LWGq1XN+9VHNMi9rl2cKdIhcPPKCOVaTJkX1FUmCTc0VrUeu0wnHPEHp6Bve4K3orbAawGIICrXY
Fq1lij6xFg9c7oAbYOoN7rBcm/FC5P0mT/luFxhczSPr0dawC6SNgefC6S408UkDL2JtfDAh2jgT
bAWj0+woEtAwy+QRoSQ6n9oZks/RP3fJbbJqqlxUqSqshTpm4LipyTEbI8HLkk6vwFN5Us+jxAU6
QfSKOuxd6zBWphqGxMfDaCq7AlPy+eCrF/oSqz3yOvZ0xjX9lh1zD4gMz3/6L8uj6EjM3JRzBBWF
X1LZ0kB9VSMuTuIAuB1imfa4uRF53ScYsV6kQG1g3GJT5SBE/QOHbKRGV9CyIHjyOaYTTUAr6c+a
UCiZsgsQeEZNTcPZW3GBJIZDk7NmCANALWa7HfkCdA30TeN3sS2KptVmXc9LPcJbhCMSExE8CWuE
pagOr3hXubXJRwFapa7Re4WTck5noRcNJWmlAGASvU2N98JduJMGxTf+MttsDEjnZjAM8hcz2/d9
K42Q3WvYEOXaQEjdm/cTVMaZ9AdfijYKzZ1Wmj6Q3Xw6OoZeV5NAUR3xgYIp3EusNsz1Dfs/Us1E
gNrA5z/2gA5SOBZ2/FxVPxWtAobsiwyBl999Lnl2ZNFAPJulRpLMI4+3IRqyxR23BFkfNxN0nqk+
GymFEmo3usZ1gljwrUtcyQf+1rvL5QCF/fD75vyRn6CDYFdjgyRzxBuF8pLGcjh/4cfnuVC1J/mr
2TQf/PQ79cpTSN4y9CTyDukSOhm1pBu0TPeTpy06e5fbGZCqqXLkj543/IHyxgSIFjA0qXYYw+7I
xv07S9xY1aGaUSdrLzbSa1ctqVwTJtJ2emU3sXCPNmBU+3Zp9eQVQX3IZv9ofWxr0LVNBnJ3hAQG
hq+3lDfDEvyF+qRyKx6JpmV6JoDWfSm0HRfQKJjBsXk7d834rsZP5CeRWSDS3RVxCojpsErYu2ft
VcFZ4J8fybGy++rislSQWG/tmeL3N+ad1W0PdikOOsWaSnkashptQT8mf2ozTz1cVdzH0OoIzPZg
j5GNY4TZ+7Mp9WDVmK6wCcAVfvw1OudSXElKtIyrEv1GuKAVFWckPuphznmgmEXMxP7wZZcoKtWB
FUbQEGoqpYPVhkFfKQ4pkHTW8MmwvczeVMOsdTiTbVUKKpho41ZkWrT2URcOQYdVmUWUUjEYnkZ+
ttcs6r6ptnt6TR6BlgiZFxV8C7pViPvJ0A+cTVjmZP+H5geo8Yas46VzaTQKSlg959ggugxuKvmO
xeO7tYgzxgX+sWUOlaRfhLObyh6l9DcyEQYHEjI0Fe0v9U8JkuoKyEQY5Pp4Es/10z0lIDEyiofm
VanP0NT+ij0QTeR/IRS/M/0e9afs+Rfaj2u6osMhiTKE9azHKYGmDmFzu1vWAzdCy5G945aXDL5j
DDv44LASKgXAqQjPszx83wlBg3k9hjpNcfPJB0AoXIspG017sb1ajYc48JQl3f859KwY9GJzZFci
ekdyZxV2vBW7/aWKTdjEhCwGkpqCwD/HIxJM8bcndr8E0I1pBekqKxA2XewPPaCL0m+lUYrdjYtd
vsbiS5SiDG2PJAggPInuhSLsG1XCpsrrX5QVuxngJVAZqgR/ciWcSn/gpW9OVikIfZGyQu6Q4wh6
PM9VUGidMjP8VwxMXACtfCAjnW6mErmAlfQno+x99JZquNaFOhqYY1pE2gjrSJmN5P0jNHmgZNz+
a1dxqIE+IVKQ5DmTvKvCZ4AmJaOD+6tc5nJDwZFZBvEiMEqXtK+AxY/z5JCKnnznlarVgNbiu0uG
QJWKm2tVbpuKkRnV6ny461f+tJkQlUNcu+3Oak3KzI20Fb/FnNY7iVoJlk1z2qW9fZYvgGiK2xXg
Gqf3rLxplUrr6HkbxoZMs3vdWx3+ZX80pya0Ui6pTkGBWtlz2czI7ZXRcc5YfgFHhzuhhrhbECjD
/qu1cksY70sEmODgyrMN1Xh4NOM0VxHZCMOIUyppYLuFpYCvlKBcK+ppFvdPZGAFI12uXCexMJd5
azlqT3yEpEOXntSysCnc2NuIdwvi14JHsUw9l+Oy/5jcr9nTV2Y0oiScWIXlv06aBNulItvgVFCd
6FlUZg0NTIRjMRIzeG1E5Jz25HjyPCGv8zAz6yTBBHu27mg5f18mZ5fLZcYts0PUjN1opT95NnaI
SBdQEQWAKQcAoXXgUZLYgUqdn4MkoshnsWPWUDd4XrpCoZ+LUdfNi00YFxInTSc0n/D9TlthCLoX
VA6X0Y9O91T/S4PvLvH47DMXSt8iSPm826FEZBhKIz1XPGdONb2dmzY4hzOGZDJGZ3RsRrfoK+Gb
5wQJC40R5HLGXO0q9uU3gbJ+zFQWXyakOEhpxMbIEi8LS3cKnCwaZlaUR5s2t4MTv6MQIfCAVpmi
olcw/6gvYWZ6MXaTYvYfrWXVVlJveyH3mDp1NQKqwXqxg2NUrfCpwJwQn2iSHtvA2Zz5VbFzPVI4
+i+R9AWx4GjR/ai5y7WRQ6Ql1p+DJHqDX/03J11zqKdv/flNmA27GhTakJEL7gdAI9xG5n7pZP5o
ZPXNl4g2iFt9ruhLL1sBk4cCyQGFXD/NDGY9zWA6N9gleLRFTCyu1+isj0E5CkLOQFpdVQDyMLgG
SR/9VNIsyF6Y+EjrxoqY4iTEGeEuur0MaqyH5fZUvwySfu3klYrnFEDeCulaeg9FQiXxUZyfU1Xj
UWi6TTmbKlXdkGBUlnAB5Petgt6aoq4Qa6SG+vwAMkmexO/JXJfuY+LrN2qEYxyqelv19+hVobcE
eT6xrvYOyYOt8MSCk73c+aSgzL/ZkI+Dsv1EK8MzEMH7J/3/OJC6NkIhxVlo3UoSUFJJu5O37cq+
UzGblL3O5buNKHbzElbJc/YCt5oi4y7TjP7c00kAJxo0zQT3apY2lmA7dYvmIRPKSOhhyuvRXOKJ
WJxI5ALoWpyFjypP7cb7kj0GuUXlXdQszg7ORs4hQtDsL0GzxkSWdlPQV4tAflN45IRm9KDvGwuV
oPmxTgzCIYntyLe7XV7MlJNggxoTk2lDsU+Xfpv1SPoBx9dfinljKfRXPGzBBWev0AerhXy9pVKS
9MJsOTIxvtSiE6nSgM79kzx21aKVDh5p6ZfcZVnzGRy6bEHOI+sfMjUK6qsY/hny2qLO+RsKElpf
yftpA/+GOiODd3d8DK9MWcSqGb2ay8jivPOUj9kvuMAcAfFmy8xGcxO3uPrPr2K1hDmRfOFTHymH
7ubNaLJkHz/z7y5zFMZmV5dXeCQ/PrcZhitjU9KnA2KXhDS5K1nSvgSz9nphue5i/42fyIMoKlC3
GoejmyjeLg7Ncc6No4v4AlD5NcR/x/T7mYBE3ohCpSRzDCRavCzMk+gdYINJyp8lKb09A3oKW3Kj
dVN3mkQYCf39FmUa1M/23GaoaePa2ItjQWSyjSgD+Qky3uzXenMgpHeeR9QUoDdycduzKnmD5lbE
Oqco12d8O0STQvQpl4Z4Pb4s8CoysFzKkmytHesy8A8nDLPtuezbu+gewAHwpP8dCYCkSFEsORXF
lNUaVs8dQ5gLVDvyIbxWRTFAa6sqJDKZKWFUmVJ+9KIBIx5K30GVWfZ72UB3wdeXktWd/WdL5h7K
pdsAwOZuO/jQO0UwGi35ZQqrQny1Nv3Ku/G0Lk1gf5Q8KtukcAFMFtdb0WsT4mf39EVDiVw9mHSX
mjuYhrgbU6mJJydD114CX4yNGujcjE4z/n2VU+WNn3o6ZMsXGvNbPbwUZ/l+kEfNKbcylENZ5wit
62D+mPQ1aZ9DQPs9URYtUGglpUrEeNOPT14oyQZUgnktqi3o3ZGr69XfTb+AHPD2++ISTbOkdB+k
UMnxYPuzwZMaq95sAmYLVla5V421toIUrVjLbCLX4tBTYR8OX/me5fv/USPy6bcHOn8jRo22cVbO
8b40faRumOKfsGOtsLzIfqf58pwd5WaBqv0gFxGcGJxWLDoytQ9QPkYKK+WPp9hTLCyw4wL00/1z
u03jPGkL1+MdIwITx6iIlX9j1vXyIFjZbq1YdkuvZsgeMupSl0EmP9TYCvFYLU0e6pKQBHhiONUk
8VU4RyOuwgA1H5+cbmYReRSif+Es3Og9XElk9JZvrwvMTPe0l/PCes0QH5mjh3YQt4Hupqsn6gam
bjUWyRiptQ76ASdwneBpxeEnY3+FkEjhMYfPbbrg5yc0w3U4rtQgTwANGItkuuLGjRtleyy0coMk
LwdtS18QIlufJzfaUfgl518wMzUuqzzlCbtNjYLGf8+zpJrxeveyzR5VhOos9jzcaoXyzyG48gxH
sJwQVHHN4UkORPhn28cUWIIxW3szUhhvkGwsmdA6Rj4I9RvYU4bMz9vMWCQYrawGzx/VQPSGli+e
PrgGbI2EGkx2UhvzvT+mAcqV+vSYcIwnYgx/0+6kjYzT0RQUjDm+Ppdj+Yqts+PyTFM7iDS9wTEZ
zRZB4NwMBLjcoDlk7SRriAucAyCEfcxwnhUsYkiFMPdsdSZsNsG8uR1NjKtpyGeMXnzYRHZ1uwZk
c9BHgpbcQO4D3aYlIxgH397ZU+xaMgTxKrjcH6SOA9n6R9VGqnU3vetVGxJ9uXVpn4aWCG+PXbKd
y/uv3FFEyZ/UqCN90dTJ3yL3mq4TJB5qWrD7gtELWpCJl1/0vFCqXC1H6pLBeNQJLoey1SSS8juj
El39zAepUygGJ7sIy14CEXEpuDpBSAjjgeySne19+BaivVgU98oNAgYdsbuQEY6qvxbkgpvsxu6p
l6cWDDMys00serwDv8EXxl6EalamJKfUZsAzKvcO2lvAYplGEcCas5f2VxpiVp0m6C9NAvhjkv9k
jiOFbm0w87KyuGSwOdaLqO1TvTaaGN5PtKON7nKKymITVuJe+spl8zfhnmhaffBayNUaTSXp9/QV
LJ2U7ja/Q8JzzGYrx5Tz6zN8I/RPVYqfSv0ifdf9mh2W8gNisl8VsIxnbkl5CZDmkgfmjH6W92ai
PMP0kUnm0rFV4iZyeOGzZ6UVHtoMoRrXc5SQ/AipDEzHKAIZl2BN1xAIeyT5/dyPlotBTD/53yeN
LW+9wKztAlMN9X8lvbGp/FwbULsS7FrLAmKthpfz6r8TGOw8s1023p4x8MDuqUlv0O2nzv/YaBib
xSUJVY20VomeQfF9dsYqTq6OsueiIoRUa85tI01JKnzQIiVnoKNzfQirYcI4ztEhqvUMawAoKJqi
8JVCWztwPEubeeDMmdDSqU2P3OdfGzMc4U+9zAB0wlbXCtJdcy/O8iCHg4WdvPZ2eT8Ozm60slBg
XhmMeIwRy33eUfG7Cy1m0Ox/cE0VCPPqSRxvxAF+0OJpSMp6YV2tUoLrH2RsusuySHT6K6NK+Uwg
NIp+tfd138AExiwTMoNCS/he4nJAbewNiq0/rp7ZqrELotAjkc4G9iJlUb+nHoE7R3KQbEdCpC9s
3VO4M9MKXsflRh4Dw0Lza0HV/2WILH8pTe9czaKd8rrxIDcXQgb1uUO/Bbh+g3HcCKAcr3RGVngJ
W9obFhMBjmlkf0VMb4YS42f3FvQH0iOYS4v9Im0v+tkAYYeZlExFktTOjjAXrNBQy/m5bG5OjKUo
mLMZDG31rZnDw9eOZX6oj1YjZ1/QIdXHm3IySekfDvnbJc0AQYHlDeWZ6SGH52ozgLcGN3Isr4VY
GEuiO7DpeLc/2VB7N+U2B9AhsoB9EZZ4rxOvKHyCS8OPWBUPU3y+jsYPb+yD1p1YcjvYObTFf1Qj
cclDNuXcMZWFMBojVMF53BPxl+sjcYQIDi2+zXbC1brhArWuby6ynjZD4hqz5NHKwUMfEABVLkNp
/2ANi2Y16YDjHH6vTeK3y+45OsaWkCPZprDLTbX/R7N8TQJTe69FTriC9bd1beYnr9zxc10xy19V
25/e8B+5K56j0m7c8muCrRnlUPVbbo2yKpfg/owziXBXj4282IBUeoRlZNWxEjCGhruU3pRSsLPw
OB6XWwic3oR9C1oidqDnTg+eKIW/IWMzuqWztBt5pAVMRxmqQ635HcjazGdjZSP8qJaPU7uPfaDG
9bTm37rs88Gl02r4wN+ZEEqHzBmVFenBw3gA12TCTvCIBFutVLfRRoELbLBopfhVBxSxpF0yTzhf
yruauedjV2AEoav1aqyVXZlPVLzOJmKnDeKImkjpMmahykLhKDv4v4njIy13yVKrTkAX5+VXs1gS
ph1EDw68cK+EbmDnWmy3smlEL3AVgaddqW/ZJAcjEgnV8vFMHfGhyEn4dQKtH8kChdNBh+T7bvSO
I/3no03NSGMs147giKfOw/59IsYDT99Gx5GXiO7rTg8Hjg7vJgC6/14BlWGYLYD94QqwfphbXbS2
lHnV30mqWgTyfX5GbbMkkgi0pgFZclcEZopkFQNzAxGIMo2oOMk73C7TkzC9gA+pdZWbp99J9JBS
jxu0z/iJZctMwsDjlj+Wd0bbvBwaiT6rt/92ZQpuL6Dg18AQPU0t1fbXHkXIc821ENLp6kfsvnjz
i6/m8WMK5Gxb8Fy6cDMSsGYTkjs4eFm1pnbM/TEfkYqDXLXD6/zbJflQ4OV4I66f3SdYBpx6gXxY
Di/04E6lp+5pXz2/4LJEit0gkhzJlBe5b4vB7V0v+KBet5JmJPCcl7azxIW4pbAsCKkLirchMaOE
RaEqLRZFqgGiFcEQ8cZSXZ9gzMbjpNJ12hIhlvvn+T/kH3eEnGCok9kkPHmqlhgGOQHzt29Yvz2M
agOrAJ1S4k9kAmfxmZIR3hhSpbeuoOGuMzl82YLNCpcRBsqVBB25JdSnpXRf1ZyKRaLsfvfUBBMI
thNC5ea403R9jaF400dMq583Y4B6XG0yo7g/L8aERoSWtKZLs8Zp0kpRoZxIpEa95Pfu3XXj2YpJ
hT7xFdaZydDWdPsxO2h3lUSRCd3gDkle+jdlP80ZIocjr/jqOCOaqYsZPacw6hpN7yO19mike8+/
XPotU/4UHju5sK9jZQjKTQxp99AWhO/VN9PjolnrGaTJuS54AeOg5GYwqufOXQo90p44hMOfINiR
/Ac0pejjZAN+xC/Lq8Rr7GHd+hWt0s2qOhKSGQW/XouTh15agiQf7U0ssVly8hRsHvYHEYn+s1HU
eYzg3ekKTVcZ9OqbK81c1ty2TdjVbZ5hJvDazHY3LDELgC/1Bb9i27XBWquAY1wKp0jTryX0KChd
i/2A/5Y/hvGKtrLExtMU4FsOP/ruHQZxEroH/o7+exKT/uhlG4FJFrVc4qeGisaJxo+Fs/EV33wb
nu6Yj71NrVcvddLkYTjHOhtex1QoC2+NticyCA+nmj7kXxpw+ynFNjYnFKhHVndxe9PUV3QdfLSF
pRQlL3P6FVh7vO4OrbNvXvksttZqsandf2A7dosjJT0SLWmIgybLUchq7jACTll3ELIGrt49tWlR
unNNokNu1qYnITWvneRAs5V5gyYT3ffb/qqZuOgb7jKSQjtDuEycBLb8SrlnM63EDA/dJ5XCTMpO
Rs53QYmtoC3Jw1DptzBi3iLf0ppU/5NtRste54J+bN9rlF2lKBFVBvygZrchFgqXuV9U+GbZOlkv
Pg/7Y3W6451S4kSK0wzM2A6c6FaQEcRKC/BWOlioPuCfl+VkH1UWH4D+vVIedoRQvON8LUOJ3erY
4w3Jn0pGwh3KN4IsO6oL72FCJYQoP59i42kDllBojzJBBrUhCTIi16+P2gxnwkzSpR4823cKsqUH
UpH8h9zRcZ1AN+zIsuR6x7Pqvz1YYVYsW1zKwCWN40QEYbiyuNuYtMkehGsICFyfdJGna1rcVtyf
6sM6qB5mFWFTGkpamp9kbFgzq3AmuFwYUpdgLDjg4mBTq1eQJskAUuYMR2Ahrrhnlw1kuj5eskEk
8hJH2jnp1d/f3So8cOwWG7AkPFGWST1+L3RAnvdtaWqPgtWSyjMaPRD8o9IzugsiJUhr8RZzT8Fk
92UxyNz1gpBZ0bBbtI38Rina9ca+nFQn8TKcNVDP1Qp3EwyyE6tr8KzxA6htav40qpo/afFQPFxh
0Ukq0NvVMk4It5WEIoJHfLarKXIEWEIBGnwJmiO+M3tk7+mxo+eM7oGcjaM8ktmyCN7FZ+mt6ZkO
MfjEcPaSxCHxcC0yeG0ys/QYe22tPE5Bm8fY3/DJ6JYQ8FwUzxXpX4br/Ns6uS51kSPkBatfwNxQ
r7VkudynNEHa1HxwfuVXHUQliktAfzDgerNdWJQmaWcujeuCM1a8NUVdWxItNfCNdQBSmu7TILZG
SqQtBE+dPToH0O1HDRdQ/bt5RV4JzHOd5qbYEujVft7v+g4dwQbUfwlvZ/X5PHm93btWi3FF6Pk7
iaZlAd6xCXWq/ZUXXxOpVmMHmN6HUGTblGWdWQtQmDNY3Jedw+81lZgepqRmCR4TCAInZN4UBNkd
MpM3pwdemCjGk5BpL5kU7zozMQciCVvAoUiA19LldkQzER4WjTeHvxgbp3pNapYMmEZOvTHYFAB+
XTRWKxVZoFHwTMa75dVBCOoVFtShW0Z28pPmi3fZhUddquFqIctH7nrq12v/1BtxYLrN5cknXwmz
IzUu5ZVTYTdcmI+I0hzFgIM1KfKT6CIuyC5deZaGPUtYfd9ybg3jYaQRnl7xcIj8nxfMIwRCK9P8
gPndY8X+7KwOX7Z9BhRaOrTs3hep/ePUkNV6BUtPu5dIxmDcSKJJgHAo1+9NAunNJVWdIMWQlq/z
eGZFM03rSXn7dHDxQsVrSuvuPQzSAlfhMPXYObnGMaZUUg1kBqvanQezjIZ3Q+blvFLSgD17gSGQ
48FiD5ZNVfeGr1f6bamNl3hsU7AZO7WyIQjg8zmdsMMNYnVT7QptbyID9/qOisBbDQK/54RKAOoI
8niL3Uc2ncjIGGR8cUJbYDDZVZNVXx5FuHF2sTBTD81lNtsxiiUvuDwIE7vgnwFVnPckX7kvUzk/
owEZYNte+3BTgDGBYi1y58xqq8bfBD3FFXDCCoyaJQ/OMfi/4QQUmieU3TiJ2wFTnBogb5KZ3pnq
Z9d07GEJkZPH/KycxnHkaaeXlGtjtcQ3eKj1I7egpoz7d7f+EJpO1cg1XQuj8USwYrndB3p2Jr0G
782WocP8HYo5DCkAuL9HDX2KrLSojHUsOVXwdgEGFLI1kBXrU++q9ppGN9AUTC3fDhAH4SPa/GDR
pLsVrSIQf/kCg4iq+edtsG4tHSQv0+/CZv1Tk3dJHW8vmmuJ3tpgXNHTL4zjFxmPWUqYNOyHTVty
mDTxFrwzBM2JRyplaETJXVYDMk8jBVHvxA/FNxK1snsgKfdy0bQXGTYRSV8xiKRLYUepLUTyPfAf
AFn43TB7R1jyA6nScTLqW2oeaaFnFASZFqhkXK7bMdKiI672oqnSDEdgNUm5CIcj21qqm6CxbtHL
BlRm7fPP+X50laXvDnzq4sTSLQY4ksgtkZLXQZUaCNrXwC4/GgUrSS5GjZTabO1w8jMUqWSFStak
5HzoCw0o1m48dxfUJbQKr17WvpGUqbnt6/c+asBjAA+MRoSsgu5o1gBpiyZ/tI5rGN9kgBc8Flzf
3N/b9/3UJUTnrbGyv0CCw/kyZO6Ds8tpUysAbbH5gn1adcu86lSqSUwbzJjoYMhViVpZQ2t53jOg
TQGTTI26+z7mrw5POi/r/fNsKy3q74x/C5x2JOAFgT/ZVSclcpL9EOOX3xCDQVmpiU1lGsuO6Pji
akzbc0qFQ1106hDt0hdAp6bQGij5da3D3jsq7fqLHF9d/rWHv3EzkcTDxgXE0qnEnogJw0YqNwA9
J4uMglM8ixat8i6qAdk/t7Jh2Hig4VaEOqt30eCoMaT74Pkl0dslHWbvs5RX9OAlqbYzrLAzgxe4
1uBeIgl/qGt2b4D4Di1FJB4q5VhyVkbAXwwqKl31GKaZlXy3WFZ/w2ul3UstqAEUVPxsr0TuoigL
arpGpyW2FrVDiEU1ZAuOkazaIvdCDJyc7lFnPG4wELRgUF7+dDTLiLf0uiMcwOI2DYG/RIQN4j/H
/H0x7POliWnDGJm+OZMxh/9cyk0c+mvsK1rZnnWXt/DTfKcskp0nwVXatD6ODgpsHwJk18yQC1fo
5E9v3xGUZvujkIy+aShCbBjg1264Paqb7Mx3+JN7scx78jZ/AClrtDjqYjzJwVdQYO2W0F6wiFO9
Qg67kRZEomtcNitl42PrItW1JxbNNgJJ2VA342yAEUwdwlQjZFv/gbw1kT9rREpiw5OvMK74AqmV
INNcp5yDPRT4tVxAVVX0+com76iqMrkyp5M3XQv7NTnpuComuPfEcybE8yiGs48Mp1pcYesSaqjt
8e/TG0vcr34SLADWW6TxZ7pmKM83Eveyfie88K1Ri1SaGvL/042xXBzhF11V0qrV1yLYzsgn/XD8
GUnKGVS6+12OXPeoUbKfD3uE2Y62Hu7k4jTQYKtZNWXm3s59r0J7PbgQhUh9xOjs5nFn+Tv8N1us
eF3QJJ86em9aH3/qWRqMFfX4clArQIZ0dw9tnx90xY3MQJc7JDJRbyaeaIzIKLnER+y/by6U7bjI
GVsDeqiBV49ALOX9eYg16nndjgqpLjR+wFEMLSv+KqGiIYZQfwaNpCElraVZ4Nv8C4vF13OH4UWh
J0pI31nxN++szb0rlOHIowPMMsSdLFtxSD5IVsVKl3bkk1iEHmjJ+UAcFS8NwR15s7D6gXU2JHfu
ogiaC7wweyCnaoR5IDXzdsKpY+kcJkop0zczLOfte3jVO3AU31HlloGlP7J6Owz6F5eyxpVxTUBW
u/g/f/u7/ChbLBN69eQ1wLX4GYTasajzsR7qJZkt+l+1I5c7CbrqT9XFIcmpK1GVLziPwjDv0lE2
Z6iui5Ejuzc5lLaM4FotQ3gjGItZy0ncemuCkkIKD3H/nV+O3cqE5EXsExJTyUj93HkfEFUOkCkS
MAzw33LlbHJUK0Utkr3HNkaj+ewNet+SfqFeK0opkPFL32vVgKE0hEEsy5+TtbOskKBO6ZJU39Ft
W1koCQIKngRUMqqlaTOD1kWMVkeEO/20rAvgcEOYEq4Fz5OaHGQ9jwoaod/gLK8RRWQLrP2gzuzU
tam54mO2CTQHh9EOWzb+FNszrIeel0HjdANSgYM2TMJTo1c/vNTYihLtHOf+LZe6Z930zGTIDz5I
MEenSww971AeRRPHZtyUcIxKPO25xQPiAGGZwxcWkmHHweoLpYGUPCI5dTuu03eE6lgTTY6zj0m5
OwwBcX7LjM23cr8VYhZQHWVk/k9SPlvNLEvz8UNn2wIzR1zqBW552MLtG2b5BZMnGrzT1dU+Hih7
0+Ch8+dKN6WQk6tmX27fT+53fljugK5tgnyqSSkvTPogm/jeFHK+71CWMHyGijnKToBhz8Cm4eOj
ixmX35yVyXBVxxdzVdFZvtscPcw5QzDiYvrl593wygMuZ21YJArRPDFRpjY3PINRleybrH+f4j8i
E90jXuJevobaWrsEGkbnqdzSmPkJi1SANMvNl5OnY31xCpnEa3Z4dXdeNPRKhIUt51Q+qE2jY4tw
uhaV3t7qOGfKsUUtKE4sYQUikg69HtDrzz8bylPQ6wZ4GW26xmsIt1JPQyki3JGKzMm+IIeqyBZJ
tzjLLvCjzdo2d1fVIIikOg4sJeepBocaqMpo5tJpSgD8t/LfBUMJUG9JohiqSSQA+aWQUJysR/VA
yg1PveZ0FZqM57+Cph2jUgAQ+B6Dpr7nVmktbmRUu/pAj+6YE0V4RiLjjVV24V0d24cwKe4LI6Um
0CKj/WmDX8Et2BT8kRmI2h6s/tDoHpN3XsxjJlW9LVVtvYeS7E9YMv3SXQS/rD1njZ6+588shsUB
gSJWF9x72jLo9383BOxVULIRaArmXwZR7CO22/0U3B1x4N7Fxz4+HZRYvCRpibR9iQVH/NCihiG4
V4d8TyiixLrSNaJoDOXoCc/W4X31/V5m1dgbEWoGdMbZEbk6NXBvhgsOsTz88zr5eVXW/X83U534
QMdzlqGp+/c/+ngXssNVsLm6OGk85mpNsAj6i2ZvS9jL4lXv5IScXkhTOQ50BoBPehHIbdIc0E/x
ksMgG+xAUIWGohcdafkIMIZBY5r12aBO55eaWGLR7UgweWV5ar8FfRWXXVZUMCPzP8DdU1bheQBJ
PeUVx3/+gYwBDFOPxxK5NZKQiLdmdulzUzDc7eF3Q2BmtqLWIxlTZwbe7o+kwXpx6/0Zj6x8YN3i
BkjWLBqbdAAl5QPHQJhVIB9Rrjj5EP5CNR1JxsSGYLpF9iAH3Vvh4cfm/uSbyYTsr7qpA+eTfEhi
G600x09fxP2ncVFOz0SkO+b0Do62Sem4xPKUcuVKx3IrHzFrX7+neI4tmVOro7frvwAnJYb2kUHu
ELVU/LxIxaZqLKMfTfb22+lyU6zicxgpkuXKPPY11gxqtBkwubIvJ0Aem9/7mTzpK4gfEHoHl1kc
82sD8pZbB0Ve2XiR1Iy9QtIpXQbiez+gD8J4VMqE0Gz7h6yczdHCun5GLfPve8+Kb/8LxtIvBlfP
yrmeWFDKiNcCtjwzsc0aD61w42LoWPfiyRvYyKhh1y7Qme06Y506zF+J1IX1E6C0XcD60t1vHOsP
c2/ErcIFqpGPwKDzCmBD3ksbUO1hViU9WE9/yykKpeZ9MaNwJ8KLtu+49dX1QtO2QPC7wrKldYh4
3ekAAB2szRy/wfQ3vYNb4fWxaYB0AXUemC0zqYWjlLPrk0p7CyZQxrClTMGxp5kka1RJiXmGqfHY
SO1bZO0Qk8Kd2FKdUX1cEsg7cH4Ld91MFZl3aK8uXU3z5zJMnlBbjQeLkkvgXXfXP59t/sR6UvKC
OPE9wcSM4tN3a9O7hUqg666pZbD0BpMYuaLaPITAcmxkIPbKW8CNOnynuwY7ibpYkVqhSgyjwT9G
rWEaDXyXi8A6De0yFNPUD/7AOtZXOhaXkL42UIyEJFIhcAuy31cIQ14zqvJFpMOYsCCfm6SayliB
HfB9os1zMf/cWxu2t5xKMvNydxMflwk6kPiBbAyWVzPHkACBuXFkAxO7k1Fux9jeGUM13TaslpbU
mNsS1tq/IlN7HQ8stM5Kz9QUWccVxRyj4lopMOuJe9n5ihs3AHMmO5zdv32bnBkMlU5woU6oKD3+
t9aNNHgzOjJgGe+8BCZNMx9x1BZdhCJ6u8Mqs/02BcRdmuWfo5KKwMdTUkzmcnF6104j+05k8DV5
/dBX6IXAVoLpYDAsgr4GBXneRpByV+bIZhinWz7fYp/nKTgy2bqyKZjkbgGZuX0RixSIra33hsd1
VKRR5WmEN2yDF6pmvn6D8Foz6mm87Nl3Qv+ivgqHau4XCPpJvgdChWP4wHMZibkyRQyki2xprCjf
BWJzbEBfiIEhMwNvZBUAeKBGg25cdQbpUpo3kLDogDMc1UuEV0y0r0tkTfVOvbHGirflP7BKvwpM
sanJxQPSwCjngBFAXH9K2WoVP+xPRg8GGNCpUu6Lm/jCYsZhPKV2o/pYBw2uIf2cNkLTeg3vHK2J
GfiGU8VZz9pyxIbLypp4sklSGM60e/J4p9U9/I5Qba7Z/IVKNVUgVDxWvYHTOM8JL3zcv8IWYRG9
WRx+VfZSZwAXTStr367+a+nvkD58d3p//u4hMQ9eMDUc1S+3MnXNJ/WUFMXRHBUSHt64QnZmNzQi
DJGAnzi6NJo3wMAPEuABpNikhTgdviY7NxKFRF55+lI1c8OY02jUa569t4TU1aQxOqJfEIwkryys
fsCricR6kcqOvrhZU5KMKpiKp4GSQdtx85Xhj+WM7IdDgbjZFcHAaqRMFQFn46fx1AHga0NSsysN
Tzoy5AycwzfC+4w2rE+v6BD1MIK3EwByLwXyaKr2csLPeSFKFKYo+MeWS5yJrB6ivCsQnP0mQLhR
3QN82zNk5udNA7k4IEnFphWpzv93EfZlmF1pzHy0jqyAg/+y1tHjLg6LZdE4ULHuvhAsw3XsNvuH
qKvkyNkXK6hpk4y7EFrrQu9suOKgWkhCDavyxLptEWeCqbxX/0wp6Y3UNvC/ri3NkIz1Oc4k/Bf/
mxOCL25z8MRFVxaN92/EvNxsBypkDtHHFUInQemDK4tEGEDxrxF59tqb66E977Q3LuC9jQIbn7Gj
q7UmZD1JPb568m8oJe9u8ZwkLAMLS+QjimqZBB1bHJ79HkLesAONyCOpUE79qxFpvxhgHI1UrkBt
M2vBpESqfMQP6jUPPqfWT0z5HQ9ygymPIL8GYTIGL5czcNkbkGksBSRZFqQnzqCGmRY+Z39IOyXH
R6UoDxCNgJ/ain5UM4a5Bi/GagU23V4zHelT/Nbpk+JShNpV9CVpQGGApf1HHpUxK1XBLgCpEvd9
v0TU0gmZaqkrsk8Zj9ouDndSU+X4II5s5id+PmET1gDyQ4HIx3AtOkaeo+L951D/MpcIylO4ByyF
jl+WBw8bBk60G3GYodZQGY5+MrrTWZ4oMaFY+VwCdnOfNq1Zl6CStMLQqsQ+HgMwvlRUV14NAPIZ
l+YKjxMWxpBJMtm6WY58KgY9Rt4UWrit1zsmvBnVS0kEwq1LzrZkADV+tWiO3yLhr5y4vxUuceOz
AhzI+GseFulpAw263RlqaTt95Esu7lFjfXj3jQDo1Ncu9JLwXOvWmDLeorVmQg73gSvnaE+Dim/J
ERvpGm12UOFDFK1LTIYEsoNnQsyegm09xsCQUyNzCUtXZFrX8FF8ohk9gARlWY3HLnm84tUUIk3X
EXq9OsO/TGKqolzvim6mYfny6zi2757+MnmfcvWWyaF6E56bkZjaGm9Crw7tOGKXazvwRk9ZD9PP
t8s8lRqNitGdBf7ba5EJC8wo+k2VzDxx2Aq4IhTfPdo//2tqVLcsSuhs2DOI3Za+y4OATPOgUVvk
luDYNZ3ERef01kQxMIwCsPLyL81q754IYFHNWBF8vFEsnONnZnOjLye+Z3hrh/Lp1cR1HWCBB6qu
Np5QDLO+r0XrS/iGTZMdPHB26muWN40I6djeypvVBDkH47fTAqBWOweN02YqVJxYd5TljywYU7Lk
XxvibRabn4VKAW8mWizAD9NYxMxZWBf4qOQiCeSFfefrOpTpvBXt+oyu90WsvYSpFRWqDNnQaamT
PvBGGZioqhhvB20a0fMF1N4DqYSwWJumHoj5eicQz83s/o5mGG6ExgXNXJ1hmUTD0G/4HlRjaWkE
YJR9EgBG9bIeSF4HH3CM3hC1wWLsvaZasifSulOO/XFsQLmwyh3GYI8QQFwp6UaehKCs/4htS4fl
SqK0LiQBPnAU5yEdUo1+5MFR7XWlnIq71nkvOphqJH2a4qfM9+KbRwuwzMXkd/w9nJxfWlDb4yV7
9j9dsD46NBLC/fUBtBtEth/bW6/ayhtD7I3LxYw9m8irzbO1B7JGcjTEBEJt8xvKaqmiDjqEws1A
IbF5SlLDnunj6DFvw57k2QFe3FsZ32NK35/HzoQUhdQY/+qs+uQ3bTCBDy77jL2hMew/ukfXwp6H
IGQwj6sWLfE5WyHmniKhfXuuPKebOwpr6YihEOozEph2IorI36w6vA3lMj0TN1tCSio9NIT9m3l3
vmBG55MN74FX9PhoawfqAaifX3/XDBdrhjBx+0goOxXCV/CH3nyUIEtkx+J13m+PTA8KKr0qdlEq
1MYju+olZYBYdyVDvHQny9R8cXPyX1lHLXdD1lv+g0uIpe50jLgwrD5JWhE0+DDyRQ23q7kbobc/
JTIl6HsOu/lNnEPud8GE81i52lPpruJaWVjrlkPADPU1LFR5G6lscjuPwZEvPGUSn+gbHDuBqto0
KckcA5yPXB6QP6mNJdZRpnzCLV1TgkfdsqFgsYG8qTiEC2iFE2i+H24VRHD/YFDEIpWQ8yWCYeT9
EOG8KJaXkEuq3mz5+sz4b0/VatlzCW5EYuamCPuKGFz3xX+ezPoCh5z2vepVn7F4nO7spqN0fI7X
CU7wNU5Gzk1UOdlXAd/2PtQw9ZTXnQQ0H2ZXW7cBrc/Zw+xVXfvfM6youi8nywGdU/cC0Rux5Vub
FtzrAm+RlLOoqGHM7+fA2GwNHGB4BAQOucnNM9ut/ySxXyDWcIkN6C3W4JZsg41VvIBKHyYXvMan
lqvswkegWTQu54QBk8oF5qKK2EApdlSYeoBwR4x1uczWE8x06YxUdseVbJfvI82coSDMI3aTcqyM
jhpkavTEyzjGTlGaTr1qHoISpoVYLvtN17pQw0p/lCQSjiw7rnSh8JYWZnqUsf1vGOJsRGyuLFpg
jxziJhBzBImnXF9gRPbJEoglt3xt6GlqAMB26XL05NLyWhFztSixY8owFBOui0CBOOuQ+h4U+Ky8
TxVaYE0lK6Qd+8And73JlZnD3Pc0HTbgsJ3/jWHUIfXtI2iNAglUvXJnfyeCKYE+2GdxO0OU0i8J
p/VIMUKUEJ9jgAHGb1cseESq25LFg0nSF6kolyOKcBdJyXHb4r2Ts9QUWKsgWTq1mwb1r0DrTdwo
FgqvwF4l+f+gL9KmY+DPbm1ozQODWIwJsMG0RsgMGK8VwSMNVlHolxqa+D3nNJvdz+GAfshZ1G4W
4YJ0bP6MzEAo7Y8SY/yzqETA+CvCSd1Ep9DcVXPsJXHhNxHWP769ILJQZv4VX/J7E8DruSH2FM6c
icwyVd9oaN7eB+07fAi2+bwf2yx3hhsVw9sr4AOz/zqDfuPeilTNxjGT4Y3ExnAKaYUEWGLZGLJp
xw/ft5PB5XIKvb+F1kKAZKD77D7seT0Gi0sSZnGbuCYdJHpZirV3JrV1AdBaBrJm8ApQF1xR6tCi
lhWd2PFkmSY7ZjSrwrCbdUUrJ/4XQppe8kJfNU12l5pLovFIyUSdlfgGHu8AKbTikMpXsrBqNTCE
oKQcclcnzDVhkVIEphYYYrOGXncUv2hrbx7R8F8bgbNk7PQi2P/9SxlhmcUf/078gE99fmW6nH6n
c85mhhkkY1e6TMO1fV92t8qkbWCLPbRcLeJ57RLKlHVN67VoTr0PEmY5KXzrGanwSCFKtqCa7+YY
fUSxcRNNh+lP5zxbidqaygVpiumFuRAo33PKzzRIQaLyti9sgjs8JQtmIUd0G0cLCo9yWJ/IosMd
3kBtzinA0ejoDK7GY2EHLLx2EXXeDKRHDHVuR59CW87mxj9/TQTEbxbF1LdLrpfY7hjZ2dZYycbN
vQ6wdeINGPE20I9M+i/403YhW6TomyZvb+lpeK9gl3WnW/SJPMHztruYMVwWIn1Fo9pn11OFwxzR
pJVnNKgQGyBKY/UjAzQT4UdBpMSObJca7Ws34TeBAlmb9/E3+8naiqPKnp7onGjyd5y4ev1AShHP
Chw0lEq0cOveyBW3bhZUG1MubZtxdze64ptuhxkerdT/InzBNrsWAkldLgHXYJ6SF/H5Ud+/SEI1
EQfj0iW5tCf+6KRYaGzp/wgVcOfopR9+GYIrnannKVyLKQRb+Ycy6oKpscnP6o+INbRkcdf08EfR
A00iQZ9npojN2oAPnjceMtoliVu+PBQU66CZU7DCsfF4YBYZ8ukg4O98YBYjUAg97hwEY09ALsK8
xfugL1f9oAx+b8ptcpw1zCz7mNt53qP19PRwMv34/kVn0kslvBpoDqmKS5r811HA56wwMoj8Fk6I
3NQDxaBkoaj6zDxPjDd6uZeLO5RVrG54I3mVh/2LbcRvE8/Fob9cCs9K8PkkfAnZJJbgOj0kDas8
Y2bEDARJh0g7PsjgGhulydOZC13TyWPGUM8JeObzz22raOIkc7ZNsWVFCFX9kRwoIBdn4y5/ZTgO
R6QRgOcb/aZw90TN0npLrDfQG20xaONJrll4/dRY4nh+DsUIg8sm9zMv8ZjbdF6oCf+lPolVQ6Jp
Hn1T18hGJQdyQUMfdVHpLX/h7mCXXNgQH75Si+e5TzGiGzA8aSQ3mcdLOWcvd79Zg5YtjnSa9qkz
+rnn+k79th8RDDGyKq17beIXfegs5nJrNehxr7ERosY2nFQiIJ/P/bMlEFM4AtKxJfyQKO7Jb11a
OsZIhKR9wgAfrDSGAagpfe48WfRzoJFdRluUA51Q8iY/URwCPa99TYLkiiXK2CreBkalg92UmItD
pR02l3olX/N1MCkqdQo/raj1FAbO1CI9gxmSN0jovi4GQHnZ1+NeoiDbAfRvOW+98bLqZIxGzPbY
H+S9qBGoYtfgAv+bj8ohyGR5OE1qgpAbrAgZBXMgZ/DK+8XVTozbrr37lcc8Tuf64e1bqWbiFkJ0
nM2P2q7Gd8zj/L6tm+T5OlorHPOP0/oUrp88NA6/xU2UHso+iosY3cC7MBiH82TSUxjyGuo/Vq45
CAN/mFLFV5Dqy1lDX6BOyaNROY6/INWsKKKbpHCXXrABOXut6RE+sVK77bM+bG1HwDmaJWz+We6s
i77nFna6Qni50IKnBRwFWT3mLPN2tVlQPuj6izqJ8VYnENLlF76CwoW70LbhPZXXqku+NtqhbWfP
TRYmxTkwfI0gdOQC1TVwuw2yYTk1G9oVmsJE3s7YsIP5y51ZiqZEaPT7PRQtDxqrsELypRNyruOx
mda4qKIXchE7xY6QSO8xzS/gYfBmGwo7OJl7xbukhyYbtzfZYE688u1cXhl0cbAN8GiLErdXJwyY
GAZcd5HVnDiCGIjgMGb9fZHmWQSEsftl0qSt/z0OXDeYxqKLxoQB1XfA/SpbeXOYaOMZF7J0f3Rj
h0eW83aqjNATB8LOzJqYqhH+jiQmWHcoTko7XgjUqAdYs6w1UfHOtO0Elsuko0n7JZapqbUizZHD
qjWdhmB2ELuGUaztGtBnn2LRXNc4/ifiB6eUDr76salifwgWKmmxKYz33PbKuunM2VTBJiEqSU7O
7p1SrLAitwOcTME8E7mqhjpaH9yXx0qZUBi2ZKzQCNM4sYNU/T72q5D6SUNbueEfaMdKWMFNmWGo
enL2fgBXVXu/HyFtVRF/NFNb8kCCIntyQzR8uOfTSHVcXK+1ZLrkpOsXBNriqiIkHk4QryoQiPR6
YX2eOn1lB7zXU4I0i4c3P85HYdu/jGfgEWjszXStQwGvRPgdFEr8U4SgTNXgzsacxNI4ZsyJSTlr
holRROGJottqseRDoW5WiQSs7JGlyIXzW5pwoO+o6EVe3XZj8/QWE+roytumcGYVnWbPk/uCXgmS
1t6tv5G22pxyIU3bcvbX8gCQKeWD6sf8CALbQJ8i7REetgd0o0TJCosEE+mdLLzLNAnR3ptl+WZ1
t9wwzsEcRzUoP8RTVnJAghRO5fEGiAa6qOvf8JMQFNvKN6yi3s2h35z9Es1foLv+pl6qbQ5OCkQW
lQUAZfVsMeyVNARlQcig51hOtbfs/dqh4Q54/oqV97KtNBjXE4TyRYW39IlBzjMISKdbNTd6A3X+
i24aXdk0mRL4XqcEgQvtFuRuohuzX3VAaqZdo93WSQABHo21q3ziJBAOpiZGnpOJWlytVsctlmCR
W0WiN4YRfbG1tBJlcPHVZl6DbeG6GEHUdn3nKd5sLc3OM6OEHmgnvkOwF8lJTqkwBQ/7f4NjlOcE
eeXLU/4dBN/GKBmfezZzUIJn7ely3UqrYovaYH75cx7PJmgTN7QLVjb6JSeTUpcBkNesfLk8dyEV
sP2baj1Pxw1j+Kikfn7jvU7C0ggRInFqaxCW8UxdFcNwMSSMFLY+ugvYxmew08juwNHBdKbVXejy
lKVd9RByQWdbysb7Qgi0E3aElnZ/x8m6RQp1tVJ5tbODUFRuDj7fZj+4gBOUETbdthiegYkBwXrE
6zgJbpB/oDy2g4u3gyVfzRIAhnrzt70wfDRXxKq10m68pUrU7TPythm8NTDfZxcPHJ5+Wwxv/W3M
VFb91nJZHljgf1+iyrWyVSjrObwfxVNdFvd/NZnlWz1A0Pc3uwRVq3C6fmONHDtkeiko7H56LQpl
bs2Qz26wJi4RRWdAVNOi+1L3cfOvehgYMpeRLmQcEzApnUYtr/C49P3Ejyq4hUIBsAkodHEncnHp
WBFnlzqpraPxNgLffNgSFEE+E1uyQBV+M3bXKcwntCU7x+ffX8HgvryjaRfF64W9mXiWmp0fVkLh
NU4Vq8XaZHI6oBUC8LmaZRUFJ9VawMhmbO5fTjRCxSlH1Biy8IELntDtXJvOgsQUkTF1WWgNCERe
YrtPlnktQxjBR7eLdvNO4DZ2kr3DUicrw38Ng84tG2QXj8I6mUgZo4YUEMI/9Bb/SsoniLM/Quul
Qo7Zscht4wjUW8o+x8fuxK1WURaEwOq5Qq5xoTRMnVXg3dllLRF5U2E+DRy1BS8IO85XswEzoI4o
nWHGk8LWXFLfDp+epzZp9pjD1kSJZZ+pkhTePFTcpXX9KiQSXi++ya2d4/3CfDU2OHv3keXw9ZGg
I/keDROA/msSQxn4zz9CvNzyCbccR6EluCt7tWan1RxgOMbHDuB8dVT2CWiqIpfl5WHTzUXhjBEZ
4cLthfQczmuYtjugW2TbpGaouvRJ292JbLaDiZcrHfwYLfMqWJx4LWmmqfWsT+Ig6GbXK7Ez3Oyi
RBkDvuGDBhKsEPLUgiDkYb3XD7BsuFrF+zFsz4AAvRKZiDvJi/53hPlpqNyqme7CNdVc+lu8ND7P
VHyV+hMZJjZZIkeLEbq/vrc4T47IQiPeforT7kZzrTAi7+42qmjYrC1CX/V9ZORNfhnOft7qXLxg
JxYTbaU6QNfUCzWQaqBdFQXUL93VW5nbUtr2UDwX+S2U1pP9Pvu53Rz7k5Qba4PcdJxVp+A3YCvk
21tArPeadQ2Lc9J71M+1qNPk+cMPi/+E/VklY3DCkihwD2ePwkHvH0BtDa98dVtr/QYHuPhOjL1w
ChE0wXNjImdRi0e9xZAlxgOyzT/d0YvRt7h31bWzQNNz9trVxJVxmaw+6XIJx3gKol8aWUheOWfO
c0MP5T9ArholIlnHqrpjq4ZMwJoVhQAV43vQA7wGED06ln9e5ZKnDQNYWAGO0B+K9cueghJuvX85
t3RiaiW2bSj97LHBmDe9XfByy7VCSDMz/Sc51zEVkZICcBgeVMYURqSP61dtVRfDqaorsUmDqDsV
0r4ryheftKiApsg8qWDBPVHjUTgZzUmMMG4uDzgJxl6agfhjOxFJY0vSp6fdjten1ozuU9hTGUSt
s1j9aY+f/ETHcC2eCRt+3S4ktZwrHuI8Yq3yycjAAt4tAfasfuFMwcombvoATH2EcvBEEprwgY63
Nfytgf36jMD3xNPYv2IK6ZnfQXb2MK2Efl5LzLcgKdmCeYZ5SCt8w5p2YT2TXqFdJPDFQBHDQKQj
YjLC93zX/kFeo6nxspXYQFRLgKcKWDjmS889iCxDBdPasdrw4PoyA9/+7rC0ym0wRwazh4npicuu
xnFXeoKXGo4n+CuseiQBBjl4LF6tEntyR0ABa/BrW1ztPa305tRy0KJrKEKWSEkBqPmka2jvcjwB
pdVmCiB/7DaAO9G6prSvTEjSTfUPWBqTySLd0JjhMKsZ80gxFzYYccULzQQD2VfvhWBCapW3knY/
vr3h0oWmQp9aTia2xQNCx1TlU/+qYF0DmUAy45QaRU1RT+3uNQOYszYLkFq/dW/iGU0AcQ82f+io
jhBZf9Rys7I2r/R0d2WrhijyzkEMn8pAaROEKqi8lsrdWwrZJFvO7jt4Aocu2b5eCczrGZFY2o2o
Ovil16N3Hyf7JYnNEC37UTCEz4Qns4dp39O1Tn1gn8VC6k0y3KegjCOt4PH7yejtuy52v34FcG3r
2IkWMaPOS+02JH1AZGPLsSFvl3up8m40s63i/nHfmb1RB+EBJwnvoSQunf5OcG6rJ7qPiUvOAwcy
C/wIy4wBiVNKlgzUqPAr4uTRw8Hq6WXItvNdYvc/XvPbVUgsY96XxbS5wTKWxDv61MHC0ewljSpt
cQJrwNAhqf4gnsvJb3IDrOZ4Gk3Bd5+R3+90z6Bt+t594mB5H1OplW5vmgo8Y2Z1PrbimmYkk81l
LqToYExqdkll2W3RqpE67BdMaNWjPoivUu8ETHbA1Vmde2TUGu3vAuHoR+EnkwChulAUf1paqzuw
2OpJV1CF05VgnDu+DOZkU1cTv4V1ZDfn55Tafo4ndzaTwNFlvTuAzjZ+0fjTJGMJ3MIy3Ibg0AIa
CIJd4nGRIzJk+BQAvKJq2zku+Am4lES5gz5Oa5VCiDDQ7KzznJkRFFv1Sx2rZ71strbVO5EPJgx2
H3+jKGFCaGGZc9TLfRBtwQoL98+J0Ei4IQ/nsAB5Q/jHMEmocwYHCYAvEZb0ECPK3BtsC8z+/qlV
YgmIs7l9dTIlabuY/FhFSKBmXm/giA4V18GnhgA5eahJDaK6uQti+2RnaLEzDNDafmECf6AjmPZa
Bh4YJhSLyRspjnYh2QPhNFC27Qq1HIlFFkrfB1Ls09kJ173Zr0RP78PMYMp4NgWGnEqckCRyPtZl
4L4BOi3+v5ojos0KdLaPePCjz659zYGZ4EkkFsVXFjc7I8SEJ76ZRRolrswaBWrd3y0tdC073GUZ
rnbWtZx9vWluqBip4sa9BY6WwjaRv5tJipy6hwm/BApY4r72oXISA8+ELpfQQV5JjEILMMAJ09Du
+ZR8YvZqyhAEmE7dufmCLjSSqnNbCjTCDw+asaPX5SAZ9L5mlDPsv1UJqsy3n3EApBBb56bZn+I5
IKiLiHApkcBMRBQzto/ECLgLu3Hi/f70HKhx9CVoxMwcQlRIofYGMzf8bMaEIVSmJtH0nUhZrGrm
Elp6B9WVuE9nWTYeapuDMm9LwPGt9t47jfzoJg16ZQhfGOFX/RRufuTddUXhRkCPvx2x6AYfuaf2
hGeGwYlidW6WnK20e2Tp4uSNKjwX4FPeRj54zUjzp2lOwq/T/GeA8ayEwD2vo1BjsCpRfDIty+bP
Ore+z+G1ffWteGzhtLeKErKTrS4EKcrQfMLWl0e6qh6ATN1LkLzWVYY7p5REg5bVEbbRR3hc7el7
kA+ygzROFBCeGKR1h2QOa4vgVlQFdLQ8aqTJ1kJzRR/jEPh4fqr3e2Y9OtZjazfnDDaAZmOAcipT
TxNSVzpKfZcDrJZo7p4LIRBwdU38LEZ9PY0Kj9vBAbEAE8pFgcQmWH4SsBR8MGi2oqKR96J2GZz8
K8rRzNU3vcA/Xn2q7zrFzHh1WHbs8noVPN6PMOh6iS4sLuTO27RjV4THr3Fc61aXZ+5Fhw+mSTZP
eDli3DYGt+W3+B17Ymk8Rx3izqXXzRV5F7312bQwjPOvWPw7Qy2U2r4HmHB2nAtLJkmOsSZUOT8G
tMvhpR1W+3R5xxUgHVX1UYISgbAIdVdAVOsQv4WLy6uoxhOinPiEevXWtJl1PaJbx5RR24yAYD1m
tkC7LMEtG5FwY/9ymxJo/zN+V2pdOTwioBEMgahPhwCG0UQz6+oDAJexVshSKQboMUk+R45hGtkq
q9Wb63H7q/HhLNEBrC0OoeWPa1k98aKSE67788kGo6zw14tdRl67+1n6lFXzwWXRkZ/tt7MoRzar
IrEMX5N9pXYXo6RgdpJ2FPOBDOVGQ+ISBr8P5nRNZ19lUBxE0xoa+nXxkUqY+u9YBho+vT4UJI0E
G8G1qzhGDgGgnVkSwiG2hd9hVQIKUEetZwEvisGC28PGMU55FDcC8pC0w8qPTuMJwlECi9IIMlY4
9MtTPrfHs9L+BAHsBS/THl6HBmre4vcaXSa+rLRCdgeOGXbjvRed66Tzhc+62Knyq1XOH3BBjfSn
qlhdb4gpHCPHNZ6VYxW/m35L8QCcjvFPud8e2hnCKP8lm4n3wuIEWD5NTh4pO8uMAQPOQqltntxx
MADnYCJ/HI/XTm2UC3LYTsoMhAM6EAM094QxAsSMsvfN+riMaqwOv8VpUrOnLDI5xzmEWbBq5Igb
5gCghjDu7ZXp/wq+uGD5ZxE/MEtigPJzaIL+Lk44mQuIJhF3z4DY90kicBvQ4+QEmZQ8jSSEHYxw
jtsudfkJvSdm/5B44tMzlsJCdDedKDZIZHY21SDEFtXFBSf6FAaQEtLUbB6elxPjOpX2/4as4tbJ
ydg0+ZbE+OfWq7JHQIx5tOHEtXDv94VrhsoImRuctXTUmRlvVRnPfeMj09xU19rpwLwmBUz64pft
I+SnWCuoJ4hxlhrbAgSRDQMk5U2sKGAmm++8WXEKmPDQKo/HrY/tl6fNhKOlO9yWrVa4ncvgQfKs
KG4UVwSoUF684D1Vw3GWuL/g7BE2Rn+Qibvb7teUZpR4v+Tdxk4b4PI/X3So9XjsvQi2Pe++nd7F
OpfpVNjA+nCJBod7TX9N84ZVNAxfR4nCmztz2+U89kstnDmYQ3es1bM6IsXcYCOifqjL/GjAav+W
3Kw9YmvuBuVSazh4FrQRL3tD+pYz78fEsx3lOtYEIxzv/5m+sGWk+zoNklfsEkOcCehK524Bih03
6Zb3LclJQsX2B+EaHCTHKpAffIh8cjOXOiaRvF83M0Xo/DU0hLOGPjdQUQhyrdx6WlGNWpxOJaC0
2PXTuA0zg7pfx4KeC8o/LbCBv/Fpze8k1E1/vFiFDI3W4atUyBPmI/LyKSO2AemM7OB+VgqISmQB
6tH5qB+wvGb3cxqc7XEf+4ShNoRsCMEDU1xdJ5tU1vtm3KFDbNV1S/4HtyVcF7PzqQCj4twbqO0l
R2ZcAVGU023/aRg0FLXu7bSjfz9P5VYyyUTRr6CdFU1R9h8zyxZ9epx+i18fOgjcD+1pKWELXzX3
UVhgd8n+W/tgU4vgof8bu4E9qITtGzUkKbXjZhhUqZ38S5/X+MlaslVHmBV8X0ESrNvUlHm/GKLV
mSJTusi62NiYltXtBhXgEFyQkiCbrCEU4ME497MNfW3iXv1sHrEkeSHes7gtHl+oFP368BBoHQHq
wtjFO10PUb3n4JD3ZGrIxNDaXdSgD4HwzaMjiwgdcF9/ppa/r7KD0tVX6MQDxIH7NzQ3+sq11niN
UVCLRxxIrD3GNkBTtOdQ3WmNqPPBozxM53vVDboXTO1Hv3CHAmSbRM00LJVZplUwU4/TcnW/BU/7
odAKTL9Xomug+Puhdsit/C+KjCjI3/vHcY+Hx6hPXexsPQvxzMlr2e+9iW9HvNs9szVqRjT45SVB
mpyDjjaeF8nteBQJX4ulGoe8wxuKazXLLAiJu9uR8eJSdVh3dhmnviZFo0MPml9nk5MPs5TWRXSt
LBAtYrWvhDikufcxgmq0LMCVy7G1rbO9xmqPPay+Z7gQv0mod9XI2gRiZGNSo/6gs75sjRTB/8/U
C5VJlxOY+nCq1ghONRRgukxZ9kQAv4Q8IP9nda3pPbZ94+DfNm/ODvuMfuZ6zlrn66TVhJbhWCha
8i9RHEiQgwl66Nf2gk+tFhCdgpSYvIRoHUMAV4/SxYuHwksdqxgZG9XJb8nzWdRUAZONWOgTcmQ+
BH1CBYRYJ7pYeVQJrSi5SxyqiZHApBts261yluKKWCP60VM2VTKuB1JEEMFbVdmZdDYhn0GS1YI7
tMPlh8Zmh+ypJU+bbq0u/DIeFwc6Gi+NyApWvkCJSsfVtUamLn43hsfFlzYWuTQ1UYXJJmv5gQvu
/47hUvtHRHlJ7maquehH0zFrAZx3k7J7Bd5wflwKQqBl/7UZSfK3hkL7fNrGhMRyx+HWHp/8Dpj8
N3Cf/h8+3wr28CDbhj0fHABHWctGmCdUsmfEjwsGDDyhuGfuLfU9sv5RAu6YCE2ichvCFYEYsJh+
cFO5xrI4rnFKnzYdcIwqeMuCsN0uevCkwcjtNSnVAhT7Utwg9Km7VtL0FeXJvkg+UicO/D5uDdEi
2YINa2Zvh0YCv6q14aS9varYj5gnnvAgGb3uH6TGrXOsvRN0vQkP7SqxC1q+JFevEs45GHpFjZc9
dyXldgpmY0IctBXMb9iP7ICEkxPe9pULASByaa4TK2viJCfiTshjhT88Us0BjGiq/4bz9T72NFXK
pX10N5wrkzcHZHDnnFZbFeruQsNgQ64zJ/hSTJqG70rM9MNwjEFLisK/52/JXA7K3C/PSQ3coNwS
uw5a+qtVIrqyE2SngP9uEEe6oB09G5rJ+obziwUPFQaKe8CQ2ok1Lh6uh6ccLOEPOs9RCs1xNfnF
ppOa8hXesniYXii8ZIttEH9le6tLd6QywEFqWaPy+yh+uZaNjiCpThzWXiKCaqsJmrjJvVSWTVDE
vRy2eXTB9l2crB+M3myW7Y0J6KKGtpzqOFBMDkHQYqzf0gqITrK58B6bXvVvSXmf20U61gAkgo9B
Qnd9nKxpE2QwG6n+YrTAyxbNg5zyQPTu9xgnLqD8bW2rdyaET5Dhj06kLtz78l5GfifI7YcPpM08
fmy+Ix0mYC97Ul+kIW5iYcH2e8VUuytk32lN7974HVVAZYpRI5tEYMinf5CbJMrEQnUZsufhUPdh
8sqjYadAqt4e3ZWvyRky4Fv3+MTIg+q6eJpwCfwE09rAhaYvtzcGdHTKnE0eDafL8raAtDt+bVnb
RMESFleTXtfd4UnR/KEMKO70lhgsmTUDFnF6TMeYyVAMLAARl5og8v7JTHInVBjzeiJC3YRBcgou
YDrHC5C/LUKvCTgWuIR+DCu1zWXMKP6kUxp21DikXIsLezpnF/nnJMc6hUCPyqStMfjX3aUy0oSt
GRoTmjATb8fmAx0a7n+bAT8pxDb60M6VIWk4CdG4YNnRjUd+/s4INWjfL/rr3WxebLskv8/hFNY3
EY7HgrAziyZq3B+N4L3eVOc7Tx5D4SFkqB5Dak0JKTZu9MN9Tf/hzUnxQcJjmugQqlFeAHWiL6L3
TNEb33immIJkffzNJzzbJ5yEWp2PdGz2dUXXzeP/0w9CirBtjykTH9y0Z5NR/e2hk1/QyBhIGY6h
+uAoFBlduvSRZiibh345fncQJTOGJp/5eGISktmgD1al7cf593BwDsErMQFVTDLd3nKhNJzbXhpG
gaApUA46wCg6Ald29WIL0juoEzp0L+3Rmti52kxvJ2dtqM4orsTeKPjP35I3R45yS6cWJFX5nFHy
ovYuNtgiugNhK+WrscZVXF+HHNpGYUpOtZHioQZG+I+rBxckNdeQMwetT0/TiH2KZr32aRd4z9KW
Pd+7tkmYUKKNkhuyq0RwqzxBNcG4hRuAswIYrNEPaB2HKolCUX1BwEcUHl7LdYwLZtVFmO7Me7CT
cvzXlOE1EXtXl4JD+zK/UHDjQZC0yLJCuy4/tz8gYYy1HTOWrha6BbGCTVyYozV+5iZdM/xirdhR
Y4V5Ot3Qir/i5vkXAEXOkpMmnw3DogGw0i4LetOqYE2ytQkY31zeHqnblAnLGwANnvIdN8vAd/Lp
oj8XhiJX9SyTC10tVE4mkUnDX0TJkhjuSkFiMaO/KS22oqHTrKwntupqWBEoE+QtqiqRWAywAJLO
k5tKHZT2p1mQupZ+y1XLTYGkIzjUUQTbiRyoWtDSvBjusQcSwi9UXJpmlxte6fu/2DQeGEdXBJOw
13ZJtd7dvLdNrBn2N7H5JiEcAP0gDqnNxbRtXlkHcWw/0owvhKXfteFfJwTurCVfwp0M4GJueiQB
4ztkowNGbD0nIpursvVpIt+rxXZPJ4nFxpHY9GrP9Igrac5QBdIVKnZdEHR8a0ASy2Ln/7CSSIWe
92rBB2MAgE+t9W1C1WmSpFqe4ZERSGiDNGRTq6vpjzTbh0s2eKSJsJZIuNRxJ1Fxj9r+vLBT0rdW
iTcX5ggDdVFUJChNeGNXNad3Xul3pNWsoYi2Ja8f8LI3RDExoikzIFQeiTCV7mrqxWT5V5zN/ccx
FcETLDrJSFWvtHFuALjNO/ziUdtZZmEXrjNtwfLrRkYK4m9l5nzjKUVyJfzqWkzwl2wRhSn7GGbg
h+AlmQ9ZA4nUEQPoWYS1jovzI0HpXrJkTnF9umkNwER5p/zkZF5ikg15DBJGNW4loNiXPfScw7YH
oL1PpZ1BunwnyN6X0feL3gspGJA7u8thPJtpo3zN0P+0tiTqrXLr9PVy2K2VBvN7g27Bj0XRrhFb
wtPDTcPQ0CqfbFUWNnza1CyIHCCQsmG0J9y3MXTDdeWcxLhZN0D/hm0aUnuINPmEPCuU/8i4Y1CZ
6ebWiHh5ehLcl5hHidSboRBEHjbuhFeAQIjmqNuzv4xr9oEeGkyHbWUNq6NHW16CzsmvX8c1jZGs
QEbhax8ESHLZZbQwytmEeoICCLvtbQFvsW8dRuh2Pzvi5vEhzgPT5lRwoqxLp2ds92kw7lgxxZ0F
jgH0yzpx5XBIxaahmZr4U56DvR+1aXwp8aZEkkrOV++maSSt25uEbUzjGlDZqZQ7EmxULHhRcQQe
LiGTJxrfkR4OmtbNrURs6s3ISRtQ7pxakNSUWAzgQcr5J7u7gq51EJakuH7CoPy2f7OvMJQRn8Sh
83QnEDUxhl5LI7wjs8qUpaJJ8pgeDChvBG3w3g7uYzoZpGVrp4ZkWfvxhGb87jDtXIgL4ZdRUB9l
NquiKGAdjGSHboBY88LU4xatccwKkFZQguB/4tB7jIL9+/+HzkXbw6VqnqVpQbTZunyx6Jd+P/Cc
9Ea3h3ihZLYfxW4im/zbAosSpy5sPdaVLqL74Bn4fznQcfyP5jg2O1GldI1mUfUnd09pyXal0M/m
3a46qLOmC5jh1u9G5rs9nk63+XElfAxkPV2BTFV1szqYezVl1TAFYASCC7wnPzvyeTmsyWsOEU5S
uN6XCe8fqip/pjLPnorzcTnIHxrqxgy2el7HmBgmaZsELJgNk0IlId8KoyCv6gPEvAENSdhjz/R0
niEHshuGMoNfgrfoZZbJQcw7tN/PP5cUzD38D/iBC91QkeUtWMf/+552x6rOlR/XJVqcEkZ/4FYR
7W4ROgpBirm2Pqbv2PVckpMXt6UqRyf3OK75XP3Nt5E/054agk9fgFmaCioI2K+aydpnO5ksj8sp
wj2s4pMWSUo0wNKKsH3MFZnQkp006mVtzBWJS2IQ2Eoj6USON8lpOsluuWz0UiCIrHaPbxDcwZKn
3Yb5kYj3SfnTgNLIHV/vFw3wupI29wtlXHT3MGUB7D4fNa9a+4ycww4VqzBDebw7k7pHAbRuPPJ6
gxcjxzS1q2M7wq15wzxSr9I1B7k9hvc79Qy17bYK2/YzQ2SY3q/YGCnRjSXWYkjvchveX0A5ZcjN
0CXogX7PLesOq8c+YRcxZ8XGl6Q3XnS0E7udMUe3nAAAG3hUhqXD9nT5pcXW6EX6KGEokptyEzSD
u3C72lsL+XmzZNA/0gCcgBJn/VpedCzP1fwGtpjqOU/PzxXHpwGlKRn+wHRYH7/4zhWoJT8Px6HV
oBmlQhUg1aOzlbSct1VxlkPaZ86sztv1nIqN5Y5L0mJSQaYPkSXkTcI2baeS/a0axZDRRkMo/uAV
eePo6fxtVCzsyydP9rOBRLTu2j0QzrI7vDKjx3apB3gIldbCNqOyOfI+GCg/Hj98kWAgZECu4A5r
c3nWQvACUl6dpdLdBUbLRHnLgHbmcXJ/Dxo1SxiG5waFZH1/dLyzsVmMnJJWwnUANz5ZlE0tqzsj
Cv79sTY7Xs51Yv0qWBsMmGf0/v+kjsk3EwwMrzyIa1s7W0UJemh4vhaaA1xjwqJQ2J+hqktRS6/X
KiPuW6vq9o0isGJ9lN5B3GNFiOwiMlCqkVtpxSiRAdrJOgzpR97PdFANQ5yUtyzMwFX2UDy3lXq6
7FpY4vIYj7vExi9e1y/A6oGmuCmoPS2DkllVn4DgOuuzY5nGtO4pMIUfshzrYdiEacV4GXwiGlDC
020CGssr7nV2OxdeOvCGEq0DLrd6S7BxomXZ5k+iGMar0mXLY7cY7I5oMVDNOX41bHfeNqSWoYRr
HuMTDnUVsJRnB0N8tDujEwXOz0lx/VGXy1iKuJJDql0HagCHWLaFN/Rv/+NaudKd+ypN835KdaH9
ZSP386C2oKOHkWE5M335dWuAlCKwNgX5/8b8efUOQXT9ouRGoLoyrJpjAAs1uz7Ct0ve4UR4HppW
czXO5meVuDcZdzB/2kLJENxO8tVoUzXOthlCi9U8UOxK8ZujPZP0Q75uJZjIcGG0G3mWpXQdsQ09
gQhhw6alcYP/MqaLOsDnSuRAw4ZvipLGQ/BScIgxw+5HzZsm+XIrMWjJ6xSjDyc1N1j1F0HT6GsN
FCGcjwMqdAHbjooIsI/xLfAXPKhBpGebXnsrT33MJGYd1gU2UN10cBwTDdG1VS7+1eCPsBzAyDct
X4DKiFEQRznodGYxWoRF+7mJEg24T74E9yP4kHLuNPNPrAeEH9e2Cj1ToX9CI06TSCTDerFxu+Qu
8FmP0u+xONgfFDAQteZEqdUfw2kH+JkYNh6l8P8kLeN+LaPUG0LuGeaT4zKxIXWVaR4+86cHxbhL
y8SN+2pBfCR97G45oMNVf/eNk5GjYLBj/SDlfjS0FTZuH5BU/tyWit+03UiPaWuoYkmWzrbu4HX6
cLa6dkYPL1tqnJ11ODv8LEFmKtukYCVsx60nodVadxOfDHTizB+iz1eG5Ja0iH+uEbMi/+gh6bXo
wqYyijdfajGoTYgxkuhH3pDGxeiut16GtD3kj6f5ixpiQGg3f9jYzQ7FqAL5U4d/gXWMiFZbzz+C
SJXZjJjyduUY1HHFeX0+f9pjLaCGsEg2Ov+7zdpVg5PsbAYdQrvte7Dwijpx5ZKZ9J/J6TGPuC+8
og/DTYgwLpD2EhD4Frlz4fPxikJ6ApLRWGFPFXcNcVvmfpJuqD4lpKVbHT5k/QzvYEuYQiHEl5FY
PUSLdPY7p/sl+oMKiRNQxxCF38evd67/KQTd/3L5blZyLlInZ4QN+sJuQzxP/5+b8Krin73kt5GO
G/RVmRzW7q6bBqD0TQ3rI7WJbgYxFpSdFwcq9EBmsqv25ANX38vZX4WA2UFuyM4MTvole4RTsRNL
gObkcOc4kLUQn2XmESZa2fxMyR/xLxI4pnY6CJYAExVFoot6tcRR5xqS4f0gLfrrr4nrSJjFUIeE
0v5rpXIoiI2HV9Dq2vzhMbHjsk47or7OogyhC1OvrPQvCYz0Q7ku6R2lT14ZeOHJ/Dc7QW7IQu4c
AMYQEl4uigY4JSzmRtY6H2mN/KpELdH5w1t0RuWasRWYFA6SqX/85jfrS1Y3dBAxspYjULV/c097
L2JqImf+Gq9uiZhj4GbCTwYc0rrcomgO/juAEXxlnEdU1kkA2irMDk1cn7vJxVg2RbLpHrXy71Wt
ITedRQYc2oLw5cO/EJgob2wpBKe/5Z7qbxSvI6tzk21RJ3raUTEPOyZdy+/eD9S7BishjC8TSb2L
xw41BnjMLDh0tD3wy8g2O5vNuWyUOz5H7634oEPjhKfdQlx4VOgkLcc730lKWaPusTbZeMbrShCi
l68LV7LtJIVbkrEpd/QS0O+m6Y+oWpVsW3Y50cSt5uEkn62IYyrLMQH7Y6W7+ELmugAJEvaX7XwJ
6qOQC4pmYspkKGaBXMFi/r6GWzhQocq+SWOWhGRzTUHzIdVPGfzDhjcUU+QVNz0lXxbhWPX5ebMc
QDWdjnopQQIUhUfLyQnip86AbAq43p4FeUzrKej7TGayi10kMcg80+dpK58sTIBNskesoqAmQqNr
2Cx87d11VZw48bz7bppUoDa8mcmWg31kFmII9fhaCWTKC5cQKEXzSSedfqloBRSFARPiEIH2Yyy1
gj5A/c811EqwaZpwaNTNhPqU/9zk6IaO+VWrzk789OaFMuZn7dOSGDvRmAk+0u1mqH/6/tFLt39B
sbBoLyk/h3PF7s0cz3+Go0SItKBRc6VVopyliTb2wrlsdWBCWDwT9lBEwCVJK5OVSA8707igHJvx
`protect end_protected
