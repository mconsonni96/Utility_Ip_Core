`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
btP9Sl8oS1xbfT4xAQ9NlU0c9lAKqU4g0IY+Rcqc9FDxum39E4qFAY4QN7hyDzN9QgJIlz7BAoyH
lOYhnymEc28emk9se6d979VYkzQ5uwoCxm+iVNBSsvh2wTQYLsnUcMfIVfTKXGB1f0C6gJuaOM72
cdfExAG/k+2/OQjLXnjGg6c1x0CAMhCyhf8327JVV8jkWqT8f0AAgnzliLAux0QwGRrAFbxR03/N
wtYMj4FshB7joqZZRRGb/gni5XucpnXqzJyWrsJhjfjkfpIncGao5aN/J/qZUpHKdT+9v0Akxdkd
/plMQ4U/gjC1At9bjyb29Xvx421LptoLWHg9+A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="y49Lfj4r7cwmGLv1+st+xuGotvdA1b/oGiZBF0GYgLc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62432)
`protect data_block
3nEZzdWN2XmUmEvFHwa0szSzDYK5xp5nj28222DFwRdvuAe8d2Cau9JWgMdkFOZJ16is7PPsZ9FQ
zlvoLrLJrquH4+ExW87p8q+HvsL9z+dSUooPTTbQsssQ2h7Bg3CDJHp1WEgz1sVcuBBIek4Zfjdw
PezEgKISB2xpxuiqdLz5cpzSM3lNt+y1hcQvRwasHm8vME/SNySWt4W2D9XikjNxTc2BCl40Rcq7
0F4J5s71HhPZII+NxknCRMkZePrt6z436qqrDmm0YcqLi1WYRPHj/HdJ/mDYK18DaNC3IZEIORNc
xtgnzh0jP07FOpQR29Pczomqt68cyukr6lEDKk/Q9qNJ9ALeo2ZjYu4wFYNKmyurCNA5r7Z49Bjr
sKVWUTl6bX0W5NnxAjUQsWH+a4GFCEd+V1ZhV6CaIDySGfs/eRyhHdOcpuF66C63JvEzG1OZ7QN9
TyRW84BjGLp2fQnyBqpkh+Wrl8SvMzjgevFlK1bGOUDEx1IlKckzTKOIvtj/z6jWTiBzGnXOcgVC
wjXws4mRTAINOPxzo4HqPb1lzT7wAdKe5gOhkg9WVr4jrPb43U0TSG+Gy2oS6v5K/oQRdtkk4f2o
phjACWjGnDRMVt8TKVS4qUplLPFW2B3xwhYafU36782pw+Z1gtiF1SXW5vy47V8JVsMsASvTIMQ2
4tNDabYPFnOEnWfSH5qWK4Gz3FrK2FwCJsgumGOINSxg54JmRqfJSb+Bz36zYfndiU1xcopm9r7I
VPh+U6BIfeO5TMKbHXjuKdK4Kuu+dbF5BUzBw1xBuN7cg6X6ZEcjVJra7sL8lMiJG693zq08yHRK
edCR07kZS88dXJm46n/DwuH3ayXxW9CfV/gHNblGjODboVfjpTT5k0MwmXphgw1F7cG7sQXG9HYy
frSFfYHyI6QfzEJclOVN2QgMy5kmoD5Qbw9tX/Rtqia7TO0JBFd1SUba3LVsR0mM3tx+MQ3xFxGE
x5T7kSK/WKBTpKfpBR1u1NJBDEvcH0GVHXnALR587mx/Y1Jg3XUXS6suulmoIF2TIXP8NsW/5yUk
l00toPtpeWi2Q8DpzHEQFljxItoXovSr3SRBpx85GupapA5MXqh83TfmL9B6UyIgAAoumLT1XlHt
PSxVaCQSn0qJQs5ZvakWMKOtZIWqMIFhauXkkbBTLyQVs8mbVJppYFGSIc/VflQxjY3dBfdtcr+o
fkAiVh1tsaZsb2yeeLfUQIIGqoH1TKjqNSt1Xx35HAAri40/AtD2CPnTasAOD+UUAHiGTm1EHVHP
6JHrr/gP4L972OiOCmdtVgh+9J0r1h8uGUST8mS2G/1ox/uARe8D9TcoWCLdlzZEybvNyIHisVoX
Xnl6Ai76m19ICi+vUQjwkdPFYrY45FVLVFFQMWy8skinKv3uxEuKciuCVyDa1OQMvAQ3ZA1oAJwI
mhItjqtSVKcFdtopPdW4kXLaVP4NyTD3G6HcV/q5ndZPpl21H9OyeLDbEihelK13VxNl+MmpgIFn
Rn6q61JyyAdQVtkDWix5ReR7w5rfw/T2bbeeCEMBNE3xjkv6prfLz9IUs+eLtZd2XUYRtSulkVjk
RRLOD21Py7OnUX7Kazpq99Cn1wle2rF8jpkc8nElcxSNOaIwZjOZNJevYoF5JFCi99BVr5RVoSYB
aGefjM5sBAQV/lPLE4of7J7zovC9BMthl3SoWpe21atBWhvD6hvZOPP9/QjfRB2ngA5n3YUBPzhe
63Hm6zj39nmc1s1LqMsl1gJIeYaUG7v0Rec2aRC64nGDjmJ9gsYVNTWUkLk/n2cEgPeFWABX+6ky
2G1SrXrRznniAMMCzv++uCKklyeYRKSR4x68MJSW1tSUKo3jPsIGsPnlm+IekGHR6htX8se4IMu6
Kb/Ziw7TI8iR6HWzcbQlx5sBDu+ttvzlsR1JrtCuIcoJXrHl1K8jXg6rAS2nJH+Rw5qvJ0i4gLVS
QTiyz+3qmg8RAuMBbWlpinQfzDwB3zetSBBm11JBDsta4uUfbhrE0Qb39uZ3NSTcOp5pSdAgNNTi
ykecwYEGq7q4Is+gW/4A7ZxuZ6x2EQ8y48P2kyOI4zY/g5ah2gFAZTRXiJMPsMm19YqRfxUuv01B
9qx3KrVhChn2sJhK9Tr19fhfoopBsPPE7YRpNczi62UPWJapbGKHCKhBqNkyqmydl6U4wRjjQ4JY
p0NIz5WEWyDNvwSUo6gJyH/ZPnV/DZ13Z+xVEIDRNaPCoecQt2GpYJ5kwoS99GCGZPbbyM1kvjNM
oVIQxnUPaZQ/7lP/7LdOoSvnBvmxlXcNqxwlcM+Wc/agND+lfmAuhU3OhRdz6qF1gxJoUeuvddYM
2waFXv16t482nQ3uNB1xNvRhdCokXxQrWP6UVFl5w/u6CYPh255UZUEZiV9SFx2zJVhGjGigFJ3B
t6mtg2neiopzmE86EFI4+0zok6RJCwPbCSKw12FEQ9Ybmkg/UqhObZE8uWGWW5BXj8lrCyxG0HQg
leG+QcI25rRaRlyHenVwK7og4Ht8I9Ek8FY4fAlZjDLKRx+qRYc682QrBii8zG9WQiUVH7UqozQA
fTcnFsenqKzbvi927B6CAvxdgmQl2hP5X7667Pzu4dlQujKg3D6A332LEAov1YjAiwA5Cou4xsob
/6EDxNxREBzd/vJ2zsO4CfVESq7Ize3ngvpUsGvgbnHJT2iirmLOOeiGevnF2T3r9Vc3uKCOCIg/
Nmj7wvlTahgLw+uNK7XW9F7kulRgkwFwntApMaIenUzBMZJ9yCy9pfEGcNAd87V6+tWK3DVjVSI2
94DPIDqELYCV89NrdyOKWMK+hVs3psde5iWZFuM32BYsC0LFQY7hVo/XpGXoPeTUDXD420jBdGaS
JENNOJ9T7x9opa337BDjl6MDVTVUAmn/jlxpnzLfM5oSXSWZSKKxXJSHH1015q3Is/XbmsY19U3o
4BUE8VYRzoQ6qrl0YYuBEGJi5oOlzJMcoN5F3P1aWD1cFAhAKtXAU54a6ZiJZHDUhUBzLWZWmkHA
tqgVRwWV02wS56bJi7RsoEt6/cj+xprcrsOd+XGyaSc3OKEPAucNMjqvo0N58pEk6GOrulvrLVeF
7XKZGGxQaav1USlgMpS8WQa1Ww/ebpfy5OzltZbyHCNuSbOpMHul/J4LfOYU5UXc6XA3GXvunAgi
hoTYb52mjG/hMYMfSCxVuzlZXl+hd5qx9ZK7rWO4tQ4qPzoV3jwKEHz90FRbhSg7KZ5a4cJChBoh
eCgPNe2ynF/L3BJj94B7WA6w1OiQuT99XuSEhXXWGv2dh1Q6EnfPsOGKw+vNJMMRGWHlP89IPRNe
wOyotOs5SvJVtZO6Vt7bZsNj2as+fmeePSDOH5L5hEwskwM2i/+oy8N1ENzCmwbcH3u06CbkN6Nm
8mMXxPUXxRohME9Q+qbFvvC57wga9xrzvcAvcpk9bxSHhXLJwVfdJjKBLIkuERhj/7+gqvqJj1WH
u3i6ZxzzP+lzbtmN79kWRGJQQw5galdmTVuD4F5kMazwO81X5RB3yY/bwzQxewsM1aWqzMAuQISg
Bta74J/u1fGKdowFtqi/d5I7yCJWTwVeUlDUkucaFnA8TofU5PJp0YMr0QUVFRz0Py6zMEDKWVqZ
l1k3NtRnZVMdEbM0iJxyHy1XyBTPbKTUzRuQh3eqtbNIcvNpwsa4HgMGvf2790ov++chmFAHA4Ne
PhsR91grcmubmvPaT+WLuMcoI6o8CcfuHcQPlPTh4tZ0EX+o/J6wQ849qv4MomfOsHnor09mWEoV
Wf6hHuW61OuR9ERpLbfBhlMimsfOgVghZBSvSPz8R4KBukjpoQIVKWYmHPBzD2glPcJOXSH+RzJr
u6O5HVQRQxDJ8K9uHrmTSKubhdL2h8Xmz0NFT6bAPNjKuywDs4bsZ9pdFmAwL/CHeQbyn+7GxmSJ
PO1zgtq/9oekYaxDFGni+2E3zASSqEyBO2OgTffeSN/3DG9+GNOutTUDk1rNge5occVyGz0sAGGU
L+hoXCyQzzXeC+sDn3UkeWaQcIaEWhH4Of0oMr3/L+SjWacF5tKsb8w+JzLfJauxOxBll1Uo7ms7
Ia/RP2eFgPafl6sT9sAstlKr7r5YIy3XH2NlLvli9rYbmJ5YXdRrK4Z6Lh8LuHRnC8mnuPOYQKZ+
zMBwLKAzOpcc8gC7a2+1kYw26ReJ5M2jBlKAFZCFoHkw0ElOBurnD5UF1YKsB6cW+swe6c89Vip/
mdvDlMdukkCQPhimCLrnr6aH1FULU/aYPXO9CiJaufHLbrGiaNZn3sRdBd2w+kOSM/7RtzQrr+B8
rqPa6rMqQZi4QtrXNaDMaxPKhzt9i/Bv7k0pn2oxXnf+BSa5ja/L+ZXK+ENUvmHFKWAbkDqLyjov
DLVBT+g/461dlsCuTUHJCw71SAV73ZEwGHsR4KCm8ndfSMn8qqOuIiChicnN5UFHWCqsOF+BQyIS
/8rQUTQ53Gi1Bf2KQSTk6Qr9U81qIrfdg/U2vw0S9eg+3r/9fb5FSIv6sadHV3K7lzGYjIUpI97f
MfHvreM/YEdxqlS9KGUNkskPSv5E87l/CfeoK+eOa7cwHcLuDrb4jNdzBinB9GPBgTd45J/jDTAD
11qNjspF3dMXMThnpKmXPpib7PVIoHaiB4xpx1/mzCaJmGXM7pVPM+mHLDvivDjrH2oUMh9biyBY
2qOc8I8Q61megpXt51M5J/ELiHWBUYfX1XuAaptuFync/r2zvx9I/j9K2PUXXQi2BJ7J1PTaCMfD
tmDma3aOMSr2TPKDhnlHnk4vDUYjBl2G/ZwnGPcJwyP76n98ki5sDvmAZ1Ct/pXK/s29NOI86trj
8VdmenGQPZ9yFcMAur8nqOS+vNVoafvEqOzlVwp8FG2ZBETyyslA/yp0kg5G+WVC6qfdZdt2IpCc
mgkzpx6tOq7vUhtkbP6HZIsLoC2IA/IgcGrA42+KhNmhdG6Bz7Vt8k09KsN0oLUCXkYm+oFCrioF
3orBUrs4Vs4OAGBs8JNxPCUCp4VgkQMOg+niesQ7uQwuR+KUUI1+KAwWruKEas0URZCRTACrpJna
D9/NmEhEZpMzNnr9SbGApmdtWJXWhBLiPjAlQyN6pEqOj+0i/4P4ExGdIoRqJhoQp8Hc6QpmJf3c
ZwbOzJZu4xpIFU/IKKBB9QtwNDYqgUjd6ICuitV8aM7kMQj5mfOf1Czq5GlPpyJTTZxal3r7tuF1
vDu2jw6evU9AfuVaKfm//pPiUTTNtGy7fypJqp4h39qiW+oTewUr7aOP/tYVIOhFNVqDFaKJXS78
aksgESp6v94iVYvqIjFZc9Xj7c6nfEaKrMVxlSk1+TV/SXe4oyova5WQFrMaKe8Y0HR0ilkRnlxo
DME2Tm39vwTUOEsjXzu4vtFvyAymydK+T2Z68r+HI2SzitwD4zzE4BvERY6rGD1FnKPvuBvL6yqg
3DQH53JYnkdJLH56//g43GC8sJgsf35Cciin8ARNM2P+J/B/bO6kQHbmcKvyWfJLa4KtQy3IHah2
K5pzaEwVKyUHvURBYvn+zXQXpXzIua28iNRlhgexwt1YSHpo6KVA2LC2Wag6S4/ENQy2n1VLatin
PrHi64+zSOCko+6QDMWNCSPWOvqGqRjYlhzNiyeZYaAKzKZMzMlB9HKoO6V/L+8cO7ILjU7qMp/q
Qf24TNS02tcuxuemmuE8hi2ERDfejYCwxUh9krNGxYceiGI3LngZ1Vf7E5mgWPbl7KNBUu10idaa
N9H0d88z71WxzTjq83pipkJ96HhS2/7brlNlL1XYUlgW3jNDIXujK7hXysyKv8nzrvce7pZbmU4Y
hUIEPmp/TtdzLt2Xv1WvRUiMmFxSsWimodkvaZKCrMTYVosER8/Cfqh0495W9RSm9yrNWtOzm7hr
EQAB1KzQibSKQi5rFl4ggUREnuP8DwN8k6CQuDQg6OxEou9asIIO0Nmtk1RC0GjEi+MNKuNAB5IM
IjjoIkREkNUTkwYsL0BI5JQ8Z38dPDiB6fOEgVQCH0HjGt5AG6PYGxaWjnWjTVzO7K6KG/7wVYZl
RmsrVE6CxiUnf14+A9aAvVpo+y7DhiOyoL0z+Dsquvz1gUMrrO5nhzCZPStKavkm2ecpl1uTYnmj
IOSdmztqR1tyVzwDY+rpzrzYwgcghiopHYJP9me3TdnF99N9qY8kWGDUahOuOTVBTQumkwgph16w
ckn0LBR+QTZG/g+fnqQON+PcrbtpqItKdTw0M+VJu3y0TnMCL0u01cGeHAf/2ygUdYO99s4DoKA2
y/JSXx6fNUVRaXzxbRaVdK97AWfM0PP44DfPWZuYB0inct/2Yux/blKiBqhVQ5ouRZEr4KvlngeI
/lDVrXqXQWn6SnR+UgtfmIrfaaQ4izySKo9qYqe6Fmq68y9np/ibDH4Xg27ZmvtuG3PZkiK31P+L
RkoDTpg/jea3GNCba3jg1rOP2ZPuDrZATaO/1cmOIYBtETC73gutlvwq+R80qHrlOrNwgtSF0ry1
73SFI3ToumleDdU4OwcyvmxZaa3/GDBAmqTu6SWVB4VGDqk7P7f6lVnrlHiQoqQPIAHidWY4qVpL
IopkyjX1dSDClLy2Sp9TDPMtxy4tSK+EEORG5eIfbfdwrJO+Rejz82s4KEBLSimm+rgBM+hpir4j
NNhtepwIc8u6EbQtyuUyAROn0nb81vWmfNGkW1ptb+nJtF+E+HikTdn+14LzUZuhxFNgX89NhY9m
UhkQgP+DQNCWNYrPY/BnaSXqV/iscFEaf8Er8TJRaTPy2PS51jA6/txEyfgAdkbrDS3uJ4NixYOo
hVfliDF+ojQllvX3lbGXrWiutuHPdvD9QJ0w0GevTk41tnjhAvCmp7biuPJZ5w4t/ugJooKTqdoZ
2YnYpZVg1ElmsnZEnqs5n6wOXzSwDKoGZPsBbZBYv0GoAVy6RQMdT6ElPXtIzUee/umhbJQt8k5E
URbLyj3NGKtjt3Os2Af+K0Lp6+bkPDZpLo8ztTd3ZtfT5FVRRCSRqA8qhiw1sKFxmg1o6ya80Hnv
H2sxHEqcIJ0E8CTw4y4plDRjQb/pz4R/nLjI6VWIO5XP24U3b2x/g8viMCtdmIw2R/LmE3xQJKwg
ca14dMzGvvnq/ola1WXTefdrUx6PRKLk2vItdh3f4wAM4JpHazGl1y0LGyA8Su/sxl81xXZPkDDl
aBBS2Cj3HMllIWWEpxPYHGyjtMsElTHlGwQMwEZsNw3XioP2AUG9yoQskk7V5uA9NoxnolNkzT14
7waOouM8MMTArii+aj3BcaeAtifMH9HQ5qCsRhZVQBH6cQb56fhrfNXnJApnmiJ+YCdsI3rbT0md
BdZNAvD8ORxBNd+5IDCQBoDgCpFzNRdE927Y55f2KR86gc9WiS8yu//sD5WsIoIWvYEHMBxsbQ5l
xlRlrDpQfmJvvJLR/icRw8QtsOLdzi3iHFxph4hMfajco/XA0UH9RDuNPGG6bw/aPc66sLG8coyb
OhG1c/UjDyPfE7xWRPDVRwvnHqjN5UaROmQSofjzYtev0/BTjsBH1L5VBCkK2z+wuy+d+RfXl47E
2U1/xm/uO07Lm2OdxY5PTkpZ4eDhgs+XYOfAkzIfV6mJ7oHgsCyWs5QaxyuLiBvkYMvqXMovMYoq
ROkX8sASmFVjLTY6ogJwNYqqxj81rBIK/b4tuddG7sOKAw4awY7/rNwhjDzHhhtrWjUfi7EmlkNr
febs0d4nsAbTat00XqXMC8pidtstcKUGMUjkHzEz+7Oz0WBzY3oNFj4k5jlwVy/O6XMzKnLzw52Q
J/2HF2iXa8s3Qb226Qupr8NxNd1duR3fL5QrRJTi6DhKcwmfWbNuYBDR2W/c3HRYJNVNeaRC5vr+
f0rUs7UbAYHV+4cytOHD04ok65+2YR2I8gqh4QggJP8rHX9mb3bve8ltz7MWfn/q8DrGoRzi10i2
ayk4oPkDnzB0VsvXHLEORt2yNmQGjrzp6bekfTEcPE08owyvhmusLtGR4ThESKBtVUK1MvnLmXw8
sMMFShEAP8BpMgJ9sXTstWpUbrzfJMBZtEowabVyojgEvMtOeRSi3e0zQ/Vq2Eg0A1mLTTOMmV67
4138dzaVAl5PRjxd1AEO8ownDC2sR/J4kjNaWAi3JCa/hVHkpaUPclLg52AYfZKlpnz34zNi29BP
M5pqAvnoHaqYWYmE3aYfhU5jTXyQjMCIvmAeM/2EQXXSlWXfDH8s6iJuNkhspQ78C6pjp/wnz+Is
JS5gQWxmVs6h6CKKF+my2+OwB7N0yqi7gRIQd2Fg+sbL6gDHKLXW1F/uZy/LJlKGiTfLi4O7KZmc
yBrVrHqzT1U++PYDiU0fqeR9rq/BOMkIdto7DyorJus2AI+ocWn0nf87ozscx5IqUArDUpjteT4I
vmllj6CTb67kQEcQya4C9XuHY2QItOozmbHgYMjDLeRRcelv3W1sZssv9mpjviVGnY5wqoXVFWzH
JTS38zq330FjPHP+s1ikcDsc4tyvrvGZC7oMFRVjkUlPWMfWw5G6FH2A7tzFg9aQfbXHyO5fo2O1
XKHNuke36mJqAMIJZvKI93yY1+eAjPMm0YTlMorZL6RVZ8bFVbHVqcfFJW0HR9/DLzzPmJ8rU94D
/K4nGvXFnwZtxv7l4zmOnl5XPXiLHbSSjtGrxGnY0QMJKbGxEhVWkwtr1+KfB7spYSYcWPnaehDI
+BLu1u4YXg60Al93BTUMrGRSHOUbky2fEysJ+e1f7WkGjjRBbcslchi/YbgZ4ZBO5iNzF1CkSMv+
3EqfftWDPhoVOAkMt/0J/+U2rCdph9BCMB44l74R73uA3Cl2LoY423Pu3DWa9XUX9bU/Oo21IvsG
brBgO4jJkSoE4I2/wkUuIJqA8UPFQCCclEWVSi7zV0hBsMga9m21UPf/qPFhrD081z3fDX2c+T8W
qxPHpIP8CCHKnh7IZJ29Qm5Sbo+Su079pU8XSyrcZJ5cUsWrCOU1Oj+Dh4rdN3ROohjJ98wKRyWh
yyAx3rKPShqz7ib2AB1eQWarY3uTf9XpN8Bod5+kXjm7mvvcs8FRTE41J6EfChyrdNOIYQgTIfc+
w6VuWF0G4EmYgnfMsCdIQI5d/dR/7V9gB19LIV/v3tz/GSSwlJsl8JgdkXGt2UxU2Q18FKwBxdjA
95Af2wYzvjOQrBp+GU3gtg/qgnWVEb7tbyulaqHRWBACP3Q0L5UAQ6GUqNnV53dlBZksdbflYpJN
L4a5sGIFTJiz4EeFWaJB4LU7bz435Pm95+LRM9k9L62/xj8/w0NAKmp3KHa0un22lqcACbWU+NFz
FZJkRj+TxPf5hSfZGhUbk+W8ibW95dRk3w96GQeQTHgohpoJ+wOZird5H5JrJhn5KxfQffrAYjIQ
OY1JUBazqhhrmVRP3mX/jTXzwxCaLjai8kEc/a7ZQWrM3KjbvG8OevK+B3HSyOGBFaoUbXJ4LO6N
nJyKujq2rfJJO8qWTSJblD/NOBIMf8YXNOmZDy7LK+/VQnOmO0sn+Q5qmuefH7g0y9+MFE1Izsyq
piCwOE18pzs9NDk0ELlNayQp9QxfKM+kiWBNZ89adt7SmsqRfcDjRdH+7fGlwrDMR3fSep/+HOL0
+fk66Yg+G3/c5HVQfjsxmAKW6LrqCqCpXnGpC5/W2Fr+IZtTx7Ifz6cdITR36j3/dPwLFOk5v7Xw
G605J5ADU6JuZupeZHIFMWBwvkQuWVaBAqFRu+yFQx+XtkVtZfind326IH+ji60y/UP7NP9ZIC0r
vkhPOIoDV8ZOT7Z21N44o5KMkIPWsxZGL1jPjvupFvu6S2VseMFfTr72F2/b7VqFdjm33pPsP3Ij
Qcw/D8c39LImxNBQ6UhiAYwz1AoGLDjZhjZCXqWeFrESyxGU85tCzUKsXbUoUxAvEvPKbSz0aIxx
ssJ+4P1IqxLGGhQ/jLRXAjn40NO5cJ/KqmRN5pO4wClReB4EKSXbZQplwLj6RfaHyi/uP/MHvT7N
FQIPivOvHIXdr2xsKlsH3tHDmRtuLo6xdqrTPdD4rk5I53XorvU8lyHy6XsBri/y4XD97IzEThNS
rc16MJ+BmbxSHDy6Z5SBmZ5F3eKGgoxxHqpBkQgDdpYQu8/HErH2CqfuAYgVq1xy8Xy3CWYFsH1I
Oo92bHFj9EbJK0geX6rMvZw/bV6ryzMAKqJ7kHw61uEmcvcCmlmwkTJZaSwyUSREyDfOqFndKX0Z
1hsEQ+0LIxHwaJ2oMOhtg//PqRqKSUmll5YgW67f+A8Jq2Ce7kEmdR2vNilB8YIV+MnZ8ueOiw5Y
ZWi7/34aNi0U2soxSCl98sXAjRvo9YUm5dRkWG+Q8wNFJGXpGAP6KiLMvkREJLPqJvsSMc4QFWAL
wakNX2k8HNYptdCepMMIJdxrYEnswwU18PcbQvXscm+AIY4tu1dyKazWWpgWKkQ1t2MSUIzJfaLJ
+kZBTAWaCtXIcvsApjHS2U6fG6Q0CtpY2giQobt1wicEE+AvW8s/ENHdpprYLMuUDihqbNd0dTdc
vflngKc9SN7Z1ku+GqzyUbDEBnWtiAmxubxbruYEwtR/2azM173AEmv2BMjRBOyUeKHmlZm4o+xC
crrpBQ9b9O+DR6tjmk7gEumzeppifAhdhYK5k4q+neC/QxprWlL+q8dkpsT8r2emHmGaKD7HVmIM
4SLPzM3uA7nsmuPo40tC4aZksa+lX/z8HZ6j8TvvO9UaESDI78piCBkwDmIxBSVw+davLkGpwFpT
8LfKm8FVrPcWbtM35+Ls0E/Ef0EuIFsRst77GZUb0Ry0O/PLrtL12WGNUIhFo6j39DoRlqQ1uBJ/
wBPNpsSDvdyKnbb2VJHd1HG6onC4FxzhDyny3HVVN/+yuy4wnYmzxzXg5ie1i05fbg0gsTid6hj1
E+9nJlTJPQWgN1S3RESMx5EINsI+ipmzFIlljmRyFXEblQbLbArJPDegwbk5SRSoLWCPlaOWCeX6
8pgkYfjS/SdraK0ngPtSxoh/yi9sw0/nqMrHvpdPBkFCsfxJsY1FWJA33oHeerM3W5zGPvpNPKnG
oPSoIvcKh+69dlWIQFz1ViaB+auyxTErLy0svgqFaNwnPLjOVm7fYIO/74x+sAF01VHxC1LkJ6/T
1EylpM33CJaq9Q+SMmc5G2duc+onWj+h86wjXNlsPWE0rnR7p+KFhyw0x3v0F4729Z7avJaL6IYR
Lq9vRMFiTXbrjRuFa2Ywuco0oVUjd5sZ2HgHUs72dqhG1ewCXFuWLwNItJwFSg4OpQ7v+vFlD/Ew
PUJGyS21+MPOiELpbTfQzpyvNaOkdkqgswI3EwNm8KNMI2652T0TfUDJPchnAcTL0L1XyInwPmrP
28n+IP1g5LIdwiSe+NgzP01w2Jl9xxthTmMaQ447dFjaLwlw4PpRj3OUfGgNn2/1bcFY0J1V5Wj7
62u4p4vz2E2Ay7e4k05o7M4ImvSL+ULA7xH7wpqPqXoCgkqH+w53KlszqPVY1Va2YzUkCQkXepbO
0T7dCSHwpDs93zoxJ3+THzRRYzTsnWDXAXBBYHCPCZnFcWYz5GdU826KUQcHUZS46VG9Utblbka1
VSRupVUsJNpSqJJK8dWGNwYELdGPXRLKFadt3rbs5z6bMMtVk8TpkxCt/EwRfEE6JEgFtQSKmdrI
tBjnmxcs6h9GsKypzjONOHdgQ2VgW9qZ9uFD/ylm/E6V7MCFWb94m3EkwzFuyRUkB0tuJ4AZn3ZG
h/EfrbP/nc7g7xL/db9/BIvghboam9uxxMBTT1YlSZTN8+m95aNtlZXYt97hCTD8Duq6P+p1mawK
fv0F+COyqyOUB9oDiyq7CY03YZ9IBfe5VuEgqD1hGSIdSY2lV58iFpNWV0R2TD5tD6R0nKLlzLp/
tN0hMDuGTQpuhWH3sYXIFnGEtWBhBbkoE6Gt5G+/ngLd7YdOpiQVzUElIzuVmBHINgtCzkO8Ue/9
ROBGgsrN7hDY0EMx2O1ic6qgCir31hKjwDdPbnHCZa53J1vb0A5hJi2PJ0DmqlZ/Uu/LnoVVusyG
iLubhFhINPiujEIVBtbA/AxeC25e+nWADEHab9L7Pw6C7mxbGKh6QBRH7/VRPCgKOkSDtNF0kDoV
W7RIfSqBsS3/UqdP3P8ck/+u2ZqcMB6UK5G5z4ZUYn2nYL6ZZ3/PTYRGPh3OWmci/PV//QquQHcy
6QM100TCJAltDFB58JBZNI6hbAJ3gxpw62VXEANDJCbpqod+J00BQSu8sTVlRn/g9CbSdiYdd1yx
/WWEgDhC4zohKEoMmGJxqzWIBXpvXcQaDYdYQq6fIIR+YXTb+AQtDWFg/FvCQUJIQMOtXNYSp5dS
0JvARanY5O/1RrMW3TPDjVvlkv41+iQKkT0DK3pygqmnm8Nag4YatTWPTRx0nX9ow29oJKhmLEhY
XF4Qj2VGDUvluZDsV6Wjy6pL+zv6s1By7ZwIUjG0GuYMUMI/qMtRpLt/c0WdkTbF2yhOMTp/AqOd
WZvdJUyqabhIuUf3p+/veAPVbz2toUW373ESSDHolTzrKShD5hFb1VWIhylpWg1uqCzd+7yyKX6H
X27jR45tdFuYFDR3D1gT3SbzfIPDGSQm9NO6cfc+Su5IezgTgd/8ox/fSg8aOjBwvOoJLzNlRmyK
WCEoX404ZPUJSTDC+mGQuJxlkIr5SA4jqshVA1yZ8FH3A5V9wku++Rr3m1BvfGtej1zXykRBcL5x
csz8hoq4LcEeSs8uucQoawTQTGZ7VD4FhxHuJ5yQ9Gqi8dbfGCbBEJD2PEKGsTK+xiNnOXZGx/fz
fcjTVD4XRJGpWjJBxyZhk1MYV6xoYUOYSr/PmwEphq0wab3Jl7y1u+6aho5hQ3SPf9u9OSvKObvR
32UNPWbthyboD5ZI0IaHb646NildkcXPVcEhXYR/LbuQE15KEpzCFvXtEFRBx9SOF5SPey629+31
gJ8FUq21oPpFI57qaPpPLOEwdQ04dnT4d+F7V/BC5adNrxPiij8X4zGTw+9BfixIuN+xzNhYbvAY
dfQ8qPhXPznSADdBwgz4mKn6UP0yX0UO/E3tBbAt3TPYrLYYIyUCKohx10YAVg9MWAQJSdHTcuep
mLMn4HkpZr5kwvQ5GBWwHZlOl0YQ9BvDwYO1QQ/k2vPkOHVCtkpunUPOxUTb77rCY0TjFMVAZ0CN
4pfte/WfCGNIDDlGtIKqhC7V/tuvM3qFvjHvnmUqtd1DeFcbFFJ4LWBEZ9WUB4n4tnhnTU61VbXH
5Vype05HwQcROr4WCtVDFsmfBySEQXmjHYU9CMPi17hW3f3b4Uwk2KsOaxba3a7WQpPlByIUOwGU
JnRId0fggNBn5lgPAPuvsmK96334Cfx720JU3Sns05hE3FEzXSvJVgRndggQaHusnIwWnayPoS6c
EL52SfYI9qJTXNh2UU+fZ2Q8XcUhHBl31Xff3aENFQjynmUfeFTSCclUJ9U1tCxLVPeqXGx2aQLz
fWDHP2EXGKHwbR56zP5aeGKzscv4vrZiesv9nsBcAUeXh0G2lVa+cZhGsmFKFjo3BPdnZaz3qSxo
fsa3ZUEqjP1bDq5KdelRAnIVkJtWbm+gooBxNIiEmrYbwokmIPxT8QffOQsRqVLx8gRV9Re0zwxk
OsxMzHvBGqA66JsMF/PYCC9DNOFtoN6aeJfIjgp+Z8pXm+MNho//vvpsjmN+0XR1Qai/smJQN3oi
Fee02WDV7+e0BpLGM16e6Xc4HIaH0Hvyl700uq+ZkRmVZXNZqylsr8/5qsDHXAZLf1V16NHtYXMg
xK5NEihzyaXJHF7/MzGrSZWQ+RBkNA1/2MvcwrbshaGbNYmo4aLoVrtkSPpg0Ex5oenq2i51ihPI
r/0fdYa60/JiwbFDhAOgPndQOQbGHJj/rrDLFgdQfWFyHe9lyZVz56KFc/J32yk67zEob42HvhJH
fS2zkTQbatFPuxM4dy0agDU6wi7JXt9BajndXMxEp4h0OQ+qJ0HZ+AHdVKETBR4K1rolZvVlnSij
FAqQTqLshYKmXIXyADSLxXN7q75DrsHaZls0QKVI+T07RZ+NCsugMySbAcQ/NYDHH4PFnX41j41e
bdwLsUyOPwuQsiaasvmdBm7kZmbfJ11M5+tFRAy5NLyfiSID4vqnlfchcFxCAWeayRF6DvJrL3pj
t27NNGxt6nCKWXv9ojuqpIbNZn6Iag9H4574qELjoW5yUfGUL4tMDGyfxf286Y1n1JCzMceSt5Sy
1xorCC9sxYq613VDoTpFJEPZNev4l+lPH9VtPgbUvXv59sbCT0ux6aFIUq8rvTvEbsiEuqQ0OJv0
p6AMUxSMy5v0vt8YefwYmO2HX0jxFJdy6i28Yy6JkokCzA9ccGVYQh3QFhQsvZ/7MApAsQj2i+Mi
uNVDh/rfEwI8JIoLTprirgjHfLXFnRXeiPK1U2Ar3HYWnEAesLzWeZEjSILtq8oQgRkYnRrMxvNv
YW22jeVD5HXt3tbqMCATRdvzq6NQU7i/Cyx7bXyS4pbdwIXrmKtm91bpZULu3cQ1k7YcHxEELxt1
Z4gg90eD3wHrHbiJg5xF8VSCs84k421WB2ESMUIBdn3uHoQ6S5mLhRC+X45AqzS1lKOL4lCR+wD2
wbarwIc+GydM9VsjLo3CPj1uR8+f7zdW/WuERmFN1EElwQTSlYs1dKpeh301enI58H+Qyc7ua14+
bC2Vd3/EK/VSqKSy4L6ikTLEF3eRN7j82WyUkuHIeygANXc+9BjpokS2jMB5hf40QyfPUgxgd3bK
64smSNeJUOYmqXrSVxoGTLXHlwgVMgQ0sptIW3FQj9OaivMJgUGP7otJxD2s8eitwyIvM1XB0x/W
5Cnaoe13H9q9+Z14EmUMzzEKMrhOMWgZC5Fn6+6W4/J3Dfmg8U58dMsrbdp6qy6NVWWsUDlqsY2N
DaWaqtDwtl5fbRj7tT80GbD5+sawvXrY39oLoYnEbls98Aei18rth1omXa6vPU0XUx359ShjFXU0
FgAjuxoTky74NSqQOgDHkCAmKxQw3j5poAjd4cKL2PG2cBWw5lAMGcW7EoDXLjtcVMotrR3ebVJY
Cica3uf4x3n9hSOeOvPyz8peGd1L1RvbcXNn+NngDmeGNiIgPL7osddkn0oO/hFynDccChS71lvA
dO2Ytmrw7sj4ou37qtwqVFWf9w9t8q4DIcEGRFNvMcB51Kv8zP23lUl4MWTR7p0BbkZoT1MYBTA7
b9RLBSVf43itYrZfdvvDBb4bSU8wdtVU9p3ciqWVyLMV8wnvRK66Og9wHGUzJpVdUDDEVYDt7i7z
fynoLo59QZIr3g7VX9rdKOWq2eQy4/K4mQfs5oj7SHImEgcHWZ3mFTURWgJxAMbhsc7ek8uUuTFQ
Hg/qRanU5gLNzhzwGgvNfNzBRsg5MBpihUWqEpDUVQYlD9irV5U41zee8OmXwvVLFMBuE5PA9w9L
9S/OkHVpaOR1cgxUySYeToX12t27L4JLN4Na+4p8bJfBDEJuwnbw7+BL3EMDx6NUerUbWDheMYPU
wbcYFPJcHomRzqnTfZWAYBKzgC9uc3GP879tevpF2by7Ai8B2r5Afwykk/HyrxrulKbnkrRgPDv/
m2HUtbygXu1qMoOk1AqfpVGOb+5n1PTXIwRruzdAGNqzd/MctflGJBGPPpDgGlHSkvb5jXB8iFgp
RnbM6cWPV1aYFjtwYFwhriBjceFRF3GB+0GznWxVyMhyjkdWvzwb1GplDWzRSOvDwCdEalUrFV8B
Bsw43SaVE2QfcFH+y1f/XRyLABB37XGuQSX38jLivCVBXaJiBb4fbEfohqkn0XEmcAV9hDeXZE9k
VyrqkFdhdQbnSUTy6TJ2oGt4LV4F2g5FD3GkRw0RdgMrKFYanY/mTOfJYPWQr1wjQqcKe5z5Pzt9
JPq/dciO8LbNQZG4zD9DQyz6uMPq+palswoAfNL81k3Vnfuy4o5SC6tFtL226jvFz6wK1Sj0OYs/
WgmGYSc1iKr9OwckXP3LPc4C1SqAIemDlpJRnRmoCbkjM9ArX1eKvsIFnGbFA9yNGBI+iCYt0Pn2
12PwBnBEDOX6cWjXcoD5XyEEckK6OskzOilJU2SpDwcm6Vrb/YsoxOiKRZhrXPbxo6VlRVOsv9K9
8ZYfFHgZQav9rnthg6u+oafT9wZ/r4z9d4p02VIzYkArdy49QUdaPpwxQOKUQcWzlYyjlq4mraiY
WuA+z97r+SYnKAADSfni0+HEpBE/TKDk0Bi/0MYDYYvUYBFUKgGF1bMu50TZ/X35s956JQ5mDN2Y
V6fOX5GYDt5OHwQlqJcHrsaJt7RuRVxmDh3At8WPGRtIh88keu5IIBnQDOeLcxH/FQ73CNYMXSqw
DaaLGgxoV1Vje+EL6zPgid+IcuwBFkpZNqz3rAcTwbfRSjy0T2qe/9rVqJW368+mNkywMMm6zFqr
azLhLi5r7w50tzY2rU4XVLnxWibOVJASvgfbotLX9PRSizsvgcQ6vLgQPn2RAbpK1/u9Pq0hMlN+
EgGiixiLB5E5Sa/Ek9tQqXQ149TCX05qij816SKDVnPcRZeGHRYww5V8FHWAu6G7HjXVKJ79z+RF
0Ya57RMo8o9wXLiGkZkRexfuRmFXI+q/ryWr+4pPnoOgFHcgIZzddQHYksaKMLhr2WdIFieqX0hL
60CoGtPKSYrcDMlDQ8LXG5aq/BK0+bNRBIVuUpfH5nI5XBhlV9r4p/FfIVBG4gZwc+FjdDUDQq8G
iPz/rpLnt0bcr0cv0xWpo1Ps//1gF+NsMl0TXcWdGNTYdbSlb12lM7fx15WELwV3PbTPQ3cMGxUT
qwT6Gw/Dj700mfWJv0TJMtQ3EdsnTRy5lOebLx51S5i97yKZgBZ+yS9/s9mGa+nqI04IIX1mXPV4
cCnesIbia1GQfWdDPTsJK7tV79TD1/mQRf1n0LWHWkea90EBIGJom2/QoitCNXDdieokAIStG+K4
U1EF+7ShV8svukpgxbFxvYzOa1ZgOdk4bE3aezIuRVi5jn32Dfu1zdFPvriv1hDF3eslesBn82zr
hL3HqdBrCfs4sYCds0ENto0jMT0stZvQjdC+BnixxPoCdVdqLD3qr2xZrEL1E6hlLTlcz4qkxQ8z
CsxiYQ75yOQgdxXCPMniI5NBmcpO2hM3SlUDK39A4u7lbJAby9Dsp3nJjOEZp1j87rd61WrAST+Z
sIYZ/mpeooPb0l/+gurcS64g7nPk3OnaS/xRCF8TNVtnei2zAOO8gjNqc2LH54XbkpOCf4hU5Pde
lLoHB5WDSrNKVI1VIZKMSLulxn6KjsS7F6WUmHaR1+rzWXZ3HZmzpDeAIRwZT2aIvqcc1Wx0sOD8
RHFrj/d21CeacaBgQU2FZ7ZrXcor3ThSm+ivAg9VeE/Ml1fvKZrKoTPRx4bBxXcWwzYQ1ubyr5b0
Ixz/qQR/IFWixi8Ux2exC3CuGlyKRy8YZD61+mjLqnV/puX503m0huL59bcf/wrZd6nlXLBa/Ria
SGE2oTRpZY/oC529AWebDThWWUNUOIRVmTqznXMrjLjhNVaCuNN0XOhkbkjkCa44BX83fVm2admH
5zvmGtC6gMxcsUvAkH358JWmdlBbVd/euHWKdt8HA5o7D+/gQFZE3iPBhgO2Cm18WH9sPAwTeURR
eZx1QlwUz9IGYDetX+CWXu64Ou3veGMQHyM6JqnS96xVst5P93Gvlu2IMK51q4aeoMS8pfLpsUuv
GXXOC1c/DRuU9Zj9XV0aT7wdV6eTC+5fskZlcyfKg8HWRaH2wQ4vLWs+jQVyxYg4YxtCdaMWyB3a
/cX12J7cG5+1/Vwvg1aDaQHkzXtP/I8R2wwaLsI/jeui4aL5Mcn21MdeJ+KtTayIld70RiFuEL3M
6sQSGf9eMxPctVkcgXesPNy/NfoaaUJWUtBt3L0Is/YXbHyK3NExBKT/C+JGxMmKV0HEgB8SZQRz
60cund55ORRXfGRtzYmJA+KvoOYCo5VK4gZgfbmtLOr2S7IvXyZ9qpb6vSx0G1ZpOg0O1QoJ/wPI
GqC6jQwSQ7LWFPFvYLrMVJThYcxpRJRhNTZDBbP7Dpo2eoH1YOD/xzlyOE/TBld4UbWdID1hvaLP
gj6cDVTMAfAAnFuOMmJghDINE1xOF785viCsTReA7QZqlynhM+mhl2Hm0aJiAxUPcGQyBDizjdzh
ThQ1niyG4l+qZLgQxcAcW/FYV2bsmCsZlDJCG7N3AiGt/wV42kUDdMZND8axXKV7k+29p920Ap0/
VtW08CJQ09lZKObH7nrBaC/KaD4ZxGilv+Vy1r6KLpqElrNnXuo3IK0eStzB9HEjq/DGvNK7SNia
AwDRuvXJwImu0gbE7QEC0ZxTMBuXgu5+TNJMbOrQrX6ndGb4/PaQ9Rw2th0QtTCZR4ptRRoGbwXK
vXISGdjeYGCMVoTKeXMGX1ExuRarET/WrnwUryu7IW55DQq7EI+g2gs6TRbubv+Gdr/ouBFt4uJN
qJW9oDa5SCZjad7Kg7v7u+KAJpBvJxIN05GxfEJ/pLfPuUrAtfPqw04fMrzUBrcIUOASpDnatXI0
CBJdPt8KhLA4KC833q+rc2/8dlBRh34d0B3uahBuMxN3qYwLfU+VuIdo0SAREiOUVy8VKau9+svq
nsKKtB8uBsPpV0sgcmT5MiAfZYt7m6WZ5sVz19/D3ESbwf02nbEzZw3vpFo3xR2No5aC4OPvs0JE
lidrv4Sg8tWG158kuNlyj77/xUPqn8F8583k5K2mRKWaFwTL/sfKa3qAXw26WVf9Hgqfzz/9fpGf
SnRWKyk8NxrKEp1Q+Gfu2ENQEc3GumW7AMncvaZdShS8ElWS3M4oWfAIHeT/vTAFGCZZcdWrwCIQ
0hnT2Rov6wTcMJzJhIU4WJDUO0LHLCk5mvZTy98ZfHb57nsUrM5gSQtViLcAMu603DyAL+Xj/FLn
sbW0UesdTUyjW8veLryxUAz4p5MgULHI+j5TCR0QtCi2yKM1N32KbHoTEano+uoZQIg/NNwq4rTq
WTp0v/QNuRMYe2/tqWx5kXVhMh7lZq3MWyb3EFdz+daQock7Zdrf0J5Mjnz4VKHrLnyGti1KUjuC
cFxSHBPPRpJwcrIqnBIttjKAr7CEjjNRQRRf30rLrjs9hDuUWkI8BCYlJrkvlOXTdg8qCbv5unDs
yGYHmN0RDO0RxUKItT2WdpIRQy72Vcaf64qKF9pxqHCE69Xlk7BEK+Rx5w0kMelcSCzNEpX/PEZL
6BfvhlA89vOoKO4xO0pLZdMtPk93aoz6tBtf9Y4U7R6Nk+UzoUzZC+LNpuLK4sdSp2Ixf0zTI/7a
6G3qZ7rgmKSijg1UOlxOShmGFuHvSqPe92P0PIBPjfNc7nWjiNgd+y33zUrGDYDs8TYPosIDGk9s
0jghwUhPgt0/sGdUXyixhE5AMpwAxEZiUMf1VfGQGoYzlbLMaGza594xUd1CLbD6TTvgmHT/n7db
DAFTpUmMMRnlSdzus2GOHmwWyAAil+Kd2PmF+5JNM1s8S2XHmePlNAmI6QX11z8vpdhP6Y2Z9pcc
NWhrGbwdFfCinTf9zfywLD+PRr2FYjOIseOL/QOa0ytbmGwI7Gcb19r/I2mZZRuR3aBxsExAVlvJ
WxkXRxR0Xmy60m/qeL9CC8m3khukU1i2lPlsB4MIIO0JRIO6M0PFS6nbw1x9/yHP0cuxiC+1hAMU
LVQGcpsHVvvvFlI5KkBp8Fhi7L871RquLHKjZBpl4540hJJwDt/kG9d/2LoNlRP1juQ+8wiLkNfM
HS19SzsiEp11ZoeZ5cH2GXi3LIBLABHGlPHGyBsCuEHHtnNnwutxEUhgNFLw7e+wMrIS+4fqHeXc
8l0sTOhDWdyB4qA2ylIMfU1aSDCvVChUj6Bkxc+8W9+GV2tg9/JIjrVld20bSCglfalTtQh8c3jQ
Dz3pS24ohx7yAB1SMhu4N6MwdiXGW7Nf596Wxh8TsIqsy8zdNiD0qiZRmUMg2/UgjuQ3Ke2l1tBu
MhFVT+UWiHzMPPuq29tMa01sjsUSckGCNV+ggO5KF2KuHs+9cA32x7yqfu5iQKOk1RQq6sxGcAij
foxsOfcjwyqeWyug694i8k25zzwBwkgKtxYTMn6skIC1Q+Yoe/mTByqwhiviGWrtD3oCw8yr2Hp6
35siSPL9VfiEAcDnaQ1uJdT8LDNnCRykWYabhGEiitVtuthJ5HcnfU/U5xmJPx8qP8lTpVbYHTsP
Quf5TU+xSdEwMlqNjOJE8NADYWQSMrTpD3/eIPudGVq2lKvjfWuew/mK+7QomVBrc9HUS6vhOOTi
CpLG+lh08xiX+vX1gd70JZgAUH9VCzD68xz1mGut5hoZMQOA8jaIO74TaAyMuwJtn5bhgtvnp/4q
/EEwbwi6dUfiGBbiJcJdzyAyy8pmQiHReT5tK8KnxBGGws7Dyon1244pjJpSQokl8o9Hv7ec++zg
ZfWgTaMEgsQIuhIYw6QHvNBezP+KhnyieTZRR/plOy8YLDt0uwsxyCeV40rZj2YASTfnGo6wCUW6
tXkYnLAj9L28HatGJe1pssrYSPXsPIsfIdTr1ttYzLWgAbOvLOtA5KTW4GZKcI+3G4nYQ5xRp3je
qtf/2UWbVK92wnIXp83QcSuc7hCC5aWA4etxDuWGot5DehIuaFaC3Hcstmqtb2KQxPK0aYj3I50M
UV6Nfz+hzgg4k++oY1hNlgbFqJZu0++cR0RAhXk7fBDb3naC+5GXGEBTvr2n/14IJHpoVCorozLJ
GzI81nxMj0ducMuw0csqjVAFjVZ4bux7CrvFqRRBVemb1aPa5zi1JwHtkcNkB3qRcY6DpY6KdVpN
NqcwKc45/s0007+NgDdaapb+00cSOEj1P+uEAly//NYrkKAzcHXFFHmAB+QiTYpjXzBMQhyqYhK2
zAr9PuaIOGooBRyp9kFNVwJYxh5/Kz5OIDpwkh8pCzotVP8LxWbBAFYosMNDKd49SqXMwPSPRqLj
w4eugam12UNO3xH4VETtLJ9DyESH7Etn/7UnC7ndDh8gZsncU86FFm6CXqnZkDQHfeJv4i46cq54
i3OJcVkZxZ+nLWkIa6xSXDDeAs9VwkhR8JieF2XoSY0wIRd6ITsb7RPI97vL75Lyqbggy7g8dKXl
yzHR3BmTRsu1HUXJzQpc8VOs3N3g2VmWstoQ9Qtv4XRBHtEy9uRgaOeTHEZDef7+noz4li+OBCrG
bYFWJg1j7AYjKqj/lrNUKWapS+2644fVrMU3/j92yfGtlm8GDwxIElL6kVVUPckdL8Ye8XPO6Kqo
W0Kp5kxd38oDEkY+gk1TkEdvsO+aMMgN9ZaKQlzofN8dCfl2dDRQteBrG+nPKrffvfvkbjtYSbUt
3mzJK9pt7ZPePUyzt7HAtS76F73VAkKpTNO656CFG6PLBk9VYBBPPj385+PqvYWZLA1aLmr1gmSe
uHe83Ji54J1bXNA0z6W1SsYAWNTPxcIIgnkDYWnsg/Dvzx82lFDVYUNikYVIP9TOFaWB9fAnsgeC
Mkr5MN5OZJff8Pz3CU4ougQKyK+zuY21fvVOC3gARp7+0lfNedqWt7DHDALGMRtrfCZ/ii8ngBPl
OSCZg3MsdIJN0g3uxUSrWkxpdFIpoNxWjrY/PcYhASVt0xdaejZKqkptS1LeaKc8TBtf8K8c6WXx
X8thkMRpI/RocoQCMXZ40Rm0cTKamQQujv+QKA0NdxwBHPjERTWUBhwTI/9gVO/oekFuup39pePf
UFX9E/8qhdQXXM4qbP0Eph06KhIcl66UnwudTNSTXRjoLlVdjb3sBpkMJW/TSqPCXnrck+9hARaG
RugvnSyPNN/Iktap+6gCAquCF1OCqZN/Td2+Xkx6lKSQyg6cQchu4lt7zsRwflbIoCxwRQ22nMTo
aAd4XFZhMxEzJbBzyeBwKLiM8ULwL4IIu1kov1v0BGmUDx7U6gyMaP7AOy9TjhW8XQH2J1G5k8wg
0gbWeLxhbHt7YxG0NJ8huA5sqYNX19dZxf2ZqgKopG/saRyFT6/j0FnQJ9PVrLpHsWM01N4bK3Ls
q8KCzM9IfZvTbAhEDbhBAXNnLNq4MJwPvnndNiGCbCROPl4xCqzfXykMDqKUdTy2stufhcjNQmSu
9PXbGPPfNnDpQFCvML11yZ4/CJBTIkAwoac0iZ2pGfQKOsScJjA2M7AoEkZqUIwI5YQ4LwrWUMst
6QjZxwGSz7NzdUvZMmCo8T62h9RG8ZrdrsBFTvBN0aFta8SFuceiS+g/iGifSSj3C6aCu7ihZNwJ
fvK5lqg6jERTvGuROSyQAq1geM+l2DaPYNCLSsCkXsNWWPZDLifutRiln6zrckYI0LeG4tlL/kac
pzbDFnak3Qbp/okiyWFOeVHnA+6nwgXCjRTw+eCF63J5hNQf1r+5SXdPK3kruw1U6X0kxqDOM9OG
pgBDWLagdAA928Jei4bF1+9FlZ85mDFzm4xAyEscHkgM5wKQYDlsEw6wDgQ5rS+xEDc5IyFPabDL
/jqgfqyCqIQSPjNlurUzXWAgS7TQ6ngh9p4vMIWXPFEx5GIWxvi+A0KnM8JvDvMIGXQ9Gg8/TEdD
Apt9QZfttBTEVqeZtM6UUzhqunpPxEPJegLUC3T2sS4hV8WWEiAxtg6kXNMBlQsO9fL4KTOGCWQm
p7zJ9lJYW2MJK1FGg03gi8HQ7ttlOLPzDMh0lbNrJ5YxFVZ1N6aFZIuGHXp9XjJYpjgppOKmAAef
rKHnnzTbXi1JLTq165EF1gF+gRNuGi9lfa7BLF4Ah8KYwL5zARR/nTxojK4Ta2c8w6IhGi0nGWIJ
5NkGXVxlP/ZNgVQlyEjBI9GVFdWqzg/7MvwC8yHt6GkYV7knrEHWQYOeFZpr5QHZHDtNob9qij1F
Zrj1OY8Uy5i1mHbu+iCJYGtF7kk+pdQIuYtnJsgkXRdmPkS/TGnVja2v8nRGtkI2pbCjflwXykTk
6A1FsJzVjaWiVdXbY91XKlQkcz73ye593dnWJCICkRJ+t/I9RxEcQGikFJewChRyQSkJd7EhXhQv
Mu/PHmflRC3R88ekEEIARCxQgRRK0eZpWbvNMx3zrPyL1t/uALII+VeAe5ZomjF8LtRZU2mz53Vt
QrRZraKqDDkz8ye7W8p2lo7VpCbbc/pIM9ox3B/mZDBPzPxW4VhyLNH7F9wHSBBC6iIrRdzR31cy
bp2UeYdmBEuaBltlpfMFVUOQCkBjjcfQ+xcois7kt+fipYEFlnKMfunIJT6CtdeI9F6YneD3IUrM
bWXSxBZ5EAWXCPhPi1/1Kfqu8ZQzQSuQ6XvqB6aAIAr6gZ0mDEailTvUSRPZ97rF3HQzaj2qlxnP
5Z1gQ2548QFddURR7cN+9nE3Ho6o3PHYXUY+Rs5TRe7HzEOS/cMBi+D5AasIASi0NcA6Lr/Bflj6
NHe54Wb+cmNwYpw78MflIS0hWRqe/X+47IzJV9MPJ9sDwci2bAszZGKWQXx9IKJ0JJ4SaspJxdMJ
AiwFUeRRV6VqlcRYrBMET2SpaEhjf3Tue9G+6b/LC0h0it0rhKhMFvZ+PVAzZ5Zgcn9X+V30V8jn
gwbJhe5jIp3CBSCGADuW4hdYSKglP03DkDgD0MwX+/JppSOn2n+OH7/zoz4uYeXDvMndMN6O4/2+
Age4DKhZ0O5a97nC7Bn9lrl1Y3NqB//zKJZTpQ9dVaeXzm2oeS6ID0vEIjaSWS9T2M6b+Q4twqeX
vZn+t4CIJVP2vqCSQF+IIlRcr2GCGzs4tPIFZIIN8MjrJu5o0iqRg74AZqBnywAw+bMC1FLTjnU1
autzjhLKYFgELfkdNlrUm6+rYs7EItlDF10viAtQrrmqC00L0Z6e53OUtVvcL8crhS3KT1oPYXgV
NaIA5+WjpjHNUUzYGmVmM3KGVtOnTtbRrVs3GuJ3dKqX70LGm9gUGJbj+w8wbdgFB+Jk3DNVf9qh
nAI23kTDwLyZgQA4bgsIJNKd2AadO5uHy6u0Ke05Ctzbq5aO3wX3rd4YufZqzdQXrEhbl4Mdjn/e
Y0LzZOcRvpGDB3id35L6GB87k+apsE5YeWrT2glefd9PKBsj501DZSjVgHMBtJSg9z0HW5x3VTOe
c8+XJW19uxTWzuDcA3TTDB7cj2+kdQt2Yvf9VpGnIAk1UjG5cCdfnI8ejFkyOTtQKo2OiIVmMJbo
NKJFXDl0K9TYp4inAfx15maCheoTovNyi7RPn8UYMNThsPEM0SE3CST491bwtTb1RXcxTOHPMXQ/
vncw7GkPBtsBo7s0MDwJfjRoLbo/jpKgTfEi8BH86sKeD3T7rh824HaRp6K1xCnE0/mxEEWAmg9d
TwzfgNM3M+X7+uBWYbHX39Wj2s1E9DofuD83hfJeKR+M+XFkwB6e/8EbO9spgCFF7ZCGhVTipN6w
RUxLasXGKCgLjwCX1JQiSvs4jAKMCXKrFRu5dMSqDicAIAOmFgkeSOyev/llzyBbYvKME8+PMJoE
QXZ4xTtKJXOHKijKsMOMk1x/jm6SVcGLPl73xbQv1zRMvWk9tYBmn1cSLuQ17dhMu1dhN/jFj6TU
Gm6oI3nUG9qOSjdWQ9lYbGiYIv4I4E7WD0zlGAgt0hq/7nrf6jsZpTzzn4DUHDDsEa2ygNg1UE9O
e+urFglojdb0iwgVUBVAxZg4DZkWpHVeWXha97Lfa1RbBt310GfbEVKDTfFedje3+Ou2vZcm0+gw
Gt1um0Zx7IzA3mLgUUZv+asnksVT3TO7zkbsIjImnsLj4oSULkoiUy+3D8Xk00ZM4jb+91d0Uscr
oOgkH6QtUYgw8qI90RxR+Z5Rz7l4XqJ2lCPM687RpzLxNyTajhel+Kt0tZ3C3UONB+qYdobkAeO8
Uye/zKxpy76r+CJPumIQa0Xv6iXO2FZ+2PyEO7jTnui77u+gz2B3zFumSQ/Yl+BZFVyXzn/SVCdE
7EhqfxZnsUJsNM93tnY/5YJ1Hpcwo9NPxQ8okdKcjF5xineS69cXsV+pKUYzsa276qKnIeQ0HOtf
FyGmJMj3xWbhiDzqIFTmL5OqK8znaDf/ZQpIslIFbuLNtry/D30VS1Yrq0dWyyxvoV32Kd/NK5uX
/RqSE93vYBx9KLU0pqRWxjlf6JGlaX6fjlnQ654qIahHOfuHO/k4difNtzq6CGNJA7vF+x/QXnGh
PVVhzTtUBuAfZtChJgJONSAQwZuB3XuzsOkg00UXSRUeCM3oA/WYLf8KC2uUMIL3NEb+XUJ+Qq3P
PPsg64AZzBgSw1XauaIzlUP1fBYPyEMSbRmAwK/SMKuzWpX655iere5dute5Wmf+RyIY1MmUlOCL
0SHxdK2jf/xh5wnI+kBLHIfIxQjH6FgGqoiuKdVwQj8Ez4cyuHJ1TgQgP/LM7UKMsJgywggYu55n
f9RqnuCvnRpU38Hj6xbV+50IkK93+TTivPsx7snr09ggmk+YFgeS0DfD29pnV03T0EdvZ6YodhLV
9b4ptStzgEv7aQVEEEZew+pUrz49WMNVblJFeE3XP9m4Y1A0W8+tChvV3kJB+BJmGx2BxBg9tJRT
Pr/iz6Hc3q/iDxaxFAHGapqMEwXh12iDpwl4MMysAM+GcojyujgyOS9EPCOxmczu62Kq3Hcwe9qF
TYKgz87gDMNLmX/OQwpdGNQUrOMGrVQTCfmx17S3Qa/nH96pxlKKNqvJcZ2oJ1bEhkCKcLW7qiZn
X1h7kDIQDhopLum6xvLmy6149qb0PzGArh7m/6QP7IPjAY7GpfpjHNaJ3KzESzIgMnViGjsJ1sx6
DQ1tjvYS2ugqSp7hHmzwBIWcgDMF3otAxKMpbzIIA3FZeBtVqaIU878btQ6MPqTo506gP0A9PKfL
V4ET2KKH1kEQreJysddrrhKyneX/MSFctbVWkwBtrVzLo+S9Ie90brICV3pcZE0F3DsSdATAAkVj
KemeqHqybSVRzlnpYMs7CWNomlasrwHlnaU4H1BUOrD2asFqIQmghs5xCRfIffJw297CvYYgirh0
0RzcnLWfn1F39BPMazwgWp4T2ATUKjt2PpbR8VSPu9N8vyGGuIx1JxF4FXbEA6qgSIPE9V2aKF+Z
uVGo+O/QVwA/C85ge9q+7CdTVDA9YJo3ilTmIvOFHQ16GqaAqqAaOZILv9UBrFB82wNpH9BEHfht
2WpngU7A1jf138f4Q3QC3MRM2iMERCMXewOe4NFyV7sZwmGlCUx/9+mlOce56YF6j+EJz2Qr9o8z
hAhIwvOy5t2CyRmgGZ0hO+p3rjNxMDQeStePbpNIN3YcmHpNbwKwg+FDWQm5GwtcWMSSHMTFVp4b
OwQxXJJXe7JeeCqWEB1cB/wDAHq5qTS/xbs3jKGPoEUmSs7/g8bFXaXk4/liJoUQDBnsMP97MvJV
745+OFa5p2uEvTuGCT76Tg9OCsplZeTf2nAf0Xu8atpGiITvDPNjyb1bpeEF8JaSkjhKAgH0F8Gn
6sXy9svoMd7gYP/0rcTcudtKaCuC3xoCCGxG8U0llAwlMGpFOMBxmBBR21SEFPZoECT1I3xMYrvs
tcDwCYdEp8Ww/igDmQRqJ5qn0QkQ409cBzZQM/Y5fVJB1PimAI/XpiVVL03aF6RALkapMVkvQ5gz
PJ4i1t740XYS9kUiKAsGB1MmEZ1uZQwvTAvEOyDJFGdaNTkHdk795pw4ZaJbpAmrAK/Rq6vI0xTY
8SyeFgaUd7WM7Lt03g2dlFIa67h99Zcm03KoLuwPzX+S4B5r/pnsQZ6f9dtpbo8NY1iGTxMPEXjd
aHO+wzDL43GI6PZqiy48Q6EEQtRpONxB5k5X+5WkdlH7b/xQkPOUjYlGoek+VpOCJWFeT1YRrlFl
/SXsbLm5j5/LRps5sYUgg7y0QdoaTHDJlEiSvAOaM+4xKLuOXcB4ErtbryZv3FC7atJajXW0Nz1G
A9xOADL4fE0lRpxOlxd2FAC4UYuO0M9OjTjzwXXlFiW0ZFyQd1+CLTXaGuIPiaG808TalHqy6vkN
BN3YLGwsSiPSoFl08yITp0zXVf7vFdZDaqDkAT4oshCGs6nNLtMcW/ex60fe2TBDuhTCpxq1/VJh
S+F2MNGc7jDfSBPZiDObtFOgld79lB+aG08wtDGCNSt8R8OfCxeQYYcSXYNXEgcI2gOaFgc9qsuj
jwp/7cc4p8UdzSL7y8qGoGy51NpDO56jI0qMCFhD3QBb/DLC3kfK4g80J+6/PCLK14FN1Je0vsSF
hFLArGerAdYVoXoxThoKqgDSHLds5C6eekSbtesMcc05L9yklY02GwpkOLgD6AbE9RUlI0JkUn10
NlOSM+xLe7cQBlW8KadUu5kan1IKyOCS9azN0DXh9aSIqR6UAmzDK1j+UAvv51IdwzE/vmfN2NGd
Y2FUXl5/6J371cWqsDdqbNe3MeUZPFVlaYlDISy56DzipvOSuDyFgDe3pFSUXeGPYJBWRrtUh/pf
2T/M5O8Pdc0HgFs+lMsGgyhM47m9oekQBTZNHujJMgcW1M47th4wCZoBZNJRFhTbA4Th2IW/tJUk
6LPzXBK3DksfkCNDMaE45cXaVL5e3G5MltLnweG3YNm0ByrQzROYV/hzH31Fo8VgJ5RchgwPeZea
9Fzay9DtaHYL13SPfNsBnDE1ykaPrWFVeKpfYmwBCrJZEdWBqjNNOApmFMfrnDlNAL9t66W2H6gy
dcLd2/g+XxD/4SCH6F59Lm7reYFlgTYM0EiUHUbHpLbfQa2CYp9KnE0ZQc4UWxTGzxsxq5h6YktS
wMeuoEuKRvdFPXTaAI5zuVBMe+5aDzpCw7Xr0M/gPtztWCR5iHVRKOWq69O074fBslC4TA0kdxOc
hQHnrk0DxwGRNgwJk71fUIzLlAD5FYJGK9VsmXOZZD7FDVzIsc7urZUgVmv/mTccCfuwEdsRNusk
PxwMZayWtUk8WqumBxTw0k9rpcqsGO/NthqXWRYWuKTrJmkC/biIaxHYTqP3TU2GOa6/MkBEFWL6
MhNsSzbSdl9dELHG9acW1bkx5u7Bj7N05E4LUZoDe4sVLi4wnNVPMQAGvpv4iqKPOfd2MDWssv5v
hrE07M64vuxtqCfCeMga3wVkWLgPlwlB7sZfQ8CUZkME3yWmPqBvqFHv3VFr2wvAB8tOGQgAie8z
e/0BbT9/lBs92TFdb9YaxjWNW1pkcDFkZmXmVhYHjbWZKY+BMtKhMgrj4mQXBUmh/nZRwDfUEIae
aOzGH7pGyo0PW0qfuz69iNUlQ206+kK2W8WlpPufJF8y+sEN1pbf4sKp2lUMZg4AHwU1SvcKdA3G
NSvuVCP9y5oLmNvaMbOWT6I2CCj4Vha+ypprP0yyG4//FwsDQEqx4thaUrZbtWPYb7acFetoYoB4
kIBU2t22VeI1YRx6eTph+eiDsGUCNHkyU8HpCo+HxL8ltx81lghCBGMtDEzwMBmV+NzKNHivpFMA
p5cPj161nnXcISRbOhzfNqwbhbPAw4KCxlFMzlu2JaAB0b9ZW8bindrTxGflCJMncy0LzedzeAte
my37Q0VYc6O3O5g6Gz6cob+bMxykOpSEwfzE6VczZNEwB2jP6J0Vix0gZZ0OvBFIhu8JXF6ZOeiZ
kXzvdNrL7yQiJoo62nVdsWqfszvZy7z/rWPWBeHFPpvvy0P+qojiHq/NRxHwzIlBxOL6Ql3EpPEx
gbU1ew0P5fXgI4ngmrNJkx68lN4Pk2mKYvRSsNqBGdMz3dBhiNPd5H27xyx3B3c9k4KU3pae/Az9
NnUulFQ6ZkA6oTV3rFV5oN0NVWfoFYDlCxcgh1ONcFPlswBKWl4Qk00XvPqWUIydnl+VTSuszY9y
Seq8o1sAzZH6rJ+9U3vjWbrgnWNTPYdcHOUXoaqhCGU/XCHAJ3LXHogc8XW/rQHFLeS1M5O7HN0K
36bPyqUGJjg0NxBDLmZr+JBHYJtYKAtRvwVlFNpWRwoHoQSL75tQGWkIP8qqyrlaWM19lZBMuXrm
NuVHHJh6ibpuJrDqqKuEvQr1FXXspwqvaMbiWEhIbViuQZQEprJ1IEbsL5REq/hQH7ji2ZA0NDqf
7jZP4lxhzDjIFq6hMHmCrieblqugS2Q+npxafxuhsMO7fZwV6GETl3HJkOtmsU4udNQlhJVYct6K
/9JKrF/2iAe146Xxistf3ZMKUnkKwDd2gbyeG/EPUFevuAuZYFqc2w8vgDJ5u/l9itLdx73ieI0e
AvkXFRD8cYqRdSbCa/k5O5VA1cTerk2JMBl24NX44Yn8lls57it8Wkz+PyImoqpFN+Qhdh8leYfc
Vvych6WJRrrkvZq8oz262ytBt0Gc8S73uheypsmE4DpHm4C6Z3DMDVab5uBZpr6H05yO/+mFC0Kl
ueyZtGcUaV4gO9KruJU+GMkZFVg/VYRJ406N8KvUkmkTKbKQPOhWCTPNpO86O7aFOeAwFKyGBVeU
HtSwiT+i93JQeoNigaeAf6pmARFZaejvXrVx0mbz4T3j5ZX39V15/DkoT5BfRyFmvG+dQxplodHp
AIUp53LjnzP9MW0f6rIZxF3GZ50jSK12x5EQ/DeEUBdGJdOvPAuohZDtcfGXmW4i02GQaY4cjHfY
mnPV4JbubsSRJuJoWaau8T6SX0LWvGVnf5FFDVSh0C4n9gsxwhMnOzZ3Kj6UpFNOlphEMdUF8got
UmBgrd62Zc6n8D7gjocqdc2DjKLWPgU+kxt92dQp6G20dovLW3NtGoDsb4H7sJUINvXWA5WWid0F
T1vsZORc9YgNXd6T3SxBeDFUOu0hOHS4vnM5KHQ0Ejga+s5TYxJlh8c3jeCxsxILcumUB0SwIYk3
lgt5n/hvrz1MPkhzfZAa44pn2R57ClMKiFuJPa3+NJsAdsPfOMyxKzqcpJ3y7Y4u7alGd7R9GjWy
qEBMYql0ekGGmCQ0TL4R4JBvZmZtUG2UzQw7x9iQAw7u16vAfZYE1h3dJgRMeo6U98DYiZH1nxxx
YC7/sTeCFHpl2D8xDr9hfHsotvVcYz94rZ580WRa+baAHXybLoz0/a7R7YmM3d/n6gC4v2OAOOWW
t7DEOF1vVVwyamKGcV4sk/4+EKV7NoOpCuKj6zV3e/yYBGlQakY2QbQu3wHmU3PIQHUxh2A92d0s
X1dRz1LdZvFa3XdqQh/+g6GgVvc8MBXm4skVSfCQOMEaDfDYkEpg4BAhCj+qvSpuaXQz93FMVIXa
JTTdGrhl/ypqlHSjE+KBUwUX/s/r3BHOLfEWLHF+RH2pemMtvujtzN5OB+orH3NlmCdXsbrVNTxK
a0xMO51j6JNw/iG4qS752EpZvpUmPqpdhbddnLlFHWrbJdC8DXgKtG0m4X+iyqbeDpZRvRs2AN2w
oaKdoaMkv+rqu4HoAgUU+tz2d48UwYtxaCicC9i9Pataw0ygrNF3kUaUv8vr3zPeD2rlH5ooZAYH
DpEXoLJ8DLCqSLzP0xSviLvyyiSAzgDvUk+ZOa096JquPzcDzgLvcPbO65MN/WsyA64m+RLykHX0
khf4qWnL6j8uFNQIhjid0K2anhG2BYgSj3av/C8R3uX9kUIy9SHLf9dvuKSwZijz/fUJnKugdHWf
h1Go4UsBEZbDD05kn4MScEY4Ml/PpHrwVOFtYRD5Y/V1ob5FXRAPB+fu+Yk/N308slBVi3LU+QWl
ThjBl7VVlAOOx7XjfYkbnp7U9oCywpH4qqSicbtUf5FHQdVm1WWPZfWCY31bCqM54LuchQJ3xjk0
ne9KRKerWWB2PyL1504/A3vyXmeFQJ2BywQvW4EctopjszlFVh8/pRQLv/H0HDV1ga2z3sOXD/FL
+IU6hKsfhtEZ2556ggiqTJ2SL67EMIPcT/7IhiDPCz5IMNOlLgTBxCtZYTrk+Tt51XGGKl0lgHtZ
bJEq8dCCM9MI2skSxJOFWgV5le4hsyDL1rf5YJbIaxqm5TOdM7bxfn8VracGbE/tuz3jgXyUVfXC
pw5vVjtdSBmO8f8FCzyZdm4zgvq/NG5ojVswWZT2ZNKx9tUXBDIPsGZtGIU2TKwRLbHJ5RZoJ0/9
smPdClhENF0pqnRoJ8fmFvlHDexmZJkaNNDmDsgg+vxKZhjHy6THOvbwr645Ezr8VBtrMZRB/y0m
xxd62h2W1Unf0Kab4zZShmUhQdjQeMRFggkVmxR+KKCskE/Jez/ig7ZezPIoV4ETTfTTzzqfxHxj
WNYtTrgSjRbObzKYOfqagKNDhv3Yw4jWAxY+kK3wTfLKdjPAY0joazFSWsXtvA7dNx9Juvh5Ca0o
5Ltt7TRm6CYJ1l09ATxoOTgWbsiIZ1ugw54/02N8XHO247JwMwP9CPgHuavqHGu7Jo4IekzmDoVJ
pwfYDKqYgkTBI59OjtteY5wLDTJiOK9MdaGBwmHJXwJM80JNfkD0tTOfqmbJPtxKGc6C8mjQOecA
Ml3cnQqVtda2upkyHoX+j3JI5jct0j6W+h/cUGQ7ACxzKI/jQ21KHR2VQpnioqDfKNMka9f24Bzd
464v52p5x/35HVudwKqPWbe1IrbPKTEHILkwFMV3tyXiulLd5nBrrDJZngOsdPKiELj7J+0n2Y+s
nGqkCr1F4e0OcjVkmD6EPv0BUU1h9Tjwgu9PcxuV/ghlAsFBUDIZ8l7fhI3PCyu0SJTQdeIhwmn8
TRp2QNwd6LTbtXV1ZvFSEje1XyNZuLyUAKdVhZl73gQlW6E7OqLaoutEeRLZvoz19hVMqTOEHm7e
Cq8scs1mz9CBO7PjlaEd0z0ZLNLoDWU2mzDI/zPYQXBBFMmKAwJ+LKAS7c2wE0CTN7tngBnUfato
vFNlRxY5/zd8cEWGem8qAyX3CkQma/AwR/bjmbNsKATYqT7G1cK1yMpyv6lqZJG7RbslsDlTlDp3
x58zr2m2kVIrsFjx9R68kRZMOE06VfBlh8BVLqOOsa6JNwt5ieWpPH+XzzjgTDjdGXuZYJKi3wMA
3zW5ZQWrIVWE1mf3Q3BQJQFg0prahJVwF24Nl2sOw8lBfMfcQSeux6CKGbUyWPIYvUTLJtPHwCyi
YZcIjfgjALFbNm/P9C3fALouEnugMug0fJMhMqd9hCv0Ec0EoT8XjYyy4ciHVQIpxJBUyxOHeYDp
vwoTzvAf/Ba/pjHX97d1GqwYUrw0QLQ8oSe+GLUXWB3Ot+qrKt5AyQ6p04BGULmCvJmyRI2CX/QF
Spf1CtvgHHgr5ypYcygO9me9oTZHi4FJu1IGZYVQC1sY61MljkkeQ5eWVpNCKPLLY+KBJ/HQY2lM
libgSR34TiqW4sOpQuEsophMPT84XIsntGRNGN48DvHG50xHCLsmx3kApugYdywJybnin8QhI15/
PKZVjvtIIQ16eIjgwwM6Z3Jj7AdMtFez8i7aisZXHmWfcnw7lLWDv2MafbTSqU5LIvXLjE8XA4E3
EN0OnMTavl7yu8r086Vlzvz7ytKU4YhUV5p0qRkRyK+W/hhGAwpsMC5Xsg0+3byw46uZgPOtWiGU
rChscxfzEgC5RbuZgCODRP5NXm9UMolDToBK/1AaIfJ71ohFQj3aTTC9mICBAEmlV3rTDWm88Ppy
HLwIGj9TXsOCwb0qHdrx0vIaXN6HQZ3TuFhdpypYznFrdoTyX0u9WrpM0Xyko3qQU/SaqcxKs6i9
vtsmNvg8RURUU/heK4H2PmNDgigvdXSJBsU2wH91h9Q/c/eey4AmDw+FHFyFO4rugZ3oc0e99Vsx
xFK37t9aKGV6Nf8/tgZ/bumru6qxELvBtHdzBp7LrqRypOvlVTP84BJMbUaAtWcCIwImppm5PU6O
+DgJxOGJLjujO2Axx+kfIqNMPxMGHfe/w5L9iS3ps2lhH39MBSEdMMqjCoNdM483FGNskuO0ww5C
iYuc90z+Ft9rMTEF1hqykJDJkpTzmhdJ/YxqUHC7UYjDDrAmIJK1wcfocHCZlvrP4DhpwennyzWl
0Fz9zglUDDFGyQX63IwQqD8ONtx9zAFAVnlI/7HM4M63cQ9+LUapycfm6KKVz2x8P49QA4J3l9xA
PFs3ihZFxdKRF/Qh5SV7UXTP4wst4qEZKIYISD222U8Ef9NnesQ1zhZMcXzXIsQGMmBDWcg/3WZb
VDI8gx7dK0Zd4ZZ8MPwZ+LD5pTt2AbLZwbcXhgq+BGtE/FH8Z+ngNV1VHssNpgT1u/9EQ4Yb1oHW
PYspwHjSxIqJNYAOrtu526Ki7FsVlz3ADI+HsF99mWR3fPjRpjJoPc2SRB7OgNu8j2Ek9FaxRP1k
jiaYNPXuC4I5958HduNCoMhsIfc4vTILNfxovwIqoxhwytaJgSrp2rqG1gmB9pcK3fIeFdJZgjfZ
2Y+jjoxM9S0hM/y2auHFslR6izxd24SJuAQHlbvcZrtjTlMubq8GA8AocgWY2KDLfydb2U/zhjow
1A3SMI6ibnenRENkd1cMK9ZahmN5jmWg+Q7BlOQsMFcqFEE9ErVALjX/G6PuwsAnEFib5YtWgWXO
UAGUhBa9hb+/OEl6mltXaH9p90N42iTwnQVjdqzr3KlzrwO/5mDX8YUM7uMuhNkg0Yf2d46Kggmr
PU86GWrGA/p83Xl5LD19DLFipn2bQ0py2fAnlpBDu/Mn511+sMFripd+++rLHKuFDwvi1IYWfh1w
q4njz3b2QNSlBwlFR/52r21vH42wgCB08Xv4LMUMk/Y+tGvMgYXcZT2ycKtXIWGz3iqEE92keKAt
wvUVBVxvHzcy7siqCYjKzgXZ6fBzeNemWhHPxAmo+kHiF59RIauv8g5JcOECv35f0DAPySb1M3EA
2AIWLYphw54ySKgdEbVQf/wwr8LbEGZzsgSw3JIexZBJZv87C0CbBqei20pgPbx9zSTTUboE6JJK
Ir6lzHYuSvH3IjW4VCYzq3Mw5SzgU9ajRZ5kffsOuuGyoXBeLMbOMVw4jCR42Ji29HUwKXZHdACu
NFICwtrdNuY7MVsrudEcxAEIHlq5DoO1oNUBIVYBswANblg0lf01jEd0tMaBCqKgw6krn2uXYd1I
/UGHubr474JRMQacuwsx3xiSCCxhQS2z1t7JyFIKesSwTzv5rJ65Bq5xzNEI1zrvO271LjLOafM3
vD6MQ5ahiURe3cb6k4ztRI+aclFCrqTMwMAKjV7aAolVhiXWcFRKje2P16JW8bSsSfPGcwBeUNrn
8Strk8dIlEXV1om0u+HNOsnTLsFp+cKfhsaveE1zaa+hyqdWJADBksBVoKQgUlhINJpqEbDl36yB
KCVytkAUazMa8QFSUygTZPDFwdfhe6WgBZysxwyvFJnyvq+4Athf2h/Rw74QP34DX2RLvs28HugG
hpyq+wbFzGX1Uog27PsW/4k80JO3Ca3nU/09s8gTAxz/oFPYNbbuIpXuAjVotp4/547dnv9W1wAY
s5xb66pDRD4mpeKW+zVo0d1olMq4hpde1ErXlkOeST2XdOfHleekokSR5ItBO7xXZ2oK0D+3kOlh
e49QULvGHPb8h7jz2aG6I4s32rv/GAT8RgkGQMA6lGBTZfFzN0AhRQ7WQawPPrqzzlRNZHjKAONi
jc5PfbyzzhEa7ij+l2ok7h5GZPw7O70KsSJE5GxwaTXl6JWyJ5UAfrH+CgCZ2Dla+9ymAY3W1cX0
RYZgSy/A5bnLoMo2DxeUCLnGU2Sny0QTcIqonuAPJI0372BZsK2GqyWrScKNmuqs2GtZ0NUdicFF
nyEnyT1rFnLG3pfelI0enKOTc3jMbh17Md4lWBaznKPXvHSCtZnIwv2TDOjCmSmCqEhjHc8C8gzP
MQFnAx+ts9waJ06UgqCBY0qL+qpTtcGQIx1pwaPCM0n6mTV/IyLJ3tDa4Dw4kPBRjxP9zm5Ffghz
B+JX40i8NFajAyOt0RsI8dAuzh4AFoLregTlXF94C9jD+pm19j+ShLal0DamoGkuMXBtOE7l+Mgo
kon7c4reqwMc6G41WaHbXFdC5uCYG2kUdM+gr5fnYyxf6hpJckGrDZlPeUkB1EOaxtm2K/LzMBAP
ljzptDScwlmwS5gAQPosZAclqOW6NUeSalFGsU+vIKXFZj1uOM0auUDWTHZSQBjcDfU7dje8VU23
Nvb/SpC6EXDXj8akQenfBt3iffqeJQLcOCe9cG73K9k8B6I2N8tXmeqWF032S8i0b3gVWzdvCP1v
6Vs43U5A6Fid0TE4X6JgpHNBx5eXFkRIXPjLirmPojOzvf/CgYF8gfaSPv/7EIVX+VleAaaulMa8
CnsEcRUFAQ/njVp0IY04Tc/uUsdJy4eMgASJ0c+M1h6Fx23IsxBuyB4DLFfz8CUeYwF3HuUjeEUC
3sPIPeTF8pKNT35bm8+BBv3lQ+/1zdVwQLbZPc2TbiF2GFMRzlea4Dp0JtTQd5k9vijmIwbwZO1L
qrrv89MMXojaAkAxolBpWW8MGjoFNc9moh2Ct9hDTSgpfgTmmFtXsvd4cK8vcIrQECTHx+d8T2vt
2+4qbV2ZddlWJezGhe9NVqidoKx/phN4EcOKDmiRJKHBxBVhinPBV2FGTME0ODekUyqUdknA8NEj
FWSczaxkjxM8RR7/xxGDniO1d96Hdv/WfECfESWPkoW88fGU/k1FdVEHkNIJx9349A8LY7hZhBHN
nAFBWXDhIgnV1eAHICxOpeq+QcgHm+gpLVoKzlgzjqkBznNfCLTe8f2vwuUTdYQK1jRqrHXcn5+q
kQdnr6dsVmx9FHP73jj6CcrEfbKQIxd2rAHm68lakmqn4703dMfBn25Rx/6paymQWniM1aGwYIyn
Gv8ECoOgIqBrh5j87xo9B9QdjtESds5lXNEj23YCYcfpbyS4AZtI4JTHNNC+BjMNWyWglk6jyCQm
h3zbXf32oj+nqS/nTE0TprCoiirjkOdjXyvDQg5smOVLfxyGp6yooOjZTvHu/m7fDx6z2ioBJif2
g2i/5q0VP17Wz1z7BVj0TLElvZDWsGTPA9ZqxdONfxieVMKHoDu/oRLdu9WJmgXVDmP93ow5oM33
F2vexV3gVjxTfSIyqw5rfvR3XVEBTfXP3fBiNgpWzpyIN4Uq3I+C5HgSLyquuX1sXpXIfgQ33hrA
9/fMBZCX6Z4dh23qo71LV7Boo2VPEJp0rwtvOu/JbHyiX8B0w4x8fFtAyFeGE4Wk6qBn4izCp3kg
Mw2bbPzIB680fJAg2rIMVldUeBJm+pISw2L+jJ3vne+7LezSxIdBJa3mBjmJsLDmWy35AGPS09hA
a0lZFU4w0QC4R8oO0GIOcVxidU+PtMFh5W0WqWk/sSIqVPpxesx36YQHnP6Q9H1EszEgpTOIvdwP
scHQtQkWmhqV0yErQXV3Qru7Kvtq5g6M4UZb8RaeNyjs207b5TegbPgSMC4o1bKHR/7AdMIwF7GA
ZJ+Nsd3d5E3W9L2RbueOuvxIf/bsEtONqtxHq5fS7bvuc5+P/AbcB7I/NV9ZmoVbWZE4xGl+sqN3
5A6jeinof0PNiq+v99QS9hR1+2CWzlw2ts5zHCaVhP6el9KU/hnRwAv+24uLlKxJySCtB9+aypNE
vDEqciudfl1ZDoBPIpCQb/dYSJodh7C6dEdseyoIOmwa7pKiBqvmEA5lQq2xmN8RctKNG+MYScKh
/L6Lf4HaUrN/qIis9DYSGL6u1+lCAfZXOoxvcDG+pkbYsSTiST4aLq37Fzlv0GIpou4xKzOQm9GC
L+yTM02Uj5L4CA0cy7WtPEKNG6wP6b3+7HuH3J8f6a4FgT2iC196k38szydIdYLaurr7UjWo93Xb
CUNv6S0qbnsRbA0IjVDBScY7cmSnRX/lAp+1bSDGQyREQZZqV4Zk/nRZs2KRTFwFljsCzzplycVJ
F7G0+6UMVWZX25aGmYOv5zS4LJgcpHbUxhaD3xwbbAzdY+Q84EmuGtQwD8Tg8cfd38oZ9zaxig8Y
kRNo+WvixSSWSUlqH70StbebhMNyhj4nKS80sPu91oIdv1h3QnF3lK94s07bv9DvvHxDE7dyBQyz
2779zYuC13BV7bM0pVHNDR/wu00RFMO2aVSjhCPJ7PN2RXN9rzYkScHVsoMZwNWM/br4MRtJ8r98
lW4H0GX1mPrrRedWWRqhFScVUnV6igERiTUEO//+f+nz7Ewmdx4cNfm/4V70jkM6iYxi3r4+G3xb
xbJo2k2c5Qtw7Wzzth2ZU5kdsrJbGEc4AzGBtPjAkdp1+mjySqvNijru7HV9VKkx8FlRIEs1zx7F
razIirPeUZRSiZ+CB8eq9pjm/ajw8/XT5CglbzkO+T9DSrsSyPYEDC2yvmz8iBMqzvX7q6r7grXP
B3LB569hucyXdblnGhge6kjlZr96L2lGbmLbn6rgVTpw2zgfZ25a6btqGNoLsCwly5oJCEjmNaIM
HhWMo/AM6lf6j18UsziCU+CL05+iVP1gVJoZSxSw5xgidcIMEpeWutfuUbzuhmB9vVS8n51dtVs5
z/hpt/aWoYJ+rWLMjcJqykZMd6+T0U3UiteQFMguxz1AjxergeMJhSjjNytwIn8ZvnWIXJJXNek/
g8QSEDy5AhLnvcrhlL5e21jwQ/4q11MwvxGRYCql/GNHVdZljjSJ5DViH/8ziMSg71vFOJUlrmM+
EwIARTG1ECiOVOx4YmPsEsAJzTAU8ARlLqt/Y3MvujOIr0UrlppMNWplWnuotpBYshzYdkRvZPuu
e5W7Z9t52HaYLr2LnFrMzWO2iIVfnzIHuXQWG55i4xOj8OTYJhSHEr6aY+js9qyVElUwyRtVoNYg
d1VnR4zsT5hNAX3uE5BMvbiNWs3ThHgSul/esrSfngH2pejcDXr6CUQJ4VyzUTBRt/ZTjdJceqmn
USm2Znlnz5R5HMRjmp1n4L7GY+FZKd6lpycq6hsaKKbn9vAJZGLN88gaxJS7DD/n+AfrGVVl8ZL5
4UpkJ0XHtHDBEuZRrs+2j9vRZVKxfKJctPIJYyFm9nH2N4JiA7f8mcBJ6a7NjhZY6OnmzVMCL5s5
QgwfXa+pMO/qQXEgaTDQqq6GCJSVDKUyPIfDieWKqoGrdeP5bXL1PsIYJcgoMxwnm9JTAyt4k9p3
xzFVtTQuQfJRHLXi56pb2CZgZUlRAbTPgWwW0tPnmQEdyY9hmV44P5DDIAsAFjRdr7g97PHfdaOm
rTdUFjaTzKL+nL9lJ7T7RSKr/d+vOiua2RuAmyJ4wap5/ngQuk1zhLxnv/yNbhHKf6BwIwkgk5SF
xWXP+woxSGCmaCSyjzw9x5tTrgE9VB3vTEQ/xBscbnBP54FTceAsXjamEUxXQIyvZEM9K/6z7nkm
cSChu7tMCG4AAgMed8X/YwgraGTUswPt1RyQh+PdNUHuNuTHwnbu9AVLiCJ/izcXjfwIJfauKe6b
tyelCNELL5yoPz1pU4hvXusynIlTOmLbvc/3/p+IEcMJShLVL/XKngxqWdZddlxS2rrVgsNKL2I3
EybW1uGI/g7Wlt554ScF+EzmZuRh+wZVtz9QekTHrKhobuHYgNfKRNvojjNaljyIMt1GuMclr26J
h3gtL1TNAhcMYx6tG8VyMJAbd50rtjnM5zG6wjelZdb7l6ggtZyjwQBJtc/RZeZCxo2dI5BSfVDz
oa1PDTpUC2EXjz538f6MLYKNpSH+3Y4H3V9UGcgNe6dD4H/NjkxB5BMzZIOyjSk1yvSYrpYIagQ9
qMOuxuOKk+6uOD/KZSTnHVxNTxGKfAlBKzRIPGJPrFnJ4YvRs6RY2k77vTZX+RAKAzrBVPnFcMsE
xhpizkJQsrxdI2WguUZdgXqQoZ1ZLVzwzS4YX6R9vgq+f1Ql2hBn8n8jYemsfFHRuijSoJyRQ2Pb
nDxLDayyAODqXC+Fi+3jl7mccoJ4KNAX64c02m68oPlSj1o9Sn3qF9gQMXG49WNTHyDRj0ZJXgns
qDX2i4KkjQrNnMu8UgIA4MTzPma8ZpIOhGhn33exN4/i3YK5Vjw1ITWzIU9wA/3jUm0Jan+KOkLP
YeoB77QCiSDm5Myg29qB2ZmqA8uYtJUoTFH6Rz5Vs77KbIqlxWywCr5yKPQeRtq6IpPLDB6gEpPZ
WyzhSK/LmwgU/2nRxnG+w6bJqpYWaqer/Jf498fko/zbea1h0NGlpwaKNk3wj717kbPRrIduVHZE
ixTGtL1gBFh6U9YoniXkKsDFAoHmof3sz8GPQzhOv3LQCPG2Mse4LvP35sc0AF5+78S7PGwFj6oR
fm21bLRGBfBqv6bIUPuDcZEoWaZV6KZPy7ilqN+rh38/aW6j2T/aWAJGhmANjLytWeFfGEkS2uxi
3wZ/JPxYABwyJF5NYlyRk+uBEEtH5svFNcFFGvlCPd28DiFr/bnWKx7Iky8iHB7GG0EawcM7N9Dd
MP0V1XUmWDsVusyyqtV5XL8j1/ZBji9XZOHCThs8qHMJNcbHph0sRj5TYGBMB3hQc8Vpcjkx92P7
wGOoHuDALksdwSuvqFJkYHUUk2hIxKG+XTptTZE6kKINyn3yf84Rb81EGJwfS5Q915WMnjxLR7Hn
xj34Gvi2eXQBltiaKHPy/ulQFVMP5VlWFPfE6pn2JweAanN6BzNLhLqYHOfWA7+l2Vaj0oYExMzH
ElyPvka9qJxj82OhqA7HuqtSYvMIlTUGgYrQf20r09bwIxjq3qRsdoXtDGHkz26BAlg78ElC8WDN
dBokOGm0kApCihZEM0rHEsNlt6bjmwXAtvL5AtKYovzIr408gYPNRKFjNBM+3qa7T6jNWinEXcIA
c8tSc6/l7BwBTGjBJhiaS1CLtRNVFhy1BPwNY+muxRMxeCfydgiB2zxBVohfofQMQ28kGyOEn08k
zdjGXF1grtRRGoC3z2ZSHcTp/uNKbn1fHqYsvflmJO0NMo3/U3+YNZRViqbOVZsgL3mmNiFtOLzw
TAB27UyRRoQk5bPkBxlhQPDk3JsTbecAvHLI2WP7KObIG3Qus7XhBYe7i/4OYDuOPwP+RVhxU/3g
+xnepHLi74j4z5pl5UI8FAXDEU/X5DiBBmv17BO4acQdYDZvwCVAhob9QUzmmhhXhN4smo33d9m6
anPBIivUzsQypomLswwSAL9gnObZum5SekKEx9xR623nOidWlFDmWKmZvzZEokn0j9ppjP4x5jr7
0MtRVA4DLOvk8SC2bfmE5L4ObzcF+a7kXm2dlI2sj7m2DvmWlTuGqH82RIRa+xFWpN+Rhe3Pl5Cu
GTL11BR2hyU+wOwNTqRW3/UlBg2KyBg8+Nq9iEG7retX4Dd3nIlCMD/OCrBqGxLnENbSuyF68O6e
LZveIW/ljt99SzS9HH9Our0cJcpzbXdbZDEmjrSDX2IFep7qmHB+laAmYk6TsmiQqlmtNWRAhROT
SVLTUZ0KMZuChNDq/QKvquXQ3fUnCBPrRjToTDdOxOLuLKPcYdOohk6kpIkTF+0tE9Zgxn5XteBP
KsvPbpOuO0V3g5M14TXMwN4fzD6PD5C5De2ggufMw6S15Osfh2vlMXuOrYUK4HSazKYVNdLfxoFa
YO5NZhVyCT583e0ZNStB12MUsIg0pC0PCEC7yAM2bu9EwRHKjGlr/eTQpwd4xF4Ly6ukea2VTwmN
nHSkUrzOYcLQGm1JHu9J7wA/hqIajrLi44fF+fZt1kHjUshfakPDkhprwaCm/EnT2NxFhFxjEGps
9S0yLRp0ST2vW5jOIseDQydeiEzy3cNCp+Y9g151lr1oElh1Zz9P43slImiUx+ZVvI2WLw9XNYb7
uYu+nDgEHJ80DNDmq2c+EJqbphcpvDJyYCe+ITbHgba0KIYfXNhMEjKWbnOq0wgXDOhzxsFj3TPv
D+LAbJFnV2Sx1av1m+xbcYZbpub7GRI01IIeSa/Ym8EjHG6tuhzXRgknf4BteEyWeK+YxzAEPjvk
7Lbo4r+yY/TM1gPLN9mHjS15hHSPYSD4f5mIID+uBZ5d2dWe0fr19Zv3SQ5VB8gCnRMqVOf9G+0H
rYoQnXehAfLNCeSbELgceub5nYCU6RLKoJcwSkSA0YG44Jc7UnZGD7OjnBvbFJPjcxnCDbSrH3O5
LB+9yzi99XaRHcEz2RqOeHDWWgYm7sitj28C0nrmbuMAIqZe8C6ne5+D+BYMjeQSh+FXhFG6B74A
ZcdrCXbgops7Z4W85R7r20zPbDcRcWIlMDy4LSn9O01wnI9KqOK5iiRJDfUicT1xt9FUKBe7x+P6
hi05zOVAy6PQ9n35P5KB9QcGi4sLO52Eb2w8vcF7iyQkM8Fnut1DpzQiJkUrmIAYHNPnL9EUoeez
PfmmClM7B9l9zy08YVFr4dKSom7mBAY2HUlexQuQTl5oJNbk8vuiDZt2XyJBIKsr07/NpFqd2t+x
JTmSNr+YflhRgHEuUlU771LF7HPC6I/J8fvPLFKpehsRrUpMf3zPGx1SBZUQ17pvok53BNYlI64t
77syqUdAEnl62xAYHVNtk9BRrQrcWQFiAucJcjT99XOs1OatMcZAE78OmBbCWJo37xFTU26gcRf3
bCi73RqEKOeS7kHBczDNrT+7tiKU5r67KvnupO/8Tkf39S5rANWDi6HgIR5SYx73WUIJ9C3moN8h
e/p3xNuzp6y/3CdxuGejkiKwbSPUMTe/m1GJoezNUJcByuFcV0uD9otaUgfJlg1qjnNrM5WroNRC
C8/kvLmEwwVVB/S2gPgLsyhbn721VOpAK1oAZvE88DePB10Euec46ru9DP3/ohbbFNgxFksXIHQz
thFFcVP2NMRtpbHTjqLBmrDhlHxZRJ7Gu1rrjAdoukK6wsXNFuaE+I9RM1iZKpVk1sxsKn3aC7Ce
Y0MVX+g0sWD5zl70QJjh/BH5KhMtioBUe9+j+IBIjhC8uIWwYZ3bBFgbC3ahFRPR5XunDe5Kro6R
CE8dFW1hQ1lZ5n8X9FgjYKRoJ+Y0uDlZsCkRXK2n93ljz+Qbq94De1WpEfF0WJR9xylsg42+zcXw
+FZtUoEYBHwixPbPTlsLvVqTzeMgLEo+VWFzvAd1i0rdB3VGF0c/ck7V1s28Me7VAudsJDeLC+io
hRfS4Hw3xc/wtp1oQ6IVhhI4qwdA25Vv7PTvsxGkh64Wgwhrunb3TJN9JANt7qeuZTsOhDtdVch5
tK61ATG27K+4vjj5R+U/s42MEH4d5mPluCwudSg2kfDnZ5pHLt9QhOincmwDade6IYRQq94X6/l4
X5UFPVaFhwkgwADlwDGtKMNhLaAzPJEIDf4atePfCfWMHZ+VUznVSG/y9XBBfCmnpuS/gGdhiYPf
DK3D1obN8YbkX/PWAflgch4t8IxSJCtfTNcoTRn5RE4jW3ZhT6yYng9QosKpp+AetVkfaEP5P+Uz
8Urs1jDTSlfFV/mAMTgZAb9oMk219o0A7VwaKas/WqgB/NTmUJfG1cntSAod02MEfzREqGbuKV5O
UvvqKXCELSpiqOacGjxjMfDOM8fDQuByAcMJZHFKvBSCnlNHtJa6/fFgB57alO8a3QFrxbuSF0uR
g/0Uqi+7vQlaIYvUWsAzR/CJIhZUoVlNwjqdArjjOPCFWCJDBek7tOjx0O6gIMwBUB7enj2B6YC6
ereSPIFQ0hNA8pT9q3LYVH6Y4a7TEyFHTuSh96JnKCwW0QQ649+88iNL3ZRifBT6razdHdZrRNPm
D9sOYS2D//gNydPURJkAjBJOh7MJvfLq4BszUb3mB12iFRsyfRLdtNHecF8rtn9LWNIMJQmMNTqz
+wfR1O4Ua7EhTH6RYPdj7SGlX6IECglaPaqt/CNozDRJiASv+/wUhSut7UWyD3hFeC++wMcInBzG
Xe4veU75D/oWhruxn0+vALV1a8UhZ8uAO9X2+e/plIdX1q1PEMe/m6WPQU78Om79Nv5iEpJOpJjo
ZEeAzpTCz3aCcaTAW3Wr412iPCGtOM2zyZ9m8Kuh8fa73P2b1YIqz56kyRdITU4/7hwZqR2ttej8
f1p9oHbv4wourG8r/OFqFrCp/QsRrLYm0pOY/wDM1HlNlhwQRPFdWmqCm9gGRitG8elPaIA6LAf8
hMYRI1xDsKAcOrSZrvZcwI9qSqYyqLQBdCsF7q5vqKUI/5wgZHdhCPUCmZnsCIWNzSqyYqyATf2E
OL5PZS6xcxejUaPl+XU4Hxiui3Jbueoz/5bPl3wcJy2UFr4G1BjPr5xS2NT/a7mXhUBfQv/tLF62
Z3E+YSo7kyKyUi7MSc9e0xJqNWaRo+38XLCloeGdGKm3HZWLhaK7TWlXdqOmNJWUp8odaQCsye01
d3J43yD7cSWI/ypQentYJGOaFAy+0wsb1wuzlzk2lC8XUq/yBM/UHddRN4f7oNolTpIOYDFk2/ui
Q0orQCE9Qfph2dHa+nlLUDc3qVasav4il3XqieEHA6g72VG84poi3+AvOg5L1OFG3olGZQAZ6IPW
+nN4WWkXVVuyZFZFUwzaXA846vZsLoU4oIQ7LwAjyY3l69UwAgcfxI4q5HnCoVmbCljNJjVcbBzP
7d0U4ESCmCNsvJuWoeU7+r6f5pC16ZKDqSrsojoNHXN0hhbhXR5AfIE/zLRhHLfg78j09rF7SsBF
7Z/A181ot54oYb0Y9VRMPmBeTALNPegdMeQhAohli9rhg2HOK3rJactLFTDdOz6UCrY4gqvl659V
ihrF6TXQpDd7DUTJ5yEjH3ne0g5TfWFt0xRVRBus5gqiUXvp41ZiqEaFKYO38mOkgBCnS49WZLdG
Rb2Z5elKWnHQ0pcfS5+H2feDl1PtQP13uxut7jOJv1bwp0DqUu+2hG1q/CCqC8qqIubFEhHmCjEY
FVwdURlLeAGk0yiGiur2tC9M4Q7usiPSJGuphZq/Q7t/Vu5nNYUqkZh3PMEUEB+W8FCwgke6QlK4
polSQo4vrJWnHHThkkVjfwBkm8I34+z0snq/7MFnzzFx+Z8O1RSRPFFEpnT3Mwf0fAtx6hc/Haqt
rnBcGD5WB7Nq7ca23nw4o55Cs9yVOxbPud/0VRn7L3meTlFxGd5I/5mkbQrr8Bw7jXqtWSYh3e6K
/SnNYrSAnM0oEfzSpYsbgIpXJN/W7Wqg/r5cvUun754m6wsH/g5vJVHxicIH0aq7KAnLV4BwiMqX
KsimDBhbSyej7mWg6XnT2MN0jUd5iUnxk+k53qK6K/xkW4YKtaFnft5+J+2evWFcGsXvvkOxj6sf
co2FDVNrhPdRvkPAim1Vq9abvQa0tdo5OCKGqTKiosrTnPQ/ABTqkd9Kp6oH9l0XFQOJ1lg9NESj
6las6ykJ/fNYNZrC8zarV8sqmFAGyUoqgOOoGFn6urut7pKUo2YCqaqxDu0ZD/hSFKRcfdiSWrBD
Mqk/zQ3UbLCP+ipuSptF8eCCLmWZaBBmQKR8P0BbWICtQguub0of5CrDmD1OfAowTdcHefdSl1EP
CrpRQQlCLcmmS/aSS10N74em1LPz7lURd2FQ/UhuIo0sTPOhbnvfPQbNMtRUERiuN3cUp+zE001D
pOac+BLYx3wC1+YPP7ph50o2WMEZjQE9//H7MPAVBThHJsi+E/9iOvO+l4Om6NeCtWUiFgIFIHti
SY+xMdj+HpHThc2KpQEE20IX965TnHXxxOYUcEHFXYw25bDT/TjKYxedUxXVXpiPzEHb2J6VL1WP
KqXlRRSNEyZ5cgK1k9Unl+X+BcAN3clD3fMzrAta67RYhX9Uw+TiYKRkAqJ8V6Ct6brjk9hnJrkT
WkB5HTTbJLkXQGEW7mctPVVTZmqmmwmVPXY0NZy5BjwrjroDblsHqqs7EZqwlJtWNL/rl8dMuUTa
lIxcguUHdW0qTln70QVOnolij9+EouI4tu0AJURfB/srjw5lMdhAjTyIjHTp7N+tAcACR0BIZyGZ
7W8M6MUOqusQyDq+TTwq4JbY6jcqQ0cP0H38uZgKrZ8ALmYYRCdNfbV0XfOAdK/UnowAWfT5riYH
URBFVFad0oVv8I87yJnxVd0nA2xlqjburiOQo5DgkTJ84D0TLL+THSNw1fWVYs2E7k1pD4/ZCFrj
kH4hotMSaZb0D+x/3U2py/w/1JBCF13kws8FNvsYHjwGcHyxLijYnvfzy/uCnN+NihoaXvY/cA5p
JcN0Pk/6S0eVMb5YaTXcyuI8yCkp1bfgLszt43bhZJ7/GucRWrzvNr2TOKQK5mRnbSSRyDsqA2o0
ywSdiLK5gykkLqo4M5gIyJLf7ZHCz+KKWZwOjqSNPTG07RTlKBxR6NC02H7WXcMo4+cY0okx5n+r
0XzcbMQ5Rrsi43iWTEQBZ5hJjrTyFB92BJEga61ZEkmnKUS71pAGXgASEAxy2wOYbWUndYH9mkMo
Fb4X/QqeojbyBGvrw6yFFO7kjtqS5dOxjKl97UltCfc+L758fEbRGdglBEDzBfQbwMYJop70w6hO
TKx7VHvFzpErfPC7pbKpXSaD41bvJk6iTnHAhdhV8d8eEX0yU1+jHssv6WbsnJr+nxZiwJRq6gNW
7YHDv3TBPEkdLwBYpcFvBd3YvqKFLcQZ7cqXn/wGPHFAlDVyNNO25DHibTFHXoE+mSBXfrP0tjrK
aZ0WJMIBrdwUVAJgil8CiKn29BCGfY3F3G/8DDQ6CqdMNjbDnCFxK1TE2zwgupX8rMXjZhj4XIuJ
tP31dxhWdYb/X9EAot3j20zPYC6bo3Hn/JA7YoYLuZcmioU+T+lxyumXiuJgk1iIX7KeTuSkLAPC
DUqzk9OMG2AK7IEJsLbxAsZTL5BAavX7rHU9D9s2Viz3ETp4WDX1aXJC3kCyh4+WR9cbqu7d+GO9
ny17RgousUUQK4WJXGmef0UpzYDqNHjoPiJJYx7s4lsCf4fBHDk52WLhIOZ7fz/Sac41JpifcaKa
FySBe8koJ3WqXITjnfYBsW1XiFee73bXUulKZ0ZkuIzmvq2AO/sS/0IgAj+FO9s/WsFfI6AGgicr
0Ra8mWJGN1WlnI+5jZlHc5jjj4BMWUWVmKPTc/5HyMzt0+XaBNdiOAqQQ+TARee7xqFPynusrcrH
CVVGOiRBTCcRmlFfPThiJQJ0x/xynQlP+6RAQskPAZHy7EtaIHBLvvfmu+IXdGjVLc5vlycpdjsa
ibJ7XAVw0PYmxnfvk1A3IIGY5UzvZMSVZftSVaF/2FNBhsA/pFNK/rKWNhc0dAOn0kDMorPOTFCR
r8abmq28T0JmFWRHNeix1lFb8E9oMY39FIg1OyTJ80mZHs1n1SHbqgedLzqvUEQz87x+i4MHCPNl
W5IdiF3CJ8OtGfd3LWwLYs/TkKrybWdpp4K9NyTOMF0A1sNor+wVNm45REo4qLZlTu1LzoY1OVn9
CUcHJUAIcW5bUqEF+0LCjV4OMlAMDO3fZdT1uQSYARalXvpw52LT7dvZS3/F1udcIS//Fi/Tufnj
6b76h5OoyOJYG+brABpOl7zexyqI9fSslxpWSGRNSzP7gUUy0rxqKzCij5sWVRrEUn7cX2ojBXwf
cw5/pzbUzVt1tXvs0HDcBFX/q53nb1UQ9unMFpr1DQ8YQD1ZqKlSAah7ihrH798nUqAOIPS/FOlV
VL3dya7cp2FAd2UYjUnOdvmQEAbcK6RYcucC29sSJKkwDqBtxD2WB3VoZSuwhUwc37HYflgIunMR
pY9gd8tN1rT2YH4ZDpNuCA2C4YF/sv5miENv5bPNgOGJF2BLToTR3cLnIJYIE5CYwg8fWGAaT9jI
Mk9CgTOB5DLzX2VYNjMf2tnz2NKiKw6AqjjrKqsLNyfxsFhorE2nQnZLCig8vMku7bETsZKoWWEO
NYXT6ML5zYjUT8gn+pK+McMnqAJE9t6wTol7DTK1T+RIflcB5cBtw2o4vB9BBJlDS5JzhkQz8m4A
uYkBxjy3slaxx88skwglTPOOd4EeBTbPWrBt6Ti3Mthq+vrYMle6Qqjj0f846fhzothkDs+y0Zok
AqaXt+HowHharWgjU3VahGUmAk5p9QSJFtd2sRDHKmgkVIm6+f7mRiOgHKzf9rQjOuaFidIqbT8M
7bS9EecqE4mOO0eCtUTktZZfHERoMFn3hbWm/EAX36dRNeW6K9W2hEI+MggZxGg+I/Vchzo1PafG
1uxeKv2HzD45yxjWSlbjEPeOvAPtjqe6VCOPXz9QsfszFIhkRSBzvTS9GnvoBzOBiGyNUZ5jFfI0
dRL7WrlXTtCoNd0xNYtDEXqnesDbgFkNBeckSbR4SBd0LXIZKLn0CZlNcVTdc9BVRG8gBwJTPg9J
M1B6U6li0+GbfEKZrM/Ns8IzTdhTclWDDa/65VkCO6A5Ew8+ShVdnzAjH3cFlFXV/weiHeqv/RFd
MCIPwc28PxDffUehibsiNdC0VyeatDO3Re4TokoLNW+L81LFVBKUrvbtIpHchoB6eR0K/i7mjycS
Ath0+yfPBht0uHV/fJp7rgE2SM6XIkjlrgL7s8QIb7L7eaWkA53fQ1kelXtMKC20q8ZmI1rcLcwz
07hTU83i3xjQbRhFJfp3vuPQLGgfNbC5dhxeWi7xBCRrqOh0NjRnzonwSL3e8jxYVkPljaO0iL3a
TFnXUHf2Q/LiSaIW2nnOFXje4K8DPl9ZHudqqtF7SoLjfLkg86QogIkkgrx9TglQgvJaXaO7S4eJ
EqlfWPwl0Q66IWLZ6c8UrZTRWtNM1j7neJX/48zhB0apDjt8mNg/zMbskm0V+jcqWeyqGCqKAnE3
dRVhZsrgwq1ZwUzbmVmDLcImKv1bFrKPmWEORsHebD//WUOiPh+sLUSxx+oiAKi07BRE0tfbkg2W
q+CngKSeuVDo68e9nLloitRsFDYJ/sXNrsYcPqbR2l4LCvMFrwtR7g7KWbROuIUHplY+oXKHr84O
lmNTU/FqsNvYw24z95poXPJKZ7WkdGqwYaYiTF27BvJPqhgwnc50gVudaVmbzk5bDAjIc5UNVFSQ
jQl504oyLLVsk23G5gg+FcR2LXkERFhqsm94veadeWcL6kptYeHgOdVHqjLgv9NmhJy5JoprfTiH
9dUfAqJUyv8v3me2n8SX9PSP2TqkaO+fwx7VQbTnrwVJnQtVP9nYBJau1tiux7fBWfAlyBDCo0dD
fvj/jq71NtbRSwkeADAWsfLmDQ0q669hZ9FEVGrUU4KpMRqmjpWp+zZiQP6Fug03bXb4kEMjz/qC
UTykt1zhGZ0kusLF4hqKYme/gHtP5XVeSj1UrntX+cUK0qW+4Ts7pEv10/W72MP6g9xkvgN5gIVY
QI2MVnLRKpsYlZ94VfTNayQwswfdw6YhHkl2qA78yV1NSZt8QAnU35i5BwbZRPixIOq+WVjXM7AL
ETMnYHk1urpoe2k5zV9RMTaYG6IuiskJ/FVVDcb8xRR0bVzAL8dMlzSROUujyBFPpRxkDfQSsHpj
KNPUin5pZOmINDapK7Y15AM3XVFEIOBsgT0OeUAbs9GNqIc5TxYDjXDZLVeAnUASOwDr3bhv6GiI
zTsG9/O0dx13n0cpmZBn6siKsrQI9HmtRj9eMPuBZyk03Ij5GpiYLy45LJ3Td3Y0N6thberEcrAj
HHcqGo4xetHw2VrBqG+ZN9K5fRswZ3bYgH+8SMJTPzc4OD1eyzWcTZnRINkNl49ZAINstHnvl6qM
cKmAxYKt7NeW5CMHmK90iHerIEGEV2SKbv/AYgZ1O3bBUdN9aQhIdfkEuP+dc8HB2UwbG0B0xYBH
AdDsLx9X9QG6sZKqku13JTkD/3yVR/SroQnUrO7QYoi/pR5CciMTzh4uL8G1ZN3lthBu4T+ur7YT
HSGgf9BBym3UyHd4IZrrDpz7NfCqvyJBiYPf4E1WlUt3+h/wwXBgx+GHwacu+EW+alS7tEkccjkE
vDl6xYwpIhxXZjt39dgbXPoinV7n77Gzkvn31B+6EiPK5E1I7/Sbxtgy5cdbpgy4fjvcQVQTUgdD
8cqYdnrJK1OiiyymJ0NHJPrIJwh+T2XEMz6CT+WoTlmYtWfeqGbS/3Dd6FkJ8xj7M7tiFFBYfXHK
wow2gzCWsX7jYvgnh4l8GVhNX8zuTGUOdPK9d/AAkT1D8gGzGeiGleYe55wcJqCZNP9DeGixzJcP
4CwjspTH/DGLB32MotoRyt90OTAtWAHvGRrST5rgkLMsGO8KPUfai12sXCq0R2mDBWXAi0eUAyai
EtOvvAuhA+TVlJ19nHb9ZLb8wd4KMhW8WkNLN3Spi6KF+jD8pKUdZo9QBv/8pZoTZS7THm8VH1QF
2j9lv3RJ0PahksHieWiN/LDzjgubq2jplI1Zn1y6bFM4PQkSGbvuaaCxN3dx4Djs9v3f8OYVilHa
WXErT8KO2V7odZlqbmqJQM3+d353z6mwWBUdhXNhmqQ5j5VVIPl7HRSUYI/USoSj5ccFmEPsoITX
BuqOL5gbP+m2Umb3oPDIjVggHSgwujqk0BNrTUDZq2NDmj8SXqFnvj0NRGdyxeOH/HJVqBONoh0y
Nb+Lg9/QISnXj4JmJbtZ/HikeR1vXayJD8HstgGKN6PDOY7RXVETlYTsbUhmjix63LIeS54YJAho
agRRMKTPOqk5w99iuEOOYast+AWhvqeSDMHimnOYBSxqEe5vSbt8Qd3cUa9PflkMWZpVqhjGMlJi
5dOcwOz9xo841axqjgo1SNBnsjwNJuWP1wKaGchPYFX5AxaCYXZaH/JCLNlNM0Shg8bLNoIFdnSO
0G4lerY5xxAB/e1f+2AWgUrdVid8BEPlbqipQmK0R4OKeXa3oj4xI/dWcxakFjObChcCupnpArbY
XW+o1v3wqPb5CRTW2h37/es5YgSZ/4AoE0QFktjMvS9yVxBDbawVQB3+rrhrHSJ0TW2JIiueVpCP
7NamHYbSBS+W3zvCljlm+748pJngHVqChvzSRVP41lHBJ5U4c7k1/bKN1MXq6MUZmQuLMDP5s0Bt
u3Afo4yzf1WkNl4zStPuEl+IcHQLZGHsqjzQd7JUzpkqpV7cGzccBF1ZMA1p13NZKzALuatkbhh6
RnRLmRSxwdbF9aMT3q2+fOrZAWBT/LUaDUWgVDwvP01XHBsIiK2LEe/XaRvnYMRTpe/FIzZdqlRc
Wn+mlS85xgb4FS0nxo+N8PmaNeTRu73jAsjYd0kvrbzmaMKt1ZmP3HQGSUwrDVmuk3daFuY9Cw3T
k+7yOaPxsdfJRxIc2csoAZyrj3eSQ8PfiDQzPXMEr8fzkckwe5ZeSAEtjGs0TzwFjIM5QP16IDps
0zHKbsxwBdLhcdRBVwSQJuzzm+avr/VSfgHaVaQmkoNHdQCEnTOvwX4Vr5tIDUN+pQUAxPyGzJ2Y
1dn27XNfCr4gzOyo/6Nby3bpUZ9AZehXV15S9lLDB2b6B+qrBE+I9XkKDzfO+Jatvn/E0S8QtilR
OuOKgi5mOhtqJq8bMChRtlSnzahuwCVF5iB6jlPhA1Fgf0iENffiC4CFaLN+46/8NVcXzj46ovWd
hJjh3LLTjY+JEqdc2HP+lSiZdGkLpefSOvpqu39DXEvkoX/zAVnKge0cipXBmrU/pbft5+OzzNWV
aCPBRBXlr7jeYCGJujwyc2bnQTSDsLr4aU+Y/AfSsal16vuZFL09yxOI6MhLP0sNHZRrhBrSs7dU
yrElbEyABU/N+sun6oBtiz/Do4u7YXS0F2HUs+E1vHGAYiMkBRfNACfh6k9g0aoTjROHVOnUVeji
KJaaMIIrk4aCLUtilybs8AWgYtKyGIRfz2OS9oQMk68SosRZ7K1wiKj5NNVfOruX1IB/J0wbbXwA
D0cghJeBbI2znZkvOg3jT7PdfnsbXn2eOF//VEKPAgnC051r3G2QK3XUOe3LkFPaGYVjyptspzeY
JLL3H2W5eEoqFxuAZRcb/Fg2kTNR35WW7JJnUtS12QmK0X9O9ZSO4dFxLOTynVI134qnm5RzXjWR
k6lsfY5J/DQUjfJ8Qwz9a8cPaji4ER+J3sXRoReNiEAFzqS7Nv83hCtRx13UjpSHpLzp3Zylxkoq
MiLdj8AnSVDMMrEMFFChqYBQbnk2mDuwsEK/ad9ZL0w4cXfJ21MLN1czVRN5bsTW1CLMtkqTaf8D
1baajjzNMT/Wm+wfaWOFjdWa02s6rtt2tnQWAr42u2rfBgh063Z//RY+4ytnZhMyvRpXKJufFukk
wKaQswzsYha/piGYootwK1olU/vxyrPo8NakIxPHl8eAGx9O2C2U6CDOdLlLdCkSwHwmiVegPLyp
FcKG/QjGy8AJua1wAhavBdnKbUFuLpocNiTjUTSujmZSWn2E/aoW0qHPEUzbaC9NlDNZDoLND5XB
/JxFRANp8LkaD4p5MsDCA0gNzS1hTOnjWdGXGzMxjNFbuHunpd33uoCOVif1jUQImLnQ90fbQ3m4
3eC4QAURfFn5Ri51xzIQ+kJibvQ9EkS0faLqzN8zNDnnxvhG5Lt8yRKE5FPI0D1cqGX/APZENHfU
2wvZS8Gts3hGfO7du/Oxh7gKUIA9vv8YVJa8q5iYvAeYmm+q8wxr1+JlOt5qgnefrHNEuw7Byn6Z
MhaM07iHw+l3kL4boeW2bMvy8ZPaEJCBxYIwehmIj+RcqwImaNsiEPV2GA8f8RF7s2joSZQYCB5P
XVCI0QV+KyJKcAvejlg+xjuE1ftnyvJ1sgFqwF4K9auPoL78zhXCapPnYEd/vxyeaPW8mYz4SGje
+oxhA7tbZuaqsDqDAIjbHegkdnfyFud68fxRRIb1iARtf7CDRC9ATBz5R/XslVanz15WSL0vIZX9
krdCjL3sep4zCHEGoMlEnHWJ4vk/OttxyJwUXPwF23bkIFzJ6RzRDdh3dYqnf24Z0Qe5KxtTQRw7
edi+w9RXeM+n0FHU0hycP16dBdGrZT7IZFXZbfX5XFFo8tPFfbOXEw5MOu96XJT0TMQy5DhGLvRJ
ekYd/j8VaJx7WQhC+5ImhbYZYjq8U0KkfQrwmJ5pzyFD3YRadIc/YfgM1XxZ3Z7u/NhxyEbJnM1F
1dAzA1spldcczafAB7/ldBMOmbSm38N+v50pa0TMTODLUyBIPHOn92m93ToND0l0bNhKN+MwLHUz
y6g47IMcDAKoNq6P5I2Iajf4RmMj3f210gOr+R+Dk9Uqb6oYp/UR4/S56w5UTU5jUkTqfiGbZ7v5
rnYIMafS5x0KrMupVIeoiA9LdtK4akU+ZgBQ0zJQM0spYYiHXJGX7c7cyUwUlEWhzPOM7yyJ3aR+
40LrR/58f9EG3F2riOAWJdgtCcmB7cAQCz4IGoKsjsWwcq8MJDJpfXXEbVZaM3J7TRvhPPz41Mml
2Pqd38O/FAmIgwyVZV6AkDvNH1EcYK3Dm2GvlDgtuKgxTp3quW45s0NTDmqRKJ9+r+xXZOZ/NE+q
a/PB86KRrvzoub4OLwdXATcQUvU13lmzFzXKBM6l9nm9hsQoBsq0GfTtkzywG1mCDYQuhnuZg28T
9pPWZ3GVkseiFgcNPs6BegZe4CdRI1Ya1Fqe/W4SPvYYGfojse0vRWtjl93PmBEJzClcp89WAuie
njNdyZ916OpJYGgv5CNgK/EJifSvsnmbbrgplVeUxnn1HlbrBj11bn+TZqbijjFEY/F1nIr6GmWb
BzsoXYOZDnkwMEWFYDd/7Ty8ijXxrEag0u2dsEA6WodJLBefLiN0Yl3/Xrm2PfCaOR3IVi5Ubc02
N4VHsnDW0L/FCKmAT1ytxPWdegMgG0GUrYSx+8ryJTZZThtawgNp6SSwrvhSfu0uRO8OXcq+uzid
7d99gjFfzH8nBxyZvkTHSQ0cWONBSyhnbx/zKRr+b0YJeBgnx7KnQH7qrnvtW/+vHlg+OKQMeMiV
2w4Hy3FsYJKHm7+9fmT4KqVpzRQwjUtzJSe1CnZFFebk1Vx+DgWK2mSEiaw7BkF4/cK//6sArX+A
siGPNMF+n8l1dMJ/nZmUD9y8yp0hX0+nSBGO+6X9If0V3QcC51EXpj+O8imEI+MXvkaPkAlx7/ax
mOYcCx1eHqSQ/Iis0JJrfqC9a3A4Ec3PysGr2HCRMDGw6y7mBJcfIcsJzzEF2dwvSavE7Fi4Qz1B
RA1EniBdGPHf52Sv+X3aWcgQf6ktEzgI74JE7QBLg8bIT7dJYC25E0wB53w+GA4quTzSMsGvS6yz
Rp5Oiigf5fKEbtFq1EQkB+l+QR8fKbKyTFgKa+UmcCLxh0tycLpB3Vp7sdRuryTzPwFbWVs0lWQD
fvvALIz3EXVn18GUOIO93Nua/5Hi0C9/3ntjfCQVikoRAa8mqGr9M1GQhC11IVSZL/XMh+fcMn57
n0K/CNlQJwOaplMzBA8a/XtdFALhRfuhwKFs/VqV3ghyW5veZcT5vobgUUNZAPQTsdq0Wej57UTE
nC0RZduGvrS3dExW7NhcD7hkvsO+b5cn0LTZsSM51J7qtsWdxjBicalo61WN5ytkaOAxOUn3M6VP
4RnETL1jCqvOwH8ICV2Yx0L6+wJSUv7IZ7Xu/H9Ea0QOyuG2NnvpegIxkt73z0n/Z9B/BcpaYN9T
OGmR/vm/opTXkgNML9Mwp92ejQLAn59s6keX0lKhAlluZlSZvZnFv1WzmSABSEUPI15ch7UUbK2L
f21uHUjmbKrzmFhVUFbbXELYOdqmM5TqW9zc6wn+NvTzFPMt2m3zjElGIO4hKcn2RXgz5Ctif694
mqRisz1LRIInqd5XtPy5RC/Y9kUn3CUSuk2a1w1QboKSTpn5m3rK4VZX940m5kMb3MRNVIcS53J+
WFOTzpaw0OtQArB5EvGavHPLoqEqyMggHCiZ5hpe4dCtHQ2i2fIaP8pmUw80EGHnTMm/flK91vCf
KIGlnkAJ8N8FX24FHgjxPd2EdbP0i8Ka6sZx70KxDUaTYGWxDIPBI6Z9y4UpmvuvjgAU4HoQc2TU
2X5/tPIZOpKZbYsm7GqlKESYRNMnr6fTXt2OCr2rNZ3db6XTJaqLm0TAkQJaAYUZd3ogc6QWaOs2
VMxMg4P3Z30p+ptBHYaOfO0RrEl4hLtta5JrKHHw0U1O+cDFqL7HjgzZpWvaqHTnG5ocYIfULRff
whqjGsHG5DEezqIFo/ZNNtX0bwZjfjNKtpTknnxyz0wS8W37kTCBt9n0r+/ZE1iZdnlcE2xPPoes
gmhvsUvijlFIPpoly5kIBJnLDa6676IJ6gVX19roS6VSoBBzNW1vy94Vqa5xvhRe+vrImDHNvF1p
RRjuub3250bDzSY0sCRCIBuOp6VQ25wEdNbO5pUfKtTYS/U6pxThZaDCeuriPnkT6tYyoMN76oM/
wc2LIxd3ayPFS/f6QOcsZE2hk/UHMiwZSxOxPvUVCzppl1HK5auhgwdDs2vC6oDV5x3E5aT+x8ts
Yci3+6ynQzFLgi700iuLi3mexAOEusPY9Pe1F9yQvRnIQZU5nFWVyQ6ApDi+phfvj5WtovbQaokM
AUkfYjn50345ZBv3CodSAFadmPhNSgG5DNwQz/z+uNJPggjF+Fr/wHWn3TEZpf/L4ObdeCx9Fs+o
w8gJshiViDsRfgq2khanKVwk9JyUo+e9GoTmG85rZZYA0dycjhtcm5NCJa0ZkhH3isIUb00acTdy
nfqevec6wgDHmj9u+JVv2M45Oz8qAV5xOZvfwWsMjfGmXY5c5t7IP2deBZZJAV3ZgF9eXVh9PpCG
Pdu+hXEpDi641cGEF4U4oclBoPuS3oJ+1f2It37acCkNwb+yHTHhOcuH38MvF/gu+Rk0bKrBkl2/
dpF9i8DdGdJaHMeuwhRYeblbpZlAjIBBClRbV9CTA9NRp84/tbsZysjn3dc7CD7kXlu+DWkV3M3z
t3w6yIpeA8+3oLxm40GcXUd88A4cS5Xt36qvTrAYI+daNVfmho48CUqKIiVO11kP6iIYJhyD0J4P
ZQ14haKyaIX5ZqSKz13dbdOL8cACRrTmXZyItT+crU3IVATMN2dtNxssceacOxJv8290PI6aOn8G
otfLbVRdXsuUcHf5pWvGp8tgk3CyOpqqjnS3nRYEq5eFFwESj9Rl3YI/OMmVbCkMYuzaydR8PDzJ
YKXH6gS9FcNHlnSEdkmh7mra2inZLaSM5++NX7XjRvy0yVAtGVB4u+WmoWb4+yyq7uvd0UbrEWWl
NnkQR+yXB5wTFyJd6tgumAfKkCel9t3ZUaubveNROsoecNzZojKI57BlhuOKNbrdEs7Sqvyi+wsL
FytxpfmM03ilT6zNd9vH3tf1IjRG+05hnfCpOP0fa93gQoyLq5VH6rjgegbY3lLW98TkbcAWkSUe
ttJodvYNBhNKcK8wm21dg29eNDvL+7jWSvJ7D0Pg0eQd10JWtgEojZe76mfWS1V/rGuEMd93fEeH
Gc45oJqt4RDnbozeESm7IrmLn5F+SOOWdimCJFNmCVSnoWkaTsxc0AWhY6BinFkZtmoqkcJ7kwGs
ffZRgy8HAenVer9u6N2/n1pE8Zq1UtyLgAsrIyKuTCXuEEle/QFRdoW+PXGPcAgAg3fpxMPS/jN5
RDHryhWSqR5QHUHdVjdGuebfR3GwcKOoukBtZk5QzXmU2xfuO9VN3aIdPsWNXv8vf5GBNbbxfDW6
aDpHJCK9IMj68AmuwAO2aXgjHPm2gwbwgRzbZ2oOEXmJK2/PbHbHmn7mkc7R6OGzei1bx7hf/0R8
LUJtzHbXMsTKu1z8GkNi/xGeeht5p/zFdS8aMGf53hhfXixpfBUKBB0oaypTqMKGn8pLcm4w8tcs
iR11UiHxbtVPXYA4KqVou8jayvhAe8kAG0w7Dtkvm9VQFQnI5o9VqBBCgkDo3ubH4E583FnkdOgA
LSlZzOUXt8IyvUtb4Uaik8YjHF42eT1MJu/q6VN2q7Uo3DDOLLYdDNinx5A4pTYw/iVyskpZAib4
6xCi59xZaf79xI9S03zkXnWFmBn293ZWGu4mtpUSrDPdNHm04q22ZZX2ewJSk26b9Fb75fJ9KsAy
Ser5e4ELTyYDL2b0QXE7na+Gho8wTuG6a4jWuLzKUuQZXEUng6KSXHiJ8M4hK2uXyFKfTx/8ohQb
BpzwV5B6IkilygkggMkx/s8oo1koYVdynADo2070hML5YqSCx5trIsgDeYKCgNcVUTty9PvroK8I
3lldrGbmWxW/Cf4L1y81u0+5XjpLuo5WcL9DXoDkKReyL4c3JIuzwvmx18n5kczvnoOvNTmAMuw2
L9gGHpK/klrsE0ZDnjqf4NA4GegoZ31b4MlzNKLLJ/j7e5WPWQOuspVWFB8fOnI096jKep842cCo
yZC9JF6gDVqsJQLrWfZfmrszH7nVNbj5tHGqGzJ2ZO3qvkX3tbU+sxmjK/cS4oE+iDw7P8/S2T63
/U3zgmz2JxnWKCwK3uxe4mY9vrKzbsing3r5V6fw9X5J7wejik2GQClo6H6gkLW3TqpYs755v0OG
rBZqVcuGDD9tZjCus3DWsMS76cD2QXJQQyGFzE5pb4F+a1kzZnKo3+gY6Vdy1IvO4Vu78egihz+T
SUonv0yFUrhqi9BOQynLSuBLUYPCaY9tH1qQXXIWqTlCoxAq1DiEkhQuK3S2yGsxIB+HIF7Bo9+o
CjRyg9QSbSmMLXOKvpRHIQpaqtJ8ivcFRvhSgFW4TJkw9lHda1RA9OPq6o9+YZlhgAzCei7/aSdw
JGP3vBnGcbR0OWL25gSGU8PONR4VGfUA/wLY+GkDvjKhpJ0gk8tQRyu6ggyMZtnehp18zVC+RAd9
iMtS4SDIJvtEStG33fGSuLQZrmq4HxHuHBGtFLJTAPRtGmvDfHzKorPtKVNF978HOvpfrAJeLTaS
mbedRMROGkrJqPTKzB4jLn1NFhRY8O+WkNsQKiVI77ObLcH8cHHXPjfIGh/iOYcTb6OeE4C1Jppt
il6MAiSCTk3I0D4T4pgshYJI8wgxfZpCgoF9cZgvWyU15LMOe0rdOWZeKt1G1pxj+w9/ciCSXWT3
2ZwUD4Cr9w7zhYq/IDN7gYpUbc6KFkM8Vui/+8Okp4MD7SgiKkUAN+YVmsaGcifX3jKvaWOrumXZ
wFxeDkS26h/1ucoZzwJjn/Q9PckoH4vE10NWSwDopHhApaSlg1z7GXt2N/tVCrwJ/uoji062rsDd
UxI1/c7kY35qIZCnjAqFSLMEBa1FsiL4G1/3almC/H6aXw02IMJmgJ+JoWMDv3DekVftDRDJ6ZPJ
cQowp3HRWQ8m1wrmWS2DQo2KInthxbIEPD8IRCFQ28iF8ruANIuX9iIlS2AdZqU9gJ/2T3B4/kuE
ovS3NR+6ByXjz8YISOm0Hz2r1ZVZpSPLuLQMnqifsLZB4krRDVFV9ksE0RLRRliJ1YJvuNWHaJ8p
Tjdps3KKIaYZrsueALfFaWKIJIT+p82HagEiPSZABLm8YXNxDls7FIsP0LS8gdvuWIX7nlPwD+oF
5livxmt94qiHA2Xw9E2N/XO1RoZQ6qEo9lHl9GTknZkD2/2P4guj+WchwZF7ea5mJvZbts7mw81l
TSOyOwhgzVy/qfVgMxe323K2CHoBHJS0356gu7BJ3esdks+DCHK4ELtc5Oe5sJ0m160I1+UHvSgo
wn6sB6MwSbCezeIs++7U6rxCGFL79uewEkfixxPGDOFmqNpQ0LJjulPahDh6FBLIGp/VNV3hy4o7
8KvZQwRJ3O9h7k8YDYVyxRhXXnzDqhI2nWU2k2Z+o1Y/IZSpZkkD92H/mCaB4lrdbmTYj2OMq4y8
b1Xbo3T6yCCd+P9Q7ZBgT7tQ8tjGSbb5AxJ3DJq00xHgblt6XeUySyXQGbdmZapsOmKFlp5y8F2t
/RuMawOp271iTaflzti63XolMJDJ5w31HYpH17r6UJD7LMBBpqOwWa0in7gDkM5Sih9aILx7xQk8
MpdLsL0iEgxHTLp3rMfTdJnwWuupfDk8XM8zD0ceEaFfLve4HI0PQdxfsJ/L28n7DjIv4FnoyTvY
mde85McK/b0ju86oyuf8Htc9OKLVxXi34K25Ih30LVij37i3ADR0RTpxEK/CIj0AGtSNuocbWiao
DkC20hugBbJFfqzPuDbyRSL/zmcFJjKFOVPNfv19fl7Z8N52Ty7/KvtCbuscythUHqrWFs7uQU+O
ineDRX+E35CYtbHXwI8Y7e5eQa4l4dnKATu9zDwQgt0pTdYQXDUqGIBGSvyD5rrvHWnGHuERqJjv
YPZk2PfCOZU7qwkqb57Hir340gf+D/v4FkCFgLrRtXIlTLY8sjtfSt1CuG27dMNng8wZIVEYA3EZ
BLzr4iQiaTgKuq4bEwkzFN07a41hN3TR1/dbDrWoT/wvzDPRQ0QjQZgxPzcZ6wX/KIzYKYZ1hoUk
N2pqSknmfjKLlM1p9DTyDAe46+cL0cRxTO/u3z9clP+8NPyilN1OLiUyOoYojo73J4q0qpDfNnHb
NOK8nRczXu1lFKGf4GQ1yje9BqrMOfXvjhKdVPXkcYg1VdA0X6rZVMZz6oYIH/l/6neOUYQYvrqB
bLM1X7bOG80HtkMjQHTrdPBjk2nAJUW+L8mw2CtII5HhXYzkROHjv1OkkmofzotJWdqbJpvwLWC/
nCylpHyuhGyAcZQC3n4UpchunXZMimQAqw/Gbi5s/cm2KA1SJUoB17IFR1eVwYFbXOFms0rUNib3
ijLvMj1VDR7ZcwDdJ+b0F6nk0y0d9iPJHRyLNTobzBXOZNdqBlWCPzjfddAGrOhpFXZdxtEb52ws
6HXFwHTqYJGX1cbds1+PIiTC9eluel/8oGK9SEW7ffig/sablosYAIpBV4qAMs/lkAZZLMyNsB6w
iBXPGUIB9tXnaWPu8lEBOAjLfHi5qD118/VpuYxqc4bGaecPqtulDBQz/ezW/Jzb1o7dl+NkErO0
cRJjKN3sADv0B4aH4gTl+GoxtFoYKp0IWrKxqgLvFyiIw2RcqgvkBub8kBHuRiZxO0NrcrTCnEFW
JVembcOvO8VeAQ58g75xxSDA6IKlj0WUYR87Sn+FbmTtr9MrEzdByIdUWKVzFt0m7qWQhUCxVKTX
Ve+vCS15hBpyjDHehiyErtAkMO0Zcp6NVAC2mTy1JhZg6ZPmCoXURmKoeNBhdJM6lMYDBVrYpTbo
k+lIc2jaOkF2aq61DLproA0n5iEEGYjdZhRD1glotea/swztH/lJuPjRWazDHV5DG9QkupLoyVIj
sq69CbyZLmf2KxhSLcc9EtT+LNtMReCqx+FzLobvYBeKAXsAblT3EXdK086p19IVEJiXkqHRn1yi
u5kjxgR8KngJ9xcU9x9NFGsvxPE1tLMfkxJL4YcFl2MlgyOlLLC8XlRUz7kft/z6BcWLGYZrol5E
nlaJYCKAKL5vzf/87XrHGInYaKeu+v1u8D48Ej1Za2MugOLgQU3kItcWXYxt2t82CNtNwPnQMwly
3uvF0cYwdykbJeDsa9Kdby3axBS7aN8CkDwdFcaYRc2Ir7wBbOZztTndenCZnYpKXHkGsWcJFCcm
aAYfbk14eVqgn0mXTFuou5uE883eqV+3mMdqCbqnPwsMdKgFZHlmpwc7gAJW8OJYX7X+Pf8lDDOM
elKIiDRtc+4OJCJ9RrJTe8P3noRoHKmCKRkR20sCRhGqmc87TkG19LEHJC2K2km6i5ord4wBQx53
S6A8wPIwcOOPZsTzEFE4kSuV534DIMvQ97dC6bQj1OBAIybWLlDoUnKgS9snYW8uJiSlUc0/inn1
4DHAIs+XfqUrHnYumaDH+L78EV/HD7m76albVS85WitjC/Lw0dRT2EfmqlDZIWz3ZXR2DniipH4A
zUO7/tilTX7LpeOb9PblsU6FhO5NbBX8/7XlULkbhQIw69glUoITNn/52jzcLIPy6aaG6YxZvIHJ
gvPnngbj4pPuN4WE/jdVYCSXxi5cbP3+mWVIzdUhRYz4J+o1FbFOKg2arsve5VCJjQfHrTQvc+tX
+jaJJyVarJIvjb0WgyYjXPgz9j2Fy1hiI8R428EJoSFjoigoF1o2PPTdMGLkw2QQF/vfnIn9OXlT
NaqhC/XjPNP4oSPWoVCx1IV/2clpSrSGDqwVyiRlPMYyJVDh1iRn5BWGvfnpd2n44dG8NbYS6J4h
YF+GVSuMT0RxyaSd/CKr7Y+7smgTewwb8E/q5+afQCGNoRsae1ty8nJjC1hlkEx8rr4XnX2A2rPC
0D5S9kkFSMbtISizPsDJ21BsuGT2HMGR/UfCYbFRdbqa5H7op1UBPl3GXi7KV1CyAHtpNYHKikJY
MKRcDPwIN/4keGBC76S5yCtMEPJ2z+Q+6zfNIpiqpHcTW21rj1cfHxnM3JVgb7gxb79jPr/vmTAb
Gmsl9PxDKZUjlH9MludkSEFbpoL8YJmRAQ/u8DknE3p3ouf5KqBwvnvq0rlVbKc0ngxRiLf0ENOq
Z5CjSMSfnRnNLHnc9GaNd8V24m1LvorsE9pJ2RW2yeaJUz5nGrFQ09BRWotU1mfCnRB4Bb9WRxf7
/EKsFub07I4SM+U0Hx7xlbzRxpXGxKAi9fmz/hkecfCWgrQYEXLBn6DxiJdQu2sVpRAnBlUw++K6
vx2a5dX6llNK96ojrYwIeB/jOaAspiST2JfVjW0BijGYp9vptpEtj5OJiE/rQUFDhy+ahRbMT04K
hrwvL/KYZuYZiYQvFgmoFPE2fTSpDpJ/j9EQ8G+6awmbuxD+Fge/7Iv27q2/5U7P6dHuxr4RPgCy
UgfcsJV06Qsw9Oec4Fkg8XCLbo/MCPqEivCeGL0gbhZYPGLbaxCzwIsQZhp9PJrGPV56WyHVvtEQ
WsI2oVxDIRqABsu1ZjoHL3HtkwvsKHR1d8wUOSNe7vDBdqsKVuvpsPOjCPUz1CISxgXIpNqmXnl1
iarf2g80yYRjXnUS3woEUcGbSv1++Tux69MB5InJ0zem7VXISnhyhydti5XkMg0Sy3LspVYWN1hE
/8liL1S+ZGzq1J8E41RtF/d6XFuK2/d9iBWtoUJ/6eWv2Wp3FoK4c4FOjLvu+TBbZecm43bmO63z
S1KlvxP9kQGM1scGqSfIa1kFTmta+NaTYaye+YyLbndkbvsbq+52hSCp3VS+CRKg1ustZsrbm11J
Pn0rLji3moQg2O30xIEboY+8sjIbY4mndUcwdXDptAKZF1r6zAPhpdCRQP6n0e+pEaxuht5zW69F
SiGiFikIGqydHtqmZ4O6+WXf5s9ixmviYj35/ND9T/CL8KiwSSnaIlaI6gUv5WVsE7p9rjc0X8yc
ykmYicbJNB5v+t3ofnsMzbHfX2or/qcxyFXbF7/n4OKFre1oIhBz3t3VjnSl1u8yfYESJWimXRjg
LCMFhuEQ3n4DmuhycS7XVX6PicyFk1/nRm3pEz6A6//rM0HBd2wkX1+47K6tgXYvF+ZXGp+dfjjL
Jy3w27k5ZT4AoxKgfMzvH8ZY4HPKMjPWmfkyF4kXxdBNeSe6QD5Jq5o4E77faG7znBQIqllXAmIa
/JV7UyhNWDNNlAbCmv/xROwshGczuxxpNOh60yWd6D6NV3JD2RT8B2Dbn+Ac4WG+eVFIy34mqTlF
ZTuqBn0j/8CV+hhJBObo7Ak5hmH5w7YY6rKxSeumEYrGQN63dIC+6Ii5VKWWJSpf7Ccqw1PRefym
2KbbQUh5Q/rhSEeGZVUthi8FYPVTnVoLfahMcT5Zh5NTlVG+zH2aQNhrfespWfoWWirL/gLzp6Tv
q0CbwFGvQ1WN+S2ryiWGZOOmhmJAmIQtPLLW7+e2YJH52oKdcR8r0enkMjL0WHrhBRep66JDAaGO
7n11+3xyiCM0MJY3YpEE5K7HBrUIxLT0GKsBdPSG8lo8b+zZOtTIlushKw0nox+vdFCO8k0iy/eb
oWU62cJBZC6meiiF/N55bXXmlDFAOpQ5X3R49m0NdKj/SGsA+wu1MonhJNIqjJRpmn7tH0DlrTIG
P/AsNu3L4tdbyZPuFWCJEwXM8B9uOEf89z68L2WIn37v5G4Ug3+PS9Ayv5BYN5sxO+oJCYKVbAaI
4z+NCTJJpTG7I7DDS08C9SIBm8kwRE9XQpZ38QionAxfL9RYS7pkhmzYEsaCuSLUiout01tQ7thd
hJIsFK+gn2ahO8j6rlpYvG82c+gYkgNIjQC99aEP3rdo33FAItMpW111xS3ZzBx6Km8ejQj2rVdJ
clqRblSAH+sCVItir9Zp4XHB/J0cXe7PCLT4XIt06pDLBEkh4QQbK3H3y3lj6VTD2aEGlzhCjKfM
8juXmzpmRsqi39pKe0oDfnRkEhiHjeJfyzF5vWfoKYVAuwOv1Ta5XOlbBX9lBsoxTQ/rhc3QxuJE
lAx6CEz5cfwuHMbLpZvA45md8q8a9aN0L7uaqzcc3Dq40Qjcb3vR6yRZ9DD/1/nutcEDIs9yPiLa
bRRigtOEMScPCrQ62ixiDJt8rPvcqTSHOaUYgfrJYTx7AaB3HoZ7nxVW0NPnAo2yyjfLaJZoNp6W
ydbhzAFk2eGK7qM/MmJvdhJ4ypBS3zQnoTsQnuPsJpBm43o3jdOdgQmv0Q5n+try4/29qjTLoCv1
WpDY/ah2OGtah0aVYCswz+LI6m6vizG0yXTCu2b8jVju7I+hQyRm16EsrfodJe5aw2GtDDXWVsaO
fEDE2JRWBer8HH2aSnvU5DiEpgQJlOqPEJDDUqWGA9dfm+RZjxzgVITLnAf6OxW2LkvnTZCYXi9W
yxTuv9scR3BwlffDCgKpshRhbDhlSO15/H9KVm2Q1xrcdzvGRRKwcnq3xXaMm4izcsBq9wMyyjUj
FrLhQqwoh/Y7bstiroHehlijZn0o/DMg7/cKV4Oa/e+UrmG58jgnXGryBAgWCyVqAPqJ2Q3ewiXH
efhYG7P4/E2qznDr3VU1bc8HmjO9hFJ3nDZEjP0PvRj6OH1qWthUF+TTWSlg21oqy1QTHozKZ8pd
PWdrqp+xSIw2KmpzlaXcrnYjBAvOUz0DiOLtcf5Lioneg5McGeuifIrrcamzXSaevuPfr7bpZEW4
+7wTMCt4QR20LxQABJkS9tZO0zChuSqnaS4FMcZVvuYF2yKi1rVPVljuQ9uTQUrQQYwdAm5pYGM0
q6lNktSgN3jjExMnxST15cFgy3smvRA/YFPHDsp+r2NxNLwxuliEwGfh6vGfcBboRV+v7D6+4gUr
lzC1+SqO2AxP9tN/Zgo0oEC/GwyyI45/eEcosujLRcBHMQso82yajVskM+mWB+7da4LMzAQZC0D+
k1Ewx5/Kp2BUqZaDdKRakERQX0aqBHTYjLxT1GIWulWtg+Eb3oChGAGc+AqCGr1Lm1HrUksm/D/+
O821jabvWegmjSKGI//XHqS353O9IVrXSr8C73YtS53Ojqw2syj+5oUO0+FShPWn16y2hWzSRhS9
lvyvi+piOf8ycsqIEnpQMuyk4z9QmhyGPlynvNjtaJywyiXz/JSDuLcXaLxTlbQ/Xq/pu5FBr8RX
ENkFqzJ1g7D8beNhlV5lc5a5JLG75+xkyxD8/ezFPlJYAaf04VOv0fI0p8YD6CN2FDYaqUc8JCfL
Ym8ktgjZ1Ss2CLYTqfRB+rvVqoa9eD8eG8GYOlg3L7LCOghanSkPxYlY4xIlLgunxtVKfq7hOXei
KaX+9olSrTB0KJBcR/aUZVNvEhhhmm8U9fwRXC6lJTW3lp6o5acWFEScA+kmJtKIOfWmSHbSNcYq
2X6Jsj2FLNXBdccEjn6RTrt/2Q/cflPpFqZZuw2g0LeClNpO4VLreNv0YvIcr8GPzFdU2ZK3CzN5
sm2SDZ7jWysxuVnGKMVt56OX2EvgkWmfAXffnPex5VtXhdtk6M8uFDHirQJsG+TQ8JXdCMDg4EIY
y/19Eh2xXmf7RcmldZRzc9Hx+2lsqpG7w67vsg/nLXL8mQHZBaibLhLIRwrehJsL4mAUcFARbEg4
aFLyccDAXf/ubwtcBjMeOw8YibzFz82QiWESptcTpUgq2GTP9B5fiUXTurkrVCPzOU/5kIG2GK/k
4K2SxF48GDkWGKKPUEKUWcAHHfyaKvx1ikpaS+4cVv/U3YCz0N0d4/1YeKTuJQ6Lhrmx/uXfq5mp
2ufaYXQc+CvEeC/Xeuh0yygLUJE73Ii/QYoy/CdF8eXER8pOLZedsd+o8r9CsG3uMvZJ161yEZJM
Vv42cnLp23m4PjYzZolEZwssgZxfZSOaIxwe88Rro2GqxVSyKZAZW5x9S1Lwbt3e/3yEmBO7AEgQ
M4cVc1V3mEsXw1sxdyu/Ln8wGBjOx0Bk/Xg6vXdz1BMNDxuS8gUbQasnSl0V0GHGIwgftsUdCMOz
4plwkApiQDwZT8j3OUUvGJurWAfnolRJxyrFPaZ9l99rZnghVGDZwihMEoDIwoxYUgRyZpDwse+G
LBN9PEdxxgdjn9lEOI5pnZEfSJMv32msbVbKrj1N9hyWic4eftHgoPNe6fQ2GPz9zaGhY8m1WGHN
tvMcj0TgV5zyUDSPEvxlBQ+pN411CEhDJDd54mN/LV4ZC3hGECWK8bLjbfDbcvbntq3DjJVqaq9C
jcxqBEIIdkFSRuVMIuLJbCwXZBdzqaw4vP3yAON6vIeXw3o3IIGABatzgZpXIdBYeUCYfumgO+Kk
o+G7YtnVEsN5QyjgtA1azI5WGYPT+6jm+Jb+QScmAEzHtDT+4OhwqmmxKV10FWqkgfghanG6waXV
9FxG5+eUz+XSmZ8m3cNTiYdl7IC4//do3zT3eMtUjxAKv/7F4NuZnQ3l7l+huAEXnx/mRm5E597v
NCmcamANn7qC6F9AmgzN8TQ0CVK2hef71LHJvfXx8I98Pno3XAsjf4bZrHZ5YhZRliqKHyltFzFc
xuRx4MndbVCidOO4ji2vtlNab/yVb1SHs4seRg+hwkpHGqIj/UGz0LIueqmKrD1xvaHQnueUaGvE
rG6/2orqYriwLNLABQY6Mh7Hzi7mnokQ9TuvGl9s/PhQQx4GCb/YeiusSvJP96MokF5jENQJQFrf
LuHgapuNvA6ZdmwhP7ujz0DptL+qYOM0m0CXjrEnU/qiMOJ3Ub9oLVu4qa+FSwztfpiFSPxbPntL
kuYVOxrmNHoXCizZ2Wbq2sNFugyier72IPHBlFCzgTYjzDxUZo51bHBQKtDO023xvI0yAg0a09Lu
hHHbpWouHiAyA7RMuPrr/ph5hUAMxaJy01hB8w/g7sXTJ07I4b6ephlLw8qFySoADW3W8QOPAUUx
yQfdfXtnjUSTnsfULSuS79WTmWmM2/QERupNVYXjOnMcvFxXkLv/h2AkxawLjuDQr9b7kdG+KN19
kw0vnRk4AzYkjPFWiUYcjzHtKIDm49XACWy0DISljN1LgW5SVymSTBALWMceEXXGIQklyq49xvph
uxQnpCnMP4K1I5HungO39VEnECzktoy55dmIjet6iPGTUC1tuHn2bEJ5Q6tt0xhzok7lB+V9N5kc
DSNUE6/tYW348xM/BGT+C5vv9ELhPWrh86xBaBH2uLuPQhWF505ioBTLVRpFBD7o+//EnVtOoDIL
rObCb15hpVI7tzRqPUYQd2LoGdm9Cj67LaKerP/Bhc92DNZNcUKU0v/DHOKCz3IlXbtAf3STcD44
H5VA2KihfdmlZR0UjtH/T43sUPJzi8newUONl5qL1+Cnta0ki++7onXeTduWtQXQ7qscueRYuMRs
oElDL+dnJEEpML0M4tNKQKdD4qYb04DgK5pQgDWYA3V++ocdNEKkmSFof7ZJhrllHhwFzjvD7esh
3f1ooaXXGC+Gxozr8eCrjwp3WPbEunkSjwbA2bLX6r7VFbJTirKbA5VGunRCmncDGX4KfrViFPuC
KO+J2a/nYwYXBF62IrVsBYXCU/3x75qT0kVjd1mrAGsT9OJJB95HlaOp7EstJ1pSWW0IJQ7XYLiN
8p8XoXJRgtM62umD9h3hyB4LoCz3QRbSc3Q2aSXk7bo043sjH6G6Pqc9YLHCYdjaZhT+KlDP7IWC
NmqpcbjccAXPxAlcTjFgxuOxrAP2esuWFSnxiBLKFmwQqrid+jFK62QcVRFPOtzBpmgRQfBSnXcS
g1l92BTi3qnSN3cI6tT9si0eVXy9pvbUPDjk2+2/VkHIbbK3tfBL6vnp74Gh4dqYilgP1oKGTWYb
8hOuyZVUP6q2lcnr7eS53AlN+YqOm+abC2KP+vTX/NU5FRxsNxkB73SFfs+ukZiCMnEYsInYT6Je
bE8DfKxQJKSzdArWt9c6MqDooj9fBuy6dUjrCBwU77H2FdDLL37JRjvGNjMXsPiw9brRX5/o48qt
7TTsY7zVR7TUxA/EQQSdHD3JROVYVQkrlKsG8ejo0sgsLkqc2FMHfTSy1kLoOAMdbKV7sB+WJp1U
9ne5qfKW/o87NAHgE7Nl9rPY/+Vk7GbuvgkQoJhnN8q1L6wz5a0TE62qGWvcSBxeiwVREWAV1zXv
ocA0hMCs+UdaAQ+Rq5ZCOjyBGSu2A+VNAImz8dOo/BiWAcG9wSHyPL6vKT/adwhVJElxBaIIRKOR
7TNnpHvAYhooF5g+EJPasmTYbEJYr+d8H769CFOU5BeorqGcBaPvA8wSrDDk63Tl7EC0VTEPaE5j
gqaxjGHEsochAtzh4BpDwV8//BOf7AtS3f7IW6EesnTMcFTjtZQ2ZsQ8rmFylkjP7KnQKV4f1Koq
XTFoXewo3UYZseyC4kKT8SHN9+6wbO2qqXxwgnAaBek3hABE3tznFtOPOx0D2dhb1skmdhA80+Fc
MmbtbWp5QVYPInLCN2qGZmn9VWiKGQ3q2Y5LRpvKMD6CPIpdhcZWshCGiT3syd6ZFFcnWeu9fPhN
1WqchDptdUuKYf2Z0iG4WnOChPUydkvPcUbwy8q5s0Dp0nPvp7o3FgfRXE+zc9zsxQOR6BSE8Ct2
HEpgudFPiZ0xVmCEq610vCxhoWnb9iyLekuCQNkTTAPfyAkLsEw9Uw3Yeh+lPIs08ecRH8/FcYsu
jag40TFDZFfnAAvnvzx6DdjPHq6gOOMpMXXpIR1cXRd7SLkFVlOowatMl5PSkgf7vwO2/Ux+LxCE
r06RWKps87uEez91zRJd7DT4WlAhZdCVkVm+KwkQFdJQIHlZS8x9xuNg7yML3eVmmxZqKqSf/0Kq
gd4upcEX3mx0iYxAjT8fjiOPpCZxKZX0sr3L/DR6BECBId7Em2f9nydcl1Zrbw3N91LXww+efRfA
9/EAoe+qMta8LeIDpUMK/bRLfE4Y0R/J39QqE6ccMcgFCGe9/665VKubDtHYi6oLYws/eYzqY2FC
45Jy1ObdVsguHV/NpSnzRPvOMAbB7Vtr/HknNMCNj2bTgBrIK8JX/faYd6SN7T9I4dQVhsEIjbLS
SGAcObgnwDSFeJYkeR3RLiBdEui5hmRstCLfQ9F5Q0fD4EOVccN5nVrfg/4i8DTqr15VANWPr2xX
iKlKo4ZoSi89K+c8CX6dwD1j8Df+GkXEuPbr1x5Jn7AFPIEb858TIoP5xZHFDjQW/VCUdRRfjxQ+
4emIJLEFwLqeamzXf0vRhXKHRRarCHi6nKALa8Rtk4riqHJYwaLEV2RWLxmOo91/ulvByifzzvl4
ogpLDU3gBWdfKjrFswAUbjN1ax0d6Z57fo1s1A2diyhp04ZGyCefDXt6R+ABUIZTTNqGBzRYheTt
CwfAhOT1YPJm3J+gCfWFJJIIK1yEo6ACqwA3DqiQzz/ZGOrD1lTOXVe7kZG8hJeyCX6p1T8+sO9R
mNF/LGkExQ+ciStCis9SscDR0NLMLDli8WuOb5RefoR4pItZPmq3uI5rGEYe8ibplOEqweW0Xmfa
POQmeVXYrDlpPX+RCNHC18cxs5QfJ8tizmJVKApuWPLyMNEiYMaGXwo8hXQW3zTwZJGen/zvxUyq
KmWkS/pcr0P5K687jbpLq72eEcwup3S3U1ldnycc1lqmunR8I7jD1RqtVMhi5ljBcew2svLXkbUa
9peW0iiT7CZVcjRA0rigIx+aQwA20CxVBJBkabiNmpM3acubGuLxogfkhuUna3ZJRoVeTKI2+QUC
lMNINuMJrjLX00AcKPDohzUabH7WdgSs1qlKEoudj/bVdgjWSRD5SyhlicOX7qYnMk9VaOzgqZu9
vNhXAUxsfdkbCdX8RNLFeRxEr/8WQw4TMBfTed+UcImW178CKppdNB6q3RLahXMGwCWo8FiU3BIn
fCYNlfG6lhTI/gv1sWJsuWo8KzskfWpRupcFeMjdhtmm0Aabuo22gmLhPjv46fvW6abWWM+xd7UQ
BuC0SE9i48ZUwY2e1HsYJKFsCguNSL85OSfvPAVc7nW8kW1pkhMiPZRnQuEQmSUvat6VZk5eWDPY
g9xGyXkYGaH9LGQmVoOgJC9lAj0KHDoLTlzW9PknnldR+oBYS4Q5gB7n9GYUkl0Cfa3MatlSEQf7
BNsdS5r0VEFSTutuNrLW4k7zv8a2mY3LukbTHduGuUqPCn+Kg0XMX2tRYL4UVmSrOg+jt+hEtxWG
GoGY+OtPPC54z3mqncEwZfIPPbffVLL+kstcqCM3bx8XNIwxEAFFaRUXU0viqP8hNoKZIvINsWa7
42hTDXho+pZS7/taQyiouIhYy46UgvcukqlQ+EkjkbyRuv0TjTkddTdjUjuFk03uxsd+lu/K2cUK
kSo8o+BsKx9feEXGKmWLkrc0eHVt6ZkiLa75hkr1IScA4n0Sm1AFHhoDfv2nr2TVhbWNcDgM8JA6
Dl64YF+siICpN1EE0/+oXjka94zNJrnCNRkWBR251A/clTG1C28tVreqZyIyG8jITNfOvsVIi9U7
TWB7tj20Brng1+kfFI8ryP4sLQCjdQaKNGNLBS/FJ2cGJETVC/omLh39eY5s5kSgJL7rxUoq+52S
oQ9BnHeiz37jm+fX6xz6/ZEv34iZE6ai5GOUKKFdcLiGdnKrvW129RK9I/8J4DyoVouoTVmwvDPJ
XjmAcchSqTJoQ4EOtx1kfwKIq6wzbig0AUYoZoov6D2C/ADiNT3/kj+bho3hjlrzXF8hhWnZlcha
r/jlVnS2WSj7jFPwcOS2kiPAko4HVMt3cWiuroUerMiZZAdmWY4nRsUlJ8qpbv/sp97aMtva0r0p
o/AUiwhLx6PVQ5wDU+jDFjpHWv4kV4w843Dcf9xGdiqaeW+6Gmkf+vEguMSI3r112srJiQAXqq12
yP0AYA/Cs01EikesFL4EFMdK5hD3V2q236PakQfEf4g842I3iRykVzhjo0ahSC3KfIqqxJqO8Nx9
To516Rsjb7CZwC5zzCflgdSkvQRROMF1HCEcIJUMVBonoEJjiZDcpEdjiAZb98mVqZV1DhMqQDjg
WEWQul6JMjtgJISQVh/A15kbGVi58bDtzj4F7vLcDX9Ju04/s/xjGfu2gZyOzpRUVodZvvl/6QXR
pGKNzuLrLTLi2ZWp4YqxEqwebcd1zwN3UjdQPtPMKdsk1DMoIpN9IGZXM6N90NRVfJljBiQWQs78
Sx2uLd7fExfEdfAw/S7AtSeoXVJk0CbAwPaPLq6SjUozv9JYEXzLCB3zVaT0InRIH+uKCYmnc4qo
c9/QEUTdTw23lybMsEbM3yODH+4bnS+yhZhA93yaHp6sH3wWy0RqWqqpCZLYs6lJpETsp91j982Z
rL7SgY44rAYviBmJpiId64/Tzd2C6sW9mMNhe2E2uMpFae+Y2ALku+AqYKusQGMJQBofA76WET0E
8Ob+ZlD26TunykPqk83oSF1M7CNOKB5fapvrjywB3+8qFBmfCzQG4MofEPl/SGhOdobeGfo72S+l
MUH98Mk5dAshAC2sk2hQrqBhe2nxN+c9O+QMR6QueMYbPAWJEhTQAIEE0Ts+0liEzznhHY69yMbX
P22oS0Kf23M7Kr/WDRcNRNBq6m38gnnE6Bu4i++uczgzB0CDVO++gHh/GL+icg1TLs+vQqlFNmIZ
TLxboDYE5xj2kLOAG0i4gJvCLXszkLIA5VkyEXjSxvbHkXy4LTgdshHMOeWNv9RX+7mYd2KBOwup
EVufQEk7dk5kY2jp29jCzSW+kRw1EZfyxByB0G/LACbaSQaIyVgldbR4/cT0buwC8gYygE92DbEa
Egt3/vNBNwcYMncfq3pws9TIOpjBYHWcXcays0pOyXiFVKAho/IH0i3nGdSrh+r9DrDFiTvWk/KL
XKjU3f+dUiOgmz9ZOIvEfTj01nsc4yRQx18zEOUCs3we/FezXyHalj1nwXUgA48DzIG3JQPW4/HK
WnKnDq/CtyI9UhOm6jnkCJXqsE6zopltmFrp8tuaXC1sNYsNMVWTL+ugHQz7ULFY9IkGCkk0pXOg
XWZt2XQEVjyRlmZaFIy/enp4xccgl9FyEUfTO12yszXP567/XqGzzldjNBgJO0J6G4nNAttk53aT
CmSMszFVe3rHmkSKsgkpkJ2Hp9v8PYgv3fmXB65V8FJoytAMn+ILvV6MAbTZLkK8Yn8wKgNvY//D
3XvsVJ/X41bh8myHycnyVyzrBzW7y7S4Cvbcawuf6Z1tA+XFNztMUG/hPJKJDshir0o4TS5miahL
54eXQ1M/z4tAlnZOJaMEBaxt9LfSDvpO98Q/F2Jn02msJUgGGY5P0/t3Aej+rpd4ll8IdsJyS4ME
FkUfm7BtpVMlFLwhRyi6abFfL9YJxgBzVe/vEQ6ArIBclu+w2cM4ltDAIC5fR2ulCmEh6///JHaS
bBzLm1zfaXzKEFmf5L+bsKtVI2vTTDk+XyRuRxG83s31CvOml+0hA7SFdFt+YuamSyO+xvdrHIpl
HTnzIgqUvovK6B6T8nYHRk5fJR8NlRlIhYlxBj92/yyyN3MY4bhWStvuMTizelDSKwcd7dM4bv3/
hSYOJ77Ip32fqzd5MjbpaCWBIsSSIqZTi990JsUgVVzY1m6LvXcFu0fh/ea0Kcl2gIj1hz/+jqUo
rEDAdGaVANamwvy2mgJ/VPtkeLzY08jdczyOZer95L81pw3WC16x5wEJQon77JRnoGJVS2lo0SHz
5nq9Kiene6wVrtZ+cuVOwahoV+e0eWHNU1HkE5ChSagIRMavb6J/6ZTkmz8A+ynw5WJQ6/fpQMNH
K6G8BJtfqxqlw+h80vNZt+1kdTvH4ipebgDD6DMGoPUHWCJfBJCIh9yiT1d49AO4dBoWS+kzJ+VY
/2Ge9O8vOEYxllqglMeub+Njwt3HEhFBwdnJ8l4FG/ula+XZvs3YuU1dejn1v9GJO7Z3+hV9KVqv
H+P1P3cIFHIFYTHvIV0juM4/thmKE/KQ2eQLXv6OyqPs5IcxRmGYi2t4gyQ+QIKWMUlb7Q04hylz
u1wVKKU+urSwArRBKEOwXf71qFRD+ZQf91HoVJRBF5iRJuHXxtzghUTAyKJcRPOxMnjU8sstJA3s
4/+Khxz+DXeprje9p9p6+eTVtaTp/u19LOD6o5kAEbJ0yVmTgiCFENjdKfKW8DugozdhiQVRFUcS
wh/HYNJdzU6MR333qjJjlzYxdnu77gQuYZxWBWG4IZfIvavVz2GFHBoKdYqhVbN8xhaM1QSClH4t
RZZl+XpQ09zpJrUt3e+UO8T7fDRngVpqGFZRBkM32QWSOoKmI5J7FuLDuwZVZPesqjDfsivIyQXN
bLKXwrxEALK6Ya99gVWFbXWeLfU7FDXRu7t9EBULtSsNawgQO+SS3bSx2neTqRQ6LLhQ7i6Og4nS
yOwd0KKxUisJT6A0418FiZL2g+ZxD+DEqBKdf6+gH59iWUY1CEV7rf685ClWkFyLieZNjEcjd9Rt
/AaGnDgh5R2KRBX1UQUfugHuw41DZ7drMbenddXzDT/gTJo/eRoNWy0bZzXuhlbl6a4iYXxC4Io3
rxP0iXB0/oBz4DAVqmsWxuJKwr1Bg7+cUlMeA4kqRuEJ3UNU2sJZbsDUVNPdAtANLul886g/Yvs9
VEPKZvzoBCYHRoz+bYMx8kPC4KQzlPlmH2pTbm0+QZu/6C7zfyiPnvASRKDZhPmB2TYCtiXw7xKb
Qf7ZC8tChya3fo8TWSx0oisDZA62LyBIY2wx7dOYW/sM9OPr7qrCgz0ObCzCDoLlhdNZGFx0PR3v
hqZBKwupKas8QUXO4BePP+FI0eyEGhS9CEfzSBqgPTspNDwmiO1h09CwcwS5WbI3FPw6iTxNCHiu
fNbKVDCZ4UkDsw/l9q18mjIp22NmTGS2Lm8w8vdJLhOUgLroAypCLg7/PhhNG9jA/5FlwNFZtSFk
QcmCvgdo1fZ/Jk2j+Db33tOIRMixPEksDph8sPlQdT1kwlVwvi3hf9ntX3LHrSERNqc8s27MP3xE
hvtsky25A5n+8glbdUVXuQYhvTyZeuYX1SZ9GhV8UdekAqs8rJvcMzqWsu+EdXe1mc12KKSYmBFL
IkT5MS02+DOHq8to6W+8z3Qw4Lps7IVqobPH8D5DV/pUHawhc3KYj2XaavLs9jJgzaQ85OWn5D8t
YMyicNo/wWqOsW2zRNUHV4dQSQcFjahw12+VggJMTHdAVhWO48LWnUTG7SnXcit2/85fuSvJ1KZR
qj5zJLC9OwvenqR3xnS49DJfrTMDlOKILfRe74xnWPOZFytQItNric9E1ynXew0osPjP6u5ltxnx
OnHIgaSKqIqMnZWHyF0mR2VvwNm22CskjROeSQMH5mIlCKGXHz91qMIyCQVmmTOo5J66Gw4c7vXx
vzkHYu0WOpj522qIJCCj9s1GF0/dhN+CknWpGjFI/tcIOYSpUJ7fvh16yD8k+1fI1m4QBGEV3Qxo
4egSvKFtfeqHxnJefuqiwB/MY2dD9nHSnh9cYe/hlkFe2n3AG9p/Se35+1+uyiBhirz6/6zU6FLL
yaSzzmSGgja/7UmBf0B6dUtwzQN5let2IoxxUGuTakYNczjN10Z+VsHm0DHGBzzeaSpVjUcD6E0r
JcGnSGyEAkaI9zWks7JaQkuF5qJigR978rIWEp2CVxiSRIkxmF3/YjqSEmA173uIeoARv2Ln2T1H
/K2r/UCrGFkPmEpM6YOVi0qL45iBa6zpr2S5ZiZd3jPRWTINapaZ4Gea1NG2UQU5oivhiabrIMh2
VscEMhC8wJk+N8082A7OGK2Pgz9MUOXQ70FxnhAXh8KETqskOMOwyuAn2dOb7Zuahh3kyd8bE9KO
+ZkoIPJT78T/XSYPYTuG9MA/EqrHqdyhbXMVKND6k0MlXSyYq50Ac1g/tl9vHrm2UPGQRFUzCQxt
1wMcesUzAuBfLSimkogVTWDWgnFVjG2TNHgt7c2Bcuvz+F2I0k+XcToLwPFGgkIoufCCrG6utrx9
ChxJ/pZyztZGVjIgdkD0SkTjiEzYzi3ZJGTZ4IuQ0JeGdTvnqDspY2n5wJiJoE1sevnHiMBtA/+c
lQRiMmAvMXiKeLR5kd2DFK5rSTOmdFhX2QElhQWmMb1hgwujoHgYUqSdJEMqbylJPwsb3isas+XY
TxlG2ltSypGXpFGW3k82m2Ef2zgIVLjFvpuRtQXMinZYuU4hMo4ZK6EyadS+gCoR39jKs+dkYOTn
tKRLe9MqoLv3I8752FpW7CiTenD9nVLnzVkbms3NQHMm1rplxqNFQn17XiuDgrBgLBx0rKMrsWD3
kkFxBJHMH+6GJut8GAUQOPR4Yx2ij5DG8XmjM41vBy7Kqe0AATTTyoqPVOWOL0peH1bygbsJCXeq
+XCr3VhYnYZeUQoPxjGFCeVPOXWVlyNSa+wgrG8DpbYjxoCDPi9KHFGO1MmSzBwBziVHCZJ+NJdh
cQ6JB5nb2Vv5yi4EqiHwtmcb0R+bxpegVnBL/njOadod6V9VzIIJZzFT4kIXqktITlGDewZqa1oB
wHGC+y85z5AnOzzSJlAr9HqB+P5SL2nYeGtzkgXRgpyHk7BXLv3M2ljW2DDXrlZCbK03lVr/UPgL
rOCSPSCG0e213wFF5H/ktUqDUwc6CBUXjnEviBrdVlYCXLHdUZApgpTkg3JIgPBvJgXKyljdnebG
22KNx9oMF69Ent0Rs6PprzNVHa11xFMaouvJIoW0kb40/giF8wmF9Cww3gtL4D6eo4AcdMM4VCtN
H1moJQPwhSJ5M5RfbTpJr2112mGyHZZ2qkz4KAhek/3fDafMHsa8aNSK+4qFSMwsfjxsI2TU+SkQ
mN6VSVU0NNahoSVbAqM712GfEp1nC3foiMXhLfmIo4yBTvMHgTrGgGQizgkTKcVbdGMYDrEKDdH7
QocyoH8HkjDewLuFZHZUmz9au6DVPmOt2c3jd6NWps9bYkfjTRdWXPtpgeDchOIV7TzbiI2u6BU4
UaTgXZZ6PVy/nMS2b7sa5Xlg6VnCFOKCMT5ZoU+m2Db6IQFEqDOKKT0BkIuc9hdJgrrefpoN4Zz7
8Bmoz7QUBWJyInwU7XnkgcpDnRZn8nSGYa25cVG4zsPg2IzAua6uvpGcUPxmg8VwwcwCDH4E5kKh
hOiocuD94sRAqxutHrzZZNjTccPTwrvNos/nqq9/pbsWxxAy3ms8pEtpV+/kbg53g5fo7w6WVyYK
+huTRJsKvtYV1qfXq+Z3TkkI93XuAdsXDsv19QbxgeJ1Ned8KJnW/Przzs4OE0bv7JiWsKYQHupu
/82i6lCzqKIvcafy0BApD+oeTjxLS/VGIn6EX7tXTUCe9xMxsDMVbooyV7f7lBWxyO8v4Nw0AdTB
r+BVJNiJj7lifyzH0FbHd2CD1wN8YuaifKSFhs+Rq/gQTbkTpCWCY8vc7vvOSJKijq3xubEoSEYy
2fROfL1wGFS6E6ZMZT84/eaGJlaXo7+65dvxHBjCS5jl+eHBMMnxenm6NrtlAhlu56i+bou5Hiea
wFz4QIgLgtFGa7YgyHDTXqvPA3JV4txt52pA7CYko+9hP58ut+A/5BEBInLFSNuAcNovPhwb1W3B
ykOj0RksfQfTXIPwd9SYkreqBuHvHVVd7ITQxj/3GZ2EgRalnpZbFEu/IF6MtuxOJzLdIxxaF54/
/pTdFI+gd4Xux1e6SmbiYgQDM9T553jGhJf+nIqP8bie0EQgS3xXyRgVNOBupPdSzdi+GoyGuq3l
zMtFnvvZUXjYv60mjqNfaQOJDYugqxXZDJddbkVzSmQfiAvdazBRVWYvKmCiKfTsMDFB8h0SAoX6
rauVTp/NaVCM491wJH5ES5kvbQrvtNugZ41gFE8/nl4vQKhq0gg2aOiEsjKb7j+cTZ92PxRSghoz
1qCOsW+B2krHQxo+x3JB1cDmqvBLv3JBBOfIGVAcaF3PD5YB7/uYrdCz1weqV9SAUQXTv8pQOo+s
Bxw3GlCrZP/yrX/5ahWa7OzeaV1faE4wyc+9VcIlXQHxn5Jc71Np/hLnMQdIt2uBKEi46KzoM9Yj
S22QynLMVy3AA9tsgS7CcCui9ShByKsm8VvloXLJGXYUCdC2fsSuWYCl+goZLJD0qIzERCwv+7z2
lBK0SPXX8w4env/UYs1CsaZTJKUQHoAhhrWBz+ZCTR5ehf2xnArYUnltw+t7SwAZzpjArach4FaW
2PN3+RwsF3ZABIppQprXiGGq0TzrjpAdOBOINKSiE5dRBAbaXnvxZrJ8M+9AT5VE524pEV2evCSE
lKJ9LSu4LJiY+00Nj45VH4NwzcGZ9JeG1S3feCPucsJRFH9xgV663dzekUgBd0tgZX0Zgnyc6bXz
uORmLktG5A8pt1Uv0wWmYKJ5rasu5jRD9KKGbj5fqyDD88cijTx2U57cAv2l5sx6+pt6I+FyKGik
wGpebq76ys0npYcGaT2VRRsoy/3d9H9oZAvHSKXJvEDyWLb63xBZpn4XARFdJUgxxza097a4uep/
kUt5/ctI5S6P2TUqNfqpnOozYJORd5ygVvkcVuBIYxk0dCUdBbcdD0ElLjmil6bWHJmsk+H2S9cg
bcPkVqJL8aPUp8PhUJRctgauOKhUG3OvZJQSIpwdpetUgqu+CeVikkhRy31UIqlMBgHmQn7kWOE0
LvWZ4AF3BlaXeeuvgWMkRHY0SZcj01uqn/eszAmqG5NeyqCayfQvMA6kbpiqWxYGO+UepUedKegk
Uonr7XuM2hml2u0KRu7QsCFpHbemqA1Tx7AcMdRTYPF5RtfQr7504HIlBIcmnuJLBbRcI5NPRmqX
RE3QaULsL7SXbcVlHMaYU2Sh2kkU7/LRl+1B35nXPquP8fgyC7XV2zzRCjsRY8IOLF2M1HtJUtLD
AV6edQzqSbl/rGbzK4MtQK+pfjSdp3eK5wK4sLRME2Q5jeMGdj2zKcoaszksWidhPT7BWb7UozXk
vIr+96A4uKd9INcXCuv6yBziYqLxK2UIQjbR/VWdYOkxbb3j4B6FcshO6BAf87CaviLBZmXZwQcW
KUlbTpIn1TK50pWgwCM0q9ElwbXv+4gtD+UwcsO6FcR2nqNV+UjBtI7NfZi8wJKarSQiOTcJHVTs
nB/vlyTSGnFNx52siAFpiIrRUYCplvvzt8N9ZlB7L3ktBjwWmIr5YDO3p/DIPyaDqKKEelJjtoVH
tQpAEH7v8JjDyj5KsII6y46KRE92oEzaksWk34S7TrNA+C+cbSh0t5djrWD17A2F/A6/GS1czbe1
YQJqfNurIukwKSYjIf4/Yk7cCMyfWobPnF8ei3hT9HSuMx6lcPWASO1gU79eYo21JXcR1jzCP/1E
IC3AnVt82cUqYYehrKSZc6u88pjl8DqWhy7XwXOnIWK2QjiZGeNoM8+q4GJwhnjx02e+8/0tjnwI
URm+M+pNA9u7GBedOQqkHHEs/Tg5x9lv+DNAQ3VPAQxRp/NUI2CcNZvly/8o3GBnANb5VrEqsgjB
jQI/Xxc5mF56MPOraMor1ODp6gZUvZC+FHPlOOuGC8gNDfICimvuaT4G5P54cyjT2NYqGi/G1R/Z
wJDe7HmX85lLGgqvgvFZNu4qcWUgCT1IPyN71M1IWiejA3xwTGvTvBVZbWsonobWsxq8oXFDt3Pp
SO7YERCoCbBLmNZNppyy9hYytEDp0GpZbGuR+mfEfHI99FT+wIvDBaFQ50D/oY+tYBmRSImc8tDi
Gq3UhXdVcLE8mys0R8p7UaXw81sNznOZFUtM65R9VZu2Wx1cBiXaO3+AC/cEMCa6WxzEK/jZrdP0
Fwl3d90WvJeGqhaeUWX6ZXtseU6XTxPXcabMaCXoYq6gYLBJ3KnqCoVXJkVBpnr7+t00qxyMjGiL
1cHCYtXYOpsFr2tjQkJIJSwWbbHuwuJuPXh9pViQRbHkpsH6qacP3nxfu6e9JAaa6aXTrz6we8gL
y+u4XGkG4suVH13nBJyuJKZGZL2u9vqnArxrqk3NtCqoloOVemqhlYjO0RjoXHw8+7GgYh6DrWKE
12l6KAGthSdVaEuSr+m/x0WJ2JJLRZSil/cQ5vUPdhXsHaMsd4iWKGdYgf1qhjL08KyCr9N/rIDT
ee/fXR7I0RbYWnpGFbUsXvREDiN6pyxNzcGSHxEmQnES00r0FdGRrka9+GDCBDPRi2Rhwsbhec9N
Lz7jHqqvs5H4g2jlLVpHoFYuomVZ/W8ETb7tL7Jepc+ylmSAwPFiyuSwchslcv7zUFcPVTSh+qPj
G6t3MQtz6w6C8IWxyII1PhughOvzBcanXtiSzmweUZji0NVv2EbdkdyhOefNQ47Ne+yrrZGSChSI
PR2GLC6Rmz4fclue0QN5zxJbE+2xs/uwpGZnKsx5OOEBSKwDuC2/xMdriWKrz75ZpVGvQpMUnnIC
LJ/PHDifV/dOeCSl8MUy0t0vgJzgQBFUW+D9zqQzDIQE/jfkAcNWu0raI3kQB1hRfsnwpTxFDuFf
tqq3DzJcsN2TiNuwb+aYy3W8hivv25bRxVP5DmRUgfzWKFENr0ODhcWwOs9eGzvTBIeXQH1FtBDl
Mg4mlbZosILQaKVOnD0BekQ98G//SzkzH4lYjwaj4Acx84xg+xwEdLTpvP7+uQzs3gGNyzKq/UfX
IO9w3W34h87pszOLFP1yi+8eSbSuHqEGPaSAzECU3h05FSDq8gDbnGT0m+tMZp6VpLUJbOZKjc+G
In0sQDx9ZYPyHVp6o052OQzoC5TxDgUb9IMvZbfc2DJkqEaWffc+sV+yGYLB3bGBqm2MbLpkygLx
ViLb/MOP/eewqTHdbJqdrYpx8rbXP3R3z+zcCfWa6jJNu0aQBzpo59rZg6Usarqrl6CzBrV9TNaR
uB5kbuc1iNaxEO0lBH1VXPL80DC1iNmPnuY0BGPA3xJ81EhRPh173xQKzcsnjmddR1lRK0/YW0yr
riXtrshjJwTiVY8bDu3Id0YzMoTjUOVQnb+kLqPo2oM+dWeb+lLW5UtNLr8FWF798SKKZ8IZTHEa
pSA+7KAaHRktn/isanwABi+wyIkW/YXRCgt4+3YaY2iM7QgUlrZ5k3YawzoptzX4je6AxPVxjs4M
SWW39Wwc61GWm6KQ6SooQR0Vv2593kZrJY/WIVbOsNhxzl2Ct2V0nl3doWsYVsWTKeJB2XCYNk6h
mCD2TCnDVaRyPkTv1+kduC6TJbFnsuDLmYG34EjqoKf7XfP9PtewF9mHFgCP9cdDpFJ/ekAh8P6c
hMSy26x6MjBH8NSG3yuJwVQ7BEJOXCz98T9AVvlH4JrmPv3SnbPepZlpAftEK81/akBCnkayC12c
PTd84FDd6G/BUfyAMX7ND+ByhO69HbxLRtvb+QYHPncI3w7vGGibErscnM662IazgXdBIMdyh6vQ
056OLHzKjrQR9QAufqVUAuGmVxPKlybg74Jh06AUZ5CtTpS7EozvNmPHEGtv7IRjUxnHO61qxB03
RZLmu6g3uckfunx5nxTimOrTYgNLz5raPcyTGgihQIztyge9I+/SQRAzSIRgwsHGJMUM1l8vETSN
jbJ+5hp1vTHrNqHOR0nnzBOijWmC6rJ/2/JVO4lezQzaVK3/davUXh+AQuQng1MMA8/P3P/yLu7X
/tptVaq12VPQxoVB4AhkrQlsCKGqkWJSKS5GJA8cXSbUiFser7yT7oHDjbiAol0Y2hivekrj9QuS
h5vslcGDTgnSQlljMn4xvSKBrdv4QigmdtYnKxZ+hk8dYRZ483HsLm24Ytsuyjw+1LmaxWgar5EO
gsgzQw3KYdByvY5p5NEMisHqLyxS7lBzDOnhS+Pz/wcHEFvlK5wWFRjtonM/TgA0mBTEvzRhWD6v
r1UpT6BMRAvzuX8HVo41Juhlphp+cYBESLtR6iGob36VJUjKv5XHaahovQAhXEuVJHnyCn670LyO
GCILo2P9NIZaQxrhTpK5HYavC3GrVkv7i9AM1g056c/NAR5xOpL2U46gEqQSsvy8CnWy9doe9szl
0twPMSxs2y39DVB11+8rW50gAmNkceA8b5O0HYeETiJ+Wgd+nT+b17XXSgZAAmtNG250VJuJtPP/
X3U+zsnDFtpgpTnUhWb2OAYC77uv4ztRBHMld1UslN8YUvMf7V6xK6WX3ZzrlXbHe7FBfBEoFE08
bkXYrJ90RMohqxmoVU5TBt9VhfkPYC+1K2fCinGr02IUZp44na660FO8uxQf5OQ7y3lXpPCxA8nC
TCj1Bgk5nBtYpY14xLQmq2KLY2eyVJ/AX7kupf7VzS/JOA+52V4iBFjggJmDQjNExDBQqQFYtaee
yEMno2LhOJQot3cIaV7woqPJzZ0x+OnDJD94nlCX0+QDdCEoQjY4yd2u44Ysyx9ZL72l/MP0cg00
ZkGDeM0o+vyJxJ1jZeDiu866/kIFfS7ichCbYOxENowiin1blwq9VH3pSUcp1Ukj/SWY68v7IhYq
6XMmAE/dBHX2Ki4OveNv0u/TCbnd2pYyCJGtnaiuj7Mmj0KU6KcZbLrtcn0EuxpkIxH44VOnuuA4
t06LQi6g//rMtojAgR7doFJvumZn7lFA5AeOFC5HXf+K7AK66qt+XKfqc1+XaAKe5ydQDfzcfiWv
nwYLEZpagr0tlBZt8KlqNPfEsw9qhVAGX5oyLnseSCfkKDCYj7V9AdTWdf+23veBOOP8gtGIo7ZL
H6pgKwY5fS89ifQD3gaYRpstFczZZ/NQjHdkeSQS8B1lzihf40Dno3tNKWF7BDGo4Y2Z5k5nrf9B
77+W5e8RXHGxxFQtcBQT/Jq84B0e7lSpUsH8jrOLYUb1CLlL6WNYza648VsdA2W6KmIwCKK/r4y9
Fa4ty8VzBR8yNyK9okwfFfOwA1dMkVTa2y/tdeua3lmgkPyMh+5ZsA3+vvRZocxRGG/H3pHq1M7i
oRVhN10Zm+2nEkZPq8x2+JRPolI6Oh02fRLK/Bb2jzZ4ixWpFVYjaI3NFUtHpPuoweuV2K484BJ+
rIHuJXBs8JEAS1SHZ3FWd+eocopYfy81K5wNN4nWlTnXMLOl+UkiDPdbU9R+ToFKppc6b1qthx29
TnWvTjhaKq/VqFvPZKt8nrc30mwNL5DokqaRlKM5O5SnSguyclccMuUB8Sp3ZAz5GV3zGJGQneHL
D1XoFP4xkZdIATXJddGq8+BpAWz/Dml2PtdDgpzPbuERb/hIyCRGLqT9sxM57QzlhTTMvpo3m+N7
zTO7K3XwHIiOdLhXYC5vQfYIGagDQA1LUhnFqXd8hN6Z4CbLzhZCErwjeOGoWiI0NcpmZAEQGTQw
pqdO6dxxdj/rw/E3ftLELMotWdU1lW/ry5D3fLc1ze7vLvAG2Xy22o4S3JAc91NxBg5nHEDbA4Of
PriMO2VEtvLwrMA+RLUfUraD3NS8xQAAoTJCcHueeM5T9+iidHvnic09Hd+DqA8QOqbXMZBW0j7e
elWQjOwnV5kVfn07DdATI7aOpmaMdN3vWgDdDZAR9Mfg00m7k9lzBJKTinCpb9JH3ewCMl64fFNp
QAas9Gn+0us8+aoq1Z0djDagJnCQdkcFbYZY5NC4ZKmtojVodKrE3ujZC+fANM8+bcCt0SjpSqsV
EkDAgyw7X0sC4FDc/DCLtr8YAHSJ182Djju9UpPRPajWjIB8odKpdP0P3xWQ4dFM65YuE3bqYDkQ
1os3c8lgYMGvw1MGQHMu6BUjVfVbX2Fk010Lt/5y16GejE/xUs/PRZv1scvBFCHl7C9BmEl3iP3k
D9w35tw5GMuVck4L1O8NCZDpxujyyYVhY1t23Vk1CcecNnjEshoSnFZCkMuood3A4WyCtwsLmas3
LTd5aJ5I4O5yHqmo4LGpEbG+Wwc5smSvJO242DnDYlMSC7+ZNHPsYITdVhvqhwtB7NLO5aX9yWcN
pwIKgHbxVhLZk5PnKBMbbg4x6hp+NvKP6N/VvXaZTUK1pgIkD7HfDnaQwvnYh84B/0soRFUksSYw
rlJ7xTr2KvkGQHN35oakATdrjyyLjA0pDAb5DkS03JEDgLDxqnCO3TCIm5+68JGjp9H13RsoUycN
Tx3LSNLRsJa4ycnbQkIvU0qaAEMLHDWlzkycnnXoloChlL/mRZVQUZ07hKlz+FT94v+tQWmI3rlq
m4ZOWt8UyMRPUntz45BGPQfUrCuhmvRQ24oxGUnXScxF7lzalLgma50z3q8Gcv1Bx+PxPLaR9S6k
uKwaO/ghiTwSC/CX0vF9giQQ4K0W1o4HXAaxXbQ/oggaLBEmUv79pDxZl/6OQ7p2ZCgAWMfYMmwm
oL9H5DYOB1u8CJAaeldo4OrjZtKSCwiR87sc3p+6fpJRte02lo/tr+Hj3Gai4THA5aSspmhGc5RE
1dyZvJJtkitEoPlZBwx/Z6gBvl6tVrSUIPwSJPvuTwByQRLb2INi0xmfSfqoWSubJSX+/x9HWKSq
Gnvn3fexidVQYdVPsSmAsNOWIC0pPVfJAXh3MyaGkeonG5TSrpJ+YzOtyb/uGr9joAO6nn+CB472
TgHuy7ZFJaHjMkkZuWKXDSX+XhdbR2b+eAgEdVKYZWcrbKJCE7kyZXotYavWfoRRH6pXoNCyEoYN
3T+p/jBI5qA5dhrzuocF9ZTRDo4vQN4C4Eew0s+Fhg1KmTT94BhvrIm0uQ9HwgL4nOBve1+FxI3o
/BUzOFb5gtMWKOdVlpTXMuQpgOcF2I39ZFSH2XUy1+lqru8XVg9VyctHEyw1Hyg9q7Q6vMnySgBO
DYIe/YN6yHNYjqT4rwIe+BIUScE6X4S0h10h3N6+Bz912RZqXv5Tx9T+1Yd4ZxH4XHl+pzZrt5pf
D2HfPIGYnJaWuGkV05zicY+OiFHOCeJCKlQ6cFbekLdXPOFV8ERRjWy9v4XSL56IW+AQ3Zg+UP3a
/zyes6Rk9ayo4YDkxpzNSKl8+t5GNpAbuOpSRoJIVY5a4gqvgh8lyvqHdygNvoBD5ovCboqhxHVI
ViTDtJ56/J5YWMNAMwggYo+N2XybBl2ZUR3xws6eQt2ZliH+vxYCQOAYi7Xpzt1GD15H99/SVht+
rLAGU7VaaIxFQg0r/rP2Dj3vpXYIvq1C5elavWWT0EseqnBOlEPoRvezSux2eArqBuhVZzc1epOB
28kIELjA6KkJ5qbs7OjzXoSy8QyIDR9XVM959MeMm9a28gEbB2bV0oUbOrW6arnPlnmx7s0QI0/P
n9TxB89XnswQjEwjdBFxv6M7zfNrijMoU1AgKZu6exsHKtjBVy+FDoPui+9aOmjm1p7hS7jBbZ3u
NY4sMnGyi5GNQAESUGnbUhwPIWqdsfAPcqzVfD/g3pSwsJ6qkn5XhQdb7m+wELZu5rytZdRhlq9v
gMVTZU/M30rdjJOHm5YZOo4iq+7kCBBeHq3On+Qihv1OFnJHG0IbrPd6USXvB7KUMwkytd417Cka
cTZxKvoXFQtrCOjVKAQ1XP99mWqpNIojjBMAXovMXzcA34XEOKGsLV37LAvp+San5cFQZXAQw9dw
TVjQkNFEKbQopa5ZS+lYZS+Zi4I5ayHQgc5Cq6QWs1ECez28SLuSQC8T6t8XVwBkHkXAgV4o0KEv
rgGYe+Zf5RuSxsyPrhkwefd+x7YtwHon1M96to7ev7u4T86iQVehSMAYmsIQYCxwHQFCx4CmR/iw
kVQjzHJNvdH15yeZYsZ3NvCaavfBQ5boALzDdIh2Odqg3BD71QWNTsunQrLfA5O4oZ77iny6enpT
ag7aYYQ3twlQ0s3G6OBcvE6/J38VkdiMoRqkTvvJdMnb1utWR4AV/j3qgpv3wEB37M8LRO6s9e4I
fWRvLnOGr9PxkJlx58s1ibDLiLzliFvUuoWF0D610rlo7unr7k3KnC954PEd1gxqAW2ChyLw1Qu3
lElzEfEYFYS12l46LZaezUMjIVQehIy9GitCmYCI9+BQHbNOZ7WUAwihQzTMsSpVyr41In9h7ftO
MzBGbU3pqaS5XjWC466RnxdGOzm83Sguub8K09pGDS7AuA03gTMkFpCknVMdo5UBkGrqtVQMJOSj
edF7yM/yh8CkLJqbEGKXBIFOFo7aR8V7VIu9ehKUh/omJcHj/LZORs5pHhNJqqj+2ddl/UUt2U+U
z8JA9Oq9g+c22gHuDOLGJ4U=
`protect end_protected
