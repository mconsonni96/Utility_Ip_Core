`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ImafQ6OuGPMUWisxXUVVEUaI3Kb513dU69/1thd3vpox0ppj6ECAJFuoT2bsisbRW1cgN8gzY7Kr
r281WEO0rfG6lhqtoOTBxANewGgYGKBGrhJJqlZXONzo5Uv4zHtP8KQhiKG2LiFy18QViyxLLxki
Y1YiGNcklyPZKxWEB/tKDy+wlv2A56hupB/c/DvndrLyody+tYomzkdSQUBJTrgeUJqLmTYYOiGv
lKwBMLO7LZPq7ojT69eFiFCbeWvqc5FK3dbPNuVahOn3HIZbjdrcIOWMx+RRmxa1bPapY+EHvIkb
jdj1IdbgG7xxvs63Vmlyh1beXYNwccQJlVWZtg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ff4JJm8EwD2ni7dXwwyDHlt7dQMvIBa5B1QP1cTRn/k="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25424)
`protect data_block
Bg8kVe87nsbAFtrc14B+1UMetyZA934nFlTAA6rYw+KL53jUEAttSj5EpH/eZvRIrWYx9JtW1BDS
fK2gaevPQs04AzT0wU0S+If8l0jz3MpwmviooheGHiKCLPJfkCit368YCMr3fSKzH+fn9e+igC7u
LdP3HbLRig9ZUQ0U1PaQ/atcoTiHuErpb4lcwifC+FTUTH8h6IVMLZo/3kqzRVwT5A0wBOY9cO37
q9LzKn9C/7UW7LgxloY+YZaJWIvpfzvYxrNtQeK7cKBcFpEWE2F/83ytGKpGbfm9Jpc8ibVuppny
WgiM67V+9O9va0yPHJAsJNwK5xVx0k8F/KSmNdaId1orlJz09SuFPEBcq1xpKVdwr0vLn6wKjJ72
TC2zVBgeqMR4Rtd+lRwWVDnL4l3IsrP5eld7QdwfWlQtHG3Cqgdk6OpSUBIwtQ9GqUSdTNLM3UnK
4iTH1r8dv05CMKKaKmbHPD3TIoHiA2Wf8R98iYJ9wWMS5MG2NH1hiJkrjYEoR2etJSyX6T8gvZp2
RDd+nAFE8ktPJSDd8kTmE4qhi0/6lHnH6PvkWEGPk5MAfPEwWX9NuWNgVbMUqA1byW4q/QtIQkGy
9eWG1nhJcygapEzygzqBiQUuu2Y43qkTFE2e60Y7OjShON1tcr0MSHISycfce3TFLkPOxg6uHHT2
QXzojEvexkypl+vme5tz9LSCHXKyRhfhkEhXOJgPKU/1ooDVczvIiNo6y8PoRTuhJcNpyQ8RYvqp
xPQhfYLe71vSwJbUuE0vCmF7moKIuFJJdM+Gwst5FnlTocZP1RBqKzzNDsu7SmnaCcbRBWs+6KSb
JueQUkJAmbbmKTCA2QfS8vzXFFIWUAViTdSBMYbs4oe0N2EdUnFazOUIi+DECpCy0GAyNHt3z8CV
qkLEFIKMQ0BwoSq9Zo5Kv6S1q9nOULfNGqw88MGLgYgw9Vyou9M6TEmRs7E58aWxVEifxV2U5ibJ
xDzgp4ZxsUsxBxBeQn3UE9vVnRxdIgkTGj2Lq9J0y88r6ardW2KXWBZ094oz9S1tc51c0FSdE10/
9y3bneVE2L0XQi+UbbJZ4focdihHSYs1PCmqizOl9CpFBsI0H08ZUi7zwqrXlNUcR1evzH+kYkjc
GxrVAcLgMN7bkKUiB8ZDwOiH/8KZmrqWUD+oKnuusr+ArmI3VZwEx5KEd8IHcNzYKKJrYCtEWgJ3
W9DDLug0Z3lzHRRK0hFjN+Khv3wKcrcLO6AXQSpwEyIUa32klrML6mergy4LIMuUMzBYXMbNcUFO
yGZsiUycBsSfMjIq5eDkdgxf3GjHwVT7mKlEWGFqsRuZH0Ko1EpARpduoV5du4VyQYyXNHQK0l+u
bYqy++FGHI2gtTR87JUeqqF8/dbqBYlSdX8hCLiYwW4dkpOqBQstT0sQMI1y47T/k7h5tZnBGp2C
s24zrVlIZ/SohQXJpPs7ZLzgUgYjVcPUXldH/kQ+a1DNG9UQ7ZwYzIgf8c5kJmtMB0fxCqznrkmO
j+vtEeGVLscWjC0jkMf5QJiecn23FjJzsZe6vXbXD3JPabHb3amuXpRawexy34/josaGGMmyu55S
NFRVRTQ0f51ntF1bLYN4yAj2AlRT50NrbW8nrp/0xVxtygrA4FUAENnszOYOAKDyDQZ8l2QRd9ys
QxPojfmqqwkTK66/zd925G13367rleq6nDaSIuWx36xJMK/m6n8b4GgMvx5TeembKv25pD61OH0O
wUBpPcVRxU/Wjqr/HcVGtWAkKAgMQ2MaLFlcMF/JbLQCwGlgr02D0dVjTi3dv0LWHtyxDssf4jm8
7xf/Ac8Vj9pj+Yi/mDKjIMLREikOylDDXdDwMTGSp1McSprLpK7rL30JIPpjjKS/JQ2R7Gotxqdz
cLYw76YoPUXgEgCtoIM4Ocb0A5EapowySkqzafphAk8Q57ghD+3LeD38sZ8GWeiLaH0d8iMkF5vE
pt+4ZIlKQ1eMrXmYklTF1k6HplzTyOvgzBsq9DxZJOKm5/qDrkrBGYnn1KW+hOaVjfMf6uMfrOnJ
idzfICtvQbgZHLW+V0XoCXOzzyPyaYq9XMlcV9Nvty+Sh7rvW3IHBsLC0dlkKLTr0GYQ4Lja4jj5
Qu7o2FVmDtNHpIz6+DgIO1I5B1Zr4KALKfM2QtVE0xQfCBsmRhm4jiml8Omibgdci0OLjDFYO+LU
WNtsS8ZDXFc/YK6UAwkmkOO0vODvwu6RgC2jAbuffml5DzmEPYln+czhXqPiCDG1UqhUx7rdvmKl
74gfT8yLYNElaMF1toFK2YB5c0nngSCKos+J/+BXcqKBo0pInBN6VLWdrbqoCbzbLAaBwZ8/mOIO
FBvxDh+Q1kkMheXssSfIGOGGN2E9evt8OeZy8t9RbbpXB3uiKLGnNuEAUzKChL3bfCpXnt4aNF3v
eFTeO8p4JhqcQjR9drLuhrAimmzcghAmXb90rjGJFANfUyMlEen/puBHgIZG8oiDigJnEXjEadsw
ibbSFHk/AbSYELH2FGu/vbK+n+rNVFW14Jxqb+TvQqX0twNFLBBWIuJotZkr8RIZ46JJl2M5pcYo
LC8s2OMbGjSdRKcCKCT03UH61tyz+LQeIlY71tVbJmarvvGVUSRUxWJvUrOXlvCyPNbcpD0Ovw6D
Y0w0LjHygYPnhu2I0l//o7UUoIcp3NcEzsxcpfpbnIr78EX4mpUba20ygLmY1qXXxVIr327Qt9L7
LJ9EiRTWQcQ5wlfbZnKKg5gh1gwkkwyM1/ZLoPZoVn0eV3uplnf4cnLCbh0pEm4trbs+KJ9pi+A3
Nx1KrrHob3+1hfTaRtycFejrUcEaKZP+mNcxVEFcYOHfMBI61Hs+NOI9Rw/T6J2/+432F/mda46p
1+1WFk7T+ZlgDdYJReNAU1k9CrotdOdV3PsSDE2Ya7e7bdgVvzU+K8LTywNQONkchWVy0E4oNt9D
l/BFfIFOezTR3AC1b0SLdrFw7Uvw6NYE5MQb4vZe3YLyQNC4NBLRIoNKe/30gENuDzCZFsujhfLc
J6r1an76YBKHVPUb1gqtDlR/4F/jtZnGr2ing+MajTytQGS827IA905OGR7akBmzK0T8GiueY7lw
a7I0fgJ63EGsUW/snN9QnarJ9gQh4howGFryocnFf/SLa0/V6TW63lmvs+sT0TV9EONGENQDqhrW
oS1aipFMBXHdKvbZTNG8y1cXCVx3jm0OIr90GigAXzTzvwzF9iIOUbqzEelZWw7mWaQCJb2xRGnU
ebeW8+bmcIO+lSktghqFQFpwyzAOSBX16z9lurpny7saTN5Lgbc64BCjfR4mw80Z3KS7nC9Nu6Xf
K2e51oBhEyeKiTVeMVsruiqYHmDJuHDSkfvZ7X9oVAe4LrehgeTgoHpZOLNG/CtljkPOtxZoXuSH
8+W7Vrf4sQM3NzkYBCID12tYchA2mFKhwJDhrIaNkc1096G/07x1LOhOVsOhjww19fGfmB8BDTaF
cKQF6GL/KTFMIwU/iMLyH/808eDdZJlFOnyuQBHerdoCpmEkCIKqCGjve1FupLg2Qk3ewjI6zrwJ
TKt+AKdTTOLyaoJpE+r+viYqPMgqAx054cahi6pq35W5zQUa0Xv6tThwAvOH/ZOCJhfzxfMaU/MV
bxowMhf7g9oPrmH1N+iDHS9L1rl1DxKK4p3cy5uOOdarb++7d8snWMc1RstLgPCfSi4QwW5CWHYV
33SBGFSI8FcYDtc0PVy5TpnvJSEAw8I31k0coPTT2QQo8rqG9zyRd65ah90HRftt9tQ0mupl2jJ3
5lvB2Oc4Iaq/xAYDotbEvokXvwqG492fYj92caI4VoBwh13tTcVO1o8BDSd4p62UnGUlBMafWlw5
9NRo0hmDLUj+maS9CbNvJvre5TGOnOIvSN2h39RdY3AffUogHHBuXo1OQMcW4SSJmE7fuLi+7dWP
TiLahYZMSyXzJHBA40v+Z3mzBB8xlHL9XjoGoERlB1vmTafLrDfJ7Hd05YUsaLpMmpTh45KhkSos
gvwLE95e7pno5u8m9wjnq+E+uGnKZVgBwKo4PEcIXa0sagqC5y9TJgIWnXYO3vlo3ORAJnwEfrxo
arHrNgJIhKv4Crf+gDiWioiYB83xo0KDw3he9L420pjelluZhpqsA4xd/Yg+lt0dkygYS+Lf8qvb
ba+QFScI0Two92v8pMH27D9OGslNYAJkAOCOXu+RBz+16PSrcfEXyDl3X2AAm5TTV38I8UX2ufUW
RJEXoe6iXQUYRM+0pM7oNw2t9ACwZwJe95duteGVIJZJ4y6gJTHtHjO2AuVo8XrLJnFYoJucjEpv
fNWWlJ1ExaRzEyAOgIrOBexs1dqeoFkFwleWKIG4k9ZZTxccbVJBwSWSYHmmHC89FR2AMT9TnJyz
gcBhJ28MCyThb2qe+RHSIGB2njr8JI5di8oCBqqCRGgEFNyiAGTgYtd9tRd4Uj9hpcJ4dDMbhFv2
CZUgJQwBwEOnkhiOqObUImtWIUlEnCO3K909kYZ0P8rkcZpyCRPxVt4aXYJCi11HsYSWR71HCy9s
x+wUiIKGZVWwTx+m21/5LIbaD+3LUL4lhwcfBl4RL+Se3q9n+T7TTcER9/OPpPXol6vidAE5YKHg
jqWsvuXEeI4lO8ycHkH+LdNiBJtM2lcEsxuj3E6UvCD0b3LkA0ZAjPyfr/1NI+is1Pve4WxMl2Os
ZlnkTGgJGq8ye1L0DT7TLPAXU8xlJn+TTBg3CxnmxoA/zFiN+CVsGp1zPxM9gyvxNFbUTxJ0bLAx
NE15pvOMcAj8Hx1BfvvQz+TX7hk0jvYCNOKUX51HtG9Q9hATdr3FvZtMtT0xl/HW1ugZwMA4IYeS
F9mcfg1+m3Ix9EmbZmvbDMgivyFBBVt2U++8RxtQwSqNNYpxC5wzjsE0KI3fAfHCj2G/2fIAEyn7
WzLbrVAZPXqXX4NxnrHaaBdEYTMqRSWCgGb7c05wld6uYWjEmJE6BECae/HkGIza1yEr9ZDM4QRQ
/7rUIKN3NBUMF47aBV2WDiTjE9k4IF4mmg+S56EgWjYvVZrkTQEFD9SAXa3OVmd3oPMde50khjik
fjOjBKoPf7uJpc1T9jhAjtQ99IfZlxdRukX7Y8D7h6oEnMuQdF6MtWdoKFmgdFLF0+S5m83COW5X
euqm+XwbIv9IlOcADxOAhrPu2kFL/XB7H+LtbWIMct7AMtxOtPKUTnrFq1ZAGg8I2GT95Vlh+ugD
9tLptoC9WlEpmQW//Js0beqn6ZuuNQxNWQSv/CSrsKdBNeOXOUUpm6WYeCKDUhwOSec3z6l/eZns
qEu6W7oScd8jnwgr/GDaHjYUeVWR0czL7gqnxEsrZUR0zXCw8nwaybUkUgIq9PNQq9UD1koiK9pM
gHKR4tmOiucoFLEX3reGxnQS4caBjb/CeuQqBFGwvNEfMZDruaIJKMUVjt3pbntN5DMHdVxfgvVh
teVxN8tV4byEDB578sh6Ib6gYMbLTL1WCTU9I4YCciQh4yu4Q/G2E4DTG5cn1de533V13VqBOOkW
WpXwSe+dG2LHn46gLBSX/za1CUEJ7T9tfNqQNHal9FBnQUG18WAM11RHUtzsgs4QYW0+CgiPCmBr
XgmXQ+QBjnROlcUxTjgIYMcOrRwKETlY6w3RnyKMNLSLi9METeFNWSlcsQFbYgNVaPK9bdPZ3ab9
ckAqZ6f3HuN1tctLVik3xlOgm5+4QsmhuU/tM5Q8RJ0ZP5vPSTlGIdc92bgHbSdWP0Ww1bAKwU/7
mJYT3OG0ipAsJkmqugur17PpAqj3ezVf8uP/gWqSJPLwhuvFaeb5h/O7y2CvE1/oL3lHZrhpxmBO
cEv8JOQUV2CU7kwR5OICtIhXbU6ROgDY7YNKKR/rhAd6vKhmpoN7NOA5eSfC/b5Rh9XLByfE9stf
nbTdi1ZZP1wvYG+m9wkWLoEZzTHXWDdzb/cw8duuMhGKrRnYln9cjOxo6ehYAlwjn6+4ZN76YIhg
Ge0O5tB+BU8e5olOac+stjXtgNTfcZHoI9Mf7XNiKEjdRnq1gPENq2Hp/ElwzDaPWheu/bYlHksH
oPt3Us7oZm9fdLgo//oNoSVuWHdtTmjTSdN4oilXt6FlwXwW0zsAjA25UYqE4tOEwb+t7z2ggZ0W
S5QQ7Whci1PEXFda3LGD1FjVIcGm56/9HsEwaBftTdlEPAyZ1HoS7T/ycW8HmnEXdmi4O5rTIH7B
T5aOnZ1Wh8i/8gmB9QqEPyHck0fpIe2gsrPEbYff3lRWm6ylYMuyLeDpA5nXVO/zcivU2kQS96X3
SEB84zQf5jfUsKI9YRjLhLCdLrQQNgDOBCruE7I67rcPqf770DQuB+xZSYVxk2Bu3ioxGJqjVQ72
gjnW3GO0Aoo6OkjaqXsDrY9ibwSdWBJ03dtU0DqUNj6o5wbIlUJHuvPO7LVhKXQn+IJr+mXU7qd8
IUk+EW01h1DjYuE4SbeT7okE/dSftmW3hLVIBY0ogBrbmD62v6NZvLetXPjJw8cANiJehrTkNQul
ekXkXkkJ1uoommeLEygOKPvE1pYdTN9JOmwjQZ7iVSGbPObkf68xTM5cWXxCvBxyewTnMeE4D8BN
are8n4mtQzAE5tCFDN0N/vbR0jzcPXoDH1UaFzKd7bRUPXrSjtPj7e/GLOX9Kcrgh+Q7RWLMB6nX
UZSJvn/wlBEgYPDbfkdMM97l3wQJz+kgfKp9RjOX/QF5jyuBk/hXAUQbdEKX+ObrRQn3zUlsfsZf
ByzOM+gnAAljIRjMBI0OzZN92I+tceTI9T95HeDz2q6VbZr6eBDnogOspSgop93bl4XwlZ2eu7Mk
Dr+HCkEDxoIEZAtBZKg9GIB0H/wBvTml8eNjrhs+0LR7vnZPxi5vXhZ7uu7fKKcmvMoPaH7EPCqD
8St6sMmNQiQZs1dbjXQbj0+ddV819OlV6TbG6Fm3spDht4Mi6j69oucmCe5jPthDpOn4elv0RF/n
8qyrSUpYA0gMhFAU8ng9pM7fnYuru9e0ohkS2GOuNbMe/CIQW9avb0upiYEfluAyX82RE/WTQujP
FKk5sevz+aX0VMm420OpyjuRxkNlD65hrvZKJ/FIvebS24uamoMUg6x2nszQnQkAy+p/FhM67TjG
FBGni7QZN+t+8UBO6C9mlUWS3RLdjgyMmsQUCV+BxnaS25mYSLZBAMq1KFsTIj1wTGDsdpftpEx8
b0xadw5NwoGIsiweqzacfHC7+gxMXTTi6JIVaIaV97q17Th4ba2TyvM14FYDgViwQeC4PHwzHS+x
Fm/gdqbAqT1SBzgbRWZ48Tm2EPRi34/JADT2yj/h77ZEYydGOTX6D9ixlWcV/BfTRAHQ7DO2pB5l
Vd4fEJgeDi3yriO04fA/0GqwrZ+yVBQaPBXTSFVoKqONK7+WJNPeXeYerEsILjecx/yZSldX8CsU
NUjTscOcoSkklvVNUt6skfugoMazpH+9Ie+Z7BPl+D5rMlmOuS357zAUm8guDt3KBcJ4TFk+oLR8
4jDdfTL+hIh3QLY1PfAR91DIK2zIq7vtueQqQmohqaJiuJD5UZaT5BBdlFuEitmLScxnwHYbmBk9
JVwdhwSI5ZPssWgQGcaRJCNB89xZpfTkzDhk7pUhLW/e6vy3tWVqn6PAMvRT2WZZvB3s7lB7GPre
L60grWBCzvT8T5wYyV6mri+6fGrKkmS347X2ITgdSRhfcVVbbGv0TZRaqohjFAZ9YkavDNB2JNSd
adj8pTA9ed/9VzE8RlYH6+5r/0MtEo6kbWTCGEnHuI5Ght/7KD/ttvuyV/d3aYCXQ7KMXVNevQTb
fWLMZGybyHnLBCg6SurDyjBriZTFuLr3SRc5Iuv4jslfwbg4lDP1+aCUEaL9+ini1N+HACI27ymI
ZQPHd1VLDeofIBgQCYKW9KhC3+SFzwa5z2ADOlYjb7uy2YBooD5Zq82z22EzOcCP7ZRzZByjmf1k
5UxdiD/BWgARm3mq0IUJNtcibdhYr4nbXaTCqxoYIwmnsUdIrmY0Z371qlXU2m6+YjvdWxj0qc12
Lsv6k9R1PmbblVwYX4jLeTsoF5w13ffJUOFacxiF4egyjp7rrXYqzWI9T9e4Qz4/J4ssmpZmYK7t
ZhALy0ylUmWXIwGEtS4ThfhH6wbv64a+zvkQ2Igc7M1UL6eGuJb9j+cMkUeM5dEqKSZxYIucmQfK
54sWUBlWq9+jZzGb1GVxiDO3FQ9zd6zy08EV/+HWUZ0lwfptH0wwNZjNnuWkBr/goojmr8RGx7Pl
orv0Hz0zE/TJIHQ/l5tskrSCyvPaTYFXtomz9F105FqqfSizs99RLnKBVxvZgf+2y1vcCVGWqiPn
oSq8b7cP8bdBUA/cCXZw/Rq0nrMEwP3a+KY8PE4sqX6X4psBm/hzzQSvipLmAr/sT+wcqPpYUGZK
Lngb0/kW7/SRCy9NEkHjAc8Wk24ZHre/kJ9Txo2iy5Y/OfeFL3R8s1NK7PCBBis1PsVQt+n1LCj0
CedMZ8k+RSk0o+QhJXqZYetxm+aZOu5QADKAd80v9qFnOAlhBf1K/XRdkGAOAXmfTg2lmgVKARjm
hmMgP0DmwUCKSutLUUoDnn+ZofLbbOBcwdTo+3rkFwB7kpmtlTWOCYgRix4gpwQ1AbL8Vk8UDQC+
IxBSnXVUVlmHcfW8VK4XTDGOzZsrXJG7lRmDstlM3IaV9Qy+cBbBJ0iFQGdFFFmGqWn4XtFMNL2b
DQMnI0t/B52QEYhiLrcU0IW5U+djSpKPXrxSypLSnBFINbyEAlhsFkf219nODZ/NTUjzsyrgll/l
7dyteZNUttIdlw1KgexWgSjGTkP2YDde1z/v9Ry5vqEMv1JmHEe9+NWpJDiC7kKknsyBvTcdmCzK
VF0nK5fi7H9yzDv7+Bx6ieKNpoOrsIn4QRuJL2ErWlsMGC9IsbB4sPUBE+RW5/zuVN7PnJemcIjD
+i4uDEHW09PpFM4UPLqDXuOzfmVbDeSpnuNGEZAbJiRHmmPf7W36/egpjjavqHElkLKvk/9RfMGl
yPFw7VaMug0/Zx3SXKlVQn8kEWydol+BvFjK+yCkx28RZi7RimXJ7u5hlqB/+wSMIKGeWXpMMj64
Mt+UrWpUqwDKqwN6iTbXQF7UU4gD5wupmyYH22e6rcAcAu4fTvRXOGkGv0NOVNVV8Hbh0kn3J9CL
ECFfSuTaA830a2AaGfTB5hLznnu3VTuPP3ltUjiDpPRX7axWNGt8LSIkpDxu1KABdMXP6PEY3J35
2YOqBAw7ZoiQUvVNf637SFByMEygR7aYGi/9x1rITTnoah4VDTfaABCbnG9MlW0vb+UzG5R74iDS
tepPJ/hE113gmTNUc8ZEvmpVYHsURrNHrnD7OUdTpNS/223cmfE0gTE/WxJDPHa7R+Zu+KOHCPen
ZBBDLpO50s0+jWiUBBWUev4lxq1p1843J997RVNHM8r3W9NBYaSY4lwjnr2pDhORqO0G9uf7/shU
e9yaSgVJOfJBNi08lTmmxpt3XJXp1OYHiDvfKNOYDgVU3aK8XrNisj6jzkfmP4Mre/w6BtCNs7Px
BICKxMgdfZ2LuZio/NROW8cCXBoSz/u1AfXwBubRNWHJR3p+Wdps5PxfUN1aKFtkHxyE7Y4ok9yy
UnntwkzX4oRsHWChrLjiDCf7tIAn4cUSjoyY5SbVhksD7nnJkyl5/6nurTEx4KSAyBcyeAEDeB4+
mClVzp2m50e8SBI9KujJUy20jQVMWFkm+4hHTvfchAtSK6lNgJV2ENeIkF40RvyHlSRFJFMjcc1t
immNWMQ+EXVNAAUfNSDphwRgEY9Quo4FKhUn1Mo7NCGMlutg4MkhtDHvTjDKtkjV8c8+53hifRtk
XEF6Sq4C6nkXdpuZuQeY62ussUsnG4IGp4Tay0/+ooakl726YOuObKfPMAM2V7gW0hiiG7aUBjWO
d9xTlPrhqNkbdUawOa/WRCfpgMOj80VW3FjWjvpQHlhC3O6TEMSxRIJJkHvn/NXrCUVaIgz5Q5u5
sfBmp85ZX60UGfGTC4TKLDjqrjXZtr7FdlEVSL7GOY/UuDQskrji1+yam3xMFbn4Kzo/CD97Cgs3
Gn3x7I8ZrG0Rf/UYk/ziIbgSE4JeDcnRX2DTrXBuFtvY8gHrOV53vNRSA4y+UCZsnFwdRsJljzHs
Kv5oOMsinzznQdS3vqkiRzZh1E8/kNsLT8y4K+j3nB3QZhJCNvBEsGbIQrGCeE6j28UHLo332cpv
u4aKSdLOFfqNYaqgMl95cWBSLJ4+HypPHEAhH5t/K4XE17l3SvKXXStCrM1sddaJ86ID5+oxGdUg
wbUOdm/gf2AO0PiTXsaHAlNgpRYHU6jYYAVV5S/la3wiTNUysI0cZfaSdk2qi5rtPxFccFPdYA4S
eW5AH5zv+DvHmv4Z+G/OgZPpTtHAjH9pC6oNFHySYwYlHzYZ+hJrG9QP54Lxa9RSo4d+QP6t0VV3
kVCsigTsAjwfUHEYR6D4eQbvIqnMXncRCh6bHWUWGY4Rhvt0neYuVTAD3abDQXQlkWuwSjwelbH3
o7lTLRRJi4gSSur281g9f15GRnfabSpui1P3pbpiAXOQ8hR+ZzwahiZ5vlHe5a6m1Kk5LKsoYVpp
+FoXjFJca5husyrOG4+iknqgYfGNDwEx51BV0zKpJWQ0fWP+QW60Y372Lawb4AIvbCWeCkZghBUI
J4yBNprUTrVA7cKTuoQbkgyAknl41qY380DH/bL7JHXLkM//bDFFER0zwohxC55g+vYEuDnVMHbV
BBrb/7n7ksnn+PWPfBLYuGjKgpP7j3uOMgaiS1MBXKqHXP7O+rT86XJwpGTZLs6Th2Eu1/mGGR2A
ZKWXizK6raopE2LUyy/hd0CSYUFLL0eoF1Jj71FEAk9DwTum0TcnO/mmZ+shE+rTPOpza6/pjMKf
g3wZwIgfroR1Dy8FHhN7LSpYn2sBP0rF6BYsTTGVrhfi7GZAg3ALN4jR6/P7NyD15iD0OUYAiWfU
POgykkTobyLNYaWndFyvGSbk7NRdyzJFHgPy7wuRKb8cKfsfFRvBEPXrY/S/zJuQxn3/uhorDcK0
o6Pen9jeLefNbGZ+rKpW8i/LDUqyjkmmZaJj2UMETuIVIx+exD/9byqTnPHN/iPTP1AHUce1S3b6
hUrXoqOQDK9zwDz8H8xiFKbO6ymL6kgaImaE+W7wvCsnZfk2aV74EM4Vi8NiycI5gV44JC1FW2Jt
mxt7wr9qJAmlblsGDem3UgStJDLIw8co18Ex9nTY1/Wxon0TH3RcSx1/9hy/OCOFSV6KgZNueKcC
DNNnKN6v4PBvKss3sSnwai2VwY5TFORYg0G365UiJ0nh9vnOZXa0AIG2cXYkrPJI+ZDY0HPAy7UL
cuDMevZdZo96Dlo7MYWENJpB2fEjK8MPxUM7l+JVsh3XQfv44sCcmity+W5UbrfcAFiU//SKBUPX
LjoOZq5xY4Qowg9+MTl1UC55px/A3/6uTtDbg1k4+qCN8RUjOO4gEG79rqaR4pY+9sl7nV0wkZGh
Blm1T4Sik8auGjSc6vjjQqDlHbQjI+SI8dl2aIqylOW+mhoCkuT4kD7aBv387xTqoaRO1ibewXhJ
B8NNRAbXKZZgCxysp9fdRYCGHBUcNzj5irFpisCR1KrAxkiGPPOK1V9bEq4kPE+7poICvz0vr3+7
my2LuuVhfsqbqmlXLmdMjCjipcEszMPKCzeyfMz7hU+dqgt/DXWqWPKK2RAWiCuvfRP6pUduYE35
4xtp1wNrFk/wF3yanWpHc3B3+w8ppJvYfBmiCRCxU6PGt8PTBvw1mGQ5MYmSZ2PhZspsfY5p4SQI
PqSZB2h8IuJhNh5vZiD2jp1WgJj4TftXj+1Ba4cbfqs47NEQlys0abNuMWwTr/LSjeM3kIVOTILt
IIb8CxXVCWTd9QTkfAPXyVW6cm0uG7sq0bXWi0AtwcioOnW5xvg6uzboaHOcwg45MGLdXVG93H0F
dwf3u5CdAaIa9veFcYAWvbG6sn/JdqmdgOuCa33Q2wqqUpuxoFXKL46Hr9qHZTf7Rr/ke12TKm9W
DMCk81+PgwtsLHd7kwhYtoVrdDAJyWgh0475JwhKRk9DUhDJsi6S09hPqzuwp5CPSLQHTMsMUksc
5BA+vGuRhS6bMuXlex8gDU1Ta9sEbXpTYsz9EMJC7SEhK8u6vklVaUyftXgdLC0BjzfsPkas2AnD
pUtso88FrjXXF93vfoRPahifocqT06GOKsUFW96ZF9og1dxMr/0t3D2uEPhSwBbcJK2tWwnmAHx9
9iATj4eLIq0GcYmEZyDcQPP2tnxCmDr2TmVERae1zu0zaaYLwR6np+VEjbGwPJqBQsptAnkdKv+S
Ode/VTUmjuBT7cnW8B+oPVtKjtf50LkIUXfJ+GeFa2aZ5XpAXmnC7gKpf9oQkV7oSkhqfSxXKGtg
7EgZI9RHhJdY04CGjYsooOnWSQRDegoaNDawgZK2bbXkfnRp1CwzarGEOFRx6wso8tTYtnaJ0w2S
NQgThZRzckEAMhdLVAxB91KB37oKDT5S5fqFwAnxv135wvCef+75jtEWOh7y2NsO/I+CtbzKwv5L
nFBo3sSt/KZUppPd0sZDtS0ojh9kAcQGUXRGnQUPwF1JQYL2vcH74cjVV66gII8hCdeizM8Au/Vi
r52apiWp5hiMew5uUAJg188v2knH7P3xihf6W31zExTvu42nWtHMrs+FJ5WgSh5IVR3tdeE0Ml3n
JY3quA9J4N8mnWF1lEQuvUC9o2jfrF536cXYOLm23Xoo5Rc/7l35VKgL5yWlNHeqEfPQfN6PEjoQ
nBbarp9xETHkn689RnWasYVZ1I2Z5/QifRxwe/udG2FiFxCGCH2ROezz1TtpkQk2e0iN0P0AV2tw
zs/YFt7tL8ldnfFnD29EOeb3pbqW0XmwnC5pBwODdBzAlx0JrqZyqoxFLKK/JRsEYVMjc+ZbgE+R
YTXNBn8Ug807aOmYrjCn12KUf4pxqrVyXQBbZ0hfgp94vOgsvRG+nsIB/fulsggnZAsVcDz8jf5L
XbvjQi7Nq0KU3ZiUu33DA3itwHcNTHUDcH+lCDCnz3gW5NkJo+AZhsephoWZN+gOJDT45KNpA/dz
7k996ulsS6Hf7+nwCjz6+0CgT5BBJh+LRIi7awJYItHNBkRV0uVBCH9oFo6ZkaTBxLEEc37wcn5G
IG5vlQ5DmQc7eeQdJObmz/Ce2K0YG+oPITVuMZOz/TtZWm/QRzhTkDu0PaMrJHWaSwBJnwYMVFO4
vY2XuRdkm4eqznVf1nLVSwRFnYcbZa6qY60zCRoAHcpEtifKVT7EGVGtE0c4cMTH5LqElWrSM151
iaKZJH6e4zTm0cipECNLz4oQp9DGyEKOsTSfUpzRU5dag9b+OIsVOmBxQsYnZH9X4e8PrFPGo07M
ShPN6lM9+zEnTk/0ZoCF66FcIUWbp0fnYQ6Ws/L0x9x9S4P5WR33N+3Df3GWEznXNGT9FKXlaxwV
Z7qJKJpp08WHLLLEpYUArw1HSvargehIjvp2QFbynUeKfK8By+/gtXMJYW4SkfM53AZGLI0ndatG
YmnFk7EHN9MmUOIp0ml3H4l2Uq+RnpNYOihdMkdNA8Y1ZohMTRxTkAcSekbVxhG93i2q3HHK0Ump
INHr5m5hSE0mY/cDPrW8vo+qFgInUy9mePNhGcVN4rkHdtIS/ccebCwjC9b0GCYZ3VBMd20gj+fb
ndWrDmpgeoAtpt7pc0BhwxAvCAFlUIimqX2sJZw6uwR86+86jujKj7c72LagN3kIsI7bGcX8l4Z2
rdTQfoowHeC3dCtPxgkYvIjM7c/rc+YaYP8X0O4L6iixtMmE3qug7k1S+yEmWlpFUF0WLPll1MJo
n8OxK5R/DqOlLE8MUwX+5j1qpfOfi+1UQ7bxMyEyVlHOUbxhZbO+9Jg3ptMks35d9RN+LHSrACO2
qn6RBeeD5zt0RU6wSm1dnAi6nyDZsOo8SYU2f1x7ygNQIWD1U8vobAQ7qK9Eeap0lJQ45eSWznYy
Q/DlhnQrlATsTLHLv2Vjyx6oVioGrhT5q1bwzO8URqP2wT7W1NjKRaQZaKANF+rpU+1TOe4SKZvs
QSQiELPm1PzFFWDI+1zMCTWWOZt23E2HU/lcYhCsS85FxcdqMyUqUgjbM1PdK5rq9mE3mTR6gZqz
IT+uZqlEYoe9ItQ3oNdnRw1DY8mmFFZcr3TPu2ohTImGBVVMsuz2mCKWYmJYW7EP9VwGRTah78b/
nTJ9IBchuhZ3raBwGhkmqmnrDfvdJ7WY+M6bPvRgVFV2YwRPZMuhcUa+43eX5dfUqWKXhdHQYTBq
jFnvbrv7MCHZEQfBC2DaBwtchyHiOpsEEpQG+wZpjsQ4IBR+FirduJP3VYyoNgZfNy7Z32AjlW04
cMho/X2DlbcabT9OMs32XkmJscf7lk4l5ufW5hCy4VRkZBxAdj5QcSH6f679p+cUp2E+9UfSGqmp
lpSVXSlmkzZfgaZzQ/wWjrRpLKs8cMwH5Kxic5pAYipGjb43gYdG69FS13c/nia15mQOU6fTN83k
qW5M2SSr13gSCXaxWtUtOJ4wvkvlIdZiMFRie8BdpLe7vRgzBasKcgOAC6SCVB775t1kuSap6ZCK
ntLfbbnUj1FuW2ffJRcFMV28X6B/BJ5jcmNcnZgFvydG9PMcLeARu48gB4J3y9lbBDnaYYEmsIlK
kRt5AiBa9WUd4YHsnMmIDlEmSlRhOkUkCDeRpfE+YV44JMpUOCsEBRpaKz/RkicjGg1IXEzWCVOG
COkRVxQXwTC5K2sBYhbeUCNVMkzVylZKCrp8bmlYmQ8i7k9IxZquQpeNkqo1WUJqVDdb4ep0ZZmZ
qxFXIlSngRTVWnZNc8Q13I/ZAcRLZNyn259xWzi+gMkpbsXGGulDMlrifMBu667FQZl/96yOw5Cn
AKEQ6+PO6S6XVIFTLUlAL0tZVfD9JT2F3dpL4jbPMPLHvw+7LB+NUsnkXG3BTuxw/tn7GrFltwpu
9k/u1ATojEfhaTpujRM/UhKO8c9Ry6vyjELrqtcnqQ3+Zkgvr6AK0W9VwLvkBfTWDx3oiBN9NJhl
urEMPs4gEW+m96E+zSLGRmQ89VjKBFmwIKIOGe5Td0I8vEWeIRFbaJ2F9v/puNNo5DgZxl7it6Tl
NT/sLVvYgHpTLbbyTufNiWEO63zozVHKXotzbq++K6M+M2jnLZxE1cf0Yp9qZGUriD8Zj27YzDqW
GUtQgFrTnT/50je1EClG0X4vcLCj+CnlsKWsgLo2+RlxLei9PdjnK/odLWmS61FCeRYsv9jEmUeo
/bDgd1x165dOYz0KuSYI2SyAvUy+hSTXdL/0qqnMksZ5UHVx3KbV5//5SJ2sM42wMg7n9UT16d31
j+BztDpztHCioN0W/nTelv9iS7sJtUemlCizUbl4mU4gdXoLHDXkERVY6hGglWYcoDMURrl7FHJd
VPIxm5rF3pGf7RdyEqDYhmegYZR3TISbhYtgQxrRXv0O54G4J8We5xVMq5ka1VDmfxI4Z/tJzABA
gox3lQ47hFm98wDJ3z7hZchM4ZW3BY2JGLkb7qOQm3Dtzux4G4U60J4LuTi24tYD8jlAMvjrzvxr
ul/RHeNBHNsx7ro0YSHh5w4zR0zhpLoJAfSmlutYzaGjuIaQ6ybrv0kQTnYGtnecq9rZ0iIp7eso
a9Z1K138zX2hMhiBondx4CaJPMmmuw2zh3ynuQiHl25nQkKJITiBodyLa819/YvnptUKxdNZxFD/
yDDBXojGH00yOniLx72+vIMdrtebVYR8+u6BOSvMSwqfBjNj/xjFaLYX/iyeiYXdcf7N9HnYreHa
OISS8krbZnsARkMAb+St7b8QD88DvviTiRTkPihnZtoxO1/uz3jZr37AT4ptJw/5g1mYKP9dVYyy
IEivoG3TaaMhJMEREcJrsVzFDoukj7Mp7al7ADWfA/wMFPhOLOxgsP5aC1U1iEy+Su5XlN3sxAqB
NpPnt0BGVxdqk3KTXnWH3X4+V/jlW0SUagULvPCODevXKF3yacJOitWp4lhXcdDlhJo9+wkTQa6Q
qbMSjzR+nt3yX9xyNhB0rKFEmjn1SqW8MujhLL/aHECZdpKbfbbJmCKMyxJQY2+2V/t4HKNL880J
XNctk/eG6WOJvZS9UWiU7pqcEMB5oveYmTXsyTVEXuJe419QClP05S0moDK3xo2QU1jfDUNpNdX/
HoBM9dKOCDi3u5VLZEJbQTnQPp/qtjuCdzLcGbTZW9P6sqz+UkcJ1PGWX4c60UobNZmHEH0mzTut
6MSpE+YAEFfdn/5Y+rPn/FmewWrFe/2SRfbPKgQZYU2r/KqYxnv2ICZNbyaat/nqVpPjE3Owe0gY
fEJwBOvO9cMbbl28rjgGB3fWkNSuPuKuM0fC0y6CMpjaIUorUeL9vUWVoI7GWU1Bun32E9wpyNLU
2pAj90UBnbGy7TciheRgaCgphaJTMA29eA20fZsdHUjMzr8qXdpuef/eefQgEljuxmQByo95pqaX
w0Zxf96aWi04AgfZad/lob5WwriwuA8gdYZZt43hWOo2agxIpje9JILOAZs7YqtQWRimhe9AHYjI
1L5CT/kJ7Ame4zQpDN0ybdWjobUYH9LIXBBDNGTwa9kzdlLtSRtB60Wke8pF+VxyMThor/5B1cCE
G3hDjTc8bPwO3VcP1Iziy/Rkf8q6oOm1A9TWNmTksj3OWCj3mBtIm7V76tHJZfIuAfxvifF8QzcD
rkgGLKhzHCdakVTWn9M0zoULfByYDS7D6FbP8DxfLxe3blPQqiDuJCHiUIPBIn5lFNoaNS01kUow
PhXS1Qvjjo4kOr9Y+X8je7MSvN/H1DzYxPiVxnhZfr4bgJ1A3XoFvIVJrnta5FH70M/hLHLXWA4y
X//5EILK+Pq28VUNpZjkrsSirbAL5YAFGy94Wa4Tosf+wjf4mNjVU3DfzufKPuVXDDYmmphWUexZ
L+xxfR4WhLH3OGC/+imzgGGDHUEcpm/D3w4iG2eOBQ+VWLea1xqd5Uf5c+im6rvjIaam+b9nApPG
9wzDvzrr8Gdi6Vt/z0jNOfyx3jY/ZsfhD4bKyM/tgyHCqpMiRDehNaegXSxatAYHob28SWxwyn4B
jR8eWfvVvDsJLhcS9sMIwj4oC9vsA4YdbhcHCkR6d7JOVMN9OLf5bpoUFbGuLqsWHSWfWYqUDdN/
kr0BglTGrWebSAAJFglfFUwypUWXyPHmRnPzLgVbrDC+Ba5pAKBryGab67YyTpUHci5JgeeWeFDq
Gm8hTDMJNq//8H7W7dUvHtazZzcO3gSFtMtxY+K+k45Zy/asXw5pGdc7KFoUp4VtqenY4iJKYtDj
FkpA1o6dhojuxTgMP+kntja8rK6mED9vlCbTNNoPtYdyANiy+wZv8cElRiCRA6M01aARMudAadyy
FzNzpE74sjRN9GNMeX02DhSSKCFCt5AOtMcSZv919ePipoC76/kAe5bejf28iifOVFAON7ase5SW
RRym/36EKRHix61UPm56ulbMvcA2fosv6dVXBOw91BNtCsJWwio+0eCeOsMEqDE60TBFKlQZqmWH
U8cNABaMjyg3qa74Ep+fbmmaF6NAv63F+VQm1wy78pmwFftaVAO6Q0s8I2PEyIgxLN6jDgVAU34k
sO7UJspeXMbihSLcepesKFRKvozByYv2XNJMPOQ6z8DO2wg4IFI9Fe01SHS0dRkgQZDpnWRSt8ok
4mJwhA1t4sOrvZk8opzwGax/w/SzNLBcitjOYrUCoozTWHjIj5Tm2IV/L9GBuTiiNETWozWxLMyO
w0mgsGt2mPRS8oTJjhL3FJtwLwdZbqjav+WxaiUxp+4OYym73/RcVrulSYk2gG+K8evmqo0s7STe
4vNjjQEYqlgTw9WzKhE+2d+0zAYqv6V1RUAGV2vqkr/wkqINOL/qDjtaax8b6GyBPtJ9je50Pw0F
AI1hFvvcnztM++HMihQQsyjoF1S8YL3aPx6sry+RTRKb+vZJ0wg9Ruap1A1Q2OjnLA+elloFEKxe
wcVLcFjAt0c7tgtd6khpZr9mYRA/uxnmmSWiOfnccUPSSpESYw7zfM+hhJvv7KFSmtHwm1RN3x3p
QHevIR2sq653xgkGJ0C42reU+Siw3vKdqfAIcHP80ZLFspZZ0IPRYFzLuwbXlNk4Bl6PqKN2qtmq
TOIZxF6IqqQPSrUDb9QowGfK/3iq9RTxx9WoxE3af1r24a19Y+qmaheDae3v1y+FJ9vv5D0oDk4Q
wzuBpBYtlzILK5KnlSmOLypu8HpjOQUKtfgUGXLCNGiTwuhQHunhYqzay5EOJOMGrpIJm44ihhMB
aVWtmFpE1i9INDC6WKre+BE9oey45SHHtn36876YLrSMX40MMLxr+tUOAofMFErPrBBaUB1M4Qm2
CXGIXKfbAR4YVxoqD0SHwH5clWp2gPkE4f0RExaWt5RupUICdgornB3fooMUMpO7ErzqMXtjXcE9
qy4kZyBvKkdhKeCvX7ujn/52AacGC5y1QCeM5A12lIkILc6+/3Q5/DPTcXPlNzq79Bq3xiRA2+5v
INCOlWvpAGzFaWpPluMd+obr0B+zfl63YGE9saq59yLJJYfedRwlbZhxBndArJ1IiWucpdpT3w2p
FKDDPklzu+nu+0+v6Y/BThVp3JvBNDGS2/pVZEidWOVOKZcuwkxhlUSntJ/YLOqIwKAjALMS/B03
c5rGjftLCslsm2FNKvxpBZS9ISzDVbODY8hUlGYkPf9nyG8PJ4BTVaEO1/zyyotyLwrBjZpKsd7v
xMy8RWJWr1k485r1md8hmXI4Lstk16M1rzQNiXDubyjzAwiKoRZoMS84Ofcup4PxNvIZhPSO85BJ
rZJzgRcOVd4DN/VcgSt8G2La5DeVbguxb4sA/kx4TJnfdoNgAeEHbN96QwewVh7lDvkyMhkNZYz9
1nSGm9NUwc5m+N4gm75XsIHnScR/W6Cn+WgYlJulnlt+IGkS7KrVKK95+G4euqGMnj3ctEBwRYst
juHmQbFcgRyURD9Gl6dJHbTyzXRVQC7VM25cErfywdOl4u8aXZ+pTXEXqssNIOx2Ed8L3AmZFl17
PNUMrXHnmQno8UXUjiNaZmZiCDsA8daJOpJCn0uR/U7gh4W6PQN+JHYmUXxJ2AE14l0l+uKQ5gnO
MpUNuL8Y8hOWwKOEtyBVjmhoOuVM+zEONZModxFvAfUoNAcKd4SGo1BDw7xn2eactFl74dqgOYka
6iMtNRA2IlnMuYuXrid6WcZBEL7RmyoZsyVeO3JtVdx5swa2dLFZm44HMD8Ck30ECHtIjsztEi0T
fu6B+cj8vpGR+74YHYtrr5iMVdWj/JEYBlK0VGYxdZSqWLG3IQZYLsmxuolMUgtaoKHBD3ZL0NTp
KEXKQa6JDJjVjNFAjZGyUC/nnE3N2Dy4sqSBdqeHVxAQTm4mRT7EJjCtLDQJ7433GSel++9+pLXH
lNpwGmD7uFD+b6l1GEiUF5wVumLqsoBSpfXnFiVcKgjnHcBUMHp/Gfnu8x6KsMt3gParFPNMe5hM
lg4aZt8s8fGSGdt+GW6Dy4s7s6DqeTnBRa7YHYEXRi3sck6LV7n03YBorgNDe8FrQ8FDx8xZDxy1
P/CRO4GGPhLXIKwODCO7OwWzHD7ofQ031yY2+P0jxoFyqHJmok8t61/QCPbegfDInsPqM2voKlPw
RixIHnSmz5XnZGquucyyxIb/g29LoCP/a+upNkqdt79fDH5wtN2/GEWaDvXS0iqt+NQBe0VH3pfG
RU3bO/2kKqbOI6ue+CNVeLboOpd7CpWQ85MFt94OgiTLi6oMCa99so6QHp9drlprjm98+RuIiKpE
vJFm+6n7JgopsatGFPzwsqDbiCWJugKyhXCDFEa56Y8/Ks7V4OHJcglmROy8wzMsrr8BHeYQ9q01
v+BKXQ0TQknM2msOw8Szrr2nF8hPJt3WyBxJWh+G88v5DLu9auuLnRtEM/QMXFA5UZCKdaagvoCR
yKv0sgCd5DDYEvPyj9weix+dayrWmiVwQHCkxeZ5gTKSzJGK7PPvWxBgiqKyaQrFM5Qr2qVSwVHN
lecLgmJ2rAC7GOMcs+4CE5AgHktofFv0yPFglTDr7N70SytebZdPGZhxIrLvnXxnbab72NGUptSo
40DZS8je9uXMlNJ0ldKq5noKykA8r6HUJ0vxyNbNsKb+lxH/tu5DS8fdZ0NC4SM6fxFeSY4ThmgM
RIco3ZtZktWhYNEHWMFhbNGC61zrC6EHF8KkpeW2uIu/tRRMiVo5UgwOOaFNszuAyphzOXEc4E3/
qQ5xRVV/ShYa5mYYYeW4FiHRzU24A35he1j1ICeBKTHA8EAncfwqzZwlz+Cc4qy2SiD3DPITD8V+
rOFdK+1f4D5nArjhpmrWEoopDYCTeTaf7ot/VSjvitk0pbxJZFzohlcZ0jiyF233ucBpg7cwgXu3
GV3nFThvkDSYkDlaPuG4oBg70iWDm4XvLO1jSbwig52FgXJnHpqA856APXhsOV4pGw34UIusvWXD
kX2Nt8wo5ogaMa5UopPm07QX/RnTJkTETwh4DMo2KB3Wv64e5IsBhHO7o6H3MAX+2H9tM1fskHkX
u80UZh4stReYa7R174Lpd8FZp7hyTptNDZGoF/dfQiGaFoCfEkbCRKEwe8BS1a9zaUfR8ESQOfyN
gZpYFpYkFkD1Rl2qadLxSO9hTVBKLWGUeOVK2I/ff9599StRHiymFtVfx+fJcJbkuPgOzzBQGPsS
w1nd78yDK4+BXwKvsCC7p5tj++7rgCIA+mZiYcr8r4Xy9lwJYEjsQ7jTbTfI8m52DyHxhEvgiibj
d7GVQ+sNASaaY0h0ii7jfX/mK0j0k7vw4OJAzrVG326lIfL1oeUBoYFoMna2nDS4OsSfhm2ZKgGH
i0UYy/IFIeFGOTs31mqh6wq4+7Z7E09XXTclktmAioZhiw+epL+6kTbRZoimX9WF1zi/lyWLZpPo
NQ6uCT4lddJiHawlNk5I0ZGMVto/T4xi1Cl/f5mSucokZmtcee2fMdimweIoXgLMsaFLMgc0CmFF
MChUSIWOIbyaMtTrwKKThzDtXNOCbeww6CnxZZ/4Y0F9CWvn/PnJF5pL/qW4VdZFo1LGOWvEsy+X
lwMCPeIxWwDViZPAFBmaSo/q9bGr31wD1ePsj4NyeRKwsnoiNj8Y798Muo+vb+ALqBggeMricMO4
5VKi00QukNd7ws4OLdp6SVKdegU/ITlbCuA8KXRFGIFzbsel93zIseHX6/L5/PerGblMMVSNGaZY
R5t90soSe4hyp05d06K4A9kh2qQIUAp8be4I3f6tSCFes1Iu3NLVhGtZm6MGrCTyo6aDqiYBGfiz
PmouMRvIgcAp+gXuVPJVK+IMeri327qD7HMz9wwTYeHxdJsCiVMzZNWDwCpTy0gFc5pHds11P6Hs
ZoC89Au0phfgegHfsASKCjeIIdXBMvWUHw30LY/CId8P6BZkAjbvhwim8Zqu8fHYs8X2d7c3mRRQ
AEnYUCMSQtDiY9PYjr/9uzYc/lnDp9uXMaEWDILDNggomVuAIXcawcree/n/cE8NlWjRx7e4XNBy
/dROA3n1KjAI9KZR4unigRJW3cVLi0Xg/o02VcAsCmhEC28vI9FD7TzZUokUMEnrujSXFdLTJvDB
5W2y72Uhov0TEgYfb5pmyluCQ7rXypFyZ7zFBoZPdqroHwWnFw19D/qRJgV7GG0kdmSgXyYVYqDl
S3m2fmmALML1TFwEl+sOsnh69GVQuBjt0mJf+9HS6DLqXJV4vtre1bNv4Rh4ejA/J6PArnu/hjRT
CwdNFisPzUFvkukNCPisln3hivASyTCDqOTjQbw6fDZcYHaee6+x5FbLTiHqWlivNt4JcjYkSTeh
NhYLTXKqUIqNC9PbXcWYmLWRndeHGN8rz+X5JOTWYUWMKjtgxx2dOtIE5yyDVE0XW9eM40yZ/Qyj
ofUv/trqBmgJxkbpj+kwV9SoEYO7qSyZ3M3jlGe0Awxi7RAZsuTge2E3lTr5aMSQf0a+mEdExwT/
7DYLX6e4uY97eUXa5RxLVnIlGm5fMhDAkxHySGotuLyRP2r5bRgglaH+n6xuTIBL1DDj081DY1Ox
S9Wn9jK3xLACxVj47mAkNT24YqepWg6dzaR3xjnemTtTUk/4bcyLxbTJOGvATHjR/SX0gGDg8J3w
UGQrBoRX2bcNbIDu5cDaOlQ23BvczwHJhOJg1pwToBd1DbRveTd3epmupMJLghveGNpnFVyUbH7c
ttJkjQwV2UQQgLAFOuqiu9pBngNowIONGAlJXGgXY+gUjuF2RDnNzqkIkWNAm16dQgFIYx94xBz3
5P8cDrxygprA3Z/wQE9JUCcx1OA4mgHjiwKy+9ZkZp/kJFoLE/knt6N/NE7423ZSbq+6OOLRGn90
toeBolpZWXYIy/wKyWB9no1eoTQybODOLrhZoi1q0Z0/VxTl4HNvMvJG6f9ZgjGSvjRN5Y8sd18L
7ixzcD6yoAj+XvxkWzAfMxGLN8KeBsargg3i/Lgk8csrhp9fDtIEzP+lgWTHSQSwgdPbMHsOPei1
Q+b6xpHCcs4OzerB4Gm4xaXJyX7O0pXdhNW2rtuuty4nGCLEgrMAMcqOMEUIwtNxtdoL5nJ04EW8
T+aI19zU6Gnmy0sswWJxYrKA9nzSdd0lQ7NHXe4TU1V40rj+K0npRf7eSGf1C9VgMbyIscD217Be
WdcZjd2tasF614KFqkJ23G/fRfkc4yamT2tbXH4PLtvzTSbiAuChY8yKpjdrGhPJ4Jy0zLEvV7xm
dCuLujCqwm6c+kvhJsv2lE4AI0uVCCfGenZgVWzuyTiHIwDk/fL0SSo9Kq4eHnaNQGuLNt7bDOgj
VKsEO+12Ozzp5yERT93tSINdbIXLpiThwr4qSVtmr6B9Nn37PQMN8UwiamVaN5d9/KdEp3PjwpHK
tXberM0A1XXNcL+Jl+kwQ6NOEZhCkwDNqj7nfyL9oM1hcIkoQiFMu4hDnONAKXO0e8PfXVmmFPYq
pAeTpwZ4v3zcOj7cFf5XLNVSiyhnH7Q8wRX1ygrvLLQgCGqrBlPn47fJYwP39vlE911eJKMtuYSE
nGn3z7bixWHCSj8Ipy51dRb1DYAZ2BuhqkZn8pBCriZK60L8Oyjh+GEt1nK2qG5V3UIRnUPo5oBN
I+8nQd4d4r7cLT65x3sIKtnsZw52J8oqyF1fuMvO1AcCBGCJkNtn9eXE8w8hDaRSXvpTF4KOafH6
JdOaP0nfSzee8aZvn4papZ2mmi4HA8YOPXtOIQHtSzNwP1d/7lmS+TsHHwnrVoYXsZQH+rIyw32f
u4mdCzGpafucQRyDywK4VOyEbbzA1hUgQKBbKyTg1lG9wxMwmmUwIY/OjhxmXoa5+qdM/wEJOolN
hxzVlUEeC2+JH5UBqsd9NM+xndkedlCMutzcGDt8FRgrTQYIMe9uBQV/LelB7V0RA0YNpUH/Cslv
XtFuHzmr0vZVnnUIo20SR3uAFBKTbocYBSYHTtynqUSdpDzntngTLOskqQFHQ7hox+fmN1aAzpcO
8T6d1gqKv/SAwQ+Oon5aMQrujOErkfGIXW+EbEJwIcLNxVqWDhgxPRxMPCAPL2jXREQIqXIt5nIq
3NDeHycLe3RxPAKBGUnU6ZAwpc/y72eMu3N+1W2W7tG7wN6cFxVVkR+9nBe25qyzUpVwprC1BBEL
BK0UqIHeZ0jFrBDEAguxl75z9F7BVGLAj3Q2+fN5KUQytDhIfSqjVtxISs51QGjolOmbVDADmURk
kMM2j5xyZmPNO3hse6JMCkAIfnI4NdFAykk5N3PrJG/Tpi86Fgt8TgEiIpnUq9lhjheC3ToQ2jmW
Uf6h91ruTmI4TMnq9pQfbSIAlH1wGXqeW/qwxWaRadDCVOFIYJDQHxu063WSPfb6nxiu4/kqKw+G
g4WTyIoP4DHQSMKnCHq83oosu2/7DQ9DBW4JrtpcbCKCXFxX1hQpZqZAGUFXPzHGy1VZao4vG0R3
5pLU7QAUiD9RKw+LYo1rILKufaESOjaHZIGLG2yueHcK2DE/I9GLtJGNMsBzRXnSYpNxdLZvx87h
xxYixcU3q4YzdLAyTdTFCmcLwa3+FeaMTp9q5HN5Jbj773gjV9L7bcpzq3X3bMeKgxhOtcnfVQov
AqHzH0j24CmcilQs6pyDMJ4OQcQzm2bbmRnu3JbutV/MukgtdZcVTSHjXoFTuvO2xN5bmGQKlxlw
o+v/DYCNwevgTv1aoz+ZxeSzhmNPjGFUmcE7PF4uPkIT9ZJ5I8SxzH2d336hcfntm+lqJOkuUMtk
FsQNhr1jul6zVxZd6hjqFhAgDw3RMSY85fN2QTTwYft6qwXxd3DfbwHv8zNMARungAdSVx48EPje
AMZW1q+BflELcvPu3ZdYSyH66w8y22s2KhXTaFwxb6FhOpoIRp1zgtMcTeGsCSeeq2VgmsX9rl+A
Qes8uZvHFwkOJoSMd8/XZElynM00AZIqMVQEA0XjO2+cLhHaOgSua+PJufKXWK2O7Nj3iBT3gq4B
iNaFrKfUpFpZmrLVE7HMcX7hRnyDezgA9/JFBxBorwmbXzYYyK7ZLtANTrP8eE2odPpP82tbokaP
7mjFZ5ct4WoeSqnqRTWH44wapC0YJKiKg1cOLqIai2KFA7sdxoxcokxBEstAo4qXoELM3x+ZyigS
BbsahzzSDoNLQMZYlNZcJqeCfvJCi87171Dr5SGiAEJScg9VQV7wNJYFmsh5WElDQ7ltU7cD/f9a
l4sn93agWBRGU4ek1RI3xeofq4L/w4CUSUc9srVGFxp4YUJ0H+lag7gmeD/7eTutI3jmtO636HFb
VXh1PlMz6iyXKRj4/aJISk0ETXoTctQ1EfNLbu75UlymusRR4/s4k0lur1rTmJhVxO3Pc9drZ1Zr
AOQ6qR/YXlIkOzhJA8G4Ov7yqGaQMxV+aFxhMdX+z7N52w128cWJV5xd9qI5wl9ImdZxLhNE5c/l
hejXqsYyvJQ282OBtaFTcPgHnUiWhksB6fSs3heZUaI0x1PJscA44KMlfEtAMVBLlDaxOHMQywjI
JHkJF/HbL/mUQxImY+a8RcK+oDpAFkyhmjqDKJGuQVAM9p/OkAxGX+tBrB4uOFfzyA7bCv0LFOZ3
kQcgXPZpPBGW2BtEr8ol94JdJIsRq+RZ3Xx+23nCLnp+v3D9wCfx4OfHH1Z822HMm43C7gXGx+zV
VgB241QZJBd4kUuS3DnF5lBJbesFA2yG5RI5b/tUKH2qniYARem/QkxoZMV49OwQQeP3LaiW5WOC
4xUTlFjafG4jthJ4J1UL/o519zLQ/Mp8N+KMdkKkv/sQQdg1w53BoCzyxZTckGzSiVCizMRlj5ED
3BK+Dm5g3goLrlGd/3Idi2EkD0otRcbpfAqoY5c39GQ2cuXszSMFmXo4AxIvG/5IrgD+wgTfhBwj
NncV4e+I1Vd82jzidTSG2hTXoSwnFIjtIIoni387nd0ZAUBgYNRDtY67H0MF3liBrCQCB73kSXmU
/lwVHblYfHlXe63oi6xFjecnricdbGwSZnLFpHva5c7VzsTUurdws/T0rtdfHgEq0S8PXyAPMWtk
sk7Gj2H/WB4FbBoU9omOzsgoBMKEysP1KG1F89PjMSlSzqtnqiSfA6Q7B7cc8fzaG1d2YyXxykZ2
VZYLpH3LQDXKrUBHMIlxCupQ9cxYQKZsjXWI4PnY1Ap+If+rqQPk60+qMLCaISUoGmdEZ3GiK+H9
L8IwP+rW14cY6MHQF+L7OXBcglwxUDzwieDjk0gvVTJuME5MudosRTGX7G2bDxv3wlAseJqaBEpD
Gi6uqmXV0dKwOhbREkLt82TXqV7bEG6NmzTnhy6MnOYc8QItuGkSTI/a4ztOYq3VAS0+jrYBeqQF
OL7a7IhIQ45UUYj4vPkGEHNwb7CMZag/H4FK/hj8jkWu4vzCVC5DIZkZdQ7VCpwN/ZM/ATaHZQtP
gPX37Ioy3JW3dceHmIgy5gDlwk8vq7DmOGf5UsMi8XHG6x8G2uv6sEB+il41lL9u32ZeeVtE9+pa
7JQC2yXSLhJBzibne+ScBUQN0wKpzAzPjoLVT8yL8gRyUOE3SSQDrfs4BJGUgi01invROoJBGm8+
Q1SZ3VIFpe93CcgnHNC8O7EfKK+xT/iNpG62If7DRhwODMSChb1mQZf9lPUhslK8TVm8ia+rdR0t
vGyUAxEyw+5YRWLivJUgrDivD0HsJ6cvfnVZq1D38NLyVV36TaJrQ4pEEBDui0jSzuwHNtJa2M51
hPtzeaM6xK5TOdTDumlG2pckKnpEekP9v31jGDhGjCt8SGZeyBb8s9S2l75r6GoPbFY/dmgffRDE
BgXcohXNojEcvkZ1beZE4qLYfBeeRjjSTfmQYf49KiBXB0xBPrlmHW6pZD9Oi9+07cBw+4HYW933
pnhJXyxY5VcClUkBXVwF5NguWUEvVBUDo5ZKsnY9vMGnlXpN0DJSspb+DbmFTVV/pTXwHpFwc/ZG
MkA80Bia5hFnaTJwS4YaqEfUzn0mC85nmUdXMMlNUTBa0Q4I7WXivciI58fFWlNbTnUg7W1rX0XU
yG7450dMBJUFY1NMtF3Q9XAhQ2mmfNCdk4fckmw08At4doc0htoRl89VllaPySeuveokmzNJqL16
rbiqBJytAZ0pXs/7KwAoHI9IV76RXFcHPezyw+Wm87c/7BxSVkCBU/942Xr6t49Zn3ZHhe2YWlHk
METDoiIljUPjjS15dwOv6o0pxtZaj8/RjhLXOVlGGuixKAp1t1jC4pssujER3ZqNMexUGkCXhZ7I
kWVmGmsVbN1myMsz1DOYO5lTZJYg5/4RWtcDXJvFzsNfV3mSmPntSKz926N3SIMmbuaCFJO7t7M/
pJQBRT0lo4Rw1A4NFfI6Q+twA1ZusGtI8OC77fXbaBL1W+sLyeQEj8MXAP4K3wnyWd8/PllKFKtk
kWuBiYe79qp2YaU6WmOlca0k960PgK9zxqxmLajakfoxkw2r4KlOMLiFpnWLSFqk704yE/8CqzAW
LMOgKGUJwLEA2YmR7ZHZV0ZZ9BXeYKbRZjQj0g8PKAa1Pk8p0229NStjzl0q8Z0bLYt8YNnapd7p
IJjPiUeXNOqqwg5QcJ703Qo+250A9CuYzTkfK7Bp/qFzLg0E1QlXH5RhL9lmIkJXtANaYaNSD0Yc
FYxYy3KCOqu3Ljt7XhgXbmF36FvGj7uMt3BC3PNY8ns/tcAsnHL1pWBd5g3hRKRG7BHliDmwFQoK
Sc2+SzN4NUEDz8pciio7aTmiy+fe/k+OydP+7Cjals9hdUTjPoePsX+TUXMfeh89/CX+VNJtLqIQ
8s/CdvbcNosYofd49NuFqp40R+aJhwaA9jFZLNBbb81D+dMiNLa9Z5t75hqgbvFmY8ChFR7lyUhV
Vvu+s4ibWOcZ81+yIZJ/qLBSR/0s7l9BBYrUV6kPbfEysQRFUlJRHNyuYwFvhqrrxv4FW49OHpLP
Z7ZXNQe3g5EbK8m60D2uFEoJ7SmkxJtYJczYv6lrUE9NwlbNEmfo/FtHizXH+1u5fYCAzzS1M/gD
7wdIc2WM5yO3kzIl2432hLUwJUK65UwNj90zcgUgIbiyeoSadvIxxY14QEPOY55KlVjadKVMjkY7
5DGDuwiC3SoDRITE9o7TbWoqgMgI5ddCbbdYi00hYWBoXnxTnNXjN0oJYj35KZeRRNWMZZUyNZgZ
wR1HKAg+zuWU4hyvvmL0soVTqveAFxMBhXSuCs8BGlqoKzfor3W9l2AzqFtiJbyHdVWehR6UQMCn
w1XH5ChLkngm0Facwi/7ZyGFKDOefFqEtHi7Ekrn2aHvVHzviVjJcxBUw3cryYEf1RTU90Ao2Zck
47miitoCJvlWkiaClcPPa5GQ6lb7omOlgAp1L5jkL9jtnkH5FCIM56P+SAaOB6Cd67ISFIia3rfN
2v6K8oxOPzfTuCvurdi60uAjWHTkN4EVnn4/cYUw4a1mYHjwRiF4BMbKl39iGQIoELB7z3VZ+RLX
Mbh2zHT0iz+pwlAGMLl8sTvUn/A1oteUeKdXy+mbfBrngN3MRHrDJIK2DuDwtlF8xvFk2P4n4t4F
ROmGbH6hXVY/4ZPBkJHsm9DjjD7CIS+8wIsi+umpmIfmKyYuHL2Deav+QLsTKouW1e8f8zuIVW8N
5MupnXy4rKzRV7TLv+35M4s8qFbtnxjD4NA/2kIIFugCpSgYWcVAuF3z3ViUVy0nJJR9cT1IU5DD
gQskd7vPPLxaPjmjPSYKnWAs7ApOFM2/pHgKB/Bb0kKvwkopbQ/GW8UtbN6Qy8Fhsn/s2TRiZJMq
s6L35YVrLk1tmpCcfvyOQILM3j60KKxA1VaL+bl4BPqMq8Mp50iCRQjE6QGh8OwXsPEJCxTu3Rfc
Cp7AKvNHIQBr2CIoKpJPb/65h7z7TgHAH2LjOWAJq2jhONPNu/4h+49zCajO4kErekc/v1DWL5fi
5tgMM/M8lStmEuDUiHqApDooCbaUkJzVEX+U/YW4cwHnPNH/iUEXM2flBUKG90tpye0eYlFewGlv
AsDDDSRIWuUl3rzd1BLE99GyVmi462WaJcqfhF0Ick5p0k90UxR9q58QUzpNVWq0IBo4s/T0pU8B
sdraTC2/6Qc2cj31NkUvWKkkhd7uUDtgx4Dxpz30Nyj2+6rrhZ/ullXf7a1lm1ZZA1UTjuZ+NTsh
wo2paKX35ao6ZQ32zFtHWAk56GLQNv4DBgGGyQptSLZ4RJpT4yr9SadYByuFwYdk/qDHeI4Zj6Vh
BPTRl+5GECa5dnjaJ7o7jIBhOgnysxFalJO9zewIv+dLrX6o+ezi7plGSoki91Zvh9NBpFzNo08N
6ZuZ8B90mR8n4AS3UyT+enDeYzzSLofFgWxqW6S4fCEz80w4BYvF/E3yYQSPu4K7zrx2zxDAA5GE
Wma96DSp+tGOZiEaJiwUFGTuIg7UBRGKm3mRjqA3gKXQSoa0xjk2/qov0TY/S/tQPP2L+21oDrGE
taBmqE4SzWivKh8UvFXZmL/A2upMj6ceXDTj3Jh4h8ryZRFHfuI26eRcHqHL4IAdsLne6PBgwDSp
J2FFhcSDDlh8K2iURiF9z15vuJ8tS1mJtccwPWOp0LRCKAKcEFeL5wrCrXTMBqyLmG66gKp2yTYH
MHVzFmhloOuuat7nSN7NQV+kzFy66ABT4gajVKP06WKd6CJuJbkMlHYWzLv5LmgWvYjdfObVqagN
5wj51rgkw538n35GNb850IM37scSzAqYtXQoM4tVylLPDS9M/EHmg5IjU5PS/jvKrB0QYW1n6QVm
BWhXvKyxe7SFw5a7E4ZWG9ZXUraghnuypanEM3Hk3dTbyyMWnYamSyg/swZq5VhyxUE7jEPWovJr
702vW25lf6UTrgJcu49qiCh8kGzAbByYD9RY19JAiWi3nVAwLKd8227aAW1AaflrgKxo0JRLL1PS
vfQtK2bArzcWrdpPDmch4fIZM9XqL7XtSnl/rdn6p5rXzdUsIw1ZlME30nt7Riwd/wTtJ705Mksd
OLbYhxW4d+sXOsd+O86E2gZQ25uvL2LxBLZcVRMAbjrAujTlqo7ElZf/AiT8Y56NKbzHLf/jLV3T
lyDf3stzNRFxemWK107G3+YRRCEzppoC/3ubbVrvX7C6MO/Je3TWpjDcluGwHy6Mpw6i1j0qHIyE
xRwG+dYsQNwvmNSbLTbH+WC8Z2C9VDKZqLICdrMT/2RJzOLyc62kFvHZy92V3VVAbr4UGaLnRAW+
jsGoRPhvUIqPsFhvEwErbvB+UDqXym6MHdim/16zK+MTMTZ3aoKjmhJKgfJ15U8zL+AduYkOZX4J
rBYDGr7Vl+qkO3JALT+8hmbcmruH07/+YuOPaIollr1Xfr8H2Oq3De8Km/UU6uhShzLUnQ9oJ2I2
2zpp7EtzfHlc6vH85H0iVTMgZYWNaSaKywi1HnR4YyPv2nr5H5MVJ/0i9fW1CNOa1G91qo6yfj7J
LkI3pl48cMxpfEZYi5n1LKMVMpx1tUAR29Vsnr3NAAHopprDvfn4p9C9duVrVW/0y4fE6urQkdHE
mDWVg2EzyfpOhSxg6YIGo82Yg9ChMXNcbuIQ3Rnw2xU3YJYG3DcpNGvA9XT356Dvj4/MfNdOi4Wv
rxLA3XmYuY4WX0Rg6Eg0zt+5vcCm7tvV8Pa9xoUbanWwYz0+qngg0Owsm0pEWJ2z5ICJ0RQiq35H
39/oTVDFqUB/GLaFMqAUiaZ5JzZ065zazsfxzhJeEL8u1ojXtB9r898a55EMOHeCvleIKlb1S6Y5
fND+WwBOYcAcGfKn+NQuyEOpRA558oG1NwB1G0tCnyZlEjyDqfNCqoKK2UqU/7osKOOc/gHXcA2g
QWSNuAF/hsjQSaTfJEmC/F0zjf9CTFEJSZ3C8eMfEPlbuGVvxCtevwzWktFtvOYNlhN6TQGd7SLY
ysle8mBPaJLTTorQr1au7rqqTYSPevvqyycmHJ773iDVNM6Wsv0EbmJ5QTLmzHld7VIFbntCLeso
Gy3eBOgWR+TosCQh0rnMVc3BbSwJZb8ob4VaY71QdlwfQ0GZvVOC6Tlk3tXuQFWuZgOHMYu4NGpq
8lfhC4/ztTVA6IUlBPWulvrmQSpS3SYMc9oJwSslFBMMjF+NULwAJ4SNCHoCIXMtSjWVHTcjB5zG
S3CQNdqJ1oVHb5Tsrg1p/dbBlPSMm1J3njGkwy9jjVBrWZnAgg+hRD56P+EgTTxm6SMSd8RxD/RX
wplRcWaFIS1MPYeIjwOdUlus0Va5dTXw6pbf71I5MEG/Opa99vk/STzhzAyR/p376juyG8ZNpJno
WaXJ3eVpUx7jwKcbnIptqtTV6i+wAIWftXhOvHgFuYMySBZ9Q9mcA7ThUj8UBwfDBWT5nE9HOCr2
TSxIZSaWRED3T2ZjdhRJy/qA67RIYwv4QG1g8SibkmnniAJumSlbuFXDxxDd/AVY2ml7KOovud4V
wxT9Oq5q5fzonZ1U2nS5ARCxxliXKw2vBWCN+vRzgAxBAkcpBnPgHrptnT/0nMTMLvgd7V2oCoOF
2Nedm5N01+vw1K+yoDkGSjb1VOv/3bhCRp6gnkSQ1BUGmChz0Ces1AIB6QVFtGDNZxpcd6IrRr/z
PdA4GYSp8FPi5Jq7KC23ewSvGaNKDS9vpYiUrNQbJ9P6QZzC6JmG/RIFTyhj9Wp4CiP7TqGsZt9u
9/57OE13BcX/BuVifXc62l8uzzFpJeDICwr36wMBCNivW61kKOv9WGLR6gEoATrlTDCijRVeCsL1
PMAQVe9Fsv+PDNFxdRmjeRjBe5yRFhrlfCHlMlIaeHGxRpfFhRaTpLuxSLvEDEcEkDez6Ck5HfP2
LqXt1Kv959Y6tuYBcorw/7Eh+KQYE/SALagqLqdVT2Tu1WtM29mcJCg0IYIZBPzP+L8TbW2Ge09t
fAITfacuR6olQM0MDu6Yjjk/lnF/1oj1vsTur5Oh94SxNwkGclEHBplQqRiqgDC+fOM1lm1Ro0xW
2pXMAvHnoe4kOqqrNCqTICo8/aG9490s/ft3MzOuDC1tshd1sDSqr2a+vosxPBpFim5EMhK3IDrK
52uT45iZeIJwt0WqasbZGbWyrxxPlGRRuUmG1TWmGqT1sC0sIEinY1Qe5BetYLnho7rxx40euy9G
P2GsMfO2zY+/V5GJa5YsBgIxoDJ71ey2XR0PT1h/v4nSD3uyWIi3F7EtTswLRraphZNxCQ13wZZ5
nfN0Gwvy4ne1cyay9lcWZnNv+g1BQDFqiFQZaG7wTM2HbJHOmlFzJJCQN1gnZ/0J8RZd4ucVEmQv
wTVQ18WfWwjcULZlBPuYGIYIjt16l1Hi/7lDE9Si8UJ/32sz2neZ/j2RQk5gAR13BaFzWIy0u8Av
sVN98H8IjKbpZSQHzv2lHuP7EW5YzCKZzSmFdXbEo7Ch6Wzx2tElspewSwnjsIIhDT6yHMS2cbIF
mM69UwX1YHrH5RKGpZBU/ixNPb79OD0yPJDEan63iyKw62QtmQPSicojHsydYVj1Hf728k1tKNuQ
4/wnkZeR4F2RHiDva3lFxkslL1DFwJjItK83YnEoW+6+K99isUmaCUx+5PQ+3Jr1w/nl6eHyVscE
y83Zdwna7RJYuUf49kaXyOByakc/3V2HR+GxX4SO8uJgJRDyL4acbstSS6J222bAaup57AtfyTTb
DtxfmNH8dJ+hmWUkS+ATELaz6dw6R/sdDgR1fIVmYwbF9NfyV0iQwQNWBKSV05TJREA4iPpsc0oh
Czqoft7an3Hs1Jwix0ybQOaisHSmWVV1bRe0cKEOY7PqwwImrOZNdE29FInqvxIa5Txut+b4qcOP
Yxbo6j32quci7KIBLx2kQ1FywL6wzMDgmENAl9z7i1LAw2x77vujW1jlaNKFGbe0+iQroKTWnoGO
sXZRsi1cNjM0xEex4FC5/fVxZjx6r1K1KggaAlzD5MUxRr5foXs2jAefiVfLrHueC2I60QNY9APa
RUFp+wDBkUWQQ062F6uSsZhEdT9WWXLEhpCUe6Jr7Fmc0HwEPU50VTQ07FeY3fNX/WhZ76eYv18Y
HsDVz7TiBhLc/t2HYA98gUpLCsO3DOVc9Xevks9PiF/6Y/V1N1Ume3lSpfL3N0B2IyBF6HIgG/dg
DWBivFMOip9aiqkCJyqC/byzIsuPe1E65G+PAJ8X2hwED/o3ork6wtN3NA+Jon+hsoZqxoBdnoen
ckje2Br1uO+KozZeV2HL2XDaKRFwQLmJLk+e0d2DpSeI/cHw7FkEja0ESbL4pYzxr8meePVmgbcm
hXRVygn7pXitwL7jlxgLzggLzP7jOzpaCAxoZlp3lFNhnhzO5BRW8KVWU+Rva+UiK5yk9uL9dCbt
nF84xB5BhrFE0nQvK6B7MVSG7EikaVHZwrVIH/K2Rvh9YggMIiytveVEUBSt3LsUolyQmncfrpR+
5mOGAtmf2U3iKwfSE0Fpv2npxeKiI9ywdfdaKanHx5ltegOccQT+qT/VH8QYd2MRCkxbXbnaTjUR
Il9Ni3DyhE6gKQN2IYVjlZkceiLgodEtdbLCcUMWS8TxlIub7bafQYPAKNMnXnXBTzlDshQmMclR
aD5IVTkHmccZ7F/kKy/7euK0Ae6fNwon+lawRfFEfx47lNIGFr/UE8k5cF6jNpxRf9X5S1nyQWyw
NUBd/gcQqc9zZjDO5yyjE1mVLjSLO032eO15H1zASLb78P8xoSfq4oOinnw8NlI2BFB76Gov1YoC
e+bgRE8AK0eVOkoxek8Safs5sBFb1+Ox7Yn7EezeEg+vw5WUo2IlPWzt3WJKM9D2IkjJUSGiA20y
qjiJVlNm3K5hLw/mQMr/LM2inD/mt1FGOF86NsBYqPg1W9Q4DI4iZbUCts+7BFDpG6XxcdywOJCo
NWr9WB+7q5Tl2DjRncHMxSrnEZPWT4QZpXdi40UEdFmOFngiGZnMgLXLeRFTU4dnjVWhj0DLA3ds
DtVs8Wh9Wn6alib372VOCMxc/1pZQ+Hu3htUZGi4s9BOisTz0N2zjKV1VqhyLdZjYvZmXtsyf+K3
JQ4lr62OeETF5D41yumFXeELCwjg3b7y3vqyQXhjPeJ+jASn5ZgleGB6scGux+XkkiEBhrzAH0gV
KB7E22f5ZMEF3ir8WGGmpFdevSDcjGQtnkUGs6/hEnWAgAgRZ2hOS69tu3WulYGdBQdqHIO0CMw3
YzHFNQop8yQ7mvgpqou7Xile/6KcwZVMkItBtOxrJdj7bFYLHls2jURZUcqxxqN1Ym8REs8PG61K
KTU=
`protect end_protected
