`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
K6/WD2cTrHjsDg4gW1cgzW+pwdbkUNQCG/iDFr80wr08giSE7H1rPPws2i1KMwsnqnu7RlXWK1Pu
foYmajrb5SM/rhhIbGh41noM//CqIfN/UYBkM5xSn+ed2DWPi1ZEnyTSFK0KVN5lA346MJaKdSnr
Kl/sNMIBUDcdnTEvJiQlxZpH2qIgWDcldfjYuuVi/I8MSO6RRaY5ELFGw8ogFGYP+qPZlU0BXYVk
ekXwpjcUdnfBdQ32W2brESbzd7xW4OiF/7ZfHNtWDoR/dhAqhn9liQ1WZx3RDJDefhQKUCjeXvme
fkWQsy52Adb+iRj57OVUEXtDGHSn8dHBGElxJQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="cynqVDIwyFGsUqfdxvzF2vqdxV5MNXtCQ2f83LZpgeU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5168)
`protect data_block
lgObjo3xRvo0nR5bSsMHrFyYjYmlhZOTrFAD+4teO9wAWfaazaVKpk2/rB+rxyYm8HcqhjBv4KbF
0VtRwt9tHlvmzy2/Mf0dj6plCwEngrAcx1V6ncwjA6KJ7i4cBr9wGth+mhjnbBMw5haHHDlyNmI+
dF+u5ojp78vOoBNl2xmwLaLevhD7KazawlYgHIfQPe+IJiO4oV0GjC0B8PQew9jeGjwP+WYrGtPO
OjhOpoWibg+ypVLD31ds5U7vvZj1lbQebRt0OvSmWFpuQkvMZTAyEnyX2YvRY/R1/yHReBQKXLSX
Ssc/R5MdeBrKiYawduV2zzZemtujC2Fx3PK/P7/Ggxk3HZeiuA+x8ecoGhILcbqan3kLwGwAIiqm
WXP73hGgWFvJnhmdkes0yTXGWfbZplM2y2/4AQCYBgiJ7teKNGJc6vBvGWVGvk4eB/v/haiq/FFD
jxemYs9sMWBNJoSZ10yfdezMP7//t+6rMT0w52ze/iuDSpZ2zdRs/NBEgAtNoQcGYWnC7bIS3fdm
vM2KAkWix73bzb1tryJ15IJsdOcKrXqbvCMV2orWyZVnbkl6bYRbdDOsfcfGtgGeK9iIEfoyaxvi
qKb/LAoBJNf/NcuR2kkvJjE4W8N/Y7tXBTysCNbStypQgXG4HZdmodHZ8IB2dyxi9f6Z9dIZ/HJ3
XDWF5kYNN+S8tHnRSjzisfKbxxfpAXOgGeZ9vrf3fzLngQZa4qYI5+bOomZar1vsXlBDcxbodKhR
4mpElL9eXQstpDNKkTxUsTsr0uK6D4SwU6nXrpaEjxGU3hb8vKaTamdCGYuou4cAiyRNVDyGzXdH
LW9uaFOSDFcY8RvQqi5p+ZakE13mL/ZUUW3IwR/GVDBlIM9KW1Q43jxNJS8GXonRmEs1lm6QYG9o
7VDQw8/eTJAZb7trEnDbV5fCZFEkXFmlANlM0yDrfUkKMLTwAFRtgB8dAdhof4ocAri1QgQ5QQuN
Pbq5JNdLsj6Mbuj3YMFOSg/8j+rFKA7TtbHj78wyrkpNHnKClvTNeAqCwV6iMYwi3VJftJBuz3Zs
xirz6ee5CohRJqyQwAKPozHBQGAV+tCog/eylaDMF7/S0x6qP7YhuSKDm4fu4yO+1ocHGZJPCOk2
M7Jsaur5V1rYDInrR/bu50Tswdwq8S5caRi9Ztu5Xt5j3ywc1ZC9aEPVBc3JLCt9T2zoi20C1OZm
A79q6clBbcuqGWb1lOepjM6sn+/wA+cW3rA9OObQQXLutPzEIG5ef3jIbOhRBWZ7o9bLYLWicaVy
gzryaPAsdlb5LrrBQGmli3qcxVckns7Sql4Yu7WmVgh6Ls/NJkU555TSa38YMDLhZ955RdDL2/te
aEeKK+WlxrJamN0l8qEmZfLulKhj1VwAG/bE03wEAmuhSMfcBbVcqPdlWit5nt+Ij6yOMsTwrAiQ
vbaRtKiL/R3S3PkSlFEjkP8ejFtaxbq5hNl1yCuzSTZIa2pXuhAxheFoB1dmlqCp5aPhAKLq6ius
5dMd35ZYBHlw5P3lNZdQIIOmiJ+NlbiHGoy+kYO79ZdWcfuTW0/CMUp0txhs0GJ8R+ZYLlzC53T6
xiXNaVjoXQyx23QiAYbSK3eJIlRJ4ZdQJ1HAdFJ61V+zWOBpf7OLnwRBZ0qEAt0ApCdNtF5pV1n2
wCftFmWri/Wn6mb7SFnMhEjX8Y6+kFO+yVsZq35Sb6pqqq3aXAYYZN1M8JRdmjLdqeEhtpSegDd+
QkriiBrjhM6RXB2ISPe5O1McSOHSXzYCcAtQVhkOaGzPy3OyaSGDZdi1l44MxSRzEE4ll2TvIO9L
rlCMpiRjCHVQ+3HNtGCyMxen8iC2JvxX+Eo9Pq7/vogDuw7NXrpp3ZuvICUdc1vISxt0JtThfGJG
749vSWaWSkA+0HPe1TndpaSXNFQOTl7+drT/bs4Y4+5tvCNmj+/mpYNkV/lyeHNkwDB4CoRQs4C0
PgMbctIQj8zIdLqhQ3vZxse2WYp8yxUhjqvsE0yFzzeB/3rRu6kRBe6Im8ssykOJs0MydtvFRyd5
kMx1B3l5JbA9+XrtbyQA5CXwCZngTOqIXh/Bc/T/Cg0yeWymmDgH/qHRktOI0DXZu8ppx/nTPpIk
V5ixNq9xqare73qcQdwMlj1m4xSeEK6d7kmrZwlUmgVbdpYbbddXFdthDV3vb8wDfuq72KX3pjOW
ZbQ0+Iciu0sDeB4wdCCCgLo4bHtsNPhKa7tNCJOCN8Qg9n1Uz1CKpv3vmN4i17dMKUyEZw63j2lY
NaGft3GJQuedtD/MQy2S3pdTgisx3lWarl6pi7d/IHLEMlov7BvZ1xbZQbrOHtsKlZcYETC41pxD
A7BC8cD1G0I6+lMdTfJ5vdf/98lbHEpNeDzyePpl8pWL/1o69VEfOHp0oWvRR16dDQoLE9BSHfki
egfUpEkkt3M5m/TEMjS93vb4ihOy3dEB/HjK+PxwlBxpNUQ1UQH+8XKGWI79dmwLhKBM4+tP9Hnl
uad9ss8R/Ul+3GLmHlSmyAV0nG0Hd8kGrygWYLXXNKTx6er4H2sJc43msAHgf96BRVW6YaKOdEGh
ExrIo/T8ZBL0hibX/fjJ2+ok9jIZ7MNMQIXLXopjqD0qmyNa8M7rRYtme75+pU1atOJWHpSCmH+x
A2lezCxY3UotYQk5S1xz8C+82wCrMdMGASSvH8p/bAJoO7kF/hMYlaJWAkFAR7d7K5Cp+coiZZis
wtWLfaQ3Kn/i1FjpCh2J62B/cJQG6vU31q3o8/WBtiZCJiwsrwVoutUkTNGQT6rMXnhHvM2x2IDQ
da13Hj06bpv8xe+YLqOSechM1ErW4Hpql24rzNtK+Dlo0ZD/siMsOW2yiylrFFeluJy0RVRug1v0
cHezJfSpa3wS9bJeCo+DZJlH6IXj+6EU60IQVQYpkK4zO32Kaw8AykQiMh3AfpioYzXhEn87vPTF
lX3aYgVmRMjKFQHR7WJJHVScngXo9CjTzl4yRqC9MCdlo6m/SC9CP7NfAAUBd71qd/4PAMEM3356
kcCFdx/U5KxxKBDrE755jJJFruwLg7LEcyOtDCI5a5FT3Dqv6QVUtxg3jh1ZeYh7WirSbGnvOsEg
0p6Tk9gBJbDg1goUBCmY9w/PAnJqH1+NpuHwZ5YYxE8I9sBwa00fQdYVLB0pnpjGkZlz1a/lt/Hw
D5fuGjJnQKLQcNkifo8sTOF0UitPxziaQnjzmmKmcbLEH5GK77oX2DkdgNS09+hHgaRjOb3/OJwa
JRPn4jRlgpnCUvsE4/PVoZ52nPBteUPJTRlgS5R6zu7Rh8FEfTCvmhOON0U8c7K5zl+B4Yc14hN7
u+rkcZYB1/nNPXRdrUI3UQ1YrYIpoxBXmzVNqjizYbeGNfwHIbCbIFb8mEOHlHJMCSsUyY2p73Sg
N3gpOS0b5If91pJn6wXLu7CM/xGsAo1uhNUZkXCFHg+NJpdXxq5ejjHH4RQ3IjscmazJ1e9wH85s
eK1nhV7fm3HArywSa8WNWsSpGmLNwksnx5NHp+6FPnwuvUrgl43MUTz/qIV708EWj7sWCmldWloc
6XsBNN0nQRhqsh8NoQ424P1OWCmmzRMjX5Cd2WsSMM6/oAFlxI4sPrl7034st1u2XeyePp4HHuq4
rOh+OrPNHjBG+WSBqjeZikL2qIrNoWRWHImFa0+v4XRy+tF3ny7eAXE0y7qDzgVImK6cSTQo+3XY
aEvoo8dzDl2YsoKCNeq0EfX7mrX1kSMjR//aXHeqQA6Dn1CYm/iGiTElao1iAQtLmb2TuheswrtU
U9laXVRvx9kYQ+p5iTF+vLkbrilztmcnU+LeWgcAALxBGFGF2oVNhoPtz28IwrvE9Hwo5ZFwphcr
MZ6J55iQ4VyYpHJn9oM5OdI6PiRxyz2VuG4R/DuouIakqPtqSSwKz229oHCbkU1J6l9i9pRomtTr
Pq1sYqoI2rWADEXCFsnhJkEHm85H6Kk4BrEudtRPL5o+yHrheRFHM0rWjWQEqqpzF9YF9KkY/3tU
h/mskpfz3SB100ZPw+K9C+5MZRhJoyGGkrJiHzbmM9jPVRn9fZ3fMOvjefKa1UO2gXJWm6+XAlFk
UY3dzJb4sv+s2YliNGbX7lsbXquPv6Ke9xpxBcdTpgULRg58UbXMQZ5lsVKOv554OdF37IS6A5kS
SwM0IPm1QNjJQs07Od7Rg/bqUzrhSLQISWi9FwURhFZVirHSSJAUNg5B5IEd5CWis45XGuUwel9b
bGEMloSlJEoo/eACl9Lg9KK2Za91AoYt0nlGPTG2+rTgCn4YUqtlKfkFuINd3xiJSwe2kmv2zrCG
W26bmgYQo25fBSgxda8cJSJ4/Fo9ft8ERZq84rVyQubV0xFNlnRP4DdpdBPHSn54o/o6mMc6+Sr3
D7SLBzgUve1yeURWqdfDGmux8+X3F9PHtchq88oIdwhdWBonB2ZdFoWBp3hfuARKYsmt1ZjZRDeu
he6w0JL20tZHwxp8iQ6JkFNTRQKSeNxET/GsB3UggsPMKpqnoFgsa6fdTVDt/vOfZdkxvZT4s1IT
3FA1GSZlozFGY78g2P2Dik8XmdwGsIbvpJizKzMOlL9ZRminQYzuBM7vUy0u7O+BreOjpmOLhumI
sQVq/tUq5Ltvhn3VQN+NcypxsyvBZACJVLVs/ncGb/sUgd+318q4youGw4uCKnxWVHJf4Ss9KMGa
JHR8J8Tq25X6YgwDrjlg7I6p+7ZJPWspYj3KIuVhfMKgvCOvmSc7lf/HdbObLimqr2pl7PkE33QY
sK4MlFqwMTiTiZsP1fpZkelU1+23tQFqefDiBDmm/xW14OAmpG5jB9C9E97cdFA4K1dU255TbhjO
pHVIDtf8Cll2RT9c4XkubXyqrG+j5ELsW1douJAbFQyng1y6UQYSaGW4Nl7ZvdOjNK4/hKX3W640
eaNbgDpAlp4Fo/2lcSKV9Yc2DXhOElh5xow52pC30GQGWaBkYzxs1NFGFbIoTeiW068XCaiXzf6j
xtDiUjf/Kgij5FQK1gSEX9dYMjvl6KBVPwPmkCTbuIUgPLnEPrsA10f6VG8uTgG7Jc06L94E/p73
QGu1q8is0R9D51zIyulxxUy6S/YYWGHle62wP+GWRNFl54EZ5Y3n/SbkR8fD8umy9gdKmNDBc4Tl
C3IcN2qkYzfYI9DGEYj+mu4d0cgXrczntBVaymRE4UwnLVeJgNoUEixiaPITBOa26SqtbtXlcGr7
mX6PEccsN2W8Ss3JWj+WbWg9Wa6Zuf86yKSPJ4mxUbTyyMBxm0V+flpVypf1XN/Q70UgY09TYXh5
4eKI6er1RIMP3nI4R6Ppx8TAD6xq+eUMyDzSB+wTddNRoeg2LE3LpT4dH+DrT7PCfl4ean9Etutc
vhCMsK+f/0by5qbJOPVNDFC36EmcqvdZZY5gHKSk3fEsIWzoopk8/CI/TREjwP+NbBMhXJuZpqsa
JkMk4X8CxEnmQOpmi1JpyI561VR0/I+dskLx+90t/RXWDA/FfVJaN2HRoX7jYgn9xWzpmXB+oFyr
Oo4YamgoqPgLHQJtcnW/bWCLdzcbVX8JeDLAKG4uLDJtc9WhFlDFToNZ3vRbfG1YFlnmi3LWu3ql
Mjf/EvXlHOL/jDqqs3/CHkf7QeN3vQn6IsDu53ZctZjaI6slmTvbmcT90S9WTs/f98gTa6D0xnid
jqFbjebxoWLSO1Tj2fWTzAdwwTQV3ubPCnpecAn9yIOWK4S9fNZXhhoWbp8SMF0dSLgp8wWI06M8
d2HvvoV8G/vLIAtqMqdLPSnz0Tq/vHCCPBwaFWrY8BSXk+3x4osxGwieCa1lV/z3bvQzckAgGalX
G7ukmNyT4pd8yi+ABg5LTRijpFgzPbTb0wsNTL3NhaGyZDhgfg7wIauXK9kiSRZk9qEb3bSuSub7
hD12iC1Mr3W04Z7wl0aq3jkrVN2pC3nhrmyR3/MiwBzLnuGrLRJN1w+lGvEku46masJTprBN6DEN
Cz267P976LP48X2aip1MDJJoCcpoX/+kFoBwpEO1Ke/6KzmgWGHX6YI6DB3HtWY8YgdcoFcxaVeb
vYypZDTqmvA+/z3G2nbaSOi8iG4Mdz3nMzR1Sd/GgXPlFxAd5n5gWFC7ttO7LY/BVbgEzLPdhiNU
dVgsYPHKtBjwXlk2qa+2PL0vHwfs6pNf/qL17KRTGaz2onQNNg3LlMTL/Agr8I4K1bL4Gdch4o2u
eCl4Ij6evjM960gSRO/dO5vKXgBGkNYys8Zy9N0rCg85HjZyNpPkdLHC0Al93psrP+STzBCzNtPg
WKrGGnNB7GQE40R8NBkMs+OutkQWDtDTBe7n1+Zyg6nr+KcM/KAcYEGyZfZDqWMjUqtIpspBdHew
PU/xnSTzkNEGeTwBi9XYmCHT+/tTcWy8CAXr6w4bOS55C1HpfLJaK6osfUJF1Vci+rpInISYaDZs
YjCn2wuuuVJmbSHL7e05C7pbCoZloxi2JnLW+fvbGwKj0A8vP2vkXZuYqEI9FAHw6fKv15eod0a/
2DWYTGKSc0qnNF7Mws0aiPpxMHspmRstt5/dNZ8CIPxY/YcELtrdPoyyKA0AOF9BqnB7X6+piML2
WoskU0Koz6HKWlHZc3J+gHGhOCMsHVxMlDH+ekq04evH8pbscwn7vwN6IhKtd3GjDTYmro0DmCuX
+iPoWTQEteh/Ew+yrsL7y1hrCArGCUNQH76hzglYsBmLxkBzkp0VbSWt1Px3teu5BZRpsR6gGfXA
Edhlp+mEGuUZcDs5imA01yBRvqntl+wY90HSbF83+zBRxdMzV3x1VokQSBlg6Hik6NXvpOrfo/J1
Pg9+W44woqedmqDbhhwMJQE9ztuRNopnfWCqV7xdkflGFL/ANfI=
`protect end_protected
