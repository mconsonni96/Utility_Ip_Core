`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Z6jENVTQn2sQ9qVz7zKrGjKpjcm3/gIYMwy6AqAymJ4NwMe5G9G4frXMd00je7/KmexUD5p4rHC8
O+CS8Jz1Yoep5vFvHTWY5wt+/2QQaixWXbq5x+tr4UQxVN+VN1jpvYxCRsUuvE2cEit5foX+OmuH
vKtQ6k/lbWEXi8OoenJ3gdKjZZgX3Q/jqznzfEnN2ZGdKMBzVRIagKQWwmXFYdvwozt4zRIegqY9
DWO5HdnZmlDAePjWnXXhZobcGTF6kpC9BxPK7r7OBuR98wVpqRnIgssZ83Q2bRbst7834kyM4A6V
MahkaKeqt1Q1ARjRzSmgr4SesJuDUwj/rJ239Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="WsINCpOV1+tYK32ZaY/oo/z/lD/HRffggyeAl0xTz4E="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20656)
`protect data_block
H+XbgUN2hsJ9aG8g7vTffvhp3EF+NisnrHNcVfoyj3QIlo3E/5Rd0rSs0mMvRmlFRLZgKoiqExwM
UJYNVRTsnWJW2jRgx9gxmMzEGEh+qiCPFqMPA5sAvMXnBvpkpHaRm1JYBKoweoFq52Fo9g6jvUBb
m7dsGlZxrffqxM90LWrOxhIJ9KcLxQAxrZGy6LwuYaFnTHJWgQg7xf/sWU01UMIYeNVCf46PAcmG
DzFT9Aby1uv1NDtjYd/WQaU5d9wUclsnOELtVVKx5Yi4/bn2CT8u16y/pwjONeZUs8EajAsgezon
HE3DbAs517BqRUEMpo+4d8gvPE0hP8AzolxUUXBocjgl3fi7+8wRkL5ulaSGIVG5ybpgUBm5yF1c
Jjc48tp3etaUrCw5z9sKwSWO2HKkTv/C55EVB8AZYDsInDL76WU2Rcft09l9F2HyXS9lRprgDTNy
C8F7s1nD8Oq5IEn4HryveZJfODnnchRmR7gJ/KWb/JlfhAisMim7x44rHopVbe3ajDl5cvrm+Ycn
ao1AVG3w1ii1YDJLOOdgg83C7wMdGOntEiuKr0cs4hCmyrDa0wQI17UfuoU3xq+qm7hkKsHj4SHI
YwlaCa1QtSJDK+5ypMpWn2AcWJFNhiW+icJY/HgNqPRNO3xwIViRv+NZuqrRBG/TtD+GppPBH4F6
jSjbehXxRms4AkiC2kyRD672hLUIUQJb1rvepCOpH3LGxBxh3ePZqu5q95DUTTRgZ5JtATTA+Nms
p0J56QfxnywsjGFVCsAcX8dL/B+LhFHR2NtxOHG6NJpkWGN9HxbS2V0IxWPMPaEqep34NA+8aLnE
eLxgcqtn/tzOqCCTx+pobgELv3gwYeSBql4DkG9HXuwa2W858ATCYAaDl9NCBuPgQukQ6AR4AEyi
74Rahu7NrhBQM/hg+ImtZWdDUg9LUf2k+zvvtZOzKp6S9Ol0DadWQKJt/Fs+YnxuxT3pR1mCYqdF
knx32ZZPVG0sNnAysWyHJ5rX4hsyOutupGwQ7QH1RCOTd+CJPlTSgL5101NRsCHKW3Q3mZivXpxx
h+T9iax4FhiS6EB8GpQHK9WVdHOp/TwGOIPrjs+UUSIjlgpjSdloIMGh95Aww9IAj1QCyygxOrdz
utOoMdmUZ4rNm6+VOr1q3G7IQPgD+GRORXkoH7quTVKkB1UhUlUA7pRhq0QTYqo0Xu91zTcygZeQ
2zven0n2eF1HZ0QxQqppG5TVruJnEw93bAjZZi75f0ClInKml/hG12epNa7hHQZDxz85U5jkoMGI
QF1j/JHT1mQMDVLkqlV7lDynjaj3/GcUyJXRiyt0B7o38tvKGRrHxorWu6Z9rbeKLhiktDh0q2GE
AIt4R71wySv5lFouA96xOAwZK016m2WQ9Qz2DWvUp8CU99miLJzUqRyzUxP9HIi1nA4j2QwnWdr2
R9xy/Ia7fIlEdsZ2S7PhzDOhdEinBp9VG/40WcrsmU3ziQhAaVLJIARMjdM/JYxaccf5smOOZHnE
NFT+hYdMOikqLMRnsEHmSWFl8aGl+epffR6XNrwV9O9dCv5Va/53akh5Gnp0yF7LmvxjQsh5KV84
2LsE6f46Q5nAsdxbek4ejgunsYz+EzHRIHETC6oS4qujT9bBxQmedk+X2dGWeg+bQguzZI9uCNxp
p+lyx414QKmCJRd3KnqZOl2c7+peJ3TOX4KpILlzBxFtL19qB8Vc3XDPYROLcHh3ke309y4BpqdS
meQwdXCdhBPhWNiXp+y0b9FoiZmqFK+y2O3ncGxOwXf1blQl3cRDilWA+TvIMxs6mHW6gVF3dG6Q
QFLZvnOyQf4UD46xz/TU3QPxDDmfEBGgFuacya9mdZugQDC4+TSWZ1rIsqi9PlYPullV3drHIXxl
Gs7cQ1cH9A3mtDJlZby010CxCjwWVn+Do0Lw11v9pE5ppA9z3yL3VP2u3IPWI2rALj9MOz820pwz
k8On6L6vL9KLzKyvGDHmORRIe5183BPaQjOgzXUd5OIT8DeIm+ZduwgD2aCx2RA6VSLNQUjLrGMp
/sNvjXTxMajB8ntEhfoGRN+XqgM7vUsG2+nXtnrfRlLzio7+qp596UbRYhGmjkhtdzCjTTTrMCXk
nIJt2ELXVFQF+BP04+jwhlPGUWRLY7fgaVhMMfFFXcvriCrk96u1vwN3DRnjl5oYZMfnWTLKjnli
5nM446njMDdmKWoMTrpVgYIBVoNCOlMvB96yhu6RPm+nSHn8+61zinfLJDKe/fNKtlLqufXOR50j
VlGGXxDodRoXOZvNTZZamH/YuR0YZKiF/4P/EsECCq2hur79nWWAT1U3SIItIA+GqJuPTdjiy8KK
4ti7Sx3zVVdh68E7g8Df8QtHtGmFadvYfV8wHCjPAZdRf01UFRxbQL71sVYqkjpomwFLDvj6AF+8
xj5qDGBZwxPD4LNpbMMN3WZCokMPm1sXXPhUD/09zxenM6m08xsW/OH+SgaR9KqAvcHw8ilsqroc
czNlv8l6J8nnclhqP2rI3trwTwyrIkSt8M/G7vhk72ujNIw0cYiULxBfYr3eH/RGVamGpd9xWozT
zKEweIz4YOpxk96e7klCdSDk/KNf90rSSyWuGOlfCvbQ60KU4cwaVYNxK70KHqGi/KQv4lzlmQfO
wKnfklVLC4qIkhxzQY8CvfdCZQ4t3mccqEjqbHk5lxUbk40PArajmCK28jFeib5N6c2hJ22S2T7w
0+4ToTW/LLYgxeCS/33+wIqS4TVcujdHi58D1CP5pt8nCu1PBNE8NMQNAF34yDht+Tps5Mf90mbU
/1vVa6D2OgG66DJ31vKizIXKUfgR6Ng3SEux6FLt1NV/zISP/f4loMzNg0AQ+CzdS0S5v9WCOGSr
oHwLtQNGQlKPoGzQSROoEwis/Jta+/fFWBeuHbecNGApAKLwaHYKQMIdGpLygJFpIfgo0UIp0I3p
d1lij6ICL8c4Oglo+oCnHbSqp6/lDXoMNhaRNLk/f55CMHlCG/Dwtkyqhq8+AQis1wS7qKT+4AUS
q6wFE+uElTtQbVASkkLXStZJM6uA6pJynW4HAktwDtNGjulPVfd+ILxkSQNygKsgIjxYQ5CuFbaJ
jRCATpJziJQw2j7zq48Y/dXe0DNtbRUnIgn0ADllUFeU9O33EhoxEKde3Kmoez0csitxxQSE4NgE
BRkyJZUbAy+VN/a5SQpTu03d9f9ryfF3f+N92DhriegGqYVsMF3jI6tpoFmBr+24NeXVKpuNdy1B
9H2Rk/thxahrl9xI2smwPS7GDagwWAqang1rvWD93qCwGtOJlOZxeT3dZPecJFsjeBeVSMDZFuy8
PeOGFmS+DmRagQtQWswx+ZgtmfARy4Yk+9gdjH2c7ZoOKcwOaaRxak1BRLowlX1Krif07Pxg0dXF
lZVarpCyw/IEtJq5h7fd2ZubRehHwKm4QdrU5r0qdN/x6VMoym6ZfufDhz9XHqiJ3qTRnGxb4DFW
gVM4MKo95NdBzNEjXub/nf0mOaQaw8VkRi8o766znWIi0f+FrKSW4PUy4eB/WiAwrYzoGYQLZyYF
0ob1ceGzZzqe6ArhKs4eTVyWP0C1Kg9kpYP3v/TFrON50xpxBt4VplcaAdGsI4HzapoLjxOxcOuQ
GKjqQ5eBRfhBE9bNIBjRyBVo3Ocu4F1FsMbAJNKW76ed5vlXT+/vHOBdjUnGYhjkhI3Z6pgsfr6N
QfExP766CBE2nBj5Uu2h0YbGIhITOHWdRbv4afza135UDzDYq+gtNH9AoOZ0lmIHm1+oOhTMHypO
tWubFUVkGSZ9egsuuec7wJu1hydtDpAxCZYfZ3ZzN368Ugr6yUt4hT2a+B3/xSOzpXLFaneP3H6c
04L9okdJIX7YdhPuqCWacqH7OAEV16dazXd2o/XvnBv1ETXMhXCJipqhGqp1tRytjzbiE+bGoxrX
dK7HmDwSXIL1JEO2xDC1cWQ3/gK1mK8i/p4FR+xy/18OVATuAmICMPJx9rO+7ABod6Vv8NW8x+ht
dfxCUd0O/ITFIG3xpwRL/nqdbjBln8Zrl2UaGJkENyuv++d9BLkB89C7VWjO3WeObkx7+FWSlWuh
k16Yv1IXF55Ghhd2cU8dTY+En0mYGE70hayChtoQbLKL0CQSEa+tgyjO8bHHXXMFQOo2UnHCiPks
pbQrnBcuhl51DW7n/z7Jk9Psk9c2Skm/UyfhvzXcXebSKzYOlxOU9IKjDYq/j33qKNGRiKOa3GnF
fyRKrqY9bs5il5LRb6PaCnFl7eDkmeEvK3Kh/aA2n3B6/866I6eaEIp43lMgf0pHvDwIhakQqpFQ
kSZ0CKx5wQ7q7fHfwTMYhscUAtAKXHGBsQuCd6p3HpO2T6avVjhIqVOqcXkmMtlqC+Ucucs4XkOu
UO9C8pxT1vZ+0VZaSjzeplCTGQCCIskPn6AYl/Q45Y+M24XTVK9bRABeA2p5a5EwCK9xKs3tmAFZ
AgOe4UMY2i5U+PAU14s71R/1cLKvZnTpuetbf5HR5kwCdjKkJls46weMHsEWz/hUGug08F354JiU
wJFDrejZOOEDUXRHe9aOHoI1s6ESrNmRLj/0EpEfFiKzLsuMfG95KDzWT54zpYBs3k0OH7RfUCU3
yPvNP7anLRaxiNx8Y2LPDP9mAnaas1PgJBIVZlX3vFrQ7PPeQCnYauZUIVS13gJM4k32HuDuIoTi
PPYRZkWpcIpm21BB2E2A+N5sGyHYbwxSESIn1argzYwuTFEwzQVlb8+lGBTp56pG78cbBPu4lAHV
8DZRB9rQlAB3EPLwo+6gte9vBTYMdCRO67KMgxHHSwxi21njbLPFH1EJuqQrTYns7gebgIPfIARj
l0kaGa4dRJ3vtzfCAhi4YMUHEsv3nP+wVp7gj6rKwp+Ko+IqYODlCGyZAUBxVmYdcc++g6r5J4WH
ONjnYQFQ+GoOz6e/ZBpN2e2aGinHOr4mYmXb4Iu//r66fFB5VONNSoJMi/iA85hqus+Q378NdcT2
2ALVLu9K73XuBfB+OpNPNxgn1kpqA4XYyHcj8C47Esx16v6XGxGX5+WMH5oFtY+5jrt9LXhI/zIy
9fjcouxaK6j9zYwas8euyE3k574og8A/iLXeWiNTPDtSS7OIV4YnUXARF3SYpwyXxfr2qZ5iZPB6
2/0bc0W8FJkPJ0FEdmAbk3Cw+8dXtPA/3xOGnoaTRMRcdgE0VRQlTthtrrkXFBixom/SX9j22q0g
Ka4oneV0MkrndNK8yzndTGRpmfqtiKIv9HhfzwCINkkjCOIfLQvUQxPcKt9Wx8eRub5i7qxw9Y38
Sv4CTkvHlrnbRmBdQp+I4K1jY7AtE9vkQEqUsFJALu55UZw1EKLodxcO0aHhMgHeUxfZHxFRrOXD
qLvSNcj3TzoCAu5xt3gYrP5G/uRtOSTKoAZzYaEtXJqLcCfRl/o2FgiOGMZ0wt93gEDJbLlEeCyI
6gvQMvB7iKhgOxmczfMjCNRuZgI3hf8zaMkUq5V47mTR9lpKy+R3HPpPt6uvpWt0kkW9myt7ISQQ
NuiEi7OPpZqQBdpdjb1/vuwI3WRz3Lup1RAne4gdtnVJl/+LaS5V87c51XEtaFf5COvcenaf6dEA
Xj5VexLSDIcWUas3gmnhk0/Px5YgdPWgtMP3epGkuetvIQcNtNmn3cBPrVcNzZL+MOHHXdrWzWw6
nD4dyJvBMTszLZ7oJJEuOMO1kyvgyGniB6BKeb4UbDX9KZAMpUp3ffTA2RPMI0nrnVXP4WAR7lD6
jcCnIqmWZc3Hz+d17QKgQJQ8kXkzSLKbbM+1sI68MXCKIsNRDt0LKZIbIGeOAp2diPmAlJVhbfib
kJO7WxnkH0wZvUGHBchohvHUqNuKlqqTxq7FGRR73vX76PvnIqJYbJrxqIK1EKFg/A0LB2ZUvXMp
gozfAFl3s/xIGJioAlhToXjuDvygp8ZdO1GRbv8jOjsqjyqIzlG5wxTBXp9GrunkRZ+TAdwYgiY/
J4iO0FTe2lLSXx9xN8GgKtAncOjeO9wSRc8NPQNo0VOZHyhTAZeicZSY2PTkmhn2YUqgBhE551d+
2xTcoL699AE5ZShMnAVtiP5InjnPpoOZTkJKhUce4rYm98GJzDpU83Wk2ckOyZXUKaOg2XR0V4st
exPwpgDhzTFGnVSDXKYT9yssquPU2OkGR8npI2ZNAF3v7QU5ftvG2M53YVKSJnqPjKYaDbO2j0+Q
4tmyhyvD50A/a3KZuyX+J9Wz1IBxM1lIw70pS1I+8xMieatdRZSyCxGkd33QKmFAQxwv1zKSIYdY
lMpUMzVWZTb4E7B3l03rb/MtPajIPK3Dn6GAPyGtN+BcKvWxssb+FUnS39ChflKwOqJtUfm0P8Ck
XjaPEku53Yl872lrpmaYYm9riAB47IpofVPA8zRR7bLx0NXS6Hym+y+f3ebgNDjCBM/yuzcr4OLw
7MTWHe374Y5Fx0EQh/qc8UiI+cC6E8mq22b7/U2j9p/nZO/6E8I3+amn5AmsIJVg6HtZdlm4prDD
d6ofIFS45EhB4oSerk+oCchHFbFQutzF9GihIehYm00SbMdsa2DS2xN05KNDzVYhDpQtGFrzwmQ9
NUficu4OavImynQ32uIa+pOLF6L8z6OqKPyIYA9ngpJ9VCdiTBZ1Rnw6AMm4cvkOCM2MO30Y7KVx
NZuHSpnlP0s+imr1Me9+/cbN6P9o5bYBn/1mZHuG4yaMR0VD2POrASTD5Rko5QzOHVMREhDdUtgH
hh0c9qgpkPXtW131iSp/YRwwIOm2yU2K151UlEpUSYowIelwfnKQMav89yWGtL/aPLWQ4+D5On0r
iou1CLdkZpQypbbZ9NSFjRB2PtxW76GneTVNhuAPvSc9lbYyxxVAX6UzTZVDTkjJjMKNphsEnUYf
SSB2SZmsKD+eVn2cUl67sZdmedRIXgGA2n5Q57E9xmPdkJwwj1SqIaWrweso1BxkiCNl56wJsy9f
48O7cmnwXltcwQHx43e/uUPzC4Dm4YGU3bQVuTteeKfcBryoZFYRL1weS7nThU3rz4SG+id7WEZN
bP+7PqJ33yVvx12MTK8BsAbN2/vLRei2pt7bposzPpVAc5V8TQ285IEIkWVbvvz78SdI9wy2ysjP
AbVWv5KObphkqByjWSprvJbbPNkDb/u78qTqY3gJfI1TdQ38hseo5NkNyWqarVVWgFcW6JKP65EI
X+HZifaLLWKuMRahMOlZMUBIHhr+MEIVYCNEnsOM8Sgj0RiApbybDU4sd8GbAA5obN03fqm9Jktc
pNCatqnAQVgiqltj2rfWvnTzq6KxGLrPiU9F4l6aBpKM+HKu08XnTe3QnOt/UNXy5mmyRM7XC5q1
IJlwHGMBv30uBOZOW7hoMUZzmZfsIigNJq6Z3I+jLcW7zf62VaFSkqHvKIu5vVQZ08aJ9OeiyA3W
54C70ptbysJKu97MntJOsZLLeszm7cbUguhEXAALLH8m2HGmJ9WWjA7wU9+gJGEwiypvNgsV8r8F
xHGxjEZruHrd8DUEupRb77nAy06m9MMjkFq0FmKKGO+//+FYIx4aaU8SCgAvkTe+iCotkCoRRSH7
RbSCK10rUt/Sxgs/RwP6m9oU9aAPTKJm+j0pl2dk5N8LsUz0g/g6Y5bi1XF5dE8tSgkBnIjnApOv
i5AF/xD8TLu8Q+LPG6qEvXUPdBdO7zY7CrJlQyliBlpsiZXgtDwwRqwMOCgMtShjSLiHeZsYeP+l
nIpwV9dfgLqlNtzRZhGnWYW73c6pbm95jkuQK8E1s1RarWkERELKGmd5P/nkz4JeCTyeUGu32he0
nQ3zCujaoLVrNBvRMjgNr4p6vjz7veI/VRtyB5k3jl9mrYXEjLPsj5l1hQF2Yg8tBdqG75FbGhMT
TUzezkxcZuvY2V8aaNR4cNL1nrIRXphVhuu1g8+0o3PobWoG2Cv/ALNVEan1CGAo2LfmUKwUMkFj
Ifj9xU/My11brskzZ3BinEvvKcy3Vc93Mv/jE+LcmhM+vEWDU/0HUB4qRP0IAZH6sSp0sqi3mIj8
lCzn3ThuKZfqiKfWJbfsaYG54ej/VUARibjMIpCW8ALOZ7pjEz17fWgnmjNwhW5TlYD8iIBGTspO
0mlXsRgKXuc5NJLD4TDIaF8aND63ZOIE79XL2royfElAArfbaCT3+6AbItcAo3XfQNmdRtfp1pzA
XM+OOpz9Dhrxo20OjK0yZaw6jex1Tiff7Q9Xwf0oJzywUky6gb+wLD12wOXh1U+6n5FAp1rTGoEU
uZ82hfmVrs0/9FVH2ff78wwAMm9AgYzUO9DAoYiD0T6+EaNvb00yAPLcIzI0gAbQvfr5mvsHnq6n
OE19gldAxNJLE4TiCIeejfLcTXNOJAlQdaOPfPUaK52jQkJGEgkEa36IZK2FluB1kLezYz1uoCtE
KLHDJjmA7WHmhSVT1C2YOExCtjYnGxISBLqwHD5DYm9y5SBCSk86osSvZkaani99eIju26YFvsQk
JGGUyyotuDlLc0T5oTSVJIGoNbRN0Ur3cRCS4HrrUILI5C9OurXNTW6Dc/+RR9ai8bVCzU49C3Nr
pZFjkuWh7xqwYmzaYQyBoP5WVLmoY2s9M3LC4Vdf5sm7ZkdzZDSelcGsi0SulW1eH0FL5XmMuLwz
yI8pXEAxSwlfCE0uwXEaX6LGCHSVfgHlO274q2rztjCEbadG5RM1oFzPS8fnT94fOxoZxTfZltAC
Ox2whnePy6vPXleU6PBtsBLOVEvShL94XezA9lx3mGJQApG29qqDsD1t9DWszLVnQ804bKx9+xnF
E9zVjjoS/C0wKOJBDjmYF2JDJQFFTrbpWTl1RlHIqeXPoAonfbYTwOunEPLjYpvtvukdSUGfWc9d
1Xzhf8UtpSa24l8FAeOCeFneOnTs8o0XDT9gPWLb0q15BvlYOQ/eZWHJtP/jsZi03mdFgGGmB1xo
2fNuck3JvlZfHLLfZdr4k438pOfemUj2lEl7vAmkUUcKMIuLLJ9YANIkJJ34mOCEy3WEH/JTXnl5
3X9FVLGMznBeLxZu6I1Fw5cEjIrTKsXyxp4YO4lL68euGIqBENtMgn/mCzVDaggMOmXkly5K4pp4
C4XH8LHge+CbAc9SsBX4UZU577FyJxDivYHn4rMbIwMY3k9X0Hq1W7+HfHWjgiX3yR8+cdHQZDTH
AMsFUXYO7CYh9XJ/3OTTztqYzivrxnEj+fDjOK95ICCCa/P/7OkowlcZLoyc9jxRXYla5Lzv8W1D
VH3OBPCIxWhSJpvMGZKAXWHvlpY0xDxvNTQIYaqccHxSV0Kf1RmLio4j58qi3NHmJbfMbBbyHWUY
T9AuFVmmZoFxJDrDbBDiySwog/8OSaw8NkZ7avA5Gz0+y8MSdRQdRdslKEkxi6NqmsqS4oUOmkyA
v5bL/4YFZg6MTiiLxsRp8sJ/XchDaf7OGok4LDp7fObTNSAU3j1qWhoOzo73bD1Xb0t14Qla/vRO
wN1prBri3N67AzQh/0Nnuock+6J2jau17VxmaM9Gr5Fld3WqWyzm2PywYsw0L2fhMXhXm3x8PC3r
3t7DkE0ZUyckI+q0HRTmmTjj8kV93Iweqn/Z0QsPxYT/9f0Figc+QPm2Q+vtVU6cWbkypt1G7HVi
3ONPWXRFK8JVad3obtLGd8yjDJ2dZIYvaRBpBjMgCJsYN+MhB+I5xJ7k7kYyzUyIQu1cz8RiICBH
rNQaXEGmYXlzlc7lgldE0tAGwrDk087et0oQOonTKmyIKLozMikTbOgbBjGSghRbWaXm+iFYMDxQ
iiVdVmrm39UqAIfQFXGLXgU0mKH4nBmsjRZC52NiBElexSEDVGGTYJkI/nm3p2FiBOW/3YNtQKWY
ttgN4P3UTmlI9ETWdhWF9nLHVYNJ2DsLzTgKWRKOtxKrPjcQjs1NQ4573QC9OUDLnS21HMAV/CdK
3UV0BbO+AoqcoILtz/LYl021HvoXoChHG+NCWKTMOpsHrVOPolo5p5ikjsctHv8cCajZ5rPIsqs5
lpJK2qxZgbNJ8sCqdXy/qrP2gRJuQjEGeCjETGeMGu0Eqjbr4yBtiurZk/mxFePgzxQ7sSs+jUZT
WEvdCjYXBC9ZOAzQ6vNAUWEKmWh4l53uXcwXklYhErrOpfSHmyG6kcz8JMvOoYujnChWykFq4Avl
kyy0Umv8L9I+nwp/op6hCt3Ol8N5ExgRrRbMsax9TQretHBP2Mk979y7vHreLyn6jQ3TYgNROfxt
6mNES9gF4T4ixkmKU0zbDrML5Q1ITtAPpGLjPsUDbB9ZvJCVX9uK21uvs0QIogwuUL2y3wW+VSlw
xZrz3vixr4OnpwMBk+qrR7aSR0GY7mzMIJwF3Ty8AtwrPgn062ZHN7+2K1j+v5YCPnWUBYP7xyqe
RyybEHpyAMSoKLcBFukq6BxcBOmWZXX2k/Pb9bh09GFxRH+gDKQucoNRbBVBR6/IcVt184Zyq7GA
cO3IBHZFiyi3MUL7SfHDqnfUNH/5BDcIAZQK0HAHrE9eTN/sWH+jSjE//9NQMxP3D9jtdrTGv9bF
Qi6eB5nD0o08oPvXmltCDFps1RqvG57kDerzh046U+MrX0RlsjXELKuBjq1MBiZneDp6i0oJiHxq
A3pTLu5+aNsghj9mDgSEDEK9a50BmG7bQIc3h22yCKZIWk6N5KmDu4xhzzV5H6+MBORLs9bwVAbR
hGLFAjAlQ/D387cAJxnWWit/fuYjjx60Saw0ibr8syeNuDgxk3SApOtgdmFfkflOAen0+Sc00Z1I
hjaj+Bo5GhsYKMA3KgfUa6hXWN7HMx18GAKfGG33V5VuWmbvOQuTUxkD4xDEFTsj0HPO0N4kmMW4
c69scjJ3kzsq4BkFy0eisZd44pjMdYfcgGbeuMt/ag5sWuea+bzoyGkQXKn6Q1OzZj0pkj9JFbsE
wP4mg5dB4t5BkjgoBu/kOp+pX1HEEixi0plfVOO5a3SkajdqR5mGwVZY4MZdkSL/TXT3LXnmNUcB
5RqVroXzCuE7waF1clcfBmuXrdmYoohTXRGjmk2FU2C7Yz7w4Tidqp6Wb2N9OFiinIsRvsS1s+oB
ZtFNfTVbtRgJ2TqakLpCWgSHYbW6yKithgvK/Jq1llfkOZWlFHwXZGboOAtcTQ1cp5iOWzEavFEV
Vq5i72eixNYNi6g4YL0iNj8ZiC8Q/v1FJC1LcFVTUFkAm3H16YPVXXSeqhjh9oM1y57Pib2ZPUSK
uWpyiQN7DbIVGX+ZkCnDxPt5cgFz5y6oFCmBIwaE5aSR9r9SbDw7QzzTzXFem0HKLTUM3YxJ8eGi
InNnIHlECBU6v9OtmbRohANSY2iEbrAJr4q3Ah6DzD8jfo2xmQygwdmNaQ3cur8GnU/BONOzV7ob
IuByEor72HbO+hQBXpOCw+XkbJBYN0yZocZx0EfJC9167aR9GEanEq4NinFrJKDVx6GJZsn0a7us
N9uJ6wVRw5hlyqwZMzZfCI7VKQmxCK70EHYCisMr8JLdChyAHHrkEn7ppHnzEv4YQUBnF97ExDo1
TGDcC25rl2/DblUlpKPNzS1VNuwt1KeWSjz7f8AEs8qPz+bTzGoxsaFJlMuGXvcfVAsNUsM8KD/0
aklZbON86TZ6yCSZWwXDTY4Imq4uWKy2wU6+1w+HJq+Oz6xbpdCpylsu3xrylFXrT01SrKdN3ki2
5uum42fbprS0y2T2R+D46nzyFbywEOJUGQTJJTIr8yk8W6IwDL3+TYuYn93xoZAuR5YbKu4D99EU
Zb2AF57w92a0IpQXFsc3TMdtkt/yv5Fe3cIboA1AolIkEnFe2MFRYu6mqAz4oBpmt5xe+ZzhQq8X
yO6pXg2Kr0UoX8kKLT0KG3ZjWYe460Vm9E6rQ6N3S/lRP2raPZgvRerwZNgJohNWCZMSoGN26WvB
uFAjjf/NPk5bx9m7ZM4ObsfqR3autZSKD7v0XrejN14dNEhtzPxByZxVdiD8a0SDYl0WyVpjEIrJ
stcgmVDEJl/Z6IODUE91CCXcCu5zGFBffTaTn6wFg0hO4YAd6s2+mhE1unBM71WVENquL37Gj7b+
aUyQruxENzoxSqTMzO1lks9PBb6faNCEatEwiCoc+BESDlwKuwtWBSJjAXPbdF0FpM+0KSyZ8DiQ
yRkTGE7YNcTtGRbkCaSJ3eiFCJQ1zgiYNGPb4oSL9ayV3Y/ahpz8x2/r28w279HDW27kHaoSoND8
tohvDDuHhwKgVCgEWJKzI0cIC/Kbd6nb5r4gLhLIlTTHn0xTZDd4QCt1wZ04vF1m6i0XHmgqSx6D
DKVLda1R+ZIqzmVvOFlmTx7Is/aRpqWLTyPu8LVHutiY5yCsdecH2s4I/eHBDIyBv/feBiN1B0Vh
trIlsAXbsKpo5HYfxpXeL7aLMNzGVJTDEwNzGeb/KoQfmIsWKGLFipKdP3iz1hErb6qa/PYv9DAo
rc2806xIdjZ54cmdROfT530m7CvJcB/2W8uprQ8/dKtP6R7Ut27Egi505C/hvcnju0cXQPVly/Jr
TQcgiumZmBkFwqE/pUNzYWSKovHemATNoemrSpMP7VYfAD0LiZM1uLCgUw25lzpmv//s+sSsZ+h1
PD6trF8O7m/NGcA5W8QWoDBmEcUl9hTvWLWjnf7bhmzQozPAMPsmhiVuGpf/ACtzGVyW2vf/ecW9
kzfdx+vNaDO4p1Ap71w81OF7TMChK9pZWt2SiPVqDUTgefsPnOVZz4+RoeZ7c/iPPZfIeSjDPPAD
E79k1JVdtUTP3+2v2VjT6F/n5FOh2rYNGQKbOpucTjbpkFq0GLDHDFD1+sHzDHR3Bxtyia0IbrHb
t3AxbNF5z7f1oyB4Sgg5l8NBbQPheDMDO20mjxSWZDl3Ye19NLjpKDt8m6I4wL0kJqMiyWlS5dU2
z+cCzidNnM2kNO/f2VyR30r0whVX8voU8l4PpxYloIb9kDcvU4VxLKjul7eFo25le65M5HW7Qh+j
BR9KGQUsGk2bB6t3an+yadDgxih7p+oqUdXGgrd/kW5Bvl2JNVWWjsUfcO1+qY2jxq+0tbRfHdRD
uJXojyOs+jgxjYqQ1s9ggFxO7cgSbBzfAmFICgxnXGPxYpUY66etadR5onkuOCaeXDzjI1tavzZI
pfghkt9JrZ9V6H7f+bOjdLBlxE6+xORuwfak8YlM7Pho1O/03Mu8euwpIbpP6/B+sZvDXthqmtPG
6CaWzP5YJCmJOYvcWAeNWoKmdpSVHi9iCawgPVwIgypCzfT4ZeJASbBKreD6KC5n7CM7d7zHx0f2
J5wiRfXPOGI82fNsZTkTw7r9mwaAztHo8zJBkpjP58uJ1JPdKez44bNNThvejd3eAnfY27BL0ztS
kMKlsOHkd2Ow8F3EgGtctxCO0SNqTV9Wr6PVm5CLK8ZA73WUfoGqAbrD1oB8fdRrRJV1NGDRokAu
hLQUhimocTXomzhItIYhDPMegcXRuU0BEYjqasTd/jXrx/M2UtCmRyU9Hjo5sZRGM3h79BBVy3Z8
GPjgw0xaJJlz0W+L4WPBmrABx8qIwXY6RHq8yDbjB8blA8cmq9IQyS4qYV56pxSJX4NsbAeaSMOQ
59u8Ia82/8z5NNZz9toCtqjf/VU1xBHJnT8bGGfeFDpZ9xkRUixA54lfK3VzzQeJqkGmBKMWAwPX
H3AD/UopyStm+3hEjpwv3Oum1XdlAysAnz4Qd01s9YfWHIUr+iiqlbPEM3i7JBFjhddX7vDqsnUJ
QlvIE3XKCDwNyZTZM5ud6lxA49Iyn9vjdJtfuzYUsvRbXneiVdj3109Z7J3v0GC7LuYWgq7kJh++
tgFgih122a5tQ4fIEPfsErClo77szvCuoPR6xn+WeiYCOycY8qKW4wfVyo8MqVsFJJzs+zF/KycT
65qaCCOYjCi0fQgOQ8N86SQAMWGOdhm5B7cvtdJBo2wR+OZU+ULKri1rar5dnqV7imJiuK0s6CGv
ANlKp06ByDipfkUW1/qN9+oaQERK4SryFiFhSVhL45fpvfGnzgMDvWAL7UqsfHWHPFmWKWd5gV9T
39yIvlEmO40dVAQGT0+Tn+NrKZQ5RdgURECtaCWIAvZy0rI0d4c4RWDhTEPtLLdDd1PE71kmPGRO
Cj4eKGh1bS8lU2WFtMF5YT7zgPH9IjDavHyMqPGxrcLoUFkoWRgZibE/LYrE33WQdDbfYjM+ciir
Mu0o+nNlk1xxAXPyYOcpXytmf83FKB64INP9/e85MvsYJG4NEPp8lJQ9Dy2HCnFPK47L/ieNQuvb
DUbJlomkuhrqhRLKug/u7zLW0UD1VZnnFQtybZZTPe5cRSq1upcFO6YyxNqDLsYFcNJezq+Nk/Ib
FzPIdZYqT0wRbe/bkAzbLyycumgVGgowBGLKhWfyGO5pzQqN3pljv+8JV75HXOLSnNq3SU69R5WD
URJznJxMvpHcW/2opJS+53IZ0FAp2j7W6kySv8lqxenr/kTk8jXITSy5hIty+ZVeftdJxXJhw4Mw
8j9q0O41rfHxYKVEqmfbJD0DHJzHBhjQmPYjsmj7GNZlfnuCGBuEF31gVfczEB8TdDIo9IyFWVSo
7rkcgWzePMW5XGsPlN6vsujPJktF8Sc/KRU+YyHF/wKcnoSCFI0DRwZP1FhKphZ+cAZTZaeNN3X9
LdF4XfsViIb+BZpeqFo2ExOQc4m7vO7hB9d/VdmUGkYk3t84f0tyuekkpmya7ruYUL+CrrqiRekE
gBNX+ss6mLNqDW8mHraoONIPayPirpj0j48GxiIRHIXhk4FUpUKZZ7ZJSVYMOw2WYfsUAsovqhm5
9kbaj01b9iVxe161bATSAfsOgiDX1wT1HQdBThKyr5i2VQaSxSklaHKm06OYxdx34LzZBBRGYQDy
W0btXE3qnVwtRE/0LT6DT/hVnFWnYGdStxlHfZgP7ARlGfXScI3Kep5OZf8IyaJ+F2oDnlwT4Y/Y
a8tpd3O8gI9BwmaUyndthwhdJ7Yc6GJhaiGZ86oy2xTiwfVEzmpvyEXuTY6qLEyCFijCVOId8P2U
IYjFNRALDOi7j2YfCts9v78UjoDrzDNTECtIlAqAQN1EIHONjV+gbDHaVslWB3x9ZDGCGSiPQ7mw
xLRah2IglEeWPbQISXakNB4fguE2KmyAbatFzQX++tn0nCCxY9AtnXDBqY3SFjH1QTXl3MR2HHZj
bVgoL4oBi8C4tdBaqQ+HvBWzkCwJ9NFNY0/+OX1t7fXm5Isw6VTbBVHIKPK3fYq4nIlRZ+04fppl
WKhat+yV7ptxkkbQmC7rRKtYhLMciWWOCcSyoKPQhJ2z5f3yX5M/uxPCLrX5T/LppGemugqdVTpw
IrCGWgNMWI/EHL8rX/Nbh7l8h5DLbs/rj96vVum266MgXrNq3g/tmQK2UqQm34BpvqdgpD64Ivvu
LsoSCHLlDqx8h1JsaaSeZupfTGrKavnE00QAwrInIeY81gXahx9ukytBsgiMzTwP7w1Rdv827rQt
fyI2MSSTQJULWPN15/zvK8AqDsy5C+nxSDZwGjVZNNHxNgD4H9Q1FCR61L8XcbTDnJ3d9JBhCCGf
YjvgyiXH0Oe+n0sAoF+rppO49JMRyJSMGbmAbhN6L5Tvdd767TC1+k+4sKCOgO6STJbSyqxj9RqY
MJl6t9Hm6gNrwiCyk3768SCTX5y3Kj4cTWbV8oll/VIEL/kIOWprbeB70X5fGAbCl/c0F5NoVSEw
BT7PCoeu5Vm7zZxewf3Wjnpnq7NXb6XJNttiHu/Pb+aqPnwS1yAmGWd6U8hPvN3zlY/uzRZ5mykw
GTeSUtyxrir8pjKRHYKs3iFRe0Qxv92eO5KjuG35Px3upWYv3cyMPoxxFlwjxXVYoJLaxo3dNg/q
RJ2XqEJlmCJw3nwLYF88iwGZOUt9TjyHXZx8LJBtOe6kHzNNY96dTCADn0JvfTcFmg1devK0qnj6
pLI369kxIfTW319uxEUOOAeOXFTSKU1o9Vz64Q10ZByCQpWnZOsW6EviVWPhSMryFoRbw5GGoTni
Kmai5p2nROmaEZDKFIzDPvCe+ayLIOYKLB4rHm6OrYRA9MtuDU/OJ4OC/iYsuJZwr0jyQ1jxElpj
QgdRt+HgzuBRz4m5Z1L8qPjo1n8BhFLjcxHR5vdBVeU6PylsRpOyM7InVh3sBbIwwSRXN03RPPXu
/CTRXPzo1zguPRsZGpH1417Zh9wCzKkY2QDe3y/3ov6s3UWr7uHC3GLU8Po1pnjXiJvieI8yN+bw
z1MAwWRs93hQfc6scPLsXKEkdj7mMIT0SDRgNPFQ3AjsBG8AQQeqgEm5LJw4aymGkBmEJfCkBUtv
vWwYe4fLIaVNCJXZfrkDAYybB6skadVfEJI7nQPlDBJY4C60NExRDozFmnkWxqLCabDi/X9r11o8
jtoQuz+vxXinKKKxCFVThMynV19T7pRvjes7EW0h8Pite0VaZC50Im0oFULAlOYAW566oEfoW1Zd
4w94J2kTc5rZBSIvjNqTgcYzWMQ/KLhv+doNwALTKzHDNYtS4g9ysdfk3N4W2zOsdE+BA68e7Eks
cfDbUy/MeeYYE86xi88BJ4lv4oLvlAsynrrfOcZUpa/dh2F57tX24pzO9sW5+vICoMILDkdvipmm
8zRbDBwicVpDSMR1BPfHM0jjIIGnsfhzS/1pLX3+KCckW5fgEv4n2v6ncify5KuD3zfBKGqgn86E
c9SFWPQX8jUcLt2j7YQandfpaf2cYNjsD3lB5pWXEK4iOW3XmMrvsHbCpl/vLSM2beH0xRybgFvX
qTtS4bkQO8QiIdOo0ujvGuKg9+PrB0OyV8IBL5xUmDTwk9OAxJmADf33Mco43gSy/E4T2p0w4vl6
XB/wCLDZWe3b6PWynb5tvHUZ4XcVpyjeYpLOil4HcvKSUACsF2a3Or0MJxTEQDoml+jo2LZTVsgB
GYwrqIePqLyhjphcaNGiUz3Q/nXhV5Q8DmjXtZTNLRkrUwFx5dcHXjdO7W+tiJk/UkU0cstEmL88
/D/T+hIdcmFgTIBtGN60nSToxOxPoJ6gE4m+qYMr6uvYEKGnFv6F+8iK6tsZwY7lMA8zw5GAUihD
j4jB3H25WgOfHpN+aWU0MMJDI6AGQ8TY2Ru7V7bXSYrLjAo53ElaCBYRUIqAJFbYW1yFX4+hIhO6
uV9TXHXy5WEIWizIrVm4jU9kfHO9zQcC+WWmSEBk6aFR4lp9VeOv6iq5yWJ1Y0WFqLjYeFNPW33u
YfXuxi+Dzoha+IcubU2NVybcGXkM/8ONqd2DDK06rK7pUmiho/7kQGDfXHHzL1vcq+0lbis3ZWlx
F1JR/Pqoc8KhaUoNPrlOw6jPOn8sk+e/OTtIt1j+7s8Tv9S2rvcWcyak1gwyC7hFIg9khbHqTZhE
87CwQl9LK9+BEsCrR4nEdZj6xh7PnLhWVUOh5mnpKFsbdqXQgPb6jOSSTE4vSxMrlYp/ouIar2yV
SCXhqWepu8If9YiPfch8qMRtHENTY3FWIZqig1oVB1CFLXzKMxZx7ZdgjTt8HzOmdprwNOE2N5rs
cAKvl3IlKywQCjSi6uijv3emdWP2a4uGCdkM/hgAsxlTU2rt840BZGd+o0KFQPV4fjK3h4qiiHeq
4UCFYkcnewwGfLRDnGGyIIWPHhzp1tyDjlr+WDIYM3qHE6YKDzY7R1q9bZsX/OtnXdCfdjDBOQMz
UM5OS30QNZv8Aerlx8I4ktot3kLT3OURgP+QLF9xOQ4hX2K1zaJ0UzVAspSIVGZeO+S9SUZPrl98
SdGSsLePxywv+7Gfz4sK2yrp1xE11Hljnees97gkWRfVvOIsjVmfxDqVEz/HuBa2cYUZuYRLEFNy
hqvkdlD5gFK7JbNSliHVA7JHRKGvr7KStHHMm88txcYkTRr7HAttFxyknfqhvT4vcVsevQXiiMWe
2LWvdATN8lPxQwLPuVlQL2zWt6yrZeoz274KgZuIjcUep12SupP7ueR99XFHEB+iKSEHssSr5FO4
vrLtAHTCf+PpV6oe6iSjAzYy3Fh/d51+zJ4paVJbxlO+kzAp/iGcZTqkWuRqBJOcczcwQ8JxkyGt
ocm8FUrUHPgVY/V2k8ytn3nfFQyAaBNGIOiulfdZL+shunwhO3mXMcGJ1bOUYMxbJY1ltY9wjM1M
8emwqfUmHQngy0nIF/qHQVHGTCGsWVmQnRsag1zPeFBepUeYyQBkVbnIcbXCtE4eOR5v5exTIDGl
al4GKOX61GhNNr1gmbA7Zz78jR8nhA9KxT6X+VvF8X9WxJ4bEAUY2xaaTVU3wy8Eplqt1Kmg7/tS
r/dGJ2fuTIVWpeL03+ejU9/67d4OoI3LRwvoIfGlEvrwqJansi0Kh/xZihOpmMlFculYPcVpC2rx
n0F6dAESDnHjc09cLwYbvR64eV98M9qmsGPM8NaMUvk4F5TsmaUnapjcIg7Hm/2na5x9SNYLzvaA
wOacznyVGQRnd+AI8h4bBLbrL3bQkPlI7XtnUQpwR0kzUM1R5hDieYGOPo3lYFT97oRLyzq9jX0V
VRZ+VGU9YydYggS/YV/uWZp4lhWG4LtWtfuWdvwkYO6TilHbK8ke9GRX+xj6mZXeBss5/U+QYuur
g7leR6bLSivUnsNXMzB36qJA74YwCjdtnW/T6rnFriWu2eziXhTxdPIelIL1ytGyz93jFvmDCO0i
FBK3i02Rt6HdQ5Jw8CMYYXJYAjzVkoh0PJ3W2NQmOCyHux36Dc0a0D6WBwa1bUooHVsJSQDu2mIK
26DoZNdql50kJZirMJvG1nLQOUrXo4iRTw8ZvG7sKFVLgjHwWihrab9NQdH2PyLUbvofKa7xQnFL
M1akY8WmqSFavLOM5suTGG3EjP/5hQXRyNn7YD/tXaov7WyYTbnbjnVYdipbIFQElymQUcOupRRB
S11ELO/phfN/zjyS6+zfROrqiBUQ2Ro+CpPDRnHNFgymRiLFpBWPQMcCJj6aaqCfJYWawf7WyQik
hPLZ7CGRBOwAGQH6+ze1nmMtixReqpXaxFsq97thyCaoPFbDQAQ7H38AqM+DNyZBtpCAB063zHGk
pGpEsiUex8aAodSX0tALZxcWBKIgO9JGxEpjakDyQSyCNiSRL+7hf0kJkmwVX9qgULFMmII7gvW8
xnicWMGEuvS3bfeW7II8gBQT6QFFVDscG0afT9WdwUzoAdL/OHd7EsA2OkMK5Qa/bErf3+IowwdO
JHPEFTQIbMgtWjoo2t8WawA26TCPYXp0R5FoNv6jcuW/qrhQRraZkoJoEXHtHEkwDie9ZXqfjZ6f
one8kSUE/bGqwshkK2KZdkeu4QwuFffrb/IA6DruJCKU42NPznLO97144+iKVZB5ZmrlZldW32KO
Bw92BKOVfHzPM47VtZTlIhssEvuC2vWls8zku3Sv5g9onSsSauvcMxKNVFQwSF40Ye4aS09cjurx
hqT6JMM7BqyrQtwoBJNkVaqMupuC3AOM9+wD5JsIyDct8N2B7eH1lqsj4/SY2LtAAeWkyqzO63YL
ua7o4sWT5+o7+WLfyDgdzjV7sJQ2kZNKr0IvzeoJ3vXuNbTv9BAihGjSpvdHamvvucAEOL9Ohzlh
LRuupWOs9Keyffw5R72/3rB4nN0xFB8GnsWAER10EFvLm5j1+BzMA8cxqoz50Qvn2sm+vZblzAt2
hdgZLaQOAHYjiQxsfy/NDofZxwiSIhpDiT0aecJ83IDbIhNPlCvLJfQX4ZOSTYwIVfWDqyp7AiRA
zQEH0QAzcxl+0JZNjuFziwNsPpIpNw1ybXicxjRwa1ccyE9N+AOUW1I65I6jB7F3yluSFDlBhCwK
jNW0nWz/B1fzvwCdIqIdvXiY/mdg/kGcJ2ZnhtlAyMZAuRsNnQOE5CMTqOnKNl0s7qVIYIeQrk+9
lzPAyo3RWG5ph1MfntCm02P31Ossbciv6AdlgY43Ngv8tabC+sBGVJIQGFLPhE6vXf5ikx6RXsSx
QrAvoUOnEfdqqTL8HMj9fB+I4Q6xfx7Rd+gD6nPFewcOioJihe5Iw8e84OFsue4p5x+CuM5zvdje
VtVlWzC5d7zBc6TpR6vibyvOErFzuhp/HZYt3QR89mbpDjRNbm7kjqQWFVoOtRuft4AVW1uRaZrs
S+J3nyHXEVSUfIFzEB/fdWiOrrj9BAVO2pd08ZX5EBlXMGmNivY+gGB7ftImIcKDvLU3TWU4czGu
G4hx3CJ02SagxaonzEi0f6Jy2lNRroWuVbAwuaIRn9mMw98tkWCUCfEDYbv984eCGHireXW/2N19
zb3bdxKlya0ege9/LpRh30SHCW31bRoNHOJ7gScBv+gUisGSrAhd1gAYUmhgg4gFh620dDN9MSxa
un5Fy6sl5nNvUSqcos2vgsymE2f9QQqzK6b7H3y7Mc7vKLwav7M8aywQhorW1qwo4hbQSL1Hmb/P
3gH84TxGbit1k8AoJ93XsvOs1K3+RbHrSIuxrGMHQFJWzQ0LH2AzMiYw9WcOeSmI+0xHj54SKVua
yj2WrMSJurKNK2LR1G7PmPB2XVeFApvGTj1ei2C4qOUfh9D/CoCLxPB2Vl2Epe/8bQDk+6GLHKZn
qQxrn2j4ugq+9emWyacjPTi8WKeYm7jczuBe94A3Q+O9k7/B/qAeyinVBvHVY5Ad0X8k92TSkG/I
I0WR8g8t5vZs0j13RPC+bT0nEnqLo8GxOX8R7ih1AZcNS/SFdHaeB/j0ivgAfhftPzV+e1EivfcN
26m9sh8TR/MAW2qyWzQILHOqgPRcK0Ce0hae7SwOXfWATEblUVEiXyYxGmdjw7R5T/AHuEeEtu+3
QIzzhdkFNMpMMxzEFX+gwUA+h5ue/OyuhxneOAHHeORjTgiTRpDw3MKv/YAl6RTgBhhx29dkNAUx
5W+pJK4n6kuRdy6GCioT+1mBVzuyP6wxMo0GntgJn5c0WPe3K2xJ66ADm3c90Kac0in+SFFaMceZ
ekkM1NuPeZnhUtFopZtXZBNXRxiLUL/EyVP/9j9UAccHdolyBqiKxipa5E9ebOf3PVjz921FCaPN
dudCwE5epewJqXDMfKn0T0M4bCcbLZnqz3XF61Q53pr0eCMCuRLsshiSS2HrRv9h5Ud+fMzvGFam
bOsp/8p2TbJdY070+ODnYxpvv6BkDsjyPDo00LZRklKjyV9nNBAvQorF1WrANXqyCgXIGB2mDdAZ
Hkn2vZxFLjiSZiUkVi5/+wwuaCXKKIp7pah/A6hupU6wZugeKX3PvEZFzZ9yMPmnZBZd18kNDEQZ
8h/Tmc2zuFsFt6yeEQ15OZLkXsERPNEfUbvblAqrsSfEnYWen6Fav1V0GaHdZL++P3b3UlGMT78L
05f4TeQ11EI8IKcjQTrS3wMWu32bxllC+9Ar05H/pZm5/iGqev1ECBLz/Nmhrz3wxjBmMwI06DgM
BajytI9fi9JAlGSS3oiOLr4TmO7yutr+lL7KlAyqVaBfixdbvQ3SdEHU+yTyxzbVB29suq5+Hn1q
UD8ZJXpopfgVf5sWRR4idt2iVp6LS43XyyiFF3o9puWilaapM+1M6nV8XLyX/y96M/zLdU0392ZS
cHj5GXaksa81mvyz+0M4Wz7cwBUILSDpHeJvi4o+WJAR7HeX4vxW6baJ15NycH4q0VBW3eRG3x1/
U85LU37MyrvVrUa9TajRc/3d75DtgdCHBc629gn5zvvv422EdBXFB1iQ2vQbL079GRzTnO7HAstL
z4VfnFWL4eMIwutecCzk11jhIq6QSDN5l3uLlSg2DOfk+1gcDxa+Rcq0ovtAcMdAbqBwubcakeWq
thW35vY26wTB2Vy4Yi4BO0ChyrXE3pZFodqdYwhAYdaEWkNJjJZGxiqy8DMmNl5NDmMAZB2m2qwX
ibz/+fs3hJAA3RT2JBhQG3/hI9a1R1lpnpTH+gsjc4NLzi0V/OtvCcNygLGodhO0XyNdzfwhKrYD
Y+oMm2MuhwWbNgT9dWNL6Msos40dl0PuGWXDOv07ehvSs3GU1TbKoiJh/irHkQOL43mO2CUj13gK
6/tTWBJGYneeiy4o5JZ9H09kjyezuovs7G9mrYJ4xgQ6HJA44k+KNufTCUs5dF/r/Oge+N562MB3
w55XGCmwk7qgkCjkY9z9MNELbHDnHZXW+mFI7e7rg5XLJK1akDbaNQGCum+fckfbZIU/MIXfTS4Q
cjYbecWCBbeOa6MRC0ohkWoG46ZELA4Zg4qaBXEzxOZ1xmJQIVA1lVrdoxWyYCEAdWKHhwKtfm5Q
XaKXvDeV49Shyyqhr3fKDyAhPIU35iOTxVe2zaxt937HJwOt4TS4TmXyVcQhPNoEUneRlMyoNC27
YytE+3Cj06pky3uDv4YotCKsDwB292FsaGnViF2I7xuuO1NQhh4GBXRRmmMV05hUdkeD6aIhoB5M
AMZhUzeGmX3XBQHsrVM9eERwT8zvrySmsSimxn8c6MccfVIIyr+BeZjSFlNOThp7Bdw16UitKBr1
iZD2wiDoHGLyWVySsWiYMAAuLXOvwBflgObB3NQjeagnHopqCeOswx4JvvIfZ6pgeQYOS8UzyLaa
d4QJPPKYyFYfX/qL4wcAwltIoFKLqMy9xwW8ychdkak6IHBWyPMd+JGhftUIN9bYAlxl1kYR6ObI
XcORAQSHphnSiLRwwssHr28U9FqsoLi1c3etu1VwuvLKquVeKUgja/nEGJlB5iFsUWTJ9ULn1qC8
FvqOxBz3qlVk8ltJYr0b81S6f9qYcJl7M8KE8foHKWuHMuBWd9lfW6kFiays7RlDi5kBRYASI4wA
mXn9+p2sbKcRuPvhYtzZy0x+dva1l9KDsbq2uIkgGPWdEtMB0npE3vfkoBAdNuMmgS2tFGu9J4xJ
Yyk3oNgfDjChbeTf7/JgnCld8KKusOB2XLJTZFG3BAOOnonI8AGKJ/NsgA0bX/itSMpGFnemi87o
M26U5KW27fUaEmSxWPjUOU8L34WGf+5qKADCBwa1yEiAwp6F3xL723gTYuBctePLt1c7da6gqHkp
8IShS/UiBI4jeF0xqfhcP0ToWgPy0UIdfviq7aHbrVfi0iOnMC/nWU6deypXeZnbq5eDiBzeBNN7
brzNvbZBIzdvKl41mEdK/b1W09pqlJzVDk1GoXELs0eCXD4mkR0nFNiBbrNtQIpUZXvy61WUGdSb
eunVmKJCFLJupOsxb8qLY8g/PO0ysfmlAKrzdzWdZOB7XeEgHdO8weLhVFnbvPTsTQoJR9HsRqp7
FW6Wz86SkU2dIIyV81DtTHPm8vPumX+5yE2ta/1u+2ynVEU5+7STqzwar80Ky7pD16iIb/VS68FX
2ZVuHzYRTE7+YaF6evi/Ue0CMc21CDtq+dyVbJybcQoOS0HTXP+vZqTsTkGKjJVFdQyrBX8Tboe0
+N3iwln2CK38bO9mi1lqil7BNMR9FJ9MzIcLytFli+TCZtMf62M/1vM+CZ4mMpS5eO9xEgp2Pvfp
yRiGvPjN1T/qVE4dRecWKRmu+TTem7khGZ7yHirw9aH3s3/DadCvYTFy0wH8CxA5iuZbgYbN8ROO
4Gl2IC4S23Z4h5cinMXogSnltDYebSq3mjsdj9xSvsLxQFJ2mICko4oD/AOR7yUSCXNs/5MP3ngt
PV7mDzmdRbq495Qyy/SLgEgEk+v2OUllk1OMhQq0UdqC1e9i+33nHu8goFBC9tfM8pJtRmxZT2A9
IZIuUyxRcqstmwqVDPMvYSZlucPW1bMQ2kg/nodwmDTM7kIPOOK9fMdDNTOXtWK58dbEMAKVI4fO
pGilIlIGG/V/GIoLIxbtPprSxC+ElmgEstKH/QFQHVbj05e83Xnim4zO7ljw6eALLRGpOrKFZ0X/
2nrNbE+wH0HbflM8kdMpWAXLSy0yBeR5nwejTlnK664l4oMnqbfadzcAqv0ozjJASCEhc1LgR5lX
ePPsqVphws1RBxg1J4xj4XAJUaEiyxu0n+hvwV4BYiGSggGlAQsz6stHEU+A3pSA7gLnDq3JA7Wf
l2Iwbwo0IW1FtsWRaNMVCOa8Bu4obiriLH4k2ddxdrPuH/7dHEiQ4+4MZxiNggfSEDDRGFC2kEkv
y5WaQLG2kLJ2iskpT/7BPhefWSolJSJV+/6tAXOKFMqm0CMayD8wmQ2YsB5qMH0Vgsjhsq5HYdw9
23Iul/ob2DfR7kjLhA1GG5CpZQnEhRmSBTZMaMaCSid9r86sJHClOKtoD01GTKkQrfNmxf2wPrHB
haEza4JopNtfANhfpx++Ua9hcZtxxT2LVhPGmuhdpNWNDwp6lOVW+psX2NAdjjUG+CmeJCj44nJt
NQHBnA968oH7DZPsQQ+bYoAY6Habdrv1DgDu1kLnJprUgfLd03q1KI7+/deU01yRZXmGNqXNVKp6
210jK97MWjn9AW5TI9NmufXLfNAPIMMz6Jsw4BvAKSd97q4xM+cbhp6qHSjaA2B51ziFxutVd/Pf
9AYITiqmTXVdLHvZoptmpYeKPlcJLksQEI075qGPhEvwWDDyZnSlq3gkcLioOzv1/YrLBc0IVSVy
uw9rlnErckXdTP1vjp3UoaziiOJSbx1AzfiCcAxZ2EkUb9xmOqa5HQbCIYsfOZ1pomrth5wu3Zl7
ySvGB+Pb+63oFS0lcwWewX/vzztxcv1cS8kyHxPB07BmwUR9TvoSASlCI2vr6wdzV8ade9aSu6Bz
Uqnwn9ajQ/mJSP/fNyiPFiOdYhktAXzDquzrxPNILpI7EPOSxLXUipXeeamKFgcMDOtvDVEbj1ce
wFflkMFGxdtRj5MPmqBv3lUxso8Cctu/mN3pKSIOsv8FZgZAniZMecxfO54nNqHCpiG79OdoL3JI
F4fjYEtELQJBJevbks2+Zh2cYl1ZZVNIyC9sgv2AGTnGfbFSGXIsEsciGnfunYZ5t/1zF4XHd1tY
zIvsxJf5VtGoWXyYlxWZNhmtmwR3Jyezu2Fv0gpjapRBp2tFpMojTcf+0m/bBRa6v+FbxBL6B8WS
+tSnWDCdIYIaiX652oHu/Zh6XbdHxYhaQxcUOh/MVPQBPWS3Tgj24athAZViy5XkE4lGHXz6iR4M
MmqHdCSy4E3UqM5ktPqIbPnKXWdUpVX94DwHCuUKWRvLLx3lBEf/39W0nrNKKHnm7IRMZJB6w2+K
pyDeCF8itW0HFleDi6lCIXpIhBRctUttt6FVCks2X/hLElOhqGp4XbyljUPfDkMBY1p4BggKoNqt
9/NwZNL/oSx54k8PVGMxAA7SaLn4qtaaBGQSagEM2GC/LF/ThQT/mNuCOyy08iqEyEcjLLwkabZE
3fMxb5iHDNC8OaBsze/yuZNFAE+sD18Js9t3q14gdrgFtpTQgaPZHhFl9ihX3QCoM76FqRJGQzHF
rr5PeLrU7vdHFR74usITQEq4rGSZF/RZxPfwUxlIBtta+lFmvNuyObBMQOfyCxSEwuA9Ee5lK6Bz
6OigzsFGHtstBefrbnd99BRqAgO7Fd/f+N2+lwLaB7ONnbZA3KcJd1oUNDBkXSR4IFj8Zufj8A/x
KLcmMhsBpcvXWehCoLHd23K9Wrn8xsIeyoFNZ3ZCM6DnF+1lvXrvLAVTh5PnyFjDU6kGh6F60TRy
heLl1S0/8sWodXybDvX2c8MoUtLYKOgCtHZOub1phpHTMGLTfvuiKfff8JxbZJosbk4RE1ksWFgn
Uh8fsiNSP6kK66stfg+ULCLi0yk9JKMr34MQz2w6Jz+haosPsyzBe4kDZpghgakUguBX2Fy29P4d
6pWa7W/iG1H+cQxNEl+5KYQ9lepOkh1ZMdAR5uDsL75I0XaqGW/e/OpQVD6h1+g6gJBkJSc43wET
j7b6OtzPSugcQeXI+1afJVAshJvMCKJqnzMjojP4x+wXsQssYX1LlCGFsQJ9jhDo/9UOvRybQVXK
lgmJHBoyoigIz12DqAyDjKhud70kexVlQhFuG4H29m1JH+I7JdiM59tYFIE/1v4cl56YpgMvn19A
qgRmtJifWUBuc97M5n/V46XDnG0058EJEYmHHTywdP0jBVnP2+Z0j1f7JifHCPxlhLpyj516Vqcn
EMGOhd+S7/RjW80PLFf1Hni7LHBwQtIlcVcK7pdzAn7ockmOB59J4YEXC6qHrpeD8xpxoZaB+DfR
n4bsu/wIkr6shBIQOamczcSRv1WUaBcu+0y3fiZmvJm2j3xBLO+mubekyW2me5I7tV2P9ARel2f/
CA8xMjlZM3NcQkgeyngoeSIspGtJvv8eIYImHeqItw7fvSNLI2sNzWUs4inAE3AbeykwYfwHWYjn
HPuamRfOxCKNFZxriY+UVDADXfZi9m/kJFHM9OGIS5CCN8sWVMva1ecY76O/5+C5HBnTSQX6Ct/G
p8lB4EPexuKYiFvFysxcJpL14MF5ikWcMZdgmf4UKL0kyemMbSk34I1h6Ry+yIdp4UkkDctcEaLD
5qc3FVP/zzMFUP6xvQye6Y4mwo8r27YYKUcl54W7toyEaxLWrPBXLWe+g0ZwKFDj9Ly3clMTFK3J
xiTdbnqIDMr6UP4G13mErGK9AMn6x4yyeQh2sQ1VbqHzDcLZIPdztqK2qCs1bDZKuaHECGImnkeX
ErFC7prIbEpc3JHOW+qkCGkYRIN0lw+/4V0B8mmL7Hm3J5deIudUHQUc7w51lOfv43ZXEwNeBIPu
0sbI3JCwLVgqDmxoorkIs8gP3KK9Q+K4NdLjNLRROJyO6rnJ3W4DeRQaYPurqA6iFqs3kBACpmY2
Opyty3KZjcnu14Qqev145mbESzpXzNLwveowc2I/RugrJEHfNlBpA5Mscqxw2EJ6s7ljUXclALq3
hs4+bJ4PpGV+8WH1MuoQLpm/AzoGhoHPDHSQje6g3qSVUYDjy9TXdu7KWg+H2XFYeJOKEMf7YF+7
AblJMG2qU1KDmzsceIV3515PNY9TLfIlzvkwKnYeIJEQ/WHmxJvOyYDRar5RnFkIARdY4wbcgGN0
tz4c1edonXWsfQXuF/Apotk9F+YC82Wp1kIy5SthN9n78CGulRO4vLMhbysU1tykKBg9I19WRA/K
0NC0WTBFIsXKmqSib4TH+XAnHFJcVklxLaiz8xs2lOMs7ZZvyTtMCxWG2iwO374yvzQJTiq+QX77
5srDPiCBQBbbLUQ/G5qaQQ6ENot43udIlHd9ZVh+mTjlb9dPotH8wshkzsu53Too206L7i2z2v84
rpILqBzCV1lY8WOu5XZG/F+zmz3SAy97tdUe4Uy30dCAUFX7tSd9+9C7bXVgy9FUM+IttFCBTcmu
GyZcEq4bvU5tdSpMd+B/6FLsI1OOyI5xlwsf1NQVFOyPg4lnp4jWnvzyXzast2IolzZIzvpye+l3
V841ngfIkUVXKIQDq9u1Uja9fkQTH/tgiSoW68GWe332tYIw6EpXdlVHAgPLWzo46aqwtB8LaJnx
KfOqk1gFiNZlSgMp64AckhaIdheiKqf/QTQUxHGu0SACQTbA1zZbUttHirjp7x8TtZyM651l0seb
7LfJV805T+tb5fkI+ZW0Q43mMfHVqA==
`protect end_protected
