`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
QlJpMRsgk+Aw41cWq0t9Fy5yP3BA30M/ZFFgd1POCfWvsyGQlzhETRw3YcdGMLPZ2LnKkojc57MR
wIimRK2VlnBfrdeaqEY4UrRfW0PZSbmur75Nu1z0RJrIfHZ8W6LlEA4jcOtCbJEVUt0KKhSIAVw/
o8TYCKD3kvDm5gSJccrm7hMWh0GLKohSEs7zcXc9SnwGse9YFB7B68XTMsdNOdrNZFVylOqigNn2
2BaKKSvhKau/631d1c/pbm+WxakauNCzWIqCRp5nj8CIPjVcNSW2m8FHSpbDUHfCVZ4pOdtop/Bw
hzejdaZo/C+qPj8Y9Wp10t6m3dZdWDjF47X0CQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="RxotkYIscEdJrn8YxufhlJhyjJdLedMy6rPEB2S7Qqo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15712)
`protect data_block
JizMoOCLDGwzje2s8hEkfqEN3walWRkIrzZqMs/acpjmrnGnZct56hkA3pxWkkCxKcvNm4VKm60+
BrKJrIu+/VELg5ptSDrkq1Pphaz3sswBji9eNIjFTNndcxQRlAwRUUFlkD+5eweHcFq6MikV1HLU
M+/lUcCIV0XNtdJt2XgRp0x6CN8sYruBx+akf8zb1kaBIJBAylt7B1UPxPrx7qxGqwS4Kl8aWk8x
MYaYXBcu/ziuJGeAP6R+fDnd+ucN6G0RGnV/xkIOFX9O6uSB/OuSSf+Ld5sdwYGVSUd4twjZMzVz
MMiKK7ibg54g1XaYXnXBZ/KgafrCJt69crjvFJtb1qt/e96U+pGh0HDTLJ0NxcjoJCC/3Awdvl+0
yUGMWoVjMQvfgSvPQtxCRfBYuEVJZCmuPr0cmrHUONLNczvSd6/1w0IbTYG7iHhbv2/fIv6wTA46
2s1Dg8k3+mXgGXTGA2SSACFDqvKHVNl+fKRotUgQkHb0lWTo05vcOoBD7VNX0Og0WJJB+0Gqxzf2
iJBdopgNkBXLuLv+mNsgi0N/0N9OBmpVRVNhK88WmdOnY19T0l+OHY/1dTZzom8fzpstkdBuUUZw
FmQBAxEA3CXL/BQXKXW0e2yTJg8sCYG+k1IrVBsgX7J8Nsj21QnQ+2jHwHeGUok+I9h7ZB4pcpoV
LadhLPlAUVXXkdz/vFIQSJ9FxfIeRgvRAoFKcITN42GJfpYjQaGi2TVYe08LDGqeEUk76mtFyM4Y
Np2SppvloS3QhRI3LBpaMbngUrgJKKroVKLG4i5IzMLo4KpO+sdMzC1ZkhY6O0+tqwqf0/diE3Tl
xK4AKZQaMuqq9vdVz6IbtrLe+TFQd9mHDe/hbXAbmq3ARTdaxjgPdlUJ5/MJWhz1ngdySBzH0gvT
49Q65/f7yFpDrLUaWJ4BKCEx055oDxhqWR4j8MGOZ+1umuvUX710Q0IIeLfwPYTmOWrz+fpb/Wzy
fba6/IDmCIQ7cOSchSF4D1NU8lopvvKBRYq3XCpEkvN2Jm9FIK/VGSLnmH1cPFH7Aq4rLWvVwggX
yVZIpUO2Jp2KtAY+KUcTaArrZ31ih5hngNfAIcMjvbXajaWR7Q7w/0fI75ve5ExIWePqCVFhqJle
8jpgd+tHTEmA3EK6H1+UVkJPJ5QXfbsCWPkG2dNEEOPDkh+3/tW0vs+qh10YShXh+6MW5cyF4cGz
LmWeCCqlz5qs3ICBCt44t1xEIS0fneZmRzTd4Kptz3JhMlVwieOf2liCmGaJgNSlpZzJN0H7LZgT
HaJwED2DRKULMO/L7Y+rsW+GIEyoh3js6uituJK56fHOd0DPgoT+y9kiPHWbdPkj1rcWk+L/aUKV
4wYqo93PiVJrQ3c6Fx6e+QqvZ7S7JPqo0bvB+Ofw5EEvTI3v8LB3HdWzvfNTaMQ5WfQOXuPp6mMa
0i0+HGxwxBUhzNazqe4M7aJ0OJgPAxvfhwUuRTlSgFNu4aXtrpMF9xv0hrIWmbL0B16N/GRunHAu
5xz5C9NjobH1Toeg8wabdXpJws9QhAo6r56TC7e3lnJQVKjYONgP9hqd6i7TXjS2sTSRQ9llr04Y
3fIafJhElq7yKg77e3yaCAmuz4opFV+JG6G03dbjSIL+Os+nKFysE5mpWowKBcXij/p/U4nLvnWW
y5YiW3mDmtX6JfTqLZWIsSZGEOcJ+WZwbxRvna/nQuHZLtRqwOugwo0OV8kSPKjGrPpO31HjDIgr
md21njOEGocWUWriZLJzoTcbg+TFH7veKgUV/ForL8wjXCl0FEf+W71qD2ofQ71r3q8QAl0EABq9
Zjciqhs0k/rfQhCrCdrb3X+DbCl2DE15+BD9AQsCKzH6LCJ4tNbvAtqhZ9y0jPp8XuK6nkb95Cd9
+SbJlR1AmDAqDklkfp5XXCNBukpvkgXwfrUMfmgcxKhutzUcS2yfiti0zZ1zTTjq/H1clAEITzC4
KKZGT0YFUNFU9z6mjKTWitAMit0/ZjAh6TJn4lmnS6R1xH343vIeDFWgL1tWiQJGpQ/+4PM7ITYZ
r+Z8cm0oW3ODx7Qvd6U16sdUJUrwyHgHswEvTxuThVOLQt2e8gNeHr/fVrzf4lbSz3ah4dl2MWiI
jYD0rl03kLVTD4Hlkybs1sDyj/1ktc52ycgTmpoFdB+G4lKSu0ezhAmud6S83rds6XGlKpK69ags
18g+pN46IEOn7pqWE+xifPQRmgm34KHxc92DEzPFzBmDtJk0zLLa+V2fb7Bkv1/t3rq6T0iWr1yh
Pm7AiPOeiN2F9+bqia1KCMGiMkfyoIDO7XM0dQGmxcWL2fErrsLS0c36itQIZk2cOm4PC+uHk9zj
z11c45AMB/khe7zDjxsA3tBozFkQcXNEJzjE8cyjVRF+7ftz4x2+jIt36aka8kV+ubthoo27bUEx
ug6IQj9ZgIkc8kv982mwmJLBQZ2Wts1Zqh3/reOm/MndqZOeKldBX2x0jTkUBey2rFOFoE7YqV4m
TyZAj14wqSIJFXRD5jjRYGNCoq6Uck8PPAbNZf726CEGpP5sFhzgdE9/y64gmJnJtwKAy4lYd/G1
FmFuneXzSU9H3nYvEWuCmBOOUu/pL1smcMKKFob387LIcaB7wyqi6kF7CfQUD7vkz5MBElXAFAmE
mHMjagYUyHGlH7iSVNf9+LB3wzUpDzk48zpdllgx+z1t7oqYHaRKEsa6D7zJtvk1+YtXBQUu/6c2
8bif4DgeNFz/EXaG/iK4ifT3npkzU1ofOaH5v2M1rhzqNFVEKZ+CzNJR1QqEFvWSCemlXKROP6uf
yqW8NRVq0DSLVRuDXZqilomhYLllpD8asPRU0XT3L4GuBd6znzA9zhaErAisZe5dSV2d+OJurdfo
VYb5OJDNH74H6SEi4Vga4QFvEhZWpRfzNAQn524N6rvx2o2URcOrJr0h6Ay/01ZWfU4nwyGdA71o
Log6bKdWSWoJRffrAA10lRrekpCZgWIcoYxEJQJE9Z6ZXpy76BLHXbFq8L1/pNnx0XMrJKcDBg+v
RaOVNS8xmIb9Tx3fYh9pFVo8nycydlgLu3d4n5oy61RQTf7MGVAIlMs7t4H+E/5M3MSPw3pW0tWS
d2KE+uV3D7h874VlJ/lgCTs6lvIUUQR8v07BFVECiVaqJ5fMckfV6b6DqkhQF+HNbuay7SQ+ANqw
rP0nzCPDkQkJYX9xwlB7s86Us3qS4Cw8hVXWlE8DvSX++Pz20cthUA1Bnnjkw74IMgmiV6bFoKtL
Y4fDERspfV/WsAURHbCgGdnXV2VUwrK951gKYa7y0kdkkAw4HvmqyTSm/FrdupoHz8agMLTkmCXV
bdytoyvP1xde07agyzjiq7jHt0WaJi1kUkERUgYxXlAMduqEX7xIKU4uUxk/k6eAmzA/iiL/MZle
LiRH4ZpGm6NadXaUksyHU4q2UYa8TugDfYRdzHpQholSQE5HEg4uq9J8nlvRvO5cnRKYw6WhiGhp
dGmynInwdkhKYtyQi9qWv0U3XlLcGn38wzrX413oI2lLGkJtBSgfR+OSl+Usu1yLW33LNgA378qB
JzF8ou6mAuvIc6f0m8j/R6+QXJyuL1WVR7Do4XuM4snGQSAt/gPF0cDcaQBtqu/dnZgSIxWyHVFI
OdijbHmG7EoNQLKMVIUDruscBdJiWfZUxUBqGv9RLFVd6L/hzjksuU0ySRHa7wOPwimWs9OJT239
fR4RbxtBhkzcVX6DPlJHhLpQWuHoxUzhgxz1eAro+xd0nIjWYSa9d3ImCJvqP59ICIYMTIwZ1ITb
ykDC9Q8RPbNk28b30tFVfJQovKMrnpebgE8yvtmyvLv79WzsBUI8UCrw3K/prgb+NJoWPgoCLvvw
EBIdV/5d72wEZaImTVSBC5fct1FNyzsS06KntAxopwVU2d13hsO1Rag4swsSY5x/DrTuoATQi+Em
Ur7bmf5txNI7d2aJknrdZr9bTN+K5CD0FilVW1ElaueV7/Ds+B1PfxJQz9ztI1XxlOFiTpmevbgf
tD/xTQukrDH59So6/VzgVltpfyYzLGYsMfbSUR4RD68iA0krPK4g/Bfe9f74xRLNYor+9a2r/V6M
DJ/3iSRsqZOXwgIMn9ZNu/PEmg9myVw6p9992KOCcxMv1veSKG5adQVnX2QKKL0i6Qek2xM/MEGI
2TCnXiWOjObc0UND3/IfsbtKoGGAzHuznrzDtMP9OPmegqhgtHq2aetvAg3uuo9BOA1EEO0d8xB7
srzH/IKJQH+D8kQSdA/kPj+87ulVawgCdjnKWwsplzJA0LnwXub4C6DoLw3TskndfQd0lOBATZY1
CxyCqyq1G4pJzWYC6Bsh+pZyK/d4OeU93I1bEFk9iLpiUxNGdFXSi7KNgT7PVMXBcnkrkV1Gx5MB
5y6h3SoGY/Vzb5Ic7YWvEJuPSgeGGAyxCnqIIwf/gHWa07HBYLBucsv7RVKhY0fEIPCl1V7tEyt/
rkdm3GvxVR6enoXbyp0JjyeiCt9BbZWpAKrC8ng7dcBD9LuCGYNHqFywoo0SuvRvfKPkXKc5IvmO
MQI08+NGTeRiJsDwFdt0OF87AZJwlRz7CAokCUP1GKoYXRLZe6ya1ei8WIwNFjInqRbvd0YYqu9m
WLOS+b3ujlraW3zZ9HhG9xk4DIcvZPbhg4H4bGSkJeVFR0nznpCjzwP4j5Hl31WyOsSewQkabJyJ
cOPEQzv8bPhXJUpX0R2rn1Y3i+HEBuMphsb2yrtSHku4JNMPiotWlEQoPJavy/0yZ0gcpnhC5Xth
ivjgTbl8tTqzyp1tA/6GrDYgLH0mu/FNFgadHZKgXqHQZN/z4Oe4JG2YK9nOhwNHHK14JfX+s33U
E38sAxAsiP7jytQPoe12WFga62M9y76Vlto25GFd0kQQkGZ1gdSI3nZmxjyGNeZ2CrRSgY3ivLe+
trFtnk8E8+gEZ9WDN+2en3h+koalt3nFcgCbaK+X13aA9BN0dVUTYx18rptL53NnbUwaUjSaEWak
xxsruxUK42IYNnoTJD4iIBszUTR0zZQZJIYoTmS17tR83EWMsSGb9ejiy6Rrpx5goT3VUf25gmss
P6GADfXJ4wc94NXdbFzjruhee48dtnWxppIdq8hxMiIwNEb5mtTfiB3B9l1N6dqlBzz04hrk+XU9
BnF/rBh29ZuB17X3vI5mCVk39RYE9NwT/vb0gsEZjwmOzI+EgISNS/nIInv6rxklvpzY6fWiuY6M
xKb3rHwJiVheb+4n/3CucJnuBtUcD5P6bShZylVo9TrfC0+bkrzqM0X7tlSb+gJyqGq2rCYV7qPy
/sFZpM/mKoRWVdiLtH5lCIFrk71j6C0TK5BSuPl7fJggugDOinuqZlZFzQKpdRJ1XDRkl1wiK81K
J5Gx6pEsMfc9HdO+zoPw0jCb5gAXCk0oTSeLxdDNoVHwGecRrELxtjU60syShpR81IMdEaRU/iHJ
CXCyPR12RqdbJ2aonraEUeCxZBfhdrNztbG6F0brcrgGEP8uunYx8bWjm4JfGawM4Qqs8IS0Ll7t
RS4AIpP5l8R1XTZr/or9wPqH4vOF4gfmxxEBSzwsv9oOx/EjxhKOFnP9bVpIBf6RzcEaAQsFvPwC
gZHO/+zRDOtHEzRZiNXMGHbcX5plbf8hEjlnWYYtRXsT0HXJRbPA1Fbj5vo9JnMlYO4NQ5BB7ZhF
fPxqMm0T1gYs1FCcZ6kNNVocS7OBMa9iR+NoSMCRemYqI1egupxmgGTtV+dlSFgvps0LzZl73CZx
1O8TgCzAvabMU93ZWizt5qcxCq1RK0uB+orrq0E55NV01pJuTo3A7QZP30BUc7U6wkuxS3D+u8/Z
iDk8YinvD98roQYrN1TkvVRC0OyNaAqH4f7a2NHpMTWH2pRZsuGRn2oGTo/8F9sYutWfE78jfxI8
oydKXTR53c9yWXRtWl2DiMyrIBiU+Vbj215VwE2XMnmWl2k/xiMExP1NmX+2R+MJBdN3QlYQSwRX
0rhGohFas+z/AeeQZYCQQkFR/2MBN2LfcKMoX4RVq2pSg8RLf1b5c/jfozXxJIU5dJ0yu1r55oJC
txN4pIsb4+/eY1fchmiL2ZG73ois3y7ejzoI7ZIb/7HlVe9z87AeP8RAbfeb4Gnnu2vOxAxmnJJS
km7ttpv2lVBlWa+HvEWyj2+JANAo64ThdQaKFmeLTwe9gd9eXHqLgyxzSt78m1TD/GbndNYTAhP5
tZQ4eQkmqiaZLD1SkmGW4APnhRPYhOHSGUP1D/JUqaJ4+lNxvQROnIUndds34xKGis1Q1XkC+2A2
NOFYlOJoB6rW3I1EJFpGkxsqYuKbgQ37MobIiMXs1JryzJVdS51pFiJfB5GKZnR8I42TE5Gxh1MT
y2xfmT3LpwUj2gCHqNqZKEqoxlLwp9qK+LYNuSMFKDlFESjxvGzBluNyusETFGtxZXPSVcyfLjYZ
lG8tdkQ7VyTW31dRduIFirs68S7S9rdP+lxq8upi7fxxaOsKozJhdAkCqdewX91iQmNoCzS2D56c
tw48oWfTIrsVmVK+FM9CMCqGCvpO1aXjacugMd0GNZGTV1RFzd1Um3q1gSE0/5i+PPVlD8djPvQM
2IspWouWfr7OEnksIjv+4NPJy7ar5F/oj6t+OuZ4NHJhP09TGXyHr56Bw1wfeEpYW1fJpr8PBkXj
oEZ7Ygni90tbB22y61YAivlkFBMxN2wT9Hh4UCi9EygvAclSPvgqGfIfNPY1sqm/dnoivl1Qp/4F
UGVJuUh2UOFHPLABBlQa3vpUsVBRO96YcL2L6NzJMfWrawqiVAotBxrF30xB4Gf/tlMMt3HNbx9F
TpLvg5TH+pERyq/KIjmwk0kJPTSaEVlmCrKKHSHB1FG73fCwekyoeZaVv6tMO1QyD6A/+9NDk0Ju
CbHrF7fd6wDajHfjp9AnsSEoNrOoB5fPTAXWLMNoQ1kGZJSfzLUxmDplwHvIEdSFYHcuJC5LMtOw
Ewzao/wJEzA1bSu72FKLMLDJy7YdnATINKozqKUZYIBT3knvmskJlExwT6PG9pAJc+QgCf5f/1W2
0fTcgItuXVpDPnnRXrhnJlyt89f9zXjiA6WhrJ0yxrTYMhi1/nATA4Gmg0l8uhWI+7g5MAArxys3
u4oZR3ZHM/JzJ+8JIshqH0bCqEfCgbeLaMoX0gU3l2AYC5FllN9xlK3Pdb3nvpwjqbtbK1QLmLHq
d+7p5TzezW8xNdLnwFhiuBb1N3q71y2VRF8O6bg6BUokf2Teraa5D+t6QZ0z2HOoX6dzHTOlKQwM
AShVtFJJ3mjJ6Vh5fhCzGjutrXrmRo7CXCDwzZX3mGkRcq8tgKTNTvfodQOEel0Ux0i1wg88WvXd
9ziBXHEgQdLygy3/s/yUJIjc0uY6K/mH9r0EFvD9SttYowK75DvtXBPw3yg/edFJUSXKdEFmOdYV
t04OUVa3ppfCzPuCzLZ0mhf7xvIXSPolGwQAgU5uZYpLyskDeKuKuCLNPsM1nSEjWgDzqId5znvN
Ut8A5m+xkMzwMrUGsfIi80mCT5Uytlj33FV7ON+d+epGXjyCIWkFbTlCex9HKzAzoUcxlRNpjA1M
mwxjtC8VPXqRjDL5YeD2unDgcyG92HQlt/d9jxCLrXk4TFmpNKL2M/dmjM75KBtMUnpvPf1ixirx
VjfNBac2v7DrLZZsiDWH2tCvfIo1R6IjWVXdr6R1oL/qjknIIv28TGCG72RkRyxqwcILx6nukj/3
eP7cvvQWL/3NMU5rhGAj0M2/IJnYzVZh8fGZCDoSi2dJp+m8UIJGefoGql3cpMYbbca92N1u9RvN
pila1QiBfGxqdwI1zFq2sae2EEwfk97Ddqo1ccjmg/xeWVXn9NhYJiLsuBpvvIMBOofmsoorviNb
piTs4eM/M+a+W0GzzwBAB/cq3J9bHCmxWy8r1sSUpqdyF4w3F6RjJU245PEOrK9Ag430P/+TdV/5
dVSe3lnupe1FnBFZ/63Vvo5pdMrooa6BqzQazAJqqg8mdZZPItMIGRNqeWv6DYckwsQVDv2xy7su
ttgI9Bw3msywxyRHr6eHj774GG29I8SaPQj5lbChL+BtEHIaNXUTRGRQq7hhbDwg8CiHGYBz8BiJ
OgtDh5BAxdVgo40hXeB5MUAmcRRomJicQR+ial2LDIoeZvCFgJ3HfMIeNhBPBIyGLpxSG6ffHSY+
o9k4sN844Q23mFQHdNAlB+N1TkM5Q7DIQFev9mDNCBS+oHQ/vGMCTh19RusnKN5YGrt7e0tLE3q+
HqRGMQKcKQlhOIwzsTDquAK9yM95d23ttbyUBywIMmhVTRqo7GwPCMawoN7JpG/pUd+EY6idIZ5R
MKU4ypckDyL4Z+bYu0NPwKV5dWoDf46Z0TXRFUTCtkGYYXtKEoekf7m6yuuRN6jcluw519yiEbPj
88yqdje1/cxvDxl7vkhH3s07GAsZYVKGmLXCVl3VDD8R6jvgPnb/S+6xanXscvXWNcu4Vg9+Eb71
VsXMIWde0OZJJIYVYa+/BGD1PIo5oDB/V+1i8hRjm8QQFcd99eCN++qTpL53K5WH5EIsUw78/Kmi
wQ75aSVjplvshoN/9hwy8FoP7uIJBnwHklCGWgpYlYUbWxYeE3Q8bIn/FethpBc1OT2SrlS0+6J1
sSghUMRcsvRulPHYqB0v89bGRntSDqr9Ow9fip6jROiztiyJojzRuHBGgQ9lpVg9rLyV4T/yVY/Q
qdlsa/A+27HS095lBe/RJe23Nsy3NTTeRKOGZa4FXCOrFgG+XmePX7n9OJpALXaNRlZfkMax0xnE
4aZhHngfP6Vt1cJtbI4/HKo2kRoVxcYgkjtxma7NG6igG/0UXhg56xLLnAqOyDjWns+RrflI9YM/
nafl0dVpaus8yglCkFPCq+Ah1n519mvrjsxrzkmBiARw91mae7Q0N1cwgFujMu07njfE5blmzy1t
iPxPVCVulb0pv+vtycyi62PP3lmNrrwJlCGUXT/ZJs9msiHbejEUD2n0m+jQ1x/cUrKAWs+yI3eY
iD37zyAU/MUlGtXN41a0mhW9P11WVEch4P/A2jImCPfbufVpAt81vQIVCcTqc35PcTPRq7S5PIH5
r7+ZcFhhtix+3kQ/Dqk8l6aYw/jbG2bdtCIiXGK1zjd+h3Zd1yfyIb/MPqytxOAOUbX4wwkXbHRR
u9bbKfz4jh52GKdIheEfiQcKKp4RU3Ygx6Dxi4ulZ4QHN6STrbiDmKHk4CKUqL0v+l6GZPRkdtZm
DITsgELhT+FoBdg1ySkAB0JahV/7EhtOrB2yvhdRJYNQwh0CImOoiZVxk9m34hvqByXKTLau2k8M
Q3zxLrSGlVXvku8atMhn9C5484T+64R9QlEaQDlMJQbfwZcPX0/YgylK9ib+bEjzeaedc0OGRFC6
6eqxn82SfQ6hndR2AofYoVXiPd6LQghweTMC3EGCxRYOkZgb03HnkDY97PTLjc/7PaF87Fprx48C
ies/ZQAngTpU/xX/H2mSMH3anfYnzFderfNv0sprJdWIyTBUlRRgmS5hJ296jWpd8lfTkJrmw/vv
dga8aeUZxuL9vYrB+x2rfbQ6qPV78MVJvkjYJB9v2SicZYCt1t6jXnDpZSH6cm7zOjfiBKXilyXx
xgcIlmSi2qopqbj452ere2nVp05yi/C4A09JQ1axaewJ4qUTXcuhB7edtPprR7i4KfogqmMC+XqB
vaJwXE4ek28wdPCLgIGKkGm/VAgUmQ9okP6kCi/OP5Q2nNuvAiKdSNPP6/mF0s3OVOLrFWLlFXu5
aMcR7f6fWqJnP54PR8OhRLhpdLPw+O7XfDisX3S/J09nnEGNiWLj7VHiQ35ztIEw3kUVKbsJ4L8O
aSIA1ntGIf+PlPBVeB5zKHOE0LHLIyLD0opqR7GKD56bsbOHbUp+GO/aW3suEFRpEAVMLjw0xeR0
nQpVbae4bHQzU3WSPLeLt3n3JRPpLz0BI2IC+IO7IBvkYgSbr74lHTWQSXojbN+I7C3p5QNqr1Mt
z/dwed/IRZdclYMpJ2cRDTRHEpgVuImrekYIi6sPgvfITOGt4KmhlYUV6jhDdKtNHc96u3zvUXrh
iiGyeyOnQuZGuW04dwC941k80lmXM0Xl3sXajXX2lbz5oGJLtWCKcCOit3AQ5nOtzLL+O+Lq91Uy
dONrnCeUGSycl975pIi6BmWBExGPZDfFM2WUoNcV4li8JtD+7Q3h10KDdusAf+PxIpz44ZuHwcxM
NhT9qb6ZULJ3cgg0GFp6g0eAbT9Kzu3pH620WN1wkwhbwhck3UtpaxnBWynL9T7KRK3Ef3SQiA+Z
GvzoRJecpTmacEjgFmfDywh5pdwXRKj10rUpF4HOhQDTgMduyFqaN4qCZXXD21ZLW6W4aEMI0Gk8
CaYH9/q1hAjP9gQcqZRwa9Z5hPzyOCtUtLErBfDYYFHR4sGf6l9iJUHI6WNg4wo3LayJv+Lh04nt
Xp+wRaMD84rtldaYqDqiJZ10PdwDPoPxgBSBrmBA05bADhb+5NshzdHZq2+JeFinHcN/ysiufXsy
IKBGFeb5OKLkgIDoTig/W0nxl0xYjiFSVsFtaWpIliY4MxeKwP8Qw+VBA8NUxR/H10LeBSpP3Gxv
YJPl8ghctvOLIgINVlCXJiHQImaloHKMVLuzNJLAwpOeRW7he+2wDmD+HilSeh8VvY+lwrpGoVTH
kZ1zc/iRCdynvc6PnbWn1A5rKZDgN9TMvO1KLKXTgUqhxnejC6BWHKKg5eeAmmBqd2fBnkPMab6+
9EXFO9vVSOuakN7wk4fmorGE+g/UrvTslrvDTvfIXvXGQdXS76HkMaVu9Tp5ZEqwTRFTJvjWtaud
oJBWzKBgAwMFKr9ZszX7wFJDt/neMuAx2/JxMI2M8IjfTo7SSiDsNURWCYpI4drHX5KLzNI3XFUG
VOYC/RUuEqm4Dh/2LUurvwGOp8gSGcdr4DaMafKHd5RdSOC9AjNelUIMYkfPIb3zWLox/pPaLzDT
Tw6XNRURFuYyKnX8n8hm0eXXbQV8BB/PRCY/GuTfPHH0+EcvXUXcck5B8ZUGJt07onBH2HT10Z8u
UtttD/8UNK04AZl5OG4pGuWXmWAiMqQo0CzLoo4fEzaCmNT1sYIWNhDn7hdUfGfFq+LEaZ4J5IhN
JwfdrBTmJoXjHuW38DvfGPnYGKhrxhokH6F1dTO1BNZxUFCPtEKdL0zMYN5D3aiGQABFgWJR4EGs
8VB0as8JWo3E9N1GJ3nCGAB7GVS1S2eUQ+G3U3KTmKpDOY3F4M5N/iVJPce7FPbchaq+KWiUKU8m
mfxHedVcejx6pebvLbT/b6OTt/EwgVt0NNvVN6zW3eg2ICdAKYuogR4AL6SD8Jv7s1NG3uG0FKZB
Y6STht9B6/DENFJXsP+6Ae5jxk91Fh3OocurfqrK+IV3Ev6ST8THZ22kWkFd3vlQlnRVvKGbrZkm
dOcBqXSQeT7U6SBN10k0pyjN9awd78BLWpbjMwVTlPsKz+vGbKMIVz8WGy/gu0LRalj7faqgMQ9P
mKDhALktVf5pPodsy5s49YQaJkXUwpR//y2d5VkUnsmaXtQ2p+zadXgIG/KCjICo81etn4nqmiU8
WNunJ4JK27Cqt/4PJt/6KmkgZYgVViN+1goMuZIC5sKfx3POlmAoSjQbgFy4wLc0pb//61xvfWUu
Sz+KF4aWfw+8yTncfxEHdogDb4YoLqNDMTBMOTGtSZV2kkCqjkX3Na1dYPBbzjTqC7jlWil68YND
0vgP7rZ4RGOL0gM+8WWug4YxhnI4WSsZ1ju0afQuUHYoLL5xC7hgP576EcBarqRvs7LNFG+GxE0i
3BfB1vYN9fCsmiHPqGDrMZ7VYwKEQnmKZX8gRy3LkvWVrnupf29VkQjlita0u5asKPlzwHJOWJEv
tA/tIfoNYBtTC6VL7dbpljyuHovMmhPdlWdg9XBABj9cfQVJMQzlHhmM3xobijE5Q4kpjqKjMaRa
fVflRoSA/SXqaFRej/MnryDzTG3dnx9ZGnpQvXNP2omB8Q/1AAtwrUfuMHo4oezebnE70nC8EYqu
MniOtEqZuaq6SheHSNA9QtVjSsBv5tfI8auY1ubraaXxe4QiyUulj48+teuIcDVKVGL5BslomAPa
N1qeaQvQgQkKzUXAv3sXPL/+ojG6aMx4Dy6DnjZ5JhpM+7U0o//CaiPhCXzhqzGpNewlJQ7cUbJK
T5rUJFC+lPzPWuR01dN+NQ6NWKnT9XJJKwudXkZyceDft/y8rE44tjCkXTRtz+/Vc4iiHcrQliCL
tpJr9xWSuttRTODi0xRfF6it91pZsNG5whKjom7TGSPbxxEExpjTU3oL6HWhhlW/laIGEjwVFU6P
MIlWZ2r5SrvW3TwbsZwNN/TBTxznxzBiarITORAAVj7ANlAo4S8X/grQNX3CHhHpEvjGHISIeGNJ
bZW9R/01MfErkOzDpWkecT+19vao9sop/ZCk6XwXVeZrUJcmpMKY4/lXGXCit/sRpMs6aFL0azRv
In4hzQ0YBb0lck0cgvEaA0mFCKdNkdjhMKGxvppt3qUCgxQayNlwZetPjyvYt9Bf3A8l6gIg1b1F
Z56iD1jpuj4od+qOQ1a8I5mWjw3ZzW/oiORZU/EdAvA2/T0Ej6DPTKMUebS48K0Jz80Y3A/5LhK3
Nr4OWF5EQJQDHIoXhwQqxQr5wyaaiS2A6LOj7JM1ur2cWCLzZIQkP4h69LstDsW0RrM8LW2KG/cZ
jYBchVv67wNalV6EpgGivp8yJ3FEIg6gI2IdSUk+kjqs69Fqvsdh5bIJA30dYsfUg7BCgy8m70i5
gHIioH3RiaPLJQ3OwJ020vwBMvmgrt8+s2WjyCNOSB858R7wEFYkU7Jlq++k/Zo1+xAT/wIG5Imw
zEIU0KFMbL3mexDn13fxdiu1DRjN2/u1cKNnmmUOtFmweOWw6f2XCtMMlRTPD/QBFh0ox05XEAmn
boLscN5AAelcmJG/2QD5Q1xp+aW8ONEKGC6nS3Sup5RgUYaM7jkXX+0dWfQGEQAX1h3wAcO4+5Jb
GQgluu1SuVGB04d2KWv+11jiab8mx/WpsRyYPhMWVKgZAxySw0zHvKrya54zRFTBVRK7ZP0258sw
5ENodfS0muHoqy0dOLQmvI5qptQEfhlAjzgEEPe+D58EmKyTmdmaVndh+/al7ZS9LIFVcg7PxDrU
jF+vK4tuJmU2M0iWArtZsvOr/Jno6nJSBS+MydU2Cq2o+DSHkFp1kDKdZjINKbYR/2+e4wjJ8/bA
FTii1mZaA/EunsoymemXaQ9r0aHh/m8dMWNsGAiKQ89HY2+UUC+C83OA60olhhoHJictA4e1MExv
okIjSbRW08uEWKGhMVOrnf0Bossq/8xm9zBCM38tZfzr/YcOIw0n5eFnEyUWKcABB1rJptXpe8v1
Bs8g7FdUNfo7AB2WjeNrn5QwlMcguji2ImWAn7kx3tHykm1dj68yLSrhQ6cqZrMw53Kylk1K4AAq
u5VutNA2+ASkNOKarhrZmZQFAmOtEAUbvOP9O3g2VGfn9e2ac4ux+lSN80qQVhaFaNOkbdgPOgfb
yVULOELWEXzAvUPHHxl4Vksa6pEjlRlFoYrdCSJ+ez+T3zccpX8zXo3P2ZdsYstaWmX+oPtYKz4D
VDwv1GH11tTP2NoAPOE2UR0NXN+X9hv53N3wA2CjqRS7znypaENMNvmbss7WUQG2sLc6dy7wMjam
0CXTxWvYYhPpzcVN1iMRifvcVKU9N+m4b0zibNKdlYXI2tsQMbtGy04/fDYEGFElYFvoOs4JJGsg
HcXpRh9t8gbee+iI7IjLn98v5LCryocsRwUGze5A9ikyKmQnFK287+6f5kff8ffM29d3gNTKTRpE
ubcXOhcHANznbbQ/0Ug6Yte4nCH7Gm8VyhCj2KWEhm5KBEK8baCwzSZ7tlB55R75ZjmuXkZA+etd
Fhjf4gYNChicHJXW74nQCQri40vEsqNN6EzszpI+MW9ZymepuyULuXo3PIVbNs0dtQq0BsUFBakZ
uUK0T0Cw4JJEsp3PoZ36r7msnK0IxfkQbDa6xS42X2/dJRnwRCw+zs4292+hQBUGN6rgYWvSmYMf
DgWJDwAehCdKfOT7t/nKsN6qyDYpqiHZ5qDRP6iexJew1t6grv9619kwavufObmQMWlBy+pE3+jQ
Qk2QYWXv/rpyjtQbyTXozeJueKXh5akDkPJhiY6fEz36zoCW67ZvOza+DA15kAzZ8RaAFI0pYckm
TkvuQH5fz0NkI/uurh+ckh3S9zzj2vXgTYJ+0n+dX+XqBLjz/+fze96Qt6Hc9hU4n2sa4PuPa+6w
uqKexTcKg1DKXe7uBCONyLDgMoZRjZ+w0YE4VDcQGxus6B8MO3L6RXJVgqMSoiNwvlH1WkYo2ftR
1lxtMB48KiTF3xK/SaACm4poFR1tYQn9D+nNebbc0EgFWsvpnp6ZqplYt1j9lvSyflleOivq6dIG
OOlf8hq2FmsxiftX1JJjxM/ehPoLiFhmN9Fxv+FBQZmoCDsKP9Y302so+ZGY0OqnwAuVXRBuAlHi
FhKJPspIBRsD6udkJgL7TOV3GwJ5mAbCVPX25+KN0HYGW2vr68k8dU8ynK6mLOHGyuTcdCziuJ9S
oe22NFLQP5WR4B8kHRcWVJIQ2K+sicnH3Pfu91I4hN1FvuxEenHK9puFzCdJZD/TJhiTzgjKme+V
PxcVXlHQ65V9WR2Sm8ZGmwhtIF4Jc0kJ+NdtZDwAuKheulnknaiCtHjIb86Maxtj5cB2lazStAqc
QV6VV+TbOGal8qpNW1ht5PtrWXR/2KDQCTLGJHYGWWfdaPVPK8Wdgp1d3HHGySgFcthOslYQD96g
K9kzEsk1cFDsc276FlyAHmBLlgt17JkPvfrQ0ebkI1Orgul4wb8lmZsLl6Jv//cXDDxGH7t/Bhs0
f4y4G7JcwOFCjPm8IYKtSg2A5rqgVO3ebNZ/ah79Ex09oyUA+oMJokZBWRcIs5wVPtZe3zgnYgIl
/mtZwmLp2BmUeciNQFzsvGBnGWKtYI5GqTFR06aM36i1DLKAfccKQ5dZtcYDSA4XBYCWBe9YIUeE
HHczIJ44wW4Jm5M3ALbLdgazRxgsg1GzcRO03EcGN/WMLd2LtFZiShJ7SASHk0dCe25KBskG/DCI
ceh4zYknS3TG1LaqgJazIVTTDv0Eb9Fbb0geIyFU7w/S81iPaFh+UOXPyKA7J/OAIPH9x3B8m655
T6cNdl/6TKkwejdOhpk1HlbUBu8/YfaFgu9WyOmkWqqmol+y0r1EDStcVFpeYyJD++YRdoP45D/H
9wAwr+F5r+tqOjJcVwVPSN443urxS5s/SekSfBI+8PFr+zlOhK2xLb/PrrIGSkPXs0yCfO8jv0rl
54XTfiBNUeQxvWPanqGK4Xnn57QczkD9722biShurj1g2Gpe7+CB8K4UsXsFyeXam58dX5g73PMX
oiEVSSfLi2gZa/C4BYlEihNVpOMeLjncuNO6rnileSHr31wn+Bzt3dynRQPRp8yYLx0NX064tA0F
AD0+pl7bkNRmPIXCULzNzeys+K5vzXYBStydux2i+3nKqKiQiDJxq1Oyx79/BWeIHMaFdkXmNJl8
g+7//VtuK41byjRGxN+fUrjplSAZQmP7qg93Ao3FN4pzS3hY+0fYr8uZZqI6twae53LTFnGqWMdf
Pf/rgBAHNHKz7Ke+YyQsgKrz0vBmacw131Q4mW1HBOmdOAM+QACip8j9yA5eQPNuyX00XkgRAE28
BbVdJGSv0D+93I+4zNc2fpKxoeJIlyRKodUlMkpA7dAF9jvIKy/7CzbE2VzYbUGmddjHPA7q5t7u
bsfVGOv98iOz5NetgGGBcbHBuoBtkbMADzQMhMxeT+OOrD/R2ThYnMemtWIkpEDQHu1GIA0HCxKD
FKB4cDrZiL+BcTFRflor319s4f8JLbFcKiupawoOPrRxZQbIohG0trNPZzz6SoSWF6AildieDl/u
Bp9bl511ZH/4CvxVknLi2HN9woTIMHHrtZeq+fxB5K/KtSkTaSUY6/tg23DnxwHYc8IQHsjcsbaE
FPkj1TklMKE0Ez/XHRujnYvI3oWV8yrYw+7qgkByEeFd4EIiDgZI3UDQOnT8X9IurElZu9RpbdG9
NeoNQRQAOjmPC74X7aV4qVeUsTVwaTWjCpYtviVr4u+Vr75OUP8jVXhkbjhGz3xlaJ666CiSrM+e
BBryNlBGeM/aRpMn5Xy9EkW6O3DRg//xjg/LkmgNxCo7y2v69BtXSLeSYbIl4Lcs/7f+V76v6Snv
CsTZMFT/hmApUH1CEFZVpc0pu5Kj6Oyj8HO/BDhhNw+UircVchCMAPA5bbA17RuCVWm/9+4xS3Jk
Kzh6ZUeXeDhh8XeIOtWeI+ZizCLPB4431UYC80dbjMYPSDF45jD3xP3Fn5mlYHy5DUhVTiCPOyha
PN3Wr7LwsYTJPbUP+IEnGKtnGnaCb/ijbKd1kTbEEe9l41heoPaGZ6elBfsdS09V+wipT92Q9yKa
voHkT6iLv4NX6dZQ4XlcBF8iTe59eyXOjaW0S+YU52Kk5ety1c6DTbVr6+tncTTNzmzlojttb/oM
YXpass6eRubQv+T8yd97GOZAJsY7cb7SJ5TMFiVXYL7rqF4zXFZS58qm38tcpkRS8IWGN765mbQX
9ErI/MBRESYt6eo7i6Ywy4iPW1n3mgJIGEvDQxljdzUKcx62SFrAOINq92xPi47/cN3d8g3sbE+Z
Fqt8IPrc2Xy3Y23NPmWQgMS6f0Nx+SFJI1RcrR5mmimNIKFqK2y0X8MC5PHFdYHNTnnX5TvTdK1e
cjoOvkLdCY1W5hkjCjwiJivdJNJLJn2LxmySS2iTNVao8U62MJ+uHCb1A6WqjfuIQyAU6PP6c+Ss
k4iZhIkuHIUHi1ihdc7xzxLqf+GHRiHWlzDqPB7M7PQWkPxG9WM/zvRQePym6vtxVRyebObTY8T4
UgiEO22iZZ7AOYoOA5nX58UwekAPyod2FBA6xklmz6Od6NXKc4Eh5GE3jByHCoUEyOkNjyG6a7NX
k/EwtFq+e8XsqGWv4Kz5cLcQWaS2/ehPb92z523hfTztUjsazWZD1iyyQqUfFklNbzfe2wu5BTHg
pKmoVV09Gtx1iUxA45zWbXW7CtN2/63zpRcI5bESM/66AObsRD9r1+3K1MXHr5TMNnqLehr/aJRg
Da1GtJY3ClVSYxCGN8cKKuN/qXmlCv4Rv1jYwiVFcu/MGfsBKTNhy/+gnX6ocK2boFu6cc4BAxt9
6QAiyQehCF9iIUL2xYG2PLecZaKbgNimrC7OyBkenSZPr/nHGEVzw/SIlO8X6DzCC+WGx9lM190l
BfxDSl51g2+9laZU3r3eZkvcZB2xDDzUrFblZIVVVaYuCqz+PPZl4e3IMscT1jzg+SfD1VbT5Hok
XEnjL5gQ5IBSGz6YctKOrxNMHyF59VwKLfs7F6VmLse9wEfNaVCczgcegx7eheJ85f+7+D3QBTYu
SHNI/XtB/ZeszlSyoG6QZybA5RQSQKGarbEXpq4H0I9QAvKOwLFngMLqvhf01b/46EmXguZR0FR2
Bf7LQLBXlL4Q2cXPhuTjB0Knc+INaKcWLnMgpM3bW0VlHqt2eZLbElFQpr1b+wsFCKyVl7koi9pV
n7qMJtIgmp6bGnjCZqDJvve9+qnD1KYbxTznVYy1xXRpLISfT9oNTKUnkCCWCoxXq5KvzuUSao5x
9SPcnCOx9z7l3NxCEQQJbsyqM9TjObR/1AM+LCRTpflRv/GVDBsg6y3X040QmSmzjwPCt/E3OnFd
gf5q08nmA47bqGCqJj1As1R7BRKNm5QCzS91aW+G6SS63XC2exjM0E2+j0hLH3x00/qSJMpq2F/v
uRufEbeXcH2ImsqhV/wckqgsiB9fmmiHuq9tK19dVn5QVkHkXGRjfuZCxSilrUf/md50j2fgZ0GW
G5dIij0+aCcmYz8iN+hm98IUWyMlHX9SajKp6Qavek3not/GsTiNiDFVLLiSY1BgDDs+xy6w8SiY
OCNTOLTr77kT564sQ/Em+tiYuKTqnFqYa2zvV798HZSUWvJvdrdqMQqFO3PrJS+kzTLN5uRt4zsX
EyNv+IXAQWL7PQm2zXloG7Yy8yF3me5ozFWJ5csoXx6S9O+3li0l4J1nSx/g7BU4TLqSUqypVMYE
knub7DpJk1FBWQMP9o7sqoY5z/iQIb/ITpw1P3Q/F/wIv85uSumUBaiFFND1hVdNI8WoTLJOC7l1
DIJTS910uEOESYgCom1npmsqxItlp62RGdhNqowUbeH+I7Xgd6WX3QV6vQxK6emV5hMgzxoUpgl7
1O1VjWoF2+kv7apHPUyqqBfj7KhSoffMWWCI123IIRUa6HYi9GxsH2jrqE+SI1v7Wj9mdTP+nUNJ
ZRfQcYkDbywq1T3bqE58MZnsFDBFTEDWn4Y+zXvzmrwjijtGhIy7e0Y362YtFKexlYRAuZSZwfO0
yJc7rVIuZ787fCZvWwzjinv0AUrJdMW/M5CWFKQswj1y6m92bT+IyHvlXigY8xqECyiBPtxXFW8A
9rMgsU6iLGYHaVBCiGFJL2kPMq8RMlIdsJo3UgYhWM3UzK/f9Q7fDKsbYq66hkvEJPlQkTU+PCVZ
KtrMeljBzak+ctTXHNC7ixy4Kyb3b0yFbOhYkfNfD0Y/sMGOvK+sXZ476jcneAlja7vUqVu0CoO5
8DUfXu2loRe6m4njhrlLAe8fznSHQxtJuhjd4QbAb8FljJMfmQdVmu914iXtldLilydNwqurqpxJ
up7Fmt9i/Byv01lk46mNnGeL/M3+qKMoHO1ptO6J4JxgJpikNBGG9KZ7mjlnJoSvK+9F8AnJaFmx
W9x6pkgIfUTF8jC2I0la41qlC4uab+p9//C9hV7I40ZSnwT+EvjcOiTcJnZivdO5PgYE/ajH0Oc9
97e5hAnfnNE7rVUNdK9p+v/3oWb+8l+ad387hrClLs/FsrWtcxLeL+YdvLxOmj0Zyg1rBRECaPDC
ANhpn2cje+306y80Hq5OowO9nM5gzlrF8P8wob+YBLrcY6XvHdG4TU0/hAQ8rC7Tb35r5fxUgVjz
DVZy+bbdbbodbLM9FopiHMnLL7nl50nTqD3nqh5Ima1uSGLk+6+2VfU8oisyVolAJ4CYf2mipp7z
zYgyc3pOCpTp+HxMSk9lsb94mqreIMYyTwwvkGqMl5JRZzEKwYJNZ7QihwxWLOwb9zVNSZRoiZvZ
Z+FFTkupYYWFCVg4uaqyrcnZ4iX7rvHz05xV8ka3BqJFXF4Acj8Qk+qgTj5EEB0HKxjOUbTd7mRT
lpA7IArUgLRJDbTT/q0by1TOyjYC1u2SwWdfecJV0dyjA5RIPi1dbj61WxJIdD20uSRGi4ozNwQ7
IXCDE7hWFbFz5sY9AshgSGL1/0QUqw6/HYmh7EiCMmvVmrONCUEdJ1ZTMMY/0NmOtwf1IUlxnYDv
Rb2Tu32EXDk6PE1K83wflm+BdyGtKfpfjh841tMAnHAGrGrZQ7N/QcIu2fx5yjlEY/k/MVW/nYer
yjMrX6fYnQB2/aUeyDRVRDsaC/QyRX7trj3lEpB7T3MEp3NphUg58PiM2WhSHT1jlIx6/k4TR0O2
20Pmm0oXQfpQSFfM9WD1/dsx2rjxF/aAApRrqXrsqSckzV2X/kmBKFVyooY2x2r+q/cEUUcQX/eu
oL9aVHuIHYewcTgcF/KUsWVhjb8srItzNGvPgFhedfocdxU2fjWyXev0yzwKV6ST37dp4Rp23Cyw
NLKTqKe5X1dBPLtZ0xg2rXP3EBvEUb94h0TAvoNisyIMp7gvkUwA6/2qikEGJp4YtvIdkc6r96Kg
Jnk9sGtkGB8Ssz/EaHREGZNQ5Rrs/G+1NA78PffQ/bSZFOegvwfYKXuBTPnMUIExwTgs4kmiJE6b
Tp9HJ0zLxXY7bcpO/YZu28PxapyJvTpaF/LXNPZqckFdwW4AxwDuRGfoIcfBOUZ7X+EbG2B/Am9P
WcLWNgn1Lg+/njVJRBhTEjsw10MAfE/TZqbsOCanrUK06ttOyeoV22g7TTauCE8qODsEGgNyUi0D
SwMYDCSVvFvbjTsP9NM3H2d6xR0ggQJFE8r5RnLTPHBrolmuYevBmWl61EwTnmMw4OoSiwUWTXj8
QHNbTuyNiFZLTlLOGfnUFAy4RNaNvW8czMOUCPNCagxvc0YAm0kSWyZumgKnkf/TKo4wUNixpZST
eoCzxAIjfhkoBhv3HWE6WHkI8OKDcNAUor2LJwYVkSZhYATHGG/CILI4lfvJNqcdq7pM+NObmjSn
PTxLkZfW1iyIMn0br+fRZragAb8jx99ZxeGcxDZL9qyciYD0cOYmzo6vZFYukLXmQbiZiQzicPGt
chvDEEUQSTJpB2zFML2WdKX45Q7gTV6bnvq8x7SjdX+fHOqmTL8PJCcVxcvXyIljp+cq740Hl16w
sxr5OBTRwKUD9rM3mttkIWf3TvGa/BYkEgONPsz1AUUvadr7KckO7U4qIIZTSvt45dtZE4xq8UZ4
ajSigc91rv0SjodCYaAld1gNrgXovvWxp4lBD0lsyquIKTu5/LnBNMrGX81B5QpwiK+P9ji1poME
TMeGlOHnhFrI5HqpOZtEjm8yUSL1U8a3Eeynmx9ErNk413U3MKQzFORJ1UZroLxY/lCYeZbUlbLo
bCeURQvEH4iS6puROVb6EKQZ3wJN5XCRe5Z6ZwiDMKD/HqsoOFfx1LpqAu3kyLgO/qkF0TENjZTJ
UWJOR6LYqCmkupeNoTlflnpD2bTfyJtOnsD6luQzTwlliIWh6qPh2yxqsIQ0O4tt/MZacwpWnxBa
beXch0/+1ZHpvIWqacaeQAqV039lHAc4uM4qGkQlBlSWtYhyjQ==
`protect end_protected
