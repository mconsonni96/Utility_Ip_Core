`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
NXQp/ScONdpualhArNZiVbdgOaFx0LS5vQisPApZVFVr71OY+tR1u3EbORoTydixrx4fIss3qxEh
isj9P65bYGBGIlmkr80jYOvOWizs12vEKO/5isDQ/8CLMNonqo3m8OPMb6+SRzNz4u9m1CZUMd2I
O5mCWHWShDyNX6b8W4S75a5dKkAx3tI1udgcl1L5RHV3W1FWAFfao4z81BmzKPB46uEEivpHH7nd
mJyCxqJMSMg1uLU03OsKTgSvv5jQb6T5sdQiPW5nIFWgmAViA8o+25krck+GRVCG5xQXf4KWQanB
8bVrcA/sYAOFFTA9n12u8EZ3gh1Hc3R1Dwc/OA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="3XN3XWPNrbm7XUkXhqbOouWuwhl/9SrXJ81fTs1qeI8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21040)
`protect data_block
XHEGTpMiO9TfXr1xaVfYbrhneePX0mVedgVySESjc5QnhpUjNOnMogN1i7kbbs+hN5UWxdhO4w6n
obFYlfiO3q0k33VSHig/v5n829GAjchce5nJiZPJ5N3mordnl/WVhijtrnrBh1WSbdYfuIiGKh4R
ZDTpFgmkirASYR7xlkWw1pHu6m++dor8IYjHWyrWaeGXu21rjo821H+0NrEsZcm3ra9sth67D+bw
28stXVZ18ygGvPbrAipU1vdRHAhPKFOhfGi5Tu2cZYFq/DHdg7P5GzU+ImN5iFV7IFZRUPM+soaS
hhlx9kaEA/KuvVLEWuVCp6eqdzL8tcReBEFsDHaTgohEN4qiGBSOWYuKyAqNx7ZguykroeC0DMA0
w6fUPttXxJ7E1T7KoXHWbfrFxww4BYbT7xYqmuTh12ciYBNPstViU/7O3K1LkMZZlHE1k1TUKlR4
R+FWzLlFdhe8hEZVZt4ig+XddMH/5NjzfP+vRy4NqW5hhXWjEW5DgW7VtBfvsDhl2wkPxqiKGCpY
uXNk7JYhbaw5HM1UcTfWaA2laVSPneVKXvd/FtIjh+VlOxVS4PIiTUX6hK7AjHDIwgrXS+D4iNCY
e8QpYWH9JaYBKGQQsgCPhQTeJAaVUHdaTTr5doviAkKY1WcDF6APsGpcuha5Sv89U1W1cLa6lc0D
5aukJcNUQsjTgvu1FWKSguIaF/KxKGTwsuZxFaPnwsGJagYltjSJcwguqCe7GPwzoHt53r4YrsTm
QY6HRKynj7xTFwVf34jkqzTAk4uIIcplFTTt2TeFtCNLTBYJnq2d/usKA7nAdw7Ixs8AyiEvnJuJ
2/Xv7kO21Yba5FMM5jDy9znzSXrNMb1PTGgcP0TKdyKNsKBKu9P0Iz6zasSxqDuieS2hQT/ZTT6Q
Tx6aJsb5Sd7KKUhfFqQnwuT5AtmSbOTYcdGRbax+nDJNzaNL+nOPSj1YZxNBm7mfZYs0NOlnvV17
YDlY4ogq/9mkoWebbisEODIUAmNyv4fBOCrp6f/rmHtwHXgnNXIaaM3R3Cd8VNogW0nTrsRUtpLf
RckDUxGo3IzoqPrbRBiLsexTDQzyiptHYNZhKMsVUU7eW/mDC0UyONRbHPv9lUt82peqd5Ky2Tr/
a3YcAEQaH5woyoyf0Z4g3GDNTDf1kLHMFoHyua949A+blNEjyWF85p2YyRQr+zVoxFqQMzbPnWJ8
geFob3DnZRBO75k27WCqWA7qNRwIuPisMsNfRUt11htXSzRb5PXrg0jAHdge82klXlmECmwRaz1Z
raZJG8IFwOwZn2UZ/6QwtTk/kpFBWwy3rtAVTB65DPllDjhLNy2XN3p7cgfmP3e64MdbmvUJV0Za
RXBhBIlfRes/5Xvx0Zmen1CBaMyrTMgkeyJT+ePtKp7avu5OikM13QXvyLfayOwq2hZ7trVX+KhB
34XVY5InM2Kd/ljAfwmP1ETJWyt63+YistQQhmYOiTjMK+ZUtktRk/AGI8YBgoznCgIqKcXY1xzq
dnh6v/RjKtiWaL3pGybVXqfOkr5x/Mg0c9KWgMUODLFROxsOnu6E2FyNpLDzyn9zE5KIllYuequc
5eSP4ba3mztyX3nbFwEgUR3Ka3PKO0schm5qxxkkF/gN0V8WadssHm/WJCPejpVZNUE0MkNX5i93
3qY6nQQfZA/91a+wZHx70o/oUgayCCtXqhMHulfPNQPmPElyi7f+DqHztNMVvRe60pb+vgOZafZT
HpArdOKKx8nUUrcmsaZ4FmP+y2LsDGoOIkqE6I7PMqVbaxKSvDXSuLTvcTUQVzFfA1ecF5BOe88b
aj4dyZNVZ3koiBvJMvoIH/zZAHoGdnNHEESTNoq57K5kMjy7anbU+VHExxCwkf+Avd6tEmPHy1wI
5bxnZ7zUIfWNVpcJuiDbDpqU1Y6ZfYcyRES1R4EKoQx1p39nVo1gij3XwAGEyn1bR4FQW37vVjJR
+xhSXasClDf8rbodDz2hNJeS0J5GLx+95OgUeQV7hk0rxjjgeHbWh5NFcZTC3YOsbGFiZzFF4Cpo
96h4aS1IczhUNNm3II0CdWrBKPfQB8kSsASzUIBk8qOnifeP1J/evFUmz9ZQYke74blW80lTPc7J
SxvrXX7KBrb3jfgxI3n7knx9GqBV0NL9ZW4LqDHyF3m5u0+y1AZiSLa9z5nX49sj5PIPf3sz3YO4
wu5YxOR1oxheO/auWml5zwTAKmoY7oX0QDKdgyb/qepq9SuGLnt05JHCX4yOafrFl5lPJBT9wyfr
tCUUndbnSn7Fo/83hWrnlpHs6WjqvDch6jli4LVeZuRBHMLhqU8035uCpGGntX4v5bsqlbOu+pPg
qPKLrcLtNVx/9r6MmLY15k3hhjfZHUs9bMpEadcusZL82J/fYMyaeWLWua116L3pD146efjSGuaJ
B5h8paQW2rszBKb4x4P9RenX9OAoiN00T2gD1OW7BQLZixB15TO35gHw8su/4DNPCw6Qg5fH6n8c
gl2Kr0r+zaBIOSRcJTfTr4obxrOo4U1X8GZbPoO1P2sz91eWbThsBbbKX3nXA0KhTUamIpDooU8a
lvtZlHNcAi7BF0Me5rpVap1xBgZTw80958BPOoBSxsyJ0IosXpcd8fMJ0dJcEY7WDkLNKBtKaTjX
xWeu7XQCN33RXCjjlBLsTqZBxjrWgY/ThgXL0x6ZyFXfjN1o1qEYbfvd2L+u42s75gpr1K0BpbkQ
Rh+i6bAqurdoEiUO3WREeU5ZL6pP9Q5K4qDAQJiPjQRauvtKhLdVPB7AEUr+aXiKKnPH8Kr0uGMa
MRBQHSUVuk2re/4H1zLCJbNjDDd7LsoMYxFO4JedzpOPCFHx3hclvc0XcvHJMYRQSJ8Swd642ugL
3hmr/FvUD7cwaAoz96X2xdfwIfiYzbwpjwYeU3MYw19TnnS4l36oSQOPccUtrjEwCn8d1tnaYcMk
hetIjkBamQ24cFf3YTx5QDxXQiBIlQFqnxhGjfBo+vp99LXth6lTwsdmypTNOQCv5E+N2/B6Metp
1ueocf/Ajg9rcqOrxwZM9gkAqF6KeIcNTtrYxIWhuGXqtrvMQgwkhSVphFzUwZttdzB2v3LXgrpK
ilrQ2m/LAB3e/dqN32ELmGX6sQUoAkLVNTPgTFEqbdOorRl3Ri8Sz01420uO1OAr5Mj79hiEHbCj
x6NnbiiQXzk3YYMRKaSayQ4idmcBtohH3qj+CCALpL62toSKZN/flY6dhldPqO2SZDvSWJdTikBe
9R0pP7VMVpROA9E2eokt+8fe21vI4N2Pol28OMQpJoyIMe7yQOW6Mhu7BkyMwC2fa4bQ/OYPGKAY
IGaM/1mCyS4+k3okqgcHTVXzqV5ur9XfUxx1sYWXRwtlRd32gq545L91eSotUlxDid3Lqe6xPcei
TdYfSCztAjNgVEB6ilREGjzvbtbxg5VS/nVPUK9bW86BJHqNHTyqvMEi+kAAi9P4Azj3rcuG/YrZ
qrBHlDE8IUCsvTjv6tsq/Z4xTpQhwV4FwQFTVY1fOiQbJKlxktlxpLudwH9NhY72RY7g7xoPYr+w
LfwP1hL9tq+9FPawh/t2Y/1ngQdV+742aLz64X+PT51rDVQuSYQUp7qsPqRupv1As+JAZh253pqL
2qKQcRNMxM9Az1M67IGh/Padx3LcQgLtLmtkXiz31/YfaJBAsGN0gpxA3y30UuM2QctOgNklfmpn
kfV/A3yBodTVpQ19Pqc1TmgOtHJY1xRfAf4VLRIIzbpkHDOPGf55tSFvI6F/1Btp2QgF3EMu56Z7
YDFp1XpiGKbKneNr5/0DioQlnWFAP2HuCDuYLyMm1TXzDk9IqsceXJN0M2KudhQXMJMEFoj/QXbl
PDNGkRgN7aUJrCS8JhLXyCxc9Q2QjGQ78K0Kv/zbhZ9j/nnJzDlwXq0guR6MCBajhXnMIHFiB+0p
f660N8HeWsd+WY6GQlvWUJoaPda6tYHQ8ZbokhQF1eeZfd3EpLs2/GDDQSJx1P60QL+ermpg0ajQ
Tw73Igia1GWzE5VjoR3vwAatOL1NLTCbYv+xRSrAybNCRuXPXqklWrr2GNm7ZR4pI1RGgpySMypw
bA0YxQBkuSPk46Er3VMX1ZliaScE2z7wMuluLX+OM2FfPxxFwCdvkCnXqfzi12O+65s5d/IJTnvg
Knu7s336AnqpyvhW3H8bqbmoaG8kUTAZNDqm4U9hHPglqBn/VTOFjOsWn1c2DQt+w5kiOO7oCTNT
333AB0UepwMr6o9v5hLcYNwltxqaiTj3LeDWWhKC8VD4CJ0WZdz9Tx8V6euhV6Fy/PVC2K+fxM9k
UIPbA8tlIjajUSiXlYUdo4wYWe9qEaC+wIrL05dSNRpSUGE1zMaKL+Git/io4yvmlWdokyB7c6MX
b5Z3lKj9bqtsVaiEASTrxaQKE8zzl5oMsGfPPl+7FlN68HN35P+FYGY0zCOgLfznnJWpZYWPyavc
PJHb5X/41fJI4hhs6RPSV29Gpsv541QNoV+WXz+QMNVBDCB62cP0qvTyQDYpyrVYUFATV63zS6oQ
ClVxJcrf1CFIIaKU+Aqcw8p3OYu2US7qc0fQTEQqwHUX7ZU6+XNSCWtPTBLvhMNIZ9oJtnvnUyWi
te9oyOsN8xRLoXmr5zR4XevbdlXnw37ujTg0CnBrOQzMdvdv63qfi8+EYVCtLQCNsUwLPW+fieEU
dQ1peWaTsZVviw0yrUKfsbDqMwLGw0JcviSWEcGFMsPsip6DkJH5VYfXg7AUa/E7f57PLqQXAlO6
lJFycDx9benW2dhvjEKUCBS2HuedOs+KC9A0oQ7xtJr95puoEV92F4KvF9fRhOcaw0rnZ5q0cEq/
SrzbZfNK6fkYsnRE4ROftRohbP5PcOAUf+0IwrH1MmUV6oH5ta9ctcFBVP4TsPeHJRVV7HBuMBdr
M2XXVJ+yxLf88u3G5kQ6PyUQ9rCSHDJTveb/EDCoref1J7jvQv/b7gM/XaQQtLD8eUtyb5z/RwGL
Ok9fvXj1ykJm8L8nsEmPQxW9wInqI46wTsbMPL1V6Ei3IsqiGn9t79SiXtsB9Nd9GdUO/9dzf1NX
q9p22rZKzLSnAGqtxTMs+kNa2jkgnkU3zZliVLyO0Gy/eMSbfphYKi/rBi9i1nFnaW+jFIDNiCuh
gr8R2mg4fxn/z6IJm7CvCRizxSUaGhkXxk91v6FJy5VmiHY+Nro79z6jA77Dv8AF/bDIqBma1bw3
UFmzyY3zHBcMC/YJnioKDVS1ZYYWA3EBSK11dhG3PwtcoUDGjO0PuAVO/x2tg++1AVCOMLiEf+4G
z9yorWfNOWIub3T0u6BKf1KFUXrmuNjDmHD6JJ50r/ALohAuxbwFpP5aRM8FpMKiVDGGmY3EgXNM
wxISheBWUSOC/B2zNSfO+nXj7Dj5fuV89Jn+iJ6b4yrDHOoKsbs0F5cVUMnOALoR4FaDVSdyMl8h
sLRk5qBRhK/KuUmPvaDqQ7DOjDCz41jBw3pFJlRXN18VrF+BPPoIYuuGXEeySz7JIqj1E1GoPiOg
a9yy74dLHAG9fU+0NC1TDKrTohXorpqQ9FnS3+0Ez++ASAeaU/Bv+4laQkMyLtEFENeEKwXiurQr
uFuCf9BO/32Qivft++FDwBCK1/z/OkaNSvcrhevB/92XgLbyKTh2G0PRLOVi0FdJ8gsH5Z2/O2JO
76U8zIWZpj13FNMQD8tBsSAVvpLjdIMisjyfzeyZbcPk34eJutXbax6hgCX9B+e2CD1uOsC/XzS1
FxomkEFl0Fd815+cp/ZJVbrbE/IXCumTpTEdyUkwVVh6wOqtc+xzryRxXqr0KFMH6+cHVfpv8mGn
jENHFDTTzXhOkr+BOcgO19VzGah53LWaCoI1C2K6UxsMZfNdQ+31qRLN4OFy5mgCegUUVISaJ/Gd
FHi3GLhblsqb3/slM92oMiwDK+8z4vcfi0TLTiKjPJjr/O6MWdOnTCb8PeMwUH3ezVLGEpDkcMDL
OgPeGNnb65nwPud9vUVZLnt1+0rl2S/KMbLDT9gZ0zRvkkPNMyT7nbYx7MDBPOkVJ7/XS5A3Am0R
MQgoK14y+8ccwKQ3jWL+gfiV7dHNqFwesoX867E7zHDM+PYTaXGDB9FsYec53B5BvR4sXRp90jGS
fURXhCcX32SkIh3+Hl15Igjy56hlHFyL0b+lP0tXWgxw/sro7VPysI1X+F2xWyHGElowrBloX81x
l6daP/DTGFv8HxBAWZZ2fqksmtkCd6Ka3zcM9+JRyMyoGm0ZfpK0qRJakDkH+8ar89D2ZqnKTgHr
duqW2qF/UOkCSe1wwfTiivMP9RDa5p2vfQOye6wbr5/FnbGn6LUk9T0NTmLWZ4evUrEEz3eoJ+QD
FaLwzeOIW65rmlS6nbxt/avbE9NCZqwOLTtYeR6ajV9QxtQKwdq6ZJE6QhEGuQAozqxWOgHW3Ai3
d8ZiqipALlPUSe3UqtYPrOAMXhHUn3OmE2c672cf/Awr0usUJJI8+e+k1BxQKkHfTlVG/CVOAAJD
9Wj/RXnPl0ab3SOlw4cS6VI4+DrSolZf0SaFRRaEQc2rrlcl0X/v1/1ZME7az+YjhDuBwcpGT/LL
m0nDs50rGqQxkg3sipAr7sF5698uRB7H3/8KETqvRaJFXlYl0y2/fbb1oAhDDH9X+mYzm6KRfGf2
doUYG6OQ5dE7+b7/OyDJOhziA5uxcELDPlil33AGsoUbaeyeyoFkYO7xEwwxbWBLG91LQqiQ1O/W
7QqbCgkJoTe37viuLfU9S1hKZXVT70OYo8iOFWZGC0XGxCxg8CNGHtUXGMG3He2+ui7LiLbDVhIC
aWWvD53CUkJYGgcWPyUnKwsdbKmxJpbuIza/H1iH/3FkCZsx3WQuM8l7UEnRwgZeaDgJCQOa5Lqy
biAP+ctQbA9jbgy8R9BVT0rjvpbk2wPL0xeyGpGt+G/j3vcgRDFhhU8w7+hTGipb+E4cKnuLbSyr
3pPaw2c6fwecSGJyH1vOihgEm4pHlklvdm3ofFNAeUR0yMeRJTzqzs05JLanxOzgWWo4h+XXncgK
/22iVpe2/Xkoo9yTm6OKcU8NbCbkYwlp5ki7Y4I/rS2sjk9AhyPiLn0Qgu4bzuzhB1ZhmcBy/8PG
JUdTKNyS/AcCPJ10tH810ejD99sREZIfOm0MIOjGlwF9HNJstjUGIpffXB4vc0QNU/Xv7xB+sMIV
+zodUB79TBMuxdeQgd3RbkAajUevk25ZmsT0UrSZnIyQ4h1cpzGcOjrr/Z5JoG4WpcyFXt5JbY/s
2ugPTs/WDXFYMCv9FzylJ1cdSc+RJZ9q5xd7ZaG7Qr1w+mNz5NlNejwSi1FJYeGwVoHJNY/kDRD5
J60eMzcIBGl0mCSYPCqmE74BYuHPErlTUU9d8J+uEdGQZeZdnRvwgD3IG71EgrgiHmeGLWCo+ucA
xwAO7ie0DuEA3sxDYra2YebJh+78YQuLd4K9MBXSqKN1D65HVu75jxauy68UFVAG9qembkSa4WhL
PXOT5ZlFp6j0z2VWYgH6wTuSUs9FiwN9db3Q9iSXVEq2H33EXBPt+DpcyLbdJi7+GVCK53tTcaqN
oNIO1Q6mmo59b3z1DFOXw7zK5ZVImd2aXUZVmSLKb/y/adtJwHUf+9chz8BzFnzpOnF6XMDKQhx3
G+cGFuWvSEbwAc16yPEQojzCmyGF4ijoL2+8zKzLwIhpuHe4bWAuD4g27Gt63QaPV6CXCo1Iy4QH
+w7jen3SAw42V/Q0pFEK/+bW7nP42HifdfvjpHFL8IvKHRfhxblJLTipt84hokKu9/7BWKTU/3ON
eN2kg+KZn+WfGpfMpyh5LHsp0A68uwgQ7aHYmRWGzOZ2B43S41wbag1HqI0Ad7EUsn3DhlnAIubv
IfykO/iwUVdegNPhh2TBDhFNN6TumXCylGoNirNHFhvMD0vKLcWCXwbK5aiTx6u7ICMHuxRHEzo9
prIc6RblhCBWvVtgzmNbuCuAV+l4auIt0mZI9mHEVHwQWVtfcWejb+e8n4il8exy6yZuRdIXfuW8
rGzACGYJwpaYeOr2fnPtB6CWLOvrDrAfUkEhkJQJ3oWdn24DBg5uG6rR5ssXiZlnKVMh3F6MdedQ
iWAG+QjIX0vOAc9RS67kePxRrDSrrtkS3xfvq0w7QoRPt7H3s/3rzmD7PjyVfJWdPLaeEUVNVyeP
k5Buj/3QOCGEXaG9J/EwM1boGHYgNrJxlE/2JrsmG9dTEPzE2qNavgKtVJWTzyiAVPjV/zFhjpQy
N1Kto7M9hw4m4ZCM+taACcjezjsdPuElA/YLXQ1ZVRO6isBKbBo1HKR5ZWOZwqGH8EMtZFVYFYIM
v5vOaHr7wn4kndSV9lRNbQVyOrvf7qPmzs9uVZnEAAGjJk9WpsfPbzl/xrSYo4N1wLs4mE0lF3Ks
nzFJw7UBg9ypOU5rtnFAzFDazJBHSd7clrgP33PHH8iaWuKI+vqTf9CJSEk0Z2rFok8ZNjMGQPWp
qhQh+PsaTup0ONdssZkTsWXB943944Lmz/WgtvcJlpzErjFpBQD9DTUMXqva82PTTPj1EwSkaD4D
GT71595lU0yaOxEtK7ie7exgqOsNtKoLBWvhNzxuQ8zOgueBJekhCCXdl35wOMsaX+l62ES1mNdA
RNml9r2d/JAinJqvKd3E5gBLySaRiHTschNKQq4Ue8JtFlda1Ni3w37Dl/A1eZN1I5QS4oxAN/OA
IrUFunyLpiKofT2G/PgO0MOi7KYX51ax6XJ/YiOd+YDqr8yU/GosIt1bSDPLLXzPtswLRmK5/sfm
mHhPpbUpVoEBYh6+ugV2/dGz3x3VE5GGOPfBGPonNhVqVmx0hsYoaoHA/G/o88KjAO6dF+U4rKYK
/B4cg4PigHjpa7osuxaOPXX7v2WqNgPMgDynslBFxIXpF/puIKz7k6a20Fw5l3WsemfzaiAmdH7F
3JAHmEr91i15p0aXXfwc4YnLcgEWyacW0kuOGomDtj88SdU1YWZjFfBsdcx7hOGPQTMec4yAMDxy
TQtLTq6UeXErov2TGwFXnTsgoPheEkcckKTtQbTymUGau6IJhTQgWDr4uZeQwbcQierxzDLjK94w
AbBsLwsAH+Go4+4oWh2POv2mJjbb7YVb5B7ck6Pu3WyKImuWrKXd3YIcZmKIcYAlvgGwFR+KpjHm
nBEkBO3l4OuPN5kD9GaoAq6KTvdO6LNzAlLgNaQMwmKRAkq+JFnZo+rRBZl/cAIWDlh3C6Y4O9UD
0VL/ovd6CtOGjMv11ylAYdtxYpbBujCkHsEis/eo2RTTOhhhQOk7df1poCMtZ51Qk3Bu0/kNxvYs
Atfkz641P+HJuCNDPqpi89Il5FsWO3KJpEKr6gVdXqZzcU6qig8XEK4e0tHqO+w6d/CEAyvHsSFe
5v5bXLH2lhREZr1OxXp3ZIFfZaEDnzuS691SFbozKjL1klnBOUzY0Jt7MNEFOMVbP8im8nKj61mC
ElAECsqIC5LZ+RyL2T7N+M4ddX1sugCBNsAsehBddNEacaZ/qgnJSUB4cRdZUVySuQBVh+CRBDEL
XAsyxkwIm5APmpboTnjrFQ+PuiZyFafPgHHOXHbz/TsWmHGrZoqmnrJB/WKLoUKxHwcwf+QxF8zr
YDxyJ7WsUZa8xuAC2R9XYI4MErCfC1UGKK6o7VYFkgV+GqmV74Iu7Qy1MrJrpcjkt6gsTZNBu+/p
QcY6hN5d/9ejsI75a9TDl4VCtsC1p3B5W90B3kN3nyOPl4pizsAqxOi4RlvIPqWXxYtWvn7/URmD
g/uoe/hLnS332/bWfOqEMeigI7uCAYFw4i8Vwu9pZNpDg6WSzhzfcOilzwT97VVxtqvHBvWj/j9c
q/LRgJEuRCas/zvY6snUxbDbiS3IzyHN3FUGnK61Gzvp7mxAEKpfdV+LE9KPGylCpemWGE/zqzxF
wXwpumfeQY/6FtojARQ5ProN3oDO03Tb/3yskZZ55+qJmAzBBzBA2L6C2Mt533NLkFquPWTNujhL
1P0mcr37cLoMiy/iG6KokD4Gz96umZpIaiq3ytGmRwt+jXx3xRq87JSiwHtX8n6859y/cXYLd4Qf
NXVhiD5wCh8hjoHi6nJYKr4dlZvAxdH16fCIhtMjUmAvHcTWOnek7iMBv9McKge3rQNDnLIXqGW5
m/fsdM641HI68lUP6YlQmj+/j3t+C2kDOpuaqxn5w8ywmZaWO38B44Fk+X5eoi8sTRLsUZSRF9ZX
jW2mSNdVBZl3Sdlr55lN4J8yqJQaUjpaLBdk2gxFTfxK9k+eJMK38Qh60yxWiowmy8Smpxr3xaia
AqdV0rlEIAoFhEhepN+Y49GHiMKYCSKVSXPQcugPT1NIRMlNRtMeSIx2Lz64d9eSr26FlpAUh1GJ
e/0QRT7lbwNcFqY9L71Ofi6iJAml/yXCrvt9cMSrTIcv/XUANmKk52SlgmK18pdy5QsEfptS+j00
5q65WH9EC/mQXwgRHEfj17ZRInZttowvSc7AqKnOJ45X37zX5Wsk7Fp9dZteo4alygEik5fEkaUz
WKbp09cQTwwb3CWSWAoThm1tDRsH3gl6r/apWYxOkDzsJA5mo+TY4IlZW8dDNSdtkEO492GXXpfv
wx1uZ885vaCQaEh6/angSbLiyJ5ETeAclqxeZtgEzB+gPk/lY69wgCUL8IYnCFu7WlyxMNUAzHqb
nD9j7Abeap7W6GGhJ4yXkm1xxZjFs1xFlJg8UI1Sm05+rB6CzS34Os7brnjXsjLy2K874w/BDwAz
RVhW4SYDWHcKumO+LNxEg2dAiNipEdRMH7X2uT+4k02DOkNhICPxXuJq3kngEEPCvZN+5oiox7/e
FQEIw5njZ+D9GwSFcrsjqxSHDcgJi8lRUPbwmtgNp+ByGsY+R2PuURiXCqIH/6K+c5HBoTE/JPw+
I6yIlq0dnUYUQOzSEa0Hid3SJycSJgezxZsPC0wzVDQ/R2kSadBNHwECHmOv9Q8rT6eN7RlKj+C6
IEfxS+yEvD36O4MN3wZGmcab0TGVM0oVEgGJjR4U0CIJSuKuXu3P9ZRC19MDkzNWPLAbEroDOGI2
vkxCXGQQCH96JJazUWbZSTammUBggsPBybMzdFM2KPRuOimfchTwvwfTgVebaaiaWicmgIN8yzkU
Kzr1EqzHGll2yQ481SRGcUp9/HajZFi1jaz5zvkKQsL1pDaqPw4UUDWqBd78RNBtYkIgMmhlPhIy
/+pAgxvna+7EQwHkvOgsQsYeP28IlIoI/4U2MqdfdFYqnxVWwVnU1Lnel2Kw8zZtgQQdtnILQcTN
r7PLUevIRyvRW4Fz8J9PINyYYDCI/snYMZjBB7DczPH33b8FdNXJyUm6kPLCIEHyFWANQUrN7LcT
CBHeOPWK6n2gyGsKs1Y2M6/UkD0MQy33yDr8ED56KU9bJd0FAgy9XL9uyyThSEvrVI0A0s6EkRlK
DJbrZUuuLfTtaEjzmquDImhBEiVrKrppN+Y/1ueRhF+8ccjXJwT17IYDdkN1yNCDiNDqRXbz467h
6ip+ydP97lZd7u4TdG9Ia7cqBQp1cXurmJgKeA8rnFGXqPnBMANTJoG+1DM+Mp/LnsvEDvTlkULr
eQYMZN6SUexjk+N6GCzm8b2f4Z+EZSaSmk97hQ3tq5MRhiadiIiw0cUeziHlAMmBSkhNTFKJsYAw
oF+rmo3+PsypYNb/3oO5qmZYQ2PtxBRw+LOaZHPfnrpymJObc1LLreIo5jHFBHYj/6YskpLqA2+T
DA3rkulLNHtQJnGFwqU+7Mbya4yrrWtFNptx0H9aiMqf2SQe+VtlITYgzsLvpj/nyUTmPYuM05oB
6JYueozv4IZK55zjI6fJUpRrCA4yEmMxRlWWxszsR9cL7xrlLfZJfzFGXY270hFk+8gcwEgT/bFP
rM5Cj/5Z8e3XBkrUjVwiJ4bLAODby9O1SUr1PiEGyLJxXYnmq7LgXMHsEKGjCV2vxAlp8u5NLPJf
kHVPrO7i4dTYYieiEfH2QQG/BQ1tM0SfgvDEJxd/Emt0kURZRftXKPzZARTsD8nOQSbNgtye2iAh
Qk80K/URI0xd8Z+vcP7BvWy2/mo0F4OOf8JxGWvsFNrnT4kTYQzv8/a67KDdP8Q7/QrlY1ErhK94
hEwAdszIKd4vUO5IJrbCloJogLhg5FJvscnUK3Mq4/mg1Xap+tNIWtlFSz2JhlTnIWQqnGJS1aL6
LciGqXecRBfbcrpv9r6I3nG9LkPNVeAbNWfdBswI28aNzcRkN4nBNFfYA9mNVBD/u9tk3/+50zdO
f4W46q5TDPL4NY85TU6u1YeZErP2iKx8qVEgr91BbhMtvm+z0ulpC1AAv5m63/Q1G9s0PWjTpu44
I1MdqOATwz2VPsp6bQ3CRB7CPjRAcSeSKWM8oK6b30He57kPbeAyCWUiTg/IU1kstd1RzCyfy8Db
riMgOJYNQhFb3/ZoMO4LlhLxUtBLm1f2pt4/C1Om5RwjWjM34F07ix5rFFMDI143fViQphDqWDW9
SiJxcpPwKvq1y4RDUz+13g0uWwdVCn1E6/ugK+5lVBIHH6Q5S5QAu8A+9xlE9OI4oU3KLjDYra89
jkATQoVpx/rSPrjYeiWzN/vmUPi++59eMmVko2lz7G2Hat28n4ja6rVCBCec8viipBsHcwJt2Ds9
eGiCmvbrM8MVAOH7z5GyDu9NjxMEP1ZITEDeZjpBfp4H2Qd0JZfz5PBN0EV5mAyhc7jaOAefxmRU
J9BKIjwkdeA930fkIrbAtG63jy7hT77iUVQz2YJ6fdRlo/w+OWdRGmTowDGKaItAtkAfSBMLDPC5
xuQx/hO00gHN2FgDeYx+cVzzj9yGcdQDZboUXWbxMOGkCMTrdSpI1TAPYncsn+dvHmm+aH5NcgBy
Q1cpV9mELgHa+1Y+xdbJYwikh1WblUucB9ZKI1Xw5GhnlgipvaKh3nEQGd7XbLwJDCV9q58Uh4h2
WjTMC0YrVZP5R6/tTuBMiVUggndHVh6VdpsqnEPqJTcWXgu6uCD8+5mqtVVnv3jFHLFTxAmg3Qye
nG+mHCU/Vpx1XhxyJc/uY5xnVKXey+gmS9A9QqTWNNJmFQreDvlS3hlLDLIR3hiCFS7dAjL96Jrm
sbEuWFp9RqaO5eywgPYXXWkzPMz/BSLNHfrbgeIaDzLOQls1bfQRY43UWKmjrDCzRdjFVMDH4ycQ
6cni7SXvtfmpocAyG4hcwLqj1YaLgfowOd/1wb8fBDFG7i2qL6xE2NNHpnE7d9ZFJeqZQxKPvmJ3
ZfYQ4tau4uF6r3NF6JfoBOQormT+DzVnuAOWnJ2gdMYLJXr0CfIwjOi1/HhyGUy0CVdP0letoQOO
wRjoiWyU5aGzT2iDZtD2Mh0tBPamkI+ubjMYulhfQE/TrqCtQNaUUhGCkfNNh1b31w1j+dwWotnx
kVuWCg9ku7JzrcpJPN5HiBRJuQtf+72rBCCqeZlAkTjYgOwQC+QqmplixosKZKEu4Q15aLRgyfc5
MMZWaInRz/KyKWXcVDN0VRdb+lBu03Vydf6FJK6Kp4NXvZ7A5LGrFZEBKuvs8l/SE57etxsV0Hnf
sVKVXP7YxLSC/rXwD+3Hyl5VCeU1fHo5BEWdvyrsfNKZF4qvZJftnjeucCjmlI6TDtDEZijO5ZGm
3CpOWSa43R9pBUW4ay6Mr1dEJY6gBC3skuRw9gDCY8jBPP8pJCNc7/WrqiZ9YJN48lzlL1CII6sY
0BX1DvmoKrRQcYhC6fFGLLNmN9WV6wbDPLyp0h6082HGlPTg5KKeu3CpisIoAhpCepTRXGnEl92I
+gnpNQ3gXQwAu1WhnFMadCpc3csjYv3yE2G1R0vldAGl+KsgwaneGYLmgp/GFBKYLNq35RMFFtZO
5MxTsTfQqWDpgI69iOWXuJxPLb01yHoDXLYaXdPNjDnSUS1BLbEW332RAHA34U1HFqQmFTNnRTML
ujKXuljzpuBeEZz+V/1IMMz75OCTY15FAT2CpiMZYJmXl/Vhnby69gHQKm34Pl84UJJj8UKZDsvf
+rM0Ib5rjSYCo9YoEIen5Zozaa22o74CCclBb8nOcvzfTYD69mxCZ5CW/OtbJStEu4SCSgJDUe8f
H/C+1lbXKxONQaTEsSWLBtGYfGP35fBx5a/yoiDJl1x1Raff0jMi61OpqQTY+0mWibXXkcpEPOYc
1kQCfV66kg+7E4jgUiRxdyrSv5xn0MCcsK373ac+Na8SHehtGVGmoEaqWHZBGOI2YSJ1TEI1qRf9
uVhgaKpV3Ff0INfdM2SKpBoIlIU5oUInlI5wlxdSYOlbCijFUNcLQ1m9e903OucaIL9pUrd3I7n2
1p2XR82GAAwCUY7lkcO+M/RaXlpehed5TC/5o8CURGwwngKaGvBZcpULLHtMRUgKxF4uqsnurlS4
ks+Y9XZsHUBK31ZtNxpUbUKPSv9MdyxvlkAVob4v9gNq9uXbikQ4mW0fpV6PwHSTpKALXloKdvdV
1ERUL2p4yl54WSkbc2VaVl8Z/ZDS8VHv2sWZOnwdNpAYF6qRkRaYCBvbwuxv2qH0rzQ6WEiaLIal
bndPG4v+7shvG2S1wERMcSAVWmfKOXksHCMKDPyjRpP0sfDvTTHngIstHE6yr2XYxPPaOCOcOH6f
WPB+Mo2TByt1SuA5fDRbOxfxXybn/zZ+hD3hMUQB6C6j7rDUAq4BcAUzghLj6cXMXR8qV8bpgMDL
UEYZcXrgePyZi+cUfFIWNXlv32XMo9ZuxcVnRVyJPPQ+IOLQcKa2IyvoNXTn2JnGhjvpfAsI6PZI
NMLn80Va+WZ6A37oYBwKk5dz/Gzmstov1wGpYy3+wtRZ0Bn620kk8bivhly/usUKkwRAvgqvdHWp
+MWwoyM3FQtY+kdO4Dso0wAvS4Jk5bXfi4pl3j13Sfgh0dOdk47+4J3mtniT/l6886QrjmuKNt9W
lVi6u4zEjkwv6/cIoBWWTrKnWkamwTBRkn6g0/40FymuUD86BpJRIJieK1tSbrGhC41NSvF+aiGu
iBrb5R/dXQwYDkOG4vGWDSLJ+jwLYVmISjdIeGteMeP+/X4XdrSSIBO/CRNRm9FPOSRLnlR1wGNW
DXZBbOQ7WFRO+ROgzE3+g/M8dsVG+4d8fBXbfqVs7i+xWtgtU6MWjHtYwQcBJFbGCq69oDSxazAk
sCF+tIBUVd1lQ0YaB9c8BZjDJpk+zVu1BQcODeD4kbdRQtoKXQoafBSNpwH7x4t20g95syJ6awU+
S52px8SgTVM3Ne7YbBqtCu453ZYea2pCblTfnE0hVVeCl/Wm1RRd7WrDI4ARE1GbJtArHOpfJkAw
ZOuk5GUZQhmU0efXjHoU03cWlxLfi7kl94z8Xj81T3m6npywY/dvqO9ia0mVeNyFjsOrF95HnrkM
d9c6G8Q4PUuyT5/Zqmpr6khtxEziUMW2SQ4+I+CUL7G0eMRxhVuxOt7w3+W30Couyij5d9CjR9Rc
9iKMZL5G5uomLJfpjy4/MJMAOPhbsnEVGMFvPLTebMOZBWYInAjHDzvxojp8mrGyjadUNAnYc1CH
HI1nE1gIWH8g1X30zvnqmfACIaBveH29Aks6QS6xR4/gGtTTDVvPSBVM1pcabzmfoJDi30eFmzK6
93IOBqj8vlJTeMXp68lgF6CSC6odRxnT8Ml2SYUFP6YDOEthE4kCraMARrv87Pt87eB/vtZILtlA
nrfQlG05W0ARVCp0jB6gnqpfuSabRY43S6ugyMD8YY2/Y3/4iYaTjdYy8GUBlDlD7OBlAQZByIIC
+9XmXVmoJkU1BXy0ljiZNM2lRgmBcaYQe980x5qHc8qvBu3tIusWjfEr62qG/2gNbQtUyTVTBoON
MjTpz70VggNH+K09GAoPmROSjRtbDUzIQRGClo5G8qyliUSgc0+THi0hiVTxwQqxbWpeweEi6aDv
7W3Y21UVrR4RiZMBQizWFlnJJwN27Vz/pZV25KGXEf4pTCXwzgmldiRFihTfJh4nKtt0Gr8wkQc7
XfSLEDpGkyA4SJAEULZQXwbFPCrFASHaSUGPbDbDZQZOtNg5HXYVlXNgdUn8xmVx6QD/T2dym+AB
sLg2PcmJOBiJcfUk5p8Bq10ru1OXfMk2aWMDGO3QkidUMLSO6whLRRr59X5Ffn6JaRYlyFXUQ1YJ
U6Ma7sqeH8TUDPqkX/eHZedfYhxwxq+cmntzIx/+rPLUqquM4d79hEYsRthKHku+ZdPLPWAVRxkh
U9F2CsG8hW+VKpCOd343ywEqcBsEB6h+EcVmdT0sWExFAJyBenqCUtqRJwOVCJfyRR72GLcSL0XA
wi5RNsFTW6nEC1mH3ktvPCI8aSJDbpysMY2WhKYDxOCCbu/r1woM8iZsvMz4dv6Ca+LEs5YfgiUw
x4NnvSgCQhgBu8vTZdrvjnbVNu/Xbi6iTpIBxane1EMbhofWYaGIN7FhX+PkP9gnnVa8ocfWD2zd
jPpVvHmfu0yIG9QuCUUkdPNE9fveS4gHFY9Ww1d9Ujdd457T1qSJGJUWGX6VIkyWy0JLmjRKjyKi
Qj+B7uqZaMd0phek6hrFZ1bsBAYhl/jYNZbETe5ONwGFCXtAAfUzBovCsGqjicnCW+T5mVlVWla/
z5c22tunB6R8BZY9xcoDZCcWDzj9k76QnJGVA8gP5nmwyLpYou0AyxQOnCaBFhH3msm/80jQjRAP
DFfhA2W3pp7MZWk4ImoK3el7xa0Cij/xn5QMjUQpMx3KzDfqqayrXLMDZGLZ72oIaF35SfiE9G8q
5BqZ1O0/rGCXgArXaBygT1uYjhvu6F+16li0uZ5GSRbNQSSdhOuWY1ht/TwUQerwgyPJQIm7zh2u
Klo8ui/muHShrwWqZusG/2TCEUBWfPcdabfzTi0YXbDK1bjqXJanXDZi+NJlbT2/nGt95ezYbDOr
5MPNbLjjJOrTxqN4oMg0ko78fGKwney2y7SwOOVvaJwmChF1aYgvbvyPwoOjCNPnuiWSjsIcA40k
RQNSRc/sbchH3YI6zpqe/IiNonxVTaAMGYGilY7gAwmFwdlkg59YMviDqwx64gXnc5VMHMFyIZ2C
PstmPTJZaBtAUtbKdc8yDzOEkXQp3LTM8jDBjki1chVIXvuHNzmdlWRhtg80X8JLwU3nx58mLgXR
nZ6NmhCM2NX0/IB+EBNvGVYvG74Ju5xA2ljtXTvQIU+dHfhNhVle9x5Ps64KmmV2Pqu/31OKeI7w
2KQ74HbA/+h3a2pBsqEueGaYA/FM9bYwI41GR5Q0Z8s03bLVsuvAOWmnjAT9Jvur6l5SSqhFeyi2
zizSNBrd6/KthVcS0vvKfVJmeSUV+phjkaG4xaNWi2Gc+73kVnHM23WBDbbLrD9e1RPkWCfCWTqp
GMp9kIYSrsi+gNlQ7CIX2O+c63yZJmtHTxtbLTiYzYBazvzTmd5gqnRCy6AFOyX4UBOFbhc+Ft2S
Vj17os8vBXT4CAhrfM4gr7QWcthJ3YqNXfxiB/vJVMhbBWEHRi78U6J/5OOj0TAM6hItOpYYa6am
t9BIg7enkQaaNG3y9/v+ojVzgmAOupaTWvnC79ByNPFoxze5FEf0QwLoivA8xC1sk10JD9WM7pi2
lcC/4rCIOqWFcNKtggRGRPEs0tN1nb+C6gTrtdTk5fW38DiZQSG8dFcuDI/Ehdayh9fI6GRJgaGy
d9JFjrySTi18fjquuYIdPuD5sUHy6GD+n8W6f4h872fMXdEUAbdOnvAnVho+SRjseCLpys4vQKG5
Gr7p/jrhsIHRXmwzXZyOww9By1uqMCfIQQOklZMrkwI9lqMqrnzCWSsLZxKWuS62U0gR7YvYILBp
Mlbacw1OhRa2qotZItOoPLLx0bsGKNdRsc+oE2wpESbOrriVNGTnjlGQnJsYsxcA93Y/NZYOdmH6
RT0rW8XJ4kfb6YRtl1nMzRs4aY+ec9dvwtKmcao1GwfcgDJy1iuZwOTUOMKa7Ed7WroEbd5jWP9M
phhPmeRNiIDzP/pcmDpv68S3R7yc4rfNCQAxjuW0rhpbwY3tdYcDmdP409bqE0L+ShC/4lPgIkcT
RUKWSaOFBTRNsN5Ia8zbf8+nXQ2j5zJ3JAw+D4E9gSvijsQXrFKTxpQW4dLUebnUFkosvwGe3efb
JzyqRvW+HGd3KrLzGEDQaqgFyfwRTkOTWrFpg3YJAVrIVm4A2v4fTfssYzuculaGcqlejaugfSxK
Z/x/rchECEkoeSVYQ9FuBKtKygoi6Z/BxYG3vH5A11ZwhJ8aup/j4ibBNlhV9B1A/glZExMj9X0+
IWqrChXC7OWLZ9VH383wkwV0q0jJ/zMlH/KJKniSg5NpbWKMSpkYDN2tpTZLn+1Qej7zxDPe+O1Q
9fta5TPORga94McqI978U2OaCVL0ViuqrDLC2HrK5Cc8pKWCwJevIzRn6LT2ElfGt5FFsAXEpDfb
GuteRX0+ZLBjB92ii0D3Tim0vkxHNalSpWunmS0A7AHzoOtDra5x9YKFK9fiwZs4DsgfW5NHxGrg
LgImg1KetXyBgDQQ28kkg5MPBZZnL0X5BD78W57cLkMlUJFm33eW0x6nDeAt7r3lJe3f5mYiWzwb
u5xhcvEjoZtUvAqQ3pE6gTvLZ3z31512iIUvVrTbADrkOmR4AQ+nbH/m5QL/YXxuXKNAop4s1B3K
YXAf6AOBZ95uP6atbdzuMCL2nIVEFuFC/d2DHoEjSISxHrmfK2M3NJiRVU3PO4/TcnTJowfvhVd0
js/8ZukzyZFXNDZeP8kLvajmeLWsACQI4ZAR6UAgoeeYfZgMPTtE8aHyqdo2vJOfrE37JTqkYb3F
lglBXRj0s9jJtp8rUlnRtIFfPxkDNkr4WYl48Cm/KzhPUn3AvzBVzCyI7KqEEBtxUW/tFEQV20x2
1i9l9CvemY2E7y96w5SP9rnjudIaGmTKGLuFlxjX+3eygPf6916Jp0HYPDQV0P+CVI3q/BbAr4Q+
WhpL8BJ+BkZUlwRGgZ7hTsj4HyCOL0v5km4DtVm7MxzU2f0o/THUhjynNV1Zjs/EN/AFd2YtjJYj
ZVn+9JWQmMuxG1TeGXzqb2f5QEiikcQEhopZ9ExpxL8GLSuzCdIzpjVwWBleuMFvL9Y6Twtnw36w
S00nOQRiBLiOAiHj46vrw5j4ZxzG0W+Kt6Fg1j4eJY0UGqECG3pOMHPYb7GW2gg/5M3izo7CTcWs
fEkCMwMeA1/oq/i1/Qzo7kXegUR7Pgh2pWhEFTYuMnB2gpHMRAK3c7ufnOFd8PGk7LUYQiTUBPON
w2KePTv5p3nq7FNrWv1pvtmmuFV8/oWiMfVZ9dT+lGAipL+5B954DYW+fV0Z4zVug2Npvu4+Nc+l
x36PxImpNrR/+1MQRrxvD9L+6Zlq/0QCAVuN7BrmZTqNEL1PiG857IVE2lluR/HS/egod5JagINh
DJ04CD9F5kUFsxHQy5VotH4saXmtPCd5R1cm31GJCwZ3ris4hQ7Y3oy0kBWeFRkKCozOEZ4gdp9Q
LEgw07DeFzQvy2NjvTJ2LC9fnQViRADRBl8SfchURJ5EraPJArb0OX9kJ512CBuuvfJtn4CvjW/v
j4zHVCMvkN4WFHECxpib7bQvCoe4km6dY3zwXqRtK1e2fzxd4XByKfNhKNlHv5jPLiTF/9wzZkOc
dwhfDLbYPP74q+EBgq2aySTmlnKi5qJmyUoOj2N+QGzn8B6S//0X1gMo2trr37jaizLCZXiy1CM+
Yw/IMnXiTvWvGqtP/Hr9kXpw9tSCgQjDdNXeJUk6fkWhCwPCmjh/opSLDNoEdq85uro2Pxr61Ttf
uAvWuviE9AySyyZq46qItHJy5ZiK8wj2ZpAJOHmqN6VAjU9RLsjsoDgcmyn4e6xEeFZENWEy6EfW
fZlcmJZsDrGr8r7UGFKDh5fq1S4wbQqnwFgezZeEJ9uiPb92MOyBHj2aMLSw4IbqFFfbCwZsAORu
WphtaWuKHtcSr4yobnPOP5c+jmh9K4DhiQ3vXjdG6HZ93e3URgiyhJs3mWFTJxXqd/72nUQTtCeh
crSmAzYNfVXZXEMJTwDMtpC40TO2HtBNRnFN0GLF7pETK7jlY9+jQSQHDZfRSXhxrfRPIRrmOeko
snC8BD2fklKj3NaXwn3sqr3RWT9HlWvNamRXG2NgDNVpIvNhU0uHZa/Zv6OymIhuJYZeY8ufiv3d
uHb9u221zljePNLs20graQ0C0vskFk6Q9G5iEoyLYqCVWrYRgXWyccqLDnq/X5lc/G+LdKulsK37
LtH7+Rx5uRwU0whzw9iUJcOhzXt1iSmn9KftCko4cJtUB50kxClA6MIEE3YvXCbhw9f3rzq/nE6E
p72V/1z8/Mk06VtGgXjzvYpbZSU7kxu229a7T103YQ7mRnrVh6Zup/VWY4sVd1nc2LckOeJVxvoo
eCM0FSIRUO3IHrIqJUoVh4x7gcHKlVdEhk7Im0/WnBOUR2t5lkDklPgHuyk1b/T6x2kAP4iSx6fM
KtcCYLltonIMXaniVokSZLAvVjl1ZJNGrNQgTX2weIHDDiPrUCWZ/QBwkMXnFIACm/XsqZq0Wzgj
ib+Hd0myOkds6gwEW4e/qVl7H8UN704BTempTxlWFK3eRtCynX7th5SFEYLKa+nmtZFXXu+BfwXc
WxqlEzLZB6ttjPxroyHshu9Dqv+gf5vj8hgiPSn4/NlsT+sKdXXEV9zL61bEj9kgANjfxLHWgW35
agqA3zdouljNM6GTBIAtEoV+l1iCisXv+dLboYxztae90r0CIpxWmNoChT+uCvTR7W/xpYb2o61l
yg3FkotqU5Vce8QIMncoBPBX2tW7bv63fMAcHAK7wdE2GUstK/vuBl+7qw50sa6L3ktZ/xpE6a0Y
8sSrmwiJRjScu+gusvfo4h+8cuDjWmhwD9yHSkxr3T/A5aAcsffJACE/eYNSnhHldAnibhORjhoq
7eg8OR4/CB53y70RSxyiA/K/BwfJojizs/MQkcsAJfOQtprKQsWimtOkqxuNxFHSi26Pq3uyoGNR
gFSBe0p/3E5rzNApthPS8ZnAgXlzbAGWnIdluIs3IFUZDl2CEYsuI7y0QhN8IVmzNG9rbNU/i/4V
C3IDax/05JVkZh2G1oE6+Z2l+YeDVEzzoycdor7PyYmeBKNCxGmqiXac/k6Aikv4/W5S9DqVlu5S
dYvI7x5sz/Jn4ME7+I21TMUh4LqUuO2r+a8T1mwPNbMbZNwMSvyYhArtwL3ZRDDS/RdLjjKn49IS
k4UALqzZItqrboAVZKT4uoUREKeGVH41bRfOE5BlbMdNYF3VKlExcmPKxaMBEYr6+AthPUFC2o6m
bktCOUsYk/2a9dTTyHxJ1dcPjfmLCoBNqIZ0VzKyjYOUOHBFoGvCN7gwWL4K3wGPUS8dkq3i7Ax7
oyxqaETnwSLhDaJwZJ/z1uFrBYaCtptOqG2tDJDskKiA+YJGFaM7A7G5N1L2EQG9Aywr3Ri/zjm2
VmZ9n1m80pMsMjY02VWFExwVX7hWjUyke7LIyBNpi6bZ9bMCfP4dI4NSV4O52o6vNraArei79v6W
rWrQK5toxDqJbagWrRt/ARWgIm/efhq+NlFG9jPxwA21unA6RPNho4S7QngLs2e/hvhYuKfyj59a
Vou0lqKyDptUSnaYoZewzyWb7J83IVW4vDK3u+3UMi6wUI1HMit9nyk9srQ0Zj74yydZnmByI35V
42BjJEmbkogUyBexWLnxrbgOOnb/5EdjkgsFwDxD66HLu3TI3zn1+mJoenqmeFDygHi+fgMMPMvH
At7VTOt6h7uH9B+E2XBxoeicjKcpXA+Fz3mfrMVk9cz7UrBWOm98sy3p6YWofZbayuuG/0YxwL5z
H6hORjNpx7i8eEwk0qXOrpe6RetxeR3yLpA6C0ppc9y/PVXsiwm7vkNiJpC8ZsmKHrg4FhvC6kP4
toD0yiEzVLJBZgDB545EA00VcKc+RihCRy1m8dJIBSvJqlzqZWFIEe/Z1QTBNdr0KGz/833SDLMJ
KIAw0sj3YJemFqdXWsVdDSr1YnnvRdpCSXs/sqzeBbpd1XHjew2znEzRk9zrEy9siGMI/RBW3kcb
ov5cktm8akltlqatF98nAhc8kSuxQRk+HJxn7mxpL8ihrfYTC9jhg27ptlXw3J7ZE12/mCMuupXo
XzXD7ZaVEYRHNcPR3F1yxOMqm71uOHEsYP9YbNyF47I9asCutJfxsBokiGdhvZQQJlMEfS3HTH+5
IutAtZr9RQw5Pr4vbGmeiVb3rAjRFfpuwb+mRlEub5l8RfME1mto1bnUB7nnxZ1w9FA7sFLOjts9
ZDW9KbNfm6kgTFxFn7JcfUhlNCk/FmVbj0bQtClkC+u6E6DB/emp7HquxxtxwzqAlIgJ/nU0yF3y
hoZt6a91gC7/MVT5H0MdVDFyR1pytaZRT7zqfKf32i8YADc6jima2DYY7hlrPpbuFLD7n2SvQAsI
7jRE/L6l3SQEo2glJXhfQspY4+zKsnKSCSrFHZstfjpLDAnZdiUMBpTU7+33c6R8upN+WnCj/lUd
SuHnucN875GBp5NOyqaLbDC13t18S0UTB3CtujfMcmxihtJYUJKiVOPdbNYu+6iPeBMRJlS5lXQ0
R+dlY3FmaMzlszPLvUEP61ytH3jrXIs6QiggFH6+UWdH+qysI6TxfbRmDNdnovGtq1/MaKiGeiGe
lMxKX1FKbgo7YBUO+FF3m4M0HdHay6OMcJmGaeiy8S4DzHUdbQPwA9TnD+pHLQM49GvFI74LO7s3
jKqWH0lS/GlTVV3WhOZhOrPolAIeluRZZz2Zw2EY5Vh3UVB5F+nzuo0M7E6LS937mbUOtuNTDKOX
kedLqmaBeDEhzrFC8WS40sQnD6abQstr4oVHBqf/UM/WwRwS2vEt0QdjChAIGZcSBF3Xmn9xleoT
g8Mpkqsbmdiv6FR8jytc251L9DHAeen0Da8BTX+t4rAVJL55Pun1a+FzRIWRy/aDAQK35aRNb0tQ
d1DE0HG4LF9QH9kphqaeCWHSrqLF2Vv2P9r8ggbuDhxzBk/Oq9AUra5B3doE8aFG3R1PNfwxiN9O
05FZH/e3rShmm7ioRM8ECpcaHJwD09lPw5Pl1UUtK2Vu+aQ28XHBtpu6BuLdYbm+XrIcvpHvDVKl
agq6+lj+AFg6c9r7+RZjxoYQMielcdCQJ0xmvt4ooT9A2rZTkt/Tcow1Qgik4hgxbPE4SpTW2me/
/g/QaWOjYDKkpO+TtSPsVzM0TxZ3GJZAouzrZquXjl9/C1Sgl6EME0aDX8uSf9Tnz3fqNFkw+B5b
B7aRnlhM7TVh7/dhYZU+Rj5xko17qB6/K8tS8qxUxOugPV9Wce1nynA/VOOd7glbgHRCbN1SeccN
wnYgM2GwpT7DjCqHXWBCGqO8S2dDPZkGKG7O/w1IjIccrIpCw6ICTghW+3xMAz84/nGT2kLZELMn
Jd0Iq5SZTdQpWxPXV1rcqepZze8Oso/PCmAtcjTrb713/RegeqEsLEG+t2yWNNdDUxllx5Y3W+j6
AcfA1Px0cC7RsTQneFi4YcCy0BxO7fbv4j52hQ/b96xJO4MHXs0yOb2Wna8k3Cud4J2KpBTbGdp2
ffPC4VblMlwf6EJajaJ14lTZgf0PWEeVmuoQByA8F68wjbs9mCkrENovmMs4henA+dr7LSpl5yzN
rKK5psogCd5m32CG7NmsJ6QSXJGaqSN5VqAuuJsJIJpJbn2M3KuwDE6GypklrdWcq2E5RzDMPCVO
N6Qhq+pFPb5XDtp9sIsJ1WuxVOTEEwaYp85ddcS0cpklvIJQ5UwqLfKbTtIy0Qi1b24I2go5e3kK
75IzJ56Q5stYc01BQYEM4e0w1AUSEPnDv/+xGY/iF+6cqIwWa4CGR7gHUF78QQ4txe6uuTSMYFfg
tgUFR6u0wjvrbRABAPkiYXowX69++YV5p7i7lldsOXPhQWnMd/BCWmBQKcBToW3lq9ZK1jW3ekgH
tbHB09mmnBCt6NwKDu42ksH/7Wo9ruD7YZw5kvsMPDLDug+g4wSFono0dODIMxSgZ3Oh1tuQPP/g
GVfGCaJLgM2k6ETzf8py9A1bsmegjmWIYvRdDpZL9MK3Ln5JHxd+zFQ90kLfX3BY20a57pPXdl+M
PgHGKhu/ApS+kRQCLpvh5nfJ3omuGZpq/n8tQmTVeL5OyWlSYHjbCcIz9N3yy6jOd9ke97/gjdJ5
arQxwm1JPsnQDAteKjKwM8L8sxcNDHPqpr+6jOXWsTxNW3YtM5K6t0pjyFWHAtWc8nqMA91V70I5
xPHbmoL7Fyn731e1ZiPYZqxOaoeqLwZWhJWL82wcxfxawv2e4O6WlguYPKWxG0cWIdXePBpBdhjF
F4Yo0Sl5nwZxTv969J+Z5gNpeElASrnrxkq7ll5N9opLbBuxSz2askJLXsWN1ce/1l8ESojoVlX3
li6xFOtUBgkqhAcGvbt/4p31KgEoG8Mv0/U4EbwOIxDg2Ep+vJjUaZ/grxL+p+5oihbrEQE3HHDS
gk1VjuCaXiS0JrScRbuaWDqNmsNfV8b1PQJkY6zaz+91DVTVxMen+Q/Knkbu7XNZc0KzZG5yxHGo
thjZJ9tCnppnxc7JX+Iqw1l1yCQbHawhu8QlpZmXLDF3Rm9vZO83PggqT1SG6VG5hPhjNs/U9Vgb
XA05qf4s45zDMOHYoeVXnRnArTSX73CSPkb6fav2yWRpdHuSVFOKdGPMS4cSof35X/Qzi1LLjUup
LCDCSib+AQEQzy/RhfsB6Eidu6aydToQmt12McXmt+ihGCYkVWPnQb7lO6xc7LYSrqRAvotKnW2s
pd6co/f3sCnurg+1Gip0Via6GFLkU2SZcEtYJ5ybJ5RjlwqubPj+G50Hk5y0outU7XJuZ8zeowFO
xgIf6D8Exu38X4R8OXWP6cn5PqT4L0/gNmGuWfGPRgou6FuyWcSAsXgU3yf+zapdHhedz02DxkIO
z10RvPIgJP4M5dJxshf/fzwKGEcNHzWteKawAnQTf+ebj33fWy0xO3PaCr4aagryJxGBTQVo5ua3
orlJk+MSEfGkhVeeLVVYqFUuhwdH+WrVQiwGgrCJ9r4Zudev/1kH+YVy4yIvd4XNiOOU44ObCA41
cZoZolL0L6E9aqK5w0ri0eNUprY4ZFUfzaJX3tbiMDIrOOmoOZz2V9PqhlEnoxxEo3uwY4okABEq
bZZTL5RqFodoCTIUh5xtO8GO0ZR2fOH3p3npRxuoycUneHpW3KtMVhxUem3ZA6VPhPwpixoVNVTR
ib3yxz0dbfroaWgAnQqCNiHtBq1oO/50WtTudxUih9mMnM1gXg6g/4Ra/ARhmL71HcOZxXUzDC0p
SJb1X00MlLx/n5k+N1t7NBDn48Yl0B9WJZVNEjzyr7ahsXGl8cGkQh1M3qi2aT0CDkgcU5KC3GI2
aaInSlsNK+VHBpDX1IQspFgrmhBxzrv3PZOCUUGhkNaIVNGbcziqQ3V7sJi2c5hZCtmlPHDdCShr
Gs7tXskEn0Em6iJmiuMRb5VLbg07jzFZ0U942UAf82YgQhkSyqiI6sgZhBy8mZ/QAMh/RMNKmg2y
TseS2Vzw07xnngH/lWNtt/9Gyt2l/uZ+ReQb2GnUWNpq8xWPKSfcCH2Mmq/+E2R3HcmXgUNDEzF+
eVnsiU5i0OM3ijC01KPtdXvjACLfVxoIpH9DT9CZyQnRaor3mdzMZ16UzVWuUz8ssLIswlmRqWRd
XKO+Qrlgr6iWzyn3B5UJ/dyqdKYkBBECPMKhbZOr6TAuJkHB0/cQbaIjtnvp8cIjD5RgoFbWnT54
LrsRBB6tfGy3XBdge0jAmxWANy9dUwhrD1gvH60G2dVGcyfxIxrSou3LQPNzN2q2QXQn6LLsX3uR
Pmnnj2G7zKWFM2ZBFP9pGNNUlSHFIPO8YnTfHCxyUXTAFY9Azr+TLfPlYZTcr1yTfHFrCSVE4rkg
NlBDr3ilo9jP7o0XI3hLYAPNqgxfVXVtPS1wtosm0ZOWkZwOUXMbrZ2EMs2pWxIERXPEg2PW4U3O
aGnPWKkA3H9LJsyMNiwyGp+Uq78tam0ikSuBvVTAWqPu0BMELWRHAsKD6xomp3o5G2B0TKGFhy0v
cTIqF3pvs6y2HBnBgEmgIbF7R1TWOuDkHP9n5VLh4eO0w4B2EgrRzhY6l2w7iTZi/VqW3ZwKKbmL
RDbi1O9i8YhwqCOFfxjRGLI7TTnc9ckK1BgIy586/bvZPGpkiMxB2s6HHP87dxvxTxLwA9u3U0VJ
bXj7U1tRKYzRCXpWANx7hDnL1J5AtS2eOyk7v6CjXj6tqaClNei8IAIKlWfpDHWXgJb9Qj4sxK8d
XFGz8Frl6eAasVB9hHzceWwlryHRk02EFBh2RddDzuLUBw+GBMfx/vSRBxz8ge8kmuqN0bFeqlIJ
m/R7HblkTjsTBqK/2PhHgXeaK1Dlrjr2JKEe3n6zHhovKuQWmy0pND+Hd7LB7QadjutctIm6a6Rp
cXCWAzRK7bgZIH7zIpuemF4ZU541HurS9mY/rDHlpGAj9BFe8KrFyw8IxiR0NWXMskdSUVt/2SuV
VGNwW0+EyQ7F+O6zwSX6Ha1bLfzxTz9ZIwOwiHFRBp8e8S1maBio7bSKv9LfENlX7tAWP6UgSapj
n5STPM2z6Qp2aXUTvMyfQgSPAt07G+8IwbjYQRIjegzE4P5r3UfhRlS5jjMUXSjwE3GtgMkcTrfc
73Z1P+mZrGXpECmjMi5xO4uuCIEMm9Rtp9GJ+rBlmqqsPG4YrDa4p3SLHJclqRYKoRZ86Zs0bF8r
+FPwc/RyJa4SrBcdHjEgFg/XGDzwFxvMRTkuTlpyJ/xGa8dBUiez7hQuDcD1pROQYH3wUPXFXp2J
FO3eGlGetrs3f9T2BWUOh2in9ghVCcWLjmiKvebtsFI+WnmWqseiHqOXmcsx51C8FsuOXWcfEyaP
WG8HlN5aQs4XQZzKH7HBsbjJVUsCnxWNc7UUH7V1DnckD8T12LEseuJLA0kgfBvz+xR3grZYRBOo
6uoTRh4JBm1TTzA0ukOdEasN4vNj7/t04WbwI57sQCf85Pws4jZ2bYlFsNpA5WWEL5sNoqyVZ3UP
njnYm1jakJUTPltcvlErc0kHZtyn/9zpsjC+tBRUbJGdtD6iU8nUkKmcT4cuoAyo6ai6qRdEfAxb
R8rihYEp9vjn7UnChLVGU/zvdTgK87c+A0kS3rw/w75mXuYv2K5Py7QlX/eCmj+pLSGH4ApzznKQ
nxRiR7P6J58LJk7wFqxF3vqg6jHAkYj8P033FufKiB3pCv9IoE1w32Dp2ZOoakh1tTxanQAIsv/e
mieQVn+aEyAof/Vv4Hu1nCkDRfnv0wXg25gS7FMZ61nZX1Fh4hyhrjELKjznFue/qvakKwPHT7DM
3pHlsDQY2SEXkHQHwC0gu3UxcJOC7x03bqbdK7iCwVz9wQ/JPYki2jeyL9JEovXiHqVSJVzyN6ig
CmDFjSzf4oWLY30EKwOanMgi1dtP/SRZVLC8Q+Ed9bOHjDKvEXuwrv94k2ydDCMBCF95NjvO2AB3
jPjxE2EKt0axc78yNTaGyc6SwZggRVXXb918JRzTU+gMvWRHOBRv7V7zz7e+JSpOOpcFjNSL9nLz
B4zklU/D0URkVCDJnfwKrIv8jwmRK7nR9LkhXgIUtKs9Y07OoG0Cehjx+uGHIF6QTkPaMkh4CibQ
mPdn5mwuotTJcJyQ9L/hA8y36LBTJAUx2shLa//tthzrOWmsgyyVZISF6AGySG4VJvmR/m9GkURi
XKYfyHKcjaDAlZOReEmkYMkcPwL50bfQRkU4EeO7WEcG+/29mCO4Nu4jpmYD6zh5H0fXJnjgUyE6
WEvrJhAIEB4dlsnRGRQphCL7mmOMgA5mrBuLhF/zz3+Uhgzz++eBFFDPlDNoIt0cT/sGQx/DcpMj
VkPiB1nIpXTtGA2PIKBU0JTkTfVsB+Ef24jXo7WipT+L1sV9eGMfPYEqIEGvGkjRePvevXjHY3Jc
xAoRLVEb6g==
`protect end_protected
