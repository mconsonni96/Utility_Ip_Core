`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
sosLoB9VQvvtqceJ4J2+Pu0iH2xK7272LddZPhVTC7vjx+Is0r0R2Z6xiq6u3qyCsXa0Iby4alHo
/Z4aznRGirD5hP5TdcjcUlP8HKF+Bsbo9hjN4fN9+4lqhUPjukZRy7Tn/knrmIzK5Uqqka2k9fSn
4LairYw8jT9CtIUZROdEtSxU4Z9YIR/KY2vhCeD/o53u1MUYGNGMPlIioqNNmlKZb7HyD5b7x0CL
PY0ZNOm0xVgwhl8Je6HEiPVN4GHQ2z4l0kSp60ZXyTJ3wx0qVAsWnay8AiwfBlgMM9fxL5QJ4Lzz
kwN0qcy6QLXHb3xYDNPpGBrLx0VS0Tt+ixf8GA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="nosF4qn+aMvwF5YMVc1/S5Q0jNEOw/5GDi/bt3IO39U="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37568)
`protect data_block
YWSoLIudTBp009f2ruVOLEdMmToqt7G3XXX15X6JBNBlKa/Y5kx2AOlNlPfHmgmo0pWEEyMdavbB
1SAOGag/TAkBlLomZx0yohJ8y/rKkzneq/pkEXEFUE2FiWhbPuRXhJgo8LF8R5SQLW7DSsELN2op
YEWcukyNe2L1V9fJrmqHzqAx07n6lkW3wf/T9HEM2nvdTcIs4qJpvcJfZrxmsvEX2i9bKkgp3PSc
OjMxQ92OMRkETKAWqGADhFSHbECRTARNCdg9yUygX3V9cH9JsFH1u6rBtIxVBrA/aSxlEvz39Q0p
Z5KGfpAqgB8aGCgWOCst/JMPNN1pKjfqnbC/dpJyKBDasSh3gLU2AqulpWe7ygA2E/mjySBTJB2l
+y442dDrgTzeezjIhBsl/lmxrcUFzr95szDm1qVdiPzYnbc6f668NaVLoRLJw2j1ue0lvLfxDven
bqwtQTAK25dDmqm33BRaxVAQAaDkG61UxOcH3Ny+pWqbIUyu6dw11+29pXdlwpMR6B1Pg0jVIzPI
yG5CNY5PZTUHAhXVnRRc+d2ZTAUydEEd3jGBuA3rFUUPLe/nJ8jj9IiCS/hKuo1r0Sv+HWZMzq4c
sPXBfZKxc0aIMAU3/B25EXzPsj1ieCgQFMkfZwCqFnnAwm6VdNcSTeA9alaIFeI1vVbDw/o170pZ
hAeSYDLdQZQXlcOTs2eqKEolJox4fba67ArDBGQ9cdYh+OfR7coSY6Gf1ufUsANJcsRpf1Z6WGvx
VHXKgJW3W2878DFxh+DGGkHFELS9wNqyySwtwv/2+5nyFJlP6J4REPgqrZAklK5rnX7E13139g+7
i48904m/1/l7EC8NadLGSm9h/hehyvUoNq7tU7xXRIU5DjhLH7TQL29Yi9/LZaThq2HXdZizzjVH
7ZG02HTB+FX/XC87K8mQRDx6JSDfeC0wWYoJbVDCy00o0TwYuUAxwECwXrfbb3TP/Zc6inf8kEP+
jp3E0h9nb8PmT0LZAbpEVS1hePD+n6ig3NGKAQ+9+T5lD0PzzdrHXN/cZUPrMIIcAO5x+oKmcceK
eux43JKCBEwKW0goI2Hypxk+7hpLTSwLkdmguiSYtfLp8oQtLyluEJ9l21J56oapBv8sQnnyWf+3
O65qt0KVT1DAEusuG/cbqsyFYb7AKKkHAnrGUyDrmcOwirb2m0zqwU7ZGUiZX6YGAbGbY+36VDKB
37fJAbXaI3EICQyFRWFK6s9mNl3uWi31lqUsc3UAU14yg89V5L2S7qihpu/LhZzmI6AHlmcdz8vQ
Uf6lR53KlF9kIEim9PDKpUjK/8HFjyZ4J5TB7tsK2XOpwRhvnRpigr+N3KuuBOI4EXQ8Hye0asNW
dAMlN/jMjkTRbK422hzTk5S/gSzzigXTY16ivPNuLrU/0irMLx1sGZ1SnEwxKT0fcqg6ouYYttTE
TPtfWK7kaLJ1zFLB7tRsJux0PKkVocc9Hzt5O6MgwtB3OtN0s3rVgz3bxjhM6X50brpVyeaeKIxq
lgtPhqu3fciEYuDtVAnDyS8ycFAZIsqBQ8vqai+vSQU8n1KVjtg09SUxPvlxeylpbSKYZO8qLXCg
1E4W+oGtwPp9Rm4OoBYpqwnY+doVuEvp9UO4HrqeFWXq8gEhfi5hjCHp2K7lcUTjlJFuZOxja3JS
+uguoBXKfC/Lly9IxSeiMTd7i872SYu7MdJZLKGyrMP56TZw4Kzg4I0hwBO5nx0Rvff8ufQnOZze
x4tLV6Zl1+1+HGG0NH8/jbgpNF2//dfDP6jYeLW/Gl0rASSvyymVx7yZGQWB/xR3cUoetzHVocFE
eqmACZEUaPI5jLgbJ8W+vLZrRYm8ymLmrtjc3RCCh5uZHLmCztRpDPL4P2YWilEglaJNE6720hI1
2PM7h1YXCeyLu1ac229P7j0TKKuvHANZPKxZfzWNFQLlSkC7vVHStMc3c6XrrBJzp4Sv81+pQWk4
EXC4B5yOdC+6/muA5LY/Nut50z1F7xI4O/Dxu+dgzLajKZHliaUL0MSTnR+IPP6SE56l1tK2GL9f
PC+i16eo7vmTeCZOEORCPV3iRUpbwK7TPjYJQ5JoBkSwpiDtdBo7ATfgcli97HUJLVmQj3Wrg3Ng
fcKu8K5Q4MYjTnus04JqxXlXu3/uxAH25JQDL7QznC77E8XyR50Ym2/kxxmPkIk24/9cPgCPzcXu
TA4xiQvQ3DmxwlyfZr/GfSaQ/7VZfh32UIgHjw5DTe+jnPL8TIU8rDoJXsMO0USJwq1fT53yJJvn
0KFLmqEzLd58TMGQGCLJeRTJQTvMBL64K+POOsy77t6FC+8pmrjyg0uz/eGmkg3teP/t3HLQD6p3
/NOHIcXl3vPrvQa0kkKNvg+db0ZrTUQyfgnqJX0+tA1iTKl037kOZCK6L6mj4FPMREro3w9HZzDJ
+8+jr4tFzeFQDvFX+zIbml9cN7zDe6XWe1q/Y303FVYTp7VgmnPOVkUURRvYQKNg7BeEEWHBDXHp
fICo+q2mwN+fZUy+1i8mfjRtm86Y/kZaqx9+m1Wn7jdMJEiGzdOHMdiL2CtEE1E+uGm4HNvU8DVc
xGasCOij2ZYtvIBFMoi5QgygG4Et1J+RjH4v59utvComxxeEwnFO9WicKcQPrS3ILvY/UlNgSlRb
j7rALr7mDjljeeYQzsMDzgoQwlNYogqKViVNl1uRa1DN4cK4mdd6PF2w1W1CwIlXPmsvSlHb/I+8
fihI+/J1koMjSbzuCOJxGeYkNzHEKXOOwLgL5j2EK3DB1ExIZAwkrSpXXqjM3+YvvWS8rsyAEuBV
XXlhzuAwH1q9bA2hgZGYbXPezeymRdoda3FJy6fm5XB5UlDztcETNNV1BsmiAWu+kyEL+Ai0Lahy
rRR7Wpj9GEppZrFlxpU8QOpwT0UIqYlyvbh7hMZXSvVltm34fTjMy9fCVD2c4nN2WzBFbgHUnzbl
URfVhUw6T1MLHiEHQRzecUWvBYu0OyERAhAwMZuMENad+jNyHGR4TZ0mqdkVXmvJWHNauIbopBN8
AyUo5r48b4UAZ1HYhMUUTTlxtgSWXyOV19cyCFBXNWqi4cTQpXI4aPIs3+2w03yPhCRl01xlQXyN
Gfgs3CgRJU9eSIpTuCpBncFyhks5Vjm6cnesYJ2WHg40pLZFDA+FvVOHgKMu3vQVYb4d5sP7Xfse
YVmv86mdhn90muCxsoMwvQFlrWiAQNyulyz9XowYB4mE+boyO32sEl6vieBIKNZ2Gk2zztgsx3js
Vin0G31gZ/+AAxouSAHIuVB6J5I3ASxMew2KFlo+ZDr7XUHIM51RA0Mt+EMSKpk7yfPf8VSfuIPt
bW5V9MzT/zZWLRe2NVxLI1VUxEQkvDxYajpg1IE2kWMjNcd5p08eWGCWCnrmRVSwkv3rv457RtAs
gIDsgS8xMGe6X1kiQmcMl2qarKDNi3aiqFWARQrDfBFSRrKz2b5rsL21gpbBE4FqKWrTX/nN1evD
jngZWv3MWgTo2sJSstl5KNsrm4qEf2wyzniSNXCnetxgOyNdBKYOQTFcA++kpsyCsJEVJlay9rEj
wctuMZ5weG/twy0bOaJpw8wkb3zIFMK3r1+So6j8M/ArAvD2fp5Z3aCUdXjBZLJ+AV+N6R8Vv8/r
MvsjOyTrQnYxX6EQ5i1LwrjBpMHeSLfUqdHJ4VsvAu7F4CH2utnKU/Vf/Utc59AUNPDgEE5Ta7cg
y06EBD5QANh1yzV1zdL4Wj+29GffGtAXX/qgiJsn3GIqluAUGUbX+x6fGHPdvrxqhtqpOVp24/d8
dgdTO8e4VnwYKht8jQrJ9q6TH94e0wBCN8Rf+ElQyzwBY/Wx/suhTXRqdVrnIneo5yScTV/wyK64
fMwr62yhkva7Cn6FhU8ePFzjydL9Dp4bUae+Q4Oi1AlxY0g5/heMdzogCV/eMrKp1m3qffJdSNvc
IdIcLQkXiAHcJtZBVIjOcyeMFkJavHexeV/QhIp4FtUHt/4szMOWpQnw6cJ58vUOS0qzqLpp4kaL
PKf+5SsTkyELthNF+NZ3FJam8to3n1ptzP1FvHFoSAF1t39b2b8858c5oppQfuLjOwDSWt/KZffh
PiVybvYAWtIi2AeNEmNtV1pJgHjVsjcc4I/Dxxk9H7jnILjhNfowFvc7Z53+UZL0V+SZ+/EXZbJA
rQPFJPA6j5rxRaNDrs+Di6slY00aH6hiOaWOOxnxGaOMuI3oOcDMeZPkdrPV1aiB+QCuIReUdTt5
9FJ0hA2f5Olcwg/0HJRZQiIdcvujDNJmWr5+0dx77WSub2ymw8UlR6WKxg7rqXP9vRjowQUK3nma
w0eVUt6m/L4HPICYfmrej6WVc9sW/p1+BH3OEd/DKKlL8MJBuCeeY9m9Ez5e4abPdXMKgLNKRSIa
2iWuG1EE9dXI9eijzUUIlGXDlYYavs5CLZdvA9d8BPzkqv5B+T0hrIjYkYjoVvw3P2wraTKJgd2V
55K6sYN+eB7R3PI86Dkr2yofFpfHQFs2jIPagnNZLyXl+c8Oo1CA9zLubJPgEvKcFqYXFdajXXRg
kJGoB8vEIsgYiP/scsgFMLP5FnQcnCX8S5a14R1sOBanHLoGHEeRZl1m0c8MJTVzM57QPrP4DP3o
FJeF2IfebhREvLRdC91fIagyPkVgHVlRtj7x4Sgz7/be0/XkHBgXPWjjxSkyrvCldc/VNza10jjY
GIkH5NGpRCXyXCy/A1Z1qKBAfilseoq4ftOnfrIEjCGDLPDy6QqpDlqa2+y7ixtYftr/z0pB88S5
Zc5INf1RA2QeiKW5t3ZpupqgMJpcElwNgeBEtdWE7j0xGDg1yec9Ho7LyJzg0rXv/lk3rPQ2WWel
6oa/bIZbsA8vhJFWRGn8YJJEL+9/QhGeHp/Sgim7oMDMiYgRHhwc6SdLZ4muL3P9POntflVWj6+m
Ust2Fc29b6ACxqq3aY6UiUMGuQuUJwtJQSobSS6C+/O+wi/f8Mn+yvTvCpjIE9/UgQ19dsptSube
sHdd82518+g25ew6Ge2KNn4+q4iLvAOFK45zFprclVnjoFUOrX0mvkwU+c4ob1MBota6n1Qpf7fI
mPrCuVtvFgFp65xAY7HlhMz5lfBswaSfUwG58mjquh4z+SsbmBjDLikGi6+BkZBxJGj8sl3HFHax
mpyw+JlF3/iQh7TPnap1EqqmVZhS1bB4NhsDt5k+y+3wRT0SNssZWxEIbeKr7hmAEi4JIrU2HD83
t/Y8eAwZ4VpkdMCY1k7G7H/DPF5FsQh9052xKS5+ksweYig3pdv06z7md/+yp+Sfy0ro5Gm9I/az
th4vWnkWNvFGiQzURJl3v8xESm9qIMlB1lpe2i9mlPGjbGiNGLy9zeZCYoZ+2k98irKT8pS3gxdH
ww/y4FH9WSJVtLtlztwj/3GFcNONLvNXlYidajH5OGN/Cntgk94O+3k4bNTfDm8gi3uKC/IwkxUy
RW5d0j61GZ4QlmGFeMzg37jrfX38vkPy4ztb0hv906YHhXQNQUdYwPnUDLaoMfVaR8aWXJMM/lae
2D6WVDGXI95jkDxTZhEqD/H5BQgfo311azJM1abnEIj0JgqSnOKsohrC2pzvig3NhmSzTmJ6avBo
FeD03HuhOSj+HRdi3IGY0hTkhOT1QPtKL1rbujAT5XdZcAXoi6qz16ZZTQK8D8PJM/0wWUqexgSr
f1FlsTnZ9fpYNM/GkqxZtnhcQp56dLAKb5Mu8OqaHeXuVgDMKk78aALWym9jmgfR24bqkYescwWV
VM74C6l9p2Rd/5j8lKDO/VqV22FeG5Sarl0qPx6bbWwzqLROVm8Y7qbwu+Q1wo0IM3EvehEGKszf
DeXuvhSGA6VGKDMHulC0hTex2C43WOh+rafRrCJTt8XPEy9KUQSuarMS39NdgUWH9n9EpiJYVA/4
Feb5ne6JRkrGNYXGBK1eCDUmWcGruX5foWsaisppYf8LBOczn5vqWUoWp7huw6vVE/OpDQmmuNTp
EcaRUTn838ogBHxDiiDSGqX11CZDrhd+bRZCqN1zaGAyGgnVfPdwRh7u/47pxfxGelJU/sRUVEt7
5dfAB3z5a9IOdU9Y5wJ1eeeD5QOHVdgTCxdF4aaoHbvVS1MbBVO+XO8Idxl/pVLY9cSNcOpB81VI
VAfefy+UpD9u5Tz0nw5pQPZhxLByn8C3PgQh3a9NL05zWK/Sd3rdGFBGT1+JB+fXCl3XbqXc+8FY
mp0fCDk3zaABDrMCeGJU/4vVdOO2Tsc+LLsM+NNc9Yjrjgb/dVz/vMIyOe2giUZsFj/9AgCIGbjx
B0lJyUKBVmLfJ3EN7n4qM75P51uPqEKyXpQFz93u7f0CkqSzwBCYRDkI0KC0zWQzn8PV3yfvs/Nc
Www17CCPufVZpGMxHpljzt6DPecRWSkUTwkpJefiDHD8hK9r8kHfrqOCVu1qFlG/s9wr+LFE3BY0
HNyVIZQTsLmr1c5jp1TklWpbU3R/SjSVo5TycuIALuPF1yZsGRM5bKwqcHBuEFnrIEl0H0do7BS6
WnsCA9CTD4EvQmP7UQ1IigO3v3w2XrPr9nYh1a6HzzU+KsWvTUQy4YBAgZSazkDDatAQ7iOUGnwl
iXyk/L3S9zSwUTz7xee+jItO7EVQfKS5u+tvfC8JxnYX+YSAVClDC6QBExDAvWpMqmuCyIl1X/fc
N+Zz12bR9Yf+P4Z8WX3KPcK2h5WgIAV+5X0D9Hel6xPmhi7O/zUBrJziDQl/snRfAvNZMYO73Hed
wM1CWUFUaDTanlec9FkaEbSFdolUThfhoFqXmSkBBdENBeLV/Yb7tKlTu4BIc+cfAw77AIZDNfpL
fGOvXkABC1wkiUK7pPiJma06o3XUYV7ogFiVIfNa9Oyr/d3Dqn1HaKJPGTCx1PP3PLSsQuJcEIvS
PWXSn3GzlX0HtHgcvjvA+8kG/nX4OyKjUkUlWRogePQg7jY+/rghnBINFBYXD9O2AiMh+rL8HWE/
VkC24VPsn5IE1Q2Z1SNRBCm90WNSUJ28uq7DgWQJqsmJXF0baV5X4udhRPOQaf91qqCrwS1BIFhZ
wfNLp8KP1tq9Eg/OC53mdpM6N+bLgld1FS4HjMP2GCS+yw84uAoGF0DC/MSJRN22skx8syM61M+k
e3+Ogdf46l2K6KYQqtguE+KdBs9uKks9K53UWpRXI4vp9vB+SVSF/pWSHLhpfKnIuuA/5pFX8ii3
81kIdyEvkuVhTnmfxL+2pV2FkqI9jF7OOzgrhtjtIlkpAGXSO5U4GJTCN8dWwAjUmZVpP2r3CzDJ
UfwyFstShgmq7RorAhgyEG9m7Ss1m7w20kI7Qw1dKi8Y8RLNgclI39nBt+1k/Cs/si3pdnHrf1Ns
QwSiS4AvaqqCTGYS+4Kr/3s8/KdcZmyS3UeVJmM4UVjsG0mKu+kfJ7+E4tcZDldA0JbEqUCcWj8P
kDkL54bhlvb2HhCsASNv1tUCppOh7heqTNf7/v1Eui+X5l4U3hK8Io65oznezJumfKaR3fOdhH1o
QJhFNiis3zNjw+oT//gD/XSU2S8NSE4bsaOj2CICr//xqUuZNDLnR9Dno41CFMXqwqK8CZ2F6bbz
U5QXRGyJOcPeHfsy/cURSSeTOC6lqBfCMQ4ok+jYTYnVQco6ZddUS/tnlCy+OzF1oKDGDPpabGD9
xt+JkOdfeRnSWi59QaZAV653QS090T5uZ9e/omAes87tU2qtALi04fC07D4IoiYQCQNObXV2DZos
7ydvAMXv7k0A0RAi/bypZ2AXLyOKUD15q7pZWB6dFEshfX5cr291jRvp0r4lc16cbCxV4iBOpkov
CcYFYwuxZyqgv2NAFZ6MTCz/N+f9ZPbVAifsfPGTT3Cg3sbfDexrIbrehL4oLrl6J4hxvPSQi17p
sb200eAPlrrtXZP17mLRShDvmpM2q4bs1TYc4gexIo46ugXUMjh0kJSQR9w25yLXyByronUHRub4
Mw2Nu4XhmmSPAvm1HsKdeR8alr7YZKN/JfWaEg29sVkTGzIlwB6O7dp5pah3jPKDbp/Ik3nsgTO5
DoE5uk4i4ZR0tn1rPpMkI5c0OyPhSc4Gu2pDeJ2svaSFaKZKZUCDYnI8BeXwRAXJw62cBR+mV01L
JMOL8xT+jBhkwS3wWntfJAhn0THjXIxYA05NvZt9IeAAdpLsLTXLXh7MnN8LeZmP4UIY0yWPpvke
yKoRXU03OPnh4XheSCuynSqfE51P2dUlOIzmXhIzBODZxI1pn10x58gpKbrjlSy/N74cgXeUP+5Q
NHcnSlMevLa/OQliNLmPh/yW85X++8w9uQGFPHkQVvVPBry9sQi9jQD/9miIp9str88EQyO31Lro
AaNxMasAgJHMyG6vEAXXmam3wL+RZxENvmGQViyvux11MjUNXf3d4TGAmA0bEt82T5ee1Ba8Rnqz
Eo7FkfrJkAjIRAG5S6tAiwB+VA0/L6vS3DoabzsXuBvu8oMkQBWp68PHKHGBPcDFS6PPdt17dcG7
AIjjZ8FRo+Mglkdv2OrLO3qxH/xUXG9EIAvHHlFh8nSzF+X7olkuybChsMC5lOU7S50BmJkq/zc3
jP63BSGhxThJZqMcimA2wYP7fCtRPt36jtyc8IWSwNDnYBdZRVQCrD9P2gYLGH9S6nBQYb6zq2ID
w/auRTSTpsN+UBwSiBpzCTQF0E5Rtesx/Fg9EOZnQYG0L7VK39JnjwtR/VAeHSpBgw7tuBPCW7Ls
lXJ30sZ8/ZLxYGRxWq3RfMYZ9hWTg1E2vPQFp/yA3vFETqXkMrafpiLB5hu0tjKEjsmVcUJy/h39
pu0Zl9Sf/OylTod8yPrfY+Xzk3HDlHXYdkgm7uL/LXgAgmYbF58/8BvTH0gjSRCpiZSXfcdd7w2f
xr0LcOWG7OrdDFglH62foM7ifinV0zI7OMl3rg0hxBEK6hLm8PWcCm/qgP4PuYrb1DGtM/L+ZEgx
sru+ATTvxZ3DMJJVCdvHgyTtEoIjs1EhHBykoWX7+MUH0KMsAWeJsgogVyYZAgmCDn9lG9M1ntuu
OmTgEbbpRkJbtola3vjXKWBpN9mpKZG96JHwc7DtZ2k8dBXYTNApvx5B4P3FIzxEwnuBTNlquX57
6/8W2cF4gvZIlrXkIVUwhn0PDrAU6zId4qBgdTFe/3MKnnPGcyzOqQl5N1LxRTp/RlOyf+n4uqfQ
iPoCp43KTwdF8TYe+Qz8mqeugF+tm4leZC8YlHEW+oSu/65uEMRratIF1dNDHeMzovUArpBRIDoq
tWKvN0bek0mjnSgCufnk8gutAKuPKuoSEgtmg2VVcAUZqDwV50S8dYxblcG6KPWy4ZodaxmotMjS
vqG2vbX3RpBVCwdy4Mm/hbHUt2WLHhEOz5VjTq5PQhraF8acJRwxFNT/mFquPgKudw6FKrd5NlaP
KZAVR9IbdCMcLG9lzAN0P51s28RSQXcTRPDnj4JwsfnX3ww3mVhdCAmkGa+o2FUmbqgWkMMF24OF
hdQ3ofsYnLS2KVXfYOZyET3l5L8S5rtGC8YJFeQoj0zKvwIuuxrKqLGv9tjvBG0ydfxNUnGZ+GrG
yBv3LPhH8XozH+djQtn5OqNaMZTYkW1981Sy/p5P0VRhxnYZ3+kKm+IevPWiy22uQ+MLzNAHf1UE
E19y6S7aGbylgFBLNLbIutX7FfkHv7xG5RZyOSDUpj7/LWa9nQArfyHYuGKyfLjfH7U/YdMWrYAj
l6OALx2/BdP802a6sYAgJ5lF4FkFSUmzZ+8xhOQ0/rVOgZZ4v3HXnx/BR+nIG//eoy26F9NxwArz
334dUCzWloBgOyJeWc5Hg4/57IY2MVhyM8L2PNJmkNOW1h/APOjo82gMENEnztaV2ffOClyYztMU
XFPuI/Df3MGyk5WLQ1E3dnpQrzDojydJMLB2QoQQyMPM9i5CiwJ5mrQ9CXIuKzsvsnHGh4vtl1ih
ymmq+AY+S2vbNVrXxzqatg9lrw3v83izHwrecE+lz+vi3brNJTh1CwRx1Kb9XcqQ6IvuL3Wyb8AG
n6EXu54faj2EzkZlxnajTfhBKvfR9V9uqtSrW9TBLWH6yJGsGM2/Bdst/QYJyjjKXjm0We3ehwkP
IpM/uAzD96/lZu0eTbDBiyePgFux90uSLx8HxM+U6xsf+B7jamUCG2mnYYf+QovFTjoN9HOXhmnl
et5gA/C9avq0hrl50eqTYdv2iASgjvhvlevTE44etAiDfHOpPl8VX29et20TFwBpe6NZmet5dh0N
/PuAe2mq9kcZsJAjljBD54z3AzxkJc9mN4uYA9K/fFCHZHPukon0Y6Sm7x2jr8CPBm+2MNTawjyR
CWOvLnlqa1tO1tVWv4L99DG/j3yRMCPZiE2WJv+ke1jNdW9+FrnloQa1Y0X+kHjlhgy6wTCYb0hh
SS/EKLgMI9Wk9KUTx18M5eJ50F1Gr7UtBLKnaLpit1pkJmAtEYAhj5lQd8bg8rQ4GoUyEWETnsYI
2dXXbBZY1FCaHiQpVYp+SH0Di7YagUYkN1rv/9Fk6a/eT4NH+9kdaIZpnGM8bcPsQWy7UjQFF3X1
shQBgCGEFCNgTmJMd5S1qoCqxf3WyPYMz0/eoj0m4zSCAPwCiPTDwMsnKP+v11vXfvoRgv7cZNOY
gEWdczXms8fotoWACCPEhJJvnhKGf9CoB2W6P7gzjwRDJmSXz/+LT9t1BYXm//fa0RojeCeKPytm
4Bw4pzj5ueJjYi2C1der9sWwTV+vLlUhmfUOuAcKywD2qWqj7upJoVzTp/tPzrjPHiDuLmitTN5S
iu7ok5ZxHLihhQOE6LXQJixa/RHruuTxGFtv5rRm2LiE8l55paUnILxXctr5Ztpcj57JheOVkmG/
MxjuyVsMsC7Q8EHW13tOHhLSriH6TiMpHiKVvaG902xqz7P2ba1Sbe6WBN/rszhWSB1eQAqeDrCZ
LnAxryuB/9FoHYM1tdebcO3MgW/tmdtBVqUM6Bj83/SnNmpzFBoujNbA5JnMeVlbbX6NjsOW7TPG
eb259B6cdX69ActhHTv2DpsLk/B4+0puCSxrxsylIB4T30ryOByyf+VLnjTEU+1x96fej486Pr1o
XJR220vezDSxZD7gI2EpLB960vDaaqIge4W3gmxu1BSfVNHKPkEskiO1vSD4SzMs4tw32UFHmK1e
2c5FAe+1sVL8T+O1KayXs4sTSoeMJopZKkOyvBwU12JZCu6ouEcuGhk0oD3rnF5cqg2ozBn1+s7U
yJBt1erp+5BChWFMs2sRjbC1Wham/aD4l7ZewWfyDKql99IxfqXo+6BqziZ1X4HST9U17Sfqtlx+
hGKAIQXjuX95036qxWadoB3ITKwasKC5JBatsBMA4lU+DlNTLRpjDiH5Psuut0FYTYRK/xhcZ9O+
3gI+V0BnrCHi1DLVzWghVxv1+fnDOveMwpn5E6LtyH5u7otFYSFOfWCFKsW0uiFv17s8tl4QNUKc
HDin7jZ25ldNeJXmVOfdHpkEd6e64kCcyJkB/DBpnR/Y6fwKyBLy5EsAlyD+DMwHTZyqo8RBq7Nl
dV+dS8Q4VDUdeiz3SGtOjk5uANYu+QAdjk5CwJi++t+pzX8Aqb2G1QQgPSgPDUtwHRpGO+bAUkGI
tgohOX0ZdHOFwe9c6WqCjkRNQzg186xA9D+3TpICn9DAX7IyoBr8RsGXusCbVaM6BjqYMKTv6ogf
zDCva8x9VUziPvPHSNr/UmrpNnD62PnbYoANy6vOZJEROIYG8jT3WJczuqzG7Qm6miGPrKZ8ZbGv
/S0YuG3Nkt4sS93h1gdSbg1ohCWp5xCc/rb5vUiN7e1nF6Z9kA/U4zYSs2NikUj9IlOBDpKJlLcG
mPpsRuw04DyG/7dvRG+d2YiBZuPHzXB8Bry5cGM4yFGhP8AQYfypxUlpnFwyTYwV54RvO8HRjVJz
QC2yfkYv+1I4QfsJGBkz00Jd56YkOdiMjEB22Y/4zmQC+nAQvy9DaSRYlx7Vg+qtNlH9a+RypCpX
r3e9ScMex5kcZj9sbPunQMxDriXgGyztiGeoiPICGJEWlqCbJrZX8xvarUBfGxHlbr584GdS2iM1
hF6OAaOieGbNhEelNlQeM3yqDR25Eos+dkFR7mpq49mGNQeZj3Vt2w1Z+oy+4XkE8nbcIFtJF1OK
C132uKeV1VDtZvfoQ0f/Dd7kSGKRZjKpCYbq238wx37LyXs+VS5URCDnGQCxpDmL67tfkzneBOlv
yk4Ke9bvlLTOqrme6DEJDDiSK8o3AeLvXS0cFXcv7t2TDFco4moTdWtWyuRLOgvpS4wR350iRnTe
esDfUp8anPSskld11Ea2mdnOl9/WgrjkOsBWcRuZtvJDvXInN0AJUdoKkmSw7e4mz1TMgpNMX9Th
xI7Z3hOOCRbNaXd1rJ2MOo14I3Yu8/eSQqP3uSbvHATjXyDo5R3uOW809uOM2uJmiryBNODEVyYt
jelKonll2xusrYy870UZXf5w7WT4vZBTsajVtFTcXAj8bqOMfYTDxoEUUgGNoLvJxgGGg1oo5bSW
8sKyfBx7qhqrDv/i6J9bDCiajG9+c6K67psDEx3Lu1WdhEVY7rZRzCrJVZugZBc9vN6RKt+/+han
ywzwL8j9e3zxxBAggfN240flO+acb5RusbTuay9C/7ggVh2jwZPAnMq9PVXAMuA3M3dST6kHbgSD
mAbZXwOWrAzBPqRsn3Cse9ElJBVeZLuR1YO/mty7/wNY6cyied4xBbhTPzN7y/mqpIVeys+IGClG
EYYw03OIFdFAadH4QJ2eZBwU4iZfvVtu2ONKdrwLs93xiI4JmyJYTIcobXehllaD9e/AqPlI8zg3
FhYMlPVGuaIuWRW4ddSHCFfVAsTGC0edlQX69rOqNBldnF0hn2Rt6B8V+Fgsum08hgK0ETLTnY5e
DfQrEjzS9NxMa3DcLF8SHbgWbWKd3pad51oP/8gMFLC81M9Y0m+D3uYDnlaSskJktw7lOD1sKSvc
Qtol6IrpF8ehvmsSPDUSUOTO6aIbavo9S2VU+Fe8XGTvOB3ugF0Rn2Gbk3Osl4tzwEKdt1tIDRYS
Y2DdydtCrsvjfrLEmvaftkx52sA2+BpkR8v8tUD7tuXL0pZdsxSlHQ2Z7eWVeB2lE9AxHlLEGWKb
/BG6vP17EiEvHW3/B++BlTSb4E6aoFNdjI9/SNoGXi9dXWWNGsdqCCbFYsFqb0GoRLa6Q14N/bXv
B1dyalxiEkZnpRs4xsqckPuUQd2B0nl1d0N2z3oEqtfjEuka5vVVt67pakxuYDb/K7tvpLvLU/dY
JebARiBJwXc8eLsN1O7bXaNSYXmvnq6jB8IMakdzL5gYiy7tnl/wozQvCmzy1x4FDaLlh0xwor6o
gYdsPowUUBDgD+NME1Llr06g8ogafoQ7aSuIwdNkcnProKtDhYd0H/gqp8x9PicXpEySuvhVK/nq
PAVQKrPCe6YMoCAlsSS6nyOXAmG9+Uai1bij9AOAhpPIjoK1FzPC5sQ75AZ/erTLFXmaMKmHrcZw
jDpPwlWSASQCSwodpi2svWd1eO7Ymnfyr72VHWiIla7bfXYc4Oc15VGejbuRTDBJLKdQcIFZT7LB
qf1PWm0Ela7Pygf7O7LX4ZqPYNLKlFcdALz3RpQzlWhxOvOl3GsMihNdaUqXAUAdZPeQZfrvX700
RyNuhv6TsgNkH+1An6NdFaaSyQ6DTstWtwYrU2q58JbKpNQudrp8DQTAobmf7zsr6V/SQ8rQmGbC
OYb1nWBvUSJfxpO8sBTEaoqFtDbFfKUcXTnSusm9gtXWxvZNw2U+idHe8SICJaA7UlCa5r4Fz1VU
T/eIRjSRN2sU8qoN9m0efvwGCwF6Ca5TXMICaQhBhGksNtNfPSrkRYHmaQVaQiy1M2ZLJCPCLEck
CumY/zt65HHXwHUVMR/sr3Em4526NthkaXx6nfJhE5ySynSDQ4tLxKA2WX0t0XsTmCmXqCMQBoG/
Pz+65sgnaWdaKmUYUiK0TJGAUmWOFeaVfMMCWVRLHTohS5LkQ/qJBCE7/XvZYZm4x3Utp6/Pkx7g
Yub+o9JBQL6iHwAnyR5X4qMicuphdyF626/gdkjoWka5cs2H5AjCekY4ocoUrR1YnHmBgjesBcWt
/U+rsgb3vc6AdSWSxxrFqlNXaO5DGJUqKPuE6UTS3V6Ivs4a8RUYSpEufXlzGGZ2CiqJPV1yQulc
qbIGzLSUVpnJVYa0XonnifYK1HrpFds/o6ZZi9hchRQvVEgp0QeWUtvyNEUaKsrAnXTFU/bg9pDz
dU6cAL8Fxyb5jfL/yfkwr1HAK4v1oE5i55et9pmHNAq+Nd0tzJMES62fB1a0PCV4YE9EI6lEKeeR
hkDqla1vNvkbqxzfzeXCvn6e71VqUoPz7ikR8xX0JKe8IzXhP9JpLdBOlX4eYeOR1ui349tEU18z
YMrdLb/cHr/MHki+V9/cCck7YTcq8eSORG1YSn0hWmXlUWM5zloLRWtER9+MHGy0g7ypp5CC1fa2
mseBYaV91d2UJta1i7mYyR3OAM01TZQzHeqb5Z5zyw1w7mDnUaboqH9tQGxLedPsuHtIyZPYO6SD
JU4ncOcmBPMKu2BDVkguDxtPbOsg8zZ7PcoBKh5H/K0CvfdcluZZdGtrGNw/NXxW2TNUV9L6yI29
VdI/90Kwk2r0b4y7RZuYjwjxod+X2wjxO4w8epko/Vv2dvSfHRbM69s7ijjROmHSokOC8gs9K2gy
1T5Xxh04KyN8NqAyXvbl5go9akFTx9dwpXrv8l90PM7PFpQrAaDoYiOvNWcvjiHduMrqHkFk7Lse
1IQkLPYnml//mHAhrxFjFQFLbaiIggZ49lW1cfRNsre7nMGlrwF6FpJQXkofZ7qElekwK61x6f2l
iUmfxdfq4zDQXgOx7eaomuvA7fSv/3acvubASbLISz2TCAnEsxZ0StXsETN+Mkl/ZQSQ+D9sjJO8
EYrP4LAwmKEla6xeWM3fQhu/oDw6Wib2awUK6/0m7/4/1j0NTA0ZQiUlnNfLYV50jQcgX43wINYw
9nm7unHXWMfq+7RKOkcT20HRs6sevaTI87GEGf42fwhBQDIA71Imjko3h/IcJM7kVdq2KXiXQveL
1Nx3HwDx2TQs7b8iaIzbRXUZj17cllyW8z/dc90GnwU10ABfInxA5Ysbvbxwe25VZ+ic3jGybwVJ
oa6iYvweq/1WbCetldiyDDICDCoX7EDLWv+K7fWkSobf5vQiF82R93ej1Das0fbZZCNk4qkEb7Qr
JfLjIeTe91N1WDBkvS/UmeWK4VWjMJeMPN2RnQD4HrqmnlvyIJBzI+U83pBDD7QT+zn/OMLOPxeH
yIKtRV2gfpXsCADVCJI0d+isoKP16F5ytUW+X99YZS3erVK8IXnzRFPVGOvSJLdrJrvbp644H3x2
pekXo2ZzZt9jnpsR+uDnKFDr4y7SKSk46cKqybs6/WfQS0sNBgxSkQUpevh3OR6VspA1basYwWCF
7bUDMvbpObdQ4HXb05MOe1gchByrnicGq9OWWYEmJgX7Dh+zYDI33J29lRXHymt0197kvO++PiFy
lXpKfjP238GTeAc88rCputME6piLAHO2tK/KxXFhujhATOP7YBfI4QIwyGzMCiseNEAyFmR8K8nR
xby0+xb/ZsMYAu4xI4GZuhUmhvR2J6YswqyeNIqHTDSvpttCcDQkAJRI7mP3WwmqlTiMJnnWYWrr
eryU06HjnEqMKcmeBd1KtX5u2Um4KQgxSOT8TMJ2tc3CH16kBIZiTistq+hW10Mm1OhJr42JvzYc
SJivM2yleji2bNvq9SBjS2Wypl+q2JzHz3a5LNo5wd4w8us57xQ4t/fnwCLRn0EGnqq+F5o3FNTQ
AqJH3EUZOG6CylzMfiDBQZBEDABXRpC7XqsQwwO43b9PxUoQGXmVZD5jht8+W6YRSLZUPcFTt98o
v77CGuu/L9F13psDg7i1Y0a7IM15TdscFPLHi2CFqdK1cT0c8wf58WcMBwzWIYzBSRMcScUtRHL6
F1Tkgw+TcnCvfMghp0ygcXeyPopIglGItv16P1A/Kn8GqTRUwINra/e+NjAqjfp8uemFrKfVOvYa
MCbrPA2Sk1YRGKHBwi4obDM65sC5KHpzdtD1vu+C9iAWcfeYZXizaMFyaxJG+xKMeLyPd/PzqBbU
N6cDwFp4nwWdwIcJ8J3/Ro0XCg1p4fTXT68ToOfqzn/OQk07MyUSuGBQIyFPuS0ehmiaV702MPRL
6gYghacMafdK96zVb7jizCDc9EY3zcaY2lssg08/QRrzm8vHUVUoLpVfmWvRFVVmLLSd04fiYFdS
iiDZeaTegmlq3IFdWyfQNBa+c8cAZjM07x9QgICLSRi+dJC0ruKZIIDbU8RFge309Kye09+HMQoM
m0XbEzIf3tnm0vAnu0ArR/YUJZIPv1n+wsFGgQCa+LQPUF1WGmx6MJEU5M4ZE294FY1fepiEsBlP
2kNCUsncmAcB1YxigvhAgMRhQCZi5rpuQ4FRw2cssLo8bjlM9scbtuFLPOKwWjQDVdbHOsV7jR6q
MGQlNiaYSaIPzGX2G24p0qlZu9I1xAmvDtv2ktCDmElTyjRl7PcZkf0emAOcEpCKPA+SAwDyfYpV
uyv8gllHVWcfH09Pp1LxTnnP7ELdRzeCsN3GUCtkDYBsI7gTNvvcaiLrxgfsjhEu7DOSGPGgW+Vb
+n3CT0u0O/7YXkmJ6WD8yOa3u3imbLVWj+AJ7XZJkrNnsO6PVVHvqKiKge6WvHUbX9Ftcy1kkIHk
o2bJ6ewdbF0F+n6RQb4vkGmpze24sMy4GtJdY2a9L2ucHcroVo2IdhjB9zLeghN/W/4s0lpUXhNG
DiNgTvNti3+LH9pRtrME7dAJbXF7Pb/CQ9yt0GsCv07aoCuw37jTG/gOUqW9GPoiwGOlbkJos1i5
zYQHJVu84YfpKHkCkJVcAbljTonE2dNGKVZgUkKO4XZ/GXXdEWGVCznglT9WIbaovDkAhPaUbJ3I
dvN5Pcga0sJn10iz7iJt1Lv3x6SdIl79N8p9EM0YuBuPPj8LUcv4tUY2KWWlaYUHZTMyTjMvfzdd
wWQH9A1X6q1px5QYHhEbfNwsFPt2ANh1cz5K6I7GqPE9QCo2e+yW16y1d7Sa+oxHJ/ww0bWtOEEu
brkxkF6PIPUHRM8+sNCboD2Fc6bqkBSOTBNI1EgVz3JUuug57oxGLUlqURfbq+sKLoMItWQMa/oc
ei7HkMZscJNZbc1KJ1J7RJAEepDTuC+TxcuSRiSfdYIj9mPg/y8EAgEo8p176o0S9hkAqOb07ia9
kSC4OqQVv1rUMAi1D+8JvvoAMVYV8kc4kByKw6gY3DPn366cbnPR3VHpHi7wRlwJM6owyPobWOz7
D6k0H0mqnCNDyGQGKuohQXBek/zCA5QX7WunpN4GRIQprAbWlPdP6CF58uCCGRtgrrTR29rOQwcL
Xl9zlYbEt73YxArYAjVbqmGykbTAvZPMT6qtpHZ/7XQ0HYLn6Qa16iakGBBPhPQbXzyjzYMH2OqY
MlsiMbR0zN/dPJYowC+YAXzQ9VRBH+hS4k2u00wzyBuTWDncg5ypldScBv0r7cglYJOkZHKzJ+96
dXOGWTpI1zX3cZN8xaKKqrCKnAP2E8t56CrqSkAHf2hZHaNYaEVcXreBefk0nj1xTinGYLTmyawi
hsJdLapOZ+1HSlydZL/r1z18bRu23RJyJVZC63q0h514/c7p1cwWLyVy22twbNisWIbkIU0l/Pb6
uwVd/9uUU0uKncc/QEvXf6TML2e9WAkmI7xttnSAXv9WXXCc0iOkisE+6FPgvWVSg/c0/U6ZFDEz
ASmdkf4IirotUF/AvcODWjNqi8GTHm9jTpREUFObXFJPMGhxCIHY71BgCJjXUgffBZ4UTxLoc5W1
ERz3mxOlWcqK61aWE4Bh6Pg+3TTwNgZyLTnUXqEAbh3+wifp+/s0Lb/CqU//aHjaQAH52cQ0f7nF
F/VKgrJzmWgJOphen7rRK+DTvwjiZECAB0Bset+bl1rSESkWKQy+a0O3VI5P/YZCzg5Gp/eKjEU/
2kmFBSX159f7rczxEEIUbiCqhO2wmS9Np8u5aeuD7Tm7SCxE7qfcctRTwOE9vycNCF3c5XfqaaoM
r11OPj/WHZagnmnqG5oR+BXdFZovWst0cjLJ4focmTtfoPKOnDTl81hvBNmGSgR2jiY4ssUTsE0A
ZOLWKJezxhzx37VPCGYn2ieVABEObCLDmlJsRWFgi6HpLlT0pSP/GQGHDAQ1pZ0s/WO0/wiQASCX
84BnyGIbmEjf3XEq5dHYUnH+GM+QNSjIUodQP0+WJpZmxLoTjT15XAlPVO4tQ1T0l3LIch4GClaQ
aYCwWVAZCuBNgR0vG60ZEOm8ZsOcyLw4EUyT+kh2tGeBodc7ktKkLrwVS5ogsrNM0omnt1+ccMJe
7/jrtFolH27Ln23I/O2+xr1s2hYDoo6cICMbTq9nJB6hPXV4lNjyNscsX51KC/dzVI7MhEtGEiK4
UqycAhii59HB4g1ByWbt0lP6hS9YrK89Iq+1wI34feNe7HNHHFEfq42f6nHCPzqmjvsrlNyrAQTT
9P4QmUBPN4vwov/KZVjyqxAIXjc0FQefJuaPyF0j7+DPHSlqZFmB2erv47d9YEjGEDrZR/j/u1GX
gXrWSj8c/S1LC9VcOhcuF/TVYjRIymTVdyCGmAhGM5ZvFrAhksJWLgh0yV/oAIUaXQYONjLVpWr/
sq826CIpiz3ZJafV6MjIRI0jznFVVuKLc94vRmxObCyAcVflgkGqjzz06qq90riC5/GYv5iAS8wL
235HjFlhSiKUZQCq0NReXz5Y/dSR3lR7bsgdGvemRhaAn26Ksx+DxzvLt8hV6O6b22TgvtReT9BI
wS3zdKzrHkTOxEmAWaUd65ndu/6p1/jLW98TKqRgFWK/31VZScXWRTyU1Q4Qcjavzbu/fijMordW
YQNr9H8rJimWkqod87eaYjUx0YpH5vL0QCMDqJIwokgkEvn1jVi5pPiStQbarXuJpGjL81U4FeHM
o6/ZBrxpDtl+v4VP/bxVjzd+BCnmxaQK9+FTppE2eC7lEQqCe/T25gI7SUC6KD/3HQ9ubFk5bNVt
nl3wY4nfIK/wiuvqEkbnJcK64/4chI6RdahXD0+zprx4W9Oble/u/jRCBgDYtEGkZmnkFtBiNJqC
B933GgvO5kWWCFu3Bsp3tBdD1CWKF0sabRDp+H7Zy9A+SXHXgEXTdww4Sot+AswwfmU4JMFnppYO
nJpKPfMddWNhCxZ7jmSEDlXD6XvSabvifWgAzIE7d8lRHXIU2++bmEftCJCOaMycTT1FutZuiSCM
oJLCM7UN/ZNwfPvKWLVDyftNF01d7L/yglLAKXltvcUfijjYU0ESgVCI+w9DurrwBo9nN8EZ1R3V
XgrSZ633qaWuOlWzPj953rbT4w48y5AU+k/H516YygaaBgF/8pTTOLvZz8kj65ct8Vyn95soFJRt
tcpBdgioAdQO8dWO9UFxYXluCzb2RrHFDyFRW4wjfWi/4FvO0nTU8FxoyNoxLYktxFQKcviwrsFy
fIqhy2ymEpDI4rnlyi4qUEhiBxo2W0TO8wi42wdgwLrp8RTYYApQMqCZyGK50BzkZ5GB8PCejOfg
2xAt+Brn+qVw9SYBKa6VLiEXz4GnJ4nHiHWoAdUMuwvTGyai0JOe+/rG5U0QKrRjJmxNXYEniDcs
RM/xtV6/8fSnhwrbYsikjVytWCDcwHa8dkzkjFuW+mfUU3ICJWftZDaEM0V4PVF/DZwHi4JkJVar
0UebYSdpG27xMPtpViMXmCEHofh4P+52GMR0mO8gy8d0JOTwQmrWJGvtq16vCAcTABKJOPeMj0Dt
wH9NKjvdSpEPrZ2TvHr+5vhwE7EykERXnyYDf/DQGJwIBcKUXo+PZiK9RSr/P7KBKhAOFbB4Klp+
MEk+JqSGU5a7+IKtJOqzXksg04Yo5tkJ1xVhA4CPRJZ1DZi7srK24Z53jTPBFhFQfXesdCiEj1t/
Z/j454jMwuK06E+/sOfadpIyCPxUysKC5qvc0IHq+Y5mz/kaQfjCnjLlYg+A3OYpL2nxw5pO/Kj1
Cuj1+boacSz/BT8D8TLbo/OWVgDHAcjdoYpjGI/Bu+TIXlnNZB20hYv/KniK+bYpktbHJWYlaFEY
DkpYQ+MxKmpj0P0r/UBdgjdlOcSqAwS+rXWVmkWnBFfb8OjTkhb7AtgqN3AQXesYjBIP5hEV7I2r
JI+oM6F//srTxZrmE+qMKCyQW+wSj/WLXSUJkFmaiMwu8JLVWJd5fkviIGr9Mp1G9WVKqsuyP0ii
sxsBV578FeFn1VW8Ne3eY05NRg+BxhQrTsezxs5H2UAgIhl5ToXB3sLlgbqdrmLHJyfcybjHOCa2
JuzgGd+9MpRniUV/6eRIpHr9VHtpxM3jgjYV/FgSyooV1eXshYQ1wEPMPmdXPMup/k4IPxxg9waY
uWsxQzx1FJIruFs8Ky+kL9yiuWSmmUDtwoYMUqN0y7l5gDLpdT6I3FCrYvvCOx+e7gkAE9CnVaoY
7AEKS1TEgQH8yNEwL6YZ6rcdXNLBUcIA0acPUpx3t4PXWgFe/mOZXHbhETVCvJxuofoxDAnkN1yb
eZRULojA7ztA+CBDRK1IkK6DCp5T3PyKieI31KtyKlm52gMI2OAPojpE+bn/TIHHEwFnYP200PsW
SInvRyLcgG50ebce+YE3oF32gD0xU+I17lA6cIqI/4OGQZ0uN0sAeN+rF5g2kly3lMoBJ9/c30h+
Y6NhlG0MkjKcq+dU7jMt43n2STtbBz5DLL+75vXYjxL6oqKh/1kvHksJXwJDF08xyDjM3NqM+xsl
c2FoYrAaFZHl+pjevsgajGYDmeKK+kL1OyNVkpOaL7zipksYFUuk1Vlp+5KoTvnrXfLkot9aqJds
g3xqcKebF3zs5vFIvdgrKA6WS+G5UJVxRRhORigi/0OPXLfm6xW3xfvc+0Z5mTlqczKPTzNFTpb6
LCiiefcmh1yWdk2QG63NlQMCzemX9Ygk7JQEn0KnESWwZJGbu/GruRbzRKrWBeTuGBZxjifAKZ2J
bkN+N+0ZIfLcoPfj+hhTjTQs4507wPuW8WLmmEQUgSwY+Fcvqs51KQ7K2lpTGjmlE01n6UhBYP/D
OHpygywPLmSh+HTTDIyl2S9ojhd/2JC2q+lqb8+izko7f2F3mqQPpefjUGqlNkfYQYYDSq8yfYYT
BRmq/KraRoZx9PU4fKXM24LZj9AruTlDMQHQiCFEIFSFFM7Lix9nRKizVSQU0ZjJmOrKBclqnLDc
WLOrB1/qJuaP3RoOCH45jREn0mJqQTyvljLhwXbU/PNnNddqV5g1u7lnoGb9xIfuFujCCisKXsy6
teciFYK5cH+3GfT6eRdWvRrDq5s4uLN9DumUAocgdEVRZrErtiaCN17F2xS9AUIXiXsCVr+BCrGK
XfkPrjDT7vb18se+2Ui/I5yPS2EDBY2JJDj2nLL0FSFtKqZ9DPbSFwhYTlDU8ixTvnzs85a9BXga
GO+aFGlAbH9KOaIGl1DJfyo2rxTUMbkkyPsw6ZHD57rkmar7fFvcG4ov+eL1WMGKk4t+NDJJl8a+
nZwGyqyHP7YBOoUUfMavhP9ZalErdiia/rwL3Rok7ryTnzU1w97LoaVomBi8Miud03TQ/g09Rknr
WBoRP11/VgqfmWTw6h8q7Wh1hndO7dZ2jlMQUQQMkp1PBe+vrxC5lCMbYoQnt5SAfbPfrnWQzKoS
GQ/ejg900Xi/T3IhGf2z6Xak1uBs4p/bs7hs/pB/bw+WP3q22iI3j7w4gPQPSOP8n5dKY8CWFs6Z
oqpXlJP1QA7YmLdr1lGFKD1uQ/Rfuhq0jZyutV9fukcZx7WjFhmjHQmP545UkL76TTDd1F/xuCdP
uSmTHqrFJ5IkgrxG4Gqs4jgfKydoFqlQciVx0qo6YFmZI2/ekleO48BFtia1rUOLZeRK8wUEzLPr
fGjd0muAcZp8xy3FFSOfAKjg8Q14TnFp0XDEzA4JCJ/4ZMMfNrS0cOUKkhhDBOMaElqh2dZJZo3O
36qYKXwaK/sGd5ob4SLyT8MvjWPa1b/s08r2Xe6Y4N1aU+Om6kro2DJPtDZTg9wKvxZQe6eZ/ys+
OqEJsMzaNm8NECcoTIWjqGbbpnus/iUbgd8GP5KW/uq6IkaKqt2LYJRzh+/ytE8c4dYyNOIE8bDv
3NP7W3gR0agPAViYxFD8aqXGaJPLb3gNLgJm7/thXVG2GDyAV2tL1JTU+/fKulQ41R2hh++BeifS
BWPGXRthEi1kYtuekdy6Hlcrr1FQ3MT8z5PvDM9nU3nf/bamznKbArT3Ow7GsJ5fPWlD1av4BliU
+F90oWyc3Ssea0G0wa9raiGBI4OdHqdKlsHebU0x/AcAAWCDPm6Atc2AhKlO5uc4UPnn9t/U2sDs
+rukaJUZ6QMvQCbMid1XDL5870bp26kM3/bvwQmyAjbs/3y0KSTWc6F/x7/UZFRae3IQz5gQLF/H
yNZP5wA7Oq1+K+3WkG562DmMuxbxsZMNH14skv/Nmxev8nFxnJXMy6wlF524MSHCG8qrp09pSwK6
aTazh2CUR+dxUr4AqOzWQMrvFtUXXa0qoGIZrnA+0gMTpe/HMBATDuqt9z+WQWU2oPzNinnwe+Ez
B+Tsa3LtqW4hw/p4ExkduIME6m7FaNmnVTAId83TORngErLzO/KiM685jd85xf0I/F/YOAihvN9V
5XQLDm228cqsJFS9dFU6N74oNQMqKVRpDzdHOr8LCvSvGsVM8aFfpNWcLisTuJJB9j2l6Fp9gpqD
x5DN+BzVc0t9uogiu2o+rGcrjEX4PHsJmnYw/lpisIjZEZPHxJBLuueazFsYR2rWVW3/CVGhk9f9
9lu0uvNGI7FhmVb2XYJPsJQ5tAkTjhg2gaMeggiUb6uDM/9lJ5L7QqRE13XdoSgfZFHA9cJm3L8j
rRh6blophiCDX2eMl2Z5+Vo1K6DvIeBJmSn0DVivpcqLb+2+4f+I4xU/qSIZt19mNituoV7rR1PH
+hPV9/p4tRj4eGqV4Eu1URIcxZcYKyuhu7lkrpqB4RsFEaZDL5tD8/0MtiVmqL25qCBxgGew2Pju
8RdTr5aMvzJv9wrmYDj342fC5ZefmYAn3veW7f73R6jYwclmrvz5Xh+0UqxiQsHQgv4P3UAnWl3D
c2gcymMwLUjYldPL69mETTqdOq0WhFDuR5QcLrbhydZ9cPuNZjLOBBYoI2pzpJszf/elhbQhMJrJ
Q3zVacU/kPH3dtZF7UIk8Rcuh+uAj6jJstW8PC7omgktf+0tmtM1FXXqw1qqQd3Cd76kPnD3bSH/
QgHqmKYni7E9I824ICIg3wsyTRr+XqGDvxoa9WnunzM/uFUtDny04QgS57/NvDWOdcg6mxIL8TTp
kMnK9nG5GsEmyFWysobsQRqK5jnY21BfGaQ7a1j6VXGu0SenYf71Bfl+usGbXS0LmozI9W9pn/Sa
T/Sf0OxWj9pccOT0KV6nrfJRNqLSFUP54eOUcKqcquR5/65pfIuqWCXoM73anlz0Hcmeugr806zW
wkEACn4yL8eG+vxoUII7RaxNXSbx0jP/cD+ql2TJZaALBHIfSeiEUnsye5j9j2A9mVLUPhL1ftAn
w2kggw+4B0KH7IsECTsFfEnuNH4rZPbglFVoDe3edECG0PNF9zOr5RHbqSp72PBST4Mq0AXuDHK1
6ZhZvoNnJPjRoGDGjN5eDMEV5/pB60G87VAl5fVC/7yzrk6JVfWk3zaNKIQk3nHUvyPMHeN8KruM
+3As/vM41qHd0/ugGdVj1w/4r+lMUaEw9KxCZsfqmoJhh7fPuR/tVeWo7UXqymZp5oAuXB9B5a3r
6F5QMw6RrgRiaySrXznHqlx7LecbzsnYgnGLRqKPcgIWdzMNn7fWFEjFiZ+Ve5c517bQKK+1zWy1
sO31f4b2RAb9rqM+8Sxzw9XwiP5DS+pT39d5VcJ1oiiHVLtw/0PEYTlRHtzqAFv6qr+xyHxenHrf
t96T+N6G1TU5qtjSt3bjiAeX3tBq5O/zQPMxODUstpYzFS7EYgcJLMibh3cynfaejJwRgUl+/sQg
ifUX8AkrYPX8/wNt/jE30LbjYy0NHlR+gtT8aMLpoyo9OQ5yekCjJgQ+KhiOftM+WEQS935AbhDl
ue5eBFeRhPalSjJ4rf0xq51mJbu9Nb+6DopM1E94nZguq/B7NBifx/21MGqLcRQJqTbXYamno2Hp
VJNLvu5CqmbzqSYaPuSsevstGh0xKWgR5yu75yWc2oA5kMSg+/DDnf+spjAWi9UoCNJgBupXRwy1
Jp08pK+pwRZZevDm96owrJ5JeWu0/Tq4lG0Z2uN175ErG8i2VdWQAnGlekxlzfPXXsHX6+EOxnTT
EkGpMGBhONyqH+wi+fPNWXPi/TzjHpWB86g0wt1mtGl9unpxFmY6dxhI1S7sqri8hgsB3Wt3Uv/q
M1p4ggwy/mV4Cy2VC748dQ/GbeoBtZKp9fZ088W6qEUgX6ut4r0M7dWW8A8ibGrAntlDwovWMVLI
94hnbL0NoGzIOyyz/ieZDOUpzVnq39UZYfrfyKQOGtnxtueYkEspV0T0/FCgiJ3ZM+GaLZ6G+4cX
MV5m5zvdZ366r4f8o6Rgco9c2AnQE2DmbK0Uwp5D+jJ0LXNoZGE81zxesJcPVkfXQgSHZFCAURLU
9HY+p2XhYMuH/PtyuWWad0UcY2gEH7C9enqa0wlCV7Jiz3zEWTfDAhwpkIUldgdny8TqQe7srLQd
cCNk86Nq+qrWq87kgpbpIU7QAZc6LJd87+vTLYIADW+nhsKE7GNhB0BfnZ9mSBevGhsfYos+gr7h
mvYASJKCho7nVu2Qy3NCl0A04616ulEmToeGILqNO9ZitjHvP6kJGCiPtPa5YN88nq4Pb0jatMhQ
ZGksbfyf7SPKmW6+Aco3i4MvUA7W/mxY1Yy1LRVTfmwjMlYvqrlkzJgNVNtEPQvtxrBczq/skC9k
7n0kHvBdypGa6KjNQystCkNSN0qvjbmD1lIX2BX78a1mQaunpIjhk/zTLt/jG1DoZYFgQcjVKBN5
AsDiTIliHYYmssNqD0qvNmcOAg+eNcQfFQfB0GGKeuK7+ea3jrPUv9M9lQr3EvaNcvk/gQuMZ9Qp
/l/4VW2cP27EqjYarKQJ7IfijSNXGpinsoS/0IowhQ2EOq4zP1+eMzvv1kVc65SVpxk6IE2dRtVn
a9BpJOt7ZO0DBnSsqI8af8K6AtQbsezdJMPZeY1E7/7R96ysO13T2COltYYO3yY39jwveKLm+sfi
ca6+4AuW1NasUJLITwNhWgsBE20ip4+9cjktdtSGs8RZByzVmCzflzYBUY9MjPq9fxZSNWvDB3ef
gkQaogKLQNxwBnPwjfAyzu1U+EFZmzO4x7UszlgvNCgw2tJ3fZrljJl1QJ6ycwl/vLIrduRkY4+U
BJ2UWakWLEz/XzM9aUfzXxtdg+Bvlc5obJd0A2766wwE7uQ1v0+gXQa73YSCLSI8FO/44Vkb3/s5
PZ/M5506leMjvPvvarekaAoChW269KMRCfgkJychuj1NNAmVxtUqRytsFR/LxOGoRtxeagB2hFVK
/YEY1ALOykPH6EUVl2QoMviTWjOY1rhM27rj4XQ97FJmm9TqC+DwxfPt7LGhlxfR/zAzChNZWC7I
vvEuhIM7vwTALOqDLFEcgjTs3M6CTvG6jlOL/BVoGFcP0taEngl9R9COImNtINalOce5xwpi/fVb
31kb7UHUJMqJ2iO37AKzKbBA6IzBHojxbK2UoxAu82n21J1loP3WMWrJxbxnLUip6L7Q7gzJvVrZ
39ZINa7p/0CphmuHPZKGWmEklUDcYTt+nDvheyO3aKO9xyddajchSdVwSTN/rC79NpDA0FNV6kcJ
pCAwtUhAtD74gFN/8oxctkGgaDJGRYIeIheu77LGluULRRu2rKbycnsFpyP+URbICi6fh9aqRsv4
FdsRIoPmV+iaTJbEGLSGe9Nvtyxhtw4zvtfr/20hCN8+jTBbQAwH7WOrNQsQbjc32NxsvpLwG72j
aYtCjulEsy10JOI5npdtojB+LmDI/DxYeTsQ/OBlMijbifMtajCgHsM4UfPYkHmebHgInkET9xId
ifQouaZdeC3zGOM5TJxo+hd0zOXOk7vEUGlXso8QgyhncvoJxWltLNQWefwlkkaHS+O7t9WiKHfJ
s2cGayeIiOL9tq6gXe288mbN5hCvfDsRP9nCJFQzgLsDAfPttPGs/8yQFIs61lhuvSgJptuItcKX
/j4/QBdoKZWrbxNmprLV0TPCj4LUVoNar3AhGuS+oKR5/3BteLVoTyQCKwLr8LbwcqUlHNmmkgFo
aORQJoWyFMXugLtfY10k9SIMjZv6B5t4PcccodXlisgRMogTc2ADJl10WCEcHqmB+WAN6DTwwzok
u81bo0NQk+SBOGuUcrwiS9euLEA5VtynN5BIROAHDGyJTVCSAAog/t5Rm99eKoi1VKX+OIcrB7++
NZ5kgeXf58VkKTcrYwc1JccTBB2b0MTp8AfViT+LCIW6RlMfJ0aCJCiqyB4FZJcPK+IIiXewgKrv
gfXtNgElo9vJ6pcPcLAWd2bYA+zdsluoyLq02E6Zg9LltxO4MqVFBttT+Ze83K2Ka4S+XLM6soET
syvlsaU9ceyKZVr04napS7mffNoqcF5BTb40J5DtHQiZ/F8ny8UZ1GUXFasowyGB5oNoLA1gKIWv
Y2ybWRwXYyzXCmQaLirVoly7FQIM0RdArFcnTZUFfIiN6tN5w+IZWDs/hiPjoH6ucHrE6NypNbug
4zjcmHi+0wJqO1nP9bvefcLneDTU/idftTWNfquiFiAfk4yY0s/CdkhB8nYUSzM53aZXPFpy+Cyn
pt78gBvgI8yzvQZMnF/3w4/UxmjFr2u2kOZy1YvooPndGyftTWNfD6XVvld0pp8zSEBAXXFS68co
FQnCLZ6AqkhKGqJ4qa3uwrXz0Y4Cbkm9XujdG/X/MUKYbJt0fEjNJbURKYQ7nz8Yl7jOpkyudnjS
9WDONai8JYBjD9FRKLY0DVNf8lB4G7i2oz3wom3nl/e15jEFtdGajDv5JZFXYAaO8VbYISAElz17
IZBWMRdOoIKKqqtLkzVvlCpY1Slgkn0sdoKEBaB9ViAGxUXHpB8eflPrXDacfw9nB0Vv/eDDuCbl
WWMQszOkI8ve0AlHr+PYIUobyUdn+cRhmMIKJoyDWjUpwWBpK/3t7srhym8b5oBsQR5hMhvx32Vq
wASd8geqx5YmwrfTd4h3P66Nx6nuvoS/wzMmhKQWqdSyREBPwt6mcE11F/KKhDiOhpF9O163NMd5
vO0Okh7nSilhmOm6Gr8yPOVrsMsuYNp6P/muFhJWWB8XwSnM5Uc875Pnq/R/H+jdB0JWUwshqdZO
NjqGAhwf1VPocaaCDszoqdUt+4khRPcqlnIgkbtQWj7QIitKgemsu7Tunv2nQPXHG8kxY4ZN6geQ
QapT7knQnz5v248Xzf9J5/TAJEu9f6TkFu9A9zDtn44x+jLQ+2Dyf/Xc/u8+vLkUx5cfFvBFGUA9
kAx5jQGeja4FcTy/AI8OfoVcBVX0K03nedi4KFuc8Q55jQTIxojSUDwUfxlIYyO8mhNG58t7H5XZ
HVdE91pU0vxkSEVOb9vewHeE9JCzuuRc8cteCKsco7EElxc74jHSFPUJxKdsVtEZw23RH72+ywvH
3zoznKQDeYMoPjipxG9vht71Vu6yNWPBxyIUnXmZI/jR46qTRFvtPjihbQwSMAIdH83RfL7+/dm/
CLlRyfE5+XHeMFEFf1dUJGMkATDCSu+R6si0EeZ3t83V3XGBCbh3wH7s3CuF1ZDNgn/6NFZiVj50
9vc6AsQ9rBWH0baKGyKgaG5Kk6L6pc0+7HT1o6MD3lBk5g3eOpBKp3j8RaXRs0xa7NA+lmigoH9i
IQzwBvLCgfgebTVOf7/KqTqrXupM1SOXCfYcegc+ZjnvqKauUyv7Wnd+ojKhFWYQARGilEiWhdg3
PIJZPIm3BY1aIihPH2IbR2AZEgtjYKiKqM25Ci1nB0eRA1/NEBGg3vZ984xe/fn+ZpwYNOJQWUEv
Rp9QWkCwih5cyL4lSoIGEV91jA3IVZ05LewRkHEcBK+ZfBAIDeceRaBDR1wCF0ZzcxFwKViAlVR/
L4NTZv4iuobVSMx3b/ainUBktAFlljMsF6H2J1mhLRWZGjx9LEmH7Pjhb2KHeBAd+c4yFF/NA5/I
F536UL3UmMCG0yLK8Uo2DqEXnJcyxuw0K8ePqjx9q3paGHKRk2FmsU5OuHmipIqAxircP9SuPc4Q
Pkq7+mPY7i2PZzicG3RV42MYaxgPSzpuux9jNIRDfPRZUbxoWONqRSJRkhN+uvPk/MOvTnRTnKTl
P89aP+r6rccU+VFXehDGuAduWZBPmhxmtEdXTEcFCXQfn8PPZf2TJ6A2ZdVLJQzf9DZiGZCNMuzu
YnUByMuXzkkp4TuHXVmRuRm8Jw4pcTialpdx+JImMvcict00BOt8vKCTRn8iCR3PBOTZCIqc2KXz
7GmIkxYlKpAtwcUlkDQyCkLEFJv+SdLVq2uWyYETom9ujJkNFXDBbGNPOMXFRCYh4oZtvwfxyJDN
iiotTb1hvFsXhj41zFuWWcYIh/S5g3gNIUXR6jYp/POjXn4G0kzTxLQI4R8XouhgZqbd4BzXwjVJ
GXfRvtzVwZRMnvT2URAlQUynVR9MuZUBgQvy5RJ7NkeqTBDQMM5mP2Ynb8j6ZSB6mwdMR28/nc+y
o4DK3sAEo39LBNFY62qX1OSSlww0NbIR9SwpxyJ4JN5X56QaPzGbo0YN8sKrkSWcZ+ofmz09WjIq
FrFJLnRGZWPH9s2eyULNMs/qYcBjVOqmzKZQzG0Y5m+5u21j8YXuQb54BqRAPwFLEmKRwwzOEKeg
tvi4PuJq5t1egwDLlGhubHNO/Dy6NnnV0Gb63ab9BjgAFUTPHh8QLAJerVV755Pbg0ibxDiUBeEt
wBMq0ZEKYxbNCv39KlG13F7sc+p3Nc/LJ9K4aZj5lqsxZOlXbKityQfAmY/DElc3KWjmHW9Ahhhc
lxaeONn2fmNE3JMSFlneEeeWYEyfH2CnUbpl2t6raU3LWD3h8BUcegvpC/WH38y915x6ouLZm/k5
Yvz8Qn9RnqJULgc92tcitFOzwYuoa8gTiNCvzIlPm7Ss1M9goF3al7Bz+CPkcSEFM9q515K6wI4m
SmXkGqEpD+Sk0g0W8p6TSIDSocjXikJuPykhYtylvsFYDsCKdgFElpiNIbPy8kVr6ys+A7mHExy7
HU41w1nuaOpRI/t0s0ba0tmOy4ARIaolwyxnqfaX+wylpTvUENCAYj39UEo96Mng9x8LYvrlsw6q
tg7GFniPkpcdurlYkpsK2z3kCpwbLOyu0R70SuUCCHoEd5Dkbsl5Opvbiw8oqF4zHHQOkKTGn/7C
ptPwSpwOHG4oe+SsTUlOsLFfBeYLMLNMwEQ8NpMh7qsIjTo9Ktb/ZSJRHbqvoqtglsq2P9+ImWT0
FtzFj4ABSwmOisdwYuVtAg0nEEvczvaNssfVISbeyKxe0XFaEbZ/3DKLQTJLBOJQzhjxMaaE1ljH
tAI4JPRVFu072Y3UXV9uAb8w/Iqri5VY6yRbm8spu4L6CHzzf4Jcvvu+w5CUlF9UObXR/SxYV4/i
MJk+NEWP++nIfny8lsEivcV/HwyA6I9QrSgphiPsP1QOaTKpqJtWYyDgWOMil9hsInQ1tBVgH8An
tvt6r6Bz6yZoGUeX/66rL2vowiHi8clbyz60+y5FpCC10lftzjh6o977OYqQGg+BHD+pDUflQrQS
d5B6WeJNxnQZtN9Vjv2OpsX/lCrx8UT1CqCmm4EApTIjvkh7SCggwmFR6vIwzKvjOEWpB1uRhmwN
fIxvgR5Wy7zbTqQQzf9Mg9fRgIvjjs2/QPsiUtUhDi2PEAc8A5hcbQE63HE1E6rJCHGmGgxoAHDC
Ur6e/7iarnt8Zi/vEWvhPZN7F8fJJe68eXRQzYmR4SDjPZ5zO3gboZUz8zcSZbeS7RskTZqr47/x
1p5i6Z6EH1tzXf9MfCgA46iH9OvSMQGSxcgFEQa38dgsImn7ngEdwD7TCw5vtvHFcojwDXRK3BU3
VdrphsUoqR3JrtPEGTqBNsmFJht06Pr3ASX5PK3DvJTI/PQD3IHN13d+FaX8XoWxRJJzjw+NqV5n
1+nQZXHTmNh/RCYVZXCebNy7r9Dm/phvbBJuzlVH+9BMk2tJe4q9Ubt1MkmdjM0DneEaSnFXw5ii
y4tEoKcI9CAp7qy5/2/wMbHs2Q6B0EjMvzjSbQbmW/hrBjO83fgC67mQYEi8GIF+4kE++nTCnziw
1bEFZPdx3iC0kR0fAXGtY7n/Cv2xcEPWKhgYWvlMAzQiqJAl4AX4x9EThycBt1W/zhYajOsnAFiU
lUsjUx9+qJ5QgK32WJmt6kWLiCfgSrW0DJXreq1QHQt3HySozSQ37p5lJbWwC+EROD+rz0rinxx7
Puc7OAUfjM6IHLTqM6h9hKX1JwCr/Ha5kXwYvMICa5fdYLSnPvY6+QuLwEUBwDm2Pg3P3KX4gJAB
CRD53nHG5KJjWyjzCQMsrdmgOydL+Gx5154BnQKPuXhiRfW/1QYDJxnf2wykGOaaibLRJp2ISn50
XMVCCgBGk5ELgoU6P+Wp6RrX4xJ1XC0HzWcY7Yo8KX7ZfWCA3ro4SfgeWxq5pGivUygO6SLUucmg
vPCz/+9cYJI8QQ9uf5zpWscM2DWn8fQb22Wd74sB6oXlKFbk8uX5mVoNzFzZbtnDEg49E4XcpEFm
IKTS9zm0Jn/3oyalebFWWOlDCBxrMu+gS9dmcYcmfbRrtKCckFKM4oC6UKJNl4SA19mcXyxjxNbw
L21jIIjmPpmsYfx9vCx9LbqlOlKKJPYgBqNQRgjZXh+lyZqnZVVkfjQXNGRRLwerYZr5cItlTk1c
Wvw9CbkTFnhgz6IXxyOy+xGosDc0uX/xVpcPoqXc9GH4w9d6f5aBeXZu3DJv7XjYqbqKXUgUlU4L
bG8P/Wh1yieDF39Fj2Iu2gbwIm/GN+Tb1a1jr1+CPVywiAK6nj4PNZ7TGyB+xXZeBLunfCLwUR73
5oHCim9+bfG79eyXBVQtlj3jUORuta6To7ijiohzyo/LLjg/CETpK7My5J/cmV/akbvoGU0HXqEr
+C4YlygPpPsSMJ4H4s+1N/A+uIPiFkmplrGbOp4Ugq6NaT+MZo6JJ58nWfxrqEMjVmdbnFN+cccC
EakR0sUNSfSeKRXiqXQCZhZsPzoKXyntLkgRqFhfLq8sgkEhSI9iV9CUSJ+mzu0JSc0BzV0Wt6KO
4lD6/wDupXXqTmzTQQCuR6DffosuJU78YsoI4y1uQs8tfEEu0iCy09ngbkY4A5Eo5yV70x1x5rqD
NDhuiBe29snT9Z756KCxC/TG6G7EA+0j3ixPqHaX4xEj0gP2wFC8nzAxjxgyLNlnWJtofyRE80wj
RmbvYB++UnwPPEPE9L/0NNBd/LxSxQtrP4tUdR2B8EqKGau8YW2TDSPJCt50hzhNb5wIdchqVsJw
f7U+ghZ9/H6IWmjp+0qwsZKLFbQ/Ox8nCmZ+AuM3EYp1q5Gdx8JNPisXmv+TeL0Eq0yFEkiNfeWD
oqrd6Htl8sEPYT9GOb5beG00ikJ5yLnRMvNFpVrxb2bOib13Lruh+Seg6E6yUUg1HigxLtrS0DcX
+qNgl9Zz/CVcv3NifzG0dOMBQpLFHFQADk+KTqnWjMVRKgIfMV55w8YjepWAwp/iKWZIyn3msDgB
kfxPvHL2x/+3RVKnANITPbhUGEklcy1UrUwIrj7VRMaE7SqXd9slHlF9Y7wI6g/IKE1ZLnml1rJy
6cC+mfj+G7NHeByxh+1gbMbUTeoxdPs9DWluXM+5wowkFjStobesFVznxTVmZk1PEx6wXapbMyhJ
kWU+/6v7GaO4vwLgHgnWDHYyVwHvJFdV37/JQlerUSEgPUZ9HdkLSei7HZto6Q7coWwTteJuyDFB
REHsPPXMAvv/NaO8jyqG35QL0Iy34N+RBSnx3k2l7N2zhhP4ivKZCfY2WmkZbQBKJ+Rm6H9xJ09b
/q/x4oKKqEwNE/AoX9P2R/aefuteoFGeGAW41X2+TJ790wjcXRsf0uzXqshuXVxzKcuko7+N+wm4
+xH/th141JCeJNtZvSHcv1KHMVdUTjsNuv3E94w6wp1UJ2X+T5S91V1i01tpD0EPMENkYw5JBQIG
WPCkIeN9Pq2eYskKDv+l5RuDkhb9uUNbhS7Tuo95uosu47RG1Pau3BY5zOAKiE7ah8jqLPpCxdBO
mTMSgHOuvu9+4N3dG53myuT/NzVBP+BFr2C3+7abmBDXeqI8R6PZGe1Ci3rN+8Pdqxu2hDasFncN
UdP8+hZrRL7b6i0Mw1QOLbVYCpRbBhlYHvWwCzlDhcgZjEej2WURmrlH7PWfaJTK+dmHe2KsEsWg
9NhGi73fDOIlVWM4J4DxJlIZeI29VfNmW5M15HPAPetb66uO1zB+46IKhk1+hq/H9RmNrxDoZAC8
Pc1FGJEnOKhqsr7POgsDZLbEML/tbccMn26yMDoPhLd/KCJU7B3SfxA3CQjQo0WsJg5t/na15g9I
yujc7UBq7CXK5gLDqBtdmHx6ZnkMWhNy27f8ggnSMd3Tmud1NtiYzSkcoWPd293IJsPtPouJYkql
9hkPfx/I8d4oa+PEz2Dcu1DuIzHzev+GbgWzbo7tENRUDpmLjAS3PaUzuaqLVtsFIeHBL1rob/La
BOiEoo8RJga7OQyd+N8pLFmRAJ+cvF+suUr9+ZUtb1e1YQKCxksBksmNur+N5+XB+MVroLMc/rnY
B710oQb0bd/Z4ggmwXwsLgLIlJaoDY90nA/Wauj4MIy26AcIpbx0x4Uwx5NAyttii2qLPjSCrr3S
yq1CqZ3TETlA7+d7i0wFPX1rK4gABwF6ugmzt5GmDxEhRxSc441OnEtAgqxTqwRy6ui25bubtsbX
2DGsZeZisuBYFr74h2KdEWET8gFp5+6mSy2HSccIRec1nz89vCtwNQ6K3oP6IIYqXdFQmYPOvYm0
u0rAdbTEeCqmOUC3wDPCbzRpy8fU308xisBBB7NbxJVDE7Wv1HjQhfMM+mDqlYI86zaPtScWHKbo
aCZt2KUfz8/wJ5sjk1IOTQ8KQ7UpkLtLuwNdUt04ZH0tlkPZ4ve8rqdoaDbrkQVvs1xHcO6o1FGl
TqpiQJbCAle53Aycy3xvxbDTyIRL9ZCgSJ7ail9y523HedqZ8AmfoH4QM2h/9et8V5+wM4n0/GDM
V8xsJqWPFBsQCrSNAXdBtjqOH7TniA9C4+NVxeiPIghudAcphT80kNTZPHpYXbfW67OYwjl2kWRE
K+EoOW9GqsCSMYDQ6ui0KN8K25TCUg2RWugyGApWPcCP6VQMUkcUbFSDcaQinbBzYGEOzk8P2kzh
0GgZ4jKNX1DkN/6XIHoMpNDdgLlxcEtTy0qiiAApTEz0SQlN2dCKDynvBGF2dRYb0nw1jMhhaWkk
IhKZSI946YRG1n5qd0bVbhA5vwwfbA5T3/7qhAI/IJo3i39RTXULXdJXhceOKWhTb/kfJ2z9whMK
4RH0dk9mcfLesH7tVFthMCHUtZQ5ZPXz4O5B5dKhJYnSX5V4tzC3KRpsf+rJxrLrDwqEpW+Nqm+/
mcfSLrrVzPBlU8KvIW9QQ+58OQRvcTpaHo0XkgGR+69in5E8eRi9/kKb9M6LiW03E0WnkFbJShqR
GxfLG/e9lFSO+o7u3iZGzWEDyGv1Q+qSdiWT6TKB12Fy9QN0Tkayf2dIQ0LSUxGKqqwthERZNQ8Y
0CUzCbnv8vsnXgUCGwdJnv9qyrEPZ0RdhjxLBM8MzDo8OHrks7S/mis5XJTbn3JUQz+HXoK1viTm
/hHmvjaFdQjUuvqEIV0iVBWs3O+b9Vl/bMxrBNAA+FFDD0uUwDi18t5dMpmr5Nf5Kt9HG4kWCpFC
lQ/295oMuzSX+HFEYVEIpPu3GVq4WlHDqwpCCYEqVKG+OCfy9FzleOQiWj4O4MKuVpUG2veWZXAm
iBXsg5vrxD4fRDB2IsVIHtuiM1CkGV34W/Tr+W+OrHAHlRN+9EF46FTER3fxkiSoE9I73LogmMIJ
s8Fs5CQwqEoh+BduiUS5vblwsW/mn8oe0Mun6E+zWVgDS6ULLD3JgNVEMby03PogCuG0YIWz2UJl
eyTkbPcFrLI/uuuUvZMb9f8XMGRkdmNRfCIbwU3d+X5/Krojke4YARXXyvgX2v0ntyOz82oWL2cZ
GOO9d8GS48EowYGWQAOKnRFphe6oc67NWMpTZcQZv8rjTEM51dcc2bXFZ1BNYt5xarCHoFDZhhuo
JT7lfBLSuskdcb0Rc216aWe7QNKFQIN8CsDeqCsKVHjvZAuBWcFxOqsulei7VMi1tpkv/HtKgvAh
l3Gi36PgPs/KPOPZOoS8e+G2gIA6klKSc5lGsDzXPgvSfE/HOqmUutlSdzsKAng5Q+4qkL83LLsV
7NVV4HXDUXUdZ4NGaWYrvQ+a6DjAN4aUaSHM4mZhCdqPQTFUkBS1ObAhNaLisFQIp56hhfnLJjIP
sbrNyLcJkoZbUB8r5/WF92yIP9kQvDaO0mk4p+8MQWADqP2EKh5EtuG3ITR/1sV+BgfXgMv0UjQU
aPdQC86ro/DCloB0z3O9ZrPHalu5IoybsLA2R6RKweGTJn3L0NG7wSUWP1CrKQwQ49m5OfH6IiSm
QahvTcUi9pcxY9rjLih624zy8ntklZIKrpFjIz2gZmXt/wV+vDqWQ4+9VONO9DUYOoGBIj+RskeY
pFY57LDh72N8tveMQQTZrJxOL+nDp1jygfq3SvUukuB8mlcOD7FYcFaGVEAwjNyh35W4bNFV+e6j
2WDOWyxZjl3DiQBZ3hgRBsHC24ii6SXcv1vFLTZW3tFa7jciqcP9B5XqFQYwyuO49OkhzzZ8iCj6
OnzDXdV/RT/0qmttpcmxIIRwZds7VgC8wwaDZEG41KyOo+xiLXvU6k/I3ThCfMScAxBlErNR8MYT
bgLRVKvJa9Rn7xIRzBZVNeECZT/XyrWIK+2eyzgQnCDr1hdEHN8/uvPXbvF/Qnait6mCZKpvDiC5
OMgdQV2iXZ9Kb82Ss1D+hNQPkT3tidHBfDI45taJoUosdehBwyL9JLJA/6P70YNGkhO1E3A90ZQ4
ugjMuIdtPd62LjJQg7mK0blQg5ef6Jfz39B0Az/vgtNa1LJyZ3OR0lOd1Q+5rdGC8xfna3FVBdYe
njsmb0LlqNPZtPT73FRX8OfrmrfGtXNgCm+ckzuonIO/Yf4Fqo62MESEdx+mI7GIPfvfh+DheCZI
mBpklJVM3Zhkt04n9RlLJn1yoEB3EpuH7hGMardRoZCVpcYFpUBwbxfhuJc1CmxB0bygdQvZprGG
N1CiNC3JzJbhMbue7Gud1eReGEkrpxChtfqMN4AGpKbb7hurZyfHDdeXkOmzKyyhyYp3oi+ApA/b
aXRDhMOIbgy6RAoKn5Q/9JsbqTknihrUgNC2lQGNvSZynxLNfXwJKn7vUCQhKH9+6uhh51FUP55P
Sz1F0fRKd9YbCGXCZ3wi+VYg3F9BdA91cwWZpMdEF9fGImZo+8d9Cw2BHVa/hohETiSZVb4EKRgS
gu3402TcYPmdn3XyCMIlOmaOlk+5F5OvEvUoxSTxUJVxxQwIFuWJKKDwLMtHh3d+aViShOF6MReY
LMm//t9KxSPv3g2KIxosgHHTORW0Jn6a6DEdbV+wtVHUgpP0qISETDL2LHQXBISiCvosCV5NTMGO
XL0ZRHFbafwbXxU0EhddTZSOnp5j25dOXCfZgUR4+6Ycln6YJ2KfHdMwKrAawsMsDYUC9NvKy7ZC
SZKYPP+8dOQ4ZdVIyoLTrij+7fWxAYsVvG7FTZ/xDPp2fdyCpcW8A/f/GDkRH1pHLGsRT/uDTeEv
pF1/T0TRYYdvC18ji7ZX5+P4m7MXSwU8OPuafuuNq/VxACKiVfQUSlOIsXZT8Wsbilo4yADLA6RJ
urB+rI+EgDdGrxQDIY1MN202/9J7ys3YsUo6FocXeL633cCAJ1YVn2/1NFjAE2C9+iDk/huG4YPz
xlH0o/rCnx3aa8nQx/g3GXG06R74432NYAHGb6GKvye1KRdZ+r5XGHgo7cSz0PhMV9s7kkGVpGTp
O3poN5UpDOwbcPYGOYqwHSuMt2aQnGUb6+Z1AnkxKFP9WUK5VdCQGp0wXdHfyMxtokPPHY0gLls8
0pXCrBRAqDn9Q3+CxIrwkz7abg0V/Y61gF72+L/BZTDlr7t1vKVvoEacnRmbzEEGP4vpcfgngXeU
gyEv538xFB1UVQKOzz6uQ+65hbDohrw1VtKjvz0HpQDMvQGiiG+ls13CdOG4aOlkFTdn9IHngqvG
dcWKtoUM/QQLQ3O95cgrT0FwSIjQgJogoV3l8zl9sq7j9HL8hdtl+W6K50ZeveMYzhfzLO1ZIkJ0
z0sAwRjQF6b6FLJuM8fEjfIuN9P28aCSh3WJmMWJ+Xj0sJBmQpL4dWtb/C656Hzq8d+bPKuDJTzO
g8CgaWF65SOE4RbFq3wwr5J7rM+L44aWrL4gnKOS7wxNlruMkOSipXzpARYYA8C8v4fV0yleoJYH
9lpu9tLzkxJAi0WA+LJowKjEAXgLXco62GxJjAKQFY+x3fhXNWTDK6ZaVvv1oO3ROTurLOPYO4Bk
J3nPxCJ/NSmgjcSa0TXxqnHuGuh01F5TQpbdItThVdr0gaJdMSExZw5TllXjEXInoDmEU6Fhp6Jb
kSIZrZ0pVBjVoOFC0E9QtsknXb66rJOm4IbucL5NXnhcpbsgERyBpCQNhWWLBz5EJUdwmQp6W7ZX
awY1EqyquxSMzGKdnXK1sU1rys4sDzd6X2kyBM81uw1dyqtYlsjJEgc1VdZIWOeaui2K4iDOGUKH
FUVSN8+IrfHE8tv6XC2NWMCv2W3W5ODO3qHCx1OBmAP+Ph3DAjsVRwVcqK56YCRM1F8S0VCcm55h
trW1/JbzkFzkv/hZhmD3s7eiowfNrd9OBOeXxPUVzlwlY6fNN8qGRZ68IlWyW1cImBJfLChhJn99
xmSTCzeQAI/a3wIgq/Pz1KdWxXqLBNiDkjAhp4AAYkXA7en8cVi6kbsPMPt4K4WC2bts+gpqNoPl
SOGg2J19P1UlxmaT10NVGPGUALJXyNA0FelNhOA5UofiE0vo/iD1KTIuQCteWENCdS9NuQmyQieL
LBZuwSiUluxNd7UdOKiZJfXAdIQwkQyWhTXdbERbVHQKycokZ/zakMwSSY/RByvixlTOSmCMjgeA
0nd0s3qbTwPtjJU6Z7XtLjYYKBjwktc5EkvwXLwYODoXRo1cesYSK9gAAYfSGwghBu1fYeT9YJcx
9MrMiglhP6TMF66HpMoz2bAf/74j5Qc8KoSvLZadIJstCs7Gqvqm4dm1Fy3jsPPL3oO5NbXL1j8O
pQ40GKkSGPwq6SJkI9f6aY2fOL0wAXVrSYXyeKTQsgx+6BaJfTk3JCDjhbJposUoJ+qwsbzs6UB+
r1Sp4+K4jOfkaeb3RorYCMxnAhRBgOFY9Olx32qk8iUABkBJqAxvrjmnZXtGDToTBVz4qZnHU03M
qw7fP8S8G35psT3mOcATWydSctFDoauev2/1Fj2G0Modk7pzYYfmMRHFEZcVougfSri/ls0ODOvL
PBs1C6tbKoUmtq5HqKGkS5q2Odi8Z0956l4EGcV42oIdUqP6iAH4QMWE9CXV/VGerYDTyuZZ9BVO
Sxo1QX+1nNwcakxh52R5aoZET18OMCwPtMLJqvm+UEkvrCPDdeqiehqb1UmId3fgI6BuBsPcJCRH
nbZ88y7kNEJhJ9pgqivCO06jhr46tuEGgXI+x1botE7EJmu4Ur7yvOFDJXENez430sFwnOmwMwxv
ekN9dAkRa0GLLYp8lLPZeeCA/Gh9mEDpzD5xEknNs81oc2JszETfbJD0QJ1UYbRDT1O6vdPD/4HT
4bb73L4QEnsnnzfn7IArTyFO2V8MsVAfCN/vqdPf2O/lqdqtDCdu/xHtcQzII1w/SdsfaM378soF
/hFBFrUXWZ9fvK6X7/kX23DrTvXEs+UDER3ZK0q7yT/wU8GIBECJLvTeB0aHGpEEEFQ17dSVfsNo
BWvVbhifh7r6Ft8XAUp2lThJW/AJ/hp43NF7ex8EcJTg5JLI8pNTZyyZjAYZPqP9cVwLMOp5VI92
cEhMq1xPPBswaslMqmfbBHw+HwXZlph9wZwsH2/bG6ewOIfQeG/tthfQGzUXN3e00IK67zbMxM6i
bNYDVChByDjbKconTjXxRcIXxxHghX7fNYCCsjBAM2IlQPdnm36rrp3MoeZG0uZ1RRiKilKk+Yy4
gIlie8m5Ff1y7ox9buyrzgnOT6QHXa5RSbZgfv0ZbrNIuVLg9Fz5LKzxmRmhc1AWCt0ghZ5+h08E
Dwd+j9/pka2rOyD0p2pxX8o58unUQim/7XvzJJ3yOfCMlgs+Msv5o/uB6KukEEMN1vDQzxCwOs3s
pk2df0uXCr+6eoQAN5Bda1Q/OEVQnOPHeixu+6YPWPw5bhpTieiLNB+5Ho5I76HM6Dk3u3Boj8sm
F+EasPQFWXhu5mlNe95zvnkIpZv4Gjv0IMH0eObztROQUWBo+BdCHO0He2CA5x2vLM9qWRGGUuSy
pXLFplVKRpR/yASDJIsnscTxy7bV8n1FkEAqc8py5OS014YVH+bPI0u3Po9alIU8GDHfFDqnvYCz
ZjNbFvP2BTP5dJBUQfXyWNaZWoD+iLYQbzbW5lmQ8BelkwfisA87pB8IevF3MtFv9ifemTx0fGjs
kHMJ6YFm2C0Fv57pm582Y5uQbkRPfDG14b6Z6vaUicfpUIbZnDmk9a2zQavIpGVC3Mt5j57gyB52
GkDEs09/F1nvquYdEuxnjB4mInkKbhTT17OH/lKmf21RS2RWw84ConkkfqGUtm9F2Y0xqTv2tvGn
m3IsxjBL3snkVmaNDJvaabcXpqEa3G1zKUPypyqkStYeiQf3nc6bzse8PT/wGsaPYR44ba0tS3QO
TOLvQ03xd0dmbKauETklFAPScAo4Ej4q8beCXSRZ9QLMwYu54dyesNeEol4ru+Pbp+GWCicEPnu/
wElwukG4++RqaQNvjWpsyEOmmGvdPdrqhs9C3n0qPCgB2AVobJIDJQOrQu7IQwiLAf2ItuS/d+Zl
IRjbMA+EfrfcpFbUCEz+5A8WHhwUO0ph4TeeMdAq+WV275dz7DOG0ovM0GMoGqfiNB0ABNywFaqO
lqHFN09H/TQugav/YmUWx8Xk2ENtqS4k0s3O0o8slXW5o3FbB94WMLVqGKVXW+3dU/b5lnX6Tred
fRyUc5Uusv7MiMhzbBJnfl70Z+hWs8G1crtTLiSghaq4gIFQfm8UejeGoELCKdFew2ZwIREB/Gxf
IXF8/odRqWG1zydJqw0n30IhBsWGLPPiarGn/wFUa/8o1GTCICd1jnlmcx7tOCLQDaTXhhwFn7vM
JhUajDZkw8iGAOUdHhrX9xSXQEWPGsqvBxMtocNQJDLs3SabqX+4vx1vrfRPTJT5Txs2IS8EZK2Z
L3vypQ4mLWvgSENbdjVczD8aDtjbGwYaRvnPoTNa7YovOsVbDzeo61pHuBQcOwu5ZshoZcO9i8Ra
fB16B9ntUZ3rKQkkjBpdN2KPg3aDaUhMhI5XWLlNhwyOQw/AhCqQn5+hFRAgcvPlL721Y471sN/f
CLMsmQPgpTDwpH+omJKzkSyKBtQ8zdpMitSFUcY/6lRiuGQrOhyPeRQP4TOlZ5cEfgydDB+QWyOg
Zne+ZZOyQMQ2GL4ekq9ESdiMhoknhxIqr5JFENa8X1heOwwxKgNc/Ma5geSpnMBoVPYuLtk5lIyK
50hNsdgiU8a86IYD6nnZ0TnsmdxJH9/h30n1BYZ18jX6JhsNwo9M/S7Am0cWVBI0it7KXyrKrPhs
d7hVdcGynAttsOpgDAv3yPskTzt4r6bxf7scCophpfmwPe0SpfRQq2NVTYHJib6PoBShzNtxUOvx
N0wAoIx7J4k/kCy0PnrTE5ZEZKetAZl0oSjClZ2SMM3ugJOlwYk94mfHxMPlCUIqUKxvuiIeNSmC
0XRI0C/P0VEoS+Wmk99q/DaPwFQy0DTD1M1Q7B0awYEvnDFLZ3qvY2P118t9lIp4vzD3YlU1uxNc
EXacRx3OU6JPxrG4ADvRIv+eNQlObsV5rlsZhijqrvW41KiR1lQ4zyGU+F7PH92iJcULgCtzYesK
edtKbFlICCcnRfCOU9e+i6NpG4yi2A/XagIEvhT9vpYi8xtZa/utfWgMU2jSXzlYyuYRxY5qyRSM
xc3Z1LaXNY/DaNkEL52g7Un7wXxln/tNe2Gl7lrfN5BPriyYOg3Zpw3RG7HSyUuC+vx9hb0nWw4p
1OtABKwi9+BAmcJrZ6UTooklT7pE07jKcI+Y4GZGifqVD+oZvzIyte6o/ykLlNZpxM3DxBkp1e5N
1D227YeoeNGmsrCnPwrbMFARcWlStrC6wngykfhU2LN3Kk8an6Ucm6qR387wBru6umgLnPJBwAkW
pNJbGiydkK6VMRq1JJNanKSnGdEIIwzHFR6TNXt5yRLtnstsgHJluGSBJsjs83e2eIAIEYq9hF+y
Unzi5WgTXgVZ4HXPLAVt03U/ZRRvG1ekuyItwM06gGA/Puy6sMrGJBuadEYd3FuYXZdC7b+97zJH
MzudFoIhUfmLt6JzGHtgi+3ubRCl/Ml61nLN60RszjZLvVI6n9NlTlnX59JBo6Nt6awKxtIMPXeZ
YayvOnQ7YdEFLkhQEqkzPtAkKld9TUT3spScuBePPPO+5h0H3fi8ghwHClntVMYJfz9dt2PBNCYM
eBne9RPz0mce/sJ9bzuq8QBF1rvlY8VTqgOTJdo8L3Do4BXS61cEDzdO0JkYZOwxoKjvnnxwxCBK
gzSeXN7NGFj6cwZHdJohQDfQxiv4ZX+xgRI+27aNTdKG0k1ZMHsZeEk0JzFDOIxQw+fJfqLubuGA
+WFYo6BGzkjkoArCpGNls0hNzs+h7H/7tOVtO9qyzBGMxZ5k6H0i8VxoJDPJTAxksrKJuTX0aHWU
GNCZVbrs5IS7R7EAEFMIQRB2gU19Zgp4yj5V7bP4AOqCtqmK1RB/MInZKAV2I+FSoszvDgm7oN7I
ZMdtdR2GOPh+eotCh+JlBW521DCzHEHr6yE2jmHINM4faGubHG61eUX/uFs8rkdArWdICkUH5qLo
s2p6JhdooRLED5sFTRg8wq4oElkY42o21wzJKGRiPsxHYqEHQKHeTOxiYxF73s9/bpem23RsgCWw
i084ERWyrAp4nxDg6XVKKTz3ln/7oLfauHaxyiVsyM5EKRkO7H5Fw2kgOfDN4zvpCfeLU9CZfJqy
XkoJjEFMpnjGLrpqofXNTz2Xij9PlVmXa7Gv88ay4YBJYOOWwNT08kD436al/Bhu//Lw+Yyal14W
1xsS8jg/nH33FajS0P/NQBejWyoX5MVyoPrcYTHf7NxApsHZi9+C/VHUOcTHyCfkdbf9lHn3oS6J
ilQBE53HkqiLjlgqSWaOilN+3fjHAcE2IiuB+loWR5jItsqH9zoD4kXdJmImKbsG6uA07ss+oMkZ
BZLUCRbLxokQGmLsCaOJSW0Tyr7aapVcyRprPUm8PNUsHP6gvmfg3QgFeOUnXXKNHXvB0g01pWYf
veKH1gdkpSzEzhfT0WcofyO+HiLEcTu4HLEZIfQDIp+xC3roaMJ8NwCUKrtelgxC26xBmh7FT86L
i9pLwzcYjIQGdY0cmwrBNPQDXv66s5nTleVqzKNh/qAeAnNFY+vTgEu1rMX387sYDZYsRxzkaypp
Atez09WAlcOxgL4XB7IiFrYuNtqNT5+J3aZXqVd9glIbZ+WSfNF3NZEUwUxXdL56H5iMcpEA0Crt
XjB/HB8lCvlUsxF1qLRnFBtM6fku9YI79mTK2PhQ8KORvciYj7Z58Fy9I2BIVayhhV7yen2aay4l
iCbnc5TBmRGcrhggI5kOTBrmYcCNeXtD4KBtFECWz5CDsdram9Hm+W+FBjquuxKIN8lKskpvSsWg
hlgFhely/dkAdHoIUnHBD3cE36rfjk+0y+OONNrVnzeCBR5zrtiT25c9kEktw3Sv9FhDBvhworo9
d0AmWORu53tso3P8T7lxwxdSP5kiQd/xnGiuQ4hKNzcm+mQB1rc8ZJqo6AoFfJ7EF+/K1YIue8/V
1iWKfL4AmxEQ6ADLH6XzJtR7dSX/9Dl8zmUYOHlVlYvQD1ZXHqoV6Wh6Mkzqx09ZsfXJPMbqesGU
qVP6Xwx2IfGlw5mqDLNBdYyyL3+R2W3dse66oQxOMpeTv2GIOczm6+EJjfBOwx64DgKCCkyukFci
hNn3Xzc0NInjU5WNgzBuUgV/ANYFjCp7DAq7/M4prVaD9lEiW9G7dKQidngzM9MIQyHYL2L67uRp
fDChCTXkFxFMbyYbiwH1t5kJHV8h1J9EleAKe/cNM2gcwXXFG9esXzwYIWd8M3FiJIxR8xJ/ykct
swiewDLSYgCRn5r6XbOgyTlDa7mA64gAwialCXVhDw7zy2aDZObfz/CsiEg2hsfVudTlBHdLv/9K
gitqB9WKiE/AD2Xq5cU+H1cUf4hPqaJyl8wmgA9Cpm9jn+nO3wGANE7Gcr/ZTkXN/ffbeKvq+Rj3
75GNIWtdIIkBn/6s5njcxl2E2fOGp8i+uZvbay8sqfg8JOtQ+jqyYCVINtuZle4b5bpOjP7RFXkr
YbMemaR0QkMEczJYf+Rtuy3TaAf4gPWyzXZq94b3bv2l9boaIwtkUBa/bu7keIoxkl9hawWsEo8C
Xf8u7o/FHYy6GWZ3xMnRTFQAsoD0IEoZJhs1MM+rgRlGEQzirQmRp7FkmsxnbQhiNrONvNrf9ZPw
8m1LeyFm2lTqiH5xIpThQ13xCho4uwOf/vaT+mQu4UqP8Lxof7c+6KHBEBNX0ZyyxluY+1NNSNL9
U8fMirif0aJ4sLpCc0t/6NLH0qnT5ntoeBMo49GiBTLleSrmE3/+R5/pyjenENSfOxZB3o6ZDA/Y
Lx3+afTYAxk8Vy/dXDVymkCnBffzDd9FGrOTc9oAdN0GA2Kel+h4xMmPFkbpAksIMJOrv0G9WEbK
1pzVcq8IJqyeg4TYmJB8ryI+lVUiwdRIWyZAH0XUo2/IYPo31dA1/LWCWOnOp54sxULSbCSURGWz
3FWUeGv0Ysg/8GFheaRXP94vRSIasusN3NWZiE6zYgO6T0QtqVAapFWC7JJrF3jVpM5gA17ajJfJ
ELiiBGDAHk+Yaqa/AV91zg4INoi7O00xQyRWI0CRjrqwnJylXBzGGJdQC6zdPrmS9VPlfIT4872B
f2Ijjjpv0pR0MqA3GqJwa+n2Qx9t4RvfhUFf3kOMN9zv4EjfwpMwk3QXWuFavkb7WoRTsKobKRzR
ecGnE7f2blgRa7rCHUNd7Ug12prdXLsd8kSkt6ExYeXfVMV1NX/vouSJ+gus+WWgkwjCLqOACWvl
5KlvS7xlEEaUnMR6hSBUrfPQJdqspOM0zBgr1KbWEZLuIjNWkmCCZDVnQ/RT6bMuPVegbFxIU6X1
x5ndaPchGFCWdwpMHJUDdK/9M2bkbnGXOoj110ipXP8rDe/+FVlTozXsFdaXdoXuFuCzSbso/Uys
kE4aIzqgrp0a6RYLWlVgG2mS4txVgC69mIlMxD0XcwIE3hS4705bz4s54S9j6LASMTwuJrn4PswR
TlDKlEvl/h43ei0UqlM5fbNMQj98hAF+C/OPj0ZAekKtMwlKQIQ16msp9lkgoHj8uVYxEZiUG0oP
xMxOaGHHlXGurDAi+3Z40wr2AI+PrUqGzzu5LlQMyEo4ZninICq+0heJwgagBafW6MqEZNRHdR23
myUnXyPPjd4pJOxIalUxlm9AbgKL+kbIJknP2j2hrt9DUBec8Nyj7tYm8uwKJQr5zKRQrj+Jv1c8
RieLGTSDf6RwsJf23KFguLuT9Ehq4p/dWw/bEpZcwYimImt7mwOZZ7rK/Q4tEs5uUgrO/qVdbkNm
kts+AE5AiI+k7upvs6PubtaAzW/OAsrJzbSnIqjD51aUq8NAHGlR5XFQsQnCmiw0neqPRaXGetgE
7G9c9eHmrqAucEcYLzYcHBX9WKfgp3ZQsBrQno4MCikxWpCYZPOOO+Gr6MC/E3RwH/SJ0nVMizYr
e5XVRqnmp0BNKfHyUGYxRHWHah4kN/D53CCOzd9hcI+StLBq5PVb8Gpp2hcJdpHA4Mg65eMpJ7mV
9UJMDgj34PGYWQASpWpckgT4HT/VuU8ysA5ankN8TTgls7wTI29iUWt555KKpcD/JbSHAar510Xp
6usZMyNBAAhjgAoNzUcPsrMIVk7goPnOAGZTLAIHzcCO7uLZN5ilP8WAKuqSs7izKIOuhH2zEvJa
9C0fYhVV2uRUhBJhuz9qc1EObyIJWUCmDV0PG1OGSevCDCiSveDZ3Ep7QXQvHOgab6FKeEaB2tP3
Jpe0E2DjNOlYUTB2iJCVp1oLdu9lAiReiO+7aK8MTmQd/Ry336NbQQfebLMOtdIoOegJT6pol5vV
WkfqV9KjSTkkqsyqH5eQobHENP2GOblHuARIwPEEqm47t4qgGJIoHCPxD/KLENnUo5g+Wa2MmLmN
uvPfwz5SmMe0/VkRKtAO6e3cn3YDgeRi6wrTdkA74SKfKX+bxtfiLYY4gWqqlRTlQ3C/aKkqAg3n
ZbgvPHRGMDu/qh5DTPi9M7W/BfokGKyqL27lctcTvzeMG7Jt+7tOS3mfRU1SWh5NBw03KKDRCaBt
WNgHMZOvqoLvbpjd0rLSxNJ53Xla8e33cGAMlc7/Afdv5tnQIGLtoRirzqSZpK88PosPnnM32n42
AOe7onV+K3d2CApm6MhIpEfb1hcktsCEuSEB8nzVOvduRsrPzZDgNRSU/xxau9VjrkdnPG9xM3oR
Sg1G1DGcyA4o+T8FxOhm5y9E9jYQinegatFN7ER/VHuw9bCaYi3Ch+gggSOm9MEq0A78VytzGFpz
hcZ5hg4nZ3AHuk8cnhTAvxP0mmd+YQPAgVrWXZl2oGnAIIH2QeOU8fYv4Frpm8BS9BIjVvNLVvmX
bVBxGeJyRqR43Iq466D6CicpkronSPqU7tx7u9XxAHIgipibhTnd7S50yvoBCXcaQX42h3gbugZ9
GlgOxzmjLhsNTMMFjv4tiv0cH7cu1dhweSS82uoPs3i9+OVHdF3erZZdziZkuLl/8PmOvLB4yun+
3I1ULCKu38iKXyC3HyVmubfwg0ypJwim2lvMh9GGjpiZ8UPVizjfDV97QCOLgBj88T8PtXy4Dqfu
dRXZWBMaR9xflZa5Zyg605pRmv4/YGpyUcme522jgeHLqMZZ7c5d1BFuYFeiuHBH4i4Po1y/tjih
tm6W6OdIIuF9f8QB0lYlPg8yDyVqOMB6E2v20KBb/aHldUpGol1x4sQH5lFc+kAADrH5poChETPu
a9sAq6yX3ELMyIevzpe0RG2YuLPNZajZb0GZvJvkA8JZ7p13jV7RkSUKkKSszutDEDA/bYAXYvtx
HezGTs/LU1xQhOQvRJ2zae3D6cKkWhfqxXK+pCIu07RZz2wvZ74MN5lAN/VR217O/KFDC0byK9aO
dO9na78j2+5pSSKjl3TylDag27pxwDPsHaovfam59FTK0+e7foFjplyySJpyHp120I5k92b8Jbsu
m8nnPt47I/cBu2fdJlgDrM/fghhKYIjRKxjXnMAuE4zEtgY6rawpb84fbmPEn2nwCGHdTj4UI6dh
bnvuEIIqvoxUYL3fZQDZwXYLedaxEC/rNh/1X5/z82FSxcXIeZyUiKtZ7gDRTJFcA0RBWH4eVwa7
PIYmES30wEU3TvvtMkMsDCLnGjB8NZdzbD3/KFkffTPMw6bJygsRQSt5E+DVmj/NklFZuSvmm7tQ
r9wMhGGpcVgzS8ERF0gB4fU6+V22kJanNGWUAjpFZXS8AHROatakVxJcDeOFN8BI1okH89QjIo5q
KNx5RHIbrYZQdYjHH9KnlJIM+ZJU37SpzybO7cCGVWByPFkLp1do8CHyp04RD8X/Zfk2SPyJhZhG
YlaWQEMmDJgG2nMMj8+qbQn23daTo1XrK6BXcI8wUB0l85DjDK644akji74L0QqHYtEhN4ca0QFh
21bZI/qkFvnHpBv4Op9PzxcFLagy8HuyZ8Byo381aPaIOLF0XFCgyURvfGkdGz3ZgSLw8b4baYzi
kTJcF1EnvZxOLKTy22L1su/a3TRjGhqMxHcmBNMQ8hN9daQKLRIm0iNiLoke5EjPSZrrZ0ALFGru
p3H/x/7KtywYdmZl7CNTv6eR8La/oRwoZugidPABkl/bit6l5KL9AT+JAx0h8qqZ2470ItsGJDRh
wum+fVghTK85BQsty9eWZNIglqjP/eYqruvAu5SYfQ3ChTGYp/FRXs/hq23RYMAdSdqrTg7/BJrI
ek2xxxJL1EErzvLtPg0DYFKQSC5uaTmsE4hY+Xd2SawB9CLGjQ3RnKsKMaSv5mizm/zqHc6dWZe1
JIQntaPbTOJKjEh2/MyXF3lycfm8u0dDJ57Ns14nKwMC2Qg3Rs040Cch8Ylm6d9LWH1tKYRmXKiQ
OV5NQ3Pe3B0R1PTho9FAq9X7PHSVhizqxsbcojQHK+j3t30FeJBEcw3yC7U+z8nJE4Z9p21d6Fkx
guvsZmgu1sMYLM/GmFs0NJDtjr/9NlE58xuy1ZdC1p14c/58lAbsHQPY9Hlfx/kVjOFmA21WpcdR
jugn2WfaHmeQHZ1Tp4CiaXUMqs1IIAaxsYggNiqjDt/WXXNkk3yjZaTKxxk7w7eTipQWW8JEIkNm
W8RmLAzywMtQp5fkArTnMHnqPwN6WqgBzlf4CQiY2zTxY/nz4UYiQ2aj48A64QSEOv3h+ZsuzdRo
2MfIJ0XIUhKN5dEUmXSqlf49Lfy+9hNt2EwkToU6oOngVdHLIOTQHIibqjLz+EJMblYiC1yVJDiT
4A1w9F9yAVAYiu30otVZ6jcAssGDwaheQmvbIrshqmdHwehJ6dpwvxC7zSCQsPzIMTYgApLV6UWl
3DURJonP+lua8Vv/IqWcFAZnWaNy57PfwunR7z+q0TZICH2rP8EdcyYd9ZALibL0Kyats3dGie2e
FoiZ1RpEw6PfFiqN6P+uZrB879eP862c2DZ6/T6qmhB5flOLEtiLeLmW2w9w+x0vSq8nPvHjkvhG
V2BM5DoQg5g16x3+a1pRmIWuD3T3ZHrnokMalY/eikRKVeyJCb7KwV6tkZdMlLwJ4m/C7WCN8yBN
fYvw462B8YYaiNDWLTAVeek3bJVMAJkoDMFOMOUav0DLKo0a2KbQceiA2cNay6+FHL7Yc6RQY6RD
lS1dp/rQP1fWaKERfxY0md3RiW7qpCEN/1WU7TWp5m0B/F8woTkWTB6M/7JvqyWOVRqcqmSWfXFA
bRu8Jg/D/knQR55PzTPCCzUWrXZfLKdxFvOuEYfZynl4Da1MhRBs/xM7CeuYqfho6JjfHfcIyICT
nJ7VKEzVhtoQCUcY5vsLG2E6XbdIWIkyXR9Rr3vRSBnNvKNYS2e5NXkS/clQvs/Vt/i672DFtiYL
bnpBGaq01F0LEzzIkJyL6+zmsQQ8G1Grw8h8+RQsd9WoZgFEW5EiYjnsJ0gwiJIGLmYARs2PebnG
enQjPUO+xt91ykQld5OOmkQOaVQTLCEAxwQpPG+SXHtOYK1IQANswsRl1msYE46qEx5LrDGT+G9C
s2VKzFKSIhPPwPE+ppk4znurEn0fO+UQh9XLnCV7jZwMOZ77Ne3d14/guk3IDj+iFUbxATZxuqPU
0R2G7m6FX9J1Aqg7kVG88/+OtR8CuiZkSWCDyin6dL6z1UipFEmXcmA6QwoMAwfvjOoWwbNteSGF
1zZpqYMA38qY2i9MXjk+Fatdi+L3mb07jsNzgWvuc9VwsyYKSkhyZXqjj1KefmoMoJkH/dff0G40
24il7CAjeKKSnZ9QGF0YxwYtwJIZNtQnweXILpkl1UfG90OgExMYyTorURxft3Lc1SbdZX96DAjs
GnZQ/T3yqUZBl+M3R7HMf6b9P07b/7i2duxQ2MEuNyz1CYHelimw2WZCH8V6XgfOZWwhlCesvIjO
oSx4LNhRgdL0KRSHTzRDDcfnO23RpVBvprWIVDuO1ya2DI+NBO0Ry4INyrUpuDk61qFCdniXYGCN
4v4FdPf3uvz2r5td/mxACK+wITKoZijqF7s+EuDD5HL6vOKb9x0lSiXGkQTMCmpBpnEhxo0ts2mV
dkFA9hH0lVfNJ/J8f2PESWnAkke39XYFB9MCTR/AIpyytwnTmkqhs6d234tNXVzGWghu8Bo8JepP
IFpNIMRPp4HiJYWBLOUCDok5hk7Sy/v8kWCfOJO3YW1ovIgtsSu0P77A75UYHDveIM6K1nyPH+k4
SxPdDLF4Xu+rgas1p4gCLXny0aHkOqCYTfgvMUCHSLhV/3y8mQYsFHVudhH6JOHXqMPEc336ZYSQ
ZV4fbgvPXh8YzAQp9sxTmzmcsZWINDsEv5FRRYunxvcPhAxkP5tMDnB4Rv1yCXXAx+kEuJo9J4Ja
wkVRKaIboPxe3+4UAkRmWkW2pMCM9pcgnbnCFhIsmqojKD0cRSBco7ynIoYZGsZc8EWdkxX5XYbN
tFl3BuIYjjtWc8s4af5dvvQtjf0Eiy+Y35gjU2D5DvA4P/9aInsnRd6yJQngEh4Rq3vIVPTFTB0w
9pEiKSjR1g+mm/0JjTx0e+yDdHnrf85X/vQEO7dSTomgaMRwllOuFydRhl+7EEUL6wbzcL4i0vHO
E/UxzDRT7FThR0KUXVeksyurLufWCgdz7iDEkf4w/Mlbb1eef3zrVHuCdVFdT8qJ8EU0JjhFKMly
+hWVM6GzV/d1vsRb556cu6p0nL2XuNDptpeS2EF6N31hX/0L5tfXniNfmyqs2XZ87UtG4S4tkeuR
Hf4/c2e8otd3s3BXphIlu3btjVbGTyjdsEiuZBwW+8m/5UZpSEuwSio1EoRWsqddV9u/ulvOLZ/S
/ODXSkWlZR994X5g9iTPq1l18j3m5AuZce+b44LK9x0MEIXsOENUOjC5pcKKQpvAeZWXJnYZLeNq
lqMu+zFjNI3h8x+i1XXph3j/FZws9p99FZN8rH4yECZiR6G92oU6+2jSyHsp2e1DhhN7PUA/w/lE
KgUqcKWOYGisOBUSdJr/kUK3iLZ9zUPYZIfjVmX5ArYzosIUDNqUSvhRInYfIoomF/vVREkcRVPZ
yL8Jli0iq1oGOQuLIuRY9oOV3uORUTtkTna4CrNVSBPLF7ffSIb2obIwVy/hXE0Du6/i97zyj7If
U2E9oY3fw94jtVYp8DWMtiBjju96Unln+5jGZqjI3rT9aLDMvwGZLuZPVLQ3dODfntCjTMR0AkmV
3YxyRDK+4gW/wPL9uSo+lwbjRWCwW65x5NijCIgq3zKgnujSDyFxrllSAkaA+B+zB0Qmh/wwy9Q5
ouUEQcvmzDMAqm6zxePgRkSn2DfBC8Dm+qdrIPDYZssWEKJLisKDZhIstgIwUywQPXgL3/7wruH2
mXRlMyLza+6M3iPziCVjDu3N2bUaw5/zKHRwTrY++ehKunbuNmv+KKOV7luDQ87Mx78xcFHngOoB
UQ3ChpItyiRTThg3hYYNciP/HsqzOEvtBu2NOeWPjxUqyNV1qKWaaWrfZB+TfhfINBJrG7FdlZLl
Kf67kN+J/pmhuvRZvXaXmrhuWRKqL+a37qE97vQ56d9nSsXeg77MrItt5puu06QWv6QzRrl3QA8y
3UixK9jYCiybJSUVIqgveD2mHud9E4eZ/7Z2N6RGb5eqh2UoRZPJnnA54r2D6ejvHWDFKv0rWh7B
33zWuyk=
`protect end_protected
