`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
oFMhUYsqtGubJibjcC7QdOrYXy1fCrKM6JuPTwv7DqgpuwwfPHMzLPu4BprrUkGyUravnZ2K86Ls
sy5Fl34Hyf2xZR9J4ouZfV8rWjO67ZWIpOA0skT4gYt66mkSv864dPXyjatvgPx4BzeysmacNgyj
ULPGs+eMDhKeikYvclCFmysCKkblK7YsI+LyJx2AOeqt3sXuyqswD/7eIDFnDOtRBDQhTC8QtkAn
4P9omPqSYOkcHXc/KlMZ3Knggw06s5QexeAmnU4Ir2mQC4E8+Y022LoyEcBKMPfCrY7NWqw3NpvB
c2+qoF8oNHydncubnLemkPVnq5z/SEA0yKxCTw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="E1cQRtGsQuad/a1Eju6URZq4g3YJt2WgEfJseu44f3k="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9104)
`protect data_block
mrVnQ9lksAAjyXfVhCexvaGVptvmajZH1vJe8wtTSKrnAUvGl4cOJxtSk9gjA7mrfc+02hSuAXsX
rctLmpNWClPTJ0Y33/BYgIiAAVUXRH9AWlCV1WZNVJqlTMdnCSPG+NADhfWBp/WFxovyQFGX2y//
RMdYZKdC/TdzFS/yJzdrJ6ckgVY+j5L8HKHnSEi24jbkyVH2buqnyQW2eBdCOuOycbn4H+w6grfd
D0ZLpSxI0hwDiq6W48o4ceqAqS5QhoAS+YKDo2TuK/yWdZINSmH43h7A1JIj4LBtUV+yM6lbVeiE
qkGnnvDBI4lHpSO5xXOi5s5bfD1nwRjQzafYWPPkdzgFWyDJTgeCm77G7XRcEbr9MkHF1BIB8OEa
ule6ka9ri8tzWC/fNcle0A1qca+VpmBNeqK1Cptn5H6CBsyNywUY6ypbokhc24+dkIvgkI6WX7Uq
7WVzWb8RA36z5wK1DHshz/SZx59jpu9yScD666JBp1qW2pZ6+/7VnSRsSZ9Bnglk3YrMQ0/C/1i4
MoKlDOaH4+iVD5vdmcbadd/CrO/vJZhRGCeevlL3/jbMRjcnIjwNATrVZ0UwCYc9o57don7k42Np
Nhf5LdiOYclOhGbtiT7VG2MtYrKcHJHBdRYStNbWm/dzNk95TkeLsQRFq3C0OivLdbBAZglbhPSV
F2xJUYsk4xZPmhESDaCN8Z6jJkTISZlC2ZDQoMLOd5ERATH+XNOJfVrvcPGK0HpOxeJ3iwybN697
76cFZfj3A2KEGg/drEX54URd2qy1TKGV1DLa0YpeQJu3fKfk2lzAIqIEyh4mBMe7VlWR9JPnrEC/
snO/reKjAhDp17KhQSvWDn/brw/Hr6RLTVUISsPyLyMPUxCRpaU+vgHseSfBO6oUOj8RHX8I3dlT
agQnRGXna/IjkAmAM0b2YXIurE62Rrk1qGGfquaPTYKl1ghiK9DorVNSBHHVNNYD+tasTNBVKKPd
XR5KuJcIYKss2zmqZdNRuYiWWlsla6KPvHm6B6BAkTDS2sFItI5zrVQLh6aSDFk6+9Qz238ofzSn
reeAtX6uYWi9t7KrGb6xjdifIq2OkUOhDlYGV+ws2pnw0CIyzWdhcnSk/ZdMCy2eZAESrLXOfv0C
nNfPO5x/6yUX7uiOx42iprV+2lBRE5RXhYBQNOyhcp6/mJW8dEYhIBrwnGKJaPMStJRTTtPnIroE
9hn/kHTeEby6cOsEMzThELOM/P7Yxf6nPBKbOzDDR9DBKU3f3OV40U9XQ5xOVUF3ditlnJUUFvId
eXPXFHrpCVCD45P4kjXXvphM+F2a2/tAwj9TiXVyZZyLfPH7pzp98jCAct12batz23MWsA93rq+U
4DJ/NNrGZqdehzR4BhOr7M574kc2w6Vz+fvYxzwipWkSz1MPNF/2GJaYXdtEE8hQzNgBw31mex6y
QyBaFsBoKZomJoMrLZ3unDeFT5keYnhX6RiD/o4GJDP/Qrk8FNCXWr4AHN0aMZ+xoLq3TDApV400
tHzggbBXktaqquY/8pHVDIN1a5deSBZX0CtY6qdSndCZ/PRRemYUT3JEBrwfbqx24IuaYUgcHlzL
TvAt/mzfwn62QrgALcWesK+8OMCb8PXpGnu2ApdtB6MEIJKOBBGjr8WBecViKqboZWGCsW6Smd+7
ZcSv9YusgKVyUkXQrQxxTaIkVCdu/8R/y2HLZvyYBJwVEeoNb1ItgdflmH2ALfI4aDmcHzzrzg5y
jwhMBwvwagjhb/9rjq4jSEsxvpt+fiR3MzgCRWFciid1klN/p3m1GxoO8zz5IIzkiOByd4bxY0Z2
VDth+yOXWhD2JoPMSk5VKK1MYK9LnrmYQ1Xkmm3lgVahnm2qLjWCEQZ0Zr84KI5w1akpGVi1sxtx
BGktxtX8fkGLxKeY4lEFf9LjFT2hFmXLon/HBYXmrGVWBu4PKVus3Otenw9ZhkfN2q+Xqjeh1Wjq
oAkeadmS5SoojyeUxArlLNYyu4Z5lMAxT4oCkuwBdqANaTYZGsipNJjoJTTLJjD6x5H5bN1B9FN4
V9Ul9UIYoOQN4TMZGnrJ33ObjpsuKECDEtkseRQPb6PlDbu8fwl+VWRnXPyXeqh3JpuAkLehLIN+
yHJ4WT+TJqTCmLhLC3bxEPGOMkfq/N3u3c61m3FrEsgmGq6/NAzXcUwFbwf+owAlLT+u4JwlJQkf
1a7KuITOLIDZ+KgGyknX9W9DmQGPZClyvi20Rv5Lk1sOx2LhIXrwBKFdLtIp0BEIBjOuSWzjGHjE
Sbtva7UyC4TjEthyFaVdhw9TJa4lRuOWacGTIKj1GWUBGp5fb+WuxRPl1FKyegoHqRbeXqtVjjsG
2POxbcQSGnjynESdsbTx/mEe0TXl2keQy7DJUM/0UX5A0whYpbdRWjEGjQVpuYs/5immnLami+1Y
9vqqLcXRytKFopICP0JZAteGuk0nSPibPn2WF+peth8K6yXVGxZEBatN56fmXXNGmepnWDRZi5xA
cfhmTvcptg6tYlxoCJgYNeuH2aooWTfdzJtFe3DBZdJfL3O4bU99hK9MYIr3O1C/olbLGTRQhI9v
MV7aoTvDcZns529N/dxOoWQYSxhFPChErUhlHLY0ZnbT97c7Hv81RtCFiohinjadN1yxbSjrFGWD
nTdzC2K3l+Lzsl33jF+IIdaTN7ekSUs3ITHQEBBEFG7gRmbPYmpm21Rz1w9rATlssV60XPnyJJzq
kB0zk+g6fbWr/VXU6kMBkUWJ+7qTxj7XeHyFWmHKh2tgdjKVY7M+s3SJ3xUzKIIi6L+ju99vxLj6
oMTmn866Y1rs2JKSZIBuxpjuyAaQPoeX3wSX3gKg/fdBagYOUL1mmYezMc1KvyOoMW8MV+CAvwak
BUQlKwXn65UehAgNX/Vc7E4O5FZa4MQHzKh8CCUVz/zN9MVBSHk7CfpRo4BhmXsttnW0BZeXO0k1
oizqjj6Jc333GGDJ1YRBuT/wdIclR11c4xtY5+Vsp7jajHJsZosTWVFLGoPMl4hfxLdiWSHsnES6
ihOPv1RryHG/U4Y7+rYKlbBd+igEXbMjtR96eT6GcuhTmHvbek06+ceovMEyFEMTg2P7WglilA3v
4nNxkTQ9+iuhDE79yT6w8oi1fW9n0qyCHbp9mLISTd6EzLpCloozjAvT2KDif1ykpXPygqhktLeL
ZuXpk8NZWIZBIUSRSE0ZqVtYtw7YwG6PV2koLmOLBcKPZz0YsOFjUB1bV0VHuKe1iBvparwR01po
X8G/FEOkk9wBmhh2QTYs0RqDCfTT4fLtkDl253DfaHsEgAYZ0eSgYYtDyIqPmzdGfBeuXORq0/3M
hRWDava0W/s3+JZ8kKhEUtaQ8jrrdMK5zfQr69Dgz5zTcXUiqwN0cVTXHciVBYc5L0tzmWKQ/6EK
l9xTLmkgiQMo1VyVh/MsOw8t3AqKwoIDqespAFVbze5YszcoZnVG85Tknky2WZbDxTlWENLyGBDP
+rsaS7kYHt4GwfPDC/2qO5gZbv33cmGLbcJUa6Vfr0rklW3ys6WYEr+dcwZD/c0sPYqrs9c12BZt
YpW5pu/Jr1Pc4yW/9E1KqNYBtGuw5nujDD+0EW+VK4mc9cHQSJvemxpjyIVwqU3w///TugnO9Mh8
OhnbBM2EjR41uGW2yeRiJDebaC6dHCoFaTMsAWU9KSyX9cwrgoTrOjtNAA4HS+UPD9H2+r5C8rd/
7Pb8RCa7epijnveU4FirpRD7ZlYZpT/j7wbdjPeJrwvXVbm0tge33B7/N/wDZj30o8EfSbc4zyet
x3uMXotGzzgTLLjlxWXLDRBs1mZRMM2wvCSuAf2xzqs5aGbOE4S6lcbm5gxAoV7qvew8L+FKKbZg
dXRbGWy+CK3VNlOriDC2wecyzouNILOR4lLic5WkwdfARYEZlLpJ9v/4kcTRsPNoigA1LRVAAIls
/65nbhuFiceQlLEA4cirXLQ+2TN3xKn3F3XM8QC7SrQ9xfYZpF4XZrW22LduDTxjItFJLH3vbeqX
ANVVa9mPGZ2L3Lz9ub/zKgiVF7liHz+3c1kjLNMic3JbcYBhjECytMRVHJYmtRl/wNZ0T/8iLmzz
PHNRDN/9T4bBES8KhBh3VOmyZsuXNfsUgx0RyFvNk4xvgn5ZIJV43iOP1GL8KSvRtF4hOVwQCCBA
g6qb+DM0r0gCTuX9rNk2hX8W4vuGsC+1Xkbv6wDAAf46MymiOm1LwBmtj5jBTF3bcnWEvRggw828
MTxTzi/BVG477Vy7JHreowBeUklCqedrNqd0xGBvgSesThg9/UBq7vMDfEl+m2b/FHax3TmA54fp
wzskvqEcmx9cdVD/puF0ihaTFlOV3qrX0/UdXfsM3YClPaa8VNlShR5s7+Spe6uY04Oj0tpPWNjR
ZX01Tk2+KlgMFlS4kHvCMyzaIRwu2DxcbppyJ8tJGlwd/ctWsXW6LJ6TvMvACI3aMGPl9+E+PS61
hCDfTLlth8QKBzoo5/5JGckpuqqNzsifY5QOx27DoPu2k4zee/vN/5K3Kp17OxqxU69bpjO5JdLS
xVyGGGg3qbWIXYgWe7WAmCfPLDQ1ComhOn8rgeD3jDHHefHHOjr93bXWtrWCgzWGOfmcTCE/h6+9
Lvv2qkOIw5vTg3Ugw73cLXkDMSQ9iiEZFqaTBiobZVL5kpR4YQTTX7nwA9+JG3T5dszzHc/G6nPo
jQPzJ0E25J/5FCElaoAJQenrX46f/kM2pSjJ5rl9cCzZO+FdKiPDOCnufmqZp55Z5cs5ijITjqx1
j6nv/iDrsh+z+EFDrn6WXFKFgg0VxuaI5QN9tDcQLVGqbJfS2FzNqYYmgMfvYz/Y7+5IyRYqVEl/
6w8W75Q70LNBIkGQQrbZSotHm2Ox9iDwANO5LtPYW1LaZgR8vGTTZjZO5rCMcRDs7iUnhuPXMHux
YaMHVEwrCTNwqi/CNsXS+UwNi4bfLPCF78MD/TUJi7Wgo7UyOYwkGQT78tKNAJ/ChDnGVJTR1MIU
kioP7oLMpUZT9IxbRLH+BCpUKhyNpyB93hNaubj7MAFDFkMnKiZmZWEIkjAysxQ950QF8+3SKvrH
oDVrO/tfFiGowD6MBOBUpO/MMxRb1O0BOhSEBL+8w6QpmLSVigSSRnYYaSMACgudtyAn6hrDkow+
bhiTG8Dksppu3oJA7nMtWXeLxnPMg8pEI4lQWnGYTM9aLe77iaOCYbhy/Sdfev+cjq4CrR5UyxeJ
DXCE/LGzUOeSdRB4GTD9vAztOMpPizOM7nebJitNIwpZxFzm0y33HEh1jSg3exyhQN5YG7CXKcx3
0Ve0dSstMoq8Vsz2iBo5Wn+h0oyekVQyfQXFXH+k5qjfdV5hd4WWUg3sUa34AzNooXufnUBMw3SE
KPQZDuaIeQNRszd5ecYUIIUNptmU2tTi8JMFtDeEvDX9bMb4/I/nUny2lnomzXdqi3PFqGUydzBf
BbJBo2KE7PguNFx05MhwWdvGJe8E0wK2Kan3dS1h7BjmV7MH6W2VNTWkJS2wrYW3wKIdLbuqX/mU
u0CExOu/8rAM/FcCK6hIQqdJQpmyvUK7WOdAh5OYLHId4Db3WUTImq+48v/pWhcRqlb6kJGkB1MB
myemvT/E0O3+0yNb/1c5108dCJqbtkyDmOMHYkwzYPD/34wjGUdOtSJa4zJirq0VddiMo4PQ0usu
XnShyEsV0IgQFbUlcGURl+hH7jXIp0GImf3kaTq83TjtTkrtOHkaS4pcKHEdFTqoUt25bg4SXR9U
U34+QLhG00kFheFNtggiA3gmQvoG3D0kfR2QdikMOgS5fsu2gerj25Jo35tHyVYtdU+eO4D/Mt4a
2Xw1/MJpXYMs6RNnUGoER5QbidfqCtl2g9uupGu1ePR7h349es9t2fxTgJ/OwEecVnG9QGtyKqEX
PoKiqZzAJqNrHbqiHt4zAG5iJMLEGLhOHa9m0+K1TDybp4FuTf3ejc21jRQND0Edy2lbW0X5RySo
SoZYh8oZl3uDlgnsH+uIRjgxnfIHXNdWpyiT55lxuCNJbZA3D3jeTMTuBRhv2T2x1A5I1ME208gh
Lsxg3uqb7ClGuAN3ifRkyRCh+Llueq+adayPgw8nmuFfp8GzJpQo7HPh55uYf12ws2V5u6ZS9VCw
kMRVCbtRRqKl7yuuKNvlDja2OGnO/DFQkBtyOkgLVLgMdhiP35wD2+zIHfA8LMH0HoNFRg+k1DBX
yZ8GT6dLI10F8tlLE6Zq1/OYAJp2ymElsxugunayK9P5ycacqyQAZvTcwMlaUI4nkMli0w/WfqFD
iKBWSOGgWgB4+/vyzqLItyuAORa5xTefLHoPoU34qU1JKwCwEMJrzYPI3OOlES2MFVFZiKrvNxCS
4bCk0F/H7FHd+15EgB8itbzyCuLw2W9dnpfyozWeej2DxuvBxcEgAgL1vjvR0xA2z8VZOOaGTky4
xiwVjZgLe5enaxP8WuZqzi0zZBqHYhjeEeLUXE5rzHrK1+oJb88gBYuZ+CXy60LUaDYmnnmtwH7U
mPa5c8aQIof0f+uk12cJdK/56r1xBdN4ZBdCE3N/hNc/ia1EWbt/fQDjng5ybCf2B7d1OfwQMSvi
gln2aCOHL00dEEPqKaUapmdDX9AYIJ4vtkAzJ+sibenvj4pC108Gl6J/PHeqEN9H/d2f/o6FQLlJ
/TFzcU+krRkXe4Cdg9d5Phlh+Hf/M7ExdXBCCDNZT4cSt7SiPHZuhUoBep4cJ4cTwQom4jv3zd7E
Q/f+R1vt2arsZ50Qz63xbs1HcNXHVC7QhutyqEDkIClVKQlz9tL5lbgCVyEXPaO30EqlWZSz8hBt
Ug385JIiDxw2cfin6/6tS0eAAyhLMZK7WpM/tqEIf39NZ6JQcTQ9GRrSbXGD2YKUvnR9hIQIHbu0
2cYqOsbgKXqPw5a0PUhMus2mffSccuH6Dl9FfZ3TWshEp4YIn3XxCwP3DPzCB67uXum3WYWr+l6G
3cJTWFIfatENta3W2500gKL1CkqXS3YV3/XvCCCRYL3cH7JeuV6GFkbOtK2klR55xWbFl45VdWyO
z8TSuYYPNbzYEWZjd+wi7LPZ5lUG3WwGAK8X/8dZeIhaqJZKo+wk+FzXtJlGryBIIn6Y5EH0ehXB
/lEN2gJLGci4tF9Avn/aZ7QNdVoe0IUNj0t0xps5QpvO+kEPUos02ttvBMT6Wi2OOeuc/GVIXUxg
qeP+AKfZL/Ji5AtEbs2LUU4o65Ydcu0pAQQ5VDEO26Bfb0ONiTfLQnSzaiENUpBBazZAI3BSq6Kp
ZCkQDQKdoSjhznt3Z8cEprzwr+Zu7ChbF61RF3L8275JQg8c/TVVh/MwNIqmYXWTnev047nvvf+J
CtKr9YFad4fN6RtUJMYKYuPNyvvajFfZPOiuH9GvoiE3b70iXilcZtOd6pk56sKlKKOdcfBHUlIa
xQuKuuif1B9mQbvx947QOAxTKuPKsxo5fUJQp31aGH/3/iCeOjwcuRjitn86oCCDPPl129gsChLM
5HMhHxnFlrB8CgUEfp4V5VFSM0uwzchz71+JSics/5nwSjpwokdg4esuVfo/xz2Qpz0tBAWwL707
VoFZsAp3DcXfqXPtjNSWmwen5CTmYyylTVlw9e1e6qzmZt9Oo95aby/5PlBhlVHoA53/WKSw2nTo
SDmVMjY/hSX0n9luOApZW2QHojRPmhqArw3Gpuj+Ib0CP0Tfs/sYGbUB1U0OkEkTDEk6vuu6OeCC
c1gg/fYpaCe7+t/g1EAHy/AHR/4x71jAACmn5nKy89736zgl9f8yiQkW5PtMIdLAbzQOO2Pb/8BT
r47R/SDpzPTKbHBFOgGlezF0EKkUrIyzye2pUTXnQXyUjTbme/+1oYIw91NxKFbX8AuFotuNwMCg
El5dG7B6JiM+hrp3q0T4XrVJGIrDGluh1fPh9GkX81poBK7suPufTVq09DkGKUMBsorV66JtxnQu
UeDBdk7ZG3BhenLNZwJpCjFYqJnBEdhQoUV4ZHqyt1TrUAvqbficreymF0fLZm07h82k2tf++NN6
7SPuZDeugw6Fi/2m/PxYdsANyxOd/Cu+lg3fUmROvtnl+Gj53224qbmRwJhiJLMJpMLbUxUN3QjR
0OiKG/J2D547vbziRuA3IdY6vSkYXy18Pz0GNKwqgssm/rDfu3p4kRgwLKKIhWg2QQEqCJWQiKrs
bH9IORYAzfP2yry9aXS+FveAhSOLtrdy+xtU/783RjoOyG/BUO1FPbnTQHggaQ7OhJYIoL5pLv72
uYF5+bw6BTxi5VWBtreQeaYA2HuoNTXVspMCZlxcs63RqIJUS5ee2P0U6kJfD3Z/6ztCyMqJdhuv
txvc5nC1rfQL8BMVQlMVeR9Cojm1a+TBmWyYORHlY55EazmHQYjpRqsDFGAQdgdnwTBuC6zIspxF
iyAf2vYzoPIaRveN2QbIQQh4RnYMleA/u7tTusXIx9jcRLiksOleejUBhxSp9PGYohP6daArJvu7
lW4jNrf3ORGZbSgCT/ONwJCOVzhyqGvA1jsgIz+L6JKmRRjRTnbw+dtfORcbgLOx7/fRabCAj5LC
pXaGWfr9nzAky97P885VkyPKAAV64r6SzGNj19+Qx9s5oC7/aXYJkwSnIovslzLZJERLPs074TJE
DFigKmPLlShjN7Jfgolu/pqBMUs8eA+UiNwrQ+9BPiB6/PdrGpBtrNrm7GDv4ksf5Bc9rn03wcb1
7/H8BgERSUvXCHJcVuQGUfZTTHpDCZhCNyXpjmToadWOsE0K/Zscv1HF+n+OVI2egtwTCGT70hgp
HJpljlEuo4+yED+n5vU/EE794nWzhqwM6qftN7SgRqHVzpczmLHr1vnzn6rp4xSuHGwlxvp1JLQn
bpemfj5LYzXIDx0mIxCJRotMGApjGAX0L+D1Sznk1XSi0JRqKMF3nlWlODoBo2VC3GqhLwkfvBK2
Ysrvirx/Tphe4aJJyziztecPt+tSIk1v9aEj9P7UdNai2vfFvuh0PRQvQLsR9ZZK4ouoxLyKPk7J
6gl58g0Ij+nEPO52wfv+Xz9RzrC11kJ7f9mUNyZ/wdhFvF+5y3ykvVnbSfFLeox1lKb90dw2U0bn
zsoLZyiSe0k5r7QA6zQmKOBvzBtHpDfnTA58NH4Ox/7dtmKGUiJVXd6Yq97ftjzDGIgR86db9EME
/1jXqeW2AH36aFlkG/GDJflucFirKyR+0U531asRjJ2zLMYABA1egMrAZQGxWSGjF21Y9QSHVL5V
ScSgcAr6raQbldB3ablcv1DsuVyfmjVi7RhEK8zcjcSl5Hl2LKpRDNraRm3FwbuK7ke9Cek5gEJi
mN4T1LI0rYlaVbuglpK66Y4si8MEzGJO3fxG9o6evJQ1/OJNM2YoLIb0gcc9azbj7sRKyOVwFRZC
0eESPIDh4ys4XTJ1EKXOdxkJLKWDSmvFflWVWeOnahnlbBqUWUDwj9tGyUD41A1dqJWy2Gs7IxvH
vfiTVWNLX3EPWTSFiy4XsWxZVrm4qEUemloBDjT8QvkPaUWKiY3C0woOxUcF21fg0DxFi69dZFB6
aWxlUeXPpmK/oBQSDORr8+xTsWkSlmhSV/FKpHZ7rgT9TOD38+f898olTzpSUa9Jezp+zE1PIcwl
uxtHF/VMctCzaUc6oTY0BFMjUBveCjnKxBQKQVefWcexsMKw3El6yi8lzZEMWkEGMd18waLAQNK8
yJtIJFl/4h7cZ6WsPQIDd1wmdrOEbhq/jLuvn0E6JRNpQiEZyZZERYdMSryS/V+nOTFANcbxQW79
Bq+IYBprmnAiFfvap253E9Um+OxObpGVj4QB8S2yAzhM1vN5u+JRrnKCx34lmpfJeGomFFinQwBI
oj/ERcTiofBU1OD4AUSqrVJtDjn5dNEPe/VEzqOu3r7EBTtVLDAKsUUGuJN0tUFxltQxTo0CfWhB
TF6wmU03sJKAMAxaSLPypx08ohlGQRqj/7L5Go4i/VdhEZZBydUk75dDhMNp+FgjYkOB3AjhRhMj
Z/DUEXH33+xE2w2fFikkduxH1+e5Mmwuws+aJ9t3KjufPoxQ9c0B0rvwwBnIVrsftymT5xQRsu0P
9R1aAAagNHFdhMIh5Fo2x1CiGjQU6b7DksJWDfc5sM4e3WR0vYy/OevyZOP79EjnD5C/ICkYgp/s
V/vAGfTTYQkrOiz2dHYgFXNcbvXjxIMYS8p37sM4FNCL4hhkaoyu1mMPP4aZh0tLwQPrXvW5tw82
xnjakMrWV/cRk+c+OT4i6OHWfPXos/akWLaBhO0GPTDcUVQVku9K7kcgXwJTfiYDChnbm5apXxtb
4BRwf1fIxCRkutAKZu96Ya2F8ZWHM68sdK717nd6R96L+j9QI3ffSIl2YeiB8wEZosIaN48muTs4
6JliIWpZ0F42KtRX8HYbWZ+nQ/mYY7ngP3uVPx0Bi5naeQLcx22k7vTZ5z1wgN6+Ah5dZOovz6o8
EhqBUeD4JKt0rgrjsawFcI5EH69vGLvfxYsSs/iZPt7hJWOmXXD8i8KjJZte5ZXqv0l75N4ez/1v
mbUg9V2V6GAPXsLFEOe0LbO4cNcVzhs3bKd/Ws8y2ZsOMYZlcbtuV7QgcI3syNvos5i2ppJvR0ai
vDFYXm5H6tORlPjuaDTFtVpmz4vrMQZAOrloi+aeETggFx9GZoMHuShkZEhzWPDDFj39FaWPT48L
mCypTuiWx3LxHqp3HCsokCceSVb0HAI5LqjtmdlkWRy9pImdGsIofyVBS7b9d7qaC8FssFW4Z+b5
ZHj67pTiL93sm5k7LR6z8RgFBuH4lve9hiEGgWA/qqtpspl3yaxp3V0ijSSCc8kRmIV/q5dGm3lH
f6mNgrBLNneXPxNpCDy8YGPwmHAYUSILyxEKK0bk+cgmRZIS7xVAxN5eVe8/9fVaUu4jP2VuObgm
u8qUdicROMh4wHMqRsfF6tUq+fG1xucLqDdEHoZNaA+Lv7wLg+OM2a15TqfzCCm3qSa1k+TI5xN1
bbZOIM0KkSSzCD1ljVH5O+W8ETJtEPDlNI1JKDxckXFNjxyjv8MbYRu3YMBh3dKEchQm2ObVLOST
MJHm/WR/Ajc1Qb7grU4ZbW/mJ4kAcsFQFxKnlWdxzHmhGxM+o0t2Os3Nj7u8ZAlgWAfUV7+fydDc
vKe4xg3ENt2X0a6PoMBxpGNyR6Rkk7/1Ss/rDY7vR2T7C3f/9A5Am5S98RqtsHbN4hYo2eRx6+zJ
CZJgAM+ruxKOygDxSmtufYlNVFlJQ9Jywf2OE9GOlilRx4m17E2ys2c9Yeuh547CDu46fbnc8Elt
eVq87BIQki3W6Fj1qYif/xxyV5UDR4uPGM1I8JeHiLo8e3/RAYCNELx1/Ir6HMGG03pfHL31JZQT
Ov8n4mNRbiSqmJzMdfDAcNEp+wps38790JbT6c5GMr0TCSXjPZ+4A0AlOYcTrS8XUmzvtWrNsDGI
b50Ouv8X/3eLDxZAEJ8Zdq5UNiF7bMp7mfwVSJKrq2Nx02ZAANPa6g6R7RCg1nKNVEutk48ycjk6
VAYVpCsmbeQ2oWIk2+JzrN1GpRiwETFgIhrxNbhfeIcItVa69ktmwNA6xCBTPDPTPJz122/hraFr
GLqrhOQTWDOPYn5NvMsTfc/QZzf3i/1dOmAoNwZeHD1blbjbwQ4pMyPYarw1R2kMi3gJfAh/frJn
COxO93zk1WwxBGsl63NMW0nCsJwyf1IjYNXx2RaSiOLGNsQhu6eNVnmoXuSudRccj97vCn01Be+l
kpd0h76GC4vWa0Y34fzmzTKHDOImT+x1y2auElyrs5oA8EzkdEsSwjylS/dPmax6QKXS+tFebfSk
khKdns9YXazUVVnKk1B9lt5Y5bJhg3jXkdQbLHjMNb1iqb/7Dv40FO5S1+zFyyj6eSmE/4r7PRnC
LYdZhK2j9B3gJA4S1qZLoGVtMgVtNw6dJ3fPq725v1Ij4TbFTe3DPoMtq/9iAhuaGXXqbY6rQs97
nV0RDIg3tHU6Y2eiYO+/zJuD0TgZR7gVpI9gkjVgtS3Cc+FvOowzu33jMswkDdW1tqEKEH8FncB2
2B6fVjO18TbcKsj4EpOKaoSxMC0flZADtQaI1hlKFDhb7W8NAaFhxCo=
`protect end_protected
