`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
OR6r3PNyn4n9iyZiro23Lh1jA5iaeFp7rjarAQ1kM4kMLAvXffvhoGOlvaesEbqUMzqrK+JGliXg
Id4UqL8DMUSJPtR19obQuln2IDfbbHOFbetddWXoJaXUtNmjJioCgkM/TSsMj3Xl66VZ0/L9G1j+
0UW9fwP0GNAhX0ygzBIjSwb2R0rM1P1aRkvH7wTTtOIt4be64fyZLVXWCqH4phwJU4gQ2cphtVDI
lxwCbJXT0l7YAay88fYF9VFNlWd9AhI2yYZce2Fa1s7TBRmc880mtupYCL4WJXN+F0F0X2igHWyt
RiVnU1TqO3nFMmeAYp7po075NPB1+WSoQ5vaRw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="zXHiLNpVh4SAO7JRyxUbSw43dJm0kHgKdrdOqhbDwr8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37488)
`protect data_block
/ndINdYdFvinalfLAwSXe42SPSk8nt7sxUepL8IFizlLi88LJGQNFQZnNbpqbCuFTtuFV2z6n+wS
x+bqLDVHs1hl8wl6VMh6fIK/j9jte/J/u6JfyhH/t0FColQxzr9EeHX5x+FEL2CtPIgwjsN1eSqA
xS63zRhiauUcQ8EdCacmeS/aztRgUU0A+NAenzazF9yW+qmV6H2yuzwyKkNgjBkWUVSRXlpXiu1s
+9Dk+tiq1u0KE/Le9ZDfo3gKBlEf1gKwPEN+bxfpKHkpC5uheWDo/Q+7WSw810CIM2leDNpu3qKS
ZfHZkYhmSl3/Ngcl49lcSpbukypYJNbP2V9yBkVcBAv+fK1gp/Fasa7wKCSz2OmLoiFfI9aVKzCU
cQunoTKl25pCEtiasFaJBW4qJX+lyk968lK1s0xDRXzAZcnDbuuG3H6lexi4+DaXSCR8IFmteGOw
4pNlYFnPyCAnSani3jUwsRhu0oCUTn2xh8mU5bvit5tGXS8iUoko/aSYzsdXtIA49OEsGgaA1e/X
hjEG1cKJcVxBYMPX/lRpvclFRInbJTnkwy4KyxQcl54aYhtIg27z7eonhUZDjTxMHVUCAILDftEE
zaXwVjPNh4CuZNsiLa3hHanrMuG0rYGRkIZln0PHVUhATKxKDq6t0ZxjP3c8bwg05K5apeI/TvuX
+67AsnYY9/KTDuWyvp1e+dm2z7x0GfXzy1EFHFXD6Pnic+84shPgWblt23Lpi51zkYUxmrenePNk
SicNMWyFCQNQ3rt2cfBzo/0Z1NRe/r1VJac5HVGOAsVKUQvLQEcGOymA0QX3PRTGv7SK0XeKa4BK
u3+4oG9wW2jweblwPUk7ovWgNncXX2lmeApACu8GvQrtC9hNlTz3TKJf6AlPfV+X2QDF6YoDlT3p
3N4W2XYNgxO/woXsr3KqHU5sJXvmyorQ1R6XINGEQVVfcSk365u6dbGrlRdZSTnS4dXHM0wJt7ya
mVl8hDZ/iydGqGFb/9Ahs7u40e0biQQrbymkBHk08rporu1ygWJqdF/PaDYUlCtgRYvQOGB2b7qk
cByDm0xEkLQ/AtJf994qUXi22/1zTBoyk5iX9X3K4sLt64ZE8D5aNYgeUhXR4aTC4nVn1uNfl8ZU
tZapfn21MvYdV3bCqdJPTBSLaCSYK3arBrvqSy50s+CRFYJv8FZKFM1PsYUKWj6a8qJ4OlXdhvL9
EbRBGoW3wWutdzobUgWf41igy36FzzVnpGQRPFvNlrN/Dk8nyT/+hz29aAYB8ZJ7UVm+0qFv/z/5
68NCtjH35ezEvhOkpm715oN6isksqm/amKyJn7z8MToMsfhYp4++N1nyde48fbP4g0tqa4KtrE6k
d1GOSYxBSz4Mb+Tcll4mAqi9uV6PpFTYH6hl1t2EyR5iCt5LpYirOoGhunptj2urpv2flNoAEJwo
W6IWSyCKWTNSPKwfuZrzEeGsgb34BVtnP/KiN8+3fRryViX4NJR8A43yy3SWiDbnrJ5RRCznBQEj
KLSalvjs8RqCpbcgAhsMvMCSyf+3x9ZHydA+Z8+ubTWI9cUngpypKb4uGywgV2hMzfJNZjZgsmEo
lx7kw6JtVgUQX551vxxfkS+UY7EIoxtKYHAedd+aR8+DEAKHRDtjJbdHZKHddZVqFGSAWuk73v9Q
O4vqxhA1dSppG85PXy/0ipMsF0nz1fX0k48YKTlZ++c1L2hEfRWHpp+KkwkBo0VMLrl72RF9yxxY
RlMnAq0szfwwe43X5V3a/8p4d7CwrrQc/Y2LbEkvxOeW7UHanZ+Ph6nZP8mKfID7Zwrf6zTdOz/p
iB0fx3Rjx6zb9SzWtw30JzWugwcb5MsP2QHpao1lc3+68EFb/DgSTIEbiUTlkrzhQVyEqVLhUte8
hwAxlEHMbwqwHmPu45nfV2wl21iFi8btHOCZBJQhfOGrF6PUcu72K31nS9zygDvgIM6L/8O7EN3d
HxpC679hcsKFOaenKelDWEtonuV54JyrHcDd4xi7qNuW325EoDPvwOTL1pKoPlbg+5FiGuxRwNck
p6gor6gVEPwNLlmeJt33QOuinDiN8NAgUWB58dDkXg4dEBCQHhovXf3tbhhBA6r9yIvNsSmzdBCU
+wqLnFCVhlE/8MzLe/mW0luR3V1GbAGdFX67vS23HBKqROpmwzFG+VOsC4A2cjU1gTsPjkKUWrAV
jSmYUGYPMJJj7UO5dxY4/AfBCiKK474Zkh93wMg+CQoKVgG5tm1+IKjR3iBOAvZv1LxkodM6tPwZ
6Ba+kXreJhZidBMRDYKhmu1Wj+XI9t6aV3+NaULMLD/debjeA6ypeqWmEPOKirQc8ssff0NVcNcG
q3h4b28DD4e+IUTrjTgdFQXYrKcJFxyfq/yTBxCt+xGLsahKhdijjxNp0872FUTZo9ynRNlcTZcx
BNThSOTvVj6aJhA3ZyX6DTmi/GTC+124n/swHOOOwpowS1nGxHB2SEtGrZhqnM2v2DNzh4VXxwCN
BSMjwemGC84T+xn3/Jbwv4L6H/2snC0ydLR2sRGhAbV3dEqTjvWXSIod5SrZu8wGQF2huNJIvkkv
S5I/tlju0jeR9/OrwdAYUYiJjq8R9YN1YEvdukltDLbDnJDQlgeGdJX+sBZ62+T+yH39fdXjzQhf
paIsMb4lVRcCEx8g/pB7ZY4RvuxR8DMJxeJvoqIPc0YJg/wqOkqzlExnTug2iOym5JHs4jpgIhRp
wtbPM1izhnGtqnW6lX5S0cJX1rtZFhHPjCeUGb0FKwB/MFGnmclCVv1NxaF6YuYM2vF0d1IvJsEF
8Gm6AVoqCwWXaKoVyfvCnHZ5Ql1XhQfIj8g2vTG6+ze3Kqi7nOIkv7GF9wXKhY7QEehCCxqAROdl
kYiP5oUYmD34OtrvmcvDr3JDHfVWqwe0/DFURx92AXRNaf+J9e0y60owVcQdTmzn+Yy0jWvwtlPW
yHy0H2cGAll/xz8qy7KtWKpuLEBIQh9QIfiDZYAqd+R2DsFMTjY9raEbz5LQLAsZjh2zORe/xQwd
2svTHkcb4EN2/+8SBxT8DYtC6oEkJKDA1hLLjV5MScZ2qBdlkCwLOvGxcyaWydyHrCY/4XnCZnP2
drwXbHRC+c3V4Kglx12ZcxnEJCx6qwXLDCog/6oHdLk/7boIUyi0UHczP2SBSfE8HHng+VwNUrSq
7hFgy2UXjXZHqYOO6c2sdqdZJxzTewTo3UKwT/YxcryK66YCk0NTQBb16+b0Z2Buaml08lOsOhm4
VDlcH2unVF70EOh4QRpgMUtdF9/mnSVxcujpUDIy2PKxPINqWGm0ysd86JNaohEtgsUl63EFy2A0
jh6AQ9YS7/WjNkwbGNP2AB6ImzVHaxve3g0fulRDGR9CVyMHFwN7cwGeQAsOzOxvm0AZ+e7vLu2o
b1u9aTyHOUH1t4qkltHxCKxZEznU91gtUhzqhPLOQKDQSXKqXOEeGz2tT2E6EAwQbd/36NE+lVee
FCbi3KXVtJecwyM7agTnRM7ozEv3E7IkOUXtxZLsF/DNlwBuRlUhfCl8uNdUz9nGqqWIoWPvf6Rr
5DQefzxEfUDrjpxP3aVqgoW7VFmbB73DD2YhrQfArbGay5IbNgNNusSVH77GrWSN6qffjTlh6Z9E
f7Y1E2OJMpN+b2Wk2Tt3Gz57mKu4IWaQBIhP3u05RX/XpzmKBYHa/hUJ5rpNfRNlz8U7nS385on+
/UDxgWVUZpzr+ryRdc9A1K+T/LMhXVCCxbW3Fp8ij9rpGUy7EsnTjY8xqp7OYKC1FoYIVkcADiMb
yUnnsufWUVon9+vbuU5bzFFDEbS3wkM1ygUA0FmJu0W4jOu17OsnpykDPAibzDx/+bUmWJU2OrrC
SZTVi7rBibuhPA8FTtqMnF1K+8bnmwM143brZiAz72abB4VNhNdr/XiJZBuADL7euQR0edNbxXea
6ykYKvfuyEWxDi961BPlxsOpCyD0TfBkJsU7fsosNDfKw8o8Gqx2/Bbe4aTX90eLFj8+yLPUUMY8
/DD2jUJ5gz5H+MngfSYHJn3doQlaTh6KeDYCk7Fn7xqtvJgydg6vKXWd84AOtZi5kuHjRDFDBIHM
ajcn9nO7XD8cnoOLerxtZGmMumc7zHorNZ8+YGaWh+Z3mq6un99MM9WhDjstg03ORIU1pidBrGvq
6BGdehlsByQIh0khCi9nUqSqqKIPibAERo9fzye9cYcZgMxli9YAi2sYPHFc/kg4kFge9LEPJFaL
Sxruww1/QLgxCdHG+P8Vwei3tEf+Sc0rSxCOEo7PqMkSWroaDtKB8MQ5dCmJPTpEWb0AsyhB6mP4
o4C661OfA4IFw1JNF/Gce0QC8V751mnkAWBClUnlRrVhG1+CofbPIOujmTn4CjSV3OcqZmWGAY+V
Xp4ocFb4yJFSR0PWSJs1vRURIMRICEqB2+vrmTC8ptzRYX91Q1n8EgqTQi0HvJKF2VLh9UZMHBeO
fXhieBYOjCTZH3bTCDu33KReSlEczVZqjfR9jxavCXd06/0NUrtozzde50BklbaAsfeK58zfEdac
6OaJ156KtW393Z/LFV2Q0ojyyJkIZVSbnONbLKJb3k2zgngSda0AkXGffxCK//sHWLH6jK69f38M
eUCAWvxFBZykWo04IorHoCJ4/lqk+ysfpaqClr3jdKCH8O8bbnW1bYauCI8rCMzHKFuBUkixuJww
dnysvX+gGWbHv9P4VEllcRkUv3+SQ9V6dEdYgaLzunokS+bhIrprwte8iPQmkZv8XrM3HTopJIAo
FBq0TuH8xz5mXnlRQOb2rE01ig5XkSqlWPZVckCgysjaI6r4v44jr+RcE2RU0cLsCgS1zr1lp5yL
2+IhWeCnjKJyiYKlKM1Ol/dpuK0tvL7WLkct8+mvbMX2Wfw2fzkeVIvshYQr3dGGb1qs2Lk22Z/k
i+1hcsnswHOpFqhKqh+rZwY9vGRFxYgFf5jclllOADnLlfUEjMsuKwwPLvuR9ouwcRFHHgDTIoPd
vACkFq4l26d0mlgN6g1E3NOdRCGYpXwoc2StdOyKy749gm45m2gFnOrhm0eyYe2+K/BfwgmSgEMS
5n3bjwDEqy0BwgyxRvRn2Pq2W+Sc3cHnsfWmHx2rwKWh4FqrjmFjlkpwrOoww43y6BFMWfyGLv6R
w0Y56U5vA1rJtiFJNjHpD2K5NAtXUk1xEn8p1x9C+aJnegqWODCX74PJFOzyj3Y8btnN+tAmL7sB
2TO2Si9RyXjPYfhiEw9GW+2A9J2+fvecf2R0QXfrEVIc1HNZ9JkujsjtUpgm8i1OiRkImex87o4t
kUnoBsBDjuBiWBigleTIiIY5J5hYDm8sxyU2D0cyoHkcRzsqlC211nlKM5v8GIQMY8dks5xb/HwV
zoxXUCkNE7wIrBnkcPUOr+rQkSIe+zHTjPA5j2eUraXDoysOdU4U/iKnHsDh/r407pYMDPnI5FWC
FTqGacy01ALvefcmdEekcnwGwiW0SBUQzTlD2xmW+I20wuaU4I430panvTASI2gIDIVdWKx2Kmj3
XO201fh8LG7XA0A7CAEZqQKa2LAy5lc4RTqLtTrvivSySHSdoG5f/RFynuq5wui5N2SazBRiFqZA
BbxcAh6R2hEPDsOVSh+hCJIxsM84mdxlXx78Nbfa3ImfZSPJ+MLH9OivssZSvEszIEVlZHwZjFrz
Pn8vXM2gCoDYL39isg8/TW474oZQp/HXFjavKwfVgu+fhXoUFTt1/d/+qDm+YtsuDHVXwgpC+Odr
oZ9rIalLtf57+VwkMa27k3OHc0oCT3MThsxbUcErz37wPeuAiaiz9ShWyuY9wvBpnAC8yAswbApR
37SAW2I+kQFbqtFA1iZKnOAnsf6djtQcRMeFhttfMaHSsk4KgwhVUFYyY0setCT/N4YdTYjlVHH6
anaJFvZy30n3NXM+8UMeBqxU+pyMtEoOGKNGShyLXw9K09N2V2atbwlVt9cARmF4Zb8zLRR7x/65
d3bi7eymd0XRLtt2Vj6AEjSYxDVGMiiiEpGjogx/BJzjRmo89vU7RZi9IJFzWiIodmRCpWy4gAeh
UpAndE5seMAHVMi3Z0c//1ZeFiBpLqVmZHgRDzVc/MtvfTdF/cY1NQuhNff1JAFdZe0J+XtwF/GR
hIpi7YrdsFMYGn2cjXX2zP6zNxL+RUIHHoKhPZHYI9RyF7Ifos5Bfr6K9JAoVCmV0+/KlwahjY02
4gQAeoVpefAJN0/I3UVyN5E8+bFhjNaLKzq86A3TV5P75FcF34Ofu0EoPVe9iZLi3lQc11Db+uD3
pW/YaF7dP6UYmUh/HzYn+DeR4NW4xaCcawbPMXkV9Km4YKJaVLtwMDoLgL/LwtnuKrHtMo5lVMqb
NfQtq+xQdFwA2Rm14SHHepLcRWeyIEGOu92V3aPUTzH91l33whlGF3UCxOqFhosSkMr/3UYOroJI
NK6zjk8A9SVAu4Is3WGkgpkPbU9f7frR33nMdkdvaLMQSOvWtRLYLIa3bJj42l9zpfy6nvPJgWNa
1VP5tCE0GoxBti9We9ThgJEmaBnf+0mJKluZtROSqJjmwlj6TTy0HV2TA1JdV45cLZVsM50wVD1d
2QjmvAf4uArJvDJu5SZODOTLoiDjX6ZoYNAj7SRjlaJPV2emUirDME/n3hnyN17RkBvihpKBTB5c
z2CzXE0gABy+4fXILSPvOuoZ494KISctNPWAAtibyTIDAWnwfkVhTpZ5FJvTScm4OedBAITPQYEO
COwAEr7WaLmugrd7WxxfbyEhLRTvG/Y03g3PIqwMzVMu/OtNDamnjAzp2QPMwUiNCYtMF1y6vrUN
vOiuOsEcOV8UsY7QhEtCW0ARGz2XmaBpSkS2MyWAYerg0Lf4gCi4NfnhPOeoc8AR71pYDyO5Yp7m
22YVcmB013/ZuwkndyFFxe9d8rHMCCWo+BasC8YlLd8WCEIlg3oRmhC8mRmdnGZC3HTB6PHqNs78
ujHABZsn3XuMKHDvmCOy8/IzaSqBvXbtgS9ZfzXeGdmhTO9ekNdZFcER40UvJKqkzMpBsSqY0fkN
HhsoIb7q66m47hp6dww3o20RC8jRLIpkFAmsHYe8A6rrJo5gwSe7Zmwxcrfku8OZ7VZYrRQgqffw
TXFjIRQCYseiTdofZOpzxj8rDRCX7kFCu1rd98o8cPrFFiSTtpYqFxaxkzaqsPWxb81RwrhXwJMG
RHE45OwVnFWkbUZ4sAsOfXFcEKc+SRrS+sJ2XZpsCdiegZgg/UCV3id770xEn966RJRUkJNuqj+L
xxH1L7KdByApF1ocbD/jXYDrRlCbUu7WEvu6KGPGhjGSRmPtzfcoNTLS1KwR66j1vgJvOZAywkts
u704EgfwJO0THUUPFKGtB2Pmn3RPeixP2daNYgWpGevF7MHZH6E1gyQynWS+DIHYCYrki/Mxvw7h
RGjDJQlJk9bk8yaNPZcRV4HS4ErGginN8q0K3waAUcsaAGFTrqQ0QFtxz7/GRboOyCm6dE3u6Xlp
I6nJjc81vANGnXDLF+3qfmir1L0pOxm5SNYjhT/qKU+Zq/tEshK6dC12eI5KHFaULJg+8lSvB8zz
UDV3OLfq66/4A36TkNg5GShNcO1TVVELCd6b8l9S+qjgqaMbKv7eTtWQ/LnfzXgxHFZnF3yTpOdw
VYk/b0Sn7iMf01WacNXCUdZvQsghlseab6l5sPkHF2fqp9ZWcsNpVjGiTaQnUNbiNPco7hku5oSf
HNQRor+X4soLVih4a6qcPJxNUQlz9wKhqzFKgKcDFX10wdcq0NZftg3L7lWAE9DldlZ+OwUi2JKS
O29n/Rx46EyrUOBvzP/68vTI+DsscbtGjI2lw4ulGIJ5KKlZzHE0fa4HFdBbUYyhWlH+l2/PVX4p
yuKqtVjIV7Lj+9kNwjrZj2mNkVLzp0F8RSw7LCu+7a/X8v27lDx6tSbDMrp57qqhTmmcrJP1cCnC
n/3PbYfiOyXFXPY8ntD7wtasVHY7VfeKq7DH60H9gHS0Gfqv0EFWvMB1gJ/CuedbtvEBbAQGaUn4
w8soLErit9w+xMCjO5b8DMKsis9NOp5uFrBSzT8IqGJpLiYuSVQ9R4CH9N/RCvz4fFfAiFvEhpfJ
Taz42WedzJMDPIf9mP2giyceDGCRfCVNb7dT3WvWqb2sqFHb8QJ5oT5YNEguGS9tTkwbZUDRTWQl
ZWNjuacvkxQfUoVIFgiW7j7cFWPWLIJykMN6dmDyocSjYT6jT4f9sTzGyEadKisi0YCgp8lUL1SN
+n0Sw0u/D134YGpEHyEm6NY7eKpJ393PsDSk1JZ8Q2yrcHCZV0jHn1MB7R8YIMvi8rEJQ/YS5Kpu
PhwSyaqJGxtisZ/6C33VMBJvMwGkxRlQ3G8eWVw0n8DotMKXutVAS/BJepPRrQFknHf6gaeMbZw+
Bxz9uQ5hEXVcaGyJ+tE4cEUzj/aTqqsrVWY0auT9Oby6b7rS1g0dHqiNbUZD9oV0LPfXYMrnxbKc
nVShZ2x50iC/sxqgtZB9hyoGgkUFKGs7hN+G4KTGswV7/boHDgR6143OjX+wbz2phJEqnnQ5FuxF
xXab79DOJ4gBI5yamDISvRrGd252P0DfFdTqxYtkIiAg7QOftpLosDhpuioBImigAVL9d7/3tpbd
AmK+TYxOFAs3gPLf7s+K+8afgrHSKZdAbfehuxPIUFa5f1YVT8/5KPCE4y4iJsMdS2a3fzcmTsmV
AXiKQVEK+O/7OoU8iWXVv1kqft1EF+yXf0wbyw11EFuhwIO13yrMtvc+oCAQ0i0eLIFuZkz2424b
ppLVjG2trAeYKyfBYOCor1gjI08Jdg6mkw1EGCCcR21CfwZlYlhpJGvV2nUR3OWwfkEABIVlElGB
l5rX95Y9JWDI2CP2hAhOn9bNSijC0K+gSnDorrSLpuNvTzvSuV/1vnRmyRxLELkvy0i1kOA+aDrU
XwIYQm+3R0yQSxYnXEebiXsOriGXD8ojOfGe81q0/8aXQlIYnqKHu07J71mCCGckg8609HHUQFyM
VVLT1vRm0FBUFgMJUWaw2y+7ZEavHCZGmLXPAzwSUOGU1h2ww/jxQCJvThdmqgw28++GlbA1Psd3
auu/z1SXYoVN4N7IlXgLpa6SdPVbeRb0v2E7LDq1oLIzxcwSmHUFb16SPNVwQ5m5OKeLmnISCRC7
a89ItZ1XVqKsW3FDtIbLfhDDYY+sw0HCC0SgbcdMIzbpRe35sKn89PiNdSbbi3AnXijBTp6j3DwO
I2W29JTStn6xOF1lTDsdQ7MPEKcTkOIiltKxN8ptf6sfXrQOhV9dyRoSyo87GyZLsg8fHuo+IQgm
sZcsd9vuVYnW3h6ZXtgOytFryIranyBBxIMvIIhY9kdswPeeSlz56ZM5c3eNbrJ50R+Xrfx3B9dc
Z8GQ/ZW5/Ipd1rRz5N5lCXFcA9g0eG4hX6OFy3aI2CyTIRMZAc+gB55839Jpj5npy4/Yu5w6HFsl
4ckstj/LHAad8GgVEIEKQKX3Avn//piYsYLDcAfQFdN34BUs33J8kM/wMq0KUCXGZ4ZxoGYbwXF+
Q8BOPC2HjaBhFG7MRdpKMtrl0raW1AfSLKVam0ki+VQizFkM/hRe4btSOdgF8dVp8NRzo9QzHaDj
4mnzIUCeZn2wowCDIkOzkPfPM5cSnmtiNsbbzS5IBFDpA7h7MPd9hyQBFuyaQdGvS1o7x3smvntp
tKY7nJ7rLhBRqC9DbFPDjdFSs0EUQsLzEMPRTQ8IhDhiJJ+CWdBKtsv6TkMLQY9C2P3bBhXzC7Vp
1+fEQv1hzAcye72AsCQ8DU08DcZluM0kACuYdL2PP8dlyJdNuXRu8LTv9vbUoOYwFhYG7sXFCQWc
Hjek/x/aLlUVnXQTFMW7Cfq0AR6k22DbLzejn9qnwhBO1oihMaRdB6aSekWGvffpGwnF7tGqXglP
wdDxOhg/ijlupKJXi9p2gAPZvSsQkZKUD7dXnH+ww662U7vkINi3dWaZd+tkaIJ5ElYg0tFcNQ6e
mdSu8mK4GH5ZlaMNv8I5yZlpEjZMDW2jzaKKgNszytFfQH0wJJyrR430Mcuzf6KVU0sPJCH4SEIs
QWs6egmOZMI+BweYNH12jocncSQSJtOXhTjnMMaQdL7SSr+XSDja42U3pS0qIf7JXmi2frvM/MxR
Th64I7e78kbUvEtHwvAWqOeCoUdj0ChMpZtg3ehOAUnWhn7R8GiSrD2spTJlHiMocmxahLFP/NCh
QN9PNNH6m986F54LBbXRjWAuCsqRZh8jSLZrbIEJ8UPqfJ1RaDhS+7Nk1s7qtU2OzOhCh+BTHv9v
xABXsNuB2HpOcAfEMXp1M6vjhP444M+oFGUNLAr+YjKdBB0HxBJ9a/Vpjw9FI56mIqcC/7aAfxoY
ytnHwTcDhbKD8AIMgCpbJjqm6Lb64Q9SpdrLmitTC7XLTHj7kNW5s5cOhfqqhthvhCvu9TFnde67
CtgSMmVM03oJqqiTqnn18oUtnmhuem61lMLKXFl5C/QhcitePQov2CamC3uZnEUuveVY7p3mUSwd
rbClAUSGXm7+sCrNQ9VUfKYCrGhnUgckaRiZxTxzs7h5mT0Z4iA1TO88ZAeEjfyB347VoUcwIX0R
MAw3TJchn7tXBFiAFUyTeY6gBrCcWQNaXU+jqZd4FdHccPk8bL2NWz+Mq9jKLnLdKiMzYSCtFQud
kXBAFUeXwdGDN0tktQxbcksEMsHlKkbQneHBHJ6y8v4YWVqaQN2WnpmzAa4Gifk3UmNTxTF+qEBl
3CdY1oum28CLnPzmc869Ftzn6MmX2Jwl8tX1DXzXrkGA+Tpgtx8by4rbJIgKZc2RKWrTV9j4Irij
9PtZsNeIrJnzZ3NcpvEiCNFvOi2vvYXHjdzp10O6JnAnKt/hOEzS9oqUrkQjWixKHh6vSBIR/YdP
CLBATT6fZ3KN4/0qpFcBb9Nps/Zs5hpU/hD837pMMXL8kglkmWS7wK5gTKWVnI1WHmsbhgf+vp9w
ASlFZ9qpz3Wh0vV0ivjySBwEjFSpcYDlL7fM5LjuRdcuqJDumP03CJNnwhzTmbeIkqfWdyzgP24l
UlToPa3f/r5E0JsxmUej607Cz+4Op9Y1yoQJg5weUcMNjLgFI2M5aLXfvOjOu8Ahz2sp1iRbio1K
jd8f2AzbUk4IDjWYxy8nJ3h/iJc78K6Zv8IAh3zQOlWmI4o/5NMgr5tPTGgdSrz+wnfmvP7+7JrK
QVMb8aiSSQkTuDWIcGhJpgt8DFZoRk2VtRYv/OT9qROXqzffGCPabmpAVghK5QkSS2OlOY8joJRu
a94dJA0QpaP/S7n3z7oRugBdUWo2ssr7o3vCecYmqYSo+Fs9f2ldrlsE/73PWKXfggeH49LLCbVr
30pYfHEUndGEwQcMJTCWhnYjDuad+3GUjNymQioK4eL9QgiXHxtge+8L8DXko1v3Pw6dmt5YDqTM
R7nCIj86r0dhde8QddSHImV2WDTAWC/XKZsujTJzrl/4RzIh2Vy2pGWLkPRM8AlGfT9wu7I/1CdE
NgiCKr292hY70HhuYbkxv7FgL9zln7NaP51yXxnNJDaN/GFJP7KS+XEbbQNN5YcEd0KVJI9Y1Wos
ncHLDx2m6ci6++AukfdPqI4/91mhWcXZj8XEzfqtacfZ84GcN6AtefmoM40zwu8wGurmm2otbK/P
JcV7GnV0A42VQNEVcch/LkQvN2lYRowe8GX0hEhgYBUs01kuVm6s8tG2qqg6CphvLi1+qGuoQayy
tT9Wy+JKk+VBiHRlHRJlw3jE4RlzP5kY1tLgQw8D+FEo1OuWTOYfHoNSyMjlFvjdrwPAEvN5A0xS
8Q17VYZN1zUDNUU+9iDd/M3CFRDgwj6EXj+c0nNHUXOAIGQ1/EFjmE0nTNa39BtzT7+DKD0fxQiS
K48hGfRCCAgK+wrpiqwOMCrLtu3YbVy73vx3EwjFTcQ4nalzCW3QIJQv7XWN0jKEBFJ0iIXYkW+t
ZfupQTR3llq1rwUHgQmgRzV55ZXDyUECIo8ElG/3H4MA2cuqZDAafsRK6QcIFpeyVQHKdGyCyv/R
Ktthjz7vGIjOeg2rFnYK/Ra0QBEYzCLmyZOixhtwphYGQs7MguytCBF0gGk7FI3/ej5ewJv+2Xxn
rBCkFTRhtgbAiJ90c7BG7cUo9mkN/wgZFNVQLfbIjnJ88CuT0exV3dxsEKLfJDvfkWBLhwXF7vuj
Usw/arlvwae7K93Zf4cPbZfCaOgYhitiCnJXk6XsgNjUkJUuGQrzC6tSpr3XBEw9GW2GyjfgUGFM
XDlRP3IpJQcZ49ZIYhVY0IOiVR9G6chgH4VMnjXAugdOpfwBYXWZ96V6TFUA2uY1o4G31Bdv/PFU
NT/IFRAx1pVUhX2JJdFk4b5qDiWldGbJ7RJHWBkP4EvlSqKvKnYgL37Ho1ysCZ5206H8/VQqev2I
T4wq/OkcEWY22fpfEJ7dnzInzcz87ILmb2nXYeb5MWCd0HnHMNzNxXuUqbhCsxbmfV3uYBru7eHx
hqi6ZlP3LRzTkVVSYxj9qxDviXr7hohDtwcuGzf+n92dwrhaLJmLUnJDvXR5QVjWhm/hg5/KlywN
3IVD9q6FPJJ7cGfPQ9YdYPJIl08DAk6WhlSE5sDIoWigJuAXyhUKyadx+IHjGxmi6le6N/mTXDIT
iewhPRksB/QeHhPtyeqK8NI0jg3rQ4lLHSotE5Lt6/jNKwdIjg4gvfHHWvscXrJTfqCAGlTUEIqk
MLgrX2IgQ1i4CK7Yr9SjLtvrnPowXl5PSEnzwiyXVHY2laAehloPMlmHWH+YC4df2yTrcXEnT+35
HBuPu5op0+kQAyXoN7WXEFNS69tVCzD5o4pS0Zn4w54iZXLlPwgLEPAUE2pXsDUGeLSF7VCqgHKI
uVE5RWxl/ndXIsXaKblFNhdrfwmeMkkAY7Jsx60a7UC5H9jpQGL4Znq66Pkd/hYIvF8FM7nuyQ7P
4+8ZlIe20/NtTJP4+slWyI2yjof4WgdD2etQs0OauNqL3GAwJjBlvMfzSo2ncPHPDF6vMoXZMF/1
Wz2kZasiU65NjE/W3A194qVCGfSw+wQ66rmR2NH/kF53YbfelYjKtit0973rbzcsiBlxgRShVyCE
X5SWl1etdrW7r5KZaCb5Z7/lfMZcRMy7sdOoBkqyXhMxvfBPTjd6hCEI+O3fMnhzpPY6gKi/Dd5n
MTBlh+HmAKP9qoSyLIJgRuSjf48Fv+STCSGDBUvNb8MrqanytmKSMLR7YW4bfl4RIqesM9f8iOkD
iFXZHG2aGTHf5pTktngxukjHc3zlYlCCqp+0qT+UfLkPYH730E+1apds5UFTnu43r6P8lPyFl8c7
RzomLbLMKmG+sM9COuwLVgoOIBRMlJItDISsuk1G+x3Lq6ehjDoawVkZ6lXxYYnLJWc1guwBCSHg
Dtwih03+i4Y49Og3sVN3hlr7m/H/YYo7sKU1yHf3EWSb+e/Vc/Vxk7Ujly4esrWJFFuWzIhz1qmv
nDg68rAO338VmWZKnK4sAx/RcRTWngHoOXoLDE3HXlUi1w2TpFmHpLediwA3YJFPhNVCERSf+iox
NmKEX/1MFejBjpANPgt/9BlZ9nA2bD4RmcWMLcZh97HBauGJkKT74tDVSB1qj5lFpSoly9qGFrcN
Q5cVDjr6HBQQOEPf8Y9zi5tjrvXUJK01mmotjFsJGKk+c8hJwbecwpeQHs4zcJBju4oVQ6ee7Ijx
4rJnOw2tEsbk7TsEb91C1QOI6Uv8F3OBTnQ2wk90YRlB8Pagtyw4CzT1Iv5uOWoV9J4UHTpDvLtf
AZTUPvhxmxDwPPT2PT9Xh5MUqOWeWsPNCEKwDHKZR5yGIF/FYgGv/Z97AzqJa57/Q5ce+ZBdqjNe
7WhAubtgHGBI9kxaIz9Zc6luz2P/Alp7ssKHxO68ZFRrgpuhCDfrU/4E9V/K9iwEDa7T5fn7JGVI
xiUxmAE39x30Cl+LmqtyAjwpup+PC0UEHgVSXZb1VOSUE00fK2Dhz6iDfoLFqtpaRZxFl0sEYAs1
QTd3Ml4cs45itnS6N9CWDaX9YoQLpHqarVZ1Fsukeirc6xvoNzD0t01jQ/zbv9rMCCnauwwv5eK3
JPlg6clxcziOB86qHBWi1fqTQKcvC51WSmotB79sNPLwUn1VR8nOsE28QfRtzrOkwXJ/erXaEwhL
rsDMVxn5JA0VoITleBtmGpKnb5YdOuahSkSBoxREbbPlZa6fmpug3DQgGosHZJ8QujyW6NoUL14I
V1piLVcTUr4ACy+43QW8pqi8NdF1pRjlNjqiGbUkAkKWxp9dBPcZPCG4XlP/UiVHMzEOZysOhfmk
Ty6E/bux9+1mf04LjTI0Lmaw1QLrGC3VaHMRCDXU4aIAglWdEKU/LvuZaHYXHCXyQ446l4UovyAM
EH7YbkrI6RDjPULnvd0/vFZeASe1IKgFxuNi4uGlxh+hQhYaB/lRdoGDCU2CIUA3hXWgWXCFfeCH
ze0iRTPNEDa0fgrE4GqRuNCcfekG//8JHxXw1t/MoOVgFdzlPiHmUPolEzTwIu0BPEdd2yoVeCas
dcquS70iYXRXgPtSWMPRI1dAgA7/F7MQiR+fKAoOlOTMs7WmjWbvO4mKTBODbwcKUJDWJM0vcDe6
vdEvmvU0JbGGmCPCnF1Guhme+kaNJU1FoALUejLZt6hxQ/oyaphgqmOogA/qii5V4+zQOXtTTplF
3VM60Jn/iWJH4Wn2V4mE0m7WukWZH1IR2YPDOGwV/cTvrirJIaSpoUlaC0YIMdUAu9qeOGdJ4N14
7rqj1cn7FKFF/DvRoYnYlZXyKJA31LAbuEeAipskw+0yKRNmmc2TYbe956iTEvbkGXpLYr/HzOJM
4wU60l0ifUFoWN+/UgJk291l7XFMpIn5qtDDOhdPu31rtlBQLXju6OxDfkXMrxSTPWrxRdyqfMWE
zCCGfFQBNv51CoDx4bq/mRXbcAg1+nsHuWIFlJkXoXy0QMYnxnLNbSNwkKhRMmaoYvSECVhgZbp+
jDRrfaUqxwwUdg0oDgf8RGqlq/8BwTFbQFaSZRV1/LFbUfhRWyCfEnqnvsjnJOyY8l17BKa9kcpO
TTaHszETXwLuZssGxk2seTmjOn8FjlPAlF5EobKOPT6dc2wSazX3DoHCHN3xDtDM17pCejNEMcS8
sWDDTFitTu+r7JqQ8WtdpD+B2q+rHZLAc2qgz3j7RdnqBvgwWBJwKrfHRgJhADtSFhwThdj4EOw+
D/81zqvwWkURXGILwrh6EOPNXJy1Yzg8HtrYLoCZWtl1vwPJnCnQg/gE0GyL9NQ5q4tIRpGTMovI
IFKXyShKCmgfr6R2kvLf2hQj8Cb3OkxgT2i3jEITqU1cpI32gcIKOP2GnbYcxQeBLUVSq6elEOsf
XxWXM+pIzSh8/OHS/AdBh813RlzbB55PYRpj1s0eCA+NKyblOL6lLhoishTMHnc5VlEdh2hzyiDo
VuEi+kaLHvfryfpeTkk5ue7Ycr9Fyz7DDIsTUaXmAuv0zQTED672U5V0IuuJaFAM54ujnl3xFKn7
S7voTg2kHB0n9a2gWdpvqQqcEzNXcmkoJYJVKo1fRK3Igti+gVQonZhGQvIdX6IKaOWB8hQJEbrn
nIw0SFvDNlmHUdNJGxb5VJ/hrDcQsuZYD24h3MFh3tt+Kwoop/oQC9HJHTDS/po2geP2qjFrGLWS
nciGd/bWJTYNoptwYuGfzDb6XosBGCVqfR/2wOVqo/OmsBiKTH050Xdr00vg/8D/e+mvouVOOShz
vLEPTw84kgprgb7tFT+tnmN6WkZehQ6Qo9gaeVe08UiE5pMlCAIj2tiXzwJBHg101NbnhW7xirlm
eqmrUETT6/SPL+Suh2rix5txJhXbX45lWz8kzet5oViuDRCE66YG/oMQq/dxZtasDnakWxNuWVEQ
oiHxsI1Rj2XL7d0Y4YT2KImbl+MD/HYNXzXoImGUga1qG9r+BNl7bTTqQRhv3KObyAUSNbZ/jCFg
jF+mrRbebXUHCgobBPNHfaYoDUr7cy4XuC4KBUZsO7HpAOett6OsF+4lb7CAxGSCwHsJfPhi5DMe
ht77gpaa0wsWniLUscvMd0h6+zU/8mjuePpML1AvYKE5ZFZLlQocUaI+EF0WF64UuwTMnC2U6SG5
j8+ClVt2E+/O4Ct1lPYHbSvtc6dBEFa+iwjwCS8FFaNcgHFhC23CnUv10kMnc7XexXS8yVnBKbUY
0MsPS9oov8bzZZU0zBDNjmnvL4CiV1weN5v7J/QI9+eS056fXBTGjWqqT8XL3xvXSfkxQXQHRAGh
KBjw+T2U+LWBkt9nriqP6dxTIVJtcsL+UBdoFhE1hKUA6fDvd0HWlmZjWIBhzk+5HTex7D7jikO9
m0BxrwN8NinyXjDhziMf/n1WWzNmvp7DKzzp5YiT1wBMbdTEUWFhM4dplUJyxiVZXxBVEFSDgMvU
j9POBKKwDS/iPWREeuIWRVQKDXMWarWCfi3UrYMhVUG4briH4TN1RF7kv4s4OFbTVIJHmYQ2mVmS
xUpYTM85uSR8CowMv80o4msnGlO3RR8fNbbm4LjLfLGaRxJvovy9xn+wfXugKk6VlTAOp9LLpiwO
+jDBX+IPNJNdkWedxfADNHuS8JsnIbyBdd4EuH6XBe7F0zYOBykPfzUSq+nCC3zOqorpWmpc2MmF
FtcgJbMNTrAsWQMuOjT6VDKgo9UgB+JRorTDpUwUNcy5XPLJVONfWoX3WeStffcoQg2rv8NPOYll
CtPpIHaG25t08u8K1v2+6tMjEQUiDULFeIQ2YtQ5QeZMoLufwOW2+kQ38GVecfG3QxbmbznkYwz2
skldxmjffGLLvVrQ0GVzOcMAI7vpupVyXWdVp5fxA714+rOSOqnJgfcjkJfRft49xbjMS8E4253I
wVfgd/wPlqjzqCDuLISDc8+vsdVNrpDN/MpciKfSAeDS/J/L+GS9I5jU/olE1rSyWSRea/yd6mHb
dq1rsfWqMNd2efprq5en0K4i+fbg9irrURFZPdHtiiikoIuXadzJtTB/EOpko0c9f8hUu3pCch9t
NWbo004E11jRft2pikx/FYamnA/mZlj0ZnS1j3WWeNqIg/mEdYwGlNSyc8POQGuVJPBeO51XrFHI
B1TcdpZjRBIv6NAlE47WMWFRsLf7aO0GOUMQXnBXeCKOfmzm5ffmZ0B7D1bQPwRDAVluv55hOIX2
A6rZMNzq8JnfdNgee5aSQSvJKlAvOlc0uHAQ04CZFfcM7RCj9q4p2nyL+5mgWtljikjD9DsS/pCN
3+OZRKf+53PLYoIytmCFoW0vB0jDveY7u8FJNTBwJtpgIwfdGN3hKQ7NkmTDKCHNwhjBsipzo7g2
VAmi8mdVnIAWEwzPB20dN3YPm80/tMjoAzcRivJXm+qsmEsPRQNVRti8DkdkRU7a/3eASIVcTA4R
ZCIFV6rvaDWKrTGRJl4i6ktfBDi/i5XzZ6cgFqJ1lqiPWoDKfUIhnm6iJHgUcf5F4P+U5bQ/971J
w5Lx7yo6fJioHYOupglZpfAG3bnk5l8fN6sMpQ9udNoJOoPq5GVPIBJdzOJGEe7+Q2puDYv1Lbj1
8WeYdbcVdUr3aSXCTxhjIIMOHLnRjRVDS0kwV1WBGdagjOvA6NQCs9svnQp9kAy1MNU5TqixvfIB
pw0PBLPtKqscBMt2FurosyIRN20L0DN3/ysNlLxFQhzzDz74qlZHZP6OT2KcNMdeUgdMDzCK2ZwB
ldGt/E8wFdwYuImEToVgn5LDvP5cs3S9fvuDDjSiibOYSgu1vicu5jX4ltBQBe8opxoj0/jVCPNJ
/hbPTWE1r5tiP2l2hapDYDewTjWAOfDBMFsotUki24aV6jBCseUNl18uYZ6or1OtYnF6geK0ewOn
snUyAV7xoDMCqbg2T2X6Mt9UbO5RchZnBbgwjGtq5NsowMvZCEn2curM5TaW5isnnZAhsj95qHKU
/5ZEYkJjohEFhd48sHfO5kiT9yr6b6VRN+CWE13Tay0xaCsXpKef0qNI5oDqRsTBkLwt5opFwOuA
05/t5ikPTfFx8uec4xOdBFeJPYkQW6+UtnLPNwKdK6DiP54vEL+3c0ZdbtPzmyvIIIwAtatu1XUe
THggtrB5g/mxmbiHxh0qWR6l5aGuwcDb+ZCii2/xKM8BjlMJIu2PXmLeYIJAQoK9tnkvjlV1ZSVg
sEncao+UqxR4xIhLKoio8SK8VXkbeGAkjxLwD74ADsu6jwSfxcS9qtXMmnFj1Oh31024a7iNiC65
IMPzAmGIQ7/KTKOYXG9zrBjDrDk1irES2g7b3BUXFUXxoaKhxUgxn+j0m04AyRgtThyJErZHxCih
zvOOWujpqgPhwtDScGFsozMaEJPIKjhKE31TLq0L1DZIZxMENszghTdS/yesacplp9Smuy+TzzrT
ckWHmsnvjyi6HqmnTD+0l8LpiAasCNp0Cq3UG4NYlzME5dYEHe5Y0rVvoYy9MFp3emJ6F9RVZyGQ
3zxrngkcIFc5fSAkNaEtqMyBm585ZRK4DIKXDjtbBp83oai0OlCaqGmkn0F13qGICFM9adUenJXi
g0nprPXKTrIWCRRUlp6R/KqNZ3ngrwJP+KfLuGUtFX6uqpL+rsVBJ3yRRsJZFHE1Vi/YuF+Edwmd
R5WWlB2VfpVHgAUOOEX2dMeR4WbJky5UeuY2ZoiO4xypFNxk8g968iixY5s/mZbo0umFRtx8eEfd
VmI719QS+5cGtgemXW39kCTL28HplF/avVIMQ2WEDs84o3Ad72949A+CQdvCrSXq92Ekj+DaL+GU
V2uN7roIk0pjyRLNxBctg9hR2ikV63wBl4D0gPBz6pcy5zt28cURW9exzkCKw6zHvaIcsTrLei7X
tPeMBjHzd1pG0X7ErOZkM8TJhNk9w8wEhH1uGkvgnR7GrqDDwzZ0vLNcSPWnQQVP7EbnfxqJQaDK
ocY1XNEz6joCDmwwKFtxqzxsbMV3Hks6sqBx6njUuRukP0XX/LSHpUGUzJpEJ5lkAoxiach/XXwb
F0KRBjaefXugm7/VgtozfGaUWInIRHKdkuHqawf4mfxKJtKD8vKLpQgM4CPOdyii5uhOTyj59llG
3Gd+ri/p31Xzy0Fh65zYvy7aHJjr02fBVSF8jiEJlOTZ8CDxcKoE7HKrK0svVSTRVhlILkWc4X87
B1lAMCQ+RkUlhc6ZAQEUXD7jHsMuFBy3kFImdn6/RMpFiMdbYlPG7grwhpq5rqOtMjMONMEpLG0d
QAOnQxmGd6JrzzxNEtyU0/AmSMUBlJruFXAnk7cCQ1+5JyUxwWoCqdl28QBusYpl31gWygLo+Ev3
CGJPX5w8RbVcNtKUs6mpzORbwE4RXBhJFU8iEx0G5zahy2hrwJsfI2eK7dnsJpllKRhguth9uNAK
kcEq07Ff0ioyFjiPe2yfeqz0ruXa4gl8J9NciHN7WBx15GHQa/ByYtJHWm6PUY2ghndxPFUVrAnL
tb4Db4cCCRNZvEC746tuXMFl1xOFZZTsCAsBG9BjbXPgeevwHUNIe4QiTw5j8oUBERSOWdLdxHvM
yQSdtWHFPMBWNeCGHOMKphldW+ixeTSY4thZemY6JcSynuPOjFzJh02wTlh+jRoM5t/yzIz4sv80
vI/elyf97cZ5+zyLnQbC8yIImQZlhnd2X971R/bKPwIa1l+V83C8NxS1jzKeyBBCDCrqPjzG+ZYG
qqjpgpr/eoYqryIUy8KOU4iSclFkNbDx083HMpuYCUxLjM9Zf70fQihO36qE0KErK77KEMmxDc3W
idFQH9MNYFvSSpI64W9H8d3oauScvO7Pq7VEwEwWGBVIHJmJDe8rEwTTJDt4DFJ4E1AZ/bLmKXk+
7GZlWtET5v13aOFfR07UTYotXSFYo+ECXYaDyne41HtInLA35mJiGaRbmEOtH7O8VV9m3APPn3MS
apENpS00hrQXYRf1lZiJUT+0fzASJA41IMo8i04dC/oAsPmLsrooLHMeGFkDiCPMAYL2N90NPENH
uJYcnbVL7ReIhXbIWul+jKTpPyiXRmNFI5C+J9cfCLpFjtvRWe7bV+0AOrIzxZiAUaEZoelC2FoI
blKYUFXJofaiZWszDtIj2nKOfN2H0PNEL36Ri7IfSr1uFfS5ME2D5hFY13PK5KSWCZlrYjKYK1dw
4RbD2WAMvFb7faV/Z2lEkZLrbhuqs2RaJ1wNl4tAAu9B2UCveeWyrNJVrzSfFGzk7TCa+tOcNC/i
yqLxe82zZfEGvlqNAsBacFAUNzuwPtyY2f6qHdyPe0znZq7p8oHIa69E8z+vUbaiVZWZDBZqp+Os
ePNZ2RcYstlKj6yV/iT1rdsLut3mzaal+lADBdcZJOkirStlXlQX9old4XJ7hgLVQLSyvuvEfPly
vF7kVoIv+uSiBp2mXQGakeekzER/ScMXSxgifyO7BVYPQ3QSJ5IUWD4LgHEA8RaB7IibwAM++2Xx
n+NoKMNb3Y02xochcyKF13CM39EQSjr92m2jAPNH9qCtEAazzpRkICsgFBw2JrkWjM/tyGIYUsT3
Z2LvKuoE1tUyvzRlZhb2Coh2h+4hN963sPZhqiApRQsmJM4YrhG6AC9WIE3is8qq6/7k/+PsHb4Y
1ZGALdXZwyFXonP7KhEStMRkercR/IkNGCatoxgU5pwwLGAxAQ3nDAGQ7iQuZBHOqTSCjxnzFDGF
IP8AE3Ke4eAqp1ztNRvsWyIsF/NoBmAgfn2C0fHVhdk6SHdV16J7nMpBCQlITsbCWazB4vtISn09
Pl+JjV2MJxXnEOnlxrwmEz9xdHyJ+LJuix1uu0/MWiwaC2Qpy/J5gNax2KK/GJaQI7KYyfhOiLFm
/pEClG3q3tPmq99sCreuYoF7mh9II7iPGFFsu00gGv5qNuCtRkax0OVNqSlvpOqEpG+qC0G7JdrN
VcTWMiWazSeEXUNcUeMuxqNp/jp+xKrV6ZzL7U1j1nPvH35Skn1yx1QYQWPv/vS0qnm6vQMkVS57
QL1gwICPYPcrgd0BQXmxIYAJrOz7t9uWHzTt6vT6SHd/rba2ktYclEuPW+CWKIXPLBbWzWtR5rhm
QIPrrkMAgk5YuxCb9ZPgqabOp66K8/KoiHGcgxcIamkE2EJyQFzm9z/HYZXHCPl/1q0eGlUNcB5x
vUgHf5jSi42TvgRDnOvowB5FahkHOlvAFktq3+yALbx+5+NcNysv/iYDAEKlZy8F2S+wDeI+9irp
N8sojZbv68wMHGgrgjwx613g7W5tuGTzx7Gox3/va5JRZXC2DNvajIeIU1cwG568iL0IcgHSVa6X
m3T2PZVfvgFcOZziiRSXmI/cuKcw7gacRwDUuHJI4GmBNbO3EskwMwcrHoUDbW4JMXoqUvqbXfl/
PTYZw+lUUm0rKzxSl/Dy3agYLFevsKB8CTEEq/482UZpi5uiLoV2TtGBQNt228iiuNAuOWgiX5yA
Nuq0t9yQKFxwzpASgDmfmG9x/UrfG0LOCjsa7db5oQ0a5LSj77w1CaghzAfwy7WZyBa5w/omLliC
9KcEbRRYVgbVN6GtCZp0ub6h5vMX/iLtubGtTi0vKx8q/6kbQPsqbviww9p9fjOSFgdXDp1W4wFc
fEEBflqyOGivz9DrsDFxgk1uXRRiGDfPBnvc06AhVppr2bvJ4iUCPvpW9v6Sso3JyMbL260Q27im
xR9OCkVow4UPNspg+pvyrItzE5KCk5Mz/s/xtAHl12D0nrRvI4XN/4FA/wLE7DUySWBQ/8hUCE7F
lgIbWv0KfpJPYA4Sy0m9sP/h6fKa+t7Fag8SAbnHuBLVSTxDayKSkkmTeZCXkaPR6Dn1XbIb8GZO
LcqFk1HHKy2g1SWHMAUe4vRYHbWm8gRW3/yJ9r7hlpBDT4QMpZYqxBlY7OIbyqxcAfnl+swZhSBC
svlbsN6QY66JDpPLl0/y6wkWIEI2ziB8c9Q1rq9fmi+skgugfBUE+MAgct/tD/Tzf9AaHhvB6u8b
yJrhvlovGW+iNpnIGKpvcIYAurpg/dY1DTZ8rFzm7xhuoggW1IYCdpJMHqS29zEvS3hMg9oQQZOI
PTeXVCxmOksxKwTEcLLC3yy8uoY66coa0zDJjAkCAcxsUwWZpS4dCu9KKlJpgmAQ2BJ7OigSP3F3
FsHqGX376LAmySH+YNcg+G4Or8Muth5qLb+8tBrcMhlY+gqk69O3qguYQdKdu7eQw7ngxVfgCl/M
6NTL2lFtbfKSbjzh06m0P6oqmQM+0d6tk8bYgh6lk57pf6Snh9mQcFBy6is7EdRSG+4RiCKotybn
UZ1auD7bq5nJju8o4vYS/pVw2tFI4J6S03s71eEQPn6cZeQY/ocAZrFxFYZhhaWZEftyw24O8Ydn
FA1ZEbxaMeMi3Mj4xZicgLOLdYzeWuGsCGFVKRm1IJyzfsjKzBHO2bSD4qyx0s/SgYRJLO8L7VDq
J0gdIUrj1pl5ZxNK4pZeWgQju0QjBkAKaVOjYPTDIf0ojqG6xiyQzKhwH4jXiKzbusrelM1GZGnL
Erc2aMeGoDvqxoYI9GTecOs9uR0g64pHJjoRabG+o39aUm8pZu5CWCRBCXuoqlYVXnC3dVMeS0Vi
+aXpC4Btrhy8fW2OWPOXItFqcZWoxZe7dCjLBhWTX6ZKermaeM2xx4apOTuu7DJpLEnF/VKO09vS
yE76SYdlTw+oZtlhExJy4fYLxgs1aiA60Z4sURfzS6pFdpcCs98V8FroROEivyqSZAdz4ZRlWvum
AIuDG+AHfxks2UrMbVzWJwxiYU3dRoXrnaiVPHmxKPF3HmpnL8sMilzDT2mDzkjalnonvL3BYmr5
XrmBorZpB2kBEk+47Ee/DM/GNgMLTJgrTx3Z31VjqDF1uzLYqRP+HSQy8t268GB+4T8ZGplaG7GP
sQRcwHFlfjzxj0NCIVuwldrtH8z5xbyAPwqYTg8x25LDAOj3n6QS9Ikf0UtTC5hF2l10Hh/ghKjp
c6946QLy11n/48fbp+YcD1W1ttGWrYU14vKUgymhYBvTm2OZohlWhsdwfhy0bzzpAdSK3Sh5rOyM
FEZUL9JBoe14PUkneF1jQZPzhtvehtb02z8Kbra3L3GXwTkQ+ShVaJP2ZoUagaTlv3h1XbTCJCKi
wnFYVruPpDV2Ou+s5QYJ/3bWIQufdpwB6J6eaYEPCuDRazWuKrIUopxUfA30V2LnYkOeslhsU3TU
Uokz7jGnfBvyq//XdjxaA727HlLgOWLuoh4jYaQeKAaUar9bOOyT+0GNg1JmoO7Cgobu0zaoTzGB
alAyZU4puWE0qL8O2/dhC8HZ7HMeGsZYTQveUVQSzcRVitNyo5VhNtUUQio8RGar2KZwOhO8eZV7
PjvYXjRQmEBCn8qcGILR6rkLvUfbmXzNvsd83uyUoCrcoaYZCjvvCSnun1I5hcBj520ygPclL6/Z
iewFGnCu09FCfRMom4AqCljuhmWUXWgPEMTk3BQtgcdQXaohlndJcuxI9ExUcdi/TehYSBDgsYK8
efaEmCL4ZpHwwqjIE0YKx1RuHnp3hOvi71HDB7iL1xyDfUoZ4eeTE7MousRO8ILHf1IWbGGXWOQY
U0EIDSYe0wrCpVMOrrhr9s6Qqrc/T/1HAhel3ofAWTdnlJ9D59+Y35oweSC5GMPn7revCY1Zw/5b
bGNh9oL+zImGEY6c23lyghJp+TeV74JJSIBNzCIZD0vwOE2AcQVzFAiaBwsGMRub0qsxH8/gNnyY
AF0Tk9QYLLNr3PFxIAb/wNGVpXNIOVgQJF3agOzLL7CHlCO7B1PfbnllvG3AZTkLIEljEneskmws
UH4cimyyO6SPqNztIU6VeiUsXXSa6nR8Nb2iZcjB52010FR8hKOoT1cxEz1KGXssqWlhhTKVV9Nx
yHjQB6YOOQ0nIVuBK96ZuJoT7WoWRHSiaDx1DvA+mG8nht+8BaCJmQAWrxfb3PHa7Wa3k3BaObjg
Q6L9Kpp6WNtz+/tUUiDpaMkHZkpd2dCfa2fyB6gWXfSHUOLsDmIeaGA+xD+wfp6cHuStRHw/1rkg
NgHSluwWUm5rVN4YgFV1fQjmd7Ni5cGs8+blX1jIOO/1OC4ifx4XQ4qWoDY6tJcudj8tD5M4MdYb
Sc+7/icdqAzPXMHZTO6vccl37rDBbASsFGDawIBZ4TkbTg8Pf+X44IG1VESU00mUZc5kVUcy+67n
hNbclY4lLUKEANEcj1SPz567Kzk+umilsBhLdqHg4gZ2nSRh9yrkrrJvMzKLnaTVOcrBmvlZbU1h
qN4VeUfmimuzSJdzAy643dcJtBxknv2HNbuWXrCZHAd4LKzUT/JKbbP1Zk8NS01h9b0Vm/cNefdl
7sMX3BY89lXnZdnNZJIl5XRHz6JkkGukyTTCneHghBLixOxR9IJm+u2gbfXa2R1vgneOTJ6qwtPI
U0wfhpGCvfcJ1qsM8AxSX2a0FCBIOorD6ttLSmp/SgdzJ92HTQwpAktOL2RpbtYCd9pB5/t2e+At
xBOhEVnCT+G1iNVQh5obVFzzpLXJo9nxYPLH5nXGFaqr3w0OleB7N5Zw0aLgnsog18cLscjzxQbh
9C5D7EStOvKJwr21xIzQl9ObdDd5vmatAULw/LuX8xzrmsGrYGdZO2Zyen1/w2V/ONWLI6iVk2mF
CfADXG1B12rQJohSa9oY7gphKfcFXAAzEEMCgDWyjq68ZZtMIBvgWXdIPTEKxXO2VO6W5xpKstDi
IG+mjz6YBRkZj//bcrNTPN/3iUCCmuyPN+lMnC8K5FjUKxYGhOKAIwwSTtNQS4Fifo2ati/zNhyF
dMVmeeITypcFBxKIAWBAxpSj0bzok8HvmpdNeQx/YRt95hKWnF2AuFRqrkDjuYnn2/1CEgcgT40Y
rFXrMpxIvVV87+hYgo5JmyqQsBWm0zTwnGkomvkAqT888hg7o5tC13jS6wvXGlqAYOBVmi/dXPOh
oJ5ac8DMMtkjNgeeRuoBWMLvyYm/YA9LAZYN0PED6g+9p08uK7tiKxY/tczKPPKeLUPDVueiidGb
83njoAhWmAgZBBI9TVsYHyT+lZIVfcnZPT9KRH4ofNV1HhOHyxHJt7KbsGTRNm2HsqShFvnP+xAO
f1hrr5Uoi1eGYIScfPrritzi1gz5lYjaM8oRRMWjiUcEFRiEGCwSv61qrr8o0HTTbtNpOfYFkDzH
Lo4Uv0XuGMH3D3k5p7ei7grkkz9SS+c7j0z71Btyh5tLDs5Dm4/t+GiZSJ4RK5ajiczbeeNfpPEx
j0+3yYqEwuUsBOuRv/j1NpIjV04euULdudq0TvGeQUkhPkE+n1Ob58YwP+jkqcDqkOzIG1CEscTd
MDckQndKPzmfBaPy3yG9TnTYfHNMtELUHaNsAV1Oft3FGLpOFOOx38fGiH9xFkZgc+/qG5IYYb1e
kYXhKFN9n5B/NrNfVi3CvcUxhH1Jlkjhn5PhtU+wKyTj5NGNUrLNlz5PZZtXnfvChVyX0sTLIHk8
NugDQzyAnIi/RvWedGYvVMt3gKi7/NQLeBGjvCanT58vEIoeikpjUcbLqh3EXGqjf/otmGqYt6Xv
y8W5V4GwP0tqJ53hB2jtP7B28eIgAMfvunzbKUizGGnSH58mXZn1ZtZgZq9oafcNfeJ8LRYU4WQq
WHD+6eEVYTxqkf/TUsmAAMCJ8IUum73S4dSK7EhUYK/XK1w/Lk9mWBPnCwOe3/4XXoVFiOIJlF0d
/D4SxJzIjRd6Sv0PCgeL86AUN3wTzeuTG1h3b18xmIBXWSie8qbLoZOKgW8RuOVuuNnDnPibWhBj
rzFbL+ReBK0mREKDeoinlPtrRSjG9NG7si+8vOJBUGn0oIuiFElohHI4F/Biz6FUu3kYtlFuFOy5
w2S5QQLUJYfYu6wvzXVQdNB0c2P6En8uuPlVAQjSd3Y/GoqEsSA85iYshNi1RJYYDajyJD2UteJ+
8bAv/ooOih7l1IaP5LEvleOp1Y22ezRWmVQ2G5xsGWyMzfqxrfJgBlraRmQygxC2YUEOusoBI+Vk
WrnFTlOVKe+AOqXwdmTPLSdgXdn6Bao8SoHMYjM7iyG44xkx+C1VpjtToh4JPgcBH5J9M1wbHyiJ
b4QPeSzLCfuLwUc47CaNBi3SVMFoxGFADFZKnZWKEUMqwmh17etU8dUyfVViL5oLY4MrxUnq0sJC
DMdRBonBbRhbrv4VBs9fIHKbo0FhOgmG/fiLQ7pzBl5B7fFQnGD8xFcInRadHy6lnfAjnpblM9EC
8r3rWQha9wQD+41F/iXKAkCD4wF4/kD4/WPoOPnVV2jM9HnO/qyCqyWLM/3tEeeuRls8Jf6Sfvgd
EHTRwFwUarqIr+8EbHbn2xKxU90T6h+MwJco/oOOs4LjOQi14gH4s9Jql26X3K4h9biN+ZZo+FkS
9Lwzz9Wu6DigjexaSmm1nbn8x2+ULT8E2AwLaVh2y9wpz+RrZXRQUHZ6tRJ40Pin2FjJgF+o/Lar
HH1pjC7F0qztLp0+vO2UD5bomme6QZGXhqydWn8XYBK7s3lS4qHftcLrxIbG37vi1caq6U3dByPO
9k5DS7VNA/a467A/yK+twv9x633TrOMwMNmsZBGLB31bc98I71Z2Zz1K9evzzENiOgBpbZbXLXQX
c9lbFi+Y8ch0hu31VREQURwzzBFKFwUv6S8JiWAnWQWygtvi/YGy935l6NfOm/XQKG23hIer3sgD
p30yj0ClHPPpw0sxE2nP+Xn9GKO1SGUEw5ZOdhtqsdw3xtyBkhYBHpyHCFEKYxin2ndqnnNPfx4L
mjv5YEZb2AZkI7irvTG77XGLRPV+9j8ZBI74U1alkp+dz6PiHJKRQuJCZVA2fkbuXaFq2ylI+shD
iPafGf20CmkcjFM00krt8Tk1TEKYEpai2joG+Y+A0Bh2YmM+SwXBjbDFGnSXzIswbuSNsfOmi/vz
ojpiIGNkhH2LAHAc4dNn09ePf292sxmASZeYOEU3WoKc22bSa5oV2A7qtZbHXDLOk6huWzqVZHs8
fXuIKnz8WupyIDXsdk+78ym/UkJ6Q7Mvn5BwGhSdEYIdYb5Cl5Qto/Nu/h/4Gn3QqKZNXHvcptfh
LQvZjte6do12DPxJIOGofU4k3tUE31IZiPx0V0cv0uuNHdiAuQtkfMADQA8Nr8r+jGKoyhaiTQcm
0sG60h0RQil4kFAxsdzX9o7iFQRFfqxzxs4FbggxLHIgoNIlkymlxOBJgW1KirfOr9eiqOKXcGIG
oIgYXdhDEtvGAOqN5hRw7upZrAMtpdv7gwk8JHPRPF9RBrMvKoDMZWI9TEhK4r1NY6jjv1bW2Luv
p90eQcld5v9bADmE5dL/LRiXDwzup5ST9iSw96dqpHSVEf4EF1C1Wq2O1JCsP9+vIVcA56DDJeMZ
Py/Bs/pvJofcHCO66qGY5rcD0yZ+P82be2OoljiIhIHkJ1Ud1qKRzhpQWbzV9Sjhr13ggweySXNF
lQSPxBV604VWRHxUEhvyVRnkMITrC7RyR2wrMlKp/gf0xMXA4Y1bx68b0zaHl7asoevnZTJiXlor
xkLIPw0DeglCrquBuabdoumXFljxV+xAFk4bVqYipksy8KSwsPOaAyNE7aiwBrsscOPyqVEWs6Hg
UjxMp9GPasPvFEbT0GndjHEC6EKMV7cTubttb+wFuvlEk9/n3TZ4xd5/KjPmjwed2HkEjXKbclcn
JZHQUka00QOtuN15Fp7CJRLUPCDSm2DPznzAejKpWU6OOmFJg8fSh/ycWgsQteTxJWLMn/DZjlxz
0jVIwY5DITFxFdQizXvkBxu8oRpI3LwYVko1fO64m8CBz+T49y/Ej/BSWCzOgctzmT1N+yeVMEJp
A98sFSM3MQxu8r9CJVMF52/0f+KXg347ILc7AxnIsc8RIARGW1cFYDYJtD02dbm/k5E4B/0AMklq
tI54/YcVHkUpgL3zeEO0yxL/yCTYSr6NmZBNt6dUERruHYxkAfXJUHJAEuKgzoE8GLUg629twzLY
8rv1xnndpITCRphPgnLQ6TQmaxSWs61Vw64B1jG6coIZC18l6vOyTmcmGD43lKNHvZVj4Jfc8KKc
ZIC7eYnKGCREEDqJzJaZU6z2px8m4pG/H22O9s7lg8jar8DZ3c4la1nFQDcGe53kD1fSnBoWDe+F
tbWwSvxz/NnUBuJV5g3Aa8GYc1XOe37Sb5KgeMyAeQq2DmBJxtWuDjJibRUfkf1OoHZ1pTSFhS0P
vgJRdgnNaOwkOrUxOddfNmON3CxkzuBBzA2cF4Ltj3QYOBAmHqewyFNW+2p53Q3fvNsgaeHDRBUN
VEBg28tLiGPM3OvvO2HpdM8uukCd2qLsIAI8lWkSHWEypOS71cpyxZLW54+Gek21LnZ2VYRC6pFG
wRh7EuR7X4GPX/Dj3nZTpMrzvsoRsI88gG4Wg12E/pXfNMJdIZx29GMuFqmuGs2yRk0GyWcJtpbQ
J11Pn7ud1IAIZdycCqA10bSN2XlDRg1un08d1YKEc9qxpJsAJ05qSw9X3Ij6rL3vaq3QVkZfaDdF
YoGjmNAbw5LL9ds9N9wKK9MxmTFDKso1uRlI8Dz/mfKmj5fZmXQdzIlWZu52jdJs04YVPXzw3vo6
Bs3gGLd/0JNv+6r3l791dHGj5+gqpOQ50HZZoTKDBXITimcAKcVQK8K5MwwxDfur+KzOu/qIh4BT
2l3jxEQ5LdTOGOJOhqfhXjnituY/mPEhrGNGRd7OFCCPx/Vk+VZhWNhloxZJAcyIWJ/9uprpa19A
G2CifmybJPClMEUUgte5GaPHpRNc80cTHpaMl/o3y3dVjW0Ve1K/M9IxCVBfLKGmov1o4s2jMdt/
VsuB5PI2etwO4GAO1bgHlPTcVGuCM4Wgog/cFqJc3RxRuaGF0oILaDD8BnU100BQ0tGlRGmnNpw9
M6rmyxPN7/AaiPGK1Ac21gwx2pOvpppjuQDajDAAot6AGicssl0YKhoFBhnud2i7VuH5nmxvjye4
KujmKShHEvjGIf7e/iKfU3h4Atqxthi11L7ylMe0IV4g4n04r++TI5Ru/Fy0pc3g3QoHvf6Rkvt+
cV/Qov98AyhEuhD6AT4clLnklrDyukqteHi+im4mAiLN7TAO2av/I+fSjkdDnmQWzigv9DG/JTBj
YtgdLjBQte3P1mBSLE+Ou6CS2k7ABi4HkCb0vAa5w8pREH5Xc2NNvmgHoCdiO1r9VrGs0MP4KJT/
tzS+TlpVnY1dCUlQu5La4gqtbOyz1hDSr53eC33a1SYZjpuScyc/MXuVNTV0+dvKTLhk+Dw7b21q
neO634g8mN8q3+2JV166Z6d4zBN02xwGMXi3UDwUoW7xusIjejM8eMasuZKo+YOQgp8mHlpk+ZBy
+9ga6mPQLvonEdCr1cFnRg7oRwo0+I+JIqLfHuoZxUC4lrtizYKX8V8CoJvO6dSgMaFD5Dopmtvk
wxo5aTuHrpddyvyTJZ3wByRUdeDJJ7wmvNJki3ysae/FQNSw0qvqaLnBZWg+PDA8lwBkDw7kOtvp
yYXGnCixEh6yYkFwPAqQvkkIqiQtGssMNR5f8gCwbpsmo0PKp5SspUAIRt5ZNo0AqIjEWXpDfQEu
VwYGFajRJo7v3VFCIyUNaQHPrQxn2Lob/mevhzQBEln6bpHv1zMuN1IjPU7AjGHoT6wDZB8YG7ib
5vMnGx6K3w+yc0Pfu38WvmZ6qrxwNnucecp2htNvWDyGll6EfXezDFtYKf8PAgx10q2rC5hNo4lU
sOun15EkQIi25TIzNSQG42iEdBUKrBqBu3wIgFfUpsOzmJiNj35MY1nZ3Y68DUGNIe3l5Tyiqxsb
xhvHTJfCLKjIk4redODHt1RfIv1idUHqe+DO02AgigOxhZsXjdzH35dwEDboehvqFtVbXIU23xMF
M97PEr+PktbZW46oXkGaoRvwHlMmupepX16I7LMS4fVjoh8qzmqSa8jpecsiUKQVLeBybwHQgqeH
akt/Jh3K98YgVlBIDilByrujPllkR0V6x16HLzWFKMxp25ZTfL6o4ZtE1B0u5OBK/v26WwOeFNC3
ksJ7+CDI0uGtJxRae1E7oQFjO89DmczbC/UGfpZcZDOv4HLN5JdjJ2oFqmqkYCfNLeb02HuhT4Nk
eiK6W7AFoNONPDXnEkFmGKfh6QRtqxLmrRKTkua469ALjmydAMpRZCFqiHTj4D2meQ4i4oSALN4A
/xXvJJndXKtbTY2sfpClzvetlRR84xu3sDeGVe3ZOCPqrv+PFT0nZgBYsswF38AyalBsL4wteAOW
L5MVSYPLzde+84x4OGBXvT4GEELjXz6HN0RvLUiRJ4ZCDQgrG9S+wdzoFpKFBHZvNYr25Xq5UEF1
ZZc81DLIjfYv7uFJmIYErcDkFhRKL526QTj7xRrcdlPdnwKSndAFHsALLpRL6DnRdE5Tf91eSxZk
DAFp5UYtRQm9wy3Pv77wYXk8SRdIPw21IooWMiRU7KuDouGFVYSzCic3md5jdHv/8qVC1+qZ8M1l
FgI+6KpfIs0F6/ShAAEsCoeoiy5lpFkLlCUV4G9O1yVp6lLtOaL2YRTkEAAM85/Lm4QQ/Mket/d9
6wI0ZlYA0VT/7IgLmY+zbEIbY0ndx7g1D2TbE6ViP48MRG9Nkv1Kcd7jU8TdongPtEWD26QByvJe
NRYcmkQycq56xYjG5/GH15EH+adk1JYrPxwhhpxgPd/n453oQVcKgmV8uzFdo+84p+hpX6k0FYPn
Cibt+gEz+JOjNnuBkK4RT8/y3u7KjlRY6+vuaM6Bp2gepWUyatrjFgy4V1dQ4bJU5i6BTt2MwiXr
N53cIQ6/U7+Ct/3Ntqq3SBiDHKKklpjjDf8yr4BAyjx2JWysXkrheGCmgitRCG9gEVjViJaD+u9b
T556XUrQDIK+8qOvPbXBiU1li0XVG8k8IkynriClNUACx1+MBdQgcZoojYjEDba+BvMRQNTFLr6F
UxHtA36ijEu/c06Hwk7tq0tDHHoe2YjymQCCP5EwlFQ8xVItsF/e5yKcbwtC9U0FMpB/d4HCz4SU
kdCc3fb/wFLuqz+6sxXOUoomNqCc/hE1XI6eYKHCEuk2PB+8O0W6xdgpJ5jo3+bG4SpGOn20+GgP
65IFr6E0N/6vg8W8RXaETY7HhAyDB32BpX0HeqahG9nEQqTxdK0bSYEUo8T0G6GQ9KJ0oWBZR48w
DeW7eCZcZjnZfV2O9Cw8EbdbH8OQh4lYKgUC2gNFthYw+fm3z31Vq8KljSPXjLGb2XWt+WIHxPIG
U+XiJRxiFnNqpcSjpsVJKYsfJknafT4DYRhLB2DigcUdKQIL3EZpTxdvVmhOkgkpEv3iibZm0suw
JPWjx/rX7fsHyT7yUPnMVki38QPQBKOcegMomg7okLqE73FR/EiU+zW9BwyPRCSMAFBRcy5PJiX4
XZsL0VeYqbb7aIzs5Nso1zhyUfZGtgB0nQ1B+QbunaRK432S2nb6C2EdMoXnaef2f9fdLp72B+ob
UIjUVrPbKWGmHEn3ocmJ6h1yrdq1Tfdob3zKeK3VzFlhvLP67LG3P+7VQyoCkgvoS6EVm4uSjTR4
H+0XrYZQp8YpzFQ3ZZ7ant/uMYM8sDli8iYeFF/j2Hvuim7W74uHP5zJW8bjf2p5G7Xl/H6Xw5ea
n9H2b7+dc40XBy/ScjSeT5RSQ0bvotz0EaYxojfnWvyX8LiitcKigAW5MjPShzd5HEaF2Qq1yteA
oNMmtqfwa+GhoggzMAo6wcZdExHI7soBOeQLEa6BWPeVCXrszmlUzM8y1p3PnDXhJ8aDgEODCyt9
qgabm/p96MKadr8a/YboZFAYXNPU1zw6bKyF3k60Ir7dOXd/P1DonZebiZB4UDPpBnTKTD6medYS
gSEXQxHXPp1DDgKbvVwOkEWnszma0J1li2OMST24K/XxNHQ8l3JcTRfsDvIDhj7ArIalRP7LF2ub
EL/AHMfEWRX+wOHA8b+JWllT3agNW5ouLcungQnwfoIWJJUUWQ0cNkvmYCStEX0LURJzeACVrHdj
TJD2lSwaPOMx3xKCx8VtxcNVVbJ7Bziq9Eb/X2hiLT8jGdEDRhry1b0y+cURmRtx8/2iVFxJauZ0
oeuo4YnmVeNP7bT83cJMUw0aS2UsSmVweURpIgh87hmCasFukrn1GZRxZchazRk2qRhR++Ufx+Mu
X3QN76ZvbObU8YKD1Aro+y0JA/7ELpwIFBlDvivVw5kUwgyonz++NbjbwepChLxui9qhWXqhV/no
+pyQtlV7JR7EOa6kj2lRJr/IfRVeY4y/gRi1w8fp/E8aX8Cft6/QC2k2lVoi4BZXmkujlGvfglzc
EZwIBTqaAH2/NLtry3zPJy9+i9MXgFrggDA0ZJjmf9IY9XVuZdY5VbPWUr6+gt/vbLDjj3NnGs+q
CHCOytn/TjJC7/hYiHwBNipwEKB/cnDbtliYC0lPFRKiOEZtZ4nPA7k8Z8oDX8Y415AofmKbdOfX
ws1dmN1IoHA95LWDfJgirkcNSu/8LRRBUsIwaUZ5GEl9YEY3TC6hGkGiZT02EOGFtxFjkPD10Lfp
7dxqHZ1xfrBegky2tlMa5Uz9bCPSJkGyFII6E6nfrWHrohiyIjp+ODCQnn5G9uWx+YjVTSQKkNYE
DbjoEMI74ak7diRphXdWDaSj1ctr3xcrrGm1dOxHqbklr2v26DTLFukx2MBHOg22zhL6VkuiQA54
Djv2EwTPFXDQCnohFKUnYIFpazU2n3Pn3Z4PTE0IUO/czfBdPP8Ls6+B340BG1WOkVltJKKoz2DW
uvijJPP9DQ2/8JvdofieHxSePQJfcEx2ceesxlqYXfFLvnT5J/QRPwa7S544fSCTNTxa51Dd1wuT
lptHQmrbF/G5vVSJSEoOl3BA8P8gD3ToY8lDd6HK3tRpexC8sVnwjsbykwgJOeUYPh4L4NKK8evC
iu3/QttACLTilFbqorO2lA5TG8ejZqnpytkpXO77Fkx5Da2XfZP1oTTSH7OV3VMEAhwEcqa/V8y/
evuEshgqGLo6mh+mpQBMcrMF7VzCvqgbQ/UoQfJrAYqqClYtdL4XO4luZ9ZpUGfCiG45UckKOoCh
XwTwt80PJUM5qCRzI7HS6JA3ddpQE2CBaruNePFZ/w46jbT3WsAbX4e12Xuy3jiI2iFozpTT7H3x
fev72H3vudb7RC39AC/fM0kRfmWhj9Lukc0d3mdk0IKRPjpJA4ifdknmtLjxXEHLmIECFDJVd66t
DOi3yVcpLSTUTcjkqXf+Qv5wJAl1vILB5uTpwEorCadzb9Eh8CZa10pyNVCi7ksMUZqPlDfTYPpG
dFt9X3Jy/i45i0paMWDCuW2CXwXw4yQjxDbN/y9lbBJWNNvYQq7q+FhHKtnTASq2V1wk8Spm3k+k
3IqZEly1kFqyOTmicUFoFclHBXyOQXr9roY9E1wisZIGtjOQzpD617W/khErFCgvRKFSLzTQ3u18
XeFPiK4AKGCFf2r07ql1XwRNzFWoe/YDt+NSC8JxXYChgbD/zuBClJjBzkhWPKnTlhx8S0NI0jme
I+stRB5SeRmt5HxSCeQgmZfgQx7LHkcK/qoJOey9dcwNPOggfw0/dZxKXgXmnC1fLGTNXGSe+Zyj
RXEVwqpIeYlHj4TTzrVTkwvP8YgSBhPjH4FFa4fkaIrj7AhgeNlQnJ/R0fWIafB6FhcUf+1Ktkb0
pRktVE+a4Wi9HpH2Bmf+DSVq9tuzVYJHZxnXBWc2MZX3tV6zjKPui3eqPyGN3//syC/AJ6XwgdtB
ymXH2rel4EpaLnQ0GL+6Perxv35OTHgIuw45x7FuD8znB1APq8E2jvpUi5HffsVAHQdouz7+N7Nr
dWR5085ybRvYUb2qjFYZtW7UcbcckdoFicedD1+8xBgXyCnvWul67QCkodpJkLHpHqwWNEwu3ve3
GMZtOmvOqvaRL/dJGKFYsTS23z63IMhHwah3bO3TdaSsgLNCvFTqd1QeQUSrYRlDf7k2NpfA4/a/
u8aeArGuXcL2VBvtVO+d214WFE2SJIp02W2IfBabMZmLx1IrvPUWrschPR8wfkKqMl9XryagYy/H
tAVS5AX2RtxE/69y8+I1PgphRrBw0EhYfgVGkrz4h928zeZbpYlXxgAvzARqkXuF9+/olpgyu1FO
SaOgigbNXE44KTZPN2KQihPMJHqcWLLfFWKbeEUGSIF/aMAZ9A1QW1SHOdvX2zudU0TAumGaY4WJ
nEDT0UlUnjDrxyZGlLajl9RLU8ovpEp91N+UGLo2HnW8IUNrannh6nXOwDwLBSLbgSxTJ2qoD8xs
4iV1ZBoVHFLE3xLqeLoAC6OZv998GFVH76Wl/dM6yo/CWlURs0E7dcKwK+O1eYXhVXMXTOcdL/ZF
ClELNIn5lysV9RVUaWWWwv2dt3c780xUumad3P0lIcxDiiRkJ7FISDjOKOatGrgztULrRXA2gA09
t2Xj8AaXfwGzm8yAWGHkpR4JPd59LfXBnNSJryVwyD2BmOtdsKQ7Pl7EwfQF7folrzzwBTaxuNCT
FREnlgZtDduUNsQOEL7UyJuqFspUSOZhk0kuLBohwQBj4nuji/W6sShvGrdo1cy+sfvKGj4zXWgP
oT2tb116uhxWM+iPRzp6mdZAdMb5nbd2IyelXEAhEyYLFeH0fOMjnJ3Tcku0Nq/sckTJ2foYY73g
k5qjTk0UsFGREMzu23ojJsbZE0LlVgb6vmzeTBfVAeIBK+o5T8s88n8Q2V8EnErvIxansDOUB2Q9
gQbA6iwq1J0SvkImt+jydFn/BERSFDPLI5jEFk9uePXjaBaeA9tImYDB02/FEHiVG6NWYMQTbkSf
K+lJHVYWS+d3BGT5f1XuyXkDyJN04BtEvV15NRw2iY0OazqfAFTN3YPA2TiV8KxQ9Ku3BhKVxxzg
yraw3xj/hHJQBD8a4N6LfkGU6hQvWOJJuj9QSVFy8gG9Q/Di0NGOCp1YGOsQL+A7AcfFqJH4ulUx
xRepNMJOoDWxnkE3kicgP7coqBsinm3j7oE+Wy46iq+ZY93zpl1LYPX3512Q/4ftJWMXIt/slxgT
d58XUsFPSidxvsbpUV6d+UPVJCV//Jgg9S7TQvkwadpBS+afvmMaNi+RLI5QoG+r+O6Y0wZzIAlT
UEBpiJTjB58n0zQFV9LcmJPRBGeyiIgooYlx95oFNEKJ1exFUhpsnNoRkrwZnZ1QMd+0JlnEybUU
FmEMlOQHevkkd+kQU529ej1Nn9/l62/J1SHVmed/yZVi5abbz0m0wlIvJ2lFqNZXs3rVKDHqIpFQ
7JFublTzknutIYIOZOx6Jc1aI7XdpHqsH+HeJL1zUwYgpzsNu6iPvQbYWCY4x+LM+fUIQHymIa9h
mA2UzFt16wTBbzfa6VvWlqXnTnqzisnxK3zkVc9x2hAm5gb8fCTwODhWMUpg6O0KfiByAphH10jb
fTLU2BEJc+qGfniRcrfMBbWUq4O3qDAyaVAJdk5/GhosiEYvLx7tSsl2+UDeSX5p1mB3zxG209R2
Gy20QWrJwR83kKl/FIihOVRK7owL4+0mOGhuFduhZPVxibh+oJneh0PWUxG+ky5qUhv2A/CPVQ/a
k9FoECknCLPN+xTfeSAa8cW0g7a0cEzWhkrCS/4YAbie1mEzsx798w2oQoYHFWE/cZaaboigPnwx
xaQ/D/ZMjG+xzTAFJULLH0Fw01sV4UU7FhjnNaJSPpGVx73RG1HyKPUGJBkdC4mGM4un4jwnEoDk
gaZg59rlHK9m+D+GsmPnwWkoWqIDq+Eu15NOPhAZPn6fWPIkx0KHBZKHya/l9EK3H1vaooX3HMLk
lIu7j4raZnRfjhGcKeIChpSDToJBUCnSbFhUcPyRdFbzN8ztsOR9Mhz5AN0381vgN7fuJ9gpyBrj
zAmGfCNlgY0+7MFm4WgpIEpsqCY6X6AnIbdE6dyAS14ZeMe5bXe1/+IW6BS+QDIk/4fNh+HoqKrG
PzsNiXEotXtJTUHz6wFQOWsPUbsc/CXimykATCABFt4Yv3uJFwywa3sWSg2ThqtdCLenPN/gjtSQ
Mpi+dyv6IivYuU2QGbH8x/ejeTXoImx//YTL513lN2H8q0KKiXH53fpc/TuGErLrF8BZs+VjGRg2
gVEz6S+wjYrovmkWxfTuO93+p/RgvYGWR2Kc81FnmhCY2bPKtAyirdUUbVFiDpc1E5y2aAE7Yasi
nM5haBWggMVrkqJkTbr0wtWOID2dXo6ZjCYRl06YLkhMG5BFB18U18gvLxdW4E15CWMVA4QDAdZB
RALY+VbcTeS4yzljuu/nBp35t40yMz5TleJSY4UiRHjfYImpfFF1zikQnHzha2jIyVBHen0HEqjE
mMgK0THkdNRu+4gCR4yxm/r5zw5Ln5lxc+JLzS/D/1AUmWbE9U1gvfY0HsF+3ewQSclck8Po9dNs
T3Zj6sDI1HIDgxyiDJ0aUhU/2FbP/J+94tTPi0rkThBJG6k1Uw9zHf3qMoFprJ5hVznk3qmZ6CFv
OfGk6/JHCRIfMLtA3xeYlFXdn+v6y500OSb7frEzGQDoljxO/GOHTvwc+YNJynNj55deLjioUFAn
d+eObra/FFkF7pAP2B7CDjIk2Smsvr8KRUY4KkRxgY1nZc8gwdijsLL4Ver4a81RTZiDO3KMhlch
qQA9VgqIggsnE4fUb3q1a+TLnLGtp3BztkjA+omsNKflhxJHEbi8NUO8rra1Jr8dqNGpDzT+xDKO
dcQHbsPfMF0cwg8ki3GyvM/zNnUrsgRZgfR4fLxURxnLRS27k+Y700+6J/79CA/GGqDHzD/NgfdT
2vtvWD8t4hZt7T25d0CsuCWUQhtQPTeYTCjcU2fXS0FHj3SBjXL6i8YlRN4eLVaUW8L0B1FKK+9v
CbrYrqNrglPVlx//hDTf1gliPj1cOgc9jTQqa5eOF8yTDwCvwjajTfkZUjQq5cqkKhCYyUDfPCZZ
omyPP+39sGgGTIGBODDlZ6tKlA7G6Q9eEw+f+kYwEHdOl7yXPGQT1NhJHxv0tk59GMZolJm71HlE
v8MdE4xbTWeaMlBrK1BelmQykA8ZqbD7ZhM+3P1A2VFBPlLfXmdQcVOAX6JEbd6d1edYtEpq41Tb
e2y5QiKtlbTHbybY/bk2tqwOzzPR8htMdQ/4SF6X73KviON/dbZH6/XUyrk0hnz2GorJsd3orUMg
zOqPcuOa7aYTO7sOyXBNZCvWA55JlOas4VVN51Ay9A3aK7/6wkUEWrf+O4HqjJWDQ5HLTtWm8nRC
LBBzS3tvUDfoY6k+iKM0UuKF+ikX7dQZO1P5XbBdb+zk2Of81CGmQGYcvGDuhm1Cc6crON+Ur1iW
7AX/T5uoTd6J3TwLpPIdIr+ENwzwFkrNLN3l5KDG/rEx8N6nippRJmyL0IwzWzwJZfkFol7ZMyes
4JDTkW9dfrwrgh3o3Kx3lkZN9zcD310DKDW3WkDjcazt+NTCvP9gdddP6QtSmgWhpy+CQDu5jbpn
CaoDXTQmbwHYCafJnV4oYL1l0AMZH2fsjbHo7FG1Nwul2PzRIZCU6VPTB6My/mubI/SIp8916+dH
IuStVMs+CbqfefY90RsZx9td7wduZ5TezO+vWIpiPoITkUiCUU9C15nnpvAEVqNbgaFpRw9ZIJk+
PTmGXXxnBEeNVblv5VKdCPRgtbebebj8KnWkfJw5HiiRCbvFgC4fL1t1Kf9GVyPlBRw3b29ZxxaP
BMrsVDVLZBrW3XCwJAB3+BnSnn0hxK6mMEZZ0PN+fAN/DqMxIU3/cnlcUpBYDJ0Z2cLXGZF5ePVg
8g0W3r7QBpdQ58cWsjcenawgjwDHp3bFESN06hy1y7jnP/LYPCw+c7iXgKoEJy42A+hJscjBACHV
xPJhaO8UXh6lqNah+R11lEdBCdSjE4VPi1uUtwFgpgb8Cg8EyApr4Y6oeUXg/1MhTpObZIM8EQyX
PItbVkwFHcpiTDjTpgqN7Wx6agZGiMW06/ecXLobcbnJnNr3dg9N+X2H+VVQJw+s2uFrWB1v5r04
xXcP5MHofsx/UAt/bHFi0vvJ1wFovrJIEOkofPiRwco9+RZjjmUQgec9hpw2o87OMQwwt3AqKrqQ
SB9SJAwsHAGIcSBL8YbpG/2mJWFL5Gx7wDsMexvD1t20/Syx103KWhZHPFJi9gDRCPXnorPtIA6/
BRfOpqd/P9kA2jK631A+UWVngQ0khuLe020u7i8GzMBRRx0je2gM6V/ylRMdf85hoECoetMfR0cO
KGzspD8WV/RI8/uH/rNiqpvlvSCgnk+oazFjqHq+LkVVz83InHvNNtgPICwK0vzyV3OosILx1tqH
/geofl05vZDCHCtN0WQtFvqyl1NPRIQ/NgB/veYQiZoAkFVOfjkO0VJ9cP0Ekn3r9h+eUN4MmdLR
OFhTGqZOXqMROxiuN0XcsHGe9505ptXiYF5glTJk4Aa+G4zNHCCulQodu5cY2NCBvvYcEDKE/qML
8cQ5EVjdQ14XFCGg+Qhk8YqpULgXaqHnpSOLI1ZwOfWGP7/AQZVcOGrsMN3v+UF6Jdk071JTiLC2
edNAB9tGCjADJh6gkX6A8TOJKu2arvBxdiNqa13B93/tcTluXA6a9mnsAzba9UJqBvXhqWXA2FHs
cJrKVTQPmNZYzinICe/OJRM46DWDEPp5o4CuUOx0x/ssHmI4pv/JOFNFOPLNQTZ9Jusr8cj+a6Jq
etGCUejZVqw4CIV3rLY6/UnCo8P43HofYbyCQaqWs2WkEl/MQYrfelXwmLSVgZmPyHpBw5a6wSiY
toTH/Pu7tOhvbrCNfQn6XsMxWHArXdgLtNtZUFuJ7qOWFnFs8SMUk0a+KXHbyBoLcz53iVPzHteZ
szwAGHM0EzX6VdURRu6ZjWmQezF6/hFaiXZAlZ9ClfBK/pfUKwcMaWQeKil+p7fgZD8HluUyV5HT
3I1qZTlGOSlkIIXDi/kUdDY2v8EFr5Cp3m+iyD93Txi0eOg1Xs84x12LLUvwLFxxrGZy0Y4x2NUg
V5YaD5Lr4EH+Oebzh58BFCqA12zyl6lp4Seq+vXj04SQhmhRbbtn5HJK/o70tHZBQpd87s+gXjJr
2G4J1UJCnMW2XSZ+i3QHNWZIfYWmM9BTg2sagVNNs0I2wtktS0mOk15gzbt0hkJiuRNjtUcDwskP
Pn+hNRPASthM1rx8CXE/5J8fPraGDSq25/tBLXjBmBWLh3IwXMYQu4sWK0wcf/8s+VERd6x4Q6QP
8+MXXnjhgabGv10oyN1MqYSLAxwfV2eQOTa9lbdAvBiaA65Ec3IPmmJjIVfXPbc4M2195KKHHwJa
d115qdppwGw5BaqPNkSKZ4eD4iU2MmDgGNVHsWBs+MaMY6/SHmGexl82Js1g3Ir5RiZGWMKwR757
iVnU11IEBS+VaHMoxFE5F0CUqBtpvZiS2G+KVmjNSDq09QyF7HLy4fkFRt1hCcnQ2ysFpc+HtP6B
dkuzgR59FPtOPgAUIFb1JiP15UbNYvMkfMswuigUH4tnRMMNA/G/ixKzMzZs7p8mesN+ThWIbgU5
weVFduZvWkHT1oFon78ekUZw+yTLzV01HVB40nAjOOPmwo7M7/gvHHj0ulPkw0kmTN+y+j0bmGwy
I7fKLIBhK3bI/mho2n5Bqc0BTQE/SV9gxxqJd+BxBNmeCrSJOV8864Fv/fOwGTqLpV48rBdFkj7s
wSOIvOK0Vscv0H2xdObuzxo8qNvaRRhFQezLhldl+JOxhRCkd9zk0iVpL7gZfhsEfWtEo0zE6w4m
+SPLGkr4gUJPFfGocDLYoCqo1U01cRLAgYsqA7UzPy5kPO+GPPXkr6VqoVIwVF/wbXblz7p2RRHp
rXK/FhSy1f6/cGCfZ1+HDpd5FBScpU+rRLRmU3/4363JZa+RX5UpW0ga4ujrVoVDMm6O6AmaW+Ai
ydrmESSr5kVbbMv+0RpVl5HPd7je6tmi6jUkz3lhyFoO0Nl3ooK/XtK6RzoEJ4+GkXYPXq4oFHI0
uk8oQnI1LoP0WufR2cKHVon035U9VH2DZeqVsaEDJIBMKf+RyTi9c2VJi9xKCNps9GNazNVd4Xm2
oQuQRIOjakg+oPShONPS7y/RPlKx3FRAIKp3ticHJyJPq/KGasjAVC2C3b/wc6en0Tp1eBrN5Yqy
2DFv5wV2Wr7J4UNFeR35wsO0IEqgzE47Dh3hLGPjZUVxgEfY9xAukMAM6xaZIl8V+E8FYh6tn87g
ehF1c6IEn47GVVd0aOcFQr0SqrkKi4B0l2Apfw0PtKneEd+RxPt7PdZhTj2hRSGmRH+Qih2R4Ded
zpxZMAsgpmiC51NVr5TMsPmdF0OXhVDhnS70b5eD6YTklseg0QpzjbfaFNqql2OAruhgmvnG+Xi8
vArCp205G0He/Vq06i2TxWDmgB3JNx0O5aTQ8WGKbo5kjpHKSzrrNQqeJD+rmjUpuJEzzz9gEs4t
10vCcdJ7QT9j0I9/Qs/liSpgJK6R+w9GF+tUYtRMaX4Nh9qPuMEIhWEiAsXzuaTpcPIX9tLX04fH
YMoV2ZaokdyOMoYMHOtumoHH3dBinQeBfuNyW6uoN7izHT4/AMaM//rS2yvlQaQfajRXS0Wj7n5w
BruHCj0vHnJh3eY2sVhLbHNpUFsOfBOcfjH2J8fq3GiS1yWTQE4ieFr98XjQb178lxwgZr6yYabp
qISob6RfbsIhidqK+8ROneZ39QvOatU+TB/vEsTrVAzHB3UR1oThCoYJ0VE5aEOrbyyT6JBSWlYI
L6WL8bzrqXsdMVoO7tlymjSqpzvFnsBmlisKDhuRIXSbHCZae4Yo2pAg9GcMeccvqIIzvRTZWMcE
eq8Flr3btNAoyuNDW3AcaurrXtmiObA0MZ+nfZcf+EFeT0SkwDLAmzOyyOjex3y5zGhx+/H2gyxd
qj1w5O6HJoA64eHiw3PdeKLIag8UOD836XHT7lkk+sEWeSc5vVFJbVu1EbBa15xjEM62/TMSNFpd
7nh84UMmkLS1Z70UeGS545J3GsdWRdVeaTVR321CMVBpWDO2DX6JGahuPfP/bqXRrqq5Ya+jdH24
SWjFTySeVoBtgn+L9gGjm6y7yyZ5L6KvAXhAsn3UqZcKoSBcFOhaTnvZwuNWbpw1aXGpATpVArhu
E1eBzryc3RVpsb2ovZAG/7QnIKDd7Wg4O2MWYDo2KXqZq2BrCJq/qTj7OsvMal2C8ycy82q4nR/P
thzxce8mYkDtI5qljGWDVAa1yYdrQ4DyMkb/ZGD0BKTrWq31RI59zF3jwhpgmnd6xcU/GKZsfeOH
JB3mNsigVRQFu2Jq8oZXN7xOawLfjrP+xsgzMl+eD+DTxOQQ+h+ACeR2pgymcA+okOllAM7OVg2U
TzD+4YyQADYCly7ElVWNJPEjGEAQM5Mw+XfjBwAY4DXqUJUYSeJJKCSvCxT2HazR1nOJ8Pzk6w4E
ZvSrWmCwIouGdl1o3OQivh09HKSCSPUlaB3Dtg1eFJx/im07/h+YLaxEIQ1bsz8mOsZ7bsrXFmK9
vFz14mBSvSHcehGLcq6S837lojSbhVT23Znh3fQr9J8VmPGXNQ7i6cp3XIY5KEyhCSTGvJNN4UNB
Pgg3ZS5pYa+6rWNKTfH+8i+0xEtrD8+kxg/BYY0RJSAWvorOOlUAPf0NzG240bfzYJeV/YJB8dqW
9egjL+PiVi6HMVqKIiGgVEL2LSsFjAbzFmBDqNmTBebrHahpaFtSE/c1YxfbrWf75q/Y/UD/GLeM
iA96d227RQzWysignJgJPU5wAIsw9GSv6rwOTHdB766Th70u+wDrQzuiAy462nCS1wRG1wZpra+d
qwbpHDM5LVUrrXSoveXX4RGjXoCYNd1xeVwQWtYpdKMLL2lUG+HioACMcYBdVcHzhL/45Z/r1kmQ
Efksh3vXMQUrn/HOcdzNXm2xgBTQN6KyOt4C3bKzePtNT+j5RV1ELu54N3rgJq3pmQfVIvAw8iNv
j0idXhA9/HGc0v1/PFUHlQJQ0upM5+g/7K2ZMspniXsfg8vMeuG6UjH+WRGDGTdDXlDU52t5+LFv
FW3alAwqtGtiZKxcxqP7AAJhlHPZpARqOaa19JOkFhRH6SKMCNHyst2BVmwS+uR1dwLeGbTKxYoy
Flmpaws4i16rb9dZn39IpaGpcp0Gdrzy1hdcq5y6S/A2agy6ZaXC7c6wTvSg3BjV2EgMuR2o3r3A
DTvw2ddwQxXZxP5W854Ld6ieJrtg1SkaoB898Qkh/mTmA+vv4w/tD3zgvAlZURv9VU/px9wqKQRy
EvCh+mTU5EltwVLcWLeK/qkCnXhJSi3m1FBcgX2U/CxaIFtIxfhPmnRZGpwicdh5+88Sq9Vil0ja
jx+dCRBXKaIpv39TccWIo9lvMsmzhi/uIz7q24UsOOJGwPrrKWG05LSlAzAeBqg32Fp6nVsvEoWJ
adTEzDtWNJjK5vSek7flxCAMrqJjDxdTnwMmx+CxEOzeZ7FCgtPfa3e4cVx243DFeHEGZ4En5o+U
ZZvoLT2YFcXVazg59Ma7UpW+O+4e7x52NaD2MD1OT1wW61feAkfAdfcZxU3BSfYvec3taKvNHN6W
Fus5a6yDQ8yToIABSa972yUdpOrFeyQVEjUwaU/P8Ft2khlo6r5r+jX1agebVbHuQpA1W5VIBKbC
76arVwau09vBwuHbDyb3WbZWVXsPoYzhk8qnxhg9V2x0nn2eQNPyth89QMN+nxmcoyRxOr74eJF5
lpFbh47bIS/oE/DVgQVGX93yQgItHz0+Xb7llob6ydPY8f0DC0+kSmd4u5jWAPlu8cmDPF/iIgcn
iwjGuiMCX2mJaMwUnnYECInPcY1BHjDSoLbrA/kD6muPuvRSbmZsI6njUooIjUbfjZAqvyWIkHHP
giaVsBk7jG5z/of9w3GkDqx+F5MSLgxdEPKjaFjsjW/1wrZA3CAycDpvu1yTADuWT2VY3ykvYuTF
Gaaj0d0VAMkyRc0desENOs7iDwEqchFPlmcOBMsTZ3ujto6R7jbIeuSdW+HxY7gpC+jkYJBvkSEq
R6BxUI/6zSHeD+8L6JPMwbDyZg9EpyOyPSBZYiWNCKcxVu/m3si6yms//xgxKHWGSQ6RG8sOys/D
rBFCCogcfOtg6fwaS9vOMkoBY8JenA6FRkxKGJslpBNDmvX0kRjZy6LL6PaINVC/5TvaWYVWLGZk
34waqt5ZK67GU+r2YNUU3NY7UVR6j6QLqWmCSWmTJWUYtulBiso0hY942xp5cojsxpovFMk1iN4L
HeRAdW+wU27e9VP9mwn2wcgx3baU8iOVoaFaojF+T5Zevcu8h0ok3pOC+OXRljzlSnjjfoOM23tV
lPXHOI1HuR2PXCrTBxMy3A/2SjhA77vfIGMkBIxZisRaxbBizaroB6xyn9PaBAEKIQ+0ie5l6qMN
YrJqbKQOnZlTS1pRbAJqPZLYXq4K7dK5NLnGwDNJzP7QW0gAoaqZAVttC4lZdmGENbiEihBuhcVI
nylGHrO/t5up47l/Q/mxQW7g7N2tHlu63wsTdqTd6Whc82KlonLoB//8zYvR2ffPKbhCNZvWYDPe
d4QRwSKaW9tDYCJ4euO+ZpATpsLe/I3pc7MXC8wGzPZxRu/5aaGEz1n1j7tiuxra9XfilaK0Zd8m
XXTqgsbo9/zgel0hAgH5SpH6ZuMufAPr+A9LwPMc+XWNNR8U1du9oJlzyCWg0gxlV2Tl0KoJV3//
44SGimB398XY+DZnitc9VvjVJ/o4kEX/ouTWQeUIzswjkfg7/x72It76/Qo2shKfpfrlXx9V993k
mtTeN7iRnKDMiXnBYebByoNVfmTa09R2MZGOTAmngjcTvE6EG7L7C0FXyK6SQdo57mAOY0BlrqqJ
Cu9qv5ymdxFmNlMWA/KoxIae9f45bLVcYFqbUGGttIrOgbHX3DMjBC+qoOinZen/1LXQpXhbWmdY
z9cZt/uKbEIUBW9KEawEz1fVIwwreiFDVEnITwNBMkBLhW1N9875qhYR3RDk8LD8T5C4gKEUdgTu
AU//LEo9uewkUMR3D87tgu2YyTZ+YIZh30n+YQ6HLVn/Ti780IhW9pE5ocZoLLK5UmEeD+CieAZV
Bv9eh/stC0+tPD7oFa/ElyjTAxHyWvwl6/rjqDCE8JoAB7+KiKHlkcCnYEM0KbkfMCCPrjHanz4s
t3ecs4zUnD28K3GxfwCEdiXOrj3tsTwKo/C8ACwZIwtHhKd/hzqsC+BXF5Q4ajxAiExAZRBZMLN7
ba8XCb2W1siXZf1RPDe5PkIEkbhMmaBUzAamkICqQMZWZ+n+QLFHvLMy9vdZAOwNSTJVFH6KXKHA
rOfMFaywsr3HnZGkC3HZ1JAphQshU1b6bTheoA6aa4pxc0YHambkG4ovgI3WbbPhwdFC5i5eyOhc
xW7WehfFFy8WMhDo6Sn7ZiuUnLQJsc5mfTFilHeU7swVgT6b/l1ujrea+D48W40D9/5kPSJsXcsZ
X1ihDIGWIz5CHeY25xi/fj48D1lrnXgMwUQmX/k7lo+qRHX/F0nUg5Rw+HM2gAYMaVZM5ZAUg3oF
m9/nnvtsWb5dYN/QH8DlYxXPZ1nfChPgmaCrm1vNwPV0Wl9giEWGMvLWhaXnsZ0iZAF66dlFm7eT
tmdYqkIV51crQl4PqkRsj8vl7Mh8O5xJOHJl7+L8/C8zvsO0himuxQDqYjgsONh2q4QlRi1txk2e
oLVNgcUtDMaDPjcxEfg/5u4ct3BxuUe7rCaecc1kst78z9t1lieSAu5amnIdcVgMdXS6fVQZ+xbX
6oBok+1sQOSQ9r4TPKSHLGSmjYfM3e34EbAkGwvZxz1bnXluw/L3AgutFp8MjKhn20sHp0EvFl6B
XNnSA/dXd1KMMPelGYDgLtEI5GL8ew6aHbWEvK5+wx2T8kNwV7ATSpE1OwMiSOf630h0wslN+wdz
1IGxngLBxuT2T/4AGIkQ76VlpSyZ0kpUZzHlYSIjKIJRyu9Uku4dh2ZrSrOv5V34F2DrCmd2wBAU
ipb5hK6n1JvFkexyymNCNi8pLFEaRNdKQruGmN5uuaETsTRucsbDC4x6N6k5xEsRr4vAN2XEwm+k
3iRBO34rrudWCf1h+gj7Np09Kqjvu9sGmryOHZNp3jSU571kQJV/D65vpN+ww0rB333pgmwMTiPn
fOgcKok2ENESwosHM8kWlDPjYC13PKLelw/m8EF4C2AcWmfUkYR7UAuSxBOkTM1nKPQg0HfqEAZf
4/EZ12lqOSRvGkUtPmxhBSrfbwzy2QJc4B/Ci31Sl0TsCBIm//ShuV3SVkn02eex0DLEro2B7SJJ
LO3DuWz5GnFcIOiKk9QVkH0VzsHgMyemlMmoTCfxpdWQKZJG1ZEXB/1nD6bY/wnEzSPgC/fhXD59
JV4XXdU9r5LUxDLpuvrIa+zjMIPt2ytF7Zk6H8BdQADJkYxkbiQvxc2SuodA8FZqP0Wgqc/IUz8Z
WBW4BHKQeiyAaAeglijpd8gqzADLvrdXfpg38Kp3eVjkqgKtipq/FYZ6eoakWPtNqRXFPpAo3I5E
JE5cM26VehtKcdqieTG76bGJIxAUC7ewfQ8r8WnxCrTqsKT3wv4nzuBdLXN3aeEAXdK0LOg4Yz2b
Z9kqa1jzH1lJsH+7wRaipNfaumxiX0IXcgrb4RMh8b0Dl/worYV8wyGxviTRerePdLqGjQIviUoa
XaFKBXioyHBtYpxV3Be2uamft6jMt94DaFr600fmrHpugoEyrFTG4kdXL10klw0IerBzxSBTJffZ
fuwP/g2XPARhHJjNfd7+YHORhbLCGOBeW2Z+VclQ3BkpkOcBy+G0kJXqA0X+RWmXw01IDvK2Ayrf
RHff8vCtEdGqPMytLRH8NnVMHhC7LY79wr5Xxjqu0QW4/GDn3PgV775qOv5rPL9jOTe9/xn699yl
upRTY4pV/2Am5JMKj4fmg/djAYykUahtZ9PQ0mUXudjWNfXJRDxiZpuy/JhuKVbBn/fL81KVPddI
aH0KKm3lO0sklChqjh/DDmklUZUrFfGXAoaykT0WtLI5ecaCKvI8ReGDMWhNdHIr8KKBJWGBT655
NeBPM49AkK9EP6EvpS7Tf36xPS2CBZu/d9Mje7scdBBacP8wlcPI+qz1Kw7RHOua1o5u+EbZivqP
lfmBEu/ZQ0DHO2eG84HjXqkwfxhToo7z7hn5euYWISmg8jPF/WCH4FFPEB7oMmovpWs5atbfWjIk
orQUvwUMupP0rTzmkM4+UAV3K67906aanxfRlVe4AiYrzFKQuGyKoNAiNGgmTifNrIJ7A07Krutz
1G8eFeyBZgwXEW+iTZvREeJb7NY5rNpnIPzDNUbF5MUlUIBCQj+nMLrkrPrfYjCYnjq90gxm8Jb9
98Nz4fn4tAYqYg4+FuEXXF+IzUMONTRbk+jo4fHJ1KcSpm3W1CyIugh/czAlN/CXeRmnaiQPdyxg
iEn0eJ1K+oDMCaMprATvIxsu+KOnGlAdc0ZiJF1jlEg9uQfxqvET/P7ba4snV/23ypCEFNo5ypla
GL+Teph5n21ruxKIJ/Im5BhJPKlnxW9lnEYntNjLfkv5V00xymRN3wuslAqJW3v+n9y1wXewfrLK
tWXfu6rA9di5joeN3RKk295nd6ewyURs2wHgHNZU5cpk/NquIMWDM4F2AfuzB5Inv/hWLO9+GdLd
l8coVpXw+RD8MJN+Ixyk8RKcnzNYtl1q4pAd2+BlIP+LHNmLE4Z5SC3qlHWO0QNebDr4NhlPSKWL
XuDVBUzezPjKxRLlasVxeTARAN9fSagkwOrD8hc5G0EwoNEfKSLnXtTKl5ELWHQK+BkA8vchWZWj
nKfLThONW3NCRmnEEv7d64t0/UNC2EUptD8tKz4qU/+Zg+SL9aLSG5ugUAbL8+77zIDrzYTOC3BC
euz0bg19cQAFGARybD365hP7y5wRUw2M43omgEh0SLhatiMy298uzWSgyftbsfeyq3Zd30zdzKsm
PH+zHXPaMdw2cM5N4hrR5nBR6oxJ4KbVVqs0e/uRxVUsHaTepvvE/meQN8lJavVBl6F2hfD/R8oZ
fRE2kfh2YSTZoxQWVbkPfHPH60SVag7I9PuCxKIWAzEMx9uD5kF/JtgRt1VHWmH7OcdCGevsPkTD
C2ijD7o0gNPbGPCjdfm9nnlb5ycgzIsrYTyzFvis9DI4147BUvSTyyBMp9xYBNQK2VREAyOntfnn
AGalJiAsv56qDUyVFM6zgpqZQsBby0t8l3PlS27q8nrGeKM2+7S2l5zsZQXEBxRHmDiAFFmKaXNM
r/3XF82QtQM43y70RwnLHXoKL1lunDXIY8P9edy5e6eY5l/0T8LU0F2UlD/wX2f1tS00K8sZgtqV
oQekDpe9YgZ6bYKUInKdbTCbZORdO0Uo7qA7LecN1Z9LMTWgpFdZOQdoRDXs4o5aj3zrCjtW3103
oIr5tLedc0bG8dibaTXV343YC+rEFfdq3e6ee0ZR3rV3Ey+gD/S8zGwlfpEIwVMuB1QQ5baY4X8g
l93cVhJRx0b45+jGJ6zcu/bqUNzh9/ocPjLxKwW/lenMxS/OcCarJ83+KCWgjjuyzI5A0+4AmKdV
cP6XKOTbzFODJ8GsIuwnXlSxcTz9x6yUEQUNzsiVUSI+gJur+6wmGvt9aTBy1GQ7Gg2gb9iYGtW8
xWcyzHbE/1u0hdUFaObo6att8ChyFCX3xqpRM/cJRxK8vWARZWVP0NT0uIEHBJLwxzs7HXV1DtaU
0l0xNOOoGEfvoatNyaEPjOT2BBaNf4HixtaKRONS5FB0RVTxgNsxrm/0dBEAKCMClFQzlhZv1SJT
LhhLqT8TzIwTWv9eafAW+QHNc7hEvdy82NAzSo9nMfFKYGHIJL+9IUU8e8jwjRUHkhwY2LbGsa8B
wyJLEeh1+vAlk7v9BORVY3uYqIQl3FrxvxRGAxn2Vxe31uTq5QVJZkjFf7jn0pQ3Pk0BoiATOu9p
q438PxqUyt74xxA21K1dSTsN6cJKpLwOf2fiKMZMJEI0vyEOv5UGiPeeY3F00enFqAV8kmqEeIhD
tMoouuy05jQUZNLmlrVymakZ80omh0masfLEf8tG3/G2H9V/dxXUJobojPMWCRiVpztm7NZZdo7l
y5ltCkCrpvlJB8zhAZDfjA9WWTy53Zh9kTCDJoaA02EF3BEJwyWXclxV6SuWktTJTg1KugryVlNW
uVBLhKEAuFVgingy91Io70Ym3c+pxR8+9BAcISvLFuwG97BhDoweil4i3wlfW31A3sxU+4cONnCJ
6UYEWVriJTx9JL5m2XAUEIO6ydszFAAy4q4AwiGyLNC42x+RIdjrvx0WPPe/ltOlZyyJVI8JFpmu
hX+BX3HAEud7LUEkJHD9KTVEV4UESzF8kF2ZtDzxYaAmWzhdfXnjDujDngzUIdxyrSmfIqhMTz5Y
i02Uxj5W9sJt+ssF4r/wBS7/hovddWoz9bG9MQO7U6AYazMdKTgIMsrOJUkj865eAEBAt23BqnpL
6H/zYZ5PFWI6xLOyfMXtvndoAmS2UpGfvMjy6/5KLRIfNbxPtq5oMVaNAqYZgMOKsrbYr9yqYHcZ
2Hv7heUjNTrh5/cYVDSyjVKp7aIliK35FL3xnpWecuCpNwAQuWIMUpSrivCpMaXk64os9dK2yGre
yai1qvcMkfLVYiIee+8y0w/2a1FNu+UbgOId4JmJqm7KYB7laaISfA5551Xyw5QQ/YKMG6KsvLMU
iynwTsdaZ2r8DwXaNWiikgSzst5GD6H9Q/5BIJ3msZVjZVWg7TWlfWNJ/uhM9K3ikfxQfuVdJwMm
89J85U7RnOeSlscNXv2SIOxMQpMTdKM2NzChMasxTlr0gTvVichYACwQPVFFbvzoQhyUjU4IaEMY
bJbQPhzl/lYghZEu/AtmhgolicUTEPbwFo28sf6za77L23nFiN1SCEu8RGeDa5Ck+zP9XXl/QbrO
rDwekk414j+QZ0PgBZY5L9nkbx+ompHj9lnaZEM9HWdh1TRJxt2csHQlq54f8lFXlIRsH6vICim5
Z5P4BixkS7x8mrPyOSmpj7qs+UuViMu/pvozf//8VL5CfSml5p3Jp6V7/odxv8dElDr2gNawZynA
dRNWuJK2/YtxVyRGNjbPIypKoZRGS0rREiB5Iuby4eG1ct5CKRuF1xVYm1nNCrRWWsnl7SsA1frU
sTTuYL49qf57BQM+8GNbN8SdOAoJTmUXmtSoeZWpwfmsm6dYvu0yM2YNjYs5O5oyHzvcm2DEVZjR
uFyjGyuK8YGo2HEqfmcl0tO6up0yNmcl8mRr2LLcICgI/tOnbIilC1F+wydiWomuwwgCjNBpaOdd
5A2GcFCzaEIQ5BIh4aikO5nWmYk0Ri6XN6uTPPo2wdJYBEXhU8DhMze7MgLfXoXjvJ1OJbVTS+iR
ad/aYCIQAe043dY0D9QPZ73eEm8vX38+jwrgJGy4j5GDccscHrseTljQtozPP8bS3H7wPudn70S7
VRG9+NnC0aLHPA7GvuThFa18xcZ1QsCDTyKJ4+5q/p2EycbxSENqOK7WahAr9Ng3eueSQNDO6DBb
+dBQdO/vJJaUxBRQdGzKe50NdyPSkSQMtIbbqZz+msL7WgAP6Dcmj8v+l+Fkl8nZni21BaJ8tneV
Wa4leRBgdF89EC+Ma5stskp7MR+7uVlPBRztEdtGpYdJJCqeX7kg9BJtz39PZuSU3UmiC6LSNudD
nrtlC2J0FlZifWG3BH0iGq1sL3kketomwxpikXLj06wfX+s08xE+vWDWnVJg4ain8uyKg9Tb/GBO
x/5yWaGLhFKO/m42cuepUkNQw37BEPo3OwmDO+Q+PgJcc2vr5btMil2MHr6W1RO01VSSb2oh9/8n
yc5cH7N54gYUPZ0kCHQLTx3/wNGIzaN1bDIUJ85eQlo6uNrErTg+
`protect end_protected
