`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
hOu1FiMMIYi5J+/YUdXFl954ufKtSi0tHn0BIX5c/jJYC1+Ru7xLDEfK0dGSL9SEJ/ZHC0IS+6sp
eFCdOmURkt9MCETXZExuqTS9sEtIeCYVkv3wkN4peODvdPbcrlyl4RnLWmPawnvHVG6fkjJ2P6Y1
f57WGYbiLr0QkyeXf1p0HZ336ijdQhQ+sGen2G3IHkTpauENW//tIfhoHeO7UeOpRd234qrNmlRP
cZG7Qd/eWvYEyPYnZupDXq6XxJjhH7nV1dB9+mtqt/4cAieTdKohvQIKDC37B25F/h8I7Pwe9sul
m+TWJ6dVtb/Jxkd09xSriaxFjMd08cBipMyxFA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="aWfzia3LR7chnL3lBqAQ5t8aSOIuxHTibva+Wg8scjY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128096)
`protect data_block
RIeccM2Z3cMNBWYzMNPtba9fNIjDDYv0PIfecPyfJOZa5P2NoTLQlOktPnxkpVHXaOhSi7cSvosz
GcF0q5eudbwACL5NGTP8Q9E2evAiXIrfs7h0LnnqBUEHIkd2ntbQGuY0ob0qK4fJlguo9YHwYplR
8RUhYslFgtI/ACxO4fV1So5IkW0+bVAYoFnZ8Dp7GhTcUl2v0fgANOT+8L6fNA3Oi3fUa2wIktDV
5ZgSovqPo551Z1yh3Fuk4Qti7KtzCQZLYVPZhN2j8hfd762hAUMeio0y1tLF+4tw7yP0BuIE2v3d
+qXMZ4brCy59+EJa5Diw06Wkl2mNvnMtF+4LuRfR+4rDMndVWYmzvGxGG7gRPjhLKaZwc4bKbyck
P2S9YQlb2VdrAa9BPoOe9UjsPXTQdR1/769MVZvJc/LAka5/XOPlTiISGv1ufASov4hSAC+Tkj1K
x3hB7G1daQhWUhApXlgENpOMq5L0/BrPwMJ10Uxy8uklzFYhWCHi4QxZuE28Lq9V09aFLFRwThRH
4DHMcqCU07ZTrlW841UXWmOtK3/xGSMO+Gf63ussqH5OgMwHayHN8rBpmbno/ZVME/LJp5TG8jml
GVY+qBMEY5/QWrQG1CbLUsditZXJfO7kDS8aUrq/qE7zt5D1vGKEaXYvGft/2DJZMJ2mMi1S3Erk
qLr1HhY9CJhNMYKwsLF4TB/KFgLAxuPJPPFrfwK3IpUkbn1pYbZmVeU4gMNIGea1pQFvoVWEIgkJ
XhMjQxvguVnSi9MLcAnrP689tBHgPIfK2wU+NvR1fGknHBgsVh89hrFt1rNy4KLum1DNX0AhtPTo
7MbVqAluMZe0e4CJYEWe/s6kPNb8UBRlavYv7rtvYF02OWY7gGzWmg7kfDB8ZVr2l9zoqDP/7P84
UR6axsljn/s63kA6PZdLrmDi6NXrrA2q5i6ekr4aDqCZcOAPmMywUgaM8RVxMfvwN0g9DV7wg1vW
aoK44D5MbH5Wq4T1v/PUl3y5OCLpU0/Jcc9Wj5t863q00cz5uuLC6tDXacbItRvFxtaZjQZf4FO0
Wy5Hjkhu63OQwtoyLvdaweR8F4o+Q0BU7HXG3Moi6inJuifqIcYcvDFpIhrdig24CRRiOXT3hsGh
bXkOyzZQqhCNPNawbE6ImrEHHFCfp0EhU4heX35tpuvqxxasDDo0933LBywMpd6Wtku0v8EeQwN3
nvCRRCjTpVUr2kLjClx8qRYOyD6+X3qALuQwv78EVge4iu8Q8l08b4TTdXUX8fxbPxKZKJ6OxWwS
F2m8wT39BauqNOGl5R5vvNXApyCn1MyaMIM/fEXb+i38BprblpvAfK0cLJkxTHoSYwy4LtZmUz34
vG/5eWB0XB3SqqIPNp0HMeiytcDdPiFCuw3tLrKL2TrhfZqBSlWZyqHvRzbDvIQViEVLqBwVkado
EjGLtbYC7EREifG4ykCc/+KEBhIJ/EwrMMxgT7Fim56vyzqWxTbvVrlNkqfXGIz8Mv7AZAbGViyr
t7pf9YtEYLqn+LQFHO0wU9IOH31O0ORN6OS0GwmxGHMVy+or0RhuNlFcrpf6wYmzb/a2CAno5yh+
uw7De/FlA8uYd7WYiqoftb7bgdhWmFkc87+JKaYnGQgp+DgRZHa4PKyDT8tR2HTE6r7VEgC2Ws6T
90jCiiUt4S0HvdPN/M0oKhS8V6+8FsZuO1jlm+371woi2cUBy7Zv3sk+m/lVel2by5AlG99ySKyc
6kZ7y/Y8qjYP3lNZl3/GMOWz6aQEht/slutetolzj2m+n+l2fg2/AUJR0rlg/gJkpL4nkPKQ4/g1
uk9hFht9nZrp71o06327XWKhBpG10mQH6RsBi4d6mnPQXwitudmb7KrAHrvlzWNaY8iMb39LYgFh
IBe/GKl2AzXxG3xBRf0Zhici10yXNqJRnJJqwGALiY2+vSH1a1+eHs3Xyski7Y+ms0eKKhbHk3Se
euNHDrx0ceM/hOKhurTnAo2ml42XUnTUkBoVbsS0AL0awgT7PJPr4GkPpcx717yu9pAt3zwhTJqZ
bcHpLkHN9wurCSuFeBGIVht/dE6as5ZFrUNgfmDejD6R3KvdImQAEMkGEtAu3XJbiwRcW1cV1UNp
Zp3MEGUMPH2iueJKQV5hsep8MwEific8ledVCn1QrgxJ4JjZFqn7GqFKLaQZSQoqzW/I1dsRfSwZ
nviNt6WvWRhYLvnIm+2UrVYoSO/Tcf6HbNyz6e0YKJiVRCxqnpYQZZxtAhzrYfiOzeslu6pLigmr
/a+8xbWWihunImqaIRrmAewNQFpvQsZA3trIWHJ7AjbV0xl0z9zKSGsQG00Ey7ZMcIESUwF9wtiK
SSyqJ5wxb16NNoHRL5aoD9XUpaueCQXFjFbRYs7JUjpLY8x4rKsr9Ovk0hTNXXIsrcaAEkweI+0R
BhXJC/ZUf0mrSzmX5k3swOVxVsndlx+Z3h1a0Tzjm+9beoJgvPuORZF4YC+wvyPcF0tnhbCjDCTf
2+F6sfpeHBOclL/Oj8QHtTKe7A+zlwpKDP0mcU2x8Am3vQbxub8WE5XqeXcSOe+XbfMB2eZqTI9a
MDpQ1/ky02Wat9Bn9h7RMmv9BYJaDXXfR8iY0INp9SWbIxnWbiERq2M6U9AYex/9Up1djnwi8tB+
rYN9KJZNWDmVACA2QrdmQhp1sCZBu+rzc8tMHv6lZo4QssjoIrnjqKyKwl749j9QCDSkUv/xDMFu
iNdSo/KOjEX0K60QCqt3W5OzWT2FzK8+kQqxWPROIztylzSiS20cZL84mj0TcZPpXiIeSgwDjp6t
aXko2TaRYdy6VOsoxebephMwg8B4hM8x24+XANFe8Mt+Hktw3RYsnAldKv8Jax7e3s/AFTIRpHM7
JqRutTj5TcqQv2rIQ5T0NGhZEPWOfY2XNLg7Eu5VLob61Y9gbgKI+9tbTzM9aE5r09A8MPfAK2eE
K276hVchMldRhKuimGjVBP49ZA9ZQhmHorM+KWNfLDPwKELsw2s5M1W/rAI/KSR8JmAzH8oy8W9c
npTQnvADWVplTS+8Oj8b/lGGFOW6dUxxWjAJMpnKPXZwSbNH8icfrhQMTrppMIVqPbTjAoQxuQpo
AIJ0I+GGi8a5HBE8V0PkhA0Sc54D0pEnErAF0vAdYHqHTzEQev+jmgeFxP2WlPK4yM6Nx24grpb2
qAnKmqntQhRu/0opfI9CvZgT1VoBfmpn7RMC9edWNHe0qlthXzfRPP+/F7W+UOgQeXLtL2U3Nw8P
xf5RG/4JqYZMARav+YoF2wXf4kACDb1bUfB+Co9cru2O4L70SOMJPPRV8s7FYOukURY84AUPQPoH
gGNLoUU5MgojAPxtOsoizoyzP3MGwyHYGosq69bxUHrpH3OIB87T+QLXHd5/fXmCffK6U5kQLB/0
lKPgvZKqkYJBjzXlSvLdIowd8tHfuiB5w4XwygR/gtks3MsjhgSZXUBQ6GRE/rBSBGnGhqfNSkDd
IEuuMY3ZrgTALqrzqoDgcEofB1fjT0Q5/I7A+IyE0xuH5T/UBe6x66UOTuLWycLlIKUpj1Yb9eUy
gBEzBz4zeLQwhVMXvWUD/Rc2fhGELiQHu7wJ36vsS+nLJ0eyTYYBBvKE10r+hGeeBc/+AbOQnqgI
49HoMa++7FjnFXKglb6NFzNmPrZrlKjFl8By5YzUwr8FqWxV+r4mFWc/xgZwFyx6jqmRt2jQQjsp
jLBEnOpM1Pg7rXjuq1kOactuGTsu6E09avbd6q4fegjbsPsa+tC/BXg1TOfA7Pa9gYoiiu7kuPrI
SUXQ+smOmvKVbz5PomCu/hwDToAJ1qtIN2e2WYgUjaIniHBDDoWJjHlAGCMcnwwPr9FMl1hwbHoz
Cc9vD4fqnj0Lb7ahayx+89INNZpK03XTL2DXlU7RC/aEia+L+m4YfGvr0g5aQgREynFvM0okp0Rb
Fk4HCIV9kOUPfVIKoTP1Rp7X+nV4MltSw1GMPH+bMGDyDwMaZu+5PIy38brKVsyhbVg2RK2Os2+0
eaP1Q4DKBjSqohVsQ9CUXfbDW8JbSqhQLNfS+5bvEeKK+r7q0KNmpBeitIW1z8MKM6+F/1XO4ndE
SVkJt6pyIFn6EoYujioyLS0Vt55+etD+44lLhhjEpH31HHmjnQPp/eMoOGqCPfxrmH6EnbTJWdRo
hyXOonNQy2EN+qZ8yv0L26N7j+SjMKEot5zVQI8XhiSTsrx46nDj0S1RpIICDacro08e+RVfqnQ4
PYtVGeP8fHdrQHzjDlf2kXeIEkbdEAZp7sVUVAgEkwIR8pnr8Q6PaNwPvQFuiLjPZDBfPcmx3Ib3
RHIJga8AevnE3UFl8+Ut7bFPjz9ZQRX8GQqyECfmza3GmDUR8q3IJm23/Rl5gwow6AtGdK8QqiN1
kEhRIZugEKj+Wgjal1dQxgjMK2UtjKLVrpz1/6iTo9LYlUKu+px5RxzDHgDuK29ap1Ux5rnwrwjL
Ji9C2a/MeUPTyz0rAcmhEgC7vYoc1vA38rGc4xZ/zJ80AQD5GH5jupIqdHEjo3Zdo77uh7qAl81d
Tyv2nd97Hhcc1F9Zrd2xLtdDjRXWu6zG4EtcwemInFsqKfVeLWiZZtrXu46ywb7I0IEWHhoSGY44
pq8ASBoz/mwu8PcGnVMf7wQWmADF5rAUzA935DfzYSXnxpbxXZlDwEHHsgAm6f5+VejofrEe9maz
CluMpTL5/ySYuGKnvWTb/ZN7GcGg/vu1fIJR97FYPXftdYLBFEQVS2v7VGCFUKIED4hxVvBgZxwv
h6YFlrA4cqKcUQvyAdMaAkKJBpwopbCbmtVQ2FeZ1KHmGdHTAAmh549bvx2Xp8n8KEZSWBoWjwKN
BBpqtPmqfFdjiDlfDQAhp/nmuKXf/uC0RfJLy0e/3W3YOnF2iKvypMSYHW+LF/AaJs000PKYX9wC
spjwqWoo9iUHcjFc5LwwNzPSL/WAYWbWW8ByI9TyVL1WmkKOM8OUtiU4O6DXsYTirCzJhBmzXXI6
xycrYeDlAor7OmIVmvlXAkAy1DFaYXgCDqXGaWjAqyBOrrfdlFJ2ffuVhyTexjT5Rp1iwJXtMQAW
6xMjEJB05XWhCN4YKg+oU53Pc441AWuppl18necXCgdwei83c57YMKYJorOhJ/CJH3O+TOdXwfF8
9uuSDh/TpVw7Q+Ptw5sAQkclAkN5TSX889NKCJUm4s5JykRhy17qQd6aA3e7l2dHj8Zvl2zBo9ZD
BDF3jM8Rnm6erqOdMauGaOrSorCjEvC4iwa+IT+6AQJpDXRRH+5kFuNVQJBldYLojk4NhQnpC3NC
oxvC6B0fkOa7UmQRVlqVMHRrfEv/l75Ck+s/p33D+0vnsGxiv6KQI5zytipJtjhZ3HcUUkvNfIsp
wSAcdvNnXW9iDPoMi2HvamEreaBFOGtSdkUDxcgKWxn+LFaWI9ynK1nN3644ZnTM2yAgf5pZLj00
EPZ9Zk/wZEL1uZ5f5R2+SaL4BQlNqgJfnOv7EOX81g5cMDNlc3L6SdDOLzcbbWJepr90uOaLBgyi
UbMBgPLPm0lE9mqK6/JHyo5IXd3esIf9QSfpSinP72xzkUcfjdycNOFhjXJZ5u382fhO2qXjMtLv
rSFlRy3sDBlBPWHI7IQ7cd1so6mJa8sLBRytFGMMMtB3nvHVUxiy3PQ9MAe1Mq+ohprerTu10irt
5wnM7IrvHt+boTBX9J9jI/TVwKZ1+uWfggvHlSuDBWMuPgm87hCzvwP3Xk/P19K3hMVyRsppxlk9
pJmIVHlh0lMsQreLghvLj5BW6vppvOVJGLsGyRgQfh8xrX3v2T69nFia1JpUhdQrI07IJ+bOzMIo
eBhx+citVdDhDULyhYB9i8zQF86Xqz/IhAPo+8NgTSz60Fkywb7ftCZffhjg2Droux5ZbrCfk2kk
QCMIlGSnk6zdBUk4cQrJDuuxgszxSlbv+9er2flDnsT7FwQUMuLIXSs4fhu7MYOg0TgC4haXZt8r
5lqILoWBne8wCVkO+0gp1LBYpizIixYktH11ex00aD9fQuR/Njmu87EWzwyHwdVhcqgTnvQ3rDLP
qlUi5o+XLoqrrW+4BZavuUwNPYnrtafyYX3YxxZkFuY3lEhMI8JBCxcdUQNN3eLIoLQMXSdLzeaN
4e1pGVPEF031HVQkje0p6hR+4oWI3yEXiPW2NhsvpzJs5Uh4uAT/VIskdScLF1ioRNWyPYGyWhfs
ePHONxCKiOrDqZjFpj6OnpEYTVDUxYicSJ+qmploXrj9rDJtDYulNEDOtVE6xT+DuQRCPh/A417Q
LTvshhlTN58JBi1jBurp8iyZeuE2wnO0rkSEW92S3KC1Slx53QZLtUHK0kf9A9QfVEoiL1m+qbY3
7pjjj2CmJwv3L2Jr61uViWKPZNKM1IdnFWNh1Bs5OidXdauziMgePWxlBhhRX49PpJNTsyk0nGDX
Fv7ULCMtfbEHxYBj0VniPwcZ+DdktnOdnOXQFen6SpUXLA2WrI1x1izGX2XVG9eHG91ORVvbBnMJ
mO/ItgWqV1ZXUdPKCCtOhc21s22AvQQgPLeLthCAY6LdRwo++46JsqND42m/t+PhJXCYN6BED7ry
yMZIyiJAPmGQKX+3QI3YyumtnoGJRIL6Xk0RZkcFnqIPZ1PSBCXuMZjygk2uc5Sjt1UfLescdQvl
GH1CItKP96qJr/x/t2qpJNtOwfSP6GoxSSchIgkx9CEax7s2g0XG8olGsaVLYA+w08RXoVMXWstl
eRd1pCz1zOEgT7R0pSn3NsszzfGYQ1Cn/ddEoLC07McxOLaVNE0ugt8AOVW+Nuo35l/dYNV8etaT
0hkROse2cpRYlJgCLfuqeTyt1zHHMnYbp07nG9WBxW0eiPj87LXMSiaNvsLH66sLEl+Not9sWflE
/HkqQi+I7gIC6pXjya1e/hd/MZcmQnvHN3MaKNkwNY2b9EydjJKgfkme2mS749l/N7uixJwtg1yF
5rFClvKRzxxARZngvHp9LBnIcjIPWJYuoQvrGtT2vhfcTh+dqT4znZSOUvrKoUe77VcS9iytgrf0
NxqCbNo40Yc8om3DkfRzVrS6lsrZsok4OXB/dKBkrua8X8SyQ2FpMP1z663IwrfC1dW5Xwor8S9z
ds0wZjuKLeLUWMxgcXHoPeK6/D5mnw8Dt2eaLmizbdO/Y5xO8ORtXPtS9Q9YlV02yyDxuJuf65sG
pITl6wjMbpXzDshr9X9484iNKXJNVD5iTcSv23WyDS3+F6TGpJb25P+pV1bgQmXKlA+N+1Odg+Mm
S70xNu+NR/U9kr9DJNyFbtLfEo/C4Frehg5qrkQQwrw66XzYBmd4fpDbiVjJbZDxj9NOQa64FzN9
zDQOlS06jZAQLxtxKGCFUYuMSrlbMRc5hPWyjfnyQiseNETzIWWpq/KBpH6ayHJBMpYHgbNN0zIm
Vb55nBosf0+uy+xtoi7zMrMv4ba57SBKn3NOHUlyDcibr4AZ3fAWQjn3taW/WLxmhvN7c08DIqWZ
vnGsVQao4AaSnT5dDAI91+H1n9Ov7PY85gARihlAFnIuPZ2CrzHxXlJL4Iwm7J/xUcDKG3C3jTWb
ZgfIaO7gd/5VYSrE3QdTrgE4D2OI5B8O3MCImhgtrqQrx+4KPlcEFwEd1nvJCS2wCTw6JxAQVk6n
hXJiq3MDnSQhZfOlpMNOk4JljmIXkRrR9mq95hgzvCQyG6H1x8PRzA7hp5sk0FdEvW2bmTn2FUDn
+68GwRdzTTdGQVQQp4zkaPgWZJjOrQiJQ4RNlwmmJ+LZz91svb875jlrNIndCYCdP7lcftvgtVKG
5H0kCFPsn8ZUYMIfvNfYmK5ZZusyqGy3ZwIaFHPi5S+qOM1P0Iwt08kw25C1rAGQ+4ESPzhv0cJR
1lQWVDugh0UHmJYJjZSYMuA5yW7DDjoA+rdK78uR+e4kcy193/MP2rbqCr9h2CRkUAeDZsXxiLbZ
/6LTtN9jlGeC0yFtdRaTS0szzKnib4EhphFyRAemVC6mjeCC0CItlDaAT4wROosmO+lbo2g0xNqF
7PxsVXKH2pw3ewGHt8v2Yv1RKuK+rE9osYX0VMSS68BNVBejJbHx/ridHobaqJ+GAb3AMKBtoceK
4KMht2dPb1nR5i0U2kZnnKwBPM5V85JDViY94IbrlsG9pNp03bgpRF1YwN8YzPJ4l3L9fCi317WQ
oeTI+DseCznAGJhoSRHpArjTHCje9ojeS3mlyAvZcmB1LB4BJ2hzCu8mhixpDcaOCUTGnxFo5xmu
YqnVkQNZtOnvQJD40glG2JVXlulrwGe3M86unp2rTOxprmVktQg4xzq58mJgWaRKMS2A4PzFWl9r
gr9WVfi6CX9qVC2filsiCguf2Hb7MlUKs8PPZI/ddIPPQceEbNtUNcN9eLlqb4MfFimJ6b0+Qd8W
JBfRXApPlr1iY1dS6LdUzCGfdV2VxTUJ20KP1unpMwWuTPKPsteBKiEDDXm1zZc5+EWteqFwIr/b
9RHnGxV9f514z27eRAPHe66G1BaPiMyzg46fiEbhDduSY9cuKlEIWc1dLZgYs9RRxvnRPI3gYi5J
qho1M2wjTucW0nJvcCL4jPXVGPWNj0sSmjQ5xYjhPNCB6jyLFdLrYdFALZGm1sHhU04fnMkG1qxX
ruGi2vr5MLBUWdr9U4GtgGHnZp204D6GxeeRd3O+w/eD8bx/g27/JtZjiBE7NQsCwm734J3ENmXn
MyFn20oa3nVjIsCXWbISndhvoaGm1x0ZlQN4tFBjQr1VitZ2EPM4I9LVJcNkuca/Ix/D9JSSZfwa
7owq7X5Q3smiKZa2m3NQeC2HSh15YqLgty++ZeqiH387CZ3urEn82Oi5vkhuvKx5ga1duUVX8G3v
378ZutEtdE17AzKhbUJbr+zSbua3bqlA2XBXwkIZshnh+LqBiUrByzeJO/dOw7OtrhswKoKfc/Fy
hhUXlRBIjJIoedSf4Ozx5lMbth6HSF2XmhN1hzjQVZcYv0cuzH7cbIb1ZyqeIJaVCRrfYG+11lBO
1vIWItgdxdDdiZI2TEur9dkr8vKFoisyCs5QO4BnsA3na/hQTSMi2Snwe0KikRWD/PcmJTnij2pc
t4iImV1WWPV52WA9xTs5NZv+qfjL3uHeU0EZZ+PbbpgBcJGxtewELSFl0vf8bwWcmcFfy5Hc/ab+
xH+FWiV3ND27ZoDThQuWv9SG+enCx9jvuSjArHLMir+vO7D+DfsbUCC7dv23TxPkgqNL9YEU6Wxc
LdwJhCHTh9v0QUiaSvNPNC+GPzJx5cUWLECypuh3ulrJersTn3fG+UMGqBRKlidpu/I72eodbSnK
13SsI0X2G3zMOhtlQlNTQ/W2OaeshJrDOMvNET1Mt6Gbzp8GXx0ZI27jciqxxdukfBcuDGgEiiqE
JYEZR8xtWVQnPDqUhjx9IyIZTwRYMhhCofVqfg9ko91OJN7xZ3g17Uz+9EUZqpgJSVUPalkVa5I5
xhu1j3wvxMM2gtuWeKzO7gwvqLJL0qPC4F7mm1O322l0YwEqjMaC/fie79eUlNmQP+Zgz78WCaj7
5F+OMhG2mu4TSPS8D82bpMLDZjhPCHltwz5z3F6ZrAGDhEkk+gTLL7kLkoEvrP8OTha/GwfF87Ut
TP0/+2cQ7R1BV2gzCc0QjbbM62rzof76wvgUEvWQ/fw3ae4SvluRbCZQLilE/cJ4/Dxifi/viATB
yJF+BFltF4BbRVkiZ+ZJlbjcz/p/WaoVo15c8Grw7xtjBGP3pFNKFNuNjgUV01zz2q4uw/5P5p1+
GPPm/uJalyqa5L/bBmXEzPE59SM0cARqdHwW9svfTN8afQzWrFw2HqsxCAbGh1+99F0CL+3r7G9F
R+2IZEcIqHcfhl3h3xQ3R4SZRA7FSi1H13yuHqY0eju2OPUm7d8VGLctF++S2hv6WeyPfOXUyavY
OS+Zp2G3BjvU2VKv05WsXCfnOH/YV/94CJ4G1yYiO0E7jQ//gSXLuFOQSf7WNJ0gjOeJqgWBXORL
H8WyhxAhKM53TgDqHqhwOX59Rbw+8yof1CLZ7eLwTioSYfHr9u/EqcGg3FdPz76VzrA+etG34FSn
uSHJnAWbhh/gOlzYvUX0Aapftpcqtz1y2PETHg15450qHV3hHUx3dfRvxNjRzNXDVVej8t82oOMA
S2YpZeCJ0Bg9Ue4hu5jcW/giM2sQ+mRmUjmKYkruAkxA6GDgqy0nvSdGBngXlRZ8IIaFh1EK/h71
Y23ldoqEkBJK2clXkVk6FtvQ0cjfj9QAekTDQR7as/ECO+3Z+ZPBdkLrmfQJFB/BBuWgfH5M5wQa
v+50JYXrJY5vwcd2KRAtfbjsjqB7kvKQvqAvfFn6187Fkn+dN2w5QmtRECwRI2p2piHlmiII409S
9lz5ZtT4XXPebQC4CGYmltg2jFn0zJMZBU0lAlEngtFGLQvXA0K7jDlqfTCK7van+M4aOLag+yId
yFNyIIedE/S5NFNxMSPO2rqJeqKXkNW0pL9vPqHFLZ7wnWik+p/zIjHfUeryCur7q0CW6ikQnc3R
v/7gygW2uzLNBTNxIqB6xXDQu0M0N7TPobLJNDeHG/xXgSgQspozBE1MAbffZUa20pxDLZKdvL5v
EqvY2D4Wj5QtEQE1bqWWrOCplJRBI1W+3R506j8WYnQvA+SiQg7qAUy6Km99m/YN1JCJl2QtFnhI
+aw0/2++zw7GbnTPY9dXRNQdWd+WScWE6+MbVh3kPAce5u54AnOGv6uDsRhxprBa6eJdovcPiLvr
IKUx9Cje6YjR3Ym8oY4TgJkeRwAolRo3k0ykUQfGyP1AOv+zQvx41i/ULkG2deMdMfSRP4iDyd2l
o9DjPzMcKuQt5sI6yCeNk2PV5m0jzl2E0d0vnu1BHsRCu85KQQaHQHbdUyBv9pvP7F7MlQoSTo21
S1Hco77iaYZlw8cXIL6r93AMNbJepKfgdVOMrFZWiUloUT1oOUaYMvOxUKgfDg/Bgr9iNMrNb95T
QIla6oLwIPnr4yZxZ7l28QCoA+9/thF+IcoGLH4je0aN6ggtynbSRlo47HK4Vth9HLHH24Oc/VsE
ICiSW05GZic9bN1XmRgR0DHqKFkITds3dZDv3Ekp1L4mCz1RTKfG72ONLTkBAqwROSH+6XgsRf7K
rTNMe3ccCDoB4R5NatVqXXp/zGF9GZGoo0YqL39VpcmyJOyHmTRlokBexYTqRzFw2NVvICDe3iXa
ixTdQBOHOKGkN8fIjfQgX5D+oiso58WRR7t8rUjybn04e79/NdU4qMsBumLpBTsc8tN3GyKIQz5R
SUw/IueV2YLy4wngmfYvuyQ08IQalVD0ys7vhWrFiV9h/v6eDV98MwjLZL9osiiwSA7qALMLdNAr
xTzNFaExbha5jwd8uS8AAWFwxO5NiVQbgqfgbDYwH24t7JXnmWySoTTydqiv2V0C3tz20W5D3DHu
SdaaYSGsnbyFUWirpGYJ26MH8bR2W7eIsg2cAA1khcb8HCv/PHlD3ZzmMIzwPGKIocnyJzBrhLWo
KbJ28gVJSn/4WjrPA1lAsXho+1PIRp+x0H/t+IS8Mwg/Dbxk+6kNei9WcDKxqsTzRge3nJTLLiHB
cO/J7k4lnhvmyELDdNIoWuUvTSTUHsbL79VV+9QiYe9MxCZAiVHHdhi2R4xz7AtZlgGxAB0mJ9Hp
4GAhZsFJV76eqaH/c9erLJfvYE3CC+ZiqfqEzCVW2d6TZCFYuyFkdZ7c3wfenzm8uyvo1LCnCfWA
Ada8ycjWGfRHFp4OFrlvpfUMBKCFmx4OrbSgN6rrUgbOY/olOUUUDAs69GMVEjpGbiOOFuQIz0Nk
EOYtZJhoOsuVrW8T3PVa7HwfE5iYDAv/RcnSdpBOKOugqYR89CEXyKJ+tMk0+yO+nAyVrjgXaBY6
qbmqCsoxmQUTG2Sguh9dnpriagTcgozlMiI9x1JagWRexC9UFs+Lj4I3FMj6dwLWbsGXcgmtsZxl
bjJcQOB1fclcpIGDH3XkivzCGxdgz68cESWCDg7rd00kwB0onArFtly9uVOn26HToTI++CJ1+uFP
kqvwqKzKW6FcqL5CXVFACrluVO10TxKbXGs3eTMx1sU1kZtkHy6c0JQPC3Qcv0XW7ya67Xz3ZQDD
y/q6aIhKosGavif2kzJOloefN6Lo2+Qcy0kR4S5OB0CxE+YkfS8JOtWL8iB2cdEid7Pw9r9W6h6e
Uw/r09g7lKGSlx+hS4QnG9WXOOc9rvlEYYhqnvrcOYQ+pvjobMaaoLiLa1r/mvrYzOzNJSqn7cn0
DMws52NFAWAvl9A0/i5TCmYTliNSM+DvdXmAR6CDyZDPzW396P6WBve78+8QblGI/GKyekRQmAxk
D4eKZyXoZcrGuGWPURoRFX/8wPGbNTNjYkwBAPT3By4NUApts7pMz6shI7wsMvC6zEVK2yrmIhbk
YNYMh3I4fnRvO0OILwu2CHyPSchdBm/TSdaQO7vCKW/KrhdcJ3o1FJpcwrW9Z+S+/yUJ1mrWNRTV
nnQGf2MVv7KNqs/mYOJDmLnr9vWsnh2tZVaIxqmi/RX3CGvarLExY0ug4Hd+misUyaRjAiHCeoDc
3OvXp4WxXoHVjRPW7pqrEgkS8JdxCKa1L4KywCgJTyuaojyoazviRwekelD10VjrPQ3hRjeMDCqz
8F/KINxwnbi5wvgoSFDHKMZJ9X5LdKTBoQVJFW2tDBWv7rSxZsABIgmg90wQJtlW9NmL6MORysvA
IERY0QTn6DrUbEPqBcJqXGfEOyEPx3r0kA/AwL/sezf3L9YnFqxB+olrEBvO31J+awJ4fGKo0pNL
Kqeu+Xzsa7vKG7nzBvZniu+Dx3l8peg3QtSmxKxP1SHlm/j02sLx0O6bAcwBPs4ioPCUSP90lkym
rEe/uBCiKcVcI/NV6bbQUl/esFDWOGlXyzX9lPh2Ko6lPHTGQgQbOlpq//d2KTKaQ2faKhYOhAg9
SVrkEqJ+TxV/X9gq4Tcxo9oyU1SqSQMW0YXhIvAuWUM6pQ2Zsc9wejFU6NxiHmQ9+YsAcUQzQpxW
/fTSOQrHY2+bI0fU+MzOss51t6CY59rCpubBlVSZR8Iai72jlrXWq8aL0lLIo9IImmMkM5ZSdx54
lL9Ngci8HOPdQCeyVuby+dumb9SiQKVVOHZarNiJjW94Pemm3RK8ZUmkIkHtm4qV5B+/OHdXc3f9
Wunzkfl8BPufqPapajn2/Mg5CMOG0NKaVjLgworesOO3igPYRGlVO62P2rvJR4/bXuPiUCxD/FbU
3bpuHxVYNqAo789a2gCjDoGPsH/NMGmz8HviG8FkWxOyryQQWdviikIAU+nqzPVyLmoAlH2KHre9
UubJjbQX//tFmH6ww5KPweMdJ7rCfNyBoLkZt5BjLZCjtwpJq14p43fY65O0WwqRxEjTX3sdhzbj
7OMmkq/jf/qdMOIPu/MTwL0UAewhonOi47vWfH//iZqZx+6807largzBj4Fg+k1yZIuMVpY+v3LZ
Qqzs9dpbAobz9AbeYkHw7fC2MJYn6AsnD2zZbP2K2S8CAjZlRKEChOA2iwb1Z/ojDA0TZA+UIQF4
FJjEZa0wxZhBsHQryzNg7XgTWapP28IQdvG95M2lNo2hiyq5iLyJ2zyN1QSM+3EuKXAuKEHG+jnD
K8hP3cSsBYgEvfUE3zaI/c//bDx4KBwMT2EbjTLLb1wTpOvcTj3DaptAl5ZTwiAQCqvV9JaYoxPc
ustYPacmZsLMa1QIRfJeh8cXEitHfoD4XDY1XHaDZQ1OFuFweeT5I82bT/sjcIAlIH8j/SbFzkE0
aY09mGpwdRTWEAAc+nGy5uxjrB7LsEzL/nf28k/DmtuXUOP/giGBXD29XcE4Ri5YAkl+bqfUyy2P
xO9ZD3m3nsvxyfkPuYFpHizl08nxBxVAyrAuwy0331wAlLctvSM6x/6XJOfKuwSl/1spPQveSNtj
FwM5su0xD/HG3MZ7rDyDW3aWdCiryTW9nIvw2JZPgn3jYK0shOHaxmaWkQdlA/ulhdOI6FHFiyfm
TWD6lyL41AIdbUVlkPbzzc+48NPP55671EPojyiSubepwjt+KLGymLjNLcgFwQ2LoKLE8yoLps1f
PsDcurcCKxPaAOif5vPu1XVrqj+fDib9o2vJb66oWIUqk5IZnaz7tJTHe486Aa7138QkagU0tLg0
E2NYVL73kkHZSQHRFXD5sCoy/91Os08YumsiA6vTR4QGGZNTtClIuR1uCzzWzGHGPNZHJzyD5pom
u2VNeteQS3xWOSifS24s6oW/vP2As8mYXE+7Ih/mimhXJ5223eVo95XWKtPh+RQzp5KKxScnxkcO
TMHM36Nh8YCoFzNRGwdDi7lz102TQ+4mreh72v7qcX6xJDJVbyhYbEzzcCXHz0OQGqL3ZIsK2RMx
WhdzUCrQQTdw5lPXjmIqjCPZGy9wpRypfE74nWGWwUsVLoGFVNQp4AkEGNF3J3yDaG43qiaWuvVz
YjvAA99jT8eu5UZl7zqVi6VQu5YHrY9wAI7PXuhj5RTbOj3dzZYqk0UFOUDhpwVWfSgkCPUVNjso
A3W7YCGTbIgb1AQfZ1WHXDBOd6q07Y/JXw7OWGjhVpgZMsgGLN44729B89hQWXPpmKbmF+wIrIXO
dY2kQwTgs5m/oDhhfIrimStjcfFZa+Kh+FLXjSi/Hu4X+tJq3KDwhnq1e+7EQHiC9SWVoz5iPFpP
+avhfCVrBx6nCL9DrfNAPDN2fH6OhgE/5zIYQ6Rdp6+d5cztpk7iNVW4hWK7vX5BvPZheE9F9zyX
/xyWk2mFaTjUMjUhXTqofBnQPpMzwCEU0nExVXGYmdKhv9x+rQEOMNsTMyzn1uWw0ZTwBbIE1p2y
CW+ItyUbqCpDc/V1AW5lGG5geJOttbx4e03M+lMX9yrK79mAqK5AhPy3q9PAjldvFXlnEx5iXHB6
jAhYQC1bTawkGMNT6AcmIegqlC480tFkkR8jMLfco1Qv/6X8p5uQVXjSNQbtb0EeozC69eFKH9hs
3QiXLNzi6gQS+ORNa3om/he7HNYXGCSvzAu+5KTNdbIfNB6ha4Ikqh8L60Qdj2jSIa1RriO78lAx
eWnAtf7xRGvd17a0dunkfMm0LszeMd3M4ZsvPnMbjHg7+cOF+kqj2l1HqE1E/HeAkJuQs9nl7Y7o
swSJkr24p8QL9LwFyKHjp/Tp1VnjfybzrNTdm+XILbxtYkk4neEQAhVFTQCYQOla1VK0dy7f6eMV
8ULA7hWEfGckZ5IKWqeUHqTjTpj1ZDKRK9GfsGbEecw5YkjA4BtJdvkhkaY9EdjRG8SZkgZ2/g0j
PZFWU/5L9TZ/rlXhSMmIHfmud6jGaMuy07/FgM7TNNirdaxoECdwLrFdfhX7fAmAuXzsfp4EEZb5
N1N2taLegjTRVJoIL4/nyHl5lvr5Gbj1UK9QSwYF1PROBAlEi9MU1r1M0NibBJ6FP/WUxvi6sSMC
ece/zcbm04aPl4UsOejBuJl0E4R20ytUXAZzPDKKV9IChPJZAr+2W9EubVaBsoIIiJHsovOykqd/
FJJT7xDUulXdmYccZ1xVwUPVxGCV7OJQCCZcCRO/Ces44lo2Rmw0mMVfLUEzMZUFR0Vto2x/iiwP
zWShxF+PsevvDszcl8pVblVa6uzeUNsuEl1Ljqfkl6zMmZ/Tvl1136AZmmj0G9AvoiD1sMMlC2cu
I1i+wk3rR9UchFNLu5rMOQ3VDNlVJl5rTXlr2p/0DhnbAE2xAD0QdzEZy+sd0MCF+MWsmGrJ1Xkc
lyrxGpCE1SL0Kc1xF2dNhPpRipzQzzbYrdYC680Sc+U8YKWG1txtDRtxCvGaUayHsLB57v9IZXo2
+2UNpxOPhowq5O0N0WX+u8fuxdLGXgXBPECG9PhhVomS1c7xR9gneSyc8OMKfuxgHzseANHxODiy
5t+Oppk3DPJM2B1fXjSLho1Q9JtWpGqoypiPFzBmPzA/AqexOQo3ypz7TrYWA6OlSTc9gH5wYpZd
oK86aOAHZrHeJix9SM9rgAbGV0I5w+RlvCSzfEhfBy/s4L6YR8UoiTT5dIemmmLueVBI2kGcXj/p
ZX9sBWO48D5jLfUd4DNS+mXsKKbLykCqj4KczUqxbtTRT0fgH+LOhyM/P5NgHTTUundx2H7ysSo+
2JsZVj/shF9zNG19Dh0FiIw76q02hVamDxXo+Mq7Ni5Lknwnnarft5GBAt4hqA7BDZffDrS+WGDx
t3fE9Y7ELcRTAdB2Ttzs78yI8Df1yVSj+T4KF4E8ffE9sBB7MMKBtec03RevabV+dIr43alDFJpx
KQ9h2UPGaIGesrmWo4DpzmRZlSlphtz4jRt+hpY+wTDDEHJ3UhAW1SQfVh69g+o4xervi1daPiXD
EgAn4kFHIJvA0wzXiJsgupWkEr9SI2crnLjHsQ7BXf+RFwo7pgIKKrqQ9fhM0W51eM7tw/k/IBWk
nSs5v6ynTIQRuQefJ2UZbDhniw+RT3DD53ZIZlM/rlDpaxrRcIygPCS4XjGbagzo8I8mKsMynw/s
AzKIz+M/VUFJvMk8OY4hc3SLyUO4BL/o2ajDy9PHR490QYsOWvoHeR8hRDmk5AomCY5toD3Bpxgd
SqwUFya7cLKS7pNPZn7mj39CdW8R4/jz7g3WdX4Lh4HCKItXWrvoMTWoFxTJWrSe5AsROt8GS09p
ZNXsoSEzK6d8cnafvu3Ib40Lyl6USKrTCZBdwh95Tisl2c6Y22I1pO0rWCEW8mdF+YsNM40Ftvd8
yeETF/pnA4Jr8bt3NQK002GkuB1o3qwI97Ohl2BJ/jZ3DmaUgGrEehoCasph2BDOhbWeV+Nxg69r
ujZwDnvdhKzrYV8+4bhqpABhcpisYxm98sL1BkTLcj1aZcK1azElggMBaiIPdnaN2CFDkDaupT64
eVC0rWbTV1TypFX6XjMB2ZndetiXJJdCTMmxz9cvAd3ERj605TtmJNhI2fX1kKLutBY/R5OTFJ9W
F6u4fSCV1QrKe6k2IIKN/F0pABgCXaavleP58fACj2NbMSoQxftrs6U7ruJHMwEozSeMhemiJ50J
/fz1C4RMvbouN065sSXr4HP0+K0rVvliOJzHYh/VwzP3QHUUDYLNzlQ4hq/wGlMosam0olZFsO2e
jf1mNFqJTY1qxIusZuKNyY5B1UlSxSISh4Ef/6/s2VQSAHNew27EJSIqnJdo3czJjYgcB4UX1vTo
CrY1tWPemyYXmzZsMFCyzSHpetHjgKwxIl4Uso4umK0piyvPBB8eN60ahF8NaQVMY/dn8LDVwFHz
qYRyLaoP612z0NQnY46ufPbaR5WlLuLy0zQROVf0BaqIN+qCbfXCo6oKIkqfsLUWtgqT9mHoIl8g
8kwAl+oSW+uMZqfOqncsnMo9kOtOwy6cyDhtyUGJsfd1xZCpHwURmq6h0TblWofaMO8e+sccs7/G
/YZ01RB9acPrSWJ6LgUo2yvZ7SXaGKOs4Hlyoa7qIPdczs2TDv9Ln+NW3xAkFYKXtqW3lIiSYCJn
Pb9dB0zlD+3dwvLcIGBkVawuZ99EP7wj9or2HhR/Qn1kdjurjeAgN+2YCNVjlUjqg4hSOTlpusE5
DfnouVXETXTyRSVK4zPSlNy45fhw0lq2Bd2pW9hPr7slOFMmuC+YYdpeTXu0/GrrceHSgLtGrDdW
bgUZgCyrW1nAEU2GeL4KgS66vPpVKq+16BonvTmh/pj1op4S439NLgfDDkJWVgRZwc6XL6ZbWeGQ
s/2UBzPDR6wxqM7Gk+7F7+welVbP9qBxJUtVcFxJkQ632GOwwFf0g25pnBD2X/I9cPa0fAFRtugY
2rMRfo8Cqjg6gCPg4VfdYVP8Km7G/3MhbACvKTEd6OyDoN3p1swMdUZ/YPmKy/l9W4Kkdv143U4N
Moxkj9yj33I0M07LiF5b376sVsumWid09lGyBwfITe6vQyKVsjTHS2wY9jkdpZpxTSGFft8GqPyn
1frVHI56MK/KJLSpFLIRRXNKuixNTwX5po2GAlVXblHRdAqJPg759PRoEpi8HEgf0lTvQI/IdFRO
UkqCCPELlsOUhEyuxs5lGQdU8ZvNojTQmNK4b2V9d4gSNBdxcF2lm/cB9mOTWyxxiV/VtA6tYq5H
QR3twFDN03JdVY4+UedRgLCJYQCzPNEquby5ymwCu5tjtzA9W2Y3it3o3f6/Vypln4t/IstEKneX
SxZ/1JjJkXNryLgf4jibOuo9xG+x0ECKXhwASn5XanCrFB4Y1D/KDVWMG9Bb1hTC1wmx2tciAM+R
FIcMh1ThVZ0fvX2n6vDr1sKY7AhhbMdjYyAta73u6fItTGSShqg+x8vtqKgaQOBvTLjzlre0z6Se
UjriK42kY0rWuI/MytdydAg8DtwG7D4UnBz1ohqyFIBvTRFaxwGHlfZa6RtPpDCD43QlXcny2RQP
4d5ux+dXbtzXfKYMXvfVZngUYDpAC1Ozwy82v5oLp/wJSEV2RZ7v18AMVlrWwkpUly6TUdJrVq1V
wW2Fe96S2vWxq22kU6mm0Mi21EmIl1R4xc/Fjc14cHJfvyhxpfJ/4jJMCDAkuW0/kRrgZk9rg3Or
608wUpWaRH6V3FzJ6rvCNKDc8eixZHXYMKiumJCN79E06jOxHSz9C2+V1GWBKRMbIs+TFoOBfob9
uJq9RRV4BCpLWe3zekOx6mT9hWGody6Xw+nX2vEIORSS9B+wLswUEt+6kcketZCVAuLfyJtXrk4H
M29uXTFF4tbLaFpqTHKw6Lz8QK1S0D1FkLOV/zKrld2wpalJMFdUlPWDOPyxCeGd27CUXW/jMmdr
KxYDwUZcaxn0ju5glVj5iK3BcqdSF22eskp4VtEM13MuBuUb0XyDRTkpHvADJsIp5mIQHPslWfnQ
MnXul+NBrejjL6OQH1U7lXW4zZpVvWHy0mKiyP04hs62/M42OzRZqyLW2sTyvCSKS01i+4V6U87e
58JZr53HySLGQf41NkfVAcFavJ6tyyWVa9A9oGzPVjrxHPdzswv9wSlBqN42Ks+Gac+qDAdncyh0
ESNJ7B9IMLYGVlTyT/ywbL/uMO1Vho2a7YJj/R8zchFs1wmMoI/hvWwIcM1CFJJhs+TABA+Lhb/O
8sYQJiYmNrs88ZilanTa3mhBA8EOj7gFRwTPHWJfX0tiy4bd8HVfII2FNjaan0AyJLLpght0e+3b
Gk72gFY5BREoyukzVlr6N3VFXGbELoRXX1Bpy7vgma9PSLm0RcQTnzClTZOmL9JLrlE//O5x1FXy
XZhPisdu2QQt/sHEHeFICa/1VvG8LMRNLQbL6THa5+ctIOODiIQBvxJLfcFNaniBenO9AdRoESHo
nM8lGzN1xLhdAmH5dBUMveLvosfXeixiBmMVNaNCgJzR3aKRan09saIgcZwtef2MOus9TcHTtGcV
1gxIRdS1FlebcqaarIhlzuOPZ2EFjwty7CkfCwhFBTW1AaEJLD5xT+8wwiKQygwr3VIrgQJZURDI
zWMQddF/XzIALqaPRCu/QMlyTabcR2EX33sZTYCaVcH1roCdeHzo3k6K+66Qn5r744ertE61U+wJ
o2lp6+nvQxfcN7UZpnwPmk1OTGXeYQD8LqNmLFqoMhJMzEWrp1SC8wlYimKi8PED2VFpqlOLHtYp
2YRUgAw21KULuqHhiq5Kb25Xirl5FOPYVRpT9k7rQA42k25dNRVp93FhfRovxJBt35c/56kMsSMR
4P06WMwH/7f62oXkSxWD2Duu+0L0KuHrMQFqO7+G7IxUSBdrKh11fedjSv7/c8CibL08VwbT/WQ8
L+A2x43MQoD4R1bAabNHhbClSYB64O5JlGk4cR3TpQzXg3/wUsfWip8eECZFLoVMG/jUpPEfwh8c
+MO+64uVADhP56FK0A3ZCNMK8WhWodFfcVUASOJO1XFXqKkqEEOM5GuZRAWaMsDGR50oNdRhMm1V
ApC1DD6OheU9MIDmgo0NmD/uTn5h0FxlSY4vUoS08d6ibIsdzDp7p7CTxe7RAK1Mkics2kubtI2/
BVTKbfaJJWfPlIE9uCjFHAsnQLRt5dNBatF+lCfYjkK0e8cTSr1sUEAu+GFHF14YWP3Hz0uYtcCM
0DAiAyy7Pk/PNkQm2suKcpaiYAWb+vrY/plEPzR15pKfmDjPqRl2rKCnwS2hUfLxa17UTGXejW4N
Bp6M6ljUdNRu9kG8FT4xIyy4UvyoKXOaqEzP/QTk4HB2A90m9HtUZjuJwhKV3VAKEdLvJcFBOFi5
BsJUDgiwMCC8QbpRzo3UMOOl04ZE4g6J23e6uD4z315UGIDuM7gxkyeCAcetrwWMc3rElOniMb8H
5LL0Ex8xx8Ylq6gykahKI0nLDhcCLFzlPKJ21aoaajn0ItcJp5hBoOc6ZkfB/uCY6NPW7DWtWhQN
Sp/iXrkE9oU6YXYAEFQwWcZoAOiTLw2uOyRmQZwN2MCwnAq5lnDt/to+sMEb4ZnwY1cdiaGAKYdM
ot4YuMVvjyzT6ivFeVZ6UnxrWGBiGPuvTuXL5HmFFFgwEdiHGdszTaUA0INZRaLGPKHV7JZ0l9mV
VBLuYV2MujFFHxXC02baVOzDmwaGhrkAZVoEh72BOtiqsBnz5Bj2ANpLk+yYWFXiFm3/FQhv32dD
0/c8G6VtPtK9piIcBxyh+wczsbK8Lw2IUcltN9h1Wt5SjNlTGW690nbX6WDZ5bLFgt5uRu8Gzg4b
qoA3MgQzN/r2mDGRXrIGnGHYmk9kQYEiLZ6YNvbcu0T86e0yOdlzUMkJ4wYBBDu8QEkQvVzvORwW
qcARJTNV6tfJAtaTTUVy93kgQx8rBxyIG6BbZ0YYUd1rnNWtgGfO4cCxLtJTZ/a+2kNd5uv8ch9c
QG4H9ZH42ZS6u/wi44ghdSmI0IXyIu1CM6Ulv//fD2nrXp3t3mZ3g4ri1D2eblq3V5hOG3MZWPWD
JMAgTl1vj6VMh+0HCLRZXZi/gbSpTCTxIYxAu2o24Ecgfsu8eZu2V7pVYeZjbA3S/4PZLucMWkQS
igv9Iq1YN/l/9a9ieFW6jOQI7IQ7NC5Kh1C0zF2fIS3+FPf0O01fyV2SoCGiXhCJ8wZez+3+v1aY
ge0PHXY0bkSyW/Ay2rbFHEMZJrElZnkE5G7tRZWF03IrP+8oRiz69ez09tyIXCOn5KOmo5f46EO0
tDogTvTc3TXIzoX9Cj1pqMRlkYjhv90wI9hd/fBxTQ7eNf6sVFJfXnQLiNakmDLxCBsrbGrnIYRe
guUd+GjtPwBWq6o+ST0RFKZ3OTpbCLMc4pnTj1n2iZw5jfqCbv3WpA8ch/EmYeHmyuZjBN/otog7
ny/Z/vUsQbTINO2hp3YJJQUmm1qqOiV9T+LGsG91YfeWkxp0gooCX5T4B/pqTZO0W+sEGJl+OeKo
fgocDU+r1kT6sNK0rmL6yjkcAa4F8Tc2CEXsDidGoEq3rH5bKf4yEatABt8QHs8n27schc90dLHy
s4V3EgqiA4AU2bfUC2xXgQETlXH5/qrJvRfFVN6uYylIyymH1QaXcen4rblQ9oXa1Cu/+Pflgrq7
tm+UaYsMAqhPmBWlKoc/o7pD+URfrZ/kC85CpFKisg/xy4ZhCCHEX/FvvGUXB+iCBCNrXO7gFjBM
QRm6Jrt8NonFtdS+7x/nNREHJT/qQC0VwSrOODszoF4uXALyOFcpq//9CW6APTopYREmUneLXH+G
gOckLUdNIG45vjyXq1Hp2NgTB2WG1YGBe9autnQ1z3a3dWSy6ipfJbnfkP777Xq0THqUwospmDLX
IydhnhYjWj8Ga+jxy6pwbaurxQFVqQ4yDmR/bKjjfHl+TxB2i7f6eQizqO6q3BXI3TtJlODxZpF7
tOQb57wH3LizTQVbCW9iqL0PAwwyETqLMUmPUpXY256BMXzrwUr0E7dA2wZpmZo4r7ZY8aoeumvd
38pEUpa0fcPW998+qdY92UkAFecDWyrJvZiibdT3GrFmP2IniKsXoU5F64+zVcWsI70/6ke9Hzi/
W3VZVDR/o+2EOjZxwHqUhgWyVkRoh5fSVneMcHYV+QVXtqhNARueHQF3qvyh9U+vwchzYrvCBlYS
tHZZ5+Y3wiummk8naxFrenGcWGpyGKxDCYPKvapAHHGUMKvkiipBmSfbd/iZSFheC4OKgX/d4Mbp
2/bQkoNm08E28/3rcEDg4Da/K9eN9rcENklxUe3SX2MD8wIQonkI1O8RLQlcaIXHAynjl7VlGW1+
cBOXPsJgtkn7EuUC65+5Rzv9I6W+h7oTQ7tJdR0XyRK4aX+NPyaZ2/+ze4+ooG5Nm5AErWm1JDHp
cV5tMveu+V/ketdusUxidhCzr7x69GitLS1Zd+OCpaiEhNoLUGQhSgiMUecQU8F7dlQcMH6FmcFt
hge0kLcJO+MFAYvV2HZPBuHpGNdBaG095TdtC4yjWvegPBGNNO52pmePnWY3bkMoX9/Dbm951QoF
huHRslVTRatn1CJPKVYZcPizdg9y8Y5fR+t9XPzIcbeaEQ0PvfCvxR5WSE0M+PwutAHElUywqCn9
R4xlpSMIGfFkkrRE+bkLv/sGV9M8ksKjNNQ6zzUTaMpu6/0LXpqWUJnmK3nql4KNqcvwCoIFnocy
Q/fu6jcOj9A4XZ6gV3qvaZvdlI7SCG+dGYKTwX3K+AW3z+dVKNi6c3qL9MUdUAAEyrLDnUAmRCpE
lcrLGtEh5AZXEJvtsEwhKzXQZRQdWGMBsIXKGnY+QIKI9Fml74zYd9p4bc+EAQQCN2ktEKodBguQ
/EGp9haZ4+hqjr8xa46AfAwnKK7ms113SEnyFTs3SLYvyGvvwMzjfhaNjrdavF0knceI+tImEfEd
hbrhB8OUltKJ54cDgiGLsCNRVSUVp/IX+jONUuOK0/BHKZbTpSNI2HQwXWHnnLPoCusjIeF9naIb
tVtI/I710JCQHFKRAblJrH6YRtP+ViERb6C0IObQdl15mOR2PTB0DpYlaY9II5V1Db5P3bOMmPJz
Cvg4Qi29swyPUXdRhNXwzTTpxBMWr1pIpA6OqsSL0tA0f9lqVRDd1J1SJL39jBHggwqRXyeWH8ew
oRHA2BI/I5w0bAi3Zxfm/vxMG2BDjp6dHHk0PLl3vFbTVkbc+BaGOO9u2cNamtuv7xWtone8wDoo
5imitbrcoDoJMTIXwhEAFk7GaxxufyuxyGAu4nonfqWQfItW2LRBfyYw6ZF+hrBeJQGDzmRlTqB5
7RAiB61wa87OHFsuJ2KOHeATKwlSdQwl4tUYN+aRrd25l97oieGqO8hSOSG6iXlkxj1IbjZr+lgw
MvHeo+coEDzEjGGWwNthBtHDpqm76z1lzuRIcoxQlzo16wF/2STmo81RHE0ecY+m6jsneI7FlBg+
VkwGTz056yrlC8Bwpl06qdfUIgA4kOPTg5J5O6+p9CsovvKx2mM3EwG2b6PPGkZGd7u9VBS64KXs
PDkPRnAPkmcbHj/YMkkMowhVG+77x85O8Gor1b3MDLGB4mvggrqaSguJea4RuR/HA2F5tQrSBs0k
Y34KPMHX5liaLJGpUD2U2Od8x/C7Jh8P5Dawt7l9MONhmaTFKtMEMqCT1M2tpUJN90a78FW77KYM
ZTI3UJo6HL9udJA7xa+/T07wcwCum38Y4TOJ+QGfe2xGYZR3TXid7S+B9aaj+90cT23QS2ziCMde
eBKYHohZ/Iou3sz10x8LKk9yKmKNQbrvayv/GB3QYFf5PCTQHHASHFgm10dDYR/LCEyKbdekTzdt
WfJY6bY9bpkPNYfV2W6QSpLoFHLT03vMCYzEAWNcaQiP1PrBMyFdFPq85J2O46sbnZf2IaqjmOq0
P55wQ+rIuKlVrlqfk9JGf/vNOBS5pLNNMR7vKBFjli68NA8DV5y1VO3zj661CN7uOuzbC1eV1G2I
5Spfb2iWpIG183bq/mGRLzPdgSWpjWh/7LUsqg55y+2LRy0Gdp7U2OVSDvcYP+/APhQrE41qTXC4
sEghaFgmBIyDWg9rsOsYLWsWXqzQ2vI8aih8yc94LeEHeYBDzlfBlKUC0UuuEbljKjEgRta4rDwS
wZ962tcRJL9LwQ3OvLmPK+lnlVYB70A8MlqcpRLSEOUvVJEhWmmqdNM+iHPg+po6I2KHInpwmhUw
08i8R89xkkkQ8xJlyLvI4RN706PtlWW6inVtQeCknHouVMODFka3KVp0pEFohzG0XVckg3XAatDm
bokHfJ8aelBJqat8r/2+EAd15DB2UkJmhw+acGq2seeRNS7g+fcfl4s55k2wUsgaE5dX3zxC6H5H
tq2e7ehC/wZZLdtBrt8gbgULJdzS+i7gw6mtQunPme69ZBi8+8eRiQNoKlemBrMnggV56luM7ey6
NENmVV8DXJRw9LHVFq1ZojB/2zd296DcFcRO/phWyj2y8ULyxRVERgn7Ab1nLl8OED7xTovhrz1Y
VxHsnLGYBsksDh8T8XV9OZ8tT4vsFECLsIXg5s/z253QGxi7PaVN46vbaGRZyqPdn6BazeoDtdep
05lDNU7d+Y4lbD9r4BiRWvpmYETcF6vbseaZcT4n8CXKFiVI9C9gE9ivmSN09LKURFUxBGTgJsM/
Dz+twmjHFiWNCqL968qv3TyXxl9drxN+O+1cdtcvXpQlxTAcwlsACLfB/n2Q/s3GqaZXX5k9t2gp
BLwV9p7v/QeFxTsb16b4Sbydh93rwzYNkVbk12JiqgNqnda9xAyR3ZybKmBzBcFRP4FHWCR8u9qQ
fKrzrg5IVcLfPV9LiPgEJBlZSTL84GKAhEbZbLqmMemcB3TeCDBbQC1TbC26vwwDcBIWd3vH4aRV
/Z9dxzKoZRRLeDYq6GqlLBhshb/XPMOMj5jiaoNhz1hp7plvReri/SZF7E9il4crv1NGYFyQdb97
pKntxi5igLY3SnEWpxMxDXQuOXp9c7vi+I4vmNoM9VLsymYd3Yt+2ZBW4cRMRQVDxm/V/7fv2lYl
ZPJc2lifkAG/m2ntK+SsalucokNBd5U6mIiiK78vNzqnn1deoh4KcliiWzGBf3MaHxLKD6Kqmgo1
zxxWOYJGJl2oASp9W8TR1DcmQcdz3y3rOb2agV+DH3HY6chnaERdc6vF4H4VkPgxtNF3t+ZBNa+d
Myoi017Rizk0nkS7qgfghDOEgfl8Y3ATURRZdN2ZDeXHwEhMv6MOf6rScT1zbN2MSq1RGe2ryME6
8ssi/zoaOADfFh9S7vOzCHf29EikVvUNyH7YpSr8/mXrnhFimgTOgxofWqe8O/kXPfQ67fznDXAi
Dm3eGXIPwfsGiYcQrLybJVZpTJySA1rCzv/JiV1hgY7EobRzg3pFi+syZ02XKN5MiikEgJg+y3/1
h24MmD0i/BZPvbssqfRumJsAu+Jkt0Jknyz5keVo0jGVT7f8jVehsyW5ug7wp/h6lCEpgHBoPEx2
MztwZw/oABqxHI4tdYI55RvSWw/NOqqebtdE1rSf6zJZLI6tPiB+llAmPXSUYot3ZtZH6jsHvrsx
blYCZDlbtbMwKUJozcaDsfnNmU4TaTnB6QpY7lM+HZvBjRpuAqYw80+wIoe1N0AXH9yFnZVtYNPe
z4W3eX7VUNSzPAhrLPvntJ/SJi31m+/xcUZDs7ONzXflj/GUUuSY0Yn9CKOtCv+Eu/V4YcLMvAFv
gJwUcEZWLkKhTAUcHOhMCEev80oOuHbupgCu7VA3Lp3vkiZ6Eoor8TyXs5Yg4lAkHCO3YM6ziqI3
dG5F7Z49dm2xo4+B01wO47U4M8zIHIvduSZNrkVw5JRRsDgnUa+luuuoI9LNcg9vaFhHOUGBDEAW
e5I3i3VgiEAyjUNfLnlosRI/K6+ZAwzFNZP7pRF7YT2OTl/1zW9L1Ua4odAlrr3uhgysGzOO72uh
Bk4iuhNAvcUsdEel8zM8Ozv7lbyq+gGcU+0Shk3RLCOacZebjQRyY5ksBdsHdUGvIqqQLpAAUoPj
ilTzX5QBPSUQdV7tutN9hNsQo98a2DKer26Z86UFAZUMZXct7HMhfIQpZOKub+8ASlak4cTxZDXe
VlxpYAp6GWIPQtmZtF8ckcrHPjGLTmxfbswmzYx0McV124PKcEJ5OSEOcsvK2Jud3F0P9kyUsNf5
AhIYqyQabx84VUfRsR+2bxvpWinYCoedG08/uqdNLqeNngCYMH8dRZ4tJEoL3zB+i+EGVSRsVgpd
fx257SHhGmB0h4xHgOUBx8WoubcvbFXnxkg/7d1ec2FzGLmBRlKqlgqg+qAbpHe7JEdX5e2w/nWB
Va5nqlsBGpgowxumfIp7oykaG+lO+T03G8jpdbtQq3J6wes7gEAESdKRsuON8gnSfgjU9KXiCAzs
217rIf9RL39g+ZOmUs6LLohY/rx484eFdq0r7t+CX36gq3+A27cp2Wq5MxP7hRIZ188RM5mr6YYk
mJOntz8G6oOpcdaafeQMuMtqiwbbgZRdk9vaiXlWryQTQLwQD4JVUBClHo7DWvweT5Yuv9FjgfZY
dttQCsTlMa92/pGZyH4OFDel9YzVovvK4gEGe/R9s9utD8Ltg/EDJw2h5xfkFx8xt7+8ILG1WgCT
umkK8MOHD8MjajIjDykTroMkcJIxjXMo8kbBr/11mNpwQ28e0OeRo5WX+R7+CoY/7g/SZgBOBMCe
bOX62UIc8eqZUySPukX7nmUTwXImvadvxQ5RuoaszRSVJMob/gypb2vYe/spD1pWDY8sIP7mJXHO
WXHSLu40AxiQkw0enyTiUkS/bN0Jwrh83nZm6T0vGxXpthjwLCETjixl9a9J7x/KHlMFF9GUhxCA
xEoX8EVROBebkDSDhnYjFPjWZU51aVbhfT5C3HUOiWcxLm65ZE/LPg0LGJynse4dh77+9IkogbsX
I8qmAcVQLyRdEblf2SQJCPT9gnp9o/rJzmu56C0JB1th2z9Sr0SWiy7ooCj1PpQnX0CYY2dE/enr
bRFQ7Od9XxFEC1qJ6r0cZFcZnvqAbg/klpIeIx1OzlubD5EaOCzdHEpS1dgLP026V1FuLeukWFSg
gKGb1egpoQ38Atynh+fNkLUCsdowcZjTEdchel9UOrBKNl+fdcyvAXHV39SsmKvMCvhh2WmtdTCx
UGwpD59o4dHZzguod+BMz7oE/od1WCrFWUDsq521YoQVxC7ZiYVGRDT+GcQG63204g0GlSL4f/1H
b7v0XTr1FTok6XO8fi7AcTMpNu5ZnE/Dd+5VnPg+ND8Ktb3ZOR5VgX4EJdE5ITrtb24RG69oF/dN
ihIOE1HlNcztm4xMBc3vi9dAZxyCvIM2/5T146XB/miGb4rKnzNczMRrWxa8GLQdqASLVH2T+tKx
BW+cimY+jBQhRv6xFEl7qSoV3hngsltzgyJKHON2e6ngg38n6X4vDGxODfS/wXYY4egt5gcIbp6n
JLKXbEYpvTq6xWWIYkxdWaBVGiAXAjGj6zrYpHmQYhsF87c9x3XMbq1A33OhsRsWIKpLS8PEB3PM
ONeSNQh5J9P2XboAeBLC3/9U/L2D2kyZMrF5t0GZYaM8UV3vxqi1HRacmQN9HsnocoVUQR72n+ub
ycd/4P5qt8NPmXZF57/HsyIzLvn7ad+rqRbqzlq9tQpXOVhvXh9DqFrVS1mxXv5VRi5d9enERb/D
x2UXuYOBq3NZ7jGhLXvoq7R5cgx77DZLlZONohRtksbmaLeR0t1d/PNqLZm4uBGDwG76wCXnQUPB
iLtIatQL0ydm8cFVk1dTKZmA9V+g+FLneYAdxMINa/B6oRaPe+SjAfQxTzxsDTVrYj92LjG7QUam
oISBc1uGS7w6ep72bqs1fE+RjWdNIqQZqSbCG9R3Un1WhDFwS2V5f21OXK6CGVSD0MilFJzRUK6m
OScpeyW2rI3KLBLPd9B/oHIKB8JzrFnivO0e8d9s7bMPXL8iMnAi2JqF7rTz5Aeq1xcnRJ3NckNj
luDG84TaB5ZvzBLFZMQSbyWi35kLO5tA9Ghokb+JQ2qdr4w5Klkhk+R55CivKwuiQITGL7PjGXqP
kfFYN94xFlpfE352VKZOZYJ3DYvbMH7lgKhaHGgBoRvFuIthUxgt8VCD9FJWZ6tmF2DDB0MaANOD
pvHn2UlYg3SnqNZjsTYfKxblJ9FuYJ59klMOO+kKlzxyC/U0hFOh5U1wcbYpNbTBiUQIfjFvwgrl
8pZKnTRXedhv8ydbOdKjxObgDbk09uWh+f0H7ZkahEdioMwXOAkLnAXVMrb7c8hd5O8V5nA+0syZ
dbqLST5iEQQv7erUQZBHTJd7YenjOR0fTMC4dWliSLbBbPxGVPcTRm74DqBA0w/+gjHv3TmKLsea
uBhuuT9N4Nhn39P6wdFrNH+FBEDIWP+cZao7vLO03DLRgqjChF14lefag0Mm1cEsHXDQbX7h3z8f
RG+N0aiK1nIgT02XzI8pb/EYHm+WlDVWOeOO3YoNe0jOGTwEY5mPq9XmOv0enYFH564sSy7xPLnU
gL6nuGs1EuB966tcTDXNDX4jQ5iQZyjvWDV+P22P6PShMcN9gddEh3wQmEf+gFtj/ANnW0A12fQw
d+Yum/f1+XuDfxFagdaW2dK+HRZP9Covgtkmhyv1PjGAOR9XRJI+BLKUY031mc9Aya5ILng+GejX
Aw6wl1GosoYD/PNMOq6dCmVZAoqun6OspqJPM6ewCDLHanBQun6QeasLtyk+9HnEAyj4CvknK4z/
faef5sIbmQTXI36mGabjOzYS2P9HSHmcTBLB+6AdS3e4UZglRgbCtcqiWUjpcB+HNTk359o3PpcD
o2xwob8BENemXLuS4EOXgYfTqwSvoFxZ3Fo9d0KQjraky2sHCThKadGscBQzeLHN3NZ98h1GI3s8
pAL/3gf4ccKfsG/EMRrLYThhq7b+qW1NWb2Se9ZqotrlyRauDaqwOw6OLtM8WooUUhjWjieMrhuP
qp76xlEhC1CBMLPBB0Y8XfD+7jsm0sq4e0HfrpZnL89BqoRTshvHEdvnKRa3e8jMNE1wi2rZgzTG
A8c5k19/tiRDTeTc+UvBmv4RsAxTxKQ/Z45P2Auf4s35I2F8rfdLwHJjDSJwBOndSru+5o7cSfhc
yyfX7OqJC48xAm51x1l9zGbFveXJKxql6CyuT2JQlVK6iRvZeShTbmszGyQQjLH5t0DSmwJksLEX
zaypjFViH/a0juYj/YtsuGjFMmxYOOWd3oaAJIVd0D0V6RQyIy54DSlWEIris5Wn/p7UILpXi6B1
0sbuq+Ua2GaZPesl79uzc3XyK8/OD2E8jf3enefPHbQwebuql0LgVuUEFIjxhvRD7nWbzaSx7tJW
n/zleNiQ6FkrWbdjKzuMu0Bm67KuDfdH6oLrlgc+H8RzQ6mOGONz8zgHgc+vc0Kvjjx9IgKJNMir
8b/sxUpRErlgA31ct2MI+Ew9sy+TL4ocWYrCLKF75m2Ab1pnG2YAYkiJzwtG3Wojd+Fsukes2zz3
C2ewxolB7TPtmriB9OCMM9aj5ZFvN6xsW2612fasWL03aTl955qlJUfRQ+BX4/dyPaIkuBlJR78g
k9tp2OKv6nr7UYd+Yng1PqFr3YKgJrB3kP5vMUjgAbSj9pf4RZuMZeWrdSwPP+LDzUwPgo1LOmZc
Q/OP3CffIeoF8cxn9UtIclphsxm7N82BFgeg05BZQYhf46Cfy2bDG2cvnqVy1PR9okN58SMIyWGT
HsSRFSFksDMuBRgbNvqZ3rdQAkRYSXQ+2SN0oorYML29DrwOwPJOjBSWX9Q00Yb82iNJuRD2YiTA
KZdCIjwJMvC34G6cOMjIW9o3lPka10Ha2ogyS0MgYRhoAyIygXTBSxmF43qOrz0lX8wITww6iO06
6rtGQgb5S1uCys1SRpgreOCpW1jOX3Y37Ne3+XB9UNo3V5ypNRpnQxJpEAFEB0ZResytpMRGNt9m
7B0BTl1C0MrsfATBnZ0xiBfv27GttqxUmVheHBiOwQKJEagh3u5VZYaH/NW1hPcXq4/Xf+2onR8Z
GLkqfbAegKbTDvrjviNGzlVgQD2a3lecom46DNtMA0Pqbn0ZUNuvMUVMW5CMabTQL30qFs9cnDbB
zAlcYAANWjw9iDcLi8/rrLaIczHbS7e2/Lj2Q7YsVz3+zIcZPmXzR43S3aKab3/bo1LDTPj0orfL
MM0aB8AotUe3XefGwHDK/v9yfEcTp9kHmJa+oCrH0ovj4hXrgmnGcBeKYwXfhq/uhQguzlny7Zzk
uDzvNWpn1N4V6Cis/LQERec0GepnB0tcMRQtQiTCfzAKNaiITEuYFEdBpoWFGb7QoDicU25pEZb7
0IzsDcRgRSmk/UP7xU8psn/n4kGf2zlf6je9SiVx8TC7iOk8jEcBkzUVo+ao304Csbe85shQeKl6
5mlRDDxTuxScm12w80eTeMW+NWo3bh5klCxa1VcQyCxE/3Leqo2kWQxW8AHiCCMptbIPELGd5aVX
h5o8nJDNpSwxrkxFjY1irB2DEmYUSe5mAWvqtWGZeGD7zX9bG16Ji1KsrMjzAV/6PaY+mGBo1HZs
rgrScx6C86MM4h17hoULmiW/yoa+uzldNLrou5mIZZkliMNEMNbLiiu9vFSVnzh/SXrewpsn82WN
H4RXGhspClct8Jwm25pBaD1qNbwaM6sa9KFwmS5OXnkN3Nh111Ihbs76oSqtq1aMpWbnv7U7Wb9q
qRf7s+0yzEd/zj8tTLwMDSdHRf+7LYeXtnpziEoF+mdT3TF18qFODt0chnd3Svu1kxl8tcwDacMw
s+vBTdpeV1829ltDxZtNcDBx9U50qlxElHa9HVap8j2n+6ZRoKrOr3Nf4yhw1Jr4GutT841zt0IY
joofYTYPEcuGQAhyLOsqMTN/3uRJHMwgGr4zc9v9a40c0Yo22Imc++C8e5W8HvMyVezd4/TbPAtb
BQ+NROvE+eBPjl8ya6YqWsiQZhkyjIyGRoxDL2NphauwKdUlLcNE+DAYfBDo+zVpiooTeE7Em2JZ
wEah88vZ1j7wtAdX3RJ5IPcEozWhewe7/AsoZ7VUA5yveeta89haVbblKw1MpxoZrCRghQ7SEOm2
njhkXrix2nV2K3hh03hBLLKnoX1JUaL9cL8RvwAgNz2ojYKdJ/G0fjTEShakr2lPx6SgC4wuChtw
i5H1CYj+fAm9FyziodqN5Qfxa3DFYD3+pdxFOBJYqID4pnBf8W1z8bixHYh81XMJZNn1s36ssWeP
ADKF9qht/SMA3kuNzjztQeE/FhkfTffDiRr24tOyABqIuT5kkuZcYb6jCe7t6nSNVV7oAYO80jDl
845Jvw/Z3dZV4d05XZvyETtp6MoVclFpazIz79JOOzYuJfCOy1Fzb8iMTLlXdIn/kZt0oibFnNnj
eBwlKRXqtcsUvoDx3hE5ApIhxYrq5L911FRS/mW6kgrZucw/6zkgaHGNpZIqamCr6uYVDDmsIVrd
LdNqjMOACTyVcryahT3ixA9mg6063o7TZLJlRJpYvn4tmLs7iPB6zz5v1K0ICodwvKifGo6UcR6+
5JY9uJbU7I2ImREriIgfxByeFxqFkm4LndOJslFOWhsi9tAKBJIhZxIH49PoahyWlVZ5yjjKMl77
qGK3bbB5pilCz8FljF1szJzES3J08YO7YZLSgVIc/ifJcYzdS9Jqa1gcFF7slD9XFdanTpkHKtMR
5TIfwxi/iF/k+kmDffsum9WPMP6FXn8vZryPkcswe2GQq9jUJUy0iy3VZSyz6yWJm7qXt0dT3kPD
xEYb7WNRUGryAvmyhan3L2Can4YMnXdQJ1awDNXgsiKDr9ekBq8vtZLmPlGt2fEvyz3aoJ++vufV
rEejUWGRwpn8RlhqEVTayLt/Zt2q1ubAU+bueBLi4OldD46te+nJZ1sgnIVkG4XFoAYLsC7qwTJN
Fpu1Bn7uEiOJauUBGZJSHM3iOO/FXy/Z742wwyoZB5CpnbnPFfTDlGkD/1tpKwfnlhP0UXmEUmaz
p8QyOow4YlEaARWgsNyVf30tzpRAaQnwU5T6NONTPNSl1n7khkKcSsnamvz0gvS6L8BPcwVmm80Z
RU++3CpPgbXtQ3lLiM4HYCaHARxD8d/E89HMM/yRMI4D3lIaC7KhG5dr6iHH3Rs61SdsnHcr/7mU
Be6sPTo38lYjfDk0CaeIqr0YCXj3/LiXDSHSSXRA+VSNwhgr6vhgTXbKtzyd6DGV4CgSANsvlyRM
eZyJSxN3G+x6DfSvgA64cb7ihzeTRkR11uP8S/91swmBF9RVtcUbLzMri3R4HgEJbCB5ga+bCf0P
TuANjqJ8AzulJU6qsGY9cAuiyMW4pDNPXgKFHlfTan9ddcEHH7gj3ixrV6q+ris8+aeLb6da3DS8
SKtupeyYZ5DlyddzPHbcwsSoazRp00EJuaStoTYm4293cE5F8IGTAjMjopzqBO0XkU6771Kn3y82
GyrN7Zf8fGEhgfxn2vP5w9WifZh1utB9m5Hj90LcdrF9POZVFLxVownWQ1D8HqGoQNk0Zs9z8vL+
+3CbG4DiPYqzEbMVE+lU1uwW5wlMgIV/Pmw1saHQ0gJ6hoYVU4jRJ8rZTojnGu00sFKMF79SDVKi
B+hX6MF5PxRQGGLyV78KyBF3dnjOVSdYi5RlXZ8g1uWWMzcBrekKUx66ug2/fsWvU8dbtMWYh48U
W4ljfMTwd5ftZzotNGW3GC4BLpwQjncBllAiHJbTBkOPUBnC39vEmTncuQyuIH9h/47vAXvzLUL/
u1LTHZV6nYVg17rSbZ2dlR1rcyTfSRLiYJZz6ulthPnuhbJFy//MNHd9o20ELCCg8XGAnBB29imC
aaf5DKEDxIq+KwBDuK2xWLUIEt1Dpyfv6mCPP0LUdgcEbDMvammyxuuh1eb1a/4kllGlOa81cixj
C/rwFGFltrrcFCNyOJrTRm9lEdkek6WssbnpU2hDcUq89+fdkjdUD3pUXCbnawLC91yfCHYmauuA
LbACZtU4UrOwmPqfyT+VMa8aS63KVKi3l0SKj/RzVc0B0oLOJxlb5R9YhVabAEC3+AD5IScrgWeq
uUlggUKgKvF7d8kGifF5t0YsvJvzGT1F9stjRV/e4FwU8ENKC6fe1EVjnxRnGiDwY81dMYTHYOav
87jSg07DU3N4W0Pv6POYjKdXThbYrtZCNUhP30qeisR+e+cYbFQlagYWb6vD7oExQFDRlPa9t3IX
7BUJ+28hTAdkE5KM46o9EDFaFx0n7zaakAE7hkoUUzRCEoua78eC+KfeHBxCTdwJMO4rZddS1zIP
T1Ue69ffFCMu5tyLdiaW8QKKT89ODslu+6gSAODfFM7BxI2rXZIyUXbRxZQld+DP4Cu9oGZ6PNp0
PEMr0LBa7lW96GmsE/OxJSldSYj3Q9Z4i69qIfiG2WI3/Csetgrzbhok+PoE1yNpEy8SZqHL2hf6
Whf+t0X+2hfR1CE11iTZ+yFvvRVlyqIbrz2aqN8HUwAzvh8Hksvk2NL6vnN/wf0QlNivLBiUZhXf
uxA+rFGMmTNZqb421ci4QzrCqFWoxlaKf+lKJiGK2g7Th67+/cU2Ew1EpzdLA1nPT9SO5KQTyB42
2oyMHZHatM/6Tacwb0XvOGCVsE8dx1qF1FkzTifcqz61HxIQJzgo9DjdQaaEApGLyZPYsLJ++YcJ
TcPOfOfWr3co/tSI9ZqgGTWS2kPfj/ciZEPKMRSNE5V9NWc3SrZ55Cu+Gq8tREConM06zRcl5cU9
Q+IOD1NzyVUgpmHn9mZ6tH7v+qnvTXlAL0pJBH+1t+slsB0Pog1JL5Zb8j3lwIwHPvsQV+jHGZYL
kKOzo1qE7ADNvcoXChaiCFEFSlkg9E9IOgNpPQ/JC2VEsXsRjyWY1qstXPG7zohq/75OFISJY02+
Fja/2exlYUhotQ7Mvr522y4yRVmLSWHkYRi1GMvqsvL2Rj96XB3KvYoeCgl4fv4NlfCqll3rQWXF
Z6giAtJ1sWNlUqL6jE7ViVhul49dsqk0nhAvHBfY9Nk2j7eC7TZl5ULfPrIB1FtZOrDWaCvA7tvm
nu9n1690I8U/zyHz31W11nSRh1k6SwFupA5+NcvntjaCd2FrYMIukxSk/kZJD6GfgCIor96/NFpb
dCLXVx6Ke1JWbn/+vwfNiBm9dtcMLkiI8jzKimbY5nUsZZdTTCWJ+XPgXockZ/V+RUSKcYRoueLS
fRYt8kkWeKHbTPiP0tSADbVp3oRSDID9hhD3ZigweV8rjKeCf2yAJqkio05e0+XK/Ew7NNf7hDQj
M4NZXeOlqrhF8YjTfV54xSCjsmIPZuxH/HAUTJ101TOqu3gVEgcHKIamzvd940yWNegECwTSfJdA
AzL650pD9LtGt8BY7uW5xibn+fuqu90nl4bF981SWkZe9Z8knzGMxZXlf0XdJWP/vqxNc+m7VT5W
Tc36qQKyTGzjxzYt6PgW+OQz7wdNqt+uoQtdlkkGFtGVriePLuQ5pJUOdne81hla2sFfwMYS0LcJ
+dO93Xh10+0t8qESDjDBNoV3AslnoBvPXKd7WrVkRfjRLHzfv8CEmYvnktp+b1aW1JzSDBCYFf4y
Wrk2iBEL9DkLtmDTdjcSUcXnYldISdwi7NNwILW0lap9UkjSHa9pAvLFcXnysKZnUzWt55QyDuMB
xMhYlSk9QEM0DYcLUJUBP07XfsQyXY3qXKl3IL32rgWpBoiGsvma2UeRcYXWmuFG41bGiA+rifpi
cGpNYZ9vN3QPiJHzfapkNjBa2h5IwRCFxCWTrMX5MmvtnR5/EAjI1DyPblyq67ISTLR8NZHutCcj
ixc1X5Iprcz+OFP/IU8QBBIuV0hCz3ArBc2FTl0Uz8Au4vrKxwwYMqZUaUagip8ccAHJCxb6lwoj
hB4Y/VNTkaCpL1OcfjN776xMRuVT76I4C3r6UCHYtIFjbvN3wFSmGHozzae/6cGBhpy2GUx8ck2N
zWWbRY/UfjrdMbLZ25AWJ3ns0mOufS1ErGm+6kBrF5eY3R++1jzJlWYArtf+hTu0SMAyIMeap4xr
dnG3CkYqqDpr+YWq9q57NaHXVKx7yyHGZx6219AJXSSxkcdPjZHozh6pxCdW/dBnF947jZlBXI7+
5XSlbNOseRLIEu6qrAUfpS4jI675gEuT0iYrSa0Rz3m6S0lUn6s+EUtykvREF9TL4XJE9JmGUD7N
tCrCs4XAEbX1vTdM9Nq6sbYpxK5doPg56GcnCke6yxI+1bjGPbzT0Om5sgYDnkUBIG1aE+8F4XXd
Zt1kl4NbptldX6kq8Gaz24ir5D2urWdr3uyIufLf8dvX6xIYVODK3FYO3eGEsUTKJMIv9gBnhxhu
ayRmtsLhRqXQHpaz+xcnqmeE/C2cSAZPmJlxOdroaci2H4m91Hk5DmCj+Yx3nNj63oGK15Ipdhly
EX5QGMDTSwkdg+/EDjaREaN4IdVBj1LzGzA3M75l5puQyduWSkRWeGhGZEo7+EgrJPAvPNspxOGV
0pN23wuBwRHlUj1f1Cp6YrZkvINrWHmgdY0pXzBb/d63D2ORPEm4UbzmEmJHK7X9BLcFkskCpBuk
HGdyixA/XVpYMn50rPMZvL6PO9SqMBntv/YarGYIyUMdWLwAGgVSrDx4v6+4sAOelU7D7p9zgrVm
xkInpiNy9lbKKnXcmSazJpOVN0syz4RnwbhJaOfQkI3ZaR2CuD/r4Dj5P2Ka0AoR1tvosxJvylCF
LywdEn9vwMZRABzNVNb5Dju+T/xECIoT7/iy96/XOcSrgdq/E4OpsHV4WfrV0/QVfvW+IAb+v/k5
gBgbfFvuwQ7YlIaM8FUCqOzDG/l7yXpAgiRWvKpee3vSJpe3217zP5xOsPt7ODEcodxRr4nw4eah
zfrArr0moP0o8TWxdZoktlqFB1zhUSbJTCal367Gg49xpEB605bODYfCBZnWoi0A1WsighmI2ZmI
wdSZYBnODxJzVYPDncc/EfZdXncBo5HyP2KYBn93I+EcMUJfnBuADys0p2baoF5iYETIhpsKLwzk
A+LEGB3sOC5HX9wSBTIXzL1IEGsEGwP5ppHU8nV6L5fE8AMIMreu8wG96hTZEcJkICtuYHT1vaDS
27OEqcBEumOvtwpGmElU+xiiUt1xQKr9YlabGTNz0N+SB5d+A6GWgr/FDgnUnUK+vCcqO4dI767x
xA/iMzhuYafz9ZaOP6IEzPK0N7cdXI/hpF/TLUnk6BlVbMtXuWotiH61ZfWXhDexn7wS0JLrryTH
KNk+5aK7Ye179k4qGtQiEF6FckfMzzagU3a+h9pq5WHfAeTa/az8KPRSg4AljCaVK5SxMY4k0dM8
DzdZjNqewUMadd2uSV9A9gO1v0V0R5AqmG0baDsAK0feO/sMiio4Cql2AXm6X0qu4SfWThrXiHpW
AX0pViVCidAxUZzSt2F9les/VPMnvOpuds8tBzGbpkU5/w2OMrPmP/aafC1Laoiv6G9MGfvxzqFM
rrwfg+mh1EqzMHMPRQU30eZAjZa5sNv6NBnAhTtSjJGFT2bdRqciQCO4foHtlkaiYkUdUYqpKesT
afXb+3o63Sep5UnED20gvJ9PtcQtDC8DwfBhs9YMozEy9Kg7BzICYhyxKoV35p7fPJdc2nUh1oBP
Y+04VzAviPi3AaaQP77AZfIy2rkqcS6R5Or6tESz+PXze6ovXqVFmVLNLcfU1fVNDmPI0LfQRH0H
W/te3R8iUOjnJPDyS2KJ/kDUMN5zGV7W3CtiIjd/eJc5fn+rxq5GEUUXWKsszltk3IyrWmOZoNow
kME8Q0aUYtOFyfUdbyzvEl5wKcJV6E3iT+fw2xHce/MZpwPCyNLj3gD1sIYfBemoz5BTE/8Xs1aS
RWNEMJZCP//FndaRLvTeVeCIBDhH4hmU0wBQ1DWvBOnobWdryQNZdGHrayLEGMcNjMtpqYRdm6wB
jiJD2ONliO7KDFQVpBVcO4TAe9M9efPV4HPwGMT6jcwTB7K3S/dUkXFRciFWhqOpXVBESWSwYR5l
xLA46Qc4mbtljpO3bCyNew2zTN4ZjBa1y4JagDKwSCP4BYo8BXsWO3oC0b+m5HQsbRq93Ju53dih
rMuJuTvsmteiz11XGZOEy6UjIPCgh0HTtS1RGyET5A2NZHq5mnUICIHepNn5WRBWEFGVFrXBtX+p
05DFaPpYCu1Jfazr3Qbs5rUqF5onRZ2zM0z1rNujyKrL7go1h749PmzejJJhCHPc6kicmB3EzENi
JGyeoHGPkgC/IbbK2DcdbfQLin4fbaGa/VX65V6DVU9ZfI5BL/2z0FHluGxkyuVaS0u/6hP1FcnA
WBDHt3242q9FONhmKtKgMG1u9EVxBqa2UWME1CowyiWgSG+dUQf9DCPmQ8QhpqMIHw3u5Wxbnh3+
IeL9HRSOFWYZliJ8Ui3UcKQ0d5br28L60m7/xjfQsfJvSxOH/+pti9Hz70wyh/48eD4erTPddBqa
DaNpCkSMFiJMLhow5/SsQjPko0eXzOhoVpz7pOx9Ij11FQ2b9BkT8zniUkrU3hQJiop55taRHENe
KEDRjzeTdKq/2oSOicMp7p4Bn35ceiRLY+/7fPFcbtCHjuvMLIMQ/3hgXtakvcrum1Hz7+QHcN0I
O8sTqv8Z2tIXCzbjrv5VYihDO8VK2QiZF0coN8QbUb56OsddK6U3FdA68bdtICEbyjcFbjv9Jr22
duCQVFEOvIiBPmXU7wsDhQhZPr4VCcdj/b3fINCsfy4OSSxQDkKGjrDYmi4mFnWc9ekICRRZzyRg
khFFvznLq1QdkWn03CwuhiH3cgouLzytTkCC8KQYMeW0HkC/TNWMnRTHUnOscdiMZSba20fHn7GT
JQblikqhWzePuWQcyI7/WwGjWhqntG3v4Vst8LdSpwy5gV+o2pzNsxoU6HpA7UW6KKKJAdVF6K4f
2zyYxMoiWflcjrtOkoa1k7Kd0hO2Po/jEwBI5+74U6VfFdk2z2ltH++5CCSnWotsv30/WRGTFeOh
PPHQQg3a1h3avf0ARv3HG2pDR/aCNik90sPW1O9HcQJcOwSu2GKUGVuPFKOjrTjhOPhhcHRwWRs7
tWYq9jACKITXUh4r+3bI/j0agzvGuznIpLvql6vZdq7cdZR6Yab1A4LaCEmSBe6h3VYmRxr78FyE
HbLEN5JWwGQOzoQQcBV0AmErUI7i+R/6ikm7AV/5OZGIiadaUjQynTG4D6DVB22kawvnRk8KLWC9
1an3moV9jul5VsbUdzoyj9sUJ6gPs1C7K58maptKZWnf/ug6xoXd20q8FG6sXcNcrrMvxrH3X1j/
TubYR7vtrUt4Ci0yp//+Ka0Dn9AKeEGfcaTaSufUf0j62lhOYVyX3yJkxPtR+23GxGEzzb9l+0hU
TL8xqsejPU7cfHY2wBggaV3pnr+eDDqfh8GxCkomYN2UvSoNyNm9RwJOLjkI3Af6vrWXpUPLqPhT
jYYhRq8RmEid7UGriAn4pNFo3KJVAokpIlYHFW4TiQEOBhY5WA6hYxiGrF1+xWR/0YUV3HuX3ArK
xsX062prxjnSVNx/CcWzt6/2PGPyTEuq52Erzz146iX+4329CwMRXSPtqcptV/eG6TBE7F6g+P6F
D1C0BJkTzN5tROMpcyS3qJ3L+2fpkbRgY8AkWnOCzhIlf87KpmHDz755SgNncagLJoExkMf56CS5
ht9NeOKy1WLIxGgYLmM5Y/Nl/utidwZNweCAC7zDD6hrKNgRKh+4qRFGAAURJdu5mErSYykxPmRR
A+doOzZxNv4u/7MA+C7D1zvNLsiuvmwiM7VpS7xtMzinwx17mW5pxESXVgVZqvStEhCCrifZSLzt
vuNro+ATFvsxI+9SkrqNB6cxWQGb7BnUH1v1IdCcE7tKA5n6HTPeAA/W4mP5BoLL27s+vpORmvQj
qVsHwTDz16hjyBojJhjFA45+uDG6BBT5zv6TI25WTpF8hk9ycGKNCBs1u50CHXWWwy+a/HkaKPa3
n+Q2k6sw2Kn1QTSkiQuKoBLguD9Mt3neGrlR7ChsMK3qu4/37+Q0dfoFpdNvugLcZv8BV5x4IXoA
Zj9bUgbTkE5ui9JYMWuJsoTBhdW/iv1XO2XjXmDc8qDhfq16Lye5r/Ptk7ljZEWg2fPgroE5B3fH
WRitq+6zqNrlMDxHx/6Vn4Hg32A9pYD7zDVL9lEaDJtlR1V6CMGkRMJBZve1c2OpcFBCjox3JsYH
NUiCXArmRFz1mWGoMZjPQ04rxxG0Z74ldi4HTOGpMJ5/9gX8Vzu8TzCT29B0IUDCeIs+BQTDbg8y
WLN41C28RaMebek02t/cONvzsV9w/LJjniEZpGc56ziPZgFrAXElpdWqJw9oFzfdWLCAyI9sCu96
fnxQf314HrkpSUuzjKtcxsHXAO+0tchGXmoY6iDQGYvoV8kVLmX9cDzypinnj6+izjptEyHeja7u
CVpuJiF3d+52PCBKwSWgmDH0k0QS3T/F24PkHAGlUAstDS+HhhK5hXjJUnIiqFyWten9VNxI9xdU
rmGDG1pM7GiQZurjhcMIwoUr0x2FC72iu1SAYKnVbNozx7acMhnt+L48Q5nuXhpOh4aIm7FzGxX8
hbK4q4SrgD83ejCIt2Ss2yTRjkFW3rX7lGhmb7rHnAkcTe8g+/wCy3bJS1qQyGuXzJKontF7silK
YtWP81Ulxxo0HcFhwnzmq5XNpOm2JyyJZSo4OIcudH1poczv+sIiRrFxKYiO1KzNafDTL3PdiF9k
ykhJz4zht1ET+3SFroC0SZEaDaQjmRZniickHPw1slGb/72XYd4vhbiXdNuKag9NOthNMSJyDRD+
ADkW+un+A+Nww6G1kvb+DD8txGwC6BhDXz8h8+ZFlKGcKnshCmPxF80NBTTd6U7wSDpd1IPn2hMB
mNeyDJf9iG8UMeE6Buolle0iGwv3BuMJfR3scwO66qTeeyid748JpzviZPjEp0KVi/KdY0inGgUe
mAYw4m8+Eea2DFvI6CC1+2qNyGPfwXTGM9tiF3jLXnVtyzGov5d0hGHCy839GjQ3LsguGJzpqTCw
X58KE7VcnJHPBdNlB5HleA5kufwz54OgXF4jXVYYwpWVOdhyXS9yiCDl7KIGhbZQYeLGIOTMmIla
RGyyxD8Tdo81RLAJbsayLTEQEVLXuDFEX3x0sF1lJR88J1lhUhrxqVzBlKchWONwmwgP+R1xejHg
IgcNVCEtvuet5CnlbeCqprbI7cji3EqLSX0NKOG7eWRi+XPAwf8i0CRfX7Eza/VdBvb92XG0to95
//Liw2EPiV7hD863hjPhVq1xOO73L3vFo8pZiHTOCNK8JLFa+GDBl81rvjaLBI35G9R+aWo9iVtn
4dKdt5YvWHq0wLbrio0UkMBPh11N2TsNXai5Ms94FhE6RwRW4/UDgPSwlSYpqWuO1YupB45WKHFF
j/QPYW076clP2fqj2mVTpqVs93IBsx05R1tuB+lgd5csM7+n/fgXwtgVCDCe87WfML6QeoN8o2p1
HRnR7eT80dLmi5blTThwy0OtG/97cj5IWjEXXOXBUPTqd8CRNuAXV7D3pkvEUK0F6w+FinbpJc/m
j0pynDkiqG65L1ZghBdv9PELTAdvkh9YFCAO3f+xZvMphhlMeYeEHox8V+YCAt0obRUYCT4U22Mx
2GMwj3ZaUzfMp1HNwfSnZJ35ex4rsKktiGkGkXkVQx8gFYDaq1yM7KLaKCfZQYCfUzHB8UYa1STl
JXsA+zvMfgZ9Qa1Gx4G2eG7UWIHovzQB/+epsTWvsbdpl5I4El2dD2gA5yQZaunGVw6GmxFJrwzI
rhpEMHfY8fFjREjqJcCCBmDjfcu/qgw4RyUjM+P049lWk45koRuTVth5pLE96LtNR296jWXeJxfH
YlLjzqYLQ9U0uutsyzpUT+gdOGQ/1pYvoWx3nml1wSKFdP5AFjm5lcQxNgucIXdNxpwKtjHsZPBI
pPbyF4UtiwML6yS858XOv99fhZC1QNuZUYHDeIZQ7SLanRIdQX7CN9SOcEJ2A83BjvmApsw8Szki
NETM23kx4PrfkQIEWgfZ77wJZ9Z7ItX4jFxosoVlHgKmg8DGS49TkQeRrl/URkGsMg9HH/Q8tv2r
0Jdm+5P4Mnc1OGNHYilxekY0EaGZ1oQat/I366Y/Jem7zlLH0xrktvhwzk/6FCgKWz5prdiocRFO
P1lnfqux4BS8MF/huhQx6OX+6097k8ds/jZ5fGedy26/FYtME6h+OV4CsttbBgPvlfqMFKVJ8uRs
q9EP5xSIubYebK7pwR7bgrQonV8Ub2uJRVQsl4CydpfuiS+WygmvjUi2ZtbvSWjz9jzSgBR2vuZe
FgyGf685LU4YgENzFV1DaRiED4CjYXLc5pcTzxI9Zk9pojAHHQ6/VFe4fmax+eVEwXjGj79DUxCX
DvOCTntlES7K7YuUgVtFExP/oUkAtWtR5JNXe3Rgikj9DjCVWCAqnSWIIZyPtSlpoMeTJ0r6sOWY
H/H2pvPuPARXo2IBoyODuW3i1+AMEmS+6S9HcVOR+9Wd82fj92UHr/0fGUOULcq5NZt+elgjnc4G
794IDQIXMI/eAsTqWatYFqMLL2BrYJVYWPYa+VPlgWlVaCdOY/7zdipjqv9Xu02bBko77C6gtEBb
5A3XQw1QVWPT6tMKK2kSWGLuVEHRdVfG+JMZT59rOUelTP0TVkQv6poUIYLG5MPoLAlSFPM9LhoX
2mNKpjQ9Ivlsz9eBb5pQd+xj45h88Yop60ghLsGi6AdJlP/1wqsEyqv5Jn4J0B+6iKKXzLVRlYY8
NSaD44nBy4RYKneHnnsrLtlARSGzr/cyGtp2tHKulajGhIzANaWARqQ4W8kkUIP6SPwGquuOR2r7
KPfw/WT/FDaQvygc/vGxf6k4a1/um8u+rwP9xhxlwmasWsyPpbWgqJxEl/J1ZPiAIkVnxhVE6d2L
ZSInyqOu0G09iMxnqI6iM+ahfNxc1Lh+JtgckWQNcOKn5+0dbzsC8dh0ZVbvFNtbbuNQKnUQb+y9
rH2fRmXuis77YM8G2eqzuSbMyiMW73N0HzNneb8ld76UnYFkngEAXLNQJc1640bjvz19u9itzIOu
U2xscZ02FvmSQt4zA1hme65FtCkTpJkrbdlgsryef4dciX2JoXV8QxSD/BVu2ksYS+vh3LI1fM92
qfDsWwVrMUBnjqzUlQg2R7PzWLFnOXYBq6G8vWv+uagh1RUT12JB8lS6/y8nS30+YKdyP9d+R6eW
c+oc/ADHvsE9ZhF25R5qql3S1EFIldMl9+lji8Gmu3WgoLY9Ojh8/hU00/MX3WX8Ky+6+pumRrCp
tMrGIO/BZctu70MqMqRSHTrOF9O9U8qtUlZeqy/1LKdce+Pdp0bQxh9lzF/r4Bxn31j1vNMoWeir
YEEO5dISkztBxkec+UjLyBWq5ND+NI47u/KsTHc5RlmDhGdB+MtiY9Py8o6iBA1bzSOc+0wecJFa
SjmIO59AXRJCqrDNaLwZop2kjAyXe6mnmFCOQnSI/D9nsODU404XSCk96YUepFYCVCy+64h4ovGI
CghMUR33ehpcS8ixuasFp+6cg+e6R5J257nUiYHb6KvZsG8J5YjIgnJVJE6+X6kjvFTaR6pt6bgH
+ooacx5WZJKc6sBSXV+FY3e5/y/xCJ3mzHHjbwGzzvTaIBQJZSxL6hDVANwVofwGV+y/XYmdpK3e
W/u5JwZS1Clg057lRd1VSeZVuWNboDWtUmnmFdTRKL+F/c0gw5IOjt9jE0rk9LOWoqiX9SNn1QkU
yEyOD6jS7vOhtZSVG6Q9tYld8bgsUCdJJWFsJ1GCwiKOPU3kmDhFpOsokGttPOnOf22ncjzyl08h
exXX2Kx0SL7k+9YBGiJJGrL9SeyRiNWmj30YPktt9o0hoeIPbzvY/SQy4btpx43rBn5SDCzLB1HH
dTFYMAxMz2rkN2wgWjQ53DfzInqOwp3DJtRDjKLOaVITtVKTBuCfrPZZcaekT1KdTcFXCvU+M5y/
uzIUmMJKfHVutWIdgVt8M7bW9XuSTc0/sTXyWKlD8S5u4n5UdN2ayRrp9666nWHea/QzcrB5cayE
xPuhT4DyX3pA0ZiPc9Hh2sCa1E4F0ykyt9N3FN9X+tuM+s//kyMzODdWl+a8f1dJvZek/laGgaj4
S2Krj48kkw4mjaIa3t8JySZtYAvlgGaig7E3QEZ/fw/KF7f9/3cFKv+xR9LDCvvnRakfY7vnEzC0
ftMQO451jvMj7rVh2/juJU+6CtS8CXaGeb3367Rrh5MTU2JIi2T3LUFisw4tlGAbeiAODrI0Hlq2
OVHmQXNR6wK4C3nCVs82nEhAyvHe1aXkO+xAC8IXJbURXBBI/cdNbdIQ+Ikwr6LOAkRdCxz4nXDD
VLYwhTB3FjzYAkQ9QHUXXOdqyXGXYy/yBCVdhEKNyb8wi1gCH8DHgOOZIrBI3QN7UwmCx0Bz8xIR
q5MthNKl2Xxf+Avbv8gMoRiVFszKl1sCeM5bnhkBlyh28zpzrrCW2QKsRuUQ/DzM0JixtunluQKs
5mxR0wrKYkql9ZjVeipKBsZy5SiHKKMLuqtSIiH6pQuCtdBA+ZQbTlfch/7Rbu2NeHXRxiKEBwPN
jk5alCjNoxiKkujEZFXXfjxwjTMcP1oFK5dlcx9d3nC6jTggjFtVl83lqldfK+4EJgB6u243jIcv
S6MKzlhAvYSYf8g2Ex9xzSQkDN94EA2VOyzK3R1mUnF8yNE0k48HvY9Uww+vBQrf2NnUUnObL3l9
759dM4MquW5skPypocaRjpptgVbpLHOSYNKR+dEI/Qm+g9bSX38k4KTyyMxKtz0TQYfNzieOqKKN
wg4es/I0Y2uGcv0ozqpVtQShjmN8SzEjP8JFRInnOG37/cL+ND4v0qUf04HwyrJyo4Z3jgzlg3kn
ZwhwCs3kJ/S72JeH4qY+cv8y/eSerA3x6yNaotMLVnVy8SpyA5HrrxdIZimyGTzP1fqTN8pJu6X2
dEgIgAnSIuwfCMZMovH3XxF1P1u9CVNZ8rz2DPpub4rQFqCXNSLPUk9lBLakLCSDjmejWj+yE9KK
VGDNBZ8r/gsd1oxHmBGEbrgwGeCBtGrEBTOtBPi2rZut7o2NKVmReasKsalP92fA4VBoMT8JhJvV
KROCH5yCEHQ7FZTQJgAqfEkwNUGLov0HqfEq+m3f9oRcvC1dS4popGq+h8HEEe6fkAPIaZAYHlGl
Y7oRGRcdnnlOaj6n8LXJsBc5QYyB+TVvMrkqno2rOERO9jH9Rbm0Dw4KxIQir3mAYJVILD5SzISC
Ee3LA48JBySitlN9vX4gklSy8yXlu8jPskdqrqMQBQ6NcCkrJPDddS/EnteDd5GO5EwoPd9xPob9
rnyFZ4WlZ8HJ+oH6/Nl7u4+GKArw5qc46Wb+EkHqhex7cwAiYVhoWU6yPI+0bTwsOshaNJAk0AzL
RntGg/U/AcmLQVSfgOUi+CNLakBTbUy23fT6/sC/u4M7IJH7o0lnWVeJ+9z0zpkqV+wGSdE9Uv8H
QG4S8nbDcRWL9eCny4oQxgAaGv0dkyPN1QMthjFfEq+4+XfppPhqWKp8TT2pFzprdzTxbLolADiu
em9/UhO6EFTtj4HY8ul2gZCAfq0uNS7cyXACBI3FqKVJl1tlE2U2LrzPXFR4CKNm9RO1RaCQ2XCU
Wpjq+oSvUsWBdLmtZD517JMXqFF28+L3O5MKalmlNsMGk/XugPDwOTVhZTc1+alfpuD/F0t/hPND
3VyuAm2PWCoQO8Zkx7q9J6rdGt5DAsbsCOz713jmqZwHoQm+/Yhwpep1mDLm7kpMo2PqCDk2AAJL
yDIC+Isq56haFNS64jMfrP0NEcq2rZGagoHCySmR2ov+Ap1hD+dOjI8tN/ZxK/f2HklY8ko8qieg
B1dQojmQExMNfsDvOD4B9dSbX2eou9hSKjD6cdVZisCKoifpUNgY5JDfw1KVP1FSX9jpwIAOJN9w
FhbixN3KjzNOobqDx2gdCrP0niYijOCwEP5iNCdG3eHK23swVSQAQFw5A0m8sIf1ebGPJuvfC1lO
pF/IcRYnzTZz75NN4Tvk0AythAlJPuIg/cwv7umRdT1VKB4ADrv6HjO3HAgaPwhGKNyknrP6ULY/
dN5jqHScJ9PYSNX1lXyxthBZhva6WUP9f9HmPnY6ppNp02StdlPjJAo2cSDQGil+i9ueIWwWtVzj
CB91Y6f+lqmHa07qx6aw8Fjre+p/9tuKa04FxeP1ql5Q2HToliPjH8fZMnv3qDCD5LTwvO1V43hh
jVvYA4Ur7uA4ulEIG10eiYEP5FjgzEmJDtr0HUZska0B8xF+/vy5OMsNiYHHD7MDl7D3E569iReQ
9HVEMjVk21FwnMBObkFA0EnIfIwebCN6rT0GIaQnUOxkTJzK14By83o0Xllpb4yNkwENorEVal8A
O9kHAGwYevijCsheM6N45z+oPDdi3x5yxUQADUPKB8VlFnVbM8keeSYvP6Elbikd17sVPysdVchj
teZSW8bQaiVDJVEjpEzh9B4Y66XV714MvtryvMN5eSKoH3IIBpNR5d/a+Jmzy4BJQlmJB0rp5gpx
lO7FqJuQoFdNtjF36yPAAhozYcIAKi+SINhiHQpRo4H/69AXxqwM1LBmXdgPrtO5fLxW2wci2/9V
S9LA/rV+zhpExHkBMA3E1s67FcFoYziA4xOBPwBtFVQoqlHzT5pewgUftP5b6FeGH/LKz2dAZKR+
BxlBad6Bjq3zprT+tLkyorHBVnPcM/hie7lJlKZhz3JxFrBDdtJKb/t6jx/zRpy9pD2tm3PRFidm
TcLYkAHd75Ynba5uBBqKcVhz92ofHdYnD35t6onfoXvKy7zXfVdNMNVFjZuJ+MknyUjlCqvx5mJc
aNkmPB5+XTtl+lBCJrnLk5mPeWc6UGzfawlHodOyXar7pUsVu60E0IXTTs/Vh4wvSGwU5uBdcy0m
cHfM5GtxZjN5buOifSmisog2JHzIjcAFNJUO//xAVf7t8c/hr0cU4R8Ci7czpJxIKd+aMLhNZ+Kl
YNcXuolTw0E21j7Eb5F5V5K7eVyG40HcA5PWR6/r9Za+ycHa+z+i0Jy1WOd3LFMjm3MaAT1+VQ+L
lY3Ibn/Hxb8fzywm+ikIi5IwBZq2LDrprsXjW7patjGulV5w4Qjzmq2bHOeFWsxk743Al4tctJMg
RXirAnKg3RfY1PkuhNUXIRYCJRPKor+HHdBmp6u6U3ajpIarjHA/2oqhwmEYZQP2wsSQnLXKz9yB
jzfrZQedhwhFcX5igIzVzASfVhM60NmL3klSAn7GdKctFHM1S5mD7iMCagSOPsNwC5wywH9CssTg
2giUwonu91NtdEgX5hse/M9x7XXNT6Fy6o/S/lLjZRM24pjdfQFfDNmrFrywGXAtuqzX3FSAwoy3
3C8NN92VY84TI1yfcfdJzGkXttG13pNSmu7xGYEzmERenR5PvbkgY08HE7n7cpuSVfkDezVTIQbu
4Dwrv6uR2x4N3eyqc181cmpBdfe8+mHal8o03YqKsjGs4707gi8NHDCgyVoH5v/eKyCDTCH4+r2m
4o6Brgwtj8eQDjdJiK9CZA+9fenGagH5c6kI6/5cgGGdez9KxinLkKdnG90MWpUDEevOB8YtfkQ0
Mo4B6bYJIW2QNPPW/gVA/VQ642XLB8GLfg3H5H4bpKPdk9sm4SVW0w38VX/ZIGCukJmZ+zmfJssq
IAAY8ekbOglTsuXNV1ZISWHY6L2v4kkcFEFzN3XCTusqnSTgDMbhhDM1kF3540jzvSv6DgkFqJQs
pZYcAPsCgKfQY+kxk9j+eK5uIpTW4z5YXA0jo5u1vI67MD83ZLJviVqwpGObMmf8+LfE9g/g1jq0
jZvJ0TgoQpivAg4IbcQlMthAlgUKEbCEnoxhLKETtKAdUYseDtSyxdpFVlas5U6w5OMb++GfhreT
H5TwuW3Huulw1UixSN9LgX0NVnLlllBFQAOkf6K96xmzv4d5SobNGxrIgf1VKrYKaO9NnfO7RjpP
gb8Jfy4984ZOtcI3pguOV1Dgh69SYyzFnizY7W3uYlcyMXv9G1CbPrcUVOlAeN8t8fdtH7KAVXYN
cZeXCgs3qHVQOLmEeehbqIJOiBNBBvcRp9bxbvMMJTOA/KTZRz4HYBa4cAa+gmshTQG9TeGGWTRf
SISuhhPQ7I3ezRiMUtdyuXQtKb2eL33IxuVp9b8rWbawqTNLfq9EcMlbRg0MW9fuo+x55Y90w5rp
rZ2a2vJdypXtD+kKXDrDo9Bqq5J4os413Hmt0EEA2c1zEGyoTfSigl5RUviSwO+uDjhhJmvE6tAa
XqI33ZYvhe1B1fuMNH462qfXIDlI+00E62oV9SmzZN0rSqWpA6JMY7qQZdyyW61HoZzsQcA5OV8W
oZ6rbYbJWkixu4B0dmkuaiapLH9Z+AGR/fnol49y1rfXQehWb8+Lq7T9lk9JVHWRgz8ECkvNQFFE
X5phxFtCAa4578gNND11Ao7VTF9N8ybGpr+SELrEvv4AnbXhh9mvdNQHviDhFtwwu4p/PkiTUKsq
pff8Z1zPWGj/vDIbcPeyZYKDx2BTLTXN+F/v/0PUUEf5V25g1YGiJLjHl16SHssrMS1CdBc8r0IW
5w9a1t/ZYLDMc6165+7oTzctTWP4CIU+m27KA89twNVK3PEZB4Ko40TM8n+TMByZwiv2cIBxOjgA
diXYMAMQ0b1W5EjKdijbf4itw97BBMGG/ONTLlvPmhgn/3HFhVZp1vznxk8c08edbhBNy1/QoBrD
6TINotX37OfLCZoR7cfBNqZzOXgo2nVIQmN5xqqk9OTKfxtBRQ0SW+4cGF2NYrMG2W1uUMuzbpG5
BaCH5d/BEYtoNnmabC+6cKINBnHg7plbMobf/wXLeXmMOF2iZrofEI0bd9NYoJsrqEOBwnD9k2fC
uGhWljYEo96EfUmNilfq0GgaLQNohAY/KHe2Fxhm3Y25O440uH2BkdTIafkNfsRzhDlP4Aykpn8Y
IJM2/XEqawssK+qnD7ea4ATKqaH0IYf1ZKeLV7eA4GfnWQ+64d2oE1HfEsgYrlnF1w4DMygpYj7y
XCvh1LmtvkoobmIhlRMG+yYfkUAbpQSVh5DPzZjntAR7gUc47j4yHZwVtb2if0PBO06xsQ/0qzNy
nRHB94FqLgJ/Zzelmfy6As1ahJ9/DEpR2CrDKEHeSWWzfahfelC0NuZlJX5/GYDq+oUdj4j+aPg5
NF6Rug1dmme2UNAY50+n58Fa+l+TXHDk6qP8Eh/PzO/2RfYOjLVW+YEXEMGjuArmzAXrJKDiWj1+
triXq1g3YMxs977G6BryoYkbLWoN81CcMLCnk7YL5TqNcE7/rWP8T37DYU2CoxlZAmDC8eYDZuXT
dHM7tT39Jz0XGqEH2dMXMq9L/FJZhSsghXU8sg/2ItflePm6SshgVhluiv7Dc7FkEUs9g9YVFr2y
sEnknLM5Tlo8C1FEzxCtZOySqwmueBHwOp3VRvWeZqWy17WLtiOv6IJ44Vygip1sXlwblRJFjfBu
jGEEf/gITlDArsbRBK7HHpZdW7qxKSfSeAusWXgdqvpKtDSKCQHlGY91x7eUHJxvPW2NsTvg+hu3
UGToPeV2MjA8jollS6m2Qcww55k/UT6CtSJcX0M/ijBbqX+HM7O+zWSApTSagQVSOP+n06UhORJG
R1PqRaviq/po4/IJ5ipyHOih8H0DIdtWSazfuy1UA3N9XIlH/fX1je4GqKKG6fhimdWbuRDBLjsr
7yQXi38Uo6s+XVoASAz726u5zEbpTnJJnKJfhDZBPwSitYnX9KOqfIjXeb+x/GgZPb9YH/IENfwt
76e1kef/zrD1QltDoRmULcBdP6Sau98r8qGGllm6Ik9DLww6stKBidu9VlFfupdV9G5yhy/F8ml1
goO80IkpNojFqyromrZdCAiOW5T5Ubr4pI9EvGcWBV4naiyOyxoIKcuPgMjYHFtQPPipaKh+OEOx
ay01McJlPYVcHM69h/X/IJW9jqU8PEzLW3QwQerY2a3m8J6ie9HEmyKzMHbtq/1dqfa/7uYYt+Ui
pjZwpUhj4lpuToKsydl3rNkcg5mjOh1LZw3rX810LJniexXVqR0KpPLuiKrLwMOf01Jf51HBuxjG
hCZyBdRRf9Gc/zfGdSJHaBNHkvZ5OX/usun7sxkOmjZnqMYLy8dkkBBKpD7yPWombJkNZCR/xSCs
sqnuLM7jn1AvZKADxmzjvmOFjTGAFGYKFql9CrWYqOfevjDotgnS6IrsXOLPHhctlE6tRSAZShTq
hNVhM4sZvgZINr6KiECEYZO4QGMH0bYN5iONWrMLCgr8LvSi5Tgi+J3KwnxWYMjEmLjYJtCeOs5l
NktTsawX9sNO6+LmvR5ZWX7SWwomjQt132dBsLr9lKY+7Sz2dRZUfK2EXLMTGx2gI2HV3IHwZv8i
rbwsUtn+utsBHM0j+gl9qbs8pGksPUErvOQHKg93OvjXtrBAEXG71VpZKtOYyQ3Qn1nnO2nvH5BK
3LyeJ59k7aDJRI8h+YZdFvonYWDFRBrQLZD0UOJ4mOImb1Vwq96UpNhGXO0aBzTWXiB6oNwTKpLY
2DQ8xKgAVFAXmjSYeC4MLFe7+cupgGdjGbRCdfZyTVM827RauuVBw7BvkIKTNZQGIXuIO8qltTK4
JTEjCYLm3nfsjUuzlE2ljYMh4pBK5RlY0dG5YJOj1u8ohhP62ElK9gxgi1+9/MPo5nU5mJK9mdJJ
jx6d76aywMYZCizZsfCeMntjHTJ+Q0pdHmvsWu9bQro2MeW/uOaxj/QGZo7rGATWUcNO6lv8Hs5c
fHPz8SpwdfsFEILYst4Bz4fKVAAYu3E87IABuHeg5Jzh5q10Z7SaXIjDfDBBXnm6E966PH84YRH+
DD20hsAV0Hqg6/EJtxqb1gWg6OTm7C0PI5QE51tDaCSBcF8NomWAS4GzicZm4qqwNS2eUJPkfu3W
PPBoKOrPE0pDoVDtJhf7ku1wPUIlGnQZ4vbIoDMwrKKyI86yhuPqbavQg5xH3jZryCQ6o7hnVmL4
1l+ExSkcCdz2GwBtD9cJ67EX0YIyUGZIMZ2U4VeU+dmVT38JnCNnwDhYKzxs5FzYJUIBzNVbiDRq
tH9R/qKNUxT2S2L17Uae0qvtz+fmFnAfY12XDLmfr6CqcAVV94NIAvoAcJZOmdMLQayxq575C1Is
+t1q/aXZxvzCrSiBbZoVrUCDzBuPsCeLW1CcqPKQHSQPY3kooZJ5KsbpQJx8zJWLbRBPE3AR9qyT
WF2ZRgdv6g2bAbi7skMX6r32PCNOSRWW+bNIBbMoh+bUivlC+0NxMJ6yaiiTazu3luaig6DZBmiP
TlaAZJCzRVuWtrWpKB+qySaFiZIf3tEALVaPmGB4QjnXxggKwwNEyeYw05F9h4GwxhhqZrpV3NCo
IgNMdfigvJv0t5bOPYsKHVxaSrJcBV1+ZxRolZQQlvMFrk85jB6CxgTmaDKsjur2KP+4MhhoUJSa
2m5lCotWUwNRt7D2Swx254PzrsFdKPBcTKrN3hEURH++qUf/3Ue/jIWL/DYR97qUR/UMxNL7AwI3
yG9bYvbqaKrmKFj3dMPWNlet72KRZRNkRJFuayoEdscwV0naEW94kRsnxhL1UoHwGF/t4ddKTqcD
p0ypiWZBsKw0FpVLq4//IspxBiT+igPXR9b7sZLYyUof9qfrbX0pSG78AQwYiQUzHjcQvsARZCyG
V3DWL1P909t+MbPJ6Mk0XJgyNn34ZwLLJNXWkaFpsCuOLlrHadycVddhpawQq9JO9DvPuNbr2gm4
HyYD5GdjW/FT25XIeGRl+S64QkPq7DL45e2LJUshbA5alCNgqxIaCmhKIq7q0hzgU19HHnVXc1LS
g2qzgHRtMnnQrlo1Zv7aPV4GJOLzcqWAi8TQklJQDCycFvb2O0ytRWWM2iE2dV4T9eTRkFjjtf3e
n1obZv+BY8eYZLESWVy4k5PF2J7NbEAZ4x2/UvXIAHp6OP0xpv4SdTVXVEru139YkPRRjyxCbMLl
R3iY1kZc4k+QYXBP6tw0IDZGA/3C6qbz2/IO8CE3vDxV/MtQ46AwoRPXRabhblDQSTO4/T5ERBJ+
jz068zlW8fxsiR7eKtbPKcoKlt4jOhZ87E0czj/vfJ4GG+4eGnIgmeBRqgdRZrS+Sl/BA9WCatKT
IdyMbjN+X4wdQ5+kHWYZL4dyWL2yJ1jVU//GnBRflcKDOsy9jobYZGVt7WnZHTRdRKJ0keq5tfgb
t9dt2cbDojlMXlow1R8ZDbHITJD0SPTncrWJsYIAYzXncXZMvbDX/ZkIQShuxOVvP+xjrzL3/cGM
JpPSQl9va4wd1frJmgmPBHjylWmsvkbMNmXlM2GADJRQi1E9SIBt3JHiIxKSWjGpX+8UmnJowEYp
rS9cm8HW6wIkV1iLmWnOXnZ9Z+xWwE2BorLO6qBEtTGDSCUdj5qUDYsGRTANlBwOiUdH3tWKl6m6
HGup8dB6eTWFzc4H3N+NYODB/C7CpIVowaSIiHK7GcOPqag8n/uXAgkUs5s0LA163A+TmpVEA86y
TUhsUYyjVmSTqkn9JJhk/P9BuAPVtB9MLDSMsFHjT2yE7RkQ4jkIn1u3fTH/48T6/onAGPBXCfmf
KvTBE7/Lq3t+nYLVWgfDCOfOSq8vQDzt1bNeFLLlQaIJoktoOwjxyas5oEqIVegMlXDwD9z1xicN
MilCQt5HS8c8sYsQAJP0rI2tKAMpBf3j6Q7Q8fh03Y/vztwj3+X176PzWIkX9obXGRQdKjLD1KQ5
fzcfu+OLZrH4+DeK+JE5Bn00oLk8MmoU2vuGXXgC8A78FLoXUaPplfz4MJKLSXn07qubH6S7t8LY
BMmrTGpRd/qwK+Zpc/P3yJr7j2A8589EVxE7vLr0vcTwF1Btvf8xatGs3cF30RFI+kBsFy8n+lkl
bCw+U1dM2Y9iNN2Gh/FzRoGdE92QbIMXR4TtPh2rPKIZerLcDXr2EqS6eQuFgEIZUsxiOscq7YEp
fzFHi3EY1CF/vwuLDwp3TziQnxrUvcLlJEGuLZvV32wdXT7Tk4xqLPK+RYWsJcKOjRi49FB+3QTQ
N7+YA7XSNB6nVDrgni/udKypVPJx0QRKm0sLypyPAlH/EDt1Yg8TpLAXkB2VZNqSxoGGBCElDdLJ
ULeIWz/5MZmdEcINEQkIegNIJsIgQCefk+ephuTHPaJ+K8qnF/bQJLoc7iQjCCj0MBPJiXrXUxB6
bU9PlDy4U+k+ERxNOw0Tj3OJSRrzAvXeBTGx8zVGpIfdwSpE5FdiTChVIoAvjcy82RK8fFsAFIDD
ip5ReHoqjHlAmrUt5R1a0egOm4M9cuevl2V24vXRq1mSp5nma2vXqaeM13YZE7wpn2girIFqGd7a
h73zSZ+ARbR9c06jIgGNw0YOVHRgKk6d2x3w8luak26aWS2w1tJ650HFXLxC1CNCUPIxnKzWT9Iv
LO6cfyuvjXWM89+Xo1F6MBufaN2KbplaCBtWW/daM+Soy/aOYew292uxQhbYT0xf1u7cSouFU5ny
R4WaaHiFfsbuePzLM6NciNdli3TlWBzot3RxYe/oiZBAeBsaa6UgOZpaq0avCo8CrhaNcy1UADGw
2doI8NmezAqzNFmusUWOK0joF5U57DpwpzwUbytxHfwnSxtL1PX9eAz1tcQiHTV5t9sGvFzh7va7
/p4wyVXfNM2Cmgp6HNZzPtk7PYSHZE9XYE5gd08OpyDLOagoT58D3DrXzXN+LbK1RCnOGkKEGoNZ
ZLOk61Sk2zqqkDH71kAow7wdr+0hA/mdLYQYa9C4J7JBqPWQok9vZ3s+w+iajwjoQKyQDKwxpv3T
x9Ri0TD1OCv7kSNm7tzgQXh1zZ69nfkGIo99qxlJDpsiRx7XIaQRyw/W5OvR5S6em/qIZm+Zpiu5
rtUj579YwiPDc5EOX9as5hX6E9zKPOCVQFJ+AFv45Cjhtpkl24jV4tx0hmQ3Wz2prgT31+OviY5V
jMqlshWJp2Str5WqSx5GrQdkDDplhJ0t5qABAKa435pr3bYAZ6Eg0XdYN7XkJr0qPjfhKcQrwMy0
82PkqDfcaKx7jpknax7wzFVamt78+NeT4kwTTV5jyZlIm8GJpZ9WFMLGE1OtbpXFRpCOwFn6Uo0i
ix0cIfrKqv+r7IdbkcQwhPIN/cna77ec08094muuVvmCpY5H1aSB8ctnZHOt5LvYbF9B5+2fzwEP
mZLQWSh0f01L/dYL7SPeCq8cMWGQWMBqTKXGeE9PBfBJGI5E5TCUaJyO8d8mI6DzCr03XPpIzyEw
Wk1fSz411GSceEkgXYgIW6M4ekQCtEgoey6c7uRW9/BCviBh1zpaA3Kjyr2nUEU7sv3Wlb1rWtxf
n5yT3m9uOuZIEslb93jISBEwrMteQvZCw40qHUMA+LGl1FpRqYuZi7dwPW5OcFWBBPEvEEsWQdrx
KNU8JdgbUwNuo8Th0duVostxdSNcaphLPJcRdsaO5hYTkVEboXMdZfXdcWBGeVFhBCUkDXpo6f8k
AILYhhQl5HTshLuo+UnoWD2UmWrpYNIou4h5x+6BnvUVyAKHdarm2TWyWRq0SICEgqRALChMl+KJ
uatltc86Fo57oMHYesaxbRlfSFX7fjCv5B+6OnzS8NQwkl+ZyXzsSOxKg99psVmt5v1aEXNKmWm9
IeRx9I8XXcMMvwaZNbUlzGqRbj+QWLHWTPGRHGGFYF5c2IcdnQXh/CFjihsmyPp4BrHHxLq9jKWr
/3/Xj67QUuVGwfvwUnev/qt4/YrUXEJlRGtF0Vct5LGSPTfUpXTTAioPrRd1vCblB3SwMW0BLFju
bLjGaUpTvMkAdiN7mvb4XH8Ct5rJ7JKWJzBnrvoMK2B4fu/PnmV76S6GYb4j1zu5nGpvhr2KhnzT
ThbeoNg/BwQ7AoHkGtosQLA4Nwniz+pFuD7iQ3eGi86ir7wOMhhPTtrEjADuirb+ryc6ztZvzS2X
ZO1gg0pHCZbX/Y6G3w5/pKcUmvm4C8GDQbhhkStgc3to4AQ1n5yI2HJk3woLbN1/frqNjyTXJna6
1eo/hf+Ml5b+SBYf/TW++HSJoUdOuk1MONUUum0KELYcv2+DeipQvA8jIA6RUkSTL2fdvwABrkmx
qPWKKGmPJfupU3S60bcS5L3SRjF/qx32ouP2E/uYCGQLqiDfXLbl/nr1wirDyBK+bkZTEjSraTow
VHXzRWUh8eooj9x1ZHlANQ/1mmstfzBHzKZUW3CqN7o3yYWeFVGr5z+IRuKYa87Q7ZnoM49zERf2
ffTWvGV/PynAyVGWie7gythe09eF4Ym1UxgI7VIEp4iYTgt9a9fqxSLpWJtyj7lhbKufNfSFkAne
+utqhaeI6P069v8Y2juiGTYFMdWGKu+lJJmjf8TsU4Dls0JgJuK4ajkc6afJFGCIKlzvh8BOOulu
xzzk3a0QOqikaMq7zgHVl+XE9v22BUqB1dtt0OcgtT7LpdJ9RuZpWUmqZ68vdazH2tJh07yCgVfK
iP8DhPVXh66/RH0mq27q5SzbtItogb1RcVu+IbBaQ4OpZewbT4AwldjLzxIwQYIrqVGaVeYbqGue
QdtmbuggD4Wz+LL515MxpkiKFsd5OZG7RwxQB078dgHH7kUZZ+sQWpTugkQJC4Qh1nngFo6ILE5Q
n+pQX092d17LHzFfTKNECg/Qj9kVh/wYRWcC3GzyPpM7sJ74BwklDEh1nZABftkAYb3EU+nShCEi
Ll9LZATsVZD0+L826X7MVXGE13t96tkvWT5rLBEys+0fKqQbEp5tYoDd++gzPk9I3eJU8IHrtiw0
Dcrgxa/BxGnjC0GGLg9ZvmkTPcLBK/PPePiZ8TI4Ymv5rdrkCPzgTM24e3ENpYg2+UbfV/xabR6V
avthM433sjBszIj93DRG7imnJz77mWnPnrEoNJl6Iz3zYArKroan9hDcR3ISwSVMUsoEUpAo4NNA
Er+ID0MAKfGA9Tydzgsl7UgjXJGs2LtetMEBQwpTR40rmoKuygt01+aTvXYsHpljnrwjwapSMmMO
J7RH9T/0rY0tYlBWM68+uSko3kFc5lUthTO2CfMVaJyWjWE5Z9Y8HlrldOYMB/hgF1dglAnZMLl5
G5pjoCj1v5TjEn04W7Qp+CQu2kf8CrVnhEdJ8nZoBXp2pN3XHXX+y9RMW/ICyWkP+a9iZZHDCCQ7
LvbT8YKxzV3U7GvlWNFFzHcnCXZ+sm9G1an91SjYusmFYPjcweT72dyQ6Hdz6GxUL5E/k8EX5BVC
JP1asAhilnBs/7zEE5f71NFcICRIcZDn2RkVBzeVSxCJEthfC0vS6fEShy44ZwaxkbAzy5s8+74M
A8/csWjtFLT02y46fcN60WCXPMEP5RLCe1Lk9s04OEejuzX1GeybPZpaFNZ2YVn0ic22SUp/k4A/
yLzdiTSW9g+N8WCDZcPtUfaBmeWuPaAN3TJIz0iPN7p56COgXh2td1zXqw1II4YuG3Xfq+ruZTzA
2x6V2OJ7mvXPknn+KWJMmpZcx88jBY5vONGbGZ5JrSvtaF3LpDahSmiZRuFV+PTefcc1QqHSBAyq
V6Z6ftJBSMg5OIXf7KpwKfzk76K6X1QMyagG3UPjbCehSuLHtF80TpDrAtgmIfh3myqXpt68kosx
f30eB04fH6chKruddd/U+PIDVXn24Rp9XU8vd4a9Llfy93xPpy86T0f95HYIocHGclZx+xrp+42+
GAa49W6ASCRWkmKOuzizA5/ios2rjvC8q1sI3ETUnqegSGLSgWtnfog+M9VO8hjXI7+n7KfVMVYW
EvpIjjBykmAuO4oXaZIdfsScDW+mVbvZZdOBF7b6x1xa0RCatNIs4Rvrr5061pg8fIpX2cEGg9z5
ImVP34WrYpBqrEk7F94euZoRLAZNGIB6hHsBp4un7kJo5RYCXCYHAWSXPHK9MV4e1KN/kkEVieUp
FQBsZ+O0QRVC1e41uRSKaVVup9k6gG7NFOzxl6/+bx1gt1ndnd/Wen2az0YmmCoEqY7QnHOOH2Py
KSUucHgzECgYoPlFvPSNpM2pbOHLJ0eR2Xo6z84kGJtnMoJe6CmVvtaxRg+2Twqa6u/Aqp+6TZYr
pKzoulaB9uQk28dPZwJ/qigSNXXtHMNUNAOPRi1Gl6gJrs7XREyZdAFGQSULa5/dVR2dQ2a28tsb
ICRqRFW6RM/csb3TX29xBLzk2HZVe6SPSu0Y16Fgt2p7MQoVuedWUqwcQ+LmZCw2d83brLTB4Pj8
dlQNyR7jhrY/nYvbiIOBLng5rM6MSdYnlELRlXouckZ3qRHLCXkw7gcIXerh2NngC5PlBxdlykEp
OYObIf4wsB975EbYTIzoG1qaSlinTUD77xEdG1TQENqqfk5x6XLtClLUYWD5GaccjkdIK7dyMaDu
BBBTxRkhpF0mVpNmPIZzO5hbyclDq1tI7kTxrSQRB25TeLI6OxhsBJo7Bp7Tv7u8KBle/FwVtGGH
DMQdaXunv7WqOiF1DZKAD+ygn0vZ03q1tMhVLdQVJRyvl9uq8+4u1eqKwPi7RemtgssBe67lwzEx
827PnuOqJC59PX1dyBnl9eiShItU/1ex/ChRXczOhFHKNoWDat/r0jnLsJpRPuATkm0ctFik3y1j
TUhBBNDzF7KejP45gyjGz6cRqjNzdDgomc1Z5Lw0QYE3kXCQd+DpUdka7WtOS76PgIXttTc8yCen
Y7AiY51ZgymoOkxSx7I91jfvPvW1AJ4bV1uxvMWmkNSO+wB6chf9SLfbntSXvLPIBFrgP43R+rwo
6FN5+OLIvp6OqvrJABZwolbEjIcKXm/42YmfgWZfR5UvukStRGME9mtEGJER6RCnOO00OX2ykaic
CS83ipWg2L/YHO9Qiv5LBdnrk+u9WsxM9Y29qfvEkUDpQxb0E/VTvCRt2EFAdq7RwA309t9yIU4+
GdsdZr08wd50HpwepzX6FQqc/Y6xsAo5BPEPpE1aHxosVr6juHpssYSelqO+Dhe59G5apNh0iu8J
+aKaKoAIaVIyNjmvugHeo9wtrt9c581TZ7QZXJZpQ4dOBy3s8z7oJL76PZDUlKOPH9Qzepm4z8rW
EkpggmaL/g96gO4nvGlatC9wqmzyLbJEkOsopPAAj6OziAVQ7HRZ1MO2gD2oTpYMpaoz7UoMy2Ch
WrGzAG/6jRScFMSkuVq0BFlpNiW5g4gYpxs6RpgyAI7jwIvpfDthhRhQAG9eqJ/fbPtRSNs8f1L9
IpIYWINzwe89hgXqsfZ9WgiNmmsgJHAJWjloM53R1MPlrZAml2AFnQqrcGOAlKIBIDrZUUQ1K+xk
rZ4kzNDAZBX+BCyZSmQh+Jp6K3qPz6EMkk/RNJqXuvz1H2VRdsEd1rEQKtGgV1eFqznndGfF1HkS
ChCo7aFuxhLd5CGb6MyXhPcvyqZmkWWMYgpsy3Red0UC/ZH0p5nbUd5zbmBRQK3jR+7dIta6zOTo
yVA+yo9tIdbFbqji3oUukvRQT66pkI5BoacDeTLl8vylzW2KhKCSQjuCQMZYNZ2jReKQ7WLkhB5Y
VFS23yAzcNcfVr/DXfe8POnvJtkA4alJ4OQpV0LdcPDuHImQzdi80G7qG/scOopeNlRhNuqSf66Y
4AT3FheEQZ/DSSU9fp3AR+tVrHA4NNAjng6eGlE3piK/3SC4JTc8y+Kniy6HwU/B+UUkPZL6hn+o
2p9Twqq4k4UeHcORJhJS5W9Gji/TiKxkdAErgLdcMDZqySu7k8i4N5fr3UQK2PwgIwMdUW3JrV6c
4CinBaBqNQZkhNyV15IV4V2tGrA/mAwYGkg7pslmGAOffgpTh28SHVX3ezvtyVBmIvykQUZb5FS3
UH23uIsfV6cYa3KcfaEFKE9Yq0MvZw8v9xcadCgjWlWrH63Pgg2dTG5aercb2wQXuo7CPOh+PhOI
jPoPkXYIUxhsOVJXqgcFt0MRR8TcOfG50nVNyv/7Gm3R0x+YL3ky/ZGb1SyRww6ZIPOrBbnT7ngK
tMl9Vixh1xg0fwVWMpqOrpMD+atPhGmV/n5u0a9JEY/gitiNvg9CyPrLpO1yre4v08Kg88sDOWmT
zA7bpbRKcf3ioTWxkDOhYEe1fxdfe8BNyyLfBQwQesmgfoozq5fRL5VGn5umMkHZoPcbWeTscuLH
VEb6kKysUXfhN3BgBS5tSHwcDccv0w55whYha9ExRKitraT7oNNJ4BSujYT8K+JR5THhmx+wFTox
8i3qa3ocPUnI3C/6QFz+pJ8cLt3lqMKKKxaKSny6cmnHaKoLU0QLrY/m3Ee3SEqOL3KBleV0FyFW
W5WQ1Av6ZIyEZberNKvb+lsVtyJtBdm0yBjniUBp+RCWvp+O7H22eGvG+wTkmLfRgKOto/UZVOVP
twCl9xlrN8KDaMF0JIO3pLqptNL/YZAEAQUiNtNY+VXyVlegmOF4eZV0U+M2Ciat5k7isCOC54g1
Z5HtFGsxS1kwJJTuV+tdAsuoPg6OdXlOqn5kicImDX4YSQP/hZquOJj6DGVLl4zWmBviWGWhNdl0
EDm0JVCEmLgVeeXfnDg/PYjefIZViq0YQrbuQUXnhIurLhIK//vGwwU2/nna9lgVyMbIZMNpQjTA
23/0FdM1FkW+lze9RVPvmF/3Q9slKjcuksTo5j1n6XxXd1K5VC7YkK6MK59RMALGJ4rYEheT3A9U
MT7aDONqOQq2NQNHw1j6cEpkcHZGhb7VrX27vi+pv8V/T5FGScdKsydhwUZSr3wDH+EZL8bewp1Y
vbh24PWhw3z3vrWh24y58Nir7pBv+nmuA0mVSO2mOGjnyA3T99vYi06JuzNOc/L1LNOQCNT54OCz
qjcGmurAlqc/QXgvg0j7Y8UaTMEEsadds3eW9Ha6Nb9YCY4wXpGuv2RJ3VYKgyJjp67FyW73Tu3e
ULn9IJhtzC6DEh10MHPcH/VgPGjn8GSBCZ4beESt/pVKjgAhye8lzEKs7Tm/uTB2lK2kRsbcyv76
baZjtrIjDySb9zwx1TFh7p9UHUXI/AKB7gvFsZY95wQyC9C5j8cqHQmfSToa3mBHd/GmDFlPmOrH
TaFGrYkI0oqtNIABbc+C4NIoMDhzB3468/vd1vruTV8VSS4J8Y5D3FYmfnlLSNEaxQNxuy+vXIe9
u0ek5HOjGvT1U2FCae+fL1I1kBsqatuKhLFSPwvmzhmtbPSXC8mribcwzEWPmtESZ1Jro7rUDg5r
gBIA1JmbemfYAaxRdDPDZUfxBAthA7OxNsaRpThcVXNpMH5ChstuKbhQ/vKNXTBjnQmE/PQMhm5E
ZJ/G6dZLBKA0k8N2jIX3YIYlAFFCCh2Lsj670LdcPvH61olXxL25GhsyPrGmIPBcw1HnYp+XaPTk
N7Hl4YxsiNtscICqtUgB0uT8g61RfHZP5M+s1EpcPoPyafb7V6tj13G4gC7y2pBaNOWTwrzOklPD
ef9wxiPtRnohYKC54xBByEcSNQBY0BZ6huocevPoE5hd0ELtPG/W+23ngDYdDxkSpcpZwwVH5qIQ
+kKSWJVzBrQcmBUBlYj1Ic5qJ5FOsYtonrjLBVpPZ04vrAdXq2KCzWlkbpUAb28ZNah0ZUbL5oVp
mOuoSgOJuRESff+mmP46xZolJd9uTuxCDfPU7gs9SXgWTqdByVIGbxZN17lW2DKW2fUvlIWjzRbR
DYRSG1fOnB8inAEhS3eMxdRy94zS8J5euNInXxnydEtdAvfvyOFJWNEQPkAnwXnVd9qPlsBj9dNi
ZvDfoRefoSJN+2QXWbaxXEZArw96HlWshjyo/MYQl1wvX0u97S0/dfI1QRJX6pb7OgkOUMZ0SVGq
3U1MQR7Yu/EjVbhE8i64r1HoQS6yVtuQGSle9EKWSO6VIc1iIEEZO/jHPSZx+FEs/JBNCPIYJ/2f
gbTidyMMuLAIsma/p2JZozn0eFNjnM49FjvO+llYlIGH24A6WR0PE/haIiMwbURzq6kL/g4JyJv5
1pGzqEkwUYy0S277RbxS3yBdeMr+QRZGClrcdESXgHF7QsAZAtU4TY9/nqg0TDAtOLc8GKX4Gv2P
aMPYFhq0IHsFjomyjtWRYbbofeqtXnqu6Mo6yjKxgSiDwJPD+Mn4AnrLA7L/oeagVNXpRKhjO3BX
ll0xifPWmcyUt7RSByR0f+8c+i6sGbm6nYup067YlpFynpX+gr8jLhu/ZbxuUxjp+wHWpzTh8g3S
2T5DUV19M4cam72LEwRRdE4Dc3ffObpBzFVPHzps3FDvTMmP9FR9YXIeSdG4t06VX6Kth7PfwX2P
IkIYs4/mvj+VkkscqAjI1+NOoBf7900jqk6Wn4innLdODo9vP2J7wjK90T9gJqoLo4F0Vc3m5H/j
aY7ZcoqRzBFoeL4HSfC774T9CZyIjVYkwb+mdHp+m86TUIGJEVUrYWY7LdQXaUKNaUV/ZEynjXBL
QybitYUE1wFJTjG/7FYFBc/x9rbNh0qX47h8t2QPVPF2RZwFN7VEoLjeB399rJxfoHQeUyxIofmO
+QzcECmbKmeuQjak1VjfNMEDr3AOQz2paolz5B13D9HHzA7UrPRMAc/LxWFHa+i41ovSObrxPgH5
Ma3YpYsVzV9YJXQFd/5r8QCXWZO6YKWk+czdTXsw4Xm6Xo8gBiDWIyNCoAMekcRRKBsrG4AEUXDr
ZxkIZkMIZqj5vb4Bey4mLBKGV3tkLgeT1FQPH29m3/ULzv6DHr+mfsROWvM7fGz4apEtUTdWlqEe
boO+wZwlumtno/D9Ta2szCpXzFaJMgWExShQw/oPMWxUo8ZLeQcBOra1uJsjD2GFyo3fw3dCoYva
3XvKagOhckyDFNTfj/IC7faUWtKtQM4mHDkBss5/5MmKsfapw74UrKglkqmIKQ7ScEMgzE4o/sYB
9XdKGNTFSrB2xht+NbDbBA+nFIQWKlVSZY4Wx7D58vDbsU5EzKRNEW6qp07Ubv+XlMw6tSVnoHZ2
ZlZuhbNuig1J5V5YyJ2PyBJXa/A6+JkHlz7ofWt0Ic1aaYS9g7EeQUJpEUpBVM1D8TzgtjEYx7x+
N2XPadS/YRkZwQN5Q9O3nrh1ofWpJsOnPXD4Bu3OujS56LupgBu4taUQobU1af42jQpQSTpn9aU8
v+fODg3C3BPiRfByTn0Fj6cIBRhsXl20phGbSgN3+qWKhhPKF4TcIfis+4pWXAaUHk4O3t8P0Dhk
3JAVH6+fSHymXMq4QJUiVhhoE5ftgwLA0QQjcFGIgYbx8MrrZCaIrPeQWeoom1OZ1lsUfdoXXsvz
J8vKN5Wj3giQW6inE2LSP6YhbOgvdBDSN613mNbZqwP6TqMhDFCWdHTs0QrANIDgMPjYb4RUj8Kf
ml9z5v7bMdJ330Y+tcqcYS9lGOQUw5mLu/zBpN0kh7q0e9/EhxB2ypyFRUteDnb4IClahFXSLkf8
7pRXdRPuiSd9eo8riCvrdIy/x73HK17dkwaDc2NxasudFZSQua9FN7Q7+3ATwqAvCsZ8IKqLFRF5
vEneFQJ72bCzgSLkcmMuA7L5Fh3qj9hl6RjMy6NPUuYPj/LaqTo2lXJRektJ9vKfBI0cLZc9w3Ns
SU+U2uhwq4rsPUL7J3RvIW8e/7GYVOisFrCKiurCDhkzadC3t6J+dcS46LDq6s0DoOgQrpSCLqnY
5WU26D9i8vmfxaMwjA79pIqIvUONr+yHTnDupyny08uNkwEf/jv6U5o/ERJAKqQGcdlmODdHgcxD
G2nRel5K9ilnpWTC3ZVAQ1t5tQ4Kb7F2+PJImhPtQhzW1QXw5MRGhnckxsOdMfh/IuRw2AKWS5wO
MtxggBSCcwIbpZmFThCCN6lMHebFOfoJZLAbx9XJjJ+uUaUzETULvrLrKwBiKR6ubpH2dipCMtiX
/Gu9XIpPOZR6bW+J1fgR72mXWBduKIyz3xCAmBAbZOcV6//Xdm/paFd8G4N3nRNNxG+Sqt/gxNMw
hF1lYATBKta4eyxuwsLs08AE+gTfSVVUFfow/VWS48/9021TvzAStX5hhx48WSJu9aTqW+eC/FZS
KOpJtf0JpLJ9H1sAERuotaCpTGfU928vhsWUiO1joE6J6i4cO3U9VbWdvZX0Xp9rStm5o/7vuJXQ
NOUk2PhyMrFuQP9w5QejnUOUY6cuthmz7hkLw6RrEnOrjJMJ4IYToLNDRJ6c9WB1alF/4vtrjB66
tkwbJthKedpZEvSHC3Ek63jcHBKvWxrDnWhunMgkYZHRRwTwcMLHrHdFHOTN5LrDO3wluILxvbLg
li3NovlywJ/+By0nRxSh7m+L4VGUB4bACEUodzeYk6xAL09y6+V3t8W+0m1rHP+JKqTUmv8YLbrZ
mY6678V3CJBNhQupBDF7m5AawOfxTWejDaLX/plItjooFTGdRoO2F5vkeTtKiNZUODIa0liHwtgC
SdnkJwo4prs0kOdg509CV8y8ertbfabHd4LJ/5hQUiy5zzX1usB5PsJEg9G5QXW42NfC4R8UwuZD
6No7Hq/tBA5OC7pGnJvoyM45eqt4R9YBbtwUzYqx+rEVKk6M9a0qn5eo7wSoJNBMHy3Qw/5SahZd
OGwV3WFDYZZn8Cakw8vPEUz9mi95zJqbT7JdH+8lBsFKkxDTgyWzroL9OjAtapItZoVSry7Ct7WK
pqaUMd9+LmwxmpOmn5YJwJBjKcG+xSm6jZ3kPJcAZK3K25VJWLqvSpeUnCiMUSOPDYpUc9upQnyq
a3Txp6+saoX28q/sNg+IllLGaGrOpoNHehQZ5lwJQC+Z+oht591iK5jgnhWM2IIS3jj3a3vIwuBH
2s8laQ2DGtfwMRJ/KtLVpD/5FdkaAALd5ubolFQ7GWrFQmyemYQ2vW9qacFLY/G/qlNl9BFvxih3
Z6wRudsWIP4+BgDLYj8F2T9ub+2Tw/XdGLn56CzG5mjBJ49bV09QEMuaF4rl7E6hMbmnJkyNDsPJ
w5NY1GbMSfnx/HAVvYo1S5XhISsUXyXa3dy53KOWKyYfsbQzPvDQfg+m7gKq5Qk5XxEJlJ0VpzK6
xCCN2SIdpeY7Ei0pnWsn7o1aJdcRlgELpQUlh3ccdqMmn4SYxcxIK/rpJwHLWTsokHhIvKKeAAI7
YWD2GLzpnX1eb3OWoWgMbdpSiUwdAizAvY3oXzc2pqHIa0/s6IcKyrwwtgjXMrTaBlwNSpCVkBSU
ch6Rh734m0RdxA0gU+e71qDTJEbdVXKNFQOXPYdxFFHb4RQV+Kk9eyvVU6JvX9SqBHnRce0JXpLB
1BwNuK3IZLKWsPQ0DsH4klKE8xZsB2s7ADFH0Fmqf/nHRzjnZhubZXIEfQUFEw3iaJaJOMzYUomR
XHDIpmva6zXm4+mM8nD/+O2EyWlWXz7g5eochVfsVXTJR5jssigV6vrKICDwIgF42r/52sTseM01
YOQzGvCp6bk5cidKHOl3kcPLRGoxuCvuXIBkHksJpZuyAVVqwYXlRMCbBXVmO70xVtlGoVCzW1LC
2tJeDrL8DpLqQZqA/jtW+bYrLmu8xRGDPe6tn1mjlK2vC/OOZ6xiImePt5RtUs1WYDtmvK/y4zq9
MPcabwZMTmsyM9P2EvZh70fmlAhCxbhCBBaUIndH+iSSgs4V2+ACnM1r8CTQypa1ME1A/bS7Cm7T
tH4aj9Gf8H0tuyG1ETvVFlc0K3h3eK8lAyukBvzyLR6+MUqFVRtWZtucBU6UCHuSaN4m+MjKiJjg
RRFhU8u+i6bbVuVRFMSxX/wpIQ1dUnc4Em3XZlhVCvO1G0fVBXuOVoCSlEQb0lv8VyXP3qQZ0KUa
rNmAxReFjDDnwiw+Ab28kRefHlBP3D8qgmqpgfc7I5OsOhY/38IoA8PuBxRwssJBmVfrRR6Nt3fy
P9vNZt1zPG9xvm3kKRh8KJb9KQMP4refggrjY+4Q7UPAl+qhgDxKJFnmy9Wsu+SBrGW0UzbwXTXq
u9f31PUox47Y8Ysyvtq8wsYpHcXehD+z5RfcL9LviInbvPLLQ5EzK33RGyM9FqccwFOAruBV9Ide
xmS6x1dGLHxIV2xxF51mZPQcS/Qk9UgTPzRR14NJ5sf42UI5FVR1FWA4j8vhIJOtnhYQwOp8Y9Hs
y5gf5CzvmbOGL+0CbSjFWUvkiMYUItfH3Rk655uWg0xlS8YvgUVKkxEOYlOG250HBXbLJfVcY8YN
O1kXJbJ96kL3QKdLi9VndO6nNWvykxSLRaP4nNWEIQz0uJ7CakbB+90oXu0QYzgruhDyMuQ979Go
kwWs8gArBiv3I3L26ZgSN8r2sZr57D8sfMG9Is63bF0N4+MrG/PwnipvNVzKbNazdg47D4Y8hdiN
26UP3sxILlPZGC36nxsKSXHSNxUQgafbIQwei9txs9iaHzuAdy966lpXor4jyQfpPWm8aYozkYhy
xLDbGJi3KEOnW7NXh+dphotjqbRQE6irU2OXneOewORrrPY6bb1kmV8DIQczQVaT+17uV74avCDi
+32nQ+t9jr77ajbsInNUmKpzIUsGfQpaZM55QIAPtrpnJroeHyrOlb7Vt03CQRDcY/x3CTYQHbR/
wtW1CcGJz+Ht72dq6/skPK+3OiBTKWGc86Guz6vD5q0BtWe7za1f4g2pZDEO1NUDtkdWqLGn7cHD
EKUIQNIVZ+J9jcqBYroaRIidePXu4TvKVweiwyMBcaxjPe1eYgiU8tkWarjOhIL9+8VcM21s7ZzO
0yiTOzv13Iga5iDHMY57AmZKBdJcEFxVxIzppUg75nrbxOCCnkHYVg/m+6jo7KEU26qjhVBq56dJ
MtiIczTWpuNgqzA6N3VgoBAn2lNEo2i0djJcmTM/3SqgF8tlY2mgksepFShZ0H5PIfPDWcZekXOD
mvT+x64WIdrHjVFwZF31wnFDhMry3HHbofK3+nwjbcU3BCIRqycd9vCClr2PAIe2CJKN74uPVL90
U6imgy8e5JwsZV0rP4OTN3rOM2qMq/G0qWAyY/VoA2XQQeligt3jDatacwEkq1Rjv7EMrUM+Yv4m
KI7RbKVQ/4SIsJ/i+57ohUTw/DljL75a8UAkiDvfqA3MiOeE7PkZcL7XNBhHFN8brfcFyvydZDHE
tY8Y1bElBwBFWz7Eg/joXY43u2zNezIDhGfKhV0PJySfCLH8Tpr70Lzk95wZMTjwlR0h1NA9gIlx
Wbf0a8lu8Ij5pEWOJTqe8nVSEjqG7Mfy95xWhEzaUHrdJtu1UpHY35zGhCJXqZHHsYn+NALlXgoH
TUT2qWP6OA4B3EoLO7FBaAFGfV3JizUMFKHCEiDoWETj1W+pPNZvFK4VMQDbE5meN5cDDjecBFIz
PvZGn5tdOJ0i1GpYfZDMIpxyRtjuvP8uDn5SpjqEHIQbl9G1CgRX2tyiigDVBIagpZo46Ka0zE9B
AifgnJ84QaAqxvjsmQH1/sg6bZes0pCx4fPlmVwC5MDunC9GLa4wjcH018ux9qWSI+kD75hagS0h
f8MxyqriGfMr6DeGjwdfJzruHUTV7Q6prmyLBy5K/Oxyn83QP5PlSOYmH8w+J58btdNcARquXbWN
ftxcoq+EcQ6hVbIHwicvi5xWWklhVs1duwyFLMkOlawN8fuKgyb/7rnSMnuYBbd3vKk/xE125QGi
O0THxh/xuAuCWDZ6eNbNJthJM+OCatTGwpj4LF/w5Mly3FIyU1YAIB7a+cvHw0vETExcOUZiROZA
mWE5YkdsSbitubhAS/Z9J3TyZDaoHnvXaIhL0bR3WMHiMHLG2Iui8QrPxpxRIOuhXCxno64km13M
xengChK2ArXhGugomADV9AeCagP9oEyLb1Ia6PRNBiBYszihLtqRInx867N31mxITIUfaB7tthhG
DXrbPee67DHJwacHJU+mCj0CYt3SQiKwjsNV/+xzlneA/jSlBBIVcyRA9bf/3FqKgs/qebKJq+/5
/01l0LvspXF50xyccx8O7/qL5xJ5JTXpqRH5BIFXpsjzDWilHGfz0TJ2GDNieB7cTeG8XSd3bqnP
l23n2r1MN9k/CrOtH4BcpBsPcA1/ARhmZTWJLDgWcpqeJEBf0dpDcImmPmNM8Np04il6Yqthj6Zg
Mg2brp5alPrYrjVkFSoaOmaZrRiNfS9fRykkwLai4wNjTSVylITnbLorWyWdjvT/FHh0O/e+02kV
qkGwNrFajBGgL42Zc08XwfzZXbaZ3QM3SdpLjJChIbTihz8ebfzOyt4IytEA3XhodS+0bkHvGXGP
LJzE1jqD63cg2lFdXEbp+sYXn2+LcELqWW2kSZmaU17hqBbfk4qmRhcsBMMZ8/gSxNcvc4abjr/m
Z8KOUVCLpBwVIApxezyIm5FuCkTwoCx1IY6cGZu9U1D3JwDX4uphH7H/KGd4pnlqYifUsgUwOG40
hCZyUNNtE3d1QogP/pnSG/ciD4cgbu4pMDeAZeL03+T+Fm9FYZRaq17OPpWzeBTakySrjAz9Om0o
PCx9UBD3L158TkAjwDijArR0roNOCUfvkKjXIt57atNd+UGBH+XoNx3puCoWq6pHq2JVxWVOrjiL
aK8LxNC6Mlhb6mfO3TEnYUdgMXQqhr0Tl3Au4GSEaDEhOchv+04lwF4sfLUvUxQQhWkAvvvosnGL
nPVikKjM4Af0Oi+Xgxcu7EHOLHhXvgJJRKeiOeGuw5Os3ryqFk5nn107MTNAMpSe6iG2RgBmuvKp
f+qfZiQ4DHbrw1D325YrdKUZFnEStSnVaH6ge1EkbYKYddc+Vhevuxe9F0wkLu6RJvbD8mjZJzUD
vxMh2HvmOJ4i+lNyobJxG8hVdO7d2WpEtvpZh3rBNtZ7TgK5y3RgI220YMBcPkVTWn1K52xs5Ym7
Acfx/PDqJuE7ptgESFqBhuUZMHwhWqlzlXMdkFZCoabnRugKvyEexsUcAFDOdsATmF2B04oaV9lT
qO4q875dF8jiI0/jJt2KvKGIvB/0beGsMf/hHjskfcVzGNv3ubIvt31eskB/CUcst3q+i+z2uRku
UGSNfPANf7bE564xL8bIvbN/tsMkIau5gpJdEXSlECbSEM7z8Rjgk9FAP/wbk2ppbiUgnUwwgFOV
y3sFvRKxV14csbbp3bB/ORWkA+uMwN+9pe7o5YsHCaSJab6E2ntmo8crNPt+r551YxBH67YfXZ6y
NoP+svX6/QYq48yhrRzfwWO2eWohhXlXMufOWJcC521o9a/Bq4i48wC+KNR2yuxW1YfkcNur4gcl
19fq3W1h6M+BLfND7Fq8Wxg8ML585Kc2KY2Eo0oBDh+cfmB2fTTwT93kBvo2uN7E4SwpZZzYTjJ4
4T6528ChDLOPmYK1h1Qlu6bUeqLs6GKuKkScy9LTRvVhAcwNpTFDhY8XCgLW4EHAIQnwhVJk1MWb
+e9F10AG5BZKQbWRzM55DdA7ba5pleqbWU/QGGK6rXgkrAKKoPPKNx3r4rt/YohOU5DAR6yn69gL
v53cHpg2kx/gfCuV8+cfJI7ZhyzhAJn4vIGNgkj0TlEmO48NwXE0/zN9vmPdpKx0zuH/uoyberQ9
ZRvJmW3ul++/bW+bItRa3zzmAEDve+vwE1JYAWIpD6zLk9HmO4V6balPQV3PIAqjKpZeuDoAL8Sn
da/UJ6hfNUbo/e0zkConBwcpK9RMKdOaXiU7zIDRAdaGZ74Px0DdCXrAmv2Hajux5sunOr0tGXEJ
zGf4xgOFTeyJ9xJrguSAlPolOAKyVO2xTAz43T0VxTqQdjpKAp1i+D54pUZBQRsBTvrxj7p2/p+Z
upHc/IM73LMFh8MyMVsfdXTZ2d2DxVicuEbSJY8LQSDFueG1RGAx6YMkYrmJvy3fGcCNcbh4T5QM
j61plcpSA0Icrev4wc2hX67BZ6BQl5Zv0amGYT8qzfBayYPwOHnE4j22y/dKqlxv5OPD8B0SDH+Q
COca7lmCLg8nXoPGq+RWoCLz/pCEoWaAoo4ZoE+aAECmfGHRDa2OcuqI7Xet3WQ8MTTyWhOQ06/7
wgtM6+RaO1nGtj+ev7iI54bOxFn0FwxFPScndKzBuO0DE/9IklBqRdXqCrGgrO21l6EWeylYo0Z2
L5qUsFRwATZq9AXkJClSspxJ3xBzWaQFOcVjlTltGvzvWNEWyp3nzvbP9klBRLHpBQ/UhghIGJvH
v2cIkxvCd601q7Zx7jqpezT4grMk4ATnFIZuD1AeEYQByhDZo6pDXiR+Pjy2tG3tnD9THXMtPdzh
oAl1wFaExjITJe/+yzLdaP7mg74Wj3eQzJ0IrXIX36FgUnk2wRXg1Tc5X3Bw6+Fase5AZmELiOwS
FsdFSZ+6flpStAjCkkM3OD89ZH4LDp2nhEo4+0DAbqhqEnyg1K8vNnD5iy/jgZpDaF1PT32dUKI2
2+hBlzdgzPlvkeKCEpgIfdop7ILkB9Y14Nwye6sSWWkTyr5uAapLlvm4bI5eYbDEhv2BfEVexfCf
eJKlnSL3oA4m4scF6echqyrZs2VQjBi0d7xxD1fyYcfIAz2uM9LZxRrW7DfiJ1vL88PpW0tx6zNa
4FSaf8Lz2g6yPnVIcqzzmYSq+Fsy0xEYOI/pQQxFiTJlR39/16XVLXObmMPHpOgLd/oczhfbVHuj
xKJtHtfI0vOPlKCyhwqQAiEe00T998Cgz/y1Mb1TITqplZ9WK4+qfQSsY4yiGaP3RdPHnyZ0ZceN
s+CZwcvyNPLypqKd08XwajLWlpZkU4Znf3hw6CDSukiIHShUbcOOaRbBLnd+hjA5TcDHrnqb4h9B
tKg4l/m0E4/FM8U2QTGoEeYKarj8cih5ZmOgKnuAU0cYodpsXftbBHeLfywu1r3ezjNWBC4dcigh
CqA1XMbZqZuD6fO7T+j9OXYpAyMntvdvFTGw99IYOAIqxkMyrpEGwQsn7BxYJuUU4Z8ikPEk+ERw
42gvjeGQj8urbYAaHkKO2c9W9Tfjb0fuyu2H3wV8s3CIE7aleqBKbs920m+vbLHwwVMxLW/LlBmr
QBkU6/Tyx0u1IzuxdCRD9SFDXmMzqBOn/TiKND2jF3udhrm37y9BNG205exn1H9D+cIjxn2Kxe9M
Zr39zysRBrURDuOneIqBk6ErKSYDskRQ3aCgss82YZ1IHVwP+zLRkNuVSAkvcqPKodof8U2H1gVJ
aSVMhBask6Oj18Tu9o3ZmZJe+Cah+7jDYhfCHu9QLMJjkc3fuwt8R/Fq0k7KsIMxBcsd8jOSl3W9
p9O4ZWlwAoAWv7X/WJbwu4cQF2w+MkVGOfaYT74C7r7GHxm+6AeTeGlyanqAqdHjjLuyRlSxARC/
Lixee5N+3Ge3BcYoCWrjdmrEjUChQwmNLAwYxL23HR8COA4jzYHqIoSN+cfsi2qGUa3GbCV982Yv
rsPNHM+QAY93i3HpnGTyHy0XEC/PYmn7Ql6hoCGU3288o0YZFcKrPnYlKLzTSYoouN8vwTdP6XN7
XowRiv7SuBFIwnsrEMGVA4t6Q69lI59JsVLeQ4Sjtqytr79hyWsI8ysyOKHfiOR4yBOdgV10KfT2
vAf6tnQdZCPG78KGv1RA3Ro2NYBvp96fYzIV+YsxtF6q5F0TaZ8c3dL1sgr4SJoVB6qx83pNwQqO
SSilCTiZGRNCYGPsxfq84VWRT390Lu8QPq3+z+qYxqqd9i+PyKwAbdFQtpXBT4CNWkaXKYpBvxAZ
3Kbz8PmuRi3h/aECUnKXUbTYUNBYrkMgnfnK4IDshLSq5rupzYnreoALcwGNW4/8TsxrxKSqcqBn
EXj/UJF0hPZ4iP2Wmc8k66QJivNcUS2aM2hoF3A+vi6H+Wjp0/Snnhwfi5I9zDHdxaTqSiP07JSk
grSMlCGPvRa1BJ0LSfzlhNB7UCZxcvVJLf7AYKUP3zC0+MZ3Ec5aQI7zXHia8zemJiM0dLRyGjEd
VOE51Ar+yPS0U69AfZisT9Xc8SJaFcKNCb34rFhdscScT2VeuSp6PMmUNkcThUvNjWODxB2Oceoh
k6Cp87wwr5bwr3/bQtpdzLFvpHYxLjs6W4ST52fTQ0iXWXvHSEqDwjtom/0pmFahoDftW0r4+oYp
hpFInHx4vh5etm+Dj6+4sZwITXh4a2JLTP0bQ1fjf8I+p5jsObYrltTbfnJld8CarP/0u4Rca5Ok
IWgPGAZR6XHRm3sQkZ/rGLwcz+wcwsADL+7MENk3hiBtGHvm9JTXQHAUY1X+BF7w22RvJSYeOwiN
RjOE00ztCN0+tzNd4iITVCZrdrC5xpiTWcprYlBIPCzc3FfEJBRIjpihxaBVyd3nYQ2hQZ0gre8h
B1UowPmWGoLlqi/09Nq3Qp/1ipfdUoCtXWSnUhq4QzUnoB/4+06QGhsJYKH8h5hI9leHvBxV97xh
spUpnOYmWtC5imAr2a7iMYnWJVY/jOxR0zGxS3QOrit0Df9JUZN+catq7UgJsTvcaflvKgmtcI+R
If8NLDAUhuYAYsHDIQwHLyNq8u9Jw8qKmgzowD/P+xTgrFevk0PGxVCfvWJ9g4pJpFidGc8zM+2Q
4iwbjzb6IS93iSpXclDmkEReERVq1kfqK0k73nEH38gCRjghU1EhU0z8YuX3zz9QEenGwELdHwfB
dbXuYWSWfn6koXnb1lkZwqf2Aq7MXTNldzgMU4h+ro04WSLWn1m4J8XgzNfQ79MH02L6eo8KAtf3
tPCJmxx3YRoia8P4jA6yELDu1KYSeexiMMufM9HcE4AT/etSqrsJxoz8YKrE4KJoQO5+ZmGlcmy/
j/vare/d/+6w4vxb8tuaImWiksbghL3NfKHlR4afyl5hc87PQ96leImr6CG96chRWLEp52Ebf3u/
30viNwzOJ+yr8Fra2ow2iU3Ki7cRycw19pHQ4FDT1dFntqpP3RWlG6+W9APZ5+IMurF5VHUuWPI+
eXSJAeLGSOyj/Zy39VVsZcSvarWT6YGe6ZcKBeNtOZGbAlqYrfmBU/jEtaYsXPgSmX0TuDmMe3CS
Y4C3nFAmuvq0QdDAkzRSn5sM42PXVnluLVFmnbcFZyRMA05+PlWpl8l+9pAMCX6U/oITg7OO+lSm
Dax1mZ4QXJmgOZblycI9H2yW257EFneT4WYrOllp24NbEZLtfVHPuWaR3tDI8kN4fBncKhoeTo87
8AXfmyUbjpbjYASfSnI5fl9MkbmBQvRxS7P70O70qihWaNZvzamEcCWDiZsSc7yZnsdneEmNIKig
04mUFTCV8q5DKZ+ClNgCEYJ15j+qw40lRie4zETo8DQjzzCgy25w5nHC8kuxVGstlaPFCSCLH35t
PiqZYk4RD1WH0cfB2ZRstq8gAadaOe6VLod6sH8SqHxjLzWQtdy5gK3v5oSXGsDlIkfxebaf8MMe
rjH1TyQnmjdsMqrPnQKqp6TK3uq2F8PjG/MP1mNjOWp6XdIL5kAk8RFGX6BsqLdxFJtFWleHQsGC
TD7f+hs4Lsx5ErHomQBc7TM4bJbIHJ/0UBJmnlIT6ERoF9U4ld1HMR3fJu3LU3OlVtVPt4Lg40hw
KI/T/9MRpHIZ4+R7VDvU12OVu94ur1vqDQVUP9yaLds76qzfmrWrmi02c5F1UG0GZqaEvMRFIKRT
rbb84sIVN1VfO0yKcFjR5I1wIGgue1h+vy0R7dmUg2GwW//KKi0yiyIvBLolpNFItLYxYtUq2qSU
7qprvuuJca3/7O4zH8yAtuMprr1odk44Gqr9V4eoqfRKaNV9p5ocGtVlmC0RMnsX0AsFz4hIOvAk
Tdicq8XPFY27UagnhJfHCW0psVFtwoNkiHe9wkmtg3GR1VXUj90gmycfh3UVO5qmuZ82qnklCpTY
LdhqFjgJzk/Da7Yw/hmzYFLJr99ouwuTGDLgjzuTDY1AiuKik5VrzTxxmEhFIQGUPeol4gMW/wN2
VUpv62dOSvZ5b5eWi8rb+28oaVnRQnk6Oi8O5iLgM6JPmyGcNCLXUX9WJ6rt56xsrlamgTnxMOkt
x4JeF3VvcubtduIWzQ5w2WtXdJAsx8VyZSZuzR/lbBf2trzPv38h9mjiwIxE53Mw9mHO5oYT0CZM
J2fScOD74lZc+JratEpHPgLF5pLxCK/TVo0v/D+7gF3IMQyHbGxuyKDTJhBOtaa/Fkb3QZPCUlFe
8ncHToTqpy9OzsBQ0pzUsQdtJ7VigTFRWJzae8EDrqK0ZnzYhnngJJy8rWNBzp/KQD9WYkEFLCmY
4Ey6immA9tKSEhKmuNV0SyzN66+lZJ9d4CWodgiKx7MAwatJSZ2c9q5sjRYRpT1lHpJQXwRFrvZC
cCPb6fB1VHrJROi+irJwzOjUgpcoU6pt2tnLEejsQi3/yCZGKwtaUMC4wM5Zty28PmsA/DvXRiAn
lQHG3gSmadI6PBWflJZV52zfCTyyIUBE8ADbnFYl2qfOCOZ4NEw7QLcZ2OdmiToj7fe1zr6dYHZ4
Dfh+3H2vSvsOJnSyWQvM3TdI1YQDfnL9eMjjBIBWIITQ+58wh6JyYXhuGu2nCb5GWgqeEbJbVd3g
WJAdMwpkiIylJNznzsMCnFGk55jT6BYsdN7mVvamW1feGllhwy4mQ8QAwkXQSsPaKLz58DoiAXto
GDln9h5q4/jcsXjVN0Cahc0+7m7ZqY8LwSDznDXByWGQnNxzXOI8ObssJyNVbGNDgPLP60Ag8Vzd
Stfhf0tG1OImOiiJnErcYvvhx2XiPtmuEYuFf+QyBTE4vejamWAyoZ+T7Cnkx8gIjnemFGnZ2Fjt
ntvuPNRhGq2ZKndGWAHkSe2Z8Ln5GJLZdB5dlejOt8MgLTZyVODpvS+BXa8On2gfrDMso9ZmnBol
DnGri0hCwE0lLbm1k1PqfZop5m+yPFNVMMTrp3+vDEaBlCYDPB+QZWg+lPfKt2hy1uek3NEXKvUZ
iZUOXRChJjYpWhSrIQui4AESGWb4aD2aPp6RQfPpdwEnwrrup9N1a22/Awixbugvf/QFsat5mP3a
37/UQ2lnFvXVXhlPg7XZ/GqpOzF3D7rR6bWAXKOrTbhwA+/RD0zQoiyrS7H0B1zPBNKCve0sHCut
PahJdESmu7AGesR5tb7WTPvfJ2AtKUCGsFIZAYsiL8FfsxPlHnwtwatW8yAKUkF0CkN0lu32iNro
/bRsIaNhhLn5IceLsuyy675zuifDicgkQB3AdesrgePOFHOgSs+8bXUWd6ybbikh2Z+hW8FjNu24
kf0/WmuYiCkdFlssgHkWsIdqt2YP58/z87XWu08ngF1rflnvUkA3UaOwpyz9p9oTlVyDP5sR/p0C
vbUPhBD7HrdJTIA9JOahgpANBmbNSpQsEDggkjyhmZj0BpJC5WP7aZH7VKQUUoBWEnoY+YkU8hKA
iVfRF8aANxq04M0OvyH/bTR3H2+W8W0oIwKLTqWTMmMxY5O++ShtnI1YJY8MT0vj3fod1j7UT5yL
puBPEuNA9SnZpzBJ5ZBbErzMxZ4AmbDVWiYzSOEmJXEL35d8FdSk+juZHjmRaLwDqIyoJSAwN+cA
4WQwB0gmoPQErRcwJmaXw8C1eRod/ZZXmnrqMYHS5hy8iSlwSt4i1qDBQoMUXILXIEtlfAMm/+eE
TVdzPKhP0/kHa1m7H/gD3blZbtFiht9UMHyU7+yMR6vb9W+soyYr8K5aG3SyhYeSWz9MkKQUUJIr
5gP6/DyvpHU+LkOnWFOvr5TFIjc6m07BqztTX0wuQlQ1sroHkKc0s9dA9gpPiDUV0VirUTmtC7g4
z31R9ppT0aD9zlBENqptmQz8JrcxrWLspI5RCQrYCAmOxjMRe3nChQvuG5hP2/8xQLOdMzjnMm2j
hrhv5BRDekh1HKF9KiwEga8EY8oSazRWdjOPu5L2hcKnvwyb+Zw12Isw6e5ADB831qXkJoeuNRTG
jTkqb4M7g5yweGjonvEWyYy7fsbv8C1IaEp12flW8hRNKr/oFb48wB1GvZBgxowVybFIUy3KcfZg
eErSC5Shi8Rnw+KH3tkLTVOMzX50KxM2vzko7v+njI+gOpBCe7f4Ert8FxKpo+20UutpmLvClqsc
5FAXGrrB9tMYFHT7z1D4Nz3PVz2T/w2mq5XoeNopBGf+34YaXieM3EFPEZQ4kJtojaJrHW4LPnGu
80GpzHY1Mwq33aVI4qCzCEE+KL4GjV6TN5O3nD+PLUuTmzGYspQhiIAvpOev7QRg2L0xHEpSPzuA
RAYwVK0vsQTI9qxGkxssU63E/UQsdanGCUEIEDNb/gdlLm+7C0wT6HzxNe5FURhL+7bhB1orBuvY
kbJSZCJcQqacSwPwoliASrAfF/XJZNaQ+yx52G8l38liai4Mp+KoyviR+QWlcoDUJTZZ7EVof8om
K1Xif4uHWom0KHz3a8kHC1jgP6jpyxyx072ONBNCAJV6/1KzvjS+8EcjJbbCq2kmNrJlM+JrdF7/
1k8F1Z0+dof86HvvT6tUCJ20cm/jyW0eGvCuCckMBL3C+b1L+r2VolA6ikbW0kUG5rozn2eYq9ZJ
vOCsi6VeLxge7JgcpjDOk2tBM9KlJ2DbJ/Jw5seFRzRPwZ6snFfw9YZuiSOn6qzecvFlLZQYxgcx
w5yFeSuHpSePMZXgs2oPPHV0MN+0XJvY31xhesmED+Qa95wNDuLxPIvNuQBPgmaLHBfbRkfiQb5O
kxN48BnytWtmr4/Qns+x+zM1KPXO0eVz6+gEPsUcYGlhdf5ufVJCWKlx4ZsHY9nWFQBK6p02N4HU
Dts9arLOM9RBPZsn6i3ujJvGVyqfqaTL1d3wQwX6RX2MWi3OvIjaST/lu9rA4SYwup2wu9r5OCZA
LrRGJF4u9tl/cps4B3NgpQiyEDOm/fwYSdemwJDePyTy99oWvneDCcZylzZU2gs1v2KR81tftA5n
TJZUVC3X6IfSzZVUZ1Lvt0Jtco/R7xGO7Vz7XWBGTd1noNgS/+QKh6eEfKNlhL6I7y9T/gBPliMt
/deikZwpDr5hVaMZBztaTVl7Hkvuh+xidTGSv1CczWRfhgaSwOBE2an3v7Ge+c5tZImVfLvQlBCG
mpxxTVKZQ/exgPn/kJ/KhNBRfADSAzCjssvJBME439mNRWP4Hlmq1bBPI0lucEMvSFXb8mU4xIVI
oW/P5awsvaxo6VzLoqwxtdSy7gEFovX4RS9Ohmdo2UmGxg0qcd7LFYLyeLPixM89RhVgEK/cMocs
O1NfGWwLhtU4vlufHyH8MyIYGr8rqJ3xMQgDxNGVbNULV6TGthRnhYkOxHTC4vlih86GWmqwBrb8
5p5BvXdh7gb7+vJ26YZYjBBfttmQnDTAmW/v5+AJAcUEgX9gH5DwpaKzpfRpluxIrFcqNAyVDpgm
kRODVIHVZk64RgwgZ9Dg8wLNiv+PFvLXXrUoVDhtN/nfOf0Y7VkY/jFwktnzv/Pq055WlEBIHQej
pEwnKbOfm/NqnSlH2Hy4moJpmZnFTgH8LXE9Of8gNhzxu7RtqJto0xdKd/Sdj6v5JVDGR7h9HBMJ
Z1GRKB8oKrgoYl6ufKfik+tNwHqMaSx4PpZm5K1YHvNke2hMue3aNn0UCLVpJzoG/wtGkgKUcQ/G
q9hUhMU4dJU89Afl6DdEUEsO0VY5ZMemvN71yfTdsNKuXvzifoE+qpvoUNK8xnrGwIAU6y1L9FMZ
+PD/O8CuSnkuG452l/a8KhGBuM+Hl3IBD7Hg2WW94UgyoG3jYzHcYeBCy+qgqVAeR+L+z8gTKU9I
7aI6aIbjQfnaKe2q44v0Z/rEQW2JNbdL/JHVsXY5BLbhglM8ISFT5FKOmCVHGLBPsExaH72BAGmg
1HVnaFDRsqiWxFPXrTK1bUD7PhGnZACqQDP74pmtFm59xk2jRYShnwFdOYxiO/AbEWOuzp6kGJ6v
7VBDgCNdwhUg1CtsiDZLv/Gfu6JE6YpiUCwUCaFBBfndWO4sA2QECaXLGI8uRRjZcn8TIfafy/zG
JlEaalXL9//wHI75+bY+HAzRwMgQNxrPcCKPj21p5g9IF4/NKYocv3ML0Pn1wcktgraDeV9Sxj5L
nTJT8EVh8pKB4oFyUga7KuHLWntesjeFyZ94Qtf6cBdZ0TAir21bYuTsFzdH+gMmfpMcuQZoPM/T
YHKNsp+E9CQRZUkqpQMYBW45rFZtZFeOnrD16zWE3eBi9JWeXGFRX3Ffl93Shl5ScXVsf9Uhs0cw
npaUJjcChgQaQ17Bkmao0Y3iRJyP3J/C+yX2WIW1DFyQZJthZJCg3mfYio18lVqsoJDL+giX8paO
U4HsM0a+m+mt6uRE/eyOkPMc4iSfjM1bzsMGCS2IRtlsrRWpah5OGqH+PtfrS+KXbTKZvxrYfzC8
OzrqpigEXi7dEOxpW+MjHgoOtuv2n4MilowbO3boBSGR1kXBkvzygnyo3wBjf1hLBbeZ2pb7d33W
tHZSPAdjL0KTnadDPfr00KjkjFIa4iWDv+TLSY50yO5t3LFrhVUGDt+i2qWgLxUL+4HcnEtg02g1
mmMdEeRM3x3mu9DDZBaWKAVh3a1q6X+u3qK4w3+hRrtZErktR/SetJMLzeZpoEjHuAb7pmxngNbH
ITOu3QdY2lpUwBfttyKDX+ypArZGXkU0LO2+lKjI2j1vhqtXoJwbHZK4cIc6hmaRz3XMimM9AQ2P
1sf0ilFOpjcG/n/Qb37PFfMTvvf/rTv/pn2QbWyMUjcxRsp8mmCPs6YdmClCc9bSYGhsQXUGX5Is
GJDU7LabbcBpWwLSsz3zp6YgfRib6dwrRVTr+YsxlO+N9UFfIovuDvNgd4C6PlL7z3ieidLdMgYh
cGSDAnL3Xg3UlOnnPFhEo99+spj6ja7mbyZDP0uYm7pMT2Y0Ebk1ADcsO5vPE7NyoNP8xR+F3ZEV
J1j137T/54bCpbTFtKDUdYM/0cCY9dNyLjKYMjUoe8+EF6Ad7ZyINCcXPT4gV8xGGLkMG31ti3Ld
I8XJhkO0gBedBNB84Nz9utgiconTULg5RxqGoEjYaZ393i7HaaykewTEe8GuqxG23vmbsPxELrLt
FIIPKZdVrlV9I54Oeo1m522/5LaD7I0hWuvHPREkPhdaeGmacCFRTGIfkclKpFhtB0f8oApKs6VP
M5c8TYNTSGLJMRu/1RTM4/9/LBDTmx0HbpqzS5G2h9vc9s9c8Syfm3CM25TnEyzkj/Fzg4kQM1fy
640CgUDhnsGE2eaLc4khZ5PZubCpwSOTFWvfe6Ob5sHOULUrfQJMHto1IKTH6EmOi7ZjS14SGpFI
HpBArz3JQqopKhfZZeC4FR3myjS5WCZFmAOTivXPfOjc7oxQ5nfsWzjRMPoM9ho5nKB11E2hL71U
2eX1kz0VZsFOL9WBijHFu5nxdH6lYtLdvJyM2ajmUqmEoFAan+ca4fg5gg6Mne4Cac35bX6voqMK
l9Hl51Qa16xGaBCURJaVJkoJ/KDQY1SV8kwhA9kDi3d13iJslZf+Lglg/yEN0CQoXOMsFXgacZzz
R5NwavSndACba/6G/AFl8TiOpsvnBlPKfm0iYfJE2ZC6qaN+KSv1Z01T48DgeovrA0gIgX3z3ULk
/tIP44RPvE1cJ0KhByNwUADSLFFHSdY1BmG9QtZ1kUlXbAkW8WbrrTjXEZuOhASo6gP496W73GMK
9Pjoa8R9XQAIig6yS8DL8kMal00mhLo2At2TmyPyW1pHEvJBTqC4W5Uikna0AluPFlsLE/iBoOBs
RoTwFV9AKu68OfagZWVjieu2ckSiX+KQZfN+O9ZeO9ZX0etSEiLGC4ciF8dL6PRrEPFT/tyzJRyy
EdkJra2zxB66J3y97Btgmhcn8pz7CB55SFMcbV2QzdJ9+kEZngcNPeDXxrtrw3N0Cxzq8nTgHZQx
Qpe+zs7UenRexcJaBOrjS4JvuHpNENXLlzX4tHrgnGG9ZoxojOb+lTRe95VjQQ+M6ArXJzJyP9uw
tmWsipvsujdFrEi309DAVlwUzTJowBvQf9wsar6Io7gwASR43Ygk5tNXmUgvQFFCl0VmaljqyUg1
3nMncWk9PCnLBzb+g4J3fNSZF3vUHmhcsZIwd2SnV4wuUoy25M1jSOzIW2D76bz/uSoTZgRu7ETY
U789miEDDQ5+l/I4kKhhi2DwEKz/8javTH4EwPibCJVTZbBYeuWVpwcQ6ac9zHWmOoRJgeaWh3uO
THvsAyxVoNnbFl9IxTsSiIWrtn4mX4/Fqa3kqB82qG1esgtLkL/3ht0bpWO9k5byyaB3jc9qOWaL
bvXfDiSckrewusnKLQpeNjxBWSSSOggAnfMRexJV99t26SThEQpTMzvj3K1mGUn2/B5lOSwyLWaw
fMxHzabDQUPIAAgK+MMH+PzR22K1Lqts538Ca/4TvYGLZAkccqP95o2YT2zSb7BlLdDv2TsBhhRY
l3b/pKxzi2qiFnKNhKQrMu/zsX0I5SY18Fzjbk8JNZWEqvP5O/pCDABNKvqjDWJ/OaqOozp+sSRS
pDJ69oFx9YGEn+0m54kSzrzm6htm1aIvgcEr9MF5wm1b1Zek6ZtGUyC6fZyy4/r1+A+PJIeg/Qt6
EaZRt1B4r9Kr48kH+Uo2aZkX0uxJ1CayenxWVNymVZNIZBwiuM0duAjRJ04tJdBeSCZKkGogIqAd
Z+mOPHGWTfgZg2fgxgKmTd4gChxpQL4fiMDGcl5E2q38V8TDWWcjYBwb3rnq0M0QbimmGu/kZ4yW
8hB6hA4N4n9LnnA2Fx//U27IhJ0YXCnjZGfmYHeJkBtTDWAaYCl+SeSfjSkUY/RsMYmxosJSteyj
tUqe4iM/lgkZQmrOWi64AM+edGEGrsZ4uf7N/+htqVKpLs2RDJn/goq4yo6YtbDsXfW8aG2T5t9t
/L8UfgqQ+pFPv07fj4UXhdz3pSU0AgN1qprDLy8tQIt/3NKuW0U2Ey3jxfc3CHFe1UOUUTvjbQt+
OgK5nbxJ1Is09MeQVt+qbJz4Nzh+iXRDFWchfvzhzYRsHixoOehLHAR3OEnKob7SS9jcSB/j8IoV
//kmxlyCfCoka/8PqNL9LNSqPIFm6PlrAGoIVdcIOHvdvkNtHpvyYVS8BAipH8AcmgiKy8X8ogHm
RvN1Hgai+2JWuqodEVLtQPWjIN7visDlyvU50nKFF6RHMdbNPywzw3yHE85vfHDIRGAFlLyLRPC/
MtlZ8PR7p6oNBQJl45N07ulSpNH0IJlUFrPk483oWNUV5TW/d0gZo0rvsyB5O0/EODYgZxHakfyQ
+7XC19mZ+enw4A3kwZNpTKSHPJ2iT00V5l1HCeGqiXjBr+bfsRmTyUiaJVwfoYBJwkMxYeVUHzh9
O2IBk4vKkok38/5AI6BBJlOL8RGJcHh0USv79nMtlA5cE7PkdZ31Hl8DEGzvPi9u8z6DZz1fsL7m
5aamYcpLXYfMxc9xuQ5bDfFQIonPMkgypOVk8RTbz1O1r9csfmuKocCd6ry9x6tTYjRa2+xkkznT
zs6DW1pM4och1AZOfILdK1cvmkeej3xcwnXuzoLctcJSgrSUAiUpq9lZ4utIhXQpKZgtr9z/V7SX
rTqiWn3Xc9xznRVYKQboCovIZZuWIFO4CZFjmIyLE43t2vdwkp3LTxP10wljebZMwULfYWI8Cl7i
x4Qh1z1nsGggRBkqxyFnOvu+iYT91c4A1IfMMYP0oymFeAlNZneU4G3wjyte5FpHLQ0K+GaXHBOz
2aADqY1jkqGVIVPxAmPTrjrfBrUUvAumwAwDa/e3wWECPuEbmiPS9SsIDjFhoS16M1SoUYEPH6DN
+y+LPbcIvbYUdCzrdRALQh67ruLnWQ41OlZICtetJur55mDOczBQzU/PkFj1BVpqFGXUl6wce8J2
Pct1eujqtblHf4BgP7SJjcctsDbjW92D1pUPXVtzmChEabWmK43qWbUfUkWP0mbLOjtYBqDzWjfd
PabYbUWyFZTOhkMzZaR36WW3gBTp/7w0ujR3Z5iZ9+NqWPbGKo6fw41usHlc+WoYARFyBZhbKDDZ
NqAw2pcPsY5S5KWSoCJY/YsJT/fgYEVOz2csFNzOMBLnmrBvcZxLvjiCqhvAGPlW8O+KknSxC0zG
7DWgCrv1jmCHcYB4MMKiIZaICD/dRh2XsB1Ci4pr4lUmMWmW15CpMCLXt1/raO3YU4z5b34P/qDa
wBBknkz87PNLIQAHprCpE2+tZwArvbsebgWoVNIjD5jNrp2Tn/FAuTMPpdmCTqatTXxDEk6k+pV9
Ab5eRw5axR+t6pG5bp1ba6CUgzdPGFQzPM9+42t3g5GkHyOSuDlANedOgMiiTriBkcHxOyfdVUOV
eGKTVXXdEUzZrxK4J9jIf5l2Zu6yKNpEYaagPySm7/ctz4/lx2pgZ1KlX9Ev1+JEZcTitQ3XgI6w
a9RmFVWJ3TwHY42S+6+rcYUQuY9yy6mL6JMfrVm/10yJx9+wx3xNu0ZxW89SYS/PQTc3rAg5EQbV
4d2sCMllSuFV15p1zwjM65WBond/OkgXWU2PXtaR+bakFuI8GR81DJ6EjqZpYufL0Z09TSAInivk
5Nc5TWtO+xtgMKpignICSBTFBpRTvStZGld8GiVoMiZd5Jyd7lQqX8Ywpf1md1m28+Mt7fk519EH
zJ0Uuhtf7d1mppQL0poxhJegdzq963bWNhRO8AMtBIZvOExofswX9hRKRt/XhUlDX23FiUQ+GSK7
gD0Ex/EApQFhWmlxhenKISRTlrB5EkrrXCc3FZU+lMRZDferQtx3SwaHzjIG2cKC5siWmUfDCV/R
g9J5RqyDokj9pgBe9QCBNb9+HYm6FReKihx1oDKd79CM9wG6pRVI3H2F9zL6fsFPwW4oNIfddaVf
KRsrFxvlY0FEUnyZQd5T+4IQQ7GMwPImikN6u2rU6OFK+r9S3+mBOKeX0W18U+0GnMdrsSB6ERlb
GQqS19jliGKTnddXsdNXdYZDjLy4dtOR4Fcv69asV8rvr5nfhfeBlnfLncgjMDCsLLqwL+2UVrpy
37pspz9QWPJm3SpucrROZG4ZwmcVDGFpjBimAeGmRNj2wh48ce2iPujXd+ihBoQBmvmlUIgCtEM5
VAyL05qS1tqL+PqKd3n0Cr1FzNZiX0sNuRFQlrmC9w6bThcngtJiZqpXRG/MJpwIq89mcEpoAnnd
Y11DveccJrIKkPQwnnFPJayvbYdyojBUnAjSW8KdowEykw46uNgSfwNKJSLmlPP5inEujAEmrbSy
5stuU6f/ne+JZ1dEMLP8xf/NSnO+fhnCV24VLSq35iOHIe3RSvZexWcc54i3Y6570k6cqiKHedgW
OUFwRN8oIFSpBYtmd/MSX5PggZno90tdCsdIjJ0wNp267cxZ+EVQdFXeqeEMaoz293ls9IUiuI+u
kyv9k++8MvTjSzM2TbI1Zqow6V3xky7k0vkdC0od/hlFSpHhGf9dHGjy/IRt52+fcHhWHaTC+y3W
bZv+zQWBulzMt7LiNp02dsssFR4mVS4WHDGyW2Bd6/OWYfMd0R2opTvhKEguWiwDaYjL/M1vLbEr
oAwK1m2Kc5cInMaIgoGhb6FpiZ8xzAMjNp/IK9iB0PecLMRTUSej5oU1SZBpeDH6Nkug3lrlB428
X4SQVA4e99Yts6pMAsL4mFfxopFmybM4hY+Gs+Q/tPQHHQ1KALC2JylOEq8jKPY2yHmPM/sf4PST
3ZSfFbEHWiw1zQAkPT70HHPtHkDPe8gPJnfY+IXwnjEdR1cLKav+5jFXBPFN7zfmUwdtX0DQOZKv
zP06NWXg7LSxMREGYARqODUC3Gbt4XHu/mnvYBIgZfICmaepF305lsBNuuufu0xf/EZglDyVnYEn
B5eFDzcHWeFp723rRmGNQ1EbBMtg9rAE7BuUiY3/MXa0QGU4cb+YzulFRHg88su8Pbwla6Ww/lxj
3Yso3G1oMslwnOJXOCqkfpAAtoH+0Dt2Kg4bcu9zaGFCu+ZXNPjAajYycWa4T5LVxpM3V/Enjjzq
cdwhtI7mtf7gL7Jk/JblNUNyCFEk3wK5I/K24Xn0j1eDJMG5KzqXISA6qDhm1W8yVBrz+u2OVSfy
32UmK+oAt7vKyYv2pfZa9l9Bgm3MV3XIEdthJ19/YD0cPwn5Nz4JVMuL2UDTruVYkcqfYDP+dbUP
1C5Dxo9+npwmfDNO9JvDMWvKTwMG2VYJtEEIdSEv2dEwz9rV9AG6F2hKXywV0uLGzGTOa88WdgQv
RAQrCaT/Z5jvh34mn2l2oqoFP0+wAPvft8OJVxfkrOghwuSba+PaTfohWqbpWYC05yjRRHturKrg
9PtVItQUXckZzuv9V4ixPKgxJXTE3YvERNVu96dVfkd5J4Uk2M0a5Gj6QI/nmr2TbuP5BBJxMdh7
LiA6ZMW8M2y58Oo60K/r1uXmgQtJ0ydzZzrWLiVFQappL+CHXxsvL/8T8QabrW/ZBN23h6pNKZcO
OFwqVjmhF4eO1Vq+U8RcqpfjJna3tCBwQcz8iY8QQ0QXO33+V5XToPlwyiiY4h9rWUe77oQ4Wabm
Kre8sVd2XGq8gEAAdz4wQIiA6uKt7zeGV9ck0v2YgDR26SLRTtaL+JebwaN1JWvZv4SJ4r52lfAK
Q4X9VK0mNPifIOI419aouKEBxn4U3+Uu2kYLYFck1a1j0ukaRY8Qa1EIFmCEYGBvI3reui93i+Et
NKlpbbkRe47WSlgE2slrFbb/mt8XwmKm0RTyf2BHlOOTEHOy94XgPfUDR8u+1/3Ve28qIRaxax5a
RyhbIFvyzayv26Xjqq9lLpvyYwCQk/Sdz/VXmTwB3HntldleWxIFG7vQwhb9D56TVMFMd0P71O+B
T7SIIRPBwT12SJzC6oL0Nm3KjviZLKFDfqNMZFCJrz5g9i5JG/ULN8b9DhLKkLH1PrRG55fJX4zc
K/Fidbb0XWYXacz/yWfyi3UBtZlz80uY+fa6bCPRi95c5GN6+mg0l6a2op8wpiSPuMUhvt7xA4YW
Zu63jBNhyJNQKncSiKiqjChME+H7K2lnfaOGGcZVu09ecGlJv6nej/bdHuoRhNr03sUKuU9uPyco
lMWMNh9cK1MBLzMi+CG1frXq6XX+U0fsoBFvFLgTkQ4GlgnK90sgLM06l7kQZ//q/XqeIVqZfulg
CJ8xOaU8YcacPJJh2cFJdzZF9NAhHCpQFEi9h5JZ+hJFKDYmAgQsHNgEhx/QlV7U8lnMI7MkCDab
13ER0BTLmUY6gKsLwDTOwYd7OcJwv8vZTm3bi0r20Pz+rG6dJ38RhpIxPUcxBZNlYHYhNCy0A5r3
VozawMVFH1B9ETrFUq1ZjcsbOfHNxAr14gBxgFx0PNh+wbfbbYjuQonyj/EUuDEFq4hjSiXlrBUD
hmYumGg0mFyyohJ+VcmV1yjCFBR7PaSe0kfkokg1CDfzHVcK7SCCYj1BMr4BlQAs4IFCYLEcHrHi
1bcMHYz4VLwuvLP0lOQ+iJ4mTKyU4hyi8Z9V+UipkjJvhiFsrkDepk0VHUrx5oiTo1RmRQxv0Cnv
cU252zuTTMk47+jA0IxahF1PXD1nRmprZuCgCLVgOzerLzlUXkrST9axDcoLtPD9XOMyz1oET9vR
rt78Hu7pfpKQbquj/LEl79E5S4zEcyl/GLuQ497ujph6xz0nR9uEXV8rUMSKERk62BnlTI3PceIV
6HOUW/q10mswoYF8ekUn9oXm7uZ566LdhQiC2a4EDNgzDL6reK2HGEF4iaEIQSwSKfFn0zVw7/ev
VnZRV+NtG6bP+5j8gsSOGJ8fhGSBLEyZQngN/MgSz+Qlcayq1Kv59eoVvKBxmMBExqSYah1w50CU
C4vzJA8gjVtcEca/6UtVyvkIKA6417160mpA+Lha9LCmtOgRHdblDgfpRrF1no32rwMrscgxvR8Y
wRQamEG9PWzYrXg+V5AqmEYor8SeaoHMUW62EdO6ie58C3v5mBLRYzYlvRKHMPtrAcrhQG/DD2Fw
4gPg0mmnI+cEaofujeZ1FifVz+DHAQJbYSaThdja/Ls4+wbW5okisnjKIXuI1slaHtZpnqoq2v4U
F8ToK62ioHPTL4wBgV7pbB5d6tdy4O3a23LhgdhJWKv5L82I4eFbMUhCmQViDpYCaAbpSqcCcLUX
B+ebdMHz4jtzUfnBIa6VxkHx+3/Xw6ZnWUqUMT7hIyFt0FNVvdxn3UB73BvRigw2vv8aD2i+kuMV
7CYwoq8/bYLIXwMzqqc5UtOklTK8Z57VGibycrvBr6nEzwjbaideT42KTzqInxA+yFGXFZ9mBjmm
GnBsmw7Cnmo/Hrx4yFMJxXNEEj4otxUjnVp80zcTzC4BIr0G2G6KEy6wg+TxNcHXzb1DbuEIIRdL
j9qj4LP4H5HBE4i1k5MQhE/6mrdCAdjpdkseCXNE5+wt1yzy/keejOrqnoxiJC1EXsVPAiGb0uMl
qJJDIKANyn/g5WF8omeQAGtZHmAsalOLCsYPBaB0yJNb11et4NAoKZWIHgFGd31hyMAt8GFmAP2n
nEun2uiueLgptrnQZGD7Ao7c5mWKQcISWrngJ+oAvTTNFOwWuit1PmbUaXOywXrjYCwYNyuk9jeR
PsbM8bUdFe4j5APYYVCzSvXNzxPK74PfeyDcMic7UP6jIrCmSkfLE0NDtwVAwdBdpJX6u9t2O3mA
A/ODwlqyC/Fs5+3GNgmlz8DIDIyWStbJaget2u+j/leZJ1gSeoY0/IXhd6whB/+mPo3u7SB4D+u4
V1FjnRxSV21MHYJNEVwJO4GDUtMq1dNwJhW9G+SNiKB6v4T8AhGDvWkTTXW1K+KY0JQ7K2CCBhMe
8qFSZtytjue5q1IgM/fJdJRKoQQyS2Ms+krmttxT9A3OipNvmAwTn/t6J26ReH7PwBvJLhZlNS6E
Hr+N80xuYAr3Hqh9YDXoBDgs1RvMdfC5qrV3M3tnaBj6qCWgAAsS21weyuzncgwx7ktGoBEPOmbt
mEBTbbf9vBQgQ+Le1DMo1u+4Cyk+FeAE9weSihaymXzyG/0MaoY15W+2VYlcpJrr3+Juu7g63720
3TyLPXYJT8DyeDcMu499cwrbCV7UZMsVfDNSzJFXn9/pqJkb5P78RbKV2VTy8wa5VcmGgeKm33Kv
EaZ5eYs3J9U3J1xsosk7HkbWiAAwyOTYQWmkVnunTw/Tink8NioBSyj974zPiKV4KpV/qH3Q+YKG
CmLSaLLLf/hf6mSH9xf2lIQne+QVAwW+4mH1g9IjYnEapL1y1tpYRKfa9wPaTOgpUpRwh2JwKeet
X3/d5zd9IyjaIANF3GxRl4IOkKpQuW1mDDRBWK/VFPdaky+QT9DrPj0SWDPqf7jgPP4rBXhC70uR
30vW7T7setQi35Z8dpikpU8FY2VM2sQIaT+tgJJcJRn6/T8HXLp0UZijhBIXw7Wkv5vd7Nuo4TE1
7j+86rS89f1BbVR19nrbQ+EczPw7CFKNAoPeCi5HyfrxGRd/CAn7ucRdBcTyFVInTU0itUP1W/zr
MSponpsUGfUazS3Z21kTo0BSMcAFi9SDsQnv2S2VS7ypbBl08pYIjBNCrIzKeDzjmNiW1xNw3BQy
goKniRllMkysVMu32x62kbu5CaJ7UsRPOiTIUB0MPzMIgcqyyeM6v5m3bqESmGkGTXDQxflJOqOF
N9MNxXUJpqdzlZKYST2nz9+tnCbMbUV6ZOgX/5twabsbRhX1p4A1id52pGG3AiGdnG7bs+4ZF3d1
pSf7Q+9421IcU0L3RvIRcrSp4b1mROzyFmqBqcgRC3460uvfvx9Opc+UZ/iFHyesyiqbddNms7xt
w74O2MSUsHahE0RRCQ7iDlBXfJOl1EOkcKlUs6aJHJ2k6uSFE+LYC7496pS0YMHnzaEpXCjivEHL
PZxTd8WHp/79+QFtbbvU1a0HpmDcM82TTnL3H2BSG8NtWg1ujXKVl+6kAkKD3Ckvd0FHfDIeUcYE
zz0OsJ7fUExsWMN8Bl+U4VIZytoZKGTfJqEWDX7kquUEi79HyJdoIHF+RlE11QqC0g//LR6kT2nH
MU/TZ0Fjt1mLV9FqPGnHjnTaFKVvtc23pgK4eHuZvUDRjvBL+pGn3afyfj+EumN+LpMbIe5+u4VB
NIdEzU+cM0dCD2cbEfubW3dX7z+M51GNmkUXa5M4wCV0hG/+zG9v/pNJyjaWk178ww434l0pwxOv
IQmxHO2+rl6TqZvdiVuWXSWcxhz8WIPqthvYb/JPF/pVy++ODzJ9XeYhW2yPY/DR8vwP8f9LUX5c
Xl3GhGHUQVALozAvKkx7Qcx/umNpZTotUlvF4sJFXJpNbz33PyMMwL+TXuCgXGYfSDTcezfqXh18
OUx2arY6qBk2iJDGfzZaMTOy+nHNLPVrOT0IUwFYg9JL3scki649unti3oqGEP0Tc4gXznNacfiO
YzA8opn2Bt88J5dk8dYCTD+J7V3kHcRJMBf+zevIkz6W5rm3uiaNPLOtJEIhKxopAbWaqoeiso74
GvaSZRvxDrabLvcq8dgv4Xh4NJ1wRHsHDbUyZszUAYqBpN4G7yJtNWNR0qQs/iBv1MbDulENovxH
PYKGP9O4k+TQbKQQcXEl95ExF++ukBwHVw6dgQHJAW4FqP4F8P4M9AffJeYkN+ZDZGZDyP3RzYZZ
qVaPmJCzE/Vc5g25ESNIxj9RtRWSi7ABa81X+qBJPMeDpkb/Ldi0SC1mlcvvmfs9+MR1weFzj7Ly
jrpjZP/OoYzjRTAAV0lmh9oibxB9ioSTgElWtw7cOQcrYNR5OciVKQDLWjIcUfIrQ1xLp3kArWXD
jMeQ19AAbZG6SvVkwVub1CHLyrLWXxhwQGTx5D0gVmXEob3gLifmY9ApFa1bx0jOQ0FIduF4w7Oc
mIP1YR3zr9DtMdeYNAMte8UFD0I5Ix4P4o6ZnHrZPuKapb365Dr3A8xBu91UPiyGYsqoisut3kiQ
YB6DHRE68CRFwdq02ni2I5VvkPzIaX880UfRCrIMLmAFwerDXKyWvMEZgTg7oh6wCLY0BpPCW3Fv
GfBt/YCPnkT8on7yd3lqvS9l1xefLAiLq5/EAe8kQsM5lmuH30UJXNvaF01y3BPOh6nAvracPWEI
Es4y+zj5n1PhW4d/pGRY3tHX9MnEOUJLaUGkSmsmF4Xs/KXyy6PwCNA729MBH2uJiwzeTNLM4ns7
Z3ioPCmO8BjBJc/k7d5T2B/6TjXjcUQUzoaqFsCQBcsfZlb9XXQCBXsI9thzNAMceAjaLdMox8Wa
9nBgcE/kNEECrRD2adtRK5XPtKAkelQG/iahizMZpp6rY1z8IBkNi/1jlbTJotVXy9H7XQWoLbI1
+3ZFQJnymjjdUUI7+z8siaSljGrrHNErwGnnmCFCBW1owX8DEZ0R72OND1F/O2dT40IX1NcXaPOM
y64yghIKLDL0cRpub4+6UGr6SzgJ1JDnSz3RNiLfj5NxXitenLOA/u/GmmAD/ZAcdPuUx1HMzdA0
n9vrIJBHfSb2as5mq8/qgXQg0RB+pZVBuXmdkt6tqC3gGln7u+1MVyopWJjlDigX3lxqdiBxVU6M
sg2b0p1PcY5JxW2x1SskfAZd1xxpMhMLGTJNVkkKE4RlXs8woVb5tdZhTbOwa5YMqmaf7dP6XuUP
pAKLt7t68Mwx5MVEY3r9QrmoIFh7Nbq1e+weRXYVoiys8zXK20nB3XXOyKggJ95A2sjn86lQin/8
Xyx1ac6560ehMeddKEUoCrElAacQv6DGwQuW4rvPgiuJ+b0QO8dhKHxngGC1GWw0KOxiRFLo0beC
8S5nFv9urvsN4K84eyXcDC5K4wdBVNfkR2X9Je17ywjYVE8OTIx+qGyskZo+gtAd4UOucAO26EeL
Zi5H7wf7V2nNzAsShwr6OsFAkTLDg2lWoQTcoaK1YU2dkxI0fJqn8n+7OQTWU1XS90DhLc40RS45
cfjhrI2WnTC4AjP1IMHpZff3lc+JQZWxABq/dHT7cGNKWUgDYJG5UkObA7TkC5hjiWIF0jXInKHX
PT3I/2T7iTfxVtKsATCkXZ1kMrciRkbvTm5gMxv+euhIvj0r38EYKVLaTxhOsQ7PPnnshJG6a4Fc
9bzqZ9lsmYHDjJshJRiumn7dA36IcBAHuJqS7JUKTucO9guH3aoz/O/lelnaOCy7NnJzhubcK2bC
Rk5bKgpG4vtyHP7TOpP9pLcbQSPtca4WK7LBrr61lkjwwPdkaLKCxIE3Mqae6eTzzqD7bWqmCaiE
3zogFqCTXEedt/eZ7siGGQjdcOXkhlxPptI+DXYiukli3B/crOoVNyRyBPvy+Kah1mFKalgE4isM
eiKXp7vmQCOH4Mze7jLUhBDMu3Q7gNKcaRNkM/kA5t53QuFoc2enxTB+zOHwRaiBXuIfyWm5oxDg
kZkjY808GAGgnXAeC+1LE0UeOOumpjg1xrKC4EXXUzmloUpbcV3+ZbPflwP7XvXmBZEMPYGTyfGG
njpT/W50ahYFxRLwV6xvx1dtMB8P7blEZL+Sk9F/wiTpQenI6ioqc7nW4AMkLufBLfBiUX0gUb6/
tTXNqiKara9tJew2SakPknwkKAYdmHK2hdDOOihusJkcpl0Iityym0qoF097A3ANzD+RJS1ESaOD
NWNzwshogfkGEjyUkNTl1F1vJ7Zd/DCVuemJh1cWxBExOQ+Ces+9yRhXYHRKIyeObBjGXnHLt10i
kQWO1KGeUO8u5X+bSCTjzyfQS+POLOnjm4LclqpzVZugzzYDVYi/FjoPp+ZYyvt3V2Wq9kicxe/b
vgg+S9WR8Pv7u5lAoSMJ/IJ1bQDZlrmowvcC8DVxgRM5KKJZekeWwBkk7DfQ2hF282qeEozMz3fS
pWx+7UOHPU7u3tnJexlmk7RZkQftn6dm2SuV+Ae66CqqiI0pBX/VLHXbGZpM9tYV9LLqOcLtkUNs
aZMPDZaOiIRaxoZxpgcc5scTsnzkHXpEOKQ3Pk2ursz5+dtElQi3MpAN4vsW4S+5Ojg5Hw6E5SYp
+uw70yWCdnLfXrK360tIsJCVQlGvShDjkHjRoZO612IMDfrdCEO7O3kNoS3ocQkyrJfOZ269lIv8
epQgjWvm8Sh/1u/EwgLuykoIk3P4fRwHyMDhJMw/PK9EkeRp5wbU2IYIkIzNf9aqv7DCuhiCOqvE
ENSEK/YiGkKd6RtXQpz8isR8S2n+yJRv55//sKSKTfPs9qWCaN0RLanFlXKmhPnO9+/SdlGR+Qbm
RGp7AiOUlqrAGkjisW5QUSbE2Pu9r+eAgY8gd/Oudd/mUEwPfcRbnj8DTrmJDRtt2izk6hIZGD5Y
Vw4Y9flvua15ZTMEAAbbljtyADQp77zT/5wJbj5Sv0JdoGW9IKEi8AsLne2yNE4xKuruuEBrQhmf
VWBYnDMxOqyU79D6+pjpJph+6d7cRkiIJZQQfSCwQyuj7ZkX9JCsQnrb0g0ET+EYfELWct+ORIUF
kXHE+SBJaIRpG23jhkOl0vKSE5z+ffZMcRBeXpE7NBpRg7UuKqojT1IGjOcjTEmM9p2KMFFrSrv5
zquMHEOw54aPvcHnG/gTWlLK2Wn74Vg5M38wgu4ImKbrwM5ya/aRE+D/xaRuaRxpM95YDTY3TiGo
3th2h/2XUjgWTgpObxB/Nzc1mLP0izrLzIPfkH+YbdVecQt3wQRhpnaycmxRahC9xoEkUe5yUx65
6Tp4oCU5S6r8XJ/8eItTSSGAiCvz3apV4rR/pPB9qgJJH88x2m76MaxDJQe8cVZsWHAyKbPL5ILy
FalMw2eGZHUrI1u700dPvYC4o9V2kQDXdoWfm3MIar2sACvbTY3NItlSNKmLB1iEDZaQDAPiugiq
TT/1yctNUmanOftlQTHvPUXngJlSEnqBP+L2v2kfkXy/WSr4+oOGtWFngep/wa4I2hZA/chrgFuC
MwJ07XGTYYol+7nv3nxh2XJDR4sy/F2AEebJbghAesK6/+9zdEACnAkAI1ENjVrLHHqWFuSLyNc+
V/cIBkV6q+miCR2V9q8AaicRGu5UX6K3ANymZ+X0TSU3z1w731hZgl8ujREH+214IIninGEjf1Jz
INn/7K2rFYR8tG6PAW5wZmPNAFIPYCmjLaAusOd818MrCAWx0+VRSXrY4wBK0FfQQftk/bzsSpTm
AivWV313lS/1OkweZ/86lV0urP1AwIFg28bDxrguLPD94xECkGFe2GrkqmZBDOHaukvoFftNzsxk
RfaDzKgHClKsVaMZZVklm/DK2m+VqLykSBD7blepo2ak7mUdzVU3BBK95QgkSQ5qP1vYh5HLKVVB
JbEbGcliSH9Gh9BB2JY2q8gzRys49nPek6+mDr6x0+AeiGYKgXqDSVu78LarCoUSGxbx1PE29h6C
iDxz7dgCC/oWLEso6wP4NLK/89TUJ07CnK2L+S5Q2+fVqVv85YXT9XfalCV+SmlJw2uwtdkYOOhC
lDwRn6+3b8XmP9murYZvy6JqE1wfd0mB+wiGuriyathRjlZpRmqT0NLpaTBJ83KVBFTvdcj3l7p6
zHbhLeu5QWN0GYcq8Kzn5MKMR+2EJfm8twsvrJCtm2nI0Ofk7UbOxjxZ94a3Fo06BvglG/JPkhKr
GtaVAZ0ipHZ/KizbBq+0lRBBtemv+8PAt29E3SuoAwKUEQpVqog3UOh2j7u7YRuydcAdryIMajfw
bvuwFUtcG3PDU5ZC6i6zSC0g4/+s5tplkeV/WXMr73pERwTVx/H0x2qnnH3nODzCWsKaL9EIYejA
MXfpDTwWt+xkMK8phGupFD7M9sh86YbVTSleCJQyo8W0w0Rcu+XfjZLWtYjZL6q445dpXkokNtjl
FykWwsHwXimaidhdbWoVRnicrO9DguNlhqHcSb0z3ozRtxY8bLYYxvhcGXIEAAjMwzy1dj6ixqAS
e3NXhV3ZC8mSFo19lqM9x++4qKabsIDvPI7Ic2Ld0hzURdFqx6Gv6/o9K4butptfduJpLLpKdOn7
Bt19yfwfgeC0/ooTViqGJ5/DPIwQ+GmLULnZvpwwI3zzyIQJELIvnJcVB/G0l4rmjBYxp7Jrydcd
rBlM4TPy/nPREZhR0QqUJtVYERrtxn1IL/06lV9zQiqKDyxnISWfxn+V77phsLNp6fC4flRa39hV
SFs3CRkS7kQutSOLItfGK1IyXjyWcZLY2/4YosDy6UCz2GS+taQZ8J+rjdHLVi4BX1tFNYCH82jC
H/wbWIO/ob5gM9o53NcJBK3XM31TBG9pJQNe+yjjoqyv2J/LIsEvzL7dDF/m0CSBWsOTH7JxcI7f
XvI1tFCShvSGe5Ym7+KNnS9CrnTI69xTJbFG/GogD/sd9TqycaHOtoAltrXyDpa5AxSk+b1zq7tN
y4BDSpZ7IKF1Zkn4RfnNhI8t8ee+86+xzZXBtjMJLQRw/jBgolR4SbsVKfAIAZrTCSe+J2sD6R+Y
Wu1eh9F7MwD2MzzqrpLx8BqsQa3Gro+ANo+9TTHME9l+rEImVng05vpsT1NlrsPlAv1K+UZvZL/6
8C42cYC2jHtGqedhG687NLdXGCYG5yfljSlVfw9wu6NBheRxcNhWPRTibWv6i5ZQvhEkMSXJk7H5
LX3Ba0bAa1pgeTOdLtNrbWNwJTTmXfnlkvtqfrGWzAJ9lUYQaVWlSbGvA+LAPX844ydNVObfZryu
LQ2Hcx9d2nUj3nj+zlQGqKuc6iruzaKIdLzhKmnlJu2Xnbt6iFKG4OHNwGYyGKh8cZugu1GuIAW8
+AvPy4Lam5tARqjprsYx4GxEjCZngTKwLaEQnWlsMMEcxgOX+cIEOBdx7WIwKCBGvoO0mh7LRkVg
+NcWyUrcCJwzCZVe7PaVc6FY5N9Y+mFkbxF42oyr84Yqe1qZgXbN/Lo7hKUE1l5cQVGmxrvXgBO8
Oh5OVAeG+Xnn4KA1j8viypG85vsoe16NdSleSGoUkd40b9RVohaHtp8bd4AVm4rgLmMh0Fg5FoAN
IIDfH2I6MPLTiAArdtTbrbHlqWTQkb9g48KOmlf/99yBFuywC1OfUHZ+w6rJfXPJTxVdxMoGk9O/
ngumOVXPXdetbek2o3pphWCod39MBADhmWmjS/Q1xF+nt7e4BBQit2PFqwk53O9ZpQ3E6z3sKr+v
o0KqzqsHbBNc2m1/Q1ZiQsAwlvsZaNNSEXo1u5v9ccH+5YuZe2hobIWm9vNEnWAOFnD8s/8zn1zx
MmtdAqFc+TE4EXIM+G0WF9QrqujiE9eyI+/372Gqhm/0UF2n3bZoCGpcxBI+eo/xw0iV3fUWi3Vh
Vi3G8qHJ7m7r5uBcgStWE2C5v45NS+dlSFN4ZM34C/y34CRWkrpqmAMqDS4MSIrRoaXBQwXNy2J4
MMQ54wUK5ghuqiPBha7O2PiI6FB8WLiGWvlAfbZJC5/N14DrfDwaNbmCTXf2DVeiqekKoIQgg9S4
loCR0a8JHmR/+AZtP2OScsEOGYhEMdzXdSJfZW+xFTknNYwAwI2X5CGvrzjLEwNTMcahcs6H5LzX
JHVw3s1trReVYlGTYujtmO5dwKfMriOeiGyb4M3iY1tAFFjg2qerPbn8JIXgLQUpoPcR6SimhjG7
LGaJ2GUYxO8WbQAOiOmhZ9Xm8R5gRU/GbymF0LTwB9Ms+f/jmWwm1gezpKbO6oUEQsjRqWuN4I4J
kRtsLs3hbT6p5cRBBTIhkwrxZVoKZDiF/KJ+6le/kla50fiDhHetRbhi7uMGzyVZhjK0OB6n1p0S
xrl9BA+cmwTgM2u5jWeyHu2iif5HPaAZ1aF8q3gMyy6R2aqKNs/OCTyr9jA+7CwBYyj70y7nXDkH
iW+gKTnFvGzeLfM5it++D5qLNo0fgRdT2ldNsEurePyGiGyz/vKztS0UjGr/Qc9g24p3Vz8TDG3v
HmAOsJN6eyRKChPeQJFRFRMYFHSxjyV4tXyQL11GeBbsG38xFCJpfw/y0AaO8/JlJZ1G9HYpbSSG
ZBb1x18LUKW9m/Bgjvb1MsPEFUDi6/IdlnB4BU6cY2K+03obW6L+HchuIcM9mcm/vvkikPXDhCP0
hNyznyu3NftA4hJS8mjcHu8+0mbWASs7p2sLiEKcyfc6vtMHPLT/JrKj4J9FERJuG5hH1Qs1DFGe
xT8G57M9LavlLKwM30w6B2RqcEw4yS/7BzOIBu+3KDwAyFK8ORqL6E3fQfA0LdMxLyOPYyUgoVS3
QJj91OJxnTwjvuMCWLNBRjVf9FJyHErdDfUPTVQ70iIL3MlVR4nFHA2ielDB+ZCqZGFYYc+Gafr6
jgXJGyW/nURY1NsrzJc8n/uCFzT3q68aVWZ37mh/c6mwxYMYR7CzW2ZbqIuSpwRbDGvYZj0+lLtO
YwjmT+FaNY4XnBOeAWzPFpOBEJi9fSbqeKOwja3ewWSs5QosTSXv4zi2M6S3VVqyqsdLMT2ixIhr
vBsEKMF2SL5KvFp2veU250jtv0q9UORUXnLltzas8SLBhPPoNgoql8T0A55JrdTXfGzQJcKYa4QX
GB1QarUdVj9DkdSc+2N3fL+pG/nqzUo7+GLKiHVVq3OJrHKgNvJ0LfCyLXaPxgxpLp+EeSA5fzVn
XY2dEEAIpw3lWst572vtz89XGqhQf4xkDhZ5vInjKmIN73WsI0TkggOMnRrkiNXwe8lu+989Mvtx
VvI8XcrJk4PcMetMgKv9jiOiGGZj/ZFgPjWkXRjrSpkFGrHBfwD0VH3/QYsdwqtbEloFZkT3vmIc
Hvz5fOPbG/ZrsnhSqatF4HQn+v0XGDnXcJXe9iyveytUT4eZS7InZxElZk9LuwGJoV/H3Iw/xdjR
Bd1wAG5z1mvoBgTIdRnFcGMUAppnDyZeDop6nqAuGsGUlVs1itCs66c6jGDVFxCwmLREHL5H0Ku6
Ph0cDYWrcHKfX/H1iVmtbO/FLhR8lsbbctwZ6vfItS3BEtRj11enler4byN0fwiUTucL0KNFdDtd
QXrZJteQgybMB8lbIcQX3PoLtSVhQEu/r+OL/95orN9mU2XWLxAVWKlIaaZwfj9s/aBxrGbj/O4r
BQxVV3iymwyyWeQSh6LUD/aXCR5VHqoNf+K21wl981eXttktxV5Ch9y8Q1SHrjPCYmaGM6tRB5Wh
1T0r5OEJDW0UQTLZrkAClo81jZRSNNw/gCSQjmgecigNm6DLg5Fz3R6GXvIiHJFvxU/D+uSaYvIT
I6rkCYDyR7jiT5p47Lmei1g920ZG+5WgmbGgC9z1DlFU0sxWjN3HSbKOfRZC9hhqwR/bwnBXw36N
ftaN2pipdFbLwa24SrnGRA2is/S8QpNk0uUNA0380Wqa45DSq+sD20/WG/Uh64X1h/4X/Wkm7nVL
awot5e7ANVI7x3DJVIh15ULIjIIlLmFpeQybtwAQwqI3lMhf2ln7EQVmcBDztNl2eSN6ChaP0GPc
4LmxhisZSBfDRsbD4+8WMq+VjsYuInFULCtTfx3HsC/3yTRCL9zkYJZ5kqGgO3BrOuXRvBrBgbB9
AC0bEc8z2GTl5yGv7ZDY3zztWeb2+b1xCV+DQH0O2n1MNsEsFYHTJmiVa1B7PAO6byzC6HMZpHbU
M5XhcMMAkPYh2dIV/7m8lugYL8rkMJyGWS2qMl2YgfeS8MnCGqYnMys3ia1/mpLAxgPPlTbIUdaN
o7LtCt1pN4xCl1TAbOJJHcakFUSLrYZYnBGRwFdPv//jsRpCCaJj0KEy+hhIemWGhmoib8cx6GgW
ciztNEZP04mUMq+3mb9FYLhryvimY35fupDN2N7Amu2AdvqLJIjJTcxjK/ZvXu1hv7SB3xCXetoc
DmbFnDX62qgbcSbEZgWCOUcrrC17PFuJfxz6Ha2PtRSrowBCbeJV60Q7W9UYSwi3dk+8uQgtdgKj
VZ5kLEhnbrTEeYvUxr03Qs2FuNmsmF+kAltkHk7P4+RAuLDIbPy9i00lE9RPHbkp6eK8An+g4FiJ
KlYHEPHhOC9yivx69rgHTNppMIamwB5eukdEtHMgXAyfBF6NU9MkCUdxPjvVu5K/Au3GB7AwBVnJ
/VoFcBkkjZY6zlc15XCrlaXy4e4uIxp9wks2iXKNoywBMdSQj7FSYFfkxBHX2d7YcGkm5IoWJ51X
ltzxo2sYlCpopqBIQHVCXvyQ5mQY0zeGBrovx1wMLCSk1cRfQqz2maC0di3GLiBFV9giIKyE798W
kIVJNXmEidfc2ScwaQSd2KHa7YZXcYOlSiUpLkRrEzNMmeArlc4xa2wbAxFfapB68SIS7/3ATpZ7
OLL5Ikyd7usg1sDdWePCYlOm17gnOVhfvKRB0uz3/8iJ+n5RPBKfe2K+VqMQ0PbhaPh9cGAKS0p6
WREouaV0mgGrhmVLjXgsp66AkQlW5Y9SRqw21pKvmbY+aymSeI+EOiuip9g5HdQOvvtOfaUH+bBz
sb0Dhgl8E6fLF+ykjeNlG791dSg2vXkX35WS9N69tku/HSrjASSnBbToSSuitOpBI5aiG0Uyp6so
a2CV9NcWN6kQOl1Llm4XwA6DeudZeDWOnz/WQ569zk0ubraq40DpEuQ/87+oT3l1S8qEBSWq1Zy+
UT4oTZf31CVhZ/EP+K0G/1ZnHzETSQl9k1WFLJV9p2m3NzVsxcOojuXqT8MZMZJZ2GctYnNDbpia
dHP6yAY/sHkLs8EJpXnvBw4amTWRNxf35GNCjMHasfj3zmYHotNOqHZ9BIg5ktisH47LT/Lmp6zS
EwM6RmJPF9byh6bjXhZvwXGFTpw2DVm6PlFHFEpzFbH3Owwf+XQ7xeVUrEPmQ57yIP8njtEvusmk
nOrkqjaNMjtkRjZ4h1P2wbF1FO9hXLWNyNclsOaiuSoCdZMbKJnX4bPgUIj5yxM6X99ithc4ZhtB
kMwQReBF7+kyhcKE/yv0vS4xv5hHIaPr7ZUE5WWrL1FtlM32zGWJ904ax893l/cKXvu1o5cPk2T3
cfaPp6BtwltuAGDxCkCpWuTIkqE36BEGvPvTfEQAocTs9F2j6dU0mgL/zOuOrdo/QRuUVSBoGDub
MpnPVbtvtInogM4EJKwQwTwuJqlG2UvJvIgv4Mn4Z8q55tdRKuHPeCeaSbg+7KcEfXwAWnrB3U5y
pN0Np7ewZs/POz8FpjG6Wm/4PwU6pTmjlUSF58OXdXXD7WmSsSQiWioGBRY9ZsdTSFEq8y5ofP3q
tt5jnZzAhLEMUwY/EBzz/FgZ6fIdUnRiT3ixLeNzGBpYN/Hiw53jo6s8BfkfMNcs4SKwzdV7XBMV
XpYt+8eQKZOL0NUKCANBfPwlpRPnvk6OtPZPqtr5MQ9HPtM7Zw1UsEUnulpUp/8cc+iY57khIsXO
4i9aaZIm9/RkGmvS0NER6qdwdkCwXIiUfLSuBx7mAbsG396Ad5JSHuT1aNqj0aSLVSfgSQgYYzLr
gFm15jG9UyaCaMgTL+PtQpyir2U9F6MlKr2Z19ZAzCKMqaSKkhZYLWdcQc9DocnLJdvw71x1cmx/
FfBUkcYLw7PtaxAdpKqPVCW3jblUhkuRHw0oEwa7RFc8uQ1uFX4tEJg7PkQqRY8CBGTQVxjCRYfW
G36k2Us8xtzVIsqYCwJXgVCauv7bW57i9nWdA+G/3dP2gnY/TQHnfaeQVqLhjgtAriZR7RNRLQPZ
ZrRcddHnoXMoRqr1+y88i5N7Mw2/kIluuBxnBSDxKvVkFWNMq+H9bMzM8ztAWB2zPTnAgsZYTv/O
+qVliG2WEPbOgQTFn1SCauCPxuCuegm8+BWvMMdxuSEeEtUGU5qQeI0u43KlPb5JNN4Am9n12Z0p
3++GnYClWouH+PU46GhRzl3FRNsB2szytfknTOMhntA4aU7CPDpjyHN0YLepAcfk7zSPfwWwOgOd
jaHdOAuScKqQqBfxtmnLfGltCrxgi+Ze2E9MIIXzYjQnbncwT9Rq+qcMz7vy+/NiuwiHajhwQlDw
oXVAtDAZ6/PlF8LDKnYh6WRIH7hBaQTx6Z+rksz3Tj9hElbQyMKVuiQ1ueQliYbUFy2+SRWYhuzZ
40gApiwu0tEnIhgz6s7vjnBmk9A2M1Xy9O0vLqP91qr7Baqq3BcD75ifRtcPRA5WJB6fjbj5un6g
q6IB37ozXzusoiY6/1XTv2cG+FK96vb1wy9hIJtxngO0Blbdrixr/+UtN6sggG94bgBzrnOuGfsp
jNnPyFfVtLm1TAen84K5H2PXr/jAwOO05bnNTJIqryMJd6a1TS/ZYdFZWSyQAnyKPyQJfJYj8e9A
FQ7cR7MAUgAJFlta6ohKGpRVdsKbJ5rZPc6JZqyHwQsk8igqlK3JKwlMAUbNGFkr3p2eN0Okrek2
XT10ECqI6ES0m6FWWdk7GU9CTGYWfwn+VbYax1zhQUCW/1566j29MD+TFSZhK4d5nzFKqJJpXmzk
QzghyhOYO4Q/92fMC6qgUfgvh/ujlaiQexAo5mPJVb5b7d4s2qOVptN0lRdNLUVUhD1jDt1oMHIf
PFWveJl7WjIGAyhZVaxVDmF9G7GMcY93MVxgYoDPZIH+mly2MComx2sx3l5+JcUVbwYkymkWnSRy
Acp3aKceMvZiDjsmkt0oMdD7iE4N3rcebNOcXDzdS0pwmIUJHMwp7y64AKh8jieX2gdKYJVeObpv
MoAM/RuxArYBz0FRJ4BPdjql9ZLB23x4C0m3M8Ivmj5GxFcJ3JdAS3TXuLlDhcygIyCM/g5gcYuA
aW+44+AZteagertxc1D18NG115Ejca6wOewciIEs5fg8/THh74SsEnsAxfjaWMgeuWJPLBPh2tMw
/PhYWKL49opm6lEmoJs5p97skBPsQ901tSQGbnDAYKydGfoMtq9yJY4NGcg1bs3y6zKtIYws2sUP
NLbGKmD/e8Fv3sFj8lb3omi8NuBQVKTt0HBEe7Klukkai0cvIjX6JmHl/pgiGH9PXtMnd/THyldg
K525B8GNxip320iHT+Jyt1zZcuYxHL3Sbx9MX/Z8LYAjHThuePjj8/n67508EjnW/e5I5UytoZbF
Wmbiw1pE6/n2igyZ++Ew1RQlf6R1ir7IQqCXrsxvl7NGIJ6SyArxFNbMFLHuGPp9o9AC1aPcDMfL
33+KFOrJH4V2Nl4TjJ2ovCi0N6G8HhmVB2UH8C37oAnfYKs88bpJeJ/d23wj4udf+nzD8uxbPXrH
NN21upfBtOdTByk0qro5G5HN6FCrucJpXRZb2dcd7pKCq+yDIzlXs8v/mDZYgpzghKKkH+b1PWJm
rXFNlXBcpKA1qHlPQWe3Wx9iKBu9w/Jx/ZGKJbtlwhwD+QEUqJth+4z3NdVkMozYDxBxja4IVt8D
MvqwbSIgYJ7lnh8nhs2mSQKBhthvRSXc0toby5B1lQ+OxAGmqjMJEbTM6fs5W83O3ArZzqodGE4d
AVvQNPraxYBkszqi/4gajpqgbBLJxj2XYRs1aSn/8II57YUCLbvejCGZegGfn4XgmEdm73v44PcC
p3enN7A3eaj99Jw0qBpv6iCIP79+eZ9afThkNhF0Pb8m3cIoIqk+yGAMgmCtj3c6LZJrZCOEJkJ1
V0J1jR2U9xGKTdCktX0/+hgV0VUviidxG7P5bCWWShjFG9GxEc4tGjDGqx8O/ZVCHrg7HvGyK78x
HCIeZ1qB3VuMeAmelZWBaPVnpVNURWizigULBBDDRsq2Y6+uz6QV7CT+yxrm0T17bRR3Z+13R+iF
UmmQErCOkCfE+4PMVYM7y8O6ViAEnaWJ1mTfvWkKgr+/cf+dC+zMFVctQvnJRV+55EWia8fNPbvx
Qasefdzv6oUDWjeuGGmZDCyxfHONvuV6lvAL6K+biobrP22AgDevZBvnOHPMt5kEPeneV9jCTLq8
xbQ1uMJqXUL/yrpVp91XfDCcxSiOJGo0KclfynBJFpdkX9M+Hu8wwmNB46c9qWpXa/bfV48LiI1W
zudqbYPuMr/tmOuULGa46OgbzI39AaXO0LWAScFR68dXZSUfiR+uNhAt041smF7JNoOkCoUPZRpT
NGX7bPkJ84RM8yp07vO40pWpfzqbnGdS3D9hDXNI8r59BOkngXKvMSfMkuElXY97eR9+NhAAmsHR
aazrBZHdYUS+KPk/a3CfmXNEMg2bTo+NEvnIpuJy5xzMhZwlsfEFOw/+U/GULJAQ9xyFTAoJIvQz
fu5OWpHAhubnlTaHWtpUa5EC7b7NVfO8VMgXYCDg9tCcb1RdVS9NYQk60hMPs0d1gVT7xYj1Bl/Q
DSssauxg7ge8kjPlssCBgqKQXtN5kyg1/snqZlObxxSGelyt2ilFzcwLIy+qcUl3YIbTVzSgtKGq
5B1/J6XH1pFRUqNLPdq8Oa8WdMmGIJQyD6HkeVonAN+QvV6le9BiM0AtVDN2IoZHYxzCKFtXcWdq
PFtG1az50khNJUtobeCx/R4j2zVjHU+ZAhVQ0dJdKk520aoMA8EnTMs3vafqvZhB3q10NUTbriRY
MMSs+WrP5TPG1jlDBRPQykD1+xcoTRqd3sWDTQMw4t1y4snjSCG2/nK2vy16QfLEUkvwHOIx9sWU
yDimq32soeNZ3KOqNDF1oC4B2jS0rirSrDLCZIC+wKVt5izeN9l3BN2w1ukxVwd2ZsU+R0rr2unK
J+EyeXuyDPLDcXby9Nwd0fQ4dgF8pqQxZP0iBP8xcJkJ6ztK7249VUb/FeQc64Dzfkz3zWLMKPLb
lnubEgUNf/33FBemEhBdoqlJf0ryNfUn9aIawhSLxIVhMvRo/RWlLqVvCpT6II6wwdgSSOxPaiPr
Ubvad0u00D14IUf3IGD8Xy4Vun9iXSRx/IIbxapmUgVXX9ZhAUDNaQCxv3jNJsD1H2Ph7sufVXHK
C95vJsMocjCZW5aQEKXs6UcWDwBv/N78g4kHVeyUpi7WfmJHGf4J12rtu/BU+//dg3NgvamASuvS
sz9XFwrA0MT4sLRzR3WO5BH1mrzvFSv+iTJw46xfwXy4SbKPaOxfZlKVEYmox3WFFtZhNM55E58q
Qe+Gnh+xcUsu5uriV6h7hDydCgFl4G6yOEq/duXEykm+IXU719D1lJQ/Edkx3AgWDee2krSd3fHV
hkx96k8MWUhq6iWl4925mLDypKC+t57dJJVgILIS+ixVw56ytQhC8BKZovFLJMcBVKLNAreigfUW
KydR9DLLELbMhzN/6hG1QmazrSmPmBiOyMeZQCBaCTFzTSZ5DKLjJR0oHyBevHDtKi1fepVVpHeO
99zx/1ecv0EkySGzPn18q+o3N0xtbfPAlkE5jbuaQxJ/oLE+QPHUcHQCakEGFsWLAoHjV+v8/EBn
P/ThFty7uBYBWm0RTuLL0pVmaf3lMAbaMaVxM3/GVTGZgtrm6wJaqjMRTI8bXeJ9ltcLtYgtUWms
PJBpU/hhq79VIDDzvorZScfW4KjyWSEX7g0r+yipttjBZhXTth4erc6WVD6aIyDzdeC1c50GxDwg
83fhyM3gn/GdcI1DKGRYtpnDzFl5gbrVrMLeHeDG8UZ5TXMYT0ulE2OlpiUXPuyVEmiSbWE6X9Wg
gR+8V0ReC5roMiqDIUP8fRsALdC4aaFC6FC5HWukUJTYijWdb6W0iXnYsnM9YftUQK+7LGeFTXAe
RYNLf2TJ+/64QiY5FyoTmDzE8VyuSUWPwvNtsJFFRUsbLa62/KoHvIkMXKQWK65xeRSIhePRbmd5
BTB3J8EcoCPgRQSNDe1SKZ8cvl7yvlmmFmZWOeAXatkO179/ug8QfyZ9thCC5JSMTMhSXgs1Rq3f
6v5bXdZXFgoBYA28waNZbjUiN6WvTu6RwnHClQ16FNfD75/iUVDRStPGc/ymtvkk4TxMD3yocubu
TsTE10vTVEod6zeRW6KLeuDxDz5Zaiq1LW9SOy53DfK/ycd5leNgpkqfxpiPYQIdGzcJQWDle0u7
SADjYqQPqdoeiNBUpT85Y9qM2JCWT5uogBrgcvwiaVCStlEq7Tjv4vuiG5RSeTz/XUnhcjCDWQJj
fXB3OON+OzGu03nOuBmmiCJFDiF6e48DgR8fpNhdrL4qxKwxMGTWBd+oSHdqLeKNkRE7nUyMetbD
FUqyouzCPu8Aybn3ikBoqsG6Cslxe/oBBI/EkLmkIhcCcu0Ce3lSSRse5TVn/5uLk9Wv64gCwi1u
QfrT6oupfPyWLjlewU/0/IZGGzu5UEpybRuVTrFTY5JPpwvOuyzRGxeSCZUe7uF40FaTBcsfH21H
dz+gK+EhFRC1XJ4/HLpvCwlulMgTUCYItUOxXGon2N8bwaJ+bSYu/RXzheUon2iUxRb4KJ1diWEJ
2fWrTGKpnQQLV47i0YEeXdjOWJkw/79kyyFSacBBOMn/QDRNMxiVzSaY2XHTORwol4fxyllxaDFH
LTEz5s3ygU0BE39eRxpmp+bnkWa8xVkKscNsfMHVioRMzqfmU15kXnIh42w/DyMVQFJJJ4YfX6bj
RHJoU+mMf3y+3AbscBwn+DuFmtW9tYvO+ka5uA5bAhzwCR07Nanrjd2FSnSZmz01LqeGKcsoL/vG
fpNEkTGAabPPp6vHe7lvE5IwLGtARFvrJa0Zu71arKrL4oYxwHr9c2VnL9vXsvl0RhnkIXZ/497t
WxbolWmJHcBsswD/zT+hfhklfDHyNSOuwHMa6dyDc8SDcMq9r98Ya/Ba/yqv6eygqNWuapAU+/li
X5niYGiBzF1hgxLt+6DEJHdNhqtK1VB57RJQG9h4zZbcVeqv+2i0fmEg1VTf40uKqLQEjYaZmdDI
JZeOgK6tJ5xhXCJqEsXOQicikBDZILa7xicD6XlizIvX+JUkyOpJznig/nnnizZPc2sxTjg3Z0gh
xz64qdQy9NuLQvaSkx8xPNz6yk1qiynHPJwCVnPF6+7NhGazmkBtLIgaO5q64e3OF801e95LzEBQ
l6d3LefliibIPjCBj1T28zOVGE/gBZZnyBYY0hUyx6UspaAKdhMSnhSisu94JdxWAWKO2jrBW+uE
vjyJy0pSMnjlN61GFU/Haz4FWYD4bKQnkilEVcla45GiTqle+OcDwPEpDsEmKTwJkwzss/vh8Rp0
iavm9hvCoHvx0wf14fczT+YCPiLD9Me23fcmHJLVHt/Uhkx0Gw4OgLXyaSEzOpd7kLWYDeZXP0y8
Qg5Qx5TwS1VOwLESrn2nniKRhvm4yR626cTcY8GtRDLfZXbVTdmukoFZIm2qCm8wnGz/AlpgJhZT
AmN91+HX5HXPsfDa/HLrh5nwY595kmehw+Uz8LhT4EgCKvdOsrBQ16bz4Zekpqm8QT17dUIRjOEb
D2fAIXsEgG/BBZRcmeRWsKfvWzWxajq27khWtr5d0YQT2fOzgSmPLI1JI3mah5EVZ5agBzk5IeeB
Abn0kIyYAGg1Zu4xta8TZwNOIYNHL8PpYlEag7w0TpIzDnIdmAQQKmYwwvO9Yjt8WE//NqhiiYrB
mJdpyu0DDat2Nbim+r6nvqZ1Epzh58+YbeiERZoRFA5Pk0377h+D6NhOxqU7jj5GgDDzP3nTg49R
HlkVsyEDSyQ6K9FA0JfE6TRUXf75uaGonouda8myQVIVMRjyxoTVyrEWI5tanE/VJy2+duzYCMUi
gGCiupDe7i+TPF2pruRlnGEyKQxdljv9SNpSSVJqmSWztkIT2td5qSWnXRFt/PvZ8K9et6xrmmJ1
XmnilvbYPi4TWoh1SjYzfP8IwUenzt/4g4vP0igrZyYiN31dPZS1jsXSGWWgRUQ4sfNAqQBnLz+y
c2P5huj11lGFTwxHVwMBETHUtPhnA9R0L8KUpQapTdy1gecn0i6v8BrcZNZKC3PsKXpM8S2wiXW6
agiVIDgOqNxxgxVJr4/boOcCr0G9e01oAwanc4sFSR6efycxKp9Oj+hh3Lz9Md3fg5F025scYhp1
hg3V4RzuxraU3yXpr7pb4zDlIcLkS7APmfzXAxWR/35g0YKt39HegdWwLFwh+LLYJAM5bV3C9pi6
AQ6Mo9fIQ+Q+9qewWG5cldK3btcj8huQ1JAJF+sgh5myuIL9B78V4UVmSLJgCaE3p5AXTDjBDrlM
2mgCfTJg+UmpEC3Ya0esJ4tljF7L+2qM4Uled1CycQpvv56uTGD4V4mxdNWQkhkrkEv2RDN7f2kt
MkrYN4ncpa/Zh7Uj51I6rEhi0hGMlOkv5ZPTxZxMAC8lGM0rM6QEDL7cAGvGm5tIyoOX+dUJBjO0
2LRedJ695NVvwBAaEXH73oV/X2TcTCmLHT0Upiz7XP54HiAOUouqXYmEGU/jH8cnz0GGKSQC8pky
WGyfKPxX5qFmC1otImbna30mrs2I5LyJwvKl/hfpYBdqeVqz+NGPl77l7nyVw+W+xWmlyAVsXpUk
ZG16JlZpnocfI5iuXp/kp9ScOI3Vx5EcGY+I+98J63OEBPuokZyvinmhQYRjnS5SmtvbaR0U8ULc
IqvtdC0dfdERPYxxlcIzdpDVwliqG0VvTokrbFzw4FxkzkRhS5Kkcf1Pm25SBUHjv8SELWdi57H+
xX0nlSGqXawYsoC5kfVpcuhR2ca/TPRt/IDk8GWeLA0/3szvk9q2AeB0wkdBpJb6PvVvIfO4vkfU
tPwR1iuio5WTiwXYKJhbHGeavZ5Vizhjg23fC+g+22DaV8V2OYkiyj4Yrjzi4ge51cNBNsaHkFve
iqfaGIE44eS6DIWeql35q/eXOimXLsmYuMIMMMaQycxu1Z3Qq97Xe/okcEPaI4QUgLV9PNUoX2AF
lXtojk6NTnb46KiqWzOqaOhXcB2CO0R2/D6HvG5eraccpEcnbZ2LJB3in8YrW34B1JRtmab+qW+S
55Z/7x+Mlm9wfNXjdVlxWkLZ4y6dAripo8lJcLBpIZ4+77Uo6A3O3MMHUUAqHcQPGw3fHkaz8bjg
4SLWHpxORFFWWoT+byD+W6ITLpR6zYuoLvF9MF7Ewu0zZ9jkfWiTPWiOYf1eqxih6Ze3+S7irZ/5
8kDV7k37ODK5xjMc9NU4eWUppOV1Ms0eloBKYYOET0w7GM6TtDNzZJgwRxZSWei++b4Jwxu0Rt1M
5xKd6TpdFfHTTj3GXhKjq0ieGC4vkQ3NouwCMcjZUtBGRyMvxtjOcWbcbHcKhtsXgQnvyvoaqvO8
xUM9gY0NvMpz3ah6sx5qqxFSPYno3aNwXHyDegigUXf3VdxHxun2BB6e4zInHZYGgkmqNSMXhKx8
maheL6dx2/JCYgxRarlYlNT+mowycm73rRVdPCgI7f4pIv0QPsmbTWb2yrpt4xrzQddhm/BUTXZI
rcjlgkoyoOtyhh9doIM8xf79Pj8vk2LKaU0P/A1rVij63d46gIzwJhMRYfQjinapCm/CPChFcEhG
q8hCUGfnyVA4SNjaGe6Z8VejNidcxmXcRWQAtyt+57w4W2Y8Up6ySOEf3BMDW93JRMm9+Rf40Z+p
Lbv+XnUgztNNmtPjzqrxONFHa4a4K6r4TZfnOPy2Sy7INqX9yB8xtBetNJoHS26skgBbnua2sq75
TAzywo8sqcly5GJek3yZPqpAaqNKlmMt7IhO8VLmpBvCssZRx7Mcs3M0Q4XEiTTCJBkE0CTd2fSr
joavUL49OLuzxVfB70E+C1c8Bjpuz3TujH0wD3UpzMVex5J2oZj9CMNhadsWJK/1bsePKrGrm4PV
IK76I4IF5+0Iz6b3/N57ZHuCgbQ9gziNPDuvAfCBLsBYOa4M0KJAa9RlTl4AHjhBaoTJrfwLBvvd
2GkW4JCg+L5HCbG9JCwAJ/TjVPB4ysWuP793dvMmFlCvn0yZ941t+rQRZ3JeUJO1V5aEAGUFjNqD
xc7bC1bxUmevpWYe9wdEoViR1SeQW/pgJW5xXYnP3iyjrIZ6j8xk+9docBmLvaCz/jq1o3qn6OHH
MjOPAWGzmgIiWCyPWGoT2G8Qo7/NqYYt/Kl2CSar0MFCN+cF3TSM3ScyFx4s7f2dWHgC6Uc03lPb
lVG+d5OIUG2BFSL42q1Kop3hue49Q/S77p9c5/AltcUN+lhiP8YEQZz99w0PyQhW3IhrndMj5x2I
mkGvslXxjJItUmTWF7R6BuZpvUWw+noMgkM0l6n4t2a1JuEWqz5FygFudas3UeZxq69XfklFVUBi
Z2m8DF9zOOQbRY7D7QwGeKpz40m4MuplDJzb3x9NEQA1RQFnb0ghU9RJbiHTg7VDO4PaGf4nxnM/
IT01vVAG2d6Ggms5UPuo7NbERYJNG6H696qi7yhKkIypiCp+5yZKBKqyYNILhfA6ffkNKZvT00lO
Xb4TWHNG2LvbYg1aVBCI2Z1ng6Jy8xJFaGjdj3OJNLhgTNvZIjLd2hZQzDvZFKX89KjpjGPVYNTk
igDxxsIfcVOMJO1vpLyYpAOfGIHwCzuphyIVAQ3E9dJBWWJXZVR6Mn0YXrnBxPbWP0dC5WH6tJCx
AzhU3bRKs9JMt92EiCqXrRdd9mPqPvma1FbucwCR6gRcN36DhhnK9TIkokhgr+uBwDADG32TwdZd
Yzzt7Ve3c3yEom5nRiLmREKTinqk4hoG6rBtVW8IYyspFMCZ0oDgRuckiM42sCneH7UdXA/7/3BW
u0zdgpyvZlCWORt1Q2e+bnJDQIXvTnkXJFuoQd3Zo4gogv/HSczxuHHYWTGcZkSYV7hTuk7MKo9T
8SJ0wM6HsCPW412/VX0aqxSdjPCyyo0rMgCBM5XxSLvvQeKDYSVCz2c03NihQhJF4vt2EXVpanAw
zv8qVz2wBfZ4rINKT74Tq4x+j/emBvZ0HjLA7h1u47aMNA730jbzGQpLe2x+TZrduxBoRweXzNgU
v2FHhXTQ7UVk8G4wLSy9T21jW35Nqlt7Srx3WONq0QpFxYuDbjPFd/2GqBfPY6yRZ6NLIvRKQ07K
zwFNKmCUKBe1BP03/T1VhSrvBy6faFT4KolcuSaxIQy831OsTPHgr9hLqltLI7iFxoFlbBybcoRQ
EPRB/GtsLSAj0E02pW6sx/OqOnhugWg4n924z/JeQSUwbr3E7bWwa7RXAlzCGJIeRgZV4nVE0+4+
juiwGC2++K/d+Hg3dbLCSaHHFn+lYUMU2u6wXym/NUzgJsJY8hXnbMk90zvCMQp4HXLAsFopKC3G
WdaLNeTyo7MYV81AZ7UOrxh17RYyXHaEPi2i1KE/qioK+he01FfMzF+RR8U/5QUKdl2xuc7NrC6F
W2nq+XI279Ag5vIjMnizfhwAq9PfL4YJDSoRaVjN51GbDFqJh4n5qWuJNQz4kcGcIh7WqKIVC0cn
DZ1P6DsYDY9634XYTXgO1fWfTkRdXyF4MsCTIjNBA1G3xs/CvmrumlQ6WorYWXYxsarVTkq4HYPW
WP1u4awAXS5Pak5/g70E6Ax++pfI0er6YN039dRJ7M1P04py5fkPKpyv2+EeqwOamKrKDzTHDj2Z
m1EtlJeA9L7SxyM2uFXPoU5oZ3G/EK0bwc3wn5agyipXCZkSU0uXuzaV7n5WPhqvou2XhjrPNEcs
SfmMTKPgl1F++N23guTZhe17rvro7knzBt79VSFEt7xDHUjn7p6FmnmZ91WTss9TyUqYXqrfDuWH
WTg0u/NWu58Wmzcr4QfPu0bnyx18Ti8sXW/uTJ3biYmb0ANZK3gW+C227tXtf1FuyuGdYTigRmJL
iFbyudS6QZqx752XGxw1EXuPlfUFvEkjV1bONN1lZZy+kZ4PmemGxn1UPMKK4n1a2B6kloQ5qS3Q
XZZiSRHgfxyZfplJDD2Iya6wWyofo/h4omrH3hcQlrSX2i6kIITgi5WgaJey0eex8ozFPqa85o7M
48UkBQAyJqKok/OLaP992PKxMQJfwtU2ZKrwiPQHAfcmVpqhiLv6MleciZCbODLN8xveUuRij8j9
PB0xhubotETS6bZw4//vUAL1/CWZPQ+6OhlBOh0/+qJWmd3uBPRAmqVzBOks6kFIUp1DzQ0Frn5F
PQ8GeUMn4G2NQ0dx+gbebk4yLFnlCHSZNXqrBIDJwmPCIidUlhiX4/l94GB1wqy2rjDb4r2JRfdo
SLLLRIMwbbIYqwzq6/EWB6GPds9KucroJrhl5SC0iAGgxTmr7Mg29mOYjWRS3hgGDy+/V1un6hSo
dYbXMct+iv0CWLItzPAmoyN0GIGMTFEsk7Oh0cHu5vFvBmtnLQG2zsNI43n92058egvkaJiQnawG
NLrbHR3WiS6pAlOACsXWK696lapC+N6hDtblaiOq0+P0sydd2iaSEZQmbd8G9/XZNiNcoyHA4b2G
q7I414kEc9jqAVzvqSQIbK8shdUC8vq1udfsI9L35HTNNC6bymkMjVle3oUTrdf3fMrHIrpiHctf
yvzYET0iest6PMeB/qAApEKSjt8C1i2bvsZr5rKiqm46ZAfUS78LB69JCOQ5TsvNSX6wGtWxT8ml
m6gkZaSHLl3B7EqCfv3JD8R7qWe3Wy1DJu6sLmsclWV8xUJH7rruEPyzFo6JJTf/leBLGMtthEZv
FZvu3Iy9GaF6Ud4wQvuCTxBqub1msyWC46l2xBtGzDcRybrod/NYshV5ssx9vaoTJoYg5ij0yyIA
38NsKPpGNkzFZjw3pvfqZok84sNLD6SUe31f6GdUKFYVjBZfvQP3dBpz6EJnZ6+t2LB9cmcSbC/3
aJBRbIBZ+U5RqCc2So4xCzoS5++5jiwrkZyyqSHxlxRywGXkz2BuJ/Kh4Ch0KKw+iK1XaEdVBf+s
jKaxCrvJ9n7aObaMPC6FgPt5gnKrzOdkYM/A2MQS5oLlErpTm6xgWbDLv1VHTz84X4K001DNoD4J
cGpij8nNXzg1HwSzRTFaVe3oC7l0QK9rzczpPbGpSIE7I0sM3BLq9qxgtAFgBffXu7UA7r33qysQ
/wslfcPZaWCATqRLyLet9a+dU5be45IL3lu2Tzqr40KXA5d9VYkeOUTSGojPfCR0Q21Hr38ifDop
BqGNdY5DalcTgC8tpGxz9LgKRl3knNVf6grc4RYv5Z72YppUGfpsYfdRI109tuY0+PejzfKP+JtV
oHyp9wZJy6Q32rJKieEptsiFfQG4/nLnHwhC51hJQzCzT0b/rZ8yuNWighravZJSnNOAcXj4kLS9
clAx1CpFxSrBNtkSMDqn19uQ7hfHlwUnXsbMrBGXwhz8epaOKQHrqwKNgea1uNuuAxIcRrHQsJwm
fPLy2LOUYLVxf/Ig2G/O9az7OyS1zY2TtoMlkljOFZYXJNst41ge0PqNdXdHGOInRSp1X3/x6AXJ
Vbr2NlUKFVmMiru5cDc1O7f01Ggpmj1UISQNL765zWBCAhOY/kKcvb/JJRsDtjmEMQCC5m13ON30
1EBOAYwm3fRmgtX0n9LnxBztmoyK8kANTmxcIyeiHM+56Zh2vEZ9HEiSjIebSEdbDwIMOJXq7cTT
j/8NcmJ/7RScjhY67D6e7XZgCX30vqmt+CZmYzbHazicVsCl0qeCiOie02yP5GscObCqNboogjqh
TWtW7EGxbli+CPHC9IhAe5JgpWSjfyddmOXXAd1+KHIRJtK15GZ1WTlvphZsx++d7mpxUh7OOgTv
SA5pFGoBsD5ctRHm7l4YGCvd70wKkGPMoZurR3IkeSGRgY4ik1tLHmIzKSLWmcLMGWT44fb0/Y6p
fN7zktTGr+ovOJHssROKrvqiUINvXE7troTmx6Ghm42mEbOlLpm/dFdOi6Iyrxf/os/cBNMd+Krt
Qez/ILA/0E0bTK6UfWYeuhhNWFo/CTXEmWxYzn/p+vYutkvwseGCghjNlhPDZkXsJf8/vMDQqGW4
yXw/jomvy6FaNU4PWtgmpPJYja/CCC0sMBcgTxt5fOLTkAWKruiZS2cxhGj8W96FROBp1Gz23xNE
sy50CNtW9JiXLIa9bFBAxLlNrWgzxbgOBla9tYdKu6Vq68daW0B92jJ04wNA9HZ4hl6ZcbYv5aMe
CTbPgf4FMXVGVvbltzbExtyHNcG+az9gUIsLpxJ9W4o15MpzBSnGk1qfoMnx/KjhCZyjXQKyM8BG
YlmX8DOvVT081wvlnyIYzmO9NUieGXYRlpJzZPSyJvQOLefTUt1hlPHytKgSapdpYAEP5RsaZtkt
kts+LxODFLiWeftS47Ec5cfmLDKVE+5pSV6KVVftby8AuU6L1WMKTk4uwIigqbtudEsSzoBTekzO
ErbXOUkE0Iak2rkrpCgJjelqBjlfGjNa3oTYDB+vTB2Dpnj4rYtwvhZxUzVgmnSKRn9EPGeXI96x
h06NWAIxPsUdOQL0x8ANk9WI2Z6o0Oq33mDnktn6vhbjUmMbzxCiKubKeyoeGTCgj3PlLL2S/5Bl
6mcP8GuYXBJyRm7sahIf8nVyL+Ht969okISZ1dlkD4BAWsmG0uvKxENsDnaI81j0lsnHcXk8pEVt
Qk+wqyD2LCs1YHwbmqeZf8lNIdw2LKT2pHNhk0yWy6M0vQ37VqE30DngjwuKvZ2XCUYX/Gwx8kxh
A4QqCqcqnxcgGytmonD/mMOvNUCWJD7wXfSo9W2Oqde9KJlYHh1wrfaVwh5G/b06RKBF6K+9tCVy
QqrW7h/nL4ok/t4d037Ut0AT8Ls/O+RbeVKPGmFY+e/tEMbiEdSiR06iNYAmOcRohG9o5Cq/1xF4
0OoY5w1tNfM5QbBfJW/3tm7dJE0pUJpFWIckN2+KhrUm11+RsWmQX16GTAl9JrLvxov/VsIsD0QV
/zADmx0a7epyCaIithlI5VB8rPE05rP+FRIa306pevThNdtUkn/HNliEDxlXmCd1OBJQGCe1oMIU
tWOCLlVqxje1EPRkYUINxP8zbOIfVUorBVNxPm2ncI2Z3D4w7DlrGepZ26phzgafVmeN2NxyK+bP
i9ur/dUClGlcKxUdQ6eZch/2F/HYL3oz2tpeewNA35jveThdB2Urf0HWNZqasj1VrKKmze0bIb8B
gd4H707CW34hnq07AEv/Pe8dNGZ6N8LSLtihgIs7sKn12+pf+Igb/jL+9xcgu6odhhYfzcn+r41l
H6L7P5GCxuV5hj1rrRBiEQcE72WUHnMPzgCklLQzjEabaN5u72ZAD9i7C8GOK1U7BZf3ZAzBZqDt
CrZmCgNO3liE0A7ySgR42Zb03lRyU+5nX9R2C3+vyzzlxAWunAfRyp+e0IKr/2Es7qV+ZD9fIs+z
fBVl2b+8apEPV5DYkA2WxSBwq6yWM59dnCdDlXxWZH2ve1xkGd78jVpDVFHo//hNHNSw+xg/WcDj
g3xN0bQOjEUvhalJb1VDBHP5w+Ar9OeaBXuVwnbh9i34GAIEj0gOmcZRPg1U1eZqFHs/oRsTk0ID
7RyYrE2yahXvLHWyPMswkavRfHF2/fHpCeb/vV20gxy5hjwvtvYzQhw9UHJ1c7tDpHT7EZZdsiqV
Sn4W24HUfvoHnLm8KKi3+ASZj2GrHW1OOH+S28EZH78BkCuL3GHaknK2FRPWgA5bD6gAo5eFSCUP
oxc91136jbpo0n9LEeVe+xGMOA+xfKVig4B48Y2ZEGRkrtk0goywerhp8HrMTiPsSX3glyDP6ajX
zz7XqVVw9U1fDBexJlc7wtIZhGjmxToA84536vpG8ALcmfNbmXsdZ+p1AmJdPzC3jbeS05EHrydG
PzW4NG3YcT86ZgYwh8Uj2e8GUgT0pmZ+d0TgrW1BgIJw+hTXmE98zVZRm1i0hgJVG59qcCWewf09
16w1nxsbOlF58nB37jiwrJEL6FoglzJt/3sgmac3rShrZdQagMeVuWCmnpwGaqxUKsh1kKTlynZ5
MaXES3ci0YX9Cv0vBE1Gm2bBuSadXH5NVpPwbgk2Ofw1RAQKuiqAjWzB3EW5J6RS3k4QFUXDBSwo
1Th9/6jaWHUP3GOrY+A6rsbFraDuLuwkATIIusUAnu7FIAg+HmUHj60lpPyUv2T3GjarU/6GROth
Zw0HUg1WGw4Sb75KYkIFEiKxC3Qt/4M0X5ySK1tQ67tTvKdpuDYuzloXbgs1bC+yYlKGpGkUywEU
j97gt/nJ1XppOYoelqEnIVMksHqjSfccoRcsbKWtRbU6WTwh8oxObuVbdwqCJqqAuaTUUkGDmDTE
MVLIsX44AjUpJ9aE0agDPCnNabdwzS4AcrpQaxz0xq9k9dsAKKPNyXkV6XIjlsFINkioAtjuC27L
jNmzGv03U95LKEaafC6Llm/fnE8luBM8zCLc0znu+O7aCoFNYDJdwd9lFBvr2ymHCQXK8A9VPH3t
jMYw0j6DBK+F5mMzs3GSVF8/a1el+9BM31R4GoCL67a09R92V53uQrYrtFIL835LT/bsFMcV0mg8
pxmNDd6R86TVJqkUlQdvg5+/avun3g+89I25Ojt7OxpBpA4S9RKFgHRQsg/hz5TLhR9k09/VleyS
wmBfKDA9OGu5c7rtWSzipo28mzW6Ym5D7p/d0jD99oFDUoxJWGvceO3LbQ55cTR+KG8ak+U+qvFC
8cZH/ps25e/NZvgtkFTM+47E5Bdysdc2oUtgkZC4Gcvx1Tqwbnaed5z18lFaDaC7wyi9ZIHjT3uN
fii/dLWkQ8RAcfdM2Xh+l4xDjMzdmMmSkgikW1pE+IdVUOqId0ze2JAJsy1bzwIaOGT+RxIKFhDn
bClPRPeZYaXuYiE64Tew4Z7SFrj+KHQbiAxgQyCTZOksCNoUALRgAEcgxh0jKwFIPb9uRbDR/iLa
QqnD5EUmJ3MaBkSNGT2bCGI6o36XiN5z9Mi9Jz33G8hPVUGBNbAJrurKqj8u52y5XqVLZNPjfjdS
JHu7/bq1IeYlHQxRRL+evY9a6DyxAsp6qbJIBCo9DQf3pOLW1F8DQskA7DZPmCbEhtisyWWrhbfG
zoynRJwtMu3FE9xKmFsaNuUs1yffgr0uKLLZ1/2CLBtEOg5TluKy6z5WhX5DmUn+k4WSnFiRazzx
Wgwl4Nm9wKn0Bpv0Rgz5kForR7+12Oytb9guHzFc1VfOoO04CZ0/jtwxFulk5rOEXt0Hp5nxO8UZ
t4O4cSxEHZ3DaNJizo0oxRBhrjYet73ktSX3Ba9wOE7Fo1SpTFXNS7HefDeE24qgpw/XHm1UT9+5
qnns1RE6niRkddkyOj2hsJJ6EoBkwgkcEEQs172JaEQpbCbudJuKpgYYygtYiC4FZfCEKzuqeNYe
kwzqcPoUeXIluIbggCkmKKPAfRZAc1hghkTob7RyG9NdP+S+LWEvwwdrI0bpD4dpAjK6gKQ+8vYC
zMB1rSsS4LAmc+UqsRzyg+e8g5cgRvkGXSGUoa9Xhb5tM0WG6zUd/i4UpcIY9FdKu87uyZrXIY/y
CBA9Mvm7S5vEnN06N1SB6Db+JQhuMmATyAcJnU05smCCQ5QtkhWIWGGEivPpqSClB8NU7CXaI5z+
wLqY38E6VuW5VL4EDx3vFm654lv6O8khw8E+oWWlKKjI9f+0sxLqbosAEvPxa3Y2Roo8eZ8QU4sz
UxSpI+shQSRLhM5owiNri7dOlSO091Hj/6g2EuHj6VMjQg0JrJBtPTwidOG0Y2onzXpMWnuCq5jP
ApLbZpzOV483EC3gKGJ7JwE1dNDjhIBpyha4Sk5regKBjy56SlyGGrkbzs4ibH7iSciWgUUYKZ4T
bywXtaxD95sPW58qSbtFczB5qH+SoaKA8yvnOF0gw/xK3EXexzKd7L1DLXT1ckoBRSDezQIAnSUM
pzckqgqo022QUJ40huHAkyjcWcewK+l+GUDA/byu2gVJdx42k6TmrCPKXkFy192wWFFIePN+CkRX
s2KhMWj5m8UtUeRwcf0kf+7eWiGvK4elI2ghx5K/nOhyT0nHZ4GXTLWpfBhkcjfTWciHc4qBu3Qg
WIgsL8kAl3AA4RzdYb/8NGM/mox8wlsglco3OI7U0/ww7BFa7W1BNkw8W3kGZKQsWf+VdthOFqwL
qoVnzirg/ds2ZfBwV0gk7vTzmSM/n76gfKxlxlj04LZdZ84u4arjpvLQvSgpoLD6fipAHaNOu+WC
tlLCBdOXFkKP/ixWfN9+zBM+wbUSRWG6aG3Mr3Knf6KNrdumVZzyXUBNG5KZpqFoAIGy2b9tYRbB
WhByJQ3GoB21oVzUGZVJDqzgaocwn41mABx0yIZzgMbibkbK6N0vOu3LfX4U5wjGyOca29KSDH9P
A7P6Fn7kSBcbUcSS63d4NMersJ5Hhpw5z60X5eaO+VUO6izTTTBsBoIlgC+Np4S/vkgiVw+sxVSs
VXgd9G3V0YHadgrGwEu0maWXk+FbYb8gWX01HfEc0XtSypBStXbBSMi7zgC5tpjy5vZzHDwKdzA8
f0Yi9ox0wjEJHIsbQB8mFe3v9zCFf9eslQgJlcuipl1g8UO9Hh1WAaHs7YnumwJ5AbsC0msKtZ3Q
+iKTEosllv4wUz33Sp0Mg7iTCHKDp5C3qQxIOJvWM/OGs70A5nc4yYXJOnzhU4JMaujwF03jRFgP
vRNWY07NMyEiBtlW8GGptZAKmlg8R+NCRu4tBJyDrfmZCtMF3gW4Y0QkbsAwYykDHdyUL+D4hsnl
bV0IaM+AyIzbvm5QEXFLFrWWdxsMqYEMdk56DVbrDXi7B5WyYmfBmnOpIuTzuwa8s/+T3C5e+vb7
olTP9+moRWCUnQNMXhSzIpEg2fVXBAAad6WdV+2eJdmblF8YUO8pj2cgRIW0IWpb7UEnq1ybrIun
U9aaVNPMa1/lOscxdEeC1IM03BDYhlIc3DEWaqFEKkUTI/DLblv9BFw0iN/JdIjxDWUa1LTuOXiY
60T3cftIYXrkJ9e5fZnvqBSOkjrbSUlAteXxiqwRshNoIeNmSPfRucCkVHkvdK6pA5NU4HBmCddl
dVrrMzY6KcoPzMMY6/ikhbzWpM/FFiD0KmRIc8rdwJpsnqkle3KsrOP/BSUaAI4HvFCeV9BdgpE4
BxNDapOQhxdqWn2swVnbMUYQvErSxvpyBLzJOtOQvzjgn1BZ7Ugm0ePg/M+Pz49Hbs2+99RafSZd
gbYeS/A6vvd4DLnBWtxf3TyZUS5JRhvLX4qqjUi3VhtgbQujHyFJUUT34jrbHZ9BbpUz9wVXhpul
vjmDFUfHqPMf/TvRgTYjfep3Y7TmNu8c0JhS1TjQxvh/GEWEMu7DpnwtUE++5gekGiOCFe+y3cyn
UQ1RfkLGZmxYbKImk/dTKCxmBlHusewcS1M0RWpqm3/10mIHQRowQn8/elQ79g+8keUgtMFqx03J
2y7myWSaZgo2i44X3z154ZhPyma5bPvy9P6/PWkFqk/0dwsibVQREYox3Lrd6JHrDSb5x+vqw05Y
Dj4g0OR3tUSQ3v9uTSss01p7MbYq+I0A5W7O0DA5DwesFYnHIVgIMyRi204eZ3xgBpee9SBHaMeB
fhAsMxIRDwGs9UQ8SMYGAksG45ky6oJzXvxinqxHKeYNchOYnfSU9sLblYki4AuUXJoVwhbSD1uI
RZrwghDrPQpqFHo+N0NmRPk15CRA61D9XUtLu1164A9fz1ZSqksS1MkG06jcC9aYcObew8SUqsyS
h2ubjBMDh6UpWtLFhSSVLvmw1qi4fCxy8ls4/Dw7i3alIsdCyMJJ/n8afAX3fnAjwMaes+ghcIE0
/8+riNn99mJwWRaoGi+bUSp+xZ/kUv1HE/Qp14xwOUorn27XMIg17+d0vktJaMLLSS4QyoVf37Cr
4UuYq4cv+kVkjNxoB2jGzDT6rUD3ZJgGjTKU9Oj+UxVDlzBFmlG93lq8JzEd6axoUUQXTEAfrvbb
8hpoWlhnhFRgCsW9/sMUkj/kMIRiqky8klLRbxVdAABlo81wV8vOroVKjDYUN1f2VbhdAi7ovHL1
50GYY7+Eq+CVeryCFY3IpQilO51hROWfdIUbigx3DFOilutJvp4XXBW2JhCijIT4Vk4v07b13y3Y
BF05u7marrUImyGD4DxrRSsrH8Zo6zp0L5tnBwiDyu9WbGP3o3r97Ft1x0VKcBuIzBTHVH6cCT6H
VDVtHxMdMeCGaNQnH2o2JFEuViikxDVKhjUnnbf5I6sOcixzB+0QKVJUT6a5NiokA1KP0WwgZw86
lcOrSCKItDYiaC4XXQFT8nQCG059U8sGExIehbaFKuEklGU8gg6mw+Rensu//rpxPAENUAc3jezu
W/iEmdmFvYF/qHOxyOnDk9vkA6/WmhbEQDbHoYsguQXMZfuirbSeH0dd61inxv1pLVAOIMPjHK1S
UxXzyUFE0dN5vS7sh9x5J+PyJD5rQ7fARykAQ+23PZMN225uObnJsNh9r6dwA6lWOYBxSx5jJbMT
aXlsCPA3Bbnro43C3uL9c0wEVn+WHTzq2M0w7qXPPh6BoeAqXEClMyarFZf7H4aIi6E5aOp5ejg9
Ij6M1196VyF42c/5A4Kc0eZfsDO8MIOkRd6VwF/L5vwCFlj4bcxmVgNguyidU4zyK+gUGFlreF+X
cMhFud4h8SHoJR4a5l3gXNhXrWvk0bisoaLalpgkPG704HjHc94pfaog1QaMcum91Ja0OuYH2kiU
V7zvqiFwe+ASZmoHIPH8Djz8ltisLO4Ca2hYvjrVdGhHTWsDtuobIEqGK9Fle6z9imAyOL2rZg8o
MikUygCLXBQ2lqHEXrKLChxa53SRfqu2n1XXQ22NuGyqyA3td6qUQdSYGb0t+Qk/e/zSjSqVF7/+
4BGkiy0jjUkLuGpfDTOb45T99317dE+llpK4NJsjMPYZsY2LCfz3W1ygnMiXrueuASiEt9Sk8CQs
fXB4hTrFLQpw/X4SLO1E2b2b9V/Q1LuOkJlDofiJZ3ax/6pVIwBdMhi4GWAxgDlzSJMgF9BK7KkY
OaPWcIAN/cIuQeQ89RPKhBdEvV1+fjaWiMenX/XxMr9+UQB4/3iDq/NY0CBsVKyYgfSijdtOU4xr
DYbXKoSIUPf7LQTb9xkPeipsCxwnMUJCNkhOIMJmUmTuUNGc563BaZTWEyorFhR5NtNw0CLfEA5a
HgRXjbjYtF5YRyUKMAEm+WY14xwIbNHnlt7vqkMzhhNfvFIk5W2N1eTFP9lrk7LEqKw3M6B/CyMY
Zttg9DSwVrGdjzc+whcSsDBmgTMWWeNUQ3tc3WeRVNXUUVpeuyKo0l2/uD0qHCaM6jZn/Hy5oHIM
8Sy5dZrPFRlTdK6scrc8dbbTOfOsyqsNMKek2LW3q/zA3s7Piev+GfIPijKV8AxFLmjZxEAdsaAc
qsVuOvT3fwA3eJ1bhF5M47QKF4c/1b6rNy8nJI04T7jnZitDEXHFhSGNdiaTcyisvlEf6HMPkFhW
dHSfLAKdGInPO/p14ZrviN2NwfJ/GYn0PmK2j7x60kwSl93Au34E52xPqyjU6C5N0Am7UzQiIWoi
jUf/mixeoBMs9cjTx1VJD19XRGGerubVZz2klpmg0QjOd5L9NcnWY1qkXJOhD0CMgBd+lXtXeS+M
j6bF7WDAD8IJpBWTG+kaDvaAwm/pcBrzVMiAWiLDWfIUQIuw/cz0binA86JJxcCI+o+NZHnzMEHO
UVoEW8yfZ997XaPTSXQsvnMHMLvC88i/qXdn6e7gcIEP7f0kZ4lJg+s5PdkM3bApgMVxda5CgI62
z768WDIQuMpV9u/eUwtGCjzua6AJePMfaInTEYjqsvRshbllxEs5WlU7UqnM9KbfDp0K8JBvnC1j
fcOoiiVSV0OZ7UHMe6R5rEpfhLu+e205UYzMzI9BPiuzCDKll+9kqouLIVrsywwhKoujcyNWNsv6
x9ZNxZqcLgNDzqm2MmJ1gImxz4kVJbK3jP/WxOeK8C1gFLtjvT3+/+gRbt8mQbirnTvZoTM2L5Yq
MQXpquUU68H++m0+Q9uUq6whzzhiUOOPC0eF9v60woOTXMpvoWA8m8XL0frm+FSVZr8vd9mHQ/tZ
yIM3E9kR1gy1M3FmLJVaww+CztBAfiayhEHdd9zs8RX2hhwvCugDJ2O1/zZctGFT+6t8dNZz1pPn
Z1/otjmhbz7k6CXVBVGaSwNi7DMTknUMrUd0KbcRRqsSNM1w/7Vsahm1BHJ+p+bjFJrIjXL63uxq
Q/N03QFN3Xt2Tu/0zowdbo3mrB3H1UW4z5Rv7j1idNrUw2h7TKj4QGb3uM5nif0120pl7KphlKNO
fesHcSS2D0UQMSEAuq3RKiPvWHnF36O/coW7+NYRbqy02FuTclcSj8kRv51uhXG98Ts2TEVdt0V7
1JwwcI1Uzc5etAYWhtuIy2mjHFG4dErlBX984qv/OxsqH2YoBRIpajRx4SgnETsQpjYx5wfdEm+c
TDMFATzAyTzhX6y8KTVofe01a+lsLG0rcfeVbJQ3yUfCLOQuMRiwTt2W8RN2D1dwbSuzdwvGnKzf
mjkaETHhWBYnmiZKdCVeGqfNR4hRO4x+YmCMbEX0dkQ5JAR9K/JxclKAhzsZT6BZ/BmMb34lp78V
UMf1REruKKWl/xaIGTQhWVH2nZQm7f4kdV020z2KR830yOiYsaNWLiHWFFMtOd3ACoJAI1d8xMu/
vG+4MtBxMDeKLiZCdfpADfKTnzXtgqnAG5OXUWKNcLunxqhOKLyEENI+W+baQX+748uCttw69lBV
ExKnemh+E7jCoLjBOtzzOaokkd32aL3im4uc7HL/rXfJNN61syaLqDDju8AFK8uCq0PvW2Z5JuK2
osSCPQheX3TAEWIswMcI6vgdEJCyYSxHRD7mNK8egj6dDQsUNDyck+lDN/cGT3WyesS7goi3CfOC
4XZma/odkgBbNmuzlSKhUzQMXmeaNaf8YHgpM0HmKUiaRRHcEaILvCuYN1gbQmZqa8Fn4v8u6e/P
fi9wT6h/brPnW5M/l32ulMIzw1QQYs6wrXWaWZGiSUq+Eoe5nCBdVqm/3zvxF3aCy1I2BWcM46bX
UYvamlIFZOCv+o8ta9Fja9j3YYjw18pvoOfzvZnThnmbw3k/hNH/+VR8DwEiDbuZz2vw2Sj5L0W5
TJD7aJSzl8QGDitR9UuAueVvUW1nD/rOh3NvAVFDZKAap54Q2lmT7kgjOxKmRhMfGtdhXh4OAugr
v9yLZDrB+QxLrFr72V5gkac6tjWSw3ZJE56TEQUW4+1I2A+FCghmbC5YbvT4dMJFj9Ocn9HvrUFn
hRRhFuTh1xiFdBJKLoYfGUAmLmAGcWMU1nKMBAZspQ/ECTE1Y13Qtlz10inljoYVLJKhU4YMIgIA
rmNiRFaVExuhMV1N1EZYRrAe7otYNz5SsphmmgKHtDKnk0KNT1hFGOhpZbmGMMXxOsOyTUAAZjZi
mldepIwAGIv/h20aDICBaxNEo3Yh3kJtomio18DZRi0K+ykKxrpxg4Cun9WpnFdNd/MLgTCnbymR
5N6ZNRYawihpUm7DF78hgKOMfHInM89Fb9onnDzpOlnwW3uEeaQtqgtPbuhoPAeuCVd2a7wpWjDk
NvMPa8GrUhXTzPBUL9kOoPq1xisWIVPhm/Hgk6DmadNpcYGSGSVqlsG3ipbHjsQ8nQHVRvfZieOG
9N3LZWAO5sYUYhF6C9iJYmfcnKh69NknURstHmdujmPq14ZkBagKxDRlShMQl23RFrf5OJlFU5FI
NdKoHQpGdVYiOsoMQ93qMAaYlNFDCL+SRdwBHRzsPxKpKWKmXblA2Jvaq2BOmPDz17Nd7PiuE48X
LHrctGc1UA7ctiitI5G7RsLEYF0XmV8/STCacLI0DpxV6rd7Hi8MHsVIFE9RwMqlX000nca+7FkB
fZ6EUWSwjJQp/gpQ/9tPTuHfdMTOzCL3OEMqnu3tA89E4GiV+h+3ywfllZjU7LLJf0bgLoqHCwHq
GqCkXtY8NVkwGgDBL13KLTdFu92uMFuw6mK5m325VrxG3oaw/saO6L3W27SHhlgYbfqz4+/0ECJ/
LDq0TF++rMrEVZn8AQsnxgYPOzNuMfXlHZYgwMWMSZKXp7YkFisqdeH4gty1HeCAXvRE6YHeFLJt
/PE2VYWU6qNhtWjqPC4wItosgPexnwJg5Poy02ZvPZi6c10B2+XfJ8zPfYSUFiuZal8zAPjtjRpL
kFxrfzS5JnAw593wymMEzzYPF3rzEkpYUC60K4Bj+SzzNGCF/SQFWlzZbV5+Z87n9TiVlU2NKpGk
KqJl6E1Sc543sItMHTuZUoa2to19uWetGwqXZmGMYO/j2MiSypYRHQmPpwilRmZIIbWUCmvd3Hek
zEYDWsLXZS6RVK9/vCfIk02H7NHo84M+JjBeHQ40r5UgwXWmL0eYGznSIV4Ksiu5EzFx78EXvDPA
M1XNi4TDUkr7A1XcFUAjsnYdpC8CJOE1BSgka7dn4J16cSHAX2obKdxcaihAEu2ujlmLTv1m87y5
KA942JSHKfuczJFsEOPC6c+y3lgPaAPVBYvUoBAoHOzjr3hqp2YKcs+pJRREAMM2dtzqNhqTszOy
UGcmAenzfzc/LN0OpikEmufVXfAJBKkEPtAWNCLh2wVpAgxhgyX5M+QMWiYd/wfcSTj3VO7m/nOi
enhgmiMzidkTnWaVLru/bOCQJmENaJwG/Vb1YAAZoZYFtuzANqJpAAZvC66wwyUX4+Fi70bMHBXD
guVa8128fxE/7VyrWj/L+ZXpcJWfvCG3WhP0BzB8ydSE+mBaQ3ASIU+p0yPzt04MmbplQRIXXDiN
Ovx7MXuArSbp444SUnd53hOxgHiPwyK3wHtBWZ9yGNWjcaiu27aiZ1zaaHOGk7f2Ga2Q1brmNOas
7XXOJVtfo9DGfPLPeeIJtC1tCRZbdqBg2UIeKLBE7+Fr8jSbnMUzNL00PJYHKIWX2ng/1xag1Fz4
NIsAlu/XMSMMuODG1DLxzIhTBD0QUR/TE/LZHRNSOrpu4nTXFr6U4xKuqO/YAaBHbXvUhaOVeywk
GAO1ApRIrL5PxbZ0mCrnHn3UtXwhUPjLBJJVX8bGL08pVMgOUePrw3pOztHtRDArCC/jY7NlCUA5
LqU/9nbjf2kmKdkl/y0g9uM29br7JcRQYtnvOzoA0klLAK/kGm/ngBbmTK9JZzRMEmc1oRJPGFin
Jm1KRjejl5D2YAQU/s3uAgeaD2PBMm2nKfVOmvTSViASWNVce0KO4PXztyAcmMwrwiOJyqN6FLJl
RXlufIrxZy8C7e5P8iAjtnzUv0EIG4GE9uRPV7ArC5bh1k20OZwIcF6rlvO8mMDjwHBGZM+LcPq4
sMERttPG8qBaR1E6oKjWU82iH85Axi3C2p1p0UtvqN6g/L9Rx2zjLNy4OHebLdDcugky5x3RCf2T
YlmstJJncui8YhFhvj8dE5uWmRxt6GE0pT+nyRin2zvRY89Dd2d31n8R8+cAYtGVGZZB5hadmq8+
9OvY6wmA4zJ0rthMlc/8uFZeh2q0Tk0GmgAsc0mU4UIKCTqip+iP0GAnqefgScjJKiofbrktZTo2
NDly6OlB7G139z4avXsdyjUCdjt7Wgxye1PCOyTkANs6daGwRkCABD3ljfxBdC9zXZPMubTpIR2B
F4LJYb/ZMRGgUgZ3rMTUWdSUycGEaqKd5GOrCTetlCr90La9bmnGMrvkAwhj3lMIz5Odr013XRet
p/aHvSXLEE9dT9KquHIQWrvRH5eZkQ0mZgy1GLABD3TPtbP0M9AGIAeUp6l/R9E/lkUxhB+vbPW5
onMh+bsC3RQuaFy7UUXl0GKZ/UJ9y7ixHNHfuKWa29WT+C9Kk/6lJbtSSOb/mxIfvZOWWRnKMCOc
LWtv2GzYgOHWNjFX5tIYTwjQFBc4hLtFtmKZlo44FJaCT/jWwH7C2fK8aDn/WFBbQ5lDPO6v+9N2
o9izBXaZPFf3bwVUhw5DDDF460xDuCP/sXeLXIdyHGTGoeOfKrPPw4VAfQ8ILXOESJc1IV5KsEZH
9elRb57RF6GDTWVY6wM6/ibph9jbJeu/KTDQntmIlU8ODefUm2pDgF2xLRt/kcwmiOFs0d69MSTj
9Rtksk2uumXHMabTouqhcNIm6pFHmDCRTp04V2koiv4i0swvlThVzTsw/ObvGHAauWlwp2H7bbR5
UfkqlSXAUd7efXWGu9madzAWYfnqhzmOCFusnGJ7PyopzL0zo9DAoierO2ntKVLAvB+2TqYngsC3
rEwYN/njzgvFkOAAy2WbDDWCLgo7R4MI63xyeY4j/xuZNsu+a2EReqVu30CU9edmq6qJYIfTPUlV
mAAsyZss0dZg8YKFfIo78evbKwS+KVrG6zLJ52g2s2KYH2ihOY83BndjxnaYmZZdt6uo2nxy9RzP
yEOb+hLvgkaf+Sc4KKr8qd5LyM2aKY+/Vg2mbyxxYkFCXfC9S0pwcwhqIVo0LypeXmVaCxZ0M3XN
bUZA12hf66nPMJcCow/FqcF59glpX20oNmfTTH0Sb0/H9K4dfun1HYhznpH2zKY8LL/vaaXMLnCa
geF7FxRNECKIE+CqcXw9r/y/C18EdcG2Fv3lkB6qoUf19rG/SsvkhFrbm/LkEgbhdKDMJ+OXFyKp
bUi3eCON8qTww5F9hSrhm2szHrFYOxsOzSuCWjnsFldL0g5pRV++cOOAJ4+rQE1N3qvQIfZDJv14
Pm7ZXBAFY1mCWT8bBABCa7muEGhhwZExGpBHmecGyPfGdmonX3izyZcMxjFIFqmbzDNexEBDxBNi
uvaOkiOdIpVqyOChFohLSSmA6ie5c81S3R8+RqA3ovlzaKu9wbRmRUOd48EIcM6EPO6V4A4t/Z1F
gl8UXnIAdFe5m9Tp0bneOm+UJPsXCtmv5BuyWoJkyXTMaEJ9VWMEELmv3BCGjWXbudgfQ1AzvKcY
m9NDE47cNvO8aIkUc/QlsX+Z9zsjIaBMmwybfJE5jZa9MJY+/+4mAxrNljE8WpOGVCRY7AnrA+/E
k0sZT31aHNV8oBgMu1yUX5Q3YSQ0lBdl2v2KqpDfbAVBb3y0++wp8817tbfB1s6RgRVbb4q7gkQV
0fSGNCBpuPoW6t6DRBsJlGF39FaLmbS3LZPNwCp4xmkzB4L6T+ODRuVy+tQBnMi++NlASqEFy6oS
hLnpzXNG7uAca2n4yw8ZImxPMx3RjZkHjJkDriFTWXuIxFIOAZPKNGR/pmJdnHmuku+bmz8Vsgfl
2t/oD7NA7X3G98HiEVLp/z+NJQz4o2GLBJTzmlTZvHHBqDdMHof7WZvJVQvkQcM50umQxfuHiYiN
7EMe9MrqE/JIKSRCUPt22bAV66deJpg10huOe1OiQoSHMYjFeJJzT0lbI80XQFk3qg+wyOoRf2U2
GIlnfXn1Bj0Qr1X5EjdYvL5JMIN532WUAAjjlVODoVG4O+qA9K2Hq+awmcucXnv2LDYPwRxCnSj1
aXEYXjcVv2oRijDFiNX67vqub7FBVwSIZ2NsQ6Cip1gBo5Su/pgHvV/uUzMnf5O7g7yfQihWrp41
EVcpp1zePQWaP2qkSeUbMMxkBiH+7IG6exGoZ71bJB/zM/NwHUnlHRIsVDchphP/coI38bogsK3N
O/LXzajGiN+PFg4jgxkbnww0nFFTSulFdkDMZPRv5zWvZbrwUvN7BUNJt1Fd77/Qc7lK10h6j+mM
TP/2EuHgmh6y9dvUgAym99NiDpwWJoHucbWGSuq5zCHhUhmwdk572oa8doNsU7XuuyAzUDZiuChk
o4dzIBa30qrRfqGgpHHhYgMWbctidHWObql9Lo+S8d6M3zFuOHV8ED/gEGLsIyLs2iGAzjohwlxR
mcgql8zjFenARjReB04MnFFONgO6Tx3S9y0CTL5xbGldWZmPw//ir+OzwOVIfOkbEAYmV5rL9Hnv
Dn94YsX27TuXxshV9Tz/f2Gp1B90EKBTSNn7wKY+n6FgDk13UqUGcGT2qTaoDMSCdySN0xA0Kqu4
HbKekzcWgYz/aJGRVOCLE10Ps5dnEBj0imykrgTRgpIq2W92xkUFZjqWHptCLrKn26wL3jXzc+ju
f1D9amPomYqkgEdKPMYezR4meKrYwcgfcNmzl77NzdOJVYflDglUIB1L9gQlIK1Xn3p9i0h9mFtx
pyh46wTscJ7uGbVCGMCcVSbZtC/4MYms0uHBtJRqk1jMJLYFiUUcexWVAkIis1TnNd+8KcMLKUKY
eKh38iDwTzK2huDImLE7bkEPIT56jE4+Ad8hN0xhQXP1fz2gidd3ws9nPsx/EgriVrLFPGd/9DTi
eXIgFNH/ruKIbXr0LY9dJyYxo/tD8OMjTJrU34qN2bNrtGuoISHCfRyxU1TqJ8e2zMlidyllG659
igxUq13wvm4QWM165HkgIFClD3wpReIVIbPXvLQiI3n7P4pxl5aMD1fipkyKUeidWIIBiL/Um5Fm
Y2Wch1QbvEyp8zOmkn7AgM5ztQO4mWjSEd0DHYsltQrxaXGkT74uPGd4o4n7WzaAsgcFnz+8v2lQ
Wf0Bbwz5M9NWLC0GTaq83niLh1t8Uu62CU2/sW4s+B2n9Ot3TxWm51N8VuY1Wr9bUE4EHX9ErHSI
B2eqIVxnSgmo82aI610nguiPLxgvbZdoPfOWhW+cAT4weBNMHRSsPqVVL7Ek6Wx6xeDrlNNlU7GZ
5ilVpHz6wc5wxv7vsPqzku+wj2VYHapCTSL0YkrDLY1dCqHLisvkaOyfVYkorI0TWDZysA1STW7p
g+B6xuJXAcmYwbR3HzUW30ReJOEfT/dEOtPovuoIBW2YZr6tpBnCfVyaJMZOq8dU0LHapqtE405u
qAPX+4JcZ9CweLD2ayIUCmw3MMIVihAq1+/usylib+VOl4RQzj3xIju4AvX6F/D20Z+HaFPBZm11
fJR++BvdsQbM5miS1QxFboFMr2Dv2QK3usmFiJdgPpdYzZ5FKeK8KcNAJjTX4MWn/efQPFkZbJ4D
Y7rVIVDzM+MIo6a5ITPimezqeOfsbZJGtVMykAYWuOHrI+Y3WGk3cxUCEGAgae65pzwwJijRz95x
aAu5HNXRMuB2uVgJEY+fzrVFeQ2Ejxe9CqfOwI6xcG1jnrTtbIQBgCui+kzcWsEWA9qwRBVfR2IZ
awxT4olrgG+0Cfnwqid6kaKNwiLrvm7qglxVqF1H7nyTA54j1JLj+UcyfceRTzCxpMJeM+86kYLf
pf4meu4pZs7Z6EPIQMGqLKsdy6Z8kM2y/aOStJ1hNdhvt7ElVM6ORnA03B7OG2zjStTMgt0ET5gp
A1gWDZtt//EodIFdNEV5FPVXHp1LvO/U6OjedKQ9GWa3Nw+9db6Q8YTxN4mX0dukfqnkQyGrGUGI
errF05DwkprnhL6GqP7DJyVrNRa6V2ZAyMv/sLHfFyo+Wp+mN3wENsSmjaOsZ3+XvDYEjoGkdTKy
TofXa5b3Gb+NKz7J2zbvVQMU5wNHbkPtKSNX1TTQ99hD03e+Brkub7Jba4JKQbr8OLf0fpdpjGbK
PCqLVJ/6multuo+JeGPicJJDXwavpItUlUOClUUDNZQ4gl+NINM79TTsJQm+yzmgM/iLZeidx/Fb
wVkBA75o3mNg2Ne/rqKQLteBdJeb8tbXqGAeGV4DMHWzCdjSgRXjtERkGAstkuAUDYOxzEAv+NwR
galR42/K1Bdapyp9akiaIUwByzAVJNBFaIriESAPmwVVCX/AmxObEWoZA9+m4uPwGe2Q1hPYXmpr
XMc52fZUBkQM7fGu+FmW/fY/PYk4NuVV3tvezEGLzg4kv3/Izt90pKBHtbm39yRoTbL7Xu7fyfvi
/1iunelPKAqfaS1X5W1pLizP0BoMQjMUh7pH3NJw+Wymo723XZ/URa4T7+nVBfzhRE+oTcwdpmLC
sdX2EPtnMmz3lSuKKdPbAgbG79LbqK2vVug+9EQ+rGVkdrtNY4C1ft5qFbkSYmGY6npaJiinICc2
wnWehZ4JuxgSByGMfSuEAb38p1VV4Ob4KjERYPCMyV5Nvi/jApjvZGBLfzzW0fEk0ksWOzTg03PK
+g/ZDxlQBoWySDC1kuw/gjvpbwgTJqrpCA7Tyj+QAdqqmPxy1LpwdO1r9fZUTBcRNdAoJ2WvOFD/
eTgqElGK7O44IP13p49GxVO51v4PJPzkznAICzQnwgtUMxIGSE/6dBwZvtR35SYQuJDIZNuS++Bl
cHEuZQauAA5zkIoPVzDODCl8X389nQIAXWd6UiaVC86MOMUhA+1mBmw+uQ8OwForBvknQDnmaKV8
1CHfAqDJZZ9/3nFt88+ORkSL+yf5oU4h6gV7vYtDi71hcZDmyVp5eaDdUZmVMeeFilSk0XixDETV
iG0RWezrOvAYnTR+xSlUwQTklQ35Vj+2je4iZP8TCDbjF7y+E7f7KhSYJgQE3nGA9JSWv4gr5Py2
q4a9vQfsvo0JF7rub/X3eMkN/HaphW8z+0jr2Nhs0zkvQU+2ikCxZGGpPx2leBAM3j90qP+JhNwo
f+ZYvy4AY7uAxfWxmR2BVPMp0hG6MQhJAwfQ+wMY3K0gTAbQkTxWD/TpEARqu6qCBI2dnD4mN9Tl
bZa0gRSHpRIh9mYyxfJMQv1rL7gAdXPN7bGHQ4lA5y7Y/8CRvOosBBq7jAM08UUpRasYOKFw+mVa
N+nKMxHK7dRUDF+tdUNg+qp3wL3KMfMmqceaEjCejIyorUREK+9Ik7WgvRnsYB1PSfrgdofhbLW9
nhPrv+A/Z+5oTIxgMaPuZfo7tYexhovjypVIttPmVw3CRUMc4JyCjwga00qa5kQPaBo0HSmbbU9G
Nl1AT6fUZ7yWsj/1s8DjosWK3zoTxCVVbEddXq99Oy1O9KmhvovEZSzue2d5UbOGpenXLPhmcpuZ
4WphATjhTPJHzGrfzQS8f2x7wBmybIlwk47s1EtLxQ8oLvH/E5uqj9IzL/2CRGqDDOMz7wZo4YFW
GALEfD1wb8Kj/NvJnfy618VYF5c8/xf46Vy8P/eg+rFqSJ9hxOvmO+lfhqaCftIY3zusPfN85ecz
cQ0QRSIpiPg5sTPSLh5Ej83sbnZqlZw2yxK23p5L1di1cfL7SwRGmM+Z161J/u1b8N5XVFFkGcDB
lbneecyI8EFI9tjdF5pV9Pixyo5Ll8pAL5EYdvAAyoVRjm64qIr8/55IBAyfthmieG+SldcCFTp5
sCnsIYdxkFFQ4nxwYz4OWKi9Fm/gC7PhuIHq4CVZFNuQV4BUY1+klaaL30YpBygjLCbwxjAYd4OO
ey64aITMb3axHLzaaNOH5LWFmt/ZWwjCst/KCKNM+MYOYoqivIscu7vUZp0NhthmppylVxkLnn4p
Xp11rkE/qC6ANrmqDLY37cceDPxmRpiNyX5PE4MZmWq/5+Rn3NzqS3zm3kejaLZHt0AItJUB72/z
++cerHl5/LJMt3N5dKdd8SoI4Og9D+Vi2aqgBE85foh71nnvuBE3+bvGi0mRCBOc1XWuJUmEZEIA
cSFpVYHxxp8DorPsff7hC6tqe3Kt/E9QzdL0afoet7zs1niPz70jU7TKIr6WMKP2y6xlUm070qfT
cFd4/7n2/mKWoEFztgDKUR33/eK6iBCqAnTiQZDK/4xL02EeURGMEeMp+zCs1jQR6eYZai1Ztk6c
uFzWE03NO0njkgzCh7jf6J0q+U3HTSm6vRL5NR9eL22pp3vdiScezABm1ETg6N/kXZlg1ySjPAuJ
inlh4ANEB4NOvdf1mHxy/TPJYKJp3PBDaA0B8ILL2pYyt/9R2Ke+YUbC9UxWpVhKn7cmV9rczwMK
buupjxabpqyvQtlQAcYLBScmkS2at4saOQ2f/TlhI7gM4fj6qMX4hshj2Q5/p8mpxT3pRpVya4bk
RbhBd9V3PlPiRDtiN6EOJKTg21Fre41ZAZunNrfqNJa8aP3RlhQaxVzMtkl4HKvSln5TeQy+Xfo7
qgbaiGTGdc3Nen1VRSeAUYXXq6uNxqtFKmb0WdiJGCmn5c7zz/wMhUTJyfb1KNlG2g4S4iZ2MdxA
CJsCnG/0YWHPJpbHpHsdWcULfg7PAEXRVjO28V24AXW7HyW4TKm9bOMkT6J/Y3H5+byQ5bYvxVwz
y3ptuds/AA0ksmBKQtxnK0bHFXmgT5Ub4nVdhK2phzGEaMp8XHPtWRP5+HdZizXDdsTYSoBeGXFe
mXfzOt1W9UGkPYRHX60DMb3c0YbZhDbZrUnHOyDlzy4VyJasJd04SwtBRB//4USbMx4+3MdoEd43
4wAH+de0ChjpcBcTpXYU5KG0gpWkVxSm+javaxpvif4hEF9Yp/2DqiaL3b0qWGYfHhIW5eEfBbGe
3VNJtNJ5yRj+aGyamK3PFVKMwkHCJLFYF3OvlgcooP+HcJGED7kQLbP94GRjwC59A7ribdt5WNhu
ZubTT+tobSQDN5o/mngdsOQTYr+h+Tv3ESiVBuXTUB9sNv2vVB/6f4PI0YwV8/stIkGLrA6zI8wa
1X2EJ2MCAy6IxJ3ShJdtOqg4HytGZG8oince5Zsx33rM6XSEfQPMMdEMbMQ5aur+/sBaRm5RMIZw
3KVt0Dsa02reAPPqKgLK5tiKOhiXa6vLH5ekVXxN/plbBOMulEhcUiFIzfv68uO0iMCQGAu26w16
3tV/Tb1DfZDaYvguSHAXCL84j6eQpqWpuRxXiSJ5tERce6VfBClZRgjCRtsKfJ9648PG6TNteImf
ZmF1Ougz2ouA2Oo3k7eRXzQ7ctiATVAOp0qiE9YCEQdldKLJJ2NPt0xNnbPr8QueJM5NZJYHF4sk
f9OEUnNPKw9b8SZc5fCNDXglQ2VQan2RFiA23d80OP9YyzX+KKgklu4LoJmAfk2dCgFBKdhaj4lI
aBB0MBIqN7sADnd1JVWaEsoHuliya9WBXHZpmxkYYOTsn7HzIl3xDB+x4h7mxOdZDNdXe6ZpyAjH
87MZKg87gtrLRnv508kN8iMVHOSzpFDhXfIqaP4RvxlScpjIWPaLV3tDgY+EpjQ6rQuUDVJZqeOX
mwTm3Gb8sDIWgOSD5K+yyy/56quOSruLPqi+ucVR3hn+eHAPNfatlCGNLtic8YbcCKszhLoHCtyv
qFuQIV1Q3hkvEdf3CYsU9ovm8Hk42Yow5/JKNdoFr89tLSUw+LEgXpVOHI+F7uA9AC42kEnBgJbd
t1h2sVFsYuyUqH3dtDs48n/a2S0rYYeQq/AdXXINHTG3HyzZaN8LrIC98FIJEUGLXrBlX8xSanOm
PjkZx4P0vwh1oqTTxE4biGzMg2uTYKtihrNrTSvGLmUZEovAGt/qfnjpbls1SwC1hPtbruMttIv6
EjdrRHudAyGHzwNKtm5fIPOXtGoMbbX1t5aG9f2T5EbMs+5ajfQdRn2JN2sWy2lGOuFrdWCb82dO
pJenRGNomVVmMPbEBIpiiDkJZblnTnRPTGrWH2MCM72tR6M6vMDS7U+GnIvi5k5WGKYNnPQrkH/n
l8uQb5ac+8V7S47aLMnQhONEL6++gzKCf+FejdXhXNZqwvykYJwX/3jhoAZYghRUp6+hayDoE9PI
aujtEIZ25Q/5ZnRu+oEVTpBjXQoxlFt7oZLYZ9fKG+0iI/eQYBkg0FZjvE976k7EL4ZCNWlRmt1E
qnsxv0skCBHWrAOrYB7nYwj90c6mi2WNqSIQTjhs64hSwtsyFo8DDxFHhJnP7XakSJYmFE9pTfGH
nrwB5dEiObBuOg3hnaWW2viwwFxu6C5KM0W0it8jHZiifmganXUWld5xcdhXTXepNrccklYZj/Rt
4nwUKAk7FE9QENiEDQrMEOkcciTjqJHzHFKjqgjL5unYu4E9lyoTxZzGE1X/pDRFdz5pIGxUFkTW
kCQKBJuCU6w3N11J1zLxIrzy1NTId5DcSIsHr0yoQWWRHgD9TQ3IceGMcncS46sUJXsP7o68OOeD
9QKcf+OlcfUATVXfeMSSu6TCJBKnvcXuC0DPI/dF7bXXTSckvN6+Q3zVjXJoDmkbkiDjF6M462ju
tDwlp4GQWVh3ijtWzk2m9swMlXTfA5tuDS5YPo7f1TErloD5o82qAgA6DnQHBRMGeGy7qXThfiB3
2wS1OAbUFArLmqPeWBUwE8sA3CndqtFvZhqsKFnPy7yE7qURdlpEguae2q4HWwz34lqG2WVypxI+
oUFsnBJSdrqTajrPRWLRZVeNej8C7EmUSRTyVhEVcQdcrVV95UyTJpuFlimv+esnW/gyBtpIhAZr
e4wVMSTFAbsKyxB7buNvA0nSnNB9zZV0QYP07cr2vWU26oo/I4EH2ouI0d1JnwP8ucooRGPnSnDs
bUYVFCprW7QENy0c8YZTFUdHfbJC4xtPJ6PDHpD0wHW9fQ108LqyNipKu0KPJk4dDcxIUKunB9jw
iIhmWw1Oi4oiPPsQt7RVi3gSPZKUkk5LBgV3gSKL+1YYSlRTEdBcoMMhMt/7/9wXU179rwE8vKX6
CvVgyEhapN4tjFlFoFU+4mqP4X9nzPdbcSoHsL3BEnrvDFRMEv9sgyPQorz6//5LJXJXx9D775xN
TBJrKEbOVs41CazDVLDiYOixGLYpteDjA94zA9W10/4KbmxRsNwNv2k4b7jm+8z/hCYq8t0wtJPt
NakDyH73dSzpdiKNJmae0FYKjR7s624SIGaRRdCMdIUcp/U8gKusB3+yIATCqhLqreqcFzixSpQZ
RlHgfiBbbZPoK8a7DvUl3qA/Q51M5yYzHsMA8wykCuH//mppNCaemAmi9+SHpeyFVTy7+drKxYWw
sZcoWM0fge4cCq4tuxrHfi9SintV9BO6eOLlb1Zzb0uI1pr4siTM0ywzOR03W1uq5hQsH+uLfd0U
DQbVf+zBoKAsGWrdyVJd5tK9BAjj2m8L1xomc7p4HcBuvcfFcKIRICc2JLPkZ7tS29miD+L4429C
8Jd0J/SOsRBr0MFSimhrWom16OZ8Y7QYVxrHzk2OvyXDpb2Jv5Socyvj65gsQdM4xrZbLzFgqMLK
9RivtOcoTfDII005+kJOCIl8jnjCHopQSzE/q075fTPs8/4uJ+KnKGvReCTYXAu7/2BvyY7GJJ1R
AyNje8PCFwqaj4rQhzER6zM0gD9h6xp/1BTWjV4orKdWpibc3PzGQEKVMn6a9tX7h6Rlrm3HpwRi
x2LoU0klCVd8vGFEDDDB41KS6cSOCY+TyiI0hMHO2exAvc4hzuq0tCErVOhAnEHHuTat5kQLdeS8
x2H+yMM2MHDOLjmcnpi2fks9E3Tl/NH4SHn2ZQ5vll2Eq7sNYwrSTZE8pjV9FIUx4Sh3LCVbjij2
L1BpnoZYt4L2coUw9RaGVk2mFrihm7vg3Wunn/j5dXLo0sVV313la830pGQ9wN+wjo/vOzxDowht
GQlg0B7h25SqzLZZetMrnxjorJenMge5jxAbiLkzDTJ//67kX4xDOTVZFWx22KKvVXmatTN7WMgP
dazwvKQbLaxkLtoLfI3r/EgJ/fQerkSJrMhduzakOEevxAPUUSSkSrWjA3dEoH1o3AFvHnmxT24E
DWjLHf+CY7tOASF9ft+JtEMCaLN+WmuV8C+R1jARGCxvz/Ymomi4WSES334GPXfVZrhfJ/opgmEp
HUapD9l3ZRtr3fKtGPzGJ1z4p1IDskhjOPJwZ9WkaqJdF9LjIASQAiaKXvCZCWECww6VaRiZ2Qyk
IS8LWSf0Q3vY/6dfI9EaVJ7+NzCpE6A7h7InojB3DZkoio5nd3KygAKqRK++h7fhKvs7L9+9lllP
ZhmUa+zIlKyavEO1Fd5bsLVCvn1eKkAP1ven0Fa5DVuTKNT1PP6yUbBrBFuLEJxtDWlYWTQNtTBi
4cDTZMua5TutUZzfeMT65/ea2vjoQe0dHI8SE5vdgljU9ikKZ04i1u/oN3g7gCY0bhj0qHmrGOq/
1YdHNYNSBK4I5p9q2AyZOIdhb+EFDZYplSu8ZnapfBkMZiHkA7c9k7ikpqGdeYGqUOFhfvqgHKBA
rSyxXlAbwP9U9kd734cO1vou5yxxqEGTYdoznjMXCA7ceMpkqoS7ZKbJDy+19e/YwhsP/MGhQoFg
sQSTMIbPLAlZsENOnoVWH0S5WvjlCSKvjrOqi3I1/iu4oYwHlfSvpigLp/XGEJ+d9C/TtRSWPBcb
wQ0yr08oHYeotPJa5AEoN81Z2oZTcogJMoMqMrMkc6n/viMDgrUWJTgZOQZwnOfIhpVG6+kiASTD
qV5nmhmUnP6u054CE27prcCf6Q/RFx8LLDhitrCsOD3xPq37JKsNI4LkDqklbrexdqIAvLXwy8iT
NO1dOW5I0FkdGsNzRtrymgkpThZWFFcmeNyYNbdjed9WdO5rSyBt20LTavsKRUBv7jjMt4auG87w
9BkZAQ0IkVjuarR4ZAUCe+asQDEDifH2z4ZS6hMd3RG/fXxBB9wy/ZQPLKhom1lGP/uf2seZAQdw
8zyECMgbpqDoW8MAGnQIXXrD44HQB/lj/FHH0mARvaXWKuk98Rnu2yAQWy8aFjtIy3xnc7yxND7X
t2IHsre4uD83lycy7B0KSwkxxm3DLtRJ5Xn1gRX9qyUgFWXDsMNR1i27dzMXzfwJD8q6F+Tdx/fF
nKwDMsPvTqELAIHp1rNBbL/E0L99BHM8V1SD7zltk5KjIZd4/w6mJ1t6GtH22BpS+ZTdEtY0b+Yu
ccumSe1XHshFKeJ/ubWaax0tnBwi+mxNuY1s5OtBU/sSDmVxL5ySPlDXeABLbz7+lcki8IHYOAyQ
+snpFQteq7qojdoGl9hI0K6d7JvUuWOETX3lemXglAGnL2W+pcA90a0GH2uaguCVRxEjmkG9/80d
LsHKuBndBwKmHUAwYoROtjNoNjclkQMCpklJz52YHvptZU9/k92wPqbiXXw/ajnd07TZSvP+z9E7
rDg9DEI3RMI4k4HA46uVDq/8SGa6nWvq8a/lYK6pRaBHyRdiAJEO74l/HSZZJVGFH24hScugXGfy
xfgzJg7LvldnqR1P0X6Qv4Uu1RTfh9QFwYVzFZWU3sbkG8bFKj5fy+bt8M2lfeTcNY3a5ioVPUcS
MrMxJxqVWY2kCQYJgMeSCoBc7dTf9zgDVeSN5g5XPa+vs4/FLwpmtH6yqKA4P7Gq6pbCfdED9cXU
VbWYQeD+sCDc1eH/+qcH6WJ70f6JNkAFuPtS+Vf2V92ktyg1Ii7me8kqK/cBqJasvp5J2EI+zCsG
F9UnWvJIqoE4Uf+onem4X9Uk0ycR5D74U7fXOlQ1g5xlYxNi7ZoU4RfJkLP0yDuAIxogp7UZOSmz
eCUOHQO6gUCmZ540M8NG8fyVWT3r1uVZoBOqSdO0Uq710bhoB56u+VIsBI3iBJ3TIQes4mn/KOdJ
ytZfybyYhqdISdOvEVyV6+F8884YVgAHLJv5DOH3XEHKZ4JZYSB3FvRAtTF4g1xgSLT4LasIBHbZ
72TyweoKqvVqDkLuUZbohJZcH3V5a6M3BoOHfd91NDny6vYFoC9Eue0uO8DNNL2x3iY9aP6cs2X1
4S3coK0b8wfMHqLALTPqlStdPD0BEVr989nHscsJkWK0mUsAG6bGzr53cjvpwqsBApHH5mGqz3G/
rgzjBVlgAzgz+0hfA6O3eCDh5M2w4mmRev6wzfxizSPirsjqa7GUVQnAIH7LN8G5TP7f2vPSj3NN
etMxpb78AdZaxTwecfFrz9pFHJsWd+EL0GUzQuSgWRngfts6ynKG0j+FGev5jQSqR0STHyZWzdF+
h90aF/0GQvCmFi+XZJ7FK7gS8UkLpF0oi4OgzcNeajE/SFohKGafvhTwli55ICbidAm4VX/QmYyZ
3U6XqKbbriPjG7IgvEErGwhDQW3dYWBe3Pe94n3HG2ayIamIsb8IxaZ7kam+/ZVIA/Hnw4R6KZsm
JKdAAc0efexIuRpCidCN/ho3Ve/TQcCqTnbN/9iaKbAB9XR/f1fCqxu7nqY+ZZXBAstAhp8vnHCb
w9FpzCXEbMd+KuUv3eIf9NugmIOUS5kgHgRaZKFC+xUUhCsOXI9gq9tEFn0o/AfL5vR2JGG4RdLs
wwfIY3wFY0ag8j4IJ7dNuP6s1yQyltIzxhiQS1j+Tr7ONAyXYAVsI4uQBgr41ovhZMp79/sajlg6
30Z3rPVBfDM1S2y2RI35NC/j3uAByjPXwpdwuXBpWVnwSMmTGuGj2U9yx0teV+j1fBEyA6Qr8BOh
UR2nujZ/B/49usolsn+cqZ7xoGk7Hr3buOex8YkxkhRNcniyuCtqEem7FhokWooWym88DS05HeHq
8ALz2pmzsqShejatP83l/3mfggdZPLMyYf9cStMcVpEVL5ZgXgumcAlehN/qcWIJOXGexueBa40F
zV+nCfZGWNcLLCEIQQs0BbD9tvenk60DsmNizWeQUk/0JTkpXtMd/iyeRQi6wdecJ+qbtrlXoJhz
XjEYSWKvkAmdp4rtISD2QkgfcNlQUL+Q+XrK2FU+olPIqWDNKEdWAcXUd126+H2/i/z4SJKP4uvr
tRNbU7Aoe+Hcf94nosd+Eu18HO+Ek0Fez/AtCaEujqTqQxIO34bykJiqP9m3wPnt6zGQpCnMuT7h
VIGceNpYYCduWmZbyefwHLpAgET8VAInTzrtC4+QW1uzwL9+V0CjD3aNrPTpvt+UbTxRDJvWvEI6
/DkOPDLGySc7DCtX/zSeUxaeAAtL/AlmhJYxockHOCkRAYPvd61xrSiWHXg+h1DM4qRSJ9/b4XGt
M8ikWLgRNQlyf6J6mVlxoWAxMuKJY8XKiSxc/HDe6r3R25vE+6FNSSFS53g9nXK+UhIc+0DIokaR
PGn8YF61/UwWimcaDjavvLTD57fCI6pxDDE6AetLuorn3X3VcxYJyIb/hBeoYjz5lzMX7GaWzk/H
5xdIiAt06q3pcutFNJzDlZ2e2KoQEZmBbrlUUF2XwtRdX4V8gE5PwL5kMa3LZj8y5W60PT4LZOOD
x6W6KRP7s+jROjtUgazgu93fmXGbBPkyIeNUm0pxn1ZAPAqWj+rzS4vbfa6usVeEAcEL02+WVkIb
+96p3T4EoeYNmF2Xa4VhMi9FpQIW/tYN4/rsIJegFaZErddCDCPQ0HfruVv7amQQOtKTaEnXq9AF
voRnWabYd2o9dfGa6g6AC+YECSBOcWY3/vsewGRJpRCo02kCSI0rZvKCLZQpknu6NJwsj7yB16dx
T5NgK2SEQTZ5tE1gev4FUPL2PKS7Geh4FtvMB6ZkqjyaLqgH7WhLxbyuXmcyRxSIumiQhqSB/H8W
viwbftMn8twAwn8WlEwcOjRS2ykwTO3MLm0MmolMkzh2yDsrammMVzgiZn/qpCKXo+J6/Ywh5idc
XMqG9gSTIkJ7pZxk1ljRCp9LKhsmOrivOdRjiLHngMsxYUGC7ke/gq140QNkeM++U8djNBn1OsQn
3gMwK85X+tyRJ9aWtpj8sTNvaX4xqBGRBhznC+5QALgSlhR4+XSuv7vUQRd8M2TAZB2Wz+pAasUz
8k1tan+F9MKL2z7DAGH837Rcjqgn/LFjYx8R79fazOnUjwna3yGu3X9+dnDFtfuXBguBxm5GmXWh
4bJgT3OjLYPY96RyoU07CHyv4lkQxxuHJNAWGb7xv/mIbjCkHmOQdN3CQvrLj/2gLtLEppFl45qR
7aX0YGLtDT0wQWwP3fcJCYtAgtfx4k/x2ipiHT2dcL96hzr4FYki53e1KswYU3MtVKh7SvRDdBA1
L0EgbMC7gvB0TgqWOjHXv/YJ6TGdu2uaGePNd4dHEW2q7n/QtaMWw/44oPRW8LppCfa5xI//832U
9SjmVx254JaUzZF2yj2OxotdMbEOO920hnwXNt/id+pLhlQ26YRaahxerJycNPiMg1F2mYgtc+5o
18Y/5IHC88ASJSzpL0C0ePdNdLywOFA4H243Az32RIOomuDVJ7sUav5/TDiXJExXaY+7l4nnSeIh
5l9dOQqH7coxMZMQ3zyk0le65ZaeEyI3lpx0uvJZy16t3dtnsJI7KqY+jClRd98nBhKGO0rh/sX5
IaCPJ8nOZ8LKPsDFONPRxBDJ9qLrT/dxS0phpTgnijvG+9njDV7twGLCjK/gS/zzGHMQhJeR0zmO
kxqWOxmDSZJjY8cOha/nFz7OtmTcGYfoeahzKsCOJ+ECj+ofqnMK5LpixG/foKcM3AOGNbfElEMH
0sHBkqBhFn/qlpj3baZB0kTptV3oqXyVZgG+DZHi2gpnGTrOrhLxuQvCsTwcjx3vjE9T0z5n7v/D
6wsf5LnmEiZk8DmOKMWJtDJdWuysn0cIdo5LSpBy3G+3YLekQDTcMlBPLyO2pdsCw0h+ZyAcJxac
ewd92y4cNJtOodNsy1ZNnQg8X5zawF2wgtr0D3K5vQiEE4pC+ueeIQ5MtAnNcX0r2puelkq9sjQf
UD4GLrJp+b76qa4OBreAwQ4yoJ+8t1T0zZkHi1H3kUPTf7Ln81svyUok15o4bQZrBqL652Yt0rVJ
GB+4BWVQ3AlSBpC8vsiL93ylVHH3a1rEiaPLXMXDZaHA4zXH/DjhswQq4z9XnNER+Z+QqG810CsU
eHKMDD/0eq0cDSgeYv3zmEOR22jZ0iJk/30LDz0L5+dI+Uz8SesqdI7NSa7LFPWGORQZFGsOX5pn
EV17loFDqsK6o/hDuu59Av08qhKLeU+bpS7JZbcyZiE5kL6L5yOi+2nub3h6OPW1Zu+1Y1WjFVcW
KEC78PINoSBq3QMDLGxVGegJrc9KjKVKV1G4fB3blClYHi+aCmSHLdsgRAcyEtv5V8+H4fntTTjW
+m9vu9ka4d1FwrSxF7SmuvgYhBG4X7SLf8NNISi6gRyZKncllCptHNS2w4Ybu+RwbSaoS3Z5QbdZ
PxUdYWVboKfDMZyyem3BdJPp3KPJuINF+ark2IVzPpb+VnbnZIOOGfI+Id1vo9eWoLlm5NSXVSUd
hSkRzkPfMy2fKMiJPYxLi+RQPlqP02qAiyHeO+BulGoAvw4qha+FKfDAMFaRXkd7d4tWh5ji4Bi7
v3URDuhi8kumspXkJWlbw0+aYtNRiKc6LA/L/qqC/L/ByAeAkWh5NMZB9MftRSo+7PjXMtbgp6QN
g8o550Cju0giR8ceqBK7KqdaPSzZxj+4qja1okhCLwDHwI+iGk3xsj7uFibwUfFOtc9cSz3aZZ3Q
kRkOMdIqenmwISyy3dYkTz3faNfcsIFW4GPn16xWnuKKFv+dEvdElN5oOcbKtd1r43z815qVKgIo
S7zvVZ7GuxMaEOPEt7W4NExo0hNwcUDtUe0tcmB+G/X60r3PEQO1cQNO3FSmcyNUjojWGZRTUPL9
Gd1AfTnn11NyUOzNKBvJHwOyI8lTy3tSicrfKPc+sr8N9x1sxTIFG/TiPkzgHmfQC+9iB6a6HonZ
9BWPAu6yUKVMpS1O6Qlse1ZSFmPIzdhDJhOaLOPXCg2XqkIh1slSsHB7QZYaSz1YIwGhait8/jcN
p+JPLm1bteKKK9PxwpNh4/InXAsauE2RRflGdObfIDZlOyqXIlkoCHcttEL5JgI2sd7AgcrIhb6A
ZR13iCeG6Jrz2haUbWAeg39Q0VdKrNkWjqijsIVSvx+Y9kBvAQciDQ+T64N4mQ4/4qKvL5zD4L1c
Ls0MEeRRG8ayiLcJ+sUfch8I7mCncGqxUIsePyv9H/9CMfVDBgoXxDf35Rpvz8q2cz9e/Rk1Gch/
Z8Bb4W31leSbtBwMz24a9gxUBG1fI5w+k3FgUVQk7XPwq0wCZB8OYFdYwFEeuAw2Lpqd4FxZSaFY
meKy0oBENlPogf1XUqzJVWEYEFFLGDfqps3DyZz4+UiYjYZYbpSclDUlatxI3zY7/CHtkM+7Txpn
+FNIAcxKV/WxYPe41NUmJi0bgLPHlRFQOAOLBWS2+V9qC71w9bhHoxgrA90hq+ylrja2hQuISNWw
YEwCwwk5q5Fny/tztMt3Gfr5lya+kaMHDfdhHUfP9OSjiztGTO5rDgyB7zH8IA8CT2FqbIhRRDKK
hkoQ9WMXfKH8pA2MZHD8X380eTJFicAC1mOvXURHXsIwMtB/0dP0bh1AD5xuCN6FLMQIocGEwT0o
5iXPYeXEpVRqwcT2+8/YzKX01jufSk+COIjv8F6bD7BqsF0yi5n1R/vjMVh1/Q/XQsa0hmFUZxUP
NK3lABKt9Isawjjdz++a7Z/TWXuc7mmnbhhyt5wrOLMWXfrbbW6mwm4/uTANw53U78NvLvgDxXwB
dm18SaQypopqIv/Qc6yNJXal7BwlFE3YBa29OAvl2qG5bzChMGVyNNguokp20R3FcnhRNu9L6EJz
M42xcgoovcvzhb8sfoZEWF3eYi0l/xJo716TMW/y5oPEp0+2B4nRT0x19XleDcVxK+sAEZyLwtGS
k12k6qMDVhj4JmGUjVSaiuAyC7IHPOgYZoRt9rND6pMTa4rFGz4/UqN7TT95/SUol2VJwzVgM3ts
HtkrxgacHuWns6/FNaCCD3LNi+9LSfMJeGN7YNZt8Z8wlE0Dci1G/DL9WFJUk0bgcE+8BvpfOnUz
EGbDGArzEfU7n/ELqRwoqo1Kfav0z73qpkfU1sK01r3k1/q+Kow+7sI5MrFrmex5IjdB4GLV2rFZ
U6ApHlavi4Mn8lGkQ7Nhk3STqeaXqIefl6+tR4mciTu9hNUechSGITpvtxPzM8ij35FxNopnv/aH
RLovBxjEdt4FVz5jueCXL9Ru2uohYZ2/gXXxs5C6Gmq1+OyvR5PA490cqjzYwJv/dF9OCQHUZZ9a
ioGXaiIU1hRhPzeJfZxqa+nA0mHpgNNe0FY6BeUYh1xGMY5iIkPjMiF2jbd6b1UCdM/im+x24lHx
nza0DWaVCzeo+X2yvKBUQxLOaVdf81K5oKbOQGmy0unJ3hpGg2k/cGsKJvLTJ5RZmlqVg5ltzAUs
9gIB8uinMCmWF3JU4VekB4bObvpl1JwlRIJHkFrXHDBEOsZJZb4ueH1/yGfy+mEAApKRAlQWuf8N
EOtpokyyodxDDxlBpMXPg2I3QDrY/OU+kTCSbbSu4u/M4b3cqjdLk5ctM8Ace22Mlv+EweSGTN7z
1LSkamI2VmIL+gVYS8SSrQJXGmcg0MJNubkl1XIEsDmBnmv8nu6iA39XHScYDPBmdaBMw5LiUCly
N8J5f57OEPi8zxAkLxzpGRduHh68OYh1F2zwRtd/UpFGtZrvLpTZ73s6b1iKQumH2KyHXxUnSTVk
NhNmi87ClnjvkOstqtCEMzUCXfzLaHCuQQDsqnVTTmI2PxyR8HW6gC/vcaK6+moV1sw1xQd3cfs1
zOBWCYxT8xoDh9Ux0F6eyLfT4J5B+JQ5GVUWLSPNwu1UahHkEpblsgpc/Z0l0ou2swDtTeVtOsPB
BKlmaDf0lISanbpOtF1Gm2tPoEA8Yw66UcQRP3CtoQ4AyQ8lRzZJVIkzDuguNMid40DlKPTvdxcV
gnmxdqp5IWFqxTa8jW7hxweTnktX9MTwsVSZvrG00rB1is14DEUiMuOuBTjjbTqf0nYYOGfoUgxs
vhk+u2gcooGcC0xbcMMzhjeLvqo3Q8ML19an7YVWMizprtbx1PJhCGdsw0HSrVhhAF7Xlo31Z+aq
Xb8csjQYDMPHL9xVoheSQlkApwcRY2V+htvuBpBkta2tkiipDl01nlNVrR54t1K8b+GuCN61uOnN
BV5za9wPkKLZ4UC3KPEv0dgmNl3HnJ7EeJleXocR0Ma7Mh5AFlUO6NwhoV6BPbkZmyeFYfq/GXf5
fYGRsi6JdACAVeVIPU5OJ657ghL66KCG3w2on8qKkZ9/BSrR88YqU+lKCi283jFeDrYZuhODV8rZ
iWzrtl8x/sHfuN2C+nbIX6ts4qKUGCW26YKs9NQ0pwTPiVZHNAAob+PpCTHALO8mQAt15OK+DxsR
L2LxjHy258K22Enr/YrnxNhEYjVAnvLqyDVkV481fxMBC62WDKdcshfsGmWc80wI91sUtNsUHmZu
OcUpwe6H7g0czNq/xzqMrDU9hSsfeRqASd4t8G3/jQMI51lWC7YbcGcjz1tqX/IwmybqYInWY+UL
wnr4k/bXwhN4a168lQqaBQCLdg2+fxWZVUvcYKl87ePh1uU33X5aZP2OA0e3P0p9StQGr2gAow6c
u0NmMb0+R5YYZ2vi76xE0pWcIe0ltUt31W/QdwRfU6qkptiuyjC7hdqBsRpPoPz2qcDEzMEg+6UN
Y+q6cEqdLmmJAGuW8wVD/mCGhbR+ky0qifSIHQNv3pDVM/AmfDZqNjoJQ2ZNBh/r58Nz5r1hvEYM
Qdc3dcx3jWY9T18DjiYETUcyVaX0erlP6KA8uBPNhYLCw0WP7Gp5pTsykZb7VM9g5+2YNkOsyJxW
j85CJ1EyehEgUqMdcN18S5fZ1ncDtl26uKstemIDBk6/BDuORBnkXm7A5FqDbOyCg+hDDW0OEqvo
icyPPf3t8fy3UDnX+f4eMcUwsDO7vQY1XM++R8/WCImqoIzXkSCccFD2jcEAPdme9vANiaLPDTZI
sRzIH8qJ/CaxyEHm1ty4uV9TZdosxh0MND5jCCnHKrpGjdiuAwta2GftAFVS6ngKFANKkMvF3y24
2foAU5bCwkbzY1LL29fc6PWUWDgnFeUsC9WVbHdxFyvEfqusHuOdku4QHsqudnoIO2RQFY1oboCP
jBGsn6N9LmTIr57Fe8Dq0d68X648RgnHb3daXa9DlI2fMlI8TZR0hArnqY6RMOfn6E8UEF1BwcWT
OYor9CUWcQuxeakorsCnI2Qu0blZ9f/dbQ5eiWXoDNuUHPn56X3lAWolKFWNnvg9D4nhiYup6eYp
Sib1JzZZFXiUgbHuRN4ThX0586OTpGWt6meM1qYNApf0UTCLe2tdG76K0gjGtSBlrRUtbR0TM9GY
jWtfPKM1eh1kECOy1RCB1+3XbS6esnYGT+j7CbGmxP9NVTkjYsOo0G4JtW8lqo1F+jw25g5rUlBK
8xtSNTSw7T6gMTbIW/k7mM8B6AKql3C7/TZN6oqv0lzrMcC6AzszU5hGxxS0GL7klrXtd6TpKB+4
Fs4kAHiJDVqLC7Ylvqp5hgmB6dQk1ijCFhJR6GncTSYkO5wjItwvHuc2rQkOFUpWHSY6bIOFC3Oh
/XObUC4lKDwjWO6XmzYqCOdkQu10lOF6fKQs39gzd6Kl49JwSOfwtR4wqFQ4mz45mo52KGLuQouH
QVou62ryp1DAQf3VYTH41TprQRCndOhHZfrjAAg0GY6eAQ39iO5ARDsEjr8t2XVTjNNGOr/RwZ0w
A4qN9uYeueOAeL/CAVy/AMTK3FfCTbMKrUKY72ILDL0S09NIMSUvWZqSfsw4Eqk4YUCpn/mCKtPF
J3r1SSR+a2Kc7OhY1Ca9wHHui53LKXrcwThlL7JzBy5ggfO2pHFrE9FxSKnPxYOGoPkLZVxQDFm6
JQ25052scUbRZNe1e7nQgIVtG+2CymBuMCF9sOLKCiAmp7Wo3s+JIykq5Tytoaj22LBedCoBijtr
30daZgTe7wubBkxRuKOKdoamluI4rYm+dG+BvDxEV+l0709/I5EZz+R6ojI+XqYNMZAhaq7R2wIq
J7FHTrCI16uCTM0M1HraFS3fTUW9LuY1NIqxLkjsmKbfxT1/2P/PlSsXsiwQTJzuvfygDQnTO+Na
6y5VAIsbIvfI1/GrpCkeQglSThywf3I+5k9A7VZIT8OnU66HvAVvX7YeKp3SC1oSzYu8h2D+fL0j
mji5efk//onQhHS+u1RST3PTj2Ub8F0fb5IOCQxxV04by5NGuWeH6HLj1fGRypaF52cN6jVycIEx
CT99uC5vBv2mEoRXtKHZ9gFdiW0CHZikpctzqaVriiu1h41uzn3EQAZqvHY+OtkIPONVTePJucbz
gZMmkda4WkBlnA4pN4QX4ZlCdKHKHhJPNdLhjtvI5biwOQj0Sr8V3/phwfrbl+n6IS0LqXcof7UX
/A/6iWYvcYm3W+6KkVlsHNMQ0mfd9hQvms6OeSy8hknjxDgXzubf35JK+LU5UJr+K4pOQSbRjXXj
GN4Z67p0TM9xJxMZTp3ZxU3kNdFhYZ4NlF5zHwNk2Z9elksa09wqgO65wT1SSi/o+aN8IFfRY5J7
wsTgaps5hlWjFXNrCcLcCjxKF23XF76ImTa+E8VnKmQDW7yPqGXxIsMpEkBu1fERG3FyoBDcN/0+
PSZvSTE00yfroMA3z6Xu+iz8ocPVs7OlBlhyUlO7L263pktc7u79QI2cH3ZmOqQ+rQ6m3kWNjyP8
p5fy48P2Ycheff7rd8N6K6K2wfSq4nfutX98CfcNZjDbRpqCjlCWJK3E+64WxENqVe/Io4+ujcWg
0UjIiH7j3309XV5qyNt8I4AWc4yAo3ZlA9RggxJEhyq+4N8eyru0dz9MUSVroy8+ybPqxn9danOD
BQef6iTNbrk86qcW8Kc56/KM4LdcYXyKAQCpVVhd0eNFaCP7M11+Ip/rkcr8O9Sm+uBX5zWK5uNg
DtKvrOp0rmjdjVFcTxReHX1N5R/1yF6bzpfeJECl2Frce10tSCQYDCsVfnsKR0FigkHWpyTKoiRc
lEYwcT56GOqXdTKQo2o+b3V5AstIryLwaSjLF23Xr3YggpW4aUgZMxl3/ya8ERml172dne/AI7It
S3LUJWFxXSkBMEsNImHi3nGckyzeBm01/wgH8zrxAIE7cM+FU7zqf9mz43WLRkeBFhP/6cCctm7d
x5j4VnXS3qG0JNSpu1bT9ZhbqZhrg7ezHK+cHOIc7L6+PjtduJZGqmma4GuwdtCskZi9JNM0lA/H
ITAebVie1tDeNx0+d8tw/85rZryi5BI+6nuV+khepnakM3F+Z0lRWRaKgSGC7PRddndqbhYmVhQe
ylHwA5i0uXSwPsA9+HvfdHtFBuFQj2oLn73VWkjZRmu92qOQMYGNDuU1uXLa6gfERymDHHlnocmD
b7HmIVV9zH/S1mMiNMdOnqtZvjeeNoecT+JB8Wsqua9LNKHX1pO7HAriHhlEtelrAD0AXAcQR1um
OriSwjQXso8lTFusxHqTO2ou14GmfaHZJazPRBchDg9ulscG+lmMmaTvOe3H0qUP+EELUfyof2eX
uMm+7UFB5DFZHW1ttif5lduHQNpkLAcMeGIht07sD1vu3/2+klghasIUF3JNwMqOkJYKEIhRn1vK
I2+0Ndlh2ZHYKZLt7zu1XN1p6XFsVQXXamlNGWf1bXzbUQPg8BBwj/ALPHHrtuo2ZK5vAvfnPf+K
XzMdEC4+lVp48/tva30PuJGplwGk79z5EISIy2h8Hps2/j/Zp4cifEUw90RGeqUiCz9f1JHEjTvr
DUnOL2wcuSVkba60kJVsG/DpVf2c4JoYbwanPfY0+QIh2cAx9SsLcLktnhZUl+RFMt5HcGIAHafF
gYzGFaYa9/OkTTFSxFCxRV7Q/YWh1dnpX5gZFuG7cNRJ1HRhGsmh1tIZXGnaFuQgeIwBgodY+RpU
ftYhgJHph4KKn/MpOMkMc9Oil9lMV79EOHIHzpVWRsWIP25t+9I66zyn13sfChPjnRlueKw9RuyU
SNgJQqweCkgyt93zmc3R/4RVFKutNkgi1UZtm1+kJJge1VA9c9y/svLECYpBUiKqJ4iYwb868JqP
ZzOyofje80V+jPDeE8Vn0sZpm+sDzBSvY/u9qHQVsg6Jjat8COPRvFXeVL9VBWkxKCXw1J7KKeu2
CYlQZzq+8FIMfx+w2KuZ9f29NaPQJiV6pLtv8YdfGtlNOGaKYQQRmfjBBlwtClPxyFxyPYXzFQVe
X/2/A3f91yeqF6TN7W4iHLMjL228ZIcvm4NlLz0Ur8W45RR1aEx0WSNMHBc6iROm0pyaEzNMoVmK
qnmKI8/3V3fLSqeiWfir5P01v02xk1tAwSbHA2zfyfktYtmSLKVWoIetgqHmyARmonI+gzcrnCeX
9LtagFeV6CetYIkiSsODJ7JNm651biNYMVFyF/0VN1Y32bz+/RJcatBlpqxW0zcixVNQzMPMQTnx
mgfFCnT4t8eVavdDOZpciDYGCqrQqOqAFbgB80r/GVI/uqwB2rAhj6s9qCl0nbnsEWWibjgkY63k
g7UpUS77RumLHpPLuISpOKHVl2MAIFv+9WBOEQjoK4CQ46T98QNfLOQDd7tD96IPc9u2IQVItKGk
BQdFzFJNl2kxaAJjEPhPR0aZCvQ59PvV3/9TamtWv9yszP4m6euHNsUWFazWDANCQVjii6eHJZc1
WH4A8yhZW1oZJ6WVK0tcKLLKJsDM+Or18vLlivZH8a8U7jwpdWGIITX3EY//12c424yi3dfw2NkG
N0s4P5Wy5UgD9RE44XhrLK8hYLYrQpW0+a3LAM87g4yNq1jxL6nclM9ISwHVzc37vVUGNchsyXed
1T9GeDwRpfO7CBpcPPvJn56YXeDnho7R8+ObzG7pFrBnHkc0fi5mJGijYqTENEJ6pZbD1zQ/DZVV
DydILLSzn/ifmF1C5sKuQAkctleXrfiz9HLkVbvZ5LF+FSHLvHlszDjRUp3kyr3WzbaFS1FjyjUF
GSXKt2hrZP6ZsVZWXa4vdCCldXYezj/Zrl9Sz7NHrd+1Tj7EC34O9zTio4spQ7CKhnkqPgT55hFn
uBfJOTrsdIaAbgNyEPTkyYv/LNsGyVaG3ibFo+qMp8loJhzQVw6tG+yw1YE5Ldyi0WoQhFEZu57N
ncVIrLK/62AaQkUqMV8oGPZ79XJ8WKRkRNC4AGzpRDiRwnxWsiDfr4f/5iD33lj/hiBAkU3l+u6u
KCVP/PltmSLjxmE0HrvIAyYd3RThGBewMBSxVOlTgApzwt2HR9Q4oACj+h76ODSc031BGxzm+fok
xz5VHSPr04zihNT+tlARdP4JbxVB/7bnv+p47HZaT+JGkSl1gyAuNhvw9ZNl1CTJJlCsMAvjtDjU
JV3r60b/YUTMrjBZfhAPTwdJ3SLd7im7hN3DZRgBCSsU8IMg2J1SPtZMjEaWTznIFPOeNHBDEuiM
c7Ioes84S9TMvc7UubiHvajUjlDBiLQJfLd2vbC2GzSOreiPkjO2mP57VVvU6lR+Z8W3W8kmrUVM
0v8ho7S/Vh1QTZeekPDbd12QclDo6sW5QjV36bR56w4PC1qNpLh4PwGe5mq4fgZqd9oCJTn1GhdB
T6RNKe6oOXiPiqAna76ZQOIpROi902bN1N/4BsWXbM8qKFSS3C3vwnkKpHmsUFoI0/pGHAe9bqp5
raha+ddyOX7EelGdrpFICRnZHYGUGucwz2l1lZ/J35qBtC0wpI0ya69WWxz4jv18sKeMLb/r0dXE
g2ek/OPk9L/GGXBXVBFM4q85P6rqlXe2S9hmWOk47fUGp8BRJVuEgR3QFp2Bt6mZ4bVlSJn3gEm5
jxGSSz0BhhYPlCrRdTx+FtBU9TCED/d5IARn94S0KyfB2HVh10PrK9YJF6tqI/ntlu9DPdPsVn/1
OurOeRgbhr8YeVV2PS+BITmnCbZ/JHrb/yTvwcCpUmA7xuSVgCGbcM2sQMWPePRzmxFZMzhVPtt8
RZf9GEKkv0Q/OEcim57rkLEIhHCyf/I0/LwNf50uyFT72IwKWhbziNC92kgxB2sK2Rz9D+CP0htJ
JmrOeL2HraVGiaJauWIeoeuq0oMu7lqmHUeRVCllc+cDXNzNkxaglrkfa3Y5Bd/aCY1EKlwhdJi1
qjO5zf1q9H5JrAfM2OC85oqb5EtfxHAd8XccGuXVsT5jYNRpewzUEPVSH8zqYAcBwp5Palugd041
pgy2zzDCfJ+Vjg/a/hFa06Xpy/qo6zgpu5ePaZdBKRrs86KcstFh5HkyHt6L6HZtA5dMAt8wtgl7
aaV9TqRPPfM/d/YGBTel442RTxVlsXRg1kyeo2KtedTXBJVKDJC8F1OtXbUC/CMxdkfXNElBvcBf
5KP+xa4lMINIIHfqeNNjgo9JpdkilZveMdPjOGoe4ERxD65TLF5x3Xr3IUwzxRQRENtiVWqatrGJ
RJ0THwCpsh+xoYAm0+1hxhLMosa3dTkJF32w5Mnn2iHJDCHLqMatYnvDgUeYRWI0LYAJ70P8SleY
layKVyxwE7OKF1jGcwTnyqZcVpcQSYI6TQ1jrTP+PWmvU0oH1N16A0ZYXCkKn3W7Z8l6ID7teNYg
BEz0brQFm6yDObi4ttmkn9n13j30ZoWbMKmNeeO4BmwnvB0t1jpw9jXYjhmi/fQWihKiFjTxS6C3
OqpXGOiREOUxCoAgajVjLN1kiE6j5DSKREBNMfi710L/VCVaktJItbo2sifrQ/WEHiNgcRpbgx/J
9aTOa6KtlnZMm0SldtA0PKIyM31j/mGcQNmBrsdH1ZEYS51yP7tR7nwtHcgFk6t2luQQnZslQ8Lb
WpVO3SHzmcuhDdziHrsJLXmriKCmBgAT1kULaWpI8cm6AvZhmGNUSQWI55tSpzy/PEiW74lXcSuV
kYH+suyrD2hxJKoAVTxKKfpnkBt08UqfZg+fVAwkTyjhFeYNijbQwMJX1U4JSf9rhm8blZ4e3zDU
9faWu3KTsrOBDbJyj3SjzR1CAJUeTyouEB9XClemMeznbgPPemkJmyVg/LBjlua5vb3emhPxhWBk
ydnLIGbe46jHpijZ7OBWPwTiVd6W2Nx95KLZHZYIyWKN9FBbPQ2M3N/m4fgwjc/8bEp78fQQpTQ3
COYTPo3W3mEbNxh5xlo2gtqy/riTGTgjSaOvF1o5HsrLchEXGRDcasnigA2Zl4OzhngQCwXTgYfM
VuINZOZqvdDRWsG/IzuYcF1H1B0VOJsKlyCGfUBzICb+MIopNU8VCPVJiqeeuG2NklKgiw3vKVWy
ACngvFXYywvok68soZpDuJBdnwUpqx27Hw44rCJ56ZhEwdt14plwtWbOP4NvAEYKorq6jaGxLYP3
T3YJBVI5jkgn0CuKlGNxRBtxJR9TKQTs0AiXFnrIYyYN/9vJMpBvRG8yMNGmT1q+Qc4cCTPTg2R0
b5yRwwQfkyCCwaVtrlkHuAgWwFn/4L07vBBNYrat1HimBqqkgDT4qmELHYR/K08O5DqAU9/w3CjU
iaF79qbrBtiWJbErudpGyCOL0x4AfGLILCwboa2/79OFwgX3AyixNWSvf8DH1ovGko8kDGP589mo
0CTlte/tu1967HLn3uCof0p7qhJOFtP1td5uCtOXkBb8ieKiJ06uGZm4mr6Uu9dRSu9LCuI3OLeY
rjmxMslt8SL2G4FyDRGon9gWDz9pc13lQy5/NjZeq9QYIYsdEDHCiDsHxrgkM3klrFsq2Ahk5Wbt
GvCAIs7//YBPWHYHEURmiMK6duG4XFdjVJK5HtnhimGz/pZ0XJiKswo/pjAz+d+5YMVN0ZESFtEO
6uv+SL43oLLeZ2J8k2X/H1VyA3R5wu2IOYnXvZFIPWnk6PthyQbJc6opxX9lMck3r5YNMz1DyBva
f4MNnPmeEDP9hOVm3KNmLunLMlRP3Yf2Iiu1NKncVkqqpg58Y8WBZBG6lncnq2EB9wXNuuk0RNdi
dYJun4eYg4W+vprsKef7U5ZRVWTnq8RSCWa70pkQzJmKAHT8f7GM9y6Z0Ev0o3auyEZy+65q/fcZ
2WBO5p7sltDVQyDEIH9hsYlyp1fKPHDij5SuUX2zQaI0qSu6hhHXiftd/02yUICw2HtMzCdaTcTK
7CVIu9djbwohW9Ej2y0y1xS8xnaMudk0xO+85b85vfGlDfKhMKV9m7c6rxzPAptWvQdnseIceYvU
yOnKA5mU4J6HIHSREeHgvhth1G6y4qX3cERyEMDS5lTU3iEkxyHkvUz8A2QOmVVB6QBy0HAKEKwO
i6tMgig6nUNBr53eSm0YxShe9p+WyLoQJzuEaI/HByD/oTJSOgI9fU60+hl4Dg85SMrrHAhgyZ/y
5XJQjPfWgOVn252TjfgNO6Go1smmOUvQMR0K2phBrZQmn+C7RTZ1PoePo83NV2ApIkXrkBDvTN0w
73RQwd7M+6MVQab6iCw1uOhF97hHNTbKjkvbI1C0JIf9EpIQyW1sBPsXCVZVzvGxLz6jmmD3gQIi
1UVYuxmJPp3RuGeJxqHZUuxj7BGAmegRsicQknEuG/sikTXy3SMa7Bc7Kf8jk7o8diqgSv3UDKEC
gpco5XwDlaNVcJVVoIokN3jxCfJHhIdpUoZO4PZl5k/h1prsszZGneqsNRq/iNHSD0mfxOdPT7AT
Je1wTojyP6Hm3QpWlRYMAThhpVpSJs40LlX6HNywZlEPIfppizUsV3l6AkNbr3rO8vOVH3dNSMtW
z4hm6zYjqX8Ft/Sn6XQ+fSgBrLF0D3cMIr8ztExDYOEWTmof676YLPiha5oO7nNBs9L1feOZbKIZ
ZAiLE/b3BNSBYnYAWI/LLLgdx/WtFpJOD7wmVvM8yW5od4fIjFrw4gfh9msmMgNVRWEOZ70CFvDW
o52hXO2ky5jS1+hhhaqWJU/R+284CYulc2ew1522aOh0xJS3QJHDOezTYx4ihDiZ9CtupwAiOMpa
7HYJT16quABWxGI0VtRVhaMoVatpun1W2w9FTLLbaxiDWocXAjz3eBnm8g6MWncSxMBNWd/chyru
j800u4vFIbF9F+fhevUHt8tX66ToT0hSriC2gI0CJcddXOfeaazdQ1cIcm+Shs3zNDbDMtAxYqpm
8SfP+xBGmkH2to5ZTC89uK0dk5Wl9ZrxnQuPjWYZ8Jr2G+dQ8sV10wO3so1nvbStf8x81+EPhtxS
IPpQ6Q3UonLl6RHW87eGiaUXc7dPS7yI4VIW7mebY/uzzWJH3WfLRj+sMrWhXThiWmYdhyfIWJ1j
AFFGkrHFwrP0P66zgSimYn66nx7uocBTghu9oEdRVhxH6uFOq55B+kknzl/gaEEk+hJeHNry/qfK
tBR4D22tRvx8RVyADOGAv32hOqXotRWFZwYS8217oWIzUbGQJzj6YKcwOz6DEmMhyj7D0k1Nwopb
VoA0bnFoUgMhz0paSMAcBkdyOUlMiVhQfu6V9GxtxWy79LfhZKinKXMVjti+yWHgX4wAAb5/uto3
2t1IKm2Hj7CcC96giNPK0Z1EdD+t59uEfBQrBGWDOMCXXnv+x0kyU3LpKu7ZXsxEGkm0+XNimClv
FGabF8rzKzb+/6XDbwOIh17/el1PLaUYYThqjJ3LkyW0I0KvK3xxH4ND6Goh9zm+qlf9jB9A2qB4
L1LwgCDtIfpxzwapzct9plFsVgALCEd/vwkWWnPgpLI8MZeDqvMotq/PmMC7leZCZzuGRmzDjWum
KwuxhrACtGE9BBmmfF3r+IJMFj83jrQBH9TI377XcgITMpnUT+8SuExoeim6FXTcFxhPBAP71bet
dLXaHjnRHtd2APYSwSyPCSX3PsSYYl7WcbH9jGyUvxhOsCm+DAcQ5+TQo3rPA5Xf8HvmXhIjYdl9
mvyAyd1/9dLVazxcZ107mXrlPxcv2lk0jY0+l6sje1edRCE/07wNWYJ+5tYewqR5sAsbYxnXjOeL
SJdN51hv6cqQ8wPO4I10A8f/uUM9IdhkFI4UNNT0i1kf2b/bmUbjjc2seKN63O0KF/lEBOkT7RSz
S8vqama3V79jl7WT1qZsxwc94v3xnAO6sBWHXi5BCmg0qwrnEFJrYiN/7qo/2qH9DgZ5Ck1nZ+vm
THms0FWgprtfLyM4JeYk2JcUKkuvVF1Q8DHacB89ulS2qENSz6IDVWOYpOfad85nPJG40X8VnmiH
hOSLZKCfgS+q+/mB5OGy1Cudn/E4scrhGy8UysJJ8UVLWVixcP+Mmwt72UlEiNDCCcnSYloXYd50
o+QLrvElxXPAdhj4P7wa9zLN8F+oSb6hIsKzof+ltfsC/XofBpSYmg66r7L8S3UP/fKHxGDDE9nD
X+9FzzT5q659aseRCDUAn591DPMEH3Ny9ntHVibPhDq0dehycr6UYTfg4kettEoNAS0HVnnZdOpE
Z8KArvRQXVXaD4jVmUh6+l9xsbE5laKpU7b6Vw7DSVWdyxJwfVcUTFMDFn+d18N9KJZFs9V2PMJ4
eGYLQS6yRtg1j0pxfBZRKc5ErMX8ydy94rrprf/TAhMVszkISanIgp3jCpC5vVEpMxYu4S8+BtDQ
Q1GlMknUVAvMF9/isyVMIzYdlpzQ//RoP1y6Otfdr+F/EFSJqTyHqw8jydWhVVzwvObMDh+nMrDj
/Q1qAZne40V/WWQOfhzYfwyw/2kw/Z5BIjS8JO+JqogVrTPKjMSq5u8DXE/vb8FX+YV75jS+QO9z
iGMZ4Y20SzKHmOk79fpQnpXMB9rqa2aG99qc5mmAVSd4dw6CPFoXF7KSHFdNdkHIAeOx4gdTKxGw
pREJ3OUQ2uqCz+jHrsrkIyBUc8usF1SYZA7gmVIng1DMmtQPz8ciN5pIQbIYh1CU15zCpAhC4fl4
Z1snd+JVBZuivV5gVCBAsmL9rxYy5rNuc97Vqj10X7QzPlVRUwZ7cAs26t50g8f1ACTAmHXsSjnH
SlkPP4prVlcbqmmQx2KT148QLH51RAZxOBD0SKLMKRGtE6i2Lh8bnTdXhAI/3/7VooSCgm2Anp38
SRrkCg/yt1WqTEv9HqWz2OXEUo0t7j9R7iNiLR1/JjpShB1BEZHEam/QEouoctITT5cGr82M1i9e
s9Bn4WDRMJD1ILQIMdbglAlJXrVM96wTAhacElSytj26dlNBsqfAp0ErDclnvtzzGBh/3ImzBMTw
3xgKe1qf5QedpAZa14q4Z/gB1af9LppkZ5keMnIN8P99ni+BVNk4Q6uPYfkFwkvZZZjJVo+VOpCf
X4gfP+15jerl3Zu76QWlAVfUV1FDHHHnpZJdD4ekIXd6aYhHMHPoAx0dBgPn+zzqkgyDKTE4q2Q5
/Pi2MiQebwp79XuG2A9BB7lt/d/urX8+Tg3ud9wyzSnEHW0hbEtQytN7R5p/jHgAMNP+v0g+oW/z
AfZFrW06/OXwaT8i4qTXDZ95xPc11mQ+yh1DCX+g4DQpnr2ECbGZXzINuLAXN2nPIMNYZBHgXWFr
hG9+VeYkY+qJrtE+P/LEfBwc2r4NX0jYlf6eOA/UH4OPJwiSeYzdtcMbtrPcpt6YKaeKzqtrCJ0V
VbMVJbGIC5JGZwaM3ghP3QFCDuKoEN7BIstCGwaE1PEir4JavalXKRsfWKa4kEXzBipeM4lFQLZ5
vuVfqJZfv3I4y/MDsmv1PTt66qAfcCeqdxCHzvgqQwXVzwWQkNrgjY9xcSzXbdzRorQbqteuxARg
OhVk5SkW3D7Jf4U6okn+bgWOkpsicwlTe05rYgCg0Lj2x4WeQs0Lt0pEIXfmjF6e6KeeePAh/lP1
/GvoAOJvGJRGpd2dB+T9rhPWQh5nC3Q1KFvOXrmBt2NTTUNzIiG3rkCG2g9YbWlas5RuI4GPcm2U
sXA2FAJQL4A8mX6Jck4zUCPly+nb1MJyXz2jYjI7Bm7EO3moyW2awGcEperwSlC2fOrwUPdWRjRg
rkJ5u7iU2/43qval8lj8BG5xY8l7L2v4Inw3WAed9DOxfo0bO9p4zfYEgJ6KsTOLJaRlKwRmBZtQ
Pu4+GIF8WGcdxLpPa9Y4bOoLPmX4BlEa5Ph8/6IS3rah6PujuYrXeIsFe7wubKwRnPgy9ouwM9Iv
1oVmL507/OY/Qt6tIOZEp6Wb0tIYuaPL9z2OPjmPRznU+QpZ3AP5IZWpys3qE+PmnUid6v335uhT
JFgTjEse58uES/dzd+7sa83or1ID/og8eMbo2w4gg8eTjILPgj21pwArR3hA/7TIRqZpXr1Dcux+
qspStMIlD3kTBw8ZX4uyxSoZ6lL7NUKnzI04O12plHz5pgf8TEXg2qE36C/Gz5nCZcHf1fci8AIR
lhb+pwQNFm4zc1DqrcY6Ykdj3WN2DBKWYibFP2xKLR+zsdVAaEoYD/zyc/9ZfRgGdMsgA3WsNrw5
he4qYq+1dRBIFWKiKWafCJN66lGqloy8Bvu06GulOb+tAr4xatjsdoLD8bP41hEscAGNkiqCWEF1
vChgYc5faU6Eh55OQwPCMHqGQI0jNnm+6U6wDpIg1w3ALx3jix8/HRILCMjZTGyhMcQHW1y3a/Yl
cXp8i1JzbeSBD2uh60VkVN4L3uFCQc74nQlm2uAlUyJIXOCgwQ8NyVUKH1CWq3k4GqyXSfZ9v1Yw
LNMhP23HhlLVmFJ1W3u+3yt0S04SPPC67Vjn6GqweelsCTZ9H8vQHw2uz4rlGdR6IITqnr7NJ80r
hbEr3Re8zXtGPJrdJi+xP6EXIPOJtojD5CREvhY/mlSZIyGlbkqll4ywLgkge0phVFjeHsBqtqqx
uSV/3xn5NM0XJyhQijce2urPNgzdkXmOrqjh6XRKCHVNhXHonvc2BaViQ1wvI/2iidTAUtktg/JK
ube7J2F+jfXzveFXQwbRyssbXEBIOTr4z2LRTMW5m2DHwJ2pIDpq3dnXTerD20YX5MfdHr1e6vfj
xYLllu1JWMqqlefL5O60jVltTYcPG1N2hcxxIgDh4sf4f4zzIhCLNLl++E8JqiDZOI3w6yKIk8y6
XPpOmf/9po8gzQjhn47fovDKKWt4EdbeLq3MuRhvabjVku5Ltylx0YmL89XuKQoZ2rhAMZCAjv7v
Bpz7/3Kh9qrIpCZwsCs7rZaPmYx7OTq0EY8oVktcjWK5/ixrQ5/h3bCr53RdD2uGSzrEZE75WILq
3xFkXjAUVHiDstv8W907oIuBbP7akrsSlliHuv88WWOZATlhjYOgRJKjm7iD8YEskLKn4fdrAv1A
C4GhkzyALmH+yFZEI57zVGROV5W63WFpv3iIP8wAjNAJhero4IWkoEDKAGqxArIA4U7/KiNJuOez
pkx69yfeUSgWkwNk7+HP/u7n8rnbShOsZGUwtDxK3GoPAnsIjM1yFAF8P0v4ZATX/QbDKWtCF7xn
odwtz9ni1S6UMs/kaqnwRXUaaJzkW25GfVSa6bXVJ+TwlqJH7g6UF8sE4UKJ4ZYN3G5uajpCJxD1
z82GJdgJ8qo9LMBUza2LH2dLy6R8q/LGpGodGRJtYerl9pSx0cFHfKWtbjlBih5NdpnWIBs4ybpD
DkJS9ZjGLUH9z0jA/57PFK2/8aOULLqMBF/lexfWxCL9usKz3BPoOHdndgIm4E4RFem1uvmCOaKF
VltNaBNTvTJSgKhctgTLcABYZKb3Q2//39H4j85RLc3GCICBcgPeYH2z9u6d+llRApqxBD0acMdH
nqpzzMazKIYe0GAAsMcdQnriawRBw1100qf2e8G186kJXkQ8uz5x/5WCyitDZL+yEpr/5hcrBEYZ
GEYBRtM+ykynXIaV6oXUDMLPjH1o1OHsFdD2JxQEJOYAFyGG2ZFb0dxgqwvsQpMQ6UQGws8vVDhY
rTeYdh4+Gcq+lYd0AIuBIAfwiZUfV74Np6DdY5jGaJfbwzwQrJdY67iR0llKPO4kUxTBP36A51HZ
HofmPyY+IhFOLQ9uMbJUSFtn5fsgeb6wHNNFEddxDslFD0nmel94fV3CUaorTA6Mwc9AJrOBKbLf
KHXbJkqjbyYQ5XwG/rSjV8Exvk+2OOVlHk2V9zBww04i3MbsmScUjCWHNcfEkuIwgSNa6fGvSL1B
RgNN2ANfPElhtlBoPBwsNXC4N4RNL7mk63E75SXnrulmsKaSY++MeILRlY0fGeKX4RETCmhA1nhw
ESbNrGQdTQMfUotwAr1z2gFmg7SfbyDZjxqbxKfAPmiaohzBSXUmxO7plV3F8Yq5WGx/LZSEHB/4
ZZ8BdRF/yGRZqcvuCqkCT8kQwhTwbp+tOsfGrdWM0D4+MZIXgZ2NzsfZnv1+RfiKgKZcgQxjG27/
bqm/WP2/cpzPKPdV+gTCGa7LklsOmZEL9VxRNxSW/xtjIDM2taOx1t73Cau286hbi1TNbVKGePRD
OLVNVTgSLwDAw2/tn0gICw98QYmpgJ5hcyd3jFHfwDqelMDIYIiBUTjXkveCCDEDvYLj/tUwd7ZZ
MKwEadX+IdOfkfSLDKealB75LOi4Hq7RxibxfFONwjo+WUJ4/EdXqFdJLYfd3oN2GE+vQnP2dkLL
1SiP8+FmHnrjRIl9QPatSpG61KwlJLlTaXmYuKNbctZ6JorBgkd9oHmlMKJE7Yi/c/fHuMHcGMUT
5hwmivnbhX73pzrk0SfXSxJ7LGkN5oNWVPsWda2ckj6GCGMh+i+Fr5BOP22uU0zuQGXOKZCm4GO6
PprUQgY7BUZG3pyHxE0wlaEtCnEPDXnSL/VJiS324FqggPsMJhuK0n/droFx2b0sHg4RRJ3606z1
3TyCbpbERtnZyEPoMGuzDjJJyoRGtlyECzHqtnTwjxdplersbRlDZ1Ji3s3L/xdn0kaIGF3zvBRJ
TN663clZecYmBFqz8As9vcLlIQx1zahoD2oiJG/JEhMO0eaFFoK2zAZ5LdagaTpK9/eaj/uM8qcz
Z7qGdO2j5G6wzqZRAjlWXqHgub1sgK4L5U2d92QwpodpOD35+vzDSCMa2nXaxhVcRCswW5T5UYGD
KS5eAJLJDKoHRZAxgGEo3uAllMwNgbzdTZXX07gXueP/VcpMiPmhSjYhtwiLyvqDDHIfILQr4tGa
XnImzeTV5YPZI9P0nGOVefOWbUccedBuM+t95bqsuA1oU9jxQ48uuEKMwabJ3ZewocJCdgM3caTy
gMvLxwioFHtbxQtPMYYrLbY+m96c3OQOBJBf5AvLOm1qO+AlinN5TPZs6Ozl5rEST8pjmKjMBdri
4i0QRq6hgYvBPYjUimFNTp0x+V5E7V1bmo4ReWkkE7+t3FM8W8xJvdyCWG8C3ADxk3xxf8wv3LSq
+PHuUeCCEaa1RFve/F+t6euWL8f0V28a4kQrzsXAaFyEBFV65h6EBcffK8WUe0UCWF4j4hnPchOu
t+49Fhpkeu8Uptz5Vyt1zcvNwz1snRnL/vp0VOPlulC5D/rmLoRU8pvymjFRZAF+ob9F3vq4dzId
Lgo781b6sERKnuMzNFu2gZ3iiKmiELRtW9MgdfipyL6w61RZGnci7uILZ/M7QQee54RkEgaxThNH
GxK6k1Hi6ePZ8V40GOfGQ2Loz/Ci+wubG9ceDgxfWiRrwo4IL1XbFJNX6l5BvSE0m7nsYoGAvb/O
lBSvN1Z40gM+jMYhcGaBdOK1onm1Q90DyCi7hEL0K8oF8XEg9MTBotVqqHWutTQE2C7KKg1VbVYJ
kXFZCRbT4ve3CHbz61DoqNVNIbtxBAx+k1rRleMdcwqgeNauYocTvIjTib0KY9mpueLXCjYIgJB3
0gAUB6HXbAKxAhqRYSFMzi6lYg5ESjMCSU6QRwCzpdb34hyS8W4GMHyO3MMhJi4OsSftfmXIowjN
yqJlKLQWiGtkp8q956GQqxRdwqZw371geD8ZZ5yEufrbwPowiBm5wYO84qNUW4/hF2TzAXt+OuAU
rY2tGlXJwbCPb+nnbJfQ+At2WjH3oUC80YiptfilUN+twNRPIPq57EmcrHFhe2BTzj1GVBnSftLa
8x6DBeyNvZtPuebodZs69R7D8tecICOHzfIo1tmfTGsuZ1liovRGpDA5MDystkIAAe4J3bB6QmQa
3XJIz4SP0U+q96SrQ5MutqIiYqle7pWch1KQZqm0Q8Jd/jKvZfg6qGuUqyL9DRsMT/vQ6UxEGP/7
6gu1DoagxA3WXbaQilPfTPhRRApUXU8OxDZXB+/um3mutvQXYZtm9iq2LgTCk56p5qRde1DpaNnX
QklcfyaifKglOpqf7uUYlnJO1FcqWC4g7iVkkSqMZRrSE7Hjagdf9fLTAaHJzDH2oeqz51aVUFU9
r0AaY/rJ1d3Iyj6pdyVGuzZuvHyf9DTVtqky7A7lCDrrQLMWw/tMhy0G97EU9Ehxm8/x19SmNZ3q
7Jdn5MoLWWbuDOVaa7YREP5746ekux8EqEhsnNLlnVPKnYsJ8mzOcaaprR0yUn2pk8oU9q0TDpT+
Lw2reAiGioH46GAhNsOCugCvGp3tPCP5/aWzUfgPf9ZjO9q/0yM8vihjV0f5nPKBEgcuNh7jOMbp
ay2xSPFjLyRgC8LmYC+iL9eWlXq51pAuwoJ2uEZfVTqhx0LhZULSUpkAO8dggfWBpYk4y1lrHm0e
4fx/jKzu8DzTxSctJSQ4snPbVRDPbu6osZthsLvXM8Ohf26BR5RSooNAu5Uy6WmAQFIYcReF2Bcu
ykUfvHMFeCl/6WVUiyFafUMUwbDSkHhIdpa4NU/k0VFvTiR50qQPFvwrJI30eBtie+qVuLKMB/Kv
Vf1oUrSB83KWtZ4tBf7Xz2p5GltbLlYTF8kN1WDnp56FhGplYm6E68Jlgt9zr9xeGWgZ3yOvmrRp
1QXVeRQ95IhMwPiv7D9lmwjgn43V38giBXSE4edku3Dt5+5jTKml6cSkhMIlWiIJKfHN3HkpbN5q
Kxrz7hSDToWv7BIT41eyVnOCPUwCxTsiLm9GbJfPVUQM2ZhuumiLKViqtToLQluSTCG/wMl23vLZ
oDNQGzi9E+ItMeFLy5Bq06aSJmiJd+EZIVpz+Tsch5SP38eDV8wxNlusZzhih9sQO54hV76+/9HC
87ptb6ZTQlQutNtfxL6UsVROYc0F8AjboAHUFRV/G7Id39CvklcOpoACyLqwK44idqPOVd4EGFmW
VnEM9YWQIZECnWUHVlBiU3QHFxDq1tVCXqsnuenkMaZtCLu0FPtfWb5wZykELI93KusXalpzSbYY
epKl02fpcybbx+VTJLUEmZXhosBxulDHS8zQL8CCzBsIP3aehSt7vll0b8BkkDfz86vDHV4kEbL7
+bD73NT+MniS45HitonWA4QAmMXeShgMPiIvS8lAkaVX2fkrg2kpsp8JUXDj5NwolhU0eEi+uY5B
xnXND4S2WyYFgv2RWE7SOqVSLn0yzYwg/MBgpO2dZ0ZCQd+rvF9eLtpdOdRgqkJZGcdF2EVmIr1n
f5YHMzkoat00DOG9iLW4GrN3wQ4GdR0FhMOJdcsgKhQbjwlNwGM625d6QqblGC17SI5sG1JetKDg
ylyTdjp4vC6QeInAOPLsvv2/320KZBJ7smH6PX1eqW9KSEIr2/izEuGPdkXyBDCbQR0Az/xPLdPc
7TNfDron9Q1mRR8HTV6wbDLCMcBibgc9G+2g38033+U4w5xYqmg0HuONth1iXttGE1BPdmzpMdUj
4HYS88dbxSDw23sdzpvhYXWuIfWqpkuEjVas85c2jGC/KdgPKysSaXxLJVNqLhTdfWzXhfwth2ME
hX2RieSvysq6gSEIkevVD0S01Vzu9zE1b9ZQfCg1thQgKET7OtC7yQ7NaaUokGqnYZMpFRHAe+TR
MR2p5tcOnc5P7duyn5fNYatF4ueM6b8J1ofDAUC+DRZb7czqwQGyH5QVDxN+SvQ4G7V56nGVoxQD
vg9dpsZH/q8qYsU0X99+lVr5BmDkIFFZDlFk6xO/NIokzRzLKcA9uQlnJeZ0Ftleb1USSImsKOrA
+rhAAzROy6qVIqGv/NsNDCuFpiRojS/fIqjgZAjLzjDxyrw7FJqm7qLNJl7avpYnKMWqh6hJO+YC
NAF4U38ut+MvsOEhUrko/7U+ZlBFFKT83pAKgnL8gWBIz5NNFyLh2T6S/0Co6cxG9b4yCx28Lmqg
CKIcoXX3LO6Bq+TFlGY2Gmg6nmQ31dfZ4pkfNrl9sXJAxmPc9Xi9/xCSUZwhzJX/F4WCNWo9ISe2
7VRefGm5erbM9Ed5fFaMPs7ZH+r3Q1ko1sAaNmhPHOxPY/cKyu1G0WjLB8GmJZ0790aaP1cVXUnQ
QBjaFUljtDhSgAyZul3bSYeeqF6PrAQTiUNKe4E7FMixJzYWBsR7Z31EqfK+piaWiPPJJav633cP
IalvkaXrHtKWCCll7C6VHfrP1itoTI6/Gbv0Do7+CAmJ6gg59uVi2ntYu+h0a5j26bmkEhiJuGbM
Io66h9Muq+zQHCTb3dd9/zVEgs1Hc+tE9v4BhGNzesFG3CLns1TgrdP2Y3+wAFDvcaM+0afREowN
qxq/hnUexJKvvSe3Bc0Y1tklnOCTyNX84ttudtpgXnJysTOuSu0JaiTZhRhINaAjQTN/MgPREZsx
JLhnX4HdskEnelRi+AafnbcJyOuE0U5JvzpOTDSK3FkGhCEyEQvTtPOcM0Zw5p+6DKv5VbFWAtyz
sbq7/YVgQ7Yhy00MtUerGXQn6UxcGDh0kleotc0FvoKlcSHBZEazEoOARzu3WzfWKFyrAOZGRHPl
O4v45auX56MODYs8WXCVSeaFSpXZ/HK5OXCdGKdexv9xobDn+DzWtjozAJCsAUK106WcmayD6PAb
6QN1qSm7DBgEXsgKxMFe6fFuA2B1tWGPMY4qyfgH5AQDUia4KRY0Ija2Nrv0TGMzHTDsADlp5CJC
flfJgCBuB9yuje+D+1WBFudwTZJ4/w5gYKAz4LmNpHqE7aIbZf6W5OZf5KJF7XagURbf0OZEhIKb
wRj3Lp4i4rMbIWIwh58SWh7B7UARhLC1x07iRBxD+Mf2WHZMKeLZ6RwFl/KLAFGB/IOwQ5wdnHjd
1vAvUtQeWU0DU8gZ4AHlU3x4f1MWb2jAhA5NsyrAVMdnPzj4wjs36JMF5D3qxeQTremfzRf2Xc+Z
eETxV+BRU89Vj8pLKM5nD0yRUSnjZ1YsqGtNtVm+GgnZpu7QJ3ujfFjFuWX7e825QXCigQ5k3dxX
eyyrcGl8BB4b6WJPbJdPh9IowA+H+PZZnXx0gSYm3+joQqSWYOaF3TJt9Kzm9hEu1y9XspiMgOuc
1wXOY9SaN75n4mZjvplhEUno0pPggDYTEGTOPf/4qOkj3P6OchA6/dZpr2xRHdxyQYYQ7A5D7YrH
w9ESCvRdnckINB9jmHyLD3XiItgHRgmmbBjh8LmqGF5WghyH+Qnhsb2agdIbT12NxhAIMjDTuzJG
THj1kiUTetDnq+WSpU9h/CjzRxDHRoI5V1F6QMQ8unM+xbqmjCkWk80yv1zQ1zQWSlwohxAmGDio
QZ04jqsdvCMDDuy/S5f4WsH19SROc+kB/AAHUKzIQk8BvFdCJNp9fl0DFYrYrkFxuvCNIVTq1aRf
zqF6ZTp9EEqTuOETc6xT8DBg1GZTEoPwDx55Gfh8qS4FRQXHYam2NR1JT1Nm8q/SX13xdSbrtwVj
FLe1waq92Rd9pAQ/tehhR2bJ+J4sVg9fcEoBzDJ9/dDJWbmcusd+Ktf9P7aolhI+XhhlyyiQLhH3
uvuYbNBdN6hdEa7cRf1TKsYguFcXyFBDa2nVjpVORzBuKgMITTd6k9ncjxP3XRUuCAh/3WpcDXNC
MNgAxxfmZwzxUnHZfWrFkPXdMAszQVfy+HE8HfAiyTXzCLzJ8FsCCt55DpWZ2wE4LoRGalGZH/R+
i/p/KlJcYh1Y1rIw8hY62RH6Zx3OkfRRmXztMJFiFhOlqaW1HG2rYwO9OZgfrLfN09jK5/Ay1NtA
xNcDgz8ineCW4kYUNgaPtwg5jSpo1HBmX/9+EXLmwZ58S4Pa+tHEXd4ncd1uhYL1dkKSh01VuOjI
ZwseIaRT2jNtskhNc/TbCTGb4Y0lpKWfjTpvBC3dYb8cXhFp8eKcuU1AyPkdkX2EMAnD/6+NM0V6
NqU72Z9Du0isx58SCanFWR7gOv1RoRJ7/p70P1thj90k/aAZo5X9eEo0Wh64yNWUWDyrSghezvBz
KIsNDGHrML9X3FV/xncgjO4CANydodkCmhQEw64UodLZ2xrNXXZpDf90siB9762CyGYjoCPcfk7E
uvrKUwULHGoeUD2f0sc+9jhomumGWX1RAmJJQXVa6llhlMJ9ikF3vEaBDLbO2F3e9U7wSI5Ut5ei
slJANDCYiP5lXzO3jFhfQm6S6ShCp+10f/b/BWm1clS3eVMYFG+CNLmHDl79FXKsSp+MjH6te7p4
vFbOQdMfSstRHAVP+s2L1wPjTE60hl3innkxyuA3XYHahda0/G5boblQo3R+54An7LJkqA6bNyBN
PUNJ23N2Gb5Bp0cEWxNgIcg2RgrWUBU8B1/Kw+2ynPykmqGyPiqjRZ7cmS57dv3HTxnc5sNHpPAO
zVJQx1zHZw75zAoxB2cuWKB6JxeUjkdzoKydKbA3JJDX+u8UMN0RB6PtApRjJH4Gc3cJOT8ew9t9
acj/SSGF1OErhf8+wveJI+vDPtZYhQSWg79kaJm5WRGJxq2P9kljfGpXStiRmm3YRHQCTRMeqtLM
TQTLp0bnu6y9/jDY6CfTzw9FF10JZIcK7CaW8xJwpdbn/9e3ognc17uUFd7K8A0C9WE2IF38OLC6
ArXLmMnUob9v/gK4FnqCjCmco6D2GWUXlhjxaoOqbuEBHlu7oFJNfwH8cKMHFjovCg4ZGtVwPm3y
1z5zU72AKtSMvNKV0fBI8XvVEMvGZGcUcRVRLrS5HM6vCI+QWKfs+aGZeZmvFrg4E4DpFnM2WJan
YlX7/5YwK/kpjlbeXTprTdXdEdATbqgWoWP7a/ZGTmMFjsxe0A6E6p3E29RjM/ZqYAox9iXzWz/N
4CferJhTU9FghhJL6D92AJD3rnsFKLazsXMJjXgFp3MYvM9ktGTLPerL35jpONbke0nD2JIya/DN
V5IcVSn9qxNydORlbnr/2SqoGPveRQp/Lz+1Iz94BeWWot13tSD83SGZNZeg5LG1mqc/AO9/4+s7
XP39Yo2wn5z/ClH60vA9aQrQ7v1VDFD/GvnVPabYa7xFexHZARdmxkKcrH/OpAc1rRdGpttacmQq
AQSoZ9kk8YhJVyPOkLtqSRWrf1OzlFEqL3WQMrnJ8akaoxIk4qjIiizC2xHcGW/Yl4XiOaytT1i2
bE9ZJe2R2xRyJNvnBNT6yWbcTZHWoIYPALOnyvQZazwqSn8O+PEJzYWiqYHmJCHxzJFOgG/n1xJW
CTdGo0ICCOICkELlLY29Mnaf5AxBX18ZxW72jTKchn9u/NfbQzK4dNJXnV6Azuy+o931x9PcQ4eV
pftRrBipwncseQ7X5qIt32QxNOeUNAy1fwgne6e0AffD88s03urTidaZM7PdJHgwVW49ASG6wWkz
6Z4aa74N5R6wm43uPZKet2ge6329t6euxm6uVnPqlwjFY0wcsbvKVeb0dVQ1sCzBuZTKlGhdxp6a
oT0CBIi9KHZnCFUqT4S0QzjiTKdgH7ZLxyGZynPRuqYk7FZiLBfMxfi54EkyjZvlfQf2vir/VLql
P2jGq/5uY5rNPuc/O5D5dC62Qy+eHjG56X9zqcbHB2XsVBNUDVvZuTa3kcNCufCdxVA/Ovf5VpUP
rvtDSobD8xhInVlsdI5Yp/moI+r8IWovvFWjKjlAj3peNidRyU254w3HpOj7s21IolRsDOrLHiLK
7UM9xkvqq5BcrmU14ySx3u3E3zogxE0nukzG1uMrBvasuhVmBpOUd9P3bxbCZglM9oLSV9KK5W6q
xrxxI9d2TELA9ipUf3n8M/8rUjUoWo3kqQ7gBEt6PmKE7EFkcp3r9dG6Sg/L5srUIvs/QCeNQOem
PreVULYgdANowIB4Yun9gwEFfL0YQtfQg1JIf9fcotSHP26Xeor/rLaxL+Ir4J/DQpVc2V+mL4H2
Lmn9yMcRuHfug8ww8N2RZhq/2xKsVJoZx+ZkEePUtJHas5DXjUMxBG24uESzamD5WNvaE4FBJB22
xCpYsW6lhRblOBSWPmvShJuOPtT3y2OAXolc4UIg5Dp0FEJBEtw3/5dOGQgSAUFeLvwdrA5grvNN
B1r0YodGZqQsJRvNNcur0SNKvFvUtLEtZjtscbh9l264TYO9k2q1ihh2+bbXT1qSAXPypk/QB0Sh
kTNjr/kL5RTtJ7wiNzp9gjda5DcqTYJVX7n7mDDQv1/1Gukk6OxoZ8D+kIhxiPGUTPBz17m85Lpx
EgKGNkrfB39eMG3kB3/bRHp/en0K7OMgovXEa+TA/25Cp4KO2wcyZ5W6HPTspKBuop0CKaZzcFcB
TbQgDDgoX78qrLAFfLC00oVLI5Qa8xQN2Xx4VdNTnCtCOmDy40U91vt9csLvzD1aD+ME3oCEei6I
oyjC/fIEcO3WTgGjwQQoha0Rz7Rny5XCfp6pdzTewn0W5Dbw2lyiwbzKVBByuX0OQMERz7Ml1F+4
B5HvRU1VUE9hHjQ0wGLnTrFb+W/OEfsOwGPOgTw8wLMhWtyhIF+8Z/js0TbYXq2zTh65tNpxAXuf
LYnRIqY6u8dYmSF+oCFUx1vhu0hL9t5mdxIZLN2qbQ2UJ4ldxYWSU/fEBzE64hLggONYmvAHuOU4
3viyHC2FxlQkRTA+VBJmgQjSQ3vyK9ufbIz8y/nnIgUlch9ps4t2MUFEeJ5L/CTHAPwFb7/PT6Kg
kVhCV6w+lra+SbSHiWXvGUw2pvtHM2cSKt+bb1/F9zXk4KnD6/tgj3Bcyvqkm6uhEh4Da71Okbok
hWFbFhVS/zy0YZpYPAfwjvQPJo0m+2nYQdcd6oAIZLUuyH+XgoUJftFnUvY9NjQVSZxGJ569CsVV
+nvTbdlheU6hdfuYyzKOxyEm2EKMvVnw7Rdf0A/TiK2Mik05T+wqUahHLncyZazI+oTnA8icHDEk
LejXkRthFM+ACNHlIrNiledGsfJJuqMt/WDwIxHbieJ3U30pobIvqhlbuUD5sWIl3dnowA5EmcYC
Z281WFiSIUw7McVeuuZc0SVfTAUHrZdSyUPloi/1cZ+MYpAm6cXPq+7ptvJdM2JSbqU0sQba6kd3
0GSDIlvLkLSxEbqtDAGvjlpUjpmg6YHfDp4z2Hpr23FzrzlJI1uh2IiFrEG6+caNsGD0Ihu3YNfi
BSs0bQMgbQwgwBRpkAfjcVH8dLNfrJzjWAUPmWPjtUgXoZbab6QkL+0zo29Iol2SPlnXlFA9eyf8
UGsAOyg6C+OisLshBr5sil1koHFfBjARDICZZ8tfNB1vjd8+DDnqs4HvYWc28YwWAw023fB2tg00
n6+3riuCMoZiiUpQiyXDznlXY59ONMXBCOnZe03iScdL/z3fl2EdRIqTdzBUe8f8C07q98HHrdIf
mRDtQBUZekvKgtJpWoFMM2+juNdk4droouPXsxEGv4XMHmmG8eCXORsyk61sTztB+uSa0CIewjdT
Jke2FcLyNGKYe0BAGCzqQse/hvTndxxqNAI00qU57H8/cty5fbblbvy+gjEFQP2SLcweLUHYEyjU
LiHsf9c/Bl4e1fhnqe6K8QV0bPJ0VtXq9EdIoxALL6z2ifikJhDLTNdTNrUJeWi+3Ae51wwfVQoU
a51LjAO6W4A1JqOXdcDvDNzHWKTzVG8NJ9azjoZltVVjxwIwiz44Ph5moaXchp43XCcqUunKoke4
kW6ZTVwEPZqx7sqnlQnCc4dTqYTVMGr+xf6cHZcgR2wbZfMzwl24aVEptcDnKdSy2Mx744c4kaPv
e37HF3dW1FOX8JJCAemsAp/9ZxkEb0ofXK0versjbQnxNUcyFSwDeaMP7XJNmGCZuBZYo8wEhpe0
Ngfp+Uu5/HPi5DEveAySUp9J3EtAtXCSmsZu2SFmeYREKuQneQ/e/WaVu678rolnHmRmx6ljNT3Y
60LPc0i1+2nynq9afYodUexToI3qY+9JgfKiLlx8t7AJQ1tK7JI1JodTrh57qnj943wPWAHUWF31
efbaSNtIwSdkjRfgI4cL3nbU5Jwe8i2rkqlAspqEO4tCuWjJc4ukqrE7p2race1D/0+6PFhJ7oyy
OkRxhEa+6hLSkZxDgY5eJIxzRe3jZLgc4zS1QPWQthv0qI5lIG0XpRkQeopVkpUV4JaMOKnNKquq
To11jg3s42EPOvLYMzjJ3ruvh5+uyMHagl/WEsUjcfW77KkCEXR617HnjUV51+0ZT0gPjdOoZeT0
wHpSBKPJOOhkp5nQXdAYQoFPR7xpRx6fnj7ppPGOEI7nf41JHb0i1LWzSvxYoixbpOjPqJ4iON9R
3oc9g4q2FoPUrvZnf4yZ0wasj02fGpqHcBnol3JIuZY6L1hsf0x1iU8tAmhHDzqp9yjJBW2UYlMd
bSCfXRx7dDPM/saCdTT2KIx3xJwNeqbDV3qZLqj5Y+puN1E55xYAi/nhXMUhgosXhhArbe7J/5t0
VFsqusmMaKzZ4oXS/LyYeDINU45UWC8E29wx0UvjR0CIbxnAWC9fiAom+wqPzw/iiUFcAQX5iMkf
M/ic0jQ9k/nlG8Oe2RzlBDlfeIIHRmP+2eNMNKoQpOWDTVKel9JJX4AD6Vnq0btEsV9/9WmDaC95
0dDdCuUpJKLiUuTR5xY2udOvKPQFVN/baRthAned7pfwKV9FyvIqX6C8GIH1+9Ga3SDtmuj4sw4c
rr4s/HYZt+2rmiz8HsV8Bo+gxrPfhZ0JVsGnuLaHkskOslWzBZJX0LhpspVEay2tq9XYd/LxJouk
21F+jgFyhdhnMsdhfb/WE6fxW3GVbaARdOqaIfhR99IyDpw19DZnLqzFi/ugGXiMn3+IUnnEt5w7
lWPRNMpfUknawHavqy5n9B5TT8z+qdV/D8FCMiBaw2JuyGcUHWlCPbAlL32V6Z9piCVhwFPg/LIF
9SLRZhFtoXrKggcOTM/HC8H89jvlFoTGUbzGuI6vmyAfOdYADnIkdAS4ZbV3hScbvSq77cm/fzA7
GY/uB+6++vvR1smL4a0pUOv4p9ZD1E+Ka3fderIhJHMrsdnwvvAFfv3RvZD1xgVtTPUf1t2b+Hmb
m5M2NbJr+eDyZLoRtOYqjIRA8gNYyy7i5Lu6gWleCo2ySpOrhlLTEw5Ope2dPax3dw6Su5mXEEtx
LM+2C1vrPdPxDEh3+rLauV8viARETRjigs/921c4l7pKIzsTlswBnyQxMOJb8bcIzdQawuz09/Sv
8iCxchvJoe0x68PFoMrg76CGrDKWWD5tlM3BMo+b2xxCy1ZHjpBAvEt2trZxz5mxLk8TrEMyxiVh
Ahnwi52dwoHJI2qZIQsMJ0saw79t+CaQc6wZ5WvDydGBrMI3nV0qc7XtdU9Ua5VQyotnatqUcX97
Sz4U3xGBQH/uOHZ1FrJTy0sbwP/YFdJXZF8yQXdo1+fYIKF6deLtoPguFdu6j48J2T6xx6oysW/a
IDCNN66djFDjBB3PqiiBS80TDBRWdrZ0AljbDEfcALFaFNg0TfLbTNUUCdWU3V6zXS6+ANhi3ioD
iLl8ocTxfGBMVz7yYgXUwN+l31Alnxjz90MuWdkZ7JwBJFfLCOdRzS3YMPBxSS0IyYXm0mV1PfKZ
qUJM+29HDjbYwcZQGWBRH6mb/hedDvKUgOYQk2nKDf27346LpJ5anTe8UBNwP3PNlg2CPbZC3njV
Yf6CN36EvRGjBeas+1Q8/opxZrrGkjVFdk5bDrVE9105KgPyxoIVSvssDYyOP8TFCX36sDrcxhBX
NThBvcXYB3nGjzl7b9DKQzcXiFJBXfowhSlzf1hWkPrYk34dV/rn7vrtgb/r4d5n0SMI6HexyZpl
qXQQoY6HcO8i5A9ldZZCio7hIuLAQBXCE9lL1u39s19WahuOjTB1EAHCD46XxWXdUmUHeZoDMQrn
jDtz7Ht1J8pLtg4fmcF1+OX/aFJp5Wxqz//5Gq9tFkvshfNGI/t3CmLXRIYUpwrkxsfnnh1g4+vL
OA7Gy+2eLRSi4rCf3/ZuvCyCBKXPaBgbOFcAWeKH7cAviFRH08RFLEqIg56wyARIXJmfahUsgvOf
HdJE1f+ctr+93Y6vqUKqKGUIqNrfGBpYpr3TqtMkeHuM7QKBjuzAX0WQn0ZhyaSTenkYBltk6cMI
ZMrIPeDNYIMAQH2LBkmIIfymhxIrLingflKZ8Jkzx4bd6LsmURtrSDC0a9SQDBcXkGbKaiS6Vtzd
r+A9yJ3JKhuz770opK0/j6dGH/OX/9ZbzjvmCWqz8x2JkhzMDeA5xtRMtUl6YhRvbVpz1VlXdOqX
BkXn3ETERR/HmZtQ/ps68vdPaDuawwxRiNbEbkAbpgVVcG/QNCSY0JCzHkQF6cNz5OZSA/rTen1j
jUaD4gPBR0IyFaiZNp9Uljm5NhCRBTfGQSJqCIFaOpRhMmf+UIc6MoqEUwaSLmvZ9iItlVqWXzKM
PGQwBDrIuzYEzzlmQ4RuaXO5ReqrjU/7nT9Ad5tjE3nlsjdHQiCNFOkkxA5QlaYu1tiNF/vGOVMI
GgpxuwLdsPnYEq13Od0xqmfXwNFTH18mjKau9Bz/M2CQiKDLYgNWDhvbB1bDruR/cAI9riMinzOQ
SoJMGeLiEiVUzsGehq43aUDc0SH4TTrsvc1NO8JTPuh00GHgLk2vhRIcAl+sYmiW9hbZ0+qFFljy
eUacPqiBTo+YTSMVHdUKHKrovw5wa3YU3MQOwxseo3qGi5fjNk2fMXQT/olgknwWljyC3emEIKl9
Slk45TSWE3UEhnD5vjzpnm/PbxMljOaebklQ3GU/9zuYb6iHA21KBFw2k5TovAYsnI4Nv88LvLk9
Les68A3EhbBZRpQIr9G5VyYdEwBHvL8mLfeWVjHPv+k/ggsZpigV2IFdCJRY0fX0OhdfiHvN80YN
CaiaA1reMoGzfUVdsFaBx8gQ2Nio9U5PdZciTQBjlKYShw6v+fI122ORvajbkA2DVCSc6aNqWHjW
f383+63m01Fmy8ZJVNdoidOSBRHAy+yVcjCSgmYdmyr8OuTmXO1fZkoNLEu5n6IKQR07ZBg8/G/i
yJ3EBLCovVxnZWz4RJoxOTfl7TEhHGuhjnmowvzGJgcF1/CnQ+MZaFtMOAlHbpv263UobXu73S+b
Z3G8cVlkdozC2xwlqZutS8+OvbXfOMNQO5yuzfu8G1XIGf7z/Vvz9j2ic6WZqz85wfr0qYH5PDlI
TrgnVlzUiw9hF7f/eVm7UZN+5k8TSNjE65qL89/GgDgqL5rfL6TpOq3Hyf6p6SPg6+8o6UrPmyjg
UTsujG15gKy/wdafUbOYSpEJ3xPtEphFvHB1gFkw+O7TT0F1f2SOiRaYJMIpHUYzKUDvPhD1HR4N
iTtBCjtlVRIO7myemAjCCAqH3D/x976SnnqInftio/XMFM7hrk3S0NgCIQo+zTUJ8NiAn9BElSdi
yg/yIVpWm/m+8O8Nmq7g3m0W9kSnGlG/6GxvYbLF5AeYpBM7MZWUxW+hFbZOQ+PR+DozLzz/tlve
yaQ7JhrpqfUApyf7lF0uGZzd5wrZKhdTgSqsgv4juQ7aEocvCxNrNEnW6oQqo+3zH+v0KelOMDzP
XcFY+2dnynNAyrIkuD7tf3uSJDFBxSqxA/z2vDvQ2KarUl2qvboRG0VA7sYcWNL8qhGfnKIXXYCZ
9fUq09dj1KbINihRrNCsT4CVc+sEIbx1sPUh6VpvuRl9wErKjlqzP91+HKkUiFc0UilFH3nJFZp1
ZCM6Euy8hZ4WOXyb28UKzgfIZRSMg0D+UP3FsuDaSc2a6E5aCAuzpElLHxzln/JA8gberh4+Kog1
fBGb9wUuWIIBqUMXGnWYM71jh3HoaL7kP2e6z0qrCMp3MCChvXksNBrlwCKWyK2me4QPeZMYPAoH
Vyn3HfHIZdLjPCxcdIn8I6wAnA7Td+Cx/x0znUIEXmOu9AnxWjJabEhg6b6dd3YeN/8iqfhC8kYP
rFQPJTSmARm+cFzAfSVbDPK05LvoNK60Z+bfsqZm5W0gv+yG9woeRtMHdTismLMuI499FbZ8FG4a
pQ6Qq68kWwnPc2EHvUIEL2U0WzcPURVSX35BzhrnQWA0zNuUA3y9xJzjBeSgqe2cUwuWVCTnzX9j
i1gMTxjVJVjxP+TMeg1CvoXJMJiDZ2+Y2t0Z3SP0hPvZBIhegILh8pJaKsvrvfl9I1TwnRYjxdDD
irYxI2fk20g4bXsHmnNNebkOu3ZEXwQuO6gDU4QhyQZcrABiDwGgM/PT2eKeDomFgg1/ohPDQKgC
bPUz4oX3eVppu2oXxRk8gnUZ564iv2lO75SftfE9rGOgsu7HTLgtusmD77Gucr2+Pe0eEmpcIlpp
qG7VolU3XYqZG+SPgs78388unhWGT7U6lO/kX3AM/A96GCbEob/QN5CDecTZIZRsVCP8uxjSexbt
3xF3EmWEgMcyFuS7tgifLMlC0+ZBOpBLOTttGq6+wD83029g6ycPlSpGyh/TUdALJoqeU55fGP38
Janrv+/goCadTjixBXfmKHlpseNjGgL2FoCedk7GyML1Zwu8M4uoWptLK9Q+7of4isaazYFWvYgh
NnuzykeSMdgnES4cLjtqoatQPmuqowuLaGasXsmXvkM+eOpSc3sjHRlTgUkYY0n7nhp9EkRjsT5n
ySTPoMPYgeQz/LEV7AUCCf2hdlkdzzYmI9hXnhAsCspY0l+eveaiVYGNLCdIzWay1JOTCj7dFjzB
JL04spjy3hSL3kGvZ5trMwVHgwKchQgVof+KPPNCZQsvfmxjWXPzPhQeVY9dEr0HArQVHfRD1pDO
g5HMnUEmk4lXkmn/UZw9J9I24dEP17MsjCJnZf7OyQ7nccfWpcFLe5kKAY8Qpx9vnhDQIcmN51gY
QlsNP2tfkFV8ORyxJCQui5WPAqLuQJkxBvUy8k8qyYcvmtrzfBpJ7V+4K17+d457igtwn6NSWOio
6RU1NsWjt2UoL+Pno4wDgExuP82y3Jf/6UANmxiDWv0+ybQqb6Q4zTVlhu+0nXFfKeyoFEeurbJu
uEyplKhEROks0cY3sPsRqymjKQQpyQvls+iVyiKaILel+8rurMnrzBwIkcliW52RwMLrhzFtEw+y
X4RxrDx/5NVqL9Nv55+zmZ0XjTGCBeZPi9jpFHa5L3s9RE6zaJrR69p9oj+/uR2IE+HKPoL1CmUR
vDaz6rw7AHNDk+1BhtK1UN3kogT1w5zEv9lbRHo+NKPe36KGBs1YF77igfQiCP1CIgOfwEDXQtxn
4zTPi+VtjlgbowyF3QImO1VegcFeql4c3Q3oXEOyXVG9nJBgObSFZAZhRdNS7roUaw4wYjYBp9zx
IBZfNYrnNlVZY1lNu6yoJzX9EtNXI7ZQRcI83klZ5xiL3P2+aQBbq0mj18ethEoA0s8YwND1JPFD
WK3gkslNw3aQw1TJsfpKdB4XQ22+vg9P3x3LQJrzEpbcKYH+t2BBjy3wMMNa49OAbBncxsfpxDzy
41Yb8N0V0+bPd4I9VqAFPRe8TWAZI8AzfqFRbDIzobIMF+fFcsv0ZqkXRwsSNIn9nYStw2AxZMc8
Ol7CuSH2pUJp+06nWHS8SG4YKQ9BrguLRp4CrGf//VeI5pUq2n/AQz+740bnxrDqW82Ziss1PRcX
fgwiUPXrnMv1fUOrcCd5Th0CUc6FQmouFKHNU591+Tzfls0yCTd5papYvGBIxyNDlmeR6h75x6IT
udFiBvWnXJqz0Yt2QadAYDNEd6CgOwQEpcvlYmqe8pU4l32wfJWwoeB38SCZFgGmFkEJ37p37tAV
/K95e8SFWqyMDLlOR2HzI4pzXCKIO69fnCkNcgp5tGT4Eu0vvc5DJG7/UR5iF7Gi5AYeQjmI78qZ
o1MxJsxr30kirD2YBQHIrDkAJidDSElL6NS+TIdKkqWKYVhKa0B7R/DriW/y4lIAAf+dwPoMxhlz
idIlVhHokF7YNE3Cn2GM4BMiMtx00A98TuMOmh8DVILf6n25AOEkuETZ5930JIZMjrUg++kNXTtc
os5uHyJuAnj5iFjvPJC+0thxXlT48YIYmGMkJVS7Q/ycEeqkZjL+gRDcZLNi3JDZEJ5MG2uuPYYt
NvSEjLAMqljSyEpgQ4DsdaRCUbqeJlz19ipvH6nbhQ62unj2Uq/0n/ivvhV2v0Pz9SK2i1OIwkSC
tV5pTLK7GjwF90V3+Cpy/kj4GSmtBQ9YjV4P7gfw2OsD148qZeAkvgOsqYttFJIisH1zVEb8PgTM
TfrrZK6yCSX3GkoGq21/1CZQEsxrhuXTcFSEOaJLf69xOKGcHEsfkoYW/6mBL8I+2tYg3zxPYAKr
ywY+T1WF2yKFzTNE5aYTwASFk/7DUCz+fqzQt6mzcJLEvfyRigZz68wGDrxYhqJsXRS2QIJjvxmS
FacdJoWm+5jushva+9Rzq8UEHjNrvrjHP8d2h67ut7n/8V/P7srMf+0HHPmpafh9J1nFhuy+zllc
ljZs0a8qZTpn8e8jL9xbm6XvRjf1ST0je/1L9MZGZzN3/iJvErdZfDoW2QF6LnNX0qUgtp8VlGtz
PMySWZryYDQkUO28gT5t0X0YR9Y22ldgH3bHsiWATfWb9A5PvTTXm5AV4BnOkvu5FrgjK3TaBlGQ
bO3OfoKMAYCTS5huSy/fBFegkKvDkrkYz7VezIH5yfYtY4nlFfy1a+nqMGysWlxdMeQ8U3m1ZOd1
atMfWMnmfBRnwemXwJKKsRrY95hWhx79CrOF6IiAH91CYyN9tw67bcyk5Jtf6Zch5TbkdFXANR5e
OK/x1Gk7Ds0hQAtr5y8gPJFbp+ArMd27KOqd1viFImGJpLTVT/VqlKyesjZo86UtuuyCm5zI/SDo
oZ5RRQdNYM3uPvcYsrWxc0FsqIy5z3ZPxlS13ZNyABeXdEfAjii7bnMl2ev4/LqkpMpgkRQg6oQB
3x74hhEamYnvwsM7SeTZeEXuCDeWPzsvrC0R50nmdPCjTSb9Wzxj2ASzFEnGHacJyFDqlFwBR+Dh
WH1xIEMJUEdkUwGzO4sc3o3hPHey3kzdyErVgRj/oIHgW/lBrTd/srH603ij2W6RjA+d9S4wXXt6
2GVMQpz9Tn2ZeWAYkD/Q/5w5L97vDGhkVUDcbvQz08ASxKp3jIef2vFnIAnA45ojG75c/rbuRimK
7qC5d1pykgb+7prnmLOQQMXqcQ/r3Gn7gStoQuOhRDbMUmGfTS/R1WVca8VENIhccUaYsq3v4fx0
uzC048h9gFKrwP+Zsq/8UnlPgJN6fftHDvb5vIsRIX2RQnk9IHTElXtE/G2v2mov9GPktjz1ZgKb
qF2NFL0tChJXtZxezRGHQoaDZa8vQWmiBfTNuzlhq4V3w4SoMJH3Q9iIF0AZZKOHoaaQWNx7wDaT
PFPImTFblX8oftoaxvUzQUORQuRWg3M9l6wG78B+CM2YWIKRfyjaCy9/jDtCSsrK0UsM6f2Lclt4
dz2Puxka1MWUTeKHb5vv3MbBIBeSRW9zd0f70lygTh8j1QvNBr5GI/gy9RivLUas7w5LVAF1oajf
agNTY9+nFKuQ7ipMcUjbpaw+pE6ZoUD3p4r2p+s6PZAAbZiyDrSdjp7/oGfmxM7mYgxMEaILxCdU
r2yCUnfMmYZhRdPYEtelLyrclZQi+kPoJ/lWtKe/6rDvZhNhcWQL/nOij5tzLLZJwQ8aoIN9Esol
BjS3FbgaBa2z+aTvmbEHuQaObncNSCJ8YevF8+rF62/Ut1wDkGle8R9aetZhoqfG4hXft5IP5jFp
JPho/ovJD42t7J8IbRLAlWF3YDy1nbLPKxllpWZXWqvknFQ80X3tdLsvxqRcDyus1Xy7v4GmzpAP
kWVEdX3w4NMoR2CeMpCKGXYddE556kH8UYm5Cy/96POxN7GH5qKEghm9U1RlbO3/q3hQEQ3SXvyr
/YknNDVSa7hglCZtbOKLsebmkuEgYDtXMhV1fRhbrvxdhbvvAlLvp9YejnIZq21eXgsBc4DkSNt+
TDe1vpGqzkgG5fuEWiQEfolLkszH1i4n9bHr2MegUNtNAnypuI8Zkvx3f6k4ojU1dVP0LRF0k+Zv
QFyhv41Kv2Et6AcLGOoRNSPmpvj5BMyzb8qdPfmhMgBRBD+46PvLfKQahmNGbwOjMzwVJZvrTTjI
1zLZzEJPDrDld7NXMoWU5709Gv3Cwa+KEHyZM+FRuYdVNXvOz1dNIjGplEV02jzg+P+6k38kv17g
Au+TmKRYkU+6Y/zHO7abfhDpBWSjwdvGLuoMEJXpMBE2zlgCB1EhhxPHnzn3XEKeEWVS1vq55i18
keoekEfwnAK0Zor1GE2xx/slsBfrGO28eOzNeykwxZ1MgFXnqEbtVTJMlfCTvQWkviNjcK0Rv/KC
5aiVcA8sXHFSpRaho8VOaZR7z5l2XzXqyaJro8L3RdYctmJAg2EDdxsS7n1c7uSeoDhMtBe+0VS9
hn71jzcQqPWsMEG7hnh/v84lO2Vt9Mmv4rKQ3zD4MHpmSVTsDn/8rismMDSkDl1KeGZM0+lmH0Ra
Hpb2u7Bgs/s0xZ8OnwIL53ptPJ3RO+nLFpYOw7RORCZpS5//xtxhPX1F1Wr1EkFVKjvY7YUjPhG8
9M+CXRvN++56QLSdjieT8QI=
`protect end_protected
