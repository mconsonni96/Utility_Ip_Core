`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
N3kFScdcJ1y+3X/DlQVjIuKov1bOE7RCYjWzVsXlq/ndfcb6zy3unz2zKmbPJcaBmzkkrzWmHuup
xLUhpZfecmElpEqlV4rmitDpIyozscTbFgmQCZ/18XSpqhVUJkagqrDxnzA84bavP9jWR99CUpew
MXUj0f6R+/zmJd3AUFkW34+1Hl9OEeb2rIlXuW14o1kQAx3fD1dwutuxUoc5qbEKdqaUdJM97WW4
9RiwciOLGDNBpMp8NwnD6K1nMtMHNnMMKpgSILF+6y2N3X6Y0PCaj5765I43I86JFCtfgl778jVH
ClFCxJLzRfnrPPA/CimoGMhIdD33rQR9KPP6Zw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="xkFbXToUY7aOtByZX9Rrh9RPTEc5tDtEkF29dkKDEIY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18368)
`protect data_block
UJDt+CBooJ05DS21q2tNnoGIaoQwqPK/Wh/H6VBvwKrn7SBqRA9oF4tlljNfSyi+vrzcQobGDmbq
plqQFrJCVUUJGp2IB1HZkPv8aMp0HV/teiQM8SEgf++tDOg+Z68YZdGts6gJADaHqRkMz+Kpxbue
ysIRM2eWXkS2BlXRsU0RziPzqWbQGPBDea++L+k6JIsN2XH5yP8Y05vP/a5uiLoOoIuz++4Wb4VG
rlX/e/IRypZRg25q0QDLjCo5RL2TnXbJVOyUv1+FPytN5Eyl+DZz7B5owH1Ag/A8XgY0xlKYjpM4
D0cOZYL7zuYGpPFe2jyvfj6QNMj5bzcjMsTnvu3zQXKbSjCcfnGz8Nxtf517MY2Z5aNsfT+Pdpjq
CybKVvdhXsb/1ywqQOcda29OYLibuirHG/VitLIggprqMryX7R70475CEthjZ0yLDYzCfxrZrwy/
g76YKnJpG94IIrM6UlvFwNbtfMw3feqozo2gROMaWGp8HWpkDHtMGkTKvwxGsFWGt7YBue9zxd5S
deEeViG6tgjemLipZ0NiKKyBLPMIrW9JWXZ5sM0vhNMGEXO8luNxgjhQi7Adq6Emw5FXNj+0sWUB
f6tJcQPfSz0U9CB1AqaB694oxQ4AtNgnHtgnaeCtnmCOtNJ/9MWqHG0AM7+vTt8z+TCrxgyFrZ47
QOXNHKmnhoxaWvDCvCPo13BWCr/aSJXdFwIdUNce34/t1y4kIm0dhFI1EGt6T+nPYcG/0z6jIZu7
+JXN7gmLCUYapIhDCoTGvIsy33zxruXFFB5bm2A5E+97FZWq9FMpfUdK/V04RhnRcoxxxr1tdHX2
+m/PdVezJARE/uBqq/fUfLY3SmA+c9pAZCZbF1c3xhOuold2NeFL9b18oGFE5xQV8NWEZ/P5qrYe
IzJqQW8qPOiju9i4shdNCABHCxEGzQYAb2jrbG5F9IfC4UziLXZ3bG043KnaIrufq6g7WTXIHx28
l2dHHK9+CerMr/MYlFZuFkoeEy4y80+WC3RLo1UitJAcBAtDniuY/ZVoE/X0/bD4JVyzvRxg2ISY
4ScCp0P4jAUynokNEdKtkMSQjD8Op7U+hazFPKwfX8mEH384UyfcjExC1b/AkveffTiqqZXVsB+Y
ce3DNT5mxs64st7p9rz2nN1ySbedojXL1DmZImfZbxB417Eh5A+fZ7/LLIShLZLosbQwr9a0AfwZ
MhOJ1hRd+JCHeGNrx7Oej67H9CpN7+7wppjEB5fIYTGr68vrICNkx9t6x6L3BHLnthESGA9+2RMP
M3CbzhFSEW+sZCILttKO7zUcQ7XtStEotyC7JR9rwBxhyTwGE5Cly8bY2Vlie/4rgCwFkeGDmIdo
MpaIuCKNLy59vzV2HKxhiBkxg3zFuqxK2WMo1CNhh9OFXLZk5DVfXQszOVP0z+tp8nq7mfVvUWuI
k31tmwT7CQE8apVDWEd0w62hNX3WfY1BJBkJiGEB8A7FVjyVlSYabqNpcQaGlSi5IfPMBNEfBxUG
+YaMgfKS97xIVyB6210GlO0fSv8oxlSJXH0nraBIrW2sWAbDAHE+Y/y55XScL5VThrGp2awuAZ4D
8r4GSUn8rW5xDwOpSMJ2Cp65GyAUJZRtfzY55GLRUb72zvXbCmfNWyNIyQtNVVUisVILNmBzNs1F
J/Vhouwl5FYJ1rQOJbhM7UjMEj1uQMlAhqwn3IG3wlnBJXfjGU7NpabN3hqr5YOIKxDhv8xqsoOv
bZG3HXn0aI9q6u20NtdFwVaZDmPqn/6AvxZ3vOwr1E6ypx9IyNgovH8EgLz0aXmV2liMbI+FF/4p
mSJr2h1h3Od6bJXyJQdpmYxaimI5OlBL4Z5aszklXEZVyR4oNIzMX7bDY4EBLSZomydhIVRxiWhy
sZr6eSI5RWFL6L3PUqxt3/d6dUNywjUrGvD5St140icy2FhIjNFiooIG4KhF4r+uVjLhl8VOcMVL
7IKxMDsDcj3QjBicQgtGyTbUr5NJBS7PIsXu7O+iv7sIVU0I2ayfzBX/4ex/Ez3oNUwFruobIniI
1jz8eKzGwZl/0lYVzeXCg/+0pwyVbDWQfksywMYvie7VTv5wrl6q4FNN/5z21rfaZz+RNQts3QVb
ucGFdKUqjL4AON1M2N9RI0MVOaijeyjP3eE7wE9HpxEc+De2ZsFnfaQQk9aTu7GvLW0V8NAtCcOl
krTRdvNdwvRAqa4z6rfg/W0DXzTG1h8HCAeKWx9EDW+JKrVRqYYfrG1yi5eXL6qQw43KtyS49iiO
+gJ9sJ9yTS3+CdMSYrx/Gv+4Gy5Jpg45yNkXMm/Z+8tN9USxEujZIyEY0gG9kMmlevTG5LU2tour
moERXbWRbVQVTNa22WprrPfo/+znTsE6JsuK4iL6HV8liDqg1lVCtROe9xSi+wHFXUcjjdiGVpMx
9dO1bVFYbYcHSBHrKyTQWEvdF5mLd30ZtdZVwGgFAZVphLq5xSxbb7CK13KyEYPx3MJyQj7IlcdV
/cy5tuLMoelj8RbdJx9m7JHap621trjED7jZ+h24EldJl6J64jhBwoHWdVxWWQE4wiAbL9wH3H1C
1A4AGsamR/SIfEvtxgqxeVJtHPVmU3CPIF/TJiNEISFC4V8ZWPAzGhOd0nOxF85DC3J5f77ibWUQ
lX5bDDgwAYkC1LnjsKGpLqQRK5O6U5eJmllz5VgHUW6Qn8/VG8HW139YHsLABcseLhsPt7DiyMXr
PvrD9yGkpYnE+rlVGoyItS3ll33f7oRsfMaA6srKffPZrNnkhE4b5rBZ+SbUQCYuldhduN/oHENx
ElwrWTdkeDhlZandIy/Dmr+X0P3pmSQ/hilwb847sFymgM0as5hpCL/YUKs79gLWR4qBBCO+/oJN
O+B537lMm60Ng/rF2hVS5J81gz2pfjBodbwFAbaHNg0At8yuCNS116RIR3v9Yf5U+JoRoAV9vnNc
QWUgJbu0Sy3dtyvOqilUjqKiYfUiZ1ub2HCMbpORb97DeQvIcRjegbp3QwNxtPyiQTUpNstfwbkV
jpq9H16FTMJ+tRP3CniHLjD5/h1B+MJ59+AcCpFinbQVP3eTj44OYmucgxTVH2FMHShX10bpPp0K
BkC+fewBvSAdSqT2iLUGFHddMjdDbw+zhI0rGW6BJVgJYd58d6nhCtJ41jQsz39W9DQZFx/6SlMd
6ntokarKpcvxYTGxvX0lCliiWVeX9yH0g0cFq/3ndKCbEdvZeFRwh5meH7Maqho0NoWJrHmMno8l
4ZlHN2HeTjKVS6TsYUlESLtn5A48TFmC2TQGsvG4/TEYfGf52mhCkYdpuzJsKIx29cwOOG5CYmBf
hvWdGP4aP9/gLWnrG+df7vocXqzkoaI67ZMMeGljtt0VY/7EJUysSV8huCWuymUNSBRB2Ocw1DvT
6mE3eXBYK2+Xx/OGEu6Nb3wsRg9NA4dRIU1xgPXxmLO8Ln58jPYvcA3rE92AtogeQRxqQpmVwkYY
VSkqSV2r5Oqmf1KcVMTnQ23aPmWWUJwQTTJXeBdNpuQUA9Mh5ae+E7laOsILxGJu4ESoAqT4Mr1G
1gs3tSuBQHJYN24Qz4IA+y2DAvn1Zhl6sWbzMDKc4aqMFzvcH/i38xAudSgFgezjAQwm8bLQ0I3+
k2fjzA4f7dd1JK3O0El2BgM6lG2pSn8QMNuG+FQXzTh6FnCq659h3O6dJb8Z47UalgXNgGRvuZpZ
YGGy6W+r6LPnyl0Ncr5LPFBoKpr0RwyTaMrdVhwmzyPRNf095VwxTtEixmPvUaaia+4U+2bd27z2
QmWaV7dMEbged9MYXsq17IzN85zW4P/dOXjGb5WmU46C9ldwD6tWW7tzOFsQm+vCbQr0p+iiANyW
9IeQDQ7bln7JTwn7gbE8QC3YkahwNPf1QIzuecCIsdtirGoqlikKmCPI+dez7H7AwRnUD11YMEqn
iUdIoVWtikrYpbsxVvaPWki91t2q+gpZxu0BmUpsv5WdNd7Q9ko/loHZH8I83YkEI1epElItpnG4
p4LV4WrYUvk59ipCkhR0Xf9R7lXNPrHcbLBHTdtb7KHGGDK8Xd2HseupqDjPV9wa99JIaKrPAZGi
QdxR8EMWzx69dAIM2YgytzTFvRHzIEP649klBHn2Jb/cF56PDcwnH+PHqhNzfnq/VaOjKE5QCtDu
TKgRDxDUx0Z12UfNj9+ncvXKBvS5/lTptQw2FNta+VkchMvleSeqVitbHu9TxBIQiQ7pEYVjkbYn
FCdguyul3bC/dPMHc6FK91ezCQ9s1U9T0Oqlq6rjZMJ0cFtU4SwxmUASqrmBKuG2aVm7gNa7iRVs
jCaLBF7044scsv4dNWevlwRDiit/XnCi3Kc4peKqVGh6OX5+SllsqrJ0aGhZSp1hvAJ3oHrMvyiv
8nnQcDhkqO28HL0d0amBHt7z0GOSZusbbSabtXXjMbobeAKK5Cn7w7ZW/1bWuXi0aHOWsYH96aJX
oS0EeSONjKR/SNbxFs99xPj5a816jiixdjo3WEVDpSwBJQa5++Nvw2oQNSVYvPVGy5HYkOx7VqAq
DmCCbr1ErJ+RRHyrwEc9NQ+MUHqAryfraijWUquxWQ2ontQYP68mzXxtsbgy7YyVd0kXDm28fXxR
AnNXNpsSPkf6/fVfWpdSoi+nzDUzoGrt0L3fWAad8nvAICRSL8vr82f6CCCZTpC4/9XMmdHWFZZJ
h/b8btTiZw0KPObOV+fBiU3tjF7LRjSfSe02leAHakjq81yvlnAiOW0BF5ueCMWTatGM+XkmZSQ5
wkwEn6FayG74EQcSgvALHxkn5RTAlMHRvrOGa+U0Mn7K4bwi8ZMYsNm6WM1KCKcXN5ME8nnD+jcI
moc86oGS/v4IWNm8rlTXMDbI5IbknJTi8SfU1MnTuOBbmMvz6L8cC3++qrvVfdbRPsr6Zl6ud+Qw
tW54UFvMvJGVB2Zji7hk/9rYT0ef/Cwba4SkTtFWpbWTG4iWVCgnBt9Thks+ZU/59/1PqdMOWYGC
tk25tlNRG7t8lojl/dTzSLBwOD2Nn6ez9Gj7lV2zBunX5OQEw+P1/YXF14OWiQS3Q5z4RDPMBi2+
10exVcfZjBPR/8JnG0zrz0uq6JvMMO8JHuQEH36HMbtsyb6YetDMmq62XfITuxouGVLDvYKQN/I1
IAjIlWCgTbBtdrtrVJV3uyI53uc9FOVcMi+/J4XWYbS7mg+TYkoNM3RhVP3QJ6TxhZeMPs3o2RVN
YjfNbTtXSDd52J/q3weq5sN7kElVcoWiCtqju2MBH6GVvXCKNkfqwD9cKuXHqPjwlvIHHe/ghctP
95vitScgYW11eyleFrjbXN8hPmMkW0MR2tHGyaFxlP8cmMwG1I/KFE5HQ7Tb8fThDuTJsNFykYW0
8fitvTS6Nl7vmfDd/GZKOyKPrNnCxwPs5YcYmwW4CWC2NOAfpnfe03yl3QGfuJmWqrVWAwGNe5ol
kSr/5dRBLM9PbF+dl8m4NruzNz1GCiZbVkRzbUuMQ/8qyq4BGP9GOOffDmdi1+hX98J6aDXSNjKF
BHjXopQ2LXf6AXRPQrxzhYwJKl0wH+sqIn6pz5E/b2mQ7KLLLzY/3FMoY8An9aEM74wDFswPcswU
q/YdJiLAsg2U5CPjd7zgk0FzoAgLboR5wHZQjQicZ5hrbOH10e88suDZFuqLtE4XeEwlhK3vRb5b
n4R1qsmr3pbLbSqWP22qpdVXVoRJnHoTOolnLxrXJUqmIbY35eTDkRHLktsdZfAgqnTxoEXwTomH
x7D3bqCH9Y1U0+VuaJKWlviSsI6KrykZvni2UzEJHRi3iWmSCuAf9xvxJ8KhO5SmqVieM5+Kj1Bq
faDKJBwH503lJTVk5seUZEP9ZICiGV8DXkv1+2JqYiMJ5B2ZJYiVOOMLpWI+a4auOSjDWZlV0hNB
HZKYh/jo5U0u5P3CvLxTdTY9mk+pnX5RXi3TrL5AxDWQjSmuFtGXuuSqStBM0UELTP3Rnc7d6X4n
JJZmpSQq53IOjj9XuRySnPXTgCT53iHxJd9H5iHojITlo1AvO85CD5PockRtZP7a41MId25FpSKj
QdrK/AybMqXbTImM60lGUT0raFOdPJEn3sY2ktHMmEKaOVQfRA/mWHmocx8LZ9+FbGpQ4ASWD755
+3VvoSf5Mhv/bhZv70NJTgdCsM9t9fjBgahBqgin1V5uCzBGV6e4pLzbcWYxmtfGPFFpbw5I0PQa
AKa0P4+Johi77YTTJHOfBz332NzP4fb2H07q47RbAcFBSxsdcCJgLfzOwrosPgNPgNccDLT/998+
hdboO/4C8JkDWV2tmPLRoQvZG/aO0U8yZRXFD4mcLkjmofK3+9u7ZKW/KNT4GHANMqNtV0rMY/m5
DrJp7dPoM2+2Usj4uLLJ/40Iag8+7USI9j22Gd+rqnQSfQgL5IlYh1pPUd6YrLldsHioJpPYVF6R
7HF/5texd0obkRMDvVShcWQGEPygX9M3cCKuq0I3R7ZgKe3bnKrlauv07lmRX/NXCzoaXT9oDLl6
ygbkh1Llk/ZDiIVe8G9TKcR6Yqzkjl244OHSlTygb/I6VTm6naJyntjE7fvMRQUfqjf8c3vmNtkk
Ayr3AGH2OggxigvJL+n4ZbD5HWZOmP7lMERlEntMTWb6R2LDrBXsohOREwZ0DIpwIY/JhdKANVfc
qfdiCsg46qnG4YiJUZX0IV3ESc4e8Rac90a1IVpy7bzYN/VzVg3j9XwzubwH7gGQ3ZFsbPSJbsGV
2RW/8aLhK/kni/8mtikFofbRC8puChPEthlW+xPrUoj2azGxOD/UTNUmTdPd8qAzER/rSdvKGETJ
U1b6KKo7y+PD/9wjiK6LMaoA1HQSeHiBZmdvDCKy3J5MgofV+A9gVfmbIa8hMG6NeVaa6/2cAv8z
WpZo8QIavbSAGQcww+0HIhpUab/YIhzOsS3gfOOyANCCKdX65crYcSWUGFLeTWldX0FKh53m86Qg
I+2nqBixarvAD4RC0RrTUgGLIpk2ij/euGnIsNNwA0RXY7z8qB6IrGsNSUkkRvtTYUYEE7FC869G
Jf80gJRrG8VXFH9p1JrjAPErymO2KKO/MQ+mnJ6AsXnKyHd0xpefqzCf5DECxhtX69cyktcNDaVJ
H9mJIif+OV20PSoj+D4umvtGl/w0Z4bK9hR7R3ZLxJgsnnLzZD5jgS+ejP2lOXxDCfvzuugojq9W
TjZYml7KGhZqszKYDzsBH86CVsUQM36P4L/rMdNwBxoxopTTANMC//JMKV31iqZ/Kgo12BahRwAx
1e0uAnK2iotYyyXmnw78AvZncDuR/Jah2m8/BDsjHP7vmgb+FT8PI8TUoR9L24iwXn8hHi2GIbpN
M10YwN3khkPwVuaxawOgmCKkpvSiBdc32pHSFEWDCEVSzvGNQq6gbD4O87LCX/4+ifY48h+TikLX
xlQ+e5ABXa38mdUfY9k9jaH5oSDHDbEh4d82f5vejLYWx7walalZxALmBTqg+3dBNm/mMZmY1768
TLqCmxq58+rUAnqV89ul3LDyor48FbNFOYlL73sEt0/v8kqsOvkwYKMS+CCLvFCKpUsEtFBRm1vr
Tp07jRKVb0CBC5P3AvQOA8hFQdRlTibdVryStkQEmJ+mCpkVs9mPatsdcbtBUfpqVkjmIpLhTWgh
L5tfWSxISlxvrLjWqfQE+r3S+LG4NCY1Cx2kqnxku6Uxq9JvPsxNfLzfNfKiXF2tUoJA0zrg5kcB
wvc8/OEvPY2EP53mhvJo+Gx+yVjoomWJIITEB5qmv6HeJUXkPfS60ruCPXg8SGWjQxwkg+iLsuXO
pTQAUJgZHA5HlkiSjvE6Saz2RisQXxdmVAiu2VNF+gWdCl3wXzG9Qy9QbVe8vSjDMyIb2XM1mcxn
0ZmeMeBQ4FS429diQQ5xDfynV9m/QpfiQzZ+ssdxKj1GdhXUBXfStKo8vJxIz3JEKnFow3stCnQE
/8PpjSz8QsFKCD98GnKFuD8KicVC8znFUkgR88nYyOeiM0Ki+PD3N7o726gvOhIk9/UZmKkpYalF
C/f96I6SJ0wE+f7N3OZdzslQXC/ykcTsFSFo1w6wjimzoh0Zq7OsdWtNPkqA9Ms2sNFpnGBVJGFX
vjI59A5zPGXtmoG+XV9QsUT5GzLA9oNo9E308/qyvMaaSz877BiW2+sAAn3nfL6wDcTLctZLWDg+
gBXxq3x+TmHyYGpryA60bIVs30y1+pyh+j2cBFPukEuV3aaJrGx7Rj/MgtaRSdz2P5HgLiiKH8bG
pUQixteko7qw/6mVtlyRnrHt0rrSIS89rBw8NR+UQUcFv2yD2gXPLRScS5TRFBCGvsbUWnN5WABJ
N0alf8xt6tc+Fh/4m/sdLKANzdYJwZQ5aFVgxE/iM//Gwlp/zElyCTrjk2J/MotSNV66Ru1lAgsA
a+BPvrsnQbELt/slqBvcaKydf2EX5PnXpnvUi1L3kJZe6B0THkoV4eIkCoRaxUem7uZgjR+R6UNC
iPlKrwOXWwMeIPb6PCysz/uiYfz2uByXlZVxwxmXJqFxC85XldtLamGY6M0VQNQLFDOSE4nAvsIt
WWOcJWaZEqtwQz3auK4wJY+Hdg468X8G+BKs53mjiU1UMYmWOKO0FaPSy91XR4zZOMATMAZV4SNo
ia4XZ/UuB3OXoEm3CoNhOtFwGValGCqs5E47nAhc0ybKW7mYSMt2Fn/dGlKYRieDWNJFETG/W4iV
35H/mgaTJgIdxBQphi9dhNbDpzMD0WzulWtPreY135AfeaFrUMjOHpkQWoXXl0PCgBBqcBQrUTRo
nv9dHaDXY9uO1MKbfE/ZLTV+M1lijAHXE3zvwpNuVO4MtFJgB/F+sWAHLeqv3BgSulII3qCEsCgE
3OcN0KAjLvXZAvJSgbyS7JTk8fgHm6XSohri/K4Ie7ji79SqjseOZNHh+uX+pGxe9QRSmWZ8cKpV
DdBOhgNY+6giUd3EJr8P1Vf/xfdCdq2AN0tfRi1yYhWPD005j7GVKaLhjyxQlukpdlkZXSwGBLw0
EDeJ+vPuKmYeBXQYD74D5Ka54X3M2lbZejyiBZUZ2wiPkrKqNpyBmnWz0lKYEmEFMrFRUgSpvyTh
UCWAsllQfzd09Uq5JYJlptkVTAl+5heWq1l8L7HCd7inTzwHw4OAl6WEo4N29oZHQBO5O2B+IFEs
GyMfrsFakbSu2PY2YTKbgILisE6b4JJkAxf5KJqFxhDsxzjMQMU+zEo5yJZlBOXf4SZmtWnBh3Uv
7Eq+t+ceeDAybko0ytQX0tcX3Xy5B32Y+4ADivSveHowOmnxspVvi+f5dmbTQp4gk0/tdnOYlToT
y3f9VMVKxeqhC3K+lYGWMtBFVT0vxq7pl7bUQXJPWzSJfnlh0ai5SpKOZyDjYNLqsRe0b7F/gaBB
/l2rhj54HZpkABfu+MGXh6mbECS1dnobW4naopN5hShs6g6rcUVjahnc2BDzOeI68tZiOrkknYxS
DD93K0GmeYPYlqB/pFErv1HPkQvark/m9eTLUMPWIJIQ4LH+79IDCtXRKXd4n/QMyrnj1PH71i2M
ANf1wU9P8gHZq3/u97crPxsSqvmVLKArMzKMLhYI64vRNNFbwiuuTrghuPa2EQFThw3NDwrmwteb
5FkWkuMySaUnhIO+TUp4xDqzq52eTdsmSquMMyHpewhwubz7egOxw/EjGGnNNZvnaHwCw6kXk0dv
frZNL+So2DtZJ6Ma1/W8K0iPvs4rPAUVTLtoMD03dweA5yJNxU4IgeBBPrPDXJFcI55bWQe1/yzn
HPslr3nHxn8Tp5y2kcyTBH23BKPHlJpjQ9Mc27y5HrfmA6PtaAuPjYVH7CXAByinz8YflhcUxp7j
H6g0uj7Cuo7innIkKso0qSmgAoivQjKNU3dc7GmTqUdai1PrBzrz9rjxAXsf021pY/0v4aCYt922
OKZy5mGF2yAPJ42hGvGPHpY2niVBdcHOs2IAGDk47stlR/SyKkUOJiGb6sFgD1Q5m3H9dagPIWPg
fmWgYHT6u3FDZkvQOfgrH3f/oaTl5i0m/WwiOxgwtaIi65cFsUuH/1IfVd4LcRS4ZwJ3WbWnYmqZ
HkAB1v72Q9+msiscMUE4EF2XZummGhGDRxqDwPHx6S73ZvUev5TAKB9OMTrInfAMIkoC/3DkBQF3
rmQpZ/t725BqeYn6w6rscPqtM5ClA9AwpdQf56NkPXJdQyTEMO0uHQqaPq/mtDUwqjZnO0YDzgv8
Gq6i949MavwX0IMZf0YXqPWD+1jCJFX4e4gaKTAskCIxbgqVcNIVHXBHS6WyZFS7hWYTGs4iio3S
GymDddkfCBs9xIyq2rB1DHzWkNZMiCvuL8QNH606nY4/9AqGnJ4mDI3VTUrv25Buzn1rg0Ttm66D
VDXpvYE1ECXlJ+5kYdrru2QhKLjl5J4f9uTffhG4wj5c/5PNdjbGHmoTzHMZEK78WKDyX2JOej3Y
wROz7oLt1YPbR9nOUHCTFHWVO8YZ8996Y3c9z/b4bfJMk85i2jLJH1iLjE5QI1c/it5t3tKnkusc
a+FKFaFvEYr22895xBYXcmYCwx6ZedoMQx1JadX9mIi+cFnGnZfxNFHhj1+gUIZBPsswoBi++OeL
CyL/CdkvJYqul6S+ynPTbS6ASM/NMFRwo74jO2mc3GTbT6+lZPAacZAJ9FROO1DXGQRsiE5PQPMo
HI/nlmnyUUfKMJIfeS+MU9h3j7/XCdHyAbr/6/clJaPoN6q2e+JfolC+IWw3MaJW/grj9Bi5T1nO
0N8DnytHB/P3m+tjqFT/nuG3Zmlg9XcOqC3mfXYkmsWh6GE1j+7dwfoMyMA1c9jaOcmPS58wK/+N
ZMjMY3Jy4ZGL840dTlCboP2Bl5MLxEOTTjeyZnltZyFXD+jJ0L61xE/5rabg4iZW/iW7gcKrs1c4
nRr/T4PA8eGWLMPxkM7vKCDKG0NhNSKybRrkT+AydcOtGhdKSA+cdAYS4D/bRzOzJX5Nq38NXaTJ
k9XENgGvi9wwAnMckGl/6GyYuBJIoM6n0QNPAM2XwYP07Jq9YtaHUSVqKjo5tC4E1v1k4Y7gMkdD
R0dHqJ3Olb0dMne//jzJClTKLci2NWatLjvfbOK1hFQjZIomnBjoWBOVJ2RB3D5FP50Upa7BLDax
iEtAGzkz4qymrNyMk9IjjzWr8ryLJvLoRiCDDOcUu4xA535XoxuKz7PWUfkF0wdSLP4O0R/OT1eT
6Ht2dBBkMNCAyj1RUFtL94+sbsqIDVh43orXit334CZIz7/CbzHdMhCBK2cgGlpoF0tEsviELGuw
BXznSvwkU0KAiJuS/GG2rQGuG7XCjmsamh4rra4+JNa70Gk+H64vrD8rOzd3uqZFBTJfaimRY34F
c2CGXHS81ZkM1JIM4Gqv3jVQV9AET0HYkNgYPN43sF0hADf2grC3YdS6fM/pv6Gu1u6UlcFhFfaK
coaARHgcG79It3rIH3tmqKfiWW8VvOyaf36yMazze7FE3+zDol3uikWwctUaC79rucTC/aj27PjZ
iXbT/GVzh9F9SXWJbFh8A+UbEc9ckexjfvQD0uK96tiiBLr0zLQjHXwAVCzVF166+sqKWoxjHg8S
7jPbE6fXvKQBSTsB81B3YBY9j8AzSZ7HBnPGzXo5TLrKhtvDku6ZCUCaBQFLVkyjgfv1F9RjMXDR
Y+Y5nCeNacXK1fQSZYJtKPf0fIHYpy8kbVo+N5Yz7EGSAs5bhuA92tfkh9sdPR14K0Ex8B3vTmg5
mfK3u0HNQAqch+7wrJyBeYrx6o9KTLBkfXVjcfjnFqEAShbF8NcIhYGIWFI6bpnj1nMRU9cftPot
H8kMl8BM6FPjTZZy4+t3NxzscmXTLPdZblpCXXyW/BnJnv0ngglCtHmrtH7EaqebujCjWYO/hmBZ
wpKabOXRe4sv7HJYu23ZBcGyAx1JdKgyLRWQYJ4QBbVRQ11A+9FR7ddZFVyJEQYcEhFo5yyVnC6y
kGJ0el/b8GRifyBRHNLChOlboJyIK7v4ouhR1GwN6iu1OFHAGTH9ALOtXaXg4H/PkDQESe1VyP1s
k1iHmCUZfyoKGvjXcZQJp0FuScOszaF6tbjNxaFjGD9WcPrrWI+zh4xbOfrDEZaaFtPssdGM9vsZ
VQI8jHkaD8JQBSIKWrmuwJER3WTwQAJgPsnPVShm4iphKtFJ68mzef9di/isjUcmLmUZIgcqMNXx
pIpRazF51e7wacM0loC+BrEojKZt81QPlvcQ3cPM9SraEnpU+4NJtAjXP1a+b+esYldalVFDSPSL
zX4xUsFnub6NzsxR7nkfvCbNQPnhEErDISwP/a35QhGS0Za4hYs8JYp8VYSUqKMhmBc5W7ozeon7
uLqE/NXrMnduE47rO6eE3/E+zt5t7hjBCXQu3RQKcGTpmYysIrDFE9MtjShiMvpSPxHK1/hVopZy
p6mKxyr94z1eo1MqpXDYDBcZKAWzndaZLXa/b2oIipI7O6JdP6NZnwwgUw2KtDkr8oSBL/PAqaiq
futQdAF9IXvtRGTVaVKHvkXbwzRRs1891b+4pSpqoMYWwzeS6ATlRajb10nQZlBCwsqcOjlJaj34
rrxyo9Ws+wx2xmxuglTp5oxt3/QWoqGHmoiAaKYGVTniyMSWFRBJS1D38nCXZgLpgWyiRKYrhdHr
0uBFMNK87C3XYjVA4vnIccRlQAc9ZhI17XjdPlV1qBwxHbWPqrLe8JftHUTWL04nfCQoP75xllwy
b8460JY9qlyJIZC1BBr7dXsKIaXsXsjostbYVVlwr8kKHTzro++oz1w49Or2QO8Mzuw5nT92aqlg
T8eTIHgtxZxRSDWeeecg2xqBqwQI3lB9vdqwCGCs8ugf5YI6PtxNtlUMkqHmpWZaLSu0IzbruG2e
y8SXXQeX+Dm1aZiKFN+5m6eEm3cGss5/l9XNdGpjAdhpL+r2KNCOWjQgiC42ZBvPIqyyQguuKMp4
lAHPSmg8VSa1aXapAQQxiw7MHEnYf3tHb4m5I/Wl6MM0iaOAHqLJZPCMyHzgAzJZ6FcBiWo2xqTu
LQTH5RcC9i6h0TK2maTN69enhvhS6HahNiynY6qkuGDDLok3dS2pmTDbEwM2s3RFb+HfqhRyOeLN
HTnZ8WEeJcvr3ftunnsrFAvyZSkILILomnt7Jbaz9wDTFWG9qU07ncJtbIYby5nIRoRrbuTyNp0b
Yk8AQc+jrv5SGh8S1dI64AXd4W21pyRDztM2AW8JqSyi05Z5DXHLfsAS1NwQl4KN179DS4M75eO6
wLR16pRkku2/d+fXY8Te2pK5a4v+wxErPlkyXmEc9yuKKZSBUxnU3amIrIQFFRQLm6BYfQhRi5jB
RmddodInT2UByZvGA4T5xwzIan/o8/+nGb7AAQvez2p7mEKAm1TI05TABOXmc1KAVp1HyAjmiA2H
31Uvd4samGywrFKG71NnyJxybWKBh593KZkUxJtOb6wO1sHAp3n6eZ++/kCOc/omftkUTOM3N4Rr
UgJTCuTRAu2w8EXIqLalk45lbI8JJ6/MVuKtWB4Y9g28VqKy58g2Tdhkst6LEM195SCv2Pwrdb91
89y8ERuXn6xQbaALM9rrNzKGeSWHpIKMtITrIdLqj6vw++9jIkAuto7UwLz88jscCk1bY+o7X+kM
lvVfItnIzg4G+SrQ7d6By4ygDh4sATnIdNzpP9gnnGE2yoNMDQf1F5HVQAsaVz98zE68K8VDMFgk
IgKeN3bh6u1JRgYOvjZKUzzg+a5rPWVSR+nVWNpLhwxF/J4dXDSo0J5t//OsLzhabxEjVWzYVpCb
h4FuGHsKjXGzPRQrA62GKg5Xjj8WDJHISMV8OPVtj8RbJ/mB8TihT9jJPUZL0HIjCpN9ILGKZYkd
nSTFYSpX93pddsfzc/eMF0IIMqCnZUkzjMUKj5MEYa/x0Uk8OcMtdG6HwemGs+1v9xQUiP45UNRx
vAgnlOa/RO24B6Lyq5sDSGJvT9PgjPQqdvSnY+yoZrLPUKIjWWGHY0q8YhJp8FWFr5wGu/paptSp
dPaQNKVh6r23MoXW0aRK/fkfYlETmJmKneamUTwbmro5uYuunULx85qeqtDxxErf4vjX0N5jY7Vc
7b73lEWIViaQP6I7t+dOddJ4qR0f6emjlL031Gaj7rF9JYLH1zU/WpVqdGaNAWZ1QyrH1X7jgWkj
ZwUZKXas1/3UZoB3uhBPEyiQlJNK3Ws+kq1CfAGTerCCKC6Z61tGWBeQmdUGfnDcyesSlkmhsNoi
8CFCWPHI2y5TA0SiN3F11uCWVAQM5/rbwwd7ATDCNsod3prtrmLqh9Ce42fOMjfbu3VVQjw1YkAr
EBzDxv7pflVYJZQACsRx+yTghWTc0iZ1YLvcQ7FKKJWPQmAr+2dIihcIQWkPhsXS04smgh0FI5ft
iHNsZ/LncVbmedMjVd1qSxLKmUgq42Q8nllAojx4gASJ+EQ8fcxws8aqJrKELyCkKG3v0q10M3sM
/ZTSA8IDDO8tSOVTJycWGEnYOBgESaI+kGjv7iKlDSHRk2ZqYEaoyGvWc7L9fi7LKNcksJPXCbNe
Aq0sBLYxwBfugHqmHFiFcKNByEp1S67Hrtq2PaHqdq5SGQY6AQbdTryYwbC3MiBA9ggpnFGdak43
1AZpWSp5SP0h1VGI+NJ7qH2RHqNOuBA6g56WVGJhfLjh1ts5GmVsaPDObcoCZ5f4vl2/L8O3/j5e
EhmCQT12WK0lP/A6Am3G2E6xy59CGefPtcG00oxPgTZKg7hxE7lMkatdGld93+cvHG8zO4zVIEQt
BG4EQUDff0/aSEn8qRMozZjq27Ooo3p2BeS6sNGWOYan57tvaRiRvmUlMDeBSN1Dkl5w0G65Wcce
3/FYDl6NLPMWpjfO68tH02sRoSYuOouzIX+CIskWgz3DKLJ14ZYHhgABWlj41ZC/QIU26ZCIvokB
nrFwrAyAoYaQti7urodLKr1EizD0f5afkO7cQ0uju3ElnivzrmlF1Q76OyyMTvn9biu0mYIbu7FJ
mdvxCFKwR2VGXj/FonW1dzRyXa9p7uwpNRUsd0W6vMFlB4jUfM+IoXpE52sYEYbOkTt0V5K+wBSH
T4JJIVAz0Pbf3pu+CZGWQyHVJRZWjEMKvv3i2yfnl6UGk1VME1/qFxhwKP5fEJaetDilp28NAPNf
nyl01jd7tNUTSsT2vv+v9i+Yl12q284N3tfcHL4qiR8MwDV4B16myJXtje3ClG5Abt0hb6BtlhqV
+D+hUAmydPfjThBzRAhozmcM4H4y7sSOAR3eEeuJWlLFo54WZo0OZRb5MXFlW21VF60Fzg4R+a0+
DVdflcjfQuOW26IT7/RTIeMf3CBMVfI55B4ZPg4kecLXVkd+xPB0DnGYpv5VTQoOq0d246NImmBV
zDTtkf9BZAwqav5RjS+/FJ3oSxsv9Ga9kTjOMVv19M9eH1cz0rx0cO7z6m8RpOazrIuWZbjubD9e
ERVT8SxRk59KGeCh+cOkYsa1if6IWK4OuIMCPo+/DIFrAxLH9c/OE39Bpp6ENYQpa8/TJ9ztvKtF
IDRyEM6fuAFi5K70cbKDtRKDgZNvVnonx64BvOR6C1jmyxTrDD44psbnIoEyNn02GrsLQJFgcyzP
mdRocvm4+NDq8SC1exp9ck0iXh2ksnXU8s12cGEq8DmQEP2WddaklCwan0rGCukC22UKN/r7y/wD
khNpo/1VYPG3jVQixZUZb+Uiff5UGO3mOkebz6vvNWLy+acfpAr7jMc7Iif4U9v6HndbNhNnP34y
OPk5ItnB26VgQBgpo2/N3klNORRANUjl/TzT/rktwIOKtfP0zLIkLesKm46ydWITnS6gLrn4DaDS
Mivoral9NK51DknnEney5D//HJBgfggXIfY5exlRmNBr74IEtEANXbmz45EcHavku83rcGDgeL0e
iWsKmxLaeKVSKM8tCZ1eqHvna4axCeDHKGlmj4UNMpUWmptfiCeaEjqn42INWdLvlbacDDZOyc2F
QtLf3vEX9wytcUyyf/AsejXwXS2bZq3ijTWBXOTRQYnNp5N6zDBTeB/Q/TZrcI9F+w6cMYq7Jhs0
QA5pX4t1CtEmWXP9fbIyTJD9NAsGgkRFLtrQ4LGNzEqEhRr+6Oko5EvPHLdnaVWaKZRmsKGDwlQf
3wnrZBajt9Pwae+U+RbC73OqdhUprflpTETSk5WzPye0GrWbrTn4vd6JrZmshUzE1zDDeH0evXNL
u4JBoUUj+DCWHkvzBEJfLzQ93K/oaSwcEtgmlGkZx5LGP51kAIvQk/mRgg0roYjxpqvIRJpkusXB
+FqGwaoaZUQGBBP3NiDF47nGxWsf2ZyDln/5kkw0sfS+UyMS57zGYxLBmz8GcS7qzvUmHbmsyKtG
z7wiPfEVulAFDFfFKaoNEpBE3vx//aK+dizA33pJ/jX/ljHOt7iKIrelNiAm6B4oJeWux0z/S9hA
SbCkXJDAJ3/zMJGASl6XrPT8eTznHbdoUitv5Twa36kXYuxicZpqIqC3jse5e8iYgQh+iPWf3qX2
bb3/2dkGFThBmmNOiXTljo01U98wRMKz3qrggHXO8+FzDJSdYmPiu69wqs6atRdyHeWrifWwRUpq
uJY5G2Da0iWVbjI55H59dpvmXyx9QwybmvG7LXF/oqEUJKXcg3krctpYwOA2KugznobMdY8odi3T
ySrz/HFTfTEOhI60TvBj8chGn1ehXtYSrJTgBopzPhvjF8QNyUy4YxkTxpIFwWJoCOUNMdDI10OC
yieTsS3doQpxIly9xFTKa6hc6KTL2XkjPAb1FeOfrRNQlPUxbbww7d39RIov84SoxTbc9db63nGJ
CHPdKcX5Ui6xA7ICk9u2vTCrdUInx16+xuSJCG5VDHX8vlxOR/gVwWPbJDl4O4NpPxi7aYe0SDp1
8EHN/dceBWx0V1rGNcpWjsdnYHgNKpIWWEKD/00MwnGVV0QM/Uz6C8R/FXDP3KptkVa49X/3axki
iAZD/f3wEUNk72OhF5zwpBk8q60xTIJJDcfZyi7klCH96RXqDOmIdsJci+P+OER8fke00vfSCY0q
5Gx4bSuCOxHONSzWgNFL88ElovcWbRvmqpaGnvgb/pVsMMwPUFi0FF6RlFu9m9ZB8uk8ZhEx7g1t
CYju7T+gRna94CpfjAhAreuzQUBOr2KlVRlaK0o255bWbwlJ9cpKQlr18gFh0+RbK7PBMY3gccuF
ceb5llYLAtuB6z/4sOpjb4xVgaK74kk9M2lX8IQsoqMF3cR1CiYYCsr6i8d0vSdZhQEs2LCeU59l
tQNRos8btaE6HPhATSzAOTWT59nhG6xwXr7W9IBM+4GpVJOc3J9ep/Ih7OmPBTE3c7d34btbn7nq
y/xB0/aI7pUYakjyoMd1f+KuFb5keYH34Cq/517VXLCKo4rjpsiDyjUKqW/bQci4ME6qQXyv9KdY
w0Y1bShJtfgrzqnattmW86UZ87sTaKeHleii/Nu6fVAjUBsAPBOFguHIOXO8ByxnruNHe4ZwL7/9
lrhLQLF6pqcGAdJzrtpLyFfjV4mS4CzLbulaHLJju9idJOQXd2XEhEs9wYMrKiZsDk9drY+Le3/z
zkKNWrrUGnz2DuG17Oc1UoNy91YgXnBJ8Q6Gu7Jggf/jVrpHrDf453tueCJauL3wx86lVcla3XGC
ttnzExSCsJ0xFmvqUnAWD2R46cIDbdRL2mh2Tmlrh1hdbUF328wrxzl/87vUR3K2y/GJAR8ro21I
8aQnZNdhH5Wyd+a2ygiVoGyyjHtBg5hntvKqCdnWLKts9CKAGToqpye0UjNZcKxlsJqL2SOUNRrr
Rhw0Rc4AHc6cGm+mEkOETYtoJ5sfHY4Zt6Hl2kpRThdyfONR4hRe/tkO7sD4HM1C32lVkCIyAt6t
GmyJjJT8HHpQyZxdDlDHY0Y+FbYX0kDtrywBbSUoJuqb4ePGi2i7ks6V95Ny5VbipEY1iPjUVxBv
oEjV/aujdUf1j2HrgXX5C+xEQsu3NuLo8BEelM30Z+6dbZ3ErPiNEYd5HfVhLPj9mvGlgBbUBsab
u3PFfbeZpfn5QAWPsUbjFrgxuEuj1CYb5TcUPE+fxCvFWU6XM1kgfj5tAvzPrgSWbzromvrCN+Ub
AcHVumSzHbOFVFOU0WqzJi/BXCpuY3uv6+oncRTv+PDGjyPRdNnhoBIzA7vLOy1ww0L1SV8lkEHn
ji0UNpr5Ebu6DJj5SDw145aECCbMSJMESGWZsBNJrvITotP7ieF+wHS6K9xud7rlK4kZv57cbHNl
Dbz49J3pj3I4Lr47WeV/L1g8ZV2IAoGCPD8PtOWK43yhI4qcL6f4L5ZZcKbnPhzL7attKKjivTIz
M4jhumoHlS3dka7PZA+6xaJOMGW8PwiPFirw3hIH3mmsfE83LnJtDKvW/fJXQvNdsCUilgT3v2yx
NJmf7EmI/03aCyJzH0jrHQWgKhCUaP9nzTJ7m2F49vyJpSi3Hz2dodbmIZWsSpBJhVKqyoTfTeRQ
eQAD6/9wAc9PhXSaIHsbspoR/ib8HyNGb8/mfh3w7wEc7jukq79N4pzUYnSSsLZSKEY6giscWZYQ
l+m+DTglR+OEWNaaIqYv78lUBuTyLjNOX2JhmB5VYp32RT4qiN9oTVACYLhUzss1/gbP+hjKl8GL
rsGJxGmtJ6aMezGhRnccS2ElmlbTcBSYIkDu2vwusHZUkr2kNG00AD13KRakUDkwg9iOhUSwvtKF
2AzwCNYxciNiv002Xher6LXLLWKfJzmvIinaR6DQKO+bHFIT0ps9CGK/k9SMIFBBEkRiywlcKDi9
X57sLBzFLxO750uYR37s7q9GbEL3zlNBtbRAJCPexVQrsREtW4+CyAy5ofDlPiUUkS4nuKozNkFC
UyjoqAU3HvE1Dzn+h3pd8sd8asidHjKcwEpQYnvESizA9OOlpvUmWXc8z4XtVTvGEFAaoWWHMdcM
rgG/wvznxVfERc9lRLB1RtOUNnN0k/1zVujuj0mvmc63mNSIy3AVtUun1GffOPeSBkd3t1TRwBGP
xxjB7yAAZlFuhX27EEYqCEUywDnHU698RZ7RgGBDFWrEXcUdRG/6rlIPL/BJgZhbYMG7fuLXGFsQ
qN7jgk2CfFgN0ZrDANOGRpK90gaVBQA5SDyDQjnWNrtKuWsu0h1AOB5HKlJKHPfM1NTp8J9iuihS
csMv42ojo/k0t1CyZ9m6wCk0R3r24ydBZv5WIGMbIGsSqnwpDWZc1eDDQ0XtWmshlrrteEP80dFD
v8aD163s5Vs5oC6uoZdfWOWyBAHzOFRtxWNfcuEIqWZTDv11V34WEWlKyAVTrtk+jkPuX/iFAI+2
OTh69rk8A3EdMc3LQbc4o2NneR7fIrEXoeexm9OMACsRYx/CKnNID93Yl+Mowt5b5ABrcmgG+QRI
erYsFEZKLmO4tmM5kRQdxzFB8pBzKgdKQYwqhBp8P6GC5Pp2zDwWzuHEF3/79+miItazjKsH+Jwc
Z19t/naDUudQXb5UrsJqqmIkg8U5G+ube/1aLDjwZM9+LFpNNUYkn0y0zGt8r729r9ZX+GRBW1j5
KAhTowNryNTzqVEc1WVtbsiZMbrF/hS/Z1+yIfGS9Sj5SUd2JCZ5C+on1+j8ShLmRzK8lW+JWTNW
/RcQmowuK/IvSnUXq1HDRnp3QVAMGk/+Prz8DWKbNSuvvjJsE5LdwSNqUL/mpR5QvQsjfl7A5H1d
GUfh5ezmqjTdVAyX+no0KYgYzPGJZ82Uk0MBWNniQKOuzXCUibaQdkz1G5JS3YCB/n2kSCquQtke
V8+b3v7q2gruCLURrlJx3YnTnaDfcmIWSXDJGyVONk2nyEgPCuLaX58tFST+AB2PCuLdNJtyO/a+
b4sP7Bm0pOUB2ZLojNwsyBSdqsnXsrhsQ1SUtfWyhlnUJnQ7UnPc5ZJnxinFL7er8pKrNp2q4d8Z
aFf9h1uzDzDHgEoRkDZ+rtvCYO7xz6hqEY7AeM8DIA5LZcMuHt4E56BZ/f27RnOgEY9y0mNNGYAr
xoCjjHo/MU9LM20ceppiJ1nWaREj+KKgwPe5vHvf1haWPU8WCXwX6v/7sm853R4GtZ6PPlI6R+FW
gESIcCXE2KcK+SbTdIY83p3jq6W1nkMKKrhfOYmur3cwZzNY+BczVwF2BebsW1Fnjybu2Sj6Pula
Rl2q7J5JpD/f37DSE5d/krVDy2FFxCHVCHsgksxd26JjMgjI1M/TLJmzFEWORx+/Zxolp8bUs7gE
ovzWD7gUQ8NsRiOkWdhpoLlbkcFzb3TXsegtf3lMwyH0aWLVSRZQKTHFEaqhM4qvonK5CDE4Al8x
6Sf6L20510PoZp+JIsvbf5BkcZuRo5xlHn7IVDtgMr815nDnT9YP+fIgPK15osL/u+KS9Ij6INBr
YC6LHH+tC2QEpa0t5+puP2OAfJSez176JZYncz2E1uuiaXkwXH/3ajwgndr6aFxlzLf9FnD0f1UZ
dTGpUc+h+6/UzRVdxGq3yxn8WJI4oYeFYGyQ75Ku5KbgrZ0c2Hm/gIaH4Ji5jYRV0GDC+DdGIGUI
77Up1SwGA1vud8GCiNxbtnlZQ992rrxUTpyPgNhuWtSq2UROUICnw7qVNvc4pT/vfD2385N7jsFx
diUxGSiJGCiAMbO0X8fO+1hLUhrSuZUeQKqAUkVwT9Oc1OkBoJUCoikT7Mu+xnWz5rW/fpjytYBK
L9v7e8IYi39Bzy6y/PXaTYXCq6krvr8YttCTRU4dtdexAhargF8xOXiZBEiMsLS736p5dCmeHsUh
u3YVBEQZE2RDsVZ/XU3kNzZoIsnTJ/2tg9B7qQCsH74oQGbJTZTixqJ8/e4LVWhMAdtHsVuy8bly
utHveDR/71FuybL12SbHgQRuyoPPs0LMmwMUlKMJ6dwCjNfJtE2Hn1p598Pp9iKAXpLvnrfHPSS/
u1ugDdbOjUGHr4nQJgMba9xqTnQ3cypSIb01G0GAVlIn+SlIsZbvJn8XGGkOBvRKJXhy+nk60LMc
0mVJ8QVo82YiqFQHb7rWJmXI12xqFgTYkpnwnrJSlmthUR/+GltbaU+CKR4eSqUxTR5E2O3+iwF9
TIRAMqOo41HLwhd99WUTGE9laatkFx57WBGOQGE34DVKZfg9/qLmxQCtWuwq1qJFYtk5ZtrivI1V
S9uaj8PqNvXc8ksKQ3ypcPgaSYqR7JnA/3IZa6E4TFjrxYoczbTTpmOXW2SEjR7Cn2OhKwR6YR9o
s3EsQY/Rvz9bNtznNGm1+soUOYSGdDLjzsU2kZ988fA5CA9ubmS4cGOpOax0wTJGKVJb9OgFKgPJ
4LgPki6rtL+IJjmLVX+BDcUflbNGvw71ur+18tE0r9mGe3NGhOlNd66QwoCrT+5HFCrtM5toPKGM
u0t7DqaLF3t5Kd527VAFq222rza1lmp+pe2528TGevBgww6qZAHCiUaxwdGYE1baniQN4Y1J7T8v
OhrZ5Hf9BuT5OvCp4LN8U+YG6dx7F/i7i9ocVRiZCcZDxnBFdR2qNBB75iH+rPuYZs5du43+OTaN
MScBIfNfR0BW9McdQH93PXNY3IUBKUMXcbZoY8bj3plmMA/MKV2Z+N5DKaDNRt3WuFir1PfzFqYm
SSZoLVnnqPazEwxZbX0uiK9d4GI9MbuEasVORzg/GYgfWBEsp3zOJDcwWDnqhDpklgOF2joHHesI
4fYFxuvcycAv6WDdjVKFoM48DyE6gmlM0afQEF1ahEk9D8plX6I2T46S11uz3BJuRGUf6rSI8LcF
WJq9TaMvH6nPPDnmnCnSPK2voMWYMSdOnHTe9S4qrzZip+rGZG/d55veDgykHGu+XnRN46wwKk9z
8bsG8UkHuiGMxwbptkKYLNyhfetFQgPQi/wTmJUevfzvrNeFAARPhdVk2kgEZ3kAEPcIaNtwbPP4
E6kXusx+4tFw/0CeTxz6RCrjnwvJvfYG0h0zly+k+vrbEMmKjqYv6HsaIX/LsPZ8cnBft9PeMoPA
jVH9A46XomGBQDBVCjSPsiFq984Su/+xBmh8AWCnM+E4bDFoRrLQsUKvQLYl3qA3fOcwaLAeU+zx
7Z5iUOKCsWl0EetBzHQ8BPgTysCKhnP6CqnyUtiofsXOu1H4mvmYjjqAJePw3gSamgRumYqjveVF
TYMrKfJH5j36+MkM5ewXZV4rWUzYv3hKI6wyyva6p5/H62N7U93CyKia0iBMVw3Ip8owFXXOBvnX
COOZYHdJJCTYxhAhP3WLvIyg0lCta6WNS5baptNrRRJOAkyRkl97IovP+htLI7CxHkGIa8jQInnR
VrbJVtuFvhNEQS3jC+/OA2Xw2cIjWlC5L52xx1KjsKk4M0IsFO+wyMuDJ7PxDy90IAJjnUhYnH1E
jK7/gncpXDDVxVyL5ScbD3PGSDYu3eAaM7E4RPiNkrJT+a9ygKnnBTJL3qi0/N9gF4f9W7Ud4OGI
jfIySjyUqcmUyqrkt0BTMZDoMIHhrvC5fif98H7oIQ0CpAufgYh+l3inq23Xi96CWzZ2J9Am1oxM
g7JDQbxBWNDtHwnx2aesRtgIsE98Jd/hf2uxdRDux4UHXLDud4x7PqQe3h91GmYarCZ8tCo8V+/Q
e49kLRG08lLnsgTmzexDQZX60YeXyKaM9XNA8ppeXq2NAjyUvb5Q8RR/2QY4z4VoYfB+n7bmH7YR
u92mPtT2L7XM0adCYzhCbBaKNaKnJbzq6nb9G92nGBPY9Nie/dwiVXmS5ZSGufyFsiwfh5swV3CR
ALfaHKMQ+8bjRRb2prGiEuYn9kS2J8srDYxufKFnbyg5BuLb7g1jJf0B6vQTJDAuv14FV3uppYCA
WuYNOQfuNQNnbLHMjPmuWaI8QLh50+hn7KM190UpkNxzlwNUASe1opFnc0pvN9qO7NTMjGT2acTi
iX9IZHp6De7cp83bdB4wKurYkSZNB6weVDTh1r4lnM13FfVIvDsPVkHrjViQC8DyqPKGuvJTDgBm
bgIyAOBJTH/dpCG2xuBhcGrmYmMicJkxf9uPM2u5PBJU2RKgZv4C1S+a7JMzsMccjsNi+QKdyWkg
7vz/oSRXe0Pyglpv7qM9/aWDc/quQIUE9Lv2xLMnYJjaICyD48JFgzRreu7caK5SuEnTADfN4PUb
NKwxTmtWw2vrszV2SXButi6eLIPmRCGWY6vBF0+S7uJFN9CMysFEtV8cDdQoM2mcsQM9NuvYtX3l
j2xGJpZObWgV62bqwV+kDw1cakemSavonER0qMqgQwj+QAYk0At757MRouGXAICaOLBVrHbTnHWV
SoD96skRQLCHv6wMFF+GoEIWR0Jnl1G4+R8bThO4WxiZyk5/BVLBHGt2WH9gnhvTwZw54+tRQAhf
iSen/eijju6AXEv/NTOM+t24T53Ympn5hxxzXD1ETBTwlYdxGvjuzNCDjvnBJx3ghIADvgnU3zGd
Ojqk47aYH8B+lp5rYZ8Vz73PysvdFHmLjd71b1DSN+baa2IVz3j1hJjnA7ejkX/c9DG/iKqvoZb5
gmCBTCrPiQw3+O7qKXkqxkLzckA2rt3kptg7bIF5/fajLsBhXzaEKrdlKa3VL54THq5LQIhGv937
etU0RLsg2d+J5FI2uLRAuJX3MkHPO220BDUQhdU69P5vbiiJK17MxK3ZXxUO3dZXkyiOvUGfhrQp
i0oHsca3CUQdXio5x97H7r9EHuOEtpXm6BaD6XD8A+0gdNIj4iGq5pq9kACgKHc7+5copvzqTuN0
NYjkVK6mJagTXh96m/T2onU5dnzPCX+rk7QOwUSmuIZMQv6hqTyXM8PJ27Bn/H496zwJZk6nkLHP
fba1EDgZMTeZauix2hQ9al8ACu4HatfyQWQK9G0hJyJ27R7bWhzh+8YqX6bO4lrvJ1g7sx3oYnjx
5vF5U5EZST7sjMqIJAQ9foMXV4kWNszOBxY6v42etYFDxOKL+1TWppNPZJYcfU9ezJ8YpcWE4M0X
/Lv9QXSASq9J03jetma+I9+7GuvuMuqJTfndPfn/DbU1P8oH7cb0k6EY1smkQ6Yo8mRwZlVGf577
k0hd+HXpjk8lWNL5BNPIenT1sZiMraf2ELQzlPHhwjXZqLaGEd15n9Z4hkCaiX8+O32U28qFBeXf
e4194CfKMYNPL6/z53Op3CvL54JjYnu9EVfWNHcQ2+5qXd35HDVDS6+affEfpc7XQqL5nM88TDFj
t/dEd0Co8nmQrZCK6zgCTSnjNOJMSeRY6zW/sl0fAvIatQvqoS8qzpuTZpjGuRGxMr5Yx7Q4u32q
OniPNBw8QXcM2USBTLhgDTeM4HEsdU4OvTPFi0irlcZEzxLfGgEzVh/1x0TfaIrdzFQN4FxUHCH/
9fxeuPETKHyTrRBf70l9MsJhNpmOVFDGOe0dH3KtRaJVc7DFhsmj48vdi5JDyxZubw+/dt8ls1ZT
DYup2R5IjQ5hJGeeu0Y=
`protect end_protected
