`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
f3hwMr0K9zJzgDIT3bG2mKyPLfLy8QEowmMzL7vI35cGb+DCy+2XfPwmoUpsgpCeCuTU0NJwLHoT
Imr8cjEnmK0+PB3Zy4FpM6INTqIg8ZTBmMsskKPHgXASo4PgeXxB4xElxGU0FFq4Jyf/WBJZ4mSS
faUrZ1aehGR2ERS1TG2zBS3iPw6H2L18hq2n/Dw/oPURoQZ1qdcmlmrmiHa5qAmXoIHyxh309tWT
jVN949RtHg31JCWS6RtDi25RKeOuMi7g3DNFci05imXSzUn32o/St7v6S5execniigG5ROpLOnL9
v/8C+A3c5LeDP6zPdHQQorWx99CUM4QJXaxT5Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="CLvkpxAqTaPY0nYTlMj4DIY3zCMwRAC4VbMU/dYBUG8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 130800)
`protect data_block
aTHAR3T2qp3xeqr/zO6ZUs6dKxyoVW6GDQQmwweJG8WHfbYRpsPXgylAfiT/93yv9d2UauqjZvRC
/HICRYEDkrkoduL79N5fdBOUMRB9Y5VL4xXvQeL7792AbvQmdjQizr/D/uthNatXzcRHEUp09+Lr
ViscrXal6pEEM2S+w4cyDSHTgE/0GoyFA0VKEPiRi4PSFWN4ID+eM8TZ2sdMtq/B6rz/7KsVxsAC
tKNt86XokoCtlGNQj3LJi51w4Rm+mxwTA4H+FCU66+8i+v+AWxCOGDEEkQ/8dMpCzQ9OdqjXTKm8
I3qFLtEs3RsXr4vTqZbf90KexGTSSTwzOverAxJlEuT4VovgBK3Zsb3oHvdcHmBrJYwLHDoY6NQb
odyf/q80R0CglsNbWl+KkkKRCheiRd2q2vyWDiHXD1TnZpc1CusCyAx55Wr7pDqNkj+2FnxBxPO+
CcBAu+rtDjWCd+CIFHQxY+IrvKeMSytkmXyRZE/i7i4B2dKJaJjd59ZMCKyhHioSpDRDthJ+K9bw
hRVrp11Qbu1t13gVvx0tH20d3RAQ1OSHHm36BF5LosBBeegO6rTqV8HVG5fdEzVRgx6rFLAcxGQV
j7lhIvD5PRrbRudm2/RaBEDIWxKaLBUVI8LxCppcGuZVBd+++FlxYVWcZsVxO4z5FDK9ChlfXIBl
F7ul47TPdQxoBKNMNS8dctzSeIUlY7NwiR/2kPIvB40P06lOBn/2AXzYgJBV5ttE6ze1N+2BGlfN
c2P3l3p+X5sUcAg+8YMX0es4IoqrGOI3mRV603xkleTqCaoIt6q/ARpzm4OR0Jc5zXO0zYWQDKOH
MlwVldtbrt3MiXYpKm+MU0qYeKregJnc6++RBzTzjD8h+wI1ujtjMkisOJBui5mwUmFBo3oUOSd1
6rzD/LB/ewCfMhOQZO5BuzaV9L0C9K8uqhQHGElDBcAhqhAJTbp7Ov1v6ndKt2gDyOzHE4uz1gsD
VqGS09u/jeuXtVtip2DakGktZj9Arlq6eo2bB9yR/tGniWMYk8wKwyxD9eXa0+expl/Q7dk7aMWQ
C8voCD74cNICgbhTQu+qARrqza9RnNhC1R9/mBMS8Da4veJNX2H4vQ+2sjbVXc64JEH6fOD5DwGJ
wQyZkShu8gCNNy6k02RcylJg05GBdO2bI3U4qG52wdfSb3epyzdVFkathcP5TTmP55/Ux9ctKcnn
5SKGusrKSRZ8/iDvRKARHhP7FF8Uo4xsOt3hTjU8OHl2tHQl0CbcL+vgGp+9U1O6Ib64Ph2Fs1i+
236dchN9Y/6JmkbhvfIIJoV7cMJQyjcA1RujvIqBmVN0kCvc8p1l7Auyfmjog+HnHyN2+jI3Hl1e
CrlgKhT2+z98OSIKJZSROiy9kDCX/VakDttAcFNSW2nVMhlbsjIa9BCxzrw9jqovAxbKTqabs3IC
YR3JPQLF1NBCkcCDpy9Tv73jTJy2Q0wDhQVleQRyeM7eKpRfWPWSiEW4WosvzIE68ZoXt34J63v0
v4SC4zT/n9wCnvHx38M5JdBaztDQT4P8alWucywvtKVTNPF5wzCHLC+5auwbFeAwnlrrvmKNbzTq
iIF0d2zEIEoBV4Lapr+AXLVXeSIb25N8sdgvwgYym0hAwRp5Y4O3MsLJ6Dvn7PCaQv55fqyYUuST
wkh0URK5x35u5hN4dC6J9I1SOALeuu8mhlGqmXvret7rzOMcviHk+9v7n7ORZQYRK4QgadF4JQHU
nw7qFKN9lrvBTaIQ88xbKrJpNtiiuHgI5XihtAQT3NaWGCtHNROzbcHNsSjCA3laB4e6xMqiV6yn
LzFX2kayhPVUeXLrm/khW7YehGyV9r6u9asl7InywE5OiBNZlpzM1T8k4+9KAe8bbjVgCwkmak4O
ske5LvHZg64OKFa6tghOSPItd1064znTe3LiOvhpbMxNkpIEBTsVcxM7eqQq8OQXGqEHvRNgxZpQ
2EPuvG8nxV/OJVznu7vHFsc2szjzT9XYXLyaFb3it4Zwlk6Az32L7AJqPwOQWXxwVnLlDlFxQ/S+
ByczPgBSGO6L4QdY0uxohDTipJX5jn9gi6ZqZkiIkkjBSeVFoSg2bdbwVX3FnHEHM9Q/geM+cgXk
5xAe9VIpKhqNwW/RelmK2zQw1TS+UvM05WHqSbSx0nc4XRPkZZ3z4pwuCUL7rrYZJ9GKQYQ12ciK
QAVJiN/sR9zkwyUxjx+DOMSkRtidgvHHJQXCyRW9PTMwjpILR76nArQByoq8gV7NBslLU18FDPbU
PEgNoDCwlyORharmQ5r/N1ztHAIy6jagiZE3L63/JqAZUHiMvr6ZsC2bnmaYWSQN816so+9yxJAr
WSg8Q+mxAjTPM84F1dLdJGSnz3JPmgP+ly71lIeXBtRQdZs93FV8JSxfrs/L/y2KxrwtPDnfr7lR
CUf/09t9p73kC9+QuXfQPIXOhRzm8sibjf+IFyvE6F1gJtTZ1v444ZsQQbL5BMaTsgqjTxH1bVCt
RXqTXXZiSW+94Fz4kJOCYp62bm2SIi4KcROqkC4wxm/Ur6hzkq5Exz2auRM5Ze1gFcUilvsYad4I
tikrJ4ceL7x7UFhT7/JhoA5VfBdjdh8iEI/2EzTvnxkELhj7nJKlga5YmAkqha8VjHJhu+SrDTwT
+FJmOx9s/9dGPPev5hUjhWxR7jJgKg3dEyzn+wZLKye/niNueC3+igXYPvHMRG+7BJ2Je5WMvhSy
XisCRNM6+8m1oEGGzAydALe9sQicnqI0jbOaf7MDceMqcPuT8S38zxWMfD340+Z4jeOYwNqiGwVX
HD/Z/Q19b1olpy2e42EMxvRqzYGxmMRL6CvavdW5NU1xBNb/dnPCWzd+9hyzSTxmhcPQdTUUEsvH
YHPatOV0mJXpcFjbUii3g9lNQb0OG1Kd6ap1IP4NESdDCFRpdO60eRhO2CEEWEMYpGRRbHCc6C7T
KRIFa7odlfo45wZNh++BfkNFkHcEO6a44D7p4m7vYncRwbx/fHXSXcTeJM3/yE3/ZK28W4pVakgp
c4pF+ZwZ2FZHsCwBpNNzaoWPzUbkm8jxoPFOZcU7LDJfLiuE1+77nxNS5J+KsDlgxqqJB7G6pzDe
yIl/2vFvRx319KKFPgfYQi5ClqXsmUnQheFtepqapgxvEO8iqw35fgeEtbl56ld8U4gNJ5hca2gv
e3JCedDEoiYLv7sGs7C35XX1oyA/t2I/x9RWztK64W/bOQtHsj8ygk/s8ZuWNOPqrMUjvMl993P4
fO3jgrSNlT16tiZWb892bg052r7Ye2k4YjxtkDAhPRXftiBEdUIQKjasyozn/e1qneDadiOaSgGA
SGp8/FiV+LtglWVPbfSHCzrO8YLqeeM3F+2ld7+XPnFwnOKqmrTNoB1j/zUzXb9te9a97QKB9ptm
S8R0vQQ/FcS6l7XRMOjHI3m+5XntzwX3aRPIYZPQBU7Mo9zkMsPW4e+Aj8Jk6aUdsCcwrDysQ/sk
zaHsbd3zBmm5RIRd5arN5HUVCbpzG3TZ8RN/EPs5yPoQp7Gyd2Doc7fwNDvYDQOHD2nfDVhLu3DN
/PjtM2zICc5dur7hhYd9N9MQhw9rIohKR+z0+7nmfiyfvyahrsq7xcAzwXj8itPqzd75mQTyT8YK
2xP7C1r9mM/wOjP8ltXXjHyS8Vb+zBItluiX6CUDf1YkCF2GR9m7sMN2yLi4IGSRYFjg3HdTKOJ6
pTtcWC+J+K6PmmDJb5hVYpJ/Yu0yx2FVxFDpoKa1eh+aUpnTHMxqHc5w5MqRQclkXh0KemtP3jnx
rXdkydJLuODTcl7S0ckKUViTkDpDj7r51L6mYexwP/B0mFYlJ7PfsVa3AmN8DR/BHps9e3C2pnFX
n4W8D/7hnB/Ec2OdgApNWjKr8v+XXrRi/rWsafJ1lhOjRcH47UZTW6ShHhf/SnQfpz2waJWcIKpX
omba/rkE1TEXPyNPBlgb0XJk8z/GtojtSZkf9luBNMux1g0r1OiALel0JdXlc0a6TR8Myc/eyiZK
HBw9jPn3FoRsiYcvUSc33ls5nBu6e/QiP4DRQ72G7GSz04UZ2rugV8Q/mVAHTXebN8AwIn9EJOSz
uk68EQdn76fEakJOJPg0E+wF1On+7vHOQmVJovIt3sNU0ma2jKDJMXQhUn0+ZhIpIj/5MQvGz5AX
ujtSjCpX/CvtYQuuRRWuRWtVj8fP+nOyuCqGFA9j4FYQpVRQvfnBLxRCdUH+ACfmM2GOLOQKt+7P
UvgA1PHNAgl3wrz1zf9P9zPNuyRKlXOjS6yF4fKOI68zIbSoV5Ixc10bAizGQO+sK8T0a68vfU2r
fuoNLRvDWuWoEhJjrZkE5+C9yVXEZGxj+M8hYSEwCRa/6QWXGF7d3dJXG0p7rrdCYtQsFy10cscz
SdqrkwUvGjZsTKxFCEVblw91cd3HNwVcqO8/4Z9koX8OFh/0DVVMhIoOzj6GFWnYmXa6iqeLW0bB
8QqkJpaQ/dEEJHAxygga9Qx+HewZj5a9+V/LkSv+9MAWCD2xmrw6ukFnF29WYRDdnUwqea0xvJy+
Ee1MvCunXi21xEjy4z8seOHDxMqi6XmhNpl+lTWPAicKH5FY1iI1WVvZhMS+eV4rr5gCodBRYuNg
F8aOiNZcazs+cOX2fjbta+gQmXzucFXUw/0feqH2g7/0hlg+Auo6rQxA9IWlVgGNEosz+Dz5GkOL
i8pUlDYFSlHGv50RcfYOTOEYIpjNz5zLp+LdNHWvc85ojReWp+jQBO5chwD9lEMkNImqaDHmh2Mp
wNka90wl+kOoqcDq9YmxWgvRVk8JRs10goxiw+pBw7TrVKs0UVuRL8iLrTxxpNxCh/JCZXe5dA8i
ynVPR1jGEl2RuL82Blc4m0XITPV6/CireFlmVHhEhpgs6dinMv62KEmnVCOQKRP8ayCzkDZJpjpi
p0No3uGMUW//TP5Q8ZZFSkmn+J7/ltZaJkqdUoeVRLLIoOyhCLjDdtjLqoNSnxIOBDXFrkleDvxC
R4KKsAtk65D2iah/u6R6nF/DDf3vMkxkm5uP5vvcnmY3QJC/17sQTmSK8OEpE9H4oTY/Cq41tYOD
8wneSdmp9mEknMYQjZLRHIptYDmsQ7aQ9GwWzOGNbFQ+hvxHenekCYRdfK6Pu0Wl7e10ziBNaUoQ
QQjzxPOuRv/AwgvUHdBX05voM3u7/FX71ehhFIz38yPrAf3/krGh85lgUhp6wuwp8kLxFwcwwZFL
MWCnM8hUG6kN8hvvOfa/FnPf8dvefWVJJWeNJQhgLTUStWIJxHDyxWsWrPbQNX0bYVtbzDt4Cof7
lhmGSWFs9RoYyQf1Zo/ny9lRrZdQNi+RAkUVh6ZjJx+ef0Kqx4Y2dj0ZYPCvsfKPSOXqyzuHbhNA
kPstlZvVAA2bgoN05YLBUWvgFDLal8ZjiLERfLH7lOXON/Eh2zivwX+GHNzq1SSmYuKmUneERBrY
3axosSX56ryQ1CzxnQ4loHwaZS5TjV0ZARrUIU+puZaEreDWBMOcSo6EWHjb3OlKYnCtJi62RtnK
kv1K3n/vvMVs8lRyzyWXV2BRdjgj6seFwr0xnYotislDJeytYKqRuaH0HxhNnctvJR8+xpo2EBAa
PumTPILGB0RWc0aJWsn3UMvwzSGndy83D1A/nTZoGya6/8zsRdIDkU8VCc/MHTmywP6HYxF9oKg0
Wp8mRJQP+tpp65tiYy0yY3r+kI3TlWSKQ+oD+7FYKDU9TmHNJDSATRvBejiUgQWnXzlrGS8GBvkD
p+QzT4D7jc6eKH0xOBgpZRxpW9OeC1XFr1b/nS8UUzVGW/UMsHIw1U8v96THY4L81RbZgeumFs3f
+UkJ/7gXolAiJkHRbErT5ZNdiIimLpKMLoSWyAxGdVab/xOwxgDuItC2FMMQ6Qh4nWlg8sgZPRJH
p4UUWrpyIIu1Cx/RLURhxHZ0Vmn+Ex5OM+sYxNX8mlB+uDnMG8OMHnuGVBNZqp+FGmkqVCkyf3ZI
rA8h6yarTSjFHqKeuMrxS2SMEuDRTh66I6deZMQDERcZ0ovcl5/FOoeoAUpHfL63kVr0SdJZyHdD
miDynvTtqoKxmPg4Rik2H/Xf1/OqjSz7Ive5dFLzH7AWoyf3G1eK/qJumdRwExPePRInzr5HLlEt
ML5sqK6ixFK7EEWePlNRTb4+G2i1FPTVkvhx5DicZFVLkZ3VCCE0YXKZShL4KWJpPmthlsj1lWVs
Ggh5j3YG2g/t+4RaYL8fb/oRSghjN5pgLGJUo+ejIqMnJkN5oZK0M5ZKxJDivS8P081xAMzc8sLr
FYd9BmqKNhWiXFOky3g6tEA3NaGysRZM8uAStCMR3LFBsVHnYyt+ihDIgdgeWBKxM3pCumWL248z
hLWsv4ScfR+0d9vMI0qXKA9WN7baAiCS6xh8EMkyfO3BCL/I43l0BTdmldwvlLAJNiBSin+miWmo
6xqNHb0P3X1z1RjnQT0DEXZoXskW4cfRr2XfciNsbl9zRgaCyPg3GLR4tLEluTzEVrAsEmRxTAny
XbAUe4ZobjDeio0AT+5ATtK2ZUL3enASs78ZjCVrvmjk/SuM9IE0yEsB/jRpK22xcN1Uv4BKKcFL
sfAbZfkwq1yL39ny7lImp5AKx8h8dSCXRESzG90jc5b7QaAjdoHpoMjA44OBT3cUIIDdIZk5TC3W
491cuklvRtdwFrFVGCzpfOPNvPYqLamQjW9I4rFECfN/xZMpKoZn+kejB/zFOQdB+F55HLdFI/90
9FRptoJB+ybwIBUAb2PiyOvWYs+U9a6SfwPk1pEM5kgb/pkOLfg7S43PXW7oIH/Q+gChlx/kknnr
M4N5BBXpX9naVUycPQxfPYRK8NFUKIUfCaqlgK6zeFC2zJLyKOMtS0TRHbwntoViiwUjWNY8IRCp
B8BlFyhaNkmKWX2S7Nd7sGNxduWEKr8nBuLupHSgz3ZyO4sL5QUX4D9Oakd3IfIPVVn8m85jnNRn
UO2yjVBigLVQbWf1jrF1DDnsoM+HR18W/OWLBDMRXWQ/a07Vf5tMvJS94VEqOEr3pD2qbCg2lr3J
qyKyLBlfV+q5LqmMEzEEqJa6MiIxjOH1f01ntkUuLJqhKiIXModLQMDyFeOC743lx+SUgWZo72Pc
xRs6pij8O+KXwOK3GPneJY3Vlt90Fab1IiXghxSN9nMvVIQtf7Rn8gqA5dsqWfStmVcLBot3I1dt
ijkvJ1CnuIVEIt+XVAkjvBdVOlomx378Udzip5encrUyTe1PucdoU3ah2L5Lu62xb6C9n3iOPF8W
wCFgSoikpvBeBGFrMYld9NgxMyZju/orrfxCvHyQcm9lmhLYHH89gzXUnBa8L7dcocFLVB5njQ/C
TBWcwyN6tW8YcGK8b1Hu6IUuIe6bgHDei7izf8kmOsBCgmbVGftSeLOOQOmWm0eIzMnH7bpGNkse
rA6XdIb58FCblm9UuZBG7Q+QSjoiuetHKRyWcUb8KH4O2PhCtUYgnyAOTlW4lIITgPC1IWHh9HHp
cDbt0/7+im+pIMohV5+tiX4PkL5Yrjd1rSeUKRc4MFG3ScLBC2C4pmeXEb0GTm3Cb3YP3MsQXUh3
O1V3LK/M/sge4j1PaAjU9QW2MG2qLl9cVLOicupaA3xjsS74UvagKRmfJhVuMHHxXJPJIgqu/PXL
B0GtBCV5/DjG6xaPAWrTfEv/0/3dLq9Bw+D65fSy84nolKWkRGhMxt4O4bvHjoSlpjzTLZx8MRwQ
r+pDAfTQaOp048TZYoi83+PtccAcAiHxEtOOUOpx3RIfhArtg0zwpJp5akDe6Nt9vHPvpJ2A8o3l
WWalxrXjGFxJqghJq7+eeFpzCPqpFj3p5TkJlTFMWyTqdSfInUVVy9xL/ApjYUK6jZQPwuA7nBYS
v3P8ggPbKxqFoMvOEl5ksVtsHfABeHUTyUvvo1ik59iWEe63oJOz5C5Zyup6fFKJE8p1Jvq6KP3+
dF+eOzkzzGpE21xG33c0giNFngoMie/6aJQVaBo1v0SkYBl+aTqmZ2/Gal2skCIMFukbSymnf19R
tAo1yfzo1BI+b3h/XrV54liWy6XO69QZUIUW14roZ/286SJaslpm7ezbPDgD7RkDh6TiDp/cgh/a
dtYd796AxfxMtS70iW1/a1+8jCeDLypv6c1/F3mz4ErMsiz/o+MIh5YilDTtmlMGnsWn9I3+O78m
XaNPQhnXSr0xHG0guTpoZ5rtypw0jdtB+qURjSyg1s3bwJ1qRZK2hWXvli+kxjeoaOkVMXybxCpa
c4QeHA7sRKjlCblG9GjXsWAKRxns5ddVGOiG0MkFeEFUmkjeXzrjUNQ7GtYEfS2NrC2ku3tZIQGD
xE7WloagA6jqQsDySMxW/H9NrX60b0y2VbDoXQc12R5FKj49epIsZ+FBCiBQmoS5TA/ndmvcEw1z
+qjjdMeoXKdAhm2kIHjgLY7hDvRq7U/h0X7RU0PaKb8X5J9U+Vge9whfrYLvg7aRuQSd4gXq+rtz
yBd2xO74VigjB24vsFK8G7ntNYsXzEmV4GD3UTlaeg3V1j8el9dSd4E5Mgx30t0nWbqVbYxDKjb8
Qb0nBa/+kk73IFwQf1ZhlhZ5iVvwannCkjTI/LQNSGmLtyGt20vc8Wj7juEmNrR48yNdIL6pMYGs
5uGiP/MBbEdXDZj9LKcvfrh3LzmkYO3llvxaYZip6eCt2fpvz0vySD4I8V87dizcGqeQBf3KrM6c
BW8hOFmAxRBbVzVsi08Vn7ldnQojJ/HfayqtR6srynbLMFEfj0Bu5XbEoVT861zBsAKhtbgd5syK
qRUULmer1+bPeNxbNoqPFHYyuy8kzWE7LwlVOTRvkrjZCC1FQ43NMfB8OtcAmKn8kNFva6lyk3If
WI9CYAeTWtDRxjMIzUivkK0O1+v8uSpClaPrh7tfByCxqCAlDOBhjdZAxSVS+qKW4vxUpZvyKQ5B
yABsrX2l6by6lj7otGAV3x1/eYGkayAuJ8mQtATFvinfhKgR9CiVvflXtEVm9G1o3sNvyfqnhMAg
Kdyiby6lv8gn5CMSKcMk8e4F8lZMJQO130s7pE/M+ZVqHHu+Jb3kbZ0my7MTKNTnZBj36C2vdtFY
CdkneXLeTdFIXhKKEx2/k6mqsjZd5Ynpu4xrv8P+90qqprv4yz+n83Yh8tvL9SY93lR783iCPP8A
60P3srh+mmKKyqnJrkt9OUyWp3YdfdFGDRwKfsojNfTeAap2QJZVuXIMDBk/LtoqSWKjXCcU7hsU
zwBeAmOsVfdqhvrQbWYWj32MIjJk+TLz2L2FHiRxcGqOZ3vu37V+Mm+801EEeQkCipiyXq+ahvuz
cmkIKtTLCfjYGasljIoqDDNNKcyr4bYHYm8I4OQMi13JQQ+G7hcWuWx31y5Xz5HWNcF54MPVJUi+
7lDonan0WojVOMdla7L/mSIm6FfguyyOFHrdGn5111fDIeQXQhb5qsSmd16Q1VDYCV/i2DwFyXEe
wzOqx7x0OyksluHa1/tAggD9ZrIsR5za5FeEImasZP/ECyFIqPeZ5ehmOrE8LqItI8UeImSFv+Wd
B9gAxR3QHg3bWwgd89SRMM1Xn9R5FppGAa0pdsBpy+5faGLVJdmHr4sZ00pE97E3pvZm8AgivlVX
IC6ubx2VUq45/AP/hLf4gNpTAWMs+lvhzZWO24koGgkRJrrdDn2utLtrtKp+PAc0nar5WKEOFfwz
OAcUOTQut7DqEs91BoTAIInIrakzqUUs9jWSbyf5BILH6VEpjtDDKGzlNzkN7BpvCjOZNI8tSwO1
EAtZuFPDikfRY0vm0BANYRoXfQgW9l7lK8EELZhLNmvILaYjdqjCcZ4llSOuqPxU4qGYNogIjkyp
NWwOZnsc3f4mq13ioPcHiOc93cPjwx+i/hBmkJdI/Y4KxZMXtjrDqRGSG575sV991PJ+6Dlstydw
Re7suNakVOkwr9V4te9F6ICWxS/p8RORZoCF65K0jz8F9ejlhN9W04tt/onnrU1oLT0Q+JOjhM/d
iCg8sXbbi3Lz0z5nQckbkSZTD0LlVHVAhiLt9WI7AWrgs1Ig/5OoAdbUKj7GyCtEgMLQItFRR0JY
Tl2ACcMDLxWHMGkbys2HxLj9Cyu6T3e4NtNBy5y/VPNKeStw/f3qKVUyBrZjRjFqvCxZeAOQTGUz
Xa/Cp4MHkiMx12WClXWm1eDJ+RX2qfGsqX/og25yrSluQ+5H0c86F6dGux7q4Bxm5Q+r3L/eL080
2XpMLMaldjfSs8vVVs2PUdW7jSNuNqOhS70m0PZj3Wv2FhEBdX6RhcX0L9Up1wJnrdkPSNmVgRn/
9cjq0d7u5pvSSFnasgiOQ2ulpxW6AA/oxEIRI4XYG41db5qhzNlNLLFWhOsUOs7m4OsowWOmFOu+
6n7v2swAycybq+QBKJp7i+AJ5Kx0rV1J7kc3FHuq9L7eiLQ8VrRwH81Hfv+8RJRwuCKipr4sC2R8
dHl/wJrbdCxoDW8cIQ+fCzanQzJlDBFT6fNGS0vOT1ILcFP1OEX/DRn7gz3KPiZIT+eqhQJwgrHf
sM07jjHlkqMqpMvmyzx6XezX3dOOMk89Zo6+3orb6xRMU9EzoPQ13+gEBpa9MRNYEon+5NGYg3Ju
p60o5b0LH+I08RcsZNVvongbZl5mBiy5kXzxHYenzXectTBNzAfOSED5aFK9Tis3rJE4KdVwLQUW
mmsPWKGQ50ENWFCznPriO4LRYN/24hpd4OsGEZc8d3UUp/vsAKU5ppst+trZ0Cex0LirrwW4MGQg
U95Nks7gdhSlyLQVF6y6sMnP/2a6mxP/W6JzW/b1u8n+Pc6udiQgUoItyiyaSekeb5+4DHYX+twd
XWUuDX8BfFYlZ3MDuyoRei3DHWoBseQX33VxRUXoR8VnsUw5u+vclwZSqAOP8iuxxnBwZdnpvsqk
K2xfWEfrl0s+yWXKF0OrCY39e96t7+vxApSC02K/ibMxidv7PDYj7YMnMFPP2E0KawCRXetyozZC
5OMnBlJGjfyTG6Gyc4pQLUIAnLlVNxUMIG79dQK86Z0Qr9fHxgoS6brdJNU5LrGYsAwB052oG6Vk
sElE48Qu1sO0u3LmaHCu/uVTU/aRj4FdSBNlAhQsMSwDlKRK8hvKoG3HBtIUApQ9aEOJpt0JBQLq
G/LaDU20x9iLJP2Z+hs4GgAYmFKaiqqaE6QocVGcSRNinylu44MPlmeVCfxcObVPkNUVjH+91JYv
4mkMPVxwAMuarxgXbsvdTETi3lv8wUBLBPJ4QVHTvRkLCYd6LYpz54pQ28HuT2IUm0v2QnY4FYlP
clPFElFusIay3onkfF/quF9jMloG65bZkYwvkc4CIkRb1EgIQBir6kXb8352hiHij0FIfcEKfIV1
z6ZixxNMUawJdqk9i1G9yAuP2W3/8FHUoQccZU50Izc3Nchx7G50kdvnvU2xYiz9RkVDRXlt4Jt+
iScH8ghrSOthB7+E9tIULq36XGvs7jhgEaGSb7uzqEHeC1McWjKaZc95j6/6UxA+IPRmzEbflZj7
7Kl+6XkLaLO2sm2OYXNVF6jK08CspgG5rI2gb0bCAT4EoFH99kvN4buroxiVI/ZeKww0G8msFwmc
SF+PLiKbR6tB+duxanL/U5ktCFoj4MjFA4dSTn2oOuv7LqFS1JGn+8mNu7GJIl9qIaLnUyqYG9et
X1eN7Q5gcqc6qjbvDucmJSgyvysnHP/vM7RQzP6zu/85rrfQBiFmzDfdPRUZCoqJ66Q7+KOf8gLo
3Snxi+ITW4xBYrburfsydjQMw/a3ROX3JefFjk5lzEH2XajT3PSdW8r/+KmJ8S0T09Z+RcK6iIMg
YnQQShVDuF2pwr+LxnNFfmJnggbY4FHCXAJWLwAXi5emuHaOkkF/zGHrEx5D5RtJvvgcdZZlaxgg
povnzRlUFJ6azJuMpjDhR/ziy6SsRQEyagIOYp+8dKWue5zNgE7HN6i/HUvytGAaGS5MWvqw+PxF
cCeQwzhnP4EfcqZuuZl31z3UE7XofSQYV+/+BrdNj6ZpsCaPdQZf1JF4Ec+YzsUOpvOrhMQf9fRv
RoWyYcAT3bm2AZAVs7VgqI8PmhvSSU/JgZcX5A90Pk2g4dWB2tSXI5ChLupgxdbFd4utYOKY2lpt
mQuQ3ucVzYSmT1TH6776bA4FUDK8/1D22vCSTh/odgz4R2yGYH9psdw+T4ZNs44Fso5Zd3biUxPY
okNO8uwAjdomCbaBonr6w4WvLIpSNeZmCkopa5nodUKop29tUSu2CsxWRnDIw0l0himzZ1NyUODP
XMPkNDM+O887CxBMaSVt3TPIORTPLjzA4LaET/ckRH9uCbpWEzKriNk2Rvr3RiK96Siw9/jXNcBY
4kLm8EwfbNCb+cnmP69z9HOky0KmMA2oTj+WjoPX565EY2dV0MEAerpq972Qul1r8KBblyEBgpzc
JMlQVhmAYrq+TSNT2pWfw6foqdzJREL+nilt+Q67lisXsrX/s1ANoqLHUsa6xxVuBTUcLVzHdiys
SM3yEBU/GpNzX6w6fe0agzEUmKps5tRViCk8oHpeKAXfoC7WqmZ252IkGYjREuNueFDHdDzjs+GJ
nhpBCbofWDGuDi2Tkvl8/u6r/YDhBNV22yWakISAnun7bjqBIU2fJSuh1UVMncsIO/N8A10WxkH/
jE5S2AesQLWWPiKyiKChFdfDma3MtsCSEOsP/XHWdjCGoP9LCgGtS6VE4SV8m/hpa1t4EZZN36hk
eoYD9IcYhxnc52VlGbRt9IH1bW5b2YitURBBmOeCq5R2DKQmmA+PiY2tzdVNDi6Kj6YBxNDTUH1D
bRmd+2q5FH/K5oqqNnhAy8RKjsrnBxw3SQgzaQOyvKNHWvRsZwuWY6c+0rsb7zfPCm+H0OqJibTV
dmcVmquXa4Yea9XYPo3ET+6ecsCB7AkJs67Lxwg1vQLyBhS8eSjl+grS0YXkV9AX9KdU6nZm6rpp
rHhjPfTb4FzvFZIi+ct304GcrbocGe3oBqhbPn3DeqdRmTpZkpCBYP7ROFxwOAvVcJ1LnCiz8CCl
a7NqV5zMynuYYflNq3qPQvAR8+ZjBgtt50oz4I5Fis6r4Ujgpdm3FKARk7NEFN68b/5QiXz5yeye
cLruU37pnPYgomemIrD6QfbhsHX50J9uSvmoLikeYvZhrKOiQvAN0rZ7rYW5aYfOu4mXVGTkZc0V
/eenoe+izvObD4dFjFiOUnZ1mgdOwpRV6tfYGUxMNxE97xRKcDZ7bCzgHz8e41HucbKcKn0f10hY
Y7u0iSnoMBcgoFhMzIW7pzrUUcg4956++yqhbtZaWho6rIYgrFdK7zwpkxCaBplwKsXvyOCfY0eY
MEXNAQ39dyGSfKAYji557iSvCvWl3q3gFEGrH5KKOrhkgXzkQmMMcrPuTpsZU/MpSw0mYx8Oty1s
RhIGSbMHGdHbOhjYdi60VT2G6CPwjj9yBrVahtRkE7+w7kZ5msdJNRTq164Ekppr4CqwWqVrL405
vl2v3sYklqFYNI0Mcljqm/GgFCilvFQaXO+Ow+iFQESGNVF2B9XpMuX3rIdooPbUGSFtBSvLszuy
r8UHfKy4Lad22/hwyN1yEUe+8JF6Hon3rT03aMqRZbGFoM6QZc8pEKlgs9LxtSp2k7mRiYfcVjIn
vAFNtL80Ed/PmCi5oup1k9YAn3vpTjCz5i4uZICbBG/FVsWRWkP3IuOKDv+YwfbKFyMJzlzoxZ4d
yrBkr35kv1NELMmMaCAIfEa/qhkdwLlnnnERiYlquf0hvCHbBRWOPx22nMk4g4baO6n5fPSaThJB
n6yZfc/7hN+fgOc3uadGSkVMlVuNXqhzlxZt+ByLX+1zXZVhGEQvCBTAzWiQCDrftE/P3vcQkLOB
n75QP0p9oouN0BzarkCd53uJ9oRn6KxNej3kf3Ggu39/QsMrefyJa1Dzr9N7s1tYiRIs4fbGQN+N
Oz6csI+Ed3n7Pf8QreaatXhbgYDgiMBlf39BpMxFLVmEwM73nrhDDers9kHZwtqFwSGn9pRnt/g5
0TQduoOU+pdHITiUqm1gfJ405+KU6bwn6w7Hj8CDsYmbrouTzPnmC6ig2m1DH4uCNgFX5ORGtBva
4pQVrb1D6f4Soj2wJjd8De/J3SJu1ezhLeHXfNR7Kj9Viw6stlnHByg6OZDT5s4G+WmrfecZnCuJ
zjz4BRHiXocKmqs5WRLohoizjsVv7j/P+9hfIGIT05tLG+6zNHfBNSbmecwf4WNBaw4/JQYdvFWr
MVSEHual+/+fB76okruq9sbaRnlqFz83LpEGpnrFOSlHe5Yk85aWgk0yGn2ljrNhmq8t9wbfxbTt
yQ63hhxEw2e727NkGwZCFDWqOdT6EDR1fHZ2pZ0yQ2JEaOvc+laPR3TnjWHbjzk6A36E2kRx8HjN
3CYs+SmGt7P1FCTVHedkqlJeFOwGUKrVc5HThlo+BUmftsikFmH0kmvT3X8vFyNJ1AzAgTIpu68j
hCK35DUS9E1H9go2tW1STfeTH4MEv3b1CPaP6TCq4G7C7em+BArHZ9OjWtoh1NMDsXo5GdVxdp53
i4Qhepm2kpNr6UTWOW/6OqMnE//dJsHuK07hv7rem4FJsfYhkn0a2YND+EZMN0GELLNlljo0NnOE
zstEs9QoE7qpaNQL1gE0Mqh0TU3L0k+v1qFE1kF8tbPyQ+HVsL1JWllBjO8XIWyBR+kZarAkSXJW
USqBLFVLGYlshe3ZmzgC4Doh3uW31b3Fo7bkCdDPP3COURt+Q9/4rX/ydusLG34+02wcUSd17o/Q
4R0iYy0fywHLohBLlBl3ozDRFXUfxL8WTlbJeQugN/HcK4jyYOK4xvturwjxwhfm0OAA3hWntEwE
kpM0j5gtueLZZuBWjCfvJbhSbJSb5xwv8uMQx+LG+ClyVfe9FtJrEJMr1qzSKZlVnFV1FIKVCwgX
eNUUBMTXA47id1loZV4ee2uc7XX6BUcXCWOsdipH390APkNILuejL3qo1BZEf/chMgyrjTUYEibm
iBSjGYZouN8LkTp+sd5lYnUmby8QRErJSZZFzv2oG4VV5ay6D6YVFAwVvHfLLMtvF06ZoV1Oxrbf
oQ/+Zz0a9ncxmOU5HAA6o8zE0jqqEWWE3eSTenTx3DHDAwihtKNrIVCvEDoOD5uerCaceZgDuOnc
RtpyiTXbRpjlG3JSYg+vNYIXISEt6XjgBuZEgy03ztv9/Fp/LT5MMR/aBcY41SjQinBD40szg7kK
Dpu5MSIgzAUGrBxWPzbjTQvZtLKWT+W/exg4f9/G/WU7Vn457WryI7IoECBxEDkrLZoI40TTsYbG
SRExQQg20/4eeYwkbpM2ecPX1lF5xpIBqvgNCjZmmxlFF4/l0Sl5vVZVevXHfjpogNUo/ugL6bKr
ulV0wD9CfYcDMNXJCt95FLX8JzkSIir7kU/I3zNQ6SVKcfVItpG96lngirsjpckA4WZdxH9EiBsz
5P3ePBCyxAWMfTuPetga36ZYOrhWdPflvCFLMWQlSjqcQLuRaKNZZpW43p9vfbcZ8jQpTsbIFqPI
0PjDQ03Bx30h78vnDa2epwXoGKK3zFiDHUkAJR5dhafW3AE02RogmzyhMpO7dtLub+sn84U4X7Bu
y/z9aRTvJBkQ8oIxtIdBmt4OyxOxHeOw8+FaaTZEX0t4ieR7meyEAeFQzyw7OAWczhaVYKImDCyI
MDlm5vLw58OxHjiE9KwG/fH80Pk8cFAHWltQsWaMTSfq9Lyi1kKtzeW/yT4jFRjkB5/Y/J16nXs4
w1gVDRLRoaf7Auda+WWxsxQ9AXdwiNVgeqtlzP/XAhjXm+ZwjpY1lA4waa8dXhOvM//dSuejevVr
LaaxFkH0jRdWJJHlmJo5mFcHp6rQVlntVc45/1gOUwZKLN3L/WT93sAQ2n2CluCVPuJsHQvdBsPS
Oes6sr4tggiNaljJGQSb49CW/NO4McBcDEQJVzsIy8/1a5D84JURuesqICadf5oeEwRPwhgxUYqk
4iaEjKgO/1NDAyiqxkgA4W8FdAv0icQoLUmLpOlCZIegv8gSq8pGuNs90LSIDgaDTiBrDKauek5B
puywPtp9nMwCzG5sSW8akzdnRj4g79V2Y4CDtq4dM4tOQWlXEtt+alv3NZbxZV4DBGOqkZGzokuC
+QfxYMQjXXRkZHO+fpAPttWfsZnBALNT0BSx8JTlwn7vYcVsmd+9U39ZaANtOw0jlqo8IfchBA+Q
uxcs5gnKlpDp4EIKl9VNADAdR0b6pZ8sqLZKtnpYYqZcUqvz9sG0qXvhBlhPWA+H2lu+DVexnD44
EeBFBAbCTLkSEkjfFIGM2zz7o+PestFBNv4CvCA7f5ZCmg0HQ5qESCZo5+NvEsVu+pYTwgtZYrY5
AJSPB28o6ZayoALIoDD9GmzlsiieDM6JULLz66Ug/FvjtCyVE71rL0OxTRlX3GzK2p7YIO4yJAOq
6NXC/JoS2k/l7QHSf7HI7PSZGh3f9j+WTfqOGgB5mZTma3Ce3OBJk8JrmFAM9BwweW1KqvtksDCQ
IdXyR1DHdhP0HfpcN3Bj1HrlPA4npb85i4nt7KAf4qfdPKhF3eLPNmz44urPRbkchBklbDITJEO+
RLrrnWqEKUbDHLHMgRk4sRb83dHB8fzffVXgTgxURLaZhadkxebPOuQ/W37CKJOpqInwPpC2CtEX
/96enwQQJF3rJ1ZVjiK/5j0GWh87AddpHf+EFf7kNMVDE1PeVeCkIe8/ESIg0BEy6v9nK7g/fYFp
FglQdGyti1lYWtN9VYqijgnGXPzl29wIBrpCabQn9KhYVBHJ38oTNOBLhlHDV9A01jP6KDIYYVY/
DgtdZ6qGSOKmBwGm5v2gli+RSS0McuTzON+8k9CrYgzpdgynvTTdxUe0wZCWnC5C+/77HgmyaETg
/djNRmyk8UiD68agyg5tucZlzuEgq3UScxpqP0ehX7rjXca29h4TskeQJ1dMTKKVDzN+3YC+AtZU
Eskq42w1rP3cKzS2+PdW25wJZMY5gVldm3oYYLuEQY0t4UTMSSWuxPYGodI+728ivgxenJ4GnoYb
yLnBBNnIINBNnMrGdHccCJKo/410TbXS48ER3BJ9UyPxVROKlIJhzwl5HcI8kgIiyVEbfyyDMIrd
SeNqZ+PVPkG0ErPDk93N/d1Au8odl2VP7GFzUkLO/9gY93VbAgUGX5IjK0DHxg42Est2hLdkdbsO
rcns6U0pHlL921YFVk9lQdXLXQCzwkLBs+5cFh8HeJJIrd3x8H/wO3lFs1QC6/ck/zf/R1kCYfFS
xvvnaky3Y08OQN0eaTEXS7gVeOqzLRhjLHtnn7iqdQ7VxCKtSDBi4E4WbfVbBErs5HabOOFYXJer
QxtCEUIgw0tdiAGSLmT9x9aTlnQ8RqcIgEKDRM0jGyPIiEUOdxm+DMwGnq3IYYsvQVqN4KAAWWyz
ngqdMHwpIBcpgHx5JSmJBE0CMgbZSv7iO+/8Im7cZiDw4r1UhwcjFNRiJHv3RMq26j/IqTXmy0Ft
VbLeNl5kVDMGzbiCQotwrAQXxoYFjih4KIVzT7A7dENNbooGgeg0jLvGvrevxio7G3jSzyBlLWGu
v8CifUP3SAq58RD/Wa/2yWVC6HTg9RUlLWdFtTCcpHuvuCO7QLAfPrRWskl8mFlzHLghdCKMo4lj
mSsyoajEscO/TmgDyym/QU3jYyC1nKKEanWik9z7Sqg264hHjaOXKyUnY7o18dTMFOl9UYdJqt0Z
gSgmSQNhRZDMTMbf8xU6HuCvnZmh6zOijyNHjyCOCMpxkHPnubWuo8D7WOoYp9Pcj3dfAPrCDI6j
Z78ojmvczjB6fjkfyLNW0+i1RASmoz/R/1G26shJjWBvdwvW37ZTt4HkMmz15MPr+DBF+DnIwTgr
cvKrp89wJIx4vt4JHJdWyU1zfvQbe3QVwl99Ng6RaQ1D/MN8YZLH7OOYReJYscQX4aIgGPiJlgNa
4uqmb36klzqu2k1F1x8PECIktpR6XY8vo0fvVPSPuRKPZZOFZsxUoj3KnYO0Zf/x4ARWkBbC6WSK
Xqqv6TF1ZwaKwxax1Y8N0aG+MoxbJVj3A+Qhudfh/Nh6HL7FEmFnGYMFy83+LSUPI1KnMfo4Kqyx
kwnV01yWKt7hAqidwOSEkrBI1RvCqiRNZCWG2BzJq29wQ4s9JjdDf65ZmXEpQqap4T+Bs41s1n4a
FBX0eSqxuhf5VwGKv+W3EISIUF6GasLN2WFy9CLU4tZ3rhEJlvMuIF3XNoHOs27nHgijc3nWjj76
Jt9w9hH9dQe4LZzDq0yeI1O+vTR626egO6mjcF4IJY8XcZRP96RBPKH5M5FWxHgs9gc6z08jTWzq
1d1PclZXaRGBXY4Vl8NV6fQHrJTA8b4DgQ/WAYK8LqPqWAKfzHFa46SFrEa4BwDtaV/Vam/HoLMf
SVsnYY8Kvmg/4xOymVhsIc5W2KBbpNK+QOX3nF8rDUlP5JTkmaRknZctxvbEijAfBMZv5iZBydTR
yfID80WFOma7gsWFWhbexiTOnzmnlKT0Jk0nqRMvvY7o+4QYqw1Ijdq39fqB0UQnAU+Cf1TZNjnU
cMvbrEgwpyKylviPAjKIsKLiJtVK0U3OgIF/n4TVgGSXCheMfTse18myeJtN9hAxgoQd/m5WowEv
bbkA3hCMsnil4KyQg3nXtXVP3WZOmBHWp9hFLqoerL5nvL4jKxQeIIBsem0yV6PR1Yf26QgWyV6q
P/eCM7gKFt9Fs7mink82vG5waEa3fdtkyKjNAzIzd9ultN6NJYmubRKwVh5rz3q04h/bP8jOzmt0
njCzyT6gkS28VWvipt/t7juPgSsOXiOUc4AmS8sLSKyjH0HWLCrOBoXw3dcxJT2yp9PwRKxwSfcJ
us7p2y/z7wYeIYijiAzcs4yKWq/Waw5gW7So9IfDMAJjLcqjw5wC1u22qGKq2mV5KnrUzA4vqIFm
v87s0MPfM0RPuD2f8RxQAR0hlT73fiklydjJ3huq16A59XO4IWCxGPuk5YPX6qaxM+pvsJDSIaQ1
Mvmh8cnTBj8hFoMfvuJYK6Lfk4V0DRJ7/euOqdWqKQFNsmXYYsUyYOM1gcoJ20G2DlWIKY6/nhu/
lhGMb6uwcS86MW11W5DWVJFjEe4BDuGVamFY/WbdaoRqYra3p0iSdhCeAtd6GBIwRSqsGZmdI2ak
u+k+uZ6Rysm4QZsf+wYSG0wlQFgNysk7QmFPRlrudurOJ+NLbXP8rCLrTy7fAVqbgdEPrdwY9QMe
51M3c+1x97OtU87srrP9WDkaoWGNWlJv/xRQq9s+XUf2lRKYpn49taRSDUcf2mOaq8F3abpRhlS1
wqMnVbJaXQHlePe+TxjnN8/q+ztzLVy2O3KPKsl8jFinhrYMaTIl63qAbqWSh/jqQW2KWFvVi4jL
xJ+fiZbeaEHNZ2E1YeO/qKsc9+n7LvikdtachZGm3IiQDrhj+ZE1MEiSBi8UxtfPjLj1KJon72BH
C5fNViJNtybVvS/TyDnq7mypsmKbF1lpQHjuwL9jOhoABehhOHvee0n2xcuLUxdGWiEEPLUvb1qh
dD11eJkdiG0UGUJGy0sNE4hG2z25qR+ED+ePlUcoripOSFyO6nGOFFbYUCtoou+yDoopnayPTgQb
/TzOmFyd4AtfBlV8vFFOGmcdtXtSvAeRDI6kmFV+Z73c2CLZrtpSERQiub/K+h+MvqTtWGAjiUlp
iIK67I6987mdJ/UIJ0OKH4ynprp1RhtpO5ZQh4fckiQLlaEULapi93xRS5r4SltL+UDpQgmKzlsJ
f6sSraIlddihGO6oPdaVLd/lKkQTrpVhFOBgyMfGXB3Xlwk9wFIMTU5xlFZp6rtu0hQCeOhkdRK6
4fhBHcR87yjbYIaNoeZM02MbxqFoU1GgR96zwIcOBc2yr9CMFfVI99P63/7mSPvnZSqRS23ZTwmD
rtFZTDewR4CKU0Wkmg5LmwtwGv9FwvXYnI2N1qUTELomXNKtjieVJxTk7AzOeLtqVuT9r3i9Nxjq
nvUC1LQ78xDjARQt7TLw5cAA3BbYuSCDwoxmbSrWPgsTjTj+s4ut4eB1tp9yfB8AdWxr12K2suzj
+vlSt6TyfBKKd5QIg3sgU7k3SuXJtwlRMQA2c5v48TlwKpYhpCSwGf1ndAhAfpETFbyjPg3mXsyj
nZEf79EXXLGFLF8Xw6Kw7lZqGla3G53Ra8kZnKTfv1Do09/9W3JOmmm5S+rkTtCB3/1Z/eX/PQjC
reNsJfawS4nqZJ57B3+uRWOFp0YBKT5W4GhdE5LeDeKWSMWxlWN9S3WfmTIGh0SMbH3+AdA6mp/Q
j4OgSv1P4yjQtp4nShYCJ0DXHxYDW1e1WN5rj/vxxZfuB+p3QDi5Zn9swQx7o40lGbiaXvBrP9Su
EIq5A2bj4l487ij7TzSvF0VFAHACzJlJ7AXsVAmiJTYA8drUqpA0V/1NLKC5KGtd19Nxg4lquj3F
BZkz0bIyolx95M8J6XoO9iLvZthbJNJaMvoC5cQu2Hur0HdFnb+808psjiOSpweLKio9yGzaWfZV
TQE9T6vuDV+3vmVLVXV+AEmkr5HwBLFgCmSPAMorH9Pq/HntE8bysAzkaLy0sEjqTYLmUMTBozF1
q2Ib9p73GXTaPLnCY8HLi4cSzTsnuBVAH9Nky+iM+2IvLoiuOAIrChk1Sck2vGKStrqMDf0524QY
2PpCdCmAUIt2aYO14ski7Us72R7eeD1mcp8pCZJP/x1KCI1CSnwEVtfcDBo/AxRzfp17Bejk1Xvj
UB+maSzQI7wykL09/V2git47/2Am8VmJJGhdwGLvU6jECL/6MlmO+oNfDSuApKXKmtKQdcJerUWx
iqgqV9wXXcMN2rH9aweIUbErVLq/0fEFvvaXvb2F+ALyoXaKzcaBBXOZ7gyZWa+C/+NUBTFLx6HO
PAl+R3Se+hcrdNSVJXviwAJSdtdtNFC6zHpRWx72aTnuMdXYNRFooggLfF7f80+wM/ymjDVbYXtK
jR13mm86N8RgUxgY3Kv/uG/2e87n8hVajyIVibXxggD4yliO/mX3IK8zWti767bInq/IszBZCWzI
fSPxYiqgtwzl8Sc1TybWFn7d2PhH1++AWP6rETxOTUe9JNpaW5GyTOaZVXNiZEIEVcFqqJs2iST+
7LicIhFjiInnfhY80gev7E+vrdt+ajaRFjeeVT6wmGVsUkobGBfvjEkpkS8UYIMIuUtNATE+eEFB
9wzFeHKndN1xwemCMIS32pMzxTwOkjNztgRZpbNMS6XggHLczFm401tey30UpxUy6G9ASP4sgDSZ
Le2FwYnh3G3rlL8JqjDmsN0+zJvi9S4z8rsGg1Q9XgDP4bRiKCvf6/hE2ZqmNK/3pp+m+5dLhIxt
zdaZpKPVGupgGr6pJ6OPsWQnTUSCC69Pb6rT9a4eaOBnjV6+0CQpSuu/lIva2S4wV/QilJYMCzbu
rCgNcMlXyoCPztiO3JAK3F8T/wbytfUj1aIxjyXk84JM0cPWIKkwarnnA8/i4thWZgsAz5PymI/g
5dXPn88Vc1THUKBnIPIXfPWIAXTloUzASvCkG2ZcajdBqlAN1zuDjEqDh3azbJARA1fZ8q+6tD4x
VYF9NJo+/FvZKk1A/8V8QGS12w4T+ezqLCwvwVOW8BxQCLeuJHXIt7sbumzF5Ym2Uso9kiush6tC
e3hp6nCQuZEmv2UoET2UwA4LA8PFqjzevo0srHAKRAX+bX5wsrP68vUmf8zcf+57Y9fswL0HeWsR
J/MWySn41HAc6jciam817HNgYDTu4AjbfLs9ee1ZES+f4whJRCdoW40sEjOJ0IEkUqAYGnHjtZy1
aCXWth/+/NjcjRaURlWDO57PRWSOW+dBeoTUP5LgfKoPxti+Pt9wZay6Oj3KBXUXCNrEnWuo/Deo
YkthiTwNnK7pyt9SkHCkE7UbJMGqC2lHxnNvVu/lM+whLOYGqMxC3DAewnqpWTz0QmBwpei1NdY5
WsdiA3xHv7nLXqbEkRlq18rsQShT/pfAej4zLaewSgGOKRfXYQAkyvBIS0xGGuyF3AyE8kWcbhNR
EOkIjgJ0diVwxyTbx/hJ6EFNE3m7eWvjWgxWzVtGcvbVfwzQ0DzKfVBy6M7hc8t4fcnY/iVpxilk
Oaa/R0O2Fehso8FMtOTciWtqfy5VA720cNlLIq4xgTpXnVDk9S6ryndLAJBY56PiUPTMMhQUz3cX
y/P3cEUt5PVX2FOCuAGwFgfK1acZ0QCzzPKi2oB7EBWBgwiJ43+1F9Sd1CXC5yC4kcvnUUNHC3kU
s1r45Qr5ZlkK5eda6reFYiM2wPPMcrPqH69sCyfCRNztTGSO9WYunpPT9n33o2QuJrmq5HBkDLNw
1DZZGnsKLC0qOT0joskwRrrL8XjFyjdZu/8Yq0aIeYF08MB5uPKlfU0nruTq4q5IVEcBFO+1eY7N
SZD1iqlGRmPUfyOxjLCozKm2qMKn0/W22hIIGCwNxEC6NM93dC+1AdSAfJtXZLvODhiy4SND+/7M
Vuvyw1AaTi42dqKmSjuQhRgIzB5f0XsAGmPxOOLYg2yKBKvBX+15Nri5CalphTvp7KMbe/KLwEZ3
X529ebzRx/ISXgQgezutcO7c554tcIeVlrb3DbcOmjkV9HgNrOZhzISBfUco8ZDfdiXez0zCkZDI
52eG+uAQ0Sr4tIreX7DJQiEZkWxLVjKYtG6fbuPPtFvZO7MZVxzz+NeGXNjDqx9oD3RDgyM0/4Ej
cHbv5aXhQzMXHa5lgyWbDbSyZPgJJW2fLnbr/XWRmmHtw6VYoAkqcHKa65hJ0/BDutoFkSo9p2pv
2ORURCkuUuf9mzbVBCkSg/t9gSnBTYOqHGMBBKgzcqx4OlBT8g6CxJN2Y/qHmsOnRd5TYT1p1S/2
4v7pF/OuUZVv0kOKnj2nFwIlzlBfdzYvqbVnU4biMYclDdoYxpaMaGUkn8yXURvRyNk5JQ3tyCQI
gldz7GY6ydxvt4A+LBjOwGytwyv39khzpP6S+p/M+XJ30+ANTnMUWuqgNDGDCBWMKY9+F8tDVMxC
cAK0RVGtXgigmE+0+gjCNO2yKhx5Q0flCpd0YKNduSFfReFYe7PMuqTpWJJIkyNsfbziECiXnfql
xGqRZzADMFxfLIrfq8m4dPZ2dMMingzD1hBBwD0Qq8xOYBtrOjnwp3H1NJWgUmBertAch041js/6
95Qbx0GnmKwZQmq8nUPb5sg67A2MiuC26Qqn4mXxbeCJwekIYgEBWqOnrRvtcwYqo9/NeLA68GbJ
IwOkpWdERlxAnhZtsgtHKZWXsnFXmT7wQxuffHfGxSDhsiAsE0ZHPdLL6dhWcgHdoMHoqUBlw4zw
w0ggXgzcJFUTfk34a8nOj49Ua3NZOTKpcahBnSQgod8IwpXk8J51Je5H2oA7Y9M6jtsNVeRVDEyM
5it97xz1/IvyPvbESFiiDMcDab7rtInhP3sxTPNym4GLbZS0M2cjLMnc0GRg/+B60SPXx5/N5G8v
ssePN5RWEKgnzzbkB+qrrEeTgik99R8KMg0P1QeKIzISvrC5Vc5Y5GkLEtHVCJPpsrFgCTklTP6E
Y5PO3rYW1e+rjoZy0j9ZW9Jsw01JvgBW2dGdyMa3RGGk8B764sGo440DPtOmInT754llmToUbTec
CQcYp4dluYddc02Gg58xq2rl2j+s/njimtr0K9KY/TTSsSlkIcwMEYnQF8VVvgMMJBT698DemYSJ
EJvgsmjr2n5WbLTrLCxsG+mqohbLvZ1GeT/Qz3p8vIn8ycno5HQfi/HiFFCtPLWhPstePjxbZpu7
RoHBSvbYzxuSO9oBiwDev6c7iJHBalVqDZCogkFCqRXNQ9Lt+zRU/jWWe7RcCmxsa/tYjmvhu/Is
eCRt+n6lybrdk+RIr/vi0tvGu3bXiVUSQH9cdsSkyiv3jXP3HFhzE/YFeXF0XXealwnRt2b+6pwU
zCgQ9QDYGZLhhG5OgP9rlo+js/H9988m4AsLudfgBqHQSa0r4WX488UQPXzvNpPINgsZQwOLSZIn
DpXqNHnsOfEoc9v/ieQUJtoHYbjFsAr5oJhFqEz9fS1yhl0FfnyJ2JbzQ8Q81O6xvmBXSC+CgIUm
aRIMJKZwxP+hd/CWmQTbjgxEYmYSHmazSUsNtHBDtW4KIGYq21J892b5ZrBfCMuHOvbgL+25M+7R
3V8GpH7d3epB/aAPP1DjyqBMPLTKkHoKbhf3lPDNin+Ii8Vbg7coLIJP8+wVY/5J41LPFRgHkAnA
V7/Ab6HQ7xmHYrcxMzjCPDH3HEPP14qLIpqXZ3RXZMDm+bCmpJzonwjEhEoqHjtIxKxBUeN2g2r3
CHEV30XbzUX3MqwdYGLeZvtpqSiZ/91ocD3+5vzxXVBZBdVpwMAQDhO71lynkkl8lClEJfHPqQVr
P4xBvyCKoHY/OrSnaqZNF8AReBFYn9T/3M8Zbwcw/cjQeitQXf53gqreggoylS0PT02XFHEYAENz
FhP9BSrXp5Gpu8q9N1kUuxniSYyCxpbByHbA7QLbLSQWT8+Pk9AD/mO7Y3UalRWxyOL+baLvPtsC
6Z2o1/kH+A+d/6aldYU3ll95a9YJkY2tIF/1OsiECEZCo0HETjp8ZGYUXQ2c4Dnt9jXdALsmzp6s
mJJ85gEia9nFQofnqYyuuD3WoPXD83hg09FzRk9zWIB0i/y1MqDhbrTvY50irLBSSCwy0oJqqPTI
dWAOfzeQD0xN6j0cgH+ew4Ts0rlUZwrprXf4SUHVbSX35XDOsni++U3GC7BaBZaE1k+/+hGQFBlU
yjBPK4eEoPpy00EbyKpPM60u2S1gvOhGCDoYmJ7NFFfBZKUp4bIncJtZfr0iko4dLNH6UK3paRXd
tuYRd11jlWDr+5LydvNsXg7ITy0e4QpoT3uG339E7duUBDHfn4hMQywkzd9/9CAwwFISUOqau8y+
Wo9x2ZiAPdHAIjNKDk+L1N3G2V+UegypviNjgoyrmTTaIBHM6+AJdy5cZX1L5H7zaYR7wYLzwlce
6bHdc1AES1JJqMG+JV3Nsi1pkt+i4JCUR2wI/vVCSB+DINQ7ZHJQimnrjxKzJGW7VNld3XVyuWGk
ygciaBSAfS/oySA9Eel2Nrl+Bq39AfHdITtLpQ+oXeqLQi78TgV9Tho5aEMZrrBofUO/9nZ2DKLR
PNHxhH0jdAWp3z0Wf0vT0SVHqv/en09o3eNyWuqfrMDObui50TAqVFB+zoKbcznuilbE5pncTm11
oGwhjK485a/g+AuTR2O5g39ZHWyNAcy0rzLgVdKgqt0xQuQIhzl8vGxFLsrH1VcIOi1WNGrr1I2/
UT5as978l7gGHspw5gSiK09xXbN+fqFYk5ssYX0T5vEMzluSCdUilEcV4vC5RfP7RJvqlQR5Crnu
uIl7rTSyvH9YNhONOJiHn6FvoRxRTyYQqLlLLz6TADBqx4mSAy/8sy1mbuCuOFmxczA11EWahTmt
EuTrM+IQS1+8CnNaVtUkHIl7Evk4cx0bOhiuiwODbWP7/EcZrm+ZKhQe61HreCKMzgrQb1oXAuqo
SOMjZyNH6Orw8gCyszr0vEilFlL/T+beglzyVn4IBwc8qAPhD3gNgu+55EdVyKCVqB4eTexO1qOw
HUPSImawkvSpT1SFutjiZ+nUUp9S7ZblbK9zCKew3IHKA4JI45euLIaD4vE3YqFUDULQVj9du1gl
sJY2nEnLS/j9TmAgC78T86zUrfj7wjeDF1410CaCe1MF1q1fd1bUTNOpSuJoBmNub072C1HOZ8AJ
tXjLWZ4evJ/xvgwg7yMIOoq9pQSSVH8wlFRpaPYHqKAKywa9OMRppfNCLxtau60Vkv+yujrvAJPc
OjFFTOkN1TVwXgRga7YA3Hki/n2YR7M0fvHMbNrX+qzwzQdl/2du8CzVvPGFVHaH1qYr8Vtzfp/K
/Gk9+5904p5UNR1bgqi6cYLJhxpcAtbscRVRG+dCe+JOuIxfIj88UMPy/WVAcbyXv81I/M1mHCwf
oBhEwU+Wo0FWzmv7nCAboMK1CBG1LXWLDe4WdjnBsZAVDp41VpsL7ktgvU9KEuVgK7287ZuFHxim
1FNq5JVsSncnrHG97PrV5OIfpq7Y+0UmMJIXz45kiNvOKQzb+f6fwV6kyIUuHV9KFeVbvDQSKZFH
SlX/1FkmK+04+iIUjncNwbHnl0o2NHRPFz8Ji8XrbwxzDBYHRrgDeBALB/P/LkALgHGe72LoRo14
Hv6AgxMxKtg77h8vE+pfxkNhaMpBDpdbzDWiIKAL+qTjL5FqgElN6ilG9awzDJs5DXnlI2ndl170
RWGIv40ObaocZQ5uXRZC2+WuhN2Eo68K2nUjPzl22G5m4XgXDiTRn6UZySbxJD06hPOkD2mzbauP
jyej3ILZZQBWN5xQtpFvcnDbOjbBIac3t02WOO6AeMcgQBe6VYAARKM90A3zGGjkt7b3yiWE4VVA
yFeFLMiyS3/KAAMPvz1f8y0fFTTjvEBVsWNYKR/JXAtM7ZUPGpe0OMQcNJOHpljzHoFoUYsPqEAW
LdFxMN9X1HIlgs8as0vb+UyX9n7JZ3IBurQHzT5mSDKXb5liflG0blCQa2t7p9aNGFJ8ju9LnuRB
HqXD/sKWhgkxdwCiDFL3X6YJihuCHyd/b/4/Ad4Y6qDpvP+yDokLqm1DIeXd1Z+DkNkPy0Gd1WI3
X8EkBqsFA1kAz44QiccSb1oLE/mipc5bb22FsdPJiDAQQrK+fo/xICttlkXDSMepXTJCjM9II+YO
0vpotmqt4O05DBV3PjNiglGH7whASmKe7mJ7WAYPXeV9IOtks8juu5i71Jt84VGB3rVZnjxyIDxu
hnAor2N0xRV2qEGGlcbQHUZlnH/xAxvklx2HupUJHW3pBHXQism93qSrLXwJTXKbbj1dg0e1GLIx
9+LSP3m0np55tMQA2kzAwvZdu0S4H2hwGDKrbnGaTxzLhqUWCDVhkEa/r+qFJfndLIvxgTEE2NLO
/hL0wkMz5N1w1fODABUr9GBGHjs2l2WH5qzCMxYbWwBmhbnHUjkzC6lUNWXq70Ee8I9n66AjTzmo
/p4B/LsHc589NneEPE/g/NHH96/w97ldWkPilMFqAywVpuDO9HMK3nMAM9KjkyUQlRTyzyn5+9q1
BDz1jpM/w+GMlQNyktFwBAGUiJV3a0ZGGHpvv4xUANh2bCACZ+24vsV9z+V7O5Fp3IPk9xKM3yJ4
2V2TJzTrGoBazDJtsIoCemVG5jFYNkgHAseM8rvIYWVGvG+yCxdF6oWEvg2DMmeNwlcLUv79iczS
fgvEw8VHGjxySd2bxCPbWCVX5VQCsM3FAYEwupjwpBJMzKO0WftFhUiq3PZ08FjZ1nZo7fZ+RkW0
9nfZqA5aehbrJxcYOxrGA2XEH+1nXNvsMbsVTpfmMopHM0SESQB+T3NYOsUiUkRHF5zS1evOnsyS
AF6+O9dWZCX3XA85R4lA7Q7huZFv6SPDFCtdHJlxdc8rBRHnGgDDVjOsOIMiMfP53wsYj9q/OTfX
YOYkJF56iSe0nFjxMBE2iJEwdMW8VYvraOwnYTBbNYHZk1m3j13anFZfe9oI+FaAkkzxVnlYeWvB
yzXJ6sExedWxcwCHW5fX2G0xYJvLcSzCQpVTcSGwMI9MSV1GwBlGzM0vFhOfZqGwDXfovcQhIca8
z1rgWBD/pRF5agLtgFs83hRmqVRGRllRIs55qLoOL4nBZAOPaAydPsFmHQnzxbgPu35ObowTzAGd
/+FB9jeSKKIP+jX4d9kigvSGGjHioP1CiyCXvBMQurP7bbyYq1yyxCBWJEdGP3fGRAithxUKaXho
kDHrr2SkeNP5TsRsfBIKpMIIJYkDwnievHrjPAlktHPJepDZEiRHYpwRDfkcl3tcpOdTXtSqPcgh
RqDnb8nzRx8H/fkJT1dzfIDW8vKomCBcIUE77G326zJsrcUxjvo4WBUKjN9R1sZjRitJYBkTHP7z
QYpKdYnBvoUMZyddaiUIKPp3SUZyJu53bfgQDcr1fOGMejqfYX3nTEVsnz4drQfVMVbxLDP03NTe
/UIMZHDyLzM+xngiXwOS5AzxMiqwDDU8ZV6PCL6sNOjI0+SzbYHkfLvt/0Ae8HEjBL1QwcqqRQiQ
tadfRdH+ILi4vEjUnSygv7wkwxo4/fdJxHHs/dU/ToTlYWrrjNjOyygyg4Qe0rUuifz7iCaf8dL7
ZNEzaxV/sEFyPQhL/blRERj4+h/sD6IpWZniETxV7z1fSaAp/7PmUNTjhBGK/rwPTZRLO2NpsX7F
IzCXKY+bkgWHPsWCSpB20psO1dbq5MzxL4Ew1UAlK4huBgdR1IoHwSS4DebcA6vDa5kk7aTkXcJV
9rpG0k1Lz98JNBfJP8yTfUPPywg+37vQnUpzb0Z184oRC4fkarsRQGln4B0n5gKCrba3GTz2GDo6
NY7d6I6W2o64l+WD6y+teShLKkLChKr+HKnqfEKQFLHR97N1IfEMppbdS09co4dMRnf9BNTdr4YL
25HtWHd9I/J3GyQ1EclKPPFZrkkqvKPdCqfenYSh+7LPt+34Z8mn1yOHCrL5IOI7idQidmk63Vxp
WJBmKki3MRDUtHT/u1lX7XIvCv+EEIkgirl0MHwIYzttnrwxe5jGoGmbvByPu+sJBEfPXo1ECBOM
35wq11DUpJnlClrF9GNdLCsFKs36l3aprVrDhdbnXxs5oGRngJ3o1Dh7MHSMwBLNSPoWo7jx3zpG
9CtGHNCCMD5EPCcjwmwAr7KuSzwKpf1NlMNuSjNVzCnnInRDS+HVAu/zvnzTZVeqRzWgpHTrEgao
EJeCeDYkB92ePlpQaUX6P+NXeS6ATLAImDjP8kxFzx927aNvf3soKSu3lJ8pWAVV6ytIzIUYLPfS
vyR16dQmhjeXePxj4Rhn9VtarSJhrUF8EqFIszBviJtzeAW6rPJBZo/iCTvhSfdi8UgQ5x5dB14J
jRCncffrGt7umWEac/e44DazNZYO/uaRV0pf2hHu4Il1XBNrn00dqfIDPUgde9vvu4RxUy7TVlQI
lJqZRHKhg78pwcH/ndghkYkEwoucMoj/nM6Huj/Tp4cwQu1iYKtqK2Z6Z+Bn9UHNuoai83FhagLC
S+W1i7mjXzls15nDOobijxj4l7Ke3xiBmSul+cKpPezIe6VdklMZAY4JavJb3G5e4q2Bf5IRewqz
NYxQAOF91eiALrdEWqjlAkf4a7FMtYE/FnxZqhmf1vaeBJswCnyWDgfYaha4+Rf7K1AZMWXU7DVO
uPQCU7EqyQZiwlIJtqJo8lFO39z9nGGC3Q9Il+JkZbMfEN0JRsHApFtsNeCt8FYMwhlcY6BdysHJ
SJgNCyErYCtkT5L7Qk5l84MtS+L7UMQP2ZSWEaqcr2pt1KZMrz/Rrd6ZY9fCV8bDlwx5+FeI+p2m
VuT+2lcR4FoNvxHVHLAIoOorPWZAv8ZoS677Vdib9l9npM0XF8pcnohWccUuXBujOpVWuX6ak0w4
3iogLsO01yGc7b6ecWfjgCHiaOqTsdxWtp1Zw117wjG0oHZq+HhO+0B+RzKhnbRvto7pDEwMDlj9
dYUfPBlSNJfOaPkfgeFCByNTHn2yf2H7oaEXYa6rCvp+/EIJ//aCkNnPkF6OJY6Z4DRrggwtVSs+
xJwmZu9clBGZETuU0VAKkd7ACMBrNT8XehXaW+ek+CHH03nqYpvs5iqMYW9xG8+EjxNfMrysvzTz
trA5AM72suJQs2AiBnJMojqkuG/0WoTrnX02IoyFt8G8ZwdciFkoKj0lThYfgwxNCAXeds4fCWkx
JvGpMW8VH4vS3BKfdZ+gkGvKEPFS0fmK0KBQ4HHfIC9Q5leh1vsfFHT+wOsyVqdN38xe3/Sahr/m
uuhdtw0xPpggcLuoxDL3vF8QZwGdVdwhP6zZ8vQF2937vXnq0c37vpJ1koqag5Ha5RACNstNHUPw
fB9K6y0SvfgHAnXuhswc5L0kLMIhuI6PJydx6H0eLPqsyDZ62Qfpgdp1EEpOivwA16zeoRdhjalt
tA+2/eDXe4ncEdMDpZ198WD+zrlOAUtqQTZNEybdYoqUETSoQONte3Wm/g9N0UAPHMi82S/SdDlO
qJlZHaCdn5kJX8uw6JcOquXlvsgzvP1cLJux5a1aWbfesqum/bUy2EDYWisg0v5/0j3F/kylbYm/
GLltZ7JOGClkHSPjxvBX/Jnm5ojk4rVa1Lim9li2/mOaZOzY43RApBv3DAzCtaJk/5QDb+ysavB+
cdS/ygQli5+OqrgkdtFLxalpw4WsxWGIvjZxmhf2TldywEqUzhwP383j0eX45SLsZwKUw3bM23Pu
J6aeZofaCGowFUkvOdLDLqgJ8fQgcn0xUjlEhwd5rN3I0kX9lyPWetWemnlnX+mAfInPER1LNNjk
egd1b2C4RbzROe2XtaUZilPH4D7OvOLU/JLquQ1J55PxQC7ZJX549yZToiv2PXzvgpZ48j2Mw567
zhlUWasicF2WuU7L3fzCBy9BbzXvqfnSchsLKvRZPVkukqdIEjFvindcIN5qWRMDi4sIndwq2R8k
jW+32Y03as0mPRGA1b6uazatm5dT4j7y6Bsiyx2K+a3kOLxFUBN4mzUY40FI+y+XOxQYpvdF8g5b
lqhCjyS8EoQeKwOt5fbD//WzPoZk956W0zhm2Ea3sNNS5H95kLBuLo18OhoAW3wI/Y4Pbl7Djete
1eGUaqzi2aQmaGfWncfgx2lqiYG7f/fmrHtdINUDdC5nteAzjcPJt8CBDa+v6tKgLGtziYtlJHr9
E4E29F3/JCobWQQj0+wY/MmrE4XH1qvni00KHXgilh/QHMvE4kwE3ig692VVjbLo9FvqojUMUvWR
UMmVDahVpP1W+NOOG8KVNfcBRbByDfKdssXSYCoktJXU6jssqjDlfw088SbvOGqSupposPl65S/j
CLRTKz+Jj/Tu+yWX1yaQWo4BbshmdXfWxYDamifyupEVTMl0R/XAVMUBtVZDkG9nhhc6fcOEAkN3
/N7cWvuZKqD/Tbl9iLeg09/bNF18nMi9If/Kvkp1E1GHQddhdrkdl2jbfuVhPPek57CokoXctOOT
CvB8OPuv9Ryr1Xdof/y6b3va/S8CVcQf1QPzEwwYj2BAGE8WKEPotKQS49LEC46BriVHv6PfWjLd
3yA6rqgjVh61Qy0JJXHb2c0vfiNv6T772qaY1WYwCyiRvyg06gN+YOH/sZ4mkLWJS0LwuoPakxo1
zwR+f9kSDyE8EsMt+f0SbnhAWJqIsjFxwEKYnwzkDz0quy3ODuexFGyWqxRlwCdKSq491Sln0b5B
O6Z4yUIVytmCnqFHDHL/sSkCqLNzP6RO4BmSafKvVEvYjcDUATKYrfT/JmzEhj/s3FDHyUh+7kDs
CbtQnMfk+PueWeVQygHWAW7bm7i0W5y7E6/kxw9s1QndNm+TNlUSEbEz0VeFGIo0XBsVJWWOk6nZ
zN8wpgf6PAnKpNK9/040SWAjumvRe9R1DhbBodxs5SMDQtohYsJb7CBrxI+HTfvh0XL5Ul7spOH8
d8ZT8i3mrS/kdOWZ7voC9WN3eQWJM8EgZSdwt0B7d+pGLeCo0t4OXcHFFVwWC4XDY9QSWCS/l1ws
0JzNeUwLxXbOnvxpl58/QHNzPKYQC0NuDCAXDir/yu90vGlSn4NmTm4rHMkd14oh49h5qLA8FnEA
Jmi2hae0r5xoEG+Tfe5QEA1FEEmzfMzFRfLl93YD1s4dKLjgey5obh3oz06mgWFOlLE3OmN4Ed07
67/f5cNhP4NHESwrDAQREExZ0cujIi2ke0tDHEGWSLDPh/qGi7kMZlBgKpT7k6PVwa3U25aaY6SL
HNP3sMcK3X6uziPzemZjIPUaY06dlqCMwjhk8zcWcQuX7+d5urK17XYWeldiHnOjbLv8Ygg4BVpM
gFTtxjQyeegsudo5OwFIOnsIlwmWXF8e24OQhdKONURkWd9x/eQAhZDnp4h6tqRq/NNHrW9cAhY0
A1e2qUUnIlILKfo0G+ZGbNfWYThFR/o0bdEUVmDZ5BSpuYonrFDvIjtr2DKaKBuS2GdZt0MWZU2i
0v+beLv6+H2r5FkY6isED7rn3Wr/ZStqsFhQ9aYfs8NSttLj2JyhNxDtgNEXo5/xt/uhbGqEKTXG
KA3KokAMukRizibuMbcarCqMSrJcOULriDEyGWM2X0qPsjVUduA5oU9h8hYcQDa0afurbzGrtfD0
COS5J7a9u70fy9tqFc4+SsdedREcDLAwUmBPCv7eGsBCUp3/24n911Ss9NmHjtzhpE1jqoHjn0Wm
GIy3RqGHeVSQIRtB4ar7ZqCgiUz5I4cnZOPI4M+ilSat3tlRoS/Hb10sMqWCQ6DN3zU9GabV+ppn
o10jx41BzMTh6p2kH9xwWCXLDkML0PigpuYiuTH8NrNqqHTByKJ3PrNb0wO/ZLrzzTWP9KvNV4z6
LsjhZIQpuUjrwsOny0Oq/lQTQMqXt6NPoWhL9maa6lLJH+/NIPkR3/xRde/mpm4iWxN27324F/pg
po65RxSbiTsjMtLqsfUnvxtPxCaFryriSuDQiynoPtSbfIDkvICJ4oiJhJTK5ufxYX+ge9vPTMtO
+8Eu4dKXZmqsiXefYzHsCyDBQh8NIFC2d6inh7pJ6r/wXOcoguwNpHFWjuebSpdniSLTU5/PkddY
jQNfv4YplTMgzm4T/ZC7eFx6zZJWSy7JEjugTKSGFHPnm9u5+t18FfRJ5uPWnwV8mFi4O67CKXBh
iTZCWtovM4UAMiHhby1NCQ4RCHNuukboTXqfFCAiwWatvwl6YrsIB5a8YV/lqI9UE4auKDyDJ4w5
4p0Vk9Wfr3F92tSUmTi3wS8XMx8JG7RPQGnothWwOASWbB7gwFmG3llKjvrMGjVr6164GgxpPCv1
2nn1/Oc/moswKGOXoILPZVbMniQ7SQFJwvUU2I/TDTWKXSvH0OivBZ0Ia0eSkGrjpW14/CIOenNL
eHFNfRTK86KjW2AjyK5/CoLn97i4kLLM+7FIEKstzGebbXHHtUipMQiNDQeK+D8V0esQrfZJa9IW
IUFaNzKjxJ5VN/Bm84K6rXgmjreXnI8rkypxRllJPzOxCWHig7gsj2yexP9rgMaUZx6EHYpVKg1L
6fvKkl17XW/BHF/fk2fvw9SNs5wwLCJVqjdCjHvxDKFS1mDkZfAL0MLfFZ+H8KI8mBw0JfskCF5y
FpfuM2rpbqi7XXg8K2VWfLHT5llukoDh/j2s2NxJPkTKWdDjq1XciatzArLY6lZ2o31FY4DQEQx6
9fI+p7S0h5Y4o9UypoOYlsN4iUqshRsh7KFlwrPuWf0vZh8aj2YJWIK5HOoD7Odsn6TaSP+s3Vtr
rtAJ9o4Vye5TDkDInZAJPqN+Ab3RxjZ02pt1Cy/So1Hm0YuBjNNuzI+4dye/CO/sGAQmYei8yY8q
4hJ2xvTQ7aPS7k+D8DsGa1O8pcB+RoCWpSODIBe8ioodm0U1VXgWMI1OUsH6144sGQrq+UvesQS8
3jduK3RLbIQj4m44ZpdTSLZYrNWrkc7VOdXJbvuEhp4oxwY3mwk7XwMOyvI5dCFrDhomNiDhQ8DE
q+vwmXBzP0tO2H3R42wUNt1fjQF2Z04F2EcmYMzVOpr/Hs6aM6rddO7TCrnvVKghJ8rdllQ6dsxI
9eQgb6Ha6d/NF/VEWi+nFJRKrDcrITCumUf4x35cYFhgpXUi7TXYe2YbsChM8PN+/StiTP7/RSkj
LaETndCTwlUbF8SvHnXF+LunIHnTxcMUoF00uu5eBMTz7RYXUj47axpZ/M6XfvBoFqmCe2UXg1fe
o+MWtwbfohmitNhXLR7GA2GnjP22QteRDNOtxquT/x/tSyT4CJizOZ2t2tcgkTVU20hIOTxLMKEc
4pqXqFGLXcGXXa1+MB+El/XuiujSU2M8/C7EOh/ZLp8qStcDGTAR6wfIhJ+O3RCxG99cyVq1V1mP
bbnVSyDq65M7OAX0TUgEhISTPFXgouTg1I3RIqI+kAIM06ObNyN111vkQ0D+zfmtX1toXyd/+UDq
EN1Yxu4IUuZR+ud/kugBd+4/xOldQyrD59rB6h7/vEwvDwB31q7AQKZCytJG0pSWpVMj8LfYyK+o
Kjf1Lg1XNMn3TZMmv0bnDhUpi7mMnnhchs3WptkuUwxCqgUC6dOrMzMBDucUeTLh//4MEArDRG71
uIbCu7D/x3k4KivfczsLthJvF+bUMD+bT1t07Ymd2n2NFbVCClCWKPy/P9TYbMHYIc8XAMctybMl
XrSgI98unSR9NB8EoL3IQ5GSyUCqybpMS+/+dtO+bNzOj3dxyg7pmBU37s9W0WzirUvaH6bQ7V/s
16P5irKoRasxFXKQviY0jCEnsxTGDLKcmY+xPHv8NQ5ccLoVVp1/ymPziRx0pyRIMK/C8XntdffB
pOjWPhruJseMngLD/SwCOhFffTY2jaUVcgMZjs4h1NDr1IcrwtEHqIWcPZx+WrO5+8CrQQID/0bC
hcFsBdNTR4DLcGJQRdtIZ3mTp5DJVJf38TVOyjpRYZFXU6yOZhfofoLsHFSmwSTdlSn2oeuF9jtd
AL6PO2JkJeApI2RUgMsw+Gl7vB9abhpo8OtmkwOYy+M/wHqzyQgCRFg8SED7wHNflIcLo0YNknLH
M2Y/SN5gk1x9eZoqnTR1AgonK2sOxzv80sntz/GLF5MEYHnpHvuVfHzozvAtTuGwCznogifFJ0tZ
tZ5hNtAl05qZwTJEgil9s0VSrEVRJJpHgphuhf1+O2iv/1iOFmgsxGFKd2XXvCkQZtUJX1bbZ7Rq
9PoSc7GNrxpX4IIWwqkmpggypJSrD+Qcns35DPc4+SlWKxc4sgHhexQWja8TsUYMbuVqw49Yu/fj
m2/vz9mYy9W0XqUlwAGLdLppZCxvmE0EiNUGdo6hgZTrm5WW5fFbcda4L2tD0kAh+0rp5ENkCzNX
BV4chASAQj4AQlknIeLaeYNLwpQiRE+uVXgRH7UASYQwToBcqINN8TwX/0LJbroSFTgLPjN6Pi+F
bvQo7ZE7uNibwhivcMMI8DwoF4kff/w1Qoeir9CTjQofCtilq90jIKQRFHjGYzLo/qx0HD4msRyD
xHLYCBShDIW5djlxgB7XAiu0AGqDZvJfYerfUvT4IhYHU8/SM8pgai7Cxdd2CYV6obTOxNpQBYHE
4WY0ayAVztX5VWXyqgArzrTuxyWwRXn1PcwwCNOEhQoiW3t3kAjB59xmV8WXVCoTYXMHxY3YOpv3
bs/+WA4xUN2GB2NdV5RFGidMnVrmbHhdePX43OocM3c8kAZnBear8WFbhhy2gd/XVOD2T4aaXWgt
qHIyZXr78+NNiPs+iqnf+WikheQcj1HAkcgRjyvKb0c+52G3PP4UCdjPFj3jfu+TEM9rTAe4jatz
Mf9zyfYx+4IOIaUT1tmd2Sryf7ODcKmObR82F1piiRZrZihb+7FJ0JrEzupyffANwNENC9GSbMMi
rq70rZHMw2VEOX1WjL1aHRumi0H4ObRiT4N52Z2DnmWZB4js17Lzye8mZnPCX6X1abq69YBihTt2
k/sOQ7qIqIkR2toxmf23RmZP2aDoyVZh9P7epOIJUIxXJwm1srZi4Z7XD57n6xQnTNu2A01k+mzq
hjvuKfg5xkTbDgHuLKJyPNIIOeR9iWGYwJgIqKEBIv2EjqttOKwixjhYk+mTEIpesmVcbnKfIU6V
rCZVnHAEFMBuzB2FbB3wUoZPQTTSSoQVGZP6YcA2N7uePehrxv4ukrlqAYvreIPAMOkKUouKKUbT
GSUKgINYSDMiE9M+Vb7j5BQ4Aur5mhDs/GU0Lio2QvNVEQ6zWXzPD7Iv3UJ43ZjVNxElCGOvjgGT
HhUBKdfLrTuflgWa+rG3hAlDGhXKivN4GpInJlh0HZ/dG01JdWhba/RkZ/UIPbJUdhLN/+vPn1MH
RmQ14/yK4gI/OUs1Hbj+usVw3XbeCZ8OJ+gPBmfsHUa7c4VA2ZLjhtMnRDP6iGn9Nyjhky7mfJec
0BT1hQuSRCUNJAWQLG7V9J8NRvXw5y7VJfIJyI629cKpWXHVbTsRq3FZcPMJKZ6Ub/1VaiDle+V2
RcLX33llXOl2/iqwA0803WOYeEPUMmQuFStI8cPFoHa5NS8HINEE5HCUS/XtWFBuMNtTyqJiqIEm
yDlooT3BhCtDCNUlXJUrxTI2NJwrw+R6Xveo5r0NmSGk4u7a1OrQVeVcSQxk+kvBbSO7pwlXiPgl
vDMBbp23wFDGpNpztfk/bk21YpGNCzN8MjZMyESsigegzsrRwFNhk/VkVVAymE4TW1lv/drBnULn
L96wJMGMFWcjcFMCaAtlw5iihYpMxtf6MA8UeBjBl87PNP++d96liuPOML7n1ighOHwRRJzgBwGs
szE3D24zTSBRRJWnj8tiiq9lnwuZVlboagVRYaxMVpHLbjcLlyWT0eFHrQ7IWLMtukAt2w6gASBt
lsLd+WI87kEerH5BTUpyXQOml0ygxWESdaHj11SG/RvHvDtZrqv9U6tduZdWImsQqKH+yd6JIflq
ePtQMmG4dqR5AAVGhu2dN33XrMWzwbuWdDUcniJcxYCFBktelxamIXO9YX5Z4LlA1Dn/TqWl0GPB
sZAVV19F6S7lsUAwxTQgsL7yxZ3k7Fuxt5fv2cPIve8OBZBrAx5hkP19xmhRX+r04SchKrEZ1wwi
fjB9xhH5AdDuwfRNvEd13GaSsxTPDVM1AmvRq+4xkI+fT/RqKouNW3rvTrPfuN8fwamGgC73KVPt
X2sIIMwckvK5OKn+afwVnSM5HszU0aeW1GhBgFQAfw83Op192/5kyBrzsnC4CVr8WA9h/O5UpfU+
Uk2rZbgfngwMuwgoVxLpCOPf7m2N+7MTygSw3Zt/NLrgJ65StGxOarv9JeXo7QKlveFMifRpWh8+
/SaEmJsF6Aq+u6y9E27m6iEOW6qPy36/Jb6TiwvW8wFXH5NTmfUet6Vkomv9EZUdspfAKMffdRr6
UabdkQC1fycJ8ZP1A5GhlbmYxtPZIkXRbnBPETD60KUKuhaoEwqxM7PFvCA1V7zJGlplesdt9l+f
nBUikNIPnZl2RIgXFdHDrEvBJ0pHnMFvSdtnvAKkWbBTCp9eitvyfeIqLZLsBZ4MU+1zQZeMBYYo
0OPU9LB3ztvHbaXljw0/xnoW/0WHRUMq8EIQCvRBsuSgftejwTFmRAryOAskJfXk75fz35CRpBP2
lTXfHLsolG0v9aZbkG8YcfrAaqIM75C/SSDV6orLLfrnuTsYPislNyussq495OpqicAPJ3Ljxzqb
WX/Unkdj0i1zZxyJ1udHr85AmAmYsSD+1Aq1kWGDptyDTE5MCKBNseeWEd1lPQkJmjDhSOJuuISo
6KX/f14vcgdlXgkayJfgQSCS7FGWNn6eAhoX8AS2s4X+F2opxumEdZRl7xkN8UYP2payDct69s05
NcrcuCU/l+yarRQ+laNUHQZE/ljFW8YjZ+dhU/ZJ+pof/5SI7Ub3VZj36wZ2oIzoc7BYNc4wBO07
WVIG8iNz+tA1tqk+4HYb6xiZGG6BlMy6hkUX0/1yYiawoa+spbSk34i00PvMzuHUTm1rmyeQhMeS
c4ZHVM/Nzb5VnMHNjjp9faIPvcuyiMWDGJ5DkiNOJtpM29hu5+Pks3xn4Z6ZjZBGVj3koynkdiY3
meVPHwxtu3NDkkk0h/EBDoDdM7Xk062djr2HxNNqXpgnBg/H3aZ3uKVtBrj8h+2n12GKR+Rh/agg
iSXyH12SfKKu5oFbjXkXQl9cnBAiTYASryHnBUroTXN6DLPYmRZ5YbYkuRFKMogqrmvL4q1c0IVn
ZalNJvwMvmzTiIkn8wU7wq9Er0M/39RlE3tOO9ZN05L+ugUIO9p7caDgjDvGpz0wt+RVjXabv923
y8Dfj+sXaq36Tieu+XPb9w81Hv6wy5LYPxVteXdoAvnKK026rKNt/yuJ89eQ8/6Pc5NzdYXkqxsE
P2+rVUhC+AcLTTIUtttglfztp5XDTUr25bXzvqxe2YTs1ZgEe6Uo5gnQd2XCBAt9CWCAV2Afcg7w
bfwG1toPwq/Ww5K9NS2lbidlCElJasHMrVjx4zM9UThaWym1T5JGzZTUFFFSOnqdPwHiL4WNUIEa
fkXGulaTB+xN6M02Usb6Z4tAR7IYiyborZcfiVtR3/Ft+qy4bjqKkGdWN1VX/qleENLei9FdQceI
jf59524Dh1ifWL6mcLH1lslRRPdG9ciDJlk99cGYHR1eVHkiAH2ihP5Xp5B0ipwyw7wLyQc6uc2z
3f/YAJ2kLoBXsXrq8i81dook+NK6ftVU+SnJMZEon6hkOXpNp75K0qyNKTq8VeIgbYxZTRBPd9ub
So5f3OMhH7SJ3YzSObXW6vf/8oGYynz+SKNK2csyA43rNBmwZO07/xYN+YOhG4c5R/TdWI/Uczq4
2jKA1A+1L0HJrjUwXzeL9F5nTLKNNXxpbOgwPbTQoVNFTV91bIjXIqjGNVKtW6go15YsCKhOd365
IBVs1ttE0CzE4nzv+eVAGXgdVs4sO3GRb3MNn2fep8Mf8V/y5bCHkXYPeSwEOzX5Sn5BBHm+Ac5y
y/TZjXDauJUkJLvKjvCNlbnqyqUc+WimcFjSoOxIduu9W/JFFCnQ6A7JNcy+wCvgWXuDk52A2wwa
nxXVhsgaIbdCIjFkjYocSPps8oVRpI0+nrTz83IQeyaXc2gmkVGlfuHO0QyhoVUux3fDK/wWJQYD
HhxPuA2hU3CgeZZ6vWgQW3XdBChJua2/+npiCPVnau3+nsWCR/aAA2vSsQxyMfUSnjBl7VOLJbcQ
+wQ9jBivucJB/pTriq4zY4+QJNGXqum2ni2xV2nQ1u7Hx2WM/ZZfdisRk7wzrve96Eb+/afsluBt
uD6tIClLZw23idvzU1s3hDMw5XY1gNGNFBjoBn0BkJ1h9BYzhKpPl6QKEQV/mudcHxrTbmCgJHg9
Fo/d3Jp+ZGxsi2TW4cCwXp7ZJr1O/q4u/vqzaJTmGbmxRZJzCeNgVYhTEvWC2jvRjzENwsaRGg2r
zuLbCK7kYdpEXv9/keeNZtmP00jfwxF3N58xdJb05N8/bnUNWNTFs5EKFf1pTR3v/5jP6GyP4i5T
pLbiPelKTsnEBG82iSqCi7oIgAK0bG5JGAZBeOPFbrFdthyJyNexHkHHTGkTor15sQOKVa1q4ShW
HqVjeBUs06wYdoJlDZxRXkqTDCLOYbhYYe+hHIkP5Q1TxAlcnK/hnzhLg8alkUr+NFMaSNNgtFOY
2tcr+5Ab38tiUA1Cm0PXhb+3ZG433QzXlbJuP/kAqsZdAK/3UEwJ3saWP6RRfWPyHc6bEt9M0rMF
5JFMd6pe0QP68pkx8SPieVc42XbMeZ7DiN76k6E5Gi12bJKDmKKb6QEZh1+xgH94OiCs0pXdc53+
0w1W5O+S1++DsOPnupR5vzkOs5ilPrAMF4kmtOBZPolS1lZhtW7jOFkrLwZToOSDsTgV2csytRRA
N5wDhWa2bOJ9yCXM3A2vw9JPWojyVge0tymAXp/A2hkeiqD2mzFTfjIY1CS93PxfLOUP6ZA3GgII
iuL9uOdUUiOM0Gy2tGgCf1vAC1lFwT23CWqr29iE9CuyXSHUJaKs0+6j5DpodTaLM8tgHd6yuiPi
rw6gXqXKSU0xTq4kGpHZ1A0pxl2mpz8zAq5yxKJqb9wrKYZcSQvcI/sgGucsXcIKuOGvPtAQzPVB
CVojGKiXWKXQPRPtRVsGiruU3pd21f+r5H4U8IekSQkGtRXnE+G2dTWwsllJgl9d6crUYSoltbzy
2fE5xeeLey2ZLUMp3WXDuiIoq97DPIQ+NyxBVyN9VKBkBSSLviLBKKfeQ3m8E6XJSSB37TNCIIsu
uid4X8ZfFyFIqb91MVdW4i0GBjbCw/B4tCn7TFbMVV2lqzQ22fltbkV59uOuqTRFORX+FUV2ZwRU
7u4N4rHIX+eFwkllk/SNQWf7nFFF774J+fpprKa3mc8m5ro1KkE8BcJ4Gk0VRor+7dmKXqwvJiHt
m/IS9WkQmTqwTkzcmN9cDn9lqMKfCSz7LzbCxQHMco8N2l2F4QqvZ3y8nFym+pxH9kXle3dN4WXS
jOxNbNmWfQV498BihQZ8t7XZJKE20JpMAIv0uEVKpGqZmCtF7S24Aris5IotW4BS3Uz+k+Bz7tgu
TGn24L0TRf5+mcyAMgqQXxbuid83zdhPFph19cu1mIIVZyu3C2gS4T3842hE9ULQBUnN+cNINDRV
vUeQQHp2U9+XWNoQtizS5l3s268/5lpRtD4vFlD+A0gi1yGJDZQvH06zdyjpdlfs8Ub73Vy8aHI4
zj7gO7CHI+KdJ66ydl7vJPSDGUneMDTCu4XIK9qRg6U9H+wss5hi2DgxKqUe0QAtu7SvWmSTweGP
Tk1y2ol4PyMCvlOZ6dKx/uPLr/duCpTMPozo039FKYlC1Z0kxTgce+U/r8MfOUDEPrLICu8ttxqV
qMQ6tSVgv2EWTWoTQ9czilcXloVKs2cXrnOBR7qdpVTc44JmVpwovyePmpUp5LPuIaumgpaRwk3e
iS4lZ7HZKdNofR+VzdWCJt1xHLY9ixKTORcOHxFD4s6JvggIuu4Ld26rU8985xFIwJfNCnlPTGew
obieP1JC/yLQqp0gXv0E7qPaF7knXFnJZ9J1kmjkP1BBFXpsvXz3eT6uucAT/6NdQUXBYaHJVbDu
L9sFvF01gx/BLYHptghUQpD/O4o9/EpKizQp3Q3d1JIbe2PN3TfyWQ+y0iql5BpCVt6pNJrI6Akh
b1MHGjdmSYxysegQIBWhO2okpxPghT8dcZoB61n0Q8mWqV38Cl1Pm1JRc72q6RPLT04BXQkGXBCd
wImmBGvrfL2CKhFXfnS6o0J5elIQVpDhRCRIfWtzzdRIuIkqmLBdtabaCkek4qqjTQG/d/yZ4dp7
8ipriC9V6At2/g6ryMRJ8G2WnLHMr3EOz6ZsdDqd1Fto/KOsVzbd8ZfEituBf8PzPwC0ak9TAl7c
M/8cWiOr+Sv9FnWk/5fPJ1hG68VJ2UjUY6qyhK/aPqs3QkQJ5yEXWfTTMPbSZ4JZWhkcU1JdL6uV
lTFk6y1R9vBc91gD/4Es8Lp8r1uAfxSa+R2KxSHpDMQ1DfOyLOze/wr4kwajmvx7kBDCMfYRF+eU
vUwe4Hrzdr8U51CAz6+jf/s3eWP8a3ggkB49r8lFyJaf+TLkW9FBNncsnfDZStW9qDd8vF1dMr1R
pW6CkoqBtEgvUM1BYkYz/+BkcfGukzBP5DU0Hdot1B2/hCEyh+lZGWd/S+ZZrHNau6PjhMMq0LUD
JfFAVBX6W/ITTABqQDqeuuN64jSYaIab7nRO37U4d9kBEILXAK/++qJWuzeY41DkJ1u+uwTRwrGl
h/OV/LxDn7VhxNAvKI9FslUOOu8ePZpICwfZjh+IMFXBRva1M8UIKOyiq+dKOn7YusjNxQnqvonT
FObIhnlA61K0BKYBHt1NL0zubhzld4B+6eDpJOQx+sY3XEdwxAsilcJOWirzPwPUTixkw6x+9C9Q
8aIarb0CQZqCqeF2U3Po9Mr+PKv75BU0Wc2WAl5HSJvUzxJa7FKB+T+N0EefxA9QwLe5R7nEgX/V
cDxCSMmVGlhWOn74bDmVofPM/lPu7ZozhZ9Y2HIqttA5FaQ3VtjmjRkL2nALkbs9HXL5ZMbZPBaA
5RoEirLltMuGFQKdclFZQDRTg3XojzDKs3dv4QsUGNzPQ7sCbwb89bHX4A1AR1DJsNpOXRpIkfIn
ndV7m+tIwS1eASVtDTL8oe3AGDvdX52qdHTCBN/kELyGN6F6hccOhR4DYAgY6w2FbFzJX4KQozzS
TbobkBuIqFlBXBHm9yNIMD4Hr9d3XDoNgHof9xeC1WZIuIPlWw8gPVZxXvFdecVS6dN93NJ2bcPd
vsX6YWbAKq3dRlwVypo1uunNhRi1FUCAaxwYNTtCkY5su92xxaa+7UXnyNsP7Cwo1rsoEKIQQM4M
nLUZs1Jh1vepyqImwsbp0OB5Ed5z2gmNvz5SJQ8N+qoh1tp2+wxMx+jpknz5a3ma5tZlBPUKS6JU
fNarhNoWiSbHOHkIzon07PZrUoRK72QKeDjfECd7VXEcP2+ycm+8+rUWa/MGVvlF0vHiwiGRURmi
ger3GhF++DWJgxN2aANc89dno4CDPNxQUF27lGkvRkHJhhhIrUu2osVEWhBDwgv9kH7LRABsC79P
4HNWn7FKDEd2+yNUtNmms/F48lY/C4l85ipW5c7XBPP+aj6cj3N18tMmum0s/AIsSMUc6p6oWAHT
6abxAvENrTo971NKT2l+V/hJseIVKFKNbBb3Bs+EcwRqwE05LCWkgClY9890bFkeHppvt7R0vgML
ezC2EmLz2gse74+1vdEckhKN7z/WcktAhf8R7r24aUo5WWkVBBmZDFBZ3lGkQs3i1wu0Ohr5uVn9
6N+ehraxAMZLHZHyq/nDvJd1lMMJQWt2HhIv9GtN5clRxstF5Ls57IgMWw8JQHJpHLoWc4+ENL8q
FqySy2jwK3p5jG5epsz9y2H5v0KdrXWcfDpq9OrrF8PTjHsKuvkpDdgh9DuoHveUTcX9dMrsyU2J
AKuwdjPzJjRQri8somahWK63iGcMl/VnNvEVrNYz+9l3p8BwkCM5cvxx64Mc0LJHmMxXChscip9U
jHFWa88Sg/G7dm44t7R07tYbr07svQde3tfy5wPBYiD55SXpvxMCcvdnZh4uIcuy7nCVXZNRkqml
0jHHlwCd9ej1VCNa9HTqxXG9/FIjwYulaubZdGuggO9gxnr4fQC+AZsyiB2T3sYOyBj2YqrFMwC4
O0+JLe5kDJ5zPGQnvuocOsNX6r0kwrcyz1+NOycjRc+Uk+L8LkJdeEviJQ+4Z4ifOXNGvb1EQQLQ
5/m0/GMUHeITtPMxprgGitfSs3U9rNmcsein/8KHS3ZhvUgW+2tSbX2EBA+YRgw5fktj62uoNngf
tAgTaBM/T9qiQgV7SDSxLRiIFEoGp97QK12cvBi35JcdYZvbfjosEag/CgyEFDE46kdiSpTdzDZa
yPKnI6DM7v9L0ysO1/Uv4ejumLxrA0e3V8BycXxG9+XT0S4EaedeLtBXDZYL9OJoNXTMgauGLYe+
WadZ7hYTw+843dTukHavrrqTyNKZP7aW3Dta9Y3U3bRiO7dF2HHHsgzXnp0OrX+2BT1oEkxrm6Yg
2qwf0kErwSlu4k3ZAq3cU+RHQorEDP+pdgJ5BS6EI4505w8nCLjLCJZNkSHmK4Rm5SyK/ftI94Vu
viIU9MNOS9YkaXZMCn9IxF93uSr9Sfdcu3//7tB95L2q25ScVj6vTAcFkjh5C2uhGBEGlE34dfbY
t8IJDVM9IQcCjus24Vj7a3U/45dk7wT05pNQwQhNglnn41vwyaGgLu5LxFlJwUFM9cOmcm+UWkXV
uey+3Ojp72imWkwd2jvoKlF6ens3WRt6J0mRxSURKQphF6Kczg7i/sz0/DOCC4RHIcrt0wDcNpSg
+RUxPehE+jk6E1Pbyp3QY5F56V3q5LZG/yjyUFCMBYHZqvUfkEgjNZIhaAkFJNJc0MPg60a/feK2
YLid+LP7FsGTaUqonmzmIqqMJ1105FpNCcZO3y+7gYmUMQdtv3bsKthWHS1XycYJHT8cGqrfNb+s
3/OKBdRRUo32Gy5+exp1wGOeCc49Am4sHx+HOpvZzR5FRA6m9HXIkGGDQojztjrs43NS+yfmKyau
BvYWKFqjHT2reqXJYj5i2ryybUA7CY/MMm0uWTR36WVHcZww0r5LAJ9liTeiUVUhqbSIrvvODlZg
VKreGPRgDeefaIzEwr+szHMKz5CIL6bo4IHIRXDX2RhBT7JXKMGrafuyghnAJ5OeKKiU8pSE6Dgh
xXRgP5fxMJXNXdNwYGXQm4ydsXkSkmwlysD4u+CArS+O+WidEqgvQh+ikPBgfGfLCANwOTqmBetB
anAw3vDRLEw3XBZW50wVNRBRiOo9IVn5GSQ2PbManac6CoIFovNAEsEYqdgmiq38qx+4BK8ZfITV
GP89kJKAAXNElJjrFi6Ien0+/rTbCF/yImjO0QlOxjJR5u/LgvL2eYKK+t6Pzc5k1QYW5EsimbYx
pA28nAghXHfA5izEVgLKBa24PUnwxJLbTISg2ZpRlft1BF4/aNx8JD0TBEun33CXkbxGGUQukjsp
RWnZnebPLmyueUdsYO6ll3RApnV2rmKs0FBa2X20JOsdnnTahQDa/i847/6jTmf+glG+nIddxgZl
a8m/M+qEKho9draHXuaXCxFlffbn/5l6A9ycqpF9clXkCoGEAq4upPTKqpV6PpUeHoyjZh74UoQc
M0MZv91i/MRFthuR/itE1dMsRkekxNH80bb8tESbniv9SbJMd2kDANaPGcV8fOxBUZnrmD+iQik6
PhEJDSd/ORIale65g/XW4oFx/pCtkHUQFsNgAyd6ENUIabj5vgOy7yhSq0Nawu5PP983xNolfoBK
2hHPGZ2Sp4c7iXyN1RPPrW1ksy/0jGEu2FistOjJxBqh1IbTIgSp/hJwXo4JjZQ0V7asMlGC156C
rV0pbEoVvSQ+v4ztDhEC+gxJurpq33l81iF1UP+soO+HfIArr4ivQ/gnt3nYZBDl8Yn6MYubANyL
T1lmEjTwUiQZaN5hnr2yiDQclEw0Q65JvGGdWI13QT2Lo+7+irvzkz9MR57mK3GDC+8Rdhz22aLm
SatfGBqfTAApWQQc5or2Iuep+neAv8fiWpR6cWJos8OS/5A73qrwpaiJYHReY/fZb5thig4L11bt
AHcyeD4DuQGagkx36fxdLYzDAtV0WDiK01K8se0oPhebXCyLrfXGVkmLa4eOxYywpELm+/9s7BFt
Wjb8EvfnpLzooN3pcHjFPSI7EvThmX7VYVTES61gSy6TzEW+c4un7STncGgul95xZWfw9w/ByreZ
RneemNxr+DaL53pjy+GUf0ECAPOCL6LuM5G5T+uJXLNrQFyDnFtIv830oJzoZT08bKEOIMTBc/w+
Yhueodg6a47Noy0TunFvS19Z+rm+VdNiXLSELlPXu85AqkSDBgZ+zrgy4UksEm5RDImq8mOSb0o+
mUpHUg7nKjGQDSJkvFZIQMBetvph0Ix1I71NLDPeWlyTNVyMYgWXKFNqQ5NUPBar6rz6T/7O0OPs
HbXYneP+Hf3Gv6LiIg957Ox4sTMPMdeuOOyqIfppBw5bwzpdrrCImQgchK3HV+ALue1blIYf/jpi
ma1O53zsanfpJc1culHOXjSyUwbnIOfcBFI4U1CHUVvJPfqoPDKOGOAj7JoLL4iO9RT/t7W1okwg
KvnOYF4p5rZVH+V3ki4akMKl3q/E1uoF++aK0wZWLwyATpjjt8FmbHfvIckQ2q7VtEkD/R2QwypV
RxkB6TTVkSdYy915wN6l65fuhoDHWklOyrQRYSaAFFF6pRD++o6mXoSDPHpj48TuPxzuFBFPPfaF
aHO7plcv7Mzv4MPAgdQAvyxMyPJsjclrbZioyh4bnd1B8T580SQv7P56w+IjMCHwUrLleuA0q/Pk
a/67FiCJ9oNfxrSePmOU+/dVNYf8AUBWKiuWQKZPe8WWkVkV5cIhbabfE8dWz9oCRcj7LeOxwWSb
ki8YxRLbdCXiLO53RbqVBLkZxflbsRm4StL3arQtEq4O0d+B4n/phmK3e1eiLY/nxmtCPgadyWB4
AYNEBZOR+JJvIKcF7ugNYK6FH6vLQKzxqtlfd/g3iml3zGyh44iO2piZJtQ/yDrYXxv0kkoJJ8yZ
7DxX5CAsAqdghxz+hfmXHU0R/SXkZwLlIKplTKATrPAQuwv8BdM/78hUQLc0SN5ti+U7o/oSbDLs
uQsCBCt6WmU4sf+zx/iu6XO0TlOoCeN8WwCd9EQEF8iWTJtz4VxTZCfVVcD0cCEEQYqLmCbcB5jk
NByUzQth63EsRFHlVDZ6MfyJPxf/pCcNV4zfRoD8jS8tQBeR6EQxXazYodTA/+IcatJyDiwLqnyJ
bQq6fZfc2Lt61OqtItkQB+IYfW2g9hqDMqELnlW4yFufzjES45H4Y0HMytYAxV5rzsJ4rEkFHumr
eKCM7F1YdvL2Im01CzhJd6Ezlf+JZskj51VGjidetWATJ0nQtuKrUtDqjX1rCioeGiopgWKPutkC
qBnMMeRkq08SqTR6xreFxjG+qyOFLOKIyZnB019V6sTSvoxHSuH7KQlPqT7ikxOr0FYefuz/Qw0O
1vQyYF8l5ZWLcnVaQMK63L4TTxhf1i0XcDHh+6/houFLRHPxeLeM3Puc+fTKwyDcS8QV8E9EnJKb
t+6a/V8XwAeHTUIRpIPpcSvJ1Sfr9cp+FvEBpdf40vtAbbxcs55N1aG+otworcyuN2EISONfw3kI
1/rdSnksGyA/aLpCsANGxNZCJ2bqn059PeavktCrUAvD7dtWGrni4822ulRVZbFCjSMBhrmm6rMH
RQPpfNjLSi3uOdk73pbz0xV7KBBDABhB323iUBUAFZ4ToYlyNpOgncQXKrBnxvWEAVL8Y7N7+Vqb
qC5kDMuUxOpFW/zT0XrxAbxnK0OoxTMFX7CxukjwHqsJzqq9Wk3X2aBbWwPEvrUiqPfYrl2lNEzM
siUV+bTz76WFcPCyWx3qxXJbq7AHD7bV7KHIt1//8TUZ3p3efj0+X646ZAHe6eNdBM6QchuHO7ui
dNJrNn9vIEnWf9dQLi4HdtEp2NygOR5xp00wKRZs0g3KUSWLnuHKDvrMOzYiM9+AiGv2g6xznn6K
/4oVpyUS3rBCPJQZiw+vXC4BhdJ+B7AVVaJMv1B8ssZV1tAHCc8I+lk6mtP/bWkCZnA9aGDY5ra8
wbWka6xkVUjx4lxXimAPYVGOxamxY/0a7O5M4DrJbwCqMZaY4ymA1iYgGWsibuzmTf/QZSIgdKgr
HlrhwBHDIfxgVjjvDlUSMcodkVMTY9XVsic0p63Eo1EAWq5kj8Os3Gbu4v4M9HE3dIR158bdjXqO
3TGrhRqGF2PVYaq7ngDOmOg07ZGaycxCH/YVu+heIKt3WDb5+4aech/v9ZPsJ7AKD2X33CHeyjby
QHxBuSRiv7INt8FYy3uU1w75JD5tpknGpr9mpqB9zlAJwPsO9NNwWw/Ebvnj1kA0IeliA/PuCRKd
RkSZgPPW8EsEC4RfZcD1qAWABw44YZajtZiq2XuRnYBVNcBp/PiK+g99qf8d1rIddJbO6zl6T2dz
ew1e+TvUw1AcDFsEFMAPPAdUEol4l1abQJLO3gKfS5AN7ef6z+ual5svrSmBvJZxNQAAQAIE0UPY
PrH/VqK0Fc2PrrIuuVQ2EzTWACLBdvRh3Sk75BK9nYryG/dKzjAp3BjgTQWJMirjiqFneaLHqQXP
PZnF7ajalyBKrKsuiPT4cXEDqikgoLBqZb33u1Nd1ByO6/zttMDJWcbbkSW16DmhljIEX3fo5ufA
7UFAecCB4XSFi8d+gRdOknsFVkDRekW6DPUItrnOwwPyDgWoVzYISEs4abIED/vfKffCzwr2HSFC
YP2RPZMlVKk2USFWijnP3LTlUcCS1HJFNIYX9V4Z+cwEofdmgnKwjiNZ0gNmLjDu0gPzo+9TfCx/
VgpGr58oRKlnoNSoDX8tqU4otb4CPwQwBRW2AhQWTjeVCMfEuuTLLN5PYBau8ZWiR6eSmetARu4S
OcItUiyXkKaz9Z3abA8cv+ZwjH67lrPgwf9F/0ns+7+DV6OuQt0WSCN2fN4m44lzeIoM/Z72ILXl
boqbwJldXg8tORRmcxKFZxILZQxTEdFgqHUoj6eX3+rCOIrC/HaxSg4LlGj7qJedjRvbrDpWopGs
FxAtwrvyuFDT9r6KmEZL4RIooeG7jgJkSid8nxMUYIDv7eRcHVeVjai5YJip3fUfn3vsCnamhyPa
7WB86tjGPk21qEya5je+z4Dx3fPc4X+/Yfliw44HwgIEL69i5gPYEDmRiNu85JTRqm0xJ+ihBtUj
Tyhka9SHf9HR1Nm35isu20HFoWYBAB6nHC10eUSZNVoMGMGy2uNOC2llnzsTKnZlgJmBR7tb7Ypi
p+RtvmZ4b/p1q7plukIkUlkwE+J22JsjGZpetjBJDm3Cw86nDlboPmxCD3gCp2aJl6whCUkX40NL
6MlwEIAe2nuwBZvQFVc7dG2DqduwVINnDuWtOBZ1T0Gsh6ht7wcaEuUPppfsdNw0h864lIesZ8VW
x7UQ5tOB5TU7bqGU+ZpsNc6An5gVxDCdwoGa+W3fxkw8vd/WDL61Ex0N3nKvJCCrCADohawYiFfG
ytZO+pR5byuivf1w+Ye2i7e6UOE2V/xJzjVxHWJhHHaJNjMu9FSXzTpMVSvvL0vRNa5AUF8wNO68
sexWV/QEjJg7bBgf/1NXRNKM4mRYr48KAIB0RxfSGSr/xO0hYcWuWZcufJV9mALyjqZSeiTKY9Q4
Eq584WP1SJG3lOiOsfVSdfgr16tQacgCauTIKANyzk5V1mPUv2wMYd4ETvXpXqNopm7ORwqOfRxg
KqrwjJLhmjo66g3wq0iRuqMauZ25EaAyBJGnZ5jTcBJPw4qducGNuXzCkKHDVfKxWZ9wnO/dihNE
6ABrBgkk4A18vRFyeC4qKwhMtD0A9wsYxPwq9dspwDqY5dqyOlhSA4fpQdyqr4uzvJzPK7y7uUUz
i9uTyoq1eMXOaH0eATwg88lFpXjOJSaw1P+aJ8gQXUbiPcgx5GDzPzYI/NRG9oLBXEgxYvNPJcOl
P0VeEGJ1JAZoceD+dEQr6ltCSBFOdJWpKaZ7dLVMamhcuN2pqF6gc3rNmjnJetXoX7QU/93DC3j8
PsAjh9MJVBwHFiayBoWZ4rE99gVN5C82vjhiVQlXs6ZqSKR4l9I1NWT3dVFeBsD8PRO5q7hxqkwA
oGoVDh4FsfvcLyiTauCEEQwUfQs/27Y/oT7TL/5DQo95IPskh8IGpIgnwgHI0VJDHQKAI0Mai2cK
doDSuWIuPuDb07AhAOC/Zi/xeqeW3eCX4I59ikzQbmQzldBmAgU40V5sBAVHZCISFbTlZ1VIA7ED
pb7S6/W/pu+vrAMhvUQ/kcK7Yyta44uoSNZ5GUHeIEuAqc5g4+YSYX/XJtxscw0+7HRwQPaS4m7/
i24sRky6fFvVn/CZaBGPC6s90hy/nm0xcSklRLYC3wDOO7fnFYeTex7QP7xteInDoNYirawTGzaM
L+/xRkXqGhfenESi4dc3+aL+GEWTlpU2tmIGMjWt59E3Sqknb/yPIlxEGOHNIgoH8HdjAXWFGJyh
mCwj4lFmqlBT2ufwxwd8wtbas5mDppBqUFNb1eyTmgcPrBwW5hhGCuQ71DPNyLvSlQxVCFLZU1a6
P3tpDAS8rig9ewoMCc6E5kJwbVE0LKnkgifprV3eodOjoXyQqLjY5NmylLG/BKUD6yM8zdtLq8Q5
e4H3MA8M+eRP54K0BwtMeHW+X8U0CgkvL+hMJGT6mmS9pJVhsQQ5zOS6szWjCNQ4ItaHZc8663d+
sdCoXormXVlCZbJkhE5G/PjP38AdBz1FNL9JYEYRnE4lLeVQ8RWbhIIbOpl1VO64xV3iXlAFE9fI
/JGFKVlSJ6v18/b+UMyrufrWQY6SMf7B3JKZEhmIhl5jCZMxuem29Kb0dQdUBMb61kShQmMDfdaL
LEcabUDbvNVC6L/jTGyBfpfD81LTCHCMRMPzK1xvAV8t4f1ce0KaVVG45A0Wlxx1v1sV6V7fHUn/
UVRFF4D7pgioA6dpUN0nt1S3MMmewvlXBEspdCDCODV2GQTF43ZFeYVW4D/b5tdf3qdwWVwrXbU+
IdR+8ANITJtNKTSHYFgldJr0efD909bCFWqCt4St0NMaN3+KUdch2oyGQRUmwtJ4YPzzUUcf0/hN
ixw6ibMs9EtNdi7/WcHnmO5Y3bJJQyLggA29FzcdkfZ5mdOqZAb3VXk4HWPDbVdeiXELMWLA50jh
Vcwns+y4pwNLqb1AY1dyCJJg9Y7PSLUa4JzlOQdQTRq+GLMpoSZr6Tq36RXRyGqLsjJmzWUEu45O
SS3QMg0vmF5MvdQR7pqojzYtrD5QoYa4eiK1fDzMXNFfZoO7xw5B/8t8s1Mmpb2eE8OUpTltn87P
Bi2/jEoepCxHz4Q4W24RBTidYlsr2+azcp19ZGSpWp2HQkImtdbSuzOqhfxtW8V3k8fH9cGpdFug
acuOYb/GuNBVt4oqfcy6HW8mvdyrSfCHi9/8NATixC+o1c+IfKs4G4ir5ULDsaymFGxobH4xJMSM
S16jamHKPr8QZtvo1//khIT3ydIl0GNlqk+89efGP3I1ygIPUOyR7ryCkkzEUAfjvWgzM+rLrt8r
9ymUYyiHXL/efIQ7c3aPnaNkRI6tJlPM+TX3rfJPS1JLxcP1JfOHtDK0tE6whd3H2ZSKC93Yal6x
Pj02RBuHVtMCD1snxtZF9cdvLMQAJneO+9R73aRMW98I++YJks2RvxVlUaenZ0ncQIUYUPwmwtk+
cLW6TcQt86y621eMwbK9/1TJ3gVQ7u5kpxtHTa+PeR1uXVay+fxofaFYUxXPXIfBwjG4d5C0MDkg
2aeeEJt1XZBm+ahDFk9NF2Bn5Glmb1wwB5H4lWvMNG8olVLO4J3pK/3VtEAaKosKcLbFYE1mdFHp
16hBwkNO+cZsk+QUxoKbh8R1JgNKrkxMCQb0tdKSy/o1IJEmFpLRi8kZp+tC+kSuEvPfkkuedAET
6yvuJO4lZVKtTMTDLhd0S5Cw86Fs9nDZ6NJhfEa3uug2/1Ve7+VrGdLmD/l/s/IUUNp94cb4W0JV
hHcjVRPaHYFSZg9UOVC40xRoEUkbUI3DcFD3IV6b/Qp+1tBE3TAkTfgVzSvje/tmnYue54WoK3fH
wh+01/3rKqaA6dpsqGXTZGbPXhtYd4InQRQmeMwiWt2FLnxWqJtqIeCtyvghxTfHKeeA9Y/RuOMO
Xv34DNuNpSiTk4hJ9VOCL7i4P1hcr7nzRgu4nRJYKgSLr9TXrWUGqBFlbqL/7rqG6ZaCCVstitA5
g/ZVe+LBEAmFZgkSUFk3TDvtOyeJu8l6T6fFNFO73a90FxqoY/6AEL3O1Tiy50Kiz0wNbHTetIRt
MSuK/2scWSz/ry5pEqkIV+6aEkv5a1vTGEyVrxck/Ia8fFgLm6dY4XTKjiwKWJZrXNq2pco+vtxc
zmSsigK5qeEZF2Zq8SjxjSK08uN8BqFsT/ZUhiebs4xlJMLkN1Y5+gITXY1enGS6b4xyTb6gShWS
No8q36oeo4+JEohAY/znJ8IcWWC/tCG99sbekuiuPYx5HzdhrNF1xSAq6uhBhdvFgeVWHqNG7s0O
DB1Xp6gguyllywwwgl+0Y03hCPbC4x+DL86/nun4xv38iu0msQWyLoD4vmlQRYmx01vO/u7YttJ4
n1OjGoDEVgs1r1zMFL+Ax6G9ohobXOYqLMlN9UMHBZ819aJ8O8bujCrueFVpzRg337gAZtMApVIl
4fi10V5vDBVsOR9PyY1JWslGYr4YIdgbLnAVhVGQf4HMuGiQIoY96/jXdaEEDShiYU1f9OBQJ3PH
xIaU7luCxH/kG2n2DQ+gr0lcn9FMnPXD4p0p6g+XZ+FDN2iDPFkq2ONjjtMAW1Mzv7YGKOtHRcrr
h/vXMz2xxjLR77QdvZzPE3XG0deIC3SCnjpBmDKBFpshavnoCnx9akGJe2A6jTdUiNO7gpVje+93
ZoVQatVtIybd99Kv3gudb6A5AaoeyP/OXFjRGpOH+xz4RhY9ImZ1x+cyNbKoq4jtP+kePbL3tzv0
lSOlTRahkgDNqZe/cfkt/BI3K7vNpfencZSpOr+C1afVJFSOGEArVfIUy3WNbpSSpW3VefnT9pga
iqvCxIUBAE/be+X1udXwnzGqFpQATE3OZJ4swkcb3ktPtvMh85UlGyohmd8E4KL43lBIYaGDBEnY
9NSiEtOJ6k1WD7o95giDkpU3EmF0/pibyYAjmXEvslsJKkTNsnCHBpTyVeRbOABys+bNyWYWCgG2
nGbNIBb/5QLXsIUfIpyeEfv3s7s52Ebh6ONJXF04PThmXEIHUMy4s5sze1WwrObyFP0p9JCVvEoA
u75shc8/YRHgQ2HNRLEAWTL+hcrWpXPhTqpj+ZuWDP41fl8P8XO1KkbdvE15XBD+2zxQOm6MfbkS
YNcAOW67EGz0qEcOwZZ1p2Xm3jjmeoHN50O2rziVFUlZ37YPK7wqUVsn4OdMcJhg+2eMmZc8Cxii
ibjzfU46GEm7jw9tg+XomGmvodQaeY9uDLVnsrWIqHIX2lqm2L6mm037w2iARga3BvogSpCFgLtI
4UUEhO7al1ca2Hc0fLwSCOh+kfNk7V1LRNF09AjMBlBZ+ZS5Kz6QJbAFkGErShJnWFLXgufZvpHO
XTJ2eWamn3/DMtZsUrktpeX7bR7e5b5l5BrZsoA49lFLU3xgxaI9GVLMJNWTmptzz1CQTfK7qOpV
2PglBVd9CK+O81hw/5VI5ISXYRY5/VP4WYDafFcxRl6v5l6wSEfRpfQ5sHhjqYIyu1w5f8sjhrA2
o4qjw3mxFWCwwuV5MN6o9cNeLn0lVf8wvn82EWWTo3IURz+hvMKm0JeMf5AVJqkLFDXN3Sn/pC+D
g7xsuwgPOcDGHFVIB/Nko7k6CO7GarfuvLgYPk3RoCvA7R3FtO6BtD5cl9wR3KN/vyko/Shleyyq
sgr0xt4path3xSfud8soQ7+pzdSZYUYM4ZunAW71ZjR96W+mj28pqunhUEtTAs3fxGirSf+O9E8I
h8NCoe6YEvwAGpMYo/R3r7fGRSrD4/ZCHGujmaYN1+TBIvDd32hYi5EcY4tsoLl1P75+9Afs5j0d
kATOS1DJwcfCv9noyvzExADqgEfnjuyAhHbGXQ7MTSYJK4nPesp+V44BDInggNBcFgnq6kdf81YM
MQea6EfIjZQcW2bW6x5omLgArXN5IVpOY60FIHwLi4jwaXxEYH+80HtkaCMO7f1QKT+/7hCDGowJ
IVZOjwA8DNzP3O90HNC+UIar25kI2UtNFJiHKIYtYKcSU5mpGRPDTSBIQ6mjF/sraXF9cBOAYQEY
FSxSZhYy+9XhI9pZ5DG5JIYV+19uRPnQfAU4tGfL1MiDoCHwB/Ztp1FPcLJU4dXXp28M7vWaV/ws
/kbc9SMoGXcFWLCL03ALxDPE22bOA+VMpesWSHqRWyy1q6aMZ0+uhOcVUVJfB6e6NK6cKvGd2xFf
0/bIFagn6k1RuPPU9xU2OCUWuZokKJCg9a3HqpmLCUgoJzstdtyTkXNvMtxARAFNkjSx7amDYzFy
r1trP6qS4NvEtu2S/Nr14QqazpSimEl/5nDKLpiiY57BV1Ly8tDPSe+b+Ouq0QubgS1QJLP8kdXa
NkbBtF3DUBVlaJFug5NqswZviWEvYafkp/UQ+axeJPZhJowbxnSFmpsNplL5I+BmRzKdvTV35txK
gWxXxuBBAeQ9ifaNf098mmmWb07+ITolobEXgHn89c2M28j7uXn1hLLfOf+Bx3oDIeuzkbU1wJ0a
c5gyoQ/iD2ol7Ra9QIVm6Gqo/Ean5SnnYdf/pnaVkvSlFk7fbQe5cKv8YDtCVi43uz2AnqHgmgqw
0RZ3CF3v9Vfrq3tccUgoFqCYEWa4bFAp1XLUxl4dnTKuyMgeiuqQEe31I3USfSf+cxzZKhnIA6lW
O5sfzOF+9qyzSIgVPlXCvWlUVpMkcksA3BJq3EfVYbMLPyBGnL5H1fTlUXscYparhSydN2zNeBB9
VU87brmKEwQhdcEsFMaeQ5N9Ixesv9iyEr3gWtEo9k49Vil2APWFfnPJD5f2IPpArauKOExK1X0m
Yxjeb2fHu7ljpteLWiJUchlyg+7ZcrtQU+ztaw82CBCavcJ+MuyGLX7yya8JowHsOth43FKEXKaZ
WuQ1GG3SP6yw5Jr9KJIFPjh9JIgbGt/S570LtYItD2VyR5uJ7dkPo+Yt8pXDm+ta6q53QuUVw8JS
cpi3yr3z3JP45WCTSVCiZdPRE0nYm9Bd1lNviL8e5NLOiA1c/V+oxWx3af7T9twgDIQtBPLTdI4z
oxyJbUnbt3J94yOtw8Q9X6K/xkHAl0AnbYsNq87JAkfeCI3Gl0lhI5w7Cjd2RIcRPB/XqQDnM2xF
oglpKq4AoPf7IzXplWUeRyeDnrkToECmtmplR4OAm5tvJu57LEl8O9WxV8zIqR0d2Ybh+Mr++y6d
Xu/JxpH+O0aJduIHYRsTUNouX9PnLyVxFFFHmcIBZj8bv2GTVlav5hyriYrZiDdsUuVQIneZb3fZ
cCldfzu2oKsLznuKa7Hf2Ez75wEoBzsXpYxJoSQVmGXZUj72S167Jbsnwong08UlInPO7QcST+uU
9flpwaUzQRr6Go91uirI1lSEUzrOLXawTAYgRHzIVVPpOxD4z2hYxAcUlfxRkmtKmp6pmP5s+Dx6
ecI9SI79R7flGvMVXBPRBhLiAtl5pSkFKl/dAV52iNuwEWNqWpxJguhRROO56PxYgRqXQ/FYjPpv
sqqG/8/IRn6FyPReL+UphompCSHL57PhytzO4SKBYC6bNbm/BkbL4TXJVIPzzlD8X6MBBxL3tJHy
PQMhkHSSBAd/k1It/a+Jx74ZVtOhHqW+AzQEAeNixiGqx+3wlrnYkrtm3/6AYKmw5oIPpFMegMv3
IXi457bxUUOzhXzoLAdypGUlSIAqyk4SsBNAij1Kxy2AGrlyjHbuCWjdXjfVTE4WTjqDekal1+BJ
Ee3cxv7doLisaYtNjLDpQKAA0MFsjEDs1pjynSlmoNQFizoUBcBjXsOWkkdmuDCLUM6RNS63kuAO
BgZ9XaPJSDSmv5kF+5QmC9qHGQL6bs9bjDTh/+5KgXOCDIUfME0yeY48fDHpNvXgR6lAcCtU0FDw
b3tqtHep1SKJ5FpMYGhuCgZcq2RUU1IcKN3a820W3WfQpZsxMBQWk2gJJpgJEDYjnE9xLdREBJpW
qtrF/BvjYlMBiGOUfiBGI/mgSKPAS5TgrKIXoQI98VD9/U6swiyr9/ps3l0GobziR9Zv5fPOUKh8
43XlmiQrMYPtHwyLpn25xrDtkIvG3qY4lrXX6exGzKKbOgTjXQgi+kEAeC1GuytKSl9dlkDuagia
afrg9CiVTit0Si55oVJ2BOy1Lxele450duxcj8CSfL8tcHXNltDxpvi0C64TyLaIhJ2KJHaqe7RW
yldErNgObWb+oaZ3/8MI/tooc5ENXkkOp+WuFQWxC9wx3XcQ1+K17FhxYnOoruAY1PlTBVmkT8tt
CE+kyzP/m1oj10E0BLqfDtQINjkRL62IZWbbTLk0QxNhbVcDMUu9pCfy7r3CKQwjyhEUZqZ9gf4l
H+7QyyK7YBtM3lV+6H0ysJZKC+Kr7DwgLEhLwc8iMAfLnInlbHtxmlJsU8v6NhrO9AAqAnUE0QqR
JoJVOH1YR4YClG+Viyp/4NabbRF4FK67pbKIxhgnlwxxZ0r8fsNLHssLlmHy3iWboEJhYkEoyjfN
bxYMSPCYY20hjyOPGv0pIMPj+swTgbEF1RoTKeIYciQQ+10KtuAyLGthixvQK9wd2hYm/xIvHCpL
nbxjuNtFbIBJrxtIy8yxKDhW0qd6he7tHmMc3b1ng4BQLiW5PbE5KqxoTaPpQ132BIr4N6bb920B
k62C2n0YzBbDxzycEIA28uFYzWwifzrO/LxLKuQJ4cbKu3p0jnuFOjGs04LRTsltrbdkR2GgzVJ/
6qo3bwGbtjtYqaDepJTVDxOL1QVeYIGVCSMqDPDDV80rUbrwmekbbhRmDwdb1OGJjHHCQ2u0xEcm
Bs2gBb3x80sj22jEOp7y8/wwb78O1VauYGNqpmnGijHlFoFmNMnOP5zK5c3qzknZLWtv2qJ6MkIX
0+rYyEvjQyujq3ZEj0heNKP97wEs41kWmZSxFEa41mf5g4iMeN0+EKk1wA4t13kskAtYe+OfmCAv
49eR/P8oajlun8ALvO/wn2ZZvsbjq9Q3eDcgxRprCbsUrmtFQ3CSY65vsVbQS9A860ADkOLa8XVc
fOPOY1k1Lg5yrKuPbcke+dmzr8ooI6UlQ+/htSLXI6aSKwVB7YIyJqKc4Jz0pBlx/IwO5OE33HgC
GymJIhi1ET5JQn55He7GdaSNX3yUF88lMlkiV182H3DZ3UgbBROfqONiRNlO1SNWJUcSlWENkAIh
0ml7hnf0Oh8uMKYuC6DSPvvGZGHIQiawysmpSlrg6suzlVpT7TEnUn2VeBN44GV0Xi7YX9bp7WZ+
QxH71hqVEgFY3xJLqmvwMUTbOHDUk50q3J8SpSvbdF1KN3WngPdol0P7OKOgb1cW+b3BAAh1ytkM
naVuZVX1ESJIumiWwlSGvlEH21Xk0w/tohsy1b8Z0CarmGNKYMsxoN8mKxns6nxYMAiyNcaBmMj/
DA7aV7ppFj+MOCDbpnNgiNmE5TYGyPojXPrLQjoF5pseid9H0+bQHdDEQDpEwzBWb6EqsEr4vewR
q8yrs/StRLpPQu4prpw8HwOxJ1RnYBmbsItA7dNPZW6c1sOAf+/VV7xiFtdqClsYtup2Yfp+/KBE
oTPjRaitPs7L69aV2qWsCn4zN8gAKdF8lPwrrMLPU3h6GWgww+IFzJwrgfWISaAF9pGJy9HMbx5M
8hznXQG5lJaaAkSAX82oD5QC2DYUqbP9f+2Elely+XnIBoCFWjH34Bljmp+6OmcN8rTTCUv8BEkE
vF2/Ga3Fc3q+XkAgtRIDb7w3vI5Knqw7suV00zdzE5zo49ctLWzIe/W+R+6UxbPXYIW8BXibxbhI
tWYyB2n6cQbRxC9413nGqSZJlE4YfUYcTzE+zurO+Y294kAibZFQuzbVZ/eUrBrWxRAsqG/ICccg
d6Eu04lrxt/IUrkj6PxI0IckTtaOrsHrxqJa08i/+MNqPfILY5aGVN8yBuT0ncTAbsIJqC4xALQ0
VSpb1iPAcAfHL84+bAsNIWUI2A/Z9EaTjJUYYyk1uAy1/gqd3v8UEA8sB0uWWQNtQdBa0tESIr1T
vSF67PweXj7IkqVu1okm6DtZtjyPv+O6skie7XwS6JYcp1nXHMEFsyy3PeHmHtDmpGyCLpvMQ1sc
qc6mnntZsMdkqrbS8J1R8F1PYx0KFSwFQSd3HRfvIvzyPqOPT0r3vpx5YfRgmxkxnRfG938C178q
6ne7IxRE/B6dQpFH0UW2P2esGWtCpJEDC6xuPftsj3p0zBxg1JfDwKIlOvJrH4Z12iZSLtCixFFO
vcqt5dxaIU7+ufEVz6rnfUVzqoytJejfCqaS0DIKfufifUlR9QDEZ8tfSPU3V4k7mrP7z0VYCjnq
ArUZ2yQ1toVhO8Po6E0bmuskjwaKFd6GYbOwNQ7UnuaJEFi3WOV3ipL4gLCSE1ZdfGo0kCC/CQVc
4pQ7LAfIgCQQJNOP0Gun9gYsO/8BqCxikym8iN4zmUc9ATYyqRh25S791mNwpyNsQFd6cxSeB8M1
oSQKp/m6P5rNfoOydi6qlJm983Oy0KnGm89qQG3YQrlOJVbMO9z7zsWlNFLk9lsJ6ovMwnSA/H8O
Wx0le19xrS4h+vqlRz7tl11cj8dKFvqFWLDYt4vG6S62udTE2OOx9QST160z46BtNIMw5C5QR71F
Nn+iimIDhJabujnJ35TpSkpimStfj881ihRDwwTnvAnchen99gkrrZll/U2Ujyy6oYGXq4wopWzM
IVNAeo3EV4XhE6E5ALg+MxJZi1CUJsqagrrHUfHKDB3EWl6+XVg8lSoydh4J06l5Xd6FCGmRGgYU
1+f+aezF7ooXjrBVzDeHcYvEGV6LufYxVr5ehSzIHjtkx+38BKF2K7VCiyjn9g4LsfKFx6Uwuq+Y
koNH55gHLf6lmcSiwbZSX6ffqAW2xhR9EnBAkOfUG+FTaZskWlR3v54mt7nHJZ5znDDKhxzpnz0P
a5yH+ZNEVH4iBX6X8ziIGe3MnXtj9Xp/i5a4zZuOiDjeoq52q1QX9SZLVRo6ZlfDELP3FHXhfx1q
xTx3z6u8MMAwgDOeyGM540xN++BB3sTr79hJydS6+M6RZnOCt/Kb8ZAFLM6VKEOojyKEX5bUQrM3
/4wFFBIbirhaJJ3VR7UNqn6flTOw0sCHhTNKjaYQPv97T5jnjHqOmas06Sl+uTu47R5DyijEadsS
5VpceA0eqUCfr6t+lH7TVlIxpso/R78btmHqdMJ0GM9Pd//+x2Uw4QBceCpOAGslGwmugFas+Cqa
QuO+01tScCzPa4okv9fqxRewyPGDYG2voA1f86wQH6DbSStkoQL2M6rockq2WIZc5x9HarHIiMcb
4yhS/pbZISh4bckCWsJ9/WlUn4W6TAXniVl0kRCqlW//xt1kdk8T4rWFBMif3zo3/gQNZKBbjrAG
26fypmWbdZzMYPTq+X8E7cwk0y8MUAKFKbt68MipWHkRICQPSm4q5tjEovRSqJJknSf4evvFXHw1
Kelzie76HzrhlueA1rfHQYaT+9SYMjY0gUlorxbjrKkvCDNeBJmYVtQSLaTm0zStWVpKIka2zI5O
f8tVFhafAfm9ultZ2hz/sTMNzP+lteCwcv7tkJmwaIxzLfWJPz1dtDOLteoiQ8An8xQzXb546FPb
a7pNshR0UiMmMRDrjkq6hvOOFQahl53Mg0tUp8V5ympZfF7i8Ib3w+LKztvlvkVa1tzQO72+yTpN
4Fxl7wCmOrPJcJJkKbQ2pt/st+TMFfHSJPcmoV+omd15iQmXzk2npzeOU7fIie/Kcw7evPCU4sFa
jKkxQu59PE6MAPFrl6wBXTgxcUH8QpV/2n2ho+SQnGP1VmC6v0LpHBHEC6LG7ikN9BkqJpE9ZJlH
6GK6L67RBy9clvkhlQNQpZnt+cWFZ9K9kCUwt5vI7tePCU0fRcrsk1um8pqWK6Gd53oGmglqFSbH
ufSpKXZ3tSAbBTv9GZ1veicEd3q85B4MesrkWwHsbeGNJyhLfdCL1jeKPBwA9hbEK7IzHnlEIKbq
PVURKx7LBrneFCdl9c7lU6Yx4l1oiZkKtAr/xL393OM/Z/3CJLRBzstrgFQNlhClWq6uB4Km+S2a
I204wzpdnIA8abZgp/7Q18NXgur0jEgnDT6M3VFM0I+pFX0eAKMkzpVB6zpc2w6/INEc4wEk5pTE
SzbCELbHU290sTzCQLOaZq0o+YsMaPh76JFaDht0vGjNE2UJniAvImTf5oFuw/QaDAazxwO+l67G
AHvn+vtghr+VoaPCn2RlKlwPrwoldX/Vr0+vykhu0i6MWtb7/1l+M4JBcUAwACMOyTLM3286i81b
3QIjgTxo2pXxqGqtCgUKSuErHBBqzTf1IO/iGJeIYtNGerNNxEWEVnqJMLL0vBQ95yPma/FLikxt
fLyLkIWSC5R64qqpxgGz3jpO1abt/QsYf1KrW/Uz4rnIwT7Co2y/T4hnv1q3pEvojc/UrmNMzcU1
+tsrvyayE74FvUY0jfnY32o1IJiFUkoZWPJJaBWlW6SoLOoUmOs3bIz2Pxc3aet7EYn9RsFEL2ZF
bfRKHwniRiOdIxwR75Wf3nshdcBFg8u8/q7UHNAWJE+zfyEoaLPXfAfqCny2PrG7vMEtFE8azJCd
vrJsXxtuCC7Xc0S7VkkCYzcbjIBL2+R0JUFdJHAV/q3SG8uNLhXSieE2INWyfc40haUf0yt2ChW3
i0LWewj13u6yrE5TEzeItJEMUoPlJHf3mA0mGjxET3KV4xHJuh4PwOuBPvUXtLQDiSMhr5Csi2Rv
xYjmYnk0ShG+UvCN7alQhcKsymJtusTG7mTjNMzO7XlE1Nj+2Lk6BH63Xil9jHbuI2fpvOJzcuZl
hhqYavYwY7uRJl7FYy466TXJd3nMrp2/g/bRWgJMCZhRy48Q1bmu8buBI2TGxo97ki/TbuAnEpjE
XO0PbXzHD3wFbfnRY4Ed2jpqaYBF3zkPC3WIdXHGpTe7fVrmgyCvHN+3VdteEmenJ+mXdQ8EEllx
QKT6szhqAsIDsF1p008/2QmwAynwNbMLdX5E/FO9Q8rffFImzVnapxCUT8+Y89NbwKT0j1RzHK9W
siqw2zFZMq75w5hgnMEi7I0eNo766BvxmKo5PMTEBnxzMFaHcjqclIvc6RHVi3JhQCZozgnW59Hw
r360bfHQ83XaZyLpe4VRCTP4XwRTBNxr/oyp4q/o3vc34pp+nTIA0lM/oVt+FFth/qpeOJ9Lo8uJ
etLDCR/3tJD6Mqq7THQCSAwF6PbfVRitv2K6Bh62sdSuTHmF7oeK/rd+Mh6bA0DKPjMUaIhmhaqA
ECw7wNCVqJO91Yr5ut7Z9gB2bQFP9nKxowv7WG78m684JVoVIJkMIrwXMGqtE2tgQCgldk0JH4r9
kmIQCQKA6mKjAq4ZzWAb7J13+geTEflz71bw/aG/3/s7LpmVhLZw43ESpalsfamiaYxzmuYKudmf
UbO9NiLpdpXIY7Ic1J6Lv4lZprBWw1fS1OaGYmVqhkc0a/KCtyKC1jk6gr5Wx+bTvY5sNIloXrUy
woih8DNMebf0/eTDxfHhGLHGusyW8BbasAfzKVY2SXm67azFsgiRhvM/hmPr38bF/4bD1G6DhB+L
OToyk+ieRvdcDYoVH3QWLEPxtYtFnF4upHkpzZfAUATTLaBZwYDDouPw5s8ddd4iRQttZl7vIXSa
sRsA4ibAiuBhb6UPnYRm/SQUsd6NDc6xACZK4N5DiYfdj2N4a4rqg9CDTCtjy1WTmkIvoQibLT1+
ZCTgeG3crtUxQwr6JNxXUhYHPVPrjk2T5tDv6nM43lAzx88CnhKjM6yswVvGQdCPzKkNn4lRyucm
+TJQI/dcHAsi19byvD7AjakelMT0KF1JWOjCIBOG5CHQXy7EOFfFG0k0LuYAWfG10atwHdEqQZNg
Be6kNX+Ik8NYPEVVcx0lV9yyzlFPmLNZHevuruj9Izv2If2NJ9P06U/t6ltQGpN1INre8kMUhJhy
DXZnx1MYUghEgr5tVef2jpUIQ6dJ73tp8jen1hVIgFWjD70cMnC0EINz761t9pq4bZ99LOORvCj5
Yyh5wj9sAhRYeH+u/jhXJNNsTHW8/MHEkLovGG5uVQf4wIUEfn9Mg8KK6x3RlKw4qQW5dGzabhk3
bTUV0q8fMqCoQ7YhzwMAr6FPVBTYCgCdJXYe5ipnKk139I5LmSu6cGHvni0VvxU4wbmkRZfCjU62
EuJxUwHuFkfrj+pjsgSZqZ58XNp0iP0rIdgxwXLkuieFrh04WBTAwT82xDL0WOX6PFbkY8an8E8S
e5DDmwo76lcm1i4O0uImAHe8xWnJY9+TcrvlzRQ/ES+iugmgyklNjPCH5HskRQBuMIQn+bGBSfb+
XNUAJfJTtb7ycYW8N0OQ9l4c7wQNbDNAScN9foqfCxLPbL2GZhk8jEG8M9b5PsYwJ+hwBZE7byqs
a1hcr80h44O10IQ8vFzp7xQJhuOOqucytZ1jnCKvqYDLbcsw7mnB/3Lpa6WZyPQcj6gy2SPNBbDX
Dbhlw24PhXsFZ7flBv0B7kr5N1EfeSk/bedAizgVsbS7ggpkSl46PtcjM/9xaEI1oJr2uyPa4a5q
NugdxoLhYcQxtYPJLCNHfstM4m9hTHgZEzZxgG1rzhtzR2TwybQIIOsnDQYll1dWDP1PAEJSffHP
eW1y/pqOSiPVfOVxLhYKZJSjaP16RUFQ+isIJc7BkpNS0BGWxws68bxBIzybd+2bb3z8fS4dQ9pe
7z64P8BeZJ5/g17YTv08rHC0FFSxHfTDGykjdXqM3efSYIlsQjlQnvUmxcGhp76g3aTlpEbjYhOq
Vv55ta+0+V/wwuyOPH4CP9KhTnHrWRInNwHPM/oxtK9U/twmzlYLMXx6KeyUK0jA9TzFXCqMN9lA
q/X4gdDCQ+J16ExXznezVeOjP89ECAtvr5gNvXLb00KCtd6BxuzvRe++bNVWO/wAFlWT749Syzvh
rhpCbVljzOm8P+yzVcsc6upJeM00kWWwfe9X22/EbX7PQeA837RZ42GMd4Io8Uyv55QNLuSTJlMP
dfBupxQQZLWQrEG/2lT4VoiYP8875bdhyTinqAW8tsP6JT3S56gnSy2gAj8I/lxj9JKXDwmIn1XW
HmJ2PGiL9518UCozOV9xO0BFKW6N9YnhKwlLmN+3w4bNmHLOhFyAgD39YpUquDdpY8kO07ZhId4j
glXo2FG/RwPIM+8vEOtZmKMgG/1MpSA2fttjZyPQmpSaTd1owcLxP7e8auXr48Sray/PVqyEJ6Kv
pAMFVHl6CA0xXvwYuj2csy7c6aQqV/Nxx8mj27G4bxj4JW3+ja89R6GKlwtEPSZgZ1o6ByiynlHP
sJ6SomWvIlrul4HIGyygIhcX+GCmc426l/rLyvBf9ybuUXO2GFp538jdvniJ4HZ4y2nIeM2tBRrI
8bogULz+oKi+kjWYHtTsJriKVBgmQPhY+FZeyZ3eWkpXLTocOXvwoU0sRODgxw8VHS2lPSvNtGa6
CIPODclRgpFciKqyTh9CkpejwS7+pt5cQYfTWkg4B/3KVArhbffc9hDf31YSLeDzgE7HnHBCXi2a
h4o9Ddrhil8ohJQdsaXd21XJj5hczVYRXSmsILABm+Twmbdh8ureKIJpAEyjZ/vjKCFVRXeFfCR1
N8ofyuT8X/eXXRSzHq+puMBV7wR7GCJiP0lzSd/nRGfK7TEXchfyX8zY+QN+0Or0MPOc2v34dkPc
jsXoa5itn/l1tHQDPTTJHckSqgBK1AsMzuLwP4ZbiIXzYWC8N5wcgrDNXSYHOtbqLGC6P8EObqD5
9Xve0KhW64AP1m1oE0fwrV7RLNFE1a6fJaAvarBcoNS8Yi98/POA9N7smZ3ooJIB1HOWR4+0/1Oc
tPzghmKnSPiuR2AW66EG4+Caob7Fr0AbwkxdNY1gkmtKq66KjQyPTzpdc97dxbH5FB8pzCTW0AUB
KCMXOvj20aCPK4xFP+sC2J6UhwqpiR/hO81hkz7YSFWJlmfD9GB8mL6fpAZAV8UVRylwdswsiE/Z
TKGrBoTB5xGPRSWXBGsly7JaOmPjMUwuT247Cx1X2IhHqecy/P8hR+RWC8fxvGwhu6YylrucBpU7
JPQjXk35AK6H6tZKJ2RWRwC7bTolWw+Uvk+CNRiPvq6S/MoOBvbyqcnpYdtbzJzGmXOiDD+zjj+W
5TNsq5w5RD9HI/WnI9wghR9U8e/xAbSHQVRfCVa2WGU/691nqk6vCeAO/uDk+KLVTvMgxbQQi6WR
WHRbyjnUVPVKBMmk4NSRD6Ds7klo0ZgNSvedJGqtAkhrrRDA8wia2fSANQCQJB0b7OJD5oWCcADJ
eSAVne9yP6EQCjygwjMyk43+GOeOyXYPBpACyQsHVCJKA1vB5Vq24CNxo4Fqe+b52d7z7VRf+E47
ZayDrPGCqAh0/2jO2XxIHtKI2A/zGNJ/TYwEkGvWNpq5GDdiosp2pXZ+epQZjRCTfY7n8MEJB/1m
tKoO7LeIk7roTtCGwWaX5AlljUZIhMSiQA8uxjox+wlAfEbd1f3wqXlcfTwxK/gY3vM//43r0Oqt
0ov0yEuVqEv7ObIoe6YfnLMPcvPL1G+XaHRLtpa2DR1l9LSfWH8rrMs5Ith5VztkoqAFU5jph+jA
IWTnwl9Xrtc630EC1MNXNRFf6rf8JTVs/iTdfT1QmcquuUrrLMd8Rzghg3LaPa3+LWhEKtU/w6tP
LCt1HY+mjLwIHjp3ti9eNsIX/SpH/jS0Bl+sBLRY0/YRrkdPj8Tja0JRJKNA0QPsb7WT85/33k+s
9b7jRasZYS5cBV03PZ0NdzzYJQoW6V2s/C/ChRQ++NWag9hEPN9Ewe1+GBszLxiVGbDzokmJPZ65
4W7yP74VAmGRmf2OjuWy32TkSAuMErfB46Fef/PMlksclObtnTSaIB5ry1YTm5TANTgauZUqUMKI
n/q3NsPJ6vsy8ogndLCrb+XJkZ+C3eij8YSfDyvS/AN+lsuZk+tDP4bUEispNqYV4hnCYgIZK5c/
KvMax/kjz4f5w/SO8iuQMrpEWqxYDtKXyCXkLMDE+rSFIurDWDGHAix2ubet+CoAr5znBXMxx2oT
7WJWmY7UdIEQe4DAnB/jbiUPh4B/dNQODtmALzAPmkO76Su41LTgp4jWfYgYKtn6BQZXRYJKFrhn
G5sUvNZfMTLXwiqXGH0ne1S3Bc4pbvy2QSaitn8twq8ZCpWjXTL3OHCvPQqDj/RHikoYmN5SASIc
6tX+Wb/KL1ukbrDqyJGeV82yuXw0pm7vMa31rz7S2ZxEA9RdLTEUTOPZzbNNWYC6jYotlQNU91KP
/mq+68cX8ACssorQETymeN99rwC1aOUDKBN4Dm9eDE5mLBrD0bpMuvex+XnFLiyxguepmJCuPT83
XMrKvWzcr6lmyP8IPYNavSTAgM+RB9PpbKzrBlDVTaJ70R2B0Jl36OmR5nHLZb1kUKbFJVSMV4o2
gCOVwgc3CrhIDRlgfgJwlkViWaWqHghE/QB4ybZFJxdRA9Dwdkakzh2L2nIJVnQv6JeS6cdJiiGp
hEFc04ZZ3ssk7HrK1Kr0YCyVHFXqZBF/xuEM5HKqvWXslScce54sfpJZHq4nYn/P8U5DoFya07FC
MBN61Q/wBrz9iE/2ScTslBv0geYiSaeKat0fSrQiY0W9z3yr2fKkQDIwVtZLZtg2N7hTP7E9Ujnr
yvTG67H/orAjOTlBrAa7zG1UEVJq1PBXKiu36J6Jm3wwz0y2zlWN7JBuqRWfaVKay+2pUeTbJvRa
ydr1rpoqL6beqhc1aMDzIVZZQSFBTtDoMB74mgbZl9MzBgMIy8iuRQo4cKxAN3/Zh7gnVHIVeYUU
o/YuXXUiBBIn1VTh65cA/a4GKNmf4aBt3objP9QLMV39ZApllMexcYeJMIGarclnl772qoWuydc3
dM7Dfv5ioJxdObR/1j4GSUuPaMM3ZLR9Uh3s3+XMYovajQCFnLBxASuCstJaUOef2oULf2Q2nZW8
+2C2KtDW4o+UrJWJhB7+axXiqtvHxaNvViJwgsGDB3HDCW0pXRRdYy/REeeYuJnZreU6jJs2OTAM
sB0h5nD/x/tJJwXNrvX+D5gZbs9ss+9oGLj7zWywAgXU3/6G1wjrDR+ooswHeWPqcLgdrbBkPAmz
5IP4DE6Aw/WDd/uBDv4Q4C9LPqUMaT46UwOWpC5n4GBHCpKeEI62R6JN4PynECx3MXYuIVd+1wHi
qFpnL9lbdomnK0rMMoCvYl8uFtD4isu168LE78vpZSSGnKBAMqm12G08jSteDNOkZZATR26z+3eP
QShrFyRXzrzYprCiazSK1X2joXA98nXJwyY7leI+747jnspj8rCMNh3wdAmTbijcBUtrt4dQU1L5
ek+KhmuJCQxJUf7d0Hqje2YmCen/sYA6jGjw9TCXenoW7/VBD25U/oe2A9C/d2g858e9MtzwficY
e6Gb/Q+UsJjfE6EOD5LMzjQjbszQu17SqAFdoMQyaxza9L9HcP1GQGVLNtegjqq0eG87ojQX+yc7
1kxmjICeBQPRYPyWEI8uExt1PzkjzIJsuYqs1ssTo9z9u+DgQydkf4Auf42CVi1+Dw2YQotq4PoH
qcp629iFdfm/3W1crQS/JpWVFUYPimChcNa3ZiEFBTw4ZDn6t6zbaIbIsvw7+pdr+YJ7ku/CWCeE
29cX9lUrulV81eTHyDd+rabX7d1C65ayyqK5Bw75m4heFNg4Y3HNaD5yngSaiKipt1Iz9vigqnut
TfLvKsLdhLk5FNnpTDvSYtl3HitpoIxjwH6zAbTshK0oTp5lqvtquVQQ9yP5k6/ox2MlZoKqScWR
CNDDYbnCF6ZUvNXPrGye/E77xX3QCiUgNvjOpOXSKuMk2JLxJtHHRNMtUproYMWk86pud67nmCfP
YnEdJN4nCLpr9+SnN958dO6+wZfnT56MV6IJAAhLtP1DpmVfJYt8P//aRTi0V8dbm0HAi8MK8eM8
0z7ogy0ZDUs1e49GKZ871gae4l0hZc+eBJ8sQZ6HfXFUFLhgvXWo4/LIxkzj7xitpRFzHtbBYohP
sX3yVwxM2p9wKAbKGkIawYFOJpyDcNLVHU/EaWaubAXeGJOJAfsjJeEShMDTqon3Co3u1kaqdUIV
AZWFwyaeVARKQR14/I+MsfljxQnDDG6GWEB+lYjfMRc91JGSoEcnbcrK6eiI5SVQNvnh/iGQqk8P
XpwNBNkswLiRp9IncIoWPNbx3Bk7vXVp/WdGgYnSjHlaVqmZx1/62Hys36Hszj+tfV7AxiB1/W7s
lkASFFHFDilGCWGB9c3nWu4f7B3Dt3sb5Z3meCdrXt6oJusS0H90hVEIeKE9ZFXIElPAl8BcTzEf
/KbrSH47glKjGgPQKaOSWEgmgueSvRVS21AMZNXzkViFHaftyBoEhBkScWm3/axBheTwuuApp1Ml
k/zBCShRcA398AT8JtykxK6SVFpCHfEIWLo5DbMfkDgZEYCTtl6kiVDQJNw9raPOXoxvG0VZUQgS
h4HimRw+wln8zQvNcdOVWtE9nwpGy4l8dMCjwr1UhgQCwalYUbAxfqErSLhpLYZvBdCBsJJURQ/S
QjpE/a6h0SGUFyUSgI26EySwDI7klZn4i/sTYbRr002tUv0sR5NIdx9YGfWHEXXPjxAoIBvSVfmr
EFvDSNQ4MNp/hceUcwBXRo46j11fu0KXcI1Pu0HkHtAg213xshqsUWfRnoNsEyQcs/e4EfxZKciZ
cD4K4W8iuEXi5kzGjXTX9N8PX14iUb87I9DVlYyTCUeQWBzdoxEKJWfxm2Wet50BNxSQLk40A7uZ
sZt/ks8No04ItgxDkPdoTLOKgg2hSH0fOQbgUYj0aRfFmksTl8SeK/XzA1Dn+lwmwr9vn2SmkTqc
KCVOJ5ysopLNiXSrT4JKXN1Bx+GkQ8ilw3ICGyhbNr1w1Wfr5c2G6ZT9oQ2zvtrOM4kh8WmMgjJW
1SpihOn1mYIYToxaWAF/ViX+x8ZPrXqfVK+LlXFEV+72I5eU2cTbtdcKSZTDQC7BWLbeeaPUL5qV
3Q1pY19EQbz+g3sxwrqv2G/QS65EtAloWcNRXpUBmQNKEldgrkkZ6N/KHCXyLrp3mR00Z75y+qkH
4oMAPwPJ4zcSc9aUEuGpmjp5ClGrh5q6EOnTpoDGc56XELG/hoFz/eM4cULNcRsaV6F0zUZ0EIW3
ngBLuBmpKZOK16fERJh36Y0bvL2UerilL8X0tPvWOZ8f4zmFhcgNumAaw6QiTrhrBLCK/sP1bQRr
dJznIWp/59XvjN7QHwmuKQ08hhDz/JWprehkN9q2UUnrysDS7DlkXh8vjZ2mf1D5mI6howJIC0fk
tdU8WAMun08LHWtg6TtakNo84AohSnAXGfFAQ86JeBOwfsBG9GS+sBrVH+v0zwym9P9sPLiVi0LC
eCFBJBrXN/dQsbinwOjIysBSI1o05X3PFxamDmnmOW+gznUEGRELepQLL2cthQJrv4do6gYEr28E
SHW8hJ7uq/rymqfIOSetCo3VXFQ3YtAjVV0AvcRkWy/bDG4TELSBz4wEnyt2cVCncU9bC2AyzqHi
sNAN1rPBkY0+kr0pqTM6vmwPs+qdeHTBR/Z2rXhIkMcBJmLk2/XXSOrTirsY1Bk637F0opnJdcaL
Uc+l+QLY566amobNAiOT+6Ox3ZXChPMIfZ4XczpCjHD50Wnnr+DYX8w7geTgGIxK6WLItFFeGW5i
2TXMatY6uILtvnifaFW94Fz8MOFYSoZFVUrA2lIXO2aAJax+gVUhmKZ+ku99hZU8x6RLvTxoA7YM
ZC9swHpH+2y4xyUjV2eiWxqgOVVdO9tvKNnZuOdULJeoSXh2a5tLVo1yjOdo0USrBu7ygTrRHatM
u45Vmuh2R4TFMbhBAc9hKT6q1nU22gZ8YFn8FaJ9i+jPHnqc96IdNMmS8pfEZM+SZ1a00T8ulKvf
o65XxpxaXMknBI+9HpBaxf7CJ713PNoLrd3nwrSxSvLlxVoxxN3RmbcAV7xqqr4L9V777L3qpSrU
f7Za8w+plSq0qkOva3gv2mGFzSP+LZdN0WrdL7X6bxhhnZOIIQntS55vkh9vDNVopHHAKE9vB77E
0jl7N2s1AWPGXGeaxP2mvGfP8T231TLd1CoVeLzEw3dsNJLTBd4YMX1KSrZap9Ms7/9HOaLSZ2b/
n7XuQgO5x8cCWbM/N8VSfk89eEiFIlwSKLKycGgHlYt6eT8KnmKVhJUi/8CVixl+KdDKUrQOj7U5
pV1T5FxsaMp2ZZMKZjT1kFkp+g6Z8qGPcFFp9itDWSobAZcnEvHfB8TYEBFTa49M7A0XoSwHk+zY
pIzOqi6MkCp623Zl9awHKOgsALfHIt63tfyLbkCOcncRtVL4lqhS8D9nBot2IKvnPDwjvDbtQK/S
5RJnwoGIfX2k0huxntbrQmkss2pgSjLUQ2qmKvmRNZaqP9cSq+UQX9OC9N4j4v/uIMU3pYF0jRa5
D2Fj8fS8B8wJVUfF1aN/LiEWhT6X+7H3GLEfkzBq6FqOASVYoYmxUi53pjtYD9i8Pz8Idnq6ZW8y
tiYVX2HkbB+brG7YAPc+QvKShXrrQvgHdhyxKGlhOsrL2nt9mX8F8lVA/WDojEfJ0oUrRAF7qVN8
9SudxQh7MGgVfMN/chYFfcR/HTv5HZyeX7F8o6zU34e6R30brVVuKnjFw3Kobde7jXrZhWhtZUko
TuYJOtCnxHPQNm16MRa7YRt7wsYuwrK42jW+VdPl6DCGWKTkgsXgCuzmgcH0++ouxTO8W0a75GHk
3NyMH9sfMI1Ze/nW5HXoaeDVu9iJLWEhY5xhmQFXr14zhwLjD6ztDWdHPsabEWszDw6XhodW70U7
tgY+pwWArZjvqpLpHQzrPnAzjGDwvEj00ipGiGEyoLWgb8oNAF6n6B/Bl8zwd2JDcb9JmLPpHHkb
OeiCxuKwYK5oNvu/gVoZME2BV/8WUFEYET9WouVupOIxnmrKka/bKPbKPiyWizbpSQukRMHb2vhd
owl7G1nv03PRuphUimk8bxS8sQ8j8h0B920oQm/QJjiIxrPuHalap1kIRLccqNpErHVyg3UW+u5/
koXNIbwzP2p/wBxNfIiGF5EUID0lbnB5soGVdIsncXdSn/LS5C9XonixykZ9erSg1RoxJbZKH6ex
/0Q2CfA2rbqjcmD1EKrLt2k5XhtYEEMpjw4CsvGBRhpevRem+rdiPEdXeqIN1Tmdlk1TxLCbcsZE
b2IP9yZEzMaUaj5WpbgcufUuSFFPj5zDbFiDVbju93Dq6s02KuzXLSKveZ5J88670tDJq4eh6Z4P
FzItMi5NRuTXy7Xd4QU0k0dBAgIv5/Wgv/sCWz7JXEWkjtlwdhPnnGELqU/F4j1Ay+Q/joH+2zXP
CA0a5be4WS/6LARdBWPWX9Knliy6j9NGzLpMiq6s8ysPkBZkGARzxcTBNLLrVpTPkR0XSdy9fkGP
ZAYHjrKQzFzUsA2Ag8ivwLm1FscaVL/0jZBYShrrTwFDNdNH5EZoh14V4GuFw1/hjDA+yn5fbjGB
CR9Wztz9O1FPJytbmyciytBVcL6vGKv8xYdagQQeX9KXWKyx5sIFsUHWX34AEQffeghYSMGL3EvB
EEJQi5veU9dOC4WJxtYteQZ4k/RgrAT/yuIvNslZGMhbd0wrXKv63/GNjUJxrrqSswv4rKxFj7G8
T47i47de+WaEkR1OyuD0y+hbMsI4FpH7GbIywm50raxfwfFgZEOaH79/Jv5Fy9JbVW1RkL3UMRVL
uBVS9hm2poh7ZAxVGc4qja4LotCbzKnPaYc4oC3/uJ5pkt6EnlMokTeLL+TCAZ22U+xhHqel6XU1
LePaKPGaAaVm3wQfhRM4pGMWedYXjsLLOkxTW3KI0OH/EaOsPPAcR4KC0/6AVsrVvs9srXIeNNAT
XG2P2wThlG7uqXGkDezt62igVKlrueJE7VCoUiiI8VwWjllHxrlawxh2bkx3i3vVz2hwDWKWmrXy
dnguldSkPcGgKzkPU2lWPqeKF0P7dPzQf6ahQS2etFJGPxtfbDmX5ckXowqVSPlsed1O9kOlq9Qn
HNUh+0nWm/AlEmYidB3IYRBV930IJlIyJx3BQGIbg/nbDyzOcvCx0RFvj7lsdDhMzoPEaw4VLnZa
VZfCBopXMWiAAkPU2+mWJPOe3eBJd7da7HPyncJCNwwRHtVYpbXsiiWmpGGtHzDwQ03P4gm7LchG
FFc0ovt8EgTMONTJcUg4nZyamoUr7N7Du5t9SqSHDebia50Dd71jLK9bC58drCnjC20L4Db4E/Lg
A+OtYKJIbXmKRcEN8TEXf2SAMZyKDdCYBN05SxpQwJ87f7ft3iyF+6DadJRSExF46MuGTTZiOdSD
ODqWTFl+GkrJ3RprLplxLAOhnmM7vIanMRnR94CBzy+WJJe7zAjFBjxsLxNBVa1tD8+pjJ8v4BFO
Idb2jGs6IKPitA6U0eMg6P5ejj4fhwOuxLIn23CMw69KHOzxAM1uysBC5L0fcDF99WFkl/Bf/uJC
s+VFXsSQZQW59J7WDZs9bKBijgMi04ubk99l0neQcItqvoz+dof7v0c6uLfd4DO6vLgaELgbUtXp
++FXUwX6bNDvgTyPpc0jygOuRwlRKACP9tq4d6wayZDTbF7b9r+uA8zt8pjz4SrU+PYGQ4goyIZ3
o0bWw7F6myDTafOLWruGHhDNkWY+6M891KDpl4QZySOyWhZ5DU2hTJCBGedq3pmGFqyzpNZo4S+/
Jt3gD9TXSwwH/i069nQUZW9192K1Qnb1fbgPyWUYeDAGH3JWxuFTEBFfvYbW4b5Wm7q2OwHli6gJ
a3luxBw0bUSs1SHn5PS5nnlcFNgNhSkudYCw/WdoIjR/+kthIpDTwmnG60ziBEv7ofXYmep8HpZf
Q6l2egWqhVjq5VW8Y1677wMaDAGXRdOJzx+XZXvptcqLV+Srczp08cswJkxaHbCdypCPtWFeMv10
iC5KBBSA3mzV7tmYQ3TevIxuGjAOfx/c59zHZKKCQ766KwZ9dE3aHejzgzO7eoS6jF/CZ/zC3NWD
H7jnrEprcFd34GMPbitr6+x6M96JXMZWkV7ccOefKuszxQ3VY2nU40FHW3Uswu67AW6yOXdxYI4+
zQXkgDIGTgCEiej2HPl6mDuHoYMdEXTZpFEHi4IHSJeazz7abISnP4MFFg0Y3eEGnFg51ubVjmps
Dr4nnPCkWcBR7yKB1YzrOuJSLIWVNZq7/7UBu/CMhSvQE435uBkDDFnS+xhuNI7ru4vYGTi+G+nh
AwMxS4XVLiR03Uvs7+zFWQMiNRQYw7eG63kKNoadwLyMONgYunfVFNNNmAO4IE3EYy7a078iB3tV
J4AdWE8JJUWBBEMZRI06PcCsUzK+4yeLImQYtV3LCWhoZd9vyg084ggL5cD+mBQA0Gj3h3/fgHVc
2PnNigBlsi8d+VllE+rrtRz1WaXzLK05Q26ch7DB1na+nCy1QMpJ2YNum6c7W/vYPQFbz3mK+F49
vUCuidZuDyLdn/aGimsewVcWXvMQbF7GYLMWtd8hX+kH3NZPeUfj8I23WdhyWq9zVXz5VeHKaaN4
853Ao3vhgdz6e9R4iZg0rii8KbmPlxHJjh7rqCvodeW/8ywCSSaYMe+8WBLuCjjW5UhlhHEOX+wL
Kiyb/pX0dY8XJdpR8gAFmFC14ncgdiuIMWcbfjG7QzlaDTnLjVl9kDie4GE+PE/nStFN+KtLopqz
DhMtj3T8dejyHUa3flF+W8jGSdwGCaBLu6dHfyIBsEGBHHe97/UPzq5cUvQKThmtiNCuCk0Vfwxj
NbAnrWAcVbWL+3a5tW3THDZhFg/ThjeJyWybfqKojDC9IbaI/KXvWcDaozDXg+IXh1sZf1O3zOF6
gCAWU/XPW2BgXXoA0pKTkckoq5N/mVvzzDsX2hwV3++3SPYl6HXLq8Ox5cvqAMHQnVhD7E5JTiFE
6vEGbudf2q7NBxxGlJyFhAFZ+VvbYOI0/DC3+Sl5O/lWuvOIre3fn4rwk/ZGPvE546YWZ/Y8FPuq
+N/QmaByvWbHYYhODDaxcxh9mOZZA4eUC7cuDbqJa5QihNoibSkQLeoAe8Y133vfQl9FLgmOykZu
q+SjXZxdm/brZ4z+uXTjRKa9QbamS9L9Lf4GNdUn32JCGCsnKgHvuyFdRef8XeBhhTd8QD2o6yuV
nMflOoMkQB7hPnqDzCzn6+rvg5yKwXh8ZgF28t5dOA8aShJ8pytyQPjqrxpPngn+0sbg8qIz1VFv
0FKApVubrrHhhACHuMeAndOetnICrh8Wd8gobCxSKlKzkPdcvBu5RJl/PMdZdmND2TaLenEhW5jQ
QB2/J2cOMwmV6oJyGXSLNhM27xahcISSis0uTqpyn7Hku9JVp40iZFig65XfDW4r5SMYyRAZupAw
zxYRv7gZ1aromXK55BY6j8CAWoRx+KEniyqc4wO1G+SB8x++X20IcbCVdTg2weTycJToRNhxA45h
nSxqmn5WLrW1SoOov068xHjobhPGDnf9GtgJgWW6LSxciKpe+ng2UeqLkwE0was85BVw0CKJLkeB
lNUOx6PZCIpQ3ZSAxAxE09f7FyFR2liXb/R4b8tezUsjPhVrynNvY5eRuH6jgReDmJfL6HBwnx8/
Ry8kA1Ew6qCZ8IsdVHp/IdaLREze4zgnsHgYbDnWEEqMdYH3dnqvs6v07NAsG5J8d+IsId61FlpQ
CcHTMl0IV1qxeYbkp8VdNmaZehdA1P7+uvFBT1NgBckyuxTOwSnseYPTMyCw0xud/16bpY3YTdIE
vQ3cr89t+12BZsFkCqS2Mg7vnLGhWUwEKGhVI1MDHImFbcbiJl8kPj/1R0Gke2TFBLj6ljXO2qNm
AQYSVu4eofYJ/rQMHsiLTSFCwHqdsqnYtdw82HD0nmNF4Wn01lv5IVThoZon8IFfD0fBYhodezQ7
6ocdlVybxhSpfZSFUzbY7XQqiRaQzFPynqZrOQKiae9okSwCW5dG8whJ82e3KPTiqY9w+KjXlEe/
629Zt/yQqOAvm3z4OiCdpRwyvWCo2F3lBV65slFMKg53bqvtVnmQXtVF9nRJNrY0Jpuxr/DJT3nC
pp7d4t6voUcSUP7AnfcD3IlTKQz8gHbPvXFp4u1SZIdhTpOXmEf1/6bB06naMq3zUVnk/ZZl7ME4
YrBb7xGriT65+6ko9Ndc7d5QIPCiXMUS7knmEnP5xr8Qn6J6teALyPsOIG5y5XRlV70MURC031iZ
oiVpYpQgoc/kmb9hX9T9lmMSIdvu13QTTcZaQ2QQM1g8E+XokHnMttC4M503O1siYKUIAeQofhl0
uELOnHZ+U05gZ01zVuRn7E/2ju7oRLHicHzw+T9rEu9LgpQcdYGXFrb0NwKVqXgLND7d6AeVI3GB
JeYHpeRPn/os/2qdgeDXdv7g6RzOzogbsJH4SuQEvkUVDm7zz6YqcEtB6Si8vFagLd2/A47pQ8Mp
FhwMqUlp8HBUW2tMAwK2VKck2xyBaO/CmMJ9cAp/guhGznUxtBetTZ5dcki0iUGXFgD8mlbb/2Ht
9mdDrKIxkX6KvPOW5W6GIzhT+V6uwxcTOLlqOVs7jlLy+8FbImCMdhzBaNd2kiWhuBwryNIoqxjw
gSOpRzdAwfE/8Cbpf2aWp41QYVIjKEa1mn+I2sJr2xUBqh84yPeVO+UCpgIeImGbkDuPXG1WZQYZ
6OiDe6XfPHU3sab2YTYx2nmtUtCE2joIwrq3jpSvO0UC7OC70OifK6+AQFJk0B1unE+fe3aFcVRZ
UbWHFMEEFfHXe+dmKi/16V/Sgx+VM09Y99HirNTamUUxcdV8TPh24NeSREk5KXRUsl+eeSJpDu49
N3dr9RKBIVoMkbXxmqO3FPfd4iByojYMksVQqrWN7WJofttDkMXhQCNmQ5VUl2exeJv9LmyD8PcL
bDh8Jtf89T7mzD6UamQNVjY9LX+XHEqAY5/JBhrP4sTo4LDV/qeSUuQugdbJQp/Nl5jvYvyAJRAd
ZJnLkk17XBsBBuw6uts9JO6K902H51LwktrI5YAq8+zJ7BNqryCLS65iZm9FCpLpQzCRqJlZxmZf
Lno9+LYZr6QFP5jqfQUdkDy8thFD6TIx0UvrzO5vkIxBYh62UX6xMusDMRuqm9vmGxXlCPeNeGIZ
4+yLwiXZ9Bo65uTHf5brDZ1QWE4sJU58iRwJgeFGsyWpQKV7sstz3agVO+ZQYmHutTvHZnh5KRH4
ewHC9Hb5wGUtc9aTkw4RpBoKdK6vO/kjwM87Cv3863+GMcmiw/5DvBxI27OtnexQewlbyVgCQFbj
vihvCeQE+2c0fgVHrWb4EHWJHWQgPg8DPeXsH/hFRKA2VtVubOn5LIK2q7KkgLKK97ZGv8IAagFp
e0RVjFiQYql9IVHKHaP8HqrZATTMSRGzPFm7bUuamrBGJz5X9gfmyXXIXHHK8Qbv6VOhb1GRmdVx
UpQQjkvVk6SboBoJmXBhcYYKAlC5imrdlMfXWUQfMQnT+MeeyAsDSI69r+A7kWT/a7X2yZ+LpYNm
Yg7tpvoy7lhyvvtZT7/kYGoOtEOLyM8ov/P+0Ue9YtQE5OzVm7wFZCVtID6r9MEAe4N/0D59JnAA
CMcatXCdc87IYLfQiguPs/ACKw+ygw+hsPTH3hnKS0sUOj+UkfcuFOz0OaYju9qee4lX4tokoqdd
ECL8umv5mmlaqSG7DPl+6JPamO1c+EQb7IufQPdsWXr3qPYEe53lDSpILyZOsuGqNc8q54DiSauu
cCCjmISTfbgIRsKXixoG+T+e5G8y6KwnEWYKrn6T9bIVDSTAEcXZONO0RFEqs05tWGeFoCDj6tMD
Kw83zJ3k3giKD1tg+LFewv66SGTrAZvefqiDhXZFSQ/YiXPoTEwF7uvXyA3Nt5YEOjZt6KsWNLSD
l2MDc3N/V5iqn9ZEZ198wsQNETt6/p8BHVt1H4Jxmjt1DmtLQRK5Vg9uVSknfVkJPxjr7+3ABRI5
ZAifivuICeAIAQ82S3WZg6Vr4J88/oqzh7FqsDz3qjYRA5HIjCYThEXaWBMm9iqeZa3hFAgE7cqJ
AZ8L4UxoI1Fg2B3rtiBUhMJVdKoFfRFsvnZib2uFTp5dzdFqlL+ju9IOeh3We9aTC2gw+XVSS/2S
92HDtJCKA08PBnmY0XEny6I76FmNr9UFmSyd9SkeuAx/u/gy4o0L4CeZ/CBvTwFUS1vHlb2bTm78
c0aKixNLj+i8vX7z2MVHEnUkiIbU8Vw+/isNigfrccEaA0Fe3xcC1UIRlpnrgQ78yX69alUT7SQb
+hkrvCqj/XBS+tFGxYi7a80InnnqMQexrlVBtNZTpmtsNPfvhhAsukIptdLuoeICdhlL/qg6Fsap
l860Et7BOeMoqtZFgmAbXUClERAOFgcfmYFE6QKyMMd7KZWS+QOMrilhVXqECni/EMRIuqVZwuqG
+U6VSdYBs7DaB7AGItlnhcfybIB/jMTGAM2VlO5+cgy3AO6OQtU3GWKUvm8av2WP24T40ScJPd7d
pGw/OGOHm6wFS1OXWqEkE2LmykofnERS1RiC8FS9LT8/AKdKUVUvsJG1sAj4eorXAfVGiYIXUUk2
YQgrRQ/KFcveghxqy1E6ghNyUffdJcp8FR6SRerCHuI6lIl+4hSxeZMMlJ/gJejtk130sI2qgM4d
RkmDZlRIZb+lFD/J2czMurWPcLZ6zCnY+YQ5qLTisDEYfLwrErmc6i+NK4kBumetggJyU1Bt9WK/
5NWoKaVohmSxbtXhcPA+rX9p3ebtcZAY90Xz7jyi8WSpn7/puNffZ7Y+FiSpmGJub5OJfx7USoTa
YLryTiVu4BoDx/uRuD6STQQRxFjwvuVrGjAasukcDWqaASaUdvvrHNLcW2keFOLcInaGQzJuhdG8
CSJGlELl8MZ4xoGYCUeuJPSFGb2DsMFon9nP0Uj+mT8DJygCWLeD7GaA53Sugp3stMMmDh9A9/4O
9yhvwugtd5c+NrYUCswCQc8HFH1epSpbdc/I8mpazOpvajX6UZfsC2r7s+It81MQ9xyzficVRRhX
spa2jteXjfJ/HLf1oYM2Ap14X+8e94PlI6fhg3qJICY6To878qJ8NlJzEV3IrUiEevD5bBsOKxIR
pTH2xaNgKmbTgMCuHRaKS5Ok74JC4Ta3uwd7xWEAgGUa5xkqgjY6u+PPsUncUgKiFAE5f7zV3egb
/y4XI1eJwwAkczNX+Bd1ZW/x/xMxVB/r3Fc2YpyRuHqPkZUT6/5FRIdxx8HYDWKzfTST4DkJuhCh
xDD9Id3f/pkhSc66H8+eE5RUMQIMnxG3JH06FRB5X1asT3CjE/QUoQUCcSFubqeBkKek6/SuHhiR
K2F6atEC430D96ZdfHEdo3SqoADhbgvYLgVDc4AEisaPWNed1k3OU4Favg7PHnQb4BWeonHyvkV+
kIhyAOKWkMqlu8LI8d/m5h/2zRLUCr7YV90WegnDbAq+0BDWu3kDu7pi6ofht4EFzB//6Vt9h/e2
6LfDNfchAzj8mWuVa/xyT3CwuZrOnBgqW5icK+I49K58qgbyyQ1tIZIkLzLDFyRsbtcj5h2OWini
4IqAMszc1BmIjf+A/X8Qswyjeyq21UacyweHP1M1/ehTwSS4W5kl9j535JOgG1bv32qM6aPNDHOV
XKBr0L1S+r+47mL7vgcLmS0dW7KzJYRet9z/BWbv782o3cb09eeM+Od3KYZYCHrRYS9/EK99ozIG
idxJRVOmvBEZK/0+5aZukgV8VtqAjbadyprAZY67XRckMEP1Vozmn6oJ1wbM1enJsk7SVhl8vsR6
Gb9YT5not1/maQUpfqcTNH7Y7wZb8/jaonwRG/MB0PIhZE31gfCNxD6wHMisbB60FM0KlxdfzSer
n+Vb4YRlMZDPzSN4lP/Ybq638zTu62nJk1eRzuYNcLVeaOLRpr/wauNCSzouVO29/i0FHDahEAil
ZP1Ha3O/DWbZJhspc0HTIhNZFASnf83w47Aduf10izWHhkOQfFTyZo57H21nFwzkFjwMJqZ8RtVY
Ul/z+6Mb/L1UgvTigvT+LhPK6niB0rnTmEo1YWZ0T886yZ8JI2z0IHnjKc25E0wjaVA1go9EAVFF
lsmyrduQ2ph44vlnCx5JZUHatTQWExtRPgo12gsYMi7vUXDDKi5Ur9YE+CwsoKdXvmVipITwftAW
z4ml4ST7/Ymyec775Ki8UgwjgUsdwDUJlGXDj42GqxxE3zH26evY1F0P1yYMDKkz9cUN5LfoyAwF
MEAQ919ZvrFqISmD33qNTWKsE0drh1W8FOwBxOL1jdwHRaX+GyhIldtsoeTSdufFXBdhTm/zqpFe
vntXQlLgvlJN+dweMnUIpWr9UiiUxNR7/defWtmTHWfXCz0tllx+Orx3SRd5jIEC8msaCckGjhff
hXxk7aNzytczCuAsteoGapcU7ItOYY/15Jb2mYvxcFEzSnn9tTuMhl7exPvc2+2rDguKla0jsD+B
EMvJ+psQPlBlYnKZY1dquq/mnxSzo5jrWP22mlL/ixXFVTpzkRvPEAmkqUAR7cIXZs0Glrq8LdL9
Hq63BcxAbvacFhQk4au0IkjCSkoPltywkZhWr9nlEr78F+vR8ntd45+ODs8L57SPjhdxMA+p9rCF
OJWrP0grzVDAbvJIFs1PS4ncEoRen9EGjFHdTS04TYwjkvHIBP2pLk7JUZZGlcfKieYi/ihPetg3
yfysx+spWqUvOOfhG/9POhNiiN7d4wsDXfXqATEDEcYFB2biNFzmQk1jAkmfRKnbLE58Jn5QEqsx
+6iQp/AUWQXgW+P6gOJnyK9yhbEjlQ0/75P37SSdw5n4hbxWt2YKW6JiV5pnMjyICloVKceANB7e
VPDtIvvet9Aow/OUCLtJwCU9rAelrH04e9vv7jcrhqfBje+HGSk9OI8ggqve3kCqEkxhAjviqn3L
DzKv464v83V78Jpgnlaaexw6/a1DzTDUDoqszNKn6ZYRSzBl5nv6VqnvCCfYDlyu8/0D0jNfSeuM
/F+T+yQnOQr/mqWegxDPcY4P5Cl82jw2IKqhZfrhQVMq6xtrKHxZV28Bkqs1qzuPH1zudpmFW7XS
plmfrLb2rxPqT2r5qM9V6D5qD6po6OhvIU9Y9C/SUl3hGmcVHR0QRM52Hwv1m4VwAhe2ZYab/Qsa
QsXQ3ujklRHjXR8IOntojqxFU51qRVos1dVVkJ0+2srVrnfJZ3PS50RzMeCTa+WIpiRr0z/Wa6AP
VVel5rfjtbisaDqA1DbEK8Wn9LND1j+5X3+YecM0b2yVZHxAaf/cayq2AoItd1PsKobxQFAPt2Gu
QD8AgNOPXnp7R4p08OLR9OH7Vz5OQE7oT8gxL3xJ0tM4XcWyp5gRH3QaX3Ap+T705BKP+qjxOaP+
39Mt0EIV9et+aJj2jOCrVbspr2zcchGMNjMZWhZZVbuPfORrzRR0RzuEVsNElNBQHFNZ5ssIjzvJ
HMC1Mh0NJqRNLX6JMUudMFPqhj3GhgPDWMS9LEG39PHwWahPVkBrowu4n7fNE2UK6qwcjxEYF5dT
Tj+iGuA2S/p2We3+Jbzy1Z1av7F1fdktRTTRDx5GTz5N8BxKrYE89aifbrlTl3zVRne4JgwAzRQh
koTIxfdIkQNM3wPUCT1Dda7kZGDVkspztxACZhSZ8tCm6+btoVv3iFEHQnSQEmVG9zqPEmyo2QjV
Tnn/QBW5TZJUzrfVNCaRI1yqWp4gCqxIXqwa4zzXnHAJ3Y7KUvlEwr9SW+fKR0TWHwtnII2H3oRb
AWddNtK97zY/KCrjgTmkXEhlOjowYP/bey+IrOoe3N6wAKs0lymcmyWcDiGKUOqak44E42pVvo1u
QJSGEnSKa2OcnoFIydBdiwllimX2huSqAjsmUQoHISe4+BrXSJnxT55zDjNyRGAs7vQdDGrwFWlG
Pi+g2hYf4c1EyubvhwU5nAfE/cJ/XKICB03fPW5e/EjU+m8g+J3qsPD39DMVEKzelDcctjmf1Ycg
DfoJi8jU0GYxu6cNVxUiNGNaVApnweLpF06W02e06GwQ0eqnAHqH24rWNK2nCe3wzZvwknMKK5Uz
ikuE0Gdw7ELi8lygb4gJfTGZL//S/mdC/ypZxYWHn6UI8y9aTh32lSrH4pfXWGvRptFNlsfWWlQa
iszoVhyk1l+/i6ZuJxjSZli+gC1joY7mq1YcXlJfVEYNxcl032Z3VtNzuV8TTnxhF4ZQHzLRS8+X
pzVlgaQYlpA2dYKVQma8zd2riBH/QQE5T404IxzdwmqHq9VkWGjE7RSaEG5NTCOTQfogDTxEu8bQ
+AMi2amFGJXFQ5kqEFBs2HcBbclsueM5G6zyjU1gkpjSVD6EDw/7TLCSP9tOScCpyGzO3yv7G/5a
TMts8WAstFuGcqdZkldSfv8t7znbDBkRsAvXiEuK+BAUlGaDl/O8is8tGBbkpchP7L0VKZmGX7Ag
CLCTU0H13kwh/0P9tqS1OlR/akyDoy6ZxOjW/z9JzsJMq90Fn+QGi84JyZDsNVRALgy1yPTQUUZ+
ZPkLSjcJumRtStNUxGR3MD1jQXCmlvpwJYXYHmsP6XtCXyjgOUngZsuZgtqnKk16VAcWIBw1BBJt
vBjQd9CxTMH6gb9diV3CrfzhM4h1rPH6BT1gUAPulkkhMjKFly0wvp+OTGU7z6RFxADMKQ2eZnEp
BwAss0mGqHe0r9sk5VHqWyu0nVbkPtkFjOwQpE/faUvOB6TLdu+pYBvLLLnO/o2mthO8WpdT4XjB
HZYrnR4M7BBzyO3X/vfyzefMKv1SCUFClvMXVOEwSkRukE8MtUZsmX6R89iBHQxWOhevtgkU1BY8
cahw30MnnmRmcAa6IUo+/gwiGQQkRx8DIqwHYmylwtIBYGpiRmJ9ASxmmvb6z8kNWH19r9qmQies
UtgVWU2ykbwDbbEkIEgIoRaxs7yPlWdcOMHGvX/VH8IHqp4hzgXhtpcnOSh89RmknjRRgq9nKTro
xgE/CWPOkd75uAqUgEgkOBFf+PWMgb0IU2MRTehKCM0mxg7XzQo0LzfxCdPiRGjcvq/bbm5PyvSF
Pq6sHgbklLpIO30FprNVhXfZWgOj97Fpa2mSayArhHF1x36cSIMtnJI+pqJTMeGhzn1DfZPxiHRm
wgdO9uixFJY9U8ZqsmyuLRG7G2bQqYS9vSMRREsJ4uQsp/W5LWRCvz2QKE8H/yd1Yk3UoXwmCBEf
8mGXlNF1YlOZNax6mZsIN1F2tJ+qKeTm6G+Qlt5b/Te0tqipQm8aiXuyGmMY7ZlIZGR8DK+nzg8Y
Zg4AAfTr0y97ZfhSOkdMrrAxoiSDlj9yHAJQ9H41V8CFpkuFfqyC4kHZkhp9qL9ET/EWHggSYSIX
JWcuEvW/CFRdsauUjuLiuhNFj1wR5NQxwPXEZ1YI9rrcNK0c5tUhaDfnhise2x66CV7OaJWJKrQ3
h6WcQVA5sReNaV4S9HqoQXvvMOCMCnNUt8Hc5Gx4eyuyQkgrFHhKDrUbFxirxZoad2qFJ/z0K8me
55w6LU+Ir82LWXN8PKwZRah8OWtMtYe+4JZ+yayq10hMYi89IJkjy5m6OQ6br0LwnyjgKvcsbnb7
3BhDQdeDNzyxDLQtLZkkyYcS6nzkhbzNmTtz/2qbZtNhzPBEalMLGnhXRkO7BU1QJoAc7+5PRxrj
/p/LlprB2a7LB1ziwP5A3H0b+2SdprvYDm9OOlx6iIBYVrTvN8vX1QUxGIpN0YcCGlhrYxdKdcyv
5HPSiXDBN3gUBwH7uUXoouQ7kbjyMm+71p1YT/fScAtQpk5IxBl1OmyaDb6on4Y/vmaN66pbRhWi
eNqbK2nXLQuuzSDcXYujLxA7S4TzhLb5qJ9uYbK/bhexPFyLr17LNbQkOFqllLXNgy/styrmH7JG
ZjF8mvOHTzQbGD1+gBWqwbl18fJpSAeHm+NleOosNfRmuKXEXx7GcmJ40qekEUBTZ1bXLaO+qJUR
btdoO+T+IVOF6V+DeXRFQ2aJfX7eIxL+hYrloMA5ckE4BXtODZR3P3BXNdu4I31nBhzBmNGPd8wJ
69lz8Wsnc9tLfz5WxBOPDxTvRbBZdqdHtkwedhZOwPfg9Sr1ceHlYg/rJ1XlB+0FsR1SGE74U2ng
enj7FgUO9X9Rza0A3mxToUqzaZukp33KEt/b6RjAPzOiAFwuY4y/GiKwXLxwQ4CZQgOh1pzZ9jzW
w8X05dnz53bvCJmcusd/w0/BYhN+YxJj104IfGqhLw9DKiwb4EqEHYCcGT1HtHH4KO+R4i2516UQ
g8Zuyqou9d67crQ7hfwdY6cXKjqz4IuB29mcYUCK5wyUCziFh9PYT49TCU/emwv68ho4nhJYpjBB
VLIO28v8cW8HczZchWK2Kz20jCVVN77yrSYHaafk0Cu+YM1xgda+l2RxhOW07S2c47a20+5bsK6n
X8Fj4Q2Bcr6cYHA1apheO5YDNHSCPhaB2lsGQmnKJuQSWwgQBCUFiiy5ImjLHDi25zt5Qclud84x
RuAIqiyobMuJU5KUs4HYHchLUwzbU3bXEr7QYYN4dNuRurotK7hVg7KcSuz4vVWft8DjvKa5z8Tp
sPy5K/ztv9PoYFBoJW+cJbuNUYIOOpoGxNeSJdzBQv2NJHBvsxEKO8ar+HYop3WOqDz7i657o0Mw
vqMj2O5sv6ePSFBjbNu+/ELDdoJpl6sYuhZo6D+5AKcDMEQ8uZZl+gzUKkxErXnKuA23PTlZ/GkY
NL+XNuASDD7lRY0tR8scK9GENz/laHhB0O7dKP8kE5GSCOqVzlOIknC1HYRvxj1zUgMM0ouc4aE9
1YfsWzAzjQ53NPfwze3JofwnVcMl8l7afC67fkyU19XSOUYNiuiVVQIyjqhuMQf0n3H8LqFOra3u
dlsznkctNc87l4CFVLpwZag9hl98CvTUXhkL+mo5zhhHAP0DmBtRD0e8J9mAdcKlKZXOKHx6LAj0
f5M2nr/uuZUei4gehS3Fl79pK0XopN9ApioMe+xgmlvLUHz96445cxsRRTX4lfZi3RZ+pXAhpMaf
T6rreFoYsV1Hepeji/b+5G2lvWdPqKbAD7vl0JbzUgxLxEfClS5vMgsT8/qkIiajJPcUaZCgc8N9
AqVB5UughZaO3qrblQK1vlqrozzSwDDw/oqRg2teK7m8Xn2BylrqJQR4wW2g/NzVZHFdjM0j+Tqt
UkUyC/hRb68rOO97ZWIppbEJGcCJuMRSbAnIV7xwP1LAEMkn0biDYsy9aa57MKBsqetY2zweY9eE
exFgAlBS6zzwVDwpompI4Dr/MEMpoWfnaOKwJZu2DN2DWglGgaV7+5b4LKOUtJj96379WRPmW+sz
707qF31oFbVAhGqrRCs1teSe0fw/YCYp6v0Pys3qPHUbfzd1dnZdCwpnAatVadBVyVhifXr/Xs9M
OIeOzXq5bHI+DOhl75m4JReLggIqpEKs/+iUy88rg7vyH/uXXyBEKpc59f1OjiJRHjeF1HIiPRpb
+p5zLMH1ROFN1/8lWohQ+RLP+Rvin02+UiZgv7Gb5opjNrbtYnm7v5CUxlPEkI0nlrBikYy2rY6X
+C9Y3L4HHI3E0eZ0P9Br8n7tTo7cX/0AluVd33ki8FbGtKVmIjhyFFrloZYdqXcsJs+CBdxoHYMA
IDb2Th7n75eh6jTTbpb4HSBYHNObE29rjz5HvdscT1pDr8yIBs+GUw/FHRlTs0rL6mSMBDNdMIh6
IE2/4DHvzqyDEnjPpHYrnN/LvsXJ3BkIeDMYG2bdy7CClJh+kcV7bAPRGrnIQfzi0Nn0jQ7bGaZr
m/4Rtj/aU/SYJwL54uE1bCSX/LTH/ungQgmRM1aoF7fVGh0H/j3rv/Vf8wIwlonZzxIwl1Iui310
g2/rEMOjtVheTVCqGPYg7g3+IHkSplnVrzCtRF8HVn5LOxuMcg+SvhDEV6HsLg/gEuhoN5GwXqUz
bZ4sGT00LeYL+PtcxR2+GYWaigDEltjNahMVe4l3CiP0uml21/QErlcVyVsiSBR2VQDEJvWpusTE
ziq+HTbNDD7SR0SpzlCBeAolwHM6WkZHf933WGas/1jO+VFuUbHXeeX2y1j7D6c9TvZuZAD5P5Nz
dkPRDPyv3AwfZ1cOskMKJ1yAdapWOsgdJh3HVNc57MlFs1Gk0rlyns9gur2lPKKr+OekO50xV6bo
g+0RlW5V0ITuStZ7eca3eOZtsXm7k5/lawR2VKFkOx/h7f+RrDYL0LvKGIhbarIoAXIvofeFiRmf
eHkPQtJrNww3bzcOVdWYWzZeWfPLxi1IwHnKfaZx4BJcrVolJfZzdcgXIpRpTgNxrFvo2CPbFnCw
fNXjkBMZWdRQj93tlxckuXKsMa8Sds1fPwaSsZldBo0TbIKCNAs5s1vnqC+cEuoK4D9XT3QV9Hm1
03aar+TNKQfoloE1XDe6ifCdCeCZDrqIX81Uybbq9iwgtHQr86BAYi89j2Oa7wlqDoId4L2GN/Cj
Qj6atwfDXNGF5Tw7eJv+IJeEbDwH/4f3cUm2TCmPV+MapiMIdJNbkqsR4qhbjqf1rH6yoY26o8D2
nzucNx0QQSO48gIqn9kMTKm4aBZLuHtFC8IWQOEEa+yUQNNY9oYQiCz6VrehiwtubvpoyC7BbZr9
4xPT5D0FQei2vfyrKdNh33dUGO4O8OsWX+yb/N30xCmlYqIUsWWcC/rO3X3A3noVS+NGIoZ/JFJJ
TuiYDVbRf3AGiFHPUAFIn81sDxtHt7qvr45p2prGzg8sleyYVvaPU9IJ4LQu36RjUxaMlVRqjm4t
fP1+GSpW3TcLig+6TEo5V7LN+p+KIauvYvYxrikf26m0Z7eq4TecyI1WXqL9tx75r3tEYeaUquft
Z9SC72C/6v2YvrpwT2fgecPlrZuaru66Vn1hYXPjdzRF+TinqCoOXLkKEFXRcC3MgE1x0iNOy13p
kPHkgRuSvHtR+q3Peoo92RDQ2II0AdqygURyj8y4neE0paZiGFeilvd2Ohd3n5XvQwcfLgEMkQ6l
cAA3ArR3kUTFmr8l+1vpoKfWQTG/OoXQY2wRhX2sDCUkCntEfD2Ab8yRGrEe2n33f5m14hRB0Rdf
D3IFwAFW5FRinokK82Wl5wq5Nhr2AUvM+36634Y9iv9Z56eBQvCpGK0hXbKle+kmXiTsKpNkJldI
uFkf1sSPj+BVyvQl0UTeuNEyrzsJj8fY5BqrKPt64+gQSWmh0cNyHpNkVLKYwlhBIKauldN89SjI
BMUE4v6F9rchdOgumQOllwsqTDq/+/iDc+2bcTbxMAGZ82nWSUSAWiI7DROMx76b6hn4gKfKPIkw
AXiMB+QzX+xqQWDRZ3a3KCJlKtNS/W4R/cJufyQLnfcb/jWtt+nlTuRP0JURgsj9/oPOdZUFnu6s
JhweGCs+LV+YIh61bdvMqklj9H75kwN8USpqNtd35OWax0UcscspGd5e2kDLdhtA2BM5oDY0KyFU
gQ4NoCP7FhnQ+l9XKjwjARQO1an24sAGY3Enw5zZUDRTsQEhS61ldEtk2K5GdNC6GZbHCB7kByPz
2CUMXeYD6ERaP3IkfhiHjNJTKGkQQm4MYijaxKrP0Y0bfS+Sfjij6KTmgIFJsb2anhyxlzVGFeJ3
1ssGu8AGQXL3NaknI15dzLSVVOE+tlx8fKXikAsPHJZ1xxd8BH425fvd0s0OK2PD0EZw+w7SpF8r
QOwbmySgZ4+VDNum/Plw/cvff/eZ9aaw86SJ0Cov/g1Sv14IfydrBwfcE4dJZcBKbtsuoQYvTRz/
4thTsfK0JjZb59kTK8WBvLmPooczrUinmGk+D+NW1wTJy89p3e5If8b4oMkPIWd2bVIFtZ3e354u
iS3VoRLdeop7m253gMldNZcnMGkLyf6YMdRAfMtk61tONaAr1+LsIt9CMar0ElH3rqiiIhTWo7V5
gSNVlehgfpMNjMI4ynG/NrjUeT7UtV0K+r3svr3OLdbPfL+G5q6vOzsIi2zzC9ra1ScSd8QoZ9Xz
Z2GSDJhTc4uIif/TImIY33DS1uQQQIXnqTJihhhc2muv71PRgpZWEEkcxRPFzoGd0ErUs5OuXEdE
pMMseMfh52iwXSMfbnF/cO/TKG5/x6MA0dnBDVAWoI2iuMVY2qYjbWgsTsHYm++QrUinpkotuQSY
wBmmeS4wL2nVOhQ0pkMTSKdEekTxAIaLeq2yTF1TmxmZE9IogV9Q2vYekO8xKsFLSzqwpo2fiUZ7
GyIKPBEUkcMhOwPv0LKW9RZF3KKoj5SEI8JmopbV2zzkoUDh0FjX5ouZdP4vdwLArR+dyXforRD4
BL+/XxvXo84VNt6NIdjmDX3wsylxasA4q1Ev9fVytpmx6YIR+ZkVDGcf1WkeLJp7POILScsuAxMi
4fJCMGExHXxMU2hX7XkbVJc9kND3cOP4YLp8MhJPE9n7F4lPphRDpaHpccEtmAFJNZVUb11Bs8bm
umQ5gD/Tgsw3qlS+PE9dHCRBIwqadzMB68bMXaSJkQoWpfBRFoKsfZ3C0NyqYG8nqVoOye78wkk3
xGkxsqdHz87TbcEFA/3VACSTs5PxgoZZdbGow2idoze2TLEyQ19gUOXeN4BHh9Ij21vf2Db+nT0E
yri4gcYpmzxCicCBD2Uf3oeW6U4d4juYuMJecZCls0v27aA+55InuIpJYrvtQmpXYHu/vhpgMRHt
N6dnMrD2JjJmbQ5N/aGGN4iGGNaUvbav68mmGmn3R3mRtcAuqq+P5xs/crX07xZubpGjyXetg/+4
JKCmBpKeLVdvbJyIwHEz7SUFkV4+omepfKXB7O0ULQY8d+0eEMbNqHULgoMQHTblV8uLrAlv7smw
jWGzz3CqT7VRX9fF8adijRivVZEewhkpWtFVTyeo+/hw467hutb6Zr/76r/qWMrPIYhM0kBaB5Nd
q/vjrdmEkgeoTuUd/MpXbMpQXQRgEEnA3VKOQrB0iXHxBxg/LAqOdLhszwEs1QFE2NukYJ1m5JOm
l87xr2RljkILvCOdp7fR6mA/00kz09UvNCuKTMopTB55QT9qD7gquuiZHVm0Bf1sgBTcaNuhp+wz
zNLWal6Stv2bUYBMl3k+B4qJDSQWXRqREi5ykCPSxQwonwNFFg+jEh4qxRX5XhxMf2eM+SgAQdz3
2+OcA907AbT6pxl+AZ4HOQn106dg60wCO1q83/aDkRW100ke3YoqhG5cpy6T51bJOze19E5TvECm
p2j9mzASZhJqZvyZku/jqayPSPsze7tCAOopEcAz0Jq2jHXNNXIBb0ZAcZgHpvzDn97LfqvAkTjF
NctGx4T/p7qQfB8koEaziQk3nYEJr2RzHTvRabuMtpJZH7QTa2QTwHucHksJXdePXc94jjSf26bR
OtaOcM7LBX3Iwd5AHw99j4ZNxHMbHWdR1UzX2j8kH7BZZuqxpl8F/Q9ah2LutK7GUp4HAM0qRh9u
znmEbLi9k8zzsKaRyPOUb7Lb351xEw7ku3VvPRf7WHxkiPtOwV8xBKWoQLUoLq4eY1TTlNesAsiD
+4GgotD6JmI41uA7CYQPxO7oWbja/omxYPJBHQJdAhDx2G9ptQ9Jqh2PTsyYqzc6HzuU4xX4ALSP
/xi1Z7WoGvrRUMZuaf8eGb+uTVNUtfZlaJzv43EFHTnguiKY1nge4a7dkQPbSYHYVaa/nCgmmZFd
VvTOSzR+G9gJZsk1ccoKz5ScTkeO8Cw8jH994kGDV4y82jxsRtptaSSvlOlrI4gZg6hFfa+VX8XG
wUN4k11oqUAueChNNqgAMkaEoh2vO3yPW/NIIlgcDKD3q5B02b1zdIuUdrGUm+f3tRJuTDf4KyTB
QXTNWpOs9CWbbCjjDHgn0u39hQ8ZNJRiAX4msx+aCy0ueOLKAZf9TqQ+rj4P31khuSXlhfRnflwX
RDXhsi7qiYveGaetUKMULjALmV24spdOCcaf6ryQqDCa3FQ2A4kXq0jpou6zW1urDyjzHAiqGJHz
qcQ1UzwL2nvR/lestlNV6eFwgq3XYg/KSoXVNtkRtwOQYRc1P9cKCChnM1epHAxAjotXVWagiUoc
JHEYAQJ9HAZLXIm2w6IiluILmC4HpZN7/3oR1Hpe4kRfIkjObT+UsnPbeE+N8rnjCSSXp7TSzKQM
Ne1hzadh1jIrS4H6F5Ud2NnLM0sS2VCC/caYTQoFKd5YvodIWeASt+lBmjUWzu/IYUbFpD0qD0V2
U15AzxRr1jCxURgx6sTzqnCCngqefn7/IfrneEXciUCbD6c9jz5mrd0Na8fglmbeosvxcJIQgnro
/EvhWaKVnGAenJ09zfgUxCNo4BY/RjYHDAqV4LR2DF9zPz5vpw0mOTed5NhDoHleTc7mFGBPViiZ
SbMsIoll1W+vdIRYPnQG8w3XhtB4Cd5WsSwo8LyRTITnkn/i3HMCW8AWgdlC0w7CHFLq7XTxALMO
/5qdhgkWkpA9uaPm15yy1RwiYSC6ie3MLsUsXt04WjT7vQuK7B06syo0vF0RgKUQrriXslSeKSgw
MHrtE3AGv3W7qzX/j/gY9Hyrq1eGn49wCQO5i9zbggAvdjdTb/FHKWQy3pDPTiT/dvegQHCemGga
vprnexGp5qAesgP5Ss+9N4cT7MJhauorscP4EPOK1aKNvLYq8o0J+tV+zCLq6O47wpjMBf3RbRb5
G3nFtBGhgtvb6JZqaIQIIGUX8j0k+bdokBfCFu8XMAVDVP2MIZys6+fnCHLb8s4MKCmkhf57YCRX
GAQr4ivWIUAQ0sygtJw3jGrGavqyOnoPEyI+4zHvTGFtSbJs1w+DAdfjm4pJJ9nyod0TajzvFnS5
Eydy0DbxD89/PucuUv+oDMLI2jP9pN79+uBoCB+14oyu6mNo+UkEo+gR8sMcMSF+eH8+ev8PN9Lm
0Vv8rDRoUksJ+1iwOx+l6c7IYmuXBl7RZw/IQShuiR3EpQ4/VPChXtPs9F4YcNj0HNCZGrl+Ruw6
CDfLf2Vdydgi651VODJ3iNI4V+ZdMYvVjz4xULU1S4KfxUNTdlsYaNnOBZNbw92348Qhpcy2LHti
TK5raMkXwWEQBhiJ9/2F3hHoR0i0k74ew3Ub8x+bp6pCLsvqYBkHipv9uz4mYJNoZ46MBFCfPIBS
rfRkIS4tGSOuGLI8slCakHAxzll8+UhOPsou+zw/RbGKvGe38fFxWa39GJjIbeLouZ69uZQkmc0I
FYAyGcHxJpObq53dRGLvabxeh+kfFO5/p7b/EVQyADb46Zajvw+ri7vY8f4cGS36ykDVDZq183F6
6yyC7BQWD++Wre0KZB1wWP94KAT+VY9gysAo+mHFvdpG9A4h9eUBSEeTT0eXU8MCEmrZLXphJaaO
X5wxBSDDo47opbqElNwxKgnYYFK9z7MFZDZ7jXgnKgj1xRehGmsbQdVGJuKGhznlBhqEEmchpSH3
s5xbDOPOa+0zQ+kH06N96GCNoc2g0QbLE3BgUYbsgTp7sfkDW43wMNfmMPhLv286QVHfhojLfWnu
nRBzojk8foEK0GwE01YfNTI+JyitEWcifF7e9FsDyLZGUiZKfCUgXfBnwxN+g1TATKjmi8Qie08t
sf2SwnZwl2qXrEmbeOa0ytUH8JDvU0qR4MfYgVsL2LFsfYoFWEaGKo4n32a1mTW9QbV4d+QYYw7f
ztG2p0h6u/p7cWlp8g9GrM3uEvrafoVymIGsHzH3vCZSfY4ncmzwf8BCx5CttDQu9qRZmMYxGyKX
bmlTKaBp9nRBgXblHHHG4bDMq4Nek+zOSBgqZ8kDjAYk4wsYsWDB8b9XEZZSwbjrMWT0aPCKpNW4
UptBMCsXboCvxEGLYw+isFUxnnc8Mx6NVWcCQ8ceOej3FvKcQ10EK7uBImSZveE1WasT2b126F28
dYcoKLC8ACwCiUEtlUrMpvphf51KFEZzju/KLubTl7qQYCB/hWjunb1r4zf0JTo5K9aZVC1T0aX+
+WTc+MT9eZkRL1pKI32deFgPI8VpY8B6I6IRP6JFwQVNsGsPE+QGZ8PmrsGUCC+pu43mj6hbN3XX
pijGBnQHrNAV8H74OJz5owlw/oMV9AeU9RxBZrKPRW7+g2jJOUKS7QZ3IbBnZ6UKgMFMjy4KexPD
Yla/YLO97nl5uC5wz0ux1mJWgDGAu7k+fUv6Nhwv2yy3IdqNz4MV3jvzbrzqC9bA8N+CAiLVOwa0
NkM1Kovw7r0hWuR4LPlCS7QS1SGdqRe7c9RU8HV8Ha1OqSnaaAHrvxhPCa/oj0HPBDjginrK8ALO
U0GuGeOwARBw1hBOZULGetGfPPaSYVmb/1MCheGR9RhHPjahzzoIOZ78mC9zzW70ZFz6oFYnY5Wx
hQA00S7ZSY/nX0ueMEDKYDGf93MbJANjf5RcQr+VX6NUt0MlamIzFM6OFyJF22nJJ5p5GyhLp7lD
PKqAsAoLyfsdD9yClRmknVCDmd9iw8xe5WowNoJDOQ45BjONrrPqePuA99QJNw0XhPP9uPzRsCSb
LN8HOHd6G6ROM6R0yKg0LD5ExikdhuPgHQPJS4x49VEo/mQYGDcRV/O1Cwe4FtzyWTW7Wu0LAz34
22DtY8X4AmKZN9jPms7syY0/3QfqcxXsp6negDnM6+CkhGuYQoeqo2nLCa2O3BRatkN1H41JOYmH
d4tMnvMHD7cHbb1BHYVI0vubjvy9SXcAHvn/pWhd8/JmeJBnn5WA1ZmhDQpgrx3v29futGRL62sy
AT9nf3bLUxZIavoZVEHWp7/zcsiW895qrvJY3isC4HpOA/+HKwvFxBSWJ4KqMqFoWdgWq4+EmXoa
EZOihyWin7Ue1CtCN5XdLa8tRjQ1NBHU5XySf7Bqw9n7zaFCf2VP3Z1zLP5sM8tzwvITN7pxdT8n
XmRpLisGSF/vyPg/x8va78covzzfkyySpQC3ag7WUhbvrHhdS4Ji70CRic2gfS7O6qgrt+Euu5Nd
Td7qHJpA6PsFbbE7kbmiRwStnGKYdojpKmLSXtgLwz0MrVNGxIdZDMfKRs5c+2yOuqPgsEid5HQd
RnJvOUPZOp/dAPINg+NgbBSFTRi1vqufil67eMyL+u88kUu2gqoDonsPph785DjiWqJjLxQS5NWr
aLomoBgwZGfiq8qwYI5WcMKJbU1BhfQckAkmzbLpnQMlfc81F3RP2ZoFXNuyXMhaubUru/BeuqBV
d160bgvXUh4gFKJ3Wbf5Qv40eVXgH9/u9jaPQK0fUYDxOrJBbdFUn0M2ASVOROLfUphmuDz5FGqk
XOjvj11Te1nLKyFCWm34njm4FBBTZPldung1wAEr8KmDlGjNwWc7b4kNJEDknu5b37AyymoYdodE
IkVoHBKS1B6Z1TtjSJhgfE2UGUcwLHjFDoSO2U/z5/GuuFkvOYRfZjv3SFqGQIxtT8jJKvAibXq1
GHhRzlbBzRQblvwxaeCZ/zz75sd3WgMJC2R2gZIttAUUxSXm2GFX4b2EPPhdxcSH5nfKyvGUo7IX
+YQRIxJqVD3WFgnmEoJvMQTOTYnZT2d7g8Pd0r68pK0w7qiY0qdpDa2rZtNbvQFBfQp9deb9aNlk
ivXuuJ3rSEaxDQWsv5hXIqrPxXzRkfqpQx028fqtQajdr5h+q/7G20DX2ExOAm3eMIvrmRG82c9/
6D9ewzGRyg77+IhssSfRO7Pvkf0IFttZ1R2JYIXA6+Wx5cgSZqJ0LHiOTE7p9mWEsjV8ABQA0ysN
WdCWtvol3rWU+9gZPaUn24uxLFoyDbbfeZOyPYTMd30CwnHBoWKWwSbUDMvOxECsdVOfja1XzOzu
7Q5z064o3TNkzScDwHFTewJLTzXaibFqql6zFFSrNKoBuZVLTzLwIgSeg5Cbk8Gh56MdIAYJmnkM
/62/tddxyFv2n9k9Y+MCuk7khp6BpaFgj6ZzJwFgh7HseYeKl8JuHs1C8CdgS+VXGypQCf582oFM
l/oXpxuDTZX/muJAla2FmQYvzkGPNLtf/+XiarnfwZn0ss6/SfB5AEqfVQ5cXPebKQmCV0t8d+th
KGpB0/lymbboSpTtxGGfOle5zHXECJiCreVPTsmDTouOmTGNRH68iYCFarZUcovpNKTyblJDdeRl
ttDT5d5OGXWSAdaL9qwwo4wo2/DV6I+5NXCyQM2/gEyoD1/HMiyip1/+zveWPYeCE+Li+FX9YwH4
kKRmBsPacK2O5gTcui7u/jJ0az2lN2aTM2uz/AVPeshPGwmeJhiEva/mzk2YhIn4xUBfyPuu4P0D
6o9vhISTsY8xie+Ev5sRcEMU8RE2AcHzyG+e/nJgVl1vAQ1TfacJbHyJJxExzU7bFWMLET6E/1Ye
Sp+IlU6LS7jTFkDQbuUAQec9y+1ZnZeUy9H5utjvjLFW06JqDSrPmTWLjY+9JCJlQ69ILAMm51st
ysu0IfeIefcktS2hvtEKu3oO7S8+MopIqytYbACnU9g+/p/gUZP6rYhMuRoRrdXkWg8lMXV3zHmy
/xnAGeDg4h9wNjSWNaLmrwIUjIICR/nUbkUpIIS/VVBQvF25KMw0QwOVBWrkWcBkildhIzD5ZUPn
5rpUFH/Gcpj5fosY6x0poPcabrdmgAVJazSNDdPoUCoDOmBvMCMlGb4z/bD1pAgPABhXhbWDTgcT
7cANuNyQfCS0qqv2rtTptbHQkB6N7cQqhGwh/nfzzCicJUTS7pDKhKRs1O25mFWNQDsKeF7y/pOR
SwE1HLuls30qWufT36vTlL1W6XPuAXrRTzPYneKArSE8Nj0FxwrXn7Dlj1k8EGi/GNqkbnBaRZcm
cIHSP3MJmC96Rp8JixgcrHWt0Wj4uUEUfbPP8yCNZyCNTG7Laol5/qQHOpcQX+gq397eM6OQyccN
4v4TKObF4DXug/9FeMgcs+sSG8nb4BrWNK+BMhPKE9Oky0I9nHODJBZjBTcZ4w4YQ96Pv2cdodn1
N0bI4M7a8815TSLjUA4KQfzpsARW1zga06v0M8jwrVTtLxAKaMvdkn1LgZreR/M1gmZM6dqw7Fv1
oZjHMCT8k7yYswIYfmIddCJZT/i2oCznnTjlqkt/IfxslnH2wbiw/j2S/9TFeMkklmILBnnuWRY8
X4oZ578kVwd89m5oyF1LqYeQO0XXgNO2rwq3XAZ7aP+pPjHSkQ/Xy34UU5CsH15kLKUXnU72O3JO
Q5JpA6SqW5sI+O2ViS9ABhFJbivfT5bx5yqnKNq5DEgKZuJ+Vjaqg1aAu5IS1g4Cs+augvmyjn+h
A0qdn++yFKw7g0p6+TbFlEDwxCioiZ2LLicgKQZVa8yKbEzl+LKAIoLb/tOdIDWFI3RMt41wTRnD
tRPppBP3c3GXJaLYyHlZtS8zPp4/NQke9qgJkt9PPONk37Pj85M81gwIbJDZxFS+LQaO/fxB6ujG
WqgSRdeB7hk3yjiauqW28bxmqptUZDtHgjHwyuVSTaVgCNHDXea6Vy1cVfkWEcqmstgO2T2a5mN1
tZGd88SIVbcfVxJ1nmk/9Jt8tRhbOvOVWxJnZg19sLc+8ntOrPIrBgHW7B7f5gRwb7gcOaZ5MCGa
1slseMUIIhAzkwig0eGZECy75ak5hxVyK/zdYmvykMkoAMR7LmmsoE9yYdGcEYp7sa7LLdjkCE0T
hgCBlpVLYDir+c07cEPkgUuvb+0aD8t3DpkaHHYdkBvSzJUUbh2D/4dmPUECY9IJHxYdXQc1kWzL
i1oSjXuPuTGeohxqZNUq8gFHjZWfF6Ru5RhjZNA/BA0o4DFOSVi4RZMz3fTIYYy+hKd5gR97YfKW
nd2kUvQrm8R2caeLaaFB7a+DKr6E65s8IMIP5+bpUbk4DtKNusPGqmXN3mpjH5QjEF2KKr6QEl80
uLYZKR2Lz6y50loM0IMeWsDQFZYvJp2BrWlyKQacOuQv7Z8E51oqone7rnm86CKrWnvM4HRKiy5q
ivjQswNuc2rSqwCjnxkyHFxV6CbdSLuWKbnF1ojnhv9uqCGayAgHNALj2V0/3py8OvpYS7UYA5vb
bxLtAUfsbnnIHk/Lupsx9YL9mBU2KbRz57ZNp8Thsv/fKDy49CAQu6igvFGT388ZGqbitf9VeWYh
VMZDelbSdO2Q03vXPk1DQy5I5YVwQlRFtJdaU6Z1kL8e42IJcHI7Z2NYCR7LFyjsxO9WUtUUoYgY
y6ge2SsGV7+yDpxNM52Gda/jkBw0ZBnh5ChXKUWvu65/S1dEkIQUKEiDbf/vJVvlooOaXuGBCZRG
V59HTsYP1C3xAPjQGeJDBA6JGY5zllkgkokUBGmoXNjaPa9hdFnm2T0F3veXN8fOAZ+ywL8m9sbu
UNN97pl5fxnj4NH2G36ZrTcmdRzB7v4l/TMS3sCfkg76vIoLf1ZK4E8agCn940CC9zQNOsy2ZFMO
7k7PT3X1fNYsvk1dCn1y+s/HAcJ20ZaCjyge8zCHeLJGrQBFJx12G6bVvjJq9DJkYS4+Dhpclgq/
OSCiRhbR75L3rD5/R7A91XeEeerVDNtKzwkPZK7RAfl8seYrdK1h0+kzr7iPxc4mN8g4Gv+CFBtv
aVSj84Xho0tBXDN0HiezvxcukKHCIvEV2GkLk6gMcd2Yfdbl1NnPVkFSW2CvqYdfbBA/4oRfM9if
cZwVkEglPOC/ZS8BrLhOESswM/jBDwLjB1cvaFJHDGUuSmivIk6d5xeiGvspf/HDMhL9t52NY7GZ
ZkS2yRaeOi62CB1ocS3AYu+J+iW1VRhbYYRQFbzPyVk+lBOA7bipn2LMQGRYrSTVZmyXIJ4Hp/oa
jzdpnANXn1UOlpfP8WNce+ycBOkFIYnXjKHeHstKPgByjsxZFUxhrUAQ6xS8QdV05i3u0QHuI1MK
l0b8ahJrkui+8I6R7aGGZcujAiy+s5PRrA7LlocmtU8UL24yPd7kBqjtwXsWhwitfsQXfalVKy1N
5rnzH1f1Vb3uQDdIhJrHPIvRHFRcF79dKwP45h8ieZUaHoqIb9V2Y7Dxj4UUeg4Rmi0jNFzJ+R/G
2oSWp6wKmE4mJ5MIvhmI/0aRCYMF8gDfiFL+i43WTvdkbO7Ytrsi476DRaggdKtoE9gdOkuHJjow
gbwF7LqCUIYcoceJPWJ1rswGDkmcriWg/9Wu53/A7j//1p1XrhbgGX3REjN2EBolzKn7Ns6eg2RR
TqWrZ6Uqiby+CpiadWB5bgxDamopqxVDOlarTrQh39MN8MQrgRZYdNuqBZAA855JhNUm2zxLjQlk
NKKMuCWSm7cb3KhZPKycf9tVKNqBaG3v7OOQHReFYVJ3N+yoxKIBVhVWJVFmIEyJ7RL6NaoOj9nH
bqN+DZ4TicURIWzjo4dbHSMGrCEJ3T7g7pVFwKHrN1q6dZvqgRdumlV/Ax8vdqwSsSk1tlLbvpC/
XmwQVOkqui5r9rgXEzHnN0P3PuNPFpwwR4UTuUq1zPC0ttS+G1pYg/Ji+kedhrPgw1aWRMxfJwz9
0zTnR1Br/lLShUNPRL8ZQiXJzWjnVSyRz0uZ904qp0uZMN4qf235+v7AJWwtAmZHVQsD4lI0N+1T
0plAZ4EgCs4E2Vnly090N05P55oVJ1DiylJeOyNp62J3JlbGfE9N2FufAhDNEOWPUSm8zsOMDF7K
tal+YMewgvxhaepQ+LzTD2XknLBkVPOAN8MM8uvLjZu78iQtDr+fJmOZtgmqIeJZOvj3OQcSTCjM
hk1HcT884XsjntZ+liAMo8Jl8FbF5OgAGUgmLvF0DfejyrjhBHVbBNuBHxXIDayO+UNR+vbYmtbU
k/OX4qS1umBQLQGfjTtqKqr2zDeL+BxJ5R2JeGkH4+ykz11Y8EpX2CkwRK06EQX5Gh66LNytbR0U
KEcMM7BL3z1MyQ4TraVV0uRpnFM0WkshWUze8kgq/AJccGH3q6eypC1upx4DNXWvcJ08FvW0TXuc
v51BuXRTOhwuiO8QPWYo9i1h02o6xmftQ9uFmUP4+0LTE5kKxXFfZsOUYwzvKiaNK70I9uLvP7z9
Fcv/UlybRUVcTG4KYFoUdrKLoLFMgT8qPC2N69Hn75b/0gt50MDrHgYD/Nh3bkKcvnyIIakKMCT9
XezOMd0MwdpaJAD1kUtT5lKToSjFsYLiBmCS4VlATy1qDV5nAdHzVkJQlfPDIdkzYzb7a7zzeddG
Pkpq0C+aaJ13E4OaMd1KHmImZPsGea6AxNwKP0qw0rrIkgfXdbTGArj1mc2jZaPHhsfCRT/uY7qL
j1DuWj96Va0t8el2fbhed/c94UNzVgSTdSWLwC5I12Z8Q6PQhDM7R5m1mHqQYOOUzRZ4nKB4UaXU
Mpr7mUQKNPdoFr9tTI174tyS9M+Px+VCI3CGZGuGQiepICMrOEDzc/5tl0CDix+XktJ8Olg9bicw
PcTfpVQEyt+5ebLj6hKyNrrTyXGes+asEI5yFtpJWOeACzSI7361pXkgcTUWC4w6yvS60ikKj2FK
DPNFUm1wC/prQwmJn6SFrLV6qoFrcOzXsW6qSErV+dgJqXckNQ6poeqd2NmxB+HZ3gEnV/zHwZXQ
ZG6VTAqWk9bfshYsE9twT2ObuelcJSG1xYjGtD2wDNvvolRFjqVufKr9eJ7pywPryoEyHhgDEbb8
852laD1JgcbOt1HVFuUsVVVzF58pDNhqBu8OcvDACGEuGKpgdOJNPpK1uq6EozEAi8FZ4bimOCDJ
5u0GI0laomUBlDSGcS2XmzTYa7S9y+ldXWNq2hGLrKnY0OJPkgxr7+V5yR7yuVS5dunanLlp7/Th
Si90sOpR7RX3KpAajR+xzWJQQDR6unlSsOU8R8q1U8XSCHqju7knKFMz+EQkRCczvtJkDz7aUZY5
G1g6PeJjdJ1xp0pW9PZvb93JBx6VUcoNnhCzvRX2g0JTdkHk/uZA3TdkbA6ZluNy6BWDNewx+eRV
kACyyH500vHPRqQLXLvap5tF+NnvPh9ujO6QrdntyXTOo2cCRnp9dqBABck6m/rNLwGVvl81lPEU
ueIkWfIMrFuxktbti6yz1GZ8RZubh4ucn46md12f0BfVEIBUZefM82gU5VWxVxhqVxqBQC4Ztrq4
f3Yvp7BQ9q0es5Wa6/4VuseEn8dUOdChZmL9Y+gM/GhriBZ4y/RyJyPqwvjIWVa63y9SW3oi9yC0
fOiPVe1kk1ciciJJLmbOVvfwalqUgOv+3b6S9O3YOEC/1d4JG0Hj/1ddQN5izS+oeRxZCD8RJKvI
9f+2oAM4EI1LK34PKFj+IY72444gX+vpO76w/wUzQJVTj8qQqkwVelz7ggeXLUfGDVmQJOAeElD5
dB16gmZMIoUPC8SEY61aojx15Dn4Q+u33QdKTCIPoXXodvS1xhMPh6EGLr0LZlYJLsXc6m1/dgWO
PFTiJrAfUIlNRVvbN4bJjAM6K2PL9Mr4LatQo3txWeZTq2592I43j3Km2iiMYp4IqK24Q6+0X6dr
zaAFkaGRDYp1SLGrulu3cUi1LGALGUqSbMf0zty8EGGda88xEsJGEgE5lOfaH+KKNqc5/H4yXtpZ
HzqoXOLJ8q467BnnquXoLpBZXKCJL9GKwmqGv9oY1lHCsztJyp8EzZqHzVieizlics3fePLcWjju
2vpGVARli1o8DZOFfPfm8tUJe00nImivc7bleSOWnjs4wsQ30JvjvlL8YdVx8cKI0XJA2NMKW2AK
p+Zju/2h9ByPNksNiliqZlzXYEIWVwLhRYDufo+T6f1Og3uPRFm9m2+kfsG2i6FSFGDAxdT0qAOS
rIWSzwGD8PgSM27jLLT5dgoOxPMokp9rMF48cvCzqaGh/PgVryXlsIkZ+87shbToL7JItqqEEUjb
G20zJERXEFF18TNZYq/CitHfiehjpvj7sjZomzdLoVYw/+hayVirDQpq3A0k0l/RBr1aydH826vB
Ok12AE51QwFr522Fk9f2IaZkMCu3jNs85VMsSF1sSHTgbQ1Dcr+eX+aR0UjzZjhpM7o5SKPWlIAd
gYStBVM9JrPoQfMbe03XCTifPJnILz7RE5zCwPbz3rdLU1pw8XDArFLJTUUliFdfUOdMN5MPhI8/
0O5uQJ+6Ztp9OS2sDXDFwR3gg9oNpTKtqHriu78z91pW8x2zmQQz414uVTPY8d7k6Qd85eh1w4Hn
j/md4vAhVBx6bpIC+f0kIUsWnMrs33wLoo+XzrzjqzQMIoQZKeguCdNvmUIXLXWd8b1A4k3resV8
WNJWUhgFuX5EbZrO6Mtgm6/58enmoDxY3Gbjqaj9i1I1E/zijhM6ikGOHbxRTm9a57w2ZzirHB4S
/hOEp57frfzLSOUhAG4cRkxu9lkdNRSAI9HIBNZ7RgCbkfjmLk2Bi89Gb/7v/YQKd6C4be4QgDEG
8MRE/zT6RbJXR30iUKkv2cJ7ilrs/oXLchhTRYAm8rFyv4X5dVSzHA5xwNRWRspfJJluVDXP8wx0
q6e+o6bM4ou6X95GuzpfkVPRPlFnVz9ljpVV1a7lXweF8PDHd5tcbH/IpK0cwSjdMbtLvnpcNDdn
ooHxAruvXLHNP1x2S/u93JDz20VL3jvV0/wOtSnaAoW9hXa399z06jg1vBb23Ycl7+Gy76crz1pm
CcK1faDw7NMcWymUMpuOdjZlDfiITFqZDMUJAQx499dZlREUC2rtmecVQJ/EIk6THSzzFQRyxQ1j
zVgCle5GEaLMfZ4oHkUSmRk5d66ojNSA0UpwFuF1jhZXAS5QZkPMCR7lIM1+6X88wozRNpNIE93A
mdlvDS5fUMya53+9Wo5db8sSIPw0pEkCv4ikhsl41RODel4Psac8e9EOeCEUYUYgUlDwVe3SfQFt
RSaDrwyfU7pU4iKnsXqRdpy4upPLZv+hqmRdkKma9X12FrregH3hC5bxtweGL9YF+ySOP5KcLK4S
7d6XXW8fEY5nr5iMFy99J43Q1WZB0u5fYuOERnugivqMoCBufwMOGEMzJUi154+3JR15s9EUfq9G
XeMnrTrl5Y10bhNR15MbSd7hl5pCHT21wDUorWNGYp80eeUt/n53POgTaQFQHn8EI2Bd/QSIj6Nw
A7SdiAjYd7FhllfUa6a+97bllfLV4oBn5onEpuGgI8L6euSrPYmrts7hdjn5KO7gnNsFdge6V9aG
1ryFzW1rd9frpxzZyeJkGuTsiN6f6Mrf6XYevl4VnRc+eEN1wzHPx3Ivnz7fsCKFjVBvWk+ohNVG
GUDbrtH/Di3mNt7ShnhORiWzPYcudQ2m6eKiF8C8xuKyIVsLyFQ+q0pnO/1K8yriwE/uR4Oxvw4+
qY6tBUSAIarKhVRjBAwLdzcl4Huwddj5dVZfXtB8K4eJCG9aHNYqG7IsIO6DyPmW8tyWJiefZcdR
ef4tGeM4q4BR8RzIlRl/+U9Y8ARXyrjid/aXxSjm8ooqO1wmgdWyVPQZhsyplDn+ARfSeSPB99l1
iFGOUv48NLF+M0XxT+hl05np/y5jG3aPNZQ4VNufyvpswuCu6WglrIfZjDcMkKLbDfl6WeY4Hmvq
76PgtrU/6+pM1duinScB4jthz+f2IBSSDk2tFUxtQUVAx3u+/ByGB2C68IRvnl3nAWupGQzrsSNX
+H1xf9OIeuAZoYt2La4gvdXQE5R6sRymb1NjuMhEkYo90PSKgeMxPmkzM580ibv4RTGe5r66JWTw
4EGyqSGqSzCDFk7ZvrqyfdEOldF20Jx91p2GNL5dhcva1t2uWnNLMm87yC/y718dU2SCxMpLVWOK
XbLleUYAdV4CxFRoqvJpBpVObgYJxi7pJN2dkaXhY4TNq3p0LfF7eYlhZWwCdtAAIWbnue+A28Qp
4ClMORmiJqbNDAXZdqi08FfeJvb420zNTvr7fKtcheDvXYtvOyC/WkVo/kmmT7V6ZIacZC04iIDM
pYYp76JVqlxpfOsrStRahTJ9ChO8rFBCFfhNwGvFur8uIMKOLS5S5ZN/AA+Qgf2DfqhXxfBnJ3yP
XXrqEFotgXXthv3Jgp+zm6cLVFacFzpKoCxl2esvs5UAsqv2ns7mKVWPAhkg3MshfIbt6qYDGwoG
UDNRH7GpVNY0tXMlo719gLIYWP0ns0oZRT2T+FemJF+GMzk1ENWhRlo4wUvirby1Au7hqUHlPYtU
36+VREHzCrJbzH1dmnXkt9bnT1Dmj+Asfkeiswbp246GXxMFRq54Zpen/9f0zKSrUXRGec5ChBir
yIXH87hLN2SyBhF2lhoGTEc5Gf03M8nZn96ovLP34UG8eTpBULIz2UgVHRLKhsauB+xAurICJO4b
mZ1nf36cQ/7uGa2qX8TrI5ymwaAJnJ8s6YCsNIIqBbynVorrksRlKnklxx+1VzUHKita4ClTuRRM
fVzNCk+SlocemfRYNtLDuf48FsJK6INqAgLpCLuQCW/YRNIv/f1IwXjaK3Apw70gEtvGnx/Mul8m
FfgTGHGkeJ6SWV+pSKAkivTJ9rX8NsakZobsYlw1CexSmrFePgTGWLVWrmOuhy39TILjC+lWyXUY
zThzmhUPojFzGrfEpn1ffgals6/Ci2yWvTanh8380Z3X518nk2+Zl11qVEXR5BAb+NU8APuaPiO+
ATwoITrllxRgqiMsxjg0/oB3pfUQxD5wubbeESMuheI3OTRb3tdTPsaZ9vJbQ2o3DlnrBPk2wXdr
qNvvGPzhwqtVlY92DTUhv49rH0YGrumhlwK0EnR9zkNVrio2UZ0+jNOe6PoGpL7Hi7YUlvYmSEay
yJ1OoTtPt9Gu+KRpsDwow0RTbvV8963zmd1FOsQ0odKB9+DulqZS/qjDtHH17hcdZkBXBs3nhl1I
5tQaz8HYZgnjqnC7SoyoVfU/WL0OMVny/+CUydgInmy9UP6StZ56Kpe5RyW9YqjsmOjC+ZJf/5Ug
5jx1sgzW2YBz63cxeI3sjGPMf/9KXI18IrNzhVEEdFPIjQFsHKn9oqvyaIsXKD5/2lFeUrsANLJF
l6VPKsn9nTOzxrtHTgb1iVYDh1+R9wjQZ59rgHIe6CFAeR+DIHPboIJALeoMRpn2egV95Eo6jRG4
tSn/id7CqPIBVg/UIe03azB+EE4bs1HGwVzoI5VUm1AvcYLV+rzZAhfHdn5GgGw7LcC4D/qbmbYu
+4sV801mZ6QqAzgBv1KQ7JbgVI2/QzQNyuEf2e/G9uAE4SORC6FBWuhUk5meG6jvWd6aqz7Dqwpd
Bp7VS3eJD8KVkBd7YpYFXmEeVm8kKBYP54/GuYs8aO6YkHXjORVL8dc6tx9I01nkc3j+wj8MkP27
0vgs22L83+puLwYJjfofiVQt8xGdtNvc//NSKfOGpLRVybt1xUTrX2kd7XFWs/ZUJvhHJIkesctu
cAFegzB58VkghZyk8Xlnmu3cvsh1NlCs2HbuOF01R/RYLXMGQmmTWakpBedgF9WA/2x/P/ZAIloH
SMfNd8ttD/De3vHIMC/gnSlete//wdCCGufRQLK0SMxFdqIWijf2OSqUsgZwM6sqGH+cC3MMZHQ5
9xMLcrE42qZ27F7wU33iRCkAdhhXdbIKzMBXCDDP4dQAyAVhpD5/v1brLuy029Gc2Iuo0BUS3/hW
cuWQVmgMLmcSTnuz/+x0bnRWpB1uIqTDh6NKozjhX1gU1a3Z0A/RVms7i5xfsK1nlI7KjLQP6sRa
9UB7s8TBe88eIZmlVIzaCZOT2OPq3CX+bUjxMW1+6MyJOXimVyyt1MoWf60Rk5F/AraWyB0hiyJW
i26i6nHZh9f/Ge5IuNLyyCX2HC5J/RYUxu9GxXtGGwC2cuz9J23B8EynHVQZfEwtfM029l42unoI
jw9pPgmmstDgtWuniE3FnDQBBgmGSji/hibvKPcGNyEmK8sNFmQIrLL1R8BivnbCaWybOF8m8UJ2
MEcpLhTiUMtilQGwiL8wPZ7fu8RfbaEHOn700pDgPe6Kw2ln78znPuTRc8bUlMYSXVSpJj5MqWXU
gaT+pzwGu3b1xPnje1cdka6HL54m/4s3gd2MzAjojehzJm9NyAyPTtxBn1eVinWyGNxsqqSS207Q
V5z43Hh8JmS/eosuC6C6sQxqmx/4SU88QTKBEBj73M+Tiqqmbx6IqMyllmSeNNWp4HO3+p/0CcJg
8ApJjHloAuhwBG5pQqRRkmLdz2OOAIy8+3OlfgYfpXArGjauNiWn4CRnUyD/eD0Ujy47jaPLjift
cZwh6ReOnIz82jHBnCEeMMurXfZj1ZkQ8cxfE8pxHoyKEXR/frOzI7FEPP/C0VHOAnEur+ETkyUB
XVkz4K0UxqzqNOHk95b8ItbpseG8mBgW8el7rYs5bxDklVfrGVcHtK2vPizi151bDsTSx2mGT5OE
XeU8k+vkRToNfwrtNZeLKIfOklrQZWwsf/Of7HwORziXK7NteN5vpJp6RqNDaRBCrXeNU0fK4ehV
SEH+0HVYweKzQVmME3tC4BbhtGL7rDqmkmGLgGMDVNaVWmh8ZcpbOHE5N3dLfgbNjr2br9cYkx9B
cquX1dPC6N/x2gZTsQIwfxDTy0JrwMiZJjLE4V9TidCPtGBZzV+qk/yplYe4rFjm3uG5uq7R1Urn
zPPEu5nesHMv5sgm1UD2ujfTuMTdAdJiamb7JiD7sWKds+qBtR1lQrsQXzV47udE+bAMA0bnFCDV
/C433g4PlVXcpyzGqe3RWMT7trGaKDSm+EQ5l0wTqWasoHRdlV2ffXyJEfLpDpGVifgyH+1LMjj5
1pF7X5255KrS2In8o3AVWvd4Noe2sHjqPajzcM0iLDpnQhIEzeSKnTmgWAOLUNFFdBtY1rrbUqMl
g44zkmQE6FXRBXhZahfEtLYE7sfD0c320TUwLJYGrlj4MPOUiFYhwYCLvHD3Gwh/1sajrFohnxmB
yLGleREKTgeOrLCWQP3a3R5jZM57DB2FrDEAr1GzZmazByq+N7wlyiNM0XsbDY2DEfV0i0s9zMZB
o944w7Bs5vmjQE01WrTJ9LjHaJm99Tj3IwTeXn+osbKjQ3v3H4TB+ZUsuQ5g0myzEFNjrkjpfmBb
rsyRL3qRhrYiroh6rfcsIoKQQPMcLd3R68d+1HsLLF5dktXPB8F86FVNxOafctXccUa0cqlG84ut
psjYslYtIzgyF0wkE2aiRgGyOQcHaSl53jZSwdQ8iplX3u755s+sPxk04rCX6VOqjiuNfzi+qV3t
0CxBHi10R4kwZsJUJT3ADQrhasOktDafY5ZGZbhEgNQzz6cgGD4UljnZccbc82ZwpBTfztbC2CTh
IIkLRQK237JixiFQ+28qw78Ggc3LGLnAJJSv+aOdfZij9r15r+PH4wcupREZfVyEWUoNKTxChxAi
VsMGeWKSwnRSOaSF1hiYHvLydmuQQ57CbzP3iW/H40GFLIDY1ObdVOOcuSeIdFB6ou6tbDspUY+S
7bWIRLp6+BNx4R4fICeqNuYox4e/QjdDuS+ncPLrITp8bhhHkVBPbPA1hjg2fDISaiSAwxJ6f71k
UiHGK0231zsdnybB55jCdL1ngDWkXslxQXQRfC2q7EaOSvoQSqyfb9k2ZP+KnktorWqixAlZZito
9OBUu+wEQR5K54cCAgbEOyTdn4zeRbzUthtf5c+6wCvEIhyQ+GVKVWELrc5xNVTaruKOAQH1S6Gq
B1UbeeICL9URqNBWg1DTF+wfuS5N/j1jVfVkI0+1naAwUtD7Av0vL8d/fhhsJQH95Em/CAsW5X40
zb/gBoJECYvF09F18/3ehMJ/Ppj4T7pxUsacMMTmFK3hg+coAL6B0H2eSqZarahb+wpSPgRicrBp
j4iP6pOWAa1KlFUM4yzOVvYmPoyVzot9WTwZs5CX1FiPzYrFR2S1vZPiq1ANDLpvzVcrv+HoTZ7u
P3Ozw/G37VfupVFZ9RtVng31AEjwIZNAxQuZYzEpJhRA4jazaiJwK3jUnm/lsydH+oK8wKOE7IPE
pA9qNA7Evnyhqv7+f2qcNtk0nDpDecOiD42aXPPJg9hv6GiZY7/ixDWtc89IWnE2EG2aY6Yih6C6
RlZQcl1BrROsESeLuVBrqQ7kuSuhFK0IUp+qt9KMo2iN9scAnFH96tVe1mE0Qut/P8ZDuwWKy5mz
ZMjrfOwunsiiAsWCriplBJgutDiP4A20jPW0cYWxdUKi+P2uRo9PgNT8h7MKDIuY6amGtL6HZ0SC
G9yR2hbVcTnYXDbu78c9odL2Ea1BDD3zkaiVXiRouuTSED9pysO1FqJc+hvK58N6eM3MMh50Cb3R
bgiCVr2wxPcB3UURpBUCnCsqrhVuK5E4vyeYinIUirYbxxOjOtvjLO+q36x04I96eDRxLqUQ2Nh3
XuPOuDyP5O4BjryiwZyjZfrwNAEt60ichpf+Tg/voiA4vdAagJfTCtpsc7vqXYg/pBwucp9evEt1
kW9U3uFs9ztQ4s4cFfV1acOLH+XU8ljDLjy0pRhukn6mD9whGIK0jN0sM0/th8d4wcHS7iUy85R8
L4Divf/sp5tOcFxX7IRlQaBNbLIyhrvpggsXBXgSXO2Q1/hVz+t9qidk2jJ9Z6DAmazkRG9Z51kD
KBEHJ3qUdwCW6pVV/CekxWjwGEAeNek/jpAPF6mikCGYs1Ujk/rTdn5wQj9EteGabiF8K8QD2Ksk
pQbaHZlToW7A+B+dzjQHlWByhOkALVebK7vUI3owvgXYghDJZEqtTRtS9FTtyl1H6VM3ox/5DHkv
t1DBm2FnJ+cxTpUsN9XeJ69RrC4MsUijfYemi9F9kVxqDj8x8yz3fnQ+HI+nAPMHhGCqnOwmLGaq
2VWQCHYzTut6uIY1N6AL/pQ8W1Mx/DOexMMcucv16x7yyfvPUuAysrbKaxq7B25kZJ8/UKFPd09q
SI9sCnTgrcvNT+oh1PBBy9P+T3wYRwQubUYc7luAisvhcJTF2zl75rc7L60agFRz/Ilu7RiZtW/U
MZXWQAqOLdaPCIW7/I2gRMH2tcreo+DJen3ZIsljRsmgxbEEz1LMwKagM+sUKaIZ4RjweagDyCw6
yfmhzmwVlv/DXZjJlr2Xi+VTe16FLYHkYQ2gtNcmITGJHiEi9r25XsK2QiZIdjbBjVVmB9kQ8Qwh
/Cz28JbPoUl6jkBGRG9Yfy4dhWMsfh/guxdbxz42+ZQ5ZxcraePtgqxdJliFXM+myGkyy5z3mwFF
nxcXq1MpcUJL1WUXhZgSQQFI90qV26UqveXd/AmXRvUKw5t06xr++N9KnfPCYEwnqWEJix4LMaIS
Y3ISPWyQ/xyvnLkTw5s5+lTzC8en49rHpsSyUcDOiMptGKDV8sJ9I4PhVv8enjB6/oTu8dAvb83v
Ytgj/VNtNrL1JsigDnvQj8WEywa03DZVPzcUaoLghdngKIRIp8h1caeXwiCr6b2GHZr9LSm/l9z/
1aWGd7OYP8PxA5KauCj+fUNmxCqtJIIJw3HOXHD+0DADT3j0V4nkFf2JIrwONmzAJUpGcwZ7uGW5
MzZMDgwE4N5bxQvpZaM1g7FS2+4oXYxRo4wUue6/BK72QOnzVOilPyX6FBvZqMH+Q9riL+BvoAEC
eh+fP+3xum0YZ3B480zCdjkf3jrq+WMC4EOeuK4X4yYIEUgwZTL7984A9G7n8k6VArEPRqvxEqQO
0SeQdQd9wlfZNEZzeATF8YM9ZgW8yRavr6JmiT0BYYc0S7iVgyuedv1v3kUSLlbpSWSwxtF3RIIm
sUmz5VwabIE7KNf3pVw8QBf67zaLavB4KdgDpeOp25dsB21ROf//eQFuEnt+la4pnNpvP1mxbcQY
wee/xB4fWBjldF3/XkSO9W/SLOUjk2VAcrKC6D1F9UfmQrftMFaM8/vI5pEqkvJHuT0FF8ucvzNx
L2Rpl8VTdjkRGRrrmi/nBmcfUiDRfG1WC7mJYc20uGGXBQ2s9OJtIl/lJsOY+Phk9mNNxCgIMy2t
niPJbSzunayA+jIhNGDqPznyQTn+RXHcjxtrP5Dlj+Ys2ksB4ryVmtU89ds/5BYSDCJaxayos+i9
iCAv4puImjvdzLDDBM/QBBIfoxBFhZEu0zu9dAdUmhE/MYhBEa1B2Ty1DzYHemMuu5vB8A21Gdc/
zDWsEn1gMO0crhMvWQ9NtT+k6uBEchhD9kgv2vYfcDbbyHrT/+7qZ5Mb7qO4sIYcYq5941GU6xHH
xjp0FCDx0iSSmIlD1VU9aobeh4D0TB36WwWigT2pQlj1+JsTSWX2sXWstOLqUa5ak2VqpTGLeHzG
aWxPcQsNa4DroC6K691IsTVPyYfETdlbBU2k7BFd1se3Mgufq/WitCULt8S+Hnx45Ibwbip0uwM0
D62mInK+zhJQGxNL22MHEYSZ3Qjwsqqd3ENJ3b7PXpK4MwmiWsZpFRgyp17m9wBFGHtfSrfP5DGq
sznxxUyF7d5lFRkql1tUeGQKEdwi2cy5t1Xu8L+PXbm5sm6uDkNfifO/r/2QNet7REE3R9CIiMkd
xdvFVXN7W9t9ERBYQO4r/WcACcK8YppUXguZty+n4We7A/5CkKh7RR8o0d9yv1H6OLm9ecOS9S+f
t9z1OJ3zPbrqy8rql49DpDl08yP9FEWAZtLNNjJfJ23GxP6QsrkWowMVWUgzn0zqod67Ibk/j3Mt
X0Afqk8srWCzUY43krPq+Kd25UD4xarKU4QG0K63+WUFbQUGpgvZ6mehRzHFbqRWb0lMF9iA/e1Z
E+tZ9tiCqoV3RyODpv9jBuHWickgAhSNSH7Ramof5SS6H0Uq3iUhprK++MiwV4+AXooE5rN+eRqY
a4mGhWgxJgnzs//dWa7cqC2eNrqk1k1SIx7j+keIfQpKyYddyVxQsLXhFDj9I4GWt8W11msVcDSf
duhxebY86Fjt6BLxYu3uAfMUeydlYkit1YHQ+hMFsS3Hs2c69keUr5y98K/sKLK0pz0V2rNTQmMR
1bpmOweqUE6gNp4LnnGBQCV+aYwjmX6bidR9rwHLMnVpyIN28MtL1jghLHIhLG6VRV+n7aZIbpbC
OBFPtP0oC4w+xYjSt8kwFOGn+c5rlz18XkU8pLfAbTLmEATTZstlga48a3InYFX6zsaQdLTY8AJZ
Cdur9KT3v2AKICDXQreHy82W8IvCWHMvbswkLXdH7c1s0qranTIPlrQB9/4Ln8VJj49OS+sgoM9m
sU4LcFtPMAE+2OYBwvXatnvVZwH0Qeciy4e1vlV4zOCgA/uI6iuqydiH65b/ZE4wCkJjkTudA3qp
usF6lYAM5VreB5pWVxOkerDGWCX48aGOTCcpt9NtQXQUTrpsThLlB+A1iiFKbq2I4BCfc9HEe41O
mHnVIBvr7OlqckPEd7hmtmcV9lDLxsI5HoXvhQBkmhInYO3Z9/3MybKaQAbltPzN8i+XjEOONtL8
9hA7rm4j755cg1HsiJP5Ufk6PGivjBfS1oKa/rxxVlRm5sAxtuRxMJe3fF5rQyjK8DU7BscMfZTF
Zk5O4d9z9FJNQys3FV69+APixJaWct/4SY7xw6I9IBcJ3qCF4JOzB1CdNtpWpBTfULCcJ8RAe3QD
ixXBjGjv9eP5IeI+gE4EMRN1N+3a6AGXRKKQLQutqOxsRKWIsH+DNaRHFhxJ7onaUHNOBs+fyHoU
zfAMirVc8E1in8yUOUqSeaKmEujL2H7Eq77dHqdQRulIEIo35bPggI89xG8ol9YlaSRj5Y3X6/Db
z9kpj+Ldzdv6D/hECawkF1YcUcxkGW1pLaJXaaOlKRUsJPuPPhNeWuXoiVQsO9nPKkEeuRJ95EpN
L7ihpZFongNNqDHMBfnz8Aowh0kx9L74usVpeg7qhjfEH3+XVAyvRqmMM1tZ/xaRFqVlkGLJuL1W
mxZQwcPqLe08gZzfglfBZaZZ2j7rrZFSy5ZIrY5Y9ZsAHpqgeCAiBke3pQOdqrgK0QCeMgwqlpr5
xdnSvKwxkUzwnZJj281rRwT81LzmnDDnJYZkvyAkf/aiFXcn8yv4PNesrskTWb2AbgDXT4XtS9xF
CYucpknTu/TgTwclC1nwOZsHNXPoy5wWWWLnA94Zj0kPwBJRU3IGNgSnFc1hKZCUBkJcDACN0Bpu
/i3Abt8fINE073DMGyy2g602voaxHcBi1pa1KysR1XnMtBDr6O1zM3V7malUOYeEgm3cXyHfxOHa
RuZXVg+pctqTm7AwELkIosP8MJxDIK20D5ISg8d7aYwCa6rNutjTAtNsKnu466PXZzaU/YM1yTQi
GBPZcUFUzdBQt8mvK1KWlW+8lb4+YAa86PudNNjezNI7xe1SJoSfn4GCPBx0ofAC2eBRK20Fi+1Q
YaoX3n7BKvvEBicCL6VMhePSGxNpZ7x7G7OU8+ZqtmoTZiWy1kgbRIDXPvMKkw019/j29JCu2cU0
3YjCGpt/o7yyqeJ+C8VCqYZYjiUguRrWemlDf4q+kP4ntu597jGNO2o1KHV+QJsOINeZTbm41jpq
3K5ZtEg/aPBq5zQvahvKQq/UEkIisQ2oLF/Rqq2KWHRbrhjq1ynxNwdxyKvo0jRE5vqh1QuG8iCL
v4lR2whsEQ3el47JiMXLXD1MrLOMsgQjrmFOCHvcOLJuCsJEl8V7U2+pHU6T9hipHEREvp0ohrUD
zdgyFGORvkOCYr4/Cs1TGXQWXoftHLsn3uL8amtBBpHk32CyG4lh/h5073X2ZBid4LfyQPXI5CXn
TFgIz5ij2DG4zLlwnITxOQrtNtPNVz/O7hd4xr3N8lBo5K/DkNTtzK8Gt8/4K0ca/I1Y3L6jHH7B
DYbWRyYe5jXRmHzFLUMvE2JLcD9sWxz8XpkSb5xDtLd6x2o3F+AkVyyxzboyt7uudJtEqqrvR8Ra
xMWdvtRUKpuixT4fnimqS4vvlOaz1enl7R3NTPYlvOF0XFSbDkhODfbLGvDpc3fGvUPdisoae04x
ywSEjsKjz2x56Hiet/kYlTCXB/k9o2j7fHmoUa1o4gEFLysoy5zoWge/r8ze+YCcnp6z6ZydC55m
JZVnZWWvtGH8QH2/1BpIOk/gR9H87d2YdchEcNuyLiQ67SPazmTnsczZyu79h+dFlx6Ddrz3s+rt
J7mizpKWGJnfAT/aWWFGes56wpNpYolg/SgnXVR+tAGN6kYOlC7r/AsrK2K13AqtXrVJ6j7oA/LZ
eXlUfqdmcrg2XF75ZVBMokAnNxIgTBrITE8MA5DppvRgCm5hsIKJP23E1qrRJ+6irbq/A0e/2Ecd
wxvSgwGeH/1h0VegypT1+UFXdxjIlpvptS5IboB6QIU4nGicB4bdeUo3pMeyj9V5xbmuAojmxYnJ
4WUc3du/aYFK7JJBscAKwjJe9/j20wzoss9i1SLvOYFegHUd+Dja2GEnmHeugu/+PVx2wf+dgERg
ZRMhTokjsvPY3J2YiX4p1pvu0NNwQdOPmbSGfECs3iYzc7i13XbpltvXrb20LIBZ1UDs2NGPJtym
/HPulsCQ6ozprKMf7414tMSQpMhil7h/LvPGsm2fcPzbPU5nOnkvnumUVtXGqhg0oyi6EM3FJ+aC
5LApOwXqRVnWKVxLHvmIFaSw1nYM1vElX2kdEk99aylK4AVf0BTH6e8P1GuLHtiTm3+T9L2acio4
9P7/9mhHrqSWSDdvMTY45FKH+EWdczft4+rr61IYfp2VghnP9eEUsYNc5q6Z/BKJTzDM7XQbrXvK
Ohwo+3KoN8esl4RQevvnEau8shlUwidolm27sFeQT6eis5IEGJLdoZ8ZDrbMIQUt9AxM8u3/MYsq
P6l4QbFH0NwRg/SfWkUJaSw2+kzejbZ4jaIBIg+PSDZ3dpsN+5RhlcVo0VVo2961Sodh7zMxrTRf
6paxupcjAknI+oGkDiD11zIo3OYTl5COcjj9VO6GqEcnM5ddhPvi6PmmOL0dHL7Vp3j5gJ1QWrRB
hiTuUtmKxYYiFqanPeLk/CuQdYRwrdG3lxlNnJkOEbqy08rdPSuekaFJ6w4EkHMPot7o9vS+ZprA
xKF41hHsZSL08CJDmelpy+KDWda69NB4cKGQJr5GA4+4H2RWOBUShhKGY90aSgzVjX2AhLLvHOkJ
Yxei0OSqUSb5LO80Bu4gNBpQlUfSI7WXjx5Bihep87qBMzX+/YMZ83YECw3Gvm1quU3kFbYaxkUx
E0K/TGUqbIChdwEkDDptzJty1HlmEiOwkIlR3dZsuk9P/CHqATT2qO8SKRm1ZRjjLbc0XvhZwIxO
CPGtZvQEUdoC0Q2mKwzeDshJRKLTzNh2pGpzF8C0V2Q3vMK5gaUjc9zx0j+Pj046k5KS/c2hecMS
gg3hJEeuOljWEaSBam1UDBKazH4JpaBJSE/upHdURnVkPdwGMQ6S15uIzvNGod8jTVsiwpipHE35
Nl2sM8RPRKj1s8rk/D4KjIQm09Ikj6aGlJUKeYDrPrn17jWV5pPvsLwPyg5ddOk3OiOe/Hg+9d78
gxmGAnrgUdLm3TKi1YsdCooixarcFPMwp4KqcLY0YQPrHrZr8Ehq0Y5qs+FSQ+poRIRtRJJQ0kaj
2I7RCX3gcKJaa8FLgG+PEn23yZGtzti4XLZQaf+hSudY5TQ2Smi+VIhadBgaJctYmINqA1J6QiTm
30Q99sCRyb9Xgw2YTjVBCEui1HL1ULVFhWYmJrgp9iW0xKgEhAL0LLPosHf55t1pIpfmyTl89Blg
9VgtqFFQCBEPz84uT5F1brckyaPoM1zuVwt2GJYJ6qbC2xAJeYDkgwbp8B8oZRgiLIkp8LmF+Ajz
nle+iRnYUPYCerrrd2IIdnW1IAol0EgnzIWF9Auo3irmwWE6g+6701TKbJw9zGwT0LiL6Zqf6iHs
ORpfkbLajtMztnYIVE6316qZ+4I/1B4teE1lVVqzrUrT+eOhrHz6x8X2j1FHBUSmaJ7Aaj0KE9iX
48M45EKupvlQm6BxfmziMFjkQ78NE09kyH3yzanO33cUozrGX/Ig7I0UlotYV7urTWj4JKQjwDPO
2xiggTd7Dl14yZ3eAiwnAdYwpUq/cd0Q90nwwHuFCoZY2xcrZy+dBHINdAVrfgtNsl+nTg/rBJMw
/ag2JaLZpFlJSXTijojnTb2fyfH+wZCxFfC0wKDcTBTZ3GUG5nwI5b5wmdG4t/xKh+9G8Hh2lnZs
XoaGg0fq2MHa7ALwlfhOUqOzYK5UOnO9ZOwni30N+4njjboUoZe2gbN14IezIcEleW7QTzMpW8KQ
nmT7S0CeRDrzxNWpGG9ndGiuqr3KZE3Qn7ggh1JATaIjHnfAxy+YNIGBBIsvIYLITmO4GG4W3vTP
pFFZFXqvniIqpN2YPTxUXldRc85Bve5LNrMSFM+2x2L32YKs4WmOrkX5L/1UUMhp2DpeK0jrxe/f
uVmPmPwkY0bcdYvEoP4XneLskOtNsVEyIXbOAJU6DL4iolycF/Pjdsw0MWuw8azHYXfKb2pgtVDf
A9YiUh3U7uOGOd53ShlPiursBZcOqq8+Nq3DhOcRaCqWV7OqojJ1zOXJqYGLLBEKFQyr+Zl1ky5E
zSuoTEWBZCtUAUMPDZp4Zb6fxPeaI7CW2OA/R20aa8fpghUwHx0ueVq0+VbqHfmu0LvKIjHcdSsv
9DggYcohNa6tH6VppdGVEEBBMlsi0azuDnfDQPKAgiv3/z8OIlj3PC3d/sVo0ndSRieQgWney/vR
DugF35Tj//pToavYizymKkbpR1SRV43GyijmA8Jsnvtsxa+JdOiispy/zzwPt594Uvn3JyaBc1NS
W0CtlRftK8N9sWfIGF/XfF2w7oPa4S5zpAF44J0oxw/obx1ptk3+IqIXHCmAOEWr0BwraItKPlZn
nuNYYrIX57hNS+EiyaCuWVxQIM1WC00fzAP3HClRUNKnOB6QZGEMdTTGIg/OfJOkEcu+Y0mnHHgh
jNYXgIpqqyeZvO1wSKnir/riv4bsfsrsOmaYs6YjqWnUqnW735vbLH5YwiblyA3PmFz40jC7dbqE
Ppa2XxmfziszCUiRq3i/7vuvH/zQWWkyCu2D4v851uS/AdfEvtXfJAghhPKs3IRPCY4FVWZnnNCu
oqrfTDYzw+dv6/JIo0uA6q/77kV6U9FTAvEfazyeCWlqEg2sAKJz07ovm3KM/rdbrjEfH+pSNmPn
a3TF/vec+F4jyFxHN9tWLMy7TqsRkY/3eDihpGPi6kLQEz4DpDrvqiVjm6xEcpMFZhPROL51eIHB
DJh8Gme6d0G9rjPRd1vCOdL43V49fhNxYKO2Xcga568LhjGVZjHk+2VUUx7qUbWus7z9M3xKZifO
k6HLfv2jkTPOwPsEfhog7Fqr4SDXqJxb6mhMN06GZnskC7nxd4xPq06VV/6PGWklLifvhBnWHjyX
4+pKof3HecjkNzF2xqBFEwShARLvgjHl84O5+Yo8FNZ1sKWVJEL//UzHPBVTHVXSwR9Ctb61V0TS
UmrOhZ3WH+ErIJDDNZ6AvfL3iDokX4f+PhoS0kQ/zDZg/88BKd1reRGDB3+eCbRcrZ8/htyk17q6
/QNEVaqXivWzve/35OG0zkrl8eYVe5/fqwwzlw+7+J4fL+sLjn+2C1xwfMGpuKyzo+hOc2rnH0IL
ZKJwPEvi/e04x1UsZJdyhbepnzRO6rnGnCjqmlRubZcX61c05lsRpHawxzlaB8ehOj82yPXSBNK4
bRQS4S0stwZBRoM+nrADivk7PIrtt1sT8VwkyCBdlt0pErX5sxkbYCOy8CmLuluqy5oDyUzGA80Q
EgSy1a7kEPFZs9+AiuPLP3+p9Vys5PBD3aDUkTTNxdplgqtfZ96CmbcoUmI+5z5xWINXqKT8/N2V
XAAfNismCQSIL9eAcnnAsd3HqBNEnXV62Ym6RTIdPesV0TLEXtQsFDiVNGgStEdCHLjyQeMu10dJ
qa9kqjNCvnkcEHH+81z/J7Uh2Fyg1c9RC3L0umanOVPBOhkR/ybePOVrkZANE8hj52FR+iljDCUN
OTSaE6p847PknLGu2HRQEhOVTJmdLWQDf+NsAz8g2U2IUTCTnYk2xvV9Xh44+liEISAh7ddTotRe
T5XEUx2nH1LNE4PD/JzKhggRoSwV2YzNOHpBDyqdzg5cT5dqzyNgpGuoMjLaVwL+nzRYa1eCe/LK
LtntXSCHWeAevjCKj5qjOkHEHbosHg2hnmNBg1TuCA6HSs14OoDwUxVUg8o5jdxoiZaepgthZ5k5
ZFZJn9El8anHCu79TW5A6cD6v5mltoTYLlySP/0hqHrIBA3aWojHDez2Q6zBKrHx1ar+sbO/EqNe
mad1sWy3fhXHUZ2hcAMKzh+BKdAqK6GuOwH9b+4zQ0DOJB9LhS8Wihy8eWdC74YLAQJZ8FR/oa5V
uJig5OWymqViQ3GWhMDC3LVcAxi8XBOElzH5qmr7MWTgN6O819QFr3zhB6s+rNSVciOToIsOYAxj
7V5OtN3TGMnvceUyOxsf8QEUECOIwAy70eXiSxb11O3MOihAA0ItFpK3lwtS5wt3WtNY0i1J35WF
ac8Z5che7IwirjUFkC888aLNUdkavaSMK1mAR/geBpO1Wk53EUUxC0u1OBm9TAxQF4o1su8GrFqC
OfjuhjIXx2rfv3s+uiftLbbPndbZHyDXkpsHTs1NOiRLnpqaWNsOt5M+5FKFWZkrCZE0MW6w9UzC
5bN9ebXJ7pdDLPIfsu8AFoUMX5TgoCT91k/bLSIf24M1npH3duaNsDNk50Z/NEzVK3d1luf5YZZb
DJKVXs5XUFMdyWVXpfeSiGFIiEjIX0jwcmDmF+5vcFVz2zG027xAZh3oVf7tnEX9LbDhehPaCIkM
Ct+ZbOToeAYV3fu/LQstvV6CJ3hZxa1G3CRzJIOt/a6tHgCcTKJ7jCMlA74AZIv7UE5iGWSvqVxI
WlKuAhTTxUNbXe6Cp57xe19o2cisbTBV8gIImjar3wD7l8waFf8w/gF20Thtl6K/kPcsa5SCbFq0
gLKQdJr8I92G2H9HC/DzeNN6eFiEeUIyYTfAjKNv559Ka1T0JFHgiQljNjCTmQSlBXxzTE8cxdU0
Oa1xjkpwUsyyUuBzse0y3UMB+ZIMNd9SBoyk2o7ixi+CyImef68DR3Bs2UyQFrtTTEq7uW+Skwwq
eGJzmn+HLECOVaP3W1Vb9Tu6kJ323aj2fUfyim2euukCP50NT3zhLos+Z4nV+oCyQ4Rpbz7cxfuP
FUht9YAj/9jK3KxfKJwBs+ZRzJd5y4XYzlTJIa7/evIYet5egw3J0LnB1X3jet7HolfHE1b/TB5H
qFMbXm7LmJqMi/SC+UpBcAK6WUcjT9rUtjfHzKxd3jDEw6lX01nSshU7CqOrDKb3e8Qavx+TjIYi
00RNE75zL7C8dvbB4pupI+990jt/7lCXUyqk4DdYN1zFaNtYHIOrRu567H1ja3QTupAmKXiseiL1
pyN9hsNUVHSDwSn//61EdlICccXnwmVNoQhjjAxXuv8KjGhvJRa6aTf99T/tHT95pMnAOatueeCF
5CXMdGt2tmhE1WRN1g7XJNDDRNxNpQGYwFk2HZlMQRa84gmla++kK2ET/5msfP227lXXGyRrHZP9
cAMl5zWzLgPtasFCjNYr3NXcoI65xvci7ycq7zdX5vtp9m2zl3bpnMTo62uaWK9d31S2kZo4NTh0
2AdqbrrwI0VAtIbYfjzDTs37QWSkt2/VrqqhHpZYCZmxaiY0X3VNNyJ47k1nfuWmDW1BMQFDaPr8
zzWHGrlUAbG02A21/ueHzDi2yOsADmymDdO80d7kSCU2QLvUtFbCQoIMMQM2tiF2fLakApqi+C1H
CptO4EONFjDnS8RIP2kTRTtqOxHULPmlTwEJZbTwJUNFX29Pb1x7vpix/M8OfJe2aTY5UidC2w0p
4Eh5bKiV1euA7RfaN2KU20yookow2SQ+axQZXx8eXJtoDSJZvIvGtEnnFoI7FgUaRywgSTpFyPfQ
nBjJcUCXAX554RcHDkWrpFeZE7TYk2QdgsLxttoptZJ5RKEJkYuMUb3W0THBuFjuRke4y/gYCfOV
6PAL6tiNWeJ1YtTnSGNPRCss8TuQpYtDwN2DPDzaDf9+iiCqUMX2swK8pSCW8S0PLjHcWj8+aoMt
Okv8iNaOw2BAFXy4Yg1WfYwDHad4z6tuxEwrqDQYKXYPryMzMYUulCW2Lu70+6sORYcNpwKwXKlX
8ul7DYKuSy6pWT+Ww2MEBHJdmeZjK0xHi7de+zOzD/VawK0uzMDBaaqZc8eR6/XLWvP59Rk54Dq6
7tPbw/8kID9dwaBFnY1UGj/zsf/G/Ci3JYSRnzB/tIb2qC41kqxUY6VvwndHjt6mftGIJ357H4sj
F485GDYTlnDfKcjLeH8GG6DkF+S/LxQjY1KbztNsc8H9bbxAQ/fbWXJpYqjwN0e+jgMTHQw/FjC6
/SE2wGyF6hhr6No8UZOXBrNd4UV9Po7FwNd8UVJ7f0A+SLG8NfZoYCoEuhdPugVoLEeL08A61dOr
xjwdQidhZ3NU7NAo6Coj5yS7E5SSx4cUuiKDlHWp+lvmbeiKuiKx02PpAtfAR78VOUY08DpvLiBu
F3JQI0MRHqTbLn2Hw+V0/bGPjceMDN1usQkqhVACsOCkERx2p+mfARX0iS54dcSNsglEZy7jDg7A
0H+flY7dfmx1gxt9A3bmAEIetiyh708Un+NgnJNjlFTjQjCsp+DcBA22zohwgCqxWbQR6VtsV3b+
XONkEkNM3uk2C7a4MaFSx7XKeYiinowDA1ACpN7KvtA9KG1miM4Yp3n6z7eZvDhMwKtllng1QsLq
BagzIMHiQ6EcpqTt7g0mHWp4WlYygBmbVUlrCqgXSwCSFvgnFwflvBGES8VlTyQAHxnyDZ0LVXXr
Rvy7GNW6jZpqNJC7FzAjizTHXvMwyJfEIYenJ00Z+MQlLwv54Re6sGVMpmk49lLAavaFH00L9zq9
Mbn9MSVUegHFtnTyrM5eAm1pVQ7PqSQvZXGxaj2Mbw5qSdBUyAEacmbek2Hf/FVKqMMqCpbbNRL0
erzE87OTCEdg0zD8jDK3QTnqPxhEPeNtbQcNPKiHsqSgUv8J8W8BLt2bGw/hQurcOVeTDL9PVb7x
h6VShSBREsxsJJQPr/rYT9YMJvogWOWT44dxTxWbyVCyI6OE2LK5scSn5Lw115yycFKgGiAUbFLS
J1XPq0HSYEaHjtgp7ke2hMoj5k+gI8W3roEPk4QexCT9gBX60esY0C1dOWi9jkLKvxrehTsUVeZ/
vRLzb4kH/RmU901+WsVIkaTn/vTebqPtZnNLP4+UaebO4jBdz/fh86aFGnUmMnAODRvgsfchXlgM
RKbwt+uBRBbEgLeVcvti67g6/IeG3TqvE7BlD+4dW+wNyaUlZpp6e+J7F6IEIRrqRABV0kWT7wrJ
HIIvJ3v3YpCZ5wSiWS686EiL4r3mIFpIaQCchvhUagDMxQvqGnDb38rhAhpxUEUy2vYn0WXBcjWB
BpkaLEE/c9yJB+8HUEunHjsJYhywZbB7KRqGITxfhUyP2GUJWxRI+zhfywmV+v6pUMWn3nmVsPJD
nXZgjFmP5uXE53Y/TQjaNDiG35VtD1WyttFVM+3HqZ5bcuRzCvAc6q5l5NA0d8efqQfUSbTvh0C7
5C5vAW4wEfCYCfoy81YWrvkS/wmYMLKescTlB7Z9x023/uTWZjyZtiYf9K23hmlefZC9dYQcPGdM
ZgMaOVUH4Gw5H6BxBLkXMfPC7VCq1zhu6ZoT7w+rvZk0AgQauWls94HwXNbaFbEQ3j1PA8lNf86v
7ie5gCNwYMvH2RLlO9Xyww7Un6rHSecMST/3r5b3peSVuoILY/u0VYgsxUubdugrUD+AIOv+f007
KP6ooQztYZqqP2vZBE5LddCCbTVGrFieFNYer35Tcgfi2rPzEm6hHX95K2xwbqCF1fgkvsoJsjek
3td4aANach8RH7YYiCgWeXd8mG0si009aAEOgssNJZ4ZjdVeA3zNvq4CDQpfobJ6vixTTGDnFAb5
cAUJ+FQXNreTRGOwpbNHUCc5L+E8ZyPHJbbtbeRQ592NW1ELghGK6aHqMDLpUBSOxtjmD4+o9b9o
e07rs51l4WpQkMsUmIhywuDkLLzE8iEEoMQ+NaNA6JLD62tQr4ioxZ9uGuGxmNeNnaKrp4tOySWa
UTzRpmuCs5sHUKMhxFrLyp0EGq80EFag7QbsoYm6KM+6E72P6nqJgFi5kvB950kf2hJQOPjNSbr6
J5aDuhc7QUlkFxYsNWqBHgixFAJvKM7/2f6tZhavQ58+pUYX03thVgi21uML5tELBlS1o3WpnmCC
mkIpza8Q4LTpWIlWpSI6okPbfMN7arM+P5wmzNuj4d6LXPk1aI/yPqfyPYALcPIdEd3zG6qJaVsS
X3A5dUbkMh5K76dEMpZzAtH0w0NKjP7sr/xKgWsh7mJfq9vg5FfUh78vGwsX9aF1sJOKNmL4JKkw
rBhIMbLcL4wYesd7W+NWjGEyVbY503hgVpedELUVIctPl9tQqFUvDfOp8wffyzVjY6xxAYVdLIgu
jjMZHBtBMH1GHf116qf5L4+LLQ6xiUVGBMVWC1oOmJwIYfYjK2WzhX1ufWml0oAxoWNRfuLyRX2u
RM2DaDAQQRVhopb6va1NCDiKt/9EolsRkzAkG9NeE52LMtDgwmpwiEy/97otaElPBwyIW+zHvgd/
GLZBWyr+WvjGGel7QlleMFMIJJ4yV3GLlfCpxb1z4wd/gdv9BP92BbdzeMxx2Kx8AJCm0Rdpki+Q
34qUiLwcdYKFRCumkdnJ3FVQ/mzUUnyDy7xpXSyWzcHnn1R052k7xjUBi6+KQtYHBGNfCcnJEzdA
ikS/V3M9sEl40jSGT0R5RN6iPbunxnyhLyL/ZLa62FTslBJtXpgr7pby1XRNaduits5E9uwYlXlO
p5WtCZ9iFvFgOZfK93fesx+r0jhPc38doTo0X9yXg1whOmVftilkeJWCHcdDxtGozPB/eUBWnHgh
wGEoOYWZROXyet4hJkJWw2SF0FFOzFahsu/VWQJfjs+8ZFRH6dhZwQDnRs5w87bRJzF0yuKD2Y3G
0DwoCFNp5S1WlVQ2wXBdarvA4l4tq0tKfMqOJ75AvDZfg/fZCy1c3JVsdks0VKTG3Cs+QbbKHdkE
ERZJrjEFuoXbiP0kBQsg8+0kTCAOwKvTDeTCaa1gajbuL1Y2sB5bW3RNnGEmSwr+APPE3QBcdeYN
AdX4Fd+16RjY+P1SLkGZbasVR6k1V+dgFKcFdPZOHADfvi481bJDRZ7DYnEK9B4WiRfps3yXQBJO
5d9f3SCZkoo3zlZDuNzXHSHv4ugyHwh9UueoFFO4undjMSbTG9BRWpZIxqgwQ+Nc9UFNhDV+DAjL
BhLUUMBwL1z+BLk7lwprpDkRVlHfmPA71KqRDRX/9Kix0kd9lRQTvk8Xm2VQteeodprCzMJBjkBr
SKcw2uSq1oePM/0mMD8tScJ0h30o6vn/ciSq4zMReGfLMy+tDfbXWksuNVryqOAMNJz3Tamjp61k
sFo154I2hVK/vzJGUqX+celcvRzbTYAgmw7N5vLFBBCje1FndoTBVXWcvKB9XY7HJvZa+kvsAVVJ
p8LCHN3pCFjqks4sw7TdX21om5cvRZbPd9JmqyfenEYBOVwV0K1wJrerOCr1++5fTdFlOb2n2WBa
iQg1qUEyFSH0Pa6s4BJVwXZ+7NjYSJm3QbJtyVdPoUXuu9xcVGARhI166t3Ookn35gW/+Wvsit8z
dI611zZkuKBVBnMkfCwrbAofMVOqY55gNhe6C7tdYqDqftrhdbz2mitkO/4Yr2xQB74Rs49DI7cR
22rTk6w+0nhoGHN9T9BHy/vrJBXma9a0pB/KF4H5LseJsaIOiCnctOOmA0vADX7F052D67+XxNdT
a5TAZlasvbwo+k4PIfJK2GX49B59tqwMLrLg0vEgne3r1T4ckemmbuJyC1j/iQYodlWZ4MysDaw4
68JONdVsafuw0ErbLyQFyQtBINSRohCsGuLX7XF+J/vRuDmk16wquc4xZPsP3b+QKkKb7eqfdjkd
1ANJWLiD0dN7M0mNYZHjMT+wx+HGVgi/8R9TZGkQf57m0LggOyAPIrCFXI288D8q4KlrokQilSnt
qd0cIMYt4IQN9Dl9NIZDZ3BbXTGKNt2IjPxxa5jABt9xiHulPXD5RA6UzOz3EbaYhXSYIkbgylQn
52rKct0xJuCYAPDU1lujJz6Dwd1XYhR10pRa2XdXXMaCrAhECwQ4sSCYlUru0TBfpJ3o7+Nhl9Et
mM1Rh5kLM3XHkfIG+wiVOuBqmcwKGHBXySSkllnyPsUnar0Jc/QQkWa8TlpYRTAmQT2ghFRCuyq3
4cZHowlE7DaI3NrIFH8ypnPQi2KTJLhOuA3O+BhbDTDN75xRYSfqrCNbk4F0oHorB456ZIpJgrwT
Ys9LMNPJyqaUE+RqKZEUXZozmerHbYrMFg8U0TJh7bVT2KtXbPxUCicEH9x4gqM9LYPA0/h2KbIC
F2PSa2vuHwxerRXJ4kndrbq4v2P2sWDZC3Ljp47Mr2LPxQeCbcs8+iH50MEjre8W1Hz348wGxriv
SN4EXc2+L0+MGtRnOp0lVohALYRK49y7BCDE9VXUatxThC3TyxNpFdgHCRXo5VzZ1bX+4WfW9VY3
2+tn5e4ytBWvsfztvZcuMc2BE39cBNEbMQICGrSYxmr45QyDFFAu7Bw1Mz7+F/FRbOg3qFGnm+vV
tY+wQvVNvMzrs81gHYqLQkgDtF+eKkwIIFUcADuykCazYpoig2JCmE/GZMhCbwEBSfWZBmMoTYmK
dIxz5lD9W8bz0jG6NmWy1fLYIsvn8tfKy11jl5wepAGgZLjaBJG2a9d6OIWxUr3GsYQAnCdsk/+6
CZ77O1GqrW44Olh+vilVnk4f1mLj/4i+2Y6TBxcVwOL2N5DsLffuCeqpBgigh6A1mMj9i8GB96Bc
3nOWXEXrrCVG+506EGDkYGxn1W/HtTe94RTJ2MDz+LVN/4jSDMC3cbh8pxaW6jlXZFG670N5cu2U
gBbrtqJIWf5okC1dxYxajEUCDVCmqpThfcnPMVabt4OPqBvZ5j0wnRnIT8Y0YFM3/ZsJqj0bQ8nD
2CrrnHrxcg3i1YUiMfRdiY5I28Iss6J82lGObQwZt/HmqppxXU79Dt3nl3GxbzOoyvDUAfkLi5YU
VCH9nQP1VcapWDz+jqPrIPq4rJtBAfehxc3M6j1GXq197cpv/wpTijO4PHnSODKCCw6RMKxyZiSd
K72IeOt2nZkTr2xdtdfnJmu9NmBB+R6ReOM5gLIHGHfJxv2KjMxU75DuFm4vIYP+h6c8Lmyy5Vqt
OsDL66olhPL/DPJEYqj62dfX9vF+DLxQnDot/TKuCceZ/+Wk1MoL8XD0tMuUormTcW4qS8WAE44G
cBGuDWW6xnfT5sMxy5ehWRNLRIfg0hLT9I5E5rroKMad16pVVayX8TJ3YfHrjciB01UEiMo70qhW
dKCapeQUff7ueQRa2u4l2oe0v0siAnPA4uGUJQtOd861rNlI1ib5rhoNBB+NnFWFXsK6Nqv7rCCM
7RBBDAZikAjiyOwmSfzpAge5isTtp85ReoGcJjaR1qhKaYFc2RTXejsZWjA55GRLJYZkl4VZYFcJ
23TEbyOPERPMF69sy6GsL+7rfjoKkftZNPzKJSiW2yCrB+MzoTfOsJw/lVJ36ftrDp90xhQdyrRx
m5aRf7U49RqxYE1vtqayV70k84kWrkQ9lBS6KAM3QYt6lQ6N9r0yh30RNLZl1EL4kmpo7nJsePYc
6lqwFmOkzLuSo9pSbiU81F0Iq10cawEvdh38+em/6+y7k/kwL5s2Irj/GBONPnpIUaCLyZESprFw
gtmuQdwCYAjsXb0n1P/BECaSJMJXZjYg3aKGq2FzCONYRtvSkFo8Y2MtnieSiuC7B2tuFSCWgeJj
PayDrjyamTNnFHOuGNgq5T6CcSSQZFUGxUY8fsNISJOwM8W580OGEB3UXJ/3Xz31hz2EktD/CX8F
qCs0a2/zohBfFmxZGf4wqcO+JABqvIChzpsQmFvSb/UnRs+63tCWxf+kj4UEIhEoi5ZCBS7npl3M
FcS6q2IZApYkx7JwsNkMmikUjrKoJ6ZT7h3/w3ywRwta/d3WzTUqqCSYfh7L2um8xfdzDELnzrCj
wCEif2ZUNrl55AQ+l/x0hnnM+EBOIc4mO4sO14X2MwhHdOSALzuroXZrR+uvq3gWtrjD5VFr2RmQ
hzLsAUndtioH94k45tY862iNf4ZfreDdWMcyUa6xT+0Bjw2YBxOWBRjih/K96shmbXQY9SvnBVgU
U9sbglvWmOhBEUG5NXPnHv8inPCEAfTD7gbq0/TLwHMgGWuChbF638MB0MqVzsd3Ms3qJUg78PId
KALUyl+3VeguqnrJFVzrJOMCVdF6Frjg/glUMqBug7I3m+utg4Hpei3TCRmlX93DQKte3rzdqjmG
PBozjb1tCmBtyGaOBoFdbGKeuwP6ZokYz+Cz9So3dX4Xfp12KcBO9ERHG+oNBSUGS5aGs0I+DY/Y
8Nu485DIH8EY0tv8DbxhDuldtrgjehHLvJp7U5QUH+HSlPr5UUIH3iW7lJp+IS34OV0+YLNDVeMP
fZNWTawdm0ZMso6s0Y2Zuisku2ReEhRyAOu+Xm7nWjpn5SMykMZdiWaHUcSwuNTf7p2vicziqij1
bJDYzHkNkfY/HwHNJuiUgaQQA7qeVAu5pGOmA8gnMKMM3md1YxSxKe9IJcWuUoHWEfkucu24tyHV
3HDSXyz3YZqYnbZfHyNo6TnEteSFCz7Aazw6c62gpykf0m9FdBI0YAPnpvAk9J/EPjUa8iT54yGn
PCiQBnllryC85xhbVOzGCWgBuCFzoouIjZDgQbpvfpVYYltGn4bMhRcIAjynpIBg1gY5n4AkONMM
ZdnxS83fCLzdrAkLkBKpfUrPllAhe5dmKYEO5FjJk7kJAZlqCvc8xmdRB4Mle1vbZY4xHT1ZqDBN
yvaxYcbxZkMSBZW6oVbApcdUbw0pXA0fJg9u5qc29LKhhk6YuEalx/eCwfmplEOvC7aCcGftpWS7
3JGxAE98WZlaBD8xlyBumpm7PEtr1cQ0S45oe/FBupmRT/tJLxNY3cd5fF5I2fOR0PZs1xfBwBSf
lUCyljfENp7RNDQgyXMZ2veZu/frotZWfH25VaKG1oc/mchpeT87S/9tOSv9QgGbxAS+Sieg3byy
rdG0EIkXgdLygc7ai6TX3ejEyR4ka3y1O1XQz2IXHn8VdY2WchDWVtot98QyKChi1Pg4rhwE3LWT
21Ph5P8ICPmY8ajo9Bepk5yb/4jF6t2STVyW6Q/uD3w/SYdO6wdukqJuARAexFA2cJSBJkOBRLCz
GA1Gpv1GuDka9CbKVTQMuNK8/+DX6PIJPUmm7N9JlP8yitLvTdm0Gw17bA8rXUdNuEV8hnb/wEYV
A61AUssQ7C4I+ZVAilgksE6C24h3zOMq3XHSnNluXjISZmlZ4zUGX0G9wJ7ePJgI/hoe/Mic1nrm
Mh76e+PoloIy+Yq9jpdy2SSq++CKt0KTQuxAZEx4ClZ+wD29CauniKHxHCRN/sd+2+30cBclZfPU
mYUwqGUkn39YPcnJ2cyWFhcyNQdjBN2+ucC+pVMgYTTRzcXVomG8oGhFOAI/iJLHMjkoSKdtLTpD
M+1g/gvXZd3CdEB3eZqeINK+bWOevsr0Xim6ejOU/oQXG12K1NwUnsdghuFApKfPKwEn0xIAbdxw
9QbQlxNydmTROfD0TqjiVBQzkBclQW1sXpvgPXkn3NBBjuUNpcIoJ7726kwHGP1YZfk/LGiSRSiI
vXf5HniA/DGTt8SSj0kYeUgulq3EXGZOgp6VJkxOjErF6Gvk5rIrMheLzayMuFrn7N53cXX+xav9
hPP83eHuNp85wI7Rwq8C2f0Ik7lU+6/oCS5Fj+iSXNz0affNJiuZ1U61VMYpVR8zD5JLzfTHm1xm
kRs4Bwuz8OiZvXr/O8Sh5j8grtDSqMyW/elB0edIVijPsWhsjkqb7sUmnXnxCH5Upqzxc9UL7WHH
cCUDDtq2Suh/rSkX95zG29rrIBD5ECofhDLlRcepnBHCLdpq5pREsuCY9ZO31UTCAjAGaqJTzGeF
OgqubFMMNpZMfFPRz2sqVcUF8Lh+pUkNWY0PKcZCEbYjxUbjrADz+B1SD8liAbfzdrdbg6ibo9f3
LnOy2OQE9V6ANIks9KV6L8nP8Du+KvCdJPJME1FBDhPBWRBxEi9Vfdnw2g7PGg4MzaeOjIfjwMMa
OKL5uVa0nAe/WJdk4WZpMTTURpUtjr8vefuWswufMgSiABNIFdcnXcdY70TFQ3zhHox1RyVRWJ9B
BQkBbwSa4iWmWS4/ij1NeEQQWKbJw+wtFpE+hZahsX1YFsN8G7LKpjDdmGroxiO7UoHKyeVlQ627
8ilC1SI2Wo7V9yt0gUXKJsPVVrpVKq6OF4W8OO7dbkd+/BLd+HPw+zkxwdfbtupnJmWiFk1Jd4Qv
dBR96b4zQLcBrecVTrJR5b9yytTK5fT0ZoFgPqIA1ktWzL9AoUF31bG2iNaav8Pxu1kQb0TmvrAx
7XgxMErBN4Hzj385y3VSCZ/g448P/WvqOk6ksGUH98mA4nJHhwtFA0lkwardVcmUZQ3eckZDFGpu
F+WTbOSpi+8gv/J0TZrMAIrak8u4ohm00KxVugoEQVx877HZ2T+w8T9SLUUh11LtlA7MK3vwOejd
CsOzZWuSIn+ApLYL3Tu3BhMcaSz+5lU3RCz2XOEk6xPu6SL3D8TnZAMBpn+h9ouv1Q0bErTcx44p
rF7fa2TK8KVzzdoeX/hQPUenCv4RzFe2PgNL+YWF/UQN20euFIVin2N2pLaWmgV99r/5vw8PiZuL
5iPaY4rV4lvza1jOLESaPNNP6kdmWC8tmQ+hQD88H/MctgHCjA7OEJqnz+cqqnlbJgjlaT+Y9q5W
N6GuRexO5RFcJ1Mtr8pYXYPrzTVAVuv0ogIakc80zHeWs51j8QT7yGJL86jS3FOoW3qzYgPHFm2A
2wAStbp/7QDHHh7qW6pargPzuL3uOQO37rAUtoPAnGIokCwjBExW2IACVwq59CBHqp/y11kF8Zw4
xZRG3gI87YqZC93jHQHyIloJH8RqOSTkNZrNZTREvtc9OtK3Uc6vIRAg4AV1YtIneVjAGpbuCksH
IbXJL3u7Z66wDX+u8TMkoEGsT6p/OndubFm7aW3oFC9ifW7vPjknW56Si7Z/vg3FkaBN8gsA9U5J
XfiK3tNOGGXkgwkwSg3wLrr6v0iEUXlTjflGzOd/tqrjTV2otZMxHWB9OQuKs8husJMHNbmE6OOI
CDj4Ix1nD9EcEwRi0GjP+wbPa2vLPDusrHXJYH1id0EQpgK1DozhgwSFklSdECOsajDLL6433v7b
+g0788z3kMV3RWcHCKgiM+Kq9SuSbR9CyfCahRPaDds2aZtde86zmewDJKhbTs6cWBKYKD3kHN4/
a18upKVwLf63R7iw3TFFxk/gnQUhDmXagCg10Kc6W0/KTLOMA7sPowaE8elvlvNQYssKKk8BNG1K
Zupfdp+MckwSJtX07FH7KAqWP8YweuMHUYc1qv8Xvf5xWb9/yPT7tKJE+vyk/v55oEue3CYIjTeV
QNwJ2MMAlK9MYO194j51d3gI7/p1Hr9piF5Y7d9uOgO/PKLmS8Vms46l+rZ9I5XiF+6YiQtu7+N8
zFHy6s1zFKzRQiH6PD3cKz0nzuQgYEH7N6qixHSnqYpBYFhWCYiFDNd3+skKa65LNQE18NpYD/9v
7n2/CkmrNL9l9n/Vxi1jMHa58AAYPvcGvNZaqtudxMFjptvbx8p3FNklFC30S1oU/nnzHVhrnAgp
524fTxTU/+v3BJDRYhcHTSl0tvIo4DgOx5GFa57zqmfz7Qo7AGzGJGNLKOlEfvqiNXuegA5he5K0
9XUDR9LK9v76IsO329XVsyjDXcYbbozO31tO0PGdMZDIUEfZw3XKaHfD3YMNaV5tSGbs0Fj5UI3c
nMGJkEdZeu89B+ASJ/4pabJoNZDtqXAzbfDHgZnv06pntw7qaz29xtt2SyPzXVDghWRiyEohXUnU
9dnmtybE5egPMAr6vh7TL01aGwDSaOFpEycovzYcyhiaX/XSQlMmp0tuIeSbZ7fi0PtAqftZq5BV
uw76CV+kZl1TX0nUgNBhOgVtIqw1BJapZQgmVGzGL1orOEimqUFo1IgD1s3SCepbCNzF22Nz1ChB
tnJ2BW8XhamuiIjBM7wNJU1KWxT4zVzNDheNbo8h4yYQ1O1EWHgVNNIK7pMfxglzyYfmSFVPcHnv
bA1pVHSEtg3Dwi3S0G0SmmqyjDJv/xlk8vJpw8FRBjbDQKfHtL6IIWGlis5v4C93cbNThnhZuBhm
3LK1V9iVQOuDvZC7HxLHAUReI2YjuOi5oC5E33xOTuVIn6GKJ3hUK9s1/7Df5muWP7JKxV9ghnu/
K0UecVTdAd5F/Ey77qsR1+KFzkuSXqGFGROE2flIZaoFjerocx1vpt0T1OsxKkzPCvu84dSVoxj7
rPL1gLk4n25MuB38qImzManhxvPqoqVOQJzo+OPb9UW6gqtqJjR7O9Jww5g+3FZ4W424xo8KbY40
tEPsuT9GuO4egeqRKtaas08d2AoRDQNlsUSfgjzmVUb8E37olxHzpGFVvhrg42XV8HzvtWHLd1k9
bEtjBRZbuYIH2Nkp9FLVs29/rUx+xuipR3k7wyuu9SXMzpJKU+VdailPDqYX80eBx544x2jAvtV1
lQf/1zpgTd/JDZJo1wLQ/z+K0FFmAZ1Nv2VkZ2oW0nAyPJyqJyqaUpUQRruTYCQ3KaaSZuzhidWo
EoZ+0xdaVZSFzzYmht9hyHwKqJ9qls0+YuY6AbBozz7qMmfwD7rE7hvBZqK/rT51frTuQ2BgPL9f
bDsZCrXcGBdGRTCVOaXtBRbNxz2Unvg/qToPSvrIx3u9ZdXRGHCCCgSZAAiWtrkfrN84oetwbNgQ
3rIg3r0dPvm6UO5Y0NL5vDPeJfqic/Y3smtnYFwdUlGCHLkXszAav8db0MzheIXMKE7qD5WnkeCz
cO5TBByqOU//deDOsF/5yn9uaFQsnfWIYwDfOcNpm5VQ6sL2EXDKNgBW4PtEWkRwc/gwlzgySU6u
HmDT9/YjhDUDw8YwkH+ZO9vo5U11/uBrUX61TdecVEaJcJ22VQ75QeFf55Xag+1SMLyRagN37OsZ
b2E6X6XChXRe2UEK6nejzq5xj+c6dWACpl8K1e45Oh8lGNt+aAVbIr3DTaDUBFb7iZqVN/AyusOF
dlbi1ff7gNvFKS/ljP97x8D15RXryfEubWpi6XLkr8gSRvzha8XuFIn3ad2nXsiPr7UwkMcCf0iX
woWYoJylTcwM+sejclk9wgYzcYnLct0RJgan6Z2CVgXDzeQTGUHMwWaFQQr+ikz7GgEOwlI/CCYY
+sbZaiCatOGe68NrZAgei4t1ruWo10Ry9J4cBGpz5FHRCzYWep49UpI0LhtGiGq1OetryZO1IAnS
0uf7tipWg52NlnnwB/pxt3F8wSMoEUEpVCG13kLaEo5IaM6ZNJHpU1QIOiEcvRHlID6qapF1XHPo
qRkLMO3COgzYwkHT3EJ0QY3/cXy5FrLIveFzhSJRNBgbGaR9/P2LyxDukTRldjrA5b/I0pOghQg7
0d+wPbAlF0N5y3HFRoTvb8uxnxlxayw61OboLs+ZCtdMuuKTeKtE4bbMsKbBVVYQS/R5t4TIpYOZ
0tcdYopCMiZO3vCK+OU5tJGnoazEOQ7rbwyb2PHWSsXwHebrFCKeDIwMpn61fhh6AvOnURYgHcFd
yJ9wEZAJLjaUODRETSVxHRLuSHY4lYNE4nUmxRj4FJimU3hQ5S4m0VBB1w8NsOKRmtvqfUk71opN
0SHZfuhL4y/fpyoYepNJssZGjrMstU3JSPEUTIT4JHaVkyojma0KCxw/hPnfDbRWaNXvmF21PB10
2sei1yKLVZu3Adm/j1/WDzoRIejWh9T2FTin3WnRSY1FUXIgrPHMIAlBbPq00S3FyCtedUkxU8Tw
XnNcG16Xre5Q54VvsgYDuC9de06bFvwJnmedL7BZPcn/W232TQIDxIgFm0L4ZLsJm/GsAqCOcE7Q
m8PpBw1I+Xq+EjeWvPCzdFCiVKch0POoTfffycbMf/E3r3A85RYTF4sr8Ds5jjtN1W8gNXL+e6G/
P5RDgnm26AIqG+AqrMzic0qFTGRLndfFzkH+rq29GoA9Ek3SrchNAoA2AtG930diBYxSqdRRG9X0
/iHs1NyH727IbZRSJRZ5ENym9JhWVaDtAMgnCs3OyD2dc5HVwH7BDfXDGQnkezdH0wB4G2adlijm
EI0vl90aRCdeGh203UvoOdHRWzfhWqa2ajB2taMB59JE3eSCrPdwDbzain7C+6/gfPnwZTIuqBXw
0svM/iwh6pmSJ4KVtL1VLIGCsxE4JCu1UGTT99+HUZdsyNZGHmbaBKG8vhUSVPQP7UTaZkA0ByCw
426QDrWdlXXyC7VTWG14ZXfYipKUh1WqjGGn5AgDcqtbtWAySS2Zi+c+G4b/b+J4/VgiirD45Wl/
VeRduXTg4xDNp7t9mD3duJS3+fULlFjYGMIoZjTy2tQz283mC99kEbr5X/9E5Gyeyxbzf/5WbiNC
SOgXHy5McaWn2Q6uSgL8HHRJsAhE5QsTCfNN3McCdqzwYdOcHDkmBO44Cg9B5gnoR+x/7Ez8cdi8
i4hxvY3J3LjgyEerzcQZoQ7vbfGiQw7wJBF8l/onw6fk/jDwCRK6A6nbA8VD2siKIPXZJc+NG0Gk
NdNmTqQKtDYkzDnHhu2zjPxOYCfBhO8Yc+OnUgcRBeQ+nTXBPAIflgFgIddYt5nF2KWkuH0JhTaB
RuwdSwAA5zGOev++/0+eYr/rRuF5Oo6hjPSWQeymzjZ/EVSPqxMRGvue4YAg0keQvREspeeJnAb0
+BhqGv1a+Oi2trxNrXgWBYby6PRjc4HtnDmyvRgr4zWHH8MAhApkXdCQkn7uq3rniK+0dBEHSEqE
tKo8iJBXCpYv2szdq/cPk+/zwMQ8jb0j03BQ6IPAxvYcRbGwmFol5bF6gnFncltpm1zk1ugAo+pN
+pjqJm3y6h6t8eGMprGElGhWaq7VUoi0FP1G+U80TEzZBcPdFt56I7jVUNRXVYNI9+Kr6Yzs2Gra
kflEvIcBwr1QDHYmgKLSMZ+jyooVqTYxr4mPjXYU3LWlIrPdEi5ScSin8HrPk4DKZNDY3r4/NgO+
GymibHGQ1/MDFcaQQOhZXwV3mZ4N2dyxY1gsUF8UY9TxdUqARCLkO0Zf4e5aP3y7LDQzP0E9smtr
bkeDvmuWwL+V2gtFCO0uFVoyoFrhISoJqnRajly56/yVxN8eiJprIFPwR5iSXPS5SDurgVVxq+gz
zhD/9F4XluzfJiKBmgSzYpjSFmg5ejfUWRjKtUS51uiWE01EcKhjgwvKEoCt72zCPQo2lLWfnSfi
+0nYub7O+zcAF2FJ9E3ZN6SdY5S65eAgO3BGOudTw5Nzl+BnpsxIg2vj1drrgCmpoeHnVH5BGrQB
1pGHOXmonIkXecQ+Uf+v1MUQp+KYzOQDIZqK/rpPNhjZZKIIWjO/SURun3z8IUM/5JdLEPDCNJi4
JA5AcHKgf2nLG/84T/McQhAgs+q6czWmpGaBMWlzivz7PzSgI07tDjSv2Vy73pCa9C2oZx5JvdCv
San9JlwupREQZusnlDNcQxqotsFswsM7wpFf/NtJ99om4+LhTQr8HJBfhb/XQWzXuTHZpgszJF/r
bwAJOwLKX+WhCC9UBk6rs/9WtRhsOK9EWB2XEsDWm8UfvJUSBYdVgd6wO/ZD18rwP+82QIqVa5fM
exydv6nUS4j5O0Z99qMEuKywXW6Lf846h3L2XmIEe8NMpDqTkEqSRG0be27AvkOG0kTsXiI7j+iS
Swk/HoJ5YjQ3re5jCvvRygX8/BShtEGyTcSL2zq88yeS/2q9KXYw+zDA7VBCrNbng1sjMpBFG9kz
ZLMApzVxevw/bGsiqDJok23+9qz/XRNSdlWS86ya8y4ZIaQ2St0HbDYh51NJT2psug9u8X6ids2I
eQ0oH4+cNvdSRlwQZX2qhrZRn/lCd/dugrx7zrBGUifIH0TUDHE2zoSaYxOBPK0DHgkN0ReOXkym
rw8Mqw2iO5FzYxN0+qqEb+uiFo4Pn58aXZ9fByKiRUpnDD/5ij5Xd1RqzcMxxuFtsLkpxKzaSwQH
KUJtajU+Ijij5IIKYtk/DGDNPa3RpWpznd0LnFqbI2C3UrxMnqLF27h89fd40FiIeeV1ToJHQj6+
W6YSnU7uP1JdDFfSrHGj6grYJt1PEIePjJq0Yemwf2ZbsbiHeEJgIvfLW0H+CUO4ysOHVlpBl+Of
nHOTGPPmHSmHqad7mpu+uVXg2gWriq9yXiz1fjRttRcO5A7O+ON7WmmOJOFStD4iuQL44oKuluA0
kRI9Swa5Y77YIHgcostshQwoVTgzg0uDRUX9A3FkvGsA0jF15GaawQvCqwMi+gY8PH/db4D6Zqwf
zzgBu4yg7n6YbPBgJ61BTC+T1USBPjLMJi5ndgCFtSlrI6tqyYpSvYrir9bkaZTQm1O9DxmM/c77
9d7hFEUFymTfDbD2CaUSEdXWiD0UrnDziBy/AZ5br1lM6+rrc+SrKCtPwVGP/vJdXoeAMsOwRYim
2e8sMD7teau8lkZ8Xg1mNgVN6XxK9ZMddz7yW8lqTUhujVGby884OcW1/oxptOPqVxsYauBtHlEd
fUOmTw31h+PcYjvAGNkAuwhYXMb09CWMd39kUQ28R3Gsm93U8v/yjHrWu9r5ov8GPARBERSYTBCg
/8vflz/fVO6eEaiEU7x9D9JTp7d2XhEHRpPAmpe3dfdTlRb7cStJEgFF3Z+e1S4s6eEIKySzXw3F
EE78nPeM6fdvIM/lU1XE+QDtht7CRxNwFT5S+xLEbsofrnZbdf91IdO9F83PX65t6BjVEsbXG7Xs
1dPqu14tL1NhxpVhcaDEIE1CCAdWYS/1uqPiY+JKkYkzQe+A1Rrhlb/9OK57IXz4/8A3bdV76Wuk
jHBjP2t9uE8re3kxAVtdn7fp6ZCAa1KnIQzI4++vLH+8iZ3lNVzUPJlmGFh8kv1n6F5dwokyDiyn
AttW2JYpekl8FTeynAeS5ati8R7mH57HaMigPeCiGMupb7gLH1nG45mhy1XmuWS+Moig7erdjl0D
Xpu7xGaFREETRUCKEJKqTd4/ZZe74AJYYpaC0eeKWFlcGj7meiRa7YfEHOd7aNOnw4LRulDtcFsG
3Nq0NtHekMHL+DUDwAysKXyF3MrG6uUJ33j6R8MSDJYvlLkTea5+Csx7AOv8DKMR1413Kkddvdyu
1Rzju6Xl2OcGL88JpBwCvwnWA2V7tXNe7IpRZCXuWM/kJbogfLdSMkyhDqDBbtrqMkynrs7EP25J
9V/CGOOT+DjvZtSLLlXIYGLaFK8c/e+79/NTqRIrsissdqKWMw/yhwUww5Ie84kXDgao9ae6OEdZ
TNAI4qS/X4zI6WhPpjinc7QqIHdij+vNYUs5qRTjNTZb1r0fpKhWfFJEvADMWrq5HCw6aVviwr83
byd/kkGgOZYQFpBRPvRY8S6lBYQLjt4YPcOhjaKJMhdu4+W+uJjAsatTxldbN2e604pnKyLTSrVv
8dD1BXQBWYBJTgz9K+OEHAqwGS3b3/M0HmU35AxOiABW0j4iqv6WepM/NMMTdgCRAaV/W7E3rNC+
Px1zAX7Gf9mz6yYPQoG+4dYdwUShF1Mcm3P89nR+ekOHOdKZpfK98UCCI0sxFEm6CHh32ALdjcG/
2gzA+TaDZAg8TEPi2sfEXIUy5JnD6ifuCu2ocfP4JmMgURF5AsRVUyYBdzcsY0jGa8YKj+OvBqS/
4tQyKDgO1q/GIzlIXqKNEoZ7pt6kt0/ay6DEiwuSyul10O8KOwVIPcmkalLNM0dnsijTwyNd6TML
nkwRyroNYVNYbbsoQB9BOdBzlb+sOPuR5pnIP/GMLhnrP2kiBZPvztsKCsFt2CaGmi3ur+pkZvMs
RSpDTulE7L2mWwtc1L70E/O75oSou0s7gdF4/1VgD0v8M4DKGcqIWhjNHatMOKpbIBlFZKN6Js67
9+3foxU2X6+Lturbrjujm4D43IXlBvXNjzFf/vJqsqKhTtiKQnfm3DD4nsr2EX8xEbfZtb4acYXo
mVbAgKB8Cpp2A6/QP7O6E09cXWjBXngU3fP+nPDMpZ7uxFhS+U09kJttexDtU5xCbFS5otO5AH/6
sD/m+hBika65aJMd9oJUZ+OEsfSrmt1YOozzGQBXCCnbv2MSZpTYilb5tiKzKqaLEGuYpQ8Cr4IU
8SceVmH2FZX6wjnTXuZuuwkY1OW8G88BVlwVgfDLROJTQKHrOTAxf4tadgiFmYjjNjcYdDQjEjym
CPg9mLg+nYClzRKWK8jfk99bj6S0T9lmqVG+XVoUa+QDLHsISJUq+HhW04a/J90Toj0+0HLmvQbQ
jxSm/HIb7aqmV0hLh2GVFU14tY25vrWsdYW9IhZGKzb3BRWLSoj5NyhvmMY1k2xi97cQbOjQ6bVb
94eINabuOeR0ildQHul0ZgQF51tlE+q/M2HBfBGTaJLFyBKvYPf42OF0SowAT7kryEEwayuifANp
MGhHzoPDj1vE/pCEbh7/+gb6X+1JZZQpGvxbLQ1IkTq+vrn7l4ihuuzbG3PObd53iq4tXkDLjd7T
Cns7MGvyM8EdK2k9VGwKP7GP3lk5s6CcatvnLL7G00QCLHul610W3J0GaKDJau4tFCuzPD/ESojN
bepHtoz9jUkG4EyBtf2UiS96B2hOa1b/cymnM5DbnY4e3XnQe2R8Z1wzrt9BzYpvrGmALB30JW5j
eqx4tPRB/bvR8+wwsQrPFUHN6j2FVcu3BUFQzkNokK9CnR6OHWPTQMKruV4s2vXK76NyDqiO1fSz
mkfHnjyhP9WiJRo8m/aY8l4z3J7s/H20mJahhdZJD+mcje/tQ5W26MeRZAqtEZSCy4jxRXTZsW1d
QVVU/QcSrB8OX/hh3SK+DE8fOH1RVPD6Yq0IjivmmGdYHgODspO8AjgHiCyu+7acF0XuAHhdFLto
wdcy5vxo5tE9O19NDj7e82ip651fbaOn6x3rzplLuYgD/eunEor30ZOMmc/FIfwEECIWmrGPpHW/
5DJyKfrRYwWAaGclrc+f6ZD98PCGRn/z0grvwAZnx0lwTEgQ0fhVayR7QU1grepo3JD69jX8nfxY
tBWxoSvtg+UvwgN4s20Y2ENKGzjjpcTk3+ZiayXApKYrqhlqZ8q1pVjjlXOFpAGdO22aW9R+TZxi
kZ96ADKWYzfqbenwj4zZtx4itVwOqeuFHXpHSjZg7F2i2FCiPKB7C2XNLPLDQ2IBWe0XyX0kyR3v
tqcMGYpMcFVmds3V/jvbr0AAilPxz0tcfNKtu/M2ZQ0diWAWceA0xw6p1tv++yCm68wOJEbyci1m
F1GrMcdeNHQjP851DdyT900b/weOxxiVk1HCkcx1PzLkvTqfw4+fb21GSUhxS51biOH2+GYY9yOZ
u+EZyfExVpDlrXgUZGDHxQLuv6FtjV9uKqYzoZn4/4H0207NC5BzV0PS538CXa0pzi6yHRILHoGi
yvcZXJ5pFvLpR8BzCrU0jxKEkZxMqVvjB3dLVCZ63nQ+azYxO22YET7jHRSTb9WbcdvWvnwa+zKd
ZHUmiEV7X40yiR25NMxZ64TbjEDU4Mgzm830Js4GkVClNb9tJ/4/NPkGKSCv0QnUwCx1mzd2cVU4
vnAG7m6Z8rqKaS6UFt3TLL27McezqqOaPxUnjqi/UYW+Jeb5xE5ni9xDkZwEH8sqhiZ9Ua4nxY7g
x3qGxc/waLkLTmzBdBkkbR4hYWdqFTlHiqVQksWjHvRgXzsfY14dBnlCfk5Acr+AjLebMXVA3/77
zxvqgmikJYLX88znmwj/VhyiOYTviy8pCkHVvzE24dadgkj6W7u/OcwO5TI9FId/PVxyjFBmatGj
sqnc3wMbfauWn684oDk40ksOTVGbifxBEltQ486O2/ig3Gcmut5LPPgexanSkD8YvnFHFW2Umzp1
GzzyoS7OwvR8ULmMbgT5l4oiMRYDD8GdphX8KpnX0rcfB39I8boNWaeA9X2APa/QUl6LxHyJJADe
WTRWQEfOISh2MzSB0zwOT/IgzEQ4HL5v+Cydk+3kVdGAoCf9mU8QPe9v4TeLAgMwxpaSzGIIjm+U
dd+KbYgiK3Fb7KaJVtQNckFLpdQAQzmVZaD59FHsq30o9PHLInsoApMJLvm67upJonUg1HvnN9MI
HCKGdq0Dzevkk7n7xJDiuQXiTO3ykUsitHPlp1RVrPNvTGAm7jshyMtenbdV0IZAeikYiY6RfCAv
oQIHFFH3E/bXUHfLAR/PWy5mOe5I6lpmys8Aw9NQfwtC1an05w7a4mSl55yJHRMW5Y+EgSdB0OUx
PCUg0w7jQSNJ4Wp4G/U8qlL4sxbXhAr0hmUGnVu2k5x3/EyEoeUi+hmOkVrvDoiD05R9uufDWSKM
Ctpkq4I6KAh3r6GupTVhUDOslWPWK1z65bgPkaQ4OTExrMLId8LtwvOAsPUgWTFq4BgMn1LScO8L
YDk1Klp82rYfAz7fsHJDWGE62aupuS5gJ4w3P04D+BtwVbl5aW5z8K4NPSRPLpQ278DR2SSWvc/g
OVzQ8ipua5IFUIUpSRVxQdBLKdX3iqE2PVRrp8vONAzULqEvkFNSuPmvytEzAaJnFf/SAF/eog53
PyffvZYzWFV2z15cL1egOZHJa86zGNO6P3QcrwoPggsTH1SIN85zJsaglnkyTcUdPO32OeQUYcEh
km023Om24kh2iEsWo3HDTHcOLX4MkR/3pHPQ/fxDyA65gxB9cSaBTG6PHmkRPlrtU1QIMHlFbaE2
q/XKSB0AK0bDMu386ff0PoJBt2zhIPnxy+RjYmv2HuCI82a2PjLQd4v9Gh/kOPUciPttt+KMmY2M
dK+Q7FgnhVdF1QDJXwQ9qxseSaFGl77v8X6FBLt2iP/ak8f7YKUQIMin34dXDlzTyghBDl6nbnyn
w6T2D5S4gYA9AzSaiHqX5mjG3GHTFEBC+eIqWYkLju5hSTn+9h2mCBwi+X6sH+d3bA+Bgqs55V5I
PupWlXJ7RcyJuenTT0/piqnWN/xeWG7mU0xoUtKFlRV8zT5amy3//Lw8yC92nf8X9DHegnBREGV5
QJjyu3WJAtSzyywos1INN1/G0dEwfjcFMAokVfGVSONNPQw79Lj+0E4U8PONx6CdiHkDexOmAZzK
2aud80T3+7IcplJzpmAymAvjkqvlIRY9ZYjj21/esR7gZ1aqf4Q4no3HETVDdSBAFQJX3CuBThOI
v2hJM3/gVzuig6dj4fd/4gYUo6dy1CuXtH3/S+1QziiG0ekUef3fVLFUpfIGbo1iOy/k/CZx8g3n
WJCfC0FPD0s6xFTAoxxHJlUTRYZFNBvFp1P09Lw2tebZt5Wv1d4D4rrrGF94a3sVN3FX30aKy6v1
KlPgN+rWxJMj+2zheEbpzaZcWx5nCL8gJ406FNfBBqf8jjqZoYZN1xTYMS7Te9tktZGuCvBgS0ca
9aocFA9Ls3AnBJd3lZ7mdV+47QPeCgvTSy7hgiApEaRDpTCbO2yB1YpJYyLDISSSLvQmaHBjqEpJ
kR2CsQLjG9NRmUB8JoIwvvyzietFN6IguyUFLn8MxGovC+gQAT1+1cPnC5P0dNx1/ZzYW+0NYbRe
3M2/hFyOHmxjg+wvoGB88XA8TeHMLVmpwK26DbWhaLQh720G7+7vHFzpt1xvTX2OckbBi1Y/79C9
Qvuu4wwt+h673g5SzQ01Cas8CRHnQYCTXBo1v7OIlKrLm+XZNFocst+Ke9x34iJOzs472QaJKVlK
goMSdUpLpVnW/PRlRw82TdSFWr8uZ4CAAQUI9fbIjWkoWKSKNdmJd9THGPE6Yxc1QWXifE6LCg97
gOzE2Y0eTCL+rAzYlpEdgWbprjlrq57CVw3CtI8mVVXvHcgFhgHvVSktYr/lHs9PNJiLOWJRUzpN
jYaZY/ytZIMzwsaqT2l67uX5p7lVD7bM7XgrzkUDCjVso7ujLQG906ikDsCYqFt2R8qZkEghjcmL
awIhU6Ux2veGsTTDEbSb/wHpyo7rLV3NkIAX2Jo/I/I4Pdbs7v/NtaGQNgWA5n7MVCaGAViYowJC
ojR32tVFi7yFxkMTVMV1gg2cl2RfRTrBOqX/N7subWkdkIQ0IXFOksQSDuRSDUvYNC6LbMf27u28
hLqf4oidBJlV3uAyrlxZXvkpQUIzaZdxjn04UMeNkxpOY+b18CATNOFuQkxS+0sU89yQaBThyWHz
XdW/rSAgVJW70FeiupJDB+MRnPW3GcPEulrE8n+/pjd8Q5D6m8F/YUkrbrU/u7t3/5LM+bKwXiIA
QRPOGuK1GQqmTVdFHeCOGqQbTZ8RLVxyM71po6BkkKwvL6iS4CSFYBEgv8vx4XxDLFKUF19cEt6K
mPFTJ2X+fcKyi2rzqsygb+DGvuvCtXVV23bT2kqlu9tD4Rs3LEXx7uPfeCIkBctVSH8OEimCwbfc
i/79W8ilxhP7T6tnk60AtPH+Ir68KHx08OeFRXAuBIdgSE26YHBiccdthKJz9LLRokmkeAMqgz+D
YgiIUPY0UOtDMxBokV2k4ud5Nz2GsR5+NcbwKwacRyng7xB3+D507T2vgC1eeHSpvu8GqO64DjnG
y05as0LpVb9nU5hR2gsuk4tQ8mR6JHKT+2dHuHfC9D3A2Y/PtzfRxLm23Shei7dmpafGyiLV8QjE
jUQn3YSOgNJ7rveRuzgT7oRH409K7mtSo46HolygDVqD8D5DWCtoQ1hRY4DuZCoOkP+i4a8J0aaL
cwwfNFr6SVBRZaS8fAJwR9ptLeiv/bxTuz2W1S6/ztmCe0Ecc/u3zHUhfwv4uuT9lNpV8cwGQZVT
F0uZXrIaUFNsYKe0X5ZaRUjV/d1FJJWUNJBDV8/qrnnv7t/dzhIV9u4LKefFTnOsS/r11X6hhzxO
5ATnX6FCohGYElbIb1cfNxFumFas+5iZt1EYh2I/SfzHXnjXBhGpPeWHGw7C6Y04EilIbssYBj4s
replE+xWLh+v7yH2gu7BrhYGsvhX35iOObkjvCTZoHmLzjWfe/JHp3jUu5e3gTDTkv20wavIRXe4
N6ow1/GW59uDHeDaL3GxG621tBw3rQhbf9n6dQfDm1yhXOak/8ZTBPDbTVReJtCLSQhDH2ZvZPcj
u8whMIOZoE/KIsrdV0Rn/SA9YrfZWn76IW7jSOfBvr66jdGBK22/5Xfd5YFGgqGMe43DCxnejJnB
3TvM16qI6bZxHob2EUjfFf0NNkrvSVfqeo3ifzcK70QkCZCdefZYW/kUHIe4+PCXW3tUxd9h4UUA
bY4ve/KQ8dXrDuxJUAChvu5zZM7AtBMrtR3k+ZlMb7aRJLvzFHjQ1feVsvTLK1qprL9kziEhzZEp
splNAImPLW9M78Nw3cvDfa9gvthwTRsG9O/4ckWbjMttK5T4ve17PqeJBdPwe0ILe+srjcpqdHhC
4bR9g8qa81YQeYXKaG0bsJn8l6LY2pIISUXSSvK2WDBoqCg1/XE4DkTi1V1P7C3gT67Ro/0OjAjI
nuJI/1gsRPZaGWqDKmhCOFFIAgIMtM9tEU5gc3781mpgWTKppRe6v3bgx2UfxfNTSZN+Ku5S7GXr
ftEm7+gPoDhNk+aXgdliMPGhLjtcJ2jCzF/yvM/k9gV/esbtH0XhgyJqa9plCagTnBaNO2HXPV0S
QyjXFnuEdmcXr/5BhnldpaLZI1NMeA+9Q6UFdcOStu6hbOSb25FwJJxl8+2yD2GHqFJsmi/3s+H+
yqlQRaqxmFTNn0iJ7vtft59RpF6rD0vk2Jp9oyAn5yu2gtivt9WwMqlEJk/1lsebWSXyk+GgOE07
M7m1LzxGtQU0SfkRugjdz280lNlgagAjCNojlSVRA8qI/5tBPMsA4orrk6Cc5VXlfDZYbj3s94c/
Ox2ek/aiGKH2JeGh5AZRW4wsvC1jbe1wUXRrjKXkzA2J51o64m4ucGNfPkNQf8U1BgsC5IfUT5vK
ImMM6DLlJ8HRb+ARDItJbhDlvgBNkszfLdmBe+EyOGLxHxYyTcQs4Z3ZR3NWzOJY8UdBlBdBl5BI
aoZ+w+gFznPYBUtXt/3X4pifBVDNpCLk6gmH/ksa8VWpauVrCc+ymlOXjYM09mfU+2ceg97z4gpo
8nuNHh94F7oP29cNj3p90iBb+3PBDew0D9JnfnqWqQK0GxmEwAdAxzL7ZJisqgiATix475sDlLtp
Uffpw35Zvy10z3NbBdnf1r/SqSUdwxpMl9wjS8XACCeqF7H5fRdldjV3rLYJlRrTPUMlo8taUmDP
mTBaFYwg/UV2hu+l/Z1TMOpqHV7uLxSJonjT1IcbNdH+ghNby5MXRmJjEWhQB5fqzHNetT7OYezc
GEAJumlgjan8jTbshH/20gyK2Ti8iyzdOIofwh+VVv3O6ueYTrFSvsyGpKeddGc4zmK7mYECHfkL
VMmF94jkFAE2trVEgs4RBvWMctkFYwRjHC+CkjdoZuxUhDsFA6HOEDq/49jVLRAhHQe45QZ9hyrw
XA+lwH9lsjtZtApSwaAXUWS6uUU7QDV24945MgCHnPkqoduuMF0O/oqKUMqN2pAomclXnIGKSDcI
b/9gd6Rk5QIqsCve9emEdoRQCgHE35sRcSBBl74UUjGyjhqgND9XzI2KXsloBmf+vTbhrxDNMSsj
ji0h94QQRWC3CMy36eyj6t1A8UV/rm4oTGGbJ/wdfowSHUaX1bFDcslQQ+Pu/0tjOED+6scTtqbj
9ndH0TUNL5wikhbaYdacOSz7CWV24Y7aWQvzf27h6X5CRtK2Ruosf/sulGtZnGfnQea5kyUxebqZ
ljuVS1Js7hU1IJyOaNmQ/W2cq5cdCcMSbnNpevJ+0SRC/qTWfbFk4o+fE9BNP6UaPdutf118aygD
jYtDnE0+qxq2fXz8MsyrR05xcN/oTU03fcZrXv22YaIvZnYo0jmSAKOs/jqjZL8fB4Ea2IbdBFfk
rHeGVlWDr9A7Upr3C/sr+qg+IVuY42tATp9xUai+txfVR1xcZxKWpB8TzrpMTQkZ7F7NpnD9a8X1
CVhGBe+FEFeZpu7bXFZ43HcEJrB9ULF6R5q5gcsvU/6/j8rh8a8l00y2X3+ZIg6yjekSzae70+/a
HngPC9p3m1MdMV2gN5+JSCJKRnKyStW5oiLGvQ5b0ltcEyRcRghsMPT5vQF6eYarQHnKWKnm6LhB
CHvXpCg35zPAACQLpazD8Swm6yW1dnZ3CIB4fT9gmxRcj1bQ6jpjG+7A3tZ+H7u7aOfojJ3hPaOY
efKOGCjrsyTuJ2u5JHujMckyiefGfSnHCoURdC+NGk0YfI9ByG8Bh4247I/ZVbR+EOVJTs46OxUb
oGemhQAOQuOKm63xkZFqJaSoyB61mhOUFgB9BKcHaPZVaPNlOXvCTE4qarlyhFRxiz1KcVajqz8v
u3/lBxFHqjFve+BHq/zijp/JMOrd/2CLoDw9o4EWD8Ufb9OND4NG9iIAnpv4p85P8lz0NOW3efTf
hC46vABH8wd/QcjQbdcVKAXiqv9NNXU0Fv2z4fYwSdQ6BORI0hwShDEM42eUtmqkc1ewbgc8HGy5
c9vOQ3SmSbQetQRRYKWFbC5UIuH0AsTf2NPt0oVni64lqyxQWAtEhltlVZDZk1/wmd2nPyV7mvIK
nQpiTyzsC9ASPHDnDcV35ysKyQUx4X4EQkAmR6fxYC5Ad6lzS/XiPfDEhocCrxVyp7rS5nxRizqb
cOSWki4FIYujK1o3zETURHxa4rOCZICkPBIxRMc0gW/7wbZwAEKO+ZTRLhExuwqzinfNdVRbE2Jf
7dlafJNDCt8pIjVA6C2X61bM/Yp95eMVcm62yfPeR7AxoiBynkLMUyvsszD2XHN6e1NK+6x3TwCF
7Iw7Z04r0U0317OvVQd6x712/Uzb3r2erPP96jvXAduCbn22knpoCMJDmHIFN8nmcFJbWBLobmaV
UXYAUJUoeifHdcQLn02XqSeabGogOM0e6KvlzWKwHzK7Xx+hXehHaitO9Dn9fKgAI32RSYgSnvLJ
+HlKb+vOcSnF84v/zDAOD3E1isTesj6M8YRLJxxklkukpTMoY0XnQwC2FhcTRqlPKRAhT8cngT0t
bQ65bhTUqPbKS/gXt8KWBtP/ZK8Rk7xrLdKx2NuPemaQnJvja67pGWDOqlQOJOKb2XAPQnJk+WxB
uHp85ohfSCAZWwCqID5SHAQwX3tjZ//B36Di48ddwcF/hluGk8IPXXt3s1zQZoY6Jszkj/G+4luJ
0Jxv+Ekz0hAoxBV2GuUgv3GwCtgMxzueywnZkFsCNG5WTJV0tcNRImbij4BUTJih8GCqN1Pai/ic
OAVvbmuG4IUnS2diP8FLWz/6NarU/LBJt1obxzo/o4DJ0otzAmAlGu7ikMeatbJVqp2H4NQ0PQPh
ChyaIHTvw4BgwZOF9oOpxYx6g2acJHL0y3FKbxuUo2DUUaL569b5sSSCwB1O89AdC6AZ4B0mZyv8
+QVVjqUsHOGhkP0NxWi3FHViBlGhCoviXEOsRx6LyTP81l8aKFEhhZrImgufXeys95VEbXpywtGj
bk9uEV2fNxxG1sfkFGEjL4bfUtL9tjWJYMnvO6yQaO2oEtNAu1/PIAJOPjYLxFloRm4B7hZ6dnTp
2zPDm1o5Y/8OSeHKZag1nNBR/DiR3rXrBt6mDiVZBYBbhaYqs5ANpaCaqJwPgHbu5AnoFyy0KQkq
EVF7JUk/cie/awuxhQMq8uEjxFQExi8HjZ15NeNyuna+lMcsbCH/PLZ5fTQWwnP1apk26Dc9l6DF
AaSbUkskBKXbSsMPYvTkX8XTaoEUqcjrhAcm6el8sQDTSZadQAHACNfzyyanOARyCBgEzKXXmJMd
TBAdPRxAECkcbW5hB5StPhk3m59er7pwxEuOK3olhsjccUS5hNk7BNlH90MCrWhgSyyHvTaVzj3i
KXrKTWYrClJg98Se+ODFfrduZMf7snKRQllS6Hr+AR5a9CuDUws6X1qAzDzcjQ3EW/BdO+TKREj6
RyZYMvppTm927wdI4GfIqOt9urg8rNgxpf7vWdAaP3e0w/9OY/Dfl17DI+2sdH9ng4sHsRhCSVD6
HNM/GSZ5Xl8g+xZJqsJmUln1mcnjHSYY3jX5e4ewy/xBLyHUi7ZUOtUpUL8Y4f41ULj7uQnb0MRz
ZqzmbC15jIb39WsOIF1v64HKuvJ3ywL0ThKJUFDQbhxmCCmTvdHwfPqfmZEkB4fWACTUft2nBrDB
h692Ylfiz5lU9nGDiKXxzmJBcMLGP9Gwe2vtroMwJJEMHVvoptE2oQtW7DU52NoMlJACjQZ1Zpzj
MG8lcvnsQlqMTt/f54I5aVRepwn5+VwT7O5TLPHt91KTGFXq9acO26h2tEqZ9agrF2Rvo3GlsxKb
Sa3QXoMl3uRsiGbaydCY3AtyFDQEm8XUhOdn71BKpAfr5GG2N5qBv341POal9ZxGrVlyLoZfm38t
L255fQ3e3iAi/kcOnOiARpIHB9qyHM0/L3iI1xGY0bTxxn0zYWQiAdyWxQYwu8NfVBmxPLOpBRsj
Exv+0g3R8dG6Ln8cGbGjg43en8TVNdzam8IcFeHwkqpFPbSJWuVtLi0y2j4zw2ejIoTnQEtqSGVN
fJMqfHt+QHo+kpqbMPfQzaQRZMz9i5PvdCPdX5ARzxNZRqk3/SLncf8ESomue9sR3QwJXFtPY5ao
E7PHxJTx6DCu/y5jRi6c0iYFEf6EWWYNIMdZyHy2UmFOumwb0HdpIV5xN6EpPR6MfFMmO1LSpT7n
Bh3Gtty1+sOyCfvhJF6Fc8uPj3OJZ8rleOZ6EK4gGc9YJZm5rnWVeef+j5GybDFBVvsYYn4nD5Fk
RjNu/zgeik+a35Z6h9/zcdIUUNjGB9lg8Jcx5/OC9zdMZbOnDRBqkaHE05a21ArztESQCiVIfn67
WHekofRLEqnajfFV3/pkL8nPvr2AoldF6kWcEXa9ReKoWIRT2abjBSFLTDa32M/cs90XWxwiKVL/
6REpG7n1QT8obA3qd0771FB8JZYGvBYDHb/O7RtD+gJmokHGdAT16SYWsB7y4JDEct5pcdNWscSz
gLFnFyMI5HVjgzZcAFGik0QOqWEiULFti5gWclygTN+94CPXv3HyufQDWtxGtWIeIfsHqJ/Xpd/s
1UB/ZS5q8Evuxz0sY2Hcy3OgG/ZHf3OBZ8yWMpabrCE3RlDjkiS3R9Win8aHeZs3P8n+3umXdL8P
Ehbup/r6DASGh/r+PUx+0Ibv/BpEiobQcR7vn/29R22GWGL7GBqsStatSougXtefOczfY26mneNu
HyNIe7f1WDgC870tb/Nd8MjQgkikfwYv9Pgr53DdCR7jVgIVjazJ1sGDtJhAJ9L/B4NbrbQVVbX4
2rfONnm1Jra+VrIlyYNM5YehyMCjCxHQGycaDT2s/EsNVNKB7SPWDPWykWk1nBGaM+9A+uDDHLvy
elkp3DGfjUVeN3LWWgkAnowJRR3CenVw3N8c1DVWlt2uvW3heI5EVTOKgVyVFcWvPi8TCX7OjBgT
laZM1kKxxhgPfINryMBrFzvDIpLnbIo8R6Z4LlXjVQ2cFZyaRqfUDNgpTKdTLFV2q/MSOulT2iuv
PlliJ4ecyGBj3A0jYa5fxeG5ZCsD84HEMLgCzwRGhfVVwFBSnHsd21beP+cZxH61goForaNLVF0n
Vh81SlGiNYBIDIIBMVMNMN0ujS88KDkcMkdWsF+EGVpT/jUId/1IimnCdaJ0U6weBHvOHJdrAbtP
0inIj+CbRWAknvvcCmwQHYXKmRh7grWhWH8p0hTXDoQpie9DWsbfDUvG0h9Vreu5NYtCebLOfeUm
AMkZqg9S329MWBFZxpMueaWrYtmWp4FuTtqxFOoyYjYlIX160UZ3NhEMdMrCoksTo9TGDWZwkp7A
8A3xyXNXFYcCyT9QF5vnxIbeItU9FKUP0AzTFr5Yg5KWOX6isCHPP3dO5MHEU6qCPdbl9FxwUVQx
VxLRhw+1fLPI8/hQUZi6wmgrORzJp/viVx5qGTq0F7J7NnEs3y7QMW/TCJm6cAohMMkvHtLGURId
RjB7ZuHhfvtyUMFSV+aX40BT00FJWANEzgCeBzTF8+1lq2kfv9WTHh9HLxh0oCTUBTfva9/62N1w
MqRfbA3JxFUrfmkRSPnROOJTy+cm0vS8RImZWpqdvUPn3MpiERupDiQKt+fOL4MOlGeoAjPPG7be
3XFc+4eaQa5Ye6H889DcOES0uVNM7+JMujfV1KOmF7JdbCFSJnPYJSy7dwaoDqiuzHRFhw+RRC7c
rtlPu8olOAywfGUYo00LoX+sXRm3bjEvxNjgQgeJUtGgDBERFaL9aS7u/jZ9V/pR72u+IaYy+9D5
FakT7Aa/mlhzR5/0MOYET3G6M2ZYTmrhWPVfvJAX/HBSqymGRmQ2vHEXTnBnvIM/64L3PG5fSXiz
ESrf8CqV9PwbkRSjWhA7miRCpxgPe9EZxHBYUHl5GQ/JYHh5K6OEe808phdiiZMIowERdWm79Nk9
7tGV2sOifimbSLVAOFXOrVsaUEKkSODt5P4pU0HQtgDDlvI9KTcV1fGy/S0yjwujgITKtf0fHRMz
Btk5x4Z0YVH4qGAlE1NqEV+AIjU+/RLviNClsmIPvZ2KB9606eJLYo2stRgIEEvtojR9pKm41g/M
LXMGrLQnTKFVhwA5QGX3yOZgUEpsKAT/tuptPXyZz+aOunw4Kib6EFC1I/tVGhNzUCo9Wo3erDV1
V09MCUfqaNmJZnwsTST9ZhXYkVg4KoJ3wMnYB6KGXUvPTuLYNWOC/x32RWRwwyRMT4x7XKXcJhGV
k85zOON7RsNWC9CnmrVybIYSRErpfDQzDQ9JcfjbS+rV4QWT8uJrTT7dU9/LJ4gzdV4Zxyj+saPz
XStDpY5hooBRjU7nrowCWanC7Ql1tWv0TAux57SKWyndPQTdg9+wa8tjFkqNuxCBbQTgSSMbMxIS
hhNkHSPYGRsg3Ty8hOOetvZyA6Fu5wPMoKibdlO1jKiOEl0SPTG3wgAZNVmPlc4/o4ioYXk0JfT+
gyciLzHJFRPj8tHS10jey5lig9X++s6D1xOfYy55TQPrzlGh0lOitQVqcjbN7zLZFmwKYftnr89f
Wh+Q2uHL4YPzjPpQZPb5LgXYeSWT3UsrMrBEttGsCrYmzwF49rEhoD895P4oXrevbWzTmzD2MOcX
7zlpXEADCN+Y9nUwqwO+eRAvxeLTKJwOvaXE3jhRfjoKdayKX42SLESyZhSE3+YqOH5hpYSKn4ey
OWY7h2k5rM10MUy6+dWY1snPze0b/dVx9ZFdn4fJrDM0dAci9oRxhKy7Tpy1//SgMqF2TVjDzJcg
BW1tGuTNyP56md7op3TtA5+ok+GzraCEDKO2RjGFFJ93WplTaUIVptWy1OQRvmgaQVtxIZMIm4pG
SJZMvk6Kbqencu9GDrS9d0ppajBw+F/kDrsNOvyuiGjJXkmjmGfRlGpt9rhdNdgnR9KMSG7KRsNo
q1dwaZ7vNEY5P+9Y9T7OsSPJLbLYhr6s6Bpp3ul3vMkvFeNh9WWBu5YIef8U5SXtAn+n77bimIjh
MqV1vfhQu6+N1mGYiGOz7bwsWtG7Gx01bdAjviDtxJOorBf8uPSuGpueDNXJtePG+GS1ooiLO6of
rBSmOX5SZS0liPB5xSMgt4/HNHuMaZo1yq9YBsV/HF91ac3lKZ62/UtQms9Xjj3sqG4qHJPJ7lE2
He41Hr81MjBEFW7IjaNaVLqLIFspjsoDjowjbsh60OVUyYNUQ8GrlNq6G4k46dfvCkVz+jaKIdjv
jR2K0OQeOTSfo1MtyBLrenzGnvzhjoKSgiSYZwakdp2AHRlSq4ugImNj9FikGAVkBh4tzdzgx0H7
9+EPwSnfy6DBSOfPrsp1TIIIjYtt0JXBs2caN9PcMpJBJI4n/UxbdIDfkUBqA3X6pICK/PXFi7rl
PQYd+qAOFHj5RHimGAxIeJc/YHOgkzcnAOMxbdRBMApjP7DXA+dsLGQRyzCaW7TL3FeJWhU8EeTL
DQx9l14DSwfI19wVQaaSpqHZ/Eg82w/0qkinN2NEAHL4kT9fLv3OjkBbRl5DLr0mdN8fI4yEvU+U
V3RaFQ9c9yeB8a+Czr0hbQ26vhcvT9NG7OWtvdkkcCzMSW1kbhuv1Ybntd+sKbTRgUQ+1UoXtOrb
CWYyezEREth9tWjTmLHe6PqtGJ6XroIESbDYyg9mLrGPcXpzwEo8K1mZEikbluXbq+wKX4kV0lKj
PRf91c1C3Cxli8izAvwfo8fjnFZXrK1Usv8iwxJbp1qfPsVMiuBXoklACBUwvDA3CKHTaKX1EgIh
HGQbE19MEUDqvZ8hMo9hlK+mRe1O4bvx99u9Y4o82JI5NZ42iZytoOyXRt0Na0OxPT2XZ4sVh8E0
7V5xmXZ/MvkOI450mYEGPbezUE8HW5VKZWoFZlt17XKpMwayo/Jx2tVZg91aeNF2M+1736Pqegi9
kkQDgFlFgXO8S5QP/w2/vdcQfiHR/KDszyDNnqY2XTbjb8doMJnEPohHNObWAzTLRiV9HSKYmAMA
nfU6xANGKa31XQfmzrl32atBbTGZxgGQ2JRLj6WK5mk/uhj2cZfWUuEAAhox3alIzt9eokzjIbuY
RTtrt14q7e1lVyNWmsDq0qesZZy35sR7FKmR4+mSnWnwW3EEUx/iqza5q7kju/jHbSVJItRygMBY
tcgmDN4SD4mhSkflxPAiPnSsZUC3rfXgI0UE6sI6cRjQ8yse58xEuxUuGnmg+LTA3fQHvExT3VQX
C/qzC6dHXyKOS9etYvGaMfzoJe2MxN33Ele0ji3Fd+bnbMsATt1Tl2eXdTkpT+cYiFP+VPgx6xJG
vod713d8XpWbMr9Gq2/681GzA1f0f3nigBUtOYkXgWSvpSvMiKN8HZr2MRxe19GS/1UFjjy5OOkb
lUMqJC8P/Gm40xg8f3Ml4Pzx1ngjtaUgUMC4EIB8DsYaP8iH1ZGgJihyIrub21YD6C016DlBHjDa
cI99+xL2It2EIEibT9bz7pItQ1H7kilzH+gXduByO/GUK3gn0RY+dMgE2JhY0k2eorDwrC5DvcZK
Tbn803u3sPCKnRXmoGM8duRNgPqZiojaMnR4tyV1W17KstcTFMbH2rKgjRdPwy4p1ebbfuMM/qvx
r+jLhNnfv7/4F9cQddxL9Sd3CKdKgRuKhVYz+qLfJzasCq3FujXFajZoWLrFWvc6UT5vXxFD4+Aa
k1vGkWXkTqIDfTf07EW1CURN6d61F/p753LjyWr9qVwzFMVSckSzd6PgX8TLPgFH74o7GY1jYYAt
tXB4oSm8Z+BvV3YZCIYjFmqiTkunZpkWZRJZrDyg0UsAjqtR/7l40ucp4hDOw+vvhNhdfG+nWI6q
ZdhbbQ4ZixhTotbW19gbCd27FaXcIChL37DxcgRYD/YRYhrEGjcCNgyrX3qhpSIXjqbulJceHOeY
ICKpocsjREtJYmGM42+8TJlx+j+gyJZtz5M+MmBXgozMmINumt7+vene7pYh6FprHvrCNKVsmvZk
uHgum/FdZpC9/QQL/13O/jHKc46q2CfSSxgnIVIteSo7bLPNxgIQXsrSTg2BQgUIVI4kOIf+cOgd
2OTAmVySTff4abVLFIkW9HuAE8hHMXqzAKgFV+4ud5LMtaLvYcwIk1Lglri88RGAj2/rlLgNqKsh
wqQWzu/LsfQdZJzr/V8m/X/3Po0eldQ8rpsD25OtScY2kJTfs9yTQNcxxUqI8pZZqbkPprb01ZMe
ZgKF1/hkERZkSEVcQeJlDVoCwyw7dug8EgGZNsDrSBhmU6WS3NTRHvP3+PxpVBku6ynoLtllxwi6
BOK9O9LeNXdAMmIbT1H20UQhmbQU10nusDk3w21oMLXvU+u6/OFxuP/X3f9uUQQIf6Jdmjniil06
isAFt9hWTJUHrgl92miLAsNzMMOXX4x+8NcUeYn/9Fcj0TsEUfR5ezQfWUhDNSP37o2GAFvlOKtS
WoJsDO/1GT6gfptAVRh8BZK3o987NDM2M/1AM3xeV0bfgMeP3W+xgleo8wVsLAFBpS02F/AfjJYo
zkaxWnAcGOrHfIRQq9IkhgStNAhZHv7YQW+GVxEb20t+J74zd2eiSY1JqkMgvHvRpsvQGCo65Jb8
QrzbzU8CH+eyDloSJGMeE8eVbTzXhUGeQrXRM7AHfRJC/Mqs8fAkz3e3AKS7hOS6mv1hliOIGplT
eFJZ7MI/TQdgkRRVF8DZbuSigkZ/C7f005j1AOZzrVPvbwbH7GYBRR55eDzWd15Tqbl2U6NZkDIw
ZDk7V7XE8K9uLPUleJDexNSmUhn9RKgHeFdshqB2n/9O1CK9UZQOCvK+lgA47UaHmvsfvMPO8Un4
Iyx/AoLWzFEpyt+ts31w/XE0WWGwxEAdFDLNAvuls4OCRo3u/+oMqT5RRvBGsPTVElERt0y9SNkE
u/HDhkvy4iGTGKn/aBy3DIzjrFFnyYtNMjSi8f4Hun/sglMv47ayjP6g6XlbcBaWv+rQ0jX1PIOt
yOv9tO978bvo379j518fQZGeOf5hoxR0Tm3UlesG0aC4NHfhtwVukRZu6EoqJSC52JlXQvVhZ5UT
RLOeEbWGPBkbExgybHeplEG2U1X3wlECYf1yKZfP6mCVCBMNfFjn7XVN98MUifRBKf6sQAMs4H8D
USfW8GCxiDttLEA3mgXqUqIrmDpGft8+svV93JUMd1W0VOm0i8Sfp/pKFv3Bx0br9vgfNe+OkPNw
TdGdjdJUceQ0gAXQonYoTgOu7Py+DamqTDlO3SYFawyERAsliYK6fUNICk+zpK+z1HnLhbD/WgZ5
9fvFm6aXdbQFcHt5GIhkNtSyhg/8qauDMuJWOLsBGp/7xvpuPq2F9LKikT0emdnDRyt3TPT2HMh7
S5BoXExqCjzRcm+Aqa8tHeg6gVNRcehle5mi49QgSLHqeQUuEXXbBBaM9vv+wpkaJX/rWzUUCN16
Caoxh5P8PjBbxmmalJvmxbZxBV3pbv/HgjxUCWZGTm+54FWdd8OcivnC7K1z1h29WTl1jwi4lmF1
QtsSRakJ5tDQlON83P8b7PrhqwBSVjah0plu4GElPO2YLNU9I8Cz6xw/CVqEAcWiDZ9V0us7Qpuy
mbWyR+gWuNISf8/yZ77CLrDWUrLg8AeDiw4uR1Hqbj3TBIlu5E8FpWqKNej2TuZNXVQFk41a5vQ1
O1FgpB78iybGhbYsp6O3myoO1WW5SPwPDUKfDF7FN5X+uAiIa9hk30sr8csqBK8jBrOHXIKGDWEV
wJyTjkOvjZpjswZ66j37XfCsYcF8eogKvQmGmKlCRM1phSBsRAtBTF6Pvv8DwiRkJvLA2w3S6Mun
og3AylYf9zkDaMjfeZLWjKc6yPzC78lJm0e1Hexc8xPf10DWpNtKJpZelpUqxDgkJPXspV3OEpIC
XYy31pwzCet5vOEe+OTp8GNO4+/9naFmOY7YAyDlLKJ3cHd5ZQGPsb7eW1hSkK6BQwyeFruhZusv
/9Ur0lNXz3VkYYMYUNVJgebP/wbZatQ9NDgoCYnVpjtsgPWZchWXx+pGRHtjtIhOlRLy7PJiL6ZS
/3bZLOzqP7bt7k7lWJLgYdZtsJrHlz5cKbNCNELtwvVeE2N3lm1lb1k4GA+04EihbKqV707e8xoK
9Ul73SK+vF+cwixtKu/I26GddN6RyvCyi6iL87pfZBKtHGNVZILlK44HR7YZQJz/w2FUZ9l3rDtS
m6Yjf6M/NM5YpaQ06vh49HuG15aBj7mXLyS7T+mCI8O9Td2AW1A6MkmU5TpNXGVHXYxBigTF7VdJ
Vy5tVgDKrKN2fCt/tb0Bz0I+m8nvazJYOlpCB7/06HrqcrZi6dY7HezreTAz6L/IuyUGmy+j/3OX
kIBnZcjiRNR2lSXlZ30/QnjoBxxhux/3kjzwsNztCdvgtuXLVuEBruiZU8wdfUp8CE6fkQqvLRqd
K/o1aomgkBsRyHd4GHDNjV12Nhg0hczYqzZE1Xc+VN5PGPnQPoSWFyAIZip0x9cGYNQH24c6ni9R
KKBjlh1SRLf5Ki/Fih1wh/np+cVxNL8p6Sn6t1vRMqy3fyO2RB0TS3YLm6RzZ29UQhC2lViL7o5V
6fZ9c5yV+VYUwQWSpLyBE1XXbfsytaBGv8Uq9yXMm8ZYZ5+RQxdc/tQkFDtGluM8wxIIamZsK/4g
jq7mZMrme9zFetKh1a9UNc9KgzGgsmZhxUkK1QLfWv+KAIT1KOxpkR59LjoLlMj/z9q7Gxm1tkhu
B0PAQknXePYaVwgJ3fhsli1h6z6oCNNJTiiV5fQbtoUaADoICDZqp2VWs07CMjBnQyBUl+1vyV0I
Tx6BtY/8BKd0bMEtbtyW+OdGV7J9AW0dTr3u9wysIeFm0i3snaR/MomgDl926vh5HVWRApgOaQXq
lrcX2YmOTatw/eimilsQzH8MlXW8mmdv7B5YDK/nEkoHL3tIFiEAKgtMavwPkEH8NsG2U8+M74QE
NlcuQoEmmzxiq5CUpIYioEkLETQsCWvG1kviFHZXImB04KNpGWER/TlBnOHB08So3bP2TDcBp85k
0w3i9Aquww+C05gw/okAZdO2/mMYqt4DxcTfKnzgVoMmTZaoUniU9QikQ6gnFqYT919DQ/hikcDy
uFPMRAmzmfSjk8OEDZp31bj8cBq2evy+fksyYv0KYahuaDOyzW8QMdJxYnWnvp2RgjBgpIO/0frp
CDQzLRCsSPgR7SMHRrtJI3VohKzyDMnk3Gkiwas1gEPmNCLAGzwnCq816nOOVdOQKVOCmJTbfmTc
cR3binvr2+HQ1ZvGuH7/QDap9uQQK0rODjATrsqyfVvdwYmWqYpVyJWtYKo6kMFoM+j5M43v1j7K
0I77eSRKhh3SySfJ2m0k40w45trsISLWyvY6l/Qx6hY3ouODlexk8QeMes/YUSC3NYWUsjEI4b+5
CnLoc1I82xyt3TziLR43pfwFFMzrkU8e/m2ixoTk6NDlHI88hrzum7cFwKvcoKE3/Q7NQqskymsr
7invA8j7k2nfifF6ltxp5tuzge4WmWVT5xrF74v6EaORz04yBP0clA3loOtS+HfxDPDSIQhsPgRe
0E7ZwsQQhn1ybvZmVoKDPnR/MP0Jc8AMXDkv+Sb8I5PQzadJ1Gb4zhtjnEOA+cKyQ047uQQWAHxD
XtGlSFUniEpJ2TeXZ+ivjLc0QIXhTcjlnlKSEcE/q0TzOOsbwYPYtx+47I2cwVXI0+knsrsXvjI2
atRbbvILUsBeBhs4QddbEAQ2Jkq8SZzUa61beWverHLGm7ReV/+5qKQgSo5zAZlJoNcBsTo4AslH
Vf7ZrX4MSUVlw2mOXIMCSZiUZofziJCg8RNr9gNDYjtwaJfaI/mdvkQUuT2mk0vHltIspA2cN9M4
BBf9jf3/dFV4Ml9iKY4NRZzAM27FiBtSHr4A4DEtrT6suQX3M/z7/KAAo49N6B44kTwdnvALKwWp
9beOx26E+irul/HS8RQLyfqaGQuMQpAG8kBRZmRdaL5yPaaMjAdNYBDEPfbwbdieDyRI6ouPW5Si
tPOrc7xKfswvhLIowuO1o9UObE3gzi1gQQMKCK8ZqoatMWa9ONmTMJNcb1cbvC6QxDlhZE8ZfioF
zdsgWGwVCXsoxmnu1M75nG8ybaTZ2r5uuv3uKhJuLml90fYe5udkOyE5asxLij/80hud9wZTzEHH
pTFTO0VQ/uEW0MrfffTZJMJLR3/ch5dMJy/dz0sPdWldbCTTNkdCN4to7o8jBVHknPSPsFXzMkgU
khrxGALcS7iA/qdMnPZPOMyt0nYzr5dzPaDvy1DSSFap2q8c06nS893hQ0OwxDLB9s3D4jb1f27d
pYXEgXvCm/8ZBRb4diJzqku8eQTWXfBuviL9nND0gpUNnFEdE5yaCsRsIrq9jgXCug5nyprvYO36
2CTbU4kKOyKg/aOdnNeNbjdW/632WsNfc7bVOCrTtxRv/0Q6Tf3mykwIDkFP5PDk4WTMpKBcDH2z
RTJ/rUL19FxlvAPxD1ilrjSaGPgsX/J8wDYJFkz3YBUXa8uLL26Mp+V4kPdnldC7JtfWt8eOA/fA
sFFe4T1+UsU0KMWyfZ139vdYTm173ZDtakkrmzK5RgBALU1XCcgPMRr87LC+Z7OKSGtnZ8zDGmR5
/LBHa9a+C3bI5pyGTxfxxfjv0bZ3fY9WIhhaRA7DbY0CslNasWbyf2cgwIKBrnskT3ZbLmXaDNll
Syc48aHBrKJ8KnCsED6COlhq1SWH9kH7Te9wmpQ75WmEpI9EvvTCqyA3YzDztUxnpeAUUJFtgnJL
goGJZWYJnqEjtrLsvw8MN+5YbLF4rEHG0km9avRjo99CqbnbgkBFSunkSeILBVdzRD/475A/63Qa
vQKqobmx3el/1Cfo1/DOethfB0MCZ6Aff+HSAjnSyGGd1o1aK3FPsZQdJ0HwS4yg2qmBbA9VSKzT
ntRgdYDot/CIw3dJTo/8xe1H1uIGUuRcMfKf6h5kz0b65vjPiRMpl2dmo/28OYKKbU6l0k1ISKGq
3eJ95CIcdiuUDU/cajkljKznCEDEzvXTuD3aXS13uK58pA6JJBSf2Y4U0EwRZcwEQGcetdqorEZj
h6BY288jPVclGtczWShcaJQUtWxKOUqEYCRpjf4Jj9k6iv/YI4s00Yb/dzDKyGwy2hJPInt2wnlE
jK9Yjl9B31oO8vEYAGnXt/jcnW0vN0NiMFMfexFaCNPXyI6zoPoqYBXZKgBSvMuk1JhiwxI+z1nL
5ZaTV5e6kppbmWNtYjVVf4Ar9qEroxXog+5aL/jnkv596C2BGH0xRLwe0aE+VS0RKrG7pqGiMGV0
+K4wLCcDQt6MwhNTaam1oFtdnPmyiLUX4qBXjHPUb7uiynywTyp/prwh/1qh3aSq2o2WucBp0nL8
eTqPBOoG42czc6/+MlhE1MWM2LVjaCCfDcESQ5MQyHvZc+FEKxR8iDgAo+JN/5+ZAs/XMg2x9XzI
Q5lUK8npvBqN34Qn66HpDDPZrkRBAsi7qoIilatjbn3SC9gNkg5GzcDEVSlhzIdWN5tst9exCtPq
OoOrDWrioqhJn96ZWqkg0DWXBNca0xKkpEGNuCHQZfU9iJUqMqe9MicgW+2xDJIAjcEmaQ5pqYYq
9V7dSBzv5Bc2RXxekQ+J6hrsOMnnW3ABZyoH/sc+bmaptLb299bm5c6z5ICnzmDlM/R5xSFh7wX5
pc3gtQWoEtUt1J2Scv0wxqFcq1HGfW/vSVLGXHuKzGo55Q10wP5fCMwbBLoB0y6oGHjkclMiYJvl
xTzJRYVgvrgRXtLNZgpQtP2mTUFVpssoXapipdmbfJVb4KWFcy58EVimlL7HsCzg7k52jP5bOnxD
Aq+zFKK/RxWpN8/KqOzFoJDv1EpaaGzTXjJsh4Bx9wrg1+oqkLgLJFE9MfZLqLpfpLtE2iEZ9CJM
CFyINmgerpfHxFLxyiHlJMAaiPiMSsIrSBGjK0XFLnyj0e54R1rR2KAeVQpqx10yPVyOWuYhxRTW
whSMlN89XDWKsMpPrDNzT/9Wy77B5y5tPltwuZ6ekv9ACh75a9BPc4VnitLWVhWenoS6tOeIXep1
2vFmxhdDDnim2dJtU2RoqMKRZlWeiG5m4Cl4Ll+UyF3Qj1vwdIrsbDbi8wKvzXXLRgLRfKo60Cu3
S3a8QXbtiQYzVr2mfrV4H3yVS0rRB04kxv7lNXeh38bR6YGN+TfpffRBxlot/ceHqL1o9UeuH1/t
i9WuWBvwexhPo59c5jht25irT25khX1BRbVdDFtqW5ty9rYnNvWaz1qIIa1IhtWZMBKOP7BQ502w
LgnPUh5oPHT+VzwkFy9/gjeaEv+c8+2GM1N9abS6BehoFD4ysCPXRo9eDBXeWRVRQTfgdxhELQy2
vjAQN6atZSK9jrg+BOACfFDpMYRlg6s8gw4zhNY70cNNxagr9bBLcXs21VCTyJ9yxH+vf6KqtLgD
pcXFzlARulSRi4/FHeWaRebK/TWHIaShc6q9V0pqvabBqBIzKa1S6RvKEXlh0kjQakkUYKZO11KU
tGBWrl3eNGsmaEgXGTNbeNhLs3i1S9Us2k5VyCHw3PO4ms2vJxfHWPP2iPmietrHlfvDFcQeC6p2
QH+VkKKSRWOacntnVcikku9mRS0BMfGd7V8r9Y4mGNcYNIXLCpV6GyaHSBnkedZD5CAdztj0UZCa
uiplf7taYnOeowe7fdvq2gS2qKEhPjLcXuXuDDl0tjtAsANYDmVGw+xp8b+cKiG9KpbldMrfyFnr
GkfD4H7b/GbTu/3eE8G6yrJDUjKCmSHyvd7H+wHbDX0pv7RDoYEsx0LRwRY8nm+QP5JLXyJQQmCg
VzElXGjtiMCijDdarS9GIotFohWK8Bg3Pfz7FP4cO9n+GeU3FOsgL6h0LszadFhfpAXq07K6Oaqx
UsvaxPEIsnQ5LCmjn5a74J0rlBeOSYBfrbvi1xaDoZkUiwqhtdkYITL/XxB0Ug9u4Fu2mq4ThyDm
UqwSFW1Q2+91zMjTjlTSbwJuPe0WLR/7YA6OWZFdd+SejI3qbe2C01YPQPaE95kTNPZMIiiF0axm
yG0Fc+cWv8qKhSHLve0+49KC5NAsJag94pPjOZOLt5i/DkqqVfEHYYpHl+64Q+zEFZvzqOUWuEaQ
xRiqXnspIQxRlwOLOxgeliUzIuoaEicxdLUrrLYQO/7eIz++OFoAHitjpWZ5AL/siJYlTrYOXCdr
mgc6uohp+hWFRJ1OFUfoQP+qFPrDHeDzS4mKUU40JFEjTmIeD2RD1YiUY7z9QtQeDLh7oWysCAJy
Ltm9qk6qxtTahSFG6V8++j0z83KaMHoGrMD0Bmiu9Do41LO6vk+NmWL9SV2clbPTgvCjT62fxvtG
yQ+K/Le/WJh2kuNRhfxFK/npNfSyGghKGvxuA9rlhvhu57wCVm+LfD+ZtPQ9ea84PXaNFswVtbAs
frgWShgGbkPuQXzJ7zli4nxpwcw5Vy7EPoJEIJftvgW5SKW9PTjZ1J8uQgfa91xH0W2JEeHF8ksf
fNP+ipkCFPDeOsJyLPNHhoOi97MhrN8efXB23916+t7p3faJ+lh6xHp37+CKfCn0wKYExgO+23e0
OXjYT9b7IvB0Q6gQ0qQXluJtzqHxnBK8qNdy2ACsSkBmT3stgUoxW2y3xc7kWDC7zhMnwrf+ZQwA
woxXF+CRAowmeCPODtE3w/Nh7GyqY91lY1idGr2gcCazCtiRVxrGEVk5qaBAI6eGudgXzGLqkSHa
wRhBrHVxZgFPERy7VpaKhG4bwt3s98sCMbvfgp2Ub7FE/QL39ZSwgNTiu6iXsBhPhG8ywJx5qvcI
8RnLJ1P723DH0sBrI8oJ/mfdA3xDYDjJuoFpHoqtmvIB5U6gY4je6ifnFQcRrfmTXBlJijXU3I2w
gYw9ibw24Jc0WL5KNzZOh8N7xmPQt/SzYPZ84QvgnsaeHAmircy7DnYf+8E9gpMBVFSdz7cZF/O3
onab7iE4s5rMiCvnp1E/t/1KI5yXlpd2GSqFrVW3WU30y8unp0uBVKPs81CfalKg2UbHgppMmEE7
SosADeX/qyEEzgJ7rhmfsxSaRldsA8VIqYn6gch/tRp1Uhnkx+JAoj6/OQhDYmD52HMwBWiLo5qd
umjNXnFxz6M7Ot1YXwOuTHOp08bPN7W1C9HBv5Fb/+bpW24MP3ZPsFvyIp8VntAG3IW/A2U7JkmY
yVjzLy3JYbDB6G9XafKxb38jbVjTbkWY9/0HFggBiLcexotlmRwi18sLtCjsQ+g743AmI9guABT1
jZzdAZz2Ggiel+sMEWBF64EpSotqOjW6gRXBgtltznBxMhoZa2ByOUL+tVAnUmCKmdABTSJY0+cd
PUM11zoGTCDaOHluGJUxH7CTinCfRulPzmnvLHxotDgg2OALzkVwyq93Vd2qshnEKRM2trX6RfHs
SXn93D8om88n8Lr6SJDi7tZziRov5yso9jXyuFrOylbB8UxYPvmlr3zJrUuMI4Q4uB9D8QU/TLHQ
eHE6fxWk1vgytBT5Z+2Fjvr5GsC1mwxN+5DbWjhmXKDfxBwkcvWZnWsBIedz5WEVo0D21wOEP+aZ
01oecAYYmhg+oRZx72Rkc9kB5ZV99l8JHV63GULcQXHYuG4uBnaJGM+0GQt7rPwW2CNBWtvsrPWD
iojaoSjleBAm3MZfnzGoyNwFQ1RHpXQUUrt1ncljU2nDaeUeQuR0B+WY5jsbSnQIYQRLGINYHNiq
+QyvwjYVfatggE4D6cGFBZgcTPHUeKQEt+9fY4iCuqiv27VQVuPe0LYCaEemygj4N3MALtWEs7KN
iBE+uQeSeUfLwELyHJDYGmBA+MpPCKZADVkDueNa7ODSr2EjoonmUP7kxGEMmUHgViAY0AdGO8lN
0baAG4W43Ln2oSqh2p9WEltNBKMqMxmiZIeIQQmudtT1PukDiX/rm1FIDM6r7xE1dqUoJSCuvKP8
tqiPbEGfGdWgFpY6PkPaf112v1tZSGuUlED7kplsGIX0PiS+wgM05/CaBr/QoxjOFfvX1Bkq0ViS
JaQyYDhI/A3XgKskBrdAwz579M8N0j+7CZAUEc49M/MnNA+Wzrv0x0Lc7jIbK8CUdEtwS8aKX0JD
5Ai9BcMzSSHxrFuU794MeOJrcIg89wCM1aNkwepXmFNlmHyO/hs5TIXnk9g5516FbPxi6mRln28i
qxZxHcRXGWyULNwf211H0ODdFLCygE0cD3a1h6HgbortKUSHJqOTPCPih/qEUWK3PE2uZW80ugWE
rYybY8fpgYt44z7lAbjm4FEpK6t6Mk+nlhi4A2i1jz2pvy5IBtD8qEfyo1h+epAYNBAI5yLQgBhQ
iuaWHHQrujNU74p4oH3gJkZ0wYpbJfeURKDOHb1H8DcLLKw4AzTfoqD6pH2Xeq9sP/YHSIoprkI1
+aMqgc5KjQwkScvBb4bPU55qucheMdVDlwUPvNmb6kpAEKK0hoY6ND6BH+zcei3q9vCMK/9ma4VG
0QBBT583CG7poQ3fd58u7k0R1DuciRz1n2AJyH6FijBEiPbvm/+YX6v1JnqV/zCJcKZ7CPyWTjWJ
Ern73doN2RNy4Rxpy45Nwnt284FowNaKlFxAu8v2C1Er7PUKsSzF6e+FGnHJxtYLgXWsj5re8Yn/
lyVm9I06CTBOYzEC4sxvMv37GoBeActB8wBZcQr17l0PHKHvgJeHpwFGWlOCEx3788iJwqkyiR2G
fx7jp3ZPIXuySXTPOkkTS4etD7Jf5vb8tgNf6rkYUGeUElQAA0QEHWhWMbqM7MgJfKjZZkCrYcsx
9HW4sTl2uf7M1zLtPmmofhKTTvwY31ZqrQjapMZC61OSlEIKa/TTgo9tyXqBrtE6ifKQqWek3HCo
5YiEnj4AzGrwfy644leo9/ynVTmgD+1XHT7AynUou3bMWl26Q2wF6k9RZKAoy5CwTwxpXeA4qFCe
9Wvzxmg+/Czkok2M+LbrfDmvxCBywFbYle9cIHeGBRosiHAjDWBlz95z8LsShpLkeTKynTbK18ta
Koh7YRrMdIL+LliDvV3ip9A4qpnNcf0fQ9yNLGwb8vdRL2fFT1IiqWt3+qMpSbF00jEHnl89Re0P
NO/oubpVzfpH0/FtgGok1v3wpL1920v2313YcmfH6Bl0kjEw/WwWUgmCn9V6ARwJE4wa26DKYkg6
gjoLpWXrTHDUuQl+bMnJSl3llGs0d0gLzoEmwEV0En31zwc9NkGz38GWTD0JNIEa4tFmy/x3q8IE
rscy33+i89jE9XvlMCA4Zvrekk5TlbDaer4yfCEeZBIKnsFaqjz9SwcUkJbmQfWU1X9uN99lxfhP
3MAx/SSpzSN4J848L2ZVDaHIe/GkakCxNJJR+aR3yonFepWlfGssUbhRjGT3vgql1vx2lW9pkftc
04XrGZQlu77YliSsPserJXV/GGZmq3ZXi62sakeJsGtvEBMsqIkOpBWAO/J9TNW6IUDEu9ZT4t71
H4GqqRz0csYt/QEP9UxjFXoVhjT0R+Wn3hbxwfm054yQblXJg5cO2syU9DxYYqEBxeQlqEb0t1RV
8GabG4FpGmkkZ/ujds5N1S1+N1ziQp7g81YRF51XkKg+CDI3JvsprJnbsW8AVBcZrXpXpQXQFbum
/E3ANwYzxkKA7LksVn3L8V5ZBvzey0lqJxPoy9wejQJ20yKWeK9/Ga16bLYZoM98QBJSYsjO9kyi
+i3yda95SnAMCjhL4+D9bNM4mgJvLOosu3ZkEc58K9puyzS+xeQPGkoOzv1+iI+4ExdlzeZWy9WT
2pU/GDWjbcY6XMux82dVA5JmPhTFwi1Ac8G/yi/AqNTeJbuCw1EyRdCMpkBxNlrepTRJu/jtcat5
jAVUMp5hM0mtoAm0l9N+VPbnWkVJmoDjaYfIdNbjs4d09bycP63g381SkobWE2w+omhfjtfCjbbT
+Gm5CUOc94cQuSe1X3poEx4zvKSak+vUcdgFbXTicQ372hi6zdt0frALflrwp1FgFOQrcWjAKjpH
WLQ+pSE9tAtHQTFSqUdALW+JzYuVgIyD52whJ6YEsPHJlVp8DfSJVMul8CvUiECgaQ3EYiE90bX3
q4csiOU9lllUj2p8yJUia+yMt12BQdE5sTEahByd81mchq3ifWMUrhRXs905FzGzP/hirFe93vnT
H5K4J8XpV03PBHgrD1feNc8lNpCN461PnHG+EMldb+re1BEpXC3aPbWKPY8EZchjEs1BWsPEHTOv
bClYZ/ws3U2/97vHS00nXuF5yqo790BENyIvyH6essbaBW1pF6vnnhsyvQML9DqNzbJ/xvab+FzK
RwKrEjb04hR2MA7elG78a6kU652lbw1Mv2od7AMbJ/2rSScbHPij42DgT+aNq10+Y7D1EgpvYpqr
voiuSp3Ng4oNunwa7ZXP42YKBGU+TmKEKBE81m1/tXLJpP8eIOuWRsbmb++cNjwj0KC+YcXRGWX0
s+NPTLbaRHMQEcsQ8nR60cTo3U/Rym/m2g0Oa+JShbTlKga80R9JZIsv6oeTlI6zX+NBgSUH/Ukk
o5fyJUTQHhosH4diVbJ7ntNqJZcoz1rpeqaO+H0act8mnkVCX/6Edxo3HuILXZKQZyHwxGr32Qzm
Baz4D0DWH8QlER6l2CaVF99IE/XKyQ3yI2O9FrZWvFiWHEjZxNocshHYC+QBTLnQggSZJmBu++i9
pyfd+oK2NONDXR5ZqgiqnlOaM3UdnijnX+ZYD30ZKKT3GNBrZFz1UrtWS9u53nKWYwV+v5Kd2T62
rwhfK+v71jz59/4HuDv0PKplwN/NAgqH0Q2eiELFFgEA0Ysh1rA9KsxyKRq9dvTGaNoup2s6sRu8
9VRryb6cutvWcVYgPTro/Su9Rn1/rtN7W2E2u6swbmyXq/0svSRTWNs/SJoTtI9d50Kq83dDdB2W
ECVZ49f2t9fSVfU5TPrsZG5FDVyM2qW7hjiUYUNLJNBQQSHzusYZ8xlCmRiwk5DDC/SWxklvrdFh
lN+v4bLyKXluiTvxT7VqR5ZltgTHlkCNyW7Iw2LJ3v/IvjNox1VWUpvxgZjsk+KbP2BrEM9ucDdu
q2TIvOBsJ95fJJRPYfuusw0gR65QcwOLuxu2lFtGxTZG9ME6cZJS9xSP+vmsXbZoAsLKNCIXCFjg
ImmrFdOicGLgl4/+aFSVwek4E55OxkKudn141PSc/jsGBYoqSxMluevWIoqSP82V65Zxu/emYIrm
USnObz2x7W496/thUGgmBrWtl6UqiU5j+Ln9raY+IsVeDIlOIGmMSlsvUJ7UC79cPY+ppycPmtwD
8iBxFWQmgNPuugsn2alXTbqtWhzgX4tXwvJypvOhOyrmcHhmMSjNoEdqIz4YJtt7FVzn6JJ+6feG
wzir1qcVU3b84e1dNatqTBO5OmUssaPDIehQWJ32LrVyjLMZfclc9c1kCUnuheTPdErCLnl5NMVd
sBTV6Z5zL//qOzVJffIDYK7jdJ9vINzYoVCoVnPBEdQ6LxH5rHq5xZv96REn46tX8QvOR5IqbOFd
jp66n1nD95Ua7KbfakP3W/Qwmo4BI+pi5+0wFu1Ygi0yu9WVcGDLNBh2BHpzNTnzqn2SdNr9cC9D
f8nf8s9WRT3a8llcN3wFTDI9vBGj1RZrHvJpvRrlQUsfhfq96gEJ4MJiabBFm7hD/txkCFwT/t4X
mKRuYcLzdyWIW7GliKo+Wz5HxzWAlGAl+QfYuK9WouYCSsVbVr8T5lsaeGR87NRLG88M+d19xkQH
Iby6Q32DffiOoIIfDUnDjkh/4Xv5nL7ZY83ooSTxeLua33+ri+EP9LC2ePGMIBlNy8RTsscYKDHs
gvQ7IYI2iN9KnFzG3TY5gj7etWAGaqT/Mp4IDrxpWowcDVHBJ6+ZKuUhTK0H57ZZKmEiOo4YIdkd
1hY9iMYHt8rHscVAjFiBOiaC4YnBslta/vxkbGPTRWZwSFaJG+jPIh68I1oYc+sM/C/Bf2DIaOuM
mo6pDbO5RWbXuW9Bd1lMvX5I/xlW2gklBFxe23JH3sfdLajsi9jNkRkssJoYvf6VZVdwfjZ0cc7c
AY8hoRgVOCPQYziLclsOxVYsiTVmR2xWVmgpj98cLIjhXHSxMOA0bxxDApxWi0uEUNwHUlOEk7iy
AH0YNa+JH5gKNzCSyEKBbh6seNQbnDzJtkIpGbTvDFWGUkFe6A+jFwiuO9s0r+ajJX9sGu7A/ev+
aqE/1+voae0Ot2E2fO7jnX830J+OtiH/p/9Okj4+OjSDU5yBK358AaZTsFFH72O6snoK0lebBlTi
LiaVuT45btkbYk/VjxboXfSK+Jlhf/Rjnfd2wPj86qzm9KyZnBlCKPlvHScSRiF5vCT8FIULc9Aw
CENPnv4UWA0HI77PM2Zm5cxv2pbWFuYGJn6gTLEHmd14KL2XeKYjr8ZGAmk9EZTe42WG8daOMw/t
46K0VGiVyFdvmMkXWMOvlYPYA07aUPLcSa+AS3RMbQoZ3oyCL0GOVm2gn7u2CXgoIxFnqKkJz60r
kwvoKKspklWj5VmkZJ0AkqxJAy+/C5jlEXOH0XdlfmRE5B7xlSWplS0I9v7k1S36QfGtzxN49Oal
pIZEJgioClDNYY3RCmGZunp3wbVgVqnrUdDeeAQzGEDuBt9lV6VmrGi9ANnjqnezmIEodQgPpFGU
wskYSglLoszlo/3jdVMTj7PPf4h0z/EavfkVBfaGqajCofAGFABBT+DNbOlafCz+/jQL/tRvqDkF
cp6GATsjq6Yf5go3wx5HDXAwpz9UQo+fcaRITRmxnl82kTW8Z25/2YfTI5hn1FhnXBUw68v96RpG
yvJ1C3mbm9LJGM4FSXNd7edD6JOcXRAORbgRn0Q4smhs4l0w7e2yOPTrvK4kJJS4DAlqmfiT3OZW
UbVM40K1cWZo0zTznbMXg5gViVu9ceVKy5fe51IWCYTdnGyA3xLBjjS7IfKxyobucCVfts60sWBM
rsMASxkhcHOwzS7hiJKb7c9/QMtTX4+ML//RiHDOh6MUxYBEruayG9ARXh8at0Nao29ASHCkhwUT
1ptR7ng438PF0KQY+SbV/bWXvqWEWFZKwtsSD7lXtHhQLTo6He48boXHY6ujMr5PZPTJM8jLb0Pi
nQX+r4MdCMXWP2MOKDYwE/Y+0NIZyRFQL7TywLCLU8xmOC6l6OCt4sGweXnOMu+DI4b2sxPtwciT
8EecxY2Jkyk1+gRaKIIEKMO6Aw7hJKXb00zZqjackxOh77OnsF99FWf46TAZpk+MRXQPLcVNDZXi
pqN2OFduAu4WgM52Tt/ASxXTNteViQXEt/U6HPFvFMnwcNCoPrdH0kivSXo3HjlTqgtST79pzzj9
3eZ8obXZTJW00nDF4E5HGJes+nhifcwrivXzjiwmaRdGiBbUR0yqzUIYNe+6Ox91wdGCn2Mx2aQE
/Kae9ObysqcJnvT2pbCnsxAEEjVUTRGUJz8CvdYxCZT+Yi5FJpvdFK54beDuG6E15UFMvK3ZBIqb
VQfRQ97Cg99OzDkp61w+niOLoKhp3xa695hsEcs9CaVdVwGNTwz86HBrfGvEEztwnRQwag0gJLYT
hNECDb9LIUCgBKgvg3efskW0/tr15pH8TkQvR7QsX1aqnA6O/mQKGPo5E9KOD8FCv37Z9vw2Pbnc
FlA6DuMvAn2mDKyAuZ7c6ikBLbWysIZMyVdnLZh0JNyU9hVmjqBVvEIQIfcQcpysNIGenWwa74G3
uSZFyc8Iihmgx7PQvq4X0gXInOcAcoGBXz2RHOq/MqnbTLLjjvteUvDDVGHIhcNn57LqPiN4g72y
/jxzQXucCkvEYmsO2+8FEJs5AsEnLfdUkXda4uIQb3sfNVUwnwX38lCmKVugCG9Pqj3t2dhp+zfN
TjbfTdV66IZe52geZH9TJ9ZZXyfRnXyJFAmi1QFKfdCEFLKTSTk7z39tq2BozCwvKllT0wCJBYsj
/oLopG69mx85S5kRI1KpibcfdIjviDIIzGIfsuW5HKj0vinyVlUGAe++qaHdD+4s0xmsIS1YDuF6
0/3lxayAZ37DBRcvw0+5V8GN4iDTLG5XIYqDmYtBQVwrwCKJVrlNh1BYoC79JmbHW8ZiiQe9ShAr
THj/wGktY/E6jhJMR7cAXsX9/FB/5eO0v1ES1miHQUNlBtvLI4jQ5HE8dfceHNgi1PH5Ix4FsFD6
mSu5FtMg1cIY3uPYti3AdS1ZLWEtuYKKlzgql1kLSNOAP9vJr10BhfGxWbB+bqha98FDSC74Qjvl
g1+F2KW00OT6ZkF3wDbPBLNc0Q1UxjzOInHaMTyuegzmCvMyub1xLKVsf0ql5DvjMmqZ6OJLQoh1
O5sRtUUQPH9Pqtzadt/0Kg67tOWBbHK7bsf5yQK6qPnBccel4s2iVlFkTe/vtQF70FIy1s4SzmFa
uqdRFlNT/+oOI50wNjLqunsJvuHQqZ1y4ECyhp5PJ2c1LufpETgNUzNNAYlBimz2BDoS98805R4I
0oyQOncG3yRoG23peVJE7mbkz23iB/joZvZ//KzRIsMZgR6FKZSH3s9RPD+aMmwSoYZ7MZFFuqY8
/FOdyikLtQ8INpzKGRIB2ylNZVzbuF5+AThQy3wufrJuzwc9l7hilWS1H9BIwtpvRZzKJqrZ9emL
BQX95w9JMHsy2/hFSzmgQ+azCut0xE71r1LGPrY7RVG14lZzRSOXcZPIxbiIeguKQ747x+yDuyC3
cvkKwyWkuTe+aajAwnd8XjgMgdooJzWpxRhyUtVdu9fpAICF6ihAq6Dv5VEq2L/A09LfgVjNjqgO
/ooZtyr5rdMvCyG7xr+u0mAi9HB508bMtCDapSaAz1RiYeJaYBgjmOZvKYgYFh2sikowFkcg+Ap4
bDP86OCbMZEzmFThokrZQd9bX0MC7CiNFrrIUMeuTOMDg980HD7gEOBZT0kuTUsmTCkKJH/rqVyq
fWICp9MrLHBkUAVycm2qP6mtbcXdudw99u/d9Ips45GV70/GgYIwL1wt5Z67Xy8FMKqhpXgLjPsm
ev4/iprp4rwHJL4PY0gfxOpMt3VdaVRFfHduHuLbzkEfr+l4eTOYKqM++IRL2RtUF6lMym/HDcbN
owpLyH43lQO59Oj3AFt6U2D+YNME6UCrK2I8Q82kji6PVqBQMjkYRctw4+7KZaModlXi6nKKX8kD
vonetsOCIZQtUEbA6Lsxu+IzBq8JJcXkJxaUo0BN2cCROsz14EaRyRAhP3Sl/WX08uo8H4a3W7KX
U6bMVG5lYmQJDTKgiKXgtyw84SqJ5miRQAM++veCzsnXpo2SXQyp+ENoUo6Ym6jROtkLigE3EwOh
HdHji3fw/e95upW+cM9zwblhsu4zQCyRIeIapBHOWRwh1AfHpGxJLLUsHL0XG9fVm50314TSXw0Z
5jiMIwWxDnvBP3+FvVEn1I02bsGP681ymvKocta6jV0ooqraAWTD79v4NTe7H0Zv3xBocH0WxW8Y
5x5btOgf/g18WqCwwjlPYOCvQ5yDqeLPxJLgRb12Oki8DgzHPYoJd+mFGBCw+f+E+aptOnXwK6hw
zzWstOmxyEFn7+0wHKwRLzW2TJyyWHwc47MtDCcuh8txt2eABexfnbCCYvOh37aVh1Ep8wJooiLp
tphho211PR4XoGzFb3kAfMckkyQuwNJAF687Ux3usbHDgZVcGrw3LVa+I/2R3Jld131+suzvre9A
0y0N6slnSA9Kp5rTpR///Y3Kaptb1A/ia5Z2aB2O3A5XVYaWBOWWEbAajMUscdnlfmfrcgN301fM
dSsY3vUl/x+Plyn9flwarEPkRRmBm6LRIVDATyfZFQls6lp9yx7WxGoex6r1ikverfvnnb/zTk/7
E6WGUqVOT5owRZ/J8tPBfE8IfAK5KDFyKc4LiSaKVu7TmKtGJaCtnUBtzl9xOfWDskZZBQuG7jm3
XJr/NyoO1ysFFbXEzCRlWdphfnzkpYy9Ii8s1q5LgjaSfkNirwYDJT4YleLdNhpcTWSwKsVrriJU
DaCD7/+Mu+AZsktStgXcK+l1+qcKZgNUG+gc/C49jPvf+VaBy+USMhqZi/oSrdc2Nwpp/j79U4xP
mcww6TZkT6Gg3N7eOOb5OCXfoGd2tsX96M2Y2D+Ts8sruIDRlyR7/ZYmB1Kox+n8ZuvjgpS3zf7J
3+A4ML3mUnVIYyl9QKRVWyCMGUyXzt8YNGV3ncOycAoWVHRuIMxg/aGNySiHtqWbFhNJJr5uPFQi
qvJEjBZALDEVufJouP+6mlZ5gUiU7kejYb7uXInNcY5vocGWe48ywiND5RkRKk0ix/vz1dyg7COA
9ktHeXEN0tJw4LB6eB5XSeceLTr1LqSYWHmIH9QMhI+bxuwvgOBhwM91lJJRj7X/E6TtFYERWjt1
YVNi1/VVDxb2E08KDyFECwQZHgPAOYqftbGG2HNMXZC7UokaySMJQMY5cjd842w/O+rCpcpMil8E
qoIQe8aL/2ZXYlTNWKFFy3EN8fYBELkD6RumtgoqlrXSrvQU7//nFwXfUaKgvz+tpTQnEUjFuMb1
ylpPGyP23zPd8wvsid1I6/CFAiHIb2Cq2E9SBHRntCYEIshPLWiZ4gsQs4YIJj4Jv4+NbCgAZFjd
NaCiA2CU4V2tQPHstAX01OHmjqeGxyG4ZG7HHl2pynmHQ8YKqTyh4PwdHdRU6+qGqyxhbFl8bbru
ypZLFKHFyHKqBC2crBtH3ZPkS8vSAckRZ3yHDoFPBggsWLIxtT1Dn8MYGciohwx4U4x/Ibi5JFPl
cTjMGKCHYAaS1sUZzWZ16c6lcAuvR4UgCZ9BBV+IAiNpPQMUP/FNskmeIbV3ZMTTX26C5Z8cJHe9
ltbDZ/1248t7GuPaq81HXe0Q4LGUmFM1XcnmscDY0Yze6Ul8j/vNFHGt/9F1pw38tzvooDx/QmUm
QBY772tlw0g008VMfiYDbH7Adqk1bB+GCC3m7DIrr+SIPbhDMh2Ce+EhxoN5JwLfzkPOilLvgwjm
AdvS9+/kx8Tp8nQvgefMzEyWimPmy1KAS7kcmIASfzOWK/wjWsuScsEl0pzn2VvoZwSy8mHbqb/j
NfuTCijjlXTwYqpCdh82cWYSjjUEJA7ywo4dNJYe6FI7QhaWAZEcO3xQBpxR4NW0/LUNlffZbCyo
XKlu3gix2+G9+GR8tWCz++PLNeFykpKXzioD81HhsV0a+DqiIW28KZcvbT4yO9A7CziHYraCnf1t
uGeCzqYvaP3OKlYZ4GSMLH965ptp+33xne2xzSh0TFv1U9DlS5zlfdlh4UHcMcpEB1vLPLlKPxRH
bN1FAiQOXIlYB164Gw4AIiyD4cykFsT/cDPBgDxrP5FwGAGj66ONMwXfMaAIURuFekQIrinvlUf2
EPkqw3/mfWaQalsII4U5sor+cX80Qk5ejhrL1p4vcBueVf+v+NWgCiEbYyd4AL+fZo/XdFgaXsgq
HipHD2wJ9kSKyFoyUX9VKQkTyM8qoNeY7uMx/YDBLGPaMaVpEzAhHYfTWeBpMCcQ5K2AcAHTgrpb
31fiOduwDfEGWwZ5roqF42bwBHvigt7nGnXoNzUUmauK0x/ifFxSzjhfEA6hGKfCwK91YNVvh6v0
VKWh0n9IIBRDH+4uthXlNO1GhInMBdRsUlMTd2n7OJaTpGp5WBk6FGyGLStNEKG5Z/mafd+xRtdx
RCnG5IQIsBFMCfLGac/+IqVyCECdvaqWK4aHjnG1ZvDchwuKI67ZIvhYZQAzUZxjQZM9ku1pX+7Y
2vwK2FNWcDoddwdOToQLjpofkT23MtWfUAvZ2CvDzMwTont4TXnpaAx+NIpPbJfic8dASvlLHMeA
XIgSfGSo6hf1KrELsoZTWJJhRCsTJ1xQysjDlH0+7+O5c2ej7qAz1U0MQQ9i4Ur+9uhH6Uv444Nd
W/YVE2FqPPsrdJPUCRFLW9PswUsu9Th1AFc7XZdi7lzOky+nl9XfVKySU6Dk3ferQRykziV6qB8M
bnvXLZo/CKZHnDe9A6dJHHUxoMOQDgFYxI4e20xMO3wF2ZupJlR4myU2bFapn9lAgxcP+J+DGeuf
naAgsN6vZcapYJgLv8vM+eH6N8QK+3cNfJGOpxdlxTn2GZkD+b/uJ9SoGlOdrQ3+5vnWI685F/pd
Qi1IWwSkqP85EcmibRCwR3HLJ21UNkEM3FLd7Xqll2nAxNX5oW5ekio3IiKPgq3g6q2751+v3nhW
cuhHdw/oqg8Cb/jhwV7aTsFy1yr2B5mKW3Gw6DiipIznjkbpW0srih6gTcY3sVswZ2CRxVSuVOaX
UK0wUnIveQKzOxgYQrUUr8uQJ7xwVG9D0YC0hjS65c5pnLhHTavSHNGxmOdQuKqX2r2xJyiJKDDx
RrH0d+zfu4Ec0XpSseI58yPQfbAql6Aiqn4RwY/PX5eTQ3uk8pmY+cqq9ROx8k/rfbS73ZsdZEf6
QfMXHovCjIDa2uSKmZjhv0bHqkJ1YD+MSKDMrUqgrz5u+SAz3/1nQptC6TVDZViA7cIw8sAlQ7IC
SKNg10/HtcdJ4RggnyIq+qRqoFDf+EXgnEmDUHFNOPc3g8wNe0cDNpgVUF32Z6fRZwO4OiQp24HN
J+YXaYQeLsKoj2O5F2OgtsAxJd5v1sU8s4zlOlkABDyI+KmaVu2BJprKEczZxpG0zyOhTtHJYHeN
G5wfcxnPUFq4BKUbCtnW6OnJlJY1D4Drxb5Mz2EPmlsapBsOpear5vv+XYKmebKiJLSbxIsleKAQ
zpJFle0pBKXXhE/JhjA3oi4yfh2+Hkm+QJJkt1DjPpflsTTg8zl1c2q8Jwx4ww5Gw2rG6U8mgOWX
ZDlrib7An9/dZy+lj+K+59H8LOn1Ej4oo+70mwH0ypyvSqpKNdbx8MRdLS3m/Q2HAH5+PwEXfs8c
+ybTZKYZsgTTffyl55wLHTGqu+Dp19reb07Q9NMz4ANezET1d4qs6dJ7XPImshIt84yvpIYL7Bzi
bcLEsGUyG2mrLEPk6ScSW+F0uB2BDVkbAVcgg9SIdp+1MxmQwpxEZ7RNSglpc4Ibdj3E7bIbHCGC
eZFesjayDqKQwZliqaqZ2UDNQg97l0KKDCVKf17aRnQ/lZ+9l+dJd2XCj8Lr9BgoS+4MEcH6fcYY
v0JwS7N11K6EHejuAu0OXYpQBB63M7s1/8t2+OIj5/K6rGbNPn3QERIZhT3s5mzGmXoGp3xEuQ/s
cfPPR6+y58AU4uFXAC1WGAAoPdqPxcBfN+bLnGk+ATKjpVE7j0YqYCwLgF9R6gaLifzz5bjK6Nds
ewZsTmRWNhPUvy7BzBOb+WZ7I6JnBYh3CfNMiKciyDW4fJB69ys1QEY8igUbiK4W6OsfCVMrLakL
o9s1K//CFk+SyM1MX2eTER9vxcPEUnkqyouaIvCJvYeViIC1qJ2iakca3cYd3X8A/I7koyYsiGsb
pc/+/H214hHEQ26oltWMbemqUnCeT9fK4CJUQwIMLV3r4Iy/zvO7qBa3V6gOqDL+DaG9de9s/S8E
WjNVbO+TgqI25PgrLmM0O9jCgeJJAfIYudUhwO0oE9Eac92N8MolMBJKy5BwC7PcmYffauONXh1n
ZtQYUPt05gdL0OpyBZkxUFjJmaBWcs/yBWTk2QpbQAtcK/Ovnt2tMYRvZgDwAu+gAEMDy5mU3tQs
+1scne+TPfQ1asCsAFu2BT1ntm48eP8GMdhzhSWIZBBLNniyu2H65EShLEK8ib/3lEzU2pvUqlKp
J3l7bNjNvU/XPIzBiaaV/wjQ6aVH++g0jghWTX9Uw6dEwJW/j2/6SaevzIUfYGHqp+wye+I47KUa
HUE4uQ1tDiuN5obesVEf66cwn4SNJGOhJwFZuj6ZcPMYZqj/gjzU11ZbesqJ4iqClgAhuzFCk1Sy
RB6MiIOhjH9GwbVgYZfw/vyIDym2X6e1MSwP9p5p/VDtPmYC9poVJuZz9cwy2RwEw+c7HFM9iKUO
3H8/9LFpT4daZ+yWSF0GBN3WeXjE161oIM1cjak+kNoeYv0n8OIJSUabyRdxTgDAdvOPx8nNuqEU
tjlcoUKJ38tR2EgVd/W8SKvOOtCI+cniNtbGmIPYo8BsEEXFXWRoPVCVJOkFPhJ1CSc2Lkv1iCLg
D36Q6BpQBY3UI58XDfKiRdi+HFCLsRE0hlvRpYqTmbjHXr1Q/kIPz/hwj+pG16prrmkhW5GU9T7u
h+ViOYCjpZEQ/dedwqVw5LdmF6ZzQ+VvC92CrgAh3KLHru067jDOtifa1k85GKhX1UZeQ82sy8UY
qZRfgvbpEbZi7pCu5HwtJLaBf3cWzfDybiJR7/W5hEv2fmBQxyYnYu+gc12mRs8I1Kl1Vc7cLFlI
DU5iJNd9KJoZcADLXaAS2PnX8tnoiVBlpIoxnbMyHUtLvVvVSuNA7vyGq+nmFoXMq917lpQWhq2v
p8JT4R398JTZj/3yZ8UDRcQpsDKHYAMpAzFXlCkc4UFY5LjNCTubL3mfV1gMIHVV+wKlViiltn2M
r3x5dELXergM9VPoco/NpuNBZdJWlbBMujwjZmpxeeQ6GoEMW9/XJLOjDgOQ6nv4ulecrM+Z8WuF
o+GbpayuZrDesjYFIuXRX1im9ShQ0Xh+wbUSiaW6GDz7UGIWopGqxCk2XNoGZEtiYZY+WsPfOEb2
sNBztZrmQ8jUrqqKvlx8wmKMm/8N8LmwNHl4O1FTdhH6nbmBMjSxrrBa1/1MpwNRI7o+7qaY/Nvv
E5OsKTV2+Bbe/3NQcrALAHfWGViUe9O77nd9DJn5AyKgD/Bx8hPExtUGSX28+EWYYskYy/nHJjy2
qJdJzP7sAZRlzAaUT7D5dTVYiv1AUqeTZ1gAVjYzs7ubZuMxzcg4XX10+9QMZPn9g4OEP+Jo75N+
DmatrXh323q8rLS0ekBzTZLjjYV1oy7WHSDw9tI1TxyqlBVun3/E91dRifABL8GtVy9aD9g9Oj64
EBJnOBnXk/wNa3eA/a/xemjhVWGg93zkDiu+THFIptLyHvRra9dJAqpU6MoVsCfCaIaWpRtD0ovC
uaCvFdPJB9WZLLdDPSCqk3xEW1nNGoGTgZzGJBW9zzvYSMi1+cRAgFtbk165mzHKxoTLwrisy/B2
aC2lB8VqYnIxuGzUYfO+s7rbGVwoga/jHf3IFK5iE4CUlGM7r0wp8e8/V9/UAGfZgX4MyL2d4i22
MNTalU1srRjfzAKRNiJv5Ft4XXmgZyCOaNe2+4XXu5+5BkkCjRksviDVkKxcL95aSOxEJqhQg05a
MOgy0BKubgCITdF7Lvco/v0cce8nbcswRLZjNKGIkTSbsLq2Z70qcV7VGpKVM37TyesjMdMr39OZ
Nu6BpQjqplHlsIyPVYG49eA/Z89Z820r0qtKl5+2Vathv01BjAoueGpKpw62Db1E2uFo+8jeiQDW
EwM/gHmXaSGBhXvZ0fEDVcT4uJLhy1et0omSGUokozpvcKuz04z6VWR6IsqWLnlKTU3PPxgerPYI
KvqcbSyR0Gdbq7K4MuyiqHAuY/2FKh9rnW6Z5V5Q3RSkGhxJdT79KIqsitwUObcJ9HPzvvzQn/es
Zj1RR4eUATiB72kY7WdMmyi7mLGgkZPSzelQmcYXuDK97/OQ+Oc2JgHcms2avn1QnN9MWmsStNTQ
UuA8ekAEu6j5B1DP6ZonHywJl6uPMIRyNviXqnI5bGhk0JrV+Eh9Y2Tig/WwFnwcElc6+EUWAGMP
Eixa0h6jl84in7q2GT1/WM3yGcSXMLHbjg3kkzQvEiW0vv+lHDRE6bV5XDXbGwQOMMoRZU9/O+bt
zRqOdPcFFQyW/ACk4a2MJhb94+Ob3xwoOBCZMlNEO+Js4UvBbI+SEBGpK4bvE7HpBLr04ZxzAdzQ
c4ltVd4lIk9zOnyIwUXTcRNwLfSqpS7rlw8Eggvql/Ua9N6rd5faYxholjM75VO5gyuWjdZp3pnM
zas4vLw1zp37j41mu4ibdJFvP2ny7Y4p4MnI1IiNCFKMGnw38TbfRq8lkRzXkuhQt8sCDhAC+lW5
HV13D/Q0S+FPCCev/wcM5b3rEhv131Vq8Hko4LUg7mM2WFVNoztCIrkYP6I91cy+uKBfI12moVWt
7cyciBNss2W1SXPd1d4oUf6R2HL0F86/jnfWItAYyjeGAKqXWCkcv2dBhAvRKRdVjFgNkq86nLC4
Y/79MVNZ34JeTPG9eQ1pgxX1NG2ZWxiB8GXIAwJ230av4qU3uQ/L/elS2hC4XeQWSApewyxMAZdD
TNMg3hsSrPRECi0oDEMgVjG8IGvYjC3J6fHPob5dVPswVisZkQ+WC5w5+0NpJgyEqnrAXJipuVkl
wS7dLZSS42dxDzSLU5KIrk3bJxLunbm6PTIKkJADYrxo1viJAIL3WQxCw8/WNVbc+DengYAaUKFM
gbs6NuUEPHUbWWyF/G2Cf+XDqkUaW/dmQZRSaal/XYnZ2ML49OIQDCc9Q8euzPmugCC8TVyiahlA
dVnGB+oZkxBhjfBQoJv9rpv5fphvGOMv0jfT6SkIR/TdUveEHXJGzbnHXuSsjugXItcxZ2TDMIXj
xdcNK7Sgc/iU1FknOK2q3pgRz0hCUxqo3UuM0ftE2gKZ8mS0gI0biz28wpDr9a0ULcqmc3fHBptv
kAxrhM2/CYTSNEmhas6SV+3R9kT0H5ztU+83GbGED037QyBu3pIG+9Lb8XZaNfpNXLKzSGaL1t80
PYE4+c+GWYZyVQSUBRQylk73MVJZB3L2Ah1QCaQh6N8DJOzL3HeAeYRiH9yZho1Zgyz3Yu8iZGH0
OLqgD0ubgSZes5taynQ5jF4tLnnRgxn9mOQ28M67MhBKOZ5y18ttygNczdZdH1qk/V3TYhkZy54Z
T/Lac37mJxE5EpYtlIICVHkYBzNYZr5zRLaPeMbAPW9mDgbiHAUJWnQ7kpNBPBuNHiW9P3wRiawC
d4LKTqNVV1LOOkRz0B0CcOYAnG6Wtm4DarG+6GwBhotidvTJ36MNDqnT1YeW4EDsGzucXmsvPhuQ
febIWlWO0E5DSBwWaubTdsQ1/q7+iPNE0sXuu5wGKM+jMz6Qf/WsLHvUwMOAa3NA9N1twPiMcvMb
N/wenE/IJcB5mxbKE8Bf7hpHv2R3DgA7V9AlPnr6FNWO/E7kRoryQyBzFNBlh56CvyQoSsWamCt5
U1mJxt8h+LpdNYNT1jxT3clIsMDp1S5fXpwWruTAT380OiVRPWKFk3h+rWeL16yhKgH9Fu7LRYSI
Qj4RFSB4UfxoVQgyVjyUKHzLMJ6qbRJYNNJl9t2n/zWWKmbWitkYYnyOxo1RIezOUpNjshEgS0T5
u2yf+fm+TmjW0uVBnO5aKmbqwwe2XgUb0mpJvTSgHzCmvG1hmteoEoKSU6xW0qCz9Sse4lZGNwjW
yd6cUR3c0SzhFdqLvKjIaMKGWr5UIAoQc1zOuXoNFDRJ4O7Nav8pJCZKlmKZcPRisHQrMk5wEaCB
DhDbomAI8qy34jgxz06bD3dFkyJGUICbtbtgM4HPPFbKLjUSKNZy9HnENDSCzG6Aqe3CYZ+YRiKI
GARYtIWNehDNb7Xistua+ak7jbBo+i0h+a2gClj2ZfgsXHkhiohh3kYb7lYYv5UHNXM3Q0Gp1Icv
uLBErGn8iX+IJEduuexqe9lnMRBl1Y2ANdl4dnqsDKsB8H7qp2PL21eJ/F4OSW3r0axCBy9MT8id
+1kvHlxU8qJ1yzl9hLU1EY27hEM10GMJ/8e6rO7s2SfuCXsQ8d4ua9+mWOYoSBFri/XtweHQQoNy
RcZs6Tj3p/lVM2+QAKEWjDXV6z0igDatNU7EHnbIaBElK2NBtU8P5rfKvR08wLI5CSN01YaJxXvD
Jqsvxmhoq2LuLfhu6F2qorD1+Jil0bsbrx7cFD3fUYxWzOEQTr6DKNqlA81TNxeu7Q0BzIEI6rjP
nhfTeqNc3Yy4y6mvVfcEHpMFZkswlks2RS6p6X/74Pm6ua3e4vkzU7tVgEsrjLbuzfMmai50lnWU
y0Wa9eugJccEwEpkFEXpw9nLyU/W28atkasG0KQHzQqu0O9lZfMpI3pfbujLCGzcv/qakn5zVha+
xRzeLaEuKPBSHGB6Bn1YT/WS+K4FhScAMOYirgwNshMqfYc+w4rn5OCDC96WINQ7XSo6ZThK8dyO
MJPp1QGLBLa9QMD6Byfksh7K7eZqtaiJM5tShftmQXpuT8JH+MBzAdqqRTQtucEtNQCFKF27d5XA
QDS3tZn9u67mdxnXGgxP5dEXSJw/Le72vsJ0/1n/+CicSCrWlnzs5QlJUtC7J+F+tSf8BUSiVNtA
sX6jtxjyXMbmWas8SCV2d2JG8pTB7bI4JYM6966IgxviqVhfxAh5grQ8eVeSsOnm3tCWZS9BRFOU
tEKe2TNPRQ9E6uZTRW33IqI3suTOr9zzBdBup56sJumAc7a9JqhLEI4cCj9dFSWy5ydibS88IctX
AwXF5aHiCasPI2sUmmVyH2NbWKvmgiUUbR7XtpfTeOEcjzMdD68azVJbkDVMJtTQQXiWE4Xakn29
Njk/PWa9iHKVjtlkevE7m8wZCgMvY8Vp2PDDpvfysSvYcnvNzEMJSOG19JtplMJ8VDIGIWTriMyT
0TGESET5DVEssZsYI0JuIh/iFO6+3M+3rmOzb7LNoEGld+4UZpBhe/4W6v5hlFsDNiNdb39uF6qx
s5J4mlZhTC+0SoxeX/FMvs6pi6n6qLRiabzLfcVIKDcJDaJ8QZc6z2UymEXo5ObGEWHzJKXTYQcC
BQj5468rR5EO3vLBRVbcekpW8ZoqNJNYlDl+94oglCqmDMxuXiCV6eSx2ZKhr/qVPHffa/6XMuiz
l0kAkrNDeWaPeAc/Butw9f+6etmwgi9mLSpV0A5DOXHKPHHhCk01oIQ3JopRY27Bfu4qE7aoCxkM
qkTioUmhpIdHy4WkqjkWQtpm5w0H1Akq3vLGbp6Mj1WDZWjDs/h81yBX58AuAxXaBi+J3OpWSCmK
w13ZEaPScoaiRu16wVDw93nxpnQsCekjozLxeRxvFnqeCst93YGeZz4YnnYTyzfcBiOoInKXPegz
911iBU3X0JISz9eU4M8NcofH6CEiYJGV/iyTNtQsI93OT58vSpQv0RSZx7vpoyKNb1rMaeArAoFJ
WR5x5ItBRaKo4BREqEC1PsJEy8FOKX8MdbI5nqjO7CzKboNjzlSRdQat3oCkRFV9IK4ur/UxNrsI
eqjv8b411trNpTtc0SeV3vKiSxWVeQhLP0cu2oBVeOWLssMQpLqZIlmDJOCxx0qeAugkuJWVSq6H
4jGDckUtNk2lQJOZPwxAGh1m1aXI8qVK7iV7e9FXC4Iw6517RFSE3BliY2lReo6tHJdr5rTCSmMA
I+tXfKU9glGzvz+RfCu5SDSO3jpQOFOjg9PTWLlb8GyLGgEN9+Yy0n/csEu15pI4cdYRiePIpO7O
S+1lIHtx87UweQL4VAdcKbYTT06mvFQzpqT1DlHmfDMJndV/kqUWOPAspPA6v99pWHvQJ0/50K4K
Mp60sGQlRztOw/YMDGjfWJU3BM3uCoJSsLSBE8o9B8bpw1oKKmdabvQHoM0c0uas83xv5ahV2Ony
jZisl6LrWGLkpwYnE112ZSrT8gbJOdmMedm3c7yIVM4EUh2fBqsgvYGyPWBk8HyTnZoLF5jnkqBk
KkViE/d8ELP9RAqoSfTK3eK9wb+84IQe3wtVZH1VWXhHAGjMk91Az2+sulveT909iyqF7WUkR8Zj
b8uVxAfIF+l5qngD6RpP5bfPN406ysHyZR6+svdH5CbpNug/z9zTQHT86shIgQIqLn+SyMZNsXQ5
G3FNJ7LaooUp5TzcFRLUPBPZPFK8dGZIM7z5cV2AjmDFEgiuJYSUD1J2lYr+OdAyJjJfNeBHXtLV
hxrEQFsNIigEeHzrvGKJqcKyGlnHIx5L/4AcJuovnb+QPrxrOLFmcxSXhPxd5Ld9M/d0MMSxtDRq
NHi38VxPLkwqJe5fLu2c8Zsxn2k+wINoow7ELbbzJeyJw0xdDW2Lhy6tt5uhR6tRJ1bhOZICGGFz
SMJSTetCwrHUB1bBU7Ka4juLYLZwQmSUTyl7pJjhy42d01+6yMdPQSAN36XycIq0inUX7r2kD4rH
R2fvCDaXUh6Wo5OHjirjZcH02xIKdP22tBpgxlkpDK7TBt6NX6SCAxpPERUBxyjlzSrGfG5nwrgp
GSaqcU9xnkaC7fpLRllqpy9Xt6WWey62tsw4VrCyja5kpvF/cY2uwhwK/+c5KRLJvkemdLddCob9
ZILbBQWRyxtEpGjZL0D6A4QJT5Aw+aCUm4QiO10Jh5717dBiFrxPxiHziGsHb/MMqIknvZdj+9xX
qNB4ZtC5cDwe5dJVI+u68+ezVRIAD1gK3TTk4hjUwv60xrAu/SKvG7o+uLqnJmCwD6glgtGBA98t
REUb5C1sxLKVImQcl2Bz1/wwokqjYXsDKRpYCpuZ+pbMa6x2/u4ESGWsapNEmhNLHX0OMA+rmU3a
2cFNWmDZz1FWPrNC41mVx6Nvs0nFl5OR+XeyfrQX13vU3U1/ALBaRu3TsqH8qeLwALXs12UDTGTJ
RftsBnAZ7JZwCjH8FlrUYpRXXbRtUUxFu5rC0uVwU9Qh76eVLyVXPbcRUR3ivhkJhoJKwTeILKb3
CoaUpOJbacFX4Dm79qzW0Z+541sbFavAaobsDDKBAFzsIiNvLOnHkqooXJCV2WBdxIlO9erGpntd
V4mBRP4ogLEIqScdPkli4kxIuY7JAuFBqU0Red3gh/Ggfkt1pxHBWbSJKdSj7kUzIw4+7vbQ5vra
nUsEvxxP54GQ6V6BZI0pFc4IhXDKY5Vqv/SH50afuEKDRlNa9pmtV+XuFBdLzKI3t0WnzjZDKZsA
5UNkgwZQmaWRWrpUdzT57PI15KdrPdGeKBgsQVEP3keGMA12xOfgpzeNmA83/Hvde7jGJN6fQngS
wZlAo6ouebSll6RJTBSCxbkD99RVeUf/oPIIe0BfNZm57B0R8CfmvmftxC0xyMvg3UbVG9o+qw+c
lo/4Z8nSXvbH2JokxgSL6XIloxoHr7XSkhrlhN21mbGzA+WDo76u3RDa5kMZwb6At3OzExuF3Zv+
Gnev2Z8/lohHfCbJmGCTDCNkJ2M7Fsi92xo4H336NBAyVEeEU+XHCXtE1FSuGYmV4VyhXkNQjFBG
ObsJ8CKVSavKmWKXwTPBDfaBsRE65a5HRg/6SDaVb7h3F12VaAhBfSBrranmm0GShZr8JMUMPvXa
33diMYmpaZPkTNUF3vLRQNTiRO+ZBG/c5azjiAfpc9ODpMpWGGHlPUXZ/PaMWYo6VcaH7VQb60DE
Kf2oKw4K9IuKjHM3DYIFEanP+zqUrc/FBL3xUU2FJoP3XkOra5I3Uw/3e68yJBd1x80hLdknTbwt
vxcoK0Bh6SnrkBOAhxJQOfz0zZL9oTp9zXlbbNkfdM6gxfuFsiVcMPjf1wwEIVoJH+jjWvts7ekt
Ou1sqtOHUGzGSeKZCIdetAMWTT3YRQNV+zRGjB5oF/dzPMDQK5rSTRFEcGNBzLeXgQHWYQ7+ZijH
jUTNj1rLl41j1db3SFYa7WSomlnIPHHmKv3BTFm9BAzJMhy45XAia48RgmdJrmysNFy7v8O/mw6D
HhBDIE4D0XLsAKXT6DPqPcHuJHQbvTC8oeOYCqKSpbrdtlK/0WjfjVv7Xu5XKHI9QgCvZhrpvs9h
FkEKOHPEyouuvzjc38ndUCd8gxUrlzzuhpg3YQMLnqO5mZJXfAfB2giO2JGsV1SYW5GDGC3t59Yn
ENm7xqyX8pdT/ecO0iHCLDr/4iMQDFdsH4phlsiwEaZB6XEVVncA9HKrNre9QCoR06qL3nXtpmDo
WgsXExZL9LUA0UtU7A3+AP00W2+doz66vNx0u2cNjdov/EFB883NHQywviMZKra9k/+hWZP7n94Z
00mpqZ9RmrDNA2aZ6/pdECPFD85vGHgu8exHxeJFDVLDhHyHGy1ySTdcEhCAUIbM5vIaZuR3zGTL
SJC80BVgdEgOnRiik6g4V9yslVbyBvZwtzdwj/vsMitSNxdsWQVO1xIP941yBmQUsUlWCnwDf3cP
T5VWjMQfONmmHpOyFV5DG+25dtpYfnG4RAPSbGe0oSpXwO5H7sNAZcFkYr/TJhkXY7TvapTSHlo6
k/+tMD9OcHduoyMuKgZiAw/2JqT0VzJrBj8jubdAyG3kFZ5zyKQC9PzDaEwmvkItqn0To7RVdvpX
/90Cton3jULujKmZR0pJEQ0+rK0akI6QL5vQrh6SBJM4lhVEthZGFsuWbszizT3gR9yJUDmX03u3
hbQkYl8fN21rDsUqk8LlPHJB3eOABg/giqrtflLOebAiacovzec6MGy0Tb81Pomu5EffwZ/NGGW/
SHw+KUSiESlKPrTlhwxUBCcBu5/UX3XizHEck/cvxiYFPBbkWlZhqN7dDbAlrWwhEdCt2npZmbde
J/BSG4hPc7mkfe0j9r9zD6gOXKUaFnZo1rxx7cN3hFsjzhpJsURfxtuq
`protect end_protected
