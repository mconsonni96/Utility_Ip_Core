`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
fmGdEg8vxvqDDJ/Z2xOXCS+B+0TkKVRa9A4dCXFradhUG+H6kQ7SHu0CjNORwvGspnX7Z8l4Czk5
CaF9DHfAFBOj6q2APdRmW6N9fbFhj41u1i/cA5TQnIKsC36SifkL+l1xXyqrbflIJmi6IhBdk2w5
BpcpqsLh52Fj1elcmV14g8jrtXpDTkrjkUFHHhPMth3+yHdJF6AcsdC0XNNurhZj4ib6m2rx+Rg7
RiYhhVXTBqn76fOHj6kfn8DB1JfFdBuo3AuO24ZidXQ9SIELL8W/5yjpU2fQl5pwfXGMKidrVLzW
bLM+gRykN+XzgXCIP4GfTk08vdhz8O03n7r1+A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="VuqsmaoOyYObZz6mqqNhNYECBopwOlTKGssAW9altL4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 672)
`protect data_block
/c+iVqDyFt83zpmOWMxMSDakhFixGseKYzcKdsivGr5+YpZffhzgVVTD3xqjLjcCGAbUGW2TNWvy
BTuyOR7IFOL4Sb34JN9DxmcKdJMp6JqXmHQGB9mP/rDRAfwB4fKnN1D32laL4u0LtCnU/aP2/IpX
z7/ULXXkDSvz/H/wU8hprh4hr+zUS2C6vhbn9eH7T0SoXAxMcrT9LA+uy6tTbE09x3SUOPxfkYa0
VbK042qvanKo570slHyecMgaE98JzggPoiBdpLbb1I9TY+TLtiJl0wpoGZzcqGuE4Ks325Kj3SOu
rQH558GqkQ3cTWai0wQ5ins3rJX5JEqq/o63tDzIJeP3tWB+OHoB3KkNuO7XvuwcCrdNoEcBs0Tc
QJTv3RxfbTUBYYQUjwTwjVJiE0TwkF82jEs0OkwsD/y23xUTen8zasL2cVKdkshwOwR/d1l1IHp4
kO/qIXxoPjosqPamRK6MV+JAeNy40MyLBHhnDlNvu/KYOM+YaWnRK5H5Xy+Et59x6WqlvVTcxiWm
gvZWZ72gbJBinrxCMdRr9Bw9syx1jHcNgfCAzQupEmq/Nk7RdBJ9YGbLK8QJbmRwae/D+BL04QBx
eGeiDq+LOqIrOuf1jFN7LLEmZSzga6AdXmaWDHjbORB6H6impbtSTyUU5wYEG9q3maBbNMQ2IjPC
/IgOWBHB80Nn7J4HL7UaR/6XPJBFPaMJ8g8F6NAn3W7ebrHP9RHyzG2+WDJkg9kAXfJr0oZD3VBM
GOCeME97CZgXXtHuY0wTi1/bp/hFk9M7h3QhJ/NdsdZ6hWOKlH18ONNEZmBEhox54kmvaFYGGXAo
ZHyRxKT/lZ1TqZ7IPqGf5+6un1Xyn0NDqaL3TT0kvPG5PMWoWM8X4Y0N4B9d
`protect end_protected
