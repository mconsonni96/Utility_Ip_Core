`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
jHUWPvHDrnT7bpyFS/jSFFHQ5EB/Mq1dzlZ10PntdgiW5Nl/hA1EJ3MsLVuZ9TyV9OzwW36vm5LS
24fTGDO/EoO91pv/nwJaHXypbY7tFnkubwVg8KiEdaqcxf5NJON3iCbmoKwXVodVhLjdgicfqKD2
T8n9/U6VTHRmag465ZIwii3VxlBS6jJgD6XRoUJGbMD9E4V3OCpOYbTRLCUj0NdwvrWoTe7DR1Ak
7cuo/60JQX21qqk7wqLiQcA3Kve/+sznU9L5cDqw1kB1o85bIpXYRkZYNfCPxHVdUciBWvMxXeCx
DMf1HdzQkf3vv15vDXT92lRnNvvzX0pkCqireQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="xXHb/JFjt/opI1aK3ULRSc7PgQLhr70MeT6h32IFwog="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1696)
`protect data_block
yo1NKYUR3r6QjssueOf/gzwCdhHB139MFmYSPosIjpGmmANzJmfJkQtSo6XFbjlELcsjoJLLx+Bd
+apTxovE0t5qZwUp/5gqQPN8dcQtUDrjuAmT/HXQa9SQAC1BTDCCvxC/hLyotYwX2wqMSbyjpBhD
9I7HlLk/24NwCciUFbiyjnMXiGCus2I9zuzfzXMhL3beugh7t+cSaZXC+UUL9fANhgFbFYRulD/O
4sfPC1OFmELWHuZXx3S5t1gUo6t7ZY8q4yvhefH5ap5palNwTRdcrb41eMYUQQGOPvvEsOg4qD2g
T+wQBnwQVfFTJ3bUD6PD4NvuLOESty2fjXc+lVdE8FyPyhEZ5zhTqnIeeJPJXEFv+UfuoFA9dZ5/
Oktav2yuE+qgRNJxwPDQ53jXlD/1RrHma4tpDZgG97mxOWbfr4ck39dtTHe6IjvnzlySPieKI4B7
SVDdbdNRXyxYEW6O6HZs9awZoqVw2Qr/tKUOGhn2mJkFNlJJ9LPfd4q0iA7e6AGJibAn18MtDJJe
ytwq3Eun7vBS5TUMtg1mEbzhkTyt5FT6jk0UEMYay4xC/OTmiKcn/1VvrrZfmDVky433n7LEu8Jj
tPCt75Rw94x/DXvBuB3lqxOvWhl4DNKCJ3Rqgu4EAbi0XIAoiPW07fgI5SfDiPw8MQNhmzBNCiYv
M2AwRgjjd83bZqWibt1Xjks2SRLUxipT8OhZIcG04Y8IpvXnu9It8NETKnlO5ZgrcEN6vl854Wh4
z/2eOPcDqrdvzYx9XgORek7C3J7ZASdT+HYWsAILF2MXIbsVM9vl8rqMwQY2NyEhjtFxANkx3DCR
w0Jf8oLZCcH9EfiKiXIZEbKR3Lm3blPOf0Bhk51uA1msL/4+pPG8A+aoiTBj8HkLhplXlyDdDnPJ
IqiEvHcCsNqdd2xlvKtjEJ496essq+Edj5CBpS8FtTfDiDBFATKdyYrLOOnWjrSJ452yFBEC8aa8
1Mx8Ku9s8eA4BPa68T7z2W5IFDX8XMZvXTRdGeqaBllPlONhxXKHmYsabfykxuMs1g6zf2HA4C3S
wO7VSGb2TMPUxoMDTxSWwNFWGXquTfnIuxUfcTTSMNjsGJrA0IAy3M9RfNRTA3j3Of6UGGnW6Ihp
DRKaOKSfxGya2bjcmhMVFkjG0x9kC6geHrSYnJEoDHL7x9Zk36WMzOgQNw9hBfQURVdzeU9U5JQJ
CWDjISpEAzt1rMi+Q3Ep8XVKiCQp5iJeWn7O3MHK73hW9I9VBW5VbAbKxIRCBu+rsYNh1z+ADIWZ
PNmEUA1QKE+Af147NruAVXuwRYG/vu/KPPRQ/jcJG5zNEPj1y/m9OZPmXFceIYLVHyicfQbHe2zt
/R+izSXTEyNL5ax+vfwDzVO3y71lspIsKQbJLUMlL7XTcTFEbtSh8aiQp86vnI3pHaWwqqNysBz3
D6WrCPzUsrhszHiL/qjtWJRd2N3qWMZBgUl+vrmaIX0flg8lEm6dnZ4niFCx08qjFopibmc567je
Xu4a4uDcZuHH+KsZH5ykdNlAHVs5nVL+T8tw9XE6v6oJevkMt6KEp+v36c+G7SCut9aiby0pVoHZ
qraSAD5gR2r5y/CRsWdAXYcz/Eh78OnjL+LXs2kuXM+YW8vEu0ABslO2UeoIgfVW4WGO6+YUs+Ep
CFMngo+7aY22cKojK3OgXFgYr3Y6x1zjSmx2Kf+tH9ln6swzPPoVlIYiFodZy9gZn7A/EOEPf2C8
/rVf9jP5B1XxH8fhcmVJRtuP2bI8HnlMKaw+RDnTC+i/5k3cJuSgs8qpmqeeYT1a2a93OX2IFE1k
xx04k9uVh8f5FsH8YNhpyMVnwxhcsBmHxzyHGntzjRhco2oNvEluJbvAJuOdCE5j9491K0PXM1tD
g4Oj+hfeJomRuUBQN+IZyc/i0K5chpsdSD6QjsrZfXUkTIXTHqsREpDgBH/PAEsqkbOq0MFHJ938
6YpCMZ98TgfkfsLia3qUyD6X71oneI7FBVJp1U/lWg3+hWlW+BXgE1qHsnmOq/BqGVrtqNxmFo0T
md8YNzlFWbX4gVS+9/lg7f9nSHGDivrTX4gKgb4aFD8ajC1jR997ZILtCljEGRn81DwPBZtfhP6T
ZZwc/7prRsOM1pqXcNbkNn0ScEUWGkx2/zJb30sV/1W6nK1qQxcOhHZHgg0Q3AEa5Uhb1chZtyZ5
t4MEfvrtNoCmw0ohjsWV1uszdCVjoRHp83dx9t6Puwu2n6t8LA75p2bhRg==
`protect end_protected
