`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
VwSrQM+4C8OscGc2yeBCObW0+puZo6I7xcMXhWPKTR4ZsN17AkBJUjlAOv4UyelwNF9dvKOm/fgl
oZiB+BlZyakx1rcJrkO5Zp25KSo9thB8rIdE+vh0qGt+aZyGSyBFQRDTmh5BJHnBpQVzUTEB+AGF
S5W5S4m0RyzqtemUUI3FjZtWC6G2KkV5DTEAkII8ocR0sH4OtieVj9NuDmuMXVn7Cmx+Mm1MWFg5
FpYDlViBXtf5kumCQHhjrFGKnNCYwt8QVe8j3wWuN/QZg0gKI9pi2GJFh0MVoCg0f/N4oWW6XdAm
9CSxd5kWYfpDYkYAL3wcCqq+WkuX4z7xhjKeag==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="7ab/dvimtg+BQ3u9NCox1fwS5pZMspfYOeEHBvtdRa8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11296)
`protect data_block
hnBxLh8uOXIEh+bOfNE8nJ5ta/YwJ4e2YBQXxLk2ccYoAXr3Bje2guI2pf/GzZWsA+weRq2fDixO
aJVVnkdpPzdu3DKi3K1A1Ltlk8GmFJiHQNoDx3chxQesIr/4FocsHS8+io27RbaUqllWShpYxljk
sjLJdWcR4BpuMhyxfJvMlbAR6y0mCusyxlxeotMbI7hvvv1ytrbK3HYTfBL85x9oXshInbMVSm0B
gejnelS1qmfGgha8AJysq0dcYg2E3vm37IKPcVaLuEQrkFoSPIj9eC3UgHI4VzsS4HgHtwTx8H2/
Yl6GDstT+Q6t7c7cjZsdz88V7/90McOCeZYEmevUiu8F9PG7z9XG2Frc80hcsCO2FBe44UCJK16Q
455K4kdnPOs3JljtIJhBi2mAxCNrCTu1FD5/eGO9NbHIAjjWyge6ZPRyj5ZPyTuPlIhJ6VclbjmY
/pZPf3rvzrFMNQuNRR3iegggo041z1GLshjUvXWUrnhsw+3d5NhplTQx9WRiHIjzAs/JKgmopuDT
S4hP19b8JQ6IY9XQeTp0XolIcGFwYlcE2uLoPoWPGteGJruc19ZXChgqraVIVyUw+w3MQL4ylR2R
I0F9JnANYGhAJ1qhMB6aGSANtgos0XEuDjpYqFxJN7d+fwhDucS3QlPPzUWk85hC3A7MmO1OUxjZ
iOCtMJE/CDeQtehncRybmoQXJ/1fZXC8gy6N7m0K3xatZVB+Dohp6p6yrvtktGPG7MpRogcvfayf
6FofxQlYTZG03xOf3nnrf3SR0VPXnn+9AaZ0luf0jPjFv18JdRzehj/Rx3AgDVQieonkhuVSmR5S
VWn9r+IAV50y59naFc5Sbq9CjOaBISXFbyhdXoHzIRdnEuSV8xKI91YV/Wj4lsxpv6l0shAs+/By
+Joexe+R27c6dhOkusd2GFZ2Y7qjfTGZumxj++QAFFcLtRYFWyEavcLAjAfjT3wUBUp1VtFnEIq4
EPCA3tZZbOfEwbcEDvifYXMtW/TIP9cKBCRKFB+A5aUScsxyStr4k2u9LL9hwpVofQVOoTGlpYTY
0ITWPmx9BiHcST2YQ3eb2B/Yy+GE1rodOC6tWq1LQAwAVOvNfN/glbrsZMIP7tx246oUp+qZXCeW
dIxBVL3Weu5bsuFmEMKfr52QisFOPXzouSaFRqu5ENxIIWmdFv3qqYRPRKxUewAB7zN+puVDrGzj
Q+CnOhtve2VbkuZtCJ0v4KJFbqFGds+Glzeqc6/zMTpAThwHbrIgbgniiuwg9tPXnLZFvmdr4pd/
umDlJqjX5NPwvUKNjZOKyGNevZm/HxvAlvLnrr7zVyEmdZYD6muuIgYqQsIGuxHdKswFhwSRun3h
376NYiJ20ZM2dEjeLEkU8NCYeFItCblPmm1xlUbX74+I/tu+Pt2C5LKl79H3GUwyWkB171Kr2o/z
zi367dLejdasydC2+UWqsmHuIDUcp933Wbdb/2zhiD1V3TqR8aGynOVlDmUB5VqrTITmNHZ3cdSE
OrB7gR8Z/s9NShbmrM3PUsXcwoAnShsADIT6pvu5CYZYCBPGCqMaz9P/PL7qEIQh8UO5P0bdozsU
XjuKz+zb53cCVJqVsQ/Be2rGyuzAObcbltAUjyuEG9oqVFU9x/V42a1QCjAuD3m29WUoQ+gQ/Zbr
tornKogjkagFKRfdwwqypFvgVFFYhIV6vJ4o73+4dFya9K5k4zr+J8Nk0gRcLfkekSvkl5f92si/
6HSny7U9exMfHjaD6wIpAiRPkqRHncJlsifgNAsuPBooOHmmN9HWdeGpzmM0LdJaV223aMyTqtAb
ndfQuAVmNtGSdSYM66Q55NG5JKJbGeiCNDTw3BjJ3wDUu1ly33pXn6UF/olCXAypJvWFKRp/eglM
zTGMw9r9ulpxp3yUDX+kmFHg3+QLefPvTG5niKm1TdlAjzvK/lKEd/O1w2Bx5hbbrCKq2ZwO9yNL
t+QZwKZPoN1GF6OG7Zd/veyTOMGIEIjdZDG2vxPiTO3E+N0ywOZqsvjWaLPl7GIeAUorAHVGjRiO
tVWkNRpg7WBWTrWJmtmuNPQmQUX9Vjz8RUgtefkvQFNgqQD0EIh9TMvmXDsBGPzGhArHrCev4MW5
facjeZA4ft2WlnsE5KFRRsURUXmw2kAFWV1Amkf6++uGgR6U4zeyd3pZFeGCo2a/gEQsMO+8d3j6
kzu2U8qegJKTYLt8IhDxcOpx/ummya7Zp1CL+Roih/HbU2d0NSTZI2IRrYxP1qWEdrZI/+qYM2ev
aDVx+k51ZHsxzvnyshLEJj2QIWC1tJpo3MpdRC4+WQG24IRxl1Yb0+wBgfXkULUo9OSANOPHjHu/
1uQPvoGT1kSy6D/PXgz9WKfwTkggdLKPAudRnUQVqQoc2giKN4QUJOYhJ68mFoh7rDplWv/qQRv9
36lujIOcwyfGX8S0jQKvfsS6FhGbY5QX2JWJV6bNipvpFw8bIXkgZSl39U/HMEQBt99EPB363BQw
WG+n8Td5eqJXVIjR9DSj+gIPz4UFVNl2gqynXLkjHJz0vwyrHQLBPlA01m8rsifsDjAMmIMNvm4y
BupWIEkMqv4tlNN7EFPnjzNpJ3mqhWV/x64U5pf6mpCC7pq/U+nBVf1K4G2urDKtonWAgWFmCZ30
CC5WMjJcaprKlwDuE/UfIDyeUv9oAaxMRNis5bSNKJnfRxam/G89mAjbXpVFTF5L3wqe10xq+BQ0
Id5RIoshHJTO1NASuUogCr2GkgkBYwQroGm9hq/T8A2XEGgy0XOAk4sy+UhdS/vwi7Ie4jfw8/1u
c33LFGteJCyYT9kMCyHogMwEw1DgSOk3nHuyoSQKoOxYqUjYhKMg3VL9YszRjMs+F/Her4yBTisX
km16jXGVTyZqk3Bii1k89vpd0BrBrDMp+zUajZaqwLLkx1MafKjpxqZmfRMn8p1fYXdRVF7Gofmz
On7/felPx9HcZ/ex2vqzqcv5jMVQDBupQXC8OXgl1KkjWoUdWE8uCLMgkxmiaQQmuKqTRg+7GoGv
/yoHSKfBC/3vrnMu+ZnyGamhA5aCMzq0gd3NI2zzkr3nnxFAIbF95Z3SHCZ2ICu7BzPlfeh+VyLF
gRDBINSXiVDq7BkdYVxAyy99ewmDXXjS0189+m8JIpNrwTzLUwo+Wfq9FsqulYm9/RuWY+23FuKL
QVwPQqc2b1f6M/M4YZOVdPAvRJsqXk2uBWBawf/OyKGNivSi/H8la+lDqdboXctwDcad7nTQONLm
HltK57gTagKMj677cGo66I+CKQGeQpanu/Efv7LihSTCDrY6WMgBR4WxLZPLBIby0YqWsmkXjuyl
IbkzHZb1wtloQz+b8cNkcZvhl+AmILXfMDp2/l4lObHRxRLQ0SsI7X7U0krppDt8StpIR/rP6OqK
noiORzBEuW2vHbcgyiCTFkKmtdWNiZASfh3d7BAcbXtBwva20X96TmBhxQ9Sg0pwZCkGzKerH7Rg
2gy/ueGA36NjZunUjiLeJUDepwLK9emFgKyTr4OO2ySnRatawC1Qkt4Q5VjILBhemxcHxUnQQV6I
kC4N8Suh99tMyQGb4wJlL86I3qFP4RzPVqvQTyAyxgRKX8aVh3oA0aV2OgtnLPK1uRVrTiTYOWmD
9hYN6RlWojImGdjlBGO0P55h+eLdOc89owE/4PVG91oK3zuRzOxGxvVAD1fm/gvYF4acOT4T3HN0
ooLaXbwJe9vBEZehOps6vYzLs6UkadXD2z1LryLOyfuHpVjwEoG9F9LlTIN6QEBH8iTFnIHkrEkm
rM1BzJkHWHeo5TNx7D6xoKmlMbdly3vDJDmaNxfUUt447kjieJI05UiJv8hIddy/SKOpWt3LfvOz
BmoWBydVYcdGMnZE039me4ie+HENlERgiuIpFt2pNajytF1tjSJSc341VfB+0ttR10Fxb8MgoEFd
xRF242C5c8BZu0rCNAk+Lr5jzSEBsgE4y5LaipPOJN2D0emgY4cZhOvt+jJr97Y/iyxdR2IZOWD3
l3rQlwlgVZX7qn7uZeVI54UMQS1Xt8kta1ANNWvFjC33z4KietXgebdDaTK8GViAC0Is1WBTQPFx
4c2U0EXTLSma4vspAoP/VA7/2k5KdADPlLxgwI+1auWtVIOdHZCzA6BCnS4zdAaA0e7Y2Dol7D03
p2uYl4cJyEVZ1r68SaluKmU6ZS8FWWzdOZJyxcU9x7utHRuacJCiXeVou32oUHbSq2Bom2bwOLeA
raKVe5RhVtVCrc4t3zUepE0HROC5YPD9NcRzkAAIDaopeBFF2ZyOBlIwobtt3X1hFk/n0PS1/Wqx
WJmBmYF+RLLwE3dnU4slsJjeufI0wwLlJggL3CSuwQCs0ue4q+hsLSpYzUI+OXUggoBcz5u8TaOh
bfUwELURMvfsLe6IvAdO6cdGGf9Gq4j3FD02OyoiwpVctlaKJnxYJBP6N6QEXBD98OxMXFNgyhoo
U+HB3pJ1eJPgcehPn58lpLfUzZLE+cqcLExOEJy62ulscZ6IMmtqEnarZ3ljA+ZcUAnu+1e81Ryo
qI3yUJnZIzG+YkEUT9vZAkVRjQO4Xigp7TU11WnW8WcZoR1OyyliuYpSP/2LNV1nMqHTVB9s+SlG
jBKSm7Fnvdua+FnzvUU1ofxIScLWqPO0U6YOAGjW2HThVZSDTjHAv7vzp2mDaOT4QUc8za/d1QYk
8Ax0daJtHXncPl4oM9k2G1yC5UXBw4q6WYGQbFL2e7SNWfllDlPZL6eEGY05w0dEKW9PR6TzIw3V
haOasu6+VZ69Sb/Z17ZK2XbXQlP53lEVQDZRSUP/zYAcP6d1L5y5s3tAaKwjKntSC1URu1rsROeP
ohqvP5ztkAHz5Ze4u0HitGaFwqK7LiNfPsxDExhfP0yca0+GS/M4xcwgRDcx24POlyrU3Gl7cMYg
APTgRLMLcHyTstYcdV+MLDg9jWM+GOYILIret3O7xezxV2JrwQcu7apSshFkJWOy2m4JgkOL0XYC
+qYXOcAhOQi8822V8GrZMRMtKO8w2U68RobhjCEg7Y3KyVbB/tpCe9WDFTdFeDE/PBX9wvOYhsIL
6z/2dgvFpT/mHRD6CU8F1bSTH96Fq9SA1fgZaSHYtaf9gTJQ7UV9pF2Vlmwy5YrP7c8MduujbBv0
CID8fHsDrPt4m9k/ehwSm+29k3wwR5PR2CB9PoA62QLGrAETSAkg8txDHGttGMvq+CYfTRgmPKXJ
4205QmcnvFk15QPgvGzXepG2eaHqAXZnvp0ISfAJ2e06nJC2R09MokuPnFIeBsunhDxB7cSunS+V
0Z3f7nAvUClecZcu9xjGX3MFzuKhLvhOHgbHQAVjuRJ/roJ0P4bPTHWI55oYeFTkEtpZiQs9+e18
JkL7z2TXu4JCvpURFyQniecFuzK8uLibXyaEfPgXeXNA7LezYgoNOTBxZ+sXZgy6wgLJjuZe2GKZ
a4TgTYXLeNl3AHvvm3+hreT+cuKUAaye93MtaM9X0mc5toEvv/IZ7gpH9rBLIR9FWs9WNBM7Gpz1
2B6c2yJUj1dA3WvHFDk5wEcLPVdJeGKc6AVr31tlkrmNKyFLruRKNjRVWI8/NGXa/EuA8VjZNXT9
X9WdivJwVvuPPn4Uhv+FRnKcv3Kl+NoAvACpxT3NEFcCAiSSMNKHXW0A+QTlZoigYaKR+QOhHqGu
IJOGPBpj6PwKGwQHDOB34D6133A+a4ajYAh/cyks5+WvzkeWgElx2lbbBtZIWDa4EebNhrDSdrp1
24XyEECSbfyN00BHphtElv9Gm4dV+G1QVQui6t9MrntYoBO2CCPSqUSVK77l/krFFLobYFfE6dKZ
vQX0TssCELrrK8ufvll9ZOTzPqJKpIfUwyUVP6M4n/xkP+gjt2DrKRJFzilR+OnuPV+cHMndOvOM
Vhnc68HBEqV4/WDCb78Jrw1Fzh3Gk1Prinwf+Jl99NpTkfubJR1T2qlJSRVIJyV3dpaUlxisE+ix
zDixLiJxzYXS/KmC446OaAI0VamNGeZDXDfbwF5bxFCSVd95A9e7pGUvt0C4U21/c7e6UBxZF1I2
klQVxojd2+1k7DGaEoUtczOgCXmT0ze2NNmq30Q5n0axTAS+p3Z5PFX2BDPcDA71sqzRPZID/ixC
8SfgLugGzlxEQgaoNnywSxwg4ow7SKFssC42MDVcPPA7vCg1zEv8pJobY7TQU0BAyH0f7K/7OO1d
/FwOIkZYtEl4ZhCMFXcwya53IV6f7p29EYGALS/I6cjuRa0OR8kAwpBq5ByMFIqidUkPhJeJREpQ
8Ao/KFxkUZVEhLSPg+QgmnoRYQlZvPfTCLodwBLYP2N0MHtpXL+gt5rbwpB7Ca8wCaheJpzGigns
wW7OmoH9v5HDMdUFkRPEND4mn9qj8eZYe495EWziHQeOcoV7U0v5qUuXi94zyLukgfFAbHqGgm/U
jxbj3kWgSFmyAUCW9GlTV5xdvRQolYHym9eXMYYmYjTWcjBQFrS5rxnGBJ+g8qBLa59Ej0dlsh16
LDNsK0Ea9M7g1HWUJy8qwbd0Z7j/yAmtGd33EbXzy743DbwOHb9panJpNpqvIRV5TbkxNPrdo9a6
gKt0sKq2ZuOn0jm5nP1qGs+EAf6Pt3F9rwICzfFrS+QENbx8jGVRgAHVZO4SReio6g80EUxduC+C
zJt4wRPOAt8BwKeDgOsb6tdpJoB3mBAGo5qlVzPosUbMkeFrFpQE07hjEJTghE79N75bz0v9kA6M
hlDrR/VCWutuckNoaXnWuIBi1EZNW5xqLnAXteH4b2MdyBuuT54at72PjYIDLD9oMR7a6ur5H2K8
pwN5Te0y+0OFgOQoB40EkNTfdDD5fdpkizLGZBEnrOPhWY3I/HMUN/+O+EgK0/hjPJFl1W6Cuz0H
JlV3RlGb3d7JRX6z24twgKywl0rLBOmC7Y/s60OAvOtanlwuPyzlI8agezndUjF7mfudDUZMOgr7
PVWVyY9+hYUEKUIm14izrc3k4123lwF6H9fnPs2nNgOug7oNzEuFELuKxMADtiltMXAZTqVszIVT
NYApdsTirKXdBzguNNb3n4h77NM356gXQyMorCKQXiuoJ8wtd2jXKCj0aoYuTie2Xi+bIfAyZGdU
adctlvr7ughW32rzkJYqhyIn+pD2zcBbIk6/bPuUcAIgxcK0gtamog/TUSsU27IXhEaKsjSIdbwC
pCc7QcLrLjVri8ivaFWU9kOhPqSaoRroVaZ2iE1jlhzbglpEPLgH0FSZKUXZHYbjLoqSaWXN6ioW
Cm5kJ+BdNIUhW+Xsnfa7kbaRJa/dRiNeAqOZaKeZKcUJ/18JhxR67Vf6AJwDpn9flis4du6qBq5D
9ieEPDi/Du13LPF2m1O0MKzcDEX13YHnfW+H0ufzmGLzY9S6cTkypRgiWDESbMw9G+ekRPpIoxJm
s9skQ50qA1adIfHse38tQe9cJLtpFXPENu6X8CAFtx5BWKi+K6FOK+oZZUC68BT9BIYXa1z/J/8h
Nou2SC2haEdYejML5efqPEuPkvaQjd2FiDcoHCtVL5Sb09D0ZAVF8L6pVhW3D7M0pbpFtE/4UpFd
22CU5e7w0MgFDAdEnD+9ERtjWpTgEk1E1uO96RY2DVqNhcMb0BW77Cu8tfAdWmsCzgQa+ef8+MLn
rwxnjIly4HBoqeYB9B2oAPJ2u9GFCM9yLKSAl1Ff9+QMhqt7mQWlKemzLFCKVU/4ElJC3RkTXiYn
DtFSs2pGV2pZI1gtr9TYmeM5CPOZQJWi4eJBTjsg1zVDvRBQAs3/wqUYp91pKNuG83Nz2vidi8Kq
2UC2rh/DEQR+TbdRnznzN+EMba3b0Sq0HJ4/+YBbM1hNd7tVpFPkEv5nGFs++maBC8mJF2czhtsO
FAtSASf4vRpp2C8IQoRjx4mIjRDuhbSTAJxknhqvKs7+8vcH5VP7i5iMvoI/W9fnYT+mrfdZ/qnP
WCJCFT5E4TkBW0NTk9otVogH1sEcd+aWLKNo8X00OIvENn7t8QqYGX1klqg4zaSIM/kQUFzOMA2G
REL0i7+bdNg9U1sObDoWsAnSagAD0Js7jd2QjoylhGQtTATBEw7k6IB3HuhWSsLbyv7rZq1Qfzi/
ro2pQPzv0GQN4G8PkhNjEp56iWQ20Pytl7pxHDkQwWAqZR6DCVcVuqeSa4RMBkA68rzpz9CmUYQl
OqwvdZ6ykvrhEv37TkTPsao6oq2pj/FQGEfyNvar674dyTXZR68uunzdDiCarm5d4cgHh5gGik6+
wVRyyUwpSu4p5jRI9Ojbn/yKyDpCxvMQZ2m8uQXK49x+b5Q2U8DVYHJHxWz/7T22W/DfLoLa4v0Y
jriqwFbWdhiyU9kf1o7QD8eC2CmGItWamZ3f+9Wjo5ICc7fUX4ZGEzMNn+Al0eGleoAO9PDpR2FD
6mJV2UFRJr/MNpQEMxMIvpGxw4fFyc4zzL8g9+y9JWDyq6m9r0oyiBAaMvJXIRdSb6sxqXKeVIhE
hLFEO6qObmaZWpHeejLY2nh88sFmOHtHFdYpCapSIu1TWmXoQJBhANpqoZarufEitDwe9kQqxEUX
EvwR6DBMijuFXhaDS17MVi6kH96cRtw32YvfaUtWCay88CHHn4KpZrK4M9p6BFVRaTLXht/gL/gl
4zAOVA9dWTq7ceZerkV8DKekGZhYEVBzvyvWUf7FFlMWUEXNh6UyVTSLyeI8ysmjX+SQGkGt8dyw
s6kiTBW++emP3Ez+Xk4T830g9ncAMlCVm17Wk4GtkSrLMK7cekrdJpE5Tf1fqAhShUPuf74bTySB
xZOooW06zVSSX5XfqkNDue+HBArbee1GO49eMPKm/MRYgqVLPrPU+H3ZnoxV3UA3r4C2NTGNyvIW
XcmhD1zBx5Sp7tFViyUig9OT5PemTI8h4s7Fz7V1KKBQVhV4soTvXQfqcD/m74+vA70gJvQi+oA8
y9c2Wgw2Ag4/jaNuosMmKhHM6x3bqMSwI/gQjwMZGZf2Ntd/80Lwju3uZ/vIF7xwsScvtFgrXrIU
j7KZf+Ne7OvK66wrtjh139AZyqA/pTytonqDZmOL0bPcAHzDaIk++qJkv3N9f3lKimVV3hrZdpae
cj670A9n8f0eigLv5euSp17XFFbfdc2RM0avRi7OsoMNOZp1oNOVsWuBL9yQJJtmqydMNe4NqaPs
DMcasm/YImx1rbH6rtQKS7JGlZQ2RK5enNqddemQi0tCSGO2/27IqayMLjj3SHsH0MKX+DNdHcOE
bmQlUBaRi86BbygKcI+0SCq+ZPDFCU5e/5wIEvK1vRdyUTsVBznbvD2IXLhxQTxBOuYSwwySJMzZ
EdExMGdP2xSs6xyNUC1Uuj0j+S0KOCn4tKX6Ft9AALKwLUitDBtcOsx7xTot6I16mPfoYA/AHhtQ
AhklLcMpIj6PVpUjR0n0zsNqLzvP+CKw3HtusPaMoU6uwzk9nZIgT30TPspbWphMq03j5J84cq0F
13nr8IA8HtEa/YoFe4VRBXMrcPMQRmvhGd1Zak97D9szWNTiuKNGhqgAD5TsuhnERnXXSgTMPSnl
+bGUZZamh7YMRf3k/2BmiYCsUe3LLeB/kVjh7czu3abxhbf2MQ93C4TWMF4oO93zfR3ZvEqIiUal
+TYcDAtaR65uEZPKPfzHDhyIyiKT77IugYk6xFybf2fBTP/XWnt4vYHSbSNKUyj/usEBHQZ6BlO6
YaVoaUlzpvI1exvduf1BUefHzhHBAZKJoq258eBNPhWfOBNeUhN8jtUFc2HUt1INZ4nGcXD1Op5U
wE7eLBL4QbXG1bpQsPCPy32yGLrBG/h8IS1vOKysQwoVpfLQPKxyQwxiXYzHcdlXGdrsMaLIQuVO
UziJw6NOWsZJrB3W9IoMkkeMH0R0ed7o2+DBs1FAZXpnuvy/s5Zx0qxZHE+nV+NsFpWG/dBauY1w
fGjLO8Pm3B+uP9ILSe2G6KgbdOdmisPbVZxHyHTOjKfHhthAQyVL+KeY4CdVBp4IWBWfs4dK6oQ5
NPA8B+Vt68MuyUu+ZBn/hk7wqXbhdyEYNGjp4+MD7wUT4OxZ8K5GzCeuMd9/FX31fIL404EwcTwn
T/85RbgoK/E8bzFeRAiXrFULiR+XewoVEzoCoIg4Xe1X+Ytl/crdlJHJQt9nSLJAX1jwB60XKmkU
E0zsoOOxTQVdjaYi2DYrjQfXIfCKMrJXx+AOKVLZ22BhGDSx06jiqXAmK1QRjJdwl5ScR8EfXS55
q7w+MzskauiNnfl0nLFexAYnkpWrLruljkN4RIty2cDLye90b73BWwEtXKX6S7niIklm1XRJEytA
raXOSRV9CKMNUnYYPmihJF+tPYgqIOjDY7jdZcvy39gtxBF9iVZwUSvNrCIj/uh/nvlsvgrHf7ME
EAGkzWaI7geuW8TFS6H1qmrkZ7X+wVJh4VVyRrKGyoosv6wQsc5as753I3FRriWl9qXbvoxzLMpa
GO8pFouw0SzPOnfNcNTa2JB9PFCH70kQYNX3rw5GTZ4eSihvBQHo3P4EanOgpquZY8J+uBe1/nAI
V6+hLxoPuBt9kfcFEcDfLAYv9fVXNHcYepljEC7B0Q/HPHb1f3s2G76oBRFrTYDvcNtXq117a+gL
VmMmrzI4xhtf1XVT0bgXba2/XsZrEEZEmQapV3bY6vLlRqmhBjlveZGapdy21jSffjFlsIO8KIUS
DyjKge/jNjChyohyH3sfzcfWklpxllCw7zGU9pSgGqrV4tdNMDE/6oqbFIl+CLz8T8KyVv3in+dy
z705awT6LAT4c6jebnXvb/dh7XpufVCmx4TE6sbllhK3ZnzQG3W/lu8GIL7/rBAfF4nNK2r1vBEs
WlRf8Sp56/b8I2DamEADPmN98jK2+PPCzkW6KtBAWI50ZsenD4MSAR/uLUxWJ5IMdA+wxbwvpIKe
BDVXTdwEpTXhH9FF18U1qmRiZxk5s5cs/+GJf2Doiq/Xs4SVFN1qfUgl1Fqmm0RTlWxdm924Riqh
WIzXf8pvykdTzLojiAjAcvuiVDxhODcA/nTV7U7rp9GUmMHTQIzeij7chAs8U3KwpuYkopqtVGH1
fRWtL6oRRg81z3mmd4e0Ztkw9MaQ+SMSuPAc54eRtj8/MEe9cUlUZws6lEHVe/WF3duQ1UeGniQg
foQwJL0l7BOpdp8OMkpWVpBO//B2uDHUf3OTLt5b/WW6lNvzGM8MPQdwhpl3ijlm7mr6mXr7m6IB
UfTlgQBig1dYJPWcP9TNfGiYtpkmRTYj5DqeYGe2ypXpqXS4IhwsCqf7ncXnDZF4eA0Mj631VD1c
e8+YxhMhIm0gfQCknAg3YNT4eGpx32eBBpKR8sq7u1GWOMSMkLarNhRuV7KC3/LCleSvZIcNNw31
xJiw/bNwfmFGUgIi5CV67FszCgH4HbdLyeVIuwxjVZZkxtwfJNGuSK13F9SE8T9PSXrrCnThxocD
rRjKl9fWan6Wc1U0z+rUiA3N4QKR+mKOBM1OIBtU7s68DvjYPkG6msAIh638+Pe26Ar6UjCoRbg7
pxr9jsDTrYfWeXHPgJMt0VxmxXDEDhxeLsaDIsVtAU81T73JMPoHWkJodYJU9r9WyRVmxp/ZHrgb
hkU/M40EPuiBtBqI6lnlIy41CPx7mD1P2YJwKMhjTUZGDerPgB1RLVyRnqVN2dZKa5dfBowTVUE9
k5oDxOSHN0pGaJOvfLUpCPOsdL0+CMntd9tU34Eb9H3ygObWKx1M+Jl0CJIPJLMPR4bBKH+9fjt4
CF+C4rDjaZOj/4ZnUVSdsNHQQm7Fu0XXHe4fvj1AQRx0sNJS0N51TO0rd+6u4x97uJRARIAXEc6T
nru5QBovZIq5m8zeTCOvm9prusluDvj3sJeYWvsbTPOdt8EOWgPBCTZZBD3fGjJpbV1QrrJ3/4SO
SdKqcEBlIbCgHGVOfvA+1beqjdDNtmyi93A1gxulVeKacqNBCyqXfZtu3I3pP9DF73+vj/wS/ed7
S4t6VAw4rA+XmSRuqXL743hnnP0gmc4sXP5lTLXVjkvi0NB6szxE0w1NBASLPrRxA/R0yN+7Eegf
vkaqjRKy29YySaXyeCjI7ycRbAXls0V5HskB/9FLyWGAaw0MFmikgHUrl7mxMezD4cljYjhUYWIs
6mp97UXQrcQ5/q8kDX5u07RWep6P4T2OWasqRFQWry0YryZ0t1OYzfnqAMlamtQb2VHEXzxGtATs
AVfdsPca4bCSkuaol4PrFQP+oyjaJR8toL0g+J2knDjRp88NGvdNqQmZhpqXqxClwtddShLA0gGL
zbR+0CLX/uwC8Vo3JMETRGwreZAhfgwW3I39U+RpIRW7PUNWYZjMdbTgiKkdSu1QUioQZMZ3f8uc
3VPcIMtHvNS+XA/UsTGHXriqP0MFqhZzTJJ+EKC4axk1OSepkoCPdccwJYPy5TAJz7iUTVIdsZiU
9JHKjaw2yV38D8aQzIfH4rXN8hcWMEiEiA4Pfud+mCdk5t1H+SvtN74feDNqG5n0IhXw4RxmjRd4
DmCS/EOOZp7QYwqCKBJZj8EIFLCBdKQ76F6r7xVfjVNnkhr9kw2yU8kiIljUvnTu9AtjGhzgWciX
TNjUfT8TeqWHAxwBE6fI0oHUt6GW8Y7g8utfs2shgrt9y2Ew93U9jgbX4sn2oNir/xw8/SJai8TF
8PN0DYd5d2++wAKdmVVC1yGyRxSnwfDzjGX+FGUwhCZySGYrElRjGoE3Os5V2SNYZ2Vi7Y7HA3JI
uQBNlE3zVyjsCv7sFu5L6bp6vGw/+U93aDMjsXwlDEq9E4p4upVniexpNZkBRAUREivalZIiGK9z
+QmPPfLBS5i+MuxAnRtUrWAyuBrTXIXNlYWQLzR4v2SphquwAu17boQQ22641e2KNp65/g33Z/KZ
09OmT76F3Rp/icsnlfQXPwfVeW8xDxHdwrrE6lEHc0cJH9tpUpSE7VUuq8P2FfzxXWlElb1JEIkO
CZnFgTT1JFWbItNURs/vmJy5ODSRAeiwJHdMSs8DTUywlqnE18xr1NH51tVKXhdRwR1H6VwrscEO
jpCvucWyG0K2up7RtvSGg+TwFJzbizXfsz1Z6OGGiSTpq63ULqzfeEGJ/KckJa9Ig+Hf5NSLl5TZ
Yl/npNe5Kp3tOg08elP7ZrGQ/cdj6Y8z2gghDj5x7ApXO/WsANcnaPLJSaNzw1Kq6lHdS9/4BuvM
ofO2Cw7Dj/LHHaNH2FT10vgMeVWwHWHQSR8hrKIAR5tEzRSh0ncPfu0zcb4d3HEpESJQi/Be1ab4
18OrUCslqcJDr3W0Okif+G+pSV40+YEo8kOZW79lCgLVKpP1U0CtoUegudbJfp2MwjvhqO0vKNcv
juwgG3ra4ngAbptBV8JePUcqxvKwUuk/JEtcfW6n04Hheg2+LDQNTVWEM4GUYw1Zfu3dyF3Txija
41rAMJk96/LwAf2ClN0L0etaeWsoWe5KgTKfhnFMlcXsVnQRLCD1KhuEf7rIeLf5lH0VvL20eSoi
euIbHtVwlwWyxsvaf63C/sEho221WBh41MKkhz4+hqtSmRI+VnGNO69tyO5Xf0TJ+2OZu6Qjsd16
bpANm2w7MtwUMY83IxAxeqkZCM1BwZ4yvZ9lyGedhTqsPOH1+tDrLndLu4CBK3tW7mFeH58ZW4I1
1JTs8WLoDNvDWU4BaAQk3y4y6G8uEBtGSjauRcZKY4rmY6ppINVL0aSqEWZR4CBoM3eXsL7dHUQE
KgLyuc7SGQZb1liIa9m0jkIt7DOxdx9qJ5GM7mNC6UIiFIARQErtNkHenVlILwc3w/lNvb8J9N6M
ZSZgi8rfGHLfgW51DzhFctOWWkwWlwwOfpeMjE6KLTmf4WEKJLQlX0qdtQz94GVVxicDdsmYLj3j
Cx3Tok1zA0/Ui9BFUUKK8QLjz6D2VdtAKD1sx3kobubsK4xsfqFdogvKpNHz0XeHLL4mbC53uW1t
JvFp0RRvKxOxeCkiqjUMJU67TBrN6jzmyNKBl3Ru+MC5F5pR9JncviZT6k1Z20Mu0HLH6Zym5oHa
u9ifCMkNCGLOnjJSvTCKGeC15Cn/E6SdJ2oJDplVl3UDDAeZYlx8wkmDfKcC3qshbAGCq+v1tbJF
4ewupUYSCShDazhtRq4sE01vRDx11NdVX3Ma1brWaxOqRIdxRUoXhk8UWM/O4XpjDb72eUhDyZXp
kHui3H6b/uNQUp+7sQH5voF8xGLjZR4TdJPAFXgxc3P4aXk809Z+c5+hd+TeNbETxnKGkxKalWen
tN97D9HRjZ1nBXmttn8caalN3xTv8b9Xi9Tgq2l5VS/bFti3A/AMDtAtsbNR10iwAxX1qei7p5bi
OSr9dRHrW0CVeYWqlEn2z2/lq4fm581g0k0qlp3Ei1fH2czH38ROcH73gwZK7D0ehfdZMeWyom9S
yZeleX0aV9vP9xPCSezUTVoTPrkJk/R/OpTb3VNQmSfIjSMm7EfT8cNDAnH59y2wckjz5cTbujkg
D3TtvJYieU+sbTjY6Y62/FnXJobxr/9oGrI2w6a/0JuUaiK+7vHFGLiM9MInp6Y0oVfNPmMjawkv
t0U36/B6udWWdpll3ea2JU6uQ05MVE66V//7+3B7UOiWzLvUyce2/Hil88qmhtYqFs9/K64uBTFp
E6vS4JKBHqgqERnHl6A229vvVJSD2IjNUZL0HcCz3gmzZPtir59ZHwKMlMnDj2RdMSVYaWIupv7f
AlauXHKXb50FJdwcJz78Mhbf3+AoGKsLRrWNx6LmmvSNE/Zgeefp8UTmHTxzHTd1KoDJCOROwq5Z
q/MHfwJvuPtYbga4qt4R823y1b9Lidys/wMTpYQmsVgxUpT7rBxuLYnPKtFOLd2lI3HWvwmRXK74
Ub8jTAvgVmCInxhbMYm1jYdmds6mfAZOtnnekgB1DsNX83JwieLQZgTu2zhKDkX8EuklpbFgzZ4P
u36XRWA8bcsiL+fuKrwZ/mCu5n+FbFeOeLGFrHQ3avbpHMZ62tE9NxeNe61wUgPONjoXMm8x0SZ/
PTDOYt6hDoGiAg==
`protect end_protected
