`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dj6S2yIo/vS9OZjRj8p9iOfzKUe1Ge60SjGnLuqXhruMvT3ZQpiHBhXTQxqqoQUK88zltFxwIGb0
5taRe/dLzKoH+UrKsZP63L52RB/ptV+3wjUdk+qtSNYn3uNeAz+SdG8YXnIxLmJl8ye1pSzK021A
8SvpbJ869XoGYIV3RHl7KOmpHwlSa/q1Yj2aNigbezbafqKeVyXQwO4XU61ZC7mR997J1MtiMb/L
cvstRgkmVRkH6S5xLIX6GYMwCoAJJnpyKF4OJz0i9BmX30gaQlWURr773c0zPRajRwfRR29jIMf8
r03KwWiPhaml12Ki/FkrFUwZObPVCTJ8VnYDVQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="UMBFxcG5XlHcxlCeakUa+SvIdCEUQXCryYrpw9sAXUo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62432)
`protect data_block
GtxEnR71BoqNtyXyoh465j/jIb/FEaF4bTY+M2CyYNJyQTkqs0wpE7MJ1yMccVySUvV9AVNi58wV
9BpBKwwYxiXVcpOGtsA8cf/8Ijp4rSXWvEyLlnHv9PuKGpTgllvOdzvHJF1jofUv80tnoIbXoJBQ
vpi0lmNp7HDZKxz0LR00VBGpEDNjCNI4bkt1/XXj/CZgnqei/6TzKilplW/+IWEYhUGBYh47jagM
s/TYvkiw4upDLd9kWDadLYIBnDkr+Kku2SH+ZF1i1+qW/0n0JUPFm/Jb0GN729p6RgVhoPN2Oflf
00Orljm6427v1J9zI6O6T2roilqtESrSQxyqHh482VqaNB8LqdFwvo7DfS+/wvm6NMg+IqUm6xPk
NDB6UXyrBnuVR77QGtsgmxN4+HHgBR25YS1eNINlAsJe8uL/qoy9ncGg7E3zwxGsIrIaydRBWTCw
oxsfZpToTNt8oYYkrIHtZklyQgJCW+8cxXNi2RsEJrd7wx+JpdK/eSmDDZnPKH446uGx81iV2Chl
xFL+QE2a6e9L20JbfC9U/v7Zw1J0PRKF8zqLh5Zq8PJvzroZtDCJkyk8UtfQ9JBiOndbIo0WEQYQ
HM94eBChRCQDVSP9/sPye/Io2SelalR5zAXHi7WqJ5FzCJE9MvzdOfaj6sn8DP6tyAOISc1KiFcp
ywx8UrEkZABlfhZqJxJp0wZy9pzzJRCu/z9VkCRN0znnim0D9Mu9YHn/I8Z0sLqBtimSZ0+37d/Y
qpCLrLk6kRP3JiIdLba7sbAgk/OqKVL8vck+UxUey8lq++0lP44SJf+G1uv558A8JET0aMDYt5ac
gSUVAnOcVJaBHhRPz9dp4hAoxv76eMbDHmQHlQsSjmOFyBUWrqkW/j1iDWH3ZKALOIWHRDpIBw3U
LC9uTGOQ0g5ms6eNgDSbstnXz4VuM51aQIVLydPRrocpMKaTigDknHd4YI3UD8Ih/OTGKdWmfh9S
OEAsq9CrTebAstT9pYpPlCHOwqXwFmSijt9r0IzhHCh5/8o0A+Q2l/keOAPZ8CBGi/g3bXmE1xO/
HURrGaytO5U+V08ha9IAI0Dyn1k8IjvWLkhymJ3XYV1W9FEo1ktaOh7WaYEwzWPvDe93JTr/0NAD
hpP3/X1txM7mBy0Wmd8DAXVYgMT/l3bONd21mQ4bmk3uvQoyvSnBbgqVXzoh0ZWxVrR6SzBrjUo/
SvBL5Y4qkFIQaRmQmv5bij1HvWcir472fESdvyuFhohzAfDkdL+1ogicbpL8vV0D+Lg2DKlBL14m
XsDoweglHVN1tw/vWsCW2v4kcn0hO15QHfXilG5iK8cJJZ7NAXh0QMUUFSMuC6BSYOOoBf3MJqdf
MaEa10+62F5LGgLhT5FMIWcmkKvSRNf5VyIy3neEDkI0YtXyFqsuNx//s80xpD+Mkic7TiOpPYJF
19tuMp68mf9NBgnwIOHLMHMgS3V/cPZBiaRI3b2oqzuNwtY+bcXTQxB2qcyNfzxAxTSWoMg98zlA
UgF21AVH9CK2M9+J69V83qNThqc6JC5JYYgrf1lsnhXZP44jnFquTkL1LB5za1wwJJ7L0oAYKC6j
7XOHliuki/UYYzwwVPphQ1+TeCi/bCjrjmqEKH7eBuckEr/D5Jag2iiBH7KhpD/PKa86skVtzU3l
dbyl97z1JtIV5UmA9MF0QliNdymNg5QGP9+E1djPwy+/Z2+EHNSAii6hBB3otYX2UVSOPYLnEYuU
9wqidgDHoaCUXW+0NditRWkWfSAz8ae+esGAIET/btjr3gQzY76wCT5O7K9tTBK5wmz3uLw7JGra
vHN0L0c53SKIndbVDQOkOAKFswilwYYRoUwv30bairgBQzqOqVsO2JtsGBgbhsKdkjJnq2L11WKn
MfE9vD+ERS10VX2B+AX8wvuoA/cVlhKvyzQMlAGTN0+XLyVUkul5kLIqCeJvXmE7JMo/xP7oniph
rDYR+OTJf4gVBjZxXxH66FZl5wzl2N3PWyRMepFWw1io002jGkcqRx5BhrU4ocS3wPNhebf9C0cT
hUtvtmEWOuzzOYsHbR5r1sq2ExBxeqLtjFsYdLSQdkLeQMIC3sQdu7cUEPN9J5XoeOdlHX1Hqn+3
T79ZlPCt/LLl1G6wM6+C5FhhWcPRmEMXm4SVnt+7c70GMASD9LFKGuJIZ4JX3T18r1ncGeKEdE/0
qyqBLxT1LSJLEPH5w1yafVfyAdWFBzZQ4NYVft+igmOd/p5M3bmqKJMl5su5LlRcUw755xYG63VG
DRu9nZSg2TDqV5MXm9E26HJmQi+pIQIbmvqpFPakU1oNBpwv0rg70/4SdrMvjLTI43vJo9KCa7u5
NONiVy/7B6QeGVeN+4eKqHzVNhEHmevy9s1R466GlvGCQkixY2xn8RhtynBtt0h/pS3VD1nM8zlT
PvCQluHX5/u3905Z96sNPfwrKsqZNL1FDIPva6pP5CuuXA8MVc6VG/PC4a6BZgsIaI7SMcA6xzp4
5ewa04JO+382qtpYbW0sMWdH3kEtwgC2gytGYlMFgFiXFiKh/0MOl634au/eWkWqY3P/vXAX5lHX
B70q6HBc/LMwEFT25we91K4jFId4veVp+RP+43AYSYY1rk4M+zz+5pZQRxIeyYXusfEqG7ZA0LLC
HRxl2UabET74KmSCIngSk7NJ6gYM26lNaPNLE3b6wBbhW+JSeaUTgBdR/lG/TxvXg+VlBaOaxpL0
yqx5pogDYF9HjezeKymEo81NntowUNX2TFffvTGk1ZmGlhUtVb8paLdDCODsydQTop8b3qwVkbJm
B7b0XCY9pH08d/XaTo4M3vJ8JCswO9mIOdHCkXo1RkPrIlifYT+17MFVEfHpaUqRzQE+HriHYSkc
nYp0mLY/zNxbTiNU/tB6te3pHP36TqL0ivOZbuxOzrzidUtTVSPLIEskYUrqgRxsXEcIMMAX2Qv9
GsZEHx7blYfX2pvR41E+1bWZeDPvwH9fIrxLFJn40TshkorTWGrjAX/MmVj1m9nyvlTB7yFiIBq0
n+5OWqsYWXUrHjvTeCEAwEeVywSfNN1Fn8T4XMtS9k85VquWoW8BBh8XSdiUxlhr/V+bvW87yCKX
zzcvit0Konsl530dmosNbWyZrORGFXqjMu8eZ8wHCetwKXRYL/TkLsR9wqimL43deTlHWB3U0iH3
FxLICjfuU1V5wp2Noju6ZIoPKqyHvqZ41OVOV19L+cXeBi6CS5+MqVGtLnsgQNCB7xq4rGsGieVG
KHYqPj9TNKS4lB0Or1qgxy5L+DS3I48896lsfYglD2uT7OiTSngLdEQiVf8TeuFvWHTl7wgk4N4q
nAsMNOlyKT/Kl1071k0U9BtWtI3Vd9bIH32X7p3HCvLU40P5dQ8t8m35qH7FedTYH+xPGvxpwFZw
rXwAS30hHVj+cxdgyY1efd1pBE7DhDxQsTCrpHXmtzTKNCw23joMU3BT4Kc9l5JSQmtjm9sFpJBQ
MqjNE2kaB9PqCNeRRZOL/Oeea4cQYsXUy1pp9cdRXjm4pq/cJuhZYyoSwV2NHGj1znR6dG6rrt6r
/QvqV9F/BqdL0qQmBjO/NFufq2TvJyQXYZgqhehXHNC/vtf/BYeftjDLlDE1OOpqTPAcs0vGWZ5L
0fBKg0qYu+NCLfEYHuB+OwteZxnv/4LOZRIdDCd2p0q6dU6TX0rhf/w8zc/gCQvuVJ0pGAWTEDmG
iggjuuQ5gwWUeshG6Mzg5BphrSt3CRfXH9zgzJMhBAiCnREBWFmxtRIXcxed+4uCNGe06K5xtjKZ
pkM4qOvBgDo+ViU1IAO1Nl9yv8o861fC9HAs+rGheiIXt+NjGKvKr/JQDG7ULaSHpjbfCpCvTlkR
L1V9JW/VlostLNXZv+tFxc2tCkqA6ctepRsIF4scDRNa6KkZp5zEuG7wv9myxnetyK7N3WmbACbq
DnRTe5oRsv04BNQhtiTWdzNxxQfyJ1p7jw3XyhGrvgSZ9A/ouRvfnqTFy8X1x+B0Spqc1YK6r9U1
3gAOOhwQhmN6OI9mxOiHMs2bvovLKbdD1aTkkDwcuxyesS3foyLPGfeNlSbGUDcj1x2pr0qhMAm4
giHOMvDSTrQXuWKymr9//yNj9/lnbQfQFDsXsjTq0FXfrP/ryHuh4b0sJEXLUGZxj6Ih7MIAge0e
RKoFd872hqd1a/lEeHIydelNpJnH54Ch086fQhcq2WUAM5KzqoSlvM3NrRp8gJJBP9DsiTScaVUW
xQRxfiHfKcOHWV4a45cYNQgNsIRoYluPxIS33nOYaToE3WBuPIpOkHPfDz3maQvpD9VQ6kwSJHVB
6viUpzt4CxLcbw/VqtGN6S7E0e4l+EYJSdgwwwMc0iNafihBhLW5tllu8hggynTxu72DeLX4YxgW
RUPfcgU2ZomqBa0Ni5NPnqXxoXanX90RcDYe1lR9RC8Ek9iuHzxIjn2Y+VrsbMy00hF7WseSaQjy
s3W6b8G3Y35pQQGVQAuHyTMI3GZOOrZijkAkqFbsyj1vZsV3unyBx57Cd8rpMfryC23U+xoATU8O
JCR8Gj9tXrR7fXIilvq5TgirIvUA0wbN1WsaBW6CwGObBEaXRqJAKnF5cHaqLmpTrqz9DCNGzSOv
EkDz352ecdyfHU2QetQZDEPTbmIGw4YOFqZ+DgD4T4MKQSJbeQk3Lp1zW2P4HcX5bsfIZkRTrRAB
MSBoYXkPzwJ5YKFClrCA+lbW6yU6QnUcH7qn3ulBr6WFKI6MbN9XDhYqfBOsrSG5EQH9MgwvMl57
O3qT9cAEWtQeEVn9ZhrccEQBrlWqriO1bK8Y35nKtwEVcs82pXJUQLm71WT3Sn8+nEbY2mcP5oKx
FeLU9dbst5jD+3LyJ9367gHtpOM1lNC6Cp7ageXjdZ0e76A7lZz18fPaat4yCCDNmr6XkX5yxMzE
+nU/zUfTHoqsaTw0iPEjCcCXeL50EWScEcTBgBqHlXsuPchLQmAgnMHBtQwgFZdWgJgE9BH80nig
HU/sbjI0KCMTF+oxFTJAOxcCa4966ich+rs0swzQ8kCBp4Acbvo91NognQyb35Ga/cAKWtsqPzTe
a3I9OXXjgWeO2wAusmS7Nn1Us400VJPzZsbe0irLh3YVtCfgKZJJy4QgrO55z4GTAOTAAWRB3eM2
BLzY1cM4MfYZ23Fy+9S8lsG5e3GFC4EtKfKkTmauP9aFWGE61qTE5jixvTTP1TChjToo7MfU8uuf
2BwplINJL00dwb8aaD/6RbWtjfRCuOkKlLdmLRswiikdDVZEKc8iO/uOMYDbXoxigcMDM9EZTJb6
mGnG/0V9pa6ZZbSnJVUesZRQ8aOVcfI8cQbyTRIufFz8a7E8wMi7O78Kl3lYKnCB0ESUWUKp50YN
4cZqkIyKDhuiv3kd8rbxiniOdhBmAx9BG6ADGxo/UxyEdMlfqCq2sXgtjRFxGYIkBt0TOwPeUgMx
6YIsOOkRIZ+iDNIJ571Yqs4/jrnD6v9kBYXa09XYZLfXObM37RF4tu0CYFXrOTcA6znNqgot7z5L
FSxt61DlfxRWB8c+kPmPlRhKU0zFQpTjybLgr8jXdsNlN7tD+YmQ0Ou/48KdjpUEYBlIvB/7/Xju
OP5M3+Ybi+EdNG6sDdya7BKbB5K2BX1hYddlBZ6uABLk1tcWmWDfkQoaSZHZaz6Nz3oHNIO9eAe/
T74IeyThJqjxufPAaI3bujb0CGHYyeQEbFZvAXfSbMad5NDuyMBaDrkyR6d6pdYnGw325bAPS5Gf
VAalQWT+WAOgFa5zXR2HaRAInBE+swDRonmpRYQXslM6mK9ceXO/bPEEfz91rPLeYEMRtyXsRL9n
Hx8csVFxi5eSekzMsEJ06LuoRPXxo1cxHqaxhHPNpCjbXPCJaD2a0MNf8gEClOipcE7gHTOpMhQs
jWR1dL1WOj2pbbY5qRjRuoUKagVYgix3wtuJPCkXK04SjoJfioZHT+k6wqoMT5j5Lwt7ya3/Vs5v
CYOIxhexlYKRr9ud8G+bXeXzEVJ0nYLOwBygvsmjCQD0KZlSR+oYXSVTH4nJLO16voq157+cT7Fv
t4AwXc0OJ4qv95g9X3K9OK7uklGNXOZdrSXM/SOCf/fFSt5/oBb2ZGHfL2BOsbEcegRyMj+mgSuV
DIkj9oRMVlT16WIFKzwsCKWoLSkCZFhw0FA2vr+98FNYKWztFzBWYe1LlPLLyWrmzAWYRzchsaFM
kJRXxlDQluoYGUbn2LAygS3R6hwc4OMgmFCJijfh5nR8mWpvCeyPpz0QLO9SpkEJlcG9dshFw9j4
a131xfCDtG8sfYT1hbjxeZ2FelB2SNObtOC8THLnp1iPqKNtDG9S1vLQUQIE1WIo7j3VUPGB1gUw
4qaSTo5DBmXt5fYWCOZfZsfP5AOfj6XyEEwbEaAEFvjRirV5oOz/jAI/uoVXUxm2KVTOXBD5azKZ
sea7A72Y6cCWHoKdh4YFVbFdTMgXFmDzSh883jhPiJdwDo3HAac3mhcO9zRpbjn83WScRdHY6v03
Sx5VWQWheaSgFpANh8RX+kMY6FMcj/DdEA5SYbUpRhCaaiIPDXSSNJSruyanqS++7DZ/bXOuB3j7
ljthzxEnCqxnk7be5o/zjuw8YW7yCtM02pjDyDeBNW4Yj1jdfeyDCwn6MC8svtgYp0sjzSO3rhGP
3eoUg+jx5sST9WJHtPghMPnfcCGm7y6JnvUIzVA2uNT684bNeKDSySGA78KJoNSKomS1OzisZ5h1
0zA9hxmT5ihauZCOGFygEdADeGaD+Ws9kyCbr2t+pl4WrCSe6dF8gqblmd9nWIUyYyEx3A1TbRIY
j1zrOlrjoWHCEUkCq3mEYlSV6GGTSAnyxlIA8StOwOSVM+CPviPM7XbeqbIt4lPV88IQzfqAkzGG
4XOAyZhmlLs0aNlCSrR4tTcOkUZEdXprVc1BP1B84YzYYITHB1gfrKPJCGB8rgHaHRAiaamIqWpQ
kUdQQZL8RVHqUqw139B3m2E3jV2qOhy8qJBOg/hfq4RHuXRuKRas3mwOSyRR2KiU7bKs8EAtJlpy
bBxGltqFF8bSHBXKY8tbNt9qzwdKHx0YWcnz+gVeG90XRbJqm63ItzmLdS4sIVCMqvCjtCCTuSOc
N0Yy/CtBauQRRdiwcVLM1rZKrsmGlXefIv7M3xwdJYfYMhr+vmwk6s1NUuyCVZn0gpiPcxGDWFrZ
pZD44hTLTClzYL1QbDGVueMOjsrhp2ABg7jAB51j2QSL2yeOvRdF7jUEZX8/eyvw3p5t8n+WfMJe
gxMPQ4TUc2ywv4zln2sUmmm2wHL9j2lQoPqhEnFNWAS/wau+i9m8a/DU+SDosmXthzTN5l9gEIAM
o2K1bRoXsyMiX7BoK3uhDgEOtg0BhfwN7GCzJmWzqr++XLRl2h/LWS2NIgM+LnT4uAUON5ABxj1O
oVoxH29xWv4CNroSuE+MJLnuZtkeGFEP4omdvswzNT021A8Bpl/5uvnHBnBarAK4T9Jy7ZubRtwQ
4Xpms71VsfvqQtdmdwlUpCu++fHpG0bSZQQhVcTyEhgWu8mMt2nQ0Dyx0Iyy5usCyiBmJ0XR0aWI
XdTPdehJQrq0z6gRPzgSIUsUS2FXSj5UQ8ibhRxvcfQHw6LbF8A8X1PCRRhIfYsVB0HwhXWyimCR
5FoC9Q/7Tk1v9vxUbF0AhxhAcKfpf4DHOWzYnleOQy+blPxI4kDWwlhCJMKvmwQ96wlVZxmbx0oy
VLIj0ZqGMhMAwCsiXQtrVhMpH/gglIwe5tkPLmMGvOy2wk7SG1fSG+F6M87pPxS8Uejpx4NYw5fY
etqClv7PIKMWTgHYW5bBhwb6fvG/us7d5P7evIJn5gsg11ZtJKsndFX4Rhw4+zbg29t3EtKJogbW
7oNP3hWgpw82S6bVngf9mYCttAZvdiiXiTpJ2dlJ3BVOqUrKC25m3hBzYGaCdBm5xTUtK2tWuaRn
PXp5VwzPHzZfiDPfWLGPn/QO3zEVEa6xS5jkIU8naTw0FijivKDOcbpCGvPCVUpNKqjkNA9pPHTt
C1HawChEra6HIyhxv4KumRmlNoEhC2FaiWs5coPIIOrvjKozyjScnY+zOy57q+KQbk+DeAQy3uqL
zTWYGdowGHP8rWv4viQxVNCRbhP1fDa6ur8ES/xMa2CnHi4KlDxtF+4hrQJ6ZTTHE7MwSMVXoW4/
F0JXxswJKYZFJ3PgbU6O9NFs6GkZ6l3wxAWWG2cViU5qCQ0oE7y/4PxpJIu5bJjzX4Dma+xghn3v
CRk503VgceTdMygAmPFvs8N9IUcdCSGOl9K0Kpm2VhmNa6PISpokeqTy4tcRp+BIcC5ZGlQkh/EI
N+ABHjxNNOJzaDOqvyrww/hEYdxmacKVhjzTQv6f8PJZyCd7dM2srY9UnNzaeWlKtedKgqi9SgMt
QpwpmC9btr3HJ6mQbYP6HoyXUwA9CX7ftfgDX/Pyg0w7PbtYTfytV/o9mGz2sb1MPMpQdAdv4HcS
JypiozMvshO3mSW7I79l5ABQxvTQS9FkB9jYooWRZsNZYEuhL2B/TKytZkmT/sm0WTpt7An9XzvH
MM03NJGKh1mzjAHT+QuWJVxTJLnPjIIKdoVIijg46h3g2FddTtZUa+bXaehkdnwPQhwqhipeBOZv
SJhlAEUjH3aphpH0ax3/x1wsPj37qgaAdK/gaPiPn+5o69++mlBdvngtTmo+sgZLpWiNDBDd5r6c
4RZYBu9tuF9fYTBWFqVXX1UcnhI8H/ATLzVtsgHokoPM+QpuuFZqLQCEVJOeY2BkQDepTic2xMZa
v1dx1PjnSALd30a4GHoLYUvjEoMRQZZE4reVh+b+3yhN3JE4VCyhcPjntvlu0r2P4sPvf1ReRoa9
eo5WsvbEWCsq0BZ8u+5Fsj78YCsc50QILCpvY9ZXRRbkHQpTCd6ZHITObNEplm4YJaKTc7bXMux6
d+NgeNUfi8n5XHyNcK7me8Zwuj0x4HJsYUjmsAE4iKBANLTaZXX0tMEmTjiizlulAkcEvbL/at9L
p9119KzrvHUuMZ3o0CMo/d5EDorMTD5uELB4xrLytQggv4GM/9iuLAql64cHjkNc+sF/1GOsGsCP
HzwPLNJHAZIWjT3z+Y33hxVZxnxE+A4y3REvaqBWNhpJ9fI65QDIcFj3JQoVcEBF6+YpCSwBJ0MG
jOXTkDWof2xZa9vH+zpSgD+XgT6Pt9Vxa64omNLQ3XBBsoYVLJYYKg/9Ln8J1vv+SjYWfxHa/fGG
ipfAU9t7dzUfCkTMA1iQH37n5KnAVhuec7NIiOCH08sWrFiQNBoEvvCIcRXez9g6dFlYaBHkRJkP
lbp2HLUZ0e+8GX3z2V6CstPl7lUOK1MqedRqnapulOktb/VezsyQ2ZpcjPpjfR1MbuUJyYA/OdrL
ECaTmSYafe9MCwfuHJsya+Bgx0ru6UzduxXwWklyfkY8fQ6VMFXlGuxSRfE/HoPUXuVHJhuCLR5s
inIfR1zvkwK6dxolBhzxJBRPS8W447NER4r2f1+hTHlErFPN/9+x7KdiXP/NBcWnp1VxO6x4bjSu
KI4Jqo2T18OXellhdSZarOSsyiDm4sVYWLJIZrv8LgG8m89WhfsEXJb7SQXbm1554Q3HZUHoPy1S
6ydxegK2/2amJDFDeh7w/T71HRX5p1T9v7ZqKRKJsZUV3EcfEwDJogNuMQX80pnvnq+inUZ9Hq6D
8wjJ40dZiVoKfVlOX/8zG5fJoBmYw9jJzlqzS+lTmB0Xce3mo5Klrhu+k+GFLxG3s36DOcLIuJrH
OBl2aOCn/oKWViaOg3MvCmjjjUZV4Zq5ch+LrijLvzgTriK4Y9DzEQ1SMeqOF21lYWxwMPvR8Bab
mgPl0ezAPG92CO8jZ/ohl/KLZQTb9vZ3Yc9Oh9XYQ4F1RVAh3wYcAmT2ogGpW1ilIUr3b5fAmhXe
pGLJUBokzkD/U23NZbl4dQFbisUPIknZeh7bb1dMiWGyDpK3s+8O65KNT2DDZrQVyv2Ie79s4SRp
258QF7wLVg65bKH2kVpHU2QnNKYtConuj38uY9FN1zUhfrUugFpfa4VB4eCEfWCbRQeRuHqjY3og
b1dX9HLqjjamAaGdxO6Don6wNGLkU27VAgVpKQuOc4ykFief315dnfptJij9E+kEIm1F5aF4LgQK
lG5mJVug3hje++iG8lOAjv9vZBSH+FjUxE13uLIpKmeHO0B9VR9/0tiBtEPOntvoyzzfvVxveOYw
HdQi2BwbGtKTjs12VNLxavYwle41x/rDRec92cnkzT0ZG5k39e2V8cDcB7iCaO3KVZyxecpx+MHn
VjUHOKh1ptQP/3ouxfR4F6nAm+WhVKUfnvr7K3Hwl+InmHcltFvClAVM9nXk+GwSDKVNkwbwoJmt
ud5mmKxQLAgJCXoo8kUfnVlqqlfW6RwLGsBQ7gyV1fCbDpUNlpxACMYFwAGbQv7Y3K6WNZDoZ/R0
Ue7xKr5+oYdlVqDy3Ab5jn+EOwsv1fjcxaKAnBclQFzfaCUW2xhPZfkbOb/4oev4OeTh+kPEw3zs
tg/f+vGDuo7VFvrBkUPK9osr2lzDCPyIKiPvV+4473pNB9UvxoD5GgyDhMxt7Qcu2U7+4rRkbCEr
PUe3N2dApVtDjvQB6+7zzridaXvtPkXW0K+YkN1Xz9CiTLP8bHH6VKpbHCMyOWvfIxl9L4iWBSu7
tZeKLq+KUbv/R7L7HyzHO8RR4s6IrY//UYPEObuxplozEwEqT/HlRdVy633cXwdP53PvYvv65MGg
uYmf8jNOsUbUAG7ldT0lJm6GcAVpGttZw5m3R6JfCXCSlw/MDBbVSnZi+483saD0JRi5JiGhqdJj
rE+TlHXWpPRXIBiV5DiI9XfN1BSs3ntJ2NgwqSh7gRdp+Wtq77YucyN25UgmXtSAMfOJpM/GbUEz
Ol18/dxX+qzwko4g4DEudNz82c9RrW+Tmt7WDDryPM5/qyG6zsaTJDD+1W92mTQC7+PN9qE9HZhR
9ZtCNLuEODnDYMLOR4BMRnec2uzRRMU6TgPkOrsnp5seu31JzevMYMRp42/htySi0OVB1sxv0Soi
hyOspwVpm9pq1DGX5lkVcnvNA2JzQsNBYxA29MzWo0pVKVTn/y3ibOVeXfbjMe36/Q9vaPwl5fd0
fFJyQfmBDvCzRhGnVKcinlUplZuKyQ5MVxmk518qytrk0HuSt32OWX5FIGQZK7D05lEn4K55+ia3
y+D59q/icKYYRhW3K/6cxZ0Zyw/peLnMCAbrtogbwCKT1TLhPdFvaX024g8UyInHBORQSd5xP/NV
6lWKqX/S2tuDJ/RM1q3h3kb02H5t/o9RF8xOaGHEUtZRaUR+QxvO68US8lIZ7qXPLuqyG1PtbLp0
zGpIO6JzkxkCyR9WQoKyFd9o75y5zd6wo/Dbd+cyqvAJvpr642xHvoOSzlRuNBLNVus93wNYYn1Z
O0q/jJZ+7rA7W8jwSuAtZ7wUX0bWP6Sij76GxrIUE/Qryjjhd2Knk0ao12BCwFRJKavB26RE0vti
m8TnHMhcSaRGXiBrp3TLayb2vj8iCaLmEWQ/LgO2iSGBo5zl18YM5AUZYYdwHXXzXwcgVi/yYll+
dD8pP+lJS+qWzToMfB7+8qu99G5BbrjnX91UAbtMDI2bdU62kjYB4bnzbEgJaOJk+h54pTGcsMPR
XMU8TYub+ha4iuWybatO6BINZacLTVbc2CS6WkKLfWd9b7OQq/JXhlkBoQUyyVNxP+jf/YtxAAhq
gqYtT2U/dHk0iQEOPvVvyci16KM/OwVz+y3Vi6YwpxYKsoqBtC3Cf1Syawf8dLz4NjA2iYuXQ7LH
5T2YBtGujsqlh3c1DXhqDkkAUaN3o3zmmX5v80dhIaLfMDTh1Dr6j8wbZtMcoOSzm6QhmIrLbiyH
Xcy8g5YszMjXDQ3dBl4YRxBZaXLRcLkpw+fh6PeQCKsUggovecCzJ3p2O3t9NctuzV6Ll0QJ9bts
NMnvjs6BVuwWlQgw/QmHe+5EwOkBQsK3AkXjPEeYDAPKn6Mz3c2zeAzFYSP0pyDYziiS1tOtc+83
KjXHlC4NhY4WtIMWW/NvjSnMaNG/w9KpjAipiQpb0CfXYGAlweQNgFVWpIytLEkWH2aCNAHwB77C
4MyxNs/gz6E88B8xjqju+rx46DQzcqcRBvUjEHoYmaxAoeSQvEZEmuxEbkouR+nF1GB7ntZmXMow
+RruPj3quR9t0flF4eYh5RbIpVxPeRCZVFNJy6s+aLaZmmimdUTgIenFudLBguDZAYhavim1FN5R
ImT4+FbXaEYfRqj+Mnv6ziYEIP1LE2m3FPzwklLOmKlx0OvGqDt5S5B1yX8MPn0+LjXcGM1aQpup
NHIZ2I6UWeKw0gS12p020iHvTndySuaYqbZTWNpECwegHlAYbtCrr9nKGcxUS3izsAdDWParu9l/
bEW81tDTuT7k8AVmlXrAA9nyI8qTsdhdgMjqYNPJRsNQYJcsiRdjHL5DALzNkqjl6qnMrcV1mrp8
CiLHmlHhbl6/PGthAwgOns/ouOC3DXmzGFW1NC7bPd7qTp8hXYZDzMKfnihnIZO1yN97doHckZGW
MGocV5V7D5ZD7xM3j1GktGeeiTDQt9zyFlQAoVvzZ09QN4S81a/Wh2T3AqX+RQ4n6WWRpRTpc1Do
jeJm6nRFoC+zD+llgS6K0ocoRl0eYudw19kFk2Dhbltkp2Cg3ZheujcDGjUnaEJaP/V42RwPCUh6
A1/OzhBJsD4GxqvqD7JDo5WxmGg27fNamXPNQjE6t6AjBOG4Li8rAUArR0FuaImbyVm/5G0DeZ8T
pa3dF3ijbnlNf1jvscPN70hWhy7TuWEW7Yeek1qDspiRrdHXWzNVbTVdpZq0aeSQoz/Ryd/VWudP
jLMaoD9gK8jWxiyHVnDHYs5h35zjfn/djdGGbbkQrWh42/jmsJdraNBCtjlWR7WTOED8MrBqC//5
DaboCl1DwKjZHIaKGcLHo9Bvha9PPYJOdFYZq/AOQ/ul/0/0RAaQutiLUrecQH1moS8cXyakvAYg
qIigLS9P6bWmaAdgygxNJzCHFhXXAUKMk9WTECUQhNQvgCUWrZE50wkbq7aBfbp+9sMI+QONhiMz
+IfKD978Y+00FnuZ1OsjWFAnHi7y9j6pmTnKdXrPKMhFK8u8n8n4xqeHvwhXlKTdPU3MmHAQFf9c
BQ7/dEw4Ol8s0qgqBHQI26VAC/xRgNaqnqn25lV3uipRZIPpqAnPlX2p0XRZVFO15E810he1hIys
qQI+eRBsrAJjzQCymzKfcacEbW6ehrGIHVdH+qiDpE2nKk5/I6qI0+CyzUcrjgogezkFd1VU491V
5h0hA71Ntq4+3/45tDf2P+G6m0BVsLH7nMc7IJyBN4Zeae/mgsywg1jLM76JcTwJT9u2N3mTjgLz
bOEB+YCm4HGty5mvEeansTdqe4yrodYdz/XzY035jABWIHU7iVZaP/4SeOX05SxOrvXh6mAOGTAh
NTrYJu37UimD8LpMDAqkXdLYNv0K1MZudwmcZowI70aG9Z6JeJrAoP7X7J0J3iMFPDINV0rG8Taf
UvdNdC3P5DzSAhVr+JJaW3/U9fiDc3AUiMqx6UiWG1sBpUf+exHEMZzJq8G8NjIcjpyIp/QEbvOL
3cz44hZnBqlXDf8lEdZIEfpGM0fCNIE/OOKV2G3UocOHZ+VSqhsdjlTpcWx0olOXw8PjlzHRA0mZ
c+8vz9uB3ZxT1mzLBPp3X5u9gWNzUuUFDO7G1bRI2ZQSaiggkBNh69pCEUwtYdOnBBcFq/UsBEAj
KG1L4Fohx14LZe3fJPtUic2GFgy6IJ+SQTbXu2gJ3xABpZslbVlMYqoI54+m0djUAGR70+FjUbl0
i4JTp6p1tAr6+jLT1IQN3BlrXm61LTHfPDba20jm8g35bX8Db08LvHRo48nz3OWFwoxmhgc8BBQR
tFBaO6jl7l9XeRfxs3I9gEBqZsvDDtQwW9H/yVVWcSA+T9MqW+j9lDU4E08EmdEllUmKB5MZboh+
UFnQXN3rl2J/57zFRbyzjqNKQ2gh9Dci4DvJ7cSIW18Kqa9/fCX4/NQA41vTbMgQVBZtOl3dN5ig
MnCaLb+ym5cVLBDeZi8azk0Aacpqi7PXy8hUhslLoJYylhpcDckhKq/yt2gaD9pjY99fp7DkuAD/
liuylICDUms+Wwht6epZT1etnO0puxzkph9DA5ylgiXqXbCxiHtQMCfMKJSk8ARo9ZWm1O9pMixN
UOJLF7AHY8yziLQM87jZ0ez8YDY6vbN1bX0Qp/tuwC7mtsQzGuUo10z4hHrJHv+CbqFSS3Gs3i5k
nn2DxMl9rJiTJluMX1AQP15TLH9msS5OJlftEi4WCxtOPjbNWk/eAvKRsw6wM4R48ftJ38IXdi4E
PjjnyWK8GjVTvjidwua4d2xlXLoZxgUmA9MSN/GJK2A96S7OPvrRyC1u0AOBJxlj+CvvaLykqo7U
mMpkWA2tb9dHC/unKhO1kGDMhV7al7JJe7eo9g+4vr8mzzkV36se9zwoBMhPlvnRZEYRzygCA2yu
+Es2++gItUyS+0cqSOnoPs83fps0ey9mGDiIm15MrN1C9qNJsX9tnn+eHezjBpc3KJA0et0e/LaH
uG7snLISTKMSBHESoheZqMjYHCg9Ra12rwod6YNBBCC4qV+fhpiRPyL7kudJcB5gFbnhaNVT70Rr
nOP38CVt/uNNHotVMmYIT6He9pIl6xOQhNBPiVSRft8b2b3ExtN+xHti3vlMNIC1mxTKgsQDd+nK
CPAL0WoZlwA9Fo9zWrdQ4rvmL8PYYIsnFZ7tCwtCd4O86QoGjWyJIDr5U8FPyX15dy0hHW8FOTkU
IBEGyKWI6wLeQUGD3OxEamBd6OaA/mwqxCTGuRVAld2G84wookWBANB/yjWaUO3Th1fXWb8Rnavw
rxpxEjFg4h1p2W7/2g3O2lWa1BRh+yjKAo+zuhRX75Mw1kHT9Qq1lzq2S7+a62jtr/SV4gO9eVBV
gGR7mKK1HZYsg0WpjDhDTqDxibK4NzyzcpowGBSB1TQC8g4oMghCUX0vSLE0NX+FXIdyxXklT2OK
4yQeERlQCg4ZKEBl1v4b9BLOUFlSow1rhcQnVUsskWIfTqTmmNr54pA6rqzwE99Hy5ijaz2Njz5h
HbSOE0wGZKPP9ajzOQAdWlcfGF3LOEO6h3fU4jV9+HppvhGJ/NTPeDSP1NDPQ5q83xL+kKykz5fJ
LE8YPvp6/CbevuRbbtaPHuYE3Ppq52qePF1J5xi80vppnzn6/CBmyhavDNR6WEhEeTXLpmCGr0fE
GCUAMjqWwnjEYLxO1tMz3MAkxrYwkAj4a4j6a67mXj+ad0vTBUukg/xLVIjPs9AyGgc2aFWShdAM
AeM6ENEu7t6qyoWcZXPgcFUY9L4+PI+0f+8LjRfqlfo2UYD3sbRNkRMY01ACDBLaJWOo7rYaXnQx
nu89sjLNnV6Ui9dWw5ZErh0ZDy0uT6QZVYddr4FEIyvrJ1NMBXVa/0U8Rq8ddT+s+mJILcGGt5rT
d6UrxRjmTVPiisEQ41bewnJc6OCwLdZIsgRE0hB7UMmYLneaED6xMIkogr8C5zJ6ckBQzBB6F3sd
4rsVUhQ0AGMTo9Te+LPm2IXotWWgJmEZkQvRHJOKoxZu9yerFPXbjlQR/k1bVSkJguDQI37n27jF
NXRGa2djzywyEjt6CAnHy6a6kRImLL8MUFmqunwNleRBwjvO5UVEasbUbVb0dsnQ4ILMMWJ7HYrO
DlP5xbJ9z0g4qYIFfbVxD/RGX2TjZjN96mi7A78kCk14FyIjYB7DYfVp3SxWTP/fGkscEBKUIEhd
E9m/KVXIYlJiHxbi7vJ3OmAPuH0bMoU1JB9fePRa2VcaRESDCxrO+FefOGc6ZDZSol7QGZh6raoN
UtMCKIvIQUgkQQUY2GjaaNQgk0oXYCFqz9KuwBYjRcN9Nng3Qr+spxI0oJ7F3Sa3MAVC1fSrT57K
qwE9eNHboNsNfkgzsZw7XEP+a+ZQT34tpcF3lpcCbya8poACLl+Sn61wNrDZNTVkdszqZ00XQAcC
Gc6a+RFhWVH4Res6qdAXLXiRruE97jTiLEpAfomhfdPU2uQycLJwJEmkiKn4wQEeaL2qXmMlEoMC
ZjULYi97YkY7aizKbJMrXFO0coAAo2rebpPDcjL7uoFZ6itUCUP832LhO4QgZyu78yg9mJS/Wv7P
6vCe1wCa2cGHHVEdgq7VPybPzYzCKIl+YqBotx+JuvQeTXUgFC43P6KzIrUX92LuXcxbf1RJi4/m
fyVtDNdk/tN/4rvD5a7KHA4yX02Gu1ZMbcqXd2Z4m8Z6C5xR7PoMJfJ9xAu+XspFLXqGfSVjMmE+
4jJN7uEnx+ZHjjgRD5q15+zfoprE5Aj0wwR9ldeOZU8ThRkhhNyGcyOsfZen2XnMu3TlZ4TeFmCv
/xPhAvqcNIl6gsPRjRJln73lYOY52tFjN+IFSB4sb8P+2O1xXobcsjqZEEouAz2iGsSynTnLDhz7
1QtTU61Zp0ERJJtKQtjpmt5xn0aYVLC3UVw6u3dG74ntds2ToV7qsAzgoIjBljDHJv2344OrbQzB
BHlZhLuHOwFKRWXn6hmxKaPlsu8x6aUioJ1HJJhmTurGrfwOwHaXjqQqoUr71FC3lXbtsH1mY/Tg
h+/rbn72+DP1z9YeEdGV9hXgcwrRwcFIZ0Yp4svXhgO6KvNQpLHHJibmWl2aGOB7WXPjaKW6BAtQ
bokA8p+iTxc2hcKOw7vBybEhSru7vscIGRskFhxf0FoXoGMqlGqvJQvTGzBVfsqEfq+fFPfAroVU
XcVzh5/UhKxScyQrYCKE9zh+H6C8DYWuTDTrfKhU3GyGwAA3anWmKCIqoyPcXW+P+irf/IwVC5Qz
el7SbvyqWpmXIHgEZaXuzuQYSQ/v3UN2VKxcyOA1zlMmwJSnxploQd7Y+mVaftHiyy2HggGie+TY
KJoyeN/C+KnADQ15Clvkbpn2jN5OjX1us+vFnYgm72+YA/joxlNC1M6zspLma8t/Ql2zdlDS5Ort
9Nu/89K3OBWJgBbEcdv2uW20U1s90Mu2eJ09S59drMy60ll2JG2zNnF7PL48p3XAGEKX2I+G04bx
j9EEt66Z2j2zIdx4a+9g9gNsX1uaQaJApV+64/TKELHuhpdQ0nfBIhY7UfSn2dymHn67OqCmi2hc
tt5xvJLHU6hFLOSvL1rmPzmtOO251PyyT8rSfaYsXFwZkj7ATs3KofQzLSP176ivkkO1uLKkEp1H
GTUklSw7wXjq9okHWzgiAE0ngIRZkJFychGsDEw18i6aRbkyqqica1mZjtUp9816CM4iYL0Q8ZXM
BSrdYozAorlhsU/SWXTpuCdzU6efu+uf9pNVyoLiOhErPx+nUPBCih9KLZURF3Sv57ZBR11gbsXm
vpZseIrcjvb9BUNoXDEWBzPnwnBukc2WYkwX6qScbKuOU8X1aFCKZapfAd1iiXWHnNrQBY60tlW3
3OwsxRDSpcz7q5dwwL5hq5gIu9J+x9KjpNed6mhuITB0VtsBX8l+PZ9mGOyZsfm1+/iZIc3K+1+G
Xz5J76LA2bdlIuo3B5Dqhi7aVVKqZW9oyBhEFK134lJYGKe9Abn7gbMuGjBgjxdNOwB8pyQ0Ofsf
Hey6Xthbzxx8k74Fks79ZJ/c8yNykmLPO5LZD4yWQ05yxVgxYHkWqxOSiZNcNpvL+ymZxoA7GlGv
eMOHBdmJCQ2UI3Ba5W0RkDsbimnN03xNdWa1DGESyNrKa6h26fVNirQNZj75gEzTvZiBUXrU0X2l
ZiBb69oiamk2auT4qGGu4SAGaRndrGXVDHxMK9p2Q0nYeJCJK4H7QyqQzRBj6mU4SF8bGF3kcjSL
31VX2Y9fNWy67u0WDinXPaugFjCLb+qCItzDOoMAi8jau8JwM/wCYxLIvI3AZC4IymQPPfklLb8Q
6cVi0CJkVbVqakvTGztVLtIh/otdiuxcUFSdLXgjgPQIOffntQ4SojpxcmkPDrifkIG4Ncb7uB+s
PD2KddhzQXfBnCiYb5+8kKAnJg7uQYNzgaAe66efoiIncf92kC/Kva7GGLUA3P5Jkzex/PZabSqu
ZQPVyJXelIRycS9chf7VplRGTK6emFzaWXscwymEzLpd7JTioWVgD/Gyg5YwKmGGrwYaBOOioLd3
FZ2UQwr2cfc0tJmy++OvMqAeA8w46kdMIvu8Xy4uzCHlaTpPiQIP9EJ/AWCz786RUcxjY2uC3ZyG
BagDw/VCn6yWF6/icQ2QfEQXAUpre2bbIUxEL6m9ew8UXd7daJcKEtfrcfQn0I2x62IOYSk9EGX8
AQwidgI/o7dj+6ng+nDN3e5/PsMfSDYxvnMMbw1rb6Hfwmo3T6N1CUb+nRTETCEgJ1rqTcYNofdV
rrXdfaN2apzG5aKAQXHSocJcYt1uubVnRMetkezI3mXbZhg4N4w5hdt3QbPBtF5iKR+brYLOAgsY
mNT46XEd6zP/qHgYNm9Xx/fPOFQetiF6v33iCW6acEvHDYaXgj1nr7NrSD+MnLCvkYvc/17In6lh
s29naGJ71CgolxINV7+qHETP4T+Mr1To1lxgaEAMUcx+irsG20guR1h5jnsO4sbsMoNu6wCiW+jX
4Vc0drguiXKYLP9L5beX3XKeavVLJCqMbXsLuiXPKpRTA8eeNK8nq8NJnyNKvVWCXxmQaPJdIJT9
V3WJd99Lsg91cLs/jy9vhvZlSEmDfxtuRogwwPXz/aZAFLAefUj1AzCsQjOc/OWixBiQFaZGYcVp
GlryAWC5ouIz8hrQMQZ44lGfL+xQrw5PbElNpg7cydOdwNaLq1JCt0amsrBO9PuIvqcHB403qGOg
mZk7y9c3SvTTxuWJ7n0XIQcC9ZcrHrU8Dui/pbefCZlS8TNVC3oG7nJ+IPsywAQ55NgvOQvW/Fq2
V/j9xROU+44hhcRiCyibQZi8DKz4Erm1noq4pL7GFzeKbUqoi91eddnSXEhlOV8zJ8UsAXa0jxvp
/X0ikKrgV96M5glXkAPXby6yn5wjgp80biocEvOYS165OUV6XDLHOGpGmbbowl/UXz4B9XLLN9i0
wP8wvljezjXaApK5NW0XakFrSOiTZKuPi6/Y5zP3IyneOxUlCBdjAjPKRYYzyH56+u+TkG7+b9vY
hhcfd3oCczWemMhytQVGjNpMxLOs/5UGDN3TNoqB80hG03gzr+qjB5DMVLC8Spx9HKTC/Tosr3kZ
WZiZOLqe3HH3EGBUiwYxPTI5LDEGGbJmWmvhvhOC3uO0Bwr3UK6YOWDypF9JlPbORrXbp0NsUXGg
P4Irh5at8M/OsLaVtelJRWga4kGYWmIwH65+fryQzi+Ql+KdvBb9Lx8ESKC5skht4pvShmnoiGWs
E6fZzgBCf/P3RhwVyFhBufPSqqK/q8n+WaYRRuMgy9o6a8N4v+8rhgBF4HHGo2iT3up1B/Lfpbdo
+oEbMdZabut2St7MSUWcKGQIn7atNsAMdpWJyNAw+1MniYfif3fpbIAOk6ffwlItCJ8BTgimIDcw
L/ZgeuvMIpcuURwG4kvxufcag/DfT0yc3y+raJqO8eHkTN4uz71A3T76J6mJhGNcopZJ7cfz+5Vx
LBmD9CAYgvb8+2H6PSgKvZmv/ZjQiLiIBTPNSYOu2FCVUuPzGV/rdXVZZys+6mUJoIOODvdht9o+
g5mnERd2/Pxs5HP18GpazbT7xMLeHnx6wITYlGtEUZLpLAt9Ow6YqaN97YsBu+Wz2atV9B0Y2CS2
A7zDGZWw31KbMgUX+dmjTpgojLecQtZGEo1iabXy5Xs1k+nz6LmI583QpUN28TVj0RtO2tF5eidb
PG/Z54skXqZ9sxJI9jqirt/1riAjiV/NvdhevEdk9LzRAoRd0fHbiw+A5F+uqGt//u3r1xV4y7NI
Yk3+GKnsmJHtEuF5gaAMMzRDv58QPp6zTssoHlKA5cMKraCIUdv3pa6yCXbi4ygG5BWJJtzq/kik
SeuzdUQv1+VU1UGx34zNYdVS9ahamoxDvvGFac2T1g1SP0Ti1COAb15qaQmI/UKFKn4VnszCUY4z
4tBLpr6C97cnWyLgk+qkxPgvRdXzUMuJnGuFofN1rGJcDbG6N2IXIQqKHXVBMieYMTkTwhOK1BdF
5qWN4HtOY6hmwY7vauNvW97AsukCy+KnolfOwfmXMbMdSjOsiUImtDZurGN9XTIpq9+KYU0pwG2z
waxHwokkpKbOIUeiod5K7HPXOsLlUyUUyVvf/LVTuPmsCMNizGQ/KtS4j9WTUmG51P9S3QFeYkDb
XR+EQwv7xHShVrBPeQc+bUsYRErd2elqwCMWwwZ8IQFZ5xohFdOFPy1vKjTLn3QO66kLf7Li5krm
9xt03XmFHDgrcoLm43vN6VXX3HlQ+btOz/hzZn1ngkTo2+7Nkcl+Emwd2wlrZ4iueSDktTb4LfVX
Q1rpyitJarHq2Ft+CcIFXXiVPYd3GqvMhx1UKz/EPva67bne+/aaZGUtRO7pKK3u6N4Y6zR3QgTN
TQKLrUgE2EYJ9gsmFlG8YX9k2qzaXACKC5QCPjeMvq3ydzRIuZD395C2rU2XGXDA30fCLV438rtV
J7MM08uhUlT7C3/A6mtA2avHLoruvO0U4/WTXn1GWkRnh4anOalshbeeadcE29VuCrwbeDonKmZX
3zlbQ3lIpl+Ms3RQsjMwdbR78e7E7Sm0TCmLIqGHpxZ2NyYUy6Z/5tg29kfuo/EJVpr0YEmEN7Xw
2GEd8Xyow1WkRQ47BzbiV/4bqRXMKWhnvCks4X+WagSWgtavZpshuztQPe2gZbNV5o9JNlrtL4cP
3RcNHxf7LkoLlkodbfQ2dASe0yGN/WcEOLgVQanJmNvLCRNqrmaLwHln1O5WcFC9vaZwrM9EQERP
dhtPLFFc0tIdLXj0E/aNc6ta8UYtZaZ+tsJ3Nf1K8wuctaAcwtXj1qEHC9LuL5BiqsWtzpUUx+PS
p0hW/NnXXMvP1vKHJ/hxkW9c5PaY5XpzTeRKoY99ZiDq85QvWlFEPiqFD2ktSyNCZC1qM08cMmdI
yNaJyINMmkUItW3gURDIs4SjvgmJvG0vvDQlzLQnZLx0pQ7bW76yheDzShZP6rus0W0IdOAB+kyN
gry20idX9HUM6QK5Rl/31NjHMmuHZjX3BporlnSbSPC89iT+8CBR1YnU4OhN7VPdBdkcGrhD51IF
ilyi+EXQmEmm643FNrAZ8DhroloHxYGaXQslwnzY7SXsP8MgOlUIKqRxUkWxRlSu20dW37SbCP6/
XLerL9qBX1r5RGhsCyuDgbUhz1Qphq3P35Vbq9j6pW/4iAidOr5FOIu0pNDeh1RW+yFUfyL3mdfS
o0Pc4xoRMnRPffKCm9+9NP+wFrovDkhyu6vlWUM50TXaovjsnMlgKOOuhRLUjyfeXL3dae7nxjYK
Pewzb4DT6rExjC57yjcmIp2NL/7+HQL7fzNI+AnHuEastF64zpnmsPNZ8TJ4HepGeWlTu6pPu2OO
j/XvsYxxkSSkZ6qY1F/lvLZihWVuJEOlFjm+4RYk0+zrIYqREpx6OpL2LGtMferK7v38SoHY1DAy
cVX5JxXCI0IS9I5OCgD7iYTszER+WCvqsV63Vr0fq0NlKhJGgSVHxNMbYHEE4vMZ7qVOl/TyCazz
v77tZhuiuW8epm4HlYUzCVViW9BQfYPaVaJFU+VC68qkLG95QTv6k18XimLF1I5gYGZ+I/R7XNNZ
zpmiNsczn9eFYHMcfU3ewg4ZhMKYNLsap5CM9fUHO7Bd4QtvbuPnKw6y0QrNcPTnTpKib8RedWhM
dWe5Qu0bdUcB+tntk9yslNNohpqU3F2XJvnS+hGow6bZq4ZXUe6xdqWZbsqRimvCc2G0U/CbxM2D
cTDa761HbhFdzWG2PIT+SiiaSjfBsBx0djtTO6eaPs7qc/q98SeoWJfDdG5Ys58SgKYsTrkYuTV/
xDiyNlj1ksMkbV+ebO0qz6SO50PighomambxhNGwc8eBuWSBDjk4K0HYPruiS5OuQqmHjyddxdw3
4nfLdEJ9eAstDrxKARZvkSk0Tg9lXZV+7Uj7m+PYFmxKJ8B/XkVrlE1EhYQFSyBurIEmy160CFCw
SPqxkMw528I63gPWWWSNRInZswbQnQffy5vBfQv9G+MEgDVh6TspA/UmVHNN5VMZE8qjCNJn2w/G
/Kkooy5g0LIwzCBA0J1aafvcOpgaY94K2JL5pXxgumLXMiI8Ziwvmg+M7Hq6OfEXkAvsgq8MhGn+
fRgbOcbVxOBqR/i/Ih4cLt+WI2zVq+cP7wSUVNGFY9yYcs7lfavNALKxj21LNjcIPNtfS4ETIyEW
Fx+sIWT13s3iEunkkEpSvjMimBmBA1fN2G2rOBmYQI/USbNHzbqBo+L6xTaXfbQhUqc67tj+/6Cf
1tZyDgEcK36gaWMjEOLlfYPI+y7eDsQM3rs6jQwaTuNQKM3Yl73sFWJpUr93VD6fPD66suH8sixP
02VahmIhiGh7jvj0NARFYc9rVCDNIULjCKQZKP1HnQXoBSu9I43cmtPQphzd+zFmsWBJyi2yGL/Q
2dbl0Jy6XX+PP4v5YyqTN8VJQXKFUzOlLFjC4+4GQrMSEsiQWwEiPAY7zeoTBfHY56Jxd8dMFO97
O1WYpGn39POxoGGokroDHSHV5CSPyYJRtY8P6m2WHN9kG3sAR8ap3033L+dnktev9Bq8LAlQru/e
SJGR9x8JsOu8ifXrhixDGoy5C81q5zzOTjRLkh/6oEKgDG5X6SQsmlD5rGaff0Iy+39YB36KFU0J
OBNnGQ52ChtjyOwDLLDK6jAPN7JBrdQZ2gx4OKZjOCoiTLSyfUxrIh9diGgWU1d30c12L4D5DYlW
NFpE64raSNeA7LtUt8LKiXfr73Z35MKWOb7aPrzZvGArYNocPgQcAu78y2pZGVY4fn84T8BUZpEg
Fz5nPuBgYn30qRPbe6pNb07xnVxVabUbTzat9o1tQFGT1A3/9rrJCnxODtl23JrO3/WHwQBEAZjo
x+kphg97lrYgsV8Ggd/Msd5Xs30SXD6h5PZeVXQRqEQbcEHPSHdXhhVEO17lju+6QEATlihzMDA7
nkP6sKDlFWFvMWBRZK1mjeH6hIsTwSTNJxdRjeUmskNs6rk8A8XyRnEBEUgfmQNkaWZUM02O6Wpv
Lr8W3frkZl7KjifKQLyTcLM3wIyWCOijTEdeRqRmNDv9lhcSrLJ9b1ZrQ5XDPNUTDfN0RydsIIgY
uwaHOc4VBtODbu2xqRr4rSRX+CoyCzjGLiaW3sXcE4fpy9BVuPNtlgg6ud6F9nrQFTOhaqlspmjD
hvwaL7YPiskUfcU1HB+QlOADXhZyOdX4lLw2YqXhoJZOFT1qW1i1OMgT4DyW7SghaeJkQ/NtVxna
77i+UxitdGkrdLFlC1X9BpRxryyWkhML8Pa8mZRKV9hvdoWQgQGHDywYegE3O6qmvrgTikOdm9Wx
9VpodaPP7k8e2kW2hiE8pWMV+sanUnABB9dckSeBnXeA4XBeE+FtUMcPMYbslQFr7mvxHhr29WFg
6cRJTOyD3cntT5pbFVUvf2Hj/6zFpvIp0PtINCSYjoJ46+wzyTCaHq1XbxdbzA1EwnVLcZA41Ty+
+KGRIKcTf3U0KdmU5r16w9e4aq9tA1E0J0FTj5lnR9I2ecR22/vGRh960X3tURpIgdkcYKHrD51n
9hbmqoOWGayDGwfQ+9fxj7FxsPNREPsArP0mUZyvelOwmemHE681xwPbbLj7DjNRR2CONberwAmH
UtApjhL/ISmCFoxDMtHBBAXUKMBIRYYL0me4yzhvkdSzXIB+OlThaffqF1sx5EQ30uwa6WsHqSVi
gBKPaEVe3Lo58DO6Ut9qP/sDaQnSVgio1qsFtMY3SdTfYOuizv+4dn3Uk6Epw21AA+Q01/oE0Dfv
vFxP7380YVpHhLvQwu979wZAI3Jg04VApXDLcqXeXCNru9VgUkWdWsyhRT5boGUtCCgA3p5fKUfZ
ZAz/LTUYxWlL0khlsiEGmdbaXB7vGQUIG2xJxm2sdLGHh/f6cBQwTWfKtldFPO3xpcsRfTLO4TmD
yDKeqG+Jwzmj5P7bqB7qTK5uBQlZv93fWCYo+mdTyhuE/vjHHMeiCibf6tJWpMdV1ZJ3EhpGJ/pG
a2yjJFo/FQWnODZ4kLnhDfoI/CVRWr2v4m3GthKpmi6rgPyt3xlKbeTxlJGHo889hlqf+hskX+V9
GVF/NuO0jEDfh57vjwXwIAwqrnlOXvv5dVV72S3elpDFSeqPqu4y4MoQVfYJVspOppu+ycpuRb04
OMB/bGQ4pvOzDN0obN04TgJ3G8jZ9DIrEZgpnC/TPp9bvROzIlxsA1vKv7VMI9j2TodDRBzxswcN
ofzj+Niav9pClR7e88upge48/AtOC8ECudGvv+AF1HeKkDGoFn2ILHxX6CSdpvdNVPt9WMoyAmyB
7wTgg3Rzq1ukq3n6bktucvuhHg8Y16EBmA3PgCLJLusVRuBa7aq0TiTkc1ST2JH5Z8WN28ltEJyO
ESy6mYcxenzYFmocHiyB5S1RTzpzoJDh/qiGq+YCi0pWYfvR58Jmxdvdm8XuzLhcMEmOIyNphvEH
ICZIfj+MB28EDVMWPLDP2qehXpR093w4L7cI1CtYX8wMDQKsxHrlVSjGtYJsg89dZ85EqvyRjFmU
NBwqvhkWcQ6u160zh76EV/T4il9sNWRz8gAE5xym2RAn3nGLt7abd1VHnsXkkkR479lgOG3bt2xZ
XRpCE6xARNAVKMQtJ9VuL0JhPTw7Iwaoa1K2yDGs0LCoBSmzc9VRzGfQ6q4ggK3ZHGZqOh95hCuX
Eb7tUW5nSbqtYy8ws0fNOYktO1DIeI30qCtOlQCE0FI6uQWW8/f1fjzJDgFOs9C9VgcSGxx9Hayd
RzuQYBj5FmLWw/xo/vlnTTQqZ2femcj59QrpT/R/sww3c10Jnh0Idq4ls5lGQxy/0bbQxSpyfket
ZrRv2DZ496szf5usFqpFcVuz9Y89thYkVu/lTAXDaSjb0kj9MWrqtKroOYTtuSRRde1prhUkt0/E
N8ScFQXNnEoDREePMVfyPUNywr01lP7tWEfVMSgRAjQxePfGP52UnGN3JtfvVyWNMRucvxAoi0aC
HC4r7ZvKT/CSjDAPEu+EcQBDd05HMvcpJARK09XYfHUZz0TbFVlhBAnKijKBYpz0cNw1esBskrVG
ri1+ig3UTnViB63AEBm+2ZQ5oC95ycpuFawI5PYkJXH7mRLWwD/t+llQA9QFqdTP9wQU4jGuinOK
T2iYfSPwlWFYPwBDMPa5Hk1OlTiEv8F4RaZX6fdERa75Jgn5L7nVvujwQSp0vDzPdkmUZwT2jXFe
FWKjV9YAkE7QGMy6j6ZfNu98TlZcjN/GgL+4Ehp6Y3u3cce+ZM2JC67eqKGkx+c0PsBvo1Dq2ZXf
5umr/2KO7HGADygwZ+eP+8R5JYaU/MDsuwVzD/BS96gjzEflSegm+n8b9fMjsDHSG2fn9guiHVGQ
oA8AIEqnYmAgto4E4shwxHVA1ZnyFy+lG2IxyGNPojbD6nwhaA3Q3ZsLH0cECRUNkwGwA1cdsjIo
z2WGp/YOpDNUM2sJ7m705xbYAGhgPrgZeIH0BvM6waw6jLMQU2N5ffDXO+Uk32eXE+y0f7BAJmLU
OhDqvV6ZLMd0CsKgtPGL5t4+fMTp1hb/lEW0oAuFskhJIu3eqLniFvSGps6+/h0QGWxbe55/y9dM
XJucCFnyyTgCCf9H+/KjCd2mUvMu7gEcPbF2hlO5edV0M5XyjkpDecJWfOjmmI1MEw2ZStfNcd6a
3ZvQmM2vwU6R9Qydx7NOFEkWz+IsZteWrkYm44vDOvbWyoYhjuZXAgHDGolLoyj0GcCn5kW2XFPZ
XDkSn6ngpe2oD4zxxWfEEaMMvQaAFE615AZEYKk0gVXwpxaRJd6scaffnKsKnuYjHLl37v22t7kQ
4FoNBG7pJqmFy6vtfzKQ4picIKdk8dtvY9d/VrAI2zTQqTvm1uEryJphr3L79YYIOz0x/2FgUJYh
6FiTpZ8FbhppmTmvVWAV/b9aazWs2lEvonKhYQPhQp+g3kkctKmNfD5+Dj+prXBNKEVtT09sLEfB
kl4bAsAidRf93fDck3+QyBeEsWDOEFq8M+PCdos8ws3h+TE7rcT7JFYT2+OCiNqts5KfGIe0I1LU
VNDWqjt2R1lYCrOtmIjXLAfrRHeBt6ibJOI5jyvhDB32G258Cvufgp+W0wTRtf11rZ9AknQtoL+W
5Zzu6cgGqHdsU+7XZODsYg4EHWF6sC2AlgyIrKYE+IWLU1D77bxRHHfQruKm4AKZS9AqGdWG5U7O
R7R7BV4g103I3th6l34KSQZBcGal5RLqc1gHVuPoeUz5pOrLXb16udgAH4sZdb4HrFRIqUl4r3yY
+MvIWlSbHnU2WpPxu6drivgWvwqu+87AsakcTWwCVQ0uz79hjqUmBR0YZk2ljs+pjxfsL6fFLpYV
L1WTh33nmk+Y2NoO/B5Q5KiVgo8wCKv3wagz9U4lE0TzgXUWAIgauaFY7H4bri2fSaXiVCLo1KvV
H0bbRIfpXOx6d/AWDg/vxEKX94E0Pic+gz4iSxX6STcrCsFwitJ0m9mKZh+FIyppnWDRItJwyOt8
IooweWs07LqPEzFpnAYP5i8ypxFS+d9hVGz+JOoNZzEUybEimdyKK5utYvSBzW/mOHYKrtuetLXg
IPc33mKknwNCFucUCCzsPq+IVXl7V2Il/QBcEFGUwrcyWM5qkFqwLz0CpUXdaV5AKUbMlTwWwbQO
kZ3mpK49FKLE2N0z4+YdrVQaKsRKY15K+V9UwEZe0QSwSPf0QnT7WMlVc7l4xdoVu96tAqb7vmIw
cgwkgCyEYU9DcgGcH8MGW/QydaSukJ0DqXJkvySxlDDgH1YMgz4z5LrA1SuDnR6Lm9GSzLcOzB+q
yJqpFxb3teCMEOWjeditco2lW0G8AFplApJuHR+9hSFswkt8XHM8AXTf5rZDI9te7W5NwR2boy8e
0XBKjeqKuyr/wDfX+Z+mDnJHvzi4DujRKIJpjU14SiMZk1IKvpwoeYyFTJk53rB+V6Vc6NV3LA8r
n4JPkwB+JVtdhM6g8cOrMCfSAURgLbQC41BwmYzk2v1DWnCeP+E5K9XMBrTUmw0w3REA4Dfq68G8
fT9az2fK/za6cyrJyKc59pIrNIokb6aTY+9JrAvArEjehkT3dO4QGdRaSXSEEZfwE+zIu2P5+ja/
C5LNwkBGuXsGNzYp86JvkT2GBw+caa7kZr50u5Is58OimB7dE1Cr9mh9UUzxyahqUlzIdE9mdC0o
5VjJKPZsQUtKftqSPwwpb56lHFg83TFDEGRcttsIfrN+2gmQYF8aub1EO2VaQlN3MNwR/VJfusjp
VKnmWoT0YKf71WwAoRUv8WJ8JOdweUf8TUfbHAuTHVD+iTfhJFIKj7UaG1XFUi+v81HdZA3Kxh6w
VCX8slT9UmKAYqBi+tvBjpPZ/VXcGV833JM/KdTlsQzsA8sY0Smk+XpHSncENbxEYn3JVjUVwTdO
RVJcd+AR0yhddtH4fSdTlzML3YOsSWT1W2Lsa7jkpQaAy2Z4NpN+hHFr/FkFlpLdJVpo7evIwMhl
OfqDcviL3QK2ioGZ95H5NSL6yPQjStQA93wYEpV8QYKuFTB13EWLPWK3kGBije8zEIADtYZi05qP
XmdEGmRr/U4q9sT2f49kjEtGXhNfMlPmG1xGr4doSKzzTYol3xKtD5Wm4Kqc+UMHu3TSZFEKXNg+
6oN4tzmhMdJvLlJjXMHZQN+3bVGA1Zk4LaPaDSybDLyZEZnbnUjqWl5XJcM9a9cX4Oi2U6PXYCMM
8uOOJJ6ENkEjYB4fuFvW8GK97OHffdIPza2hV47QVru4QpziT6YLICTCmoJXg0iPmwJVHw8JkTKX
Eb7vLNvo17XoowWPR4cqr4rhHhAL0GnYqFNw0JhSxpgGJQq8nSjXtr6IfQDg52oXolVNHHyqOnNC
wWiuyPIU96ImBPKbvPvUONOSjfzHi/q+DD17MHxY9acoWg9DLMs9nLZmYpjw0OhStcNqyRp6p1ux
GzCf+yZmbg1z73kUQwtPkt+Sk6J9pmiDCF3JTMJMyRV4gIOOyvSvKTg7g7QUwZMpC9bVt2/tijxB
EUpQfUCIq4FlByy+7Z7b/fsu+9SYSQwnJo4ml50P7iZ2+NSsF/PCue9M7KGyXh5IZ5nFHmuVH3/m
AnFG0HSV/FbGPrj8TWmEdAuuQiBq6ICuCXStK+VfD+ENt8Rcn7JtMaB1iPK/N54+q2m1HyMdSqv9
VYVblLcGpuG212B+C/oFMmn3Bn4v3VMJfwsoXVHLy4HekoS1jzKmc3x+Vx/EMbrbz5OtnQQHTOTb
uHwNqpMdTE+dAmmMIsw0PbviBhUI1RHoomm2PeTjFUHvbo6BTt007L28i7Ejyu6tDM39sDC5Rb0D
yuxytesibK+En+cmxoafFq0ozi6CwhRvQ0R1j/FYUBwlF/cIAi/GuyN03lvMIelsvvPFr2+aI2w+
goXZLzZ9ySNyCAk9y+Sa7KDgoawb1SMlqRh5/SK20Z5qvO85l7pnQpTpx6L+1YgXwgYe8Q9W+vcj
mu9/7L/OqH7LIDzbGBq83Do97Yc/Y41TrzcIVt7Wwd6rW7KIJH91PNqgM6346E6ltlgbNfXe0ggm
R/ESFfseI4BJWHisbSLic+efqkg5FdrwQSbQfHwGWVVwTVkkVVOQESkJ0E2xpIl4aMoAHgCKA6u9
g3YuCvXSpMs9dFMZ9zr1fynh23364vQWuEehguaBWRTu/WrLcdEqWtf27j8EBG++cM5YMQQSvgVS
MVj1Bv/NvtA4IP1/XY+xx0lOpluVDyhkwsabZ8Fw13XG7qwzfnQPZiVHY92dJIB8Zc7XdeTp0Vzz
hcF1h2Z7PzSaW+lhoSmJtJeP2MAyv+xzbKCaK//5JMHesJG4PpuGKFMnP4RmlDu2YHmPZ4uLrm8t
hqhidvCE6dOGR/pnl1uX/Eg/Ij7ciOnZXwuFCymkEA3p3UC4Am6h+PBYnVDuUln/9IpvCC2iWjHs
3836MWYO1i/VhfXXZiiTwWUxcXUvSRKr3okL2IJkHrBTsnuZ8GdZuhXEb3JXxJobw7Y5lsxke8mB
AH5l6Osde/qC9AC3W7le29ZQsJtP0qafpl8i+zGVHo2+6N99FZxxQ9u5fd7/St2Ma/gwftr7J+0F
AfTXVMVSFnw2RVQ4fN3ghEnIzC5APJn3+dL6fxBMnNfhP25z48sj0CsOldebi7XOk1jEXO42HueO
8GHQ1dSXUF+9IqkKZ1tLUVDslRwyLwTo7Q5XR20hgmEVUZuBxuomrBf3TzYt8ATDBwgQ/LO8l/wY
PwhYU592KYCNnyco5dOB/pXWXCt+wx891XGTAMxSAQegPa5+bx2L5yT9EXK9UqRjC6ZjeC37SGc/
ic42nx56D5kx/41OKSxNpmLWRBB/aJXOkE6cRHpnf3lI2WpupR36QlbxT1G2vdfr+nd5ythBjYsc
YKRhGTccbNyS1CafVZG51GqMbTRjtW1Xb90Kva4HjFK/51+nlGM7Cxuw0AQ70tAm9iuXMj5TS7cL
RkLAYyDRUv9f/q9W+qP1pE7jw92WomMzHB91UZcAd6mbSbJ+NJXL/EZ5SRuiBSeVNApFN347CcaV
vFajPdCJUWHxqs3sOXMT5rYqtCwgjZgRiNJ9xTSbXLedCOgFJW9tsTLKQNj493LCnzgAqysqRmhY
MH9SrtcMpZu4SCfWgWalE2giaVSJnIZ7rm/Sdtu/HF9NVOmbGX9M0CqGUPtmvUZpnXtGvx11ES97
qMS6aMDT/wdx7WtzlAaVIHNQeHhJtF6t0ehLWimn8n03n+yaT3nEtF0sh4qxA+a1ywznMNDcAHZ/
h5Gv6vK/2zmqrijLXGolhV8DU8P5pDXtlTZSBWlTBFIBKfUBrUYvlCYVEZxq0wHwMfALy3tyKr3Z
/4E95lhYYFkYNBJxmxlah552PIxp0A/1mlYLt/A8d2vdJb/JfrXI1eJx3raLqpTwmCQ5GmtoRt8i
Ju4QvbBlvRfYWHPcocKY6ff6Rwg48SuZJAFRtsrKP7BmrQ5QGxsn3Z9UPmScZQxPou+2wDn1cFP5
70pdaxpMUKn7cZHzM6wvLOSBdIkW0YIZiXB981BX1l4xQzwoY886LLZo/HOj0EjwLO0DfG9XlL1Q
TbxloyqItsR4aaX+L8tfOcJPdorRuu8tm5cQcFQXuABgSkrQckb6ciSdkqrMPOM+9ORKvOGTzf1B
STTedo923c9vLwmD7696nqX6CQ3hryArB2Hy0cBkcEup43+jgAzsjE4OGryox/U6xd8BMd9rQQ56
bC+Yk5z7mE94gyIxhH4gEanPJoiUeM5/KONWLK951HtwRhYESEFIz1zcOCT/+DWGbqQEti4QggDA
6dIlD2YvTpyuTWSw/1RgP9ED0280qJjb0Yfwi9KB7Af9AXDTwqBDJ48aba25rdAWTF3qTNZD/BEK
Vu5jEJ4kQC3fyWeJM7Q6lJPl2tve7Bi2xR04OMtyldBIcqjw7923yadg3agOFJpPy992tMBYKgsz
D5fk3aoLF0UNdpSrLX6nvVnkI/HXKzBKA8RHIAKJIDoke2o0IKuRAZ8NIimhmLH6pvsgXQrA1rdT
Doq02gT50N36bcDiSVDrTP48A/su/FyyjhUHprqweBE3VsT049Dqh4qHy7PIdTB/m29BvsekDLqq
MheHr5BqY2suaqBIAAg91GQdVqYpaNkISqtd95ou/exaOk/RnBq9QWLKF2NBnKiid1tx5GSu9YCa
EiyZAi8xBElVIB7HhP07x8RavPbEXngE7ScYngq7vcYYCrSGYagAR+1MkYcN2rDOT+H8wgnq3JCI
6Q9CDZyjr72oHr5JNakTQ/4oJ6rKNVvLTNOk9e+6++sLVAaYUr1lZC2Rwu8W9amZwjc78Ssogb5Z
RDH4VaVsEs98g+Qs2uy52eD4KSd2SyS0uCQ42hEtMYJCNsZBrxMuUHNOuXbtOwj5kAgSc0X/6mVt
DaVnBfwyEzDYoV2wYRgJiaIdH30PBjz2vRjHMnVxk0XJ9NdxQkuvfEuDBBPxFtFpenWO4Dje5dw9
R9EUcNBiTp/HWBCbFzbawwleB1XNqgQbdacaMnSGFEJcHF55nIYjw3hPxsD8Bf/2wICvdOVU6qpD
DVJFr0OjO27fENAkFAi35Xaglp6Sjj5UgoE/R3jdFNjtV68NmPysvtmd+QvvBmcSuwb2BtZttC8c
Ev8mreRHhw0pZsX1kKkkmcqg6SfxfLQrnIGRF/5ODfJ5xG+RCZLpNqLSdQo3r3Slp5x0QyPw1SHX
Ycxqi2LlAcEYu72/4p2vWhCNNoMTgwr7q91CMFdUDjGiT/53J/WCdY+FSsXcA9Sw8KYc/luzTzy6
Zrzv+LY/FcfNwUNOO/M/G5IqUrN8dqFQkbuzmv60dQS+V98LpnwQbDk+YOJY6BttpiJDjjKa8sR/
coZotGGBVyenfGfTB2ZwZz5bt45l4/6b1hmgIXOdJ1RQ2VDOoOlV7Ww5f07Oe9JKltcBnX6VsqOQ
/Dlld31rTO1fZTvb2Z25C3nBkR+/HpBVYs37Nqk5WFkBSt53PN18slZfEsk8D8bZa+CexOuGgihQ
mWERwqWR7eqFnpnurrbu00qXCFBi21fKpXJNJn1AyGhU0eFazc9WN8Gv52uLqo1PB9mEM0QzuN3s
W0kn/5beJLUe2uVW52rd66ocI99gL0S1Ia9pQAIyHAO66dbAXKliN1kAJynpN8uatr0UyGLf8sLP
72dFloBGk3bZ4QytrJgYHEsijqJ/GsHK3I1UpkciW4sinKdhsIQQxxiNufC0l2Tfnrv2nZxyr/Rl
jaeKM18Fi3BhHF5gYJ/mMKspz6yXnM0f52mCCB2Upb20vSgsgCAubF5qjL8c61fe8GsrUTmcPH7D
dM/sUzDtFWmqyWxpEo6JiPz7M24icX6MmCCBWpafBAHr+W8fEWKoypdX8UJNXCSnexCTZEBWFzlm
BxV+JJ6A1+DCXhvvUj9qBnmUireq6A3M+jPfByrUTtitkXy10Q6js57klcaPsg+CJbsbDVMvvvzt
5LIqla1e5Veea11zWxlrZzrobvWyJ+yxOaNXfVrwPXKV46lIphY+s+s9r9ddBxUpW/cy1cqYh7cA
K8zZeVq27AjHD6ayo+WXUtHx9SgEZXQclQ1cqjXzECLD2iboQc/xa2sJQuR4xyV+I7+l8LLmJdLR
r+YytBp/EBHAzB7jeeg31l+c+BUbZdHnBzy/bynRvfBM8p+W0QUUCRc4HnKKAWebJus95sE2tx3j
NESFsvU8xa/4jZEizoZF9Dnp/lD92MxCVfmPTr6GoB3HBJ/Jtps915WlgnGzl/s0tYIpw3u64939
4B5SXEwBzKXLutdXmrkY3hs6vkzKrekeAgm0x1hehi8rTfJexlVNarp6Sg73AmrEQJJegWnjjtn6
jlqvOkoMAVz5jE+ssU6LOjtCmmnlZOByYdrx4P1TYWRmiXk4XpzrNNmemjD2L6zvRf72W1GoQy9G
RRCnwZtWLrZIKpHC1SYkSLD8YWBA/V56w8/bqnYJu1EJITBWHypSCXCa62NQnZ2VVw3dHaiR+B8E
JHMYovo6NAupkiGhRvtpK1WifcMyPeNBsYm9amWcasm7OPwbhMVd9mzhzsVylQc5u2OXVnO9VQs4
8D5JfYCEFKVk82Mifzx9Ivtm6ko6PVk9DDwKbpJzimi5Yj7auWqgwM85gu0oX1CR9vAuvkfLBkhb
1oUIOpH3uPdZys4eXLfDLAmi7H6Cue3AsLnjzKUvA7oUEoHQg9oKhAa4FjUAYlQyT3Zt5CILNS6R
4efu3TfNXd1+6Bx8erkv2t9iMAvjLjhBGbtVAXJ/KQx4/UKpIo7+ZovXn5WArnO3cYDhD2s1Lapv
M4mGiH3H8k1+Lu/0uUYsNQpt+XvTAY+gnP+35qtJNkR/kuueJbhGxidO7PwZlU+Sze83opGE60OE
2tzTCU/iFMwXK9dgogYBj7NA68we5iToADaavaxlvaERMcIOi85oYhQZCpKuXlXgSUxokn63WMoc
1N1faQjVU8G/6lVys4EKO2XW5BWJ0zVRnA5nzsN+uvovKZGH/gij1IKKsLo8/f8PilJSKl+i8UVF
8a9K5r5dA45dSO4HWxQftfQ9aVUgjv5I4jQ439KRVd6Si81rWwiMDo80MvUr9o85R+YyqiPHMGsD
vv/xQb+c1iMkOVp3HiZ9c6HQNkD09dfzceKVzasmT2IgxCdX7pUlxIfCUFoQS+qob/2VKg5p1/tc
zwNOv26pS4B2u8CsSllpwEOx+NWXzVqIVQTlPZZSgackVrS+kmohKfOYzvT//nMQm3+pgwpg0RtB
pdEyMny0hLNXKM3JOcZKhdZrtGLC4ClfjmhRmPyu+lMQOXzKAUIH7h/Po5THtywjsk/TtmyovXGY
r9dbLY2WVCFXzoLMgmNO7vMu+hRFo4kdnYN4S1PnEUk4Fx4Ygxj/iVzx9bGuRMJActhUowqG9yZR
8pw4UgksvUa/O7IqTIGVGgNoP3eqKPmOGu4XJ02QTIwPsmgHsy3z3HN7dV5TH/8ibtKDZ22RMUU4
XWrLun4DeLFgbjSP2b/1wnvvI/ANRky+NZMiKLvaV9RLxMi36BSNoDB+kH/Zmyd+Pa4WhUTMq18l
qa9re2a0lSX3TzGO3Gre1v25VOyJAEwdu+CP4YXyY8jbHI0RDnLd5AJBxLJtx0UBQuNVfdsrLvom
ME/sWtFsuOV0cHCC+ZayFrsjBTcT7+4wZPfx/LSbjAY+O7BVRq+n2Rz9XkWFEkCa4ykP+ZFWOz4y
qF7FYpE0QS4Hb3otb5n1iofhzZPD1N4ArsHbNxVbkTDPoa7sVA3oCwqoyO/2f0lUN8VTeL1ejeYo
lYJbNPMWU5kb9O7AHqYabPIv9Ck9/cZ/y+5MvyLxc0c3JQNXNbgvMP7HsjNOm+Q4Bl2yTZKUBnL1
OZoKj5ni++JVLGeM1sRwWHunXe4q5czpiQcWWXEVpvI9f3Nve/i4siUZ1gqPe4ffpxlzy2CM3AHt
UP77CuwFGpdK95nMaaNTodV05c3Xs9PLUd140mxiuFiDekXbOWBxXOAPtjxT2Xkz1W+cLXgQYjBh
Qu/1rUn1AldgVRI4ULGNClBWgMpfAEkgC1V05jLQeciq5hGYanV2uV6vdlCUU7+TB1b1bNyUSKLj
j7Q0YFAXv431ibMDQZjrPyTdGAkcwHMpXzsRAh7QdBjZdtmcco6lcUY5hYV8XvIxv2ZcDO69D5eU
3loNYtzlc8CNk2/4yB/0j23++ueJT4Oib2ZLXwttqfloyxaFrfZr16EzvAuVJBrr51ejEeKLeXcn
/ml9BjHleuzcG71wc7sc64OqvEHoowO9THpY9mjdcz/bL/F0cygMKqxkUNnM6zn+elwsh66TpftB
Ks8aDCDw90V7n7sLSv9IhKpYx+KwGXIg4/S7pZncKq1LaMGEOBwlHmDxxB7jXivwgdA3L0O2xkUJ
ZkXonBY9E8FKLCrFJVpVmk2EhIh9k39EhbweQFjpNcqewTau63ZudupA6cVWXNQ1og5s22097USm
p2QSR3GfDgItDvQYbW895KjzdEjaRUapn5LlFvGUjeEyZ+JPXrLvi9vwBsHe7d7OrjL3G/20JhWc
b6PWFuNf1fI2TW4quvkzQsWCzJ7v1iWy922J317cYo26NiFQFHLty0AIWEY2FupZ5UR4TREPAjjg
iHFeEzfzvblaEHNVYZr0bPMvCbfYiXGk8M3BtSJg0Es/5xhcsVutiucA/HSXnFGEWjf/CtQLr5eX
u8XS4lJVNNKU9/YwqC4MmzlM2qA8bCeDN4orRWH9GjYcYt//VIXXSwyt6eSP3lErKdCqrz1nXjyW
LSFVDVNh89ryW5HPEfst1pj/bGZ5MyB0UV7TC8GDNLX71XZs0njuQD+/xdC5VtDuxzGMYnTceqYA
kaSA9Y88lGIbtz3E5utgcHAkSaMg2h/cpbiW5KbL+tjkZXJFWM0F4S3S0qTr2V+AgbaPR0v2aMsQ
zU/AlMeCA/YMDcjAeaenyk4wgaTVnLPvZUpvPfqx1/0ABe8Ojlin2dr5XDRlnELqztnHZiZ4O0x9
pm/wu7yS+ImQJ7Hlk7JNZqjVFxO+R5wZHPyRyGm1DLXakfg/1zFJjOYjiaTxB0Ab8csvr4CjU/RR
rbJEGLiB1J3tfneZhZQCecCz35vGitPf4KTABST6E8JWRNPKsAG88rz6Pfxdt7tXEknVJGETWGz/
b7bR+PkiRP2dYUkQiuQf8qmeU9ucsrQ/DSwzNzsXoioP7AQD+18r1z5HboCde2vXLmORhcCb+MX9
zcm6oGO2NH6absq7x3SshsCVjrRU9wgRlY+ZNAMAubs9RDKTgvJzsRtWBhlCjzIk97pqNJPb5Sal
Kxsaio6pOEzj6JtzeDd8cUwOZoPSn6R2cTe2rP8R3XDtofIux76oz/XD4/DWQX5yC7LPZlZ3j6AV
DeQJw+fJK4lrmpJ/iD7aAyqZU2FkjLZ3+x2jhZi63fG0fzcx/tqcycQuaaRDTFtnAjTNTQnOA+G5
fF7MKCAx4QkeOIB6TfNaRdRB65IS+Kztl72GrlX9xmqmV7UTOZirk8dTmcDRO232NVTjDpyU+yVG
eyRy3M3BT4/4VN8QJi43HMkUMfDAqHLiPp+vKbLQpFI3P/oksQsq4HtFSya0YDYOIRPaue+7v+re
40ctCnWjd5EkIJjvQ15ucUnENEbb5sMsFqmqaXMKAYDR2J4nKbtHhO1nI2dMm+VcpHfLBcHu0mNK
hmKW9rnAAGwjyk6csJBq5Z4EKKzROpa3WG2JBc+JwNO0igQXbCfUxykcV5Vo88ZNqArdJ3iQbpUp
klEYD/9hr7GHHX8IGPsa6hrgKMr11/Vbx3lHnuxxEgYnDhRSqGJzb2Q/GGAPyNoNVcMIT46zuxeG
vnDlz0YcwuHIkSyh5mHUy4i32cUQsNPoc70hIDO87LSqLHqfbNFbJjRrqCUqSBlvyymWpL1cqeq+
4xWfBlHQ4hSShUVz802Pe5YKy3IEz7BvVuz5+ynYZhfHEY3w5lpQbbyKAOqM2DXyPbD8iZ5tsGZE
g+kAfPsoHClSTOoOi5BbBAmhYcuk1JL9bQ3SKcdrHXdldVq+eH4oemGOs3oA8p+xOC/3JrSHrDoZ
a0Dt6gL4b1+IzPzZ7PjuhpbZ2auEZvwzwKtQkxGYvcu3IxMY/+NfnaJgtYNthaTK+ZdehFFHJVAc
Sepmj8zUEmZZieQRlqyd42gu45mqTlR9DODthQbwhxjQcm5IjJGFA/sjg3OpujmeDt5AHjUAbH91
rKph39FXygyVW6FYk3TmdY9SGxd5HyoJvpbq7WXk2qwct8AUA+ifw505ELSTAq5CnBY/f1u0T66k
9uLiE1lLptPNpl/Tm9UtBxOtpKEEwmoA8wYVeAV5/S+R6V9shEtNIR5+dYDC22K1LY//zm+T9yPO
+1yzOJNj5RH8O/RiH4kXzziGkz/tfpzvYG7WJ0GzzGmUYePCJqfzRpfNsmyba3MD3s+EL9YDcXWX
QZaVo+PAVt/COoC4XwdEqXzJxJyi50jDb4HCbnGI+QPIL8pg9AZfkWaFFHZNKkYAFEASdjGDnugz
lo4EMV6X1dROFB15D8N1Jb8JEJUi/uDpaTFp6Q1ASx9tcQeCZRHaUbJG1xWvFUlPk8Y4Ye0m7hin
9Q6k9+rQWxG/sHoQCkF1OkW0oZv7qAbVUWkMuaOz5mgLuWyHBA0KLrjbPMu6C9W8UuDZKdVMAMSR
HTEJuEvXcYef4ZtYicU5HrM/68lh5RiAs2Qfp40L/tAf2f2tYZuF25bseaOf+Etc+xZLRVV1ZtnD
Ah+ajAxaxFcdDPqDi8BczX67IHCqp8RAuL72dZdmILbEK9b43EKtgfRFRu/to3P498zyjuFAUpRP
ZLrEDGf48pchD4xVyknbiKBLOBtrgw5pLqoR2AREcWFKM9gdgKYyBcbovgeOfU+9v1ZcD8He0Bn0
BDwkSACD83PYkNqSpurf3U+hktqgIno/FsZWvWo4qIh8T/KRD1lG7eF9GVbshg/vNzVWLeYehM4+
7nms+U5mixHlbETTs7nOl/zaZyOKzdKXclrWh+u1eIawkm9K+ELLNVvdp3oTJaYLIpkvdw9RuWqb
M8ELuK0wvGvrkahnKxR/0uFz+BrjJjT0ah5ai1TMqngz+yReHJJp91uekldKZMS49eObt9vJGMt3
kciJhlA5ILWQ0FX05neBuDVNebKefGjBS+p65oQvSuw2J/ArfgnR/UOuqmi72SxpFNJAhYDo/lmE
sEfFgbv1gA3q2wZ3NhYsQGRYCST7qd7uKDjlRI2N/20CSvyLWiByUHYo/PpfyamVpUehvSFU9Yit
HBm95WlSh/UjUInVnqOonyL7IMHDL+ZqtoOiDDE2U07jhA+otFy6jDOPHxQeTxE+4rabuIZsPaG9
Gzxh+KE6G02EQDsc+kkDqc6E/rcak+0cWyRMMUClXDqsFy4/Vk3sI8h9sue27xhpIfLlDLDhETjV
r5Fn96PWW3kAbLS5kxtJ6s7r6JRXOTJrSu2A7jBxMpQhZuOP9LHMMYYzCkeyNMfSie+YLxX5SO0s
TG80CS882KZpsSFxOLj3aPvVkqvjFfNf4Yzu3v/i6VqBB3lXvkIyHdEljqRNCqk/5jS6kWMwnnyf
KPbcgUCMPre3Y18y6kDi5oJ4sdsEWTWoWfX7+XONIljihkYLV9nNc2hu1SEYCakcunBHY5kfDa/1
IBp1De6faiLkPj0xZelbG8PkoKi6IqkF2O0gfoxF+hHllWpPL0JM+XoJs9Wp+sPMJZb8nwvAFrAo
xCzYlQmUmwrD7f6nnpGLI3U6oE9zZ3UMZHnQJamncfvkQ3jhm9ZA/6yMcIVd4MpS4G1glO81dkPR
i9ovyTobpEZdUd9Y8ErmF7NPY/FdLC/FdCNzQSzjC5DH/vu6VT1wUF3w9a+sOKojjWO5KjRSW4lg
cgkrZnyxYqGxzlsrbE40aykhIkm7/SjSYuwl3PheawkjJ0LhSF2IOuZNvrPI4OhJnf1ASoNryaod
pdf4MpdUCOp3r/PkGUkrvp8h5efZp/BcJUB32wGTW67+6EntVa3YQ9YEbP/w4/fiBBvrcWaVhzpi
GHEEUk5jMpL4FSsBM7xvcdWFbowe45hJPMTFZmi+nlXpYzWj4L9t7mUcpavmXKkGvXZfFr5FxuNb
H8iudML7hIdNX9UGWcxtdafakOhKgUYCLCvESQu06ExX9oDKp14+Mg2eooC9CMX1kUq3ogG4uQgJ
NL/PgzabpYk0I3oFOblJRQ+4Ufjgg6vzYe6FYVh6uffbKgC+JAB4Vj9NIFFPlQW2ATW/c55MaA12
dsSIAf0rqLIwF1Ch7dBt/kK1BTrJwyHkaLJYBrL1Ro+kXmfoSqmxIDjHH1NbPzmbYtpFNFofIZVk
UVl42o4NsnFxPlDU2GzT3e7qKS7reg/r8lRTZsxdikQ0qJUBJxGe01ENLnlK5F5cq50MMp5/HVmR
FNDq9xoxVTr4azbLzEk+xsSEi4Axv6gH1gs75MQogVTfhJ/JP+eLrQ7SveZuh5Az6qhXiHCnC5xh
Uue76bkdWL1ioPGP378cEY+ZQTLRqWhAO0U5f4lp4Es4GhsP6VHQeAvlPrChM0tWJQDBcrxQlRS8
zA+KLW3t3FKp6vs2L7gTu63wPWBs6dqcadSXW4PaC+8lgrlSKzLBnQUnnZU6irFnF6it3jhaiNRN
p7miHzqC0E0aquKmIM0UXLfxsYCZVIvFkuPHdI8tBQpXBbNoXKzfV2FbjAbZcJgFRFIyNB3nClMF
x9FqTnv91RbGJ6m/eOAq/Pl0nCAasGH2e4P+9wz3e/u20CimgNms/opyHTBy3Bp29cqHmhlNGDHl
hYVroTSIzFj41FHYsV5Kxn2MZaBll0/39mS5nIcHiD7rNCILaILlJRnMVMs/2uA9MPEsb6hSxvGb
Vkl4L3H6AXzNxw1rNZyGbpb/wZRHqjAdf5of0GE8MZ6eJAwkBUzq2JzzqfQUFQIrwSnolA5Sy4/y
M0OI+ok7nT1sgJ/mYykVw4KkS8WYU2bkpV0C5KU8T3hyfIuNyZa0h7w7bGZoyTXWACTDp+JpJ3/B
Y/dxTg/FNgWnrRFE6C5fGt2lnShNaCG329pAaUFzs/QJ2+6FTPgWMxpv/fin+vDpOkZlXRfeoGYR
2kpFF7sELAQVi6ZYfwtnojhWOIjVPhloeh7VdOUe3j6ORVDSun/soySYimw3s2Ee5COBSTokmCnB
nbXyztgGQCcT5FMw+osbh98rOqX4YGrsGSR0N0p9TEGYE8KvQyW29ov57viAbrK+kCEb+ZhYfPJ+
ahaHfOzjA3pO4aO8nLpdn0/lBydl1cfpTfPb3TxIo+0si8/ZzzmbnZZBq3p/WFbTF71M8F/jrHuS
UgctPN55PNqdCzS9mAwhRl6a3mzcrzjcqXDHgiFBzVxhRLvMeCorrIunbIITfGdUUwt2EVOaj25L
0pA/qlzMHacrov22i+X5/xiD4Y9Gj/rGDrf65/oY4JIUsGPmxSvTTrNVNSr7+1IBnv56KpWZoJwl
oChnnGFUYaKl9eI1WbRGmB4HE5XrPZ8xxg/oCkLdPQyAQ0O+7hwUXA9AL/XyyANrjKx2S1YSo4MU
fGEmdFCyCOTRDeoTxTl57H7imk0Ua2t49rPC/hgwTXXYYVE5UH2iwP8pwMe3/cUNG8ELRMkhpgB7
rPNgi4ZVX1JdKYjrKOv0RnHHYAPdFcd1GJhBH3Kxtstid+KakNTO4m+ZyOsDupvXFucrIKfUeR0O
EXZDUvwdxXawzzYl75UuP5I4fusIwlqc770WgCKyVEFqtWy+7r396QNbR+HYPqhCmuEie47/BQxS
ghKA1kq3OyxhmGjgL6Gr0/e4yOZOpzwVYocuwLnejw5LUlWXji12ZbxVYOi532Ilp6REWrLvI14o
2omJWn7/ugGXeTrtgeBOonol80u+UpqTAEHsaAXT1m+XSV6NeefN9odLz62mDqUpkHB+X6GZ96/Y
sYgJLN6hw3MCU18VXgL6NI5rLiXW45V/2GWHN9G1Gtzg7Hfi7ou0uO2NqJZ7W88cS0Ef8EYtmtcE
2DtwKK9lH/JcLNHhw5KIwe17rlt3J489lmlJO/6Db6mZfyWFg9fOLsf/VKB90DQbK3G6VXjLbfvT
prRV41kjRQdgQnY+Nj8uZDJgepMnydhppAOHXvXpDLYWbt6K547vxrB7dwQS39joA7RJiId1U6lY
fxomVbfKroyFG/7Ji6qVrJXJ1FwsLKdSieOPmHSqNGk0hUfC98qthw+7N8D9T8P3su7yFEwmF4Ow
P6lQWJ/pJnDXrDVDmwYNcDNXPTRVf8691GEeI8jLlWPG/tvSvf2EHj3uKzNfVTGARcU/bsRsFagF
Q/d6L9gm2/9lZ81g4vHia7uDdvqagOmuaMV6N6ALRuks91+odzkLcc2sfwLw32XBGiz0WG7KxpZb
v2BtTO1AkjAC9d71dv7B73oQhGErE52v9vaEC6jKm9mpRXRDLuCp+y6b9lc1TLN/2DSNQo8oJdX4
fXcxv6atVJU+PS/EWCL4pO2g13N1NEf0QlNFc/9fL6CdN5c19yQ93vLSJ/IyFiXXprDc3cSjDYAc
ThN58g7Fm+rAJPjZYbFDNuJPe3N/Wvs0l12HB8U0AVkjsjSs6+C4q2SPtPPtFv2GBlMmq770JUFA
XM8osjWK68cjtd+kW+AYc2nTJUwvo93TNfdoFu6YvO+NCFsGLaZyl/nzUJRrN9X4aJyO5jdZ+Ug7
E63SLMdtvAo41t6aUxIIlcFTLMxYOjyhYBIHFhbSb8hAghEL8ZBgHFrA/RdoX042EXU7d7wEF/8W
7pmgO1QMK6LgF7nUCSIxauzA4JdNndsPKSElz9mJihLBsjiL97o2mixu0OeylSH9qEte645fsKt5
jTzystS6+5QvA9jLlsb0y2L5yjr3zo+X2A1aSAyXYayYsez3X7AMX4SelS1T/0NvaQC82i0z5dO3
GucEvd6pCC5vapefgPwy67+Vvw/E9D1+HElD8KzxU1blNL1gF0Yb5ygn4wuxwgasVO9E93C3sj56
ZZS70fWBk0w5FgkayBBackBRONPYfrHAC+JcJGt3mAmTMAzy8gM7FV4cMqWXpERZb1FuyERxmegf
U+O8ex35q13TQYBHiVUdmOTzLlmQXL+1vBRP5jIAsgFlVuRLH3eU7atIYgjT64Ld0leFEpw+118L
vkNtajYafhFEHCCiQ8BTh0ZH4/MnM3ff9dC/dOJofp57wt6W2xx09nZqnRUMEiZxvHJFeMVl8B2C
X3oXh00KR+siNS2eywHmqZL+wO6PTwy9YXytL0s5MBgakGCJLckO3Jz0bPerqhybWwJ+Bp37jXQQ
fzZliZCBq7sIhDbzQlft7b1dGSUIAOOW5KXDjUO2akilUI5VjnxNS8QmYtJ8W6jdwFsRoJRRL8hq
wD0jI4PGBW57n0fYU33TvbWojdKt8QpdPECCFODRc0RHIW3QLc8uUo2v2PTPjb8mWNttMPvMnzr2
rmXoYeJ1a9TASeUT6b/aqIhpWqhfUuUGpHyPHMTTc8/HHJZDA0ZjmjaFcJe4DjZIEB75zy7QcK3U
jM7+4+k2FgXgH49ICtNYQQRJNbukpKS9SY0v8xGYLpkATW6l+IwzOQnH97ZgOpCAmLmvnjYDs8Fw
UR/GTmU5r016ATT4XYmab5mtzDx/SnSixCzIIKmG35rgkvE5e3IDMceT/xvvaF1/WbdmNlXhmGmd
4z7dGn71zGqefOTsq8f8i8oBX61vP9leMI8dlOFOusII8dG7GsmU+mz47HQQv5W0oAm7UmYVbLTZ
FN/9Yqi9czWwAG4Ikl4ROzsETcd1ouE6ZLUTB1VDc1qPtqftC1hGxIWr1nhNmVPqBBJ3U7GaYL/c
PDh8T2dMA9RWe+9oGPhHtYpr/ne4NTc9gLU+4Q+mTc4oMezT/fSHL9mQ0NPL3kihfgnZP9o0aAx/
4H971hXG1fhyEbZunVsAyat5kn+SDIrSFrZqVhHyTo2jSs9OrhazmrfoqIgHqa8tiHjKNMNsURLi
PNRtBUfil5KJlgexEHj2XbxS7HTSWViL/LNtQGSo6uK1LvOi8Xe5bHR8KyGmMRarMNIDDqq6RMKC
7eKh3xzSERPWvM9CTQ8HkWPlUAs5khxi+mjJvaTG+BVX7GGTKRNyZQSn5kCt6m/AMLi+fE4Q9GEN
oSPAnNnt/SXeT1Jr29h1AFkEUCwfIpOgbEDHi6Uoq2LZf25W6iF0ZonH2bk7uHduvz879OO/R22/
eByUIqS9kzcUVdamq6cewwBKb1sXQJXs82z6f89/9z6zCZNDfLg1HJOiGg0zO6jF8saInlDQoNY1
/oNnydjEKSf9tj+0O3R0jI/3VzE2CwrYCVbrgpRJzTjkyN/uQ5YxA8pN+xdrDrRLHvLs14/jXP1J
zZMQktUVA+pYiJPVtrNP6krmbqkDXSP5TmvYYQZ5xhZY3pQ/YLPVct/8uLJjIbPy0TnhrQ/IvLyj
XV0bZDbzsb1TGY+FykZeWbtPLI582uTPd1d5bq9gCL03/hb71pwQQR2o9WiK4WSf+oUiEo/rPSOd
NnL9EtGXM9mQ8NRLLH+4sv0nEJ49ipjTiv4oJenj5xSts7kd+D1RLU/7sIFCteLbimRxWOND/bxc
l/+0U2Y8vk5X1aAqaAg94mI/PumkYi6PozTh5sbk+9J1N669vgRXxUXy/cHugw2G+0H9hRQ9qyKf
qbBNYVkR0mjOCilOhywLqqkYJ2nqWkQGAaXyXDmdQ3FCnFvvR2B4Q++F+WyVBZpVB+HBfjNbjkcL
deOEeOlW2OP+jAxD4g0jIXi6cDBlnNFr6J+5eVaYOpxlYiG70+f+e7AUp8lAANtYppUp/5/jkskK
kXTQuBVaJTmkr6w9scsqciaN8VxjTN06QdRPhPCBouGMdSdaGuMl3RG+h6rEDeQD6Wen9Xzn+xjZ
asveeF0VUaHvii+A3QLwpUoekqkNDWaaVGspkq2aJOFgsigVGCrwI8xVqT4eJcSBMykyPEPsEZ5r
zXntfXHjM6iULsaPM66qO15aq7SSdLck4V/5msr1BKG6Ykc6EtkktghQh7opY/OjXycT6Q32dqRy
bGyWodMEVfOISSSqXtD/LSbvyPn7oeUvzUBXQ/VNN1hSohSUyFSRvFeuGNxmXBtVz/lkhvLOceMB
G5q+DLAk3wW7IBF7f3szNAn5C9CDDTrTQAEfgEXgnxLK0iIiZ3iGvJzRTMicFsmPYxDNpm9SjB6O
F1tzyBQYfRn+4q+cKdS6VWim+XL8IMnRqDb9Y8LZb5d6x4CFXBZ0XPyHa5noWbMIIBlagrOOeNA0
fIDya9rDbHxngjavVUWuNzGHhLBBiRVXJJhikBUU+wXV8+H+ZDRaJVJyzEsdI25rN3V1O1zdYbfM
7glmyZIjf8T+3YpDW9KX6ZbFVCvvT8MX3orlPAdZ3rpxotx/OFUkEB7Q5A+f/Rc3k8UUaKDaqSAM
pch0e/TkV7LceOtRl7mq3sNTXz6Jm7cfLraaYHFD/iKxtIKMjMXEZ3hgCs8/PO0pbN1THfFgZWRm
l39Dsy0h/VpdHyxBnwsjBON7cVoGZ8aYG53/hAPkdckUfc9os72QHSytCIo5E0M04UJojN2QACud
W+Dun+yO5wjKNg/2eDQbBw1fchRrRAYaI9EzKBY2lvd+v/IhxD3M1e/HMZpAYDUghlte1izmLaLa
f0QdlrKxNkqjrECrRK1bctvzwmKRbi8NQR09HcU0fYKVzMDDnSBN5ZYDPu/ElscsP74rbyYilhXg
+X+W6EqpTllTuAv5uI5vGTeljgEnFf9OlyNX5e31VNMiwtkoXHFpA/qGdEWXn3N0eaPOdY+Ac4QS
RC9DEbfN2VtxPHzR9zp3MX8/OeiG3QtQCZlTZHFVQGdbDUDB4KNu0r4BBZux7RavtczwcuV/jCzd
WR1MhvFd7Fujiy91X6rR0vKWX4SnXa5G080bTOFl6iYZhgkrJabWHuSYsaS+a96EUNjLxT5iYbF1
WSNWYwAxe4dd/BzoU1jq0DKy0n/4F33++brAviNSb2/AbTNOJbP7E1HUBmk1sGjomK/6lbXfhBRu
mHYrVV2UiZezlMgUgFBEiH/ww9QwXr740YpWdiIwi9+kbfOYiTK4O/UvY8jA+p5Ir+B6aVbkqrZT
EQUHAfebi2xTxAPgyLOz2wabIS9Onm4G8I9dQyDXQKvpczzhSksrln1V20+Eh0VZXyaqSC+xr5Jj
HskNObeoK8hDTfGZVX5ePM9uv5YTWn7ueLrCxNLJFXBkuBzokrGucx4zajsjTFTu2M5U3fIno2Zi
Vk3FqmTdY3BgsNXwP7g0ed06SvVJlDFpxqZUpFr40HE+QL+mKkQkBuYSQ+ypNIopq1q3Qtl1WEet
an9EDHLy/gxqwGTMH3cEAWk187cZ0dzZJIzPIG5QqtmP+gmGwc3SE7g/+ye065yrb6fQiq74w8BN
QB0+04FPLiUWwqYuwIEefCIMUESDwJy8q5M5ETrbzHlvSt5Z1JRFzan3skoefoKJKb4ggkPy57sv
0M63eLRpxSng2nIVrgcS7flpmeD0oWNSFRCO5VQvciTkDlMdrnSIGl1/VH23LSU2wGsbS3NebFVu
WxaZhnAGHCMOzynqHm8hcbbx3lm6ckHqm32tmrx58/5ySjXRAQ/ph5erCVCOTpu7YnbZK/xv62D6
5A7c9JHjbBi1dBjd2/3BQDCKx3VjPdxvUWgt8jlnoEGjXevhDcyzKz2cjAPQ9yVxW8wMaULt4JEb
qE1x5AhWF2ODM0m1BRcy64z1hYlC1jOd+qh8oJl+RWn0Gb2IsAEf0rv7Uaew7hQBbxItMzb/AAL3
XAaU/Z0W+xiKvTpicqtYGpp4dlcWQBgKc+Tfs88F4p+XTpxKchXTgZkRwZVs3bVzq7+gsJWLZJ2f
S+LyThgl+Mu00D1WeiriinrGWHTWg+gzoEwp0jkQ5Nv/CgMMuTQkETVSppnTGwbeGR0NzCDU8jH4
WpM40Ng8JzkqgkVYUyb/zCIZ9cXDDv6nm9MkPEqu4SmbHFvV4VNWOhb0neFQWkJD2bwGogzNN9R1
5M6Eal1JYqOlEwExb9/t9LE0NW8f6EUSCYbSO9YA3NQZR3JJ56V0ajNfpr6jg2EmrnTtEiIMIU1r
sxYxUnS1O6NgeTdGFuPvvpn+RiV1ap3eugjDqeJk/Y0Xks3LzPZDB8Fn93M4pQTHRnCyD2p1Wz6v
l7xbtjSmnT09vqAf/F52H5OyMj8QbDk+MBT4+6WPzhHd5mBf41nKnTzfdHq/fANjXWMAUNFw3Vn7
fNbZDszeyapbxDQtGAUYZf3oQY/EfAriTyWIu6wjwpV7lRJiK71A1sY2tSz4IO/CsvXDk9LkmINZ
koJkNvT2PwcfL0LsRLCF8KZzuY59YT2NjXRBUDsMQVO4QJJPkqU00qoZ5nSnBZP6LR9q/ZInOJ3q
3io9marJ7IN8XcdZXeIddaN03IpFNVjff7cEeGQ1+DbQxbiFch3IX4aaTKcOnb8C5U2k+lRMvWn4
1lg1xKmv+S3Y7ZRAuXdd52vOgGRYYGUSfvVxUxELqmrfoUf6W5O0mhjG+8ro5xbAEZqpVeOxI39q
yc8NiFQB2UErWlVeppEQ1VxyuW5NvIM2W8nX1sRk2cngZSBhUZZbH55Qj0h6uL0Jhoxc7THk2H0f
RY6Hv5FhPvqGQX03GqE26Ax+8iM+RGA3M0NxWCeXpW0l92llff0WyMYjDSdYbIrUBFMI7uQ9INNM
0mT201vi6hxTj8AHgh/E/9b3YiythiAfBFgNJGcaI7osDwkZSWsuzifcYRZCEmbDnhSMUCW5soz2
YlIKFeiOBImQiGJ6BjeA1TJIjzsWamJOagPfePw0kLnl7C6Aa5xuw7zgHL6gjbSMLJ+UcAXh/e/3
cxi9za8FcHznccq7VSmAUymwr6tx+EsfmZVoQ3L2PkjEUHyqbt6VHhU1zVxC8fXW0pXJg8dxyv2I
bLIgvrh1Dt1KCw24G3VAgL2lOQSvAiLr39beIbHkML2PkxN2ZRWlFzsvo+0+7MN4PhezMJpkvXY4
YZcQT4Psuxldg2p8ZVv//1Ujk4qSTLV0+nw9G6WDVIk2CmQWc8b5xk6B12sLrWQAg1pWWxw3vLcK
/OMd3IaPzvmtKOyeAhJFZfB/8oKmyO7baChq0e9Lcwi38lTT7lYtHVK2Q6/kgGeoSDMpzTzoc00l
mf42iZUcuRNX0jMBDk/6Gz7vdVupi4CpgWPOcRXWh3ZVODFchH8dr5pKU9NphE5vTN+cKGqgIcJM
ms3vRzIDQ4Hm59FF7TfUCBABHkqgp/Dg8AXBgJ3DWVPuYuNris3PaGo/zG8NoXW2faWkVqmsf6cB
qCTmFnr4q+ounh+13J8uEsAsaA0u/NX61d1g6UTqVK9lYKwdS3p+GltvtmOzHqwqNiZCG3uWz2aO
ENLibgA+AHw5SO2rFRuyFAuIM/yKa6mXRdelxeicDOENSEXYyWqpI4v5lj76LFCskvfh1JshNEkm
9eHI5r/GfKxQmyZqpE3mpkNQ3lzapU6s7AagvQTqwjgo/xQiOxZO0VVcSqCC9aaMOlizi6rKJTWR
1HXUvAeILc6V1wbIh/MdC+KI8jOxmKaB2e7xDD1TbxYPHTkjqVXRtbbWlP08jhlYewjOrpHClyjx
7uktRNxgYGE2jxVQqMpwsXBPdglXZyv50fJ2szsDzinr8b37HbHnGUd80jNl6/C/5UXW3jZSq3gY
JsMrMRaHtS35EKX3BtAF1tkgEs2eeAcalo6iMAIhbC8KoMjbPEbzpQ9LtYu6EK2H3oKbtmEMoLze
ytU1GLJoaSedBzaOjIzRHXxdl0fZII7izrv1sYp9QMWj2d4Fb/HCxO8B1DMMbDQeIMNn8L8/OuHx
m8YWCxnrbTdi1i475K299dDp1PzeN7XhLaw6yBWA4h7VyHsHvmmUi8tUy2eZtY0j5l4hn0wtj95U
rzdeo5wj+ckDDk/wjS4pzc4UhaZCHBowaq88lY4G0QP9OjtelGjryxMHCfvB90SOUcguyWnlpueK
S13FKe4cxv+p75UF3AtFo3jl2vPmqcK+hmUjabQa7aKoXfjfO7L9OF0/PawkjExISzXh6rF06isI
pqXUS93XlSa+GC67u0Ue79iONx+F9kMaKcQj7RUiRyQTo22uSPyYMlu8qIxAmDraMHv+Ek09hdoH
JG5VunGAu9T0mVjqvQfTazKQtoz6j0bAKVOVyg7AexjP7ltwKDFA1P6I83qIRjnmMDtXD/xAF6at
rIvHjfBEJJ/vdgCBV5O73U2zg2A6GTozpll98UUUdNnFcdhtdAyYaajrhcqhE2duE0Gi/PQnbcHR
SNJn6SRQ4dCFMXFuDXCfL7n0ONrnhqUEaMYTRglPh5zU/EI5s1zNHzTtrs29yVenudh6Wd3Qmzy2
Eri2WZQDgJ07dNdiibFIotCBH0usCDoHkJuE/OaTEr7eCXxciZx1hZ+KDQ6wsqRWCXI52By0zAUy
g4QLfFqVDtBfRSGbmUujcRtGjLNtpezEzYeumXnEO70UE1JTYmho1wHUdY/G4aIjH4gwY6SaGXU4
uKhTHf0jnh49Py/CQMDG6ciGBjCE/FSvmV06uvpp3L8wzjnOqwZ1q3O5MSBrJ8F+r9+x5Y056qEb
ARMYdk4DhWYcWyPL6c7W5vsDC9Vh/2YNhYwyuxL8nsMI8hGMjMhafI9out2glaBEj8DLG3BQA5dT
stkfysWRBO1mXSMJdis4rKhKbxVCa/qMPDoDTlrD+0GUzdprhFFaWCw6VrWjBTxJQoLS2BbTDU/H
kxIuiMDwYfvzz6LlYMaEX/+7rQhloGA7+JVwAD1Z1WMBxe296lD8zbIQHhrnsQORm7vBphFSl6b6
kLa4h2czm2lzM7jC+AqEUJJt9IGms/IELNGe3Ci4owO9DIB5UgQSegOTqmO2VBOBzk/9WwntATEG
VXb1+T/tCoMhWysMNzcA9mhch9x5lPzNSQHteFA7V0Ce3rEVoT5sGbeSvWYQwJsjO6TshYlwlwV8
/yORhtTVVZR0wJg8lk1w0DOcZH77TKEc1S1f1bbcZs0LzywyxZF/JPpCs23tBPb9wsW7TaCz7rYV
Rz4ltshElO0lshE0Aq5+3RHuozam6lKJvtf3iSBz2eiFb6SJ8PIP7KNXcy+gbfn9T/+xRHv8et2B
O3lsw97qdHUk279SC/3L/a7NeoYQzM+XMaaIhv/uRu+1MgerIyUIra3+HXOao4YZLr5bQZWoII1f
Xnds5krdugHZY7occniWXaz47gW3fRZuF+pWaoTAFsWITgrtOs3ZDxNhl5jrKQCmFWJ+KNRWN4yq
Q7Z3AMJfi8+l8xh9SP8ybh2G3pjIEO+N67Mu5zCGahdYBIw96ymio6XKUJiRXJnMGs4hZVLfp3pe
803cyafmemh0eOUsdgh1daHKKOaLgXDTokE5DZL3uZbGQQRpyzEnNKembJR+/I2OUmH4cc+q/eX0
/Gwn1gtaQlAvrGvKJ8wv0JXMXvXmZIcicxs5RqNm4I+l8EdE6gnCSOnLhbQ/06QyVytdhFXWrwb1
hlPNXLBJ5c4Ws/f0RPYiJI0SZvYNoLXLG7sXAL0ctQpCL1T1IcgESeDYdU6TwziRiva7t2xAqMZH
ZJb+ofNkvBQlwUFdNwu20ZaFRFkEcpFKJzdWrRtdx7zVwPDgQCC9h0AwuOLB2iwsbWauQS1lQ9AR
NV4Ib+m9qoNpWr4p3mbABXnEiLD7m4RStIzKYiWmlMHb/x1XLnls56BlTcU7NPuNEpjGnO7A1OS2
Nrt7ehquu5AbJ4VrZOqB3VjXFUX6Ae+GnpEiT/eEcB4eIwFYWPQXGjq3Pr96SvGCuJQQa1IfGKVY
xM6EBAwOLooQdDvRUYDdGjaxKBsVXxE7SfMgo6MkVtx6LQliyirgC9v4ZLTKck1GnhDonFw54RZ3
f+u/V5unK1KEU2L0SzbkHg8NbeN/sMymriiLbpirITmI3Ajr21YnIfBllcHvyxiuhpy+B+0+ux61
i4rbd5BNG7CPNxqICjKRMmYQfJdrOn0Hlu2qsH7gkoMTtL8zU4D0xDgjt+zH80xB7UcTRFpPDYl8
q45xS5ehuXn8mNrSFB36WHn9tF9203OzEC5WqdbVPLWQ8DlUyygh4gW2NtdsbABaZHNIeYsIdaQQ
+W6Q3AbL1YRP8qt10JaKyCn8f0KZKn1FKxSoXgvCB0UTd+haYUQLH3+f4bmvOWpTo1iw/Iq3XE29
cObkgbc0SJb1isDCRy6+W0x7yF/6tNnZ2+60qbpoolOO8/ATwuHWgz1laX1qYfVgP2po6sH03Jbw
MVYGTsoV723RY/xtf/YbqvZFApm0PQqJxpX9tHqbqiM7hZuMqfifDUUyc6fSZ3TbUZ5Fa54tC4Sd
Rw48yEcronV9Zx1a5NTO+Cg+gBHPS4h1LSSAiykiPgMNGeQfaRPBV1246R9vLk8jDSQ4uwS3OoX5
o7o6zp+Wnb/Kkie3pZMj4c6SlvEOZfPkaLvQoZaT4FKadT3PGvyKP9iBeQNdmaGN+PgRgaknYuho
mLPUeB90iztOKdhQ8K/hnaHXw/sa6PH10u6ksXdWFYfC4jD+vG1ier3eXC+ltiXvDsR2/yiS9qka
HbbqhPDRP2O52Ur9wbGWFoBy3p3LE6s8fUSj+ZM4qwYnaCpig//NmVJ6a/kSP0Qs2mTr9Ee/90Oz
RIbBlfu0cpIdobjSrT2EVTVP1LnN5MBzyEFjA0bWgxy0mpfVSMTWL6Q9LAkIIkQjOe70EofvB0wd
E0+ZO7kIhZ5ZI0TRVKIa4nEetFS50HmXbOZqqDnW2PhfNq8ufx372oNy/ySs9840oSXutDJno/uT
OGNNA7mmyruwzzRIh0B+1ADlvTYzV1wgWTItfuMu43xhgg+EitBEc7gk16xuwYga0HzwJY9usgPI
LocmkbLl1EzKglpoRFe3gjaZfaWJWPKc7Rt700fc3KMH1xWx4LOWcwMo/Q92spHSmqWj422zMSKl
cFouBGAdlUyLACM6TEoqZOjTdLCpxipNyDfZBcITU1x6yKCJ8onigS4h2RA5E3P8jbb01Lho62gf
O+OGZA4e8JL29fvFJVUTmtT3pg6VXHGVC2YBbcE0OEGF0xG5z16Z/QfaEDeUtJk4hpfC21lCybaw
wGGn9Hd6VNmaKhyGXS9EQ4ipzoEZ1gBqf3p+KQ/Vknc4fkOhRsQk3q6s5Pj/ZULylpxp+bKIGrtN
pPRdOfxd6uckLJkx2NRE9liUCChjeHW0HdZ+sjfV2ciqC6uNnSfLE8pDiS584v5RWwUcSYtqngDe
bkY7ebl3pjHVVmc3JIqOiPy9QTM+nLWYGxUNbPEFuVpzbz2zVYxNJC756FPHumBDi8s2gFOf+GKY
LGJSFLAclv6F0Nx21mnMslG2VHtHurFxCyLj76G2LJvzqYfTJ7zyzN1+cG+zSBm0W5jV7vzY6HWi
sRoe3a/a89aZ6aqu5f2J3r4470sRH9vg0A6FMQIEDoTCkEFHUFj+g/wcgeQunB5ZUGjEpQkhX9CT
M+/Ze7hGRm39BOzwCZydN2o/MkFg9J+6rz3nqrt+rSvzXTU0nplTqX3zWVpa7z2in9lv31WseKT7
AulzUe6ktua0kvnMRJ8kA8JPRp/p6QDFUNj7WzVcgrJQI8D565QB15TJKCI3oWfma8Ch3A8hYzYp
wxGscKpSU0IaPmlbtGu5YTz86LDJ66Um1Aoq4+Uq10N/LFCA5KEnY9CLbFFKVV4EOxl4tBXeSE6L
IJ5hcXKzC7n48JhDXUfqjXBmpvat/+iY6Us8Zn/1HHDhRtC6fgP6zBzYhJwM1ZY4bC/KZkWbZqAN
nDT1t1VGQcgvFOhgCmTIEhuEgsBTE5Lkkj3RhlGMcTErKhz8a66OX0TNWE1wDGSz0fYROHPQvfYV
SGUVNP+urV7AlAVzv/PMjptkn3JkXocc8HRlNObWYEljGQEZ/FvoYxUGkmGgH7OVq1x1x3qKrI5+
VTy2scL8Es6YVTtF+Gw66mdXRk6K88Icv2YaXQYP0bHJeQHvyZQSPoFTPxjSK02mXLz6a4T4NG5a
QJhcVR0iiwmo2bl4725bA+mdwemxRaKUR/d9iWxFibcYCbjZ1damkBV7dTgVkfBoc45a3ndKfH2f
F+Qk+5ZfSbxnM34qHaSrL7LtZzbIePcy7sUDUkc57aJLUREKh/kevGX0fUMLlw5nGFL8+nDOyaTg
3ln7TGmbxEje8a6o1Bp215Eh6qkcq4nLoqX26BHwVnXR2PxSuKNX5hdQmwdO3Tzl1XcikXPw2HTR
Kqv3IukPP5aQUQzXo3fmr6OJBxP+Kv7b18pNHbHdGCOTBOoCEQrF9IPcmw7i3MfPZqdv/qtotHag
cbqzvBIIGfq+mH78jYGhZM+q4f8LhAY08YkuS6ZEppdIlfSUVidKKkGTqw8l5qAOY7fn17cCz6FB
hmMAZlCkpuuebLJEMZHlBJuELKupNjO2yulDrcrcj8PVg1NMnha6v2EHofoJyEr76vwDD8+fCRCS
cB28HXtU7+BNf3JM9cLmBBcBCnR60WhqVcl3zRr+l3V9D3XUZRAR6+6Jn3yVTw6nuD+F2YRasskl
5REvO0jaijTXtEXAu/z07+DlgyOWjjcaE66YdvdgqW99Tpa9qy1h+EtWzNBmxSxDsuuU65QyiRA0
GXa76GcH1fFMwbik0kYPrSqyHqYvrIae1nG5OYm1RC7AoNEZ4QRnkJaNg88CYu5SQwoZhf0Img34
fAgSe5gJJ3LGsqw/sVAyU6qMD6b5z+hFu6CkYXhKgMrvYqUGKzEVcfiGRokU/bygWte5Rn/FzZi6
C1YY0S2KkJkrUHxvsiMM/HgG23Nfluznxcb11TjrwMwzFY9M6KVJ0MSOceJzIhpVQbt6qp0I/EOn
IIBryBzt5tONChlisaYXQKJRp9GI6eRWX+f2bIxSafBOfpzsaoYG6NDvEpikR7RiQqQ3OngiBx6D
wePyHaiWb/siQD2p1onOGbP9rlhY8ySIYcW/7KiqXg3N5uIxsM5f0ctAQ4bIfqsB30tY0JdeaP/N
GJpuSSswP38EyuOycvU7BTxviKCoZPEN/CaInxHw+cua9joZyJOvwJMx44PtDXm63L3wbJr+JYCw
xlsvMWB1iO3QKglMt6Bv10HpBsy34As9aezCvDfBUJ/mQTaJXsKymwH/F6K2/6FSU24hza6Cuzjs
h5ZDN+/R0+hOp4nPLfBO8CNuQzebEYQ4pP+qPTJxeFYw7tLaPo1kIRD+RPzsNIDe+G6s3Vu9wfE5
GRZ1NRV/oquPpWamf9IjyMZScQ23osSd2rU+B2s+kPJsm1hLOta9YmtBPol0A/7DSv9+nU3+jD4g
3/jeJ/v9q/b7r6q2vz0YjaBxeip9+TGuH5w3iA33Dz3S8aMXzQQv2LsCtc8ULH2IHFeSs4+knyUm
R+a2C4A6ZwUR31agr4M1G0g+/BhOu2WQcx/R3yIz2PcHRZFtPgng9UWR7oyr4f2KS/9avInKAlur
m6grh0DMlN/AQvit7nfi5wgrGulkg2raId4DDBRH/wept1TnmAX8lE0oKdkvnAymV1RJceir7HRb
kEERSakapGLXNyKL5xQQ9rP+WwH8VeHM3x5J1t47nDBuTqHBMRR6AnmlR6o4i5MSZHsM4GX0I4Q+
1KfYRZz0CvUEQr2GUSWr49AHd52+uQvEgTP6fK5TW2SD6XUVwhMdCA0Goqu51qRLEWFd7RCW65Pw
Jg4pVY/d5tOv7F02d1YeNWANDLgIHV5xRLs19m1qank3m6ffIsVzWftqCs5KUqvo+MmCA3heCFRb
xVN8DI6XEbgDlCiBFzvTG3IEGMAMd2CZjhLHgkEOFmaeEL2VQWsDPYtOjM1uYvhCgDj2gMgLPH9E
cqU43PBcsGij3dwpx9MhYoAtOBN9J/60KXymCHI3ZpgMFVELqZhOv7lNqOwjCquOqztRAy8GO99P
u2yXmAet/mWAEfJw7WFkubImRJLIrhrSoiLFjFPyFzMMk98FoZxbBq1CiSbZzJsy8WZX6mvWtGFd
9Mida21iHAzD46wRoPeksscmj52Icy6oulVRNZzZnhe8aF4hcBSDBSPSLxiHYAfqbzSYUmqKmhxr
TXBInIU1tTHtERhhW4t6ylSTSupm7pCZfHHuSZhdDSezWwKMppa8Oyz37cMBaEmeHRX8vuGymVmm
b9wpO1qw6AL9G2VdBxTkRuh5J5HuLri2YFRDVsDMHJpzYbVxxxJZzWDyRV6AG322f9XAlChs/a/L
BkzqtVMNrRyrrGcf6/TK+/4+7Q8rZP4YY7gt6FS3XWZ5z70PUulw657/qo3kbWz7Cgwfl9gqUO/o
cgYZepW9ISgq5a4ZeH0HbsfBAVYB5qzXBwyd1ihXdSEzQ9Rv4WHswuzTmYCoh2Qko9UBPcBRwmha
DXYrVaXWIGyX5vSgZ0BjG3L0bhUelJpZXCvDQp0ynUwzxpcFg/KRgXSYPjd+2zrWkdzC0XgA87Cl
dpALyJrbi7wji6njrVIaLbotNeE/IX0NU1M4lW6ICMQZGi1DtP2uYcdgHq3zGibtQZ8+q/xZFNwI
1PZ5/ggWvxkXZuVwk9VwPUMotJ9BVqYfA1o+gniIzPtqfIjQvVAOKwIZG5ap6AgWBimA/QwZxuh9
QqfVH3Su2YsYRrkieplDk6/lX7kS+Rt8AdVpj4dhJx6jnj0AhGeMj/AUwvktujmKyp0FBkdvSwQr
hWPxcn+Eby57TXGk2WGC4yEaoUxUCFHwr35nzmbSuAlad/6iytG/+7pAM2IVBbYLxaHn3ThKhv0c
q8PpWpHHnBdjccW4fRUcB9ldaNSrNtk0FAkgfs0UdJluznFryT5tDXbISnXzVZ5XZQ8xwxKDE1sd
fj+MOmLDS4znj0gbtCdAOPFz0vB5oB1/TT7v+kzKe6yuj+3Nv0mw5WTmDVYl+yZThi+1oEB+7ugW
KiVU2Dd6NQjVkHZCmh79wboZxVZzQKEmFxk8qQLy7aTQDudjPLkSlDatZcL1p302ZgXWpXwfxzV3
jejAtLs3z68TeRd1HgdOi6f8z0OotCc4C7ziTxUfqfgjHC1vp1CwAMqW+ia62GpNq7ul6fb4wBHl
heE2YnAL7jmXh1f+LQOPOediK4o/eT50Dk2g3V50y/m5QHWpZjyTCJi9vO0Lt9nRuPwiZ6lvV1oE
ReVygqWbfMVwX06dO+l4nEFkHhvLn7QomfXudG6S5NoSiAL49x6xCzfGAl0b9c4EHxsM+xWM1d0+
YNs7/0cuMohjeIcM4oY4XIFVDktepbJDjahqNtSxcix7S/R2mvAPxWu4+ydlguxQAXCp7pYOmAdc
qpYRhhEg2o7dUWleoKmydmw4T7CVO/ra/Elv/23eGOuVLwk4Se7rI3FWGzSBgCjce960G/7MGVvR
Urakqnr4WzIo2Wv5GA/Z6wtv0EoT3SUIdpZPyiTJCHVuGSm95GYLh8Stp5Ariu3FHX5xI3u5LVPY
+EtPXWVwxwZrxLq/L1jVb9xKyp4HGq1OnMb1C0u/7MAT85ubekaa7e6hXmK43Nf45m0tOuLpsxq6
eu3o+BxCrZdVnUX+7hQUS9uUtV1pBXnR7QgFUJBylqaGVEwJPHAPM/TpR2XD/j9WA8zM6dXrc5v+
P8HrTzc+9Qz5Bj/ZO4JgtKo0gZaWsKd6Sk/xVKZGDVljKeit0WYB/eVI2ZxlURBSnrubOcHDz3PH
UIh14G/GqcVY1EAJY280Rd1Xu2Sg0Lo+mIwep/dX8cy7B76LxmwPl4VnQhZP1QlytT9rIGfm/Qql
LrxX4ZHhOSVgYkvrjVyKwp4wO4i4DQduroN0TJ1xD+b9A6BafXksktSOeS8e196oRSiP/WT/iqHF
knMykgjPbsHHedu3KSh+gXYaGwMYKNK6bGRq0F3WlQCATeqGRc7OE6CkvGMhs0zydu/QW52ifABs
Zr4PZnjD6I4nvkHflnx1+9KmmYL2Y58DpK7azt2l/ZwwN0QVJ6bkKIp55ozeIQo384syF+ghUPtk
ahjYaOvppyPgZp6olc41eDTIFGBqN1TwDK3QXoBuE6OHwqKPS2BCQNS0Rf2fC45JpWPM5ktqVFpW
vmu/fAo+bpFxHAf7mLL2cFVNp3qm2fW5Dnzt8b9XvPfdW+nrbB5yt5k15l+f4gSvTkkXh0XgK9v0
MZovc3+M7vKeEt/6DyWkx7k9+IFTCc0zhpwxh0m5ZI1CTqvBj73FTZ7nWthVGCLKRlm1zLpybFZe
TREbzNgmjMhSRrkzwi5tQHhj+jkqAKNFE4YSDvsp0+cTbvXH48a4BLW+R5ggzL9rJe6jVjlW6n+s
/fIquH7suToZ+OUQ7NxBPmiFTzvykCYVVh4t4R9CPcs9F2C0rDsBgyP8I8Bxi7gWfWfRUyDIQvSa
LZMuscroXul/r1ubEaU435TjnQ6OEj8Usqok7AU0MALYCbIoUqmO2aL9NL57xN1hY29FPfuROw7L
uB3Yi5FEhhVeUA2UkNnJyrELcbQBIBclZcHWO0DmC2IUFqpcpv73N86XOK+Xe0hXSFBpsfgFDVq4
EREjdHxIZx7UaWBfbW3MJzb4fARTGC15bfjvJipPiu6Wt0z0i2TfhEYnNE2XCxlbdOVOvu1cFUce
tMyGRz/IJpH8lmDVoYhMwQchwAkvIpf+MyPX8DNjtAsNncqcVgpKUbiHl++nJn4SGaiswc92qeQ8
+Oz3fWQ4i5F8YevJksRNDi5I9G4q7AHGr/6HdDtEHxmU9Ecjrxixl71vEs4SopFICtyRJZ7L7c1O
NZU318JnfA/fW4hSeOGId3IvgeFEi+B9Aropivl/+tORXAYy1dPJkK0+RbNCaRe6Bu7/w2ASGL+H
9BmPK3eHK9TwtATFJuSKV3lfL00OulFguIhS9elx/f1oVoIBb201m0aRLUtpOeEdbn9Oena1OWP2
vCNFhFy42M04qECD1t6cdZTJQMYjL1itoHC7pCxRdr3siK0jnsr53YeBqquupWBBRNi8Dw5eC875
QC0VX6acBoTOP+5Kd6ZW99ssPwReg+EbPNmB5fXKcDv0VRMuYJWo5giZr3p4YbK599hrD6JWhyig
B9qmhINPaUxcULJjF/sD5r1EzlGI6RvnoLiS29P7XWzI/QJ1GzuHeKE/xuuHQomLyxsX8k4FO88U
vUVFdniCMeUEJ4hDbcLU0PWKpTxpUdrqNMhYIa5WU+4stbivLvI1iGUbI20H6NCzaEJod7AFBoJw
viwrd3Hglc8N++k+a0VIQX3ZyvyjMZ3J4xJFInp4R2EasiAb9A03wdK+mykWHKVU3CTernwG6ZrH
5mihirHCz0E1Ks7bKyYss0Fz6NyaPHpqTGznSc0o88ycy0MceYXgBo7p+R9uid9pL2OfWtQhv7Vk
1Dtt1r9/u7CTHnyqmc2148lqSnAWiWJ/f5NCIhaKygn24vV3vGqMOU7lRm1uyfNrNFFsZrUJH1pt
xRwJvt0t6Ms9cDvjf/4AF7n5QkDqMKjSzX0rpQ3aooBP78blUNWd/U/TNSWKdwjEsBLEXvXYIE3u
vPkn7nopqD6no6R4MJ61tKg8IpgoeM3fcSxqUwe7R1gFeu3kcfhWB5RopGB62KvSMJUMlLYcK5TK
kFwNp/xJ27TpixxaWvCLL6z1Nf+dg3if9Rl3hgRqARktMRfoHnedzyfn+UL8cckbIvOGMf2RY8+Z
a3UZ/KESUVAMskjUYEHP9JEdamb7R2RXp2kRpgL35IZy9ujnzAlWBlylB6EUao8kqCUmrMupZ2Wc
DcTiPEUjV7pWJ03k62+P4tUPZ78U+Ha/ytuJNlPimzYsF3sGz6vuv/8EPl5G+ehCupbXeiJ122WJ
RrRR/+jg6B2tLaexLkm4uaFGWbDSnthRE2VoS1+Uurc08CmyFNxZ31C655lLC8ISJ6AEjMVfeuqe
5B/pStpI9ZRsN2kEkMfsE3PkuHypMkLz7SRGy5TdwhThs/5vB96klyP+9E7NYZ3T6fwQNoLn5jRR
Dqf+4rfFMJTGDtR/JzTlYR/92O7s/DWXgsKHPYfqIIDwF4xYZDFUnO4IjQcY3TkkV34Aie1ECueA
7W/4OMm6up/CPESrF0iFEYgXnboNcVBG7dj0CBPI0jK41UcLYnyFPwUuWMMKm84SBFJfhkdRqbuZ
b9iu/dMtAGoy1wgyr/OVZXx5soRFdoW99JOdvN6Fmplky+SUYSniXGxbzNQg3KmWkGqM5yHouvul
Ft1FwQs9SQyQVsX8A778jBXJyHx34MZcnZO+K4O3QKhnWzqBsg1s6pQeuHVswG2bQS/Msm52xRH4
C51XjFPdYIXdw9xfGTUxVios8tFt0SBWKfONYwOHyXLdej64Qh5Subqm5nzKBVXdH1ESJcFxBoAu
7jZ41LMacvmXhUz0iiWdx1Uut31PSdk2Lg6cAb5/rxnwvuUIBl0V2My+g8WaReKKpBXbs5gPDPkx
jbicVxRZKLKNl2Ltl0y8xb7rP5rifC2Z5nOHVcOgp7zlQPWtpzuEg4GWx1I4tc0awow4H2oeyPHL
o4gxcQiygl0V4Nc6uVGD0uZIbt35sU7k42zbid3BblnQpJtT7ayf6J8rX5HnQ+of2Dzkd7DNws6k
rDjjzDmcfCGsA4xFo7KB3lNCH88xhgiUzPREQVvaOdxD65P+SYfKRcwaOJIwXQM7ALtPoX9vgco9
bjEIeKzTDumgTubqpFPIdJIRR6MYSCnEfDBy6Jtwgz0lWwdda2kCeCuKrRRtAy36qJssfGT73Va3
HOJok8+uEM5JVfkpqeKnvnP1vYGGswzhn8q/zHTqc+mhTwMp9gEpA30bOopKRxwaaE3WQmaxE0Mt
oqYLWYu9kmpKO8UoCAsQNUldVlmNLwd072naWEjVGKVRqpNx/Crflwmx9/NMY7ev5ENdjABIvFhs
GXLckSKEZjVn1WhsMfF1wUXeEx7xCVfo3dqhmsCTZ0obm6QYKv0v6Zn+xrZIEh4myHBXKilzAM6M
lk8d/snB+dFC/V0faBvHXMcSERC+MR3umPG2JG7EWIxqAs4Hq0pK35f9W3E6sihc5KkQ2ivondbM
p2nHfvGMyHXAzuz41eA9gtUrfHEYYzfIdrnG1qdTV/P5TyToO3vGPN8CouL8aeJ/ypcYtqgtn78C
9nT10iG7nuBrh4jYyQqN9ysui7U90lN5wZr0ZYE3pRgUr0dZx6bvKCHplOzg20CV1VJyC/dqRRMN
PTNNUBFXdgGl8C7VGQdWWk0g8PYF1fTnuWDiwtffKG0l4KqgiC6U7lFT2UjmimMgswZpbzt7839V
pcPHqSdwhrcdt2qKg6OMmwRSJIfgncnAgT9diEIIgvJBdNSGk0S7smhXrl2wvQEd+NS+re02N4j8
0cFkiCQeIpONBpxve3NMZMqTIlh+qtmuMgXJhyCOh5xGF8SnFmKq5OeW1LXZpVazDeGx3u+lIgCr
SQkElMIr6plowe0Ul54Iw0Yzl8wdp2AcWCiehihZ9EqTcOIw7GkoKvB62R8ePXYnl83/Y8DpWUok
11NONEvCk+/a/PjwYiFgygdMinexhABSV3mAkgzQj617KXsAHlho0KbsLbRUeiAWCXIHkwhLBzqy
SNUABbjkO2qHCBho0yzjUL9zo0T+hLt/Nw8ZDe/JuYG7RgedL20x+HOzBP3zjIG1Iq+O58KtlcDn
Md+PAK3GDwaOiOmY2fI5Py3pzSEPVEy8LaAeZ0jcXiYvAcePP8AeFy28INT8yhYKSiezl/tkiisl
6yO3veQULwfOmY6pb4qO49Wgc9I2MjR+4VJYUUARK9wYp5Bq+LwJshxvS7lrQvOynxfUxrPld0+W
dI5mvQMaroVh4/+i1SdlvTFjG0DhjCCmxjZaEo0rMYPaqWhjkl0Ol6/Qe3lBggicCFghMRgDKeVf
iPCchs+Ykjej7Aty4d8GlTIGwEWdr2ixXYJAv1LVAEiaaMrziSnTGX0pCFGX/FbjMI4rZpz/Dh25
Op2qgocRjjf5YV3BGAOSCuyh/Ef+MXB9z6GXekdSCONjeoox4HKVdum4BRem4kd1aaxUrpG/dCpi
jWoNE6eId5llL3nrb2XmZoxrRc2upNxkqvGyur7DHmn1h+yjDjutxQVkN4sdIeYqhlgclygE5Sgy
cXDaG5ppaXFYwAIouauAzDU4XcYbOb63+CHjP3jiD19re5wRyTkMX2Azie+49UXWu6sbVWJUii0z
A9bmf7wgQvMvZcbAMZDB4xtuHMM9hPZn5+1bEQ9oAbScQOSaHG8zMHGaC6oj9NgDjpbe8+Y4RXYA
7+3eQ2MLnytPwOcgjXzHdRDetEktB99EkObA+wpqDbMuslAUehpp3z7bpAv3BKSgODx/U8OOol2I
jyKfR79CrH+XgVHeitLhXG6uRF5o7jdhCmZyyFzvxPM3ZPBoknbufsYTvn3EOB/ckgN7hpAIDp1N
1jzHX6IaM7c7WcCcLW5fjLfGUmX1rVTw5cl/3Eftkm3Lh6O5nJE3BRPY6c2l/MGGvsfdcn4MBxwK
0c1ibnN3bTOpQCGDJQ9sGt4y/PDS+dQpoeVWHgmdXkaBluqKbbejjQNG9EGTqzsf2ekx4vxWjNS7
FcdJSBjUpzVwbGNYtw24MbwH3eI+r3/EDUaUGmvFQw4WbBVDsRpINeqI3CXnzx/YUZqslmDJ43dA
nnXacObe4KHgJkCYe9CO9CnD7TS/pQwrZ5v5FMllfFHM4/CBlaCrxx/5Ym9j1RFGT4OL/sFThjVG
WnVzzNAh8Gq7y32RHSq6gln2GDUci5JKGqYIaj87P8Sz+Pr5Ea6/qqKgrepsS86B+pXmsYElVFPm
lM4WiNWgSVZIaxQ56MpawyLcvV+RPC42ilXWzppZwWfjfB6dnImtUpT0a6IIPisA9JDPF3BGMBy4
dCCdDD4LljqhxeWDiPr0uYOqFG+wr2b742XN7WvIXJSNVtxAgnovAw+4xlOXfF/6LyMssvQiAKES
VE0gN1xGQ9WqsI3XysOH8inYHGnReDtM0141tK/WsVLIuq1e6rY06XkL/ndYiD2z8iC6vGWUSrzA
occAxv18OsZPtU2/vNjteHHx5Oh03PV6/IyEaABaDdH6OvkDAe2hdqpfspwj2RWJco9xGrjMtkxa
YbBpijCS3y9xmHqXHFaTVaE3yIQvfi/lFZi7OatGLgyxh4UK0ZuAr//58gvhtYkvl9LyXlr7oTIg
CmSET6X7G+gRyaKR4Hf4ZX6fkA6uIUgfqndDlzPhvGk+VmWKwNWeyc6bXFUQ2i1MirsHntp34iX0
dELQhkvWNc+h5NDksIaFSVJ+MYZkdC9Rc51AO0zQerrQm3MRqVznFCp1WVwPMT0gwhMy+eWmREIy
QqPNeP6xhai1IHcczCpd13qpJ1uclNFSsSxKXi7RwA7mQaqsztDXz02IUc/mr2MvlcHQCWZsJQFV
YpV5UgIlcwvnJI8VPNiipZjeQbJX2Z6Ldu8/c+EHteIVm4rho7eGM5FBilf5v5hUPOYh4OXbQ3Ef
OfUEEwaMD86FxhwnW+d7K2g3P3rFVOQi5Qj7F0q/5i2r79HVpW6kQT0/XysYVVU9sRDidA3CP/xh
VoRMcM1ZebU0nvPIb4FTGs0/k3TNWboFw1K3XjNuo0IJnjF2UjZQZr0INk5A/RyPx1FJgnMxn5n2
xVqFftIkKxrOjc35cGwaE7VfM9FGx0Zt6IhLmuCFFOsujkDYF+KmRxK9hqVmIfnhSfG4wmTUx/wB
4I1+CC6xrTefPI1+fS7nRbRsak9eCguPRtqqpIg0pB5iMN71teM+n8kRz9lUV6wW16onuHgH4Wag
fjTve7Q2VLE2xrE8NkFO1EzstkJk9wyGv6AFBEYXC1/jVomkLv04DE0TSNyt5T1wrr/Mz04LWzJm
jxVHIOTkKnOcipQ/7sZChXsIATwDEJYibZ50JbxUIkKeHbaygL3Z/b+Inqd7pSar715SM4AJOb6j
75Ad0elda41lqipbkuQoPc8zlVU0uXhBVNxpCbKb/krhWtbEP1Tg0X6vWYQQdggWTDz+9KWBetcJ
3XUDMMNNAUo2PLmXG1X9VSh6BZJ8bG96ofzTxT1214hVNZ4AggDvLSW8B7XwB7c1IDE6Duj4m1Wa
+895csBOBg5E7dODG9pCg2pLNGnEwfZZs0t30657l2vtzf9Ufq67Yd0xk6sciKrNvNXzxEbTMJHs
YrD5I8u4gBmuf97O4ri6u12q/FNdpATRRlwLCG0pz8anLenM2VLDupvkIaVpcWpj9Bmt6Y7C02kM
hhu4qJEGcowLIUliz6cZdTEtECFcuGLfFWTHkwQ69IH2cdOEn2HkX17ktKu6TPxiZEBuVD1XXYwI
CBR9BYIQoVZUNneTCKLyiAgfCXkFQ+Y0tjmVuxRzYQF2i8D1vObkYuDJb+z3NzoG3QodDjkD7+oM
wO7SrP0OfVdw2SYXobOM8NuL29Dmqi+TXc1LxXNLdzsvIebzH2J99Vk6u13hEIopYBc2Tg7nkh6U
MjyLFGQun9g7ns4LAwlUeZT8yOPq+imNVY4HUILUuU4XcRGcaj7+4qi0YZIQOQjBPy5O5s6rhD0B
V8nXgrRNO1RS8BzPE1mmG+QBtzOc4AQFOgaTkMTdXb+MFyozuOp8DxRyDT/9FjiYW3aWwlywifpz
/h60cUOzO/9Pj9xM2zxweOhAYiXEw9niEdxU5M2joXHGrbkJp6qr9ns9VVepWGHMqsQs4bLOkzwM
3ezv5MrEhVG6JrpMUU0puhhTAIiOjEMX4feg0Tu024YFyREyhtGL09QmfEN3pM/SUetg3WsUpOgO
pUjVng4GEQiO3b2VqnbDj+ciZrwrH2U3vHamrXIUn3749m/IVAP5fF4WNWp+dUTs9BbhrsTbNvyu
xFbJFLHdFmUkVtAIj9nWbthkeVx50xrFSv8floBcuJkKyFX7n5Pgz7xn20TxG6HIxMACJJkzGhdt
3uLR2tmzbwCtJBJzWIgbxdUg73f6BFod9qtxJQJVmBzYa9qKTeM2WBF8EGiSRhzDRvwCRgWZokbe
6Srocr2mmXJiqD6cYrJ9urXD7pOjuBrkhHXEWWzaseSJjgVkE5Q8AJsm45o7rkZX2OMYlpwgcNk+
qcAxVOymTMsHyHTvuRPY/AL/37wiaQLHPvx1Uci5uc8hOcY2PlvSqGmyzAId25uwu+PRsGqJXDhq
U2zG4J0Gb+znaiGrVaO0sBNe4wIRcESWj3fBGeLQE7cNwMFz7UNLxD+9nftRIT/ZcZxGNsN0Hunq
V5wVMA2gqjk2xMSBXFhrMhSjxRo42dmVsP97tWjmn80Dz2F07gP3aa+VRAqxDUD2EZG/1UKXzgkb
w/q0zTfUvt+EOMWeSoyi2MJsmT6jIXaZQpp3l6SUvT3sNTe6fsdgl35wisyFPG/L5J5jJowx2oo7
StpHWalZWwQkd4Sw8fu23tLIIDzQBT0uYuHflYeGdaP7lGPqxoFXl5n9+Ngfk5chZcY4mbRowEJx
0743nurnUR+xp1gKRkhi2DtAyo+Mi2WlLq35hJfhHunxnRKuyrnDVHfwZPX9+ir5amzjL/rXwqVL
4KMTBFEmvTu+rQBitfH9OgdmAI+/GGoiBNzy4xWjxMrlU75PJqns8fWax6MWOeV2pHzn/+NB7L1B
YqnJzJHdnML2V1wACH+obVKvYrIPOHipsQFbiVd3OS28z6/YKpW28+Cb6Lm3bE63vOWKIC/fmAtn
c7X/WCVXQfRWddYKQD6rIjXfm4jZWCSITje3a7iNqI/A/O5OfbAjcGoeOgft/Tg2nY29VwWzK+js
uZdEYeN2V0p0ktjZ0xIt4ayxpb1fznWwR1Mmev0d8dzGXVZEIyV5C8qbA3Gtp5N4ow4u2Iyozlsy
zecyiz75erPYTyROUlOxkMuQ5PNSnjpQQEYnovfbFuSJSI9hgfFhfzU6ucVD0g8wIq/NfOtTJiva
siqoV9cbMc83ry6g49cLzZ2uxI5BdO+RBwEYnyX2u8fr/5jFcuv91KmfrkXVFoAogg8v3c+c0xhO
bxB5mW+LxdbBZod8r/KVqwzcG3egPOCKipNvYAkgp0dtNgmIu+4wCmTdc2Dve3CHc9A/bjw8mcU7
J9b/zlDDHyw8P4jq8KjGIR2qvGvUy7SQyz8GzLnrtVxPfjQoLrH5oIkM53lErbtI6xCxI5DTUhw7
+bHQwXM9FviztLv4oizVHd30LlLPuBTFd0L36F8Gl+zpKSGS+NbfzoFGWxTaAv7q0zHOLnlaCNW6
ZAQtuibJkR/Bol7QqOB1wAyqX+fi7y8IRHQn5sLDEFINEgRyVWoDjo/BA+THLLdye/Pfz7qpncYP
py8HCieC1LXG+jsq02ACE+0/5R3C0lm8J/68rXaSbp7jzGFnLNxc+16eZZbFZ45lJoBsyq0Q1ZT0
Pd4e8T3Xd+QzelyMkUpeHHyzViBHfw7qeOTSeo3m/iMkn/m3B7KF0Dujq0yIvGvKMQ3MdNrHN/tM
VqPAdQ/c1wfhePFUJvUJMjZ7Yo3JJEQcYdeG/97JWl9Ckm8E2aWzugjV4kSNrP8bgbE2hFFJvtAe
wAxJFgyv2HVwPkpLYF05rShfuoVYWZTvhb9PX31qTdfa1cIPGQvRFGxAUsshXd32Jn2ROue/876u
tpkV+cTkAnvpZjDBcgFMGEk9ry1DIFr4VQd9A7zQlBf50W0BPjy2HlRVdveUH9x0mRbfd2Es9QoF
2wdpMYkWxk5N3k6R2u1FayYVhRlciAyTMBX8IFJvF2j+537BlurhX3FpajXMJzJvgu2jwk8DWFf0
sdEJAM4ywmvYNcm4WgK7WBKAPUHtnRv2YRkVfiZTp/fjf6RbpTtWvYGqpSmpjvE9Ro1KSpiq0/4g
4i8ltE85fxyPuvurHMMOlhvB3H8kDCrk/QyTZT6cGjfDuGyeJBpVft5ttIz/oBPjH4TOl0izno+/
0RIWnS5BThk0YO/NJK0lksNnYMJwov0EWl9bkiOczb806ORmjAqFYp0HJl/nBOGgImc7T0I9biI3
FshGG8rbohdJRS0vhpfmtTheZoU1HrxAEP3oCboJY+BL/cJxyws90jy6Oq7d9bgyYSIz386Ap5cS
EwFhyr9Ci3nhXKS82cPZLNpkq10nDDXNc9CcNid/BBkqWSG6N6P2Y5jjfZUmfyPoZMqKf2cz4oSj
5Tn4xvRAzcA8ZNWW9GMw4NF6GLwHbRrSyOJptP/wUA1x7qw4uOuFlwbVcrxh5GG1YUiqIFV16rr5
GvyWwwIM+p9GKrVLuCeO/UzfxKSj6y51pz0sMN5Shy276mhzud3QxhUKkIl92XYa841Jh93xFFoo
45gXv85wmDQeP8Gt7pcMJPDUq0a2uCTc3WaCuHtH2ouqhwGJieZMZAYEPOvMGnygJ5pdyvDgLDT6
fUHTIWZJ4lf+u2KfzAf4cVbvOPKEU0DduRecCZddTnw7I6Gww32UpyHpMB2LWEB6GoY/iBbbmhm3
NUi8PefMP7a4FGtVXOquGwWGrWccGg/IqqTdm914uNOeZ5hWitHI/4wtkpvyWHms57BfBNzN2pAA
QRT+zN/6AuoRkIm+ZwduELbYRK0yPOJReswXTXPlsgZOi1sGM7uET1NMNVMEDW3CQO5UP7rJqBXP
2P6uO3K72DV9hpMJCa/Aiw4vLkPxXFnP0H1gYJh5V9v36Op6aWR83MSWUT5z7g46iAmoOri2XIzr
OaDB7fl8vpWeQ0yBmLuFrQ3oaPnSAZcHV+iDAk92hqB3S+6KeedLitnBRy1pbw1waewmYns7fDw1
fBz6hokc6s4BY1mxjzSU87L5xa1v6yyQvaX2RLFL0LLc7kkXRSpFNnVZOxjFPOBE4juLvYbkXo2v
BTALqjDMmgPRS8wT9RbyGBVrGmxPXZsJS4gXuzyO2T2xn/yNb0jKlK9kPDlue+C+WnGHCu+p4CF7
Ih2NjwTUGNASt0oe95boafQGH3Mth/ekR/QFCUBz8FV2/3eko7Zodx4wkq7LFWJTpZzwS8Tq1F3y
Pj132kUs0MDnzsHJW6togYKpa4dHcwiFeLBmb7o04azXifDCh7Ju8lRCaezvNOUDq2BfErfD32qy
/rwjqpS+kFgwJXE1XrRPdzmbhThXRA615I0icgjni1e5QC+dMKz6g1jfnGfYcMv9qcPg8xORtYM6
8Y1L9xAZ6QTELmLHzx07vriZLKSN4Cu5Ltk3WwSAdbl0OBiL1RZe2236UU1xBy9EBW6CoSNTWjHq
RF9e6QvB0DavzptP1yRlEo8sSe2i+SFgKXonwqW1W5Rf1hgciUAEDIptUMah+YZhuxZDBjl9OTkS
LQTbrFe0m905bsg7WuQ6NP6k9kCQf0zoCCU9bIcIkX8gmEekvUOLJ5wFnaE18BEeNGm74IcQquJb
Dqfs3Sl4f1CNnl9Hky8rCK/7NF0N9Woz6LlpNKHPm4jvpX26Mc6yphGJadKFnphoPN0KSvjLS9kz
l8Klfh4FFAXuKoDCQBiqp/8OCBiO2A/dJhuiKFPUvdDnQO7FAZcLctDwgl3iCrc8tbp3Gcip1zxY
gve8PVEIOhpTJF1Bh0B+TEyQcQSbT99FueBHzAk5SGCiidB7KhjH4e8peoh5Ik77v/Yy+a1ac8fj
i1OUWm0wWOQ5L4MVPpqYkfbA5uKPHrVBTJQgdLuQXefrjU8N5BafZZbL6VSrR5gsvcE4o/8z8vq0
TQLrRE2bALKldrpwTVxbVU6xfAhx06Wx0uen5JvbbshiXIgfIijCGN5wyRoAVOnZrjpCP/wPXAZ3
9MwfoAKknJbvxKRMjYToRXVakHRd8Mh58kgeqj4HpDVs2dwgrAX2Xl+1l1yzf84xiwycpqHjmIKi
I5WMJDTSRPe9a21Czc6ZEezuYH7jdQeA0IdueCyt75J89aOs8Pya3KbhOsvHiZ3/K0CSWDeVa3BG
FAojyKgnEY+pZg4aR9iXcvOcM3b/vXWd2kl3h3dx5Ak9jG+Lj/BPiiaagZca8uq5DQRnoY49sKm2
14MMkULNAc+V7oN9Fcjr8sFJjoL6q1X4xYK6yoaP05EbgZ8/qjXMfbyQTuCWozVirEnrbHopDMFd
ZqFLIeE8Dq3YiCF1nING74X8okrOvf/QeeWOrCRHWnNSVCn3p+70BLnw65dE5m/duUo1ckj4P7Gu
5sFZQgQCFJqTLVQSxzpofJZicG+ISaYh+QDenSr9eDPgAPhdgLOtY8hju+B4D+B75VemC0WWsozD
eaSOL/lN0l+p46qEFom+/E5WP//hng1oYNhX7wdaV3xjqV7zi2VNKRsPlCge4pfwZkk4rXwhDjI+
x+7DbUcrRzZCbO5IgL/jC+kQhHCDaI/3QgFGdvXDCOI+rTYlsZqdy+yJTBCN0KX+vIrcjxn9bQA5
ipC49oi8xYAcNT0KjmCZWpO2CqU5j1AAk4J1PLQ4Jw2pneDz/DFQIctxbf16q6fWT0y96MMsdHdb
1ZcZwB4RZD9MqCyToMQ5KG7R40gfp12hxe4IAAvyd2wz6iHRo4R33KyccuU9fSUFAEYJdgHpysUg
XUy1PuPbv4uhTBR6garnuBf+DO4eNJ9M+uQ22Wnts+aJEFx91hjke9w4b/nZqq723mggs9DzFLkV
rMeg1Md4pHEcBb1buUFSr+PHb7bFhqnkzdk6wder21QNag/+c0Cy8n26NAMaz5ebehrviTOg6ny4
WFAJOXTOO8/U80uaSwZWQi+NaBQfqsr3fkfLjvNqu1ODJqzJj1XOVfvB3lFGtYJsPFijmA2SKdKB
Gf+D5grlUq0e4nFMUjpHy9NiVNdGQWWiBObrEl3dCK9QGOfZ6lUmryRNLzINyWYj/cDSgcdnGpMk
Exh3e5tt+H4psLUVudnxN/WC0tdkjO3Ec1aRPsTFNsJLyQzi/XDywq950wCCj+k7QxpQsNCV3o3H
jMCA1ehh+955rOnfWK3kjz0QmDcNhWSe8/uDV148/LITGwN97F2wQkOnn65Nzj3616hXievWkfR4
PSoQaeTC5f5KHAw7h+0BACupPTid8pj9zCYJFHlAJmymLDBj/dDG+Db0QMHnFFivRvtblkehMDzT
RfSHzYU1WWP6HLnvJdhRk3CbXqBqsPjzttKLj6+yrVvZWGtkjmp+cp0hYpD39iEuRGwBZuaEQ5o+
rYwVGr2z2Q2frn9tBp/aHYOHCoOKvchjXDg0D8b/WdBhA+wE3XHaiQIxd9xuROdplE01ySgsalKy
EcKbOaXvfQ9ru97dhyWnEfge3MSTvJNbiXiUsXbvbnd8EWrWEU0yqEFjL6zhJojziIheXVyvuMng
KoqPWfduJ2IebtAJOpj6D+DniePT2U0qa+4cJK51leLBL7rqKk9G3a8v4chnI3ugdr7t+zoE8FMv
QinwuBy3uq8a6SIeL96dWwBtdMC3WZPZuBwQ7LWhUNBHymqyBw5PTO3hxrsXaxoCaXwVTo5rjUqP
EHE0Plx0SY1xneNJmFF6GSAD9aA7UupuHW1cb/vCQb/DVygxgkwcdnmA8bXGIcDxls1CmaLXH8/v
xe/oyEh5IFTMb4BMvt5xP68XM/ADtVJrSnHgX4hkSumgB4AKof/JMgJ4IEzQPT4NG0tR892KNKtp
784T8ghAAAH0DwSGxFQssOMRjN1VJkItLTiSx0y8Af37qoH525pMOcGeKrgX9ZhKcTyJ7AAytEwT
60bB0LIrb4rqzJTFWJjqTfPUQi6ixJVM2cOr3Id5XUw6F1VNWuY5NZuuMvWrqZFb96yOl9wIqsNB
g5aK6jBjFWXgrqym6y30pReNCI2BHLgUtDPgcVUtpYsAMVCv4ioPSUnbnZXrtpQDhZBdt7xUo7B+
HrkKsOLfBxZQsCOVKKZMaIhSn7QKouoV7sfv9RZG01G7x8ZK0T1HYSezPzQ58vaXY0BirIZknCKd
SdHGNuXN5u22uQYQnaIpiTA8fDXH1NeBQdZeRCSpKoEWYVNMpTPljq3lsa4UDrmPvA/KNJGJ7DcB
twjU2Hx526n38rjn15PFJDE+CU4vlBRgrW2JBZfNYqAA9IiK4iFYtSRwSXVLwf3GlRnMPFaqqcrJ
UdZmwzO5A4Y9M7NRVcPyVrapgoOMDoE5MHgwlkAz2XOp/U8Yog6kK4YugF2TnxkmomXLFd/nS5XQ
IF0e3dkL3bQjJ+5TA02wtbbUm6tgiDsHVEcDY97TLNJy/cLaFwTO4eK9k2R+Jw6otWQigUo5XYvv
tt/lNCxcWRQXuCQqSomwpPTfoR/nO5FwYs6iLaz0LyyPrq4FJJtpfzxcRFR4pIcZqOhOLevmD0Wg
kMSkV8TUZoz8PtW+8TPcN9R9matcCCF5UUOFeYWywzIhP9TbJJIjoOwNRaD71y6lNHGn8OQbfQsA
7GRJHypDdJxzkoxWNT20/kJoY7PrXUTlXnxcRfuIWNjPU6iITrKuUbeAQSTQrJ44eNtFtPW9/XKe
Q4dWnuPqnSWU6b6yX+lzZ4kgyicWBDHFSkTaGhzLQ/xvKOifmd3BIyHtnaeGvKfkYnbwmnuTBYRk
d8TfG2B7xh4aKKVCVZcryP6tKqlKM+KfHrjB/ddW6ht0B/cC+D49Dgz/aiube8xz5/Kdxe7hO2TP
rrNorYlHhFYnVzuowLpLujmjdJMjDNkE5jwL64phA+vWRuYcf5SHVu1lFiu5YurHvVnUntlVW6nw
AaB/REIvOsVwa+lL33nu2uLXs51EJLa//SjAsOQKomIL23Lw/e3Qajkx67xoM2quB19Sz685j/tw
L64QCD1qqGF/NSbLBclVjqfU6jAkGXEsBEKfmXbvf5JjYcIMFgk/HRX6NdWKEY70rWYGNl1zRbtN
2EwSlVwB3M2Sv1MBkpLfNhUt1y8xleQ23du9o6dmL7QxK6l3kvD4cH8O7TcIHpPl46iWAM1wLE51
5zlvfI9mBHzgFqokpdLdr/+sDTzolLydAJGlE/0jEf+sa5OgDSHzoiD0nc5x3X4TspdRCCcrW3u+
PekOO+k8JstuTKf0mzxRDjuHb9vkagdWIyISHE+YxldXy8aSrdpvIJdMHGaKF2+fxDpONjZUjnIn
6SoAXZA2R+s6eXhGZ6B6/ApwZqvy/hul5NUT3XzIMKVxdcH02IV7ffsmJ111/FzDrt0rMFOwIgKL
AJ3jqTaYL/VzB31JkhYeOrcsq3vKK0NcFs19SDklsELD8e29Ky84z1qXQMlxMD76FuoM8l3oBPwi
GnddvHepKp32KTigN1jTl5tb86d9Qp0DB4ZDP4/GpS+lvbPppDztFymHbEd3DYaSmiQG83uDdhiG
fkDrOFEMYZ9Jrl+bp2vQ7LTNxbKck1SQcxMzpcGln+oXIt+uar70Gy8qOuFWwAFwVJQVAO6MY0uu
sUSWlkV5jCo22WlvRSak7O3+W8Syum7MHOiKFpyGNK/WSHZzEzY4xqDDiVf19Vg4ffCxkENPt5sJ
KyIgbLu8jTvZgv6m+f/4EXqGjAiSTVnjWjItKatg7U3c/eOWyTOCs/9CrqtJOSdl05cPlFHurkBD
KEPpV6QMuP2nK+6c1Vebte4kXZTRtsR3/tR+KmzYQtULNbCwEcXzw1hiNhdzRkmdDZ/UjJoy/HcW
SEffsMp+DDuFfBZI3azz+NgGkCSm8zNng2QxcxZFBBrVaOFE3n/CGiOjjot/aNrUF6hQbQqiPLld
67ylAEZoGdW/EKSQIqorwrhRKQS7KaWhWxX2uVLN/wgo7Tpm9Z/Z1TYaoUAj9j/KVjRZ7tQYndj4
izkWmTu58mrKWSpOQ+mDmsyRq3LpL85I9D9pfyzCmZ+bgdqD+0WrDfpdziVSMDOR8bSNhJt3kro9
fryR5EeB8v9I7NTvpVA4XPmNRP3meiaTwkq3DI/sfDWuvs70kONOnbyda1LDb50rTX98esglnN82
XomolYXa34pPw5MuBWbZ4Dcon1NsyyxMz5LBSrhw7rT8ZsEZ5Sua4PHFmOZEuPkQ71GAHjPWlfT5
XwMW08/tfdpVNXNHZPZiXUbgi+EQYEu6L0d3AKfMmtJ+X/I/1L5raR3xxub5fdeUZuUO563xj2Sk
5gMC33j3YnMqPi4Cd6H1pKiGUE6QwLOU3VHtFTCGXk7+tkQDvn5kfAqoUCFyT5cG1uMbIqCh8eZN
MA+odivskY6FFzjlQKg+DtA91xXHS1avZBOWu7yMbUKo3wn/EPpz0u+VdVdIMcMrPmXjsZ4vNWrb
LPYsCq7HLeR+ufRnVoBst6hSQPBPAMKN7ZpGCZM2wxbvcg2mqVkok7QyC/8kYsFaseVYmOxK5KEe
+XKMBmKSGnaoFdQ+o56JKzE6+1/VMNmNxa0GEIObqFqLAF6vBiMJvdT7N8h06uSmieNfsuK10WEm
tDE69aA4qxbIASuLzEVECi7g5PfDPF1vt7CRotYfhaiNxd/xEZVdwreGBnE7l0wALy71tYxlAJeb
8NT8wX3DnKRfybDGVo2BiK0fqnnKP6utEIUqkz88TLtLb9uQyzTBll49QQbmMZpKSH6/Wr5BmebZ
5uu8+TPSwGYv/Pv8g4ihyvaNcfCY397lKCV8bmiWN4MzRKPHA+mevBAXxMqtMGJ7AeMGNfrm3Voi
k3qM9a8L1TNoaWGd/+BSYRKtukYFN68lgWewAWOx1ubKn2wOPnuCYClYdxCQc4YSTpT5d+T5XpOT
QI+EEirn3oAyyQi4ZhH48Qk+qnP4AkcXk9IWGS1CLHC3oD0g5NNTfADbZl6uhDbAQXYStfWBmR2v
h3YMdTWrpf7dSjYrWdiVGZ0bn3TCl0y1HuXqgCzEdsNiw+QQqIhTDvHF5FgwsfsH44c6S0Pph1AH
vCgA1twDikLMPIi5oMU+7OFomK+cBP3iBuFd6tgL70/fprg3e0Q/T8/NSV/a8XsnqZ0vqQSZjgxO
7YKD/DcPnH/ledNLqP4ikpw9FCIAAYbrVRcwW+58DDZCPx+wytT9ftfSLNL7ym6rAsS8vqIne/Iv
Yp/IUQGrXkUqoIBRTTWMuYs3rHor9y4WluYmot9brS1Hy46afHZ7DoG21e0uniOgKJBBlmxlmHLS
i9TjJO6TiXpaBE2U4EWAbbsnSwwX3HcEWLpJcwxxzuwb2lVVDzNPFcx0w9nd6jE0yaj/5pFFi2E8
+UZf4NyJA/igFmZ3+qdweRMVRqERIkZc28wcDuo2yLtr15Fkm7Dm49TSN4aXc3rHJzxYGT1OM/9R
VI0XdNVg05fQY1BOvmLhEKgG9yS0ac0KN/Gv4957X+tocmICspC+OTj3aZmIQjvAeg2uaWEpzz05
69BpYwjAkRXSQqXPMSFTuMAzZsy7fSX2w5g3ObtuD+EOeB+SW4gFUJ9PwIAX9BT5QpG/Usq8KWiW
edPcUk9kY9sDE6sdSr3AbAQGGX4EI2u/XGJkcJndW8QGkn2dQGjU8fkWKXME4BwKOgQT3siAxxGD
+hrqK2VJnN8statmJpz2AFWL0ZIcQFvL4/SF5W8xfQShoP5v8mD+Uk2mkxZditASzW7gWlUmKyQu
ZwqWxylJPNxcr1FilqVgWr7o36qlKZNCTqNxPhVohoeKB78Lye5QCrUP2HdhfcrVbUnivKj9Ug1C
yKIerkElCnc2PpNkaUBcUrye00ozXn53FtxvdNUWhvDxc4ORxgJ/zYSBfu0ejbwFCog939+z0jcR
o/RGMf+e8EhFEhO+ObQFjZ+134CbwBelFLIu92azP7GXF/LLZ798rqHi3fjPtCPDSZorkbhwka3R
jZYT10D5xTi541BWMRgtxZfgoeNl4Z4kk3ysk4ZJeVTX9peBBpGJ3Xz/nsFfuk2di2JAxmSxfcZB
YYtB95FyPkkZp63lfpKd/jPY7abGqQDX7H6a0vtLD8beN7yBT2xZuwIaI6HPU8YJtdZlbS4mS1hZ
2TFhSSuIMMIaI3mTm4etBG3DcSSjFPnnos91j618bklmdyKYTLa3X234ww2LDzQCCd7kNA8gARVf
Cf3joDr5fAPi6fXGXv5cAMO5zv+vfZCUgx5BKRAH1q2ybmt8sXgw62XOAwbg/WPSXOfmyKg8jtf0
D/n5O4vYNbGmUoFF3fEyG/Cii5v8PmtqcTgRDDwk23BH2k1U9xZJlpQ7dOOrq/fhJktfU2PP6cHb
6qf5M0fXCydhMstHmGgj4sjnLh/uGmXHnBVzrPckVR8/+OhNkXt6amP1TlJK9AjiB7FR12uyU0DI
uWC+P6gfnVsfDudm8gPUoLvFwX/R67ZjSu2EJlHagtf8zmPPR+KA79Nx3xHdhLRp1OORtEKPBVvy
PIrx20GoUmXVHaOmlgacBMiR7cJ2lpTdW3qBqjuppTDEAvi8SvI5enVxnejjTUM04IzNOltezU5f
YFpX3UdI7tPL7/9yyvI8G9v8SQ9jLTgTENAB2xUSS4sCExilgEGXca+uMTEwTK7NKUZ8vNLDLCP3
P2360Px/bDiL595DarfORmpxlixbI10+lY3+vB2Mqoi3zC/XGmGbzS+ZUh6uRGrkYcmn3V9LmVXj
ZUvHrrjeBgGl0K5WI309N+yHdz+EkTRWeEgklJSol0JjGntgGPkZlBuZNcIHzMA4cqTZTdRIQeri
fSvbf0eB0l03UuboDbFTfz1dFE/RJgtK8d6lapIcYZ1FS/CBvCptTIji/s4iMNohBmrAen9BVIWG
h5qCyAeNxOmB2drgSdCNdQ5eC6SBIqr6rlEfm0R6Sk9GyvLFQcS3HJU6h9HiRWC7jAlq4Kv6VfNw
+Lj7kJwEMLRywaOpa/PaWdv5BG98FsMyIaHgPvSgMlKvdvKcuEO/P7CN+Jm6AYB0qDR89DxU4GZo
i8JBZzWiOdcaHsdTjTU7eQexmf4SxwM5c19qqsSn2/Q6Mr1j4q3NIigUzv3UZ8i+8nMQ//Qm0mof
TP9jJgqgpn+mQmtP94OwC/y/cwHsxVOkv1Fg3J2ZLvQGnsACRJZO9HdWRtfQPhjH5r1nb40biVEW
e4p5NQbs66b+ADTAYEvLFQdag95miStsBq/FU0T4USmXi0SVpvT5bnEjyboZr+FgKkFyFFOiQ7U4
T94hgwS6GGzDpFAwg6mM7Omu2hnCoR2QKMAJbH3dxJ3n574V5cTiq31u4sRlhQTFsDYxIruKcQyZ
8F1vbZenMbFB/YTBCUaX37zMWx7HbrIpvpfORXBB/yWJipWgDU5lSaw2vybwoRcc8BM8o8jvj7Hb
fnF+jXAHOB/Sp8Iyhwe4YMoN4r+w9CIl6I1aPhjZOfSn/S6M3lmWQPEY8ZT00vVBD8ZI6UeMzSMM
p/g7R66WN6lHwp7sqFgPKdvgqVjy6ovVDx6gRh7+SrI2GLu9mRzqIhZcckntXskfulcI3mBEotIJ
Zsc58DcDAxCk5IvdTP4tf3OMoe4z5+buPxB3skoT/ZLxt3wQ+GnR2cFtV5Ru+5AmsWYZn4LcI0fQ
NabvpxIo/6aKQY3+0RYy2MCWXDMs8F1uTvGvouXCfvqMCviji6y5nD4nKZFSxFZQCb6s20fHFm4p
X/AEB9Ug4OmKU5X9wnxAOdpGECkSoPKWz5Uuda16EEbKHXEq+BDPKuC0Dh9D5BMlrxg/0JahRg2b
J2H2n17ZkiZiaMaSGvdh+GTlk3ueHdKC+NWD9S8bxRHLMRDWfkZQWg2NGPps10jnJ3SQb4zTijeY
zttJXMiw+/p+cLoimBVUANe+2OORh2Brc8mHGXbhFUsbotHptG3+OVGN131gnxN+SG0D7lGgFFze
oR4gISF3f81v4fDnKAjsxJUoEzvHAGYOPm3YjHSdQxnEG7JIwgeXWYk4h+YucKaG2dZgtqwgwa2D
eCR1o7EKVdgSm4uuK2IqQjdVg0v2NrfzQxkWDRJCK3GTgY9jdDpnuf5atzVaKSiNENf7ssoa5ysQ
tbIab5q6lcYQ+31bG3HI5Q95Zsac9MNTi6h3DIU/JXu1ukYUeSPTQlu+WSGBfBG2HI8STmBih7nM
YI1WXivsbB0lkiKg9q6ceESzRjtOa4to4IcsbDDeT4Fi/UtWO44PSzmB4SW1v6VbS6WCEtu8HJK2
Fo4rJ4MWfV4ofTbP/Os1EQRIOXIwjM8cFFRJIu5ZaVGaUhgzZefRPCHhNHltc6Pb3IzqamvWmxZi
o9nmKbp//rWxosFn24LXfgXjHn2Tzyw8ZQSlIrCITIh3eZmQ1itbkSlESlpP1OZgNkDAAwftmeQN
xZXKYPBHwGwy4ihSEQyw+OUQpSWUbTQON6f7YF/HwXwW/n9O4QHGB5hs5dXq3RLBtY2n+ueYjBNm
1ecGSIMJKzri1bjyboMVjleTY2o+FSk7/K08h8ss8CcmVfYC9zOnbz3DtwWUVm0HZPS+Uhttf4m/
JQcbqSgEBD4Qb01UAJldCcV2TrjCvEh7MRS8FBHmvwGKuVAySIAiyam+ke28/hiYkqtQ7MX8mKy2
652G80J0NBPwSVxU1PgWqaWRVFbPK6pUT87Ueh8S9mEJYz8OoZgdB7vOIuP1dghokVsFOya6aqDc
pNVRXs1Ei5Qz8wvbUS+lWX5YTZ4vRsvytdGE28CJfhTopSWWdniVxbUG3TieJs8nYnHMx9wv2ngB
gGptP33HC8AgI7op89j7o/SRuQahFcOCv+bvUEX4m65h6w/lteaKPw8wwnR8Ski+UaSbDm9bwLsQ
ek7sXYR3thAl4L/iEZCAAx7eltenbLxgV3ogj8/iHkHMo5aZWs65lHo4d8GjU0CKEvuFIUgPLQns
paaBhhNr+Y9JvsYZ8EvbLumo/qHIt/me1o4fM+41QpkPyHah4wKjC5oAi/CA66OSHz6QdEmDivpz
3rnHhijATV4DPrgNOTZoIV1lmxWzkImz7cOtWe9m2iS/fCHqw7sXsyjP5AZDKBj8SNRTzXNkaKDd
EOAfSgURaeIQ+6aihurmcUYnNW2OgYEnR6rVnl2OPNzNKek1WqCGUeDg0hvyAJKUSFRlpFHokuIV
ZF8zUtWco+aQmuJYe+8nBLb8LOo+zwZWgH1fq3cHQ9Micq4WRFWg5OK2Q+cRp9r+fRsYqDsL0ojV
pBxf2pfs2+eenV+4Y9fm84AsiyfR2n8D11krptpdSACadle1rTDDAmR/3BmVK9z4HD7JFqEZ/qNx
X3IL96PmAdwzr5uBR7WFrAHILGD8ffQEdUXqxoD2rrZHmzLAGo6Pba1epPsgJYUGqKSyXbDaxE69
jhSGXbQnK1Wy6wzwyHXntn8i8nrXgUTE6jdyg8dnPkL4V49Y8eoSDXksm7qurcC9NtL95j0RY9ro
CEGUqcALUy8kVAU7jaEHh67E4pO3L2cDFV7StQnk66YdjPKVH1vo2uCMZsVhT0Psm7xe5NhdCXwP
mo/8nFjVxurHd5wok1GNb9p5WjoVSfSz5WAWgyqr0vxQurnuCHaDpPhzESHUgzh0xKIRIHSkXVxF
ZC8DeGqVfoFNbi2IOyYOMSy3dtbDnoraDw4XozjAAo/yN7f5UP4cqyKYuy6nqxBrkQ7xlqrYcvr/
nnayBXJPD5lGe4EX8t12JRrZ05W9pxzT04IOQR0rw88gGls6KQi+S3QwBwEkBmqG4NVGAI1hA//Y
WqOQwNZrxEoVeBrkBdAtvTOYDGFO+2/i7t+khTxlJrnpmlsyFSOysw6PY3PR5ahcg4RiRyaDwI6K
v7YrTlE6mA7Wxl0JdPo/3f3k8nqUcm4xTsBeqHyzTRCobBzZXlkQRVYG9xCixxBCIpUpOoBwCts9
Emml8kz/v7fvRlTai4enFrhgxLyVnqKfdXYr9qL53yx26efK+Yz8tNho3qB28+l5va9I8UnVYyH8
n+Ub/8AXJIiw/kVwBerjFQA7wmJ1oE7VwdMiX5A7xaaG5JYxUVkZn4mfzwdTX05lKR8vhoHanIAM
VpD2h+aufkPYgPmHG5Kq6VECfQV/A739uYq89C4Pw5jirZvIJRFiX8q+5t+JQp8w27XDqXN3Uv/z
PZC5/51e9JPtDGd8ODAAVnJ/ke4mAonp1ZozEZ2kYFjL8dGAGLQ364B1zdWpZLDLW2bmoMOtuYqU
i1lzZgjwXNDYg5uo/lFiK9VtdOexm/9XdsDYqNVbFChMvmQRrjLdByJ8Uw36BBV1GMCGa1UMnQOc
cq1Pf9VwZoDWin5b879oAYv6sj1aBs39JLc3N1eXU8NSsKo49qXCe/5WqYhbFx6SYvIZGvLm4cBp
BCsZ9fo5yusfD3JenN3aJQ83EmabG7d9p3xgeDJNH4xlFl8G4hfwejkhhQonFrZhFlFJYGDJpQKC
4TR0JG9H8hrr5qoAPl1gqPWdR2OezT7XU9I+XGvz6PZDL6twv1s6p51THLiOhXZknd7/e7GISPvl
WhdTLmNZd/rP83/1/CJAl71oMcVDthI1lJDoEoE5fdlwwIKWlE26fAVQIMkA7Cn0UqTRtLGEjg6V
LEa3W1bGDsIFBtKkkZF/pg1nq2HkErjEmhN2q7d0IQ7okq+158oN/F0V6elWByfWUihfYPVqLWtt
Kkds8dohKDxA3uhos+ZQ4Fya/6B0IUDy1ZJhbaZ9nVMmOjkRB2Jh7EQHwb/9Di0TO9nVBdkW7Irj
2Jde9rzZXsWLEgtoAw6EKJaG6lCz9mBa7ssGDV+WgTm0ZzFFPK+GPLsnjL7WJBvJX4/vKAwIJ2pY
HQb/355OM6DMSIsmD/zasMgjhNof/OJ+pOlqJHhSR7vZ32ROWST2FxYICLjh7JL8nOrw7Idzj6HU
eKIIIoW5KBuXHTZhLKLmg/UnxNRZk6K7smNLp52An3cGcn5K+PvwqdgKDcotOyJgtl2wJzHFP85a
TAk2VGiWGGJAFWmhfItu/t9ZcAvqlcR2R3drWFDaEzxuHstlsk/Ft0Rq8q/deDmaWJ+Ok068NJYq
60KPG/vL0NZuv0n9xcLzc/D4MhGkSEjPeHMB/IJfCJFSVVz9nfh6DAEOOeELOLT+dmwMwoQz8LMA
Ic7vMDyJkV2XxG09sh0v8hGwgRxBJr+rIO3MLbBSrUcL59m98+QRb0aElv9xCi+gcLih/UoiTKWs
1UQ0DIL/bOOkGBfEOL9aPPsywkVmI0dU/0aB4sb1CvNYQjEPmzfAyjlcQ1snBb2qtmFm+QepjitY
HAb4HdY2VwLPLojrU2OTptJ6KxGAimYXU0j0Qkqsk306ffHQaUO6uN8xUqMyKREOJjGav2GGFd2a
zlb3dzrFhXtLJ7z4UZWas/2gxzWhFwy3GZqu3/D2q6ftP1qWvmRYCw7s1oGy+5Oj9fhAjeAk9Xu3
Pagp/v4b/OVMzWfLamffnuo8qg/RNZhVFjHeH4jZ6azJOgA8R1qMKGB6W/Ho6YmCFvjBYXQyXK4q
thNM2EI0MSR6KIisQ0qGPHLwFqOZ/wWjwdApVk3JD/ol14QGOggAYeI5FmMvfYpBVYE8gImSxKlQ
OwmoHsDDF1d93277kK+mkbPFQ6fm2J+QSQ5MHtkQZGZKVAgGogAo4XdtnnfY3Qj04xnf8eWMmHE0
EPhpS5Zp6Z5h4mUb6MQZm0TAqpcuQrFVBSVnByoP/C8K/gJcEeI+DvYO8VKkaMfLXVqseSABRJn3
xphhFs15YdB317LxXt12F/PU/YNmweeUToQEk2XqzkCEbgnCSRBzICCmgzW0XvJtFRL/WxhvQ8fH
yZWo7PtZNm5CQ/rzggYf8eaKUc/8A+hloAmRVdpJZ7kryehwTfcAg898WZ5zv1ABEDq9WcAyyH8b
Ll1ODeTeHs1/kyru6sD2cSs7IpP+T15VNUp0xvAbJ1BejHDEB/au3uR6jKxG5069JxMBTozZj2Kr
clFMB3Ihi0pCHNVxkRQ82VwY9NZ51Uj38K70bBJrPlm8lvogDJixWds5FuLObrzXv4nLBeGK1CNH
GJ4gz4AqTe/RvJDAjMWX1bVu9tHg+W/gMPwuBsyWXrE7OXrxak6AQ4Fyi7DSrc3hGFL1SbTuPxVs
OPp4epJ8R+x0wdnRlaYRIRHJBTAnJChSOgb4T3jjJEkUH8hA1k5xOju2/9e4SfZ17H8ifvzWt+gU
6I0/tQzzm+MUn0+inisepc8ZC/F84tpkYbIGPhD2AzQrtFiz9kt8EHv4zrOicbd+3OKAxAztPzOg
A7GEOgusdV1AIOCkyckfu2gM+Oxav5LL2RdLJnJDCFZoko9vpmAatfzSNbrWtTCoOp+MCQyH27IX
B322sFJIurU5ACv3yR4r2ElwQcy0ro4K7ZcShFj9rthx/MWmvOoPHjZzoR/i1Zqxw2gpPt9imcLk
sJpSQuSWiielJd3Mn5tcNpCdfl5MZpumEGY94735pmmtS59GT5WQF/uTUFVlet0pkY1s3B/Kk1DT
Pf6WhufGF236/2a19ulXFHNeD64DWwNtZ7kTJBDZKAEvrj9AC95KfLqgDPCbYeLFdCp7rrSEYNlt
8w6gKmURaQYBI9oSyDjfaLsTpfhlA08oxuqv/Rp39XcX6YNP8o6ChdGRHi/F5eu2/v6zZu72ZDcX
RHaH6O0cAR4/vl4HveP4qImrNq8dmJ0efSYgMks9pJxuUxkd10yT6voU4u0maWhPCNfj7SXvD3jj
nZL40NSi00DuIWQ5rGA80z52V/q2AG2p0hBKRGQWicVH5P99ZUJ77Bq1WLxOM3V5HDXL9LZvBBBw
yqPhHmlNuJRYegwMcuikJ7Ixj4W9+J2qbkhWXhtLZUAOXfsrAQS6VopKm2RRTcQymbvRDT1drd7w
92K86VlN+lpnKZevYMxb3GEAH3HgIVio0nI5KfuzRAnjZsgEz7J0N6Jsf7kE8Ig4ca+IMllJkXYi
I0rCwCaLIe3z7yCejiUt4OnVWcG99t5Qe2Opo2y1unR4iOk6nWf6hCDWEBzJg25XB1QG9uIQroJ2
cEraRVPxutZceskUtUY5DRAZpKSIIjOozij63e0RMs9TWfucHULgPlWAPN3cT59McnlvzUpy/Sy+
zExzpNGvFNsp+eH/knaM9Hsn7WJPUVlCRwjwsFlmJEGUe3+JGg+XoyRnIJsjV+3RvJzg3Pfbgb3X
zHbf1a006LE8q0Lxh983hoYRMV8McvVdi9MJWEighx6oqUhfBHsZ6ckBf5LfEm7kPqhfGvYAgEom
Y8NjOfWKX/QikxmEwidN4qqPervmIce+kjD5Bh4HitCXbw1NGeIq8rv76KxkjLFtJG6vmVFhzcmV
t6HF8u0Pru7MlXhtjOSLN2L6yXnN0QHCPkdCb59ooESDsFf7dEpVJX/NPUUj7ytNUwovE7NhtoLE
R7rDBxJ8piI8ExalX1fkDBJzvj+wOvMPQ66VJuSC+afBwUOPHQfidiFis+Q7eyGfsnhug0V0PZ1r
zX2RFXOy57mngtISvJxaiassQ4zBtA146YRcx8eo8tyhVnGn1Bwg3+TzCG1lCCi89oQ3hkJoCQAW
8a3zd5gEMW9lXaVGftYhwz1P042L2TjbrY/rWr1STwC+CX0vRGAcdUY0q7sR4VdHe8yUetB2VnCV
Cqqqj+XCzdcSoxSLiGKD3O7zovyJPl8osQ5w5hUsXu+xSntYIEMixUETxzvzZwiSfl5dG4YQiVqe
KGhFS147zw/lHuYb9H6/Oyn0aTXwH89CM0ndjL63wN7ULC7y5dcp+egzD28lsjQykENC8+q3XLqu
/t8LtJ0dWu4asLyOIOFxdtxjLuEt8yGNL1nXWPwZW+Ya74Sj193xZuqeCOC6D1Zxn8WUbOtrQJrx
Mf4aitHktc8V1QHKGpg0fq/HAS6KHQCnwCCSNDIvMqx/S3jQwE9bttDqH+DQh/h71RnkAB5F8aQx
qPt0RJQKoUz+wxN3VaoLumKZa/SNtq+2n1BRRRPh69dPbGxqj04lheL+o7lwFWSCa27m2hT/+5tr
NAJPA3ow0nEGgwhBSpDqSKcp2ncKQqjBxU7lgW/+muYW/mUR/ooUg80PmXDd13OfrMJrqoWB3GrM
UIqtoAzytOq/1Zt7uDdmYJJs64YZBwh2zVWn7z45ou34ZutdJYoukMTnYu8d6bp/Oqs18maszUMH
500gxy4+4tVzY9VeQrU2EIs6+LnwVB7Puma3i37X+RZL04rhTDkjf43ozwV4NYT1p6JjBIzeh6iB
L1KCJGg6dtF2ovAwenW50fB1ePFkJ4AmHF7xELgpPlvnHWGFJxMY9TRIqQcwks1K4nTl0s0HDPZ6
kTpZn6YInc00ZC5m88jIgPaLsdAuU9xvTQly48s6yAo2bTZTsU5OoSdbxwKN4EO7NKzE42aZJk9o
AfsmUB7tWQUBSC614+vR/Z2S+fsUikFmiOqWn9rkATD/lyDwT0IzuP54wnUCQmmLt+wPQ4WARR9u
2MD8oZUnBn6P9iNx79ZF+lmmeGpPMS6wSjv9+0hkZUbgs7AI0CWC3k0xfKv5ZwgDhdI156kntLAk
x912IlHaHEsXiDXzYH4zr9OVyvnLlK/laDYSQu65Rp1o20s6ZbZo982TpSNXnS/rXkARLy8ih5KD
qqlPHq4blqAeMX+y/qsZmzfw79RQO3TU+y4uUdHX9i4kWKm/nce8RMhXTW8ihysYceyfcSk4xcpw
G84QqyyQI/QNQZQAd5O5yat1lj3MJ4WaekCMwFSrxaAP1tnHHLeMhnpVMf2JvLbqFvOB6N2bZzxk
sn8ZBbSdBbQBymnbCECkvfERT/FQj6cAhnRpxkN9g7En04TndPNkztpUQE6xnhhjqUZssETC3NrL
AkfHKxiHtc5M72MSq564jTJSDG8pkyrhM6YGde5YJQZ2LFXCVaUtwuoV1xzu0Oi9o5p/dk7PoCgM
aJA49c+z4pyiAucWn93/DmbanhdBz4T/c9cIjkpjJqH7qzrtvrTE90sqqwqA9XvRFsdKmWpVIpiK
kYZ0vs9qwW1cxrFdP4PS9IcTLkbD8IzBBdDP9hczpkO5I2GZ2CuBblS/O/EvAYTttLEhZLQv+fcb
7TpSH8e81j9mM6i9qk35q1IElFkM+tfcx00LPBK1DQZdR6nqDgiSki6c0WjB4tpF19y3KLkpzByL
ZhWSZkNc2xWc1GCqL63bTI/DQGjc1sfGR1RqPxUuCwGhc5XZ4Rh1Jd5/GLpkMd5EHcwRDSH1Tyv9
LoCv7PTm21cq0rHcuUuWdIhfHyG0vFBp/XRrVaGx7pWgRIGdhULSM8SgNB5w8jXpQVJh3vBAOcBx
m+fAaZTPC8JHxo8ajfDzM4Lm9J/qG3iyvfTc9+hoHcg7uBwmAn9ZgvbJjZK3+N16dgLpvIhK9Tok
IkLDzjcHpILNR5A2U1338qvPiI8Jaa6mV31r4U8Ecq3f5kPEJkzse+HMyzd0/8svE3yjEwh3H8Do
UIT678+K/6gEKJEOt4MVbPAjihSfh47CR+Jd1Yj1mqQd1OpAZYwb4WCkBbd4DQqwvsM0FkLD5LlM
3rndTyGtnYPdkbF9hihlh8BYF/erZxhTwWAkpnysDvG3ZvXsyDpWcxgaWIOfysAQLD2Xae8aK4DY
JxMaGGxIvOgyeUeWsWcW8I0UZc9mkwW7oxhB06kmi+bQs0l0Ioitf4DNnS1bA45kxKzj8IWXKhUP
kLZFUtlaF3kRftIPgk4FODltso+D9s3lVOi1gXzC7VzO3+GeuERylHQGOq2/Jh0bzKshb15RURNt
q6l1Dz5XWyn/ZlIPg9x/JJvHGJg4rdemU+uwV5O/v589Gt+jh4KXmcg56snB2ihGpGm+loMqfBsw
nx2xN/z7VJcqR3DfBe7UyP3pTw7FqXFh/ywziXSkTn56V0CM5ER8MWohPgHjgFDH84q9b9SmEkk5
Zq9DuwFI8p6nmk824Zk0sJM9xmkLolxFZ4VSaQ/7FErQlB/W293nf9xlFDXuvzUz5G/kmhvFnxiP
gYqv2dW6nzNHaViBs8hl9deEL6T0eFbOuCGySbwoOMN7NVW3L/OCegmeDkPJZVITuLsqjnV6UNem
sjHuS5hFBszo/qAI/JKRPV0pWd/VjEiNTiQWTSVbFncXTBiMRJI/xfp5y5FxcyAxoC81fgBKJ134
k8CYTX/c1ugCQIJV7B6T3Xhs0o1m3S2+FzoFSpgV97oE5ZHl6le3DJ5UrrmNnmR7XxBLvxrMljBY
9iUhOGRhjG6uQXaDYjZMqlm3iXbN8kBTpB70x3lIpJJPokUD03/EWssFDuSRootJNFsRtcw2Cjo6
29yla5r4T/XAMwPyTxcU6ZHFLCG3EnXZLrQLZr825HrrytmPDldl9OLuTkcVApJSNIhCHjusJvtF
jK5F5EhJDVpsaUDG765MvsSzWNhDYU6nmeDkwBqt81XiccPvadHNfp0puH03HYJEcWEvk4ve5GBT
rJxTUCsTIzA8QpvQeJ5OgrmWcsAnTmROZ4iIWVRflVUObpyrz7trOlnFAn2TY9Vv6AoGZRysWkX1
pGf0627QmauNaGYFppyKct+Zy3l2fibGdSb0vKlfiyHA7GnMDQift845bvc2uG7GdUTOm7BbfgQ6
WLoqKeX1rDkc+X7t7oldUVRSHi24I4MBRbr9S+/dVOKy7fSOJnXWXjREnwdvp88KSaXQx8h54Dwa
tyT+ijHqD7lvuAQm9amq4VqM/4YwxwRXTkF3kZbyOXAZoxpYpZSCETHFS3OsF5JAjDScSCJGqWRO
+KjJCnKlwl6Qwkvyyi+IVES05nkKi2XAOx/lyAXDygBCPpemETVs/S93hU+M/2pBqwtOhvK1yNjX
payDA+pXnKYgktRaF0hLfm1YaJTLiSDYMjE9EIfo2J0veECt29FGcSKrQefSicBESMC2EihmrcYQ
WmUmzNKJbOISWTkP1mEhSAKOpRiiymbgY/H9xiZ3poAJIJFzbHVFFe+Ox6cPURmHdmg8nwiDce6B
zl/133hWi0119nZdGGwgdL2iH7dn4oGGp+Zsf17m4Kiwt9sEiXGIAjq/PHAbdipkm/SP8ZnpIrdf
cahV3KUzazFSWtdFnX5LrU1e28a+jCdtfb5XjGS0WZNYxRTitJo6nS4E1jeVh65uC8Ml61EHRRcB
uYt8dhTueWLlGYe7jzH9awPGN+kN3o57mqMgxDKNZzN7W1KHPiAuuzAoX33zjy0SfTQpQNAkZHrM
6yyRRUTSkIlYE2B+rrmWTH13trO4Y1BuI1Z1OcNvJfbHAigbKMmlsOTNO+duyd9YepmgJDxtaE6c
XHbUmWeB0taXbSPe06aWols=
`protect end_protected
