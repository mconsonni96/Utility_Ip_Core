`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
aErT4Nl6eMyd88FotghE8pKCFelYO/ACPLIJX7UnqFzPSBWRw6etiotVjyIN5qstkxFKfXZQ/Zb/
Shgd/3N7h81sfWWhvP/Yj3mIKwGo9XZPM3jyLGJ5WQbLbskHTbTqRTeE6TZms2bR0plJrc3X+I+D
Jqd03/FZLQmRN+xQPiAHpJf0ir3zEpRQ9h1Ph5c3YDE/nSFVspbTm55JTmd3TCXRt7jhefS0rsy3
YW9+n/M/aWEIxMzbNLVeutobAKMsVrfCW1gqaMvCBrQgZTAHEunRdV8QMpmi30y1ck3l9nTexqu/
I8lq1FQY+gwHBXKebdUM0qtfi70RZF+uqXfCzA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="JfxaKJEIAj9uYBELQRdCFPDJFEBuf7klNnbQWHPnaCU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20656)
`protect data_block
cobwTO6BFm9TQQuR3PfQVI0gCPjoVKkOLsKuEqImuEx04oqwtJLSxV9w9zCTXhIcSTojXbFJ1+ty
HuU+g+gQ4triVadWRoOSpvK3PgTi1TTt8ITpPcz3ovXIdhsdN5D6hzqRnuLlRVsCn30yYw379SLq
P+bqRttaSbdxDKgWK/qFTVJpffpyWw2jOMrsgq7DCLNP/hkqOd/chBhpEnU8PyhgbuYxh3VL75sr
Fr+n6whC6jioRd+ZUcO/rNOPJi7dX6fxVNRjvgLNx+S4CR3CsKVs10e9LVlgEsxpOQ/aG3KcSCOn
047EwATmBUa4sm3/0lwAylXgi7TQnFUTUaWPdXSruYh7kUefJxDfA7AEaQgrU3jQzfuiGf0t77H6
fSWXOr3iYPrIM/JiK03V8mx6X/AmMGfngd1CqPh+NRVJpdl0pxRvXTsku+gxN27IDJVOmKo0Xz5C
mU1JIhXEjgPnuVuHJibY7OOV4RL/+9f+yy+UtnDn01QFoi39F8l08D4QH/mSLCMk0uG4VdVtkLaE
TaSZsrHB2wdbALVRDA6UUXQKDv1/7tkGNi5voQj8IMqd74iFMpWsse8jFngcSQ0c2IFk/sYSsiRQ
aJVIklbwAgAwwza5gqvxD9bGznzFGzvuQvg7tRww36MqubauTjInRwgZ1GHrPWj0/e5+99wcozzL
D1lG0aQxEaDfIDJQWy2CzHwSJC6kZE2vxN/F2OM+vMx/CiSNarXE1V8uLEnt6lET0QB6hlTe98B6
hp2JaDRoq0xqNo6s+dk2tQT2hatg2YjUdw1bSvgoaf8uxSni1EJCgW40KKcoTNZS1wlkuNiY+/7c
lOH1+407TXTFUjU8ItRbkgasV6dOUPH1Il9VTcLYUTPWum+K5+gbxrm0++hpJ9Q0CZQHLfwC2FhI
OlGBumTFAwCr8bcIJYk6Zg93bfqsrb9Gs/KmqXwlXom9FuNSd39xX4/abKuQiAt+W4kyy0/Y14sZ
IqgwmpgIi+Xjvy1x1IRm7bUmvH2xDZKr8n89y++7BfnT5rlITP8ohC57zwkMaPnL8U5c+XFvpPo7
siym6WWRpMuy2Tzu+4grZ9DvjzWjvG9AHeCNd2JskHjuvlts9pPWpHtGgjzreQc6+te7mGKZN/QY
sCKd6iPnXH4KRx3za+aKDuQbxGyO72WEUVWAHZHaUUt5zSXELxuZ1gU4foyG8KUKljimw2QZ8M8H
T7XxUq29Fb2cCpWwY8MYwg+boJFuYSinjXGIfVl/NnbA0dDNWstvmnCqpWTWxEo72Lg8TETGq+Yi
2kSF44XriLbxKF38DOil4tntLS+HxbxbQ8h3QFQ8goS/reeGbGxoabbCgwKMTqTM0VoUbR2Ayilb
m6lG6liZo9MgCEX11V7G6JVSVA/1FLVgOldRJIeQsK2t6pgdRCMJCmKjxgcRIR7Fh1Wv+H7jFkyL
eE077m0DEA303YxU7KgQ0DJSW3UPUkY72hP1uhx8aXS3VaQKV5znYeOmL1BVgVKVauXSwA/rW47I
iWJMceaayfCl8fdbjyaW7V634rQWNK1TeI5QAUayWiwDfUFN+BdPbkgEizoRgYfXbUpXsnVnHWp5
umGLO7QC5IZyX0B944HM7YH0f1zql8cTI2ScLoVjphpnvT3TVOj/l9Vl31FJqzTCxVbKz6orrC+f
AxAeqzc6AmVUUpYF3obA6nAT2zyYMlEUbhzXDrqAHjvOf18SEoX1mSyJn4ahf5JhCcQnf4jRV6aT
NU5gk+7a0P+fTIP2rTvArOsJOaEyvZQrYViXhnIBLAEskWXgNyPQjnQNbMuuEJl90ODBgKyfQVCl
gmFnUAyY92wigHAf9wcWG01QGfbJ5/4r+QGBIh7D0/m640ljrIIxzQ8RY6b0nR2U8Uu07QqQoTQK
GTMfDA3/vUndymk39OGseoa4leYFTEORkiHp/ipD4guPLs0/Mbu7JHJ3mWfbDqaR0jjzGL/jsS/D
qOdYtYG9b4A7saH0vr3O3xIJXtaGSBVBFzhs2fjelyhHnwdTTuPuG2DZhB2E/tC5UIXur8AzGmzT
wKJPgYXSwL9LiMWtEJO/bBxRKx38TQlsKBR1iv7xM+Kopq7l1Qf8bVDnMCwMTOp1Fy8JghEXHMf9
XldMCDCMRjVCtJyzTdgsBmn5SOogMFjoBJ0tC62PRp7Nma4qeszS0pwODTDFkuSJjzZEHlveFOvO
vSd7pbVMVQyZejDnJlrj7NEJwoIzmU2kJBc1QyUOCyksxh+wwvod7i/w2ApqZy3+YjbaUW7kPCfV
eP7/qZ666IVnJ8OZpCeVqjAdILT92DYpgjvfayk+aJ2Ldg/KZeMwHaoTpDjUVpQAWQ3yWRKzV+p5
I+315HKPJxoAuEFDXU4ilXhfiX32Z2cqqbm7gY7RMLZHyCxiaDJqI1LAjieG5hNMRqhxe3K2H8NU
6Z2jbIY1Q1QJ0p7SA17MtcMf1Zt0v/TMAy4NX3tQ2BevnJ4EHCxWj37aVoaZwjqjGY2XzAolavIe
w40RSvfEr31wgnd5QFMF2Qjhx1Haon70Yx0KLKDhXWKeTMcvPI9qByXEHZc6NA0NFql9sr/yF3Uf
Qwcjw8oE6o3gOdn9QAktNaxiy34RRmbl7h0amnHj2oEJ3+1jJD/Sx5UZ+Lmz+r3CM12gDJ8JLx23
vd/yihgIFBXWdw/mT6Dlc4fZ+A3VCZ8Et/9FXU1W4UnxDy8MuK81zq4Ieg9zm/Qtn9psJFDF7EsH
j5o+pG3sIIPZHSOY+IJl+GRN5xBdNnZnQ0Tu/82fF3PxDiiP4RRBZtyeHycNp9WijKRBKb5IAZob
pEE/fj46vVo6jBAA3GkpjUpz+Ww03wJWLb2SjhQrkQnC6CYO5fr/T8wOy66Oe3MFFFQR0+FG1LUr
l7CvuFqcVoYI/Q7fXgFP/snhkLstAsoXbDt56C8M85KcHo05qjq6+Nw02ORSI8KyFmwGUQ84W28H
SECIxj5ArbK4caCrxo44HvmIG2A6EZ5P51hN8ZV8Slv3F8xPag67Z1ZtxzqaPcZXE4vQY+9HSmL1
Alw6dW3M65sH0nxdbf+diwXWC/MlhgUGnVr9yK/MJVdZpB0UG9/ueBE9re08zuALYIRkC0xtXtn2
HonSfwd1Ad607XD18aAs0zfscFZqjPmLZ3ZMq5RnpxJRMPzamCH0hIoUpmQaYSrdfZjV6kiaw2OH
e6sXplAg1BHXsN4oq6spDTYGTgvl8xqrKxQ0z2ErOf2cCiSIAIsX4p2uFdsHB9+9e3mMkA07gMhV
pbxJrDXvrNy663UnxcMdTism2w3ynYIiUECVB0V27KXrR+apldPw+BmdPn2krZKFvfV2owSMLCRk
+7IoBTS5wPMTsldPZEJ3hOmL7jwBFvcQyBbyUrXO2riOLrOhue0XmgELFjs4B10Er7lHtnsdchcz
bgqrsH1fwZSQrZ3ZoXqvg34q9tmVY97+vLpuUItuaVSwqWwtKQF7BuCr30uIWzXU4CMRWL5998k0
1B8GqmTe4AkT/cFLF4goSts4pCQf5MKVcOiSL2LW7hXvu7U59B7REUHNpHY1UI7z8cdTdDV/BTbn
SOx8ZPjczeW72PnO8c6Qh1JJiX7HA1gqvvksCSnvqLedUji3+2uspyb7ih70KjJUowwsqYuggS8z
NMBxOa93NbsjlkF223J8gxjpHffoy23RBGIXwBo3S/Ci8u+Ep2BE77cWUov1JXq4Q9snNCmel1qX
+PO9Uotla3LJgnIwPw8TFpp35bg9ol58JkN6vPOwR64UsnB+jIgx1rcG9Y9Y+45WwUPO+v/05Cu9
N9N5iCWoF3uHFqZcrzf7uI4pS9KqG/w/s3jJVALhuFpcj0AMQsrCcYxPmSlNnWyebYcTRXeHcBNG
ip/wcroxD3e1U5gcte1iaCI0BEh4zGRHZOtXZ+I+pDghgSso4qqtr6Q4/xm0KwLmC77rnOpDS/2y
5+d8BXT7yX2P6U5FVYj+FU+U1yLpzZai+FcDtFE2gW7ih286X8S4MtiUHOE0ZCVsmj80j6IVFbuY
xGs49epDh4YZClnjTvGhUGAcoeU1m7I/0CxiSMQnEiAuQP1Sdj2HCPZbqrQhC2RHVknrKMFocrcU
xP1wLM9mrGcRBMurH3M90JFK/1ZQZbY3G2rXdOGFsT53pAhShW53C8k2vK9BF5mFxKl7vY3zEjIQ
hghi29BVhUzJl7P6tvjZAqt3FlzALOnHHPP78yKhBcFz3cv22xgDYy3LHdZkh64hID0NSgk5V4XC
zVGTQ0yXvLzbAVPs4QCC2PKLZVyRgHhJ1tHjHbMfBboxHE+oYRC+Wtjp+1qaMUYxRNzN7TjyoV69
7UvGWUfU73N5X0cD6p3GUkb+C9aRWuC6zqPoPG0AigfJDLvK4zJzPG5zzdF+JteyggoNXrshijVF
rF9sUifANFKtm859a7EeZ5hvCyv+xrNXFGPGj0k7lWy8LF+rQUrzCxRF1am6PRyE4sjdc6TZqbLp
qEJhZ57JhJwt8O+m8pOKlTp07CccNQtGXCMLAGk2k5bC2Gzd+1bk8Jx0Gw4YjjJYzQixsgvPL/fO
tPT1TS0v124i0Pk19GDjoGC1S7dpVMexcgnzGmsqMpYjilCznwVkEukrlvddGRgOwVj+F/ptqkmu
/6UrNKC5xhuEbgBNSUKt4VAqBAm3ZA/bh6FpOMRIG5klGD408giTirpk9Do2S7ab4J1ogIQg9mE7
Yenc5QzlbiUqrFZJJFaygnSzZSomvRhTzcLdy4X9GILJn2WtljyKbb97j3J8Pe65fRC786k3hXMO
6n6Xw6ckzuIHWmIbYBQIjpALwDgYlaXf1ZnWH5vp/dteZXh7h1a3Ptog1I4s06wzw04cMNHG+Dls
KR9Jq0CXyF1oMNLr09hGOJSr9qT9Z63PWDm4rLz8mdclUhFEKjmc+s3OdhlzeHr64KXSQc9u3jT4
Oyrp94HPOpncIgObf2rCF6+dI0mb2x4xBm6CbUSMhgFL1W5qERDUuW0UFUkw/Gb0kp+V9Rx+sJg8
zubq+Lr531Pij0NNh414qAb96XIL4n/ZGNysCtrYUPeHx8yYlMkXZmoibSgd01xcKoFsoRrk1sp5
FvUdQeRochzWnqlcmYKD/fUPuaJzcIFYu7LGNZZlu4XW+jfW75BmuEsveAZIuekXWTNKTI73l4To
pzzDJ0EJobedv1j7hrQOUrYMF87IHDAcI6ZdQkEicFi9CS2jPHCtvtVm6wya1l4nAmOZKM5APtca
JrLIIjQ8CWssu1cNTZ6mLHqD4dWoUSWxhFnQlGca3E5IIBZHk49CeeThvsgk9SutOgOHKpOPHEF1
GGqNbNsynOdKpqMvsDKblOxr8mpB6FmQJkz/iLKdyzSAAhOah88RZkiXwsPtZBZYLmaHD8mzUUuf
8IK72NJIsirf3+r8GEWKaVzR0St08NKVyhS0GJAcrI8Sx/vJ/VxRp5Gi4hLrUMgJ3dNtkTQRcugs
GyA/uV2Ar0bwTLMHPOkfV3US7A5hYeG7jHHpSPUTr3T0aj8ARIlCgpsGPG6iBhWj2Gd0I2mDkNbv
fJMiG0GHc09WN+QgwVECrr54Z8xFk4QkzdN22wmVnjKGSI1fJ6fXgY9dAEgkDU4aF5JXTFd2PG2s
Mcgg0OgBcunwq8tmu/H9Hho3Ryi6N4g+9RE7v7124D7+yQmJ3UlOeg0Jg0Sj82zKsBZ5oCtSdSY6
F41DI/eS7Q3vHTuq88Y2j1tA6vCE/zFEyoJ8HGfUpskh7FUaORXN80j1WEsKajkgM4o2HJY9Gu2R
cvkQtHuD84F9x5vpV728XV/EsPP0B/kmYotjWMXvBchaM9/Rh9OYQzE9TGx+O+zed0rUs1SOgmKQ
SvLqEbVSF5hr8iZTQDqzaxZlgBWklAs5HPIDLULHqpXz0qpR5WiPQlm1MnHbJ9RobuxDNLuU9XFK
DaOLQiYT3JjpioanrvNuNjtW85mAHIjm0oHZdiWge2kkgUHvLWi9UtLSa9XPfoKnn9TFz7e30bDb
2tnGhE4cGjhY0fQDet+MMUzQ3irQy8BsAey3V9oFEVvUR2jhRFyW42oxbGqWMohuiE9vIp0C9VWj
Aa4hCLZgnPODbggHXMnf62JpjEYUJRj2tjJ1N5DvvwgZ7C/kJ5ZOI7DiFas9iPVavVxt3K4qnVw4
G8C0CWSqic6GHov5f6FVZ5aKf4+dbkw0te3gblBXE0C1HrpQUJJBbDd0Z03O+auwFQBHvRvc6gY5
m/EJJWl7HHmhmusJj0VW6HrSmskwJe+yn2N0yDPD1opNztGFp2SRLRnvWmlvr7wPulusRfIjcd6Y
2o9F1MUEHHmVW6gehNwOET4Nu9tBNi4uEOewaC8r7aiJ++vhyr/LnkXQHF7lOtGyruAqKWo2MJ8M
T03l4hb4Ke+R+yY9A9goglljFbD2R3Q4d5jZCJvQdrE9yVnxA5bkGNXMLiifTvNqv95rOtD822Sq
zCncWQuR1bGFbAVt87hpGsBtp2g4UdJG2ST4F5o7eipkS7v60YFzu8LtkZVBfCRc30IJQ19ZnQkO
c+Z7WABrz+AbwxNRuDHT/bXcUStb+OMVncRDzAiTLQuEwji+p+uGgmng0kk6rQ44pazm318Llewc
HCTCIAPYc6MWbaUihcqa84h3L1qE8iFXSdTlu7+kMSJxfobZZoGcx6F8M20DmL74H4vnfF0TyvuX
kFduubIk/KydndR9TIJCaE+AKzpH0DYopO9A21JTN6TCVNE+wTVvQBdP6KXZPazD9G/06sqc5nZk
Tj0S73c526fX3qtkYw+7X4l3BoRMJVGXhMAf1NJ+zZfK3qSfJtVjlsuVfyLyjdVhHHVqNB+kprPL
1f4TsPm2U2Zujybpgjzwdwr10wMDUV2P8Oxd2dKixmcEaQF6PJS84KD0zqXOfdY3gOJ0ynAvVqmf
HPQeVcS+4usTuCkNrO6JTSwWri4nh9NHd4s3plwTzbI6bon4E19y3jiGiRYUWEoMJc2nsJPudl/v
bCbJQkoMKB+mFWASRT6Ud1X1wb2ynTSx0I2sz5xSXdXJVfaF7xTBT0l5aJ1Q3gTPZO1g4gtJR2Gd
jC0EU/Q0+9/SXUKRHa+DfbvFXr35Si21iaKg6Cto9kH2JTXz3Ks6vR7JURu2JwpHj1tW7Dxn5Nk9
5ZJidj6LKZiCg9xWc7b2EdV2huyh86gV05F4cNWO7+rDKCPH0DZOjitKOINcOGvEB+SwpnH+zx0y
/VX4vHLIEyIzsY7UqVb28pqYUDnIVdGJB5aO/Bi0SRJI/ZiCtJP7pE8Ji8euV8vpmEppGNYmasDk
MpMXaPE5UoIUAZQ9AR78/CaimPrWcVR9dM08/28u9BGqCkkI7vSmjdiHbemZlFmR45i4JdmTrEJJ
rIjaJG5ZSyIJ/EXNcO4SZbVblGv6u6+tve9BJAYx0mpWJVh9L3kLFL/G2VtR8ctKdvSWk6Sj1W0L
fuhDOenEu5CT3p87CmnuPQnfCT4EEwklsc4PtLglaZrYsC4kdHVh7+wwJvntoFk4NdlJ5a0YLKrG
PkC/3isA5iiOmmUSrkxy9yNhPNjCHPHDUxyB6nNvVkKvlDXWN0UiAsXufEqeI23dpU82ZE1ahA7/
61IVkqLyeOUsoRuu+S/okBegflq1Ffo7chOn/0rZVol16QllmnOvLl7VV1JMLFr8MEQMsaixe5r0
2NTvl+8Z55qpwwJCm0pbvvSzQdotXf9sjxyAj1d3tIRAYLTW1WXFSzJakNL5AlQ3kMl90ghGz1uH
7EDQw0PVVIEeG5J8MZAEA8axj3ee9I2wJX7G0yIIYGymqLO5AVwOiiAx98O5d4nzhbyqAyMKu6rS
S8cr2u09BKvqHFF71XcblWiNnlyGiABbjO6mE/WNhHcPfCnjk7KcYJELkmx5/H037CpzldY2K2UF
fF7iSN/CqVWJMIraiTWHfPj3ug9Om1TnZ/idtmrlOM1NFULcCljXvL6z+PQXXZmBoozqFaCpkPs3
c1lwevqZOD2f8/t3VgNgFuaMftmrZkpvbkq8NDdBTp6DbuuCijbrIX+kT4vSH++HCgVFZYUJ5YBo
knI6c6i1zDLGEqP/x1f4eSXm4T5bq1tkM+aW+ONcEa70I6vMDsfyDcQ8znTiKWWzHUKWwAHih2Z9
dzjPbnHZFw0ze6PvmQoCG693V5r1Xz9c7T0sW4dDpMqLcUkm7DnlbJbfmbArzG94qpKgWZs4llN8
FCiVTmEat/SzVx4JrXmwnJlvVy0u5y53WlNDMQOkErgyzpu18GaZ4ZFoJbU3ox0r340y0hunEBl8
2zv3T/tUQsXT8dOcR8FvgKKwLQ/8uVCxjGjnk4cHxTySkryo5vmBKCpt1K7lWKJ+wWOgFyOhPsh9
S7Akj9Uj5Pc/7WU9P26WXAfHpt4EKiu+74HCcrNZOj2nRcu8gJYS0vl/EaIyA9QbZJrMY+CMRDCw
SI4kJXLX+LWn3X57kvpHFHBMdNJDJeoItmvY6zctD69dvkBB4/9qHMGFF0PbTY5H6QTlXYigUvi3
P8UMyk4iNbXACCHn67yCdfgg2T9Zo55jGhgDbrV1TlG2llQT5wlITMfwVx5AQ/PUJjZnNs6dWqMz
3JSoPdKczvN47MIZRyrxQxi1JHW1CHnqIy7OjNQifJ6PaxXAjTsUxA2HUxG/0zvh1srrE/adhk7P
gy17/O+femG7Wb8C0TnSThYQiLvaSRZrMkcpjx3/JFPBICC15zSq9pU94IPOH8iInxGOrdixZeg/
lYJgZKDM7D+anedMNCp4Mz1uzxk7PkHFPsheUWiq5itYp1HJiNQFMsL9q+nx4WrHqD/3s9TE2wEi
TjdCsHqgAAlnYyynytk91d8Jk+b/Mp/ABzmxDJT8jNorBf6KiALtmD1DMp1rynKfTtLrJS7mp45y
UbksOFr8i2L94+aJGj6MDuDoffr3XRSXFIHi8dH1ECqJyXqmqdACkuWE037fYeP1cMrc3XykPnUb
QAiVRV1lggHJH22P02CJR1DJbgxb4ij9OMJp0ChfGwN2desjZcmlL5EBRVoKYbiW1mDcH+pBh7dd
LhsqwKPMPzfjeBEbAD+UVV+KhVGK+MlFLO3gNfQwGyfIJniSamH8pcbH8VX1/fsE1uDJcXd7YZdO
0VI+pzz8Nv4w28kUCBuD1TryNagPO2VIL6kjRpbRiB/fcxmOHgNEBW0S7UnLIkkMs/KkRQLXarW6
kRJ4BSpoSLxugpSgtRWf6LnWgMVb6FJrfC7PhF7mqIIZYWtj4jM9NP7xfmUIM4RNvEuKILH7lqvD
Y69lVIZkbEBe1JYQhvKrX+Mr7OYx9/cBGjjKGVSMbxxnmTiSRzbGAVmtNnq0bdLddH5DjGALRouq
KZhrXkZaiTo0/YKN2CF09G3Sfd5sfZSDOMImrsZ1Bpqx7cLCAVZNpZikxqh1hY4NlqdIyrLEU5dr
UxobMDCHHzJ6vOpiGITrCnoZHuUJg1LffXaNi1JGxFotc5C3z9Qr8Si9XSz8TF90Th0uGEUH4bgX
9ULI0pOH6Gll/cZk4FnBAkU2wqKhjGjTc6GCilaG2EhnJQlG20h1Wl04gTkOIu8vnp/VP2iZu7AY
1xLJ98/Szs62aElINSf8CErh0kUcX6u3oMnmMHt+woQ+QoB2dmCjY33OcGAWNgsKHsRAbr8lT4Sw
5g+KMZehVZDFyMe++VW0NQ/mrNpwJf/gb+EDyZQrs86oRO3b9mHyCVLKoyNWKIDq0tphV272WV82
WVAy80AfxyWRJsyivswEAcKedrTB06Sxp5lzmS2+b5iE9LdNjDE27PMGH5ZnMcKzJIkODIfpF/vJ
O7H72hmbbzum5Ax+jaSxauSngDrgZVY025avToLqvGuxjXK+W9/a8rP1YTYjL7FA1SisjUm5Dnn/
MyKtH0XeEDcwbmHHCqfKAVQX+nBQ8AMuQy2oFAOlAsZOR1bGxlkPluGDYsuWS1QtM2LB4cNeU2F+
GgAbYQJzPG1Jh1P6PCzx5KSZm2vaOqxyP4x+/qJdNR+fabSAsl8/vPX7RCyX02nDRlyafxI2YXr/
EKOqBwIc0FseIHacEwm/srLTI6f4BvVdCCVI/yC299PRXr0esgCiSiuRF9y5m6jLCZXqF1TClLz0
Tn8hqAjHYMCNfxnUfiBc7Oc/H+oPZ0PRgJpLaZi4Wt6d1WCTr+xHzYVygo0aCpmMOLpB7dHSGTYH
pSFO2B2VPWTUOWtFiwcpg+775rM8ArAv47WTwii602VZPzNJow+bP2WdsqStVjNuZLBHjgS/J+FI
mXOVr+tujnlbnZhG0c+HyIoM7HWbPcI0vHQ5BYym2L1bCbM46LIYe5AjWkAHP9WrhxQqKQNXLidU
Jyo6byF2xfpcyDXPzNPAdOAlN966hUq/hap4eFDQJgOrWGCvfctYyPfzV4svQcWqSqhFZFWkXcnM
QI/OIY+LL4rAq8ycI+aIS8Wyj4J0em1uFH69RpY7pTH18zBZzjTFJw0aYlEv95AQkdo+eVXNTMFu
CTGvjFVpGN6V3IRjBWEuH6AKSC2QqqdSqJXP1t8s5fUtxpvHhKLUg6BRk9vjJJxvBFkNffcIS0cr
erSRMYTG57GdoZ/kSOvSpYYoMyLb6x37L7Ltjs4UvAM2ctyJ2ArG+n7t2dksVMLyRBA23SlBYdxh
KIf1k3fbUyZvL7ylI3flJPBf9lVCnqc5Gvh8axb/2kOzbNs3ZrE9T5uVt0t2170mGFcaoTbwED4F
TNuWRLxpDS2UFB6z6aNfAktJPWnRg4yCWnOFZvcAykflGfKAZ0hOyT4FTv0HvtUbX+jOKfdOon3H
Zw+GgIsnSpGtjVlzgcLOKK53Cya2Xsi4jRUv+4E6g6Ws6DHGhRQa3BV6XFH/rdhYktMjEOgieQyi
stLaMDALX0fcYxnp6jxWSNRQLGug3M5ttmfKjkticCDxEPMkqE6GE9rLAjH3O2T3V/8vh8S4O0q+
oajOSbwRYhrytIrbIianw8XVVXbK5NLoRZC+fSCmDPlD2NeUMsc4j15RyGnQcrmUkrLj1NZepzy3
HhN8PB7tcKwuc5zE9cHxnoqPLBVyGTLoXD983J4dStk2KOrA9mQtI3EAubUh5k4Or+dXwUIVfgtF
rFd7t4VSO/rGwMWpt7CuxVUUiquueOB5HjZhb04pG9B9RSHS1IYGBVAoGZJXkShroUyO3Gk4EPjy
zcCG7M0X/aeoRlkDlxV7oTrDkaBvHs9+gAlVhy6pbZjEH4ssvIgfL6magfM6JP9R9K4nKG/XQrKh
eSfEHM0g+QCCMBJQW4Mi4VooKmcKH4PlwkZ83puUhZmeIqDi6Mxv7CJI9pD5dtkHHpbYdGqMWRMH
PxFUgDulQh5+cxpHIq+vTBDJQqUuixtuFFjynvNRiLHTTb9NvkYSySwm67zfUJlzINYtWTmdYfc1
oejVPNBhphMTKnXh9LlmYkNVKKjCNoHGWEnxs/UxJeiJ9Z4xyS2I7FOixcr74OBTJ35K8VrIKtUS
+GtwvKx95qzPeYMRgcNjjFylaGPAzkdZNXdrKkLrpzYU1QKmRM5zGIHLmoz9yy/WBXZTqPkfKrpa
Qr4BQTaFVwrvHTcCSNJm+QOlpXnIFqb3Jt512XbghCPdLyniKT5/PIeucPFggZxU8jruIj1KOHCN
O9PsM/ZDvcHsIFnEdrwWfvKuCHrmFcqUhTNlSv+ltzgrnKa6b3yXtfJp0SpXT43UbReAPDE3+R61
hyywNjTRrOG65hSjoGOggtOadyyDeHQ42M/HD+J8x8pHciDEtBe90FuZZSFjC1Mg8X7exWg9M7kk
kNlliB0273ealWptmAhjC8u6rx6jZY5Y1Qk0U27NAd/MNwJTobs1/ZJQ10WjcCRt9t23OuaqWrkK
g12XQVTZzd6GEGpDqSCiJE3dN17UOiNj02h7xlf8R3XWXXN4wz7iwDrY1hHfPDmD/P4DugcT5mwl
hfWij3+5p4rkqUTTwsUqfHXBQq0b3ehHiMl+SR6Di56fQT/r22kQt7UPTzX/lzmo2Y70MCJRzvuo
I/gb9WrmSXzxedWef923NF8VutOja1rNf1jqBvq8SZNIUylgnP7FlabNvF4nBOXu5gY+7RLUObUy
9eaptlsf2cIEUdpnwDPxi7spdFKX8L5ODjSR7It/xcvXOPhAitpqGsLu3THI6quneNyIvTpv/1Ry
7CHgBeV1NHttV7QzIQ1B4XhGUB5HlQ/VsIl5PJMnSHcWd518qPmS6ulAaRJVXWBwc8F9YcF5BvZg
PMe6DzTWePa4cSTF9Xq05puVDlGMt/dIAzLdvSuR3PfItXxo8k9iaPOigZNdUAxGWF/2Iafq/piu
iqN4EcMlKB+Cgr6bRKkRyWaFs8Pt6Oo99JRpJyx/T1MSAJ6M1+T40rA+vgRgcl8tvS5U68a/V7o0
nDNrcrA6Wb7REBTpQL9RnShslEPI+CcnSHZ+F2alzSY5CDFnd5DEEacqwKBHILIF/BTK55+pO18l
kJBReGqxiVZUSEd4VxlNMdVKpnKoLJOVjImg3WebUSY+LhFUdztrk4MekkY7hQDf49QyA5CnEFRi
yABl9yxFK28GQYV152c7CL/Ze3liwkPNxvYln3wCeNtDWlcPYOCD+0zWHQLfuljiRR6i4AMJIZF0
oHMBZ2vL9PLQKl3U/6MZ9ezb/asxTeK5HK/2r8abBvEYeLl+LjUM+Ue4TP2467tKlMXDRMNb3E/8
ArLpV8wqkKq8MscYkcmzPUK5z/wAjJ288m5GQAJfF/ZxiAAqM4c4EEdUyxWpmEKQQKeQq2vaQzeE
Geq7cOYl7CAGHm+KxJSpF0W8D/ycJvaxtBAfzE4VzSPzoFC4phgnflDozXsBS0dbOsNTI+DCcuhJ
hImvjRnI1b3GMtyJd/AYq2EPA0KUyX43g0fL7tcSINH4wZXoNJV+YFpxhfD4E+Envjaq7BXVRVaH
5aelD4E13KDJF3jNE593Pv8wSQB32C7skOtOIGvH/UEDqonF4nMq97TIW4NMwVXeKAIALkeRSNdo
nyvEMRLZ9q0fm4ijYamYAFdL9k7mA1sn6ebo65QbXRLxRd87D9ddmC11rh4NWW8KYVIl82gAwPfJ
OrViCSny22IPdKa8dlYwQxrigw610ZaJ+pPfqCfDfekco3pTjJy5EM/DsKK0umTRAcjJl4xhSKYC
Xn74AgzxLO/QsZtoJkLmXuifiLrvKF5ai2W36sDEpJB7XrilmF3M4upjg7WbVB1Uii9DDgoieTgU
3EJnmRfnO2gHG+H6hYCz38hpMbexZX4sTtM7xBaHguzE4e53BgW+G3cy4EuTrqxMY+RgikdXZAXd
srG83t71F0IIyCRTfQgCDt3XzjSXkZ3E581RiExUtLNgS9WzFCzLUnSOQUaDz/NupyglaLRgjZNg
n+xiUYqELTFz0ryXIn3oVN0rK0IiJPmY8OyAkdRBgmlJb7iulMBtVjCg+AljdzUefNXUmX7RWgGZ
p5CjyHq2SGPEUJ4tibn2qkLXaug5r7Uh0JdiDTcX0QoNRvoy326/1H2/WQfJOvntbLwCeaWsIthD
s0ArzQuKGrQbuJCJKUK24xvOd8TQSQy0UQHgY4Ex9EpN685MRg3P/My1zCndWAJEtqjWqQvSw7Gb
VcpJ14BiQv8N1m9KAornecpn0cq9brntzlNt6sLwAntxOY5cQSv3bluoNZL4u1pCagDQsrTlDn27
ARhpCZM0SJuY4t95zpSYqEraIPBv/ePwPF2qUTAf4kCwPS/RARZuRN+kQGzlw1mC5eJ9iARoWVf5
kqQJ3gDwBx0ii0gYfYj2T7LtvdhunxgokBzuDyT0KlOKhuDDA5518p3IHwc/yjCEolfp5yegKF3e
HYe76wq+loeTWYbQw5eB3QIXHE8q+ZkZQG2BBqfZw2/ZCT/OFjt2ltqGMhf/QVzckMj+IwyKDFiz
ejUKdsuxoB7Ns9SWYLkdXB7I5zPxo0l41ZK5VvyD3OPtunT3mxp13jQHcRhbPFoxAq2FnlJnLDXV
okDE7EfBD+nUog7WIMKrg80d3A8bgfMFuraT7bejfyYFi5/0+Q3mdjGKbeZcQGNr0yBysugGFZGR
uIulUMqHWjav9ie41LjtDWs50kb7MC47nekWQiU655ObsJm7zZHCshebm9sd4DF4IuAOH5a2jR+i
oECW1KTQ9bjxM9Hc5lXeqCwWq41xr9+mpN/CzLvkmZA/uHTS+r1oLHLiEI+sSWq7A1CV8h3NAbTZ
YS10tn/z8O1raDBSlJNjG2KbPbOkrKvKuGcwKiLAxakYs2raz0r27ZUjZLTk7XXqw1LHjuxANaD3
bJYl/E+DMu+Y8qD/qikISaX1HxHNYVUwE9q93rBXlcjMOOgJz5TiOzAtMtokUGYExFAaq5j5TnnX
1OBdhLmOUnp6fdsIW0NhOCkTUyfKcSWPMYfnBi2uuz6BrDd+xffMldIUn2ZdcG+UXwi30lcwRU2r
XLtY0SaoU8OGAAmsj6nID1yW4SoxkBVupkWFo/6cMd7inKuVwlT4gOgbvhh/cRVxYvlB/Kbl2DGU
vmwF04nPiDqbEHgNB7EJvDb5Skq3gVshkjCrTGGpq5hWkOv+pi9E1Uxn1tOcpxOKanEs1B1Bh6ch
v7M4TAm68n9DPg1YdRArLm83sgUw2acZ0nyiRaMvXUiHhEEZxxpin4kzsk6Q84ET8vOtuXjgI9Eq
kKeYIsXSs1YvIsJjgxuzmvxyVye0ubH5sf+GpLv0Pd2ihaO25bfRXWdCxUcDO6zEENkaWP6SY1mR
oezvhc3xG/d6SZHzEDNwbCZKSG/CTvOUdsE1oxrraUKJjG0g+wJJJkcz9qfZ0w/WxsDDOrfHfCsG
6YXPjqvxDZ9ElRwd2Khrl+xLOZ0nfUGf8+NgBxhg4Lhu5jFKtLlMrwB5g/bCqK8SgBQI4pRPp9Fx
KDruQtbBGjxfQ9N/G5h083JIgjkRHzSHWHULEguBH0VfX33x9PsxQ0TfabjsY0mDNBojX7d6/3dQ
S3S6ZHWUsph7FIo5dukNbhpRbPUpyHFgTN28bPjA137JhoykSAiD8Zjp2iV6GR0Qdi82r9SMWur9
OS/va2qa725/sLDcODnNSc0yyFLL4D3v126fDxQ7EUZY5tT+EF56C2UYCaCEp9nzlsa90MudPl7M
a15FRnfiNVeRT5v3uTpyYMi+ehe0rr+ZzJ8VlNkBvyraqTRIahSZ/W6yYHltJ3WtW8NxRGmCNS7b
Q9f93Ha1XSQSeYuTqmCbjYh0nAIMi5ILBIWcJjnMj0KcZKnCv/KsqL7jp1sqPSJx2EepN1LHN4zj
UFja3c/icAUVK1fKxjXkqeHlYmubSLTlRn7JOGtcStKIrb4DKYziKp2Dau5HDKoMF6/IXxtnYXEv
IQC0FmRcyB16PA9PFk8dwLz/9lIHJ8AxCvwMSMRcwoETVG/dEBrkU3+hUpJYkqVdvHKdABZlxkgN
yFHCISO8TpF8tmBWAHF3MKZnm+KiBsFDOjFhOsG28wPNx9HKxIaVHJnQZIBn8hR3tXH2lz3wQOn7
9Bl4kQNxjLo4UTkD2yHdXYYyFChKPkT3XlIR0OIagBLzeF4+Ve2lWgXw19fuEIf3DFGWZ1XXBPNH
7f0I8MMKG19MxgjIX3lqaVeRKUf3EQ1tH0K4C5XM43Jm8KrOJAe5KuspM4/un4UC2jUgSGwpNDRX
DHePl4NKgIZjptT3ALyPXlicI9mYhQ3kEmS6dROoUeRVw/NJ92KijoSB3hwGsvJNbUDaVYW58heA
u5tll92ha/jaB+0ZqBS/lOzHcmPP+IGdoZ2GMqdxPU9sAo96dOtiw7BBeocVZ7pZEH+qSYFgmd5P
uV8HbM0wYrUkKdO5d2ytW31BFFU9WLshCavEfj4UeSfW0hV3N8NqWINt+jE7Ed977SyEZLsZ9YPT
B79Cv6wMd7s/HonJlOyEeRooqBjsXOZlO1S0iNO2RmAhSafptSXEuosXOTy5f4mPf8WNd7a2OSNm
WzHxg9iqVMb/v77udcfbWwir2/Wmt86aoFOAJ6tufw8lLahjdpMVlX96YVCk5GNGHsEi1VMEXWls
g/7xLnogmfPfAc6va6Yd8OLE5BWLsb8mykEYwccB1lMGpEa74D0UwhNcP6u4aRIUZ9aJ38NL3KfY
GIJ/nutvFuiyeGOICiNEyZ3JVIykrpf8F7vOQZuIkB9LLE7QmhsTnGJrqHBfFlg5M+JHGzcIIgW0
nrDfUhQUPvER5nwYpN56C1nwFkvm4XdvssGfC1grAmt0Bhr+Z6YqCztl+bfQrIiI7qK7M7w0ayVQ
T7eg1QT7b/Dy2+lyWmK4eaKK2G3/wK3HomccUTjFjtcpBM2VnT2FarMmT3T6KxiwMkwhaiqK/fOP
6VKsAIfHvSHsp6nCTadROkykeBkv41JCtLNolBP6SK5/sVuTXmbhvr+KwSVLXzn9mzCcz/cHtO0A
5lCIkkuKzoyVspgDf1uz3uNwDKIttMGESgLO3wAnzwCm4bZF5LVrdKlLrCjh2qv8dJFuWO0VVzIM
u8TTOlWlqs05XdBsfU02J6gusMhkoGZv4j7sNKeGe+1wTo28eFk4MOuUth96/Ow3FWaQ2QskUjwI
hC0xKZBxMr47iLxZH0UeoMDY+8syB71RnTGaIa3QhllbTJvuq/BljV24u48wxVH6O9jw+1gY5Jaj
cXWj/uCHM/BrTxjDetQq29wRNdOovo32yJ3PCAoxdeONHnK8QuI+cs3H8uGXf7ViU2B+uJi0NFfp
iPkvJmLCOM3u4V8IQKV7i8g0cZp9q0yN5+eEZftdDhQwCs/oMGvWVbRPp13J/62SgabZ22pOTK1W
f/BmdO8NY+oBt9jkWm5FfjF2hpgSUWWf5j1os/lqSjDGxk/Zxw6npt/T9gqw2EaH/jsHt6TY8uXh
Vy28DnmQVFi785hyLIanTUg0NMJkq7ayr686+Mn874uwJXk+RtmqW39uX159+pKvQTB4VFINbxcj
sqDKk/5jGQv2piIfs211/nvTOudI2Z7WfxFPjtY83XVbJr1tOX1EZBsJT+BZkLzIoKa8Xb2HhQUA
uqdtVLkJVOyasWCHPizi3ofV5HaYaPhmOYbtNk8/vul8YFyNrejYgIIDsfYSxg36uyeAWMcakv+R
r3ARCUBed766lrw0QltRg6pqw5fSDJKHBpVsjl7paBCwf4VB/9t+nraUHqOlbJoKOYzRVtqBnpgj
HN70ITYXSYxVs3aGPVUtlYMyEGG/bxEshwqinJh0XKAWhRM3cSAtOxPh6rPNGKDgc2D4fQGaiEEu
Cjz05YZtNlu9o6p1FKrcz95nZYcSCGwjszouFS9Ee4YJX8cwrgn14+Op4NXpukqLVkh3KlKWcX32
R4KxJmF52w8vY0kS4QjDFUmcH3jUtsUXZHnkLCLZU67Wo+h5gMsiLnyR5NZpcYJw/bNLc9LsMjmR
Xo+NEOlCs5n51QmE/Ey94PLbqddbTSug0SiwgmTyzFu0UPh2uNXYkt6tHYYSxi1uCg6wzznGwhO2
4z+5QVbD1ysMIpVqyEHgYk5APvW1K502fobJdF3s2CXI4471nViS4AILexY+QezRB530seOiJvGu
X6rQ3pU2ryjxXIr5fK+LWYK+BiJW0Rz0Y4rPN1J7XokdXTitVbawbh5U6Mgj51//qErDpq4V75CQ
r14qNgvlSFtjKkrPFZxjYmW7sjg/ud6k+5vH1Xi4O/+oiUvgnVCVSTQ35ZXcIZ3NBUs+C5j+Hnqm
somMx5Je+lWqvu29ncwTrnpUaS9y6NYHKE3xNSCssbZrNxfRQVaN8+a/Yz8gu6MDrQz9xAug05gl
wQJI5jejjMZUnahJmmfYLwwIGqc/t5GvPwDmpgnj+JR/MS0eyEgqufFvmNUA/h6CdDVaUhceq9x1
pGahcu47JRRwG2NDWHZmZhShdlfd2BovTcPT4Z9/dlxEfyL9NzyJNsb69vWM/ExvDMO4sCopvuFs
S1ykFBR8j5q3RHZozTrzppy8Nimwk8okMUeFkHmlfB8Utyzm1v5DmWKoI78jxnMPH1ybrPlw/1XA
w+Z8E4LAx0oiO/HT/n2nXkY5099yRU1U/zIBM9XZ8c1BKhhcEheanQJ9TMuUMYRe9xTCVqbosgMz
DEHjqu1tN+oSWRxCLNTHCAxVxipzYerdma0SD9MdqZn6lrlC6BRATX8GWFsWPiOum2u0AvuhB4Pb
JhJNJFxqZgttSi9+4x5M7m5briKw3a4m01Mk2Pgy/7Do4JDZayfURYV/F1rTJ5/FAQNtIcbGNl/b
j/5zylm77ctlIjRGMiE09E6dszN+5Lks8u9aCJlEZx1MdB3vMxd+pYWHSpj8BHP37uV813mAQtPK
Z5WA6dGOATBH3Th12bKKSq1KwVfiGxUW1IAtaBECHWJVF3c9sRm3v9MyOy1J5/qBwk028b/yQ+Do
oJ2aWPTrRZ/D9XxMaZQ3+ltHP2VmxlDtAA6UYaN5uSvn9DKqMTFwQkYG9hn5RroLsz8Ne50cJX5x
iV8y/JMmrHpOWEK67zVTQCzmVHo/MoyCZUor5Gk+dYv7wYp1kvSqrnC56AJpNuubZumr4MotCaSl
42wv5TQmiHxrzK052WbugUI9/TdWCUC+gGGLeZ0nmJ8HpZAbt8gvFjHt8cgbBCzlvRv8RnIlIhxB
Dppm75ICDX8+64xaOeqwOG8R+mpLgYNF9wTvJVSe6p1T4mZe+2Ld2beA+KvmTmU8bkIpKrS1CtmZ
lxUKYFlpVyTjf3NwWK9ZF/mY6IfTE7YwJSycjVQBqAwOgyC0aWVTMWjiuyoEkAlPvvQzswo6pA6o
W1E6zx3hor4C+K/Lts776DcSFqxJ5q7h/YB6qNR5LahHbe5vKLerq+lhKYX/silPNZoDLOrO9v4g
x97dcpJFC2/Jwimm7oFFrpPiOF2Q+hWd3DCubL5owskVoQNRWhpaJFqxpSqbgbm12K9x+fbL+Ri6
lfwuT7FpTRXaYlzk01mCVZePYHA1DfcIqhQoYV3vlukBU+Ee1a7Ul/gX+t43kAkB6rD+KnrrkTG6
LWfxELSEPuFR4MtKmEwLpuHGWFfUVvfR5pxsB289o736AlUGlId+TaFEnFazRG+TkV0rWCY2sO8B
n9EK3gF07E83KxPUXOUFWGLALRX5Sboer+pHy1uamX3Q/rvF4JIqGj98gA1yr53krS4E+jFq0s8+
40uG0T9gXoL7DbxsuRApDrcYk5YyhQjE889CIWJQwZNUyNVDeteSD8SRQtfd1o4yZsHCvkYCtDuY
yS5d5soe4yAnepbO0L4hSaiIjtpkOnGT1aSlYTokqCop54Gki0R6Wrui5zWHtKFLe4nyRah1xOJ9
BXZqKqke0WLrQPloJQbirsBItBWziP6VGauEDA71jJ8CsizRwjIgs+1z6nNjlngTRaiMtRBKNeW9
ShYol8Wx4Srw3Z2j001MWqxIu+fCUVuS12UUER/W2iiCW7AsFODRKbqG+LlzbGifRdKU/h6BDcnc
hKYYzPW4mF35Bf3fbwsbPk5FkHJ2Aolhuv2zWnSmLRQzK4GfUFnohLniMgG82GMoRmecnm762h1r
a4gAQfFIoHERNsw+rWqNM+qDCgWO3UGAtsFX+DucZ3VSHb5gUH+hR80sW31LGkhP447wk1iZ9/CH
x5H7MrJxGNFTYHotz4xuTIu4FIHsV29XaD3cnNYQj7P12EPMmCHg0WXMXBFy9REKkQPbZTCvf71Q
z0a+HdnLQns/VC9vFXUthMgLQSUFLfdBvyqhsVPQoHKDHl5XeiZtsa6w9diXSF/VuzfLN5si8t/U
qSZQ1VPFEOeXMsHGxPYigYXuylMvVJjqBZGKhfGualHrgkHyVigjPVTQrX5JueFccWpHIOfZXXhF
hNcjyqQLhRHqycW5K0ZlvOll6nQ6bEDVxzBImXBzQyj/5ez4dmclgYKUY3aRbOVZWYY08miA5Zxr
Oyi9OgQbfTSEbbA19zpggeKctxh1KIEFD9ufNmRMPM0p4f//7kS5MEOPP21F3+dJLNw5jm+nsoln
HFsce+K13DnX43NwdewawaoBArlHGHkWoPLeqtrfFFEyJH7515KzEeJ6Gzs/M86VaPg9EFAFpFHp
KepWZYSqna/bTUQYMpm4ewj72ysjYf29hIqHzFljhHWuj27yo6wf5izm8mcAIryMhIRK10I6aqyC
k15jkseRV/F45JqvF5TzfLueyV4GsB+VFJrHDI9s9xQ5zO3fzc/sasSyaDZSZfvid6j8ZtYRSMJ9
WT1/qRGh8bgBd89amMBVSPjvKIUfd0QLJUZiA/jshuB6rjCkHpo3jg8TySa5G6LpiELO605k9TfX
sGorG5nUnRzeye7XyPSbeKIeaeiq94p/DxFvwj/hzBDbU1ytArxgrUyasr70Y/uNYu5yovf0gq3c
8n6fn2zWj7+eIBQqG+hUpgJYDt2yI1eAcC40aQgaYUIdIGLCa1sIcWCP/z0kC41fNju8zXSxCp5b
t8VBYQcUN0Gkb8nW2/wRW0v2CNHOPTVtZleQMind2KyheqjpTMTR/wCXKls0vebFNOv9apE1Fgw3
isnZleGVX7mgmNRhnkM+f0q8D219znGl3+nW4BaFiJ3UJAql4Xp2aGwMxLyFc7firrrB4w65KYdl
d/cIj/q2+YLYwJysfeM65Pod1nMv5bH/y7qF6ZAF0LWigjSTOWXNKTPiWhQ8XgYTTSFqO6K4234e
SAephZwR0mrj19a/mx289NOAE5abBpHF38K83icTu92gwJVmUWRHsGnH5fwLAsBD8Uq71vKqq2gC
o2UigjJVrXHgCLxeVnNCZtRjk7THKM7aDJ21XK+r9gQqF80KdvG2XR0j5wJT1D1gTivqlhPaVW+j
q6yg+pXScTCdQRXHQyAmfw1X1miEL2j4R3uoEWBRailb9CiuhAtNr37XqqZidRBi7cTbC86VL0Jz
lxJz8L150wNnulDvrKvSyYY3fW3eJRjVHCm5XyVAF/Zi0tGVqFf1BQpvXdOxULoRa/gCC4M5VpZ0
pxIP96ul73NbxgDXet2WRUFjSqoR5kRQUdwyZkAEnz48GPvCXQejguKiTlaOTY16Zazc10Ojv7ZZ
0R+A7cnPMF+U4hpOtFTQGbCqrQmGlr9ykQhitAF5CDbNF0cKzn5H0fvuwjYVFNax8uDG/rTnMvPp
Ot+GFkighEihe7FNCrVIHNF+mQWsATsozSa2X+sw8iIb4+AQumbTEokimRy+60pHz+KGvVKX7ltf
nXzEcerccrrx+tFAPZLGlqmGrJOQhpDPyXGg5PeT5HWPCZy3tbZfchAk/gOi5HXgEIbuuATeHs9m
W+fk47gcdSDt3FhDAtqqVM7+kLu6k0lOVT8MdS8v1mq42WRDpuxB1bFIB01FRs7abvtcq/4HndCM
RCO4CQojc/ZhPz4ml9/fDaJrCZRyG4hBDwW24qY0Z9M/lBa7dAZezrvLMKaa/0UOz4Q6LOdi0AcP
/y0uU/y5jjZtXeDWbvJ7lWrLDZl86Pch67264wA32mBGZcgJIrlaWrBrOqGmhjSwUlZLhgZwG0JE
ky2S5GKyK+LNtPEKEVuLe8v/qKEsXxVMXx+G25nzALI++8lHU/8DDBOyDsYg6l4Vqtw+ymzeKB8N
nd9r3VIu99xXKT0srWeIdU73b0cu/ZSfBMDoJKHCb18qmoN+WKw3UyAbgXYbXMFIcFZzhKIwHp+5
cxeKyFE6ih6MJCpzIG1HU5FfPSQf4lGVpgunw42ZpQQqcbChBuWv0MAqh4lV6gok6+buV6AXDGr+
rj5XLJo1SR2fzy1frLlFs0iXtlkvWyZFGiGctxPKzMy7X50hbBwtnpUXmvz8yY46p7XKql9oSQBk
BrjVlW/aGWbgt23zRhpCg5BbkVnjm0kB4u5jHIm4p7YhxZZehexckde4eDKcmkbD8az8TmUQ+MJH
FuRH0pFdP76qPsdop/lp6taRXEcohI/W+2GhU9ZHM1i/xaYtY0Wwi6lJequnmidA3DCgu3vY7uEE
986ptxEQEqeooCgp36q8hE6H7SgqExeGJ/afzFTQExBlH2ecZ3QFj+C2Cchw++rIiv07EjQf3607
ToIXm58ang9GMTJ6wUoopPvV0eVKdxKnzU7LF4U0HJ8SyM1UJWeEtHNgs/sKlJcbiL93ccIUwuHM
cmgKrsB3K8DdxQMVhEomcfZCqR5Z3CqDKdp4tbZMXzXCdAaCwG5kSf8ZIHgIY/dHWwQ7W9B7GLLa
dTIcwey9GbYInGhqEI9iCMib2cnhYwLO7bXV+OjubNNoLK9H/qeWHdZ6GCnG2odOaLHOzQv+ZIOg
KXtTkgBCRU37NNIpplk9AP5fwgpq6YC447DCiqyGJjRZECT0jRCzHY3DEPHySKei7Myoz8EQMpEU
eh4uu1KtYJKmVpJN4AxFaUSokxWPx0jNyfE+/Pen7PCoW1hcImbbIzpEocQ9NbWL1RC80H5LTTWm
S8JJFFlTidohoYoGDhFzOsq+ERSF2l4JjyIcjhn2jOhFdqNKqRIID8xtDcph47akITK2dmZppTFl
XVreKor5C87SZZvpwkRh5kXl0/acWxmZ66sICnaMzSgZZYbCs4hWKLq3C6F3Q6L+SY4if+zAIP4Z
Rac4Fu8F7chPPtaxWOoW5BTOp4wsfwuLhddoQ6eEDR14PyslrIH2L1cqBZ0HzkNfmgrdTGTNQFTA
K3Qnh+XDT67wh2tBzaDouE+GYZuzUmrbx1wBOkMNlw4ihn574ei6iGYtObrs1QRarMQbMC5e0Rhg
xu3/KBDXPTVeZtoubv5Vh0NsEtlGBub0b2AwaS8uQ4j4k3+FBv/dbIH2b/x28FWsZk8vUKdsarXg
nxV97PUufO/LHBg1eHU+daQMh1MZGhgPotzxp4I+eIt7u7QYVtxuewixJbBuLAXzFWWX9tYZWW4j
5B07j7OM15oYZySs+ZcauKuFt/+k26RaPuegiGWTIVP3n2avtM4z4C0QIPlIgpfc+GQcRB9H5Dgv
LeL+Mjbn2XxY4ADjb90lCTOTVkzxhDVjYP724i0/0MIBm0aPRQS/9QV766tZWigtFqx8YwFUkJNh
FYikXoOEEfMliPmOqKshYqvMcgXQdXK5wc34i8EbKc3RUd28u4ItfHQuv00M25FyHhKpa+FGOQO3
jSgmZcfufBzMi8e11JMrvpqhpT+gcElYEtsg01VcWi9BEsLegPCJwvc+R6OZfZIEzimAmzqHN4/U
8EQH2JipVjuEr7rOV7gEFULEwEZJ8Ut5BdYubLsYIHQNvYBfocxdB11CLZGCH5VKCY4jr7fYM0Yu
ocAWsnTwiySY52iQzoLaG6LkUW+Veq9iVoLbRABNrAEBf04QLvaC5NNDv+kx5uWH7T+Kor0D0OkM
IHzU2pRusl8zT4XqW+W0ce9W0CO1mXP4seZapH+8f1FsosWZL+5YSPeX8MO1Pq0jKUKzDH26YR+m
2ZsiRXJr076Wlpno78WTPYvo48k1uFVBNhgl9/W7QuYouWhmI8q8nciczDerfRSjHbE2mp3AOgy4
j0uafOLDAX/pN3FDr5g2LolvlksJmhk6WFX5gqzdzuNBpIAz61dP4NIkLD/Va8PXOaVkffxUagvT
AP+tnUpOCa6rh8P7xoB1pKtZ4AIly+uU5BYQoMWV3diX/ABsI/IjFAB4dVvPypu0fB87dLdOZOZs
KgANqwtUTlyKxCp9ptPwLeQEf4v2jKu9NG79cbvkDzG7APA23oPrmjFtyqpbjTv2t7D8ygxNYm84
KK6LTpgQAmrzF1IT2uGCknKEf+OATPOM1rTJLtVCVgXvPqoAD6XDLyxx9pvo1euP2F56wBU3ctNM
5duz4ZCvUueuMXe/36Ad1yn7+YupRx27UUowdt8AJe9b4cIxSALxaaCCRFwy+O8W6/fYnxT02luF
zfWSRTeg6onqSXl1VisFrggs8wsVu1bfaZ2nieOdZSBezgISUCrwEZ2hVY4OdNbhCzDdroqObZih
CGEoI6NAA0lSO1k3BKCkqltJ+XQDTPblXEpkxbdc6sDyFgSvJc4wSOunr76THlJT8YrJoCy6K06/
8FmolfDmY+GmIo+iTuCl3fts0NHsj3cZSMeG/vRRDQunzSZDBvu1zIS4rdj7c+qK+HOYwfUQdrJO
BNn5P6FomBS96SLsZgWrNYw4Mx/S6JCuX6QSX8euthoewG4DCqgepLohgl2SP+W3ZrjjiVILRq0v
+zzx0decXefnT28a1eKNH1M0BnsxZX0mzULFev8PPJ6nDLMXusS7UF3Qg6NAy0ZQRJYJuKdxFz26
6ZxrlPl2qLTf8n/4eNJcJFsWTVFgrjjlnuIgmJiWj6vKMLr7acqtO/7FX4n2FXNDmF6D99/QHfQ4
pabh4CdZ4OSXI6kKIe2OXY/3PscR3al8WFAnd9AQvdWaA8rBYZ7QYpQveT98WggPqbuw5xcxM44R
7JNGEet8TWVwanssI9ef0Pj+v4+NWRDyuw125WrJpLz1owyJBmC20d2EChuH3VAkYcp1vYDLwU+n
i3I607KnbSP/Y9QSna3+Y2Rm9s5ZxIl5EZOAMy0ojrRhZ4+JStEuJUoaGX5KxIP5qVE6y8RkILfR
Jj/k4LHvk4P3FjCmOPPQR81im+i6fxH91pyArTLHeiCZge5p+bEnJD06XYEn1U/fgYUmUGj+ISNQ
3/nzUVt/mA8u5SWNa35tI7sS/v+8Kqms91y7id61xsUE+xiIBa8ZMZ3xRWZ4QYlKyJnbARj/bkXu
ZI6gBIF0a6wHjH8ju5cEW2TCxViZ53JemKDRXk6uz+V0Ra+wzrcR4Iqkz2/wisuJxiOOiEBWWc5g
ippkq5cozfx2TvvJ/BpM7Gx7Kd7qJ+V9NMWXI84qEimNxi97gt/OhH6afFV+ohiyCL1/V25OEYza
moB5ZjyoeI6VAYiwXGoKU5Ob8ybfLVUmknKEwIJoYavy4+0FILaCB/0LrIiAMcZpZgqXbzoynLif
nOXiDGkSLPuc950InoqFkYwut5jAjAmoqmBnOIgyt02eky/DOsw9dKdqLdr28hncO3d+GRvRVYps
VqfjD6M7NVp0gvKpNsyMM/o1kKFRjlK1lM4VraV0C+GD6s39kLdrvYDc9+7t3sOq37De+bSU9M4y
5omdAAbIvF0NTjmZ+S2tG71niveCziz2YLPbHDGaD90nCsFsh2u1Ugp3lMaek1DgCqZ25QGJz26o
llM2YOi9ZSljCtpVPfC1lANqSk4j7SloLfowvvIhKvQZ6PXzqmBsY9G6URPQ06AEufx5Cl0LEOIz
L5ZZbyZnUhq5kaj3brhnjkNLUjQAdXEfRabFOLiFF9BLuvsI5V69K6dxxx1iiiCaCXG2BeA9SOc0
1Un7ytQSUyjWiCpd6dgZvfABPDEHOZ1Iuriz8Qzqhuo1J+91EPoYFAkS3yADWXtLtPE/qvrjaKTI
TMnsGnBIoS7uGuUZJhlSnQFJq8ebOuRDQWr3tNtM/MArxDFNFshLnrqEQxA5/wW7SnZB7fGewVwO
bFRpHrVmvCJJTiwbK4CWvRp+8t+m5pXfU8lVFVsg0wSFkMwVy0/KyOPt3R4bL3nSNsRIhW2+/UJJ
9bQHfpqkOwD1ALsMByQmk1nozkkYfm07FjW6Pr9KzjDFeQBJfa2QczVPOgqlxrpgvgY9yNEcIOEJ
RE4bZXWX6W5Z7GMVVgbsrqCp0X5GOXJf8GiDeXgoFQLPIJGPWrxYkEWx319LCGoufP/jWLXryXUt
QESvnXIG0FdcA9i29+ejgdibpfjVNh5wr5eqDC6ANZ+RCCVO/HngmlIix+5ne4rNj8Z0gZiMXXWm
Us3Um7y8SgTbEeMRjLGoCqfj9sGlrOiXnUBKpOlTcIggZdy4iMFXtk6o1oQaF0zqIu0muhe1pvmr
00ohrRMM8z8T7U2ExVJukFwI1mz0NnGOJaYuZw1ugh92NUt1pEirMHJymVT9rvj4F5LTJFnsyHMB
7oJWyyb0KDXDCtH6EGWDOrLWTLRm5BZsFV0Dg2PzVRBvDRLasDKigIbfgiaXRZMBVDt196MjIuQB
RGU0HvPwJtHEmGj3+5K22HwgckfM7bLdMnmhkUM/BTUUGNJa7uya0T0mWM/RZtlVTDfbURXx7bh4
KPPKrJ9GjqJuIfEDVZ4+DwLIJmjrXPWCERmnHx0vlYW8iFezI441xmIKT45JUmGWwUeYqYCTPjZ1
k9R3I8lUvdK655W+onsMsYsW5X8R+a6z4FuUx2OLvWAFGX/7kUy9XYk15zVmk76tPHcIQ13m7hp1
ZOmBS/InoQUvbHZYdXkoj2T3H9UdOXjJMmHqzb/dQZXfSUFMR5OpH3mA/ar4/2KBLn4/FqcAp0QS
ELMBkODD1SzDgN2rP1jwHpCYU9aAElDkPQhOrFrEV/PLzIdjAC1SppKq1iWZy7owna8qoLSr5hJE
YZu+ddKLPC2YJ8/DAsC90ruDMame2HAnfx91fZqRAHzafghpvks1lBkO824SRf9DY5uJgD+sVdTi
2xa7r5XALXVAkdXPudfSp/NtoJL4TPTtaZMWX/THPgDPGMN6GmYYsrJyRS+v4WIxSE97+1VqTYwo
Zwz+Tw/DDH8YWK2EP5DOKK6Av3CUXKbk6BnJeGH/Jif0CBwgVJfEEwmUcZbS5Y9M9ET41c4xmboh
9fQo3vOkLhE+5iXUIslgvmwL5+z5VGyl03lGu/hCnk/r75x+XmSk2leOCkyVYDhd2Z83UjB1oIAa
6FMaJP7RN0DiAtZE/pSQR/8f8N6w+T853WAr98rJst5OgynhYbFjL5qZdb4f31ETlixMoakBanb5
XKB5u9cAZZi5zmYZkesrKFbCpdGpJOsRc9fYNOmBzUMM+wWxuFi9bCKRoiVEtM2oIZqwAE+3B19V
eyOHFiBMQ/HRi1gDHOdEV5f0zomMwrKY5r5InTGy/VBhu+/dA2PfPfvgopL3NMjElD0AckmLHLG4
rG2rjU+rJ6I/dQMfEhWJjn8ODHxcc9W1GwJmTQR+4tkq4kciwc5obnfy8+swudHhmUj+H+xaStCY
QpTQbJBQhqy2delkv8WZwrGp95yx2jfTCsVmXPNtcvKHOb0ROUxKJEhHaD6tnzHyX6xdhD0Cq4WJ
hinBofKP0sD5G251RkV/4YjS6foeU8ugCDbhb6dtFR14UaOAfK3X6lmbJDfk2mB+XTTOR6bJ9sy2
EtiDTfOcHcjebGG1UC1+zySRKe0g/lzwmGr0Fm5Q05xdUKE9/Un0kpXyB1quHIohUOlysO6DlMx8
VlYdVMMriyJHSyRFtvkyTfmDD8P/wsyby30Dk5UCXlT8CNSTvrqsFLWIDSyAFRv2Q0Z6xPfTnr3Y
MRaus/H9xv9+Hw6DL+Pm3FcqxjTWQwebJmjuU95W2L+Hs59xAOXRp/urCkMGnaOt9wV0WEzIdxqm
5W8SfAIL4zJEfupkSSsPwuHuY7IY5fvlVrCAGtejUuIc5dubR4YR+pZJdprzq8iZL/uUMmQpSn2+
EfcqDpBBRHIw0kvNWK1/duRT/m3mNLsBhFxLANlCCAilZr5d/teq2FFpeA07E4lKG/cwgK3Em59s
CLj4Lt2TI3wrpKclEhPYZOz/0PmTJQ==
`protect end_protected
