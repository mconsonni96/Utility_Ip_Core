`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
oupg+nRLrrAYA/XTaIUJRBDxCh78jXrLO5trRwMVBK0m3z7FmJmFxHu1hiljgS69ri7wf6dUtvr6
PnIyqtD82HghmA7IAlcj+AxhUmdynvmU6lcvSlhSnsSKEDDEV+Sal8NpBci4rdX2dilBi64+5iWd
ABeuzWhRKIS1esMjkwbQ93Ahb+/fYf8wr97wtcmiD1YIrzhyFl6guHi5o6DuUJddWKbzKbvehqAe
o+QuMxCOxJHiO8/XnFJFZJuuwPK3sCam+WdRAXXDKkkecKBiebM/+GMWza2EiuFopfs0VJN//wTR
l+pbzbiDZ2EXNXKXyMN92y1vx3Izs1NmyRp1Ow==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="udGRxwFfwQ4jEUGJsrl+/43Ef7rdJdHKCEjEMl7Erfo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11648)
`protect data_block
YY+xZNXkvHqUccGY6dmCWzGxW3QZmcwuuvH5EB6IUL+XYcBOo61GRinSx936U/H3lYUTiFEYhyTC
MpqetbttGITQQTQI7sVxIlh01WQW6kMIjP46brPxHqGPe69uP6u+GjrY0wv0ki9b5ntmaWxHBZZe
WUez5VEyR0zf+W/mt9AJesm8TBLpBdokHKC3UcMQTmtOogYlccwhFC2ulfi3IeO+7euVl9IgdNAT
hpiSCAbVaicDNSuXikd8Bbrf6ifxL/JtRzK+01b5nrxSkRVRch8MxLjeEwr+FCwxU+hP9jZUIoin
CKLYH7Gb22jVPEwI1YnRfwwnrLZzhTJOLHS6TNCkmeyrSHtkqNRjpnpAyGfluvD2ocwra5WUAAx/
G/fSJ8yEsVvrMH+F6kCmJ0+CzEr1m+EWWpIwGafIIZBUxhAkKeQQx2VwkVd6LYUYNOueBwJ4UCh9
BhEYDb7Qkrg8RjuzhBkxGRDhHWdKnFfe1WqpCwtHzjVvp2lIQH0SmgwmasJ0CY9+T2cRrZ8AagO/
QGWb0QlJEhpP2UfWGIqZ/FQFFaOFYoqYe30uuKzNDdKztRkQ2x7aiTtmtUapIN5uNWT+mGgllKhZ
Lft41/eKfLDos0d+mvolHz31qzgbQCxbq+F791Hxj9HsixTIldnAs3gpTiG5WI58meM1G14/m9hp
Z5hEkjlWGVLCu6mO8OBES5gFAfFwmOP9MsO0xeM0GtUIdTJ+hl74vH2f5aCMa6qmoPdJuvZ0flSc
ch7bcSW8D8Emx02+3Oigt5F/vYGM5V3ELOuNQatkf09F8F+pJDXyLgl/x637UgWVQzwW0+zGEJbg
PrHzRhozphWQVSUgbO7Ic54ydqVXHo8zVpD1Sx3Fxr1c4RhNw60Wu+mEF+1a8sIO6uPT4tCUcBvb
6XT2owHz9jC2FpTpYaMiPaf3hEkh0HyLF0vXfDD8pW/Npp6yjmNzeqHDI2tbeEsLhbKJcHN2tR5B
HlI3EpDsxWqmGQFMWmU+D1llTniPmbyyenGt9Z/B0q8wJxaKVOkn179iIJdU//viwbEMBQ7rzwbM
sk01IRppCqD5qQA134Vv3hJtM8nt6AAONqJoI0wR5X1p0R/quLbVxuiFnshG29tWQTo5vvzci5Tf
7EwN59meNgQkduY5kx18jqAJdfSk1OnLc+NHqWztGasThFYZ7ARMoelmvtTHW3aZhT88FKToxo+7
laR9KL+fYDZVhpLsF2LoV/e4itCM4aeeD/lTIOAzA7YpnjymZRWfvbEKuZe9cPt5+XKGVS9se2od
S9jJoY/Ak+WSGypSAQnr6WNMRF3l0i+EKV2A6daRk1SRbQ+qR38PteI+Ic6voM9H69RbfRvdsCWP
bZ0/9aQg4VtUHa5YJQpCYMNATvtGN5q6ycQVsdvf2Jfsf7GdaJP0KSBVoPceX9b3ciZljJSUXeMh
cmPdhMy5AM1ZPQdd7knkkjWJIa99J6XRCvqrPvq1yti6MHTZUZG9ELlSFIL6gQXBx33Mh08fWIB3
jpFm/iCFG+PnPlRBgAivSn/slxuBF7Wxykcpunjc5uyph8u5FENWUnsEI2Zvag7A17vkfKdv3+eu
U0x7adFKg6Txn42lHu9H6W+Xoi0SMghwtlurrHlHJpZsg74VQe9Vbhe1+vea4BgnrNXLxTQpYZYM
VlR2sMTsCTJicWP1iNXp2kNSRaAU6RDKHkQgZtPNQRqZSKYfQ0MIRkGuZWvJZzpSgQbyynMCYLJG
awVBcoSu5dhlqhKmlgBAfxp2Ut64T8gEaN2Khk1NBfcQUQo1qAaRgGzFpP5WxmWxF60hkjA+AUvP
g5nfQPid+kOdxnTtugmzlz7C+0yat+rH81w5UiN1NGjo4+n+lMPAN8dSYCxyK5NSyG5iO5S9mKAI
2PmCfuHZk26RGTOakQ6+QoLziZj1yG0fiPpMwH+eB29sRT1WQNk+ZwC+EpKG5RiElT7rH9lLpiDL
oKtuAK2IwIzD6NE0d2vktzT3b6RS8ztp1GD+uB6rFop3FvzuYPpgsIEMwdpNYm+KlJ7GjInpDjAL
DvmqfTc/VUck9kZofPR55Q26psNWWGPMgnCNUFZJUKQx9SrRvW2skRAgSQe191ipQRTTYx/eh7+U
sn+1qGjXHHDPVWLBzJeeDvHK4Ar6MNsIpZbXtjNApo+Kz4Z6nwS9IW5pok/FCqdauMVDDm5mszB4
wYqNQMMnt0OWNzuK4TRrzrTP5crbeVePdDHpUekuOwV7GaMw7/+eDEUL6vDV7g6OEnaJ/Tnw5xPE
db33yywRY3p6cY5dmQR0XronZN+2+uhseg1WeKVUlfBybpRHcorkmdSTM/eSE950G2VWKxq463mg
dl0bScHLgtNpdq9tcfCi+Gq8EiNSU/XMy5DZeCC1+6z5i5GUJhMjSIbop3rvICnj6fAHk++Z+oTd
fYUWs8LYWwQK9mSbwpk662qiOmQFgZcQSdK7MTg4EHwWjYUdVtdT1mEC0J4wRSeYNox87FDfAyQ8
Bfp+NInmsipRN7ZOr+qKG7pqT47P9X3iUaNugm+0LUSPySo6z5dhJOxME437mzb2FDzvLqL9/1ky
yO3uMGFa/t28AtGMTI1KCOcrfJjZ90JaLrN4effg+iBN+fUhkY4/hzv4HuC4ivXivjq3Vrjy+T8e
rGaUTNbeq7WgyFyWmJ3Z8x3JtEmP0STHFKSGwUKDkeiEmEYKTq1EX3hkWQE/FRawNJP+oumb/HJl
vqQdpbKpdgrWeHoQrTnRfmDT8LNUFU5ubfMu3LqaCRJJxIe2eab37ntt0f0ydFoX41465cbFuqSO
IlMCLk9nuq2ypLMPH1r5F1UFWdBtMgTnHAyw3EOIzL7Cnt2n5ewUVG3PkcTNG/h3/TW7VklF1++r
PkDN/gCcLwNj8G+IJswqzpaAvvfwRtLN7wo8OpX/CqpLL9MTO8hAIFqc76eNT1+xuYGOOuIqT8DJ
AsPHWmaKTNhjfiVIASvk04ydJUulnbahMALay4VZ94GeJ6kOsFJVPh4TN07l7c56BurwYB6/wzen
byRE0a12DAh42zZt/cOaN9VCIPVoPtMgO3yQqaVJfOTuLVzfH8yee0a/wJMY8IfDkOmNk+yyy3tb
QpLmNL9/b0tFPtPJ+8w3rykVqSTx8TV5tWE6OkkaMbTgE0jUnkBnlDVKAAjVIMK4W5nylXGG1g/r
IEOs2Svf/pdXBDSnrW2XIieuYTiFXXg7JFqZ1O+q80JE6uGz73AEjnVer+iERJp2f8449vrIqx7/
mBnRsGt4BHu4FEXsm84zOfVkP7iqCK3+GqcbUQUrNr886lrLn+GH5cP1Shfs8imTzNaHLt/WcZcL
nEc2i9oaYJJ1/TdpD9Lw2Y/MtNSZD8R72B5TtQNymp0tVgoJhexTOXCUOjhq0RgiOH26aBkjDzlU
imUsGALqdyEqjRdRbP4YiWWNf+xAfPlshUMGaA0uGpx0tV/ZzVitdvPC9JZzl8nj3bTIbY3R3RbG
2qksb50x5wsw83LR/jWdsxBOdWEJbTmgd68Nsx/b5tIRjJRKx7dK82sHTckPdyzpAqojrlILR/tn
BZ50P/dDA8F9KGeVEIoXfFcyMqaNNKsm5MIJhE5LeAsWYQnbGq3SQHCJ6pccki/zAZHmqhsh9yEZ
oGRMqVbqpaOaMvG9kIEa5m2YvhN+spMwCNP4IOl4gAtrd8tWd5G2nrHiUcaEbIfNaLYV1r48u9nu
CFUs6+HpkKBZEb1h0n+LaneiI1zpgDAIvb/yejamaN9PnEU7n29ZNzZXRAiZMVJPBDBvRZAGX9cc
BX1w6+Nnqk1nHbs1PbYJvPtle+j1RZHO/fowxvWkfhBXqjLzVsjkacTed10KNGDryvShe1rLcUuX
wIepCdlLwtkgGnOOCHiOpou5wy/1rGAkFiAJyJ0I3Fj/fJBJWOsTYHoZqw3Eoc1qnGIQ/kPIKCY6
IYOFu16+5vnPcHXgK+iW1/8FjqoPyH1HbeFDUPFz+l+GPsKsc8X9nETpmb8c3S5bMLFOEfgutx9t
bZlKYN4AMQm3o9gFaN/L07pt4YBdcyRmvv5DWxIxq9/B/JpXvz9GDzkKOTfkE+8EOldXsjp1iUhV
gwegDZwTIv37oRJRrGksj35gB8vh3xbDAMM1TAXGUHimaGJnt/EZWBS/oJNxKCynSvGkrCdHkw9d
o0OtQ9xXDyOyEZ6SRjK6kkAHhAc9/x7vNDFJ2fQcYL/p+eFx3d654zHw9KWLRYVr29mYmfwC+kDY
5Hnf3DMzTkT4e+OU28mzsVENwHh6OkZWWroSfHuK1sD3NiJ3/6CUF/gocKP0WDC+Wg+8JJnYD9A0
P7ey9HOSt2mKOBVf5a+YhYaZ+ZuCSuD1P9KhK+zKt2ggmxrLlu/UqMgYaO+rffVOKdw+YUKK5xeR
MOgJ2cbTCUZVvC+grjaM1cTikvAFGbnEw1t+Rgnpq7IzbPGAEzsNEcqx8aYjIF+rhddZlRk/MmkX
21O9RDX9iN+D/rxGgNCgwwzDl2JgA3OdsuQwazY0jyGfQ5do8FmDkL3/KgSwRM2+F5/YdAgGXyCE
I3pR1eNLIKn0O/blPn7coQ6tyMO7oOLsg1eQY8v9URWFpj7yoyr6l/aFTHHr3WKoD+GSaKsuXC73
ZR2tYXJQNPTVkBWF5bRvl6gueFklTDZWDFusmqoL4rgUS57+7GvlKv3uXwF4hy7Y1UJpt0dlg3sk
zvRj7yvnAGbRfBGkYlukbgAP2jkBV1cSSSuDJmZouwHQJ17NpSgQb0fNPtnT5k2hAzlVZF3D5MX1
keHLAVJGRIR6QDj75LrKpT8ELWqWsqosKuJuMSu7We2z+cmW5LFKo2F1Ra3gqXFuug1LqAR3PmN1
XDpd36XCVfKz4qMoFZDb/jak2/QjD2Z7Msx+cKOd5Q3ljhLNKKjBDJlLoB5qIYamYACyChhOmqEc
w6wv5mbRwF/VL5RIUIZLUPmrz1EwXRVtMdmg2lUOT9Hnyod+CxWteWMAHAeKrXg99kAvI7tUfT4s
V4C9uC4aSp3Lk0poH2PMFwnoQ329Q5hp64ouM87PdJaN7ilkd28PpcZAQuEug9nqpbi3t3ZmS32l
cBRj3szsqI6oU7gMboSQuTSxLFyCCOlgGgsyfzPDYNFrMTZnxlXj8mh2kb9W+OLk35F5qlpia67T
sv8XFEGJVUByG65hTGLKWyn/oa0rLkUTnFwCuOCP0dlceUuFQ330rbK/XFuDUJdidErnZ/4vXjbI
Z9ffZUjFttt1QL7p8ijwxDjcxhKAysPAzy3BgyFf0DOifND33sSckvHzX6WrSPdfBSAnonrqrNtY
AXfXXISGXynjDHzJaVHPBGCA1DWLhTFJGBKJK5NsSdmkH5U4g9aDIo/a/7n8tsx8w3LmAV3A2IT6
MgEVE33ZE7kSwbGxB/zxcsUqxSoz9AyMIr6cI+brvcTUq0x4IJqq43uf5SGuQh6H7UbA7HEgcBFg
LavD48LOJUma+eoz+g6R4gpXJDmenscL3+91jc4wHK9zZrvmwmBEC9MMxIR95RYvefTPFV/dN04l
EF8vLVoj1Ai1Ugznjf1pKr2qcnGyF04gOpxnMX83FV4HuqsvzVJmxvUs4rK2Xg7D7JFfq8/Y8l+O
u4AuhwdHcJWfQRsQCtkzfUqLFNqTtUYEy7fcKvy2UTCvE72axKu7vHp6mWp2p+Rs4W9hiQ3+9ftG
3ntpQ1Q2kM3Dlw+uyKQhvJc0X13MMgWCugflWO3YC99KXUxWStuxZvn9PjHHhu09r0AWinf3scV6
zxQzgE5oPEKbsYhDnGt5+bhpvbyYguDXMu/U5TS+q75W1Rg+L00/hBINMqM1C1FL+TmfrXoFWqWx
ipOI08o5yslOsuLweeCL9snBqiP70braSl2OA44o2rrbkEPacksZlPSBXmaZsKxIS647asUNUFoT
GG3I/PHUb0EWKHHgWf31i5zO7rAyd4p39VfhB9X89kWZHEzsN4NLK/EQJK+m4iE7EHl3rMPwZ8W5
ejjggd/Ysy1I7FKGGCfeDDL8+CCiuo/c7Jm3GnD3XZ63ly5FZte0WM2CRxyY2LfBZVURUvgSYOeM
62zGho8AuEy+35MR5AIi5et7TOxSOShh0SU8er5hISUnloyrgA3c4i1fB2gLou9eJxItLx9UgJhg
vEzAZN1ro4b3ER/xF5DzYgd22xILKNAbrlnufq9ALqPL4otPJkh4H5/IB9u5IxvpCpPWNRKhWDb0
bBodX0vx6tCaoWuh/oKs5A20wksIyFSabKh1QmHNpQfSo+zcguq5hViG+Q75XJ8UkScH9zjklPR9
/66RmlNCFjEtCHdEfbJJmhZHZ3HqSc2XznkRNuQfuqM87CixVi6JU5RRG08E8RMXMjhf5pt6wviV
85gdhDw242FhpPy4vxDlYNiHJZCltg1A8g0mPUnW7mAIpTZhW/13exRHvfg7QTcgjjLrTCX/tQAy
Zk2Z2RFhOmfPiIqfxS29BNmydUbXrIRUrBT67SJb9L0MbGOqg0wD7N5xze/pODI46rWg58T5p5ty
NzvDGMIn8vCIt2MUIJ2GyDbdFCAm0dUj5ecjURYJavMAfCfAg6qEAlHoKk1jQWQYkF2LNG34/6Gs
+ALPeNEBBDhgWjiqi7X4n05ghUBEgBvMeuVe+7eeujOSJO025p2AjiRb19M0ll9mER3nt5eWLN5k
saAJ4Ax8cN6Go3GCrobfQQ9OXDTbZTseH9ByKEebfjjZvR384c79rvO/PpWBynXq021D09RGyVN9
J3Ucuq8P76nT9xCnI5QkxBVqPDcnez0a882cj/z5VOWH4vqrHZWxXNbD/LRZx+vRn2E2DztA+A7q
WEx8YpmrxS9FZ9gH0YIehhM/uqAa2tT2vGtcWolCtFC1jDW7lFO7eK6go/3Hhgka/De/5vpIUS/J
/TL4gjDjc3kfDu2cZkbhbeOBkf2uJrarMt8c06Spdhgv8dFQzvtgj2qN2TswJUVLlzDi7qlUKuFv
XeIS2Ja0QQTGhqzcM3BZFxLYyUaEbj6I48oz2KlB52CSl1aPsExfoXlI7YNLmpI5mElglLUoZkGg
Ns+bN+0xc3CPKsYvM9M0Nxj62LiIrWs1Km7N6/aIcmoTrAX2SKIWxGHh/yceNO7GfJBJ2VzUN57c
TKGaFWgRzbLUVFtq+R6wp27VKru8coLy1yo+4vKAYDcxVE2jlx56TcG5QGyAGExywjDEvIaEzfEH
jUmAWHyMM2N8CVcajd0cZQ0Ee7knfyJPy2ONoeKTp08IxmOSZ547M/xHQNo6TxIInGnTlWydUvyE
ysbVYe+G/T+OCjKp/jNUubzsYwy+PyuUKf2hn5VDz897Xk5kqFTTyT1vr+vnTpZS91WjuSQSu93H
KV27edeAjwkEfS9vdYw2/CeZcxMbqLJLbb71inqMj3j4iTTYl+BxNZL3UGS7UiLbUHp3BzujXinJ
uilCe9c4xX/JbNfE2/y9H5VeYAGZ8raFi0FwR0i6NGP+mhjA/QRW7oOj2FyMGZTRdPwh9uMn75lU
oapq9uYeRfsyCOcwyS7LTAQ6WF1hI8Qi3zYrFVrtwpQPkwtk4+1lPfN+tUzgdpD9hXNt4bb7trP5
04RckNMRFwYO0E5YeAEoFk1jmxLQtUt3r/uaDN0lAUgkDUEIJ1I5hHpLNwlkfOddT3GHosCkwob3
b1IKOkkHmLBydhCHtrEXnUlMtycJa+jIVlJ54hjmQ/wqXtADrIQkuymZStzmGY91SmaSGVB2odKo
9cxsTkEvTE/oN+5PQjbjcFCtVfBXGwdHYpO8fZ296RUIPrqB+bS2ugjTM3XuNrjTuveAiufU4r0Z
/s3v0Ov00mXuu/dGWmOfZCT0m07Kn/ytuVj868WFrtO1wtPvWdIKUuIVHuofd/l80k3tK8R6kRbQ
hxb2+ARXSzK1Swrs/8oTkFz8mTAC+nX/+5JC3BT0hiR4q8EabN3PDO0qIUIfVsMJBnzRQnjsebqY
WGogZIiVPVOUnJXLIxE356rpd/g/JF2DFT4jKDCxn7U3WdW8ZjrP0uNVC92Xh6A+Oxb/qU6300oa
ky3bFh2HXXgNV6URvZoGMW9/RJGsLbxibY/2xg0OtD4CgLyIaYrxjXZb+I47MV1qhzc0BUbKHC9v
QJKDRC3oKoHlKEPoBydl96/Jrohjjl7vmlusD+CWyhlpfGamNr5ctXRHVo9jcC1D7/JJuilV/uwQ
ZREGWeOkYeuRA+TvAWllCqaUBkQMcVuaDXqOMiCWqDzqWQTNmJT1+mdxSPY+gdseVWTlLtVQC5EZ
3uxr6ILtcYAyyStw8yg7dHq2KgYM5O56pQL4QJ6JxvzDiDEtQwMRnwJ1EcfGIhC8lEkOdx8Rsc3C
hW4fJy3Yf3iyGSZqAyJbYzv2RulS2SGJodROn2i0M6xvrFYan7Nn+zjwj6NdnXDu9yJlhdU8+Kmg
kpASy9iSMEZ4jmQxehy32txQv3lpBKVfrvM4GdsfrJCeySddL+rN8PGwVgaWAl/O2x5U+YDbs8gX
FCqNrQZwR969V72NCgcawyWzz9qBVvAGHld1W4Ykcs98IuC4pSTIAYvsAdI+tNtTPf7StDVKKAwW
ouwEPMHbTHHY+lehfyV3LxWBBus+SNN9GzpxLpJIaRYKUl12QBq5fCex0w9kcP77PO4VR2b7DcTu
4VAb4cRKv88qx5ArQBODH8eAgjb0CbLFFjgIvg9jbUE6NMiblSVXD1DgM48U7VNtNEUkNr7qRqyW
NlkD+6N4rZaK6WNo/dmpomh/87/y+0Tu3nFuIlcfQMQfJcRfrNTCI4LkgjDCo7VKi8or7Htl9W0H
srMh4aKHAs4tTXNcpmk6R3KwZmJJpW0YkVyKxMRKi9Ht3mdQojnZxpkEg9HdvpntzpU+R+qTeT8V
2TP4Hbc2NIxuA9cslIMe1jvzixZyGoi15nN3nbg5xUo0jdh/0NwSVwxw1j+v5rzjZA0JQcwylUCI
kYnM6Yqo1lRD2KA8HWGVT39IVLHLl2XF5KcVix533aa1TIPP9xdBrDbopRRKUfNfL1jWF85FQBU7
ypXhWODOrG7PXmHfeIF69qc5GelLNK7FI9C8mWFCnkusPcHLvJvXeWjjs+irGiJZYA/9yDoQt1Qz
GZGM0JImAvQzAjxHEwN7K4bUXcnni2nu3cKINbJkjAPzs4Eqk59OQVuBev5sSz4OMqJ8euHQ4vAQ
SGzUSIVIW3x88+zcJjXR2RrHl8uF58aQk7dFBJ4uxZrjjrkzhi9izh3bDaTY3Vm7I5q89B5irQdg
mjeFGFmeSvNSab0h3PIPVy15OtRubTq9jKBB2kVaapWGnatVbjjDPnPxjS3S93i3gIbueRHU+Z2x
NXwdBn0v6KrUToj4SJBIlqA0lSvUUR/2LNdbesQI9gVbST/C9IQNQWdwLng8gstvwCEPkdGRivkP
L/VChr3tJi9ZIpQ3Aea/f2iZGyMG/uXehm3xXN7jImLgYxXdrvY2sI2DZhC0j1BaIKwNQUM9+Ox0
VcFD98MSN2oEKjD3/cMkPhirqCGQH9Stxq07/c2iLtX9wA76zWaaxpraiJCRM9YoNW/cuI2lG1Xx
lby0IDTtaM+3JAReEY/+yb9HhYQuJHfrohtBkSDRJfKsTATLJ5poJ9/vCGwVqvgkiu7aAIDArtdM
5p5aomVYI8dpTFWWqqt8+cOo68Hzk6alxljJwjPp5c+Nohg/COCXSA1AJbwri4HVBOgBu0Y8mCOJ
7/aRw4mPRKygeGiM3f+5FOffz9yZQ8YrmXDd81jLjwbJPfLV62Htc6BIRvIubrazrnQhaArZ5zQW
+LXx4A3gRPubAa/mHQfWuNr487YiM66ezUuZAZhe2H3FPPB7aJl8+zODmuJm0u6+5HYEnEtOZ1H1
9lWo14B6kbiNMad1DUoAx9SxT73nl6NPC0eP0LHeBPNIjcwMwyPRxQ+M64x4R6VPww3phhxBYvR7
sSqNMETyLxpVww/fYBkSjc8elpAoIhZVimNSb7Ycm5rATmvsfHi1cUwVdUzSdscEhrbW/mLmVjhn
Z2Re9IyjixzAMCfgmfbUC2CKTe90+zhKiaSgKI08xst1bUlSmxTnlrRY9Now/+jTJ9DdCU9/K9Ev
38ghA+Eqy15KGXqRYoKLpXk4TXEf80vd2x3CUwHG8wcNXy2jFagd5sQGK2LkJk1frZ6KgwcMLSrM
63p2Ts6IqEKafLma77EItytBTU43g5HL+VkdmPbj9OqPigjFbyz7cybN7mzwYqbhar3zXQ/yzMG7
sMlG2GPVvpqcbkkBbzQ8e8zBQfNkEE0dOy+ZMsrrhsIlDwEfZ23Mb0WQZR8rJ3GogvdIckNS3xP7
/5lxejezhErwQMtKc2H3+ua+HKHw7SPFuIGXIekDA3W/aFner05nNjbp2kZfzKAU8YlTLWVMp/e+
u9Vm6qdLu2x+lk7oEegPqVbzKbNqVdiREFzqkY4Tou9w/NoOUVfx7iZFMb38mT+wfYXQk/vc6sKJ
VjWvEB7U3ChPvcGM5V7Gn0PZFUfJfa6WT0OuIvj2qTY/jOfVu/uLyxVRlykqtHs4xf3FYrquJamH
qGRRu4OeDpPM4Ytpuh7A1/39ScOg5lhzI2S5ANkpIeHjWpGr0+XQqhGiMSprt4GvC/uVX157gWVQ
Q0set+6DwNP/dRQkzeFM2Xd47RoACUn67ptqkqmrjVnJbZQGozR/WaqSBVaBJS6kFFYbygD4Hncj
TGdaGjKG1jVBFtwXa/zKL18+si4v0ijLKPA/RpLzLCLOfmrRQ1wyoaLDYz4nsPMCsftlNPkIzs68
3dqdJtOfRCNELhN82LqDDsTn8vvCyQPn+XdPpMxTKnCYsRtbqBuzTYRVGxLor0saKLk4ShSlPgy7
a82htg8DzudTQN31x0e07+B2cD7p72syLfhyVKp/zrU3xUiXcNsz1NewHIIhrENvkKbFa7te4TTA
8kGBOnpnRis817ft1Jg3efWGfBLBY4BralDFA6IkH2uG6zdvz52dV12DolfnxZ9EGIRD1QQVD4+z
sXQU9XtaOkk6QZjy4PE8iNocMnlRShecJmqZ74JuzgxVF7uQFU0Vtp8bFWn18R6UPt599LixbUKa
WjrE/VcD4g2Y7d6xx9W6Io+Odfpc9KyKy3o8MhRMG+4CXuKWxN5tiJkHzyaeLTNw+xJqvsmRO5/f
iZifwk7GaZ9vUgI+mJDSkSR4F/bb8Z66EBKF69KyngVm+7RBdM3ZsCOTomECky3QL3/83j7hukes
XXPGsspwiVjROZK71rDmvvXkSSkajxO79iZAQBXk+nkBCqxCTWoSiwLWNQ67nfJE7YIXvT1JKifX
sYCcRf9MXdyJKj0j/zN93yQ6SujGWQQn3YiwYW7oxRLeTU3Blpo5cf5pWtdQ7f2Y0Im4IBNzxDVj
sT8MrJWuobU2Uo3Mpjs/uOYIkPRw6+1JxH4GVF1je8D/7+TuKEObyTeD6EQkKcpCF16nFrf2l/L0
1OjZ02+uB0SpcSUDL82Z8uuGLEdneQKDABiyh506bAGiZi3xrDpSulcaHPF8ZTZG7D/uWo4LQcDY
REyGq+xY6u2YMSjsyOEEM1EJ20eFZ724arLqf7ZaxmRqjcH7B6q0NWdqoU5S8myWwIjCQlLIBEFq
X+gYlCw0RtsUvZQk8lpR9oW3SH9VnGujU/CLrOyT5xTPlNRfqDrkKqOUZ/JuYLcO84Iva9Jp0Lhx
IoM3Pc6JXfms2lDCW+7NzgvFpvaqOum3V8Fh3VDujREa/9gew3CMBk64wBUfFmNUkwF4Ymn5gpfi
9tfIJe0egqlrbcp8iRLwQFhdu+YOrR9A8iXBxaZkmPK+dp4R6mBm2ALN+U7PJhLMHCoEkREHl/gt
S9KV3QAGcNm3kL4hnFGx2eDGQ0wZ3ImNHOM/60jTq44xopsSIpPagASSE78Es9FdPkwbtOjOeEZN
lK/wl8BsF7P0CzFCE07TCxC1/6TSVkiOWCSId7wRQFSCj7CTS/YQpKQxGq4sgA9ZKEOey5rtcTKu
JcOmD01AqYjJ//kk+yG3ovwTCusp+vXZxDJ/z2CEdevRYXdSTSmCZ3WRrOOHoh4ezZf5G2lV4FdW
e+VqsuO1wzAyhzcedQiEbyJz4R6d+Qbx/4crr9HWBpUdD+2u2Dr8WLyAPr68L+tefwDMHJ7OJY63
10O5wULbz6zRYJgXGPkjaluBS1H9GU3T/0Epd4jWpT+Rcmq0l2+B5TvBxtLduV1UJrqtVVMZaLcY
1G2QOZE8/KXga53YNNubGpetgtFyWc2onuCibkHp2HS+Fl0+IcMAphX+P54tkTBhOVYvQTsbDiUT
DupiQqpptC6ACmbRSrjWEiTR6a9sOsBt9v1XF8Kles4QznWKonMP9ghEeJfiC5ab5vI9J/bou9/k
L86oqdFkDoSLi0pT1dj0Y7aK/H0yvoZfRIhi1Ar+K2ks/hSZi4yNRcKQvKkQmID21fD4iaB5KLhA
KJzvZK/GwPE8KGua//s0/BcCPYx/DpWtQobQlYI+zbOz023Nl5zmeVkP09SI5MlFILQYDiuT5VKa
5NFx1CaehIxP7+zQeqyJqGKqf9uw/uRstV8KnBDRuIuwA9wfs0MPPPK80aLcbHqgjFL3J3MgeT+O
KxbBQTJmgJrrAGknwAE5zEq5voTyhD2AEN0YL8FsuE7cd/XAnXjakctC6HswQsCabawnSST2wHqB
9EH2tIj/v7VKGOyIeOz+bGN9vStdkgeklq9ZN5tyrvX17FIsYgFJJ0ivt5Mwg8RxGR9qe/bPvrqa
pUWQ0KS4bzZ0AC8w9pYlhNmngyCHem4gZrdbEohug6pbWocRX575b5uOWBLC/SflPPCRn0E1V3Ub
NCxUAf20M4FlTln0R+BKvkKHJDPTHfYMA8xXra01PSA76SDkFpez6lCniNu6FD1QrAk5i8xsd8jv
W3TlzX2DR8kke7z1ofR7e6izmuGcGbFqTUajMC6LCKYdI/8HMfgemBoTJFVAdGYl2KC5B6bcCF/O
r9ZTxFMn+Yd/+MyMD3t1+jxvzZPP0uoa36OML84oyAKBRp8oI2Y2n2NolWQXf5zvp8y48ttW4v67
iZ+CbsyENbcp2hU0L5Dla+diCE2NPk6i+bU58I950P5vKbHn+xivwEX29ZPY/5MNKhQXxHP2+ZTQ
MpNTnqFWvJByIT3yQkhS6lL3e/CcWGqCSks+qmEtp5y2OtymNv/yKMxb/rAPIKHk+G2qZ9Ayb2ir
kNFM4BORIKuIuWpbVakAM6E0zMhp8+bdKosC+uv9fJEQvJBN/b5DGIc7Evc3jgRTtDW20nBFHV62
IoBZTgpppiigVLYQs7Mf9CbcwL9X4R4f+vpR5+uXZa1MNdWGJX91Ukjivbijk+ao5gGePzw1pm+q
JNmD5vPbKJW4pqX4VAtq+YontVBlTNSNsswA/P46I3J6OQ0YN4lrWhuSv2dgXESjH2kfrfcUC3uC
n2n6h3E+M8o7qa5BNNZpaaoaeEkHujBS0zU1l0JNfXc6zX65nRJMOAi7LJ24j9Rgf2z0it9HoVpJ
xIWF3Lp4CR9cC41xNJWCQK1ejR8sM/768lVJXoANp/Zbb8VzBDaAKINvqbFuqYsvmZWhO1uLL0Yr
wMGw+KYSSU8cG9Z7ZgYmvrPBC1A3bzn25HIuc+GW1+aIB8A+HEdR+ni4zrM381PQnw7ZtIguCQsG
Ms7pJ7v+fmyrYxgKnPYNp6Frx6tY3zDjJeXY6++BJWQMTh5bKM0wRxiUL4dV1SuTmmhSxCAOQ8eR
hb3r56GK2RRsojkleWJweMLYmanaBu+4vn0J4H3jVSmRvChi0ZkrDDWdt5kVoUMoOLKhrANZncX6
eE1i3O+zoX2G3VJ5KaMt489r3tmv+4qpdioX3vciVFeiLckuw56VVdSW9q31wMcNzo8hX1plLLtn
s0pVfycZUKAgbrmdfj/vl1lYBLTPrh4Gn+JDJzwwTu7M+b4Y+8VviXJjy3O8rBcDT7XI8OCIlPpU
YXLwgEWEmCbjnwKfwBXih8LNQneMgN29Bhtb8gmoJtq0VGEG7pfwCWKRPR6/Fk5RN7UbhFj9s1HY
Kq4QRwcagjByacsTIKcBCBj/WS5Wti/G+SLx+bxfH1k7AMJ5IpedVo1Qedil9ML39YCdsO+y0fRS
JCev9Ym58JspxJLbaFMGqvzcJsrboCpn7gc1PJiG1Yis275dt89KgbPuUPUKVsRCfKvU9HdGXIGa
q/+3BWyyzIo0v9akjvF0XzzeM4Nd8SrUHTT1Z0VPgMLBJZmctEKu6wMOr+C6AkP8T1WBOINIALMt
FxzNGUPUM0osNHg9Rx+GmZ6+OEyYVViWXz69wvHLS3wruhMt5Xt+3JYCY89DKnJj00aKC9X5Lxl7
syTvn6kk9PZrNZkIdmyf9QbJjjkqMc/uEUPX3Lju7zt+xyWq+KVrMCBSf4uap8zmZwWlAXGxIj2r
N4Gd+vgpGqrwc9l+7zBpadudSnXOMKGbhc1BOJT2LQYxNypy1FcuUfui5x4gaIe34dQMdhP6iNKx
4av/M1W4UVre60cXWAsDk+91OFC1YihcsmTAYUa9NhhLEt0dIaoKUl3wWKGvZjxftY44J7BUlJOk
r18xIw2OFM/YEAIWS3HNA6ajzkP9cBUONnXy5cdOpESKyF5dpOVM9HTJ1Jls7nJdhn1OjdZN8o/K
lF95Cy9x6oH62ibPWUX/l1ZiIYuTzsfsxiokRN08cu/B5hMjQ8uhBStHc6dumTxb9QGvb1Gh06eB
rI1aBI97ZYclJmtaw/j8OXyvSAMdLX8AEjeKtlyKJVxACy07rrVWmI85wAO/eyy8pyYTuH5kWFvO
bpv0ApAfNgKEAjffNLGWxxM7qFlSKQdP7vVnjoy7sSLm0WPGDAP98d8AUpr+lpir8pXRx1OdkS1A
MABD833W+ZTzCpFKPK4FhRDetQvWDyv5ChTXRb6WEN1CbBEKsQpd1Odfx3QZqfp55GeYWdrit1/z
r8+Y8U6vacNygmv+YzTWSzS8UYcwhC7SRGq8FJaaCF3m1euDI4ife+st+BYR1HZOhtK9qZEzdHZO
ji9NZqEEifgKdGKvDX1EfJ5aaYxhPWzcpMFe0KrcaWQ5yHQua90Eu/73Yyt9HPWhj4VEgce8I5mn
QWQQrQy8WkDRW1MV61SCcvcs0FyK0kWMwF3F8yGE8kEo6C/ftb0+ZVIdl7rSywDUhuft6XkaHrIQ
2DQKgMY+suJhVPLW9vc6HG2uglHNLenw3vTSSCB68oa3RruUQIAHSrx75jswJCciGBldP8n5AOL/
+6IEVKj6CTX241iaiMjR4l5FbCDWvRwmunVEP05N9nKcxQ6UCn93bMTkVofEefBjXSSSqj93AWfG
8tmKqZMvHFw0CmBrxlevkAGgR1xTgrzoZFFyBCtyEkhUFVJSLLPcVozIbgQrY6v0hQ52hPZT/Lzx
tqRZHqMsuxhExrfe8pBNBq2CGH671hjtcPibT2WQuTnwuikoDWEVGhB9+yt7feh+UR2IJYJG4UtD
szUO2PFPWI+/yDmS6KlUWqAe6VM=
`protect end_protected
