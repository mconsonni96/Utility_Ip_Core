`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
GfilFL5d0mf0yfSp+IvTJmJ4e7Z6brODYHewKjxgxY8B8UmN2vjN3eDescdh8YCgCk+BFLtR7zXn
hiUwqjw4/93TxXt2g4292HHhr+zufiw9KadF382Kq4jrK9WJEFzZZR1fH4MCNqkhxP0VkMElDd39
pqU5TY5rlk3kiY26KbLkp07OUImozH3tg2VRhil333FUuwCQFyYAp/jSvKN7rFHPlStfeYyz6n6N
YqVE50ws66aBpn2+RGbizWDjVFRZWZh41AVR8MRnUUV02w3GZKaYZF3NFtjI+oliQxPDVhbYtc3U
C3OnIzsSBNZsjg451RGGAMhAUsiUKkWkMQUtRg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="oLn/FkYtcvKyYCm6segMRqxmyxIj2B59HZMNpXlQ6vg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12368)
`protect data_block
LABNBnLd3yvjTSFQkx0gRAAjcdVDRsHdRKAv4xatpZuQZO3AiGvz9yWQ5Wv6z6xSQY0o6fBggEph
olOlP9a+eutkWF8R4K4WzC48kiMSw4qdR6CP6DrKtDhc5I1CAfHkLHCM5LlO704agNBRkKwnnYx+
i2K526nyv4Iq5k1XF5VUnUiVP5l94D4QHJRul6AACTZzRicwxIjSBKPNUoXtmtrfDM4UTRQEhZi7
Stq/i6Kx3FwCC1kH1oN0c4f4WAl8MjLE6gEdf6XfiLsPIC7EWwEkEQrhNXwwOmWSmuTJ+83DM3ep
nHB24HHSRWi8LPDGk671JDZpK4rRu+xhSo31QZoHX8pl+aOwK8KNJ861q+O/wXm4pYGaB1Ng4gzu
cE8LH0WkVAG5qLSaRONqiCjM+/v2/IKNUeQ29cHSnu98KhruhNjFZol/EH4qMszhabpGXkuoogky
Kb26YH5UJ1uD4+NpLAbuT2+mAvDyvi27cVEpfOWE1U4juAgRR76ONfZ5u+TWxPlNvQZ1AdIDcBQa
vf2UpjaFtGe9LMzr7zJj0SxzqTpcVVCQ+/vvfCKdHjW7VFjvi6n4ZvilyIk/e3YrA5QjPMI+zUS1
oTv4uprFitAj13655H+aWWZjTB0GAehyCoxuj6g4WiURSWN0H+j0hsRoeY9YfpeXXLPdDS0ywSls
e0lEF6XhHwlw0Wcyv2zSScs0huxG5fIr2kLGOn2c8aGuvJ7DS8zbloa3nVq1XCdzSoUyjMlom/ch
enbWKTASNRFIrVtLZ6QwE2pJnznvVYTjJxE4817UO/R03weNtqIcJ1AUvR/HCJINl9plFqgV6uJx
xvO9hBsYHCA4CX70OGooC43RLTf/LI1wz+F3WFzentigaNIWrkMnIza8NuG3VuG8y0BDKDmRPgnz
4OuTV+DJOxAyK9NYjtYGS/8HLAwtxcqnbUWJwGz0IYT+2DXpiybokvtJQA5WrptR9meVjJkJ/CaN
sysfInVBD8ke7JofZy1qOfWv3M0HDGda6ehCPRE6eg802gCcpzhpfgapqiCFqsncTZXcczJl/Izn
+KQDFkWdPcumTvVGcszUxUl9ptj5OB+/gNVugSi719fmLE4MPH3RrFNZ9LAOZ/X8fhdGQUzx9M3P
KCeenj8JsETW0JLb8gZ9maengy3ouGA9DtLPXln4fJudKZMu1q9uJIcpOezYEkcAfP8QzSWRD4in
WIYm5OB5JWzQyhm9cxiJJY8YVpqEqdgnSjHBOyT4XA9TZQGlzBMus363rLF9ZqvitjlFQJEfR2lO
wZzWg8NQ9Ua3X0auBuQA2CfwSD0Ogjj9eXWC76yTAfWsIgOw3u26rHoL/7k9vx0xtvJ/s5dsthuS
zhTUSoKNUtIyMpWLETHiA+jZnPv54khrqis1Sh5vfnasY+CEoSP/8yCX+vNxMgikYiR5q9xGVBdV
j1t7IuOiuSDPA1BDHjdq/GARQCGLS7EtGtCUrcfarRnjngrXD8fqr9JOTPPxfTsu9pkWbtNjl219
gNGjRCEFvMPNeKAJaGlax0IQ+IWX+iRGljDYW28GAe68OtsMmgbVN7ZPps+TzRsXuRmgj5nSpY4T
5M+YjJehcSuSZE5mpHZuuX75svPxtxFWYZrSWA7iwPeVBnT3ytPwxG88BJPRexJRArlGs81SVlbX
440yLvCyDeK4ipUD4yY7toDlT81RYV2e1DAfNHikZTc14AgCG/wiv+ikTmq2SCkqjCCRSER2Xg53
Jyo/Q1ne3jXZquo3xwgt0YIQu7KtRjZOjFFKU9sVlTbhJe/+iJzzo1AZyb7mapqy/6t2zcHY6WjL
emN5dBeJD5WIynUTKAUp6U4oe3rbwf/nIleNHrInKKjnvNXwoU147kzct7V59LiHsti8GhYvwPSy
8hWpFwm9VjEpX2gwgJBJ97O6JqBo7N+eFpqzPAqWAhP8JTR8iHJBRJyPfYhwu7uizIvK2iICWOiu
+449GuWBuo9vjI/xL8neO8yuX6aIw+6nRVpZjbkbPvZGbWvGIYaoSsgBGviaZhTomP4laVqKsVno
y6fdAeUApKMnm+kQd1+dRPpwQKBtaZaWZfcc0p2+mvD5NVrsQBc9Lx/3HnCaXs9Er/B7QtFNo3UG
hSUt94zMkqzRF50IZHHlu7yRcTlGyBQS0w/M1O5XU//63TPhd7gl66UvszcdXuhPP+QrOuT+EQz6
c5DncTrzhJYFM9ahl11m+Hka12bx7RylLnlIsbNw/f+TqZoeXfQ6s7HGrQKa0wa/JbdVJUw8LZ3G
JH274nkDq46WzD4bFIxmOe9Hn42g4fIYkfc2OUL82W9rL9Tv6b4n0DHybG3rv6StNlt5UkIXLZN4
jh7+Y16CR6wiPqoD68mU2asJRZLr85PTsVSOHwT46IN6wRszbX/3m30ou+wUWVhL5+OXNIQCE/fC
VTuAKU1vG84J26XY65FoWhvhPdt+vugHKawZoG8C4yl4JxYfoImQ2MOi9k7fokynhGmxOLHSbDoh
qWmEj7PR9e88I4+pICF/bEFAeIVAMwAT88nF3IZwPy+9XXpng8thFSvy9pAt6UqrSFqckg2qualU
H+5BC6J/ALp32sCcMqLrFzhWwrUa5Z6IH5sGTJGgBeoP5Y/M4UNX3kPwQ2+w6qOnuaO/th3HEJAX
9FOsAor7mFunOEP+n7UTylr4r4g1mo+g4HqBM8sgUdqfLo/QBSgHvKincBN4QpOHgXjEABUEiRlW
1Gb84pqg8g7zCjK2TaKfU1y4IiHR70IDBGYq06I5SlNS1ZQ+ekjyy2ZGTxeNcQdKTzHZ7jLw4LHb
/UHVJ6jh6iB3N07bz7iTj2wPgQqafOHF0EfbZqj+z7CGUcBqQdjtFad4f2XPn/3siLAtyMMtzCVS
bYPNQYrjIV0WuzlUbTOGuykCBTZQLBjCaCKQo9g7KbxnhS+qY4zHXqq2+cMpVbncR2x4VDvtg/5Q
mKTWAs0Qqd6VZezZl6j4GucnVhbhnE0QfICzm1WcRAu1KvjsehrvI5OT9uyYTz70jNoRzNWS5cBe
sq76Cqju+sy3xex4KrY3YmMsgOednPDNZgAxMtLNJ2UcMgWtOK9R/gX6SlPdiFxNoXP9jusrsKXg
iDzbTp+8LkIErEBCX65dg/BUYOLVRb0+MMUyEWHhe23Zmksu0V/EFPBsek7/5aBjcWF9spL2Iwv4
wKEnu7++bO4v0JI9cwMV11yrx1L4Bp3sg/kPbFKS36rjCD5MznBstJbNcO1AEW+TMe/3wkkITbU6
O0EzicEzrSKOtQ9qIjEEP8bcVoLhmJpjdQdCqj2BTRKa/307Jbzv+pVkqccW8skcdouIZ3Od9hwm
+A2XMx3gcS7ApPeKNLQSXjHGB5k9hVN+h8Pj2VfCj/IfSjU7m7sqal/EiDDZlf2SSmV/B4HTDl6R
c8mIqCLcmnKetSyeNegozPwFf2nATYtBM+fPxquE6qDZB2fB2W7jjDfmEgSfwAydEGqN/cadH/Za
+RIxNLOe4l5BS0KNY044vrO9y+svEfStgloHcIurUdAGGVT+ypa5MudrGYVugU8RMCLh8RqOSiFZ
BqXXaHa1r8balxHWYVvqi/pjwLHRTtvNGR/oT7DMBJsOS3xVtBTBJo24KqU6ARa0A+Qp5YQF97l5
S+KMYR47IA4HEWaFBPv/Ik4lkJnPIQloZN0oYh0oTlMg4QRm8HLc45iWJEpO3vAGNrUiwRLWVqgC
Z//uvqfjmgdLMOWT2zAHXissT5d4Xz7RjWWwS/se1REPiFYk0b2Va0JeJ+SNIPa5SVTPVlBAi+Pn
rrwf8TPTRxGoKfBsVPbtpLotAJZ1Jdvs2h2vRugXDQVYNuy4S9GUYfz08p/QJ7ia7gi47ivH7bdJ
+xbAbNa58uk7BxPAFdErIBarOXMMTWEFbz0nA3z+o00s+udlQ2luSYXGPquh5P+OTjT3B++QgSnX
Dt6z0mCYV4Pn4DXvaxePZLEQJ7pvtuym/eTq3wDcVg3ETFPvjW5Oxlejo5CYfmuiA31d7qqwuF/R
lFaySz4T8JYoHoWBEUE+dus5J42qCvKhJTxlC4JgFvF+L6WWVL3LpbIBzVnwqGiRl4ea47ZJf7+h
/NHKYVMD+wEMx5whB3nN+W5f1vamxER5KU/ig//2xOSNZ4Pd5sg1kOUGeB2Pu+UywFSeUlxOT6uu
LlgSBjf7Idxpq4xfgjG7ZRWyg8ZfvIenS+ah/UHFr+aEdkRm2izNKS8fKeCpFKfmm6+frAwQtPc7
WJMSlM9xWjHf+mw8+O5FD5642atyWqJlVNW0EPSMsh2+yj2PgucZtCrEb3Kj/lEWUpoD3k1fIoao
P/0JK+6Ceo6bh+HT03F+5MdJjbVsc2Ik1hMa/xHAX9FfQblGj2AWlELpBPhUzWa/6PbnH/Mamhd0
nxr379gaMMxkkqEnA51MJohq55lARo/8a+xmtkqsb+lc90uNVuoZVEQgej+NUzCNu0Wze1JogsFl
Cp6k9Waxmv20LZp1asAScUVj3yNcbE4cppkFLjhfBtRuSnqOKJUnRE/bcC1Wuacdv5rQ7A/U0Std
IPPLI2CedggxNYzoyiS5yb+8dEOKvdqIgF1b096rWnnD983lBOgT9DAh2lJDSDNJuToGrADQHDWQ
OEmXV4wOZXUQBF04EfjAk+dhP/aG+ZpQHclIPqC7enMJjXS6COyKTInt+6XxtSV8RJ/gSXp/zdiJ
OGGTAjuGEs71F7brCzH0sf/eF9wPbYtQ2Cjmi/tHg76Qjhw+7REHpmVkv9FC58NUGz5BDxav9+Ew
O0L28Uh5wiPzVYDyU6S1LPVvVOfZo56Na3UHWBfg8kWd5pG4N5qzMlkWF3vE1NJ0xMOYQUPJm7PT
cEWSViJ/uAbf90aJH9PosQijNv4d0mcWSIcEcqpgbd5d7X4HdV30suVJB1chTAa6euIVFI/yP+DQ
B9/Pq7rELC21F6xaNJCB+cxqhE5RGIYbG0WSCD84dHZZafM29i2oCsLDq2gM5lDGZmG3ORmG6p/D
hi3KLZX0cejSVhsZ+t5Mo03HvIBAVX7wF/QuKLH+uZMXBvbRzf6V0vRc6bHi2ZHmMsIK7j3jKPUh
2Wx/SkoEqlA4IXuH4+53v/catOz7yk+hg8RJ5cFRGxnfeswEsnpbxs04mNiiz+vgVcT+6sL+6chS
HMSMdVzCm3yujBHnrpxLyBStlJ+7g1u7PcJ+1Mjpv4GJGl/l9NZ5JVcyga3z4z42moYap5oV4FxC
ZYo5vPkKrlq/R9IcXyZ7HFMPm/d6OlgxLl4OeVb+5x0CRf33WoaYyoL+FyhndDhrMDgYh8Yh6SJU
qH8JO1akuNZuxaKA5Y5Be+AY9Om2mFnR+zuXOcToCA5o3iZOKh5kdw2nCX+8ZVGznfRIMk7vTzT+
HzVnZgzQxi74+23tT1iXaIXvX6vONaJeKUTftZXvWD3SbxgFnpL9AUQVUomMruyYlOnDC3fMvEXL
WN4OWmjeq1ve5zwUPPpaElzcnWjyZ/aNLa2kAp6Wkjnm+BT7/yBNE7GJqDLuBZ/k6ovPO9IggxZD
MWA/GM824yNXxw8Tce8HXkhh7mz3U9XGb66BruA49ktemAGj0ylPLYXaQKF7g4bprfOaKyUK9c6t
STcjGT0OfZahtHpwetnkScRSvQ9iEqTA4VnKkXgIGrIlKRwZ6yoTeFwVfiTS1dHDkTFKVFtB4817
xfoo+ayRgq1XUnSOrj0wQgs1CuszozL5TIxw7f7ud7k9HO2B6X6Iy3cApvgZKl06Kv7kGxl9FlPp
759mMLDtyfa24tecwUsV8JK93g2ALPcEL/miahUVmFtcxDE8s0MkfhuLKzBV8KR20vN0rlvrzOy6
0b+rBYSVntyVCB50QQ13QQOtsqldD16G/vw1E5xnDZx/PCoZBcTN30PRGt3V154iBu2Iab5pCLt0
hDeOJ+2W1BqqBqn91MaWMr5zS8lg0/prdpfln4Ntfc0qyaj9U93H2E8QCNTSIgRkhpaGaA6ijm8Z
BeW8OZYIbh6cPAa0UqHuKVzqc+aVr8Pdy8LLmfabZKu1Aj5sj3RxW0GGWdWqHAHTfbYQsJiimiKo
fFxGK+ibw3g6acXzIz0RbnTfYB/dEDu83//N0lqks7P1a4ILEi6qfAMyCAwuXdmkBMl6xiImYFGJ
oSCaU1mQzdDsSknbZlR/PJAR44/qzZCXGqwbPMSVQs2/tHEa/vMjeR875lbs9PQS1qBgQKAgBfyx
icN2lZ1y3JqYPdtnCxqc92da9yVEdR4Mdd2kY1YuxvzX6qbZM5rE5ZHhHYnyLRGkEfWtAE3f1fyy
Rk+diAs1HVIorDpkNF1LGu9vELv3vf/KVpOL7Vj/HB3O7l58VVeDnhZ6hGYLZvXhY/55ojE2kRii
2vd/orFa2u/fAwvIRC1Q0nbBvygbNQbuqTiTwlvJTohI3dgCuOLj7n+qP0Z5POwiWQxKJ1jafN/4
YnwIHz5W8QaJFoJHbjSMku02zkj2gyXa7EBsVz0zNeXTbM+kezwUn5jLuDshOWRHrDwiMqSRQLfr
z6hMlFgWsiXWB38J6sdHrkcr2N3TsOP5DVS0hwPDPdfQCBbtMdpCusJtNPBbfHCulkeut6jLtFlS
ZuoPAIybw8Uez1GERFJ+7tCLkifJ+E1LoS9a8zLVrlvzAWJh38bZYeWoUI1jr60HnVFqL+fQt/Ph
KXembnEve7WHhljrZacEggBfu7RouUeQpvR7OUzj25vLXAAymS3NkfWnFifv5Or+UtvWS8NJMQOH
G1EUmVbmwvr7YP9L5LixAywWv6gY5/DSiWMv9roIHXyBsb02TmgRx/LpjuGskR4SHcFI2zJUV+MW
jJIsRMYmo8itdNG6elq2Uvr7eokn79U8eXMwbw7ycZbkM7SJwHNDxFKHi2cYUxK/KH2dOJrzDenT
HefFiA+HAmpOxaPLAaF8xvryvWAxcOPaXRMOHou51r1PSUzQf5ULP4+HlfTsgkKG8yFNuPnI3E+T
cjxZj7aNK6H6ZHHRgVaNRSlBOCP+IurUL95bZEWPgZNCxObUmz0dw9xBY5r6fgmxN/EZNs9TW9fi
PUQjIuAFFMuOM9Q3RPPQpDroE/im7uVNesOt+VmHTbyF9NcjBz+CaNcfymyNyastV8u9ZaDPLpYH
81vRjMfH84TAx2yOUemf1HChCCgJrriL59igAMsav98eg5k94APkmCGJ2OHNBuutQTqTKPKv6Ecu
+qPl7mgyphjaIaJapLb+W+NU8ztPLiHCXjOb3uI/h0mTzfa4eQ1NcggwzA2x+qh+1zQflIVrNK0L
Q9K7VI5SLWxIUeo7jfW5hlzaUHQt5QMG7xN81M5gwdhBw1nlasI6tHt1Zxp8Mxc3I7alULZRfvRF
NLhMPrJxw+fmZ4YX5b5lmfjLMhHeZZ9tdtHgMTpAin0qUY0eFwLbJRNgdIr6euZ2cDKhd2mkqMtC
XG89NOLNIzEvU+Do1afcAz5Kh6VcQhvbntlyrmI2n9X05j1uo8MYYLnc/bOn2uXqyS4FGux4uq2n
WKeBOxYQMw/+FWPsYgUECQO2A849iQbEk57iECY25oJG+xBXw4Zsm9r5RGtUP53VH9+rAVkN/UfI
8ZnDmAROkEREqUdB999gn0KuQ99J5iJDQBviRX5awEz3PIj8jFS8gIju+2zyQYLCCSE0wzJKe0kB
CClp/EZtG7wiZAGldN3PvKqr6wEdqok5P6dPzWX9NEmvh1QZcihr2dAOfYmt5zpQc3C78683VNrS
8a/U9XiEr2t391AbLk6uMhbAkW1f2qFiXgoJzlq4/mPqAWHwo/w2xHHI0bboR6mqcqKBSoct52Te
FhiUSEz7KtjU6JVMyleJb3yrlS3Vx0DBHWKWV6KxU5eKkuPbpYkzX6/r2EGXymoRYSPP/nbddk7h
kTWeg8nmyY7osr9jpujT1r3s38RCava5sJ0W6uMlszeA6T85B/Rv+TrA9tROSAF7gV+G+gIy9AnO
s3ZQYV09cWmsb5CKYXl/Llkj9RXTZ3IRIytdze1L3i1uiGSWV9yLuC8T0H5gRJhGnEHudl7yQl9J
J0n9R8zne9GL5XnmZ9fxbKmrEKrV5t9VIkQaycnUiw5rtBLQUenyiH1buo3BqT5P2259TEWjw8xc
PNQxhBZUf2kiQ0D6VNdaAAed7bTpNB25lxHojr0ST7O9qhRHPiJ/bzBFtVsKmyZ4hG7rh/FeA/kS
bsNNsf2vwg8sRQSRqZrA+GDW2g2+7ZIazhDPuLZUlAoadDhRWwtfNA/2MK8RcxnePuMeNSkiqqIO
KGGrnKkxQL2wpTqOwPoVu901IuPsxKgJOUxi0gubQhVkBW4fKBwCjQEW2vPdS5IglP6vZWlkJE9H
csyRMali0dSyZihQXh/MDWhxaqMydsf7r0jr0PDah0vkVtpjwY+65F1WJtLQRjq6d5dk7yaEpr4q
cu7KaxkvNH+EUWWhIyZfHccdn26mo+yf4zUwz97f6hcEKLwG4ZoBK5hwKy4E8Bd0etkr0IR+ogPf
a3vocvBeLZMSqXZmipbHYxF9LTsdzUlRG7lb09eFEphJePjIbTYepnIDyf8zwJv384yWFj6W2Zrg
Qc403L1839tHQZcSgEdHhtAHQ7yLZJIvDQ7OtH8LjpIuUytvR2ZywKxNFujnlflNG+xDCsYyU2gB
A6Krr2g6tnBTcYESG4xrTN4kVwclARrfFZrX9/UZzFq2tEb71Csr1dNvYMCKcNKbRxhH9ulybLdu
kH1gr4LYWptzPcR+XGltYVl8HNoQo+RFKA+E3e7IyoDgdXEo/hu7QxE6BbKWujmMQcCztuTFh+19
kgGFg5ZiGPIdZUef/ihPLi3ab80GXSqqFC7jpJqU7ISp75ZScQFJhJ1N5KodnjlUrJ3AxGAf7z8W
3Z31sIZkqBhVC944fLGdEPPCQAYsiIY1uw4ET1ubIt2x+2o/TsyMolThYPhaqd9YF/PJasoWxeKR
jKZ8D6XRgGGOfNAD0xUvkkFDx8nt1smLUY/iy3JQ2grvEWwKUrhVMc7dmIlHNJKe2NMCDwy55SPk
ozazGMVhwonbHk5wDEBXgXrei6aj7os0y9kxTxzitAiglBF5oIH/wZW0FpY9wf+wLMIZUsds5V6q
4dIN/jq9ScUGpwIXScgYXvgthqjEMPMFX/83S3XpoRnqsW8BweMW4YJgJZhCAGYrDVO7jLCed7c0
9TDsclwmQOzLkVqW65OGe/CJjPzR2NXrHc5AMyodHoX6M7skU8+drsBYlMRvBlI5h92PDasowp4H
GV2ObKBhlhMGewIJd/zUBjF0Htu6UMcOR58CKieCcc2QKMVoyIMCS9x+AHzNKoQBvRoHajEgMh2p
G+8vitRVz90+kLOHouKVsb/0FeNGOlcAb+MUTTWZvE4Hx4oOZkI3W0Ae9q7jaBLZWJ8OTb6Qu/DZ
eNLBJLvL9EfCCC1F+infACodUDo7Uxtat0eSyjvEO0wqTL+FhHyP3dwCtH4khUXR+JsYz3/+DRM0
jYDLsn1mq87Yy+rNOuWp7di94lzW8xDtIT9T0n4DQiVO3C/i8UT5wix/vXMEt14wW7qNstlMMgPx
wvyB+lPOwKLH79hGaVdSg4Po/xgMx+FD6BZmrFb/F6S7bGPPEVycKHWg4ip3qIGymhbc8uQUJUwB
f5p2jo7ti9AxOA/CA+mnxQkPvrbhozFpA/d0pVxEjiGB8aqmZK/t7KrynYjMJ7AB1MGsoHSPAF23
XLSiuUqMm6J4Apz2TcS50hI8nTmSeRmZCSJ1NcSabZ0ECu+FLltpzl/Sw4Uj6/UIQHdMBCZc6J/J
OdJm9gGrIvUaNWEVMqAaQ/gc4veLYhkszpS0i5FbVpBqag9ZRwX83kbHDrSQzANi0RKxBzlTS4ma
EDjirWO0bLGnoF8uPpmSqfuRElZFEeU9VxwCN8qRGOx5/eJfa6gCb9V7L3KIkRSN9bg1bxqqN+i4
ksXGBPt/uFl7DIz8ZJCPYMwSixCtPfIEmQw3zkFOUb8TgiZFLnhVMjqh6q4uJ49rzRuTTkfh19Rz
nZmsDRkE2S7E5ikEXV9yhmeNRSy0yXuk4iH/75zVGfqa6U1W2m29bg7pkHR7Cqzxbk6JwhHq8bqk
sHF90/+eZKZTaREffKheP1RvmsZPxVNGuIoYHiPFyWBLdh6k2eCo6qt822GJf/WdVRcHKLAdNOcU
Ve4RYc4qB6K+pMCg6iC/CJXNkVBoP2oshn2C6qtiudvD4b03TqbmQWMp06ZfR0EoBDwAnw4jIzKm
/hzT9UsZQDSPAg8Ed59z/PMGhVvsS4oGko0k85l0hgp0EOnaTu8ln1Y5OtBmjCvtHQg38IevHjpi
1lYIshA0mTMNjI53NZKkLuXIaDJMPC7AiXdsEvqfuIAXmET85OB4Prg7pwN0Kf+8IAm7jbwF9Cli
SX2cyn/DhIq5d0e6RPCeONmDvw5D/AXBdcUtaOhUJ1/W1suT+leJjCZSUuCOzmoRK4nOn/nyW+9Z
jQqDqghwBKMb4cMiImKVB675nJNyTHIooWv+n5jlv3EWH8FUXuwxlI6LvFMaV1w8QqZRI8BzA6oP
ZlCvsVMowc0Lw8+YIAibHrW0ByCIN0pf0p9mShCTlsqspYJcRrSmwp5tyjgCWK3OBjcxk3gNSkRr
x6VvJeUw6P/lhjZFX1V7ccNuRuA9iZqodT6dhZu48ijILIjShpcv2BugB+LpucMN0dm7m50b8idr
QhNsHdiGLNmHD6iOQ5zmh0DEROFIL1QyLlVwTwMtA0jaurvLLksdvh2p5eKQuezP1zVuwdbQGQaH
/bcp4QNGB1s+2EzPVSAzmaNLvubViz0IECltoiPiLB2fwlsPPU+N4iq+RTwLT8Guu7VeCT8/mVaL
2hT9uWCXig6qusyHW2ufjcZOajkuwlcXgQKtNYW5Ae5WZ/r9GkhCcHYIhekUFxvL/OHKxmg7mViN
XVohjxpUEtRzK8eKVxLmDk9LOOD2fXvSPsEQDmNIpAmP4sfRGH0UkDhQ582MSOiQ2htVjTIAIwTO
FAjOoQugk/TaZsYzIQlnCcBzJtpidkV1Vp3Oxc5178Lexr5kBprldEp/uJptLFttYTmOWMq3ZVkI
DhgPkPL2qXjBzjW082vqk2LIrHHdzRQ70Yq3KVCtBd1Kls5uOyWePxnh2Pe27+QUmlz4rBPlT4E1
HFRJx/PZVGQjaBxcovTGwwowtTyhao1/T4FPbpG/JYKcXnpfu40AFWUJryvEpq7RXYJTs0ZV6z1x
geXgxk2ElP73//8MpNt/RYE7yI96Y//8wGNBMLdMTDpWDq5lhONU53/wK+ODV0nE/bPHZXYuWPmV
CK8r3ri1AmpS84K2PaDVHBzzvkvuVEU9IpnZWsgbqC9nrF5rWuEgjKDYQBNdLkZodhX45MlCCZX3
S50dL+73TzNFi6NJu3raDbEDva2QwqK8gETT5jD0+4dHVEMYGR2ISDlNPLpO9UWia1L8HA/EIZ5S
OA0CQuyZVfzw2OePINJEtVqE6hzU+QG6k6H76PdIIgX4frAAb4jE1zWMLu4scvp96teguhU850n3
vUFzyLt/5Eee3Qh0s8tGxc+g1DN8njyyhyjcsgp4L+JhcZ81sg8RBQffIo4Hz4CUWkavWJgjKbcJ
X/EZCEL7Qg4+Zb4O7VKhFD586NOWditrmE5qiW0aIozosCy7IPobY1kQAu3bXfCby37JpsHaTyq0
nIIQXh3O+jVqROijtKcNvJoCQ+vnbROhlPm6pYgUWFkK7ZwU2HKshC9Nsb1UIgoLN4pb3bUYrou9
1Sh2FdivSumiAJGMjWsC80uh5TKy2ViiTp1uOH26SxHmuG/c/OFhP3FQtNPmcSXN1rUqV+ABDpBm
Qrs4a1d/CY0ytUzwUOhjccA0nlzrQcjZIcnxr9a6JWiDctFrOTOr3lxShmGmQhV7LRUjp/F+tGgd
sCurUdtzGmm7zFXOGtEohrZm8PlxD6/1iA4Van4Q37CURRB9Ui8terL24P1O09dWL45sSGJLkDr2
agPmwS3HJ+BctHfP3MzCuFC4zOhitFVGVkrU9esrLM7RP8szpIfxKvUNVy+N4w6lhUVeJFvdqb+E
NQxtQ/hXfKzTna0XrRaIpBWXX1T6k4850SFx4wUbSxKm0C0uLTeEDg6ZYqYxJh+SuN2xyTmQO94g
PS1h5gURjccz9M3HiZ4lNGTlNnDLGRSndGBAzdNlXb8WcK967Wqpn11Fk1Kheml0o2bsXndaRDFL
pjFORhM5FHbz5iAotWh4J5HAP0IQBt9rU7Qv952DJ8Tq5peIq65xqmMCV6zGARX3sxCvZWAay5OV
wY6FOroOiDFA4yOCieCFT9mYz7jiMImr6O6fkAd8kU6aCZk2460GyqLKtsepqNazY0DJkfvd1yvT
7BI8Z+ihHlOrs79cisb8AnkYbS4aQ/xdDT2V6ZsTFplTVOXAxCgpf5+D+IIeUs1LnM/FWLZKKQCZ
/NWUpxDB6v3J+W9tg+UYkGY6uRnZMhB1qSRtX7FLeSpl6eIMcob7CuguekoTaQdU4e5cpN37Wbzo
DT5+soD+JhN8bs+lBQEr+Gl6kYQxNLxJIpe43zcSualmvmsaIDQNTB3mB5gPezEkmTgGyIPwVVFH
pk1XYyr/3G7wOjHpA7Ywv07+YI6DACcaX2JgNbxHMZ5PgbaoYIMSJYUp94/33+g6HD70sGCjCt0R
bAZ34YccjfadHY0vO5p6MQyPUlyB5BIHgW3sGWy2en3PkOMhFAx2+TDWpWma1E17uM+xTYNOqrKJ
UVnqDwWNVeTZIi3/wjWMA2W3+rmmNWv+/4ogcZXiCJetPbyjUIM8E+tG//VL3sCQXgE6650neEcu
lT8Bo5zgxw0i0QltTtiLdlmiw4xiYw11VFX4YaM/EVlsI/FHBDPMGob7BxgoZfABiew5WHvyFL2j
00jDbHKb/qPW3qQ4HYOnuA5x2IbXqQcHWqWDlWSSDw5Mq5FnXaTLommg2fErxdARrYUMvQXOVBY9
S/VhLQyUvWXDKKqUPLG4euoWUGN19W/noKL0FtTJ4bwrI2PKncHHuXzPTCYF0HFz1LxgfLnvZXpL
Tw7qWrJEW/GU2wTNQx8ktuTn7eR4KnZ4TH8jcoGTPKIvDhbYFmb43eXzRqADQaT7lgUqpXc3WmCw
2MrVRALZ38WRqJtINWZxEj84cDOkn3HwazMdQgoiE0qAuF0Cm1dUFaAYxaJZfpdOJK1SOqgVFPpe
wAFW2rPJKywACT8BoA/h0yCmyHIPduLtWqgND08gtbuz5qEbq3j8gkRxEZoZySde3ATDg1uO+C5E
yC9V3nvWl0TUDuyhDFt0AI5F2BCIkUwvTjlSc6er0TN2IYq8Qqa3vu1gv1WlI4Trh03eQxmUWUJx
OOQ9wkmfcNqCLHj1G8ECeDrGr21s49FMA+VoOQ7F/dSsS20JjrI/7tH3O6Bwxwkl6v+yhaPxLAFw
zQVc5SiJghtPhf8Nhb9ZmzegPAr0PWJu2CfBXcPfhIrwmVP+o1FqY+0hxHQBai2CxzxY3A5D1Rgd
uutl8ed/Fv8IppPODEl9U/gHgXXjhCqKcHvnmnYxmgguLwNyrqIHv1V/TXHVE7eCrbAZoNrfcaSi
vUBjzzlmnLXiMddS5iwyQjzQNPeSLEGFtV950I9VeshBn6C05QKX2NbKmdyYy0hPuln2f37FEJuH
VWh5TowjgA2QUmzXNBdatZYxLwHGROCELq1UPOY5acBJTgSJSyl81/vt985WXd+lyewzSR8Jgnae
qAqvtAtC17jZ8dTJju4/hfdHWUivrCAkEWW4r5mOTK/l6+O1Hj38ZHglNCgZeZyMwLJMOwZq+alC
aruZStVTZ8OAWPC0jvf9xn8ZeTyUNP7wtdbXIBKVt8jepIBVmbPO2kh6knixzwmJGue8nq4e9LQ8
lRMBeHkSdBGaRycpBtxwrzagQImEJ/ujSu+ko0TfJa7Wcumyo60eR2hOlVOPgWOvOzSjt8Z/kfma
0oXr3/HPw5nRdYyhB4pPCwKKtLe3MOb37sWxtJ/UBzd4DktmiRXbAByGsZSb6pEyT8fTSQIS/b6f
RwpcW5lCj2GFatb62aCMAleiouvrOJDIfGscjgCdbFPIlmYo7oWP/768LU6A2qLkz8zyBcVZIZpE
5qjnW3xueBKZXtLFr6baMqgRcJn3zWYUalL2qMg52wWanOQk710kEXsc/T5Xqh6QfyHxVN/e8llP
PwK80+0izTik8D5GJTyZlI8WvR0VXC8OyWnlnJFhe0/s39u6OKOYrNouMYd3nnyj9IBBJirW+64A
v1d//zQ0kCcK6ZPYb8LfBMm+5CCBz4mf5uLjKmTPBF7xYWfHjbenDQtpp6J7fz0XMXY7yYKWS7Tv
inZ885NWHpJPufJ/03FldVKdhpVnCiYADuh/qm3DSW/Kyr7eL02WN/Qa8EZfVJ0fEuY/mxqYiFIO
TS+foMbgQz9hsntMSO4WPMl+VbSPocSdz0yiK6bX3w6Ktod15BuzELPyH1i2S8SWCmox4K5FZ61O
988Yp4Rb3wd0fYJMxrZiF4BYr3UQ/1lHRJGO0nnMR4JsjLOoTWzVrtJXpuZR/tKK6AAeKKZ11aDY
5mSpcXadcnQAjr0iJu4W/m9Hwj13uIuVthXDWB2pbVUzW1/bRvjSy0bpSKVMKcl14z6da4GrmMSO
rsSk/ZWBroeKw4FyHpUA6W5HIFdxCkqYLZfWAdc7wjYrtoJOeVBAO9/z7clTWbOP3bOuyj/2wclA
G9ll1qgYx+m+O1ozEW+JjrWrbFP2lSVnsGefg+i2KTMDhVO/jY1ZH4UAUxmzXGUOl19/5Om//Rcd
xVmL+OKkA75aT8fvGcHDyOpelXJsMTlM9KKmEp/3rk0zsgJ5xAR9sdH0L7yU4GaJpgZQ+1FpXugC
GkTYIxXrQoJdOjBYaYGflFDkAOjw12917Q0H7yV3p/TAbBnub8+pIfNbSSR+ZZ38lXiGaMb2RmZQ
5qlzGWEbZL6gMTIciNczSbUzTi/smAHZJjrmJ+d8RIjaKrh9ty9aHTXFnD/HF1/AUH8JyLSeRuiJ
qrtRIyCY3HuAHoUIhEbaXQMcT7Z/rrtC9NKC7KjKg7So46zw6bPdHXtwGZOFCgsNPzqt0EJ5cgd6
n3RjWOxMvsmOGDupccL0UrbaC3L5GKGPMsK09L39xZd+Y4Z2jASrB70lihjAYWKrlq+d5Hm19tMD
z1DLlTVQWtzlq6RnJPulZKoqoKsKbVfyzop0Tw+7104hCUSags+CO8xk5QUaD5yPuoVbakekMBux
t/tTfDhIBk0mYCyU4TvSL76aQzvbWl4iRcOYzel0XMwTUqui4p951DIX4PHvXgKhOfswfjYpKnE0
Rr5NPPEZTOjYu7kJToqaLkDGcR6IFIZJDHZveiJdzQAv7JrBHLKy3WeIlcXiio9PWObLDSY41eSU
wCDAZKLUBkw4zKwyafpr4MnbI5uBvUgowcVsMn52E/40gw5mYsMLlU5Fnk9cWvsvYQsg/5yIPPDW
qsjcFaHQ/LWvWndGdox6QXDqeZBtpO5EOhwxy7f0iuSWNOrtreZGDFS71PV8OK/nh/N24VzSi6l6
2OVFGx3lQES4iJqua+daLroDKc7/0MFePktmNWwqtfGBwoOHJzhNbzKQo1HTeizyHh8Lb5COspBQ
cIDEZflfmJ2L8a4PubX4BS8BwmBXLUv2TSkpq3WozAHj05ItzwgrYrgdH9xdXKkB9lPuVqTPbVXp
/j9kKM3QKCMW/oa91grQQbhRIYgSyt7qC1azjCoNQkrfeV31bVeo5lc6pVugmQ4Dfa6MYuNaSfAI
xHeFuGLrRQbvELmM3jk7MDrzcDVz9iK0eWW9KHTt9ohIRJW8j7UnYjpc9LuxnBagQmPExnGNHS7b
ajHvDBg0uqCi7jzACnw8NFjWRH8JMPMlsJUtsXvENC4KmQ3TlPkZvu3Y+EK2HhbUlHnqAEOJA/8f
4kWOK5KfbkDDD7PEOkIgePNhGwMePn6NLHJms8jO6WqPeUWlJZLUgCoq6JKwbOg7u82hMGKpSfEm
nNNeFK+UyhIsnWLEuuaalQOTM8yxswwXj9iN9JApKMqH8Bs1NWAryOWRfYuJSndDpkPFIMQgxtW0
rwLrP8D9mIm99yOSQm/yrXVSnIWEExGD0YCyfF7SElHHX9doOXyo0ynXnphrLEqkIIXRJPZjyeg2
L8g5qqn9QT7j8lN1gQ4rOfim4mn/28FPVJWtB52Yvat7V2DxX9FrQ4W3QT/I1sStyrHBgWPeCPHp
IICIqt1CtfbvhorfQneLU8SqNwNF7IIhTZEB90pvXqZzJ5fut42sf007NS/1lT/M8T+PBVyadANJ
WnWtfnC2PcKUTaYCAPEf/eGQ3xNEe7vrM9ilCCnCnuDf4JbT2DSuZNF1IrEf0cdN6fVl6xyDj7eE
qq6AgU9Eh0fY+fpLK6Q1Gva3dpPBQCXU92lqFPh0Sx9o8PilXL21lhaCzZrJoVaGha5Jk6GMXq4=
`protect end_protected
