`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
W5FbZFBfjmumSRWMmtxmV4MkKeYXftqBAUaXg9Fa2rfWTbzT5iUkeyM3FkXKGP09frE51B0IKCeV
apElwG/dYuwcGbuvhoupW0bgbgXjSxsg01arCM7uw8EjxqmwfDjIlUkr5RiOC5seOoh9aDAi0tw3
6agdAEuoWgcSGSgbW7h4bQNYy6/PjvrIWVlg/Lw2WtUfAY6hhtnAWteu/D1UeY2ZIzHuL3ZcU9G7
uCsSTnmXjxGG9twSrMUiYnno+zxVXdRNHA7Bq4Mfn92dEwg3cv8oDg6mN3A5RHvS3DUoi+YuFy5U
cEK0x6SBZCqqFJAwWh4XLW8arhnGL7epU+cPCQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="6z2rrG4tTNyEQ8N3B1eJZM96nzRIPHfOk7xVU90z0xg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17168)
`protect data_block
ucrHRI/WiTKoOngATGNdBBRGeOl9zYhn2snIgKy3CiMFosjuYboDr0tZVbsbSLgU43S5v45GZHSI
YfPR4vkg7wqwyPkxuycu21HsdDHrglecaZtEg/KFGSc1De0Epa4ZN/Etm95BhI7ZqgE6rGMkV4fV
PT8cLyfUC5ASRESkvYNQXgqo2c9zI/THpAFGFbMCRVpo3ZmrBA1eUvTokUF2ttjL57W6zZ2mKpn4
JW0OvUHVxOQOxofsttBXcYM3dAoYb/imfnTP2H9xH7zjBxn7hpEVpk29gRj2+XCnlB4ahKKtOU6s
hDvZLWhsyMOTEPiTlTy1zS4V9shOE3qxvTzufDWQlbRPCRNaTmcyxB9Zx/N5L++wY2GFNUwo9WXf
2VQElzzmISxK3DTopTryoIz4QqOcFNyMOfpHeHpN5ybwmhsP6j/SM+8py0PDywL+Qcxlac+T1RHW
17MkxKp8yxMbqLfQeILetLEDDTqpwWwtKPyCtk3cyZ/9aB+vJ8MWgH9SKdGveVLjCW6mABQFFHo8
GLXfMURdYVcT6o8mfp5l0Pyi17arRasgBJ693kcMwP0wa6FhBEdBKrJsfEXabvzNvQbrYOrzLWN7
IlXKhfT3Iza/uIE61YY4MJqM3Zt+hMVCIq0wsAGo/kx1n2+sFt1Ht8RrwRkIwYV1Bi0myFWKmhDa
9p+NAdIyo7S5kalS6qyNTkHOmhham/XB+OyFhNoC59pyGP41MPSwzcu/Y1MerHhssRBVqy/l8vkl
n43IDUgHaHzCh1fVaScvRuzd1XQC6bNHFIhg8EA1rdGFj1D0PpUV2ohFaUiocfz83tauF4x5Y+gc
TPW2fuBEed3EUHQ0co57bhz/rGFCJzSyQJTyBmoDXKSQR7Rl5lPKh7ichZn7jIVL1C75qDSxNdhC
hTuB0upUJWVO2ERH8Ez12J+P6kFCZnJ7c31752Ayyzw8TashR3WG8rUIk4TsKJcoa0Vx03KUfdiv
JHMIHxHcTiFttNGItzljUo0mTHakwbZMmIukp7lbhc1geWZVndu2kkZEs/lkcxqqfT4g7OhqqyJI
SbEE8v2k/VGiF6iW1jju1407CTmme2VmbKCIA/vJc3tT3CR2Qc0pZ6fn9bGjl7oLIF50k6BkZR0o
TslKPakUtDW1v5rcqUWz0pV6CDR0ZhCvA/uqFu+eIWHFLkHzDhG7ldz6jIlG92pUHc1X8CDvUmiJ
iyn53nVCSb/aIPAcqUpymNfTJCDeydiC1vMj+2L8iZPJ7lzvKIem+KfJfjXNU4zTwv9eSgadbCP+
6KQLAHWdF6Co2Y7puNxgsNtI88paI0rt5IiQOQ9OKU/UHOtJP+hnAz+yFBD6w40NAZmU113Foco/
OBZVuFpk7ifHqR/jwNCwGM1oiwPvHo4orwsC2xnVadSqdYaIoNGagk3ETHFslRBliGZsrFRTBHVJ
/72upvyJOxB3Sd7k0NpNgK+O520ZuZkcV3SJ4Y9jfOxmsDzzWR1o9zlUIh2SdcFJCD7u0B9quaJe
Beho5Ql+U8PLI9U9XO7Pwv881YrU600rWIX40SoLUrRi93wCIIv2yjjJavCXtxp6Q3ViRKFD5Czq
O4afrhGeR3WukphezcA4GfzD2ICzOhHQDXsM+bjqWbFT/GRkxVXa14+5Ut445kPRyWXUlCk6SkOP
hoBBCQDlEMg077tVRh7nkPbiE7bZQ0aw2hM1XIZL47ZtN9E4cGoIxUwytb7y3iibnYs8KAGfuO6k
q9CqKDf/yTtInLrECpbgXEtDBQc2mcmFSRDFGOsYn+Dz4cc10XKILy+nIDGcM/I6iraClWPfE+YX
fo4pl09P/NnJyiVHBMqjBZvbdrXvfEG/dcWV48Jqe4ppw1dk6rZfszt47gOl2+hVI9l3LrnlE/FU
yuHIKZRqYE9Dgxx5/XQPhgJOf6Kg02v1q4vuyFxUhEpYp4X7PipFySO8XKMB5saFNBOuZ03HkmAo
5bMpVN/+OrpYKz+KIu0bdfEcv5XAI2W+/K9XX4TpOG5IIhMZtwptSfoWl6wEXsh0sLm/EvOU0m3O
9NPOxix7CU0ifs1ovbvuI30KBOCxsyEmySzn+Q7lSkr5wf50jXgOmEpdbZQOASrd55BWXS4qdt8v
NjDGIMxlKU3k75vP7VY9y0uzUlf6p8OUlulMMYnbD6XezVILn7nR86DR067Iow9dnGqZKoa8AIE5
XAvMO3bDs6TTBvUN6zLyh2OrejhUKeAGHNu9eC6CbLPUrrc2hr/tWXV638KUY/it++JTbzblxRIB
ScnxEHk4dvlD3O4ejPYiqQgDdyCBsHbKwBklAvrmJS0Mdth5+pb+weuZOGASji4/ms5OT8CAOU8U
POvv9I7FURzr5bXgKu5oVy84kgK1OzyQbUHhsmOQx3z6BWx9JMWhvWp506XyWbwXcu/L37+ob6XO
E4CZK1lG4Rgq8OMQ7zonJaHLV9rAGBkYCwhyjmL+G271OZdTXCuYtDWFwd/1WkORboIb9FX/L0Qb
k7KXB+lhgMNGnHkZSzL15I+DG4sw2yaO3KMF5eilOqyZsI6YpgHVYAGekGOE3x5IkUvYyQWJako3
5hocsaj1WVQcyPypuBEchPiuTr8bxXQl6SfcaXFGgtrzldqE8Uh21XqOtKne7JdjezyoSGqg/PRA
UKf4twOW9GO5Nov6BKdEntRfi60G4hreMi+0nXGb/yRgBBJI7tonE2y4xWe0vEv4BqrbPcYuB1e/
FFEt02n38Xe6RnJ2x83yfa+jLkt8KsfFWD6dZncJNFPmCCXtyoooiAJfdgBrgi1XDLG+unsMJ+x5
YmvLBI4MnfJ5fAihGBCD1F5geUUhbqkNSgkBOOTsqtn5NLT603SIKNxlC169BoUvIAlMddKFIcZJ
aziiIp4AaePm/4hnjh46sbVAaOZCIHbe8lBDxWfwKMciXxEyi6NsoC8QZestK3oxZXnTYySubfHi
06r7PCW3iep5xECfExvON+JacCmG2A/vEcWsEZCYRbvCLMxXh48xwV+Mi+RyfI+OEEbYkls5xMGp
12Z+bnNxA+DOmAmFV/y+x2VTeswdhnSQhILkjACfk7TZ3Yw7AEF9pja8nRV12OV8klt2r/tK0a8B
zzKCLnmoDXfCLjdPa0H+noDtr6LrCY86P+YarmlCKZP1yyLbFsD7cXTxckqyR6Do0NlHo4Km+M/I
HN7UpFxFCcbSE/jDYO1TLc58yqxXbEET0JODY1Eygt1HokWtY3uRLA66HyBcpGVURrtBFz5j4ZXW
bWaGStVcoVUp0IHj/ZvvtjmdR/+/nOOnFM/rIM1PZQAIY4wgXRXXRaMX7fxNMm170hbnYnP3Yjqc
hb6lc9YG8CRufLk3xhtBO9JqvOZqDPW2DCsYfBmm9j2EqV0YtQNI9EO/1NtUZglKHGM2Z+E92lPZ
5fG0d8LpR/IhUOi6AyQVzE8uMdJbUlV6l+lMpeJ9LJBJEBj9rt3j8IGHdimhi3qixOzn2mctGZS8
oMfst+74BbACSGlJdJFiKAl6bgmH43IqVxou257wyJWHyMtq6WR2t0vVE3FCKpv0yoo4Ii3WpD8W
eh4fmT+tveYftDR5plZrtClJKBZgG27hfnzGdGSyta3F8RaU2bIMeJrCvLtpSWXgVDAfHTWii3Jc
PVREWMGrmFxqjZIcBILmc1Lv10rt4i9NSxRNcK/XK4VWt0Z0CIyQS0IGGeo26SnpZ9q0jPhkJOaL
8PDgcrXMfGegbz6BAm+8J/s+yTFRkA3QncvJ917xBSJGBKs+YxrTAYInmFYqqcQqkfTfSbFHklVD
NYm+egCNI1tgicxDRa77HtJqJM+26BgVDlrdaNB9F2YJCGeXpIxmrY5GwrvFSOdlGHWEHZkUiDwk
kpSuWXd1XvhN+nZZ3SJV+NBHB+GGcXw07xs6DCVpwObf9j0YP8Djcot6p1C9alGlwGfSPuvbZQCb
mxVZwVsRP3mpscmeuYpoPyL/ZP+hzypmedJ+UcB4a8++kTNuma6gowECikfeSnIDDtGndkD3ZYhS
2bttoSuB1/R4ESouMqsPgVasSwjSpXDnm69QxB1hVlqumBKV0TgJHgl8w712oyfqCRu2XGUbBfZZ
6VvWACUx30COnKq7WUYTtElsTtC9XyGi+IwyrtNh9A/dKe1VAmMik7jQXo4sg5s6vkkHPhEsmNZq
Sns0Kb2K+E7peKM/IJkv16T3Ybpl27T4QsxiP5oZ+jLHGNRpRngJ6JUgDaA1Mh8RenjKoVA4gBwc
HzVl4MmIS8kZfLZ7kXknSv9HwH2F3P1TJ5PibZr5nKqxGPzvY+97EygnEeyTp7MmLUlCf1QunYhQ
U79dqU846W1o4Cd/dtnvOlvPP71O85ISnVt63uCF4J0JwmL3Cv10KAxzJAonoslJnZtDtKmBcHVF
9v6ZA50wM/oDMa5oOYuDLMg3MHYlvgmyROujQTImGf7LJRPiD60ISbz46u3/cBkO4JfzqLKsvNHB
5zU9Vcfxj2V2LXvMe+IHVT8yDQI/WwSZIoMnazid6sZqNVpNYDiYLWOD9C+Y0HA6YgJM48A8s281
VKNOHLY85l6OjBgGqHJ6hFgIpvU65/uxvRYiKtZ+5OJP2G+WvaWPTVCgS83RKn/H+9D8fLWuvHKr
CDbgrpe4f4sIA1USjTD0LuBZ+nTErZznRRMo7ZtKjgZk/+fwOzmhs7IJxDu5AWhzdOg2pd8uaxr2
Gq04+/EVbh5cah6DtXBLdRwTu+FNGkZ0ClkzwnIqsx93D6GmmgWt5gowgFVBgRc/2X0Po4ieJj7q
m4YmuZZiVLhDvRpqBRGWRi8/2ESvGDNmKgCIApxnZAnneBUXZguhTHB91Iaj1htk7iMX8nOX+lA2
qUEw5A/DXEnHnAiztBtbit+bEEi346YKG6RhqkwkT1Y0YGi8LYeQbzx+39l0alN6cHpjWn8ujm8E
AwuFbwMik2D5EyArFRCP+ApgT2Dwzg1S1TSHaJ6ePITI/FhFXj1KBXcAlX4oJHTr0Jb7wwnDle6h
Rrn3bYv1dWIUwCCy1Lwq6NZvL14VStGJ32hucdarFuCupVqj3Cw2DVKg57mzlXurSh8mrjOHYX1W
MCP5H4Nyrarw1Z+Sxg04RhNzCLJkOAW0NHpSge2jttLi9jECUqxphj1YYY9s9tFWgZxWtDQvSLY+
Ym8a7dvjBJBeY6XKGqcR0WjR7L2NBz3XqVevTV9LMgRDS7mY1oF56Y9SnmAD5x41Ou+3RqcQcbnC
OiQ/h2F8OlSjTNvibt1frEux41OxoJuznrvq73NkYitnBvVenv6v4t4yFPM72/3CgsOu7PJtnnfZ
OiG2GcTXDNPhptdUjYEFnFVS74VwfOVTWijnvFeYQkKM1s7LvlbvENAf5gHRiej/tI4FAtAp1w+L
sJ8xkX9y+F95PvoYNo+vccgL7je1xYL6ceREXzPDSXLEPZuW/gk/p/ZLgNogHSa811oxkhHJYg/J
mfX9p+OdpfdNBx7tLFrl+wpQ2JcTXDsGbQxbehsAT/s+qfgQeRWRDBw/VFtbiaTMZdDWgkrLxeIn
av3p0/Ew+FGtGsGE6Ez/JkljwyAQYQN9NQTEYCq1vAxWalt8Vdb6Wh24Wxv67CcRxu9Qt6pw15tk
8SqTQeL8mYQ038uzde1WXXpOzPP2nqAS/1nBA8snuUHfPOoR0rJJHKAbw4cPBNMFW3TFwXrekoT5
if/SE5SW8dh+xLqLQfaN4Zi6EeqLXeEU9XF+dR0nFHQjw2O/wjtrrPfG41EKrTwtazcGnRA0zADN
H0UxiXJW04uF0W1MwmD24u9EJ03LcHYcrs++JJyAC0DBOoc9mKI3SVZPOCD3YG0ShN0E159MLgwy
mOpjG1HhNn29Ml+V36D1Op7shzJ5q1++gdHmrK4JEiIvOLM+kKp+olnEbmmd8VbB40ZWhkOWGSb2
GcZYkOQMyItRMNep2eJhX6Xx+EF6exe8a1+YhdgLXTZrz+0d3KMNjMzweGjpjDVzaPNsfR+7JY1f
dlDo54c+J2tIcnxWgXsH1FZRqGh6RhSqp3zRFRtgX0omA7UrCnX3jy4rRkFKSgmxHKwIIGyi7V/O
vOarkc50P5h63D4eJsvuGpXH020ctFj/udJiIy5Umt1gzFEL5DApY0Zlw7eMcJbSF/yRyoOE2kBF
uwHZ6HqfcfLaE4x4XCeWiYb3wPm+VnE4pk1IACiBWFHhKAlxCnQjkS3oBKGc49tqcXCKirS19Kem
bNSdufV4fSPESBj52dHGtdV4quYYQR5XMSIJ0g7tqZDbdRR1Ioncy5uYeeUFqspOYUSnLa1IruNB
Jp8AnPWT/g2GEKG4ErePeUz5l/2dlKi2kQGmIRutqGSTK7mPot2Lyx0vGniSaonZYape/lRidxD3
caBqkcFgmXQLGRz2/VhLp3YOq2UAjM4fxFImfaqdSxnZ0Q73pfhQqEq4DTGyIq/qli4kvnQLZD1Y
Bcq5CRxyRWFtS8ll4EtSyM8deXZTcuC6BQnq/0X848tDQ6aEZxyAcEKVwr2aW/LZaEjd1Q9i+Pu2
POJzTjB26yvyLE463mR/V3vsc847RljrrJQVBB8phpBoGvXb93I17edehLunirlQVDP+BSm581gE
gZRuP4PD9ac4II/qywKKLEG6xrDx691NnyGVP4CLjTVum6yjZ5CCJKU2OgheQZBule6c16VXmYAd
y93ZO75k1lvnZg6vFrzOXOnh8GXkldTxeKWhTY9UEEKknsTczYmiCU2ed8K2thH/SrO8WT4QUoyS
Y9podc7MOx1GrrmkEzgs67riJ5LCFdm6ghDQoptdovND9XQNujW4CLaX2UHpxVtgnlByOWuPAwg6
SKtEWA5X+YFXOZk21qCec4pInk3/O6eIqh3bF6MXE9LcYPad3F8hXTDZrH45AP3Fwu5CHfaqH+KB
MXYPBbgA0nXnKsEi1AN1CWD2SRGZIUFrml/sCttZa0cZo2ganBekbQUm0UUN5EmQget/OeDNybxP
5ihXdr75wW6swpQ3khb34iKeLngCY3kspl87HK7tB9QQ5yVR8ElyGCoBXsPGGghXvy9jqB5PqZd8
aVqRN3YEVWK7NOvZ8CRQrG3kIovnSFK1MFvXUa9Zj99J0J4woeIlCTmZokMYiydXL7pF+/1Tyy42
8bTbqUama87s4MzfX0fmdI5eWkMEG8ihWvCiP0tVHQHm+ASpIEFkqvqm8IUHYlFBJB/UOJCxyDhh
pmCwQRfg3fUoQp0PaCR80AwjkNsdxl85x2HZfLfP5TmULE+/qbwBwRDbhGG1vZbrbbMvElfn1dxO
/gbThardidJ2qz3+ujsxg3BlvvnvvU98nSRHiz7Qd1D3h2kzMgEKS6Z4XwHLyJNU3nQ6R+z+ypX6
BDtOB+LqvUIyD15u86viXYw3wYmTHw5PzjbhuGcAeiU3JU+tn1/n4h0AeyTB9QMUE1cMLhfs0hSy
kTMjfaVWN8FtFzjtwWygrX3OuPCs4hVQ2S+HNTONSujwTuaEBS4ITlyucKx6f/iXUvKZ9iinvvBx
XiqyQiT8oiCBpyF7wxCOtozWO0THhoOzZIUXFgepzTwLrCI/ey61eBv7JKS3VlT9j4un+yNWmCUl
fwEqRyxtLS2noju2AGONwJnYsvNiIp+i5Xdz75aUe8qRj63K+obGj/6AYop1uAFaDF66/XApW1Ot
2kC2TTIwzE19Q6c0ORvPfEV/T+A2EvZx/Ku9MB5KNVxjM2/cvBohsv3ACQpHofvMXSILM9eSEq0R
oZV9HEOXQpljfZrd9UbP8QQkR3V9HmChRYoGQNnWdYTbS+QYdcFBhcx/jieetajNUzZgepLjHirP
lO1wkptNlrGRPsCcUQYZw0WZYafeRrL5N82/4UiwkYG9jAlCY+U87FOtfgoP4fnYirZNBTmq6Gkh
sH5K+Ga+rooBsU+GSbwmd5auyHyDnYgF6vV5A8f3Cbf3KJiHLrHcaEkEUbNLpWNpgDD1Q8A5YQqU
mq89G44tHUdhtJYhcfJ0cHKzX7+CeFxG1Ek/3Hw01K3dQIkoIPYyb3ASBfmRH2NnufUsef9BeeN7
j+Fb7tZZUaKE1jTeUbHGHx7+Qjaj6B11Zkt1AXHabvMJABeMyf25qNHyiSD7YmFIsCcmiGfCTLKC
wyz6sQGtpxbnOLoxEJzrrLqaZbQj07O6tZLCYDxrsSXxujp7vqqxhmztbju4mmXiZyHgoA4/C8rS
PMy7CB8cQX4SusRsVYMWbIAW9WijyLFaPxayFKsYXhizgys5U97CYlmJDg8NIKuEOr9OAi2IQxZj
i21KZS4Q7GWHRRwxs2V8FMKvMlkBP7y+f0ta519NLw3LXOflApysqQhu/DOiCeBT9qi0v7Y63MSl
Ol3LrOhvjB8Xg1RRq04iYm+3Kuj2pnywTZG4uLk4BL2l3ZfY3MbZhZPBcJDDbMJ5mQlgPbkG6SAg
pYKd3Zhs/DEYtePEZ8kYg8MLxBq4lVvWnlsEiZVyit4065rywjMfT4uFWJuvN3/dvcXN7B5JRMqD
5avwlLMdhPEyOyhWwjJPt1QFm0neE3Zz/1zVHM3+JhsqOzHxkwfh76er0nzKdlHnkhLiTGd2HQL9
Xl7Rw97jq4J04oz8RNp+wma4mE8U3r9DYxUYJLKnrmW6YO0vM1PpsOMpOZ9jWyY3LKM118lByGmF
E7bndOLxJ1s9nMKW8zmv7dVn7sq7NeN5XwlW0BvHc6kHOZQMsPvXxt7caikVT8m0pC0zkaLq9g/f
tygxaJRBsFDnfrhqNP8bzNRCC2+u+gPLgjeGxFiRk+bhSi0GtgHC/amzS1R+vjRvGx/tXEFviNnN
3WxEs1v5fCZ+rqMxq0StYuXcT2M8MN7GYFVOcImNLi3HOdaIARiLaa3bRDaCY6LUNSB1C1C3GGA7
nxr9faPtcx5lAOHddhTUW30we1dRuyPGrVHbLOUu4OCamw1OYGn3qnf1Z7albUQtk1d2DPWoaNyN
/7Mc4JVSLoW60CkV+dGxVGyf1Z0ISKwwK5jB64EVrHSTOjaJf0Cc1Vkr11ut/FsZf+MdugpOgn2F
fhJ+5oGK9pM9nNH10KLQRz90mtfTsE93OMvyOoa8YtwNA+WuzGtACKrLsbpHyaFJ1mNTwM/sYTY8
wTNWA53K0q+19Fw952/Gvd+MBRLF9mpBc79RlFR2FdO+XEW1ny1FUm5I21ynYbawgwQ5w6lf/Bff
uk4wrAD9mCvT66xgkeFuQ+sLzn/dVKg6y4S8ezzydZkCh8y9ky8QFVo44sPvIkBw+GsiDX19bMph
JRV06aHPdNV6659pwwRp0eZytwRwWV9BMvMYQIrYhF19H5ajnQJFJxo/9Dk6bjmp/9EZQHLnWbM5
ZrhglmiO4MaUX5tdX4ao0t4yXJCnd9RzjhSW00kXZ1Rexgv/Er6JzpqB3D5NE0/mPb4YnFLgUqo0
6PyMxPlsiTHr186Kzn7iBprBdJrCrp1l2KGMGCmjsb9x7dL2HbJMJ2qj9+DRAbMTPdgmJ4E2ysvW
gAkbuUJr2wd44uLLIyL2we2wlY1fqF88E4trsoJtrk/TWc9ZwPEWxMuKv27k7m1BSgo02hBQpfxF
RFXztWVl60bQc8HXTazVyop8ZIjhfN2Gbt9/NePDaDpyQka8ZZ9WtrKPxWW6b8oNY1kK4xUxvcxO
PZxv55bwSi6iJ9+pjIOlRDQwe1BbkbU8dRq6Qddz3ItdKBz3amaPMxpvifv+/6ku6JGBZcmt/tU0
oJvKZPk5ecMEqtKfenHFtrWvD5q4twoufF4pKbB8QsSuiVUWSOPmN5jP2x5hcceNNA7cxwW0yUeg
RXjtvu88ja0hHddPAKx7hJO5OSZdwOBv3SrhKPTvNMlW6FFa1oD5SrXG3ACcG+8YLSAVGVLdso1W
VpK6qkWfcsTb5nx2WXesCC03Zd1DVUncQogK8Py5fEQD1FbXwH2f5fnQ2kmZlohla/MdVCYR9EJG
9BTBZgnq5js7/ymS3RDuWePxgqzwr9/RMkimaHlvxtkFgCloEEwdUdtB8LmUtNjBBCsFXklqsxCa
cW0oQLefVE+vXLc8IEld9DggDmdb0d2o7NuAsUFP2VbSN7i42j7Xf392pMym09VQ0I9HjV4oPt3F
ADAeFLtDB5k1N7JxW9Jtm32GWk3UL8ZpN6lNXSlfoXNgX1QK0j/yEdd9SyinCJHmw9RFMFLI00oE
6LwbFBO+nE7tJ64ba19QvsdCtSQb+/KaDT9KwnIDEr6V6/j4/A2XJwJVbJCcxKBlgb3QFyt2aO+N
WP++6MEFwrApfyoTkPhTzfPzwy2hxx0NC5XyfQ9wTUlO0Nhb03vaCqopaZjzCdiUhOtp1KmwEb3c
DuJxHHbAtYljI/1jRPwCmWSC7DkIqLhV+Qb4wuEK0YLB0tZmiUOUeBVO83P1Y164xe7R7tbfLayX
2IBYq6Z/iEdp3bRujFLJy/5sbRwKa0xfQk7uv+w7Y4gtIjT7DyZXjJyp4ja4s1VdS5WXUjJPF2RR
dJ7C7vsQ0h1nqCP6HcTqmOwJBYHvPWrL6svBYzeQ7hrQoAiVDhJR7usuj5E+dmPIxCJfzCQpqoRa
B+vtNAvqGId94c3YZ6b8YhZGjPY2jrBdVvnjDPqc29rXPKPlWWIpCAxYO9qagIMiiLHylK21vPFW
rhcuD0pd8yHA5LNHtc11cVws0dMYcgJY1y6HxiYM6xM0wsUckxjhwdLCYv35z8nlkfHRaZFhXb1I
HWqkylWjZPVHcPQsJMtQR0VK7QGtMFPcMuzKbG6EBarx65cpc7aLNAwJiWP8otv/HpANNqD7m74g
QooLZgjIeMsiN18rZJ6iWtujFLMbSCCu521S0cNis/J27f/JkTFW/aRBWOtuOFgSRCCmiDcz+mv9
s2tXwILVk6LUHIdyXD5ZqYM/j80Nf+jsMebY22Q4eLhBaebqu1hq2lC6l0ioF75XSYicPNbwuoQ9
0ysCWKIqL5/CPFSKdiLjAbNAKo5LXgThklQ79YJsRjb8B1bZo1ozhrex/VIoHAgiZLBkRdJXVl7o
bz9/g8elpr4ZjO2SEaAWiu725v4uJcnOFl7a2BScVWesDovS2ViKwJMmMqSR/HtCsP4JkEFRgCzH
pHzffOc17kK8508ayWxExfXOF2NCOtJXVJmYv88PBtfctYnwSEo6n+IOtJDvKix/mVjYDZPMDTCj
DiUtyex70GJVaq1gzh0fqjuLk6Rfy8Ux3cXgHAC/7m8d9914iQfOmq1rCnQgVAnMyBHQUNU7y8u+
MYLJGT0EvBtjTILy2CuPywklyyKWr78aW/xWwTNkFMNnDwbKvPmwFfO0GAnreRN9EAR9S3a6978a
EovrYNqrfra2WyrMxfgmxZqnNfev8/Yg2ON5tF1ZZi225pxY7tpE3TnGLVkd3YjeY/cARqlWIHas
qJLps1AhD44/G2N6M9+mhHy3ID61Kj/QaMzA532l8RcojOT/jXUsB1wCxyHDKQlGQLtjSh2ZeVL5
Q3/d8je7mJ0u/i4Zk58xWVMixrBKpuSlVRyUaG8ciiTfdQzNGdxhzUK4C2u7GFE23IW3W7o9qciJ
hkqM8lc4ROPOAhXf7zirlsZeSiRejS0g50NCGlSusdO+MwMepmKhwZMKGVVZ637zQGLAS99abQJj
7VBhnS0sU+vvQO/HjkB+NM0v9pMJIEjBsCM9lu5CUHYAYOGHAWonsTL69jJX8x+7m5uqpRGST5T9
0sXcC1AQDCOVcehujWbJneTNGUqeyBqYJWuPxWsGBPg5Pw8671TqTOM+zHokQG9KChe9rbT/3OTC
wGx6mLRexkuprnNQvgiJ0ocGacHmmIjxIUVaJNaraSf/eZ+FzyEIT0wVXuNWrs7wdIOUfIuEeoHL
U/HJj82CE3+HInZKPd0FZYkz5/A8uA+7fpKfi5xTmtZ7qbiQTxlLRcYqfiAmnlfd7fjs9eK+fWVL
5t/Oe2OtDfSx63gJuNX/GNCX7mxcxnfxkMYYiLoVMIbkz0EciiAo9yn07C46Bm9ikyx0dvKTYQNo
GI0cBD/5iGNl+n/DtlfUvzp9DJZSrRwk1bMWdK7NRciI/eWAcfFxQbixvtC2E+Ee1kIwRYBENdQk
vZ9JeinKrBBr+yA3XF0hf6qlzlOhGrwrTHq3JSRMo0D7KHakfa6gQPsi1QveNtgR6mI+PudRxxr/
mdiMh8J/Kv4mN60LlWVn2q2zw4+9ptsbKy2EL9ZPahGAQqttzYAsPXQG0wyiEsWc5oOdAmbRq3Z8
iXbszOiFqojXp3Gdo0bbaUo3VjDvBrOy/hMv/1IJZ8BOJQqOwDMNzj9gut6bvRCMKBJx+bVFkBeJ
MRSBbu55mTYXXbcQx7PUb7v86EGMxCWrydtc1NfR9dJZtpNPCBa5KgmkM5So/Man/+kN/ct127Ne
SO20Hmly8XkficoqPrU8Dd+ZwE9TttGLV67c4cQGHKO1+IC4jQnQt5cdC1XT60H7BxSLYM9ik/TH
6olImrU/nkz6+xVeztzP3G1F8VsA8d2YXLrE67bxtwOsgsZhAC8NOCcMH3EizSMWE9giPCsTQqTV
KVd6LOItJoFwqN04SgFbacYimvhjhzMxYEKCa0O9xJu5zS5BCpqqaYPaT2om6Jwu6g+EgJkPPdVP
STor1LnITIA6gXuON3uU8dsCQHORs9Icw1wZV8YviSGswdLIX81vIap6XdYEFAn/5V/0FwzWewRd
M4sk/wkdb7BGH+RpQSWkj2LI+LQo52uxywRWYBM5lPfo15c+koH8Xgu5lBbeAX4JdCrUn3mH1zRV
UDhj5RbIyuSWhEFex3+Tj6+IXLtLB/3ga16GFOfeDSxU2LNA2eJLfwQoEDkZOpGkfcwsLuKjz6jm
uEk0a6zzRbIUGGvTEx8pJNPLg1UMftE49mYt9GpNmFSjDMqdIlsUKX9mf1158pzFo9qIh3CKxfQM
+eQOd0cRXGLusPu8Pl+K6A8Y4WP9N1PJQhs5lf7Zkn2RFLOI7HyNPeHmxrO+aHH9zcx9GCPonvJe
zy/e3TzvC8qC7NhPIXsdW7Qxsil2mfH+iMLa3Wv9pWghiozYSc91eWVeAGxXx/8Txb7N98plcIOi
zAdcr5BXR7Z6PptVbHSIbHDbWxUry/EsINOdtqS4z5B+VWgpd6gQsMsWIAkp/w5H+LWZ1bH3uJ89
z1udaSZR/oKOESgBayqXCzgV2LavodUln/3aBzN9GCuu3IH3iGwvqk5fbh+UjUg/+xClVNxtqbEB
s2Yyxaj2YVQuvDuSJ/GwXqTvMPFQa5K7vFcpW3Un2AKt1g4On0OxQ6NNjqb+aSwdfgGG+dEFGjwI
Vx9Xd5hZMpf+dQpS7T+57xrFgd5Fvu6Awe12hpSwj/Ny1blls/kbEUuG0Gu3Bs90ZAPkukJhZPwt
+WLS7Acjz2PRtK+DpOejRGVfaUtEZ0DmUkMIxK8XkB/IJZFLfqzZQm8mu1C+G/UbrVHIsBc94QvB
p2xz74alQO62QGMkLd+43z69/ViTQrXsAtjkyvq9spr4nqU/YBt1MHkBok1dpqta55UONshvdK9q
kB8hJDO3o64Kmc0ZCzfFp5Cb5LPWvqQ1Pl/zPQS0grdZ2HwzBc5lAwkffWl5H6L9pZMhSIDnJpnC
QDpY+hTtScR0hGM7MKvm1F1hLXktqe1oS07Wbo0bxLTr3UdpbRK352glf6mvi8j4zhqwhaLPpCPv
agO7dgMRoTxzsSBn//i5LbFGtmWeZ/JJkhSMWpM2y20Xs8sR5Mvp/vrd/EC1YytdJJ8L9g/QlO/m
Vr5z5Y6/+LHDogs6yiWLRSAuONs9qkR+2mEg8hLJ0gWXS043XSpy1mxO+h8vYNAohT4VWlD4Q4zT
vFYqt10NiZEManZsOwtls49Cx2m7Zbd7+gFuvupquoNf4BJ1UV5pyrJpRtuWbI5y0whQJQV8TB/h
CGWkuVHYrad4FH2/IsRYbfTxt5k1nsVWe/AouOfyrK/bfiZay5qNUegoRils/vP/26QpSGBz/H57
xdZGPb5gMXUJezHOIttaZJOLDJRYHIG7xHDJZ/iN8a5CNa3U6jeRdVltV90036v+/1ZOZ34CNsUf
SrFIhRR4UKxwRLOxHEngdlrVe+7VvdwHEbRtMVSUOKGtPZ1UqHnXcLwkM3BYhRKrP2r9ZW+Vx0YU
6rQxUeDNGrmnRLkFlSDyJp0yuwypUxeXdxYPZAowfCvirntm6+xUBWF1OLwXFioA0nXEt07K38jn
srqg99ECvYe3/TgPKkqZMc181p+idfG8uv4I72dDJiOjP/Y1tn4uDr6aMgYSJbDtqOZyEaqaoF4A
txQTHo1Ut8PB47HzNbFRynnVsDxPR/yuwXqkjBp+pYLiHF2W/+A2PCIjOFk86iZgNgQFk7410aWr
7N2oXc8z1noLStgmkIuDdzZpfIun6Gi5hdIgi3JwVS6osr9bs0uexGRXgSUr/RQv3ei5vfxT1FoD
Ik/PP9Hiy2cFXo6RImlbS+uLyvmu7tMWFQy0qiPu7aQAyyhGzlpfInZyJ+mpPaMKntQZqaS/AZmx
IEIYBCWn8dHFTGKGfAFsPiineWJ2pZn2rMH/KilOmj+GRedC4pZVoLPbhE9uP6SN/37GTb2PM800
oXl3psRPaYA/OqD0e+s8r3bneWMDmaGB8+j5ATWMpZMfp4FMtutKvYsOhvVFYqPufP8t/xqPJcq5
vO/2PeIj+EKdy5E8ZsMVUxTQ5T+gmui5JAM74OxLaGZGXhgmx3OLFxNhWnzV3cPuH+QTxMlCVO6s
vpV5DxwpSGlrprXqgbLB+YWNEVgrPYsObsetna1+yfdFnjihKHQGAi33DydBLkfoqJWqAbRHabGa
r/9eq0gIZxKyo5HdtBTOYMGAG/4w9P03Y2JLY1A9znP62p5erPcNo4+RQkT8cqvRe60CIfK2pQVy
5ZiXxnYSwjaFf02Sz8bGP1GXz2PYWthkjL9ljGpEIKYnLwuDMIBtZTG5RzkgHp9AqBkD1AGTDuqs
IDyeXDvstguPQTwcyrcfnFNJH/lkzUbYGo3a7KU4hKNvv1MBG2wMzNtQNE38JUdDkKeRlB62spYO
+DAdpigAnQ+ILaWEZnfgXeTkcujfq4W08iM2FykrWb/60AlEDfk4ye0czLYTGNBiXvd8xWMNRsOL
6l1Prit4Hpacbq8v/sX9yaApZjlf/ShKJlF7vJPp0MO3/yc9UpPnj6sA8ISPCfztyLptBcVIsEdr
yCFoIZUO2jTjYizOX3NZFnVt2ZhymOR1FS0FnS82KYAq5+SSPHH1WAqY2/sIznvD0S4kEvIQ5h1h
mdoGNt3MO3oe7wXFvptpOwTWQ0dkecGBFYWhXekLN+9PPG4eqbQJMYBncZ59eN/iLNanl+RsdFAo
suHpJrpRoqythRdqY4ar5aD8VfcqKBSn7LHnk9wlQYytHjdsp+918+dcMI34Of+cUr2YlaLieDht
icdXcjicEiNyfxAZgcmSergERoBsboE+OZewi62DAFPBIi97/N7Ya6x9acy070jolb+u0Z9uYG2Y
hJ0CeDny/Ov7B5LtE3niK/7kItcSO5rLxASQeb2VCTgRx1WDCsmIHC0Z35yD2Qr5y+2Xa9Dufe36
XzjMCeAcA9iYELnwaO0cln60L4/f4iMvppL1ocpmBEHwLvcD9GRYq5mVZlxrolwdMq3fRbQEPc/f
RpoZ8d8RmGiKZpGUmxqEfqoFMVfGscHwqGLi27L1IA4pQpa1LV8cudf7HQ5VkgeGiqCog7semjAY
8jlelJzBh2Eayxpo4D7GAbAfvB7x4ZdPdtWIyQEsyiOEAzh1P51Fq8j23OwxLbO8C3lCDkXFdU5F
Nprsr6USzZud4M4SCB68Nr09SMcIPagHxnLWcRNc8VqWOmWkcbhGoNW+JWpWJmjyKcJE9CkGwe+T
SFuEipZ4YKHemcisEiRo3vz2D5+IGu0u8cgvGLm7LteavKOO5FSioxFA4vtaO4cdhaTPnuYDVFgn
bLAlmq0yIy/f5kHHdJr664Vy3JKQSezq77Q5yh/p9foCD+QPrtMlM2nqKEUuRmY4NcER6WT7O480
DBnBWE0rOVx2PYJneUemHlroA6dN92pwt4NnrgpzKFsqFbRqif8pvcEdOlop9shjbDT8fgXssHtY
W3DgSoczlo0V7mD46NHxbjJGov1VilesWBWq4CFsRlutNngQQ4Ij5ozmiiDe9Ez4iPmBJsWkcgog
bQ5yUqcAozEH+YMfdkiUm3Uz2bU7c09E3Owj1FMYq2V6NIIn6DsT3XTDPu17N3gxKJTYfVUwAGbs
g6lJ4M/tnHmPKPqPG8b7HnT9nowDLknLWk468Fx37WtG14M6/f0DTGJ2U/ciIODHJk5FYYhjZY61
O24I7c2Kkhd0LsXMpL0pi75ZREZgsYqukXkRCKpCk/KavDPyA3XG4EnAHPeX+kRqFUDcbWob81Xf
a1ABlYU6PYl2aJCXiPl4nWFwvm8gung0MMWUKkaBVAqKteavTfmK8VEJHMvdhTmrW4ok7tUJHc8w
bYnp8Jk2uvdAjoko2BEntjbl/8N7cBREzUczke2ClhbqiLlXtUyFPccsG66uky3V3LnqawGdTvF8
XvIBX4B8XDcQzBUFc2N+XF4zUjA+7bg3RmB5flXMHFZC4mJb7gYFZ8uP/029RA0MWdONcipA9wcH
jyaW/je4ym/Qk1f1A9xRvSqnSfRqfigTr2Cf/TR4o+1UccjjNPBivQ14oD8Ne/he3VEzdey2PzRr
lsD1APxhuRCD2UNda0vXTVsUsoFLd/E80G1a+/MY2MOgXEoAX9QhZNWJ4GdriylrVLN1HpjW1vGi
Q/vPy7/j3fECYfMD8W35QNxwyZRBc0i/AnyPzHLNWyLMucd7Majg5PSRteKHKA49oRMHM1UrRQn1
KZG8qcvmsd1+2pe4xaVpgVxZSv64DG06NTre0HRnJgriu6YaoxQfkJ9OA2/MNAyY4ulWEt1hgcNP
IE3QxzVZm9ADWS4fTnxCIzakjR42KqTQYZ8ZVbUTaIL9FqR0d6fZsiQ731Hd7PELhFmLO7aA60wF
tcvUDkTp2sfmfqZnBBCniqJsxdx9Ox7j0Mr8JRrsZ3oVhzlNvygb7tWSIEx5Jrx/fqqBzjH0L8ZT
82HZhiUUkGevwAKrH8FmahqXDVOLHezBr8+yf7HYLAbVWhAWz8HxwQHWbsiF52m1fAQyco82KXQJ
TBE8XmHtyroNCU7J5aDONjZyR2mWQTdNGcskQ518a3/XQyntWs4W2GsrDoW3ECN+9cDcdl/sHrz6
E/JlO+NeA6I1v1Me+8FUZxwueoe9N9oqcU/uWxFdhZZDZTgz+fZYGOnBjGAZam4hIn5SQOfwEW42
Le0bvY05Dl5kKwQgrgx/9nyKnzX3gTZatXakwHZyz99sRjIMyoVvGZWNg3fLzPJe8c0bwcPXJet0
YpXutD0zOv70oK/NkhpTjY0a5ewotbtstJuhtkqpGDGha38nWwglHwKhzgxrlT9Wr7gZ2pjYk4Os
zky0hLYOmB1Wn0Verd5VHoxSnN98P57BjUUfRqcjn7xp+KJ9L7xmfveTvUfiLse+EJgEN+q+hyoE
m+D/bAkjQn10ApAVVwwBD53XbtASH9vDQot2c+NSQMBokORZjYlGykOlxmCa1uW813p/W0nlE1jU
Jl8hlUBHhT+OAcuZ+YZobHmZfV48RgARnuT+67fVSeyJg8AW3N78+1uQEIJo4LdglCWRKrHSPQQX
r3SUBI4JSDhZmIUmzvPwMrzhAtI3GeK+P6e6uey8SLTAqwEs7V+cJE0XDZu5CEqpM7YZZlNTDw7w
vcPNSE8w67ggPOMrqvShqQJcLMQgS/O2ja86LsKQzvXtcPZx4c8ELGNZoH3PzQFtR7zIlJK32kBT
BOvkVTHRGd/wQszcXYQplEJs1eNGG36Vj0zwzVgUmTmz6lpU3U0YoAPi7GoeKm6AwVa3OLWbsK0B
G+a4piFCjFd9onhCaxi1rfXUfoq1xa0bs5eKU+Zv/KLWFGzziHG1LJD5xlLP4csKDSbkXNk54KHV
PZSSEt/pUWrByFTY/BaCiTTOtnpaehE7zjhbKxWxuU7bY51yEHOzOHv7S6kjF5MoI/gWuVcZONZm
SjiUqvCqpt9XDXkOz1AXXbXE0S/lcstU/AirMOPFodAZI9ty0zu5Px9s0Fg015rKKKC21boVgPUY
jnEXJxNlhr9d1ps9ZmWjkEnQ5Y+bnlZwlGEdL9Yg7VImlg9Bop96jybl5V+SAXz48MG43NSQw1GX
nh4fWSH408OLObmJ+WiPoC7FQ3LP4OMCwCKy4l6cNAmWSTgYv98Sk92+WEOvlbCuBLM+bilt/ccr
Kd/+ZZ6bhqRrxChFKWXwfOMEvKcErZwcIKy96x61qUclqjFz46553fCzSINi1FPdClle0vaTXbMk
D56bM7jhZtQ5UAOZf1S/eGsTDYVk7tmuGBdu4KYFeVtE4BzFwCYWtUt2tUtz1Mqzg9tusqE8xLK8
RcK99lFBSzsVqjt6kpKE1Jq3LH4QNzuaeARDeYm1N0JobHv6g7MIljo69Kcb4keqsge4DoDeR6Tv
4Ns9NVYEWDt2wb5IlWZDhEJHfvsmFr4ymgpaIXijUnsdwfCxNaCCNB1YGJYPkmmB+BeyDrvz/7QK
TMaZpCtOHb4UDCvrgZOXomK73uKAYA0q3jX+0surWWLMIthdpc+p+DbCQXw1M0WgVVnz0ML7K1Jn
xTxsCbv7JXcNUVYNgbZp+6AEE8sk5jvTK0vQhr+zEFJ7nBpOMkSrzsK3FjBjerJDTPU/lP08lYUw
iQ9BMS+2lLJ9xHxO4bOMe6T41ZybIwbAiXT+/Nv3fPNkn6VbKJLCYsoqOCqdluv1hcaRfi+0n0uJ
E7yTBXTGVfmFEp1pVjlqh+JgSufvdV1uCdyRjsI2Vo39iTtRIPDLlPMXIXhCmbQtTZmMBTpT+Hrq
toPvBiT/7i8ee+AifnpgUlrC6LZWhiEtAmIJuEaF1nlF3ZtgA+W+DkXqMYv9TocpKguoZE5gK0oT
wnbFGS6e2wtW3rSrAm/+apFi7NNmKCk2O2GgbYey/mZNDbiDF6cZvqFdepavFgEIwNHHT0+hL6xB
ZDaNru+OeH65Px9WeI6NqhwJB0k+XHK3Mo5c5TABrPgyjnghPGaBHAlg7MQ0jD8BwapWvPwuE+WI
r9BQKAPMA0IAdmMD5qq/TpXbsfyW+Bv3IAZdMk4+kHhH0Z8WWd1RG0af+nLXiGx4/Bze1yMjC4Ce
/rHwG1hrF/0/510LhChdSDPHXf6W9SqI5rpO70IDS1Y+CfE2QXs8mxHJrsfuGwQY9kPnyEN6wTXF
4ABWST75R4pTj62TQLy4j8XX5eQJeuk1ne9bE9kNOounrGW1qau5PfGVd7bETlhSi+LnjrUj0/3c
3NocbgcVNrKs5bj5RJHWULn6fQyVaRCbVmxvEAr73bdQGUSbfiUQiWO0gcRJDFftQP/MDxZNN3LU
uW3lzO4RE5gR6RPavF4kLRWAuBpf3pqM88AwCMaqvCMYh5Ni8icwCWvli1o776HxnUpwgfVDd3jD
CXrNG+sSUfs9AMgi9MG/PAeXlTqtbHlkW37OAEbzJlJ26el0ZbD+U3ICNImfldBfsj6K0JcL2vIx
h3Ki1JmsVUCG6Qal7Bttshl18A5LeaDckcaKhnuxZXlQXFv0/oPrdPBwiWjpGTAGLquT9txeSVMY
g/iVjxtwWOhQjZZrpG9zOAlOGjQpYcavyF5S07K6gMbQKBYBX5fOXi55zWKQjo7MbnpPuNE+kLc4
f9OwQsKELGNxP8HoqrDGGs1qX2JlriHdkCs3PkPib/zD1QP6a0SnhpghCxaoEB3lbpvz1sD9jDxY
u7ltX1ZTsRbBcLdLc6O8xnP4CSothPodvSF8zlWZebx6lNFv4efr3RJr+mwjOfNVKJpTd2TeZxSS
8cZ3cn6+DICcCqRFF61/kJzbDaYwxUS8JCwj+R3KT8gsO0LwOV4eYt/HjGET9/XBykb3fuwj8cjx
W+art+iiU+HIsea8tm+ZwZSV1x654dsXjZKjBXwpy4DUQo/G4EYsDlAvlCjLrnU+uBGKNDtKICCN
SUs5mnE5xswLJz/joH7s6cSnVWqzvs2euTxDoppWay/l3HmvkqbQzV82MrRA+g6C0m7Oc5uInERZ
bHYcooU5nsKLuolMAjWEKEwfPmybey5v7uw3ClJ+SkkCs13hTYRBSXJ/2VdkbV3926mtZjb2c46A
CLLIBr6CuhJPH4xCGkzm0jTXlSVU3Fxl32u5ujg7Vf1o6SZ3TEksTzjitT+LQTW5hT0EhTuEnDOV
WOgOirMR0dMNP+toualYboyFYsOMPDiLj1N9L7DsxECog7ADyUJBQg5cNwFcNjsrQLmTJuVwPEu7
mH8Q/aULr5NgOFdEV18cqtNqwrMbeiOw2ysVADg7ODBkEd5utLsiNG8AExsQGFPRtGJMssZzsrVS
TD/t1YUViNwSD7QtQs8/SfVpghGA3MV2scpeIAoLKjSz/0YCOkLBIPsPZO2WNJTkZhfcPQSVJUNE
+OYU48bmfaxAvX74Mt3Zw9jD72OZxW6S+xifp82qZgOyaEq0yWDK0nq/XvoHGlMrYsuGtTs4G3GR
6/tUZPSksZUQ4Pu1/6gwmt6IAEGmpFKFJr9j+RJUz/b7hwshgTXFrlum9zGaAYrgj1hEHobTTNTs
dhCHJLpdnA1x4bp4SWstlh4z748XpnosC4g8hkuoRFOPq3u/kPGttrjg/jP+FtwiBYrTBDbz7hhA
g1V1L0B2B7ZM+7mG+EUCdF7C7RDW2KcQZiV3D0ysjWR17Sn12R0QuhdeJx95KcZAiaSMGoJ3rJw2
n8++6oi0sMp4YawewK0D6DJNtvM04c7tXX/fREe762ug3yhWao1BPGQhW0HSF1Ak3H19cKrdd9IZ
bYxPC438xM/8tR7ud9hn9MGWcoGfXM7GkZrKM6vV9DfLL5INcJXI8i+dksFI4PpTKO7cxksot84i
sTVo+vpzFcfglKTu4iOZwyxUFMeUV1c3xvwKFWQU9UOtn2QXFiAUABaZr8Gu4RxYgl7VEvzMS3sQ
l7FYeAA3Rof/1M2mjp23qXiwRhSSCSb6We9P1i+SRj2rqBE0yz2t/y71ebkCVMJRxzE5xO8VUJ6W
46H3qgMiX4JU9KoYcV0zP59SOYedjxBPyTrRIOXWmZjxdqvJSnQdo4fEI7NKiQOepuXtkhno9yME
1e+A3Q3FM2tDEgiVKunHYFp4oc1O5wRQ83quVo9Alwbb7p8UuNqq0iiIIoxyQfxnPAH2XlXoXkZP
10u+xqHiLKg+o2A0U2FBTkZMKzPl7EzltZqoeRbsbwq/B+82tAvlCi0p36vy68Uhy1VrZ3Dwl3wI
/SsR6dlrjf+yvDUv7+q22kQRDn8TNl4UWs/oSdzRHAbE9MOTF5lkeBj4DKsq+Xhzkg9E34ik2oOu
RGozEgkqh6XiecprwiobfQ057YWVVjWj7XussgFNWa7tyxh+dXG7vAcz+jKwcEDJ7cL89FUOJb88
06ZdhodJB4IAAjMIJ4LgCnkknt7uqn/IBMmVjDkURuHhe7GjlA62ZO5xwAyXP2yMiWyEocwMSp+Q
vhC48OE/3BVRIWr4G43BYgpWk32Ld2o1fvNo1X0kDPTz2Cby9B2PatLVh/eJhC9qKmiWXLry3fG7
DmSxLWDwCc0AAV3Y9ANf13gaqso5KGgopexs/BeTqF+HYw2QpLyqvEDSn3GEBsOe6/d4MIcCgJRH
5k7s8i/Okfqcl9SQ7NwUPxEgOZzp56XvkwR2sVz3fcKzvT+XFGdlfDyShrPDVtC4Ybnx8vhLRDJR
Pz6f8nlUPQv/s8iV3aRm2XE5NvBRheuzND3vfOYqWGyRw3eEFu0CCNxohZx777dYa1OcDYL7/HXj
eEOrClkWBqaAqebnT0XiwJLAF7a9E1577Mbx43v8zXC3TIXqWFT8uZAACSA9s7FQVvFhgr6dXaRM
NKLlhkbPFc308FJqHXvmwcHj9lw03daU2XQ3uAuUqpIFromHjX9UOAQ1l1SIw/Wy4CCogCn4G6qn
B5edZGaHO+ccVliCusF0Go5Fl01HItcUPr1myuY2FOhmM6v1TQC+71vcWt866VI+kvZgf2O6nuuZ
gOJ3u7nZyeBtKSpynvbPMWISikLguwhHOeIwrbyoyDH1u7Bvmb8fmC6jLsW88E7T2m7UN5b8WiYl
nO/LGJcUqZRXBMv1ugXQs0lfvAEPAkL8HUzDVi3/Q/+gm+EdsxWPSRazoas6sb24P7CMoOH8DcvI
FQoWw/i6qfWwVBVkA8630zPcG1HV/WSlKJCopu2IL+aeNqeCJwGPVwAZpEKeZQYcsYyRYdS9sJZZ
coRua3otFXEhDDMYi0cC5UsLiSW7ToeXTgdEBoalTxbWQ1EeCaxMD+VxQB4z8O1B8C89Gq1UGOMh
2mM0yCQeLUIa3f0E1sdRqzoBmgrtGxjzKO77PD2GC+YyjyWEzDZ67kHHUmBrtTDndb3jMGC6NHhn
yD2P+N3OuDKyvdAgOJoeoj+3sgYC23D6hfzfccINtNql6D4UIBvVKcAjUwfrhAkRBUYhnvy1Ce93
7vTVRSUjqgD1Q6skdnFAupUKwnt2fllfNaYPFUCNmgDnq4ek0wVoH5yjWL2QUswld//8oa3Gsjvn
ZOZLvIgSLlMx8uXXWJdH7G1pBO3LMp9wghLMtE0REF3IfOgGP14h16OR8hAAA2Mefe3KENwjDYRC
Yd5fouFPCPkjBZmWFYMCX9IO7RYzpYPYrbbud4If0oI2KQliB26OFV+gJ6Qc9Od9fqgyz8BGpitt
CCJIZ1DVMhT2VrqGWZ6uePnhxofcJpMW5QeG+6kcMQqBtywh6O03y4/1AuTeUg+MabHtpwK5gG6J
VlnTB4OYFuyqhcU=
`protect end_protected
