`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
pvYuv8mgK50k7SxbHF7Ddx04sXc0iC5J3CD3dWZOHn9NBfY6mU3ZaMmlg5kIFTjW9PDqTc98AgV6
XGpa/zctefCmQkHH3ilAzos6R78ErhClO0tQt1RM5VWOeqycFiwr1fmDhUmZDcNyB4tfmmiLF+m4
yVVnxEoOXsw7V90pedAOqiOJ3h1pKJzME0jPNsR/FzJS9TZzVNBzOXuKFncWvdGjsvyJwxG2h2WV
ajaiu8T4pxZH2VSfgzAupiArIHQMb2I32oEw6VKi5e/2S+I0NDTGtM3qKr3aejd/SBFoRWpTgfKk
aaHhp1tdKIA8Avs7PX0K4U8QlHXBYcMurSB6bw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="NFplta1hyLNHFo+kXyq/YnSOZmu+UifrUaF+HBQXJAA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12496)
`protect data_block
ZSCq5ve24UcXzKeOwOtV3LceNmqYlo7ypilqXAXM4kRqAcxetVLJGWlQ+7qCPFu2vH/4GZA6PUqb
fr3pFzm8Qzl9C8q7v43Fd6vP17J1/+qA2B2KGWnWAGgu7H2gN3brqLcM3ADyIQ+pfyIdSwc2GOgh
F4ACL9wbWLJtSpfPyRAG9cHe1eJjCARahdIWsC+PilYlxJ6MbwVTdwuJg+rrQIgOUVqUgbolZaQa
SKCsqAib7Gg4L2nyhNkL2oe4Y8sVJTSKz20GWa3LzDeY3qXSCioShjEEjc6IifI2oIeeqiE7Ofhb
g90Efn7FEejrmymu1yXhLMlsMHnkREx6DAddBqbHXg1J/U/MrSOMq05A6X8jALPKui4/kjT63+/O
sf043kKJ0vV23gvtMbxxX75aE+vLgXfp6Ee2KyT7SP5LYDd00DUY+CVjFvp+eiC4aQ/yA2I3/pwb
7l8Xq9ihs3zkgdQuueUghx01P7zxaHsWnMV+BbpXMnoe87vY8caoANJ2DiSGVR909ZhzjV3jqb3I
a/ozhTb3ZsrhGPbVPPxAQeQzA4KQB5iFLkJ90sU9uYZCCLAvV3zvaYMf8BAX0mGVmJAxtrQMaaV9
MmfCEWdPJVFeMAUY1TjOWv/+oJqF3JpPV8Tt61WvT43DxMWR4xWpZY+zh3eiu4pl1NmNog6RuDs9
bpI7tJ/yIMQlYQUHxlTfu5kdT6vYlZZFwYyc1mtnzTxL2uWVaTmtYf9Vqc+scizorldgYS3b3Lny
qNkKJhrQdD9/nhurTp7BvClO7TwMCZG6Q021NxGalEufJkBNq2SoWR9demNEV4s06tjGP2PMkYFI
x6ZzPIQWiZoo8GFB1XpXlFdWiqhHR/B4mZtWN5qSpoHcx+q2ML8aGmnA2Q4iZZic1l2ceomlS4D7
XXytJD4EiIrrzORElyr3BijFOT8zcspKMuCz6DTOTEr+1w8kB1EocdJTOgAcPSRBzBmhQpTELkZS
SMxx6tocbFUyQ+ZstKACP4JvEcp1wIvx1St8+FOEL7EJTcD/bEjNZKEnGOjRsUBIPLkza8ps6Nfc
OtTUOqtKAZojFRV8naHjZUGhxoJOr23zjoapMzEhjzBeUNeMwTGlaDDJEGjaX8hE8iUkaAl7NK7P
TkZd1Dp6mDmdIfWoMgCNqx4WoCWnFuSSZ+lrq0wyiKTc3Odi/7b6eO2zGrzLIAxj/Ge/VLEcZQjF
GPPT6ECz3hxPJ5O0y9+tC8vdQ/7AxY5UGW7dRAKKBRoaVidFGeZUtF0nilw4o7RKki2Y4v/oK7tF
GoG50Th5H6FOhQh5y3bMcsN+kfRsXciWgpq+gvTLzxwRR/DKhGMF4VDEVVo9IOadCYBBi/ISIX1+
3ur3vN0nszRq5nXa6EV+5HjvWSP+Uckj4igZ0PlAnuCzJrZ/RhWppy+Qev1O3Dp4sJBbvTh7kM3g
Qn/SD+FIjoJvHTu7GR9EeTJTzby1UjqlHQ9p/X6RbyQkcMeynVUxQvYhdN8TfXUJF864kipPZ9BF
xgWiBbI9PHTfuWBrt1QKsdoQMEpbmC98ZQk/sVQsekqaS6pBlfGG3VXNlDi5Wv5x5pZKvXXvndhx
n8qvB6ycyC619uNz+Lt9A6iS8QSkGhwnKrFnLn4DHloY45AWX/abl8HnsqcGcW+Y1ew+Jk1p/7yY
aKIyCI9ObGbaAjfdoz5jAlCdpp4FbiOTpmTHfSmVLTTTjis+V06TI3geg8mJLTHnRLvqcqrdbsfj
oYewj6CyosRW2EuBLw4XyiTgANIpR/bMpsS1i90oTb8tMuhtLzhvc7knRfCWC8nV+a4ujfnARfee
A/JBOtRAb27vaAedcSHPjM4jqwCbzzh7ra9P8D7rWT8DML7D3xrPcPAwD6umhE0SQ7GTVYBuTaNm
WZElmZcIc9xvaeXY0FQo/Po8Ib/lFl2afEVMMn6oWUPee3+MVNcNJtkOvEhJ1LF3b0bOGgDgXXIY
IedeZKcHYDmYenJP0qwpXtvNrNVJuMsv7g6zCtkA4iHMrZXfJ81/Emqk1Ifqy8kNYne1Zr2IFkW1
JT3VYVMd0inZOvoiCExQIbeeZhZTLanrF2U9NjH4C7XH39pEmubR+jTpAvobwBah2UOaFTGKPvk3
xSwOZGUlxjgB1j5ipj1I9X3kYxyxNmBEpb9vjVmXHAazQSC+rrFwEGT4iEkTEvwbjnDV3LiGGuJZ
ENYY6udWpOqdwv35WaGDTO480WVBYa702AjA0dgrLhaDaYmCsiZDZ+mis5yuaOa0REGvzAh5jOCy
tvtxZFQELLhUroyzzQJOqbXfcQ39JYB3FYX58HVlXUYdrhGKOfYNbUgqVBxB8Y+vsLv7sKaRKouR
zMaye/rWQCiD3v25/jXfJ7eeiD97Ad9EiIP2TbQ6uch/vJ3ImcKVzvxdbLLQ3FQI3VhjceNA7o3P
mXg7DR6Fvc9yfz3/ADtGvJuH0F1hV2D1HKCcUKZgajUmMTzWGXv9LWx/S3vdO4+3YOueaGLYRG/9
Zv/Y/UqQkxsFlyUKeuHd5zwz1vm+MwAA6lQtzuXHEFb6IhPDXzdP4jPx0EZdleelPTP5XM9wwCIi
AkpBMOHYfe9iIRp6z80MnQAJ56FkemU4FA1t1cEA8wr6XTGeMtGu4r5exct98QLzlP698M+3fTyT
uN5Mp6v6TcAaNDLCpETPNyzfnkCffJAuEc6WXo/CEb05k06EcYysHN0ZZJ678+6RdVYVqlVjBmxO
kKXqd7KhNdoWXRWQqzwjfMWTOjFzUmiyUKRPaq3br0C1KCypXx1TUd+aR20IzFxLoNz03wd848yz
3I8A1NnyR9z6ZxsPUg0Fi1YztO59Jt4aJNRMQLHCTveb9zEQy8tML9wXTBtLtJRMcXx9dIu//9Fm
BhtXM1u2pGBqA4cHmOZQmoY7HGtcdYzezjn6yH02YUmMzR5r4g+Z5TnY/FwLbR9WX58HLzeRU5ff
/yEWQg8R2zIPDC5JuTW3G8hUJ7Yz/wHbToe0TI7rT2zvwaEaACox0zGo743zjXTT/ZvNmy4mxDCp
RxcKm8HIZWyQLaIj87YnTLaSd4eoA4EAWmdfpwLcTCMiPttlnEdZL57EWnGb2yFSlDBjW+JA7ozk
9oOK/thnUsJ6/IMjigBXhvVlvUKFqG6RvxZtRTfR3K3tygENd5p/K4W2KJOgbrvxCUkIZj1HWpy6
xH3Ht8P7IunFacOOk0OnkO36zkudUkEFlfDsydTyFwETZOOSbQ2MCGUt1BmooFK+tOkSo1fSHBgU
Fp4siUkURXx/YW9l0nNc2eT8g1+AVZ5wMXw3ZmDUpIbHZ2rghUzd/smhvMPSpt1HbSnB4qFWH2c6
EMrAHq5ges7mafrwGM/+iO4GfYFYXn7uSS1lJhn3Qz0hHxQ5S3gTh/VXmjragNWznCjp8QYXnrSq
Eb9gs3olj4Sj6Znki5ygdaocRp6NyvMBH+30NluQfGQAUOn8vqkQhwWKRunxZYQCazO2IEgJGbs7
PlTjR2SOMJUb3kj0xnFvBWylfk2R77xXoDS6RiNNfztGk5AXPdmZdZD1rS5fx6/uuwiwhcQ07/3r
yYxzgL8UymDQeKKmDjNLXPJWBj3Uf4it33vTzFFjBlg4A7pMe5uQ1opPTMPdL4P82G0G1o6m5+VV
XLzu+YsiiGll497mvqZCbbzW7sdBv/KKIE/uqpBUSKsAMbHEuDfxKsUAD/MPIbpaAdh4aPGn6kG9
U80e+/FAyMwGHKnJZ8CceWvebT8ARYeEeMp2WwL3BwGqPiISrrXqR3TEvkx39WidkFWPvo6v3pr+
lzpEnwXVBbc33PPbHdHb8NHzW0Izyx6fUnHeVMP9xr2/tdQtrWSar9ETAa3KU75CSAL1oxlyIxG/
RyZAocbjCNs7pmLiNMqVGuNdn3HwKF/8YmbF7pKNTJEcn/wRPiBz6N8gxZheKPz3BIJfAL0zInh5
a0OdH4yjV0QKGTYoH3seBILOeaKhA1z+mtL/FjlyOsBwMlIxbSVYzrXkGAHg4Qkb6r4qS9h48jdf
u44kfdkqbPuOEKTKKOfoC6/WsQpVyOBCIM7ZpL9itvkbCwmNq177byfllyeQ5GA1Q2xX+3M8yNEI
qIVYB4p4dYcBfw4D2PI17iwUEO9LnPyTLOZSqP6SeSi/T5bTBxH0gO+XAw0/9Oo+Sad37bkMVlWp
FwcTdcOMqflwzxw83lITCG9XT0eXi22XR5K8EM5hsmuI0kp8xPdMCYjjB/ECUDMLevV1yVcIjblC
svu4GgvmtvZuPiGr/8DOsBrPl6pM+F+fy4xQ8v3oRl384T1MTICsKzLAzrIAAP59S/JdLIFhFwyT
9bKtKSxTQaiqHzDYVebA9eFj9cY1msw5wdXNmZSA6Eb7Wqoi77A8ZIFoRopubsUU62YRz6dBto4w
6qOscFTacGo7Fvzx3y4o+3VGMsN43abF++TsIJNEQMEe9dXfm3aIqAweBkxgolS8w/tS9Mee+thG
fOVr4jZQQJyD9G2o3Jp4BQH2nE/hoPjM7/ZrP0T3cWnVRQWs1hZzHGQ7waAQn8iR+GPSCFcdM24u
pUm+g31eyTejr+HsUgFfL8cljA3OQvawtXssuuZO1CBi56GCYAVlXTdSVn+o/da0xxOvlZ0XD3zt
OZFSM2fSgwydaMC/ZT4FOIoQoa/21QlwpFRNDggDghrqtaq4+N5zouSQ2OaTfU70Zy4B1nusxqlw
yvDS0Hg+OJQobXkySPU2HHnn8ylP8vhF7n9MRnZWUXNOWiPmJAun4GKL3voYbg8f2QxZI0LKfPkF
ff5h36vQ9iAzSheyxYXlc6DkdBUpKIaXAYPu81q5UyXXrg/ny1rAFaps2l9dMzLSJSy3s4DLptS8
ay7OAOCBciijPfanOHGTFokB/6jmtGG9+bRP/Uvhb83Us9p4qpM4ICu3LnD2ZMGWOjM2FDQfnOep
ZJ572CodvxGcHTE2vu7l11XYjRwW0AaQTrh/Ucozsec1y09g8YzNDp4qzqfFdNyLrBOJp5OPk4xH
aYhr0UiWAafL18/kwNLgCOHubU8XQ9dHsnzk4H4y0Yrk6BVD6R+TAjnTSdfe3Zi/g9DhTL65Ce3I
arGR7c73Lej1dZKnTMW3Hohrm9CmKbLDZHk4PYFvWsyu5xMSXZnpfmt0wUTgogwt8Zt34reYfsEn
HZxV4vyTDORH9cl8AjWaPadMVlSU1Tm9DiC+TuJLzv+8JlkDhg2j5ASJOLvcOMDaKGZ9qsW8tebv
knHzCT1BOinboF+SLvC1v8mIwlT+I+18JL8XmRal5Gima8EEkOKtC7389jgJYZpcgxhh4PIS9npp
G4cfb7D+0S3oB92PP6j+h4OjnaCExnr+iBdVnMFXmnCyqtQYpslxCJHrvnHEza0DPMDKeSo8GdKQ
UAYzoo1fBZIsm9dnrFgq00Dx4iQIBornrvPVroO/162X9/6kntGWgdZtGF43wD8+hVazcC7ME9Me
cyPMOA9fjzD1zROnwcvxDAISLNDLSCjBhiV82rt5U0ClnBV0YQ0o7X49MT6mACsSjcveGtph5tJz
Hw/0o4lmLas1vrE61vbzmdm1EHc3cttSAOj15n9Nf8boBKnugtyee2309qxcmeqRJoj39bDwz+Zo
3dEy81GRaAEPqOIz65mevDgNUZDASKqATwHChDS1KRLmnGluNtEXeqKBipbf3JqrTqdvhlSB1kT/
njS1+EH1T0IjiEwYZ8YxC/CWrEGRGQ0vgv2jjFqFGKEL7iihKm/6l3D2yrn8+Y30sWmVQ7pHVD2w
03VYtPMoulPBJDWbJKpDw8My+gPY/jNYVFyg+ppQ+PsVH/ghWR31d7V/rQ/v7J0hH8Ut6dxVUhAK
N2uFAw702n+bHWy4L4Vw2AOPobkdxnfksmiIY/QonkZzw2A7NsBXLpWHdpiSm60wtdiuXYyS7+8V
zzIgvYjfx0LePXaGe6zl9twUMZqY2G+G+agTIish6NUCRNWZMQ22t8GhK1kRUvNB5NiEPeW12aKE
1ma62fyjUEn/AdcOLhTRByLYdEYwZNpCD9624qgwj6J21wc/QJmbctALArmMun7YDF7JTEHgD0/R
IPDKVGXvFQWcC9DDPHCRvHIX5mUW3AhXvSxExsYrzaNiY9+NfNGsVNtu2AaRyw1/HzQ8+3oxRVLl
ecjf+pP94td4XeROB947G/cYUjNW43OUIvxAmH5QNP4H6/cvMjc/YroCHanZH+Ig1aPaPdoXiMy9
zd3fnnQpxJtRuCZuqXTOKuL8cbQhPOWxuVte0SdpRR7MmlcvaywiEc3PzOFHOwAdstWpYaH2a57a
XzmIRb5eQvD417aOPsI+9tYLIbRKtMl46NEtg/xyEidsOh/mGpSYuwXend694iPiuekevU1NEIOS
tJdgbkebf3/jbxWeJNu/WNzvyL9ZmeNWa0Ed/nPmOcGAtD8LlVOo4dLaMzle/d07f2bfCCfkPJ3Z
QvqWu2Na+nMMiIMECpniaJStApPpzNRyTYtlrtTT++knlpv3M0Eda8U1okci6ZO1ZNnUHU5k9A7U
OZL/Cq+Kye7MQWfVRWO5k7RoRAiWoZEh8fpyyuatdCvD0iyF7L5gmiG9CzvnnAQg0oMuAYLz6ctc
RfS5ce6NwvC52sz6Pj203r4sDsgdHC7Hwc+7B+pxkChKND/PbQWB57EDYl9TBXdviVoZcBqW6vlj
OsAN0WlfZXSUfm7ouq5yQxxu/SghkGchQNXImCDofGxIwIxuLrMRnyhZMn2uyKc2DhRfQJuHfXq1
u3wk8ZcwPQlkv0LKn1ga/SDZZkcFHlTAzSI/HSbbEdJU/4+j8MahTkgmWE72tliMiIl5dBJ8qeUh
bZXTXn0OjKXBEh6iMQ9upAV4R3ZaBEVEylxhI8qOsXW1Vntn4GVVWxXbO6quOwur0otaY21+xJyX
i6S1eHrcqcZUBaI6DNfngIFwAC4I1YIjiz5c+Eqf2c2S129QiFwE0xn2fM17NVDDJ+8j8cfIBVtZ
m4xHSwZJDmlkDLzUSRXWlliZ6fd+y9uIPBtBhvi+hoh/r5ZELZXF7R9Nz3VpJ9HDZ7guxzYLDJH+
IqJ6GdZiF8IgPQtxmi9HwMOcfOLwgxlq9cWqGgJrVaeZOlA67MrigclKuUDXUcowH8686Nc/mCLO
cDy+CgOV248DSDRQbx3dafTf+boTDJ/tZO9oqQP0PHd/kVSifqitLuZ6Uc7CZihPKDnXFkVzPEpV
WjfjwvVYPdwjDpQ3P9MTcte2Ftl8UlE+QKgUBEo/hLDi0J1olBlxGRu84K1viQZtbjuT/5sQiyg5
Qh9wvKcxyiY7J9MsoAcPGp+W2v86aZ1lJidJZEt85ZZpXJFLGXpqa6jCA+qwHRMqPyi+ZWbYCNia
928lK/ssYn7UKcnUerBkde8z25PX2PMBEXZD7xhYiUDhLcGCmPKYm2pqk0yrzlwSolFrx6RRR23i
j6VN+uxsgTcVDtygONp7GJrA0l9lxmmtPexrqjpIcv/UkoBqh16hTto5+iym8YEvZsUsV+uWkEIm
o9brXLsmLpNrGd6I7JfeMj5FB/aDj7UGUKcBcZlOFPpkFSmq5Uq+TpLmc1vArDHTpXnrM2kVtDH1
smhvr489caLsvjV72l8htOSudOUOopAYS7yEdAmWuwp006kbI4SWQyFfsiHxUG3Us5qgQdGLQp2R
qXFf43Ig89emd/WG7U2O+JgUZVVtmtAi6DmDZ18bhz9NIwc/nHUAGlHsIbDEGkdig1f9eu8nD5D5
Z+Lho0P96V19y6ggvZNoUqeWm93nfHZNEBnsD9ZnWQck3DG/bZT5rvUCQDRELwnO/Luk+lXKLJcI
7GtU35C0CUiDRpTRmp2vAUbwHpH+eSVOAH8iwLdNDwEcS3OZaInkpeF7NipLOgZE9SJV4IYWYgs9
f0t/0ARDCH3aGQVvjVX9BHuJR1LDAEVBPhUOpSHTInWy86ritWwShnjFiLSPEfLKIptueEA5i4sE
RVJKYheKicezpGx2acoCKwIGwfUV2CfAZ62HgNx6b1dgzGTRFQUTRSxSCi5E/z6m/BqjZ9Jn05VF
AqYod9QJMk8d0ivTViWMzuI6corccha6wH1MawkKDvjEoiHSI/hTui47xsmP/RKqKTPEO4Lad8Am
pxL0fZanVtDGMqmJaAN4nBhAdA0j7NNMhOvg4/4xrLGbHfcdU6+6Jzi3UtPxVMtjUG8rr9EySyDT
RDkyXHePSd4RLWrVgHlKw5VUurx1fCruqC5frqdq7Yw+urw796gSkHTrIBSD1JAGs9PJ9Gs6Pw1d
QHStu+S6d+WmZcvvO7jLC/LFcjlsaBLWEfRItaJkPV1yqpS4cgnT89/JYEno9UyZKxlyzC6HSOOl
8W8mQOLO9oYLQSr6Qd1zrM8EnWcXP4O7xOwWtEFYs7paNNwFKJ1Jx9XBiNn1q9oQwtyFyL+j7ruW
7hdCksgJTUxk3sZ3nPSLl1Y88RA0iltWAfJWqXDjFheQpTcNM3hJJ7o+tCLdY3uQ8/DY2I6a5nyP
CKTyS8AiATP8Q3xVHUqVpauRYI4z0pbAovVt8zH9aEr6ecYGtjOOHIFbn0mtD9fp8x93Gg/1+lXZ
3+qcCCHettbPtyQdiwGmdP5klKtYaAJtbjIOXiphLJLF8lHdedli7vNYBj0/ckCGIDlmNrr6Zcz2
L/ywxK/t23Dn3Rp7UjfCMawfkApDTj5q3N3Yb5GR2HjwfnQ7T/eVRbF0ORdmg8hVZEQzO9VC3bOd
o/4XIF8Xovg1clz/0G8L33OguOeUcY4Z3LYOAv2zpHTyzJ3k0ZhsTJ3iqzW7TtMS4NtGIOObkc3E
QDs5V/DjNF7x+acBTY0XnDE95tMFrNCUnrHVtBhH98x0JClp8BbdWX2DLqrDv9CCLXJpoyhDEVZa
QWOeiQ3UaN2hxyNfs4VvWo11M8IUSeH+64FFXSn99mkfuK3OMwGmySpKKEvIdvHRISJk4b8Ip8Ix
4e5Us7skviWepLD8UgzlDpORUsujSi8x4Nh60XJYoWo19byKxTP/TEfImQyV+HoMHETgVZg4LY70
xFEOEaFNeUCmgYAdBPfChe2vKcB+OD10SuMmzFSDb6LWWlYq8Q0pfRy7WksdBFyKbOtwNropiBSz
0+y4ZT5UCrneAwaaKjlqEhnWEZyNGC+gd6UdtfL1BnjLCx9I7Mi4kpbah7+u8g8yjkqzNYT2CzCx
GIANS/Ey4GoXtbakWYcZIO55Au1WNXbAMTSuVsyC7yMWiORezCZuIoh8MWVYApraoQyzhJ8kiBqv
bHEBmvpxHDQqHftkHXvYFvPe2AvFGNs8Qb9xDGoKfuNsq5E2AFKp6rBip30xMYbwmWlZAsH/PMVj
CRrj3lFPqEzU68jex5li18ij+X4je+/Xo+sAWJeXhJ+m5trEb2WnFyo5WttRuIR5qXsk1ya1LGS/
+P4sloE8XkXiPltxyb2ZPjcqqVGkwFftaK6FRYSFd/pA2B0IM4qpRg5hA+0np+jG+AZESGQyeNoS
nzR6knPtR0breaGrUyDujaNugC6MAVpASpUB1DL/F4O75/nZTPCHDPX2+7xFDSzzH3QQGfyhLevo
TrO6DOvBVPvHONwBDceKwVIUyiGG3hiFQFa6q3Rnks8qE/9vULJaBPzYKVKYU5TWTI9wW5tmGv8/
9hXAX1B5VQuJ6bFxCfel6ib6wfKoZMsbnr/eRBVeSwRbT946MVq7bEvzlU5Lv8BsjoeW46g6IA6a
8sBosS1aKpJc/g4McVHFKgA5xOgcdQfA3Kul7TkH3483aaU2EftOtOUViWtBFUnY5adoRPdPJ7kZ
2m1aS4KgVSNpxFpBhtIdnvKl6MOolYcGqbQIixJOikHAlPP3pK9NRv0kC0c+a7srpbPh4XBoiwDA
q40qDcFtpeXtBcHlidChuCthzElqHq0DrGmPT2C57cZXkRqgrCa3wwcR6VkC/uDu6HDjHcJjRzN+
DTIqHH/2xs9j/ac0Zg038rIjPv8ZcyjqSIb8e2RmLcAGU25hrBI4QCd5xVU0aQR5z7IfcHmQKmhe
iOaAcO294EgDbgAi81Bp6VY8aH/pwhJnkXdoOs+KVGHAtSsOUYMuChJ5hCskjurwkkkD7YjwEszK
01jwhSQdHDErCaOoliEJAI5F2qzzXsrYKauDyoDfCbZbL/NTP63z2K3kokjC8LYRQ4DWWc4Au2mu
2e2yWCTtqx1HQSCxEe+ARJMTPdxfBRP6i/7X6aKNtVN/6t61fJhBgEbKdNWUnK8kQAbfJXXNazXx
R2vbD/e08QybQPmi9Oioo9KQjQbvZlxV91kb9wo0yKXMGVWWVZVy5szViT70/JUS7Br96ygPnWjj
VkeraQbJme2gnJUPKS5QdA4b57AT6A9Syx7qbld7Wa6VFAlC8pk8b1qAAAFXGnhLB3tcknrRnZXh
kNJWfo9XsLskS+2pAtFp1wqFVrPAGTiVFV5kdokcrbsvyyl6BalCdVju7sQyF6juDuV7BYBfFyH1
8xgfcNObNEgtLJBX4I+CyLcVyYCOC8nMDrPHnMgfCH3eUCZ63fNLRP8j1Gnrqz9CmYbVOBMpT91I
wucYjTdcK9Gn/5YV3NmZR9OnraxpmXxVKegaApR6h4iaNlCDH6cXdwPcEDkKzSjyw10IvVY4GhMN
brS65x5RiTEs51zucJ5CUT+HHT4qTsC4WYL3pCdOCa7So4PACUkFKxy8CrEyf9Fm7nASbUSrOD/e
skoO9QMGsDEDHmC0/ksBAU/KldXz2Xjh+czKWqGvvAbBk8x7uK7bMGaVxA9eQ/yBZ9PoAfIN8zwj
/dfhRkJK1qVbqvgoyeh8RbMuRcWKIhL8Irr61TI0tMbCcxLvdOvzMjA6t2qznZYDizKM0jdOuEVH
U9K4vT7q5VoWzyf03xya1kvWJT3uCgonFKZtCQYViMT6ZuBki1NtBTpVQBtfK0yX+2oJsXYUBeXz
TbLF4FjiCfGC4MubyV8d8dCJT8/Qudcye7jFwZQbe2rv+0qQWN7TR//lTXSjzKkUG3z89Zodfkz7
LmugWzU7SI4JO+ULXpNuPDabvqQX4BaACP9tUSuyrJ1A3iRZVLizzGxErZDTLx0jrF72NRqabrwl
2ZkIxLabLVSnkypzE1Sc6VbSHCmrMjqge7MAi3FXAZnEL9JDmz49VEpQWhE37RrPbs6R2zPlCB2Q
v5NIc9JtyAZJN1IxStrKU719UHoqyrKzPdfmQHcudr8MFaCYzHbbd7t5JbeuhqnkVgsyRTEFK4+6
g4R9K7UkI9+MQqTOncPsBT3l6KBORrn+4hratZ9tLldneZpFm2rwFkXsFA282DFAUzATtvU6ArYo
lGstSfgkyUT1BxNUmKBqAV9J2CJUCl/frLpo/w3c0FQWjEftdyuRsFNeZwbH9J8sVuyiFSYh1rFA
yn4XPaQxagmB+yhKQQN4VEFytYK0SiZv8q/ZOBHRMiMAUAAwsHCvCJyEh7uVCs0UAkp2BhXAkIzC
c43jFEGZ+Ryd8VozqEbNfe2CHosYU/xdpDlLpAHAFZhDummE2GS1qqiIVtxJjxIL9u9FEglcS+zG
XtZZXBYxDj7Z2iDnwcpdxgQF7B4z6Qlp3srT2E/Vx+WgTRkbEMfT9T1q/R7/sSiDSM5UdS9QUlwj
h3QMMUsaZWzty31J7WRDsm1sRrlRxgeIqeMWxlW/WZ9G3asjBW4eqydbz4MvlLNmZU9KmmZSqScm
vVQGURfyb5s6XZyDTRd02EdrVYifm+i5H8AMG8RoCKDWPNvxLdFWyv2rJ2bBW6mxbazaI5fB24x2
x2LMxLa1TqKvN19XlwhHSelYJkyYk2vg/rlGxM3rAgpqNF2OsxjcbW5ZFNH0wrxj6prrSDvXeElP
i3o++WDJtHqv6oS/EWavIP/X92bpji6/ZHX0wUHLN4h6k+C0XEUOIp1jO/d3tX7JgPc0jyeQ0lHg
mGy+IHjhK7KcWw5Cl9a7eOh6yv/CZ5js7i/Ct6xddoSQZemDBfmunzVwvaQ0h5tlzSGfjzScbesx
wQl6SyjWPz0hQhJOTj44M4f34XFSy2SI59mZX5kC2Ya4aac+3n3dctmUzYReickc+stu/YI3QHq4
jTRi7DduVmMiaQLEgOyNXHgVPJE3wfvpRI6toIRUMKoyP1H9ugje6g8BuC0QafdvfKgNqKLrZtMw
IBOyrT2fdeEGoMk0vCU5V8O1rvLvIHE9j3TM4G9g67e2QbsZBpeFjW9Y6a/zo1s92XgZUDD/cxe1
WU0LFrT6OkCGzTTIHb9wJKw/F4i4T9SDMFA9LIz2eoTNJgxX1ImMf4N7cluHgWphT5z7WQVmyhUh
vjbxoKpFn04+qAw3ffP4NggZM4AOsSQNaIMteNYryfZblH0CMG6/zJ+g3ovDPshD4vT4AHRIW2Nx
77guM29+ntlIEKuT1Cr82HTqf1Axg6GbjTsaMmuoODZIZB1yxRVHlAs/G/ks2eVVsffOa6p/yXEi
k/IjrOVTQrymU4MXbQaSCkHyLggs5wryZ7/xm9QOARINI7aO6EjMaesm3EzM9oMV7K54Dn5HHeJu
WCrSNJxSkM4e8xwFoSrsfUtViC8BaBc9QU88lUIG31QuE6x9iOuwA+Eshe5T3ne/HqyZbinfWmns
UKSC8v9s8j4sVV574+XgpHYqaEqeVcVkEdpPPDKPZiM51d9768C+y6nuMAjSqGjZCmzKvkK03qmy
SpZIIKdBfLP4tK2m+dXHDtHcSQAqz4ypSAhi74Bl400eOAgTWoz7WIAQDxOdTYC33Pu7viWRfmWk
CObaJjC6KsLn1eTmJKhoGUvNtxVs6Lbdn0P8+gi60SVtC1z1E8562glxj0O2PudRmYi1m1yNlmbd
MtxaG/yVSFVNQZ9z2U4JmdpRw8Te70ItiFcgc7k5eBM1/1HXkg9fjJgVl3YPJ+PnxGzaLRFf5zEB
a8JDDCrhAWtaJcADz9cwjjOLhfyisXph91ubpQatY+QpM+XcsevQAN16lGj0AozfeRCKA1dwHQ0h
DI/u61J0RmDIr9hhVK/0rz5yqZdbkNlLnUByV6z0F7h+0AVl0T6e1JJyMI/IlUmnnkkxrrnC8wql
SqCb3dOrHLOw1zaQz1D0X2c30y3caqPvzYXp8fToORIdLCNB7pfjdYyymRcDdXwJlBiQUtUnxH9Y
jl0GyY+o54tYw88s+VF6qZBibYQI2RX21cpsB5sEZ20GFCNf2/5oMjXRLSC4ogR/UCJPb6sda/X9
9c5McBK2XGBzYFWjil44k1bORcsz+rxiz57awSfaD0Be25lK56mufsLlU203+Tqe/Vof213QYaIk
8dlz1r5WDXvEmltvD04+N/1FFEA7bq7ZNHmN2YHuu11f32P3IvBKwYz6m5TlKngjewyc7ZY1hQVN
8VDPOenL6fAKYLDm25/lDRDsWrmtCcAOUvk3XB4kHGSZVChND3oydE2USyJQhrjUCb1iFv5/1JLW
F9FQjs6hi4IgrM7XCd8Jq+PxrZ5ltv82H2McYd5eltDsGF9L/qCVNsJARl4zUdtJWfHVHyegp0m6
FEIYCT58fi+T317VfA32n89OO0w/RzN64APAIqnlTUiByNs2eQvLylzOJRNcGNXQtCIdX7BlqDnB
IM32cgtD0klvQPy6aGk8BlveN/wq9MaJcSmfKuTooCESjVWfi0vUvg+rKVwQQvO0Ohx8a6EYJFEU
8ZK5JWw0QPo4/2NoLXBgM0N/S+96KQV21QEDqLaXx2k/w4ZCsjZFxyISwU9s6toJkC6RxO7o0kyh
zlZq5WUuT8qMgRlWrDdMCNbm9XREHD92Us9ldBhidYKHElOWW1j+LplqaQB8OAojYOjjDbNHfXU7
JwzMU7FFYSN2+/IosEzOrq+J65R6CMcUrGYwbMJHeyHURYrY4bIzh9oL5L2srfk+APfSmtX5LSIf
U/+IZOPxLj2DEYyZJsZlbX9cgnEgJur7TutKv/QE6pWS0890VVYTfGFm0Ys86GGitiMHchrsh8RW
1tt+e0vU+jXtXUQu6cX0BFKMEFDaDTzjrxQH/Teh0T85gLHNd2hn5nsI1sN1uQRIhh31tCjfS6EA
f5ilama/jQxi0BMGb56oeCno92/ASdW/WKQSwIhGcLOgW2jzf5oc3BavhrOYZ2teKxW5DEJEf/pP
M7u+mGLqLE9XeembL2EZSvQjHLVuBF7V8bFfSsl/08iRtGOXuBm3Nzay2hpacpoa+6gzZuY5rPWq
JrSU+QfiDZYQQP9z3gir6ZPxun1KhyznhbkgKgL7oz/CqIeRluDQRUhGOVANEF8t6QhHlaBGQRFV
XIPYrX6NTa+BZkBdh2UBNnjY44iDFuWwlxI68pwI93y5V6GU3LxWp3IbQKRv8FvvKAn6tFljSFMR
r6K/ZljM3wHJxHOn158BJUm8+zza0KRnHOOl9uzU88fl3cNDTRAcbUhV4cEVl4wA7Tuwr6J7sqvZ
fJzx0Wmrr4CgZ3rF7xoZybEUAZgCacVl/Pjak85LW2WL6GD1msylGY2HMpvfOOV5Fr7WrWn3GIoG
4JngviNmHwKCOTe7XKwz2e+vtqTM55dUoeStMwDDGNI5tsx61dWzSPUiTm1apdgjxJHkGICXDTTs
pSIHQJ7a/eDZBcy2L1C8HcHir8JRqetAQ+7es780nBs1E3bNRYXX/Qr+U7/L3AaSiX6idaGJKa04
6doUPm9ULEfAi5piROvFqbb8mwUcP1fCjXz2XvwPYukAqBeIxLaMB9dXGumLzv+zc4/FhtBnGmN9
h3YLLwFP6VY/dcClEdGWBm0VFR1YS0MFdxr6flSyj6WVfosM2WzrgRDw+qZ9b7pwy0nx/iT1xLRm
0ZWRYDf9aZvfUfgrQs/nQZmpXlx158Qx+pSvLWlKZ288gWTCTsWx59iVZun4dke5sLCnZejhSQqE
heHACTQHmLF8f6OP7C5h3pB0+gCcYPPH+t1AoOu1jKZIfTe4g8Z043cLVsgeQpASSm8eqNKsjUPE
K34HHysskM6W9XdYuZMnimaDzMUYk7Ny5ZBHolOR11PZKoJwnbQCAlY5Mqglkgm3SqfoFa3NZH8w
MjVnl79+Q1pIm5Nlw3vGwKnp1AP2cRke7oH3chxhNHEo71ZzPOWjaFZSg1uXvX3dpaWWFL5aJGJ3
vQmd8VKu3eG0/Oc1rIviRAoaJfG33BZB+A4cmtSIrpGoLmlxf2pgbHEDEza30xoFLTMaGpfh4+nn
z8IKi4JjM63S52yIUajgWGI3szftjwSPRgmFuB95ZtKByyqSPb4eVAzcPAJFoBT59ygnGyuhgu35
JhGytSrWkJs+8Gooh4A6j0jKcgO2SLTp/AjapvFJ0p7UGO/JzxqlSfqxCeW3fuw48uHa/FhJj7zp
l88iRkQexn6zfhaYtv78em2nKPhXfk0OXvfpmpLlZcQ/nHn1un+988NxOiC86u73w6WPXGqAlakn
8YST6L4VywocC5f0oty8byB+VC6X8ebbGgyRYWBeAB/iI7Z+Kvg9bUd8nDkVHJuJPuw48YQm7RCZ
ONf5ZCb+UNB9Ccq0g1Jemx1zyDD0Uk0KKyNgR0EMCQ9Z7mX4Z3yfsZzBa+QmI6dCoIC9grmDTegS
8u1z8Q1n4fQ45NHTmkXI9JyXUIF4ujkmGTPLygd0IsiTKDxm0bMho1cVAQEGIx/1mPpLKl7YhRHv
/8pDuv9wmMlvmkwb2yQmxjDWruD7rdE7JjuIUzSjVGJflK4krvXjYaa3Plv+ibFIKQCIF/95uJix
4NPAW/KtUENTrlHfOJ5IVeIzoqayzElYsJvUoatowP3i07Xz6tf1PYK6xLNw0TnLQynpKVzPFwD7
8lVStoDtCK503lr/3PqhPiIw6qLX0lCCwQ6Ji45cxRq1ObhjFuIdy54M2oE8+6TEx3+nuBucEzZm
ZRE08g5+nO2Ee7TpNANmhP3y6FCV0mszbyko/cE8SkA6TGChACJd2B3fmBbdRNuT7v7qA424Nd9/
TZ6kxWZxLQZ1ZK1v5E3sEhh7h4GwKvNLnwJ9Td4lB+iNPqsE9pr1Jge9OSDb/qZKstOY0FDtio+U
h7ITy4jeb9oz3G0i0akuYfEz+mrQzISy+qgHiV8dx1dHYVUh5DVIgTyZs9o26fLTRaA62zb2U8Fw
11BvYMYrzHT4qfLJuCrpnAc7T+Ldt+U8Vpa0KhYtPLLefQSyihBi9y5RyLzZDWKo9xVGhHyj8HyF
kuMNO1TD0RElh2L6n+Y4DORzpISf5jC17NaEj9q+1hb+Tuc0w9cDTEtPwelHCYBtkII4sYtkjNo4
LZSAtv6ECoZYzYz/gD19u++SqNfc+LDER3ZUvXAF1KrHhveCBVvOcZAdrLYCUOPyFK9mlbTgy/Xg
cTTYFg/aesLbJWnJuTUUE6uHujCqzGZF4NjmpcXyGbmcHTUBUbChHn1Me2ySV7IUEUYWZ5FKRcLU
Bo1XXpM6bnfjFR540GTXWI54Z3SYdAXoBmR/tXb0vHho3FRDjapwig/rEmtIqrU1H7finTHmdpwG
KIiFFtNuRHQNscA7rT9vYbIq7IFN6h6HWD08oKhWHtBC0AdPvgaDG7F7xE0BCubZVTFO/+cg3T/G
iraPV8h6X2mQYGtgCYHxxEhsfAce3VrOTAYTZ6jRwsUbNl3xYwv6UiGorC/JeuPuNEscGL9LhwaL
7IKLsR0RWDXxQJxaMQ==
`protect end_protected
