`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
LtPJJSIERtkec//EB9Jz/CyRjrEIiiiYc8rPY6P/87Py55qBc8GVqvd5+SCohrH1JNeIh+KrE/Ir
mTWSiiJOWjFu91jzgTicHoAVw/yaDTZ5i7BtF+Abmlz5cvpTGWc0amMuuYkNwtZvGGPgGmljQiV7
IVWlzlqq58NdpbWgFWrfpyfVAMUfYcvGxTIT4g6G4MNVyCJeI73ZhRRNVkWNEqR9MZ+ChbTYuCzW
0NGpD7NPv3b106yQDXoEwWKAcJXnCHJKo3OAFRLtiJ8wV8N4AtXN1mswFxMTO9Gq0ePWowYmFhYx
+stOXevu6nvyXONIjPRlDIaEniO6IyE8iRhA9Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Qg0AJTBf9DMd6Q8h9wDvndhGF1vFB4O0a/xWdgblSEo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 171568)
`protect data_block
D+i79zdGJ5819Ulzd2uU4IqZcR6jvLFUft6XaS6RRas9DWi840slsOdltt+FuLCwORkaNpszHIwf
KUSHCOsQcWoQX4Q4/rr3Al2KgLVZ9HqWxkAOsxCGshtX3tpDi+sOWurwsRb8iU2sIM6aJhkvz/uz
s4A41ig/PaM3Cv7JDUMdrVotK+U+Ro/PjNuBpli7UdwKsCtGW/myXPkKvVRYN+3WLUm3jTiriqHG
zQHDu1TkJ8P89aU2nF+2KLPUhcwQK+rYq476BPk0sU8jdC6Qh2UKWr1X4XK+Kq3UCutVvTgD7eUB
knBQeDd/DRAqW3xpkNsOJ80cotwdfRXcPXMeMIaSqPJqEjdIHIotBTfxzLLtrOjKj+rwIZpFhm/y
DW6NC4HWD6vbWpb0ok5CtrZSRo+i/vcQGDC7XRvnFWMR5JFxcW/O1i4+cOkpw/xaOIFvdq57Y5C2
URdCFNl7Wi7YpGlV/neWgofk23ZA7cC9cOG16eoPHwOQcmzXS9ZSWXYZZMnVK0Rh0DHGyyF3Kwiu
4bL3i6VmMsg7q1Dg6CulvrEMAHMa4FJOfuqItqj5POUSdruZFIlxZp7mEQQfYMhewJO/CCbl10/N
oSdUVjF4oTwm8ZJ3yq4DInKWxFUfsoX63CQaryDpX2+SFr/X5I+4ZEYfjnrDPRIVbGN85kyO8BLO
xRVCtr70amp1P4IFgbykCfk3Zi7jN2Few+xGJEaTPg70Dr/BI745nrQQ7yCD9Cr/YrrvdQUjNpH7
slV2XY4LF8bdqIsfruq9RKlCBNl8lGVRAtO1yZTFLGQJqibtc3maJIib3oedeN1JR3Zbl6D1itLE
fusqDJEs6ebpr0rwhgLVYhetISpPTgt1X7K/ZdwsBDUR7xJKK3YUqroJRfqKEO6lGhMB6ulSej6F
ijSzzF00EEM/BLEDZLjArgRGGvq0onLyLlg3e5/itKY85oAOdaKEf7zgZ/9nC2tmGvd0hJtME4Kf
heH+b46iKd9xT/T3YsDGIf086jzi1aKzb0l3nZnbqYUEZQmGxXkcfdmXGxrbXDZzUGILDRT5FcP8
5AEdgVsEEP9ILEwidUxwcPni/GUHdf1vJO4+0hktUZ+UJab6t35ReCBye65D7TPA7RHTTjJnRNZq
fiE53MXEV7J1TQY5ytiYoRKgCxpukadNjI+X9x4m0PM7b5cHk/U2tKCnJdPpLLCZS19zphaDM34z
Js9vxXFWlHlwmVRb8VGm7kWd4k+tK8vPhCU/hGeOLvCa34vrhzsg1Q0V86D5s7qvsE4U++v1A6T5
lAW+TBTjnMEszktne3OIcAJeS4qYMenySPjcs9FffirYULrqowNjrEnedCh9ZZGQZ99UvXZdpyRd
P4zIMKRjiQ7xRiftLJN6ItcefUfvV9V36NF2bvlgfYwxDuW5/S4shPgZFBnXDUlNgt6Kx4TZDGC/
htbCIvYjp5bHMbiAgEIxzSpZaECv68wDz0Cr/tqsMiZCTiJmmXy1PNWnfypoWdAVrt8byAB+0z47
MzgeJfVbddXG9X+DBagXOI03csFGrsdgJTPW1W0ME9EEZXajn5eHfS6k3D+qo8J4PMBt5XeVBXEU
zXIdxeOW83f3j+Va2YV3KqM2KbGbXOl6gRWzVTCdhXxsSTCXLmltRI5YlQ1YgrAx4nDyEbx78gV7
+4T77FIyhkSIEPpKUJP8RMee6q0sg7ZuwlPP4AKxls67NQgP3HcLthxF9EYr6cdPydDvg7sDAoDz
DDxkYAnscHw77c6NvRHtQJlBu5SLJFXUTU8zdXZDzKkvsvIPuZ1Y2vZpc3RZT26vzKEH/zGt7RFe
EYR4dVJFs8xyry/13lqcXl6BdWB2SHe/oX9tfIYKYN03HRiwdnc58bSELIzPAtnbsj9hJ4xspnS0
hXc43pewPU1pV+tUlgSjPVNNjH1LRG9StWu6l7T+04pakPh9rGvXWPug9cGOwvXCzFVZgnHSgM+y
//1XqlmURpeC3J/BwgstJsJ82a+Zw00vtK+emg/RIVbFq47pL54wmwmhcD7Zc9AuSG37+phlvE7w
J8f0XhC1R01jU8yMTx3uuFZH6A5cwyEp7fx584F+a6Tsnw/58X17sfj8dHTW0AqM8Z36ycVzHfAH
oviPb4FiQbADpV4ILdvVRKvYVAkjEclF8q4rF+DWP97r+cSkdKwm1AKx9XuSdw4qsbZVP7KnM/MZ
0/h7C6IM4LaPhmw8+5CA/C4vdbhvRW2wO43cvtWIZgvlIqcB3G0tGbBB1g5ZAGi/eItTQJAcilGt
pwXLfiA/Anl2mI/ups15EhNWVjL81STA6Gh8ekFNmU0wA6f4AJ/godtHrb6a6r/LFR4dYeLQjCUT
VmZEAlBbd0uvizGiUoHCq/VMp4MGcgoKlk6wKxsrPOI2Xw9ukAFu4yZ7dtdSw7zc9j0mldMSkA3y
qyzNLlkB8zlu/WuAuMSh3CEIqbFRUoj6DacrBZTxKiaaR5TEFSXijRZNCvuI0N54l3DMH8BZy/T6
tNc5EUDFuDLBdrWI7muWMEJt6S8k4aKhkH+uzGzwSaHj7x4ZsEZ5prN/A+l8Yry1A3Pg4jFCCE/W
WmKntio34TNTxmPnzu/PGztYi+M+7xuXKttSa3MeD9Nrvm03T7ebpXXWCDwMOT0Q7mxBcViCZBgU
F5rqR7IYMTOgsFRVZH3gDeYzxLlkMPCQj3DUX7RkehcogugBUdVNvPdEGHliFjNauQ/kJTEi+0Z+
Cy6q1G78XZgLFtXJ7PPZM2FNVfNlmRS+OVKdiqFbeO34ZIrahu+W1Z4V7rfOnbPrcIEj4vi4SqJg
88HN3Tzz1zzeVaTw34sMfUWO7T5UgYGe2tG6W2u+fnqngClDS83l5ziH2wuZkg9lR74v5yWhqMDm
J8HEdq+Jl8oeOTneUzF/aPUsuFSAa4ygyZ1QjDAQgCPSf/30nDn58U/Q+64d1NCT9SyOUHaTo2QN
tdl2w9giJVrdF+RwG319iGIDLdqcCCoP2vHEWY324FstBtOKnfohyPVswvV31Gs0PFX7Fzi1Bjue
fslokpe9fBU3s3o6uPhA+CAR1j3Ujg18754ZhTe5UbGW+MZrcNeuZQNZIfbRddmShoy870faTCGr
kvy5MMDGb7v4h8F7kMXfX2jaPen4iSQ4BMhyiwVAuSJC7uSwbQE3pKAcPj9+iGDXm76VOAVBJUm1
Oupb1PDo3M/akGbW15nSblVpRH4U4mimguCGibBwCwVgyYTxh7lJF8s/bkv2W4wthRjtCWeHBcEM
JReDzeB6KQ8ugcIdsB9GJblhSTfFSNdzo/kZjRlCbSvcDo8auK5OaGtNoznyHRC5DyY1Ta2Pb8I+
tL7THj0RCk8qFGV0wwgJZEHA2GSg8v5GyL+pmlEmffbOV8dSfYE27iPW72b4u/IXg29ugHlJYpTp
eqAGGNfiuS4X1sLKouJP2wMMVzjXz0mE5gCqKOqhIeI0tVGPpccJPAgPWBPJRCjvJnabV8X2XLU8
HnpfvPJ9W1oR7wV/er3ORQ9ERTsZ6QcfkuSh4y2P6zxvqF2xKTlM7p3UKhjH2vn4xEPiwLUpq0FF
Qn8Gg/Mw28zjYKP1gopkI9H1oEvudY/6vF0XPL3YoC5P38Ca7GLjqrOt/TuNuOrQJ2vXykCvVwAB
TVNKJ4YhxKeEjdw1lVO9/OG1DIeu4e2ywKMcakYHdJGM3Ij7f4yKQiiiCRnYTxq2fawBFliXAm4z
OzCNc/NpOp3JvSSGmaHAYJWqWMNi0SY8zCm0OzQb4OMLU9LAtq3UVNHAHkTx0dWvfvDp4v+zb0dB
5LJTppKUZIpJcImvCjK7anSY8R5HkWUVSjwmYoEZcE1lDG/gjNxliuKqf2pvxhAju6veEcFq7Ou2
qVnOUU0aWueFyrE7xgPN+1Rtm1fmRWgldWs0Auh9aHRvDZytwrOK6db/Obf/pJrSzxYMS9kcp+iS
6QRcHpKfbzM9vISIvfqgC1NswbwE0KCH8dzHt5M9ZrFVwEkRakVk+ZC29CiH+PwbCZju5YnwtziX
48u06vio/nIp/PjCa5au/p3wQPlbwaioi1bH2JegP5SynA0O7Kb9TX1pBj+SnaED6p464vIFv6tw
U0XDkhOFICaYslLgfX1H7NsVZYl0LI6bLyA5lT0rNdcLlZS80Y6RNljpJp/TUCOLtXyDIwCRtmLS
hRcUWcpzHiqQKtl6PeOb25Pct7FRq/E92ls4bhSgx0n8OtuRkqBhh0NSKd1DCeULIHhFzyoHsMnx
C3R7275fznHv5aA7T1SQxN0Dsgk2Aex2wDl8DlYHFgqhL1E4yiMQMcHZIVUt4CYcHCuOTzV1fElB
CKyml92UQ6iUrcCKDKsRjRmhera+D+JDAd7Mjy0rvfR3SzmP/OJbkJj3dSAnfi5BQR/aaVkeOG9b
sVRTNlO8FCZwLk6htRsgc5URZJzCozCrxSA50oIJZuKhBuN2muBTmQLnj/STiA6yLO7kVXlxcBIS
ZtxjczjmwDjjAhfsZhG17G6hIK815oEf3vX8IMum3ag7WATHBXan1yWVI30HJAPqO0Hf89Zd0JQ7
A8RTiI+vtG77QkteourPAR3rEd6ajXDuTzBBTZ2wl/soUKm+aIQ2B19/gC03DDp1PaiGFWkH93ci
EwVwDpbsjNOXMGXROFU3lxIBMmDw+1Cu61480rDJtVyuXv/tJgGnTvVYodgKRE5nJsqGkG095mrI
4Uqg1xjU4gccD+d1vSnXNqmfW68tNlUTV3+rd7qkP780zS3jv7wAhw91Lv/hGPN8dYiwVjLwF1jV
mW8k5lzDQ6uEG8OEmuIUk1vDYA3KKFzmKBvUCySIUGykUqAKmY8BvTQkPYsPYlpoU/L20IM6w68E
Goy35GMvDlTAMteFjra8UYjW4y86eW/YVUYx1nTs3f1MxTPAgHf6jxB+3jTiX38p/yrwsFPPBZ0I
oWoUcXh/Nv0VpdpUIZGXfSCEgSK0pkxEyy6b/ydklh8rhYS33uAb4KkBOAgVCEgQWyW5bfWGrPob
ADXSvTfoVG/hjtepZcXJfnhabGKtPChS+JGa/n5unAkPDrhUqbtJGMlcxBRhybre51eJb9Wjny1v
L/r10RXBe57FxoOESqYtaVaI+PYk/IpnyEW0EpxL7B3XJ76RZ/q9Oz3HYC0q0COR5UYO1zRgP+K6
b7Aga1B81aNAw9qDHd9K6qMVVIFKiuJY/wt5oI50Pq6V/1zGUeyoPLbbqYbwp1fBkc+8lRhwK5sL
NW/eDfLYrx6TulNXAD54LonqIRVIbJuDXisy9MRk6W687WmF4+ccH5eYN+GB0o1UnxjNrepvSINd
GV1hqHLF0fPM+HOPKhKea+nuHPVCobr6Ua2FJJokePywLF0zmFCHpPhSeSBd57lIBZEj+RlfS4yV
q4gtTTIYp2+BwCAtinedvumg18Xz3uEVdX9nwFLRdEXahHGWmn78S3NE6yo8++Ru3VLlkEOHSs9i
dxPpyZ5lV/20G8wDB/ogYQGK3CwWwzUhhvYeAA5tduGhLaS63t+obPzPZclHFtqsbx1t9191Nh+T
Z4f23wQjR7kF71o3WLT54RuKXpSFnZgUl+pRz81PGLwF5hmBdPmKLy6TL5wiOAWhsKB037NWtT4A
Ayn0YH1ZUDgl/YbW1oVfzBWylgjl2z0hfsn0zfxbqF+2BgL0chOSkQJoNluBXsXsu83tRUQmPl5p
2T4adY8XWaCO+XI9uSn8SEWUEjSZWYL3H3c8aebveeVSNuW+Dz1SGHNjKpK3eeUvp9xtnjwXvno0
sFQkO1waOhKYvn1OgE6saTky9FyBZIxZNq7Mp/ODyPB+LxxI4TnYSvAodD/aFe9Ug3jlJ8wmmaP+
aHTavb3Cs7zit8cltIeAE9hQQdjvo5OiMa+L7ySsJH9osU91klcWAi13iwvrsy2Zj4lffdrHOMf3
GZOGP4VVE9+fsxa7LZh0cAF1sklJgzqP4vDc4nWmZZYaOcC82bMYCBQsGmEqJ0cHIyG8FIDEJAID
gJUPTnLRZBYQ3a6T5g1AXmif2cmVSHbLzxr+HK4gB4u13dcZ+3kqZvdYP86NpwFt7oJ2fue7N1BN
T2lmShBfGiwa0B/WF7870Bai8vebWe9Uhg2FBGMxbakFudnPFn1S+r+4FK50buE21jBKaVrnJftk
pOzkNq7l+NluzKOMajopu6cEQD4FpZUOYz5L3uXto8xJV42MJxgIcB5O7LI5xi5MeTUmXaY7YJKh
xtaPqwGyiRDFIlLpcR7y4LgZBboOBfZ1wWmKst7oxf6epCbWxasEvn8h3k4Z3nkN0hI4Yj2l4VFi
tlsCWfmw4GH1h4ZYlydIKd1Lyx9P9eoN5j7v7AvmUK1VP8kgOxxoYu+VuY7MCbu7jSOD+t/1dFb1
LEMu6LgsOQYH2FmXYBj9bjo9OCMcEkXIo1xOe0OhZyq66clWYb3Hsh6fq+Ht2WZx/vrL08iJXjHM
W2K/JYP72OJTewVQ0sNLeJYoNDGsth7w+VO2t/O5nIItofR8i7n3sTKnM06RbGUuJrUm6RDLsrFJ
lPjgut4jnGvjpY9M4U0MgfoeHge922jGGF+yOGalL8dZ4HAtB76xYqO5wOl1bxHF1cL6ny4L+bg3
tONvf1qYU8mEQuyeQEfF+EVCOUZMjuXXC7BjIVAMW5HVHDlPles0dBPSjTOOf3cWO2h/cqPyK5Kf
u4XsMwg9X6sdkpo4EvFBNdU7O6eOVxHQM0dNLhuCQw5mj0QVDGjP2OSAp78C7isdnHLaRdlkatP5
W86PyqBJy5pNMzbGZDhSGW6rk6/m//cdQhMECMJlgF1sG7+/GRstV6rb/oFXwb+WmWzvSpNQW9Bo
37LCSrW7hJKJKAfT1Cfw/qI7LjUkMYIFTBBLLcY3Jy1Rp1owL3D3DkQafOrYkaTQfkCzchkjlgPB
PxaJXNwZGkoLj7qd0/LriGkjC1lWwl7jMJD57CXgU+QQHLj26w6Hr9N3An3iTRRX1I6157p9Jl3n
6rhRZhWEN3ngEELQMoxdLFggm9v4+XBqwLEGoX4mrresrYDCsFz55tSu7AQuIwqF3eBTXSwe772n
8dJ3R8oMUjS4mKrbUEuukMPO964Wgr3CHS1sUzEW6GZyfha2nf/pqqg7wzw7JXOAhPgT1Ta0twKg
AWlIOYLH7fXiBTw8y4ac0OOoMByetXG0gIolui05Jpb8mYIl78LQdNe2H3AselM+Sf8RDWt9CxTq
unhYKWQXuFfYJdmlUSJxsay7phMQxRDsMRe1rhusQDMGo8IDmHAhdN6nbBrN3f0wNyMPYvkKTGwx
tQZIkjZz4d+Q6RBpno8bFGQ3uCEqiWymiedRQjhFBLk4XmFYldwTfExuxWJf5BWzFUTABegyPFxQ
W+t8fRQmM1JkmKfGubRG4zXK5QAM1nDxmDLT76pIfcQGDJyBo72QlH+u11thOeFe+kxYMvjUdPpq
2qyE0Zba7U9Rl+dxsOZJQ9itArCuSZFnyy2pNzibmhQydsFf3+hv9GtHlrq9YCeeNv8txUEUhsPC
s7JxCsO8fs8vURiAz3K/+OgjXXPx2iwSVSg9NKmI0iKoXpex6/+WmyFF/mQmh6NEtms63FhvUg6n
6zFHghwJfr9EwakerU9zdHabvenHIh+BZRhfV3SBIgkPgbn174BULReBTpywMEUVtawbnOiOK3ww
CyHVgPCpm05nQZpp+n/05t+wgHyVr7suDuBmxzwZLQn/lxz31mH3VuGKu6jEasu5LztJf2/LSu9X
cVzFwLC5zoqV55VYNRMiSX//6bacDrEsAYzF9yXOwf4yylpBiZ50jf7CEbHyoFnuB4RYqPohFZxC
tbJb3ghXkFeRxwDxtMYvA1w89JiDMlAtyjdBlPxDOH6BuVY3bWXVT0XcViDBumOW+RuchAz6h/Kn
HvEX0ZDen+p8pgfUH4Iy2VE65QnydTi+cz9npI71iTSCjN+4Yt9YI6x/d+q5IbUHOAuaawtJp4Du
qy3hK2Sx8WuGxuy/kj445a+krqJH8unlpGDoex4eNRKq1FhULfM0zAHJQ2t+Z3uu5hlLo976XVrN
dYturuCGBbLnRqqWiOrnQ6B8WBV2gR/LrkrTjjyD/4ZFWb4EIbUDSuKhHgQTLY+Jv41pszaovKfz
HkU0cVKOH+05q/8DCszErUoW81GvMFEVQp+GfoZv89nA/gwrBlI8HRkelWcAjuDbpqT7Kaph9AFn
TNOQMchY8qO/6fI0KfUGeshVgiruNvGOr2yTgbqhn7OwATQoMfosWd+bu85hpgmiD2w/w2Bc66cU
m7VxsxZRvNQATJW3KX1WxHimleBWJ0mp0Vp7FRcBRXhd48756NZxZbp7Wu3NtKDXKkD3RlRAHdyL
PqovWdRfRcReYAtH7AVjvEZSSe5iDE+4NNzvVV99JMjop6ScdSr6NtVIzDhErGMCG4rlFKJvzSuh
d36pqa7hTfMU/W+XUqnUWXTuB8O8bYM7M7aagOD4buRDp9qoFcE+YamHDFcjcjjm39eC6hx1wfVJ
6zxiYXXq1NHLTIZ+U3xDT2a6ZwwWS0C9o2wongj7NWy4jkPShUtzI5cmTSEeTCXzBQw3lKUpFcqU
FaU9qetOz7Wg+AMfl17lR1+9hrxiYvW7yKauNdvVhGUuvpdYdO9Bzj2xzYAy+ly+JKECbZnRTKwl
r8EDlqZwm5/3GswpQoDJN4rae3rUN4rC1kl+72/Ry9zMZrNcqbIavDfm3H3uV9jvrGb2p5Marim+
TDCEXDasrVyFL4P1+HkDczFY6lA2azW+l8prT8BCze5yhKlXZ/Qo1mXiD4919IDMVmsYaIYkvxHZ
QI3zGrJP7nz2myv/JAZxmWEkMq2qT0MOFEiyHCWroF2UWfVZXlhxAAIbsxUEzrd4HazjgY2AOvA3
FGuGyUlwdmhvAOQpbniYsNgkszPpk3CHiFNd0S9+0KTs0QyOpHdpKgXg6QJtL5kQDt0McCOU01NE
yiUUnQosLLxQDjT9RYwiPk3CFgP0u04V5BY4sZvfAE8tbH4c3axF4bqMuhfc3byNs3/SGuwHSSk1
a3BTnwupUiDbs5FOnqIFQAfgTTzdhVHCZVjjuBdoohLqp8aylT1bTYRat6TdDd2AQBijr5Jcb0J8
ADGJag++Wer9dtjt0cLOkH+hZlA+i5WCwkTycaykjW+vf5uRYye/FW6R1cK4nQYMS+PwQ2zE7TKH
dASyRBF5IbPn0B6qKvz+CVAjTNqz59Y+ThSGe3WGvLQSqZjqKKcxpQpHc9kTYZoP39hvq8XR0heC
JcULRbGASuWzso41ZNWSpm7Ib1kj0ZWARlcgZBlreB4CcnWiy8xXFaCD8fDhqJwsrzRLDOMDdLJO
wn6VXRo6o5+JkIwI5YQ2+pUaK4oS3ujdCtRPowfVrYtOhPHz8A4YtAdg1PjqmsZ6Ip5YsRAbYCyC
BC0bzBP5mNETJkUlCF6ieD5xzX4OWGTl8jbdtOhAohQwa/58gUgRDeAojaROx+ovNATVwiiGxFSh
3FGNMkXhaApzF/LjWX+L97jE9155H/gzDxgPL8gCQVAFtGJoRDvjanT0dAsC9B1SVEeE/ZFW7dP/
56ADOdHLhXjlhypC8k2SuphUPfsWVHHGyghQj0MYCgjJMYr8K7AWxPydzh0iWkQwns2H2wlI5khf
p9W8Vb2X4SSAsMXAeae1Wy7zIDZOFqJ86xI7Gzd+X92vEuaCfUNtO6WiYEX86CHVAglM7Q0BFbUN
AG9g0CftTOjIZxoHY+PtNtyFcd4Itc2WosEbixa8KZ+yfN0N2ne//xCaf0McXZLIh2rwVQAhMmzn
9jIueYoPrc4ZiqFDx8xNwgKVR7WqegxhZXiQ4QGccIst4yEUpDIKoYdSqoszmUagBrXnvMhuyx86
rsVEVgI4mYBjMjuUFQNOAxVDLm2RiNQNEBczTcJCfy0Xpiww/XukKdLkCCjc+ZoQ69PyInNoLeUg
iOYM5Jasg4e9pHmgWwHXAOcu1mmYQFpI5o/mitxkop8wDpohI/6Scs5Th5IuWJ0HncEftb2FTiI/
wrlkWSlLQH2tM9VoZ30rNQS3YXCa1XWEyXwSMsBUPHZTAgUxVvfCaKt3uzAHCElLIUNgpwGDtsXl
T4OCUqzp9Nga34+geyIARmxr8sxfCch4T8g+fPDvQ9f6yXdzt1mfmthsXUqUiMPcXTe7wwS3IEPr
wdvwqgvQXYQ6/CmXFHDjt7rHd93PBz6VMxi6TKnwJzd+7PQzaUElE0W3O548ZEm5oOpOpFbEV4u3
Nl9/Ph3AwUxorPqC7mMVD8A12jc9uHhv0T5OKth3Ev6FTa3pQW4Ixe+qnBXukxy9aomyKji1jV6K
k7I6Ih3CdC6Lb+lYwwS1N8Q6doSf1gH45UpHb4R4iYAB3nly0l1IfVO2mUHMdIuQSWOMHaoUVsAi
0SZ/mvo0byLYUbK51Mo34h9xLBW8+t+BfKd/FotkisS6uZOZy7X6gob7am4kyOBvfE+1k99zkH8o
jtQDtTVgFXWd0lp9bzuBdmIiKNJwUQ7u7EMMF8FOfkmTPwKC1UQO6qxRSbhAyo5OrW68zkjzOgBn
TheKo3xYgALQ2yeb6TVec4svrN+gvAg5DemVEJn+eoi9aPCTwe2GUScwyGLErpi7+C8biVKuvI3w
9dUItxmIzIB/6ItevZm5ZyVuyfxY2MRjfsPLpap0EWtvp9atavABVPcZ8k2U/B5SREpoZt8DvXdA
Bu9C3Uf4zqmjOKMsf2jlfR1Fe23wTXFU7JlvOphZBwhvyqJPfKVLJiBGkqpjaCTF+ylD0fK9TDXX
vrstqRGJjpx7Pa+8HLQ2obSbJdu1ZKZTIMz8deoL3hUdRv6ZIDUI0kxjCVWULoBaOM49Y7l7llTT
ND+UtbMHcJh5+8TiH29BcyCgEncRx0USFHZtPMZY4a0a10//Q7P5AhtFMAc2wyTpDppnkH8gFy4N
IRDvlE8WHQsMCmlzu/6Q/rIwEV8jdfXpuJgkWL8goUbe9REQEG+K+tHrzMAsfW+f+wGJ6pUygTNo
Ia41tEQHy7M2uEU92WjYNoayAzMJvb+kCYYi68CZULP9VHNoKVcdXN+mjduCTxZIjNzGVGAr5qPQ
NvOnbII+KBYb8qeoqFrOsldZXNOIQEQnh24iw5SMCj7G/6B2zgUWlA05xHbMB2NvlyN6Hf2m/TTv
HF27yFyxlLJL9Bwgute5wOvTNPTXnlS65YPHb16X33kb7W3bvj41mfZgroPGvV3DyMBu7gM6nwH0
H5lh25Tx1sGxF1+837Xd0TvwstqjklKG1p8NJlkjVwiaQHCZw8SH8mn1i5vUXOg8PFsPe055Ouqh
wwkHfVjNrOTnznwY17Fahk5pO63IcDbTrj2rVYixPpwWf7iOfrtlm28WVE9vAg0I3xqEMuuKqg8t
5OIP5iQNMONST+gsi6DbtINUCXmJLft8AuGH4H69/K4bryXk49m5K/yhGLuIVf7aJmZcijy6CMnR
lic1Z+r3VSdFqW2BEoqLfkGP5mVsj4d5L9piG8JpOu5zWJHt1ZkOby7l09fGVR1J2tGnGLwNyhHe
9HddSVm0FVejB5AezLxIxSuI5G8OuCyarfgyO6D8ypXE3lFwxoSes5yXtq44RUCJGok9Yxm0WRTt
0fxYS/AGKSfJKuyn8v4RMUgOm+LPn3bipIfLjIX/p2y+or0fiXWL42VgYZ9+f/JOGScSbXp8FabM
vtr6njxCQMZ84Z53g+1MAvnzY62t+XHMj6dJt4Ax56mWyxV18Rj3pmDZHikadxu94x2Ggg9pnTG4
sYffnsMYFXVACltIFr42NZyddkWo78QWG7DtvTJhgBGJLBGE1L1IsTXXxHTURtF75Q8wfGn5lKDW
710cdPfhI9ia1EEQYU/RAdpmlvdEJJqO86XicdaqY44uHRn85cdAIZ7R3QtDvwUbwxee42GeXRxo
H4aHMpHNfCPKDQNDf6R0D3G4Nnvg321MANMxZb5lkOAfL1PEHDh8oi0Sq3MFa2EjhbLvf2HjG53n
ULg+84XEXMSZbAgzmEY8uX0bYCmTCveggtWldJXLS78I2IjMA1CuV3X5PUovM6OG5biLCFsOJ6Xl
AurnGFxxpoRIBd5KUaF9a3RVw82M/ygtuOBufDTcJO8MMSmpe8aRt95681uZ0rhtA5909UJn0sc5
cRNUX1SE7ExssdSqtEQwxBPIsCesEyr6196hExin3T3TukZl/NSFwmrVKHsbw5dqOs9ZSxD+q+bm
XlbRFGJb309Y5xoaTXeZbKD3f08QVLD7nLkAbLhi4MAOu6kl0BWpB9V3AqVhVx/pU1TgZ59rHqjN
47lCSb/vnNmNXbF43csFnGT6xZIVKOqj8SerAoxpzrDQwxanNC4HDErExHpiTZspRaJy60nsL6c8
pGHf+UbJMmo3uT2XkSUd7pugfEiSTmAOkhN7Jc7EOUMNnsW/VAX6IohzIr+kxLk2HFbcEbX9SpQX
fJFrbjDtQjP2Iu0TwE2xczyKyjyNbjaMdxVXmSkcoh5WHV3ASfsoleCkhdWzcpq/XSAwvUvUPQem
f+pIEjOuRTcCiZ02eekuqlL7DAaGCO8hR2Ex90jdIZNDfnu9zJxgxSFyozEJ4emqxREjNkn6P8CE
m0WdPP0DFfMqk68dKFqyl+W0KAPnTuB2gMqu4/oHhghsUl0QPwPilTTtHIwUReB873obt07eIE6b
d0L1vPG31/L4ONdPUMYTwAVqXvO4FG4asRX4f3awg6RMT/Z+X2OowO4lnXpqB1QdGotqGIAzl3RE
RKVJytg4fptXYTOKlk+tXwpHjwh5VEqG8Fyn7YbSG2svwMfzSAlGBXAblLSC++DoQGrmS/+uhW5n
Jtxx6rxaUo82ju8oVZfhghkRQsaxftcq5TFu6saL215zrJuxSk30zXQpQ3mu4JxPHut57Zk5mJal
axhOHSsyXLdcqddXJXwrCt7xYpTsfnpZM/R253uYS3dcwHJrCLh+Qsx8SgXsp/VOVB6dL+h7tyMn
7PaRvkXTdma83lVP6d9pGN+Xj8VcV1Ox5s8wJuV0JIvzcMQPR8a3WuKeOVdfNezIYJuXNqKB7fRN
4gkFVNkzC6KYlL9Z1aL/wpu/h77np9VvlDP/LD6bWiIKyIZe3izCVP9FINfa0Z+kQd4iGNi4ftuH
vXkBxOsMqdSgMlgKEzfDOFVzjM67JYkJXl3ppijwuTsGLZY4DFlv82zfFm9PCbyJ3S0JxNG/j+ue
UCA6heunQfFmuN9iYyuTgLFgoXjOyzqPYgqOIjjzcC+3+/lLW12DcRZ2SGSCPqiUqRQQFSdbtwKE
rYAca8TJJS70ATJGRMZxyubKYHbG5folKPSqUgYDmT89s2V3/x1XKK6BNFcRNnFfyiEdjeGNX23F
ObBaxOiYxpHIGPr3af12HFZGeU8yuLy4P+PavBZEu9+G5Po3W+EJ8l2qtiWegQu88rrhdhX2J6w0
ndUg8BOVFnmdyskczznYmxWtHerQXIUYfe+FXZpN+ftqouVPxZamv7aWpeyP0I0dK7i6kPwKfKHU
TAYqpJ/IYh4gQigKQ0YPI5/VaHLi4F/kU3Tsxu6JxHMbIyO9dImcohgaNSDW1GWEypJdZwWmeEi2
KvMveisJ/79MPBRHae/sgJKQlK6IX4sk+RCHBSPMx3NzCY2EHi6yWEnFqerg+h7fpq9ILUCHAOcr
JgkRoxXRs8/XW7D4waaCsw8E0i0tbLzutMf76kJsX64VACdPihWO4e7wGG9NvvYCH9CEretssU8W
cjISOChpSrf5mpV/95P8o2QwFb3XDEH/WQhD5lmqd3PqRlUJfIfifzQ4ZnTUCn6PqDpWKWWlI7tG
MwB1Yc0XTRV3N+lN49akhQNclNpdg77lQlRPz6aE+tQp0x63jIEq6RGiEXdNW8z8cWKQCKnwF+Aw
UrAbq6zh5dob0rAI0Sar/ixR72LByEfIs57oQN8P/fCfSBMvf1p1x4xlbsyyaVGm3ylKsPV0dy6T
UywkK1txRer3mChlQ6C+R4YMPuyQF2lMf9kJtunMfpL/fjW0ufWrevIK1BDkJKYRRLmQ+Qbd2o/g
c8y7ry9S5Fye5szaPDuOPn2g1CxBkUveRvzg19+w6JM0a2k8fIPSsEY/qwUxgYgzBxPvyU9csv9L
e4uOeUWoYg6RhqcuqBRZMtcGNCe3aAincoT586usRR3t67tggW5UGo/DQossfHC3B/tAD7TAUGMT
xcvUWYeRmkDjmI8cPRl9BtUJ57uEuJDHXM7FBxdWoW0/MBLK1eST/T4OgrhFDrl756q/ORWpD7dS
5a4Ei1uwnOkPvVGQ1Oc1cPZuQB+8NoqyCnyRVHbA8kXZgS9zLLRp9k+huvq/3T31kdZSO4OujYPJ
1OnsWyqmK+LSZzPNmxk0/tTA8HdUUrpAWjBRmhyEmXLBwlh06+kQw/Sm7I9oLeW+EvA65GVJtW1/
ndXffuVhUP9SCDzJapB882RipNTd7JBBFOGAr/PQCHUuTPSxzkc6rB++hiRgW+Cga9WGyaz7QVrR
7ueNtVCQnpRg9p5OaTPTcGoJdwG0L/Ebf9s0xITGLXAl1JpFLF5Mrafx0vPl5eL1IT6HgYAKRFw0
34+Gdh90lQkSYeLSNU2oeBkVVAVkk6oD0S3Lk4Yc0JoJT4OegaeXb7rAuslusRonJh43wtHcauKW
dExml3dKov3g7Sc8hi7jokWLEXrwmdlBPfj4gcNkXxnXwVaTi2BLofXS/kfrffJNrAEwjvK/oXwR
RELdfek53oxn9WWkxoFzhgAlyNFfWjuyho9YrGWjFjV3zZevmKM26SVZ0LQhHU5jwgLf3HOUpmvK
AAP0OcZLSvFJZtET5UGvqfr4jQDzSrltUrH0/mlxj/+9o05dK8RBQM1bPl9GL6aRv8mAaNd+HJxu
yVEWipRpWYCdoxZUSIJcU9zsVJLU0nfE9v//lvkalYvrH//7O1AllFtFa4T/KU4lqj4j4b5J7D+d
bIMl1PJWaQ/najGcbdZwkhlL0qc2IsDUe3Qc4rgkt6kYW510sILjDJZL0xdzFCzcFBzt8w650j9M
MrxwRCDWlYJeCFUqFmv/6eGNRJgqpaNbYiAUnP8HrUvaD2mpuM0Vc5gbTeAg/HKojSpPC9zUKINO
6iXl3ujyg6h8GtYje2Qs8wPmQNya6qmN4ST3ocWzdnmrHYTMmsw5uMj+QZnwR4OWF6FqB3H8wxCO
BmInnyIGRwTg6M45xUxGv6F7XMleD25brHS/xHNYTWZNc5hEjSlmxgVwR2Yt+V1k1fVj6YyWiG4g
nF8thZbpFiNXunD71ndcpXfLzbtA8H6MYgt1e+M1SGi00fMidW5+omibohiCvzs99s8whNVJMvJe
sVkS+hTenQLW2rIKrjti5UB0UF7CtOzKbRJJinWbT/TbBj0o/4OPdbu6s4JQNQcZTClJAT0UaCZp
ThxhpWNNmcXcbTeeF7x+tzd+Bf1Qs/ABZ8NtcXtaShU2XzRjJ+qZA1KEQZ8KRn+bhJ+TtJHj5NmS
NddJQjt219nbPbKzy5R+T1jlQEIlCJ9tEbi61HfUqv7557SY21EjU9mRxud3hs07/apXh/6zz5gc
U5jV0sM/bgwM5PaUflBZQ1J/wMHKOwXbp/Ns6Yp/nDYU46ssImYJhPJc4iV0Y+ZQsESqPjHtzOme
ESYb5N8L3XW9ZZLutP+X1Q7HYSJYtb70oOJ6sm7S2LEbQUCPn99+/0lXd/MFQfhrZvhkpYBfbd2W
WsUbYQchbvPD/6s06cysxz1JNgVKZHTvKH06iXpj7RTUfwYBRx45WO16UfWwxfKdl59fSwR67Ogi
3d8NpccIcl2b44Bn4JbJZKh0NS1Ds++JE6huF1G2Ho2jk3gGu97mJnmnHiW5FMPplOv5VwogEvcw
ScEQIbEQgWWYbEkcwkSGcMepYUXDwHUja+TVdAc7iMxtRvEnxJ58wJE1syWPQpAfywAJnP5CczSN
PJKfILQJX7aKtVm70qHSJoYcgD0EvOuiLZyVa6hp68w+K4cQ29KQbn/iGRVlwQt9hvmwnyHgoF06
+NzlyPH3HeOL3+ZCrmAJQDCc/q12Ad24g90CicZ1kO8IyT+/dXRokb9TK9Eq6H/9oe6EjTeU4YXU
6eIzGU3SdVmNZ2hgWxrmLK0rGmBYJ4F1pLuDjrt5zEvgUrIOBwdhMrXJ/hADcu9QN87p1CJJsjsm
EbKcgAtMIMAILjw1osmBbhWddSVbo4+9e2Yhit+1PNbtfjxe8aDjEe5wjoco/beT1b0bZ2+BSfuo
WLl1H3oqkRxaTNIUmp+UGMd9tbAC4sFP9EzzKCKW31nsNmhr+X2VLldz74XSgBJRfafGayMknpdk
bWUJWX8kyM5KwGcrcblvE96w8+4oDQvsJGVyuOfUWxr/i0qTB3psQxdvvDKBlokn1DL0yE0yHiA7
LAagtlO9qLB1Smu8l1G1QW1YRwBqBPP3esmNTQ8yuVADAGVjrJV2VUPwQHKGZ97Zd2H2SW49LV2D
W7yMOrqYaIzmhSvtP21XXEQ6g2M7C1FQS89aYCyugVj3sK3+ztzLrKZ2ZJEyQYHLrSC4J3vggJIK
hEjcFtc0exeH80+v2h0z5s9PEJhcUBaNgH7wh4E1+OLdlFLVhXT4eBdRQpc0ogyuyoefT5D4ezPQ
4o/xehYBLODz/YpTRNWgr2fUj6CLuuUFGCE1a3IaYPaxhmuUJY64ExOEbUXDVVioW3rgU/jiBKVM
cGf/Xu3SUmR4Y2iHYczYxYzUIO1NV7WnRzR+2C6C/lqx1raV8cVA/Paya27AHafZjvm3dr9Xycj6
EEEYs9uyl61o1GDneen68qyIOnJbIPdzOk2ZC6ZGlxlZqrlqazYwYSsrmkcR7QKwlL4RvgaLyc4d
142/LYniZbZAGiYqSpoEAU+nQFL2uMN6o2RCozI4dNI+x1zq8Rc4vNckS9uJ+pXc1bVLul3hKyd3
46NP3tz0YUSV8JwP10BQs3fSqcDP+BNK4KFqie04Ft1+KrglIH43UqIJZLM/5ZuMUj7WSkVOCONI
7MNa6XdXqSn1bIdc2m9UciIqbinBljn2MU9oA+40X6Oo+KUFMwBArW5+Z0hgDkPmGhLVJVq++7BK
NByk/wDrWj3MA5LcvkiKjv0eSAu37xq88E4xs3tGdi5wow24E69rxTh+9lnzKSWXWF2JR20pHTfq
7MgjHFSqlqUXr/mB0DrtgY0Y7q00+CNYgqXsB6G5Q8hyQB9lVzUfxb5x4e0rWGT8+Yu3U+N19PBX
nZWG2Y0tOgVLwjXpT+1bgx0VbqRSvKjJyhGgt6JT55WRhpkM4kvgZsF+0izefie3AHdS0W1VEK4M
Wi3sG1x9OE1/B5LB/YT8uZTVwBgcb0Q2RgVih/btdgMX8lroGuGSv45ZTyh3oAXQkpTWOYK8b9To
5zlKSWpZqE+BZ8gQVE0twDYsySdBB7Rx32IrAi2dnoACAJ+21dWq4Z4/8mmvb34s9n0HsVXFjm7i
bHx3PjZt0Rim6YJtVOQcG/urd3XMyQQjW9gcuGygtyK5fC2txBmvanxSmq3JsGBjP3sXwXWFzDhC
KQL5tfBFRi4r23K/ym6wk5Xh4CMULotbunx6GVkc5Tk1GlK5fa0qKqa3cY7uX2LyJehJTqH4ZrmQ
BU0MRsciQb6qS4S0I/IDrYv68Q6M78zwdJxqoLkBtUx7ipuH/APAeZlCPi7rEOGsHapTV4Wn6exy
XriiL5SAG1WP8bBlNfuMaxuDG7GJOFwHzTWFcBh5LYsLlqhuIG1S7RI7hjivGS4UeIjroEb9hTDW
Kjl1Bf+cFHJ3njSAa3KcqgxgIb3sSPMUrR8i2TkeclyCH8DnVzRVM94yN7ZSRjLYA9F/Wzp6uxNW
7l/JhMKWtlI71WVms5742smY0twhC9w3Frx12V22GM7cNRgoaj2pWr2Z3CBwvftuqvQvIP1xH1JO
9GnuGKuZJ00psg4c2UMgk8gT4bc8AoPBAeVW/noEvbHFHdLJwTe1M9QRy7stfQEq8nYGc485e7oI
VaZKOTp+/Lt8tg8sQW3qQoSww9yH49ujqQurWfcp4Z4tSRlkxlx2KlQ4JhTTefi3BM39yhOb0C82
XlUqC0C18Wg195c1pCv6GbXZOBgrxOBcQMWn8BdoCRoczJDGYFJ97fUa33uIUxRPgBNE4pU0AyBO
kFaLHR62mPxW/daXYaq773hw7WqoMDgF0+whOWDtSBMJCcQERZPqQ88s/FzYBqbTj10hMBs6S05l
j/qTBz+Gn6UFYufWU3YW69meMAVf7vxtNJ8uvcgHwlZEavIx1bIkCM1IKfczehGF1MKG5/fVf/sU
zhWdyS82HA69LNK3RVtSoOsJeYpOSUXdGmZH1NTyzkoCw5rm4TF22CI8emKAaSaypv9BGFhdkk8/
HPLgSptqVRq897cphYaq8w64KaqSDuoU+4FZ5xmkbhdQKOZbQnQbx1yW/PP7Z0JgQRQos0RNfU9e
Ovp+5jvoumV/K/R39WJLkW3kqfwhnYehrBl0gc5dS+2l7SkYdqc/+EcGVr5am6sljnFidhdiK8dz
9N+m28Oi1+trIiGxBPOaqqRDTIqPYGp3T8WliUdsNZDebqPZgUUHIQeJED0q+zv5BRCc/5B9jZe/
d2D8NL0n5T460WzvQXaxWSUkSOFi0uZc+zug6bzKzsNf/ctcj3U0P2BcQMe4pgYNlP7N+YUjlHm4
rZMHnN06lW5mk601ZuAOXhTe2+BtUpR+ZUw3f1yx2S/2uvLoDo6roeP9+LjYomYcMSGFyR0syZDv
hSacaFEHR0cFMz8xQs/dJyQx7M104JdoTlh1oNzmNja+bPRJQB4C/+x++pSWabIRjnB0c6+iCkFS
rRW8xnuUcgUUC2hxBtuZ9CjGvh6CdB4to4Cd2bXDVA2bpWotFuMvxENmfqMdhwbVlNvdTfNB2lGI
Oaqk6j+leud4ADABMCxRpQTYdbNvGfThWrrV5vJshzlJHo6aCMRJNTP7xDdz1jwMNS/qlevgmqMc
/TZGE7gXbTta1kvrygMAhNdrD+ddva3Dd8pw4h1cY9vbyEMkeIgT9HDaIVw0/TdpLRUZkIlSemCo
RlKkjZp3GSift+WyZdri6c0Ll1+ANcXwlzFHnhJrTIbH67ICmhjBpqwc4AbTpqh7gGfYg1zQYeLB
IPwUPSuapkFdYwDvnN00/cWoVfzsikYErujw5RCuVg+MGk/JTAPFNPMuXGAD/T8BSZsgYreOtpcB
wm4DxZu0AwBIro63+Bxy3VMCQxMiYKRqUy7ftj4fqHPXf5XPNasDn8rqx286JcwC434SU4bV61jd
ACNAL3O7B3m7DNXiVcEGDJJWMUwvgMFD/p858qmEwCuYCEKc5rc8EIRfp0kOtNEHt33UECkLKoFC
DDax0iNoYrDVqj2iTVf0rlY2sfQ36Hrd+a4q6fh1H1SjwO9pdMSZqM6VsGAnaFVAeMn27uMf6fFF
f5QuBPveqEIUyEKspWurSL8EnpinRzDTJK5Hey2NQz9FV3KSXLWcCkoyRcVo+ne6G0GX9e+/O/UN
P1vXx90UbIlwUWeWvMAJW53i6DueE6AZ+owO46pe/3I1UG00DF6gdDawVoP+UghXZ1hcV3ja4t1E
kqobD5tR1a95HTa8de5j3HFTi0n5tYU1FclLofDfKBKT0MUGVfj349WXXNSm+ZA2J5+aIMjElwWL
uV/QZet9MvBKU3RO6mufTJJtH9deRQJhRVtjTrgJ0L+ZKyPAv2yWsrRDeTRWVbinCql6dSqcByY1
Wf7J3QMuuTPOoeZiFBiglakjOiCiohOFRRpGhKezU2CcKT5xkDIBhFNsHZ/IjiYveQ7rPS+4A5jb
U+sU3Lpv+AdH8xOY1C9ugidvTY6UBeIL8pP5WeefMRgMzEGDti/Picv6UbubXM6eyUrMkWvT+HT/
7VcwC/8vBlF1SIqkaUEtSByWqMMARgMAhGkcdiHv6QTVw0tUcrraD0mxmrrjRohS/RU6rjlZtbPl
LnRM2Nwx/ONBDrdGaX/2YYDvDKCiX09vp686LHPIoLD236zUaeRuC2wd5fLF0M30Q0ecS0V9WaES
q34nIu5D8PsJU74ltEWDPUSHcQ5iouFWOgPc39KG6mndo4o8nUA0lS273vkqclAfhR6PXvYiha2V
3X5o0ege+5ZX5BCaCBxTnDtUrdU2Jzu+lKe8Qcj5A62ptbi9CtCuAQwqr9X8VTHgJrxGVillTVhG
EUAGi85JMlTvckAnHE12Fd1i0dgVRoUj+dgfytbYd/8hLSxUaGsnCScS2s4AwkSTYMgrVNQtBsCA
TzjBpQuUDwMCfCqp3GIKzAXK9gEziNuTNl+qGayNx7CmV7YKq5rVYjVxYYwOX0K/G/vQR6l/MwUe
O8XMBhBRPKnMWJBTELAtKPgKvk6266WtQlCZ61uWvEZUepbA/1f1tT/Em88waUOGwzgKa1/B/wWq
PNequKlhaS31cS8mPIWrvUHpAi3voSrn+zZwJmOGba5bSDeC0MENWeCuMh3rKd0WmBfpmYSmaCuE
l4ps14lEJ72FUEnDeB2Ur2/UyB1vu2imWeThBbvFACAZCSM/bfbTiP5Igx9odvJyDWllHq6KJD3Y
F07oXxLw8zlLjZaaOWjC1gOqqUqSK6e8jVzcEDFGU4gUw/TYKFOLJ3E3wIdWvmx9O3ynozvXkneY
PzTGywdasc5ShYB7VtI7pNuziPg1YB8tou/SwKqg1Aq0gy3hM7i+cyMpZUT46HbXqvUB62/c5agu
rCPpiqQdFYmg/sJNVpqJBec6AWMY/E+Y6ZqMZspIz1n5M+h2dvZk11EF5PIUX8oUFyyQvNdXs/x/
LwLw8AIInNbEyMgERUmUFrRpdyHgVS0bYeA7KOKcVSf2AVED5ByU57LB094UcyYoATTn+ScCbHbd
QUCtPv+ZTJBfuzzmyGPZVLpD4TSbhmOGQQSUa0b2iAgUWI/odshEUThu7TK/uC+ZW9SlfvZ+wbMO
mLORGrHfkMiNhQQHlxbzhL5kH/s6/MiPEZebtF8WPOG/ALzOyedeWRhN7qeMxpv2iZKwt0hQDlke
lRNOOSmVxKUNERW+pmb4clqtAJk9NB84wp+18sbCcL7r3MitvjezX6YbiJt0H4IlN5tOzaX1Fu62
0riSgI9z+AUhEhABRe5YmhCgDqbuY7Mxda/iX0EXPP5DGof2VI+NyDF9fWU5BjhPCqj4fugKwN5L
0WcGpLnuMTLcph0O5cGRU6VlulqN0Wf8J7nJ9d7ctAVY+UiBoBty8IHF7jP6/GLrep62GVzlW2XU
CS55RqEbR+A8dJujbM+iTWpnN9+ErFaZcyXcBIijTmx2w0Pu3Ql36kobcZR4oyV5v27dENWi4+t4
Hm4T3RDqH4LuRLiKHR8pzceOUcEtYfFh+AlZLtY0lXftfBVKaNwzkUds9smVBRj1bluqjCklp3nS
+ASRIIyRsT3l49+588ixEsyQU4EGfVPJMdqo1WLBQPJn2VIpz7bpiFt7tRBdgXzgR6lYSI1U4z8F
iKOG8C6hUgKYA35GWQADh/PIwzaADOADXlJl2DCMv6h/9gQx9cjRk9prdFJoWt5PEEv4+E9CDoAF
cFaFiBw0JUESNAHzS07CBKec/VylUH1y+QVAgCZbRxqaMF4SPv5onthC3Xfn5EaHiEAkIkkXwShA
XJ4d2E8HhdI7dIqIu+Z8SQa0wl47uh4/BZdlMY93Q6ZtqAvNNNVFsXQipLDzc92wojBhCBj4IdL4
nUgHuxGOxyXm00USakdJ6EpDCgNJ+C55H+acWlNqQwvRlu06755iGH+04meESOoetahLpPzyzcNP
6RNv9C2JZL2bLlBlqEVDWSPEYRB11erNso6lo05skfhbYe+JeTYxO6LtOUJFDVOpxMDLcK0JrtAZ
9LXWnaOwHh3nZKLoFHsBEybAttaC2m8ITq11vBaniaOp2d3cCjnCdUhZkW+Arn0teTikG8g9qDQB
LQ488UOxGyUq3in4RUejvdCxj38Pluypo5f4Ol43vYnXVbKPCZNfwUc4fekFek5vO/qhS+MCSs5h
7pvcObew/n86v5rloIE12AJETd5VevXlBE907vTEs5kkGQjKf+ZrQuiMg+ND1fmmR8DvFjEY1+cO
0UzgCl2nP5k60fhdfSkGTMtzjUsad1wl29G8vsmkLIssQDcDH6RMltymBT1h0UcHaxqIa5VbOgX2
Fb4FnNU1UJEE5NWBaHfRPJUeoTXfD5K2hoeB/6LDbNZaY2Wx6QZ0+1Zs8cIDQbWyp+AsyYTv6Tsh
J3HhGq4I7USE9oNdbrT1MudtmSfCsAj8ITKVf/IH+lvOu59328Dv5sdnG+DcxAe++Do1mT6jLYbk
69McB0ddK5Y5ipaRd59vUdMMLikMV962AGlpDviGvbIEuhvNGiMAzsOajnIRrOdxR3eqjM8whf1e
nejFUMX0ORVvlIhhKkry4xdPHRETpqCBWJEscuA5YRejZ8D7Fz9QY91qTBIJDUdH1PbwuLpugXa4
Nz6B0gRSvlr1Y0f2FsvXa8bTC+kHi+VCX5FmpQSaIDyDgpudmPe5eYbAPJHxYHBUF3u0poznCnK1
e4XeOhKw4jZSqSuMi995/6Z3D1jTOFJMHpyeXq6YRDh6I+7T5AkW2k6KyoeBSLRIAePZ//nQZdns
ahaH06GFnjXPy33QALFrM/JQhVCqyE8vg2WoVWvIEv1asgYu/gxTj7wqVY6q8z8R0+5VEVx6KoGP
gaKjqR27im3iBlGYsuuDaDKhs0cFKQ1kOJIv6n4JL7SEns6eoUWqItPbEplgzsX/50RSGvqxIGFs
Vkehxh+afQbi9S9Azo5t4a8xTFLdql2/61GxZ5GknCEXkmSm0nWczaw+8eNiHpHv6wp1SqPOroCG
BeSVjTyn6iwC3diu+j8mgFtwiOra88b10psEvodpm5NVrq7GlVXMt028aNO0JWLN764E3LI8Hk28
bnnxgxQbBP13tAPrLDHnFsWQPIvM19lpa/DNX6+4NWG1G0I/wfF84bNudyGl5v7w3FbKrySCMC5h
KqNJWduci6FdMdD2sVFSB7mOCKdDvPsy9WuvaJXPRhKaJ+a0KCUlxIfFiSCSi/gUnjLSl0c9ro1f
QnLv95c2P6BF0n8g84oqXkRDQORCY6FOipbc5BJitbXV8Zklwt9e1CCkN0reYjljqGJ93Ceocs3O
+rNPdB0jLyBiEnSvnViaQoSioXtkiTGq1CxNd86ScXODDypC9q0JXudq/JIPOEJ3gWwdkLJaqsIg
BdDDsZgcCV5ceVqHINFRp1OiYWA6ZtV2zkBeTYl13MzeZMgPi5IzGI6HGKbPXPHIuuRMIHPWMOdy
72zJVNBixlYFxo9RvSa1bBtDuwurhn/cciQuZQ1i8TdL/CZS0cwBZY2Nu7E9G2LEIK4PvnKKX9Ct
5NVnCt/yYqip5nbTIP8PzoNucWmkJIV1grlXen+QJkqGNhG9+hSYySkk64UjJCxrDrYouLW9hvFe
UJ5w9gQpejhzkgrnGPVicWfx/WiMUF+SF+5awqC3v+KI3UdH8X5smEXa09ruHfQEsQxmn29FRdvV
zh6r7Y8i0NjfV4ZNvSy4M6duqYIvQq1i72Q/hzMfyvcNrmKZ1mUTap1F/ZFOxnRbiuKoQN8hLc4i
1fPrIprpiik3ZYp8HgFX2R8vt4yELAwSqNYyFMgcyXxGtJu3F82MPvPjcZwXWAjmgE5ppcVy3fLp
ycyxviClC3c90iFfZq+dfWRfsV+2eiKVsPfZNNMK8bkxq90MxczSTsqk34re1Xg1JFQmc5s6TFZQ
co4nHONXfS/J0y0QYhK6n6PTgNy7zZfpODQ0HuTFqBBf3Twf1ZahmK4dwFYiQbsIh5fFWkrHUq+i
1c/69WVIfr9X3sso27Dx5hEX/PTXNs0u1jmNR6/+1TYhcOl3yD1jDr51TSUV9NAdJyOGc0EK/4Eo
GdX8FxAOZIdPqXLtsbt8WS9GygygS2lmnkAp/R91zikSOKI+HMFu0MR/LPDr2e1jt0RNRoP793zG
JUKGwp2OX+AnUWcn0365e4sdgPftNz58dRRSkaZs0jRrQUp9IvOdhPYlPMuZfZhG8HXYLIJcBgi+
5dmhZsa/2/9t3zdAnu6cCONsO6ZZKi1lR+39PuM+L+jbPWYRG+MVsi/JQApUkT42XINGvYVCimCp
q/0m8IjLtw6S+a+wJDCT2wXgZtjDFeyW2OLlR5F11Cah8P0n+Jlji4FINT+3Mz9qs4WoH35MrTOP
OP1fncPzaAfnfSP84BVY/rIooQjJm85McBt7Krd5zFnQvZBBmvhCl/zc1JqbsEzIio/lIx4ovACI
BHO/SCeU2HYy4IpO4fuL/CGCBYahRWGDCegwXV0e1kU0OcnRKBmmAqiQEpVn5q6v3SIlviiA0Zp0
489iNBio7EdL2Lp18kmuLgi/UKVqk0Q6LIuqzbKVq4s9RM7lNfoacdi2datM4q7fZNJVV3c5Z0QX
GGCWuNGxUuSx/2NoG/R+kqlRIKgH62UB2eWBdiXXjwYllQPnK2UotND9V9stLZAHfD4Feb9BFw7Z
2tM9s8xBolHPm2G7OOwsuhWtiAgS6PZ35zH7vOdnj/b3gdPeDG4ZzwNQFw+T24Z9ySeaWYl9sSVu
UFTRUpBdEF+SXifUmMvc7Y0TeJiuBnK/Qr5Itl4DgNeaXp90lIoJOyDRXwsVFVNEYJLcqqmuS7KM
TccWO8Ehzddc7eMV77svGZmqs9hxJNsJywBAG5R5AubV6qINbURoN0MLV6UP25V+M5+CPLP9k2Bh
nxpkrXiu5s675hUJco51CL1WQAHl3pzvCzt1qAXEpy3Z7tLzyi6wdePNCtThJTUsMqwzmlVacacK
pyqondnWLXzb/tFDFmyUJAKWnzpkCbP1vhpu1JcqTJ4fUNFyID3lNk36LzjQD4u5pAs4GGu6OIRS
S+k28CTEXW9KVXiCBBJt9kbd/+tnlSLqjr0gicuMmXgpw1Ftrw0A7zr1fVGZ0mMsjEsKYiiP+h3F
yQuTq/jLxVmR6cH0ZmziBLkEZkWGWIz7+nabpcPwwx/W9FIaXN267emmx9NMM3ySOhiKhWlpQxIV
BTnODaNkG5usOxln5XOIkIumdqJjN1lh2wOA86OlaHzawgiO7mlv/9oYPMOWyooypLwLHx2a6ZFO
haf75fGB0r8dqSN2ySU2KGRScDi000aZxDEY5Bp+beGTiWo0DN/Vv4LXvHSHUMPFsM9hHpRphE3X
oomxE8dMTqmgeCSMWzlqFG9aCGUQdWGILbzHxZYmRtoUKo9WgdxmSaCM3L416Lfoo6Gm5G0y/BvC
MltUj1nBr+Mq4g4Tj9JGZ4C/LMgpjKnDbLWHfFIl6NV9jip6/bVjEOoJw5Y3zIe4L+43KwM56mdq
pemZAgaLrQtiySLPRI/RJobT1yWzLwpH0c5uIrMtsyfSYfvJibkBcYMSAKA1yI24XgEmDIM1lXVG
neKuoYGoMFcd/dvSdNH5aj44bNRnb11P59Sij1u+MnH6UFCx/7zKIanc5jlMKlz/WK2tlfEo2e4x
GcphOYh65qKkKQ7mEi3njzi/RgpcqOuQFunB2fNeq7LH6ttx+m6QoaBdoMpoZjRKQLV/eNx2cTMd
7gX8lQCm6c+fv2sGDu8bMSDf4kNf/HMoNjPGpgYJfId6ZcMMy/AUeNOw5Us7FtdASj8gXbXrLUc8
L5JDwFlUtD0a3jz6pTj5he95Zf6blj87VI4vX8bCanlO53jvrv1/XAM8Keo3fZYLA0hauyup61Yb
ui4zKt+bc+DEZECZaH8O1So872w21vqUbueATle7bht7PJ4FBZRrke9x/a6LUld8D0vnCD1g+afM
w3zgXBfe+m2CpAURUu1SSkbvgCGalEpLuix86th1qBE/Xye2bIJD4YVaUmcO9k06gDPBtWdYCP4C
Ns3QxFhMGK3xtZWkq3xT20XB34ltdk5BlzG+EAiE0DZkuBsh20o/w+5vCoCR8uVqcZ0AN1Qe+6tc
C1S1M1az6ySKBbZno7ydCVAmYD23bwsNome6hhTBoY1pg1ign7EgcWbgUStZ6urvd5sLFmknyaYw
bnq+hxOp6MHikuUT51wDrexXh6DWDSTOJ0EYBUzmgjKjrxSgmsPo2BIc9pRBVMPONtwuSh/UGxgx
O83LJaDf7tii+AT2zWSHWz2XXsUb9LXEgedGf5C2pr/CMe9C5KU0IPoOEE1wcZEGV73vEyqm0/nY
VVHj0vok/DLyV1jWrv7fBdN0D69wByaR1Mu0mXqbx+c8x69RCV/M85jEpqOoh9vnRLPA81+luVpI
6UWbTlA51cqvQxr4q7vFM2uSakqWUmfmoXRbCaFSu/KyZhIH8T6ae1sb86nn/cO4f02bBXCk+5aU
hxrtAbatBcRMTzALWOxOulnNmRHMUXiOsNKobBneKElTthdnewkP9gm2Oobn5kFJzqrxQoYX+MVF
+vMmeudLssIbbR6QpAeqlk+ZO+P8q2CcKbrB5gkdkHYUX4jh/tbPLoWR/t13wav04uYgDmQwm0NV
3V5UUwxHMQ9F+dO1REN1c28riENI0Nxuhxj0qhdhfdW+WP+SvXPfTCsGM8LjpjQnIuNVhFr0isw7
YoH7/xfqxLDuWPPtkkfzvjZ0f3zjwhKFH1ELR2NN/IcDD3u2qFq1ZnvjQUGDnjm4yHKAJTBdsOnG
H+wA/iVGSItuunjIQl2Xbw44W6fEGdkwbFhOLTyy2C8KIUzlx49409Om+t2N1OWDHvBCEao9xBKz
lBlOAnGujZ0+kUyr7YYOeco+YihruY6R4dZ1SakO7VZ7YMry5oBbGMvFMAEG8kZsCdKgHKykhv8x
NtVviMdqeSmPOwwzk7OVUPp0d95qXMklkZr0mF22hJyW5udmo/44LY7G184uxCGVQ923U951UU2j
8QalUcJkCTDJ7gZh8dj2AznWnwHstuviY9/zQuDfJgHfrqDXY/QO1Qtupr264UIoehWORuGTww2a
BwEIY1VbGyA4xbI9IZighEeJGnWpuOzNflgBsBAnNG+Na86zf60UuV/EXY76A9xn//w8eoszsxX1
/cgUdqF97oeyN72O+Hwy87uCTzYz97Uq3mToEUU68riNfyL0149hXyD0uR9jEefCMdckZMu5XqZV
04MF7esnskfR0o5i9UeM2rsvDBbNaGiqMDdJVyYPXwKeOKHjAJ7S5lhPNdDhmBICgdYlDykloMQi
KTBvvI23dB86GVGm7WxD/2m2GM6bOIeIFOSO4Rpahd635SB8J3kePUjv5Sa/AuKQozIpA/Xic3ad
3t5wSGLoXhWSeCvHx02yM9yZnXHEsJrzwADhCbWYbkC4JPVvlzX7Vyh1y0+focBJblwoj+WdQ4Tm
MxifOkLRhq80IdCfu/REhLJFu4W9fy4Ii0+TxsZl4DsoIC0KiZ7smIPqJLT12SRh0QwWnynrO94t
O4KhiesShiKOIDnhEiJXoy5bVb74Y/b+JrLGKn3mP5gTOeVc2JbkMfYk8sHIL1MRPePVh85pFINj
zAMucz/8BPGpkvtyijrER9hstB5WzhJnEogBuHJRsS/2fBkCxHTtb6wb8GCSsPXy4yE6/RzRIye+
qSZBnTMirAy++hfUycg9Sw08R0c71TPPPkKzz986rxE6YU1FYk+0h4nEGfquxrXzp9FetEwFYcZq
2p6JKWge5Uf+SPzd2b/aPX0CBIZDLBS0csCT7O0ynGZH90HFGw376zqH1DxqspXFo6rw+N3zaq2P
Z3347XDVbiABMw864cv/pQFrf4zf4RK+Ofv52JxVOAi8vZxcr0dfjgmIl82IpaRUtgzLClKXF1ME
NIN5ISLaG3Mw0q8PqCu43h6XJ4Zv6xqs9a20BZP+XCW6WLRCfVXbdaZXtoDmzKcF1nvj9eFq3p1M
X5n0Y3YYwAPWHebRVW4IrQpd2bR7+xANDvvMbLJKcyEtzKSs/qxzuB84oPf7y2WrtWlXBiCedN44
khDfuwUGH/wxSnoKbyL9auc+81gw9fNK2aq6Sq4MGrZU62j0VsJxVtGhA94+jnoz57m+ItDf0fBc
UCxZZEc/ERubIrlwXbpEDQUDVlsQyGLQsDd2hEo4DgEotH3reBe3E2NJXscRoGZgxh0XYirnkqJs
AflTkQMnMKg9nW01izKDYJwmUdoFis1KQFx744b99tIZ3lcShxWT4TH1IsufQWUkclXJ84zis5uh
NSV9zL4gHz1bz0SKrSHIjyweDphcq2yQrafdRL+Uf0gCdLJIt3s+e/2VYDHNFN05AUUNCBE7sG/h
V7CptzVeOlodpyzZ3c/KChUWLs9bV5XL+i2eT5zlK4ncxRDJtCUipeCYjuVgOPWftzo8zGtkzMoy
vNTvOyXqr7jXymmWq+pKZNyUV94R5YLZKYlEJpWtCxZyqKEHEDUSXVOvwFkle4j5VqF+JK1CQL74
tZK2+14AZtX/0aesTCnpXqWmXVg1hGKgBxCHbk0aEyoa2Rx5ZJm+fl4tQKl8tJTXpMkAj25qoSNL
9DnpbYlzH7laKWmOQiz2TybCyyS+Xt3uU0MRmV+06vSlGd5W2+c5JrJdaYIXXrUfNBdcmN/mw66L
hCsq4dsTtGUQtdwPOBITFI4y+6fNduViHpeTQUKsmFnEyRkoXn9dXIHJIyOBp+HnlUdj3UPyE2Ko
hGKfzkHb4K2SoAwH90irLUO8k4vOK/IknqXikxNW52zlU+CfgS7EjJIxPVuzVnyKUKWcmVFbFHwN
NiyzgHYRVUNNGnJSATCTACg7y1CZle39LMRKIhumCGoZDjZOajDJgni/Y6mKQlaVXT1kgNkaoeQz
sPJpM8e80lx1XhHeDMfF9LLrCvMEPsJeHp5/U5AFk2nAcv5eC8QAZoi2M4TUTvnzoe8CNzhCbucK
YKSq7EExOBYyLyhGxczVmHFZ1/EzEwxTf03nhlkvAQQ7C6omTlBVnjVVE6YK5rlzmDedm++zSsz5
CxeFKgKoAqaIpp9BRv2OiuKl2DZvx6lytkH6wybAgUL5r978xn650g17bFr/2sFwGxFtj99wdNf5
oruFKu06dDudGQRhRdYFrVS8zmeBQXOFp/KE4vIwMegyWzLZVAG+W32a3yzNOxZacoDbBpNY9EZK
wXi9xncREe1WcA55TAu2bnzS3kz6GIxg17f+mpY1OguGRRdzLAI78OzmYLKB6BmloV4RrF7+Wna5
KdkzHrlKx10pBLL1u5Db6HHlNHJ8TwvGLc0v799P0WzW3Tu0ywAouwu7ffU3cIyCvLQ9a5ujq1UB
C7dt8XwPFrKukztZ1t/nHpEmqWSMRFitmTcp3PAhsRqU+HRGP9xfA0yM1ylf46yoRvX8z1mG8lan
LpnoKHtW7KhHJM2DYWE2zooPMdquF6+tiQzC6V/f4ClAJBXfaOt8Gf6bc70/DeoKQMuNxiAK9xN5
2/dvUg5yudp+6MzpBBY2FmnR7FkMIAlhenzOAgVoKi5l3nVo+DvVxGl2X31SYUJu4qqeIRajzMvG
WkzTMGMFEB+/pTBsK6nD4lr/xO8oj3NOi4OfqQ2SgqeaSpbp6z0/bjzP198YxBEpbkp3ySYGsZCv
6NKwFqfaNHL8bfwcDa+DJ1UQkASTiEMAmBv+gtzWBseYruS05NA+ZrXk5z7C+qiR6oIQz4tKR6Jr
TKlALJv+EgvInt5GSBWeaxNtXouOzBWSV8/dhpiVu+1xTi2TgFm+NjVtB3UxQUT7oBn+Q6TFkQxj
R6xfz1XoclfTQT5S9CSCfUskvGYNTWbkngkX0oRH6wwTnvBGvfrJLNBe0zg+0g7BjaBRRfSPdo6S
ustgQhl+W3ORunyaduRjbiWtaGZq1lPnU6zGCWvjlIzjZVgqr13HEkrD9EX4tIU/mpMuEsUv/7Ft
qu1rQpnYov0hnCsbW6OefzptTwDBvhi6J61HvgPWsJT8Tt0cAGGg+8jWgMJUJY3SFTNhAKmFJjC/
Ad+tm0Ki0KIZYMxoINLdIotKh+MfxgA/wGLS8zI/48QTT+4orumhzEdUJSbwsXwcS5b4Y9rIGxSx
LwetVp/LYigt/QrYIhlyDePi4OVZzQzKJbTZ6dqX7k14j/s0GgpMOWDd1R5sP+1Mo2gFPB7d/CRN
0J9zH3OGeXIJoFLyy/K0GjnGFIYx4JUJTWP/qBDzahL5JwU7AxDddWFwT8t8ZZcyDYYeSZYdh9+G
IqXIqGM+0G6NiQJMsqWRSAQ5Ik4td83HqhtLbbgZuqwtalr/RLlfPLg9eRsxOj3Zi9A+ztZnrm3W
tYkBYbbXP3oao2kWPQwHewsPgepr0OXN/NU0k3N9ps14EmfTxQKVAB/Ye+6J6zehNhD/o+5Mf4ke
fY/a0JpTXn8F9+878HIzkVAWCJvveqTkI0o0zCO6IG0J8/sF25sOh1AfzKZzw/W32nsCqmF3/z2R
W2Knodpe9CMMOzHDpOepRKoQG48D7G6h3GdEl0Cv17sp1FceMSFjrE/HNA1ht0mZrtKAb/P7MB/n
dPyIAeoI5iJQkAt5JE/bx9YDKPmaggOvPuE/N69IR24/J1qwX/Csv+k5Q98TyN080lLvMeKozZG0
pOphhz14SAawsuRyUF5w6bHy7CyVF5ocW/7wGbE7ROUM18abYi+PbiJMJ5xXoZTZyj9mEfYK4Fyq
TabhrxOlJQZW34IrXMVP48sUHS51N2rxQ5V7LynT7VfJfo3q7gRPcwaSa3NVazZj0Ncc9yI2dtZE
o6k3Zxo8Wl5QZuIeVx9PYYZCv/u9d6d/UCNCXbpmYa+iCQj7l1RbkC7IXtI7CqWJmZ52dT1zktBI
/izYl3ixWEXmuclRmHSaI2dX6EzNAzvKi5b+Fgjgpk9y3qWp/oLYoPlnd883otb+/81uLgj/NSeb
ANQPCBQzYPz1RDq8r3YhfvW5554pr7UdkQj0oxT5jZkeAr1IivzSYW3fyUjS+cyso3fCTaTyMglX
piyVB5L6qmInxBa003gXTeDFwgKgibDVX4V/W450qlcRf2DilkcSBQW8lWN9gD2GNI5RJc90tEcH
PBmZ1Uzb9uOLJ/B8MUivneDyYlhtvlOoEGfJ3NOw4PTY3Y2eyvGhFUnZmj/sPMqV/fTv1M4lV7DR
3mjtfktEgPFraushj1H0zgoqGRH6OwFS5pHfagfkrAc4eSW3MypaiI8wdM1Sdweb7WleA9jAiiZh
kLPHTnoVi0mY+PBNrpkx2IE0wdKBOyGcC7Cv0TTYToIZ/54b+NqRrMEXy97WBRv54vCDqPZG8Ovm
FZ1NvI1S6u5Y9TnuJuyRh1+Qr2e9P8pM3L30MXSwTO6KmJQMX53QrlFZF/hs81IS9xa3S7dBuOAS
ZjFuNTgTk8BqQD8OLAlqsRvIqIJtPJB5lr0mb1aauwimvweSagxvXTg6u2+BLJwle62LAqNyOshG
z6oFFXLUATRMzlF1nWSZtGskJEPTtAvuSP5cZg8eDR9tT/xo/H2IJ/ry1v/uX67RuqS9PpMzJApl
DsN5/yGQIXX7xTYB1ZUXpNxk2OZnGRKVG0fDDtXT/O9XjwCfxqDb6onzb1XPHaMgSyGYq39VKDMi
8IodrOUu3foJJgrM52VYd2vviRVgaQPpetDVRUquEONuSNPPHzT9kAM6AEelfSp1qmPe6X+moauo
IBopqwe8ZqxslYY0mXbd5LBTPDM9oovAoeZPddZyTTcHwAanY7BjdYv1M0z02zpLmnIMN+1+1mAM
K0Jq8G9NDgbsI0Zi1eSdZqL1LJdDnmR1QsAbwkaQWQCZBcOaN1+Ogx3UoaRIatZKaSiYS5ktYU1b
JLK+XChb/g6dpAeY934TCaI/plsI04R8SmhMvptlZ6IyyoUR5D99XMu7iiL8VZ3CJw6gbTn+mRK1
d9e5mudohscJ9VDnzpUjoaqlvBzFXL994YPzFtR80ipUHsPFDAd/woYT28MSHBkIZuDm/3olg6T4
rymDBH9ruCs4lf8eSVzVGiDG4SDjzoyfLcNC+K9X7M5mWO/k6RG8fsOYj5P+faO632tzubiblZWO
tlaozAGdnM2iXhlWgf9PoXW/5Iej8GMer5EYwEHri5YJIyt6aUaLADO3RponuQZ+ki8kIEHrT0U7
SdnXfpnClwus0coy/6zuq7tEmNwoh95EU3OYgTm7TLzz5DhfcojlcAgS+wRxyNaA8Va3V/Dkqwc+
LxDwNv8l9DXUiIzTkbGCCgXScLXrJsiNGT/JDym9FHZqCP3KOa5u5IVcBze4cbBvWuP52vNW+QUI
+6zmAPJRDUsKAfM1r21JfRcnSC6tyyy6/ENg9Nr+3esfrcQYHwhrIK1EBJ+D40dsES0DHCe61nNL
sQskIbttW4277YQ7sSIL1M/ABWByV7puVLlZJa/ZvkHfh6ZoGKMttaxSd76k46alM8TPCzNvg70+
AHwJbUJuWlJKxy2kyuMI5lpT7oqRrG4Rgifrh2rKeTGkNOuP2ky9gwOWfTKLw7Y7ZzhSwf/aISDD
Rq3kOkeNKS4SHALG5D0rvtxc1Og3D5Zd9YRHooFXDPJrGKlBBhM57V4i+s8XADYWPWqH26mNIAQU
5gH9V/xMoLh6EpvXf6CT7WB2aIKn3+gbHgSRomDw/UG3I3yEeBaYzoNUw0Yx8Hgpx8c32sDsMtrC
/qTW691is35h8FOdcgV0v+725YAj97SsUbmE9urFBNcqGH1rHz3vXFbS99Rd5gjrEkCs1DlBqd7n
8QxKvnYcbZPjBrpDRpm/cAGtyWKE7fU1zGAkSNqRhKRwI1aDfVmxqk5Wgqjrq8N9bUA33Ta4iEPU
fjFtKYjnucOCkzQrVnTL0vGg3DKlPGkQeGIZl/mOEQbRgdYMzuO243bIe0Kt4lZ7iRsfVax3ZOkU
sF+tok2WKysvllo/bs9/FS22Mz0hgKnesrQ5QYWz6F0RDzhGZf18t1IO7L0k7ZUFpaiRXJvJ0wRa
7GYtiHeXApTOaMWARe6PRxKwOzb+Bc1bKEq2TEJGTgDWBOYHA/ItV76ddl3v26inaAncs+oPQcLx
DDfeBHY8LLaJoHMZcYZ0QLJix8SQtYbutzLUy6P/F0KZwA4s1RMyI8hsuPUezD0WMZwNbkOKEwH8
gzOqLLgfsYEMuxP/y7erpyx6szVJFTagt1Ywp7jtndrZXZTC0/TCVO1J6RZxiPvsKQIDQmzEbLyW
cxfebYypR3zgPxxNE7mB40dojbCxFoFtj5CH0AMSdZzAqUoQbwrkrxZ9xfe+lEmjdRfJoc8d4OcG
fOJ/i5mfRyelravBBV2CC+X30kH28LTSguI/ljjY0Q8FlGBLpuxKzFPHX3X/Gj4a/CMxZrFWWnMf
ngQfPfk/a5ToKn9Lja12r9IOLl06i77TSqjWV06TjKQfeXUttHc6rOi2wnI1zWCQOUwnJqlwUBh6
bmvu7c6oFW4VRCC1Q0zXMVAwN7CHVccDTBuqbxmtRnciEHema4JUN3LhwrTzUGGS+0OhjwZWAQxj
ncIMg1xw7S44ne060zjv1aYObs0It8QIYXsfr1kJJd4bYi5GXbwFqblRiU3dZ1HHV6fC9te1mDvY
p+dAYZbK97Kjb2I/WTG1PooXRr1x3idm/8y+rjmPOCgplEQEM8tlKxqtzX/Wc7zK2sqSKQz6AiWJ
n4/wyIPxkVjoL8qyNp3r2oCqbROMIylelxVx2w8itEGtW0auA30ObnBVxVIcG+XYHHE++K2t+puU
NjlmKCG29J+IrGWyL09yiqfuvgAd3RoUksWMDfrEJdU5RhRQkHc2RsPDcFa7OghLGXiFShBo5wg3
JCyzPABy6aaZpf9MjRLKisBv7fFgXj+e7Yms3fq2Cu/19BFRBIwxMkTTKh/EJtK5DF+gQyaMTaPi
hMgzdgH7txVKzu1oolz8chW6OzQOOD35i/p2hR4qsPUjoC5gPevYBD8JypL3jtWzCliI+S9y+41X
YaBBW/1V39fgSi4SDjb0MQUW7nRSyXypKYuTwd2EGfOn8tilhsMoQw6JHowe2vm5LDCXMSvo6hNX
qalVJQDgJZeRH44Di7Cir+5pSmITDJCMcE4yS1fi4gKMySGwYD8859ebk5LYxDwk2/msHV03+2XL
z8byEiCS1BvnegVt/rqKpo4OGtHhPm8HA35sCqQtb+sGGvr5K7d7KmnDBHKMbjrMyw9RonEkQvjW
L848Rf+eqMPmT1/SIZKrRH1ACxwBqVeE8gavKSo3O9bFp41vZH2ajp/ADP5bYFcbCmEGmKcerjUt
vajxtZrFYv/BuhlT2CnzjoYsE/eufvl3CeOyBzSypksDdtr7YeGCE48dKd5clCF+cT+OhSme02hP
F8+AX5UdkdX3YvKzay50LPbkCdh9I04WN09pQHjT6kROadYW62qXmAcsgVljuQSfVl/iiiTzVCCR
16FD8rrF670j3K7QoJ8MhGgbLl14zHiv+87nvgFHfgqt4szbcng2nByhj97K1Of3+HHpTLni87+S
Vy3eH3xVV7qMIUt2tbKbMHcxQGPO+7pQiNNNZ/IlUjun/D9Y/Wujngky/ic8kQ9GDHyIhuu4D1my
Q2lsChenlaixOwUssvAfQJBq9guYFACrodsb16cz8ho34SiYXEnS8ecA3YlhKxiq0JQI76np3aOw
cvDzdX4nVUiFVlfGC6vM2TvikOx4NfSqCUXrFcgUDoy/5+rykp1Am3F+Tpm9pQbi9e8BNcS2saIV
QTf+B5f4X1J11lyDLlr4AC0TvKwIU9AJHo5gCyHJdu6D5eia4jijO+I3+TQ/1TJO1TF4Kg7cPvUS
FnI0iXOy3JGMacN18v52+pIp44zC9O8QS/BSdvwf8Kr4H6o1RWm83TPSfSzJ2n0lHNAwtZgwup/l
qM8lCyo9MnAbK0Wyjqr8OEr91B142FobJJrpk2maA8r2qZckr8M3xeCXztdXE7n6t/6xbdApOQnk
ZqpNjJPGUthlGUfy9ITBc8HNglbCL5pAGM19D96C+ZFwI0OgIR2PCbaouru9EphaxTyLPhg9RHTB
ZqyXvEPoCE8aUmjKvD3NT2hHaDvbNdH/1n7vq3gI8Dkxts+PpzwUcJlBnhQV5DwZxv4CfF2XPWDG
qOoDP5ENBktfADOM+fnuCeR07Mzd0ZWkBWlGCku+hJ9fRbYLWmTugYqcy+pWoLYGYEJNB+20D044
KucC5BO+TwzVXt0PUY/uiqHPT2iLC4Mv9yx8IDecnW0/NKFxJm0A5SoFkfXiuYJG9liWxOMEolHW
GBK4Kgd4LKnN2kcPClWOiHtUCt7jB4EWlRIkkJl89OV61kJbdsrr0qv8rdT8N/lF/747DiDZK9Mf
qCzty2XlOcjEvTJoAhcnFRykN2PL40ozhHksNUvi+XZicrqoQermu67MyOHd5wLL5XNX36p/RNR9
oZqFm0QHRlGKX84ZODcnNJFNIV7oZUYCDBVGhwxT/GdUfyzi6sxHx+pKQ+v1nHlW4ik72FYYXW28
mOseRcMAtACwdaGxQ+Z/ERHKUMDHqHbmkQkG/+dDLIsiuSwT+9luuys1aGvTWKH9tZ9m5be4neIM
dgNI9dWEs6s8UUvJpNPUwB2j2KoLtKPn60h52uxm39XqTgxONrTO99y87cKVVLvWOCHb/pLDD1J4
aDUJ1thwiIUgP3xNaXfNN3s6AsK1ke6gwBmaKFc7QJQHeVd/g+yTucFMm5nv2qmYgi1aACBvK4Zx
tEDp+ZVNL/G5GdC571uNruGaYFLrioCkB38jpuEAQPi9iIPJ9AB9hbzoqZG9dy5hNVXBf+O25gjx
MYdM0otHB3lns4YR43JMuXRx4rFn3hrZpiyiCFHgay2qlmi7t0TyenMY9WxSOL+tG4UZLPQTu+AG
ltlvR6SoIrRdbyYns3IihBGtMAuZlBzLC8BbwT7Qq3G8M+pZ0gLiHneDjuNT1lYtJupRVjzzFw8C
NqvFClcEY8Ft22sZm8I5NpkWOKcnWI2GIhUQX+lOM2CWCkcJQgTvmXHOCxyB7eDH5hf0tJUsnK1r
ZfejtcHpJNUmKTAiBNVWSylJWk3EzXzDPypSqFwNDCSdQ4Gwhv4pY6Li4Gx4v2CDukTUCF7tDabr
E/XKV1uNYOUsYPKH+AGmtJNZPYBYHfrdVFEYpItJ7aH9xx1WThTTUphMDn7gBf+UY7jDnqJiU31G
iMjLOoD1KBf3OxtYlk/q3+hDOEGbi9rS8qa6GQpRW3LR6Gl24RVMSbPAHgJK2jf3n2qygzZgBL+P
gu3siTB7s8SuegrIeLB1dLN5gMlABw+oXOL+ZaRIF1c/WaIT5sLjVmU4Xq1on0lhfNwjoqzwi/Q5
+zgDwJAptRsOJnYYnhf+RxrYZdhbrS4Gm/p7FJYNAwhjdHP+qeaG/CuDM94KC8abng4zLpx7eYTA
mxtMjVeD+vzxDSkZ+PEcfl7Yh4C9VpfkEna0zt8Bbxis6cmAEGAcfDCmkNlnteKrVv82mgnklCz1
s7lTOV/vnCPVC+B88ISAbiSENEFpfAgFkBCO+Q0VAo+/dpbOUVNBIa206Ou2fzlLGyloC4NA8tgh
kffP+ZTTJxwZrECvmCO3Fv6iK2Yk1hw0twZScnzZSQE2/LsHQXnTjCvb/vxpzWQTSfPeq7iCzKji
PVN/lkARklklwyV1szPQIyPygVbrNucoK8jw0esgCNdsoTGmntlC47LEPvhmiVmvj2cdwez682ZO
YFs9n6RFmaNp47JY695zuBD4MA/jc2Wo8QIgR9ydyum+NZ5nouj3fFCGaUf3ou8MDLmn/4C8E89E
t7S/Whom88I3mq8hfemz9HwOTnQpEa7pyDj+RaCaa1KathDAOyOpRi4Xt6AdnT1Qx4bCmThmJVKe
03uGJOuqyJgZXy22fcln4BkaqPWzJG60IEUb5iRnIRTGoWy6plQZsHv6v5z9F1uEtrMrTYo8s9Pm
phR+bD7mY7/QFlI0JPa1CwEtKuGaZwuPA3xkTRgiSF8Pjg/76kq/an3r74jea9DrXWGNCYxm2yEG
raMWSY/RqkSAuGc4z4coqJzlMA4qsQF9qpn6vOEJ3y0XHYSkhs2reDB44EOqhCbH1Hj5eOUm0XkV
ABfG0FIXYBNDD2nm7TQ5uO6u1U49hbKEvBOy7PaUsIciUz6pvgKhQ621eY9a1t+sAU7Jtb/rDsrW
PlY1X7YsYNXyugNICSufNSpdDD1nNUWxR1EMyRkLJW4ghUUUCnzmAD2ce7L+k4aWTtbuwNmUepsS
pd2/SqSOyMyCXvW8FlYHz5jnO7vakkxCwWS4+s9TMRefoKOl2XRhsPnb7MbXDADnX8MgltgL/v+8
PuZc2E7X2NfELPBxwnn9Lc1NQnHLnZp+AbOo2zD+ad3LjcWv3OY5F6NUMUIQ7YMtPmI5EKZzsDHh
RgZIGyBs7EvNaVTJjrpHQUAwOETzBF2O1Xx5YIxmYpb2qn9fp/L3I5hKp/2T3CttAvpwuZfn17Av
iJcASvNQKVbiMlak0EH+8VSAEM2zWAHao5TWHnbGvTpqtr9FiseoXgoH3WjclDtY+6M/tUrtua8o
kL6ph7eMgGZjQGI4iQ91oe+/bohU9m6z6fgK/6Ry0G0A82QlxRKit2F6hDBDzXqoUsD3WMKtSJLj
FXXTObxYEBvi3cCTolFl3eXSjz0Jxo2nOtwsIn0Ci4YmwhuvQiK921dSUYu1YI5ncxSPhGnoWbJp
wtson2fGfBXLTytE9mCHrqE0rLbvV9jgIFcDYG09N4qHqDKoztpX7K47xtEPCyUjh92crt8I7xXK
JKz/QA/7/JWpxK6T878oT9b+mZc7nB+m8ejIiCcIfVbBUg1NGAsge0lOyHFLEBFgUoMWzAIeuAiJ
DIww/76rao7GFdau2xevNQt+ljLR1FvMYicVFFFM/0ly0Qy4wIYJeGsonm9oee8ZZORnVj6GssR8
GFlAkOA69gIqkUNIY5v4FrCPyyVFyvsKtEB2+wt5vLq7lsIZ/Vn072uoRW6A26rytwRp6K8XAZ9q
XqFKsvm5F4Fv3SftdH6Y+CWkfQBfyiBFgxEs1boeqesv0asfwJwAW2u521t2iJ0EFMMRtFk5ZOG9
yp2RjDpWlj2qlyXqRrCUe9lEDQafCAw5YPnTAMbOBO/Np7728yTPpV9F+KZ9473J9j+SUxwMnGrK
GMu/YFaFh5cFbV+lQwD6i2jWIj5J8ax6S7bieIfPFcDEqQEZT7hR1gSBpIkQOrgPTlOKk0wYrBUf
o+U8ZcIaMvQo5Ux/CBBmZ6wWcoGvnvFsPolCXcXjFFsUsysyVTT5Islz2ss2vo+cdtKZwzT2uflK
zwVdLT+j8Bhv2P+kNYqayw7YXlwy6rQsP9U8gbucU63YAhFyZMMP3DlgumSBxvY1fTBguO6IzTm4
pcZSheVDDoeHx4BZ8nw45MGMTlSYu8rG+p7ne5YzI70cXrsZ8VEprBcSVfE5GziVoRkz3MLX90Fk
RXyFP61wOsVlZJg3Y9Fcc6eNzbWa51x1KFyVInH9bvByDtHC7d1+dGcemwv+osEKIUuLXiR6RMWl
NHQofywU4thjJboW+NMBKWgD/1ajzrTZYyb2Qygv/rkxS3h4FXHlm92Me10h3W4RMPsZmeBxG7mc
yVUlKFbCVnsctp+uEAOD+OzVj2aTMBNXSgOwYgFMw3mpbL+qPLIRiinPU9ZGNRWOkShGU4NrE/G0
5SWScdyOLJXyJehYnVu46hkVJFrAo5ABkmzVMW4zd9XzrFS3g8o9VkeRapXSNGR3KvuWKPKYhNZk
BfZuOu86gSst474h6mLM5uLklYfO8gBHES81M03QhthBT5BxyUGuM7h3hFtTC0aB4cwXIecoYNXq
zsJGOkCYJU5+E1/TCtk4UhMlxeCJixJkHAAjLH88qp1VGZ1P6fI+uPiuH0W+Xhg5iKspTKYdaslh
dwd3GPyIsIbqA0Im6z43Oc+Bqos7DTl5xSzIoh0NJdRVPD3oLAUjBKG1a39JRpHs2i3I535LPClL
7OqUpWa5u1Iqut6yvMEO0b8Pis/pF1ysa/003qTesgmdXIeAWQGm0JzLnW7vZZ+GwIn6IgKr1NbH
HqXk1c4bgk/afk+HDsvcbOb2Jo70NqmagDvEHA6NQx6SPTQ4ysta+0jGnkXyyevFumtb6o2Y0EzW
vrKS3JwKzMOydgG7qMFpMf7lsBGSiAY6S2zKXZvkh29yOiJDP4Z7UgcB1KVre7u5EVwTTSUIMc+N
vl7HyHW49ITJoeVk+f/QXxxqlmbUjpsLILzn6OShLlCbQTlRig87BepVgYiYiGKgznU40VrgfK9U
0nWDtv/0Cj/jaakXjYj79iKwo1XV77z9ey+KT/YITfzGsn+h3C4gj5vTroPT67ygNsP0XGNDqEjl
XfI+coAUXErwt+NqPhSxMabC7Etm2FlMTsSnQYJarjCWCVfvJrTW7SYRMn4Z12ZqVP2FDV1kTkFO
ApyKoLfvfr8KBNHAqyFkmUjAz3JkIAq0z9tKVJYeY9KhI6/+JJv1mdUIyDzh+DlAQX3vzsfTsv7d
V6Qz7tcpSqKWY7wF0IRyw2KTcxQbaDxQU3b2oQU9EDgoz/KoQBh65anvEvyauCuvV/QqxuLXgz/A
mhwB7TI62akJtJaIevvdzF1QCOg84fAuVvvBSnJsb5EdcAVmyqEVF5V9OvqPNYrUhkJWyhYH7hOj
BcJDxe4vQfFZROoF9ppxjTBkLb4umo9yT4enurxTgfIT9l1kBOFHlUW0XA2/TnF47nI9GiRpuMxy
QDTHMbLgNvj/T0bQAoKVIBnTCncR07F4NFFhhC/GRSBYK+R7BRVa+/TN5GIPsApX5kJfw4KQG3qU
d7qe+dNnGNfpa97QccLPpV9GLvSdTsi60rAHMPm6ZyTbeRCDZBkvvQXjzwrk3F0J170jpxBmSSqh
7EZvvzuiBTaXACyGgv1hEsQzbzGT6vmkDQVZMNhQWdeioiB6EvnFoGWlRsAwJxNcAa+FMaACr5EB
GycmcXqU8Rh7gUCiNcL8DBuh+706keqzxDY8mOU9793YkAbwFo9BoSSL6qTBRlJjU4fmn1WrL2sd
rYA5C6WHls5bhVruUhlS3hNNfKhNhp2tznzSlxIwTsFyW2vkJZk6L/zwkD8zDi4O4KB3JCyJzFhX
mz2VUVA01zOWqVgWxgc9f+ZWewN6eLPWj7R5NY1KxeyrPF5ZstmMgqD7D2EOgBMhIZFwZ6oVh8AC
6JaXXR4eatzBazzMXWzEIxzut530BRCm0Q+A9RyuahJo0qfMoNYVq6tBx19U9+QHK10a9qDcFRR5
XjN1NgmikNymDGeveyS9RYc6HPWGEzTEfaE9oI8dbdrijY/wWOrcbLdHni6JuZuadZ/4+D6PYbsF
si0yozlpdVEEE7U8HMDThVmqEWMAOQQpjTX/dHgFu7ZA2uuqkolBsXQdWTEZmo5HWo0LOc62aSFC
UhMybZtBSaTDjdSkV9e4jpX35okcjmP83ajhwMaG7GQ9Xu4p9Y0hTRYL+wU8WKg+HiOnoTrirtw5
YNI80HM/mShm9g77aOyngZAkQbGJIbCaHkyq9xJdjfz3ai80BZOHi8z6rzGPJgxTpOQ8L9bsECYl
0al2cYM+iBq8g9004WO7P7J6S6Q5sLh9hX2Dmd5lIjsTnhfPWcmzwh4jyhMydMo5XMpA42GEXW7O
Q+tGfWwH8srK5u82Bg1o/dzpw6My1J07OOmfHm7PVdSX2dYYBbOwDrZHgE9JhaNupQPVcG+ekB5a
ISMS48cqv5AoYjQklWSsJi+CAH44V3VqAkFwqqpvLHbFaf4he5ptg+VlDWK7+ql22QzKO+nu5ECw
RDOue9dN5u4fWyNY+lJKcZilySjEXZ85KDXUPHaYT7VQL9AXnE+Qn24WLTWz/OWVznSh/rghllJQ
qK52Pxal820Cj3OGkfoaVO1vfX7cBZM36KT2PXZfSWqs8hht17+/TZN0Kcv9XKq6qBEHLaNPNwIg
v3pl7OhFvtOKM7HL5RbOh64nhqTlGRfw+WA1D0FuFobxcYkEpqpteb9lm254sO9qNJzyR+LU2WlM
LrOfr6deR3+80VaPJrnvmVytXggrZBvL/i8+aSawUKPjOaNYoLh2ogy9zWYbFZ3I9oF2H5Scf/qq
GZZQ80W3uXw6nEEjJgCe5DmSJwPVCVD+aIa+GUPrHxZ7G2P2loz106sDcGNYf0ty8kfNs6cn6FMX
9MkhebbuWIG0DyDqvv8WC5fohqGhOYqd9mRAGyCuDlgcdLpByv0mJ2dcN2nMfH99OVUe7Y0U9Mn1
z/AqZ1aTB6L9trawykqfaU+T16t4GWfSj+UYYodIxWICUMmS0SLbnOg507/DKwkvcX1ZhgSGA6T+
eo/lR4xxit3wQ+KRYrH3y04STLNVUMRIo8Yvy2ri1BRq9B8rYAF8Eaa+R8cKfXlHhVlikKDKJBnA
InwKOQMKmat0iimr94ZO97hQJZgYwn6C9c+wwBXYH5nQqcCSkMUVI8urytdOBC0gt0Cz1VJuvgSa
YBlxW7fp/10iNeWZHySPG84q7a7zgwJo0Uj5n7G1OXa/t4T3VJ3kLOqDdxIMXb5ekb1aaE1U+A58
Vg1GA7NN/ZOy+tA3tBomB+/XBD2CpQZxXRbRSpJJQOkREkOD8+cQ35+wnguNI1yC6R0jvlJHhG9c
4xQ9GQGiIzaXmIo6GJ1xk2rt+flyQlZAXxT7MGISAKIKQ8rOUERD1wq8Q29MlOiAFRMHbOTndfjG
ViXcTleKb7jbj8ip8KpQN1a0CesNzK4m/EvEdXn3STN0YgsiB++aZz1A31DhJidhnbh3sgzUqr56
0K5eeHzc9lBpyFon85/n6c4V1BiJkd28TAAGXYNJYYjibw50+FgfjJaI22isA7naKmoLg4TeqC9f
cAhNeyPCFf5ZBx9ezZhcpohYZAJ4kJDE43wh5yMBIBmBQq8OoC2S3CKR4nNo++IG3wBicIZO5h1F
HWAlse01jpg0vdnvyXtkhAxKJYQ7FuLVt99UemCc5AJVcVJRjpy+7GWq9ZfvtxuBX2ZM0TMwH+F3
daiV0LwVWf/LPpR9Bb9QQpFstmKQ54IXok+wpXLyMW5GFdQjw6mkOIMo2chegq85PfIrO/plCxxs
Ej/empigRK7CGsyi+4jqp64L1jGGpPEOzdUE6zQ5Mm2UaWxqLesQykJ38T6QEgfkZlaLntfr932l
F61PuzaZK0o/Ok0f9hNM8BFYFCvA5mr8FnCQh30gOdb8MyKA/GOtxIzdHrjDGfAxIRhkj7pX+Uu3
V0NQjZpnhLB1pXdK9W9nkXPyT4ti8HCRJUdZ4KYleMlDWujIJ3EUPfTD0mSzPKkKFBAWLo8RahxM
QeGpYLGeR3R6Q+F4E9LVtyZ/+6dOQgyJq5xl3IDsW677Y3JI7f3fqkTLd0rF57GxR1WnE0C/um+4
KDx+apPxWXElr+S6XYgHpXo21uXD3q8+QtoONhIQ+8WJ7dSXpEmaB80iu/iyxhfNyr7WwwVp9R3z
UJzY1YPJ0dsdPxK0OwaMmwb70aIJsdBixp0bjCL/vbFQhvfnA9a889teavlf7m8N7zki3K82XwaF
J6OARe8HHLbHSO4Xkz+2yh9IHSw6o5RHGYyWZ11kkvZb+rRt8UxkIz4immqxyFl9qsEBdBLUqiGx
Nd4M+R6NgtRnYuwLfT5HoHhrKLPiN1qQU5RO2iIwxQMtqXU+fQ3kgRE7K6QkxXegGjE2zk7bmeLs
7J6XhG0TMzmwYJ+irP3RLUOD7dpew9jh53LpHjvvAj8tDzlE/QnFhPT+2NxYQWGstTwsq9oJ1KIf
gB6yakCn88uKbp20GwoVtRzk8v8/XJmiZixVLrWskKSLqiyodxdhUDwEr+92cnq8onl7HHfkHt2G
gFSDdKnQSacswCzXp20M8HWrfTys+xwTmqIuwcsObRGfkBZSL88l12+pdcjD8pGFLZLDPKzq6koX
Mse8nqQf14u6oz/QidXL8B2TivRQR5V1KyxlG312f4R6hSFBHY36psRYUW+WhSSp36dOaKwRVuL4
iojW0An4kusrin9vR30D7uV4W4l1aKtOZKNaT4mgAfmYWErMhGMywjfWoQQ0+UKxIdvnKJBq0O1g
xYTSPq2S6DGv1JVYb4sXjQd/9nWRJP1eyviS+eJ0BPol4+ToTw++5Yz6S07RikmtS4nJ0Vm9H3aK
CPlP2KHo840s7NCrxKvY2RxfUX6MVL/OZGUw0wzdPeQNZLxGFmz0FvLkb0FQsCvqrurnSZt0kcCP
EPQzKzSFB4OfuyijVenM+FyfnY6p3MTYas+NRuT0sLy6u5M6xIwjjkI5LgErr47/CKccTkmjt+0Z
IVg1OTcpyTqcMII2aDp1Lxmbgb5ttUTTemhZ9l6NpL5vYXm7QVBlslhniM5Jrt7Y17G7R9GCBYXg
cTlI+hICPj9ETJGJopxIrB+ReRQSk67deLn5t4eNyS4r5qb830WAdjTLbpCbj90pLYw5bXYoesTt
w41owioZZeThXdlGUg/wK30+9SLVs1WDKL1+xOikw6f/FVseAluk5KOTg56vD7uS25RNYZCca4HO
BYXD3XZ81UBNLVJNREH8TOPQBGdq88LJ8Rp8oPmNPSojvTIab0rpLjsmHUzE5J+/VoKdMknPW48a
aeU0kiMlJa8hc9lf6mwpDdgPAmBQUnXJcpO+DFRjLeTsZLkye2REDwefbRfEq+nZtb+ufF+QQDXJ
YHM4fHL2iOa0fGqRX/u3zPkKmo9jSAnIQpdLqh+BgB+f4dn7/PDl477UKhiPms1yTLq7gMyIydoe
qkiKAO6pakmXetPKzxSRaUzY8nsu3T5hzji5Y3kYKrI/W+Gb/b9dJr3M0ooEcy+7BbPiQ01zlDbO
eFPw704iGBGYJeGoGTx2JO4sLW5ZpzsVbMKsD4p0JfmJo5GDz0D7a5N7r6/LVnIMSXEisCB1S4ET
UM57DYuo3PEiYAELTnsEHCfoRFUkfwNQxu3Dza699nNzeIXZty8SZU4mMR1aE4iwxGHz1TQ5u/QR
JMQ/EcuijF8il0l5tau3oE9cOnl736yv6WNLGfHUGTSVGUCCe4VPpXsXSeModgiONx7nfxAyyEmD
K1zJz14getHQkKcbimjPJN/Z96y5gF6gZCiUyFAUYm2CL99HhtPy8yEQd++LwUJVm3tNFiDuHM/I
vdBy5/2lfzwE6uRVx7zdc93kfsEnC+StmpLs5H96EEDknb1a0J8yiALWOXuV4fhu95xY/+ezCcEy
Cfo4QkWdHXBNVqcZkCCmOFlAeWQqfNuXez/L+dFnAs2p1Ps6T97BSfD4qgFm6whettV/po0jR+N0
qOEyBFA65uFTDitui0ygqtJHRhahWgFPKLQWVocq+498gfMjksuXyyQC2rVkMnevLyyI4AtKSGVI
6ziadcDADiEzwAopTeJYbRrHQAab3PrweEB/ExVmJE67DtruvBgil35suwMo2n7eKW/T8Az9NfUb
BQOPhsAljohkVUztXbX3kvT0V0zk4SwE327GRmAm0kcDl8H7CH2ttmyzKG8R+hE09i42dDmepSyH
RhIfmXVQkmyG749UEHN+19cKFMa8EiWNuRC+c+zvJs6WWWkEBGJV+rNZ/OqyqNreR03XtLg83HJs
oysiSZqjmaYRk1Xe/B6sKy7Mpi8hX1QcG3onRCpCARbEjwuzb0NjQ3TIXHu7xPso7eTpbMm8Ms5y
HQbhQI91RTFv2bNR3hGt2nmecBDtkU1xzYW/o5cHdlBI4m/J499z67q1HG7sycyACZ8d6aMoGLps
f1a683fFqKQU5dnxvE8HciT+0nS2Qeek2iL/wy9AaO8GZhSibNZDnAaIgHiSUUfsUgRdD66Sh//Q
bLnHZAoBmNxJXMnTZZX8a1JuVFmlYbxIuLLWaal7fnmBygKKBr9blWMYo/NlgsevCHrDfCc1kQIr
d4NKrqyKd0l8en3kl0tJG2GlS/1fdSkPJB5zCIDAG12K4HskzuMJJ8wv1QLH711kLXdFym0qHgEP
YJIJl64Zo7KINljr8tMWp1lZKa45MqbUjT1e83WpdpfdLpstDitDJehvAYDfyu6SvunR6co4aCQJ
XkUgNTxck+z+5elpSwP9Z4y+zcJPQS7eS5pBUJypRVZevcV0RqsGlZWX+i/jUNH7gyj+xsw+YApw
s9mjDiQej25mu/IUMBwegO8geg9NF9CxeBP2RbGsF426GXKtXaEwDOhbr577M74zak87Lz9avTc5
go9spG9TEbPm44HTz5I4FwjoRCwaZM4h0QVPbJL5YqQUUGS+ssxsaTC8l7XHy1SdBffOU55YD+9q
PwsI73XA1NF540E/dE7Byk+OZbKmfKlTRMmK+2yKcc3DK1G/UEXqufCLpzaXFP1+Dh4wMLnQfwwR
YwKFLLaVVWNVQNb+y8GYvIqdGcJwwBjk1kqpHpPE1Wsp5lPzUcBpSyXr5dEDKOuzo3t4J3h1HMXV
eVaUQR22OLFGi+sjVl9OFk8V17QM9ga8uide6aDBXaRM9oJiC5yV3IsBRwc4ck9ipMGEMps1eFdI
kOu3YrLZ447jizoxZp9bi1eCXwCVXp6edL22IU0dg8ZOgirtGgLwrO40BHPilHR/xEgLtTKjwUvn
GqLQR8FtQhQAsOqj9knefdZ00lEe35JxjloV/Ofe208l6P4sNtUVjl8yluhpQrI6pTdBuZXF5ZxX
088pfw3tbEPheFFj5HZOnTfHAZ5G6wLtVdeWj/ET2KUqBqmXB/slTj0nqKnRX6CGBuAGmGGSUsHu
lqVVmF8u792u4XY10W5pZOe0zwMk4Ah8mJ2jBG/cbBqUkVdLcmYqd5qblncqUdalzxxrLL5k51Jy
+NDP+o8hEkI+8q8mv7WFfeSKBotLxUmph6Kal64BLcpxsoe895McODtXJeu+NabJ9zsATvUNsocT
3xIVlJ5LR1DvDYh7NAaHtjxXI9rp5GkV0n3xqKhB6/ApwJC7FdtzXmIorsSp9taVQys0Wb5yQL1E
TJUOj8pC29X3B1+UzWCsqpX8nywDC/6OH3QQqrEvr+Ff7dBG+t73ie3LCtlbQ1s+4PKr2ob++AYu
rQ9hoHU7wSUtkjlfiQehvYfIAPZ2R32SX0681Veg+8tZgnAkIsNdbOymGm0joDdaPe9MEtjO+fS1
cRaX+nmJq2kCfT7JwQsueI3HdgV52Fh+q4pBRjhvnfa3eeC7Y4b/XApsoL4d93z/iVSp61xi/55W
nKhVfDUvQTqa2Dyu3xkgzDX3k3vlPMDgfpq5qF/wFO7ldm8qC0sbCCK6qLsZOJGrYkXKD8sY9ZhN
QnYnLN9DCzKe6lejmU6WHB/YC4WgGq7KjHeBZ4k3tybcbs+tJD321BCL/wnhhH3SnbSyymIRVrFB
22Gx/YBJhJDTNEQXTepBhzPYSTWUH7Zam1sxlLjiXgWDl2eFEs526bpiaH67ZyN47IJLZ9Zjvcm6
1nxSxJcZGkvIUqixoCW1+lxXDxo7C0JUDGip6CaYi097PU7xuUth0l+qZaM/uxnMcd8dPGFw+rQt
YvZj9A3ovjcsOiSYZCjEOoUj79Wh593Rc8Uw69cQJIu435oEJ0+35Vk9vYoEJkTWUW3RCWuJYbeI
ZpvSc52xunHgvVCxqOoL+19ocVZ/fyjkkOVapZPD96v998IClXfVjhrfeoSK5zNWxgJ3p7J3yC27
8o0JFv7ArGn1vAOCHXmKulQciMfZ0ueG+md2obiUH5ZDminXrvq2gDjrwUaOOoA+0MfrhTlEtMwc
jMrwR1qloR5kdGPvoSu0Kbg6LzIMv/NSU9AfDRgYIL3jOwSfyrqanuMr3+rHogO0hqY1iAJKPNFg
/mqkAqyXzcfJr0HUQOA1FdwKzzwthuQnmXWsRJBYTh6/DSERthpWN7XW4cnp7Vm7D/k40QWVCDmq
U3xAmk4ZOgYMdkhQEQ0tl7Wt5wvyv/+kwX0B/XQ5F90gBcnbCWl6yPbGYyipq27xHuTbhXrrG2eF
QhvVmVVPTa9vUlFuprco14JWAN10L+PUVW/hUiZABWfAtPVjN/FREA7zbmvVDfjFuJZ/UOJ9YbzY
VFPJin5XbJa2AFdAU4JBGuZ8sKgJg4ssjUkjDASixTBdQmZmiAkeoZ2Xmvc4erhzwwMoeZmBjgxb
Ue90LtVfl4vW4H1yVkttJtP3Z66YWsHs2F5IBCVYgnJbvPI05uWZrmdViTOj3RjseyBzpnvAEKTK
5l6b9ckFaWocHUw5EM2pYGa39ZLuhlUklwwNP1JgeCL1oBFqUctyaQZOrJF6eY7T/FH2BZFiq6P9
vMk875tuKUm3GKOT1oTYIL9IBqd9cfuwLECcS0utjUP9wee4eCv2MzcG6zH172drlPq9VkUCXmsG
MHY+rdHJSrOmGjMD/B3B+Lah/Uu/axRJJ921h1pRnyarJRwWePAA3CoKoC9NxoXn1tnKBmgPjhv2
gEYt6aJn/MOry3/TP4lnNCMeef0euKWiPPj1yCv1xRQyf1EuCuS1P4jIzu1JoJbTpBTkKzAB2+Bu
jxcOgr5rkQUJNzn8cVGeoQYjdWlfLIrggZEFo5oEHuBO/L+acnNPRC9odPzXnpNgPXgy74g5Mbcr
6eLzXNJhFL4x0z8vpp+kazePbWx1+Oe9Xb/NjO6dDA0lWaKVcaYRcXf5aCwzRPJLbW783xHMfJjq
+t/rImKpPo0h7lhegKc7D+l0m5Nw4F94IFZElWBDaerfsiCeFas5UXGIEU3KZWkMz19znHBmYDiH
TPwGIXD8e6Fd0HC75mmLTK5NnV5EHKXw3Wbxy5ocK5kbMSqsa7DkyJZX/AqeS1XwAjuZ0pmOESRT
UdFbfFSDnhKut6xH5jzR9V3oPQBhJw8gp1E3zlORPrAbOoE3SVHLFpRKd/LFLewKAL9PYJWGgWIB
qi1vnCtUbguXpMODrUS7BNCdIfYwl1v0uTC+fvNhEorzdP17TcZpj4DBhcQ+LF3MOURTvUFqQQnE
TGdaysMApMcIeeNlpZUg5PABGsMJ/Vzm0EyIqmlrU99C3spSsqYBvvOiIqmmyc8c5WGaQPy9E6ro
TCGYYtpdkGT5zC87oMK8QWEin0w50iWkbKxEwK5CSEbDIBZCmtm3bk9gbFLLxWSPMpY2lDS5N2+b
znRFx5IpbCqLXYKXmMWmGOw2tgbqng/kwPb8NFOyq8pSCD7JnTxBKpspuOxXOsBap8gS6YPhX89p
GQ1ELxunm58ZmTnvPTQAnQkNLF/iFvoOI/Nr4yomph1o7ClC/7NAQN4PlMt8XRz6BdseTQ6HbcME
RRt+9HJTRMHMOg6uGj4rLFABtwit2tBUuf6Be4BSBwGkTtts3t8bQBQVeAeteonCvA6iu5RcVRe+
a2a8iyF9F1TYeiVRftKArPtvKdWx5bej5NrZhaWob72iEBOt0Hs5VcUQ5VXjJE5U+XGHQWvtttwg
16GePnpTCNQbbO/O56iPEb2ueP94II5smg0wduK8uEzrwPmoEoJTIJUpRGUe8xy78VRR51JN3pNM
dvYxPnhDeeowWDSsGkFGk52/eqzjvvB0iEbZ/djq8zKfAv2N43xFOjsx5+nExIwAD4TYBdi0OWk/
PgxkFP6wK8hIAB+Y6wQpryTv6DK+7ro36LnysY85d37EYOh0igRbRLXU4IU5k6qj6MlFO1yPmAs4
5kply0SUbZkxRsmujCpLV9EWowuanwKuLPvgsa+3yf0YMKEvHfI0GFaFRmqbHmGtPbdtuDly+gDN
GroauY8YoviECD2yfKt6oy4L7BepWmX5GRDaw2+EVZ20K2xEh4lvJTFdMhqg4a4y3nUGtFsdcW+X
aTu1TIE6iqeetkyUWlZSVDrmQ0zH3OzZ/Dc4mVSYdMFuMQM6Bd+laC8XZhPTPuffcR/KLS5br9+o
VGjHqnqLz0B5RoInrjLkYjfzQ0TxBLLCBCg8nAAxgXIkQQF1WiNDzKknWlDZp/wzXKJ80pp4PiZx
LZvNX3hZhzTV8ygzFHURDYfUYesPxbEDzQQJfMvgBGm9X+V/VdRNLF8qV5QzWLHS6VTdmpUnLyvA
spdrZudBXrVgoBOsDRnEC60we1v9EDwIsyUx8rMfZLqn7mE3ngVPUrYCGWiC6TmJ2zi9Cga9aTc5
QaMLCfmbs6yhOVM29hk1Q66PsWLkdhWmBlbPHBnUQa9SqPqrxJ3lsImf1RhCU1PVktmGCjeyj+h0
3phcrEhAdU4TJx1Io9ZB8rO1x93lQeyStXFvaNz/EzDuVEhlv0wy2fB2x5ngIqYhp+BG9wY6UMCl
+71y9Fj+XQZ22w5/sNZiTLklV8xDakloApEGDD/KrL0VzRuPxRnzY0Xo5NzyuxsPhG/+hOpLqYM4
CeFs5wcJjQlVSeog6DRk4QzdvMyeOFjkhKuNSUfIGgK/MayKCLqi/G6goPE7rupdY/jasjL5xprZ
gwbymJxXx7Dr2z41z8vacNW4lso51rCOA+CihrzHNWwCCUW3vWHh8b4Tt0asjYsZiFBube8dhN+Z
883+6wL8nw3lJtEDrq5mWB0NEguoonYw8VPgiQZean3bvf5AlpZK0qs3xIzhdLs4PAWXnZ31hFAI
uEldMzeweSvDuZU6bcJiwNBCP88BqF9lrCATNpI5W8eVhiSv+OonqwtijrIV8G0zYbxixsvKiowC
Nm1c5mnrChlBeCptIva80s7LZ6g2jl3mTLy1sKBpGLQbS4SAycxUG+CZaQpTbizMoKfSe/5gqOSE
erkcIX26K7wZH/wsZmYQ5hfsZnQZ4/psVRIve8tIHv/c76L9Ih5INvs3Gw2n6VGj1ISBelmaTlaF
/0lVVfIvFbIfAcxz1NYWYqaI27SXIHYqQFOtZ2el+foKW7uniHz6HIf0g40tgb+Iqr+NiovpGtob
rJxI7h3WppKe2QuqRFi4uI61jAiiS06doDRZSIVtk7+dJsj0X7sHZKfLmbLR7kzVgLq85lLFCJXy
pKw09mMs8zqsc7NI2JS8r07ZE4Zbza/MGnawpUnF2ci/Hmk5ex137LJ2BKzVtRaps+4aQr6P4K+C
dY7wmb6QVOZ0XUXzv5OnlBTYSq8FZ7QPCwyIowgCCgqisCIPfbq+F9Mf/Kxre8LdKNGgJ6VCF5pT
fvWZfxPQHT0lH/2N9SVJhm20pEEcgLDtnFikidf5wwWR8I+/mmsZr+ARp7oqSJuC6rjLH4jV3R6o
X941xMAe8V0Q9PSNNBDKiRqM40GwCdYY+c8O0dnU4Mn6KR9x3Gh0a5992awJxXTS1N1LzTkrTS19
l1qXCzEmvkMoupjPWwfOZRTW+alVRSsjjN6wDTAuJl8CJZs2AcaouuIw71y5vVvdGkIkEEUbAoeY
tCVBZtaSZzoZswzdTC0WaRlTSaNvh8Bvq2W6V3K9M3jctY7zBxRcOOUwhzOVfGXW2Iix8VDubPBR
wBYC7T8WRfTy2zJQinoqHJPYGMz/kMPkxdMjWWPSzLzYi98afJv7uGgG9fLnYJXK/0dyiuWpumvF
uv0O4b2H6gaYqOHHJy9d/BlG4/DI5JYl3HGHUgSzMYetpfK9p+vtqyG9pm0mwQcqYjV93+vY+kPG
lOeXpqdgjPotyr0n2x3EpwRcYPZX+O3nhYxkzevERn9kGzJKjHf7YSrQGFobhFWL/WZPKD9FB+ZY
K+qCVcIWyXhyr+54YM7RC07zLZvO44w7XpMbBUuxXuxDLLOl7Bcs7PJtApEU0wIZtYzeKTp87Iww
Q/wap83FjhAz0pZQHzgZ4dJRMEH23LOwL1Cp0lIweaYQHJZ4sOwoaVuZyS85TB+G0xdvcl6PgNbY
WTded8BKPWHOJiwU9RerQRiupwppvWnqbLWiaJTxWyLwNrM52uW88tdqRI7oc8EB35/YN6EGgDhH
YHIxviW9evZCfqFcHUThusVOtbNvVV6EQoTIi+TsVdhTw7hH7uvKOywInZBqsLTyJhjvuZIUo7BS
t8IfwpAHS68jga/3/05fQD4OUyuC/yxP+tNwvHAVQu8dZVmph3BF+EPRYJ8drCgc46gvOPCW8cbx
589XtahwzbFtsUz52UCxLFhYkRtQPnfDnYmGgpW4oxkp8hNsiGqzXYK3fNkvB7tmV15JFPxXRcP2
KZ1FXwJSPrdYahna6SMCYnA7/4TbdgHDr/6GZ6MLsKYL6y9VWZdwdm9P2ooysUkL+WQn8uSO6P8T
94SWTsmkU9qei3MZAYHATzOXjkJFoyAK90rf9Kp7agH03J5gmYd/RI0+9UzAb/kxtut3Ep9w4vfd
h10KkScHXCPinbBG/5Hq6eATFRXiT1eWxupH/ejJwOufjfdCSqcZux4ROJEosuWTh9w+54kP22Fn
wWwUgFAloIAHJw2al/0PfpTqTHVzKq3r2aLl3y8XDixKLgPdridhOvPkROMYkyeJkc1mwW3tuJeQ
mMjTdOzZj6gaT123rzTMXRKKwjvWfsnrEgiXJ3povGPd1kwFWx2xQpR90veC8HEuH3jej7ayqdjH
5sKcvog1KXyfN9FO/q3xlUaQBtaaiedGBJKS+BRoHmJWXNfQx9C+4cpEPjVUf/P0u66FxeYWQYxO
m1F76RtiwYUqOrXyEd3CQFZdCfG4ZMdwQRSqSOVn3rWLVR94x6lGBxnXb7iFLUg/iRDPh1PeFbPz
kzGISzHh2CGQbJPCj1V9LTrCl29ifCruc4on9UknT4jyXOLkeXXopzaGu+iEH062ERBLitRkH9IA
nDZx3dDhJJkZMuAe09aeqw/on90l9ihSAG8Ttdu901eFbDFkyvfT/30/Epo53wU1PWsr631qk+CZ
UYs+QriwYMbS0OsoRAV+1/DsO1qqA2pqro6fYDUJq1oVAFm2UK9dvW85Lg8E9WVgUYNv3SX+GEGi
dy0XDB67LOEBXWkAH4YiVBD1NU1JJOChPewuHJ7nrSGpO8kt3cJg+UeAFQbLtzQr7A0fc0lZcRK6
W5xBd6mnh9+4eOCZtU5KDqM4It50ryqUm82F1D3vaVb0KwXrgb9N7K+An4QPFk+1WxAH2zH0m/9e
VoytiNYnO6Y7rTrE4yS8h1nDHlE9QQLX63poFHRWRYvLqIFv0aTZFweBmlKMJuGNGjIqDRbVQMxO
QijMEUwxGIzjsk321k2TZE6WgrFG+xlGtvjwXtNXIFb5d5iFIaDuJmMMtnFxRxuagn1Als3CzCWs
Ik12/D69+eBmxedCjE3zZmnlu6omoDy9I80IEFM7WT0N7imIU1Jc0YCoWKVeuiYSqfkFtOxJHNf6
jii+Fekyi5vZZfRsNnoKCRsgYCynVE6yfEkMunHLphVvzmsZEnv+9tNWZ7qR+Dspmr6l4lQuznYQ
cjfYHG0tfVNfbnARHuhkT5eLD3uxDbrfFClsDEhsXdg6M9QzwqlHHbVxrh9k2/bOyVgMLEEd1zti
3qaZZbNPz7Iy84+R7Il04z1o4vmkz/781oMUZe6i5oHSFzRDxfvqGwh8myLEMK5o5+YrBI07MmTf
aQTJwQS3ZUrhNsswT2Ija3gM0BiWbw+IgkQdHVMPBqVAcc66/TSqHnuM9N/4On0bY0wVztnE4Xtp
0tNxcC1fmvLk1CaQwrZQch4r9jlR4kbxP1QFiP10T0Bgo2BrwowRHBKWwgMXEuJ9xKUfDqkqG5YP
PRPFC88/a1MilSa7itgxyEbb7yfVwmlP53piiJVs1Q1E2Naeb9M7+uMSpLKHTvtLv0SFwUhAd+wO
8zZYj6GxcMPutMAo2v8zlTZ3ltgrDrYcWeQhis0XIkN7I/dGiyuDy0hGK4Berq5pw77yTP7LL9eu
swvPRidruFqyjhIUDrzrfcAhKH+JnYSkWOiphIMkDJM1T1S8k3ire0qKJ6UT3+sjts+SMjXsbiKR
yYtDeMdAFFG2NpvVbZJVKwxgQFCtSvVPPJ5BR019EMueQw5p/vaKRg3VOUdjVLc8LRqeyLrj48ds
Tuu2nc0mMqmHGzDhrICCLeDqL928e3SWOJe8N7jlIqWTRaEqWU/Rsztnz1sZ9rVaBnIavsHl3sE3
BfU6YfKrZJv8+sYSuLhC93RM6hluQ7/2jtRQhJuR5OiiWvAoLNoTnsfJvCUrEOwkawMcLz/20NF4
xNSAVM56HBsRW7iUB6aoWNqWq20CN8nP5ycuj0f04sP3zIBOlFmkhUBK8WC9+B7hUhUyCJ6aS4Gh
i33tMpAO1ft7s9yF0Z/4sBhOjGaXXvV9M6LD4zpZKDJEbYTmnt3aGejptYC9RxeTsHotbKyVIVgj
py+uK89OPh7Di7IaYGQ/LidGOoGZQ6xTq3f8mSPR6ryfC7wGs0ri6OBQH44plpAJT5joAwcd/Rbi
lG3pl4cgPOTTrgMGuZ/FKif1L4YO7Xy3vX84zQFFYDIYiwj0wRUKDhOX/nqCDaOj4H5cmebwilBq
5slnE2htaUG/es9BoNoDt2aj+rbZ7UDgzPsyn7QbvdTo4unwyHJgaZrl5yTvJWNAbnp8d+SiNpuI
pB1YRBCW9FLKMsn3csK70qWFZ42c31kGO/BFL92OmFlxhwFrfzIVbNFwRkqrQfkuopJkv8EPWmWm
cFn7KeqsjNFZ/qjNHtBr9/gL2eW4ZLVQsyBONN4dow6z5FFqBYfOE8MBbfMBM24KXFB8mkPVDiZ4
t0+Ulv35fa/G1KJ6BJx5Wo+CSTNuDD1h+/Z/QGp5tFOlOts1wLqyZldhQ8uDtTWGjrqyZIlW/Qpc
3Jk6snIfT5/1SNlGg/R5o5VU6KWQSmQMAe5oBpnTPQXixmeqWG1UKl5piRiEztXjw94XgKJPMIXM
awiSVAU8EOU82qSKYD0y227WBsTX7auSvek88Mz6Ch/7kJST496orKt5tbYuO7sBtjwwbFGM1Ujg
r6b1LKaykOXvCmOu44F9dcqI/CVmA9z2M9Rhv4h5q9WCN5zKthC+InjkX3V4KqjKvc2erqerV5GI
ZWx/1w2ldq5R5whTOxxb3bY9pu49freKAsT0MiwWLnJRQaTKKhkSmEsk6+c4Irc3gApfbZsd0a1s
nvi82GrbFHZ6Agjs6Non7w3MvW3Zw33er0E6a66IrXL1OpES7Cig2QDu1wt3X0kIvGKIU+DRTTTG
MN0nrEGTCvBn3vWSs+0lyeOj9ygnUSBL5PO26tm0ZnRq4oRaCy2adVQLRsf3PwrVOFdnJ1SmetQT
XzM/auljAeWeSmUkJDIBFcG5fo2hTVVBPWK9CKLoOtFa+oljsg3uEXk75R5p7lv1Nuxeid9Piidm
9E6nXOWW0CTQ9pxu9uf2WvZpxCr0Nze01r2QunjEt+soeBVr/HA7NSW1MGuw9tVdS0lZnF69DmW9
WtaSGZvuw5ssQfD/Lg59gl1dc0WTnFfNWuZ0M0o9liCHdcb21DclWQELfLVFia1xF3RPg5DB2u0K
itCNS9SIilFpOI+JFpcGSN/MnXV/2P2GQSoKw0jXsNGf4l/tSk7IqX2Ztprv0wIIIPTV/Jf/MIiz
xs0E+BQnyTF0QINNhTqbYSbRz/nFJCSGAABNuv3/9KPliznwZvgaSP6D1+2ZTQoXHWWc9KyeByK/
8gOs4akv0dXugeDcp7SeFbxTD/dOzev2VqfpwuFA1F7oAKgcAmLgIXyX6BVnH0q7NusMYKizKvcR
dWpRqoZYvKEutN/4zXJHIVUCzZp1NP8LFX1/kmtmon3k7xGO42ZNzbTfjIfqtmlGCEnJVD8Y4vQH
RZrx7hksYmDvmpO8Nkdg0IQ9H4222hnd+O76ZGghvalZNzRsqaWRj1MLbbYgEnWVH41AMG2WS4fa
HQFSXMPnE9NM+LOeHJb/8p7ZOAT9VcvW9doNJRmc1ST0/6nXprlRZZxsl8wB16RkxC52h0vP9N0j
wW5QmqSueh256vkcA/nH+kfb+dWSs5lHeky6+OnAOJOZVD2L/V+m/IOAt6CWzTDUML513ZARVCsB
c4NQfLULL0ZgEhSA5LgkF2X2dEb7PRop6EjVUOViNFh0ZOmjdnadDs7jgVbKqbB8RpMuGVh++LiU
Utm2Z6EVDUpBRnLpRWdU5WUZko/oPWzDPpRl/kjFW7GhpiKEj91Pg1DhA0jVDjhG8kDiZzhsARCj
6ZB5pWWJRi1SbZMW7unsTKA4pMSscjF3RVQowJJwXkxnMPSL7asr9gRElNmcabaR9GtlmWP6DIII
FK9pQbALqAEVVj8HaWRrX8CxjtcPZznomdEia0eeaazA+MBcqLRinI37dJY8VEqgZCJXuVLFtBu7
5r0FAzV6GDPnvv/LTkCe79ZwUPw2ocpsl56YEbGl/YR+D2MQLaf7dD1DyqMrmqGD+H1fbrMd4cyK
DPCjf+j4T2ov5i8YVKCsI4TtZSbAp7mg4DG7FzRrnA0HH0YyKnoIcnDfEEYUinhVRxdZGXmTJYXe
mYCHDc8qJqK0DL96kXl5UBkXWkvlXqu3ffFSZR/xpxms2YURqnlcbXXw6JOeyO1ju+iDARFay5wu
sNmt0dtWVJEWisgPpXXukl3uNpNjohwk1+J6uSSxgty5CaC6MsPNqfkeaRlu9OLPKEO01DXD79MF
RspZJBhnt8PsxIi/lfftuHp4sq6P9EueynpthjlQHOIdhwMPsiZFGWK3l/gLei3N/dKncKbhS0VR
o4017sN1xVQninGhOegETyA5a6TFQK+JBFfWNwNWcUlfYFnMW2EOfrFq61ABdvzvgxfuqm99mB2Y
j8ZiCji8UQnKErJooSTsMYIJxJEqdrcTtDp/SIEGb+opWMnVcrbQVFuGSDzdrGKRIJaIajUb786H
4uZOYkBV+j/zqgpcR2F9qtwgChoViiGRszXqhpfUIL1KugbNpEcq6EvOCbPGi4Lgt8E8Qnb+NgJF
7oLSdYBKreoeljVNTXf+ERhUyH26/Zc0q1J6awFv5ixkjI9lXQiGX/vrBKGvqh6UNKgBoQpn0O57
umaQIs4I358T43RrhOOU21eRBU0CDRK+UforG+h8R7Hf/SZW7hLu3HIXOA6VwsqRfg2y4wSwisCl
rh2ATFtEf8wZHDVmS3PD6bZvUCOydzo70sosehMVIHKHyr+8Zt0WvTEs3dqn3vL3o3BqhE275kGj
SI9IUDZ3NNqOIG3AHpp3KoGWP406yq9jXwpHbpTG+cxYE8IFXrjFkUv8oJKd+xcCiFH75B04Vlej
Z3c+2Bwv9R9sN9LLRjo5Q1pR6vFsWZnu3d5Nv0dW9rUV2GaPnWDLkAJUndP032FLlZK4fQ66+/5m
OIHcDcKkgrfZ4T/krZdQ/rqkcQ2/yxbr73AzN0+k7OhHPg+5A10YwBaKHpEMHlVQNGP4oWBfsyny
8Wpqfw8O17v2ue3OdqVlxODzUq8uuUUQyrFzxDjgoaTsf8xqjpz3N1sjEPnNdJ0elJEbhWUyVGBB
YWUAWXT01DFj0mpwGqlMrR/DAc3+BG7M8W7g5g09stVOeS86HeRGMJzigRQixOh5KZ8rNQd+3zf7
fzHfdHMpqZ8PI0PDSFUWmLOQZTuLNtiZEwzzcw4+0d4peA4l/7IOEgyFHAMOXYeTXL5cRybkts43
IY7n86toSCFMJtzZoqeFt7/MnSTTYpN7tdgNWjt+2Y/cU3D42WGB8aIAIICKoB23MvIptsfxogS6
kz2y1OiNGeiBJ/zxHdRaxj8/+XxzypYShu3iTUYTUohgZnmf06G+51aaWrMMpHkq/JpgtMEe/mqX
lX07C06N9AA3iEtUDGV/aCrTt6Ac7GhuV2+z8rPCHGFDB6yvPOkL11NvkoSz6lr1eflQQ5A+korG
wHJUPTpVy1XcG0yKMZo2GFibwVwGtLp9zIoVL+44As4/3MGRGWSxUY8axs+vUDNcSrMZLByiWwHP
Oo6VsoqSbGnSAZ/C7FhXIwOxEKc1Oq9CPyLKfoKheiQr7/rbdFze04N/RFU6M6e7SImb/8srkSzK
qxlmkPlNjeHok7t3pC+wxOcwlh5I4dX2kWSQtCBBwcLHl5ecVTB0xOvbNl9a+hTK2RJiSa+DwLQ7
Uu/zFWsmA4cP4TatxZvf0+QOa8uiJP5VJy+5T3huXtHUAlXF15J0i4M0PAtbC0t/R7aiIy/v3TtU
oR5rbaEcJEtLYYXeY3YL8IaKH7cK7MpdIFoosbu7BaBQwuF+XO9EahES1hJmnuBZ0IWa5Evk11L+
nG3ggSeQhj4uSpwBGZLjd8qcOQAmYxfQKaDmz/MLw/F+x9ZZRGTYrfLJpnHwjEg+NLb4dVreby0d
vAvTXWLKYLqhOqc5DXYI8BH/UcOl90qRwQn4hNBdFS8XNTLi3mhXOZFx9GJI/FO4KOuREJk9DEBP
Htr89Gp5KSITfaEeOVTefmStd+Jq0ZOC8aKnwoUPRzLtcjN3T2vPHE2Iu+l5ZG20drlSLiWca+Zo
eagMGe6U6ps9uh6lsCZc7n0NLdFs+BP01qdEgInA2A1UkQBgGUhDdqAEOme1cqBuXW+YzNnCaS/q
1fuDxiGa5Rpfqxu0TfqQGwdtzzttNELaY/dmPZYv2fUDrjzJ4DKMvhNYrJ38CVmj8WpNdAIuSv69
UymX1ybJ+3rABI7BGtlH1cwFYbF1QkirG99C7jKqgKA9aUrVb4fAy6Mnt1YnoMuO4+UMXjHdCaaZ
jVCkCumeQ3O31vMitta0jcmSY3+00FpW5KE5P76ssTQCEkoGox/S2Jvw8dRfLs5jw98PkN327yUR
dM6v+wDNr/FD7N8QnF5BajP6sJz5FaI3bVTmjnX8xkJZD6a46PBNr7ufH2zcQ7XCEibhn+nqa196
KD1N+b8Ht/R1+fYcakJZFLwEyA6IxXkk6XnMKVi8uI/6eLAmJPmdPLQ+LmDe4YBMzLIqCpU/GKPD
sa87wlrdAXlOhLBQZoaOXTE8+vFhk9MAqVQglRmnaZkXVQr56eW/MHL2sNjv35H4eHGeqW/nCZkr
wlsVZ2tpJQg9Wgs0IzzOvihoQnPdoODv7TYjlaQCkpfXfg+98dDYF8XRGZkWUUg8m/03e2cX/nbb
K502uqgYYwD1rm8gTsEZbDRBwu9HCtRzaBExY83ukO9wTT3n4zqG6khvE1dlh3ZAiRldZCqGom24
AffOKX8thGvnqVfeHeSuDOPuslRmOyDVPJJGVYGOpT5yLsPaRMhgXdRw3rdk2EfLQDH7VyU5wExF
bUB1a5wXvM4QsPKlm61TSYid4TBSNY7OjzzTljiZzJTdambidGDu3lJ/7hYNZae4ODN6jAEi9Few
LXMnHN2Y0d0lod/UPeep4ZCHnPooHtbXbtYqbipKV+7Rfq6S9EU8oNrmT/kM1Ew48HxIMlCqY4sp
LNI6f4aTehCi4xoJIXeWAoufXpaq59YfXJpYzrAThb0gzVfP/MGSjcNGu/XI10SXxIsJDAU2S2hY
r7IvYu6EpyMKnSVrtw1zUlpwotmpT3b5ToKeU6ne8lEtrt+ee+YtAD8LjoxjcIMnqx7nDTELWcH+
E2mx31U3Hop5m/8uGZIRVlWXXPocgXK52eKo2ufYaEHspkRleyYBTs+EPqAgZ/1pMdZA3n07jLnA
s7+tLXja1thQPXOQ+c54B1jx2POFp6PFnOe99kEzHcdOJPk6hTM4Uk4y71hXWLHQfY3WEdZcshh2
Aw/CXoc7BGNUAKJUddu+CGZfAoshuSH5azM9o60ojBC++FbJObNuLTr6lS7I2HgoNJLg5mPNCAbt
mGy8gf8nm5a3G1CmNv3nVp0IYvvEGT5CVUyus43scqRpdZsMnc2pR3bMnHyF2x1HAJP679CCroTr
DgcAbZejE7VORloecIO0XdseaPl6g3X1u2bzNVDbw8cdkTVGfbZwBdRTZtSln1vphykK/km8ypoh
sGHD4yoKR27C7CwEPvKxgaUXh40zIlwDuYPTCJ45L3E0I8pUsaARng8UW/thrnmfuT3GJqrGttbg
H+fsdc534p6mPspmfb5jA8LF/WoY/qstoplSTO6WuFFpriMXP3GOLc18QoE93XMxoAHniES/Kkn9
qjxvg+0VVDAinGTeICRZc4N5C0Fng8mLisJX0AL4R9VownhdIzR2PS/n15K9G5cQV0xjS1/izHoC
XkkBN4tmvsW1xQ2tIDG4xpGdgh6PlvdXNBHw+vXONlGkNNxRsm541jC1HLe1udXGNzcx1zU7Xpz7
IaQwxi5TW7uBhVup1vAeeG7wDzQ+MS1XotWHGNig/kwvBc3l/b+RF9KFFTo8WCloO7sNrTNDcXXc
HgNs8bj0RAeF4sWWyk0BtG8XjbTbrCAK7iPx2NqLoK2KTHiwz7MZNpUQMQWKDN1Sx6WGNxDhLgvV
YnQorlCaTDAa+C5qLDC9drIpv0+2wwZ/hlI7wWCRxoudyhTRc/hJTe1GBeCd6vAxr1eHa0Abp5jB
7twwPckRejHVinbK4663LvuC7oW0bUvIpFb6zEPLxbiVYQHG54+bdysRub1BZgz2f/QAXaGVZNmE
9EYIedEhaH2T2ROZkc5lkVcroMot5HGvp0Vm0rYwxoRPUlvTFKplEX5dyd9TeNufxSc8Fo5Od0tp
Yqhsks6XrwGq0/0pXSWSAzTWUZGe8FL5relOewvpqkHqzb9rkJMY6Q+habdYhmZCJvGgF975EZO9
feUHOG7SIP3U8QQEtJzSFjs3vArf23KojR3elmGlh2eQ/TDzwQ+O3IzY8tqVOJYjfPcVufdiOPAy
atcsHL/CM9p2k9XWtqcCJnVpyhSDDqQ4JGWX1B43YKB7J03pK7yLQaLycRVtE2/NoOX5+qooRfq1
LnIRBbcrd05aAizog6h1ZzPIaG3ItpxjGX4Nodw3R3hHSp/9jrPFF7mJqQkmI/7JEaNzZkYtur9m
crqX31RibgJrdh/RdE10tO4KHJjauTiaV1BezT0Tc1Hsi9ry0UGOHPeY7klUN2IMzAiGdvOixLhs
Gkg/++j+U5+1WrD0r7S/rlYnAkIdg8+WwbNHXGtdE9pGIHB9eX3vlRFpobINRjD7eHUpoTc2qDbc
PG7K346tWN+4fzcALc0I4V4emJ2243184wOlwad/mlHBDBRJQoOYG6vXhETaiWAzwslSjAq2q0hU
eWMDQ2qOP7r/qlxc2513hWy9s64DCEuqtJTPQs18jS4D7YEvEDoMREBoIbiuhmEwxV8v3U4bfFqw
W9DGK8fw5gf0Kz3kPZRSqnMsxhQgsHYlIf+Pc+F80nUNjxqf0xSbpw7l9mLpovl9XaNl1weIT6Wn
z4nMcc75Yu+6VWqlas8RSjUjpuSQDb+rCdBihGh4e7M1Qva3BPvtD0J69SvQD4hOYUMYikj83ZRS
o9zEgCzJgMFlrqsPrSfeRIQ/eCSxztsoQNXiFidQapld91vomw55sBdnoL37VUl79/bw7H6v7/uo
8GOK0qArkhg/RNtxV79Z0GDfwVi939R3CkMW/l06J9Lyt6BYdKAwsWYxGVngs0HLaHuOY7fF+Bpz
vxAwVqhZJq+R6XE2fu3NTPhyCk5Rwvu2oQtlhFPGBoH9yLeUPtrukIh122VwtpLrZuwbJtLmtsYS
af46xH1Wd5LF19gA6S4dOK1AY1LL0V0pK3ogbdhKTZp/dVZDyzdJlvkYOrY2y4azy0GqWcp+i1ql
7zn+VXEoAVzEt6TqrUt5/qg7Da1QXi86BTTGJ4fr/Pr8INUXq7DuMvACtfYBZRfbL0N0uW7hVO27
8D/yuMpAUKGwu+T1HNulp4G4jpUd1hHmfFRSZEflzMJetoqF9SWmRGYCArG3LP0VT4S3dl0dXTo4
wSrq9ObpvkWV0/neVVtci7DhRn8EBZhe2EOp1vcj1WJXRZJXsTJc6jCyli6HHGPr+k7w0ZgAk4cx
MGBMO8ofXWfXSdL3oegOn0svXYfHDaDBWXN/Jq4sBrLYbnxbMAo2X02sBw0If5pbDXTiK1MgeYWZ
S/oFR3w3aCjm3h3yDjwbag6I9zB2ncvZpLKkebMaULHXzrnb35q7Q7LG5hR4K+30h4jLgqR8uTUy
UMrWIXwdZpjverEeHMTbKkIJKdbBYtf9xojdFHwVkXQaE9YyiTjjTrvdXg4HNs7KErdXxh1ICtl9
WJ5CQEocrk4FLStpJSVhz2mCns9K46ZkspIpwt6HSI/3pPJV47kFObWgXkE71NVOkgTk9pSfb56P
NePhVYNPWSAUe0I2RCsqtQpBwc0TOfq3nThEJpqH5BNwMQOr+0D8KUjyXFBObMfBW8x1hCJtNuYH
jDdkkvSeF7l6nFJ1uItzq5elgWIBjoSd8O8Lqm4SpMos4vsb8+4GzbUwalTwfavEYhc+SqNLDiE1
HTGVwW6LSsFcf8AAEkE3ZzhKWEVbiwlrZXZ9454s3mHXqyXVRjpNelfvOU11gxz7FEC804eVj64m
naUPJd9PbKnVJ+I/FTmdajMu+/M/o870hlgkh260f9y7XARqHeDUX+ZxVB31eKK3J7EtQWWWOExl
kOTJ0Cwf5EFDhBBaUu6EWPZH2sXW+x9bOqWWG+RIAVERsZs4zsu7pG/Oudei5pHT3Hc84kuCaZtO
0S1Y/ZKFf88nBfMLVkvsFee7vtIGI8tWhnujcex4dqXwAO87jMFweE0MjeQxxedWhUE/ouJFg/6+
oCyxfkiSqEao5trkmr5nD9+oPprT3WDRHywddwtIYUfVmpcKSLWqRMkKJiUgm5H4izVvVoMA7rPE
I0gP5Cvg3d0zMLbCnWlIw2EEJuOGweRyiSeGAuPRQEI9fKG5X9MrEv+qGGGqNSmGD5DpK35ieU9O
apU0+ym8/yNR9K+dvd5+SbauDHNm/FrlYsNJNMnfKcdMVETjuMkxlGMdPSZh+gE6w4Ex9PQzXxtu
s123wMIELfEvpHtoMXEFjllo6YCePqORzA6AIEa+B/wf5PCX2qR2MN6xLcS2ggNL4D2toDo2Vilu
r3o5uQ8Al2gUI5EQohX7F3IGtb+p6D4doszranlUKEUgHVgA4Q+9+GD7Vdf5QwvduLTiz0vf/Smm
8sLyQAxPpLj5YfDGTomFtIQpvvcEJm0uSj+cK2MG+yApINMCEBTKG6/Hu0A4PPD/A7gNfq3qZgMG
PQlYmaFmNld9+/qCTts924PHZo9vV6z8i2svu16jiXVW+s/7jVgZSKyUBbxWsFa1izFDbuzD9elB
lAFWRP+n9upusd2uDp6pFgR9/kYivVId3RGRTL0Wfn4bYB4AwmrfU81F/alu3rfdoCnuVtpBcpJ/
aDkplV515QQz0d1FIeevfUabJxU6kng4fiqMUmqOaoPGNJ3yrbiVwfJy5uu6/0HsoASWKDoeCnN1
Tej2KYsCkPV1nZ4zhNXsGvAEjHu37QhWbR9LhSSUzC18se9gKUyJ4JCimUfaMyE6nr2cAzPcKMUm
kUSDE0VX3yeSAMldvZmva71ciIwaE0AtZ3hDe1NXwFGciwyf/3W3LB3BPMOJLFqDhnsrBUm8S8iH
l3XxSTsVpC73xUtX30GD0Xh4NKRbtAKkV+2qcCopY5a+Ef9tbP6hgq3Zy2LKsEhboCyriVRx9ggL
mH5WN1cKQlaiFXojp9YuBEQtdCSmKDPIUbDVR8u9Vm46g6lev78aJYMxHtzqesgakZ7EcYxP1emM
II9U/SOw4EDVsKlNZRmhVe+iUUiuukwVlCYNoKvrfBhVzKHKk+3qXCJLcXHPu8oBflgmJm8Gjdhi
23kMtlyHUjkfeDlajZ36v3OQGUiIbE8jf+73Yf6BZWZd63zzY4ZbpcBvGhS0qOp3AnmR3e0MSwWC
iJvGUeWbtuXFVTj9FiFqxuBCV3NZ2+80vka7nXagcmp4vNDYX5QaLSsteE3kwMZFXBz+22t3W+hR
S5SeewNY/naTh41g/meITDDJVR68UlL/x5zqUrPwtfm6P4aPL3G+sKxgcxZMAaGy7hkKUkF8SUER
FIF19aKlatyQzr/Rv8gAAVO+RziADShcx28/7pNHKO74qOf5oJ0JuibSzWmLQg624MNks6nwOYys
GzL+xW9Xudy+L5bMT9JxtYfeg2smaiThYC6WLbHOZR3VcUPQG0pgV+I0NkCTWya1IqSYWqCttaNa
lj4maNKeV+LZ+7wM+pf4YZylOU67T2CJWwMWgtlwNjPpNL3sSD2/ApVNSkiGAuedaoxTfPsZIFbg
RZrlL1d9U/U491ZzoVkKas+duRU9qTcNHl5NYW3S85hrD/mPDjzr2VhbgAx4tCjgDJX+hGGknsZM
mZCM7ZWMlGmFPdzIQn5gRB93+uT/H7DF1i/atKGCE7+7/sZFGj60kEIGu7/47S8mRI5jYnmHEVrO
1bdN2A33kDBTCTmMeB9oA3RgVxOuoxefdQpQLcKZbubYnSWZ/wjezZl9iftnf2L6XfdWA4MMU22d
RgBhuzJSiJdS7ovwlnh40JQLF5Eiw1Bs4WcPbY6THN/F7HsdPWjZAwIG1hkzV+Hr7iSK1QRfasPV
UcGl4+D9iGyIK8x83/JqKP2ISWgH2CvBU+y7Sa+dMQYoI7AielRr0lDgnQJg4Lm88n20o/4S+MvW
BLQIxkpQzh5VM9fKUE3tRA9LzL0SP0cCEyjqVsGW7O8DZjFDsDbfkig/O/oyoMhJWlO/eU19zJsw
nMGKr3EKZ6PqaaLEcG2b2XiKU48mjOKS85pdz9UCdMtacw5zBiuzaVvu2bUW4UItOGj7bgXTuceA
bNe7A8JHet0hq9AAD9B02qdRVHQC9NAcimY7K7G0gmVv4gccidZ927i1tfdBB+FxGZh9joyGWyYU
iDkMVvZMcWMIcBZEOCgT1xR/RE5YAR21TzoQpD5T5GM36qvEucjc2VzdOPXr/MyFvoYKLaQxsw8s
42P+GNZqbYUfPGW/jVV65z6Ry8Prmg2qKBu/D4cPBhMVM2U0hcLgRkzAZG7dsQl3RIn5YcSOiMp2
O8ksfgyKFOX/yxGcJkoA8rZWTCk17jv/TkObnT2eUImpIRf00dhOBU2rydHDpiRDDJDqsMHqML1v
hdAjFs3mzKwiHJIQjdelDvKEgvQ6njZB6Z2t5nCaHzldlx58x0NUaX4n25NRZmU+K8rF8x/LCfTx
/m+GksoWaiBXEW8bkTt53EserpV5o2dFCgFY0yLdKTkTo6umUW7IxQbixSMb8R4X1fkwxG8kDF2l
4G2X7b+y/8ZkoyExyLyNNsTSOOoejjDASBgv5+F/JN2OETNCVojphBx3fjs+nMRqcuzkmhmwbbYs
Z5SOYtkba7b/Kfx74Ckk7suZfZ20Jpke44ku9tzbQQecVWssMaLKxcrxRtoYW5bMaqrHElFlLzTQ
/Yoz25lEwSmmOfd4OmrQC/MIGmJ3v3XYAP0ev93VKvlck3uBz97FgEzVDlKblZMvR/H/V6dtVA5l
lLyvtPBJ+YVVFG7duir6tb7ZXd67pncRo5jycY6Bo+e+qX0Pmcub7V91e1R4i3bvXapbzAld2uAk
nrwbnn3mhjZz9PabjaJwjLj8+y84vufDLAiLSf5RSe6gKIuQsPWlrY0pgMa6lhg5fzMokOWig63H
AFtgDkySxeEL6vHEK4r7HSPEvoHOvPUTDeYpt1Qv9THyOxjMqNCoki3S2LrKwfbyLJ05hK2EVNYs
DB4Ws7fxwNqD9HXe/qKPfqrWIrxMDQ4bAjfvmGm9LJqyCLgj3y4BoQjOnfEx0AEiA/Zcf603a7La
zV205pPXAh8laItQYv9sdnjygVsIlHRIsYsMuavFdfP5qIzVEWZgOnVHDJicTn2pTkvcuW5zLTJo
J6E2xkC1snxIyjsW3i4wIbBb5wZ0ig3YY0soQ1UXWfckdyCWCDu3kbNRCITpzoLiPkI5znYNdizy
CAGDc15x2URMwtgJqsUlAwJVZ0YXwvwz6nRVXpqijzD3GfoWnVdylQTzlU+kT2SqJuXiujFSTOI4
c1yadi9Fm4l01Rc+A+hKuYurtIQ3DYVLbtQn/on8wtCmQYPrq/yMAEN9/aDgi/lnc1maRv5tclmc
hfzgjSFRbNcwkzQiCeKC7th6T/6KJWGAntfaQgc10kUlILkT/uldAWkDBODAhRLftz6HxzSpPs++
hkos5Vd8GjlKb5nZsYnsamkyo7QgILpz/FpPXd9mtMDewUtGy2G3PD6eZiClMsznXHVFkWpqulkF
Q8sHv/Nkc729UMKJQ1N4oKGsFNVSy2GEi2tOdKGD6jb8ayjSJo2807IQ6F5pBMdSGyJP2momZY9Z
JwNHiTJz8w36Gwy/il3a952OLfb77/IVptqcPRC1mt2avaapM1AVPrc8QXT+m0CISihuV4LRRkz0
H4WOtkvcKt7WnHbjgWEupbBADQv4aiQiNzakIc/+z6NBCJwC1BNbkmP4VbHnVZf25la+33pnkh3I
LB+Nm0g25VFM7VflUhG0tzTk4xqBAQjqahj7scOGQjGV+4aNLqDRXtSBZJDkvnsi9azXhrcLGt4N
saCv1zhNq569jLITt3cWcmTCABrUl7ekMaBAaoAI3XPnLNCCWpwYdbS+rkzYqvBtovQfHfoa+eit
pqXcNfMSgGkeDNmSff3Tp5joviWqgoKrgi1V42iSSqbQ6+1nD8240v7B6ueJbfg+Mh2A8o16qbUX
5sYh6tMuPxT2/2KzCiXSNAHfq/vh4yNuU9StqBNQz2CBk01Fptz9SRFkc47TJn3PUeBJeyFa47wX
aQuIcsXX7kYUCEKn9f3GW04KpvsS8jcog4IseaRHToDBKhvdAceqAPP49+QMkcUqOrXk0CvkocpV
X35BdNzEXBuiuK7sQ+tU0wKYfzSL/rCgajN37Sd3LAyCulA48a9P+Vr3msz5AiBVEpcdlseUFdYw
VZVEI/iX0X/uMk961Kcls9RSAgVddmnuNTdeKoJCN/QyTDWp3TDZl3s3d3rYEZXbvcI+8pYRQhJh
dW2M0HCpCNdGvKv44S2vFyX8dHzLQEvBNvKLPOmjCZYQ9S3aY3Uc7DC+Efy7yzfXkRhEm+V/OiTE
lqcEXSJVWnIgFbeNqJwpYTY+3/xcnVl3KgCcHCw5EvZmFhguW6ga6GpdTbCC1WIa+W43+FTDO2Ta
h/tpjt8ZqiDQ31PNNnN8KdQhXw3nUOXKxABW9eNvULaHG8C1afjudl1VIv9BIQqd5SbnOY5tbnF5
Hmen/MWSlwLvt2Pdg5dk2sUe2uNN1Lq/qT6xJXzyOniJxF2ruityYv2Ngqa/PnNFcxGUCx2OHCWq
I++pXp2t0Sbvp4IGD3eAQbSo6ijAsxYqcilt/yjl+h3ap6yqptBIA5yGbhi5yuVR6kW8un6BDA2A
yw4+cdqhFie5R1S04m7DZJNV9o8LrYDsbtxYq3YRbmdPmmYg4nqzw7vPBA79tfBX+yzMAdLifCvn
6BExQ31GYprRFWYAqNCdA9EoSGBsFF1QNwIyEDicRPKQ2PQMRCUbZ4Xcw3aEsmfWD61cdQ3XLhkh
hB7VnbStBZ9Er2IaUUeMHyicLLFqaBpAOz+dS/oLtY3+YqJTDSy/+UKFkGwx3r9/LqiaBc2WrGT7
Hl7JNCOJg8p8rNZA8C9HYGfjrgOWgElV0FKowlFRe57PQjB+CHRVDLb2KP66fzjaMjnU+DDv21MJ
6HkUidfyAN8KfafMZ4C9IycuEy83pwYy4qmgvAbUif3Ye3E8UAXWxzlt4GvwaOOynS3kOTwGcA6w
UdK4tKO7EHbZrpYMxajDnLXST3IEeYPDXw/j7EUvtVqYmbMb+X3OYz8PVw3+CfcjLhScTBHIAxQP
84sKwMWyoPY3LgkspFY7QFd9DkeeJW2Ur2yeYLkvJdn0GqmI/nYkNdRQM9MBibH5XBefhKFmUGLv
+wZzyE8WDkHOI1jUFynqyAIXyGZY95gukcCGr5lvBfCFgmsavQPv5v9swTDzB0Nsl39aZEMEMIlH
noq4EB95fpb8E0YQlZU1wiUJzzFcf2oeIGWQi45HMRmqBMTsTVRqQcL0lO2+xHfSKZydunquy/1r
qsuOjgtg+oIkha4an+MKrKE/d9rYmTz5Odd/ybVilUmY7CRnvT7SB7eJeqYgxXs5a8gfufP5VTsn
DR7XckCFE5h3kAJQ6rgg2NWtmADtlZ9qW8H98kO0wDhKGvxUoJsvArgAXbZqeCt7OvgXN1BoN/5G
qnzUdFRaIL/u2Skezv60TRw3ZB7zQNY3ziYmqksoQnds+s1xTueYcdpXFloAJNrVw85uV8VnoQ2G
RJfGXpSeGg3atAFBvH9BEejCxVp++DkRE4vJwYh0G7aXbajmvuO8iqzL5QOh0At/A/NuE4s1P+2m
KIQBHNphqE2mPO2InGw7GCd5Ey8nvpDgvPu+9RM5qVk9m1qVwHrX+NMPMGlN45jf+FPTcje+6zU6
7mEychp23wE0ov79s2sIhff2KwU7NCNSh/wuN0689wkLJklRfInhxMP1gjDSgORSjA2Zeaa8U18y
FCm5zERAq4xrW3zTr4ptyywAW19ifGg0zFPFTjSYfL/I/KtAFrv3FLSrKlLbcAnwUgm9Tc195T/c
2XLmIDyxXKNvsGMXzSiOkYMnpKz7eBtMYsxApLKuSyWUWgmBje2HcpaWhNJom5q8whefelyiCE+K
+rcbYnDT5Hj0TLBECBZCdKj1d9PXawnhoFK+1dzXR2VYFRB7srX9uMQXQuz7+PS+O/+L9s3o2mny
hYatcpK2eB9c/5ZL28PErxzZ89lUFgWt1oUW1jhNXbsuXXeJxlL8HODBAxDigBIhIbjhmxiUz40b
7O9cZccq4ulY9no3V5K21/H6EWzPrSI5w6kfIfIiu8ln0uusaWa9tr/knkN0lSiN12hoLRAEnecr
shjyUu/mO5FgxlcJ6jzkxhO0iVevNsXVE6zDy2WDLZKaqmNdMVH5Jq0pk6q25HEzu8FRKrxksIMe
6UjdJhnA42a4T4tPnqoACuzqgoXpaDo7u7/9erR4v3Bn4wj1YQG8c3d41BaKcZKeT5slzwF301+O
GN4gg50sfy9qeE5rTjJ9VfO7uQy1bOQuZF4sMpFD1ZT9rBDh12c9CBNWWJ5wjuXxtRMeA6TI0pOw
hw4rNDA+g5ybpkoiho/XxQZfCsQu9S0hIAZYJcZiQt05zL8Nj3NXCea+biYGYPhUK+ip1IjzNO95
7SqFcGvyaIyqAWZ4Y3F75bB9W/UV7oqLpcQVMMETY9VQKXqx/YbsKxlN/PMSXqWXxPUn0w4Axvi5
/I3TtOv4iRlWx41U7rPeMUDRMUBU8xshGSPV7VchIqHFc0WE9H5q2f7Tcb63+PLKW3EidDMzxNZW
IhV/k6sxaQigndjzS81e0GZIdduze1eUDsY958OOLW5WZisknBWU4tmZ61K7ETP58ePipRbX8nii
jW4TZrvSVpt3wdYUKZ6xEXWV/Nv7iHyt0MBUk+GqlMF0vLntVfMxbHSIqmYab2cDaQWZu8jHIlNG
HKi1hCXg/N3eWEaNDurM46oWrC7Tq7soFtu6yaaqku5lRYflmPwdIDKJw3CFGuFC511m5Gs6Fl7C
I/FGcKzAtzbQZBuqS/0kGQrjZkp1a1/jVHQXrFVavkDQFxadrmMYkqboXYk2c5Wm3rQf7HLDiPRv
+xTxle3ZM2uV6gJkhDZNLLcF797md6YyKrY6hdMQBbvSB7o9tupLWmZSo41h9YcF3cmiEbUCp9Uy
z+2R3uDuX5wZeNFXJhZW3DN9ZobAvRggNgdcSxThKVBunISlckzl1L+l4FZpbWawTQ5pzbXmNEuQ
eH9eOJCF4jx5HBF8+BqtDkwAC9UKGTdLpDSoFHrrcFK6itoe1N85tS6JAa+uUg7+cOZphKtVd+Y0
jkkvFZpL93GBqE4pNk2vYePXY+L2HkOa95kKPt8dxMeMroQUVdMYkx70hq5cK8tHDiUTXO9cdmWW
RP12oOySd3c2WUN4aQQfmbMynnTisDkHO6IbcQYcsdcIDhtDxFcAm0wU1/EhgC+f9ZyDIfuk4bNM
WhNijq9jp2s34rugzZvHhmzqQSLo3Tq0GvsTEoEGeMrFvi99rqhf/VUFG2G3gOIbpK6Axr4Y89iM
rqF3v9BtOz80avpneGUPLOlas+9sRdVj7UYjxknE7g2yB63scsBBR1QgJxB3/dtiFL3r2hsDw2Ri
a+Kyeure2EL69f/fim2B0tiC6JDJBqKYJwn5YuY06VpbJdmtj0H3xO59hHUIFYRBkCCfs18mZ9Hn
So2J36U+jmn+HfvdjARRTbzFHlPDZ4hZEW8K/GPS27jUFd7zqX9+CKB8FUxsqSKrmWzPCfU75Zij
tHAeZ8ViYn8Nh2P5gItX/uJBrY/EtYtYkbvA8vTc4xzo1txNAoRymTPHExhLDsUG5hS2rbZhP0+H
4iNQLN4sr4pUbniFMKNU/Ol4j1E3so4a9uq005lUYcDcAM2BG+8EAx63LNP3sesIRx9Qpcm/i0qf
xK/553pVQj41YeUqVQmFfgt8nOd3MZJYBlLcoGkCEPlo27fcCVL4poFR/v+uhSBnN1zW64UjxaFN
juxoKWMO7ELWNqNnxOWlaBzcs6INR/Qdkm87qt0L/P7hnx79OdvGQ72JvyeEwskHMsHXT67Gm3fL
slBWFZ/ZzxsmBWFu0sty7s5R3PHOtnAD3rY082ZptOMlkMaW5PoCUHEwi/0dcVFVWgL/X53TfUbe
xXOHjvmLXpnStAxR70aDpqYtZAs1Q9a7lkzpFzUeFVrTV1e24LcU68963e+EtRJRtk/YppbGDFvr
KXLDNy5elnuEElJhwqvDbVnbC7pDjcBSKf+a85FIgsZi0d6bA4kmU9/HKQutb2VXfVoMIw2Wnlxc
YbcuaZbQWF1/jViWJ2V7JJCv/J9Mkjrlw9aYzgXEo71fPlaOrHDbd9u/gZF+vW7eUYiCMOfBX0nN
tOVr78pF8k9zRsS9kPtmNyFL2FPAvZ0Z6ptcMpWS+PR1a9wboKCYV8JOuYoys+5TxHq6mlaDrU1D
uGwWaS984Fx55fo5yT1FsUTXpTLyLAJQeILINRrZyi9LyScPdkz64MiefW7bpGeCqvbX/zIqOt0l
hMl9FMsT5GbI+KHT0ak0KvY8oaLbt73r/chhmd+r19KSSdXKuOQlExJbOeKwnzsYGQqkhmIw4dr3
SrCtmTvVlTJ+jpZCYw7iHRq7niJsYQJOlhfgB2XdBJtWC1RZ1VQmY05QDBEJgCiyA4WFG3GqOBDu
ArG9D1ltmCy71LG4uvemOahwRkgfqxWx+1sfYoi3qtur8INYWZMpCRldSg+Xk+MMbNaPU+VtH9Xg
8sMl3g3g23ztkY/Ooo8XodmrOGix0Sk2MAtCII/dtLrSb025UU+2fdQH2wZ+Xsr4XQL7eDAEnGv2
Pc9oILgMJBKDTTd2vaHv2hbXE8v4tkxSuEl0ThL/UP5CiteT76kXQUKoQ7ynOdDzssZEw6/QGStO
oh4LgF0bgxhBsc9r0Z2pe+I9ioASbWqP7O9UUMA7FkgIhp9GQStdzTYP4W0q21AFz52oiCXBuB87
bRi/aG42M7RdCQEhc4jaxIw0nLxy5icDY9ZwV2+Q+eUMwRpbqs/vFFzg2jbLLFveznPDe+CbVDYq
upLbV0bVNw4HCSrKIIx3g5kJIG29GaO0UBslDIl/FLflCT5ScZNzoV9pmMphed/2RtkcxgBEcPO1
27PTAlahojZmmqDWZPuTUFfC9dR8IYzQCMKX7ppAUA35aGmS/huaXm7zogC7FjUC+4+lLLu/MD51
V/YBCH27HM8SuzoKrn9pUhO41XnlXtHe1+nBlAepLy14Ne2KLKDdRgUaUS9+GLiAMXln8QFAqSlx
0ACOgM6JtNLcuha/zRNz2gjpIpmXjpiphezZZW5YzG72wngLgCXdKIb4I0rAH3Oc8brkYHde6K+s
GagePiIFIH8t3ybM6GRvj08nyq5dSbEfbCT7LXeB2QymF4jA8ooGgqzSWv2Dv7J0/P/h3YWbuEdx
4Rd39UvU7NJGWWQNsrDE8xA5UHsuMbe+TSAMi1hZj7ka+CqrApE8MSa6Fv2f6MYLmkBWyLr6D7ph
4wtVVHy0kEW0NrWvX8+WAZcxOLLVyyrPDMzc0h+yaWMWJrmcrFWi/s4/tSvdxFNCgCQWmMMxmkQC
xE2L1ng/t384fxH8bYVxNol161U+GCI5M7eksMC5O3mv/+fMzJBw1IC5h4iMHNesHfsewm3fSVXR
ko8r+ltPgYeUr6rH91m4r7oD6CcdNmsrDNY9Osrco/aXZNqmkX3Kc8OBoDcG5N+4E+/kYru0r0w9
FhCDAC4xQfgIpVqyzO6tOuoRiIaIeZDYNiDcLApJ9rIfMHZ3m5tHtcoRyDb4MZStwXSNwPIOnMrs
6Y3tE/d+hjdnqwq4M/p8ctZghNbeNFUbC8edFgDNjKxOkGib783Mf4XiJVyuCPlDvTrZnHSFeSSu
uWqOPVvPqTpoDgTFGVj7jQeQzFc/t2APRgd8Plll6dAGnLFaFr4W3x2T0sZKCDGnlF382zKhjTaw
NtJo93gVdULjut3TyZye06NJyYn1fKr2myaZJud/lPOjDm2kS/3yGTVd+8IS/vdEA0Px0LcxYk+4
Pvj/f7b5/IGZx+9nlO3vn36na5NmFDOiRARvNu1/G5rBrXNoVG93Ez1rpThpbcZqh7X4Dnrhvz9D
iqM13LhTdiqlAJPCmPjuh1zb0GDF7V9rgPqgj2yI36bctFiWHVAJBjIW1l8QO0qyzMK9Z3G7SJRs
wJeoLhOFYcDnilp7vhFcARiuSNMpo37+4fOxJoxZa408OXJpyMrasFD3Qp0zlNa+g1843Hw5qFOz
e18SV0fjVJ2OnbHMlhRocrij1/PHIBCYRoq16qHttQ+9IOHffFDOYumzda2bbTKL11WaUuyrFfzF
14+VwT/tPtVJ/q1wowSsuDptW4AHZM/UOJKxGkZIXXlfO9TYL3Qiz5dOevf9crpFO943tdtzsiT+
xHFdIP/Fwh4I86kcHRA6EObikCP6xubhVfcnkczYHdzZrPQq4Zuv+sMU+m6Gnxb0pERhUOnsYihY
Qw4Po44+P/V+5w6OXSrwttc2gRJmh8g1K2MYXsI7FNWk/5kJSMVoqy8vipGQvvgqStIIoq0QkyMx
nVkN9udoObQFAR1WVJBVVUhIaBLIviXbVMKU/wO7l6TTqqSrjPwCPzB+TGP+qOSrtJ9Z+N/utEKX
XLFP6TRTpNS1oGolVrQkZJ9Id7jp3Er7P21Zdp61rK4t1PRhaPDQhwl1+16TcQtrJy69xbM5alzi
9ckbuLX+ICTKDkhyefOKqDjR8etlTDISzoHQEIznDr4XU+ni3A3ZcVqds+uKYOJTzdUti2vo+yxC
/mNd8DtCaytX5tqBRqjuvEtgW6fCbab36PsX4f0hBqXbFVWjN8AFSwBtGT8zbdJiTxBEgEcZkoEg
bhd8zoSGlKmyi3mE/7KJ2bhImTVs1lMvepTtFm/FzlfQ7tdVA9IwM98IgX7cXpEyWkbEf4DBp/Hz
7Jtlpx/HDMPrk234y755mCm4y1EDR4nsoYcBUm6TDMgPz+ID1FOn3GboAk30nKOIH0Rsxq9ZKrtP
3hy0Mf4Q0zRgjwJTUUdRJ0ZjDZMVIHhDUuMWPn4nmEutMP8GyBYnLvM8lZFsHER+On1LJ2U9QcqV
eqKU0Ikuxbmw+n4HYjfx7bZF0tkqRPE9CAWlL+TJWtOj/QOrmsMwKAU2+dzFfmtGZvWaF7Lxwf/Z
yon5HQoejMWwr69skJYJYTHfTaNoyFaCeBl9P17fC1WfavWcoPVzKPMtGp+c7zjR9EuhkLiKlIxn
1MbDAgZAxNF8JG5dp0girnU5guYpsWneixqeEuv0GJz3p5dYYCPeTMe+5iVKKwg/VCg/yeJOlDNy
0Y6pOxcwgCuXklAxLCb8LFWm+8ejhcij/vaZp7EAzcHgUjvEFRJME0p0selAEZLqg7KsXh7Lz6Bb
jupvuXB0BAh7bp00UAyBdT4YQnJ7qHyPFSus4kHrreowy8YHS4APZR9YJJJI8QQo94m0tHKBciq9
DJpJjktTgmDT/XNzZnOXDgPqftcD50LuC/lfHGPWLSIfgctCVg5Ll3zRCVQCkAcNCrLaevcQUOp6
ACY/NLgz92+3HgCw/K2hX4isH4yklcenBG+0bp6C8pYY4xrhGL1x/LxLB4XZIxQdhqJqZOmyfSDG
4yk46igKkqzwjpjzv/B55BH/p5+zYVvxHeIeQjUP7SkKddDa9phSIxm8ZPlweZzSOk/nfWfVextz
mkc8Usepf/da9MxOL4BKeg+QKoVUBdQlg5C+j31Or+v+03/g5rkOvU/kFlch4BxMf+n4M7hi+awO
dGKwC+kqAJcrQ/Kr3mED/6hKyFxumz1Fo07tCRd7ppaa+rM44Rl+hF+aDBJMMbDQ94QjvJrzDQfC
5WxSvd2/hsJmSlXUVznYOjORB+B5779n1T/+fcyLtX1rCvjOdW5ipR3aIQM+jkvdOorxqqNJBYgr
ALmlH4GC7OKiJ4w+CwaH+NmQyGow0Be6DkpVkIhMrM93TVZmUxoqjNMuP95fLMMa+nyWggDJ4mqZ
m0jfskjP+DbuSL3dKplT2D+S2SNrvnjBui9nv+Sj9SRwx+d/raGe0X05n77v853Skv6oGtRSQDQY
YZ7hqbadNUDsFU0Y5zygNylvFM8YqATqWlGxRp46t1HLkHYhw4X4OmpL5uXbeRQTmWXH45hD5Vni
2lseQils04zXlwZ5zFc5PHJgqi67QtY/NEQRQ059svNF/U2Ob2kf+UGi71UUVnpD1SpGDojDQuFf
bRMERNjFw6BR1VGxUcGWFF8eDiq/O4Wn2GPU7APQRc7SLDO2Bri58rCiHYiHrulI2xBKW5NTwgS0
bt8CZmzuhCdWsn15dXTIRu2KWmPBTRUmtNMojgtDrNyORJvZnMa7ofnW/05h+b/pMHYdHFZVYfIv
TH6si0x8Gccss9AuKX0dDhaeaYz38Ztn46SMIRCBQiYMA/xuZqMbVpxe5nYnYYT9RP3jRbpTVcxT
TR7yPdMaxK1+Vsohubv2DuQE9VbQdQs95T+nuS4JmV6TFUEl168V8if+ojwYKKkCIdqgYDhQ2N/E
V7ohN960UGtu8dTzHCNxsGVqUSKEqxsfS4KYh9eYthh5jFRdqGvEtCTNSdfNCKhLRNFR6xFomCJc
a/MhQ8GSlgDGuYzt9aWTqaz4t6SK4WNSPkaVXdXg5vaHh54hmtND6yvt+KcaW8oJHzl3dWDyk2xM
fcOiwZLU1zAZfBOUC+hyx0tYZY1nF2LQPUnr1zjq2JZNQyxHsmifz6sYf8LF0ptrs2dHLLenFxbr
Q/LX7Yx5IctCyD0pJBacfUndnoEzDXagHbfSX0cH/ioKOznMAEgJVRoSDh15epDAehe66v4Rq8sf
E4sDfLRnl6M8LDDqK6ZNepcYjPgZMUOeCNSkWYLxeDOBqhMlPeCwbFWITR1c6e4oq812HnaRDeF1
ww8XLgKFGcpen/wieN3uYJmv9cQeXCKQovmIKZAv2Xk4SyyKtqoir6M1e5RhFKs7KzHCv3R4yhPk
H92Fy9scphoD6F7TBsc51AYZ3TWcSihTZrTJKMaXhmNuM6aK7wA0z8hnhyaeR2DiqvXU3qPcT6U6
k8ITVF52Tq4XbJrGvEPA5RcO/p9Qn8Jlf5G/1s6gYWX4u9yz+C5RiCwv+c82b2R1TLlvroiEzwuo
m8EVpNJ28+7lZtUXr2OO/Hs7KWyZq2PrdxN7jTgLkhDa7LyeKOlW8yu4NUv2+rbA1GEH88eGtMwi
ljz5tCWL53ChpFj3DkJAdhA9e3QR0ZaypeBbrhlueMvXlGHKE8TOCCuEKae5dBD+f3wfCaHPHdPP
GA1ELMAa5o4r3qBDd+eIGZ8nJ9beztIXN3+M+cu7WZ9aMAFJfmco+6mQ/drXwXTE0e50WjcKIfw8
hznn1ZhAFFc3PUUSgLoXp5ZE8uPgNmpQyPQixmPE7DFIi06tgvMo3mYmHXQ43GMxiYm8pAfQvHy4
fl+anCg6F8/S3xMv9Fse//47kSLUUq0QbuVnPYndB0HzgcYA+xdi+4YM9fWOEbyMxJSIwBQmTZNP
3GeHHMyJGPkVqVCens4lRx6ZA1D0lkYxkY9JssxVjNUVpgrxqjFD45+3jQHrpZTdjsQQ6dHFXrWv
GTe454oWTZpr60QKXfq9kUnb4jb+E6XhuDpoDW569fRTYBoPkIPEhTPjIM7CKF2DFbBUNrX5H6oR
aogZf77Uyisq6ZBXGwwWJwgZAjQV5ESOKXC8Jzr9Q+OcXuFIn1YiYarneQWHXwtGlCn0iIFSoLti
FDt8CNKGmVqyX4t1EZ/ZWyX+5Jq724NKJhLNL2CE3OJRgukp5Ft9EFcKYj1nxEYvNcSfKq5C6Zji
oHIlJ1AHCQMw4viExDPHwfUDwwcaCfc50I1vfFwz75rni53LrWkO0q9FooRRMa8RSg7IXCnDCRlp
c9z18cAKbVBNL+2ouJ9TcgbN0/XEiU4yRwvOh3vhr+GRevsPXf4pbOeWo/I3dTVEEZX+FZt/nHZ4
fNbaMUtvM091yYgwy67HViqo0N0pwxzhYR7BuxNKoyqdwzh6JCnjlgPR3FQ4UJ5Ihk1u8q9Q5mI+
8ol3klWhbs9MJxn4dANfvrmRiVN+LNu747+h+eoSZeH6h3gFTdeReD8ty3v80mBcRjSZbzU/8YEP
5+X/hQgnrvPuilvwcAljAgPfvQfhDpN3mw90k4SLTRKIbBVbn9cG2zhb4chQEHqHPxu1kkpLZEe3
fjYjtNDmynPLwh7wJhgoSrGYhHEYjqkSsRDLYylBABHMf8MBJ+JuZ+B8wutoWlki4VMhsG2O9u+S
oT+3HgtAVRpDgbniiMlNr7Aq91IEQJ2N4KAAW1XL69kVwrbB+SpMYsFbbBHJHaodtjvrb7IO2nST
g/+8cZ4E7G2qYl1zAr/PKhzIQtm/I8SJkhl/7Ze4aBinjaXLYUlnIM6Nm/mdjzqWrzOFQU5a8eVJ
M2/ee4+s7uTkvVuTB/l5EwUjhO50sZLxOCmD9tGvbItBQJMhM/LZQGAWtM0TT56sBOWdP8Ezn7DQ
5B4iVb2rwQrO/e9u+0eDmD6KWNEc+poyAnSBQY1FzGEH5pREizNYBvkilgrMRQ+a+4NVdNVkKYqT
K/5madvyn+rR7UkoO/smVNePN6eGJWC4YBAMduI6DtjplmwdDF0wmdEudzjBEFfcNZQBkp24anCn
RKVwkwTyJpuqusJQKMXmWetfzENTSEbECq0u2hQzNZ1URv65s99RiUiQ9UIvjQXRRKwE8xjtJ9qR
ZeVyWk3SAmUTzw0GC2TkUvg9uCVdrxbJ4DmnCutEDca7X2qaOZhr70FoVkP/gu1ogfTM2oyLfrI7
A2aF8gjH0EcZL2H+ShiY8WqJPLA9I/hCmym4o8M6960BIUxOkhmw4uFi+bTWBfo9kHxgTyxoS6/1
KyZH897gPOfWLC+Jd3vS1UZfeXaDyatvpMdARJDJJGOZBWyKaiqot4xH2sVyAzHzFDhqOze6iRmN
tZRsiv/nPAqOYi9bCRDxF5NxsW7JpiF84YaBdqN7hP5Z4ez7EqjQvrwTbNZcqyPcKT1IpNFFUFG1
Kn0YPIjotLDlBPRHWToUhukvPfWDnY5giG90OqStOw1EvTfvTbx8tttre9Co3AvuufBZP/hjYVhh
+Ga/FHmb4eisa45jkUhkqJ84/3bapqcgoDK94UDbX+lytRTOLcoSZiDJnbxVu3dJWLeBsdZc9g+U
tY7y2WbACTSZsw0QLFYHVaUwu4JYnvdfLqbq3pqbiP8TRzMwk1IKUGZdnVFiiwbhjY5VxNsVAPzB
gpf2jcLE1CParxKp6Fj1OPKhSFqMtvh94FR0Iszr9U9mEHXJMuWRyP6wNwsKxn1tI2xZLwSCeO7Q
opZfL6NQNdrs9CpVGf10Lx4uXSBDe8Q3HHiBT9lRa7X4958fkqSWqjeGGQ/HFivKAs/jF+LCvkq5
MPhJeuOjq4eXCpe4/3NuTXPslvu5dEtiSvypQQClXDRxy3P2QAiAmBoOkbrW8wsoSebz8gmnUHwt
ekezG0mRTUBiGoQLfnJgBgQSClkt96ynZSBG1puZXL0h2KLTnFji5uQ1ZyhwPnJ1kHWku1OjEiin
uSnppan4byYwMZ3KMHQjl2lxvhcYwyAf7UQeUoza5l9K7vtZ74n4aNd0LobQcOavBPsXv7VDDRyU
UwaZxN57aiq4MK6c8+aSxmiyKDqNFpWQmi7ZtryMHcWoFG1w+67G+SKzbmKybzQsUxpv+fpYAmrw
43OQn80sXwEaRn7wCQImBIrmt3LQoupVFegZxylYPnsfs+bGjip8eSZA0xXhtr4fvN5usrH27yry
hmG8cMmJJb0M7yFPa28sNciG2XSWgVzF9RPOjoRr+tgG7zj4qXKRvguqCtFIukFvYnl0jCTidDGp
J4Evpc456K9StBHetORfHiYnA/e75XN/yaVaHjAUAh5IdBxNZ/xusljvIgFje9Fsg3aOQiZAHvaq
msGOVKUb5607gI8toD0zoVM9ijqYZ2BW/xMyiP5y/hMnvCWvwoQGq2E3snnWxZTTkBIFuIDcDeX+
lKlnupk6IqSstP9QCY3WG0NHveLuvAagUHLmJwQoFQvx65eU7alFw2MpTZugcBZkx90cj7PpBScP
Z48OcZ6JIvKTzomR4CGxzgi/Igoh1AoehndH2WKCJrvz3rTMNxX2Lyh8xWqB29h9k7SbDek/Q6K3
9XSjJswkTTsJwlNSNMEfZC78hkDt58t3RoqdJoGdsgM9Rjl4vIz6dH2XAJyeKQILx6vqpW3RvOLf
BIb6p9WQFzH9N2BC+YbnCYEqC4tzOLadpvtHRtRwprZiYNuZ99OYxT3pYkztJND2/eIGbhbTiinr
ZUw5ppe/CZV5F1c0bG87HMvNtQc1V5W3MYSno+9nGXnWf9zhbx2gXQ+PxGNELmYANlpvzPkW0Y7R
ASfSydANdTqaPKhspAIeIQ41Ef7nePrsMrfI8nqX4wOY+wTNokGGGNKWwD2c+xAv8kaqAxW4vbiR
2iuJhMsw/yvhodM/Cb/MorcDckbAONIB6+Suc9IyG7qgum+MWWWhvVoadGI0c2ZDIBWSzCU1fAsT
5gCRsmMmuqQJ9kfEVIaYF2UHLv+4vQKMP+hZQdtgbHTvmFu+Ks3vNudruabjVeg0b2O1+VQpDfzo
udnkGFbNv8FXpKs0FA1mJispi4CsXyC+QC2CBCYjTm0gVRYQOaG16VEx7NP1fyhPIPvLQHxgJKz2
pZE2A5mnIP1CTdGGy82GL7/RhuuVpE7fyJhsVPOK0TN2hhvQ+cZebmzWy0Wz9HmzExmQHDVAqpIh
XBA9Syl+rqKu7iE+wQqWWkOtk+xlvC1oRrs2XcdbMzN2festZOCPk9yzhbaexXav4gRTL3aOc0jo
1EKiiZU/TlMMuK0BQwVUUfeMBbcBoc/3aRw12EhhjZgaYhE7MwnLZw2o+vO+gLD1VBIF4ljSNo4q
hh62Hg4HkkNBHv6x5sTsdQu2EMmvi8p+QT5ICv9GoXvOykZtLr0leWW1u+PHmqJ2sXLJkfEixkfj
9/SSVcSJdJgdUXct5EExx6uqJwdYXV9QgO6o5w4IORQGNvGPlwtySobTjTsBKhCrinzzo6N2njkz
jGZe/Sm1Yxh3o96btuWBpw2vPslePHH/lC1DdOxFr0y4GhTBhG9iQRFZ1GX4UEHR9B8hyc85JM62
rHYjL3mQAhLGXBXtSApNDu41AE0Qs6AmD/Wzo5cIEet7glVT0UeCWh89DZTMwthMMjkcNJ2Hdw4X
TCZIg+Q4SDLtLuRHGKZ0xxXXBWAvrllpyilFI6RhjtkxnGHSPTmzY5QO753v+SaFTBViN3oVZJty
kzQJWw3F+kJ5X1BBjNohExxhUWw2ROSkB64FX/9HIF0Vn1AiNP6MUih58F42H4OXe53T273ilZAP
EzyOR9gJWDXPsWc3TaBQDdY5tYbA/p7bjoC2EuMBLmyc+VDavTg2LGMaj/TqS7UX6AxX0jljM/FJ
TJLAywIsN6LRVGYb+pxeN3Jy56qTKTrc3ySTJMEU82tsqNb16ysoTiMjXDoELPF9dH4x3df0VzGf
1n2LSMsRwroWc9yablQVzeLZRppWeOoP5as3nj8mchpsYh1sPykl6Q6kbkjHszUW3pH9KaBy3+s0
qewjoqFRO7QA3rMoUcdgAt8RIzEKRRAXQxcHT0U/PFCdA2o/1jRiTE+s1S0OogTMNMGaPQfgd2Kr
cv/nLXWLsa6GwLF0czrDDGSuh/GFpz4jXtzvrYay8AezjqXrdDnHD8v+OIJ7XDqjd3IFMfYoYcDq
va4ujtYRItjs0Do+lA0j6NUlqD1tAcWRe7A3RFzlMyX6oxUCv2QopW7L+l1kQ1vZDmAjSDYrfGjT
/sMq4y4Ol0A1xRdMqeONxReAzNLUe/T0jRaOc6LfYKLrNOvtF5G9g0T5fEc7UjYYQCm+XXPoX28G
QxPFuCqhbbyTUHwV3tr49njtUAtHmef0MXCsUgqN6E2/zkwncNgaOUjdCxm+j+vll/QmXK7gDisF
By9C/Qdh35RzhcqdWfIOQTbRS+janhvHVJXIJImtEV0bHEZVoDbXxdGA0Xo0IlaGylIpTVr2odlV
hIxe9J+tTy/9f4TJAYf/k5nWk4AvksRzSyvVZnV6JHNJketmuhAiYg9PZMyr17jX0pWyl3E5WeBi
4ZS8Qaxri63o3Pya36Wq1+a+ULC9vxa8DMr+j+kTQdfmaejZaX2RSjo4ocmLGv6+yigK/anbB127
N962r8BGMkODXbH3TQs40J59ivqoqeQ4xsOMDfkRL7EFZdYdeKfYGwDIhzSysk4b/Cy0FMf7xhq0
un5AKoCRTZVVR0R0e6dIkol9AZ/eNVlrI6gDHw81d1ytGvyTD0lYBcbYWfnmtWIKLaEJ7Jz3QvRC
defCclFORpO0KVtabrN+7kwuYfT1oRVqYb/T+TgB4PtCXl2UCeB2sXogSO1nj5/6VqVrFyJdB+IS
Rgygxgo4fY2HpSYNfXvhNHXBqzHLniecrgw+Ze7ovxH3aDgbN5KJNy6v/WQnn+z0mPTcJ8xBTZ2T
DqlG6obhnXHPc1zYZnAGSH9QXmOyOsJAiu+XOA8bdifNNgIkdt1YmnuKoq0O0Hz/Pt6owMpS9JgV
ZcYwpZesH1+U6cFm0bkQoCih4lYBDZ3XpmYBm/XTc0TA2VXggHuJppzntBQ3P+x0eJzpzDGvbBVa
HzCtYgToceJOpd8Ll721h/z0+YSd2I8x1vNbz5poK4ODVdHu69eyEdb2aPTRbSM8VFzJNJ56sJGl
zCJtCrTjaZzUkDH3QoW93ltLKDX81SaMCOCGC1gWDpQzD9laz94J5zansMDCTCUnP3O4MnRqFobQ
FQp36RoJslHXFTTVUp8dGMLpG7Q1xrET14Tys88D9VObKhCdzUr8RRuIwgIZIsVOnIXc3h/27AI1
Ql/qP4MbtJLmqZibcbIMKQ2V9Smex5QWN3q+x5U9UdBdgN4+km7/sWSoXNsMrYs/l681hdAtjx0K
1aQJBYpFhy1KQ5OYbnZpIv9Pwrrh9JBXi/jLDvXOtj3S4hs/gPRD5zfDhLT9MqhGVn+/X89LLTcu
D+HCHfzeiz2P0SBGwKKY9Q8yPsmL5vhwAkte4uMAaF1kwIKfPVSdoUVQkYkuVVc6nwAZaYcSce16
08TBWL2nXyfFcWmkAYuVrfzjkqXtCf7VwepfnXEu6eGhyyA3OyQDYYmhyXfPBvE/rtcxntCMvLbN
aJVR++r1SE2mVlkENkDMwGIj86veA59uXprFlaBKa8Cxc9GYhu/RyEAon2hbmLQtmFRyevbwSp7X
Eh8BGJ9NQ7sPGwdqJnN5SQyrzJJERSsW2Hect21tPIVqTWZdkrHndEltmopUYTGXmc2OL371n15q
Hh2uVZGrGxXA3YMOiDlcMKAoCWihNZvFdVC9Qm8TAzZZ8CBlqn+12buL0ERJwRjMxGarx1T/mVFN
Da8CxkgZ9N5iOw1AexBW3X4gQDsYtsQuxz3sAnCHRnBS9b+NovNbX0bpXrZuzEu6SFI8YKE9lxv8
qboDxYBsh8VYHecA2SpmNHQgut+nGTHukPtysISzS5GGeGg19QAAXjnSjwnd7yAJYPGl9JxrHgNB
QHM6jbCNPSk6jiO4jC/sOeSL9KE/V+AclnHrDCs7dd5plAK6DZ2Ylr81EylZD5dwAJYY1vOocZrd
pzAMgXKqz9fO7xH2AoU0uo6a0tLkpD0gQvdG2ctIRci4HKA+NThpVcv7qBmOdPK/XqX7LOcYqulB
ctxjEPdRydGlFpXWJzs3yxa344AwBd/cmMdQ0tsm6nERxWF/66IOeq2ISDEkdfvA1PQjpkW+16yc
1l0PE/zjLhg5j7RjlBaBEWdkGEU+K/oQ83Uuq/tv4NOHKk+XUK3Gw2tJtrI2fJYiPuxFZ6SY6dAh
2DjeHWUPpOibupsWDApoPdbWDVmXz5GVTOZGuHAYwEFosMNjq6/1IhyE06HlwwqaxRjHW80Hr3Ej
ylFVAmqoWEzYERu8e7G5olGLhrqfCKM8ulhALgPZyZEblVknrpCX0asutObmBeHWaYVi/IVhd+G5
HIzF6YK5EfuRtFV8zLcpxg7dA0VMErzT1Y4HRxNkgtdDoynNIB+3CtlqP/zr+SUdOedGAtzESn01
kuX9b664lde8QEhd/VtY0OI8vGfC6NSgSpwHz8La/W+4j1G1ujtXC6lUUPtqfkBv23/gJbZFpN+Q
SGyaa1eP8XWvDO6Kvuda8RyQw+CXbHWyaTHYBAM9bRMmG9eUqTGxxgPoA9P8HLvlsCaj0lP1q9ov
Jlimm8AIcgDnv4QYtJwGR+CZaObSI1X6hJOlD1YiCJ4X96ktDVM2ZAi8iefWTa+zid2goue8tRQd
qbaV+ZlMYtVa+hzUvl1+8u0fkWcSmoKLhg2JCDL1aK+3OTIQBLMNes5rQzSGw+IXEN6KI5lcpV12
thJ22oJOJ+XAHfgWYWeLB782CnTKywu7UX6ojzmcGfwyNj5AwvRLff4DlVLkwp6AnqsY1LXed0PA
y1kKxtYQTw6pb3iTVYBcTrq0JHVH/en+UkcjIy66oHNOnKIVBEZnpAEZgu+tzJZeHohYV8qFF8P5
W33/htGQBCKgjFsnstx5S25VZVoj+sc0QhraEedmMNu3vwgWXAyTlpvB+bnzLBb1kUqAIwePc9Ja
uAGxr1mcpa1apyVkc53uEKvA1O1qFwkKl2UKdd67o1CT7TcE4is3COTknY39KuL8uZqUJ73HqeBJ
+cdfV5ecLXpcbgvgq6AJQGuv2/Ja6GfYMraZy+lTH6N2eXTVGlAfYh862KHQE/Ss2sT79QOU0kbz
fCohGXRm5FebG/Ms+Yq1tgWUH06l24NktzSHNfKAMKieGHUyhRnewvlqn2HkLKo79tHXarevxmeh
5NJRLDAgjCXKh5QgugAYL5/m727NQBUuyXPViyma6vGy9VtdOl5XEJ8zCZENvCfjy9bOLorLABQR
S3MZNa2Az91gRFx1QkCtX1kRf6u4nsuq/CXmRnAdTYN7NWjWr61GWY17EN4YWFswDqOaHfR8NVh5
QeNCoXBpBP/6JBns0Sdm2l7xPwrNfOZ1bVjJwtwgWxee6hm+u2qXmTYecXasCNCOxleLyS3EtbJq
ZwFRat5lSFPltoO3QkNcgrk/YOvEaTcjeUCCFSzYONThUjE6m/ZgqmoLeeylL+KlZ69ysxE8u9G4
V0t/60U7BxjVwpEXc0+AmA7WdDozqp7E4D8C/cMMefmJZPjvu4We9iuLSxf48L8rD7XZlIhVAnVh
OleLkiEnFl5IWYl6cVb5DOlYVH+zSzBUplhob4z5OFF0bIVGRufJfuwYeFX2lbi8qmt3jNRMM/57
/+lxk5MShzCE8i5QBD7XssVHPMXYo64La92x1QaUD3tNFSHsU8TArKqtd0bqBXe7PytX0fU1BH+K
cYHczrkvysmM1O0eVFxDjDfZamUxd5YbHP8CwPg7NTKQv56XYKjgp9XVbr5mnESAcj7aJhvArRwr
L0uK1ZHE1nKTRsHDtK5xcLzhmjCq3hfJ3Mm4KsaaFJv3wlWq0d482ATWUV5GRfzCEybuP+pOqmvw
8Efd7nS6hjKieyeo2v/xjh7zeANPwvoINSMkLlQKwaaVFXYRKkDXmtYv+JlDFOU2c6fGBvMm0H7i
2M7Hz8Yj/YHYzViJCeWmvxILJCNTAGVFiaxcFap5rgA81O6YxOpkW0BoxwDkodzc9HDzmn5Pa2Jj
xgfNb5yZPzegNiZobeRU1wGuwo+LC8Ul4aa2HcwZW4ZFgFafcYsJHfydIB9iovbSjts/LvSa8vVG
k+RBEcuMohbDRcMHOpVkh4eKsiHZCA3pp5StP0yhf57kZEIIZPdKd4oySwynUGzdpNcuM4gKTFx7
qO5jSNddLEU9FRlLHtO3uL7qzWGs0GWyRXKLbZ0GuGG6uyhVgPgAb8MGIcrGrDxHahgFmn4Ep6zb
hJNGf6DE5noyAjM2XZPnuKb4thYTlLWklPjj435rTTUThP42sFwAbS+TKiVsw92BLa0iUTHYpunr
qCsRdpFhQTMWwEbIzoYt0SeyAj3bFDwMDTbvX9v/YAhdgEPhtXIdmFVY6zo/cwtdhX20dPi0RB74
SVYkUw5lKid3+FT5sNgi0ptNRsF1GhWqRmATEvUjLi+f0cQVzytYfFGOCBxRw5uyBnFEX6ySb8As
crldkXAxSJL0FK3oLDSR9ii5iDZ91yJ4YF92pOM2fcP2hwHGivqxynNj7rXEmmmjRYtUwCAMHf/f
UDDOHTJ58IzG2jbPGjaH3kXwKEbzQFrMwcZuJLB+mLV061kxEz3l/OxJuypBkPjJalIkrSPQdKUf
3MLx0/y655FQzDoub8YOyWX4lpZlkxwb+440D1mH1xHae4KI8E0z60gbssZHNCH4t3GB6x8nDFnp
8ziAYfzlDwCWQ2OwLbUfozliJAzvgsbfL2tkt8ijNELkXWKoXES7czh/QcwXqK3fOpkomDKr7IHz
BKrSNTzLFeBhzRQ4O306FFQ54mQwIG89DjIrfVlhbVQCbYKVqdf4WAxsgLEk7g+gOlyu9wwbFaFZ
ow0xmoIpWPSHtqY8CPWOkAQP1NK/m+XlfhQqK735jZEypFHQcNRhpLO9mMky7WhhhJwn9L0BJHna
tZMmODNqZaVrNi5iUm/vhxgAqWzW1Due4w40jm/Q4dSkn47DtsqMGcHY3t8MvNF2gD79BtsfwlgY
D58mAM9hFZQ2gGZfAVIXjnAUJogr/8BO2TNHJMBbE8akopZuPIM59VD9giauAANMZFjBAQR6tLTP
eOJFN0nOrNfS8xuGh8c4b31cgvoPb87aQIZSjRLHQAgu4VF0Igwfzp+N7bDk6iZemrzUJ9BrSIVd
MGNVAX+NerKbfmEteYC8YS+9gdTARXjt9io3ed8watS6BK/UIKwQ1kAe2k66RTc/HJZztnBhW4FJ
gYbQDTJhpf0uZyplabqTwbh9XwzhyqZeVdTK3yYO+im0cnIHIyioqTg+0xTxbq2+4WRdVmcBAp+h
x8JhdbF5OtA30NLzrnejFDbyUjkq/SfLcawis9jerB1eH7rYLhrIHA9jOq60w596UXUiVroetWr3
YskUvKaA4ifBXFMcqDbQTvoimwDiCdK13w2Pwcnt7kdPTx0+bHzEkr68EaM+2nxUITFuRS5u4TJM
DuY2eHV3dBJ6vuZmzzJDMqRV10TLL8WVb1zG52tzDT5t/a6b0KCdRxd+PoiQ9xR0TOtXzIQcrmwr
zbSX0a2UoO5p9pH2gDC0uALhUzBq7At8xbeUj4/YrRVyT9SeBmVd3DguKSQEJA21FlC3TO8guXVA
480PYuFqN9Cu0EP42jS+tNy+WiZDHWOvTLqtc4cEjWEJ83xdugcMGcQEjI6aPtul7Oe2OQOM0YjV
EmNtWWXS1jrntFyGC65aYFIOS7R3KawOPPt5pg2q4wDr2+PDyReWPfA8JZv+Y30si4/j+WnewTG+
r/HNEHjrEK6M2h+Z9dzPfj3gqLI2r54aY+3xLc9wWSQYFJoLEV0WiazQgBbtyIPms6vu2JPq6AD5
pJL3z5hLk59iFQ5OBm6ctyEsVvhWhd8GmbiAZMwgpylXy/cRZSExwACWTBK5LzibpEgQQx02BD/e
Hm9bjN42PLXOBvOMSk7xbv9iQfyt9h6Uk4VLaDXze4SRe3eSZ9iVTmi9bnD4smsQpv4dPxA2GFdi
Pu1+hHiJR/ZCw8TJBwCH/Bl8fabrpWEHdqQMUqcvVxwUxtGmSL1aZBhINCGQqZHGBOdWz3QDl9ZR
2j5YIb/fvFhTu5dHOSpDY6WExrNy7Tu+D2fONO/S9LgDOzud49J0GfhcvtfhtDsN55MJ++nEfkvn
Ds4ltcwYQc2bYmYDaX7QKnLi2MnTrywIEdr9Nwa9WkrJbKyBCMNESGr9S67L7WFlIgxJDgJV8FY/
cbcaCbk4jkpFUkik7CnN+oSoxRc7C7cQD3qGzWIBe6SE67VrPnA9YdeLzYh1auM5tJe6khk0oCqW
mNam/qTn87Gz21sE3RHTCU2OXLZbBXH0TsPTDBcd4SasLq0HAqqyvk80IEDT+tO0ZYOtRlSkuEVJ
RHzK9TesLUsydmR38p/1phzD7aOqoQsajsei7SqVzArHK9WUT5KrKnybIMNnIbyFqHIK3ly4RKD3
qZzDWrzoF2yAcRZ7azZqJGb1NLRY53u3Z4ByFAx6hxkMq7or6Fe6kgk/xw2VWuwJFX6zAb2o86vB
6IS2Zk/eNF2apO92eOE0tx9Boo7fmYx/c8Ise/8J/WKgmqnZcv75DquzODCsDPC5kJOz2CPYHW8v
a6sPIrFQZ4Wm1j8d78rJf7tk9SF8y1xlg0J/dCP9SrZE8d05cSxyDcUm6I7iMlt51JgiKaz+joa5
PIkhFTywYIck8zEqr77TJRtO3QyU1QTjl6LfhOEJCRkFj2/txRIU883dH8HjtPURGxgxT/cBiVXd
Yjd8d3RHjhCFlLiB7V4d8Pn6kjuBI9rLl6hHqtJ2Issckrg6KjVYBwHPIMODrxnwLlnLbwNjv+MY
mCfUsI0Tr4A4APw1o1xP8RipvK62i+zkitdJvw5KMJjklqpmYpH+jCU7kEOOnKuJhyfV6R3YFJr0
20YdK3LKlwezGeZTFkkye8cEy8qTRIk20jn7zq/VT+Zw0Bmr+q5Rzk1gE57VOGr6LNN9oXn7buMR
g4hzPVppM/zDQhUIn+KJqxZKJHog03aRMYH/PziMlK012VVBxw4Og5rDWf4qunNKx9CpI8MuS6M0
H5pvWf6pPGmjR7Jsf68Y/Y5m/Ow1BIOP8qBkXM6XqJZHdiQ7T18dJyh5KCZOsSKZl/pBzHQxM891
sUdPCpyXVBAQb5hM2pme3EOkv0jm4/3uUR0nKVUnCIKhp2fRBpEodWXc8VSi2o2+I2xtpvzIT+qD
GdThSEtpqe7Y1tiTeoCtM5fCGTo6cyoWdpq7dOj1mYkdQd3Fv2MLZVZqKh8GCn2FbAWi9HI1rwYg
iSeY5SFJO88xTOFLeQPlrqB4yO8MQMbsEhY/Rh+M8hq9mt9WI5wqSE2XG+kZTKKIJuSewVqHYTug
8T+OPdTzHK0L4bLW7xNRXK7f7u5hxk0g3GWndhoUIex42Si9Vt2Kjkj9oqy32BE82JRd8AHlvDnC
fGwdc//mflG4SbCfzsXHJUeFP/hzZc4Vri1JfTs2gM9znDDbfsAaXBn8k8ND1CoIdmQZpTfAMSkf
saNJzvGbIroMLLZVA872sq5H1+ZsytlGWHzwgpe8jzXoneCvvRYclo6mkfXDI7GHlprrPrBaBxSX
y+eIQN/jDkC+wxS9FUJeeKhS5DyYE9QAoWuejfMUsq4z4vCrmf1G+5/qK3v7wm2rx+sVj7wW13al
nnlvURuSHbVGOOFMKWnE2G4d6tS9XXegsBCuYkV8OanEYfcYuvLjE/k3UbNbH0Fo5831+ZaKL29j
YWhnuXIfnq0HHKY3YGDj5fwRs2KMrsGUHIqks43IRJWMiCoaXBn9i9Tr2ZHL4SLVPd8rdKDvbst+
/XtE2a2N8sxuDUFM6aooI/hwjIUdl5qJPl6GKmBe0BXpe9jMyCmN66EmpF2KIK3RRYm8mDTFnhXb
eQSBidQ9OZFxGJTbFUv/g7yhcX+UrHQ54QUyQwj2jtZzYa1Tr4Cp0HHpO9tyKNsiOEJL0s5L/dti
HLunQIC9UVqU8TJZOxtFSGLdQ8WcEUZ3Mq2yEYmWp/2JrkRGAwkX3Z4K3MuuYJ6vhdle/bZGOziz
PT7x8aTcNrGrP+0MV2W93fyFh44983xnxC4qNOMeZnY5q92yCTyPKE9ZOv4ckNbWPayjzuQ2PEMU
7OqHsmfvMVz2A/ROkzTAbAmNXmkubho9gZ17renr/6Wckz7EQx/CU3Nxg6MRP5VCZnQRlxCfmX4p
NKfM4Q05J+/afsDvue6qFBLFyAvyHMsPG4XBGahQmTCywEgCj2KvjXjeJdH5iV5EN8EDdIsJN3sw
TtaJARvmjhm+ejQXkuX9tplAXzqpgJxXdGZG+xbAhW9MIQeYMKprlExLtVeTartI3LjtMzTG3O6r
aeY+OM1iHsuwk4YZ6/0z8+tNhGYougEyALv0EwedobiwwMkeMuUMcbxPg5IiUz6y4dNxGFoLrwQu
VixQd94A6+1rtQzzBeKwhDsz0blpOzBp3LgUkQBexXTac1AnSBwKIP2dPGQoBb8R7FD7lI6FtgGI
gfQRtLozEe0w1G3ZrO8iTJoXphj+oNrqi5WfZJH5arNBPgUCjMUTuIOqSgD3WfEGbTFi3yQ3H5Hd
gACh9LAA/Q35xF8IauXRFoM70P3j/rvD35tzSZprHAFNecZYKGNbxS8TjBt5w+fumtsANYmP8B5V
ddQJDWy6GesLft7sc2or1d5Ub5Dv1wgnv9/8fC2eUCCBpa7AZorDoQc8yI8k3aJHUkisgK4D3VRM
DH5eRbd/RqhPnoYqeQ9dRj+4rWdbZf+unVHLrvtAzoUITDfjcih0xISaIpzUs16xW34DtBZ4OEiZ
lb9D9ZkpLjHT+Zar4ibBUeTtAPMzWEfQjzzCsxFdrIERnfYFwLTapy6qChMqE13FcKHvvOkgKHfe
/wLdezyJhv4f+d/Ukk30RXqQIqxngfiykzsMOndJvdt5L7Im8OdxaPFFH/JcoloR1IHejPLxPzVB
cUA605vELrDVMgOgnOQDUuudPY7eLUdFwtt+lMospF//jFtObMA7v0i6JBrMhzabPNgOdju5i2Xy
RFVmQaD/++63RpQMvbUXYXnEeQmpH3fMSHMrx6gLmb6gWF/dSr1kSmB7z0lA/n2YBj7RrM1fHGzw
lDLMBurhUZ1Heiw/PKUmi3I9D9XiT/I+yua4siqMHQNseQptySsUnAKXSq6+vWjEQ6YOZSjrWtpS
Um4uY/TytrZlSnoQuAX3TW9dH4if2m39Q8ZNqDwRsnxtL86wrVi1a3WzEXnzS/R4sPwicgFdVBOL
A8pUYJTf5VL1L4r2eS6+lx6o0of6/m4+csLwyFiSchU0rM9kX6dsze6CI3edO2bOwP55x7oIrQeN
VXIC/hGjDagCbxpavWQvWd3ra8TRLnpQXpz0tks2UVXRxRG5Keshnn5YDLsFseE4J1znG4J1ggpn
uGKYE1ACvgVb5GciOZjMBR0Tbq2TDm5RYAv8lYiFLXG9iBjZUnp5RAgkcORKY9owhI7KCw3tUO80
duCWmfU9+EsxoYyI6L3T9H9JV72V3AqmWQvllACkkD+5Uw3SGo4FZ4qJUIsSwEllZY5cbT6lAh0G
PdoMlnKKQeLbgk01BmPEee4pHg5E2wK26Gzj3QWBfoFWwDpBkVDc7xUs6z68Sw6avEBE2Pma3Quh
8oR6p/4u4bqCmf0ICP5AXDt9rA45JxgQ9Ei9+yFmXENqW+TxekB04xehYZwfKvKYwkdthc/yAM5u
hntN8Ueu+W2h7mOXs/1Gq9ISOPcsG16k1BQTytpNFff+anfE+TcxD0ML9BZ+QsANq32LlX0N/4W/
VmJO+5s/sNEWfO8T7u/MFJiWRO0uic+9629UP/egB0nWXys3b/Xhua8SEY1BDVuMV1JJdW3xZWWz
g3SzxksITgfcKcqPi3W5JofFkVmPjjildD8wGxpWz720YewjHGppCqJLeW+48SdF8IWTEnR7K+WR
Z6oAyopsjj4jfhj/Kd6Zq/+T2xSEXAgmOB86xrqcaA5jhkqfTWLEp0YGo5aEJewoYjDHuW5268Fl
1P34bHXW/Q170EFzlZ8UXLFo7egFifxVokTNh3PBbYvHRZVJJzctXI3AAy7hrUjPjvRc4Y9VWxc9
aaTQN9cbaudiIk7C/nWGO34BOsTCkf2hn1mkd60fd0FW2mEI8AL6iMiCwdtuHMkRsaXzCMQUBPhD
dp6xGJ4iy0Pn+uw8CUJdSiQM5YU5w2+FcxCydHSLVPqjVT3WdU0JctrMEAdighUYX/S2Bq3WHxq8
mmL6a0yPum4fbI66PMFI9JoqXS6jQuGtu/l/b/ZMnACYcsb63HCVuiuRiNBCQYo/U99opkSaUbJk
Qh1fRUcYu59gvFxQ/b+/v+zvJLdUSv5RJIa6HKSX4E7LzHyuQ2ZkDYMSKBu3tF5EaAQM5FA6li7T
ZkocmyCDdjqC0MiA6VXy1vmA5fvSAvVJ6K5jDH99qKYz0czRCxkLz6VxM09veJFRInI3k6ypiyQY
Emxi+pP77leh3A/XHwQY48ryByoQWkzrLfH+eYvYW9aV7FPZOSGJHD+vlL5QwHy67HMgl6QtYFi2
jrqeVbJbrBBn3H4RM4/YIArUJ9cRRDzUYIzGAq9uC85uPhMsKMzBga+f2/b2as2t9jBinc5OWqXa
2fIe1LkujOJGazue3dsvVBoJc7Xe6tJh/lEBcx2woPMvpFuYtwU8x1vRBjw8oaHzrfNn2OsxA8yb
GjgAJv6bKJz/RwKvT1aR2fYKxvq4ZkaP70Yh6i2MIkLzDlgv1FF6TQPUMDw8P4qUzwRTFCkYwPIP
Pb0zH44tJfWA8JpQbzFJct7GuVQN3Cr71F/s+NLSH5y1xg2MfSDTCYFn2b0CeYZl3ltb25c/MkUH
4Xozm663PSjeQH1HoG11XnwtX5KmL1VZevWbryXCfWYTyoPUaeDyOJBpTEgXQm92NKi5gyqDsYNz
pvmd8JuLy6Vut+oI7wZOV0OplZgrWitYdllSt4R0qxXDz4WIAYLVy7K8sbK+qTlCP1JqKIbYRg6L
7giomq+f1WewNvCrq05HzE4W0A6wjAiNoAYRAvlpAZLVQxT3Ct54lNOsoN6pVAYb8qw6fnJ5Ni84
6W/tVGyLJ8JS2+iJYD7xqhijUdFXQb2lzDDxAq7yto4P2rl8PiwsWe73aksfI2eIt6hA2Gr4Phw6
x1/PHOInK4BddY8e/YWSAUkY15z81VhvngsvPymOsc8lB/iONKIue6bhKe7sZQmVPkBQn4Qpr7oh
8LebH1/YcRj0fp1+cJdtJ+lm3ZZR+3RPT4uyewblIOHP4a/i0O6TqB/PqH5SQYD0N3feyo2zfkE2
Dd6t73Mx7KHJTRVQbX25IBMZN4Xx6hnnPzGAWRR3WXTSyc7MqAKhcFMSogKfjNIAgabUQQnsPvWL
pNqe77Duzlb94YqM7S8mPOgl1436WeLl3W3jbxvrTF/MvQ5G6orFKgqOAykEwr1v4+uLUW2VrBMl
vbG3eBr8A20BifGlvP9qC5+nMooiOTDclrHwAWgMuhBGI+KPQ71sqgnIx9H1/AxKmJK+BHUUnVkY
3JhJ+j4lJPoZPR8a4lqOh3kgSTXEdK9y6uTEVsmVgysmHnpvF6vB3d5QpGjxkAHsEyafBW5xtXD8
/VqKz4dimgzyXv2UWbpZF5910XZaB0Li7sWqf4RavotI4HHunLzbh2fQZDvqCjrAalY0QBvnbcoj
695Y8m2uXVVfQVu2omLTavJWCPfMvBHFT1dGzimVXoZYJ/bPSOZp8aunD52RwPOmAEz3Xc8HRk/h
MFfojFhD4mgu+Fyg5Jg26Yp+rUcitxr7dTnMdYEzFuCd1ZISAGSVunmH1itncNmwfDIWTa2XmYev
KE0mQqKW1UNsfYtCJukIGmDldPM+p/OwWyn2fd4Sjp9pQix8IQ9oBELWXyWFL1NAuahvT0iKxzzZ
Gl2r1SsB/N9kzxmC2a9cs8nlRP9PQVrPNckxZE3HjuAWd+VI72n4IW0DM0xM1Nd0kWBdwsEMjCct
xOjRtLf35otCWmeH3Jn10MF7TMRw2UsZbiZx13ZVEL4ncmOjUV5fxHeTVnluM8cxO31A6OK/CyH9
osDlfurWfqwyIf3FTr05xyFrbxFYFvT97ulZdPmTKSDuWQZzAPJYl8J6y83p8Obgpqp5LldJmzYt
LK5O6ZOX8IqxYZvEUc3j3iK/eJrNhdcsau134qpqqCu6UlVOU8o8vmk6FmSndlNap+RqFpWBPutt
kPd3YAMnxaJ4wMpMHA3RW9pdo4I6ZlEg9I7ekCx0WOEVaKNtJzKKVEz52hnFqti0mfVyZZ0yJXBv
rd0aP0K/VQHny0LwkMieGT4zvcrHfAUP2eP3YK6PC8jvI/GhSesPmpezaF5Y1+SveryUdhzCzSrI
K8dzURUuDALQhe+W94jCnzXRZMw6gv2mP7BQDG0oKfc9NAsGaKKDKReJMM+Pccz0eHjASC0NkBKq
6JaHRHC1g2eTjqik9fVVwgrmwE5yB4KM01T1u8VI7xL7FcCfzJ/e62d23WSynfSPs0r7N3PxLisl
hIWN2HblX2Jo7GYIdOuZiBzlkJZSMOs0QUxlJAy0p5pd41SBHDd8th3Za6VuGhrMzSI7QD8spKvP
Q24Qb536gG+vbfggi+FlndMzFX+ddFaiqibKjoFFiEroI8mx0m8UeUYqE33bZgrkW/kiFofrRqQS
A9+lqhGQg70gS01ygY8F5L5JRYFH8qqCgh3y2GthH5PnZ01+4Z3P7mZU1I7iu9B5kszgoZUe6r1t
6RIzI6gqZeTBBHyp+u+fZUJmWbT5HkK2rCsa1BHz0xwSxNDSfMGV724zlbiF8mfj0F6Lmmq2Cc4Q
q1mVh/nLzD1tnFpcqd9EMHiHU5AloItPSASXGZonXMQfiT95QHSghkA1cYZ6TNriXTvY9yaHviRF
nm8R64q2veewfjQxSDX5dIATvrLrozfuR4JeShDmJ7G5axezuaBGrR+3zsnJPiUJg1zq7zauCrYK
wXc0NS5vhX16wLd6RfgkgUUMcepNjK8Lc0bHUQFBKQ8ZTd3hJ6yPg35yagKDYZIYi53rbrmqnS56
lgCyzdrlcM89qZolBOPuKUJY6gt/T6uC5JM8lRY7e+N2rgXLF1mS1bnBr4obXmEt33gpzmFEn0Ij
st4vdQq9FV9juvcnO3S4d5eW2/tQp9tYlZI/rwo1tes09qUoQAv6faQhdvESw+DGFnZLzw3/H4pE
DkQGBiA4aKIPZ3zgA/O2tLD06CKrwie5NTxB+GQLBUqX9efYKKvy25wnnyjlhbf1mqth7EbGT0ct
RG78IQOzDb5jLqpO267UvHypz/497UNbBVFcFEoo8f50L3mY/pcYblqjqqBVHoTuixrIw0mFh7Ow
UNJf3writD4vGpnfpj2u0tNck1S6raZ0vf/8wnkD3DeT/5LWgUjyfzk6GJnMTJd35ICV6mdWXdZL
Wskhc0FG71B3uTRl4+Oz2Kaw1TUv6l1UWgW/9lGEYl51/IKJZCb12AoeEan5lt0MCEezEIMFK861
ZlGmQTN07ubBMp7NIBBMOePibWwyx4xVudLlrX+MRvMMyjCiINEh4xS50PmIafwr/sdTWya7Gug4
O+g6npxpyH0RibJZGhVvItzRWxz30qNBNZuLPu9FCTMmY3Xw0AJVTWZGADr3OmX4xHaOgpQXAWxZ
YbuCwWHAc7ANECnN11oE0SfCtwu5akfnv3ni31Ba/bDX607Uh72N0b0P+AqLzdNCO4S5sIOx8ku8
ZFwq59DFSS9mqdLUTsuaLa3FCr+Sb0QxWnxyi1RmKANoYwgo6mZcKq/tPCD5oNvchroQzjDyeZX8
LtBWTJwxJYXDPtzNE/Pe/x3UldZhw8R2GkgMbYMcfK6hIoLtKB3srBONsQiS+hQVQpRsgXumMUjn
Xl5isxzSpT4GK556JSWuKtEMMm3/p1DeHKLBiXGQ5h1GyzUBbMuM8IUD321g/GA2l8uje3rzNi24
rQD83jB3XYoBK1QUu4ES5+Zw2tGzt9Xi+poiwSGy/7S8LKF2RiiWx7vfccbB8Bl75rVf+686O7Ox
5F4FiDa5uBMS8xBMQyl09n4LH0ryRP0xEAUMre6ODJGK3yQinB3UneIqTyxpdbgzlfWXfelsiw94
hnXmdkMazJJz0qLYEjLdLMpLzkybGZ8E1vVq0PeHMH34fnhcZdIiu8cCZxiKQphaIWs1FFxF9wgz
d5R2SoxemPAo1JpEPJm7jBGVOvCTxEhwVjTPolWmOHWQBov8+FnnVJ8CQDzBay6DQKSKlLR0dcIT
b3jdATm5LmuvK7j/l2+pw7uxSIUTuuTHLbZsNQyZRfpFSlzb05FxAtwuPBMbVDCUlt35YXlk2N6s
R+ay/mLOBmQUsJ67pnIqf2+ys6b0H9EWEcjchINhuJcbIOOHOylqq9L5doYNxrpSn0KydW9+ENt9
afNKE22PKU5Uir4WIcR6Pddx0T0Sm8b7C1nA5TG8okh1kgU/K+tY1HVheAoAHxjUWIdKTbR0pJaw
rmBMOMYvnvrGzJzWTxpw3LA/J/JtGCFxfIJYjcKfT4yk9pE3272ACVOqmO2tv4iCtwmWl6OdAVA4
gtFSjio9kucosU/4vLb7lAmWFWLJHE8+lDOmDerEI5xwhiBgkJ+p+DlRAxlL5iOPWc7dXUljWTvR
vMJQTBINNPn7eOO0W1ClgOzvJR5lmwYCxj2TlqVSDo8qILd5aSISwf3aXknXG6Ze6MoXd+dfNgCA
jnOoI+ZGWP1vDOPuf5bcq37dMxQxygY8oc+ChiGYp8aX3aSXhoqD6PS+XUdUL++5G/qA/kOKGa+N
98LVZC884AMHMoAbznuDyh3l7pREh3iUBRcqc0YiGGa5KqGR22zi5n5o1fwqnmUQptei1UpURrYZ
2g4MvgXzsHrjWKZQEOLREkDhNglskGB2M0X2IsBLxWF28ZiF4XCmytQIXm6wPGWTi+RJotb400f9
y7ESWdjYA9viTEE4a7ksXUxS/lb+clq9bTe64yrl9Z3KsgTwbhGszuV7WMPHQYSTDzi5tuj+xYy8
2EM2DOj8oWd5w9oIYYmQrBO86mBwJYu7ani5FjMjidpT3pUm+sqY3iFSNOVevcAPJ98QesXVAw8n
4+mIgOLp805eUuqZsE0ZjICHd0a5W86tJYojPeI+7Ed6rDwIpHwZGw86yo55EIUST1A38RXgKDUi
CBFlkTEsChrF0pPs9QzujJwT7qb391e7hOJB8sq8jCYk2eOkrrH6EszT7VJCEvPMRk9BdxTXwJO/
soTB2RiooFF38SOQcw/jCp+iiy7oni8Jb7gW7xIk5Zmc0GX1VXePvs2d9v4MgxL7D42jaeOOumM7
hGEzut6ga8IdUNUz0anUtzQgJ9ms1dwZlU42cdZixpNqUxDWtsc/uJJ8yXMykGRF5mLlDhk+ufQf
YN00EB6PjCcWPAzpsKMvhqlSh93TuHxYL7gsgClRoP/T9IAZoIMheq28up2oP0V/1G//pbIxibkO
9TyxoZ6dtXqQHA1fdoUUVPX91TIMYqnW5TkYwnDmcuAEpTQEl6HK3nnuEFbyfn0dMYqeaZIXFbTI
ZPDI09TcUn99D0T/fPRJfuEaRaJntHufew6jGShAa1Jsx3txQ3ZyR01u8/tP8Okn9d2ffdH6e16Y
c91X34C3q9JHJfXTPv+mP29/puIltMs0SXIeKjIGLm4bzFgv70xELmH36KfXBZMcl3kufg5kQwza
Qe0plPrdlafIZhqt26vc7equSHMGTnb5I3ts73nbAuQHUMoF8pnTb9+SSGCazwRMvKZlfjP/3JWP
cFcItONH6NtRfkTL+vICR6OmGzV3Z9FPBtrHG5EUqXkRRY4yi503oak4XieIhAEftKwUZeNGXPMs
Xaj5yXhN5psGBU8Vg+5vK39Jx6OIyUENh1rgliJ+gDJ+8G4E73Ha4uIhJwzVwsiiPU5nDcZMqGxl
46M/WS/NvkfwLgu/Zc39pEpofaxe1oq/gFrTSBC/+yCYDd2Ar1hhZKTwiM8KDh3J/X1pb0E6J8FM
5dBaz7AtHEq6UD/GMpd9MoXAxKkffs4Ez7br7GnUGa3ot7tabsJwrWq19YnCCyjMu94q7VhhaqOX
IvgJb4o7EgsZMOKUkRJ++1zxU0dunFUTFfSDMf7+e++Un9FbOUL4ZRl4HHmhmR4+eI3H2x4wX432
HD/HOb3H4JNuiiosuv5facFmsLn9z0C3lUytmLT3xoIvQIkEjYrDKjK1t5uq4l0/abktbrE7iS4o
RJ3FKBHOrlMJGdQJJc2q0iGUAzzkZBy+zgobtc/VqVgfZt8mOB0O6yp32oqtUWrKQKDg7ver3aTb
Q/8dhmPMKS7MJFf/EMWOpNZ1s5kcyYwEdwBR8TaSKjJBGJRHwEPm3CJYAxX9FTpWOlqz3WAoNchB
vh89PC+A76RWUuxNOh+nqfOFGI5602zP+2BVb6rGfogb5+R7vqn4VFr0vNeNiHy87LlEM7ebYRvq
55kpgOeBhZvgBfg8wr5GYscwANheBRY3SBPSuMIO+ZA6//NadmhvUXqvWq0T1vV7KgNPWFpvm/Mo
xembSWGhuWexYEEGbRlbyvQSokFMS+M37H9cDZqwXkWzqRwuy4WeHLqCxVdc6kE5lKnkKHklmCNn
NiiLR2sNC8DHl4K/oAs2yWOC+oWCwlYPAKf8M7iAfMG2gjYWGe6/mvmxnB5UC0rg3yB1nUtxu+2i
LzUB34yO/D5Xpp9T3GaZUMSk6gOR9LKQJWhdM9jkQkfRaAOjTYUB1PRyQ0BGzXa6aYdQ1FRZPfpR
4KssGMfPKdMQIS1uwWOLVtnG34+bjHb5AdBFI4sNJIJ60HQ/X0WVp4pMDWTrjSPpC4EBbi9sFs7A
/P3Gng+3Z3x64Kz0TSzbjiez6sAULCFZ6CFJCLpxojlgpVwGnIU7bQLQEQixtOjk4efwhK/qPJsW
BAizNMYQv/+5oBEgBxzHz6pX6GFBnST/sqTbdMJWVJFqApqwMn26hQxIxdkvvLovKjuDm67UaqmH
ELkOMAN5xUwz48X8Fbf8sS/K3SgCkq3QT/DHID93kl3sC0h/1V/AX/a8gBINj0G6pY8AfxlE6z31
O4sj0N29D8eVvMR0ztCsJlnRulCVrF+ZosLxo4rnMqKg3/IA5GgN+LZI1spWDK2bLtjcY97a7Xki
Q0Yp6ExkG/6XxjTROZ2XDDDkqUG9FCqYGA/CAPmy7FHYpiUi3zgvpyiQH8KXMZRcD9eg7RBEpwvE
r1bTZnTn1Wdnk5ZnXY3xsk1K865pbkKkTuPkfNmyk/f6GgCdXIYktFPlouezgfzyZJHxxvVPCoql
QuXyMMCCLM1ns7Tu1YDA0fn6s/na/aB2uLWP2TbozGxPAU3JFSDprotXMZMnuGugI/SNBQIk0pDi
kZVuIw7O7uFXtqADiZipSB/8UEepZgTVYgyfDqjQnQeNPOBQ1+sO7OCIgJJGYqC+bSnXWVpuEsZp
PxiFls0MQ53wv1a4pW/UAL28PqcNs4Dyzm37mmRZ6ru6xrj7Mq/xIN3mXr8pbNkBRYBNfSoLprWp
0Xvb5v538ra6BZIbRKMu6RtQPgzau5OMDac2O03EDXHArc5Mth7NzRf9ENjt3/KajqosDCRLvKdq
6uKmOa1qW9iEFKdV+b/5rTxBP9DKpCCWpx7LadQyGar3HCxjfbVapUOxs3aEXRJ4Kf2aL9bNIGe0
5zxUAhGH554CckZgOAmuYKd8N2wZPVNarDwrFV+VbMcmNsWOf0RTVe+nLOTbn8GT7of7TpeWmd0p
+eqZAdCW29teVipsieEI+lQEhKA1oGh0kSzNR/KsKW229SXq5XPJEI/BNMNdId66EVO6BKdoK5mN
Gv79rpj6NvAwRg6J7QIIBp6LkB3PCpQFiGDNNCgKNHFe39LX6qMol+0lFlRyGYi/YAn6FLWzYOxP
CB2turgFNV9Bp5Qvi8wlnpTsurtGa1mOr4OTotzazgkgq72TIjjT7sFeEriimPs3rKYjySTnrbE5
Rc14R/hq9hsKP+4Ow92dJhHcCt/68pTEvZX8mOkibCkBnD4j8luizfGCBKN2Vd+2hxQKPiT9fyrF
7YcDHUP42C+jDaDsZdS7PNpviSsim7ttfN5EVRD5t9mr9+YdZUynDuGwj9jYYKYb+WdB5UifPj3A
i3AlwNypHPQBVNBbcJOYPmvluf+GCJ5KkEn7vrYglQnghQRpgZvOXLEiXweP9n/ueuYhImy5hQ7P
/V1knO6F6ES1tAG2RctFKffATT8jGMl5QfOanMGFmARhlC5K6wX2Xs7QzZVT6Ux4nv/YZe4JjnUO
/VibhFWFqXWRqFhaMoVtx/HFMwRqmmh9walRzXYDfjKkM1dbtLtkqWs3yhHlY78zClPUwLA6Npi4
qZDpFw7PDR0WUVbsWLMGEXrQICIIqvLZUmoHaXlRutHNwyGPy+lOE/BFDrLN71ikhrEWB46Irhq9
HuE2bzIBufbFyoGT1uECRVSOu4843OzKzEQDiXP+o0eWVKRdCJswJ4wTZwh6KbPAZ5oFBNfvuVw2
yYH5qO/1sMnLolcOUTpwC0uTYEQQ+laC8deFbpmHsAbI3PJ8RS4FQ+Xw5BJpmzI3pJujD2015jyh
J8lkJFcLqDnvfIk/WHbiBWqx9PXxwPvu+99fLiBMNsRRmo0vdHXzNGzdc+7zhQWKzJ80dpPoRLAs
al2Z9sS8NwTDEFV6JQruphUSzbQb8RERK2jNOK8CdDq1Q3JATGApmW5zm6Pb+9JzPEdvaxAp3rNG
cgcIvEkU4ck4sfc7BUA88L9JLuzy2WIezIb4SpzeYOLaisvFgdOMMqSXU9rtwB8ChyzVyqTKB0t7
nz1SGFXW1VtbPLGjN5rHQ1KG0nAD44kwW4mjVTNYDdEgySW0DuAVs42jhbepEYBreThmv6X2DlNq
Yj/6KL9aFgzoTJsIZXKiEaCXN3kESUycxZWV0UOpslRsJl9bIE10lqqlCHdE2vhyUTLn4LwpxThE
ySTb6liQholn3PqjfydzNrcJDj5e65LuXIN9PcS78fW1QpBB1UotP0/A4BeIh/49+lfHhMQdesVv
dgMEB1ugFCQKSjDL5oNHD/QMFDWcJ1NfKcLGHvbMDR3suu3fB2b7VGsJ0PCg33plMMA2uhfRICNy
u4Une6Fu6RE1dRXAXx9wQ2mdgeNl2EpxPuo9tVrphyPfdZT1LI2+T0NTMqZzvE8Xo/CKHqHz0Voh
qZeijI4G2yVVmGMu6My9tjpeWFomJztaPKg4wDU4wM3V5u3DPtGR+hA17K6P2wWJmGxGEag/9A2j
m86xi9o2vV7Ss2JtK3RMo90gx6cKRxOEZiTgbyA6EhLmiySxMzZBIR+Lz4ZBaFLW9Dd2g2LDFpeG
omsc2gM00lzuhE2jlBAt3IkIR9ZD5TQ7TgYNsNeWfgNcnaUFox1MVR48vJDBtEINuJaOAvR8y2mz
zQRCME7OhFCrTtP7LQniGMYq6gAF4zTIu+VLUeV9ILVFHa5Z/zDyhDZoGK6ZFZ9UOC1I1cTayi4A
Tg8RZOq8wrNif4TJALmisE5bhHZV/ccgJnMrGDWMM7Z9IuTNOe4uRzow6797mMVakX62W+4l1o4h
ybCeffgcEhHMF4vJUVAxdG+jBW9DfEK/qoDORpBp4I1PqAwncBwJoy0ZhWu5JEtkdpEFGRJ0adie
tEJYJfBTyjJo/rfUHqCVAJ4kAsuHiu+6WYAgfK5MG6RqqtmppoGFtuc36BPJHEK5HZyHnMKj9pqM
2oToNdFNcUuDSIPdiCqg4AtM2f3mLmMPaNjLlI8k5GIZnngIun/0LiEsa8D0zV+NJd9kp9u5jtZ/
j6PWhf4kY1/5YJ741KAehYvBh1QBFQTanIfz/CKzJ6WTNKlNZ/3lGgI+x2dR3O9dOjbri6Y9D5Tl
Xz8idDb0/36G5s0du7SQFMJJxLkqTitZJ7PbLT8IZvCKQuE4eDWIqaoR4WBvfo5Aww1KIxq5ujaE
h+z9205HY4kjSeRI2B/Nrvm9Ujp5XOdAqVebNeYTI+5Qua2OCXBoEo4uzkMe7h98cCuRe6eqhyfe
+rIC7ko2rDbkzU5E/C7/v59FuKbvQliVAWMZ8AzWfpEjRGYPI9n1hOBPA63xO+5cxG7wQTL6Zlcm
OCe/9FrCLTO+9nO93e3KunqQBMF7xMNhfXdh2wMMYRH2JmAGssf0SOMTNuaz+WubbcW6v6Hj2Yvn
cRs/XsQ4n5pNip6KZTBPRY3hiKJvIlXmOgsEtH7x7OB28FjTUT6oU3gQG0OMqbqjs684YoIbXATe
J3MmpTlok3fr6sXYWVZOvkbPwZ8b/gKIoIRabsOKqMw4F7MYstZZYNyAYrTjhBUaggFij2Cljfyf
VAV0FujpcOR9DYzvTzx9fVwc5y4x0pLt3WaMj5Ta0964z+rL//yL/hzV3FKt6KifSqb3KzJGLQuG
EVCxIngCNdAG37jTGQ3wb8pmwvLxN10zHOEXIn0XySFEXtYAUpEzf2Fh+aF7k/uJ9qItCzRqo/O+
W9mFbmEEMIMAFB3vb7/PRAom09GwDShqKQCBjwRWssr89A8LY8+NlX5KoKIMrxxmQF1rdw3oWxaH
v0/SFX/jvJYw28cB9K1bYVMTkcc/jt3YRaQoO+yDwz71b6e8ZO0NLSUpZBJRnOnbc5ecaNvnfm9t
EmaRfI7bQ5LzVOxARnk3YDObPLV6DfPfx8dn7a4hKlJ9qAqjiPZLdL8gjKvXNmcye4Dqt8rwugrV
c2hiYaVpB3aD06os7oJuLXcardCFvSxoIC4XDv5D3QDFY4DKpiaG8i4jLGfLPWHeEeB1fPYQkGVo
ZxBaCGm5gLK14kHCYBtJ2Mitmk4yyWC9q8jv5G9ohxR0W687oBiWZp4yhemWCBi+PiNertEKpnEK
ICokJr4Fixm8bJnvlq5o6t1jEIJ2WUkQCbopvLcVTpk61wLMH/8Mt002zFgprRnhdDSELIRXQ429
kqmAg7XXdQ0EfTBa9ettGSUCgRi057iAVuUFc84xm+YPZF5Qr1Up6baiKte6oV5cW6zc09FNk6SS
+/FIslZs5XMSoBeqelKRQ8rXdrsVX0W9jMrdgk6YPAuAMSbiBR4QvelrBZ9GrlNT2VuQxXm4uCNI
xeMiGaOLk5yziRIs/swDQVRfFS8jKleneLMLKsGiwa40zqIiq9W05+ngjpFrS6gZImU7JP/3Hluu
4vlE3Vl5oo03mVLQwjbVbJ45VfpHhkPCOheUy09cf3QrvxX5nnzVZf3sWnQ9Q4nz6dH904SdiDgy
WC1HJ1h2/Td+gsKKnxGxtiyZ4n6v2GR0cFN+FFTDXnm3x+ykGqqW5mfVy//UFKynuDZWC/g0mHKe
FZ/b/3hhBRiEcxjhydxFXS4aC5VL7g6Mc6rZdIwqZXg4MybVUYJRpKTHkQYjBht04dMbnL+gfhNX
8yRCb1+6JBe/SbZRuG81VAbXMuCU6dk+C+1CIQiVdFlrtV5paV+OFUjlZPYWyKE9OGC+C2ZAyZ9i
Aw15tORWvBczmPdJJv7/n4mcV0zsgTmYzfAZljBGN329mYYgLhWioEdnl//v0lciDyLc0RzljZ52
g7ahWiuqbMMsTnQV5QGxlo8V26bYrKdoELJLQiYH8eqWlJkOYgwRjuVs5DO1Zdu65mjlzT/cw082
C6/ayv3KQ7i7noS2WGo0lkFFz/GmYZA5pwqTGPNNNgm3i35FijAwkiBuCTD5n1+BTTb3YWUgTZPw
3ekw6aRThdtJlcqiI2Gm+3GV4RrkqHXeR9rq8M3IACtw3d3dJCYH41+0x+B/n8NLnTCf/yiK+U5L
9VWubfSzQ9uNfqaJyDbTiUs4TN+ZHozQBQAb9wUKJORhHPMVHR+3HrjM/T7wxI1N4wJ3e2TOlq9X
BI8iU4YpsOOhZtGthBZGICJeUdP/qPSJiP7wxgziPyilwjvQrOBHRyk+1HXo3xI6gcA/CVFFlckZ
ETpM3KwINzyBZPxsUfTC/2p7rGV5Enu9CFbEVLSoe7kxK93oFUY2pWHM9GdsqhX//xkxKs6nCL6S
kB9mxpWQ8dPjPlb7pZ/G0NCi1pIGkiEuMwGusLli9pTj2m8xpWMLWpM7U2b2kooSdg78drX6XPYG
KcSyz8kv3rxqTne4x9EWRT0Pb510NNJhkes9DJeCeNFBTNk2yWTw2pgP+2EQwpEoTeouY/E856vw
kBDUp+/mc4canj/aM739aPpsrEq+eq6X54TxDeuQExq7LokP+5FjqZ1NagcIrseJXKrvRvFIZInj
VpOG/dsFg/imVA7yc9SFAWXkY+5L2vYPihdrW0n7kWoMXDLXNLb31BpYduuqCJvP8a7gzff8Hg8S
fdrzZfhOyvltlAUKvXH9wbwLoMXvYpMVuhTQ8VVP3VrTZkRUFhWtM59dGaME9s010uGIt4Uz3j67
wtlA9hUuTg9wcl78KnZkH6u/VhtxyrDTWZiELqAXexBEJhm+r4qo/ShJbKAYnRZix5X9gL9bcstR
FzYcQyAX1Cge7xg58NqtMf/M8RSIteNWRMJRVFzeQVkXwGzJJ1HfDgGhgaWulC8RlbP14mVf42NI
W2Eu1bzuEKp7Gh4GQhrsnadN2lFPZ4iJLNsw/Nj1UxikLW6PVT7gdqzSkjc4bjVMmTOrA00hUIuw
5R1yg02sZihpJ/Ha7NmdbUWsfWasyIlorJwX4MBmzpgoLKoJtdqsOx40pj5SCWf9Q9BvxCtC9LO+
aonAcvi2Tvw0WzXeyf66i+cSvjS8BUbzjtNMb//ckzt077kdgrUVEqCF5YXpjaJOYlvii7RccXf8
8eepksaWe/tQPmxtYdfo+UJByG7SiUOpxa7s8SjFljIeIFYJaAnFF7RzBOknEOCbcoEOlrMiYk3G
vxXJmU3+MMMH5VAfwoXlB85ShwmAfa0iOmcJNkj/lvtHclD7ZLSaPwnthaivQh5mnPjiIqGBhVZ+
2uvxaWb9qLhaO3lY5CUxAWqMuFp91tI050amJWxfWnOVM6od+k7zV9XbKeg6Lp6IVBtWg/V2OTES
lkArehl0CZhnvsmKjmlApTcSnSncZ5A/9GCeONgVxeIfXQ5CJYjMymm3K0/Ytv+iw5QvOCPbbFfC
zaN++gq6QnnQwrATfwo5ptFajFinWG4z8dG8RZmAdJQ2n4yzQ6UGaEWxLrHzKu0IWz8uOF03P3VY
fl8f6nLTjcybNC+oisa2E5g96q6igwGGLAX5v0VehzCeU9uzcwRGhTSTXl1gmntzeoiPPBVtxj+w
VbkcXrqt+uHqX+LNFtMWcQqvGRF6QR7Qvq1Hk44LfR4USpr/TQAM4ptC7TMNr9EGfb3f+f5boaf7
zPpWbBU38J2uqu+GfaAydjy6PkYdnrYn5ev7b8kB9V5BWICPOFxUVpafKljrZwbwVNfT9cZcUdLU
UwOvPCNYCaiFDncV8EbZyuXPHeZdMJqwCrz2UaJyMR4ds4rVOdDN9wtw/RN/OEPrsXZPtf0/2fvy
EhteJk/0eUxBtzgXo0lVt6DT4NiJB3h+6sUBtLrZrEVLoox9jfojAmFb2ZjrmxiXu1nuLXUAWWlS
tBsqBbJZ3IWy0Nkt1ZYEt2jxNqdIipd8osM6zW13E7nMpvxLozmkvloJqTK90cG3YsppfmPrI4KG
wsOsQeywZvitiXE8/3tkAp1HIa62RztFF2bH2SlxetZjg9VPqSZwD7FM6Yk7GPR0pn9AAwpqoKGW
pYwIyXHCHy4IApBaihZxWzm8wK/9HFua4v70nyskMWno4ipkdpkmOS98AcRRjEX10PYrwxsys2YR
rM5rryiaFoNQrE1wpZRQxYZUn+P7qSqPmhc+/LffqDTuDoL4OcxIy4cp4nWqThbsBPPKNhVe1lvv
DVDxk9Q358YcgOeYYIlGaXDOam1VqGlXHMTVQCc0TRdCWWLswvJMuN5G94iISUY5TtFd7k8l+yl0
x4b0+SB9XJFIjaEmDgZTBZ6biZeHEzp+eMCzxPXZFkufeoNOaowtnRiIA0f72PXNW7duNfI7gYxi
jJzufEjBImG5K1UmYnkmMwwZrOStdAAxo6lDwHaM5SS8r/vbG4JWGCVGEPL6tDqQGKqmQvweiQih
1/6RFpyYCgXKy6KpfpX/X112RBlWCf1JntiU22qOoL7XCYaPzOr457DUUeNSSizBu8PRrGb89ePX
36SUqf+q59iMRnLsZFXriOXrK3UlFuUWm58lYYlUis8Np3XOrbzEcBKVzd5hK64msWM/RQA6vMFA
+pZMXJIro/zxYJRKLnyiFnq3yjU7gByTnm8DIoppa/S3vlZk+sVDtJ1GkGrh6YGYUTlFpbDOUSY6
RvuXa7f5QXsi0gfmprdXThHamguPmEBd/HF10dAiPKFBxtJeeBv1PC+VThUeORaTa5anSRyrGpQY
ddHKW4k0c0G25hssdKLIQxZlLPM0eZiQ7nROMgSN2dCASA6zQRimhRbKS1HnW+tJ8h44BpIfp61G
t54+hwON3Hu8CSD+Qs2QLuPcVghbn4jvZl+8rUJ9S4V8/mUCNj5AjHO+m74WXDzkWq1dZIy67OJ3
PGAIIsm6faaVPVro7AAu4PjylzKVrM9ga32js2CStH9Y+KRuRYVspMObSQpeFF9qTx842JfgDyl1
6XDg+MdA0QVyYRl4tdZWpzf0NHYXI6d/GLNcg3BnlY313FK8/Tvx3v4Tr5aXTi9sJ15Cd7vqpn9W
Ox05VBKnmH3UKhW9BhrkF51zaUHo8/PV81B9TRSqnk8RjLGbAjj4/+BEEDwdzvPHvDNSeaKnWKRm
gpdIjgIVFSGQoz3otbL0QommnQ+uTqHaput5YHN0S8Qb7EzvS2ANBYbG8Dq8Heg4+F/D95XeybyI
OL4+elM1aAvVTG7o2vvkmge5xLYL4LDEZ+c6B7SrxPHjJYYbM0Y9UiwgezDEplho4FNMkYDTqZpK
Irrznc4wbwtNzC611jsdSHJ95DuMcN9XpkumaSvs90ZfdmH4yNY+4ObxM7VsxK8z+A9EDFkhB0wC
H3WqVyHErd9aaHBdcm8pgGflZKDlLyVEeLs0KEVGmceVAj/cl3VHdF73O9HwfnMHDSTUJCWg3Go3
pUyvnw9iRDNceGlo1N0VOUV5zqT5TWbNUh/7LnpVMjkz/xCGoUVvnnj5X1q8Kleh4GuMjTDVCTie
W5RO2Ink5hvVgNViAjcmwQn72/43sHpAie8GtqgK3sIJ3D7zh1Z3Besk9jpxMJIdKVEUp56+7B7s
UoBaOrLT5kXxJqrQbcPjdTgPD5z/4YRatSpzEdIzDMCRIXFLg4+DrzHxya+Mp5JVwMjjn+87IhS2
VSpwydVoqsyBNu8wK7UmP5wj6Fs3TlqaMJesTDToLUaMnG9Cvx4P3DT9v7Oh+xQQaW9lRExppz87
YgGxMPncxw6c72JwSEytQOYz0pqvc7hPy2axusLi4i9/GqnnNLh6rOkcAMRD9jpAQNagGgW9gtkE
tUhFfjz/IR3wcOxeJAacQfigYpny9UBZcPeMkO8NYdO2sXaWUljJSEqHt2LuHexjRY2ybvtfZPo6
2S3KoFteVC667OVTbrTIr1MwrPCwgbJiqMdhTA5js4NU4xqf2wEt/XDeFWccLoskLodXJ/RfCJ1o
KO2dFI1nwRqRoYJGihopiX/+Y3vaf3QXv72+DbU7MzGMpJ8d2dWaW1LZyc+gca5WilrvaV0OXcKo
nC8kfNhjfYKeZeEwdcHY/Jl2gAdZjJixgFAi/vX+3CBAHKfF6enfhNqXauWH9nolJGWbHsjw9sGG
SkHJydIvD859A6bdlsmZM+ctfeJcn1LElheA9+U0yFdDi8ohQx7fcFsVnxCE+hTZL7eG22lvd+X7
shWBYNaeIxgZRMko1v45q5ZXpoe+9id2HUFIXLF6UCmDw1LVF178TTa5BUmBM4E+JJ7pm6S4zb+3
fQSJ2Q/nUQj46uEJqZ+LqCwVDLZRQh53hybNHkPkSLrygVWvF+k/12DAkgazIPm0ToSpDjwJwrJc
6B6UwNw/PCGruq1qnvrWxlYdcErml8IRm4JpnEf1DmQwJYp0oFRGFJVgY2SuqTQgMMu7OtO9Jrh0
bR/A1F7+YYcQKbvTtCDpsDPpwv3Rrpbp32rLlI7doB4V3qxCaoKmlLSWGusDFsFucf0N45Ho+9N1
ZHEcuzRGlYNYxdTwoLnihoqHUzDBwfqvwX4r6ct9dyPGN61fTZrAgCsU/33tGkoErxuHANAY917P
1a6HgZZ04uwmoZtFGO39/GLSeDtlY+0hRVGf8plbWcTogrxZ01bs1OEPkUzPKi9qtJfS8kkOzU9t
bvHAxeaev/RJUkjUxpUcF93P8F82O5Dw1kbt/wLdk8ZCgnhfwkdcQch8GaD4Q61kr4TNqEZITHoI
EkCb/ObJI/k8OG9byW12yiJmoC1O1f9xdMjBPGG1c/Qhp7pw18B8Ln1507NTh56ENagzoHusb31x
mRjmQQFANmroxZYgopPYXp9WYUqVjdTwTUk86RQ5dCBsHvsieo7P1+icLVSpfv61e0OohLLIcDdw
Kt/Q5qe+QUrnT+0wmaM1mMD/YBc0PhE+j5wzOtAV+nBZompxtLq6jCWEIpRC2V9hoLfINTrFcdpK
3qq04HueELhgzZWHLJzRMnCH5TdFHY9Jr9QZB+J/j++3zl4rCd2UFa03VQ6EwcYnahM6UuxVPvas
CvN/83kJTeFpaFLDQt6L3wFRuOZdqwhqJs2E89eQg4+pJXoFTMvIreOH5CR0yyPi0lKfS7akUjWg
KetWxLqRMOOULNJPFF/bMBNlslrTHZnBqCpE8kmm39jq6kSyWfHX8GtJ6L5uRqtVHDc/m2P1gWb4
gHtrvGPgEZ1AMZqUzTem6sTDeKVKdiJmGEsxX/IMJtNY2LHGR+pHaoOdtAbk/1F9Ys1hw5GSxi67
X3QYukVd6O1k//diKHUIRS743v/0pxor+LYP1Yl2dYyNKdFH0FY3vmfEA4O9fH24YwfG/Qj8Cah/
Ek2/omRDMChTDdawrkdnbLkBmg9i0YDNfDMqAE2Wivdcaek1wNMLLNpuKz4ttSx70EuxNp4KouCF
SqKNnuMzH7V17aOyxcQJC1ZwLSq3TFgTGuL3rUGvZi2Q0K8/63idFwtOk0/MOAAyJvK0ntXjDICv
g5Z6iNB1Yrx/2BJBILijd5oSIXHsiVqa0pqIsm7Bk3nUi6Dlhm8M3QB+DBCC6HMNUhk1qcFUI3sH
6asofG1OzmoEijMWuXcPil2KR0ZvK8RrhsJtYf+yc06x1f9C89HlMZr1YAMNPO/JK0XOqS6FRKPs
9tk9qtBFZ9HWeBzOE9yQWIUzLzV71gB9sMyBEujIB3VhRKKzCLP2npxZIxsfObPBI+Io36btO47y
zVAtJc1iEqT8UTZIa4lu5Ki1wdybBwNBY5F3i3KcmX3TTMePzRC+2w1uaH1586nSBKgv67BtA1W1
an91u8BZgNagzdOdYO7Ij0cjD0sn/zLNFl+FztTnWoqQt951MZPI4oAPdqBKv5rg5VueZ4jurAtg
ASQYZouBU5vhYCihxzFxJD8AaTZqrCmnrmcCVBcRyuJHkoEtqRzU4cAlRpGTjNt4xRGOxEctsKX7
gLAAYgU7kCtCFhCQn2j/vUDZFAx0mMkiKrGA+I0vZ449nUR+4wXr44tUk/eATWp1M0ZxYE+Pl4RV
XiaBnFPs6KCLXEYqBC1m0fLqXcgDhF+OS5UM6lFgJ3A3M1TAoyF0Iv/AyLZ0ST86vkak06wfY/Cv
xjC+zOMOi5PTLJo2XNtsUBLKTYruGQ54M19O6R1Ie2hG/Poyg8mABRECmpn5ZSo1Lc7LHXRixCFZ
tgOOPeQXU8r9v6Ja8hjqPhoOhL3Cj0wOvheQI4tFuI4tOuLMPVaM+fRBDwJWaXhF1bFdbLSMatQ/
0ANZDTxBDPUfbY5sVWqfpOQ+wvYH44xbgMUi+tThO1GM5HSx8pWYAU89FP6dBo4VZybkHubn1are
Iib8eFkl3MZm/G4lnZl2oK2xQoo0cbKrrkDd6mWV9CkxRftmrwijNVBmwL6WoKJbJ1VPv4eySYJ9
CnNrGcOC8G2GQcmZF++YW+3MXU1IA3XuZ2KJYZYdcgCmWhZcPY+ctzkwjkn4d3eYufbvcHrXGcRz
HZkzOkosl6ztr9RRn/GtCPCCX4r0C3NXgz6U2xIv/X22iPJfjR1WV3aPjWMeaThWpwiBtZkIg870
0J3USA4cLhnIn7aNNh3ZipxVEj9QZmgyaP2+Vzu9vOa5K3OVhp5C1UjUqoswy/hrjrO8Z9QK4XsH
8t3ueD6r3y5ZaFiDu6r+grzeaePfKmVVUYTIgJjXt6lsWRcB5FPrbZraIhjeInlOf4005Rlqieg5
IgNviGb/pFhaW8F+QZCVwypOxhXkxt3qNom9hlOPXsFMSmURyr+Tagq9AohZKlHdQd9mk0e5fNSK
jR5n++IcujWvmhD4UEmFbmaVd+HIzTX+dz90ZeWMoFSiwyA5wd7tGOxlPp3YDZRhhmgF3mJLyEIq
E9mAq50gPzdi7XS9fcG6p4KBZ0kIRVCJhrKLnZW3/dK3R7GpvXGTIzPDjjx/pipSc7G55GGo7WIu
YQtb0YLEIQCCXF3oVq5bZLfF2VA0Ayf5Z1/+7/l4yAGbhXbqHCBXu/Gi67y7HW6UswNzmXSN8Lat
LNxiP3MAXcQ+U3WkXRnRe3/2AQKoxtDg/VltmAJpDouBw2u4ABuaUuB41anmVmgnpQ5x8S8gkHOs
3RtpsTMRv9/XZUEQkiNp1eL6tO52vIRWMGIN5HdO/X9jpkrNQt7P1HbnTScVPRHt9nMflQfjt25W
hcX7w5ZQFRaVfz/525x57W/XGGRJ3lZcNeaUx+VQIwlBOu6ZOxxNNdogpc9X0zcRX9SwNQbGuPYc
Nx12vTmXVQbs2orkw6QOoDV+B3vsqTR22fpOhhBFNQ3EgobkSHCAL4qDzgSsxIsCmdtR2yG0hO8D
jBJri75pFkwBk92Hom7JO5w5NetUg66L3RMqi8Fny64nXZV0qLXvsLzXEhsXpsdZIZZIXekPCR3O
xbTDQ+TvgpTSO8Y5uiuNQ4DBrXutHPuOtbe5V6eMxTUHDU/wbQKl/KusNifLQPhPB9nCb8ptyeCV
L8MMTvJ5vksiEo9be2o/OXFeRsHY5djKn7Q7oawMZ6HtRJU5VYtUM4vOnmDo5RWZRo4499AsdCZv
tzsvv0e6rp1ojB38uhv00e7E9KzgQPDxL49YQ5UubK7uWCVPd3tg27egdnuariYeBvTE/ky+Sc78
MzZ3xnOrhCsuS7anI3JRJOIdwaAcZ7/8Z6/zji2Qt+2k9PjBICzwL/mnm4/c+NEse0wc7/6Wepps
iWBTk92qkKoql7NILgAebEqp2D/VfGxQ6iLyxgOgL4nKlwghDkA2bKGpYb7buFIKEbnr49w21byq
vpQFdv4auny88dAoo2LXcl1P9DN1EuhVbyMeiA0b26b6z4i6+r46nmth8jDa/FT8uFqgC3IuRLgA
2walbNkOfMiFpFuJciW+Q86DupqkpOt/EA+RoEpY1qjHcmM13JoK8hXv3BrLtfSeccNSVZCYifgj
FFHdyhb9Jw2FOiyIKZFOlIzZgjbHpP9Hi+ztnFPf2kdwfismsgEG32SC6ntE88Iq759ecIt31dlc
EuUBt2lyOQ0tOBtbWf7DtIHiRFgbXHTDx+GeleU1obrWGRqKwPrg24S1RKlPuTmXBGxqMwl0ZQDn
Ub6pwXan8FYtUXR5/1cXFp+GYEfWA6AULIkpva170cMIWD/TvJq91lqKPWURxJlbpnhcMljKj59e
Sa7EF02MYcMf6oiTFlimBkX79JWDFOw8iqGSsmB9ORikwxDgXG6RM14MuR9CQaWY11pD6LcIdWGV
zzTOTq4i8usDapEj6LbkYWLLQ43W+Z8jeZiC0EN9fcRrJbrX6PI3CVPDVx2fpOcvwWNtO/yK1ulI
GkcuYhQhgT2ZwcLwRvxViBqiwybm0emPG5L6l6OQrTrU5sddDNrJh6+3oeLwFKSSU7GtKenn2Xwy
Vj3bpvs4NnIOwEvaTszSUA0aQ0O2ttaa4R4RjUObPUj97Ebx/hjpX2uwY0QaCy137Xubs8xafGKd
8u7dIzVCq6QmG4CwmqWCz7C6HN7YGcCoNeJakxRFyDNNheKZsaLUQ1UWvrAOFvj/tCG3Z+WNz/ge
EMY7KQH/i60RGsbgZ8rKR5rCyX7NFhGdo3C8E303B+nMEPRClz0tqlNZ0LT+hBAD8GnrsdayXxmt
hhHzvVETYEkZ1M4MkvuRX6sGFFk45UXkNAMAPD31gydyI3J7oAV3FIJDnSVHa88ZoqCkj30cNvaO
070aBDTeKq3GJYb0YlE7M7qwUnclmPN0AqjvyyxkuuMWoybUZiwC2pBOhC06ydvXTWyGgi+3Uv0y
ygsJBMXGqhofhYDT2njD2sFnqozkCJnGc4DR8hXeZiUs0A25rayuhx4YgoI6m5QKKc9ylYx10IJG
acV1uUp5+FbPsLnqu2Ng6pa6osbKay/MVzoyC1Kl6XG5Pt8xWvYs46q9xzkDF0tHdIoIcXgmU9/b
GsivEOc+7b1RCnuKL6Xub6/DN+S72GXy0CxpxsEtspEQxUtvjBMdA4AOO3EYGzznCusS3ddGFFXN
IPktTwGo/CoDBBOYZqZxbyoWnU/stJ8+CTn+aBbI0svRUutqO4zKOB9JTcBgNBoXE77boboYdpWq
3AMNzQUpVV7iWsjs2k1gQj7rbFduGXIugt2VlXEDs2vppiKGHhKF4Se4UMDihwNYypO6Q/OD0L2Z
dA21BUfMVvaqdFLazpiqPN0zjuspHGifJrX+kraCTEn0QWA3iDENblq5yXdBXpEjukLtXMEC1g/T
CK1IPLa1w0MBjrjzBunL+x1A5KsH4CRQeBq5T7clq6jIYcRdXkN4evlE+voage9kxsIxVxNSeas8
2MyFE2x97ZaIi4RTXdx0kbgBdQtKxTnqoR/AtXFqL4mqnZZap0flaRdYmt1gEkAqBiLw6kRvbowH
5zA9Z3bjeZl8QiaQBlmdFbKUDzyrZEOkb8asapptzOvQCjVxw06i6fq+UqdkEnr+rYfbPzylum10
skrLTx0V9F7F6koyB3YHMXqyE0VSIRmfZ8iWlBWC4kac7mqJKQKRDgYn/DJ5y4DA6anYZ9C09vbj
ecCTG4pXl3F5RRgnvQlwAvTT3Bw+UOPv7g0pHWlgTj36qjwwjBAlCpBcufjnIpLdGV6B7l7ehGNe
mWf/jaTtdprzebA9540IYqaSVVor0RhFjI+eqWX/IHm7aYLamuHKnn9aED9Dsss4FwMRuz9EwVMK
nv8MvN0+hhlnR+lwqreNlUMLXcMqM2eGqbA8TCuly8kemplC6JNyROwSjWRfUAUdthVNYkN+er2K
4r/HpXvTbdQAszbbBF0RMp/hbRy2afCvcdhujjNCm/riAtV9RtVeltdUwS5mCzKDHbRNawlDew7l
Z+PP6p5E2WB8kvuG2DEi27S+Nkmwj4QFmzcp05lW8SLQV7uvjChduhQgMLOuaPjw+2njOd4tfJbQ
sWgqLbeJjntm0V+c7yDRlpXIPLZmtp+Y7CizrFDwTFlixVKmuSKqRgvAFSkE29unJxUQsa6VIWxj
nVGqJtHV+mzo+vYYxwMyFI6sGtmgzzmNttcSaakkq2fN3Io9bc0SV27yt9flKukGpG8l/crdBX1u
TkGhB0psDv293miC8PAQt155HF89QfQ16u29JUIMaQGR0Ux9g3Re1oGX3K3C4UY8pY6/fzKzBLat
kAsqzzPCrdLylDx/6zG4vLUBs/e9CYht0/qED14o7GCKpIqjGV5SNwVzPvKvKe7ONr+Y4HS0fN1H
Zeba5tmuXn+juEp62rI1rIJle/I3b8BEKXV/TokV9/JKBt6azrcGL4K2pDBVSOxM9Wt0XDOoxsMd
OrGGfHOBdtbnrfqbWQUqjSkTYaAh2m0ZgTrIOZfQlbVAVokAdzKHO0QRpLMEIBYCT69aKQBxYsYd
Ap5n0o53yhMzNx0No/RK9Jcf786QK3rt2ItJN6DL3lroIpKpHSTKWBN4wZj7fqgDyB5JaDPWQwkV
0dzPZ7T4eWZ3FkSshC5bgjfL867bdHVWvOkPmMvH8d/qf/2cHRdL9dB6XGQ2pcriuHoWNyQsJvxm
BTTmUbdWdC+1JmWkDNVVv+bITMFjDzaG7v4AN/pHftf3r89mC9oAvfY78wa9w6ukqRB4QrP14W6N
QDSoEyIcWfF/bFV4EHXVejpNuIVxuv3SJX3a1uNXwCx/oKcu5RraTv9TFm6QObaPnP6wlaY2diDT
GLsqKEZUiAbW+HTNjcyLrR85TjaqrEIgIuR99O5n/LpfOJIObgFI4qpZbY075O8Uop8mwTaHYa2m
JIOsE2dFm6so5VndFpRdDgxPsaH0hHvOG12PHFRIBHd0ae/XaqFddWSxez8jOdBtA/Vp461pHxOf
P0aFO1zK1e3J2s0p/l5GXpuO7YK5UntamCyAxr0rjrMCMV2N2kjLnw04LSc1L3q8aFH4W8/h19SN
Zy7Ih9XqqHe1VSSetqIcJWrNR0/4fQez24UpXfR5FUINbpYsYxvZZjRDitS8ob8QlmnR5Y+oof9R
5h17OmmPm3L78jnXe/1HB1cRW4XnqpviewH8fZKXBjaHKuBZ/kxJPJ9RTU3ZBF6I5gXhVHn1ODgm
57imERNLCrXPrP7XCJum5cYubhRRYbXBO88exG7nCrFcpQE2/2CsDl3ht8Rq8UogIRdozkg4P8Fj
BouPeYIYO7zM9uAdoJshR2BV3r7h9dmQ12ycean2TJKJhc6mxcUgxrq6xurvJaPv3ihA6GXmmK1P
JR3ghxbQgsYqxIjWI8JRV+boEfyqGqbF1l/tG+1yivIE/fyjkXkGEYEzR3i8FKo3mnn8nJj52ox6
lRQ4qfOlbVlXHD6w1kOioP8c5o/LbE+zh/Gxwpu80/NBn9VGPMntdcX6p22swzBTvAMtg82u+51w
66WeYY1OT2+6E77Req5UyrXO9U/b3za0Jq3cVUTNEjKUyWL1wW+3Jiu1kQFmX/HsCXfo5piB+SPJ
G7GQA7WN52U89YccE3xRZHlUcWzzI4+EXiT+FjG9glouJEP/CrM3jFxPtN13Ow+8lHm4zRefwCJE
/vWk+suwZYcYf1NtmI3sJeaZRjCqjQ83to3+QkqKqlORmncbKSCSBtzNoaYJo9UaNGL6jBgw87AA
4X0RhsA+V37DaoFhqcCvfcfvyopglWYhvq9w5qyjt8GeyO4mvIEOGjUVgJCz6Y99eHr7gnIDZKBt
Jh+quKCGSkn3xzVDndIosodKif7QwyXADT24o3GVt8NydpUChoCubWCGiL6kGWNxdx6WZW8klqXn
OzhXCTa3mRmBBWv2n/H+mRYbK4n2qAJ8xfsq4BndCcFxF+3JIRMgRRbV2b6oUCxsZhpGnvlQ5gY3
mf420WYhzKClmUPmDTro3KjMlEZXKkWoy/PqpwcGGCmmhX9S5QaGlJIsVnwOsYRX8gKEapJjwS+c
xgZ/oWx/CJkBtYr736GmCHxSpGJAcTNIbIzVDY+VLGnJjzQO0nRI2joSeOP49nXHa1JZxqaTlz8o
mYTc8qxziiQrZEG9kWj4xoEbYrNf2u2rCWwMSLRLsvenccNskokMzjCsjvdkDw1yR2Fu94Ah+WoJ
Xlun0eDAJPgVIIFLUWb5/6Yaz7gyZW0OYAKq9HRPxX1/t2eTtKuyNxCM2ON2vafBYHdjrorLA1C1
NhIHpgx7zQJiWRMXAnKfpfvuSnOuwGC6/2UXPqf0J35GUHeJxInTqMjCkTXsS2+AnHA8CVfcQiO8
5DyoIVsFaKgwhEp4ASR9BRq+YtclBN2rmQ2J9cSGt5T1XwDNcWZ5QBqIwMZbHEnLs+08WYI4vQfM
5DBTJwev+roMGY3UsFE/V//tRJn2KM/WW3ccbA0nwOWJINA6AX9gEBKQfPFCCDD9zmLMqXQiODxm
00hikvXISudRZ29uBCyLScqMyqqpTrXnea1275l88ZOIpUzv1YtJOtpzSlg6hb4gn1Uo3AXox6LJ
tA+xhZmTUTxCliTFIk7I/wfHQ0NkVjDiwe9mPKpq4HSZXDGpNjMuSwfuzZHGZBFyYWWowutcSKPA
bQ+Tet+vag3+qIDGjgX6sUoaKv2h7VyD7cuPxQVj1QNyNFDaKilx0g+JKzrTXAnrfOV8ZeIRh0q7
5MvlSTg0dAce1CsKEXH6sS5ofi4waE+ix2nMon8GEcMD/xUS5EpdnwNbmU57q/XH+Q4Qj0DVno2e
zdkiP8ojzqU+Tjs9rkFnfeUXHHlfCNoBbQJo5DLaSotsiQ0Bhz3r+5+9POQwKoMohSG1FQiTnjsM
K0jawJaJftkyzIOcgago2jOe63tWlO1qAd5XDoVsNEl94K35XSjoDp19HxQq4Yt5p1Cc1Wwrtgma
xcstc81AxVLVXei0GsdJHG/JhGQ36xpMGbgctPtmsCb0YF90+onCMsZ8h2eXE2ThItEER8bsLrj9
TWzgNirwPkBLKf8J16IidGNfiYF9ZOkW7yFJPGsDWsCGH9t4iizlC2bbGx0jQV97CZ9Up98vqwDP
CXTrXN0ufDGJhI50cghdsA47+sOQd7BZVMXTcXSMDf7YeZqwgBspzCUNGS5g74HrSWvJ4PVi6fYC
UMBS7V12aOZpUA43TjeeR5JhwWKC5jCHKH47Xtqi/DB2AS+gnp3FFfDiAM2+5jPPEgBjxP1imClm
vaU8MUXMpu6vKZd26D9VctvY1fVzpIPXoq4rUGuSvAX+W5RnKmQhzTk5KVazupPCO2Pvb5zeSSvD
ntxp7jDFV2IsvL2TNcHbSBk+oUc0a9fsh5GiqsGk0k+tFQXjYzUIiPkypuC0YDOWUv/7M2dIXEOj
iXD+fgRDoLu7kfKPmKsy9WcKsgJ780ugTvTubjm1bt5/iuSzsGuw8UZSTQZaitSOw+Dj9lbNrwbC
SUooXd5PwvooJYPe1KorB8OqrGsZ+7WtQYQ+aS/Js9Jll2292JJPPpR8dW1seCK61FdIHzxJoyqa
h3ePO92e1td/QGSUIj2anJqvyccMqAbY3/B/SoCa7j0AVESAAI6i9t+JLMxBoPb8sId+L2MHuJCd
O1/eICe+fJeEZZw5khHoY5n0CIKn+Sxj56Hp3dcpI/3yBni1shZ3ijj4elhJBcRK+Vz6mZ3nRreb
1nIt0set8KlWI8IllPWbFEpSk3q3w3auvFTYTsO/LZcBDc9eE029qVWUIv3WDRC9NaxgNYQrrgwZ
M5dasywVFsfioEc6YXsEQIgiV+o4LQpoDx9XTrehkFF21wGpiWMIOvbHBtnvkKNFE27v9l8LrC7U
YsglHG24IdQWJa5lMxit0HSFttUJHGVmoK+sCqfaGAs7zaefkmyOfGJ0azM2Ap3eOmfCAOSkGZ2R
ltlQdutRr2qTzGN3+aaWtMwistK+ibBURNa8qUI/d6GaLj+zL1+wbyQHziRZoO2rtSx8akJlxJ2J
JutUrCytnF+/vRRegxS4Wp6SZc3cTNoPsjdeULsjSI58keuVSNlWIvcYJO8v9EvZtElyetw/1wxe
GI4QyHd+SQDSf/YhrjHT52CWh0hs0BdftIChi0NaBRcjozME3idJ7nK8h/vuJG6IK7N3gRn9+yBo
70W01qe99lWqM/Wh3RrelJK/3QmAefBGt09xQR+X8cnmzvsL/ji1N1yR7QOU46DvgpDv1rFR+9Kc
n1+7vK6TV61Yq9ZdTA+0eqZufmFGxmhOBNE7PBp4Pv4igvJGjERL+c5I2/sVW8glc208fHNFIcVE
LHj3l6Ucrd3zK12CXrSh7CSwZ+VE7odCCYu6W9pzOxdvh0001O9GDpYqSHBSJvAnWwmCCvcckp5W
AkTKxArk93sOPlnyYK3v9jNPw3X3nwikbX1OXeOMJxXUahxIUOFYKS4F0jdffeLs9VkK6IgeRsYE
GqL44NlbJvXsc8bb2xMhrsmHITeaAA7rDLXE9uAN5GPWem8xf2vkV6ZIp7Y2X4aCQuusFVo1ROjG
Ft2NGiVxljkKyP7899nBIVQXvItAcESH9bNhPuGhgJAa/UhPgqv9+4x8msVuPhY5CPC5ChzNSxAG
ulUHvofZXcUROlFZsaEX+A3q+qVfM+OXTA234fukTtEBwi1dsoAWPj/df/a1WG6liAnrWL3b2K2g
Y3wOwUdIEBhPMEwcB5QGZPT39G8cfiUCsRCRMxJ1QROv5dcfJAtN7ICE6+7a/sMhtKc1MulgIPGQ
XI3xggLB/AOeujkowQP/87yXdghZZCUwwIsCNH5IPBTQ6e1jnS4Z1EXOGiHoHysUstyL8izF7AMR
kSbwwz+mUbR30F2rO1ylj3n68igg3s1E1StLpxcJNhlAoWsn6KjPOTPBYep4UhhZWljOl8AxvMTx
VFbQ2se/xZlf5Rg3WGbyUzLlnf06KzxfZNjg104D47n0B9M9JGur0zimY1zi8KVMk7/MYMwthj3P
3qlZhT4cU2kPnDYj0zMtzVYIcjetJAeGnbBfBKAjjlL95R0kWU0bkH0RTVbFsPq7MStLuSpBEXla
MxcgyXle9HqP4HK0YImihFok3DesnX2vPjrb6v6RSKKC53sGy/ZyECCo/1PF8DQ6+KcJr5Y/Xb1c
Jv+ftpzpXcIJfxNtWJsPN4gCpaDgAziipSuV/3Tm1AKoUgd2GSjC3VQCE+UN2MTYdliktte5mvAE
b5vIclWRExSie3tQuvUSPHMzSPZLhUIUshl+rxG+qmWtQbMcsNRc68BIER7IqdhZJdbpEYe2YfO3
saAj7iismVTr6QYJy3oFt7lKXbG8mEo33DmUv5gEWVNcB60RjtaVtg79XnBq44yGJgqk+23/3PKj
H3gixLIwDjgspOEdKW1UMnIRw/sz8KMzjutRll55pJnB9aXA03hfeyfJ/XcLGh6o4wBVh7x8i/Oj
DkXh9rswFBZcuvfwXjl8WtCv8/k0RC/1HwRGssl0eLl7anCVletys+TwnBM9J5WBL1l1zasRlf+B
6z3jX7iFVpQs+aBusDD7bMIVWFQEdcjWt2yHQcBJ21kqhcQefcqC9iiMZGaKXsbcsBVec6rTvQqq
q0R5o12Hn3iboVuF+L5JDAkXBZ140MT8KnrBHrLOZeeLsBfCwl1vAlcYTyzxlHq7YEBrokQOsmKj
AYCr/OoArMouMhuO7rb1oqAlbqxI2QEnq3gfhi4fsRneFuWNqPE7BjxaUzFw50Vh1MdCK43MZxxm
eT/bT/aCj3R+4M26KpNfS1RmKTTqFV8Du7fC6xTku7KLMmnQvFGuVF+yc68vsyvkCkmcOGZ+5VtT
VX7ccqXW8A/RNVoi+KW7MZoW3dZm2+rLzRNGgUrWeD9iYI3gWNq5QhurNkhc30QapjOO1pEJSJ35
4B5F4cjjbAaXfg3vcJNPlK58jwhxP7C4EYNf/gQw9fWvVfEZ19uA60H+VSZwuXq+fYnRp3p0tAtl
pMd0UNzhAhqo8lEMlnyU/vg9TsMwo66OFKYJjQeb5UHHFEoSB7q8whVuxu+c8CGrkuXpNy+7NQjZ
Jn6VysLPb9rs2wt8Paj7YA0+pxZc25joHzBjlB7U0yBWUVMgLwMlBe2gsseQi0h4GH3iDwK2FOf/
TYVT0osFuOWrHO43pkKEmFlVvLCwS3f/7hjf9ENDZeV/xJUd3nWgvyZivr7eXJCHBdAN6hYJWf+B
ewIHs5rH8G9kYQSvVvII/zBOco5q/0A7iHm4CqERy7oaWZ9t24jX+i4e8DRQgAoD6CMbwbrUbKcB
6388xK1UgeFy1HZ0O/5QVui2h5D4Wo/M1kzq00caPdTFQnqCddWZNJ4WPK1HkMrH+2CZy9Fme4kf
p8tUIRRofLWB/QTuFqKGBS+rSjoYhgdDSZ24vZXwbNOKSq5bKohj4p5gOffx1BOWZg0DL3skCdld
cyCTOVyH99IyZ1TfwhPf0ruOyXmdooCDvLMIm1ANKATuQ86qsumLc9G7SO2XNA1JXii9Q35iK6zR
mIkQj0GA+CP1ce6U8vrlegkityYH8bIcCknDvzctXmak/QWrb1yIttKKIWP/15OYgNUUUqQtJSzK
RDZn0U/nNuK/ZxQjdTGgyNWPgo1whryQy8HSVJo2ng7QcyYZye3JkpHwMuCdWmmfoi0ud/i8hQd+
rb3eRZ3DV9xMrSbQVEOtBax7OF05ILc66zebaVJRqJ8fM7/1zKNLm6mM8nG1p+lvp7W2ilcNk8Mp
ntMNNsstb8e0aZAVWEhInSISXB4jhfktWstuwQMx+5Cb6cT/vEqZvXwLnYVfTtAs4tkishhK1kYr
VA4KH863dyKR1cFngHmBkvxgRp7mJje7nNNXTu4A14VEUfnaxR0jr9Z8ji4AHC0scfoiMLmc67I+
Lm6rSWmb5By9HceogYmV+HA6GE7pQk6ey9f2NZXZvEhXK7kFYzUJV+dLm15zoh6aC9X1N9nexsb7
a9qa50d0NPThLcBtP5oEVskQIx4oDXfiZhi3YNQsBbc2n911zCZb/RS/lu06qAjKVu/4HvjYSO66
bTXaeD/72SsOjfuVunwQGWUMNWcdC2RAC/vBRmRJdNC117/XZPhxBUc7n8EWpKV6A9jE4PdggLvp
PBEjhxF8emoxz7SeT1ReK3nJZ+HMtiDE1di2D91YISbbHXsh0x/CuLjXEgYuBeftpCWexM2BqbOt
7UIR18sC0nOaAf2gqaEjlsvVhgAuSJmciels7sO5cRa7E4N8YBePiNp6MqR/Xd11hxUAVbisoiUU
9RmdPai6xPIXR8ZwI86RMxX5tTn+VN7KuGlOb2iwgmhEi4RWosYbmq9pq4RxWFv8w3gUz0+pyWGF
BHHAeIBHDAGGp7xpyUJxvaOgdIDRD9fDXhtQ0PnB66lPY2+1S3d2Rfm4kaGb5INN6Ri/92+gVjNf
ORLazhD6CY7EPLSa2AVxpwbWc8SeC9Uc3nInam0adL0CVowMcEF1YuOuL7feT+a0ZDrTtgUDDA4l
vCX19fG1YierTs51qCbeaY4ah6WFvek9kUXQ1/K1Kd7PH4YrRaXaf/ThtVGfixvfkIKfXyIg+Bvg
4vOM9jggHNkS89C+9mflqmx7X5knmtIy+btdmzJcYs3gR3uhUUXUl/QpQUAZkDr95wfELLJ28A3/
VadptVypLXSxwvWWMmnoC3w0Vz1hM+fX6oVbEEJp1RFuNUDdol/57p5C/S4os+guI8WRTUE+XpQu
CESCCGfN/k11b0cJBGHONqY2khXphL+gAjvy7OCtsYJyODK8Dn2GAnG4tf4Z02Q1bAD9azDJPvl+
LIKSmjktyfuGJE5MckH/9RwfdcUV5R8DgF2SDh4hmIAwMjyCfrLGpOG6T12BkwsHCV9DRw+p/g8Q
RiQdEvOOgR0WzGBgVNyQkOrRXIcbkYY6x0HcXoRShqUIGmHe42yKxMKCjjNo3tiiuSOVRShPxOV5
URP/3+y2G9xVK6bBI8ouC92Mti2GQU1yK3SJnQyUEDk4MB0dj1aJD/OZ8X+bLLUwKL3yssiTwkYI
FnTGqrlXv/ea3FgHoK7h+6vBQwnjkOrFjnEbls4V01B17YYpcsMk1GJ6x7JTBwLEn7jYHAjGkDyg
T+MQkOBJajc13MCkDm7EMYuB6dyyFifMuViKmGrxDivc9jnetKCq27w598AxRxhVV5tG+VzHQV77
bU1FNhpL9xiEhAcrxy0z5esZwOL0MjTZUFYS2G907PKtLopxTLtPtRSsM4uuwkvrYpxzLjTVBYDf
wuQVXEwRolNEMn8aUJ3zq87ru0Sk4Zp85WdVoiwly9+1IV89OLyEetI2nWVZMU220qyah0YVi2OJ
PpdmV8FHs6cV+/vSYzZ6q4WmGTv4IsR+GvjyWBJt1mfMiE5pMYk4YrkaoI0JrRzhzmgXuc1ap6dl
FpF2eCT/I1yMxJOdE+w9cNMvJqidnh0zTuea1UHfN9KYpDR4RyQR9MVcSHCGfklrbbJmZaklTxtg
BiANZkpqxqglEJuzSiY5TPSevStqvtsCSLtJDKcvd5kXinIpYxsr9TAPWniVY+mPJc5HCrhTEFlC
OwkT8N5bGlTxXnfR3ylx9iQbI0CaXKZvbva9yPt4nW5bt4t8ADMf7Fjd8nmmj2BM+T8qcP6p3lJl
n6OmSHJB493R7tsTyKBubEQW2DdfQUPumR5Kd6BLj0r6xNT0r3d9ZiB8O/5v2g7pi5HbiGP5D1WH
yJlCZ+jEuRFVdvMyApq+BRsWwGO5s8R5dZCx9Lw4FTgs2Cn3KXOsopXG16s4tMGazyhvEMUh+kNo
Zf4dR8igRJFrZHmZfAsP7rJSj8nlPnGy7Ew0meyX6W4jpUyMKsB6UW3oVpwVOeCqmlXCUwXZ2Qw1
5pJ06/l88lEa+F0ptD97fWRkAbJ490pX/inu0YAZ8EDswN+0aEO0dWCpywUKLDAW5RLGbBgR4kpx
+D/cQ4LoancxQ1lWGteyd5Qx+SxMboeLQrth4fZ7bB9DeX5luBCl3ods5an/HlWPOOC8EXOIRmYy
QMgCCyoQYdlTLmVZ0HWsKp6K7o53bMXr/DgqaiMoKNQNlZXzT0lshDb6k3IpICgU7jUlpqooj3ff
9uSM7zlxJLs6e1zvYJADvf8AEyRbvD7fnqp7RjYdlJQkq8QytggkLR92W7mm6dNpnrWLn7ERsmiN
YvQ+Y8PzTKfdo2prg5n9H1xE6zO4lsNmOT8D3VvoiQB0zb1EKS7dPj8ZE1BHNzAwYZLAKtUNBHBa
3ifh3+KCqHc5NkYrbojSKtbPN6vdseur3Nmrh99XyJ4C3ZhvUrQD90psxQ80VCafYyLfrmlD9lqk
ToYj1K+xtmyH+zwfu/su4zPcbMPR6w0u8eocgiPtZfY9uGE7/QdZ/hLsSnDJTmamFsrXDNi9mN//
JJ+QWTKIfgPJBhblTioa2xFgll0bvlRCzMe6vpvEVNBzbB20AeZ3GHU15mXYJFDulAH8SmYnDF68
hCTluZUJPI3/N9gMYilkePht9yeCU/d2J6wlXoRZs/jgQK4FeqTNhSeqDHd4/W4BWSVgMApOntB6
JLfyjmAjyDg6Q6o6d+BUCw47eZZrJ5BHONHWRhJOKMT3bBMqe8qUb0bAA2oxYLSsk/xjfcJQVKtT
3NFybWYHQWD/qjTypVBIsl+FjV2E8oC2UGi1RujB26SIaQpI9qyrylGu51YXX88Z8x8OUzYOx/Nc
crfSTDE++sudkAuy/64X2WwsGf/cZ8UpDyr38k/NixCVyx5S9gf5Rxvhn3BL0hupTpBi/myRAs6X
CZkqjmXrzSwJDrgt1sgu2eteV0CM/S135+Jhd66wS2qDdDjaTqORJDSuQzylXpEJKrA3+n1sKnDA
p/lV/ToVJT0X7HPZo+VSHddegYX0HO6eD+ZHrSXC7hk+eyqRWZ0rkIGqFx8WGqbOWa6aLd5OCK5/
uFr3nlPM601qxDUMvImbl+qVYwC61O4NqY8vPm8hIHpxOBlClNlAFmjgn9OtJAP0CcKjtn3TO0pO
pe2XIvSbzeJXmfDKlXAVWDd60B8DNeqD+sW6RIRfybewNbDllfQw4swEmWM3dE3NLc+zeVp/Hb5m
6qas8buUO/KiVDKh9qlFU4LSfrai7sNNTzuIxXO3TUsnmLQ4Rst4wDcrvNsxR347j0eKUOgoHwcy
rVObDQiU2Sgi3pqIUsYFteO2virjdZ82ziQbwGuVt6CANo3gccx3dZ7skE7a6AH3b2kKm89sUbvU
nEHDMxKz1UhuFVbtCO+ReR4DwqVfjK94yGJGKnlKKMnVpSX2qz5dSRw/eDE/n5lFEURrp6I25hTZ
tFFoajrVSvN+12OwhyoIuOufE+lrTmsTEOTHNKrGI8+EORN0f2vKUyVYmNolrb0Qo8/FUGC43v+Q
XIM/yWKpcdqm0fli9PjSNmAitm0Qimr1voAARaKVyjWeYE4eACV3R9xTWUHL/W1num3yh7QFOvKU
7ntlqtfifwmaD1XNukJjoW9psNZj5zgfaxoHFi09xTinK80ztK8Ldh7PVLepK9/IVvfC5dvTejVE
xZoEJU/vSIcJLphk00gzFixl+Gs4O/ULH9jhbu2SVKAnq/UN+LzdXg+91bVp9yesuMtIichjLew4
AVMnZ+Djwqc5AQx5vyUaK0SSPMORVdiK2LQPKhyMIrHOVIMcFRNVER9AaUH6YWVjaeJzgE+hyVMp
JM3/OXnu2bfP6m3Rl06R6qhhnYuZ6vIr8nOf7yowJHzC81DSvY7A23AW7zhafwAGiRALAbE/MmcY
MFRXjZynhultSt7y7ek5m2yDd7zbRKJqs4zRWPi00TWqqlv/g+triUr7n6hRuU/wlV5U9GCeVvon
fM5qO32+po80GmY/pQ/LxvKWn1DGs8k6rDDTz9Rb9pYEc1xLlem10oUOdWWcVG8pDoENqi7d6VfX
H0ZEr6NYoGwsyx0JPP7KRObjm5p3BR+nx+/owm24/W6xC23pfVDOnn93LiOodEN4AD6VlThG40KY
5rzsd74K6QYf8BctKNngtKFuiDdsMxtTpzZPmFe6VLIx+QMfjU2C+FJ+fHCGnw+Qi9CaR+2KVRXz
+UI5uxopo3Bz5aY9B4uIL4xa7ibrGHAE+7S/6R4TwZOp1fqN6rdYTOyjGZnn16lTqkbKYiDpxOW0
1Qjm6H8MLPKoAfrtcNkViyGIpQ/xMhbsfMyV+tfXxJUolE07+3C0Is0R4co7keg71yggQbpvB1Gu
pC85QUd5w+UBaQ4icsHSj8XQMWfTyOjcvzkiIkI9nLkoDW4uthnd95gGES6yAvXZ2wtLohCJiuQT
ZkwdDf2vevAyiL31NrfemxsPRjrhBKiAkfJrB2Tf0A0CcHPl5g9XuYlkIMLlFlu0WEWnDMSQ8oo8
1slHIcvgD7XCqf01mL9RnHqw0OkyiagS359VgYMm1O+6UqAwBSDPf/t5Srs7oOMyp/1K3w4k0Tht
X3/LvhEEuDTua8hukx80xNmu/SmEQhitRfrQprCOXISvPSdCzchYBdUw704SXoIrs8o1Vfx8vjMS
me/6R/9eXPOg5mT2S75PNOQswTFc71Pui53tzQw09PujBc/xLv4/le7aircFTbB9FbPNVJBPwTCm
wrt4ls9nM/TII0Jf5TpZcbUPd4plGP36fXFkMG2CV8SwlOdIjOKkqhfX+SPncWuksQ927uOPb1ks
hX1Y4QpNWJfPE3ptqlHJKqTOP1u+N6szMaE2Q6H9XirblZCQflonFCsbFXkteQS2WTSBnHif8HDR
ciBVIA51+KWPpme1uiko/fN2lfF4MxC81gsb7g3TV76xjMV0xgyioVshuXHUoZQ+h9hG6lLZ4pLF
ZO1UZqay8HynqdqccqIvzsFF3axIbWyWM0zHe+Q5PIGhOHyCL0xRI2uZxS6RzCyQb0b7wHpx0JNg
IdRSgK+cH7OIMwUNKvYgzofYpL9PQ4Gnn9rD5lF+GX9r9lo+sPDyO3FGqnd+QBk2LiEi8Kzc33MW
VSUIPkMOHlsjTiMUVG7xxKSaHc38JJI3X3Q/awtA/ApQZA+uoMNm5zLggl2sRcuIbeP3q7WnEjja
FW/tUhiF14WKEGmn5zgcsXJnfAsM7ABafr2Qjuvf0aPjmH+tJ5ljZIUBXyDiqZcOVT936C+QxHlN
I7eENmvGcmXm8nDC8aU7PR9UaFWS+NIZd+C3s0CNw8byYu/tnjJFJdtd0XCLqb7jsg76lnJ+/NnB
cEhLo5MNtdU5ZvmSV9pIFlWbtzsc6KkstsPrKgp/xeO6p1b3P8KE1GCv3dFfil0aPJLrbcYQAX9y
As0VhTOL+aCkWIqAB7THeQCpVqfrTvenDORaKS6jzga8LpygbkWxnnJpmX/wtmIjPs8YHe0mYm0j
YzBeOo3P/xr3BPPnpXZx2cC2YfgeRbSrv/YD8WNrYW28mEhtui/halHsUXvzAFKx78dTBBKex9Uf
+yDqugSt0NniDnWOeZgwdglnA3//uHimJCzNoNLG1Pt3uICcIccgJ+NtwZDWjXFKkPgSLookugeU
LsC1jloK6cbZjh/GBtcQGyKusdRHvFA9JhmzNyDSIUXA/oGdfziXDM6ThuhoUrK2T01HrpBptcNb
LVrNaAZPPLkJcwEAK+Osg6uNOSkNkEvh2CQ++uM3LCzhJSTocasg+8BWedExecIeltUrsjn+K9T2
VVznWefdMBgTwOk5E0UPm9HcN6/24vNpUZufD8FBJk1oBpLsYztnMTWGAVQ6JGDrq491qhadbpoU
ADdf9ADwHq9ROrJfQZyEQHTGXt71aV5+yxmxhj7USMiD/l1W8gx7FN1u8FlRG8hMDvWtp50637RA
GUxH6QrvsL27MDFS/fjAJ+4q6zdIn7wf37miS7au+blcwf83KSFiBrtWNZ8GWFBOmV+nxPsqHf6v
8xmoVtUb7b7cgoDGzQZUkKWI4Plsxp5GTpv0UAmBM35O9vHEuZCMe5boqNp01mciJIm+SfvxGnSV
PjcIOJlU67Wkkpxf21IkMibRH4rHoZ541SWf2pGQFjMMNP43RjbkUKiNxaIPN1ueIK62D0QOgEnT
xFcJZKHYB2Mug6jYSyMPkvH5eQE9ZmjD0hh/KIw2o3uuLuZBnHTVFOmKamCWW32UXwaYLMGQO6Nr
d0alw96XmWYciSIt+IAxI/jtQhiqXaxiaS0O2Md1qCrxVos+2ORbzln/hvKPCIYINsQx4pBovrqZ
OMM2wMC6xEDRPOOg0gcoyMDpxAe/LrY9AcsMkm1lkgP1C3MctdsNHejcYIeHy4NFKhgMlsfYramE
6o9CLcjWooA4MG6Omw6x2GQwLXnpXhALxIcp93gnECDRfJ0WijbBCVJAiJul6qHJk/OZyiFoTmZ4
Gg/tnTfcPdoF62Kz/fE8j+PudlWUojB2Uk+Ka9if4f+PazyNpQqnDIBeApWJXe746oic6k/FxgFU
zOOC+tD3hn6oGP+rwq/Kxts84Abhe0F6i0a09QxH0VYjgkqVQXg47pEu+DKTdW1KL/IMDJp48VWe
0jBOhnUb6h7G4dvPdgfh1d71ZYR7I37cOePjOZKOauiAddZh1B7ZGZpx2D7J/erWRjfVTE+W2zuQ
Sc2e1a1ZSZCgEuvV6PGapuSfRq5QHgRrIwt44oAsOTkQPwgrLqUBUHtXcBepOWRWqmbFlszpD1o5
xlb6kNvC67D5mjWWZ00qcg9WkyPptoJEY1rK1pfNKp0nNTEefGfkl+SJ+ywH3opWCdQLmTjJFfbe
FgmMe4D60vW6fXxOvXlc9dVI8u7zL4vOqgkBKOV90lk9QI/zBDC5XYSioS5tuPCRSQ8KHhj233ja
2na/yCnwkx1Ba/RTV8ruR7gJw4XfTxPb3WkJTL1EVT+1hPpqVFWNpK7oaSmwVe/cWLXjFDX79lHU
b/1DeaKqUTxEtWagveVdAzxC3INqiL82BLRLnuiHX+MxtAR2aLNKekaPZuPAxiiMxEa4WDV+Jkv5
fXS/rq68ylFnz8fBwO23K31DzkgMWBJ4wkMwoDe7YBZOllOv63dS1rqwRlsF9NypHf58QBF9uMo2
xT0gsZm/XaqDShRRlEQWGO2Q0wofR2HJRtdH5SF6ijUkP7+sf9cR2hDTnKlzdrSms6JnUQSDQFrQ
YxChW9XCzZ9Qe/Td7kGCSgeGN0fXb+56u4bRVynWh0xg+ZYp3xS04zwm5FRZ7ejFKn5UX82IxTUj
Z47F0V2CfkF2OE54G5IU7KdgOL5oJZfuuCEstubFzo0DmT3EdcSigU2AB5Hrw4lKDGYg+sGpNWhr
K71g0PPUhAVeGQlSO09v+Uy6PSCMaGOsi4xPApjy0YMa/AOaEA3OS9+ux5wZ5pMPY0uTTzdHEa64
sYoIwbi17ie5zbul0N19QyeWNTMt+VA2+Hr2pf5XqiP/YbfPupQb5ZXJSMZbbhteMT9Dg4ZMitYl
Wk949lRVooDtD5yhzy/wdceOg+pduJLVOe3Z3Eow/fsObD/Vw7Z4t8eCI6n5PnPd2H5LmS4NsAOq
quiCxUWjBhhGzwEDB3dr4krIil2W1tcdjojDiN1mPeE9j3wFjHaghsr2g1dYIz3BcRiBNJ1mHty9
A26IQUG7GSdvtktby1gKsLckQXYjgACF3i6OaHuKvMp4GkdNbZv4nmfA5nqDgfGhSPJEPHwROl9O
+sHxEuuNl+veAqRg6GF4dMgTfm9YXlxPPIajfF02rc65mxg5fih/uxJz/BbxUT8/PPpUHXOA0Fod
UXL+TGL9LHavWUSBBZ7OdJEUoN5ZScQGmvPX6aXLt6FsB88idpJDr6SWitqsb+gwVCcJtwS6c+Pw
GoFOlvV/u2XxdThsWdh2WEvHBGzxLrZnGftyoUio0Ij8AlwrYUx9qWgdE2CfG0WDgcXBqT2TOnVk
tSWh/JYM/A/uyJ10z8FKmLqlVdFp5KZaPFgaqZbHSTIWpDMYjEnQobQpzoYAnfwMARR2jJ/hmPy2
YuWPOKCkMe6GNh0lDAAhvnqaJlE0Ju4b2XVJZ7bPttF70m8UrhenLD2aNYqIRoVzHExqvgwrKnE8
3Ga5nJR5qcZaM8eUtPNi3Bk1eg9BaTnYhfhS+SLm9UVW99kFbpZGkSDM6+upLOHHeLhkW63nydEJ
oxmoZW2tYcixjXpVTZ5rQmzI4Y4ersTOujGF9elPIy5IJwN8oCiTrlByhcgoRWzTEzm5OQCd3C9r
n0bPq6riQzO8q34bEDasJjE/1KkD/PRhLJW8CHY1dp7LhDUhYg9m28C4/YSzWl7AG3aiak3Uu5/T
LEm4VxqRRzIvFExFM8ZQhHTouGcxbXD1lUJWpA4mc4ptGjtrxnvQPf3se3lywiO11OnetK/NnOQ1
3Q8Y2Rlzq4/OABMD1Wz6ld0B32+ShDHyejFpbQxfv1xQsDMGZSUzmf4KM7kLRWJeg0hpLPXj7BH8
E+0IRzK1EbFppxi2voEqxHQ42S9Kc1ePRzrF7RyHLiuHmIiv4VGfynL/Hu3enh5nm1QlsW7XoO2K
psMUyhc80xNTaLegaX/qI5ryq5msQlB2swdD04lprM20XYv5ypQFnjqp9J518HSGvqgDngyRwriO
2zI7LBaCCSxEGTH4DgjykJvp4nPadXipgv+aTOKhTKCXDU+6q5/ey+PZI5bhZXKzDvH4ZcoNdEaZ
jkD2Z/bboR9NNJU6Yk6wUYtkzcXgIOu9XfpEiEFydhJWnvuE+VE2a0Unnng7UbrxBuV2MKODFBA6
gVplCqd+gkjpL7DCzuJShstAZwzNsBB1kylTXMdLx62yAMioiPiXg1KSMLx2KlbdW5XK/cHuE2+Z
PM8HCJ1y7XL/lSzI0B/Pizshb5i8v6b/ueb54uZHtc8wJnnPeVuUDfBua5ml4JI538yo56Tzs1K1
+liC+BsQGMdaaaQaFEgJ7gwTyfi566JQJAESjeDz66Teg+d1KUUbZULS2VreJY2jgUr32kKS6xpY
kK48TIJZtIBgYLDE7I1bA3hJmnsLTe4SgSjKKZccw/i/BvOFVoEvrNxpJ2Ug9YbMpajJIsOInHvd
mvfyiXwCQrVoe0iDvacDIJ29SXXVFqQQOU8N1lrFvZLm+IZO/CAQQ4DCJeBfCjwpHSx/iE0B/93G
ihmmrqXv6cmTQ9yB1BAWS2RFiqagzfaYiHeKkF5AvB5hQEhQum4/TncLTdnKWmgLXvdCbD/h3bWh
Xq4jYkYKifu7CIXa8H1tCku6TQUv2zQh/sKVmtFDwCDjA7rEzKCE0IW6XdihFQhgwZfbhZkKirHy
QBDytGdDxhrGpmKojS8b2hhQszsUK4JJzA2vnqeBdU1QdFwXxd2E8vFJqThYGQ6G8MfMB90g5DzA
FpmT27y9FIfYsx9ixZIvOxKNsuVeoufLOdJQrQQNmuv3AF+NMF9FVwga5EXxVFV0ladlXfxfwiEM
fKaY80Q84U3rE4vJ9x4bLRBXM3OaAmTawowZYbUpG0vM6JZ2wr0VleMuk+VZQzKkRbv0ief66hMv
JIHgqoNs11U9pBtKVzs8j/QnsvwutgSMMBBuAkvSADETn4kY8aqDbfOCo3afJ8gg+yZyuzr4zxu3
/vN5eEw+QHDJI8CTEf9zVzOqPt8Aoi1MJgxL4/iiLVvUdvdpziJxlXsQc7v0TGFn90lLUQYn8oSX
Cc5S5fchXDUCVD2uBTRtzG9XhU0O2F/0YkVkEDyC+ct+o9txB+fzV7b6lfwMSrXifceljaw0ON5+
wriqa/8z9gvfZc6uks9kebsFpmcalsx3ayWVGZHyq53iBBP+wHNNzsMZlNc6K2Zg9qsrBHqZlM4r
fTCdx2K0H5QehFBGFjIJZQVPH3e8VidSEaDukWY9yShP8x3SDYrd7Thr+famstCqx2uaolATwzfq
cn01yB3LMrkDF74uOscZl6Dpote1t0uGWpTz/1MvxzNS9eLSNS7KU8AQPUhbqFxQgmc7s/L6V92S
b1mkXpujZzoPLE0uq/2lBPqSY5NTYjrbvPm6dVqfqtiL/3rP1xrOlB53rROzxuK43v2p4HKJ3nsK
HbBhLgrDDXifnYZUTnttXkRyhkWtZZCYQK3gusU37GNPl12WMujd5mtvtA56HtIucPEL9KEjDWbm
GIA36imOmqDT7Idb2EdcYbh+VwQBufk088saZGaXweQAfIYNevMrduJeZ1mxP9JAlrvIJMCzQyo9
lgKrdDn6a71glC6u6EBocG9OfXuJwuhN0c2NJAMbThGFNTrfcK41dbUPJdZBq0lewS5ALi31lS+d
6LVpZv6bMsuc/FceaF2/9DYF86UTXJlovx8x6m13UyJ0RFL8j4Lw5idFbm5FhvxEXO3tIU5rArRR
nJjAqldeizgRAA3nFur0Eus/c5ZHjFabGbuFUxCbM341wDQ6zDy9S9rZP8NljOJe8Cbzfml736qy
CKHzkoWLqF8cj3yRhw6Qw5QM91G5bQxmgGZqhF9Y6uw+D+c0/Vyk6NnoryH5uc8NvsMUHMtvBDHT
PgmbZ/9ikkQBXp7PchcsL1H+sq0gApNLq+rHoWLMXJGAVQ6YDnGOSmvoPYYvs/jiCoK1HqNMjbmU
zCMjN10wViYRiVoBS184WcUTpMD/bj8PZDJPLRnhLg1KSLRQGwI5/nzZlNTryOdc4iSTuETN9TlY
Ctc3PqG7YeLQc8UUd4Pk9HptJ87lTH5iZPTSiJ6A94LAq3h7X56uaFERIGATeNWWRyKGMpQbtB70
QdgRZVB/zYxR5hhVPrCr4PXEdeQKQnm5jS8UtFuRVrmcOgYJH7OOaRteWXYpikAH1Q8A1ecMVHX7
Y/rYClnyR8MhevZxVT2SXgyKOGROxQzIHJk8c19WSHzTDO7Vzo9VB6tIS+G3dZivaQqb5RrwKOia
+IEzSUNt0nHm3Kt6KNS+9p0yxg8TbAI3AdLvhnXfxXhKolsT32nBZBeNdkuTdzSZYbjJ7DQZD+9y
c0AOGGHBJgw10RU9+CV11kxfPebKnE9GFeR2weE/hW+W/PUKvBlb99eqL5CAVETwO3KbH+rS3HgJ
lbgQBg/of4kKFyX7VDSlbWBJrZrksuRNsDk8y+vmlzEqoIEZIPyMPu8S9jBciyq8TQxjdb5fKWVP
+iIYrCDDUysC1bTzHHKJ2pW5IbDOjjU9AxbGUNbT/EJHnD7u9sERKxyLTTycYtv2NidpEZqSaoPq
eiL+cd/b1m898IdEHrjxULxEnEkrw37EEQUA0GcFx3PylHGoqEIQKV8tBpkg/uQ09+8yC/vTo0lp
5DzoCci+cQz1b+Pw1n76P96BFVdHjqVrZApMMk0y4CA/mo+Iu+wpLpvCcmPzbEQTnKfMvJDsjMBb
6jSugrQp8D5uLug8cQZA3Sb6DcvJlRcKfplmo6jZZSsl1DldQ9nCrNAD/rcCitjj6eHfA8ucUdwp
vQr+k1VoqSYQ0YeBxHpKS3W9qe92laG6rPCa2Fzj010MLtkz0D4Ff6kLeV3dXqsbeTouLb3tgujF
LE4WPLavHSw0U3v8IFEhRW7aj96hMb3S/t+BSkRrSA26hjFijy7SqtmOdspRHzdpQcahKZm3O1To
mEK4qJdOIItPgoEQg3k8fq61xHVpitn2JfHUWw8dJ/3FYEXHhkWucl5/vszWJT45R4vioGqLgOjQ
Mj7hqDm1Y8VTDUdtQG8FhbosADnEVOZ9D+Zdr9ZitZ2PtKKuQ4wVSLZiSfZgcrxweZpSCbYjKkkn
LctRQ1yu/Onfx9LXeLK4/rKZpdTuFMoMjHhD7trrFQ9g/XBdmR3uc/ry6npQpd2U7WiwWSPZr/PA
KnQKC42Y8qQls2qcA38hLnbmrdNWj7eBqgaXs9RPMofBwizI5D1ARwQUDGFWCMc7GtDAbirvFyEY
eCTs4l9XLqGLLXGWI4Sd5vQeUk9imy1ec4hNtugvHu8DMvofbysat8Vh7o5l5YvGw13+YUai7bW/
8B/LkzF47rPcGGnrs1cdytGcRvcJSOntBqVIhAoih7H0TcHJPB5TMeVGo4Jv92W2UGwWSXeQ3Ufx
LhCrBmNu9dt1iHpr4KVB1Kv417B7VTgWUjmHE2XeAwPj9MlO1Qh6s2q+YVLqZfyIvNwVRhkBPa1l
aIOzCdtLkFpiB13Ep5Noma5JxczzwUuyEFj5B1pbBnGhuomw3ktJMzkFUGQIQnI0NbtfzhjyY9O5
mk2ADy9vMJzKj2WcmCCJRYS/1lI6EBQpHp/tq6Gq7AQEWbrVkWDnO5IGzliNcPMEkbTpzt8bvbRD
t8BeLWz14BsdRfq484uS2WFRasPzkoIV0Tr6Cq5GYNae6oLybQo8dsHaUyatlyZY9VC9s+TPwtlR
SVS231q3TFcOLPgxTbnYnJmxLgzDrOCJ6fKDM9T5SWODN7dGlzSIeOG60u8JjBP6dquJJviynhHl
0ZZK1riBbWL6p6sw26j0YSsIHWJkfsb4azn/kh2q+5sXKr7qnTEfNT6xPgT0LZKHAMV1Gcra6oeM
KsCZyGQAIMcXTbPQVfJhIdPJ3MdlOQa7rvl8ngACoguSvMlqLS8vgpyzlj82xqgOrWvK0T8UWRIz
9/Oex8Z0pCqCex+GzedPojgJYwKfPBkZ3rRfJgll0IOwoyeqzIQHhdeQj1r2CWQ/BmvBXIEDnuZq
xF+UziuPW+ppuWDWpIDvMotlAz6ZcUioq7RzH5oXvWt2QGjoZWJRldH0cfIODR0HJhp9xrjEDFOq
t2pwqdFDxwIUtOJJksq/UGyb69jhMpwzlGiinx7Nx5rhAXPDSrjKmAhJPUxZguchyVHN3uTUn2ff
ip+caD9VEwu56niMefJVU7bcP6mXUH+s9xCuC9uVOUE34WC1LOhyOTvHOGckHErvev/rhlV8eTHd
OcxFVyHSzBcq23BjyeYUGdEKa+WUu2V1exeGKWAw5g8fdniZhyqwuHyI3iP1wE9j9ThXDLY+rFdY
ai4PvsUUVMpkZF+TG6h6uH5QPeMXDV3zTeTE0gj/mxuObvTeRCRkC1jCxc9yEQipalU2IXlGNA9n
WYeIyLPRv4mm8bQa8UJPgbUUNsmKV39yjQ0HRhnXJdaa4DiG+fu9BYyebtvhKkK3SPPigqtXn0QM
pEPCakR1lETZ4V+JmtZlSBrLk5v8SieS6fm0NyN6U0PVDzmYEtNdYRIizvEP+QGIYwwW6/Sb1hEm
1WMW26WanRJQxGhOQrqd5UgNgISk6w8fnJqFSzUqyQ2dduIxTQjR//SaRN90x+oi2AiVi7emwBXS
cqlgc9E4Kecm6san2pNtLI258oL2KVHpsawcZ23sd/hJKkDPTHfwmiHUdL9cvN5t1LcGvj9nYsrW
fNFuCjCUqppjFpOsGqh5/CPMpAAhsg1l51r+LZS8sC9kmzKubj1V1HUOystHvv+V4dEJC236/8yX
jTtRlUwQeLAPjAKEtMpwt9/X0IZchrnGJ9yram4QZNZ8Xa0I6rPsCr8kdOmQutxSG7EOPbbiNHaE
PGl+1EYBOSiHpPTiYGIQh21lXQbIXTCibOgZukeaO00ejLKIhp6b79hcnfzkYQj5SsW/qJ1lWzQw
0M3A3mKnreWDGD+JySVsHEOxuSYyn0B6O0YTi+3l/leBBulmzGlnwGqa2gxOGY2Tf2Ar1zW+2WiF
+AxMJGMQVAF4w+UNcAV626VBM2XCx6WJW7rAN9rQav6lEQ1MKA3DvDmwK8F1cybyMzpJDhqH5ZsD
IAK3CEeP8L7lP+ZUXk9N1OTRMI9tl7dtzvFgorhhPwQ941My1TKyq+jh7ixEi8ANQJIZe0QIIYz0
5URTQ53U67SkoLA7F6YwJGOgEEOJ97+322zrZqN4EZ814z5BdhEGxYuVXSa5QVjy/pO21ddOK6Jq
4kXVwLUUuGi1vbp+p6rd4EidsXBu2jgEcrJew0hhu4pnpd8Ck/MKB2qaTn2Q2/lo79hmokWbsmk/
K0YjfdHQZAr02QkjBFInMfLa6lj58UOjSQ8bWulVrwc/vLLDw6N6r4YgDnEI370lcOCSORZrH8pe
ayQA7NR66v0h4Uo2N2vBwv5lTj4ikWCJCWvwKAxIwtOiLWdjRp3Q6WpZNxkcgbMsolJYN4Ixp1nI
fHj+usEz5Wz6lS8D7Wvbv4mIDSEsF/qYIExLhfH201KTLv96ZWZX6WTbBV0Uahtn42D+tyDwVwAq
ppx2jR6IZyp/XtNkmC26Yo8mS1dEm83VP4WZ/xtrnh/TorfcFG2x+fJQI/D1L/rgaMRcA+rJtmyC
H4MO13+76i5Pf7NiqNruw2ym8HKawVIhF4bCqp5mTeFQUpgk3SxFUqOv6TUkLeME5E9EPS8vGJoQ
6kI4dQanCSFvlI2N3c75fXuzUwFF4tHQgkqIHfkB1PAbhi6UVWKKySC1fDo9uZKBChOcTqUCceoy
j6nVmFSkHSK3Mo+K4WeB2zNg7Mdz3QE8wjU38B3xPe78IDUoBITeto9d6Ar1ICpBFmGaBFk1TLXQ
NEfEvULi85aQOtorv+ohhh/JU9sCqGwoRaKMVCw4P37hJxTRmMufLzZoYfNlVwEF1nAQPAlECoeU
myMIprLxaa/CBpu67PJc4rRZFuf3mNd8jfrdGTsdYTpzZxnKv4no96UAEY1uEgk2gpKxlzPj9t/Q
3roK3z1v87xApSgtFaYZy+w322HiELU6FOoKwUA2VoJOMOKqT4/UY5AE6Cx7EWlv9uyEB0SVwZS/
V9s7A3KlRZr7l+3ATVBmUAziBr61cWx9aMw5eY1xVhwqxSD7o3RgNHh4wKGm4llgpAW9et/uKh3T
g1/85fwK1nFMyHP1TGj7rY+3UKzxl/cZeF0HLmSpATaMNhvQT+2zEu5xPDcUPs6R1a+5by12x9oq
b29ed2x5WUQ0CBvyYl1VUUyagvFzL2ehi4RK/lzef+DrBTYfKObhJHGTGor/TZNh/Pxv3ATd97Pf
3LJwoMkxQIzGqDZDtnwDYnqqm59anA3pID/hdPvoSbhNGaozDEq5DWD6Hc2vDAw41EmXtQOEdpC9
OByKfyVHpoQIN//r5Q4cYrT3TLRJ5LjmvWbiwcMMDMIl/GD3MkcG+yLPRchYA/nyPEne3bNbphLS
1ASHA6Ds9+V3RNVCs9KuwxLm+Bho9Q7dtab90492iIMduIs/wKQtQBJx3iChIyAikpL65IgoQ5Zc
u7Dq2V1qyOA2b36UHxv9ddLA+6pt26BdU4tG88EfIgVVNTkHjaKXTByp4698+0KTgsveyMXBEd2I
UkY31sY416b8ShTDERIkTCZzbGrhg64+W0BOZKwxMPaH09BpMCEF2v4WdT/zqKNyD9woVUufWf/e
0O4PmoHKu/66KsxI8Etzib9zusUJls5QqLs6hrM/CjtNk0ugcbC+RspOJ1MKRSMqoX4led59BkIJ
QEs9d3toB0USH3YgTQSLPOMeWQqLOrXdS+Lk90MXLNZpbXo0uTREGFNMdvk77gySvLwE8rHhal5A
5IlJWx1BYGBGJ+UedsdGks2QpCDXtJMqRxeamWQ7uWKhM0ge/ChKvcVWE3mfAgU0iP6EKYIji9dI
paRhs8MSg6PugLoSHw6YMt1IvrnkgkcHTjvPUWkwHEn+GJe1PMt5yK2tywdQSmdk5xKgH6X6UxRt
FPmp78mnKcGnxvVZBAy/zUi4hWn3PsC6qjdf5GEwDNtnJTyFHGXlpCMiEvr//w86UC9aPN9OIZld
ig5wZgwLJ+M/aszob5OI2ihO8uTI0iZCsqi0LcQ6mUZi3rUqkb/gcfCXbg0zlEC5F/VtcVYIndZJ
siX66Ym7HkO45LCWaHN4mcgIb12akGEMtV7rRJ09bq5SGnWkaPsvB+nvVDub+gaHArJ1kpxKp/QX
h4XWuFKElOGbTab+/8o9W8dx6DfYxXwiQpM6Ft+iE+TZcXRvWEtCSfiLx1ugIBSCk/f+0g9JGFCm
u9H5TdW4jLDY6/XmokOktc29bTsLG01xagveaJigFizJaaYDAXVtDl/QtltVZQjqotuf6kUcHBc9
Y3hrjiBGOAdlgUgNwHPI90j/bRzZ4IsoW+Oq+j3iUlHeqgzpdbogOFFEINYsqVUQRY/Tyga5F+D3
x/zZjhKOFU7R4JMUyMGS8L2FK5QwAm+Vyc0TAwMynm/HCpmOeIULyXSEJBs/TuVy6pak6z4k55em
uYm8pwyVa23/RBjNJn1jkRd9oWIb0wPTngmW/05MbBFRn1Jx59hF9EC3ozWE5wKSK0pmxhGz69gR
tzyxFKIgqPkgw6QR1r2YTox2byzJitEaKD6NIKzKlVb+0rq49pAMNxGGafc18E28KFy3Bbk8aIig
tmx+LoXft/90xYUOcXDlMEREyA16ipIn9Y0Wzqe5NYyyxs5qcg6YgxbzalIIFBx7EKSQtOTrVOWj
hDb0+wLuJ9Du4mJtPPnqfm1+7BnQQiSLRaK67MRxh0baTT5yr0llElZF8cc2QrX3+919/7nAJDF6
/j7/7Czo6NwHpmfr8d78trGFx4AoZWdhcePW8ylHbUFbYwFqV9GnBy2B1/LAni7KG3/fSQAu8rkv
QUp3L1jE9GFCUq0xHLO8bZpaQS4jPScLxmV00lb1ZYo7VZX70zori0A+uQMsM9/8SE/foLc7+Cmw
k3beeDgFgBFPHLL0Nk0f/CSU3J+hKEb6NRa/wf+O0fmNyeKR7EXEgfLcoGFoxUgHWdgqu+Dxf22u
CTy0Y5m49mJJApqFFCgKrL7ZLyzSLHYDfV8HP98aKp/sOyWuAXug1ecPWPnjJLls7eywPPfabGGF
EtX4EDPi/k+rLR7v9komjXEvxeQMB4ZfOhOjloWG+siqGCB8FQQ8zX66mGJ2eb3cHzw2xlzF3Y8c
/mHqRc8zKSdGY3qZ+dZplJp64wuUPvDITc9BqP6Bf5U0J/SDf40cZligYFkPhXuHNecRwfZq5Ub1
lV0E9S8Wzq+AaxEDPFDiIZORE4LRvnKvFrXHpr/UweJ08IXzXlOW+TKj+w7C1+oEgRFkYq1mMiEv
wXjELdG5plMGNcyjxsbaBBq3P0iKF2JBree087oxAGpgHQyOhb2GJCT6TUyKI+BBqXe6yZR3I2NP
SeGw85HaDfBPFVj1qG2Z2QD7V1j2v1snZ/7NOzFIK0d+VminwxaTfcc+d5fFZLYAR9FAj8b1L62d
cE5J1GtR9sQRvzC1nPYl4+AauELDTZ2FnXAX1uIXLB52kUdisx11addXISCFu5jMwQ7blw00jdH6
2XDaXXKAXljgZXcNV0tkbQpTtClf9JvuT+lff8ocOi7rR2AXaaVjaNVuLUTUJ20bOSP8pfcdZXa+
+vmTYmdsTD3Abbz61gGirfKX6vj3lp7UOobw2PoXfe0bgMIguczGk4SfzQ+QE1e/oPeAjjiZJWUM
1gEslV8fEweNN5VKjjNIagxGrY6JN2ntrjNZAFC4MEITIwVWKGRNE/aFNmCLCSxo4RIOFGlkJiiv
TxMLng10x2YGsCeY2TxoqfNYFe90WdspPUYonlFOWBlbLlpwoATthikEObJNq0yMli5uI/231Dmt
Wr7zUKGiJBb0OabH86ycNJ/IypjnlYBeA0voD5fbgzjqUCNXAYH4mdqvn1mY//kq4sJk17ZfX10t
UJAxbhqiTfrjqB2UuFFRhH0pFjYIj/1gpqBMMfQcEmO4CyjJMt5YET0jMQE9KdnI1lNRrt/FchhP
psZLVM2j23lz0VpAJJZze9Z8Xm7Mry0JpSnT/XeMTCCuB1Xh0B9BsKYyMDajz+/0Q7MNlnhSitDh
7PskF1MLu5YqFxvVdyhklspCYwAdM6M+AlEfdF3BDeB7tUowHzfdej4QH1gAiuxUChF1YiovS2XN
OQJnfcX31ML1Uc92xMNbKRDZ0dY2qaNNd6yH9OBGLEeNeVm21A45oy5balF1PKap1ya0PSZHesrg
+pzegQNJQsXJHZY7RuC+QptRSt7McMun9/Rix1Sr0WnC1jE4MTM2TNcL4QxQ4bsA+sXlEcMD0b5a
kIEvG7oxZbziqIxnS0C36LzinJVYpHksIqfgFrzRLOH9ai0cKG3QmGoU77+LaJOUZRGoatcB8oxm
QnaR1g//U1yixzc4fmxAolKMdtcMfMoij5vJc0NgXZNk3VRT0WATJ79GdZbhuUMNQiGIwTXaUVYq
y+GRIgP3KHtnF+3Sblt2/0tF6irrs2lXVn+mN5ZjIKiEoUkWJswhUdpi4bHd8z9dikmaB9ARnmGl
4HbswvMKs6x/Lxt15D6vjyVanRw8CQRo3w6dKPDQBvjd2ok0Ces5oYIuTw8ygUvDPM0RALqt1fuh
eYSpNsjjSAcIeni4gQPd3kZfgSQFP5tXA7CjW5OqfE9D+cspGSgShIaUbs/XpIshpXxc8O2xlUls
4db1MbTnMX5soHd6LA9mPBAk0qxbfMyqmSpN5GhP1QyvSnMCVmq+2gsZLJOMXjcQ7RzcNSTLA9cf
Uyws8KpzJrQRcSEFpNntHIEwBKK6kNyjoQKo2K0AjbiwqtTDxKz19B0BwlqkWzggwEnQ/q+p2KlK
F9ec9F1x51f3AIc7/aCSbXzcolmulXgMYeU2gOe7FEfF5fjMW46XqHrx7Dy6XA8Y6hB/ha7ksZ5M
GMeAoAhmAvPw6OSPtylKrQ6o56sKXQIWlMw3kxZR5UczP3N8p78JbSjOgfqARP7p5ycmvF5soxMt
o5bXL38hAhUl600j86CsrRLkj32313q9Rs3fTS+YURGiATjMH9pQoPGbC9QrovG8shIk+9kO1RTO
IAOF3uI7UK49OZ9ODc7zzXNC1/9ozIwFCRPdxtVNAhoCbuRJwKKG51qY69yMwXoe7fLeVsoNZRz7
OMMKUEapVqFFKd9nqcH/HVHbfSzKk5lUFW5tuCaHEKQ6NqZFKyXCZZlyWL6gnULbXCJsjuh76ago
4YWwhYhgdSn4R/P8BOhpjNF7wRdHwznNvWD5xuME/NmmN8lJ95oIAvmrohnJR+UIFZ+ZnYx/I4wz
JLQQBBujrxo5dYf7HAwiVEY8lNzrZVUPuw8Ssxj6iCaknNZmpiYYxybAg+nuBrWW3mOqVz0EpqCw
/MOyWYNZPCnPaitccVvS0BKEtf916WHcPkF8+1Uqly8j3L67F8v6V8+LbTzaeVvahystOyDRH/nI
EdMmr2qQpmc1ILs9hN9j4uaEObLErxc+NtrhajrC5ojQe0x2NB1kBEULYQeJiJT41XCB5pdTe7iF
Ly8l+EkNpbWbJWLu7FtdLIep/PQihH5jQt/eQ9Sm+18DT14Bi3ui3fPSLvcm+Io19WhvdL7l7oAD
EetOTg2AlTCdrA38vnEgGms0/5lh6il7Uyf44WBKa2w5Qn79Iw9htY5ufKav6zibKMI6pLmQgGWr
HkX76TdkNtqnzWvJwTO4LiV0uobreLvR4gb6IhnYtm/IsCui3pnOoTczZrqA1EXem5lvA1y0BnLQ
KHW8t0VC3TxH7w6Yh4lRaTWmMtGtTR0NzFH0MZsOKL3my0FGgIcCmmPz2++Xp11ye0zJz0iNuhDj
Yn4j9+pSVfj4Qfcl+/+nAEFd81gZHL1EfT91RYycyhD6qdjzuxOBj3umRf0L2B7dF48JljtvivSB
df8FpjF9jG8VFx+C2E3rwXajwCYMBWlbjDvwPcOaNHDMXy5ebxVYBiU015VMXLBUGCMGSPMRRA0j
Nef9N6oy83ZWfYoXkBXzI1MgtVbAx4jwPQGs39TND1NL5JjDrv8CElg6IPdWdSEt+ilD2AEdGVcc
Z5MXcpUQ6xTEBUUoRCaT4vEpSSJy8mo55zp+lQ5XTYR0zErXgzGx3oh7jvg5tTGViRVuIzLi0Oe1
kXrg9BT3pRJw0IiC01vrJJgVJySZ/ObO5ceif+UHCxHdJPuva6yhmm2weKOdq6CEC14wbHPic9c5
Y5IvJxfUmKj5Sdbm8AC6DyQrvFwLCXqmAox56kVkFE69dfBfew3HvBLijZ5TvGZ7CM8p9WP5lfm6
7oQmhIAJvZOxx8mLVmDK2SP8xqJ2+48el0U5ExepxNB8o29spZuFgARvLxzDHS79aXsG/neRaLcj
X/j9dUomkF0TwL+oT7k/K1v/oVHA1FQaNQCJTInYmPZfOv3MFA2U2M9DwQZWNn5WzoQTOVdyTJ/V
f6Rd81HCphwS11Nqqun4IGw6zXzdOd5qQJzPPZgaY2m3OhPb1duP8vFNUog0HQtOwcweUyMszQYF
4bVk0VX5oi571Jl6eelTbNOTJ9CnI3D7wI65Wi5pBAKNk43wOe4aLDgyXHjTJcpQKQ39hrWQ01eS
/kjbnacUIFe0wNUWdW1VmMB4yp9Ub+2hMQgo/sKjzCLMkNm9B23y4kUT3ze/C1BxYB0IE+A2BXIl
E7BWC37kd0ojYLTQQhRxDY/nxXUx3z+usP1JRKLlYXQm4YZ4OY6oFbTp7wBu7Saa/Hb1djqwSRK9
HwPtvYhuQx47CfHTrwuVVERzOu1zAET3B9LVTZpL1yjnj2UrXV/X3k+xbazjVAnBZWW7ihIh88fS
LGyNhv9ZXfedyQH31SKwATc/dEBrHjMA23XrCh6GILctRlgihRQbNPuuFbVHsC2u2EZwaEsqS+ex
zJyEVdJR+sANAGDKxX6BLfP0B8ysIfohTPu1GBT7ZOVb9sk2fqy4LcDPAJNkLZs/hGnUVQwbEzl0
JHfBcbZM8mFw5wbMLIXNFtrdlel/BgvxOScTLGonYcIckXmb+tBe1X0vda4TLYpvHjicAXrMMyyb
WSHGYd1+YDClUAUtiM87Q2tm0axQ9pSHX2XlhwY/PX0lavd6Mz1WPzHgHZBlB/OwEL6hjhyDqaJE
nJO3/QHbq8kgjRWmeuvGMJZ4Ekb5mBhHJrQcKuptrBsW0h0ORIeAxyYABZ+/Ugx68hxsHFLTs8JD
It7C2UiuLWI8yI9ufdphDGL6ot9tyf/56iXWJfpbw174Djjicnma5AHwGa+dB1CbmK4OripipsET
Yrciw+7J8yXw7+RPigTKE35I6GuyTeLalfP/hcRv2scFzsAASmTxUZW+cbWSSGePuHbYVq7YesuJ
Y60GYfw6uBKK0H9Fv8TGbyENpgR99BihD2PP/bh91rb5KoAIAaFICnU3kZBJ5CsnErJsbXggjQS8
iiVeUkqCfkwGIksEzZlnsSLpb2HUD/EIQ5+UUAeJ3gpOcsWSNuBlpY3+P6ThlmkBYPE+hJzwmLYD
9luHJaQVXWEMvUrY0YZfbp007G562+wibUzjm0m6C5Drnge73zI2Ux5WzsBH4VSE5Bh6qhM8BQ9s
DqrN7ql2PDqPYMfI98Id+nQbgT7Tf43F8XqMZM2OUWfZo7MB1z1RhgRVeAoWpWES9Qd2/0VXnwAf
+66r6xXCviqpO/3o2GrW0jpdwLuwKKCDlj0y27vBUPMowTaQASHsU9lLzSbJo8rdbq3+YhWgtjMr
TDQfNugC1E/5AZ5N8uyWSzwLw7HwNnhvpxYFG3jaMqdNs1c6QnARzELgLNmIQtXQmRuRQRL+Vsd6
upG2WCw1if3MQFvWdKKtCqIWQhKGOb754TQ2h2BMFDiIbpotoiPvSd3EmlR00MPXpxSoB4QRhm+D
fAun7E8KrsFKSJL3YOX1pwQSnaoU0f2dws1GFxGgUBz0b5XoH8SMVIEHecfPrzLMohhF4sYzBtbl
+BUOZriYgoCr+LL1OtS1IqiQ7WdxDFsnHbCZ1ZKPWWWZRKyIqPMOnvqCNrlLuXLcHUyl/ejkCQ9M
kFeHXOdGfDSVwK9wZTDi8RGna4WIJ7pKkHxTgNBYbDpxVXoj5snYRr4Ry5K25xKLOGCVN/bQkmzM
h2o05ljeVktGC5N8FKO0OL2REYa56V1ZBJIGsjXC0U/J85EjvXfD7kEpyXO3lUICx4KhF+bPBLqB
1NR3pOF34acUK/z5P2LDSbNfaGh1KHGcRz8u537Ebw/eI3N8xwuY//4aw6x0FhjK+4DDYx5galiX
Bb9QV2JL7oRJWjeI9TSOgg6MnlnqlaL2YMFDnGBVaOu0Ppn3HwFY/QcCStZepTpBlv7G5vhj9tN6
M6Rx+ttJjS06ImmrvF2NOkAzN5vCOjaxXVh/QrPZkzk3ef+F01uJLhWqGbixuojPwIvhEJgIBvFa
eheH/AHhUpl/5P+p3QtiDUof/DZDsrOfa2VTagR/hytmHudD9GjyKYtArq3J4OnxGxCaqu1cO03j
EAiSNLpyoNSBx69ZKkJDB/TK6uw0bZWUIvfGWFixF1X+rqb5D+IYmPBHXBhAsdqwpmYb/2GtDn9w
PF9I0KSuy1969cN02emGvX+ZjA9XLiG7A2+5sPoYiWgDeDUQPH/1f01jVHAVNr9PCgwwNkIWaXAs
mgK7hXjeD0nBcmI+EzwBsMZUd/V+p8oXAvTOHue4u0ilsL+Uun+gq936xQFJO5BPlwZp713sNIys
739K3uzuL4dTNB0Eh5KDeXvhKMpid6Snp9CKUR0pkaQbr8Rf3pRTLmoA0ML+O+QAiliq9fgF9+4B
AO/QgIUP3WVCe4BSVfBmdSpc1JMvWpvU+eXOqWq04VWOIZh8qvclX1eZU/0Porjj+KNBNjbuL1Ot
5/2M+RPOfIF5uXblKfqnNgI8UeQm5hJ4iL4TqF0gC/9Rv/vvPfvt3d5vIJtZtAY7AAccbfHvoco7
DJWsSK6nEUOmJ3nRb2SCWfay9aFJOsW52CELNF3jU3UbGj2Ur57Ydo2d/wMjnjFOXL5jAqwMDMrj
aFSXkh1zqGxBcBnQm+lUWLKQ4Ln/LchLtcgLpDmIUOWtPWUYD2Cvp9CDGms0Erc4/QOof1SOCGUD
ZkHiHXcu4g4FpfHxO9OnujIO6C66ydMTzPTv/9bzbOiOgcA/KpkHLqh7qzCE2Xjn4K0PD2SDXTjE
5DovlKRtE9kBG1RMOgzUHmJNM0CzGfUJ5ndxfQc8g5eRVa9W4RZmRFpb5Sn40MSyqgWQzxKxO6jf
1/dYZ63XPvNmv7GEW7j29IjlPq8EOe5kwT0OA4hpMjUD160BrUY6ogX2O7DkbJsZaA7waRja+jwz
fkR9IwRkbxiBbqb6FfisIIqZOyRjQQ2vW5WpppRSb/CpLXbKR0MOyZPcfukllNjdDUQkFI7IwfXT
GbNCHLZkf2yZyFdfqVPWF0zLU3Vz7RNYBAsGE6bRxQf5QLPIY1InCcWFLIbBK7L70+dHS3Er4m6+
InAPN9fMLKRQ8F4wm6k4EYtoKAO+C6LALVparlvAEL6edQTMI50CjQkUs0oExQehAMTqNCtSnZ7b
NCLaHVPo0UimQbenFrnmiWndYYikYBeMQCaG8LPiad/b2L4+iorA1syZ0YpMjNLBYw835xo334Bq
xRhG96m26xubZtJByVSELXRPUXcRxSGoO7mqfqVFtXNq2u19RSE8Bgj/GlmSU1mqp0f9FrvIOUub
F6Hu9y/quYuhsboPUTL83AnYxnxVCSCGiCsCeRg4bsI/vZJuwYfvyAzWezQCGbeO2hXSZFlV1SId
UIwt1u5ZGvScfLjWKd6Tx0BTfmVtWzm2MhjTJc9XMXmJJssVI0g3fpZkhSt8FJWNmC5XlA0ZrJ7T
SGqdb7eiSO/CNcKUJ6kjrQPxuLE/SP7OPQu2os9cpHnEqg7/XLDgOFONByyLaxmhwYOc8J9BX4Xg
Esg9cyLyLf/UwjjGTsAr1oaCltdR3avtgXRWUc4hfJaeVyBWL4f3EU3z/HevF5X6SCH4bHpkOnMa
VFbPia/+oECAmplfp2k2dH1Tv6tf0QkHZqJHsVCOouUwtsLWNtZDWoYDvKBXmTjuiz3dENh3VgDf
NTgAkF+Kmk+2D89ja2+Tut2JwEi+UqtdUJkRZTbRv2CBmhO9LJjL/XrzlpiH09Wb6XDSn5NnxYDO
fFrtxBV7kLzVCL6xh5YJlL5gGkwI9lco2Q9N8Nd1IdmfPcj4awp4JCVNCd5gedUWhgK5Mk4TFZ8/
4kSb5I9im5ugCVV5IVlBvzAOvf4ilmqBLBmq4yrL1S9F9EKZQXgOpi1RUAjkkTyzXugAsQjm2DpE
33f71Lvdj1WLcUWkS2+OOYhGv4PR8Q2ncno1kuVU70TJZUcDHlatHIn77dczAJkunjp8POBtxKYT
kqBMEZZuTkluTQuonUh2CUVixk3vLivVI4VKtNWW78ha+N2XvRDo3njuyPQ0CvC8sim1djutc3qB
2CHFahAziGFEv998fdKdxdpsKxgBvhc2iiIb51Mb6qpQCVWvnOyLTpv9gK4N/3Qqo6aagTmdKAgk
ryAmTxftZCVwVUhJVX5tTQIduHHpVutz0O09cyn2idc36yGUw8m4sHkUiYL5q7BSs3VVjt6a1m4A
M2Wu6NhwhSXo8ooaZ5PUJo+aXveJpoYS5c9731FkyBr2R4QJ49vvYm/FWv8Vd6Be8bXZDaTI3acI
tEStC3W6jJ6e/ynxqulsb663gP9uivlFRR6jY/0Lfzfurut1wmRlTMqtyUK+1mRD+8kI3tvZKQqY
famea3UBWVQ34cjpsxy0XUG1e5M3yKT8gYBopgU+h4k7QhQ70bI/HLz8B+5NoBZv2aOxeSrb+7nc
Xs+SJJtLzJTqE6JIAvqgJ9G8D40G09nE3QghSu4xyOfed5K76ykQQqSc3Lxbj2THOVj7g2LBVswW
PiDyHKlUJgfkIo0ARb+/C33YKaPL5f+XYJ9UR23VoptF1xfL/NKlCOD6LCl0XlBKpxQZPx5HcgcK
FpLqVY9h6uQyWK3OZV3GHE6/mW2jjh4WVXusIWzrZs6QGUXbflyoSaHlgOVsU7NQaTZ3jdqSAT6I
Cu3C2SFnnusJCvKroh5eovb253glLYlhk/uneBD5s76BowGorI2n2nux3ouNUY41EWH5nhUNJjoS
1sxbzYb7uoACFjcZBvrfDdRemcIDIolXzu9r2ptKPKUGs7sfr4fmBxU4srAmLjLg1Fb9OmXnBxMQ
2vq30EW07xSVVoB661bhwCBKvJ6FT/GKYUv8wb3q3Vdf+iBRkIuMjblmuQKJlyS6DYsyb3Df0TR0
EAd4LeKNeMMAl6TFdxBv85WcacegkQujITklWPJwX2/7/2V33qE7dEHIGc5TO52P0+SyG563MGgl
wXpEHO/2zJqxIqJb6pS2whabWrDUwjQbfNYUJM2eKhoaMh+0T7J/DSOVF+GCmUeSFZbbwFpEcH4j
M4FTiqBrzTkbhH8KZ5SZ4gAHkPsHJp5DcbwNWUdkGNnKY7R2y5RZ1XGs/9do44UVO8ezf4WXKwYf
TMsnh/ZDf4GxFrvGRGgQp0pURIwOx3mHYvqCHH0nMr9m3uvBvaU7ProbWsadpIo2HGV+sxHufVk8
J16kN9hyv9ITddP86jeWP2UkaH6YQ7/wG0WsjGBr/A3+kGI7G4IfQ2RAiPu2lh6d23sIngj+4HXV
z/cXBkUM3tHd6dsoG1Rs8d+Arzsn/Y7lLE3nS96xVBbvdGwV/LFsMacBWbII8D9+CXeEuY4wbs11
8r8wGIEl4gsiaY0i0CTtxEgCbaU1fWIoxMNWiDoPWcAxvEYdSBmR1BJYQB12eNQfsxtPKCqK5X4C
2zWyhc65gbISNfrhDH7M3yX21ve1SgNsQzDjrFL7SooxJr3MB2heDB6Dx7A+mJ5p15DgnAEe+J6a
f8imSOYvNiX85Y3YoIGRM81ygbKbi4AlXAdAYzzF28YKm4hS1UwumxnjIK+pH1ekibZYR1HaqbBc
oC5t4lIbiXCFZZ9p3EgG107ZdTjzzWsP6hPgWL9O3y16wdAhl6+6n9SSNoLZYhJv75usdoX3FosM
AA3WtRY0AMxZvFX+YUNXsKzwf+Df0upzev4kxliMGERLSd+kvxJzwwYHOW53mym/4f0duAvP4uh3
YmeFR1mv0C3J4SdTFEbV8K2eawYZHR1QACI/eHoAbdPOltGPJpbKNjPZxEEdlrrfjnxjLppBU1VB
XqJf1DdDDM38hbtph/cUTMi2Cdd2tNVb6+ExdBBzyDfSkO4LeSk2dFDeJ55hp/nHDPFQPYdTwcE/
iupOs0SuzAf6siyOkeIRttlP6yugg+fBBapBiJhRfs7KT4fccBZwtmhCDMzbhjIOYfo79mtjY6EP
0qKl+oE6h2dEUoSxYHLa3bVS4DvAVvFOGlwveXosoau92LVG7S/xTK1TK42uqWmEyG4e2DMgAQDA
l6AMUnIfyLgsPmtG/Rd9MFDA16H1IxdpEpbq1ULxE8iCcOXh/KjQaMz8AOIj8BNqwaLUtuu0iTwP
Q0JQxhvpyYaVjz8ocOhQmcU443DW9wu58XfYW0XkmsgwFNlVZJyQf5R2LC8LFtCtDwb0f0mXfyvR
e18HV7P38mLCKXKbBE00AOJuKS8Diqh7DDVSXSf84Cy+yc5z9mYg8Mh7Puk7iqzBSlz6SNJySZre
+jU3u0J2qVgBo8j0pPliWHtvqMAsAAeKIp/FCP2KJoYp0+h7fqtOv4RtT/hoEO8vHR3rgsUNesWT
pfz1TdmszenJulfL2igd+grbwlfUXclN7ney78DL4hLKyxM3d+lJ0VKTGghQHem6vxHGffEne+hB
TJgmxrtBSgZEWqVEMlGrfQfFumllBZziZ6WmaKnRVggY7NRyZjyGG1jcBq7DJoVyXDW5M+Nn9mN5
fHG9YpHFomWOYLZQ0u4TIH9e4KCjyl2hNerznPvhnVdiSrZZZVwFQpu8cdYr5R0kKoXWkJG9M0Y7
hac+pQ7d3GfylAnzphA3Eyt3GvMRqoakQ/3amIWbm3Jd/dOsbpK4keXkIYLz2/epPcm8otM9I+9/
O2PhjbONhlxnydKUcG+L4vFDYE4yQ69HBzG4fGK36bNKUAJDsqZdFwvIDi1e6uEJjtjuhbmoc+L/
pHMjMBM/VMB5QwE6Bubu2iCOYyXFRD/QAPmp/6Y3mVdfCgF7gQEhRfcUGvhjH/mvaTV31570QzGz
8GixLqqbp/5ihIcyd1qF7WG8cGuZipApSHi1Q8G9lwU01U5L4vernywgnpNf1Gvff8HTxOIXRA4u
v6AR4O6Afgdkj56a9/x3y9LLT8VR5m+/w0+EROVvG04RYXNV8Ot0QyoYNLdya+jS4ylMEesQbPYc
36/noWioOUUKEjx7LvXR4oPSlH8TAUDW4GGWHMrp6Q8an0exkY7fkrLOtrfBelebxbpYe3V1odKf
6cQZARcOPhJGbCoj9sTqH6pcZb030NUka63grXiYtpiCXdnDz3DiMYejnp3GTVEoed+DbTejGo3a
qwB/chBfHl8v0ooP726VHOVfLfLyn2t1ES2bukiHN3M7v/Jly9GhrObPIJEMy2uinPbb309kXNVl
+AA/anAPumcNFSgw9Ts3wS5PQLbD5DEuXstTR9yNSRrBvClaEvkJD6ZyjRt/PmkWVTPeYbg2zOwK
peukZ4F3J3gqIQ3SMo6JTbA6fr0kXOv7eTcGRCdTVbHA9RBYEyBDj0II1VvE9aUzrORQZxz7cYD9
bAN4Wc1oiVNECVKIqeHh9lkEvqsEKVL46RbHJJatLChEtCbpy6tD/mrcvFQ//N3ls4YEiib9KZqW
qItKD/S/F34Laj48aSTe3NT1+C9sywXU34R6QEzp1OcdNFEw/9Qbyxq+UVIvPANOuNhn287Ugw60
WOCZdTwoO+ceACdHb0k1dJIedGZ417Gppbtv9Vmkwr+yITicKDMnPzviws4c1gURu0j66nWTnLjO
HWlVj0dpC79Dh+2InBkbTc0SU0fjDKznbtOOsaubJcvmEIxaTKI4E4JEv2P1OclW6yKTYHkPV3Ok
YMCceWtbQUU8Ese9HlHh1ZaJcqaXwVCPst9SZXfS44fc9VFwiva7roLDHseY+P04ABkL+V28MluI
9WeVFeje2VMEaTVA6ULjMv8/8zD/+4txdmVQ7+YsLz6AllIwTUe/BImE4LoefFWtU6l/38oXfIgF
BlwSWumZCNR930wwpbedmRNUbXV5lcYsgW7BcB9J48DiMvJBB5cULEXqMWB1FflW4ps7D3ZOgZay
2WMDodDNqEjNSBFahTJ9vKYZDY1FrPHmLgRgPL1IozLCCFdEC+IS3mqERS1GbAYJ9+2Op0E2pzKe
C45ldOWVJ0ZeNq5IXeapweAwAL5mYcRz6A26fg6XI0Rmrre1ZdQn1CUvJ0junyFU7GbxFhhWcPAt
nyZ+Pv6DIEFkwvRE/PNm1dYY772Fxha7RkLCIzT281T3KV4/qhbOxcoqeZz1Cm6GJaMvo+Hqv7Js
az+pKwS7tbMkwOZzNhWVrNcQykDgowAVR4fExQKPsyR5vCmVUOgtIUSBc8yZdT+/VeW6ra5MWdu7
kWXrU2yGpr8kBBZtp92dc9A+jZkoYCRTuqThLYD98Jb4AI2Z+BqFpAIdnMmK8VSQ8u8u/fIP5wTp
0CseJ+dRjZ4k1wPrfPxBznexpizd+Wl54zIClAgBHZMiA1EadyecXAhkUZkbAiuY3/13WYv6kRkK
MLRo36Q3tMq3wcaGP67j7OuRaTIzJBDIcgotkGLJ7ORF/gagBklI5x77uvwfdEon+ULoakK7m2KQ
7Y7LwMVmM1cm1nkzY0ZA2AbrjrF8eAWefW/RmtIukUqDkuo6ul0PRvPGhxk23m6mRl3cIs8H9qNc
2bGCYTsiDENGUEJsa6Tc9BEIyoS8u2uIM04j4FuXIuCGr6IWJZJURDqf/R/pvab6vmvohHhd9Ce7
XgRc0yoOJn2KdlSoRHvHh52C3W9HBkFd/HvxlHyDy7+glULOmHWIjW25j/nPB91z3wwNZBtx93AZ
ns6zQ6sv6mpNjLrbkyAS2bZJHSXIdzom/kxrBDgZrx79ts6OCD+BjOPLcGd5lIbH9kQwKHTrMvM3
M7HVBaCNEyxDcnk7yyGhxqogFT6Sll5UdgFWDqmVCD7rna9wYmsTtk4QPQZwiVx+6IprK7CrxZFA
fMqUgV/vrp30p1Ga8wSYHR07gUay+iQf7yXHGXJKcpyjcKzw0Q1Di9z4wvdiEQTmzfYF3pRmLfb9
/EX5rSDuqg48745f8EywuM9xpxiebexqPFIUNaP1MDeB4JMAYsvnhT+EAyZKvnoEANXqRMu2j6OG
9b9IE+zROn/lN5UE3ASMmd+U/5ILqYN2ic1dJ9rpznVh5yNTzBrjEIxh2F9wxxd0Tbn+VG8mWj+E
qoL0CDBRgk4cpH7b+0xf3+/nqtZ/mYx77FcrIbKZs1dhYaVCKPicfp6p2AhSgiOPbjT5V3Xdccd+
92JrzkqJCL7ehvHkFeIeZVcw4kYim8um+H7ViLzY0uGC9Ga0MAS2+7Fv9lzx0mDbnKIl5xRSxWDP
g7envGHnOXLD06iJ0bdBe6JdusEVLQTKc0dkEH69aoHDFtQ8sJ0tHH4lqTvLUglpkonEkpmaTn+q
vgz8siAc+rEe5JS6qsZDERN2rXq4eyF9bveF0EO61MpNeNt72Y/zYNnEnn8xIo9Z6ctS0Y718FAf
kVqEgIzrh3XuA5xr+8ERacNSjZcBoDkvM1Z4bG7ZoxdUtMxMCLk/qEki0LbW7VZV7tLvXWszNmO1
9oQpZCegDdMCrdcgmWwGFUv74znMqtZQnumKOGqQkR2oJfRHkARlKvLgppslPBvCAvBtsfD7cqNS
cPRPssMilV/ON5cJemy+/bcVNOSEvi2G8SL8TnPJAhDEUE+6B3BwdQJLHZQfYBFmOJMhnVKtvXi/
F/bpwgdu4e5gSY0YxScyJX3kRcm9+siemEXw7+OS+R8zmBwl1YxEO+QyqSg0guIen+j7AQVz5UtD
Y/358hNo2cIEFEB0D1vTK2kDpaZWI3kVgRDASCU43ZE9+E28VMPh0sdSXskrYklzwsQ1Cg6mLDz7
DaWuSIC0jG7m0adJWvGiJ9bIv772L4FFXDWqU+8yf04H/t8UclSHYlecdW71t1n8BGhIjQL8jryD
fx9VEdoMH9sFWvhEIDk0CC8Gtv81MW694BiOsQKe5bCobkfK+J6FTzDZufngerUwOuYvChROg/d4
zjBpokIlFqu9BrPQbnRlCJK1Ti4fKOVkVljYC4xxX71Kbl+PWSD3zkWGRGYW3EamHD8oi00/MTZX
fA3nxEspuFGIdc3ZNK+oEROhZYZmPGOjPg3wThpLFezi3epU6cRiON3UdpUMB18LIJNEwi7yqTTB
J6ZkOKi2ljLLHsI8bVsR/M2kMKR70reZjSzT7k9moX7Ic7lX5teJQ+A0uDP0glFp+RkLRc81BhZj
yV1ts4lCTGS0zpAok3kuN+lAjPiyBC3KL6r704v/drqCcmEQgzOvhPPPKJM+J3Fi40sgCc10yk5D
+Vxig2js8dIhI6lfi+qxdk6c9FDCQdv+MWeB/YmBEx+SeojU1s18dRriGlTEIFZtFTwb1veDWzGr
YQxbiOl6F3JGu1w2w00/5DkesVtFANNMbpEHictJvSCiX+UvosPGcd6CA5FUgYwzr/orc7QANmcH
mFWlKKLFEUVxg2PlIcdA5Lzeu3P/S68t1KT0J93FEm3pkVkhifwMLSuIE1OxP0AYAzsoozffzrxV
0pWhKs/QFLj+hyIE3ayOYkJaSJ13jdbznd51GlFg8/mBysl/GnbWcpiRee8NNS5Ay8edQ5sgG2i3
NHPEUDL/ouXTk+7cEEf264C1j/pxFF6iS3TNBde6tjnvoU1sS6zRaUD/uoMkf3MyFNmzbpdH2zGT
8Q5sB0n4ViG17M1cu44yMzdbKVdP6QooyKwBiLxIMRir1HF2n9fVbJJXcRFWHOvNfC4xy99bIqYe
sIKV03VhQDl/rtnzJxn2ChGixvwgaHmc/GUOL5tYmbZbP9/3M18HpbLzxkBvkJ6+Joai2UsLl8WP
BgHKCDwnQ5stLsf9XnV8vAQR+UiIHaEdcc3c9a/zcqFzRkz+XinUSq2vCmBFKe8c6pdMETye8xRr
4jvAVsT9NwEuvRAu3OzeoN9YxXgxXC+HmQoNNM+8xu2HbtyNBs7/AEjGM7Zb9A0o/8mrk1VlAtTN
P4Mii3KcTvlqTTMyS7UjXodnW++H7o6BHv/N0rpK00gfAc+Qy5SIYiZxyHZ9UBt2fY7gEiudF0Pq
rRvYXSlmcQOPiDbosKon91XLyhs5jKs6T/q0ncywSRPHhYJPpJ2zNb20rfBPuAb+6gw8FN/SHQcV
sNwkAjDgdCv6pAy8gQFPQGwVzb4IXGHH47rAl60LZgIcgHoykXYWXfHrzAgNge9n5lMNzx2Rz10q
rmF00a87zBwENzB49fj2gtLDiNq5AC4ntMxgID70nITnv2JxvmSXPUTbWotG3Ln3A1kmkCy3Wzg/
KIYHDmCerrFnJAc30thyYyEZf0F5BGf+50Rw1QVukgh7xoO9dIak22R5kerkE3tRCdtxGlXVkl04
MlnwHbqk8pCf2K2M4DM1JrWDIYAjuttpGVY3r4d2dk0fJLGutCJT6k3Wt7o/EAvnmuPnvAfwMWtt
RJd0Dhzcj+IZt94bejQi8Xpl0qwnNU+JrOxjGdQf97l2kIAiiIHhVcrkDoj2zGBCz7kvU2uYPSxT
XNXD/OCd8g/9OGSnUtpcMBLxkVt18Z1iBthFcqi3Dvqh1feGUe4SqeK2EzQaVNY8p0C72y0VL9+8
EorN5d59qPsbbzsOHlGlOsutNpW7ZOe6vfdGNQazbJ77GicCx1MsM6snUpzLd/u+YODEX8J6xul9
dz/HtaPyFXt+haSn8Jp039VC2kHfVQGck7nWe7Z7Mo04uzyDwXWiEM3Qf1ze353oo+QPSCXWuseN
JLLz2GO5LHdpjv65qsb/fBLoh3dl0bo+qGslV+k6FGSFyTkXINGMNe3jS4rrmfbl6+Etkzv5XY42
kLFHCoKl/134xfcE9jr5bC18agBzBdcbKw5LFTccYOxpAckk/aBdaUL7usqJH0zpTne4H6ds6vwU
bgg5BUmmnmYTS8lWL5piQCKNVggCA08obefMSXi0YV+wmvH0E5lGqneaAhSGwiq+9cI10JaFOxhF
d8M8qvT5kCWUNkKqvEKcPBqkZ3VlbulHJapGR8RRAel0FPupVTyL1EE7RL+tFkG8E4Ua5QR8tKzf
tSrK9ezfzik9CMhv20vLPtvdd1D1LCj6xLI7OT6FlnyzYJv+PfRLZwY8XEN0R7KRsmi/YsDlSJJ0
Jrvng8UreKWF07YkiJNhzpJJPzNi9T+2nTPC6ps14F51yTxC79CaU80XNo5ZQJjfemN9eogf2rA/
gAxXtuUeaBKFgQaYA7nFqVHGRjpyz5F1I8RC3I6OpMWTIiq/vfku939KaVCAqQfhZsYDk0SMTVwk
5SpqrCMPKB35z3OYi1d+w4N++UzhAkxwlpf5UuGLXlOPHw9ybWZLu316s5c1BegoEu8jcufOvE5z
xHAdT6HBmC46w3DIGbAEy7mHgaMQSbo+4sJwJ6gmSYr1Y4vv2UTIZZaWIDhiL/xCPeVv0KpPAtxB
Jw8CPxcwV6Th9W/7b3DjnHxwgHv7Tu62af6m9fYAPF+8So5UUJo1Vv9/wsK3Iz4JxBTM0IkD7k+6
ILYa4O+Ym8PVWOpDRzDe7k2U4fwYxUZ+689KnKEPN7K12S0Pit8NA+1vY5HpQlpzWzz4j8Yh4C0C
tieB++As8IvJfn09hEBNW4RsRFQmX1KeFO7nJSLCaYTt56X0fzqs2b58K6WwoSmkFd/HhHVQFjtT
bJG2qyevFrFUmOZQCPRBwYEtvLfBvIg6JrgOxdArnavH1fvYCXcb1gbGCwbYFeT7zVIUjXG3xfXt
j5pmmst4Px/VSqIajPw7thedQR6p9mkpplGGe6E8eVcUCWPvj3oo0VMYTMl/C8//cDjUdLe1bDtp
7bKkhf3kWcH/W4QUsXYPCAer7f/O5vMl7wxpIGj/PmChOLV2Ztz/tfO3aik2Y+vPDK+BFVW48WK5
xhz5WiV+GOneochEgPxqJna04B3qjz6Nvg9cSBFUemxEbsR6vvkui8RHhiY85mHttSvxy0gpfMlV
I0sAORZJVumjt+wWdZaDlBd7EW2u/S/64ORSXkkETwsohHWn6BHF+3VLecIozXtdNxUxwfUwKdvR
wIdU6Y62JxjRjDRJrF724bmfFsbsTdLIrsbjnox55U7T8AgMsZNrcMzLBxouZG3yconieelJ5xRg
Jvthxh9ejXpmxu63s1KDRvqPUcq+Af01gNlNK6mHU8beljskJr0hyFcVeJ+uzsFKoLEhBq+SBSt5
p2kwL8INVdeDmWT74lF1xQIWvchJzrRiMzMpHqDgfDo4SNPjTOQjwXvgVRoVofKsH2yrc/KpK0FN
3i/1ExvRfnXib+PX60vHzNLkfJuE/eNoDnekLZwjyrTFhkGSu/StvIwVl5Q4FKCRvp0HFv9wJwl2
KjNuywBd7cf1G3y9ckpVJw4EE03138NceiRpoFk9AQZd7FzEuKpaPhPXztKUJvYuAuMgiOd64zdU
CT0BGp34wWZrlLBja5kViVUl/YsIKmNSqijEJPc3wUF8YvOeOLNerJ7kcyvMEtr0r9JM4M9sT9Nd
O5gQKy637dbT5KzHjm1awdGppchpGKeOf+Jl1r4vyhwaDgqOz3yJjJxqRO/wJ/aervbeixVqbVfm
/DhZCNPhJa3D0C90XBFxN0lt3m55y6mc27uW/y/WVEufCD0Cqfsx5epL08lGjCm6o586+jo+wLhF
WWIkrsBRG9ngOmavei/scsCgJQE6l0T7dZHXxUf5RfIq/usmpjwIZDaClVLddPP58xTvJnU/m96z
GqwpyDvw/FhpjLHLF/W7zDuaBgfwUgF68Yeoq9Pu7wqqtiJ1ZZVXmfgeeBWluFgOe/Yc1Q84WI1w
nmEnvCLXvh1j8yPwLDAH0ryhslyrC1F0asJbKSLeuhKzOIe3JwfbqIA+DKUaSiSlAJI3cY+aGIBM
rLx4X0siBEV1qJ0GFQnOVQYN360IKKvdWZnW0T6EtU1a2G7jB1Sa4Ll/8sWcVSrpTR9j7VqT5+yh
479LYzQNK7uzc+RvGQ2xF73I3nMOPkPOE+8/WgHHxIyE6ONIXwYNT5QCmn0go4leGqNxrmVkSehz
/ZAOqrIoN4BjKugJ/Qolnmuox63QhsJMOT+qinxLctyi9tdcfB6po7xOueXuftE4I5+YwJffacV6
EQApvUenJEYCOISKFyc012Rf8rq2eYNno4Z2fI2daBCe26i4R0mRj7lYvoKM6tiCbx7ub9pD0w9A
QHjuSfQBQhA+VndOKZS5OknwGezu4sZpnXVe6gewDUvewDtNUFOk7/okS+3aJ/iPtIYtRed8rdlu
JVHM7HO/N+VUgPmiUNtxw2XDL2Qxv+VUrvCCxNXAadsv/x7r0Z4ywrEAABQkO71XQqLxpvh82r5k
CkUVAcd0JOxFTHA4RSRnb2SkQ45FsSC2EDLro3kemsoBEKp8qzWbWtkjnaOjxIbIc5IMQVt0N2JY
JvFIWjCOC2hZrrChOILYtibE+wcnoXgfhcFH0v4h3/VSeEBHldIg9u0Utwm6zNAkdQ1ok8bdi8eh
9Ys4dvgJGjq/r2c2Kp++CENwAH2+G7M9By78RvfRcMubIurc1VOiR2qeYzWg+wRQNHLrwGPbCEFY
47iT5MHb64JN07Zea/J3hFlPGNHzHge2FfoVSxyEX2yskOcPChet9LQgQxQggdabmfdnoxC4sHB0
9M7OxlRWyUEmLtbCUBATGBa/P4paVpb8BsDFmv1+wJSEuIrvR1Y9pZR7GNi1ergkLRdgXa0VieEm
bK/Ek5qpP3KjowIin/VL2Fxyv7f+8HUv0G7cPV6hR8OmOX75llogi4Ic51HbZ4+Zw/voKutJCj2+
j7x6GJFD8z2CUJxoyvCmTLx688K3+D+F/Fh9I+oWq2/HwGjlY1s+xBXFKfVGjYvZcpTlUkvKPG0W
JB/LOnOAEfEYwWcyYhjmg/fF72iPinxNUTMXD3cbBReDALTrJp2RoCTGSHLzIbhFeEnmDQ3RaAwN
O5hNVJ/l7Yf/ebjyvNXVWHuwDpRCRHDvHHsDopGW+yLsMdBEx650pwxU7VyS3QsG+7PIAmto4Xel
qCKcHrxZ0lSBeKagK5W61MrufKPf5UD7rwWt3jU6Pce5MWldLIhCD3NILxxkuMTF/kDrK73KeOg+
Evmr5cBVDd+k6TnLDG8BCC/dLtryZBVGLrFi2AD6UAhG9qacRW+hVoDHTMZDk3Vf6uQ5FLeq4aMQ
NsNkOGzLely6aJOM4RKdJHEDzV7VYinsoULKVT5JbFsJj0/+JtabYKvBl5chSqrXz9nczW05jtXC
LxF3in+l52zRcGdgm0wwA5UxPRLoIDyCw8eAepay2wk/l+TkZNVnZzwS8jSsmtbi6oyKJU2ZuSXP
Bxf1Mvs1MdB6iYELoGYNdVQmSZvnoNBp7Xe3/ZpicHmALL3PZI2EyQ5VT/i87pMdW5qJbufEMvpN
2f9oU0HRIydQWBgvVdbUan1B8M37sp1NmyaNEDAX2+jDziLkJE0TZ0vQvucX1KU8/oOVuf8feZmF
ZsSFqTIKi3bU3rOXSJdY9YiKbYQW0wdrABYbK5fqDUDs8Ok/1cYN7Kck1zR42+au4ycSK/ekToY4
M/1xa+rTIGG/m4S3vmGtGj3zK0zt7PsUZS0gnfdXcaEfh9aLZvcx/r2ebrA+Rp81itX7dmK4Y/cw
2accadieC0QA1OBodFwyo4envhfMq4t7s3RqVmn0QNr3dJWnayY0deoaR9MisPZnaRiW9AVabIIE
0scnFcBFkyXAOKlpijk8ysa1SOaGBxdx8JCcERCix0WYyeVpkbUA38ola/bJRJE1zryETjZlQd0B
Pp5//tcb0e1l5CjOIdjndP1FyQsRJUp6T94qK7igh4AjXF3yM1s78qCxhlymxJNeJOsLKbQhiLwO
svOPhE0LKworuWLcBZpzT7xEYSmIIg55qkFz5YZfdz46KJazNVWKPjoYXPQqSSYZq0nL5kxxsSlF
DOeJlsRNH1TKqOWBSeHXDc91X0LRoz9MttQeoOYYlVfg9vSRzYbzH5NqKNuTIPKAZSJ9cEcdeb72
YIQPYaaKPWuF7oN/l64yocijTfSDRliXusN0b+LnIxm0hfkq6Jjpm38gj3IabScyMkwwRAvLYFwj
tRuGB7wB7jkoBGD/tIsfc6zuNqnttZk9C8WYfWh3E0tUJeWB+xVp5rNVGx7cgqZDMS7kG6U/I5b7
KF2J2T7W2xNZeVFtNU0j67873nTw2ZsETakPR4XXa2xRMf6G684IIEGNdcrse2aspnEe7wnR7iWz
XBJhZfHTsUwvhH10D2r/sDeCZJNWrlUgbEFvDUMdVKWxYBrkCtQQRLxr69LgKkD3xALkT2/xTbVQ
llFi5q7zm+1K+UccL5hvGBONlDIdIVFix72vA5dVTraXxKrmIhNj+3WA4MzFPOHP+oXZwBKzzv8w
KyJg7lx/2/UvP9YrSpHdFLPgoNZDSUmrM8g82TW7wrXKl9FGu/nq8jjK3KbVYNlttKsoiynbDZE2
r1ftfWAuIqVH59u0lyx7UDI9/XeZ+lIZ29DIHqzV8mP0csxj5H4poFo5GFOL0CeTKwu4eRm9ue41
7VhAjBmL8YL1vuLs+DTlG2eUc6OHbDGbJlqeoj6eB74F/lo8AE9OB0ZiSJ0zqka01QSW3NpfSSof
aJf8HKVFrSnJBWlnV3ESOu+UDCoWzKK8Xtf/7dmSnplnlsmMB0JMv4im10cHlgsWY4SNeG+qIrXe
KZRZjuJuaoXRAzX69A8g7qkOnbSEItIiWqfnqdu0uH/JyF7FLMEX8MoHFVwECnjLtkoYZ6vVFQKs
He9SGTyz2q31zSrx4VRipFALhpFmG0NifRjPxRTFshvtuLkRCpB1Nq6WtS+V0w61Mt6gygshVzvu
RQy8Tr48qCroB+1sp3TzxPgF2Bur19AjJU2VMnNhZ9q212KxpbTMHEc3AHJnB9WHS5wK+bTH0luY
vj++UBM0ebtrPiR34UMJoDcq1ICqi3nSB/Aj5UQqbz1n1xGfMinfBbYW8skbWCw3DuphY+uS1gt/
DhRratFKLW2yKgOs3LAQES46lDBaUIVXHgfafhJIIMGTFB7/6gMZ5s26DDsW8x/uxnmUHFEoDOjw
t/oyd7zfl6a8LVX+sag4QXH6CgaPEUHWfNwy2LKpigSmUgOSjdLgOuBsl33tCzOBj0HhyuwGsjdb
TAcI4TX7u+rXZzgMgxzAgQvQfw29B1N/+3SKc3OW/YoC7y1XV2qLVtODzMyb8rzDy8VUlcRHQHDZ
P39BS4Failkv07LFFvgKzOw1kjm9Ff1/jzIks1cMFsWfRCqQXRqi15MZ6ws8YiBLn6Cs/pBhc+kz
itTW7T06iJsG9vmwAaCjEvjjwm3aIzMXUDMScyNRWtCQnhNV2zlh8x80T2CWxCNRETbQNRPWvjB7
caIoueOswaZZlSj/yqzJpk8+gWph1phb6WhHFZNfq3TvSFzI452M6mcIG6U6qe6xR3jL1NhNSn4p
b0SEpa4UjnsPtszepUBkX1CePhHc0eRzkj7xS/hmCVAcFAPiOYngNDz0hrIMXfRAUzQkCmso6c+o
uW9mrWypBiOwyCQ2NSdAfGV6iDHYmML7ukHdbAuKa1PSeVYkZ7biGHXj9Z2dPXHFAFfy6L9Jqm2z
zkJLdwaeGUvFc1Pxb8CHuQp3YoKTLRWWYeGqMFVziDLmmSb0bXX7TtvAO958RCD/MIh7PsuPRjbW
nYLRj0ZGnfINKNpFFVFzDu27Exygwd2zIM+0fC7xB1TKA4Y/bBfJKrcj89jCoXnmBa6aMjwOqEE7
xO7o3rNtCu2vZaQ6dCXkCmsL5B9xPlVpovQs0RBjwrWzKgL99rHU21V85tFAUhwT2JGQrwauxdgQ
o/ukk4+HByoNahm13cYamw5jgFpfXcbNVnoyZmKDxxXSTF+7Kbmj5S8n8FCExuZRQ4/EWIUtJduh
AKA81mf0CDbQPz/YnD1IihyW0xL9gPh/2traCXrD1+bL8eFElZY2UP8LHeUeC0FYDO6dZLY7Zpu9
GWw4SVTX1otWdziyTf1FY50BrAGaH8mP9+fzguqF7PCUMduRGnS5h02W4KP+QQ1xRjx3J1vF56aK
8uO1XsGJvCNXL/R+/kSptWPF10LpAQDi+x4/r7JAy1719PZjw1j79CbDqZ9GkTw4HQMw2ZOgxOvK
+E469JNuH2RyNL64Q47tqQ3wWDKy/9EbuaSCl22sIQC7kdx99YhvB0IWbtegDuXnsh+RKSMF6rQD
42CG6iORHQOkhaxtFcz53a89Ftzk5+Yn2NZ+w68riGXMJ7GKa8ny2MRtT1wYUEyRCjwyFTUb82Sp
O+IS+FP37sR5VKTSDPM8tFGo2ro/+s6uz2+Pm3CGcQpjCV15RBLE4VI2wpfGUCdDBvmTC/g70U83
aqns+ADABYA2joWHas6ri6wOeTFSRQWecsReQPqo9aeqw60xFlJp2BXZ4ePU1aX0bwnWwhHxWnO/
5Iav99G1qBROpoupZdTV+4sXuneZxTOrvNdXcomx0tLM5FA1+UmYjNPdZY6mUxopqYBDeQBlS5eA
cw8AUuxtwXuSyMrgBpl6MMaaP5VQUgCmYllAnEI2SWmQfp0wFrVp5IZYu4oDNZ+pyxIeMRdndGGf
1IICqppl/xV47UgVqzlSIqRJCWQh0qUKA7OvzlPDOz5s62jyHFIolU7OppO9zcb9U4jorteYV7sr
uWMidFzlegkimy1xKmTXZiPU69bE9XumOxLzOcNppQeE0+5uEWwhG6yPXnkekWgcNk3HSw2JQbFx
jl8JAw78vqjSy/2uAVD2FdI88+pGBaeXk2vN/IqRDmFP+RiJN5Si1ggNujvsu6irXioLQPKUPzhK
Pqo2/TAC06wnpXjvclGQH2S654U4jjdByQdDzf46yhQFwiHXlyq8pvOi9iq6SkUUCBwTuBfEdMUy
VCS90ftk9f0T3SP33pgaQ8A/PRGgSLPX+N4JNO4k7wCUyb37AYAlfda4RVghCUrESsyY0Jk1WLio
etdYFQxIwSzUAHNLSHdA0+iGxUlj5F2Q5r0wZMlAmtmpY0d8fF501gUD7Rwv+s3dEE44ydO2T5q9
wva983+whpF2t8z9mr43Dq+oL6QW2Rz6Yqxaysxv7Aba0Wn3S5UYJyzwe2TEctooeKrt1TZL+xcT
fujXpAXHfJ1+cQHXPub1EiUU3DNmm+bXO0BSRM1P6F9/Lg5dZdLrd0ot2Qz7rTRgMQivmzHm/krV
AtnMJDJRCYImVYQwQW8NrXKB+DyJ+CoulkQPWF4LncgFng9FH04FiytxPUKYEv926MDEScg3FJUz
snW9LPVUNhi1vmbTTOu2H2jCUM2xI1uWj0pRmyeUbnBW05eMGIiyeqqyMOpXVhTt9TmrD/MZvcEr
etOvgcnTV8DQLAHdL5sEAvXY87jeXj4jrYawnLnrKsnN3vT+MF3ungYOcohqlfEWv6JM08kvv0T7
j/0MtMxsHnS4XmyOtef9Gzf00TwPbkVFkatXGUPIdDGuCl4KY/REEUAN0Jj9yQhoX4lITJ5cm+jX
f3RhFodAQ9Poh8TqJNA9FumO9u4EYOd4LxKDrHUJqIKZg2VjK8a4Kmnok9lQ3Ozotach4XEfFE2K
UJ77AwQ/SAQbgzSe3TOZs1fKsLUGWGOPi5jzkcxvsWTbmUI1VA70afwFkGJVphTNK4egCgVRieI/
KW0iUdrDG94KSmu8A63Cn6rQo6ymMAZKokqp4g/jQb/VXZ7+vHfc2LvXiovhdLlbF4ZtFjKqzCey
T/ds7w6guHx0PDyf9Tj0sW/ibtQQzlzyt8EJNusToE6SC5xs76TLePwUStT55ER7gwE6dz7el8xw
/17bIos1AiYrFiI2aZaowdNArHxNxYPs0R1g3LV/OjExMFIjx4x8ke7a6CPnGX2od5LN5Ic3JNv0
pmcseqt5N2S6mxHuNsuQhfaysmgYpRCN1XR4z3Pt9ZLef/NMhZ+aqX/Y5rTmkoNh5uXYbO/g6/Hz
dD60D+u5nRhHBA1LmU9dqXurGGxqMozMdxR7/Z4Zi9PyxnYN7SFeM6A7U0Pzy4cJy99xnEZgPpwI
fQh9nbDmxauYcjZCYyzqnTkpTplE0e+xqlmuzjoo2WbTpS69U0A4kCnxH02PSiTc3q3ehB9IdY1C
JEbeb02ZQu45YxYxNC0ovAeE/2bMDSV1z76b7Pub9d8tLwCATMIU77xHaP6o3M7ZsTIcBYZ9+XIZ
NE7hC3tNfurFv7FK2Eve6zJ9nw90RBmu7kcaxKgP6kOS5ArrzLkJnihwqMb+dTXfxdVufJZvRU0U
oAqMicqh+KJa9ivvAhmlulcobAXTJJHifhfxGQDmlLecDfxcPciYqrrNLu8LkwUq7NbMwTUpw4VY
s/cJmr9m4k44Zw2czF4w89rizOrt/BS97N6wth+sRtIAfupK8B68nxuFMBaZZnHWSZqU7TkR6hZg
tKW0fjcfepKU7yM6k0+gOGPt6P3PJIcpbqZoNYlxDBnsBk2GayM00fphaAX8Rirpq5iiZpaEW4Al
a75VhncUk3Y+nam6UffY8/jNcMthoHqbkP4PbkOu6M1FctQRu7J98O1cSBXvq0/hz/rLZAub/2y3
dIiuav+oyTOiyuT1sECgdwXdpdYXy3TfC21xQud9BQXb4zDXPagcsL8kNHuz855i9dC2u/cH6O5T
fT17aMNenvbi8TpC3ZPeuVwHDXdOvIX9aRUrryszD6Yi55M/rkOjdZql9tL4XRAytQcNzeqlnJfe
7wuUGTbo7c9WxGu0XJJlmVQdSRHyFLs5g6IYTv0engsSfuGod9Y7PrCz20T62Dd25ZWcPXQXQH6+
rL6dom0xZdfRrR0rw/HNyupFLb5hAEqyKT8QAq1iHM6PYwUTea1IfzRf6/9tz3qte5o2SL0DhIT6
9MlUEw0Pbv5R3iHACfDZwVSilFAa1cmbIEJSp9cw/VJBh1A4FaN6Xmpijv9jkb2PI0StvhiQ5V0k
caPzdrciZ1RT4nmVtLiWAh+C0ZzjBorWpOhiPCz9DUhL4TBk+sQZ4gIGBMsWYmqnKmgIm4wKbCbK
6rpbPnJAf+CctkaYCgD+erdE7gkAI/UkfE6XXKKasyen0+seetNXzjsSl5XPJqHtbeIMA8gGwazV
tfeUio2Rw5DifIxLZVw7xakcUuTwE9WxNv+6LxsVPhNAzx1ePaCfu/Ez1QDNkz2+TuA55wQthby7
RNOBUKK2ywtLMO1SC+NDt38gqTBU5UY5fO3MnwuUgN4JSXAdWAc2FsFkjJ9iJn9h+mC0fQxhhHCb
ii3oHIbS46mLBMqfMSXbrfo3Oq3+RyCXAbY4J0oF5cyTgHakqavrQYuU5wNTMvjPVvIxUwYvKQz7
ozHlQAW5Jr0r0AgYxE3wTHIbsFFbrSi1eE5JQYDL0KUIXLeZJ7M6K9Z/y6/ROCP5IZH71HLO8/bn
+mZVwjJRE8I7xVIJ5jCvTfxj1guODI6yn28K1J9OY6PalLnTmC6Y5eFwvrjRlh+mycICL9k4zZjy
AkeuilHSd11BqeTLKUghFXhtLhMUW1zfuvK8l7PYrjcvfMkTt7u75sHgl09Im1MUVvWrHH/Wmi07
lMQxRbchP35wRIxA44wZwrV5OvSzN1Q801BCora7z+tSyIc8SiXFZ1revAVxk0ZhokT4l/HLzBMM
VKlg4lVAwaid5cSBums46wjOlz6Bw2FuojkL+8epCgcv813fGpAg+yFTHmiIB4R/dfm7VLZrrnhO
S7JdyznkdYnbIAF4BMJqPi5y7FcXqo4TVJaZEySrxYW2vxNviVH2cvqHmS/X/2jrES5/VnP2FnZV
0sdaTsdm344VVeCNJXfJlSIsDo4yluxSdO+ch/F+Zn8A4RWMlISzyKv11TfBjn2EoHN3tdcQEtE+
2Eb89CMe8m1M7Ms26XnwqlRS1evU/GrfhpPjmCh2W0w0DTu/PPHW4nh+4xXP+Yiv5q4/CD3f8wqy
RxblltQ0qA9wGBRIDYY+evoYh43dU77k6B7mj+iTNj2AACO/KcOxc/Q9CcANhVXiIcvvyvdSGB7F
1kGoO5LUVbr8NJevqev+RP9YLEa1+pVJCLXD9qlfscA4fp7cDXh+fqJgiTCXJBzEvLcsYQI4vq6h
i0N18CobM9nfoTj8jfsS/BvtOS7Gz9Kic9VdigHSexJ2t6RzcVptMxpUc4ZpVTIwNjRXHfPN6LJx
EZW56yrnSsyxQGVHmCSvp3ThER14swpAz3hxIB1tdAquEaIrYT4nxA5pYRWpqVANcFajMpOrf2nT
lyGJePkb8qjBJh+9Sq9g5+8gikdJItSDDxhwbD9dIBCjCWn4GKzUg48iLdRuKhMlLxP/f747uBIc
ipHayRn4ji4gBrmhQ8pUqM+yv7Hqv9iJjssrImlfeED1pdHpzgmkvhVYoqruah86zdBcUzCTa0k8
ShIbZocliy8chSCjbpfxBMYXoboUqDtm/lJw4pG9Y7/8HdGr+V4RP6fS+vF6PJFHVZU9joE2QQVB
6gVAToGdkXPf/ybGbBkb7V5Y0+5y5kwFkmP0gSrXpgz0Rh59KGD/oqLNs/kxdz05wvWokNz4UI3/
pmkiO7bCsbGoWpKW9tv8DobMENkvS3Y6Y8VXSxd3r0dtvcdo+7vHqPR7gNoKdp51XiQuRARlr1YO
E+jGIyfrJcURldUp5TyLXiVWFo3mHzCuuWeRQasESB75TWIL1L33OhilFh/6XoNlkaS7t2HYoglt
lrJVGFW2+VsaYEv0+Uxg37uy/X7GPNTEf8SAMPTpP3+/GXgcwWSoYRsMqwvOLRj8MUU7PXRBOTH/
WWwywcjoEKeQQyqvXOiadbkalkqfQS6LnxBazg14OmluLMzr1xn1FjXvXhdU4Pw5/FrwQXOux8IK
04B6smNncot6kruyhrWSyf3eiNcI+6N2pWwOMqoLwUiswMIb2y5E6QBC+BnT7eNpwpOr4KtAMaKD
LUDTPZk64aQuANJmv5tSQ2LnF6gn+WIwu4R0MbO0L6TrWfqrnNyLoDuQuDFRRCLstnFtFomXv/8S
zqAZfOKrVJD9pKbCoXm10eoG6rjfxjLz5+TZZl4jk103t4FCdQ6zH5cW69PciEcpPjEQHvdu9Vqk
QBExAfL2czT9LdFnROQuOX+vKUf3WCPSMXBIHFQZ3swTY7FdJmZwJGI7l9fGhtW6RGCMIu2gF85y
1Jbz1gMGWAXOFPPM6tgElgt4CRXA0sDZlJhqoWs6CT3mIs3YS6B5cODnus9idwqxWPy4VfZ6ArPC
+tY+h9puMIpGAiMlRlTDdYkyQmF+4a3wKaNRNenLWllj/0CgrM1r4f3pZWtdS+YYA4T0Kr6Wv7WI
Vg9K94EkopHJTVnr6Zt1cjeNo3iTpw2uJ7OBvD50fNsbaE5RKZO5NN4YKWDLCr1IkWjwrdysuWw8
9YGabQIwY1QfDs2dRtmFLz9FLW43eJos7LLynXaXJfjcGkdovvJWc5Q+CALkTYjANWHAPVXHWLae
Ou2wjTEXDxvP/ohBgsWeDwov1sAEHh+Bck2E5r0Uc4O52oSLVNNR7ggx3g6EIAN0tkFp1WVSSRQa
yrR4i9dfdZgG7deq0VXKLSm2SZzRcfOrPOvT9OdtPFv8m1e4sXqwxAIVIXO8vaCZ8izKaFV7hUwE
C1qP1NCw/bwTgr/0mUOJcKog6vOysVSUTycA5YiNPzaWcZLypPht9CEOmh7z7V+fmopdQG1HvY8p
GT9NXw5eB/yspirkRKJnSLSe5cLcsjaje4YJzxNf3xlzrh66zT3SGuKpUNT1oCTw/XIVwvMXKO6f
LP06bto2C4zfclTRumgYREZoOV2d273Kf+2SjeZwTwrdf5a0Uol0h2zR0G1rQlsyygxlfxe4MxHe
e0JJaL6hYrJ+hXa0hCYZDqMr2AX6FG8p7GxvNWvRny+D/cLHeUvdXVSzF5s7KDYakbpbfyb57AHI
dKbP26gqhc/r36x/+cYILB5YXskvfPpx5xVrjYXCRQKzgYCAl7nIIcIbc1qt8aVnSQqMlwUSYV53
msmgbLbdBRIf2ld9WapMBwCl36WmcQo+WGmDth5bb0rv5mUj19rhomH3wukIBHYG9LYTXP2zjWaz
yCcc3MLmemzbSts+SuSvsbPnq6kfnNo9FyrGCLth9aGZGhuR6sw6Nn+oTQs4zEl7oklgRdHpoU+3
AIgS6aWBnEeY/FCWWTnv9y2A0ObLj0iPxjKxIweU0z3Co8qg04UIh0BqhLuXmHQyhnGYAyBg9jUe
rkNRDcigQ2YXAVygIyfWBOEpNoz3mmOQHBB4psHa4/6l4RjiVIlGn9oquY5mNTpDu4qVbs2ErSXq
0k4P1k69CFINgVGPDj4ewHSkipeD5hNIVfDnALlLF/cpDp2oT3Nht01VURy4LfcDgNQpumSD9unM
0e47+OoqDNuG6/md/LsbJLkFPKHIBu5OJ2UuGQQRIi6fvitu+V8frKmYLuGRuGo93bx1Pkv319BJ
KJwXrWb4rVcIgI6c8USm3qZo9W4WDkFZ62KcXdi/jNMdZUtWwWSWR1+tYfJx2WLmb+ueLHVYyERU
8nnQZ79x690BoeSk5m+j6nUGNfzcR3p/WG6cCadv3h9A+bbjt8zPvgjMWbOkj7mo5czWzhBziHbF
RAkavD5juHwALsAoxksJZZoDhKlKfQmY9xK8CpoQvyQIqwWcQbRRc7WZsIM+cR+/CKhmDE43rpSy
dsD6pG9uT/afwYJEadqqqaaUyECtiFGDgDsTK7DRJLoznflQbUWkKhnH5bAD2LmJn73hOOoXhQqi
NLwqCeAJPtEcPJx1CQHsSkhFTqUANyJuGOB8zMeS7sIKOvHfRVtuokS4P3x4VUTgaJHq4vwS6+Ue
JjIrGG0u02zmTdlWIZCkQQB+iHn96U79EiaTpykxbQ2Q+QztLwU/gnJDADHTf3+wGTylSEqa9P9t
YTap+oE6vahKtefZopMOAdqNFQpjmsd/5/vf96kf+yBKgIM9aB9pdLAxvGQRtQK3BJ+DU0PLG/aI
xiffuJuaH4JEatNSpsWeylWAHQ6gf4jn6XENho8o3oJAu8+KX3pqAB3uLRUWfZnF9tZznLXQgmm5
dwSmCncyFVDSFekm8F8DDlevAa3jDZVoC0FIwQzsWkLbS1OylQwDG/qwQpk0xfQYQpSAEQVaLEpi
Ip63RHRlHdihJxCf7/Y7DMOyTEg7xMDRO7iAl91yU6jvyCvVZTmNNHXc38SWJY3vtgLZyQXINO8W
pbr0kg/N+jPHLweaOmpcRmtnW+cgZWjhlF522Ejn3edEDWNpJ4ukjodR3rn381zgw3JzJd5h7kWx
LfRjw6jln/Vtm4rG50DKwDDgbS9F9nZDP/Pf10niOBfWFtEubfhEBLJ0T3N71a6/IcnsRFeD1XAU
j0mkQDqYr3Jvn8D0apOeCP1Wip/Y48dfy8Fosap8g4eAZi6WCafEr+lUyuTpU88UCCk/AR3tBqkV
pTcqDcKpRa3SbiraV7osNHUNXNZde1OzQaRGtiWq85MAfUEOb+qeF1aDAx7q6XLemz9GC1SIMZzE
ewzqh6V7rto+feDCazuo4LEBG9XCocu4qSFWqBAGKNurgUwlUgaBoVmA0PqkI9JN8rfiQU0mNnJL
/83thAjcfEB7PAoT7LdmgMUokbKQZk7qWBD0roFgPoI24g6rK1uaqL8//4n3Tub8IND3ZT9HsfEo
gWk3ODoXb7TGW4zJfEFZ7MGBLPr2wSOkvFk908o1zZnR8XlKG5gE1VadvoMui46ZauX1F4tIBngZ
j6WmfYvTO0WUIXHPt1iKaPIyGaJcL3srVcoBqhse4DZbV5LQVmykYoySwviyvJK+uR6+neTZQAN+
4Hcm4dRfNHt4lXXnV+S0t5pRuZw3qeHC0gqfEvpW+a8fk2u2wUujeIiiCfUgdSW5Bs6LBbSCLJko
W5q7Vc9s0WHN7j9ZFk4mGXjbVNWqEh1sHacW9FO2T3i0xgcB06LuLOHzSE0DZlKvGwx3gL8USjXK
pjvOp3K0Z0zWkbYgvcIvOeSjyT76n5SCAhyWHLQKWaGgHeQbEnAEN9W0WboZ6u7q9Re3wFjRX9Z6
UstbEF9rJLKZ8l9XzHu0Xb0eBVNI/3w27K/cqPdpxM7H6O7S2s7ykb4KBS8crzyyaW2U/ev3L4W3
iz+WLXKPAeFI23u+vRKSnzjfzjj7zbm4QGqqDL3mQb1HS2S+5KFlj/0H9OGEIbouPeGN2GxRCoCL
3xygLXNKgkhNSa5+ue2fhsPZfUkQlxJ5aDpmRNdqqvP0ejz+0TN9IY8goyAbfnPzdgR3T3LiEZZK
fwI5VWPih6ZxTCBRNLJ25T+JSvdfPXiy+oDE5DlAJxl9eaT+tGtxTQ4ilAdm4o8nFAPDbjuxCNxx
6v+Mj8rgVboi8VZJdVaaMSKZXNZxTj+vZWLgBKXU7vys2wDqSyS8U7xFq6y4Wdr97V4Twp55Ul/F
59fR9Iux3wehnvSNE/Ljhs0w7CdwSN6vskb/t6IreuZ2MADZVIWNC96nKby/1KySEtfQ8IjrUNOF
pUS5DnHNBWUs1FNYtctdnMLVNkEGxTQOobMFaewSzF3e8woBTGsLumpazw6eu/hLACwhpL2jm2Pc
NloIkhxITvfQn+9nAft0Y9IkWNbtTy+QinOpSxXk2+G3Ji0TT2KkC6OFM71rHNepSw1sQIsxcZlU
ll0FBKFzqomN2RhnyD+mg1+LGcptERP5M1s/9Oxy8ZEbzS1ABl1cEb82QLeVNwbOE6KjzUBZZFut
2CiKzQ6NB+ZPwBrlTqnzjZEvUCcA+wW85/RkSenfyY/2r+D+juk2944w2NysJnPMhk0wT84TNy1d
s9O3ZFxJYpACtpSle3dHwx0CnPbnoaYmXDlpEtGL+sgDjw8nWRHW/HIIb0ZKlI6SaRMjVBSB8M9G
IWB27Y0jI8ck70XjxfX0LnMhojg04O0ztYiAGdEmsLn7U0j4OK+Kj+YLwjkcJ+KYCEG/RrCyN2t8
wk+wAxbtSpbbjPojrQNoeoPRykRQnQnCBMxsKUZFDAFlT44hd9waFKg4Z5zUE+6H2U/kkc2fQZyu
Cm1fYhV+mxiPJEA7MFsItvCuPZtGM2l2Yd32Jvp0ArEsqvCfKQok2kbGD5dUVDYrje/+V4aPe/4b
1yPK/vFw+U4QsGipLZ/eSaqUJRMP5Y3MOldli0CnIsCsxuyhCshCrcx3+22hdDtbsjl5boxwW1E4
uvT7Yg/CNYZRIk2yIf+qD1PvRS1tqjBJdkiJtZeqtkCs9Nz/Fvw9ksLwaMOz+uSI1TnKOE3LxFWa
rEpqCtrGwvB2WljcsyKr8GsAv//UgW4/fA3DNcbxeQrI39cSquvj7nhvFp+59c4r7WZZpFSFCsDR
hx7GwN/ryUM7E8om36Hgnnxhz+zJGbQthVr4Yj1XahoXYFhRdnlky6F291jnSonrTF6DrT7rcd/R
lsFEY1ZZkep2LvnHxeHHGNA6ASrI6s9iRsyU8pRh1uzVdu0SkIDNdWWHlqLXX7wiz9eI3ryAQG/0
yKLzlu90wYn8C1wGxb1UjrwxpK4k1wPWF622v8hfhNyINU9UP+tKn6mPtgGoLmsnuuM1amdMcshq
lljk6EPmmobM3LGGiP4CnJ/qewZMVhO5OeXOJReVK5cGH5JQy+ZQ0sh8z9UnWdTASGEmaEwzx0GV
gZjQnUe0jJxynqeO5CD+3cgPHXKPNoar5gDiEQ4j20tYqox3HQm/c+RUqXQZ4lFEqRCZw5dmsCcu
1IicIRLMPyz6UMk4DgugZBNce7Yaxm5WD7R34lVNC9gapr5nAvsnVUWqy3LogTq6K4iv34zwmEmF
qVZHFWJWAf/PuKODSZ/nf8CWG2ICoLafZKz9KPZ40FPo3r9fXuI0Bsm0x75D627MqxOns+Yf/tYN
3Bvslx2kNTBkYOWJEdczCTcolk+KvfqpREiBxZS8D5l9m6MuCpEPfLpDMXl9GNlb663BcQuc+NNs
1XswOOi4S4TKYDLYhQJDN2EebJNHl5tSm34zKMR6f4/6AfUYaMJ5qae8KbKSEl51gKQ74FUswKT7
9KEmoZhUWbAzgjW9NfYUB48vHm1iPiU8D2LLxVrqMkiiCv14tdutlRQnAVy8Jtu6uBYAFKdM8mKQ
Y+yXq8oc053PrOyK9Fflg8Qd0znAlNOELy5s4hUfAkCVSeDKFMtS/LAUCHUwZvuCsnGvCOX5XOUQ
Z9jU/WhkUKU0U8XNBLschkp0Pc5KzrGRJYEhY7TA/imU301yGbbW2HU1ubqQvUWxAhwwRAU6aoD6
6BNLJ0dRH/04AXF8zPXm8j7tD9g2SDH8ZCgV/GfqllCLFcWuwgZtgQRbOfNLs7RIQXqIbEAPq5yJ
rbZ6E/TQn2OhzJcakNijHX2uM1nEurmCCS53p8+gNFjC/xsmSP0p1pi7Q136LdZNNhwThCCK/5D8
naCnKbFaVE19y1bD/Ftl8vR1BgtWJA1//4MbBZzLviMEYIioZw8RsDzvd7poa+XdqKJeh+0zYUk/
VAdDesL29uo+3IZ3EGE3WDT/+vpOGR3uBZIuVbgJWWVuwzoPL2alpbdH5QnbkCJM9VQa2t6/MhtM
ed62MlxwJ6KXDbiVSPQIXwaGy/ELVNuMuOCWUPxUkiDKMw5FQFv4TCbzkuyjpa8Ht26h4CdsaUhO
+0eI2hQdPAW1oYHnh6OIxxhyBPFpxVNf0kzNL5X0jUHlrVrmYb711yBOfJxezSH5GnlCYsTKWvkb
iDLbOLurYaZiLorMbAPn5N7P7qm2sfb448hgnbkHvTJc3Hxwi3GldcCUTuqE87aq00d2czTuxclz
EvahB8i1amBnqbAXpDfohKVdIhihIvpJ8Tt7dnc9FxuHMwcOJxnEXBy1jCUC1oMZ+yaBgxKV5Za8
nNScWrDZtW43Mkmy/zTXnjrVMaIfBT3wqF9tyepx9ksCpcGqeZmUR8NDgTRxY6qi6iLS8/UxWnZU
1R6iV8zz2jLAiifU70yNVHyOo5yQ25x8LaKGWE+Og4fXvsLqUFQA4cLm2d1yKEKfeD47OTI6a5Pn
Lmedc2XKqGKmDx7GIEbvnaHYO752q7olmbv3F75sYjBXpMpbaAsKIyECzN53p2SKUw74yjiBn0Pn
1w5uMCASXxAn+0YKXpTAXkYTk82Pl4Xi0VO9QBwc+c73DCq+pmH+WoWZZYsKQeqwIINlryGSW2Lp
4zIDNtURBS/hAR7z/sEgWLW3khbv0pMLA5dyke0Xi5TSUAR2MAcOa976z/AHnWJja5K5DQqbeHyz
8scUJT5gDSysuVG7696+EVT+k6Idsy9ZnsZ5lvmsDbIpumpbWfQU9OKwFWNeuJRz/QGqkWPDWJHl
jFK5qZqKHUP6bT9j5aA4Y1iIpauDRIU/b7WlKFzBQ2s8OU0yvHZsT02A5hg9PWLmZOxJx7M8RCWQ
AJV61vfirq8sxk6j2qaiMVWY9hGGJF+D/huX0h2LxaBQU7KNv4DA6td3bHkEC/rksmtY86hI9KBe
vnHqBIRyeP79tmbpBbX/tnDWmR78c8R9Gvvjl1mPaEzv9SSa/0ShzRFMofWHE7efHz9XQ2XBrnyG
ejbGeXct/0floovzVkrdyGf5X7ko+WbCjR8CL7exG8pppzjyAUIT4owUJ2dJTN7feYJk7Z9/wdKK
aRh773KT+dkx++/h7kHRZzNpGWuRy13fKTuRwaTbNdr2TSp2vFkuKkm1LsXsIUIfVOg1g+kYopGx
xheOoQMZ5dRqguzDJM0ce6OkdlzZeWKeMwDvc1GMuGvkazpDCW+OhbUQx7rpLjOkodE7iQLpjCOk
NUxhHQPxCpGcwEydOwF4kVuJXGnR33oeyhtJyu8byshmwbYpehiFoeb9INe4Gv8l0QGd20c4P3hU
j1WUogddryyeoI8kfPRF0PYG7rh8kObg47GCRwdHZN+sjl7p5G9xb9qDAulEPEdSl3OskLmqTMJn
9ya/CjFrPQKdaD5/8z4n8Rt1LQcnWoUNeLFVZOeeqKCyGFErylAzg1iBPcRQBQdqCu2D+NsB2zLe
872I3gRHCb8LFIpwqRsGUlBKMJm4IiMbL0E9KPvIxsS1YtW8mjJU5n/6UwHencgRuJVJS4BFijW7
Nh4ykuz/d4+6ZLdtW9N3hiC/EAnmsuQ1ezJdC6tjY9MW7J+OjANXwNExDr3iOEunx6AKRxauXO0a
m6N7pxOaNZI/+RMd4gcN/G1tfbPYff3LHZOi2RJJ1mfTk6T5fC56qJY/gclkO/Q+x6Tu4bGtSRIf
nFOFF6RIBBe/uNuvsyPPxT5y00dU5BsHbKdXFahqLgygg8qAYDjkXx5bx/Tyk4Q3YfJikpvuyq38
dCalTCRIIznMj2TDseBVv3hWv0Dpmnt0F6nBQScRNpX1kBzc9d7T9I5oV+UHrPdY6i0IlqWSto5W
H+FApx2XPjlvEUowXYiaoaeDnl7DmNWCp4guIDxTrrYOvn/Am6gnwc2qMU2HHbBYV108ds3Ad+lB
MHmQo3WLtmjVsoPi2+HOZmONYTObqOUYqiYqm472BTlTcaq+S3rIqrZKHMCTVlFyMc/IlM2YRXiN
rKDQvHymfXE2px4f20wbB1oUtM14TlB7ioIWg2ymaxkVX4/NWWiLoXiOfOkyzz9U4iYyply1sXf6
fbOjpc4ZchYKUohVlSy16jLbP7vS7f8SY6+3tH2f8fYNDN4q8ojVJw92pKtDKra3zLyfbfXBxQYT
Fc4wBVBEklvp7Dx/9N2B+xHGj4Gn2NkZGGjhvBnKQcvOdVDjkfREBr8HS6fXz4yuhb5q6lozM6xy
GMCT0+G3pm6O8ACezJT609zlC7Mjy15shCnxHxOMNcRZvIesC2gfeaziFT9hoNpyDt8ookczI9fg
aq7IeNksmBZy4vNFtKp4a15LvCI9dw97tD7eaeAnjFuRNJbYrhYxSphrJLceQlF990NaTYpodgqu
Jkrmi2XE1lFRQXk0ywVYQ2YY6vXNPpOQCfSEAojlEm+5NwBEd9ikE1brM3oiQdzG7eSe8kJqk8+i
CazGB0W8BfEZsCbsx4qvG9QzL/Al0511GrdaIj4J76PhMLddRyiJS2safsdjncltKI//LatDNbzZ
uKdhiyVJk5oDDpopz2ybSX/bcnMw21JVtf6EYwVw/YJiqARiEBpAnl3Hy3cIch8fsVxYI1ViWqss
VF0nbjTi8IICESmuK+abj/EjMMkn6EOLcCnLTmKiG5xNxOHAhqjgpLyZe94FetTNkFcEY7KlQblZ
+wgZqcw3tn760VknCugEPZOK6u1ekP0r5JPK0D+cwbWZqqwCTlVbQdXJv/+Zt+pFRixOa1bUlGMl
Tkexshu3Qgi4XCuM+ZEPmhIfi/0jnX25m8KysRdKNR6JDiXXJuWCSHnjnmOFcF4DdChAWYnM194o
yJF6YmkaZR5CMkuH2DraxaKfMuUBFMMcAhShpeyDq2Z5tfi9+SMax/zUrOMfjFzXdx4JJEa1kcqh
AoNf9MwbdBO0+ulJXcZOZOdLootUjR+c54A99KKehA9ORgSp4JvOcpHf7SHOke9Ha5buFIqYWHCb
M1Vei9aa/X+KEuuwv9x2+LGMGFZVWLBv7OUOcivRhUd0PYHtcY4AQTKrIcpmS6zF+OwBb92bEpg1
4TiAYPNTvlc2SbUiuohsNpHuxTabOxsO1tDhLsPPwBRd59KbEIY5Io3d4ZIjCniLsfMpmkk0IzyN
R466eMcHJR4YRWAbd92ZTCZ52cXRyqXmDt/LtsRIrZ9o83S0YDVZJ6cNar8DM7rqGBugO+HQ0QMu
gfkWOHXPKgKwYSYcUvUhVGDYVM3JW+iaI7Ia4t7xrjNee0l9Ik4Kf3+pEXd9UvF282Z38vVRURNt
55qJ2dL6aO8kxmRhjqMKr9qRtyRf6MNMPmFH3/C+Ow8vd3VL9cwg3RHRJRDGNALH44NX9XcD9eer
GkUJbm/P6vHehi88xJgx8nwBgb4l8wLlqyD0rxQaiUlUMT6Urx2fVntvZxATnfbEAo8p49XwFHXB
GhUDo3Hoa7awLhDn3XvftJjj1mc/zXGx/H1Kr58DHdvhv2aQE6bXY/B4JlLiVkpNsLJ3M+CtepiD
WSxGDuz6fVOUk5yBO/oNvPFj2K8K3VeYhbIZbBaHmTOFGjQTcwWPu17joOH3IAG5jOaLHHWCZqsF
3F+46TOp/wTJToRLAgGuiVYphkc5ghL2y+/zFSQ5svarj9lfc7Rv343jH1ufVlRQTnWcxQLBTumr
74uO4bd44XzFPQmSP9rZwBFfSIj55P6SE4Sa81zR1SYwLimztuF43C1vK3wP3RZDdzWv4x+/Xgqb
XAXMxv7VB9IehMNAztF5cZ9d67NfPq3hsN2gG+PWEtBStOOfUoOQFueN7+r4seWRpbWpT3E0iFoF
WsdIcKPcch9S5dYz0skRSDQ9+88PUMqGuKhwAaE7Ih8twlkF2SfE+DedmK1mocQ4RHe6rvOXOpGO
bkp8qPSMEky9Dqa3fljGtp0quE9iG/hCsZKMP/p4XNA1WaoTIjNU7D5GS8Ril3QqMr86Sglbv3ff
gVrlJzMjzsmvyaozl+n0Q8RA9+YMaVTFeKlqRDJ9CUSxLcato6B2U90a3RjrtFAcz8HDui0jeWu3
YZ3CDtrPVnKnenAud9OzRcOXRT142U86Ge9qqcHx8ac0eauXwJhA0lKtWgLDnDeZNvL6Kl3KSQRK
w2hEqZ5YuaUH0KmiYKYNT3ytV5Z17UsZ9DDBkRfvR8r9+Bp5Gcz97+SQz5XNjloE+uZpin5vFVWg
dIbmAlCdU/2dFK7BONbQuOSIWWcD8tHC+tesEXpVc+N8owsYn9Kh4iUEq7HghkvUxrXCSS37U6Y1
DMtooPQ6zDjPuMYsbEFLgJVzUGXie1SKE1SMLaLJociocxpfum2RgzQhmv7wT7l6GU4h8fs0CmUc
JBeLjoYkvftgfp4tjl/zZPxWEtZ7Es9hlOi7GLJZlVjC3xH3HdLfc2pVkpmpCrq2VUZXOOugLwuh
EWdliDy5uHtsP8s3CUixTYkvQxGyUzEGguoJYXZSrnz83SefwzMoNTfTp+7ZU7t49dYfDbGnlFPJ
BudsZVCAXPgKBMN6dlbei2Ed6mzrZwUllFnt1TTUlPRdV/VD/t+CeLV5shp8HH4wm0eqfgK4Tvei
H4mBd8S4kgi8OiCx0/djAuPJVnn7cSBCmgPl5pjwF2zD9EpzLzUGdzCNFq2Ph/AD0bomV2/JGr5L
17lU8rIByF8mak/G0hJEfnn5ksQYt+AIRdOraJqcIt32iNfwg2+xXgCt86KpuudQHQto8Hea3Fi5
OJChD8iP2NnaxUIQzh1fWaNwb+ocSbS8ceHCo06c/farBkFZLFZkYLrJqQm4j0qup8sXIHpq83Zy
4QPW0RSFtiS7KQw9P0UPuAlSr+nIxgrHJARZu3NQJaAwrbBCK3jYQZhsQFJf81dE3lTZwI3yIxLS
pZ0k77BjJOrRApMugJ00m8trYUyEOUeirEgOse0dB3pufohoyPFkpqsR3z7Qog876ktkINff/oqe
yQ1g9Z6xs9kZl2nVpEk5q47w4UYpb3tG1CrD5EVdljtO+mrSz2DyWhRzFTasd8mA3k7N1i6ZZ0ec
N7X19XbiyKvnU2eOt8mMUUC/40Ht8HfqwsGyObHrNtlVKMMHU8BuPw04vybHkTVn81BwnD8rDUEM
Vp1mkNX1QD2OJ2b+/rQb9VE+Hi74bmubLcXiNjdBLhODoA90thW5kgK1thxdGsaPGfU/OvJLJipC
jq65rbTRCMLJqFsNaL1qCJM/Nn6zD0iaiAZ44zGyEHHOtp2oodAdNY2WnMrKue3eehH0kKJvfTi2
6LLkBnQPW4aWbz7UJTOWSnX3jZBiBHNWXL3YimElrlohIwJGr7pDJVBOqHxFQrCodMvqWrbHXMM7
rQqjWwEq0MAL5QQqRcRqDSWFqknce1Yjjw1kCmtkERfGh3bBKYsdZ0vOSpYGYYezPD7NiZLWCEJe
dhDW8MDcHTtIY+4Jhr31ov5F/7z0rmlUKUQ6v6hLQevZoE1HfAtUInoHdQFBafrEUIiYZeVSy2DX
86yOVsoNoLsYTBok5G6FV/4flTPjPceTLO0TZTdUY2P8+dydnhitxmNIVGgbZI3+68KyLBZU/PgE
e5aDHz32XDsGOaAFg1GAmeJyVqi5lGBEBbef6/9AEgowfzQLSCFKHJpo/E/0qUiKc8o0WBCB+Di7
ZR73mBdReUQiV6QA7ZB4A2judgPJvnZYxLSNRTHEG+lpJwNOtIrImDLknptfuVMED1BHU9cJRled
e41kBFV2Tq5fUtsSElmE+N7K32xF+LO0hW7SZ849SwBWe0z/omDC7gncwdTUP0aVIlt5WSg592QZ
rE3nB3azAvMhoh8kEKBFdnPQ6f9Keem/Pr68Drk2qTcU0eN92X07j/0IllnpsU7EDcmzYGZsl7vx
s2X+AsaZISYjXxglJpHtN6ayRErLIxKj/N81tqGhFQ6HpWu768d2zAxIoB+ugd1c2MQretYRw56u
PvjNsAeCpxVX3yUnomo3BkbFQRCRn+EcvrNvnESCWo0cPCVKXixlc+5y+38KwB1wOqQQGSOhuz18
tsbGwasx9iVXGUZT6PQiXgwo3ZvLLj69ojdOi/QBWvrhc8nx3axZUjG6JA1+tI0YSUkVilIzYC9A
Yy8qatVjyKFQk3MDYDziHWRQX3mAo7z9UKDlmK0du8/p0ZUma5V9wYPHgQwatg2pBBSDDxVMTi57
Cj9HfWrgQWArKAB/xiw+6BCgHGRv/Ijdho3HUSDxJNr9Iig2jPufz+tQAULNSUhwjeJYgK/Gxwfi
s17zpqwRfGoe9aAizixOxk2Feaaau5xq4qA9dkm0gbhEF5O23wtWxgN2EVlrcOmKDgow4K0I3Vwe
jhheXAxhHN2kkqpTw/IQeD2HG2cEkDSNwnZJkfgyEmHlyoEkdIJVaFUAI8hr8tcdbNibqDCW2lgP
mF3UuaHDnBWvCAEVcnsRFm1JDkzJLjiauO1w27Q5CHT9nivWiePey6JE7WjFsk5z4yW+pQWMAwqJ
wpXmDFiGnTWxZgdPfbGIy6hs2jBbWomOYOmuZK42CJvyVcGdYFjjMXsSL9w98dpPUuomeuxnlZHw
J1iPauGPPBtIab5VrFO0X0vlhmXFctch/a08yqPj6nzs0c344YnPSag7FVhLN7etvSvWiUNct41b
7Km3sfz9PHgQyLhPx4QD69m5Rx+aVwG++R+xcdEJDgtLYxEoRP+bRmfXHrnAsZnhfBww8na0XhUt
vrNIHXB3q7MbrhnQ+KWUKjiwi8id6nEouAUISXhzFh+OlxfONNdIReWY4Ti4+o/fvbuKEz98pvfF
Z0iwomt5/CEdsDbZIwNgn1tyZ7uUmLsUeyZHijdbwDjGOzPIOT4nZ2r/2nSpXqMqP4IP3iJb+aZ8
E9QVRRu1L0rSe6I6estC7fbbDGbgEv6ByIiaLhnjk5mlBBSMra5hR8N/5ZFeJi9N9qVVEbE/d1kK
P34jHIDloUQhjDSafSrYAWqcNQfRbtqVSn24EBFM5fwwBJzAJLebyx26xTMkAk2830SE6HAXk90W
BuaFfXaqNX21QZnwEcb4Gfv02BEfoYfndLYRrOhXNxbnn8GxCNoNgtL/mHOSfAA8CKAOjfXkFV+N
Ao3j3TZs0lGlKxwW/NzPXqfsjL0gcxrYPTWE9AII1lbpTdXtecMWzvvfpSeg+d+g/TDo+6pqsMkF
SRbHRXqF6g9tqrh649ysfABJmjBDKcFdeoM6l+O9xFYWZrCvjMW5uE7hi5H0U2SzZmB2RClEYQLn
kxxw4iUgfHl6M5nQdMEvDLvotT57G5XLnNtI6LTVtRfjuj9mYlryHgP6R/W3emyLc/JmiKsRa97Q
f6drTFMZlqR1GRKZYYRyhEQgS7DU63Qny3BC9ghRSckD064Fq/Y7O+VE3OcOBhjpXqRWmY6irvaW
J0nj/vbx/u/PshtOsoItZ6CdKU6HyvjuJMistllw3Rplb4qP/166lmsY7YCxqYtqz/RtFnQzQkK3
RbdlZNiZSsKRm9ItGXJzVwnzPNr5e5M416ZYFQyEsmNgMmghJTNj1RkVQYUnAevpEn1z9W1c2m6f
mPUYr4tbEfbD+pRQ3Oo1OaTyhWMNnCBzFP4su/hHH4J9+TiJGisFaqYPMP/GtSujsuTX1Z2CoQqV
fJkJAZxzuY+okKoyMyg2yOVXlYfiSo9lzYCvJtveBtwqOQIhJcghqqb1isvXT8szWbXWZs8k8dSC
1hdVoBD3QpP8RHZA0dEZ2vKAVHAHdSRWseyhvjuXhy1O4Zme6c31HWiePB+05JwEh/Kve9VAt+vW
eZGgPgjvaQ6y0f2DzpJ2wEUL1bkFQvJkxx2vJPTUYaj5lqF7lS/dyvTGYj+XL7KROo6HNSq0i5n9
CFTDyTmQCuptKxCqgKF3zUG5LxZ4CS+uN4dOyUsJ8XusrLe89o7cJc8JC+xkI8/AI+Bl5cqeFHZB
knVZp0qHCCh1WMTN9Xv86cyjPJ6+ydp7xvkikTDqnz87sRzYVX3jeRMIJmQPDtjCZhMYhBVCMtoA
bOzhVnBCYlue/+PL6CcQ56rXILzBv+3TG4gf1TmBcedt7bvlhZVeUkvMQuUhaeKsGipLXdLHrVYa
Uo6icgO2gBwlJJv9s1Fzi+RpzwE1dsESt8ylx5thM3dcFPhV42OJUap8fcLQuGILglI01yQiWqDb
sUVAMY18XygVc9SXkdUE73ZIu4h9BO9CYMPFrQ8C+QhEK91gFE9lxB0ULuiL5o0f788mFbGL28Hq
Cs05Hhxel7L0lWhtRrY5+bkngLYuEuAL2EzsvT7YwS85TF/36tc0mXf3UZvwKm/h/btkIEn3kwpH
M7TcbQfGQJJN9pVXPkh/2yGsZ210gx7EZT3hBzmzpMkIG1QEOd0kPkE9t6Rpkyz2rDihslIlj91G
1nXnaDHYnz5f4jubp5eWCJrnFvGbLeMmPpynC4xzwYl1Nsz2+UkOdHxHJcyiJwcsUv6E1ObikBK5
Htwo0Nwmqvi/CZXCD0x0oi4/qsMVsrb/xdkEk8487k7weiaJbxqclKnB0Q8/tkJjwPPWyybswlaZ
W0XO+GLIYAVGzzhPsm5BhcAsrbybnX4rDiPtzrVhi83FzvuXq4a5pwXjXL8y6r4PxgtqAqq/R4fj
9avYdu0tOAmt3/rNj0FzV8wBHPYPxGRYilFLvx/Ujb5xt9n/Mnyv5Z0GxXcWmXvKP0T9Q38tGJYt
mDDwznMQZZEzjSGcLzqSGQvyo75lzM8tV4Y3YKMLo+kkgj6SIK3WJQChG0tdB7bBr9m3zgLa3e9Y
3oTt02MbAP8cVevgvmK+mej5SW2UO0DtxMKUqw8pUxc2I6df4Ubbm+++P9FflCnwlgYnvb1wPHIx
g+XQ1/YVht/gwdddi8XzHieYwy5aLq98Ernx6VWi0qlbxKwAto4BHE7WYCrCwrGc4NUkpB24jJag
mVtluqbZ3kRGuH57MiXtlSxmANPdGXH6cvdezF++HcQ6TbshOY/GODakO0dEahTx+Q7FzNSJEnYl
tSW9iFVHvHG5co2Ow7oGpMLDe/G+lJvj2GD6MVMh0QVcVdW42D4Y0jrkqm1MoMjanVo70+Fwoc/r
DL/R5rKCJmCXK6ZXvdvaeyAK8x6q9aBHWOZdlvshJhXecghGhB7twAKh8JYGcczIF08cX3P8AebS
y/x/v7XDvpy6O8icKvyQ9+wC3mcZxzKnI7AxvyvVtCqJPNxBjXzh9rKhobbBvipJiF9cpMnBP/OS
rv85B9idaVgpM5EWxmVq18t8oDUUSLUwKoDpPM0WLrX2o4z4+msgd1TRkBTCOFq3vmijfMkgxFic
EFUN/9TCWwqw6rq7fhKp22WNtJDe/WGLWPZK/BNLNg37hPkHy/a6i0t2/URRBZv2ZKKwgkCQzozL
6V6tAlEpkhssuV94bYD44Dw2hulABQVyGPLsh06DhM4WVk3FoS3M5yepSBPyKBqWVrHUeRSEq7yN
4mCmPfXibI/OpaO84a0p8sv7/aB4VrUjIcv8f8DlVyV/cmTtTgx9hqnZvtaGPzaF8MUwo7iUlLkt
TYWHYDCYbHoY2E8PRuZ483haKOGYX5KrOFB/6/lpxnBSgYccUl22cHjAd3JY6S3mxNleb7vcb0VQ
sBqUkBfgnD4pudyJ4TxGmiSwZ9P0ahB0RphW6XI+oB6sccXvf66636w8tXgctKQEtsN77CseBh06
UP8zdzmmGN0XSjr5Us5lKqBvdlCIrgdtFl2/9RlCA0+RngAUw++6PEhl/fmWy0Eevs4XC7z3ONJZ
e/Lfz408zn/oc9GijIL8AkNwatZoQ5YZzlgSiADfWTrE7vI4xCawRtd/2D/ZaQ41SCS09uiZCpC+
BXqX8v2ov4qHAWpvJEeLUa8TtIfbaLk59bOcSgaFWs9Q/CV4XOG5TWbz/tBjZxH2evrW2XlsKKEX
K0eReuiblM8zEuajObLqE+bBceMX9/nYYRUwEkuc+1DlN6NzhDmVZ8JDXbEjBMQ7ya8Faf7IDnlO
oKK28lt6hv0PiV+BRIKX8sRTwIfCUtp5fz0jqj7KruNBTU5YiBXOzjGt6lcF7JM85yOmYRtS7+/w
ak02xnfEGCcHVyykbNHZ2k5Ot7EIAfPMHJT1MNeBWntkTELh6o/NW9jkO0Jg3ewBakfabzTAku2x
I/Ud6KlWEjmvUHfWRESaytgWJd6GLyp2qIvppel4KokbEiZAFHMqSITy6+UK+rYD8Hf+hWpz1owZ
yA+k03X7dlMOrvB4Po19++PYVgnVC74CqDTBLuh6Ob+O1aqfdX3Qam5Egx9+7izUUfC2Ajn6DFNt
I/Ip8ZN/TTguL6R9erYEhdrsHqhWUBb4e0eZop7W3GgLiLRsZelVHNiDJlVmZebAwPlk0o3LIMH3
gzhCub2Z98gUi5SBJ3V99yPjlQ0jlK+11ZYeO+yVvZuKjE7Wf834YJK20O5fdpPP9VJOtJYe1hub
LEgRcTHpEGWvy2z6gvJ7oh8ghVP+bJu5GNQNnVB2LQ1eL7Xusm+DrXTYH5+daVl0ec57rqU/HE8V
Ubr+4Pa+vJCy6+zsEJYNwaVv4XaZhSz67tEIDkxtDkRzh7LZeMUjsVl9UXb60unz6MxWcJrrCbm1
jceptMiN0EHjL3Jd1BZ0EHuK49M4I2iK0r4Sy8ZLGhynMjd7shmFWpWSo7k+IjWT2NVdaEGiU9hW
LSU0chRDkN/mLDtcVkysuwlAEPjX/CbfU7jdyFU+o6JE4ZsQ3RBx7oGIm6tppmdRPG4/dnm996Im
Vd6190VtHY7fNXqSq1TGLSpKyYRppGRNpGfW12iREjkM1xXQJmLbneI2tsd3FNtyhVGNbhuFBhS4
gL04kTcv6j9e8DxqCLBW3uZrFmPuGxAR/vC+ZnBO+NoXFm0+NuSMD7Sx58YeLb45anoOeFJZVWm6
O7W0N/t6xFRNq/wW9OPlqn/2ac6TxqtCbEXMK5a/ptIl5EQksMDW5HCOmojX90ESUZk2xxapfRny
rE3+ti+G7HiwMbBiduISVwaSgvBrllpfCEfpquDl1JAt1GA552tkmoQEvxZ/SD3GH9SYLlz3yDkS
ey0tyPAmaKqycbBmVOZn45f6iJEsA9OSWaH/8rMgfJLwUe6qw2VckB+PZMS35ds542fHudKxslQh
ffXj4BGafS2xpCM5x7h09wbSw+zBx95dnULFLYAzkXhdXDnhVaY8tIL67+cfD/gP6GT1vkGTDRQe
xa9Sb5r56zAd2CHfcndNJB9n4MNE7BbpuMy/nFBDAdf4rnRB9FGokiOvzFEVBtI83ydLiA1Bn5oP
iOnPbgmD5ZRoMv4hXPls38WlTSNKMtBlEOJbltdKbziYkaPT0zXzUBJN6nnSKudFSCi9FsonZCoD
piXCeIlwfuK4ZdY7IuhhMSvHg2coSAid1h/ALSwx0pm0VCq9F0vx8AIDgQ6fRZYFlaqDZZq06tVf
DkodJxAOMRH7oVugs7pOQbQ6FfzI9X1x98F+HqAMq6m+ttPswADbNcJOp3gqD2j34ftRcYS6vy38
9I6knhm1Zz6TDnvtzD596oNM/0jRyfqea/3hbxZYZLpGiblaDju1NrXkWNAGYDEZv7WY6COvFz6P
Ff3KiMKxPOCJuVj8EH6W/oQMTBjHHrlkyVv5O1Px6CjfZ1rAwXmUsE5kdcmlZZljENs6WO5EsjvZ
jwpxYh9QFSvSZ5vPklvt1WN/n6aon190w8iiZR75mn5QNUyMlv5kIjynTq2bZOX74mebLz9yUyxN
nNn77PE8kGHMXgtEbuQ0oTEPEZz7wmSVZF3su2Cu+YBRj+M8COyB7bheJok+dpm8aDH0BBaZgwSO
/qmst7lDoTP/45aAeFJfSKlQLwOEVuC5shD0+gwRFdOuTu3ecNEyF4DmcjsMyVlcfbHatgJPwFV4
W11Z5CoHivhn0TVlFZolCRTymzVc2V8YIlGKCz8FPgOWz8z1oWE4WzRUK85SRcsVnTGKd9F2h6RR
+cAZKdcm+zXIZGnXUowK0BQUuWxwacNol6CzGKXXbK0xLStY1nwXdyZZzfvx2PXYciwLD0eC3sz7
vVPZAjoS0EAvj5PRPOnb5PgsJAtIDjPbgcLXBNlWtc2T0DoeDTiUbEqozsPCrY8D+sNhiM5SMonB
X3/uV/jV9MJzoOp+uaxzWvEpUExWrEda6r7XRa/TWo2ZjAtTpnY4ncNmFZbNgWaBHAqzD7BQKQ8/
yPNx/EZQsO7TgQT/cicjjjvebbUR2b1+mxyQUq9uihp0nnNcpTC3SBAJewLItSujHZVKX7UOB1hV
tVs5H80N+EChm21qRzDL2d2wZW9JFaEPBTjaObhrjNpkqrCJYejcmqHyE8ugjsMSJnQkZMbQN6et
PCQ+rLrIvlC7Hl+WzwWAd1fX0B/YKPYIb6tpU4CMYX3hsW1vLSfRiXysuHESEfBIOa69VHoVL3b0
ZhHWCngOfpno3OLBMo9DxrNDhlU/dzqJtRS6ktmau36Qo6ShmOPZZ82+4/lXU+brwv+moSc/7HrJ
rtq5CZ5RbnWN2eUnAmZEy2i8uaD+/ryH7cj0lwO05L8zIlmeY4V237IU0kNvp5VJ26DvJb62plO7
3fICvuOXqQGCQ5DVkW2+pEaMW56gVWxJ/lazlxhf0fCD2+nmU40xFnggjKrTMLYa4+6sOjtg8jJZ
kX7FidlUtKLEMiu6gM2Md7Jzj9y/tFevviqdTjqDpscmC4LwW4xzxDyHRtpMpj2i+I1tUifjM5Bo
dzXfBngYwRMswT/rlOV8zyRpqvCxQsCfd4aMTDBt0T5vB12aZOMMqjN6wLHo6lXzPrUDh5EM25e3
C6WuBB3W9zqmhI2d4w59U7age3U3h+RZrxfhDCIxKr2axket0hYMAtZVXnye7irxmxkpjGHck7wU
NnL0FTjydDU/Za2iLumc2pdTItZde+/e7qJcTMXvVxcGl6dJzmo+fbZwSiUWu1mTFQL1Qa9Tr3yS
MyL/oglwT36KoicTypxWh5s5Bj8y/uqCpELRus7KnJmGY9MKoFZHBOHXGPvKVlZRJO8WBXBcSw/l
Y29Mkpwycf6D/4gJFkHLMqRmc/s5kaYgG4RgU6HRg67//EHFb73cejB0Nd1sCY5C+vn99mgGGOTd
Omu/CWr4dHhmHUH+H3NKdOLez2Yx42ws3Zr0nNVmhZXuCO62dSAFRIkb9ckjLs31Kalkm0y093V/
IUtyN0rb03u/H4Aqe06RQwLgatjdTB/hteWrA5IsWN3xaIAgsl0S7CB8mRecdNzEsyYew0JmAmt7
75FwaTM9zk5BEy9/D+zSjfzUmZ2t1HldXk7KLaY1Dq8IBQcz4a5555nakRXBYh/xb+NmUDMLSkw5
br5xuQ6u/dcTBuxxwUyvrfDJ3I83AxGWnDBe1riu9LRVjeCGaMGMuRzt3Jh2j5KN7w/vRBUQoidG
2VoFQCBN1kyY+3VqAF4n2mRKw4ULSdGyEKohttyM+9r5HReAIuo7pKSUEcd9XiyNdCRcM5rMdDTP
xzDitcvlLDq3//4Z8I2CMpnngG1nq03pFVgKcHpWv3Mccnr6uQXwmLKfr2zlMEHsRcESpqUBy6O2
8sqV3COTCNVl7/TbemmPmuWEqQBLFkeX36QHkQ5Fgo6O3R829RB55qy+2sBU+FhuGjnJUqaGse/a
ouKJzlnyyr+eCH1gp5zgr8yRq1WUAkeQfS2S03JXjc3lhhsHPxniN61bB83GN0npuw8HLyjYugqV
fRMNBU0Y17kq2Puk17v1lLs4OVRhr/D3Zq0MVv0sWCxVjkSQmyUevrtG58SV3bFiIYvflafKAhGt
zHMHSUc5jcpxn2Sqnv+EUZXRPFLhK0I9IuUAlhZKEKBaVCTG0DmIDgYHCAcFgt2WFdCEgAvfQl8k
sOhlf/EtQXuTkz2ha/oZwSivfJcmJVT0hNeyrorgHg0DyUighny0+MmYrRW7Ti4S6yrS2qi7w3yx
43t1dZCfPE+QFgBggEuUfjdI8Ztja++03fObmrEpNdXAdLxlcf3gOf9dEy7Fmed1SG9/Fm+6Qni5
KQsoWOBAjagGD5yb/qwv2Kr7SOKhktzIn8DWZK9yNw4SpB+zdLLQNzW2XnsE4mAuQm/dB5Dx3512
WNOmC0IuL3Ff2uZdFf1OnzwUsK8XEIsoDqhAWsoJQPadIo2ea72wY7tKnMqMxP/Kdd0PL12Gyj7v
eCCxoNI0bteGQK3bu70QNvo9rDBtDJ3AiWMy/gBf11T076Iiw9LMr4IHpqUd4EIkfKMOyQr6bT+N
yXHrwKd106rbTpAcUzGjd2jZovzdw/Jiyx4s1lhrIZT9ZdJ7kM8PK9Y/P00ZLXsHYdgdpOHm4ueq
Jj8DXZYOwFvvwisK82l7qesWzYYe5gcV02fuOg64BXL6yIu5GsEhxTBksaVxp+eGxLV3E1rhJ7fX
EJ4QJ14psCZdUcykhdM2zsNsjw/iclAQLBzWtfh/OSkXv83o8TYW1aDuovYMB7r46t9mOCj+tju8
H8+7OWvb/c3DKp4atsP+nlCwqLq9ug1Wsal+ZSrBwkYrCdc6h+egsz7OSlXFXQ5V3HbHTpZvs3pH
YlPOqQoX50u27LVgVS33N1IYSXSvzJu5f1NH9pfK6BopmbcUYIa7MrgGWqH0SzTZ1QXfaIt9JLRT
yvep1CbUFT+1OblDZvZUujg6PkzJoN65UekLrsVYrfDNPd8Y2RcltpQ6meCo5QIVjDBdIJ3xgarl
sSgC0H7p1w0fBZeYsmKXysZtRoDatmNFYWhVMaIMiQrSIQaamAp+uQ7ZTsrorrXihShIFlYu+uYH
/sC3phl7RQOTVNKYkC8rIujfhsX6dSEua+DkkBYuMr3T+QdHzKbTyMatgUvOR0niJCeMNPfV1/kY
7VtQ6yW4Kr6JMJnjWToKQ4AiyJEs9eMoSBpkg3nqST/G288aaePZ3DnvvVU8gMlgVuD2mOOfaicz
TTe9JofkLOhum/vooGekz5lRpGGD5SrS6qwKbFBptyyzkB4OwGbKFt94Y4dxhm1R5AJnpLMNpuCa
j6l1oy/FFQqnWXDiTYwZ5N+qqu2gN0WK2fSqAuHal3jNJlEkMpRHmsw60P5ETJ+ZhlW7iQGYk07d
qxQ1/T4rGTxknnteHJKHc04YYvFFPwmDfz9m0PdXelpC6+E/NAcLfOINy78/es/2Gvu18OIy+7ii
9JRFifMuw3ebBdmf8z3/7nq1pDjSzSAhRBEuafrrzN8OfjRF9xbF0t3gMG9FB+NgCH8Hu2gM9Cx0
mPv930JtD4/EEFZG/r1x4QDPBlZpngCKaLV3vBk/JGln9XT84zF3UAFtTxF88j9Z7cE7aKAKdR0b
w7i7zZe99y8tFAgq2M7IxTjBoCgt+rWIsWsvnhgBA5BZ5V60IucjkunHNA8Zn5GJe4HgX/gXh1r3
YL+zJSXYCIYol4T16VMUpF1unOq5Q5t9ReDOS9S/AL7NT4uCVBGp6He6MbQ1t6kGbDnFG6ZAVfOA
K9ZSr4vWE/Z2qqxBgHSsUZvxVYnoRXXQ45mN6X+/fScA6TysRYiaiu19/Ms0rJFN1sRIoodPzLJn
d6nlxuNggkuRJtUkxTx2w4cMK6X/ybAcp2A/A21F8Yy8b/c2Ge9Fsw59btUFSP/45t+9IdjBUkbD
1uR67eO44md/IXYDMKnZcd08jKAghfr08Wfu+bIyt/FOBMycguRYyLhMvc/NDhrF7RrQWhLvDZIZ
HKpEWNlQreQXuDhKvo1GP4FN80gsIAfQnA/aF30jrs7rBWmjb9sng3ScSmnk3OKg5Qv4sqF6DdHv
HQCxqpqHtZHWKefgDg9oHy1G0E56Xc0Bz2vzywnxSSWMBcLr+RS6EW38gbWm8zj/KduHOvEzXB3c
NXVoba4jlCDEc9r5jmlZK27tuP+IQ5W8EcV/G5e3Iwx6HQfdgdabcle9cONgCvoy5R2Vnma4R8EE
v1rCuToQ80DlqoCY5btNDvlNS1ifGp0v+Hlw5wyxt5BlQNeie6GFsMe7OzqdQeQtXNOo62mHvJ6b
Tm+rDhWefeNYM+kTCcbT+V5tl0NzHFYC1ysxiw4/hmLI1a1wh0U6Q2BXZcl2TW6+InfIw//POY+Z
bSBtsZ/2wm6uGUHuGMxO/O1HJRxTGxKY4f2FhmaZH9gpJnuej++NlP9ZhcVSQo9+jmhGzYBIpKEU
+cIFF5+L4tlfqfcSERwo0UrIVAeGtdOMHSURH3+zgrl2ULMSRGwyCXsB89GDppEIp35G6LMjeHgj
p2fhWjLgV7PYK104O3TgO27COI2fKLTOkf/QJ6/rBBMCZSizMiWApGbbwFGUhgUK3czy99hF2NSp
n52iFlPE9Vp3W+TVbwXkEd84C+g8pu7+ruWyivtbjWd04pMXzGCaYtZdr3nmBYMj5ApFoCLux2b+
dE/3GcIcVIy4UpnBUjddhTEat9uUAFiMaJz6q1YwWlcYulf00tp2cEktdpaFOX/kMpg+DS9WbB5R
s0ARsc1QbRVz+VG64UBDgpKE5Tn57As68f1hzhbYj1g772ViIzcL3BxtLrQmRMCLORseXvgG24ar
dVF3Wm/s8PmxouPPGFXkDv988fSq43IP8UixxrgHow1tmeAHa+l/18EIQ3QjA61ampNk5FaSjTtE
upOwzM1QXVZPN3VrkDtAJd1aq/YlIemqF8wD9e/2hL3e0r+Sj2zyHOrk8QnS0rYWiqaEUp+2D5gR
vs268RGxyNznNU5u8pCKg1PGVMwC8PyGDivoNwDm2BMiiMw5fNAzLj73Iszc1lA6kKudB/zEuAHs
0t3sWPiwuc2S5lSxklaBJSmUtAeXfUGZ5cAlG1pq6LyY6PO6HfZQjSXEXpI3fhcWzkW6ncYMLGu7
lb3uawKL6fiU+gcawia0oSVCCSj34Z+NQeiKU4X7dLO17G/kFU1kjdZVM9a/HGV37HFpYA+ZUe/u
N9eFvV1goDynfmzY0wzNGhcdB4DnOEq4gQht8t/SiU8X1E8jY6aWcAZ/SlG1lKKkM2B2Y08ByX6e
L+7AErqYxDujkrT/RC6q/eAgOSz1gw5OdfXOzsFJYG3c7DKxDoXmk5KbjeMhBDo5PPGAtC+7cseb
v6K8c/QAIW0NH9yDdL0jTP5g0DDCgpjEo0BJKInlS3vIcXVEE62Ubq0DQOj8gnZoBnZJFgNqjQtY
voB8jERA2CCbkVP6s8pIUkIO9pzDbUoXcvbx46QNbNdzKLUDLyON7kLMGgia8FtAUFRpzAcPMzrs
6qJJ45LLhknUvucli8RlfPT5Hdx3SNyviGKgQ3KCQraMGwaiIA9pF26323tgQTBGHt6DkX7BSI5W
GHl06xECMA+55usRUsgsozVYDLK+rjGMeC8GNQGJIoz6TdO1U+CB5UeLmONUAQqBgRDg3e5ph3QA
8LKHeppzSznTgJVYXED5IeZLDC/cTZkFed2kVF4atBRvvTP8etmzYHL3Ok/s1h0sfZ+6sX/lmmSF
+mNm1jt+KJoUNhUrsBlcFqSiRxsIE3LUim4ZpiAKFA9oxiR2fbkXP3PcsCJEDVjue4DzVtQeXngq
g0bAmoYaJYCuRT4eQe6qhGTElySFgg50pb15qVVjz0hIUIG+jG8i2khvW8iqtk4ouGwdGr3JbX79
XxYJZhr5XsooydXSNMvduxBGB0nnR3JrsX2wtKRQIpmEzC3DOC4cMeFvk+0HVsGpsPOGuZh4/CWo
b27TIEk47wcMUmxcJqJFB1m+Pj28mPzRBhp0P0vq/U4TA4zWgMZEVYXCMUru3G3U5RuA9o5n8gbl
PHR1TfD774FZzcpw5Om1ekPPLTeHCDa50W2GyucezjguEJuTee5De2kIBVeU0XAbixR3546hyeAk
oWCTX6yvQumvZxHwFyPR2p3Pke2gaJeV+JNrR4F7ndvp4MZEM8LArplFth3dd4oFIWGo+DZk+LVj
S4oq1N4kWvnSbXSn3hpAGIdtL01rtguzgyUp2Vd/nUBUntVCMoX2W2VLOTqL3zQPEHlXSnBgPfjH
qffW11rwlr962WHU/4t2O9PvGfTCwmAjg7SEWk2cA6I22lBGlQyMaivUcFKGNSJwwgLFh/ADjSnw
GacJz8E5xlbS+klW7ASac+akaEukIsu7por6Vsyo/IgjRm8dvCaaik6yOV0mej6s7fxFStCtfltx
WsDTFwPqrLoiEodgz7kDfnWelWLTAhJAwkWxNFz8YST8pWa3UUNCyErI9CIfVwuzQqpUctNeAzMc
CPnfVKdTtq2WBeuA+W5MjN3WjkDsaOZD/8sCrTfsSP0nr08z2DM82GNDfLraOqxo7/l55STwkUMA
NNlKmVjM5EbuHufZ5L1//Al4evSmkWpf+pmFQnNWSOL4xN9giaoevT5d1OFI0g2cW2CUSwXDpnfo
yMq4a82uRh9b6rAT3OsqCv65OfPx+0lAtZjSpfAqS16KaXMRoTEwwhWzEa4av5N/CEcGg98M73Ih
O4TF7F2QJZTN9S0OSO/BGV24OOaidrOvGZkbYtVjCPv0rxzJbgbSncdQHWP00Z0GmDgZRfGI6Smv
Gps/KgWqCFsrM/aSvFyJwO4gjW56/CejlZk/g7PSYAuIXaJhl+TY7tkPTGQOu4LkS+FIuVzqoXfo
qzpeQJ3/jXELMzXME37U6/XBeulLL/sVoBYY6W5q1GnXDnHqnW7GOYeTW8AV054jaAe7sjZ82gu+
4ooAZR+idh0iHOLNCXqWhlCf/4equuKjquvCCicuZukBJ6sOZeCL+Zol+RG5RK6Vb/GsBcLmMAT6
RDo4TCdcQ7PEWASlLNKPzI8TqRXYhiotltel+dGXVXywb+Kl9RQEwfn/T7jCsuPWg6za0yVwlVMl
QlYoShDeu57zSLa0ewgMJGzuGnDIvtQG4ntoiiAjcu6Q+d9oHRD+tl5trW1thZP1EDwkDJcPl51q
IkCJY8Ik9aoyO+99h7jIUMvyHPEkVNqVWOhjtQwGR3wi0b4PSgU/a+yuFrLnj9iFmiVesK5ZSxH7
+xrYxXsxUCTR3e3UbfG9ACffGpgk65cRlrBieV9UoZwI3nL6e+d0PukWyWPIjhI9e7gRMUWjpVkx
ww1A4K+ITjJI89hw+zZWeGaZYEqsqdulMu9ChOHf5MqkoDXSB4PhLS/SlglLunXPy4AFwGUafbLT
RUvfvH+E9ard2PnYv01ddNfJ3PYu9etdObd+wqvJLAtdzF5FY9rkLgbhPTaV5meFBlrPqsGvxo+7
+Vv//KuaidnVyrvxIAIMZMIUzqV5VfsdQtGhDCl8R/0zI/SuQs1PUlH+JipUUHpyos/jkYyBPuhu
yWxIzks3x6wvGLeZn4+MXD+/MmmaDX2J7rCEKYRQ9NsMLApLh5VE+EK7DTzG4i7DdaABCBW8wu78
pdLF8yKQAvZZ6kupx6TDqqhxh+h2+IvG2623PwaUuN6CImxHbsGMAgrrECp/YSOhJmjvNDn8CloG
MEXKETIhEcO5dcYGrAr2kNiHHFxdQmuv5kP375dEyYNr3f6kZqnmLAXVb/SByAdTNIloKEKFo+9b
V7kT5B1eCWIF6iNhXvbpWBWOrRqXqbXkycNRmNQ7X1Hl9Pj+x5xe4lT1FdV6CNrWPcD4Ya0K0D43
4C4rdRfwZyaRKKubNt/R9sbk8exa9SfMI3Qva6z7YW5B1okM7rGKE/8BM/uT4+SkhNeauW9KVPzY
EHl3lBJGT2lfCZSQX/NUayMQA3BDbo71KJGgUCAD5AhKHYj+wwlPfvXscpXX+sVEFkAR5hTjuW3X
ISMOUO8sFHkjVHw7zscgQjd0wgsWm2cBkTwINHqEE9bksOsdpoUU4vW+Rd28erCwcT5XtQyPJSnJ
51t+KrT2ax4lla93Dbgxm8pGe+TDFgXttyxdmCRxJDJv1Dd7NNLnUFOBBR3OWTKuEFFRkt4Xc82C
J4ejwAaYfoQKXUrOhiBFO8ghElObTFsxzhNaf1RovkrQjo2uVo7O6OKoN3IDa/oBkzgDnkYH6zMR
aF4+v2P+odA/t2qDMENHBY4qoPYP/6BqdznQKoa3DpVl4ceWfxv/Qs3L+NA/128x2/cFlF91GAI+
7LH0cjLIox4sHK3/F6a919SgW/jtk5FGJx7y+Zh4I9GXCI6R+vUGfmsdUj0uTAQFQPAuis5j2Kl+
6hMyQrhxn8RCnAyva9fZ2Vb+miI7ZFVF6tnrG0ggVH2vaPxheQ0KCA3rqt18A/9GUjWNNcMQh3WB
DKaA9xR1M+aH6wbRwcz83wuRT1nJVQiD22aK6LgH/r02VuxL6AlaMYdGhs7cAKVQbxfbxE9JFhwZ
PE8KjIl/4m6JjUUI5BYYW6Sv3LqTxqaUiaH6oeMOXAmLpg/WavOjgNU27N63+6IOB3Y0ha478Usf
DY0Hh6cxe+c+Y67gn9TyUnkiR8Ui4ubMfhTnD41LYw9CcqIHd2Cjmkw1Te2MhUTllDCM9PHsSdin
oYl7rOcHvFSGhJiWmS8wy56FmpH5MxWf4AFZylU/IA2lUGVoGRp65m8c8rJ1IqDdg0TkrWP1hEh3
3H9fxjcbxOUQ1YNNvLg/2kA1ox734l3tXHXgGc2CD9Cwn8MbufbKjWzO7I4/WFfNwh1U5FeoRDKl
26qPiBSaXKQcZq+cqcqWFuNolGpCxHFNH32towh1zIjyKiv3xDa1yLypM6jg6tVoiyooPEFgiidI
goiEMPsvybfeKd6tX9lv2p2EdKZ/+pRjfioucgFyvbu+awOADB656X9qTjRntIILVp/9PnLxmXqo
tqIYOYBla25t4Jn0Hk6OcepV1G0VSVbzEU2DKOa1yEirbTpvNI/bkL2IceWVlkucxi9e7ZPBgYkI
DsI/3ODJtaR+XE3N63nuAdwesDHOX45EqM3HlS33HXsgrgj1H2ZCxspPET277u2U+mwO7DuQw89q
QfR7sVtQoTfoJCsJSdmLbG0SUlxWdieMQ4gQajSSPkxFC3Qd5mVT83q+whJlhR7o/FbSomncbI2i
O+iSEB7yJag1QLUdllVdq7VOjUxjF/v53XXiBx4mq8PtijLRH03350mGwUGRX6PNHJhY/9boxO+v
rhsz6gWuSYv7/50iytwPGmYhTDaitRALhyq5TsoTBRQt4P3mwaX8wWxxLgsZX/7yE+jIRi5lblYP
nmURUxJ5Sqh1bCfKwHBSxONiCeqkzzLuU7nYXrliPAmBo+WJtzpzuEgKrQ183pIfM5v0d4sn3gbl
YEuwJloaRzRmbfMLzy4VtUXJYXJ6fU1DSRIBs4uPHlIpPppf5o+sbC2BpxIeQhmZW2eThEvy80IR
60XCDdJfKqMUQj1U/G9E2/ULUral/xfvWTPdIwgvh7SX7B6999Kh8APdX5ikWGNYnUzv/AJyBehi
9Jxb2qCJB+2CbOJkbxaHlop3tYADf2+ay1PIjZ6S3QUiJg3W/Cel1a7/HlVEagUApS9uZJWy/bpL
2lBozVMEDlycGfHMeJNkpHAhEnY9+VhMW8g2Qdk3hLzFMG5cdtdA+xy8jn94M9Ssfdl81KFPcYEW
+0KJiCDvi8xaKmzo9yZyOPfol0yXLBv2ub6GXN5XNZZ39IbcTMcnQ9vVpgH2nA9QG2dbOZ4YDiEF
tWWRZxQYg2XUpX9HvG7T735bP3Gqxloao4NCTsz8TCJDzhZ04BN1wUHSdmGVaWv+3lLPu8tRGL3m
5x8yXbDbKDTXV23enVa+f4bwHq5xiSTyOJ7pxM+LArIMeSSrZhNClY0MJyreJ9IDCdIG5294jqeX
mP6elscWssXTugXszvFzB2wl6g46MDKDlZ1LRNdM4sXC4RXdiQ3vrRWIHmYoWJzVXyd6TlmHLF71
FY+q6JvASv8lXnbJ0VZ1G1fihOpvchIyCj42O7t1vDeZIQbjZG2MArxCLAG4k6Z2gHGCjF07Yhw6
iBBVSDG3MbzCj6qeZM2RhCLKr8mL/iPAyt1cuc3M5D7Zlbx5jqkT69z8PpwnyIuDr24oF19x5xKA
4wEdrGIIZUbT/hmrz1wJdSfpICns/TVdRIUM35r17jRWfgltw3wBKJIxEHiIZeuSCa9viwXTe7rX
n8IEOYegx6NOu0RXhksuXb7VQhOQsL3zFBoZE4cBF8+fs24MT5XsUKONDii2XoiXs6NmUf9AsNhx
9kpdT8896z4bJcAIPbYFZk1l5A6/Yv3jQ4pBEVHsk45gfGHUVNekbpOTLXZs7SHtjrVYngtloNbG
HPsUbO8JkBLsuXMII959q+LCrsaU60taKYFugsgsv+roDGkz7NXXSb09g67Ja7xYEpT/ZC19oOvw
ZBudHaXyZAA0IKHvdq02jvnZ30Opb7B/AVPqwnKrDMSK5irD2bhz9a/LTMPlQHJ9vGl3Putp0XFt
fQQE7p1x0niW5eBE+MzxkoHp7Gza9dcz2NW8S/tRsCvibc9BJ+gnhT/hgxzc/B0pFh7eB+fW5LMt
Yj3PsE/4a+3FCPuhZYGK10m7jfsgx38x6pNqiheZzenVHuV0XhZVQ3g1DUpoNxOkDfz7XZDvsOsh
rF5St212ceFQY492xfOqZlm5t1wXsWDoeY9NSmYE8uT1PM4d26RluotHgppkK1OVcc791Cf7HDnX
vZdgSswXZb/AoPYO+eGsNlaaQVoHtHVOW+mLgw6tYTm8krTkjkWoKngtuKyqLV01uhdrEMwTGwBv
v/GJUuylKk3ns609RDm1yxxE4DuwjF8Civmtin1NzDz2vxeu9ckY3gYvJFgNZCWNDqwRKnZ94F9U
7lo1oX/ynlAken5Bgve2eKf4pJnAUbAjXXlV/ceKtBMp1rimefulIV7/iJgGxo7LHDhV5eS5TEYN
b58O3Ml6YVHmJLnyQx9DU6F64z9Ff3/UXOWvzxfZbyywpqss1VAtK6WObZgg7vHwFqlUHXx7peWe
jma7sNS730chDv61DJYeYhwdak5ADYn2EVvIqQfTcTHBKtgZKdzZStIitgk2wPObF3tl/gT3zpoK
UuJYnUeODfwT6oC26cA+dmiZLRpzsGvkq9XHFOqBudUSVXNoUIkUEHebcCCfZURml7Yqr4BxwVHj
3g9EzeRE6Z6Wa1fVkwdEOI/hxNdlnz7hx++DdjwSUNDHtPgZVBEjxOLeTLwiZmDpATWLNd8Q+x+y
9TmnNE+nbtaziTvhvt80aqPepi4d01kekNBTnm9irhTK3sY5TnjvIX0cDlDpNJhLCuxz5BiDUiUR
fHwk3K3z/4Be+PIrveZv5952S+xrGFjoZNzAcmUVQl/eI7rRe4LYAw7dnvDW1bVu9f9uiWsepMMe
cesMZSQRfjlraQsQg0jh/wNKhYL+epDUov8qqhvANF6Tx362G9I4L7uLp4S90mhVFRjhvEli053n
jTiCg3aFv33ANia9XfBvODe8iT4KnXMDeLYgLgfNNfjtsPBMyczgY3+DEF79o0ZY0d/pO9dVdGV8
BUE17G4Y59fGLqAU8MN76aM/qAG/+QrU26ZrIlnMdX6t+2q5TEZ+KHcBHd5vyX7Wwk1fSBatPi94
dcIsF/ZiVx1A/p7gL/0tYG0iIaDRwHdRRtjD6J5xu8f5QbEXljXV/x+TJTeH3yUkMZpA2qwp0gcO
mWfNAPTcCQxTD64gnB5JB0US/Sq1l8N99R3KNetHmETzYRld/fz448aQIAfJuiz/Zz6La8M3/sw6
wg5CWAM6mwt68WJBIlYDcW+5/uSSYCVkqZWgRhjvmAFPfXXyf/geWxpFaTcXLeIhPQUGxTvabjQf
sQ/ntzqc3nCvEX7RTOP875itlml1IylwlilWd1MBLi4P0mwyKYe5pYMNvSD6Jfmd58yBnwN9dmgo
sg+zQ4FxFVey/jajD4rAc4EEz96oIn4b1bkvBQOyns/R6Is2dGWxSwNxF2lwqchZlpBtVUsz3ZX6
aqKFYKxs2jkSeby4HQdRrUwLWQQGMmJVAKuJDnoD6ZiA2ONg0fWbCirgDno6KsAALqusG0r70svO
0CD2daEsJtHml3bFiGoG5n4vUVxRss/8VvDYrmItCH6u2ACmUtOfafGUFiBCr20Yqb3QPLnINUe/
DHgKKTM2YKckHugbyBKNL0SH4J64VFyOVKsn12qILd9wUinv0LefJqZQ043ht7Vfe8C9M6U4Ejvj
Uq0Z+UWT2Gp6VZHpZSRrSnHmuWgkJlFhasjCUlBX04b260dgpUjYuaWy7WNUl2LOtVYc42xZTVCW
VA+au/q2LM+jPLZ6nB49gani9jUv8bSswq3f6N7qbUCt1zpB/rVfrQBMPpc3Da+Koo5rR5HGskqE
x3lrVADNGKjBuj/Yp1hffm9znHdUfOc9Cs5ZAxvVRl9xOAR2ij7fGf9j9BnUPYsRePnBICkt35Oo
Oakd7Um2y94f8mSC9gH4wM0O4RNJGlo/Rj9HUsYjMsphgu33duLR70eh1raUz6t5WtJulylX/7WX
/Cj/RPOWVbPGxO+a/9Y9+MDEPnGB5u1X+R57EXn3d63MSr3CfBynVwecx3eKAVLviq8JD4ptn/yF
1IH4LezCPNSvLFuza3RpLRw0hb/G4xe1UhUatORpTRdoJKTUt5loUHXHgBUGclK/6KrIalYjMOlU
T55NAVcOSldbTEAd5CGW3yLql5OSv2B05gsFImf6D0r1rUNk5fwuNUn/pjna0PrtnkAduyUdqbGW
TOTfvu5iXepNEUCdWJ59EUCYxakSYZIkEBr1du6hHWbLj3qteua1XZxBoEp7pXisVuZz4i79PNsX
I8LXrFP+O+2P3YyamK3Fa4Eb48AD0C9sbhnbwH59Y69Aendx2s0DxEIH4LNdZ5Cv8GTajrTX57J/
7v5OJF2GildT7qAdNyTkqt0hN+V0FgAA7SxhSVViWrkM6YajOZ/IhumU+ArAbLxRyWy6ZSeVJcKG
TOqSyZwZQC6Iufi2eu9AmsPzhCvgMqLahIo7OCPm7B4ZrgYDsKwleqC8lKqcjcbHGH2vL4QA6zRO
KEWy8htPli9F072j5b/m5dZ0nwg3XynGVjymR5gqc2HMCbCwxDAUcQd+Yel9KZ7ei99g+hGOgJ8G
KEXjYnhHltwURSumYgaGAhe76tbDqmkDjcbbLLhQpT9xcBjtFt2QV50hMXVbj84eOcYyJFqxY9l0
FznbgVDkmHyBEgiMkoWlwRUGWEMpOcotcFdXyOTMdpVUbmMmucMie0F/6QLPhZOCHvu48Qxg9L3N
qTnRy8yglbalPBy12Pja3emKHWWqYJ4UIRhNOfNoQogVU7wJEaMd6zKkv/FyyVGt9vdPWe1a5jKF
8ufSh/T2Y0z04L4azoZGx+X5c4dD0k9E8EG4HKV7JRXoxr6mwfhJfqMmsploKvaOmXHm2bJzzftZ
uA/Ne98SmTosINkIiQrqB+uaM2fnKoX3QI4yHAJHN4XZk1EOQ7sc69lRBfFxxZIc2vJZuj9zJXtX
wi2vrtHfzcs01rwCF6uc6Dy0hJ55ddnX/K3gkTvxK1ICWlc+kWzhD0fNL++kQLsovkERRdIxD1ld
jq3JYvrJ7R0X+MtdnaSo8RolNtbL5WRMfMlzwPJN+pvBH5qSEUbguJQKMchg5dNd/TqaQX6+UHq4
DVtWl0eln7TLTMU1sWz83jU7JR9EcapX5jVexf47aa6/fI4d4bm13/3iqR5CBVdaU8pxzPTHXe3e
z7ovdgRgm9zDbB7HGouRRYB/cErBwVbY7qntspXb3gb1+n6mZE8Rcv9Dc3RDBXvEPlKtosUK0Kjd
fcwej9zbznYpLWudJbX3jDpTFwnD08Nt4PbhvYO5zG3QxIOqyoOb7bDsFFkBq0hWVinJVSOSoNlo
Y3//3MnOE5kGqKYzIdUiSSsR+zFgnGJOQ4RrCw5XXGJCogrfaBEpgLaKsrLMvg/V2r6+xsp8+182
zpDUy3WRA2aBaJ5YqHOKbmyOrQxx6So46zpmfNtWkb5fG2E7diA7oCJjrZ3p9wcaqYpuScqeORCs
ldKkEJZ8W2oIIBEqZPWhKmBRbfoH/uZzF+psCIpA+W6oQ6lTo8BqgmQ+HnXOev2HM43wwe+31vOO
skEbtOdfKwVPAe7YNzB119BYjFDS7ZHCPp8i5OttvGjwXpwY+h7ghtV/0xDsdIciM0VizmJplE8Z
SZvBWFGdoJZBrXK2WtS7b14h6ZjPJuv6WPDgAxWrjiGAtVgATKdSygx4My0BnWElqwEi6cL2HJJt
u96WIcdiIGv39p0fsn24EGqqPZXldabiAchIBGn5bp420bUmhNN8dABco5mP/qcSiTYPpVf6eCWc
1hbqoTJkxtlfd/7Vq72wkfZTAeykE6cNWxWxVc3NZd7LR7NlDYhMEa7k2Fdxh5cutwJ74FltE8Ne
2NzN05HlMRyEqDf4Bzx+eG8y7XnXK8iZ/AQq6V4e76sWrT6FnZhYhps5p0iqcdS82oKHq7/vi+w3
Bj0r5BQuNCTYRvPShAmAPaNl40nAWa4v0lMsaG6uYvo3VIGaXTLsUtbRXFYvOPRr/J0x2jz93UUR
TJz94UoVVHRYbb8hJt3d2xlHo0aA4W8C5jTP5j47aDu/cFHGaG2iIG1nZX9SwkeEKu7+7wcJb6R+
66HWnt4CPZVzsE+dWglkHVwC1PCeS/1imbwQGMhrMxhKn1TrGZjSAKZrD39rqmATz07Zj+crN7uF
6wxu6LZxOrZGemh9uruykoTFkswdGpzqIV5IdR0FJ9FQZaUK/1D3IN1cYTUUEF3Hj0OhnIQPU3A6
MtGj03+cSzcXcthjBovNHIw1yT0EKNc1TaVoNyHbxLx3+yPlF2mqxcTKlmL9ifKcthqhfz6msRC3
trlBn+TwAePw8L9sGDdPG+3UlllJe0VmTxVs9sJA6mgYkr1mI+HZhsohffHOk8CHlm6Ho52B+1hd
nwQqUgbC94KD3MjNHdaJpyc0ABhBVd6jApJUUHI6ay00w8IWQwSyGmHmdMKxjeY3tnbOj6PfieOg
rNY0JvAE/afiorf2AEQHm1uJBGybqPfcvZFlAiX0DIY1mI2wPRuTikT+PAoC2Gr2E3M3u+5SI398
kJjRaNAhRir8+njgeQmIp1NhZvNJafgTkhJZaTh8njtQTxDBcnuE6QR06dFVQ4Vur5d4lDHbbLga
7sNGmTRyQGqDIfCgzXWUg8ItXXlr27mewicE1XiWyfmjNavugGLdUeRQ3fxWwv7ux1450ZjBINfs
0tzJVnUbtrBIhiTzT1Eda7btzZZUp6UTUWiuL9hBomuDw6a/TypMT00g5ymhx3vVnEEFiNAvsLYf
QIJuqB90nCv7Jx07tgvAjoi4V4JB6QgEFObnJAoV4o+NynvAYQE2oY4QGPWX0K6YOHRylhYy9ytm
zqG4kdsNGrFOXMUQtm+++L+XrfB0TpAB5Sc2QkICW2bbRPVxPT4pPTorzXmaRd58dOHaHsPxo640
ayOds4ouCSXo4B7v4GRwYQcicD9GrwkYu6bNzlzF4MvFMCBuRxdreAATS8RGPEqpoMC6dps6s9Hm
zg2fTgjzgyCIcNIdrSn0WZ53QMIE0C2pfMYlC3swoZcuxKHc3Eg9O1oCI9RHu+jq6ksio6i2rEVF
9YNAb+9M8hpCzOXEAv0W/VNtXhbWZdp6ecApRosHQqGyOlypzPntN29uN18l7rj3BmsORHVwT3/J
q1V9ev2Z6IdiVC0gR1bcOiMD3RJZp5Sfyqj1uY4WuV1IcCDWlh/qIFp3kK6hXpb734J9sTUVq0Ok
RG/XAV185mz1GPJBno+z6VG7PwOiWzl6MdOMDM8r2j+RN7XYEcsK9YWlK2LMXKYNajg7SfSMD5Z0
um89b8+o4O72yJuJeXIws3PzmTibwsR9/8FY1kmZQnDb8mXFki2f2bxhmquIH0lVicuuCszjYhEX
S6b/8el4EcdAHIoFQuPjYRNQQL/W0lswvRBnJ6oDKJ2J5xP5v5cEijp06v7In1DLVZlkcRmczxAd
Co/bAi9ZifNaq9SKF5LoccwGhiUiS5FAGiMC2A6uB4i5Jk8eavM7i4Fp/olVkqCJ89/3qKX+w1X0
Bn5nNpYUkUs68ifYLkIObHXANKc9VSByLl5BcjM5l+4RbUOI1gdzN9wgzZTrXshOBBqynQ38f6mq
EuQoqDPUi27POaOSEwwbCr3aWcjLgLOsRbCnJZRhgHcJV0T/ovjNFib7dSqnyMPEWP9O9OPDAJiJ
i+VkJKOk2WQ3ciDDfpT/aTgWDC9SLmCxbmVA5+oPjEOq4plorsHndRs5hzomJJBOKk+4uUgwenuo
Vs//1F7ZrC2BqxCd6q5BmIO/BgKgeSjexroDURHEiRrNKYjLFdphP6j6nFIovXzfc2aTGvj1F7QU
1BwMyDBxumCMD21PN+FyMUwoTXb8Qr3pwiGk3fJ+TS5Ky/uwqyL2zfNcaIzfjH23SwkpUfnLTHxB
JkgBTzsufxQN62ZAp+IV5iqUgzKIFQqkRqdp7rMGFO4xpbZk41d5YhNPWzHRN4IVfp4tPSWO0huY
OpGGHAjpyy7cW401SQ/8VHplH4pyhZlfTsdz4aclMuP+kS+QLMepsNrtjPOELDvz5qX0KZOyTMZR
Lkg99cfSy+1xrLcE/hrv14OBBGQYyK77NmDuDei995Nip0iA3yEpZde1RSQggOI/+L0fWHtNxzfr
qSneVVZckV5YuGiY9YFwFOcRT0vLG+j8XpwmBH4SD4bJdKeYwt1b0YuVmJS3R2MYM7EbGF9yAyXr
0KUKbOBM4xvl6ujUUCPrmRR5TMnBPxC6vJlVlDNapcmQk8+8WaO7zC/2S8QteffipcuADKhaOMqu
F5IjIbQycELpcRdHqFFWqAzYfRRxCG1jx2gxpGGc/8rbU6jwf/hbLVfMbP7YC+vj/awMummFL4MH
l7qgfVPoq1rmoqY+jQdV+vXpkZHQPxLWJWboSqyXAUtB+QYawesMYR8p33dYqj20POoNMu+00hu1
4RS9oiZ82ef9dE5s6J4m2CPAPPdlVBdB7b5fqBFffKqm08WEi1y6G9MT1DHg5ydbWAF+x8cl/ArJ
w3VrNcZ1Tg+m5e3szHHRaMlipSlRU/69OWaUiEUIaa9Z2tIZ95EVLAXlGZQ3vzZbbBeH+Q9JJqYq
qRiudK6pLYFkG7yz1x9MMl9s1gno7Q2PpOW7cbN3wbbzCaOBrdGyduE5T4fRuar2pWkw04hXQ6Uv
GjpgTgVBdxfABHIm2qtrRE0uB5z9K4IKigU67jrHltXMEl5fhUmjew32qg5/w52frxBGjtVzELkz
ehKCqVCIiDBkwTV+oYm3HRbIsVWqIzbUtW6HMDg56GhcByVwA8lgFcCO8sd3waWrbZy9d+TIkJVe
hxPPu/WG8sytFey7Tb43u7UFZIarpA6di7Bl3vY/V/3jmcjNOleoKkvHJiMosx2kPq1E7Z7RoMLE
IHjCvMoWdcysvqcqScOCrbs1mS0A80cDkf6PWCnNFutSGaiyygZK/GeEY4vOm2pSj+micri+GhLP
8caUdIEwUeRKXpxLkHR+vFiH4jam2wQcXEvPbAGE9JJnnpoeEASuPuctKwkDhAKmpGPX4xNWj4v/
kYRbGwVSvrWGZmJv/wpdQOt0AcaA21M/EbADTVCCubGmkA0exympXggFYDnDfjPFX8B7Al0QhMxd
PbEaTNp3sA9MrktsinGvAHKD030ZEZSEJpr1aj5I5+N7hvxeQ7EjMfEeKQvr2/aefdAjduUqtIMa
KEKvtqtOQWK6AqAdlHvr+HUkjguk02CdxkFJJC79RvkKyvLvzEEbHSj1jZcSavn/AsitCeyoK2m4
oAZoWbm1qcS3sYQ9qV6jeAa0uNJeNnQp4nTFjnbjp+zp0DTejl4trUzJFJv+C2XERsZdIJ2Cp1Et
tHR6DFRxGNztKTvyYNODdvIDursGepMNsdpJgf3FyI4+7yEKeLgujlklMpDwroCS8y1n5jewmwMZ
8BFOu1iDrT3zMehN6Il+a+ChilyYQ9uUm9iVaWysi5cbIRVOnJcKmcDx5xmUIQJA+innC0fXNs46
WH/MkXBA3HRIOxLZ6/vfvkgJ0FcAw0YGb1gCOuC5mDnmB9Y7Fb4iEVH5ec5MwLNpYWnOH4+UmTSd
WM4XL44Wrko5CqjcvpM3bl1gYT9VEWQsAmYawwjvaPzVAAmL7yM4hCM9Pbueur5rGCMt/m0kOgin
176YqNhHxT3gqdwJPuPRZIv9q9qHbGe56K2pmJsN7KU6BbPR+8ghQpJourm8MLwmGlYM5r4i8176
laM4+UJBka0faf9LS/8lFLWRpNMShWW3tU+PxH7sOuzVjdSpKc4WxX23XiIs73mHUBXNGQPPZZM2
Iq7x3Go/A9MHa9KZeLM5QhjGA0Kiq/vbGoA0rsLGhysgtadK/C3bUDFUfHlVuqivqCvMTGad/cvg
Vwk1nYmkXqgy2SeToPvihY3JxIR8p4l1y4MirRRVCQWbGmpNmEx2HTaWR3FxEdWS1WUoWuG7Fn4n
k/RkBD+uu2Dj/fdoDxcIWgx+efwonUOpF79L4AVH2BfimK6bkI91+U2N7wwJDD+MjUkkAC8w2kJ9
ckpkbA0vjFMuCn16z9nnnwqT7IEirWCR15vO+sVArkPEEhiNk8/+TQZrwMxzWdEi39h3KpWQfDtT
LMPcj1iEbELAL14xLKnIhocJ3EAbRkxxzvBqJzQtNUiGdDp2D9hlSi0ttp/0lG79i5u/BYIz1Qra
ZQUwLuCbWKkbKuifTZo3LbBgtYakIIbr00yzyby4qsQ/ei5dyPuQqsUPdWfqMm0q8coTJoJv+h4P
rC+bENyYyxfx05vEi3DDgwAQq4nkXKR8jU3mwoqLTUAMAroUFjnVQlb4wObEF92Zpg5LYcwCfD/e
LLa/ZMg9Rt6nZMJO7WrPsxGr1xQO6BC3u2o0rtAue5IV0PUY2gEn3o3ssXpCtvcOLjkFuysSqgwp
25Xq23BsQu0//xBQdhZ8LrrkGwghZDtY5AQcsTnpGWeZ4SWsH4rov2i3kAoa56RxCymzNKj8q+XV
FsINw+otSb0xfI5yro0bnlfyGkvL6OdKcJ733uNsVcZlgVhO39Ff0pIapyZXrNDH5ssyCua8L1VK
mrpncaSVLWqAOWjN0fnNqCsiZajvNFKWbtMRx0xpj5smu89ZoYbVtAliAYA2D3ScA4H2OHXGHqO6
tznWvc6gaUr5kpfKun9j/ly2qa+9yLYeMJPuxpy6icTTGT/mY/08oCr6qKvpIynsItevRMYffS2b
MDTDRS22yVOvzTZ7BYYXIprLzozuylNGcDBCzc/OLXR/zBk6zD+lyWMeWx7BxgveTdSOC2L9Bx6Y
btYKPcShW9ientZR+ckESQnyEUrx4putXuKRYuPsWoTgKnMhWiGRrgd7yF70M1cjddbbXjJzWFRb
oINL21RrF/BUdxR5vKvSABUcqUJYhiHKn2sxxbXekpz2XBn1zW/NwgXAzxY4hBqyckXMMphjNs9u
invKLUW5HR3Tt7B4X7MPLpKeMIXcWmmHzLQOUNaKknemMlCsGLdY4CsIhQURwI+pqkw1+00H+1RU
4xYj03/M1Ogm8ijezXuY3JSydV/2dEKN67naVH7m4agrSi7MBXFe2N2ihfWmolq+21CGAGJegqmq
8CmTELzZGsAijUoMTFxA4KFPhtTLxBdc+EMcTpl2IifOqE2JlHp305Mg3EtesoGhddOVH7YCDvVC
NNhpp7fTaVNIDPb9v9knAUhUgaGIUbkjp8FfADY5cFPf/kjGkEyHTaEqsdJ4zzgn1TXz9C97ZdON
ujH/1dGUd5O7xFd/IaB1jbcefxQXmsQ/TtauyYDMXZ3v356Dq+zkFsf2PAQH8FqN5FB6moMWYCYL
Cqjt2SEi1hVQSxEiVHL4E/RZABGu5Tf/sclILIBVFPb82u0rmyvKtMQbDXs5dVBuywACkcEei3To
paOMIEm8HGtCSQGIqH/cjJAQ5fE/5xFUHNJH8E/0MjZvJ7ceuT41dXW1L1lpQZymSVV5gkmgrwlh
QCnRPzultYWa7RYTPw5NqUxZC0zHFbl6SYF+HDfvBm+IxV9O48HaodIUVBBMWDnosD64Fp4RDCcf
kBC27NQXJiQ4r6tvfmzgU0VrHgKuOGL8WVUCweiXP6pvDDMaTPb9G7Rt+rXoU0mKdzXSMnmoKRAq
pD8EOwmxyDW58XXd3/2rfqP9WeF9vwFLvA5bgAAji/HApsi5yTDFDHAusMNMhHTDa0YpcAZwHRh9
JSAtXpBGcVY7N0YpWh2jg09ZQ6ZRq3S+WuxOUsdyyuPoswfWicJkZaM+jUlGL+oX7O5D4kG23WRp
GMoLhfELEBx3W+MY1HSTQ9GcX78hDc+O2JZCZdcjoIObfpnY+7rhS0fjzhZsUBJMMnIwfszjCEJv
Y6BZTuhFmeWD1Yl263YbXP01F+y8gQ669ZclfGRZngmBDcqgsXGIJRgj6CA5hK5Cas9K7Qgmsko9
KpJpMZB3pWhAOUk7NuV+LSqdFC29rU8GHR9zbFzxyTETlGm3LyTh3xEm2tFAcd4OJeEOcGbJMNVn
IqxU/edvMn5kXPfkqtEckiatGp5dkASIAfipzb8k5V5fxURcdS+AobHwEZsGNW2ns3qRM1oBZ01i
biaaQRhbaNafTMJV/aBwq9myyE8N5UDiLt4W7bevL6+3a96BTdifSwF/IMPwVOE0Cv5QB4foTbtX
tlfVmby46Uk8cm4ZHm1A5yPA0HOxboCUsYiffbZwQMMxFQEow287kLyC5/b5fXWFOZhwd8C7fAFJ
JIPnmRbq0zHJZe7nR6x18rJDO++WXg7MLuNSssT7Ow7czfkMTDX1E8z1YX68dGu/pwdN5CoLsOMs
f83G0UcYfW9oOAmkbssFtlEBlxRK/hH2yGAxJJ7vVl95inRTwHc+3mQuQeWT8EfL54iRnrjNXr58
GmLqtOs9/UUdAlnriX+oRaDS3TfYwFBpiEMOw9vKIvgtsz5nm7JIJCNCMgfqiyZt6NwdMJ2WYd3n
wxQFq96B7ET4yX5N2pz+Y09MEbntaVnoMsXBwbpoLWiG3HDiYTo0ypZqUfakRpC5yxFjHlztLOL0
seJcCQxldGKvV5iHM/Sm611EAeR0As7y1393nbgZ/VqrlPgc20uqgadxiUsS5R/0i1tSXKTYAPEx
PBufpy39d+wgKxhtT13kNI7O+Q9WdTza7VUToFTAUwWGekVZ5PHKaV9Q2IkOVk14xEsvUFLIsI4U
3M2j14NMckY6PAEtLWIRloiyRjdhjPkhLH/zV8P7+Ee534XaWGEmbTZLqnXjLnuVl26ett+2wuTO
5p9/2J53G42Yv2hTcJNGM5Hp5Gs5OCM9cu9ZIbWWmDN96ZJiNnmonr6QK49JwoPJW+kbOt9uplWw
xYRHXYDKJhCse4nMfQzHOfQcxedp72BgVf5x/sObGV50xbpSAu2qX8MbqClmW05tRnS97e7C2r1N
chIRIY2pU3InXSM8B+M5IsNdOFAPAGqCbNemofUWFb7mP/EYzCQ4hlP95CEg4O0cbdXTNz3N1TPo
qk6UG4/IIds4gThNGADszTQyDy+70CoN7UIfNaCL9XFHVil4xMKm5/Q6Z3qV+T2P1puJSDqXi5LU
I8XZQSqGAff9ArfDdTQcRlkpvq1zOAcwLgmWx4d5rtU8kpimOoN2PKdtLJTt6nMNE3S68dbo2KpX
L9d3x7fYJlpmAZKJ5UuGAcib89G1TH9IQoaNSGddQweokku+oYzoEVbuCPJnz1PB2muWNYXx/OYi
UqqaUhFJ3fiYne8dlqFlg82zTeCVNM2KahLlELg1GOm1nnd7NIOn225bygCULwJoaPiU1mK3VclA
Bcp1lZCadJQPGockUb/aNl/dBipJrKZJMNmpVemSmhET/i4JnUd+v6/su8mjxO25qZ+etZfNgYOn
sbusG17+C4Cu2djmovGlo+LztvZXIH5ornRFuxe6219OtNCSzMiVKres+hIORtzS+Z63Y6ik6H3Y
aY7X0xqEC1A54M9MhnrawuY9ETFDtBHEKQ+egrVI4mtd8BqXMsg05gJ/j2dvVTLR/h64CX4XGa9s
YQVfrBa4f+j9jGva8TEU0TUWEnuunHuHudfqgyeInOllDl0UoUO1h1Oc0UDbgZ0PTGReK2aBbG2Q
H5024gpXBuKX9TMg5pcMfIA/d9g0zIVYMZBLbK9GY5ok4qs13T4oXV30ogE5nVOvQP7TVbeNBbU7
qm67feGymX7+Mp8a1P4Cn2K8P+JFaKj0vVmXDsTVtXAwqCM/bd4mRoExi6caUhqzbR3/BN3p6/IO
1bSLqfjUBSKSYd2XMwLeCfM70XdFFk689MfEuoJ4uIGm+1ZzIt+9VgpGsSip0Mhtm82Hci3qua1X
+d+yNk8+4c/OkRNYNbxRf9ivKBX4NQ9tzVmkSdZajxKz2d4OnxPEsuyQ/XFsSRjpOJJ/I6OmJcxU
MAeFcGRlsmeNBmLhoz0OUpT6Zd/qiTttux8d1B//dbtt8cTD6O2tSQOM0mBDWYaL0pWL+TkbJQbb
agYWpM/YBW10ccH+EWcZhV4mCxc1yY9G6JnARSX4ZvqLSVvbgCsydoDV3sdRsYv2HKox6LiADY7L
JsvufXriCRWYhurNNAxCwcxIcWI0ho+2na9g/xI9Q7WXRxt4zLRAZWTbrXe9sipHXIV2KrJnY9iH
mooi+gi7jVRDRjDoFwMeeebmnUoxTqzJo5QsiE2Vtxr6eaVdQsi7r5TouI9P5vM+0vwC1IA/y3b1
FZZIc0yiV0mcF5CN33rYzeBjTdt4N7fd5o1+SYaTLSbiPosZFzN95gBi1wo7YhAYFd4FFyiNIh7R
V6sKQwVVW+UijIkoW//fNgefNXA9BWybyx75MkYvBZfHlC0uQoue4qvrfsxWsiTONNiwdyOWtkpJ
YCHADdb8Cy5BMJM8pvsz/IcK0vxEu9VUQaQha7ej14x8B98uFq56Fx/6wKMDDU9ri93M4/LVRIS7
MmvPFqAdtPp6yp7n2fGXOuMjDKQWfRPoQ47/TT94FS7oVMTHoG40564FYfSqckyJdwCB0FXT2Psk
Gpxg7aHGz/z36EVGz9/et/cBHkNuwX2VWDbnJ1AO/k+OUtmKHlUTHsFClx6I3+TXQH+YCP1cEQeF
3oqqqFr5zFDiVa2SXloMBBNtO2uNgTcTnX9UjTeqaaiqLKw5zERzWyOSMWxKtVChkxImYp4YEQaB
euttSktEc5HsMx5aq/LMhJqI7rbnpxn3Dn8AvFfyowoY/hTQ/+uWPk0YIaSDJbyPDBuUlHa8Ffp9
uzFWgIcPDOz/16dmdZPdu3cSPU+Q5FaaoxRyD/wbN2+oRhUVbtpyV91ITC99D+A+VG1vLccEYHkw
4oGPsUB02f4W0S9dgJBiw2EBamuHLpYKh6fskeabsE4TpQ7u61HUgghZXKM96ElrFzsZhdf/Vj5C
pA3JY6cEO4ptJhpB8uFZcjhdBdeCFr1fA4hiCxpUNiPZbrmkj3kM/F2aRaeGqp9pD78jOftMSJPe
Y8pMha92BmqhOQnLiPUSg0LjwTGwqvHduoGlVw3kDH0QEg1n4B3lDwy8vu+s4RyWGa0v4pYLY5Hl
htoJSS8ktR4/jZEZfiPSO85KbL56bXoqGrNHXdYAjQN36BOkymnl/iJJ44B10KOHBeVW3pmSh0e4
jPRhNGlLyLw5D8ZmVLXPtcXpB+TguGxIMQCCVdlWyJ6YKrk+91jB7dp7ZKl/5NIT3e2D8uNooouv
UHccTBpg3BkiCsCNm5QQ/RxPBuMBa7wHwAR0t5hzPllSO2zkbRp5qAGDW+eEogmungBFAlwNiSxt
SP/PGBgbZfpmvc3Q9KqLrmLmchx2khi/eZxEjpbATd53XJMtd9ypOGp9aidjvMJ8JthS14E82LoM
KStpCZBf2a6ZZl0j4lYXum6E6+LcE0aE76XC/G0BdGfWu5WM0hmyRudC5t/9zKSZp+nq48JRx5yI
hCpkamKgcj3XfT8akszLFyPGp1NBaouh7JOjqZ2+ejkRN9jE0FZjUW7w0inwZUPsVHj/JCfgk6CF
BkdBIGNJu5pcauH62nlH4aq8YhdnlDoflflc17yoC4ZF7hKOdeuHo4ZhCuaEfICuuGpgA6Y9Sy5D
0uycz6jOa2IrATTqThRMmWHj1qhbBhH0xEEquNN6qIjatlQcuKS29dnrtNS7KnPfB3B6VeVFle8E
koqtllfcigMNufHhS3CIoZsrVzOs+MjX6aX/q1p2R/fAuBwGTQnm1/D2eYfoyVmdpNgOo2QjyliB
cP+pdjCMJ3JJlqScFerjzlghAAlHDB/DAQsSU6khAEjxhaJviLvmpzpXOpFmCcJgOr2q5gMnGkJr
ItQPIDyeSZC19iKPiFpatSjAcBD4LFGvi1t+uBTzXIRt4QXAEhMC/YZ/AT+iLMxm/vJjmzhKzEiS
JltrgCNfXvdBmVjLTbmKLnMvIf14peQ2jRUQm6we5gkN2HBWCiAXVnory7atZHxDf/5oOXv6/srQ
ocG+CK0huT9pd6/N7Yi/Q0iN4BdUOyrHwlan4wQXvlZtBeCITyKbYFgeolsKJCTBYCurreekgPmF
6C1KsBEXoqWJ+M2vkR4NUcnAi4QuIOBC6pcZkZJqToxWTgOFIpl+Gjrg+SWxEN4/R0O98XgwK8VR
5HXmxm0SGFZAaaWAtNJuTmGz/th+emK9C7LciDQYDaOZspHlvUQH99ptYHbKiuIsd+6NCkopMqky
9AE3dko8UVtSTM8+FOSkyv3Jtk9OxU58R7zweLr9jGU4QhGGfxol0OEfTOoRhH232dmMHwKt0J/c
p37FVrFevPtpLnVwmAV8RCY8+BXXghKcO4HEpjK+uaczJroF/RbVWw1r2BuqyJQPxtvIG5NjMQ13
dmXL0G3TRE1uzzcXMA+T6/9iY27uKcA+WHF6MXXm7D5FtuFO7ALSnmciUP5ujG2LQBZs3NBhmFl4
Gmc0WmeVAQYR9trMEbDxFokARBzXiW+IVzbQIxQhYNO5zNG05OfYNNY9ziAnAwzAw40XFAynWVgY
oXA1iF620t+KnAdAxr9vtq/A89d6hr0mk/b+7mKAI9lGgkQYa2sYA52l1npGa6uH5YHBHRL/mngf
LeF0sO5yP+VqSCxBmkQ4evJWoXTon3OBQLMh4tpj8ITfxOTkePqlNQPjPDsQ/uEdCuCm3gEtmZy8
YiB6/Jlv+FxRwP26rY4sleP5FzAkddyF0Y+eArNr9sFz9wDZ+dzcxmXceBZr2N8zGk7LITgEfuqt
Q/OZqblJpnEfZZ+w/IceC33hyZFTtgGRHesMkAkrzaf2CMGyqRj5ou/6Z0KQxyCrVzASDOFFe4pI
V6aXcSb5LgZJZb92vxEdslsyZGDCIVdrL8/qIwznS4cvCPOwmTL79Jlev61Dh83FK7ILukAgM+sg
z7a6cwp6Jt+cZagIty//IkgfceEuJwZMhX86LLm/1ouPVJhnCQc+lXstDpxMiFq7IHKG9c1tQFwm
0ocSYTFmLCNfmELnfoF9adrFeAdf/QYvMpLX57mX3aMX0OJcZS7CPxmTiZ2V5FR0aYYJ8GMkBGeE
fsj82p4CbC3qnbp4h1rIo6Rzfq6JTiJaiq9+wDebDz/8QzEl+nuD+YfpsLjRPGlxol6Zv9uGSH2f
fUaujg0mUm1Jh6ilI4VIpO/2s1cJ08+GHpICZeFqzPt8UeTSqMSSw2rOaz6PmDBs+2ZzbxORVqyS
UT2qksTKAYjAe3MGpSx6PLAsbhfpWLMXAx0pHfdKeO5HrAo4gps/hCQouga+c5BAOSAz/+Vq6kMe
hEkhh6StTQ8sDi3DQds9tFlWedM196bYuMW2hEHgAnFHvjdfx95nm3cmhjHexCvUhjXgUbYj8/Qp
ppZSyO7a3DvOstsfVcFELuhDXeEaW2ubpc1e0cHXq4XRbOK+NtC2+pvMwz66gHD2Nch8E1UkVNtE
wMql6ZAh2RN2T2ee6c3TQKlt4uWusYAmxqb4U07QOVFI4jQaTUKrYu03S21JlzH1ZguBX8lZQnHt
vetj2BSObOtoKc2zW9LOnLCouBuP4WEupy06t7uglKg9rxoJjDlXQCpGQKNevUQolO/ZGYS265dx
7nNhupauAPlLK/NabbIum3/cm7lSxGkLYRrsuRk4dfc1+bH+8hUqV7j8Tw9L8kAkb3PgHHbReRyO
b44tSG+hesXMpRQslbOfm6pmrxH5aU6+sEpF6bCxQdKSJlb6565CGa8TSzEVtqL/CB3GuxL7iz6P
wENKYAPP+Byb0zBrvYWxPMHESatv2VRvZfch8w3BX9f3s5g3EgqLgwgiM0KDGE+uYNDLh8CgsVXh
c1bpLow7lgulvaaA48p94GC/HJoZg/JPvQ9aHEzMcKGn/PnGNPV6hwgeyoV6RQm8nsQnEpJHpLPC
Bv0giM5/wjgcwnH2bI1fShqmqS/t6JzSz2nYuz6DEsobqy6y84AYDOnm+5BNQ1+C0wcSSl8F5rZE
YqmrDcqIxuizFlvPQJMIXgsqM2IddgF545tuhZ1dFCLEAPZzPRkhy5P5VArWDRLFxP1GJrKIp2Mt
UHE6SMUe7cp7Ow2w3KYJ3jhjtuFIStAXTVa/W69I14D2oLEjLpF8hpf9a3t2nOtfNlDek6wsxUio
FpbkVK1KyEEu6W+wMfsDefjGl9Fwt9l+f6qCeDqw7Gn7qRhExSlDr7WDf0DgSp7aqxWXna9PUQs6
xQWdvmzqp7XV8IKtech/uvVTq10n9BPQ8AE8o7dyaznRYl8UMmQPDf4iEZ47p/ShBTYOkAgLgA20
Hox41IHJcGOB0VdGUj85s7q0hrWr3wiiGQ+FUXiJGZpChjVNUtE4DQrv1NsmgOA35FZgbOwNZld5
DkZs4P7YHvRgUPQ/o61D6faN2qU3/i5A27RSE6MHjlbsn+K0jCDO1ICcWquTRF0AsY0OwjwFFNI4
8wO298s+LWUihaUIrHltx46X9rLW0CMXhdoXZAnv/JRKL5p9t388pb12MyGa1psw15tHHBNaodNk
vqTfGEPAVEQ8ZLkzZQXtSiY6Fr3qsQVgjNbcPzCDgcybY7u0l30+Ckjlpw9lQg0Df7rFcsK4uNAC
cxJKpnLMXPlazejslgNw1sz0q3O7B+lICDZxsYJ67oC5hmbAJA9uJmsIVLlMWzAB58l82enc1iP5
NikU3B59X1luoxLzPBrsTE4znDiwDnG31eTRKLmWajzSSPgcDmODKXqeqn2RZCEfciNuv0G4uX4c
Is8qBRXvTSXv2eoNeizTKsZNfuZ/cMDcxTqQuMaiMkd7ggPfDYen8ly9JpxBW8BM2QQ4ZNG9nPp8
++X+v0lt88bhNl//PD9yXfdFZ8FjwAM5yuO4mPX81efjo7+hYLYVfAG6g6/6q05ZvtSsdWUHaiVP
BP/ymlqmOXrGxL/n9l8lxU2iLJJD5QugRtvyPUCwKsB0TEZDN0l4kTRDV4i1vmue9HXcpNrt3vNA
bPna957YjiyWpsIAa9e0by3l3veo4Exbyo/TYomKyo5spz0t4SEe0x8ChPKd1MV2oU7gcncnz65e
uz1p69vVCQZcJJaXmmZyS3mejEiGJsWsdJFL0PJXAJn1U6nSqinhVYObN8HkM5wXOmXfPVyoHJbK
/kURjKhzg6m2YFaFEIh2aK4ri0uns2DzKjHsc6WxXUkweDQj3sgrgmkdCb8LZBtqdYBMQcWz/MLc
e0M8waqeXlLYkrQJPlL2PHkI9fhEIdnEyz0aHpK76ZmM9Ob7U0vxTsCqEVCTnlMgqoxamD05LXPu
BpOgWIjC/nFHWYUaokOo2LAGHZ28QHlK4kuXYxK6oa9moXHJ6bipAspqLLY2Piuu79LgSLeb8iSL
qk7J/mB1QhT61KsIuCpiIvBLf1afUoEBdXj8oMdv+kY7UA7Y28Ckjpu/8wctfBWsif3BIJk8mysI
a1xSFhV6uGpP/m4bsBSHaJZOAtSQrCXgnNY+jZtQwk6/jmbh52QM9GLRLuCvdJwXrdnHa8PFpUnM
Y3EmvmwcPAd67+fDiBgpWD3S+i0FGBnEqxHOzL2wknVHGKIB6xAxSsbXbY6UVlCxAeUlf+I+XELs
A7BJkSAD/NMSkTq5tNSdiL46FFPceVpP/2LzJRpyaKRsmA6YE7vJ7oC3nXh/lbeTRgS30J3GLq2g
e9Q0imboXZ0I2Aw78kGbZ1FxTW0DTnxut0+Fh/CK4xsZye0UcMbaxHk+ZqWSDOAGvdzJ6VpupP1z
Ml86HF3X7t/S48MvPovkw4XwPl4ROJfxp8SHxd2+l5oRh7Xc4mI7l2TnZ1WwbIRtN5ngVmjU4LVB
f1WoydfCcCSCWnn3djkng7+v3VTTrIIt8aalP3gHzqUm1cWR2EuTOB3PHWvDTYL4Ns7cV+olHno4
9iVoSmNT5n894hZEwZiGHMVSY4Flf7zqjrypWU1dbz+2Op3Ypc/SPQDAOi3jz5Xve5hoZy92epqs
JXV0WqEMBkRrYZC2h/lnC6fL83uKfYrRJ1AU3VzoD+Ys9YYco4SqkIfn5ErKZLCst9TdVTntqacz
I39fltxNe0nFbIrMaWOk3vtyvwB0ckko8JIa/XdyqD6bRFziEnfEwtwkU4gj5nhwcjKi0wHr3I5Y
e7SFQRZ1l7ny8mvJX5Ec5nnqKpXNYHikZHvDWr7N9IHmFVodRFFNf9VDm52Wlwb3YAJTIqzNy3FD
oeA3FZVPTll/l0uRWKCZIHskVjhlSVtQsUASKB5r4AjvxlzpQaU9Ew88lRcwIFimGClj9IyJQeTn
Yxan0bDlBdeFsox92W8CfT1ECQYgXMIOiMMVYXlBwMVL3BZqpEPVMIJXeNJ7oxrlMM/0M1vYoEgI
9sbXChXQ6ozxcSS2EnXvRkzXFAksEfpNdCLoxok7BBaMT6mAPDw0n/skIVxHfqZnwrA527H6FL2h
9wtRgWR6vSFudt/unDURDboijFpe5P1uwz+RIArL2Aj+4iQ53Zekn7m8D4cx7Z2LUtGdMkO56kcU
+6Yc/YGYOXEEnQEzy8x9g2Mx8Qqrkei75yUw6x1o4IHYwfhRpCtoEagHj/3J9GRC5Efshm3+ugWj
anbC8Gy/RrP4wx/MvYydicVOq3sWifG8IBtr7FcdXYAtNadVzU6SJtRVdhnfPhIxhjqSCtAbzVCU
U/j9KPPQ5p+hnBNpUDzRXyiEDaR2ls9ga4jGeQDHTsKHaPQ1kJQrPQLoTYTatzbjTmWBpIA3SdnD
vaAq1rnfjWCPmak+18eiGeEF73U5ADrvMxL8L6k8vb4TJrqy0QPSnFOWa0LUwoUwVu6virwtonni
noAZuScOIZ21NhQoKAq5f5K7wrJj3lpjJbktqlrtKvT/E/h1gKo8lk7pxK5bkxtTWWgCZtfaTUFf
0pFtFp0pUUPgIGs6gvhz/gX8shM6feSKWAYwdwwY6T/+tIphCaKS+wRafWh1oIhnyEGxzLxg2wwo
T3cmmau70r8BFnr752ZtBRe2SeJd/5N0U/o0DGGz3bwZjOC6lFAjzomLDQr4zQGvhhhe1U6H+lMq
eE7zkM4BPXpA0zXVd/rYWsb2Q0w8lsaeifO1w2O+cskAR9pCoBH3PDtUZgZys3GJcEAtKH84Aair
xQSDVz/dRRbCpUXvW+mz4wNYCDVy8M5geanNQn55OjRY4gX1FEWl3uX/+uojRVLPtWC9Rj5Zl9Qh
1aoiNGeAOZDrngQw5vftpwEaI8dZPxyUVe5B3viGHzlJryuA3kyQpSV07++ftIWFaNSIsUSkd7/4
+YZlyieggBQlMtmHwIiWIF37upelOrt7HgxjnA2xCSH+QKIB8Pa1pCctm1udq8L+KCjF5WgN7Ac2
8GRexSlC5ED4eBLGX6x+B0HoCStn0WP6vcDUyq+ECJC6NPm3t6PKnBR4H7ZAfRVAUMsQwc6/nKby
2DDp11/pNtnjPRyueLgp07k0KEBtrbEZINwH+bmK9HuxPSj1l253hstIvEJ340uUJ74OakqmjWCI
nxgIZmKJeXfYqvBaXlUF+qbzAtTDVzcpgSUAKBiIwEp7/kT40tpjPI3ImwLz5lShrbGnigfmpNGK
HHKUvePARKlyyIeq4YxGsxAZtYeJWdkitpRRuJvyKc5+d+kh0PXm4GoX8vWUMIFZgVlDWKqpLWCd
AxX+xB72vsbFBogZ1Lc9ci4W0O2k+Uv5OWe4jHcAlpRJW2warl6soTm5et84XpJK2hkk3oY1/iZq
RXsED05K15him/srz6iLqvpY6Gt4f7jJPsoAW93Dv2G8+T62nL2JTZyXo+8Qog8rVbeCYJJ1Ga2H
niqJzNqujtiewKTiSzdY1SH2opIIOkTZR41McCHLkxmFv7EfNZLuSmclVgk5REz8WTnSt6XF9i/1
ykoYusvFt1gynnkRJ9+O5JyvzW4GGpQZNdXiTVKZPEBE5EERvn1SwFsRHRwEj1L03Y7g0hF27lVN
m67hUsCQpv5Bs4xQvRJS+5LOjkgExCB6L+k67IDQ8/c9UFVr4UMnJCVZZhhjvEg1zAwK2jt0LALX
fkdAwot8ZvytMxwDQXO25tgfEfXXIpHYhq1WnrHl1wsU0lFE2sJaVs2RnJMfQ2SQXT8LWuURIYzM
87Daxr/FbzBnNAqEhL6iEBh1S68OnLkuG101lOzwoVANOlRtWozPIcsQcAxQ+PEaqaK6nByULNAs
VnT+NTfoFTD70me6Sbwpss2ebf0SxPGgCgQDiNyibyzhUzcuj4fPCpSpN+2z5QftUbUxudx2bz0v
tX3KWby1xJOLE41OySDG7VyBLruaF/hfUzrMf0BQ4XkVDJTqTncZ2nPcmMPKlpUyYujCaCzczmhA
TbrwcC/7P8kpsJv2BBUM4dfa+0QZP7Utb57VugJxhN7FyZNrkPETLrCam9QVNMVDW6R3424IaQPz
pe5CmDvIRDGF1N1jxrftW76EnTNLd22xld5QQJjLjenP4WnVZmKHTG88qszBzE6Cbt45wdQjrq1i
94KTiFsC0U0bTaMrVjtsF3ijFueScMXaLWvGuDocFxixkcs4L+kKOyIy8kqqKdoTtcdX9fodTZmU
n3ac8LdllP2WBi/17rzZMTAPR6aJZ7k4M44TX3/qWRhX5pcn+tBWZnxaSQvFVjdVdBdgNPO8GJ17
DxHnf0FOHh+fvvfaKWfLnRcWgz0zXFS42BX0i23NXlq6NkbyaEOqcBTnFzX7nLNhsFwJ2tW68h5P
D3lhHLyQYm1R7C5Sod8NSW06kaLYelhtj5gZtxYzXanxV6XPs0/I8awiq3v5v14Pqsvo/Z9lW9Tw
i0lkWhTNdBTtukCu0XCFhS7NM3rXWaUIk4pv/SiVZ5c88Ytv9cAGOxuRko6OJNtasejOBu+h2h8c
lzpzIBgumTdF0x2MU9heu7R4GAGDYqArm2Hf2Dh9aDGNWeDuBtY+N+cxAoM5jQA0fSR1UylIkvk/
TBtOv1qICKmytToVE6CaV7FsaDF1lNdSjqlIsa4YQXcdrqVyCEF6Aa3IK4525RPJKndiFr3Kxt67
x+4K6/mr/xOaJpkXy7TZxVbi5+S/P22xGrE852Uu57w/8VpJn6dD5rLvqCK1UlkO0yFwUzZwD1A8
RlVo/BYCp0FzIDlCmDNDwo2auIcIZBJzq/KhkmjguFrdeG4mzAA/hdkrpul3XjrZRT4cpPmhzM9Z
h41dP8afsfSG8diMUmgbCsVdYMPAHpKj+cO8sMl5DAnkzfQF7yAA/9QQ1lTxrpIP9bZvTRskaMro
fRlXUBYX9PoTPJBBu55NzT1YlQONubJOzJyevoEAap65NGO3WCww3oEcXDZWKywDLLDw1d+6+Go1
YIufQK24ik0V1ccumlD4G00kFLgYxQHH7yvfSu3SY+AKJPFpGcQGiLZfVfVct/sewjPwUZSIF3/e
ymeoCRViifFr1zSWlt4LIuCF9X9iY5fiDC8jWi1/68ynsI1mYCylswH9ydMrD8Q73v7ZWssdcJXS
QgbyGbrtlcrn67+bInVEK06ynfnXF5S7ZKsTsxtanJjSr1wWynKbZhBx8TIHat+FJoIULM5KsdIb
AVe+n4TEFWq2R8OUT5hW4pFuTKl7ynL3i+TwuYyKVNPI6T8OlOa62ftrz5ixfI0bqVF6Giklc1mh
18yAV9lc8xF7YX5HBRx15ahexDOaSGUmDDcdsUIgTtaed8BnBRwqBRuEO3auC/lrvWSPPYiszAf9
JSSaMVoBjAi588vB2mh1lKAqHTHwlTcN1+yC/3wtEuzOQ3o7s/9AQoJ3RftSDkOuRKbeJD5v0QVj
aHa24aHDpdKFTOZsBv309xiMhLQ0iAjTOP7xPVgfnnhtbKwbEDOUPdQ+4117EPVcWlyKwOcW/trF
T7AeBMyYVgO1iyDpwpFLIBPVr+VuLgwB4ctGrHfqaWN9kEnC9WeXJWLxm4SJVLoQHsP2qB25P3OH
0sPUZ+SmHT7WmGc0OW2iv57jQ3eL9chKQH8tEdIOFhiHujAjgitw6BvPffzAeoUX96gNuGTolX8n
VN7PB/H/b7UhdKs4QiI4JyVcDtTfFpPqYa2WsM9CagGJQEPX1VX71z8pa2JNt9CpxRPuuO0bOuUS
k2jY5vhfMFkVhZFqchug2+kyBzdfrSfJjR2duqBYvZrjlUomEHaXh1FHaLfnenxRvdoDbqM5m7ez
T8s8TSpPbBp6Pi0sVKxPfKVlRlnldXqa4vGrnZ2q+8aDPAGZOedfy3J6St99zsoMO7UQQBLdwZbZ
GkkylWlu5E9umva4NB/ggY1vu0NlDulIDpcVxgZld0WKBzVCXxGh5OVggGRdbyhbPDJARqn6OUXj
t4GpMr5J9kS+TFv6XTRan+1ZjS+BDJoD9SnJ3tORDLURaCUot/y5/u9A+yklsh+GAGm2nIJP8vt1
N4ppeh2Vc/pxCn78azhyVke/PT8sNYr5LNudagKkLIGNTeKK5bjOYmUF+NCUNMNmJJcI5LuIYJec
YB7pbWpBvBF4kYYTHxMAWVvN2tPf/qtniBp1laHvD/wfd9K6550DeOdjf2jn6eRQ+FhPmv1zroCF
APIPIzwfjc/NW1+1PPxk+ZdzywNUgJhRRcd+pJfBj/d5vBbWK8//xu1pKnflRuGV8SZRlg+b8F7I
/m6salTld6emG/OA5vak7KTYF7x3qt9G07x82GH9QVrzj7PYekXO6a2CYK+7YdssSoVPrBrr4auX
k5NLo/wo5BmRNfcoJSb3ZX5Im9L2qvRkh2TCLvW9PnMXurfdQCllCZ/K440Y2zvUIQxKoW279ObP
ya29NMqQJWReg4bVq4aAXoj13TilDjy3rCZciQZDP/4SIYZFAAEwCc5r4lXv1Bn5Sw1Q5JxS2TpL
Eu21BYml4iQgHYXSjpQr9i5SuDLwbjpF1seP3kvkVyqpbDcF00jLaIyMu6tg61jGLEIj3+lwIDtl
RneQs4nun0ucPQbqF2nuX8TxG+nNvY1UuHxPGo8imPUqS/KlF+HTl3KprFVPCsdEHwE8BaRgMiXy
wsEhV7YduT+YNRwh4x9CTHpM8J7BoB1NIntuPFmvw/tf6UkPTxtQab7gHNTbAUet7Z2uM5D6PRQ5
Oefh/JNkgUtZKFB2TJsj93MLwd3zOROF6ZbsCe9y8/z5LPQuL69uNYO6weB4xcsAgXENp0sH95NM
b7XIw9YUntyFo9xrS+Hjklt3f1ZVEzdtP6TsdcdsfFaRta/QhO2sXxJS+4i2RSwV1fZLNDPU5UhO
HTLZLgoDdoQfoCgu/egPpAVF91hqZH0P9qqnzBCN89+DybhIx38xRFSd4vrQR+5c3dBKlKjmcDac
0YIzZcatun7HHBM4NRKC7Tp27s+8dOJUkzLOuez6WsnbhHniIV7v7np5AHDfIcEZK9uOTXiJXVcd
GRyR/IZg0lUZrg3OQklcMZWU5LOWl15ajecKAC22AktOhmQ3hfDVbSJCgzSvPHY5b6hqsMoDDZNV
DM2HbgczQ1v29l1MvpPWA22vJfij7LYUfzInfZKJ3OnGNjyPgKZfCWjhEblWp7nZve8T5xnH2xIA
r58hbhygwIp38zO/rHQFxlQ6bgyFcsgZB3mNnwMsUopzAUYZMk1DmkLh3vekfdFF681KnkD5PNP9
KD+f8m8Zjci+fLPI/y3z7SssKRKy9jj9nsXXT/1KOgLR2P8PRN9jW2vwxlyyGHCe4XPER39C6A0e
HIFcO2FU1we+/C3wAiU5O6YraPryoKiBSvNHyFuoWTJ9asN1e/6IA+lUi1ad9aTvaAUTLy16rQVx
KyEQGHxvokVlQyG0AiZBLBjwTnuyHjGJ4MdWyrAO94UTeA0L0icKyxLLWcD8RHmBMpOYjonGnavv
FUZJTcYXLwqlEf5Q7zlJI9TXk2IJgtWBaJYvHR8Bu2jUX2OFaYXf6DQIuE7u9bDTAQUjaACHzngB
IFhNLlCfyEnvqut3XHuHhf0iJXhFs0B2/RU1Mx7rmF8yYce6XqLnZAkOml9tDW/cHiEnzA5XgeoG
LJc7g0+tGUoiJVc24JiPs1Nii2oifEzJBwMYAJgjSCzQrsbWQk9gS/saA0exTKcXHNtpRuAbcraV
N15iuIOsYzoDCehJPkFBTrvtC71dBbshSao7Qm7Y3+nSBHAgA0MKvp20dOnk9n5fNKuDsAdwCrxb
WGiv+lUU3Q5hgaQJxunjNVIeX6XyxyUapvmPCXH4MuZBvYpR90ss86BSpPuFAXl2xQLaqrETEG08
KZ7alt5UsAAXOUiaUkQiNkISSCYs1OgW0Xglkni8EX1r47tRKW9ksGQODqU7IXxpoUTfXn37FNn7
73JQz42RDhmhQ8c9+KNe3wW86z5ENQCsCrf02ejIixE5/JgAcEDIx9aX3vsGQCrRBXhrtuKfo1L4
bXXR2umjCPK5X4eT8+PGNQfQcE/7gVqR06L0dqJfOraQTf9448xzIf2E9sEoc73wyOCHkFHQSaTN
PHObhW8w7WfGaCYI1nD+//pYEGbAY/0c8wJrvTMb9JwlukxJVfEyDwbEoI4+CK1yOjlftX0B9Czs
0hbKqkE392rx8DvjNnqcFsyrxh9OL9M9vYzAdv+DE2hE0cMSDPSEUxmHo+wHsn5XrxSIVH3ox0JQ
+9BL7uI1gjJ26HtEW+lm959co5l+mI3xf68/TbAolSBZ53ew77olGfTXCjn5lZ50EB1RnwiruK/b
+5IOzo8fHzk1nqpkRfaIZyHnO+WkGunE/Lm/f7/gl1kouSwgBzi23hUzhjNpFb/isN8XzuN8wDxL
K5RQC/MQq9gd+eMOLd1QUymWQofME6TLvVVUMxkq9//RuJYebBUKHHiPoFT2XP1eznFVNMwqIJld
RCPYoAeAnMoP/AcSHsw5Db09K4BE8o8GMI5P5aV/g7HVqt9/q7A+BfBqFPFIUpCJd9vlUWGxV+i5
y9jmlQtMqJDfcIOxcz945C0IuUnKusB4PUI9Z+H3gG0zYlLErVPyZtp4LcNzLw+7bSMixkgRN3Ss
XVVkGLq/IuG/B05GyFTOYAx3Yv/SWcGRRGrRNEkbvCGSu+DW9yTDALANm8aA/OSC271qJvVNCfMO
it8sotUanFpNTKkkI2c6Kw6jovtP6WjUoHRV+EKDYf+Fo6otuwFVNZgplWkuSizWhZ5+fQ/wSf2S
zBTW/ZQA2MkXFCnGA69j3H6NI216bG11wZbW+XGuA5M+UCqEFH/OjB1xYib/Ejk26BsyLtDT72qa
terUF8pbz2a8kUIpnNEsuIBMUCW+QADoC2M/DRYwbI2iw20HXfwtQP5MC1by21deF3Gd3IASqymx
TvicCcAyGGVuExRc4MfTUSiXORxTlgJp82ep6lhMsi0WmfX8qGMBpS/DX/Dp7sDKbHH9sT+U6Bm/
1gQJhZDpix4NcuZxSmnLlh6YvX9vIbv6ee84IUTWTCBYF3G2Um/3ekGhD0rxcjyeBqR0K+fM6At2
q091JAztEKD8BWaBK3iq9Rgb4XvXHDUl/bGGiz1T9Lv6HkFpsGt7aaoOXmyZr8/P7mK+Pf1Zjnae
y49TevHGy0Vi7LNjngKKGtDLEn1pXq2h8mLZhMwibH0Ibj4w3ZARMgqKHjiULCEwyhLdp82f0FOO
LTcL1UwZcCetVAXlCNIHivBajHT9d1EhQYYU5DL1GgihvljHFO89eqPfIvdVsngaJkMxCP/thDOG
cp9pBamwILtfUKSEdWNMU+zgqd2k7vECov+epy5zSG5uFOGFagoiVIAyFYXxVIys19leewgZVjAT
oxa8IsW7cCGrUpaortS9fLJuhErTQdCg696+hL5xnSDsDUlOwK5JMZJEhA5alfaMGOX4TwqQihQS
8eaYMzvsOh1GpjJSDElpb54qd+8UkmfOEKzArTeKXeeKcpC41D5yfpW4fg+0BZjYHyaJHA7nilfy
cPr4Eq1jqA4vW+vMZj/tqwtHzarzX2ecZ/Q1WFE7HmwcfeBDuB/qGFrRsSty4O4aNZHZysE8T+Mh
me1zUAANC65zkLe1+o4fmT759gUJ3xqze/xDRPwI++dUv9t4ZHiYmqCnNs+YvMYROVwfQncWVZT7
Yl1u72wKpShmrx5WHKehHoASU7/6vXSm/1oLjK+2IvNJxSKy3IZO5wW3Cwa84OH8CtCsItd87/lT
sytrinPISGxJenEYNUwyS5Z6z525hQ77GP8AL6wLfruOZJO2yQ1zdwX0wOeKxUNsXh7ViWNSodkM
K1Y+jRrBo4hfOwxsirxK1UKLJHA3nX8CdeBT23t5o0y9dt18A8ukWWMqhD4YiSMsKnreW53tLQIA
5fFW7+x4KJWMRKNAlhKuOfCR2CDqxDN0fVgpNckNNLwhL7ImOCbld3qszzwQTtp3QlISOoCmVfdQ
tcLCXYOv3+Hi50N5gpyPGAfd5L3z/PPnviCBDN0yDOCEF9Qw+Jyk2EQdod+YJDh+5leDyeTjopax
0g/6mvFN9NY/T2pGsxO3cZLVmtT87A1LD3YJGlS26Lup0VpGq+lcAK/ZPR8D2hd4kB7KrK/cTu+X
Xtt0s4gJlHVVm4czELJquwVwHk3/qxgoIK/KwtEKMK2VboeeDkYwDwxmONL9OjDJksuPEu79Sv38
yH9QRrqgXtv5Cv7LoUinZBU9EpFdYWJQJAw7oegk3SiyFVh4ZjPPQ0ALokoOnVv5ZbBdYF3LPgQu
J3zuPDiYVElnLPKJcnL6fB2bYlsnwZ0/9BJ4nYheTRmGdfnVEEA4KbZ8LoKSCn1u11Nh9Vykg2mr
1llESY9fXlZTWAF2sg09g8yQM5RApNXHa9LXwDWjLG21vOdZV7sPEX0eHDqj92XAM43wfZZDNEsV
kA2N/rlkajlNG82C9wwiguTVMrU/wUNB47M4xjRgQZObOhZKVp5CED2EAtiIY92lW0m+TFo1OUb7
2w2oo6egT3joY9lMQPB219VAADOd7s8rdg+hLWkPbOkGl60PL7F3LO14EeBv7e/keOe2BBQ9SZrE
VXQKyu03hH2Ca6stKkeINxFj3ERQJOBHwdDiNKq61P8xhhWJbALXGk9vmjxxqu02EAidmfXRHYcU
qsD/lG4KloXYndyvZUY8Q9x90H6ERhvvmADsOtbEwkXCz8ayikVp8/teAQU39k2Qh3/wMMR9NhFV
gK/WZooikLLL8OUWi7c3GXaRBclFL3HdIcN1Futb6r83YRAhy1+tV9VdMa6C/STtwlg+zW823DHZ
JzyTJMbCD961bLonRdQMBNAjwN90Ow8V2JM1gG0Iwygyiuc/kZoiXZw2EWOhKKfClwFHA/c17rR9
2GYb9ShBcTjmuhSlf+FN/9dJtEaMoxazC9H4KVGIinq6cAFHhizmeZaGLXWII1Da++MmoOHpcIXP
7lrjIZSUYKoEY/UiS/0ERQJndFwYrMac4LYEzoTzXu5FfT/218QCLQXegvzAR2JszOXHYkZvTBTi
YDxCviglhVFoeYOS+AoUPwgHVMCjxeCtd+r11DBuWbwnZUwDcJu9U3C8Pjhr7IXLZIIBUcEiapGl
5j8zC5NumPKBJ7+q3et5qAL4DvGczcGJ6Y6dN0PTWbAZY8na3Nf/WPJegWEV8wIASdP2lrcrNhzm
Y35AKbZ7uIl4gkInIlE+NJ+5CItn4V6TU03f5AdFkO0nfb0/uR5/BP5MuH4MppD4nuQM6r+xubxY
YdNeFxfk7JEvpjyxsRYOBDvUfM8R9SLejKcW81pzbMloagTsLABIQdTlgS9gLckj33cN48PNj+PA
libTRGPHmFXDweUDqpjuG99rYVyKuOhuaHCMXf9uJGG8vpHjDtc5UbpyhSDiZThpFIC6c/br3YGc
xzlCOpZU4VqBedazu9nQnmozK5uyEs0oAqlRsGVHJiYux8+UgKHOM8MjWdK3z3BUH7uGzzY/yYb0
l2PbkWZ0WPFcJc1rjOfzYH04fOJvzRqa29XUfj8YxzrfLfB3gaK4wucoWMUHR7pGwpuDPfj2O4/o
ugsqLqqIdUCgyzTm5ppwX+bsqCW2iQvQTGPeRsI/BRmVTklfQaJY1DLuGeOmQajBKG3yz8TTd9+E
hVV921qnWunk9cfgQszqwzdFY0Pb+5cs8myt4U/X14pRZls8dB/Ovl1++D6gT/ZlUAFwPsIeN15y
PoieVRn7WmUZotwSCyq6rMj8jW8+PHG1Gp17QemswkY4LmLpcWDrpUl9yrvRv/bRMEMRnQyJUzUu
zzXVw+FgQOgtjE+/K3A2pduTTV5vt6nGB9AcU7/JBjdOYVniw/vIDX9R8LU20qs/18SRYANeaB6F
gGocFgU0cLZb/qtqxNsEmGmg+sOH0xKCuC/axc0Th1Hs02g8l1oXAjMdFWWraDSx7qMyRpWhr9Ze
achAwZTxkluAl54tSHRS7zWohy4JIrEKV9/ph1MlRJYZJKGNZf3W1qy4jBaohdOuN/73VjPNEEqi
fHuD/3heFzPd+vuWQebnsRS6l6zOv0qonkYCWCgcWi1lucc0Uj522uZ4nkEr/iGD2QwUcFK+Wmmh
7oa77FTYWao8Cf+xlM4Qer9fhmW47gHFPE4axVR4SGGqmifThx/9zjW1nRvPj8Nm25lN1QmC0TOr
fsrlUyuxJ7nDYr2vpdy+tJGg9GpGohEcE3XYHiexht7YmTKSGfnHosYjd7OxeVjX6lNNneccLmi/
QKGRuXLMloxqqsRAKiwI+eNZOiDQHsiEQs1H8wIBPxskGbNDdswVQCZSMBgrS8Rg3CmKl3BBsr6W
Wq/tVfsEe/Ue4lYPu869IjGAUVWe5zI/dgnPAwZSVonu++eVIV6Vs971SFFPMWk66m4kaJe5lVQS
0qu7heeRO0UUEyK9Gm9aTv2fUm3ZhB/DPhhlVuGn7X7pg/qQm8d+dd4mcFhWoHPxeHvgQDhcTbmw
T1Jm/LFtAgUM8GURCpbYk2hj9buMNhj9Sb5gxBpr0uR4W86I6DJMFCcBrVWG2B4K9FHcmz1Wvbqu
sVj6apWx1NQVIX8olIobG8FXN67kUD6tk9GAOEB/JuGH4m0pCLj7X5eL28qcv0aOJBykCGwCYxzf
SssTXi4Bna+ETftwGf0gA6NderYMkkulc/YUJugk1MCvBlAwciBlDKQeDSdBGDNcOwU0WOra0PjN
125g4MGfU6/RncqusYoWG8L/X4l9KD4qeKWXlhFhDpAU1J28wcDDUSw04wg0o0cITXCWFBjR1xeR
G4qBmMynEQ+rtCn9QetNoMuNWflDdXzT63Bhj7g1SgDlGsUtmD64sr9h5wOL/+Zwv7AHlVQOW6Uk
vU0qn8c3mpMGb1OrPlKNrTT67kF/r/NNJVyH8sAn2fOiRg2s5q4Xya4YjHUBtNyK+1W7JMMcSKJS
KL3T+PTEyGL6Xd2dhQwdpWse4jOQ/E82ntLbf67GAdnPna3xIh91dVaYo8Rc083fs31hxlbJE7B0
Sc/xSk8qiL70NIkVHnjKJAsMcfilCE3llJ94YJ/mPQBao4pAZkxCqfs6T3CwOXsPVTCMHsHcYXMY
pnRrEcuHyrUVsOu1dCG91QowmaHgDD7qXuQLTTi8Ti38iZYioC0ZKYXOfWxqPqLaDjg85gVpsg2Z
4jy/+BsXDLsurb0Ymf/CvSiyuYrrchAwI31Y7+85l9JJHMSTO/SU1E2Pkl01Jiop3cPHZhHzGG/P
xlPJhJoJN5xa5QJ8nisvGnPNbiiJMxqB3U3WC5ospOk7Ig8jBvhcu2V6GgVDOPtqvV5LGDvbhLru
SAeQ7Npmkvs12/jt8aByhHcANVBLMNg3iB/vav5q1oX/x0ozeZMXvWL9W0E2aKFRh6xy3hd4oZjO
6B0tp7Kt/xgoh99cvl9jqdzepv9O3cKxVg9pDm+sW1SIf6rq8dpHLnT+4q3LwPaGVdiuuJyhK7Uw
WDr0yp/GLfEuE41Cyd+jGodzJ9/qFaN1d7PS6dnZMH4U4O8YsRnBTPquK4Rf0kN53iCICoK4FQaX
UxBTuIBk6IoMunytDSC1yhV9N+VFwrmyoklI/OMmZ+Vec9fCC35qQGCM6tWe2PaozZeZ6s66NL83
08WYkn8lFko0jhomePgp/hsy2X1/5RoUDM9TWIC1B8TyNqGNrJzI7yM89MzYmKwi532d8dI5gNFP
wNFR980A5mZ6gj57XO3EDlxDs+Tk9VsHikTUpfMrzlguTtf3e8FjdY9SoXb+dcE+VZ0Q/2je4B+o
iC4TDiVYTuFlROp5AytDBBa9j5nlMAKFkIMqWkoE2R9kDlRTTmisMQBxhguO27Pa830XgHO4BeUX
ggHOvBzBL4d2yC+l99hpfQq2O+AS1Y93QWqiFfP1DVyHi9Df4kNawdFK/+BCUqYqgcF67p/AChkS
IIHOx9+GJJ8O9PgKU8PmbF39JmEZCeTkTZx+qsva26SpASj+cbXumyl85TLTewkcoqaA6IIxRzdB
+b5rCJlekSheIENKmqRQYW+ty/Tk71zUuVw0mP0YMUrOfiK3nSC3bzVHrL5cmZ/l/eCLLuGUHAxo
lDY/3uETF8KLnNZ4q+kD3U/bAoNWJUfYZenf6jx4zkAjuIO0z4kSO5u1VUdHEur9WdTjZnTRqL5i
s30OpcB9V1IVBDa/L7dK+JZU8Ay/53TyzCgE5Ttyn2dtWrSayUlB7iSYPjB2YK+yiViGFadsNXOB
iAZWlEwdI/hh89h11ajYGceHBOn7VXyvthMUBy5ytUKJF5+srs4lkSv17gD0aTby58v/EdnObG1C
u5HJAVsssAjEGi3k1SuDOYZ2WM282+FRPQ462oEv/Wg61tkxAV3J/g1nMk0LRpaXpERDMTlvXRgt
O8aKL53DbG56W1RpqiiRkBHhxtiTA+b9hYYj44Ik8CJv2L3uIsWLnRHxfeH9WPSJC8i6LehlG8SB
3Abs0qXGZfJg+rMNJGJRYa/0NJBC3z6xpO7GhWByXFNrXQBX3hIsT0Oq8nxMeJINW0HIG0JRRtqV
WnPBvoLkaT92O1zWbx937sDiY7qKs166nJqk3oSWxgfmwZe8thuBhKN9GjiP9GLC4OS18/e66oiv
vtIEFouok3J6GoBS3hKk5qd4OuXKILdUf6nL/euyd05BYpMUaN9yjJ/zxg214JvIMPZh0/XdM7I+
+gLklTZ70rOkpdPMpp/ZfBkUETkcJllG3HcNEB+mVA1Q40UvL0ThkTiO+0fApcOx2hUCbdPQCCKf
A8tw0N9zqqs0AnIwNR596ebQ2axQ65bWptmX2zcgdqf7d1DvR7RXkjfzq49plOBv7zyx6EYLhLWd
qlxbqKh37QLOr87JJgnIHmWRChWGyutOSyGWtzpCczFFbwe/UIWDbUlKlJ8js5067CyIDnrz3ENS
8w9bYD8a1ahJvsLGHsymFRwZryXhDXoJBQdj+C6iLDI02TcXPOmOICf+X9goCXO7C3KZz+0gYYgO
L0OF9ItiG+Brl78zgwp7avbuzKWzbyGsP/rRkNv7Y2lwXF8kljD/KuIc2weA5bQ5EysonnerI4er
ZGb5Vv5Tw3vS30Lec2zRCfM95+FIYusI4ywmGFUBlbcnMl7UHERcYTjNR3ZWIGhsW9Kb8vy3gvnI
Ybnc8qC8QFyl+Mi6royvjY26kEbZi3PBs7nq5W+vwYVTHF5JiC+IN6NFBGUaqUrUtBlrkknxAG1o
7mzuUJxYWVnunipPCa6nOGKJF1CtK7eN2NFeAfPAeHYKJFDb4VWWNM/N8ASaw6jO+tAWFM5gjEs/
76XUTMh+JUTd8VY+DOI6S6k3POL507uLLp2O1jBU295/xc911yWDsH3TWNIPouwOQZTLxh+I6KF6
8R2yhj8LI7N6bZhxvOMnqOFz+hDNi+npIiRWFizvCYtkwCeMB1Fq7x5ypLW4BaJ7Mt8LGH2kMRF0
NTPrJSb9Nb6Z8nKX59j6iMScYef2wBEAPt/XgkMdUiuCL2knh4EeEf0v2kWgOo/yEExBZaup0aPn
mW6lT8182m0BBWTwjJZv2iAgl12NXrCG5mcRgkVRSLLZeC9zIjxFhOCQOY2DuKsfkPwA3oo49u/t
QwAhFXz4fWr7DDjoCK/987c3Y4eeNdr6wjD561PUcpfXgCPU5rTsomRya7Cmi0lThBZy2RA1laXA
Hl1Ncr8DoTGauZuKa7/W3JIfg8/uI7uL1F6ECA3xQ2+F7V4pjIfrQ4OkWQwxhTGP+v4ghnLi57Ls
6i4o0HMGqqKRd0iDOp+8ypiGVIO7sNfByDqK4YYIGkimRoDDTCNW4afEi6G0llFlIj61MtOgIOT8
MJsJ7/tDJ9DKf0tpx9q3+8PW5QfuGy4Z/0lmlxD43+Dp2KfcAcZApb49I/tNWsmKFPf/8o5i69sO
IUTwGTLXdOfCxS3skXjEwC1I2j5lv0eQmBaFEBreoLERCqX22YEvwZ4B1tbzNcdMif7VBhqYhBvS
aFEphsQB7MAhPuxGNLI4rQiY2LCGc1DWxeWMUIe1EBur8KTXk7pdy48s4Javq/e/6FSCezLXA0rF
HD0huIQWteRhEXENukJcsmb5E0iRl1C1Bgg4z6CGg8xLKECusVhA3sl+j3tOIofYe/4KGxrKV0e9
R5OYjt2K5rcuqBGSWLLLU96zXU3AoZhttdgF5yTStVzT57xio2oQ46HooAPbvlq03Velx25L9ccl
pzF2v8Nxn8yBo2ijiJtIMJdITXlB+ysBo+v6TP2sjg7aRoXaAlyjvtsUwycvR7GWGlSDf3nMSaDR
P0npOmH8H1cwjhIKIs4z+pcXOX+RQO/L7KVPAz2Rkq1kB/NB089PDxkSmkma7F+2XfwUmrigQzYC
wdCekTWtnnmQg9RdjW+oo3UlY9eBBbOdUA+0dHqbXCsytZkzPO16GIDuuFW8DTHye7Gn47DBU8Z4
70GQ2Kw6Rm+o7vJgz57Hd2Ok6Pp/xeeDc0cE02C16M2R74rayqoBpjMxR7H6r3by4PqLsgt4rBx6
FQeaP1BrbwRLSc4MDWReFuHqphSG+tJmhpCXZ7A2HnV+LkxbISiquVxc6RtOPNTkXf7/4JL3VjFn
xBup+ExZi+j2vE615ZP86sn/z3q5M/whjpcp4veelbWhGAZo3S6VztIAyZ57iHlNCYFzT1bvYs4i
GAEeaUukpPvFxDkwp23FDspuS0alGHgkd8x6OBbzjDUiVO69e8iDmnlnh7QQ+beHafVvHESjcdY8
gx7KDNwN86yI665qOyMb/aWMKMeiCEmDTy8ZFUMgkgORQVnwkfuKzPwqjC5Te6oV2jfaWZ2OjyWY
oDmSKhhuq42q1PWu091AF5LdGfmNRUJ7X53X2dKBrl2aEjMuxt6q5PzIv4I4mFb/IxP2EzT/Xu0O
qzhNv2Vot5YciTg3VzUOeorRUfIYQALSItQrlBJ+J51OFaFL+QcLtz4Qr27LcVAD3lH1sMgeE9iZ
JW+Cynoz+6X0XzXVgTRtB8xTQc6JHg1HdPCvFGpT+KPrw58tBkYSeGp+4RCOQQrxYkhC2bU7NaLu
uYzUY6bu3EC12/Wqvipen+BaO8Q4S0rf3+W1fdMvmiaBuw9nERqEY5VLzbxmqecy/zeUk27wLXL6
jxxG6EmHo50iaurP3RnfKQ+mt+9+DsllxuK9PJdqBUjpRthbtsKuay4Y5ZYctB43s0ma5GPRCPjQ
1rp2ThrczOiPAD53M9Spl6PDN/s7GW4pAtdRJVn/Ej2CvbjhSQPGd1wMY8e0xD8yhsrstU9qAk45
5lXqGkcxTSG4IYAhYqr+D9oIh+yjzFzl/EenGrmYvZJpzK/NfJ6LlvViwUiGR/6olJC11VFQXhYT
9C5+X+VD6GZdWcA+pwmcckHScs6igvOtF0RvXyKjm9lsGim5WXq3sE+/JryXLXoEjrH7N7E3Mnnm
a6Dfdzr/OqsuvcZWcP4Rx8YuBYN+fTTfurhsjZr+eU6GtbP2L/9VPpwAvxDd0HMLRUDF53bQfp+U
dEvp1XMXsPMjRczTFFkenkEAyjnJqcHgGFpl3L+RTTDTiB93iYIHbVM48R9LzrUHZ7ohojPHD1Rn
HsXXInPb1L7W7xO8aF6cOcMUDOv5CyVwUx8GE9jl72VY35IbUo5bZGpeIHPOmismisOclvrWGXfL
Jc9sUQdzNKHF+joHtQ6HkFGe1UE0i8kRglrWsyLDICi1RCS9sYlMhXXosa97eW6sKSValoTc9j3a
BwJT4ouJTnB+oj68STYAzIstrmJGAQYGtw0svjhdcCE9HILWkef0cL9syYIJrB/Hq3cBhumC6Yi1
YQPFhwnQbv6isfftAqpM0oWZyv64ohIFAHr02gMYdBlbnQwNqDIH2ZRZ8CUBI+kLgStvCz7TtEcj
uPRiQVnIAZVm+kV+KihAkeFpw2wQcIa18bgMvLXx5WEWufYJpLndm0ylB77//pG3RcXzqfpge9SX
0NqpYbB5TcVEnatxTwR7WLWlmWzwMTJuUsD6wQnwuRxcLWMIsCZdjJsy1WN2GX9E14pxbp106SdL
yu02HG4dbIFEaceY+erNBBNdMqeE8UbkNg5uLZ0OtpSQkf+8aXyyUIGw9FKuW+t4ynK+IFe7nqpO
P8ujBPwI5SEKvJ+dWn+tfbOqdOhTvwNFl/y/In5n6K7RM/vU2/edrTng73PEWjKViTSGxgN9H9Di
C+9JgmCQ3GjFmD+0lTNwv+TbGSvxWnSSHgkXt41kiuYCZ6VhafdHK7bkPVHOQfVwLd0ihRaHjiSv
75IjGFhNlMD6i73eam0LR71+W9wIzCiAWMVUJYgidMCpYa3zbmMQmew7BdWVAlg5RlmtiyauYelj
XNerGSqYwdsujKCDhsF/ed0gG4SKtCYYIiIq+IetiCWocNkig8XWB7vTivUICjbbmsIJ/Azs+nYJ
TdMtTvlNS0GkHFK/+V89chtKyQ6FI2nNurs5bg8myEVD4KHlwzhWWnIyC1vVegODlSmn8tvfChWt
Z259U4jTL1IT3JxPumZIhkcT7BZBDeEv8XFuoS9wLDIOJPFwNcRKzYZ1MLJMRf/Gt8h2y4TpvRGO
FQ02MZRt8Ys+5Hfxb0xuBxu6s6M6Y5Ztuc9qQviDRwTdYUABCym8Z1LQTwAtfFG0FHAf4uSWm+YU
aND+CCIB5BLVrnFuStnlaafLwc1jRh6v9PFwS3gCHTMElpdqc+WdhqkXCYT3CF4jADiXWXlEzcDo
eQoajHbR6k219LStduM/GSG8aaEFO5LyBghXNV6rupS1ujb0wcuwzgG54dyF7Jn2gj7XhAKnAJQR
VnxdTS1LQ0XfsZr42+UiftqC/1nsdyYaeqSbQVtjFLyasm+wVFMd21N2akWGfjb8z/OC/iSDV8Ic
h22Qfyn3pjSTEGQdLWBHyO3cbNhO+Pr61Y7QvtAqqehojz/LP7M6OAHizqsOEooKrbLtk15GzZeV
+6DXTej29mhQkhK3dII+2MeurI3F+FG47tScKyTpqNsuBLmACbnoMFo6k4Hlou8gBlLrElnhOJ31
yLwKLJMCDxLIAeaSoj7DDe0bdMW1gGS61iByhE/RHm7qpNTKObBrsxS2AiHev1TaWS7KusnK3jyC
Toj5m2wshmFw7xkIB/QVVIPYXqqeUCobxhCtl7g/FTKsA1d1nnJNRGZphjHUC4zRqcR97LQb0q7w
sUi5lWSCfgm06bZ9gdLljwReQWnH3y8Y82VNpGuCNYrQJARt7B3kbNat8xUFl7p31aeNgT8A1tKC
buambPYlo88tns6aZMICNCdJbnUCtjzyX5Otc58JievBrmOx4iTL84uJ16oxGogmBsF7c1Zz/SGd
jiYYubul4oxUWmpW22IecwXWS3kr6OPkFbve6JLc6pQwUweDBO2DtSkanHy02YvPKvQ7+NWd080l
l2b9T5MNmk/Ru5QwzYb+nhMJXxG92OydCOFjy5xCTYWOQnyGHYMyZylLok2JPOGeOFAcHhrKCp9T
KzbbaQVbC0/LGojLOGJw2Dluu850lmqLVeYAdow6vsmnUTl9l8reQ0MaYxdE/J7Sf1L+f/ywvP6F
dzL4dnTRXx9H4dWxKRF1rH2KhuQ+t3a95Dsiee6c9nZJ8+7eCNefHq3hWsMvuFHlucHdxPhvcDZX
naKVpsYII/Rv+BYGo7LiyYsPZw1+b6Xmsdl6A6aR0YOsQzx9dcLAQmktJRCDY1sMjRnnb7SwizWk
6VeQuTZEha9J1R2ucBB6VjdqdZkqKrCQh9RwiSRxHukt9gGkQQa/uJm1+mnYrAlSi4p75Fo4Ya84
UTgPWhqc7gQycvEQUq1wGRWSCD/W2m126oYB1u4t7FwGqOmm/idwgby1+6W08NA2+WVUnzzLLYu9
LNNi6qTAx2rCdotw53vnZNHHnVHGyM7of3SY4UyS74Jz+5zvcKik1VmMGPM14nIE1NtmMutn+xN5
4UiZffStuZyml6fXdghgjrIeIOcH1ZHJKrLieyvKyUg0eNqC7+LD56uvvT5eGC/xHL5ZGUO1X6eg
j84n+CbOjKRdV23Q8C5MH4bTFBe/nKAszkUUoo212Prm7tmc9S3Uwl5Z/aSjNbpRDx7MIiVHVm/B
Z4feQeKYj2gw3Q/VQXXKC47K3CePSKFgAHqySFNsgD+YxDHrMnjaJCy20XZFPvj0dN0xDTZ2RDCZ
DA4/sLiuW/Rd1GXSp8aIm6djQ1ENKfdfbGAjxLMT6IHCbQ9fKGIHP447MaLHjgE3pHFtu5EmIo+S
ZLUlvc+IDvTxJjTdj3r4meYHvmVfUTbwmB6D1WoaM7frvBwVnKNXqX6QUWbW8gZNbeRDq9O0Qu1y
y8bY/SnRTpR9fTib+C8XbrihzzKOCV22m1rZvvkWKw5+dsGbb+ta2BXZNhiyljIC3rubI2fvOGT6
GmobBXfLZdjyKMUPkbEdDO1pQNOI4D1VeW+PNOiCPm19GcXnBwOi3GhUWZs2nBCCBoXSb1Ri7dm6
Wx6NAoqRsahtHQ/j7rcXXemWh3ZIOT24/dC1Ins4caOe6d7ElWpIY2IxoCpWJbCivNGUjpXMP6ex
vavYAbAlRxzXDygWwQCm4/vLzx+4H5sAsnlJDWxPJ2p6rivod6BQSLATsNhNaj2Ped1DO5eSj4uT
WKk/RAg/9A/PVhMOvYivOZN+AzQPsumCiRnV1jP7dnQtmtBGqO1cY8EZyoqNymx8pT6Wc53GmUeQ
AA/tAB1Vvu5zDFseIx+CDCTGw6OU8lFJdSKzWleNVBLuhPXmVitipLiWqjQ9LQnArn8r0me3WhMr
rFmIY71+zyFvCtpeuHB/XatcO+NXtff0HSbQ2WMdysE2uTLoh+HzSn+7J7hMvjFY89wS4AsIQgBF
FQYgfjiYSPHrAssAKN1c8/kDtyAoaD69hpflGhuYml/lwe0m4iHHJtE8V+cs3edGGhRkbMngM1I7
9F8MIfrJkh7g5AHnk6xAlj+Shb0Ghpd53K5mKJ5OCs1qciv4dxaMnx+qySp4/BebI8XsR/6s8qRl
ikqYAySCYZyx23knQKoyntvLew4R/sn+ZTCgyx+Tn5ile4Frlilic+z09M5uCHbubl+PMlTKpu/t
DS0i8i/58l/dzRh1v/nPgShYEzRVVz25+yI0tUrYAWszVy97u5iYG/ix6KhEIh2Nho2nyhaC3lWZ
n/Ie3agNalDrhk3t88HjiW5R3PqZrlTSPc+ty12Zs5oPPANrmV0mB7nCELEN7LfNKSAsyspye7JS
rddGJGEBo50EjOdZuDEX0pxBxk+DaQ4gQTpLThoITA6F0Lm9KuUHQO9XQwIPPUETqQ8WKjMVqhYK
APax2quLnu2IZndA+jTd0tmZImRcNiaob25dFDFhmqd1R8k7bxwY5nV40SNdGQvRlSc52G3aIYtJ
XOGDwEQPJneL81a+CRiu7ddRtPda9AqstP6CcNXQcwe42+Fnb3p2nhaw15AdaY8Nj6QremYko7Kb
ifCKa2XahX3U+f7K7pe4MIodpR6u3xFxJh6oASGbeh8Ald3EhhCPLiPizHh1LHJ4OdO9ptLxcH5G
5bN0NDifEakgbjLGenoKbxjUev8OO8vK3Jrm/yayco6Fk3zQi2UCFXNOVol7sa78iotqjDX+BUbi
qby6nhKCC5a1tJfS45vVOl3h97HICrKP19j2/IIj7PXGiIz+d2gyhm3CEWWiPOlAuj39OZKeLFh8
tVo7DRzXWXaPFDpkX0cm8H/HCVMJREAKNNGe7hI8j9wd4S9HX/Oe7EiqudtMYWbP9I9NF58UwaKs
cV9dQ0+NfR0BP97fJMgdmJPr4haJ6zRTeezDgJbWes9hQtUMU+RjHD8uwgwmxazvap5iMqpsT7yP
fUTYNS3yG4kDRhKTpc9kMMkYaX1Lajn1dgxOpdejp2XBJORxJlMhMOS6KLJfLvaLlzn3RXFw9SVK
vPWpECDpmSib7Z7I/t/hmJmc+Gl6ZzsJuYZWn6iZ9JkTFzb77Y+G+zWMpFvEIxCNJKHHlpv+BANx
7BF5P3Jbu45CIKhoZjbdvOzEM0ee/I6/YogqPeKW/d5Okt0694vJR8m/uR/uY5JMBlemLmrNdQf9
x4ZL9Jz1y1/0/HSJKg3e0yoKjuFcROYCe1XAs4HrbkG+C1eF0zXKkXvJzffrTE3baCDsB+EaBs6X
wADoY/YgaTsio9MQUlkObP88A80U5Q1zz4vt2GHW9eNYq/VnzrlyMageKVdEyIt5CCh9QlpPvv+I
hG5eUZhPSjE2eV5Fz3y80cnD/DmKgYlkdkKfeATcUSGUfpyBovsECxwGuAWR/n7OFKEDH+T4cshu
VtURMxD6YRC2oturN17JV9hqWAiXl0Un8xzCwMwzGo0UbWmAMHbuPB4/N/OLao4rdW5YKc1rwtx/
7M0Wl7hRkHIvRWu9XSfvwvE5y9W4VEYVrA7ltsW/2ikG6qIa7O3BbB5zwwjSR40G/dVtWuJxbM6v
5ojvC2jCMeAPLo4uNLlXltnoBZ0WJ/GpDL2KbkKJO4zL0FHKjp9eHKlYExC5gMaqoeWl9k6E2bvr
4GRWkDHwXrF5py3SUcvaCjL2B/XVubGlGhUxUjF8tDp8RyntONLQGfoWZfzL1AdeKfTkK9z1mMt9
CYX8SLebf9sI3vNm0lp1A8s4xxYWH+R+AxD9tHrzrS32M7ZQUw4tA24u6tTRQJhLKVQZxcm5CIqM
58sQUGhhHA6US4pAOKEVtydlrliyvcPySbRcNHwdOf0QUFaffJLCzratdjpt4PgAPnWoYdcdpQPZ
8smNuYxXed/z7kwNM20WMEuf2yah7nl816Puz3Nkc+HX6CAN6gy+naMqWUYo53glsDOXJq1VG9WT
YuY0UPtws83L7+BR2YHwJe3GdVoK4usZRhZuUnM3Plt2jQhv/gEt4QOu/tu2Xje5ODhc0CC4eEXf
6pPoHInD1WJ7ZFDHtecAcmbYkqCaEGAJID8w4178c6fd6vrqz9OD7cQ/MFZrId6b0oQaqfiU8bmh
mnNyCcglKHX2ybZfXDfMC7JVv8bkKlp3/stUwzqb8ps87rtA51pXvOPNjboVgPU58/OP61eGRjtr
eSwnYlH1KE/OQ+W0qxeGXVal63SU8kTvLJpX/S9Nq4A5Gn9/aHmbZnGwnkBpmJRKGRkjyRheSChL
cnjuZiZ4Y5ajwTF2h9i1UbF5veDCoCDZtsq25EVVfN7tUJMIvquDSv4dcLg49k6g0hS/2UxuQH1A
p1b0KwPECkpy3bFMvNEc+Kr4y0w8dHqAGK46eLAt3a7Dmr8uEH95EvcC9MwUOLQG7wamakld55Dm
kAP7XrCDJ3NQ9DuAvKTe3kw2MsMj65jBptwL7okR1mXfjekoARzTdZkMh1Cq0WVKeJVa8r2jF8lG
2MSsu4hLFEifrAvL02s6/L4pw67eFcgBLxuh4wHy7zwB5FgW5WfStlf8qaOQqMihbTkwXnMdOKl2
MDEfuLH35ocknv3cEHc7b5G4ncznjsAP3c/IXuLEQSisKshj7LRRRxCd4LDeQ/eOqRPVJxr0x0Ky
buR2NkKKx4wRhwz+uA7Gyp591P5sCTbZFZnmUlxXtjHVlLwtGF6Y8/BDHb2dY16eW515YWSMfwMa
F68Geb9ZR29ufinWhSeqX6SslpfwrwwthZ1YQIKjWljtkctU5v008hpoMXyFkjduE4UH+Ed1Bqtl
MeY/ilFZEv4JmpaRiCs0Bq69zgImEqzmb1XxCP/OfG/r77dNjhPBEh5nBlA0uPI6Zzi56RIBUgg0
ZNKktrybfOJRLfnhZA5bzIPm5pCBYw8T/FgECscxGuTKP/oaoYVb+S8a1SiL0aL+sE307cGVIv3H
xzU1/kpsvFKJ4So/KfVNhOnf/X6gW0/SEMyCaver+cnPtXKB3NpGD3E4YdcsNd0Whm+XOU7QB5I4
fzubRCe7sE9whNSDrkUrZYV1Y89GpqJ1Dqk5pcd9VHmqvMS/CEtKUk1mraAn/MfnRkRrjz3OjyMQ
UuVwYWOExn8w2cyCXXqWeMbvGY/wMainK2ZuvZ91kBQGaNL/rn63OgvFjqBncotPGIAIzJ4xmoRY
xTRHS0ac2NPtBqTHLzr/pLMSG/olX6+bbGXktutWsPxV0jeOiPU9HdhofSsFslK7BOQkRMpu5Od6
PZ/SuPqTln0N6uJS0XcCFbBxagL5xdBh4oCYiZAmbwymR82+joWIrq+5oFV+tbzr/N4jtRyBBbOt
pnnLJCOsfYo8YXGh92DCDXb2Ov8/Pqcf3aoGxD7TqzG389SgVctFdjCP8baEhHdjwb4n0zvUvw==
`protect end_protected
