`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
kT0+6zb/LcwfgFhxXQFK3PEuoz5vm9u6rNhr4cnhMxhXBMwS2h5oEUZhM1M2nmgk2gRLJuT2puYu
WmXIl14Qv4mC8BzQGZiaInw7i9LQAbYfODgYufM8I5Bum69OYRTqSVC9j5f3EfhFHZrmhjNqsh/6
HO0yPRoRKq4Pmi8Z6DyHdasidR9cZIwbQsMkOmTw6oSqrwwaX1WBei8aoHAOtq0DuuImOeP7xajX
c/gWQgSyk7CfPnChhuy0Eh9SCRU0BLa7GC+CJF/DnJfNxdVUJ1qFutmeQqT/xD+MM6VTW7XlYyfk
YdLAk/tusdQttrAChuE8kWEzzXPmwxOOGEfKig==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="JWPGIckK3yqkWfrSIV5LQfCuTTnqjWwhPwbYmBGO940="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
HUlJBBMcr2r7WLGDsClFFoyjWwdIx49oFEf4J1ndqkD35Ci0aNWDS09eMUjBkXXZsqWpWVelRAsT
d3rV0yMjJ+VLBDkRpG4Qo/pZHSKgDNV9TOkW8MRs40WIELrdv6c2qw2d4510PiLxc/Oo/RpL0frx
ST63qn7zcgHCLYDDOjgoHsa5grAnnpjkewzvPIgWUfNcdTAfzYix0yzO0Pw0LaHSwUCvMGkgsA/H
LNR5QYZi/hFjt5/i9py8SgXfJJDS9yidi9E2iZRVeIfcUe4NiKizDof5CGFefYFLKRPtNdIOzbCk
MkfadJFt+8r9BdZfHVshvRtGL2HZbYG2Mrne/XC3Tq2uS5evj2XV+i/+xFAau3BG5XySFDC+zjix
khGHyZ7IHvC0RMxhPMMLbxhO5JblaLk+EEFJEZ+KbEMDyaC2OcdmrgxvF2S91t4uIXSAVVoMwh2X
bjGgOCBt690MQ5zlQ/roO0QbiJ+Ug2L8cPaL8jDBb3FFDZChD9MepQZvu+vgP24rhmsJwFL5t0h6
aELJhKOf0F8RA6h+g9xQPwEEejNjCapZTTCT1c2WOheTGU+mOOxDPIxmu/DvyDvrZcstSSUMZQTh
3M5DNlEhKHd6orrzSJZV+sLRB5SRPtl6wXh0r7pv8DrjDUPUyLCkWw/qLfpqXSp7KDgcbBJJLsxv
vSS28HXtkNYdAnKnLB326GdWMOT1LgfgKVcGMMUNsQlG+KGRibwwjV7aOqXyQXS51mqBUHB6d3EG
Aio4c2mI9tF5+L0WVJNaQmJ3tFAybMGDVgPphTiEijW9vuspA4pm7czrg/3dizLuO1E/LHDMxOj/
1W36Up8Aog07JEf7hNHjJqiJoiNoNfFca6deATKR25SyJMTgbvk/Sy/91ETyoVl2TPSiR26PeMbN
ZwSl7mkscWGCw55Np8A/bIU8P9DxTgAzETaBAAh1SdE7hycuk7l/mb1E4jcHISWGmUV5/RFhBW6O
hx69IWy8kFHV96yLkd1+zUG6tnthHpAWOZY/1Dc4U9iohQcagOtGndMolhqaeIS79cC1bWyRuPbd
QUbvncs7IYoed4ah2wYkjVt1W9t/zi19jMPs8MeOcvk7aOoR1LcuMKgSmlg1FMAhl3gxzYsAvhuK
lsv0R9IBsDsBVhhAXZU5NQS5DaFQ/t8D3IoCfQzx6pdTceJvMvXWuYyN+HlxazvRCJnpVvWM0TOY
Zi+U09GgrLWNtZvdbP/eUK5RWFn76Ne97FXaMVcHDxaPuql6TcW6u+OSB9gRLmXCBvkLKEoQ4aj4
flgajGSB5lNycVXLIWZYqlrxGjlal0mfbh16jXc2qoomF/68u/XmEovfClaJiB1/kmXP3DCq0BSX
X8gHsUYuqVrYnReLTZGD2gjUL33I0wIYBzbmp8vbcXgb/Hjb6det9qtfqDupBVq2Fc6s+QsRX+19
dDv4vsR1XeQ4jfjHQ+3zixJTe+LRh41H88uHcaXZWJmrfWnWJ/9GaMlyOHZva0aNkjAeh5r2ZDgE
nTGfP5T6e/DjDkdljzZPB4aNza0zhUvfqLGejCpCBVVfZydwPxx/R5IVjcSj/l8D6sfWc+P5el5A
YB4+vEtnZDkhBtB4jLBkTN7MVEzVsJpAFB6utk6P28Z/pxLk6rI57vH6rFJ0J1K6uTpjvgRJQDJZ
py12FhsSjad18bEoXOcLfMcZM6HfpNffWWlV1JeBKXzEnGYdeiikx5qztIf8Zp6zBCVm9rz3pcEx
4jJ5opNiZ0UvdQa+i4S5UbjR6gS2ar8u3fwobNw+kYQSFjd0USZIK59WbFnD8ewogFiBc45yCc+o
rlNEy86yREU+bmfBxjWVqJQuEFL/6HUiznFfb+90SBKUk37HFOM6E4QgKQzjMMcghA9zl8Rr/7gE
n+dOlBIQMydsyLm8zF4/P8XuvmLY5KEbdYdY1nC2sjLgro0lWGQo32JAVNFAdnF253U4nB8bVvaT
lIa/gxQSMJsKHYT2vlGE1GHCPVFRyaOwD9SLv8KhdYlSHwAWUL6/XLRpZK35k0BTcnhhy2pf1hLa
VKs6jE1JBLVY6QcWGlbRZo9o89KSoCRv7b3NQe7RxFYM1DictyyaQkw2SLUDjAiyWl1BvedhWqZB
lugIzia5+q0CNsDw0/1ctt/eqX/vH9MsgdoJWtNSIIUlMr1H1gVByXfdlWbbfqSLgz22OCoqQCfu
guKlfxnZeKAqOmP34lde3iCxfzYW7bRltk5pIcHLOUVpktxlVg9mw+Nu2UZLcaMsSAvy0wTLfpBq
E0CXF9H+xcpF/VMVp0MvcDcREsdSWJdFUhC74IgFWF7CowJHaPchB9QRUExDweQjk45AOYQT5IAo
V6jzDmf+fsDmNeKMG/88mnPt5dgT3u+lmnQZaP//0LM3MvmLCXze2ROz/PhgcH6DGpIHj+QVa9i1
79hUlAwlVaW/T0VDj+HfICgRPe7YcGpEI3VuaVfyowGtpJSOFCAnwr1yB6S6QSz31FT8UmpSsn57
KU93+QfEFiDalO3p0JBHI+0UJ1KGyyeBEnOMXH6dFjV7ApgY5vvhbKqHsKgWxWkc81Oye1EYPoXL
R7It0qDQF18I+GomEwLFwJflYRfCVZTk9TJpZJTjGs0U6KAaJ9P2D+YavmZqV/5ZEGUAVkgY8aR0
0Kd6BuxlulnLdgaoCeZHiHgr/yUdJLVf2KasQUHjL8VWQypBJ0fN+RGGdJEHqi/TGLnPWXDnwVdz
UCQ9k+uI8j4pePMVs16a6oqMNsFBn7hLmV9az2LVvgM55Gs0vt5fREls+pUvQacEQbyad6+P/Sdd
97WnVjPmgyrvfLibt6MOcZXGhF9KiSDVMVGDdUNf298ovaFT3RB72gjv/I6W6o/aTHTkAlpnLtgc
llCMnhf1DNcKnc3lQTW5YIy0y4q7c78+WB5oJmROa6cJ1e3TXhBuKFPyT5htTZeXkGeQNaeuty4M
SgEEyiLm0Yc87an3ummw2Yow2n4suJ/iBXRuVy9ToRPP/jsJm6/U7C8YFJjmgVfm34x/DMMIckew
cfW1bSi44EOzrGYTSqSh1ZgrLTVtiGmSytMddq674iEA/3Qd85BQf5402a0GFZ9fqN1XC+kI4zrj
DlPHHnwQJfDkINlowv7utZD2e6DKccBfGW9JTr0LFy7Z+1sQqYh7sgdUHu0CYqv5B1xYkGFYRehC
siyLlIDyynaM6Mg8Srx21/E5mB75zcNPJfTxevhXbo9QDB3APBFFJEV2EEmj6vP5V6bRk7MjS35a
QAWEX/i1yOdjjbbRlde01v10KbKInMPaJs4rzoze8YsimxaGtE2l8NxKw/49u1a7ym3e0Tnldm7M
JlC/jupcEPR+ffXNcT84WP1D2T8j594hOwFy+7K9TtstZc+bx122BiNRNOI307lM7yVkV2yOG/po
trLhv5W6MotQtQ7uvzV1iCkuAyFrdzavJCEEiJa903i5dl8v+zqNBCAn3PCUu7CvrAXUe5aXLpfE
5N2ZxoxniIHTmtrtwPazehtBRXsT9P0FVNA6uQljunjovrx4+Tf7/j6mEMNnvI7XRCBoVLyeP5On
vgJ+iZ5xhjkpkZlbpSlNtjETQNX4+u5GJalNjgtY97jRlCmGiMTVjTAkkBUP4+PK5Fu4gBuqJaLt
ezMdRmDkxYcJm+ockFzUXpX+/J7pFXdkC5XIT1ev0cKnA9cPKUfODU+uJaNAbB3l1EP41O+5ddOG
RYmXa5Xs95CuHAlFGQyVBbu72t9czGiGf+2BahX7QAWE9lG5Q11daP+NeiX6CctYuxc0cDaRXHH3
TORFx5aLPq99cw8zeQBXHM1703OWsqGQ3VLol0OAgQ8ZLmsCNfUVonDhznHcWR2Xn7hYETyA9nAT
oCq8Ch3vmMkFpgjgOd1hU9tFJCB0eBFKxjxwCaSX3IjxcEcHPHT6ZpQH67pU8+kBvYvKg1Q0ULzn
07lD6/mu4Wrx8TB5iFgc8p0HqvwCZB27+NDPkL+KweH+ebmEcQdO+daP1cX/w35cbC5/na712Meo
QzFnAyME7tXrXKu0K+41+O46kU1cQMvTiwN4FYHYyD3cirnwKbkZhIg4Ws9jUrY7OYh5w7EKiBhm
qbnm2um8JE1Ta2e+kiFOvQph3FDc9/HFa32LpJ7pgX82Gw2wgtjTsAfppZOxiBXLWtQcRaSQdlem
ZFK/9irXTzAKl6aeZGrt4jR02OzUBCdAAUC1nV9wJ3jg+bxy/Vg+XT8OggXkbtki6+hLYlQBZuaz
MTMG64ZkGFEDKKS3D2qJine2sVJz4wPgEsX7ZobVMhn2KUhVCtV48PIFwzVrWL8793tFwc5gQttA
KNzBkKBLcfDfbg7wWp5tqwwXi5OAkwCHNDOaFDKYY+g98qrdrvPLuUUlAD96M7A4mB0KnrIdL/cf
wiTtNViA0OFrgr77b/kIsmUqGys6VFnr3rdTPASjhapNozkqdGQ9HAZcQQk7eJMpJk4EiiN5RmYx
2Q1CCZJW2+XNNhGHCnMAmBpVnowDDjKh5HxIuWf4BoLl2qs+POw+VMFbCOBtLTvvhF0c9dcdUyOG
GN6Soj9ATFOIlXvwN27ypqvaOYDOGeZapnXY4zlNrgpZAzYgusu0Zq3tb4vhaP1gtBawGHOlHvcR
01d51XFVSN/u/uYfQu34Q7V+XuoFLu5DGM+2M+IsMNcd0fl1aIx4xaVcCPeVrrO5qFWmiUheLWjq
V001jIddZPaV9T7ZwqtQZvxj5/QRvT9CNQFvyre3yIKG2GSrVugkVFCRJ+pgbEOq3m1YCtG5dGGG
exdcGFAhMlYOMyzRTp0/ZFP0ZQz3SXKheKngINf1XPwoJnLuKNYawfkUXRk/iHpA62bLQ480I9iX
C3iZkqK1h7eZ/x9qlY6eP8o5IxlJGuiVpXfDq3ny7CMhJAmLsZUwi5WUHUrGrog+otHdydQclrnb
qW+BstIWZ/quPpqcrXz5ha31qIDzEx3qoagNC8DC088BjD32c+Z5gEbFHgulhWeMKMI7+/SLHiI/
p/0Qv89nOD9a0c9HbncwQPkkYku/zF8Wv1e6VC6JzEZoEzEL7b3/dCx6QogDF6oJFr7G2S4hMGdd
m72aIdI/SRCqEcFfZ3pv4u9S6SFgUnSEkHsGtpdQHLfuy71AZXBYJKhYhOm0lL7nr4DZWVn+9nbN
+puL9YHITGrKZzIzN+7qZCurvFiveXLIiYQMrQJ67KIeacjRph8VG+DHQ67ibZDChUkP0uwUxGHW
NY9CNqq0XnokNcXTcra+U4oGfEYhWPB+Me2d4GPOk7xOJt8Nz8OIhsXi+fJE+RYj0U3JbhMsGNQW
0iI+etoEwBwhxZqlp3bJQhEjfz9UUOinqNNzEHvDwmDeaNKy2rDxCWXnbieZAeW8tCIcnSKBcrDr
lQ2U/+/ka+iSTarpR5f5wHerNKIitZ6FDzJXS18Cd60Ohh/CSx3N8R0QkHUV48e9UYUXsy5Bjp5a
pMURDFE2zJ5P7+BK47NAp3zO49UGef8OqRcQmTZHKxDSPqD7Z1J8JTFjsQ/7TJKHupPMaHCYuPkJ
bKGkROG41gV/BgpPE+W+eVt7NJgFgwhh4i3FR/MnKpy82i2QgcOY7MYP+MnaMjNnQK76eSgEAYPE
jw+u9JjWCpnTgUdKr0l/H1RNw71rrXIS/BEE87TPVRXH6h6Jyb2SRYKUU+L7CLXqNI5QRF+OTMsw
Dq9WUYlErIYExkBYBgo/XZRceyB4smhRJGE+Zb9+J860CCIizuwAC2Af63fdbJyTfobWmebfla3v
eJ9W0tVhybBYCP9zNmZqFUTsBabGDXHoC9h8YcMQb+jV7WAgD2ysbehwgU5Uok3Bd5WzXdK9eV2Q
0BhX7ZovZUv5qJi7biqzJdH0GoErvv3u/L0UU9TK8rkZ2DV7hNi24q1K7eEoY2uO4KH8tKu2rktQ
FfGRnnlSmR8VgP54T/j2bnQ3BlKwb9ZxYUVOG5HV2553pZKRsDqOOgmVY9S+Q4fA7kA3IhiB499/
af2ZGGJwzQ+jVX3eHjWeiJLrbo7kiGkDPikPq9Bsko7vU0APVgzm9u7DEgkDLmZGqM0HGhIGV3nJ
on1HS1m7+0dbB9sZ03JEbdhRKQedDA130ugU1w+Z2bHgt/sR6bGNASwIF5yD4RFCqSRPEjqEP0L+
Jrz2h5azq+NWNFRfqBT05kyuiS4KP/fo9bkZBV0weCRlj6VsCUjPnHEpPOUQnmURc0IPLnbwIXjQ
iSoGod/5FETOQ9WYYnXeJOpLUxW6RasK6mUtOa/LAT7cwF14HqrvCMKKMiFlUmmlsduFlkfyOyGb
F5vKRwfSnQspHXHFaxOcpVurj3HXf6MUl17kVjRoAm/pDWLnT6cupfIT1tZ2TFC+AEbL3sd1yCXK
4s5HFkt4q0vGb5SXKh+cL1AuN0XYy+Z4ksduRzEbWqoZRRr/Z+bJoVeDoWpGGbn1/ZBs4yke7kIt
CS/lNRXSw2Oow31CbLSP9PHQBfFe5v4ikAnYENb15eY0Fxg6QxL2+z0sbwMfsVrErsat3hXROnrv
bdeBVVaJ5ifEnQo6JatfvWLW8xX+2EwHSQw5RkmsayJrILEDC67/qnCn5hKc+sINHTDQUBAs2G+J
l9UoQPmUAlyh/6s64aAv6yWRv1FQmxnKr4VbdkSfYkN4v2T/VGCGHK4po3SAVXiK/LbuXDfWex7l
HpYGRavGmc+6s65zdpDlyA6g7zzAk2riIFX0IgdM1K8BwkbAlSovu1Bt96vfFCfvjqbYbmC0syEF
H+djnBwINqKln3Pky3mfNdV9FbcHn09+yUSWSUeYU/5LGPe2sWdCSV0jBKd5A2LL4SBsStPoUujL
G9WjgH4fTtSvk5rxhpzRLoT9zd8wbXmbXUxL8NJs2SOWGZVSNJWbXuUJGsm+cS63K4SXaVAObVVG
fIuONI2WYKoMbZ/DzZ24MAdu/BJ3y6OnSLwoIIM6f+M70qN86Sx4mscxjsv3bZBvm8gZrfNXMMN6
PrgaioDEQxMdAbbsUoLV+fdINnxhlWyk1078lhCj9BLHu0fiMRswQNU2YcSjxYN2U0PInNTO+4IM
JAm1X+MhUKS6BOtDj4XWhOboTtgxCRIXIRKfPsBFSnqFwGFdQll0230tIFoHmTjCVSVJpkrcog0F
UNNo8mEg9DvuDl30RKV7P//7Kp+4EFYfERxmbTIMxCoK7Hjjtx+9ajzEoh4Yw+LqoBvtWU8fOMpt
t9DirPjevplLSA83mBtinJ9JlCDoPt7n1MCSxV7nuIwiOWGoZi8pVn0GP+9GoBYiTRpfCaOlCabZ
hu+mtADVYaU0AGK9fJY5hmC1kLILXxxTwSmvLQK/ZzCW42b1OKFIIIrGan+JzkzX/mbgMigVdMWI
b3nhGoBhk+3pCb5ykOVmFwtKADdxc4ICO/jspvfFM3koFSBQH23O8ih77Cem3g1i7n3z9r3WSGwY
n7rXnQKijs7maCMQVekavo4PFZy0Khnxq5rrcw18QTpH9Rjj4vfuu+Q3qXVtGQEfO0E9C9iVf7Sz
SB2cBODzV1n29z+9RKLbL70LxtIZI9CbO6dNTk/w5rQ/uKSEx8dlbyVv/tOtLyoxRwfdsz1gzz1i
T9qVdxBTAeg2CcYRnPmc81Z2kduwY6imD5kr3kXQCrLxHkH7hagNhukT2B/R/vw6QvQESSV0OKzU
ge5B/QD9HiGiqhWANeXr1aRVvwq6gAs6NchFu+IBIDpDNP+xLleZ1u3aTZPFxf9kj80DfeGjEtMZ
oyFCGa0XJCNfdj3oyjCvZZQQMyZYaktj0aYvBSuzbCMxmKCK2SxJVIYANXOhYpELvfJ0RG6S58xC
FRu1KQ6NB5IHtCUwCC8CedP/AucbtSts5IC0muGBPZKEu5eECXJyXHqwqZWPK8UkajqdFS1ljfy6
LYYFpsgBiC/TUDceB1tkMC0S0j2kiF0fuRKGe1Kb8ho45ja1iJ4BNMgL/ieQyVfww2v6Cx94wy6u
7F0gHlIgeziRpIA+8FnTGmLd9DW1RVhKMwBWyDe4C9d1xkGi+Pb6keHi34+dJdtJwVUuRnzveDoP
jeK6fQMIs2ZnzcngGHA3kMGX2rgQmz2FkiXCYPPH9Cm8f86fIDVvzAX2gKqVrZYra+AITJ4r1jH4
Bl2edkzur257AX+fp9TcJHFxZFkCozHfK/0bDW+YahTTUHl407b+yjOSKp3aymbhtXKMy3i8e9m1
ZldY4jFcWpIWpSnXLuGQwr3wPD3QBLKFYWp9iFB9Dk1h1k8YwYrKCEwXQkhaRL3GjkPlWQY6wv7v
jMVptBYaBlrhPgeKzbv3Vluh8MVSPsMPFOWC+3kNH7IL0WPZhjuCamNLE/dbCZClRsu2g7Bf6bFj
d2duUJi6t2sZ8tNCeBzkmh4WMJaU8wgw84DhmvqX5c7Mz5P7iIQeExeTrwNQv8p2buw1d82tNG6v
bTgC8FE+hB00XNsWdEVo4mMLcOZU1+EY5PVgEghLn3nulQsLrGrxbiL73xV5/q2xNJVqnEMVoHHK
7aO+TKNBfqE+dgnBzlQl0cf+339hRkJcNcta7LQU3FRV7kgUCgpbbKR8V6WtLZWwrAZ/IsSA2Cxt
3qoTqjR2+I355vnSsfphwCqvPla1vqT4vCq5aAQDYEKNOfw18SzVqwXvLmrJ8eqL18OhoOCoUsba
5EcbleAB5xeV0jo2oQTUQvHGKTj296yryKiiIv1dFuxiQtBXH9JP0IXZioWvaiR1Wl/SLwZnkuz7
JP3+QMgyk9L1FZCifkfcG+S21pb5S/XKXoT5xc42c5TN7eIz9cWg+/GquJLzsGBNNBTzAnXKOWKr
IHlkPDueVWFQy3jV8ESiofL8jbiz4J4j9sJohHBm8sCwB471fuGEyhl2zYLxIMx7dVKsy9ptiYjp
/gOmTS6hUOv0+rAaLhdga+lZuD5DaTFJz8nEP3RroJP6K8YQ59SeBdTmFc40kv7atJ6zUpWm2x0I
YkKdjo9KK7eyihD/mOzr56KeDym/1x1QGeXpAz05UmNVn6dXIjFpn6HRbPOD/on1wFjAnwt/D8pa
vjTrXzybpM0LphhNq8hML1JvCelE8mnXeibEtLRliNKO6A+DJvjpMqcRDn475ralSf/R9GEQcdIg
u0diP6cY+s6b01TxY4O4ltG+BxmPSsNjPWAVQ7Pu6chiLnTRyAb09Aeq6Kk0KZK1gACzXcX9+S4h
0hrwDcUZcVO3zFzlPoQIX+hBbOxJbmdK5L2Avi51uM51ax/YnC2fzHcHl2HAQoP3k2o0W9CDaon8
oVuc8r+PqoEatNzTvJkBfwHU5xS2E+LyJ9UVbufGZgo3Ca9SzAzJdTJvlgrOailwYC5SdRKP+O8L
o8dex6jXAxTUDRO49yW1NIzFFPxSwTmMZ+PyOmVRCj7N838d5lfTzPJSDHfruIBd/mpF62PVLU6+
ucb4+I/FPRL2Gng134qdw3FVvNkW4YYqYcv1GHvvKTnw8u2DidZZYrzLpE1ruuABXPqVVQ6TPsev
7y9sSkNdtjv2VGnPQBPq5FTLqprWhOz45j25+N1yschrD6Nrje80vZIRWm4oq1G4uXLBBNCJwJNd
HDLMzLJ2ZL3eDaMq9eefrYOWza55Ufus1OVEjBYCKGYq1lJktjvqCVETodmQgAzhLQcDxcSvyFKD
N9Ed6w/gxIavCMS5lTWOjGNRmQQQAaoRDtIn0arexhOaBQkv2tdt1mfeb5QNJIIkFriCKix57LWT
Q5U10RPufFFm00FtOj2oiZx+NKBMxF9nDGIQI+etC8Dtn5k1a4PgjRykVuGqV8ZP6+ssd9YsIJat
j9ODQN6yTYzoI1onk1i0gKqH3yUYSl9Blk6Spu/USUtTYcQ2Yg/0j14UXpiGEayEMJarT5g9U7ue
xkCNwcGVbhqosrPNFmaBX7SOWBChTdACJq8h3l4ZNRH46O8suDy92fTuIwI9GWtaLcx9IdPBmnXt
BzADWz8RxFtkqUrUl7cw70Dt3XIXbZep5VkX6jXXlGOH4INAnLaRTEQK1FzsrndoyPU9ekqXOSS8
H4SesTZSvRY8WDrrmKnGRiYlara+nNSAxGHmWkUMU/iyPifXN2dD+HkbeOUTNxrEN0AMUACwy/pI
R27bOgZTweFtgFxb0UpowQF2h3SNYNUNYXZAdYerlZe2m66v/CS6SLKyyLvG3RdtNCwRXxInMuWD
s0gp9kUFq4NwpN/0vuEg7rU+/WRQlxKR18SosXcIIC027r6We1mu65tRZOPp+IxLLrmtQUN4zLIM
YBWaZDXONZFkLKAIRhu2hsN3zzWRokJMTyzrygj2D8mbkytxJk/VMbRstwChAzs/h+weMZBfZj7s
SyYnyVzGXt7vIKp+kMPTHz4mgV6SwphU19KlTLZyiGcBI8lpHUQw4Y1y/bM/lP0HIOe960f+O1qC
0GTL1p8yt9S9gT0QqtRWetK1OsMMlxS1fAfx7sTOEtKJCsG2lrsftn4AAyeQnh3nhpdtrJ+Mh6lW
foFakamuFE9qb0NJuRyKh5+1/+/CoZ3NflWOv6WQKWTBoAbaSpm3ji9zutczmLWbqD9XDeXJvUm+
CPy6obdEtkX2MEm6Sc0RjDx+pUXosFLsy1GjV3q6NMrbqBFmrtm3KTLbd1fiNohJ0fmP7zMVQTLY
Tkhl/6klogZSQrr7ujJKIEcTxwADEnQ1as9jFVyZJq36ketL63uYPisSpuhc+FZ4qplkKeJQPMdf
XGjJvGx3LDEuL0qbLgrShk2kEPmb4ss0Q8IzK6LLRAuSAliDmX487PDz7vibCjO6/DqKAgENjJzD
Tlu0n9LG26A4QXXlAQzNeTjwlhAIxgAXwuIXiU5JRqtnlN6Fvsw2+qDdNc3sLp0ATzP8lqrtIHue
QPj1y6ZI7seseH+QkKYRicD03yv/9ALjT4tRYHK2NbGndLgrsAIEMeYezCgXR33wM+htoXvgt+0c
2xgSFZEVZMolOHSgL4FzYkTmr4dV28v6NDjIKuvTExa6wTAkljA0hWCYymPgXeNaYoFKaPDWMJCp
fZigdN/9AE+55LD6B2SyHq5+AI6Jdvy7+d6bQ+73H/7WewCyuL0k3i6Q87uYJQxi7ta1u4eE+xcd
PgiW97TfQdrMW72xjFPyRoaRn5ya5cTbKnntenBjHLvG7tYmVmX2pGYIkTFdZgyirLiWUw2xvQUD
cehAHUcjly2sko+MuJUr1CZxbsirbtCypImq9J5BxWG9cNkwv5meq/nc7dcKiT3UIzG1XKpNeSu6
BiCpHziS+ED404x+isVkgie9xOn2xpx+hmw0cmHEsKOaX4wLDUAKlZ5B6oORkLDgtdGy2OwoMzf4
rzkgaDs1U40zDniuAbOrHFxZSomch++Bim1yJTuHqx6cyPjF1QKGs7g+nVj7ZR6wnw+GTidNb5Es
AiGyr14YQtLhkbhL0huefBfCYsyJUVqVUHJss0BVOu2u7natbIapZvJ6YSE0m9zgJ+n0iwgCXsrh
lXhM8ZhhCWFjbG1dZ3H8TWVGitDAj92YGqS7ixAE8nM4KElRdMnlgKHe2Be/Waq5WWSiTr5wxF3y
uWEnpZbfAIWIwTtdweiBj5O3KjKNKpGvC1J1TGONnPyAqW40x0a5tOb2aWvmTf1onlti6yj65W6u
AEuRqNB3Ru/0xtoclUJ5+OofvBufFdF8fzNJrAikL6mwkLt62aqvBB1c5hUZc4AW9sfGlqPxCFPo
oAoQZ8kIANOPPf5Rtupqj9o+ZrhFq1QIDpafilP/wQp7MrkaOzZNAFz0NO7QMyd6mZBgljdDV64x
vFbn+ih1WXqyh8jN7A+mhtSn1FVEk2+6RPEHVWBAXd9GbSJJn79JL2HETNQdYwQ4XRNbYZhGOFh9
MopLMPhMmXkoKEQ7l7nrm75qDUQPEkCmOT4M6CIKA+NZqVhR34zeXBAMslz0+0o0NgkZxtT52Wez
p+b9LpnP2KkgujEiKiFWhjBDnJyt/OvLvPehgz3gy5gsFEIJDReGiRinpJhi3llglvCFQdHgEcZ9
vdQAQf8PYxIFce+ruyNizC9nxYuC4XqOLkqzXXUhRt7kfYlDB/RYJaNooTeLRqxoJufHHB6tn+aL
2L5bHi+Af4mp+eZlPe24WJWiKc/z8J7Dj2gnF3z2Gs2qC7Y+BSuABrcVJyDEEs+W1e4uH3VAMrwr
q+4IeLu2RaXe+DspUBapIclWQ5XIr4jRLcbJleLPAMJGFb0hBBtu3dYgWakMNpm/EaCVSYQB31TB
lOFlXR8q9V23uaKIE0cvgyvp16CWfGGgd+xGU0/TltRn8l3P03ZdgX7hgUWCM/z7MOWhiCGkfGdK
gQ5CPlHmEKl5XO8ANxjqt4iUb/MqMcZr7OLTe9LXwBhyTAqh4lA3upgNFMrMTbKJv3weLOT6ndW3
iTFQFHVXt0r66GxXK/l+HLYNSLl/mDAWwvRl+IWDe2h/Dk5pdtcMHP/5MjRVJmLZSds61rz4HUN/
NX2WOnUL0tKOkWU1oqs2ujyWYIdH+bbkujGE9xvaXqE6oa+PSxfqCEw76Lp6qGsPhHwtbR5Q+ZCa
VgaCfZM5/cCKMiR1TmG6FH5hUN4zbacDfnCE6oc1BB6UFFIS8wVv1WP/IKBNTenl3j2L7Ci43MS6
Hg1eME4ApNXCKs0yOxlz01fNJGL+ir9LChU8ajMQ8q2Bb0Rrj8b+grkx92D0pIcHhrgjVZddkBGw
9uv1GVnfOZhEDnjbuJqRMxaTo1xPsGg/teeXoBfYNadZZjpxx+gIukfGNBxfDKwId3kPrbJFLU57
s1QmhOoXqYeoUynTM9Y6Mte9ZyLYQcXNF/MI1kbOE8uSfDfWp+B7hwwZKr+toTIPZqirXtP+Y50e
Gz+ay7diFNzBtA2ZnTlNcOutVbSVyeSw7O4nEMvktCv/1lVXQFO7vBnj+uohwVQz5kvMhdDerDw+
5YNMQMGDkjaMJVm29eBbkuzVs4ZJfghX51RZjLgOrnUiZExxXMMom/1bnLqVchVwkJC8CWyqx+iL
dscJtXBPnR4rLx6NuxEhZGkgOriqFHQAunnQGYLr7C/lLUDqCE798BzJGphROIp+KwrIkH7FxMrn
TcEkF3Qlvh+yR4Xvl+qZ8Oz3rz3uPtg4+GYwhbG7pmHvFtx2NbEYUeEKgDRYp7Z5C14ihE9rs2M6
72eGIcJNA8Ikl+M303Nwhw1OmQ0x/6bZzr7mOWOOme/wiUbDvtBSxGX3DKFHr4hlQrIa4IDz1bod
E9b5yddlr2mtb6Ius0DwZvALu6kx9p+VIGIoKM9Hqw+P/wn3+D4zSfyw7r20johvRvU4UEPZO0FY
PmueZ0CGTYAhNTjmgzxWHU69ruHHD3dudA==
`protect end_protected
