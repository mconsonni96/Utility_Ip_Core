`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ZF2TSl//TIBq7cfr+0d0s56xE3K3Bsm2/dyFhenJVj4ETRCjXSzBqcoZqvzbUP9J4PTuUHL3azzC
LByYXW3CTClI2q1yly+BkmqzFvQ/E1FlspDnWqd3VHv/A/mVNM7RMranDCZc2cenZpcQA+LVPq7Y
IshkhoUzC4ik+TZXIMnIBrXbab1vxqqa07GU1KTtduC1pAxzM0cFt0ZN6kiFp4eQnXFw0lXtp5PI
0vLLi5H8iPs1MuSWh3y6psfnQqGbV72A6+GvNtLz25VNRbJayW67nNsN3qxlqn3zIdser1UzHk4n
7SYCJ3oCU8hWw+RADAqJojsv45058iMqH6n1uA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="9MfS+0qzDC/jCVwAVY+oX4EKqsrZ+/HPcjZwOkQCcCY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 385344)
`protect data_block
A1nGSUzbc3ngtdxEfw96wvfBaeIPyVMgeLgyt7LGsRj+msfPblATcMxJc68apGagPDzw27t0idPt
p9JYwgThnmeQPZj9GquwM2XYECdS+A/vCIu0sRShCL74BLccLb955Rn06XYgL+D55Yud2CkRaoIF
4v6UhB9oSNYoVw9RrQJq0hhSWh2lGSsMNsJl0r6fZ93mOeLjrWauZXEru0TyboGLcDZGXKzAZYGR
3eCnlc9HGfZZq1zIyMiEqNsexCyGNHkbbUqUV3Hgq53L/UoMgZwkTtQkQc4IpM+LoHXFpAKx/HPa
t+nX2eXqZP3ROmfvfF+Xhci7gDUyqAI5y7gxt1N+5mPnsXgzMBzRZIdBIx8bhq7t5ZhZ0fEGgEx7
dcWvYWggtn3jBvdwUWfzq7/tGV2g7YJgPR3McE6m2UXiO+pk46nTktrrkKt9NZuMRfAk4edJmnmo
hnhUwjO1TyFsPHCC71XOf8Rfdkz7Ec5fA0goRVEv0IgTviUxoBNrsvVu8iUUgwvsnM4fGoYh7J6Z
4gbKOvqRek8HFUHbcuanEHFBndVMT1EMCbgd4qVe0lZl8gOCsiZZe7DlFNDbenByZXav6UAJ1FBH
iZtddbzFEfph+L6SugmHLZ6zlpBk7JcC1rp7+v07vtocAyFG27tumiIoIEW1Px5agsc3OBkVdyIN
RExh88OufEe7EXLluUia0rnzDGLZcTntc69eiolQPopHlQBY+ngt3psWtl+Z7vwZDWq/dr1Ny3ku
WMGniyrgBepOKrwUkhD+f7a47bUuM+o5Lj2zmRmAsGAXnegiXi0RvMIsVdpEtW2Ivvl+HGG94yuD
lckgMpCUvava5UoLgltl83fUHDW8GAK0i2C6RZZaqdNByCsaHT/qD+v4xltHOzvsj81uQBMoUFMz
HPGdiO9fXdkcebAD0so2XCr4ijZe8EMDugHfD0BQRVaDa1WmBRKldHk8wu8y9HrhtNs3dMpnRws5
UkGFhEkI5343LRuvm5l13yMM28a0ircYfNptE0enaHLh8kiF2ofZJepGKADqmaom7yEdHppe+oC8
KNBkEcyruVpAA9S5D1qMbCjArgm0w+v3oNtNjRCxfurNYWG2NF7ibDQDj1wip/VJp1ILgMxvYQ21
DScHMLcXgRELlSwt5I0O40HYfhwpyGRuzUY/6j5ytP0owCfeX0jdby7yfYjq7BEVbs+SjgBG/GV/
/bPdqqV007H7bunvmiXHgnKN707RrSFJNAdjSKxpUfVynBbm/PDMmx4aI1LrKMZv8hqLDAhnrAeI
zvfHuwnSj6vdkhyqiA5LYo6RuDGzTcyiakoHmSHKJmf5h4OSEzGxXutcLmRgwEnj/wUH1p/HO20N
sqo2EUpg87Lqpl2gCtd+LCyPqYXAmBJs4SqaSXbOK9+lT4C6S8KgyQowe74lzGB1b0oiCKjEERHC
5SIqPX818pNyMKymkR5Lv/BPmn0MB5CATLvCE6fJ1qG6NuFi8Q4sD1kVAU0DLv8xADfvIkpY7oMs
fl6dJguEr4rYXyBpw5ioYabe99o3qVg/fOZWVltqpx/+Q/y2a2OP4pUpsbHRh8eVzBhN/Kn6W2BY
LW8MyzUkX20+bN0RF0Plo5lq/eoRItuAFmNXe8Mvb0gIiEXVnZtMVlw349UbczMT+tDBcqnloM2/
ZOB8hQchO/E5DoaIlRHtr/Vae46B4TzUDkLqxoROs5Qt4Ls/ROO0Tkpc031xmhROEBUkOkR4SulD
l0jJwnQkUzWdekbzLeAXlypZUgxHxmt+ioDFaC6uwiKtUeWuedO/59ajl6dmj7lQD/GXyFEuZk4v
3XMCx+FWE8t3uPigwiafTLiv1n5PMq5+vxcD66i8nlD83nClGW7rdAErKtChO+N9x0L4twyxjBX2
pSDyBBRsqcZMWzKkDSEFtFY6xOIMz3fiQUuvn2qrztnxmUZEXTFWCO052u/L6ZeWjyh0VSUlgxOM
rqN4E5DpG6HMqVciCd2IVl35W4/uZN/kBH9YZ3C+ORndQ9XaPBPBhrjPbbFIpuTPKS4Ugp/pngEu
rfn7XOTruRPPNUu9Kevce/B9JWWfBluSSq4yFoL/907rFMFnRpeh1R4uPuS5rBj7GCBJLVbYNKN6
rAD4T5SS+fNAXEmhjRi9ZX8ZMzJfmjkTzaFwd3EuHArJ0nbrJsNaJRs2EciGkqrrE6ev94lzGIP6
6GKPc3ZN4KyCN/yo8zJ+bYrWxmhLMzHK004+v5BkUjiQTprZoOqvwcauWmigQToK90/kk+f3LH3O
2oqFJxZZPJNKE5Von7UJvGqN2bv+xHKAeBVc+1s4+eL9u8o4YY4mf+fzqNC8yjfq2tYfTpoq7HmX
lj7fzrjiCAujWZE6323gZ6XpBFKbMWzZyxAqSjKGhNQeLV6wyvzvUFui8YXri/MQE0/wZeodgPPz
uhqpP1IvGzB6i2lCcL1gGIsc92SN8v+Z5NvI4/rTQUSDuW9sjCDYXLNY/AbEXCp/ZZ+/zwrcDVWZ
yMeFHjQYrQmySsOkaiBInRhXP15ZOhpRrSBxJ9iOSjGA13N4MF3ayNXDk6qZZxTmlxesfb+IPDbW
Hm5f//JterwXo17oSKBtOHED1dMvyy1ocgpzQiXKFuyDfW4tV5b+ycFOpLyfXljtHK5PKz8K7A25
BhGJvaAJ/+wvu7qPuuiZsm2FmAC1cy4Ufb48hf+QLp7PmxEE7B5Ft1JrgvyJOX5bmDtBr2c/ZY12
OJkcFAMInk+8AES3116oVJkf81ZPVhAS5jcVKfZZEugA6QvL128GtdwVyEPxeQBSYgWG0hdsvKt+
v6kRBDqhSDgpASwCk9Aj/42f+rhacmiKh/e4AZFdYX2ONZu5hYBo63Qn9jgGx/htl6vyJ4OtnPyY
oVS6BVofRT6+MqJFOgBBINnE2ueYzXmtDVqlERsvCgsqb4CcmeZSnpXUdwQAz3RY3PlGLwup9uoQ
LDg4rqYc1mE+7bjXHhWNYLQTT64coE9SCTdViLGxchsGZTi4PQNlaeNceZcfiWmQmszr3DkmJpXY
GFdkBJ8GLAaXdtUKoGSEC5XppprT5R1yxUi4HcKJ32rtRqqbNUBSLshgxZWz8VOLs6YY+mD2ROW/
y2rFngMZiBcNSA7W3BSTipA7h3S5+JlVcPSBOKyYKXZDv/5AP9xCXLPAam952tD2bEq9/6+R+M6C
IXQkW9I/peLXKlhrEpMIbKW+LtMoA+xjxBLhNt8WCWovyx7eVPBZIcMS3UUM4YTKulGb1/7xPy3v
Bu1JcL9V+aaWiN2DsTMH+Gu3h4u5e0y4a65N1k3AZsxxZLa9NE+aBz/dnIo1hpkVsDQhE5yeM8X2
rKBETtVnTeMpKH0eTlJWCS3/HxQ8BEYlRQ0IW3YCzI/PPsr8eNVpOWD6B3A6vtmge38NCYx2Tnix
3TYMmzCtYjHOlzQlj0VKt2wO117F4pZ/ED3X7i01KAGc4xe4uKFuMMF8THFRwLe0e/PRetw+1QEH
jZ1o0WaTxl3Grjj47vbE6VfDCwLxFwK2Hcxi/2pzcxG6Zq/gSVGTVN6wMri55Jcdf/8CYTe30m72
UdqYP6ZSXKyOJJh1yu6tyPUPo1xVXgqhTnIKwJxa3bMi+fcQqpX+ofrE6CBzrhIDULi1PGW9G4Vx
P54vsirEPw8i/EjgQuW4LfFy/q7ClIkx3ci+snS9+DDycmXOMni8enYE6EAQT2Jlp0MVifJnZ2+2
uwYG0aK/w2Q/ZLs9IE/B8jOY/vxQI+Ph3O3tCltAknMbfUbZ5MP/HxpSY3IY/VOnR7hS/Na/A7/z
jhDmj5PfijYWffzQ+riPW5yd8Kdg0m2+J7ijlh4AsioRvfnyt7GgQViyK5sdJ21Bh6e4Y+ZaRW9L
xahqpBpw0B96ZBkibemGZnmWZbk2uNpQ4miraoXgOkhGm97wFhiVeV4V1g3lIQhokR44JABdsu1O
LvjDjji45gVQEsgcDzmLmvKs/scLDQJUtapEvCm07kkMrA6GVqRYYnUFTwjjsaV9LQIAqHU6BDjQ
QSlrJZnepyd3fWyP4tai2BvIhbE3CLU6ftUpcTEYFNWLY4LmCDy3QjY3DpgFvLp+tpMCtaRbsoCf
8lyACmY/yYoA7EecPL97kiCHPUdgcM0TbAu8IEKLXzuxIiOWDoBmcAmWA7mwE0p+EhDrNAkPYBn8
G5RDaGrWhbakiYGO2bziMbRj7s/BHSV48moGePhYCgXf03JKIeNnE5ZAJQagFHBamGSsE2CzPo4m
Er0VYpwZQq9E4SHIjppXGDK+VRYBTBbgB5eaHebs5BeSMCcPvQpGFMnR1bhhB9KM4rPCS+CB9h33
dukpcIHI3aQOS9cVLHVxrvFRmGpu4y2JCEVMpiHPgShAO23gP63hd/ykdm6/Tj72iGFDI67rtiQP
bdflnOf4MbSKIP6JYSB1/C25VsuyOR7DlvcLGCgHUJcSuSVQMOEvEdEgLqvOIof9dGihQhl8GwHr
nu/LhDzLrsbsEOsWbXnRkZVQ1hJHYxqvgRz3S3iTX80XbDfQ3ADwlpJOvwFz/ibndSYrZr/p5Diq
pe8ArRdRGyYCoTezAc7P/l+v81IpOAqVghhhkFM2jUiTXSc3CO1gVKOwa4Vv0iJ13ijwwdjAK2Ie
QbF3EfHMZVlbkdQwW5siaqypfF1p2Wj6OMbXL8ksqIzkg+NKvi2RxCTNTouEqRxCfggwmZU389mq
GwIMWcj1gaRiKywi1QRvvA42s3YQWnVw5EQhyDYOojvRIcI+06qaCQWFTENXsD9oUK9MloXZVGbx
9jiDwi+6AtmZhofruRc58YZYHM/Usar43eHW8S2eRu0P7fQUr5o6usfHu43O6G2TsIB2Z+/ddHR8
MSTcUuw7jR6c9cehZ8ApjehgF/7ObfmJKsflSzUFvehQg+vvzkgYOVfaXAsy8x9cCbbhF1TkQjvi
/EQsLntarpc/M237d3shMEwwQ/wDDm9zS/g3u22qRrE20yIdb0RqoFLUO68vfUpYuBywIUIBG7Qt
TQ4H953D0j1+YRYDoMS5jAvGAYenRyTnuydhVBPBVdhRlrmi/kZOHqJ0rCcglQsa9+SZJ6fRMCp7
LGITFZrsl5/Fdc9lXFWBklOsQHaNX+7ueTOOdOJ3PGiPn27GRByfyF+cVUWKq0T6s1XAc5AtuwbA
LmyapFzFNkAZoYQVU7uCVIfSTUVnx+Uu3v8cp3Df2HNfBQsxQFzkcUCmSh0BwqBtQWBw2hMquf4I
VsI50MlPcgzm2zESymKVktojk2+zzfSAReDc4/KppXdvfdMRt+lRHlzQCjIXLAyfsuqZv3rB1QOu
1/WLzk7O+SrJ4HhQPsnLG8anfUxZX3qJqZt980f0LUmXZ2iYOUnhprpe7EE3dn+IMblU4Ow4do3H
A0jX2i6QowCPE0KcpendQzAHePh6T0jMSkHVzhq0/SW7X1xBNSaV3lbBUeuZ5aPFCrk8J7ugfp5v
EOT9PJp3q/ai0OYn/RPkIHrVYfFUGL+tDe+l6bfh5tsy/o9EkZBxfmDBAwxqPnHhBo6NyV/kvzGH
D3iEW6GrKVLa79drHV1ThVH89PCPOVW8NvZJgq7B9kBYuKzgm638g0XgIwdZ/VupfxNxXQb4KO+V
OuvD9L++nrY+2dwTfMdGqsO+ArEK7ja9GSYbRrmo5LMC1p9NTOcynUlI/QrfZBTxYklyYW5x55YH
9SvGHq/CT/xm4/tAMYHOLsP9lJ4oRWc+3/zcI8QG0hHuYs7MlUI2frNPAtU6cmj05EAV7SMrGGth
tJwiVQ0HwRfQK2o4dBIN+EjQA5OxU+IuG90DjR1WuoAPFnJazzgfd82FO/16OtQWHCRksRNoEAYe
wNTPz9MmfXWGFcFRAq0K3Yo+t5+xZRMGAtRHLCIT3OXnMVPpecC5ZVRbK/jxu/f2tUAXr6gt47el
Vw1fm40Ad1CyCquXtm0Cnmnx5XHw6hrlJyHhw6SXb+myh+4eY6AidQ/4g0JuQsYfkAD40pfPEma5
EiwKZu7W7LOIV+LAtsDBidN9Ewsjf2/aAGWJFMAUhs/UUSJtPYPrKjVo2St0gwL/4O73efWpgJBz
ON90RQBse7pLERXvT96NVulDTwWe6+NEcIQc8ZJ4aTJ10+IIsOV5mHVLcoQvmTqjX6RHU5Dg0RyT
KvbiioAy8TW/F3n8C4T7psoJRdqkmvblGWYKk2gLz47LYfTFKvdMJVGT2hhWI2JOwgcuVJFjchIM
REAn5j4qyol/+Kavo3krsfImmT/8X0roKvb1WDbR71nbdhVB3fo79IqJr+K3Epg1xqmfdDQQLmZG
1Vh2ame9Vp5n1BcdfWZflArmCxWEdESkw929ZPKxs8CahGoJuPzx8n9ym/ufS5upB5vlNYO6ZCRR
tBhMWfmGT/31bQ0p9V8Ir4ooCw9Jv0f36jn1kvJusiy+mFN6H/QNVFBXDx3/DnuwHN3r+mr4ine1
03a68tE3YIrlIrNcMliR8mcIBNffGRD0+DHTkpw2OVXiJRroLRXyfO5LEzUqUm/KURBDqYO3HoWR
SxbpjiHwniW/FfGHQcra0tlHMPNrVcEouB6/GTo6onI5e1ze5bgf7sCrwYEXySnBuOoY0BWd3m9b
k5L+kLRwVYWEhqBMqKLaw7ssStCemmlJ2IsvqiCzhKN8HhHGVw1YlRF4ZBMRCJGaKqex7c5AyfIy
hNtaDBUrdMMok2lGgYfBfAFoDnPMm85MGYwgFRSTfXg9TV4pC+z/a9ggyxmXL1aLOEFnlLwYu5U+
ELygDGDwMH21qSj1cxHUz1VeYUEdFhAOuXqOKfsDXBJvm+UI4tNM4OxP6PRQaHEsI/3yY34ExziB
AaSiXj500pEmfCaa6CRsIaIdk0xeEoOR68fcDTCMYBewtKKk1Ns1oAhS0eK4nTMaz9MU1ziIeA6b
quPtPGLPniBNl23X8eHFlKtEJhYftolZfxoaWPyEW+zbsHKbAtrwOYVC8rH6nMXt9hMWsp2aH/hR
x/vDWJEjKuzOmPBT9UIDtDrK3Dw4p68W6wyKn1JD659dvSlf94AoKXErmb+UXz/GxOk8SXmnAuqC
KiGxW9OhTmigorirlb7pYYlA6AH1sLvCLRQeG+UrDaOUimREHNrIIlzPgTS6uFxl9M07WrX9TTof
PhQNp1fumJJGeUuuLk7o6i/nyFIcU9CHExjPIMn8S73c1DzyDMm08hBiKNJjLuA3lvJexqlzxWa2
+nWxXuvQsaBKq+l19AfsdH9Z9K85SDLQ2JONDeh2cb5mkrHhIk5fUgFEAgnLsmVGlVmex6+dSm1p
5aiN89Q5L7H9N1ys0toU7q7UXjU3yKcNnNH7T/QnFedIPQcnn6fkqLKuPZ3v3sHS8RDZnTvhteSA
drJwh4opcVMteQdexuvGQKIMBi+X1+38Yw3HaVeY4u7U2Ooohy4x9dSSQJulDLNMQbd+K4drOr7G
0tdvYykX5YkoQaSY+Iucko2T0FOXPmDEihpZm7RFcL2+ktuynR1d4yeXIXcj9b9Ajc7+vrjLDV5i
k2JkrY85l2Jm+FgKpMg/xmRb5Ih9mQKElrbM9JkXvhjlyNhfWBSLT03qjSfNPjE8LMMJ+qs8033V
Q7prUGdSghY3rspSGjANZ2ikZNS2pWNN8q+xKwqIDdsmsOi02SjKbnw3oFEhcFnHM3E1yH+QhDnV
eFv2Vljhsqm2bN2PrpQOZBE870o/Bf/PQAwFQCq843JTFfZQpcyQ4UQpyE922gcqSh87mfcGT5mH
T6Xds+0gs49iFn4P6JnLjXK7qCEZVF722ElHyRr9MLSkM4EfUTQ0snPYSHT6TBkbYT+O4Ci/Qh1h
p235+HYqiUClnACWj00F1kiyul6fkuhn8O4EcHc3bMTvBiJ7weqUS/jyogRlch/WHv9XXzJrNJw8
q+f6ItjaE1IiVPlVzPn4jeFn9RSrLjMBdwhi+wfB7a2JAK1bUGr7kjVwIKho8eKwL7A6bQ6pVaUr
Qn9EJQhDZqWNPnhg9xvGmhyoZ2HFjps55e7jRVSOP1tkho423dMGxbk293MKgWnEa/wGxEFXhJnz
X8L/kY4hxbc4glG0rrPAn9k9h0zxH9y44zsQxwQgVWqkUyl6ZNkyIHXbmm4BoYOu9/efi6LcYUs6
Z+wIW6pyLpHjTXCFPNWe9jGPIzc92QwMhtHVtHkg7Kl6qm0PJRd80PuT+L+xJA6GOjUsgFq+GnjI
NAvzLx/rlTU9TUF43r4amcVnR8n7g7Mq8RnUskc+vU+LOYjFWUXJeqdGSaptzlCJH5NWYjy9Qzym
duMHBEZ7hiY19Sus4jwqctVyFkKttUQbl8oZxpiJovWFra4Kq3DJZcAUHSaiXDtPDw6jNMdIkEH9
1ppBK8d+B7Td11syhD95NlAJh29Z6hEmkPirrHgVl7nbHkc+6A3313clqat+/jLy0Xx1MSrNtQE3
hQUVlCUjoGitU/BC3/xJBx1XKNrwAFGa56oYCXcEHVKA0t5/dCtUzI63mlkDQKg8rqcgVx6xJrBJ
xYWa/s+YEnLLAUTAg3f0oag7mCnwrKwKr7grx2V5Dv+G5O/kJYP3rLndnt1d05K1Yg2lldpEEnDl
AYMIfyyGEwhLaUsOnSTht7ZirwYByoShu1KKQoDsObHHy6GRTewImwUmk68OsmE2W8y5elAvf3AS
nLfPkXuhUBFb0VIwibdum16oUSQ3OIrNL58T8bfMx2NcD5Y/r81Msw0SgTz7mWP3LzOcc5KfM3wD
5V4kvLT65BEwaON1eROfgmlp9utlwAYunHhLPD+TnU+rNsfB345euDktE8NZSrqeKOUAVx8ZewGS
GcTQ90K9EHA14ZeDSY5RiWDfVyoZ5rFrOc3hNVE7iBocRz3HZG56xLsVbwhPvSXmnuuCJGFDLQCh
73CZVoSXTKWW4mdAM/pOLaQEqhHWMEoUeYolN6XKpnySGPKSxdVm7lReSLJnzJd4s9DUTp0lVoQJ
oS1BZQZ39aiZNBkOz72sU/OT7YACX1zu6M22i4xz3jTqCJm6ytIdUz2KpSgMFMh7av5GV2bRXKNY
RG/bVT7K3zYm5uZAavaLPpnpQeyZ8+fJW0O4xknTxmrDPaY4Mv30twSV9xJdMmNq5jP5pF7acB7n
KvTEy3uIIALTfD3Qv361vw/jwMOwRU5IHE6YAU+MUQdCdLfDw6270t1v/J0/1jhQwBN6p4KLDpH0
VGNOOinckO8KfPiS0NSxoD9cPWTyNDGBv8cTJ9nPLI1OJ4vrmgCuFs/mAjYuQrZSkOBP/OCIDcYE
qBwNEOoE32cNlTH2jkk2zBQYxcLBlVRDAyNGf1xQDIaPATjAzb8jo3aGmJdE9ON9tx88x1K5U68g
Ceo0WFcsJbauhS5GwCvuSgGNaMeJiStetmJy8o3Bbli5PRdB0ULJpzYIFfEpLDp2xt/YSO/U6XVW
CilILIg2nnB5F4hGHARGvzybQFaZKepZxfCV+db262OS6WzmrSv7aHnrqYPH2tLGf5CIipWYa1fL
dCFaulFYGClEpm1tPEw9PRvcBr8xhkQV4jaf8hSxyIEd+tdPbt+iFC4ZucJv/uHpD76hmNds69Tm
/nQo42HPALQAl3E0Oo7eCQvVcM4yux9CWYrVWxq4dIM76o9OdOVR1zxiFX6rvZUbLtUkMNl74Vz7
3t5PdZ2K8fhENvPS4pCjnTxIovURcFxcLQtIJ54E8X8Y73QBihDgDPo/O06sdoy9bshOu6SZsgY4
KFwS6CYNcu9h2W38muJBfVK+K4141Cmcq7AID1wH3gOquWd+G1OxlXqQ4vSqNk2Dz51k0UK2HYTh
ER0ZODU5pHD+ol/A3YUtEBKDaUx/jKOnF1CUrv9YlFv/kHuC09ysfnY8AglxJ1aT+hJxyB+GYp7L
sB2Tz4bX5t6AhRAApE7bs2VTvuOWwMsIYs0ffXtTfL0IJY+kCgdA8opxOBXrtgKkba4TBd5U2wJj
qQEXP2/BLK7O8qYc2mK46ibm/dVBiKs/1ThTS6gRK9TdJbvGp3wKLOS20GIenpISMej+3RVzNMDO
cfpwYa1uEGti2RXhg81HPx4LyN83Q9IBZuavtj8U0sH7yPhM10nM/AkNqqX3YBvaQHtmKicMjbI4
J+2oIzINN8zkj4teqlaTyEbeBi/rzWvfGa3MZbOBcT0KEXXFkNDNFr1Cx9UdsXRibuKIifnGlbMA
SVox7Xv3gyUz7HN0htaxK3U9PRdel4sgivJuxKJQF7xDrGK0tp/wUeVZQW53PjtgxaO64M37Kb/p
bLqGOhv8qyRQnL7sy//7clxnxIQ96px6pdMaEWdoGs2muln8Zn4LPVq4zhwDL2GUu4fU/EbCZzfK
l5qjM0ogc5PWwALa8i9Foy16gdODdJzNk95QiwDc4OaLxFCWJnZsW2eaQ4OJgIbZ7P+tA7GiBTOY
c8Kb9vTssZO8L7he3Dl2C6GzlIBHOG4BkPuC592vxQwFlTK7AlD1EkI4Ose/1iusioCHZiq8F3Ht
+tfIIZ1fd/YG6i1eJWgaxGl4zSJRmZ27gnE5p4BeeLk3RMThUQ7b4WgdNpwc/Jguy4KPt18M3son
KsKLH8PD+FRJnnq7M9SYFxUOSLWdiy6zVDxCi7h6g8ACIIVnkWk8fLNan9sKscasVTJgkBP/Ju6x
eu/rBweZhjCpmXiMhSmMaL42deG21VlT6PYCLg/q/qvfedoyLYW58jbf2yA0dI0ZhnGHvNuZd+w4
Pw7tXLlAsJA3JAKWiFygvHecReud2pJqWGHxvd3PM2iydAgy6gzEN2C9Xin3brxTTScD6NNL4x2A
odpn5fK2pKWkPvPuY61+Zn71XzUuJ1MrG5X5FFfxPiRWV1qFenJ5mW/GMXjNuDPtI8e2Re0tdJKg
Pa6ROqzAHeccItuoYUvHM2bR15Q+vAaVF5Ynmu//1i1G9J8CU6/nOcQ85bI5Y7ltwVR3dNdLEXHL
wEwypLyU97R8vWo62hk46dVT1ZVwaMyNhhHXZsyRvyhIK17gma3lV54/8O3O+POe4ap2aMG1W3t0
rp//82wqIqNUodfecGZlvqKA+9ZcmIUfmaAj6MGzXr6eBF1Lkfe+dlyOwR4WcFDzAxMdz+gKPrLb
AK416FS2FVi1dfo0J6VZiq9aLmlzsKuy5Bten6eC/RvCPJQS4Ls8IgZWSyA4B9485pdVxgzw/Eg+
HX5SJm7uUKxnyQ4jvPoxulJd24aV+s6954bth98nviYHRCohELfZGoSLNHXQG+PKknf/jfk302xM
BXhfKmjMjR0+juBK63xzQEF24rS8UlSVDvUJ+2VAnA8K5rgbXMERJoCAMW2fomnOBSThju0MgI3t
rwbg99CYGKFkgLjFPIqILOYMs7xq5frW0XWf+vAtMyzaCC5ItqeExFi37Pjr7WPSvQIHyuyDVQIp
nnVed51AlsjB1cpRifSdszxtt6Pn/ehc+aZlIab0jor3Cc/7gkGgnpgoxEN4lY1HGkOFs3uGbFc8
tAn2ZUEZLT2l+iBdNFLf5T4HhG7zJ0PSptvzgZPIChAejxsfaR0bshOz7n4cBsosypVBF9JoA+/V
sdcin3Jt3rXZjEGR17tf37S2BBwxEO4sV7XxcYTJaep+b+rB7M5ZOid+i7EXM3uZCuzzsJOjpZ06
6WyD03bytruBqSVbk1ZhAfopIaxWjB2+mwfqiyq4mKmxwPOJx/eSvAMd1krkDoaakFm0veRIti6l
YMe2Z0PIQ/Qcp+MJVRw6AafaiBrMb97CvvKH85BKYZibPyVusG0cMqxRqtaD4RpkwxUb8+P62A+7
hANAVLkIjJ+D7pmLZBbq93alt9HRLb8rjrIlzTl6DGRS7t5k6Y+gVy0ZRqmZM+AzgQ8bp6HWKcTj
KxVAacgBr2KGDggaqUBWqg3sR5AEIp3lylGLKoO3V3Qb8X8MU81NUQxguIpjZzSxg6/WpH0TL6Vl
Btoqf2hzFI7VNLABVkW82Nirn6CAS36+Sh5VxqsgKIH5+PvqyLLANyBi5XESH0BBOTpfDkc+y+LI
dFkSIxqKDiGpdi1i+ZwUT4CrajGUyJ7hs0vEM/CM8Sk7ca7Kfp0Mq1xxwDZKxJ4PvGByd3+76iwD
SpH1fU/je8/wpCmOU/aW8JvVSAlzpLFmxfdHEYGmu3wQrNmIgLzzNS0TZ06eWoe1nxf+1Jk+mhjO
HZETWe46GLVzQDHX7tQgCN9Oq1XNVFE2maX8cvS/USBeoC2NeANxB7jQLwYkgO8gVPYMB7bD1pVj
klyDIIGQAFRiA8+sH2N60ybABCxOvWoSqZbkb3V1UL4DHtWrlMp8v+mLLu6d2ZxtolhpBLGFGPdB
0wCIPWQK8/OLwjDD65i6CF3djBMq86GqBCCHViXo6VwBUyzV6ZBYcrs1EgEcVOK1Ug3sC+VChAoO
8y7+9Fa8qlYv5cH4DidJ7X717ycrrkKVLqlxuYpFbSq8TnhcU2RnTTMQk7ZLo0RL0BYgqGCXQ0cA
TCOWNIy+5j8FUuPSXcxjSqL/eVx/MSmGJhsJyK6hBoUt2y6yvJsn//E3VkY+HykkAAn9i6X+WhZU
J2g2ezX8wpHVQbIvZUU6Gs2hOvLpU7Joo/a6qsRrju1yPa94PumdX6j6e2B/XJexuJvE5JHFIALI
XySnmpctJ1TO3RXJvO4z50dwNUQr2iYnNRxJoB9yp4TbLZ16t9GB0oqj0q7PQq46CDk22+uhPBou
W+lGoHr1UoqQ+F8UYzm4f/yJ5tS0q4Rx7qFp1ZIqR2MNvUSkVLZzdKrVfcxapEOcoUJo91gdXpy5
XYXXwuhqX0rAHWInnIrI/JlvNkMFhy6+ak1mOnANeCd4yf8HO87FAjEcCKWKlDv4EnShU8+M86KK
Q52R+Gr2FpLl//xp9JwWGP1mcTrvJqhwvCaXUCDGuL3iSAQJM12eVmWTu/56H7F9O1o4pvYm9dSN
i84TEyQ2rLgdaHDY5lUDdaL3sBuTWCNJ6uvXOry/ND/l+6eez4WMNi++VvZHEcEXbGHVpq2f0VkE
CLRLWzrYiGvIt2Z4ckx95C4yKS851d2B+qXp+fi/WS9RKOQZQcIluMQSXNhSsbwEdoSl3FIsf+7h
EkChgJJbYPS1W823XWvx+M9GqEi/T2IeSl5PJcbTAlRR0fW2LN2a3la5fMfxhTU/qRZrhtV/lbQP
rUuXmzX/IOQzUq6UCmflHIV4Kh5jTEVZwWelu9OP6Ys2kUwOL6mA9f/bHKA2X1T5jIjfPCoLIsV2
XDUZiDSL0krq96ZT+CwffZz3rBUprSFA9w5WMRkL4JFKReVIMTUXiYXLPbhmJZsPCw37sYTxaGKM
nAD8EXpBtPfO3fzJUeVHW3iBdrwEypluM6MC2HrKhpYwfi0fMo3NGEueup028hFvuSXdTb/2Ff/G
lEgn9ftuJgt/CKi1dbUm8AXApZ3jGxJSA/7YNxUtDf0ma+BmudgPgxL4mwdzM4PK7NfKbfYFYRpy
sYoHrb391hspGMBZxhG5ug3qaeLDGTPCcfHTUB0VTi8jyBupFy0WJIiNoDrPwWjqv6SHWB/p6ziQ
92GCtyuo/cLmqLvj9nuzc5oA/5yUOSBO5lSsxBAavrW0Z8/g398T5io19uCHbq1nrtuGAi4YtLHW
bSVp3qToW7cV1gpeRTs2NsSuVan9kpkdkHe4KyOAnMOhK9EtLWOPJzxarU4IAHnx5lohFXrXRYKv
SIrW+n/bFvepU+lbUw4Wf1wJZcukISGqwveYCD0U4+HgYBubiXCSJ9jo1dI8SWNL6xhXlS6hu62X
CVNQoLxSmSTMFE3tE3F72x8z/FPLoeNyXSSrj29zpJlqKrd0+5j72gYdJTyY8+FIfPPaBGRla9nO
Ae0BS1Uyd6zA6z42Yyyyl8P+ZAwM5WMbCb2B7Vqf29yiWQ66JUD6Yvb3N5PlvD/aM3VKbBmC9srT
u6DFBaoAE2vZ6mgtq3Aj/rh27yLI4QBY0urM8m3uoeCOM/e6SeoEoJajEUthnkv5B7n4y6j0BuWX
R2c/LkuZIUNDI59YwF8fT2ntZLXQpvXv7uWtNQTrSo4tcKP1hulO0SzxG2MHnIbGdmQW43EzTS2q
DdspSX+ufMS3OPOunZk/XjYwdov8ltaOzoiVsSXqwcftY99SKp0aarqR0eJdnez412dSpZKsTECi
3lwLLMqtrFYtgmXobtZGRIFy+79/1yvb8flHQaJv9ioopprjru2zZvYnd0Jnp/3/uJ5xjs1ZNujH
5/MJsl8zLHhPBlefujJtPvbNvlJel3EdzISozjPtHptiJ1gtDvSGAIfRP8iOb9vSDNdmcJUZHZxx
ez3FEkGZchXdat+EnsjYr3u/8kSOePUrG4AT3LvxlonlufVCCpxLbJqfAWsRcNb1PbpeaoSn2lvd
0UrK/n66OTDZiS7K9v8HBT+YpiISHMoEA3qeF2DieJZxxYdEtYNZ9NYCbPtA0E5NAv+EKedcVMwk
S1tMoH8cMx4VQSAPgP7d1oHCjrzq+TXo9+S/Y6fjXYpYCjBnRV9T3uGD96VXLkrpOQi599uwjbFb
DIX0DGChMDHo6FjuxKKcpp83DJ/5ZsShtiNmVKhGFwyBzNjAmuqEfohYHr9v8RPqCrx3Mv60zcxX
d2kaKvOxiOs0pG950xUswlQE1rW8f5amKn0RBw/2kQXzLybhgwLLtnjgINDwbVeVQmDxgWA297RB
F8Uu6dF1a3yWWB/UrJQ1J6Bi65sOCKLarQCLgGMhlO3RKmjHpa6bJGvWZ8y26Cg2vlK/GtoN5kOf
+V6+Jim0qQUhSl1LLnZPy6l6kQZVi/pOc66HUHsJZD7WgZygN3kbUtmnoSwyyYy7d5R6PaJ+pUsK
IQKrHNXL0jaPxejq78GI5SaGZanNDsoElvQMRYPu7HkkYK5l7pw+KouQEEGhOQKsWH73oolBk9xg
bc9XYeP1heOC4O/UKTRBqnBHsqCurly9EEeW8X6XNvMhLHtCd/Hbq7SgLe1Gk3rCG0GvqAQm/wyR
LcXxqOuA1G621n4UpSvlPXIDhMzZZywNvP+S8xVddKGtc/c2DW3LBjZhAUnhKQGsXSaaBm2hvMk9
MfpQHDHasyLZgzsENwhZyptwYsK5+r1pw/E9OoK80NEGFwmOhlVhwkOXlvlyHCLi8JHx+HhKXYfJ
JzthM2i0MM08SOpuwiUjiQFDuZlxywtrUOaJ3HYdwaJQkMyZHQmXR87dYr0rQ0VnWmVmlGa+nukY
NseG5XiOzuS+qdFdix2rz/TPBpI6n72KBFJOfWMvIV5o8NVwjcAkxOxsiEYdx2g0mqiM3BA0tNJ/
MaWeABBLqhzur8sxTuty6T12DEXODBt7gpQE8ij+VhVYzEPIeyhr5YXIho1KYTuQqtCZ3xjjdelP
IZ4WYoTHYd1be+4Gy5Bk4Rv7Q5It8bM0bJn7V1ALua2Z6xv49S23PGD9PW5gkLjMBl7nxKKbcnjy
MsY2P6tPYW4iazHyCTizCEtjPOt4uBdTWINTvzTqMMIhus/aPl8ZW0WOgdU8x8r9YguZCaAIDWbm
JL+JcI/7XZT6FbDa4m2le/+hqsLJUp1S0Bfp4EeUWDFAyDEhilaxEeKSPMoxfzNgtEJ4YfwjYhMy
rzlz8c4cC/TEma/hosKbv6rdsxtfTy4hURdPpigEGL3lSe8P81xWOK4opUovcnzosrq+eK/4x9AM
REwk1GhneaCqSrARGX+rMbXiyjcfFrd9xmixlOrttl3emcmvU7UouIXnDTa7ehK4QGoHKJrQxkIh
kadoOkiQ6oV4GZd2kQpBWjjgbJnllcYLrFMlVftZ3WZzlx0eU3pu6rLsjD5PA8k3qTFYEEnHQfv8
Rfp080KIBf8rMjtU4kwfpcAPndaTrpPhK6hwG6hYLZrn+XQY218Ob99gJ28nGHpdJZjrWyM/4TTi
pdw/u+ak5iXSeZIhz2XvohGLrQTEW/Cd9fDINYINP8hjaihK0YgDIGKedCg5EicK2FKlZyaTxt+e
YON6HNHro9nyXlgwTNlm1Ck0Tt5Pz8n53xEFGIwgGCgj5EsZfYFARLW8hIkuW4mfqk6FtsFJqELw
cYTv2osh93PyTiGvypY7q+mxqyZK6S72KpmnGsUBURIQs/DBcncFvcTOp49yHt0ScbfWqxzI3LgV
I6whA4nDMcazKj+a4emEU4g1xblm8Kej8JCHmBv4mdF8jLNf2fYAts10YtKSp76Y8sqV6gobwghM
zhEyhHUHXlOgaLOwhrRqqkPNyUf73LzIsaV848LPvg52GBGkdkKOCO9Q7DlVg4ctEhMr97Dzb62G
XhgNvvPV79Y1nL+fXNukwMKgpaHHsDvSa7geNZa8KaAZslfUYT0sW/ctF6Ta1y0J65rXk6d9/NMc
g59A/tuWXr/PQ+UiVPfIpYlo78DQm1i18zyoeBMyChxHEkkoAmA6mYwpo3Te+CmLiF5z41mwf5vW
LBf+CpwIG9/JeX/EMG9jCym2iCXfqJozBhuMFeiV1vUw2r+GP2JA04ZSAGY/sceLwFcIozh2AYsH
/SiqNPggPkTPRtFGaDPfQIcOnZSo1xbaXGLrMox+mghgkJPtUw5gDN6/GN3z/XxZ89DxMqXaJDh6
Ui15koYc1Kvxv16uuw1q6tbjTOGq1IjogklEezpO4Hbu5JtLY86PPAIjMOCGQgg9NbF7wgE+MB8p
Zlr/oI2uKpskKP+tnSqHWGLCBp87jxE6qXkI4s/V2yiKM6Yk8CoFlXpOIeex0pVLjB2tbewnVyEM
08a2BLSF3xOGDw7670AVicBK1vN3tMW0+CEycmq7rdmD4PxfbKw1wYcYrEBykluXVqBlAd/Cdo1X
CRgB2xpUWGsz2YCs39lNXnBnCaTphp7GPbJ9rCYwFEfs3QwgY9fzyJfknStk821PerXVOj6H+V2F
cRkKZcrLTwdXhkpl5k707IzIpX2L9G9xvQJ2noNhyH3ZZzvkrXiKltUkoSOJYM8Yhd1kvgnKwrbW
qzRr+5jl+W4XCuytj0vM4hqD2lhyxZ02F6htdSyRDLFAPKApE7T3nBJn7jtmkGtOEPqy5jLCuh6X
o0ak+5y1+FOJwHEIkI5SGEIdZ3XXhzs9KyY/pVZeT9nVUD1sixzvYftu452QZk6zv7zOTMaBARuL
KnUV4ok4RgmANK3PO1JWicQdnmV/Rsp+KnkrpWQdUOVd3VtVTNtAI1qW3QD6bGgAcQbOj8WoPthq
4OlUHUjEouo9B3m38zC8ubk3vIX7HVPqwWYy5xJykodcVEvJyzziO69IAO8UwTc+3pg7ZGhYvlbg
dV1FdttL9+XFxdciIQfs+8e6Z8dV4NAnY8y7FJd+vFxqhi1nq8MpllqQq6OtUczj5M5GkvCE3EF6
lcCyjA5NTVgSBJvHxKSmZZKhnEAtqqfxvlwgfNe557LiDV+EUhTsgWTKzd3zOmSj+jXWW78jrdG1
Q/DUDBqHHwuA6x2PirZJwR5ZbzudDhWssns7j/+6Okuu7EgAB67NWOGDRPd1gedsaddJygi3nd5A
9EAbMHzzORDJZ6g6YFnlvRzj8QWJm0yI49WSr/nhjkFNngs8bD0tZoeWKiR5Ei2vSANrHbjOAvdU
xyRN5SrNeRa8h9zuFWrru/Wb3x7M0GKKGbaLuuxjuytVr5O6ZFZ+QxTa9LJNysVpTPJp7YusI4NI
ttsRZ/dRo4Vkajui9mUKeSHFDigO8mJLQ0YnLzajNeap6eei6IDDimN7BLEvp+KPdwMNITWks+YV
yh2dGd2wVAkr5EFn1k2Qud6XBlWSXSzaHyThB9HsRcUCvDJjzjHlGhhDMwkhMKAZ5hgbxJNLe8V+
AhCPUhrRlLPaI39vbBKROV96eyu5YVe33KmlpKdtl86nsIDpcDXf9lBb8I7qmt0StyZj+26Fbpor
dejeny6Omchslmg8lN1UEhCj8I8DDoJ5N0eKrQNta9uj5sEIoTuNBUdxS0rkwJub1VAXW9Bnhp8c
ARpBB5XDdIVr2axHyiTIhZEnHRNLyQvHUVwtBjOmLY5X24Pna7f8idaquHgZnjd17hI3JJUSBPuL
Z43svr8vn13TGYEPmBKu9KMzia1lHqrrx0MpG1MrnOYPBzUlPdG1SYVbqNWUhJLDTZ/FimmCgPzF
KH6SqzWyIp/jrFMFUeP3nRrW0aT3q+50NSGwXyMYXkpvTFVltBTniP4bkNrGlxUmlpLWeHv5q1zg
GLNIxOv+fFOwUZN+K9gesoYylvFq8/veJ+a0aHwrqRQ3gwdkc7kw7nkVKlQrvY2s39ahHsjYcQIN
FL+EomyOzse9IVjltkdugHeYQgGWT66XjoE//K/sC8qRvpp7JgWrE/UwpLIS9QHSgOSxT2H5ZRdC
dciBUuVQpSySqdWJcU4D4doz6XwTYiqFeBJje6vPwHOGIVYfBiJG8bFzWpeikBbDOSyL7OjT8es3
CNJvaRTQt+k68eJ8D4WzSigeAby7O6OYrclzPO5s7dQBl1b4tnJ43uVkFY42YP5kCbgcoKmkHQK7
jBrBJJzl31bJVfyYi7h2/G2dK2UxXicDxllSXh2ocdjBiBnbZHn9ED5k1K+cVVJ6rxCQhMZsc85K
DV6tR0G/USKM+r9BYf3cAC46A5tJWQuGPJ5gjnIa5K/r7XIs5PySOPffDKeNj+twBdlQsGo0UveH
FMVm7h0DzhIdTEE6G+HZNGuIoFzqDxb0qqi9saMx7X/qQoqomMHJ6+HkzglqeX32jCyWnEvjf3C1
nka21+N8/BhsJ9mRrdyIRFrMHeEbqq2FSe/LdXQtWo94HZaIdDRlE2DngfLCtA/JGHc5H+IhLJCk
7SrWxj/msS695sZnusI/wATcWVKJo9d0YZ4tmPxYiSThjXEWjxbgEbDjuqirEjsxomdQDKPo+Ph+
8nvy7+rf1FogNsPgILA8RGPzXMlIjqSaK5zsi0ndeU+3EvAXzHk7strypSCBpFVoinkGzoAa6dQn
zE/tvFKqxii5AYadpzajGl3gipuIkRllo1/spnbsQkAJniFgLqQf/mefdpdw6umRbZxlHamwFpdu
DQQ8Hu3PZTdWiBNasAOokeWSBA4twm4/ttSUXvHs0Cks5YIgpcfuUJWCMcV/HoT94xL798x5E71V
jkUBZSyjxscWeyg7O/8ZQTXeAFPWOuCfYAgnczv2o+YVZwcHq8vtyzCCUMHlfr87k4sG1fRhlzku
MF0ralkN9jqiliMubo8sxo9Vs1dM/LiqKm0XQeyYx/pO5Pw+Dl1rWtRBSsZPiFCYirA+YvdovYS4
5ey+uPXK6DAgasqq0USMTOLfVwdFP+1gQQsb7uAHJdV61Hqcr28TT/eX6d5/gxlpN2v1pXzncjcy
TlQHyIjNZYphO/oij/S3Nd2Du5GVRHsxfuK5Z+ylfMsPS0kPtXUTk9wFHcFmYTBPX/pc7/wsRnlJ
0dYRX5GNOOHbfnTB4uX2b9w5TkOiBPZt/etAtfHvC5lGAZZpQ2v9fhyKWyebSVA8cOisOrnoEkhy
ng6qyHx+dW+KTJodh0j8Cd4DJbNrlu9JwUc/V2zLbE541vMRWDl+bz+xY7/3obeVqPDYtPTBBYB2
RCkr/CA/RWkkEOGR7+9B1OOcezpnyfTlE7VPXg3IdObYJGr7DF/jmA2adEChdAIcrr+fw9dIQbbx
IOE60bDovrlFS5MvrEfaFAf7XmFfiJuJj/Sk2CUyMmEpH6NukQh5bv8fwd4HXbzw2YYf2ZLOYp72
uXPXTO2q/DgQVNDlkFKrcFcIZ2vawMA+Rb9guA8/I2T7BY94ZqpU+fz99wgw/owErBWxkWcQnNtk
LOHdPZKi1oLJleABpUTlKp29N3vCuj2UgSlX+NKNTcvUyHTr/H4gfKCFLOzBRKV0ia6Ot9DPdFTY
xONN+/b6JDRlYpcTSNL2ETPUBVh+sgHX3TadtVgDIRQTyVBmczXxuRFGynDgYMzLJQyAU4xCMkYw
k9QoDslKth+Ja/thS/IqGAmi0irLUtFCIB0m7w2LJXZjSzNcnEaDME8W4tWHVCK6Ddlp9R/4m/fM
tyXj+sqkgn7/G5NOHwbmISJopVr3SpAyKeJH8URMXV+TMbMoXeGTh+KAhqhMFZ3i1AZf0rdhaXzM
ugaDwhISKFVvOOTSEoLZJ+W9A+oYSezVwMwBurRXJM4Og7DS1zhQQiUI69qubq1Y8nDUtmJvay/Q
mX68L62+fbc7TreDDFmz9gF8qWsxahAN9Y25Wn8haswNpH/u94PIlm4FKt6epWVNUsfg+BGcNox/
gBUJYFt76LsEbPF/gXfIvzPS05UEbsbT0EsbLlQ+KHN4Rqe8lYCsFVRq2Y6zbhD8mgAGeae+XojP
xGDc0WRki6oREvA5dwJT2SxwOy+tsrkP5i5XZDuS5nS3IhJ7ECrP4bpyMrzgNQhBU8tztZ+woCGE
CVEqonhkY5ni3EHHhTG91fpMgNrJwqxZzLLcqBRw+lOCEuiiBG9vsYcQ6ErlUh9dLpcKzSeO6Tf1
e5zuN9VpJCsVyvc7KZhiWO5PT25JbIgZ4BAxm9ERnQBBdZ92vZ7cjZsygA7S3grkhR0B3155Vsfs
mk/SYb1wZ6Il7QIJcZ4o4wQECBOYRnF7ElWT5BSYQsY49583agLQwfWsa55HCXtPkugCPw+2Gb5n
Z4otcGE9j3H/9vP8x/BCjIc474EcKv4V6YTOQ5N4lssMeokKt74eehTq9Pp/GtZBCQYLyeQR0zrE
ms9Rrvx8NyRBWaSy6yKYBdRtBwtS0zmrU4+hryTEMIz4fjW8V0zR18R/NcwKNm5o1AUyUQJ8xJKe
hlf1FcQCibt1KWxY5XUBdAjpXz0ljtyeJOTaF44XaohKbGAaSxYMFSt06xXSk2QB1I5uvoI4gc5z
TSTe+UzumF0BTts2vukunr/L0TW1ga4iT8PIgggbPYJIZTXhpxVie9M6GnloslLa0R25o6mQ3RJ/
qkqN0Y4WKAQB2gDkn5HCNA3MPLfjh/Z1CamtXOME4a0IUnNEKWmyHebR0m7iz9Xr5sL1SdIBEiLf
pyVOSbOLiVg7pNqGYZi0Z4sqyN9qjxDNBchWewRrw0e0ccnAN7oqVBiYP8+/njQ2WngaH0HBT+1R
bNjLE72DcjWiNa0y7sC4TbP1PR2vbELGHcAj2mHxyQgGtNX6CZpN/XnFlfqfktMH3JSJwSz68Qga
8t9yRPU6MnZyhjDBV6ufrIwF1Yq5kkT/ujlLj8RNy5uavrHf+E8eGDDR5TvtZx4UPXr3ZNjsvfqN
VElNq6PQcptV/k6vKvoh8SVHyC2DgeNByniyVpxShYZHGrXCq2Ldrf2qe8AZfzZoqIWDP42lpKtN
ErWHgDdOEL06p8ECsLMdZifkWToB5sJxvkhTwK+WSyi3l6+nzUamh7E7hyBnf1poXGPtKldFi8po
0U4U8/+s0wTHJc+CcmQj+rIH66IeEN/hWf6/dYMFPVyDFVTWYgxq2xJFKPEKKH3WXnNREcXQHc/p
i/1JUbFr+aDtiyUBOqCdYG6tb4xKaLeu3gIEZ8KMNAPIjIBZ/bpS5wXpzPocjmnwfJL/3gWRj3NP
7QSdJI5zl4m8qf8wDwxTgJxyHVdFKgMRditOxPGn26p+7UUDRkQTlFIod/hBx0TJcJhRaty/zabq
PgqhGb6peHDSIQqPgUXyLCS2OLIPjM0qD7kvKy6ilBMbF3egIj6JoTIrhhwkVHFsJIZnacoPfJJm
dfX/3+LJo5Yl8PYda63IkV1GJNonyU+Z6k0w8h1S1R1nhMm2EfHmyam868yyb2Jfbbuu/77DLjnm
TaG/yRhoz8P4cgqYwp8AUTnjDpGRejFrNtWLPtx7xdhJ/wBUStB9pOFdD5Bp/qwk49TNmxMjYybA
FWmAwiTvYe8ONDX5wJaQdgUSgmqKrFtxkkudXb72ZjX4UEpw+2lo78iR2jhEUeUpM6iX+dCBjgzG
u5WEptkOdpa6uJwjGxFRLntukvK3iwjqMPqzRHUaB5yZziJt20TYZdFSHVTAhvXTT8TRajyMSEfv
+PrttOGIGInBm4GdIWDOkUOhhVL8K8xPIyO+0woc8uJqzoNvvslGc+IiDJW4aEcRJV0OBsca3rFH
XNSlyFok9Tdx3kt38lbkQC7s82QJ8R4oLL916G9bOUaGeMqCrXHD1dlJ5OvgvDYS/68LYV55cDqk
VxKI4/GSevxB5Oz6VWxTEeTGWTTBd1DhvzQaemEU9HsHQokD6vHl0TFhsvHLJle5fnHXuTO81+1e
OBLXJCxn323aYgXIYb1R1MteYBL/l0DgEI77PCrZOe/DtdQvSFT+kQqQk8/cWGJt/sIrK9BY0YOi
p6pqGZp1Ke6EBDXDz1Cbvv1JRqvJa7+krU6TcCo47ckXe8TsvQ7/GT08xqySIO6mOnrW5HU89pKA
d/2kDik0UYbGnut0wA4oylF4TMKtgSUzOlrUA4q7z/Gi0eC2hUnCJpRqAjSq7+AcruT1YAXk6q77
a7ZnyBJrUSfb4UqM2yS9IIGmPv+7r7ZkAKUnn/Z27RfSZF6O28GfH9WAivQ4b3N78IcsR2KRH2Tz
GgVqv3ubGM1r6RK4wCZzraJUdWV95aNZ3p+T/vCFF2xgU4xmPV93rlkb47J2N63bjH0na5OVeUId
vPnZWLeREn5o2wpt1lbB3OO0yXZPntG8Opl4VUaBBgP174FjlfheNnCQVi7Tgos0WoJKj23jQdkp
GlgTdsLMzp+X223mFfhpWMhg2fvl7vlYA6lPKUTPUgq1isinHobZCJKLkMt0AJ9P0fRsmZVkPJdZ
9eIrAxbdLrFNQb06stMISiVMJ2TXjL29EUqDcE/TqE4HHhjphtdPTIBlz7LGqJ2/BeDH7eEkt18s
IowgWRNX5J4YvoiPJKSkhiuw2G8NJjFd/2XLX8nv8gnK7QH+fZJz+IDjXTtCawTEQ9Pz4ta/P98Y
Ns1l6ztZz6eLcjiIm9uoqxfevEE40GM29b7Bn3TC91OGxFagBmiJTIo1RP88WrBIeK7nmRWoZjVm
6LeLtfp+cEkJvnYUPGq/G+hbvEXvvo5ub/2+AdriYqwkWZgICC2GJukMor6J64yFoLIJkSvxpBM+
BErx5rfNIcmsVG/2rf7bY/XaDZxzuGT4pe1UI6N8zrF8WEdBCCivEpPQycKsLKIWR815D9X33UgT
9nHmu1nz2QuXIhk6FJF7Lxo+qSAaIKuUFys9byyrsLIF43Xig0Otnq4r1xdfZ/c1qNCT+HmOfdOC
7yT1zEjUtrYhAvgtb4G5veB9r2+TuqX6Y68A0LF2ETofPVcl/wdapX0hXw5uFLRfpE6cy5hUUmkJ
Wr4lN8FO0kwbbzcXlUuuXIkX0HZSgs5Ly0TNmozPFq80S2eZERl4LbxVZzmbtqT3uGE7VIaYJUaZ
qh6OGDVlTApyPPJT/AI6IiCT/1l6ZmBWmVcVa9wuxaAkgKBSJB8serO2SxajcqNEo/UA29YCgwSt
nbflSEA3eHRc3xbjm/yJve2RA/sZtUisnUyxjUmQN/g8gBtXoJAF4bx8i0CwVakWpy6fxLouJnZI
A3hqeZCI1qdDQbNN5G7ak5TdVLjLABM9cLNfallUUP3ISaMmiUzsEtpufQRL/L+KA0wcBLHi9Jj0
MYITJLKLEyiP+GYrQO6COaH4v++BS/xg7+6nKPc5GBvlPOYV0VrrlFLgl4WZNgoJTE6kCNUFGK2K
pYS5ageQDkRzskZfg0nF3NfhcxLCJBiar3am2/Lss/xXb9fC+o6C1flNKcAyDeEo3PWX6L5qhXx0
+3YOihCbrP3gBYpKzOyPgWRd49SEGs01UOOr19e4/XjE4gz1q2Q80eaHYWtW7tJm19/oyRWjr2EJ
DIdOhaHE0z2GHxS8WxSTM6ZJrm9v6OL/PY4kR9MFhAy/6gyDpmA2cZ5CMuuAnOaQ5PfLgZRjpAWy
b2pVKktsgmBA2KHSHqJ6tGlLSfuZxTtdBdFMdfjmOhopkWRf0vY3i7M7z1uGU/0fGKUOMeDHqSG+
cDgeb2iU4oHeBM7vR6RJgyuxGpMS2wDOhqyB0G+TkPfAhxQbTjwPyO6KecLFeBZ+2sE8dx9fVF7y
ve5wzvhz0Ux0Am+Mc8CHEJeTo8wgPL3HXL798RdMttD2q2Pp684uCsWNFYt+ix+vGGxakz1UtuEY
AvBDQLIEBDF4CbZjTJgzAq4zMSqgAMbTHct6vR3FxRoz0Xxs7b17MKMNA1JzMRuLux3xyz9fcBsn
mcJaBHl0PY3Au00HmCZkOlygQS9BBViBWlrwxMcDfTUAy26rGDlTSe/5W4ATjMhSgi8xVFBAUVN9
6HlYe6rMATYaa1wJA/4HUGDxZ1U0ifGe3givPTteC/2+/ADojJfh/XCKSKQ7OuHrUONSr8/dC8hs
jJMJ7YpO0Gr+q/QKn90jUBOGmFOFOqca5pDp/F5TA5tNrhI5Qs4oHaeENino6JOFZCmgfH0UhEHj
jbCi6FxhgAvvJwyng5kPUKLQ3+n8Qge4bpICx9Vu4lVb/Ujnst1GMfludWUikrHpC82XWZ4ULUdq
jz+kkvwJ+0tSLd3+wmMkDdKmkc3I052U/w5KrthLEEaa1ZOZpGXAcvZ1uZEpQ+fDa1rirTxvRXEY
9qAZu44N8dU6OT4Qep8nqoPSIqISVCXBgkPGUeWoqZO2h+TyJtb1l7WSkrTWn4GgHuIGzOkeZSkl
3ObFUoovs1DEpUpKaltCx8lqntXzzlo8+19bEDnVEXS0MuisxU83r8mdaL1bVAoJBZWRvShLYD50
7deH/yaTct7QFu+Jgu6nBiO4ySlghOcCi63Kmao0/UvxWvIFVyMnJSomSpzKBMix4ejUas4bJ5Rk
grpmi3G9Npfzrh3/c2ZIH81YX3f+jATFMaWlWdlb3qmC7MOxzvtN7SBRZTEI31yzjcSvPkOBin6k
mHW73X6USgoaRpmQO1c7Mm7dCvzFIuqDGTpFkFX6OXPPxy8YbV8HbeYb/Hee/CV+II99AtkMkBYZ
iA5A1jddWUqH+/93oakdac5aRexVHGpV17/f7Rfkfe234jPAf53v3I30xs2htuo6j4G8a/lKfnOk
CivHd1QwFtnrdretw6pF1FRgUs4SZs6BrDiHX9J3MoMSCb5zECzHZYBLobBU7nPeUk46HnoqgFq0
DNZQPXOkl3PN9L/j4TCPEIJySgdZ8lygYG1LS7ob9jknJpzQOySx0gxESCfECvlJDOPP5lLnq8yM
bxknau8FrowfZtVyb8arxNqOQ4N9ge5YwzIykQMg0p/31h8CGlLWqkmlCt4ykVYklmJUHXDHxrBT
qKSCNBF89LvJmuRE0E1XDX2jXuYwCeWbDs5jYmn1ywr5vvZFv4zferJkhi5zWpTYdhJwlDtOG8DI
dgyZK28OfA39dNqtqTChGLZTa5FnvGfYjBFoq1pLaUSXS0XnlIPeWJhpGW2V4TbqCzDN6KScfJbS
ytJF6ZDK7H8dPT9bPIlXCfUw736oIPr99ekJeC4BSZbwrl45ySQTcfjlAv4XcyfeMpViFmFAn0ex
r4CnL1nDFEmkRLuIH45fV2fW9TVCXT3X4sEi+698z0Slu58+Sq55r+z2IyVjU4s9Vq+aVu0YZdUd
uKI9WiOYF5yrI0WtRkZPJPdw6gI5N2LlFE9djSQ5HWQTp1gww5kT4GnLHKM7f4/8xp+l1+TjAkAq
jhieonodos3nQwYX4zhJwQbaIjn5EKOQYZ3+A5eqFc9aUkpgZDYdUvLO+zSlnniXtSKmAwBQREvp
uwjVDuWeLjujFQj5lV0GrTdM8kv0fMVrqPuv3fcyCvqtlo79caJlRSByoAOPNo9lpYdHo639WgJu
n5qtqpn4wtjt7GnEK/LDoMgRoAFka9f3vbQCFU8qvHcJ6EL17fKPhYNTmFtDffN0PHNdTOXopAtS
+p0+AC747owAd00XLemHdGFUZ9zTZKjYPVzUlq+GDLeomIhurp1JjitsR9VwAgehlrJEWp/Bf4J8
LG+ZOCxBMDOnnHaOsp12gqcpdqnjxlJyM+0wpMFCyVVKScxK0yCkGYKXB2pn6WzgDK1mTT7O+bDQ
PT7wZ7D2Nsum2PFUmAS7pPUOlJBBdVMiWkdRY4rOM6UcmIdzXJK+sofHwaYv5hq6w4hJVKMOyTXs
t+v6lCRt0SujmA4F6DmGLPavqgQxz4Lxj3LVNtSudTJ86zotx3VPURty0fdPiYXhn+YEF4nkEkxE
xP1eMJHE5Lripjfm9KPuEJLkOJU2Edtu9UwRieNB3rRqiOXFERHR5aK/TXMWPG3CCUjFaqaJ1GQJ
6JRziTDPu/U/BRDPk9yqwKQpp9A9GiAxCebtE3nyhM+6l8yvBpnizMvS1Yd+3txA/lU+Im0czLbH
E06IDIIdX+nsWmjqBCIpZ2GpqgqcOGRJUMSIXhAunC3ipzxUZMD9K/adJm2Mn8D1rEoL/g4eoVh9
lM5U31ZA74hHCmLlLTH4M+HGTQB5A4c+p9E8173WObLGXuU5dgTcRPvl+oJ2Ahl/wmdNaxwDVpHc
enHKbjDu4pqxG44/YJ+DPVjsEK7coQ3w7IHngaHkR+y0OMuUMtBNRH/dh8Jd2G90H7hOQVr9uYnT
vtFW9jLtjNsk4JLQTUYCHddcy0LBsSkWsdpEC9s8u3misqyPx++ETRwZ75lK4HZX/k8EUOohYpG3
T6+3y2Ng3ws3l/VY7dktuKYpnvSLFZEmICedQoKC6l2cUkDXeqN+cATfx/bmR68NAryDxpSYEdS6
RtaIvmDAl+0aFmOop7uovRhfxZJQ/sLq+dTI2e1fPIK9hUan+1CJArfmnymSKV6yYiiquyzduZSQ
7PgW8citAKJ0YRm0JKp4bWTHTPOGTeOH1jxz5NAylvDeJwzWEQDrCkSqGvY8LKh9M5/IcuuawNG5
OVblawtvWUgUvjcJ7+5FAez88YwBY7NRTZwWOkG1dj+RfeoqTfVE5CVzknleLDdEF6bRVVT7aIET
Cxh93byMF9l5ValdwZrIczYUgiTtwON36lyDsOC02oUjH/NAtvgOCUTYP7TjJh5eyse1t7t9jzBC
y4uwo2K3/DqXGwAgwYEs+5FscbV6i3ymoeIfvf41D2NnOFQC6ISNs0nhIl9tMA9O82qq1x317hde
0th83Zax7W4yaeeu6XyEKH+DHZtWZ0iejs22Mpi6ihdcLFOlX10TFuzW6nCwXzllUG0A/u7M7HaB
AnzqktK3392+DG+Ev3Wm2G76TYIeGabRVMVPNN2jYOvflOBtVq70aIyuCJNbV2ldbpLaKSF+NZRZ
iiqy+PryDRh9QHoLQ4BzelX8A5Uxq5sAf+ZEkPBaxf9LL1zi9VVxapAt4sqPK9p6wYKe67pmtLNU
UCNVJRWSQiuUvWNKMRncXsUHpYZMwilGAVFU8jaC9xvCM+2HQopeB3x0R+51hbh9FzLQCEcn6CIc
giulKjuP6rrZyLkFrUONOF6UQVOE4iQWmNWDfA0Gq0PrioVnIVvM/be3WqtZu1/k0CW7560xbdjT
4LG/N8PJ2VyAA1pub+BjlyUr4m7LFxb+Fi2PAlTngQA6yRSrTQSe6wmZpEva9dU4cBcBtlk5peA2
oi5Fl2iK8SI6Aia+oZ2aWrTLPxnC8ctNbvcwT0zIC2hfHc8ZGfgsqKEf1I3effRZUPcmJsYGPsGt
Y3Jn3b5joKVXMSCOqRCS4msOCehWgNZqVirAphY3GgCtqqYoiSfgjDXAn6ZDb36T77AlCFQPEB5t
gdnhAXnxgne5smEQ+xiB2lGrlPku+B++EsfjPfkPBNC0MSHlBHGTwfUMDPTilyXI++IfalbwLkrp
OK42G5Ev4UWYmVuWC9pup/mDFRrfegWIGxG8BQXVuoEOyM3TjerktP824Lvcn3BNVppQAKxRJ77p
Kzo6qU/F/M2F879Vo7m7fpzWq799S9Im0CqsEs7wfpIOkfOc3KENRmXUAWkfR0YXBtUiHI+BKGSC
2NH+Jr3tPxn6/2jzHJONaKYiDDyjrmB2GmQf1Lzf5HrBhMLYoHaJYYflv+TGqk6RGSvvvxgp/0AL
3amlplqZgDgW3loIxH7Zvzg/6cD91IXnRYXyB1i2SQN9VEufLia2UjCFg8oedZMp4qUoRogjp0A7
msWYz0UYwyMX6Odvp9QnGTTYvFhKCsGmqsOB4YjwHE2J5Bd4duxI1p7z6grWz77N8nI7uaaLSKOd
SzH/Ga+JZPrrdLlYyElXAf+IvhF4Dx2psIlNmK7BA6ncH34DzsqtYLBLm0D5L2QI3kM1mYrLVo+b
Nd+ZBAehjChnK9H7YmVoHBddE1EYfXeJz/KwuRiCpvzQroaUFdYZRy9SMEJg8MCaJNwEFuXztt+y
ShF/qRmw9zwTYLNtjAr7hJViBmUAFHCwXNT+GJtA4Be4ST6gB+W6KYhoh5LLO3pMb12UNTRmCezf
3ACvIJsSbp4xNFmIuvtgvj5yXoRiHXPVKCIzB5eXk9v73qsgjCPBr0ThDrfJrKU72W9seapvrr/7
MRW/j6JGJJPMFiWfsdj+nVGec+LpzAA8tyL5xEq9vOxGhfgxy5vrqph3nk577oPV+XBqLHL2jY3h
iCO0Im6a2kTtRTWUzCrfLNyUFMII23ItaNgJmr0neHJUJiPRIY7qFgaMrAIY16wQK1tjvkqzFKMC
0deoPHSvy7koJa1iJDuXNO+wq6jU14VjRT7pPgVSkAvMHQCFYYOZX1nzyZ5KEQBZ41v7AwnDx3Yr
vqZw8ZtGSaZcMVpoCaZQJRwZYTS2Xx6WgdqrDEjkgJriIY5EZGkvzqNElXpvGfvLXvgvHr8jWKoM
lvF7af8sMcZsDWrFGgQrCuiYDGQbwQIa+3r2gl7KsRkJWZzXkkO5ly5EpLqLfA+tCned+OgiOWdN
8oTpjmIgt6Yi7gAguEdAbAoEdIPdl8+SmfQMvcHyZ5qy+TOF/IOIrsFca2phAl5x+C2sbcmkgNj+
vwUOjQqC2EcNeJxVNryIdsaHWXUtRFKOzwhS8t3dnBIMCSjuTWsKW0qIZbZEyswQuUS49g3NqdJC
6D8yGNmQec56CNivSN4ty5ZdArS+BjxkjjltjdB7dXirnn7WXqlDHisjgFodpwZqM/GGLPMRLKcW
7pEOGrfL2Eh0z9X6EEi+BENmylSAn+/EaookH93cmDQJwjTaL7GXSVpGaX3659g/TX2LPbtX1vcP
onPY8FqNzXXxddO66EsD7n4brWXt0YABRVG2HDcV0sS9TZcXxKp88LPscMJUl8D5I18SsmGWxg9V
BRvRYjP7bNarB7eaazlbefT6oGuhq0kzlmGxHvSCrKaqp+tq1ZJbhMMevBU3AuL/yWv4vkGtJfew
Pm84xJqx4FlmEKyEY64vQziqPYBfQ9kUJWs4723rFhFWhwgl203+Nrlq3yG1VLdT5c07hEZMHdjM
V2J/MnviPDkrHjR5pzx6qT90N4qc9QXSWN1PxpYNq+5bq5Mqjp+68QZ+bM3OFkWFDdBAANWasQuB
dV1zoWXD+ebh40VK/qlWhvK8DaKhmx+bTGNJhJfNU6oUM0D5+iXfPf8qwYL3nfe5OcbCL6DIluGd
dEMgSyE1hbhBxtVTyM7szt4Wuhva9ce8IUl9AQAaYzGfhYQKgMa9GoFU4ktefznoZdhYz9PLVTFm
uHz+M8kMjADubsGF+DSqGw+fwV2U3RI+n0v6A3SlAJpmLl2AzUIdYz9godsC4jjEJO2NRzc3eJH3
6WEsmvAtXP2d5Fw7/HzBE2dcTBlnJD4wo616TCUxTV5GCrHjP8YUwXn7tvBXP5mr/E15F7gRWxK9
bHbQ+H4fr5UjVBxTFf83nq+5UrWii1Puw5vbw5KYSGOkuw9b37P+3UeR23HDAlFg3DwDCHJ+/wt1
GciEYM53qcEEdbF7kbRSK2OkNWxPfPqLp/ed7a6Nq6+NNn5SqSsMjHC75R/kqKQ0FwEEUwwC/Tqn
4rAwRJy6/eRANdvp64T6TM0ycawLv+ZJkPzK0QrzLW9oW8WN2510HbvvE1eQd/oWivV27blaFtay
od+DTnN4rYC3oYbY/ycGBjZYfKz6MfVev+IdFBErwWL88SBDHMKAFbeyiv0P9EVPNcp2NMAbZxZi
mdUWKpSuAJbro75uEipLLGPJF2Kog+i+/MLQxoFme/vv/sLy5zrobE7PWF9b4xzOLy6KngDqp+xK
3WmyjySbqC/Eh9XPM5DIzMQnfZiLHVtpjDjrrBevQrpRLrt4O9lxgTVby2o4E3yhX8E6LYP2V6OE
TmNIUR/RutJ/qRE+AyB688xmPLYXo3t9XnzEFfSFA5RUUYtj5ibsJNmXRJbeoXDHlELtGOfbwVSa
k0QcZPuf3/WjGPEGr6BjuHMjRVkYzQB9H1sLoha0EvBrz5bT7MzTA71MKDmlrZ2C0Oaz885OCNJy
bX5spPhuf/ZX5BR99ePMkD+iDX461QeyuZYaINl6lkwwpEH81TolncYzwGPIswPQEiN1TTDor5UU
zzfBb7Flo9CMaVs821rZYZ95stk7S12eGjJ8SpANKHWtt3u3l3ZO0hfxtZ4tgNJkXkg0OxoaZSl4
n4xSYnnamY5BybHkvQ94McS94B+uwTOzZW50jJ9acEFG6jg2IJOiTr6/kbDGtN3ie7semuNwOa2J
WCex88BPItulf60FyNcYporbQZ20HU7ptL3vytoGMXMWQMnap/1wDGO/qiwiTc4jVNxJOZpnI+C9
XuGmpudT1q9Gow+eT7hIDQZWYGd+QVPatkqGZt0L9cbHpl9tR2AE01vx6YWoBuiEiOBFwyWvrBiv
OkTPxJJnM9Alp0+54BwW0uyI14H7RMGTJCO5VnO6b/tejo4lF+MN8W9AaXixheoMWjTx/RGYFUYu
gX8/PjmQpcaHlGn1Jd5v8i9MkPKQTplAsJsoFjgS2MKnPT1dRxohYWHy3gQ/r1C1TiAe5V/VRlyf
NYkO3BgDAtmq+CnyiYXDYRPHHwQtGX5g8xmyLqrHK378LaNg4RvRT558zAdyCHkrz7FLYYsI1K8t
0J6yzGTxK/C6TaeCcOna2HvBtdCMw8/7oqCGHNVzYdJvrunfIErDjKU0SckaTQ/jCUR+MrilLx7G
uH8EpyN8Czxsbgxby9iD+KZww+alKNs1kLtHB+9UHYI4U+48dr88sVuBDUm+MWqisTiNgbvJ4f5B
k1/JknAuQw1ma3J4yuJcqFlUVxrH3Ts5nk7bANFhMwoHaw2i3WMSOOvEci4A9T8QBfBjiCTwJ+l2
zPZTZ7PZp0t/SlN3u2kEioGmdYxMolSrq5tJs/Y4IiTdW8vxhOzFdB5GqHhWrW87tLX8OKaipQv8
CEwv5TeFPgGslHnSnqQLgeAJ7rpDvMqt/aXaan4+GZvGcHzzxv0xLdZ0l3tncIzaU3/6YUGAD9NO
HNDtqYTeiM1Bkzrv5ukvMWQsxAVCz8PoRS5yoIQY6wFhd5UrTs0a1vHN3n8u7612e1Be9jU9+j0S
zgkOkwbpKIB5Y+cxswN0dgmnEYgchBHmkHALjWB3RIQnE49miDO7nolxu5hi5Rw/Y+SNlIkdHGHc
Imttw41w51l+uLlY4qjSEspbJ/itMivY/gmbkMo1WBbGqhE2DYzuQNk2NkLwxuwruGBtZm6VGXYk
g0DUuEeCE6qoeDOUXw6lMVgRCx4PoDoQkcF2adTMSY0CXPBevFfrIRwPwRZB6LGQmRUPnC15/krG
hWOpSw7fJB+N7wyaeaV3T9uNoGZjG3VdGCAipDhq65itCFFTLx+3tkWzQ40HfECCoVEeg2a63O5J
k0WHRh1BWJ9VneSXtwKNPs3mBXqnW3MQyVnBuEIs+8hSrzzXHehQQ1UY8t2XUla6rp3ICe9kPNjb
l9rTyUFTD/EL1RgSnvse0qANgpnEfg+bxgWXxtjJoIl19qWCWmbmXxzEkq+neH76B3ReFY+xtRdP
Lojr80U7uNLlrJT5OLDTjmDakv2wWqU2sVF5I7Z/ODpauljeR5xT/IQdXZTsKGXtQc4p8aWw9u7B
JWWdMrm9656x6taRhc2BmIVZaR+C83YW1nAyc6E6kWtEJ5T1R6yphZOizf++PzXH2BX4YTzQ53VP
NBizUGu56lFqkWs3amJ/sJY32tbp/RnkoL09W5ofEwFWjLQbfCIQxHoFRq+quT0UKfGcHBcMFs37
Ce+yWUGjgCvkDSiGkn4BB9o4YpQZSnP3mBveG2a97BvN0cgUkCwxlCgVrDzmE/Bkt9qJByAh17WX
7W3izWaUY9CX0BKa2dobS75vfbxeBq0MH2ydx5IAjb8xaa8iRAaYTMiMq7g72w0IKzL2LCDRwfef
FGKx0UWQKUfOPOriG4r12q1SRIBBC+ZPxHaErru56rc21ZmMGKwM3fblJaS3ZI0cLwaVX6bXaLsV
6DkdNPXs0n2uCy5B+sdyq4ioIAVhTluKT4/gZGXfFw3zk+3b6HEs13PW2aSq5Y3mN39R/Nny2f6+
PJ8U6teg+EnqfGn+JvJuIfPaZtZLlrt0S0dZQzViObv/71nY3mlcAH/D+5ThgKuk44IICq/1tkrN
CdlxItVWnDInxgvpESbSJOcawdEN76hkE4SO6mYRaNLDOSyEo6RGnBaCB33ieRXz8FyZbU9A+f6p
798B8lCzREz1zdO8bgLfB/w43UdtY5F0epuOhI+lL3waEaaSCg8k82DqolY+XZPrj/zf7gFLiliP
7wBD+aoqjyPMWC1B6/ZM1BaDyj/CL8BUmH8LfRuNsHjiG4LM7Z3vYjDcEM+JRACXo2WGT0Iiw6Eb
kery9IbjsIwYV7mEoDgokk5F/70uBvovwf76X7ccBKeg6zBYh/4gheD6UeEOPPhfxLfbCOuKw4ZO
o9xUfq7WW63zWZugFvCFgHRLRNhiOJ8UqoJ4FgDHd2MQ3jYWzKcKYq0xkMedy4NiG6agP0xQGuSg
3QPA8p/cDntmnQGmxm46+4l1L7dxMB+qz9DIoG+LQI/6cFSNIY4Sq/vaU2qZGy4YfAFAbJJssHHS
N+c90epwfWE14G4SFJlb/jMZyENcLrv4hREVUG/CrCmGrdXth0oQIjZUs1iFBZLQj3DfpBUjU3sM
p83TxU2346pFCBp3dzGGsRCt5fphzwtsUONM0FNqjPogaJdAsx2Ucc4sAt52Pyv3GlnAL7BXUZT9
DluVSt6z+25J1bhERtUVZUpbMvpbwbbse6FumH8tiU85DSpigLzA1/ky0zNtjILbcJ7hdCBI2XCS
D8QCwMv6LA1DNmZXwCCo/K8O+7lwKCuTtSl79lqCAfge1vtnrl3QdOUCi6pTZ2hHW1Pm0Q/6bntf
cpF2CIxstAt3t1xrj+SPSu9nvcRTx0wJEFaABrHh24XLh8mni89+ResulioBqix9HTe5aNsF4i9D
8X6UaIoZikk2iNyjD8eUheP8jZGW6HxFBdY7Qxceinycy+IOBbQtsL79Jo7Uq8iWAdmOyX6Uf2rn
e+4EwZHXR7rhbdbzcK8u7FnR8D3ZkpGVJz6T7+K6yyBtucj6or2qd/sgllUDQfnlgv0bsN754jGm
fIJMLqC/xB4lAMjOWwKOMUR8BY5LDkNWW9I6HmNyAOJfQOpNDHQ31bTTacjiq2427OZW7qVP+frd
6X+sFtDRndEIj/o9jINJ/78WlWEkOceRD7DO8EeiRkVaBZPoTctPwfUFxWEmmlXDs/WnTRK2W5/Z
yxWdGF4BNHmX5fjp5D4zMmaR2sA6ooAS/UAy8AKRsmlIH0f6ARyZo5Y9CW5H0veGjPYzNbdNHr9P
b4thmxoxzi2Q9N3+PRWY3R+J7Ua0rCMGZ0L3JaH8NjKbpa8CsXoK/ryexepNaKE8YBB6retQWiHf
UHK3LCd06SSVZl5/b5U49lQMTBZGus9KHT33PgtbI6+Wot2bFiGc8iZShURJynCSfWfE4LpYbz5A
1sZasNoMwj5afsfbcajXvtuLAJoOOuw8AkkAkR1vzKuLGp5+OCn9dStMxT1W6Q4bk5SryyGWC1VF
2TL3K/oMJntZVqMnmpr90K1lKtPPjsP4kyD1NXB+WaIdcfcL8WeOyTi13x2HB7u2Zb7QT0i/C5uD
vjqUkdN//uiWL4JPguU7NKHS2xF4L5YoQwhHCZAzxNdCtvt48jSkM2dirxJ3eErjzFK8f4cDiOiN
PT1/hMZakX+M1XG7lATjpJJslOVFXoY1Xv4jY0Sda/9glyUhCsYw9zDWt0pjHgUPZL6vTHZH8pf/
fbIIXbrWIR4W0zvLrg9dyBM0hbSgqis0QHBhnlkTjryvSz9+Bc8kQneTZQppApOlmbECWpSrmSTq
QHiu2lBqSfBQDyCZBOSfDV8Szicyuh3kVP6GG11p+gF1RD3uawrG0PH9aclImCiejIMbWqQSNT6M
kJdP5kCrp3SBnnM6Vxs8jLuuyNKyd82dQs4lcuZLfU93glrG5fpWEzEhHMNyOt+s4ovK2swUTQjE
G6iCXHH3h6Q8raX6R+bBQ+/xdhGXG2cw/YnfrZgSbYa5SGq2N/dyw4qaLgBYULlwtnTgM+yRONRi
sa5qaziLGhN+btJgtoMWFWj6wvzCft1+9a6zCrO2fpEvyNxIPJ2rttY1ibPi5T17d7jMxFVWLhPz
MzQSaA8OrQzhTvei+nOm0nwCDpHFVk50TAYtoXmZnWh8gxSBuQp7GyhtuBoj9a6hE7h6g97bSoKj
TP2Z4sI1CmjSFzvlsEUf5J1G3+fZFEDbgfVF//Ov6Fhb9ORnG8aYUJ1Ha3onvUSMQ8ORgPJXQYGz
8iuuBQuuKa+rioZmzExU6UuqV9R+Orwin5SHJdC35Q0j5suRyfTqns7yjhXbNMwceEXI2U0ndxOH
bXsH3QRkvp4Tl8pEDlvWIt9Zvap4i4RjvFlB2t5dKlA44D7qm+KoraMTJ8+aPcCVUQeknXKKGkeL
cCadp6oc5aoLNIbxwXhEWdy55325NCvTLDiTNKbcFyWwxXaPC6K5Rx+v5t3XApQZ/MwaeHCrZrOu
GLuKPtmIZd8lMqkFvaTcbUWJgEColkOFDESZMtgcDoVZt1UJo0gJvjtS0FUHMSXYHq+B/+yWkwQ5
Qw3RYVa/zCmJlTnbVQUQDAaIADmgFXvDe/Hcx1bfDiqqmfUetA6h+OVvuUdc/cQrOiJaLWTwqMB1
E174LAa11Y9LLNwXZRRifjHijClz7gEGCE6+JvxeTw8jqY9ePvKnCqqaWWtp3HP8i/Nf1/ukDcEJ
mrVKWTJ2jI3Azn/7WyQR6YlmH2DsYaNnQxdEEjwGrAUvvNM8uER48UqPGy9ppwegJXFjOAOpda5/
DW0mQ0EAdPBfQngbVp1m7bpGtrpqiEkwVfKxe421p+IvSrP5Ya6mh2lqCQqmQctCz3Tnc2vXgVKC
TrAdEIeYsBnnWHPPffR3bg4FU9cqd+TpmFn0fGeQGSLfAU4jMmFGLTwDTp/bNOazgXnwa3fBwIv9
Syh/OMljE7OKEZnSuwmZMydgqrHCM4XDRwd4ouad9UnIkI3JEI5qiLZQ9MC51ASAxAMHhC2sCfDj
/possiwGMX0NofhBGKh/UpW/O+DyG7iwe2DO5a7m0lLlplLiS5NbNiUwdZ7rkvg63jYug83W7PQZ
59geQvOM/eMcrJZrnKe378npeT9K9qkCk6AREgswL/moZrJ5sx/lUbZZpy1a5oSsORnCgqHjcV5d
f9lZhOmu3vVbNlm/bir65mjVIdKGOxfktQmEBY3w5dNNj05MR6jz5DorfuskZcXA9Nzn4j8TevPJ
F7znOD6y5CaazUNoYgoHDn5aoHb3f6HyRQk2Dwte5l+/05XCGZrpAgsZGgxsge3k2fQNfvltsUOQ
+s2WO1j2N0Bx9idqMb10YHOIxLnzagtZfaGKGEZw6s6AmkQaiXslDZO8kSg97z4kpUc6h4K89Wai
ll+x2Vs+iT7kayfVGMJxxPchmuANosVjwqmAw0VBnPjXaOgJ5kK1AujgiFTL+R+5gK9ab3aFLrW1
QVTxiU2GWKkS+h6nARrIobdYS1/LC8tUacKSJxbH39T53YELipdBRgu3OrGcrxv4ALORGTHUX8kp
CSbxRKT1V4EMRVJ0BELe4OUFNHKKQv27xOA7wAkeR/Akk3jMeIWVRn2BJciaibnUdTscYgcQyCkF
mqY3z6vZjmo5GgbWVfKOn7DB+KU8VMKIg/uXTRLsojSGNJBUCz1RBelJh62X0Z4qjTzIAxwjyoQP
gsoGUCBvydQ3Z3j6NgUuZfl6L6PicPaqR1ZuplLb0l0QEzXxiSYbzpqJ0MzD71ZYO4DqP+ls41xQ
/cTUVUtDqPSFolCbDEvr1OIucPOPgEz5AijAc9t0abCu/O2Ese4s1GF/zZW2ewQUzBcJ/umkR0YH
srPEbEiLYYxMJzLhL9/sFyr9Bc3qY71BHIfHeyvgXbs0c9IuEhA12wy47OrfRHNgEt3RKZthnXKf
KhXyW/TuymiEHEjl3s8U90sbW+kjF9EwUGqZpU5Yx1uKN4Bk1mRYruCkPkAz1D5CLnZVzLLDq6oj
Y3HdwN8bxdNNSTcVal4se4ayL65hDu8F5VoYoc8LrFnrMdeIZVbLt/m75I5LX89GZA3S/Mu82ToR
mCJ8/V5Tq1nRZJzY/i+8Vx19igJ9vR6NBDoPbriSuKhD9/hdShTb9pqtRR/9KTGxc5ybLjwZF1En
YYLBgNcXg7NRWKwIrq3uzzQQDplyLv3E91A9toXzyxAWTIdR5wmYFiIBrnPcDjslZYmlr03iUOTI
+EtyXv+AQ39T01vpNtcAOfnsXF65Y8VdSd2Gy4DT9u6xYruRtZkQJKBm5PTgX1tgpE3/P4csBPOi
zIJIOMC+swFEgMZ8orbxw99e8puwhLQD6VUGEPAZTLtb7Ef7Fye9twWyMQx0NmO2SFscpGfiCVlw
cs2ZVQHO1/pyJEyzKHa1XjOx/3TZvifQC4+1MSM/zGiqO044b8KrVOgvufXHs0VkborsB8SldXhs
Sc+c9L1wpteM06EeXTLzq/Mp8Bk2xmFY3lTrRe9hl8i+DKdANsDlL+pdF32GUVa/OmsZ8GBdlGxl
VW6PrIuAedXRkZqBYGzYZ2DXRvbjApuLp2izAzC6B0YX5Sz+sru+khm+q/PUT7Mqh+e1sW9bGaMK
sgAI81pbGxrzWrrN6ZEqU70G5d2eimb2uuD2lniiazbTJCrLYIGOYIVzseEAJ9IUnIwcCJ7CtnUs
hzSLlFFC/QO5zEG1mPsDrwUhf0B0D4IRhWIbg7jz3GMf25BqEYZ/Lwe4zQxOTKRB4ICMDmZD6qnD
cL0C1d5SMUgLkYgp3+CQV8ECJvQX59f7n+x8GWERJ6pePOM2hGA0/Qp8Lhn8Spg0alRwI3NHmbpN
oM3eMHAsRS/i6Ii5XeGO5IQbDBgvJdOqAHx3Ly0fn46v30ZhfvVdg+a3P4oANtZv5oEAtQIRSuy4
sFRudCY06y4LCLpT5Ym+8Nha3xpDYgWh6YJi/lsfM40YfFc5gPK+W/gItS18oA3bLh+pZ0wPhJh1
HCpHWQITvOt5XQ/UBEfBQ6AmBwopxSXe0m+eyT55xM+aqWKrrFXy8nDglVeDbQASOZPcDZ1V8xSM
d+rGUb/w6d+CLn0BIFVSjGZiCbLM9UcYZ3lIFAwe8kVoWZQvxChq86ctZ6Uw/KGDpEMRe4hPhfQD
be0jNdoKQ6dk5m49IguVm1sL6jBQlIKhgtSBTDYYD72GAVdppTeWCkE54xeJF4NJcjBusunJAz/G
3+T8cnNj5d2vcPkmOGsIJln7Csm3RcPXUAt8HYdabaCCXha+JmYoxyJ52ZeUtNAcD2JSVYi4QnVK
Tnf733UrL0+4ltKYWrR6CQsSfonPZHwzdHrf8/9XIclPb4UBzPrXWMPnMkRoLqHwZfxahuTGDoaa
wa5oR7ktHj3S8Z84uDs6QBLN6Eimr6fhwk7xUquDil1ukWTe4RJiuN9Hi4BoWsHfzU4uZpdh6FTu
REZwOUW9O0sHJU1+JDIa/Ygsf/FWhOMmZVeVUGDNBZU/QxRlsxVblDw/eUL/ZMXeB3qXMDylXmXM
w5C2lCu4GMrnAV3k9gGdzYf9tipM74shn/c1tk1XvFDpqbhZXZ2TKHYAtwcsYAIHqIiesjxB87cl
DoZYfGXs61qLAHuWvTNpOTWW+o58ntZtMXauk2hK4rcG+4goZh7RxFkcDzbLf1aBru+HPRaN9EfB
tkJ7lbmT84v0qzWUgcJYMsOFwLgWXgrzT/kZ+/wzJmWTxEsYm/hpKcoQarmw28H18VlfLgR5DOr5
dffq3q1MHntX40/SK8jXZQKoj8L90SJIbYiqHBvjAGPy9RUC96Sd9POpU5bjoB0YCDDiIdC5X1+1
lHyeDoXqmiwjSUFvMzBlTcQ9hs+KCR/KuKSi833fUdFWstcEvMoBCSIHthJA1SM/7Q/MQRu5K3eL
Yay67QXEX/UCYkH31X2NCJh0obwrmJLhMyUIz3mnVVE0kaZv9RaCoMzZwzNGYhHiv3sxdS8kIUFY
4vy0095wXkmyXQuWYQxWhVOnHRmhv9F37Cjhv7rgWtP802sR3WQitQOSOWyUQDPY5juemhboyjsZ
sUXBCyLL2AqbGMcltPalTQSFm+3OTmJt1XE+lqBIJoi30lkIpnEkp259ap5hbxcNHxtxNHrcezFE
/uQOigXfSWhyfXS7rmKp4rEtuApmvfpDxmBP/SmZ7q3RgdIpolNdI0PpE84ZLK8MtVIKVMs3QsZR
IUxJUz/+lDuPPDWUlkJ0j7TaW3M5/2m4D4ZXLDoSKhnPxYnPSH8fk/pN2Pnd1Hu74xrl1GK/zC3w
WIiaDXuVFF7ziIPl3T6+gYwnagOP469X5hyJY2FpxfcT7SoFj+6cMNU1hY30hOvXcyA6/rPiBuYt
ohw2oONJ+BVHB1Br8o+pzLrTgwdAnFETEmH7R2clv9jmWmcPeOcAOfLn0GEyVNBkc4HmW0rb4XZ5
B2E9T1VO+uhN4fs9h2sw+2QF/vijjXwRYJUNbAiDGpaoR0fz/5hf8gyVZRnoGi3gznPvXBuAVrtb
krlEaX0ozZ84DUxf1Y/ApZl6T6AOsyGLB2owZodcKMaknsBMFhWVWFJsq5SizGqVf/20KWd7vQ6+
PZTlizd8cGynvrjBXIl6GN5ZH277QOi5lJWuVaA2H4+ByEJLK25gSDM/VJZ0cFoVXm1zBkGcwpBj
x6ylMSXG1gGcbI7leDndrJ2aYqGTSwngL+1iJ8wvShdTEfKxOGfiSHbdSEbhHtjOMHlTlkeL+Cwt
bD8sHFXcYTcd+ij9n+OpPq1vxw0TzdzbhELkJqiObfJdfdqC7zjxIh0ahEcHJzmZEeZJcN0jJb1o
8o5Z+Ez1d5toLI2+GAM7R8k1VezSD11IATSwSxZjjtkgPaWF6jS3VnInTnjbZni7IWVm7+2+yVQu
XGy3/fSIOAWzpKFKgXTu7MQ+fgUJVFpnR/bIW0P56PUX9vHwHMmWwfIiDLyIk3yTGRQZqGMJ2TlP
Lz+FNtXI/UegIo71+kH2PD++qRXdog4KWYPgVBB+kp2ngvWnYGuAPSFPMb4EHcab5HVaPbz6NvS2
IWZR8a22MHDjFHhMgurls3Z4St+6xqqgMkZQpJz9CxVvU0MfIGcMg5uThdswUb4EMbN2JOxexmRa
OYwhBzK3P7IgU7GrndjPD47twfBaO9v2OqIoIhTJBNZ8yYZ4mwHsd/ikaiN8gEYVXXek4KBX9AA5
HpN+oN66nqF+u3D04K2nQOa1uTXm6fQ7wW+1t8LcXl5qHqDfE3D1BsekRKQiCY2w04pHA3O33HxU
XKmB5gQzFj1LTPGdk4OoFoHcl1HlJgxOy0+MeHesPMSckL2WA7HSO6mvdVa+AUaZrZxnQc/qYhGB
rARq2k1GU8/VqzV4P2F9OSMPkoXQWqvY0GJqCs6aEtkrRfxXezLyyL/Jhs+IFBVQO7HJi66NXT9e
Knw0lJqe8FVTZLUpsxasjGplwVOmSq+sSSMV3L4KtcGIj6eh4tJTmYRjCtrtTQOoYvW8pfiYHMEF
jBwnEbhCO93eDQ7d6sTejK6b3wpmnThBCHU3sIrvrwl8pYQOW3zVFFIW9W0Nxc+a+lbpV3SsrIDD
RqojEPd/x+7a+/GnJ5mmkb6DqdZVD547braZCbtgmCWdzovpODK8uyFFcUW8X8B6jWNtl4W04CgD
2pOkpNZX2zxgGyUD4FgN9PBvqyS7qwDvIB2R8XLC49X5OQxvrxVAPnaEqxoO97iqDTVBBgb6Byz9
3Md+I0wHXreuoNxmiF3ONDmwzxLZ8G6T6m9ihWHElIvSZIHTSEgtQPUrnUra8qtUYnwFgrC9m/1O
YvMm8eNbdCZHkjUN4UOKwEXLXA5OCggbpPDNI/RWDv409X8rOqjM3sN2t3MO+p+sBKSdZvcGzJSR
noRCYRplXU+VSCuZsf9Mc6EPs1rTqilqrZDNnD9XvwSWYlaFJnAPyJRkgt+C7kDF8gp8YRH02wRm
91RjEJT+Brtnf6kORruau3kjr+NbryTjluFgEhj3GBuMN9DAlU/APe+AUj1yjaMDXK9uI2u94jpi
c/Kl0b0AvGx33S0qvGy7Ezu0hApnXp/a+oAQrzUquDZcaN3t+GE4P5j4ejrZ7EsN03ocRRzbJGJ8
GmaZcpmf4x9hR17JpERkgUEelLNAEqtdJjE1BOeDJpv/Kx/Zgt07Dg9d8ib7ijPvN4YTrukv6BRm
AqxmnWf/vs7i3rc1ytFh3J/HSjfibdm0Ku9FGddq0ANGuqzE736cLDitsuc8vo34dtvxUDdE99v8
OBGbq6ZfGQqLnS2fzK2y2hl97CeXCYCcMCcijvU/lSVyOB/PfxMCjzJTe+VetZast6uMVcmsavut
keNPmF6dsW+dDVbzVL04/xNx2tWGKJ98E13IuXVbJ5IkU19tr0orlmcqEKNB1IhVc/W+18bq7hjm
Wf0peysIv2rjAQf5MZ73KZ0gBgw0PWH04GtwFdFismuelcJdPrAEItYDnvRswNCTQa4BLtRjTTL/
V2ixn3SwDiQmJ/XuUYsJ6wFD/8F/70wzKUl5xKOUm3zCyvn85p2dlcVnOpil76Gyl6urpO/hw9Uv
ebdhxqvGbhW3j9NpQ6oLErEdeNlqZ/eI3D6BR+v2SkQpTBsQ0a3usfmP1qi7gkvl1bILWpIocAJm
A4W24xBkiKF9gh9OL8L2HhwkzeSGaYPhCSQ+l7bAZ1YflSbrFNt5l9kSN02vd21pQaBEapOOOknY
Ca2ooBzhnyQ89Gxv78YwYYKW4mJ2LD5aNA07SYM+moeP/OLmufgCaSmd6iEmgzo9axWl27g4yI8w
hjhBqUz5BFVzxvkPHDQrFo6cK7Ek0Zs4ItqOt14Supz5zMMTLezSZ6h7WJD18MeVfs00pl8Q0Pvz
dhjuUVEqQ/x9fWQX5qPmlQokfLJJ9TSrPnIgWTDn8QkQjawDJ4wN6gjANmPc2O9Sel2h5ZIWbFFN
GQgGKnaOT7FSS5r0Zb97wsUHsmqgqLTKHSATF6ozmWc8bE3wn5Nzy5RtlxphjWpu/ij0N+FkvaLF
6aF7nuDV7juERvoxtcS2QQesq4gfHrkeVbaTvaH6bjFEVnIBcAY25IjQSt3VO5Wk5ilPsTdD0/fn
Mu/dATNO0oBXOQROomwjLmEIKUiTKUA1TrJfXhrvukCATHXrQdPk5Stij7GeGv/Rq6TxpYTM+4vE
dJ0WWmZzzlNzXFBogUG1m6T1LmfVgy9h20u4BOOD9+jTciR7hzUUAIVKhOBLJgXW5uhTLSVra1Mi
qXmKSxxOc749rlUvmmN9Lf10u04PVnjGuFYz/P7iTW9JjWS3zifRv4V5goDnQ4uCJhqt66z9DI0J
LKQCVMYaL7spcpPDcM+adeiEXGQVWWv/5JyH8fU/5UFpv/QgdXZL0JhKwCBfex9viamlv9dZa2kc
DtEO3QKc4F7W9p10W8na9YTHaVGTc6nQwCWo/1Ia6Oo0m+GybDDcLRow0kq0Auxf0rvV8KbczBjC
igHrdaa17U2iHT55urcavngwITcOdKQSzlIw7tHHDEQoqHse4hOUCD7gwnwDaCsDg7WyCxbHU1bP
Sy3rxfqXsZ72dCZveaP9R2oVX93K7TcnzCaDR/iVSw/DWO+VT+ihvDv9s1wAJq9YeCc4XrpIphdR
YSVx17k4TIKTLwb79N/6i5t9jCSxIqpfxWuhTE5RU0zAsjwjJf4ce4Ghrt5p82MyVVt5x8wo6x7h
BZbSpKvwf9mpKnt/IlfgFITwe+ogOz1Jc56FoMH/8Hun98t0SLSv/XTFsQ9i1yew6pnFOYxTa80h
eEG+MWkuVtoDXcSwVwiZHbUyMU5VeCvB9ihsd+pqFqgfxc8zN0O84JfHnumV7wmomyCy2DO8hQc3
7G7l79//TnnJD44+hC9doFBicxR5pplD2RSXhTkCh/NyTBtjI3LAimM+Y0PHbzRqK7emNAiX2qEp
bRZKVnB+ehEZxkfL6wQDja9EL9npPgpGJ2nkttQ8jWnqcUJD3UrjMhmU9HRCwmliZef3t68ceck8
B5eZfdyd1e9dNg4R2D/MuNnouCyNb+LNc71fRxi6AGjuKvr/FDIuW8csJW/GEMnkYSuuRP3Q/9vV
gT1F6ZXUiDlL2tJ0MZaKFKhDQV8FO4GiLEX2FlbmT+nms5RCMDBD9NmB/dJZcZAwodkIsq8iBqtF
9lJeFN8q7a7OtwHZNYCDlllF8/05QIEXeEiUMFQaHo35vIv3pjojmWYUSvKj4hRCIEWk7CkLzfKh
CFdRZ3IJmaKna3z2V1HV7Tee6lIIR7H572K0k7WOfUSizbPyy1eu3VHQzOFgVqFMmaY8N/hWwKP4
Z/21LuFiq6lB1GCedQ1Ol/2UtxbZboE3lkLtoL9seuoAeIiqMoSjDMAN0oS8KPq4iIaojXWd62jh
qZ2ppefD9oOiS8rjJDaosHEZBn8zcN4l9w2ttqcvlTFxeVFh5G/pNQ7++q5E2wHrGKV0ZDqjGBHc
SyD8g2wSuIl1mZ1bm3Xq28weExTVZpQUjEhIsWZk87yLtwES4wx+c7i3C6iGF7+c0qyLHKWqYiOC
VkVb01gLE6QIRQ3w6JHAplm7/3Fb7u7I1IwFjCV62XwDFCOOSjPHCdTTmvjA/NwsSw0bJipxelkJ
ymys8b/WBIVI2elhos3NOH6mHfHQ1aB5SDusLvj7ppmVo5faFpHHfKWAmj/72ICStcFQFSLqYuQf
K6OpIqV8eqb2EeRcnmAvEdsaFeBqMU2g03kPvih9Pr1GqhmU3P79anXWJyN0cgLTQad+wn/8RCXM
NlrTU0iKH5oSHd+TcfvqidqvzZ5OtUXN7vbtE1iv/mJ6J6EgXr784tkQVDUiyU2fwYmobGon9zoJ
D+y2KzP5lfCHYgMfZYmCkSaYJyCIQkJ2i2zqFBXe4ylvamXp3WK3txsrZwRbUzeJ+daRAJzByhq/
mogsa6b8VVpmvx1goG519KaKSw7bgWMTjsmuyX/mJ2fC48xI+gR1ckLPZjU9UsfWi9GOgBrZ4PHR
eEO9vvzF7Bil/GAlo2dOMYD0CdoCVblYKwL77fhCaL3KyNv8I/4p8G5cXDRv+t7stRHWWy0ATMA2
ZRw0uH0arhXSw172qc+UXfT8GYXbzaaNxrXHnVVLHnJ4PDzQMjXPy94ADlLMrQwBUI5dJ5dZcybl
1O9GR+WqV3qoancNNvUc240H7Zpp0uG4nBfMVFHVJn0faVyzXlFLXEU6zV8gT/8j8Ka9jfKYqkOD
S/myMR5ZS8zElwTTgvz2gAXjRL0YdJRL/AOpmfABq31l2rOqEYYsGxJ0lTu9wQqEjBhz3llfRchj
5YJ9RZlSm92BSGKEk85QdNjwUJfJvHHiNEn0JvjW4wEBjBavqH7k9/noU0HWEBeMbI/4ZpYOq09X
j7Ht0uz1tXbod7SMVjbnBEi5pHDPPvbAtm6N500khE/M3W1hfI25lJw70Rl3Xiiflq0GhgSyibHd
wONfuZGvwWn9kvB8xCZGNTdPf3ytoLgCaojQXsaap8i3LoGLs2GAfeoEvoKpEHFcDeBAq5zjU9x1
8B5Z5eRht2GK7JiUxj8RVBveNHU+CFUBibjHrCdOCzyS/GExiy0iAudLATJIBFpDZkyA/6+NYlHv
1y4uoSDjiROmycTbW2c1AFDJrW5/v81Rjvxd3jbH4bmY7+XRUeJgAwbE1IbIeDSbshNzfrjVg9ah
sQTrX12VHDx49NMO0vEXG9U1G0RkmjETEjT2Ci3v8I+1fxjujH0DQS6C3rqJOe4UavncUZjOzVGi
3mm7mgblVOrM2UvVEljm6hN0AgJXAGzFhJmiY59CY1R1C85S4GJKhrpzNbF91OoC7IzdEK48X7Bu
2h5jClEyyZ2kB45te58xfLiGC41HTKYuhAGlaua23izSeSu6FTixNaUxgijpeV9CRBf6ZlM6rxMk
Revz71nsvgfaFjc54b48xDO8iFv4EYIZLvqTRQ8g2htV/fMaXpuQHRAqk6X/D2OVxh2ToN9ncJ9H
8EL2T+ceb+Qay3lVysbtgEdbWQ+7REbMIiZrShpqpP6s0Q7VJApq9kwgp5YROz5ZcREGCighyecb
1LFT4n6bwO+c2I2AVkyI1fKWP3DOszpLyTPWfaoyuzHRDADOXpMaSX9fcO6PTJouyyxlFo1pZA+W
EBwf+z73Fiennr7+2UnOHy1loiPwXj5pNqY+RNoA2ZAn2gI6PdfcDC/5Dc4npADFI86SbmMlG0x7
0cVA7uqmPYtaHtkCu5at9FjEBT7JjdI+gIBdVV7ngqN9HWYobjkjV49J5QPyYqU4d7Z5ATVrVevA
y/Q7kvgZLPx3TX9ZRc7qQwU4B8wyNTX39k83BRl8Vgq3sZup/39zTPrHHOhERd6Y++kMWrILbxld
ZtPp9BjUVtQ3iBO8HKREA6esTPDJXPwWLJmSIR/2Ye8UlQofPgySHNexF4ME2AeaXQnvs8UCIz0O
gp4dvcbxZOa//EBKnP2dHO685rTtEF4PPvzHcC/VljJNf/LfxNCaHTtNuoVs7V/cRGd8wD2PdDGa
XOi0bfFEDw5jbcdHUiMWr+yUh7UAkHL9Ylk+CY5FVW79B3PKAv2fffXNcpeorsL5IKHb5QZHeaqP
17laVglufQ1A91ZUYh2jKGnVIdbbUQflB3TOoaVinCdgooDH0JFMzGVuxPweawh3cGsMORycZXNw
7l/DV8jKfTFlS5BeWL+dsJ/qbaqel5vDHvfS9EtIIh/eDwzf3XV7Uce8Mhj1rCOgIxENCNcmar+9
shIbrgal+qzAjrGR0jgY3yKWMcexhmqoURxpqxTwDbDFMSjuO2l+7oSQdR7PiYxWgpFVve6tVT9z
fScB43Dm+kbpdCQOAVSAKUhbdGJwyX0wSe0hb/KBgrpHeVv4kpCfUXfJs3m1FKmfzFK0e5tbYwrg
kuhShLaxYwWYyl//bd4GR383dg7BsKKsh2h2Xb3gtt7aye44GaKjRpBsNgKrnYqSnOw0iO+Qi51H
UbFjn2PCJRemSwmuG3DADGgzjvO3lbAgL3niZc2iO5C6aAk7lXIlXJokscE0E+rIJuuyBHS74VaU
JTB/6MO6ZqnV9VIFNLGLhpI/n/4sD6j4dNUWZJnoPVLoL9SfLgwIPehHLCGroIzK21ADa78yYA6y
/tpX6iUKt8nypCRfAABaUWrfTNzceEBOnHKqg8yWr5wQAqEMNBwHWOc0U5mDkXzqaZbWY6cJvVFh
Msk9YAzrQOhEudwYAANPcyHvQNBkTNPb3ue0ujiStAYYO5BDdqkyBs7Oq+YvRkVSHWx7IlqeFaVl
P8S3ftXpfKHbkCjNUdq0rG9dqHQZDQp5LIuSxbV9OPAz4CMOjNzofDo512MKijWbvwd3GlEnHfBG
jxZwtA3O1cyz3fhUf/aHotPXDMwg3BK3oePQ7pGjTo4ZbTCv9ZirjO87O50b3pRIgCnQ6QQ8es3p
LWkQQLBcNGExkMkdShqDgz36PeYZtf6oz5Fvbh15QQXGSk+YDtHL02wNUQ7ZG4RJbTvCL/qfWWc9
l7z4o9AnoylObOF31OL4s6micpfNxeJUYUQ54wgzDbC/ukaLxRse+Bl/8pfmAnnlXe4CQwtZXyDY
Hpfv+esM1JUdTgVAUqR6T3Y3xAYk26wMguOjk/4vl9dfRVK+cLX14SNf0JvAuxG1cHuLDKggAeWv
iOc1HHztiAu9z3/AvulmEJ+TjD2dbymEs3mJQ4wPZegpPl9tLowl2JuSdIiJoNZFnDo0MD+JoSL0
L4CwfQgGwtgSvnJhkk2odEnRC843kLJW4CMO6ZtM0rfoVv1hhoizcR0D+qdzBjmT2iynfsf2Z1pY
AoB16taucXgRZKRS9o35d3JJcDhjs1zz7ZMZbcuU/NXKCRmfmN9w0FIZMdsffuFFCyi64UZjGKK/
zgv/G4jlv59lmXMloYN8xiuFNxka3y8iGagd7EKa96wat2aSqAOcW14x82cxeGMcqLz2T93kpBsc
2v0gfHhhuquzMPf8/upaO8FVi5G9WoWxjsX2d+mIKOy1N0X40111GtGW6XGU8DyIBYG264Z5WXul
M96cscO4vNBVQ+zbU2vXwkdBlTI1Isyg25pr4RzO7wJtoN9m9U3tc7QKUDeUzrVYxlcUTv+10XTB
PYJNGRJtUAuU9u5AQSFz4Jq6zPpyruUeQpNb94j4iZJbf2pyd+Bj7erdke7OKFvy1xFr3Sv8DcAw
wDKZqitRJnpBFGcqs+ee9eQTRJS7wXNwr2xwbKXWVimcy0KGoGkKdTPduImngURQArpIVAhk292A
qCLmMdir+SQ+OFQJGNuzSValpvPxU4dH2udBI4ExsHA02eSxsYxJVIJs2XixFR2zBnkYaMCbMpP9
xj9iHC62pPhXr4tEgzYj5a9VC3iWdIV/YZUurxt+ybH8pbJ3/VjKi9eA/HVVTGBCQIvROfXVW4U+
2PnISR6r8zAjJGGVX2weTcj4Fsbbx4kyUnm35PNXbTkbtNgZOB/kTi10Ds9sbAkBSUa1fdxA6SeB
XYlouCwOK4gL00vQDdpkUZS88RDfExQFGMQgsw00xKLjPAqwyJcHSSYZy51nm5k0mEUrv8K3aJ67
bOnYyPuagQTkOo5N2zQxW+eJ5wPpRObOwYP8xWOTzj05Lu/ragCXXLx+unQL0sJpV41P7NhSNtdS
9o4gTQog8YNpYTxsGOv6F47tGEbGb9N7ArKCYivalosxvnJOOajVrFMSrJ42gFr1RqNmW6NnZzDy
xxJ0lIRocEe1sCtrrrjQNAanXKJy8FtrSesZtRZZ6PDb/4BPViNpjmJI7JWBGi2Ie1HziQC9QiJ4
lHbxnOcty8wcJnQ/rNhf8UX+oFUaOEhK1mrpEvtS/te/ZGtlgj9PfegHl+R9Ozs0QIbxhod19Yd0
PzpTri9WGI+J9k0LrHawwxQIwQ9zC501XdF6mIrja0o6ixbkTHgIS8kX/pDTXxqcJu0DNarEV5lh
m4SR9TC50EyKHR3cXS85dHM7BGQnai6KuwsqalIE09/fgrGRGWw8WJioJBnSq+T3KJi4WwRRvjPp
v4d7rYkwvUhyZ9sslvOERf35yVHQUHFqTGV3g2DWFA1Os4fYUg1dkKwIoB0sbleY1529tu7hOTka
qQut/Z9XN0s2ebAmuDtPZDfGdIclFe4r7IVfVSZXOO/we5wKZ61gzpBdyy1Ouj5rECsAt748VDMO
hNeXZr2R06HnoKNXnwB8ckQAd5w/b8H/4r67BZKsuP+5ItPgnegngKa8Z9TEAcaLnggXbSvpQG8X
k4hsSa+6InlY9237t235H4Vo5bPuSBtU1MKzmkeAVvnozw7od4L9m6ohozQ2PPc3HSYesz+q1ovY
Mg5csKcb+YVqQhXcLhZE391D/wrjorYJsvkd73kMpGwiixwomqV1bRBiEF2a3xLNN7cTOilvlurh
DyG7rAqNNWesVylq/SPctrJDnVXXBtdqktjn9jqbEguw72T4Eo/uj1gS5JHQ2a5qw74NLGC2SIO/
4eJnLYyrEPvKUPPcCkhlH60bqmCGJcahciVKf2fjxxjCRdf7Dtg8scKjEKpE2iDdxzMCYKW6ttKS
dT3Zh/bB0n6ZY98Hra2yzw2VCXu6rRwWjkjPRH296MYtDgNbqfj0tID4yLqu+DZq96YxEnIKQph4
KYwzk4gLk9aNDNXLqdZDVCwfat5Nl95+zDOqDIGnt/D/y37fjD55AGX5TP6C9b7smlUufpywGHkV
r6Td3X5cwsMBrZPpXs8viw2hkQiiOrcvj5zUVByqtrQ0d3jlmsQaLwOml29L8dKty8DUJRo04iYF
LWlLrT/OQI0yvy/tmjF6zBkbA3/8i/cRytTrcF08V8iXjHx8GmgEu2fF46yClIRjlzqPKlemTpBt
pyTQgW7ocyc/2sI7pOC4mijmin0WhBsMo9IYjxvLjmqzT30LvnsikBpc4/wCOIuKJhfcoVt74ieA
9ogDatHhGa3JcYQNa9PqnUm4CvzXCRZIAyCnthXu3LfQN7v5s1Jt9nbVc/OlwoxvoRiXOeBugfj9
ztVhyX1E2Me8K6BQ7sBvILoBtFlHdOpSIUTwJA5KcWeCFa4jTd2rwlHg0S0WijX/mYReyqUHdlFz
bAaGqgGgxUEF2L7ch1ZD93Z1TyO+cMPkl04gF2axDFu8lP3nKMGLM8pBBkkJ4ThBliWt3wg/u8jM
G9lUbsJoyUBfS7ixG0QJf9KomdryCBBNNba+JQb/LUlpn89ezxsPy3VKxdwxKDKwJzxdjCba0i+t
s7fRSkz4dCK8wtZEzhgzRStkPe1hBejpbQXKFmPXgYlZpE3HmIBbfdp3L0PG4HUuqf0c32NjGDtJ
1jYMEhTE6TgmmD2+Ss1kYiIiTzQCVYExvDwd3KeCQnUSUuv4Xr4zSW3iAVfsgTFgZc7PyU14O/Xw
bzRm29/Tq9dW5gYnO1rGTUf4rNPxlNHgvnrHGGCPuHVUqEYrjn8l5llC33MceVj0pMFby7cLz0Y7
MPA8h2O4G0AalzYC06PjnLiUmZR60gpAsMYJiwo6ftawKTjOQ2IXqIu3F4Fb5vZr2hc0IC7ignlx
tJemmbf0hJc/sjZ7masrYJQLys1kmkZH+xaJWqWBgqZNXlOEYrOV4LiSRvffmmXReFkMiLYIvUj7
YP4GrY6UKXsaa0khubcmIknCizzauh3ICkFuEiFiYotmb8P1CpWtV7/CI+/7BfBrkQBigeRJpJ2j
Y1xbqKx4w0RxaySpifq8aHd1hCNsWwzBnI4vakrKpW41LXWatmdrpcmRV70IbxTcZa7boJJkmnMl
i6L/JTYpanCZKcwWbdupVxupTO6cIVQFmgVYfJI2uwhx8LtRVuHQ6tMP/a6OxFve/6etSZoMoqdi
VGIJ85TFV72+RPvcQKyXf+vDD4e2sAzQuGdAWVq2EpGQfPJ7D68cbm1l1OiFbZlUoZfim8rIfO7v
czlmuSzpsDCxFa3B1c/93ed0I0BI9L8lJH1QhuKRUR3osH6pOJOnL5ltSitxFwuGy6OPiXVjwIek
53B1F807T1Hscx+LoXJP0tdEEKPb5MG5THw7GJEnVsL+fGQ9ZiUC8GUvlTcuy6I+vgtRQMwWrHBG
hUk5OqE8ovmTBWWs7CMO78sTKZMYhGywsgdjUUAYXCvR/gq11DxjCktZmPmMhRWXRPxh4QYUyypv
K2rZbozwESJSi2lU6auBLt57JQDfUyKP+m/l3C6kRq86VOLaidC+wLAXXCnVhXKUaeR0LQelNT9n
GgnO/cxqKx+4ylkokRaIVeKebFk/G+VqKA6hH/5VNUBBWXAOGAJW1YqLrWQ+VPGfTifTcFsQhSPg
SF+WGdMolAIKYlul4fPa/80k0jlwZ1tee2Wg1w0+fCMbw2lVKrfS1ukPhG93sC14wa1D4GxwUN2N
p3N0uZniYVXkTQxGN4FywJZh9xNicp8xrFw72d75Szc5j6LJUOf8F0/gZr8lmpyYBhGlcP2XuVB9
/NccWoUH1lLgsPsE4C1Ssm3MDv/u7H7RJItROqzhI0E8+rximCCa79begtyfyNrC19PWvciaZQEu
oox2G+Fq+vFM8/yIyyUner02kwftZjcH4CSdHCkqsXV4A8zWFgePoF0t3UJ0kpN9yjQFthkzHEwK
KlWJVTBW5tpSWed0hIo7zeDtecTidqf24bakMylFicxHTXv3gIeguXq2Zr0Y3cSorSVBtYoM2Zps
25pDGTo9LERrjonfzfOGDo2Iot1mvp5tBilC6gBHb6/gcc3KOzlQDywvNEIYpoWuZSVFPp887Cyh
Ts/XXVsBPfjpJc1rDJxWbEomYCH/lqMoFvnsb/yVegGV/y6cdixwujb/52HS/xTbcXNmG9P/ySQC
5ZMAl/VVpmMm05Q2WcNU05WoiYjRY77pAcMJ+LEDsSe/DOjYrxvMDfnRzdM5bvgcA5PP2Xkf2Vj4
4s4jvF6X7RRtY//vTWCNkM8rR/of4FUlRccA+QQrQ361A0HxMms7GN67sZh0nM0CdB+1cY19UZVo
Hj2KcIKRThPsluBDMxNJuCIx5K/tTQKv4NOtTLW52fOiqJ7pRtsbpFYxdeiWipMqgAViiTso5uf6
V0cL70h42Ys9dwu+31ZcIeBp5sZHVLiJd5SwtvrduZaqWJtg4d7P5gy3Pr0PjBqOi82QaxjwKTxV
vqnblkoah0llvvM6q7+OCUEUo6n6coyOJx2XQm/Yp9T5eywI8WcmbkmwsBf4GSBl2I0wZGmLPQ1l
SfN2cv3ZdEXO2+5tHbIlF2Ny3IPvpg/sY7xSZg3qUCSzFDEx2/buuK0+sdQZFEpbgUamVDIgjIMz
4fHTCgy3VNCIOKYYbiuFmd4ANMzDGgricM8PkjyMvPZXHeLqOKD/GBl7MZAaB2TXjirE+thA6h7F
BS4hd+lV4fcgtrQNWer3fE1HJ838Gnxyblfue5rUbSAAckNJFb1xy4C2IU9W/wz43/ArF+1PFPkm
RRx3+jGbKyVwZTFyknHpRUDBJCFBHitiRW0SDunEE9K8vCKTIxj64xoRHFbAX8TTxq1U7F+05Yqf
XJjKjs6vaDY6kw+o0jAOCeOOb4jj0Y4Lp6hl7aLABNe23b4XDpeE8FPNLET+Lq6UbiJqVzxgY8x6
jt7qkJ6JmKSz93tq131LcFBpBfmqdIbpsPLeAX5/6HvB7LLdnnX1ASHzFQcEjg3CLeVt2tJvmncg
UxORMOLCxwekcTXEzekdeR8kl38fHATtYvMVIPRzegYfA/M1dmPHA8/CKdL+AsdDTEV2KB6qxAUx
93nhpCyAY7yvHT5S84qyHN5NKYUkFT2zcYDZ/GDYoVbNuMk27kB5yUk4wY0JV03wW/5P2bdOVUj8
4fEhxITBSWzJQdhqo7+RpEyxBl7kU//uIYFw6NQD4wo0gxjhrTGIzR/hsA5dIpf998PCMrtAJ60u
VTuUFrYgBSbvrkDNTESkgBxFMSdB+Sk+LbpH+aov+h/gT8jiG9vGUIuI1tHmVAne/vobINjefMkM
1x5bkiaKLob9ji5AiF8swj7ysU7ad9G55Cl9jMZ7PdH8a9YaQhp/jWnR8t08sb3q2GDH2afoLozp
uZEp4TM08edx07W6rnwVVuENpVjHNssbBnOP++/YVgojViKLjv0nVD8qf4EXzd09fk3CsNKA4UpI
ieSy0gvsHTTJUbA/xRUxHRtm+YjaroFxjYbWRYTj5qpfZK8tzV4AVyjKUsNxaz8RC1EfQx4sgkw3
KlyVk/RhbFeNg9VFsl4bZg+4t27MdL874R6XYEetGx5/Q80hUGQBOZrO4h2oLpfoQLFKrEVXfogD
jg9PEwWHaV0/ssCmIm+uGpXmELkstFCZ68IeHUcksVgT+lkQxYTHMpL8Xigp38QcgKD+XDDtkI16
8UYVEfwLpxHxpGjlj/QSQ9QJ0wj7cvwt/YavtMD/FvnZDW1OZq5FDUmL3A3cPZg+QubH/IqHqn39
1lqkbE1H1NB0b4tGVRZGVG0AIUPuui/TXOfGDQ8fWl5OpQJIkUln90iPhZwYKD3OYzrqtZzVHuh9
bQju7idX5mb1rsJ1jClHrbVm9/2GrKwSCHnsdi4rNSudpzvWiMj5L0f8x5bY/RzqiBF2sMk9dEiB
v7/qEFk/IFl2IGZy4bYYY0wHBZ0k9PUwSpbEI2PIymnLVR8nkZOFp27X5f71R4ueRUEcNa1fhFE4
NHxzVq5sWP1yOB7HX4WcQuXAXJ5WPcMGalSXoSopadA8czUh6vUuXu9LMTz8UOBxjOyZMFVNBQA9
Y1bx32KX8gfKYpUwGKSBGWFJKMCHDwmxpIAZwdWcSo3g7fh3x+Me/WMilCVnTD8CnC2Msbx0vxw8
duPg2QkIGB55I3yLzS8NCVcZiJGHpVa45fG3HMSbUNedhaL6dLTJ2PmJrltUUWVfTZd9S2E1ilJ7
piectHibemXyKSHVwMpUT/ruPISluCt1JwXASgYiPiz4i0RtYbNt/w5TRRMMbO6LribqOSion9n/
UyIAz47SOzie7kCmQSlxHJwj0Pk9CTgJvLGAGW/LznEzoWegaGCGvOA96/DYxmQUAAG9BFxtsGHI
CxZ5BIuReknwMVE5peBRL2AU7urSCOYVph+JvtK6uBP3y5rw08fiUzCw619Avy7cFFnyso/u7Gel
vLTRqK3gr4WUs8GCIcOPBahOBtv0LERCHTL4uRKpxq5MKSWg0WuZ3QC82O9rXyx/t4IDDbxl9Av9
jKO8HycJn/YtzW3KickjcbKmkkg0PD5c7mhEmaFbgFcB9tWoJV2QgMEZHqkp48YoOGZFNp/NRkkl
1bXunbEsRzqHSaUF1ZIZRTV3qNHwCYfgoa1D/AOsi9xNt4W0sXTWsnoCSRZbMWrB3IqJ3MiYuHtf
9kX7UQu78HrahDYQYYbO0I0WlrSerGuszVoghvYvVl3qih4+v+3M5n6mMzXVDplIhUaMxJogVqgg
S4WkUK4j7RuHhPMXj1u4yEW/5mgB5SsWav95LuQW7s8g1ZbiohWIAXrSS89Q6K8h8c6FXk8WHUKN
hhXNxl0kMAHNohjJLiWup/9rmvJosWfw1JWdtrAcBLuIWz9luZnzRYarcaNVdL8zhOpnGMgOgyD2
8VdcYUbub5SBHV8HzANsQr/c3UwVbs6osqpRUCuLwUTgAkwc0apeUSwzT5rhOSdWh51fmG8Yu087
eLbRDCY9xOl1cloMIoZoy+LhtaDgYoehrAeVml3CvXukwa4RyOEgXmlyrWxJMFFnh5ofgP6/lngP
qgfwTsj4u7IcUw8TeIeq/CaBZeeVsm1trKYv4QRn8xoo6PJp9NdEdSc+8z3fxo5WM1z2yUQfnyJV
DjHQS4FDJI7SaxzVn503YN//YGAwO2RD5gi6gV9/J6G2MAKhIhDKmi3dryly5mun50KNmy8/Dng3
ujyIQhbOMLOCcoeCql8nE2Eir/ZRBIKQU/PL5ppf+B8V273GCMpVXvt4dvnMsWlelbpkxp1k70He
wUoRzYepPGw0yCS23egOhtuizj4wpip3VJCKVTee4D9pFswiHPaEruur0bRwraUKYBP8Si13B7sJ
WTlzAv+WbCM1IQdmbnpnXCXIueD6N4sIYRvjt/yT9Lg3xty02pfF6IOBfcNvjkGGLgstjiYYf3am
hb2xq9YDFoPoCoGxu/pCi6uZwZkFiV4ARO7Npo1tss2Iq6TYXl3YsZP8C27oCqP1u0baCk0N36H0
BEXJ9IV6aMDkUMxCAgc9uM9Av6NrFO90+98Z9WggfsKckU5qpZpHX2tazATte4LWuVmmlW7/i10C
XkWtupHi5qeyxtvuzlg4xWWY3pjSoxy4UNeO97vjYVqiKa9rzGGhOLSdl4VA+RT9gFpBoYTDnmkH
6AX5ZMBndQZE9Ja/RQk28CJYfiBWSr68wRW/zBPy/Vb6JtlgT8MfSq4uCPHzhcFDFpSQSTDY2/Zb
xySYOKqWjc2WKP+98quVidJnUZmozu3l0Zz79fiVVn+v6pES+wbbHRyZ7LFDsZCvVsQO+yWx5bRw
HunD008CNfo8RBPg1mEOKqkfBHjiYHl047JXnmK4lEl1Iuo73Xgeky5o0mPmdHMsUWcZ9eo3rOq1
aMsdBMbYQ1bDiguAhEitS5TpkKPE7sq6sRcpTE1u2fF9UxCkyBaQyiGuDzas4LyiXXDLNU2dvg7E
zRU2DwQ5snBpmw6r8SvRd79BNixNWB680IObLonif3Mo4iFqBBCUUa5rIQjBoZ3dy90A/jeFn/qi
haFKxT0vj6jIOSCsETePDTi/zbXRatvPaMXZF9Dt8MS9Tlkv2kvWApsuc/BVywUcrjIgO2M7K8+e
1xIzLm9UQXLwUQRQQmJuMf7mO8X+3ie6LRU5aDwhr6yIos7XjHs3pLXXIShf3B0PjF4fveP9dJFl
4qF2g1eQ0cnZnMqzD5BtLDmQHEDIBf7KLNc/frhyzMnYzF0auiwSoM5eYTpZUHC2rkZ/Ihq2i3V8
RxO7e7ZKiXJ00co92Cx6RtCCoCqRpgvGCmK7o0fV9ad1WAlPSDkUbfygr/H597JfZyo/1YjQu8lw
Jazqo0nq45oq10XxbFUOyDmT8GHJm7NQSxLP2JsyiSB6Fy1MLTfK74lOyyp2R4tFcAvvpsaVHV0/
7/WicX9rJPoXthhQ/moooTgrj6H74XzRNgAnS+ur5ZDTDqQEq6JnfCrqb1EunfjU7nVginw2RMJK
yhlmS79zAJsfxkhx66OOZ3E/qz30aRkdt9iwIBviElIQBPV1qG9JNh2+0HplQpkYjaPjlpITiWqJ
Q+E0KXBAYz+zxD4JmObO7W8/ujBDWe0mfhOdtp+0ccsTD248kx21DzgaI5hJCs84tDxagkSTZwGn
l+z00DM7rhv4fstt1TLQvdo2nMbp93FVOvdFJywhA8/odZFK36D1GXzEsxxbVzvEOAIDyxdrgfGE
8+ah0Y9KQ9pC+3Yf0NeztxHh3K11plX0aEbWzrTP3pinwkFhnVAbOxGXdFEEO+wBjfsF5X+o2uLh
NnnQx2PIkMDObCCjPf/FPwnTdaOFIimVJy88grlNkErszHwbkaQBb+Y3X5Rs9EX/vGo7upMLLhGc
pdGblghXSp8Kd4UGd8TfoymKBXye0UAkDAIL9udmyXl4GhHGP9+H/+TNOpAvIht98bcHHco53mbI
srxEQlVzs5rjUlbTViEk+2bb85bP9AhJB4KBH2UZqCF/nybt4NY3SGb/dFdYVOyjSAXnY1PLy16X
o/bSCGF9jUzQwxkhysq/10MDrSWBUGKyrj3ty8oeGvpJyUwmV6eCJrFlwRVAhDKn70EG2r3ed/NX
nWsPqTfK3c0bF/EaUigOPxHF6i5MlJPuVXZGBGvOkeYu6zKETCWikD69BDhLgL/vLBdCZizOESx5
+RtMWN0V28N8/8bAXCMzAGFxCkonn2bwtfGOJU+cLI4AQY43+KjB4/8LEsG8mfqadb+35sG1spaj
JJjoSoijuLRnW8Byk3oqSkGBTDwv+rnUHoqcuAQARu1BvN1ykI80fAh7hxV0aXANGJ9jONZL2pq/
qZg7dVmOaFgbiIjjUDdPXMYtfH5OFwep3ycIvpTpmQDv4+4kKUF2bHL6tVnTqErMBoPZo8B1qles
pl0u8wiBJ1westFFdFqUbStBK6GdaW/kPEY3g1YnqTKDM6DV5ccOnSj6ybzjYaIlDnPKXQt3DgrC
0wz13mkkOqXzPBNVkG92XTR7JTH3YHY64r6f/OQlizzAnWYUKKk4HwxaG+alFt+mCFnJ95C7apQt
3IK/9JTnaQRkApQqKhodiZ/Kz0RYBlGBtSP0dgwruTfiLHgFryZ8RMa2DNDVm8V39vygji6+3JsO
cyXye3k69UgoDzrU3UAC/WEX+hAX6agJL50tVqbeXuMIrA+aKuQzqQhqnpk74X/DYqbikuB35mCT
sH4TxFcPd0NgvBc1l3vsLr2d7n2dgIuhnwKzeGXhHk8BipLdxQwEnpUrNbDLhkwKuqTNRdXstTrb
u4fIHmCQRcK1CusiLjnUC1x594LAphGFBNzdk31lKmkNBhEYxLG++DQy143fy9l1GWBB7Gk2zXeH
hEt5PFCt/3O2p+dMLByxo/HQi1BvEPKyGcHlhABx1PFyAMRjzNl8kr25+BtNX5ZEVTOD15jQRqrU
vJ61z/b1iV6uV/LZ6rUI672ZNOaVN+d24dZZSiGOy4oPXx2lFrG67XP1ciUAIRIMY0AHMlKUspkW
JanKAPhMBlytr+r3AbbovpTCB2Krpc6xqtTQsZ7IkPAKC2kZqc9EedQQtCUHZ8bJWSI5yBohHnlh
kDbH8vIBadtxfOFJziRiIhOZcGt/wCl+QlOBq5uWY6ET89qwSfas2tj6s/4Y1d48q18MSvzvczqK
U+WJjwQ/rBNLUnl2JFri9+IBl9JS0F2kSMDkNnGIqLa64pUZWL/0iF2iifovou2JBgI2QW46DttY
Nz1ogOyxgeDlUB4j3AAZTmjo1AzLFL4RxfuuWPDq3ODoyMBpeXsItHLtk6SB87h57qA1S3e1zD1S
Zcf/7cEEsIydqM0KHJxMPT3plUTB0xSpCEaiJ/jw0dF263Saf0SdgDCElAUo4uoSH5q7Vscw9MQK
gdWX7uCNT53no30cnm/mTVU4BqzP0DDepBoD578UmvqPgclgzlQnkWT+1mwQZe7TBehQxxilGu7n
GclDEnYuZmRYITVVpu+Pg/55+2+0xUcB6dGa9VQ/UALVerqzAlwzQ3rTXV3hJw87PvpFTsuPT42C
rKwhErBFrRHtabb8uJBmdFIQLCM61mGzokFXihMLyTyecISrt0KFz59yllNzY/eJJsOs8lfUuAAS
qGJWlXdCQkm27QEDvj7WFI4p9ZF8NoiVwdMaZn44rOMKLl4aG1qU3sxzYZmb/FXOG1RtSUYmNzOS
3xS//xF36tMbB8WMAAp/9yxof5bmeU7/5U382+UjzCdLu3a3l+/XbNcGg8uzxuHuflFYwIXRhzc8
skXjxJDX2ftOaZBf00u3KB3qjOLQo2kkzo6NcXRlpnZjTnT9hzQkN18giqR/npLgdmxPCcwoIt4C
C8UWxclARJ35LIDh/VkiXZ7nSW4cX2qPcPTDJUkCZ0lcz4fJtISX69j6fXypGxGjmnJT6zXxT7gV
GOM9A9xTzG+LFlzJjYVkGLk3mDehR8ZjkvDrpQGBHRbe5mdmQUwmWEXJQhAGxRV8iLNfKt8NfTXm
j5Uej9qKDF9u+5IfJgyNWT665r2WcU25zdhevM1WuLZDmeKHoZjcQns+KKXuF46tFQ38q2ywXrBW
pkhmaZOfS3IkdEYr3Gp70Qx7pWmkUd296wxQQbF3awwSo9DJ1APaZhos81rqdeOZrZHGzd2PwQx4
b8wOdiHy3sPVW8WrJN8RWIY1TQb5NQ/5wwCgN+Cd+M05vGsdOds+PQEv/ihDpKhpDmR3AB0fdhz6
EwOhwNVI7+jzL1z7W9FHOV/3AA9Rz5r4wxnY9hVs9PzuvD8NPDttKkdmjuu9c2DjA/BKr+8QJEO+
yjx/InbcdBz4ppyH+fmzZBWab/oc3H6tQVYhZ0HLrE6R3phQo+FMcygKj1Jyf/RyabBrgPPxBfMZ
lOfdxESVHhXCMacbSpHB3SN7E5Lac4f1UW85CPXl1dD1ZXAFJ3tmZCt0pCg6aQYCpFawnZ5qyHYk
M83Sbi+YZg2o6/pbowTUumdZnRbncP8L+H/pjKKdfwcLv+B1z05rfdSgSLpDqK+N7ZO2G6vbS3Zn
vZJnqxRasYcHQilLyRDIAmTk+Hvwju21M8vODMkCIWus7FgX2HZ+lmQ/NW9WWWIRMlKi38DfORyu
RG2RDFySugrfqOIotTKkEnAy1VnP1nNto5G3XKNHm6gVZFP3yDCpbKu5N8U+HSMDgJ4n9tn/Kkan
Y6XQotSkodtZ6XWq+QEGJ995IEgtKlP111QdKQKSULPZojO4w0bpMLD5fJ7JdHd+SFPdzP3Tu4LS
75vu51dpZ4prJYKM7owSkZKwfjFig0iMHzskoWFo2wEX5V5X3hCjwWPES2NViIwTqBIIYIjkT5sp
rASnS1sDjkSnaPAtPXcw6tiGpLmWoUITgrPGnZHbmVEMfHwr4tgQr3yELESvqiLQRSPkkfRmlYQO
V4wNYN6KZQoAn7NR4GWD9B7yyYmdP6jjzMqkdkBxX5lcprb8+oIpx4se/tIX/ezR649CnqND1nbo
Q14SyljEQMQYd6jht79OWR1IkgLdNFS26Tv58MiSEirJDHzU8ksv5KlpLlbpm4rYBLxVv2POEGTO
skkAXMUeypejoJ5EtEkkyR/2SdAgRAC3F2G5/YgsyUt9rjDvoyQ9kY8iVDTDkDLUC5MQ6ZlzbJz0
sGypfoT/nS/3q5upLpNQGTOtS2gJuHrpcWGy5JYWIoUfAQn0RnQtEOgxQPf6lyWj+JuwP0YJwOAt
8WaxIDALVu00Ny6FSBbS7rCoH/KEE6okWp+8eov8yzb04eZqVW6vFPBEU/dYIhiPQ3fav/sZs/pw
lw52fi0vJbDJb5+cOMdE37wRqe4Lw04W/xR4MwBW+XQHLdcyzvU74f3j9ayZAaMQO/8KGG2jNd9n
QCMvv1QJzxd4NFJdpFpSKx5AOdAKgkZsVSF0b3Ntznqfuon8ZexUfroUiryJKVy0vXEfF5ETGm5p
r35SdFfRwYIs8dvanh93ohcB8hPInE/DMrVGQ/SHIQiEhGb9KxuGnnyuxZ88l+eJyKXp0N7KUbWi
Biqo+Gv0EVLiWDjXeCj++sk4k5PKhVB69yFPz8mmqnQaVOSWyptnIoyRdBQA9Hm6Zc4M0GGoUt0K
c+sWD1hnDzImGk1u9u1qxT+NoKYd4hdQ4jVlp4xIi38EfPQDkKqfyfUvNvELtoVvxf8701IYVNb/
qtfvOXQBe2yHrBGslFlTFQoRJCdryBQuy2mbSI/r75eMpwY17zAqWSYvD5S3/WR2C7t1agFpCFZG
ytGlsJAAoUpq2MUQSQeAlPp6c4OyUDGo2WPaHi7zg+h2ZQ+vb4N+Bjd5N4GZ+0lLkjeaodKPnHDQ
6d3zma6gxo+pa/1fC8V8Una2WaydCWjlukMHAFGM6RuZeqdcRgWWKWLSzjghFlzA5Zh2KXjPoZDG
EtTykqmCBgPDQOhcS1BUtnjwNZ8ZWP3R9Op5mOWh4xCFnx3xGTn/ZWq8LCVtvLpUESXTSjLIYxcp
0DvwT5fSc/wtk9u1Awr3X9cvMmBLrLCHDmodySxSZcqbROrjkyRhDMNmj3n67CyAvSNcLsYMoqFs
H9IdN90CirUCl4Ui7jYvFTiuXD/vPyMKSWxmWcaaGhoJfE933TdSWq2hQAEyHdIsaOizj5rZdJNk
qPKX3d3T9aQ6DT3gZzi2RvIrcOyEnMw5OT91MCuyf39Wayc9HoDj+EVNR/oBoFL0eYs/ztJHVzuH
KPnh7bA5ArmM2+4WQnjyMlnBNbdW3FP1xEKxqz9+62LSEWbIpOyjyUEYGcxfvcjRyK/sWgVksow5
yl+ODunuohbi8kyH8ACSQEfHRU4qTC5pBugOv9one8YjrowKtISLmsdn86IS8hpAV2aTyafHic5n
sdeQx4ZIizCZgkq1/Sqp5zN2hRtiHc5m+kN7QL64AOET6CuEP0oAB7/g+l8k3Zjqip2gGP8BX8Tm
lRjkNkveRKxISL6xsKicNaG3uG8yRgNDvfgqr0ISNOEi3LFmG0A57g6BBJbonOSRTAFj3KJMryAn
8zaESsG+PxptqtIsmS2jqQsP87umlVUHkauvKIlusQ767i6Ojk4PAYSQBL3QQZCPbwjGax3WtQbt
mk4e22nTGT35ANMOciKd84sKWBozjD/Mr/8wrYSDN4wdX2ZvNBNA92Vex3JhnxWF/lvjdvmGAPiO
y2LY7mipOl75pYGHfwO7wavD2R6VMzHd2FdwLVweH3Tdu+175rydtX1AaBig2Za3EMoFBTPMz+oR
N3SsdVvP2Gglq1/FPHgt7QGUNho5wZTimWRvOK91oPIqo2IG7ngLutHCXCIkejjaDqHJu/ijHehw
oB7hGy4qxETQhfxzIdt5Rjes9n/R8UnXb93nPhZQzTFmb9hjceMmuVetqtwR+VoRJKcV3B2fBE1R
JA3seSdyrrJK011q2Z+DWbkZRemIRelVwEWtz6Ryrpnl9iK5bLSdHy/a8J0Ifa+hJB4f2KPfcqpF
hsNHnlwTQOSgbgNSl0sguqfQuj3wnGLdP9kA2Qa5Yee1JsZCjIvdydzsKhHTeBGd+fj5mOjkLJW7
FZL2qwSe9H7gwC3sMtjH84zuKr46zropQrKqs0vUNMuZYwClhT3Y+gJb7rk2OfpCGgUZFDaoiNyv
4nj4mwZSiQUe+21urD5uAf/VaAoNYmcPXljywz9g6qBhb3VhrC8uWbJ5ihEfQQFivR1D/3Z+OSrC
WbrVwScxHTOhayQOJgwerTXgY06a3hlx/xrNyltBaa8N9Y9S7esiHV93RfsBHHv5rJ6dUYHQdzeB
YAPrBSMpxLLuhXksEK+ZddneamfVlFj1uzx8dxtqE505+q/798eAC+7jFaYKIL+jOEq+KF58VvYp
sy7AKALPQ9WDMxA+QTVX2aUYiKlxxR3pHgeijUj9d0js7FebbIytczVWn86oaXSsLqXpH+sGHDu0
DYqY1OqLXzxnoyad9X58o96b1jzaCN+/SXjnL5vO+KcelMiBJYxWAfv6CKPqIVB22Eppo17AtF9m
Oy1majw8c7sx6M7XIv9ONYGIgjSGKIwuic3M1pbUSbrBxL6yg0pKuwQpM8zTkf4wF4jAiGhLzlGy
Zk2J0DVFP8PMywdVmZ39d5QfjVBoI4EeSqLDnu+x6kQG8FbGFVMhXAGQ+IWl4jQ3uo4Mi6eZ1y/v
NxYsK1+EmC+vrwdBy2HLbj6CumC0nV5D/FSxinsTPK9vUJr/J75tZbppMG2REucgnklWmis/j6Tq
ZAUseqwh+BEQITzv8ZckiDTTkHD742XES2Ii7DyxbK4MIMW9b2LiPE/rSke1/RdsygKI5T0CEkGk
x8xk78mJZc3tzhE+3GzbljRDc19b0yQHZAGllQTn2qhaTO1dppH8z4N0bBzk9NrntF7TaAcgRxIS
X56QYAHlz1H1W1K8vKn02iwE/HQYk1qjpCTGO1H+w2wx4TeHp4Da7xeormhRo1mUAW1GSi/qBx/V
A2JL1bcAEuX6FBR9AxdxXsVLVxLPbCtv/1kp6yoihucNGgi8DbyoiGy3Nu1FKAoZNxv5HTqwQqAH
ESHIJR0k52pSMB6CZB2q20o1HUY0cgtKFy58fRIi1xzxMCYyWwse24AbNh5NxNs3qkd0CAOmjFGn
9yoRVjXYVy9JTm9X3rdnnlXJHv5gGa8etP4ibHkHMLK6LseNtSyrGKqPnlDcwT3+bq+Upa353gIX
FWL0akySTZIXi6rO6x5VNqAibOo7WzPTlbEkMyd1qAQh3CR6YJi9gzf77uEnhXPiU/Loh+XQWJxA
XzLDVmeo3xn1YOU+In3EfwoAAeHEEFsBwEbs9qAWvTTdOywElMstP6CalQEkK84/II6qCITDoTx0
IgCo6nxVDBzpkx83BL7aIjKPX+e/qBNTkzyLGQlDInZ7XbvAbtmAQmCYUeJH5yCBWVL64DVE7TuW
DW8qe3JKbdoE52P5kXSUWFq8ZjYf7p57ocbLzvcSpoAloY261HTfYZ8XwtrySYJyRM2DTKyT7pHD
29681/7DGa4QBzDviH9TfFlVOmIQlKL7T52m6OZw7lvUz3Dob6QRADByEwqyUhgwCxNq39tdmxdR
knnV0kec77LR9CtQIaPfH1fuS8SXrPRiy07zWTP2pODkc09IDwTfzKcZRyWCx3ppwec9bgDn7ukB
6BRurA8b99HkjAVw8o0mnjuWErznMd1GV+m9zgV/POZcRvvI7odY9T/QN+aeU/E0urAxoUmgqNMA
abRtUiz0R0m5D7cIEDtD4LRvPJ8rSIK7VcjzWZFMAP9WUh1OKBRf5bIdWS56B6qqecoxEyy4j0HX
TUkg1qUXCGzkk4MYM1bHb5XIE+b/6328TucZlBTcL820aWi0hYbHd1IxOTGPVYm5iBRlKfIVslLA
SGMGPmWdMwpmlvT5av0hsNnjW7HGdpXmhZWObXOFfHOQBNFSR4RFgT7rognxWGYwziqsYdvyH5gI
JRGt5QhTkwm+7zWgzYl5LZQjlyAkfCGZm4JYnfnGxozTj3q9USGBlRbDhjhbidfcU+a0BuwPJjA+
BmPpPsjbi0MQN4dB7/q48t/WY/f9TRBeKQGJ9qiY2ET5Du3VFK1oOIh/r2zKEzW1SkIXRnzfwr8S
UZIW+TvAbWo1zvWB0n62XtNH2fklnc0QT88iINgYH3AsOrZq576WNXprBwk7rZ+joTgOA3yiu33u
HPePMab+C920/V7FwL7yharv5Zauu0Itr99q8K9qJq44ZgZi1DexyyOuWk28k54zys0nfBHRHghQ
UcS0E6mcY9a8bu7Ra/a3VhwdGajV83ahcEgXkBsI8E1l2wpeorMYxsY+D8RZkvrKl7y/WH/HAd/r
pFutiVsuUG4xGAFz/vUlM61nQrsWBQe00LtEZOCuIX9Pku2ZQaOdOGYsWuVtjIqRnlqqhmVHm1Gy
voWdCbOcxk7Ph2Af6NZGOykIPQL1PPMMqNaHgS5BgHR1JeX2u1PSzAtd0HMYMumhoujr+U+FTVv5
QUyt4MMRRQk+cQZg3Tm9QQ4p8lGNWzAl1yzjRQAivIITIvap9ff66wG/KIs2QZcaA1ZWr1m3LuY6
L+sTON/h3uyUTuc6B+McszSsC406H6S+iT2S4QelSSFQyBaEY6nwz8Yp2Zd6l0skkXld+BN3f/xd
Vk1nZgkZfhd//CLmqclfE9nhN5awuIGv7AvKNKUhtD3EEDW2HZAEkevrc9Bl+OT8vDMRUhO+QMpz
vGl+WayOtIR8KeYlGYDD2+2bvJWCwOTu9/uqnA/c8M0hwK/y0cdTxt+SqeLy+4nb4wpsMkWGWuvh
GpsDeZFh7Sk9yGKArFShfY+7xj0EH0yPBCfuv7pN6brVJSuOKlazNU+6YBQcKiF13tWwmNv8yYPJ
/MQ+8Oi/vpk7qaIsydzxtrYl3NUEFJk2h4/zb5Lqjqpo2RFRMpfnX/JzrgOJjULqBRRMjFwopXGO
UemErgTPjzNzOgQ6G3HjMXTcm893jPx3dwKX3Bw4zkK/6vSKVknWjHDKnTSCINSlTooq+tXkM17r
0shTCzcjk1RD9BOIyA1eN9xqeXcCKy6DHlLr/4W7Yd24CdKGIaOoWKJqhxVCm3NMkds0UB6ehfDf
Qj3OsjEW2ei+wsIywOTcLIWcEpkQd5CiPXmX368CFZ/m6rHn7OYeV+K8mIVTeinhSgCH0lsKmjYO
cGsrbyPa+V9erAD71h81/orLsIsovNQ+q4pIjkZ0Oo5fGnn3yZIaoI48BeaFsOweKz8rT5WjFx0J
VWTe3sldQ9q2jvJv2d3wMUH+ptqHAABVeSfLoUmQRvLyqbrzyl+X81czEauPjzq/I4rqiI10vYEX
t/GkXXq/cHC4XFiKdD0or9+MOnAurFY9f8gEK9BLRKNMlHnKKvHURCZFepXo3OwFnXWNfRtfesCb
IgQOxQ6sbKtH+5vf19iAIO4K90TG1oG4epVDMov1W9xxvlsh33Ne63MYLUZjU6sWooxII+HzlWbe
ETFrElONuNhoSE7u+cy23yc42j4mFfDPpZgnSF7lDOJj2u51Cx5Aw9yl4pO4TmkRX7grRMGs2You
9aza3lY+bfjRITUGdEnmLOIRFRTKmlyIyVXyo+ZwxIH6zr60SLt+v/Zp+vbM2CR+/OBe9h/Omi9u
YjVFyAsDV/jOEi/cXK7CQemQV/mVxYTt0Go3XuUh14Inwxn6N0syWe7DWN/gvGAw/kOYqyRXcYWm
hUFoC1J2YIq+mCbtAAbCcoLp6JfoV9owAczBTXg69ulvfVuZsPp7aXucpj7mx8REB6ylj2nT3To8
W2JdKIGHfkp9YIrWnPgfsRVvHzotj5DiAy/yzCV0EkMSvnKjTPJI15PWzZ3jFLc+Zgpuvhdvb1AU
SFF0Y7PAfKFjk4u+u/9LL/0Bt7ftV4Qk/t7I+uUa+bOJ0ytUyucPpRC9CTo1XNn84XtzcR2kUEb6
K+5ZoINOVIxLY2UMhsrlnw2AmSGayHvksh2rUKmwuiZiTN5Mve3+CCa5S1IrVSSdK6Vp83Rls3aE
37VC/M/egL/hhh72Yk2FgRHHGyZ5ciYsS9qeJwfFzxje9SzEm9N6+k3TC/r85ClN9qAa8mU89Y8+
e4IYCGC2PY014nSavHXSM0JuRWQnv2uL8jhBxN8lhYmaQA8IFqo3YwYZcZ/FNMiMIhG/9DPL54P0
Ad8oc4Tn53TQwdX9Jc1IQuqteo3tJiigV+cWmIOAHmcCW4YlE2D2/Nbkb9UpFm5o3jedx5FV5dNP
4QDaf1QhcxMawxpIzcJ7Yx3FvS3iEJ62dGypZ5Xpdbr0Hg9BqtSQwVYNG/ajlQNR/BzKcf2MIDO3
sNNKrRaW/2cpZdUV7s9VC946xhbPCPznopjMAPpoDjGckidUpBgWS/ueh0vXZk9JA2Behtr7xxIi
6eA+FuZY77szRw0cgWl5NlTPmQw8VSzvsAAc1V3RbNlfZ/p4s8KLUV0cY2+/5RtV7bdbVVJSlfN/
VYhXz+BEP9UY96okSRPBMOB13Qq84ySqPSk3favW72OWny/loeWRVZyi8x9NQHnO/3s7DDceFzrr
R+thX3xXZT3bRkHXtj3rFUU5LeKlbJsi+seqR59gCTa9/lj1O07y0SwRYFS4z48CPfp8oBw+d+lV
RPeu5Is8g0/EV7QtayJef7/Tifn0xb5RMsuyIhZ6FkWtZbvyayS2kzN+TbFCyhkd2Jx/98UIGjlL
V0cz7NGhhiYxOpdrRcEwX1DfqrwcVku867OohpHwjAG5tLToJqxrEYW0dk57yZzyYwIq1xCsSfL0
iDEeU6GlOnAvDPUwfZpLHRXgXLKgFSqE5dLQSLgmtiabJGb3ny+cEX8Hyi/XQXQXraeDDT6fZc90
wj59R8G7Y6WLy3F59zzCZ2JD4YjFQxb8hmm/vWM+7lyVFk77uFHafO++IsZafDSbLvEYRCUU1N60
Ms6z09ZKJ3Gqxpjmv6FR7vXGV/zzHdPhScQOtx6C/XnT2rcf11CDERoiBnl0f2RzJcDRWo2iFnkW
e8/RMAeNa34tGJoJmTPD5I2SzglcCGAcQmHatz9zBiEeUCub7lYKqV/QRsE5Y/38S8xShzXkt6g3
kQPdSKVk4CSE1OxlQ5lDkRnj7ce7b6vMtmMONm3VIcK/RUOQSPpzusNUGJlPKBPusaiJmTO9G6Zd
mWaeQxVlFPnGRkvdNLG7+j+35mFzVuvsA/GnzeGWZDVHc5RLJyow6gxhZIDVtidH42g/NnLGIjuC
shoj6a5vuP4S/mC0pWgrdxfSkO/QxzdxXU9L78nvxLoMvLk6xn0cb8yupMGO2OKE1dCWzZK+slTc
q0OM4ILoWF7YAmeFAY234tW2LJVnB/kJVImFiAZyF0mbFhTsTArvbHz+QTyE+t2E8rFXOTwQO1YS
dOwmpAMbXK3HDtTQ7QhSC5EOnEorTnkkaGaN7hXiyOKuizh06bOlJ781W+EARxjKnibnPzLikdc6
fOSBnxZC+PrNd0/pfUn2K1xOPjDZsPsD+YBm7fhkXdyLFfFwfLnQtWYv9/85FAXBvVA9uBwZTYeS
NevSXVHUMCTSUPyaO1SEZgyLkUcCWO7ppzLMDZvZmB4TrJuHQ0H1sOsdfQuRSTnY7GBy9GtVSrYv
up+Jzj4FzWR03hX2sW7ORCZpvUAvoDXyOtaEVDS6DPuq6x9Bqh/p2q3GncRfmgqcsWuJCU30oP6U
Bp2qIuojGQEUuiDfCUVtxka0HCmKp+geL0kbxOSy7pENlyuqrnRywJ/dKIkLkspTOCRvbrzEhGPj
0h/BGS1gsBjC665NRlZH8//ZHVEbC/BojwBG7uLWjHDMw1LC36xza3qL6YbQ/AA9fhGYRh9DwswX
WmW/y38+ucre6AjuSsDMROIcxhX69l2KbWlOKms0T3knaxES9FsH/NNTp4euqQjOCxBIYVAq3y/L
wwv1+HxSkW/0Dh/q23MV4b5ZzTjVzNbs3zILrkJvvh67U2b4SJroJ/zZtmGczkqQSLsNc0E+i02p
Xm3qlUEUcXiYUeXFaWhriFkF73pcqeGxmj1mcr/rtEcrIjinYpvc7exTaBug4avZ+vNJUnNrKjci
CdjmwQscWkCMcox3htd0+6/+Bfu8FdUrIl/r81Brxden55hHANcd9UPMV0RgHx2kS60CHDY78eL5
RjZv4ZA5r+U3S+malAGxQu1tfwlAC3ORSAL6icPHryLBNZmCX/R08si+jURQvDbsQIBAr8rHcDwi
L9nsidNTJxJVRWrGGKP3uDOhHzbIUs62R4GjZdHEKeagT0HRiRRMQrEh576fA+LV6yIpEI1e083W
WYWdl1ItOLB2nh+EjXaTahICmh0t+AxM04dP/Toh/q9/l8nPTzFsiYkM9p9ydc+qhsAAPNLnNGqP
0OlRhrHMKY2aD9uRGzWZEANqm+8iuZOXOUmVtDs7uUz5Fl2qnOXM7U5R1ZCK0XrY0SDyfJczNzGL
/NymTnzpKiBs4tyybD4FB3QBpkG9aZBrIBh2CyH/1cHV34oedbc+f59u7ldO2uMNFvOthy3AxDOO
qUKzwLFIdml1XV2b7GHB6ybdb3KsEv3Dvp+8VOqC1v6AfjnaInGs2BIeTZCZ3CZhy3MixQotrffd
Jkz6sVy7jgb8eqGMf0bikjEpdQeWof52BCp21ZrumANieu1hR8mbi9BQG7FjK3q/RCS18yxpIlvC
6pB9+Y9PrnoxVh4puWRDIxjnfEUHh2h2aHs/ZA52/Z3jsTqnvH+/GVluykL3SaksCM3/OeZJV0qq
MBIbqPdDrk2G0Cc25zctQPRTndapJvbMsn5HnE1fdnfD9PH0/NXw60dTfVa0eTj8fck4XQSyhIm0
xmekwgLHP+HAD1KZJwsvTGJhcI4PbimZGX2rZSy4q1Nz6KN1MJxSqUsS78JFGK1a6ntDo3ZnAXub
4HqQ7qXekuzOg0kR+4ZOD6ueGCTFVk5J+P31HBRcSgg+JWULligI3iYr3ifBaLUUnHwd3sCXZcZr
oq9vJg1f811OAKnt1pxrh/52YEok+5Bexw1NRPEdLXkPXCgvwsJWssiPFJiwegEk1CuJi9yX4Q5q
pDFyZMBxU0ifLWQ5raWBlxj6q8DQgvNimpviHtKV5uIstmxKb6noN4kaXUnGriKAx1cuOHDcmwgx
jFoNyuXqJH6TU4v2pl9xf1Q7LLFIJMDtpeC70Crh6lwowAnIpBYqTgxRfAueyQyrCG/NGy4AEJyk
+t0EZPa9YxetaTxzctf59zmrTtD130NCSz31+tTfg94yCjvVpliKrX3Drwt+V8YoWcIiNXOtjlIh
LFHAlGm2vHZpzbRepSqYsw+4GogHKqIU182/IkLcj0QMvpyLzc0HluKX9HCHZy4jgtlWm07sVfkP
TgMsm/xk3bpRVkLLE2GPvbGYl7x/2kia/gNYo0B5qtTJ6Z/wIoC7XzZsMrfXJi5yWy2lGaos2ALJ
McS3pGvvtK6AOw3Q/zINmIBp3gjEKKIUPoWA8gBKgBs+9WvFbKHr5g39sP09kQEH9H4RQop94VFq
Wvpn/UjWML5wtP3Og6KOApHsWu/5ZojhFQjf2QgQsuoc270wVboofzg/iWknB/tjIuvT2/+4JGVR
IS6boVtlxrzoyYy53A3x8nkFl3PzotRlushPn3MJWwPxQU39HSULR66Q2MaYdgnKvTICI1DzTdrD
BNIUJ66EP6sp3hFPya7GI8jGVooxEZEE2OrgRHez+6n8YQX0bSJiiOQUuIWqKhEEDEyvE8IGWGLJ
DGI3CBncDd7ZPzEy74OKEIgn0gV1F3U9p53tL+9CRMOPPUdZqug3pn3gj0DNyMAHaPxZNwN8//4A
AUGAHzMT6VH9EncOK3inveyXZkDfKAqdg0qKx00qnHTZ0cRWTM3GWviOsW5hM4nCsfU1kjhoxdKL
QPNB08H2XCM0ktIYus8I4Cdq+WIGJPZFxrsLVTaNQ/GWE3zovVdOH4hR+hI3yqp4+Z7E9t+SIFja
JxgQ2o4o+fOoshSASX3GCnLgmDW3j1zV/en/uDzkr8KC5cCEVkHPg4ZwR8hUgEWFWLiWTegvtAdg
29t3GC1b7avwDx88vm6ntDkAOl5ckvl06eKZrfC16+0+dr4HcIdZ0eESgKfVKokjUof1v52372sm
x+8YsbnDIXMpFaDSs6GuGDco0kqKe/+X+jJ2TekZHVKrfue5OVE5jtqTjc2TdrUL6DcWI6vg2fnX
QXYpwKgHgHkiWrgjj4uldQMTWiKv5icIiTqZuuYKSv/dmfYhPqqgVWLM4Z//UBsqDFimQZvP3Gjn
mYP8ASA1+X7cLbYw4QXVSX6aCfcdg7j01K7CtzHkSQjVh8CHGdxnU9mZY4sMo+NCdxdPq63Z/7kN
8fDqlsOwukCl33zOgc32L4TjtKidDuIrGFZ5VmChpX+XPtAgZ1eCYgRu9EJQv6tExpnewZW4P24S
U9wlfndjl/Nu63KMf9NFGhpNVgtBXk/J62dM0jUvEYqtOs9gAahfFNJVjBzaxKmt40/xon78Vj8g
OD3yId7FPMrIplW53RmbkaBwrn51OMJSuC6wcXyENAHlNjwxRO1ktKUVwj/4np/XLZSTabC5odWt
l2PEkcD7JB3U7CeAbvkhNdhHHqeS/lVzMVPAj/v/wN+ohMwbu6Ig4FilX/6VKhdhcmW5XJ18lMHX
7oYXTsS8Q0h9b2ELI17a9ZtkaFfBSVDsDKRyLpUSVFRpXvzDDRPTAVTkA1UsRWvQrAg8iUEPSP3w
xEBNxcEDb1UkfQC0o/URqPyJdSz5J5bl4kuWkhkiIkUmK7o98TZOVgxbk2ckGJRS7P5j2Zeba/oY
9TKPMA7sN67X3D9OnKcTaajZtTtoJE30Xwk+jU5I6CUI7xND2xwDZ9lgW4l9UI9NUqxgIy6nHIiR
0AZIRWXQSuwA3XWgOkcoe4pyoKcKggyt6PbWiBXiYdk5qPiIy3ca6rZeSr1xrDmibPiW2cckqiXO
3jyZtfDRloa6rwxrkfXudDRq1/T6Js6a1CIfEjv1SFKUHFDBXR3x7PMncP61lE7JkqiU+do/T/Sr
+Gfib4nNZY+puXn0as5eKUCTPBeCRokceYjIOopgwIDchGNA/eUC6SuVNvkttlTcQPAJ5cSyVAYy
SXvl5CCtMnJHQWb+G1PiEAYVojg4qn7/pAUSLens1oN4oH1Swjr7wbP3T4XOYUSvsJ/Mrgu6iU+r
F3HwujFHQidBK+7W1VuYXtx7mOePWhdQxk0cpgdwCNW5w0dd9EU2T3IvdsyCJZ8qiuoIIBJueEgE
vB3Q8G6gL5vjRGC1ZKWbyeDbtUxWf8Qm/aBA86VnTxHtV0G24B5fJNtT4b2Jv5pTL3cC6ofM6A1I
taq8cJs3bEtmnc6tDMqxvOwk0O306QKa0M/HZOEztc9f6vqxP7/IBJH9noyUAE322UwnoO11nUub
QTG7kwKgXrgvVAokgYBEQd3s8ZWIXlNRVL4/mJZzXccpC4BftaqlLfCXgDBp4Q8BMwMahB93kyRN
tZC95TdONQNm9fEty/VT4zxIRF54nZ5Xm2LdAfTfTgqmlTO97TTP/sfTy3MXCi0H04m3jbhOofrf
I+9IgrHdePJThB1W5pllb6OrBrOWbQwl1oJ7cb0wbIHxAUvCKshfIdOvyNlqL3lpUyLm5b8RwMUD
KzuwBAFsIL8gWc8GsHMqDYMQ+FiqUf7uqbrCcn+Crtp10llXZgc+s39a0SlGVOaxAIC0Ghy1nDsF
8msjAgcECr7tlGT66RyZLnQdYa9TDyeEw6UuQE4a2qjOpx/+oe4SUfstz1VpAUo6BduS9O7sde8H
/Vp+OceuuxrhU0gfkPMcJexnYCNCsc0nzysovds+rSKdFEjeb3ITOOQEThkbQKmiNW5aLdtCdNdC
GPeTQuTk8sMM7IPVPtLqNu1OS27tGpSgDMZOqyb5CAtofOvBF+Ws84vgybL6Xji0Cg9TKKB9EJKW
xOMCqwaKp6AFOpVVya0Lpi7ToTWj9S+THy1W9+COd/Kuu/68eQ8VFb+v4kvd0eQeuV3BXEMfzmAo
8IRifX0s/jK+ubXEwS+Es3EewrjGcl/gnmpjIwbLf0Xi9XhXqMl0AJl8bcTvCmt6wF/6lIg2iqfe
DF/ZtbAaiBWwSkVUGEgiqQ4uUHIJVudSdfOPvoG31D//6QAZbCMnt7ka2qsHqVOfTOCtZtNFAyRV
SzZ4U6oUehN6MeAoXdCKrk7/K3A1M9w/ITPB1rsVOoGYpG5y+Re5FFPhrssZDQPh7e4d/BeJLi2J
nc9zFYYVc51mQTsiIKcFLiIEdeTyzk/uodw2lMinlKBqY50CG1TYeSxRM1Y4WJzOvJmrRH4Jw4Qv
YGkc5kI+j4Fq+cZ+C7e/N/6qIbNEiZEpkqwPk95vUiRnUFvnWos6A2keeK7AwkMPjhzjWAVmoT2l
M+RydfzWgYx/3gl/q9fj4ZhaeK/ndIfpPE4vwym8WZCiX+yuU5DKNy/AWw1foa7PCvLWtYmN/Qdf
12f4REzMN0eqq+ElR/EVGL555y2hnmxZt3DRGtGOGLtPmojOtyKNA6wm6ewCON+xjKi/3HJdTNwx
XeBk359EUxHy+sxms6cR7tpDK8Jbuqkvscm/HXUBZ4bzYpVkqLwbCqqeqcWWLe6+EOSv0x+l9Pu+
zK0fbCWPvRwJwn0R/xyegSJOTt8mvq0jecy4zAyZ4E11daNGa9RxpXs+gtbg8AbTjqqqnevamnIl
UUGXet3UCzg4vzBHowNW54ScQo1YCn6rXIMKfygikxdqgtaQyU+xLqUT2x2amLgQktbACxkv8n0r
5fVW9b9sHHiDyEiQOaUU0YNeG4ZJoNt4BqtGpNgvh5Q+E7HFRsqc7bX1TJSr9oRmLrSlNiaXnpSN
e9S8S3urP6Ruk87Wvl5kJ3sym6dwpQLw2cKXKWf2d2uQ5NG8YNuIgPRMjLmOPOFCzezoGSXmemqW
262JaAgIisrWGcbAy7D1kucw8jNWdSlCeS1wA4cQGoM4eD/WxCeyUbLjmx/tz00i9/LXe8p0+c/Y
gFFKKO+fVoR9VNTgnSf9C1gucYwWB3l71snm8wnddE4fsHkjpT+/494Fmeqp4GpWYZ5co/l5zcf5
B5xGV8sOcNnNc/92481tJb4QoNmbMrMS+60DiZ+Nj1G9uylg9qdUS3BT+CtXG6PQysk01l5duRdc
/Jqfgbg/7XzuMuLRkepNhnSPzqm4B24fzgtcZV4Fm44DAZAUNnryCJb7H71E4IFNwXOw1IVKPQAL
FGwmqXpyGjjyTRBzX+ag4w3IVVPsZOPVi+expNMPmI2Ad5rlf7pco1RWukaaEqGW/wy1b85Sf8wE
OdJTAcxGM1HkJuh2zf9ggKXsm77lBYW875SsF14/LfWl+RCELTBOgxWh6cJjpVWYucpo8FYsOBOB
eqmKURSV6rJilcYrjT4Yq4qicUKplnl9ji3n+WSTB/E0+nQx5Al20l4gIuSVqJVZ+H6ec/EucRsB
hIzjVYawgteBQLnLccNwvqafbb9fugwUR55/IgkSEwcLMDI9as9+aOdIwThtTjk/iyH0ySIndu2e
zBL7fVJONJeR+ZJL2YjArRZ8L9b7Dgd9i39Pg8qiFxXJReoTRr9McPnXrAnmuE/Vfb7sgO9+rpIU
GDP6czfyNNTrZQboRkj+jALyOisaWGSjiukJs7t08PYyn2vGGl6wZkE4wThP6Usz7wW407TOgL4c
QHGC2icPof0c99ZwMGZ3ETcYJjLgl328XsGkDfvkO66TJLVF6cSDSGeGI+RBD+DldVvgLqbRN/2s
HNoJMBF8aoMniylSseeYob6qp1SDmKudniEmV8U9fYGjt+Vx7hKq0hIRUZUY1EQVUkiQEW0A9Rsv
jKPDOZbUXxBjaKpzuQQjuyh76JxQXeIfkEzIA0lCLfudDurKM5R6RWzVzv/crAYwjhMudPDvCfKH
0byr/X58MxdGG2QRB3B81gsIS64TuO1jTG8dwOSkxq/ih55FT1Q6bWOISkkV1mavpcYP91ZDfHeg
5ec2vPKhRSwDA2jQ91WWiaaiLEucQR9tmzlv1R9SK6Cf7AWD4tGsjZ36QW+Mb4ZfZ7+dnpHb2NZh
X9JMmy/Bvs+9FQSUh8SQUXa81pQi3Yr+t2BnEGVX/w685ntxI39xf+jg+3D8WquEyi5DUS0U/5g4
9KvURvAR+rNb2R/lbuPH3hG4Fweq8YSWTY7cAxlbEczNs0BwzwF5PMkrZ8YHsNE4gKG1I2KWxaPq
535dV0k1gsQp2yWKOG/n9DI+l6Nk1xY7cF1Tij9hkqglv3o/ouyhJdcuKBqgYvrFwh9zZdmytOR3
eXpW4of2mwhZSPLGZIc+bhD/0lNZtdQIxpYo97XVG7zMYK7pwwyPEh95QazZ7EfyuC2jTf7JFYVJ
2jtVAGR5A1EndljGNBNeYORfncOIRWUCZT3u94HOnRBfeJNtjOg5tFwnUDQJxruUS1bC1zAuGpvB
I4cE6hFtbB30bJshsl1cXxewgsW0/GiXJ6dYQdiByjE9P2us32Q9WoXgjiPXh+74GWqaelKobYD3
cV4PD6J6hp4tIBw94rWwGveFW7vyBFISCKKteEl10qKwE9TBjyX34fh1Tmq1N2KozlWGERxTYuPd
z8FdESTboNOUiPXVOSFrP6lVAGBrv+NeaMz58oNEyDrGrJ6C14NWFxmcOpCp2O3aaLASAQPVZ5Ba
y0YJ2dbeODwmfHHIcK9JOABsCqMjnbqTQgCuEbypBQI7qnu6PLHtXSM0QLCptURkh2VGn1ik/PAN
VfobEgdUTnR0l8M8YLVP7hMIA5nSvsuh3cpylNPVvZtXyB3CvQUGhl68yznzdJIO0Z25raQFDg9I
JVFizCD6i5OIBqkGk6FidDkSR7lQKdIjSoCreOgHmv0skQVGnavDZP6454zdj7xCd2+ROzUfykRg
m8N6seOg+C7m3E+ehRfa7RguapT3QnotWDhi/ii1UOPi2l7KDI5XesftilP8W8Ly8XLzZzAcNG6J
AYEBNuSbh3xrNQVTshLYICOsxuqOJvxIFLEO5AG+jpVsbLfwFF1usRTIu1UOwER1+AD23tVd9UqU
XiWCqQ0/FEZvXTp8SUnX7dwAnknwV841fPvsj1xCqnFY/QX3C9ixkOP8RB/RdBlTnyOksfnx0cbJ
8zG7ncNkBHTJ5+Jmq4GOHtY35Q6UXCvnlHrfWZ1DGeNrzVKEfBoCJ2oeKeO//sIsX+xAvSHuNyiY
kfhOBHFESQe9wuMZ6Tm28DIA8CMV0Kn9VxRSU/xaEFNBDKflqLBnT7Gh3E94u5GJ5fkTff/2YFxf
4gUjgyCqSwOi6DV5yQBYEBIZRew993HaW21XgmvAUWM3SZjhKKQPQELl3TOHs5T6Sd8mHQcWpyc9
FLpIwbZEXgc2yoItjOdwXUQzMJ0bYSlu+1IaM/awW1DlihRx+5GVbWj2xjrXybT7E4UaEWQzz0hR
hDb1FoPmwIE/bTSPduy6fz5Ky8rcVkcIv7py+B0+wb0OrgxPXUNdLLrJyuWo2RWLCn0Vr4J/rjsN
w6dviDTJhL0725tLVeeqe7sM5vz5B9ajgYc/6ZGFxnJpqBrpfOd/P9Ib16w463QAKLSDBKIk4ew8
E4TEcz6juwKRtTRgX5Apjcm3vemOc+YKNQuMTsWAgYxXunruxFhYEBY7dJk6Rdi+U+ZhSTXo2f5m
Q71hCO+uWNjLIm0k5fTK1JxgbvXU26k3jMA15NIoV/MYzOn1vBz89vvyGo2tIMKpgXvFehqK3kpj
nxjaK2p/rYMA8CR1vvAKdllsTQnVXy3F3456XEMgZ+7XrVoQWtBL0r7pdZr/ebci8nwVo2XrUN5j
bRU4ZedgRwC3ZkZv+0h8KsESxUIjGd13BLHB2oV//uBWpUYoYka/Zw53WUmrL/3ytS9xz+mYsgh5
PWzJWeiwwBLbZZ0qOex1lmXVCUbjioMOQ3L8UAcnE4gf85MI2WiNIkHw7Xs1sMqa/Dn2JL9UNaGh
ED4IIRPKa95Tvr+FzLspHRsyeAaBTx9Quh4YxaD5yGxJhXd72FzoDyGHNMowhDr5A94mh2imKNFM
BgARwe2tGD12OBPPZiaPmY4ih7WI9CAUUCfmm6Ln1mS+xdWb2ZqGuGPp42kKO4IioMfFqVCD/FZY
ouBHkXPE3omIIyanDmdE0j3z5yrj/6LNjJzEDCt13K4AFllZMW6XWevyrtCDpHMltF6xwWhC3crL
zAD/0G1lH2fOAPlVVaUu/axNXScO+VOZyoW1DSUFkRyKcvExt4ErmCv+px6qMJI4V8suENsnNBjT
xegSr3p46fMqKCqVNIJ8wXQZpbEn8j1QtCrXaGGlZKJ0lXIByHJc/Xoq6Mwp7Atf59eIWpbqSRX3
8jcK0KDp+/z6a4oogMbyl7d/uqmFEJDIru2u4qDkU33DS44YMn3yKMOtQWBjxuMtsuXK9b2PFkkw
C37x/4QCvVG6z21TjMuxFuABcOl5qd8iSPrOo/3G9C9+QVQ+717gfEL17aI7JrSY5SBGYPQoF16j
pbmDPS9LA19FMCHuSpRNElp0T/JwgnpqT+28RgInl8KMEo8QFCgYno4INU3s559ANTsxnLqfveg8
jeA5Mz+GUXAzQbCi+uxTHA0RcNLxmwCNp0kJaNW718NKwvQtumTElRlPHgoQ8gXdRyUrYVBLsmbd
y+txPd5gIanQUSWiiSXX16NNVfUynuWUtTJ/J1qi4ea1/2gFL/KrcvAdifdc3I/NVuf/t++MQVUb
dOoQfjaULdC8kJxnOKN697IvLRrtfd16UrprjLqFjqN/t+OQTGBItaJhmxjVE6NtVv4GfbxBXeqA
dUUiR4+viw457HBsTlFcyEm6rw0UGgbkHbON3VUGTCDE5AHCB+eJ9VciFh0q2LbuFygQM2snxeaG
pS33vh1VewVyUy8rlIveNftZnQ5AT/1Q4vAYGENX+BtgqC9+waZyhhhLgWThVgCBm61p1iKe3B0L
TVBCjmdgpKrEMqH365WluThlZmbAnNH5MjT5zmW4R0k5QHazBDvEkLy1cmpJ2QKBzd6CO4Yxs4X3
NdU4NbjxxOobGZ4kpgkQ6Tu9TzIDq0F7Du0FZxx7J8y3KRnaK6yYZrUfK2BVBsyF9+47H+p2NQu9
b9Qe59bwi1dEm3PQkwFkIhlm1AIHQ7F57J/X5Fn/VDa71I8s8UP/dc8gZPozjHEewbC+1jRaz75z
gJJzuvwmmKk49aP1yf8g5DM+iOGp7rQBH2XUmtmGfjCHMorBpPwPG7HJAMzxmcNkgTJX0rm7uS11
WLO1J6TGMEnr/N1SD6nTQ7+9AeuYflHSHmBM8TRYcAIqMVtxwqGgL9wq02MZHS13TjLVWbpiTyYW
VdHx3G1mKGC/0FZRI/klq0rxUmy9ewwvtvUFEj/q1MXsclk3sLxHvuxVZcsWqHA9YK8xRAF0Ia81
Xvg8I7BYg8mQcKcK7deRkURFD+FyX8O1JGdFgf8hvfuX4SEH2cFw6CjmErRrm2SsoWJi+m/twaGu
IvpBT6fFDlqlnkQonQ2m007HnyNy6RiqzjbJaD5pb2MCCkv7wFg5YUiZ916OWJVL8dI+nhaJ16fk
dhTWVnpes9yQuzTy1qmPRMuxEy3ExskBN8CX6uljczMbDd0GpgNJ4R4xldhbWNEsg8dDZ9avxm1z
NGTjl9WvMdV2Khd90b9+npCezZaq8La/hILo8wQbDEE4hruIUjNFJVwLfw/DcNGOsvLe0t8I6qBN
ZhhlKMy1mxRKzC9eEhgZ/MYiixPzI7HfQ87HoKb7IP34LKOo7oVAcTe+Pd0fwubVyLO5bwQ7uy4o
EeZ1x0NZef2caLSWfdJfOSBQPU0nkLMcsOhyJB5HT+D2RbKY8QnZ7TojUvF3H6ktMm4LCOTmAg0p
VvueHAMY7xfCgxWsWj1qeR/LCKaKjeN9eZAHTdU6B/sTB3m7E8MLZuzAl9pfjEkKKWbELd4FRGUS
tcCu5DQKj1AFOch7/maDUe+T/Op15Ij6/wLtUZWHhrvZ/Kq4WeGvHCHMiA6vsiN/hny3XQGU0Znu
xRIpEb5RuzoZl05zalO3fByxkRLNB5u2eyt/qu7XmA+NTqMpteGlogandhSkH/N7VvuaQZy/R8a+
U1Qmiq1WXblBmgDIsLhPsPcZmE0SvsiK6ViVa6zlkMMly8MlWMidjguod/7yohPNK+vIwIcpkuuw
3lZGE7qEENF8FR0eMw9jLi767BuCZW+iOmPMEWfsvaAS37x1lX1daNQ5Iu+UJqgP1eAWhL0XKXas
Dzq4ORgVDfxnOCVHROufYvVUJ8UgOxdmJ8M/x5ixj+nZCzH7oxdMlRuISw3yJIB1W8aBcNTYMhmM
NXKsmNkICShNbDqTY545JTja8bQi3Cm5q1ddQo55MwWQaANWmZakw12FeChzTEyMjPTQ7+UAkezg
8W2moBJJqwtMaNP9GeNotyQuTz8g7FuZunnc8MLaWOpY5KRsAce5QqLXJXsWR8j2heg2mwtxG29q
ZtrK6qZ8LOnP26brS7XxvP2Jx7wXIl0V3+q1Vnyo5V7Gkk1SPsgvKQTd1kc5kGNA+A3nBemoJwFy
/kTgJnoMRsT0ylUOPLmrKG/mS8mnlUneJp6rkqOhLcQMbQbn92RDltVLd2zKXSlorJd7cjYffPOW
2EmxxzrvjaspaUHXtDUs8KlWAKZv/37Z62EEpXKN4HozPezLhxSF/+JceZr+GdMxzGOg3aY4zdzG
nbuZSM8YERGt9j7IX4ZCZ3vEN475bJ6JF6F4vf93nQ7eDnhVZJYzaZIlRwMjWtuqwU5tw49YTgrd
T8LLMsZUAw08JFbgylrLN4q0fzIeDaqjnKmM8pn7B8WpsGlw9tDmThA/BDWTAtm9L0t5YTq/HxXh
ZAaX25eTlq7+esZcrpMeQiwCvJ1klt/O3Q57N1JbLmwxhVbkU3WA7ZIj4/NhrlCk3JAays1LYNMd
2ZZsJUO7aknJ7cKbHVpSbZ6TTos2Fx7eSkA75DHpR7msnbTaVAESWROopNL190Yjjt0iwK5HVpao
rMdybAYcd7x9ZMyQ+/KiYlmIfaF/j7UIJYqVWkjawA3XSP1Et9wB9IXpS2dajworWmatudJzTiEp
tN9zgZsTjd39BlULAuxJ9vSZMakfLHXZaXilkwuhyYCbaQ15iMrU90NeXkEQ4shSHEf7YQODQgnz
wo+gLEt32+YimbB7vx8NwNwI9aZhq25L3FQoQYBNgQnoHunayO165c5+4V0fqBqs9EXHOKBCv3rD
eRiD5Ym+zIHa7SpQ94vDBRUYwpJF/9mC2/6+83Jk8wym2deNHDT58dGyfZziWvMPeqBPjTZL41HY
8kWIlYxgnMZ3ybRJppJ9pOZK8EMKVLOsXFFpk9gx9UfoVqi6U6BAZNEcO/Ds35snY80z5lG7ZSXJ
qdtRILHfVreE5aB2uNhBoGKUbXxvSE9brAhWHcIKwKvoKy1YiWpk9EtIuntPnzpRYsN/TLsCxGr5
/rYE3+0jrKje+s6ly0h7k9lWRRNosnl6g3s+gXcbp2CvV2p7Sv5dqLtc+FGYjQqcbbBZIVaW01pj
vePzwsMyMs3zN7jQQ/ihxOPzq5kI/RB0mGfhfAITXUGQyqtVfie8qOEM7x6Z647HIj3N+BpSlcLZ
Rp9TERcmNpuh2dO9xwird6OmYOnVe4GROuO1+tK4ikJyQieuSPOAxWZqwT8IRmdH9NPf3uujBDN6
Ptn24Lg4h63GL3jV6Du+ffXyJuSKnWtl/WPFwJ0SO11uUZIFFDgsl+Eh/LX0gJJu6yu71t+wu9DS
UvtaXUwrFO35GrqgSPUTULf6PU5U+QgNdPSyQWdoNYC6rFWSVMS8rUSKc+pIlssjPrlJ0vCSGQYO
qsTQyITlmlHEztt4pBj9+WDvkWc9W+TDfHVu0SvdWFJBdVxxfBzmRGz/paXeKt3tLwP+5AqKASut
Ork5NuV3gLo3aWRNFwIKMfx3G2Z4+k74o7Nazt5ncruyxti3IFxnauJtLRNRzMzp+TaIkYZvwP5B
9GnphqrfbnV/LpErZgN+RfjwK91sDEg7rkiECTsltf/fXGDXFBM7MbyEZdtJKyV/dAzXkt03NXEB
5jslp7VF/S1pkyPD95ftJcUh8eof0IDOhJnaYWmFZLQrGY7r0mBU5MOTUMwQzH8VYH8oqCM6mGjf
eNGxgEvD3+icCgLb4VNtr3nzM5X+f0tLV8qUIZAb9rwOyvL2FtAdZDVgLKDM2wLpFJYJGIExxosz
spQ681Jpsf+JOMiRQt17G7dng6wpvm67R3zioH/Kz/cXWtK7ZpCoox1iGHzvswItDikMXIsuEFK+
1AswM+no7BM0ZzijgrT1Kdvn1mQ6SNGSxT8wHAvb2qg+5Vecc51Yqc2vOoNa0klz1mpDyF6UiWnh
qvNOad5V+VlXiQXCPqLvnPqoQO/VhNUfYbGIoBG0ToVR/YR86jxvk9++G1t4AH4AseHYWbsz9wfz
e4F/6QX1bntRJADOa1v9HXkYzYoSaAgFPS0nV1iQVjql0rQ9B6XWEXEm2cnz0p0KAG8SDG1HL+zc
CwHStHYZzHL3KHfBjp30mzYAtudQ3Rxnnklz8XP0H8lISva6tFBH8vgprcoUxDBQbDza6f+87i7h
BJGNoMU2ol2xU2NjncPpJFRRNaQAxyhgbU/SipGTpXqGUBZmgg9w/poFvhHTfqNNFcYxo/dFWN+n
7PK6wnpMhGaXPMlnqKvvOgMjLcZyNeBTApRp0TVLN7upWK24qOlfUAagt+5AvEXj3nxb31CvGAc3
lh6jogvl7XFo9PJ2QBw6NggOy246x42dOXei0T/bzznBPcVceki19QCoMApCOyXtKGYUfUZOoWkz
4IaxjchzadvWgUEIc7gramICrDHx1wEuw2JP8WACrwC3dYbsJOiFthqwqJTBZOxgp5AxiPm1TcnB
2DJjcfm2jWuR4iAHl76voix1avQ1k3ZMViYEEjM6iZ+D6bFN/nBy5cfXziLFrOZcg3ihE2fw2Q4a
FKsB69CoQnfDKJEvE8Qgj8smDWg/rlHWRVXK+o0pqdYeW2wgek/rVRpI/c5jthtrDNl1SFpEJL1U
+MOPdEFEsGozPbs7OX9O+CXBZt8tvsJHcFGb5q0ba4it9hfG6gPXhc1/oY5FPqsTgX6CJHYaHeTg
sdaqxmrsOofBmEdRJR3KyWNpFIBfEdLpE2CCDnreazPRLtY5Dac2oS2E6vdarHesLWmMP0u52SoN
pe4kmp07efntJMAXeKLATYBWGtEK+SK9rNyYK/BkOye/yQTzpfDBzgMV/5AeZ+GmGgPGpeDGTIHz
CU2y3YEooZU/rSPcBl9+lbiEvDFGtvbWfR1AegwLkIuMDkoPk6xPrlwjoiZ6JOl6ONN9CTw7L/Ga
f/eJySNZKxrNaXkVZ+YK9hw+ucRf7Qa0vmdhblhKDhFDKT8WDyPo6nyVqY7mPWzmTTLLOG6Id8KR
0pl+i6B0w4/UD/zqZjwoLeCTDpvFIvP6JhLi/VrTGhCwr+LH97YdhZZk2Iq/ASzq/PLpLl/vPgAH
vhp8nHgsG59kz88tIBepXDVFuL3qvg+qXrvP/35H+9jLfHe58oIqPek++FdmrbQQwKobAPanIz1j
AibMj4yAN1o5NuDQtAz1U0nLYa1ZIO/T17KM30Fys2jTQ4cc9tgizPN614Bp7AiiYM6IAow9Uf6g
BQjJTHDGuZRzako3KN8nwmd4fO9HICNZf7M/nLubhkilPGAa8EJypHDTLkZ1Z0NpNKxpZEDLD6rz
0U+JIW3G8DJeLHmQ+x9DUHgw9hoP0LmWf2o1zt2O9DuvIJkR0PGGnCTrj7b32BjwNBTlQUmAFJ3p
/0G7r/dt7WsILnMoAbsD6oPsy64gwsu1KAgtOtRCwlc3VKmfhfJ0nLUjXhSO4VCtfzTtGzQPRJp2
tK1pIIR0XSkkUY4eeoA1oFijEe+pPisBjkou+J6WD+Ynd5zuWxn+xPk9H8ToJJ9uSgLO/iztY3lf
usc95Jch6u7AbM29bg6KZGNIlblns3WD60SLfApSWKH7JuoOfZyBXUW74VVkoItW+DE0xOlajOne
RI4GoCmSXDjbsuQhM+a3GYqE14UB27kB8RGG3KqksE5GhwcJzjuoONUt3ltRJjKClr2DtRTxj7/+
HwKGzaAEF40F3f7S/0QAjMcAiKsQTliNjcMzimU3qBD9LMUegMgWIa/H9FyYkoj3dAEUewSrVwwZ
NneDvfLF5lhtNoB20sIwH8F5ThzOibLpQt9qYlTrbAh+vcxA+qYINPxMVFfuMGUcE7snGif0igqY
zq4YsiJ1Akc6aaZ/fzlG2eoTPqwPChNlmcadotIGN0Hm8FQLaSQACpN3IAcxWUpH5qHPbOr4+E00
4jqA2T82kBFIqu69rq95em8Tex+AaIeqEAS9u2VDSBXbZpaLFXeWNcqLYa14viCzJttjULpW8fwt
1lpoT+UKVJMPit8RP+IF2eksecg4/U6B0d6VWRjkZL3Yg+4SLZVmRwtE7rAVt/ERUiGYl9MGxT8C
uEC6jRf8r4m/zPlkbHPk940WD3mVSlu6H2J4D8cjCEBTQcoh6ksb1noqyXDNj78a34O9Xp9dGyed
k+W7S0iUih9YOeTIQ4i+FrxfqD1nnbJMV0prnom6a4qEYI4kV1iD4SpGfhGz1zMoi+LB5EWeYkCU
91uEorSlXIxepaxFQw2Jp/Oma5bBeltzgB/S/J77T5449AeuWI/dmuenmOdgjp5RXmsi8ohwES8x
GIZPx9yV4S8OdQ8SPY09B8Jjaj8bJsPjxVc833il5ROvKFaRD2rT1bB/dxrGRH0kkh7p052rUWA7
BDxXkCepkxvlp5j1GOB7m13u87F0Xc1RfFyke9SeduXUAhHm4A2YK2Al6oJfQdJ++rDrzldTz2UC
Lx3JB0xtOTVDLUxrMu7+oA3wCxNu2Vu+xhv89EgVGqgcyuO/l/O6ZDMyqk45Y0IlbW0x17HTRw1A
CTVYcaVfQ2zwppCB23/lH8WhM86BEnrNkqtW5RXVazb70NsxejXky2G61jftpuTtN7Q2kNrrIdIy
RlBg569Gn0whTlFSuI13Q0bY5Elsb84laI/5Taf2GiCrtNQUi+79OBYMdrxyv7hPKDHHFzlOgvxn
Z/HiTwvo09K9GQobcd/No/vMXTBV4mYeEAwjqaOtCaOI7K60vyXaKzI/nAyYOelrz+PAcMTpSloe
BFsz8AymZF9w5k8dPXipJtMfHWm9w+ATy7c1J+I/tweiuDmqB8thTGc6jc/04ZmMar6iB2qj5Ghq
UOD7im8dVK2KzAGHtNr6Z08/eiJggkQdId2fHbrbQ/GAy2aR1oEyDzkMuICC67xBiOvCjuEv8FOZ
0etSGzE0JxPLLvAksjhFB9IKJ2Ph8lAdKSwcg1k1JerxnWJu0XD29LHUjXFoEGfAbyW1rrrYkhx5
XWYJ5SXkq2TE2ecJLq/cP8ZeTn7XD002XpxtuqbjuwdvN89eVsRcuejm783EzW1nPeHBAy+kuFTB
MiYfoVlS5i84SZsvAheZE6uZ7U5pJJ79NPaYD3/n4sHy29L7h2RPk+tyi9tYHt3wpG9wpCzIprQm
PCIsjV0J625Y9V7VIQ3flQyFT7ZfN8ocWdObt7a42+WCq69infhZatGNxC8cR1i41DYNz+3gBhP6
kHStQd7shxsxf4rwXhOGUvkrYGY18SrlGw0QTjN7zd0Brx8n0+w1vpAt1iYKWEGCBpYz5lDSxPuh
WHM1RDdipF9ODDndDjeTDqn9ZxFYiYQwUBBWCfFWg9Kkw8oLauyXzmyJDRmPttKo20MAs/NRor6E
OfY2D8SmJqNhKYUtw6KuyZBar3y77VsaQY57qWS7+v8VHHd7vwgPy2wBu8wqxJI5b5KrLys94/bU
o2VcYVWKlwjOLQjKb8Y3daUfCr6yq+v+rKjaWTmtJWKv5rHLHXv4+fzU/dKaE6pc7mJzIPiqiFR5
L6Np/Nzx7275CuSM1XyivT9P5Bxrh/VW/NOfKmflUbDDwzvofnNR+ZWAryr42x0qezL946hADnS8
lJdcIYKSaqTUMsy2kzcgmmQ562tydvcftQx9/71tNh9PzXbd9cyGj98A3lUA2RvztMbruN7J3H2o
2Ptah4u/aHqeudr49LgDToitmlAlVWAo99Cd8suicivWwt3zbED49GUggCI6K3dGA9Gp3WMiaHix
Ghh9vioqkhfUko5L+LQJyXt2ZsH1bpGuNzCB9lIsylWIepfbKcnWNhC96XPcqiFHvxbRC2HAtoi+
QftSUOkRT8F6HtQR5/CxNIPZBA4w53B/zry7ILUAyiw2i/WYTWMUykgcffcsvCb4lwFlAInZFNEW
FC2iwO3DnP21aJsm9GJhw7RSHOXWMQs2X0Xcn2hWasvWTwlteq1ZwsSWCxk5bYyVQflCBegMqm3D
GO7/2zSd6V9KAtYzKY1uE6JI7cUpsQrTEuENf72v0jlTp6Kp7HIsKQQDclBPm5sjgwo+60A+jQDz
IHh1bpynm42ZvCP8T/+DuTBIfafNv6rR5vCehiF7qXxI9kqCNkLkjs7NCwRTrBdf79kCpYL75mFT
JuvnerWjMnrFMi/a/0q28tMR3OhHPp8eiOom6FsgFhtgIP98u9ujuoBfm7nslKuhTtPiaZrSmApr
b1kJIku4aF38qVNfc8lVCHvNM2nFJPtlL2FwU+2ROfd2BhgTCXvPV06ZWY0p9+zdiOGAlsF70Emw
D4yB6R4xKSrdZlC3E+Fatg74n2olibMyDlBU6/kxgxdQjrwhAFwF19UImC6bWJN4UAxSRM7dGT3D
y2u/gi3cUmizR32+KvnZ3yQKC7p/DVEOBs2Wdtajjd7tmK+vy6gLEicCIYahgmKg4Y9ZEs0pDbbf
uxju3qJAz52k5Qe96QJP3AI88gsnCleiBu3Mzquwf/9NlGYgErVv+ZbnlvHU1Qk+XES0a7YpSPH9
iJUw8cG/cCw4ebRjs3il46ANxtg7f+nVpAMjN+TqoQJiwRZL0/+X2Gy30iMuifPSj1kLFY72C1Ms
18Vb7moc6C3Ent0qzeeXmoGIwAA16H75f7t4u7remRV1wAYqQ4kGyOBVIvMMfYOew12DSSAW87qR
W7hRr3YPphmpJ9eJluHFRVrhRKB7oaR+kdJ1JSPBuSztQa9T6idH8myaN7pLRtD+SRGKJbzlKwqS
j79L1DsMgNnq78sVV5n7oK+4E5HMCY/v3vMvDw+m2vS94UfvLQG2uRH2x4/wpkRlK30ManAk6uY+
DuVugjUwQ2Ys0Xf8NPVAZ8w7prrjfhS89BKdvz+DjvhQMlgK7NccufD3306Hoi/Pir0utW2eG1A/
MHx5oa0flEnJJNbcuEpY3RUW3+Q4ryY2rBWBIdBtuXq0yba85tDMhKvfZWJ0KxdR4WPbrFDZaJ5r
OnMkqzVR+MusH4D1U6LC8G6LRHtLS01rRItKGIUUTIJG3OApsAe/rdEDrZ5QpFzQMR1zDhhgDlYM
414o8rQpkiAKAnbeERFoGtFmTEI3PrfGL+0X1stwGaFAPkryyIkkZOSxEb/3sufsIlvDX/MB2ieH
ZtZzVPXfPC5HARTY0dCVhWyjT7fBxgCv+ZK4mbrQa2K+Ha4uwNArjqZTYXzXeVsJPaCWBytDh4UR
EayMvw3Qi17HtzWnxe+k+AZ4Y8DTtVxTyLgcn4OWZarVzjndL6ujnZ3JaUQabkxzhCt++J3/zu4v
DaeCeuLDMkIafQioW+uxTqeO7asf7uqG9eAor0ONr8U5D4cpfLgLVcSW85wBL1Ht4B0ElDI2UaQh
WK4iTI3wwQ+Adi8ftcl7HuVBEG7K5Ge94RJgNYhLikdAFir6E6OH1sKNwoPzmUE4b/u2fnePLGis
yGw9O+7yFF+vsP+iBzLg1kTEVUZQaTAL3gDSgDuvN49/9fqC0nqxqT4TPn4QVwXQAzEXBBwmoDy/
Jhx9NVyWTX6ZjsljtRoHF12nJ+ayNCzYqqMLqhvaaRTOw/J3BTMl4aCko1ME15wVVXFMBPvdi6GM
22GXKY5q3yOBYh9o7KWTLaMB5PlQuh2ff6dmpjsrTRN9FpLxT3ei/wNlGCaMo6bGc+aW1LwTEg0+
avC6ZjyWSpXUkUn0E4oeC+HGrL5/iOsQ3TyUrZ6W5T+ZtH36LwSqUeurL/KIzLyicYxdzkdfGj+c
a8BuaOGiw9yOaD9OZenyFphZxGSxEbmWpQWKycvt/eqO4zNTpj5HqrGR4nl9lZ5w1NXoO2QmzlB8
6kZpMCqMX7Cc9IaO8BhKSpTH71K1Jq5qb42/lr/qk7PHDngl1cvwNj9yIZYKMgbfJtQe4A7+m6bW
ysu6osXKK65+yXOpYE68EO2qv38BuMH1grSFA/mmtV95MpYDD49zErbVjm3yCCgcZkUAii3V37dJ
LYCM5vTOn1yJbfwFb1RzKPJTNPk3zK4xeWm2BnBq4HWsBH4064plPj1NBtMUst5CP+k2DGS1BNor
QzUuYqcrSXsPKc2J1Kw6wP8QJXFYOj1fFpRLyd+fRzmSEsmPixbHFejhPj99MDYY9ida80SJVSVx
QLHUQE4FEh+JHqEujUW3CcbwmLt7INxwt6hEHu5fwq20cbrhdZsEbiIk3SzoDd4zRi00ymAkWGxw
STLDkOfnuLJ2jusVJaQjmcv7w8huEVvBbuGupH5K2p0NKynk+hkr7DNAtWsD6RCSdnnFWtCRgQHZ
b5APFb2s/aW5sCiWXgzK1Pjpnq7VjXXS20QJEiQjPA2rewILevrpu/PSNYXhSXWimTgRkz2NNguP
sk9iC0DPpzNJ3poF+dx4FiJmhPcOIULTaeqP7Sv0Iqo93vfW+0qwVSuhO3rsZR+KlmluvMyNTJDj
6maTW6zEUEtUdKOQZ+JZzYQxxh/sxKVHV5GsqQd0Hj6WKk9TKEdxViDQ0v7CQO961zDVzvurx4ZA
43l3d6Aw4RFRhN5XRIseLrE0KxtNz05LJfvBDLCHzeg08PU02BLDseHuSQzOfkz2yDwewlHyOqqP
mbycbKy7T+zYReMH1vDOPHVOBf1FJ3ym1fH1l2W7FJkdZ1QTKT1AMQPjXOFOtMtU03BMJIl2lGt/
vFlO56veRioY/iiMKWzhDCpiz582WLKvrUY1pHaqftgIYuWITrn313M0PQloxb+x/2hyDz1HtAYG
NREOfKDlBQgtFSITc9tYcpruMKKoWYi5nI8LH3NA7X7x7D9yfnFE2hsqpImmsxCgkO5EzznV5Mpc
TcMDDqNJFs8kv4/XNifoIrmO4lJD2mFzj2EdKBplARLSbCiqFBw++mZfp+GxKYmRVb6b4MV4xAt7
KXGC4TN6jqyATXsNKlwQs/uhceIBfJBr64ZBhxVL45QAH77k33USlPyRjrRgpi5B7xGVPK8aQQRq
3vcz53R7xrIsCTf8fQPG8OXwpv4nPpDxFX2kWfayII5PS/qbqXAvgZAU6LnK8WOqLwhLFSIo7ufO
TTVli80I6ncUuM3s+dqXc3oI3AAs4dC5ncYm6jY7V4CsjwMeJUUwgJw2RGiyKD/mLRrAUoNrksvP
9M4jhZZNIFwMLCvZ77lMzlww6Ez02UtDZeiEhw4F6o2GDwAtXAdUndJRxbhCeuh38g6mbSipcjSD
Y6YxHgZPIPOvRByCoWlK3TC2qm4LVEIx4hF5DyBC/0z9uUbewEGbLzLm1ExAIZcCR6jUpYVP4skS
dQvM5L7EXx6b6VbQmtzuRU7YurZ7e6/XraQdCgTvwDYyQ4p0J485WsUtITDSiuiwRLrXLG4NSvhA
nWOKUHXSzBsAMxQ9vskFcezSQfSGsk7QRlxGb1K/JYJ3Cd8TZ3NINFNDnOTc4+mmRNxFm4/7dqfb
E4iIU9/hXX2alKIIdyScC6vDjhDA/zavvIFxzm5qybpo1hORcI+P9g1ZcGU+8KD0v1O3oUJlU900
gFSICLw3zw760KoOx7HIz8GallQjviZqZ7xUC5WF7JEkm82C7N+Ee2i/jRojvP/C12pefWAR1Tz8
LPu5izLUwJ1gIchkCOBXwMlZv5gJEIxa6sabNIvNlx4V0CpOzsV2MuPwhOCQnwfYtKiFHDH12wTY
+eyGSmJ3Gk5uYJSvBM0IqFD1yCTkKuX7RVzE8ImIa/BExKcGLok2S9DPn19TLN0cosgvFl5VaV+Q
N5lXrVwXIWzOuu3yNS/vj9WvNKN1v+3eABrHnE/s1f2teiV/KoR4nH8BD7WG+VNS9rWWkpDACTP5
lrdzVnAqUN719Oq1fx2U+7jobJteQMz0nZcP7o+DcSr6WVh+aq3wOqOVB9tjeYvuNH/twwjaoC71
WVCCEW6VUUL4IH/1OQdoHepeGuLiqnGtyCazXbrfA7hU2pme4jXCgtmTsZ0tWRI/PUEfLC+PR/pw
Tj6CULkQMgmCVcEi+Sleyc9hVrBxAdOoJxblkQaZoAYZB/nyVeI290hweXSWNYsiDRk4lrJH7RHK
RVDc2knl3gmhIYaFKn3zUXgt1kh500xP/RDKHNaFZ7X769XIilvyZcwZZkh2b0FrG7mHUSDfWQx+
XE8mj0lOhuxQfw7U5KaKBIkbERqrcXwuXcSX29GxWYphULVU7G7li1ivcd6bmtth9Z67hNJf41hH
mH37cGT7qdtKYenJTUhEu6E9ah1GpBO5xBQE5QBsc4NgYPCYpTND20Uzxhj1JHv4cFBjs9nGwudg
9Hjep7oMbHLxOJLhegCSJDGTwqq8n4Tw9gpQ9mWon4DhOq9TEMxjhy9+aUHCdyoKDpUsxGZ+Wh+k
Xl/pshsUOQQhvLvWVNfQTtOZIhvtBi2G25r5bvgiD2eerl1bQv/NxtkXCrdNOClK6Zw+R1it1nmZ
szO7krs7HsBCjfclbmIfQ5+jplfElMOfk3Fspzi/q0MYQAYmjHIAg91sNHyPfr33jETa0fmmIXlI
1V9lXKOptoejXMKeCLl8KBVimCMDW3wKHMA0LzEq5JkAtNm4Z1nUeooDrFKNSWeDgfSWC8onj/9y
1pSzV58W5ysu0FX8Qv1BiTG2FGUR8d1wXhUXWLazAh0XYFQEswV6wKKZBrbybg5XnvOXGTQpD6tR
1C4Hh0hpvKnotOgjUPgyLabUgI+kdkwxTjj+LExlY/tslu/jV/qcOZ3qolG7Ifgye6SXSmG32GFw
4MqmdZwbVgy0tSyYOVF+S8kGB9YSwOeQbuvTqcslzhYSAO4lzruO57oiqUi5T55cJZCuMQiZR7Ip
MIaDWX/2bWxfS9cNVLCyY9zTr9kJ92m2EE5YzyHmm+FqK90RNIfcBbCzOegtltS7Qj0tvHv9e7gC
eB6hGZnRqE8eF30/92DnRYodm0GaU5uGcKOifB77oTNM6tvcn4UlkpuGGm31pqVlb3LMj2CRZW9M
749qpHnFEytX1pSxUAY5CgMGg5R4fxagDnqMllY9zU85Q7E8aV7gY9sgGd8/cjEQDA6ukbkF1kem
PQSfIIzWVXlsky36HZegYMVXbHfxnveEKZBVfwESsO1mCE6KL91WW7TOc5fNgUStOVwmGLBxptjV
4d0auLbufYbJOdGl3ArfQpIN6/MMAFjhDODj4KE/O7ojtFCxbj62KTqr+I9gMvZf3ruf/gFzOfLn
gtZMA1Gc+lfJj0s31h9rvV36pUJhYW26vhm8pa13ddwRUa8QSvEnIyB3aM6dsYHCRtD8DavAqnJ1
q8q2j8iHfxBRHNuMO4+lF3Zc0and31zyCwjRXA7x6gDVAnCoFPKioXDP3TavbxcjDSGP0bOzoL3o
kZgcuKVvlPJ5ArxI9x6HnzYwaqBnWiSZPScVDEL691pvftzTsz7/vq3bfMH6QL0FA9XnOf4DQjHK
BE7G10V3qvO+jEIoHk1kCB5zmLzFLUJosdkU6Sw8aDG2xqgfs0HB38A0TvtwmrP8eYGYO2B3Hqv+
D3gqdghOawcJ0XwTarP1ebnoPmO4KWmOOW9s1T4xQ/4tW++kRCfdfVLZ70SaeeLEC/JIwkLS13Jz
y6ZgfDe0KlKkKPpTAsEpdrRZjnKIB29E2bRlBZMVSdNadRmmUC92Dg3bZEf+pQQynja7o62QTZcp
XbR/qJPBb2BNpOC2Klt7fBULumYkPcJrkysvBJdpgXdCs0vckCaxDjJyK8GtkzkdSSS2vdFjFWJC
IC9zswPUoCCre5/LcFON1SI91baF8a33cx2yh6rac+qdyfAaKUYzDWF6Qe5P6g0huiqfVE58Qni+
YlJ+y6YQyxbmevdxMgC8lyjmppEIlKey6TxtqYdk+eXHVGXwAOnKQP+ikLhWFg2dBZHhoNr+cL1u
jL7WfD70FnOO6LmwpCOdkQeXsf6AVKtTgujUhWgQYR6TeCae+2BulDkdy1yAO3DQUIpUX2jJQQht
C4/ONyKG5iGaTpG6kN/7xeJh5q7FKVLxm3nJu9HKjR5seNYh6BUGDGpoOXrrhTRx1s97NFS3gSl9
ddYtAjdB5NVta2c863NpxbV4CFIaftl4B/6khHFVECXCPS1rnmnpQIr0nNLYDxAf4NJunPZ7OOsp
hL/FSdVvzB6qUC6bnKrMI/j/OER29ALy+fSfyb8Eb5v5WFfrH9/xhpkEMCw6k/l43HX+SsuwQ5Hp
Tgu4DZzwoNzLhAWkDJT1oawNfnCDOMCZkpCv4r/iRK+C5fbYcx5Yl2rxkvqzHXR/zprjdSZKcqGl
yMEKmN+xZAPWf0qwrNObUnyTGV15Xpf6c5U77fQBQIgnqETT98rSae65smZ8hK5e2A/TfdwVRALl
175fQ7CWthn6dbTAC+RMydj7b6Ay7NgXVLLyZ2oM7XCpDsaej+pr0F7aPe8k7YXB6WoNkTLaCUpI
qFWKGccysSgPGi9D791VXo1pfZvnosstIlQNEfw11dnY4PABXQK/s1q5saD5ZufpFVw9OOeK6c9N
2PQW95ZI4oKml6MoaTh1va84oDw2b/X6gRXkHT1QMxwXOL7CtTCp5f62tnIRBJhZaUhuypvKZgC2
q5S4T1zAFGO7DfIo/oB5gM1vJO7LCSoSgVgfOFK47VbM/qppY7kbg16MmJD3jpVihaJI7dHa2gtt
zfpfK0VNyAE59iNhd2z37T1nWyMIfPUyywtf+JD+gJBd1vz3glgRmZAt0mXoo8sf1H6kKDh/byEW
7KzvZbQuthuUCBg20dJXhwtN6MnUOQ74w9OjbiscRKj92xLr5Hw4aUHikOQPdTwW1BW6oMsbuiA1
KQaYfvUP+u9LbMTpEFl6AtheqThxSH5sdML6NkSbX9quBBKrBVsfuR8aHizZZ1DBFKqJSvYgROhq
ElY8mNNgkV5jE4q3e4mjfVGPhNX0C+KUOLk9lL1ig6atLGMF5lIHCAV44DHAxJS3ecEhKz73jPhQ
o3mZF2YAANhFpK0UQeGEHomtbcWrdkXMQWloHwzg7HUCFCW1LXs9aLpLY2yAlniOqZc9HznuNWVF
X8kTiJg8DFYVYCZOEY7n1LLNHp4+zmiTwYg5V9VQPWMhLVQVdsvK21XPN9T96IQV1kHntdjozSLY
kdelhhH5WvfLYFgKKhXhCXq/LfujucStU9toLZ5xiE6O6iFg1QOLEfbTM0iTLlzi1NpCHfRLot3j
rFPJOSKIl26c13aH4luwigJ5e3m5LBcjWoF9SC7fIOs8zje73AoO3ErtVXBmiG1Dt3MA1HbpZaXd
fyMlhr3SfIiikE3QO5WxfBqP6h3JWCRtgD32yromIK+9cRMIj4DGuqFKIZZfCsZWvMWqWX8V9hMh
HX5COoAB32Q0aylrG9PuueCARLVcz/twqL3/1PaVuu6T9E/jlEuEiT7BGggXBrtQrwwv0refmc+F
p+JVqQqn8Jit813wnh3S5ommTACcNgpbDqcQtKdRKQZ8Tp0v3SDQ4AlrsHrAV6Mzxv3tsMBBKm8H
ZtIjFgYrxFLw0B/+mzIHaBKt/U8jBRAemFaqtaDFCXqIQ4afjueIR2VthIl0W/caSZyKK1+5wkbp
MCYoHv3Gw4wDR5OYdXN6KjEq7GJjmZxGZB3XQbV197HcX+uVocOzvzIgydfdrGhpl8gp2zlz51sJ
0+tg8Gv7Mg0HsRdje4idqQJsgSYgU84is+hZ4jNxYQ5O0kA7/Y2yWqCbEoKFveK7y+Uj0R+jJ/Mr
HBsos0hRgRQh6Dhimx644tSj10kkje3zTOQ60o0IFg3EKaTYGp7kMnU+6bl1fasxFs0LgBc77d0F
svC/G4qC/RiQzn0sr5fUJvYSbJJwkwxN8KZWeWEKoEeoqR0H8v1Bxif+B+aWAJg5HiQ3ql4rRE7A
LuabHyXGafPKH84UbdnEEukTinIjlj0EIoz8K1AvqzrKwD+gxrrk96a3uytVf7T6bXK1q1+5QWQj
AZbAJjdoU8NTPbXu7JMwGcS53d6ei42pKmetMO/14ufUliDgmr0PSq6LfFz0yZQ5O3mGfXO2SmPI
JZ28oSbJN5TfE+wnARK77IXhJUH35vNxIfJAfxjwUAHTX1Lb88HIWvldUUn3t97pb2KQ/ocaLDAY
DpaoOni+TGpH+bnAGdpPOkhIfolkBrSNjFP+xQXYOLVocnwddyDMq5Y7lZIjoJx+kzo6m9ZslRaV
meykSIRwUp52A7M7gk6GMFxQI03Vr8vA8Iay8Qk6hEbWcH/xP3H8vqJSYoNk3sgS26qtx59lBuuE
HHYsRXJsMDVXsXCSuxSPB/r/Z9QA7hRg+QyXUFOUN5wZTVGicvRFF3F38xaW0MXacGLButeNLB+Q
3ylqLleJIrenJHnOlXHNt1CzGAW3i88wuPfOzwFu8hPPq3CbXCAxOiC4W3oACCTcg2A4OhxojbD2
1hFNC+yG3xIww1xF54DNkIDTEDLSHerB/3HlLR1HuRQMWdEGxayrjpEb1DpdlWXyNBSQMsu37xCB
KPBpbhNsF/4WkRaarwKsf3GinjzXxZxZlXkOl9E1i0mw1rSxMqa8vm53SxqAWWtpWlu+LPqYlQOJ
szUMVjQaXzZ8+85AhHTnpy6iGym7DvKZR6p+fHYAxYMAftAsOwg1ujFDTsYHLPJH08GBCDnnxkB4
5nzuH5BPcMiMnLwjnws5c0yUW3lXBES68ZaVbxeZnxDNHKQimK6Y4eWLq/+fDYXV8LoNppMaruQq
ixosYOguzsCcZHV0AddjII0TIp3WTo/T5+9UCVK4KUz+7woiAM87pMjqX2b00DaegL9JNpLtmB/x
a6MXgxDsotDRuNhpJF6INjIyulxPRrkvlT56XsUOqYKKsmb4b95XmiIUVCZ6TYt6qXBW+gZ4QsII
G3Iut4Y6szk5a6BNtTRnvVMBaVHXFoo4E4nuv5//HBp3hBHk9nS1b4sxNvMl+xN2hGm+nGxanUuP
yY4Nk9O1LF8ZLMkShnxc9iWkqLP2R8334TffYAk2pRaXwcdJFEMX58qijTK92xshc+gnSqP40eYc
KCUEKI7pXWnhohEb4sOZ+eB2ELUkMkSrc0diA6i0Qj5QHUnBHALh5AhgA/Xdn4a9oRNGZKuDH+VG
3gonCYW0hklvFd7mp196RevfI2uiK0LK0xkAxoyBRTcBzC6LVoOXAtn6PmZdvv8bKRv4cO0J6r5s
YIpHrxk9e/8RML3tO5bVyjmp3aEqSxjypZP0Dhav0samgHA4yXssAZYq0nzrhvDhMzTZMFX/8H3x
61wde4IdLsvYAq/kQsksLxO32hdhDkwu1wFgZS5DHAF8yOV5TqX7SqiGe6EpJLTKJBvChd26dmk6
ChUIWZ8XpIP+9l+9oAeA2QKiBB8prGaesURYZGJaloTmL0fXq5k6s4V14KNpizudgcNQ91Moq2QH
edlK35MoT+f/lazz4wOjO2B9sLOGDyJEVcLJk58nPiVPeZfCmpxb7GLOQRBlIOYFsE9burplOSQU
Zp8/BKuHbwa2fCAk951c4HANtDNrOPAwApCddpyVE+S8JyUjRsSuFzCQw4V47JAJ0KWvvM9XVu2F
RRyxFffh83WOcmB1M/unH6e1ioBpyBAEIzH9vgYxAM/bdumKZe1rPXCqPobOMKoqVs6Do8gfpRzw
4yjC5U1HxmFM/iBCM67TBWqZ5a7a9VdzXnPjA+CdgG/JyZxLIXsgjC8f08toJUDW08A9BEgebLaW
Sm8X2ngkmIFkOzVadDvzRs0mESnRUNjmZWXXgfBGdkkXl2CJk+IdtYsL8mmRBEf+PqLqVmSWcJas
wOLzO4yHg7VZUYRIgqyPBZt1V5oKpqhxLuwHwB56UPtmIUhazVg9fUbNVSpMBp0A4QBd74O78FaI
FgSs1yNaGYJu9jyprcvGmlhwV6XP/UH5ezfP4vNUkw/Q7ZMW7dqw79cRj0sDmcjdjuS33pPxbbuQ
bZfHQev+w31gC54BBNo4QV63ULBXRrqBQuMzm/OA6nH70z7wJT0Uou288ro7ywnwmxREy23Rmyqy
z7f/EtAsex0fpj4nHkFPGGyp824QX0Vwqivh+edr/cv4rMVqebVBjPF5kNC0TEmnSFDqIiVzxzco
5tn93JUvLmL7l7IJ2/OUz7Uxgn3hecMIeqO/EzaQ2Cp33PjOIlPfNh10vxmfeRYWDNYV82TvsWwr
mF7MvIkT7JWtw6xWKVXB/kxq4TwA8cY/Mb/pbvw93uJxO86PdMvEz3XWxYzfubaTyESQI38dkFzq
dySDxIO1clqPhhFmLJLd9CdjzWRugGeXdsmcQfxjPadfX2FfyIQm71plu1K1LocuhpizM4FCJ8fj
Ao32tx/MCIdK1esgP+5mt58f8Il8lOBnQLqyXeAWXfjbRySNi8mWHCxKD7yjH0uFstuZ8yCf5Luq
yzZNj1Bh2MKUGmyNExJYv26RyajRZWVEzpCrjQCDA0YgL1rVs4lSYvj1rUJw+rMVHEdNuvQC/cUh
VjKeXXDwnWGfMiEz1G1sMDUxnGS4yU+xz9EFMkPppTbKOShOZfDLEqiujKS5+UfGxa0Qy/mZyLGa
SsUmlSNpb4Bn/hLFkbr3JHff9oCWo63sM7uZ8SbitTkuyEWRSn04z7zKDdMSoTAsC/JEA1mJXtL8
3z0b22ClEwqjh5RDm0m7wHyoNj6+GjoDt3tIOfvXbpEHbB+BvTkcVQRUmQB6ushbKp42kWl9Cxnk
6vkps4YAlmMtgwi1hYVleepViU7rC95O7q14/j67T5Gv+KRe6WUXHcDmz/2ifXCVgVyfa9J58A2y
gq3HSdzYfOrZYnJeH2k9k6i5YqyDK446B6uETWeDd9heeZ9bl2t1yI+XLUgJ/cX9EEsz/0ycdi61
ciOpa+pfnq8Q9hTR7ZukPRDlBL1Q5olbFSt4knJ4SqPdqNlmrGVsFi+lgDYDzzaSM25x0zvRuGvM
ec1A+dzpk9wn5f/xzoPzNj9Hc9kJjGXEu6ehZYY9GqQGCjFZ7yzEO7e63L+nxrb/fD0YQb5+iHMl
g+r+MjpmLNlYz64H2Te0sWLm1Xcql1h5tFD5UTuqczJvL3kt4GOCg+1imk4teAeXsyQ1LpHjxsMl
XP/0uexS5+MYq2ESQziJF7eSpyoV73IcBBveORR9HRrEPVzahL/5zhNWvPTDXn1WD2wIA/LSyJkf
Eqe1yFDJTRnd8My3Y4x2iPjuDeblabVH0eGKz1cxeCe3eJOR7FDuL/MT6cG3fSbpwV8lu7g8OSVI
eW3yw8rGFuzJ9RMKiq3yEzuDagPvwCilTVmADQV2BmmRBeStpL9dAGszifrn/wcQCj1eV1+dHqZh
NfOu7CQfiX89sdxlpHiNAQiVVbziRl1hFE8wWvz4aTr+4wTZyZl/aUmjJ86tnlcpEZBTWSBmjyBC
eeeXuQOubzZNCZN2MDBbTGtkjHnMd2WyjJDe6jIwJWlx1A+Vl93fKYNu9ZqBQD8unmCTm0C94g8/
ogx3uirNbxQfexkhM7xAyMRxLUmn9Xj7P/BCp/I0CgyF1alC4mSSy4eInuyZeKKAtOaETwUmyIZ1
rmH12539hiJFoTkvXCZjWjiGblXmCvMeNfvv+5l2qZgC9l2ZyuHqkXdV6HDhWCYiMH7JHhaIzI15
eNXdFVisGgejcq+nFGKnkiETupWfJ/Lk2YeKVx3hFiVfmoDytQdMR6gpKqSbmppKE0glEN5BQ7Rt
kU9T6UUvqfBttccLO1w1evOVV06i29mWXvle/rZKRO+AnNB59oc9tkbOhd5eYQp43+PS0uj7p7fv
XdFN/2GxFsctUdTrmitY4X1P3WO4KV/vCNf/CKLbXsVwjYQjQxiNRnh2g2zzm62eHR+586Zus3ff
EDmLSWZAS3yNbk/kUzPRy09TE/w6/fQoACTgcvY0pwVTKyPkuV+VoMV1JbhyApYNWTghX2BHROab
A4wA04YDAc/53le2c+/ayCOAw89V9trQG6Cs/bFVqWFikKEU/JGOsuHnMsaEM2jNIKEqzdtMVEHS
RRs4+0zeV7DdqihWi/cdqy+CjDUhb3mG3bVlr/C3fwsIbtcBwDOa5jSk71n4lytfJQDBH/zaoIzw
pxezC+o2eZKAzdWurl20nQuDgoyoanqwG6U/aSO6kq6M4mUDEmimVsldrL17DVFcmoC2UeYg/0Ty
J7nWKxL+Vdhr2IRQF4JjN0fMIR4rkNYdtoi+AlrfqHSInKXXaHYdjJXYnAxMdDjzaPHIh0ZFIXLT
M1WTgVhev7kQzg0ze8ILn6CPIjr1rF5RkII7ZLXy6gtR3TTmFnWTnqUU1qiCMLY432hIBsc9Xkvk
fX3Jls++JSTlglViYjA1LIbuOWS1pEdDkLto/UO/JHu/kOZwFd3PE7Okop/Vs0UwrQ+oSdzEtcuT
IVAGqA4iy4S+woD3zusHVL4SwY0a/8hI7kEOhouZWUY9N+lV4HygnN+wF533Tda5HqznpNg8/YXZ
yL/Rby0j5yEAlJal5PtjiYjGR8/in/edPU4f/ZqOQfDekE+U7+yrovP/VsUITc1OeShw6LFvdrGW
66LiUOGsGqQ9la0uAGZ9ZMZYbGKeu0aGPX50RAq2sEn+q8QSbsDjnvYGjbjKKmuzey3upkeVxoF/
aD8xDz9hSomw7IIz0ILBSg2A7acYVcSTrGFMKyYzXZE+zO2l6KkQn98cD5082/h2Qf2wnYv6efrf
o8Dx8y0FULxKq7gJHqOjwfOLNj4qCSlDaQXOgniEXUMJAltKIbkQ/+qnI3n6aUeMgPIphy/YKkxO
IbwadkAhhVHF0vpcYDqt3g1OLZC/G9TM/wAdowW7JB/nOQoaHuWgMp5vwY7AtYVY8/8tJxrdbxv/
74ID10S+bGivo5kq92DwGi3wu1XxVmxMAeXbMzmrHA7qqJCYZPJ2bf4/3plggbquosnJRlAVaxnA
gHN7gnF8oPXkGjhsk9MQkUiIviiMEsL+O0a5LvY6PlFInF+biVGqnlUnBDvASdilFqTNPjSHZ7W4
RpzDZmY738IITg36UHv9naG1KVPHwmUSQowKMSk//oiEnSfeYlKXORQkcGdgoyjONiiXMYDC/IwO
XkN2M5el4AuUjHycHCQE1QEdOVVo95mefoohXSJUQsYw9I87rOi05jxZ+zw7ef/zsgKaXd9YWyNE
3dcOWstVnsQA1PDR+n9ucU6xlA0LJhyhJKGtzXW2IlDlgaD66ZDj4u5NqjS2eBPCHPq93Ml5GXbd
PLaBvEl5Yk7H3oDSTme33r+GUwJQG1LSZP98AtacOip42iDMWrMhMQLIc577CfdKZQVDIug/ZRIw
TWgWlxAb5f4OOWcdCR7QofeCA4NoKuapqyBaTPUfOamttJCyIzqULSGzihvHy8N1dH7xJ21Sgdsz
TPT/3hMDuI6yjLOuwYpBS1ekk67Skv5pssExI20aO6/ocaFvDyUoG2uQpyE11nczS/8CmzZuZ10Q
l3BkTDmMsBwgszBqjfNHW65xzewHhwkHezm0cOM6etsz4D/Bja1LapEdkLOIu7cFmwCgIIdnbKgz
91FsYjQ53dCZAGNK7/axnoK0BtR0qZE4fpuKyU/SQsY294XOS3kalmi6q/3yAVGtb8wvVQoW0G2C
Rat8WSe9OI1uL2o/YiU/pwf5gNDGEsTDQefv+23DztZz1doNIuhHp/FJZFmyBYTlXIVKw2Mu06Cs
ciHRKTxbVysucGdmitcZjzsodKNA/uGFK/yyxTBo0Bo336c2dL1zRjjvCSfGDZSAURXfM1fe1Tit
iTk0GFOo6nYkvsmOWSnsXX7097Gt8xnvodsI4CKZX7x+xV8fJt51RTx8uR6bRWQcqJE0Z92T1EYt
JZH4/twgIJPQaWoGzXXkRb6BUm3IQ73tPxaIrklDy8FF5VdLEXaTxYGkOwcNKANEc/6m6pXmZnHG
cuQSoiS/m1O+QSJkZL9wqb84RMpLkURiEsvrr04vun5l3qh7rRIO5DiZJpIgpdmARtzlc6sxrr2s
nz4Uv+1TZ+K70ijOH7QmKj+vv2vEyPLclqvjbYF1h0wedqmYXMBjPT69kvM+bAzFQJaYoWyE8GpW
KDDmtKxU/vOQeNDHttUddm6Rxr+BqnLWAvFY/16wIWa2jal485xZ7RqLgVk4+JclSbW+UCeWoAHh
fpbfvMqfepVX8wSaeeGqgdBdCl/MX+zDWeYF0DsFsOugT+fwpNNW3CSGpL3zXIokVEO+QxOW7pAO
2eGlUbVCiN794RkZJLc1yUJqADCrvnfa2DuY1KN2dOG8unp+akP5jxaEV+nT/M/dex+qShHECSTf
JeBLOtZC1WIFgxwVviBxVU+wHGjGG427Gyh5ek+rI5jWWoVj/sQLqzI6r5NoNQLqTntS2WHIM+uq
9pQgOaN6G/6fiTDUj9mALQxpX5B34+xnzPPvY/8n79QXJ82tLYpbQiiHKXeFex58VEuEqmmycEXI
PorYDFfH8eTBSIqF1kIzZaL+ea8Fy9K1FOx1AwvC5/Wl3g+prZS52TC3RSGri9gYxqHdXpOf50kG
eCVVlv9TGzwFlBoIqLoBYL1hUT5ylsgT8mnnrk9gVSxUJ/yxMn2DHn7y9G/bftbF/HBwQN+jNq6O
E3/S3L73NtkZfJcQWxcX/et2NdE1iJkaDlIXyW56JaLfOm/HExGfjPVucl3sc3Ne+iLFZC8x3Gd6
s8gff6p0aw02yBnjYQEw1c97K0RjOHuUZETsqc4/+EI3po5pixSXWjfq95lnaXA37l3dFIBBXYFh
dT6ejyAlmWAPsq4Q+VGkVRXMliFgMhqa4m/bvKiV/S1h3lynMG7LoYDgo2BiqW5G9m0FN2EzESLd
1NpdHGmEoXf2DVXs1iSe+t1Jc6uD5/GZ5liUJA3imaEurwStvqapB+xHuGC+oRLmxHHYfbrTUKcz
RYCErPZLz2jYPDd1k/LnjP18QpqcPYPXuw3JDZnztcBa4SZxb2LwU5L3zg3wSJTCeB22SGyis5rN
VGFfKrz+GWxtIVDp6TvRv5gRAtsleLZfFkWKuYpqDR0wDUgdmv17bpf6E4G4xuU7QlRr9AdB0mlm
48VgupVrVjfi9/uZSOh/K2y24FPVFHaG0BEqAiPEP9IKti7hgE1+hrRwusIq/YUlDhOqYxcbACbc
Dmd8SF9qL/pY7aU1C1Upwpot5BDQB76uKLP7zMmt9ij1YTL8QVNNzbL729Q6v+7tyZoYLyKhMpXh
VAvSwT5TsVjxoHcORPaXryl8w9mJJwXWah01oTp8zqUDNVQZDrvuR3bzD57LzqMGjG3k8jZG7r2u
5/Gs+G5dIw+cPnBo5TanXMM3CI4zEIcmXKqACknKlbZi/4CKVZ5abu2OBAPeECgSD9iYG3XvkDIS
0cobOHN4mf0QkIyhbE22wuXl0uC99AaT1RVUmhHeoSQxQv06BsiOo8OqHU1Qw01dSaA+5NFLj8O5
KO52Tp0e8k1Vv7+3cbmXOQ7OFOOALllWrf4JmRjn0VvZOAgZEl05Ooil2/Ztw0NdehEXxvqS13p0
SarC8RYLyqbBuUP1mJOL/Mnu2yrDCpD4CGVvdyKP37CKB+14nnAiw8jLQJeslQGRVyndncOOY7JN
dyRQzQXExcfWM2NxrvGPPjq45lOTEukTtMhf3IPsK14/dHvk+5JtIpERMxUM38wyEFfWM9qbu9xX
/3CvGmXHDTo0j6KMdlW72ePg6ZywgQDMegwktksr4U22qgAeetNRuIbMj46Som0aVQuyFjFv+xVR
/GN53im901DKlVBuD6Q7sHgAJBbfsk4AVJwGbWU5ki1pDpxktfxO+mzgR8QUSD+z8i3f6ot1x3dZ
fsbpcA0X4IvOLP3ocaCwhVRDXaWjpTPkddoSt/OhhRtHU7ve/CDvX5/XqzDneAFBJ4MKkixS6GeL
p2KtYP4dOS/wkjHxKKq7e4yjr3dcFI0vjYbX06Pren/hmvXhpCwX5RXr0/XrVtoRRHjJoMgf16F+
D6uNkcp1Ra6H7hXM1rD2r8zeXC6Mqc+dBJqNRajJIfXQf806L9DxHED/VqAEklLBFlxbyACBROAu
HVAEn+9sT3rTDr9TB56zyA+qiSXIEPPeF/PN9prebkKt72UjMhRqUXmysfbS6yAigCog8OU3pNPx
p8cG/uJfHBdg1DDPZmlNELevZufe/3jaRWyYMsk9I/K9vg8DBNNPHSYV4rmzfVf9XlrC36GCtZeH
zW+nkwCljsYJlNZ9pG1fhohmCGoEIylVqYIljxL1K1dLvphtISzBP7PB0f5pGm3Scwigbna1rkor
ZuEcgfwCoe5cS4egT5N7PzR++U66mdXcBOuGPRTVFQLoh3kAjchFgd8jwnZSFm/+703zpfNzOpFV
hngtT/zO072qF8dEyXdyWcOx3dSTUdwGOjIzyvt2ktGNbqWMNIIPLG8zdGRxz45+ppn3USoewWBi
zERMw8ZTFb4ApPUFnZeRC14BFmDqatl97op6fu8t86VUDwCOcWZgGdt8LYXSyBAnJOIBtxo1zyG5
3cD5m00HlyGMrccS4Nvjq7dQs0/EpxjjksVfnQLB+fASDx8xOvuUqrg71wS0gXOgfvg77a4uGpXg
GY8gbln70SAjexPUfbxU0S7W4DCCIayPhvE3sALfdD6J/JrowaYZ3OvtcSL6E/nrhQye7VJn+P16
clYjuFVAqQXhMu8+psO6zNupo9wyr0dIq1zIHNVlFi4G+N43VMRNN1c1qtmR6P8APa91Jlq0vEUe
C+wzv/c3tN6s4qNRDAUJkVBzxYPFWAdbA9cP8d1DkqDD+v5ZwtKLZER0ODczXEH3eEku1OFyp7VH
WBfgfWJ5P/TqvoLw+exZ7wftGF30lIrS4XHclGy1b2qF5VHrwJUOwQ0E874uIh9uLM8STaSRKSu9
Njbz2bfPAz+I5rdCRx5oEjkxMA+c3eObcrFxM1nHODXzkjPz0QWnCjHVw4exzQLRrR6HjsA1F9Ms
d2HTcqkthCA3MF+rX+utmLKrmeJ3qDWYQ8MXq2uM5r2yKLIFULBgmVvBwSnyJ6xIqtG7JhPUolMz
ypF/5q1wvt+fwaYRXFmKSnoIz0TECMePaVvy0uQIkazrTZVdT9TINh08RQa2KOOZFA36Bn5BzBZV
14YcwZdvOlJurTgw7xY8IpgCfFW5YH7cTqBA1LpgE2xMaPc4C2KtbDXmRjMrfDgvox7XbGJkQrmS
eWsTOdGKVxcSCLGPy1kOEI5tKCDhQF/j2AWgNeSBD2+6+euKPtlsy6WRnOZ4JhZiGb63t4emc/1Q
01AIpiyP8qRWI6TNind5baeMKPPgE8It+2UUs5E8Co8AeS0K9uHCbQ200g5GLhr8I/oWNwNAJVoX
9isimYE109z6IqN1fNesZ50D4SttL8OnG773jvhD3iP7vsB1b9WSMPiWSUcWuF8UJC3Qdnf1tYpH
5EIb5Q6higalJURYqFqXwXB/W0J+8JRV7y/Ryn0YFU4WuQ9rjsKFJok70qA4PdtF5DVd0ERUQh73
u3CB6WZorN+iwA7rathVb31jd8nj0LeRyqYyPIixBdsksIfv7xLoymGoicmK/OtSqD/YmtqfSgCg
U65+MRyB/DXFsuwXfe11C+dqHQPffEMyo6DxdxTmMiz5cABbSCfvb2Dxm8pvK7WR5AW08F06N3Z6
/GADjtHBcn/kXbgZynH4aJ6FAKaeTMdqFAq3YJuVmlhxrqhmDY2QnVJytV10KyKxMelTa+yObW86
WGAwlAHezbrtFzSFIeL5/1+LrH1nv9qrUi71ws/Mew6czxi8hMYqajMlImH2XpVWz3WjDqCJOrkY
DewcGEpoq1On+umtuZLl9Z9nWF0Xb9s6bJWoJJwcDzMf7OIuNMP+CcWSK8GdUc7s1neHITUUuylp
CVOfir4PvPcRSnfc+HuVKqHZp+HIiyb27beUUxhlSouvaMGsNreawFOXwYYtOqbSSZQSNPhBH0gv
0QA1FzDYpzLQ7N0CNSP73WQrRkRPN6uAA1dUfqKYi1gcVCcYzrD3DvA2ULKHOjTTF9Qs5FUZoIov
qjgvfSJMnl6KmEyDC+iz1AZFZmau/zc88Qz8pgOW1H2AtNYjv+uwF2CgqgXMowj+7jtd5MoMpTdQ
4hQiYXkBqbKHp39W4iVRMsYhrjWEiS0whw84aVVfffRxHFYqpbJsywKSmberfWS2iahDb2CD6enk
HEhN+p9MHq4EcKxTcD7ez+vPYyVakqsAhNtPULdi+mb/XsavE9ERgIhx8KGbRrVnJFsAwp6YYy3A
Dq0QyLazdQm/4JmIZTvvLXf4ZQvtIqSCkC/BVX5a6akQ8Epk+vY8vEyI+qnUeO+W5lDY4AEE1/E8
GYO0EGlpCytWCz7FohSkUNTUlPZz1+v/2Z13KvXLc+wzplGwGLyR0QyFEUu+bPGzLYmkVZGrcwPg
q6AC8Ev4/XSSH3KfahiqtS1avjOTz2lIOAUugrZ85UXpx5hkRtwzfGC/ppFzaT9Yh7e8mHCTIY4j
dfjGrgxmXcavv1PD9gS5M4ZJjYJ2qYZqh51GXGp6j7zhgsv8m6dDoNAeVvwuFEWZMPU+33Tu+Zp7
mUAgk0pojGqy8m1j0yjxAJWhTMaNiCQIOf9xznhPCiPV37thZwByHiNXu3DnT6N15wx+/AHIkU8b
RsGDoCPwYqt/d+y1V8+gM8+R1uMpfWFj0SmDozB6gDFhwmDK2s74B7gYmSscch/XKNqXX4HoUQGz
6aiue0xqaasfFrNUYnH+oBuwAhn0n702WcETzcm639HUXZDfAJrBn5FycVdz6OGboz33nqGPF5Ss
+niFrHpfDB6T9psh4xG8dUDvgEIS/0JWieDk5r+mwR5FOGtGlF3qLpru/RFy3JQZtLI5nw7wjEK5
hq4uTxqu1dKwxdADx4EQFGfAopQg9vzyNVKg/TBBPC8t7psNt9vBZcsoUW+Ow4yraUhoJyOryWJD
GGu5nAOLg3+/FcGYQCYHjmpCPaWt/r/9YW0zgL6RlY4lNFDKBlc9B91Z2gmkhMEF2H/ENobD4t0/
6M9pvJ7pysRSQ8ELmoQGU6u7FdoBSBhPyxs/RZzLrFOhh6gcyY8SAyJcigcdcaGFOp5H1bz1p4ET
zrO7rgGb1tl3oePSdLTcZnb8955vqtWmNzNkZb0EQU27lNQOAcBSiWN+QMGhOba6ssiTBm7Znebv
Tr3s9qTROZmnMyWz+MWxr5+NPLWynu52veP7mlDWoRTufOb+2G5Uv+/hGe/tqSikm2NhxpBrYI+g
RpvUhS+EK52PxtGNK9lIVrJvPrh4l8Mnekhlzoo3QIaDd6XyobnrWPGElPRq7oTxcWpYKhmPp/p5
YXwRTusIa7wGqV5IQQLudNRpawugfBe3Irqlw77DcPVpZ5/IxrCNTv658E6LtIjOe5KTB6r4dKpd
oGYJVsiAlxHQThr7nyU3ZWvGbQDNCyiKRlqea66oPzGoe/CYSbe1RmE7fVgbygQNm7hh5HwpGiWz
Lm2zU2JAAIbZDQhBAC5VOUJAd9aNRaBozMFET+01wa5Fbf6RvQc3lNwDJ5LWoJVLzse7VLQpZt6b
94I+27/G/ABcQP3RLHAEA9wYDUL1lUVKwVdnNmVz6GSukysTQKuj6WkTAdzlYPAYChF6UC6tCNwO
sda0w8L0x+wARYXUrsVjd0fVj9bQ2RpiImq+AuPUXuLLYGq8xy0kjuVurcVcGeavUW/XgX8uRzGu
/Mm/6DFQawFRkkAuGorNM2ghtQ6plKLnM7fGEBnDfBSUdRD/ypjZY44jx2LTnl9bGuIz8IYzVQDl
4rPll5tdHBsCNS98niyHvuHhMbx/jcqqXhP4Dm0ZjkUmMjkIOO/HNxfALj8EikntfDIuy5buLwmp
D/wV5gumKq40Zyi00/Y5X3URR9F2mjhfyn2v1bT55ZooOHZIT07X77k1ZX23VKygotniSIhicZ7K
ZNhqKhurX/OmWxs5F17uRnXpaQiHl6/duizNqtWf4V4U4WzdBCF76JebUHIzZmP4x/8q7ofvyo3E
nOnzO1PV4QkBFEUHDehpwPTKJnkGtwB72nbK1xZCvpnKi8I918pYh5hRGIgICtPbxek8R/k0UpNR
d03+6EwlC7eLsAauCRlxC6HzfmtrQ12R55swHdGw8+0fyMJUVNd9JqFHyXzU4siE2XSOxVYdoaMH
+JEvaO2X6+Pj8FrN1xQoA/lwmHJIm3+M9T3ydMqEiOMD94SLZdFPfNH/OxX/mtspmsEWZOFjuhdM
Q7jTLKp7bEP6oRFjHXE9dknZJzApyFvRwjxh6iWvm0APjUlRiPZrUBG/PoWuRmvwufyNUD02OEMK
VAcssJ95Wgh0VjsFIkkwlvNaS14zj9iKibgA7mRkFgrl18+1IuIWPNSEyu6UPPiZGKtuxwYce1xl
LzPVj6u78CrpJpVPdVg5aLGKc1yObZPXndthiUFX8hzsLo6dW8hMt0iJuhyJkogq4+qaxrIDciU6
c/FGYvU76vfjLR38JYxL6rAkTdqPkF6ZlewNFpAPkBPZFEgBLp861ivgvBR6y63Nm7XldCMrolZr
GTrITzXQ9GmqveTpKCXJTSq5vtfVwNRf9GInzrxDv5VAP+ssD5KpbX0jF4M+ele+zPQpeHPjOUPk
7ElKROizQFG+/IaIZm6xebGCU+c19D/h7ISzyDGQIbqrB9drk/Hht61MRXZAqZOfrxqyyQzDu5Jx
46xDqU2q8WtF7G4RBFBw0a0HPoGiwHjl5U9gVpoQRHHIvFXITgSv1qiK07pgsyEGmeUEpfDXir4n
cbvGUEwUEZ7pbiIfRpvQRJJLf9P+3u9y7gGFZIkqbBU5vJWHdlkOginxKQXU34e2DVjnAnEmnauL
i78z2DwbCPGXQTBN6Q0kz06SwpJvA9vUrI6egDWQehW8ODIGlbVFgMETWb5ikExstZMPDV8Mbmf8
5Mef6hOS41wIJ4W3ngA7kUB5RgGlEC94WR2xz8CZIxamzU59/AGHpaCyWwP33d4RPBQPI9OhzaeB
o/RLCFOusXmG3pE635r6Fv8bWSBzHsoOvC+Hbez6aoH+n0EsheOEe1m/wcj++cdnfXjGsulavhgN
+dd0Nf/68do61cIlyrcdTeaC4RC6vKv98Z+wwW4LsJietwcOT9yVqlTa4icvuOtQWsEl/VHhfBLl
MGcomAPbN1QoHBjz/+CkXaJYe1t3md2mah3OQrsywT3ymk3nTU4GzMg6iOw4gWgpLuAg5TFWAb+3
1PGw4VxxK4TegBhR2x+xy9jrHlETXh9BePYw6QbMg/i0MADWW8Ho9z2fg8zKkT5Jh/l53PVuH0pz
YrVSnc0qOHce9E1STlyfNvj7bBY46Z8a0W+OVwku1RVoYnNizM+iUaXTcNNQLCQhwP9FvsOKg2Yc
VTADYCg6MUjetUiu7bc4g8ZjNTaYkSmU/c7eZHVoGrs6qt2TCKtcUVqE4yGQ92fxHBWFjM3TCcsl
Pfree32EQ3/JknH5R72h1FplJuBidzazkGsMfSzLQkWIut14gSlYRNCqXAAp/CxgntSfs5hOA6rP
BdmLHjQasXL6r8CiWj6Gr79qmoklxQ3q7Se06tI7A0/V2SLyo/tXG0syG/IY7lpYxxRPzKtH2+sX
kuc8JkShDp7YaygDk09ob+iP11dUeAZlf045FiZZQJk6kWmbEKH2Wkgks8wsCP8S6QWkX7hhFJM3
m+yvlvvoy9tvNQJv0DXL/j8b2zoeYjcm/z/uU4iKmG7RQ7m+lp8UWb9LKCzA1Jzxmud+PjCiEqXK
1p8+OZ2Z337U9Gn1SouqSJTTgQ2aWnZCePe9o+QZ1bib8MGAEXUObAAq7TaxUYvjy7pk5UTlQWYW
X7BII926VF+F/xJcHF36GxnDW2QxLfny2HA0yVgFg69BYcVpHs7n9oMIQwiyjSebm8pP2jXHha8T
dgLIoICrgD8s2P8DLg+ClFfRMUxhUv7ZM7id2nroyFaFdxqzWwgvIN6u3Llim+4aDmhLX2Ua3lUa
NEkR0P/erHB8k5tPYZe4pK0lN5trn8kDIpoMlC9SEPNMmfWrzKxi/NMK0YYgOWKJUTZvVR+QZMP6
9nubNqWSh6UvgpCVzzHAsDLkEO06b2NZJ1QRsA9Q27y+QK71f1V1F4lV3aFJ/lOtckRMMz6KX5lL
4n5uuyyNFxCe/iRa8rL1YsTqJjzS1S6Dto8O8mQFOg/KdKuwJmcwubLk4lFkRVLwZqrIxc4y8/tB
iQzHXBzeeyxWSHm/F2BgYCFscZdHbo5kJRutUdFRAAfzdyRfm+FJFep5LJgGkN1HzujVwUYjUOTj
GHpHfeGjEkT5hcoi7baDM7Z31pMJA8FMpXZ1e3DmvbTxyyWKluZ/79Az00I2ZtGg3EAw8YvGmRfG
yuloV5lGoQn8KcGufdFnhxj4+gC/oNtycrLI1gCIePQ8jbRxHcVCa3BWFBfCJFJqCz2ajy7SUpJE
WowSiX9p46V8hg6N+CHkOiYD7GSHDnZAxnsYuxMWpB3CCd1Pg7H15NoHceE6t6PW/s1MNvM8+YZ/
Qr2na92egXMBoU5KlO44tAK+GGRKomOnOscCCuoCzVrS6mqM0JmbgZIDNBb7t7q/q853lJgJWv+i
he9ieHeS9UofSDYWkanPj+LaGiEWjctbd/QpE5lRzSSGqTBs4nBVKUvKlOANA7eVUGDCvsbCgK0w
JtwRRxzRzwTe0FNmnAN803F6TgE+82LgpAFRYoYUy4IRWChZLxTDHESKExStg6in1M6r1RDDAnCB
sjVd8wu1ig/be+VLimB0DdRbO2oVUY2wbzEWn7S2q+ZZpmvRIxgTCAaF1itQX+suY71KuYK4Prah
zsL3WeyMlueoAUFS+pCTykhx+tCkKDA1zxvd/TCIXD1mLmphCE3STVdqn2+qngS0Bd8YOyBP1IFD
SRxSb34h98Kr/866n39cT/Q8mXMJlddLhQeVZ7h98+wSAdAGtKB9C3W7DNwQKc7tJ5gzeSf45MqY
UzbNOxkIioVwxy92wbI8jOoNQ5Am7phgV5EkeAEgrRAG0ye4HXHY++ooMjTj2+hnPz/ee0eI9bG0
00qku0PlHtygpNgBFmhm6nSbstEtmlJWWUwf/C61O27AQCVmMmPj2hoQWM6tF3Afp4sleIxVnzF9
s63NLZNJc6fnAgcSaJgN8D+rIDYxIuU55KlxRGM72LJip4bCzfmXkRHpSW43WyahMMUhAU7PMHsj
ykMcEi0QI54q1B2/XKCKcywsF8SeUywAjp+ealT3abMOdY3rQhDVKEd0VSr6GuT3TtJNkJDiYQh6
aCB+MpN+zwPe1TGk93vRhw8s4xL8swWWdkmBW5jQOq9E2Dr7FPduW/OX9euofYErln8Z2hHgWPg9
58K2wBb2bztuSfIxpcikdBaItvpaq/1NLuBrj7kCN2oaJclA/CRI4s3kHib2xz3bX5eaWIKMS81v
ktb1x7Jz0PupsChCtZ65mxMbpm3sIKW30djIpPIVUfVcxtJjjxpyr1ulwCkwojp4cHIPX0whuPRu
IHqEl8U+KTAkVg0WRD/GUkvGCGGOYp1BhuqZsKR7PPEP0asGiBiHD0+7G9dB5lsyLh0mpCNX8qf8
/MHEhR4A/oy6baxzwtCs3H7iHCYs28TIzxAihepoPuGgSRAk2VfaocYZuUTbzZNGCnB8fmu7efCK
aM6KoQ9QEpv+GGKVUm57aeg0/HETD7SS1594rqscVgEVEpa/Z0P3p7iE4gabdn0SfterrEY0UKhY
duEWgK/mj/MEt/HgEFgSYuG9qUvvOVeGf6zHlR2UJv2dZ4vHmeYEYBJpU7i2ksEcTsl+bI35BhUu
s3g1X/UsvW7mHPQ2jBAVhboKJa59jQnHbjL+mUwA+xfdcRU/wfIXxliP4Z7IvtoTF7VNVKrwajcp
/dZSQBNo5xX95Gfu39PvYsFdNTZ7YKGqFbhPIMry7fqRavMzg1GCMJhtjFrKvrY5VveHOF/gBbON
abEK3v8S/g1623l9V1sK0m+8S1BqbVTt/96j+tBL0Qi8yu3DPoDYiZF9w3gwVznrt8hqjY2bG8TT
uMDGgybyuLv0Rxqx7G6G6GrqhC1sVMEWBQ55ZLFA2enhFgVi3FyHM93CK6uZPkN6bkThNyQ0P6Tg
IO858dGuXtBE+9fuFkEbLjbBhfyAxs00cyxDqk2THx4DN/76qIaem0KU4zBxkMRjfOCnckbTMvAK
3VNsihODHykuglmDUHjNgU+5Ws7fF5WCS5cb39IQh5PaTWdt+IFfuQ3K8eBOioaM0JFHE0jnndG6
4arbUyTMjNRbY9yFKy6yCnVb0ISzZ0SpDLAAD+oWXYDjEufyy1Vzy6SH9XwzmMoE9iPhjvjQhjCy
EkU4yvzgLdY1h7taukl8QyzvT9VD0avuNcSzzyZ7BX3OYB5ft8wB8yh3PQ4PU90Run+YuY5GdIPT
RBCNQloXVxA8v7VPO9XkLeQBiP977VTri944ZaS/YlS7Ow4dcrM1aTzMCTIhdfuHMWbcDFQ1FwiQ
nocin8wlt+ERypcUgN3la7+jO4aIXDPjpnjisQKoszcTkH2MZPZ67xje+QvbCfFRncAPTqR+fDf/
voZ60UGi/RMc5WBM488NyIjRtn1TuTsvmnDzf6yvdQHFJmm0jE3HMndSNdjWqT1/FNhKOXSH+gy5
yM/sQ7xrtPquRZQkD2NaOh0MYNhj5kpDTnrRKhoE31Ia6HDq/A6QcM9dXBsTAPWil0NvUegNGIbn
rZ5GxOABxAD17EeHtM9bTHX+hfiri1PS0VMWfjLZjCnR1aO2mgv3wh957J0nWp4EMAHdmd8v2P1l
IRf9vP01d2DrLzDbpSG+bRC3TFWkpjfaOpzwpZY44Q1kMyiBtnnQkTFFcVWgCAw40PcsPsaB7KZY
UW8C5nPy38tU7hVWB6hHaSFV7YIG1vAG7qlCJ0lwmWpE1FtDGC53ZyoMCMy1RrjyuB6yH6iAofe+
IyCKahZuSLjWZQ/TFWJTFBYnSb6JC3vnwQ7hNeKe+tzAbAnX+wQU7+66c5FqN3dUO/n1V/YcKmcs
XrzrhIavpWXlJdb+r3HbjlVNloEc6s9C52pVl4DFiiyaQc9uDlNl9IIBY/Hh1NBiukJyToIgp8th
m2qq8vWSmXjWHXzMc/E2ZynHKqo3n8DaGSGNPTjG2IlyelVUgvI8mak8L/ckHnRRzUCsRnf+sLJ6
tlmO46HQ3TPfRpeJ4lX/5/7x+KTiPSll2U7oNeBNsLjQDqvtDuM+B/g3S4PFVQl8MO4qmd2LAKWa
e6xyJxuTyLOMyYNLUgoYPqRLXEs3XxFhNkoiDg0U6x5+8jqRb6o7WhwSHSYjXPHg1YMcghoSrAwv
y/u3sN6g+DCzSMazPHmcysEpsaK1In1xyGk2xfpq+VooiERX8OboVJBLD/+pbyFV1AROV8NQvyOY
RNLa4ixUcPkYzigwb+rdjvh5plEoc1FnZR+4gTHB0Zq6Bn2+i1LCnrKNwVCWRqa/8R6/c6EFDDj3
IWkBaw9OvlbP12iB3jKNP0JQN7jdCp1PXnMYd+4fYzYK0LdEWLHbtOKbrKyDMEpEFPpv3kqEscwQ
If0dRs6IbkWXHSmLaShSOQEHSt5nM3RCWu4u0v9O5Zz18QCrvulnpjjXRx4v+vqBMLoGoCtrXj1m
6qMSeLE0TTK5B2eulNHZeSb5nwhOPkUvVOa+VC2bEl6GG53zp1Kvd/lWrChwvISpCEr1IabA/H3R
ROq1WNrcM+iW50CB6xN2BfEWQ2R+75kfbPX/STMW2F3gFKnQDmCch5I+nP9VoFPAAhvE3pFW/uYw
avuYG0lC4Pb2U6aiZ+61+jek+9MuLCGqg8JOsFls5uSKK53VPU0k2I2MvqpMcAYg0jRWli+Y7dxD
I5mWrUjdCu2i/AUxbNDw59FUOLM1l+e5I2K63/KBAPCXVyueR8097KxAJL3dVM2UDJwi7S9XONJW
phLLlWBrT8VrOvJbBD7g0NsePZIbPpNgYr7WT8L1mUT6NNwHrtqU9eXrmRX5GL2m+fgmGTo8kJnl
vuyhaLqcxKIwEBAh3OfM8UfCweBfUfiGCtXPTYF/T3tZfocjZPH5Ldb8wK3ZIaEURpGjQfTuxMin
G5sTIYfqguLjE1NjBI2jEHQ7WH7t++kXRffS/BOeS/kPtq3S1h+lq6dCbyORDXIgFIfADzN375Ka
sq9oIfmr55a71CYCMpOSduQKb11ckFtmyG32fzOlHTuLjFDNTNC8oeSp/8/7pv+0H6vTs8FOxbqZ
bBs2HFIHPMR5XtNyR1ydAJ+IqOQTGo7cvsRT8VbP6KpmGdmCBFIa+dPKN2Fkl5Pg0DbYJsAInSgm
3cwp4EhFkIDO9+IrUKp0M8v0NT1aLGOukfhb/dG3hizydy2t+XmAEdcaHZ9w8TvKCEjbZVqXPSq4
9rF+6NtBgKFQvbxOaLLZo+GUOn2e/ZuOl8Zdtw/PBJgXTq4yTD2nYM3TJI1n43cfmRgxdpHZusy5
pF5mNdSiAJM61T1tHOpMDZSFNPV+46HYK/EQ8nd9IppZGapjurdGnvRWMC1pMpVsvpC8Rqxb/dGV
IBBUAaAKnPyN7TS0ZHIxyhJQbpn7UJju1HGA/Tad9F7GDiMiESr3U8EAPxAh6YRG7VRdtVDDdDaH
YUz6ZvrVSMyHSTinHXV2cawm5XYbOBdPgeWTIU9tjNMm4NXcrrrk+gIgOfcGzpJ2/lczv/IqhFeg
LTtARnZWEatuqIMj0R6o3dE8y74xz3ayUFqVQMPVqGc08VNEA1XZgEveNngkLVsPhzTUeJq3i26E
M8rJvoiK7RjDYus6w8EnDIUuZBRqocL+jw9zT13+1QrV6fUBqOBFXHuwa7Bm55ofbt3cUPeYz6Tt
CsO/AB+expfXl8mu98q92GYZ/kaMkU8UtX2wMU3cxK3CAKLQOoNOvYZX0S1p5xUEqyKI4YG5ytG+
kWfYVKlEIGrMeaHFZ0GvZj+/b1W1mgeyNDpaUIN1WRhClZqUpwTLobEJxd3N9YVVrJi+1qnNMc/0
1ggH0C8V0frC4Hqq3UxllfmL3z0+FH41EVbpfvP79/j3jt2R7e9sybDoRNJumrVUX8r0GLvogeqE
gcuayVdjuoBRb2AgtNDOcnpEOPQVW4JPCWZCd2SKgriNHc9g06Rxn1NwJN3KT8Nv+DkQ0si+nz0i
SVUzfi3cF9flSq2YEsGYW6h00UjWQPtkGUQC9pN+VSsm1SpFKwXZV/n3mCcOgyGccTBZmVzCJE/M
AT60q2r4Txz5DP6rXB1ifMW3gEushtnABSqX9zhbIEQfkSoxFCtKPenPt02Ii1o53mQHXk9zoErE
vXlQVHdIJnqAvGEVizSBsZduEv99YxU8kuRWw049RUJ9f5k931tkrS6Hv+P3Aqb2OXckpHqmDVVY
ed5gqwkVZ6WGGEMGtCcQmgoIgCwW2qiYOEmGRlhQj1W9MHpw4mtYgAdaq8QDcyGkRjYAaf/dPr4j
6adKslqo8N1onHqICOfkdY1dVfrIFMHtZSqaHtoBKztljmp6atQIqZsjBGyHEgtuHLHSiRkdW0r5
wmlGHQ46gsNZTBHFz1JkJz+d/uOouT8fqNz1o6J44s8nzpn8auBZZC8fDQOhTrgtqI2JxwGRhr6N
s9ZiZe2SR1IiGHTvpKcdlV4nHIhcgqZvE4iO0lYBZsk9oJyHf2iAUUVjX8oTdjS8TIRrzJNzTFBY
rE6Ra/sCnh4XBQK7CzTqMHG9WmyjXBgpNhYejhllnP1epL+vfi4z63zo79Rnfv4HltusXvAV9baE
0dUEULnnIEYrWjDUbLkUsriT37b84TZh6ICXkY8ZGfm0TgNBjh8b8nSMDIkMjG804SQ6wKv72eOq
1S+P2U1EpUqKBYt4rc+jGgVKPisLSqt0OjDn9TVJiadoVwHGBjvLvZK88B09mn+xMuAw0I9av1rp
LvVwSuZbF4abJ4dTcIFVMv4ATcVRBuFp9hAE76pV4NvZJIseyZ/uhx7GnG9braMjeMVvb/C76gUB
we3D7ePzlexHsPE+IU7n281XcLzaOosW6AHRyImoXxKHMop7Af57HVd52uiRI2lA6Nxl5uYj+nz0
wytDszIzZYGvM/MdruSLgm0UGNa8K4r7naCybOKzpqmjjqSNy7vGThn8dTA6mnIkmnrMEbIHr9DA
2WBqyN26YI0O1Z4jAZaskDsNQ/EiCQSo80NbExChycRnGwO+shiHyj9F1Kmw6zlc5wcYpoeRI9SL
ISUb7GiUJk2+IXARjgPEMt61rk34sJd1uR4mDlt9X3o5SNUemxGaABxN4dssMyaHW4AEMrp+7y4Y
8GHRMP/gWQBh44UB7hH+JSPdll43hDL4LivU9pla5JYNbujSPy0DEOT9qmrSriVM/WPBv0gk5gNB
SWmz0wd5XvH2hQ6j5mGzo/D8PeJxPKL0miVGlaWeGdvoCxZGZbAZtgt9oC8zmYRkYMJCi7xud2l3
ZtHuyXvf/77EW2HbcVj33yLAZVejDE/prHqxmWsP57ammDydn+MwhnpYTvH84eI0MVay/g4x4Yiy
SN5ieZS3Bl+OQSs40TXEwMGj85lePpt0SI2ma7zao7cPYuztZkygc+jofGBhOQrQooH6Dbz6/RmA
rhiH0p/fEIG6wHYgdOUkz25Yswn7IePUqKIMvJ+z4oJekYKMSHyvMyKExSMKHg83VXWydV77VQho
2iWGr1JtDX7/Va6sBV2lfLZ8apdXuuOD6hDzF+hbw/esqFowTBbWTz/KEB8SdjkUVcSXp3oqACxa
pfRpynsrRwpZdmuZWMGGFrplIUTMYe8W86jty1zBwHo8uzSwckfOQibKG95tnP1nZlyS2f/iG8a8
mhMO882ky1tjzcq3g8lJcpLWIA+ao2Lzmi4hjX+Wm/f1TXZg49qYdCXGje4jIggVWbejFq7+Gywc
zveOm0tBpnTV2X0dyrXjN94uRFUzvLSOxPDGed8h58BEpi0CIA7ZiNMytjlNGKo++dpJvQM1pw38
wtRbhf0DXTmrS3DdzDJuSeeaOV9PMC8/gNQA35qGePhyRDeQQjw2SFGsw6IdbXIgoWajniYIQgIK
iIj+lwpBgS6ip8AYNDl2C6Ea5wUNCH3OL54dqn08DRjaEgjxHyfWCuQdV8x1KThxssN0eWNm0gIo
C1l1Xc7TS4fOrkbdtGaDe4frd0aefRorx0m2vKTwVM1IYA+dI/yu45Sq+XQYUPhqn4iaCfA6YUax
4bhUGQxNVZWPzuTTfi4PBP5kii4WVFm3D4IDPiujma/jbJxNXQ9k1aFQfiPmrLSVSNOTrbzKto9e
ZohsbHsZWeaR7kXIQKBeHGih4m3O/JnsWYniWZec8O8iBxhs+lbzWW4etpHPGKR+kbFANqw++v6f
vLOxiXkbGXiOi0uHIR3oz6gIQoaOLTXhjYl4zhk42hvgCtulNXXmJivwlUqZpwZjG8qX5kxnhNxG
RFWxUKDO9IMakJLNsGNwBMAVKgkb8Sr2oqu5hiI8jdddt4LHBlp3PqHWz5yLtzNoR2X7EVeLbCNO
1Dp+UyVCSjXoCztelW3Dq2l4UoM0sqW9JoQU0PoXYlWysm68QJtd9t57YkXu1dRSnMC29WWwA7fo
WzQa1nDC9KR4Sh/2ye6EHU4FVoMj+caxlBbaSrU1aWC+mcwaLR4qap+r6bD+kn4UKXt22GC76vDG
DydAOyIJkUgRBeXtqPLo/weDEk8hchja2vwKuWx3chvfqB6Fi3W/XBVIJAOy3pVTPrVL/vTY2Lis
yszV2SWpO9w7fOt0ddiFmuTi0B/uGVfJQC4ZhA47VoCWjFk0b9BZ44ufZAh8XIhGw9r8H9yNxMUB
MqGd6DS5DteHajQGFaz1TuNx2UbR60PIn7+XFo36ymkPA0dToV0j6NnaVt+SsIZOgOP5WyyZFLHX
dC5rtqqEz3kL8DYETluKIb26P4HQ9JOdtJpkftb+Mz/tN+MtTTZCSIhf24C5VIHOY4wAPKltpH6b
ubjKtMHSV60m4btGbISy71W6d/farrqQ4cPOjaFcJomtIpc+J5ZsClW0z03z7XZk2crdNQI2c4oQ
AFG+Ii037e7mmQsS5Gz+b4sW/41UphuX3k6c9zN9vwd9u6DAhILeM5zc8G1iBrzICDnNw6cb4Y/+
DnSTJVy2YfddtyT96LTZBsGcmw0cchds3M9vYjPOhBaqFLvPCJHjKEE0yW27JKujGJJr/tXoDybW
uRfNSVNu+sQNJ1LVEqPTFyFFFwMo+qjbNck6vrWpnjcPoyQqWUpDXBgZDh6R/52wyRGaGaXm53yC
jank63ie1ueC+THkkF3Xa0qnFE1Nyf8VEPqJzrnTsLF90dnKal7RGvJ35Nk7t7yUlgbGlGwhCDNn
Jxh2Key0ovYML6v0qu4Tu8+4bSE62WAz1vXsGEF7US8OmkjURBCkZ32vfC+S+Hb0GpOLMsU3mAqL
OyqfHx5cWge/I8zMqcAKh9ZsAmp0jMS1bwIGt3fQDtFGXmbFQmcapvexL1nXWiyvon3tSj6bsPXx
18OLqMhvsszhAHHnuHW3OJkgBXb2yoSlp1aHCM1JJIas7yYk8rqn8HRYjy+a4hVgTLpzjAf+q694
Hf1szQnMhtcwNWk2pSdEAH7TPz751nR18YNMa6+HgazHfEl1Mfn0WHPfFkChgKwGpnCYKmaBWmxN
rGWR9a2dYliigL0msBQFCnjQ/3pvXmRJGuQ52A7bEsSKZqJfKJsO/iD0vrFVWJz9GKHS50Fs8Bs8
QaM3uqRZv7RK2ar+8kTxuCkV6gguCW/tlwMZsvVrGhAiUtZHGNGS38AU7KVWT/1IL8CWPvUVh5fH
DA7vNKzI802UbcJWVxJCaF/opm/4ZWbhOsruZya9xHf+vzTmlyjvllgAWHh9BS3MrC4pTnY1HSBO
kD0id6ED4tqOf55BqgTMIlusB7LkUn++cQvPSVRnBd51TTDGQgczw8yjS9JKF9xDWYFaEIk4gWdv
UCpXj/BS/+lH887WVTaPjMehCLnz/73S7qs4Re1t+UAI/E6aQnRdeL6yPRP5xCvxTnfOzxT/mhKJ
pBoMN9oEuhgQls4EGQHmCk2tlhBUqbauSo3tQlOU+2pYn9QhJKL7YwOIU9rQhNjD+f66Nj17p5KF
ANJOZEhVzm2Tod87fxz97oj8kPGlSPgQ9soE2xBv4zIdEY15MBDMjTx8YjqADBcWrX3/ASI294ga
VbCePDwTn+ofutWF2bT2NxolF1VRJlyaPEIn6gtOSi9j2jSoRHw1vk1onA5VeYRNu9taskcTEgAv
O1JUxODBacSHLKoNzWIvumIYDApU7QmKdVu0wSM7B3LpRUteLrzrQCTi99RMRVXK5Zr5JY2RQA1T
YQc8QQmn+QR4kIf2l/xBKweE1TZjBt5PfGzDfJsrWQTMBSGgpQMZEFht/zvuA9Ew0kF+ObHnRi61
8vyAHIcWNOWrsP+7+gLiPoce5qVuTlcIICVbQLMwKa8wLy5lBYluAMsUAOqbVSj21XVraIzi9EsW
Wj6mPYBkxPG8ZIdeZpa30+s4OG/HIHHw7ZgZ7lA/wsPZ2UDuqlNxB9YPb6UM9OUSaMwPfajXsF7w
s1VvYehJacKRlGwtByXLT+SNibyQuaKZ79jMIqhcBXfUiEI9l9cml+Aq0FTndzzoncoB4mggH/Xn
k1v7hPZ7JKL9Njeh0sFfNtVQS8RbHcO5t7k024dGid7PYrTaV51a4UTnJup/bEAUw2p//HAqVjd7
fKvLJfViptWt4PT6kkFxGE3xBgO+JLAjiqrRdMf/F601SdeLx+DOla9WnIAFKDPfhvBm8OX7gL6w
SyrR9mou1PW2AA3sKTfGexTYkeQQu81OrcEUwtfiHyMWc/OvB2+jNZaid9IhvfX9mwZlX7YqC/09
AUjfa8fpsy/RslcmZW+UPMYzNC6Znnfo74B3rnqzR5wJtPzfcwPWcuzJMEnKjAJ8GOdqc+5Qo2N8
nUmbYqBwmCAYeemHysCYgzpZwryNwLi+eaWYXW+1pTeawXbWx9eITXJg5n2qxUgVJ/noMQUAIH11
4cNUlZ5pIyjwt1yvhOOK3/b95z5ZRVRS+XqWShL+pMnwXy6b5WUKJ/52qsdgmlSZrp7M7twUOsNe
UZSef85dYNKebyP2ODFM70Zh+LuMK9GI2bV7wELFB2LwzF9fT2s5EfEvZh3BMw0PGPTg605X0aqe
ol7QoZCga90pcpBgZ9mRHa+7LGufiSRZPMX/qjS/VE40m5P2L/l8pjvkTIY4i5JewIedx4Q+8C8w
O1AU592CImuM7G/fCm9I3rbgJgzrhBkrZ5q9Vvm+dvIwb1w6r2X94/HkmpgOnPq/ci+je+k6HR5y
iukrIr5IUsYHtbCxXqpJGrnNz9uKnVah2bp7/1c1VadJLcwlJceqAsHUjbTesZyaYPP/CWVQGs7r
qJ4PyLh2WirDulnqZXVGALi59NvLf5OM/TvZjqvD+yqqjxSkTa7vRH/WEjx9qDvySLTWvJ7NsQ1J
uzqLNhpVSaWKLUopAhlJQPr5WK7p+UprsY99tmNHJ73qJnr8pjwTScD+NQ8UXokk2A6HJoQSKu3n
zfJEbGGrQu0I+1jBQpqOY8um9iKk4lFpiGBLPdyw3SgKeyRkG+gw3L0psqq/OkCBzSy+scwOHvN5
cgOG6JxMfuhcdSY8B6wniWL5Nosv07IRe2x2ELqvhpUluG2Mdhb9ulM4vZHoKWkM28vqQXuiZRtj
fcNwSDjjXClmKTunmoawLNfaa8IoGvJ/iM3vzNilEtNE8gwpGBef06mXs+wRAjwkJNjUyIGNKmXe
JZt7NcqDoB0kNpWvMXLpEcn+CiIIHpgWYNr5kBUpmEpjLbo+NIEfoE/BTSpxRD8s31XfXLgEUYJ+
pf7CCjThlklltzyJ1t7ikn5dbbWKSFdVevq74+14VR68vRETW/XtxtM7NvCTbzn3bQDF14k2mZME
mQk3oKhH80Bja31QImae7hWOlxkVhXjPmIIqE6lGulWbKcP/hB2u9VxVGrFwbKgDuNPm7knIUqw0
bFUKVSPijExQkotDut0940AVwS0ne3X66HGn4/r6g4c/2kszjto1N+FNQZruUoTj0p3rwNi4pVqM
Dy0TtpYR68QmIxMjJm/rr6ysCdIJSyRXSifaDTNOXj+p77u7hN0qR8RY+MlQzS8I7D6/tVVa1k3D
8WU6pEtZevScdDg6U9yuHN7eSpmm9587cL0Hp8U4uJthDiDFhjnYxtz5IkyZCH3ci/9c3lmVumdL
I9Ny8hwhflu5FYVa1XGkwoEVoCVV8LF52+At4zMpi4g4Ijbrol/dxBMRE36sGuNlgfOc0Ba+27bY
et7uHGshD91l4utcjEyq2mEcA01B/PKAqWdfYK8OdHTvOdEeUozyKowZ4G2350mnwtA2CuX74Mo5
RPUDkaASJZd8+/Xplfe4GzPOFA1XMQ5SUC+vPL+44fsnWtO9KXbGjRVdLLQdwvuo37pIKJFoZ854
Nl13dCiMGTaWBsYq5CL3zHQYlCfNxb9S1w2H6zsWFBeLwf7Pdgn8l39/DNyoZzvESrjgH6IlbkJ3
2DyT7c0mSgKZUhEZwHPjuaWLTJ8s1x8Sp04NKb+QChNHQ0qLvVC3ohtM+fm2GStQcGXdnOF7dIra
KcHTCU/nJ8sKIaNzglXgcyI7h37KPfzlDIz8krYx1URVoKF7rQc6U9YUm2/OWk+JKiR131IZ+VS9
i/mDvXHitmOzdiuFbWcdv2J0rTmytOmIIcPaOhA9frRVD8LjSUTQ41A8w5pxjMPJNJTlWoFv79WT
NU3pzHpO34IJ5j3RE1AwCveaOxPMloTmpFo3zrzxVInTisNrU8/eACRrPFJOcQ17xXz9bii7QjBr
nXtGu3oZKJQXbnN4PEcTiaMsgOpTYWig6Kbt7qzJuztm7Dh/023UnFR4hKjN3dKe3RHpXjdRnhSO
S81HmNv15FokWSPjN6ptls/ccnGXsttkP6XU8xtF10gCMkp7EnmcEpy8ByMAE6m5k+F2d1z0nXRW
7CIVi69hcUCf33vox+mN3oKWcIz8pi772vLLuLdqjf7paQSwbF0FiAPCpPxYTaJth1fbcKbbU8Ty
0FeRK3MuKiRAUj/68/67TvUgi0e3qdeJPivJukJTG0Og+bTTHDvPbjU3TrXhG3ZFtzBKNkET9uAK
D0YjuCGYlZ+lfuYf3jaIcu7VHWnOuQne28jknLxwZp+Ni15jOnvpn4oLLntckJcG5li2IViTymgZ
bI8x4XkGJc2ye3ni1Y1JIARgTwY2dp0M0wwaWrKplCANST3I4pRRY2w0OVXgfbUo1YuoIrLxHCMs
DF86ANVxq1EPJPcXpLDuzUaXCCRFwU7qks6Z5+bwpLqsfeIImgSTRc6Jug5KxElWBn9Mc/qRDjaw
Nt2bIjG0EnHCdKJnVRIUse8O4Cs3a8G21NCmKXQaYdksJI2z+++TGN6RNfej5J1wzuwEn1t7/7Fp
0luiCpkdKRlktVVe0xVnXLVFsWBXGsF84pSIRHFjRZsPIPfjjaeCqZFpw58U0QXI3rWYe/Xj2gPX
e7gz0f4X/ED2PlniADn5Zyd3ryBcbh49haF75EWE+wVfCZaKkaBSM1GxdYbX95PbRlyO1EEVGkXi
gE4X4Mt/ue6Se691mwfmH7DiwXzJ5X/p+j3bfQbmSh/c5X0MB6Rg5d1JD5414fX6TkCYcz47w0I/
qvSAhXQflUb9scLwESgandWYkdb/dHgIxATG5U2kpLnGyVRXgkIcSYfZ3Fr/0T76BO8K4ROcCo1T
F7HhuV5IyxTM9CpFZ7If/KM7CFBvXLX4/EbVttrS9DDvnS6fwsJoAUO+CAm3+fwcVg9D9eLi3l0z
8G3Md0eRj02GKPv02ttJi1OjCHaXDmC4rrSHU4tZB7NSQB5SRqezUCi17d9zUTnvhl7idic+3G6/
rX/iWMssPiJoXf0goCfxLudjGrn/hDjgiJqrtBN/0FrntfGPsnzZ3A/PLnEY3UjtNk7onIORjuNd
vNDZEfjc0GlH4YsGAwX5PSwvgf9V7kPPlNKrqfn2oMSP+9GobnOT2QTezkuayWAqbTpIGRNvWl8j
xrOxbIe2F8wqMEMq7rzFkAeY1CmFknBedTq1Axyni8Wu/Z64YvtO+JMmqy3Tw+3yjzGtAOWMVvCX
aQ965W51IIfV7QiFYKmytaFBveljerqfRz0+Kot87UUqUkcw6cqYksqt97i/RgJ3zwt53x6x5/PI
Vk34CgVgLTnmb3We+LtfyaxX0dTIBJLi94alIOnsptz7bNWyik5g59JO+AKxV8KXnMwPqdswBt1P
weEVOlhSTdKCpBjbUbB/jc3FWy5II1FwL3ZedUc23QEDfyRkWYQ2jbQBWcPQPPorop6swZfCVZVC
PogmhXLnf5KRSdHwheZMQZEU1HyhsAM7xySbIU/8Zh78dbg/fvNa6H7Q6yv+mOh+lVIoh5JYRdJO
7DpwtiMq69tus9ulKsZTPqOw5b2PlmJQ/cTotgZaPreB+p66hQb6mKz/INKr7R5a8ch48eNTo868
wAkd9OklUcUG9ZuTC2R84VU00aMSiQhnaoMYVGNvD3yfX3WLCjB1VxCPjYWamz3l0aMQpvYHPWPc
pg3xMWQPTlsnSOyP5wgX1zJNWpjAwL4aQ5PP7brFb25ayy+gv3CGitM5sQvzkJKQIyE9lIWmozSq
lFLV/yuD1WXvoeg43A6N7YIT3ebpdbVNvdKN1l/umP+dC3eVtY2ivS7VNex4P3NU5NttgSfOrkLA
su0dQExK2UYI54APJ2R4NofkApzuqaaMu3KPjKCuexLI7x+JbIjbvZItyzDw9lTb6QcFqafYXUBw
RhRXsi0ATL3G/NyDFRNeX6LxWynSSCRgtc0qisWIYOGqfxiF6Uhl22Q78Abg026tsaZBJZAwE+6u
PbnQYXLi/p2axZSj7Tof2puXGFl76ldR/nGyjjJw+XN71gYs4uuNtdto0F4iVsnp6vTqm6O6egAQ
e3cn5zAtyYLxcs+jHgVIqbi4k7OunkmQZQjJZpz1TsCqsJ9U+6mgOgeoNZWaGWrnIl+JJIrIKHq1
8aNFGVh/DlcIcvj9RqBx0V+sRDJW9a9+MfGRvnt+FvvqhjQqP3nlnbMhb1IGsqgh402zwgNhEIHw
4VJu+TZlkjG3JqSka7SZNSvigl3Oy5Rh6oMs8Jc5kZD8jlmtHzT3QtT1Lqtt2BA3Pv6zgSkQFNcM
qK95ZsDg9WQ5P02ig7aJAKzHIUUdKY64Re09/7IXyPPtCgRQ18FOxpDIoIJTHL3MOZXo2d0AdirP
gcg2MAYqpastEQw/LoaQw+8gmww0f/d4bbo6pw8R1wdn3q49ENf/40RDikAMVzAPa8pWqIJZpsKf
3MQEbvkRLYn0ir2a9xFqlGc5I3UBq4Ui/N0ci5+cFc46Ywf/HSinpGd2B99yD5Rs2t7BSzRviVbf
KKdJFp7i1qY5IhNi7j994nIFkDqkiTy7nMYxetJjBDyLjfz/dn5xHY1/W910/NUkM3tRlE5mSzyn
HkYpH7Ptmshzk1eURiuXjsMceJdHKvqRVz9KpCpZC6xAgiwy/hkZy5LwKtOzZLi7dARIoovrO7RJ
VqOv/e4rI7vjq3Vsp5g1xbXKbCbEjOuhtQL2g6sG3qwkgB3nuIS+WJrcUYG/nrQrHAd3TMtxuHQp
N3USkYYUq406nQtkmf4+tapbFKE/XsZ/5RKiB6GZrZXK6LiSPz0mUDzvkcWLaDBZeSvAlnoqLMNL
dQkMHCTsWgsJyrsc9rcCHHNVYGb5X6IUTCH73NwMaz79jgbNZt8/zRhAIe2IkEu+YA4ox+sv1fEm
WU83mF5SoS6GtoiJhTP+//wmpuEh7AOb8uQdQw6QVfDG4yaNIHmR7lmOSHPW1TQiKSN6dayJJB/d
TquU5s/rAQFzOSEuOYUb/WMIExUjJlquezcqzWuyQiRxDGyDKJ8xmUnyNswWbHTW46TEssbuO7Bn
R/hQvb8RSNydijMixzycTnxZFs2ewPdqsJMpcMS4hZxdz1AQz4F/km2KgrpyuskDYzyBwyZbArdl
qLYjBw0D4aUQHlBBcRMPcyoqZzhAHBRgN/OOB9JJAtZyTkiqsxHPB9ARs8I+cQ/aMJR2jYYKu/Rq
eY3PDgsP5Q3qEE/gZWb56lymLQZK8VmJka8cwc9ICK1EwAliTepiuk4L94DvYvkLijyfQA/yFuCU
+SuXkKEEgPW7z/R2cyoXz8eWobGp4UPDZ7/ijllU4bTEw+ODbGHpten0Ukdz7b9YF164hI9Frjym
zSn6wZwwEFQn0Yieiyi6pnViDJWjlOJ1hM89BK02WXUe9jkdlysSc1GSe/1ool6J4Ehl9yfAvgVm
SF4AhpmHPHjfgNwDs+6ClFzVDe2axg8IJzHDNhQWNb/HeYVB/q0dX+MYA6Ra7Nz09itlz4Mj+vKZ
275JadIbmV8muiuy39cygjSzi431woP/PX+L2fCcuzQyvEO8S61N23kp0qEGfkLak5YeUmlndeHG
YYnQTjAM3WpLAlzY1syRQ6jz3ZR6y190ezpdcSiEVwbd7wj+YZEW84dqY/4kNxh0UGn0LiwnSgFX
KD/POUh2n69rRYDWUI65yfH8+w+fzRc9TWVKxO4ALIuFpIn/f0XrqUjktybKJsEKBLZZ1KFAhbit
ogGvxcYSWu0X5QHLR9vPaJ/JX0aCjmGx/NqnCzPMRqiJ54vQKNY5pWzDJM/P+zngum26a6KsY9W4
ZLT2oUbJ20LoXXm3ky6hoPYr7teQSKH7d7Dc3BuyeSUu82BCKeL/UQn78yc72s2whNj2yOgSA7mf
e8rYisDLGlaA6jqtQj6RH3yPMD6ZKK3Lw8xHjXF4WSPstLeGfsl1v7at7fIBT0MwVWPTtoXTHW3N
U3DdQBOwaBHnGeBxKpnjXGl1AhSysJU9ytwbFlti23qtzVj0eIOriSzsfUJDWcN5zDv8RwCwBgJb
jO4SzWGELISpcnytOjguj7BOsbp/jOmlU2VkF4nnA6jjPhiu/bThNVbMs491ODgR2b4maSozAnhd
MJZ5aNCNY5bGpJuA1T3blx5iVtxTDiflf/az+TSHEnIuWxQjrep31VtzjZEyCgB5fkMeHMrRF3/5
+s4BMUoBBDgegQc3gGDDIHpnTIIgvY0ORZch9SuDfo9Ao5mpFND3htsz5GSkiwA0WerkZplFhvHP
rWCgCxmdFXU/7Axje8ervephLr4e+61c6CgrUkuBuAw/l4iJIyFtGSgiJkij2XF4wrMUYvwPd/rR
PLQTDsC1emN3XhbsHVOJB+kTQQw4+P7GvF+HLoY61f7x5hLRj+eQ3l3xtGcNmbN/7WxtovQkRJxW
/DUVQI0y8AMW2gauPDEMM7XEDEzEgsPBJuAbuBubvGJLRbNnYOOzZpwMjxgnqtXx9flvK+axKl4E
RwCA7dS5pIGfGS4JQJwhC/FzynFm2wrNMi99Bi7u/7jrksloEJ3GeudkjAG815tEmPIjfp+TLXcG
c1Zx2hVKy244uRUhGKWxVvcne9eCzw9oQqNfPPsGhagVI4/u1UXnULkvhlcXbJpZ17dvrsZgODO6
GM/UEblGYWy8+li97bYMyxrC9aPJkmtPEFyJSBBuJU9PkoeD7h4v+VkWSFPzTv+hr+EfwOPgpmy1
5QWveiQvcKVSS/DRaqlvEDi3xNth0RGo4W7ylXG4uEjK+VyVCr7RabuHKEUmlHbijR8bJYIL9HJa
xAV9iJPTZ4x9okXexX6CGSr23wX74zccVewyD8uiWlLpS5zFQmHFySldwmiwkIbFgOIXbquaIyii
ngc6gB0Sf4zryRxZnylEKYxyxT2/KiIDTCUrbLIyf2odGVoQ+IWDjB7MQk2ybi2XvTxJ6IrmicQt
K8q73S62oZYZcJ2/C4wJU1i7v23CEoPCJriJOTUt1vPqlC/Ezh1HlPLQmQFM7+IOlxmT4Taspl2g
D34jASyfb7o6vHRoCaN/Rb164Z0HkcIveOIGgPEQCLbdB7TnFfjQ9tGijyjazFp1Y3GyAG3LB3/+
9rCtsbMsEFZek+8fsH0S1+DjoQMl0o9ezzC9EtK5JM1bEwzmRGmhAlIUIziFkIvoGbNZxcXfpmud
E3mV6XyWsYOLcvO9fhtMaD9M234bxO/EKxlhdrTjrg48v01DsJKdLv7rYNRa8CtxkBtg3tdDTbUh
HnWE1Pt7xz2YNWcEmzsJzpVJWcW4vlJmjKaa0iIBWk9z+1LD1CEBqnz8HES4QeeFzzsVSL7wMJO6
iVg4lE3nqbLuswc1PHUTv0PbL9R66EzX4MH96qaJ+VLIHXqjpw8/HcFEr9P7Zk+IbFhJerzgxVNv
fxr8DbIlV78cT8cnrCLNkf5d6uD63j4sNxhFGN4ohcOvwA92EGllfvOkSv59l8NSPe0CQZ7HfJ3h
cBQlaBcqjI6re0dOeKFv3izRAfQ3HpBFzyso7jQ3tmfOBmVc/k9CHOxiHuMJYUsy9cnaORM8nZYU
7VNB3/NOSuQX55xqN9/hzVlQYwYN5UZg325OITpJ3SOAvsgpAlJv39kO4VJCNTqD9zDtCRpIRdxK
IFNNjuQCABQZhBPYsqgBVqKk7Y8a30XPxoVZwH1UpRFrlOUtm/mKrXcRYiOXzp1d76Z1TGwEKVdn
74kUscU3WFABfdl/Xm0uATOw7yOQ6qYehRCQbABmAMF1jnmPSMDziJKp4pecIJTR6JrDGotfNmgz
U/mJfB7zKs0ZGxQKKhbNACJETgPar6Hlx9m96mMQvJPBlUnzSvqpNTNcgycJZwbr7990IblyUHDb
R05ei5S9eNTtqACyQjdz09InqZg5BE7ibMeZ+QboxauLiQdYTz6qdiNPqwFLxmkR61HqJ196y4Up
d0UjHnnpRw2V5TXnCSaCS5uVvaKaB4qdhHIp4tuUpfFNSClcCv6VXQE73fhOph5zfqgM/qWErI5o
np0qVTBu3CS86eJy9mJ1XVySlPjGO+RxEn6IeYO8g1aDqcvYyjnuGtwDRkwf+wdxgSrVbY/jLucA
tFYpJuO+SZ8pmFNaxZU3HauiXs0oU32NFuxxUertfSGQGWB0Webvy6PnMQxREV0GXpoRSXzB7Hag
EDqA3gjowqZw1nQGlLC42gPmtkUUPsb9s1aGSoWXz+CQAitA2Qw1OKFCqoNT6o0g9eSi9q0nwL+H
kyQBMh5OIjQyLiSFy2YKBiDiHj7n1NkziMltP03RUoD1JV/PaRVboW8elRJzerzRwnVcvpBKEF+1
xDVZwmxLZC0I4N7w6iu+y1lSGmPvO/XkvH3XtYlZPnTgStLeq09mAmTuuniBDrfhCfzJsKoKhjS/
30Qd5QFYJF0ePnM6CfHnjckmxVl1rLrUOSuqineEqMYmRKe6iMf7DiU0BnuoVjg1/Wyncx3oV6Z9
IkYEqDVjOARfMb6fqQeiXl8ex5rDk8rmK3Hh3jRaoF+BdbjviIIypc+DJjpmBB+XiU2sDC1ZzrKq
THpLvlVWNC9ePXmXpTcmFrTSZcKPcQLGUHcuMPaYFATVA+fFhu+22zamsub71GwE9Lp3Ru53TAsg
lrr3r5/03D8FgNh/2rBEnhOuNSrnR38yoFoBCh5Q7hZI/YPd7LsFjN4SRT9GsZtZ5lfCUDRQqGJx
gI7yl8p0+CAsWEActAh5qVTL+wHJC40D2QGPGmHrNV3HoZ/0zzjF6vuJDGOP+ec8FvhNFQ4U1NzJ
aZvXZE/0Qrf1URJcyCky+PkQ49/Z2/Vz6t3TEyICw3NppN1LqNT4Te7F78+ibNKWPCEwlYkE6FTi
ohN8dAER4tWOzCWLSn/wfY49RMM0LQPBwJJQ58lo5ydABeX2r+CoiquVxG711A8/c/WA2HfELImt
NpXipj6qQpDNi+OGlDbkJbmL1D9QnmAPiVzDF7Q0nTV6sI17yuJixguvFBQXyGCcEFG9mDvH3myh
WePDLnvsAaNlAwAixCMQ/wWzMigg4HEzwJPlnXu61aftYD1hKEkooSfRTESDiKQ+FwYbepIKCwT4
urXksyFyec3JoPvkk7SoNir1Knq0f2qU7R0gwvD2BlMC7OoOI/BTFMlSMvbjE2Cy5f8+JT9I+C/u
LJOc8/CUA7Jd2GvRsDgNUhzW5WViwkZFlS9NsWtwfitXYu/tYS0zzdmqMAwiJaIcYsPtQTxGVrth
HTU48OsgR2JGFJfj/kURpusqyXxCi0LJIeOAruC2kV47zO3nvQggUfVz5fWJkRBtOkiiZdVCGRDi
0B57xdMQL+7AvZDqbHiDNOT0IGQyjjw0l38cgbr7XY2P0u+AgXFYwxW5CshVM9UF1dT2RkKreumd
1J4Ciqez3Gpq+HlBiu4RkJxGC98walAhGOhsophhQZESgSHZ2v36iE9MZt7mh51KPB4hSv7n66fE
tRNo/NFRzeKHvh1WbFrEaBvu7DFIAkDopp89iXkn2hFcygG95UAlaCcER8BD2tqc3uokrfycuaNA
l6cVJkZJczv+Y8WKtGzJ9ex3RVHMWHJ/GiMl6tbrDgxAW/olm1AEsyhH73brVAPLZbFKNfvX+ICk
KBnNyi+gt8x7wNH6Q4NwZoiD5Ko0yWIAFzKd3dzsc3gcsclUQ4ZqRgfMlIPHxpFnRR+3GRSAXk+v
f+GtFNxh/CCZ5m0HGGk3aqjhRCaIUV8e6kAlKoPHwuSMRJ25pg+bt42gnZwsjtFjS2kKm6mHlD/Z
iIVA6PnYZbCpQg/5yDlHiPTaNTr2eR/foyk8VJv0ioOcY/qqf2uNMGgrr1nPqV/Z8TItJIqC3/e+
5SLC0MFS+OZDkQrxN6YAUzo+WFxvSaa4DFbuonKUpp3puAWcChHov/V78zFO+Y9ORptD7ytZLgWh
tpn7OIExwX107EfxqNzVVYHOMVew9b5LDebTYK6aS2XKyj1u738TmUrTJfaos6NZdf0eT01+i5/k
mu/pKOfw70zLorJu29AKwFFd08RiqC3DhET+gaVYkuV1EEmxJVxyXmmt6PdW3SKSE2INDJIVLbkK
rCxU3i6A4hy22OzQAis7gskdL/okGlMXL3DkYq2v6SrfTv66qf3hSHJpPDvtxuENxEQ7FXTKogu7
7n+yNcdtHyH0OtsDOr5g6mnnn/ydeAsJ6GgjRHmrfVHYRGz2RMCO1bJXquRQsWOzJBV9EQ0ip2A0
62Isv87k0Gdo26fWiQvHtDknLTtrZIFTKbXWU2U/FGAmSco16/9XzSd3wP47GpbmC6h9stIMpuF0
Ut1wJG/BfG4uH7MWmg85dNij0vGPkzUifRg9bOog+KmEw48Af7BC7sxnhTh0p7+xZ3kIFg44cHvR
MDv4AxNIjyjb2qBY8qmnz62vVIoBOCj1iaUuW6PI5ZaozsRamNjSOgShJ22N70faJB2pVIfqBaqV
V8ib29yllvwyDlMYo/nrabwxXhyIEWiR3BlbJQwk4PgVyc72X041gxhI+LFCE9MaxfdiqkJSLOgx
lYoUi+UtaaSB4qHl0IArETo8bC2BMhbCcVEO5OFuKVEbOIJ9zBoZbvHGnLCaF+3ii/eUE/Qf8JD7
CWzl6wAR5TWhFHmLv8EMiTr3mhcbAaEY9YJLnETdnpWsvy+6ehEnpBRTLeaVGKDilLhCuaCyIl+T
fTl6SAaTqctiqQJtVYgKN0DQqiiDpUf2O7Uo+FqxHvmV1AvKJWviaBBJNpxj+dkCqILcKddEVIEw
+20A7f7+y5qscyJtCkaJh41BQre+2/8wlJymPgYHood44xxyOHlMsduNaz5kklxIVGOMX4HG5GhV
xCbFEaVU1nWuQmaFll4MftYPwtZWkaO/iMmE+3kFRvk9QzcOFLbePoEsB77DzYBmblLKtIZ+q/xd
zVOKNpdKVdmcMZrEuKL8GLDKvABeHRbSoJeX8g1s++DNqbf3fGOMd00vdNERyWffoZjUd47asoZ7
wEnKuoBAvODjbYBWl2plAO7kksip2zCM5+u8PrMDe6r5iULoN9JCytfSwJLROn2W/JU4NXhmM/65
LMo7brtQ+tXqGgu+hmF3Pg+AEwUxwIwM7GHrma5cfTD6pKtE2uc++B5LoHcao9fi3EgjnZJ87Tax
D3dT5CRFylX4vqQBA+PrEyjrRmABpUk4DGgkBJQnbcK/KJ1wqXmza2odSBhTU4ZfMNjir+tf3KeX
LRNNliJnYxbUo0ftBZd9SZ65QYaBO21Jbyz/G7ROSsDKu/I+vRJrgvwOqkeriETXYC5L0rzLONze
JkXt1at+uZCNsiDXGOJ2GoHOx8YwyDPXz59JffGI83ZLDzY4JHOA2mJXzOCT1MXFF+zVT8kHj9q4
/btimxEveUyZiGYxgetM1ooOKdbKdEPTJFdWicMT4TcTUdC5RZUeDSm0DOi4CWaJctq/z2B0JmfQ
PBjbuUQMCz6LZPomxd1rKNG0lr271V31QZYYg0m/E9ko6X06oCzrPmrWRgRZydW5BooNa6WzinXZ
IJgNQuqEOfh97u3pwMiqpg1ZMAmkx1dzcR6s6q/wIs7DPE0JLd3ggVCoktWvEPdAQsdYCkLrjiIq
gFuAeuNx36YBMtuW2tdKAgVsJwekaVgeA+6U/VNwZa+FLMOSyj73qzE5k6FEIvUbsf224BQnPrG6
gMin/Ktq7FLcGE2+XLRZLqvfSPqd5Ru5dS5XmBLDncv3m6bD4y/mUwFcJ8Uhbp+eHLPNFFO9nEvz
oNPzFteuuNKiBvlorRS/fdbYkfKQNJ7pHzlK1GSN2/Z0M6cyXD8T3NZN2H2+mxN2gvS1fFtrGNUy
AXIUBCI/yMHQkAKW1oXGWt/KQRangE0fvYWhRelsyK3i2X1V1pqpx4KgGhKKogX0y7py9HPrBdAS
801mDsYl2tSRamjIVw8hx41qnlrXX6eBZvuklTumFcoB2wktRTnRgPza4fJ77XcyGdI+HR3xpPM/
g0QIj2XgBFhEdOsRcDR4s7m6xg2MTJt2MaBRnPJNcW2xPioSONUMen8yYgI8pNf5X5QeOxjWwlQ6
dqVXz8L8/ESrqK6MgoygMJ3nwpwi3AEdozLMbTABlb44a3w79onfHYOG1zdI1he86sNo/QjmhF0s
MG1wg9atHFGUHm1NZJRd6r+iJQ6FimmCPFc3UOZxiYgCjbf8fjySUZKTcgy3sNCzD8KbeFRUOXAK
sNP21Ife3flM6rsEJuMmfwhil9QJpo+fOpaEPsgdi+6G+LoO6NcX7rphgZinRZdXiR0otkU4yZbH
Pnn6H49PbJCd0mkSr1DLdQk0sSkQnxZV68Fh+NBlP9KFuCTGUgo9OlAo0YUlgqpoUGuzaWWU4PVc
1JIwwuvZAKcn5JmZkHQAEQPCEafu3pn4pcRSwu2DTsGKWz+AP6xfEs7/3Lt4F6leaJm0nlgG48ts
/L0rmCpc6dEuRNtsAiTpZnWJW2OPvbPUCyAmVZZW4cJVSMX2lRSk4CqD/byVM7iufEQPA7XC5kV7
Y8Yvx/dtq01cCSgvleVSEggg89w4SDAyXfwmTQzbKclC/uGM95eoEkA1KlVxPwMt9xiDrh1QirQW
DG8rFkOIT9Ppv/khjFPL2I9trs+EFCCT1VpYRqr6qrqvnUFumr/jbdp7DzgOM+2PAYtXCs13x5UI
Om72TOGHgxn4Pb5+BHUqYKG5oBQEgnd12tLM5Hte4JWY4cJIdKSjEJ1aYaCuP9MSth2SGC140EM5
VJnEA9rx7aTlbNHX0xhtxEAHqj3cASEUTRxaVitV4dEUKpkKuSKOm5EbelSr0bCtlP675lnyJe4f
gRztPYNxKn3aoWRe/LvAxyZEdqMS4deL23zkt0IwBxN9+q7vpe6td1FL/GwbM/0cKTyJ/NG00Yd1
hy7wojQd53ptzYjmclPa8izKHXfRZChxWHThx2fvSliq6PFkYmiMBYsMCzwicbH2VBK+qTRhN/QV
DdwnKZ+aEDo8yQNv2Ugo6SHfXnB/D9GNKQsz1N9QccZSsiJR5xmiIA8WOeeBV5stxE+hRbDnz9Ml
PHzYg5ByQuXBXKdKIfUapoy254JC66T7vJRk9pOiB5dTlLXfIHCcYZJkbvpnbYeXc4yd/vbexw7b
R3jefwB6fNqsY6QPxJxVikdfY3qjuHQr9e/iu0rtiZ9e0BtVCCCZdDvnlnyvZAtA/9Le9R7CJLfC
4VAwjQm05FhLAqthXO61rYhw3VXUR8QgWrSDKtytQFt4Oak0kn25QIXuvDrrHogw4rV7LlE9YU5Q
mLjpIMTwzruzWdRefRX45Ep+38wDlMK8kU90JCzK9kFq49oGrCuhP93Jb3eImEBwQlZ5ELO5kWto
s92Z4BSYWU6yO44SpxOjJUGOrWRoVVMMCu6X1TiHaBpyfE+jSM42ITaGeyAs0P8wFNCUnSHR8sKB
HgALkNxWbOWiEDLYz/W2QpWv4jdbpAvzzu2yLcL1Tbg+K2aP57Usyjg20N6nY/w2+sgV5D+CCmU1
dQQb96n/kTrNnkVG9yTXYfD7YVvIkhc6grjf/8kcjdDiIuK0IzP8INK2YbUTskGszhdvQHnMvuMu
NfZFaK1Z+/BGFruLUzp2WCKDuvWRer9PlvxZxY7M0yPLmzbcxT19c5qxjMvem7ezvHSz0R5MD8z1
7bdalHfF+btnycFb71dCAv384Dn9fV6I0kkimgVSg8ZRXKs428gvGi5fkADkU27QP0/1bmA+ofMN
dDjiNsX+b7j3+YeJsQN7LoanRRBA5PrDtcRXfmA7I893e2wKtutu2IsX0WFuBqoIiymtB3/ojGhL
TKIig9UBgtWU4i6OiqQ/3Abt4P2KszOXnmfQeEB8Oc98wKZ+LxYwyY7bSYCCBflbL/hd/mNgq2fP
tWgt9ZkBBnTmbc5Sz82BIiDbk5cHYqc8myXfRGEmx3NdhSFa1nOmlAmQzuGCekRtdO+aJRVPr4iT
AtKcv4JDYpao1at0ExKkA/HhXKnkAi6rH/DIAKrzjKNfOSP+dwHGSbaCafkk7Ye8BYHqOH4gpyir
pMlDbWjM+BMM3IA/DO9ZBBDrXPZ6fbPFo5R706TX5Tpg8ffAoBTdAwf7AL6O0QZGfuhqtnVChGOy
F4CTqoEUzSXK/Rbk0xRvRfrh9rBVyp2VBGbuQQ8VlWIKJ5ERc+zgzXsPhA79zBGqfpTbhhZJhDUc
zzVEsPjaRpv6iByCHqHFN1hj06kZEjLvJjfA3KxMe6LY7KFwu/8w2F1aWZ72QODi/w+cNHwqXLXb
WXgpiFYofQOCrbJnsRvW/TTtPZLiEuP4sAifRFr8IH7YxQ+Wdwggwc+xHrmm2b9o6xVQqvTQrYNC
gkAXxWMkILcvucNA1SPzR1U2etcvVbxC2KMAp49pkdhDmQj4S7gIymycgL4s1c7vRyL0KkoIj2Or
OBc9AxqHEChlyXprEZ74dQg/PImp3dAbGmypAoSYd7ONrp1RzJtRfghUJ0hzSQDIQlB+8TW1jdmj
+t5c2RRfCMewn2Sz9kl8YzhjmX9aYER3sWhsWhugEcP+XN9OTJbw2jCFy3j0w6fHIFGzM6dR9Kjl
TSP9XEgSkUY/G5UF+AOoC6NaZlWk0JAv+Ay085IqsYjIsFM4e4hY1WIc4j1n/3eewXXDDIrxSszV
Cw9kRaCLf+8VKAruli7sN5edO1+Hpez+rKQqI0sBiAajcOW+8JoyGATC5bgPZZGrb+Oj0fuv6Xny
ETMSlnVXuNv09dtDsLZr17cjz9nNvA8xmA2VqdNpLgMKATdL8sVJdENSfWjY6VUl0eFp8pBy3b2E
A3p3SIniydWTljIweT8i769VyaKbS3XwDE2SW+By6q4Upn8wKVKuMdrpNLm/+4OXh4BDvpBV+YzJ
f/yNFOxH0hGfJoAF7wB3S1Zf8DUwh60K57xMui9VdPho5hC0wMTPnaeGj8lwwlh3IGRw+Ibi9rra
cD5anAQCZkTJNcuxI5MurPE2nZzh+1P3p0Y4V7cyjDLhkRqEgs9nFoa7wS1jzmZbrjEfSXyQ/pjF
nl+2AG1OlZs37VBXSoearLLNyPKWaAxpQ1MqtC1I08bzvLM9P+q5+iKWKDPPWlQAf1HIw2Y5t/3l
UvM0kMtPruB8+LRFyL8gf680sMh9G7u6AUxY596Qs09Y83MWCeWAMp4Hn5dWpJKqlqVZD78XOmeM
a8/DekPrhZFt3LR64RPdm0oA1CVBfqD25qslSqz2c/sL082eTNoL7O+r0Jdr2xqRm/Dgy72agqbL
t10iYMLVGRB1qBT2M1CcytABVIozd2BW98DXqoaAgSvC/gQnCRJLAjnIXVVjvd0gWYJI2BPyyKSZ
JMqNkQu78HvZn8uDAczhnamPA5W28ijG3Z94y6NKANx767fHEhPZEkhAbKXrW1QnBY70EUNT4PlP
vw81ttgqqd6JepIjtkQ61y+H0xK0lLdWTkck7PlV96X27hmEHhDMdpYbcEci1bDkxPh30d44nkBS
CEYr++Z8y0QtMYztD6MKWMvb2wJmpCWKlQgarfgKmKDey/a0Sd0SXkZX63F83jNHvlOJJzc574bZ
IS4LSaXaHw6qkDGVYcJ8tXkjn/y0yWVHWCnKcH1iA3QmTa04lxUNmTexKM4CqSABB1EFsePsKpSn
b8cnS4QcOkixJ28PJ2YV6MSpsJ0S0eDjD8TgoqjbhzgYCksFPgaCBc86mINu3mD3A+DboE/u0s2Z
WnSpSOGITO58v3M3oxQsHbCvl5c2yVjdEKsbq+8k1g1vOQTZaAW3AfmK6k0dGdpjm84ddjbnnw/D
JiCgEgpy6D5VMeKne9NcEGJKRaj6mu4Wik2xs47Xak0+QojewI5RIc0mNy6HukjJrid9Xm3QuXMv
h3gTC5FlD/GLO0ILel6BjSWlJRbVeRmretZmh+qteR6cJ4xtJhWOBGPOIvrECNQeAiOYz8nNrheI
LLQNihZJbY40V0A5dRKlMa7Gm+2wrDZ9Bc98jQi/dos0FovJeNv+fZVz2rmeKO0L/cQXX9fVDRI9
CtNSmfqY7wn36A6GlMJb8JzdDTjT6FbtDKVIMhcahvMyQfDfCLwHP6Hf634d5BmC8B+3citFXmzw
jdJw1DFrdTGBG2/HbqycLucNUaCWsceFoPioGg1g4kKISEE5XEf2op5VnyWjERW7dk3rAJe8ovix
BCp5hhK5Nn2KW12yWmeRtYLN0i+VNyjeMUtyrEHTGjB+84540dUUvtXgv37l2cgSHVmkMnqzeHxg
A+SmEaq9DBb4fAkBNzp3dcHVI1I38jLc6U8fWWyp49yNjo4UJj4D2HtdAiG7jz6oCEkSpiwR30rx
od3AfJifBIl95o58qkJHoyc3vfKRhU5IbQ+vwk8H8jbItB2q00G1QOXk+hG1HnCw2rAkTd3DdI/J
w8CunUUCr+saAKKrD7QKARvEcRUwizPxzG70xPtOgPrQNhF3cqhBOt2rthJ8m7FPFMFvZYq5VAMg
Ok3/fEgUSGuRQloXSNzqQ2PCg32X3Ys62sIFuLySRaIyzbChV141pS/NuGwU3y4WZGBS841Lo2E0
gxl8HGC/X99uJobW8yRLChpraRGEjFaq4KJ0bFCYQLXabvtgMzqoN3zTMuf0Mwx5pg+3C2hRbpoc
70vZdSV/Gm4ewabioyIccOkKxy8xwGBVRzOLyXq5uFerZPxH9tO2g7l0WC3xZLm0jXfQmwf4gk8x
h+JhoZyxyvclc2NnAAjdBUsijwvKCb2dyHIT8utqepy0/onwFAiPj9wXgJAK1/snxSr/71RuEare
RWkR4s9J9gvBEHW4jIWXCgTI0Y16xMhzS4aWGVp53SybN3W8TMa7CuYBIJ78/YmHVyBiuvhRSaBY
5Ep6tw2aJ/pBUFt4ttIHAVPgzLKmM+kCRnW7ygP6S9ESbchw3RvFFAMPgGNmCIDCaWGKWaGr8cxj
cY4Ii3zzpaQ7p1rVdKfpY9qz8Y+mqK7F8M7xZO7RnMiNzrCh4C3pM5lUo9z1xLfRSUmKGKzOx/MS
bQ6qb9GGClM0NL+dMX2ifHBbGINjOnpkraPkeO2XON9gQq1FeA07NaoVCKrwWvyVwBRzU9Qvbyot
LM+RT3sgd7MRukqCWtdOZIPdj/PHco3JFoYtwbVcVUPI+1tZ+WMUyHKpkM+voXyVBuK320F2XyGk
54RRknsHHGUiVUZXeNvlFauz4jhR7A0pEtMZwhKc+q/tsv9k13Y31oQ5psQSI+bMPCsLaCYLltsV
lJipgGLKVeUTQi9NzB8HDn2yKkHJLcN0jtO9QeLAJ7946j8Wq7po30hdhJvTWW8F04ljcrHxx+FW
Ou8C56V8hc4WOrwd7oV7N6GiGxeIXPYrC+Q+FnKt3CvOYY4OaKXodOoAG0siLpMkzCPyfbDbUUHP
wueB4MAs+BDWPYHk0mXN8rl3ssGb8sict/JYHNk5xpaptIPIXAl6BCV38z51Zxs5GOvyfPPB78OI
NIUpz135wLRq9bWuXOydXGwKP2LoiQOw4IKnZPPSxOu/yB3cFqiSs6ahh+D618D09WlH8lMD7jxP
V6p3cJNFiJ0isPjzrS4/WMnn+mB0qa1jQG7UQ/+IrBjW2Wc5s42tGSlrZocwHYCGvIMywx8TezrX
0wKu0FMXTQ4jStj4MYDFCn+lbkKGF84Wy5vzn0sMRk0322vHxoWR0ilyHJZ/3eGcNOA7N4AJK9cg
qkTvFC9ZRlQ3DqVagTlIj8Z2ihoHtAoVF5oOP8gzpI2lXFPhsSgVWqTORRfbAW2T+rNA1X1fSkVI
NFZx4UHGdnsSCe7ZHwqRgt5vClsm5OMu4eHuyjy5kKTfNIlunpD0kPMk3QO+CNJ/27m7E5fDa/8M
CLCh3W3IhkuAjTlan/yydgWUK4hJfCC9cZBSAG0dEzUuwcGLeLq44PWpVHdJkWhNlmcTxYRqisaa
GT82dsFhM1usx+siwGNDl4P95+juyGjZ5TlYFDCyaSj89cLOmS0mprCt6Vyc8SisqDtJcTQdl0bj
Lzn3SdEmNrLtEtovvIta+YKPI/lqdSqjjxb0MFxfs2BNo8ENiKjCv8pM7W/lCKeUC6u/d3FESQ4X
KWV6eGW6aN7eLQ5p4ifFEYKwa7NZNoDGa++qIe3I8P05qoVBTxKYrSjkzEOlC4JG6P24fwzG1f3X
N8gU2ZbG+vDZXGE+ymRn3HFDz4814Dj8iV0RX+DyOpWd/1y+QhsphhtmYJLpwS1wmciYGMZ7HYBt
xZgbQBOONkcA679XuTqgVL+6LH3+kKRMV1ADxwaf+61TRsJm3eqZ84NAoXQODAierAS/LXZ/WbQU
rkW/YB7lkTCgYlFrkGf9G2WCzvuVhEyeiDH18ggX2QPdtGNSHGeapAiOpipO4CJFOjX0wIwK/QId
8ON7/vvF39PO5O/E/AW437jYrDU8XZ/9YZmTls2ZXV7L54bGZlYx4i8mx2j10SIpTCEa227WyGq0
BoS1WbJbP+loaD9QtFkHCAPfrKd1Df1mYv0b/OytAM16CQhCPOfHoVpH47V/VXSoyP53CG0mMYi2
vJrC8t5LpbciGWwef77CgfRtKuyKfj3sWBy9hr+0RfKwL848Qjm/w5z364XDHc3XdQXsvaKYhYPb
IiwTAyKNHs8w+1BS8eUxV+AQbN0RjOadwoZ5JpSVURo2ZM2WzpAy3zmhsV+A+fNSqNQCG2KzS9LJ
VFp9st8/0GM4itK3OxBHa2YWSR8ydTJ03xnchurG8cpLfFfYdc0Im61MS2qhkCBqBVBlEtT2teR7
3KdVrGqoMhnU1PF7mP5t6BGeFH8M/uD1zLmS+CW7X5DqopTrzk45GUYTuFPYkJa9KppQ0TSeBGN5
YcP7UWiisXM3ia2cA1Y+hEizP9/7Rui78GwiWpCvqTYomEubAG5yXTv/2QLXsdgrO9BRG8apL5do
ayMkxpdgUUpsJZC/WMzOhzSo4HQdHUUsHjccEThOUjHyr2OcUyBjaw5Hbyj72sUgd3ORB2qTZUGD
tW6zNdJDJ1J0itkRL2/y1adTFK0UoejgfEjby5lA+EFHUrxWVD0u7qXTCB4r737ZkFPdMSaWumzT
F2hdAjc4HVnWS3wE6jrzhdWunexEq1riPbTO9yAbVs2Zz7rsaQy4COtuPVi5o9dkHknDzF13uqSZ
XW5cm3W5EVTji0SIP+CJiI99JJ+vSRGFuIwViYL21O2/evR6gTOrb0Tl4FD/FkKOSDYidSOp/flm
fHpyKcknPNcAUbcqJ5DFim+IMdU2w0bfcTV/2x2PshS5Kb9qqZEDwtIHw9XVp7huxaS286hED4ja
Z3e65uW90pKcTrRhHVrZk+8dOgKOSb0pi9HukwxgsbG0Ei/Bjwmojn1iKN/+kcQS90oSNuEAxVJ0
iuQqtE+8THZQmM2jYWH1VkXejTHCRz8U0MFkXp2TRNtbfD9a0DQmJxJGc7/MtO5HZra2BbXZc3lo
SJQhJ0HL8625J3cEt5x5OOIWs1mj0NYTayHGDVD2OPwyTY6kBwjNjWT7dxTB4BapefZksNohhGkD
9T1MlIxSYYC74rCGqvLfFo7MMqGWx5pZYq7cO0tSY//uTTYHSMwD9ZV/7Sx51CTQJqRs8O4xiMWi
OjMjVQZx7nQzgFsBsMDHy2YmyzgNg2++rE0+cAPpsS+lwEtxZ7OtuTB5mw/OCFhqUJfKR9FVOkFF
vvWd3sNQ1jzI/QOgCRZTWtJLQcWkAhd3dj/9m+0O3AaY9DEvU1cp83pLSEnzMorDfoDYBf7JMuAW
OAzsI5UwxOVFWmFQb5JD0uX/wtEliumotvmXqo7yEf3xCA/F+rRc8EhsCyZUvxVgWhXcULx+fad5
oDTZjdpu7/brMrXqFRWHIW4defiKlsUebLZDSrQwMSzR7REpRWVRRKEhMMOEz1cz6CSMgsZQW1lQ
yRdZPSrgf3Jgtzr+ZYWCr7RsALYGQ6y7d0P2VCenaEzMWIFSXPO4MkC9CfXoAicJjWJ7EjdKvqWE
dJpoc7A4us5RG0jYIRSSaIB5wkEc/QzYkwog11K8tXGUyGXiMoD2thNXqu4qvUgnJVOYXeTsQ+hB
5LzZojbdfKZm+Eop39hHszakJVYghnncO0LYYDuztBu9YtwnkA5HIyzpRNtiTD4TcS68GodywXM4
geo7/CkIUpa9c8k9eE1gGh1VWKkYqA9t9O4eKk70gR/Sm3sdL//53LflXY+LfGvuFhtqq1+d8Dxc
zxR5bpTqUgqpreciaAAOGjdjh5UP51oml/sJddnQX+DmW7PZ8eXGz1E9bRFjkBceDmN5VtrtgsyX
chaW7XeWa9aBrRAlysBtqAOxeUFyYNhpC9NJOLCSfedzS2HDICQFG73nMW1x60RqEd6wtLWUgWyD
RubrWBTWxAQT0A806W9R/KMQ8WXPH14FtgA0jCH/vhyHGHbIItXg3/2LFGsNCfvlmKy27pK5TUCJ
66XeWyuBD/5HQep7p3p8cETwudOOgegEM+YEa8z/AH4PwEQOydlxCNS6UCAbjTRXgkReNcr66RxX
eJSLq/kHWgIotEtvUV2W2ITsyZWwi/OH4jyEOyAsiyr/LTd9feWPtTHVPnIFkV4tT2H4vHqk0Ftb
a15McJ8EOboh9VmYlTGpvDDyiPMXnH6MGqT4TB8IZQXs66wxerojuO9g3DCpzguEQCSUIJ4AP0ah
VpK3Qws5dAy7PA1/i8BZEtIPWcL6tWrc2CQsT6zGTEh8RYPO2y0n5HYOm6jfhhLqYfMn9dXD9gjK
RzovaamyNRwS87LXcGJTXnwxMmcAnrzmwXRATbx8uHmEJamqEkwIsAtE8Qy/S1zE43ImBFEcq7/Q
XzuACj4/cretgkJFTVy42LJyvsZLLka6FSyHUje0QIrQcEqeDf7d4Jy/VkOEHg4nzlHFjqpZ7jR+
M2NC8YgkKk+dceMQxxaxdeKlruqqyX+r44+PUkznwh3bLDOpnhtgDvJN0iEsIKVYaZ7oy5aPZgQn
Nt9YNaKBwWknstjtczYHzpOZGx58xamWW/aRCR+4D9KBJcEcCuW4fCcfJxlnRAtDCV5gsY/sipkf
ie30vkbxgE6suKlanQoIgS7OcrHmkotwlfi8j9iCA8Ya0uBwaZMlLGCpJfNDefbOcK9k/9uTUdM8
poQuWa05uF4unH7ipMA9pRXa4LOOe4EHMa7XHhx/k+/CL7PbnJceh0dki8WT3Az0g74cwAhc4LEd
0SQEtDIvQA2Gubhrfa0oLEX3i57i6ex3O3+g3iMUlUzeNhhieTf/Yn4I3+Bl2ziFaXq3aol4TRI7
qW4JEMo0qmiQCl0Y1KOsXrHlFedDdcWAIFBPg6CAVYhV8Z4rLgjHrycd7f5VGculTVmzC9/AozV2
pZJEizLGf57fmTzvdUFzBy+SsEOKcRzgwF8bIKZlEtFV+Yqz1IMARfaTDa5wXmzIrMO6oXpXVW+C
f0e5JPrmA577C9AnjvxUlhntC67417IFBw9LRZibqa9OjVgxGImZgXIjFiCzXaFLjaiBaReCEzRn
SE8ZkSPEI8cG1EK9EM90KIYiUXznUYjdhSMrQcHunn6EDYdIguRVxAdIBREG+j3i+/FAnfMNnlLy
4DPzoygWiPuc5mWXkH8XJLNpd5QSb/9FowDDZsgY1hBnpn0kkH7qS4+jy7HoI5oAoV7IR77VE6Lt
0Dg+A4Fc/XCjQpagq91UVxfJZEEPByTE1TwOGLFlMwE6W4yASryPHQshbLpA/7T75mujk1qU0Usv
avTmbJACbNHVmVS1AuDJ1ETZDbsr6cW18nU3sHBDM8pHErWgu7fqijezfcOmKYVjfFfsNYruR/Vs
/qkh17FVUSOCr/Kr3DR0vuPV2DcljAIv6NN/MWudgHgyAsU6rHclUF9Lxv2X7VBNm1Umz1FtYh2a
iYmPw7xPuKNmKSgg7HkLP7IeH9PXmRrKIWO4Q83NolqR/QCIzqZWEj5FwwoKsyXjxhOO/WIFEvYN
wvwjx2nn/kS0WOZRPmk53fTj1G7MBppiH3+SMYPDTQagRDg0IaONkJSdkkfPJyx9llzJamuTprwj
Wblop3qtiSnzOsJgEQyNth7YhvKj5bZerOT8lTbGcv2ikeamLdkYEtV3WM/mwvBKnJCl1UYFxIez
glDQPngXmy6ju0RqaY8rRiLOeolC14hKpVrsJ/57eE7p78GHQ0M2HKtKkx0s3ScV6mnN6+29Tum+
G3yiEfWJYVAGcxYDd1TS6bkpEiK0dBAmdTVvlbtGiEOeqO60zE/cwcq9eABzUmJGbc6I4u5IY0Io
VF5utg2SVV9xfLxTaaCyk9GCpqkGZacniNrsOxzLO90l86d9qh2I+Tq1F06YMYIa6Wmx2oO6nDms
rFhWyAqGSkDOF9kKIpJoOXN2Qm/qogAEo2tkBuoL2zWwkfH/y5MKGZ7ngVJNsZo5byotsuKaL3hk
dXwhnFyAublHqi2L+zH7ZYd9uZ4YBRJUkm9VpXZZLbyTvL5wcc9upR8kAMHxm7ChkHEP0ztNGt71
ldvscYgiLk9V+BX+01jTcXN6ZYPQjaufBZSzRz92f3i4LaqPkzcGS7uGHoiwhWaK+/2KYBno5ID8
oYy2QYiJ2hiPqiscyCZwz45eim5jZYS1WjXxjxk6OGzYayVqDhd7K0bu8QoFGQE3FrsWFpjVst2r
7KBJ9WqJd9aGjinooMlPO7jcKE7JmRM7BGtMQq4/Jie5unI6l6E99VT86QNh19ORBt69/OOdBi9g
F+1o4UL7Dqm9ndjgaWtU9++VgSZWCtNW+VzEZFeC0Ov9tc0PkHNy2DBTk3TfqSAIWwskS1uP/hDR
gSMb4ldWYIWDBiagdWCTrn6Yja8BFMK6YkiQWT1eetv7LiIo9k7XtPJPb6NENVrC0KLOPXsV7F9s
sefz0Kbm2APNkdQ1loBjNfRxYMecurc+E1j3pXcJyaBSaDSlddD1KvuQxFpq8EmGq6S6LQkI/FqM
leOD5Trw0NMpbhuxa0uHwjCfEFIPNGRy7z8w5t33Kos5TFKgtYgbRcA9n55g3sryEDYyDFZSuvyt
trO+HhJD/N6KnCJNoOzKUTGhX1ZS4LjXrDm8+1q8rNXujEVW5mb7Q0Rj+COkzRmb1jvOlbKQTZ8t
4Bq5R/nsgGjOSWepCreKByCh4D78s4q4ZiDf3zOMzjv2Su684dzI8ptwXwifL5WawAg0SBP5a9wj
EiRqwgGVgNxp8pQR0mG7EbwoGhuZpsQqvv/Lo/gnCPIv2XYYvr8ENvJchyN5mmw3SuYzTAnMeGS4
I/6lOrTtF5woGKSZD8iOsuxUjskcBTic8a3yQ48fY4XooIkwrfq+Ydi2lYTKf0qC50bDM2Kryzbi
nIDR+QPD9sj7SaXyLhnVACISOSlhur+gz3PjdOosZZeve6fpOx+Z4G+cS5w5J5xX7mjaBVZvkl5Z
rj2mQFOkj61CyYe8+e88pvm8ENujrNq58L3zNeunQCoX6esaRUSrl6iar4FUbREgwAJo7D9u4OFz
Z6JklrR68v7ru/AHYFLbmp2qNUtAVjjp9VZGPV6QkFxIB6ueEfWZIMzWPGWebTPIWZ6izQP66131
he7A1qk3yuoaLX1U+OerUDNzswGJ7R5npfzwzrREwh6UOExFWf7w347yItsz2O39VarQ/Dj+XtKt
3QEwSwPBo9P4aT9LPxR/rIAiUFXpeQbOVggOvPS3xuoTZSoZnI2GeOUKaedqLEmA71EL5ghOAEXJ
FEEzRwTJAsXom4gB19x3uPfiKjrJg1Pxe3X+jKNJ4fUaspGaDslLpiTs3u5Emy1FKn5xDXKGqMhi
gwT2V5SD/mCUWnTJURA12rS1dN/0BLzI/d5wx1AYBMzBNgA45HCEaQyBzuK/H+eme/+6bqCF3Y+E
NrU+DGh7eam9OLrEjYPfuMZQySO2zITaONqDD5x2Y2/b8sAINAgf7PvUOeH7riQZcjaSRIvbCE4Y
ce0hHQLZxW4dvHFnb3Oi63dt4a83uCKyYAcRntW4o5CL10aorhtJlmk6XFuKmHJtzgymQ07b6kDg
gBn3JlQ3eEg4hOVqZIZxoTg430N7PQHNL2WbOZ9FCmXS4PaNjwlhb1wnSbw0zwAV7I0ZHg3UDOhZ
ehnvaz1xzt5Tscm4GDBKvtvKOmQAzQ2qCDnCiGEgYlDOsuNtSILaPLfQVpwmxdyIV7mjh8/Nc6rc
91rz0botazbYWoIZX6oBTYkGcmiQIPe41WLm9WfPIyyL+KMIvI29OUzDW6GKD1UxS0msPOC+/oNN
DmW5iFWsjVORqN8W0Ai4dCeDQYMtqm+BfUyc9r2GWG9hS3WKxYighxN79Jhf4AQ25M17wu0HXJfh
lTy5NZIljT/gyqdZTzpMaul7uk3NTwCKp7kiTg//goXzyUbbIMIS63W6aNEFlSdEQu6pBfv4NfAd
rxY+PzddmsABYD35vOF0Xi92WSX5ynGlISxMn+qlTOfgXNivfTU+yu2ehWX2bZEIYwtIA/dNvhAu
hAe2GZRO9xpXHhN+nKPkwIeNbtu2HB64b+AL2AhIc3u9R++HTISGof5e6CHTpvyupZciVnYiKw1X
rFQAp4wdzgJhBjbQasYYCc+9xv4lk14q8ozhCT3slUQtCncy5gdhtWQKqZLHeyKvx1AgqF0Lq7NJ
XgDg+tZxNrMbkY+boJM+2a0tOw0DiivGSSbkZ6loVCFnW+P4nru5or79K6RxHBhrdAXSv1u+yxLv
QmMhpWM/PFuajSzuCPwJkYE3+s7p9CAsAF+wTnQTgkMW3Qrbex1QSzXogXh4QmBK5rkk9C8tyFro
V/bhZHFD5D93E5PN/lAqLog8HUi6FHMQLFZzUoelErkAKkZNqgtxY76KbSeadGHXZ7q7hy0YCvVe
7KmIAM2a205E/cDVR5OFGgq+JHpoOuAJbj9ETwdQHCMzIvkZWQ4JkO/1FE07BNXSEaN+GjDYYGZC
9vRmk7Y46ES5N8+iX/V2N1sZ8ilJL0gLD39jI5gkPzFTq2W60XNUTxBTT24hBG2Pqlwg/MV+PLw2
SNjO0+wsaia1/NVSJE3rjksgKbwsT6yEYQlbDTkda+pBAI/wYU4Oq9jCm+yFrXsnAenM0B3t6WbZ
+bedNsuTH3C8mSfXk0xmCKVoiQ4giduvOIykCHPnFitvjQrwlGh65m0suMW1umdr87C7/UdDYiVa
wMCnDCkqt/fO0ryImPVZp9/XlCsRpC2ZrABSJcGwlzrP95ats0YycuwVZtYH7lt7wVKAVwP0m+KL
H3BR4NMSmNX8sUTzyUIEe0mOK54UCgSbvkO/lunIUHAKxE48J0CR8UXmdfAwsFzKlf78FoVKCd5e
n9GotBIqcLS1M2UXU86ZqTaxIqsnbn5gZ9jJjXVkdLU0is/P8OssRd8M0ivyDqs4FF/Pw363XJZO
yXJ4RnYGw8HzyoScdjllZfBZMX03MDIc2wN/zgbwhp3/F7Km2/IQ1LdZfU+P24c9jc/b/CR+PQfg
wlgyYbdV2uUQFIi273ermmTr7NC0YGq44N1IGrZwm9IblM+ulmlSUYSDniHhMbqe7tMc/miXP7Rf
xl37FzVYjCrLcPzkVwpmTaUXziLxRibuYLQcvNuxc2uyVUBLRabElXpGpNQeyArtNZ3QDl+6aVqC
PR1EwvcaJ3AsvY4i6ibMw/DzUHIPS3/x6EUAVRrzzTigiW0PTZ17qF542KEiF/sUBEw0V8kf0jsN
zmEt5IaMWuc6RpkamRBWRVxceCC+PrY6URCOSvgpfAsdDj+a2R0mQcTCMnVA9ONiNZk5jdX9c4UY
Xwe5GpM8IURCqxc7VjsOAN6R+VVo4vg1Hs+ryQGdcNq94QvQSpMbRqsuaN5oeyyArKQelXVzkdpB
1fIERWWtqgWUYgCHu+dsdyYDKD4mBxFddpkzJLmtkjvcAlFsQIg7pANYzPXKK3H6dtGxrqQToeg/
DWjgb7ZsYpxNV83XwUz5ouFaylkGFNnFpTkI/FLIKgKTH4ySmufOnZq2lBD5i9+xl+bJApGnE8ds
jauMIltQYQ+XF5JKJRwAex6jF2Y0x2hWneeTsif6xtHJpiT/G5DDGLKtuZugWrtsPClvVDKr0O4L
Rx1jOlnUFvcpPfX2E8bpargLAuumjQqtLpwcqffRdm3YZNdamhQFu6+gZCKvlPA4cjBJTE7gjBUs
TAbEKngQkQNCZNPVWu2HQqexVmJ2ooosJFlogR4WUop8/ueSdm/MGUrmLFEbnz014dtgcrMZQuvc
eaSShh38NifBlYusYhTR7FATNSSyZ/8zpV9MVe+Yi4slsdXqPlg8TVKuFAMQI14vsF4eiblfYjRe
y75vAbpRVSIog+FQ8tup5L8w3JOxEXMukWAi/sKyx9KLB7xJ1GkHkA/rUawL+QfzRJAR6+C+Sf2h
zmQqN3PZAiwzjxeoEANd4aTErgFldmf5KXYGrUGkGNcsuX23fiBVEzR8BERzFqyWh1XLm4rCYzvc
tiwBoAPChx6wwCPRhJaluFxEDhHA2VbyKiMyimtFdS2AeLZsSo4hL28lHT5eoqQ7beu4mOKRmBjC
J+hn9JgWQUx5JqXEwu8hpDnsQId8DO/Hr+wT1q1uPraE5tMqz9e7bjR2R5Jenp5LpaS+YTqIQuXq
S0AuLfDA4bGh5cuhnmvhtJnUzUzChaeekTDQaMizdByYPGODWsi1m/hkaNP2ttzcuYZnvrWeyVRY
L00Gm/tV8yJimWBu4Hct3c42480I1oqn2C5JlMXVCY4ia/btx0nWuZoAPxfJUt7kMYBMlSbk67mx
58vSfbicFvapPyWnqjje4oQqfM5vLOEUupsgMjzEWuihnb4vPDrQbj9RXQOxG4PFjkB+LXTu0Rpz
8G9SXY+S9J3Qszvms0FT8cV1+hUGPi+h+QXYLnssPBsKif1NJQplehCvJCdJF9z9FzqdBrWQ9+3L
Oz4IlGwAVd+5d4rmmeMmfZbDJtToxSUWm8Kndru3VF4mAiCePdGxTACCw8FH+e//kVXYiiQ+ci9/
Qx/ytmCsMZzE+A34BO6p0fIatKnUCAINP4XjSrBcU0pEpbDi3vvCsB31GIeBvmYjtsAw1s1xsMuc
XGYtxhvbkhyOZ1bOQiJE+ztQzRYtQf+s9rZUTxS34rpN85Eg7S3trBhFH7wJNnZi41+4gMDUAkhs
/BAeamMOGyoW/vjTcE/UJqE4yfqt7jHW7M8wzQYwjsKTrquW3Ox5/8Lf/09FlRJxK4quiA7P1q1C
rVBCFl3jzv4sV05UJvAY+cuw23M6uCoga2d8+W1Lf98TQK84VQ6ZSG0EwqS4a76BNgcJEo14SFsH
MRdFdczsVHXoMPIC3EUyJtKx6aGyCRCTiWS55QvOeCY9GlaUBqWRcQpOyeKEKnO1NfRghr6Kemo7
2jFuqysifS9eFHCtBmLd8yeTw8iZUuhQCinGHjB7TSWVUBROaMqDizPN3nuCSBacVz+i08NZeiQP
Etzxmd1EH4mM1OK6/OEjevNKVnsCX2DMeFLTM6xZlZWC8IcQhHLwd4EhFyyc2SNDh0UZyyuOE4J3
OblzPBCp2wszldZeNBNFd611XLB8lfTKEhjbvmTWm80wXnHp37PePK+u3psoebF7FkehAMGB2JX3
6aHOf/tvBKBV0gY38sbsonSIWN7PCVLQ+lv+3oZpGhJtBWdq1PQG9JdHJpEeAFh6HNEikRMlw1Nj
GhgKyoCUkTGPiwaGa8Da7PNIcKrXD90me5FYlFpfWOD2n/IUTn0VhXWuz944SpSDXUOgs23TakUb
IGit3fCCSloLUlG5Ol7SWTQHHttNFqOoC9ip6DL2+TwsOyooegyVhA/i3voYSznUS1+eNTQc5bKf
lHDjA7SCxFtHVKj50R0dH8WsCgZaxyqfa6wclkLiipMpBAngprnZqOkP2jpKNwA0fNZzD0OIcPb6
YT/xfuMZt7cxVM40l5nX/FPWWhK4WZ+UvKqMpbFcV43AEkpXf6BPQ3YaBFpg3kwXArc6dlEm14q3
9Pn0qenIIzmrCe+zadgKsdC12EWaeVMjZjNdodqW094/bBb/nvo/nfS4gI47npeOnD1/ymEG7r6Q
WNDWTwVSdXHigRZ8pi4Hl/SS+r5XAhLn48yfm5nbkTmt4s2gg3nmApHxoChJ1sMriBIUbdfNLnjf
p83Z6MOPzU64mTLu8QaKM1XPxGoQN4CjlT6bbEQLwQkH3cGvAIgHkckP1fc6jUrYhhCuFiJeZGBz
rH0lXWpU2Yc63HLWWJGoyDcrgKJAZ4Adh+dIoaAxqUl3ASceXKHv+NxoqJKDrKRjMkr7bjGSMFYo
cNTEvjbrkh+vk2ioAChMe6LtO8PATbQQ8i6CHh2ZEh+cmVWCAjnwC3QeFGVRrEPr/Ybsw/Nxp86a
+lZcEK+SEWt9BAxMS+xloVOkjYAzMDYSC15x9jk2Cgr32eKQVQi8RKE2JC8/9RVk34jRLvcPpuRr
dp8+kc3MMqOQ60+kA7gr/GQzzBepjC/WrSXiju7FmsSLJpqZq9zarIT0m13ymEQOHxFpKld6tIcP
pyKHE+MFKX554TVgdcNeZvTjR4WsRR4vPM56kxtEbo//2tuxWXi8MoW21AR1NecUh0scvLcVDqRo
8FSO2570gKYuwqwRA2ooR+Qz99xshuJ6MGSgMcRP0Bq4y0O8Qv23IjW+HA5DinDHQ4gfUrVxERAk
PGrA2P+566iMksgujqjYg1JMdF2YKklm7IfZbzoZ+Seqz+DejpFERW9WfkAtn2Vm1dTsuUjhrj8k
ohYoR6CNeDFDoehHsvV4f5gqk0zbzapatAyDTl+Rf96ffBqPviwEl8C7K0ewKwwVvx5LPwW1hq2O
3zw2X66hJzcVchQT6PVJHdZkfDWclpntxjPnhozeOhAd9TKVEpqSS57EtpK/zSaOJO7mT1EQ2mav
pQcSreGT3QFJ0fi2rzAVhJEtTgvWlqFSnSjPuELHMjYpc8YH2cNXK/cNdtkgjfgN9R37b4fzYnG5
oyb9/lp9H44xYxHzOBHuC8dyd/P11O4bsC6CzHAioXIx0vrnmqQKIUu6OHhT/sFQlkvEqNHT2kW2
EX4d3q1lCYK1KKUNDqVXtTkBD0Nsvg5CBa4WljJO9CpxyLMUVD+awvmXRqVNJCwyDF65A2qhLd+H
z9ZMJFzGgUyABUP+8ajmdIr/XP2S0nfSdtG1OMOQggoxqR4i2T1BzUtg9UgTuOnbKCyoRLccQ0Oy
Wl28YHmvp1fkYw3EfXe4imdWVC0+srqgbbgjshw+BUpJVIuaIOXGEnlS/aJY216vgd7PGzsVchoq
bfPRYVXOV80xQQaG+u8QV+jLg5Sg+t9MyH5WsDlB4+Kgo29r47utHzXkDxTx8U18DjSZ7rKaXfKd
L02r5N+cttUR5nQtxytBeBWTpDBTk0/ov3AKGcedxSCSJWLlaTK8CMUfbhFo0q0AdWZjYL7gYA6i
+TtucvTJ6XjZUTJMb6k5IMoAAWrAjyAud1kPsU7E32gcaKJfQMu/AyUvItLaOjfTDIjhg+LgrvpL
yNhIru466sRX6j26RLFIkhbsriODPmToplcEvh0RG9Ian3ZQK04wesWtj2y/uK5IyZ+9oE7g2ah7
5KYKUoLyPELouqy15hAdhamtyW4SOHKIF8sIBACHRb89aqFlafw8vL+GwumNiOgg+7dlZJ5Cwwvl
K9JBSMd4W96Z2kpeFG/2H2BTx0TwIENVxcY8jwEpEm2UPHspU7alyCpTzWKNIpEY3h2BmPJQRVJR
qfKSSw1JBERQ6iAdPs5uv56XD+6kdbLC/jtW0wLA4D8NsQS8PP9XP4E+Sh1veozAFHaefyxtq/dq
xgaroU/hl0RIEX9tp1HTOHtWRQjBwirY4dQU/CfcZd3wY1LeO0OBN1PWxoznTwxdHr/k8dDj26c3
R8zYmSTxMId69N8EMNjJ5JLVVUa/lhEZcWIOIRBaN2SWZ6huOrKUNrEZQ+4bj5f2NE/YWKWjuwTk
1scSDM1dbC5Rjrr/z5k9kNtggdlqEJpSx3i6Lr2KcceL+x0BpA7BYzqbDtwIw+ugSIXnUHuhL/Yo
bsHrwORDyTIRlFCUfb4RR8Ys4U3Rxbo2rYq9Rvjkc0Fgsct4kDw03aGmEVJOSxXzOKMytL8Pao69
G8GfwDvZeY/7K9LEzCUiHjZA4ZS+eg682HCoN3AMr+yuq11AlJYSPZJLKc38CyruszXsavlj8PXG
dd31QrOXR15xz87pooSktM1JlociD9ROaTsMTnvXFl4KeE+us5FzSAWjaOvAJSB/k/IDnd7I4aaz
KlZJ3M2yOnmN1ZPXDhq7U8DBM//mVLTLnimX7ZMhVEF76TXE2A7GgwOyWk11hQG06lj1PC6TTTP/
X6E49lu1s6Hqot6qXj7XHl4z1pEyu6DLUcx11KWvlqaIJ8dO4lnJkJrUmvYdwtfhBpJVNtJ3HZzw
AtwqAo01ajWGfjUWokxhWcV8cWE/YeX38kiUAhgnObDr0CC4SqPBLgcyfeVKDZWtVeYxTwUwyl0/
uxW2p1d64Lte6gdgAilo5fwPOwAUIsXVjcEaWYmwvgMXlBMvm+mgjckIDq/ylRgg/yRjDViz7kpq
EWZYmc9mE+IFdIbKl+EY596bvjcFK3hLHsDtP6n8AorGNpObJeGjHXUjdfQKWurtwh7hgeqH+GuR
f0IxfTvryVKiu5WXNjLqoS6O3+j2joePqF/tQIBaRvv69CEc5iQ4LpG33UVz/gDXXDlRxHgvgMkO
q53l+M0cm1MR3/D9eWPdN1gUwhxHmNdjKaNdUsKXBYGVDhImSUDXB4mB14xOxl4+6DsnsZpyC5d3
13ASTc6CBnZNJ4omYf7M73tbS7121khBicKc+oPM/rUx6t0+nIHlRbsEeKx+b4QJZufWrUbUDzWu
AW202hfLFJlYujFmEg2r/jxld8rqr3KOTxPdO4J4VbJ8HE0ACTaKHUP2fNRFsmXnoD6uqUkHv3+4
+0pqAn+iBHH8iAtnOa2P5aBY7TyCP0K5kqg2CM9rz3z2YFjwzFdLfft0f2AMSo1sKqLLwhyRbF15
qx/nkIM6RuuJ3ioMC6096Fke5RQJ2a0owfCgpAXlakBBKlKY/ox6J4EZtIXWF9wcE6hWDkZf/5mh
Y7CnXgIUGfkVBK9DJUI05JSOntxV453MLaT2tPztC3qH1yF0atShOIBi+NhNUQHc13tFiywKMuFq
1ebUry5J4x5DRCufRsZ0Q84sFQqcWKVyi995RMqOmEB/FaIvotMnI5jMGOg8HAtQfWD/jDqBLE3p
svBwTqfrPm8Ph/nqeLMFmjUlZfwPibpbq/veK/QvUYy85oqTKjDbtK4p5ussP9C6KtMYuLpe18qn
JbPnhCdNXOI8NDPVo3EVOVaw+a38YchhsgKJVdK4bw9E8x3XTdD/uo92ZN5d6Wjlg09a6vegJ35D
WKGXgikBWAJ0fMg1askJ8GXtMm+5Wrr5P5A9ummDfkb0kFyVkYjBcX5spWEGB7HGABgVVbzG4x8U
ERzEfA9YZWEPVEXWs4RCBizRjGxxtYTgRAhkHsyy46DllZiiP5qG8dCzpfPOZIr6ntnmyEy9Lc+v
YeTIcfaAsUrBlDFLYsdRb0LhLL0lsPwJGhwvlB9pl96A5F4GrNEnXl3rWiYYsVvX7V99pvJ4a8yH
Mlf7mpb4GoD8NcrIboonAnKqVsi9ZfDMQpkoF43fDcynRF4cfp8NDdjQ/byXCUTLOe24u/8LV2be
2y+EXvHH9ndXmmzR7HZaHqbLBapgLcL879/Wu5kYGC866KxAiFF+jFO+F/SNY3ykO9ITfiOtixBh
uBHqcxM+wqAOohm8h6qchN3og0mQ0OTt8buLE9492VcVOg6jhGh3/utHcbEhXRl+EFxfHtHeaUpI
cUM2feOVTf7Tey9KUOF6f1qc0s4ro0wGdyciYK7+abJD2zTYBzbfB6KBj7VegQQuIso3jwWk7qJF
fyoOAggTSow2Fc44yMZ1povopTLLi2eTsOM270CpY/nYgTIRu31EZzKKBwYTeGmux+zkhgeCr+0R
AT5aB/vpGsBPOVn9Yh5QVS7YcC9gm+BTOF7hqBeO+SVjfg+2cxOcHIxdCcSPE/IcT6+g0q3IJyvy
xgrk2RQZDt1ADnIF3s/uj4t7qKhLPqRJgPuSkROI5rVmZ5lUl4/Hh9zBX9dXPvqrJxslz3htdaN+
X4LKNo7CRK27d3FQABH8hugHXyyVfYyHCvp9NRdYxyQZHFGJumjXyNDt/5ZPCkcyNWFYM3IOPK/n
SaR+NbdLdVtuhqBWL4utKxtfyoh+BmPU/WN69pDuLjak/AmFl5jcgxNXA9CEgeJWkbKvJHd+aAI7
996YmNOGb/xB0P2O/vh2BxZVSzzEP0y3wARuC3VRziNoDKcrPa7ihiN0xgff7T+lu8xdMDWY8pu7
CinhsDRpFXP2CARN0x7RvATqa8n6J0+tn6gR3/gg1UubNp0+TAgFgplq7ADb35rWP6JigD0LCKcw
QPGFTp0Xm9T2I5FPUfmxzuzpkkPGf4EZzwgd0ZZhS46KCy3XFK6NN5Jx05OrzvOJJvXM6UMnFTux
a9vVXu/QicbHW5gJERMcPOgYtxrZ933SxNwpSdZwYZVgUnSAikuvuOsvjQjmMtHzpZ57SrSR0Q7+
H8xdhQkcML/pAJmsy2uu/62e6JQCyTyci/tG8jgAVTSPH1hTJq6VyrSgdCabgyiEH7hfE8KBCuAq
C6lpQRnOlszWFRsfahi5ptMA1R7ED5vopIRz5LT0DJgVrKgJockIfjNCx1geNlkJkWWd1CbnuubU
+SSwytjsZrsOM1W8+mfrfT5pBIPssL8SFgwpgQtzfAd8cMmSIXmWsji3FCFBNtXUsizl/aUnWJzb
XaKgvfPn8xZHxk7uzvd6a2wVvzcZXZodW1uWVW2hjsS4MrfcKMRbLpfLwE4hbYyvSqlZDrKAlc38
EQYxQ8YoxEWcjUWhV+0VBqrDdVK8/Q1foKPjTL63jZt3UoQUQTv1QWVz0rgudrx8mhOJSLpKqmph
3Q734tVoFEHg09RXr/FQZFUvDYcm1b57PMLKGf7V2lVaJA4hzvm/LE/1CNoAeL7B+ppA7LBZKSxH
ezQ6quRgDWb3XskNUZl6QhjTEMsGXK/X7f1dW56ortDTXSTOHcUvsO3JQzc/Q6igTUPsHrfSkf1I
IAw282lui2XNZB6kB6PEnb1Mn1GrV6PAvrAbGD90uzhsgR9EqLTAuwhw45OgVc6fgL3pC74RgvQL
MpINnyRSWl4CSwBZ8FtMaH8VVxvIJWd8dxpCBlq3Z5JYthMfPlSVc5rNrCrJAmh6cibjlpSuxHvJ
bUvNAYwRMMKHSjHSqxQT3LUl7tr0OC0e4RUDk8T19b7gpnyWfdzo92ZNvTRnXqJvItQq6oVktcQf
RZnpDfPML/Rd645rb0ltuPCJBpAppGT692z+QwzhPufL2kRqb4IjAt1k7KsADab2GcYQLAhZl1Zr
1QXZP8elrpOhl37AjBfBrQEcdC4m7b868LkUMWcxJhmH8sQyH7EN9mSe/zjDwVTjnk/hyNPRPi3/
a9OTDIg9TmuAGH22GV9Z9d3F9YhBdEGmR6yFhud2Bg32XVnQMKHOJvOlqu0NOVNgp2cOUeuvFkT6
0fbK0h8S8ZtCouDcxCTBmNolND9Mac13TYy9vf4Ks9xfhgGUpWYkIOQyNNh/7WuhZGfSEC13Vf82
wpj3Vldk1Fk4wMeBCJIaokwKO0eqCNB4l1q4P5bU+WGRYr57Em4whVeEWScS5V2mDpxq1PRZgWN9
4FqHUdUihfA/On9Y3D5u6YCdDWkwKMt4m38NlIkx99IJurAHpt1Mk9/Oa2Ld7Z2RkWq4+GmnLkjE
4Somhot//YimIpjXcClEtmLgjuMgOnryMuQ1USUHVcZ8+jA0Sk6Vx/8AcjI9cPteOuvNCTzea4ny
mfbcY6tDXhl314SwWI8aMRc/C4GutnkiRMFwg8KABIsuUWGAWmS8/OTgQnI3Bk8ONp1eQffnClIB
aJaBReiMH6sA3MmTjpUVpGqVaaOXYkAOjwovqODVffBLR1HwxmMDrVFKbPBxbmb7VQChZnwwkLSE
s0g/Yaj3QXNNwcT+4u14raiOSR8qFnE93XOALPwyMU7sQtPhIZ3VIhJBYKX5QLf/pye6fM0Q1qrN
iNZ+4OI0gaoOhgeBpVEDL26tFV3GMEVgazWmqFGXxRhkgb5wwamu068Ek283zsCEM88Dyd/9+ygk
bQRcWlh1btEVU55OBLw8L/bVpDLMrMlkcCz7xdi8waQJSijVrWvIcH3uiJchPOewZix9QToCiOsa
bgBzv2QaZ8cwl8UgnFE5pByaWSLblIy0je1ZI++C9LgRbfxDhGhEvCXOBedYz20bTVJ/KwrxdRra
aLOSdwFEClQjDUz94kvZ7/Yb9V2F8l4PAYOnWabfW/x8m3/cUVREUTNV5ESniAVg5N1edxPavtVB
Yr9H8x0LCZraZCLRz10bz+ISrKS54T152UwcStAjOBHKVzkTiy60PePFzp6eTWEgTnnsFKpve+PR
8aqGt+V5ysr1LsAuGmIHm2LDJljynJuHwMQSQcqjgtO5xWbErbfXFXnABDKZUgQJAjkALqh13XlF
iFjjqMN+lbWJ9wXVw7n7abLU3GzlkXd+kwmqbpJ8EGfqJruQhNcFtvuWJ54ABmoMjlM1hHLrBmii
/InMawBOndxSZ//+5Ri277e8b5mrX5bgJ1KhbZHQMHgIo7SBLzgvEjbyEi3tfh2ZHHSTkz9tKfqY
wa8klwHAEzbM91Q8705PXMUonhwvUy/CIW8t5hfqvVGUfzxvP5kcE2uoIsUR1rZX6XM4bTtzqn9h
WpZWbt4w9c3/wcL0vtUYqGbxtOg8cPDf6Il3XGI26lGMgNgGKU5SY7sn856+/5rh+WRvHb2sW1B/
sUvIt6XzhcxTd4V8/DxybvK/QqQUPE1wDptM4EFiXa0p1x6oGRCeYzcgZvFs0rs09YdNGeRTlK3u
eNmXyFWVLO4ZXqZYwNrWeoDx5Kd491Rp3mZL73lJOR/3IOjnG6HnIcvVuwug2py3ecvstjOMi3Bj
r/UBqZv/+pGkDKie9p3RfVn2h4giwPuK/GbD613ntZYjCsErDEnp/aKgqiBpZtEDubNvoOebF3ol
HMLyeqWyl465WtzTNFC5AxchZmRxUFCBdVn5ER8IpG/DwTbXxst60rZnSlJkcyOC8/IuOUNw3xDX
ab6UIQhOPAg3NcHv77nGIUZk6pRgJylgZYHMsV2JGO5AzpRhf/Vy40SXk34PjAFNY3VqLmAdT6C7
hYMTPrnu8ZBZH4LX3EtEdTjpDPFykqCJTHyyp/EBtDRdyHaU1RLtYqy2bIxD0Q1mo0zvgaBoFLYs
fWF1RRwBG6t3+F0aCsy/EDFHqjSmOFmgcXyuDnVojgKjyiuhapZpOK9SNwlXY0mfrYyE6Q/IQWF/
EMP+9O7NSU1SlNFTGkD4M428DWxHuAT8SEirNedQC778Rt6NWHDKadNjRBtIvH+1z5jO5ycBNADB
RpjUl0CGV1+cy2jnrBtXUgEI2phJSpveaL6LckI4UhdmL241PyHndEZXJrn2lSnC2/o2NaTOXoAa
oehUW7tyb5dpZBr6TRcVCdYSmIsV64kNcaBDUl8hXV+CZjwhE/DPDNVMAHejCFQMSFwZoHh4y3De
QvIOkgLj8vnjHrZaFv+OXEUWQtIW/tW/hPFAb/YF8S+xN/W/ZpQTvQh9kYbyn/TkWsJ0tECXQPxH
rKD6R8R2ARYCG/iK57jBQ0GVY2TSSKI5o7SI+sS3dIlIMio3vMIWDda+uw5GE0xo4Xho5jiVqw6W
bAeT3SzTNgq6/yYCSdpEI10TjEZPzt8Q1G4u2881vyFtqECAvJubbZBc9t8plqmRxLVfAEq709No
dOTV2tY2SuMczspVy4Wv8gYpwTCMNStm74eBg4kEV856jTsHZEU/DkEx+g2mypWx9OWZDzgDV3S6
tPJgi5ZnIZ9Q40jl7YW6RvuVqHhK0TwBQHpNauN5WgtZ6MRjh2xwPB79YKRXrf6wRv7j/ZEO75SP
zj9Pm9o9mPSDXhYmrMpDMlO83dZOHORqYeAXzHpHmAF71JoSpif0zY0oXEzWdBAReJx3k1yzYsWX
G/s8X4MY+a7cj+oQpuksjE+L6eNSWShk6aVkrYu9G6nZ4KVeaSVg6ZYuQZwdPy9Rdq2263E3sAX/
FVLhuZnwXgXIzQRgDzpUbRlvdSdb7oVOQ51vwdnq4jf2ivCoQmy/mGIrlwaKmKOkoG81VlebLacj
iFjpunk8eYH6OeLLixf50awlSE8bQG+i5ixUhU4Rk5yepFOX11x9TmK4ZXLs9NljmYHt5XWftbF1
e+lt8x1wbIlIicUxR/plZVGsqrskSGb2xizF6/Cn5bPjj3knE3ae/AolG3al3imTEPOkzAz5CMiN
MVf9w/TyxT78N4gLUg6et6qbj4qr7hhEs7l2T0xQ9Hr4aAx0JL5vfQ5szKyOWqi3YlbmB87Qswqb
tmUIrSVtbwkqJtpNRRUVaGbzLR/VTrsXXzpy4ZETkS8tlpmf9Ho0XzLCCNntPXC6pVUmWlTG+yAu
FCwgmAd4KIwiLPweFj8LAZWAc+0BlWg3czbS4J+l4wf3vg5Ohz7VDSwPk1bqguDlDe5/9llX4q/k
YZiVJza9+nkolrctG07L1ZLZU+Yu7ItM8DBjZAgMXQ1/q+dVr3qpQy1TRL6l/gNTLK+BTIIn11L9
A3lhgqdYJF+ZJZAeRDzBStV1NJIB+IVbjX0ucb6Yl2EJcbNLrd6p1u70Oj2PuS0qhNm3lJrDMpjB
UjINLjrUMVNeHguVN/RKcNMvmhs6J8bIb19wxqvTNLx8OmEZWxYi/cG9iyaiBZKhmrJ7Tq5vBicm
333LDyqmoLicKYdUnuD+iFHe6m4S9015v8x/nWhTM4ehqAm+YcP3W6oC8JHWadaC97o3F78fHg7U
mWJTv+ysfmnJ5vKV5NrW1ilEq2/aELQ/zQ/0v2wtD3W9QQeUEWbqLeaCeDHSjixeGn6lwU9it9q1
QfCODneue2m3QWHjpewMbxTJgv7KK1UmbmyMEOiJldwTeeucL6XrrJYR8Og5nhDtg/n2rbAQyaGU
yb5Hd84P+5Boy2h/h9jey9sfGC7jKgNjRBg/OTrymdv9PI5Xh45g7T8+nhlcx1vXVkYmWP6uzPOd
o9HgkvnCh+rrvm0wXlJvAwLtpbX3AjrKLkwwKDEb7nNCtLeWCx0/HYnL+zzS0n9You3SOxf330aQ
emmz9Jhpk4vUiMATvw1vZCf5v75GlKGJwffhf6FzOnIP6ZMIGaj8V5HvOMXjGSKVUjO/ZL0siqIr
aDJ3x8lkBVP2q0Xk9JnnLYOVVtbq+ckAmuMdHR1oD2dxEsRkFh4Ia05i2nex9empN8gzdEkHvEcX
6JtsaIuV7B/hdm4Ue0FzuUSyoBKgeNroDFbFhzPPimND5ItV26Ay2UyLFYjeYvlhTm0rFFFefkZO
FF2UqvqX0/0ifgF28rNJpRzOz7DsxRGsyvEGSVIcREpa3RPZpN96FV74Q/2kKcUXetfa9S6qHTh8
VQQx8p1/CqZpfWb3KGOXaHR4AgAl20knVRLudb3/rrT+FYDh4YuF2Ha0eo58Kwa1lRWrXFmughQz
LnX7wc7pBxnmZpYzrk1wyN+jeL7EcaAGTbxXePYl0iLZfAyeFojCqXncazb+BmMYeotZzoWg9aqp
UWz/Ufj6/fVXyo4L4JlG/Qn/fM0crXTGIQk/Ilet2irWX0BlmDIxZRTKk9wNxGAOt1D9DD5v0GMF
vae3Tb0niRTWoEPA52E02Vacll8D+10zrK+QqoWbGXqdliUXOHLXSG8fI6ZRhwaVXpynvmvjK2Lm
xCu7QN5BRqAm2LQrbZqIRMYgsELmT42enRixN/W9/iwDe14VLQ1zJ7sqO5besJKs6PwM4b21WFFC
bNHF8xVDk+6mu8BHUwBg6ZjJMhDu3PZLkvTfSg1kbfiMDm4LydpHk9+yty+a5U0aRbfNoxURTuRO
n931r5oEQ7A0W7Fu/DdSb0ch2LwIiRFBsXLUwVL7VbGKqZdVrWKGaFXxp/uAsKfRI8+TaoAmR78I
yiAO/8mD9Ad6v1dffqsmOhq9AMWo1BTwfptsx3JVKNUUq5nVUwVckH6QSQKDGwCnhIb1vy0Spjkt
8TxvPbLnj9eolQkSNYpy/oO7NnwzsFHo5cvONioznhSBillxRHK+Emln80qll9V1/LEYMl4mWhYC
y7QeeY5fOi2Xwhwom4Dsc1pHMIre9ojyPLydIYx71efFCIEJnxCQZ/w3NbkpT/MU7KBJSM9u2BZD
JDiuCapoxRNBjptJyXsoByxfFknH/B9EYxh18eUH5yU9aBY1NI6CDmgPWZ7iYBhMSBbV9tQJzUAP
Mknqbw1nAWMpAWz8/veSIKWDf0zhJwy418t/CuzL5Ro2HCqjhUPTi869j7jMTK/aWFaRp8w5ijZt
wThlGnYFkc4GlEYGx1JZdX+E9XG9KhaK+yMGtiqFERcjo7PusD2dheADu3c10Xm4y4+s64t1FlCH
3f1ncsWIJAU2UemSGh/42R8W1zaCz/CmlCwHj/YY1OwzMdJkvWzTNAz7OMQN5K4TT4tP+661VT3T
Cfy+QCwKEQfjQT9CdTwtBsE9M5RnQq7yp7E1hR7CMjez1ZaSet5m2raiUGsMVAga7OvJBhEH83tm
wpahNHNUjyynRjCSFvw/mBaWPu2oeLhnCayUksERYnIKd3htht9gvAmLnPFf8xk9ROm4eqxv3mYa
ULa3cW0vbn8oDJzbZ0lmKzKRCGf9P3HKkYWmHz8UfUoPTVVZZOcKfURqQut6cbih7mD91bzISuXH
bvYW8SHsyo7XFnw2HZHx+TDvM50x8yI4MhTeflaZnNh18MkI0IwuojXtgMPLQlpH6C5SxRBMbzlQ
XFTBje8kYLU22bWB5STKGCkhgea4h7NAB7a+0Atg/NHuAUD+RMe7/V6hAfsb/UD1sUpqpIn355VQ
RzscgjgfcyVvnFVBUkxek5oHramB8G0BnAVa8COR/nRAZANw90yLtWOyARKa8S6hHZb06LtDqcZd
AJX6+6UZ2y26qARHLmdsy52ANqskhb0pKp9rL1fh+hTrL0MxdUVuhLqgTcqNWtoH4wdtJfLAG+PE
V+eDCWmnpDxTYxjG17Z/+BrzU7yFRzgEdVoPb14yAxxGE7CfgkZg1czqTtuEvkKrIdgvkI5pSETQ
9bZzycBscgl7gClFvzmny4/SmLoRkQeFXfWXS3uszvKBTPsQP/1hoWlSNtJ4ks0+FiwPvh8ji3QA
9wmKB7RniM+lMoipNkl6PSyUxMr3PA+In2klqV9lRqDd6fMPyowel8aVJ08VtE+7TbIJKsPTTxCG
nzNB90rycgEcmT94QJd2ZdXK2Fpi6LAZtRFojL7r35NJlAe5bPj7C1/rgMliJrXPmQfwM/br8+tP
/ZJHrBzZjhkE/MfvlwCEoT83MDHrQkfH9piBqLmY3XuIVPN3MaI3Wu4LSggm2UOAkVH8VL3nOimL
hWAxw04v6JbPLoWfR9apL0sDqkAca5tCper3G0BipjFVRaYOMnizKUZM2bsC4PMq1oAXS/71N5u4
YfvZCGy83LH0wDm23wgaTpijQPLoRfx6D8Mj5MsFixWQrm6ImXsQkeSLdZrPxzo1x5vcO7VNyt62
TjDrGqK9/xpC8d+yssI2xtqnhGQWe0PADhSPnDzHQ2s4sQVZjWneis7u2ANOtKEzDMr3QuzaaZqQ
siI/E5Nd27zfPEr86uS2W/HYFtxeNQDY53O+3E1S6vD3S81HsIAzx/HCF32cc4CnqEbM9w/oVukc
2CY1KyRoo45W6ZHjHjPrP+rByoEtWAnKizM0wJLModPkz3DwDnRB7ZP5JO9D+RcMJaTohNm2vOK6
IQ2iHjL1wRaYm9pNZzmytSrEg+xqSMAPNm+AR0Ews8iqv6k4hWmm3622U35Cs7+m7EQRZ9uSDIWl
6d+ob1+2MmpttabPmX3owsCaf4byFwrN1AzmosndVCXCWPuOQnPm86YLUzhk4tp0S3iJXwYz26Jp
ehebyvUIKaPUi8VVrhM15N7xy3ZtSkbyZPek8g5hegKaEPd/dAT7QESP8PFqcYDD2kpcH4ArA927
oOB5ugGt2WIaaO6OFNFqyAh6mm3/ChwC597vxbgXVb2F6Kajor97kGsaKRPI4gGXSEo7I57kGTu9
3bfGYjwMDQFaSp2og0Gj1sJCfy6D1xYs8p2socj7DoWtUuyRTsFWCX11USdraFNfExedHkmoGUDB
3Xzf3OCL/1W7a6tWLjFv0ud773svqkflmVYIDeXxsXW3xPUJ/4MvVKXNMbp4pOkkOeJ3z0vOgvVo
q0Sdsl1spK40eZ3roOnS7geVGsc5SS7QX7eX88fL+5gl6MweRklcYgqnifV3s3SGyBIKhphJTxPa
VtE9njxdly0NAQ8Fqb2pr6fuc2rCx1QGtKWd47GtpePP4xfoj2OAziEff418bUJyEIMfM7vqe+ut
hDPwgRbH2jc6EO04O/CGz3qJKUJRwJ2g4ZEZSjbhV1Ef8WDRMNXQmTStDL83wuOJ4kEgbk/cl/u4
MB6Q6kM31prYcFChw0pF6zUWzADsydSIlQGTPHeeI/Y/yYLeLtAPxaO+njFtKoJ2IHXJHuA4Ptuh
FcRoEtIjxYsZOcyRhFFBkX2AqYkqTz+EUxmco5r0BX+qpC8AfxH99B1fXLHHsO34p75qAfm3cv2C
b9608DTdBYs/yCwMSmg58p8pf2h1I3tmMJeuHb+FZNTfqTlilQuybkCh0UvfEAfn2jbEEmMrtICK
qWVxmYZMqXge+sCGUzVBzWvQvCnVyETMzYM+BTyiaj5x5w7wPQaJzGkSYW+ZCwaXC5JgJZjb/vBC
NtX5ae0jFCtWiH5X2FX3nYTJSzMR73P8/VRFVqMmMegO7vkFlW9SMzXRcGS5I4xZcT+3z9oJ3geC
KI6hr9e+bsGkSGiYQ9n8Xha3+PLHswsAM6Oa6++cpgzGxvtg21jUZRLot3ZiowYbeVsFFE9pwBHn
1s9MEkG9jcc6ODSM0h0unQVe7qQYYpuqv/BEQeVWGHyfxAI8YMRgcXlnNWPhUwmFYNRycTD2wnx9
YFHtbACRdPuWd6TyChXywddtOnKkr2lcaZr0OnlJCnSYgxnJJ6g8mgmTxtxcciXBAqNiKIZ3+1xZ
suALEUCR1Vj28BelrJOwm+x7sfq1ECBPlhI3T718TM9/prOCvsBb15ZGxCvrFt+Xza8Q7I36D4RA
E/tuGkbdJRSnlxiY9I+OTNWGDULjLpyHQxmyeWpQlqqyszQbsRDsgxElXHtj7a82Jh9vFLDAdAkM
17B0ToIKpGUCo2EPkV6lwINXO6mmpdsCnX6m403UCY3qCu7Ov06yNMtjz5dDz2bqfg6Hsbq/QH7u
Ow5YWX0JVPio6ZodXtxUgiT8csXgH3fTc7z1CItIDGNnohuGrR1t7GR1kCyJFQ9nJAkACFUJrLor
OoxDA4A2tpW8ZdapuvV9uIi1sUrH2zTJ0PqBZdhz6c9jajDlgOzFv5vxNDmpGakVMkYijHEE/SiO
AY9DdEGSBIt0PujWKPbWsK0r+wPyFcKyHJRbTkG4udtscGm9myUak69602wU/u2C6BJPUVb1vQ6W
hBru/2wMrpZu1863w4Gknc/PHs4r9zaBOuUo3CHE4DWvvGrVA63vp28fNfKQ2EyzrmSspl8jl6D6
URtZhXco346PUmLaUBHr8qSS2x3esW+6IkXZWASfijTf7uk/o0Inea0gK4MTPRfGzvuVF93uvzsF
90HTBI8leXirdQhtfium/5yJHKWz9X7vtDDc72Ou7okpEv8artzxmGQoFn0M+7OhsGqX+UrZf0tg
V5idJ+lzeJvE00mif1TeKZrDCJWs8UAr3vpKOFH8d0OQzcq6FH+FWG4IkS+nLBeq01eN9OvJE7tp
rEPudwYxike0YDjUzVP+wJ7ID/V10OixQWwsICUh/lnwIKcaE2/Z7aGO1sgl7GAqKEnXDF3VwtiE
ZLBi/l0+HV+F2sN38yDXqpxqucEJYRiBxeN6nFhEMhTWYDJJDb50XFXqzpqbrobFFC3UtRGxU3lH
OyXZK+LsPFBgBOAjTvMlyTQGoDJNN0CONAPyXczpEisoSgvaON9QvF9Ie8vfziz9O/9cFn2BlsLM
bl6ZdUFAcOzsa57q1a5fjBXJ5ghqiNUx3mD8vGCoPqHMSCiKq4wr9mjn6Agn6HksWAIM95/iy6O8
OdOgqRlb/0jP03tU8ZlqgqbXTrQg72s2Ze9NwNU1/z8nR2+Z/Pv1Bw/cVoCFbuX22yHNS0T2day6
QbFqzYg2wTmneRGKlqCIPj/DGE2+qKcG4L8hlVftAz2DUQqxbDKhJEa769R6+h/OMEHpjLditvX0
XS9/5DzvG5TKZlWCPTN5YJ1GbtQ6NW1hbtTarwZNT/wCrUtoOo65eJ8p8xjWHmCaiIr4KMG+mfYV
ewYLD30Mj4CTVsJtPgu3vOqTRFdDOTTIjJq7KnvoUCqlwQwnFYk9b1PtHZbF6GaWYJhi4lTmWfjr
x7lI1aAhuzW4XmeiNYIWDna230+mrcrNj+F14XnGybpGVp72m3OzXnXqqI/5mIgbxwgGwV1aD31A
juE0rrNV/ozgmBK5vy55XGtdYEjX5RHzGMSzv+FiQPnghrFAiZDzvIXT4BSheevVLdaeZA3eR+vY
XKB0FjgMzNyRcbcYAIaXeHM9TIxGzJMmzL+2qRN+t9r9synxrhfJz0iIE2uNInHdli7MRQ9FWJMs
M98gbkLeh7Sk1ySvn8jtu6YXRcK6StRIixhPj8dRUwl1E//DjtY86MhMJntV9jeHHeM7vtexwaeX
aD2udkHlwYDnPHGg00V/Qak5AuymDQ17OSwrmG7BIIIIP9Fng+IVeq1tnnIgJt+pFa7xQuu/XaAG
R0is/vm1uOdQ0sSfcX+qagWB0oO9Fs/7p/EN5Am+u9+DXkmLpG4zLiCmS0fhrkJeeLuQASonRBiy
jAS03av6f0NXxjWjsNk5zSlAGMOHFE7wzZOttpYECoVlHPd57uEEeQE37+e2kjtJ9tpSB0igQFq1
MBJz8xfQvkdXV8vFAac3lDKXV32+A/0yV3As0prMLYCDzYtjNmK2bs4s9eXio2Qlnsgjc3j5boiZ
26PlCv2YLy0MyeKynmip0gZVBNZUYc3LfKnMMLI0lbINo3v6q+59Q/wr/qf8TnlYRChgpHxWDXPz
Pdo1pOC9hcH1EYOIP6+nNgHH0ybpIe7a6lEjFELSS1OEYNSKiS7RZAdOUwji3emgra3quWM/utll
uUQn4BciMLrtN9+NSR4zcS/GXB/luAmPSjUYvXTbEbPzUH3eCjnPmKyRe8BrCVhF0kcW/2pK3npj
uldYz7TIohW2y4CuqklMTqF0QPszMzJHiGR7tHcmOTMCsITlDeXqe9xPLoWR/vYkhYPuBoZX54Gy
Ii2iW4fLGa6vNCz+vca6ob0K8hO+ZV/He6e+8TjhqmI7rCrYsiq+gMBbv1AfsxfQOuPsq236nPSx
MCZEXGh336HKso2KmJQ07cbvMwTSyj8YBJDTdRQjGFOd7ZNneJAelOVOHiZAeawQBjMCQvdJKgc/
bMy3ez0u6fxRh2uXGt7VP2NKTG4obOSQYMunmo7705gWkufn6Aeuk5QgFaVlchnLIw+Zpp156Kzj
TMkoKMxF+1qcToG3B2gM9ssITCku9zwUJcnQGUfeAwnqB2jX3Hmw2c70qK31xQn7K9TXkc7cqmiW
5S+PszIFE6DswbfjQIJlLuYeyMnJZP45pONIEBDF/xKhQtQBY6IcgZQrtB3q390Cf0WxMggSFFpK
NzheP+o8RhI8+47MyXpp/24pnFv4Nb1T0KlDEAVN0uWA/XaK1ZlktKG1JXcRdKRuzcj1UArdgX0h
CBqhom6ceG/c1JcdLtOXyiMCE50BkADCrLLwSeLVoahg1j4R6MJy2e/rwXtcH8ny4HLza3bIK8Ug
mGFkQYKeexTitNjp2k9XTC3OqQmqlH4V0Prl91nzKBGD2ijYIgBkU1AbZ0Lhle3T+lwlilUri9Qp
+f66lrw3ujFwR/5hEp3cLM8emNDe2pzrL2tTbNQ+qJ1i/tR01sCfeba/pizCWq9koITpWW4z9i5v
tjrcEosS8IlNDcCnm1PLx7qh5G9SmXBgNhARrvQwx5LmfhR6zyFngNBSr4Ccw01vVHHdVPCB7mfB
F0hT1NVtVNSBJ0U3OEQ+GzgLlxq/s7arKPXlc52P1rui5ppKiQ2Ue6pCaCKQ6Mr6GHjikkjcPkxg
o0Zw/W0KJTPJtUNVWhZB+FAKFIdiKzzDKaCt8PjOu3Xl5/3LREb/biYRS4/YvGFIPzWE4pN4l9pW
t4vr3bASM8oP3xzIoXv8IfENF5X8y5nGNd8lDGfl1+KbihTZWFSiVwbQcm1ml4+xmdvEJzy8SiR4
SbDlx/0ksd0U4V9B72VW7H9Ti3sQuO1yHqrC11CYTx+asr1GiaP3+Ob/iI3CcRO5QgeF120OYCO7
wedkKOB6Gi8HxBRV0cUofFo8OXiVU9YQoUmnmrRVeEQc3EGvT3mPxkVNwMzjUxH+j8rvx85iSs/9
EVWjyIOuTT6ovYVuNPZ1ZzDGaeXMJONVxrbMBPYuMftX3y1lqQP3C8vegZjWs6s8eOAgSwPlBCkE
4Iq5srZD7bGsZVNOWaJjjJevGnHmzubNNrj84rJZTk5NFIxQtlMLsqu1qiHt/0XJjbpcLtEBU86g
xKJWX0RQMhFJOJq9deySRI0aRn6o7DTyOdX/RnuqnKX8oitUfMOVaR8NyzJO1PR6KvakeoLwLuRV
p+XGOitkC0iuf2pVGtfB0OfjX91DxJjq3XPlWVMdVjDrTEJFXNDwt7PWVYXajWbuMj+CNMTyfy/+
C4KtNMNvAvy8MXI+7yX2MeSeUr61ZDORX+HVj+DwJRKUl5VNYC+71SmNkjaCHQJvc+dwScpq98Em
M4M91W03jxeHWTQP9/8HY5F5TitTqXXZNIuRZYAmrb9tHCYQq8nl+xO66xVMpNlNrJaqHmCqbAyy
zcq0FRjlYR671V/nMcniB0g/Sw2yxGlp31UG/57xktyh47UXNPLFwofbSsGazMADI5SmE/E48efL
YDT4be43wdHd7TiESF74Mu/QNRI8jsp3vey1mdGdOiHdq4CfY5pMBaG/p3QzZCvcDe1DenYDFudL
pUneAN7op8oz8wLjmOGR3u+Fyca8M62GewMe1xW0iMJzonI8hAR5uU7XuXQZyKkzJaEi4FG12TY+
mtHb58pdX+Pk8r+31jT+Ie1zrzP7DC5qH/ly07lXh6bN4/8Z8Y2U16pwwmRBkbyCz+RTgqQBsNVG
sXmKyYY1TuFazhmDzcWN/y3vf0Hs9BKvKTw6hf/AQRCaBuAEe204T1QfUAQS3JGJarXThpP2VXi+
fx77Uw/UR1de6eA+HnZ2e4Y0h4EgmB1Jik9yLI2EEjUnuDv7I963/H312ToilxpF1KLICZZl+/my
6l426i3PDdQSScVGnYO20EX5y7rLHT/I6EGxB2c3dbaDklqnPu7eBhJgClYNxWK5v1rBz7VKTn7T
TckavRjUcbFCGxdhXevzaxUwhk1IlkVJVstxVKQN2OP+nLhwJI0Ym7jdAg5DA+an2lPyaRn4e2Lc
3oB8xPL//kdKbcHILq9p0TMFVdSVN/VqONxHuNGqr+kUYz9u4fmtlZTDLAPJlQKsAhqcvjqFV8wS
8m1W6MNhNsTT0bljaPu39zgU9c4aJGuHDWfe1p6XZQ79e8b3ehwn4rrDbSAIYOoOa8pSlwiS1h5o
Ht8LNlUsHZ8eyNSAwCMjI+qzxljFMWoFnZ7N7Sed6KI+B+AN2zpnSh8Ob1smbWXcKmaBsTJRIjjt
kz62ys3JXNrurmACjJScMaqfNbnuST2SkiaSnHdh14edCv5hkCCXeAUtXBEDzxMKHSDQnQTRc703
LFM5CsjSb6Muf2BDP+X0IUskLgPFXF/Xrv3supNwLzgQqIFksdY5ToCgPeKeFyuBpWS/vm0JcJRh
p9vfi4D8YwiVlWvheLl6Dy3gDsBej265JcVoHfQqTC3ZMsuHLQcX5ED4N+eBuD9z7fy9c/6UQ2jP
sbsx1C10AD7xR1lY0Dl1hB3TEz+xVZyBIi29fVKCPt6tyR68Odo+hCIlnC5htuSsCRFZEWk3uoM9
zr/sAyPps34L4HWqfJRHG5SVAXmAwuMMwakfyWAPpfc/frCzLL9u2gxBGnqEPQSNky/TpojJIqzN
+foN8XqOW3HlfxqYUb83EbdvUU+6DznjYwZLAVkWNff4RUixkCbf6YcqgGR55QKPY8pcq+BjM2DR
gQC2YEEiFYQ71+EJTFcCEQLUVKmubtHofC5aGbAJucjdv3rLyiR6CZNBGpJ7UX3FuI3zXeg535a1
aWQzShW2rzmHxUAIcEcnHnG6B7I3pvOfNqvyyhO9OtlhLn6dUXQlLar87x0IiBE6t05BzfYc6ZoS
c+dRDR+o8DjKpqsn8pHGjUfqxx4BMtu8O9uWOEX708ENctJ+4XHoy+ojB2aZhrrHYSy1uJ27vPyW
bhyCRktQdS2iubR1SqY/7n8aqAeWOOpXl9KYz3UByE1kRbqCk0xe7Ncn+770gN4UuVet+hWuywHV
uK97Ew2jiobvg9k4zdXtp80AGCNmZa2byl6nHLtOXTTPZoSYKWDeg7g+f+S+AA68nU5ebXtSG/RN
BZpRugeJK/twcT4ig6KHzArelle4dxn5Bk9i5yrd4xTlevulIk6eG0xC/KgrWaz9dlr3puNwLLgd
MsCuwx2AuV/kZ/D2hibKfeRQY4vSASAvY4tOmL9fqsJwJMQw7jAkznhLLjRyZYUklb5d3DbIJXW/
9Ql5WoPBkhGxcurd4aE0ZNQ+g+CRrV3Jsgr3Yrg3FfOHgbvpfg5RgcqfMcB5Gof3IxTxYGKvqoqD
7XBc2XxCnIDmwoFtyxdSQZtLHcbqs29WGarAxvm7er9J79K70k22g2XMRcc5eIMH/B5IibEvrRGL
gok++xKJru4jAFmdm9QJRsIP8bbhJp2H96CZWuX2N9OP+KJgxdtXbeSMR9RGEjhvoUk1M7vLKUgQ
RadJx+j4YDTKwSdWDDtUzGukTl10mRGUqnQi6gijw3s4u4I4ZHCngc9/KHyQCC1w6Gg1V9Y80qO/
J9sBvxl+kCvLBQ4CP9Gk1/bibsOTgrJeBQj7OcglPBZXbmwwnNPuZ8UXEf3NtefgA6AM+I5hYA2Q
vX6ui/hhUFljt6Hd3Dr6c2r2iFShBFFr6KFhBYFrBiVLdQrOZHqtSy5+9Su1CyQtsvXYPmx7xIGa
7Vw3PAqBmYsRI1xL+H6ukzTNGUYjUBJZSyXtNSj6d3KgbW3BmTwKY7Gmx/jMvl3mFrINFRHEKaYI
E54V+imfT3uN048rlqTuGAXX0zImbTprOtfv0URRKGAk/5aW8H6+6775jDnk9A41Abs+95JzFLsM
32xW8h5wDEcRHkZRXjiEuyafb+vi/1Vc/PegLwrowSrtJfVXRStlQPjBybKxJZDpZKxIzc74ZzUV
joLOuaBgX1Rc3rIXGPU2zgTA4H/hcpTYnv6avwiLNIf4SeupoFmsohVWpBC7AOABNqP+L/3rVktD
BruGVInTFeCMUi9PEOh1CT2nbGL0pNG+AZQtP0vuTQFOJU+X9nmQw/ixY+yM8Zrkmi0FBz1PupKY
D8CP/+hNyJcrVeNp+1EmqyapcKkBSRA+/w90fl2dlZmKi08aQW7L28WmxdzXt70Pfk7cjyxMeVun
CA7D1BVgF7hBqdUrL5x5HVfIc0LgbMeXsaFCefP6Wd1zUpWSrHG8z45aYHfQipP7dM3hdJ2RwI8n
GJjFvogQKNq1QGCpL03yoQm6qoZq12lCBm9ceZdpKpMVIL6TGckk2n55wpytlGrya8VCzeEtms5d
GVeAwOvwo0QrxkElQk3Zi2ZacZkFBNctMMOpYqzXeeAuyb/cXpsl2fKncAdWOowf6knaEcA+Ui1A
1MYGvyaAvvOdDBOjBwtzpJCfL5Hr37YfIlzemZWke1BcD+sc5Lh28Qs0rPdcQCN/dh93HEOZYeZI
QwPNtEm9/3D18y8c5K19JFHxkevVicdXO/f57IvzimNwpawOVz3lDcGil3hZNOn6itMZ2pnho/Kq
HfMQW50iHjSaUET+5EJ3LXT3qCnhm53ljT0vU72ajLz6qVvndEyJ9u1CyAofcoYK7mTvymv9KQXi
RhHqQLqaB6t8CRRw2V/rEy9iFJvajnRVLpLYd2hUseHt0/cVV28cnEHF54S3YM4eMFYwSju5lqwV
mCDgaK2oCkz3HkESlYtaW3n3tsZmjIzxHX89OoGZOVnytuLQ/ce+2hq5HU3rfkd3O73/a1gB8Lez
4dW6CLmIC2S3StgRGAtbmKdvzWvgULNLMzAB1saYPA3AsGR35PJksLiCaB2GpCMhbAUFfySvgpeg
pDtwQ0VHZeWvwYHr6UM8WQ9JjqW/3VznuUzIO+8rgHVxptzsXxBdoZT89n+SnJ3ln7QTggX85aft
aZb80gpSxjXcZW9i1kmg7rPGXBUkROEttNc4I8N/Vh/qxIdtAifiFowoEYdJIlapQzjtv7MBjI7U
7o9rzDnv5aj9BtDUZ7CpJ2mEbs0GhqzoSwkeoamACAE4qTEZ5AxaVdkPx1e05uzLPsFAMrPlg9yw
rBtbKmnn5jbd1ROG+fyfXsPUJ9Qhg4kVqpLIMWMYWXGrrr06a887SJea05/S1/w+ODiVHpghdXUE
vZiCsUEjEIi1bffMThEPSWWbCrRTVudchYzHcuDkTGlbfWXyXY5ofa50yVTUyhv/SZP1Xry5br+b
NfoeEBWZI5nlP1Nlw2IvSxNjii1Md5eVOzuGs7o+i1OnSAwEgg1NUphSc+bTPawWywW81ZlQP8r8
NhKzov+6s98umrl2m1gzVsnCmayU9ew/JZT/UYA1XyN3wlfN9z8k37O/faK0ayyeo1aZFFmIVERg
UjHexMLyKF7ZWx5JVTbiLIjlLMFbhDTFhg919hX2pyIlGwAICq4HKY5BmKHIbz8f9mOXM1hupRmZ
MWjNBT8j1QwAB1QEpthT1qdoDQTmIHkZbFLKL9IkSXXG3h4uwwE6+A1XTysM6DTCQCT3lXxDcY2F
UH8i6iRke4YgBXHq05oIAJu4AEVyyMpvG9oL2qBhbp1aHaWMmiH0UK7rzM8ecLADsNyWABib8geo
ceHOSP3Zq9RqXaCnmFKmp+Id3FVx5HvjAovY0pQfgTeucd/91Pp69s72v6l9TD5+2ltVN9uZMFdP
Qu4FnoAhp2vBuoJAPTvPIXh/MxzYWHt0JMC77rfee5iWZxCA0t/XO4uUmG1GryZtJpgTnoiQku3d
E1CmSkj0RCXs8Ek0Ee9ApdpOSR7RMHfFwVu25MlPbvm8p9cJn8r5sDNk6dXn3r73Kd2qKkAbqBTc
thk9DnTMsrQ9YbmKwTxGp+juTZyBboVYDzp6m8Y5PkKvh32kpsUsqPFCGT4M9ChsxuEAp8yXLP5R
5ijrPY/LFffHP9YEqysmzRvkw8tZkyaWazEfd9TGKniSs2ZFWq3IcbRrR/ggldnFnqQHZvIbEBJN
gx9Jp+9HA4Wk1rpgP5Udeca3B4iibBswlQRkzItWpEE4QXYhB3WTKOYbMKWGGg0MiJ7Ee3jqlJwo
HTd2KGa1Q5fYknC4g9D/kunQIy6Kv2+UBXn3hM30WigUIjw2Ln8N+B0b6l8ah7zz9ebjoR6yLXYg
SiL2EfoMQlkADwKjQRI7n6yGbBpNYsIZHE0+3cRUxYO5eL5TO88aABk4ybO7YOpSmLK5y3ddncFk
TNJFM+a84s2ilA6/p2rxMG+0APorJn/A4P5nGPUTljFkoKFq6LfdQq3kiNn0Ff5QQBB7I+aIHlKY
0kF6b+G6m0Un3jap13t7YN77wbIQzO8Ax/Nm31rf1b95CPQixCbohjf9it7ny+Fj2Uv8UmX9bqT9
229ZxyQcwx2PcLJXq7aFv+93kMSHHPilyhtc8dYwzZ4+w+mxWy+WNDz7pzAgt9rG2fYK6Oc2Egr5
/Ozcf4KLu+K/DrMHuUKxXasYJVCo4vgvGUUPvWjQb9StMHuyLpQgtwOurO6VJJPjoBmkzSR1DmOA
SI05oM2T+owj5uXqp4hsTnM0qs8lkIw3tQoPHun+V+jE8/K8ZbqmUYENQjPFarxl9LVOB+76M3fW
xznzFw16tlTY58fPo66mNyM1z9PW3Uo/Hbofj3FXQ20Bn9OlZRDjbxAjFWfg++pJEjYJilSGOSYk
s907eY+55FMn/QMwk2wtoNVeim33F+ZBKMxvcalxKWqYJwMIki4SRn56omGsGAKnKR9BRH8mHGq9
bgTJSKVlTnMZwbrkvtm6eirGvJ2cuiD4ojUSTukz4rANSKL7hCGPwfklQYhgK88vo6mSNzrIytdg
7rG0xneiwJ1LzGzUh6jZcGVjXtZxhywIRbpdkNNjnnYPhwDtoJNRW2UtjziVIysnvsIY8CpSmnRo
yF6UiPj+GW2crNy2NR8ejeC+MRpyWww8mnQlvj2uBIW+CUYmFsaYdZ06cWLE2xxwgKEK4hMOfmFI
8VYYShAkV2U/4QCWkog/jNVS07W2g2LScLi9OzfDtcyCHCpid1J3RfKsDTl5KT9g6rGJYQjGpFcp
5YS4RysOEEzoNndR6YDH/p+kSVw4mtnHdAP+vi+ORNalJ872yhPNMHGLRu5eeI2eiy+UqpaCdgbr
dd71Yeh4Z1M7zAvpYkzezEorScbTdOVbvpTL09hVzpPe5w0i2RfifEQCZazuMHyPIouQin0gA4MX
3hq7kWmsSozLZcGGEYs8k4LyCRM7B/A56SZeJTjm7fwltnmSKfSORVSfMNQEjd9gKxWZ38XyiYDM
9zt0KLeCrx30xyGpMUnsIqhwmroy2FZPJp8r5wW1uo5ebd3GXEdue/AhUWPAAo+VtRWmqLRTYto8
I4dUXPFkHcjWfwBGi/4wJ5OI6kVvWYGbLTI82NJOAihzyA2zRHUz/JwqoLIntWfxsISomJ2ixUCy
bYujUo3aduTMW50fToEozpyZsJ3b1bGtTIIyW6SvPjZvWFoPCLD9C1KLV5S+hyOSW/NVBU6eTXm2
F60G1eRPbrB56BUYfAn5+TR0X9Fdj+5TrfTCkhnVz7zHvL9ooNXBvzGgZSi6i85l19FqffN156sF
3QsDuFCPE/NDZqVRXS+zKN58bqRaeBtzKa6zBAGKJ+IGy8w7AegVHBCw41lI9Cy52xeR8Qgr1VHe
PB4E0ZwtKqBheAn3zk3mo2YebWlfkamwXnScNRYoYxr2ziDw47mWhhyw4j2plrFeYFMt3ifc3+bP
gxEwEXNwYaSEBqF7AWj/nxkOrviLHniycx4toJqvwcjD6B813USs1k22JQwjA6/opd4oAnANY6aI
2EF2Mig3ukJT52JvQuhjgTdIyvRW9ZzHmPsOZaREfnuzcormpjOJ24MCxZURV/MYD1N/JkOkZGrJ
aG1FSRipsGuCo4DSvVey4+XAYKDw7zbqkzkmShnvj7rFS7e1GKHeSh3aAQWsIeuVKZ2pWWz2WVfx
reU71Zv5VA5iS0rdsNtKw5FeOwvw7vfgjHnYK1E27UGmID0l3MrGOVTUorGa6B8KvgEyPlwxW/ZB
U4QzhEyN9Nj5T0vmjnn2n5nM3SnDp6lAUFnplZkbP74U5a77Pg7sKCgVPfxojuumEMamy3ASksXH
x5Z7ccAEjM7bV0GYhaBUhYPj6G9biM4PqaXdatomnJ45UBAHwmTlU71DJ+MNb14JeDMiFBSkiMAq
5VGqHouoR5Wp3bOwM7zmzHs1EMYQpPYtAaEEAuwC2I/bCc+oeOX0c+D2zUBEVyWKIPAUyS56OiHb
OuA3f+/yQNqYjW9MbKTf1uUJLfgAEfVUaQFkJXnuMsiUbP1oQCTbmCSoz7WqPDdZ9ejZm37EvBw2
7uO2210qi8YbruTebyCTuy9nZdp/JgH19IEekJvEBeA9t6pxzb7ZWDnXiPQsXdc1LD102fTPDc9X
kSsGmE4Kp0COm+aeiOBwZSr6YdJ22MoqdK7NOI+a3unIVniR6A9MIxmkTSsUYSctbBIHeInFHTnj
t0NK+0uePBzbMWxvCCS0xTgKRq5WDn1kjfwkvQ7H30eTsk34ahoKCtHpB4fDS2gBvAJgCMAZ24Uc
TceZUgotIcnj3dfwUOV0nU2Lxkh0pcqTMu3IrIS5zcAjyeAfSVc1wxbuoqJx7amNaIuYzYpcVSSB
8WHb3DtaVo045MwlRVSjURTgqC1B08WHtNB6twPXJSnf9Hp1ZhicPi9hijHynOyVgDE7/rV9/Sr3
z6CC4URicrdbRk75hQphXaBb7HRlDwQD02vUxWXL/Q7fbXc04DkgLkV2ZXzMi9isL+OQCS+ls55N
fQ8ang57/vGDch1mFJS1dOmS+3zoKHGkEl6HcQqEhaweOxVMvU4BWbppppZp45iZeM5FjhLKeQzw
HvF9s1s75KdWIXbKMIrhgF3o7urE9JCtRVz9AyWF1au6gQ7v7qDnBhyB5SSpxwg8jgagPfV3HAoQ
tyGData3wVp+5n2FhZvzOSE7M/PO/TXAorHrf3nCSuFIUgKpiSwbcTKROsdB37m2EzavXX28jVhh
m/NrBZooLE1dHwT5qT5FiWQp3w+xXfomn0m3nZ82pSYk8DNoLdlPJUlNLTGyKwIQE9jbmy9dqHBW
eQfumtn+Da7QW/gjtcURyaLM3oCU92F2aQcwXzH9ej14FSqEDjIp61HQcXuJYC4QcqoRO/+76Gsu
MGlKAFxTcOUfJ02ll6CZ7i6odv+KO9Hhtv4Zw+cJLP85estaqCabSW0avwJ/y4M1ZiwOFzcSklRT
XXUNvrpE2yS+yYTUmVgpetunYYHFaCxKIR1cmisCcpavVD0DLNG5CriFrFnFwGUhw+A/0x4u4vDo
cHVQntxzsr4kUVGfRM6Hto90g898JD1Vyym4fRjhTGUj50sAet+uELq+JmzMQD77n0QoCPPF8yeS
/hxxMl5Y8QSDC2tGdh8VUQ/SaBZL21bHdZv25ACsUcVq77ObAiQqm9i6jFMTKHK4pgro5l+PI3eb
e1L5rsvdNR9CgqSXAPvs6G7ZwkS4YUvJFFHf3PpFOV2y99Rh88bG07PRFMJiGnxv+gw5pjGAeHzA
C3P+W9dL230K9zBUungvmtOiEviZKvjoQH02wKx6ugKMJWsYL1vWpr1b0aQbEJsJyon8kQ2Yhgtu
VpUso3zjPfUKdyDOkjtfnOsLNGaA0rCqrBxc8P7A9fHb7qtpJ6z1gtSnkkuJ2eeLe+4IoXOjwI6K
7ogU54tYUjwPOJLwlKCdbQ73+r6PX0jIDndIPKsXwo16d8Qptt8R/3LvZShrP6q7WV9T9Hg582ZD
D005pbaH0qqDLwVNu7jaApSNnGWopI1cA+CKl3k2A+JjPmjR5YKDk3FM6R+TYjulQ5u9uPJ/VDvb
oDwkwF6oGlTVxRZftKoOvoDIqSchuydad4dWRnFPw9m/mo/bCRw9q9XtjNtAzqxiPnzkW4ZyINuh
/f1/8A0fvSEasMTuF1s+PfaECzE1wa6Zjq6T7owtTEYRZHGyIod+mtwdXBOGmsyjVZPt1Nsydi25
S+5XC170sq3hN8zHJxq3D9nk+Cnv3lp6drlCrNaS55k4TxbApFVS0GyrkPcqneqkTlW+u4wx1+UR
iT8yFG8DaNZ/Y7PBugEoo6db2yclmU0YN7tO0zzBCxSnfCQaH85GsTnHyyLskwviwW6C38sYmFz0
VgukZJO5EZzqJpfkPtvEydjCS6PjyHA2Gk6lP8rDX4BCZzmNQcxdsbOJ8s+VihSghc4uzDhGIjDI
Y0WXCfNPaysz7VEILWSsNZLt9TiWu9lwiGEGo7u5YX4/rBYNYCFJNj2ac7TReAygris9OizsD0Dw
N9zbguyigXj9OUS7pUdIR48MPKp+b5r53j2dmOcCdlJkAryW394uOfKkBRlcRfoVgeDVAJPPOMGg
zuFmBbSyEcmmDOv2YWqAxD/rRByC+JpR/7oLZ7bjbFl/dP++W6u/6tSKgPg1YT4pgdAddC5BJgzk
8cB2wPwCgB8H1solrSjy7lfuhrkHwW7bm5Rh2I4EwUzZ6g1WqHKCPApgkjJQiu6CHTDKuL03ktY2
OEiSqnrTOBYrd6whmIspYqZjCO8eAf9r3csJJbtfuqcjdCL54gcqFVxNN4AC8QO9R5cE+2mDNMuD
UrXaZ+ELHFq7LMr7JMS+oVDwEVIob4voNSeT84uBCamoJmRdVkoza/5tyUEue0hdNTbhmsiaOR0n
2Xl+UMPj3YSdzm7ixlkiGE6ybRWpi6JxvNny+bgqcBFr/yGXFZ7EEjTjbIatnBLA/qDQYRInZSdb
5qQJcQLKH3eTasEoDAgddx0ItROFWsnfrHJecqq5SymXVQCAmhHQbeVdvhNXgPxMF5wzMFg4c+f1
Wxte74PW8GsLJnZIZSoA28jnSTrbnvKQUmK0yb1OthKamApByLMno0sPlBJgDm48tgT+vMWIwojH
2PkgRo+bHANpv3ZmGbPmhXpICklDxSo987xQ5wlyxXxQeCRLLF3QQixZSAGmgwbsLjfEjuUBpPYs
s4QtWRd5baiequtAZXxbATdADZYJN4EME1jGNJHBjE5Qq0qDngqoLcQwSz6RlS67ZHuaRE+1dP5B
MWDfRX9Jf4h9ooKvzdyicLrluXZIW7XYH3M4CMlgoPaG9YQScgO/6ctPmn3aawQGvI5NnFRD8WCN
F2dHOnbGCmPq6APR0G/X4IcT0hnBAyQHFLklpZkaSfkafdu5dax08xkcxjVkvVFLKcLGAfYpRcXU
983oZRjhqz/2VFcarnS/r812oCg/54/c53HRSWwGyY8A7Jkkyt5iX30s75Rn0O6FnaMnVDfxfhr9
+DocsRpeJAXyVdIYq9x7VXCEgHsJ93Xg6gP8eoFQ0DcitgtJ2ygB3xi9Vtp1gWkZhU93n/68/GRu
inKNWgl8X+gNh8uHc7Jpjvrb4t4l6VLvzGIFePLjuxg1BOgabLVqIK3DRpekhung1phSDgraUUiL
QsS2cHZt245NbXDTZuqEk5qSzBvaC4/TIsMKHl7lZqY5UpWSpbdGDEa/d1Vf1Y9ojJMBMan5Lfmr
Uj5yasgdH10hjoOC1HaAtr+C1AUN6morFktCnN1dGbqZC65WWW5JJQ6pUz1jaO/cVwibI9QfHAHK
NvHjhlorVr8kv6zLZ48YvEzpuWunpce1fAZzSY2iXcLh19iBwxQybhhcALQypEF1GVLBRp1/LWXi
NU6842Wx0mFXWxiHUC+f78G6Ou4dhBSIF9ifapY56lVbQUjNu3TSpJiuj0zpVbiygRNydaNfb8iN
7HMZ1FqYZ7377B4VjpvhfzsO2YBvvrcgHto9MP1yZaEaqRj4QM2Jfo6fN9UGoK8KjG1vv/4Rbbq4
iJicjkR0C0g0hbrBvYLcM0thQyiImWMv96CaL1g5fSOi/2VObaf/eRJJsDBhhgh0SMKtlJUDfE2O
OPy29Wq+UH8eFm2h+pFQUdaZOa/4hIZzDygHIOuLIJQPsif+KvhxOKetpROJAZiqYzbiwT2UJBfK
PoDURCCc8P+EvIX8cMG7AAp0sL0CtRo8oWQg5vsJ2aJ0jREsESuu/mjQ1Uom5TCDAfwWnWP+E3C8
LdUNmto27EO3X9bYo66qKcMABeAjT0CoiY+ICvmtv5qRy/9k/KWnCLFR8xwNaMmZujVPzIbsjjce
t6FiSBr/ywG9uVTMUivOM7pcQRTQgtMFxqEQLQsLyzZAjLof1AYNNmei9ny5ikx9jfu5tNo3dGXy
PTcIDsAt51LVAvzDWtTmGIUXn3NUSIX/fH1GhGQSgn0SfOHSdRFGijRYggoDX+OZhgLIUPMPY7/+
EQxuINYrk8WKT/jTZPtlCn02g7GIQZW8zMK99u/3Mipb3wwQ5M9NTTbdAOnf/bkFoQVgPIw2Hbof
fcBHZeso6pnnjIr0c3QGspid4/SJORbus7vbqqNqjV+CQ29uoteVmn9bJZigl46AGOdTalGDV5yr
6NMb+JQiPpV1Cc35zZ7CmN/PMDkk+UOSIja/MQhrQx1FDgMju1/gembA46629mcMi1yw5jQNbNwq
MCY7tWnfrQJI+gRZ1PUlnKDj/NgWZ5bK4J0VrNJOv/a/p7Jy85IsKQPLcseubKeADCbY+6TsDd8v
kgfd7jPkWNIRjpUEmLblW//Qq7uyr4+Ju2qm094M6t+CSmU5P4/vTS6wZ4w3PxwzdtFDqeJpAnQM
cjAw67s4Yhfzr32FH9wIDswkf8Wx9GFVTVrF4FVVCX/TkCFRto0ejISXO3/EwEJD7E1lOq61B4bt
xaLO5U7R13Dm9ltzzmhD5xfa5pSUf81KpllOAAlP6/+VRwn4hadhdrWTwpZC5PXlQKrC47G2oeKO
zPByiSw2d4zOWHqA8nu3bPHNm5ZB6ejJHgkFOEEHD/Nt2Wc89sVfZgmjuvuj6RGGk392iEvezo/z
vO3m4qo+hp/kJ23u+sKDIvu6EwgknDDzrWD3sTA30pv3P0a3UWpRL8PRAo0LzBmVH+XMN/PzQYVZ
5pxRyKaPaTLKufARCgDHOWItl3D+0b6t6i+izZ7icU1MPDKtQxwQ7IczMGNtGvCSV7u09lqEXCJ6
odfpfNDI/kbNVn0KhYQe+MuLQnRLXKK6q7kg8fQKGDX+4i3p50J39uO+HZK4FMJ8YcdmMreV2K1i
BfXWCALq9TWHEvySfX1vANHf3wTxHBcld9guHBClQXGzEooNL5WKjUGIiQih+4zXH7UHZRyIZc84
ZXLLrjKZYl4CmwNeVUxNMYD0ZBS5idAfAFjiTiiov+OQIQSeuIP4zOFCfWH0uHQ7eU1/pqthi119
FM8LGd1NJG8GbLgr/ykiaZPOm+lJNckbpQGMTPIl/mLr/Caw7fl28gW8uc9s0aG2KDbyd2/rNnkl
TLhzM2cCcTMn+dgeJz6+dQ2av+mtKJjDqjIs7vMatsPRsZN178acD5jiNuqsUr4YJgTwKsc7ay6n
XciKnxvxt7FgpY6xJJ066u/I498cDw01WMK1kr2A03D+Or5N+o11XInk0VT2kpLr6/4tVFW9qvYg
fI0yvBeIeYif3g06nEucOdRMDd84ChyorilyzEY66ElH5J2b21JKGqQgKF5aPslchwAMJR5+Hd8C
mTJ1EAiRraw6WU0KD/BdlbRsX4Zrkonn3C7uXNieD8yHLjat1MDnQhlBRgrVqBw8U6/EfAYleqIR
W8Vmqo19xEqnu1HYmHtKslsX3/h8w4DEWmW9cVAKGeV0ACzcUcWDH4BcGRz+N61LbenyacScGcaL
xdtSYLcsMZTUy1Sss8GSIWw3nFfygVM5Mz4Az7l6yJ05veZdM8DuKDwuf7l5yVIXXMeRcrNMzLHV
r24NG00gtLa1yLCO/yu1syNGs+yy93Up1iQapEIZUJREMKZJoTRHHStSmeE90fVShG2ZKFX7gLP/
5BmRdZ66XAYA5X/mWRJU9N+oCja4su1N4ErzdDi3Oi0oeLI2o0pZyi+ZFoCYQWwhxAC7Cd9uhZAS
seNModhxwJdQgEun21S+mD3PYCsYawU7DAp9Ts/HjCXD/74lEhDcO++aWTlkiMoaOn+EOuiDVkCe
bddkPW37VP0bC3LlMxXZ+1lY1xqzr97CbwSTc93XvXvIsuwGo5agaug5gjiANwewAWXOnZayLLkh
Fro755tsuqAVaP2HkZkHPqVVkV1nD5Iecap+OGu6x9L5PcQvWa02ZrkpBLTb2GbSA8Q9X1yj1/kL
Nw/lvN36Mqztbj5q3NhRKz74QZDv5l643EEx9hcJth/dZaCoNn6NzdGRATv1aL5XXJguNQejosTg
WEvNooJS728UkYdJbv/w+B/J63fvGMA4W67APjfIiOzn2/jKEdDD64hzNO/G0Dv50a3VktclXz3l
IMC/2TR7vHU6Ix4MzlKqnzdd7jcjqDS8VnHSrNlSdc7PS0nq90ZGgLldfksCb0dYIt+PxOeFoETw
7nZqfCPOGEPicBLMvsRaVpnZuYGsrfpzA6HyZXdygLMy9T63vJ9ViyRs7hc2HARisn/u7XYUVsO1
LW0PrV4turKDU4U2NtrSqYcFvI0LQQNb8Bx8bAS/PofLog/yI5mU0drj8gwlpSaFPseGAKdWIZYK
ShyAe5564yYeLZ+aQIvjgjJ3dFlQofi6e3gNQfuVoggoD++8bur4k+6fNEV1cotoQXXQwEtWlaGv
DYi6r6esdcQwC0i6NsRzOvOdDH1oAVFBO8EM0AJveF9eKhIgG1Wk+55LwSNga5ZnrUOPcUpTNDEp
bUkGIMk4cnrZuqnOodyHNAkoRMmEhs2S0vKFQaTtNQiuKYFtTW2yQ1MJaGprhPYIjYD0z4tpB1z1
JyZlpdb8sEHrF/JZ5P3m1GHGyEzih5yQJMiPCwnPCMl22R1hB59j3MFGd8OtUQ59VTOaX329wucn
D7rFFKTf9kde0RdrBk5oc6ILvKqRgWOHoaqo6W533CwdzKc22cpKPEYrQ0vBReAKsD2i1GSpP6NF
46A7Uxe2gXkzwkgub6saE0Fd8P4Bd9WOnMU6qudxfW2flobjE0S7CgSKx8ef3vpwNewlAJACEieS
ErKffc1TjUfWa1YpB6KGBl2O2av6BaWfERSVxJal5ZOea41doQWgpWT+N8AKUBpL7vozTeB6hRiY
5kqnY2lWkrNeTPlh5yF2kBrNqV+/oanuSbaUBbQpV1VN1crnK9XnnL61IGETKU4IpxmigwYZaT36
RW1NpL5bl3+iMDxbE1qbd8WqZOq80pRQHXFrqU8TaYX6+d+m51PLlD/OwCDmXHXFITJle8OeNfBU
QnibKoXwjA6NDKttgiBEn1KkGZO4MvKDuNEY/7JqRoJAaZdcSBsoTWQs0ZLmM2zCknErt7naj9CC
crWnJwI2iJDRoR/ieVnZZD9uojcRU6YgSdKy+Oeb71fd0hQycHxZ05KDIid8+Ynd31aDsJSibsAB
ebi/cXgQCRvSYFrxjS1ckDs5aDMJVlfTsd0jrc+i5NTW2YVGsjOSwFt9DGRvJ9qSHA7iSuX8d45h
TY28z5aUGNFnunq5+VcO9ilRV63on6Mq73YzT9ZZ4Ewp6NbnAZ8ANH1wVCX6au74vxdCV7gTsho6
YuxS+4byHtp9lDVdUooY6leczB6JB8TUoh5ePtUZSJDsrRzM9TpwG5aLWVoQk4wzHslrsU6J4WXL
NOo1Sc1lncnTIB1FHvBAXkBtdD9wmIXZdWTGQoeSSuBL7FD2NIKFLllzozaXXQUT3P1sxK1hH2aB
1Cyc9QepzJr5+GzxwuZQYbGBtIxFm1UPlLa6dgHHZBv6Vp/vdXQuGlb6SpT3d+3E+unsHttxNobU
qnaXyimdS2y2ySBY2QNN8gQp9YcH6X+1Sn/dtDXbJDAFL++37iGjhXdX92Nr4OLDdTORIRQsw4Fm
jAIurEeHvo8KOBxyNQnenpsItWHB+7EOrpnACMN0GMmp9qC5uV0U9y9Hl0EXCG5+W6NGd8W8LVvD
MddvPnPBaS+5oAPprYYLfFo8eICLDyBiqZp2Wpk4ea4ppQNTIp0FUX1J8d0s8ew/G/bcZRFldY+F
kMqCuDRktqPv5Wsjmp6Mq6SpHc20rTPt3oZ7BIqidAZ5d+SSH2BXD9KifO7NcwZW+I7dvuQawK9i
Z8wSNy2W2334va3gGL5c72rcYlaBUW3kOnTVCvdGH293zSVbbZdbv9mERMtkvvwEvLHaZ/hp9Tpe
vW5mkc0I1SQF+L7tEt3n3EL0BQ+Gvwr4jjyWnlhsYdl5y6hPnxeBUyD3eVYHsgmzQEqY3APzVpD7
VTGzPVbYsrtzVaXfLTtwkb/mFEzTihYUyq6VNojU5ycdePwc3z6YfETgrML3/htuDvDR+6i7bgdR
dk20PrtynRL1IEUkjevDeZ0DxTcs6bWgL1ZAwL9gw1oqwauGQFpTOybflITfnT1LZjlJ3XBeqZIk
Uo+7PflW2pGNnNAbN5hbKrGJhT9rsbfqvd9vxqYe2zUbSl7XrFzHhm81d555CGPaqC0+imC8On7z
GPkwo1FBcBxiZP9TuDcchpR8AZ/IfoD/PiQ6JrIo2dgSv5Vm4mlTu5H2TLqtLSn8a8Xf2eN1xRKi
oNt99/IwAzyezR3kXTKKZ7pJzYP6RAyvA9GRJn0meVJwpXwgXGcXllWd4sh/y0OlbjjKz/U2QYQZ
Pxp7Zey6afsHvmDce9qT4a259pkKJmFwqGbi36pN6umUQbhWxa4JMtxZbG2+KhuqU85AmDFEK6cj
G0W2oSkzuFhPSJU70XT8zCrbPCdlLAhRhICZTG2tx/ERHQFSb1pDSNTdqiy82XosFtO5DGaeHBDs
aBmsKoOhHIq1eJ+w8AJ7uDCLn+dr7A7jmfRYtpy10GCfV6mHxnMH1x9WZPNb44UO3Hw0NGob/aKM
H5mwa17eS4KoEjwshGgBKUPKoeJFqIoVi60dfUPerp4AHpp6+6OTphfd3+W44ZMgFez9TXZLJ+yK
9zziKvI+2ySQJl7weZahi6Oi3p2VtbLInAR86ShPjWZrkeUqX5nSE4afPaIMYh4mbvuu0e+nm/ZP
i0fwtxCItlpkHxJC8Wdllp8MVfYHkAqnVaRsWpEcqInrUIfIqtflsosWHcpVBorFkZK1IT1Me8FH
t44Jf77+CYvxlgyrG4t+fqqzsDp9sW7PnFAcT+Feiqkk+Zm3toj8v77JflfU6D6HOXGxANfavCeA
TrGoAa1g0pwykJhEk6jlv1e7D0ih9cs0doLc72F3nUBnbbB9ZYse6NJbFiZWOk8jvR3S+FHNBUXR
lfGYaaKmsiqM/M2o7QsFYGaLtsloYzCGY9fIpsb8PraMSy2AgP8ccfec5zePegDlM1P7wilOpdcf
N2LDIz/ZQs6MMOOEh+hwviHgoTpd7ZMy4mWKn312be40VBiXQjC+ZCs/EHhE36ep4aXh2V41lpsN
BmUiigI8hxl3OtX4Y8DTovjy7zb7N3L7iRxWgjiWBRYFH1cY7JiIJGjkscfTlIqOwqHYye+o3KLx
EV4mFEZHkUQF2MziJQgbBNP2FwzcWhMK+6Gc7Znkbn5Rb7sQv303WRRcizCErCA0NsKJyrPJ7WIu
ANYaQpCc/mePtw1LPMzFap1uwHTHQm2mjy3x0WWg+EsrMm6kZB+v+/Tr3lFhaYEZQLlZOU05Z6iD
cfxFLQi28SfdkKOGpBrcpxY1VuBIRBTntREvHRmwDhCHOeoNEKQkOokNdmU9TEcqX8YWkeG9m06P
MpJplUl3RNR3jWsCIcLebPf2zPTiXiMA1EWhMql/HX8oXrsDx5aMhgX6uBfGUwI4WeQbt59lxU5S
K83AJNQ2dUIBPXt5e/eSBBYLjDpNHLfOsxgSNXfi+4Aj8465uWGJRNQSy6sayvEsHlF2dpmbAT/W
R3dn4PdPZpRDkwYHjAlT52shCDhdQcnvJ/rP64NyHPq7Pru+6D73dvB19/no6iCwWsR43CayWsuV
9yqXXDRivwdOHQwZAPi/GW+Jn2hWC5nIBKPrut3DTvGvbXFcg1dKi0xvHxnMRZg9iKJvWPWhuZkw
14d9bX7kyWwbhpA46Q0eIj14m1l49VImDos4JMgls44SJyFBJp/s2jSAhtVG+VfO4MiaClYMCM8W
ZExE76T5O3krWjxYwFNqCPul7uTnh3G2EqWephmshlcvA3DEsleSzDnVfFDbzHbpsCj7bc+Du6Fo
84UI/fr0NVIBwGvxlmrNObsZNQb7IIYIdqLsQAJGPPlr+FH9uv7kSYdTWOjOp9r9/i2NZDNGuars
yH4dVtHEE90DdPUNGdoQ8rECQ4GDkqhYs8zDSrYtviMqlOTF6CoHD+G1A5c5TmLohvAO5OXWfYtc
HCqO/R6at8oHf2EaOeApasqb4uG7K6uORQq3Lt7TLAc19MLTiNzrkL4s5emBUMNYadcewBJnlYCZ
HZQzBaUrX7EQ2XxliAVn79SMoOLgxfRc2EpNYOJjbupBsK5dCR2xQ8I65zYWzVzJP0j+jGpRVrBM
+QYsHgbIEUAQpvFzuWDW6ocKLqLA7nWFNq08kSrDTEaxXlYlBJHxfO1JDUap0dCnO85DHdbS4X5H
NTRCO/5Ye83zQzQMpWdV91mAFsnQ8FStFCcZk99ojq5MjulwT1Wi9UGcPVYaUMjjoI9XKmSXdQY4
DTr7Fw8i6+eH4CP17jQ1WDu5gWu6ISHIOcq/pyOZoBA0L3m9QB2Dt9e3rTVe21tQ4vYDiDVCMMOX
RMDDMobNGo+lPc8wXK3VfYFYf17bqVC3WEQbhNs29uDVJ7TiaHIKwrE5xm7+sTLoE8cHt9q66kUu
dp8a4+iSs0qGbBkwEGq1t9TcWgmdraL/0qGAL59lBonEg5ktBNuEM2atPTN7PxCNPq5pnlDZ1jmy
G3jXjZviJqAGsGZ2HsUgab1qAbWObfq1h6yJR7Gx6QHY+QfNTqV6WfCv9vzDNrfaIOGFmpw7uciy
dBD/3I3uCyumJyCZLbEDkosvdX3bG6qCAkIQLRcYuciWe9hS4FhezZW4ylfVO5GdXhISjPnCVjpb
K3bp/rhRD43xBzifdwLptQfeZqXGlG/x5RTVCxgVionLXr9QFGNdweqV9ZlKbndHo76jTEWILCMw
p5Gp6y1IR3kUoPB1uf6YaTwPhhluldBGb43z8F4CwoHUKsSrvnA7dgDtXxOK5f/i7OwaWEzU0Jv8
lg6WXu2TvdSvAuPp3asKLAg9whJg/mIh4huv+vgkrhJ5+T1ybvBb4/jAzuUmHfUzqjXtQxheDgq2
4vs7cFkJeQ7coinrfmpr2ZjO5bWtYwfS6mI6b5+1tZh1CEd4vu1H4zlGT7KPWfMIbp5b0myhOzHS
UyfKPzoIWKanvVUDiWdj7/2DaJrzMmaYTsQjUEC5aN6dhif15x9MxLSxaXcYfRee7r2nCUA1jIdT
WKtT58L6bADkwEldOtWxRjxVcjxvBjVjWAf0Qspa8bls9RP9+Oig1FDT3wBRJDM2WohcxiBbVgFd
vuH/qhDx85IRecPNNqikI5sYSFjLiyc9BO9YJ4vrrSp/Gxs2XEns7hrkWC55uw84CDJ7xvHtGkbU
BPhAp3NTZN9trJciw2bKirxoiX8GZgKfPNSlb/QWbNrEYLcsP2qg9LykU7rAh54MFKyf+LQflmnV
GTcEE3PyH84Tgedp7c0oPd1XEJVPR5Vu3sfdkgyTd3daurkAtUfawVD9ocJgV+w27enPSxWPGxhJ
3t9ByuB5loBZKEBb2ev6EHC3F9WuLkVy7uuohbdiWIiI9pw2kdtjPqcHhxpvAL5dBkindBIkssti
w/FtTT0II/tDLnBI1DjBvsiAgMO9LStHzsjjspYPuGZ5ez68aZcxefNnmQId1fXfXsuG80WmGp9U
hldwQgJVy27Y5FgJUaSSsKm6kaAATdpCXWFVOHVW9LNu95ZAL6Q1K9NVSjqZIZjF7FYET3w6UPup
31JJSHR1rZsJ03Ctq0siUHJ44zdmDRoYxzHqfDW1SHh+qjBnRjYYaeEUrvPik0hXxLjn5Z5mQIT6
aqC5uZUB5yYsv4fkWTXjvxF8H9Y/jmgxpbeZPMywyogBGO1t3TVWs72PnviDB1cYSFPGzgYpuwGx
t+KAni8QyrV7n9s1rJLKAn373e2szqrUtboAqSqylbEvzMsm+4Mb2jEHzfJiO9fYzaqsK6gjmk+W
P8zODXQW/Vzn0Th0p+J38VP4ccN1B7UdkyfM1gbznDEiLFZDDDntpFPfQgXichQiRN0tvmXyowoI
RrCTcUUuTB3XnL20bXbpeZaPyUHobvVvWZPDnX9h10GJmvGGKVwfFnRyntO0YtGoj0fs87RaOLHc
YUd+h6ExQMPtwiLjlKcirGtxASpz1vzjObRCpW6AcekS40CYoz19WY6liIU4D34VPDiT6HHkZ067
bRYpHfjcgltp4vSrXyXPIDWNIB5i25xQR+HzG3CTAJxXFeyJWGz35yG5gphDqv8te4A7Lcx1yltt
9CPVPEbmn84f4A7MglZes9gwr3rfi07RukpbJxalmk0hL8kvRDY2VyZ9qagpZVgbd+vjbR+8g1zB
lW6dbJx0FdY6jqOkc68eXjHi+H238Smn7dG5k4POh1bFV8w59cI/F4dAj+xwouKEpgt+rhjsyoj8
bUEbs0pXVk/dGDz5YJk4ED0UqDkcSTKlNYCDTgYlBiFvesvCh+PonCyR0X1xKJduwTacdPDmcUFX
Q/MoHABKqnE27ZqQsuuRE6v8unXeicPK14BGOusjlm13o663DWIkE7iTquIzyt4HonxPJZh/SXmO
8oX23wsv0DlfIjZ81imSI4mx0z50/nSnvB/So4NDYZZute4T8r6sia66liOzeRcS+3HRt0GoUQlt
mJ/tloUekhDDhe8/m6E6lfJLufURE1BNKafikkzDG9Zou6TrxxRgeAoOAUiHkI2QIBuLa+8etO24
roBq4vl8ctZ1LFber0XrJyg4G5Sl9Z9zdNgmMzD7YiU8QUWTf3Gkn1gbHoea+wx6eJbTNycOfTnG
YMJrDS/gyaQgx5x+o+M+3CmovQOXHflyjJUHP6Hi3VzwiNTmdjB1pY9iYjgoE6WzKP0UZirNreCe
f5RLDWJM1Shgr84pUoBjCxhsZEOWvDgRhabiD133S2A2IJmLtf3T5dPY00c+8l/Z1iUMBnn58iy+
jEH1U6pmON7H94febtHtkUmpkKMsONIP/c4YASLX/UNEIRvg/1nE1H/MMIW/8xP+Oi0JKIbp4afM
3StuvldYAH1xtzkjCt5azRQ98DMAhOpc6onMySVRmYFSpu+2Q9yhR2TKoMhviZN9NJgCiqHu5zBm
/o+jJ2eO1aURc+m47HVKnN/IXmw+zaG9R2HB4/ZsSzuOProG3cSwFQiq8OBgg1QryjwpWyJKw5LL
XEsxVFB7pRUJjCgX7WI+ERqqCd4pd91sJnrj3N6qozzLEDtM0XeNFo1sD476SX7rpSxHeKBuAzlX
joa0KYt8fFEb4GlpVS9dFr4vnT+nI1dzW8W9ByT6hLXcd9elbVkxvGAn6VQCeCruIFVRR206VWQZ
asnhHJw61/MtB5wTNRYtmFN8tRiS9jmbcMWlEAEfpl3CdTQP8n9ocZblxDrEbiEH6RR+lcTD31P4
kNUxsNuyWQPW/a4rG5uP0l67gf/rf0VwNqZbFJaCujy57hE1CfiznlxOR+9gOkROmH7uYHiNs1Jt
5B6m4rPYA48KG+uBpM1Rcii5CZuqAmLu7rFbjQzGppSa2L8onxzLWsS/kcgpZztolUlBmo9Il1UP
lKJnMjXM0Dn+WVklRI6erMTRQHS9roC9VXAa1jWvarmjlO8LKk0KlVNN5vTMfz0r/A6MqxM7qR+e
4kW2zieKXs1OW1oVEL7EhHdKiTkkjHCSzI49mITAxO1KNXyeb+68DZuRuB/zfVZsI+Hd4TOMl4m8
buYc44IQK6yiejOI8wgsApEQevxfVuusmjfJMra5izPxN5RrWikR+OatudVMqaSoayTvCFYrdRnA
o/2Cb/NQKMLQJfDv6lCSYBuCXAa6sUV1zouzWxCyTTVbIkaJDRmAv6DzudXkHmUUL8Xej/Miycmc
HJeXDr3sa2EvVDW+ow6a3CD3Jrg2EDamD8GIDP4As4GcFIDvuheLDJgwjgSKBrHbYIQlymITVMf7
dp/DT8JvUL6aLqFjKrZDb+FdSEaP+vrpJyauGBssPL9oSsTESK+BJYm5IpvDL8drD0EsimcKIxsL
/XH0a0IXKwqWcNxrEyQi05pJtxFbYZODLgaCQWoSTmsAV037AIivktntiOP2D0nCSz8V/4L3YE9Z
8p8l0uzp3eIHXz4uFc1GLMQcKSUiP66HAwpWPjmgpG40F/L+LEYNiLWORzFRKT9KNj+umneu5JnZ
npz6jDF2PVCd2wvgVetKADhd+NOhsxDEahcAEbGgBo6qU5RuWkzuIxVXG21vikgcnLe4l0rNpiTg
BriDSf1SAD//iox27qDn2pz5Ppy8Cc8a0G5/VSFLl2Hj/c1p1f53Et+dmPpMGXZj1aP/+RCmpaXP
e031i1co9FIyN+ovzEHIJPcJdy+90Vn+hHs5HSmol6KIz4rXGvOClT27MaGVi1bftRmzcowQ/YJA
Re2EvwlIzQo8VBwvMkRE56GSxg/T3sQeH+foOT2NTbsRm+B0yRCnY51dCfs8efRfO5DHDZINONSv
79vb3JZCBeNANBoE/H64kkRNpnYueBGIBR9HvR6yEAbSO1liHPEK8gqyxhJwxVWBq3oYiKrWQNIS
vrBB4GmIZoh2vS3pNx0+7khrd6qePhJwHoq6EIYZuImR3XNaWr4UgNwCqFyu/jumLINC76bqwvFU
uQNTxCtK1V6Eqw76zPv1wD0a9fYBOltqmYlEq//eVIJhwhGSkNphMbyTWBUUaQv4Zo787XlmtSJ7
+6nKpgw8Y2a+WblAkU3IyYS85868xEBiAztSQwGDDNTYeZqfjG0EiOrtrt3xnKFLK9JvgsGiQUAg
/3a+s7k2l2q/DA6MM65spejiEpXdhmdUM1gxELffhJVGzVT7b29ZwQZe7yJ5paJpqHX9t/dir+2o
wUm3AK2vKdk6x3KghbjfNwwvJOjC46VuoM9uLiA8JZFqerqNHT05E3oNK7uymzX1HR9AtstFCyUo
Tk500caILHND2wRwV8pL7xM/jNtxH+h9LgMA/ExY5SiUW1h58DZzrV7q3HCnnKSdB73C9DW0y6o2
oSmCPfLYb18/N2rhsry5BIyC8HJzF7xrT8vBA6pj5arHx+1DFMnZ1er5DuF36W3NBWj5ElycO9lM
4kewewftVHZUW2GC5qObD2vrMJnyVSeYc8NHs6VI11eEuT/mXrkA7rhuHnOOViEkatBtbh6DCeX5
Ex0ma/t7cZ0iAasg/HO8h/ufWcXdOInsQiCD4i4QmDx2kmFSFzBhnpMcUmc7YQcjsmYlhWqF273r
hXMXq1mB7Bw43XP4MEhmc/Na7p0klS89ClKbxW5A+8XnnKqQNig0Iuz8EJYPshZsgUcMmUNYQfAz
4OX+8cRSuRTrABeCLjmHTklWuTi3OoLYp/FHiXshU4rOy9vGKaM/IkYDQ7htyqTs+W5nzngkEhGt
S/HqvU6/UJniMNsxcT1cnSSSxLI8XGfLU+PuGChYRHfDNJJS1tpQubThqLjw/Nt+rWFKOGW7z9OA
5qnj8SF5Uo0U/2NpQIJyVhzEHcoAxOOQG1bK7ONbYrNsjTzep9ts8aBI6leA2vA3H0e96e0IjkKo
XUc42HI0VdaTbZTktNZ0XEa90A4ygSsm1MbZtUFscvz5RFdHlI9lWYQ1T11qXvJ2ipEUqTS6f80r
Bjp16FAaHLaQ8bB2raJ06mIe0SLAMVL+UZUV8nln18GobOiaNlIPGBIVyzuz30u88Kt5aS/4R3DV
mSq9I1wUxpjz5EtemGkT0VDAMpOZBw3NnBe3FUUbRgoglSw1vVopSs/XVQ2C1JUjcrKkJ0DRAwGV
MNMED9GP6d9wyW9Q67qH7pwoKdtNSI4edlLTL4TQB75w2TcO3yNel/+kmlbKQKVMjdcThSnff9Wr
wDS0lwe6/9FUf7mH3B0el8U5Cuseevq23I5+BzojcUitCK4nhQXL5FsYRV0GV7L9yZBFsvSqohgQ
DFMRpK9kGp9kK+3tRfVOwAeGRMi/LrpHIaFWk5NjAmULOhx9Z60dRDznTQjfSUc2ODbRLii97+Q7
wRd3XEiMBBfdOBPTSrsDIBwyKtvTP+Dzl2zsOp2dLXwYy0q58JdfoCRMTpnxHX2ShZgcUkLAqVPi
/T8bMRSkEYetTy1jgyf4QgaEcTUKhLr+ejN4c/B0UbL8Cfx7kwYjUxlAxMOlYipXn2/AcaF75Kh3
qmG1tsucbmj8RrPG2r/lz1suUal3pKCwNF41i4OH20RhFDeR4rkxewrTmO0cmiECxWcB6RptIfET
MAb1GRwfu5Rf2LOl4HGiGncgv0xZqwrVlwwBs4CndU/55vs0TwhDP/m09k7rJB0Cn1Q4OSJDrhoN
xEgBP871SPe20KeHvfOisy7HkL8u1ufSiIXU213bQNroQ5qMdln5oALQtdEK3fZg8AVlggPs6OuI
FtcSyyYDhLFo040jqBrOOXNsjaIfmkIhyVkK5G9x33XeKQtpzH5eq5iUFt476AoLY6fbHHmq6rcP
wo/6HMLSiFybbDhVbl9PkSIl+VL3s1h6Pp3rQk3+q/n4pnPWsYI38GOu4Uu3RSXwznjUyRwzSsPn
g0YEffBpH0ZV+qVP9rV3dCUfteiJSKCVb6lClE0pwp2ITv7K2SF3QLQVlTfpj1K7/zOCDPi2SWNJ
/C+p+hZeI6s8m4UpCMJdHgnoo3IVAuvKvTFdsUBbCxd3Np5vdgl6XL1VyHamhxspyl44GClygJNY
2TYG8QiQYR7wdzz5q2vD6xJWtrJ5KhqAURSdYisviaABIPexti92NMQUFe6GY2ZYitNcwmaOByyn
dgcuwg0uXoOVfNgaGu3jnks1GLqaEK7lKgGzQ3+q70Bkzg2DxdcJsXbnlNxYKeKXuvIqQyXIWc+3
dC/RoTl4LWt9eQz+ckYLYRf/MXOXlpVtVTXfuLQ16jdcHD7SkxVGRJWLH1xmPRJFTcYLjQrW1YVr
j8rXpmcrYdTACpHqdiKC7p6qAWexzpPgtLLPbHdemQtr/zCoi99AJ5dMSr0aRvSqghtRxzv9rnF4
ki1z+dkRHpmHvs2kLJ3FoS1XZ4ZHmmcr4SHsbqGFZQOGVPE1oix9m0BfawX3nwNLc5A28kUojQlf
YBJvYxmWH2XL+UaiYXFS852lFrXmyjxhjGGm6+sz0X2ve6XYGRVaZP7wp2aifxA5QTfHTlyyjcZy
nR2PmZby6tk1fRyWKunppeS9Wbc2nE4ey2vy2qcJqITNttdsknLVeaBKZYCWNg0ONy5Q2EwgHY8I
maTD+S//fEo8HLmi4aDy0E/rFe0m8zqX2BtKgNj1xncqff3RC+P1oVTkiOle9Ks7FZLPJZ0l5kJc
ubgqkWd1+k+3fPrckQK/HPAKhWZMBGVI5GklA21CxEhbLaL4o3ApRWDYKAjB1VdmnMn83gLXU1vP
5q5k4tQVKNPreXXAGsAxDRkIGiQyH1rB7pu/xChfhsGvyANEGatGws738DOpLKNfyO2zMB8q1bqM
gYUfOoObvNrILfLtx6tKy+HRv4+vlUNg6ehVr8qYZVWG8L0p7k60J/rwRbTzTUYl0BP8ZZ4TqfCu
7zwwPbQk59rRsvmnnEEztwWDpvqAaqLhxivThrb383bOqE5vO7KFaEXiNAc2Tca/GVTKtVTqMb+k
hxdnyCyjNOuvCnt3hbKznmRdXy06qIPns8Zws22SxCDIwSHwnbEIprXbtlmmOYs7Gts7vbO3JNUa
tf/RxGYGhBW1b4yeDX+DGNm3VrCgY6RIv9j5DJGMhQHMGNhU2zo+q4JUa+VybKgQ9T2ZOroRYyow
VwJ1G1/EiuXucRO/5mY3MSCI2Vzj9nwZOasYlV5JQ8Hdh06IyCj0GNY8saYhtHA6qfjIVLKMSsMi
h8zTQyOviQh/eqVW1WfPMYc362EMx/ixFcvuYFhUtmH41nLzzHWrLK2ClyNrDxWWN6opEZqqHnPa
/kxRWYL4Q6fAGn42HGHyv6ahzsfIGxd7v0QTNWdLAp1zMyP8Eh3D4JG+bRGPPL+VyUwKjFwiZSe1
m+lnENfKRWHeYcmZAz7w+Bqje44/kNxhMgM6gn0kpuUbRKooobDIkwIxPt1zj6Qsb/sB435hwSaq
VadWnNoVVkom21Y/GCFnsx0GZHhcnwBID3tR7434wRPKc2S/wl79gmb1g4+lefW/5WTsQlocFpSv
iMj8mVNIbYdsjwMTJdPByNgFit4yX5uxSI06o/K0pgpzmKwYElaJqqRblbG5xAa0gd+eVFtYR4VJ
UnUOEs42QGBORkeaJMkSjfsS6K3ZD9VpVXS11Ufg13cp1q+AZA6r+43Rk4xQieef/uYW+4IXQfQD
rEHJQL03ZOBzZzzgtsVX91LU1IupJ6PXgZlHAflViyug3dWDVn0K3UaV/jPDZz3VUsWbRE2th5bb
a5uCud1Ji+WmsaveBCYbTW8R2S//vkgRZZL2Rn8PtVjjV1D5Be+GWxZTWAuZBXTowOr3iTN+5lFM
8BzQtV9plGjXLk+93j7ebZ8dJxQuwhWsa7hJNA9VStrxLUiXxlOquS8+Fti4pqh3BxUmgntMepuU
jGMZkMXaeGP4ZbasWFit14bHenq1q9E/5GcyVcF+nc7yG+uXr3hNSaLxDz0uenceu06P0++UHNgi
Gc4UzpL1PW7SKWDHFYJBQkvsHlsu45hmhjl2uElKg30UMBSXWeK4gMn2UCdWUwcMVm/jMJP/iGjp
NzWdFSXb86MGVQM0jjWEgGuOQAiQwt+OUXDfrPIN/o1VPp3qgeZos95dnVVLujyQ56oJ+T29TczU
5W6dF3X+y67HK0r1sJ5ASpuP4m6bxNlVG/8AEMEQi+zJUXEYoZvzdjEtOfzyzGn99y6goq/r/Wmo
WonexFZf60g7xDbJApo7XUkRQfzTN6hNC7+ayUrVa4wxI4mpOI0Nb1RnBcfmW23CrBF1UH+oKoGu
0RdX2YKSrno5LxuMGInmc42EKvqdWq6tmUw5efDEpicMeEvYl+eCIPr8i9vkpFgSI4UIzBF/QwZf
Pp5AIlhcve9AYk/kflTRS5nJCGdWR5EY5ksMwvTGvIL5OoGWk70jLUDjSdGfO5e1SZYeEkMAfc9d
kx18Ge4Aj7yevrDUCni/jVtoBRFk8hjQKr/jThnz6bWxv1EhSe245uGG0vp9oshC+KkAUknAeHc2
xtPbD+tBAnDiuZwTWP26WEX0wframywc9ANmSUDPGkjlb7tTjw8sT+/ax5BC9rjgmkYTsLvnrOzf
wD8BSpPoqr839V/20eE1Tgwn2JNvJ5txaUWPKuxpg6JvFSgpeETMkhjd0QgQORMfRaPYOQ97Hb6f
L1GoHapdcCBH8P1vpjfSLsAb67fcvpH6Fk5tsa0Cssm6Q2mgNYER1kSr5hd0tlF/Z+614c0yNLUx
U9dFhpFSS7O4KBuJXeqL6mWg72d92Zx4ojA328rL54uQsWcR/PNEAGn3eXm7hYx8j2i+8PB4DjkJ
l/C7zvAoPiiej9RJFptdclGXfpsrTJDreWovBfrYk46XmJuDFCz6z9WXOgDjEENqWGHhEqoViDK7
ecZU9TrEAiYfXpODioRYkjQJ2Oj8w6YTDlcYVo/VXGarCs1ebQUpO3Xivdk4EEojEk0oG66SwC/U
2PCMwFX4PY3ZGF01SiySFZtv0qhBFE3Em4XxJFsZzPBX50s3Y2G4PjY+I2KTLC4s2ywIRTk4k5LB
Q0X32vx/PnIZ2RSJGfQqUiKfSlWs/bbcKh/LJZpCBTdLCr0d/ZK/obyuFhG9KO6MUWcCxhOl0Geq
7sqVnjhltplMJ4zyRzc2If0tdFc7UBd7F9OzEmhzxKvTzVnBPl9EpFuffaraaFhiojQYekFAWDXr
2+v0KCB0QkRnRK1pMg+ycsXz6TltXja8REiviPDvs1PhGOHEw4M8SiOrnAXm8UIHauUecOqknnAM
YonXJ9bDUD7dXQMRwdv2uhd7mNh6p9F+vLBuYyKcWD8L4dgW36mDg1zHwjQZRKLS06QnyxFyHkby
BUm2FxZ15bv6diXt2SnAdV4OKacsoenvjMp1BgOcgkOiI030VhTAf3eyrNFyo3TTHbZ4ypo2/d9s
uS26kvVv7ZaFAGbykPaAGGYXn0Z9WvkPbvQ19jT6EzgqrE08Xe9rZP7dxy9tnRZskhwLY7R4AFZf
Woq/iVEXwcvL9u6uPc8fWQtOcQlAWsixIJb5Sr0VcAn+9JPT5REHMKZLOjQOf2OvwuR1xciVuCdN
e9NuEWbfPD8XtLaYhOslPDQeydTbi5QYR8xODuulAn0AR5EzBwqZJIreQU9CCgQ6moC7gMzzd8fs
tpIKoB2ZWe1PpbxDjl7R7KnpcYjjfK6Np4iS80sIOb/Gtdc41EMm9PEV4HYc9Gp5CE4nFJiN1Sj7
Qyw1uPWSSdsMUTW3N86yhNxsW6bRlMlOz9ZUwU5d7hADl6sipLlvMG6fZpBjo7RFNK/J5pewvu9p
AF/gvr7e/i8RxTSzHi/Nwj84DuumdZ8ouoNTMB5iWvS7qde+dxTmqs98dPBgHagYuO1ObeufcxpL
dolC9eVL3QRG8+c7tpmb1lrDQ4g/64H1rr24X69PvPW0bc3Ixq5ca60vUsKkOXJ1d547m/ANmxY4
2Ldhr+IwMqRRjRZKkmDfhLC29xu1z67xJw9qHMOBaaWVZ4UusFSdcHy6heJ41ndcfT4yu717IhpQ
lwx8dRlbkaCvmPYT+LGmviOw9wT1bPGazAIdYLuXLAUhRmZ/GeaSTmBBnSWJ/Ub2AKNVPBW+dUOg
aSAxMU7Rk2DfBUDTF2W4V/pkfasBqRaIVYhY8bs7yqQJn7cWOH2IpWj9clRkt8BeKJWBa5YqZ56s
VZgTlVMHpoAVxUs77jm9nf6Kbvo/kDthouwbnBHci+sXBNN/rNjQuPV0ixGrQ44zvtJJItZgJk3q
XwzQB+lImLvVGvgADdHufkUysR2wvOibLzr+BFXhs4H0oLI9dDu7N83+31MltrOmX839DhywTRRZ
P/yukFqEEHCVbeMBoMfCvNH8ime445A1CetrGZfoCrReJbsmqMQEb1jySn3eVqP6XD/mtFg0nI0X
UdWAHo3stQxjct0/mx/9RyBeGlzu7ceeM7j/Mtq9QwDfQp9wARZtchMvGekaRrKafI9fqQkLJYip
xxF02nv4di1E+iD49NWbsC6Z9e7BFufhdanLFXHiH7X+H1EEPduG4yX/tCR8vCeJnXFprHbkoDZS
iXSkmMCOXD4Jlnh/ax9CwLKbSsmrN1ntbtcFAZXsJ67VbYOgZTkVQ4w5yXuAZHIxGFN7duX+yiDD
zgRGJDCt3exBbXw2slC3Uc4MWcazV9TXckItRdgggLGpF65FQ8NcLE/egk7W76hGTCyz+aiVLF4e
s7nY70AsVK02g2ccvL9r6VMgGM+Kjf1moJyk8rx2Ga35kZjeu80c9zsWTcAk41NYbya4fFutl0o3
c22m0vw9iqm3USQX/vgvbyvMJQnPbVm8ySNPWLuDCRCCCyThdlL7O0EB4dxx1QVdXJcnUJsETVyp
RANk5qY53RF/uBpQGJwXI0XP+Php/xa270RlI4NQvDs/hUkOmgcRreojUZYtkuvIIEmmhZz7mcD1
D5euj0Rhh0i9keuoryrvzxG1cCdTvVAtlLDlZk1iMPah3B59fKu6QAe2dXqq/FhhTMfPLPF/rUwm
oOAwoA6idQg/3rLVnGJE1Jr3XeRbg9mcPdqS2cXj7kH1mYqQTmye783SViG1TBi1MiZfyhsXT1UP
qqG++25tCQzWI1Le7ZcorHxb1k1n3EQv94DMVS3PgIjuLQE2cY2wcKUVAKlfOd9p+hZeEsoNvUmY
f4pylM1opkgcnWqDdoAkf2WKtDqpuo+2DnGoSkPOxTc/m8+QXx30K1x2CqeDjaM+pQPQCIrcQS1q
B1wo68cyIvNt0QwtadDRA+DFflVV6akVHpMiNIGxbh3Dw0BN4qwFpy7FmrgpDOsIXIUahT/wUahr
QPbWzAbjr4G9j+aYTA3DEP+U2miToPL0XcwZ4Swy1rTn3fk4MZRCLVOzxRx4sOpVvkAWZn6HTAnI
WaIFt+d5b4Tt0OfrHQX99v8Wc4JfZat+Aoy3sHkH/D9dJm8fceOX5NshFGc8acbur0hXsrWgeKMN
rPe1U7gI/HHp2Kwv5slXVFjnd6OSyLR0RzyuEFC8eDahbu4LpcsRfGtZICHPdMbQ8ipu0FlcpLL2
Bl5sqxcjFTBIpCp2cRaZ4vCkgPq0OZIft8WZ38ZcxnRU338ySz/ziCNlABprVmIX/AnsMvPyinSc
rJaGeZi7iAKAgicDG3YktpZfGRUelCVZd3Jp5/1xpM7UKzIz38AnV2EczhdLuCsSrrefifKtu4k2
P9wjvHFfHWS5mJgqAW26Q9H2x3jLW40Zf2DetoBVj3bNWjotkKImBQI8B8diByVv2n5/0JFuRMC/
bRzJWrYOuuwGIktV3QtuVEBmxszyoM3IU9x1+VBxc4gzERv8Ay8n680XLAcW/IkwvJYTr0cMyfxv
KrB7yZRrbNS8TDPi8qPgJdWtR5MjsnMUV+SsD3B0fyITGp0XPxAz7VtjJxhi0WZEvsgvyHrhZq3H
Gr4mk75FDeMuvF6v51cegV8KXILgLGK234lM2D/v6OlsJOPd+jj4abLqFk6AnLLl0cfTdjI5dO8Y
UYcSbNLMXtiooWa7ODvz8hVXkzLyuIyadmkn/m8DbWTs4ueOeOJQ0JXPLByMhMekRs3ZGzxGqMba
rqHU9MSzd9R+9eWB6mDgZ2Qr4I3Tmkbd+5FOs7KW5IkEvCVfaQvuRNmd/ggswymwfaj8IOr3bcig
0xs6sZmr18D8NuePzfibUITRNLTVBgZClsmBSnE0ac0Dm4Vw11GvVlNT4pLYhR0ME50S4T0YP5YL
sM6D0lLEbSNUXcC2wgeU+fUJU1EtkKwJrF28wtXZQ6ic638l7+HoNGKGjohX+WzxK/wRwt7mPhIU
8bv70k/WtZGWYyxGVSBcVelg8HrOXDbqW/6JA2DNBNL7xuoP81nZKmEZwT/m5Hd0Z+qxRWVvoPT3
q9rWCfoMR402MgOTnAL1n6uvw3VzGG1nrOjtPoYqGaJ649lt1bEUq8e8QEz+m2xHP2hw4ogkakkf
uhiob4oXoALRdNEJ6C45XoBlNJSEP/lDHubJ93HChPgaVveE5z6aEpoZ05JwuFyZ9gvsDZpO0ru1
huzllqZUvOgxottAAf93wg6v90R7lR3/wce1hHeTvfYOo2Lwum9tmQ9+S/1Lu6wXIeVpEN/AWfoC
MbFfL1EBWrmGfEdfz0m/6ofvtulQQUbzEcn0CNuE51qFMv6HrgFpjQrqczJsfBJH1uEqb3Ww8Qwt
iGihd0gIvhPb6bbcFB9wOI5hOfMsczwgQ40oXW1CuC0Enm9grpDg+VGU8Zq0QNpi5+bcY2vK8RcL
pknpunuBziggUKjrF80uQOUwjM0cE5J+8cXOB96VDFLPHa/8jIbj380umznHX/qXeJm06kNjjkPv
V6TnniuIOOwYg6TU//upYuZc5AI30gRnOcsTwxYAw6TRYjgsuyLk1FZJXKfRJKZUarBcQ3Lw0Gru
im/EfwOesfnSIkLIM96Qvn+SzKLpHRst3cSvWU491XtsempRtJFJUmZlsYxrT+IUzpeKxuoQcQ39
Dlrb0hgldvRgVQqSPUAnKeQWZtVgETIX0i3M+4pCjRV75K3a9lpylTk5rBFQz27J3RMXjigZzWdK
DuJ7p3QWiPJoSlyqRa+7V0gSN2+Odw5nFvhuMAykgMfgUWhasBaLQAzuXzcmDJcW4cb65sE97WW7
obAfUuXABiZi8vx2UF+Rz8DPDOsVgGrCgMjwHV7VVT1jc+6Hwaa+2sAxQzXlYqjBCe5F7jeA2OTf
xmFD7VBkuaiX6tvjIPkdlG0N7ulm3KvL0G2Cg5Okpt108OZ53Yk7a/ZqU8M9ucC9k3kHgmwwnrg3
Mami9fNJL7HWyYp/bo3FK9ywryr4GbmOY48qvik0M+cU40TXlKTCdu8a+DkS7+SUbdL2Xp7COStP
32BsU0Wx3ixfSdsRRycV0hWHH8U2131B7GvEhEvkJi7yOMM/YkQVjFBEnm6n0D2+V6dLf8saAzZE
hcycdJ/p/JmgedH+BJ25IY5tKChmr1RhknjkaOVL8g+XKPTcJ753U6GfQ+KZ5621cxGMa6Ot7HgC
oSW8XAC4CbUlyvVtB10XadWtFLNgC6h9LpZcxQrivtOV3gXaXNK0WoALlsU/kDBZriCWchBSj/wi
BvZZvInEmN9N/GBT9LM92rXsnN+xlpk/5C+zAsSo4u8wHIpIFLbNfbOpKdWkqhII0rt6ZnpXs9rg
8DsfwOf4EuXNJaJaKjXOQYEB3b+MfiIj3D2eiU7H1+4fRHBnKBM2RVE2XZDaMTzI1EVKKen+PvIb
Ai5LQkvRt1AwECG7Y1ApymFj6sfbE6VWBCeRTGmTNoOhwkKgXK3jkjFWh65Yw9GArQtvOtwkovAE
6x2dd2qXRP3QNKm44L0+kqqh8dNzUZ8LYavpQkV5juSNNqAYWL6aPsRRNTaUe7Q8DFNTfGUnFket
FlLFdwcDdfU3Lc2M/uuzBfArOh7cLTwjMTR62H74V5ARZRUFMmYsDAcPuskqh/Oz2qjr12VOtzPG
UxnOMKmnmE6mVwI0Ehou/pnhQLKiPrY/HcTAy1FtZWvL6M6myATGq/fnJGAkShCeybLYHJPzkuFC
h2cGsqtqife4w6lEcsxhibxtjBtPN09Wrm5YA3q52/7kFB4F399R5tjfs3mwQsU2l5PK7GpcfJeK
jhmnX06zcZRoh3pBB+c4HfsdgPwmmMUCgFBv0OyZpPJ2RjdrLLE8owU6IubolHjDc5t1tIS+SBqn
xXGZhuXaEwLOKC2QbhwTRS2vntya3t815mv1A2q2z6rYyW6FNb1t6VMXMG48+rJPrZeMzSo23tWH
mY8+itBjdbCt1rohYEeqbrp4Hcx3bXANPmgo61od4Lxr7YG6y97TTZd6TPbgV9fg6/oQQWZw9myC
/+BaggtGg7NXnhyZe+dZaGSleMCk3gIjdFB5gkCWy9rIwi14kAFYkvvH6biGn6ZsaF2hSUqfxION
vfdm97gJmskPqjXqhilJ2zzCY8ptzmb61ElcrDBEkTsbi4tsyHIzlN2veu+KY/CaqwnwnWVBl6PE
20IZ5554o1ho7SeIu8M+I8RuYyrOgN4fEBfjlxHtI9l7CI1sg865BJ4pzXwrh46lpQNjxjXmeNPJ
V0GfsbTmRdz0dGZJU8p868t98CB6lKvqGYTWzw9F7VxP/sQ8UC/or42yMgjA3Ws9e7ZQVU3jahys
wR7BkxjucvhbhP1RoEhtsWhHKhOGGXaF8W6v75sOBkf7cLaUvYk0hAkXS0wLWpldE9qCzIAJegZW
Z+87PxAxSDZvz73fD/icwMQf9G3pQfp7Nb44/wj7AvtF0YIhvD8p9kGOJoVi3goFGIWR7p/tt4n2
3kaX+vqhrBVSQvv2b/89qHkLc7BrJnVTEWUqFjnoNF+YGgMqnIfdnJFYcjaIUZnXhRQQnGRBtSi6
BhmuTCuRy2MUM0TT4XwqrsurZ7J1BT0CNhqdM6HfaVGFGByLuoXIi+Kcw7DQILLojREn3WmXgrGH
KRbU3p1/wMHnRe4NeePLTVO9r0TDUjuW1tBZ/pFzuajLV03O69V+JcWAN4hDOUayb4CoyiszSm/G
XY+5Um4iXfA8AnsokNeozu7KX/Yx2jH3nY64w9TNG5rgcB/qvbwNqsUZ2+Xml1sXGwelRn6GB8JP
TptPg7Bqnn1QwdoXmGNBZRRbA2UpE+1K5fwKmz4SSzW/UKHsQpOoB7eXVLXZUaBiIL2iwqZQdSpG
RgEZcVizSzVBJLZlfxzluqzbgoUv4BUdaCh2U6t7/pRiLjGUDB0QanZ6jQM7XSGpm3l0ub3T8p0j
UJwHifPB+3+RumD9UysgDYP+JeB3GZ74zgiysztl65NviwkDacbhOPZuv/IPl2ZtPdjHvsX3HlOG
0T6oRjNIqk7qYOkRLm07ZtZpvpB398eV+oWyBWrNQrJPcE6I1wrf/3XjATbl2QGm8eAsm2e8LBNj
T+VqhOPSIa429wi76KM4YjXe/LXcf9MW3k1x9/t1akH6iLDKRqKTxtJg3zo5XW8TwmN2g6WGWM2e
7/Mp1XnEjOebuVnXn9s4Fthj1eQsdhwsAbNJfpfM/GlXhLvrIx4wiBOZLlGCO6WvgWLkMtcp0kYE
uaK4Tvo1Kxgxb2cDPzOI9oN8FTSjLGFKtpqGmDHoQMQ77qwcfGniY05c6qKy4E3pNlZufBvKOtW0
ubVE8YLMUQ7e5axTkYt/KrhJ0+0TsNcW5cuFsRV+E43zk2abXCptVeMo9Cfpnfjt71qNQyrbz0v/
iK9v6Eyt1gngQHT5HJKI/34lc24nxjt6I04GBh8ApYqEvvRHt6R2Gwwf5oi85VnFy6/BnGOjw3Pm
+VbXlWh2ZAG4IW80pX+FcCShrqbBOMPn+7IBzEPzgo9MPi7n2b/tjwZz5gdNz0iBK+yzBhlsE3KD
pBzY7T9jlQW3v2exgHCsuTDaDR1YHwDGifVIXTVWTExsHcJkF4pZz+3Nxz2E1HBfujttU/Sh2fuJ
RWahiIolNUk+MHnJNKdVwJ8itc2EtmyPQjTfQY+X49r6+DWOtTPxLOHKtNPAANJBRf8GRUPRyC4C
przPkNiajgeGbet6JPh2581Zc8x63QRmQO5qrg5RwQFGeL9uvK8Vq4Uu5h0OA/F5SApl4bwYd/Bp
7qRbtsQK1iDReRS5zRxP5Zt18pg54yae01/rK9kjvSIqO02IAlIxmfF8zQfD1l2AV+q/YJiZcUv/
lIlRTyQugU/fpFdE6dQLXu3GDN8O/VyRBTs3HCoqqhUB9NCOUXT8MGuV60Jwjc9cWx8fAP/3kN5I
BQFRZXzMuUx80FviQPlrnCH1zeneu5APdbyxU4Y1Y0herGr9WuT8ihUG9aYtaeCw3zEHe2CntJHJ
qPBmLNbESFcGpqQHc7zk3AwLPTOIqCZ2mgh+3iqocKXTjvMzV2pY8mep1ss5kut2xOiliIJv8HcI
YE8LdpigTFZEZ81E3TcUbx3n/d91ga+cqvHg7dUvZFxLKBn7CIsDj7vh9/9C7Kw2ENfHzPX5i/0c
pbZocseuAy7vzy2YIW3cCBBfs939mlukgs+hJPkZbdvEyCugcmMT4WD1VNmfCQeGvHHE8h4CLyUy
R14I5DM3AighZmLFpjl1FJ5kBkNSHtZQs42w/XGu/L7mirNC9oD9quZCFrdH6lItxgkn9lOkB+kW
XJCmM5eeGS6OLWvhl4MU4Mg6zYJSSCbtsAS9YHqSxdkq95G+Gc16P50dRBkDyQmStBbUKaFXRxaZ
jtyS+GIYhs6G9N324jhtz2YYO882tP+QGIw9LiLxuGbtXOmxuhi2nyYwJ7k8QD6X7kOETjHM5p/n
XtJIGV3HdNBXewzBlu/M4hOI0JuhrfdrOnpGeVIt/9E3AS91Evzh+ittNgaZ9H/ti8viKnnX9GXt
47gB4nBPjVT2loVWOQqBc0MU7RzTqZXKX4oisCHpQUID7A3xEA8abf5hIh69QSKJwcVOQeTffctJ
rsbR2q4OpkGP78WYg7+9ClLy+AXCnCAPmvY+azQOAVXiBtW7P36WPOKByHh9d6T7hGb+c5U6bsDr
GkuT0cpdtd2pYw5q29RqzPmQZ/kYFvQ16ffahtOj34DH8KJNOd6W1tWywehKrgsLtu0mi2+oMznL
7hvwHe5KSaRuU78lTn/8JNf2VK4CVsOcnjV7mWZ0psvefQBFgT32bWINnsy8prUJhubsKPT9xKUi
PRBtb9/K/Y/7sCvO7uOwE5E1VCUqajj509/ZBAk3Vs3SvIiJpS/7viaWvDvti5oLdHLn+e7RrTcG
2MPhQFLTCpdWwVSCGMXo+Q/UoonfsQQz2FFQ/QVzsxLW/VrQeVIW4QY9eif+jD9s4hOwovZBmebq
vQLqL/Fu3BEkXCtQex8BisHG0cOjGoxXjAFetHbh/B/mvxTSeK+OpuUrzdcYjrfV8mlwWVzKmaUD
OkmvnGoFPZqsvjr7yHC0ThjexHRszf+Ur6BGKT9dA228oyC94VZzZaf6RSIUFDkstTFECsI7cN1G
G+NWiawT8guvdKarXmFc7Cvts0QRLnf96HvP+7zYBEunebYNofQz/GDMYZwrj1Nco8FBZ8Ew750n
bJGX05qgd0CM4tVMoj9P0pCqmeo46SRQfZYO0LQ6fPpGsNSDb0+WWdZWIU9I1/YWDXFFLhR9Sdf/
fabKgocgnyvWVj+y+u8DaSqPjGz4HP5afhxR8YsEU4/suXfloRVCHmpQThoR0kU1Y043RkAVxyU6
q9MJPgW+En0oZDiqc9/iaCjIOkNpD2UTJFIC8kqZMqZ546kKm2D/606qJstQDmeGQ7c1zXfn9GM6
NXcO/5mYyERJ7uxjBewwqAbFcTrPc+SvMC3yEu7st7cXbGDswOMDqocw53njfZpO0YRBTLiU0sk9
ys0w05xsduivUDHQ6rhge5T13kcfHb/GU+VdXCVgzRrw9FpFsrZKg7kkSOBiKoH+7LExFZpJM+VB
uWWX4XdjA6vvfOPUVxAFzpFiBAlb3Zpw6FwhnHekqxI4A24nEN/CGaUqBqu59tYE9Kij1HX8hfrA
Vunu3PJl0fwcuXYcdRlPGDCnzOZltpfXsdGCroA3/bvbPLMrgIyl4rSFb202PUgxb1cEzcP1MqaA
LANWLaqfYnWwrk9DDcJ3ZnZ+7AcodgTQHIHjQrsxbswOD/19lWTX1ya7mVykb1WE/+3M+aJ6ivut
dkYt+FyHJTq8/+e3voTDG4leV68fUNL62jGrAk3fjD2YTYxi4Wx2HiiVtHOnAj8Ywdqwt0sdEVrK
I7aE2s3YpgG5QwsfunGLvPprYj+W25zNjuKWU6PE3QEzevAkaE9QIOv16jyv9DQnAqgxlEqtMW6e
1h2SjV3CF6SuDcmA5d+z5KUbLuwOCwj+jd6nuODsFPTmHIaBC0sfsydTvVUJe+/PCeAiGfz4bPvG
zMPlMpi+RO5eEW2wU5jeMAoEjjA8onlikbWtHr+juxlDUxrgnk5PFtACsp9eku0LRGHvlF+wCN1P
E2LT/Pt7vH8Ebf0xBy6DXFknuWxxdg753tThEVAQtjVT/rOLw84zSqhQ2HLYCT6NEC8a8kaIH0GU
ZLfJAPsTENX9cO00sAixw2CpeK4+T6QoWKsiaFOnBD/GW47anA7Sh6kkPNzJ0XJPlfmtTz3Y5Q4g
63bfxyzsMdPfK5x9k8Fvi2KevOXBMQrUfQBWZSxJSsqf02sv3JA5rCh/IeNfyX/hIFb7XBr4j14p
cC7BqmElGgw8QjhuG+tPDYiDVmhIAAQl9dS9Nb7iAQNnxDDOj1gOwZ1SI/XK8OmMQXsb3lsT2khe
mFtPyzKUdJD1kAhcEbC5PZqciUQEAl58g9RFIUX1RbI+WxpDZIlkPimZdxEShns6r38eIUstaDdf
pfe4usSuc6rRBoTk28JS2val/fFzNhrndSeLqHLb2hGB77/osK3icEv8GTS3YSnMpgHJ4qlHU4EG
Zso79IKJvwihbknWTi59979mHspfWzUxqXhnqyawQaObcZRQ5Bsl7r8MH+6v4ZuUgF1SOAcZovzG
RNb0t+X/bLWFTTTlQ9hG4JWnlI3QmmnnHNaXmD3DWOFdu8bXQK2QAjJ+4IJkCjM/AWOR7wCT1Oy9
iAe6zTbYmYSfxQX+XGFkMgDdidmXf+RT1miQQDcaVhbxWmmtxxzr+o8FrD18JSn3Ip/qoJbUKuIz
dcw4QyAx0KJexSTHXSnoCewNuCkYP/F3hvAHJNq8Z6WXl5cq/QWCFrPxFmtOrRk7ThG05ELCAnzG
sMQC6vdU5xdxbEuTf9EqiACDqmgOxHvRWf72wSrWjD4BBy6vCs0dPEEHXmC+9ykoGz9Xbbs3nJga
oDVPBAuut9wKCKEi2S5nbJfcJrDUWaS3qUrba9ukDgW8mc3acZNtf45DtCKG9WdV9tF990h5uLVh
bXWeUz+aRvMXTHqTzy3SYpOhj5Xo41DVPmJiOjfUV74LeadH7H9+H1pQbyuSwSGo360Ha4nJrMnF
0KIv+WFhtvkfCWhaBHRZox6yivklvTxo+pZVdgY0JZvwk0hAELu8/6yhZFCKgrFJSWrmx9uUBCFu
Rw68L8FtDslUAMz/hWZgIayNtW08RYHSGA7zaxmEXV9mul5dikwxxqghOi1iLONx21cPJFLwlWYn
ju8OBc1lkma5Atlk8CeXDCP6fhNwfBJdFvgRldAWdx9b4rX9WbaRo2A9OsX3WTxbwcBgqp4FpYJ5
dwJXKgRH/UnWMooMgBLLqZ/1/rQ+NLY2RJBcDikc+LbHr3gaz8b4Swpa8+XGd0CELrfgn2YQn5cf
/zdbTvLaBX14D42Ed1RiprAzj7G2qg321AD47VHqXF7iZOg1BtcuCrfSpydOLzApOWwr5NyDvC4w
Lg5G5qwOOFgc+lSkfmqR5kEvRNLrII1BLRWVNgly6/ZNYvAHxy3ZscHIsbeKCCQAlmNOj1tZ8FoS
jRoY2jbT+LhxDT4GwSsQqej42qty+d/03pr/YZWSFZAxzIRRncKydcoEbPux/pvPY92qRa/tSqx0
DSgEuZA53t+MDzcqDK7bg3iMAMjojBTfLvpdzKhI6hmz/2UCn6oot/Nh4cHdA8/2KtZRNfXZ71ik
f5zhnHhyxPZv5TxYSH3WFWA3B85+OOtZmw6WG2aCjcXuDnUDKSVEP2YsaqHEQvD2NQ7pm0RFegoJ
0/FRrOAvhAb3lBp21deISDOgsVQby4Y/V3OMcnDkGcbIUqQyCbsGDyA5ZWIUVEUVFqWwqMl1Y4mV
Hj/wprzCgLHWcZv3vhurfnUt4RcvTEQDcJK3UggD/LnJZ8mnCbo+WAY+aOAZOr40LjVmHN50oIFp
mmgI6rP3qg4Y5QzNbkYP5NHphenGtQBYjcOeU6Rm7x5VA4wGKRhmOv0b1xMb0Bs9TxUmvM3/GON5
6j9VJXgfxVGaRF1pGsoqjhheFJHgyeHOG6Q6nTC6BFcKkSG+F1RtzsSJMi1PJWZy42xOtvLjrFVa
2J3SD88X+74H29Z5y8sphblkkc5ohW5eTtuGFPPVcvJ0Kd+xhkuBVocfJz8ai+LoCY9IgxzyPmu3
pdh4cNHOVnoaGieFhKyJ4xJxQV8SPc2tvhWg2cSOxQbHuan/VYsMsL0mqDcz7HJcOuwduFtjggUB
op4YTpc8EMRFdjGxNqYkSu3wVeytIVh6RYhEDpScZcQCrFPl6MQE5Sd6x7uiJC4fu6YYBCqykW3Z
l1/GEeUU1hTZDMmOa1L/NPwC6BBuAjctPiQ0++RAHkA2mYsp6DP+m8PYMcsTpPNaH1i5rumtWeE2
28CysRFkEc3MN1sfkKpOe/yN1i1//JX0UwzbNIo0zPo4sucmfu78fJWWXnaQ0PAWSbRYdoQ12fw2
uWZhKYoabqOJHNb151SAX+n9/T0nqWheaAIFbWxKYEk5kybkg0sjxfn3o/0PznwM7GLuweMahUv8
mfRXkD+Q48jmTO/abD3vF1sVxPBUeu/HnwoYgdHKNMuf/JZODNBqHrb67g/gqLMfusG59dJF3BLY
cb1JSiK+DlGc+Y0kS5v4KmPoRFSllg+axjPcTSpqj+FSVQVJ3PWFyj2n4Rp7FC94kY/OWJ+fwOEO
3E7qVI4qbaw47XiURNWGs5Pm7cIzjHwfcJcZy002u3/RVZSNoY9r8a/TLh2wyCqZd4Zzazzx4PeL
+qO2+YnxaTXXQNJIUQMUfSsZdOnTjvG0Y6rbM/sfjQNAt636HHJhfCdfEhYO6rK//t9WzNgSlJ3X
16+zxRvrQHlWsNDg98Qq9+141GpdNvH19aqPe05VnviJcM0cRsV+4qrAs8VZXvt9iJ6yMV3PlieX
63p3FHvHpIg0ZvHIcBiwAm3fOyUVjiwidBQUjB0+ghWP8iei2tNt2h8c9QWpmwAUMOE+aRyg90Ho
PYMDUN672plI8Nqh2j31rW/g4O9FL0HOjH3wQWK+pM5LdqKhxL4g6kfnUS4YeUy34TZcGv5T+sI9
TYYd38XxnYySjTzKwSg/LmOlEfXmDv0nddIZQAinetzeCqQARNpGYNh31dttJsDPmmcN0K/Pb1jr
9jQqA325/Pv0nl82w0ABCphZ0IhTxLfFmvCImobykB+SvSsUuZ1KvV42WZ7bZ8Ytjjp4GBdNHIYl
Zh920jbfc7wi+2k64qOFH6cUvPtA4Hz4l7MI6zkddY8l4cmiECmRMnCl14JYRpy4YntS5HNh/hrj
oZw+TUugSFGgmKRq2R4BLNPYedmuCoPRKP4kHPIiWLVlMlZtzni7miDLaNz1Py1BUNKZ/ES9W6K7
qEZpECBVhIa4igo6SNUyp12e1nbeVYIYv9QxlJ7ortAJnlUr+b28c7AApvDbqyI+WsueZuhaYnNv
Zd+FJHHXglpTH3LXbbDf2a/cbx3/oxVJFuwsql9fhMLPH+SKfG1by1O6jYc0OZ8sfp0zoy9YSpJK
s4CFnPcoLCVr+0t6yC++JIGzw3jZDjuL9ckU0q7IBRb9piIANl+gTRpVuh/sPmloXneLO6rAqFgy
d9lJlZI9W8Kv+8LY42pc0K3S6NVd5SVelPk9NlXlW1VXnN5Pw2PI6nKiy447w7PGdyrlBVTAEXC8
9wMPMCTz7fLYxYMH/Y7cA4t2BSBlBzTOU9UYsYqCC1j8fv8XIe78RG0xJj73jwyQpYXcrf3TX7+7
t7EFSTaGp3DWHUSt6XPwD+Nog+qLYTQf/fxjM2Olftr9w64cE9Gm6iz+0/f1t576dziGTc50w4K3
wF7H8R2TVemMA+uSPfDAvdF6IrooFBHgVYYPRGh6j+XeJAWxw0tjTfydzGmZEKxxS+6EezlpJtxL
Q0Oar454GxEov2OhIE2+Y5hJcrHUOwFQpFwVKB3fZXBHsqoudq4VcN4Uy3ejIsiFK4CRkFQAdFvt
EnNECjnBQcpxYY/YqndGyGN5Ywc4cK8ykKK/DR/w2nYnbmZk7yk/XG1vR9QAQ6OKLGfTOyWr4mh8
zVam/uF2X7QOvBMruMAYSZYfHlrlWW4DbgBKC760XCL+6qI7nLoX3OiCEReTEJ7beOTlvZszGmhb
96QL5Ktit0wZpuCyTP97ogCw3e7y3XUK6mDA+F7vbXqbzqBMjOMj3OHHQiHgYeQMauGUy4RMEYtM
n/aAhNVrHO5X02obtX9fsxgZiFOD+5bheTDKkZfuUzVhcxrELvliCATuonqn3NhF/wSOe+ll9PCZ
Layw9mKMUcaeOc/XDbcIgB2C6rkuSjolwDYZW6DsH69Z/V5hs+YFKF6E3WnDumwlfABcQbEjk9Y2
7JUeaWgxv88Xq0uJvh84p08pG4s2WGuNpDMXkYO2duf/7/H6CCOF7uj+dCvIPQZwzHnzvzR2MIK1
TVE/HoLYecGFboDPcxa8IaJcosYg5rsrA4uCN/Wd9aUhsb0Di+997d6TI9DnZd2zUPRLv3meKfU/
NRtJoIMeoT399bW5t97LiXoQpC5XjYwjMGvCppl+uMeX0HGz8gJi+MV3VrRepetyx5wlb7+2K1zh
qKGkp+hUbjCpoZt8oW+GmOuNITWUwx5L5nvoEiCxxPmLKdZ6yTxCdRr3pNZ+4LEn8aoPOKWTlB9v
okclH75j8B/O0jSPYlXjBfOux4dpliI0KMAp2hiJltJpbvUb5G6v/H+KEPVHWeNk6lueI4fXc+SW
u131QarFEvZR9V1WMlCIFAbLwpcN7Mi08xM5GPKXfWsKu7L8l6fo8RJ2jBbDqfAe03vdKQe2Tpc/
O0sl/MY2bYxLcUSoLKpaXnfoIZrpn6n6zeKrIrBHFwn8vDpYC24EQW2TDPpNOq0tSdCU/b84DXFP
wVOjdYsDFciyfTc/Li38fS6ccavD0pkCYLctnYw1bAVLhQ0v7F4+HL+hbpS0MAmt1It8d5VfNEUb
79nHI6hoT3Oasn5Z/NaKLMgx1UMM5TCbMHVPe3Ra+WLqw1sV7EVb9oDf541BaM3DvFCJvtWgSCX7
ag8C9gDlQ6eL2MGfN/EURiv7oBJ4qbTv+Xep8QwrC4r2IyiGuDNg/lZH/pxqbmdYkmsfYGkN2jCt
YapSSXlv1VQb5AzDB9kB2Ym+ZvR3zSKaIKKfoDJDs1H8SUG1NuPPkv10alefYZ/TEWjHDjqydoYr
jbNjUACKqhLiFl0PD6vNk6mtPDX0XKMtDiQdElnqp+klX5PQNd9HNyAFD3sV95ny3q7GoNPJDfwk
qJl5E1fYRcQdau3e19cD3Q+Pt2tdPathC9UA2xWpy6iF5BxUcQcp7wl03zaIIocZDHbx2GiTiwXj
OfaLhqlIL7MWwpQPA6sBxtTftJ9ky/10MmHRAhG85Yw71DkNVrGAV3zhhV+qma5aUEmZaUoU7rCS
MtbyNFOs3wNHVjAaV6xYCCFHYb9gON86L5/4J4Aoxg2w+5vcpx+AfrQayjFIpQen3fd3IA5OmExS
xzac1R7UKa/oYdH/fQhIpeU1U0IlGI3PwDbmg3XMb1iK7ZtYerWobyx6fyR8JLkoJvP1Dgc/Ku/x
LTgL8B5CUKswJLk7XeA2bSetMfXimAxbwsxL/3KR5zmX+irtJfOe5b1kVzQQPOLsGStaWWtRX27Z
sLv+y9MJVQTUlXQ8Fpe8Ba7VlZqd/YHGThWPE47bNIYx/3VOI9FjYl8iE8bVL8chuXDydI5FjnTw
qqcAtPCtiQff8pPZZnMDLwiI4DsdWVjSfJ7XjsvBtnCpmWgBcawGr2m1fTa4QtRUbd4Ve/Nb71uM
7agh2u3gTBjh0fgmoEq5xI6NIqHOCX4camau6yciJjHZ0RowTqhEijw0u5HEK9NUB9IaY2E173gr
8jNTdgtV5wU3pRFPlcqnO61gttzcmpmgNNVisKVkwsV7NafJ8+Rlgex+ropknJFhOGdV/J1OwW48
5GIOKjGCa4TbQLgVvQGzNZh8ktavfLxAnC4YaM90FIpEF2iGuezI3NL74sO7Gl0Wwzl3WVvZql9r
1UukKMS0ngykgcIQTVSebCbiIB2KPopVIeIJeL8Govd0e+oMCL7MVkJxZ+Ojjx7Juo/tcG2Wk/0k
3AAY+SD12r2mhW93M2O3HhCwQDZx9i+xNxToN3En9IdS61N+UPkU2hQOohK97dJFmAii7WeRDlul
5H0I3OPQ4jZtPE3kZo89YUmYs+vHph//ubpb/g3r7JdiS3+H61U4KGJ3FoOSFx/y0dN8xZddPbeo
okwZJASWgMSRSGTyNfUv0Q85im+CYW9Ldi4yadTiiowi3AUBGSPB1ZrYFGYQwvcFCqJChYwRnMUq
9+GodCBGakPu6PDVWQ2fxVaLzBTZEoFCjBGQsyZ7J9tPzpUez6eL5SrDt75ckpJGBI1zsPfdi7CF
Tjc2Bzpe28I3vgFG1KqJGmzZASNJAmJyrzZ2cEZBRdDbJmK5ke+J1FTeE2q8u+PgqeASAyMtwAl3
sKTgtQqInQdSDl6TC3x2trB/ijSWKU8QqvIMjy0V+X9wr2nWJ5uMRKjg3fgfdnbNV0BQ/UBFiAbn
FfvBXYp7X6JLWrzZwqP2YIucIAkbWH32aE+Xe3+0luioQ73S+0Gm6NkjSTniRy8g0qOPzJWyKSVY
zRapp2xy2pRlcpCh1hIDFxPu5CCRRshVAQYnkBijtY+MZaZBeMgFRR/CnHv613JElIOEDuW8JnE5
5yKEuODnXdHo+A6YFV0YcGMrC1QUVWL5wzccVMjcG1gPcKWOd2UA4QwO7VWxRMkdB65Chz7b7TjH
2YY1639z0HxUK0dNe30kbv4/cfmtMRgYk3I68bw2q8LUAzyzxOMTCW/pQte4zFD8nzZrqoCHHf18
MULNP0X8lZf/oskuSAtRTCCcl7VmZpzP274f/PJWrpTTgS/o3WL4vNVLx88t/tu+o5ZrAeGTHcqM
ICnI2uou8gz0q6pH+D+DG0H3VwmcmZaNK5QvQnRpVHst7yrBYdsPQlToS3BUrhLiPHxUCiyQlXbz
xGIDjEXbwldDq4/TN4a2ZyN038ri/V06t6Z/Dxb56FPTTjKBjqzykqvb7v+K2bOxKLU/5pQTByON
uNRfkx2HqAq3i2XP4Rxsp1ygR/YhitLxpEAiBXpb6IgeQbtO6mPhG1iwrC2bdhVpN/plItrdV6At
fS002zs2Woo9BNGu809wrGL6A9VhFrH6P9L2Qqd4iOeKt3gwE/3/+rUA7zYWxd9TNlON9PfcMGHL
j1To4n/rr1b/f59Mrtj3C6t40N62+JMQ9ccFE4eOGSL/fl+YgUJaNcPeid/xWd3UKD0US5CKPd7o
fdrjsVkhUbVv3EkrlEwP+CTq2lgc2Ee5Ub76XozmKz9Dszga+Degbjp9yPf63OVD89N+P2S+QodX
dwSuytF4bD0CwAe/Pf0+BRiSALGfTF/0jDCROCarxyIkr6LxY6Zq1nRTy0g6GAz2H0ijTy/Du27l
D2KNAM5RrmTfkZx4VB/5XOYqa1qeQvQyCQuzB4eJdxTnoAqgvbemNsn/ABFveL6rw6tQ53RgWvDo
qbK+mznfrkWfDMgi6TxIdAShWrb1P6HoTbPPmvJFRyeWYPuDRT9HQ2G4WVMI3ZO42pDrjmx+TBfp
I6WYWN1aSMZ5MYPn5brHIZYR4IEnhslTMlNCe64Y3tJc8hIvwQkpCFnpg1lHiziOCwaPnD4wGFhL
9g1hvOs5p6Bpyg0MUvoGt6Y4YbJ3MrWX7aaHdnhBVwsLQZ6lRGYMlOgE5GOPXwSbD5+UG1L4wJ1+
Oj4AMXt2ZRpJt2JED2Kf4Ylcj4vuFYOFFqLkHH6kpNwXZZ6ps2qr/LGmkDZUi8DhXarP+r3IC+Q2
MmqqOd86ST+RNDdEkgq8/5LtYG4Y6rdPBtST0i4rVW6Z3SKuyTt6fX+/oSuKU+Hh2kzEP/VJ1JEW
CPzbrHtmTI2vs4xYH1UtGb3UudjdDUrDlEKahAg+ncurHAy319e8JtmlxMF6kIZiJOr+ehnzkpjp
bXExNzCo+E4HmFWKhsHHhhCbtNUu2ZiH6uVeQbYxvUN6xFWvv7q6KRuA0o4uVo5nGF5qCO/3yfWQ
2DtzPQrYwQ+Z4ImCNUpq8BKD8WReyqFM+0EUKbPsxxKC/8qIWE52mXFM0hzftYsAbnN5TccjmiYR
dTjcJIn9vW/gqew54DUy7p9PJvZ21/Gu5IgSOdX37fLTC/vlHi5SB9E2PVQPIlXJe5XTuuoE2Brq
q0swp6i3ub+3DBx3NK+D6/G5XVhQqOhT+GxzKait3ACF3xPc3NF9856/8+9129AhxkEUB0saTot5
bfwZP/vakr/qSu3Rfiv1pP0265cRc8qFyT2zsaqg3kCOuugtVtnWZX+CX2vtbNLCQtoJM3TjlVea
AR4Vmfl9gI0rjZBBWgdeWw2izGNYEkhVu2q/SHJpaJ6igqlrIjxO3e3MGM8UPGNsLWzAnUDFvN7X
mP6TopIo3lFgQmdR9mcrsLKRJ+9YpKAMhEyGIt9jelHnk1HqK3dptVft9Y94pikiA3vC8P03h6Hj
5mgPId1Hjo9VZP8eQcRGEIYVhg47SEv7AMyrvBxMyo8wT+ph8i4WGtFTAEP1lcyVcklwnm14md9i
NELekbcSDUooMT58ZoX4G5MM41om3vWHBu9qgM7Yc73miEGXorGLXl6KeKB4SJK/Bkyi8LJxirv8
orCLG/74x+YiREDXbIX9YYM0Hln4btIt5wE2H9iquIKQQnl672/eQQRLkKRdeBKxcQbd5jj+rbVp
pPZdsx632ERIVeeZJAhOvfLJS9dB7hRln1zKPQQsqxaH9mUywvGeuKwN5VbUmXHJPMpfsXwyPNbq
3ikxB0RQtnZ7FinMe79VXiDicxny3UxrCGrABAkqMnCfDcBaM8rKMrKgVBa+hOPAvBFIIgFM1Xbx
pRgUAbJJi8iRA7goMV5OOllymoOdNAHbQuqvfNLQlBfM5YGyo2+6dxjwZP/6mYsHliyY01ercey0
Gx4ujjpTVpVQWE27QUTyQ8KlS1nPWN+2dth2iilETX/QiET4sO1Yn//31B/xfFAxwvljfx+IS2mE
KbecaSJqNyQMsNqI7Y1GcdJyYNi3dGkRFDyfIpMDAlyeTKeuA7CxfsXNWUslPq57+k/VF1noPDVY
MkpWmqZZafifOldY3FUXM0Rx2vjfu92rC2SUA/cMN6SxmwDX3AoY7SKz7srbkuH19XT0+a25suEK
ryXX5qss9GLL49oX8iSIEH4KaCHhnXc3zhtizVq8unpS5oGM9mxZnKaAwjQ/Hr/ci3oUxmvH6TKr
xDz9rvNssA0HLLm0DqgouoEjXe3Er8gk+0I247yBI2nrQXpdxn4LOO7+z7X9O0SEF4Tdu7ewWbXJ
PDqFH3xuOgH3IWpute8LeY9oJpktQRmBVUgkWWRAWWlTvR4sB7Hoo6Dd0K6y5HtUwThO9tdCr15L
QDkSFP3b3d5V0owfyIz0q5vibFtQkxzSThqnCIZl+xvjUv6+H5fY5IhHd7BRB3oN+sdBPvJxxwl3
tplOkvC4ul3WuoIxlpYz9RxHXd4FiYKSVxlB+6ZC674oPbPlTok1A2c3DggHqWPMzSaPiy7bRH7f
dgn+ZdzYq+EkbMsnwNZV9SoQ3SQRqKRkfMO+K2KsaGYGzQlpehnr6ZyyrjPYORupMeX62xuEC+fG
nv08sPhmp25ybtrlz/snv6tJXO1Kbd04EDkHpNGXxMisbork5S+AlIGhLSkbKtgsyGjLMjHXY3+8
/f4X4+r9dUtvLo4Vt5/XbKejvFEPsMXc1/6L+dDkbTzDBMwFtGDqsOWScLcD/R0fhoD0KI7yhu/V
ptvrMeVmtq5R5ADjWJXL2uDVZUUDyEI+pRuTb3NsxM8moJEHfWdxbgE2DUsq8cJd/nQEUbDB/hZs
2+NmIVxhK29a7FvVegrJkT5fCoPTMMrA9yG8+WcCjkxyxnU+vZ7hJ061gk2h+vZfccGOSifmVJVH
sToaC/3znz6Tn/f5G8CA4XwghoUf1V8uuq2gV25NrS5qITfanT+nC62o96cscih1f1uzbHCyymBE
9pBUZFZCbxeVuvngWfNxRUGeRRfU8RY8ShnHDuO8HoBQGk4yidzwMP/DxKJrImtO3BIWMyK/6l0B
UenPmiM9Wn0UWJKRagOSX0GxWYDcDyool4OUfyXkutYQP7KTx8apW0DZEI5Pd4D8n0wm+zv6ybgT
/3/mEhQnTQDUGiw3mOMj4O/p4cWOwvVdyvfvrprauEk6O3jz7dSLoJA4f5Uu3qgr5FZKAKvT9OeS
2LsPvrpT0ppjlVPLOpMbiB8WdjXfzbxU6aNj2tLyrUVp1erD8S3w/AYM7mTEPrargAj8gwnvplIx
QkQczEFyA8tbFgJn4/GMNYtgpHWCvdVY6XZD/V37aNPkylyuJELZ/BpwXSbR/RJTFS7bNx5siT5t
wldgQlolzNDZ0Q4YIXN7AY8N6BZLhetzNCeiDGZUqVxl0mUYICkuxxITMR/05AYPLpE8QiDFpuHK
AaAkRq+skMmtgVLGGwyupu5hQXUTcAkRm+GfpAhF3o5nQaRFoPWeqvFUta4GS3Jv+XdSIrC7rF8V
sUassJWY8vbFgBYlap77jz0sWesdOAxpTvO5+Pu8HdNN7felPxnVe7+YS82AWiPlOp0iw7bWP27T
I6D7YUx+uDYyx3+qTz0E+T8WkOY8Nepo1FizDBdYdej+9ih2RszCAHGvvyPzVEUc0eSMps2F0fdl
PSf2vXXdKG7DDP6+cnCZZ9EMz60nxFWvEK6+bVSKw0sQKbuLgefRN4/U12THIZtIuWaVVYr0jQUB
/YoyZZg2gcEnDNjNeXCUcpQtu/aersXtZ+n3k0DrpEziW9RkrcZKx1lX6u+CB8t6+gPO7pLDJcLV
balQvYrXkXxXCJ2yNet3JaWZtkHPn8PkNh0d9iZYkG9Pnea5qJtT9+heaui8CKDxX41kGtpIRFRA
PsYpSHruGRRBcGiHGKrqzs/lBDoHDz129zCoRvwRpySio0TRasJCsYL7cA4imMcmZy2nI4p7abu/
dX/140i2HNcyIlwQjZ19+DnvDR8ExxMqzNQth7p3C6WrcZ+36lsuN8QP314ZLgzrI0W4XjLiLxT+
0nfjAoB7+nToUe77A0lqMcLr50y1Gnv4a0Hb6xLsE7Ryiy7RebIbNXSID48qa9CzmUkBsnASvLwF
5b/IM0aheUhgqxNxh4pzeuaCnyVY3hOyVX/ts6FURIIzk7xMg/yALExetMAA1F90K1YdTiQEQe76
CpXcbmF7vv9wlwFu/wTNqvGJJb5rafVIrlYMW/1B9+ZYUiCmHdI0Kn+2iDFxM38+bGG9YN07wbDf
4CouWdzCTKX2TeCT2naakbt5//AkgLOdhNbX8rSpwzl0qRtIVrKsopnSyqKGRdwpxX8Hhi0Yjx6v
ps/yPXgvjxE7Br5YLz0f3/zFyB14nF+aER61xlcdWzzdmircn/2Qj9kage6pB78GG1IM9NxUT4eW
gQzAYVnFwDx9q58mWnwqPs8rL3Bja+EEGnjutZhXo5qqHTGQCJTSBsU1AVYPn1cIgDCCrnOpJF7G
C6wh/gYknarfW80Hfhwt+fch9FJwgs5S+hX5jq77KGFxY16ze76afEWhEmtrsFfTw9vSSVeNcxGI
E2udoUpM6XblBik5YUyU39AAslIgHbwJKD+mXwDMZHXb3JDsH466h9sR2zij4Z3JcaE0hWrH1BEU
A4V8gpbeVXOZn6j1DbY2IsQi88eTxbCk/s7mLmcwrk63p6ocv2j7heQTW5SzPgPi/+LTBMn5M8Eg
INqRW0qBG8aBD2qRLfarJcSLZGLkCugYqCDZj9fvkODrhODzaadpS5jJK+dc+B951Pch4W9zC29W
j4MKre6GQFTHKj42G6gmlDriHUYCKp0b13Rfm4bqF1yq9JYw9UyfnbNYMLVf99PnPAkgeLTEuUe/
1v5v35jHch/DmKe5hW0hJZR0x3fQbJJvWFUpTIzojuhlcZFdT1rU+xRqFuhywAQLn+7Mia8FO4Xp
GpaBgP032myfNgNBl3WtuXpe9EiYr+vnwWfzCxOn0IWUiaYL4JIQhs7WrSWmaa0Fwoo23Q03wzC0
V/CgigTvalZDVEZ2NhtsT976OJ2P9sFy4RUeekaPqm3gfWNFzXiQlAjieodrPJZ1+NTKOoabqUnf
t0qFkFAH8cCs3mLJZFmoro17b45kmWSnVteTsk04Ebj/Cgjd5R1m+aFvYPwsMFQwEkdmCthn1CL7
0qLsIflGTMt7PR7xUXUuAIiTXedLx3ocxS5kwr/Fpf4/Ti/DPM0o+2cvvplKlc0WYZUtH4mFbW4j
3fgZLGnEjWWzKzTb1mTVZpiJzo+cDwbTH5TKpZPq2qTj8eTpM5Ba3jw5Pd0QDRULfWpAuMdzbTwM
MYkL6ry5fON9e1rKJhUDUkx5YxBbOY2EiycGJs0y0bi6SuwnkXdP/k3Ov77I9XpnK4L/worwvQRP
L8saUTVbIETQwRyXoCLbP2hJ+MqjYdWrk5mmiKFj4I7b2nlrvRKasas2tAwyq1+cLO03yzvVFx02
LvqFCSbGJRHpjm1B6e356dVPKOaqjv/pIGmNideHXlcAvTm+xfhTQVgSWuuiaa6e4ROkfz88py9O
PftcUCxLSQvGA7ZIraKx4SkmkZopuFm3eksvKTKp3wq0l6ECLcaaeFoKRFr6Tk1WBFlxRA1LyVyt
s8HbsZ0x6yarTm+kIt0GOnsqWRKw3Fgk0Z/GDKGQAjkraScFzwqWDGjajEBKQbeeJyr3F4oJUFUl
lkpyOZqe6swCYMKTSuh06qGAiZpVGkcbNL5pUe31AIOl/fPBANjX02tRifkx7h00bSHTgeRJ3/1B
kMfwA5lw9nFj9RplSY8oqB7XeiLSSs9xCz2qfoNnLAP08lSrH077Xc3wWPgY8gDq0O/3Ahc5MA3y
j7s8feEO+SXVZEEEB3KoKSS7FFXsR4P8OjFUIwS6PSFnKhHVnk5u/leZrNFtBmlxGxvtMlanvv+n
ivK00hpgtOLHQI/1Fe5U1tTtFttZ8898RBBF58O/q4gP/H7/3kziMKl8uRNEnOOeBfkaEj+XhKTd
7OFiX1XwW3go6tFro3DI7V2MkmRtsQvKEMgygG3hKxJfW0jsHiy0JESHTIRBuuseWWd402wgm+ib
jsjfWuyS0Q8jGzGUMakhxeCuftNnnM6VA0zclsP8VAFy5Fru6mpxJj70+m/nRU9g/f6FQxJpquzR
X+XRJro0BjF9wRqHH5Uo0A79QZSxtl+5G1WgMqSj5L92OSFq9RyhubxYazxWoSLe6wiigHXEPCDD
DgIED/nWxWR85a/u4lTtxmtqKkuNEnTi482Ji6Bk1o1kfCr95AzCub783knmdRUAtwzPoa4yYX4Y
Z1u0qsH1Dv3lTZiXxbF1dgyZMfTSjVeeO2WxmityV3qOSg3XeZOB/iGNYYHpyLUl+WzJJefUFkT2
WL1sqW+3n0Ip5NUNHzNBzqMe0L3dnGPNj0QK0+FoxFRzwltl8zuTiPyVWnLwvfLyat3V2/khRT4q
ccqONb23bh6uqOMNt/gDe16fMsaVtq1zHNmDh73JHyWLNMVYll9LQyjvzi00+NCtp8JJIDm7B4J2
U2oadhbVSN5ixsA2latl8+DxeigXCtJNnlQeN+V+lWrhTCZxbdHCG5817YQLQdvrP2bB4Zcj40VT
QIrGydhTL95veuQv4LuNXpFGClZe6LHQ1WxOgpyBjkUO5Aq1thGfMyvNgKFaEg8p0NkzpKgn2V36
d0/YcoFfh01ttFvSb5jp6hE+A2VWejKN4oGQg7xMDFAp9qsPyoT6DamegGxGsyak3oG2UXu2pxoW
0cOAU9q+T+ZX/PjTeg9/UMVkkN4Q3KEA+FB5EYu8wMj8pkx6SBc/GY26s0Ks2+pE9I1UB0VKvrLr
C2qC/2pTWT6S4VSE1K/XYjIVeR2RBiVALjRTcnBVq7axVvi4IKI/HzfGwhLLE6NbcTQwY9FunoD9
dYaCQeAYeCyzd2lsEUScQ9wtZS+KsvQRjAFLRa0rpu01Afz8Ec5rVMSHip8boda4WR3/nyzz0Qkp
sAaXNRTnw6ZdCSys5sbD+uNqW175VE3JszYuD3E6LuamDBgjNhee3NMvby0bZkxSK/48STWf1vth
vbY9o3oltHl9UqneDuRTrg1zha+rwkcUBit7np2MwmPySg/iv+w3cIO/dBo49eqpcm3MKqtJcn+A
S2eqJUSwWQ452p/pPturcFjh0go3HQiVwAcqrfT56q9aeelp+MKY/RJWua11IaNBuxnysJmFnH/T
3MbGJwAqhtDZMv5cBCRagqCbXCxm2jX4fn1IE9yqqjoqaQ2lrdNNvInOEfOvs3xcKAlc6fAndot8
SzUx2Ej/RRTig1Pj/JSc7jYYyIfbU6CeNdv3pUuBo/zL4dj9iy3mb166nelTfQ2B45kjBb9jbZkV
iojClYG7+dhlG8q9A4JM9vm/hgVDcbCBWTVaa8DlOXINVAMhXKlJvX5+s1QzQzkKJSjmyJoaO3EM
ldA/EJe6n/ITnnQSQsIL+pF6SqjXYhC9mQnh2uL4s8GG/h60OSr9ym/TMLHH9uzlCjgNUByzQzgS
XjorshjiJnXH9gr6v8CPaKx2HX02bi1wOjydTOGW66KTEbh7fma/0BWoeKW7LRafuWr06X3EIF8M
/SJlE/wO/QlXvNw7NtQoA44Nk2uJs7uqeY90MDjINo8/bET9tC806rngEukucRYxaq2PlTKST04k
oB5Y0CFF+JfKmmfb7ZRl2fQTPIMKf4aMuKLEfMIeg8Jq60Z2MlEMgzDHOr8MbBeF1jyso9y6M/gW
grrpAdGRGMtCgl8ub2rJLrC4Ptyw8LZwmyyCwAwbC6gwyA35BYsQk1ZM3R7RNt1KlhGDQg7ejOEG
rrEWCRpsccSzz+bP6l16ca/mQfnLcWo5ruBudblB6Sd8weBI3qg0WHR3bucl5t5err5sGC0A5+ew
5R/kuY8viwOEcw+AOJH1FsaBGR+wUzxpGAqtTxB0aImhFcrPnqDk5xCAlyifYuTcXxuBsIyWLdo0
n+larl4GCrHfSWZeqeDLVtyist3TopuM5g32ikzD+Nu5YCB3kEKsPG58/fSRNs1q3ScnsnPpSsHH
ABqHD5ZeZyBfoCjVJo6onvNXeZRYQQugU+HxNKSMYvJv6v0j97BzFipF5NienIU+EYDPqMFxB6aT
O8pSpwRyCGQy/H7GWtWudUTVYsyD1Vy8EinXprvESEDkk6OiUg/7ReadJFe0vL9pjt05pHqcqJkt
8aGAtoxgNeZ9aBuMuntPHf9qm6EWaC2sPPGQ8832x9QPS8D8fik9CSbsOYTVE6pjPhVhfvf69bn+
lpkhlo+dXGdeoSTjBL7Tcw9BjDMYyfvP5YPRmy58uQjABNvnBzQL5bo/lcc7xBZrLb4fgIZ6Cjcw
k6HzBzaNjLNwYybeRuyFZgK1ZZdvHKniJEwkZSM2NzLxlB5Ug6jpbDoKIEKv22DMLON4qf/tAufj
1FauBxvEzXwcZKqNcz2P2pLYMACNSwiHL3dGvkftZrKyIFQsGNwNY8k3tqGekFus/d6DutPBDrO3
rPtgzsn3B3IH3uZ3m6Sv1pTpWITyJ9eG1oVFIegttJEZlr09GAiTLYaRD1AXeWLMto6b38J0eyKU
orWwZgwLF8jebZiCZFQejh4CZ2X7ewMvKhxSiW+CP6B3XEGx78z++/4Pce56HZYcM6ipBw0oGVKZ
0jRSk4v6OS6uyQuEdbIO3hV3GvkvMhr9Oez1QqXNrD+AilUQz4gTXOUmRx8EZ1AWYbEUCJabAE6Q
yGxuPLL5txOOH/v/i4eiNYkC1DqIIu9HEZdyOtbkdVbf22cGVxttQh/jAkNbDh0RnMkIL3/SCcSE
qlAXYCf+J8pJubkVl83YsY1cYh6h/KQFckYdJVdTnWrZHGR51tUW/K60LjEhnMOKBRY6/Qd6A3l6
D0IQSA0XtXVXBKHC866UiPX65sth0piHf5cLdvl9ZlN9JbHoBw7kAFRxcC+2r2zsWe+fwf9RdjXH
ArlWaFCO5gxAV4Y8BMdqv5+gtuYVawCg371wtf07OfIsvdV/yurOL1fjQhHgChSQ+rhCPiXH9JyL
d0Y095zm99iES6OJsSQIjbYsy62PMyjPha8jEDNlfTVhGIj1ER9KZaIF9KA0Qf9hzWhWi4DYxo2n
qQrjTHUYQ/XlAGMXdxW1yfdB4Mj2obcw8HBIcj93JRwh3U3ANLgQfk/5zSrFy6rxS2exw8uGcT0Y
z8qcqc3+v8F2XrFh7RIayQ4somlJHvuUaSsKc8WK1uPkPSnp/9Ytv7OCwxduJl1flLjyy6dBrX2P
angd8PrOTs/VDKJH1UGWfR2o+XW5anl7fHvO0zCNoNk9rKj0VlBfhe6aVEukezttKf4BKTE2CGZ3
MZutzeO7hyqrO+SRXrQMRPDSn3qs+7Kq49E2w7NTZESHCmQ2VstraErFGUWcUDQXTsPgsRKJ336R
fXbMOBDUkje+CRyL13NgZWeI61bKLhP7dh+HHL0My+btZFVR0azapPgHgfSQ+PLQPDOj+d0ZDDx6
SO5+rgB/dDk0r1Q3cUSaNOW72YHCUnnUJjBJxTEEKlf7rKC6m8691pOKintE+H2k4RjHisMA+SW1
aSnEQaGmdsm1D4lvX7GYNDZCUQ9jx/jKWeYDAYjr9v9amnMp9qPxrC4xeV7HlFOpnN5l5RCdE1n8
cwK5yOIl8D7pnofXsQRhARz1QvviwDtQ0FfhyPI5nVVSsW/J0rqCP3K234jLmIqB9lapE66MvLwa
A2Lx+Yv5WTPxfgbWKVkbclN8v7xXqyIVpFXbZRr6gLuYMWctgZ7qIbRaNwi2t889BOGvM0M9Wlov
1s199xT+/qeEKsnYkPIhyOIsvKgPhtJ/JRDDkV5p9bTv0T14Xw4iEyADKptBrTmldx3ptXLadJt1
UzZaxqUouHPqxqRFFGxFtI5EMqOb3hrEL+ngG60FDIlR4wiHwDgYdNz10aQSj0FuRHN54xqy4t09
4i+d1JUudAfcbJ+H+z9QL6SB2t2TR2q8nnot01PitAXKcRrje1iDKuMtHnPsqZLN3MLPIyezzB4K
pEl8CcCgNEDZsTMpCFQOYjz5aUGwjTCmBo85LBsvwjQCwRRY131lYBdRVLrlfJQ0S49rRMyXXoy0
gJU+A1FA2rIEvlVderiWdz0kc5HyaOo4rDRak5EJjLaUF8Lsfs1QQCSbdmf07Zm0YU3HhGN6E8Z3
xlvEHWUvINQPjaiAxni+iUaF1qP4/h/PCuTI8H92tIXkEAeVmb8p9kAQq8TI+cIrYPBA60iaO/dP
6qdrLESCmi/t79ZtBKfPUEHO2o0FTNgzQZcqfnduxFepOPxeKzSiI557PdYNKa7kLHBq9yDPRYgr
MqjCa+CWMKj1yJKwQH737wl7g7bbB8vzoN5aj25gGylUXTzoNCbHinn2Fm+wRRWZU1XYoK6xrZWb
2oKHLLquVzeuz8/BmdJo82pdwvz1PQThC5xwp9nXn4+9Gr5bTqgeR3m0OK8n1jagRFDgLLdag6d2
T084jl5DXjcB/mX28sQS8GF3GV8PlaN/WdUEvuEpDclYS7GJDkdVGASmbgRQJpmO9hhmQsFBJTSu
PbkB/QvKNMIeAaSFQTI6wJGZgsAAfZHJ1P4xaJrxsEs6GcFGBMMsHLJTjuVRpb4l+Gwcl/j/o6Bf
1d9x5EXBociDrl0tW4RgtwMqP8qGZ32b9tdXKoVTLKAbEzzRMbrR6ej7+ntyzad7enWLzlqUwYVQ
aKuNI5ixfGCiDmOE8sKMhO44Fus5AJ8TuUxGAW+GF6lt+6xY6Gc5uOhrXaf0RRCsYfnA9XACLcx5
VihLBDSJYQa0srjeSg9703ta9IaaH5GPFhpz+7h07h42PldBhagNcEi1HA0jN3ngddzT4mXLLnJ4
EyZoQCHZOMFZyVhr4RSSe0QRZG3tQ+xvfz/y9olYDtYNERxbCK7foB/uw47QAcgJsYqsueeuLLmD
YK58aBxjGxizcUqcFGnk+sVo/NYq2/ZZCRRVEofje5p4M8qFSYG7IlwHAyvjPWzN6lvngV5Y5RGh
NU9fmVtlYmqjKpX40aN5Y8h82Y+vWDrPI84M7TIUCxolZ0LVa8xhmJoJZOCWWZIBAToMUft9CY4n
XqWF/k71ADNQddG5A8T/OCgHiFkn3sYN+Y9R9iFYTohUh5Yt3pgIQq3hQ5P/JTqb0D9dnQNQZG1v
szQmUxJJdc2E+zL/qB2+8x7l/BSBmylurZ04lSSqfZG+xx6e8pS1KPV/rn3X2Ss+gi0015sVXVn7
q0sAScLDYTd2amq39L1STm6gf9SLqd26r/2xjykBnZqASTGEu7fgr0et11DRpOrmWcWcAdJUa7O9
mSwWASZ2lcbi/a1HOa4rcl4u6W7+5tWUDlzusgr33NN9AcMXTss29GR1S5SQNTp7ydqK0bK1bv5s
W1u98HH73IEcGnVmGDHlEYBGxRXzqLGSov4u5OVFTQ6EI6loWIYif1lmh052BNaViBrhkC+GqUuZ
xrFxi4OE3XFcnsN08QLNO74ViXimaBq2GC1Ku4DO1SeaZiRoVDTRCKrqlAvTUO8PT6yZ1W1sKGdM
Lxs7ZM1K3WNnVgjOuN9N5n/Ut1rSVsTIqIQmcJ521DEGsPssIyKmM4Kzu6jRwm1OQYo6T1Zen/xD
GVx86ujuKYMeg0/WViK2/JZQmh0yebf1xBVGuE434uGctHBU2RrCMSE8wDwrnt8u6+ibu5JcKGdN
5dlx/OQi7vNX7WfK4nR/UbW4QqUslL+R3cU35CdNZVsad99x1FWjVoH94NUGR59wsnnWM9TgJM/4
QEVkqQm002aMeW6nRx3fx9FfafGz+pK1Hvl/LbZwtPBgoMi/d63cBvIO6XHOfdnxjUdzejD13Tax
siOE5/0mb/uVz2hDCH5s947lPNH+9aJtLoWSQKKFO0Z21r+rL+ffdYB0IfWXPZ0VvJlkRc5oa4Wq
CYa8HgQki7ChAGA0wkVsOhJPUnKWnYCgxMxK217sKs3d+Dazx0+X/EZiNqgTIxUDA1tQSJp4mNoe
FdZYB83agFbGw1pZiR4SpWu/Uo0KweuFTwgRAV4F9hPYt0iI+iRKWyseAeMFAR6owAIk+LqmiMcx
yglhpShG90wulsvRAKFKzWTasZGwUGGqG7abEBI3pkjvMtsXTPH5AHsC8ioJ8W1lRCDUjcAyAdfK
T0vCaa+fq47lX3kks8FUuVXYI/oyH6M78TC+k/OhWqN6uGHvrbVdjAXiriHqkWdrUtxZLXJu0SAo
MBcniKoUrArrj6nXzVDuup+Vcptj8BuOfeK/NVCGKmjCCedciWQyibNlPHNe4W1pVrcIUtvETEsB
L6c9wPtnrCUJ7BPzkAlsPKomnlxliynw9Llp4lxkD8SiErnOOiCAAdJM0BILZBzlA9Y3f+ftKBwX
Hk+bs6686onF/dp9GMWXRDjtRsGIiftKeGkTtiZuXwg/0tcDm9+chE9P/r/52KPmFbgKwfERMJrK
4pu00FQz4O02SUcraNH9KTdGi8agP/CnszqX/wQdgUeyfWVXqFj8dHgZB/8j8a+J+6w/X/g20xgP
x6KW9ef3TMxnUg85ZQFgVO/puc2Fkp72Gx2NZcL7nq5Drxn2X2otY6vQZpyGD9xfRyEtKNWyIi2o
3kLQPj4cz9khaC++FSzQ4CarPqvyq3TOum+WEMOfRx7awUN/yB9Y2QKywTLwkYl2drefUhMKHUFf
oL18VVliBAjGnJ13Z1wPxDanQUX+IdMWX0UYza0tkMXxt170jBx2ywZrmZsd1pRak8KNlAg9ZEPl
Inshyk6XyJTvofQhdUYNILDSnxD8Q8CcQkNA3XTqYIHsil5J41eVL6ni6RSbFO0KF4zIGaTlJMtS
oYTLWYimWjwTtbSqknAUoI9xcgsFwmrf7Sa/3ce1Amp+wbuB+H0idjSNSsZf8Xrni6bg346UdOXR
LlixV/VMLiSnxLuRPF/iRz8ZUn3KgV9+khyXcV3T/8i4UiEvMmHyqaZpC2K/0MpDd97I7RHyUJq8
JbMvl+EXaKeJtb4EOrFBPt9ulRY9sck96E/B+VsSw5cSWTNnd/lqJi2KBRzHBnjWk8FYlzzMvCBg
Le2OsREXaJFffsy97PllygKkrZd7/brVyTX8muntr34F5p02pUWrZnPT00nYXvxBqX8fZzNrCckm
0XFl7TKW76oCPlRlmoNJEiWBDhcebxh4UG9Ynr5/kTQ90Atmjfq3rp6QupRl8MLtouB/zyO1WHX4
l65BjfnDV23QhwY4gTm8F3aFlA0Zg17Qhlh8BziXv3OsFFu84TbRKwNA3yOeDbhNi1jbZEF7OXtn
62pB1crbOZ1wvdytzA8bVLWT6l5sG5lEUG0jUhnyRAp08lxR4zhyfC1BnDqfbckdj54kIu9ySXrN
LOsf5c2UeSY5aB/XMdW3JHWrBzn70It8M8pT3If3+Or2PbhipwFhJPS5MCNGFYkxqoEpdXHa1wIq
xdDoFcO8D1bfzp9pRJr0at09UCi0ltPAbhzVHAEjxBfrAffX6KKNpdMgQJBffHb7HWYoFbIXsmEF
8zW+niJVCEggrFufyytrXZY2h3SXiPC3uzGhFf+d5MdFacJhz1Ad+J7GxjzIv3/qRKz6m7CHHKyU
8htfJm2XpYh33e4a13RGCnW6Sgrk9Qftp/oVzn7PZSWMYx5BcNU3fuPtOYnbFgBG1tofu4Cmu/oP
zIhZ/7NFuL5AgVCiEhCmD3nbGrqRMrhMeQIFy12CkOHdFcnp6yxq8cdI1NXHnw3OGIeqXKJcXShs
ehLlbvusbTMnARbEj2hR4mgsd5saumnfTLQgkfU5EyZEKucEDeAY0eSZ9tPjwtDkv8YYETk2wSo0
2KSy4WNPnfQpw6ehRnJbqiMSjlkgq1xCKsgYkffLflmqyGZFGHx9ENICl0PdnhoLmMTMfEGcJwXh
rZivIPUPYsnAbZVAm9KK3/veUREq4UpXfoiNiEqrtlOPNlt62T7P2WFLout1MNnyqzzrVknFqpIC
v9rrxXTrfsLg6PuiyqoJMmNuvHGk2vDxJsraKXjW+7ub55a+tCu84k/FGFy72NlLYQRLldGVqSes
+6x3iw17kIRZZ2ViicFgEbOINYBDRkqSbui3/XSaW0I9QgltDVOpl9Eq0VvlyiJNu661iRcy5SWo
lD746Ne/tjU30pumG/K67HqI3/No+oUL+SibRUhxLKYiDtIKU1TLV/H5z/mqZiMc36IjnTvHhQNP
DFyn2KRngPMximX0ZzQIquUSfvRuwwgG3QQpr2OhqD10HkF4U1G0+kZfjkctbIywMH7X4r2AtZYO
bnvzX+AcfJv7Io4pb0Oc+HkW2cIcdvdmiA0RgxsU0zxllR6M/KwmSkXG5lsaCVAv8t1rmIY4se0z
NwgPPUgGrTAXm4UhNjj/xCtU/AHOpE7uWJETnswv95Pla5EV5BEBlnItGbeck5oAfKJis0GCD8Jm
ROfDcvx8esMcidlXdHELdoww/aTh3J/j2o3mHiRZPp45xEMWzFfz2WNC+S5MIeLDd78PCOhlKORW
1t5dzRQvXCY/kQVhrkaIQKs116eygkitYB1qBM/TQEi0LEaypcb/z6YDuyUlNBloF92No2jhkrHt
7W++ZHyXvMNsHODvULQO5xWZ2yP77lbs3G41A5S1gSsAGhkgt+8M9lYVZL/Po0xo/nTdKlz73/Qf
YowrPVfNOfdft09/eyM/znsQWMDxPCkKOqlloIm62OE7CURQiRQW116oabv5hjibt3Wk7cqTD0Ct
8JKLDC4oeGvYoX7cL2bSH/5xeuSCH5xKceTDZkKOsZU+PAPPNYqKll8VJftDLQtLrHW5UNPryfyx
IwDOs9rboZoSAu3btiF1ZEZzplPJ5ROuq31XsGOew1MT4MDunl0IY0j33Cts3yhFZ2qwnEU+NiX2
GnSIPQQjkUYDj2yJkgp5OzmNOV8QsDGczPI7kLC/fYmeLQWK4viS36f7nQCtBoQdkZCUg/sGCiiz
00XUwgIqft7JzxMc0OmlydHWERUh0ggdwohkNIInU5/8pCyq3i+AIqA6G9mu8ZLaC8Npve9KMdIV
0gB1VBBh+9aEo3a/Pr5h3/a8HK5uMZPQ7HQbOPSCXwdtEJ5jaHniFao2HoSEUAizBKgjgFv5C7m4
FQ8CrDrzpZhvzCmTvmEYMczf+IAQ8WMrOERrSnYNSG/ZTApKxaVjuuoKzGPXpkZAfxpsCpL3GfQw
8aSPsaXzES5NoLNMKI/y7hgYuoHqYb8FwM/zNn4Uxh5YB+UEFA20Pp5EE7OiOiRlLwwF3MckNIHI
qdZoymlb4eW4ZiFa55Vwm/2Air5GuGkfS7KWulA8mgKO8QPFjz+8p90QgXiSj6vxhDQOv5Eej5tr
BANFi8BqgH3SycWSdZsj0ytBHU/tNmtluhmQH67esz7PFLaDfTwgFIdwwqjnBOrwUkLnZrYoO3fB
V3feKuGuN1ThFvj4r8S+gflEPkV0+un7o1WzJnQ8Rvh1GXaxRvknODCDuqnLT63fYFoErFphLAKI
ok79QAhRFu0HRIqHxQW25d28G9qxmYeW+ZxxOanGHJbUdziTPLt5xTyqeOxV4YlLhMJAR9YsBzvD
IxOE7HqfW2q4LIjri72hUw5xc6gNIsdhg468H9/VlrsOV9g5H1PFuK7Ifqw6A3EMvUBqQKgwP47u
rFdeQ/P1A6dQzebILnOqKDlNbEet05st7hFfyZcj1H0zb8thoElLU99csz3SWUZq48LK9GTw4DF2
iQPtxGKNj0BvFTLC0I2puq7rzGIYmPaUz50fsN+5UXEtSL1Y5HVkMACcnbxSTLFuNqZyeeUocymn
tJaK2eYXte1eh3ilscR1jBv9MZbwN45X/hTihh1kIxMMETFV8XK4oMLD5wsaHj9EexyHyTOIbWm2
E+bkBICuG5G2dW5yIPQHORhDArCiTfV6VVRsV6w40TqErfQtb67RBggA1zRksnT42LJeIb3Y5QCp
aWXrvnyacMnJh0TxoM5PebZ2SFVY7b1h/5UC41ut0YPpMrXP4s9664vS5TaTQErazQVqrqK6yuAx
6uzIgJhh01TFPfui21La2nG77v61e5tJX+3sWjgscXOVKafgZxYjGh8amvOGFWTRJPnqU6y1OHny
MUjd2uD3pvqiMJT6OqrFvZlR+fGY873AUqYDVxoBJn9zM1OC7XYQiIayRnOH9kghzVYBzarkzZZB
WkYtF87jjy8FvKdwbwaK16hpcH1ufSOCu3MNM/iOKUL1YvDG3XpJFlRfXY/NXmwoUQN3XKjNu3Pk
LqG0Ax5oT4j/yivAEndNzk4s4VSnMG1HPMr5tTkFyZGbgjg1aQ3VO0v8PFw05YSAO2hXZJz6ouv3
160HX2tmkjiPD/ichZ+tjVzTyaUvdumlQHLlqVHLE/B+C1S2t3Xi54Fny+lDrDclnAOyXuh6xkCD
KYjIwuNcA5PnnlglMy1/2ISDPzt0R0S8RRXRKtuQjIkigapU6Iiyw0IVMxfr5YyMKuxki+CMwPMX
UFW5Gdacm+snKcoE3DfJLLs4KkKn1660/bJHHn81Vn00xcqLujPvilCLikG2qpejRdT6iiCYhdFG
jJd4KfIWhlXjpI/xgLN38AyOArXt5bkvsjz/DmX3MJbCMqapp/9BxPpM35puHMFJvGZfmFN8KbL+
NbT+mgynzOhVEbcCt1gOgAIWKYooUaqLg4LoIyfMYVv90gd1sopp4jY2Lcq8aFC6Qd+8mFvmwmSb
+2MtdBW44T3fKqNPFT+7bJZ1LxpYNMTzJfSiXo6C3ADcWSe0/MJoVBjaXyY2UB3fg2xSsaBuQ9ZG
Rf6R003rBm3luV/rU+BFeH6zs15d0bmkFTaLjDFBW9x4qL/2Zva43eoCf/1+BNHn5fnNGqN6X2qw
vaxRC5NUeiLGA7SFEi82VqgAHNvSmHrObjhMN0bH+EywiwfaWGQuBqnmyofYgpFYX8/jKZvzT2QH
vynzj9c2DfEQieHtWrrvcygusLqHroZKiamCoxJ10D3W5C4E6+IDgTXelGFS5WcTHGj+rP+kvg3s
c4NugjzVITpuQQAqPo+RSZ5hN/2F2I1CrCxLMqTY4nxe1o3d5umVgO0/uEJ6sOxTb2nPVazK3Xty
Nn8ivBnYHSKxChiYcrsd8yvcza1C+Y9/8yvdFShDiGMk0y1TMTtI3vAvifgnAiNBSG7aBm/QpvhC
rq8d5IG572K64jINlrcYasvLUTJ5R4yqVEo4gpk5f1R9PhYcLqfwEfKrd9oZs7XzUZg+UP4+0dsI
HMNoPhtN+SoBvebPtLI0WO0wx2CNYTk2MZLmWG4gn5A2LF0/y67ePPG+fcB+FngyF6Br/6SVi1Zh
o/jpB6A4iMLkA90PuyHieH7nTUaM8Jx+c4hBFkDx8dF4LCu5sXFScf2GjTOx8uVgq88LhyJuEsPT
muQ+BiBHDbbvbquCNjWgzai0OB+cngAWF6G40o0aIyP6MAX1ylwmffv14m9FCnokXqp0FEouzlSr
9o+O2uypihZ8Wh1v3FDsK6IMtpAl1Cfoenkv6lTDjfPHtfESSlvhY5Mxh2JK2hEqRl14iLBVPXzQ
yLZAnrGpxL4aAjhIwHZ4/JJLbxUGgsZtk1x4ICEbo8lo5ySPAg0XbZLbkDQdk9cLf78Y+Sy6SHh5
lyeBeMH0nw/P9v1yzEfX17OvVw1hkwLsm+ASM+ECzTWv/rjZUVS+XGTbl9EX0iWYp9xZlUg+XWAe
T8BZbO8avR5PKR3EACy4zZcmYeWJALvQr33ZaEcOlDU786sF405g0bEm96gYaecfv9EjNZAPgUfu
JokvnIxbDWckrobVIJ3FjRrMBVYgKipOY8/nCHIg6YdL5kPytK9YKfy4oePq5fDSz3Zg9sTfV5Ku
F0G6Ub+4E1VgpfegSEsM4tRsxMuAXqW1OKKJocXrVlcx5YAajXRdIxQ/DnbZaiEbzd/PA9c1gPSf
W6kq+2p3pmXE+X7mi2Lrz+/RL7Vb9u4HS6/hDgFVCKizO7387QMW/U9y92pBixNOexCdme7DFcq9
k3HiAkd3cssIRW5p4emPcoWjnTiQ3lpysLDLZhNyqQwgO8BYC3pEqj1N98uh4bMw6fasstahzOWa
DYCvFzhM+C9JS5Os7Ip8iy0Ii5UxjJnRjadaBmf4F3wy3Op5euO7v7aM0SZgYBh1cg+D4D/UK7M+
8GkCzYFrT7gdjox2Gnw5xykB+/Ny8wDi10x5Ra2rNf67H0LOKOCBMDJcmK+/F82BxmjV1lISZV3v
kZ/EvCNZoH9KM0vLriXChDXDoNryWv3Xd1FKxXFyorRh0ua0vtkOzfplYCZebJ3Q4JuesZsGksGW
5Z6gpotcagF16uuTFp5lUVUn9z/ozYlH7Kz5PLkPOpUIZjr7zukRnWlvFiSTaWvskPadCyq2rBU2
RiI+s7/pKlTQqUM5psVUZAl2V2nTLZz8yyEpbnAwCSvPoqkVMMvAO5lDNEb3gdwTlahkUFQmWwv8
6PVJ3Mq9szjPM9xxQ+Fvufg2tPmBgPvUYaiNWUw2cEpMp+KYvHgLuVFrMileDULferBl3N58vNhH
ixleBRcD0Dwm2XfAjGUXCXuKUkosFhT01x9AyuGnN/b83Rble/GSms2tWOI0E4mR7mdM2nP9tSEE
X6GapgkzKE+oUDEKAvzuu3P+uwioUnYFQfk/fwcA9cPgPmi3KEzGcBZvzDLTwAbXVsTDntRhWJ6+
BXPv7xyF8MfrekgN0fXOqEemkV0EIQ+kyAEWDqtQX0ffPPhAFxiDvEfxluy+iyxxmZJ2yEcMTVGe
bEqh761QydYzkAe1brfvcAGm6xIEJ2zwoosVcWuxAaIVgxzFIIoMxP3R0sdIeHbti9KFC9md5rs/
gAdoQpDCv/adPC8MHth1lmywRBP7LMX53R5AeimpidoZSAwA1qfdFF0ACy8WHVY8kVH8ygoeYIuh
MdisL7WxACA0p28RT4CZU3OE86qZP3KgsxubMT1LGo/dr+fCV82B8qSRV3QfbKkeR2IT4QD0XEUl
M5+Y3HBA8+dIZNcog3fmJOTskf8kZYOqRwRW3mj68omCPV94A8CyDgf1WHXzF6cpSFE9r/6jZKmo
gDLs91ozgZ9kWC/gCJyqf14vjnLkDOb24XuQNJ/YI0Hr4vgHOi9LOww1IajCbobCW69TREjDyDvI
M6P4B+3iJ3HHIW/Nxd22RL2/gEXONegkRgwqy5ES8JG78sgoyS5FFogWwjfPrlQr+uqmhpDi8HAQ
+JpFAtaCJ72mCgf6EGewYQQlwCaoiCsYdym9Qpwau8z+mkC/C9cUsXxwGl7dNqK9nzN1Er+0AMkz
I/Yj1/Nu9F1Jwvt9qMaPmqhjaXYxJpXHMA6H9R9bZe/QlHhYbHpwjnGkGiBIlf4+J0C8a2Td48p/
W82gnnBwopst0LrUT2wQ4KCrjqEFiA/BPWrMpTCBM+jDaytyrdzKCB0zDE/OcGjfGkKEVATgHMC2
BYM35fSnaaf5LOVyQVeb6UH1ZrnyVYYeb341lAzbjBXv1M5OkOa1hgTishEJTB2qdQ3uAILjP0FQ
jPOc52JyXvvyfrIQX67YNPG2C/xapvevQyBD6cAQEyTr820YRRO1Knb7PaVXJ/qYbQqDPTSDUSeG
RspGFpHp/Fo49QqVj1F79BEZabyNh7DLk/7BhzjXMEN6weIoxjrFUCTP+fDFethPJcNX9GJkrnnd
fQ9VsiG39T0L/2NAIVEsIWzYf7qnUcdhL5Pb0/odyKJZ94q32lgSwt8gv90MhbL2NACS6capTdWu
60WNqy2gHYVGRB8KWOkwdzmBq0luqdIZEzm00aDlR8h2rvF9vh5/aebebHkhOPZ+kolACpXkLbXJ
QmgojCLfVSZZ9a89tYXscHsjl3C9OhcpzX6W3ww4O6NppHAxBBIcS3mgFoAKHtrKJj3NP4NHg3ft
92Y2TRn2wU29DgAGKCaTuKEE2vpkzs0Z4O0hyPcN83FRPWzvHex8DrRR3bUolhwquyAysF06w9oN
Cvw444oiKK27y9ppvgtCNliOzQtVSmcq+SQ31e4KCcI/rARa/7mue5wbczPvfo2MDibSqrV/ilOm
SkuiVcnVYPXdtDW9p1e1HRkGeVEhCkBTnj88t+2uMdvAdYg6NhZI1iz5HIPMttyHBslO77gNgZnS
InmjJq40KYkVvZH9pYirrFx9/SU5fWQUSus9iRlnG07Z7wtUtWjJ/GYmCeZaAC5yfYJVDRoA9WPe
OrkIqbgsnDcNX4XYKeghONlVH2M3K+WIENTc1YPd+8oZ3wj6yIIm+vnRch2maMJCmWigFuWYMtoV
oBsdKwhWnwTz+IQh2vsoyZ+WtjEoO9Aehq+RdKhGdX3CLXNGL8tHYOJkO7DD2filw2067TUHzFWJ
5w9eQsmgd++CgX9ITBsZGze7zkOIXKfvJN40nviwi7OQ+iYou7bv+StbHYFhseIx1Z6J9xS5pAwN
+LSxWb7HordziVv+3DCw70ohneyEDWqIH60d2X1ovDWnscr4unJqvOK1y5JpACOCcCMTWlNCV5CT
D3llBKA1R2DBQ2VSejmtT22rUch/b5StHFTlHxusj5Bfx9X0SixYht8XrcOcAbyhGa3n5iY1550f
Npqld6FnTKWdOElzDJvJv4rOc6q2oDNbXGQkXj61ZpF/wFl7YlcBZq31oilhB9nS8+pZVX/4tmlQ
CFD9Egm3UDGdIVK9wj1k0omDV3S3HubsDzuUI2pU+QsV6JY4oxAukkfdtCHiB1W6uFt0EvGQ2glV
gGOwaYh5Jt9qckEBonXOUkcyRHlTZ05ZBJ8uXXE2LQBHzoKRJOheQurVA9kcVv6SmT71F9oqmqwM
IebXhr2QslOY9HvS+6Ccw7QxuSR7aHmUFIwZeyc5b5D0/yA4ZNnZnAx1Ortwu1YlJgHbyZsOh8lF
ObO16IvOXwL8MZS8zaoQaGJOvaa7dwAhcYYBw5i4jVY7duUw2Y8CHxmeD04/xcAbDTwnF9Js79oc
pYMblbUAMYDvi/Y4RRi0OzN3DoKNCZVcf6+wMqEhABqlZDxCoV9u5cLnA4e7nhVkxgRPgTmSG7JR
Um57DjmfZabcxg8MuCGnsIoHm0IG9edk/d1YZXPPnZdJy6ZhGeKEPf8/IFLz9RvD5KusX9mxDVqo
sjqYm6zhq/1/M04MMx0WBM7L8hGbMgfKlikjF9d0aiBZt1QsxnXkd5iL1hW0BHu499LYg0PVkFpm
yWDiiBQ5jrs125yMzMf1l8VUVd0rvQh7ookUSIvafjzGHEi8TPmdT5A95aQReKZ8/7OwnyPqqQzQ
XbfYVAJeTEHX55k33RpTM2biCq/AeqBCVQN8AwPCpmEFZZx/JEajk4/R536n/0Yi+L58zpdXwU0t
obyfXTjQkfWhCXAZhCjNa5IyQM0W5SNvdlScJPR1stZWIAKXsipYDndSDGk6jNchf+K2iJKRl8IN
y4oyFAPa89jCU4e8httoGifG0CFws0a18lf54MBt8Fw0cndBp4iUQ/qj43UpIcTL0n5iLQygYNyo
2CldSsy6ywZeTPOPBnGe7ZnTLWZVdCa3u6Ky7A7jIKlYsUPKWRF6LfKHXjSUo8LAQwCRCw6M2KQr
2eUbdjmnUIQhmJevRFabkx40j7PUv1JbvmYJo3qwJ8Mul2x3Hha/lFisGA1Yb91+YCD+ZXmMOA99
Y1AH/bTDrUj/zZ3i8l5T0sLCO3lgicvuQlKcadr125SHGj5/xGuF7kYdZIF2nVwgRWFKDnPO5ITu
YCcsWoniM7EgAcvfFk88LkLAf4kCeRD10JtVVBIoqePvL8PMIiwIPfgQ9Mbp2UV3/hbj1yCQNrKv
Y4AL5W+doNSRtB+sPKLW74f1oSFXY2fT43HeVLjk7rT7CK6sVlnY1Old1rrJgdTQPD/OOW7FA599
5Cd2xzSXv9fsPjYS7qhbO1E79zzgd3ab2+Yy6/uFbQU8+MTPFbMOAZpcSOU5vE3WSbeW9MlEMUOO
QVhYM5I2r/h+njqMLhzqlvgiY6EUZcIet53aFGT8PKUAXaFWaREtctZ0M5scdYxKpsyiiJfcYg9X
0Kl8w2J3FCTJiMvmZOIgCOKsJ7z/wcT3PIiNu1eSwGMfrK2zcB2BXmG7N04FSroDqiGV+iFYhDWi
5Ai97JiwEQmbZy6yae5Ne/AUv0oxBfGgHEUXKh18QoO+G+SS+GSonqz8lzW2pXj72WJnf6cg8uks
hUKqF0KoliZcsMvgXHpvsAZ9vVc83RSRLZrCFTTOO4qoOh3hESaulu+ucI5MCHGSxUa4VREmj9S8
D2kJWQSbjJKXB2Fgaus1LhFLxQchnOeeB6JzvVDZKQtwVDKvLOk+UxshxXpcPaeTPbgnWCcEC7Yj
SEUuBg4TfKabNk3ATSDFBPpQ/xeixd7PNX/CEvIACHZFh6Wg0uDF4HI9vg9wdr4gCcrhUzxr/CjG
j6Ui+8EhT8PJrYsgxSj7h4OfQuUTmBSll4hCryz6+ljoGckiBrGldrFxh84QVPIZyt8hiKQOK0dl
Ct/WnPPUJ0K7LMNdrN35whoZkzHZn4tMVuwAk/eQd4wY+MqMFe7T2ZvmKJ64O4gO+5XqCKYZx0Dq
yOD/GIdVZwCXAZEcYnvJ58iaKdasCJvi4MG1S25tjjUrF/00GEpic49K3F+TliuwG9hry2Bz0eh2
fbMfJ+eKYbWQvIxNLgyQdsbNOldHTGyrwoItYu7TjtuQX1Hh0q6DyfGIQtbLpI7fQezcZQD8KLUB
ujTZxbZVz7yvbSDfNKKXGx3hjxxzHaQZ9q32zrVMdwz3PAxs67FuUU9YA0y61yCA1oeZ+QkjXoK1
3xIhwq/0HB0jkH52On0Gfwcy9dp8Pfbx9BxIrlcpzskqt5WsvGHvVYz+nu0t5v6ESEkO5NkZ3UQt
Vtdjhq7enS0nihhGwrF7T2DUoww/dx5LYXHRJXUfbiQzyjt0bQkznYpgilwRc2OvdJAwHIpJi8Y4
1JtrKywKmuTWDzbDPtBl+eCD+AP1kDNu1YSirl+kwuYffIm3xRC+zVWkM2vZvKoWB0Vi5MNTzGt3
hwz+JLmcLEpNsXCz74PaBCI/6apI37Fz+CCCBd8yoK+Mov4dwvxcVj06TqLnQEgHMPqd3zANDCKT
xDAjyQSI9wm/ep4ryumZXwrjiuBJuviT2U8c8niqvoCB1rI16JnMuXim4E1T74unR116J3qyrD9Q
m5zLZmiMGZXwsBhqB7FCfmTmFLDjqUMPAEeeqP4bkarYHcHApRmjwDjnsZ3/yURHWRLkvkrrQ43v
oZN3uew7dDFQ1vZ2ste52rxKAfPrQYqxCB2iBDxd1WnmPqWK6/nTA/5zfdWTYl1jD/GUqDcTmCRH
+YQmi9qrgqPpRjt2EHT8vO2F9VSxRl6jfHBdzb5E3Lu6yBWsE5TCH0dHMQZ8y5lcl9pIQCmxuXfc
hHRXvL9I68s3xsFjhEfjg/k/Az64AmbdnmStgbm98ZIqgCmKg2DFUNVen2NrMJ4cuusnsoS0wl5R
EAwExNA5yH67wsotnSqRMeDxvV1Z9QKN8ZPZlWzj1nWEPqeF4c8Q9fDfb3+rKB+yDz7A9OKLXia0
rfv7lBFZrwcP/GHr5U1+WI+AYGqxCtsijnBPjbEos5tDqgeV5oygSlDyrzPyI3S0QleWuIqb1MAE
ppjyM7f/p07IGMEOve1Q362zgjzB/D9QFNdQS8uUA5A0/X++A0dBF4gYgR5YqR5Zz5DzstKCPoht
tMRn1XC9ap3QHt2ywDt+yxbhoiuVpMHMfDNKk5gi1LzXrvzRy4NbPwdua6M8xwVjjq6vrC1ZgoiV
SP58qaDwchYLNgtxK67TKHVvwY/u9bJk9YgJxK43o8Mzh5wD+wWbZkiLjBVkaiFQgMQDV5KgFBhv
FmusyudO3j5wohmAuYmTyTa1FlhW6hk9PkjMieh4yrhPRv7w8Dr+b0n2+wcEy+1si/Ml2oSfoTj/
r+3JkmmnRKsHIAHLbOVbFDqmHOBmqJOKNF6Ay+K5kvJXzUH7CmGaH1W2C9RHRXxlEmiFzR/Afn5+
jHzp+W6o6OrR756rBVWmlPX607ez4hYWhK7Roxn/e4fl6Eh78FfQJGJFuG4UfqtEo36IXFtrDi6O
HyA5r/J+5DQ+WJGdE7PlLQTvdibO5BFeoBVVJKDnUGsqomnWyWuH9h4+tC16U+Iq99SJklDfxI0c
5iQ1pDmg0nUFD5/xVf20shKXfhUP/7uGXqbFO69FXliXLeccRUvhsTGi21gv2F22bLzHcoHz7G9d
AHvPQTE+jmaAYz6LYkJ8l+pmgXJnfQWa4rf168YkOTuWA0Su97WPmRVlRDb3Dv5RBY5Af4X9lQda
wKv4spbQhr7Xv78zFmXiYsuZn4FEjR36q/VKs7lGPnmZ69blqPaUDbpBGDvN43c6TVht0pfL1Ipc
OzeB9WNMbybLynyb/bsKfAEjOlMij6jiRG/8WSfvR9vGJldiLx7pB+7P7+bzlJv1ve7JKneIJ3Ro
t+Ntnf1/20Z8XbU3BMQ6xgDha5jDX83M47ySvjUeR2LrG3ivDPWnE78f5T1Mb0ZnyvGrsS1JRY33
jTfJDBDJh5wrPsfmFTkPya5Pk5wzxlFRnLB9MM2mYXeINXszzm6wLJb5e8yEiYxMrfgSGZfktjVr
7EIV7fGKvnBUIcE4TKDCsqwASz73FJtUUNl5e91+mNOM2l51fCswC2l+9+MBjAc81kz/WMQhS6QQ
ox/n5Qs3Lj/1p06/JzZg/PKDAn6A1fyI+V3PYsfhAq4BlOKeMQf3159fmFGOQiZU4neZz9E+uXLR
O7nLmq0BKPz16THQdVlTaJeQxBDsP77ITa2APAROoopnwUMr3tVA3jhVxJQknZutqNx9DLScd/+X
1ISQXALsNwVAV2VRhLr97R5IH+qKahpls7TerEUP0gBs8qheKCl9dKKWMbgf42YyC77JrI0eY07o
xt1NTbfxqGe2HHAGB+x0sa4648S5jr8D3pjt904wlt81XhGnVdA/Y/1zcIR4Fcq2Ywo1ANWK1hyu
erJAa9tcejxff1mkSdFMwVubRumhlCqyDDLokIYjFYXE6+4hnkhm9fSq/TYQ/3PnKOqneOHg0qYT
2YFCOsEUo2mlmyZwVUItEjk9mR0Lp/t6W63K7cZmxBT8SGTTFnl6ef1ijjjxuizuDRLMtnxutJr+
ynGy2slzw0/kkyB4zpZbmmaItduXhNhjgObl3kTrJmHDKeiDmoXWhfUPWWsxvQtHRIVNnNa+VL2a
7KeO3I9J0iwWRMlJKyszD3H27lTE1R2KvMOYEjpQ0yK9BQuMsSdvaRGGyUSGj/jLQnFKAAy1lRoN
SnYk3tmE7Jc9Td6ykvuSXdEKZBR1Tq61yquxNcu/k+WaH52pKu/BcSgQe1f6jvrazbkhMaTSj+6N
RGxqC3LEGNz9rCyXTuPlMMABiG870qTUTZVIK/n90sMPYPW1sEZMrzZlUMcO5NYa+QM1LOg3Xyz6
MxDAysKOUiuXNuW8QJzQTX+0sHuX+7AegnsSKGItPXjZ9qzexUPS9S8it4THZNE5OUqphJCvwPhS
7IQRWjoxrDT74xzcYyuv98T1xq0mQkJUK6RLDm4TWjVRjx+e77L5+0n1cs93IRaUZeDMbCSGhmP2
6N8HYgYWC6+EsWO9HZH0hcrkuH8jSMxT2wJivkX3oGAVs7Sy7hYMh+pModVDqLq4TDQWU31stKh0
UdUZQ4Hl0P/R0OfPP2nH3pVznkyKVQr3BMTDqZOIof18cvfC0MR4KPecp8aaJ1d8sMqw8amrZOep
JfUXtEGtB1Kkw6QGpE83oxH4LVlPqOnuoTia8n8GKci5M/L1VpyJXd82aeBLD0BmzBki5U5CkTPO
pCdFu08PrSDDUJbQgpR75J3oNzkPyMLOpXv2CE/i/A+V2p17SAxNlKkenK0K9f5YO/vBGXz0qKx4
eWyTUDqy/RWfoWCfLfvvuW2Rpsw2G9iXgx4x6CXCLE2sO1v9swahHlmk/NckT/J3umFc1OsXEe01
um6Y0L/MczKS4xPY0jYObhKa1gfBSkHsLESj6Rqqdwic7h0It5P+sDWBcpoXj/7seRMkyitj69S2
ZI4oUA8CULZig6tGmayMMH+roAqK/3XSW5ZlZ3OHHyHQUkzJFGEPdlzHXU5dXuKy4XMzBzHjggSH
ZlDoNYYwSjRSh9pMez7nujawAYSWAFfzp+1+/XnE6Ixk4VnTHjx6gXvBqC0IaRxcU0CQMkHfR4zp
u3p3jE1qDYBEzzjN/C60NRbFpxM0BxdFdUW9CJEx3uPSlV4/jn9nABNZQPk6CxWS5iwjq4yTF3Pp
dclUXd85zYwONYzJTnT6yLOfkWa7czuFj+bxAnd6Y6AvpJDIT0dIQaV+ifopjVMx+EEYUhIIObIU
NO6Tk5VXDuq4IcGS1sLBB/qVvLvBl+WBBqGYn0sfAT2ZXgc2pgGtLtz5gZZXyIzc4yRBZYIBScsH
0jUXdNj5va5QHPDv395Ps5vWKzc8mJkJesncnOxm1BbE75pk4vdNtUMjqV8BWoDtsrqlqDvdwIbE
2Nj19gQ/hE1P23+MGE+oL/VgsoZMNdV1iTkg+u4TQrVqyIMCWQHiCk6ypcACMShHVs7S0k1UbOZj
XeULD5p9G4TSJUXSiU/7FqSubISOKwGq8fzj87L6vyhAgzRa/XCxfqdXU23XqHfUUeFCsXlJ9ksR
LgCcXQ3pgZo1XXwEFMeIzpmlRUJhyLCUF0ACzlAPCcwPnhxoUqauXECIN6QfO8YZ5dai9b26iD5Y
4SRz0kE9hukuFs/R5wLBIgCSfZ+v34C7kPFEo1yB/cnnZjvZ0UugmTePR+9pdiS++3eU+gE2h2uS
YfDeY0q+oXzTNdUKXdj/UMqueprmHY98H/PsJ/hjPvF4wnypn9IBForyO9mpM34LT6gUSB/oY51f
sWUxb4zItEsGAYkMyj5vr7Mn1mLjAKOqm+FMaF99lEwrJzmYpUBBmxVwK0H6Gyn9OQBz9HCAFFhM
/QdLj0IuSRrqRCKd7LbCvJn6+Q9A0i3Os3K3TuTT0QLkVFfnwGLUhowYQ0pwvnyq1VlEju+sROfS
d1gSolz5xEyliTXU3++hu0bFxEZFaJwbCxTsloZteFitbmRr1QrjUOe5LBnzt3Ec7Tjb0mz9Z91i
E3Q9qb3bzCyqH3PG2TTsPf36g+AnXct1qETA62XX97H89x358837/tVkEKP0095DE0eH98We5g92
2Asg2p6YpHwYw/zga9Ply2vl4eI446+VCUZpEQCgY9qlyD6PpLRDm66GKss7q2aHLB4VSr8gZtvi
AFMnnp5HcdkN/6w7eoKxceJacGUwcfSW7u7AC8jwyF5KgxPgeBCVkCaOlY+2EStEOWl9j/BWAbqt
H8LJZf9yH1SkUionL92R5KZ0tATC4pL29OaDu0BBpLl9IbU5TljK1DlKPxE0ZU3C2b9qG/jnKhWv
5IWRllHMlQU9WkV/zcFH01K+03tHSO23Xum2y7TsMXQXuERSSB9BLuZVRVjkFvwE/IrPicj42Owb
pv6XM2gtB+P7YGyhMD7FkkvwE4d+f4B9NUt++syoFuZ94TZw9W1YI5EU29jviRilWjsEDvpqi3ip
o1IaQpO/7L/exxxoeobnXU3NQ8igU86TUxxTDq14337bM+Bj+n8Kmrk34bBK5+TL6S/2WWGdQAnv
aFhWMYfarXyae1qMzD+hzMuzpvtaEYSFqrLvj+N89cspOCkzNIQfY9jns6scb7Xu/h75erGsMQ9+
t1kiqGXffOg2Ee9pEVjAyP7yzeBEk1lZbIAyQci5/V6p/qMjio0mhAEPPgWlsiKVq+nlQRKei2lr
2ChC13N86c/P3g94nr4sALhN+fxj6i8Gs6Z0NOSs92zEacdZoO/s6/dD8WbVNRPiNAXbSe1fBT7Y
ePaMRcGoB4L9SoDv+zeoUkTFIiN8bxqjD0WF0/GEUMx0NrgZnRXPporE+qS5OSTRjAPX/4KtXS+L
C0ahQq/faypEXbMHsRGstqkOYH/UO3RXLvbOMx+RhmoBqE5VR51HaQP9Ta5RvbUjuCpE+G41VS3S
Lf2b7J8L0g2H1dtr/1z+RrkjFxMkXhcMilVAyLjj4aOt0KFgILs8aX2kC+H6vpFGjdo6JOv7D+e7
hLgnrGXBEPrHtONllZF1vAyO30liWL60zJYwfonfCbOHzQgBb5YiaNv3TEd4VbbD134COaQ1eRMT
qp2S/nj6VfqHvdPEtgLju0U73lLUlK0O43HJ6+in/mD8y6diStgZRXiO0fW5hGUQMEMFcHXa9zUD
FVOsoGM+/yhGi8okfvOs0rn2SFHmrlRD3B3cL/emuU07l189+FxmYrd7DOpaHVIIUOCz57NZV8q5
51AtDxUK+JHyC0XFI95cAjJ8ExbGt3nhM5TADizsg7xseP+VvmC6kwKDtu+0cxrAhwZhpZ/UpKKY
gyyRZlNsBa70Wq14Im5SimvsXfU2Qj/LrHGYOVSI/HewLXIhi9sxMmw5mr6TVWbpywIWbjQnknrP
I2hoKr+XJtVOuVDY+Xe2tK/imPNqlUn2D0evpqB2O+pjqhyr9hrmseffqP8nJNwo9GI+yhc/alkU
hyBCXVeAlJ4RyNUaHsxi/50rXC6UF/P5EkSw49nAR8ikSEbwOTw6uBFZPLGt8qgZKxz5ABpSfqrD
ung34/8G4SwynZKrIwyBKooLGv/CRejMrJqKD6RMirw2j1JPwSnio83aNv1z9ZpKG2LXXq6AXqCG
mRJtviqJP427p3tAspe+s1d+rs0u8Hux4X08fIFwp33fDd9iDptxq+8lLjqPZuCJl/Fi+wVweweR
KtV3zoKhOMJySgS9GWpoqTT4DFI4c2anlKUSyPCP62/Uz3QzgRvYrEXgWiCnj92qfWqhQzOFQLYD
ZgYqmQ8Kiv1qwBQSpYt9UiKLAynHWt0wIdrtxNXZu8K0mQR3CFwOlqdHQ4Vvyx4qa8qGEt+vvADx
GnMxTf8i7wm2Zic9nby5dmSz+wi+P8exmb2p1dyTLuZBuX4d8Ckzd97LOu+Qimh6knPcNMeFDXav
KoS1OK3jTiT7CmroX0SKskyTG8HODDL+5NJesPZLNU9NtZEHtYxnAHlCdYIgduHZSA0egiWcTFtl
Q3SCmgruXFOh+4kXvlLyTWH4EYaMsWFEQheNlcoGSBvjjBUea4sF1X0+z366mwVWF9cfJlshLcOY
KxNowT1ZOGY8pqk1Nrp922IFPfxiQY+GXtMDzIKtgSBTrPtUYOlhSBVmD00ml+MTabYz7XfE2odE
atMc1Mm4FLNxkbHcahx1qVZWHOZk0EN/bO0NQmKVg3/2qiSogtFC1Z7h278CVrxHl1g2GQdzy5RT
EbwH8nN00D7TwoovvFcncbxzD5MbRGdQiRxQUGdZw46aSqattNmwhxu+yVmvY0TCzBN3hjxK4i7y
2l1T1mgq8/rV5DibErUw7gNn6WqS6YAgk6bPvYIqFl4hJmaYza5cEhAS7zSZZxNvoQ8rCGffzvLo
xp1dhZ7rKSbW5qB61DGT8oMPbftdF4a1OZHFlxaJpV6VQ9cgDTgfiLvCSibBauJDi3dGXIHR36I/
GJy0HUrTum3AWBbAskqLbERTlkF57r5kVUq+Zitg6l5q1X1DwUffR0RI6pYWKALIgHYDet8Q8Xsx
q4ObAgunHHew9QAtRIVfzL+LoEO/C9Og7TeVRunAjANQ3qDhMo1Idf7Nhp9ETuKn+1bVhuEMVIEC
7UEKBDEGqARkstai3avR9nMMGPLRCgs8zZWjXhi8LkEiSLCJ+55hYmixesojmhxVbtPahey0wbx7
8eAvFA6v2Dd2YsZNyvk+ZoeuxzqdcLcCKOZPdHG6KdpXuGG7zImbzcTmIfW4oey0LsCTNvPx71D/
WTLLEHZb2RiQw8jbpYFxDrzS/xvrGjY/GPUqrItRVER+ryFuXF/wkzTi/ipOpMwTWEttI9pfg6uH
nzASeWHCdmJHiQYIF8GoV3GOn9VzjiGfhB8UAcxfqVPg1gA5ONqkBpKwowCydM4bONXn5QTD3jmx
2qv1gIfkx74ZPlS+dNZONj6oUB+qShnRlkVzu6nHZZPsdoRxPeCg04W6/Y595pJ3NV1bjhJ2dEU1
DpSrAheW5uh2dJkWMfpXzX3P6c4QMKPw1Pr440LS6ZQCcdNAddz11PxHb0uWxmZVOizNjN9b2suN
15Ywoc5stnjujum0vDaOanqA1b62dW81SZnsi0EcSQKBqOn1z3cZE4DB0e0Rdy4QcNiZqUr89MMf
FAcp3DEZoZ1vzHyaErwHYNnu+oaKy9mhCiz0ieeRt9P/hzXKrZZSNAhspyLFf55NYw4a36BKUBIq
tRFcrvVMv/1/WsUkgci1MK5ISJlr0WNgsNuELm/Cmpl01t09o5g6/LcwpDsPM9Lvc6SFpsmcyGIc
TKkWql00g7eo6lH62kDLhy0UIZ4I51yjl2yIKm4tot6PFH3qQJ2DFeGez6FO3HvHqnXMcQ8Ije96
0Mk17oXV1+d0G8AWt+IJyBxTcM72sjzOAjH26qSScCNk+Qjr5sdtKR7zL1F4HYzgJCz1ybJ2n6lP
XQc0Ty/6P6loCSYLlE3+55dNhsCjQDaiq/VhU/VtaTMtttGpm9a6/7L8JXrMki2mAzJpgpSmqFdA
7dNCKdNTwpTAYCg4k34fbdQl+JpkLVQPJCHAk/fCSNIU8tnZkarheBrJnf8L7cdNXXKFo7QppHPs
WcqY0gI2Gg5qaoPogjCYkcNSqT3Lz5WSudG6VTAUB7PlRBn9nom1RzEF/papoqur51HpSmQtSCjB
n6JVKLErm07MUAmgjABHmHpZFgqiag4/oUHRhxiwDzmsTv3ky54dm3Rfvz5kXLmDGLt64n7eT/Tl
Whaj/KD81H238R/GP2Wyq8G7qSWqHFGUH5YaFzDnjqjz1wKo3IKxmAka0f1dCZdHqUD+tDHaOSj5
dNghLrESMSdoCBkElogb7cAOMtxjcLr54Mqhe4HHVR5p3SsfMBHOUz2qpM1stQ+bIFz7Ce0pWl9h
ymUwV/Gssu/o4CGwZdnjlZvVQtYkroJEKdp4cSz9Nru+ApG5bWfEGwtgkI9kPC53OQ2WiiEOh2dc
7IAIr+tgvCb8/MYfnBTpIChE3WZ/4w1SMVmIbUVQPO4B063VW3GgCXEmH0TO87ENIrocLIWLOeKn
DZ7slIgaxZFJQrMRDgk8ma5fQ9gNm4XxiaDBfGGZPY+XOAsCoTlKc30JI10+LwiqD6HAqhTzb8Az
Rj7GJQHS6TgAVceU9cFVDqVwIqtqLL6qc9ilWumzlkyH4BmT8XTn9yDt024pD3pf8Al6oZRG2TEO
FGhpuYfmkfQ7ojFn2gfY7qOCTCaGhGlNaXNHuLABZCkTFHnfNLwwvRnz/eqIL0hmHZsyJy64idx6
1nYitK9W6GucZsHazE3ynoQUccg6nC9bWzqKkbLwpb2VoDkrOHFFJb9vxVDbFrgsUQuVY6c4yrQ0
xaLjrbrANbHse8SMFEd+YHv0d1uoXptP/5UxpnN6LKdwrfP6TRU/jnnpeq3JhYnukE7CLgyqUixV
Yz5J0uViv+MUsZoju/T/P/+Gs0AoNTm1VWLQa94YRcmfWYT+x8oEM1nptss+Eco/K8zYprv0Sgy4
JiCPa9sgmsJ+ywnnQ4ek1xl0bzlub209UYtVItLBw5wlY0OM3MraDDgwPfr02iIZLc+8ziYpcZ25
OrJiVR5boHg0kpQuaqeglUu4LdG2n0h+T0RQsp8aBo9uF8HImCw78tGps2W6xoDGjA/fsa39/MbK
6QHQlRBhagVDA38A7B8SB/L9Vdee7hpHjk/7WvfMNUPnW1llj1+xEDWz9WMvAtoRweLqO2scEi2X
JZNLBC6L8QftyTNd/IFMKSaIfGSVKaMH2jdDx8Ty4YOazply7EjNhUfbsXNhZZKiYt8p6cKlkufH
VkG/kb/gmJ8ngjD+eq23uTP4rGRwqrOGZK0+XwpMc4QycomGhBvO408IinsSVvLhAKBYcosWTXoe
+E388rrn88/YDbrZzIlDTPg5uOYiBW48a/GBm7XG8cWQvfIcuKqoCm7Dfjln8+OA+k+BMyaoPrAm
aUsnAfghlfCLwKS0fUDjGLLnnSwiSg6rIbcByBuU1xFOxZye6VmfO7RGOOSwyPNp6qaOvukSDgC8
ppUXIfVHLOPYrNE9pmgpXjMtpNKEMLcRoZd8CTMD8mSkf+gTN89/6TZbS6Xs0QTNGrCNnc9UEKi6
wXBhPYN+erPa2YtNVFnWKegFrT2u7yY4bSpKRWLRkDhxTc991gY8HkgpHTPIfxSOiuDNTpXGFsa+
TbWC5+JfGItJ7qMgg7JgMoM32goN8GeQveCz92KPIA+EtOLCrXLnJPJSLO0SZ8Zk8S4TWZeq5Prk
Sqp51bGxreAp/VyFFr7PKZWtbzT9vQXWC4vvBOky6ATHYhBzJp8C/wgssGlPYit7KSFO2+DTPnCx
odzYSeDG8PtJE6/qiYRKtaLB7bEL87b+mWR5TGGJA6az8pGKG1cOVSSlkRPJNVAvJvu4+1234gVf
TxH91nc+cy9krkWdYGyPRSi5UIuOPZT8+fipUp7Rb9A2oAQPBx1Joow/KXUVQPjHWyqoiWhOrFC5
chHFlnQZ3DTDd88V1NbXXVJ+McZYge5NC+s1/8lwCMW82HIWUZxqqt9lzjreJw6aQp/hUF17UVmR
KV3IMzcLCMHqRAH2Xyicu27A2TYXQcrin90Jq1IYTeZwM4YzwU6Aei0ff0n5QaTwvchxyxI8Jwxv
8UBQCYaXzprOpwLVL5ezEPvf135dRgkZB+AXgHqw1uoROeeJt08Ms0Qq3G4RJnjq2jxAo5kh0TOH
yLteNu9yFXr4l49mReLgHot5mhs7d6X2UQEZEyh5rLKFBAqNfIRfD6eGdw054FQRpbNOGmqJb7JS
jqe7ybN18ftJ396Fuy2h0MU1aCdGvHVDFRy6aDHLZEXaOPQKGgre41jpF3x7S8tjcFu0knSGO63r
KEoKELXl4XlcB9J21zAuYM8KlY/8Dvqvh1Qaf5DJkKN2auUseQJV1rlxNNopiayS0rcvK4/Z2L3j
F85Tz7xLvdnQHcwoj7pA/skfAa/5vlR3PtykgmKDb5gDxAaxzVAXkRjJmdpfBoXWUgwqNvf0BPPH
pApkvg1PBIINtptGBJJKRykaswRjU5pQ2raCp0QgnslOodgJT2E7mOgNi6SLDHUZzNCdS1Vnvu2X
YNjzWh3LABN40dmexaOwEwmDDTIEaWtwSgd1ly1tA5tqP5j7Uij2vNJ2uPJemysu/542mHhJT1tW
hCD5Sl0ZE3DntQbpoLDPvPh0JqqCYr/b6YXIfWJSDnA+3ZZqb+qZpLUevAL7dKhrjuzpW6GCgGhp
N1cm2yUGohatw3Bp09lwScvxr0Hxop5DNliwpYjK+3LiuSCdpxH8YSVTW4ywdOU2gXfTyf1ZXqtX
G93ZMCydhF7EtoH9THjyFMT0UBWxBDXj9Y4YbbXvczGFdcdH9vUSYDzqfnjMB1kIJzOu0PILLnsX
7C1i5ZKXIusSdnu78N41HwFE/QvEQbDMDCFOZG3TMW7Xtl9uMi7tptvePsoUozN3hUjreKKDoUsl
lqSIleBku7vXAhtVrzy2HO7Re7bEciTEfNemi9VgXh0njrxj7CfHOFJ1TlBaS31C1Jd9jbFLm5iN
vjjz7cbrZbtGe6sP2JnOXx9CNHsWZDdwcSF/476hG0VSSgcbJdH3hl8KXbuQOqAqvOlvuQ4gcBsp
jxgcCBznq8FzucxetlNxXRj3DFgoxrB9axkWXG6FRQyf2E90E6PvDtUDNY7Ylkh2+uf6wbAmUAp3
MQrBP48AgIqotkUM9wBaGm0me6S9NeqUIdlV/cu5BJIqbE3Ym23AZRLVFLg1GiaGxzVpQYdunlUL
moMj5mL4d3YrQMdqumeQrRGQZH6pAheEoFHOTmVwhAFBPENXndX1xsjlgXdsL5vi44GA4XYTHY8a
Pl0/XWexEiDJn0Nr9nasdJbJ75BoVKbz+Es/4hXwrcInRuK2RDHx2Fgq1t8ZXe9n7zcI45gng4Rj
KTd4eU2TBhCoOh56iV4/mPD4A1U+Yn9/AvfALJ+/nHS/swJJz0QpHLsFlvJnhgDSzXpgC5jBfM0Y
R2mMIUWxb4MfovqBvEnSveqn7Uhx6FIwgnBlts5HY8GoMh1+LD27/ZY5vhRjuYlqPIZB4XqKe79J
2HG5aD+x2hodyLoyolziOoHG8o12UoeDmcXBFFpJyMVMf40FXISNUJ8WYFDXbpfagxKOnmMBh7LA
NifU5BV1T4wXwQnK4rbLLW6s85O8HWV5uOJEmxjS+WNyRmXFziBoQ5/CCmLyIHhtlmP/jUsdTCyM
Z31ZnIrZHutg0gp2nqWWqe5EHHCvg2QbEsrNpouuEMMvSfhw9pVt9mnEuKP6VwiZ/cutt2py83ol
/5e4WgmYeUlZzA5ceojYkd9j/XzZGIthHe4gVnyXDNjM2kV0wg+wOTySnAI/VfMTT8qN9byedh3w
nL+3hZXorMad2N44e5Cq4FCd9qRJHrNZT9DyhoiSauwohNia8JEQyleY1jCuCFTyaeR4IwtwqGON
lbm8aL2SACKAJiOl124Eu+2VkaRdlwgZYu6zPnFzm4AadJdppc5dgxQrIcbqhPNPbCGrpJtqFECq
xmybw823peNc1+v/s8iN5snk0bhTeOfNj7MzmZ9rf2LtCfOLm2eWv4gqaH4+x0slxc9RiuZhrC/1
0SvtfVUOc1/7sd6jdgdopWtFzs5DfTiE6XxygjbPKEYGUwUJAqdI7I1fD909lkybQ7hUJ8k4Znef
aBJTdS6fXh6OgAESS2PievQvVLKOH+6uCPAw15+Xm3JsqMRUeDmn22Zb3IjPuEVvxdA6HXFDDfZ+
nJFn7lxeUiTguYa4e1TGhAzIbwIdWJL9MqTaZhsS8Dx5vUyzdYL7FFTg52tew5eUNZHf45Vf6bRG
F56VFixX0802W3GWYtEMl50fQphiblRm7A9bYHSvffLVgURPAG1FuW33coiOid7tlkZL+UNsSZ+2
qVcU6+Il7ssZB6QOxIW5C0QDyC7T1SZ43+n3BWwD97OEYfj1j+ON4dfd445vRTRn8ttASJr+ROt/
5vxxhWZY+wguSfIKUJ07zkeCsx2xhfMArWar3VnLmxgoqItQy/pJif8HexgcJjmZr7cKIkwmPIR3
ycHVxpL8Jo6OQAgvBSbVLoI78raZWOwHsQkBnWjqAfQQwUfi6J+HY2QGpwXgoJCLW9YGn9q2iyhL
t88n6lXnfKBMCk2pNalLshHod/2wmywbjbmY4oqHeNmid/H8x33zB0CV5BGIesQa1y55UzOeYf1O
XYaYjIg7ljScF2qjK24SV4gu9qAMqViXfWksazkKJ2XwZKongl5ky5UjfQtJwCVDynm1cgCc2Ba6
1poMMbbQb2dRpKR1md6pt0uFZjY9Sw9SZk93byONP0+d+QbbcIb+Z82r/8QLf1yuDLff3995oU9o
ZPVpPxqbQ42aloJBYDAs6V2CLF4CY6dIw8WBuewqd+uVBXAlVJcHYvG1uuKAntf8ecKETyuA9+No
LoCzUUQDCarqXqA7XyEKEZ+oXrSIKgX5gw4H2hmFmwzM5AxAtoTWrmwANfkPd4OUqmBgOyVtysE7
0793NX2aVg+vvOYEkufIk/5/JJ9Mb6jE40TfXcFecY3FKtDttgJTuWeUeYX8RukZ8C/b8X9iZQ9f
pTMqY93NhJIqge7EdK37+cBRgDyTKiEdyuyR5ar6tYL+RYJQ6MwEx+2CILbantCK7u1cpT6reP6g
Ht/ExZcA1EuixXvI0FZ+M2RoxOG+yv6riGM1QcDZbGlA+8LM+K1YSCLhucN/rrW7TwrbBgepMt4m
OLiM7814nbbpDGXdkBBYSRVtJXirm3WL+xWVFcoAibC9n8lfdvYfRJpWJUN0+KiJEuqFfNQ1pqO+
X2CJ3iWBzhVMj2+XdWG1fvMAI83W6RuHYqXp7ozzA88huysa2/UrBS2LVc1Q3OLpcvcGjdyyUrTJ
iTIuUgL+1MJmybqAVBPtDfD5m4xWNQ2T9oTV0OVTKxFx8+GVnW+sQDqYLva0G/t7SMjTYV2SjTW7
YIn8SK5EGLujikJyq9nRi31Slra4qEAvW9w/ExFmGBuxkWLr8u8HGnWZZqV7ri/O14WRT4nqRNtq
qrAX8+rS2dPVBRqUO+0PZ06zJk8/u6ZgISKAkqeNoFXm3ptRJAJlxXc3g9PCuGqSxafqNKDbw4vz
toyrOekoh6ebwNpdzYQCbvDGhSi2NAYpvDACAd43qgVowktNtpY2o7bbYqfgi0LY64weQ7JZSwY0
grTX2SPmxKSP07T4kPTPYkjNaLj0E0bhEPEj6Yzfaj0QxfFNpR1Dgcidn4NzLKwnNKs6S0GIs/5b
34+AuW0ZAB9mEScKbKMeubLtLRWz8T2p7rnii4c23BCK5GCjoUlzD+B+kKUP+SF13ZDNrBG7NGmD
S2SuxrvxdRXK3PO4V0f1ZG+vQoFmiKO1CdoxqNK0IQON5uGnY0xTYAyBBEfTYQ0OA2Wy2JjmlqM9
8Bcbcb8BrZ0QigQInCRik5ew8oJCuiJoEZJbN0Y+LoeYkjD1wRzlXh2UEcWdTOksuQ9rCQgkket0
GZLcmFUbl8ZQUhZ5B/ysoKaCvM9lapjDeAY2PJzjtT5bmLCt0I4pSUDF1oS9PsTP7tM3v47Yoyom
Wr75bPjMRAF27EIpHliSrrKk+hWCulyE1+fJzm8JXg1aCsg34gkWxp3nmdoIn2OMDtaf8EnDmtLE
ozNyq9VaYgbX4PrI/MvNTC3HIt8aBXEyOM9hrlaxw5GB3w9wXyVrgj1SOduJVX4QRVUzUZ7de53N
gzFQ9jxZLhrvNeG8UKEcOHzvVQYsKr+ohGMh/M3UzNZd8De7DnUzqVQGB1Sb0XczyYZOmS9+k6Qt
9cBMjnqiuZl+/ncF4hnyVXzaU6lNwWRsRTfmd50tCwy+hIfcBsCUyQk9/7WzboRolu/Z7Lk+HfD8
e71SGGwOdyrMqpSBD8eUUv8cUOc3fmWyXdx2GtVNAqd71ewQNjCtB0xMxfgnDlBIKsao86VuwVwH
Si3lf88jUg4qW775Sy1184XhMtoLE8i+PgpNvoyUkV3lSZNRFgdAY/LnACVW/+xgyB1DmTfrKaDx
TzO1X3bcq5/Awh9sB5DWGnuZ91fneje0/zfyxu/HbpPKnhEpRGU8C6FGrMHN/0Nk0JLsJrxrbkCS
KIvrJGliSwDIjBb+h7vIjPxj34mXL8sj5PComC4JaELa8ezpFtcVAwTwyfnliEot1lfoiQj5z+oK
utrnnW/zXtIocc+5C/tR8AMbpnziIKWlB+xGpdYPr1jd9kIcedkrSRGMr4BfZCmoS8yJkw9I45Te
lJb+ISqEPF1tmOdsJ7HTpC6JoKIxF3xngtT2gBIfoftawvrfpmvFhtzdAOdV3IBhu7sUO6AZqNOc
R9bVbZJa4ohboL8rKtLWOQfLYqkDp/tO3tLI4vW9FRkc+waa3NLNWu9bXGYN5Afcazhubyr2Zj4N
caHdQvAtAsGfy/pLGv7rfOFmiXPGxzx6yhyOPv2gaRxCBDmO5WtzSl1xvQsEkD+AD8xkyZOrS01x
EJDahj2pToqnGw3uTv699IxU22FPrTM3+JY7oTmH25dDHmvFUhJ9IN7I62dTI+31ddvF+TpBCARt
swzn0cX/GmgtM/+44K1pOLseE5rlOLnPb+NoFU1ERvcUO4bWz494icJzSDLlwI2rqBR9RJvHsRU3
Wi1xx9m5a/M87TNpiRVUQcb3cg8UcHOAK4K4iZv9Q+YTe14jgSYurq9gdMaNFY4s1XyzLBrErcXD
PJzd8Liy+Qcdry1ihaswgZ6XxFbfpl1RKelVn0Sj+yz9MFtyU5KszrKbJ6lCCX/IUg6ZsQXGmPqb
+b3m9Mf2OLI2I67QCr/27ddRwMWXXxBPobzUxbWI8WVG/p0GjJCco0sZrfBPej+CNzNdVZi6mOcz
fmfPpVSmFnUEZY9hif2dWYlbH+ExjfIJI12Vih+G6Cj1j09pvePLqUnkl3VwmQwSR+nm7jeeJhKy
aDGF0HeAUHmiWEWl3SX1XvB4DJmRoZxqmL2PmGT5j35OUgE8+E648T9sqe+Q1y0tSNgsbsKrVrP7
WaVH5o4PnhDyQNZomJXlTRPh3t69GxNFCTWDJbaVzHdZDejDmqSBdsseTOVUFIJpm8tSWyMR6/+R
yqcrPmnTo6+d5NBR2op7RI52PArW3j0jvXa43XOfqRfnVmTOGX39aHIEgre9qzHl2GWhw8yoKpJN
fMs+BxftEA3r5ku7u/rNlFDkv9lhO1465WYU5WFyjQ8KPTGlFdzmrFlSSYsem7kLaUhFVavPI5TX
48z3YgfkjGvVBCZiO0stRiPk2icTooiA4cNyqtGg2HrsBu5YPt0czvPS8AW2tM84uhUSZhNcSeoI
na5jmSVntlJsjS5Q49EU90JRQjdYfHoUcqZh1bno8U9h3mzULoSgrZH25pRH3LrmfL1CC27qr0bd
bltroz0BaYtHksgD5hKNqUBCrlKN7P+b2GvxuQ4ci5LhsEsK68rI9rRXmR4EHsh/Ih1QX6dLO3Jk
+rv8PNfJZzPn2ekMnKWzVZdo2rdS366tOEHfSR3sXJ4EppDcwSwg90alyIZgHQRwxC6/Q6MTow1f
xwsJ0vrhp2553YgFPsbc37NfS1TAlOWrbcxEL/odDsqO6cnctxq1mCISURUZ+bDpaxdkubArTCzY
E/oN0V1SNU2620TUoLdCSiZ1L55ssUvAYB+1kNrNmDOPTqL0n27pO2CFCbovMFelqeprVdkC+vQA
EKhoIMcScIg1ZUZqjuwzZhOLdlXTwlqfPUeVz1726ooMLUtjnI61onhz4N6qgWvZfLhyK3m+9Rmj
QmnTOyGgy4+QdOEC2Hci1LYlqSVQ3bAUu7xW0IvrlQRth61O4pnnoG6FdliOi3FDv7oX7hkXu2zy
Zgd3l1t8kBx4sCFkURsNlV73GhDJDaHA149RD8G9QnKoI7Ca7ndyZGuBfw0Xpz76skv9Y8nHtmEf
ajGaY7y3bLnKVDrSAEifYVPIqhSVro9EEWipe7WZR66KlbKCkbd9rGMt6GOS4WJBLYhzOz62auGo
Gro8OQlR8DBC2Sg7KVswIoSYdAvNY9adD5Se95sTDOK5cGKtckzjhVFtBcPKb5IXZkj3QLXJS/Ni
MFiAwhkSV5dcEx/JanO9Kt/PQo1nqJ/dvGsrFT+fpqypEmtzFSmOQArypCTTojxWIjOOGxVOdO4a
RNUm6Ox8vkPmMh6UJO9/z/eafhKTwO9gBGTcpElJvcugGMDBL84HFnVLPLSCof4LZQq0FSHzPcq5
P8iF6qaHfvjg9HmiG/Fklew6fFR84mL+te7kAacLqn2PuZ3epqN4DCiEqnr/BTTplIauztUWUirD
ZJje5B51DCmU0L9XpJLtBWTQFfquY13gdMp0v7DL0WCbiF0eaKFHd2Pkwn1//NiZl5B66p2QdnYP
Wg5LsHEhvBhVt3o/QFLNPUttMEjR29k973sS0J5YqSlRHETuw2yWcNTEbG40Hw2NqsPqheOk0374
tUI7qNC8wL+oZmeT87ae53sdL+x2feM1RCCYNw19U+5WWYn83BuXtrsgIjEzOk97XLdwY0Y8FwTA
kjDIW9/E7zXMgZu8brDlIjZWxMRzqkZQNnXbnrCgThJY+/k7n6SKSS4zbKYiQWQtCpm7ap8CCih7
sJzwJjLyHLMRqqYnfRFdhq/WN8TeTQvuVfE5xtjTq66L03AU7QYcj3PaNMx73g9dEjXq0RElBUs2
xdxPWXsZ6IzrOgjTW6myTTxxX+r71F4VwYWlIRE9E8VZecSy3Nk5i9kXgkaDXhAMyPStJ5do6NrF
M7CDfqcfh/CQKS/FzSU+5Fp09Vx+oYEW6FvY311o9DFpZo+K2EO22KqQ7ywMFMMJOg9vBgoC3ZN8
QqSltYtQFZs8fFTT0lzcxVoKgNNqms02d7HwJav7SY2l3A2JTudEzzyrWsJMCP/lBFwHqC0Ff2a4
f+HOIP5bmlj9ULp51/cFE/orQKjZqm8HGJD8W7LoO3G+Sto+8iawMrK2BBwcbPv8D0GwU9dbWMnF
IZE7Oizea9jp+j20JJbfuZQ9RC1G95l72CRACQscm1DqBZbJn5+Iv3rH/s+GekY67FsQ2PysMZdr
RRzP48+XW7lTttj9CInHDsRt92NWW/XusoUG9Gy/KsBonSNc3G7ZbyQRXaCVA8Mzf5JQRsxzP5bM
g2MPX/g2SnLcRODLQfNsCPMzsJZIM3LmH3dX5eHfP6jAp97vDS7GGHPbE3z7HXBIbSezL1JZBqKZ
lHiXVg4NzjkHBffokr2XWadYYZv56vemV0sEKeZOYwGE9SpREcgAqFgk9Z9WbWtOUw8wqluZyQUj
1RaY6D3zxoN0KJNIj3y0BDiu3Dz/4x3DOtqa9FMY8JCjVwRIUfzwUNvfbtZT4VdyAmmfF7k9uvew
c7q0LHJSXs29d4/0SgYblfHier3RxW2jZ6VsyMSwbxsfhUICcS5Yurt9rzj7p7WH6wMnUdDstxrm
zL1H2tasfX9PQIbHC+jaDlxwyxQ84adGkFG5F+TkzA9PxQtIFRHq4/RsDSwLjWiF3A5Hu4kVymlL
sXHtQANqJugmSNJyqJtMUNT8xE97v5XZGqbL4qzz8iv8iZdbWO57hxl0xANdmrukIyBfqzBUCSli
6gCxLh73VPQOaf4cNmZLsrOT92DXuw4mrcGlHlhRj9AcNmZ9T7Y73og0Bhv6GstVRQM235ueAvNp
m7taP4KLgEPyBomX7VqaqpUkUbyLA5xeT6Vf2UQkpF4LOWmYhx7A8R9neqtdzoYMDcnaQFTPW5dF
TLOSnEFzK9gC6dvUiermuykaTJPpzaNy9Pwiqka3rAR7Zyz5PFxZXJigUckHc9hPO878MszjdlN2
y+7HnvF1vsoayyYBUUM4kLqOvRDqhCTbixCmK9nisu5PoFjhQZKm/6pY9h+oLowomOT9Pz6aOZqk
7kkoRjsteE8N/NJDZ7LNqgTWXnXjihFvI5K668sHT4KxYTg2KZdR4/GEt5WDIMWbuibeWVZMrARu
yh0BlQxr2eA+TAfMeTxyINpKqA2qXM8X0s9MJRl+m5RnWHIpTmtIxVHHoC1U6R32VK+PMtgpFMdQ
AMbOIb4QutAV+LkxsSMSi1L2yhcjyj4xu94HF0KAf4t+QzILcnJyCfwhQTQDy99LIDcW4qcauMSJ
W71JJm2WS4PsOxnx7Begk1sBia3BXLqRLm8KClqsaBsrHyaN0xt7YIBy0Sez0dzWB60eZ1YFSnSa
Ud6G9OcoeqzFJB6M2K8iQMhPX+Xw70na8xejKTwlw1YPzwguMolvsK0RiXv99ZUepkLzawZkEq77
JZbYD/wJu8wXO+li2wWbaeRbPWiHRAjHmIilijQOMX6hXN5oPYnItuL/N8YiVHgaT7wSWkXXNG77
+AxfT8/8lExxg23iGRbiSTeM7d4MO1K/NR3doGYrY8OqWX9O+qVI8q99o8ZuuCDk0SyGC4gE8jUU
rWEOxdvDyw2T+ppVOCBl/Ldd0xdk+uI3t5MaTAz84va2msyt9ZbJ0FRrg48ksY3NqYA58lmQiR3o
29EhJWOhzU3qab2CppdR7sxo82mvj+RWxLq99aI3a9F5Hj0Fw/6DDQ1M9ZkfDQYTplTjDcqT+0uV
f75ZTm0lUbJDmUr6nHAP/m6AYH6HMdNctzbdwdTeKy4lOlSCeaCRdThO88sjEbbZgOdEYKSGxiSG
4MPfa6jhl/ZcJuWCJOX2y6Qy4cEOzo3i0CCIkEEJUSkK+9Gk1E4pjA9R/hf72BJN5KpspWDoxr4A
a+re/HRAyF7jHpZfFkkX0eyOFVuEB4QPbjLw4V0pOHNqOCfpa/Zs/kh3aHPa2HdJKaMkrcLjEygw
/ISAJfI5CNCzWDzHygp+vf1H/DIVTcJc+dUxrWhjvLCLwLL71wTlyKewX8+CZUqctUEt8GM5tRe5
QWqxNDaiUV++T6Pd6fJJFcW9UfqqZJ5EWqDrh9jRrrABNQdDbHOYB5TmViIe1ZDNh9aiLuOOeQyA
zece47A2YYlLmG0tWKn0+fHpkN7+3IifXEjJ1pVGuzpQO78GhygKvBLA7ShYqdpqC7WaYGC5+i0c
D1o75nBof3h3IMW64NMPI6QrGx0FFCLeOy9/5SkMHZUz8Nazsk9YsS/QhwXKPVE6LAg3VYnwj55t
PYgNOCGbwBxYf08H32hKoaSw3F4wsIjx1I7IjGSEKdy8L5O9Urcuus40zvbmMl+1DsmIhWR8IYNv
wYWHNiTVTterHy/FJbKb03AgRK6gwtrulspkkFUO2TmWghmRClgJK1G3eatUuQ4LnwRABY7YHsV9
Id8qHEohp+HYSwtELiiIcaMbWilKOdeeLbvv+9oZJvQZnsUX+qTyapR8uqubHFve0dQHKrlXyaPW
81l+l9aJP8cT2gI9541K1stx8HtPjTYLKzg+rNZyODXzRj1bTmKJZY+KS4w+frzEDfg7m/2w3jrY
nEq7do33tj5m4Ng3SQI6ZisxpsPW8zos9H2n4a+EzLdtvvkxqwKpkcaAv+5fXbrzPz+rnriah8pX
Bilm/7QYa/2PwEJ1FKF/mKJZLDocOsqWzhPHH/nVIobwBfV0T2OGq1zSdvkFFG9cYEpn2MMkcEqw
zP+np4i535QA5x3TUR/FP6eUPlEO6xlPKMhnJC3EuCTQIvymiqPwLMXk3+N4xUvR3NnFEmTbPGAe
2kqBFwe4vCqHBuSdrJnsKSPfqzTXvKXxHmsWiI3G5B6FDpfxQxTY1vjq0aB7sve/y8NfMYzwsgrk
5aPBSKfsg6lIp+Fqnb84v9wZOFiT10d+YhJMIrZv0xxcl5Uab/bXYJw1kGabtPRZ4hWlixbIP9qO
a5e15opgZ01H1u+lIeLV/AMdzNEzCNPjkiUiUU8ILFDV/PsZvHpFtalyqYymnQ4bY92qcdmek6Ps
l6JV9TE0A4gXU9gVytGGnXnCuJZKqE52Ph+lv99jFfBCbkLllkb9ddMTn0ERL58gYuU9HZ5pOMtS
4szPv98ddZtB9ftu+U94MeuxF/jJILpbDNy/GAx+YMH7Mnla4fRvkR47z8AxKn1xI+0XcXCko+jd
4ksSiUhObF46V7at4aRL1MeqI9hh412/iY5PGpkqr5hPNTA1AO9n/GA6PV9rL7gE/oTdi+upOYaR
W4D/GctJQYxDNhwF/9GUiVtx1Pgljf0DbcUiXlxDBDkEmtwpTMYjGB8t3qCcHabqY8M2RI+q07s8
KB/SCZjvIBoU8rDVYs5gg8QTOpyFUeIf0ppm0eJRdWIdcJr3uy/yI7nPjr9Jr7OZ++2rMTC6aWfN
ECD99eUTScZMF+3CVioyVFo9sjPmHfcOlYL0XJ47ci/qH73jGK6caKIgPOiSPLo9Fjl63Bf36iCN
rm8WRL6OItDG2g7bzGLEcfsFQZtabjyZ0ukyLi10eS122AjIWCMb1yI86+XIrF38iYML+CAO57Fo
/4FC0txTcDU4xUq0MfmzGUX0sj4v7RpkyWTrjOPczdrX14wTE/s54p3/fJndYrkQHweEvY9dIMQE
UzN5JOKTW+QMoNRO1pmQ95kONiMk6+ls2uD0sILuwxj+rSygFVi2aE+ugQbqd3pbAgouJSN4MgtJ
UbWEfx65iWQEkCYFJNAkQ4N4O00rd9+sMuumx8ixSD9uo82Q7LyfcDLIu+5PO2KKZrKMwHfCDw6l
noPbLv1abgZJ1nVrV9NGwfVfLUfojFWlW0RjY2rzJiMCTWePiSsh6yWsxR8pLALEoW4RuxinKQoz
CatCjc7fZsZYN2kJR/zS4+b6qm0JMP8Yc+LH2Qn/Ex5gCqHzh5JzLuwJSa3SXkxGBUjseBQQj4T8
qQuRLPTnuigs2JIj/1MsbnCcVEy8lT34pGYBiYOnwdyAyQKbWZA9bkNs7TBDA7yFXG4Ul3XjmSZY
G17MvKlmpCRQR0TV/B1dA7ZFSAN+ybAbg1GvD/QZu2cy4JRPh1cLfoaj74bB5suhm2QdqoWmG2EG
qaNz1q96Dk+PYqSXTsd9lb8nmbrgb/dLHIKsQ7tUtpFGKRy/8wQ4Yq4MMP4AIShUjVHxI4Cd1vsY
N8kQZkzVsCR51iioFoGU2fpW/Bld4029CDpAQVM3blDWaSFs32yZV9beCt1BO38QOHYvhEMaL+sY
xx5wY6uDgILE8yar5SvtzVrreigjASzMW/T9KUUGrfyQVhz1SXGl2bPwRJof+ycbPmhgJBP5i6uF
lMpND4Zv3J+Ky/YOHAVEICEJneH39l/TTfcSLhTS2erJo0tO58Fl4a8ifG5E0iX6A18Xw6KpEoRX
NQYkW30qC2xRK1MqdgEboP/HZgHwQwCRR0euSQML+47q90hyYHr0gDsHq568EMKvm3PnKA++7Gqq
mzgtn2lE82QvDVodR6rs1f892piErqYlNGpanq566JYg+RmbUsnizEBJMK5jWfqdZS55jecgD7gH
zomG1qH/KIWx1vwBgQbwClsdDXZyikc0FCBZ0a698bmhnNLtCUozvV/rQO4iez1gLA3jbTzgmUH5
yq5iBclNFpBbF4XhF2g8bNnVtPyJOO7VMkV8/KLd+bPc/YyxqA1qwzkNdA1lHGs/aWrRzKK0ZUwt
y1xbQgUnk3bJkS/vTfIVoL4Xrrr484M7yEnYq5UbG9Dedo2+YwBOhbqXkrcnSiwrw6kgvmRDoQwN
aLFk8vnSNjZ0a4ZiCLTpr2PNVtYnFHBWFwqeml8SwtuShEnGFEJN0TdI3UhkGOtcHeUxzjl7m5Fi
rcyLb3xI006cv4lxyM9LzwbIbmnwgttRuJx8kwyrcO3hXACzlQtTX7BCfDQWOF7XvxpY1N7ZDJJ+
4Z1jWMIxWPEw2PwIKwVZcpRH3IKEL1HpfOWhX9b7RPgIdnFMiKGLPFxP2UR1w6CRNajEEvyI8g7S
EQNjNexUNl0H/kaWPNSOFaB1qtoRmLBM6Yj62IAmNBbArrSnrLA5mfxoA9oy4viXqccQEFC+41Bk
8KKafjPlSePK1MCFMxhuSZxEepC1yPTVfK/sqiIoTbOwr0lLmYI9Dk9AJWIiyJHrUvhsgYueYhvm
9rptOlziVje+1hJyGnFhiIh+e7sUKQSTQ5m+UR06V88iKGeCnEWhOKgy8vkOzROimtMhEAv7wL5+
crZFLpNJ9pj5KPkFxu07CMxEWSWJzGEtoz/z+yXBaAEuzlLx83gy2It2Mlgfa8PugX3AlNRX33wW
mq98Km0NROjvM5sxk4pklsDDRDoqI3oYFXCfjMmYY7MULsTGuTsnjZZs/qxWCNXlaL3/6rvpa/sT
sZMVSCOuoKCZEOrEMyhsYGpwcry/a6OZwz2EFJKFsJlIVjlwPgif2vLoBPOuuYnMFIzwSFLEphuH
tem0xI96g93T5+SjmdOKR006uakvoOloyV5Ys2a60a7zVihUVtnqRZXoUC69ci0BN5P4l9BLFU4Z
C/PCJdsQofUwrTgR4A7ZD9zpLVQton8GbII3/wvmsWocexlHl+X34TW1J1TklZRMmXVKodIR68Tc
U49v9HHnudocfnx9JenDmMwxRkNbyzeDsdGn5XeHCBqKftBS0XwD49yXmZ/mJnwYvHxX1pRAAhQ2
iT3gohLEtcM+qgpwOQNnsCQYNGIiMXxS9cFfwMlsfJfgLBs+/v954ASbp1YYWcWKYLLM+Yt0AkTa
XB/gbHwCmLgseGOR7qmrwFTLWgXat10AEOSbIqxzYhOI3qN2QjQyhaTJ5OhMMlzvpH1uOCMhfZu0
ywJx4JViRtzE3hrtPVFmO2y43vVo4CAW8JrE8M7UgLKZ7/XyVn7qwUJcKeBQS63aeK5QR9c+7Sby
ky89rXuIiTmqBqRCqvc2J7s1TDScOHP6MXMPJ76IgmY86j83zcCwFxo8Zft1UdIUCUgxUPYtsBFS
NmEUuXrMYK2xB4z5HEsWjTeegoE9fcflIxGzXdeY4p7MUaTlHZ2Q+X64trPwizTNYlpLk5yiUX3Y
WJoY6Z3swKAKuZXTqk8d4kVq1rqq0F9krdBlFnOEiVyxF2TFokAm0dG0d30ibwgmsbyiVrbu2jjS
uBR4GC/5PqUygG+nIEcubGJFPqaH3srJtg6lXgUfb6BR5q3CkDS8BtRJdyco/9YmOpaaZW+agpaW
TOBZLlshMd441Dix7eB7qy96rHaMeauJDw9E8umMOwSglGiHrw4K108CZl3XwglOYv2qJhyHkUyQ
uAyruWnMrRM8NbTr2sV9ai/BwdNIMY+qCyk6atjT7sHydGj+bCefNg5xdxj611tTrVy5cwrxERG6
/FjPryxYG9tewpDiKiqV0k+BFuX5/7YP547w7shfSkHApJFQYE/BUMe5bevJj6ccnnTy7yXCWylE
7hGPlHd+pJzMq7MxC3EMkzC84U7tHwlPTnUdLmPM0oJDdFkR1WJBeqxYOyfj/UsDMDvR1QijuOVi
q+X6Pm1h7Ak6wQ9NRp/H6pI4TbImIsIyXyjGzlXbq9jVmkJiFizF7b5J0BZO3ettSrHcGVTGGTG3
0K/OKu9tP6aN0iU5L5yNYfsBrkPwSDBphEVBgmtm7shE/HvouzCSeEDLaDm3YFJ4i0BJ2AnHjD0J
vzIuFYSu6XlJmtsI3xjzD3m16owkJbXPv2PHBXCsq5xj6hymTRDR2WIvj6NfSNhEqi1FSXEDruTz
wIMwPmiOA8riY2d5AVYPjc8C36Q+svgEJjfzp8hhEpKBOSsF8xuekjZlgAWoQM+juQDiF+aNngPB
MZ1IOUntKSR883iyhOxUvBHWyo6CbBOlLi2Vh5oSKaWNrJJCIRjGdOe09P6T09NIbw2JLtVAn/gc
MvMfqtWUsGTc/JBn9m+Yb2wiAu2bBPXtKKMERCDI29tECQwi+5OtFm1oGdexL/Elw62gXphieBqJ
NkfKCPD5SoFPUkkL6j9H21arK3PErRsvOk+kwk4ptEXdvxVx5PhIYUCpfVDJFJvaov/KGEmhDGw3
gRsYRZAZjxph9d55o/WKy0qZOP6ztDrCkX/4UacTzl4MwLDHP4zOEyV7NPaXqbfAANEMlUO4OVMp
Ez1+0dMx3tEQoPzbJd8oWHUSLfAYp7xWMbQ2sXUMJbf6us+y6gseaXiv+5nh7GJv3yFcv3oc+eaN
6a2GDO20wl5pNCWiwBppfIKkR+tWlqHrm8cJbzpnDIScUgWbONdJ4poidrFduFfyfZjOeAxJiK/P
tGMilYbHlScqY1AHgbHykWnKlT2z9Nim9Ryvt3dagEBwyGEQ3FpoD5TURW/afm+SWhHG0cVtYgRB
DEjLq1YdVF+hac2SZvc2FZ/4EYTV0eKADG/Hzaw3BkrabU2HZyxGLUnt2X7VWGT+GM6b70Jy5jcg
j2zrvM4UPgfBL4Jra9p+Ixx4k92qvvynd9qS8tWq6qLL9g3rDAmzJ3xpRn9f4to5AFjnf8xfCoo7
kh4GuZELMtMxJFFxt4lJgd0jwouay6pi34OGAQTugNpg/JtMFJnz6lV2rvK4Pk6UOawvU/8znDHQ
bR8duHdMm0h8vJUMBFRuPK3o/JMjEq49dq3DSOWmTvcChMH7TK7/Oxizu18FQ7rXkWgQmZ5aQ1q4
crghIzs3Ao7OQOJictRNkW9XMwJcgTInvD1WxyH+ODmUmZb2mD7WB4cRJ2UfrqLrOLni7vzInFhs
e6zywOViw2JP2sKxq45pZqbWO4BGsod/AIfAedIO0CWI7pNXg0QAnmFLiTGVUbHLZJQiZLveH1bg
ZRp9t+7FZeFC3nUIbRD7v26hg+aX3SCoa0l4+sRH8AlOPJQjqtG/g5ynNVi9qxFeKXaLDGyLszqE
yMy2H47eNwyZ7yu1+tfYOWzAK8+zP0yGUyGH37H5M1TDh1bnwfenfGNrgzQ1p9h2vmLntNIkEo7B
XBqCVzr3nHDn78IBFerzR+ayeA0tnejumcMTcbFbMIFYeCj4p9/Hxybgeamag6liMDtdHLw1T7N3
8Bgfs/790BPjMMpakRmSN0EP0fdPkmO3wkM0YJ5aLlx29u0ktVzpyLQBjiWVwaRIY0nH5qCYVt7X
S4u1N8tfTS2vb23AxurDqAiDl9zzid/29kiyCaolwI1osIQYt0zZWlC09ZFZYutfZAOkTvDprG7/
0tknzzlU/ySg5MYjZA1fxobBQJUb3T3bNX7V3/EzlJBjLT/3si1oeCL+vo/xZoOeTu/izrY6uS/H
7JlrGVU3SC0mbzJ8UiGIAjzHiIvYh7uRVn7XEabzRJZxEm89NPxj9H7OC5VOjxemaMr9Oyq0pobe
P+aaGEU+7mXgu4saoMm4i78+yY3QAORQWQDPrzEe2BeCUveaj7LaN8VWYFPLblF+aErF4LHiX9Ql
v822f8hBWBf77xy3u/OgWPrZaWApfO1czejYe0eMuPGdLs73P5O72h6PhqVvWFJ6Z2cugVo6YZH/
Mp9GRKNgKv72NH4yhAHjObz5YHKgepIAP//wza/Dok6NdzghUv53L9UB1DTZZMwy0dXz0oUaJ7FM
KspkRfC7eDWKcdZHtH+vOsvz3PcKaNvyGm7HaF609OZJiicJY7KB8D4GlMayo3mNZ1KafBIdwu80
YQjng7DKzH7xdfAmuF+OF+mgM/OvKyLrjA05bxw/Bknyv/D5Kp51mM+T9eAQGLn7wuxH+TfConIn
6Rse9CAqgrXGjHGjc2fRS9qXiXyjKOnzw1rz3RM34ZXHVrw/+XMVN9CAXDXGTMc8I2OhaIz5HdDZ
ecAYXKU7vxM6rCxhjvJO8mBNIT0rNmzIEs8sTl2SfCQCwCaK7Zf3xRlSKPJZbGf3jWqfkB/bP+F+
/1jXspQN4xQNoQF4K5UWPdQL28GVYVj6Elr8F/ya+q1ObmlBaXgU4DL9YPAnBn4VsiiFHtq97vYZ
pgJquJsl8dBAP5ukUBVfrRENweR1nq+OyuE7cxGWK/61FXRIyT2X9cwhcgRj6WTA3Q5BLIlhWkY6
6Apc4B5W3SXT1qkctiAoKSxjYkxZRHvfehMuUtHbsfBDGFVs+ktOt+SxwpJg9cxMT0uT+1VUa47b
cfNSAw+GFRyiMrTPgtbj2DaRIpAN0cF/TdoOSneV7hqPzU8UGGKTt2/GwD1DBOqWMug6KKCJ9DQs
otlEsJr08tvYhR6Xv9qoWOPmr25vguFC6Q2rFdxJdx3Z4h6yMo2wa8DYtJMWMcCg7cqe1WFrRB7A
6wIOxC13USGqMrShyY1EOzNwB17V9M6LlLX5W3n9IRaqqLNb0RYv/0Y97iIz7OEjQQxH903Wr4Sv
mepsVvT9b5+VfMQMFEwxOzyMY2LoP+fF7+RcFjGQsm7I1EceYyi9X6+k2mO+4R/gmX70tt7p7XlD
Gp+u9V/viKdXMPbC3srv64ueLyHNIQoHCcHXwGlqDzBQHKRCvWG8u4cmen8WO0U2LbBaATddPkO3
wiv5wGF+k8/5LImb7dvMuRwlZ4sD4mfB1qt8bptgCpOQ7X5WwRicuRrKqoE4YsfT/AaJtdquGKtT
PckkOLjcszkRgMA/qUSim36owu7JGQxuWFporLGZEJf3G4d3a1INeh94ptRM1OXGcvqGfnLhvT5U
xVIVSNpNi8gmc+03ku9z5VkClzlIMIT1O5jJBOzB59StpGlYWaqTGKPsCqdxxW+Wl8YWkoGJI9ib
H1QGLUbccQDuAAkTKrLbQL59hUhAgL6hGB6cm398JCX3FxoD9pbkkNaL+TKjVAk6a9m3XHKpmJIx
yzII4GcUMpNMYxIcOZUYzUm4wDuo9H0IP+rZBs81mbbqQNYYzPL9hw4QegJY+SdNp4oVJJSUvFDA
sctKDcouACQiM0wwge9R8Cjy7u/nolvFAVQeRtTsYLwJBZ5HyvPNCyM8zJ4aPIXOoFrA9RHoGPO+
kY4TOG/sw798NUSbvnPfYZv+zmJCUuujEwXFN03cJG89lUtK/5hdl24fSFqd+Yuv8r5YfHxNn4cS
5VAlsKEuLZhxpNhIjTrJWLp/cyxxsN10sFM9O9ysnkU2DiV58Dvjb1KoiKft3QewFPwqYjj2bIuz
kRhcnZrgOphSQAkdqMixVypSPAcnD+FsJX0bctD6mTXM6rQENQSn3FQ/3De4Vu3H6/v736vlYndo
tSVRsQ5LzRBF3psiXHdEgFl8Z6S2wctYp44Bohfxw4Qg4VbaRv1FmJbxR2lcfkW+FOUkEPGY6wMP
2wFHYz4WsI/zdez5NM91JRsP1+fgQ95lUwt46Fm7dgy/HD00rOF0bmF792aBZnwZLaMzsLu3NYhw
4665DO7OS0CxONHlJ4wuThxvtfa/yLy77/VG1c8LDLVm6hGg/EbVuY1PZnBvMVJBEAaZHZ5HLsJl
fe0d0RC4/3r9vnTTtns2cTmOB6v/k+kv2LFVC25sEMcZ88F8wseOLtSoVySMbBxfs+6mhnofIDtN
TtbOYruP3xKVCpNwqN5EH71Jy98ep5G4EfFY5RXsYoLMzg5ypdY5IJEpucTaqx+yHvVx3ySuYbKC
xHEcDhZioryIMCfu7H0EXioo2Mwjry96GPzC37flBhXsFcVgLiKsMv6pNNAfPrBN4XKXDxLhDJr1
8epYaF4qQFKsjiZ9vdBL45SGYzLPUffMp1OKauBxVh69hZBSkAS7eQL1CP9TcCI4CzWgPhwKFLjH
smUmAwXLgL4O41IYcUw06X3uCOwH4H61xqFtMRm1DDEf9vZgOOXwaUPhCnfdudfvzKGvImAiGXuH
syv4edhhOUsn2McAtRjTmi4FB8pR9u3dSY1TTVODxpSv60eHpSgJtidCEoR4EK3Bwt2aYe3I6lOm
fHC3phMFRx/WeBm58amsS/4gZFonwzdKKwnlboeejX+ztteMQ1kzO+M4jfByyAKFzTNQF2wVrB31
Su/YHStpv0uPpJG7hLzMQ6zGA+LyxXfELhVROQE7RUsbGUHlvBHuR4x6BkJU4g9UFBeCs5Xz4AZI
o/eUBLnbUK6PMi4/1ej5ja8f75qpk4TLj8KCVRJ7vzzfIPF+AhVqqtDc1z1+XVI5BMbVPwYAEkd/
DQAxaWfxu3kBOt/cRjole8G0TKcA/1Qdy/qce8aPpnWdvmp/hkkk4h6BdB+XpjrgP6jLhfEOAwT7
kmozqHAQluUo3Z2f6UQzflVsdc4iCx6JGMPn87cRAKTrWWUVqsd7ZXrjRzzvuat+nVVB4H130ZKT
+E4Ak3ff6ZkXRyuXlli1e8ShZOp1Uprhvc4YbqORCwDb6HpecsVWqAcdfrkL12FWefmlIbjG+P2e
KgeLHHEUCI0SChITQ3salLV+vZY6L9T8PdnjkrdJY2uGCv6B8Q8fwcm/s8VcUsAPXxAKpaIfpXhl
fNdoc2meDB80ss/BX8mrPjyI+4Da4brt3bj00eHDwdy0MBDFolOoXFYUIzw37KzUeLuxx2n7P369
TAj54jVLK8lAQiu0i4jVjS3xgvA11VyqRt7nlba+/rfJQhUwW8vCz1L7tYjjYTQn2/PPHPRQxgsi
LV0kC/oLJHtrFETnS9R1Zs5mXjc5rIcjJ331FQD2Z7unCe3INUPDOhweQfVAAzkASEzQa5ojQZNN
9YeGS+bYIFS6m7GYW38MOQT8/EJoW9UHByo1VzpoUM6/v8DgL3qz2oHVtfn7Le61cOjP5d3pdiBe
90vQDTcjoospiY3bY6eChgFLzjO9vrEwuyFgGTKRblxg2SNsBaAA4SXb/0tmCcmXmx6ff2+LHyhe
dNN0ABezMUlSCKA8y/prq8m3NWI/C0BhJL5Hj9gAX2Nnw8Dyg0/mXRFm8VMg/mQEzQuUdXeregv1
Mo7+66LIRjxoA5laAj6EpSdmYE2grVyeAiIj1A9t6QzizoAlgYeEZFGMPdohYeR9mzRHbf0pCH02
/8vq0GeZ8JpbiGUSL8HEfBusW7vGiguSXOrmz9Kz/5ulNm4rt2nt7/2cAs3AVTO0Do1rpbcoUfYj
4kYWslJGfMIDqBdxnewa2BKu9gNDslbMftu0wbX9ElEu7tqko6564ZZRenGbY0tvveVYIGD6HZ2q
XANgrOSLe6FbaXGXH0YZK9SzNAX+TaIGusF38fNZTli8c5BWYo9RE/gILil8Wli6CEENlFkhadSp
pw1bbGoXLT1o3L/vHuhKj4KlAxEZN9TVM64r7nZzArQOWerZS0jHYeoIALvFiNBthKaf3Wmyx6Yq
mAtuLLy0PFp0KU2Xu8IlyB6oH6IL41IIvIqDK2aUzfj40jIIg7cvp79HY9LbANbuebAG9kiMZEyf
pyMtqjN/HROTdWhpDRz/i6+71Uq3Fjfn5ese0hqst94yQa73Nl9Gr5iI8YAP7M/jqYpUnklQ9VJm
rekFl0ur3pv4gFoudgXBQ1bDyVpW4IBBT74sQIAfdrhbbqo1N+HJaxv1eo+6wua4FUtOqnlPiUqc
ilYIl4t3p1BryKYQkakKpgSVB6z8IV8UvMN3VHfkUgMCh7YW5dDnRpH0PPW6q/arJF4aRjjX5IVS
YpmuVBlhYHUw40bOMvYuKr7s7Fwaxmj9ywoDeNJbsxuzJ70e4XxXG+CXvYf3moNtdfdfEbNFb5Ye
iTLU0E9hxCz5y0RwKh1C0r6PMnsB5oJ/6zVvk1fz8yDatJpjLhfUpSoJvrN4InqMUwe2A+evNJx3
HJiPbBBIzfhEn/cLTGNQVmkzbNfxiqLD3VH8qL8LJ8Mis3n4SCiStcrHgJjicyQ8Q/36AWL5lZzk
Jt87XBRX6Mi6XzNB+hdg4DMMpEDLVos53VHGX9b34D9SY+lUnSjw0x+F7riZPU7rUphRLuau3lzy
h7ze/eSbVvdjb1GrVVDgFk6hTKmWU0i6wjKineJ+2k1+9sDqZezw1d4n7ejhxABFW5sd0jVJJKA2
EfAnknStpOXJWxtmgmSoRIZTUfTvWvb4rkaY2Unxfu+2LyTSlu8GDhwKIBuOKwzW7tmC3ErztovJ
xbVRIJguvYFvCwvm55D4K4pbvE2nskl6uKws5ZTbVeRIl/gPhRxOyPXdBD0v+F91mMfTL0MTrfFl
WEpr2ghCt//KZtSfU5PLgXJHYel+ppEqjADHW+/uuownfgp5iGXSRLdcLyxgajevZT+W8UCZ03wR
d6ikxNH4ZGivtqBVKTfmjU/QBIfltIlUa9sOx6xoe7D1qhz1lCWyZvdc9mqnXnKeZFMz+TgHuQiQ
65nB42wD+5iIpsXV6i6lqYyV+42M2QlxVM0gFWUoWGbmGlrGUVMDaSQfg04vYgHXxftw+GKGM2jv
TkbvNOZW2OSKjM5t//IA+8UkUW4tBY3NSeVVusOow6TqZP5+WhAFhFX7DJDMGcIfhn3dA/djB8G2
gabrQNpgQ/rtkzxquHKSLY15ngXgnGcgxCFSxG/3T/CHz2nl2iSxyU4xlrfNwJZC3VrQHBxUMgEO
FbCmnUrI2wKBAuZQyvltixXTSwGKzXD2IshMxlS5cvpNL1VtvIz43Sj1T7p3bog3N5WG9IoRPgE6
0+O1dfqVcPeRODCNPAGAho2VdEWOziu3UMkaqlZQoBl3USJCU1eoKVnVNfgZ+SUPuAIuLmgMD9NC
gR3XRZ2+uGr9fTig1V9cQkEn7CWm9q3qF5qHmi+IR4tKPVzNQnePBpyge25Y2bNf+2mnZgUZTc02
N/AlrQFI3TvUAXhC6zF7R9dDkJUZRdgVdt3J1tYOr0ZmjewLy6LftRcpYW4m7SKtYOF8x3WlzEkS
Epcthup1DN8G3yDRu9FjfMwfYtwMs07qBbywnDirBl9d9Hmm5AxFqqA2+YZD3qLYtdF2u46vL2Ad
hFopF6X7hVKbBT4x7jPKRVAOp8rmcNJNVZvDZ9GiN3dqV1U7rH+CTYz+U+98sTudwDhXdlDGlXNo
MMZi5a57jsT81+ShtuJSm7RnS6VmPOV7YmQt/gWI0mCbwfkfD0rp8psWFXIJukNIfLaB7lQSqRQn
sQ9GTrkbB7b3JhtYjJtbpY0bGfPzSCjBme6emfhhS4gM5qK+DCT8hfW+p8n9mr+3nosZ9IWrdmx7
RsG+pQw4IGKXh26SxqDnWAK5n/0/Yn8eNLKA0ZgJPjWqH87qvYO8vjdXHv3R8BR5F3X4+GLIr2VZ
vJriP/2kBqVPC/teC255dzMdZBb8UTe+hVRkCXRJOzZhqvooT9R5KVv1TDBADwxbx2HoxHW+rFZB
eSm6KSxAGrAPjjPv2gR59b8Z01mvAJmKdyKKmuXaAOr3xlCEmdaiSQ7kBBE7Z4tCe5UxNm37Gyhm
G78wTyWHj7GT/7bm4m1ej9ClB+b9UVomn0cDhBATqaW2fKF+6zC4+p36Kpyq6SaeyQ6LcyY71WRp
P0ZmX1u/mVywVuQoS3Ppy5Ro6VXKApVDomI1pBhFM2SaB3WxTDoZli3KoB+n5Wwh5URVU+DBAqcr
5dhOGTlaZXq/5iqg9Td+ygjNjVDv1MK3qZbn8TTZl3g+WpEnzjfY0tcGxGO9ibyYE7TYWBxAUL0A
SIQQe+eo0xGNVM00rd6eSV/b5He+xrFGbv+Xgs6l9Yti7FQL9vcmHQzD4QzhVj5wddNyzeZ29l7E
VTaPfjSrbN2glpKA1zciPG7lDOuDGBbv4p9zA5xMpgiiaCV2VHhJsHTTbDb8xr9NdNDQq1HK2RtQ
rB2NNogsPig+ESRhcdsITBHfWEFGPuB44SWp2G/CytqND5fsep9U4OyBpP5LoDclYT8h/D+VpMu1
TPnAObPuBpVuBEprt6rm9k7mNUhUWHkA52ZqnlvFn1IWF4ZXgd7PMr3eyMZGs8OCBUi/8NHMNBg8
sKAvNskyZh0gYDpbrN+NUDE2U+IikwaemvK/uJ0C/617wNQojykhvh0OroxTLO7//zc93nAnwGct
g+JWf5E4L47+rHtDHYmu3CQrw7dG5hEsU7wXJD7l8/nYDz3ve+w5Mli4OJW2O+7z3RFpz0hp0OU2
znnU7f1NJWYofshjfyhdaP3tnp6jrAKOUsYoucCt0mGGK0NwKq2lvUh9NLURA9cx74uMN9tuM+Ee
N7b+HWIASBex8LuVodna/SdC5Xg4PGOolmyHWSPoCaJEOsvyE2hHWTaOS/nTu9uX6zzOI/M+fysL
ffP55mM3bc64YtRQEQIf2I1bE0i/su5gulG3B86Sl+RyoC4q7DsNyl3v/15meDQp4SlX9jP0gEPM
t+DewNoxKHK2Ci27lczsYi6+yi/UkigURwnN1cRPPfZTUSQu139h7oqUH6JF7hpIZFWn8kpeIjtt
JgEAHy5Fumg6X3kIwWILRPEZvaUQKJ3UVUDadwi5XGPdEQLZulea3yP4WbpINtTmSJaPqHoDAHEj
BoITlPgaVl7epW/rL7xBEYIS9gd1FL22UJBfeh47xPiQv4vEI30pgwLoh8MNksWFZS6wZ7svHlEl
MqD2DZqvHBJS3nRjl6GBi4RdSjQD/3QD+tLsaUoNJwJedS78G/46dHR5z6xZ0umGHgO6dpkDPJao
vd0TTkpCUEN56bdt+fT/OgQdcSxl3a/TuKikV/ig//MdjgPxhIkc4KGIwZ1pC7/3k+f+CR98Xxh4
+drvBgrec+tMi9elAWRLdjRnkQfVQAePa/tAFBfbpMNt+RyLiDyyxbWP0eCpcPFp5vNiQIZgRkBW
i1OSZxR7vp1+Wwgf2RJQV8Xcb8iGe6QSf6cxBniqCBWmuS8w2ACBEBDRgTesQTi598XQEwRkjUoV
e8SDe4kfNVJ9kqX7QQXyUpRISH5ihrR5BJt7mVdah/O9nYukVBwsz806wXS0RJL9U3uvqYSd1H/n
iK5wX3Or8drOXJ+shnS3nLple7f0MGnkUw31S9GJAazlJrBkziu9H5AAFA60F8dsZ2ujKOkriTE6
6NECv5z25FcCu8AsMN94Pydcz5QW2I4apJjWW9W669x/xS0lkY/EFYaEuQiYHLA8/wlu8xI3LyUf
p+dMt9HbAQljK/PmprpbiXavXZSewEs1m3Bz3ri37lQS6iyrc4QSBH1JfDhrhqab607FnglSIdp5
CGVE43nYb9ExLb5HhiHl81x7QQaC6XEjkbh+1oQrVtWzIN4GaRzMZ4jjLG2fx4tv6kdZ2Le60VwR
2Dumm+5VflWaE4M0Mwazf4oE+yIdIyIYlni8sy1rCQ2HtUuIBJXTmsXIUUVpZejmk1w6dbuc8xPm
y6u5EPwaXFfsQGx7FJZDMqFp5z5Rm4xA5dU+/GRA/uOagk5MmIUsTfL9+ySbH48DDhRoy1bXrkyO
v4i/vu4sCer24f+v3ETQ2kKXqOpmyIqb8EHjis0Kk0dUj3npW416SdmJW8jZQd6+LbwEci6B4ckc
/6mIRG6ykyIRfZonP2blB7pK0uoulFNw9wd22h07unabTK/g8PUi11vR2ODVGoAHcwUOgVJjDvF8
AxDDiBLjIVogIT+f8i3RlYdXszsUhd3L3CHkuNl1tU3dprwyNYOvhLT3wsrp5+LHA/XToLvVPM64
7MO97YJXjPEezOQx2Ka1m1qM/3I/FFRHT9AyWR90pHG41OCEWB7EbApxL1B6IlVLMGKhsqxgA/uo
N+EyZGys+md9BumNwfhFR/c7uSihMpvyNu4jySQEcMQMTbAgb9BD4LRtW4TSBjpQNyAts0ojZQEm
ErfVW7fcj7OiB8QyjgDWH85C6+PvcCQAqWIlAStv9Eeg66QWDq1123Cc93h9KZxrIS73Y4poodWn
05pbZ3fPXcnhW65+yL3vH5EUyKOP/ffKRQSGrVZrpfuZrspJVztzYfcsVuVxQsi+7Vp5GoO113Ic
t5NEkXtAfIeTlB7zTnbP451be8wxskv5bwoh2YrAkLOEn3kmd2nVEpehzrM8emqqC4Vb4AQUEmyW
ebvuhsUWPTsOJEPo0IDzSYyexcISpJ3XbR356zGGIFAG71S3NfE8IkhzivPr0gKiFIVI0f3bEzVe
b4u0P4hrK3lmG/jC/TvZteW4SqY/jsSejRI/C1XiLXuPiFQreWcdNSV0OtvD7CUcmwIUR8LmYb+l
nUwQsbBurRmg/fYxI3v/DYGkfezeye27NaGN0YUBM26VSMJutHk2mR6iaUuurA9kmQb2agBdOjY7
A6oeNPmu/D6n7wCP30JbfjG4QyvnTb53mNP2FjkoMtSXpyxxK/aw+zdGvTTlxd8iRLhd/izaT93D
2asvNxhZNl/6sw+X+zQqnBkJwcPVeh3tgNOYa9d+h847Z7dodySIhBvsWJG/zkARSS8WF5XNfy7L
cEgIj2wSx8Kul60gd9FuvR7ob04uIFEKm9tESeaBAiZTZH5NaqRQKzUbXvfzO5EqC0eSZVMTF1Cj
QX21WRFuq2WndXC3Ro6LBpczNC7XJRh/sUs1jJEhm40npeJqTixeNYwNZiWZJkjED6onuxly7ymD
V58p97XNebD0L/K+CGIMlk9yQ5eKzT85eio7BfKABheT+i3iWLuj7eLKZRWgcyJXgW+XKGQJIUGb
2JJd9FVtTa/dAyKNzn00FWuy+EHiPxZSGCZ23sYvN9oTZRcmyBr8m5qxFtUqn2OeeUCwLb7GGE/g
NV6Ix7jb86OpMp2kvdx66/QYV0iQwPU2gITU01E7gvphUGnMyasDMnmhemNG2vgdqGM39VEJSQGh
WYsO4jKCkaDU5Iibkfnz66lPKl5xjVQpwAWYOcVVsYVgpurGhZqSDoR2AMI+TPQpS6nLhwgPECGe
N+mCC01o6skRh1zv7Y7C9MpzmuB2S5UjRXjayZWKk6xJ+ZRQOURzyzzVpNOk5W0k/sIPH0iBC6jr
vQ0ZzFgP78AlQO5AI8gfiiCxYx9shveRMFhNjYwSU3qiyrLnXUSFSmB/WKjGMvNHUg9B8RU5QrPc
qKcFEGPrJ1qoQmV4xnhinjaLeZiMj2AR8sX027fQiWTHQ/IGmhn34vcn0FP64z/XLvZUVuo4EL5b
xaJdaxzJY8AegZ8X0tludh7BJNeYCiFuGPsgwkZm+XjipFRSssCy6ALCNXAWFEedrACB9AS7yQTX
3Oikn3GOnTn07HUv6bj/yA23LLWOc1N93752piMrO0SnSc6fQBpPUGBSzE0DCWod4Z/Cvqmv8GAD
rJ9JCdu5nDMeNxK22IDHR9MyOCsxQJFU3Im9Z3wb6Zve8Yiup/ka2qFi7YKumR6GUz5ncytUzjPa
67o5Pxuk45kj9ABnguMtoSK50EK+FVM1WUyt4QcQS9Fc+qWaAIv9O0o4bPEJRqexCc7g1lm79+8F
x1/j6wv82Qw35yuFZN7qEhJLzRQmiF15LlVRn99N3cAE2C/ScedKt7RR+QJhJu54lnu5gAiePjeN
DNPa71Tuao4d4OEesNkBWYqljFcektbyUjz16LF4cigOsBHQK1RG1zejW8WcgJ/FBW0vp4++U4Hz
Rs1FiKFacF/5xgCy2Bts1mzgoagub89Y2tFH/Nsk3r+PAtHBjwWutfmknvrPNmIsQHZ2UmRERAvl
g+HpXrOqNgRB2AKcaVSQGgHRGB4EiTLZRa/mwD7krNLqqktxYtClt4x/vhf1QX7CFeMVzxnImC+W
DiUaqTE38wQx8TaMslNz1y+3SQ6y2AiBnojQq9Bo800TbCnAl2/TboGLvBK0EsF8VpIvYxIBwI0A
XXH7I1NXxPkGtt/Z/ABJM4rXrScNMlQEPAZ9guE9RmqLoFlDT5O1srLH1WkF51ZmrZh76z22wN3p
4T/ATINJMwwpl/FrpQhGyAJncaxltDv4VSvVIj0Cnu9ixBiSyh50PHkCuplTwowEvbZsYi4UV8gl
cOvHxq5lQx/HPPSFE0ddz0nCGx/hyBvg5t9WZ10RKsoeKxV53n7Q86Tw7sHHoIswe1HAflcG5EAw
bXv7xA/lmhJ6/isNjZpibnEsw7ZR13O/Hzblx0C0ul40+853G7eh9ecKa0YWv1hGhVLZkGbnHJyr
oIW3qXIF7jBftVU+NvRR1zo5Stm2cMwuPpt3MqB9AsI7Bs9QlEJR08FqL5tOqIq42tEQHW7sQvbJ
R3RQ4KiRypxzdyGZtwRiyDnnxYV56sGP4thrvtS4YFyJsor73H5i1Mq/4TKh81KBkHAo1BuZ76lc
+fPsvj+p3iXBG9Qd5iGvvZFwWIay/zqAk8pj2Xa+0a4xmOHgEwT7vVAZ82KPhfEQPlGdG+fy/hci
tW64DKUA8CthKnJhwUPhLp5ZUn+Qrr1w/JTgMOZr9Yfozy8u5scfC+ULmFe6Zkb+kOGd8g62uFLv
dnReDkuG2jOY5gZMnYDlZdA9HtBvL8Z49/VWeYYVl/dyMKHAQTDbqRHKc0qUcR6B2GoPf5Jjg+gg
6OsKmkZvNCjVnFJkmOvTOQJKg/jr/s2zrsY0qojE4kl5kU93meGxM6JGQBljJPgBHCWrZn2X1ARl
mp2TfcbNMI5QI5M07l14CbssJeTTlhY8UPBYck2Z+2746TKrW1qomVabHntIOtqY1/goY/abOPUe
qaI+SkiCsOON+7Ldk0u4Kktfu652AwMQmJkjxd+22a0NFnOtn/r/p2bNlEvokHwmNy9JLpVyqBBu
1ChQObrnhcGn7Y5ufKqYSXdqBNQ4hdvDMZ75iI020gs8fcrKypWX8JXusRwL+AstnKSQ2IIupcg6
U3/zr8Eg4HQ2l8K65b2w01QjG+cFAkPmg15so1IpNGDaB9MtrZaOlt+OfdHXdX8YKn6C74oTV5vG
2ucmQKyF/E/kOCRiz8YQLB1wFU/e9Xb1zXL3Nd05k4mnfWTYXgCnN+HckHqr69kZFYXaPMhjvLTB
a32UX+AWAElvTuCKE8R3CU7ab35KcgAHDhM7hDZrNQX7MxcajaRiyyUB8yv78ZzPil/TyYIS8Iej
R55fiM3nx7MHeh8B+n7skCeKwtupphhxsxslqW+dCk9uf3RqpCs/ANgRfOc8EEmkAkIpdumvYlQH
X+IRfc2PSyJ2daT6sTdqsbH1tIEZog3rS8S0v+Yg/u/1Jdv9uaRIFqWJHJpvVMdQAfyjhxIRC6H9
HjCxkkTnRUJ7apn1N0JwACdF9Cj8gLG9FziTEd1YJsAjqAUoIdhUF0gNjsQlirezKb0ww2/iYVxz
MQvJLNmICedfxsEx/K6sI7CS8qhpDX0WwM7C0rzsD7Kot41Du0f7gBeGRmYZ2Val6AHQ29dqndHv
euLf8pgezfFY3Zp3YLL2GTLT65VqmUjtMHlZr2U+SfALFyezg/K5nlvMVx7NLdfXbl/iRKs9jvA0
hiklrUb23TG+YNjJ9Zr485OxNBIrvJ/HQpf0r779Zg/Q8Z1m9ML1cImay5hkyNDrTWUI2rJAoTZy
czo8u5JQGWNgJCthVGbgxQ+u1at6WqmKa7wiwvJm0j/kRZrh20c5GR7O4Q4MyPdTHWjPkzwBFnr7
bHg4gbeFbDQlhiJVeWLHgzm0vbYeOQtO5/dcikJZG6IgiIaD1UrKkerOe2SaAl8ke6HKWUxMbKNh
XqOk/IAE6vitez1RJIfHZrMQw9bgB2kTEYKiXy2iiKpsXvRr8Ok9gvg5nQnRvvCpIJWtcQleo9N1
IkEqr5kVY1PkG618nFf9pIfkt4rT+Lr9nQczz1GhXqkSytg9Jsj6lLMiGDgiG3YRZ6vB2oVYsqly
H7oYWBahdFcn+6K/5+Oj6VoyQ8nTmp2HlcyulvJIIJrqQ4j8DGCwzXanjAMvTolAwXk8de4cMLsr
tSTPID+SfAFtJBKXYMtGr2Idds+Teja0opUhZGHkIEgwShmzqsAHqFRXjXnOw72wY2BdUZpSQ8fa
u9jZHZ3axoMHAIBCUYNhh9siyZTeKDhwUOB3i/VUzgOY7exjQHubMBqEM5KgmG56Ee9OW6BryK8W
w5l+8oROt3EHFSRzkzqk6wg2aGliPeeU2AMFb5QEpFrkIYPEwWKysdo6abILnnoAy6Xw90hqNuva
m1U/Iwywfbne7Dl/1Lr30+UXgCrmtXOHIROYsqjnJ6pCgDt9KHyhZmlSm3lpKihpTOLc19aUsgEC
mRPsF4J5Zid5IpaFqbIqDV7OnO1K6o82fdoRySVSb8EgGZntHjmMBj9jDQ9PJaWTo6qQ+jRifvbX
zhSr7mRXt+06GiKUsJEqipRGczkzPizUYaX48frztbCTV0XuVhl2g55VZfaFVxFY4EMxKD8txVyb
bd3xZjg7Whe3uMY1PVMZi7ZcEy2XiojG5RDWSnyKjntgy18F978gOqcptv0xPC04wRo/CN5NTpfQ
+lTwvC0I6Q8t4zdQlaUK9Uy6cAMniOGaPJUczx3NVYp7rkxRk2A0EtUgATtCS5MFwe92x5KHrx77
eaEMM5L5hL1/hisFQ5/OJynOYRAjlpowikPryZGsasbUanbW0Q+rMALHt9jPub0a4XJeq+3nxkkd
8Na7ELJczimG/3T0HZMoXw+03ll5kzXYzYpHD2ZEdlI+nUTfu4rtOmhAq6vcUZXBKNa0xsD3qe6K
+vHSxKIV/cX0pYsZdM4CSFbIJCLasi2iC0ILSaS9KrsMdFPmUI32Ajgzkmr7NNNB8GPab52HO1+r
r5p4Hbea9v2dLzA7H/OBIzfv+Eo7urBp//+bDjjnfIx9BonyvllrjOdGTBkOSyfK+1NP6qwLc7wo
bHzQRFDOXooDl7QBBf0QYCmxIAEWMTrSiWGeBxuX0lEeIhbm65Ru7ZJOgCoaP8RcmKvVpC6uPn5D
3z/scImAtq4TVWUOIZNL+VDrvLOdjmQM3EG4H/4bReRpPnkbNIJiXohIDWFmj4mCPh7T8mIowSE7
LJO/n24ePvoOM0OqGM6lOsrcsa1aiTqRERWAlhu60bQx8MkLlMGDl65Z9Py6YGfxwqijy9kEqGiS
meIkbd9vl8WAs+070CvSBda2CPRuPIrONHaiy0rLo/EJsyJYfeDqDdqH369XW8GE8weeajKcQtZ7
Srp4qZs5Cc7EZE9yfbWeoY9q1nUo6B6/IWnWUH+9zP7d0MSAQMMZgQK0cCJBA1vRslr32c9V8YVM
GXaeq5GL6piQKexSBEM2kLj9Q2RhxlASqh6a6bv6jBL56eXmwJYmpCIiNN7QOqF/Re7obomdd/Wc
UK0dg6po42CuXxZy3wOPOKsWkZOe0VnnhXf6LECK1N2jEjHX8c4KJr1B1/SlSvB49go6vz1EAsba
OA4ozkOhG4aW/IZ3Dh1m59g1ndgaBLuXhXQ6Y4tli+ltxOMGWOBJt/Hf07Mr+6H22xYV7FqULhxV
+FZnz8v7WqOX99uJ79axzn9lH6CbG6cefRbh+NToOOPKgrE6snk2JxoBFYE40KDOT+P6lxIFjRfY
ItJEuCRNYWNSeAvckkqiXd8fTBnmeYf7sGvjBo0QF2BBVq0wap6pNHPA57BSyMTJM3a8/t15Ocla
1vr6wwmhX7Ut+ZJmABTD1SYScAoWW0V5u9wwlPjxczOeRwKM37bY0HVqB06wRMOBP24s3TtHWYv9
YjXoO7+oX1UIUGc58t3flSWFybEs1KP5sAtCZsRy4hDcUmhPG/mQP74lQj3vlNLJ/EYw2R7XjbJr
g3vKoVE2nsDMtA5MWmX4AYnWr4O3KPzqrSpw+vpWVJpv4of2yrHHEOfYtOT6cOQVt0J8wWBjYkOZ
WQldOgpEFX90x4oPVRqsbzMNyDR2gPKbWj+pFb7dzt948Vca7Zk19EClxrtqVNIQLAsZmDANJFql
WFzMzlovro3oaGIVkC9dexEl/6lLSAIGFkxAWoUxKuCisEu8SzdqowNdNb/2c5kgnKOQM4nghDrg
VoE9KV5q2MgBsYZ54V1zp3hCVkJ90oQRiuLf+yuktKHsXKQ5J1iCyvyPQvIGfeO3paLarF7g/lh+
efygJUnriNzzCgLJRkpjQDkFm5HGLsQjmGBDZBq0eO0wzpzHONogX5UbD8lbTUIox2i9U2macxbB
kudwVvNlr1ZGL51UEKqAqyOW1Gz11xtnV5rzTevNH9l+AI/8ByJnRcEh1+SY0MMFRNFGpWeunwbs
syweFGtf9fZru2pRs/j0CBrNxTJ/1Z/sUrW9FRNFnXwC7cjdTnwAn3VhIic01/UU7ybq4T4TXrEr
Dc5PVwD42/TdVtqTReMtcRGvJSRWVaaJ3rA0cJf1aigffNrlqUrMHXukM999MF9s7ptpo9Rvmxun
DVUuwP/XbRoRpBtvi0iTEhEKKjY73aTlfVG5eCKUchQVecQkYLdPHwhy0PTmscMhYRPSjAjLHkbz
dh/TfM0iUMSvLV7BNuU9ZElycD0X3v/A/0zJvlgEo0Uty0kI7Nkpl+5PagfwecWWxaBnqtEs1C56
/kCSg1WaN1Vu34P5mQ+g0Rm7qXg2rbnDG3gTpzC8Ol+mo3LoW6diSG03ah7dIcuCMyS4iGDpU6K4
1TV4D03w0s0fYz41klNn/fAIIjDFey9IUMg4DU/gR4orrq+ArFPWmB0Ho9CwBdL8xGGZ0Ndgu4ne
vWxZ9iZMU0d50yyjZ4GStGivjuJp7xjYFLZk1FBjdByk4DGHO4BKg7SVowM0RjmFra58iu3mwFrB
NOVhFar8xsznXjmvpZaIQMgIVI4c/bKy3Yq6jp3NeS0/7Yq19LAXfzWAJvcB1dHGPYKKaNmDw0O/
uJbA0xA9TbKzPBwfeObnuBTUcfkz/kEtjKtH5HiDqM0ZZNqkr5D8AuLdrmdNq3hWPImvwxqP1oL8
mjJSnARZGQfjW3CpyneAjb94AUwuk4y6r1sheBWW1Kf2mFNSstfmAcett8uuKIaroYOq8IQ47ZCD
nUWOMndJVa7Sde7MRQS669FQwk/0lWQOecnCLMxA1UldEi+XMVOM/dSnsp+b8V5s+htk8Ppy4UWP
Uy6JyErJae/p0LABy1yp7oMseMak2umWre937GiQOiF8i/2pKr+G9H7myp8Vdl1UZffkOXodhcgD
GtebpFw+90DeHXR9Kn/VEOvm+z+OanSWeD7t0Vm403Dkq4qljettZBBK6jw2fmOhkA6LgCUga5lT
iFdv+XM+0TWnl03yNwnAkF3s4EB6pFkjcxJd7WSMV1iWC7Dgvh/q5qGwit6RCekZgedSOX7LZ745
Le1ZWaWF89Ae2FjoeI9FMfpgU6kIBZA5NYWuVQZ2SM3UQY+w2ep9F5K/Ugxx8YfHWTcX8JQwbueM
jwXAYJ6nsdNVbjnjsmQsOnTz8rUHGoZEkaw2XAX8kVxQ7/yoj5b9n94w6Q/U8eQULH3oURAORIO1
6fib+gKGp+17h3oxG4i8YVFoIxfNj0P+rZPSdu342avWQUo4LacVHXRov/YEdzC6mDkOOIjqtBow
sE1+IyujUpVarsQy3OnaXIzrbQf2RmS35gp7FksAaQFTthIPImbbHLJXscbqGlk8RrU+a1+syamL
JYUr8w2x9l8/JSLjs1UCG5LxE2xI18QX9X5UNo+9XSKHDADks9SAGWGYdnzi9H41BAMs1i2+EqPv
fY9j3dxXllj8J1hEEF2fmt4UnjW8yKuyrTcVfXzI9TVF5M98qjyMcNwaXr/0rGuhMRxCRcmW9rZI
nlDR9WAMekqarR3EgqZo5/oo9GplN0oP0bDTPxJPWPLEnRyeR/GHd2CwUPDUkJLDLoKojDJK+GyE
JZa9Tp0qflxqDKoR9nbu3Strc+11Ct5FDKUEeLyoXcu59cZohIUxq1JiszE7hZfn2Vr021TWjrw+
B+Cz5GZx96JkJxR3xyEfs7hMN6ARDSZ94ELWguWJubNTa1ntR18dDY59/XddZV3vJYq23XU/MHu3
qmev1QN4WYvs/czlwvan0a0AVTaEN5XE65yC5FsOJd0GGfidHjmndKAmwj8lZE8Tvd8FH6dHa3ba
IAVQ+KQTYBRJV/U9DmnvF8sao0iFRQvGEbONEoDfN6bDAEfEmYk6b0FIsflXUmPks5/pB7+aX2r3
MkU99f0T7lNjkycjTiyWlYgC/HfLS2PLVaDGKUIGvrL/MOZpAClYGQiso2tvmJvUirGpSjKnvObt
UbeEzN0XRPAuB6iOazqxw/eiuS5h15tgETmQ7A92+tavo4p+jvgwZ7dm0qdO9rITmljBlZxZtOho
lznhF02zx2HPDoq1uC65Ny5prF/z4Xs0r5RjmLDv1l4yvQc93XPCABVaY2JwhM8yHrSm6M/GHX2Q
M6sfSHP7eqWBrlavKxijSIBS/uT+3CB6H6HM0NugAQ5dKtjZb79k9wIEMcCYKBVfxkrlTp1GJoWC
MTidopCoklAx/G/1+0bD5JPlLBIlNy9Z51saN23fi2PgGvm8Z5p5YMCCoyGycx/RzsqZqg0xyTiN
uLAZItobIr8aUe0HqmxNpgP/iSSnrdRC4ZPYZMg1x/7vPbpL6/B6rumthYZxWu4s+7Aq/5qS2N0s
ApL39ONBZmjItzeJNmg2OzJ3y19pv69IpQRsUf94n4PNLyJJVv2/iUPGqTZB4+nLxk7z+Gz7Oscf
v4EVeWqIYQTuRMcmD67Oo8m0kByODVNfVeK/BK08lcTtxfpcSxKCMQGnplLpWcuPfeTRfoKxS1AJ
GjJSUXRhC06YzdeHuXfVIWIRpT9Ytm1SwuWShJPQVo6fP3CwFGH+W0JoPg5ysDai6fHRVr+RyvfT
lAeTBpF5tRXnKyKnJMSVpY4jtUT85nndB8UKYmFA+MtTX2Wk+EAHuKDEVy02rR+1EBdDj3PQLShz
fkzAUL4fTv0iEKB4gfm1vEpyVSqe/SMGFKgouIBegPBJv0GNFB1+BrS6ymiM2jjHAmPkeE5nzD67
h+GxUBfNVDBnE5tKgcv6Vu52obA6VpYVJ/WhRKPrKjPNmj13b6Tz3pp+RFHIaiE3YkOeYOWjRE0P
fdrPywVrN0FqUHglxZGDpyxTpnGu4JNv+jQ5auugNYYjiqLcAqy+WRs3zNxfqmoFYKUn0OTt538C
2R6JNfi1u0Gsmkek+e7Kph7LBy7WQllWTwmmAvTu5EnXQzEBnooVTME/IKNShMKxZwsXL3mf0IZc
ltRbc24kEGdHM2jxo7gB2jfWbAaS0eiwnYRv7pW87KxrGJgbHngy34JShjoZVZARlTAiCScyHkBQ
bnsF4OM/UA0sbTfOySDj6aAAIlC3vR/Yz3R0c7ZegQ6pLikeY/Q5KI4mH3RDf39jvs1SGY0OIbGL
pWA411+tddh3Fd8BMSgTGbYz7lt/ziMyesSqlfancKms2EcbpstAUNlqnJjeW6mZaZdm49+23NJQ
5wwKrc5foSdk4WUHzJ3SaO/lAnuCFMPDPEmIjc4Ik03xnQmRG/eqFmtVFfuM5+qAk1x4KkVgA+0H
VmeChWvksOul5j68boIgRSOp9qpqDVWlSr8q+/bXM19dBt+F+MjNAnZNuuZw0IDTfz92pSXtyi8e
/Mwv88MYx+LL5WTQR9YoaESUF07OM87SYDfIpWvg4pUOY1e3rt8HHBGZiblEakjt7n0zEBHZlK31
z8LQO4OheDGfuqEHqq7DUZeXP+ajF/9KkRm0vU6GrmtN3otMswixXQSATjTUbvBobqI49rLJU0kG
KipD4b8e3npTmCasMuX+ljL1qmHSdvIZxF9yOBcLTNNoIKjLIJhd7m9VI8yOuriJHa8bzVqKbFTo
zG8bTgi1+8MsKW/OtSap2ePM092C7aT5/ToAOOcRJYJ3cb/R94MZbz64Q5qmJJMXgk5uIZbV5fzB
BFl4FxDqvcJtYRSx5sARUXR6rTiXnTy4ULqhmVbr9WIYBLXF8XGfQgF2HoFNrYwqG/jHhr1XTXPg
ArB9ONS/2cWznmPQetmm024Ab3R6nng0aIx6Fg7tExvepK/U9PL4J8rvpLk6ubvSeuMM+K2gXk9D
Cuz75WQ0LMrjQtyN7MguEywLqLuMOc8+iozkH2Q5CCycPYr+spD+wcD/pNglRjoC9x9tHIOG2rHA
v6/0CDviqBx9hhqzu5+PxtO02GzZfPBHuNF5kF8KtyTV/bdWUFNyuZmamZ9mZimIFfspRPHS4hVo
S/V//UKaZPSM8pF/34J2MhJJAPvwXVBK/vU4Ww5zLcf0Ej1HTH5mSL2Eq7Vvy17LpVOfRe2to0IV
yPk69obwp1ABtRJodaFRAsMZo9ksKoJ96zgERf1OZE8CaeS5c2zSlWFxMmJESiZBd2qC96q6zYDk
UEofIQgTAMcI05me8aSLWv3mYGFVRbjyKUy8SVtX1JQsKCw3NlLwTPJeIm2tOnrd1Y9NYbeERGia
VNIb2u52UGA3KxqOWON5j4pmP20dNFsEwi2bDTlZt70TKv4yyFHRtUfGW+7r7gaaMPVY4NZ1mtTW
mZO8QLxqZerMtWy5t4lKGf5kE0uxuMdY7QGtMU2JJFCuRB7QVuin14psS67BtWAX3IsuhoaEU53y
vBMOwTPnIrnJqcBPSMfKklLDYpR6NXrinOxIF+bNBnR+j1/nBvz5/ncB3IvTbSLyPC/ok0zYioqP
5gX4Pnx2UbEbY9UUOgcgbqRK/LZ1VOtMC7IZZi2Ne1+2RZLaQyitrzvwIrbkbPmmP8lrz/duMr9S
G4gjQGhbhMx1U7csOxqPrSEzNh7A3yfQU39J+vohw6W14ajC+Jn4Ve02jTWFPFaq8CtpBXNb54Hw
NaTstXLuazHTbABozkxVp/qNyHSwpihrBQI/1u0SjGR95Hvdyucz6loJsSBD8DM0YEooGWZZ533e
Pu+ArAueNh/PnSqwNqFmpO/eHHfV3/ezCS45SEuzMSj11FX4Fr+lVsATCmAnkLgW9GEeZ7iBLaax
6mn6bkRVtdBS5Gf4SR0wGoPEvpplNvrgMcmOUGJunZWdAyP3x5qGO23xB1pXjr04YuJcr7FXwGKK
JWFXbdzstyNLuqTOkMXr+ZrjQ1jdqaCCE1mjT+8IVm3Txfhg/26BBbTxG0ei8tAbzfXmywvIdbQB
2XC/S9ognVcDklS6I8AnW7h6U6th7nWCVbv5h52wBNMBkbb5igiZ3Qtb2DzTAE8ZUFqjX3I2LADm
uRV7Mj0ylLaQopXt3PLHJr9pp9wEf5T1AaXJKr+Pw0Kpj1QnhuB65XmyyBFmaj/i50MKpiDJzAtG
wHs1funlybR2xeCJj3383Bnv+x6P3vMvDU0EH057nfTr+BrHqOimxY9SZdltqqur8Sla9aebo0Kn
YXJVIGPFKlYWuAysmGwTyQec7zP1KNOR1i0hSEtRwgg5HbSgWBzajNTW1BBa0h/M1hafSS4OBEBx
TMpa4JNQAqSdjOb6WPbJLr+BrfPqo32YQwt0WddCJT5oEveElThE2HaEUCrp1SVU2PaEXDJvxuVX
4xQ/Wv7X2TBXPEQE33JZBba0vXXVc2KHP5pfiOyeol6Rr2sMWwkANSyY0zNuBVlN2DTd3cw1tav+
NOuRHIJtEALtblw9xjU8A6oTMvXi4JJWcToUWOPKH5kSzof0yUQpRAJOy4IeKz4j5nF9VFwaPWhT
QO5AhTk2rdIwzsWybANPzkqgc8DvIPeAOZAx4QTjPJny+VH+gpjh/0fu1ckN5NvliRHDhMbJK0dk
mgpLhgfxmbR2t3sRQgNQtjaXnFvYfO65tgA6QxQGbUKu47+aDkgUmWrBnLa64lB6PNc23CSY2OBo
1dCiemzfLEQgtvIsDuF69w8pcvmDZsbiqC6sQk74+u3/tvpYPZIl7tAQGVVkSZwbDz3JzATEIOGN
wF9mZx7n0xV14v16ej9/XUR4oJpMdZ6EBt1dqjzvCcZtXxt01Iz9ej0X10sw3FpW9GB4l+6PkqiH
pDUjjjcFdLOqABGKD+VgsNhAUkEl00lROj+5+xjRHqH7giI/EiZCZDuQ2ncIX7dtur69pqhh6XEv
9qzviHBptsigpY1y0QvMzqJ2VGg46rFJZPDCPO9BC+1ogQj7iLI2s5h8A8Kf/NjaHMUTcr66OgAO
6vW21mSwGJ6baa7HFK5YxajjtV8P2qcfwRH5T/UUU1PNR5NGiVmIzqYu91CrhTQgpAUPCVWs/uED
r8G4e1oByhwvm26zdfCg9yMFyI5Q9OEI8sAF1yPfZVX6tnkN4I3YHfW7ZRsr4jPhfG8p+gwvaadJ
iU2ar4VRc6rpg7LF8Mdw0ZHkWDts9Rzj73HcwEK0ipapKfWspMSVas2UueaxYbWeMDoWCkahX2Yf
ZIFRQeRZ1YAlDt98BTJH1cX4QUkQXXUJB1nBpx7BjciFPvtujxp3EOMjubtXS8HPTs6J2XfrtMVV
MRZjHu5Nyr9wOuuNMEb6Js4uH40X+KeAcPSSqF86unuZ7cV86t9/kZndMCLXuIwUSNnYJnsGnUTc
VGx0gOxb/4uG4CQEMwOFPYdC46ygjdeYndK4dzk76yS9lRHuEoyUe+CvrGWYlv7aCFLfxmZ0xNiF
6O7eIKfwFUdvnw+GFOkJL18RfLaGnqpZ1zTqin4d5msGIvnP+rvDaFnwfOU2kEM8Edie/uQxJkMy
iMJpqzTU1GclJbq61dsrQ5CXG2wALu8OwWIlIDh8E/zJGTQnjJRL8kimsxvIY1FEMzIErGAr2/XL
4wZADeFXTaGOeEAG94kq1bUvGWT4/cvhue63wtDApUpDgvoFq2woS34LL7sSfPEM7WjHoPX4yqfp
2KDjp+/9k/guU8rlezFroNUgchlBQjwBAk/AIeXOcBgD/QSEDQnOd80APrwgu5hEoTpUm0AgeoKl
Zn4Lcyg2YczjZQ0fETDjgeFNKbNBfc4vLXxwWP5KH9rpDjvusOT0H3SpzaxUpx1xDhSN9cb7y9Sl
O7SaHWNNaxmAfEjE5wy0w4M7p5dGm9aH6vA0VtCtBGAMoRd7J4TccUqiGyM0FI4hRcECV/hyx/DJ
EJHqHdDNq12+kMqlw/glxyFWZCAAgT0ZI9sky0/AAUpI+hfl8JVHnVN9VuO0Vif7d8wWL5dkACav
fIVRd3ay7k7K9+x3bEoqyoDHM6LrZfoRr/AKqNYNs2IaPeEfSef5Hg11H0hpgU5eV48wQcL2fslU
VguBMF/1WSjsiZTs8U3iAJtVvUocywas6ar+a87tce2Wmmlom+6hHeB+KWd7AydPOlREpF8q8M+s
IXVl2B5EbohaKVkznUhdVcrvfzj+oBLZgVfd6f2mxCvG+XDy5gzsLKdSEtbeDMUS4OiN4r7q6E6f
2b3uFn4UoyGx1s5+4XceQchPMGB7E8OKDMt/UjGKqTUceYXuwtstjXfQ7TEva35SOG+Xito7K7rj
jqcYMVpQq6+Kvxgt+FkResAW5VJLn7A+6LVArLIIQhn1TxsVI/6ksrupRTPtK4hGy8vjv90j/oG7
2NIm9WQNiZevv5u5ou4M+mTDcw2z2fhndagMFYJLPfzkUPedzcSB09HxrEdNQtpVAqYgBzmyOnM0
1Y2x/oiKqXtwAaXqVSNbYbO3I4pUtHsrVJ74qoewGsOV7jiI3bdDaEbQXk4wpvDgp3CTL74+7o56
/w72bIlsDGklJGYVq20A/1JwGAwDFMZ2nMxogOwVucjSUVxZhR+f9Tdsgh/jl7np6RaX2j66OuNE
BSxR0dGUEKyFHItovDgmLBNwg1jW0pkS4HF8YXAdkI9Kv5oh4kLZtbfdRJgsft+aryA1o0fBKq/+
RXeUEd5eTnMnV2f3HvHcetpw8PGRKOWO+lpxAPaRigeY+wv1csS25CVRAO0kSpHd0mpHsp9CD4ry
JaVTwzbwkD0w/46tWYj36jf9HQNj63CRZ2qoSoPqhUWFXHom26B6YrtujzAtXK8zE4xyvhxdV8Gf
TUAeCHYquqYizVIttAj3/UhB3w/3xtiZlDOu4d+mqvMfdjb4SBKF2YiEdHwxwxm2FuC6WJwSX/jG
JLX4ok0nLAOvAL3s+1XBL3ime8cfeMH+Vka95lKtTWmATgQxncEtIBDqPZICe7mTSc7HYF/bwfQ3
e3XIQa6xes/CSAi/krFetcRfCedJOaFffb99omfUFaIvZmY5HnelUR0AzqmMBCbAV1tBCDUkSICD
vefuKR3cWnGOIznHGwfGV/hDABVeti/ZUWRSK8FNBP9avnyTEFp/kHbu4VqGomCdr26cOQYkSfZ0
W3tPDIv6jos8BoyUW2uyyK4bsrXhdKgiAkaWKF6bdo3b3ipKtjTSPGbgAw1Usjo+q0xLhDU3atBD
Qukyqp2QmfU+bZz3ctE4FnKWRl83VS0Ptpmm6gHerV21SiBmVyVncz4eQMhXc2Oorg+GMwpu/osq
8z0BfZE9odOQhdyRL4OP1cTuNyDFdWHyW+svALU4P6YbO8u/frnGxuVQ+QgIUgjmBZmQ5SluL8Op
U3NE6I2VlxBZUHiJXuekB0+U768wiW0xh7u0TNz4wRNEw32BhdaVESQRgvTyIRLyYZ74mK2GpiZw
S3Z7HNab3Bsyku5mz4Wjc7Pto5mOr+wK/DFkMXxuzdFA59T2nYgBYQx9p78Yn/HKbp5Hdh2eApBP
5v434+uqEtPibHpDNtMTiLHpeRLyWPJL/Da7rjEvc5SH8vPnkenc+44XvGPdRh5TXfijvDaogWVv
X36YevRKKcVl4Q2rkyYPQEjHF3UJ4i8ifPl2x9f3hzA8VxNX0EiLFUH2Am9sWsoQiovNS7g57TvC
WuZT+GDoIgFD4703eGCpMitz71Pz9aX4sj7fENGJpfJpcevvN3rce931zSSrPx/A5VkJ2wVDbthi
Eky8QJdEPP+FQHT6/CyYZv4sBJe150ulrq/KIwV3FuH1QV5VOEtBZMmymZUEufOyir2QMbBZ2GPJ
NT9m28GNEkpKGJT2YdVVhNGxcAmZJUIDT233zDnNYe36nwicXMwiGzdpVm5ajz7SQYyxw79h4VXW
4fO8Itrcrf0H+R5Czab0vNxGPkiACPh3JvAoRAGTt0UQXy6tLAUsYexMR6maAkx9YDoJq2B8SzLP
RCx0OdCYuxljK8Vf7kWKpJPXtbO35FFXs9AKzLfiiLxQGXlZF8WLu4MeW80rrsTkBDugPnfwjbzl
XO8KiysmvSX3VWNE4KipUgSC9Joz1a/G91hUMviOy1nLWU4Eamvagu1eEDwwKDxreDfto2MbBe69
Y9LNCbZvj00mIEVKUGtGqRZAr3tBTnNuFTdNJekmN5f1QL/MKzBBhxW5voyDKY7ZnuQryiu1IRtj
3mSrsFI8HrcfAuu8WtkSrn0mxSFExATVL/acqmLweoqEf6+lFcCNsyy3cys1sNxhCloroAAMSaAH
vXzIk8wjKWb3qkHHcserhaHPf8N/TQA/+5tBQ+oVHaO96kWLddx2sGuvvjtbo6u/t7Stl7zNLCeY
H09xsIgMOACHGYeEJnq580ppint7LP1aSka+MvZf9pATl2EvBky5OBRkt2cme1rhp6RH8zg5ZCho
81L+BV9wEsnf9hG52yyeKf5dYEZgKXcWVwlxeIPZHwInM4Qx6bsvxAq5t+IpgK9QpjW/R768djZr
Go7OTX5zmLsZkrxgQzCHgOAA+gfkVRRZYCrez/qB33SuG51QyGEROPCKfnX58BM8sJ+JWI/2t6Hn
r+NYVUtdtGUlGF+K1PB8g4Lh32J/DNIya7PEveVA+OdZW8X6g4q3bbstfoiAo7i/8hAoZU4Z831h
2Wj+OynVzyEGMEFDShmcEpSLKMLvB0YOo7/AdG+Z1jb7nRYzhRPgrIUsdJJi36UXh5KZNoHaqA41
KbUeAay0rk07AJ8XYDJhI00RR8aRODV9uPtl0aRjBZ/mDpvWXX0CGxSKUJIhBHe7yvFE4d+peLRA
wqjwWd7oivcpOhLRSglqiRsTjxowSGL+KrIs8XYX/mNv5Du0+ROUiBN28idPnSo1Ibd2B3yGXPCB
sryOwWwB/v/sAbP8QVSmDGgQWsm9JGX62c6Z9chcGmKwS002wEmPFwWwPDcwOicU8cVRyoSD5Cbc
l0TXKbRSQ7DER+M7LS97n2YGaNzwTZx74/TxF5HkcBbXtr39lN4o1Ej2B1MLr/+TliQDmEruna2D
GVTOsS/xGtGDjepxzqz+hhlA8ond3Em/ORWPTuyjHpLlrmWmV/oOomEjAtOAKQMiyCgLwVMOt7U2
IJLcjyWfBRPPaoOIfdAb9SaVfbMg44bCNkW03ItBohH5inLyT/zEPfEj54uTSxu4VpgmAv4Tfu0/
2a8LKoP1bWYHSs3kyf1qtFw1DhD4s4ho2Mz4Xxv4L77ADUqDcNlWajgyfr1r0esxZUJLHREC/css
H71+/Wywj7d2nBwnhnRsLozePDcYLQ9dbF2bxPfeRrF4JISCoaUqrd0wXL15n+75gC0kglChaR77
5WIcG99jAM0XygwovFmOSmjcnF+UGQABaP213rvShRNXhhHIdTAemyYEBf4oEN1xlHR+vqX8i6iy
CcFaqiAsvslYvyq2aYNgqbNy752J8RE8DOHZ/e2iln+/z39QaaCAhV7jfa9Fdp41mQ5OyszYjL1G
d25zevB0LlBEfx3ZtPeR3xdK039R9+YSBc4cS48ROu6QNKInZNj0syTK71BkclH4MvMr9Ye4rykY
M+MW48gthgCUMMVIEWsIHef0wPMAKDihuuBe1GpOFABaIid5O3BJlNRieI5Hq3vYYrpJVZBxNFVK
Od/3JFqwWCyYLvfQqrRim0ij/zCl4VQYmObfcZmMCK5G3CYwp+ag2LiNczGRG49M7ZwUWhEQauzT
HIUczg25DCOKQpaf1tpp224i2w7jVKhfKkeS6UdNWyJ8kGiJwEYs8GYw+bMkIWejRQ1QNz417A2D
v3wPp7DE74ehue2XhHz3pAEAaaV5L/AZCy31fnyn6ghMwDNzTciteigFATllgnfPRAmEIg4ys+gj
YBKJKgV8sI60MUQW8+t8hAQd53h4bivVRKo1D7aKCIMbeqpF7itzVrL2h2ODXT1hbQzn2w6Gutay
TqZ2WqhmaPGipZjRYw9jXozjU6HFCNwIiMu+I5e/fRitCQcJH4ZFczkA1Z/vXv1JUQotjXg2ZlhM
JB91N6YkDeqvRuSmx+jK+WPqd88M4vb6Y7ztf0ZmpDna4Hx0phrQdfRKbd07wV7KfgqdRUSh1D5K
EihqEf58pF9NAFUybHX4cvj8Ytv1OWTgt9dyv7fw9L6kU9hzY3zq++SuyD6aonZjW8FJlNDVrD5l
CgqacLMpgoS6elQJw2LlrG2/vRmmp9VYvmBUym6u6cqRzD8d+J9ncpw4hts53zpnjKFrkgr9OZE6
9n/rr9Cf/H7A4ZdsA3akAoetO3iisWKTcP63Y1Cju4Qhy3zZKFv+q9N8I5nCsXzuFz3iGdEBqsTu
xfG6TZXivs4swgTYNYUuzylnxCVLHigUqfz12WNET4O9eKJZvgthbPNLe9wSH5qTX8rIR03cqIm8
jEazIumlTNI2uHmAYLsxRQQDwnw+FCWZAPEY9MmrJTAqWwDG5wKSoC/vfMCIfwclwy0t4oDV9JSY
DZ+S3mqxvV+wMfcVwBDgkChXXDAkLtKLc3csPifYRHpTRDGWjWcSXIa3IZ8JHUOFzmMXmdWvAw0f
zroqifC885jcT2mOPm64r0oARqD3gou2TfHtdASuANBHy+W95GOlp5fLsmpRzWhxk/by06u6hdKV
P7UbkQmk1+4WMAYdwnJNqjSUNLHeugMNKyMjYHD17+mBSV4q/X+hKu91sLZ7l2JDTnFqXR0Lw8Po
m84WD2b6wGmgIpul5PSgWMIcoVR37KoCmAzVYZ+wTxQBuebxSfGZgt2kEeInZViQrXKdDt+dXntW
vmKXL0/rBDN5AJ0fLh78sB/EviHuc0EV4x4vHpqfiECff7sAgjkgk8UQlv6qzwleWM1cXHs04YJ2
ZDF2W+D6x/3khg0z5I4tM5wAA9xmgGPkw9SSXkMrD0ADHPDi9bc5N4dEprqFoNDKJQ5P69MGz2jL
sOl+X6G0AHYlCHxSTFyBAIex2IKsHmx4GutJV0JYuLAkpGFwetQAOCpAe7jre9TdjmRyx6ZvQ9PS
tc5CQan+DWtvehZyVKp/prUob6orgvSKQ6IJF3G9sXlbV1EnMG7U6BqljshK+PMaXLutcjDZ5/vT
JXKghtOeqypx8+4CSgvCmAKcxE/mY/DYJrIsJ6LIooKZyJ0rAjZQ+QAUvGfTwKil6ZVFDH3mUP5U
HS01cCADnqNZP+sGPqS017ldvAxT5yPVKIN7DiPzpHneYwBcwyPqsVdckJDnN/gC5VmXZ30tiMzO
SxPQuA3c8yiyxZjZA2N9dYRHU8IcFLHe/K36/t2LY0f88mGyYf3fB+MHpP7jb6iDk718t3pU+hvW
hVFHPrhXGFrkiWUGVoERGqJVQmFDgVOjeFok9kULpHwDTrwcN1EeS0s585Mjvn9fbIgf3vJJYpEO
PCM9k5PfGq5FgGcMDhpf5ro359p4GpE3rX87v0O6jm/1qN5hXkj0CKDLIfd0F3coWbfbv3zndEaD
0qxWm9Xv6QmHUDB9MmYTT0NPoOR3ozOk93EmAetGPx2sBkD9SDlnVOt4ELLxiQC5HnEJZLg0X0NF
kBMSYGCsgTHpM/OUfKsThGu6uDM5Be77BQPV1PdzbbittAZeOZ6fCLJdTgizQ8IPywSgof9q0Jjm
gLqcWtT01Kveokog7j9tDAxI5w6htH2d9ZkEHBWl3dAeHcfqnqnPHRumNfpkY+603L52bJr5L1Zk
FAsDVef01KT6nE8xEI8xpdEGB3XygE87dUDP18R3tTLrXZqIOPjafny69H6EpxIz90NDn1FrDtRp
pQJkghv3eE++xj9+atML257PAUR+7W50XD6NEUX9lT6jx/CqMrNp4Nxe4gr+akB6fwK81dWuFgtK
vZa0jIltLqaVzvuRuT4o03tM5mFTdMXplI4SUvgkLT33Gj46kyVgrdqrS/5wtet4goHaqRCibsOb
JwtbUnJ7cuWDj2CMU991efL/UAHnPqD/0nE1ZdyHuo4oY53b3z/PvJiagYten3xQunG7Tac///UG
Bsad2yULejR9qCzofdbgXo5WPP+qwuX3/Hl0QGd68LTXjySXItnCQpoHZO7snbRZOqIPWcMwGlS8
x+jORmo9FuNc7sHCqlAc+RoLlYRUYaXJd5+dBOm4inOYiF6FWOm9TBg2fUVWu5YaNYKEtwby1M/q
FaEhCE3nJYQRvEfg2SurON+NpDQc2SOxTQDTQ2mqOxV4nEpxAFFplm020mRNNLND5cjwXMnLMnzN
3moovhpvd41bzuvrmdwHiK963s2tJQh/5JZ/lqVXZ890Ng4Ib6Ja0b7NUMfnVd4nf6x532YKg+zD
NzHZwqb3co3TVy1IbKoT46AfOWewGBllEUvq0ZloN1YsXslKMkfnY9dTzJOt9Gzfd66L5237QYFb
YQ1vtCONEQ4gCcKq54T9IfOPF531TgOVExsOUmzJgd25OPWWCeku2hAYjHH4jgwvGeJg+8+HTCeg
0L7wXYtqK2U68IWMCK9V2UISM3Hq7FBQMG/NT4BQhMAKKpqYQLjQltKMfzwA9ChLARFIV012ksgQ
ezW7nYCwRN139/7LE7L7nXZD2oP7uo15KwwriYKOR57SsbRNMjoI4TXJO3KqItG51MgmCiHn94dz
KYkbB55ixReo7UDHrWCPMVbbv71VzDjIFiv04eqSuCn+T+bNDsHKBDjWxhhFD2t2LKHeYTFDZvYt
Bveb+7ghVs8O5+AyvySbont7c26AazsHS3Li9AcwH/AIivO1uB2QYZOLoiFkJmzAVR/JZAUz1rWT
NaNK23AUlf9J6OiR/nA5XmesURWePdz5rR13CwNJB7YeErdk/Tj1KXkvc9Jp31w9QGDUhz30TRAI
Hq++zv397eSbnC5MYZBS8j4brI4zDmZPPkMAvp2G2nzNzTOgOGiJ1vmQ4+n7U55xr/uyfWCKNJHT
ekuiqqHW3N1zUO4WMUF4PV2OXWAmVQjdsTvBF2xDrOJuhIzAr6iD1w+WW9bozd12LNNl63eKv683
aXtjrWP+zsmd80Pyx9Pvsv1Sec/ejEc+p8+n1elim72zwqdQdjunc1+v69Mw+6FGvNBZgNsv5EeX
+sEEKetHUdwLLrU9r/gHYvjaIkBtX9Iq4xjOHn8eHcyR/fbASAc+mIJD5g9V9iBlL1vBnr2GrrB5
jadE0RZ4hPCP/h4YfnI7DMkQQKquwN2MxGuRoQLAkNIy2deBQrOBLacq7EOOL729WZa5c81OCqt1
rKv2kyX7k46fzmH6E60kinMWJCN72s6eyJXWRDnuNGqlqFWvolTiky5fIuiUbzMPgHtsWJQUvPvf
5O8U4ISpQow+e3Gv4FlydNmPZeCSgw2rIWG4i+zRApChKTLoGrx2Kp9U4AolmJSS1jFEqfOvHR/S
3HczNXJ0lHfckz6jsx2LN8StzvJ7SVuwitWFPGszKiK4T9D27tJRrf44ewvmL6JG6JwV7eFYS6jE
RiOQ3KLkoew2q/cgDB8HWwH96d29fhRQ6X6zPzQaZ+BTtpvVbsyJLGgQKTUP+Zwcnkrhq/cPHD8u
ktxml5Ns/6dxegivluuaRx9FTzqeblViI7l6b/ACZjsHkDYGvmQRjIpHF8HP2x04VJfGuNfbBn70
MxU4aW9fp7rZNQ5R7NUeHCA3w4NtjQkYsdkmpGC5thA5hB6zkGEutN37aALFN7R/Fk7Ni9gKweR3
1Zj9jMvAg4cz45q2zn0dp37nGQT7tKkDua1Qf5cu8RGC9KT6kz4F07YzE/tcPiBh8KCG3lhLnYvv
Vohf22TKP0lR/X0vyoh6DjMKkRGvruASuJcps3wr55kUaoTXzVNIwuFSExwDeIywFcrDHKI28uw8
+ZJo+3E6gjZh7c6XBDS0mJ/UA8W2jEzGeg2fyKeNc9btZSMJEtHw1gIghld+33ULbCYYk3oy1dsW
uNacSMG2+Nh9Yc9FpRDsXf1wc4oLLI6pX5gw8j5npn5WyA97gBdukqTcgHdaAgbghRIDeCVuW7gv
CsemXMUSplgdtoUL7yXNJUlRIzWkqyhvV50gg8kU7ytEYrxd4S+pS0RbUCezwWtj/OiIkAOCJPqt
UYP7hnGtT7mYkF8dv9J+j+hdCLpA2qNdbSM0PKuPNE4g1Mha5g3HxI4iJbGeKalJiAU+iEXAcaBO
+qbYh8oXAGFsUlcQcbzRofm7a5dqmvm0bQ+/7aW+JEkXgo+eHID6YRNPC0aodWhWXtsvQbCDsIRY
GX6Pj1AC5PSENT+v+ZBe4u3MX0o0qZ/oAf1SYltHZkCYmeO7v8TppqaR+ys71ikUvGTiSwlVIjIh
HkGcv9IsFUrmAhZsTs7VibewBbFkYFtq1LdeFlg14s6bNulIB+Wnk7UhzKweQ6CuUjIAS99zIr8I
7x+UBPVxNXkcXm45Y2NSqsbd4YIrbLfpS0ce5KvD2HQaOj1wxbshPhEvoRw74qcjnaVevitaoz4S
GTL1GNnks+T9NYyQzkshZYdzgi8LTX6iBpCrPOhc3CshtGa9qCC94Svofwjf5TxAInioymwoTC5N
fm49q0/VYypoqQMr6C8Ew/JrLZ6ZfWQJhZW11dEzwyIrRL4I5H2VCRgsUd/qIZlo83CATiSWk9x7
oJS0HfpUqs1PVpQ7GHN4ZbMY6vJaJLxT3oQDMyQGU4z/n7npNY8Qqs24yUpoZhNM/WNqnSrPDOfV
z1GDEkH1HTF+wbNcueV7zdRCXAkGUky5RvohPRGzZ3lWcp96P/xINu6jFJx/LelNpxrO4NO0z2fR
/wf9D6+20Vut3Lejha0+uYgJG/LxJdPH1aMngmeVA1+pF9lzBrMmV+EOu4SGaHLhcD9ww2eyqy1O
omznfdIwXgdEEcHSkQMIng0K7Tn4AKS1yQxBrQE4FQ1ruQhKA0Ol65cKjApQayhIjBonJbDBSuAw
oj0MO32DguJk6unEgELo2mLgHQ56i3JxuXf9Hf7h9Abj7SLthWiuzDHGZ//NH4/YywRIpWN4CFRZ
CL22LfT+XeI0U0KutC9yqV3Wi0439mEfq1r4V3Z7v/CdUwBzPeifIQrOfrQeEpr/YyrLTwUkyAln
jmzcaGjA0a1u6cAmMdaRlfsTKK7dtI3Mzekssrcs6/Jjged/yy8ey5UYx6aHpFKhr6m8z/poaJaJ
zerPG82VG8VAzixKF0nmU+JwQMbnnn8cTtLkClBvfHQlEAIOmkbu71py8ljMy+NmQU9+1mFiofu4
12aiGXg34+Sfn02IFUqoaTZ7Fn8DGQHkvyAYrrknUShHNvKUJVJfSIvbbs2XiOn3ups5d4vD3B+4
JrhynngRrIj7SywK0pKndVOydjZ6RUROLcFApAFcVJ5Fs3QReHD2Uu9KJPs9zZ9WOMBIlnQDc6si
si+enj26UqwGTg4oZGGWVYmjSlBjZZrnDdpUBm5C/vWpE54YBqYb7nNEyGukHbKlvUZb+WBfgF+i
q3JOoZLOdze5c0ShstR46Bn0r2zFdslqtgI24nAbFY0yTCxQtYYob6FQhFYU5GAwI5ubQsc+8MIV
Z52OJMEw8I5ZpO6FISqLnkrcb9KoQ7A0pE52O7iolGFwyyJFQ4ZrmcUqD2lsZkMPDe+v2AO3jTxM
vq8KmqRFuaDHht0gIhVX6Ddl+KtLfuOL5osiuwiCkY/M0t67h5n/idrkfdD2tlrAvcifivdouXuV
DA/8SJugvCroYgM1qK1yy7TOXP+VM9tK9CxIDNz7Xp7QGfDik114ob4oIi2XZOPZ/8QD2RdxRygE
l1o3acPGuUbohDEnd6PEl4Vl/r94Ng5gjVtdGdaRcaSjy/o8AncjCMdllOrzbGUeatrIxiNQF+w7
T2c0dhG1uhGRO6lquBtvvqfkdtDGy8jhKEGpGYRKxQAdPHtnmhDnTV6i/8PPkz4usKbbUZ/3r5ed
P9aYWLf6shC2TEHA8t0UzIayL2QJTanyaBnR4W86gM0jPhZehKOEbXBjMs27bbXcfuekjdAYpnMw
CrQVPW0jdpjCCMpQGCj7Wg+sdim/gcTn7BAylCyKCSZqisXGR5BF2RsQLOMPxaw0LcQIqI1ng803
n1EU/nqKM+fp4IM9iYQ5WslzYSE40qNX1SFEWx1nGtHRM4wVS4EVuwcWCMuU09Y/0YPOvp29KQ80
PKjCJp95w6WPwctoKK6ncW4DXxfmONyBdwm54T4rZYUDIxnkparEuI91EBUbvOCBOfdLgU2ESNCK
URo1/Y05iOswVXv2U83x5I6P1btB8v/XqSXD0ifGzRcgREHbzwHeGCgqV9/zFlfE3kxFQjbzKpT1
mkwJNZBPos1m4htCVsPc0geTd2igjip2N0Jk1W8uhYrtGjibP33/DMEiSBrtNYrxozpUaiiFEtVe
PM+FXtiXNK/PGFiiLJqkblse9JMgjKF/1CBHX+ViMoidghKGt9bbKNyKqfc3ir062ZjLj0MCfuWd
XTygrU+pDitBc/6iMsm9QqLEnOVpX7yGQXtbP3LWyyp/nCwcvDQfl4egWOV0CXs1uVqjGsX1UlBd
uuJ0mVfXogKYFoU+UjZfwMmnaa67a4CITcMsT4Ms9MLYmiusqTrLPCYdj6mpl/AZuzVAP3vsM/1a
j1CdbgyWdCwa9ZPYFGZ+eNiZVzJ9vKQ6CeCYC7pdiTEN7OWvMAaoSNFbqIatvrtgy12+wTyqxB+2
/qP0YztIzbKqahZv04HlZ2rYX1ej6L3SrM4JzQT4hKwj97/JySGmOggPKe37q0jDD9hzSlTwxkB+
dyHrRBu8N2a7TuRbPVjsw2w7vkgkrYgi+h8sOQEXSdxzD3WN7ud59L5osl+16SKQ0liJhtYWzmmQ
XPlxpqJwSsQzHiFQ41fuBgixpDN5+kCVmiLy/KooB6/ZlUTwZPkIwGHqfzWJQ6y4rsI1QFGOhN+V
qgwCKmFeKqHRoNWbxkU9gDVc2e1sA/d2J8wSt4pxRdZF66kNy8Ir/vUZMJTv+0PiNLOsfZgCpApv
J6big6aUju1aHgZQKZOYBuLehAjAtSTj+6NOVrU+KtUJhJzqHJGOdqqTfFnJljPNcrNE5MrAA8IL
kMStAaqI7L4axUMfj0fNOY8KmTOQsS9HznFFFVrbSpNeCTV2qfvkvyXtJP4UdGj8UWTHGrX+1pGN
9AgSvAUKD5Fy6EFiSzmwdQlgwB709sCx0b/aY3GD4tMx8WnbwQ9Tb0YLdlZgWUf7rL9J2mfjyL7U
6svz7c3eJh1hs4vuMPf6Od9iSfVOIaWTzB7KuELAwpNbin5EWr4bgbjGY4CuNwu1mt/DApxkNGhC
0tl+lq5LJwPsXEYxmMtDn0ydkc1BIofEUbybyBlmpKu0ijBkJC9MkZQYmFZjrBJq+UroTS3PTa0C
zpWiZjizrHuGPOolOU4QhAcTps+kBg4JJlv0JrBbMq0MBU4rlriTsK2vMIS5vrpYymwa4bH9Nb3Z
fv2bSXaFkGNVKL/XvmIGCuKHvg8dwg1/bqNmvKtfOzMQ8Kp1Uo0KoxT6qCkwvk39D2oG0l2qJymo
vn6vQXPzNsd1ZCgwiyrxr6nsvE0D07Dbqpc3YHKNN1XINrawb6VDpVlAXRXc54IU4vGo6bh10EiW
ZUisA6Y3AjohWDuZNINsUBEWhOEisXwMM9myGG+WoKobpPNOzWJROHYaZ6Px7SaFbDZMO6Jr1jOP
3F0OY72+bmOgyXcbAdjGtYViKogBwhjCZk4zK4mjViZXPAVd73NkRsnS1gZIXFZoz/+ErxduJycX
Zb4Ku5QbQg6/N9CDSz6oRcUtgOezozNl74oHNWn6Xge9ZC6ARGQubFx2UDax0dRNMREjgr6U+tTc
bHhJUnLDVfbHy0L7tuz02OufdZI6hUeVgou9v00wgilfP/KYzxokzjY667wXkycUkhi796fTdzFd
Qscnkd+IAYJx3f9qHB3LCbEFhgUoukrDNqUZEJ65VtAWEXtmUghgQNr+6oglVAS6QHY+Mx7DSXwA
8avEJ7dozIczsAwjn1X6W9kk8oHltaoYpv6SgOHjCeQ9BjBhk2PTTLTE5YaXMVLKJXhWg+DmVjj8
PjlHlJvaL3Lr5JcRhqUfzUf9r1hOUeW0ZhDRqlRK1mwmccffumeGHx7ly6FKNjANnubCm1IsNKdb
eBZBTutWqDiaq6IEbZkJW4RptIHgC2g3+VjU4Fkx+GeAhENDuifz2SYWaTHCLazayPiednyjVtDv
tqzDDdQj6ZGJXxIZIVBZCDivxQR9SMQy0BPQZVS5fDZ3niOQoosi5I8GIxTt5X1Mwo3/hc814xx9
K1yD1gZnWWyneVVmoDZXCwPtx0C0PlxD2i6IL4ng2uNSlFAu2vHjqlY5sapIb/+2TZjQJAnWniKR
WWMlCGR/5qexToPvrSbFjyFHxmKI6t7BiajmqPreMdbTmcGcC00BY97NpeU0BpnI9o78D34so+Tj
G9Q/F0He3BsNJhh/E03ysYPTOYj5BeAVuTrKRPi7BMNJJrgzfGtt7fryhtIe/q1kig7z1+TeHoEu
Z8G7gZmwEZaMmmGMMREMlaa9JDq9N6+0gd/e/nfq2mAF0EsSzrjPNupnqqqyylUGdNA5PQ7LERns
7jYVS4QO5upcoESkcbhiWETei/s8uMd+rqH2EpTS/tCyszVJdhgOwD+Dcg38Xf4Qvm7yFAjwptml
MLmM8acfk1EZWO1X5nQxhkNYft9h3xKQK17eSQhadwtZ58U2NXiwX21jmDgw4LDZPrWu34aJ++zf
oPRvI8GgCV4riGSbDInXuyDWClInxF7fBCLUhhARM9xxUfxHsMPHZgw4antARNJ+zGnEOBPgMplZ
KnYlYaj/3oB3YHMP22LmhlSaj+69I4EQHdUaHa09e/M9ooy5f4pxSt8Vo+AeIJuutkWfA2LHewoz
hzW7j1wN3K1O8XNPEYvJPvtHw18YwlFQpHyQuQkrF2CYUm0j5dvNir9L6/h8jpelQLsMlb+uk5CB
YPI9wtaRnR3bYxQvoY9hyu9alfFyvYHm4kxzxcJY1eU2tRlIoGrXGRh6yY8rPHuSoR6WMvk5IeqS
TcilNjF3CPpirSC7ZV71VvXTfPstXPEHZ7Dja99f3MJdacSNNb4NQXoupZWQiZHzZ74iQfmCw552
7+2XrlMgt/T0BlT15AXdBq0AyRaLTOwiY9AX9H7pqEcuUZF3HCnlpg5Tki+7E9xP6VagmzYZ5ZAn
0lujTjop/SDrY0jtErf/ZA2I9W/1nV8rq1gFHN0RbDylvb4avcOQvQ3LtXW7yz9cXMwe9Qrsp1i4
mwn6j6zvglnh5DSbpSWRIa8pspiyDd47O1aBXBpFTE+mB4+uYibkhmIkUYYtR/Q3Hwv6BwXk6Uqh
2MY4RyyysOIe4c8xQxhTeDCme3kHLGf/0ogjdfd8n+fV66WeNUFOat4JZfxJe5+snxgNw4vKln+g
eKKCLIJadu7MDWaEkBew7D9hiajFi7O4Vm1n9NAZQgEZXCLb2r6D2/D3lGja7Gr5nbQn4PE3BLMz
aWtlUTFl2qTID6xXGw/F09sW2/a0QC9Ym7eRrOkRqPK6pO7Jx4CPDh0xYR4xfzDi6IO7VSikQiT+
vivRzwne191kh0mFh+YGz46myNs19Mq9EiIFKU/qrQUiEBwmbCaySDPIWUP8GIrRU9bYtGwoCb2/
AWQOX2v8LRUejEypXGmJFCJ/KvztxvvwRUUEM1+RHgp9bepIIuq+b9LPp6udQWwPU/8sKi6ntd/Z
U/S4Yt1XQ0JGcSgdIxgGAjI0K3ZDfe4uG7FxaZUJJt5gdd2EPhChgHMzyNqiwKPOZoQh9USt4bS6
i6cggtNYpw0Bbxs+sNJgFRpqxWD55sQKG/6D7cZiE9S5GUqaMvnZUmS9x4pdBE93fSz4VdxzA3oN
tvP3ZSvlGD6OaHqqAvpuoXCUWDjM6Lc2JvpSuWvQoyDnL175U+A/jSENm2wtEqevTPAIhS0cDTzv
NG0nwk7SkBr0V9xvb71Kvo9t0vgfKNMJV4AgqfYkzRe+K1nWsxuhRfG1rAJyn9FzF+WJPzXMzmM0
tFjcdv739SvEFOTbswYdoaYthUF3TiLs9BlUZ8Ik5EdFGBcv7y3dnjH4xoViH9wUtij/CIHqtuJg
jKO9sFkjt3hPTCRNhqK4UrviPQKk/TU6TTUvse3zxakwNE3u4iVVg7OfJZSl3vS2+z6U665/Ljv2
NKaq3JadbuEm93efsXzT0ijBSbkRzLYFJ5q4DAzThE+md3hQoBYJRfLmfhVI8IWJZLzEjNyxZxye
S+iQuYaBlxDHn587O7vMtdhcfPbBeIT/6y4vrP6sJ/gx1K4pX/UNP1THOTHEbFcHLpudg8SbKaY9
QMmEMqXibisTGWeJP2lCjjKzo24HlHeBSf+vwlHEZOlyHFHYn8uN9EkFu74Jkp+wlRkax8DwJnTm
fQTV8VUDtxn96/6IRUJ2kcOIEy0HCNjfdKfq5Bjw7mkpAUHsR4FyBSD/hSGgrVyxRwbXjjsZDuzu
W2FdNqquggau5mHOVDQp7oBjOlaIejzYXHdRYX01tvq6TjcabRaFTjfPNSdGNErWWfY5Pc4CICq3
E4//ylEd9pgOsjCsmdX0y/XgXux3kEqwt/S9gDMOcPQLQRszN4CHELs0YhU3h5JrqIq57eeSqb5L
oxUl7vQmwDXSUIsPL56K90U0xdusNWeAYEq/k/zFvFAsDaPWaPTIxDrmTQXcK8OFbENC2CAIO2n2
oS8aQdARicZv8eGrc/BS/rAMMUy5Bus3DEAL4N5Kp4YSldHi3QexjSLREc8sfwQ7K7UVFZmxk9Qd
Ctsg8Tqmb5LxJta4+qQDkwny/CacOWDkCQqyP1jPEmMMrxN927dnAAIbx22DSxPFcItOtuuRCc0p
DB3P7g2hTUL4Jyp7JEq84Mo7N9Q4SSqev4Kwifiwh0JZRsano2gF7CX56/KbHKMPqVgWep6Yc5oT
u2JJW87TfhCO0NcsjeoyZ5O6eA82sHMRKJ5hZVZQJ7H0wanfhh30AGQMHfsD33l5M1N2gyQovKe7
cqgSj+WZW1EYwgt3ANNrHThGnY2BsgdUaoFLmfj9CxWO5b6XHI21XzWAfgcLi3Sw3oxc/5x6LDVK
80uKqLnUZ+aKng+EUt/YGTXYFKaDJYh32gny2tc//A11GpWYMQP0hRy2Zsj+0OeJn6dOQwoHZQQy
SMFojk0UGw85dyDy3LsXr3NsK3duRjwhRaSQvcRtdPp7FDTGPKsu/lWGKvz2jQdJFtptXTL8x4P5
NeVTI0nx3wRU7e/Mbg0eP0zPTQDaipcA+JZ3Ht1WlegISBtaAdavPOe2LWF7nDFdwJJsJbn2U49r
T0SaqoVgdlZ4RDcEF54IAAWyBV6e54mSLLMk+/GXLBd8vsDWNQCVI0T1mp4hdVhjsbaxVEYfS/rc
3SX76uQVlLkLJdLYQR4X6US8y6iv+Oiz9KLN2T5U7q39v/lB7pyK18vhrgR3/CnkVRtOXSJ5Wnxk
rW3qGBR8ur5p5m0BxFJpiZMikaQcuMVlgCp+hiwCsFgKIglozeKbREOXNw6OhMV2JPBwQVzH3fjv
R/acWUUErxhS5tv5/9CmCifN2F2abu314MLpSuWDmLUAjK0plwJTEb0GmLRuIJYFumRzOqwXT+wh
x+Dzg8M9f+nhH6SjeiZYprDwpUjMqTYjMKgnXhdFjS3CJR0KEPYFZfeuAjRwtfy1A8/bRyR3FrTR
iWQHcpNxdwhXcla9mVmhQOzJATnOUd2r+J9ECC10p/USf3jgBMSOAXSoYN3DFHSAWU/ngRQOO/Wb
XUz1khjy45fviJ9Y7R1Gam6XdahOyBIuAYGhx0DX9/25ItHuXKjh9phtW2t8TR75iF81Ts2DQUGN
57PNYVco2n1xJBdx7vIQLaeE3woPiw92zXXzdhPj/36f+jv5Fd0+9WfNK/ZarzbNLBIi50ObBrx/
7DSONZiVu72QeiwSp8koj1UA8nnkjchl1b7iqWMbzenO7fscZDxjkSobcWRwObAdY6YWkIZ5Mvn+
996EvK9+DIvdRRm5ybXaL18PIguKYT5juRg00ZywAv5ORGDTQZIqfpj455Dw4d+Ks/P7Fi9breco
UoqdwB42Fl0tsyXZDsQXZRnORAZIBgQlnPdGo9kQuz3/QNMc7UsXD2hN1CLTAbTVUTqI1yd+OIxE
t/teOV9ubCzJphNbavWFs6Yx5bsi3KKjgua1mAyFi32xfNLcxAfc0DCmBu/jcLR5TzBWeGot9fMZ
+4g1VnnSt1gHdk1i4UTRXAB/Nq6KyIeIzZinNi5gHp0/ftVinlEBhLV6GrNE28Yrq/cqVvxISalk
WTcGh3gFVtWm76Yye1qFSSrfa+Im7MVz+APCivvzLhY9M+qBweze989RfURO/s6x2u+7V+GviEOx
FhMQGUUy5GQnDtTQ35JeJND/YsgXhObptfIY7T7eZCHujFIahGbkUlIZlOJUf4SijRjlT0oOpKn9
/6RwfVSnPSQSZEiTwQqQUpki067CgtfN3yBQccPfgR92n9M/zUwbNsxYnMDkNmSE7EC+OcuBfFhi
Ydy2BvOEpDn2AdyF3pXjZXRCIfnc0Jj13s7WZCSbFJb8pkskwjPOFU6PsyAf0dB7IIEITHlKp6MC
/2ToaSf7ysqXJE2lirP9jx1CU86EzwiPy6QquEVK/qETnN8oZJGULKKDHPo2rQm7fW3Y0xIfn6Yy
hyGIhw5xj1q9iYHJ+wSE2jj0R0R7mLFpnFYEZYGVBgftJH0uNiJ+lfjjkQiL8HMhTHdzQ7CxCzxm
aQQSATfRUBBQai97YOx+uf00P8Ei61FT1LpxAQUSsgGszr4HvnGHDthd9INcvrlLQDbPrTRxxdTR
0AikKzmjuvjlUcoJ38Ceo2hh1Ln5W3QvuxiTud6gSn5LrpQ4HxkjF0KHCH5yuzsRDNhL3skz1DPp
HSS+4V6fnhCGE1sA26DHO4UnlN1MY3DMwcUL8HkaW7r+dPQH2DXjv45porJWS470n/cEadFZDnQs
l+xZUFHi/ZHTZnQUQQxUwdkhygF+pXcNglvu9/r4BoncGXc2EAa3BGuRzDJ4iAPg06+ZuKxd/3yA
h+OuQaEsjkGpZZ66E28bw/c+2ocA+Bh09qxMf2v2yVkrrdhA30kZocT3F4Rg7o+bqJLybPYz+mG9
ZQMtqWNsHaQqIdYL9bCx3G77cp8VMtw77GdMen2Yt07Ar8YIkB0vGM7iWTTwiJfKGi9UhgPdWgQD
XdPGwdkPnqn/7hYKqpdPq7RZ8frQHr/UpZUbvXvvTj4wzYr7K40vB5qC6EAlkdDBbhEvITtnflMF
jRm5mBui5cHRXDbrInll71DEZmSdWI/0p764ynOk76/Hc2mF27hEps3sJHqW7v5yryMLukrN1r9L
YjqtxD7h4ThI2IA4lndDJz+1NwqIi1szCHff2YXrSs3dxxLJ1PPFQ9y+Fh+mobtkGCq/BEt1nlM5
o30kaY0aViiPG+Uld0w6nvChm2jidWpZWi0VItvzC+p9oC+yWUbGkrFttTC8P8Qozmm3DIm7uJMA
XEZ1t+wKQphGcp/F7UeexCG+p9BxoXEEmrEaS8OEEss+zHDwCTXow3Noqy/EjVOgUJLj8FoHAxhd
7YTPiA/H2tdzYmpmvOCFYkzPHDgjT//uXClM9oN7CVLAeBMz/yVcEJ35CeMTF1y825d0umbzE083
E9BJQpH4Q5WURwMn3oIN3ANNXMWjjamUJK8eYH3DbdcXUeQJ6jKj1X9P68vWgwYV0Tl+UfU1tBd5
ORkHfoIXiV7h18LXGBGQV3UIdGygdt6O0kbzbnnr0WamdpKwTFPYXyoMdGGpvKf5GO1Okr3HEnGX
sGUqQbDlWWNRGHhXQPpS8374cw0s/Z90t2W/vw9Jzh9WsevBOQg8MBxbJeT9FrSTmhcpW84fTop1
ixnClBgiA8KfSEfUjXfrI18ZOVlKzGBOwHqfyb+K3IKAm99mKebOX6pKq2yF94LbHFrUqfHUiLhG
7hjBBdcllhjU+Qt45VP/vrBXiHbVNBNmniYW3js3GBZA4gEbUw5iBTi33nNqBW2/BMiqdJ/vl6/S
i0cuQCcwXkpETidNefIZTk0gfENN3tTXbpxp/zGOOoZ6WTEIHJF8MNLmCfgNzS0xhe/d4PhkWIHU
H1BtOZDJfuI7tHyYiKPaIK/peoJ93iCXbGhWXZ/l1ufMFLqZ6a+roJimQ1thlybWD/Ky580qllC0
sRWx2pOYut8ToFdog1PxIcmovvbXAnDZhGKQSdzkRS8deHYXlaTU+wUzwePi7JRTd4Pit1Ha2i23
R3Gf6qX44u1cKSW+qqYlNs+GG50pERSKdzXQPgu178WqtikjM2fttpchygOmNDhFkAziL9oKUORD
QiHWE1pKuLWRfC5arVGqhi9YY8wM8iz9Vj7WzOP054nS33X7KGYSxyJpXjoauvoppGLaimkedqJx
5T2qC1pFUpEmpFlI5ze7NuY5TpxG191BhXF5JXmmWahzhgGLpUptuR+jX/kprG0d0hN/FuPFcJL/
vz5cKYsBxQFnAnyjdWyItLOCWhGdnoMSwqFCylUlaCT50vvvlmnzv3BorOjOoA04Kzw0D5j77uSt
zeooalrsMPXKUxTJ+ihyNQD2CzAyP/jQFBCdFZrh+aFsJPGpEtYX8qSOLxEXpwWe6rgeq4A7fg90
K+qXGBgou9eZVFjyo2ugDnlkS1xJZp+FaWGUyXUlujR74Q4rzpg3Yo1/vNOmoBhiL+ylc4nyvF5y
nHTpp5+LJAPmO1MIbKlP48ro77ica3+0wy0CJo5bt5AyyS5JqmR7di6AjM+ZHKL3fj270kZ0CIvH
L7kSlqI++LnyBBjLXfeDYB5VGyb/bInjcgYnetzWjKYRhZJo+uHXTYq6zw9nHvyfgB0I+pi2XgdX
K2WT106l8srGk4IpbdAdwjVa5a8LnPgFhytmMYOa7yw9LPyhlqx+3rOg8QjI5UBcx4fWYkXGduON
kSXrzKdXjM6KdKh8+vT6wr47sDemvRAFHHNFXOto6F1qp/UPyE/Ml7ZmDFvs91HUOxcrZjC1Ia0z
RjwmP3RBCVACQaOhR51xOi07QSfVn5DaIetW6kO2lMKv2VBLLrRv5hdwYYRY1uLcA5cj+e6jmw1L
+DZFQ4cNQnI4dAlf9fMk1hk//vLgpxjgfYN4C716ZxiZsmGzw+GCBJzJ15zpN2Xu6mgPLbY4iNFR
IP/HkPLkxpB6uAYmO4exza5DqjfYGyW0CD9OxuwhQo8YsrUcU22SEovK1VjXjf/ST3nEtcE9DgsQ
xY0hIOWgkCS/DhUd9E/aC6AZJaF+KCYnAmrJn5l+vZliZIH5TJz6Yp45edBggITKkeTP/sa2V0j+
ywnyzu1STXlmCL+MquqyU4Wt3fxv+yt1uA70gLBRiNP7FycpvvaDd9e+IW0dT2HDxSVnxeeAurGz
kPMPhjWhliUPwJJKQM96wN7vPD3q5Ezny/aMtzsTR3JSvCMvs7W1roBTR09Wk/XwetASvrIjq2Px
B8eHnXb6w/PgYEHs3U/KplM489A46gtk2FivucBPJdnsehFUpiv124qT/H3+pzjWqIuEc38qdX1n
KoIZaEJyx0fvpyPcbtSV7/1R3j3+MKv+BNNRW7X+eBWOiKbTZ2mJS0n6y0prnkZQ4s81qAMxqwC/
PLxN4EySHf/3LR4chSC8o7MlBrEfZkE/cze3FULbAglov5Ty37FJm2YUT9PgsankJ3QGjHaVJmCh
mOhWEHupGhA/1oF0fYMxsFzQTgYepY7gSsRzfVD3b/x/0dPaUWjrf37TIpnQV+DSGDGrBloYxCQ7
9WsSCiqNrdwOZbK6Sc0a/zONBuMPY3mtI1QJP8qX7wEw+8i0aXUHXncHvosv8UPIRaaAGm/f+ekR
eOdrusKl3ti9NOapDhB9Cs4s/gS+97UD/hAD9T1NMMhwXDPV4HnsYV4LxH0xLEFm0CFbm+2HXlvb
sOGDsRi9FPS6j70diL4vboeNBiG1Txe7LNsv1qfC8PFY1ST7BPqukzcVyCZw4hx2UsBs7nPD38/w
4ypMplMH5xlI9qcCtPK8vMo0mA8p1Ecr/jPC8VZTPGSLSzutMD9Zc4zmxrpnJrzCGZZiRzjrkk1q
o90IREIVFhlinXz2+t459KPL9Z1GEMv3qsJJyoPcBSukITKmLXy0osOyZ6SqRMgz8F3sI92sHh48
+utPVpyCCKdF2hUVthInkLYarjk0/hxofdlb2igCErphiI98oNJuQTrPr+C2+3Jv9+LuWwaE7eLc
ZNU5pZ8OlS2HCSvMNRISH2zkQVpctSTILqS9ZuDB9+aNN+9bSDyHRS5I7FVfA7o3cjp2LJdFJoPh
z9py9KstiHwa5Opbb8BsODwzpKHrUZKOoMGJylE5HBmsNPLWT0DWhcTvde+y1lS9e9NZo4egP7tI
1PQGES/ali2dohjsmSXPRDyR9uWhqQs0zDIq/UDoOnHno2LQ02xfpCpmu8xmuCmdY7EkxgCGe4Qv
hj81R6DDMBVtrw08xtB9xuMaWHvPOfcLAMQ4x99ZLbHH4SdGIqp//562WbGhC4tM1jBKFf4cwS6j
Oa1iV17inR5jhWIFza09hj7msRptvZHAx/JPBAYG3c18S68XF5u7sXAFfgGKCaaYf/WnCZ45jWFj
Rkr1gM7PsSGUi/KmFaf47mJxWhnQfiaurCzECR6r9wFjQWJVhq/KHHqdythtgPOVPbDmc/fLCoPj
QqUcjBPRDDOq4M7qgPKgLp5UMPRr+/BYSB7nIW5QcqWru12RcNscii+ON48A1fmQwKGXN03wS6Ix
S9+v1SmQulNFKzMoPG4tgozjXd5HWj3FKPgrGIh6/cbXa/4sZjq7N7ZXycesDOlw6gqVZ75KYLBs
sGbdC1SS4sLA10M7D/jiv3tyaaif+kHIFznOWHySY7XuN9xfo+DN1OtpTM2HKD7MRpt2dDrKloGj
c03vJ9Sch248yGVdHB4MONZbjYvmZpfQkgZtL9RRXppAJvpCwbcwCqBv9Wf23O2T6GOHTCvlN3lq
zfPuypvIRSHU8RVEgc3wUUtVXBAhO1jlvJ+TPA7kO74TPXCjqzUMShZ/5iyiaubqHYxwXEcWtyxe
GuBdxXzhLtkgYxJcOg6WY3Udw+nFg9tAinCrlbzBcktder4Q3EYcDI8jtTIc+mFVv+nCcG/3r8m9
EGFoU8O49jiWTL+ntZ2XBHcYM6OHod3s4g1XMHOUph7amqDoZmEASSpMQ67snESIBFkNddk3SVx6
L+rZ7ZspvYQerwH1ytdPhLui39Dlq1eVlyPCvCwCNrzm7p0/OJayEGFXCtrb0T6TNFejOmKRiwG7
xSWh6eMfh8B/UvcpiE7DdA2wYX34vt7idK2XzyNAoac9+xyYUUeXebz/hkda3MZuJBybc6971G7V
CZ/jd9r8f9qnWupc1yMPTf2vdgzRJns9gQ+TCakfn9I4g7ammUVr/b8d2Z1cAOg9wKUc6ms6JO+6
TbQCoHTP4ndpQ3TrOe6dDcPRf30owyrUcemPruZSG4p1v8lWvyc7QsBGx7MGxPjwLsW6DjgA0zZ+
P5ev+O+SjFyOTkmdZNvtrRf9283v32Tc28w+ZgahvC4YtMnBQcVm6/tXjgEVnfKs8FIaXGvF/rpe
w6njvU/BGunVuuLwRxeHQN/uOCfrYnaEOKV8u+6a14/boayjjGn0RudUTK5gpp/FXRXz7GqEC/au
Uo3URD1NDCFpLGKUQUo2X0iDyYAQAQFG+S2FD/p6hSE0Jfwo+YbRgiSLuMQVQBY7k3cmrULu0BD4
2o8bF/oEmyKpYQVUC7PwYU6WF4QfmN21JI8YR33TCbuNsUuvRXacRs0U0XOfD6W74OcF0kEFfYuz
+FePftCPW8BhMYzfzupr3lfdKRiaVt+RXC2Nv9sKxi1Vxm5sWiebRLm7mMpbE2/YropvVwCqNEk0
BBk509dqa3cG2nLdcOawEbjXHxfwO15GROB0Z3GjjdymLerATdPkETOqTKoivM1QWnUOX/ywDy0U
+em3TQJJvEN2fK1rEnoool+UDm5cvU9wlgddwJGqvJiWZ+BCTTfv8VqzR12fEWlsDszhoRGuB3Lk
qSihbjHSj3msxDEC4mEAjMi8nDd7MSkBjz2L4Y567MB1/+i3oDBHmvT9Ii2p+98tZJXFqquVvpvo
FiQKyp+68sekgXS/9WqNgss8t48TT13IYD7hBpcfk5RYes2ylleoDifoYKIRPKYsJUMb9UmhplnR
d8DCamRbmVJy8pyDoJs1FIYt8pv65bY7hG6tW/dVXQg/ySUpnej/NJCvktL2zf3zokECKH9ZB7Uh
lEEpCcGIadSSlYsC7DsaLB6jcTN0fwEygmh3LKcqQZxFLQlJlec9tjZQCz6BG9pNtgjGz5Dg4sct
EcSnFXtiKaSj4srrKijJ5jGt60WjJmTTbUGN98zYW7TWfBvYY19ex8KmUxSTggMWbtlx+DoLh72y
aJKPqJgCQA/YAkEkO2yjzBddt+roLkLKMWSvqXY/9GoUN3dQX3jP3yyNmpj6coxt3vtEiz4g8qyU
FvgjCV8p+TpufuNi2Ftkfpf2ihF/SLShagwSICIHF06qU1juc/FsGObNnZzH2EyfQGy+J81X2uJz
qeltrPZV+SCEcZiEgqlR9BCwEpBAkE/b/Jlr6uAhedZnoEFIrB1Le6jisOou59DwincTAmKaSmQZ
fCtKuifJD6iGrZIueeLGFh9Nu3tD5FyUqNuY6lv/aD6c1PHvISOL9HzIrdeeqt8ZC3XdE+pxhTHl
BG6Baq3RlUC30i0Ep+omzes5gDmzkQ83y0aL3uMVRzofi1fbgHl0W9fviJzNGTtZBuV4BF60unB4
0X0CPqGz/RKM7MLsWTJylpINbBlU9aE61BSVbZjTyL3OqaZaKO6/re+JpPh2bn/mZIcPn8+ZqgUm
PFMoQM50gp45aAEuziyhhKMlNW8+2E1mYFFQLzv0gzzAfyukSTSamRnF7guG/PYTw/uKl/RNs7Ml
r47m5KmE61+a7DfRMgjy5hamGTdxpOd3XLeoYih1PVbkYEt188hik8c79rQazrU1PETznwcV5rCR
zY+rZt9pbQzZrGjoEgeG1IOBai9g73usaC9uDGmvlWGx1iNxXr11YdARZb+qdChI3Df4MpOBtO3I
v3DJ1IIanGpI7aB7r2R/JLz8ZiN5IHm8eeuHeoD0dCzoIyIROsdEoMQf3vUjlig1OiiCSJVJS2cG
IBOygZ26J+600JAN4o1ENKlZfB6rcAHW7/mNx/cFADMXtOyr4N/usbJHZc+1vp7ZucPgW0PZIel7
qbVvTxHkQO6aj7WT4AYyeGbo3k4L7MtmDB/169LcoqDuyspYEAGryeLc8IEgR0uI+Z8qXp4hrgXW
cayEFJW6WBEtb/R6+/iy6cFhW+uPFVoVE08J2zj79vxc02EXzehwtibEUZ0AANsBZIrKD+TUR/+B
nixh8fTMlnKoi6qa3aVLlU4BaoS9xd+01GViERlRj9sRuJKcyHIIUDKOyNntia3VTJMv1hCS8f2g
GZx/8KaUB+/FHl3yfyeJloo+j9PKeUAL0rt18QhbtsT3NiMJNGBNd3ExkgNhe7G43AmVqYorZ/mJ
l4gQ+KPVIPZnJZkPWfIODtz2hmnHO4lTS3GRwTjxXSOZ7Dv7lcrPsgBaQ+fLADwBGAwCx8S091qc
XcRPJc9HaLf6Wk2sdkUto9Wbl+/ahCeQYnKqjW/dnitB3tB5VnnaQPWladI/UGn76W3sqcxbyr4r
B//i4utW94phQTMK9dHpKzdAqnPFii8FTs16UiF+a6PddIPrVeIECoNYFuO7tfHPq522ui/0KR5T
jOJXbUsp3/0o2kzgBtKlXTG8HuNjQEqbVAepAX53KTJP04CefhP9TIHnuuoTPsdLEfWOqx4jeDVB
xNyETwklDBzwb1czbZSYBKfkivbhpbETbJUQL5yqyRTU9L3F3Y4b2EFvYxh9aWtZA6Z3PMZKthKQ
2CCIBQJ3x14legSOkYRB8LDwW7EWWa0QWkOvOJni51ijhwq6+jVtF5esz1v6S5w6lKuBrsDDBBMm
IhYuWvMm7m6zV7uDv39rRS8LF+Fn1nJmeIlJfUJbncDhKYp+r7LIRum+wSpPeLcuV/gzDG5GXSQ5
4n3VzWFjZGt93OvLEeNh58BqKIK3MzOPjqx0kC5FpH0un9sF72y6631hUo8VMKdhvB/LmSdOCn7E
m9wvQMGXryv89577udW4EHSavNSpbSvXDkFeTn+bM8dtRLXJJ8UqIRddh1SBnDXyswfYwYGALRB2
LTP6g7oODU4rxdBkMQ58w+cca0oySClUdVIc6aln1hByiLQ2297P2QB5qZZY4mVc7FTj4m798r0W
YDvb+16SV12JXy0Bm+hVuKEnTGybiNweNeM3SpZxn6FU1iJ4DTI3OY4b6ujiFUdHho0QB3l4zsUA
L8w3CtnH1+6Fv6qrX8+PfZKjY5E57OQb96ImI/79dMKkbpB3gb2H6FxjJgUawzBVjh5m4kP6O1iq
TJ8DFMdlOPKaHORUt4kpnpnq/VZLg2LGZFOIkduGVeX+PIu79+1VnJpj0rjZorkp/UNcTu76hfKW
OQXVM4Ke91HSpgpKwt41+A/+6fPeoQffRzFpQp/Yug6akxo8WuxCgvkgt3q5RjfMdULOu4em9/Ag
ncNwRYO6MGvNYKWZW538uxjHG2eEO5GvkByXPlC7pRiEwDa4OS468v+0o7UoNQU6DYwxdWF04n+w
/AcxNA4bFFh7+wiHvfFsP3U2R7hFAmRjYtR3Y0TUcAM1jz965i6q1OlPd4eayHAu13yRqC1TnUTO
vt8GnEZSFOduMkcGFP6Hze6vikuY0E7gBp/jac/HyJahHCs0+iJTebXkGvOjVVj9V2exJISCuHii
guTGUnRqxEjkE6XCJs4gJeE8dArMU4FWL45uufrFOBxdueZzEcrhSz/Ab/SAjAoamIP+kSVM0UE5
yu1/k2nvbhzKmdGJ+4my5VX2CNNq8NXnBNs4/Cnasz+OOcXcxA8VjjLZ7LOthYsSBi+ut1UiXi8Q
bl8mGa2FQGiejkC8BnaT06IJvs+91NPllFsWAn0o/FqM/GYp72TCQ3s8aZ2q2pN5YybDyYyQ3u4E
8JU1TPWOh87vvaRYn0JWdHDQewOWtpZB1DNJrbCG8kE+ppkhM7KPU/eYJmuitiehbp6xHLYUxTN8
/9oNF0SAKT3/I1JokbGZ6HlY9FR1HK1WAE+h5F/05i0dn8ybB7+btaatrrSRoYmfsrBw4BJyxWUD
Jo81XyL7FVQoJD20hQrxJhElEss4BCoJewxkxjo3l3SACVd8mgWW8jRONRKCgRNMrDeB+x2dIIHS
j9KqVEDw97LXTUuPsc0I9IGlLocRVHVp4io5CKbd71RW+X/W1x7WfFsZ4NT7XD9aPGt+695DgCRC
qV/T32hNJGxvkMdb5h6fiLshpf899jWsVMgaiuuKiZkC57e3lILEKQZe6XAXNWs83XapJdbDxUzi
QH43JV4g92oNebLdMQqeZ+XkJ7lRcsBHRapj5bwGBN7xM3FM3X8Z72d0XYbhq2kxJ4I52kjCiOna
8aeIB2vQuWwdaTa6B8dtpKx5F8XcrLU05oKVn8DA1FZeRHK7DspgGiBd6FOXro/hFt2HmEF2I4EM
/9ZzTBV1u27el8xYpTrcRJHftbz/8FalnWq+e3sEtMr073/42bDNIjk1VUCvBsiCXJCvtBHTR6HK
kPEsu2pBgefUkKesT2PHNyUi7Bae17pCn59vqJ4oKk4oS5qrrVveHgNn3f1HqBdb4ynmYs4Kt64E
zJ4Gewqj6bopItKpLXYTYmqNBHqL5LdJ6Frc4ZVdB+0V37FeM04vBk9FR88nDJdEDSNidAw0rcXc
VSr/dCvjLtuOcMzoLcr14k+X/mb8Vr/L5Clu2/LNw7KDlgnn8Xz6xaYJ2fzwJVOXOZ7KkqYq/V6B
xzRYF+epEoRR76sGUx3DwsIG1+Efjkxz0tYfQEiUwjy0rCmYDFf6nVWxaV8tNfK9f+BvphGhC5/S
fg1/fD5dlXCs6AUDhQAquELDZSzZNLQP5zbHhZTYVKbe0kxznBMIHZPwnFQjRzo6vZNwM2m1QXx9
mAoGE59Dh/qxFH0uhonfM9+HNAjjEHp/plGorzXOGKgTIaTeKh1qCzE57MQw1PSBZiFhuKCU3S9J
iCAZoC/fiInSIJAyqtgc8//R49KmDC2DC2CAAD1nAH5qH1FhFRUDShBpJ/qPaspOtNeTdHQ3d88D
Qxfrqmw2Vi0VPvikKAQJZIbVCQYQs/9yvefNng+bPAwuHHIdtdPeTR0RP6b7KFPPZfXTeEsGGzxg
ZUPLEKTFSn6PFHoZRqT1sph6N7uf0J5+ApF1tFSPYZ5QciC1PXNb8b5r+qJ2sHarsz11Am3Jwsyi
YGMMlTNDA/eUdtAMgB7k5yZ90YqXV7e12qzZAH4O/tJEW3DVcL8fcrZIfjc9ZrzBRw+U8kq1J/4+
89jv8x7Yft8fdIjij7dCqhdIXQdp3mv0HioX4noBjvquSAyiax1QqDiibrJLnyfZ+H3W4weILYev
iKh4iGfbLnP6cEUJvp1V7UKaAPaqLggLLwGJUVSKWITeDqaBQN1GouBHwU3UsAIzfojSWoLrlHBm
y+FqAY7nAST8Hr6mpVg9QhaZkGQ+Gl03i1pjNcY4ORY7Kh7K6HfrJCjttOBIrJmTbUw6X6aVXOON
PK4rMMs8lnbvV0jqsHyns3OCXMR47r0hM7AvEKkhKqUJ3nfdfmlJ/jRKTPayiG9yW0P23Juj8a2i
VobXbiF3aGCVwChMb+FKaGw+4iOeZCxL1Zuj8CEQvvtRZjcfCMW2xl3inqxYliVGlJj+eIkbijdS
93gG7fCHl1JoEHib1feOM+tpC1H5q3rinCzthhHMpF37DnsQ2v54THDoaWfkztni0+95Y2GkNjHF
R03TGe8PAJ48N35UV8hTuyMNjlaZ+38zzJSjbjZJOEn1l3E7duvt9lBPILFrCpZwlSJVV1Pnc6nY
No/gNABHIneKs34f5K/8BqtyFFSTk7e9Oy/BkGHUGroa1D5RUdFMU2GbXw0SYjBylq0kepkzhJhF
e7XrW1b+M1UX6SwFlWue/r2X56mQLBSTWLy1AIIOTJLTF5wvxCLjcJiWwWDAhxFwx3JAJyFbkC4r
0E3xjrK9Sh5w04Dg/ACDBGDujE2hf+rrN5yhs4vZ8nSRK+dTUvHhWj3WkB1ybxZ68EWZ1TzFAGVM
H6cOPKWNXlJOsX7Gkn/j/BArmzo3pyqYAeW8yXk1WtDA5JajmVm71dRSktj+SEzUL6TllbYkRbPn
N3dmCXRVrQr3fFLYuDOWjJcm47wtVzCorPqJuBGQpq+SRTfnCAfxCCADKf4PHnsv6f1/KnjXBx+L
LS6dx7/8LqtIPcl4UhAbR9kAGi5tVx3IxIwz98ZS91D6KpAz5PFtnbfvNv/XS1P3kXVIF7ySJ4Vo
o6Z9DYkhQDEimz9nIk1j63d3qDGI3RlJgCN/Iz7vDTtDBm0KQGrqP7MohabpWLuepPDcGqR6OJ40
XGiQ5A6SO5IStuROUj7bysEbqMOC8c8sKlSQ5l2SkOX+LnRRrps+pVG101cPBNX59b3zOSnhX9Sf
Xk2GrzTpCvLFLp2JPK7yFE1X255Lskt4KOUgdTvaKGIj6B95dyk2+X46H/yAt7pgGHHurN6BIGA/
yQM6zLctvqn4g95rzapiYTX6JtvkwySFDO5ZdcA+N8xMGloSFYv8VasfJGAJmRG33ZwynhOuCEF8
YOgwQzvruWJ1ioO/n0E8gvy8ZwsDTG5P1ppGrL8sq/PghBBAZkZViL7nRwawsyFTAfudca2euQjd
GzyjlsxFyNKfFX/337m5W2004PlGEpSnug60TKsJuMMDW9sKaVoUsX/Xl8itwt+6t41qZyDwkWG5
/fRBsX1Y086Uh7UGIWTyQfMeLiut2Qru3iH6gqfRCSDEh4bLWV0fcLeeJcBXatA1b/Wb5ixei480
bbswUkvasVVddVMiOWdyjCf15oUcpljy/nKAj3WYISi82O47kH/LjOZ62Kvv4vfVodS92MKkg9MV
z5KWuywYp67w/bv22EDZ1n947TTa7Vd04WZPazLMNcI0DMqGjGB7Et93jyEFm7oL5zpqWhstFu+V
Ey6xr7DIYvRTvC7HGEsM6oipvEGNWyNKMLx4wjGCNuebhn8WXtBQUYTfhAXqRQUjcdVbWgHc9WSf
mc4WTVMMmC0KYboLiHNdo+qE7l7goskTCKICDKEMy/pokcmEyd+pCIZyOO306G7emG4CACRsxIhn
td6blEScX6hizPvRkoNG+Xh2Vrh2qm+bCU4nYMzvfzctvKbxxaFJMeE9FDi0fioGO12pE0oXNoN5
h4gbEpdg5MHlQrg+VCCPnJHSEtBYt92vX/8TiCZoFkPGO/0skGa3PJqc0JxnAhILtCawJcJ6LHbA
hA0lUZ87G7dRBLIs0JaR/fZOTsSkFx2CIsLVk9KZz1yH7079k4Nz7kVvIeBgm4sfwSEEr3BdA8lc
gToIxlS9NudG4aCS+MZpBpRKQ54fy3tV/4MIgQKbCUFfXeynlJ4Zez1uB5x3RSmyfoPIDoLZEcPP
NJqXx7niwrw5hbSgWtObU5ymxg4EI4sQXTjcDO8mXFURY5fIrf93C0xlMNlkIpDZ+TqcX4g+Ot2H
lKWxUNOzfDatVIevtYwWYpAFtpQjMUecTsQX4ZZJxvjT/J6sFgyCioFi0CAVUX2IZhbDZNlvQm/L
kF9ZYvURnmPx7e331GlwdQAQWD/DbtJfKmKQ2onH1ecNAnTU/Ngrli5rPmdAwJNFHpG8MrhSUij8
JSz0vnSLqCbuRY71xddMAbkN1sXxqs5lCYskoX3fDGjOeDxrrMovwUIJzn6rpKMnUl8Us05IrIgj
SwzrgDDfk2NrBjtEWuGtWSaseltjfxbzobJRn4Bg92Kn5++QQy79A91fzqBA2Msskd4mHk8liHnW
BwR1ihGbZJ24TxDzlP/ZV8OjPMzXS5oACmDfGTMNxaVLqraNHgsKKkM+GFeV9mKXdncuWPRKf3l0
00IyttFBZRkAmoB9rx/9E5oIK4gjcl2oQMRqh4PdbvipPLQSMqDPGODAlxYyFfSzqheqif+3rqn0
gAyIOLt4jJiSVv3NhS+R0qNjFYtefTXbIcSodus4oaQsBFLYzfArpL1eNgd6+FSHsvk9kemotpXr
JmnOyERCfwZm/P5qAi156txEDI4d4gar0MOLKieOld4/YEJqFfoOztfn5VZ16QupcEhiZlizefDW
tXcfdknWacUwmbZHSYcaD8djPDUKHRutW2QeDnMMZSNtHUsHZWuYKzKdbMgtoytFN5pbiettOj6Q
6MoF/fafmNHQF6JHFiQXmjy9Cto1u0FeX2GQG4ns2G+htkJkMsOSh5bjdUdCKI0/wLQ8Ojcs4by9
WfZUjhEZSw2ccKfCi7Hltt0hrWHPQN1/XIFRKyplmuPkjF6LtXYQ1kHOFkXJ81znf+P8VKW2kciR
aZfOfHZWMHjHUkLbWNRQy9TXdu16Kz8GTSQx/5+ghZFLvQcMRncW4WKnVTDg6uV0pzo+r9R5+SWw
LVsgh3eOuUKwykHdtEtm6B6e5CsrbNejksJrJjAkOtsnzCJ5DtN7fqhIx4a5M0+DsN1jm4X/HEfG
zPf8czn4f7sX3tb/Kn7PvFxtET2DZd9vPuTFoNz4qpBqBfqu0mCFeuxkFRMHiHCVVchdeA5OoZYb
B9n0hJbAfXjy76VfAayUvGO9cbIl8wxO4F93u6YJVVK2qNH78BXiCNdcdMOXWr+x2mE2LSoG3jdu
laGAR2NY1Np7mGLI8U4DEbBrqFaE7zMpYzFbbAEiKAgvYoxUq1ldAPRMoJcXwtkW9WJEVmcNPNr4
OwqNXlEGbnWefkCo7/ecB2WsHUvaaAfkbfz9SHXDa0QGtvtxLbW2l7plUWlGdaFL2bReKYTEgytA
pjwON3FYqTfnEjwaHKIFjJucQ1/GQbDVQNh1GqbdCPW/GXSq1h+0+g3T3fYULIKT6BPbp/odch4G
Tspc7vZBk5uo0sgIq5U2KsLfKGJiJgdQMp0RungM1ZNFjiwqcs2qE9HiqJr0XtHKsD6YyHlL1OTs
477vAB55zvfEqf+56yJLpXVe5ntUxbAxDcruYKffhTWsmy52YjUNDwEZIcQMPUsmWS8y9o+5wCbh
O+lkb6haabGL69UnYjzKclAmdu3p0n4UkeTJIxMEIjyqdc0h5Pn/yUdznCkQbSAsDpVGixSC9pJl
R2TKNYWuiyNmfuG80GIs+RMHc7uw+ts/Yr9MThtglRCxyePPWe2CJeM3BYktEp09k0hwR2ogI18s
FaAsPZirneHFkMglHL/+EzMCKOBum/k0UNBb6W5fXP8ZYP4qpnajitdMPngtnJVvAsbdkGIczoi1
Ekne55cTBDuqfTPHza5IpbPa5/RKTIL9k9ghJNR0MGK1ZtQHJXXv/hNzbWyY/mbbcV1eu7OACTBO
lGFbIXCjHSW5Vd8DtptbmurQCN3JR8oFtA+/+2rFCblrg/CY1cAn4J4v2ggGLVivSBr7sRqMNltE
1MtqR81ae5dAKHLfqJhGbR6/oHvUoA1yz1mk+dcgaW1TqNzT+Thx5PvtQLZVO/hSJjeml/a9Evd5
PFmIPCt+Exe1fJACdgZ6+SEe6Jew4agPdvUxLhtQGkJpzg0DIjOvdHcyqWfmgtXYiz0U+d71ktXb
ngS96PPguvAgK0IMAlp59GhNKWYPNQBCBfZZU38wg8YxISkxsUsaa776ietfk4Q+cCDNygabP0uC
zqfF8rhpBQQGctrKd6CCfiM7yqg3Cr4lz4O+s8lEI+DFKEs1/KnrIGqeqJvRVbK5PbCwQBliXfT9
EiXIiXdExa8B+Wp5TpCO1jCpnOs6EieAwNduaBhoQYw7S5Er58zN28sLv0Z+GD6puBlyC7/l5M+B
154k8UF8RmbCS8vi0d8TrMEKexJSkyBAq7fSgEyr0aNgWeJDyNTCOd1oC4rnRAE1vw363ImbzwKu
RJDFm3haXFYqIha3lOy+f6xPkj438CIpKIze+01stbtwMbxZR2Mepyru6YCGXGvsEPnkuOxBW7HN
62/7/EddG7Q+LbD+6W/YUMVQ7lAi25TOGBNJd7LIFctmeuU6Rcf7dNLIeApTSJB/13373fHqvxdt
3b6cJz/o2vkOp4ayF6VDy9gggGYWwPJFoKTCWqt/4EjGfdk4rQkUjK9FH5IjadV+NuuA9eAh4Z6W
PviHdogh/uFcqs+8RcjC+korj2EDN+fmqmpEoFQYpcj6vkY8NvPONhlCOAa8Vj0wOCcvN/i8OaSA
3MM4vDJNS3mV2wZcxAhZkpJZAGtL7veiUXCbMZVdH74GMQNal+9x/+07lXqXAoh25LxSz/vbV3eC
q3kXCyBgCWnsBx6+4/CYCcN6PY8gRXzcRT98WqyHC7QkZ9FPEIugGOBfrzWY4gtwZA8YGmD84V2T
m2+VyWZeQe20JDbcS5CZQbYv35J8uyN4v4Q3fNY4Fm4Demu7tEStHh/aE5E8n5TtvaPU1z09IyOe
tfqAYSmIf3GWhMqy5BFpjsvGpf3AZoVs6fsr/4kfk4bwd3DfBwhjOGyj1LTm/YvObwXEVnpwlSTk
pLSU6CzcMyVomeK2XD6DEOqqhfxNYnlCX4vggTIISdaheaFWirjYdTfSxJsArUdeadw6qMV01RTb
GkgCJhPd5/qh5/dk91yBRBA//XCwobqBnx/iDZZu1Ew9H86Lw6CbVM0rcgFUugvUM/q2/bovM/bh
J+xtv7TNMp/3NwheCTSZFfsFIbylfum0IQVdrrMAfTZeFS3mvBeQkq2qLGNoGbI9WNOLA2Tn9Q7g
iW9W6og9jfIsdvLSLfyS6lE00QuhAWvLbBlQ8MXGDP0tThRZwqgqj+q3oPWcZLmjv+PPDqSfYg15
i+QWVEH7Ga3IZ+9ZxY+N8zqj6GJWz5ZVca1Q+Fi5m+E8kW+f3QUfFeBXXItTxNZGjasgaiZxNjU4
wkZ9YdSvGMJeR+M6CBZi9QpRRxzXCRSqQIPJorCusgxz6vfKvJ558R/ETh8d9LIIcmDTWJcjovte
CqipP048d+IVquGpn3o9QFxQMmaJes3CWKAv5qRLmCsUJflIVp02zXEuV7m+g2a17RL9+gXmBN/S
89dieHDjG/wredqp0/mUGpeoDNsvJNnjnSaijsd4gEDSHwYA/24i8IvSWf9s4s08Bwk7k3JLHfcj
L3s6QxETfvEYN3msOxN2chcPCquPikebPF8HCApqqArg/+Aj58T5BnpCJq4FJRl49xuUbefYCemG
fErVAPd+yVsfsRgbW6D1l27ykeSCI7MEavNI0P55S84cRbuEOqNoJ2S4I/WBl6Nw969bqTc2jMD1
32+p1TIc+oy2YIKcILlnhMxUqnbOcQHRfEHp0vt9zrAaO9Op3ZkXkX6RIhG7IlFgITrjOA6gqhvJ
3nIUK3A12t/t9UoqRsn6TsVWntUIq/jNTIqiKa/dEMiw0xSNUk2sBs7saEpneXa0N5WnoYhH3vLD
e0+6SQ1VA/0sOlpCw8bwybTk2nXfAZka23DcvwwbZSomRlinUU7/ChBN/nJH8etcuMyLJak98Hpx
hBDcyGC9gmH9LgtVW/a9TfNCrrULmjmF/CVy4jzEl0xAKNEHKaCEUm/QcGSmgxUqkLNDm8xVMe5e
IsASP3GF+OkFRXxOtO0MqQt3HLAv1y8mC0ArIvm4xcuQvGotm43UWSMiVhRa7jT6YmthF6FJC8Cy
MDrEzBe4oWCoA+g6Q9TEKSqZY6ZkysDWcU3SQXAdVgIW2ExHGrPtZvWurB/UQAXj/13/Ss4VFnxR
bJneyrfY8GbtI2HC8DG1R84d2+imXVz27MIG/mWfRYqUwwuT2fRGaVrZiDwut0/JvW7ropAML+jF
1g0U2WquO42O9h7ZwKqPDMOrYcuRWWR8Fe5EQjY/pasihDlitSzRcyd/0YBeAxTjetFi0Td42dxV
Xj06S/lqAlQzX2AycKtaviMOFVuSddbd7KbnDi14D1EjVhAIOa5uhiCfNgoOT0GEw6KDfgmcXrhi
2Uskxf3UFwFKTYPRTQBl3E+m4eF6NG2UsjoGTFjEa7xzXB5X9QSmiRTPRmrdkl/o6xmFyxlnEsaP
WcJhB1EbzBEttpvrUHL10FOWVg54LDONQO3RlqSM5enUr1TFEDYqyqQBYtpli4MRHpSrc49Sje5p
6TQGIhr9NWLBotFjpG7Ek8Rllf1abhAZHss/xI9R3xvse0BE5M/Xjl4W/lu6+iccw3jQh/ri27zk
4cvKP34qI02jo6cm8jnErpnW33whLCTYfGFxYzV25BbHkF/khE5GmBRoDU8fEm84Li6uagD8hF38
JLhd2bZS0xv5eI+LcwapGAlyN4u2w2Y2Eqh+dZ/xBwNXV3OwTmxCCE3JfY6zhVj5hnqrv/DF1sjM
NPxxpNGLFVzp0YLCI+l4zGso7igqttLuQTPldcMFZrybVf/b6Sif2L0utwYGO0WzvIIWpkwM+ERR
Zj1vqdipHMxwoRCyATRiAJCeIWsBEP6EeBnW1AQqsdJalfMYX1Si5T8laY+D9AdDq8rDVfvBXURy
2gWEyEhQfAvk8p685xC18xaNBIoNg32vs4dobZD+oGwczR+2uve3mtkSR1sa0ELQxSSpPXDTwlQK
fxCD+vPr9U1mDDUZYzWaz8Vf7A/68v4UoVCzb3PXJCqRyJ3N51f7W2+wNE6eokziSOE1FQFQRfKk
3bagmyC6Rr5Z5hUVfXTpLqSnNBhtp8un8BnEhNFyqYJfhnbYs2miRt3xFXArG2FSKGr6qV7dIsL/
nct3ZMSDUiz1meygXE1aZe83TNpdSbPXMeiYeSZ+Rp2cMZB+Am1+mA5w8seL2CBHIZQ8xGk7z+uD
00MhcR+MYcGFVeANMn9hMkTNRtMBnxzWxJEiOlxGJnRZJsDZBhKZh0F8+2sHXw+nkydqAmwInAEf
6Cs80YTvR8zv8bVbkpAJZhv/RlB4HjhYz25yb0nmm9Djyfaaw1GZQZqfyED9qJH9yji5hv0j5s48
5AHm8AeA59FxD3XO/U5ejdi7nf1Ow/Ow4MXIQNpwDJ2ZXt54pWBjPj/LRrtR/++DzWfMIOc8usU+
3NOdUwYP+XqLyFdmufMSZ0QUwiedKKcX9eVL7jckeeXY8oOJSxidlDpaA5f91GHXd3utrEUmh9ZT
B8rbwbrcA3QStV2qkCTF3EevIcByZtQ+XXsr1Hsrcw1kzcVzPPHJ3C1TDzoNgg7hGerg+B+sSIXM
VLyAOlTOHbjPQ7t0zych3NBINNUrd1s9JVEZTBJy9tqu+QR63y1lJpGKNaH+XITbOrSg8B7Z8yoV
/5rEJncDYHY/5ltWGL3CRT5sUB5eWpYVHdREbT5mECi/nKJa7HfhjDmhAnzfBAiW7aNGjQVohoxA
JuEkdt9z2E9PYB+Kpca5TsUFNcYUJU16XTq8n3s2iTmOyOh6DT+pDUNJwniwUcW2XNk3esTjnoHq
EHU84bl40XkwMDRo7pVPM3jVjvx91TczKRE6v6j4y/RTQ2ShW9GUj2dcO5jM4p9kWq5nRux//+XB
/b3iSepVB8J1bIOzSYZ/q7RGkBL1PNvhfoH6mrh8i+UHTUckSTQmjS1udBK/Y99eBylsWSIJ/7kA
RkUzE5tDF4OnaHpGccvaoIu1Ocg2Yk9MN7ORXoARYsJYT3xqW8qzXCMPKeU5mEqeVEJG1hea79Kw
frsdZvgR206duq3dXoSGByfbeSk4jwcmTOy7BG4V1DdrP85RB+crrlaE/XE3w52NrgPjDaddecqq
ykA6ZT0sdLF04DhCGP/PayalEOY41I8wRBnFA7GDY0Xy2rTEg55DDy0PHTQOC4XggfcrOk/frmqt
NkFseZ+eEJE8KrQJgKGpCoHlh3kKh98do28KRVfxIjm845a5HbiXxmu7p6BNsBAwl8nP4MN+OxQx
9ci176S2N4lxEUJleAHJFqFvjmKPji6lYPby6MrQHszZoatAZXEVX7WLBDmZX0pX4Sr2emGs9oCe
V1IvOK9aru4XD/RLGvOoyt5PbkouNasHrYdBOnBUoxiDr3lvpNb4c4ao9kK7iToOamWV31uRYUzA
hJtmfA/obcrl3nlQNvIeQZQ0YD4Y5iNh1v2kS08yfSEcEnLoa3feW7XqSHW5k+1UO4Yy0hIav075
jldCCsIA/yKqk3j9y330v4nlp/1ppEM2HUqR1IpUtLt4THIx9dz5T07LZYY7lavqb0b9Q1nJTWxK
x7Ub3votlBwUruVzowbPUspomII8TCkHEp/UBo1uRIF2mrEMlWWYeikdMvD8B4LDzVeleEzjkHKD
dyxFzlFnFI7Ft1MB1zVAsD3RyjnYOS1Xd6Ce7X1REzu4iEzlHm0iSMKjCPcGdIHdYJ0geczCEdio
lD/g82QQIMUOlY64PiY0illXZud/4Q4bvysQ6Z8aMMs2ajk4UGqKk+Nl/Th9lDUQJ+MO6B9Ihum2
xPg7xdTJRRrn/+qzUadmgxXkNaOkYNsK60gNLr/TZKfOPB1ghMuq9FdBoHAskNm77q+C0NsX6FCk
sMMx3BE0we1zY2lokuuItYpBlOScuX7+aG2xPUEvsWfox9wgPyLQRnU6o2wgBjSSK4XnGA2LA619
en66otrr3/W6jg9tIuBeHMVaZ+mvU7orjIMCWfjnYO+XZamWsDuTfdhXoJXnJeJAHrabJOGE7g9x
YkZ3U7Ay8XWVCb23eacF7UGIXvMpubCb85ItDDGNGqpFR1BfF7JzQn+DdWk2QAjGM8IbbqIyovyE
Q9lZ7o3NkGFLz76iGfxfkjQPIV3RZ8elU8BoKa/CAh9I4h2fhUVphtDHzOvKHpfY/3QGPUdFaasY
T9Fg67QKBc618Lqb/crdjeYop1bheLgjQdkwGeYyhBeK97mbaglIewmUb10FAz6NyNfUvZg08AH3
ItkZs4nbXrXWMO4b8+0qw+4UPd9FkrdXHhrV+WsmARAsaaZZVvUmJbLwEZkxB9d3WI/eF+cXyxrs
JjsmKstv+gELxYkAOtdP/9N2X70KadRrmyqMcoRBt5kDmiE9F/YeWwmuG3EwT/KIeVn+7i6KH1O5
kingNBFUiq4YLgwBz58YPtFiH1guqkDKNP132AXSuqc6EHmLEsFk7Vn3AZqdqTnbzNEFYbv2Mxzt
+EzoVJQgsTEAqzzQ8id9qXAGUYTiIlhhRIqR/QXBTi+OtlHUyt58p1nIFGtpeBJfj+qhkNkKR6G2
6brJR0A/hkZQ9TtkVyVAAnUgh+n4+nZZ+bRPD3FOQSq+wZdZYh8BydImU1F5yxtuEj4DIGMlTfTB
uN0bjuGq7Yucg8m29TYdqvNMmKNkEJjTOZ85iqC+CelQi908x1oEiPGLfyLaC2KHc07wY5MIim+Q
Llh/km9i+NLFVauhEb6xoOnrfHi4wc4y8wG9nNAMBOz8ust+iqB7GqtzCH+U3cD78KmTYLr4wFKX
JKv01/h/YL8LgKbhfpFJLc6i1YDcXoDPlhn1de5Dy+WFm/qeFVQndkbEKL6dk1G8+QXRfp6cLSIU
ZYAhV+xh8OX2vrRlOZarMYnt4JaQht/kSmXONX4dJddhRLrg0QNhyeG5skywnFmEwOFEgc0/mrEE
S2M1Ex60cKHjRcNS8UB7+ZPhlGPXOqKzx1pTNoELpLCheIhDkH0RCycy3UmPEwGIcUu8s21CdEO3
gEWr4e8PZ/p+mx/Yb6T3YUuimDAbNTeIPtsCVZENv9dpHeZKQuP7FjWr/rwmZxj2yy/3BVUpKA4/
u0Gs+mXGZLdeUw43laLCONjhpVom0MoAF/OJttRJv9yAn9Ajy48lthfN1BaqwSzP+vtE8uc6+rAl
/iOEtFhM6LekmgW/0q7WLmxroy0eiNSIIhxHCIK72n8l9cbJBOpJGjEcKwkKuqte40wFBwir+PHx
3klbgkTXCkXk3XE2xQEK/UaAfNW5tZmHoF01QkfCEIly73geNDk+MqoBm7g1M2REC930PSJKzPpg
tY97vT6hkh7vEiA16Aop3T5mqvhSeOrjMCjrnk4jFTpU6Kii2ZxXju2uUI66nuS8Am3twVFfc1IL
+eSCJmHWPIgDpLF5E1UnX9fmqH+2JPsGw2rLyc3L5LiTIMbx3JSvalwYwFa9WKUEuzDVuaMcdM4I
ptbyx7iR/olgxKvS7V4PoBinUnEc1nld/j7s80F2W8mYzWpVvX2UC2+AbIgbBAhN36TMLcX6JakM
BKkR0utJNjKap+qxFrxAMka6w3zm0qIwiqEQOgZ4T03EgveK81zwaUNnstHByjruABj9bhcBmwWn
TAIxlI5wBNjpUkv5UX3uAXu1hQiZ6WQeCxMhTr2NBgG03vdlbub7R7IdvdQxQm+8UUpbc9hDpUj9
ddgnOq3BbO6G3u7oHzoMl0UAFhhJgF2RBJo1z1pZqB/b+QMiiBB2FkZcT3lyR/CcP+/YxuZY+3aR
fILFqupfi+PwBlf/rsy1TbHeI5U8Huxke5nPeEmJmCJnTj8OqQ5SkgJy0e6UkkT4yjznNr3qw3bJ
1hiBB5wIt3yivW4QnaWh7u8EkyS5DV43AkMjt6v0YV45xJevrZQjT9jAdd6ZRTXcoWLynYqWuXW4
/TUAxlHfZhxGGtgQrxXhs+Y4fUxNdDEbwRgdGT8142ZEdxrU5TEahY0krsV6LOGuEzHwaGT3r9Jf
LtjZnGT5g9cg3GecqcpsP4BRHgjwcTdfWSm7WZWV7AvvcwShw/TxmO296x5JWU4ukJrYY60/8hrp
zS575c54OZ2PPZCpL1T/LJUszBWFKedvDQibFkux79kRDek5CgkeO7ffO8UhIBdx824hFs9EzcO3
PMQNyPVCxyhZbnQ6MhgPsBY5fpn7rqGZRlJdrv2+zb+ma/90dgEcjzZI55SuKwuZ8+4w6VmEg08W
C8INgTCG0rHm9sbKs+PUDJijfCUK93QXXRk20OAsRZ+jWENjm8789AnXF37FneQOGYoDH8ipTGoY
ZljPTe+qV/u7ihD5aKAUV65dK0iGbnLewH3/y4Zi4x15DZ81tjqvLHLQq9eECckHgGEi2ichjN0t
3r5u7mpo2ygDAxQZ8Ln/OzjBsAPLCP7/eQs4ZvJMTRaOV0hpECaetZ5QPvEXUU7ZKDMokIMR+IOw
4htKx7md6QCnWDqLsUQzI7zxHWQIjJmVGxqFUOGo2JStEsveDAsDMx/vjP4BNXpqOHXWI+j25OS4
+cq0US9VBBcMRCbyEkJFEFblk3Jb4UfeS0VkK43+in4Bn9BASljXDD5vEvwzbtzWDcnDpAIaQEvk
wQG7QBocZlw/Anf9amliMXf4ltck+LyEETQowtGT0yDsO4uQqY2d0qHkaX2cjxRT77tOpZItT17E
2XGgkYp5yiUgjW2AfJWoo/Zo69KDFsm1aGSewF9FWol91TYNP1mB/f72hH8hAQTwAzPy4Ybr7wzW
ohb6PwEhMBAoiPA5hBU6fhhXWCwWJFVDIRTRl08XAjTTTWv2e/x8RcloUssa3b/kkMQwPUUvtXbK
qO+IfTTBZP4YCLUwbHbKvISupn/zCUPRarg0TQBqblTYnbHInZ1JUX4YsntgL5RNsDm/ha96uq+Y
CsX+ErgQ8NwF9Pi3tknidsbhuuY1Wv4AbIo0PhcZrPMj4U3AlmXZPpu24CxSHuuRthUNISAxWYLR
pwX10QwTIo06wasvRifjm0EpWiBZRYY7/ZB+JS8TCaQ4ntWH3BxJ6MrdMYzxZrOEoUyjtwcwqz6M
cs7MvP8+zGL7183q6KNteIJE8DGA/nqZUZpkf9r+xSw9oYOQiY3yQgrApFxOTqVQKMQIm5WCx8K0
vTdMRS5WELifWL7ebE8FqhnW+0LPO5yAqjg8ZLlSfFb6rMBBxgUmx9JgL8sZTFaAWqsvChRwoqCC
BtMG/pJIEBSqWg36duweRQOv1SXzXze0jKftBN3iTCMpk7JWx8suPt4SVkjI994MysVTZ/42K4md
yT1P5Z/DJmla7LyQn2dwqsKMlf+JmyLr+p245/Ft+lO0VjEYtV8AvRLvj/2OVTv4M8ssyIoZDl8Q
eQNb8ZE4ADMnErnwnKBXgPf4G2Laq3eMTHTxE7f62inbKn4U5rpCi57n4XFmmARLjZuQISb1nyii
bimxmGG6E3w+X8xIayOM1AwNk08ms3yvPBXOfq7DJw8bZpNPIwVXAOBqmhgstGXF3eph6U0GpISW
wjxKUaC/a4aIl4HcxbDR+m7hMwAKDjZ2Z0qSSvlmLwR7KsduPtBNg0nc2xtDIdc2+I2uT1e/nru7
p7FSNkaWaMFY/ijAK7vrqH3Wq9XWlndDXBLq6c68v2RTImCXQthsZvHcTCar17q8ieAf0Wid2jQR
ot5DZXo8MhmkOnuwK4d5l1TXstpaDZ+ZcG6DkXh3TwTycaywWhyALZU6Xcq+IkQamT/P8WUtEjh5
qfrh3XAMNbW49NtoZ4BnPQh8aDiy/gEauhzTEKullOr3jdaUKDIah3f+ClnJ3MOwBnk9cFeezCzX
tXy7Fr0lqso/EusNy2/eWBn+rYq9WXVxyI9KlwFfu3hftmUN6hJDE4I4wBpx2jNzCoyVT/Fh/x7D
5cBp+n96Kz5bC+iM85HkOB0in95ebWo9mzksVrlLH7FD7DrYGIKthWWji00jfLuafJCYc2b/FxFU
Xd2HGnO1uyUw26qQ/0WtO+xLyvHMTEi6r3SKwvEpt53mbpcARHbj8W+Ukrd/hgNNDa0rP1lTd3Np
36SOsOpD01JikqCuwS1b/b+91IatiYbWJiRH2Tkq0/2RAtMhZVc706XrVwAC+Bk2saa1cetwkLZv
iUcnkA1yIOyYiV6Tzpeabz8Lq666YSCilO6JT5laFRQsEgjRf/zh1KqMGZi/bJwcpy+oll8F1gWX
qojsrj9YZgoXSfyf8WIGlMbas5MTo/C+XGfYAUrcsD+Wtn6Pvj4d48Go5nRzKwOmJ05P/UItdn9y
yxkWsqMctvBAREDhPUP3sbXwp7vHDky3wWcifnYCYeXtAPTD/bbY8gYZPDUOZGukkD7zgq8+ha11
PW2LA3dVDnxf5D6BhuvX3fUTNGOvv7J6G3csyOtHURdj29Ubv8zIYNaMF2PSiPGIsoTey62sRAF4
/RSXkuadnU+iFhoR4pqWmYX7j2W2zYzrm/gywXHVKBtzwblr3nDGYg6DzRXZiQ5B+ASclqsjirV3
3P4S6suwfF0rasZnUu8ovQvwpawjG+k8pFBDu5OmPUJzGcWvVZXawNBPEpeReuf+50ejyeVE+U01
boFL/8WjuzYXK6pma0GecRfyjnEu081pgoikkMVKSH2rplpWLb4oZv8D9J3jZuwTCTamxpFDKEJY
9V4PzzphlBUgNoglwek5go6DqA0POWe/AYEU2jeD1JdNaRjLgUrE0ZdK8fd+OceGuKX5lNRiPnHf
Fvp6PXTPKk4qeypEV8LQbZlORS7Mugr21FB2F6FgnxhdRz4n7L8JuMnlf+yqmRjyRewlkk4kVH7c
d3GWkG63V+7w3eaf4w1eiwyAAvW+gExX1+MDxSuNXyIG8KsQmNU4yjjJc99OSim2zF6ilte5vkBC
Y/HHqDQ56oCey7S3+bm85zGZzAsDbFEIZT6Stz0dcQz1wbETfEI+YR7aQA6mSCzqcCsfEoTQRGYC
AD4pdV6wxffCX4lf15qea3w6GkV4kuBeyeU0FipaMewUoNJ/w+NJljc5vspPBWK1BsqaHYZohZMC
NBRa4FeZDIXfCarqwzAhQ2brA9m7IcDCGKhr9zvBq2aQxL1/ryd97eBKKabDFGTS3LDh+F8hlIBr
MohiNaBDqpSHTtTc1PWWLRtNfAko84pUu4pjhMgtSKTUSU7E6nlo98eLyD+WkTr9ErqjkCv9+7AO
avrhYWr+7pLZCWauxpbuYzos/3orLSBGhdUeACQvA8k5KLZFIjeCOE5ddaEoJ37ZzGVTZ/09ly7P
XwO399o/Ga4+hdJ3GNb4XT57RiQ9Q6FNqzapwh3VOWm9KxLy0XhxHIXnZ7g0DC8E0QSvU962VVz0
mvn0YKm8jyWszYSc+sUG+DLRuUspaSnRTl9goq92e2ECFp4n1maxSUo1Er1y/L6V3UhlRKXZVjfx
aJZyKici5UyIpaiUdSMFoVOYvS3c/fOMmCm9tn6iQh5xLeQEUWIbCKeSyUAcCg5T4KemAB7YbnwC
U++393fy1NAwgtwO5XRcG1IRS2EoitnfpOeuQhk7A5AFSaIZpv7UFyY9zLrJU+Tmvxhn11JCNdCh
TnipF+sZMcpd6YGuQnZVRNO6EAN1RCmJlxRHh1P9VcR54eB1LjL4mMmoK/y9LkiDLyhBi9JIKExH
9Tci6en1rWIqDM/J8KMvwnNhc6fYoZEP0DYYMgSGY1pPIdh6HFs939wGbBWkueZ+YQE0wDBm5YYJ
cMeCBawumPBEjnyF3IeP9Xc52y7ssUopMPEUgogO2CL1SoXHLR6B0xaUvNxyislNNeBdoRenT+uV
8lBikD5+kI7Kdk6KoaERyQqoe6GHOtGAk3F32cg0/m9PleE4FzSUT7y7hwR1MPTiPSi6GWBUHrE4
MHFaW6Vx6/i3kwe31OXMS5dpujZca6Vem8+rZD8P/61WjzfKuZcRIgb+XQQE7mex/mK49jPd0Dj/
L/PLolGTJEw5XREWGXWrRzYoj0FPuSxqBfQ7FkRrl7gHF6msDtaqsDTIeOLNL7wGjWdZs1ywMntX
0yiL/eb7nColnAeqFJipdUWjMPafv8jU9xDmkyL+6xmAKcO2ec1CrmzFdClgLQJpU5KPSJItusO+
Qv8MQ5B8UK4D25yj5YwaIb4f3wUWPkdcHfO4TLY7T6u3YAsEYL9oBgxaKg6QQ+jih1+TIwdTRQiO
lR7fWw2n9pTAuE0joRHCT7ZdLbU3hf0+DzSC4bwkOmlAOpF/rCfWfsFFo755yDWUZJRNR2eNsrLV
L/uasFXTi9cK2UDkkBfqnXp5/KPOuYAhqdMXJFOM8SnrEHDB5QRLmaOxV535bOFN9jHOrcM0kh03
rSqJF5Q4j0cWp29XddRDHr+UFtvK7W7eFhIgx6BRyowX2MJ4bFKFfO98rRiPX9To+WF9fDXXmU2E
D8REWS2jUU0IBtK4jddu8lVlEOqpa6QgwtFJn4Y6JbcXabUAQ2F8rJgLR+X5hJYUfHmfeOsPzlEt
e2ynUsfc+XWgLaunPfQfTOs3VzQittbn7FZgiPGmJMwAaL3VRo9nN8s1Ki8zMHUrwHPREqyRediQ
JJjPPBDbWhycSw3/8TqneJEcfOi7Il15Ykvfw1mcQygSAlY1ZudxXwJ4tkt4ANeHLZ8pUqeUkpak
0T6SRR8JfNPL6UNWJdvXox1G4pxG14rjjG37V5CMOrmOEkZFGMJmSnTEdTYmCkfrjsKj0pEWqXbh
ltANLhvs9Y06tTS+DmRFNZ3++jMdh19xR5k+yszQ+RpdtTpQbf92JssT3lSci1hwrx7gbM5P549L
8aoeIODD7B2drmmuiShmJ5vNdol+luasmeRYIHhPnkuV1n3GgMVbFOX+e471TenhHRsJVsgnSf4E
vAubCt43zfbYZqblKT0pPt27cATMrf3w9hSYTNkV1f/CmiXsDUCmn0JGutuc7pKNReW/JuMSsvPL
MXIstrNbzv+OKjJh/TK5UIo0it8SpTg3awEmOW8imt/aWAAQaEjn4iQvDk4D8s8jDHx3A3/P0bc9
ukZPZcXny4dkaOAo4rw1oNPhCrzYeJkb6QRDUiPbag/bLzAHsT0yIv3uyHUVAWPiw6c6uxaaHJDC
HyG6QEv2cBIfv22Il2AQtoK504YGVbmviVVXOYy+CfMWj/w0HSKtJMXeDJ57VMBpvbTxGeBXXdCN
REsLIW+3pCYqNhvsZAFhkasvNlA7i8x5D9/JDvLy2E2tjwnds04N4iEPWRkFYFWFsJsZ5TOW5Dkc
ccILeqmEshRiloMxkZ9kkhW4IBJe0Oqj7HW19d2T0OWS8bQhvrCEtL9/9ggggdfm5LQ+f6v7Awcg
aRHpM2+4bXlW7S0TnKwGGswJ0KYUo5vhi/YbHEoWQlbpwT+9Zjh+2jnO+GusQU+tW63kMB2bJbOs
31x8pvHBXKV/z031/5kyjR6Q904kEgsfsTtwgTYKra/E17oMb81t13Qf4d2uwyAff7aLiF4nb/Nz
ycLJc17q4VFKTrGunySOeUsHNfORiKTqu/l5SPr+Wl3eZJ6cGr7YrZTZOJ8EH1yqdYg7sXC4yHu4
N/tOcBlZQcFPFd8WBaxOCzZxvyriLHmsGqLeQMdOOlFymYFVtEJxD8it3/4Sbop2yscRa9dYgQng
VD3Mamrd+EvqHpXbFfQz88Yj5hB21i3IUWQPI+5h+tO/EadOKCBQAUAeOcmObOyN3ywgepNymXOQ
NiU4GAy3qczZad0B/YpCOYjbFk9H5uitL4z6IHtTj7TuFz2PuqNDFDBJzA812eml3wf/M4BRpFNC
IvyPmbZFRmUME/fVd4HXvYCUyiN9p5O++EtBg/wsCP88YTpiKdq2NJfIMSuRS/gmKxsSVGQ79U/k
0kQmQwh0urkZF4fxVpp1YwZ+QEpBP1PSFlvWSU3D9aw95+IJ++TfuFH6jsH/UnR0XDJpKC8TsFVK
wZBiTftPOaJ46qNEnyCnRawomwdQjYCZbfFcfypkoNsT7eeQOZNOMDqzhz6b1L+rQnJXA7RwV29n
4Nyx7UVFADv6yOIqvTcQeXldXr4q4NhMhrBiHgwfpgImfcAAAHpKmaKVJc489QeaJof7ffnxdDei
ZZpx2LX4pRo8QEuAA+hNZyBOtRxMODurzOKhVlsSekoT8eMibUfMlz/ItFIYIryEq+550DxGgGLW
KreVvnxZprwtdMjKtrpSexxPpw/FmSJ+Cp8wwzq7GCAJFhqBzcXriqS4T1xza01ZlPibfJOylLic
UpR0fR6QzmGPX8asBv1Q0AqabEf+vy4gx9n3Rs3CtNpz3srh8L2VcDUuDL76+EpIMcGAGygAVVjb
Ssayfryhk5re09cpfvzjoAZsXNpJWfbuBoCXKQmfbj1uJjNOBzHfTTYrBM0aowTzJwuXS4/HuW2c
Bv2Lf6rBrOqATt4MLdeWq46rS+htXdFaR0e+y7+d1xB3LD+XFUnfx8iJeZ3+3bWMdTgxnp4GeXcV
UColtPmattYPXfyv7XMRu+Slgnxh2/5GLkQJ34q0iA+BmqBMfTah2fxT/RW5XepO0iY0Cpuxm39c
poaxvgQVeZSdchAiYU6qaMbDg2UX10YytFlq2WQ8nxcEf75FckZa8ErNnEOOyjvuPPkU56tOvRlA
K59qsFf7pr2lJvWSRHeAxgTmCfl3NXVKLLiU22oUbc1ETZiMvh1kdnVGKs5aiaTIzkb8s67xYqPZ
aOV7R5rE01J38SQ4F3aqk459ruDL5qrVSprsHOh978iaGqe3Uy/NABLgpPOvoNZiVsyf6hH7Ru13
9YfJmcMMdVAXsHIqkI4ntlmZGJ71st2HFcnfvVKN3M1aABI4GQdVNIns3hW46XK8vxy7KWgVkODe
MzVmefJOmDwZ+5pigGnIvIRvyuaYbzh/f3F4HrqEHtPpJujqKjQHgxJ5FG/7pcEzvDxdxZ5CG0Vf
94/DRzjsZ3i+kfY5wbQ818bQQyEoDd5+y8tTRAb0SIy6HAsizjPm2UneUyqdftmg95rHrSjGwRWu
Bk+9SYndelX6BFpbfiVNQBYjtna08qNz8ESGEQGYZEbFd2EmO4F6AJ0YMXKHaBvUWuYQTJpTWAxZ
mAEIkFQxyXJfHJMITHB87P3DbjfB7EjWYHr+OETsRbeGRH3EVIfh0NX3eGkpQuKwl+mQd48rX3Ab
3//NYet8y37qQqjcEQ8hrD49qBhSFMeZ8+NhKUPnRaQ/OS6Mb78cjxDKTsScLcjBiuk+j8HhQPs1
yuiFtV/1+8lWmrR9DoJ4cBFfmqIToNgptsiTR5Zu2u8Z1jdTnJruhG3RsowaGM8+IjYMmQl7B0Kq
jRvG6ck5CYt41rzOrCoeFUBaeds3E9VK3UHYC0iS22/EoGJDy6GkvCcZqIRZtsjbgbvBGO0+tqFx
+pjC0nd8NEJ03Ux23aTobG4F5E+Gjj40kZ+jdtdIqfEGL2Bw/Uobrm/bEKcrmbw4Sq4EUiZi3RK6
zV0c9mhz2dQCxranaBhZ+XGrJTSF06fr8G/5X32xHfk/DKr13O9QylC9tvjpcCBgB3SUaHvrc9cF
33ttTWiF2NAX3gZLqG1wEaQaXDx2LOGv4gKzdH2+EQU67FnkI7q0biw/pQtShDLoUL+dnc5+AyRn
AC3e71IBTut0cXHlec0Ts3E9VgHFavSLcBJNYqOAu05Dm8cyHGrBaWqpu+WVfXmidYluWXEEqPAX
uKgSUiPKswTq/KnqoQ1Rqr3nRheqPuVRwMHIcV8eH4sZl5T0XSgnJ0k2oN3iyLls2TxG3DBaOrax
X3xuC9iUCWIL09k+C10SlovWzYXc7IocTp1NypzEnrjA4Fan8D4Rk3Zrfs6rYzpZZGkUyG3VnHJP
i8BgqypKQ/Pmtgg+t5k+RoKGwb6ROQa00Mq7tFUv1huPi2zunOnxkRo8Bu2B+e6Y7lmzTHztD2qf
3UOQ9QldwMxy+hSY2ADbOnc03W1epsm8/3jjZnG9AnaDpt/wux4FYWu4bVyWAeYrqLS4lICCS4X+
qHzGxtLdvtWxryN83Z+TiuZwmBp6ug2qYpVJmEkACWOv5AiRCX9kq1DmuGH/ppmqiCUgF+M2fN85
y3bvArcbzW7/05RMlBETLCwnDEtvEMs/bQp+BR7aRAYp5wEgV1wjB4oPSesniVDS11lCg6v4lwPR
ZCBZUeNqadJSpkgVtkPmc+LqzoYgs6sRgh8sAbFpuGKeCmFz9wG6otWqUlU0a12GljtBSdgDcrWY
0NqiODP61qV7gdCqfY5Nb59LFCmXoQkiX6H68/MYwtfH+t+VPzy2VBiWO3EI58vpR++JMog+fFns
+lnZpMaqvYHpBooSdz2hl79Zug1KKEOmZMfCMUiRLdzWZaoYr/QVyD3XXhaGQPC0sp08JX6ZAi0i
sZ4//hchc7/OOOtW9SXCbnZcIB8eFLVX4FOcroFpI6M8TkhgevdFAq0nnL7eNfWbVseXNbbwQSzt
E3vzjGULG7THSPYN1oHcJfinkUe1vNk4i/MmA0Tt3AdG5vBIb6LtOLxIIQpA4gTQbx1Y6oydy9+K
Ms/RLxtAFj0MIiPLB0gQLRlcpJiyP0OeNTppLGOMt3z/fc7dX2vC66E9GdP0dE3RsqnC1zU0hqvs
3KMskU7vhclP8u5X3cmmTEZQXTMsGXrsqrvSANCJp2WeoBT2/7F10g8a7ZFBALBfnC8VzYi8o94O
pCHuzCdx8hJrw+0mZpQEEtp/CNCJYhay91XYrjDpLKcOuzK2aTIdd3lp6idMfAGBIOUKaoh2e3S8
fTqNFuxYC7YOmIutsmEbmuvWKK/7Ik/H/tOf33xb2j4ZF0o9zzFOeZOXFXyW4biY9lPItIQQG2F0
+DSDuyNsGGKzir8MDie66m5G0J4S8YDrvvOFlASbi2BeRkIHUk+C+Gp6McLZTht1nlie9jGrHHVB
ClZqAXQsIONWs3JYgIkHaH1WB4iZGt5GqrzV+2RrFCIxaDzav5vuZjsNanUlo8xIWXsfewmCFP6y
NiCIYghjTNVEO0ul8TNGV61MvMFEl4plhKpCX9Sj829EbRRSOOwHRxKfAjmY++M8bXG8FyiEGfGH
FIUMORp3M9J2Eu2GaCUmea5fNrn60te8X2PBjmP6BhOb5VjoQa39IkM+EGg+dnqA8lJr8pMRe3Hp
s7VBqRNiOnB1DvmsazPYTlZumFZDZs1kioAZt2NpDgCGq+LFGsPt5gfGh36RvNe+YihSI0gj2STS
9Vu1XWGxXQxtii/BZZ5haAcvnyfaXyL67eTMcB+eI2BCUOAFH27PYbisRakN5LFiBZNQGqCOMfh7
Tb7RDR8sYuX28xjxM1DSQKGIZheq71DN9A3j3IGJMqKVQlN9UT8FmKIUr27yf7VGlJfowenWDEg1
IhTUcEKP2xcWgSmau7goluH82zWik0o8Ie/0jy+i34dHqiYTfZFVQ9sAEnS5Y0Yv0lHytacJTguL
7sj7gN1RxP9GqQfAfJn1uunVbSKenoVl7Gr7Mik3JwEzEJur/8HjC9NJ9oyegUxKLFFeQyQ9o89l
I7ufrqF0cgW8bgyiCnyvk/z2w5UCkNZbeEOhh21alEXJO/8PbLcOzKQzdbMTZ43H4Pj99PH6K2eb
g8NYCiMbq1uWF6PEnxXjFTlfYl0HFWS3kx4qc7Y4pE7Wwm0tGS/pEkp441TP7fbt7tC+bf6Cyxb7
4k4Zwm+qLqat2Ux4LATk4gYJbKczYUG0OP4vgsy1/osHeWAnsvX4i+gXT9Si2NIOGkbk68gKEHen
oeU4s2fQFA3zCr86x0f+OumX10PDGVVGGlMhDVsSEIIPenQqNdMrIOXmJJqnOambCZie4qbUu2Z8
I5qVZEeg0XjIFt/PAmxGu2BVnOBbyQWKZPykjK1eX5JtGwruTCiZ22u5xRAl/wI4DSEHIS0lby1t
aZHijAu0RvVS/KgcJN26J1Aw7AzdyTe49qiIjA6QUF35zgFkmAb3rftCorXX8m2oUsY9xniw6b/P
Zf9+SsA9Qt0V5AhYIJFr5SHetxc1O3+YGtqvXYYoQ+GYcBrdmrbNrih/NKlTBtK1a5Np7a2dZwmI
abJghB2EFZ8nrtqX6TIDH+6/4ri73bkq9JHwi9yK6mfSQ4q+01LlrtQZGsWiVz0uC+X2JAaMjsrv
Uhr2NTyCssD6a3AdTCXviHGmko1UK5L8aJG/KBhMrWN2QzkS6LeOaSzS1fPwFZdMZQSl7RM4DKmJ
IzrpKUD78klKgBYmuZxxj2Xo232RHv7IXXb22kFgHKyxJwun1ZNAMlEuTLhXjAioIXqCTpKFUBzF
vmxmShjUJfBtRo/RZdnWQLB4OpZqDP3z0tdqGi3tBfUJUggeXWv6fgQMEjKTuZjXinK0pN3hQKB+
/PQpZO+yyo8ppWZ3X6sy+opHRqGiBcOGTZRjX0OvaA+pkrnC6I/EJtth3gZQh4dXv5mZ/4r9Q+vf
/I26CWQvou4Iyk0xmKz4RtO2nIHqEJzk/p02xZZK7HEGdltDJrCZTId/gXh3ACw/iyQMS+nykUEy
u/YP1/CFWHvKDdniua9xPEdg/5frJQAkY/uKwO8JcCmOfv41vx/rPI2/5gIE26EUO55u2mM/RQol
ExvnCGO2XCxC+nBohSoAQA1vlPyaWZtLvvbp0uqLYFjZJe7j7BYbszCJ0cOY5ufgVmYNsuFZqiyw
OZgRcSbs48CK2E5sZYEpDoCzMskewP+hEJ1vLh1h7ghWaivBu972ToLyTS+9iZdOADklCqhaO5Lb
3EwzS1eyWkx85cDH6uSZOh0yk6GPS4/N97wlQRmQPJce2g8TDnLTU/sCvlh9OrF+mPCtVhQUnjgv
Mhnt78k8HVx9JZEFcYM3l8wpB6hDWDuFU6TESgeZ7yxEWcUdNIUjfGj8zDD4Nl89xKWCBmMMW5zi
/SfORZU+u27v/vOSzrGEl97zAWyyodQNm0NB+43LBYkvc17R6zdgOs0AwkdCjDJhhwDj8mxlcSXQ
LqpTe4ATXG7IIjh6geLVWUCJZ6SCrMONWM1BmBmD1zUO0iYRGqrr0eQPNbpE567HSL6TyT52nS/G
AgZO7zwJjhJvyuK3OwLKTB5W+YSoymlQgseZ5cEiNMVfx7A22fzkvbJO2mtExQCMdlaVleNeyZMF
4zQnAUuBvY2h2ammrkcu5VdPptBVUhq4syUzD6SlkOgpkCcXg96WVxl/AvaIh324H4cTrf1Bb9eC
0zM70eU/wDf6CUpmx6UUJcYrbSm6VBFITvZFOLoDWTsY33FJ8E+WNvx3g5DyrgjA2z8xhcI9sud+
q0sgByJuMPdJH7xsjg8EhfjOc/hPmCtvIfn1nk50mIeIiNz2L8s1xFC8vzXnPMSTIHE7dRHR9Q9O
TJIA4b6dE/UBkn9FHjqBRImFpfbLU5hvFCOIMzgRCWERRzUsJxlVlnyCnGJDlvI8BkoPWpoZW9Q6
7dJZCzNe/0i1ztnUb1JJis3R63gCmQ0KgUO1uFhCGR337utHxHGsptQ5KeiVnIiwhv1Jb7MoU0ED
Oq0TGoEradzCyeJ1a/4zQez24jgERxVl4Wxy/IuWLsfk+AUcTsR2yOXMIeJTEBnt2UXnrc8xVpJF
Ivhqmplf1999VjUZ10/dgi9Qt99N449XkGnmOCRKsySqRXDFyhJgXDOFyoSFso0EXdYLP1oXI/Ki
jqXovQWRRa88aYbA+HtZF+4QhO+pA2XtJOn4o+fuZC8I/y03vN/z1znPpqyETUd4rPrefSUEpj3m
H0fJI0wOVl4bEr+8xoA+xiGZ6tA7+VDG6L4XsBkwdCvEiCqhBafdBSchpngyyhbicBXAHNykbNMA
vYzXWq3+ha5YZYe9Lu0ZtH3YN6EQz/Ndi+QrM7w8470/zXunhP5Oos137yeLVZHGhmZ0F3k2qnBi
OpPdL8r4/p+4jtUHJkK+5s6MEG3/nv1g9zrgTfaK3MW+CGbV9oJofBCHWB2G9l1q8iPlrO3HeDTV
1u/45ipwqSorO9tzJmP3kx0bf8cR0Emjv5RrFVqpMYoaiCa2ZFCyyafarKR3Mg3st+XxLhCaLio5
6fIzdhz8i2T0jso7Tyv/iMm24hgjBeTNP/PxjYE2/V/rcZBSkFgcHwMaQOJKNaMd9GaqumBOaX3E
ALMYEbU/p40bpMhrf/KdbrUR4Ldbc+QXvNBuRcI2qNxBjxNfUmlUbiVr1ggXekb6B8oKJ8O8f2Qu
0RWNKmA1eAubkYw4WfkzWcIiTgBSAEyNM6frRTp8TE0z0VR0+AnNl/DGxcQumfKOpZx6NFg7+7Ov
wdAMIHMPUm2fNzENsuCKA7XrZV1dTzqwWQgp7F1HhD8nxewpbip1CwMSF9YtE3IQ4HIhB7A9VNaH
wMWy1epJrpMC8IOWa6b8gGcP8vZb1iGDWhKmsIkZFhFY7BFl4Fo7wSG7t1ouUy7OsOYgIQo116ep
ZZRTWh4PvzXcB9gMbxI8dIAkHRFdDoAL3drzExw3fX0pp3dWykdCQIUUztyvu3i66NLLP04lxUIE
q9CSvxTWNkxECbuufjOwegpXYSF999+shMH/PQFHCavvIWfgjIxmgwznf9mQATY48GN4FJyVSan/
j0VhWs93NIx2XWoD5yWkVyoO2iz56zoVp5aW+Gpz5ogZQ91ePg5qVbIf55afo3U0B48ZGb3gUSnF
gR9eeMKqZsuZpIpn9n1KLFZDWLPULt0tIbO9Wh5u9MUCg9lFZO2jNJwikR4kh6AB7/nE760Mb8wJ
GcGM36vS8UZyT30MUS0uOe/41aPNmW72v3nJQ1g7r2H6IqH6+1PAlDeZItcBn4IqDlqNXGLSZclt
ciurwGw9m597zFvxTzF7uK9eMhVY7U7F+LLFzsHLkiOGcCmgxWTLxxdyM5DMtmnGyTeh/C/FALOL
oEkxzUfZ5m17e0f20qq42mLeQl6k0dyLUIC6uTaENXhU2z/BWIFW1a01SxB1PAP8Mb+FYtFA7Aib
JfFGp2n/3VVxoXsAAHEoacwIg+rZbgbFJzD1Lk6izJZfB21Vdpqv3PyCzCDFI5Opm/w4KvKoBN1y
fchePsqjTvJRW4MJ4M3lB0MfcOVZegCWQ8brHwX2sEyqyN1UPHv4/8NpK8UX05sBVNAZ/bLfDkgH
JRDloxO7ULDmg1kl5eXRuuQhQQfDtiy2+s5lTQ4PUhHhp6wZ3j9jXasSBdiZxIDFiG0VQsAQ9yXk
mo/oHR7SyCuvucExI8NWI4LSr1v+8gNQS8XbsykuczhxlyJ4Y0FUUxbPIw5vMUlPLeLoLoMqU1lZ
4hujFc5LWr9wObaIUcm5k+01HM1L2RN2+/8I05UG9iZ3/gyqd96JPy3MdVWlK3kzIc3pYHD/uu5/
gzFcBV+4eo1z+l6xSk4nIvQ/5TjvZ2v8rmn8u7i36FZuUdFreh3PHnvrwmf5iXDmm6fr+nsWepS/
GnrUEjYDhuJc8dgZ4AqS4v2J+rrs20yqroFFv68u8RR034+RGY8mr4PmkH1j5RhOW2XiGLq9myD0
LpHY1YPHuj7V+l4+8RXtimJB6rjmi9J5GDUtBgGyKib5P8yzcHIOdY6mySTQPKNRYJCqTpmJ3vOt
FdPmKEOg6UVH2UsGpZoQyHvwm0gPESj9lLdTSTopbYuj5cuqEK6Iep+wrkSHVoe6RMnDx4oXjtRa
WBXaNLzcq/Jo1zAnbzc6jiXihfkd9BE5AZITLpR0HAzpf+xxPcgVLVzsJ/oSlb6WzHZB/vIEVY99
ofscXR+/W1dSkMBqpP8mtCdKN/DfG40n4yUa7a5IwTwbqCH86/5F/J2SsDRsQtNDKz3gT/LNzM2o
N19B/y91eDc6gHDlPvoXAeyRapKVlAu342tfPeBOBeMCzjceJu8nU5N26EkG2AVuDEN2Eh9PY7dM
jBSLk+QfOBQ7w5KPjjHs8H4OZQoA/guXaTRvUNgY+mi/lAsZN5UqXOxozDYKiPMIsJiJoponwhQ8
pDy59BNZuHPio6rdCaT73d6Z7HvP3O1zjBjYnlruDnOvlg+WiNoquXkMfxQjzfQjD6bmuVKELQZ0
7+cY1LkjQybJV4o6yEwih7oO8Iqb9IqYkfgRMxOFJin+VRBURRYB37G4IJTCc9ZD/9dJQOSEWU9L
eTbc9jBWpGGVVN8dirAdY2vdU7HI8e68MV2Jyy9c+ZVFre9g3psGDwa0ga+I+VReT8Esp/jTH5Kj
8UCyFkHBSbsuv6yt8DF9a9s48e9A1Hbketi7Rdag7YhqCfWa6cdEZqqkN+XmMj+etZGybb5Y4dQW
9VvAsn3WGCu/Vd9Wb8YsXYa/9rlFgu9b+k/bhKcw5ayQ+XkGpro33ms9lzdHAoyO5j6cqzv4dsCS
0h+GeCb4sjHVwMOvkYb9oYIUE1JCYXkz/FJt78iRlue1alBRUQ407JaApki5uQjNCf2XZNA1vcWP
q6TVi6ts0HNbqr1IkpzwjvW74v7gI2XttFJcGxUK12xahf+X+K5xEpJvoq+bHMUCLe0y0dHfbZ6K
LnpYxtvBSFzaYMpAUnI7qJCNDt/LKeS/qNah8fUsTKIVr/nSEoHtL1KiMXOknPonM5tKuaZ7GoKV
Su9QxeWMqG5Zx3MxShvlRQplcTeIXFBNwBWE0VWLxfXV3N6uN7Xj+u14gqSRYXsgHE/Io034GGCi
sCWzrmlgoLuNabY08hljX4LDaDa+ANPV0lmmu63eqVaCYT4SLDJYn2CKF4qy5mopwmhVYtHVDbm2
HAN9C4m7exVTdmV+wXxPeX8/DNoQ07RY7CiKSGDJf/5ITughGKgn5MyD7vzq4mQITb2BiEbyB0nF
4frCBYQKsW0eyDGemBo5TNBrfnmmgZejVLSV1dOSrpddfYZ1tEn4Nz4tv1iwC7FGs76xb2MTIBR1
7iVOZ06GVMTLcZLA1SL4/4+I2397VNSSIjgJE7783dwkJmp20TYb+xt8r0QDjJGFzDDrfLwwPo4O
jJxAE/Xk8orrE4bm29IuQKlka7dLbABH7JK9uRuMqQx79pS8JjukoFYDUIsifXB3n1KovTmAxrVD
x7bTn2Q4e2pBNBRHOlQoWtH5B+oELxAm7rcN6qvSfDZxbylp92WZvkVT8PEhPcOjjA4fhjWTqhMD
iZcD72wgmsyjTzH5DfEt8K5AhFyd4ga32cFM0KlfclX04dn7vH0zyILte03xn3yBFsp+S8Ki7eT9
O0ocMQ2q2UNi7fQi5vXdw2YAjHfTWF4SEBV6nm5a92mpbRoXqZFm/ATQXgPR4mgH+R55lG7Xhhxd
rmP8ATeWc9krWKcvaCnvyQiDuPQYYoGYC7Pk9kPrMdo8spLf++MBtxhxGEhR6D1iPsHMNePkiic3
HkRMcdxh38UL80a8aOyNDzI0EriVJCAYOryIUIz4ml+BHIpFr4ifV2WW2pbneTOX6kOQv6oWhhkG
pABpK9/qXidb0qjU0NTk5V3hl5WOo15W1p6ftCUKQzaduVZdXvi2xGgTQ7DNj/Gv7ChlLnTR9NHE
VscJHJDCkF5GKZUZuI4ZX/ytV6dYVXykCSeDuSOJYQDbcZvNifZb4iTDDRu0j72yLBuu348cnfxF
zjo4J6zI2A8TwcRfdR9gEouoqX6g2xi2hz2YzWhIfn9plYOQ1TxhUzlvEWuJtyZHAmlG7FqLZFcm
T6opmL0gb8QCeEc2Pt9bh1LQUqgVeXNsm4ypYN5SfSY87Ms6i6LDv6JqtbRk8qUt4tST/KBfAoDT
beXel2n5pb3raEnridSNVVV++HUNV7hcVj24LfuH+arlW7OE5ZR65ncq1xyhmgU/xE17Dc4Bjp2c
8Au6XTtyBb8434LgqUY7x3Sxm8U0cE1aMSClWCFNv+G6WVQiIbSPBZlSu7KIylHTqnxhighXORns
vcm/QVBaNeLC99Qe1mWKCG0FN1an8vsNDI3EVkyfTJZSe0/pjow8dpb5vVSA18yDYNz0wjAHQImB
5i37pZ2kpLSr3fJjbT2M1u+DMuOpLDuBiMQCv0tu8pkxUc3kWo5ihDi4mnC7U9cO2dVRLWdINBVy
KrnA7HGY3TnCggsTzTgCLSMacJEC/tbYpF46Bm416+LBfSn0D6kgueTYwNLkvvNemZqy8DBLZr1P
ODWAv9NCoRr17lbVQ1QmyYzE0ytU+Ecd9qpNDILnmzXrwaiIaDn3v4eeaWyxSCx4g/lvxSX6ue7R
42a/6SzS/HaE/mZVnAdM26fwOx3LWG8qTHleKsVOLGDdf6pNKoUNYp4nuK0FmOeE7J9vYHdHOwC0
u0sjRZltgF+TsFaVn4e3D27WmdBXGfGsXhrwiVhLJ+VndJUh/xoGrELtlPTFsHwixpxmGHZ9XtrP
iD2xWndYlFoBR75BT0wERWjhkd0thl+XOsLNntyUl3Hla4bB9h2Khh95zryVZfMrXXhVVEBoaEW3
KIh8kW8Vg8aWjVLz8Ra7MkWNwUqn69Oy2rXjf2AJknyyGeKl97yw0P5t0Bq8GvAul1hdmq+Y3bIN
htfstcCMQOzishh6Ub/AUnRHCN2+4RkV6UIM2OVx72QeIzqachAj0FDPhwCBv5y8GANPRWvnBMBe
t9F8FHHPDobczn5O3+GKF8zV/F8B0l/VqPqS9kjuogTRMlzkv0I6A123QQm+ufxhAK8zYl/ibK5C
CyjZEXLo74RSXuZHX1X5AT8LpwCbHT+ES4BsYsMmZ/bHHSzIyXnAha6A0jvkT5UxbnjhkKA12aHO
0rhOzt6QdeEE/KDyANRtRLUSOl+xSxozupfQdrFAMUi0qOzX+gkQ46Al6q4GdCoyWfsHPRYLF55H
j4fBxhDDfnVjjWyVzvEZcuuTNes7X/jsvI+ByhrHhm4WCP0Srrk0FEOxEMtHfbiihClWsZmCKY9j
llLvYet7JNflQhu+CrdS/edXU+ea/XiERv9iDZEd61S6mQadiU8VVYKDrNBHLNb3QezQ0vBplO8u
yElUqvzhfkMwIb+7hjzgscZMm54wonSsM2mgsZ/bGTkTuOSnYqCsYNgjvWOywGtzZb6GUHIwSCew
ocpHD06x0GgVk6ftv8HtpubiEltTac+tBSpBe0cBszJordlRl3FSb8ZUkundF4rwmQY6gIgtOuCc
3FmeevsIf2C5Bab5cSWWTFLTs40j5QfvNUITW3+wZU/PQxPwB82UF54fhPJPxppF0c5P5wDcVSNC
5Uw1L7+Zq0iow5FsJusPCL6GTMBmfAorUB6T+UmLhZWnpNQDQemY6DVY6iqRs1jyargQN8YDsJkL
AXqr7domevBAneLWYdADzpDU4hPvifviFvFsWQ4yX8T9A1H7+ao/Z/UvpvpJ/4h/6C888dphqbt+
BCwMVzNlDenbIhSj4Rh5OGaG6iRlmuWMWSD9Q+jv0bFx7pS6SIPeNHSZJLJeimHYS/Yz9QLg49Tp
eCKoDKClM6Uzz26VkuKiTgLEKmMDhvAiylHT1778Tg1N90pVfvDLSsKlf7lCD22T/owiiYFmPy/x
TGhrvUxrAR0rjq4Uj5pjfb8PJF6cuFvzSrZVb24NxzHYqYudllODSdQJjqMjlklScjN7gPZ8xl/L
QoExxhAuPTCkqyzamRCFS5rMyTkGurXccIwxYQni6SPsY5+3nTo4sLzp7Minp6iq0mCCe0wd6mTu
KUE/OJJTO3moI9XjSNF0l0qVpgMXvFGDx/m8z+tjAvvmxZbfUq6Y+UvjWU21n4//JOAzxL6B7RkP
6JsC/Vt3XKdEEVWtyWCBtgEs5dpiwvJCuOvA6SNqVx+xuHQxwBRh/sjpIcWe3HP8t48AXGjFcU7q
eByUefW2LkaGde70/S/EuUxb+ujaFPZ1tjRRMgnQJG+6NbPQzb8kVoOPCBqTnZUfhWyfG8ccO45C
wuioWh4VMRRli0yU0hgHfNgzltvsWja6KYSr3rUC0tSFje0eUxaNTDRyA9y852dfG0GjB2fNdoxm
iW6C0ihz/+GiYZULgp6gnkfIqRPvGstkRXdCYu0/kx+Cu4oaZ5fDSqKV9xOnjRbHpcpoIiDnKm1w
zg3uHpCugr4py8uqdgAzGlYujijEBdunXevR9kKSlHljsybxoY5YyaSCyaeNyRZ+VM2VS5+DNXbH
tCDZq073ZHdJBVtPj8xM6mw4InikvHtBOsI2pDeiJzzHzB2+LR5b/MjPR287+HDIRfnA01S6H98u
kvFNeC7damTW0uYPj2I8kt9XLgSlHD/NmBbxeq+HnAHbTWTHbk+szkaMy9akmFXF/VXaD9F3Tkht
1ka2JLB5blxWd5QBoigO8CN9p+fJWTaCDEQpgKuHwHgRc1PeuKZumCCaoQzbI+SzAq9Pnb4A0fxp
6zTPDT6LaEKp0/X8q+oGaSjnb38DQO/miPSlnf2SonwmOztEJHb/fI1NTeJTHEEpJ4Oh9eqCARO5
VEwdjkUMfjXyLZ0GKdPQHkVhKYQ1Tr4MGeOmUM9YjWPf0463SRbeOQsMHxi6LKCzhzy0xiJFTrMO
dn2kw+As3bjWUCQos1BCsEIO67H5FBNVCVppgMoHPMMLM2vME7eNjumHoJ3Cy4C47/sOGAjZIwQH
e9uqQEaShzT6BiMLjRhszolIhhHaBl1esu1vx7a/ZSm/PnyiJ0Vdfyy1Jxu53KRZQm1qcrsvi+U+
PHFSR6SLZFY107FukGRY1mVCZay0ZymaoX+fg+mub2jBdggCmCmqkk6ijdohbyde7jV0/psKe8XW
itMq/P+OafqcZ1kzkXB4StIlc7D42UDib+8Z3FdesIB6+SF4hkj/g05Rj/Bz0scXAddwclgos36l
MtnUz857+NirVjGDL0D+yy0WrpngGcbzzL4iZDwxSljTnaMQzSIQjRtYSH2BOE0lysxm6kYdBAIE
Bm4796tfPLehji7VmqaNmruU7GOl2CcDZk4IV9y2EPZnJWw+D55LHNokx+jSq70FaZYm34Usdtjx
O1kCKLmlYBgtN3Mmaw5t15d93FeThr3fO8mTUs0KPi/+tcYs2XWAnubxwhgRoJR35QfUIpGFg8L+
Lg3wR3jLG5hxmXNAb9yXkOgggeMISe13492qETXfFxVMI9JicVWJknw/q4H7e0nmnMkd8eOPCDI0
cvMFi3NpkU0MaPf2huyUP0+3ZCDANhUi9BSgkAsEnvUQHpboqHz1kmQKkvQvtlSLoQo/8ITZ+ngJ
6EsAR6bE7bCavK4IoTZpeRQw3iCV56rYpVyLAYcDCdjdYFZZcU/L4sS+Jchd5x2bgBdGkqk2VA7E
X4olxLcs8Mt/IHCM9izFOSdBQxRCdzXLbHBapxoOciTYzpqfdqatEPC/gRgFWpJjPfCCeV4eU/74
2XvY5Kjpp5JbiDjFCK6JvVIwJjVQHcEsPxvaGt9d7xJhkGF6oVhiPvcgKOup+hMj9YPwZ9mDgXRW
2opAZXzHYo65av1ZCQ47Bt9yxibqjeHMzgX4LhqduU3B5JpvJIkEbce60EKTj3jiCTMaJGB0x9dp
ImHKB2/GUGMBfTjntppDXlnJxLXCYBSfxVkoKPLbvFEG21DNiqUUFbeKLJFXhKvZhgB2LLcSOk0p
6/zmUtbpBDMMkTapJuyZRLsqKWmzNO7zfS+uIaCdIvR9hp+ancV2vtQg7Lia5ITfTzy+8a8S8fIS
yAWXznPHsPVbT20daif/dLy95giv2s13MNMvrUODpyeZ+RYdjLqyGbQBEOpLmKc05bS7pkk3aApX
rK9Xjgftl337/sJV5qXpd5GCnMMAxnv5c6wi6S36Jcr5fIm4e4bsgG+Ud/p1YKo8pvmtOLxRHVri
bf/pOHCA88mxy8Anb+KrAo5ObmccoqhjwOHD0EH9W9zIbTR7Yx66PHdQcxXaKpEuYUnsVwjYQ1Wt
1/eIAYklFKJxHWGoM6ADe0y8k7rlcJQcvMGQnDPr2+C2enYH2u1fK19SpmZiXzpSqhQuKCSun0at
bqTm8bP5vUMaveT0miGGXttI6RKhioNVvAwuHnGnntqj09m0UBeyMzdo+aQdos6BdkL61IA9R0+p
UVlyOX26Mp6fiskomEfBWozDQmsfgLWAklQ1xw7Oin7oHLYUW8Pc4iLA5fkgazyembpApLFHjD7i
ViVLspSJj3VP5Fh7OrgEZHtPWoApOkb+WcCiwU60DA50tgynVlSar6V5sfubvjLOZqK9Ct/1FeBV
qNGWQxbczdTBUFbqFM/T71N7S75EdCGfMixcGG1tij7YXFYt6+HACi4rqsUod2gJKHwimRqU3S9b
/go2t7+/S0xxj50iI/B3Xng8fntOVZEgxc4SSb77DzSsz4L9TLlUPh2f42TmFhFRpDh5AapTmR3+
PRAerSebkXrd62fzSX25cwxP8SS+rR3NatDfBfbjV4u6hKCBHehH7eP+WhKWcet9gmOyeYnM5EE9
2xHqm8QrX2/sd4RXd4lG+TtcNzr0Kod0Pps5PIEv9A0I9fbltxPpMvdRfFCFiN4RJ9SE3Afg/riz
SqIingI8bFrKmZibyZitJT+9LOPWwgiEnkv9EdIOtFW2kbnnEoQvHwXlk0MH/qRsCeEHxQ/WxzJJ
92Dfmvr0P05et0jCvAR7OgCkH2xS9XyoAkIwdqsloDYhQ6jTHS0R+X677BzfRidcVZ+pULASyZ/f
d5t3SFgIlXq1voNwpQVjSMp7udQbwYO5uzQt8oRysuTs376pVAa39/EqGVk4q8OAS3PEMfGEajBV
87qH2Kb+jmAyutxr/MGYSiRKUQTWKgfD8Enp11BgaohVDnzJhN73w/2cWG5ibQ72yINjR8QgtZgs
MrNz9/HN6Cd1kMTz2EymvrY4zEEIHTATF6TQeR8s8QhVzTr11ctFvD+Rm87Z2EadF5i8t0C3p3gM
CxXy+T9rkpfBUJmgizCfuKhR40CVshmeFh0U2JSQjYkMD9NyL/SMSMW921RM3ojJLkIAOaktPD8a
5NBsXQqAAm95cgKiNJT8YwZriyqhV5pTXo4ZGJ+uCahEBwgichwoYjf6XltT0kk2sE18qQUyWlK8
JzfxaABwhAafneFXL3/aj4ydcVH0LyVq5fFumf5kvYWFsMN2SfrhYummNDyaSEpF208WxbKZjyfh
Agcn4epRJkdk13R7aY2OaD+qP5MJ1tumhlxA0jyKocdbD7QMrYQRQIF0kcmu+q/5z5XtdotRL79S
qZh9i6lmma2ynhk22z6a/V7OQ0cHIEsgttE33xq3F9tvDGffpRMVtiODM2HzJgJPHVetlSBz83l5
gsxIvjYOZN684zKLUnBYSOsFgTOLCRziUiJEsrfdAe/Yx2vq/GBnslRWUhXFGR+qpqzEZDX3uhgz
emcbTfz2+eHD082MSoPtFBGpedhPaDprZrMtHwqB51g+GwsI8RtoNYCn9Q7d2XcGgDzy+gNKaSnc
66yp3wqsszAldBDLYO+2oF5gTpuLhgnhFIlEuPDPV3XFEdht6T8EPXt+1TteCRWf9rcCgObFrsSM
yrvXa2b8JoAj3kMwQ1mzKJXvysY+Yq6GD9XmVAFatlVj0NWIBujtapYtIvnyVi+QsgdiReUKzHEu
q4RHFEoI3RerPh9WfehsfTXXYT9mZ8KMImQS1OXET5h2GmX4s0f6VuXDLi10iMyukROH4ZoanHmK
vDH32by2aP5efRkEeNSiQq5Y1ggyqtRwcOlvrfFDLoPFu6skWR8DP6U3VdJvuFnaTy0yc4h3wiGq
/uyWEQ63MDQw8V/XV911KmQkyf7psdApRS3jnwacL+uCxiwVc+vPd5ITTPIHmQ5v3GpgEC9fBq+4
cZRqpVFvx2omStdnGDPLZtQj8fiDG+eNB0egXvWPQ3trbpsmjlpr6X4vWfQ1Rk2SS75u+dG3ZB9O
B7jtlqm8HzxzekIRO8x44amQDaLANd7+P1RdGxXwQT3CDHtze3+x4Sm9o65FuYZkOxDh52M+W1IS
/JQPSOM3N+UO9FWirjxq58SVsbo+RiKj83cGcjwhCA6VFdgAQecxYU5Uqcwz6assdBHu8dhHSuxH
oZ6mljBt4DgZabCqO0DW2nGe+cIRoZwLNBF3telAIdTbbMGWtnhNNxel3eJfsk3sAAEI/KecQ7xt
s6zHfgPJm3T7QMZ9SbaxJRBVakji6NJwoMvAYYOT7LfWJ/NwUrz8oA5D6UExoWG7HG3OnmQkhfhS
cpqFAPQVZr5jQBp0BmYkGUO7I+77WWsYD4NXWujfiHChyBMgVL/XmhNHaLwbpqSl7u+KO69DyPHK
rRLXtCynqjyIEgOxDmQMRP9/Ws6qVUZOadssEFvGhMEEfNyy7GZlREdgoY3968Dcq7xKBrTTeWPY
2MNmqvRxLcu+fyGFu9G+jeBvM9n8YjV8KFV1zL4VKucCx4TtV8k3mcZ8gbWDXF2t2N0iEedN/i8G
Fu4X2q9pfAN/+WUNzs1A21jSwIY1RsqNvUGZ//yUHv3nHPVY5zFM6jb8FAhM/7I+q7fTBCoraJw5
hZONDVjWOHooijYWi6MerLlLK+ZAmnTyiBj36vXpq10FLKqOujp71JPW38z5pJYc5UOuZnlRVjLf
/kaVjwzhTpsZCMii+6wVPsu01TkimS0O7Dj+v/UegSSBmfPFAKQx04Cqy8lm1Mi0fJVFrngBhd6K
Wf3jugC7jApgideL3GfhTCLKDSabo73cGvMrfi+aWARWGOHjoeL0EX+/RxKwdfNAFbbBMW0LveKh
CVpg2j4szG3Q+v/IcL5JghXUGpgrmMo2oz3lNqE6WxVyr2zWZ54+T7o5du90vE3hfdrV+diG+rif
N3y6AGD3jRiIc/cQZxNPEzy9sgrjusokZ/jIQkt6fMvZaM2J4yvs+kjzYEuYG03oAdLqehLxbO0S
gS85LGrT7gcIwsV8nBmiSc7FJazv3uaU/LaxjAlAYKCeJwd3I0Z7HVLDId2GQdwmmAk/1u5Fmv2/
Rdah4X/JBbo16GZObfEtnXRCygAMeVMCRPtgv4CJyhEqEYEGgDeRR1TgP49rAuSJt5HTgC1l2eVt
OZeq+AoNyXDE5aYkairMlqBmUYQnLRiQtRkwGy/ftjezqGhFclAGljhuUsmVViijNtskM15gPwR4
et1+pMuJLH5POwLnRoz0F2Y5OsZrrEvRm/I8rahbcCG2s6R2fIcKD4aTnj3vrs3fx70EE7f0PLOC
YrAZ5moc6qKiXvN1hjHk/JA6ztR2wdsCg4oXpf8H4iOnuwxARWuDniwKgXWlgTOMBTQxo901XAF5
duaLzgF2HOg0E0+1b8Ks4dKvwMzcyd/5Du1zmhzCusU3IDpBmzNoYGH40sf7yFEeesI2/JIcTQQo
VuO+e+qioFDkmibrwtIAft8gXpA3X4mAYbrg3IyaDTSLlCMkDXbtJr4wa+m3O1NSqtCY7fCiZQnM
oBkqt+dB0z1q66oFtlzIr9ZKjhFa48s9NOBXUNXiBHrqeQwm7AJzBfg4Kl9XdmhwskohSutPipRt
LMenigBKBxbM0D1dGiNCvV/U6+D8fQvcuOJUwWqtGnblheIq3bZQSd7BCTOEWJ96XPrgoy+/nSuX
l5C+irt5GTolekkk3WMmlhvtnbWJ/+31Qq5cB+mq+ALcvLz4zRuOHq5rpOBmQaDgIP6VOJ7noXa/
GILZa9gEOGMcsiTwkqUQULd1sATq2DK1n6PuFhNRcm6ys++TyvINjHmeJM/wyaJU3Zf155lrsgcR
is7Hf2NEU5kMjVy4URun1CSKDK7Hxx6LUrAn9YkALTnLHu4KfMKIISGcEYnZ3BVnhGzAu8FTfT+9
+cRZRQrjHo1ubKnnIxDt4ooTTheyltKtdjhntc0cG97hyk9Oz7MGchz0+jJPDIfZMYFKodVSE78o
JIbAx1hlUikwjtAUxPrJMfFlb9G9n11z4QfxNxd4BroK6cBx9BhjCuefOnS1vA/LPq4Ab9I4YIF4
vl0EdwJHjuNtx+f00QySh4M2zhAmm2ZrDAedD7AwzhvI0q5ZmURLo0r4NzsXMoxI5goKR/cqZjXm
8sZID6vtjQQoRzdxosvp6adDNNfLz27C/cPEmSdCjzaDZbHCZFKln7XSt/v0qOpYnZFsnAkbRh9Y
06NnMEYFqXENZ02MQ9ccPPJ5WBuzL6sR5AIrGHF4dYc5ZCHLujeZXFkQIohVdK1uvR6l+56i01dJ
oqI4532GIAGP3Tf+MeD/pElKaA3L6yTFOXAcYfnmeMbrQTxi3iYpIx1ZuMj4C1UwLexWpg8VLp5L
rSy3qIUcnqqrNXiqbJAaLanUqI+JAkwX2VdlmPZr/GNsxbLFdU5Ax2IJGGKib5z+w6wT65tfgQFR
vQSpQq7tAC9ELvgZubeB71axZZFdAwyOXwt8qGy8Q5VV30YklcZBpR2fhAbXKYVsuTTLII/HqI2+
uMnDHknBgP3xNXqjFAjbUvtsmD5sUPU1ROXWbSJre3cz8CKFyZxzmpdUTOaN77g0L2PKHHtII3WY
yLbAK1ySa/NKbCZ9QDIpgYwRPTqlPoC3YL9VhETSmilVPB4jgzmO4Ir2nnv4/+MMBWco1CvyfNK6
iNmLU2ltelvJUMq5l8MOgCMyfUj68mG5/L9X8rmIC21Gu3AtfBWjY1/1AYkS41ln9Mr2N2reqjpL
0+SuTtVbEsVsVl+l/W8h7a9ecOnKMJX4S/BYbq9D9Y0T82Q8DJOOoN0DhOUx4gyOH/eWrM7Au8Tj
1bLEyZVPgGT4Oj08zgpSqxkZ9xJ4l5lt0mS+I4DTj+9lK7uYYjZ2xcDmVmoMONHxAQt8ESoPvqDJ
0dHt7ZNY98eD5UdBEA7rCdCHQRBi9O9drTlLaA6jrNvGFR0Mk1XOiIJ9erVXcR7tj3vUzB3ADo9t
NqWq3MOAKFqzCMMPHPTxQHSq+QMSIwn/WJArXtnrrjSGMWGflS3cFErZFK1+YMrnLay6YxIUj/5q
SDecpaPErZwCwhWfa2zJjMQycVoMhaKRILLvU6ju9/WHClrSLVX+MflX99KpcSNqGFb8spwImlgK
uvRztJYPdX8tCjJCaLGwtasIEeYaRl5h1MQ9GsOM4Zf062FYGri30if7X2A/HilbNc+Z6G/sSPys
INsKLPALLq+pGV0G73N8a1O7pwSWfb8RzR1pOGi/1MtzfuGm+fU6Fyt+Ya/PHqfPNJ2bBt574S9U
4MMcSSMurea8JahipiPKEOzI+s5d0k8YuTEi6rN5KOCKJPAXx6wmR4zfyr+a6j6eOrsTqGm5cYm6
OrYY0uM4NSv3br2WR64+EE33iKiUE4PNcXZHhFfes9NPUjXuSxqGcvtf5r1tN4MmRrBPzU+hi1Uo
SReQ3rvqfw9Z0ibU+12A7tgxIYBQPkgu5W0NL555ASnfTDWIwPDek57ZFzSh83WskLjNS97m8ynM
dnif1qyfPYhW5x7PI/zgWHGg6jVR6IUepYXGOb1p0KwdIR4i5OpWba0qHbttVaEdzDc7N5XYmWIy
ZxCOryeQexG4NiDGBPO0QnFUi6pld8+yNwyOs0tvSZuRpmZKnv53dNkYiMkdLIrD8f7HVe4AEaCX
wSX0xhG9kC23/eRTYa1vG6a4iD7roFeHuhBeiIIeWM1AQqxvjv5iuXAUHn0CyW79jg2cCM9jTtNm
vN7abL79t5GOcqwobCqSB+0C2ceQ5vG+wWh4lpimRtUBk0SA09dlQS0kLZVJOYt6XO5WNXq0pyXI
8QLbv+nwwN9Cbn+g9BbE4KsJ8+PV7qlMfpwQS3XaYnLU3zD66qkIdSxfLXKofsY8Z6rvxccCrG97
8+QZrSGVgQv6mCVenmYEZKrFqyr/Fy9fhvNfbUx9L5oqYN+etRVrDrCPYJlBpWdGV93BzH/EU9+n
1tzR03HziRg+SRTVHnco0YFqBSKHVag+6Misb2P2epSwE/v7H1ZdoYgQX/SXc4uJjyg9NSRJXw4Q
MRyQE9O6kUphCFdaioRWjS5mKq3sGVedfASpD4rjITLAQ9F/d+H4N82UuLpvT60INgssGZGoW9Pd
Lqh4RD3thzWdY0Y10VI8Ifi2txTkrPt3xPPbzIoQb+4AOvQbuc7DXnzSFz3ZdG3OtrQDwn+TdxjR
33kHQI++uhLwkrYSw+1suhm7cD1OFhxAyIedSuQflI75RVXuJT20M5dQdHa4ISUXJt/Y7pV6YtPx
3Q0/OySg49KpHwWU3Yed+LeavCI7PPEopGHxRSaQW63D0T6H8aA8GzF4B1ORQpOhJ1xkxl9jOf20
VJTSfa9069nheqHXp4Bc1K0RfAcYC4GwZw/FFugv7M9737iEey9a3W9td+cRHE1+RhQqh50iv/z4
5ILl/uNBY3dDBc3Ak8T2ODD9BX32i490tzNcVw8okbEEZttLO9MHe1onDc4zIIx1x0UpckHTH3O3
HBBX8R58grBGLEyktij1nRKCNLtg2nw45Z/B2/TBMZuvI00uquqAw0GQeOMaI+zs49VoaRBrh+hu
07rk5Qb8GgngccHq6Gsqoz6UyPNeUq6C/L7q+Jta8VSmfAdtC0WvUUrQxv6PSMIvhLoMJZDm2Gbc
A9gI9YIvIhuvjfvqmK1XwF1TaWSba30SIJ6PoKCGqLRzmHVne3tGzqO4DrDYUcuRyUV1jyDwWUsr
engudo8oi43Y84+mLzwCvMWmxd5JO6FXd4MNeQ3cRYTf33hY5vYv/po0bYug/xsADKvUM74PfSY7
3/YHB0R+1TD0rnzmjQAQv/4m2CIGZHbORUsmL4mPcnadjUokIS2ToYolrDvDxVIkqLUWK61jdK5B
MuURiy2AbiHIw3P+ixT0QxaLn+q+Km24bk/Z/StcYFRLoAXsY5cBFxo5OnaYQ0pTVZ4kgJ5g1oBu
movRXDqU5f3yhvQfHvHaq6rnzR0wU2uogJhvT6Pha+nleFpCQ7MgsQICYhhZmlc8aEaTMr48DEvi
mmfIJLu56zWIbmhAVa2S3LhCutp06sOUpGWJ5vF237tWcdhyIO/FISWhnR3PeOThqdxplFI26x6F
KW/Errp225uLQEE8cfw8A1/ucFg67O11M1syV3bMfiM64Pc40o0osy8LNL2e7GRXDFMRR7CwrXjN
ySw/mvKT+yfUghKI+5ALRjus13CQIc7ucafcbHilVhPWTzfKETq1C9yyADFvHtXWYZXY6ZUcFUeO
4PwVcvnFWjkSupUbmYZ2jhTkTW/nTQG/qg8+hyUDEUXkSVfHXq4S1bb+Iigy99vhlDhHDk/cTAYu
i9udBxa9tF7x0P/uCumjFwh0Tt/tTPKpoY/s40i16NEM8RD39QBzhXhujq0AUaiR+dKf4QB9zxZf
u4ZOn/kO+E/lTs2x9I1x3tz1E3RTWo3CzXSkkXEwEDomzvvS5IKDzzvV0w3EX0NPZDK+ncrdyOE4
AYvnAItoMhvOk4vokboRNVRiYg17V0nWi0sGrrJFjGEUzhEhqd3m4zv6dvpnUS+tnqMAnYbzBgI1
SivSQJI8tAPxewgf1JnCL7N16VS2XsgnXw6vxjSoSVnWh5XCj0H7hsoFBEJwGWOhTeWWGg5NV7tp
nTcq0Huc9i5zhgFhkYHUv8edA0c7AEZIQAVaSgkUHIluTxnqQLJHlKbUJRTVF7VcfdliaKOWhWsW
JJ7wOGGJSiX/kRkNA6SH6CjgAQ5FkaMzTlxk3L2cqYb0uZzUdXVa/X/E2zaoePRyZ5+M9htQF/cv
tnDJ2U/B+7hplYP3LNQXpE4c+ggOVf1VrGnT4TWXDNYMBrGg7xW2tmhlwnuPdCBnaP3uqA4Cjfaj
fPmgd5Rq9/LUAnNKNWx42ZVAO3gidrCwIAUFPUnhSelfmYzC5DO+9qxsHgvngvlxGSWgVtc2qHOb
hG3qWgEytbEIYHw3QTA/S2IWQTm3lI8m8GVQw9ae+r35nejhIMMgeqgSpLa/VGuQT549IWVHKG8U
rXqRWfI7IOWQNzkW0xsVRkABj+HDFiCO/EHgBbOwxVoQYRO/AaHBWWHmGnW5EPErT7fyeAD5FBiq
q99J5ytrHM9ahRLPuv9ai8pNxBvljFGF89YVGh+PnMxVNxn+p9cRUVjnv9oqiaq/imUrDu5fb0aF
sNuJDKttNpVhwkd3bg6JRaaR9EUVas9KBdzJKnlomOynRN7x473GcXc3OczfeA4VZLQuAy+jBDEe
l3YU2+fPGRQ6wl5tZ0vipx8ocb+kifA21ShXc8GKjhc0usUIMhOuh86sxk67ZzmDT2yf6C9shnff
YUPls2BItN+nKgyavQGo4OtQjksdawdKX3FpSP7tiZ3Qvqec2yatCqakinKoqnBsegv8nLQUG8bP
nLtZT2EiCkLlNkOlrWV7yQgW8vDEKeXjc04g8CRQlLIAaottbfoXXXMQ+2VM8FpdM2JxjmJEy+16
ZRy37Z5oQEL2PF1i+Y+dq8lMn8z0cm1NsgNZQJvaRvIflvnI5R1RkcbJ6XAIYZD2rsRazf+Jq5CP
ER8AN9Z+5dx3zQcNDfNFPYNRYANSrlSjPqLHVXJ9KWG/jcy6r/Bg86S0BdmovBM94l4N/W+w9jLK
v+WWpeX/QCA30C0UTK5IGO/QV/oKySHt8IoxJAY0Sa44dCZrB4jQuU4xO0sLFcaIz+9hKHeIWT3N
TNXqojZalLjeps6fsGmH+MdFXiFQIduwbxrkgkm2q4abzQg5wvX+BTdn8Wr3ZYdrMqjfSzbWOcmO
zVCjK2UQc+S+S3rkYbx+kXZRGlZMC1vyYTJOMheFdEkHWTA5WJgQk6Q9jOaUcbh/4nOyYI1WVXdV
FxloWX2MKF4WIcr1C/w4/Ev55/gpKzyD0cJA3j50N0Ys5gteHA3k4cywtbmCunODuyWJWak9VqxK
pm2DMAcRgFghzE8wTT8WbH0syKuPl3pnnBRfTKCLUAdEHeg1lvccMeiN0c/pe19xhOIJSvTa/3Gf
uR0g5M6njZD9d0pN4e/qXKVgNFYnDTfJiTUBaEIUrd/90lBjkEmAOIrVK/DCazNIjqE1B9z+FI0E
6jDQ/vkNc2Pt1lYeAd+UbUmyTD80AtJmHtG0Ta8jET+fUbjQVXi8Xr1BUw6k6UoyHbuZ9lGxf1aE
JjwiWcVKi6z/BW3jnD6FmRSjl6c26rsgoWkUuWKDt+nXKBhHQ67/Qp2oozPYYKcn2ayBQoZMpdv6
l++yEIZqcYtVEu3WiHiH7kL8uVw0CUs71shgZ3rtkAF8gLODI1mzEsVSW3O9e1CB1Z20aqm1rTye
NUZ5v3Z851VY+g7X0E8HpD/uyLG/RVEjp8gZyrnMVDtxNRRs7BrSz7ZDW7rPoZBQue3oHfb0GXuE
lD5SEbuTaTX89VRd9guqhynoYvOwICMnQhy4ReDEvfUzvIc/OVgl3yv/fkMC4U0i50DXZ2zheQ3S
rigm5vqCFOCEG0Qv85AEwNlM94HhjbCvJ9S22LCtZIJu+Fhr4QB+TLJnA0QDYuiLm1GWlimGnQCn
ZU+gzFx4RsXODspK3HOy2XsBxPhs100yPvQzbmmqnjOuBoR2xFn3GfLuuc3dwv+X/S5Z4fvMPqOD
UWlwC5VA4WHzi4v2AFqoNKM0ozWz7lIaMfzhVefynwffIbBR1zlVNbfKWYmQK8vnHkTRv/fTwB5C
LVdBRQOqFMJPkPRuFmR2cCZcirg3c3Vt3PaXMDe6Lgz0ycs1OoSrB+oWWatyC84/veL542ZyaDyN
AeZNhiKGaG35PHTTYNMUfqbqM+VK+8ONym0kjnyLnrpsJNXe+C6/JSfjWrv43l18ts4ydNc635H7
Ips/E17zmXtQg9F/c10VUtcQgUmczFEcXcCYo5nLaScooSrsrD3aQpVu57pB5lKJdbKN9fsEX3ca
qrtfOSJ965eNc4dpW1086NCcYCSxEH4Vu560Iklhnwp5KDKIx3WGkWJEr/4rTZyN+LDu5dVkvt2m
qy0T8rAHDAX3D3HGZNjbMa1WaKsjAcUG7iSeK7gBy0IeXRMAbXMpJsM54bMEBChlJVwm9jR6+ikx
0zUzIutn+D/Ko+E0rOUh7AiuXzWUGEVJHfp9O/TG2W3DuIn1IIbYukW1hMu9P7TkRWuxBHUGeeZp
hliSyPxC8aZO2mIBmkhyVomvxfxUIg2yelswiOQAN3EHKcWsZQXLsfwPXGuvK3p1rSxpMj9gS0dS
utLQUUREy6J1qJpiiWKLdhq1Vn6zaas0XPVDaYbSQMvDdPeNEc53D3xgJ3X2S+sFrzvC4YGbGN7o
9SKHlPSkCp+S9hAyOSv0+7x7c7w8qWFuZumBNNMUsqpPVUnUFcRwDgOV0R2DqrzQfHN1DxH3NsYr
Chyejrc2xWP80KhxVy9WR1liQjb6Ir55UFjt3Bqatww8F/7Y/RpaaDaIaRTqMELmt/+QSaGYI1Rk
6YlSCbAwGOaRoGMcXvHF1kMHcoEcOjkvZzd5r1YkluChlPRTqK2xsgNagIJnAVGX0aS1/4kvQmUa
U1x76dcbtScm5UiVPskkExDgu2FDTg5Lp813oKbr6+uAqMs+dRr8vZvYxS77gdhD3ucfptMHvkwx
iAywoLqLGIBiMJ0cJR+rlykHNYWFs+RBhNSf9lhqzfiGTmakuNG1k4pKt4kDuZWL9QDIBKJk/zFT
3X6KRgpBhnamwSKt5RZwvDUilfjMy5aSejwB5TP7B0gQSLQqAftj38bRlSzdCcqVrq30MjCzAvYK
7XJy9OdKDSobhJGtyOsbb/u6h5MQx0sEx+GgrEFG9MuLA16E/zPdPGLZ5adA1bhYftrexk1ocYoo
5h0A/Y3Rjh9S4aHgbMpsoRMKGSVCdj/wgpLJE2BFiqELk/zl0fyXtjgiD88+LFCk5Hv5PqlAudyq
kxFmyRlOBw2qpuOxSYO9Zjhxv51iMEmubV0N3+qAvjE6Rz77qdGiwctEf1dIP9Wa9kV75b2oSzPZ
FhCvUS+RsKohulCoByOb3Lb54Pq1zpDQeaI+EAxvYtM3SapPo+5z8eHT8m2cy7jXx0C50DjzorfC
IwXUo2d6YD8Ft66vlERosRYCh7VxwW/FU9gWeDE9ZH/atuseM0NhgIpKPC89W1ja7B19DtI7k1AS
rFznMkDgvK/BQSOClhm/UDUGsZtDGaQgZDmgIA4iJ9QJ9HWxJEpXd7bdZyYFR6fhp3g/Oc0uV3Jd
Wz8BQYUaNBvRF9ULs0TxBPmZy0+1IB3CNskf8M/gzU/XFaBAvQOBe71+zDwe5r8VU/OljqPSlT7D
55qoh+yo+13yKX38zGR9lpv3MN6W0gms22V6jHL2P3SvbWzVXCOTqamRiNm1QE1STxIwA16Kx0qL
HSIMDZl5W2bVpklNoKereZ0toN4NAk6x4XQfsJLDvuzDsSk1SDOcXz8p4VTgNzMlg0lL0s8f5HYe
y+3c5CgdhiNeyqvqklt6kUTnf8w24OHHnWFy2JbgUHrvJzJCy+sgDCdkKofcf4UhnwzeH9aX4Qpw
elB+CQX7X94CBGFB3omQKSyLNWhqc5iov8W9tfy2qQzqfYdObbYAZrRszoTuUAFlY50pY/XUJ5II
aF3UZUYXUW7PEJTlolL8DH96lQpJ71g29mauW7HQ7uqKhlID3jlvvfF11DlsMH20DO+tAa/Hlveh
1omxIGYGpyCAcmQ9X5FUN7Bco2VRIHK5x4jLrFxkMIilbhemJ/FvAS7t9tuhU2Z+hwqW/UPpj/LH
fmZb4nJhimX2JUohsxec0eCgdZcnLm/fYxFzAZhusdt/HcG94wXCAbQlKMUqKt2ZSAVEe7FJCfSf
oViEkC4ZqWSA9Bvy/yA8OvKFYlUvR5yKTKK6Hf3Ut8iVxS8KcqjmeaoVYYjx01A3nhcktpZ9EOZV
qykdTBGEgbw2ArHPGsw/fB9hiA6cwJDNTYFVyT6UWKWcj0ostZt9jHXSwkXJ2VSFLpKJ6Gu1+eqo
579+E80wwZ50LEzNQQSmOCz/pltUQhRkiRXTh71axdCeojrU07wi0bVMPjk6cu+3IMgWyw+/7wy8
I2yzBDNO5YYygckA8jKEWsoHcbV1wZ7cnEWJXPqD6Hju4ropsvsuVjwR6tVeC52dYbLVA3FcVYCf
y4cfteqkPCHyiyXM6OkMuAiSGyBi0Udg0jK2yFNLSGgs+vzQMJaRTXo3dLXClsVUcRteBD00vEcj
vrZ4xOvmO2GeMqHwO469Qocuzed/zrZlAf2lnYZFg/mOiPku5jRhuj4Ir1KXefhSXV/oCdtCVuBU
kUTSPfIVfnmwzkM5PSamGG3nOrEXyT5HS74QDsXmF0ZTDt4OTTb/SnY8Bb1YVEJDjH+nXAH+okaK
n9+aVsVwSMGr6HXcUZnRqbUERgEQtexiPIEc0UYFAQcOl7VOWL7SkSe8FF0BTyaJtXjnmewI9ty3
l3dkwXoRBIgJpWuFM2YtDhxgsILR6X+wYWaNlyq8SoLa0i6FuZtKyjKSoshpwVXSPdGZbe4Mf+OK
k0+DTzntYTuSaDoi9PSdlbQ7IXeexQqM9U6mm4Ipr3r/yZZi3Ky77VgFFvkOCu3aKr4sa3lSt+Xh
+lrzmALBxm25H0TUFVV/B+epAabLlbufkp5uu5DrDM5TieaUUk5zZfFGCnwvyYp6WSJtqTWijM2o
bO2+n6eTpyKgmml5RIpq+9RqXUo9gg8cF9Ckz4hU0RLYg0BHHIikhc+kfDHlVNbWq/bLxsYtLRzx
/AvmoQwAqSX3SgLekdUujnVl64AoCWn+UcB4YoG0RHHZ3jEgsyLP0VwTov4I5bSquU+jascAxcUL
4W/Hk/OKE2J5883nJE5CzJIbass+24M5JGFvl2la+a54RjBGN68A6CWeGPZ3T/GuJK2KDQzr2jrB
GwlSQszwZi6D/J9dsFxHSgl/Zy4m0vdbHCpyozvk7HFZmXjdmxmMclmibdbkYS8wLEJXA9breHDy
Vdd8WHv6xAWYDBGYproTKoPQqCs314nhognO8/VwWjZDB5JVGv0veCphARYh0eSIMPnLcnPg2yjJ
ANagTt6mAjKdJ93ZMYcjxQbUdpmvF0KfqaQaWbKBEECYHT67hteb5B1CUo7b7ZPL1Bpj1f/bHM0e
TXl+KFiURnpL6PtA4b0z/UiLy+gij8sTaP8g1RSIKPzFqmSB5EzS+a9/VREDpIzNwpZ3w1d7jaRX
7j2VnS/mKvT8fD9cNHEEImRoYrtCgpcCBKpzsqMAB7FWyRZbyhuD6kT3xeaLfbvcmVVmiFgbefXX
Y4Am/HSoOqQ3B8i6YXa24uaVCqi6e6fRAqpUFnKSvPQLN12yXEDKPezedJ5mXVkoirOixWq9Cc/P
QCaNteM/AiBm+ay+W5O19jw1OWw+aYYPxwLjc/HhMGl7YveKC5nrmA2xWG68bmmVGb5UQzCQvqx2
bM5jm+tp3LNmMunrxK4+cgpTuHYdVh0WcUw+zaa6JazW4Z7zLq9UjsBagIt5QZvqAmc3rzQ23oqS
mBaSHWAQ8sBpXWBMAkO4HssznWtbNbozAy5lE9SsjH3ReHwLapblpqV+ddvMZW8DZDCISZOgtQLO
3VZSM+VMZjcCBWA5Zgc819Q26YwDD55p2Dm2HRPTzRrFcfwjUgNcIFDkYeCBEk/4AORKsRtZDiou
OIrDl+aF4ZT8+0D9eTohFSBuwKRJyj4jasjdNxxy0R/Xughg4NuNhwvIgUcHU3Dnj9sS1B+t+4/Q
kLYANnyyF4ZEFEuUT5fdF5W6qL1lIGbnn0QmqH9OCZPfCdBLihU//WZb8DApmQx1+3G+GZoMect6
yR3l1sVIJqE1B+Kn5kstpQ0GkOCZptRw6y/OAp0nVdcpJ15QYCrJW+WFCTOpak+zl3SHCe3uioUz
ZfmbvzQqp8XEYKPNDcNOyUWRKhIvCCWqBmLoVn3uliJYFKpgpc7O9AYfgAIwC0bDG0+O4H/7AWvM
VuPQdlZP3d+ug9PB2ug1goRZNPTxyuvx+P+EmEd3oV+pqfTc4Ir+Owy852tzuaiPSxW/k15VRnvw
hqL0cCYd3qw3udCwepcskeKPKjsLX0s8zBW9PyqcYi8p/o4RnEMSQvjtJ2Hz9DypEOoLpo2/Gxuz
rICEi9yCONbRI+AZF77VY5FwUHPwPF5xp8cw/votnH2YJQQqqOG+MrOUA7enbngL2USLDzmqeMXE
Y5EH5vqNOeGnNQoSTtXY5wUB/LmfTgL60hmx5f321ZgJhAH+3EuuGXVCNqWucF0uB+3iaDmyo2Aj
WRWl2sGUy+UlROxt8vpjDHkErfGVjuqFJPV9YNMCvIIP+ZN4zMomR3j9Qw3dFYVxFpnsTVUDa5Mg
OLXR4vn3NNn45y5x2lPBZYI679ZREbIGCrUv8MSf7TpUFnd4vh0JonFnAnwNoPCtm2Pv/ilLR5ev
GrpILuPn95iy7eX1BWctT0oLiE40bGrWD5nOYRoyyLv66fjLKS0Z7OwkPA290TIcHw2bpjy7RmJT
7uUAeHYGmHK66HZzsASapYV3NAtQanlEDcN/5EyS97BxOe8905926ibqJ27bWzcdnKsmFMBQK40t
IJ0FFn09YYhCa/WLhnv+vta4MJo+nrxS3af4upT49V7DrYe92IVYPCEvlXCaGWbU+MllCEdrD5Xy
8OqYA9o9WOwHJVr5IIFMiqW7gA7vlzV9/wnz5vcBlKu5Zx379efge46MWVrYUlTjb8ugDrMqSgma
yKbBofCMRueMaOrugqntBTQl8silMRNnE54jUWGRc/dzWIy/fzp3SZggNxKxYHSHHWtOY9RayUXJ
K8p8J0OCkFOKTq4fx33zyPpSwYcJjd2utRetKQO63eU8D5nh+uhd1lD9q/+Y6uCuZePWC8L6CBX6
hJA54GH2TeUyD1hiJPOyMy7q7oNTqRUA/QoVXMw21cJ0xvc85J7WlPjq15wNBOXgPJRfFSms2JtH
eRBLycsysA90z3VpFZi4Ta9TnMU8K3vl9+zKvXb1rgqZU6wDSczppS/ij7f1A+uyyT3cVayugNkq
ZEYeIxBIwrWs4vPhe2RND4tSMLIzQyPYy+DEa5M3taHr/cA2he/Z/5affZk4qkKCFnxqSGnHVtXe
jWPNP24+Wt0d/771aNCLIfrEPyoMn6Le/q2ghm9nO3EEr+K4YZKSGb8vntNjaK4fXyq9256/MfcG
pSK2DFyHL0UIZg+J7KWC3y71xQqtFmlEyZrFL0Ua5llDdTwNgwi7VCiIYf93EYAxWulLwIcrEdqd
nUjZMsfe3hG+hq6z2mW1hJPsRsXr7ZcyzWDf7CZvCZSLvpEm6Ogz+QjVy8UOdGb+pK1mw/ICM9ud
BPjX0+ojEWCREX5lAQZ1YZa6HZbL3aV3qzMQ2DS7CDVMdK/4zy2M21LuRJhXZlsWLkN3rbvFRgEq
XDarGlCQV2Wm1VVv9Za3xdZAoXgHwvwONiEE5uA7ZB4dsiozXeCV7FzkMSDI1r7f0HHDrgg5Lvx2
z9RGmi26YxsqkzugkFWocorYD103oDUJMgLDvFWCMNUhqa56/yEKV88u2At48JmT/3LVPUg7s/Cu
MvGjqDk4jOr7FNkNfIh8fAjEq8blfWlKobd1+xtz6clgF2LOxV6weZCWLv4XQYovb9J3uFuRKHNU
tXAKdWI5K77X/IlPQRQa7SbiZ01ZuZy/Dw/2UqE0A0rxm/eAd5W74JhzV4EYQas2pYLm8a2k/K4E
NDWBLxZIfpJ5hxhKmjKJBRUOF2VquQks5eINkF+/YKgOuV1voA+htb5mENmQY6ErIqUPHkkXFcYz
itN7DzwPPSPPrwMqzOf+sncSeZFORDOeFc4GbNo6/bhoLruBkUWOKGVrD41Zvf86gp0b+zdEhDZ+
jGLS7pM4I7EQmU9czoWqbpLYf/aUkXOveLitT63APNug6/VomWumFKrcCPvyHEtrxhL2HNaAB1fe
ukCb70Vm0aL+HfVctneALAEFj/SlmF5ZpYt/fb063OmZipVlF3B+BoJL6t9KM9fip0DRqSFcmC2W
/jTN/OevD4yqviH1o8wFd+QbawNm/Dg1WQ16Ugl/wvrqaT+9sukm9mGqSJB1IwUWzwC4lNV28hzZ
WSKJxnagVdgQty5k1nLQh60CS7yknTs7Yt6I6xyauPMo05CxkmgY7kcUZzyLWK8etYsW6niHxApV
ZYWMuQmfQJxXYKzxqIe6ICgZMgy4GWJZxbCep5pVdO4jyfAKFNbcH/bJAUePgyMxW6XRFHc8vgPW
rIa8R+Jdtr+eJDn/uqwDRtx5pWsnZg1j0CrIIbgnp8Ovp9VeIm2TC4mHlNazbnWGX6pa+lKVhlCS
IVYizG04565sz8Jl3boOc7rV/QeQOA7dmlmDQMX8W4u4QRX8/NdqUdjmidgQ4xoF8EEl3apaMmto
gQGdeWV0vkwTTbBjPnESpP5dt5d7FyCr8FqrxtvuXC0FHFzOgEDHYRwlfg514Umzlul0RKZElUnT
Uw4OMgeun2ZDNs1y0WJxjO1UmlRmEFE/Ic3P3oMVx9jihXoQokNKJnGSSBDUWMDyBLVVIrYjfKEq
Iq5OheOD5ZRuFyrUcD9nN/m0D6lyZUXVPwlrfVaX+wPDB8M7/zx9hJ3ZJUtwIt6oRNlqtHn4V7CB
F1Wo+L6eeEbS6HllU6CXHb2jKQlKfs1RwSrle9XYSZ47Jqy8dpjJc9TtmfugkpwZmp1DCcg2RIsg
e3GXZFSlZD3B6iWs7IDtiyjYHhtKFTx19JnGnAdP/yAwGvBqQ83iUJYFzi39fTumqW1dOD72mpIt
Wjo1oSGwZyc+YLG57BmW3TYJj04HoAwRnBJgnU9CjHK/DUFC88sfHT0b7JvRk2klHn0XS88I6asi
Tjk7t2PXwLK26A5iQb1I0Vsus62vx2uzJn2vjrIcdeMT9qnlBUnYqebw2Kf/njVmZ3cHoOYhsUFW
yeYvIkRuljelVDTunSqJ4MGAwng1q52AjtG7egqKIe2LeqRX/BOZgnHooAqVtv+nkWzfdv+obqW1
r+WKzMw1eqEn7BXz9p5u9ZOVFiEjSmIW3F9AtoWZJD8vJZUUYB5HVJxv4z7sTEw56bnAX/a/67JS
T3OqGYRIhEzbe9OF/mULCpyq8ZjtJZ9AXoT24xBe7bKMwiK8ISNo7VTrOUv5souZfCoZ7e7nwH0A
7x2uPmriX0w+Zozjc1rzPOM70LRZKdUzp68PpNEN8PUlgBpQbYbK+SP9c1galJ44ZBEDbdjsRyqK
6SUnWdHl7tdFdYcc9bP5tj61U17nRwC5YpFcgS72B2dtB32n9dNaOCRpxuYif6PPoZW6yomFw0DB
NyEKF2MQ0ow+YGclREXaN8psplb7L7WAzItpT2p1hZ6ha2yVR/lV5z/okJOHIGX/L+WxtRnoyitn
Mzu1RyphFy39Oz5Y8XgeZzg8b61APtsArGZooI6ih58AWiYJ8AeihBRdkHq3igPTsgiNddir52zj
aHPH3FoXNzcNVl1GAHT/L776c0RJxeiVA/oDjnPe21B5Uw6cYOBkJV8HqyzPts7Sdj/9fSxIa5Mv
164YA/UKczMIQKJAGB0hZ8q8EitXGMiEuwbj6yuaYeVf76tO3I4u9la7YHyv0epFRz4eLjGQoyz1
PQOi63b854QelUoG2giU5qwTgpQy+xr421BMwWGIipNDd2FO/8vpmmpiVcN+PygB/+jZDMCE87dE
KnKKvV+vqf3YRo3OYkci8JNfyaMT7Rw+cuauUGWpAhLEY1dnNcghkl9Vkd7gNf+9LA/bvQuRcxgz
Ictc5jsvYALfU4WenrzwLnvI+FT8p2HyssQr3hld4xhtY/OOxbedaZTa6StcdAmpVAM2oxPDu8OX
Ta0ZnAa1mY+KwopTvSn1wlvYywUX/ZB9HZrAhAQ+bimum6NkR8PidYTGnPhsK/n0S/ez1WbHpRcB
gbmN4NKYnM3T8O5nHVBpC1ZNdalBeqvFDoUzEin0hL22tCftEL7bvzQhbGWVKzor/lp9RanwBiRd
oBXtxCxbd4dz9sCAoJ3EnF/fVvjFqvuvLmPPczfWmWXAJrzTjOG73h5Un0KvItzMzBnr5CCsr10i
CmBskMGTVpm+wR4Fkj5cdTpdgYkEKXscYvJxzg1vfFrj2qeN5Y0Kx+uEmqqybWoxdu4RNIbc8h41
ARzrGXl7brHKH9I8Y20vey/6iab3BOqV4ULPFWPrEsucTy3SnveA4PmpTq7vyUQz5pJo+RPMoRpw
cN4m+AwKrPypnSNdtk/3+3IWAAx6EOHWaxUTBOpVekhXVoJzOQWTWgGPK2wd/PSlOAr7OpSiIKyV
mV6RhVRwBLum9XPzbJvqeOYDDJ0+srDOM7tiUqgvnirCmocuIGUCny74FFWs9Le0/bTf1NqNcSc9
WYMpp3XcZjrp7WNeMhsazh0BTvXU7HxSzjnr+uK87TpRfBxNfBSGcyQCX/scjlsk5Tz19Y8geW2d
iXfeSyDKwVlTMS0xiYuFzXC0XCYiW8ozPVDL9E0bRwLu3Y26R2yp1uByLHDoej1IenqQgaXBg9BT
iPnEkIVT8Y1jgnfr3Mw0vYVygkpMa6Hm40h5kxs5SyUbUCopPfzmNvo9GDKwV0KYP//Ior5jG0+t
S/Gas1yaVD6MHjxiZflvyehDV793J8Wg5U1ZwFtgvlIcwCswktvmosSaUiC71Kq52KWC8PtNFI+r
U7LHqBOTlEukN6aPZ8p12aEQNvV4oxBVowzpOmb/bBaQme1XPgDtk13yPkIkSBtb5n3Nf+DEqf1e
CxzUvp8TND1PETYIXl5jaRKmi/KNzX8VCeifiMsU3IUtbvfhf4f5et9VW48hCb/AzhNdupofOStR
Qo75omFQm08Qdi0X5IjAbG+uaE5VUPi7dYkmwa6vwwn/w2e3grfIg9sjSlDG5DOaT3I6QvJeyHJL
Z59VIzMoB38ZyNEiOGFlYiCFEiIoQrkGnN3cX1DGXmHJOWXYaMLxepIggMBP6ofeoOMbnazZfaJk
nC//ow56Bq2+guuNTQLvvvRzjT5RkZ7mhXnPVjpqEK/cyXQpccJ+dnAbWQZMmfzKQoxE9ubKyKIa
AlvZf9Veu0SnX2UZRxvvF/XnuO8znl18DWBKl7FqcghpAchs1HMFpITjPj/AGiW3In+iPWl0b5ve
5cUF2ySquPt4B0vm6QdaKJJWkZj9dDzf+eISgVR4c0DcT1gbTfUChwiO7kON1UdfSUKy4sZi+LCF
M4ix3b+15sx4XBc4haemgcVCeIZlF1reZiX50SyyjwjINhFEGISveSvgZBQQelNBpGZokg+2sW6p
icE+XFYkCSoAC+rMWpMFSjmQ6HQxp+nDFrrdgme39lszdUBLBLEcZ56uuf1Aqzj93lGuJONXWP2p
owswv+jQwSz0h6kbgSLKWejIcPsrSWQZ1o+JLwLOGf7XFXnithPvswy1DNm0FixYpy9rn7rRRsOc
Y4peE/a1MABZ/q36NDzhkBu6s1JQZBlrrbJ73Wl2mmVTj3UO6s5Ruothw9ZiFNgOd4itEO1d+BwJ
THQCmQKLqEAygo7FV+RRsEZ3JV8T+asXO2XQwEUmZ8s1gs7XojZbZsK1orJfPf7ipVOEzJLy0c4v
Sixz0KBHFOe5N4Fs9C9xPHF64eaUQ1oEF+fd79Efh6SBpZ4QzQe0EyPhKb6HYf6UxhkfwLva2fF+
0Fht8Ln/I2NY9YiGOSaUnD3QP8UpOhSepoJh576b7eqMUo+bPbXMyvcypcDSlk9yb2+4U/fKiFKg
JgOV4e43PFJ//p99eykI38wiZi++/ndCTeqWt7XZhcIJ7AvEppXbHEeRf7tafnOURH7LTRd+gdL/
VNxKQ+vJzQ0neb2/pNxwx/WousoROxQQlXrKwfBCyr8owWThZU/ibGSz1+VWgMpD3caVDdBT7AgN
mTvO2v+P487f8GmW68LfdBiOYXpqXEk0/CoPK1Z7yOlbcIvwfp82/XqXIHiAUm67QlDL5WP07gA6
DSc4Cip5D2ltnYWDz7AGF4lzyRxd5GAf1EyiLysZ7r/k/aVai1TvxbaRmOH7xmuONH1LvWp0yVrP
5ivDXgU2UclpCUuPaP1UvjbDocDq6Oc9bq//r3SIXk53t7qQf1ady/9Zu+HMc/jCFU0KDFe3LmN8
vO0Fre/9unB+EXDUNXc+4xEAjYSDzzMDe3O+cjurQ8VjTUVhTxFEurUvl3XApRe/DSkHntI8BGE4
4QHwQdq3CExu/+BoZbs3tzyykYYsJl7n+Rfu3UYSCQ3+avhyOLuKG/LwIaJMSdTQ+ZvxIY+J8Jn4
vFb/yhiUW5wIOdGp0pg9aNf2Ehfpbk62b3kMsLxJ/qp3OzqpAUFQ3eXuJpQlxg5/7x9xC65Snbxm
9rWLwbE3jZ0CWX1/lmWXZAIEFObQv51zF0MEMTtAdetImWvzmhB3HQ2898wMFRfQIiCBCta6R0AP
GnKS+en2QKT49XC7ZTyiYwACNZ/jWD0kFP54oTgCf1J+TY08y8xvMfdHmTrC8OJUuhv/CQBQKCQ4
SswNjX0CqU1xk1Y2/CRP4E2ktgAV+AYEcn9Ryy4sgNZLFIYFVqz6IhS02eWVjv95xyGRV773QKlw
+fZVmA9srUXUCHq+fbyAvfA+MmqYKjQOzaxqv420nAeZrKEmciw4QwBFGaLwAG4GJVQbT/pv3QIR
rDta6MqVJIGQb9UR+unPbuconPVie22aWHDrCm1J6+cM3H0lo870dlHE4ZoAp9lTTvEPRyOSZTFa
ibgR0qVRIBBKNuS0B4o8Z+qdmuguIQAhA/BrPzxfq1fS7YytmoT79tMsmC34OVUiq950ONeqhdPN
YrSdg3kEb0E1TBajZnvae+/1a2NYXInK8ESQOk383ciHvIwBja+Tm0Bl/Ve9rg4SFuy0cVIOVqjL
/HVxdnNOPJg0ZSTAF30Sh7qoeYYXOrr782i6Bssi14gHs8p2pxP0C6yLlb7jwIzAshVVinMp6Yk9
T3sMzb5LR46Al723j3/iTnJBl/rBA/nN8ftkuCxnlQFL5dfQulrzzDMs1UcIG/6M2YSNXzAnRjb2
bWKJL2CDAGcRjxtGfiTOceRAxgQBskMiRjDXM9nW5ZCZrVkpIAgZ3uPHfG7cB54csV48rkm6v4LE
fW4jbV1z1z8qotbvl/cPRm3eamzSnRYvTXFrudBD3rSGHf2Tir9XCWZCtlQgIYQUoH71zc098hxS
3LnAOaxpEELkyniGODdUouzM/hbr97MCEKpGokYMbbVPBC0ur99yW7Xn4wRf4V/ZPYf+KlCuueNx
QofRlhx/sVE7HOIZ0DBY8CFyt2GpBXQGhX6QEVkvDfouPBHHYc0O2QF6lEtA1S85VH3z6VckHBBd
4RuN+pGG4RngadpL32MQGb5Fd/BV/FM8aEQCqzNCKHRZQmatsoRdrcfut6RBMMYONzvFgTavlbc+
HH68UvDAyqIv2XNpWcBFsF8vIyM9vQNvdWKzWtH70SZMmmF6VWSnVwUtdVySu1XH76FeX2A/IJen
Es6y48Pm8+ES7Un2rjtyGiWHvlDibRGg2OrSa16WQcDZvvMbtS2qF1dBonQWnj9ILVjgZowfozBm
iH8YnvR4XoJkf9m1jV+wuaP7+F4uGWbMSWyj4t/Ay78SZRmTIuxaJ+UI7uNCOb5Yk3XwyNP2OAdj
fOGkznlz9UPpxWL4WrHrJI2G482HBRdV6uUbSKsPGsAYx5NlpFDVC6wTe0Pw/J2i4WHMEkK9kTcx
c7jkFCU1J1aTuplEnGbSmuuamFVRggVhm2qCoppOHWf0HmoIk42igtt78+Yo4Te5bM83jGEBq0rd
2ZtkJOBrU+TobrKrZVHevuUmv8ZvcYUQYgc2WK9SZG0pea68H2Qv2boTM5DQEdWa/wZ7ExmkbIPa
7paMwiaJIDE+0mhQQq9zmJu5RdfkYr8EUSd1KHHUqJbAxJo2wQk1oQ6SygDzsU7MCm/WuLAfPrW5
8GYtLARYCk6pc5ggos5vE+63YSJbn6qKhIXimvcUpqtdLNX6G5HDjOJyRyZBXknp4JSTRNkBM2Lm
2yXTYUgtNKsKxFbxMFtK604ZkUKsuVAKtv2CVJQSsrPK6OaMHOTEppEmHNfftMrefJLD0DxGO6t1
wu6TNIroYZmIsYiIBF0+DBZypUfLpIRuLwkhc+zOT2bvIzehCi73Cn+wT4fQa7/6aGeHG2jp8v1x
QuStM/7NdAS4B8PHjI+y0j51IhVEr0uoZAthFCZqTR+8QTniRBqlVpmJDiD+cbebBzSF2A5VIkVi
2c5wu3GevVa2Uj2B7fdkiEQcGnVUuaNCxXafh2Hy0g/dinUYJhilQRE4kDVvTmzSBzeHnLWbNLRR
neAEsyUe3FHgFjHIrxbOdx6nYo2ZXeYkw2rPLKy630HxX2NNzVjO0/CU2O+jXuiKHNmlTgE7r2Ph
blx2s+UV5fjB92ladrxZoPM3Xs++OPuRwBdyBYvkSuZPFt/ZI3Atxvaybm3QZ/eu5NJH1LoOE3XM
LTW9MKISwhbb7jzfD2fFGLeDr0qPRDzm477/OBfpLUC7H48CoQjGXVHUDGqEMF4/tOg7tgHv9MFG
K5HFKOsveT4BHcVYLhUxBI/7IEiGsmE0x9wXXjNRvShHxuDVb7q1gltt/PO7Xa1mgLh0DJSs1bVi
mNvO3QJoc/n3Wu/qXVOZmvYVG93Xpv4PdUsv26dbtyAswhgk/9CdVH245j3rbGjOYav/154uKN7Y
baWZaDHfIBwoeIDzfOZsmdT3AtIUw5i5kp4kKptjDJCkzUl2q+QA8GJpVyVuSHMvyDrdRMf6QUOf
WrKqoTeS8NodpQDUt0chvufdcUBQlzntwxoGIbnsdcpYQ5f+g8UoMljSbdZMqaRYHjoZ3vCWTTof
afiCC27cfkRJSJ9G8ouP9p4J2SnoB8LzqJfXm8XdNdtwp9C6wvLeZqUJPmflFHUAq5k3HEoN8FRB
kENvo/pKkvbkz/JQazip5NI4wGVsR2t20kKT8Jlg1k2U+HcEep8LLnAQXSTNEE90HhD/vPd+1U2e
mBDl5jfOgnrnxWsCV1EvgPV/QuVz0O3cLuT4dMBZK/ZZn6OQ9hUb/EuSTXADa7e5cSNyuI+Yn2AT
+/o7OtTPSbY07HzU0LKfbC4MbmjuuTmC1IMYop1IETEMSJ6fE0uimyUh/U8MjHeJkav3sEc+lbLi
ZSLy/zh0kmQdht/RvFXw8S3K8ciZ0EOLnJDgPNggpq12MCHRUa2yNfMyszsUm5aGx09WEz9o/Jfi
aKFEeB4BQ8vc7HSX70jX7TF4kDYmkVnPKPPLA+V/1HFMb9j7AVtYGv7qAr3qCZCGje+Q3SwKTw7j
PLlgjZwM+7+F6tn0Is7mGUbiaYxpE9/y1LjjJ+PzuP82phUkognu7e3JJ9ZKi4amETiBgSdTVe+5
6dJPhuLBu1fxbxwLWqZvwlJzgclx7OpDz8F8W+0GLvKAEt8/5l10c6PLdK8HfAh3ox5nvnKyL93N
ld/jOasWodOWpd9jWBG051qIUvH28IFoiuRHMIATV5g0+dtTRINs/gMKsm/HZVUS8rU0iJLOehWp
9jmfyiruvk1yaxgft4Kka/0nW7/rNS2HhArJKGjBovL6GZ6txpQWA9o7huh1s602cgVrIB/5bAys
bJaER+zDvxkcXB4d3UCTbT0f040QJ44a048c2AOWfM4fCwNQSdCgVQUsKDlnFazMgyfY4bchWi02
NmZA+J3w7MW2dALrmwMp42zeDN42vsMNxrYDpeY480auJ9il7Mx8x87j4/m4TBxEe9f2FGBt+P0+
mMoHDlc56GhF3xTptPgPFdD966ba6FvZwbuMtrYfr1Uh6RKtfcFz3C/E1kZpYFNxybf99HJoPh68
C9NNco3fG/WM4dZpFszICQ/tGexMJuQqkk17poipns+L87HgF+gxQB3y943oYOHo8Jv7G7v5Sqdp
azPRfv0aFWkBG/le33cEAmmpn8DcKg8CqdpXeOqj8JPv8Ykyp1CPidTPATr3xdjjOaT4hGrBmQo/
lJTqISpINsGXh3XFqDLv4aAwZsj1456jX8tLZf4ycZZFReCIXqjHAy9+QdYG94bjkfOY5R3aEUwG
kNnKV9SI2DRT8Ov9+RcDzTuflFlvbPmJmiA8QdNYfJMaxJ2+pERODv7tei4132TzONpHQohqwYdp
zlqS0agZZfYItD7Q+Le5YHQg5GTWDpCz9OgVCxbhR6XQyDUkOJj74cfWHHMXv9bn7sGKHy9K4sgj
aP3ClnDRY3T4pBj9zdL59BEqs9TioNox9P52wckieAnStuNi+Qfid2ePkFf/DMcdxuJmn9r4Lle+
g8ANhC/dQ18JZysH9sTC+lR572OcRPs2VDqBA0y8lKNmXk3SyHk3FnD5IvIalPx5acoADv4b9yNL
wn5LGHh50hBI6l1x4LJ9LVYjhilnz5e0TDO5eboELnJ5BUhaOF24vMxSTXe5yml7HRpYFnK/jELa
MXoARRDFEyuG3DLT4MXVD9LBiuzBCmTM54wQF804CLb2gaPPmVFXq8BQ6BGNWlvKt2ZeuIdnL9ew
FKwCRE9FFQQE6m47/S1HD1vb0dF9OCmliTz2iAWYd5GyxSZefvfzfBnVW4PWi8cYj8vGYnaFKig5
Q+JoBdmGhiphnpLmqUnoxHio8xJAao/zewyZL3YFPT4YHdvWyii5993oKF3AVF/5XhixrIJcEpoq
vOrWKylDhPX5+sSRY9llRgpfkpG6TuP63XRfKphfdqN4J6kTHtwIKOzt/PufYO5uLDYDqJTxpuSO
jJZmfGCQZOTd0oaYyDTnPeWH3f+GNF4aOZla4nL+cLlN9+JbxcGu293HsUy6hS8bUAJwwi4OiZZm
ovVoOnXkU5h19TRhcr7U/ycB3VcXrF51sr7il76nagWOiIzjMZGPF3Lmfg6ba6qbZeTvbKKEksYR
lq4pAY5S2oslrAaO9Pkg55u0wHlFX2Lqt7Sb5/hrvWHD8gOsmerW/WBDwL+MGHXAPDHNJhzLaLFB
2fBW1lQrYajxHTtPl8oB0Pd19XXI2G0eojTUGucFT4Fxivftt2lKSNyXFOKm3DWj+cakNap90Erx
j/sppAlhIkcMgTP97fbgqg0QnAK/sZzghP1t5avK7DUoJfjH8NKTwtpxPbIKzHgCWzL5igy6uzY9
Lr9OmJmPbiMyn0Kw5nxTq6Lzohg1xIaLbcq8D3badvJJQt7OfVWL7DAi+YnesLjq0Cs3XvQoUiPi
ONYknhM6DJ4ybPtLtaOQhS/SeZ/NAER5lx2nUYZ+ih+yRgf5YqXmID0TQeZB40k+fnYD82F0r2iz
DwODEgPXC2mdrWzCkxzD9hbNTBMjWjLKZ2YQwyaFloRoyo0TrELZ3Y6d6GKPldJlh3CI9CHiLS1m
VaDgMfpilVXepWeH8N1GI/zIopACTnFaaxatJMyEjvmIYFnjJKRTC9DBwCxRX+aZCqRm/KHLH5j4
J/ngTrAK7vpUZo2JgXAE/Rtn2vFyZoIC6uv/eJ6f2BQt3Sx6c7r8FU237OyDGunrs5diKWQzYHxK
OcEqlR4NijEvNatuqx21WALxwqSXVOZblAVB6NDIJQZcllqkLTQrqKdgNqJLXQ6RD6luv5xIGaiA
JPYBsgl9+sZ1wBa14gQ586Myn+ouF5PKsezluZJZelYIzjndAoyjwqbXoFvcxoi7/r66EZjYL2A+
YNITR2DXdjx7gr7WaZz6oNoQtt0VO/b2SvbtlR1nJmx7VOsTPT+FewBrYxS2OrqH95YSyi92mVaj
JVKCndA8u3Ctb9G06YHzTxfOikZi+M+4I08SrjXELURGTi9LRnDFbcUiU5p4CC1S318yEeWmGGr5
r+NBYojUGgYOjLB4LYvZsf3CFu2Bv+S+MoL2KnaUnkwWHsjaAcoW2GZXHdPwTP16Ys3zpnWaNeZG
ZnqPDc4on2CE8nx0hCyKCU5/3/fYGe+B6eh7siTm1Rn09fFWo+Mefs6ltQfXtL1KFOKWJ1hj+jZd
jtrsuCn5KP9IFW1FgHmOb1f11hqcGMzhOlJHI+9V7rwo03G0V1M0CnZAhIUAQzPCBB9XH3u3hYET
45QP8IA3p5lNrN2cXUMjOMU4k1oeXCE2VF0GQSGALxYH82bfueYb5KsOydWwFo21/heQK0dEzHcR
xR8Lq2+dWBB6T7D2741y/J0DJe1/JANcB2aB2eUagqUahVD4AWbBfi9jz8jlbQq6OQKgwPvFoxZC
6WWMtf2g7X/WfJ28kXgV2IGKrpyh3JQ/F3EwrwtxML4fqdbSLXsCyR6QLVrhee2XDlKK08jmttp6
s2Osiq7I50whgWeKv+sUMMR3+brmNAN0cCE3xY6DCg8KCCkQFuO7yRCIsuh/vDL585704eMYqdVL
8M6EfbTdgI8Q0BFWaIe5HhAX0zJLBx+CJyTP7/pJS39PslbGczVU3mXfKHLg/4kTEEIg5ghfQCe4
vYlA3Kb8y66QctHsPABDrUW1InIkbwW5ri11PspvqQCy6hiqyYW+l0zZdp+IU68x3aXzU4aLUjLz
yCRMJ0hHNdiW9rv1F/VAfFV5Ez+RLHUrYyUcMd5oUHBkJo7g8hvxepMaHN2VuLF5qMnWiU/T0Jkp
iKLRXMTa4b3rYAiF199edRfV5DzprLzSLWyRm3OlFjBZm9oBzL5iW3qOyV1vjJD4Q9nrJ3e1HN2q
Z4d/IgH5s/tIqVaDy3J6M5rmPBANfcXxgjzlsH/zG8PxIre3DmislV2eBAqOmpeha7x4YqiGv7Ir
woOtdP+HBx+YbsqFO/uw7VVaYjg+qQADpkhi9pj/2EZhlZuTH16cKvAFP2MpdlIgz4558qU2LOwk
Fc4DBcnuWFgDBWWMHLn7MhUMy4MlznrYE0rwrhQBhw1nEq6OvkpOrMhVubbvYjjo8gmDaUvLbLG0
M1GEvKdqO3FdgOqoC2y2u4c3IBK04wI7QYkL4j9SYLDSn+kZDuJzAPUQtW9+2+f8hsA6ElOi+24n
qntxItHWNgG7Xn123VFFuFzFzNjmY/Fw0lL0MzC0i0iCj6zvyx1/43UCVl1WMzHKAuPHtkA2eRAb
zukS6Kxy2IzItq6bE8KGcV4A+g+T21uYlmo1zftuGXogucj8Ie4AhQYGE6WgjgoKKYpRZyULbO5r
70+VcxALzrqZaxb8xgz+2WJQHu7zYXPUmF4Ws83eWjpOHzChc9COKqXU3j3a92zzSsJcTWQ/1su2
+ON+n/dxD4kHL5BhqyXCg2JEYlbgeEpLs93aNtjNmn6HFeulMQA4jSKeShpIoIjznd4C5llTU9VA
YdiYH+cEQBVOcri7PU4q+juiNQ2Tw7Ewqdni0hxANn1FB6Ehx8zHEHJe+bio3Dk4t4a51FttSInU
/wZ9h+Kj5Rp/hPXo0XueN8jK91FEAqQCHw3OOh3nfn6lwOU0qfEjX0bC30POB/CDMImmNhqR6ney
P26ZbzBFKtuYQq5zmcNfhNDvtlA7rryUZ97dPBiMXiKd4gK49pQzHSLbIs5gib9fQJjt4K88y1z6
wpTKQNrwGuVT5lgyM1inZ0NZgV3pd2g27H0uGUkQy1vOIfimeoanMs+EqEgccf76cwodfu/LyGHc
2gMh+7CbYLvA0IT9I5VEjp4IAblYTApz9MrPSvXRLndfTjgNJN3jKpuzGcElFWnKEcklOXf4doeX
2jc3XnHGw6V4eCyLsO+dgwMU4164LiOA7obohdm9+CbRh4dGIAo6MRvlBOIljBdxnpXg5gs79zxE
houbVWSZ+jJYK5lhtt1RKEzOc1EDLf9FLWos4xxRdniCDpEjiNKKm0jvX+tsnvLGPlb14JQibtjH
Y4J9zYBhNtaNvKfaprbenjbwzjxwcVavuJVRBAIRx91Y8zdjPNJRleyDwutRXyJCI7SGEFgfGdlz
GHSx+Mm1M1+HCVd890/OZRIBIaEpVnmVt2/1olNaUKHVEudxU8kIaPfIS2ZYe8enIySUhGluexKd
nIh1RTuO32Mn/lGh5Q9fJ1d6n/eGS0NVvWxS7mS7OpRssV1lD2NYd6fSF0bzAAZSQbvq7yAoalCS
JjyuVrU3pd+65B8gaDZgX2FklzhyCwljrH8Aq0WtJYvX9BigQxQAPG9u+QmYWNLcH4NB4KrisnGT
yiyCJKm1mBcIfYbXG8AFDPswWOXcw2fORcBX1hnMql5fXmHLWmBI5OtpQ2fGSbsuXLC5YirmPx5p
K3mygmJguyEPjTW6N5viBikk6z09FUVXBCY1P5I2OOWVFy0FCr2wj0P1m3+vlauFoy3GWmoTxo9d
FYHKd5etAnSk4Uh7QU+FOqllFuhRmiehdZ7mRXmo5vumRSzVKEGDn/mF8bYUlhkjaaB7j+nEIyVz
0tigXrwih+8YUxNjafJlEGdw3N6VJ9lDPj6SyiFfDN96YXqFjkhiklYkdNw9Dw1DSW6zUrcGHlgE
XiDJOWEFUMpGLunb4N9BbwRI/DW6iXhYCxkb7ieO9ruTtFp6vBkIQDwqiC8aUKo3e95k7+hYPOM3
cxwBASdrCVRJqIo+0UY8T28GlQQk24/SwAr+4NvvwDA7SitBhet8dT1/rBAPjnclIzwxr1juF3LQ
6+qJFxWlFC8eLICtD3sje8PmdxBj9XgKB4cdRSIKnWPDb9AyHxMc1+FEOAcxixfDgqLs6QcbCAa+
+Aayv6rR5k4BC58VU3TU6QhCJlMI2T+1YSVbvyv10pvyjkrnn3afFgsNsmJWDAk3TTwGojlx5qWh
Sh+mw/5GlMU/ZGHafhWMdqdTrlsNPZL3ps15ZDnXrDtpOXJnxxSncX9CAQGIIW7rhCKZNsujzxDm
rSpZ/uVIyUy8S10cYphgRiZNqzvw3KIUY1oKFmcUOl7fQ1wa+3VR1WNtJXDJfcDi7VieMAjjPMXY
32A2DCK00696xUZZk0WxwGQMAQpBA7GFgNUI/dJQH+qt1tVjIi1mqL8Ltm3z+moF5blMLmBAP3pT
1GMwB5IlLy96xhKaAic4SAB2ZILaGKb9SVo2h+kTYA0pzQSxGv7WHKErHI6sTYcVU6GeqT57AWK6
TeS/rVnYgdMpPzHiQwWwQSlzUaaFJ0D17UedRX4Y11Aq4D6CwVto97goNr8rq/BIOIbRvXyt9EY7
8WdlWA6MviVIz02j2xGv1YtkVsQUgoL5MwYtuJMKyDsa3nXwtsAou2YpjkCyZdIei6wxF7x/5C60
jjoepbkQYDb836wrGZzNYC0Ld6GO4BuAXRQ7JR6kG8qKVjaOQisK58Xobf6qpO5le8FY4H0/lV5z
HOfcW8p29fXceFTOvzyjsbqAmhk8NRmcHaCAVp1DCwhGRyHrWeeGVj/bgpgLVZ787FNKiMmox08g
SwHwNTix1Ll4D1DfR6RLBJ+f7OlkeODVTCd4qSJIkyL9QJlaLmcK3+ZKiLW5uLAcV2g8621MKfA/
tD0DYRy80w7zldDeCt8ENQn/dpDpqWdUt+TwT2kpNxtCYdLscr+Q7UWQ24jy+fDpzMRrdHo4AER8
MYDn2eGh/7D6fc+qohpdNofY7Qj7SOfmDeV6TPimosrwVkJhx4dst1vK6d8GsGt3RNByxP6jgULp
gr/CXeos+iQIlB82I9kKCkf0bP3jIaQlOOV/ooj7bKxibRpk2/3Mn4L1Y67ZXT+4h/SUUe+CWB8s
rZMK7WxkTUwMCqakPcgqSn4iqfQtDpXsMv7aORnNYBR47xqXq4719ROfWjEFn22na0MiGS1S17eI
V4MEblQG5n24w28TPFb1R/+wgqi6033Tyc3kvzvIn6s/ObQZJx0a1KxcKkGDxO9BIXQMnryUed1w
GN0xwN95vmihfXB5H8u9FNnpqmU7GV0mBwu6c5TePNRqSYBHK53Mt60/u6h9Fi1qO/XUR9kVpS4l
nRNNG9OrvRjIOWYxQWyNJwOBHWo/myJu5pVHtQwaU+DKrqZcc3viYNKTCutQosciVmcQJzYGhDCb
q6qyQ6pOHOVkV9FHjaCxr8fgwaU3AB5oBbBAoiMyR6oaq5/agaHfAWDDOVs0LPyfUKjwVx4HNQpW
ueacXiiGVnfaermX9ovHcxf68jZ321ezWMduRijxwHv02FlowfIa4mEJjWuiYmcIonr8YqJ/egKG
3P5SHkGHS5EhYcFmM53hLhnjEkz4+uEdMWQTn2h78b5gkAwdFHsyCz7piUY2bIkNjUhSEfzTZyeY
9ks04ibTmPycLJwyc+W0jgz1X+EKOxaI424P1O98NH5sFakT9x/YJN0MJ5Wj2IStS8tVpvKBo+yK
CdlevtJWUHx8goCKth4mEf/ocbb3JB9yJDN5yCBtu3Ebly01fkHQ4vGDq2nCKRKDbCIukynsv7bP
2UNPmmOc3IarLINQ6kPaPK77Dz7qoDZoFcUaF6okv6CUE+HIXWzONpog/Ek4O4/F+AYE4BNVkONy
xnQCsQ3wXrgJM0X2KJm7yjyHZgDgj7j+oTjVFuSV9glh8HMyPBMWutcwVW9BOpqaiz03kMou/yMZ
scCZyr4QBH6vb25+hElEC/eKCtw9F7LxoafX5UvD7tDFnz194mvEK6FGCoxRuiwYuWQCgpWx3RLG
qvhrSXgYvyFR1wYuTQ7Hhky4sahnpdlWsJvcn1T7X77H6+A/O9e09LkfBKJUNrYiouyJbNCmNzaJ
zLaq4Li833WH3U0WQCBfIFfoFd5SgYaVG/jpifkQMKfS6W1WsOliu41fPmmc88W72W+CMGRjBXT7
FKnTlDKGc4pRZtUU59nVqnC1fPXaMrpYt4sjZeJcWQkvf55g69eYs46Ol3NaD/0lLzAZUkHxSXyK
2BGXktu+vszXBrQKN6FIjX+4YCXhNHWn78LEXL1uwLBniLZAONenzuZsb4YYjYOiCAk54kTug3iV
e3MqrKBxm+OcK/1CjxmaDF/SE3QTXrrxN0nEdone14Wb0PRjFJ2ytZSbn0taP8t0p5NIUs9BF12q
6hfUYaQa9CsnCS72U8p80JlKKTFkKm3RbB1kuhJq3bGLcBZnkGZIHc4ztfkyxEGXOg6Iu26H7IxU
Mz61RtbqR4BeNiraJPxgS3xcErK9cIhrQQl8GoOFPPOcgJNmZtRCTdWCAKjrYyWbYDUj8B5b4UPS
PZXn6wnssIVdvvZadijUfrSikByqV1fVUChwBJK9iIssbums73Hn+nC7a/iHh4qtfU0icDA7fuNV
jrkgKxwqtb8xBoerRkrREzpYQ+xKZ0zPGRdMnqfg4yD0gh557916y7CuODOUWd0uMGpI57YcbkwI
BfzY7V4H7eUEffgmGhpUDoJVT6DKnq6dFZ1b3gTsK/Vrxq2U2LbipIIZ16RDRvxEof57UbIeV4uL
tI1S3W/lm6Pz7uYrheq1M2CEOkWQoYoJDzQU56sFW3cPjMk3U2AStLF3Tcs5t9HlBUm2VqGSWt33
mcvo/1jKvoJw85ujtLDUr8c7PcRsIWKpTp2ERKeDvK/lpNDsTbPgyJ+eA9e5+mJb8BeIjMyN58Ks
mXZL0LvmsvqXLSX87jFkpm3z+pm+WT48wHHNnYrDCJu3uOVwLaaoevykKJ4/FntVf6tO3LD6JYGY
d6L2Sp54mAlvubIA7eBXDng5a8UDN0Z3aTRT2qC2hW20BV4ncIKunSRpHoE1spO83VywXhZ7Q8H5
ihZGK07KcYpTkC0R2+Rbbft8UkBFkGbBneaZ3mdHNxNlZhvSpr1FFenPBlmIeLce6bqhUrzXwcQR
aWHOXj52cxZVill7DwDEjlR6dW8qa9hmydPcSghS5LlotMsi4ZXHT+g65zIjbP4biL4EKThfmfo1
Mb/GHspUfp0/jp5O2egXj0FO0EttQQPqGcLBWmWreTzmcx3/+Epts0TIbIMLX/M6QP9qwBznT9ZM
9hqIxZ+iGni+57F13aGIYDV/iBzQepUgdZAKncHONn9z+A0xTcRg+KUUhHM3xHTI2hHY3x46NaWZ
Rmzn4BO0D41WGP+f3MiERUPtRLZjSUttpxdSBy0ZJYEvbwqAMIFi8JzpFoADK0ak6twwRrvii4LG
TVkMBCU4Yi80p2KaBbmMczMR4xyQ/aCHnu5Pv42kQVcr/G50o0RE4dTqBNUFO4XcrETIvk4E+yH1
pk9cXfcwhxnilndLm6kWixhR22pwMD+vc+5HKmRh6xAiQVcyvQAuq9bP6kOeIEK6PhzZWcxHe8F7
RvZ0SHu37EKOZkU3x9A0uTDYhCKQ+yNovfQbq3i8GCX6ZCvWFHWQqdyvA+Qdg+UEoDzXaxZcXl1U
dRca5mvlclEDXusKJGKGY2JooseDbyoTfFuCUHfhYpaYSjfrJhA6K9bid1o3ZVgiSYCnBSiO8ksO
HgBAx1AuVr1PobDs6Qie7dFlTjt/Uj76bT25FN2eR8MA+8iiv74Zw1OuYpJO+Qxx6RpOMD99GQJT
Fq2bLzDGw6FEeXOK8njyMohnS+O7wTfXP/XbbrJ1PaZpJiaX+aQuraAvijAL+t0R9hkJiy1bVCLo
TMxTqqSGVxX+QH76a8EfoNbhdtw7t5C0T48onGghxP/mv2X8yVc6fWzJibrUHA7S/KgUftHcoMys
oHnKpuu3I4Y3ddE1Fykcc2PunmIKZiRvyZh8YwcRfIA3XKFSNGUnUaidEeR0RVKm1dNZCfPFw1sU
/DhBWxVmj9VCfugfE+Yqny4bLndMaLGU9Y/K5Gf4BCPudQfqY8X6L4kQQC7U3s21nl5qllYy8O5d
x6EzhlfvbqlQjlm5klbOC6Upk4lhbVWc1s7Eu3HwyvWXR2KybmqPL22LLFV1/jezqH+1KDIuozd4
G/CZ/KtS40eCp3o1H+gvg9WvM/PQlyCXo7b6MfVTD7+hHC82j9pAaR9Zf9srZ+DlmwdbxdYUq5sL
snslCdx6yBF7vFbZQ5NNypv5HY5vcFiTEdd7TUJvCVNk5L/u/Y5ZEwfaXh6Zjc95vVTeqPgyY6G7
TiK3Qk79ub6jczEo6yx38xbiAK6DICjyx9QNMIUxcQP+TqtQ+A5C+vReKzdwHAm6K06iLXyj02NO
719E0IRU6yMN/tpo5HZj54mgQNQjkOU35ODHabHwhktujZhw6I3bEjdwj3iZiMBzyZ7WMOZn1JqD
c6vN5aOx/6nnV1dvMB/eFRzoqpqu3XNN8X/74L6Oy76Eu7g376bTd5aZWWHLcZxYXGrfhFCjKdir
U7RszVFnmVdgOTjHosqc6aOxvoCg89sEtiM1V7B/LCmx1SPucweuQNDcJs6WPPzXSjUDcsGaWRL4
N75dJW34ZOv+ypJzIiqZofa0hPcg/N44peT+1IjuJ0UBbI7tNtYUne3R6QrGsaAsbHEsSFrjydux
s0lFKgotJda4NPYEHM5OxovhOZgMOZh8xqfydMNpmQSqnYVyzduBZ7bHR48FRZwNz+oaZ5u7s3kq
BPrBUQ+FQIehuGqSdbkCupVsc6w4sNMiXASctsM5XSK/+1Ysjyy7t51PkEOUYFp4LHFMaJUFIr2n
pXPFj7P/owApOAK10f35g86Ls9kSba6hLgISF9OvVDOK0+zcOOoJejRBkBORR+bfVNEbZkPYgQSx
k+r0VV6Wa9Fr+SVzvxgCLrDKGshNj5O4cc05dduvZs9Vy7jYXc01E2c9Oy2RTcEANrgKNu17bf64
o0ZCUFBHXzyqNZ75bGsMc40QtjhpMOBuheMdyGrfJ6zXUvIbLrcLEsuWL/FZCgqESOtWDR+T9peP
kIc0zeuQzPDu9dAAGrSGAzMPpPH+7GT1BnHhtWmT0qUVcAJOq0LcV7JUoBfKbae+OV7HmmkDdB5e
bFnCqgEkaiH4/FIlYr8ZQiRC5qqC/wiuKvy+Fa0DM8knV7jPsSSNhvrIcPRIlzACJVQaGP2eW0yx
Qo5NAXU5gbgK3pmhoT1TJUfXw3NfT4Quj05ahAK6PjdX+bXVZU43y8zb2Rgqr1lNo3ajmkcT8k1s
00tuveeXZfmONOoi73k0b4CdkHpReDa0a1SQQXxKRz9XKw3KvUzLeWElYaPmito0RIdjNNL6dpE2
5HxeVPeusZwmshnY8fPTqQx7KYiwco1OPvs154LdJQmCgjaRUf0fuyrNAmw0I09BPJa3x5v1cqun
lTDEnsJVQpndWE5lKNkDT+JbD7AcCKmd6VVsfytoJV3T4GSRcstL0H8sBxNw44e2Hbzq5vimxY3Z
0Z0noJMoG+Cs4CCKTDnLU3u4+ODB+E9V2yy1iFmh2jqUOzbnHDJwVDqYR/w+JxWE2bIJhikC69OY
5Pd8EIlWvgNLCO6DEzsWBDE9hF6CewsjuXtpzEE4aii6WHeTr1TI08ftMZ1U8L3NbWVB/4Vp/sx0
HVcbKZ6byWXixp++5o/+rH7JXs1SKJfPbgHPtWFPrd01WaJVflaDlw6u2z+61zEQhVBImUQWKgRL
fhK0pzHGYECznzcK8vgJzzx+6i8VaepDNo/iBy/wFbZMVJj2rk4Z0Smco1MzOEqdHtMWW6hJRLzk
ewBwh90p9m//8PlRF5FflQqVhK251Rb02CJPl6Xrusqa5sCzPTcuGypuDeFygWojDkr5m8RQoHeY
ngJwOzNPGEJbVfFwbcBTqZi4pe0NEgNI9BcGRhX9FYbe3bBstG/Yj6gz1dY6CiYw6AwKYjxduLju
15mSEnpF++kZyZRSTwkKB0d1CB4cDnsYFxQhrpGDGrJ7BdBXlwwql+tACtK3isgZT95v7dGCi8gz
FMZQ/OFRsWZV70K+071MgTffOwAb7VRxL35zG74D1sIDc0VjRP1hdOlonnVG62WGpmFse6HugBiQ
doS23IdcmfI+wcW1XUAutKuH64eiW70QUF6tpplmI0Q+Q6e2kRicXJtS8H7nCdqPBOM1/kbg5i5o
Sx6iKeujgE4R9fVlEmJ0Bu1C+LGUulbdYRjPbeAnH5NgMTHexkr5jlFz8vcz6yKr3f++LiwRVMk9
aJ8gvJ2C3DPbwElsNfIdvgPSY25rfLPY4pKhzNVuvUoRC/ofhSnGY68eV04lOFbKoHEEaWvKursG
UQOOKDDloawrL1mTYVsyvhEx36HUCWKGb0KKDiwmOzgP/pBtH5EhqEze6bLPs7ZQK7O6QS3fxseN
kZfj+MuYle/E+XFwGCYJazns9nVQgnEY9TxqB/bxnZjif7U5quwbZnzH06PubAteE3rfklnmqaqG
oRPK+GpqW8Q3v0lq1hpifVHBlc+WHHuod+4pg4QjkedLmd9GMfuQqeR/+PovOjxUYiWFgCb5bWUD
YfaETYLK+7W0SOMmCaM1Z5uLVKjdtA4JA/tgVidNjrUoL6DJ4nlBH0Q91SKFibJwH+rEZgVI6+Jq
Q/MiPgNUrUvGWkYyh0x5yA1yUEiOL4eFFTVS5EA3MgziRzQO7dXRzbj3o/pIGsWLojCS8UfNVNyp
g1BbRAxh56ATMKSUAPKusCh+1+RQcJ65bff6NeHXKvyB+b7eeRlsINHBwlnPI+Xx5B+TfpFse2fX
Wy+tzBC1/17s862NkRVWTg7KA2kSCSK624+5063lbd6R7/BeLQtY2xJf4U3lvi0VkzrjQQiw9Etm
S/ZftnMPnvsHISHX5/9fA8HyhAq7uBOwxPfpQFYRZeI9HrEl1hI0xq9pJ/WoYGWFIReQsHP8EUr/
+tHTLzuYNtZuDRPjimZl6eYBPVRHriQWQiSv31/y8+k46fQMdXvxbKY2IlBckGUqkx7gnGMF1uFQ
N9d5DYk2oj9cokLrTJeOizkgoN492+Cs0p09eEELtWe3IF6px3r+Sco65MvCsFlwn8CXqjlpdndy
2wh8ZqnaertxHdXqNGbuDxUDOe1JpHJQTwfsWlXAfYDVcaImXY6Uswi471IF+F14j2NpUscN5jXw
FQAeqX1eEUM32guEBin+dG/1NasPjCqktJyiFUL7iTEVhmAwJqVQsoN4NcNvllJJ8z0sgS2yZSLD
jyTYxGqSU6dFQY2a1Ok2VO0WmqQWG/ugqMmBtmoa8irOawzgY5Wd41FvsBNSMYoSz8Ts+sp0pLEN
vJym+9f9/1lXQkYiTIPvm/5BcRbA4CHBUZUXCN8CqNwQbQlYJh0gU/FUupKWqfMnAZ2TUEMVKeLY
Y1Bo7jttcVyz3wgd8dFXzdIPCjDE+AkAML8lyx0rH33DChbFV3FFIHVUzAG8L42WzxI/1zrwgd3M
6tWU95FSKuItSQksKF7aFFVZp4Lm8+VjJgIXr22Z2fJGZRE77Ul4R2PPY/Qu4lkBUihAu/AF3v6Z
djGEladep5UdeYC0MTdgNOwEgvh+zC79ls3gn0yRJpsBWKHR/1QejiCPktsf5gyNi3aXXwCQeZVw
UtcoOqID9CHsTkLFOolFtiTeSzCWdxgDBRTtqQr6IzqXT8WLVmBCw9drpYb5lKGBKostFUpD5cbc
rEDAy4OCbJEAfJo+FUNHRy2YuSqDcKWPhOdMEnnFreWlj7sqQ3zRB2fDUGD3ZJEWkgec7BzSZCF+
FZh09j/70DgQndw9oKXQcyGp+5fgKcCn8WLS/a0lCRnK3EKyQTBQyTcIQVGKsAxYL9WwkGiEaqIU
cyNgxazFPRxbUINPJoc8Kpc6CO6iIo1MWfGeo+GW15bWPbAhkJ9wRqtUVG+ohDW/Dx66Z1AueWhX
tbrGeygnWTnRdm+W2Xt68ml7m6EQfOoDujRu/EAIEBhQdYWUXGKlKl652h1nKrFHnB4W4dkOtyN3
uct38E1Y6SFBlEnT/RipW3Q2OtOHBvITPVDJddwb/C0jNiksbDBkds4mN773lh8gZqpf0c3Ce1Ke
QBmgnigi1Q14GdamLHXgz6P166lys4gNihUbNwzHQLDn2xq7cTTZHrdZHWV4tgIGb9JwPXQ6KOdm
jhXbtkcaNChR8OpUZUIKOeVdWvePjTx3SHFl5X82dDQWELdpQypQE/ea/hCAgcAdfKPGpTaeuiDq
X25cunvtp76wAcOTcfhw5Em3ZAswUxGweogoaQrQueTN6FiQlYYx95rg8JMf2XxoGEqtEebiNkjn
2L2skJmjC2pjyYus4sANlYKYbFuY1KsbELPqdHawKMgW/DrZckHJM9nm2sMXYHSa6IeFJmvNR7YK
kSR3lUBY/Yk4erP7Zn2817Me/arYewSsbqcqwo9Buv7jH9SnU4DCizagvPK1GYZHkTcEirAVQKMU
iKNkAoeFXmh1yKKc8HyXuVJcK6NjPI05LZUbeKX0j6yh4gTVbNBMnwgvdSP5zydP4x/PHaNLUrJE
0lkWG/zkyFxSFTutW1F6ZTZcW2NIizRpEUqCWG7V8fr3nmT0b8oC1PHBO6cxh/Ptpe0irj00Nv/G
b5qY0ER8kzQImE8B46n4yqqoMYqHZ43h8rUQ3ic4Ya3qFKLqssVea0TQAXx7b6kAgJDxGnj7Q5m7
PwjvvTQ0gjzk3f/rZhLcLUPEooASeDH650y6wGcraklQLfY15tDEYxOZdeblAi/Ve/GkDwTvC3da
8kkb3xmnii3jfFvAapm7n1bh8rr9eTmiD0mM5ChKfvc+l+vXXNJkv4YZoMvWtC3jmuQWzOzoKjFk
M2gUuQ3x7QDJxx+Qi0Q1FftE2e59+wMiIIoI4Dv6LJ/9wSrobxREmWlVYTaEsL0tP8/oBRLbsx9j
v/3gA3+beVegDaw3AgQ1ciJqMQrJ2du5TJ4zS6oHtN9MTmShQNWFcCBIRLwy9vowqqB069tAvNmO
vA3El6GByc8QKa3LdG+ablwkNSo4S5Y9rYVYUdrXiy0K/sPT/cAhEiYZ+yR6q918QspilaT+OZQF
LZAzTt8DjgIaG+Gt0ua2OYHLZtc1Jh8tdB7Nc3dZIXcsWRovTXlRawz6fG9uD20Kxb01CAL9B2u0
2e3zZkmBQ1QkGOv20lhn1+8W1k47F2jptGWaElV5lC0c49jSSDcQff6pBi3Al+NDDBPPh8OqJ096
Oznmb0IXARQly0r3Pz+2XZoFcRXIycbUsrPcTt+WtetOUj2y3tQ892i4FZJCLtMwUlYw8Tuibw4U
p9OMPbeeKW+6fEYyjwWF4cVNNesJmxb5TYATWPWcNJUUYsiaFBnqqjDDvLPEwJd9NrwSplErr08p
JPmQN3lObaTLIIt60optKG7x5pX8JofVoIWsTWMp+GBc0sK+i8JeXkpZ4kWRhxdqoqyzn+kRZ8Qw
e2hbVM1sxlXT2cm9yfVm2S1ZA7c5wJNZY59Qb/9VK4LkgrAergOLCX2RE1y3AdwoMxtUq/tIEmYy
Ake2YJ40hyPaB2CySgb8Pek/TzaXAhwf9Cey178uuQ1CbXl+iWsjPmxJ5gAnodtSgxMOlMrF6BJ2
2KFQTgSwityVV1uLH3CDJpAxI9ZJa4Yxx9S3nPLcLjipdWyFnElYZ6QqsPEJ/0PJCMp87QiDvUzb
mBxu0Oao2gIfwk7ddWzsuPhBHtkpu739AKEdY38RjikmcEGjgk7c6BQXRC1+HloVY8oxe1BCGY20
sQm0oK1TyHpv+HEGrBLrj+H90IjjX2C+L2P9bKwwPbN5Q8kbmEuInXVuwhAdPB1M/jF46KshWW0g
NJ3DYE6/JwfWxFPi3+63fYAGJqg2RBAAfiZlU3W+c3poKlPUWiC42WbaDKbrEAobv8HkbxGVtj1a
qKcVZPXkwbFqYRH8qWLfkcLxsuCN5ysiQmxi9jvP+BSC0g297eQUnFJyK0FLEmHle9PhHzgNxqJM
JnzXBYrcQAY7dzgWZcQpE9rxq4p9q7pMyJRrAvl1EFouQhayxVLvjeSPZ+qcrRAy08DYo5X5M0XY
bD+vK0ct8LPmn8nOBUCWPZ2GRLkg9+Bz0Tj7uHfdWKHBwrujasMhifyG3RPy5KghGsMpKSR5GcoU
ZeY/elHdKAAGVf2pcpuk+F2GJKM6fenBk0d6FOIgRucusrD8hE2WdBWyeOHdLppVlIT9LAs9+A3K
yF4oh0fFsUurCCeyZXbfZaqN4oBj4PEdICSOmuuECwVJCyHDcK/FYKt8953RyAVjm08F6tl2+70/
Ar+ODZxEqImrz6P4NqBSb/DWu6Yv9FAhUTJffkL0JsY4+1splELmiUBf/CQ3Xv1cDD5CoV6kmn93
6PexL/XvDmP2jw2RAMvmwve98zJAcauvKBUUIlAaCh83TqLavd+wDlNdDTu/P3PThX8RLVqlAdKo
Ul2BmmwxtnfS2W3AflgrUErxadcZrUdBxItbLghD6m8p2eu0AXbGKaBqd99KQUuwYj8HzIzZk9WG
pcjQF9i7LdiD30P9QlI2uagInFKiBMVSosRfiNeUeQhJJtBiDZ6pCVmYlTgZmJwfHv6bq/09ZgKS
7U+DA/dNrZ0BIe2TdCFTT+zr2sR2oVUBZtBQ0qq0YP5OyMytOCdV+1L0dcC4KuNziff3sri/k/YZ
tXQwAFVRJyZHSyyU79pxHc/O/VZBBxuec3cnfpwBYyuFEzDKCgaHm4LYVCB1Uy79BvzfRnu5lY5Q
BeHPBoeNa1dzmNVm6KRW1EhdCnybfZb96h1xgDIqajGKSzTrdpwqZDt1hKGF4J9nr8epwySBelp7
UcYjlSvBX71/3yGuI5900xEUqtPrHVu3PZ7Cs3HHZ/wq2+n4d/MpKZjK65ttRRqJQrDpbbKEbkAF
1hgsy5V1R8btMfn6o1wrOpZMnX2gKjWb9bHU+Lgad7J+I/xL9YC+SCH8+8jDeUAYyuok75/e5EEF
fAQEucUBmP6HdgNZz7nYigI6et4Uf9M32qNpDHEuU3q+adGDW4xLfLLl6sFPmY4FKaWHua8M/uEF
pjDzl6fUPk+0FWWsuJ6cnPF2Dwq8ywCviCKnrh7M4NTODLID+n5W7x8Cv7aZIbpJODpB9JVL7zI9
7O8AHjldQg5c3rNMXIe61fyjb/++yqHSIja1YH/u3s2CfTOfYELNQE0cIcIYzjnZUMjy5W3DOC2M
qaDbnxFKNQa5VxLfL0L+hvNLM8hTzHXtJzbS/sn1qxLV3aCltGSz6R8dltdJUpQW5vZp6+/com9y
KwZbK5qTklLra8c7+PCcfquWOIqJqFcu7wvtLUu4+xLQLIZM19Ln5y7V0Ma/8oLREN18C0rTl0AW
5I7qsW5YQ3EGX+mhSrtPCWY8BoNelqpaAKMhy4a8UUoaIML+H1QftEy6qWAYEgSQdviTVmi4MEe/
3QZ7RTm6Y35FDy/DLlLJJ4VEzDWmBrHjWeFhyg1hYcWV14XLrY0vRamurmPdxNgE1KdY0v4DhVgp
AMbTqEOSxaYbtdl+cKEfdJ42N5L6Bx5wCj+a2Islqe6GRUdHWJjCqhL+5iUCrP74h2NiGHQEvzyb
i0ToPE+x+5/UhAxhgnL7f0kLHCdq+0HSJpPYUsXCAkJdY4q1C4EFgOZC5ACGVFO2X9CC3zsIIehx
5+OX0g47269cDTuXYqQYgSbd48eLjP9NlVExescEEFGxCCZSUWZPbSRu9KV+oDSqvHHWY/Or4Jzy
/7gg2vH3osl035zAO1jvHELu+gy5n+IwbGwEGq3rNYtHffjNfuarhF3mazY+k2e8IA42GJxNENui
PNXY54oUZ5/qdZl4GSy2F/9wy6bCp0RYmMEyy0Uo0jSGTihFD3gxAHtl5M5bgq8XX9VvUG98APBj
5gS3wG91heVdjDk4k7a0HfinuLPz3TK9t9at+wQinCTBccKgalX9Hh1ZCItHciD8Nb1E2l3NXllr
pgaeUQIpNeGEtzvIvBwuQkxy0luvBy7+OHCnvZ0IbLQXdQm/Xi7e1ya7NkakORsV7+hjSfcvATnU
ey3eenemu6cRsxfTo9VeWFf6B/2OEGln5Gou1cgi/0XDfvSz7W9jL0N+HmABFvJAH5M0t0RHdUoe
eX8dnQkOW7i4BXF6aJSrt0rPP4Xwm0txT/ldLPqSCdWFmmUCNq7DVEh6zrCB6+2BJOFNQ/7cil5z
sXQZd6EFu8oFunhPJ2XfpDCwjZfr4S8p2fCfCsZYrM+zTqTpsm9Iswdx8Hpzwq8NpBQbXguaE89T
HHJgWxwFN2Duh0R2VDH8TcGQ9RuIXXCQfHTY+PYzHsVNA3KPsywJ4V5Gg9HA/mC0OZIr5tpllap2
c4IHbwyIfWc+WyUti3EPkwAVvfPorc46TVHop367tKEmz7qrLKbKt3he2E3XltWEprz8tqpvttZi
iMpUOShvp+UQImNfbsw8PDwV+xeoydoeohbebWGrHsaLNdFfDmuBYhnX/hSNesAfdmOhOuhDx682
4fZIEbkUonIc4kUC/DZd4PxOwZqOkpog2bBij1zootDhRITd1X4rulkjrgkNZnasWRz9dJOXV3bb
hUz0WfN9usvHhdo0j0jS/Df6v9vQW7hflXv78ARJpsO943bcs1ZWYYTd9zzhbV+8PKEyBOfjyhjI
5+2W9UPK+kAyCpeopg+iwnbSgwxwXGDjPxGucTvX8x6pPzJ3P8y/xVHITpns8Ry3C7j6J77tlZia
n/NRUMXzUCKRwe09/YVrp2v3Cdapw7fkmi/QAaVRYsAI21Kx8GSJkaCmat+z6QzTCXX+3o2tn3zw
YRBcWN5QyrfSO53IvUGUVamRL7ljC+0Ov3T2KnWM0mCNomjLkZICAbSFtK9GIkuk08VBEEr/X39c
QCujnRNiCamPKDeiNmkMfsM1mqVJcEB/AUOQN2i9sQWODNENAKp2dHAy9bj/DWusGzcARsaHYgFa
8xAFDev9xIjRGtJjxdPyFSbNTm/flI2c2Tf8bg7XQQcq+C3pSseYEsUHqx473APdPZA3oysHsNtu
QYsO1C0InArIlRH9DZze07MiupYK81JWKkUNgvisU6iZc2I/gzVE1DvpaJ9AGOvDI9L+m07s3goW
6k9dIiZDzORhEpzmZluUINAP3YGgoGuOxiqZUHoGkjtPi5yrBpa/Hek8PEjKJqQOAjVuzqXoqmi0
UBdHCMPYBA3zz6zUOFnrquUQDYKgc80LHI3EHhzr0BYM1CiScyX+E4ixlOCXxe9OS9/0+8K3/pC3
4AsbRbOqMhYXllRiWvOZM7Q10ZE9YH04FwEANfQ8arpH7XXoDJVNzZ7y03uqfk9G4tyqgtTyaW5z
d8Sr/il4WUKdASfDfbsStayctBVNQV4WjVuqhCZQRCA0hi9L66oad02icrHIt4v5RrZrw5xe+1Ha
LRXaH+1hoDDi00eKkhjb1aoADarbma1DqOeRhi8Hffo/MMjPGMe2OgZqW66bz3wvNjy3imwo+RWN
WV5GLeawenLWgulNwdMhbPTLUuF/A+lzFxvS6wgmONLgdihmqFqr21fNNGlyJa7brMrhx3XEGsyC
UUJdK0O15NC5AoQZuZ1NiuKLY3HnrHFUnQv0DEVBb+p05Wx0FPoWAICL+YqvPPOjB/BdkPx4X38q
8SFguMD0fxtUPnJu0r4xW9I4fqv4zdSFiYZRaJWa0oMHHmKsxkHb7jN9/XlBsmIKSp/TqLhwKNeF
TT5W/pQsXSQ3LpB+PAgkcewj5QOCpP3xuyDksaAGQStBA6FMn9HXx78XugfN0GjUk0pQSEiwyiFY
OdfpMQVUiOAMd96AaRYNCNG72rasahgLRj4GOlIa06FcKLYPaxurCo/uhUmY6NQ8MGEXhtpqKpiT
7IcISRHoJvTTOHwjQWNlpcj1IsFB+gLyYk25+dS6mHMY4+R/Ccz8LUXqs6PFYf7NPsQUBC4DMPcA
ZOQC7y8lqb5dayxhQ7xcQrZ6U3QAwKIytiB3FgkX7y8l3APIAS1HCsQ3h8TRXG8P5fLNdwTry46j
fGQNdiwL8/igQLqiyH0NkCh5yBFGVTLHOe/FRdfBiMtlbWp1ZZemYnROd4+0RHr7h1XlvlvyN56n
MSHc+vY5rcjs41rWF616/I0XidFPD3HYRPOY7f6WtMLCpE993N8RJ9WJqsEa8Ezw3yv9gi9bUu2u
kTpI1ZrvRJnTraN8m134Ue5Wm/GN+ifo+aGxD4TMi9PWK9tvcHAWAZ+sJc3uiKwM5yMGkNXBjiFq
UjMEuXLJwFHAmFIw75aaX/IQ/PL+ns2esktftbu6KHFRP4hHtkiG+nWlAaEQkUwMCvt5fUcHZmau
G7ERKfWVCeQ8WHx55l9JdcFAff+Q6MFfpYU1fGakGtLnKyrnXblaeMFX7ZnhFwhO7dTeE3Ofksxw
VHNI5uCr7Vu+1q7cuSz8ldrRaFEOxR/Vjolr9SBMYxDbcgZqlE2qIE9pt5pKs9hrNTNo/LWn8AlR
T5STN/7uJztboSCFHykqsIUTnbGqI/t2xGUEzPKv276HhjhEwDXnwIKRNRSSF0m/BqPddncvB8gJ
XXCUYn+BAlPcu/inFSElHGJgLn6luo+T3u4WN4d9DdJ59POH5gHHCptEet/gfY52eK/8jZ6dGeJT
V5/1BVlZ/SleSOrI8UEYzoWbjeZOXN5C7eLCymswBX0J2Gb/EDaFKLNtUY2I7obFdgXYCtVs9MA4
4wqo8C6PjQHtqvChzg1mLcm+uD5b8B+tQI7wSndkaz4pJCt+VItd2fmdwnEgx4VqmqwNGYyMU4Xc
8lYNhRXrl4/8cuPElFsln+eaf98esmOEbTgPdOtOdzMonKU9IULRwqdmhcSTXxtg6H8ozJGlrm4H
Y6kPXop3M+vcJ/uWOOT4SmdLGBiuzk7cYvJYlb7X10GmtHNoaKzNLkKEI314yiVE3FGfeJE5KNFb
4UeIMZt1d3wN01hVpZl2YsW9P5nrfJ7otVP+U4LdMVd8FTRdJOyKJNSnhCD45hqgTygMbP9jQHm4
4Yi1PKyx5xLl4TUyVmipx9yEnOZEeiUY61Wn7JpeDF5Oo3nYs5deG3SAMRZpoKpoTnAcIXOHklUt
4sysD+LhDnmtGAx282K2afwr0FOLEPhObOinrO7AgN/N5zTeZuuyX2VT3nSjyimQGPzAXtVjvkjH
BgfsntnsG+jDa0FOvoTevPhmWMW4VXRW4tha/uTkXi9sFl/LMHTYoGL0hIh9zoSm8cgHfnPEaU40
Kd6PdHOAf3h19ao7BJtDYTkoARrcLAgtuHJ2si4Bzn+GGdDkljZBbqVDrDZ9Q46kltspqfjPVt5V
c2xNEr1PIxDVqrfIdBjxdn6Qhoygc+5e0GbDOSFSd7Uy/m5WJANml98KV/+0SERtecwznfOVYP+j
VbZiNQ8fkHQaYgUTDpaUSSAt4SY61689zLqeOamt93ECqNWvDPbnSy3MlV7w1pLqVxSgz6YAZYLz
G+vtC6EMw+Y2fRQcSd5eTzzgVKMGCQM8vRxAxuodufWLJqHlY3N74IUaUSg5Fk8HpM6T5HY4PY9C
K0CvfWNxsZAqtYV8M4i0khB5EWh9jKe20VH3On88K2nOI0bPnxgu/tetx2BMOnShNuW+9iLnh0+l
Eg+kZ6LzsG01QY1FMASjKzq5VZYi7eYgQ+QDgmlIh6vN1hBdmxDkpmwSO89nshlRKgWLGghvTiYE
FsLHoSTCdsmm1dWmxofIVqskSDGovrJ/TADme/fNxGofFNJ2qLNnuGm1ngCmIh/PndwvWmc6MlOC
k5ox8WlOCq9wI4LR8V/qd/fhuH0NeW0UlFQY6ieqnHakGwW+8lXbEL5L3h2pTn++x3epPrET/Z5i
8BUGznCvS7v1RqYrqed1ig9+zNu1vnbeEiGooiB/BY+GOmB0Y0oDyztsPl2BYBF8qFYkJjUWTdPQ
HVn0LUlkc2nla/Oa+yXeJ8U/EBoj9NoonMOhjqZg+3Y8nvM5fEFcJ+fB/a2fvKfP/SYZFlq69SKK
JOOtNVonJ0Bfx3z8CvYMc15q3ZQc8/TS+3zrofom5Cck4semo/9XcYpS9kGs/DncvxN3V4WtHqfj
NA3ywLLVfgiLrIPBnmUkRXSWKMwH8d6dxWrIG3NyR9wI+dYsaPcr+wFsNnJ70Yk8PUAs7OzIpp66
+g0mqk1Qd/aFtP+uXh58vs3R2To+yn87JAbQCM57V1i35cDHLPN3S/fHBIMFExuE1UjC1UL4j6wS
JXV0QaswOI478lnaBN82b0oMzs65/3D9fSK7Q6so/J/CtBTZKa3H2HI5uMntPaWOvSECJBfLcj24
Me5Wyhucp2rqo0Zaw0HJn0LJA9+bxBBlWhMxBxKloul4aeAc7EQ3bzneVPQ8Akj80VjfExCbBa9M
IwJjv5JuQ8lvqul91efuOsayF7R3cRea0JDh8hNPhlcM6dzeg9qEaC/KcuMP3QQm44797AqlKU/7
VXxN+kE8tW67yd5y6maPYJpvzggliRK84Xf3v1wdEPImHtExDSRy03RHI3UXZAj8YuxJC9udgS28
+woMQmHm1WlJaiZQk5TGq4ahnWl7N7jneDKH93XChAETJBpu13Q2f/c9ODMfO+kUXYcjHhLiZHWF
HClL5InuG3E6BuSKgJLNkndTEzNTxEWcKJzMOBi8Zdv25gbjtYaj0N4nlaxLl8Os/tgLJsQgdC4N
hu4SxW1d/vheA47AVDRwmaxsd9wmc8XY1q9yxVqlwV+NJkW9haVCL5byx3GN/pEK32LxacLdqJrR
jNj7h1XcMRMEMwYKpN1okmD67ZTrtZyiORTswpDs5cO8Uzof9D8bbSbMUOVgz5lpumJt7wFjJnfu
FPW4171QbhnVwidRFialUFIMvM6781BaNtue2jdyWADoBBhI7rfLmNHJtKnWkVUIL6vDl8ki8EgW
KfO3whax5Y/wXmC2f8MDQaCUVPo5p8pg3oi08owfHMJv6aAb9OgC7//F3rbDehBFKakQrX8GE1eG
C/aA/HAF08e4elG1rzQ8ptw9VYTHOOJVKmbOTEoFhl+7qWzexlGmMVtl2YAhHjNM+gN6HM/Hfl42
KLZn8kkSglTnD56qRZe6d7vqPxYdJ9ENBmBwKl8dPmNibioFB2l5/Ms7oT+tT9yp1Kz8ENH5z40J
PvWhEXF+0ZJ7s7Wcwujn2gRk/c9eeoHgEYUhosXLOHWWSNNRSdsHm0gIACGGnF1xgs44Gkn/LHW4
quuHKGlyVIGtj1DkTIQMybMBCgLYUMyGGo0/c0m0ywEa02rKkZJvexAS9fYx2IZ4E1jHeTqv7pww
lR3HGfLeBcXuLWjpc2QTQLVGyvM5i4fon20iqQs5694awp9ounbvKFAokuJRn/mW9OmmZndnwjbb
vp896ouh7AdXpQPe+4J1bG8pStxgjJ4mAOnHxBYoULAEOYx8bHVjI+Rou2gzW4OB4KSug5MCir4R
2ZixMNLHbF2vLQPbu80ORw5Hbdjtvi+qqMSb8f0jCpKq8Qh1shV8A3nQkiQqB3sq5hBZJ2pPYa4+
YgJToBdOGmU8VCPskTXw80MkKojKW6r2WpUV/70GsRzlLm5se+mzyt295CSldfAmlM6JW2S0290L
5juGTtvYnBOuuZraVdytD3j56a87+i9AUUHaHraSPwZ7hBXK79FSRP1I6YLlhI+ijAX/ay6FoF0k
/cWf6U85xYh3YHBwWpw0ldsAl8sOdEjsCCeOldfqRu9xyqvP32RJAawyaNhc5ksMp/B/z8ImFman
qJvPM30m0p/hKNqfs/LPHF7lfl9L9ZgDtfIAsy+KbYME3UVyJzw2LXv9ikTmn4UJP8mVLz9xbwvj
e1rKTwO0iOdkfPCS+3Pz4KASn10cdk1I6YJYVDOZW+LeqRJ4u5YzEAfo7u4PgyOt9aKsCl0oQPYv
NfbiLw1mFPhwlSWvJMRupMfnmuirgCJpKHjdix04HPaqPg2RumncNKDM66GYg1UEahHnQRJ0z00/
ARA78mrbTMFC2qx238RHNIw1oKdGEr59u6ptHoppiCxYbgDBe5iX8uLVq/zWeJxtg+0KcO4+uo+9
yALqXIofGNHKTV6NFP6CLZh9bc9YVi6p0pDTlqscS0xdthryoDkHtklKWZh2j782W9zhSAgAVDzz
3Aex94q0VHKsPLPkWGS3GC3WgXOOkGAg794OFuAQnaIfFwi9vR2YDcEON3J9bNls+8dHCEZbSDHw
Lgztfmln1NADcQdlhvlDp/Ka8hdNqHF20eN+dsypLF19AMqfrE6M2GXX/r8Pyz3fSAreAGA+gwGc
W7gZW28gGH8SU+h/L+puPCsVxmRE/++yo6b/AZxxND/md6zCBhuXOVl4hXmMjG0f/h9XiR/Y79Jv
2A5zLfAcKa2S3lozgC2P4aUNbFjHMBNhdIqgb4nMWd0pRvuMTe6FvHNzlMC8wPO4HHFDJDsHIFb4
C0TkX/lj0RcV4MPxUTnpY/KmbVhSahSgRUGQ7LQw4ML9a0GT1UsZvKXgS8JmO/QJx03q8ZY7VQ7r
00saKz5+nCGpOJ9eit0VpUn/6hfWRAMM+eYsvG3/SpB565ydyxEeux6S42DBgaEUkY6L2mKHH9PF
WVGCF7lXvyA47TlKcrWf8tvTRAP/zCDfLvW1Iik3S+cj1A1RMM6qrCEjcSIWYPk5tCjVURDKqm0R
PhW1/5iPUG6+qJGW9oaLpAI8HZE0glNeRG145Yoikj/CYNswwCsD0w4NoQQyWUr58VTMX5PMUhkp
91PUjcbH0as0CEOPWTPBC7mbwNEpId+7VxqzNuN5jmckoEzxz60CPVwnk6Wo3FME2Of1FyUYS2td
sFxEFF5If3CeWx+jDP+mdzlud0kuUwYEKkcDlG3znDtVCg7tlprTHPNYJzFKCqoTgcUz/hp3qquu
EMHLKeJxN1h4HZy0I0NpZID8O2TczQbV41i8JoIQEHDvyM5l+alnbpSMUZL2mz+xeqJXcNot5UcB
87MJqmp8sGUKqoz5obx+xgPweCubFpawnmKAFAjSEjs53m8QJetDUR9B3Q6YNJ46I9fAGdtsVybw
vGdJaiMnhEEJjf5WoIWuk+S2Oko+0cKrZvFvYagqHAy4nc0tw4KH5OyEFRtS9fVJRPQ2mN3yjM5O
JcmHy2kB1iNegpdDsXvH1kWvnqKiA6+BHY68M6OBgIjfFVMTRfQIophK4A62UvcZVAT/Hbr0Q7Z5
0zdPWnjRhdc5zOQwcbp7vfsScUZyabeAmNV2TfwVVuPxzUlP4KGkCmXNneUNRfansxkvyWR09+hp
+GIc701k60XneHePN1EW+7ZK1OxbP1VFDdBTMFnKtdQK7HCut63ZN38QMYOEjmIUDUIwKVbjPePv
omlLP+mALxyOo2iqvYb10S16lVM6RNvKLdKQmwMdU/i7XNggDGjWAyFb0dbtrZ2SOGBvGctLG+Ke
IjV0DOB8YxbHC27yDvEvai66wN3yGRo2/ncIzgPRM/IwuCLVU3sz1Xkk6etRU1VlbO6hyP+7J8Iy
7IO+pXf7irgmb0rTfSosxVVquYEVoW4HEEcW3ZeDNLCJF98u3HDt3uxgMJyeY8wnVFSsFCu2YRKX
lZurmdZDAiZNjwE6r/8JpJj3R8QOQHe0nTI+GlbW7X7Zqh46dQHnhHTwGJs3Lz2K25Us44eTvvEO
lb/paPQn54tVfefs9CH4161UpwBbx7berq/QdlKfGY4PYs/bYiM/tRMB584tRQD39+r2frlu7wkb
dzaYouR7MH+joeRtcv+nsnHpoLm5Z9on9SEE0+/NSOXGX6lZ/dI6Yrr/bDMOrJOV7Rn9Luumx8tG
iAISSk+iXqg9uul7kF6KIzn/8PY2PI4MAefXftlRi+2b/gg6JUlu2/oFtVFqXCj+rphp8nAzHJZB
1Jn3wZm7RL37ktisID1+gdsyBvobfV1X2mjm+7YTqtoQkIDpbdt/jmjmEi6KPKKeGvMW0sDDdqrf
XX1bvDWyKffQdviZ8nbm0EXY9N1XnpdMbhPHk1ad21EvRCZcDIAddGFUOjj26rSsJUuCHHONnyuL
p+Q8bmSJxiSIGEHSGgCCuSKNS5cAEJT2WkwGfEelQbvSGkAvHhjprRqpDWLIzmonJB9WKnCmGk96
fqhSoOMpa2g6o3FUInhgKhf/UwizzfF1vHeur+wEzdlmDAo5hugj1tutnHur6bC3p9O702KCnH0C
h3nnhVxTtsZrupNMhLkjUkPrsRU6flirQpuOXou9wth5L0I6uVERSPRyTKC90JIq7ivAELbtwbOl
d+2r+oHNu6Y6WIv9UTXqjB3ohrI3AK83JtxeLUteZ8JUye8CyJrzBvIikNStSAIVKtmm693tdHZP
lhtj7X629OnIE4/64JLPtKHwcQnNUlJMGE1jfitVP8qRleJWab1tcSfU7kd9okTR2wX3fxZ0GZ4H
wz6GnO7xTaekA6Jx8x3JZoPbj/MYqxf/qlu3tIW3cE1EK3iZf0lXFvNSFEWavawH4ZfvKKbVJjML
Rw2OUD2QhSoS85cF6KZ1ou8sKiRsHRrxmLd26d+g9LqM6ruuD+ARNYLE+3qog9WQ/Gc/sqkpyS8z
qr42FOsqxLmIWUQhn9nKCrD59DAByq6jW0O4dKnkzYrgqluyZBAMY9VuLrAYZY9Lgu/3MWUL3U3d
erhNk5WlZ+q8Ssl/gE3xRgDyO+H/n/UdFkzIYJAPM5ySnuiQ0mNiOg9S/uciybnmqCMciDCLUtNo
+wTwGWdLdxBcV7yztdbtPeWYrZSqD6/dCQn7xtJbDwvBbHLaghrMVoLVHujNmjdNjYLhDiB/meaY
I2MG/tO6s9s8KV3bn5zlTxbVpZkf0lMtmPrR6ni/V01hMOXMaKLJSTfv8g5GjFecP72jqdq6u4wj
WRHRlSNDUbRQE5GIXipCUfPT50QN8PbETiGPZROqHaTxDjzlDCGtbgpvWQKAyE7lZyt9b1dJzt55
L+BoFYzRULV4TQU2EyM6/gwS0hYuQAVIBl46teA1WpueDC3Sgl4bHd9qu6jBqjvOifyk3R0uy3OK
q+KvFqo/ZU/HnQgXqQEjohSLUo+rai/293QdNI5HypYxRjJApsRzRKNgzNznu3+xTHV0V6o89c0P
71mOlcDPH2pYPizm3LKfooM/Cv/G03AajZMnmx4fl4+Fm0bi+xjaxdKJLl5vfnxaznJtdD8EYd/h
JyfVszJRcjE9O9PMLCpiAhjftY6fK9Thsvbdw8WU/JJWVt5Btf0570Ehl6n6KyN2LLUsfCwcczRS
8uJUk7g0wq/IsBMq/6sDIeQOe61Mmug5GJNAodszVxxe/njUew3J2nomazQMBcXpXxybMX/7Pfhh
80QiUHfHW7t7cFDeh6MYX4xDIEoMEOZeTSZ3VZ8quWEwpZD7cMWZHIwdQ7UR0Vq33UTIq0FcSXMk
aeEfZdJ8TXrON1pb9dSPqQPgiPWlm+v1PXChCVasmN84XNzDrLQkA353f5ilyf3rlakG0MQsXfob
20WJOsUn+ZGN8owStJfKKMNlkiB0Ch8tgZ7p/NTE9e/4oBEt3h+NOHglqfPbEr4mo9d3UcGizOo9
HFyQ51vtrpTAJOnjP22XCxukkA5bypnYrcBDGK36AxLwgn4KGAyXJQ3tkU/4JS+R6DkskNUTw1Hv
q35lfdnpMLAf5GiJ73AF++PIEEnLC/6LBGfuXOWFOBbjl2yflQw5bJhkGdMcnCbhiDRH5NU7/geR
wJJc+vRsCwCDF/yrROlgLoEsLxr29qwBUsK931aRG/0Ag/2hTK4Dq/ki8pZbOO5ME38tPcUQFwE+
RAM0xkaoQPMusipFym+o0zqdERi3yBQpfaWuZt4Fa0DYy+ZbELeUxH06E/kGjkibzXlYyk+GZdYx
JKTUT7A4WMxBPyYtmMZ26rxQMU+Qz4XlI+LOnsU6g9YpBbBAovwyeLiaZjoPqjKDvgX6hDXUAa+4
5GbUPQ244l99lcCa9DtWWlhg+X8InzRMRtmZkJN1hYtiT/HVwMk6Mpsn7jDx05HUogBc/XzPszjx
aBSNiXwtjjMvV+XGGPJ4/f0D9L/8khOoBqTDEMx0cxiuR71NUsEOW4lkVaup7uZadba4RAaWvKXF
uKZ9wapR1Rzkw846pOgZrYpQLV7N4bEI08+TnRgQrLNw14TCGPyX3HT/lr4flrF0IoeP0+ppzS7O
Iet4nty+ja6pMP+E2t7MKEdTh9izbKcmbz0SuRwbVHKxos6+AnBNX0vsWjrRdP1fXPxeWylI8K4Z
zxpBJPtK8zhDhXEz4V4j0GRjmczNGiVDIU2T/sY80JToxGsVdQDlJespporE+ODugwcPsh18F0py
QYoXoL8KFsRzlUHBzCmzRpcCAlTqD6RdZRrFizE0ITmRBADgAP5loA2R3aoWXa9AbDS9ogBQ400n
QHJm42Y9AuVs1ePxgATxutcCYuFZUmJa/Q0ICl646IL6K8dV1YqMT7xfPwYAM/+++PgwRNTTr48Q
tdmKolz4LIsJlS1380gJBSSrTtfrJUeRXSG9Zi8MKGhHxayea4qjSInNvky1MJ18WXvOBkU0Dw4M
WlQrzxy4fkeipdO5PO3tIViwkiWxIkApKqNDttQsfluLslGtk6J4liP1qT5ywwBqmL+GnMeHTcBR
CUOM5U+LfKqAyg1SWTQ1Bwh9d6Y03PHeyN2qO4jA5nuiWrI/evUldzW2IzWgxixQdJht6ouwsRvR
fdQVd9KmQHb/h1LF3wcBiAj0jvD7B7QrMeuiVuxDF6XO/wBsL+8BKF1JJ0oeVEFdgbQrs66ZdKVl
p64WX6TRmUtywUnxlJqxbhPuogLak2djQ1zdKFESjJI2lU/+ph0dP9l4NTJ+XyFkgVqbsFJ4HUOm
tI8H0k4YGEAV+eWMiX7dIVq4Lc4WIlRx90XXWUtIltjXXSrTXm58noCgoLQ5lAxKrFpeJqyHEdao
sdGr1KGl4pPcC0F86ECf6HxsfNqHMzyiBNWikbEl7eQgKQ+n175Ej6q79At1Ujc8V3DFcE8lQbRW
iO8vquRUj062YZz7CAwhlAknzgDoqWEYz9WuzxZBCa6Y2f2tWgakzK5O/I7E39dON8vfAQv2Hw2F
b8Gl89sZyJHaNNg64ETYDwu3FhNOmDPMyNTP/nFyQOedAEahiNoFvpYPwdXezr883WBf0Bcp96HE
pE8F9X33i6MB+7d1/2GFXz3X4lIBaSb426xcNXdOfsfdOlJ3AftbF8FCh63JEOTyaYDYG07yp8hx
lbHdpVKpdy1Sn1hoUtt3T3Y1Hjp2DUIJfYiGSfzvp0ivFJASZvpEs6OPJBtj4mXnFV0ERUQVUrQF
rhvtckCAtkaSyoFVD41KSdq8IC4I7NxTUAqnX6LasZ6Gq2tulgo8t5M1yYKT4LergOAsl1iyxOYS
8VhihEeiosgMfUBI+SeQyX5bGhSl5z5z/Ooi221jEwibL+6C4UC1QPIgstV7JndkCc+RWlkKIMB1
gtQhmpcuC4LBC8Y4my3zyoAFsNuBthoAolGtEdq1X+9jAcIXYx3dfLvrAtJhrMyICZND7CxJVyBQ
mEWkuqGcaT96j37TztgRUT904vaiFikQB4eAKS6M/zmsaRjcHredFcx8pNWTixtWnXldC2g1sGv6
Nwtu1hnXoGAeLU6A3fUjfdzgL4XkKI4ZTGK3LTojgydTrLSEslziDgl1qQdO+KlR/r3uE58Gsct7
3WR0neMgUd0+NTwNf5MVldMpGkGxLiRhwNC1ZgZw0IX7QiYn+kci2ncVv48Rv7Bvsa0L5tQ4n2p5
/kr1IWS2HJcr0/SfKrfTP7I9C0wpg+LlH1Ytetjsy8xeJUYyqh16QNZpXJmvWIleqzVzYMAoWDgO
g0vOWzwpUZnA4ySAGizfmDbbFtzU+w3Sc8acJLqfS509b+QwVuWCPqPcQUKVlcTKt3ag7wCogG4z
hJ0JM42TZ/8QjGU5cVnWArYjdIH+6CQX9Chtce1EnGBS2JVFztb/m7knvUG9RtxvrotUzURKRffN
39dmpnzOGIUSUtFFzcLu/Cpk7Z82k1+CFCkR3uLAmfOqLYz803XVAsPW2ieBsWOhcxdYtccnrSMe
gk9r15bXixFw3WfRkn9/abEUkcwVjPEq6eacPPWG3Fg3qK55i7N9EzX/C/ao60TLPtkqGXY/qeQY
XjbnVu7TPGR3Ro9dWGtSm5BQ5Th9l2sn08APBu/sUeHwdyGSQE3A8ajjq/VuZ+SIBlxmuxc51Bf/
OMqjv1y5IM4rBtRA2+hF2aiP4UOmoopWc/sWyHTld5M0NJ8vU5ypWx3ixqW6NL2hdZzpq57TXns2
G/AWYI4cLQbPiQo+Jd05NeH/IR4wWZphfdaki2e19M/eHN1v+Eft7U0FFBNcikYmOtYfTrxmHZsz
C1AiQV6SNWozHOvIERmYw4Rgqv0QSNPn/W8L6OLBTxa+lVGFt3HBVWGbvOr0Gc8Wx8N1DHXgJP94
6iI6W/3KS+UqVP3FJDFm5VLa8wEnQ3Ll1LNwZW1VkDIY59enj8rWQ0YsPVRhJe3dq7iy/U9ycZS+
7yGSjzkGnwIwrlIIt/Alt+TW5/3T8VntoIc5hpCVG7Wrfi9kU56s98JsnUU0zSqCuqBj7U9NCxlC
x+qx/JN0W2z9uwsmPwwUUDOvQ1GhxVV2CnznAvqMaLWAW5c1LBgpPLuFqtz8RJIWy4HSdnXXXY1a
lcpZirOY4i42qdQKxHnEAU8DusMn/lqk5ZcpXeSbIwQKL3e9dEwqKd0rjW1JVK1RgsUkHLd5KCWp
ev/0iP8L6elnCLVvZx/DzzBpaLpt/yuK+qsEmRQ13CNsMrgR32SYycGOgBgzbAQONNHkWuXauEk0
KgBzYMfP/G4BuvyDViBAFTdSyzBwH1WjhOwfYHfPx+shfhvIGSykzfhQnG+30uP22bgloQ/0EvL4
I6g6teyf+jAo4CisNIisQThAjFGNO8W8vO/JzVlLtyJr76k5uoMfnw8tH5HUqlnNcqYKxo/xz2cS
mz/Si0uiBWhFBHtbODsR+mYL/IKbijohyduq7uRTreFOkoUVlD6MuRIIE3LKSPnhiKjCelOFddeM
SbKgDkN0ldwWL6s/XbqaawBMx/pU+nZLhtPgNTl7FaVPR0TFPn16A9mRW7ravstN+viLimsoING7
Lpc7H7PDBdFFu/xo9KcQEL79VQ6dog2ulYduQg2c3hK6oR2RrULJ0wURomnfx7I2LrfDWAz4scCy
Z3C3PZ54+ev9tzRByltMkeqs4/WbKrgcDD335IIO/6QpfoXLVsGXXauLBjw6HhtM9k3uMYa+3QD9
CRrptKeXhLL1Q+NBzhLcwuqmnF2VrbNmIJ6TfVJjcl3+jfrjtl+SD1JreyIH/NDl0fkKA3CJuM2O
oVKGomrlRPElqHBS+y9VMLeYm4y9hEZKiUuqppuWJ+szhMOlns/ofu71LwFsbH6hMp8aHm3waDKU
kcijscTD9k3DNcDdqzdcR9rxTYhzUU6nxjjCW2ADqbpJw15G7tcacKpsEnKQlTblMd9AopBQBzqR
Gb5tcrv3gePDHxFpeGx8JRxbMmpk8R2EdE+fDds5xGOV61LTqQgz4GEaeBLthcEil2J9mfskbzKE
rray2GC0m25rsDjH6l8CzP8KOATvr+ihgb0qZPOyJ1SbuJQkIXJtXt3QnOrdf+KGIKyAiPe6ERkm
8Z+3D55qklgAkvjB+Ous2pa2Yue+ZQt/MbSLxkACs9T293B7KbHbFD2ytmrE/TNRUSPtSRNZDdBd
7G5olQcvrpKNKaamkmHw4aqld3/h0LXMIXnGxFhB0pQoWjuKz6T1tIXisWDwS/H1zYI0/YH+jy0x
bcEcPcI7YDDSanIlmVn/5gyk/ZCVmuA0+LCb9lXUihkRIx8g3+dUN3aTp5PfePafwVOCn85cwijA
QUPTxCk4sd3Oo/xjH3QRASCB8vsa4IFU1XNVdKEyGhDxE+/lXt4ZTAERczWpay9BjbeChOVPZNQ3
S0FZnfiKXO25hDuz9IbPx9o6xkjCcOSlAJOnFcCf1kDZOId4cgYJBnscqYYYLMk6kmI5812JGsKq
d67Tqg3X9DlecPIsGIcfCItde+LBsl5JRjFVMoONGBQ3X672Q706ohy5JQcwfZMl7G/FRVoBh5hG
zepzUQN6E1Kf1lw906qCVEBiQdKBoCAAOXlCCTciOiQdg/5DiGEVC2anoQjAgUiuO3v4cPQ29p8Y
JfqTmtgxWhG+Wxwbh/icGGnn/YLgxcHVbgdcgwZTGr4qyTGsC9OWNo7EuYpn6n9pHQC1PCIfUeQl
J5RnZUmt6zaId6jOUZ1+XoaT0rJxpgp5ZHe3jhr2dzD3mI2m8+gHN9TtwmCpI2eWWT8K1hj57dct
3iIMKoJuF1KOalA2wB0a6oT6ZPiHX9UNLEaP3eDJUYoQhY0+zPZtpvHVI4CZFaxskGQeQDdjCJCM
lgHPrpWK9vqTDnF7AIQIl/qwFzOMJEHwtwRGLkabLPC1ujD9m9QRLVWVHfeufif90AbW1FuBVssg
R3Cx1j11+HcPhc/PXgqE5Fgq/OPy0aE9p1VT9Lunt+6Yc5RxdIjGR5ZBrCVGpHxMv1Y3/Ryp7w41
KUWRDlJneYtQjIdEkKzFt0q2yHDDFjACaLSAYgXL+CGZmgDBt6hHPzhWIbpDDJyho58+/CpgMnPc
19JlEsGp1c5rgfZ0EofL+4XOdxgozMjLOG7jd2tUyEaT+vInRc9NbJFyl4OrkT2JVif5d5Ms1T32
HokCaaZy3Z3UIONblw/eWT7VuSsFifSIJiXybJk49CIV8nOQbMWYk/4JwBfawaLjCk6rF+DW+GPJ
RLfc57bgj6BnAe56uyUe9ZeXGbi7mUKX15XArCPRJGmel/NdcBKpYrhtmBz+LJzRvSt9YeCvlP2y
bjxnbZv2ZPC78csPLEPCrf3dWcRvYogfkqNoIrha5T37WPC5/WwI6TOLAuVPWq1onopTtgPR79zS
QEqEvYiyRYwnaggHwmKNFfI8vb0/2Nlsok6lR9xc7tic4CurFv2niMs+wO4pLWJOZ6+WayFg9uA3
rzPhi3ZkRCpv7X9HUXslRaJQR2W0IxAMwrYudPb8P7xqKgLdSEShP66b1Szu5+wOpwL5XqgD9t3g
gc5y+my+xJBKs4Ijy9hhA8+Ua2qX3/jpkvUlW0e1WFca/0zn6Uu8Jl/xMAS+FTBg0w/yy+Q/U7DH
lzhTf1YwZKjeAlyxk6fjI4Fvy2j5/FJCrmlSFf13GwHWlLVEme4fN4SMxJ7rb+nMPtSJf37JHU7c
zlO7UmTRjkHpENEkY+V/MdaSzixkqG4okyNy8CxPFNQzD0g0Uf00lRlENeCzo/NeZn8AKcFHupK7
hCO9CiiKDck1cKr13T3CXDsLNTig/TqI+ZHv0zZ7417lKw4GCuMuplNQOcrRLKsGvq7qgMHw8nr9
RwoBBl61UUF6hnjuEi3AGv982u45OqNmtfE+rx+nJ8ufNs7lfkEAURiRgt+p3JjdqQg5DS+N9ZJ/
2V9R+MBcnsOL/zzQCRlKR88S+HNdaGOr/BJ5IaJBGcB+ohZpdmTUdrC8u5azlLnqJMu9Qm2mS/qG
Cr2G6ImNVdC30FywLUqRGsojGFpxifZ+jrWnhPwIKc8nbZQ2q+Lbq8ZWZAgtAsIglfWi8Npy3HYP
4TWtrS4ohJ9wdPE+P9cokHSO3H7CDP8LBNygcDmeKf4p/h+s74/+K6HubkiIfTxBxnbJFAd7bztY
HsoanZcbbt1VH+1US7jcCBrWpaB4+I6aGhpZyQv5x7W8CQEr0p5CJA93gNIG5dzVe0P40NQvhSTh
WnBJRAoEwBVhvlJwxO4nLwWsPsk8czExoCQYT1z7iP3cC0UBwlvOZNyPhQu1BA8VaC+mZ7AHMoC4
6eabVG2ePhbeTeNfbjZI0nRImXv7SIbcvn4A7Uh+Q7IiTa3M2k48QwTW0/FmZ8Hki3t7hIskG9QZ
4rgJK293Uvel3VdiOfsG7rfJo9ZzdPLI+FKTh9XiytOxgVVia+dauymQ8xvYWUiJDp1xo/K4dmQb
975B5IpZdjdAh/02yI5hQuMaG2M1uLZxECBj3EQ0bkW9ZzUzufuOluI9xqG6PyShs/UaB5RSvk3r
blDSN5SvHDoIzXvXvX/mdUSy1LNUNJ8sMajKfj+dzIEZO7ca7+NRDfaw+bfTvFZNjNHyyeA6kZpz
T5+SwDKLgmpcWuVcVAljGtcvESlYjKPO+hgzyLA4Kl5Fck+29kWM74KOUUCulvaXgMBtWzi2AYEI
zyMvRp4vnTSWxvpXk6V80k/nPN854lj5a9leGA0VW0uKsuTfAkVKpWx/YrHH2/0HGn/Z7t1yepsR
DHo5weaGaGhL2ONFfkZFC1dn2Asyw38mmZmZtWTE3rchq8V3HkO+6DbIqwZFaLvMDuWsK4ikU0IU
DQ+514YAz383nlY4p+1o2laMMq9sZH8GHtgapIFumlY+M4HI9g7L8stDwXrhf7jfJ8HGu5JCPMQ0
w3+xF/yzacdb/T31W5HWNZ22y/8BLBFqNW7EhaX63g9d2Dt+c+P922lI/LClH5uoDnRruxi7HeBQ
wWwwGw+Eh0pQ8Si0dgE8QkaqDeE6AGyPlL+IIaYArA5BXtOLh763u0Gk8ueDb4Xer3qYokFazk8L
pAtU2DF570dMO6VBO9UN5bi6VonjhYiExwq/ZyD8DmbY8qu24jJIVet39QMwrKWsyLW54ZNuNRj/
SreFdMCwQWoFKTaDvKnGmRz37QLb+6IMwaadDCqmNWq6VizmpZbIw561Ykvd/Zjxn/lloPJlH3l1
64HUtuJSsuLUfIaygRdnS+2je+AtUIEqh4TsMcktZNdY0lvNTFSv8G0aJ8e8FqNz8CgynAAny63M
J84/xTBGBeOx0D0ka6CS0N2A+gQuX/WixfosrHhYvLP/7c4LZB5PTcPxahFHueGDKx89ecbgV6+U
94SK8czfuzWys9QBYCUmOZWAAlC4Rmo4RAJhlsrXBT8b+WGn+QpM01X537jwU8Bdj/uuXEUEwNEo
klZkhGd2KVYlaT48BwNRBCQN0qEp92GLSopuENBRLSj0JeKF0eac+g/Az0wA9F/MCXs7CcDojolc
bfTu+khyT3jeSu/VwsawJ9iyH27RJZFTPzw7Sx9tAlUItbMviObposMIUl3nCGv3DggMeM9RNmOf
OtM1f23SxJ9wRAOwQ2F30ULgAIQIAtdOkWJnER0H6ADZWEiKwKZv0VLFr+2wN7yB8uKk7rsnVe1C
5jVO8P6RY1j06QNxG4Lvh0ujkPXuXzpD1ynGThEZ4i24TQ4nFGbvbr9K0wOoWO0FfcPY+JdL2QTV
2znl7CLfbyxhiyStnLaZIaxiCDDXTYWSXWUNdj4xv3dPhlKB+RyB180hn7K29DKnrouXVngnPkqD
YvaE3iBFJdQMNW/Dt39BmcZcyoKz7tHG0TI+4hg1DAO8PsG3OgvKzjX4Nhpexs1bOXVXfP+89LE+
yTguaUxbFTcA/W41+npTT9YiMGUzM3QrY+6h+zH+08AuBIP6gW3Jh6T9M/uTrdlipPgrcgCkxfus
puLDQXY7Vxd5ZPAnZ8WaFDOm0FHjmKk7DtxdrazXbCs0AxrQyNFqmEc85gejWZNygl68hbCSYwv1
K4Ez7NNJLitdOzWlPhkLj1wWdCZhv2myCL+GM4ZRZ/H+jKdPGjh2hSm6W8r4r7FLTU9VJXYPXpgZ
cyzSQMsTx4uiebSCt6dj5yowaAnD78vFuDz30wuZj0TbUyQn5FZOtCqmCKKnicCNtfZdnJhXkELh
EIxH10IFKKuCGy65B3rtNebzxZbImHHop9bZdWOeCkEP05Kpc+MxYVj5ygAk9/JExwpC8MrK25//
ON3gmq6vBJvSHM7TIon8YG77uJyV6c2nfkpKk1jLQ3wf6J0vUxO1lziW3FyPhJzBIQAPqChqwLqq
N/K/VKriXd0QUb/k8hAj+HXtpgut461kzcuAgqqIdLX9Bgk+2jJsnuVL3oSLG+3/eYs29XkVAouI
EBFtS0PrJ12hizKMFBhZND8ngvhJ4qazxpkktmIJkwfRXc0z72WX5m9CN1uV/0T7WowovGxP71b3
hnRHzdIYe0CJuTMQ632PZdWHhby1cgye3pImuJdRHD/C4XJyt9GnX9L87b+xzwhNL8oJ2QvRPlyv
7InKbiHfrWWyfSDAZgIbW48UTgaYr8b5E6HxQVpKnT0jhEpCbNbXUK9jWSvcCDsUhmrSdKuxntTW
I0H8b7/bWK7F++RlznldsEV17OBOF1luwmZfwbW7MDIzmQ16ex5jtEOvLe5Tl9lvsvQqf4qEaP+d
rAuTTWWOMurYBdtvqcDJmF5eRMpkdJMtzoa8U8Sh1C70OS8B2tea6JYD2dCs1kTbdcSa/ZOUH99U
Qgllm4+RVNcBK4CoiGdYZOF0goj13eEsDwON1q+eHU5YAue76m8h8Tcjhy+iksArOkhDYFP3H9xW
qbbHCjvBkjQnKoth/6bUbuWmMuC3fKA1lZA36smXwldvhOWif0D4qlBArYTnR8TMDgoqnqpm4aXP
TUHGTiowYzbQfgngjVEEC5yJ3uz7Qd/AvF8EoPu9KbhcrGTsPBAdokScuzwba+vUnHgFpTEoVFKY
JLmPVuj1EQjUU7wfvJa7u7OrJtXvD8tBt0U1XofTr6ZWcwssPsKU5HmmEM+xMBQQqtDCK5SwhrDU
yRLD+Msj6zrrMrKXusulxBoBOFLmRcs7zaElMlxUArmlJXKoX+o6k/VEg9S0i/2lpb9lDV3Z4dfb
N1+vjGNcyak2xXfbAvxwAaBjuZ3Enxc46z8XNeg5NdVT8v1LmwMTIyz3aurXqxaxvzbyoPf9FqHQ
YxOMqEQA5TSbLZWuwsGyMgTF9pyD1avTVcUeey70WoHBBzxNH7/HqO2whkf+EMsubf0W8o1Kexk7
KClgICZQAkh+iEJxAvVu4lDIGY2y33+jMlwuYf49M/f62ZCo6X5Ptam8iyWwbYGAqbRJZ9w0wTm+
Cdj72yrnotAXk6pqlPblnocS0tH/84IOZpEE8AwCV382qS4aQ4a+hkPk3dbnL3h6+avj0usPkUdz
8tYwrRHp/28qw7hGZIb55gnOnE76KOmuFHod+3toIGTeM15401VxGdNGvAtSpY37yK+FMJXr9mDj
0WDNH3RYEAmhhU3XownKNuie6QF0wOY26id+/UnggOD2KZ9/zdeWW1CNFSU3NuWnomkD/Es5j0oy
bkyekgSFAOsVsDmElK6Y5Cz4OsRls+To0I6X9VamReHLTgO8dmN6ZGUQLddpusmS2og21MB+DJiw
olhAiInz/AUhRhCuOfj3wwF+E5+bFxmP4o7EzuNpEPKdpwJnOKfzNNROmEzikMZrAE/egMwZCfrD
aFtseZfV/l80tvZOPpk4mF36Gt4XQuLMjbx8w8STOSzhkjy15Ka1VFAw3eN7IpVzAij4WY9OPVxq
29eJG0YVQbh5SsHft3ez2YAJVnDVrS4/R3czcYOkC9NQkCxSzqN/qvqjexjqNjTr5DeM0gK5czKj
qIujbP6BOKJsRcNHm0OE/HYjy4PmbbChXPR8DWj8wqCeMQUhdoh8ViO7IUJ4QArKbUpfr/txBOjg
lxaBAK5ZZJ/TOFEvbQEb/w0frntNonEXfNzCy47iSByzrloBeSFlyvKI4gf5ox906HzhXNXHR+L/
ART1AoAtsxaxUutOss9UFuscYCfzwpSIgvljBe0ZYyBorXZVlRWTWEFmPvWSa98Hq/QN31Gp4IuA
2FR85rFqkOaTOuEfBRp8EIAkCAmNM7jNKSzpy5b7zNyP8eb4oTKWgfcrCKNeIhpEvUNOnx5pt5Sv
Z2NpQuXe39ePl1pviqOWZfEVupgu0LAC3aPfXeQ8JiqDzxUlN/LJs2D+bUsX/1JEnkWvK0x9SpCk
6lAXwB0eC3Pyxpgx6bQbGkSzgILeUh20jQhtmBksXd+Yv5zhh/ZDzdRGvrDJs14HhQaUoebpPHNo
Q9oUu7/O/VuN/Isa7szU+vBIdgNk6zQyE9ZP8yelcxSEaEYK9LjQnHOrwAisxeZJUiwBAQnWy2xi
pt7YQcJNfMkjlAFSPGPBWmnjtkxdKXZMUcWl2QiqujSDKyhReJ2cv1WR21BeAN4HfBYFctwjkCak
pAYHdOeK5D3uTsVN2H/0vJa6Rb+lRRoVhJ4q11ze/l46LzfiK92BDfSexfetMeP+zOKT2zJC0QIL
kvyOcV/Ljl2wdungFKlxKsSD/L8Woz/aQrQP6yAEgznylOBiHmbDAOpM0dZU0DIVbWNpImKOmpWi
t10Iy4x30TLOUp3yXJEG5UM6mB0Vznj8JGSlmJwuI76ZQuslQIpnuE1/XpSw/u0TIyO169S6k3Jn
2u+mn5Szk8CjvXkprpHN1h3ioyyDtTytyX3/6LP4r2gc1SUjMcuLHnt3+yJlFRAmni7t1sQam2FB
HYXYxJkI0Qf1KEMhmfN4w+rNFbrVyOkRWH1j1/XJAH45mPeUo9iJTZ8+i41LKgYDvOitTm4L858J
qeJ4ghG7686tf8XDGzdTCBl1PucBkAzqc6Mg71HVnvqBbqn559fyE31ASy23fHw6vFfa+P5E7vUX
xGvhUjbTou7lyh4owmyfItBYXPdPghN0o8ssICgwc3lxMWpsqknILexyWrufFssaqrGvVDBkONYr
PmDYFDpN0yQY2+nNYf9u0FxIUlKiMWjGFZwN6+QMX9ITIqVbboRcOeQ/TDU7p9EJhbqHTYoVep/3
Tu24Phsge012uPk1iVDJGaA/BLw+cUh5TE5r/ZI5uDMSiaKBmZpIYU+Zmv1imszfJMcTt1VYoSNB
LHZPIzPOou58VqT9b2wfQ/K3zMYAENMeqGObVopfRaflaQSZGB5UqsJy3818zV+zyRhvSSYsnwtM
bGVZNMqytnrw90VlK+RoCyc2ixA2cHnpCv5PqcJsL+UQnPy3LIqHcvAjY2zk+bHDgESPFbDKDzeP
sS96ofUnHjrfY3HlPXvD4vq8u6YodBn6yDfj+Q572/SGM1anOe90CaMQy59wQRvNyH17N18O27tf
WmbMwQkG+p1Q7ZWnn7pOx+KAwwN7vz2CK97y3WNiOoH592VEC2LxtEm9qsXV+5zRgSCOhaKibXKO
bmlEiWDbXuJ1uI0hmX0sTLecG3gCZceaiu6Bpq1aVxJNHycaBT8zOyg2ODpOwag+9or+nWABC0JI
1ADdRMLGlpR2oqU5mHW71EJxvpqur3AyBTBzJ84BvixLvhKnsoLL78F9gPxfIPRS9yeLVBRE4HxV
r02DL5v2DWrjxtpMtnDx4FNxINODAZwF1YCTNs/l+3NLyujntkgZO4aguGmM3gxoOT8dTQF7uOwv
AhaG8nfoAQ25AT24GWwD90tRUN/zo18a+9vBNr/pJGN2SX41StojuWs45AKZcGL0A2Q3AAEvE/Zx
7Ty+bu4wEaa9fD4oiSbv+gmOJzWMYAkL732LfUJV1QUT+dNCco6dM9onhCGuozS+zrpwmaEZyB54
6/8Dzft6HPHSCaMIZZelkW6WYWZ2hZpMPMWDpvI4qYjZTquGjPT+hl28JOqM0rBxL2LdAsTxXQNk
th3/dGCE5/gRt7bGQYNOVQPRj/jxcwStrCdyQOvmR5LI0cyFhabWBQoAzYpfwHy9QWo4Iyk6Nbsk
KMpsTANDuLebMBelB2bhW1gEoVvU9j0pn9qxvh14v1t04qkuOkv7nqxk/2ZFDEw/lKiZRlV/Cli9
poNT0SHEtTh+NCm6FMwnTEQqYwye8oreAyMe2rbnq5bBfYaNJnBx5DOcmwmf1sJd6OAMPApU3M7s
TNIwni7vkwBzLbL0xAc8nUpxUbkpTxQH4mXWfLz98/HuZWzg4RGUHNMmn9Avorz6edVmrLM2UDmw
aczJ4oXSHd5nMnsJkZIb6iEX5njuFj2NCOXra9XnRHTmTzXbDz8befUn36uZihRfn0rEA9b0TQmq
gqEUJzpjEFih51zSBbZSnNClf7PVq/fyVyMx3WWWVa4L15MgPELg0Rq15Kx+EXhPOWIQ97pt/m8h
Ib4rpXmCjQCe8Zfaoj2ugWfgpspUVDGWt9CRisWgzB7X8dHs6dAEre5CN7JDTecNjglOiFYHY3nO
D7v1FqhyVHweDh3xhOYl+/10XyM0Hfw96bj25WeE8UQzmJBPTJvtNrnLJgYM7lg3OClZqnfnRpNo
eAYLocEZYGNqIJzi4SjRTC6EKzTnUSQTKZN2+hdUGbl7rNFqUsqwWUw/2W57uQPCXF6ZrV3nz5Ay
XN3Sf3T3lQKBfdxwEZXQRFqNmpjdLf36BgpAnJiwU3r3hywUCfDQg3G6lIhUBy23R7PPSBGV++Pa
7Z/d6N4I8smhR/20pO+9P2Dy2I3r+S16HRhUZesJmpNwvrxx8W7tfSrjmcQm6fpLxyaH9d+s6lxK
kA4VB/2FLh8nTgY+L1XZXxbfNmSqkrYuutY7mrpUvZOJYltBffLpdIFm8g1JG/ykNeBh/YrAZqMs
joPd25wMjVDH2pRAM1ExQ/TUY+W4EtyWeoAXGSGW+Q4mFrih9Tgt13mtgrbH6+FMbqCpikBqsxLj
HtZo8f8Sn7uSnEw8GC39ujiIn+/HTeLBFNJ3PDG42JDvC/aMoeQ7bF4/cBoIftHR6mni3IGV5fgj
Iq6KzzGpPJZ6jY1LNTdijIBRh9TXXc922nhAhhWvy+81MHXpfYFPc9KxmSQUG3GP6hxSGjHO22qy
/LbTbFtbQdPGk57YQ1zSrYkr99LILLS5NZpgV4NSozft8u1D/3sqRU/PNecrn36rzo8wTUWV0Ci5
CJLq9LbvFEB+jXk172E6D5uh20Jswhzf+3JwcLra7+7JMxcqSKTHlr/6NPR95hUOvLsX7bN6cWUr
MtoN9fYiwNZUp47p8RKuOqn2WFErGCh4TXtTUVCzl6dSV/RjBwGdDkJ1tsd1zDSZ4j8TcKe0qTR9
Vj3MLhWIIEzjBaK3GGDlKLgXHtGM5fQYXOwFGuZ6kCr1Fo6mNgjafxZehHM5P27FTS9GA1ZsB7tm
JXxgZ7eWGn2UwoKne3v64kwwAlRC6DjukDJxBkGAqmWqHgTYujAi+AabljUULAMuAr38f+OPg5x0
DvKx9xiES4zV1LKnS8bX/MiE5xXPM8Z/Mk1CfceORGH0iCLNdKAgNYSd5tEqpzMM+xIzrft0r73c
7fOtrVR/h96lqFiCp6vnzOFo6WI9xW7Y3H9QYRt3SjYGPmUL0hNn6L1ODyPpRl/QL2Om/zqf7v2t
ZRnHXrwko2ucV8UFjxBXBE2NrjdqvZeoarvWLKBZP9zfKzXkI7CmSnbygA8JzytoA5yLSe24IhfI
GsXDZveJou3eaSlhgT94q/+UJuTSfkcafamSIJkD3JnyDIaMwNGzmUvmOEDvAcZQ2sdaz6QZ6DZD
lWL9DgTR36MMm01Wo+IVSqCLi0AlInTdUQhfGsmbdVkYppRUPG34sMm4LKXLmidc/9jJ/nY7C63A
p3AWx10JkdxKnIw0UVciTcqhmyjc4yDVHIb6BxK0iSa/59cjFHqQipeLDw/h293cUrqyb00dVDrt
fRb5TI8AVSlOnAIKDJt6/1f7ftKX0rvhJncs+e7TtL+kUmO7nVwHc798xlbISna9A/D9ikGkdjwW
4dZ3PSvyjvdZk0ZFBUY1KuFbfskQYkWd10LowxEN/QXq6PqmrJEMuRdULVxy0Q3jZaQ/B1+oknsX
xImZ/4rtCKCaqWnhZAjiB5ZPbe0EWGxcfWBC+NDw3QLPDD84dNzBRjL0RXxlYNhdl+CDWVRH7cHa
iS6xHkFOy8utmsz2TDUdwntTzwhUDTGQDiXYo7Wi4znsb544INE9kbqS2t+0KWZTTHllXm57dV0T
1FqA/WmgA5dSugaefP7VIoJqqLcR6T0lWkEqi5Af9RVA+gJZaao1WO1gFZ8Hi2Vuz4MGqjDgxNAw
43fjCqdVvbfA85xdIFSpM/NBjsHCN+f7V+W8e7Ugyz88nA8pNoqYwo0AghyZXaOle5dSCcOxqZ4A
22ab7jkLl4jS22EHgm1aWWasOQ8YyxUa/F+E8tPLOtb+wHR/mbTx9DSpMtIkmGbwnB+dLtx+A4FV
ZZTOqTmZSPzwkei+AVXaH89aalvocKx3Rum0PEt1q5SivD1tKRQ8fwVRLDNWrdPC/McgfSl7FmCz
CctH0IfVWaM5uaa1n5/uuJVAxJU328ujOYAxFzEFRcamQg9BRykoJVh2R8buX0nQV38HzcDuuHWM
ji/Y5dmp99+PzXcGO2hwin851UDj4zrLjSrsfFBeEIDxSJf+MzX29hseYgFMvsNIAMznwJUcJf5t
ZfCvlOu5mIfgQBfss9cFfhms+hAVi7LepFMkfL2hAYBCsxm5/FZfMfaocmoxdmVfrPMGIMNswKAX
d2ToFaqNl+CPIvbvC+0hIrNx+Thb3dmj125fXLZ+jBeppX/HrDAzQfHTdtf+vI8DOgHdHKV9Irz0
RSs9ARrqg7JkPhSOoHPCmy97G3Rn0i8i/tHlvPRdu+Wri0QFySotr6opJe43FoOwECXihoFfjKB5
tPNCF6pJckoXAlPeupHzEV/v0DsgUeHLHQkiQ8iRZOjw1tyqZi2RREt/pksSz06zirY3CAhfsx8K
P1ITj8ty1tTuyqy1fba2zyiR7EYNcRq/+7frxJZjf1dDs3a6vOBuF+TaSD810zzc+GTLM5u0UOP2
ZP+CNRbZCLoh2AjrmzYRq4v5rcolP9FHCrSWb9+yspMtsm7gWQu545HoWJD+P3Js9r7LBV1yJC0q
Bp7RaJEIZUaPnuV5FQ7DZHMCzFmwlIKrmcoqWO3R+AexEw/rNqwlOcuK0Xn2V9HfGNR9ctQ6DVn4
7AZ0LAiw7cPLIa8EF6w6eLvTV6ZvHz6DV+n2aNEClEcYc2z9uUKwkaFCc29T6EH/nsD7gakbgUuf
MO+Fz0TDDVoBxkCWSM8j1nShqpXCmh2sBUVBB5mBtHXyiKJAFmVPyOEeelZmNajX5YohgvgJEwph
/TKvpMhjO2pEDVfq2MZubQ/MQ1Z6aGVwCE+2FB0VFDFmpTsaDhgpmJ5Q3edqaJcTSFFk7lbPEjzh
0LR8VizqIo7IlmXfr3MpLtC9KAKq44d9H0garI8p5kSRsI7bGajYGxua86WB++SwsnOK/ke592TL
ardz0nC37f5siqLsSTWpBK+HPGtpqaptrEFLLbYO2gsEJ5bhLRAqqSsPbq+mprs2JGjdokQ+7twr
eLg5j+STYJPbH86bLdJBnKDOSmqPI8ap9QZk8o51dW8f+kC2gRK5AZA9yueRF381rsfNv+qrLynL
wu5F8fXuSaTIT/k7OKG/jdyC24cKIIh4YPv9pfKqOAelKFa1oyz72esIAMon29IONvBkzkWDzxqv
naO3kw1p+hQehXYAbImsrhrnwlxQOGRWA0UHs5AU6EDZ1i39ta86lbtDKWJLNkEgxYzhh1pK3fNv
nkFwcAABmWY1JkjHmVgi8KImtKb3iZbOYvGSE33/nKR1egtBTW7rAZu5a3XpM1kYPZXbe7iVAQsW
cLwjeb0Wk23jt0RhkzvxGTqrBY0KdxtJKPjDQed7rastrcbN5TeGfF+H5CC/JAEChiJjb2i7OEA7
3+N3gxaX9moX/52caaT/rOQazIQqQil+OUjoZhgYsREQ6jHqc4oF9O22ZuP1gHaLH92uDYpu1Iiy
MfqbNMJL2gjkxyVYIMDBFWP/UDdct4IM/I6anmT+ekWnVaNaelP+HcmjGJDBEHvYifQ4KibfanTj
chBSfhxHDt9kNo+Lm5CkBkewtHdQW6t/eZQRyhZJwKziAufLxeE8VuzQRsSV7qwo/iDdkBeuKjbq
zt99157R7V/UfZqTDSxs80qW4rwsjaWkI3RxMw1boWeHewEndFjicLpnKISimd8ZpcPsdq6XfC4x
sFGjI0GtIZa5TE08s1IumZXDUdDs7s9uvP8UrO3PnImQavOaUUr+k535k4croUm3DyR3STuL4mAz
ngysxAFHv9f3cB7ycDYNfOgquwl05ZyXGyQBVz6vz+M9JsN35Pq68x0kL3O/g8Dwk97KDOVhuZkq
IQCE9G97I8jUvVaSZ2qcQThDuWBwpRr+F5b89DxNKOyte0/9NXXqNzuEzExgp03Av6gUWWt/DYhy
nFgpZ0/pvCDLj2L3TATN8CxAJ03Z5xtykBkRPbOBjj5Q87f2HGJ+WdzdPVhC0r74fnCa7pmh12t6
lUdC4L0FpKC5KVDJplwZe6aX25jy+79uz2K8+Mbb2oUvWojuWgJaX7dhIh9jBowJlU0e2Xt9kOL5
S44ZgJZHU8fkNuTwRLczQonpDkHQ/kNvl8XSXa4j/eMpjTJrO9Dy5H4eEyS2qyHfWNwNwg0JFn9g
/LiYCTVOhPkHNdBw5/p1A9HaoM8yaMF4CH7zgoyxzpR5ZnVKvDdh+lNCqKdBFYgSGhM2OuLz0m/V
D3BFXbWAmQodc/YgO/LN1A6k+v33aW4eRL1sYOjlZ/wEFxQ5rxziuZC8eHq3fyZx17HYZh+wLyPM
XzynlAZrZMVH/ev4Wyimt7fZG0c2hDYKQugvYB0mEgTzZ5uEZ8VRWjnvTICHMoMYmU/fJjWD4k8x
S4GbfeZzkSKmrd7SPIWPLYumCJGyol2BhJm0YSKJmw2eiJBmBf8ZkZmMMqUGfesUQc22LaeVi5ZL
eOzAKj8z2o27guhqNnTwXkO4kMZSdSm5rcwZ51or8t7FJAi8xjAUMS5l7BWvMmKJD4UOHitWJn4b
+aKrdIh6lbYscNe6EbxX3DHw97EElQ4KvUMBOePOWCnhIKYSoSmyBisNiGtsYqVyWdCSST+w1rRp
2b9YD7o3M8kzEBywNnVA/VDjGKNSrFez8v8MCzwJtOpm2WSxy94z9ilNtp5JP78FvPBpWVmTpHpG
XPEFcVwJufOZDcRtD4Nm7VrrLDnYH/tN2e7uhRni0QpExT4SRt//fjSs40Rz8i4fMEQ5ZUQEbA2z
PSLYLpHWBIsHFacUCQrVVclpmb2Ve711U6gDjJXKiQ0LgZsRosJarrX5vpmt/H++ElYQskp9F9/C
KdWU8X95qYjoic12qbu6gaLcF9NbU9svwR7Ri6qu5dLoMOBz16JfeMZJbk0IulGIlvgCRBEFVSFa
Vp1hMmTtbqh9Tjn28ru/ufGYMJQ4xZ4Qp4ySy93itEyvU1CQq/vjnQi3yzQwy2uPbkB7WCVWkana
mntcJdhn7DKEyDVbxm4PZNt0blQSQDbkNnYsJIEOwCLDEVHG0sOIH3vLhNqvSb5toZXr2tcC9VJP
aezgVp3+DiDrbkcf2HFM4+AR6fHdantkpM5utBZpkGZw506EUZ/QmBhpwNpX6lYcQI91MV/ocBe1
9wND0qlOILMnjAZx51e/rOdNxUm9DYoQPac6pVnnNLn8rJsl+xOLOlyQfCXQ0+7Ou8glKI/0JzQi
8ctPYDq0D6j1LZ+HDpZfFf087VlD0HbTSByzrnXGfHW/8s4DdWLvxs8o3EDTWPGq1zgUZYbYKBfb
ecA1O9jEnx9/XHtZc0EMjIh4lUKd4GFb9GPd56GHosOooeUrHtb+2DR4HLViR/zsZdve/eN+tc8S
3cBdYQu/yIny+S7e1cxB71zZn/420tmJO9QrNgfVZRcRng/ZL7tOwoUcQwvyWxKvDgUq6hbRSlQb
uMlQ5eHa4UACeZ3YKeMSHS2WIM0mgKgNwKQb+P0K0tb8hJiGvT7Z9aytJYcc2K+/EU3psa4Twy9C
aAUBEFJWpaHw9WwCFjntqR0IUbaYYhm/pZWqgnO7m/mRE+SBU8m31siSVivA1SkmrRd0dWKEvnvJ
puJwLH60IpplAyi+CoUmJCeMCCa0QIiPexZxao9Gel0+VMUQmEsl+aQgj2+gdzTAitp/bxcbdJ8F
TrHUV1b97clu4CarO50FDWmzZ9o43YWSMmJFsLn8gYQdeMgQXY0DpC0vFHSA2iHP1j4l8wBZ4InS
9uueEMJOdxGjjMZ2WFbn8sybKN3koIvUwSnEUAhoAf90pjdxQ1WobZIGRyju3yPGdz/tkHTHEEFv
1d45Fdxxxf0YqLL2kWBnoq818B4p307rvUXDCKQCcdebq1gzYE3F5xz3exZ3y3peonYiMaJva9Pi
Ua86/VCOylsBDckezkAu6KKMGm7qAyboyUWHkY5PvoGub83Sew+KZ6PDiniMnlBuFLG1cBpNnrnG
uv11evuv5Eo+yMn11Exz8/o6+x2quzopSKzhdydUq9h9TeZhNuHsB8IHPewQ6LE/1qYzohR3cgw0
6Ssuca79vmR1Tp11lQE0WLpi4ppOFncv2gt3HCrYWFlsv+/xKWRUAEMG5g5TrOKmJrvyFU8dYCUb
SLuKs6GW/VgrYlxhBgtbGmR3L2yvc+BeNFaw5+z1jNEZuZZYMsaGLsGKI4Ul4Ud9ZaSss//Mi8WP
WLpbRkDf1bx2mOCXqBbWfrQ+5vrONxK6vJbtntcwLvXY5irrjcynrFVA2tGFG+Jgr/DWhwdFH9kv
4PsFLWdZ5XQR2mhmvqwxkDe04zNcXFlvVMU7egs5rUlmjfNftRgUEayStXJShXlYr4Ns71GR0p4b
Xo2BTzFJTe6s1qiJZ/2z/LRW51/CWNxPPs+lpsrB9U0Mz0A5ra/wW5kHV/sJCTm6ukewa/qUUYzG
7yWHJTzh7mmiTGSRteIdHBOnIeTk3lJKHI1E7h+wU97lfg/Aru5QZVJX0/ULWtlJh1Ys3LTTxeTt
raRzfCDXDu+RsL4p/0TWyj0AUNS9KMo+laxYrguYGvvubaPtXMy4ht36iUph+81lcG3qQQRH8ruY
B5JHIqBatfyTIeFyr9cG4eS7/RAKm8omtMpLiNSG8+vMuixkZLaorGDaOYq6CFvP/dyEJYA5LmK6
CQFYcw3wuMgJaIUGctgHRYLlbZMMLvNHvjgPLUnFAXVocABvKkZBKTRlHegTKdJowUlcKM9Rqp5v
bmz/87E68bWkhZ1XKh4ceYOvC3LEzmw/xVx6hpGsFlISsfNbAMtRD6/KjevoX+GOxC1yBV2OxplN
mqLRgJen1cfPImklLWIOfXWOYofRPmOkbQfWBC6pzmOehdvO8ObYjDK4wNi00Qd3CiiFVIxk3LNg
fP9ZpyX2wSiNeEWRhQa6zoC2Fw2PE3glVnxKCvOX52/KIrDlsyL2BAQE8OiMyuMXD+qEP2CgFbVg
w5T6p+8Wn2GpCPbqj1yy9Iagy1XHnpxgkI8LDat2Kxho0bMgP5XniDd3OEhBFLyHmGy9o5vO1I5M
eTh4Z6Ortc9rmPq2YUcbYTh1aXm+tqFf9IWP7w+t8XMbJhc5N0+e/KJCKH92uUWhvxxZV0iZMPaB
YIm+WmmYs282nABgOk1eKmaI0aj1pavFVkHHW2X5gcykiAv0Ct4WELzOZJiLqeZzKbWlOnVtok/D
KAytHnlEYcByhqaWOSDNrZXl2EV4xds7u4yyBnr+8BgYa0nYMMmSUJ5ge0dYGwaMV6Dq7Uhuqins
fUib2hAZZArIEyULFSgyGQ/QfsQwhu897Pay15oc6fCtVRlinbQ59EvqmOxzSoCNRq+BnMVKHlQo
bl3C0zHHmEpeXSjWLcMlXQ8PMLqEdsCqeMPMCyWGqN2kbj5GY697xRYdW//KCR1AE4YlvBKpCVDB
ZjNPN1iwzNyuHP6Fy8F9e20o0uktemn2hnmX+12F8nbcVZ1/3siJss67qyIVXFoPFsJGTNRN2Eon
4c5tuxw6LBIyMGtHLBDv+cLL1A1LgdJYT5j0obLn4mFsStuOzSIm6Lt/2VShuaLbjKFvnUMnCZPV
8GCSlmYQSiobkjXvmv5OLWtL1BQ68J/ODL4zFnu7PJ6OKzLgFVCcY5X/JgERNBwZzrVTGUWptIZ7
bknYwlk6d5lbuyKnIvlHK6XUiY5HZMhSU+6ZzW7y6932iTkQR1MdC3IcKB9JuZMkef+4gIzMFaz1
2x3urjaayE2DPrHDjrcdb5IBrRUhdrLHbQe2fX6Sfp9lA93xyXwNjeY3QJ5MlJXaUJDGNUoPzOfm
t+YIXQ44RiSlNDQYH8geIxQSEBrN4Rp7kYLm/nI1SyCiyChkgdlmZFEJ17jff6H3aDzl5uwMR+95
D1T2F++ziqrt1hyJEblHY5Xk+FJZWYZvh8eVVEiRRAz5DTvA4gsvrbez6e4N3vj8sf8bp+ue3aW+
/FbmvJuj0wZ7/J6obQ0LBNf6dJOX4wwNLJKgKNEhCUfCa0S42TkqJFPlaMUp6yVGNwFVBwOtuwOZ
Mlqp0zqBEM3H5JGEQA0GIkNb7280/gFu0wgIbYCA3XWHOyWRmJWHPVFq/T2gQFxm9uH38omFXqff
08mv3Huc8KgnuJnvUL6hG3IXdqA/MaHYCctOzx5TVsVw0md4bs5n3oP+uVNL8bSRZrHAfXM2MIG4
Jf8PjVCdO0LO80JEu1rd6E0V3KPDbNHcooucTn014kYk9Ko2n6TnoshEwQYi14p5dgPipW7zrJJu
8f2mL7b6vWK+y46lUr6TCgL5Srcq82a9BP9LJXcEIzI7SiBhr/wyvollKhF1G2EaDV4MirqQGk8b
meU95SITHYPi0zcvoqsA53RRwZV6oasOJseyhZ8Cwyv6Vg1YcXhU5AKpw+i4htt9bK/1LX5FEuwP
m8CVG9OTa0zyi9anPMGqmC7Az0zvK+foQyKXH8jbJ7Iu44rpJBlwvQwiI19G75o+5kCKGKhEo5ei
kuzthRopHRIvsnAKwi3aXWLawCWaBfGdqX6B9Ws5V1MRWRZkHCxAw3ZKf1SR0ausYoKCDH9IO76K
wiWJOk7EYZs+yjWf/0VY/FjpYjkvI+Nvj80Z1uoQ1b2gPEFpBy/BrYI/Fx/fVUM3Hvde0sqD3FR+
JQOgZgPT4MW8+8p/swonYJ0AcjR/PsIpGOstuzZI9iU1N6i8mh2xteEKrhMc+hIf0SPD5KWRNhoO
onyhL6F6ZpU+jlLCYT+8NVSafL8QtNAA6OxCa1R3DgCnve/oCWTr5jDYpoUw2YgDUYY/LsXCoIt6
dlBW9kdJ1UxVecUoe+Juyy8XYtWB8mU1vUr/CvQ00Yuv6+hMhx+RMF83KibPZlqG4meYY6KDLgUP
uKuOJlePC5Cso9URHM8E+DGtxMPahmob2JI55c1fAHfz3TGmhvovi+FPjyMCkGovnBS0XcKx7mI+
1FYVFOwPzBOKXKHslKSxlSddFWJAWowBiiNkdCsxWOz24kkxjoHtkJDfnz/JsfVUuvoH350wqek2
aXzYWQGam1Q8hZ7nmnDLU5C1zggCAbmvCC5iqpqsBVjszOfXphHlBdJpNZYFC0DufI5cUh/xWk9x
G9pTFHSSTm/vWY/QnTUZfz+Coay0QbIljZf2N2TirnW6JFYzKGlC0Y9MaKrkGuAR0E6j45TreLA0
/QwgB98YDTtUrCRpJuYXRogocsqODlDb7mBBAz09UmS90qALX4DCF3Kb0T3HRWnrg4ARBPCwsHMQ
Sp96RQInJ5nGyAI9E6BZDsZ12wJlGqbcmKeSCmmHYJy5ZMq+e+kw4g7rpIoRdneJU1Kk9e1LXIvh
8x0GJBk9SQ+pLI1rPyegqlpxmjDlxv1RAfDFXD/YJetWd+O9wGe6ZgmisZeoAFPF1iQYLDONU9BB
QC+u7YHdClXrNTZHFyYUiuMrgshflgxAWHkhz0pFMrghZjd/qvFqfWs/kKkfZOyzx89GuC/4Ftk6
8wdu2C41d9YWKfE+hJG8r/wRWECAnNxItmFH3ctolhmq4IPz9p5K8KtLwg7+K0Nlf2Hf7VG2JI8A
f4zAlgNMgxVntQ/CAVl93dO5wyq0004jJ2Tsp7hvLcjylZgdGErFciA8hsReiDFCmeK5Sp2ogb2w
E9OvkwZ1fVh5Ulzn7hlyblMgdJMLVkuzP//e90cLTczoV5Rhte2hxGxQfxLTFVrAQF3hqOEesBD1
JEa79DUwBCaOvMPs7215bNfnQJ507U/tsldXRRTshtbgS3eIaxOlYhFHIF+2rbuRcm4lM84Qqaow
kNC2jPUzNd9LF1H8MbB8V3xVFFfyL7lDcUbKlTOGIa727H6XWrzWebU3dfrd3aQ7oczX2lCV51pD
kLC6b0wdywILTqpLwK4fLNqpxbDkGbabKWbXAjRIbTn8Xu1c9GlACA1K3SanKvDA3IO2L5VVih0F
awtR3dtxs/W7f7DccQwXqxIwvf6kZnuaEwQMxiyQI7y8+T3owjm/fvjAcWHx2P0ZBDs8ylQAn9gN
nJmXhlzOEsv8n7KBixll0OZNGJdcsl+aU0XibUR9d/zAeMC1XWz5V/LZZxNQh7+Oq3WQ3sAUG/SA
RY/+LLQjb7NsgeEm7cNrYBsdJuV74QLbx9sn3ouIPUW/Up6K6jBK2MxXjREuXDAQ5KrrPgE71Zc0
ghGX1NNy08own+A+v3h1CC92DK3eIxfFSqxAcFmXmmqx5/EXchC9cjSVN/xW029rGs2YK6deDZs1
g0sFGs6Hp6F6+Otxzb2Q/kMIItBDfu3stfDpjiDYlUtixZ4G8FAmCg+0rLyNsHRv+kM1JWDw5vSF
XFxPdpHdiJjsbjI5OfuK9vD5WA0dzbjegR04qSYrzNNPsgnsMJ8k7/ABLsLpiJS74f8FxZDf2+0p
2Ok0tIu18QR5pv64bLbcOuL815XD7z2QW7vWTFeDQtriMUJJfhTxTlNavIiFntpvjVi+Zxk2pwW/
Az5lE3Jlsogk6+35YhYzETUqfxX23v3R6HR5IDExqdfDob2OAUrWVvj9IOpyjWww3HWMvEzbpSp/
nKjO+kzKGmMuUfkWNUFIYZBCIFGyvaGCiEL43kOwqVVtX8gwzpbfZjw6ReTyLVxeFzK7OrzvZqFa
wBij98bpFPny4G4jBwDr1gU/l9j3XYKiroUClBHzryynmaTI/SKBAcPaRAciETRJbqgC8mPr8AhV
NV1igBJQhNodF0gkUMbq1vWPzlp7XzPkW819g8b600u++Ox341IAS7GVbEDsKg//gpujkAktED3P
e2e8fBhsg0umcvC6u/P12lOHh+soPznEZl3bRD+nr+WQnGKMjeQCZ4XSlpwSRf/TsiQ+rE/rBJga
bPaqWczL+72t9e6XVy0VpqghNSjaeKPZ+FZxJ+pWZqYiHzY85VxkPezawVv2eLS/EOYd9MO/P3zY
pSLaDQuvaXhpjeAZ8Kx6aRX4hKrFW8iVHVKCAkFq9ttHGxU+pvDXdLTTdb8HcX0TdqSWdRU5/Fpq
elN6H3X58Z1MnUBVzH5nKhY8UU668Y/S+t8/CuMRHdH09bbFu/3bZMaMkzTx9iNW36tN/byqJU2f
KI6jhi38DVMXdCM8YiPJo10MuQgUISteJJ1Go1XevyvLO2Qdx5ocN1bdewdf4XZDeV/9G4sX/peQ
FLcRcPzRTvIAM+ebhJ6oFOpbw4s8C767l244rEkW2+q29feJud9YfB47AyhOV9ngsnMAY3uiKu1D
T0scaNRRuTtn64QHBsHQzkyTvTXMIT5p972gknGKIFldQI8wpyojXgGeLWmZ49KG21IQfxbGaE9P
ng9ZqNZdxTpdqV9be4eGSh8BRLGq+xyoU4J4gNve7m8MB7XWMFUzAo3Ehn86gGkjQKtBFpejrZA3
g72dYv35W3uxLj97sA2oILgQ38RJzPob47nxtmbJpeAWRfmsii5N6ZimAJlX286Jixaex8qgk76G
jK0Mdi6PHDCQNUCUOr7cOfx1YckG5SGeaslu3/BamzovPYM2QqzdibBjxBkp1PUxQBcKXskmutNq
D/hwIccsCnqY3rho1VhHHYrQFbg1FJqozFHVo70E6zRTJuh9xMyVNT7sa9/eVXdsxWTyXJqlAOFU
GnNc2qQn4uBtUig5JBegGBxiPqUYtAb8eie5/BoyNvzFQ9j8Sfb3Nh/PnPAvnf2GYwTOx1eEmeqz
O3dMJlgZcOYItDUDKVu6Xn2AgjP6OkUaWaWIBwWOQS7TnevgRVBwajtAP04SdOXQaNV09UUuItHI
8HJD5w7m/FfrEBIJWByVbaV81eoMTYt4u6x8FgRcPIiJV3HM5ccvqnAjB8qDge9C+azHQJJzotYy
7w+pgLhhjWDskaC6DXKgbIshnxytv37G7i7kiNsQaAcyGvW+Twm8U9f0WlRF7gShyUq7JOhuG7mk
/OaLTxyd3pZXO5Mjt6JiT7ztB3wntaovx2B90vdph6y1A8mu1prb9gETEZxOfgb4PTi/XrbOicfk
U+dP0/MyGznnBcqwUieEscHSduxOVy90GQ8VLocSIb0I+/pNCHhxcJG5fmqyKnM2wGR0YXoI/UzN
164kgPQOkwYGTi6RuIeHSg2KTnDmWOUVfLMoy+aDx9VUcznHXzXCFjmk5NhCSJ1YwVf+eqCn/cTZ
a13AktbAVIc5NN9YzQukfXCEBYUWq+r5R0JNwaagO7GCc3SugrjEncEMcEVQgR1lv8NZrHuNrNNj
LMyQRBK08r8lTrEC4lkLXFWaEXiabuYIdhqTua8Dpp4c+4TEiCEPzjDKLkfQEF8NG2cyIundi+/O
jiP2gyd+XRpszhi15kHUH3D9ZSrfWpkNDPaJXxJlV57FeVKrToCO2fpvdJRrrFvjA/i6csU1ask2
/3g8WgQ86UdY7otVhTnvfKdeXxz4klfLjeyLsG+g+zo3gfnkEUFcgQv6zeDvPPaBkpDfYa/ynVef
j1IcOnZBwxAOwjtgwshLRMoo2bRvatIrhRjzqNg9tvIJIWRQACHL04//Gt5azT9md+c/9IUQJUPv
sZ8UhGbRKTH5P1GzJCqQOepLFXobEp11YOqVVMj6+j5W7paeyExK4n8ZHkizP+4Ji7fMTNitYNRN
u5FMF5NBzve6zYLaN8IOU+2hNB7ztWZLEdN7FHkAmyPepIkg7Ora8bHg8IqDUZPEolnaGZGQ6tOJ
i68vh1cW3B+X9DZ9OnzIx7xeX01Z8jWEHKBp2flQULcIBC5HDTdfQWMUafSYkEGzpVswhnjOmvgd
TtO73F0e61hxWqzeiJS/lTq+kbzYsoQER+ysoIFCPWHdfXfDxAv4xsOhhuka0v4F2QsBF1Q+0Qa1
e4OWcLEbPtCIe/YC5q01WR8X4K0XeXrQdcXBgaqkaF7Ef7YjvnpX79rnQzq2j8JX2JXyiqQjWtye
ZTIQUg+fcSWizYZh61BAtgk/A437X9W2EuAMk/Ma65JFVQoBL6qk7rRp8GWAA5omMBkHRvjDQycO
xnYUYXFVduBYObXpG6UWD7e9b5fm37pmp2jWumOXAPVgtw7OYtwnMkMUvhCeEy+G2S5U/tMhnuUv
QPw9qCJa/YqYFDsR6yjJwph8q2YIgqTejLsnRAbcNl6//FZ6JxIZ9T+3U8W48Ph6xfY7UVasmkBW
4o2xMiPWkcFzYykq6tjovNWmFZL7XPboeUlVETm7VbnAAmDeJChIjb+5dA9vsQCR2HqpHEtepgJl
M1ZO3HSngItjSI2gMAzxZte2VFzNDQvXwnOs6be04iYckocc/fR/ZNOS8IaIgciWrWeLObuPYzQt
Blb0nY7k28cdFXR24AiLO8T9m5NmLjH9FTvQO9XBNc/cIO2uwQQPwXA6S6+cdhPMn4gQLOhPXtcF
Xb43iWXHy6qkApi326nEzN72GmlXYZEAyQR0SV3+NHgVxgRq4vAGrS8t97t3aXTLS8DkAltlciWe
Eru01AyTryGGWq0lFd2oX+Lgd5fjV+lErOfV8ouFkbeRSWStN/mVKts2OegheLXI1kwGtElY9SPJ
J+TqiFk34qseCdDwVEcsQjIbJMCX9928CvfYqevZ6CQyVBhN7HKD0UaERSi0Rf5sbMlGBBsRxxsZ
fKVHOvMB93jzLMypZBoZYgcdLZeyaz1CfkwIQYgnODBmffNK3/QaEgBTosnxO797+sNSFMpTaGFO
Wrn+wBtJ3LBoMl5E7znjCCM0p+LgIuFu4tr5kGHY3OYcfihdnRaUsfW+2b2gVCrvFdzuTIhBRIX9
6lDLa6Ije549XXPUe7uwAuzoFRxoyFM9YPyjzXKZ6fV7r0LGySsrOBoOrKvRnUEv5zyChypbGGMd
801t73MG42NJY6hH6JVJx2i1v3Uz+AyGhcCzBjhvipQGHrLjF4u4nN6vQh1kqBZ+QrBE0O0BzZGm
CEbi+Ref3xIumUw1yWsd1ZZXVfeNOsIFw0ao5Wyc6LYQsBaWjrYkgqgTeyqepZW5trH4pmXH+I6Q
8C44YTQyMBjaea1HowxP18fcVHRMCX3c5tsCw27jrBQi/YAWQIdblAnsKUa3allMJXilro31XF5I
x79k8nCq1SCPpNKPfZKrehChcZ64u8lKfRGLy320vVzyA5gWXnf/LV8dqQDarJD5VCNav7tv35ys
Qb1g1JdmTwLTfJM8vHfifIrpqf5a3jBHVgXJ3XmM/UID3P22T8fLT/AHkYQtIUfJA+GmBZq4/14T
YwfwOFfnqnmLHFQGiu3iXzYGFFpw7CsVP0f8W4CAHjmpeHKirCyHT3wFb6kqwlVZcoUgBSd9HC/0
/BTwcxBpHjTYowjQPlvYY5s33GhdoKd/9bQD+jgmG+UMGqE6d24Qc2HtOkOWxCFL3dikhq8hYZRt
4Ui3BF3QRPKvgo8Klou6z/zrewUiH08i4HNY/5yg6oAHl9QQEAhcsGLye188yenpGdB0nzeAyKuk
NNch5IQ2tHyYSJ8ERymgc0pPeqmbu9Yce0jghcY00vcoosR+o/TrZJrazH0gdbB3PzF/H7imlD7j
Ky7q/EpJqyoqXzSxm2Fm17IFdjRAzwjybFFR6A8mkvrCW6nzZG0thbNf3fZXx13MZ20QrLnudOyM
GuQKGStEmK2j/YAEi8D6j4A1VJX7fL9LI4xC+SUMYwyOU97QvKojWTt/ZTqveBeGd8atCdqPxCPY
T6ip+gSoFLmOIrc3D5MfErMOwZbN0rrUumiKr2OZZi6isN/iVRq0pHW/HwAtnmaS91Ks3WQGxD/M
9Ks3S4AvbEMiGvFXD9OkcxrmULFQhEGhBYU9iUWboO8YtI3qZo6Qp/fS7PTD45r+hq1HDzHIiYv8
Nvrf0wfryZKO6mp357iQLiliTcqvIa5E26NuDuUX0Hpn3J35szsA2Vjgi/WSsAlMlZsrPf7HFfF3
Cei1vo2EBprwbD5oSK8uQB9+eLJg3bHrb9kFtY9fG3mmWvvu9vXmqhGyuLVL2heV5ydHThL23KAe
o/tIAhoTtX1GlILGtYJE2qBhNJFqrIOS1Ug+VNpNk1wdMJnc+Py9lqerMkiRrygLsD6JmdZ9Uzx9
jDxg52IdSRtRPlb0DjdJxPTFnw2VxNgZ5gbpBmsj55cWXZer+E0IGfTpKlfJ4HHff/3BDxvC08VI
RbL6JVDlBRjwfuuYj2/DbYrYe7J1uwk/eLaTtZ6pNneaMlEhfUz5z+uZAI49V3L9j26x77tsNXo+
AB1ha4nkbqwyTyo137qQoikBcj8IW3k60WYM8xc3RfWi/g0gfq7gOknkzNbVQuzorUtprDCSqUIt
oM01+Vsgg4Q+aKpZlShyetrQY1Lb9BitYX0Zwi4j/K0a6v/OCqUe4ipiQC6e28+PDmfWwqHD7jhc
rn24CVfN8iVECB57R9VvJesR+5aAaIufIUU1nbe6/IGBhn9GVlXCrLD2Z23qRlqKDODCHATBLlor
Z5WiSUbB9AsDfw8zkklUq7fhrG+bppn36kjoLsgSbvPjzgDc32MAuJ5jmqdM4zwI9UkMnJ7XO29Z
TGG+99x9ro0cBJYXUGOjrONJkvQVDMdmBjZ4newyyvvixDoK44rqoq6eZlH6ahKC23NxQWzyCB7c
X4NpKoN1DdeAvSkaRRFV7hYHj8uCLGPAVc1RszaDAGumzCn5Q84iX4TtDZ6ict+KKCMaW6895XCp
TInSgWtS5lyV+j0OirU9lMARPWfLkcqxcFPNtKSGcAA2IGgzXHi9ohVpRa/x1VB0ok8aabuXAYJ+
Awi/V5q/oeCFHEeBONBDBuUxy3t+Co7ktt6TH22rcPnNFJheRQObLVoWQh3DjdKhFhhXctZHcWW/
JdctwGbHLEyhvSx28P2sdhQLu8AiobBnkB9CjPdeKBHMCElSQYCyv5BGThTyteI8jlkm9Oxn2s3s
cmSG2HAIOtI9G1P6IwUK/QdMsiIIlX6JrnpDiHQu+LkzYnYul+Y63Ojplutb4nAeArd20ujssX8I
QJjZ1lOmWPX6iySZRTThaLHNLq1efZuf2X9J60wED6Rim3Dzk6E3Ve3JdHCV3G4tBZPixzLgg5MR
1OtQe7y2DzcRsqxFd2vps7Yuc6fltefC/sO10UEf2wS7fxobfXgPO3FrSmccOmk6taNga2/tjos+
9FT8A05j1RA8l4JC627//XYhOJf39f4FMj1N6xSdBDcVDvlLLj9Zxz2qH4g+mItw6cxpW2sv4j0M
pr5IhSQcA4BHl8OJxk0mXWpgmnPMcm417EnnuES9VPcaCVxv4zawfTPLfUyF0QmKFRcreoKZXD1M
iu++GeaMUap2zxB5PGTPdvJB8yfW1jBkZ0BbV/I5c/Z9RmY4XuhkW6Lv9H7USNxFroNNIs1B7bP9
ZbZCZN5u90zA9Dbmy0QUHbIziCsEWajw9xeY01r4flqcUT+FYbaF6Xpz0ouyaYpNB0I4KCSnWPpF
VrKrXtTIPLjLRRlj2K/naQlRY1RSN3rZBSzrDx9HO3NdCXSqLtElzseCSHgsjOAjoyy1Jjuc1/QW
m6spei84/Dcf1qjO05HWyxw9dcPlpgscaILWe9bPSZX7K3YmvZZV/mS+QgE9JHxPXtb7ppxM0m6y
2EiDC/a00lYRCL0eDFQDrcp94xT/kKFMRVn6uKbjoemqFp8GoePIu+HcVDqA+ASMI0LSWIMhTK41
Ir+TTGfeam68TficKptl53AuZSyqJdN263iHzrArVJFcypLmIEPumPeRVbeEsD+a6i5eLzl6frct
UtLUbxusDRRsRs3W9qBVq96K1Fmhqy4p1jnAwL9gUpeeCBaOIwQ9YVvv/2Dh/qL7A9cX5b7tsucb
4VUwAI/agt+SUVJ+u2ap4CzZsMtzYFUUBWPrvAwxwTZ7MwcOod28HQNbC24aX5mc/u8pRo6+Bi7e
j5P9rjD0RjM0nho185YF6BnkZjqfp4hAVq+h+TSHnZ9YWLEWez0KCpXUtxKykRQiuw5idQkk/f5s
KTQeqBTY77h+wWB72MoCeDhX5kxdlqpw1qT7q3YGfWd7QNQKYM6NLL9jUPLqwKLYvGMjSPgi9eI3
VQuP6kGJ+azKRS2+/lK46u4Fl0Qo/lwtnQAW1Lmw3bTaOI5FH3YzGVEXj/D4+862RXHGBHfwhYuX
nONHGuHFFTfMDjLR+XaNyCg/9RUnjUnaEcxngZ9+ONFtEl4BK/EGL1Xq6xV5Zf1rBZnRMSUaNdyP
CuskCz60X8zpGn3tRE+d6ekMXLBHS0A0wx0Baht4YE1/0oCqNX2g9sTZYZbqGqHPTJK0W/YsqPot
3zvZeXyynA7ia+NwqPaLftFIdReTxp+CITbckRZqmlB8OhgbpMZny63rJDs11FWTQL7GNHZ6YRIg
Bbwpdj/RQBwEnKN0KNx2KHyj8rIdL2n+i4BMfjP6B0LuZk8CPK0aiqG38CJ3a+G3+uOIytpYL+eP
uGRRaRgFo8HKa0DB2Ok+5PHCRpdWk9rYX3h3XV4S84fb4fcx2m5CZ55fwfeI1Q+vS5whVT3pLtl8
urrujY6hs0lgp/LPARHfDuPFSKoiZYeYJ7p1nkiedoqyr+oV6V7fzUQugRhigVmOy5xA/MTsMhjV
tVXD4iQifNceF1TIj+dqIFsWwDZ5nHctE0F3wHjXdYxWVp85LxAvf/2/9C1hsVEUMR5mn3h0/JS9
EUNq2ncE1uqSif9I/vyr3FqpSr1MeyLDxIgfwfx21dMa4dApQIYw+S1zYU8gJej4ifivKjpO5OS1
+S615O539qYZLBohUA4TApZh5OI9HW8DWbgHxJ/5YqmhXhdg0FcGrxkQdygUQX3luX7OaQLPO26+
2DS7ip64DRXFILdcJnjbCTcciNwLbh4VFRgWgBZu9CAws89c+eeSBbUFlkloF5PulrRRkY96nKM7
yfNGArslW60nIl14suu2+70xG6rst/Iy7moPhqF3SPOots6LN8jFHccPywFpz629o/uQGjepAWQD
jGp1CTMqUXWp176UBDFR264TghgaDJgiS5JE3stsN482NbO9cXzHsa6OLvfUZF7hOxxAlATjKokI
7V+vwaMoiV8bq5yVt129pmSnQYuqMKj/8FELdpDcOw5cYbouT3AT4lhE2ogZIOHaaK3zNbXQuk6k
p7O3PXFrAzL7fpPfzLY84EeNFx3w5byqF7SP5/xqCy4eEeTofVG21IFCT250gsVzuI79Zq81LK1S
+zd8/+0mz1EeRBUR/TNV6HM+CIOnjqFyQ8M4h2aztlcJU2tkzRS0qQjFwYVQLUwEFAgMSNIFuFtR
ROzCgjnrD5wgjmweP4s4++Zj191RZNIhIMafQGdzEaAc2j9SsKEfCl0+QEtKL2Tr5/UON/GUrODK
mMOWQdcxbXK4jp+2TPSHUsDeEC5TmVnj3m41IBlO146TCnrNtHIumjpwQJ+EWuWQtDCrBMFNnWwb
2NmX+JSaIEawieFftzSjA01X4NksOX+Nr6qOJ51Wp2x3yc5zwYgRjE7UczmGqZd5raLiOoL4HCIE
I5mxIgmX4yRyRRBHiIG00txaVrm5ImzRvE7z68XnfIXmr//g+kfBM6gDyXUIuWI7uTusHIi+/esZ
0Qzb+SlWkyQoiFYzJxV3ls3DMExpv1VpjYn55JS/2kCNNlNMXqM/tLp6/E24xHkFg4eF75azzP6R
aw0bab6JuRQDijPNxtH4HCdrk+SCInPLTItW0XDWZxPFw96H8v+7fDAZm/6+TtxzUhVl5wfBbcSB
AYRz8XVV56HkkGWX/gWrN7rqJFQ88A2SuNJijJfXnqzsuDYQP9gr9pLoOV7T2MqNaiIreJu2DLgG
rMt09erMFS/Vu9/zmSHSNRzPh4jXdMX36hvdDc0UzJlm8jalKKUvCTnp/CGYglFtYTublLzPNs+A
Nqd9lWXo2xVAbCs5Qy7TOBtj/MVVi0G6+McVQtzNqneSb7thMIeBP5y8PerNKAPrp6VG2eYaYfCQ
26BlubyZGmIzDIO08oZZQcEIpeh7ZvRjm/DQLyBAXGwdYGg4XjIr431hTeeeAyHDk7jrWbpsQdID
nYJyzhpUE2BhWM/1/kmbTgu22YpM16kF0LZlIZz53Q+Pz/2oMXyvh2Js282zJ1ZrR2DnaOTcoGlP
ARW8859K9dHNenlEjWAttUyteisGr7bSE4QPVRhJbtH10/xY7zhh8hMIoaKJLVXLzKLp7BUI/SAD
3wPU4+1Wap6lKonHIOBm+jOoPjdh/R/WPSFqPvpvQ218F/NLu7LjLLAdDFH041zC+XKWxzgO9g2F
AzjFymeQa1c2qA6viC9dxhrcTjUu1pQQd7AfW7zjvX/olayJFfEbXzu+rn5uKCp+N55V29JtevLs
oodPlO6IE4pfWXo1HdGGeSMxnUeC8ghoBKJz9A/qAjLlKUC4mLoSCuKfv2DOtdk2Q8tEUnTY2scL
ecXfrNjD+64h9c8Iy0QAy4oMq7uh020v+ybUCbM9ubVNKj7HWad+WKqrNM8yiu/vUTdGgxJJKXO7
QEwKJv6jv7KxykpQQY6eQmiifPT5/JRGDGZ+NQJxzccoIEHvgvuxsQf/+yZg5xlA5wOPRur+eArm
i1RVeTVnkdxTT4JEl/Viw57nAHkPls3J3TmamCjhaJ4Xo7cy2XSSBlg6C3iB1W3oDSn372v5/Hej
fY1DDJMZwg5l0Zomw2vD2fA/ZgNazpSK8DbjNsJFVuN8sWT/1ifwonf84kIUHTE8uBT2mOXR9q9s
RO3AAsVZKGwagpLxNw8v8rcJMEvj4io2v4GVfKOxHRYQJrIbUEQzbtE8whnGihWXHwszMAOxF4G0
v4MbCyVh3zYF5SCeujqTwd3L1u2QSGDH2AEJo0kXkk2thY+lWrXTEaWU5S984jbpofmhuBSihYUR
+PHNEgLJ8eoZavGNQJXGFejK6yd9P9lfSfPSBGiOa9SKNLJXSzevy8SSP1ApaCkNJpGftoYaXJ+z
Ul3ivwQ9iohgO75NRGesmscCU4Uddf/NRKfmGP19lAvlsu+IcghHRf+ezOTf1t45klFCFfuD+c6t
MuoNNFWDp8SB7IDlkHmhw1JjioM47UfVxz6+YUjE83kP1viCXVB3IXHgGG/SgBmR/6yryk6uOetd
0ZbR0GZgWXlVprabYcpNipAMtYeNDnp5xcY6WTfSxHFSBU6NVlKRYRCrhRAv78663JgZOxIDdXxM
3Zq1T5lYRkymd83V8TDP9fSuUgszffk+gGBBiC8+Ztq/wo0vU3CiId7JpWQrWKzuxOorexZLgKFL
oD4vEuPNP/+k1FKxD3813HWfjKnjnd1avf2In4MjYxEfALeeJZ59wqUBCYOP10+Kn2pXYRIOpyUC
S5cbovouNZgMV/auIh9I4mzSs4O3dtfguADs0D0dneockw3bbwyHOCDjVUgopOVIRCQEA6FdTzpN
I19Fb9buGSKeI6GIYTJ2ZpSXjPEYzSV1UYqlan9uMEyPkDZJD42aggRmnFhAA9YidjUWtKMcnbxZ
qFixhZveqDu/cS7cHEvVeibi0xZWUcyq+eJutDjo07FG97CKGNVFAg1GDHxrR5gTGtG4BIinUJv5
By5yR2tDNkQ6Ytgeev3B/Y5ijg49MKM4U9qjqnwIUbdlS1qxxDrpVUZgNxjOGuFRbBAqj/IA9WSh
oQoZR6a+sz8+3IzZJeGt5xXzB4G0ZxpSxoIbpig3L+GXhEOP1Mg+PS0x7qr4pCje3YkMEzN1Fzw6
QxTJNLFOS7Ei2KpNidilQ/fh8+cq6p5QjGkJZc+M7gCWJ38zglbegg/DdSBLr+/vKqFx0ndQgKym
uV1dnUkijEO/SCU2pBRK7AD36AcW2LJVgtp0vsilv+mJLX+D3DiwWGXmKT73VwwMaECIZFf/UuD5
38gfRbYT8UluSdjmVuEYNuSHixU0jba0a78InazK8fcBoNm8xNgtczMQLGkoim5gbu/zhw5Hotvd
EsNgLSDsPjI1thUJPcJvG8CcZ1VkXheDRquhkqoOUIF4Xr+EqN+q7XjcNTYM8+ZDQruVX2RMxor3
5k7pPoz7POi/mc4CcEvCT738cSS+Z/8Ct1u/vTKLJ59KKK0QxmLGehzW1req3+XKCMtB7FUZ1t0G
2cOrADMNxXHGrw3SHZYZ/vfqrCKDpa4h2Py5Ev8nQSfqrnNYxJcVEGnONgPCZda7ymfXj2bOi9RE
qfYdIfZQuWnvVR8/t/00DBspl+pNnkPl5sAiFwi414NvW2BOWY3JeXeoFEOOP1mzXqiPx+jDWp8q
Up1RXeQJHKZeOc3RF2RJX/9ZD6N7tmTf58w92vhsDUYVFxkUApe6wxjWnfww1a920A534AbSSOT6
O9OJEXJZMqccklSYKKkfnu6HcJobrmBauCOqm2XiT5bnODtTnQvYbEktGGpMgX/OZruz12kh7hdc
rCV40Ba/ET8yWw+N5JFXl64vjV79h3FetzYZCYQlQMSbewlaUnKR5uP2Xq81Fz5xNtC4BDZlzyf3
i1XcsBpqGRtlQjVjYpqjdowg9gbXF+GPboiS6/SDgKlKWDGyEtXsmt3YxNjXSBFHUTUnG50ZgDmi
z6XPKR6MlExDXC7+mJCgCQu9wKbt46e8jVy/k7QNH4cI406GhEQFKIo3MnPshCNMRgPGHM/DTNJn
LskBZzH8KixTMlLFbCa5k/yVGJVh7Kr29rvVRmFjihs5VjUrYPPEDk7JcTHPyvpQMfwxtS0LfHFa
yw01A+R9M9uVomFwf0qTO+ghpwkYKGy7y1BBXyYqqmxl8eLt5cz/wuQMM3++b/BU6uxnULGoGhlF
dN9FP23hMS3Dl3u+ACUlNNsPJY78EngkJtQtyUN04Zbw8QZ6BoOi9TYohtMjHHk9HgjpC900rMT4
TLyEK80x/vrzWiImeODQn6yc47gykSaKNZDebmBQX4AcxIWHv1QrzDBn5Bvu/gQ6Nl0qbwfsw6Qq
IsAc9z/ySURV9XayRC4ROTgBvEwZjfKzK1hdEImN+jSxY6niL8CbRY3zR8xkNdA3vG9Zl+JrLs/c
ewTkUCfdKTvu64si0X/nla+W80YCDt6cF1xdZitTeVPUMf/XvlmzPgF4XeHqrt/gKnYF91ZcyBDR
7uD21w+XO93RB8F+cYrQ/N20RY3nc/I5gYgmNuC+IgOZ0YU/O8NI1zbYk4x2kdg4MBnvpP/Kv6Xf
NkuT7/q3FmnSRdzL3Qkfk8+IsQOy9WA8XGtTKYmQ1KxYoYw7p3eGFwiAe4cfTyJsMfcIUtUdBRiZ
5uKngTdV/F8YvHG/9hfFRBEVZZrwpTEAvBIk7WMYLMfWQb/EKhgUWrLEGXCGGYgh63nPs8qWAJQY
OhNXn+5XVsVGjzxPs8juFB+jbK9Z30aZB9CmjJtAbhwLuIVGGHcadsjgcFSMP/JnVZEKVQYve8CR
/jwmp+Vr2VE7LuR9lNvK7UcUpR8sfNH6Dd87wq3THR3WbkBTVmjmLLyLm00GFaGuPxYwWTfyoYnU
R0YEiBuSw6GlfqepOu3ts7TpTOhyVYeNToJUaw7jDUpm6fum9HnZgTBFk5iLBsGezmolGHktykJv
iqmMYDKZt1somdhPv7zgBzQgNZYmc3QpDhbj7DuHoBs7AxdFRjfDxUcxeWiH80O8ddCtLfz8cLLH
XoaXuW1vnbr5M1gZCG15yrdINDhpp0utlkkstOwv3bIYIfWr0HQeWuXBnt2wYP1PPgfy8q4vlcyW
w2s1fEknC+Vmew1aQKOwtpTSxiRdQ0NA3NLIUSX35jlWi4JF3w2iI0JQTT/+EuvmSMYkLcSmfPb0
5wolSFAUwwcn5/vb48QJUL1yIuVCCUPx+1mcjEo23P8pnQp1ifAkPi66K0KvQg4/JyrM5qD1sUFD
s1PA+i6x4eQdijIfgNFF3apWaT6uGwJcp+CYvvpUA6VccK3qXqN1N6O6hPmclzH4iARGatxTJ8rq
7ijpvFgCIeLwUn6dbTaeKS0L6vLfEHZhlP4ysTP5BUDoZsKNzTHP0iReEFJmFK9WCBkXDguHvDRK
l5ITa6dIG1zhu8hX+N/pc9d+SvLXPujHX+pg4ByIaPEFrz+SUIZ0TWO/9XoZvHOz2odfF6FiEOXS
opxqnW1CKKE7oF2CL43yZjojLJmU/jDsm977s2aOcOY7O7F1zblB5vWzE45cIlu6WRV2KmBBL5g+
N0gkU6EgDJiJIm1VB51E4iZBiDzkdmywAID50GOI9TlmpTHarJalZOuMiG3PlEQxYyxrAhVYxwds
8+avv+pEmrXacitw77Dn3Egmj3H1xAZ9iv7/cR9JasvaP9li8rzcTCClUTCHhM5zT2ylihAQkm8E
2BhKF111z+xrJCRChY35rJH1qACFjyizSsNjYKbie2De+qVu6knCpC2wwL1zB+fn5IC7XXqUkYlF
D2Xt8UuaPgSEpOHQxiTGTAI/fCadaueCNQr9M+2HfSVXBuIOal08FQC9h6LcgJrFteD5CCrMZ0p6
EFXkaFO3mOfCz8i7CkUJQ6+RnFt3bIUDwg8WMqNh8Ilan9lLDdxLeJ8wLQ5hBnQS8jmdrBGmLsC2
46QidAcIH7awhtns5Jv9/9Ek76BTie0CYOtxLoXMX184OFBXsPfXedyiAOVovb/F1IhzyX/mxUjy
xgpv+MRUEwQSH99iqPRX2taoLtvASkzMsgb1j1zVRLCEGLVNDx0HQcoSJBmf2YeQEWZ9/yBmab87
qJpgGIvnnN5iF9qEnuxs8Vrt55RDxsuBb1VYsoXS7PWloCw3AcQmB0GmLTQjpAiWSvK2IguXKSTh
vSjx4Xa2Nj4bCJOn6yuUWCbpDp8Gf2AzL5wYjBh5rE04krMoFl79+fWpvM5I1jsBHjtieaANrNKo
hsrQmxs9+E/29opBawsQKJYiJz5DgZNkxeLYab4zdKtjbv9V63fvUkqv3X0BQ76/4iU3TDYPP3Dn
5wKmdAUwh1rlNXhY+18dY1GCPRN88k5WZiUXjFpxKkQp/itEI2ShOlIRI9Dz+h+CIl5vpPFTVDDx
L9Oc0+D0E0LuCMIHZ7q5bqyKPfcPin0LIDxlPiMVbjPtqiTPrmr3zyRZF/0s9YqwYVZyRwOyNxAf
RQFxTX52rnCJrospCJQnontNnlR38Q9S9ZWC1Ll8E5gO2QJiE+0juNbN8PA5FCqF54dyzgqpj9Ha
FWTx78Fj1JDBuUz9otDx3TLETgyhbTe4vxsrmUVr7+YRyxpwhMDTa3Gbs6Y7kNwvH3+ZgeKd+FTB
fZBKgYCDTcvDuasdKS1XTLWarfeZALQQPnhnAxqWp7sKYDBtv4Fkiv67zgPHTYQJYgJjfS+pchzc
MN+1Ei+af255PM6osZO1hPdW8xFZq3Naipa9A3GiW0l903CNupZN2dN1fypVeKkqHYp3z5xxMhrC
5zwFM4Ex7yWPItCe5jatagQ3+6YmPaIsDYhoUI8WR+pq6FCyRiLE1bFlYvT3xZxdXJDoHjBjkOjM
6qGdghxW8IIvglCTV6royq6su/IKMahtuB83vue4R5GOdLh3y9tDlWEw/wGfbswkY/DdkDll67zI
NQLsG40T314klVuW4jP7K4lcYOB4KgKYN4z96l3ruTND1+Cu0D6PwqkSixhS0uumaCmA0seyYmTB
mTMULuuRTv+s8caxdEu/C6VtIN9aby9q24LQNk7uxls1MW3AeCqT53RqQu5klPFRWsnAgV2AIQx7
JK3STACVDzQobATteH1QjKgRewWmkr7skycKT8cYqXe/e1jMbkWOPEiYAslW8Hak9hId3n//4tLj
E6ctQDj0UxmTuW06pBpuY7FH+SuoDJcK3QmPOf/YP4LoDhbkdvOw1rIp+ogw0Jr4V0QwmE7q0sGG
dkbvI7tttTemiW1jKvvyc11cFk8orUgTzCyypZbgOzXDF+g0WdfB/CU/p+LuNYMOveY8pLJKB5KM
wndxnQGglaQ21kMtxtUkfEIo6O45IlsoM9bje3f00qdW7xwcseBgKWPnnD5jTR8xyc3o9/xAgKXV
gjJ2GpA+l9TQbj5S78K+Nzcv5pMMyuy1v6Z7oK2kNes34Vw+Mrts/v9jUBFqZgxAXOl/z/pdFvcU
R8qHIDfWmZCJPs1WpNhgFbqAQCD666KzNYFYecfUPCbfdsknhhKYxgrkrqU47bBWv2u2koOAeqlm
gVeOxmMBx2tBs1//x8etEiWXRM2172csuwh9csKbkTF60yN+koUZXAUjHA+laXLCxaKi+VTCzKUe
klTSV7WqOtPh3G/Gf1u3VxKYOMwDtOU8BzSiKdmS8TmBwwEoqUUefL1Cd4C4x+QqD6GgKpxzkNIO
1zjGN7tGBm1YAT0bkSYWI9r6MybGPLHoe+5m2/8Ll6D5S6kpdwawuqoJEbD7yTbrwMkp3cxAOpY6
K97rz65HHgB9Zd0WLBAs3i3PaCtSfX0vhtWvM424XipwjmGucLJ/Dp9P6h3N5FLe6wVC/YNWh9cs
5W0kEB18JsFH9xGcUQlmpKlgXEZEKCCnkQtUsMPgt9EpuuUpeDWS86QYfKXuAoXmGcdfN493XtB3
b8ULwL3BH/RrysZbL2T9rCqh7YCAJIo0XjrxwKvYxppBkFFhEpwBNjNOq8s3j65IpbUKdr3oFw9k
C9qyKDvZHo2NOXkNF8xOlBJbwJzOmVzk1ktDdKKxncqBCGWHtS7lyuM68FI03LfXsqGleWHbRghb
txqyv1i1MOL07fbWDH1uqqcb3eEmrtYYbELgsFSlgTxvTUF4q6f9+8ywhF17TTPhK+Zrs8bKuT71
X0Z9G3O54DxNnGxevpVqGl8PsB8cWmdtvuthtKTF7uS2nSE/3rMLqJl9WNYAWbSl7h8uwWpdovJT
ngfacDx2AYMKjeGsts/e6HqSW6D6ytp9Uh6BZfq3pZoSdPz3Jif5EbejUvoJFfl4g6BrI4kVeDBz
2XPGrkGP092sTP8AWNdjeEoisHuCJAa9Aco4wxD5qnrccNT/hh8vELFgkXUOcHW5lCXcosHXY7LA
h4sDSL/uOtPhW2hdcIoY3ALC6cNDWmENT+dJtWqF2pHUSvFqTM53POULLtzI5hfpULYHDFJyT3Ip
o4PsKnJ2IkZKm1IdwrweHLtF7XcqjUi41lB+rdwkCxi0n7hNeKNT7NE3sXqbYRQeLQHWJ5yAlG5t
TOYZnyhDVW7DMvQXMUaj/x11XQQ6gtM3sYjQtfqnHBn1TBwk18SS5ECF9iD03YriBlorpDs4pCGD
yF5yyjbBOP1NB8m0254Q3h4QRDwYh0Bb1BvMcpP3HfCIqZQC3Rj7y6yToyIjJkZ3lpbeHvLh8CHg
z4IYjHKZMpC6Q5S8K8G5p+FPYonj7+xzti0/zwg5GJTX64JGssaDHiORC2CnaxDUkOhw5+8H/htS
LbFKg6glXmNnhFIJcrXcCFZomZtLI9Ioh0ivM4Txo+o+oPrInUmd64FM/LE3hRg5IkIm9/f9UNpY
VFg8CwQcr+r/AFlm7rhh2x7hxOccOwCZsBo7AV7Gv4JqNgC+4brYSGJ4JUoh6gh5xjGbHWkf7Zum
vmswPrAmEpU0ig3GZGTuIyahzSUIMQFfzIEBLMFyfwZG+zl0qRYFcBmXSL6VDK9Ko1fgMfwzFcKk
nXAiRF/VVTJcLl8yfmB8I9Ue/EU+md9nLDfKobxVe4SDddjrTVtB0oShkMXwIa6teQPNr32TDeu7
NHCcfabR20Djvwru9Bj2frAZH+ahje+wnOVQO+FnnpRDbULXjo+rsNlBQr6dBI3IJxCsSIYEDNFc
X2Z+Ar1b6SWe0MVDVN0N88ovLhJUg9fxs6HDajbC1Pay3g0mItLL2BNJ9fs+8wcExYFxA2/Q5vFs
aKEEMTURrqWIl9M7+iLotq71XcYJOwUhdL1q1ZuRqO6nS1bULV8vHsWsUkdjyVE/Tu1mqySdl/JM
IxlMGPSbRvlN4FXROZzSpKxxYfAUMMUhGpeS1Cu6Grn06wAuWZ8bxpWCBPl21NlzG19meZ3Ia9S9
Jxa2GmP8dR+GHsRumf77M4jgJCfyliOzikUBxjzsdAVwE8fDWgfelxL8+V+Y0edMU1ZFgnGVNDLe
AmDe8z6jCr4CIQxh3nBgfFo/RTGg0Azts5EpxIQR7S4o8Cbgtpuhce3tBjfA8PDhv0NFpbNca0oB
1Tv2hR8EvC0RLSJcwC5MJdWUBuQ3r7BvVPu5RkuNs+OqCSKqV313sQaZXtNVZEZOM37co0a84P9A
mrHoc51QxA1sE+tZjuovMi8k0GrgvaqMi4Zasa96FhbRoBJvp5ihWprHmca9Pkll8Q3s/Q3K3rjQ
sgMVomiheOkAQsh8lIzx72ZnHzAB6VbnPIMzh82nNOLqRG9PixC2tWGFZtIcTHY7fSgiN18QlRyw
ggsGbZyKFVSH8TBX0YCntXqojq0wfmEW6Tjy8F22qZLZzyKKw8Jmohrj1gUVRyKtdH+Up/X7sQAD
bxrdRyeAdwSym6frakzsPsiW2rfVdC/CVixiKc0KZiy4Cprgs29SHBCraMNQ8m9f9yhKQEa4AdQk
zmR9F0ZOyKf3URBQS37LQD+KiZxR00W8EV5CwyJsKavBrSgSb7isJXYNlOOqmqJ6Tf+GDe1l2hI4
iKV7DNjgKQovFhbVMwprWiVAXLmDUlvbzk5x9AsM/BlNghkVf06C3PPPhQC3hQb6jHHsjFO0MtgH
I6E8GkKS1N3xmWj9Q7YhUAvIaTOhzBak02IT78xGe1tZFPgq1+nsUb9wUeRT8F/Qj/aaJvsZ131Q
DoPvFcN4Edfh14mUEDI+nNv0q7TCJ+g3aZcbWalDu2SRTrhcqz6F4vc6I/i+YfniR1AUmbDUHXWt
b4y/8oEpBNEvb1A0S7NFR4rXROXe9E/E5gNEERfQIkHglrtIzZwpPBA902UdCN0AQnhamxiuQIzS
4lVkWlohVH8t7OKwxo6MHYZLWw7SmNCrSzhOkzgRNd0HaaOKFBYFt5COGDSESc9rgDcjUjNffdx1
18Cf6ilVtjllKsTZGljPcwtdnyeZz2vhNXXxkqentjQSmH8yWEm+9ME7aQCyv0n/XoW/KnIdxhg5
qBgtHuDhtO/WwHzMiCsMRC8wvZ1F2CY7CuEI7d1oIAAO1u0EMLJPKGicmwpWhTKsWfrfGGxd1OO2
6Pi+H9fA5UUlpngebIvjNJpXDp8Ln79nI7HPw9ehCVGEdf+IX8jTlje0oA0Z7wiALmvIteLFfSqK
H6Tw8hnTo4kCNcAzmb64O5g+eVvcKLgCC2eHzuCkn9fDeK6SsGzarrc2rfUJbodk87IvkT44mxZ2
3vkdJX1nZNJIC53D34aDb5UinySHjn48sPrM0HhMVSc3GHY+3FAI3nuU98izyD9MtOIjcpvtNAt8
4anuTKohs4D/z2L6RjeJ2d7Ddo7A7R+MkFddIBVaP3OswKVUBIBTX1uQd+P0CGDVaWw8ZrwPou28
3RXNcFUNpcSgXAvWNfcxEcvO9vLIKvz5i0WL80r/SfoFR0lgEmDX45OQxWdIKDhzUGaCpxCEWSHB
ASN2Fj3SWohwXM1sDhAKL4L5i/xgpaAtPt8HVf4UwV3cxLxICzeUJZN3W2Dx2r3VhwDiNJNGptyB
7fv70oovPgHIOh7pJsO3U3DXpXXv0OL3OItSrgNgSup4k525pCj88ieNLtn1yi/Eb0TePbNSpISz
nLjCk5nQrkxFQo16GuaDwjXTDHyFF8El03/uy7hf3WuwbV5MnJc03dFs67q/GJIoXpFFaYh3OswW
ctEGSfRN/uExh6Y8Qgly9dQmQfBex9uR/hs/FmDwrJOgM2ajseFu4PUPhXkAZR6TZFb2zWeXF6lW
+HXzqDBwEIS0h7roPKPFNau/vVGIArhs18eGlaT3//pqqVIz3NQpYQsNxOMqc4QhnfCKBBB5pw6n
U1V8ZhSqEDgL1iDenOcMKHuOn2RO0sqVrC/BX0J2GhIMzjCccwSHxAYXM8RnrbBr2+U17QqLL1Ve
pjm1yL493vNo23Yw7c9otwMH/pTif/RLgKRoTN9CBypuQRzz78Y/m1pjR5GblOWiBtrtkTI//OkV
HIsl911OwGpK047xl6As/pR5+a9WTZKyZ6CV649xuJEIb4/kw1D7dRMw/CvzxG3M3dTC57wAC+YI
LhQfKMoKp3g94ej3VZKxByjMcrx8BBtZKHw+r183nVaYDMOPObQoouNxMaagniwasAiEr/A2dQns
+fxyZqkga+28UvF1Pt7tj2XGcvcWTROvF20JJkE58SBDKvZvaQLevNYtdmeJemAYwHfPBMpdid2z
DFtv5Xk5HJLDmk4DAQOzSE21BL/oy8RxtCFrQWdudZuc5YahRcrsafohzxwPUObN6GOZghwPNHQf
2iA0U7EoYXjoruEEdIja8qulu7CJXodYbxePKh6CDzpzr9MZom2rxLBN3JYZRpuvPnEmrtffY0D2
Yijx/ZfoLm0pbvZzLAPS2dLTKrXCtnW+roRPmeIe2T/EcEsPzmJFsCgTRrrFopRIydSjvQH01fRS
XxJo8/w3sMOUFsv4yfsTZ/wpZyX2/Y5PvtRg+XC/+9PyeqSw35eF8fugSrWTOHytoNDlg0P+gTaV
ij/8vseA1HvkpdG+ighsH5ViE5SAjUNtY4CMGZS8LTNLkP56jr8p0xz8DE7xJNV024ebIOqBVlQz
jvZlSY5hDBJcylDojEizk+eCjsAjyZJlkPmmT4hp2Tq+WqPS4rHDokMu3vRWEukMgPaSAgdtF+N4
ndf2iCMCfE5tBhU1cp511gYPxnqAr8Jimr26iE0eubIBp9siuklSnnf4AJRzfUYQW8oubYJZM9c1
EhbBM3wSjm+639l2P3wsCNBk2I6YjrPN3EBVVUjrSlhuGPPePmiG9yuV5Le9F4MAItB6PuwgKVEt
uwElbFgxtxtColXj8w3GM8URF6SMmuq09xy8wbyqt0gg+vfr5E97HdgqAfHpNpLjclqiupWVGwgJ
T19xtEnjG/K8IqXgcb0Qgmh3xK6rPITM24VpDKY1wHhpxVWvNAzLuaAw/oFI5+1tZgeqjlIAbbDB
P6mQYwlLbZ9kYVPFjOrrblYbKyrxkUMz+1k4yUUFcI2CngLYqFu9t/pRPOworgoneL4S5kD0LUC6
AKAflHehb6SMdxqyijrz0zPN8DdcY7QQ1kBbTuhSYBbhc3/nFJk0Y78UE4EvQHGGGIZlHj762wZL
xXnvEvotTq7Yj/etC4EOXDOhGqCN0fMITKaRWUzNjdHTknTTLOx0N4xuEELJarJlbm5vizt7w9/0
joIjXrdQtPHTF6mykxjBT5zqGuDyK5/+066IsAdlj3B975KP3Cf++2eFs+xGanEF3t8aHr0p11VH
MQRAi30FThxYRd9stYKv+REqjy8n09fQQ0dqgab//EwW0/NsDEc/LblBTRXXhjlUvr2kmMq9tI8b
5R4BjY7MoOaSTFL0AftKwFtn5QeF8G7fTgfy9YWnKLG0f+7YNXHa3Ld/+awHAr1pOa+ZwK7u1QYY
FiHZEt40M/bvLz/AkbPB673eJkVP4Lzrb5s0d7TR2vyGy17bx0zEexmWTY5tp4x8F7HUy2Am31iS
YxVUARZU3Z6i6Tx7eUrkqeTdK/wSS33D2VMIeNcnYxXpzqgrNV+bxpkgSjHYGZVoHMALuCPj1LA2
GR/N+/2PAQVJzTRSYk6zsExE1nFds6+PLIPVJhmnZQBO5i5xUChJ9S+FtXQ0M+v5Ib+DWyF8qOom
q1EVEhqHkchgPWbFAErOS5Q1aQNOx/1vccRpwxJe//g6w0bUX4rWTshhatEygEpNyIKyrSR9sKCe
vonjQjmUALTMMKs/RChAhPZcN2bYrd8eMEgZzahjZ/lvrn9g/CxbeAA0Z9Z1e7FrULlTV9MjUx+I
F2E3Xjckd3NwxNGLFUeCxs88RUtDkYJ91tBhK5YJdEvrT0JSyTjdogqJmYGmZzinyN27fYBz9eyv
LVn0JzstbBL16Ss9ZCXi/J+jWMvsG51LEg9BJVRehJv9nTr0eUuxUJ4QXBNpg1v8bkekUnwxJWv4
h0tTzeGDRpUnOrA8Vp+BMDrPqB0GmmGvIoBhvdNl4is2IYK455rRf6tS1sLKfCxWCkU/ZLcnHJjH
V794oe0MGkq4P5NBkjd9i4MjHnBoBhzQ9avxrOj6cBtU/Uu9ArWpZrGKvwU/Q2JRSb0MSmZGBsAz
H8E8iH8PRHV+WoJZVisEfyuwv7+jq+TqQCncJoCrDZu2HN3z7tJUusSdszf0gWXyOyEj1db8C/NL
WKY7QPV/SGOjzZS2Zv+jyPxEVx0+LzCiXQ2OpN/uN7dvhP6Mmeh70b7jA+za5651jIQglSMzdttI
Qz70oBHbIKwzUUtde/l9ozVOZCGPBc0UC7Tv+2Txlsavql8W8BDuzoihnlH4H6SxUb2LN/1B9a/Q
oe+wfqNxLPtv5xomCvu+EO58UNHpJv6dvFyfPhy8cnh+eCxDHFdtut+tPuoxKZVAUDFJlGk12+f8
8fksYJGyWV5x8Z6oblN6vZmbS9b2kS2D6+K3olLQLEArbO9wV2RH9EBH+XqQMxV9gQtfOCxDsAwi
RhDcMbNbz/mbJwMP9cr4Z97bH62Riv+R79Vbrpm15VvNA9XtnDujoip9/JMkTnezQGgyB7wuNB/W
gH97JPLgSVXQdaY9xwY1vLaKxiqA7Z7oR9W5THoO+31+M861X2z1/W0UiOpEw6civNktKQ10R9AX
7UtfI5VR/bvCRN121j3tgPaZcDjr+Zfoobi2AAnpc36eaibgnbPMZcnzxZeb2DfsDeoYzFELXt4Y
4tnUdfnQLPbFpM9Z8O305z70bgq5Nz52BJ0zMsQhoPDXsA+C0CMbcRvl0M4IuVELsZ7qpbuUKF/5
3kttk31+VmNIkw7H1kmi8hzphlKf/trpCRKcd2FsssOeNPiX4FJf0xhtHdXQvg1cp5a6w3PQ4JSA
ZKGUCqcdXErDNv1tl0TtM2YTH2HSRIdQyWmxDQjm0xPQU7cuoefQ/XBWsnCZqX4NW061MrJ0+Ii8
AjSFTv46ofHJHDSuCUwY04CL+9DA8ia6boR6pNtM//f3ZUrui3IIJVkEovlHso4p+4+erXpY7ADb
eb86yyrct8yPseWofctAJbJDJILqsAhFO8XpW1DK/94QGp2s8fzZ846ILNPjtozB8aZNeoQddo/B
Xuan43HG7+5EuY/INUT2DFkCsvnCgcg8KM1d+hP/CWT5GjD7jDn2UeWgvSU/Xl0BuDwwzi32L6L3
Nio/DfxhcSJN7lcNe4PjnmXuakqqk6AWalBLz0uW2j3JxCCHHVdoaagQKN96ll+7tEFsqtWVR+1H
fh8VW30GdaxWMHuWjKPCp4ht6iZeCmEF6ofc0EBx1+9HlZ3c19HBhcjZWWqP3WC6sp4AiTxs2P3/
WmgjDwadOlh3TCZI02Zuzf848dBInXZCh0AGj9kRp2+BznYrFFMnb5AItEwe/SeNglwIRdk3mXOv
In6Iw0bNFQQH+h7UN0NHG4OW661lpaM6JVl5WNf1otJVe8iTnLytxS7DZClpXIXDQRPQdnQoTMRa
qnEO5ryuT2ksqgPvLGJGzfS5JBXO5XbPr7ZCP2FpPyqQyeYbA2piSeSbt8oqaRNOPs2ap73Gdp54
xlMgsKlYVty+S9QkuyQpX+2/Fh+CObtjcQSi9V6JICoZJoR3p4sxidQpKUPmGQU33YC3YRMMCCHt
M6v5yw8m7xA1EqcxH+jCjB8Ky4ixgPibCUTA12xIyH/9G+1pSw68soJJJvYKSDDpxke20/hM8Jmc
QKnXgcOFl6oQWtn3p0aRkYk8boeNlDyDkDupvhRYtMEhwIMU+0SfoPqVVqVD9vVi043YmDk0M1rc
3VG9fvxfJ2fko9sKWP05Me7E+G+epcgHkN5z3ANS+YHzpd74jxPzZU6S58JcKMXBS+KY7GihtW2b
fGC9nzq3CPX9eZnaSiESqMJDCemy+XADl44AgK5qQKZ1icIOQaI0EkjyVNMYN9PeY50UOUKkPCzQ
vIFqP6wgufh4cykT6euowvdWHWkUSqYoIDWAYLks7QDroPyejS9tGM6w/Q0RvxRstVUZuhevqD6M
inEUYIx/0ahvnwv1SVu4ISH4OZm+nLeE1vjeo+Uz7rzuJmw0jzCwP4ZzEQjR7mo18w8G/oIgo7z/
zo3BVfb6X2rWIdeJtOblqy+wVyHrvvca70bFMSp9uUAW/XF+TVi8Eq+++7Rn3VmRfpNXQ2EKS5iG
Pi7XgvjrC91T1Xej9EynheIcr9vS9VKqe4mPrVHwUWMN3U18nvnP5sUNHmptTvPngbnQ6dD6Ibze
3WqkXdZA0ErFO34B6Lf22qqDK339NajbN3FbIqrK/UhQIcEi/JIicY0BLhJLI4RRkFVcvTdFpK9R
dLmfLl3cZ0H72baYzhbjQhf+k5y/Sx73JywSLu+WFpIwbhNJux88HLGR0xdp6aoHRsbBGp5djNgw
GFro2Xv8steOQyivw5+R6N/tzhUrdNNWrJ2Kl5+npkTLAROM9Topioebzzhn47a1lWnW8wxCSYFB
QWR7pNEtj6IJOHikpb/i4LRexnB2PX/o0my7UO6oT0GV1Q5g8QB8KaKXQoCyrSd0egqC7h6tG/do
URA+ps8th8yjJCLHVZK/wA/IhkuUJJZEuAQlzOY5Jjy1qPmpSuU4hnA2NtJTRruiIbsEZhoWvXa+
V+z5AS0Edda8FISd+2cljMHZ+sbKKoAWA2wnHxzpDfIzhSBOt5stAgm5gtoxotX2Ks5vpE3YIQnP
cU9CKvoOiOpfNNtEnc9h65New6wgenvKsLxnOuYgB57KhAlCN8PonNvAC3jOr6dbX0bAY77UEIjx
R1c7I3AcYIuX+b8nkf9v6cnthYJCA6Rxx4xiy9YdgH38uYKcIYSstKHCdBYuTJ9tUBZnTV4xPe3p
lqvadiEziq6fsoflNXgFtXB3O7Cj2Dzzq75AKNUVbdqFDtBA+7M7uK2aNTPx22OYboe8rvBx6bkQ
sMpnfXOIvoJ1j7Tf59pq8FCa58prNJ1pBfhpkFp68NCFUnV1KjgyxMJpVZ6tLsDNJgyn/IX3J2PY
qDMmgznZ6pV0+2DUwZbbxZ38LQZQre+9rLKXCH9DnqY5A67mOslwTcfAnCMkhqKQ0trOBnuJL1Nc
BMET5FulYdH/nFU5TgdHKuqzL7AlomuVrLZzldUf/fux2DXKm0BuPm/tEmxtKGWsNxwt/ZC4Nplf
w40XbDtMElhhLpt/ERGbUBIsuv8/Ok2zMWoi69B2Xr6wRAakh8hk0ZBJZS5w2Tw2SRxSosTmUDsI
izRu6nfvfl68sPyzNdjfELfszFvFTjwNMGpSST6NgpbrsE6yh0ls+tMwcVZq1iVl8oKQQ+lNg1Gf
inHuuMyaLKxON6O94zMz3SUpyKO6WYVOt00cVoyuhVnUvfbAksmooBHp8tWOdKBNcAcGLlS588tK
YYW03QHPaDuGu2Ge4w1cUhMBKARg3xEKOvRRH8kBMuwfxyfDPxn5f8b3tUII9vJRHBU8gRjo8WoM
txluqyGzNxbnUXbmoU3v/TLK2/wf9RT94fNUjy2Q6V/WcS1XBiEqb0ULoDa00HvnHlaTrtNVOW62
aYwXdPI534JFJhRE4hD15rt3F36aypsPDb6mH9ROK3hK6y4lYETH79eJnbnBmUkqsKwV80loFJzY
4XfaNhvplvmzWSltPM7ROGBoiYohCoAvS4GRurVCheUo9rjLHXIyA79J523jBDSurJhrDP/kxYyb
QNon3rESRonhn+XdBYp+VGC2Sq3bW7fUIFOkvAtL3fpvOoYsT35p+zfX/lO8mHoPTOo/6tJK42Qc
P0tbyYFVR1p8CohzIpU0i/r9JT0coc4UdfAYodmjyUy5XtTD772UBPGNwmqTWvSTzc9rfJ9DJB6Z
SF3ko5TXA6ifbvHPi6otlv65sP+kYhjwGvwhgAAXeuC55H/GeZZBl9F7/AgKCE4xph6nQB6/NSON
x93iSKkoWkMDeHXS9NmOiYac+i84f9x6IhRkmjBeoX/DFhTiFw9J3dDHdg3qU+CwRtIe97ZsosuX
1OYFs7JncOHVabt3gNyrHIZtydBxtv2YbFbdjk8s4FsKJBLbi4FAIIkNNT4pTN+Zw39RhRvn/lhY
rLUg5iJOhP189oWLEodjWmbjQPsfMv8HwhIuE9MH5fgBlTErQ6gGaQY2Uc+NlGS3Modj1BkGheRd
o3BED7bRvOQsbiM5DzZzUl9ZxQCNn2MrQld8qJv/jIvLd7VQiGmqZeBwF/U+qWx8umAZ62x1irW1
A3Y/OQXv+Id+rGdIr8hpzgnCw/r59c9utYtN2aKB6Uzg7f8X6dUsCmIRiIf0wJ7xvkvTnLsMiK5W
i5mgaVDdTlqQR38dNXX1uS9Hy+IQLsVPirSojptnp316A9XRe+cOcr+CkaIeH2WrWH5l+pDnxRcm
ha5c2JxP+4//wiieLxD4QJY0kRD6wWOcGMwypxjDO3eLEbZ3D1uz4RbjCZQXQRs5vIoNFsikeMiy
Rh/2KRVHUPlm533UrsIu7X95eg/b3Uu+fIClDnzPEoUh06uM/6b6RtXB0KTHChgYjFY8Nb1obcwy
cDI3SNpIZ0dLFGdaSR76wXniJOwkYOIzaqrkXMz8zEdGiLGdDpe6v2Jhp/GnCZA3/37pb/g9KMCy
9b7qP4TsqEHbUKdBC0FMe8dc52q/EHExDgItvV7UhfaXieSL1wdJyAvp4p2pcDXLM2OAfYd0D2Pu
GMSrLgu5EsK6D8n5NFeis2sC+E3cmc/nrfD6DpXG5B2OB005sOLmTtHev4YT26lwPZkc29WZvfj4
UWEzN7jV/+CNfKWCUoeYbqdRi/i6y3qEdKBiLhE+bZhznsOK3aPcWLZuq4X36EPL+zs7HeeHya5P
SaP1uVFb3VeEjSJ0tbLAKFD2bcFkoBuBzKRG8kFnXeVOL3tqU4fN/UnvF8mcmI6C+mCH1N7rE90J
AscTZjSXzp/ixyd8yDHN2prqevMHiic+9Yeoz5ItIqV88TiNEuzSIeIcMkgrv/GBh5lVG59vN66f
/RercA4A/flkq8FOnTGHUmuPIJm/5Idb2kwgEBLYkjUq9HKlptlwguVv8bWF9z+2185Ng/Yz6ZTa
RNTtXNhDcOsKBvnKOkBhvBq8ftqzp5ftTMKPYR28eEEnL1Y6DS4GpwCzJI8WlsoBiCqUubNyeRRZ
RIAsEPJ5XMSW+aEVYbXCRqthJduM1ftEK9hIIE3jRT7jhcp6+Qks8tyx/pxPU6x1xOG77/RrCIQm
aMYGpfhyNceyDc/N/tIp64Ci4IPjv2AqO5D+aMb9IkluSsAhpS5k+fvX5VVkPBs+sdzS+bV0QdzL
Ke+O972j+kXmLIuyJAf5q0730y4zdk24xsO5FJ0b+RsRbzDw5FwC8d9dEfA3GLQdMtw9bUEMx/NB
dZHF7cdTIrt1LDQvv1+C1aIj5cnr7BNZnf8AnKfogEp7/j32tqf+ePuYq3SCLbVAGIojUKhwSLiV
piWJlXYWorgR1vTZE8pUof/29Kihm+w1EuA6t43NS6uhYuklM3exiUFp8RHVbFZuHqamz2vdXzp0
aHcU4hHHHr9piP4hQ7wtSDPFGWx64ALmlG/DuigsWSDa6aJS2MhveK4+zMFNPYM5xV4dlQjmIjba
2fk9O34jWgecaFlhbX5ZGf2tdRYF4uBdtORFRTUisPDSTWkTUmWkSf27lHOVy9UINtfMMG2R5Ocg
NdH8J2roDF1OuhaAGMSjByZfKrIZjBpESoG4/0iajLVC7livvNzpLhsRCvGB78cmEoNHzucaj9da
/cGEPlDNFlm5cJsxbUPApDelmThjB7NwLsXT0Mi0Jn8ZK7rnuaCXSjIEO5XRDKQKqiof2lTMBk5c
ZUznrle+QGJ2Hd/kFgZLs8TYS4idwHGMwGVD9EqnUNFCWpfjii3p414ccsNqx1cviSnp5M2IJp6M
/TruYGibTYnyVgFs0wJk5cmnOwxtDFED+y81e7XCu7DcTQev7QPKhVCJ1FDN8OcnpkAGjTS+AGbn
CzeJSYoIeKlIE2TWLYTyI3EDM2WCL92eDF895DicKFsevDornTm7PVoZqVWgCBTSbKwnBkvSicR5
Cpi1U8azRF5YTBD5nMZuUjr+6/Fxfbl50HQ+fqs8gh7E3X6oHEsK8vBBLQHLMHv9jvZx/M7k+fXG
SjciA9VD/r6z8KgYivV1SCKBmDGdkepAj7UVkGyeBsRAV+bIeFm3/UzfnsCZW0zy5Tpohtg7mMC+
+iVr0eSWYevDAR85XaDYoqWr6PuHFL60xFBtfIsuRcYnS0DhoJOIuK7ZhdcUcJMaG6YoLY8YG9Va
x5Da7/WOy+HugHZrtB6PvA2HdcXCDhxuE3BrvygmQd5yxqDmfXAJKIPVY+lcJY9jR6rKra1d3Wjx
3EyfwyvLP43+pQbBVTfLj1gNh4rin5mMj6K6dX7wWIkpOtrUXjI6Xtlvqd+suG8JoNP5hLBRqQpy
OiJ45DTiCjlF3SGQv2ryfy74KuFibcrfXQAVqtvfi+ipuYZVlMK2ioGT+sPMw8/87Brhj7hW95Yg
OPJU6ew3E8o5ly4JdG7CpS+5pdchylkE52ur4vEBg0PWfto6uRgPBkwKd4W6Ql0zr/14K5OIwvw9
wW2vbQ6vm7X9kqLOQexUTsP5PROEvPR3RXMUec61yo5226MmWW6AKz/LqerS6UiMjlQHPS9gOdip
OvsHuIvOZYGAUIlvC4wQq9QbzCqFts5zaQXLfU58m/PKUWaf9nX0BBXakfrfCkdje1JU57qsUEEa
qw7iMKcJZwq6wYoj3hPbGc/m06cmBdzmB3qQZWuUhPPEe66HGx2tU+g0IHFP901oS279jipUbX2J
o2OpDXXj9zwWvcR8dpSI7U+S7IrmGS5h6g7njhTytbqgo3hin7XttwknzXiueWdYlwdQ0yrP4Jj6
yAURWJmMoEt2MRQitCVf5g447e5tawlKf7rVIa763FgiWq3fDqOKOcOVg0i/X2hOkHv1Odsc3Dr5
okO5z4OIIOgi5DQ8mkSjBW3wAAosPgF22pJj4dh6s/S9QbDVYMo3qtzmL+bPAUockONDEHfsZS+t
wVX5EpEki3uwMOrcKHvYK0rN+Q+4bopi+slmQ7rF9VtfwXVSd7dpja410SYyz5ExD2/NQsMkmOGC
8KN75h2BSiOZTZLHjHdUGE7AuAExey5uKPFj1XXe0LZHVvFd2NK2m/a2cgKSIQzeexoGlTbNJJDj
HbSdtQf4fkpN3gnm/4VG5bJZrJr06Q2RMIDweadAy4dENAbGs7rkFVkSci3R8sylprYTYZxYe0gR
RRmbu6ldVuo+hipQn6s2938+QS7q9cmffKqr9zFWI4KjI/mtFPuCBAfkqMU10RlsSzRKwJslEEBT
9OVA1a4QxP8Tvv39E8ELE0Rxtbx3BQmdCXDhBEOIl6yZap5pe15NntCyn26zASPKjaf/c65R8oNA
o/bZW9y/9ISaQaOYsuDFQsjnj0GOxRx0894icb1eoWV/sw5qJ2SWlie4UOUEBdp9+vWPqX87ztyy
Z8/ZvTvZ0MDepbia2MLxI4+GEmg7mPwyMLNHWZP8sb9rWaNVZHvhUjSvj/XJ+wbZzNPfhB9zYKKG
wtQyODpWloIrkInGkrpb5kp/T9jgiQSvADIKZBmwoUXGX3saPCqH2xPdJXT48CP963SOVqSXtvPC
Vfa8STdCCKOgcDey+VBNpDvdjD5FlADhkv03lv+MsOC8m8Ccx+zx1++0nzndbyvD5KtMSVmarM/X
u/YLzdBnsqg+CY+ZnHVqP5UqkE4bKlKQ8m4Oq/Ff++sAQ4mIibNDetEa5WfaDdxkopTSK774v/lh
VFkZXPcJoHuV7/5MNGdbkx6cn0lfp8lKDlkHL3loLAZm+2BRyBQYN60OsCDF23dJ2cLpt57I4xiC
G0Fu1omqXl33T+1CCHvIqhCN+TJgtRsK3ZB1ouDMc6P0oitiiYpbSmWzQEu8zbhzCcMY8uPi5dhQ
Og1TxbiHylJEhXpSLMforM8I90vxvGyem13BxxSR56RjdJi5RpTnoKDbN+kpYjvJYfcai9EsKqfB
2S+KGMlmLlvbOAYV54RRlH/W+EnjoK0i2SDk766cZePIWHWd3ysbZk/WFNXjEmGsZV9U4au0o7SY
T6de2ckeqZi/V3SzBLO5VT1HjCNMahBsSvTdFDTyTipOiLZMt3fKiE1VuNbR7T1BAGMMZ86OKg79
mLFAwCjFsIs7WYepcXnvch/M3+AHW2clFs1uVLC7ngXBnRnfyXEFr8SZYF5nmrQCFATXkM1//nHa
Tvs9W449/d7R/D9jQJrX5ISCuI1TY1kuXP9VgxR3UaDUe7car2klDAA7hPTqOWuBw85xFCvmL1mj
YlKUaMRnI1UnB8TUNDZDBytzw099qRRFzWj4cxD22Mq85Fbn15qLkF3cAFOb7pHo0+iYuCi+Vqxy
aOroi0+W5lVwRH4c4efebqdMwDf4S1itPqU0oAo/BA9jTWQaYEgKdI65Cif4jyjmnt90yQMiG66l
LI4XrxjObAVc7XaBHtiHUcWtCwPchKG1vCwsDx4yh9snIiDyzkjFX5QH+pUElq4d4PoPps99G4ed
EnzQoziDWdpBNpBT/3EdgGm8ZxHsDx0FmW10ttdMeDaDxVv4Tsei1JddzfFWTAwG98Bmj+St1Si7
/OTXFQ9cZ7Is6B3bCtLWsjk5bv5v1Oft3Fed2GK1/57AEfzGOrJttJAgV1nl3RXMg/jw6nDdPSed
jwS+s/yVc3wLr2UpN6acSXhmAodwOm+bto35OshIv6qjTirlBUKKkojb2mU8ndZ8eLTW+XlqjefG
K6V4Vt2S4jHoG7tBA6aCj5JwwABvspbP5CpdRA6fYfK77yg/Zds/5jOVy4p9+9F+1rl8bWeZwuY5
pEW6FOMKZzyApoLdinr+qebki6urZ6F7Pj0zvZ/bzCLPFnz8IXAA7ban/BASz8r3VU3ntTOgwwjo
5PtpcvXPoqPVP31iJu4Hwwtph9ImE6tLggrnUYndrG+vx3n1F7UtJlIDWoAaVJBYhFwmqfNxGqCP
K21DImLS0GO7qr0562j/0e+WRWWY3MikQvYZnx6B8w4jaNq9roB8ov3sLjmnK2q5+gFoaN6cXmi+
UYElRVn00X29vCGzCCoba05avp7uofb6Lnu13krki+WkxHT8hIQeLME17qBc220QatkMAWDWWAuV
iKLkGiZ9NHp60ParNY4lJyxbUHSz3ib/eGMQ23aA2uGWubInXWe1HslStIGfmLZO7Ki0NdOT0aAs
fVXYhftCH0z6KsL62I9nevTerDjRYesAPrpvTm7DJ9FK9nUuN/A37BMvAn6CCGTyK5tzBfng1c8h
XtwZeCGYZTEfBZYVwFsXnnlVje6FX/YdU8n4wXcYqAEbYkM03uwKYqjk6ZdXV6PCV9qVnVPdZaLY
iBpaqPS+ZTr9gGadeFpUn9WSB7RaevtLvm0XUysRaFC5k59PI4OtXjX+0OBwJoAJhdqAEqK921v6
/fcuqfLY4iA7NwfsBZjd3PTnSB9qrGBgP1MbHHSKyqaIaXu7a8U40FDD8gusWusBkQxOK7nQ4qKM
XDzkj09/eU9nI9nnNY+7ywWcxgZbfHTnmIJwyWTI4r4YulM3OhmMMqj63ZTLXzOqs6sW+R2pf4v9
J9uAKAxVwH6LOP/B+9RG+w9e6Xl6qryzJSO8ORv5flXGHHtDBR5LW2CPkULFbjup+dsDE8gKUnGp
DyEPza1AZrfVPuVgI8zY8HXC92D/Wcz5YKEZCvfTeQSH9efMXC7aMrEx0UtpATkD2oU7lCF37ub1
wJ8ljg07wgNT1aQJTcjK1jOaZDGWj+iwWUn7XquxmN4Lwnij7a/DhdDZpA0AM00Bi2KlXMzfBtv8
OQn0IlLVDiyzFR+8aUmw42hRoDfeD9ctgDlbWNpRw/NsXQn0q2hEOePEVJLwXj64sPU5sd7QyrS1
7xYreNGyMZqB9H8Z9Q6Lp/rhAIKjk436e9cjL3ATwgb+m8B3sn8Afejs32C9NcetWEtEKFViYo5C
101C17d2zi9qZaEvVULXPY9u8Rtb+7Rl4MVIVQTkBHbV7FwdwtNRYD5DxicBGKku5mXs0l6AlVVk
F2gBf8aw7MxA6jpyahTCMnMgPH3Zu6CTkyoV6tt8rDAonmmgprLFxf7ctRgyhzzIy18DeNvyl6Et
pEcdCQTW7tRGFW3Qyo+GWShNYxPL6hAQtrCXk9PYoHnay5dGQ58l6kduqsJj/PETknM+SfDHLYIc
a5rErELCylGIsChDVxdF3kF0gP3uyY4mfa00lqV0Q4IhMPzRJY2yPgmCCQx4dlyBowKZNwnSxkxX
6jv3X7hbNI8sJWQ7MBn+dSP6skIepahSW+HgL/y1chuPXsOOAk6slKTUuTILbTxYAE741sVK9keI
4ogDwcxDbUvTfBq4Gf7FQIyRSJkiUUqKJ9DC4Vr6e0/KFuTIBFmdOe5n8tPV5eKkldhcq1y58Hxo
GmBmucvY2E+8kk3ILlNwfVVgbfFG/7Q9HaisLhICEKYFHh0+/MGd8WxGc7FGeo4NJpGSwekA97a3
RPit039WYAkZIcf5srnilSBmJdKgDyFxUaDfXbd3snClCLd8nJnzHEAWTX1CNjQtF7Y5tk6G7m2R
jB5bofuDRBWi58QL+/Y5FXOQPsNyprOjY5dbXxKRZY8gY0l2aKDt8JNXHlbe5PSQvrn9zME8JWuj
m06cGHZwDK1yyAienLoyFw27ScVxE9q8RhXdrNygwvjLzc17Ro5XNl8VIpLT3c8uzyPGVIjCTQQu
UWKsCZJ71asfZn5KuRv9BxTWpjry5pgVKxy8Xigzj+HOljXwGYxnlcpwxdedLsCAb1mWpUgU70V4
ddFmeM5UTaFYjGGtrCOQkE+jo4oMX5Is3LKxKFy+IR7WS3jEkt84YtTgtopbMRdRDoTp476HznSj
CXd0ylR6cervnpBirjdLw5mwyMTc17PWVUf+ymDhv8qDHdR1jBawT1FRKncbBQ3fozrSC2/Gb2J0
ptgrTUdd4iQw9ONK3q3HDfSFiK5owSKJDRu3lSDl5tXDn/+yvX2FdmiTQINzTB6ZaRLWk5T/S4tn
MusYebyVC3XRSO1grioo330ps8XZmXP2rkGuylTCjZhAJjXhwxjjaovXHUyM7FyhTOGiY4lR7AiY
Wbkl5umScB84GwiN2KtQ14U7bjPOQOSQGyY7UgXKueiQhRSN2A91oWzu2cq1RCRTv8j3VHeZzE+R
JR8lLavCK0XEn4wNc7oEd/X+gtQpmJj7ZX9H+/iZFsytZnj8iSov6oH5Gfu44N/p8hAuXotVGXGM
ycJ60WvUGBU0kWaaB4wcEwjvPSKc4CWAVuTcoYiUyKBvZNjlOi3i4Xu/f/wDcOnzN8GzdenysTAO
Nuv0f8Q5XxYDFU9kPWvvbu9XTUsP36sAWbIlrOLm+/casMjr3Du7ycF9evfZJHZl0J02HdezVOfk
qndePL/5kVPUGJ7BbZjjwdz/RetjXuFDRCcGx6AYhkEGA5rfhhx2DbmgqoQA0iD10QtHZQFYnWwT
AFRFKdofZZ7wn3lcUOFXvvs1YKVnpehMt4KzSdXgtQ4bUgR+rZKf239YB4CBedqtNfa2p1s28hPN
TyLITS5z3onK1+Qqw8MdX4td+i7N6q5MCLco1uWGizI9F/6dcjI7ighy5UVv0L0gdh1RfngW1RKQ
W7XlG6uVFvS9Uodz44aJ5z34Jm6ierOPDfluOsAlL6XYXKziINQKcpCM3XzJTS2tlotNjjTJY21T
ZrUDSmYrHGMrXcFtHFnNck+FHcFONTvd8y4VoZvUHrB0yEAohXcwoFEUCf7S72/kvT+H7ZSJ/hNF
TC2f0IGCf9ZDbQqs2Hbntf5/Y3E2MU+1c9FmhRNo2MW/vfA8uzw9Wr75FCvGu+OO9wueN+QJ0uxT
ulZx3bMmtksYVMQbUoepQRxfV3ag8mVBBsbbi717XI5Uvwz/vmalyJPdZL+M90e7uvs9kpmFxEp8
qS5WvsTkgfSeID9hkD6pamM5LPYK72MVO6rrzspRygTtmI24TbR/x54F8gcDy0eUmMxkp4+C51nl
jUVhzH6lu5ZcC6s7b7y4O+MNVycd3hesNImbx7ecxe2P/7SZij2CuQ5Ns0r71unziRtCQ6LwXZ/l
qQNB1EyhQVjGMQ5JQTEP/x7PD9nj8GAC1+Q3dSp/Q8j0IQ+plSEL3BCuy3xF5qL7zpTIM3L1IWmm
mbPqO8odfv0i/VDF1Ka7Nu+jNZz0NF6ks+d7Mt8pBnJVt0egi4nkKuwUpwIPLYukrgPnIytF46w+
V1i3dDLV6tL0n7r3a0Ese9TxDNEKEv+uH8FbkFfuEnKgqM+/wMz7ej1UPuRFndyPYosq86WkzTEa
WSkbfxANO07iE/4XsPl/0WWWqL+A2TQRw2KELlMoo4KlovevMsKDP0rybqJPJHezVH3GZ69LXWkD
pHJF8gS8fC0MPVIGMfCF/UcIbH+EKm/TwTZDiqlXC9/kQFnvnekZJgfbn4M+WthyBU/dhSY7lP8v
tjKcNElxY8296drrPVjpmeleK43WnDmKkqS0KEx4tUfVoODxJRH/NlfR7i3ZeATAWhBZyW4sCMdR
KpgZ+XVjZJoBf2uFfi39Tb4TOfv73zlcHU4uVCiysXfAOyhFQTqjxs+pySFwjNM9y9vqXOQEraAF
oCNkndxCVF0JRsT+QzE3IEVcYKoX5K0/4Ys5zhZ0VyrPX6LiVt1WYS2aXrimeSpp1POdmWlWjCkK
CSknD+eYb3hX5seLvCxa89cbOn2xCqTO+yV9Wi7FvpHX7A6el5mf0iHrC/Ns4SbVvr4USBpUwQLl
IZGhYhB1aV5jMjqkkW4TTpV1vo9DctLWh7aOv7S0g/sy9XmA7Uv+8n3GnyOcRXOAYtC4Ip6dnAV3
LqsBquq8U89K7JI0EfQmNkDHxT92lgC0+Y9SjrY2/FRSNV7HX4URWcWBXbsZtkAgEBkK84NNjVe6
NS2dxkyQjKfQAx7s66EnZouBRRIno4gk0RBy4YjTFjJKXKisx6TZ0bpR1qe2A3yChG4HcTAD6dpa
QWt/r3p/sAlAuqvOZoYO66BYdYqdP72kRchNUGvChSabN/YVEb5Gk92LpCwsTN+LWpa+x7JNU0gt
RRX/7Et7I8NoMn/nTJECjkT6omyKzRRJdRRpHguyf4WvPcLjiX2NAUCVmbzHm34AC0N1FQylaO5Y
douhMDLOEznMqkK3c3DPHnmWa2O71kTwW39/jeiUFe65yLeOg+JoIt8KhO7PXi31oyLmB69wOXxS
iQko/Rc4WtUsU0Z2Ak+93MQacc0esOPmobkwB7gobCdIperUHT21+x0y/lwltR2pN2zQhNDN6ng6
E0samsHeWBqWyQQZP9EonSPrURBrp2mD1/7CYq2D+TCAjQ1IWy6w5Ji/L0FJdQDcGMtbo/UFzY+l
cCrqlZfbZ1GkCQ1G5gJIyiEi47SUfLAFqizIuQXkayKlVCQerttivsIemUilgiD7andd2AwfaVak
EYSxkfQg6Ypkd2X5sKS48UMaK9Ef45sggHCB99Wj4uvW4Vif37ULDa6eSu3ulvTRTAFkvo0QwikB
c1Cmhvmeuk/xF6zhfIt/A1Hz9jLt/thfk2fAnVNf2sfCWrrhs7yqtajnVT52918yw1wwEG2lXZmG
osBGdmKd2M5pdULBYebv3SERsQ+IuHgZhlMA0+bGK0KU7jgBJh4LpvvuNc5ZXtTSvio5b1nZE7zY
V5a1LdkmLKGv5bS2W9nvmOgmA8Rw25pImD4of+jHfvVZvji6gK5Kg1oOOnhnJ2mDX4XH9Yu2mTvI
ta+EMWxD8A/PzjLJ5VDzRLM2oRhUzwXc7LeFzbEGe4YZY4RT7zBIkz7ncId4qphIQ5oTaCze06Yu
Whc2LJ6sQ4c06uJES5QRM1JRJyJl7fdSrI8E7nYuKUCfnt3KR/2V0kKnNnjxSqw0Z2ES4fM706y+
Eb8hI3Nxf7S2/BoUsipI+g0q1Y3piLtFkAsVHTZCRnSpUk7dKSD0QVZX3RDPiyX2Eh6Q55fbx4Np
aJmYESyL2fQGWjGML4nmalPC2TTgqD0IRCzbQZp/Dauazd4xRLQfZOtbYLKVoz3tOJuPCFiYe6WY
hvTI/oe9NE3aE3Co4bp34Aml6yPWRbgOJioyTOMh9gzreHoHOm/XXmxDUM0uKl8Z703OmkpuM1MM
ycjymbBxtp9cwdUlKWCuNOPvpv8b6YIcQlM8jQbyPk7w6rOXgRBHNrnDEok7kazSnPciAxo5arzr
usqQGFmDqEwT5Vd70Ns2X3VdWyehUliFu7EKxWlooSvPtVth/7RzN67cfYoJhuSMhydGPh5OSrc7
DX6wyP29bMV2TJ+FmI5suf2AyNtwV/rVBmFikW+N/ta8Xl/PAlp3nN54PqbuHmm5k+ps7FV7ZiJ0
CT6wrLufsHarp/b52MrSXKtrF8b7SuvzklA+CT78JP2lH8igjx1nKe0C0/ymT3NRZG3REy2ChcOF
oz4TRiqjbyM2460QyewhjcD/WZjJAE+TOZrLTVplNE/qaUDd/T7OUUBlX7qAGV+UexFyrsxN6kSQ
b1AWnbEwFF6SgV/zsEGBdCgS6Is/9lUjLSdSRZzb6x9glUdVOROfhOtjtRa/0W4lvE3d0PXp2BvT
pgClmA0xQd190Hb1f0NcKfq5/Up79kFGbLQY7z/ujH1VarqJ8wnFiTCSpA28cefDf+p3MWH4Zc+H
UDrLTT4qsBmMzdVykOlxCi/Buv5giWOT8ezu/5Ea4DWA2YqT0PmmuOngltSmec/tHD0KP6L7IrGv
2n5KJOwqsgB9ctS7Ax+HJ9Wb/gDfE/WghwQdBOluZKxB1x+5aMznEsXqmbMuqb+7cKDwNEq5Kchu
uG3QS68sbPNAykdf2UctnoueUSibSgEuY65a7YDM2lSUAllQWRx0xhcHdVgUp+o+WhP2Bl+i1bE7
qZ3+nNumUjML9EZ5ZOreIKreuXbYczumocQUP6owpNXudQzCdkFQY+12HW4keNP0pZuPnh5lnoDv
oOYWm4dWthfDSw88SwqIy4WljODMW+9FpX2gTWcFSWGxWg19mPwY+rrXDUe5IrFxHOOhJ3pJk42Y
wBph6OiU2Mg7AiROPkgOAud9CEvTQwG4R7hHLBA6vVHaILZ+oBBZRcMo48nAt8+bzg9hA1w3tjLb
oLq+ojFmkIIMWLRoiQ7VfZ0ourSt1HwrgVNmHVLXoGBZAXJYQHDW+M0dvdls93F25fVAC6iPkgeO
Ew7KAcIwZu9uOCSDMd/CNN5gzFifAo3OsG8VL5Gq952pP3GbyKcsTMHA5gMC7VLvKm88ijWoJk27
unbAiKo/AJxmM0o81lcn5K1xRb5JRu4aAt9sJYOgK3ctJppNNALfiNkQ83sjnm2tFOSLwvCKrqB0
F04cAznA97r3vk3Mhy0gzx5LH9e7lDoIeTNHJB/K2jGCaHBKMdkqO/Ckx12GeJxpe/zmpk7qEgxT
HFwG/oMuUhmsLsH49lIxUu/MgxzhH2SCjPo4/XpjJkbgXnUrUANCiReevXTp77v/9vr05PlWC/tN
VAd9Hn5Q/+eaRh4X0j+Xvw7phVeyy+teQe1INtJiOwvVvijdpYqct7ZwjNwOD8ArrxcFoHkJhVeL
3uipq6zlGDQbTVYFJHKfNPP+VUnXmyNKAEZOqTqJc5mAdg12QPZGYHTC0EoRn4hxTO4CUViyU+In
JYT5/IEi6RRmHTWZy+nOk+2/VlF0FKCVFFmAFOGKJtQlQ7+wEKRPiWjCg9z6KFE3SNgu05dwR21x
qASy900xYZ/K2fZ8FncJ/G0hlbkKziZEsSfHceLgZqZfkjifORvihmKJ1jxvVBN20hAdhPHcQNvX
qlnMBgGltrDz32DL2czlwDWZdJ8KEsuR7Nok+ZEJpjhDcds6MOanLHh+qVwWH6RcD5OKO9htazlo
tch1ApmSEFHTSxh1nQdDz/Em55+RwfcN85rPD5BVXvFKlBGmcNq7HJNHyE7YujvswYorh96XQDN+
ijhjE/iT479bx83TdYzS0OVhQGAHQ8dMhiqhQRYWjhw6TuO1PVrtEQd7gWW0NtYJTvjwMjLuytNV
G62pE0VhS1h9FUuNOQRcg7PuoKXDHuZnLXl7MuMwSQ9hIsfhBhXw+dYXPH6LZSYRpYFBvXsKawr+
0SnTkJfbBHB+iAr63XN+w6qzg3Yp7yGWBemcc1DIkT3+UMVq3FWcqGC0evrKgN3jdSNn6v/M8ml1
QzeAW61lzbQnNyBSCg//XH1Q15wFPBQMejQkFamP3qDpYmxAPIm+NBA9FdP4B5QjmGv9zJWfMCHE
izg6g+ytn0ov7ivW3JDF2CRdPhhKRiZwyyMhGh9HkjuRGDjufRQs4x7wGbxLNnHwng4dxwxHKk18
/VMmpmVA1p+qvVnrbsjqUOXwqHmYe0GLq18LyY2hMrcuBaNSQsU9Vm3FwASzYHM0V5p2E1bdE3pY
Q7CW2d6gisi2W3j4fwnQ06Tw9pBr7ZeAvQNx9NCN86ohAzSG107ZNo50TuUu5YY+9X88nPtOyEeO
Dvuhw4w78863Vtd4UoYB2YNNtvTWKsENDR5wijGyCLEUBQvLtXi74GBLPOKZSb2VuSFpCZBJXW67
k3irjXYGoOQnhzNPVtZOYZFd5eBzEZSyVylBTn3DxkN1tKlAtS/5+BYLdo7FTJQ8pYArW6AQoA6w
HoFInxA8S+81DnK5BHX0p5Q55zvaU08/3my8zdRZ7g8hi4jdB9m8UzTrQVDdjeSs8tRI6UHRs4eY
eLZpdpHVNyKw/BANifmZnMnJuodZ/8y3FNW2PkhU1J+BSPXEY0hBD8xCcKIDk5SmiGbwO17BKcOv
YKkHqQkh7w6v2+aFCqDbsTGB0VE1cwBeKpXFnj7emkznEgcVCM1myeuhVaWoKoRnxvEI92x861u/
tQFe6CIGae9yqdPv1FRpKbKZChgfXqFs68jBR/2zMAcET1SbCM1Le/+dEsng4AKAs6NC8s+9XNwH
0zUqmaPax/5Tp2tzX46ro5QGRYm1ux2Td0BbM98sQO2ooA5iKYX1ReEDRKRkTSP31i9oDVqMBHpj
UOBV3cpeAriZg9C35Ze6yW55onfug0T93NWfMRjs4zI1LbmoTv84t18m69XeArUaznpDVtaU6xRZ
76hxvihonOoZ1x9tYRJ6JBMzrARkVjsiVt9Z6qR3Or0KOUQXExd6zwHBMXJEKXBnJbA7lXRm+YNO
sfhpJIIWnI5ORgcGz2QRD6SYx77SmDf9nq36gMfmL0bEqIlnINx0N3Vjgr+ZrNyCM4C5v14W3fha
o9YgB90xYr0EP89unRQPhTSgSQXjMSeLlzPNK38BqrRDj0st19vM637E2iTQIVVuZWoQk0UB8sCq
QvzS3JjyoS7/kuahgH2F+JEFamoZzzrv5TcvMBr5Sjwz50LirxDJc30vHDzTKL7Am/RITe7W/lZ7
Go8TB8oBYRcJ9AlGfmbqsEJnf5n5oFZW1H5AWgWuqz1LS64hLsVCWFqK2EWpFwIpEzP2uXfsyJaJ
tCPZ6kKU6/+CndA9I9IruqsoB1uvqo4PGc771sTviN22xePPuuKIcoOki1GW77yqGkcFOw5H+yVV
V0V+CtBeG52e66A8mb2NleWF4lnQEjgRf3QhKlm0t0LVL8I4Lp/GJiLgVKn9fsqO3KW/x3quUWby
8DofjcSlz5fMdah2uWKZxnb+B/Bk87SSJJ9a5ODdexPi9orS5Apfq+lOuknuz/YPgD1bU+ReUicf
UXj1UgXNzD9SydkAAgFP9mdN77O7P8Dof3tO1qw/BiYBAlzs7CLd3R6+zWfC7kFOZwuKRHe6Pd+i
wx1YEB44md4QTm2KGtKkFUg7DBc66F4NDzjzkJSzCBRMSRewZKiWtxv3Z015A9oV9Vsl6Ka6Rc/O
KAKe9x/MVGXDGup45XK5k4V076rSC1n/mSKN0BkT6eMs1XtwX1glHHdFTAUGSDTfA6/E5DGLig65
IhuI55Z9qKhCBzBbwcItMwRQTumnlB51djyHkCzh4F1ehhaizrTLgae/oz0dkgQ8c+t16gb+D/Wi
dTB6EVl4C4n6MsFcc9CZhKxiQNSKVo8fp5Y26Ucz9XvujEpwXGv2qqWNp2m/3cN55yShbSdSBEDm
Dvnd+7FqCYRrsbUgRYmsWI27j7uxBgHsbpIp4/yjaOcc/aVy2oQTo8sijW7Pj7NExwXE8TN/78xZ
E44ncCTtLKMJJzNoK7ase1JtgqS3SIQ0dCnSumhsRU23DQQf73Yv9WPmu/iY+KHy2T9mK+Dgg1Gk
CCD5rLDZJ16L4ujVglwcn8spwCG3NYUS7rJkC7qM1aUR/5noQQNFXaZVhGog0Ugw1puomW2jVu1w
5SM+BW8XE9vn34Q9L6X+MovMP5hRbl/4RueoJ+Xa4pL1Iv6fjZRVfW4Y8UTM9+JTCYihOcnzWG7Z
Z+8MDKDMiMWl7WjpKM0tu7QRQ1cOA55aKnpSmzYowbJXdz8DHHQ5ap/UO4uk6anrm2hnLvpBx/w+
K1F5DUMpdB+2y4TWwey62D/pKfjAZP0jxnsOXWhRb+JLlFi4kBxMV0+Lea0B+4cnj5HdnMT6fkD8
v4AP9rrMKWXbrb0DRmJZpc2j9guejKoBHZCcdySXsLIheVnNwcFO4ShUCcgLg3JycAp5kiUPZABd
c3U+yZ/px/wqgHfsjcox6+uXE9mNgg0ee7a5t1tFDbpWpZn3VG9z0/k90opcfRdf5qYZGSSbSHpQ
/OeV2OkCKvIlke5qZZAibm3iBhu/5TIvJcUHuVGGIZQ0jV2AE3XWasYC5rN63mDvnCzQ/twHJHJn
G/kiuf3fpnf6tOUfbRs8n68kQrqOc6/8yWvN8CT22rR0guI9zBrw1y66EJ443VtkB33pnjWuvdEc
POScM8BfS6USw8TOYj8l04hOA2DjitRBmzNzhhVM16XFDrOfUAYa8knjuB+i0aUR5cAhuK6JxalJ
N8ufVImFlg0yHRT7a5f/v7UKut5Ped+dMe1Ajz62KgatmQK5G93EXCzEzwytxqFxD+nS+AXJTPXe
lQ2hog/30xAVXXmMMLT5avYrtIaZJ7+p8ML1Yh0vsd+zEOY7S6aOUQCSPFBsiyxXGyAFBAmfydUx
fiiCM9aEoLn3zh0BIzH7vCWe8vgB+Ihjt7IsJRyfnXQXaOnP+tSc9/wAddN0Fz72HvTaC7rN2QSd
qfeQHox+LPTQz9PRZcUsGq58+UdKzNzP5K2OgqDf1+nLZpLNmUTx1fv+CPXNlnSeQezHcJKCSGKB
EhuyX64+iK45zMl5ls2KpUSCTHLs+CGC1FdSYssW4DYl42xtQX2T57T6qKHgVfBTHHb3KYkvh0Ze
P6RRGIyps1GvnNmegSQ0APuKZLQ6YU76VIBQywpAhgcvpsw0ixzc2KSH68TIlJGWB7k2+vxtqTiD
9jcF+sjq/kRxlDZsS3y5pIbppJC0cZux1fDyTXu1K9/CGzPtsVhOIRDo/BgX6SIsOxINR1hKtkcK
2RE+Tvpfkt7alNSuGxhhFT6bslBADJla5RhxK3Q4KRD8wOLWOdT0LgIJNwdnBqzjyTeBlr3MBLoK
NThix1i8OcflaGdfFO7DdUvvVD6ebjsfn6ZlPkL4JWQyeDaZd8smh9BuLCQOwu8pc71mIQuI5jqN
1lT6mxeN5CDhvSDuluuNx+pxDQHjYaTX+gynuzNz41WGl1vVeVHrjbqJAnwCyl3MeNSujpxLRa+u
lSYbl4TP9vGsj/elGMaBUsVxfPtGnUQPr1VAaUUxNSSGFWFkFFbEcW+6Jkcy3ENVUhAcHhTI7+W9
dfWBrfrMqwp2ISUMv7+Cpt3z+pHh5MxgAZQuPEi5D5WeuA6rds2eJcZQSb6mEvF5rsjQT5DvyCZD
fTbsJnhAq5tqZU0UW0UP7msNYLsKmsS/Dz06/isd1u7+Mu3ERiPitDddq7/oIBixcwkaKlKUUEjz
Cyt73B7E/fg9NpMzkv4NdFLaGoEqEZFZWp0C6RSuN3fGvPFhP87uw7hgLKWHg+C1RS8f5gGN5Qtp
LooL5zG+Lls4TsybKxdUZn73QalUNGfBdDX2eH4k4RMZpFbp7o7NF9qaxrxUFoV3pVZizENbwVIm
DE6iHZ4wGLx6mAdM68vLRFdWvNlQbFrr5BvL6Tptc1HbLCkFWbwij+oMV0DayaD8cWVX7LiRM/F/
picuqqXxPHv3ubv9OdkSSsulzHwvPvOZDvSnjWBQWZtQ//bfvYoQs+UBj2f4nznWDd3mfGjdmO3g
oEiraRIwIxFfaSzvIfNmzmYSbHfzTe8DZv7vNzPGqp5SryDeM5aJWx6E/UtKrZiL9CTUrTZk+hvE
GUjRrS+KwnXB/Uknvnh8neCNBnqTiMzSrCTFcGQvkfpGP6F/L0qb7Wdejz7QbTYGMIEjFRgIIpC3
vW/oJ/X60y0if2on/J0kV1sLaiJD2uQLALK9kQWH239ZAcg8GmZUHh90KMa3y4/QU05fc6EPrnKz
rM8O20qLTWa3Qm5A45c9pvWvS5Wv4BRE/rdyooCvD62lLOXMqH5nN3zvlaumLPVVVvpanrsz4ZGt
jg3MP8UjUYsIsuVu+4WKh+4g+Fh7z6IEjW5WFkpr0iYwxIqTTeCdHwJaaliTDapBpJ8QHA7U6SyB
jVDLRcmvWaltHGl3B6EhBj0Ccbz6U1bfGi5eCsw4UpMHxWfeYLnU/XdU2yKPMCBTGF2bTayLH5ex
c9CTP1I1ROU9I4EOtyC90TsrTuSLPamX/L7VVBIG7U6+CU47f67H3Hw12wMEC3D89MgiwXbSetWi
zoyz4Q9b003fi8mkrh1mQ7UFWZWxfkh+IUu+foSr3K1y9X0HOCudhqx+B8OWLDEfBfGrLBRLt0Hc
jxeqZO/Ot6z76x/Oe4BPU42/KX/lOKGcUMhcJvjcl5oovoGT8AlHC+Qs0e0VrPoUeeH1HZw8ijgQ
7YmnqteNPfmZilYLxEiuJYezYNqZ9CN81g1X9HKWWEFdwq0YuZKd6lT3JXKlJ2qcxxiUeB2vheun
YbJpwyaCcRcuAjISz1Qqag4LDKgE0KQqcTEltWI1OQwSBgffhHq7NMygVwz15PpgHOz8sLX4Ek2L
lTXLnwsnplXIuv2jppqa4KlTWsdsKC85cLHYBky2QBbobnM2xdHEj2QeHG8p6ZhdH8xU2kMJ1A99
D/AHjJC2CKX5cv4YJk2KTlBHuXXSmpsBdKPNrknB0i/6h43g38gAft9XdV8I2PQ8J9p36hGPzs0G
S4qcKv9/2B7Y1F01bV5CQ83zpGmZBMfjzUqNku90Qq02vm2xwpDd6oew40KbHPq+g0m9ur6AbktW
OlCOrjXz3d9FTA+oJFn8iZBX0Um1Xwa47IjLLBAO3xh/mQrkmC0WU74bTW0S2LaRkufWPeIbnSeq
vm1BTopwTrUgfrAtnDzlJJ6p62sLWvgYGqMwpMfwL34c5YzcezyW5DrGJvWYLysc1tjJRa0hI7tO
IEkrpx8DRf6cdZ9FLE0O2+uWoGbSnhqoiKfErzOKDM6DGhD3ei1v2T/nen6152fvfWHZ8y/EB9r4
y9EjV1tMLMXuBfYZcnwjAZyaKD6pcyqStMEyX9x5f6WkcbGdZ08cCpAR8V+gIMOd+Oo1ZatdycDl
HJ0BjVXiv1CbWAEdMDwHsLiWeFYXNULFlRyZhqJ+0mEF1L8PuTfvFUPbrnL1Lw/+c5Lg08rDjVEq
FLsxYr2zPMN6vr3QxIdyV32FWJfCKCJOdFEpe/EEHKYDWiuvU41GB6PttlVMyL4WRTre2em1AW7m
OJ/RD0oOyrhnb1+TgRonKngx6bSmBhDmB+OI077PdoDbVB7qZw1dWLgRugSOpDwus1LGAcg4nDui
9UDdnZPe7NNjkf7MAGk19FPgeUc6BqG8klLpG27bhpKyLUCoNq8oop9Tat2QBCsOweUyPBjHyL17
5WWBAML8zzUiymXR4PrZ+cP0mdG5GzmcRbkj8+PEpmoxt+4iRmWDVL1ZziLacglck6o4O8NE1Ttz
cx9SyfDym5mARzvNKwJXGFfqneM06HejiHlwqru0Pl4azlFUijAga/wm9JsI/O4lzL9qqxnTdfX3
/uIdLjizLc8wJL821LzQ9pEnt5Az4EW72GqsjSAUmuQnrzShPCuzCK14N/hdeXjSBOoth3K5KPcI
CKt3amCgZdhXJaNUeIA95So1qyZkyA0zMvLtAxVODlItUdj7DsQnLuH1FYGsMe2V6E0y6ZyH2D+k
mnoezXhERhqP4Xkv+xL/MRkWwZ3beO5BsubjVRESt5IJdCOUubUv49WQYwPaZBevuBemXyOAIIgZ
Kk9gS8rmlUnP5bXFDVtzIbChg2fMc3UxEk/c0qivVNYWBKenwUCCAqpca/O6FKjsSRAItcbJBkrg
DiZ9rN6GgckUVAmEHQtTP5jcTXq3PiSYCTQNwghmWQJiKIL1nVMGhyouP0U1qQdkCxjLnbb3nRq/
Q0R6jB3x29fk43f2WYTSNC4nT1VNiSegTVwVGooqT4aLMdhDDApCTTtlLuOPpOUWkriVcM9PrLkp
5Xyw+3kZt6Duze5p7Qh7dJpv/gFsgOPthrv3EV4G9xrgiyDrmjMuoexBTjBdyXVmNLyVigjhbd9B
u77uVm8qdkmy3xt8qHUb4JbUtX9A8D7oxNnRlFem+pRVkpce7OEB3Oz9GfvQPcyKEpHTCnXNPjFa
XPPCorh9A0UnDxCjAhz4juIvGvVTR/36ajRQtB1ginwzUtWRJRGy+7uoOaNv2OzyzEp5e9QEgtZa
s39+hUpxNIjyhNJuJ4vKvjANrhpACrb7v54TCT+hw5pcppx/eeU25Rn22LEj2/KeQvgv7/R7WoOo
GPhnydrMdEzM37vWRHRgUKM5m/k+NxbUNoF7nX5MVmYL+L/C2UFFoZlW7xl5VpXa6s6r0dcK9zrR
Stp8TvA3WX/s5TAOQCt26nxBY8tcHupxj6skO0E+mDf702xTVNpKq1nSngT7UPGllzzVPNDrwsA7
ex0UA8G+2u9V8e3Gm4FOxBj2aDGeemR51ZGkB3GBd2m9dqf4f25iALOLHhMUacpLAs/ZxWFHEXXM
ianSbYFap1UHOW4ryx/4cxAJuBiampiir651X4Wo3DCzamG8kqivXOja2SWSzqZPD3+If/W4J2pR
gXnvF1fs12t2bk97z/T4mneYvSGMZCfDYhXRLUkq57v9jrLBU7rKnpycSfg2GLhQB/ABFfVSBHLP
O3A5S0p5W3K11woMglddbRaitMWrSao7S3eajdqFAWGNNvxHWU4UDZynRqREaCfXr1Ietuvqypzy
cZ8DsX3iTKmeGCZ6a7BXidIwvOUJ0WDbjn4NNxh714BqBvQ/bX9rlcbOK9ldSimuS+saJV2DnyZG
GJgerUp9QyrRLTB/ODiIu9DWKjjb6CiFS2ijG03S8aSMf3sCuHZWfYy+xZnZH7JyeWbLed1kMQsz
a419LT5hFOk0KFUSK5h2oO4D5Y7JTPMvuA+jeN9OXns4HWdJe8Hj92Kn+79RbQCo3rEjrwSL3o14
jrzrFpfZzZoTDiQuPMf0iuW3m1nx+mwWofZZ5uHIEPt5prHPpvMnJFgSsC5ABfLQAfj77kD/hDQl
6cRR3JcU5lHWcEOYxiv91IBe/2auS8mXS4Qz7YCGjWPj+/oezsyp/GE/+8DD2oVr4qX45c+jo3/s
A9E8iLwuOjiBmHcUus9FP3kecDj2URM1MO9ihVK/wiTpQwzYrj4vnploDf99ye3YYUyrphYhQM45
n815q4pA/yboQ/myuoJHbOHN31qdAB+yj7KKMWbMqhRuHaorIBCG13Kc9Mvcf4ukfuzrhSRbsy0j
Y/MYENRyHLLzJJwOpH71FVNJ/T8EGaXXBaD85Of0++43L0SyrvNu5Csy6lg5gpe/8lU3nTO+7T3P
6t8PMaJ0YC2412VKR4MXuzmeyDDLbvSE8hoDE345rTD9puayv5yHUyrErQGfeo7PVObXKe/7vkgh
ToG0gg6ZfC4frxneB0NHLsxnh+mGX1Jj887kFjKuxep6P+RkUQFC/CzDUYpl6QWOdzGwZqWfNZUq
bNQmnFncIhlLN8Jfo38HHbSrcF4l/3NgFRe+wLsEq6t9UDv5v9AtFV2nYY1B3BD5cJxdlH/rUgMB
Sd2X1f32akI5jXAZ7N7RpDvggI/ejBJL4Z1jUbdopCZpvkWvXnAWdW+0dAXpYysd0SBvZP+j8pUz
xncz51cfGHbLp0Zz8ILuzloaRHSwWoXyF5KThleheoCHF7KA+6Xf+nogwXycfUrCMapxy+EyH646
OjsMooIYHi8KI2esjb/+9Yf0C2he0tKgqht3WHJNUnvY2gUC/aDLq1uyKK0PkU4zfyS9zZSkyfZ4
y64kMKN41EcXzOpV/L5eIu0844wg9Yhx4/gdgk8aDIV/bl1cJy1bHOyJXDzMScpSTFHC8n96kMif
SKimWVu0XlTiC6YvUHOBR7dKAH10utw0ltRpH1px7EJjMEPOgiG04L/l4B07qmnTljW96tw8W1BG
PTELqVxRBRFkEC6UunWKinztlRBAqqba/o1ym5QBn70HM2dLXVrInMPZ4j1zKX3xcuQmxSyLOSpd
/ptZ7YJLLr3eC5lPjOJPXtxMdeT4Ndas8J/M75ajYZFtqxiz5l9XKUWdnVzk/ftenruJqA4M/Ou1
IyP1E4XJOC1tSH62pjLomvBxy93ssHlFNEsUrwN2M1JSXqYzSU5iO3jumeUsrolTOpSyJ9L60BcA
5InysxPNJ0cuwtKOhpoIxWBi8Qaq3qqgnhhlFz0T49HnKN1DMuA2Ox54QdKQxIlrdqfLZ+69w2KK
QRSsx9N18NVILXsf25Ip9hpcOrbVIBcyKNOhPdJX3WF6oFXK5vKr5ubTYo/cyOGByt9/ccVd+pTX
1812amZZZeLw5mCwA+tx5r7FUL0EsQC0EFROk3vKcWH/Kf5REYD8JJKnRY6HatC5+CBGu1ICn3Xh
V7cSkRP/nl66kD4dwYVURsDBqwCdE1N7ToH7FPsGQLIKkP+tFGUPY6Khn0xUwk7YVKTKXB1uZ2zd
Tm8pPfsEdsTkTPrl1q5SqX2D8ecaKx4QfdcYribOuKVIZDfeHYZXt5NpsfY7g73vj8J8Sllj3E+S
nyWHyKjatOMn0Z1mYznICQkxiImHL89dAtAnEdZsfCh3YsM6PsMCPjnn2cVjRhg6+ZiyaoFa2B90
YmE4JrtA8LVCd7uw8VjtJi+YK0Tlhga9XdElzhXYVJCy9I4c3zhbu0Sty2rFG/Rpq1tVwiD7tyu2
H79nSrKGVhAKPIpjq9mw4LwF0/9h8oZMPZ1DkPePX1iixqYHBHoZnOKAlXYEgmBh+FyT2ZRaLb0h
KH+S2/hb0wUgcXXjcj+sKvaRjhr8DRhDNKAKFobdxyFcFKDr8bM+XCn8T/A97ArtsZeEUyQWsjPP
WdT+rKb7IPvxZlliggpfpETwLkRaq6fN9hyurH9W9h00r8q5BhqOO2Qak2tqhcU59FeU9zgaw3OD
2GiNY2R6NcOVk2p3XHJZj5Ki4NEfjdJrQUtDSQwQ0QdJ56iDJTx6gPqNW4Z45s4Bso97d96wBmph
zRjFMJzKXhH8j95PzfBBMc+aKCmYaFkfj0gVcGlp3AsPO0NzzXqePpZlKbbtwAyLz8c2N6gb+qwa
yuNNES/hWsAYl+GG+hcQQ+Jkkmh5gdE4JGLwPSLdz+NV3Em31saa//KxMplWlHhPtwnb2auMJDES
yJ8jSvdOo8jPKJ+IjprTR9858uhNKu156uWYtd8aRF+x/6C28f1CXYYt9mXlBFCRdYKGxD1W4wEH
SEX2pSDuXTUPc9rZ/rA+TSBEGmPiFNBQaif6y6f2lTyfaXWCnv4+EIVopnx9XhL5bHLi5M62EvwY
L0lFnxrJo155nFfG/4+w20rvVP5oy9ovNLfQ0QkVZuluKXwyS1JhzXyMhBDXzJzkFJJ7lp2zMwue
GFK+jp8NlfAdagZch6Ec+3/gxoMDweS56fEorSamnOJzT6BJhvL9+7g5SP04HJ6b79R+WndGaM2n
k42a30eifc85Ju7gJ6BFlyrge5bf//UoTGieAoSKsz3apO76oqd4PluH6pBAe85mwRvBYPsOonpo
EEDrzxs28amV6rxX9IOqhP3Ehee3aU6ILprCRP2AR3s9pK88E2E64zlunDOK4SptZUrfeRVmjnYD
vf2sKmYba/fKVLuqPPbUE+l9jUsqx5tLNRK2TK3JMb5awQauNnHMDM5OU6gG7qEKKeRXZFlKi4uL
5dCFIBLvs/JSJlnEGNC/z3JCJ/16RTTrL59267f05IC5rS5Jlh+NF7p5b48YIvbrjzGxyDt70+h4
rh/iFZs4r5aBhPrD8AmqI4l15IACnN/uEbhW13DvRV0oxbS6ROw3Jj4hCBk7vdoS0oipjDXM3WGo
fDsuFrIelJ8q2gHQwCBVHCpXUHxhRQkDfXez+ldxYumOwUlU/m9EnOt0ZuIXZDxrqNYskJDBI00a
D+kFHnF0s4fpcryJm7EPrbAQ1RVmMH8JybmvTSdt36zA4V0s35UjrSr5XSyAEPZMrCJS0mp/kbe+
wG57Y9dG1goK9PLPu3+SZfcoVA4mjLQXtK0OVV9WEv2ew6lbJHM+8wfHxavMBUTzOnqGsMeesd68
c1JO4pllU0yAiss8043idSwXsKad/2P8j13E29BLDVw00C4ll/zt27SgQIxg2FBbEHQ6DlD3RhXc
NZ64c07uOGY74IQxIbMEyuMaT+M1SsiTHkuZQaQrL6ODWBhC6VmroWwiiG7i1fX3Nvb807KLQCe/
DKMWpMnqJx7T7HQRsaWe2gl9GqxZOCDEWib6HPpDI8zTFP103katUXcVZ7LAzh0ZFOLCWlR1Pg9A
LdBtGd1MYRRLVp8E4iPonrEM1H8xamJVSDe4MV9fUtsNQsT9x8gdJEZhDAsHhJDHVTzYEFYgyPBQ
Sj50VPVJiPfDO+JTZSzvsYTplEUsy0LjhKYdxkxM0gZ1/CkI6m69HI28ncJI7DYu22lBJHg+gpg7
DObtz/KR44z4pj97DZPgVsfi784BsNmQKrVVVVBdFfg5nzc+JQ2yBLojJGhEGrCzNe+jS4qd8/Gc
Xr6uw2/5QlG4D8tjuFfJKj9xnDnKrIm/IRw8NrXwGc8ZTEEcFqKLD9SouZSntiVcr066bDKrZm7X
5pgLc4jcT2pYTkpK+sJ2l+jFENxWjQpfit7iaBaWJvFr7eDkTQSuLT9vSIMAIXVro31jlSgjzA1G
3Y5pzQJupcY1zJ7rvmieeDiKI9Qs1TT0rnIOdnVsXMiTCcsB0JSXF5zXc7TMDxohAyPsSI0WWuRi
t7pBVuQYl44hGUbdP0MEikISVuaDFmZkl0FkXJHDakLf04v80hYVU/6g83SHkW28/76F9l29kJ67
fZsEjyoHa7mpuaaVx/ObcFNvzD6L1zD8Z5NG2Yw8W+b9u03B6tZwvryVR37j4e4ONm4azT0tUROz
6QkucFYEmfHFYBRVMnJQ5+5harxzMWY6f1Zs0KYBhwM8v0iZ9SUDGJs9QaSy2Rnrxe1xmdPvfvRs
jZW45TMfoBDmy0JgwIkCdafv4s56cVLDB2aIhnL2VsSbE8X2uCKdhE3K05hLIp3vItEPWwF5id5q
tUMcz+9u8EXeIl1IJG0B65qrA4KpCtqwwYAWiw4ZqKF47r1FcXvnClpGbw3TzxefBpemBTN8sWyF
kBdh+UsUxbG6UFGmL/YRKMwg6RRKsIguejpZcU8d+EmcWv/CE5KOZlB7Hjw/mLl0773yiY4AM2OI
cIQAOnLCxCejgpuRHbsSLg9GOVBRTv9U2x9rdQ+diFv59nPbxMuy9aoNobJxW4UiyaVb6KKYp029
cMQoCXvCoYj87LoCpwZbwwRPKkxLAHnpZyFBRWcDLLLI429p8d9rJGU1txhyReWtGxGXsZ4/8nBA
+90GYHZqzTh6ELouAJunYMCzDzcFpKM49JkcIHUBSiRHs4Y+2bwz8M8tO2YAlmzuTn2wa/iz0q6d
IKxntlmqNSpbVZ1DoUMKVRaXi0Pzq6SZbTIF6B5IoZxb3OYXbeJSoBaaYOwPAlYBEYCPL/857iE4
ttBl0T2K/2ODpK40FnBSZ7hGM4vSNgF8z59+g1Wgs++WtDIBH6P2HlA7FCtKLKrPVbpitevNRMCq
X7sHRTFB/bmtt/nJk9Ey+VRf2X5tbeh7eVPAKA1dAmHZ9FwwCx9nhtysTfb0aGOK/3oPmnhtgVvE
vj5tb30/FuBWme3lahS+BuCYw3VsLULvU3hL10QQKYcmRmxDaHeN4Oe8dZMkdcaW/3SD3T1tWFcl
HMjcEQErLzNo1OsQ+LzWX2DkR3XKb1Lk6pGoRttyghKrcmjDd1q5Q449pdb7NhXWnVe5k/+THKrl
2sJoV+A2dSsQbr/FAFkD76GRF8QwGvA/TWVmW+t65Ofg15xju7Z0ok5uLn+pBXidNxzCWB08kd8P
qdfH056upE5RWWc8KqzRcBRDj8esJeflmAZs/6f8Z7Jes8cDQsaVpG2wvGY2WTKFz9qh8ugylXOq
DOM43EZi7zAZ8qyr48UN6wPZA4JHSS+BCROmzKqtnEl0N5jSsLNeXbwijA4FGZtxMMusThbDyKrg
5QrcQ47cY6wx1mXc4Rkb9sH6rC2Oe0Rd9SfC3NbNUJ1WyiorMQYaUZSOqIBxd2VGRD0o7FMQ3l7z
S18CRHpGV7lx9Aw3GP7pPdBOh6WgzSyDERZXsfqkuxw+Y32bTA75V7bVpXntx3QZjdxIKTeE4Rie
d3oG4sKQg5FeOVmdgy/RbJDyddugtcIKejCxt0AeYgweNNihp10nyLpGgbtrlheuesXzltMtT23F
jc7rS4BrZO3p3VDeHk97sKrg46YOqmMxQKRjbNkEuEYeysj625f97Tl8dfLCxLsvGECQdrp0xzX5
W1nPSX4DMvuWOTZihdCKoFPE3qATir+Sdv93OdQ8nIW9kVr6wievRtMlj4ypbUtJ6XuoFY5Fj2hH
LwOrerThFs/2v+gpLhvswAl0xxZwxENMC8hS0/ue9JeHaCIr+MPhvuMparGZKJgUYFuv1qMRmo3/
B50DfM/sSB0HK/2EjgUtdHC2ieFRmiRIzJaEjHTDN6ho0F3zMCzUrozh0iEVqv87nIoQNz4u0dtg
hx5DN/IR2d9tdLiZt7ruFGVtWs/hkM/hBxAPP3Aecko9OAsmiglgg5Vlaam3wIokD2MFXnEI6qOF
pmzXT1E37hfO17pYSISe/5htVaGAJGdqY+/9yYXhvowDiiGpaK0oBslm+REKmGmV4rRwLmX65V1T
8uJ9PMsbLavo9DgdHvv4zg4yRzkXgw6JizMZHpQXxQv4MMa0WA3wxHIrC+Rbi38ECt8rGBng19xA
58yMq1FpOj4gnswvC3ARERgC6d2r7hH+G+n7XWeECrGppJT34WYpADhXb54/gfIWWCgbtvRUXqiS
a+TVWinxac5TnGDZryVoUogiW+ZOCCqXYPjnBRimFzFtUOgygDhLVfjTGg5WMZS6wGo9fVkIwoRi
0/JiqoH6SL2ht9NHyDTXdiExOy6AcQC1xego7xL79DIzUsvBGFgAA6ZleaD83ulnJ3S+cGtwlYEW
8tUlpjkfgFj8Mgedbp74v907HMCvsrxZEbmsKadDwk+YQ/D7+1VA3d58pWqukZcV7cUooF2LPJg/
QcXbRYdpA1U18sDqu30kUKTW/8qSIu1DyJjGTBBZxLFlU4ucRezijbeSp53g+CkziFri0PDPQtXW
u1z/ZcWXvIl2e/tijhuh4CVRWvClJGCnYGPYD54DrUGvnZPCI4bF500RlOWLm+ZP29iSTxYV6sJu
DfZscJ0wnOJC1s1dLPsZqHb9v8b69SZW+nxYlrGXKAxKiy93Ii6TqvT8uF2YJw/oGN7dYK9ZBGV/
Fov3ec9qs1+yDU8rauVVH+ejPsthI7lCuqluUk+AWkxHImYrqKiSJaHqBbyP3mQRixWfWtEN9Qwj
7sHZPVf4j/oHaVEuMJZ9CCX0rYo/1zUS+YWH3YtVZ97orePKTZKuliWL/fKcBIWS7w+MJjyHuuQE
GKZzYAsc4dWAqRPenSRJxgVT7/KwR7mO0qNz8AVAhgOcJUrkOXEn5i0O1VrhBZ8KS5ppi+rwqBQn
s16P5TPT+7EQTp81o+QeEkHD2YQVY80Yb9TALt371lX5O+iZ9ImYs1GEZV9Ta+IYmuwh24w0yxI3
TZq/0nGmr1g+J0MYZgvaCHxWY2dUl2YW02cK5WwEx7kGSjWDAy6px8rKsRcc4fxUZLMKhKm0TqPU
crQtfjUiHRbgitxx3dWpu7cuh6KYgMKJBiy+V7zKhX905LekEFZ6HPuISHrrUSC9fbKQEYOiYI33
BNhcvYFUANgE8J8IBYmOmOEdR1+corpfq8duj5cnMic6rferODGAv2HLOBajNqqAkEu39L0Okli2
B48My/PD5r8DBjiTZAe3Nf83C23RxlVDusskMDlEnlyYqGnHLUb+WNmVjTkba25ZMOQZbocOwH8V
9PR3GA1d8T5m1j+CKWTDE+005roBv9kB6o1qcwO+x93HhMzmSXjlAVB2W9VhnXEOev0jPX51aVqA
6Ni1k2ohaMUVZsLdBous0m8EEJSAsgoNbHErwoEMETBMg5Mnxkwl9gphzQ4N0WkSDYTh2GTN89uk
994k0RivZL9eOzDm2tVOkD0+OmSPPswn7/Q32SesUPYECNRIE306QZgHgZohOCxCumHNgaCbMv+4
TxzEpkg+7FZ1DMMP6jrh8xZZ0QXhdKsMpRXBugqtI5bwnJ8YYZEV8vfZUwco8LFMqgxItUkTWdfU
DjxzLvJtK7BwkaKbMu0kqX3xKGHZTQ3gw2+XkqZrHf5V89GaQowgordIahmhWrO8u39deMb+cG1T
6sn1c1YwxacKOQr7IbSwBjnrmdlF57o/M1Pkd9Fa8njvl0Z5jXX75rCjvTG77TRE1hef0P/NjQYy
YyqnyIJPUYxeJk9vfCaRgGECx4OI34e7Qla19Y6dr+YIyPh/n5o8IRl001ojgZkBV2TcioFjFR3h
UGJFlZAh+g6VhNBTRKUGaRS+tX0PNbTD+o+FX+lJtAuDHQD78k6oldHlQvm3LTkjhIQezF0NWsxB
lPBZpZTe+9DvwdevW1KFP/0NUXaznEkYJeIm9qYQfVL2Cqqmkv5bxsMqti8T+EJU3E+1DDxpVMML
2Cax1qZs9a2ub0TECQNedHpwi5/zbv6ZPHy86wKiQzIRAibi30GgsZn0Fi8ksQlrX1cs/PsMAFHX
lKgzVQLYR1lyIY6BGxL3m+HhXNQRg/K1DdQuCv0PM997w7PKVcq3OZDUdNLSOEakOGdHmkC08YGI
8QLcOrOutoaz1RJDF59mEFe5kUpDSqzWilynurGPHKSF0GHdhIrXHuRHWcxNIPBNCzeqoaMiYb7G
1vl5TCTGn9c2+G81UbO33xd+GZ98s1Pvf//pEmbYoi1hjo5EGEf1ZjCtrBCjSXo2VeQ9iRG+6yIZ
WRfG6O4bvPjeJg02llwdksLBLvxPy/dhR0OmeILhoM+3YlxP+dWxPalx1HIIRIt+3JPuKE7ocC0a
UDrDkLknzTT4pziwORbk69OUy2fEwjPV1DNIvF8TLhMa8osaeObVt0+rVNJjbZaQAb8P5H+Uc3iW
yF+Bhg4sqVq2xwScIye2h+NXyDyfTIW0A52ci6OdepkpH/KQXmwWs987IY1NCk3OEJUQA5MgtX9+
RzExEU5wMtLPXpfIwc2cxBK5rMikq591OENPhijvUoDl9+vw7leN3XDtVup1Xo99zsadXYXFLTsU
3Xg9CoxFze6W3yN4LbabclattIq4yEzDRpcODrUr0e9UO4rhoHMhWqU4Kf6C+fKrIhqf0hvRgPpo
5zhCIt5di/BrQBScE8elxY7RewQGIkhXnSlPyTmRaYIDDg4xzVjal6i2mDs9vIY7YKeK6XDznqf/
+7/Rb6adk9c0O7eF5vrGd12iASFRV03RkC0fM0Acmat045amaV+UJHcWMRPrhCOJtPbaZDxVi80H
TeOVYHSy1derf55OIj2cLcaMe8jNsV45nxoFVyraE9T/5nVf+jjlesyuBw2F8bD06VyMhKadlBKC
m/ZvqO59m5eumJeir0Z5ad6V2palU5sCP/MAfgYNWdzYsttYog6P8yt/hi0t+4FEOpVvd5/anrjc
pXnoUCgdmT8M0GZKci1yd73+Mq0+4WBCija/rQskk41oH6fDgl/9jESiaYJK3k3asqn85NX1pVo+
d56skX6HELfiy0o1KaWQb+FODQ6Ra5Mq7mAcmoAIT2lZOSzu3Czo9Kf4B2FFAHrz5sN3PLlkWCb2
yCfp2e0yDfESjkP/sFcNrz9cfreR0VUfpfI6GCt1iiXwL1WJuJ87L345tkGhjhpLNBIE0r58aY2J
BW7QEISA7WU2beFgRNRno97Et4+VYB2oKwS003toL18IfIXWs06I6VshaRCt/poA8pN10KILuQMw
Hg95MVlISdjQ8EF2W7ZxRfv2G4Zq13HB6Qkb6hYM6xNK03DZpCwSNgI46AlQTYZTnimvbBATVGIy
4mwXSxEwDtmayQNe155u3N6kv832i3Plj2e3WcY1le/II1s9Jk4aet7DS1wKMUehPNN3pEr6fyxW
sRth+h4PiviAi2vmPZ7uSSbLvMv8BYRvHvC+a+o4Ba795UGxYCVTPXghUkUB0YqBQ0aD9cqvdsP6
NuZZsZUlJSSoex63A8jPVG8H50XNzTpx3HmTfGqoio2L+nSmYfBM7vAIFQ7G8H77juaJUf+P5SH5
dJUqTBvCFW59/YS320hWgf3tgBi2L9xoOXGHTTeOxzKXdQZZUyENUKPAoA8qPiu4THptnELPaeqM
uwiHVC5z6Qk4pCccjnaJQYx3baaXlvbw6IqeqIy77aDHAXmlx35IssNxIOOiV42TglmDI1lXkjNh
uceEHnBU1Ngd8Vuexmi/46Fo7kPadEbJTp0hfHL65u3Y02KfV+odlOf2cph0Uq6U/zoNS0BQ/1DM
aklZdUdvbhnoSKrkneD7CGTnnjdFFI+g3Csjfnf1Bdw+A4w0/QSGXZpJfKbzUN8qpJX5f4NZ0K+0
Z2AxATYFxXbG9G3yUFfsnqNfdUxdhn88+RJkjB6fRb3IlMba0sQvIfuRyVtQVDifE+rmgl3R/hPI
dpmrFZrdrJUp4ejEJFDlurHe0KvkWNCxkGVEv9yfdqkXL9NkoBKnXviy51W7nG7ufUK2wkmK8jtc
R5oH8semnORXMmKne2bgr9/Js6OUUEyvCbylskhghIeN+GW8jPtgyOqHgbCLsONI4YiPOGdpmtMg
OPZmEc9bl0eb94K8muJPehqklRGB0Pq9ExMJaYbl92U/E1InsMZDpVm6n/sw0ArFjFqRwxGUf/IT
MAfjLGu8QgaYULg8PZq215GMxDwbaOkKWgIRh6pY7U4CXoYRV1T3Jp159vNi6v7TgfJmcZZPwcyT
bEbDlPDfXe019K55068Pn0an3Gpa+Po3fuhztcni2ewv1suPTP5Cin+bgyUoq2kPxlTO2qQ80R+H
SlZmdS7H/wrDAho7rll0zpiMLHwaFt8NMTXV0rb87mGPJqg4onK4lBhafoI3OXJ+nUWnwsz0e5EV
DbzoiBQfJvq1JIsroUmpAEUK8awePchuUcP7cLhewZA8R7NcPzppUzWvWknQ1NCGFQYXaCc1YscZ
mmKjMxBRCBbJDHovhSp3C6bSTgz2JtQj71hyzoJGNUyMRZiDQo3023uMz8LCDdWZx94J5aAomCW7
jxuzWUAQFfxkeoDfyIw1oEqmW43raJV8rZK5yQariDqrqAQaaFdVqmjhyb0vfnEX0rfYw3wDNBVZ
dUYTJbrzoU3MDgp6+UjVdHZMlU5p1k3llFjGodA/2cA2V9csr4AnZjUbHguv8RTScjOiLbucv8CZ
H3myJ4/zwxDQsVP7npJrb6eB96z2JfLxbbxqvIzvHkdE85KRFKO2VIiawf+yItBbGySGq8UOS6yr
fy+ulC0ELQMHEFar+fb/yDKo050PTvdtoFZbg52IZj56DkwcN7fH+IRmzQfCp7Fv/Wp748sAzwxi
KYQxeADQ0I6OenjPFngvfHaOAWVdr9oAig5EFiw6AfRAxC86Y2l4tx/bA+rNavRA21rixV9nQdGl
K96epr6ir9Ov3JrfsgmLg4wTbEyZ1//L3lv+DdZp4Bj9n2IplH2F9THDJTlnwGJ28pwZ285XNCHm
87C9hJ4omD4YYmPmoUNel3Un9XJoGQPqAybDzQBHnbF/HtQEg0EZzig0+FYDepCFE/aO0EtqcY5e
aegXISafr+wY91yz44WFbBWeT6zzEv3OQ7HQvuItq45SsR/c7K1/Se/63Wds86UvzSR/UnPqJl3F
NtcLbyj/mzoVvvjbri6IxUhKNGI8hz5b2ar3KtTujkYSE0pAeEdXuL+RQF+RWzXqcr61GKEp+lCN
IagFu3RJhxJtW4njOBqH5JniobgyTpNEKc3ByjbvD1JveiZU9+p55K1XUNctBoHTC+9wnYbdke/e
Yl0HoDiOxDnkdg3sDmhxR60ZSKBzOqkrXuzo4vYbnusxub9Lbl1T5c3xOSZnVI1CgGLMktyc3/bg
qcQiOiBw0jI59ZZ6nw1JA2u6WHK0/of3ZgCBnt8GLMlVHZkvuwmDuTx4w/cXb1DcotuW1Y0IygAl
Kl1iWtzJkdSy9dJ7EayPZVFEKoTM+F01euyoxWrS4B+mID81/GNl/rGdc5ceQHYe0gNrUruyZUzZ
4J1IKGBF+f35qTijdtDRg59M0Ph5UjDjSkt2CUYM17jY/xbChSWj0cWvjR1y6n+0gt+MjyoQbHPW
CCL4lJiyyW4B0V/rS8ahiKx3o7D5lqtGQaozcjkpS2xg4PwosOSIinTvIZoEWQO6vbW3PAF5bQzn
BQXY+8fbqDFf1TM345GirlEfubpmgCJWyST/fKRfHzUGlcO7g2asLJX3pyIBfdVQ51s0DI2qkytz
m0IHH4z6WXV/43NKRxnWx6Z8MGJ+ZhHNFZr46k8uGTWiamu8eFsHv52cE0NwztplrtaEKeUA2ZLM
O4o28NXc9fWdJTMpRy4Pvwfo4Ml8mpgVQ1Z/7YFH8atxPBT6wMYz5tKAMyObhwtnqmVJD1X+Npx4
4J7pbFHeiQkkS0qkxAH7AdJkOS32sJD3FJFe6i6ytgp7V0QThjnYdd0dQwTE+01gvOJryA/6KL4U
VjKszep9i3NNtCKYjdmMCsiju+tQk5NkyUgWoxwzsn2hyzOqqf0GD1xGhrBcxbDm5OY9h6ZQCvDH
qKgwBuG6Otew62HBSuo3DYjGGjkUJXPE9trWRMogT0yp951QPqbJXcRKKyqdubi9d1Q93tFn4U+H
qwGbNTpn1YjqHvjilsRwGcS0a5WRD/mgUUR+PUsgGizsWU7dMiqydC4mNdXnO/jTVZ8m4AFv2xBV
0HplmlEkelRyNuwFj+zYwvehDzJFIYLZ2RWK3zWNnr9AMO59YUP233oGANd4DZCT7LyxUaXxjmI5
FqgVd8JeBhfE2bHi39fLQYxK+22dwJisGbkaM4eNQxY0vVPuo8yKuGQzjCSiKJUwPIzo+LNxeJI3
kluiciGB0bjfIN+glWzfjcegihBIZg9v9d7DXrw2ZSXwrB2D+UEsF+6OyPOHT3T42rVuFWNozqwK
p2+a0GcF8o0z9ncU/Re1v4TV1rXWAzW417zydAaXjfIwed/xLzpfD5k0SeAGwMxMxU0aWubLHG7y
EabkiAScTYmIt6BK03c/cZWSuCa6wX2Dz/Dlnai1A2L0OsCHo1Z2FZaFAEutMuGq4j2tHnpz5B82
KsChJ7kV9ImDMMEYYHpmzJw2hJ9TuXxpXRvCTfPQb6rpMEnMQ77IIkYf3j+P08Z0eJB88U1PinC4
AtZAYHDbog0Y/oTQybAAMFXdPhR8VNbU8Yl53Uo+zS2x94JwCdaHSvK435i+4AT35LnrMAmq6FBM
PxyB8FNy3F7uW5L9tHUlH0p7ynhI096fqFcJaPCckp0VYCTYW69JBkTp+cagerC3GfvcXSkd0emu
/pkB194Pt9iyIbCDZE5ETDgtBP7epaKUwQU5ot+c1mVDl6JwRLp8UHbyCwDGNjeSUKsYXL3TtO8T
9cWiZUIaCmgKgXzaLULRijx/lP475qcqy/GYXCDkga5zDGvWR/CYO/+MySde9PoZokV1t1f5fNq/
OtBVdfy7/E2QXlHCuO2PnJoRODqjKHV0zgy+jUFL9RLtAK5wsPSv7YhWO2nL2D38B3qDq1E06Hwx
bOwNPHjUf2Vt7XLJ2XDfA8wNCNrpCKTnSoXoMS2GoKi1jPmDGhwtnepuQN9HzVQHA6/PCw54xYl4
Zc/tXl6g6YoBR7dQCoHsLcb7b5EZPwTIc1jYr/XEJdXrNLdgDGNmjxkAjOx/8zI44LWLYBfA8Gq4
RQGea/TIxKLRe/MkOCe5CasgPcTu5itKZMsDrxr5vchQVo/etLhXfaBmDkRikQKIBq4RlwPq1KRY
IDZDuWKbSBDSXY6Y2GwYtjNayidqxUmyKwVrjXg4MjjvULv7J1pY6MP3lB8IFjpkko9z8j/vuKlc
qq2TfLb1C0B+R3vNw5aBOlzBWNKKvbg2VKCf4WkrXE2+nZtxj/NyeaQpjCh/sJYZS0IKW0fd/1NN
Q3x5LroeUGqOs8xRcKdz6biKSIVLa+zU02982tqPQ6GJXago95nlIXBmNyUX6FSCR27KB60IAVxk
6CFIuZyODRJ1YYoLqGmzzb/hDuNFynsVk1d7zvdyh+aq/pjzfZ0Lfh94ObtQ4ICnwsy8vlW0q7x3
okeXRCe5taiBo7xyHoNLhiwDvbTjbIc1tJPKNubh3UNpRQsMF9UGRlax2SopIwdokKRwVg/9fkD3
CvbrZ7se6h1zZuEX6WaDWs4o9AltNDk46ULrxnj2Y0Frp9vQuJ91mTehgidZJjC8Qw8S2rYrVzLH
N2PS78Jc6o+NfES1rqePHt5n9u/K0N3kpf/L3nMiQaE52r6849rURxDEcILRm9N77DWHf+uxEFn+
KHU51EcdKVA4qVJcihZ4tpuqmwIlkFdTHQB/bECIJ1OcMAmFtbRav4sQCzD48yoinCYX8ug0DLFx
IcweQSLzio5LMtAtN3L9CtsDBD+fC2CFNIgxjn+K+BjCk8d3UUwA5Auh32ucSyluHCL15UwG5XWk
IEqKqMZRIihNnXiWXiDM1SdwrF0FN6w9b98r/sGBe0yt8Dapc1+bHANJcPFE12Qwn+qfOrIYufT4
B17l3LyQ6RjxfhmMgx2hp0+xtuaLLdWbocJV7PS4qKfk9Z4KpGajCS0IKooKmdgalRi3t1rnvHGW
MBtsZIivFHzwIjvE8+iXR+zDq62b+ksDwmCLXCpMWHtWjnwan3iYki3/xRYMq589rVlbnYkuiHwZ
XU8jUOy87UzPyBJ78ClZtmp4xKoSooR8onr5D6AuU12T78yvQGjWr2GKMPbWVPtls0JS7cNuX2xe
LJdeR4PYy+zMIRtQQNvu5dJZCymsyzeRU7mSPW0IlPVy+OxKAOvcUHKrcV9ZAe8pS/bTq5uodwSw
wJ45L43tely/9UR02jLMDoVmeaDk99ATD1IYVzQ6KOfINx0JEaSgECffi8A5Gsi8Nx3qMLXw18MB
qnzwTCaqkDPiF1LiEMEi7U7Dy/e0tH7u5+FdpHI1X+bRlXVR/SFeB/PxKNrILmgidDW5Fx6SM6Fs
Jbw7jGwWTrirFECTItmN3lKZuLgOA73BlCwfaltL4+KA3TL4saaqJVVzbhRSSzoQf0LLktfLfSSF
sNP17wexiUtq15lPNNud4wSXHc9glrxKVv6Iv/9Nw71Hq4a2lqlmjvspEk3BqIxX+tAyTaQDNQpN
FGcgwfnfR0gbFr3BiKcwLa4XSlbxHDoVkdJ3F6tttlQAQdBybbGOSfMz8vZg0x01tkLSadqceyQ+
A7cqJ8IBSCNrqDuvxL1pe6JoFDuQSheM7Je+yyyypElHp3cS4vlf4nPh+g3x5fUjNszjot1T3kdL
b5fy3E61as9g9t543XRZhnEJEBzuebLZ4cao02YL2mWUjOXDh8Buh2tIu2GRjEluZQHslKfecLDg
tVcI/7r7m45ONj+8b0AWmKqpAsgkeb+3x1+oWpRwMIKJetkyg+rtHRzLC1hQnfn1/TpVTxmGm1aN
f8nTtS29Z1gOcm86+SDgt/P90n6p7xXtpWTB5pbgzp+xqil7FuoAr4R1zExEW/XZwzIEjYi6OsFw
hjFHU5SrYcUS1NHe613ku8OvuWmxNZ1APLD1YWvd/sNUaA01Sj9COGedX2AplKm596ZEprVhvO6h
3q0Wth27bXYKkRAleIz/pdT2u+60/Omjz0QR9nP9LjmuIlRfVOfEl6z70pdwSHGtdZvVZoJe+i6x
bJe5fBzowqb/kfNt0Qq5Hl4CUpYJGmWjnoo90FDAVeWkTe8hCCt6OpMIRh8aCegVJ/AvRndelMha
M7MQ2w+Catn0OqjsxmDJhogOZ2aNX8zcRwYN8/7exHkPHPV8wCOgV/dIpd2YHYTPqR/r/UExT0rA
xrxzZUtHEypfZ6uYBtVM+HXV2fJjZY3wnK24taOcHUeRllBexcUCvXyubSKsnjIdY8lfD0CWD41I
y2tRvZ0AqbWtGMaRY4GkCvbHqOJDJHwWOTMZ9QAcSCbnDmk3xxvd1IheBddon4WBTJnZeI5BHJRu
C/2CYXOujiybzrZM8AMVvv3REzxgIY6MrgUBcAmPCc83BocBXBGl1LW+3g86S13AJUL5X7d7MpH1
kZAIjcCHriE4JvWIIe4txfaYmG++q0dQLnLJ64Z7PGiFAJ2evQ9Dn+dYnXqpM/TzJ8lo3fbJdCxz
Y9Un7+D7WTIDVK1bgy+e54N4hUhj9z+bJRYYmgkDqqsY5l/93uwZUrkjJ5lra/s9E7Pbv17dz0Xr
yuFk+NzrLPVaX8FqeFfTAiP97n6PQWSB12/SSzndNQWK38E7dLeGxhUhuc7sbLD4RMgkrrbfsPyG
LrZEx7m/BX+fHdtlv6KQUSRSDcC0CsX82/TYVz8M5QGg8JJSab+ZPlKjYDuBM3IjHNoIoURtHUla
OlL4C9MVf8PzXhrbqLSrmgNMeK6tv+TPPmctm+A5A0Cuk3wF069XdsHrUzacKXo7XUYpkSKoL5Ym
XUuuNqrRlIQvrDd5HRVAuZunK3fijVsDVhu67IRFPWadyN7YQtdMgWhVnL71E0Mpm1jFvcTLzhz5
72RevyaruhrJKC1VnLlnxcRucg9BfjiUFK1jSaKmisOJoOizE7aylLS7Jy/bjbJx3BrA4mCatcrR
UFLXmbsjjzI6DEGxLn46bj1cTbERYAd6ZTW4fRRw1jzTrO0n2bhZHgb8R1ddMd8EGZK2k+m0ukLT
ilUZQ8uFoZVJcin1GdCe7BcQ1Y9Pc/j9zTRMn4F+vFu+qgdSUUrf3wMZFS+jjhBdaGTXvPuN+Twy
tSmVvm6663vY2LPadnyLjx8peofuYFpNzve1C6xNT9/v+POyxYrFbIc1S9722ipVdnd4WX7jbtz2
G4mb7tRcooR/4yLzfGeAbHL3bFH4ItKHXeq00YTJPHYxkXfVxFLfhQmgzqTS3ADwZSGPQPEKC67P
4m4udX7PGZSABJbedkh8454+CzSkFy4qCJF9hXJ5SykzTc93YaQ5EVfftNBvP4Q29kVy4+t/Vm8/
31RU6gSptLsfHkk6SSKZtci8UO25th+R6Wz214+zZGXm3KsSuudgG4XFYZtTwip6bQPPnUbm9CHb
8zTY1yRD4OMcCvrVKMSKLGXCguuufMYpXl++Vd/PxkBB3cmvIlmrNngWnK+BRmwKXpwfZa30aGQj
BaYja1yrPLIzXAi8sqBmzJFeKbiekZaiqYWDoNj2OgpJbhQb7WElEfQgRnGDY5YbJ2rjI2e6pBll
jv/pWwMcPvLlAKtm4dkLHf4OXAVlrGxj0avJ1iqBebqtFNAEn3t5QQdPbjWDgeIPzvK3RC8QQ3tL
VKk9AaJgpVccwLBjK4Gobiw7LPisRv9kA3CIzI2weruujs+XwezkxxaseLgZF07np6uOKVevDq+f
Sl7rj2yEF0f5Gtk/Rnxn3axwNcEBM5M45YuhYA0r5vuL2RazllOMGLefaUvF/YK8TtjDM0iTOLrx
hnkzoTZIh06ogby+ktGDSBOcIgt9FbjFcYAr0L4V9ceIZpxvcr5CkGEyzF2/lgrc9mTK6iYHU2TE
8p0U4juev1xJAPkIKKPK9JfcK/lsxs0D51no3iyKC+A9VGWo56Und7xnIVppb9ykrfPBP3m6+fmF
EXDxibWSmjItE8DuNcIPI1Fz3ee3RRfHIJUkZBwx1ca5Zu5YPYhhQxao15euZZ7uCs+STGBTZw3N
u/KJP/loVFGbdxtQp3GyKt70m7YRN10gOFa8RL/hfdgCBlVk2o3/OdqYzGFcDUVBKPg5ZqCJb6US
yb5uHxc3A5vgy3vYV7Qg0asnl0CeJbwGwP87/yhhpkbiFY2/GxhSbgjEMZu9ZLMFH01ntOPZOi1K
0Zoz0V2fhDjVAWJJFp+5IUyHkXtfsrXNaeBy6KgIVFX43x/SG39gUkjyWv+C4k8s3a+OBRALIBuC
oabyYG4Xxpf+K3FGyYrdr2iKR3HTiuz3k9QyTVjuk86S0LkGmsEgjDgBRCpdOLVi3tu0lPOEGFNc
erBQmCtziBFqhqypOVYKKgjNX7u12kd5oraL0QfiLwhwTBObZ104qhUS2jhhCwREPKdsWffs8vqe
9YJ7N3bw/X75h9blQzyN/6BHxV0tFuxHQhtBGSNlLWGcFf17DA7Dh31Hbr5JMLmhfrjkAp3VpSym
PuxNruOHbmuMZZAWlYmxd78klmJAkoFZiwLlf3h+ouv56Bn0rzC9sNspEncDFrYksSHDslOLSIGA
GB5b6jYnfeLwMtiMaDOC7wPWUL8qi9wzx69dEwjyEILPymWs3GT0rZIPQ22EvS2fxx19xJJVecyX
7sSG4bpP5J0RuyoBSudOROeEJrYKlS9IHZ5aB8h8WKTEsQKTt0EDMt4CDHkRVUlLRQcqqQrqsfxA
0g+FP+MgNgW4U9zSazM0HiH81v7niZqFz9sH3/RvQ0b6ce2HqSRAgOUB488JTGYXpkSwqsubZGEf
Tx79MSkgRBpTZH/rFqmIxa1d2cKtaOm9gQ/jli/XjmzgXphi9VVebLgQTIBPT3O6ZWCxwoAq16Wn
wAwIJGm26GxQZo4UIoDG2jqLyKzoXjDU5TfGJNv+ixdhty6GX4VyalTldyF6j3g2RADBdA64Teak
98ViEj0bPYCEShQ2q8m0/Oh9SvGhSdtLYDv9VoYdaOA3LBzhfDcrhtd3lEL4wWOVUJbnb/8PL8st
1SjovSfTJRATLd0H9RCKSP3JwEQY/ASMsRTULvXYwpNHOodmJZ3+3KvlGaQVE+A8mQ9DCddUGE0s
91/hFE9jYn0iybawBMZXZ0POSRAyxIppdwYqEcbSS/KDH8zUwuwX9ScpB5X3VW/lvn/ZHomZdI/s
uOD6mAvcp/sSsRbzNcy3XItr8hidh5Vs8MCcoCa7x5B9sRbNMMNAhp0eJX7tdB3/FFhxDVxrcIcP
+QSJEommqfzbzIFUF0ACIsINiVPV3GHify7rJfTRGtUL1DhWEejrBNwfy2K2+2kpJXLLNOViAcY6
X9hPf/sxa5F9/Ebing9msmqpb4ObI/XBrSr82S08o1FkltwqVyBWwynoMfePh3wO+EiujOwFTuDi
Iq8eHtZmceCIqsqicyO9J/ZQL9+AZVeo9cmwLrxCNJAKKOgFUSRdENumRvrhbHiBBO5rNxzzYb8k
oSI0ZkEx42l3o8HTN7HWPhBe0pNrHxob2+gJVI+cJ59xVhZ7Ey/M5h+y9FkuzgB5+ACG1CTj8VCL
lWyHp+B3AdEhGP796VqgsK6aZKC8B6Fp5eORpi8/LHjIuq/unL7nush4mkJNudkcTGH/GdwJK1ei
juCWIg//zeTselW3EU7l88sbfKBjLk9PkHY8RbjFRE+0vtBRbuOs1AEH3mWbt9wyxm5H+tQgF8/O
VShA7bxTBJaCKJw2OeUcI8bhsbx3YyK4I/mwkUFajncX8Deak+6kiITw34JYWmQrGCSuhbQjsySc
8mWSLrD39TQ3ZVAfWCbM6TJfrRFsNQoO9m0MXAtW9ZJvwvH38BZygcCW3TWPgOYAMnaPeQ/8QyDK
AtUcAGZ6HAaSV4M5UG4uYBsmtfMvPrcMhSYf+VcUBm1JEjMgIT1URGFABhuZWvMnlhaa6ewBrcby
XkIiXNRsYuSWWNDCPtmGFsYBuA9StRB3Lkor0vTn1DGpe33iFzelhVB5k7JSNGu5w8D02ri8altN
fBexKXQPCV03s5hm5kJgWHkdjGn2LqentXog1BF8UHR7w3KJIf/p5nGrQKOMOa+eCpa1/IIXYvd+
DFWFPYQSEBN6v1PepPHsHBwT16WKheSKNNbl3aeUjHLoIIwMr/ELEuaa4oI8XMsgBxNJ1XNKzTm7
sdn9UP1hngj8j8Pw7yRlQR0aEHOzXd3x7CL34djZLuO6AdC+k9fiAHvuui+k5eQQY7s9JQlk9839
ofc4WLXTNBa+fpyApukLWzuhRGXQL1/C1fuP1M4BJKUMJudlreTFgpaxfWTknZmdf/kPdKFLeP7N
Fj7JylToLtblNW+ifaAp+EtylppQzjPx2AK7pL2j+QNKoUkfPvvV0qqCimNjUkZ6gzhD5mNUOS0G
nOMb0UXH9+5huUOsJw/yU2zw3ujypecT/+2qeveZN7F+zOxKiu5Z1siKzi6ERDz+U+i5wblNmds3
yh/WCLhS66F8ioV59Kd+UAhYTDPVzqRg5+lzQOpcLtxkhwRxWQhorMUT0Cd067Uk/bByX/PN/vsi
gBrP4gq/IboWQhzl6fdJvgFe+1hoSXyDG5sGEUF7xLE3ngFNfP813jV62O4VP6QqTKpyl9Xp0p1Y
3FO4m4SkwDPiq6xZjqeYXtODi+E6+iCKcMT+PXXc87HbqD/XszDizRIzzQosRJsEr5yBHqUSQxb/
Pm1bFiFm5Am377MIr5OwjAkqfpjB3yAFl9VkIgmBVPbtMoXcDLrjz79E3o3chhC+ykGzuVQn0DEQ
t2NjgpZ0AneRWGs+4EFeVTpHsu5ep9gMR63xMYAUrgQYkas95mhoc/SB5ZJQm4QTZ4duKTTmqP7p
AmzCzq99F7oLqVz4Psgw2vpIcy+itLwtMleQEVWo2nCey57iv09Gg5+JQDVnB0t6yOfzMjO5Xu9L
xmFQaiLAv3lyn8sNrjEDBStcQl7cD4nre63Fh2tUmcEy+6w78mA3K4zr+Zx42vn4LqE8NpJo5JQG
AatfQsaerNBP1NiFsg+iUoIEFWnpHZ72SXQji4IdecegZRFVm8L/keJiD9h81KYPqJejqMVcYy4j
0KaiQjAqZhrYwvspJpfyKMxcsJNSyWklG5uCOILbd4fhjxBA5bYQmwZhKZ62B5sKVUKIsPoouJ5C
zN1ME03qV7/3BZK7tfZqKWK3f632y2bXb+G3w1cYFoKoUiFt9YDjG2EmXJ5HUyyreBmiXRWRtvJh
dFEeiZ7P6qcFb9bUsYc64mkGuOcxyfUVtHjN9aSlEk/321+4tDoyg74Qdii9MIr5+ekQgLFb3PI/
80AiPhcv/eKRc9+0KES+ewbVmwUughfLzWRNmqNsPCZ7e3mfwFIABljYN8QM6QO9SYUaII0EZXv9
bV9FVKvzO04nnexu0o5LdTSeKJNYpOm0Mc+ii19X4tkd6NmiZLf0Tvp3zAmQXqSXMCNuR454t3A+
VRSWVX+ADGoE2vQIrnph1g7tb7rfxRzRG0gCRej4ZBtEmkR6IsbLRlb1caQ6joiJBXUFqxVRvpJ1
XVJk05sMb8DnQ7PU7oWuAkxcfDu+o66ZdfthCWxkmENt9+9HU6kb/4LyMLjaSr5+kod2KCrswJ1a
v/80PmDAKgnhO1UCOyyjdZxsG61F4Ylysq63Px7+Wjn4ZoCEHcyG3fW30fKu2VZqyzGTxtBgyMAt
44vQTbazsNG/W1DYwIddMXIBtXPbpH6nPVjbOucG5lN1xKuqkdCaf5kNoj3RxJU26vdm6TJ/VEQW
KNq7SFszQBdECBy5jLcRH7b3b1PsLXAEh+ztquLWuPtvvD/Rz2d0UJWgbgv3IVF04eomoR1Zfi53
TA8W+oOaw+JuJgOBI7Lc6nOroE3pNBjZSS/5RD6ETtbkMC7FlkcL882XodkTTxd4XKRV5cenU9Pf
jKjLXYAhYtMC9I0k4u6Iwcrkq8aZGabzhsujuIB+PctyuB0DvO3QiiTilSbUuAJPcLsJzQP1I3YP
GgrAGDgjzlrTtXH4gy9G5ckTRqfrrMHbTahjJn1u7zF7nF32IsyQx2B0n8I8nqygJUni0DsA777g
/dDMpmiW2XxLQaqIVaxVeXVLp4XhXAWC0yhw2qJqRdka3KlYfbcMq2VI+IeG0XZ2Y/6GYS1RKwCs
DOjSCedhn4HefWxhuDItWOP2vImZCJpGygtDIGg8TnitJDI3DNCeNwgMuT/B3NVNFBR3YJk89++Q
tNCIyfu1HbxBpyYxy6EArmXLdGkOGSzq4ofE3Xzg5qI7VU7aAd1PIt+stg6Nsx0kY5PeUo3+G1rW
WkPyFxEgaMWHyP37JToZzzUeAIknIlZ90jAyGRd3NfatRIWIgL/mlWMvig1LLpm1yuNhKvG6YA3Q
DA6VVo/pjHqb0EvvLEV0F+4Te6OtpQ7iIqGnUUwF8iNtXb43AIbFu0o0VyLm8DIHSHbVPaWf3+bn
KgwoaVLBT7KvCIeRprqPwqyHlOUuNKpzv2H0miBoiIDJdhC4ypwDtCnE26Jco1U9pVUA5hDa68NG
oYzc+5sqGPQAVv6upSb33pk3GCDoktEnl2qGamTMb554j2Rgs5lXDxAtCoh2PS40e9lFcJwtIk0i
vqkZpB97Ad5agmr6TbxlSOsA1FuSUTpK/HmnIczSapWlOnXm7iR1AanEgqZDS3Q8qWSvpFj3LXwl
+I9Khu95DwWQS4pF1iYN3rfU5t1PB+SJpYK8l6fBux1hGF1oYMPfmQmj2Tek431awBGfYpUZXQPt
QdqCUQSu7m6KUSGJsIuqRqzmNavmyRphEqZoQ0ifoNebLl47TwsF7XCX70HZ0j8WIO0spOOCfTjE
H17NEA1YahzO2PRUiZPS++/Zv5vvAul7PpsM2E1M7vjNde2v3ZhKdVnbueaBHoo2k0stUquSVYb5
UkqBMPzVCiZmVllSSTi7Mn3A+ximNGj0skxv7kAFBQiKIwVs2cCPX5RxsgAYl1jR2VEXTaEdQNGG
H5WnAuzloo9/kJQFvyE/xpBD3NhxcIeqpkDDSY89fhRSsZnh3HKkCNwScuAqVb8hK68iXETYWFS3
WKw3l2rYl9yHSkSqpLHobbOPRjUszPtxrQR6GeZtFTpmEPgT67uCQk05SyIEDXtZywrGxvP99ybm
4gI4VVE7kFAeZNDgxQ41HGXDIY3Sj6dpl5q+cSQ9vWAS70t8cbyvNQL6xxjCqmIJ4ajhBvckRzAo
Tu2J3VoUmrIyUHuU2VEo0narsqxHRCQrVElduf+etetCo3WheGxIJFKT2of6mb69KpYRp0SWJeiL
z0dDYCIA1Ef6ozRw88jbwsR/UyyDpQxqBcNgoCL9DKb/or4k5Zrlsr+eioGckbTBYCZSvMCVgwld
eDm5de/fcisurR0js1A2jq/oosfmpTAZIzjfQRkhAyWHKYaQuXExnq2Qp61F4WqaLHRpFD1kmg/Q
hKZO4kZfRtG/5mPp7K8hJQNmmbLxbi1yenMcVIRD8xtlIqLVTgINLroU8K6HKEqbQ+yjIdt7esEV
+bpCVVhoUry69yxLVXsI8aisHrG5m2O00g01Sv/X4/NDb8lI8PIM/g2KDqlC7Bs54QgyOmO5gcsy
SLL3d2u1aEksb43yM5OcpZaIvHuNQl7gRiQoTcOasRQfEWz+qVtNMXvVPr2CZxpZhksCuq4hDnkW
qgTOS6dh7I9zXRfoedCmwJswOw3fTPjSsw101trbaSwN1rpJwN4BEWVuP1ZAptLkZOzuIJVsJysG
GlaeRjGsFZC/no/ol1IJ0G7Bnb30qn3m2YNB7YIm+4VGPPnAcMSnTCoeJG4UVaeiw3j8sYShwp1N
MHyIA+bn4t+RAOmx7/pcfQFCUq+6yA7T6PHNp/hYeLtarLX9v0L6s5qmVuNvCbi4vy4z0lInIzJr
ubKzdDpckjPwQGA4EpDF5T9D+guyxh6f5qYDtZSxJnqSeWnibafOKKpKEr17HShQeryycerwTGBR
ZAHjCj2CufRrKUmH5JcND69tlUv1EScTFxGxkPTLlxiowqJxXEb19URBughf1zvxYkDk7m/fYRzC
cF/ham03lQ4DQ6oA56cHcbnToiJHlqrk4dJd4r3gYKOYKSKNMM3hf8z19Z3ekMP5pJOCT+U9cZrx
gLiT7AG4ZDPy20EejLP7y0WcVtx8G/uFu4MiQDnOta7NNNDf18oA4UP6BhNALTbBzH0Uak45Gi1L
TmRRBoDzSL/gMgXbaXbhHUP2VwWdd9fE9jwkvPUIcvIpjB8+wcNXa/9lPRVaYh/VU+kLQniyyfRC
bmPv3yZe9fAev/7kYbFiaTeAh93Df242aDDWfhZ6h2kfccmR4lUsa8mrreqfjuQOnIUPPYCkX/pK
MuCkvpRH0sJ5jqcUFq9NJ+rE8Ng1H6nhxrTg+YIqgL+cJitRBnqdJLDShI71PjpAqbr+516ZJSYX
0Hz0GwrHN43CevlHbDhC8AIBn7+1CpWc1euRnZ+wIPXgkhglNP/mKpNiDgXWsRLn4zXa1Qa86Byy
WRjZg9HdXivnOCTpTpS7UGtbK1FkaD2rfiF94skSSVjhP23jUTK1TUCXHrHADXG1Y+IQI/tBSEyh
y4BuB0hf+I1YHxkG+QTUIsAdwPNTv6GemViAZvZiyPXBQby25JQS/AH7Digi+wLT4J3aMd2dRXu2
m70xFIqAVp28L65QTeW84XdSXpWkSE+KS3AHLzCvpa3tg1Upm4kmV3ihfAflYTVqTaS4TEgy/7Qf
TZu5pi2ZedsprhzKI1cLHjKOV3mDewSPrsgECeoaCTw5UZHul5A+Dm9ZdyomhdWSNck9NUGdDr3Y
gWFAXKl6xEJNzMWEyqEgmyqyOxpKWDkyeRx3XkQiIKAm4CsOfsFZOeeIx5tvXmHUBSloY6RXcLQZ
LqvSbRDsne5VgfTVwWkoPddp3bWI/0ll+vzKnbHhmcLt36G3Kcd8EIvthMU6whkAcd0+B5+3fb9s
GuIzkYy7/ehxjSTnvb9WzqjgBzbGPJuFCMwlM4DoApMeXsntF6d8MFm8Z4DB40wpddMcawljBbqk
doeoWPHD3q5oYswvh+zAfWqcF+VYoOB8Esz6U9Q4maibXKNH7dGplg1jVTiPtkag/tEdU+XckDoq
ExcJ3UjPfl2nuy5dZVl3hzL4UTeCn91yNgkrTKhkArPZs6Q1oHjwRt6ywVQMMMDz90VQW7dbGRBf
gBkdiQfcdTM903UK/Z+YmEgH+mpEUaD6n11daResGK90zfSszgw7xN2oDYfs7TUwHOpyUD2XmFJH
OseMSBv2MR7JWGbc0tsMNh4+LE0lew+Tx31hkGpJuy3sUgcbFMG1JuLNgbrvmGPz4KxgRShYwGBn
IX4jvOJG/ojoNNun5as9yMvGCUDMDFqKpBDnaJfU7BTogQ/eLF5AVEgIfUYBs5loeW37LFZLQzNz
fXe2GQDLjRWHZdgfTwhT7GsNyRPZwp7q1Z6Z5ohDTp7Q3K4caX0MrLW4EDHaNhQe/EiC/CDEdmO0
xp5bsfb/MjhsBP/ManHNRtwk2pvzCPDnnVDD/csWl8xskGgCoVkXaT7/9Dod+k8wviQIz2bmrCKw
tE8nCXZYKiQ1buLAf1lHRi5/wIafi1QTXe4cYu4OITVoJUpErTndH5zfbBdE+O1nWYr5483vxThh
bXJ/qFGzr8Wl+NGrjJ4hcCgTOxgoJVDEIXJS0Kj39eF0J5HqHRpkw9g9i8bdw8Snv6jduTtcV6DO
JNj+bbdPAZ04Nt9BjfwJ2PED23kHOXCrVbvfOX1GtkrG2TQyY7dfQsfDipEUz3beuJ7JIue93JY0
WlbzktszdY4+pXEk4j3CXi2pRrG0OW/vffBtrKsg0cpFRim4XNzUv7HPXW6icXdiHtAeTYB5rJqj
zcYlrAFDxI7tjzTYsvU4+63aRWZg6PH6KKPGeuUwqj/Tts6ZNWWfeMHcw0bTErKQYDBylSTBv2o+
j/iiYwyQwj+ThNbJi4DBNRti5a4TSlTPVrzYiB4nCHGRNL2Vk1pw7wZ5ufU+tDng/KpkyXa7os0I
uQSt40qVF6173h0b8RwDGwzkRrEieaUQXdRcn67VBIYG7ghq0MiECX2p0tel9EdUZolFq71HilwC
HVidfKd8aghLdplpMSfHVrsFCvfuf1xukhJOLkiSTRgsZUzTBXOcSzvDuqggwUeOO5uaZoQja2Ha
NP9lkfYdpBOtEtefmg3UnTE4Q4zxcZMJxoc8J/o8MKdEzTilozlwo4Z9purkKkbkbn9l2Kx2rafd
Hv6qdY9i4eGU64VZrvIj0RgigWwYV1eby+g4P7kTVt2vcTbB9qKO8GhzZ5wjsWX6D9MFpCWMlg8H
uYkOCiwAwtSGR4p7U878t1cTDVjirUfSTier2C2D4+wLPcR5ZxG3ufjW2GKtzYgHwI7LxFeRm8Pc
Zu2fuSBnFRMpJZRSr5WsCCIegwpEZy7nOPcxrNJPMtRKLDMlzaS3g0U4p0xLHoFcpnbqjR4JOe7n
+d6Q6Jn9ZWqAtRk6QnAsqzqsiLHjQPckMUZPbW0/PWUzS0QUu9I0qx/dczIKKhKtdtb+C7KsgM/U
IOMbqBPJA9n9GYcU418Tb+l+mieCGrTDTve/BU1PF1WsR81PBnj2DY2LpeIVmE/SUCKVt0/VeVAI
xQ6+JUp8QzV6E4wfnsQdN8vTE1lVwyCmICMnQrid9iQYlwifdrBiEphaEXMlXrK1/w/WDdLBjnaV
bnoabYuoc7NRgbV3GgRfqIbirKYWNkfr7oCEVt4tx+67/IDGDz0SdkhrAI3NxLY25gToEV5BawyI
IV0K8fIf8sIWrJli+iIYDe+hCtvMuTdoOjF0jNa/JoiSUDtJ55f3gfsP0dYU7I/nT7aAGf1dT9as
BAES89scrRRjjhq70aEQfBu2Cow43my4vAH9H9Y07nzu297fEZ36jyve1wehgLvCfoTCFC6BxA0J
WXmzHod0oh2N4p4ZmDlYonx0SWRmXxZwBU6cXDVHR4AJr+Qah60NS/r7BL9SslwL12goU6ldKLTq
42ED+3RsI/dJ8A6/buBph5V+tYW4tQ11OPBd9J1kT5ibYZGSY29/oMMQBGD1hjPq1mgzaFd/9Kb2
bcjdaI3JComxCwKMVKfGQUlM5osUYz5spy0Z1staboPHJW5DruY99Mizy6nV2AxdYUt4YMunjxDz
K6bd3lfKL85SY2nRrZKwsJ/pe07rqw1ccOV26C0dbH5jufKcf3jgpMhXxkABiTJMBOySJi5oA61B
HhxihQ4J8B3LqUgnC20ocxGJ/0mNRxHpEyJyPhhOdrFePZku/vfzwJjXUnFGNI6BiYEjq5ED4hVz
qT3W4xc6ljHLpULij56FBlVnf5aSQnFW5XSZzeeb5a9807j/0XCTujJpqNWRneMixnjYfg11FJwJ
oOyNuBGWwh88Kg4qheiiEDD2oPFegKAtD5Kx9/V0mGQtKAzB9WCUSbQ3f+6Qn72LHp7v7X3Ivbw3
6BvNwm3rqMZujv5QD92L9p5Kpaocg6OM9ugTRjhX84N2T7g0ksD91+7+b3wUgJFUXJnNN2WWV+dR
CxeO9w9L+VDKYcjpXTpN8RQLByd6NNnHXS6ujFHF45nQb6ZCxjDrh1oxKk0gSm5ppFNC30QplGU+
1QsbzzJ0IR8OAyxBRs8PLDvXcKpNZGQTqcY6oKuMpYIA/aONrsoYT0rLnDncMjoE/ELK+EuG/gdF
cRRmFqKoU6E2/EgXiYXx8VCgq7hqAjR8IprTrf0kQ18CAByd9CatXpJX4lBVXn7ROEQ36QQnHbbD
FlRor+ooIYxnYF2Si9XM0Zq6OHf0t7G1GEYTq2agyHHOJ4KDdXQ0O+Yil5+WvDAzxtGUIO8ZF+9P
ftclpG3uI/p9sGb2B1Z3AcYCoTwWuIX4qH+OMvH5FaszdLO3xcHJtt/UipklKPCWGuyYpjrwTFID
aRh3yWJIL8UwMlCHUTr4BJVQ9zJ+zngh0rBWx6UbCWb3VWYYHdV5NRjKCAzWn2GSp06IwFqyf0o9
K2+V1VJDuXey50QX1+wkuILg1vLdk6OBhaa5q+rQX+TssSaDb2IXcke5p1PcsNDcINKVlBgy9DWt
iyl1S0p8qwmLVkacUf9ERU6yPUbFxWRgtgwpkdf6hIwH766QrmTRun+GFLI1rcDpVPNMKcziObDy
vfWkEFPPWTou/7G5ohR+nvlh75i1GDAOf7cD0+PQ0YBnWq//mh/CmWcxCD4nRXo67twDhszvdtrd
pUHjcVDF6pu2D1baWy+czTyiytL1/obWDeCAxDp2bTCJ66A6fpqUVV96MfiTABqpivcC7WTEChG+
MIfFPw84U7Z+2mCEa/jgVjY5lMYc6hRjpmJwOsLEDtSHpVboSDqYiW5POPWQtBsMNXVxLRE4/dF4
WZ/XI8iW22z4+WQiLfBrxE61ybmmXfR7k67IKDETfUX9PGgmaCAh6VoNUMShDiNb5T3c+5HDgLUP
AHRtMrSZ0Kl35wb84MjBf4QfNxltCI/ZQPG4Zkpgw+wxGh9gxC3Kpcn4Bf76Q7FcIrOebvfHtAO1
/A8Nm0EFz2bhkm76/NF6k8UiatNNoheG+kpoXqX17M+SMf4qa2QWkt6WfoNs/wWMTDOX4lsZiEl0
GqOuySK52pmiEw/cMVZbh+9Tdf/+alaTZGw9Z4oJsPTXoVGKdHgxCLgS2v8dy5oIY9mtQhEIt6uc
CgeiOsiX2TdiFZzWAvpPfv+F8bjtgS811MKzJXebvsMg+DWYKE12ZETcczHXSRjxWhqnW4zFf2wQ
RLCXgmk6o35hytxoqWGK+Bd6eWhsQ98Be12EPmMEw91mpJa5pFM3V3jhG/M12/6NMs85u73b6lNa
ixPCsS9ZxDc+e9Bw2Dyh5UvAJAPtAsh3R6kVm2Fpk0KE7pkvEmc//ax+efeiuWhNpAerBSHkv9+6
iwTU9lgwHpgFmGLdoXtkBoG3gMOKEfcVIjI/m2GQNn+/oRLBzFYPtdmDoKASkDKZbpudTyUFOpfO
AD/sHdoPSF94D11aYqdQb/lfsvYYK84EyB6DYqPTmxS+AUQCLEpEHa76kaq6ILiOXsaQEL0KYUgH
MfTrjWX5TqbXEAOnwHwMIBx/5ExnzQjLD3HOrYmxU4XVrS22kBdFHCjZLz1PX37yi5le5txFxocU
F5J/OLswlL/y63/Y/zJwhFN2IMGVDmAmG2cyD6AvW/RxzMfPo4pDJZNOif5CwFcd9tDiF3PpSbZy
TobK6sE1f7EJ2ZDMIbNMLlgafxArRbazAm4zVBVUZZUhunJ2TC1jSKi0KwcsJIkzRYZX9UZFuJ1n
K9ve5zOFvSJ4H3C2qOKWjgkBMEDrKHhsNSTPrLtoyZe4A9vu8JMB7oD+astDnzq2JUFedMISQb3r
H4uV8eFKBnRkKM4LIa4h1AIhW2jr+M2pLMZKpmLH1hY8+3ivtw0YWiYuz94lgfx8wldp6voMtAYY
o9dhedpx2RcNbWEXgY5BAO/wTIM1dZ/vJfDFxjF9kyg0zAON+L+FTZwRlN8KB47jhGsqFSK9DZQY
TkNbLSqs8P4lFQbT+canYl55OJspFO1JSzlZLC/HfO6PleGC/OImWCEloMAelW4MakdDPZb9hYGC
CJfNqKk+lYvuzBUxpo0GfPNjPvAlM0CIEA0/CQICn+9uRDqDDxQrWAUeRgbVtMG/DB1RWxLqbOqW
tFbckOL/Y7b2ofY9FWvmH/pniwI4mDCcRtzwlZlqUQCQa0oIMViUUrNDCIXD4s6JM2MlH9yCndyN
RE7i9iKe0TklwwVrkKEUwzisUHIvy4XFmLanMFj0y6SKgOfLp1olt9EkQFSd5WwOcYloJggSYw6Z
Who3y7FbUYcm6miy4b85qjv/dDaqp2NClZBsPK00e3lFiMq/Y7aWITR+ZZ9B3UHV84z0wKY9ciQX
Z4FPkyPHgb9i92aQUVyq/CXmBzUMgX41wiZ2y4tOR2jwenMPeFnTBzP4pBUhc7Rq9ioN4sFaZ1TV
qblvmA3+hLNR9cF8i2DGHzAKbMwSknIILbibKrnYnKKzxHoHuiOVTwODBROIcea024pG/mXzlbqK
EFkhX7LOzm6UjCK5+dok7tEXrZ6Z2PHPaXHx3JAlJkCTHUU+B9/ZyLI3N2j+qNzN5hHx3T8ok303
sxTAZOZr6XJ0yWfwvwVdbC4VzToKousVw0sQ+LhulhGwzFvynuneF7jegtks/BXqpUb69zB0pNut
SQeovwLBoD5H7/f510pUAsBMlq1JT1rR2ryT0w0YMszQp3OLotRUra3WUalWaz2VfgRVyTCQuRZ2
BeKTjxIdDgZGw3XEFp2EYB+SH1RUqwquNoBGe1ytfnQ2lhNIMeAYKlUrD707qVta3wjLQlPrT9j0
ji2sI+Rjeb2PrB1rDstISolUUkqp30pYRBC4VTSB7r3iWik93Nw28NLSgezydNZec4vrEasyeuC5
EUfDMTkXnE3OhwguFNtqsmxNcmZO7ptBK2/vVHcluYcMK8LfviylLOQ9uJ++K5s6ufs7ZVA19LlY
CGO3XpxW//q34IJR88Gg9KqHdAbIp0JCDh4BgpJomH0BlcDnw1qhKiCGZ+pjIr7dj7mSBDUE+tXG
kMXcWWUONlDFHePLok/+Pv/9zDVL0IcV1mgXApPUBIZaUlqTUuQKPhR4KVvEDp48WKtB+Qxd9vY9
RPdFy+eXI8j+t8b/Xyuu6Az9eDrlveA3BkYUeETQH5nU/K7Br1DmjEywg7LrA33ek6ak+6nkog3X
qdY2aVGiS9Q8luud33uu2MzlwXBbk/CUB1EFsWwb4Z2m0vLQFeuJ2MFZ/c8QPMJM8z9w+mSAKPVU
c9kv9X7KG5UqPZCKIURJP+wxE69uhjwIVEtRCzDEiWEn3/3YcUqF+lX8DBSK5PxiAFWhwGGz0ge0
QS8JAXoNg98EVzm+jZVS2/colgoyqe4TuBtyTI225VEQqTHL/pDdYSa/KEWOj5zGgHJvFIIyDh2H
4vxdhDyc1khXs01IXKzufo1dn5uW6OjC7FHTPqU16QcecYFMsQ5GbRHLOKLvu1xzLGEAG2r1wJJa
NnG+drHXdktmoLyw2BjmQGdDyuCeyD6SqaEjNLzfp3WS49XmHjeyXs+vPqZbbaCDZShRu0mkILYl
vvvpFuyevUxGmRGNp5ca4cQHIY5Ybq1z7+pQdbomQdaz33TPPRZrA3eyPHCtDjlmOsfIasizMjWG
UG0xBeEpfnn3vzQx58t6Rq/xgiwLksq+42Ks/2RXIAue9M8b0k3FCBaSobcu59sfeLYXp5ZjIsqg
z3k94W9KDy+7aPnNxdnV5rqtlsbb4W5g5hRLcvNmkulaJn7oUHAlEkWHcgxTs3V3hBoBmWnegkOf
xM6wShkSLgHf3X3o9N70m5bHueWzXuC4ppsN/Vp+uQs4VMLPGSaxybt3tuHOAi9MIABXqd9P/RC7
oKTKS1+4SHWE1ZbuF+SurEVhfRLYegWsj+FeDwB6iTAtg7/XyDh3E7QicRG6ceRiU/oAwIgygUgs
vQ1FzgWCWg84hc2bYTUwFSjzGaIqZPeZmQG3LYnz5VCA28Y5UpYlqxIjkAzAFZDiY/dJgo+TMYxN
/ZLES3xwU//FQfWul0WLlQ3aKkpsVZ10YAA9RdJo/MIFuCOXysAEBPbi+GvAJ8N5Dn+mgMxBXWGM
7FEfgi6yFWUvRv0GwEITLNFgV7yJZoB+qgRjZN/nTQlpuj3mz3Zfc5uArHBZqjJ2nDhw9fJAY8F/
oP0o45g+7cVnYdDvxVbeRsDq3vIeZb7r6v7NrwtUp0wjg5x3JT5eudH12SMaUTXvzxQlQYOt0hls
8GhVfVCKVGEJhNO2mcpF59Repr05cstOEuXiKEslHGQnzFXdZlCmLS88+zIpcRiBby69YNlzCi+i
CbaKO2wlCAk949JWC9KKpmVPe2eAyQYogkJcWj2BeqdGf2eFNlPd7NRnakV61rljEp4l5mN5z4EZ
1CyudjZfHBJWAreMM4j0qAc0x/uCt9X9ggcREJcsXIQ49vubHKdMwtD4HfzbiHNHl8eBh1hIEV/d
ca4NZIw16cwaMaZzxqGXLNGNZ80D4G18E+yGwZrMP0k/CokzCzVyb3lI8n4wZ+KaXIaBdXf3rldt
dMjaGJcauP2EhHg2IuaD+h9hk5X8zwJJWVI9fHwEkYh+f9guUjN5kF8iSospA4nlfM6KEjkgEbp7
v3N7SN0A0K7257ynBlkrvNlGWreHphqgkNcOAVmjRicXZ9z8pW/hHQUMPTSAtot6BS8S3QpMKcUI
nOJ2iv620iYZb83wsqaF2fOJajUY591mTz2Pdyq7QcNOkp3lS8RAXp6jSh+Yx99m7dBHQZ4HHH7G
uG73F0EaVoKH1N8fMZGn5xipWdNpFQqkKdmvmUzKBibIN36ADkRvxszKJDBjsjwzXc4yWjQ7Fprt
0U33nEXW2L1U0Iz74J7qOUuh3T1rmfGhtt/hfYgX4HCToTGV/4YM9nhFgo3aiYtvG9Oe3VSYtoMr
UHEdGuaPeAl6cw86rOfVaimyRkU9SlOgB655oY/h3oJbr9bPQbXe7xYSpK+yL4AGSN8DI7mXap9+
YfNpSZoPYxH4ziWmjmxcJntSSyMWFJU8j4P197Q4oxWKgd2fPcOy/w65b3T/esM1nysY4FTOaeOn
dWxE/Hpk1iMPkPrEjvJQquI1SWLyqpk2VNMspPcZkqyCymvoFYaZxlxu1xh0WJJQkpWKIPWosw3c
SwGQ56BP4F/AG46XQCHRw+lID6jVWUpP+zT1yTCVQH/eiFT44s5hh5X8VB9PIFfAnfGu2dcoPDNp
ACl41cHwJvQwAfr2pawEjGzGV1sfdyHSmxmJsqSuajAMcGCmkjkCqHKOv2Qf51lTF2VjLQWfzu4x
VDGBv/Kq4XHVZpyGkRbZ/G0UJ9NAYiOfHzBocmfXgMLe1iHcF5qWEZVScDK+bs9lGbrzpleW0qac
WxAEOkbaYgEXPaL33H3vu6jaFpMhnKbqWt7Xqz1PKioFc73tRUdhVisK8diWPkadDLciqpzxHv6h
Ci3pODrbtT8qASaAegQvAJ3ywjAEQTQZTj6Lz96ITucSgwt+5LSuuYTsPojX3GDHKz/SWtE78AnR
PkbCwK4kKBMBwoNhNRNT75kahljL7tpEB+LcEiYOxjOA8EeZySCiWUEkGpl/cAk4znrZ7jDY8PwI
CbypIPSm6aVOYqJV7jd+7S16b1Z4uk4RCeA2Xx+VCaI9C2Fe1COKy7VbocfRVbxpsLjDwEmR5J1O
GdnfThtOnU8yGKWpiM/IifaF4zYAM1X1Wu3+Bo9NCSKVkzr0PQsZT58yp01lLnSdXnIJKP+jvMMo
brzBLWyApjGlobrXkiO0iGPbCn3jRrplFlIY/xfyFfN+tFbiF2LlkRHGrQekF4BXNShUSnzLkYi7
QMX4n6UW4DKDqK1NAS9cNGHAXYhiMjoZPdiKRCsTA0peLh8LlhLPMu230EZkTJE9iMYxRJq4v+F0
5PonbQN9/ydk8vHo5mGTap4M/d2CpEIpy1ZnTivJSXXKdrFoD8/eIw4WmGjPEY+dk6xXX1KR6s64
8ftDdJjRnVHsmI+6DBsKkQnqYgPbtjYb2XyVy8i60hiQpJG32rLuQuYM35q2uYk266v7edX8hjjh
xEVT4gzLooGEiz+jHgXAXox2739p49/XtycFzKDisO8Nt2RQ2cava3e8HalXBTbFbVKFREhzfG1N
Daphygx+waVEaZpfGcmVpG1Q8y+uNAxAuZboRfmoW2VEWI1bnuDMiAXAPHzlxt3mf97Jk7Jv0+f7
XX0/xs9Lth6TtDuS/2U1+5uHbfRABBcrmbZ1gOotRpLYKUOtdi3fQj9UsMwJYUm/acOlRBnrj/Q8
5x+grZTP3/9cemYurhCHntHYZKp0gzfGs6cPkd1uQTr56Tt0jI3d4D7J5J33/jSHRjcrTY+J5lI6
k20K6oief4Kln0WGxGwphHlKxjanby8TtKhFMtNzc0uS62eoWFztIepLa5IcpACNqjIHzF6MsMaQ
taFIVt4CoCzF9erD4hjQhS8xshjar3mys/l3ycsGLzR1e6VOEPgXM2BVeoK/pEK0GuKw2amgbKV4
/0gbMxcBjaO6yo0/E51DWF2XJc7a2N8a3b/wARA68hGkNJAkdtqDI5lDrGhLzvOwxYl8ShGnsyCo
oZnzkzB1uKgl8lYbe9lRmPNFz7nWOE6CS8dIrzBQ1IMXnVSsDOrC/ZcofKYlE6w7zzVp/PQYv+83
+Azp/GtEoy/piDaZDoOSKL8tt5P50ZFWa0Db9llwJFK2HABo6WbrU6O88Vda2svNgMtmiPgsN41+
Z9ARSxsztc2zi3ToN0wQo6zwi8T2Kra6honJg0XVYu6jALwgHBAVGBa21/0FJBrU30oEGXMWXaEe
BbvYbDNExgPfIFntrasdJ3uXWgzZfU+lSzdIj5mJwJl9+ZCPiLLLvTap4ViT1ck7B/PJlyTvH6L/
oPo5vkECRQJ75FV9rgxTSGuICH28C5tBt1i79yIcXdbYwbYreW8OeIP8frKVzFVzufzJ4oqt78ZF
o0NSwQZ/j2WEZx2OQJi1UC6oOTQB6j8++tGTW06YHH6a+IJE/d0kWojNxH9WYm3HmzM3C4kOYZzr
Yfrhcs1tbXVmvk0ATPJGat+8MAygAOtxcPHhfKtO+82uMLDkDWPT/0lQlzQI4wVkubMmYbV3LUXz
fHADrR85F2Hkz1MAVsZSaxLWT0IiRI4qlWFFqgDAeqVYjBJ4NMOa7MdteD6kuaEnY5OqdGMwM0wh
7sg2uYurqs4j+o16MmTUMvYvRJENy+aY5sjbE8t/X7RwmY7nSWzgNG7SNO8kPoRzvsmN/SSCvocV
9/rLAqFZ2nZweo2qGYkkcQeozvMCLKN5z35Mrti+C7mxp21qXe8XBVGZSh1+d+18O6wsJKoYHbs+
Le5AJnMOEqhIdifibgB+xrzx8EWWMCcKy2u/vaJf0lEbc3GMdezJuz7ixGLZ/xLAmY4KiIZOOADx
Nu0ZNVsKELtR+52OBDdUixT3bX5ljf1Sjc2YS9wL1hzmKmRFgfEQsaVqiV88AIV+0K8m6p8MFdcV
nngYJg04EbwWsKpFUTnhbM3BIA9rcr/4GdsirikFTmpaJ/eB1uQG1t1fjsoknX3g5Bm3V5J9dt7Y
aRBPqqQeOj9Trp/DcZjOCwCaAK0qRX+53axgApWK906+/qaw2ydTn4/Z9RjYeKu+l13qwoPGbVMM
EG26ZLMtDmp28dPsmMlHv1lhq2fSD1FCeyI47LLahBtdy45nkvDQC8t/MdICRiZ8j9W443JgFSCI
Sq6CcfIpNuAuf8r87w4f2jr1T+EQVNfxfdXfscpByXtkFStTOmtcHKeb1Efknz846pcp0ZWJafkL
WZXUon5bEMZsOQfvKku6shBFWl1dTcwB5LpDSlewf5s4iqTMw/2VJGbw9kMi9V5jvv+LLCS6D9wQ
d+bKFvz5tuxou6Rwu7Zx6rkxSTzkp9eJL617JbBDT1J9ZESgravsRKknJv5brt6zdGz+h09Ch+bn
HGCVJM2W1+AYhi2MaE4aANDqtOk5yXAL2tTofmdUvh7uQOgttmMJG06TOxpqIoizGGYBx58meCsy
lCX9WSYRpo+95KWdG8sKZ0+Jgc1kFPvSLzDHJo1MeSTO4rpNTX1iDqsTlzdEoF8FsqjYuCw5Vl8K
+3pQqOe8G1YXVQHgnUW0RDtnrhyM4ij4jf8zDw/YCVx3lf0FkvK+kjHXiq7Xsuhdavtk2TPa2h5w
hMladjxILZo8bAWg/Q4iCWxOwpSiSkr4OQixfPF3qDBpqYkUfacjO9INyRG8hoel1RGBnjFMv83H
ZPYKkfPEyZM4dGIvAo/57LWHsMhsfYDBXn7KIfLmW9rcRoGm2/+1NWlBy10MPDB34p7CdXsoEEEM
aBVQ9zM+RVTtcKgIkbfNKTPqcUtkGwJv9tpPQlEd4bnEGAU58IM9XQDWAAs8mrBDlpm+R7z3U14y
glxZCiUCeiqA48Jji8D7b+9FhinRK1ijk1Qnc7U5Ubm/2MQfckmhF0p9hXXB0/hCcvv4dvvQdprI
ovJBLtSUyzS56L40ptpHymeO3w9BYCWEcLVexQw8qsqZnhxRINVMEcRtJRkx/8KEKjtme4DXq+l0
Xt48+QIwiyr+6fKF5OKVDllLLAsmpb0hCPL0evcauXt9Ltq2f5xGC42uAkyq9ggN1R+ZuRQJBjfO
kb27XKyx1vUgqiFqzMLYAEMeXOZSltc6UpJA3vTzuYrOoaQQ22OcR2VhlZyEK+7ck68DmMq694aq
F3a/y3nSJLsEQBEFiJ/TKZwFf77QEaPa/54rjw6oRbkRvPPmCySq/VS1NrT44XwMyQt+faeqZHd3
Iotm8yr8I6v45Imsxx9CG0GjZubNr6XnMV00S5VI87kuZ6iFk/Oibtvr1ndTsIEPgUHE+cfwIy0U
dH3WUeuzsYbEFRz7bZ5TD4Jqpm+8IwO0awDWUIgWyPx7wODijmcQ2+aHChj6X4j2OSItfp0xJVWK
+vJPe4JJiAky/qz2vlRXVCmhNYXkaTtp+ka9m5naEaprUgXfwVyCXwQ6WPBwRIDKTptLa6ibA0u1
ANTNNanVH1ZD/lmR0Jhfv/xpDSDAgV7L7TxSzccvSG8b+Xsd0TGNxuzCq/Fq6rrYeDXMpd1d4mtM
AwNAq92pY2Qi2cs8WmspFi2dbUUBuY2hAHGjG2FZ0SouNniYQCM4wBNwB4XHbOW/zur/SJZuKlc0
LKoQ1ZuAqN948vZHrk0k3ceOsKpxqxFQrWf8+GTXvwVRbRB+1/NU+/fx3vGMqLXqB+1ilzDkGeSZ
/Qi4MFfTQBXJdU0vD6zUj16sKuFHx4Lh3TcWvqpT6JRDS6EKB7mGKnIjKbXC610nkpj0SQykypXX
ObrZ3f1T1lZeSH0+SNEY2AkhNl6nMi8M4GmwdM9o22z8t2oHPzC8toCbBj0P7eV7tzeBnZFD+uHN
Qe+GdphiNNWTO+gHZqkx1llAbFCMWKTtLJXggW6towGIFehjCVjBcbajFbsbpKTdccwk5TlKDNpe
QI9Z6LqNCJLf30JpZkGvMfSdqSHJjqvzktBHY5J1ybsnIMJm4bEudTuRUZEnad7WgIORhFODGZ7T
df+xIM1dvy97+OM7QCt6vgElFbdNi4zMtVXVQ3mzdQ+53RVwlsreF+0jxIM0RPUxCciml8KF+Cix
VcUg1XhAInejC7cgSMDVeW93Zx29vjLMkyhpzqTL2wqIznLJj+IMYPCuZcNFQLsNa661AY+V4z3o
+WTEjAuBm+DVtIQjmprbp9Ap4YUddtyLEhagXmJwV06kgeuXvYC8AX8vKQ6uKthyQi3ynkedaMvP
3X5tDLGL1lpwJiLTCOXL+J9x9lAwUfrarEvcJ1GL5Lrds7wfsgRRIsEWJvGxqp0qb0P5IRKigbAx
CyVi6QxZOMphGZJaBe09NGV47tzxr97ePVfSyzf1w53lQ++FyTnUo/WmTXbf47oc70vv9kP8HOyP
bhYEBaXzjwYn2c7IyDGRdqHfIWffBZ05KAaTw+Nyy65KA4UChr23diOsx/qXwgo82MSUp1hilkuH
LJgAp8Xqn1ULQdZhSHxG8w+Z1vSGdEJ+rNFv09lZe+A9hZQOkTsDP1dn+JE4d2S+IdCzTUDvDuJY
HQF2zc0Lwbp2Xn3BRzjc+zxqrUkM/7wSuCG/M3xw2FHMD2/RkX8fC6W1rSbJOicKfy5nX3DjLMzQ
S/xaZmYtsz1ha+wIR9+QYRWl8an3VFnApPCElQke9LCcEkHTKGmeas3GCiNbC3/4l/7LKtQps8UM
2jpnCqLqn+w8sQCjWcIlvvuCLYsV/f/Rm/NOfh4kkSlhl5+az1zTUfodPp0/d3xRGAKsLlkcPuxf
rJTO6hzOE4Ur1OIhB164/ofYGiuNdrEWGCvGC1IYmHaOaCQH4uxIDRl2/pxCXY8IVwRv7FM9ukPg
5/dufWS9yfleeThTPp8B8z/iLdNpOS0zeDTezxenbGjOA/gONNo33u1n/Ab1bBcyvHhkOIiu6o6p
zSy2Ngv+Izxm0mSrkJPq/XLYPQuJliV+BGi3szAaSoiviLczGpHc2CqYueJY/IJbxUx/AbTPMkgP
xfOtxlsmnmlBaLLaSb0ghscj6DoIIOj43GikxaZpEdWBRqzFqhI0UqU7g6xZOc2yz7TCmaVpSvF/
mNN9jSlHkzdCbgJsCwmpe6x8FNVxJyNpKORFKqgCu40r8vO87F+7zbdsTf41Sqtv8ZAYmzs1n0aU
Y5ch7FAbRSxk70OaNRv8D18L0cTRzVAnyWxKElAzn4rH2duhJzus/HVYKOlvTWd8Rzt5bJZn3cLS
TTZ94EoI08Gb5DARthENbPCsE6cg97kDyU02vWWDo9LAD5J3TDA3W3BGGdvpeIGewLmpJgCSwhMg
ojieEzjprozAEAcOOUsz4qM9z4C/QAdwYoMfuU/M7wrmPrZsZaX+QKMmB2x4fdxR+RgCFhDhuPh7
LovpHy3ZZEdomr5mAm3ENPgMrgx1Y01W9LFwDfXyMaWINlyAvY1uJ1DHPEGczFsMJkPJEjiSzass
b+sItF6aoaFrVVjqOUo40RDIJSfrzFeVmFvmzHBQgF2/YuV0+6Lw6t0eVjUR72q56o66jsiPC25M
rIGjuiUQCCVfbDih+MbmKRe/XK22iQJUT6yB2nXL94XH3CtN6D62dJrEQLLLrPUwJ3l5vl9JpmoB
TAeP1XrYGQFkARJHOUJJOsUR90tZoIiwIHSzirM8EDca8Bp+WRkDh3dpNWAcNGoUwxtiid6+nb4/
XDsOCInIhGSTif3a6w58fmFea5maGgLRWydGthF+5os0bPkgURdEv4kBnpRWkPq+zZv0m0GEL6r5
ju9ewG0LdjPl0ETW6iAOlPNB3hCLo7TMULtZLqV1Mr89bQPggEd+UQ9Z153DmzU+j5VrPxpPJ/be
BS8toCBs+RgditQEo/ot+U+qtnSIAYTAsi6BH1hinfdMufThimASKYsvRwPOasTwhsEkDAHm8GqF
Y+5YA4daPZri8qfNLWGJAethMCz4FGBV1zdmqsvyF9sAyw8JkyP9N3GSn915+2iLtYKQdeXTIvyg
HZVF71lfo8ozLQdw+kXHSd44rViNYzFrffuPnezO6rBuy1VIA231wCebmpzIQiwWyn8m03V+A8uh
inPJZsnkcNexuPCTQYtV6Yto8oRxk8TRFza//FebqiPf9rzSHd/ZkoVYCsDhZssXkwke5hF0/Kqr
ebaSaGNJpiR+ROlqr6SgEd3/O+aD1lX0AE8JI1RY3ebBWC8nkE0s2bEKUNWKBqX5YaVouZ5Il/BJ
qKzZWpWQvHrAVJTYSEJUy93nx32fFkg5sRrYHv45apastXnpc53R7ErRrAVqAm2MdHwfvaVRhMof
OZYHNxr/7DVIvR0ztBQ0dKHG9Kagbx6xRgiIgaKd0TTW539XoJi5US4h54iZKSipBs4sjp3p84+g
lAr073O4oQmgAsKVoECaP9ypMdnkFMfHNdklFvb3/CnJPxxlqsjl87FAc7Ye/wwNBdmR/PaWgw+K
oBZMYCzXG5oIGvtBqSoBSZwYdOLTLJOj2T9XAZv90z6CiIlDUgnGpwCiIAqpCtdvkdHal9hCqUNe
mDjzENtINMSuDopazBjGpaFl9AkJTpn5eYRfwS8aBayRN5MJPiTfPk2+vaA8a7pDSE84F0tGFOok
tXuRALp6jvlGkDSNRznsQQ6c5tX9f4hfw87yKr2aI5P7SpSd+qU5wyn3Pu/dHMm2LE9jsDGy1s6r
L295XM3fMmuxjgnGTsnv0aozoYjDqdJLYW1oeHN3FH8onoCmLr8ftUPw4nP2bbQYYdaZBkRBV7S1
FnVtuztWbrsDPXRdowTnplbTb861gnBd9vYacV9zbVswnTOlK+oyCcRVJ3U+u5oQVQJr94K5rDYv
kpJEBV33YiDhYlD8KR+lQuWo80WDumQM/xL0a02rCoYrwomsF2RfeW7uVqs1Xt1WZZQZK1UyZyCf
BIHeDw3x1Eoe2viISHFnrpgclhyFwkx4n/YCo2ZggVQ+RfoYXBIig//Qc3jutthSdeoVQ6KLaaws
5MRusFU1g4HnZcMvJrZU05zxkoZ0O23SeEW0H/jYSUsCmcKNj+Y7mLkmgJy8TGDtOcdAn0k+Ndtd
dK47Y4Azf22uctq5Nx0EcDLEF+4wEI96p4D+Eh/bZP5InJbDkVGbfUXUwLfvlH09f4ZrWvfS/tkr
YUH4SycflqYWjzBd4qRCJtKNIePtgLYL4HdK+o2vmTuPtdt0pwFb2h71Rm4/MJt4A3hS3gDxLS7O
5BG06AmGCQmBGoHqvrZpR/NmVriWvRhR74u5H1elNEbX3AyiAlX7AejqKfrYHDqx8QLBHcxcKn5m
cXsSC9/AhMxMkEzBsM+aqtBsRwMrHzHEQjbj12SDH+9N7hjmdYvFkdsLXNUEOWNevlILDchk6BrY
CXuiqkFcojMGN0w+uVrIZtd4ZVXjSUSE+WCZEmFaUc4HGAKTohFA6mOyRemqgLA7O9u6eWILlkgn
YwGWLXDQzvm3JRxPf+/iZsCjfX40DZ1VcwJKStCyVhjoBol5oqxgB+neFqbYeN7sMuZM5dOLAuUu
1yAVylaHByKYM7/kVbucPMNKnZFemAwRSDs92M7DxADH2mwSHRLiG1VRbdxoCs9N+GBseGCUVsTD
Fg6HRlTtM24sGhhNLZNrV0RMPjUbko7ltUaf4RCZsiI31OmrNeA6uVcB15ACw/mmgixUY00+V+1m
qspdU5Ujis+JG5wACU1aWIFjTOq60DOFFHmG14q4f90CrQiKPDmq+ExRY6wd5lhW1RiyCCkwZDZq
YlBwK+aNYhVN773utHabt2S++ZsTE1UVriZfCMDJg1IzpHE7NmehxuPZNbCwLe9tLZHjh3rhOuBF
QvoO+maePX6I1bA2C361l3YiOo8o474LJX21GeSAo1UDxKV7Xqx03egRWjPXEvHiIY/6jfeC0l+b
t6bbr0y/3r9EA8T6gfz2jRF2715J2Hzn7Q/g0V4aRh+/DZfGptJgU112FUYKJoMTHRdijdLl9vCK
pyn9yHkGkVKBIeP/Pg2twmWtl2EDCbdckAAgnZN86ONBYdja2f/J/m6SWpl6JsgcFgXtjYsOeRF0
rSq7HZbJIt/MsRS2cz04i527pinU+bwyJkPWaoAdMEFhbgEqwFE54HwiM2ADkgb3n4YzvsnhJ932
nDbkmIVOfvKomXrL5xGfVu2L1EeEwLcSZY4GAMD/TF97cJvdhzoIjpExDjinMrb3i158KpabEkOV
JEjrcB6WlRhIcS2DfZFTKC3rulSmcjhFZgaGJLxQqUQyt0A3RL+kOs+Nu6zEWm58dax0Ob9u97TT
rJVnTI6XafPTUTaedaDrZ7M2MKWmqF0a4m6kDYzc8NtWXNhJCRf56bH1xjGl4kpf3vJl90s4xbkm
n34N8aF0nzdP9/fmD71SCEANnmDLTQj3QvP3Y6iVP7OUKvuXTigBG6bn/bdCceA1Xq3Zq/INJQ7d
85wvjPKMpRuDmu6jPtXohJ+4MR7teZs3/YA+3L4gJCVnZvOAxJdaXCl2G6fmpVeihrfljOU3GorH
Dh4DUgr3Gg1VrxnzRw6M/BYMcZKMSD0KPb+tGA52TBT8jjfDThX6DKEw2n9CRcmp2ERfCOsA6nW7
ik/WHL4JMqhl9pX0mP0bQMLhK/8jCK7Uw22NAKbfH4l9L+QgV7BvXxPLH2rmcovLahotQmjqZeQx
OCoOPfssn+Dqs8OXVgDSyU9oDcr3hQybktA/4cCmbT6Ne49M1nHd0rfOK6xcS3aAVWRjAehAXO2G
X9yk3AYgL3LM0fIIfKnSvNQUncy3vT7VrS2kCcVt/FCEhuhbLLTdoUOdiR9FqpHQrIKIV1jkNjyV
1tPOY54qGnbXwnwEPjIYNgk4/Dp8hjbzU82rwQ4ccokw+o4o+zyEnlcHoHZk7CiEmpdNmZzv6NXS
s6kdTt9Xfe1qs2oS37IfXjZXzgGLdeqd7swciUO5uyGQNBLZif7C/oUHHmQhtql2I0C5wu2EYce8
/8uoI2wpZvaDqfrYyxfesIP0+NBnFBujUlhic5FQqwh+ImxrtgbGljzQYDDnbgKxBBHXCoTTIrOg
tGEaA8y3rIIsQvzcbFzJVpjil4MzqRk8b4DgvZSkotc8hMuL2AQo11ZkJFRnqZ0opRdUt9gxkOkN
Z9ZNLq7HbqS79D+0PuVeZygc3x2JTiqDt6X9UTXBr3x6ZODQ47sMiRkIUUf0S1Xv/XZsCWcUYoRw
KuJqKrJHkwDzSJclLCFcjVQ9PG/ZmAOM1WGPIaqpxIk5+ox+14xVPHTTup696OGbWhTozzRGgB25
L/TSjQkwPuFsz5OUEQ8zObwWICb6B2GHSKCRJWaWCIqh4Ur2+pWlSNO+13uGCD7sd0LFN0JWDAwo
2qpWE9Efch4rnzFYwHl+5KQxWICTQNHZUxIH8yG8YZoZTIWW5baMgOkVnRrM5b8AWIvqsTt402EJ
CJOjMgd3D2TbwpdGUOKH8Djregv/SKMxpgr3GF5Vda6mHI/ICgX4GdDwe9KHQWN8EsIbYhMKz96M
5XJH0Ofly+vrK9ZHhtbZlGXcppbwtuuYAmWRMDGr5fyiUuo+zLyB/09KIkg6eW5hTo16nONhVF+y
5WhCsnpcJ2MKgT/7y/u5mFRa+4ovMqTXC8kqODGelKU7HQG5RH2RKXbFeO26w4YiSljRVxkgQzMW
6vHhkvI+Ymbuy3mPwgetKCIHpsMaOxcC2+KI3QbqF0+rjHncu0t3bZn20MjzFiQQoR9rTDldqjPi
YxJ2KF5U+sGjkY1N+m6AYaYJH6tM+QxaBsWkmwf78kNyRp2E0ShoyArzUzIDac8Yc3lTH/7WxvOm
8cRFxzqW49Ld+KuafQvpJkVX5n5o2FkaOE4R60m5b6GVyk4nsttMpGFKoOnwX/cpAKckjwqilDwj
RSIx0MigYvPK8pRTNZHZ7TG9Ul0KP6lYMvkPZ9QmTAr4/rN/RJAHyFcoJxVeEHiK7XTygNZpKBD+
TmKXnvvyqqj1UYxY/bc+Hh6SEzOvwQ36pu5mElHX93zY6c9SIBsOGbBoGB7A43+8AEPQGH8/Xaj/
WddHM9gk4xbHg8mxGsBFKNrT0L7rnbMMAflS7KKv4NqZaib5ig0bBLz0rmphfHQj16eGOtVFc/wi
MApqE3iB9Rr12KZDHKOneHdW7IUb1iufKFcRHAdreRfQYgjD+Eb/IiwGkQBX1wUaPSXhWZSkFQVs
qXZW1Hd+zDxSLUUZQILlGeG2Bf1yLeJ8FJ2Yh/KK1xDwxTcO7y341RQZYyxsCEQvJrqq+JcGjuMK
dn7uVQROv6caJqsghNVxQjDBB6yL2uCrTewxJIvPZzNSlMNmK5bENerdKowcBp8PJq/+tzrkBFYF
o5IIxdFFmlWQuHbBSOC3xbVtY12ehMYei05RUkBxjjfE2MSkZ6V7dj1nbbqyvpjHL67kc/IZEDHx
xm3M1JF4Sd2eMPc3ABVgunnLxub8/cDZvE+EJTFs1nSs7NQ4+tTpIHKPMIUUxCjWvV3HMYt3sHQs
myNqw3KGVPQ7ZlY3M81IR7aomdv0vApeQd5hy19eJFpdOlAW/Zj9Ge1Ae5qhsDmyQpko5LvZPRC7
B5mCjZn9hPBzE9+eEEU37SGGuYlBf6qlO5odzeAfCGqPSHOqPj0+xQiu21Rzy+O3bRI/MHjzdNXe
3QdsKTJ20F7vxpXa15mzwwmGa56qSqSBBaO1NjfvppCb2KJErWxI2r8MoHOfIkC41hxNf5ElwKn9
Iza9iCRjjP89Oqt79v5wOPIN1qOnIEnP8HiFHSnOmw4VjN3+TNBKAJDGdTUSHcWqSZjmw1dTmsjr
/pe0WvIWGnzw0RfJxmMpC/G+IfTyGk0oWqvDieKwtULlEC7R8gdu+8P+JaoLNFFi75g8HCEmJzCf
rY/O+ao0QdYAA2PXN7U3eFOdRurhIoJ630t3B9PqMD5WQuMv3eYF7IFOYrsJlo8Le7qCZMlENa/v
aT54CKL3y9emYz92WUuivZh00Nayq/dd1p5PztPsWn+5KguwpoZZtcqk5UKfxTSNn36ND04soQzk
Tfns7NlFHaBJgDhxhpGjlOZ7nXAeRK4mLjm5YaMm3brhPDt2uhb13kfJg/Vyc0DBRD0G/gzPIj7a
SFJhojPROOWQuTkXaAfvnQkV/oJstdxhCp9hhw04Rc4NS3tzJfjH7u5eQTAfdhFbHbk7J/W4cruT
vtcSyVF78QemEIC3r0vkBt0bN5/ABoueoDwYZd2NmGNd5oRD1Io5gAnRdtK4jcsHbXBeDCAWuuHn
mbXu8QLbipqiUPww2fJSS1sR9Svli6FwjlaWxuA6kKMRBOKB/3d1MVP0/fgQU3BGmxiTKbNwBiwx
CR0lQv9NQs9uFiPdlNtwZKrEz4A9W5+UN/VbC3o2uxP1ue52sWWsEkEhlz66A786r8wlG8+CMSiz
RwlRSTa3d2JSRlWbPfSrse8MwFaekUUL8+6qgYh0LQFVxqe/n2uh43iSurSliBus+bb0xH3KcDgc
QrUbo5y31Vh1YMZ/bdcJXFh1GRVJfrQTnF9CJBDkbfp3dkUHk4K+e4lghCaOVGaud7VOJjoO25oB
qmVvb7RzwljOn67xHFMLlGtSGxajU1f29JhyxGWqiWEBZPP4FRPLpWAGXFO9uf4d3n8IpoJViSI7
c+SNgfqQQhPvvnoEFUTI4MHvWXmvnI3rY8PJ2K6OKjLpvYfR+jOp2yMeiuQ6UjDJsBkweu6GQ0VQ
PhafjQfod/Cci1bISIMp4RsHWXUmdA/MGzzGujcU6kEhUum8GWkQsrGmKX/z5eE949E6WeywrJew
OqlMIwVBZNBFvecb/RFishVk3Oyj3y2pMJtX5rr3sW0fiuocLV0hPvpmWRKRi8jFyVQqbSu+QSwm
ipE8m3aOSDVeBEBp9q/hTktlYt8a1QpPSKqYboOWecF3bMAvE3zkqpzjYeyTlGTmmZCSwRQ1aV/G
miZf6+dDhblCCfcP8s2OnRdtLfYapn7KpxwkN+JndeMMgngaacDcb5EMeaiNlrXAPhFWOCJ76fNX
GCYcZo0DwJvMqVKVHIHKmxrBU9khTS8gwvTvmkHc/pb5fg0yQ81oipAo1a8ChxONOJNLjdkPj/Ez
rPlCVuWsCWmWpacPBdXxiskH8St/H5yIX3H3EqnLAi6KNep8QNTSwtls4l3YoR5caZGy9b3QLMvh
WNlV4P9Y6uFlOGeLv7iuArNxviGiUropNxeKhz5nUqixfC+4+7sDj2qdpz37kCHtGQZbfMiVT3Ga
153j9O2s9QsW2B790qjFyiaJamfnrhSD4nbzM0KbuQNxDFX+cdmw6x4eLQEYXLN2grSZST8aI4US
QJVpDNTYAT3jmFufzHfsMnjfJhR8xeiP1cGsaz6jvup9cpitnNMlouBxzkQ8mbNmAPmHoFdMgLNT
U47gGmxaAaqa4YZePqPpqSWKxeGtTNHitL74Yx8smA5rssyqcXurCwEJBFxW3AwleaycRR7sMMxM
kzFBy88XaGSJMHsxlwwjazjAxfrAN76tiwA+c0NerLkNe7kp+cjF17jUP5H0MOnOrr53sIZjZqJP
EGRHMxY2YeBas3nVeGaYcXcFYVRcXo9Sj7gLunWB+ltNJpMNjEK+xMxt5OjXb6ep8LAam/nyyBPl
LaHWBM6agj+Ps7Ko/06qYK4LbbP/ybzEERGzf+FkaISTZy0CAe04HBVhJ9fGNXqbThzjSckg0O+H
C52/n9VtIKKFxHIYduVzY2RRNdlL+bXHk6xfsgi9+df4vjQYYtDdUQSUzHO+1+NGW23Wdriysp75
X+SfrQY0R0114YdeMvwoHmFXhPBzB++MDUN5OfZ6S4fRIaxkZxzVVkqc9AoQ2drciSK6GUpnb9Dy
gx3Klww1BtnpxIf4qLFrg9yF2JxBX8Y8GrrhTjjGh3GnpSvPvYxiqm6DeqoaIXUaavYtFVw7/e6N
9aOw8TntpeF4bDfz0EiwAF0ZcOkjNICun2cO/W5a/t8EnFQ/nFUh1opYwY1DN7EM0xFjLykz8xJP
HcM0m0W3uNMxVSQYVMVO5tEpNq4adKytb8p9qrw17pxE2NLK6ntrYPI9lsZ2dCMMI/3HjyTmhIjT
HxYmSNc2B2/QOV9DrOn3IUWSZCVr3/9+PH7Nek06vWGOqNXspwuAw3rTYsUiUYpR2XQOxjnpd2Yk
qTsfxUbrbOvH9KtFHRd8nzvGJ9uS+bZNaBk6vXNFJSc4ASYZy2wyG4eSqgCjv+ApTwbqXeTnflHo
TN5iT9FGyN6P9dtrgoaIqCWDocXEKIxPqsgnh9Jy6s7nCipIWctT1kMHFanVqGhQtLT4JSxKqu3U
ClMC6olyshZs/RTPpteOvStYDbjwh1vjtmq4ytruI5Jz93BkfMwvudIU2pm4eoDDb4aTjfHO24u3
w0ij/3u8TgEK7eMWpqX/yni/hiNaKYwR5tNQQOQujbXQV1FPQH5h5qf0BWNue181JoOK8LmdIjM5
lkN0ybNDp+qkwFcMYbnGE/r6WJ1rKdJ2wPqF5QYFOtlc5ODcTIzTKMwtzYXyATNiqCWBCXMLHP1g
mBUryYHtvfdrk3pMnKCSYjPR2Z5tVvCkwl3OBrBSnuyBfxjqAEMSucv3lC9ncTx2a0jZRKF4iItE
EzMy6L6s2aATjoJWmKUOBC3pNzBrZ2z1pPZhxrA022mqJUiaJHkusn8wpfOXHPxqTTRVqkxOKq/n
Fgv3TNdWaAg3MelJWJbisJrLMspIuvWPWxjNcFUtysOm1fSV0zWi6yeFb1oNXhOmefazOXsp8HJa
97jLsBLhjF48avLcnbWPj6BxKPyigXLP90z5b37C9EqYrb+/mJx2mBZPBshiUAFHezKpET9OSri0
WWGw4ZBWCOtKRV/znAhja60XaWW/f69Czczc4ejiIEhuphocDlLMXHjogK/bmVuaDpwwTokU4MIE
PfgtBMBLoH/cuobejxnK6loLNVVhR0t3o94MhCN5EfrOTREQpNo3+38lzi0xUVqHEHN3mBryv5uL
q2mOcNhWwF20xxszC4pgaq/7Y9eUIRCPF/cYVgnJIiFNdR7sbzo5f8qUilp/540LKolupLfvRNKl
40p/m8PKbAHst9isOS+zDEAUKT+XFmpBjxXBwU6+MWoU7HRqtSd5U6QTkNAJt9yhqR6yKT/caNiG
Uw3hSWluw84f+cxSxFhS1g7EsQrjP/wqx8bfGWc3GiVRX8faebO0ZHwUf895zwwVV3KRlGk5S0A+
tZMuvTrhuEvP+CImUUSQUJ0BZ7EAxoudhiIp7rG07etA0nNkF3L5WmtzYrjeeDekG1N1ey3O28yy
pSB/ugh2MFYTuvvm8/0FJD8Cmcdmu8O7/6XFdK1WxrDidVnd62EDdJ15OSApqGB0sJW5iqDv8rmS
qYo7q90ulFjrMwniEAlGOIKo9SjlrBvdzX1XeBV0iDeHN378SR76OlAlE7IIHPLF+wGIUZNctdF6
Ej5Zq6618JcIChpbFI6qbKcsiDlUGxuAt87fzEhWYiPmHr5NybA5T80W9Mf2nQKZBU9pkLGOJE3C
KUNt9oj9J39HmLxE5YDXMe0Tb065CQaSr77FlyLkBB7+NCRcJl08HP3XeySjD6CKtflmJ7KpK1Z/
8jiUYlMv4kmEo72w1Ef07stIy6bHJFZDn+QAmKqmNP9/Vog4IEXin6M7Vu2la8pGjajp0yZI2rtf
CZwR5/SnzboH5eG26TS4cNpsczCL0YY/cvOxxteg6jro/f0p/xMJJb2+SFVvxH23b5itv6YJNlRo
/PkiKtDgLapx4IOwlAaJMRLPXf91d3sekRORnFuLUYcrJx02gSRwCORsjPg4ix25RrB4KA+pc8Rc
B0vTf6fe1Ps2A+8rTprUHGZUAky4V2zWA69vVMaKsAQ00QsS6egsrFgvj7//ukUENl6+YEC0CI7X
KNprF1ZbtqTRySAnjo24EmONf8L8PS3Dyh1gJnCpYzYrm8mwF+13YmbBMF5CXsnXNNXaXdPA5wFt
m2a+fHysmMpb/GPGz1kQccMlWdylXGPNcIWOa3EMwOoK0syHTSGsEaTC42wZVUtYY17DKIsVkmTQ
lp3zdQIolc/yR5g/ns/fWeQ1o7+Iz5drUddeJvOt+NDY2M8N5MZDGyiYgzPQapK879ItBgz/T32D
PnXnNTdBln8ItHQJrHCVYpFJN3ZpElwm6jqFyBV8xBtlZMzmgeQKhfQ65o6SHx9/2aBj0Xo/vJvs
nmW0enTOK2Be8rP9VCsXwTokG8oFQTwrZtHUWRUvO1gUvalJwxxleVTHRwrDimKMl7hZY0L2q3lX
2InqEaq4kBh+yA8fIYO9xB3KZlmp4tQcakZh+lk4E609IbPeAz0V/vNGYsWhKBgs/YohXaLdgrQ/
tbKRglubsThU6tUHVeEGfUyUujp2BiNSbpfcUTLUO4Kny/WcgNshflOAD/6wzmM6Yiaeh5lIxslw
W7A+9Rr6/cO0aWqd1aEWE2UiWaG+VMNvofVNs3bxXRqm4PRQgydcak7b94RY036W5WBmz8naPI+F
52ud/8efBvDbczlsT8AJOweUNjCVFMd2mNVaNggucF5ijw44tWYEY0tu3IWy+2ddimW52JRY/5t1
0rO05yN0RzeYS1ujsR3Tq1q7URrBGrJhZRyWfLO2FmiIAOYoW/wMUGRdIz5FVSoPef3uriyAFyEi
BBTpMrwgE0EsjMrCCuRGqwJ5QW8twYvmwT0xURBEn9ieboPTUwei9Mc7ptF/5hRs8UHhht59qZi3
uVbZXR9URZ5kqs4yrsTH4DrkaZ4XjHw5mOWAuRlkJBCuNU42E4yg9gm64nog/XpUTiCfzGnjFnpw
D25A+jZCXOaNUxnIubSsPFfkRJzZzM/New7Vgfy9l03Fz9lupC0EYc+9r7+YY9dAGZQFpi+LWTIo
RXi/GsC2YnA2/MLP2/t5iiWEXHVqS15chzLKUaBpM5JW6eeIHBN/0RotYFCMvLvtPQtbSfv1LWfU
ry6jQTfRL0l809mratQfMliPYh5qMBI9v4k+Uq21oZIaADh21dVzoDIvYVrA7bUjUyDLvuXSvQ2i
Tklo7FBtbJ6V5KExFSzpSSrWacaPm+wGdnaKt4h7vVlOIoZS+cAWPZDr6Sli1JoIY4bbRua25f9u
OWA0hZdQbjHQWUn5Na2rPbSkaC62S6/i0qACms9c5mc6ItUJP+VEyiKYYitkwH8WHp6eQ185eFEz
KVjj1FF2n0BII1eNOCZrOVlifGfbwobnlbRauoMqq9ugnPohmody9kgqMV/UUSQwK22LrWrAL++g
rk1423MNccfYUndLBnQ8FemcV1ZF8ikENu5gYthO1ppb40Z+IK3ldkMtR/JjrATPNntjCBfkifXM
9NB66MQVlwXtRMbZAwHMiMeMCBWAfa0mxLZin6la7qqA7L79W2S3GF/UdUC8rIcJmDDuq40PDbwe
f9qZ6dMsL6hSgYaaMKAq03p01GEBxaeWdximlAbzVdM5/Wd15OuSrpHDc4hPpTm59LqukABltC/7
5x0BekS/cgbjuNLMvdnBn+vEPsqo32X/hn9fpl8YX1juW8fTl1MKJyG8nRChzPczDb1HyzmLxnyF
K53yQ2+cDFhXSJ9bBUkmgarCjuOQEEQjs4J/9TJ3VbmsFxEgUIaDE+sJKd/Q5hmMRHLuBYHdkzZh
iobhWrQBun/JaScdsZNtHs7zrZUfwA4r+ae//ggt4+6EYtd4rRJoCTSAjuRhJT9sJIQ4XyLw30RS
tihYtzns/D1pDvVKFGyrNHL7vXTKmuskBDoTna0rsOytnsdgItWfVAK0kpiO8n4GChOSTX12NSxT
AMbOoLn7fdizu4KZhaGw5WQJ76rFpvBAG7zjHmlDAAXUSXXKaHtVJpmoMQePvQQojnGiFRSApF1k
vkYJUJ0mkm4zDno0feU6yBeRub+aj6WMhg0Spceauczev+/IxgA6OkKLGPjoLzRT97wgmJYXKZtq
3bTENq/1qdt4odChRu8tgCn4t109G+wlh9wBknkyyB6y5zQVpRxmHoqH4jUEUX7uSP15WTNSYnXZ
4sHGiNix4+LvMRR82LudkNPlKttpQXWJy/rDN1Sq/3aggxqQLB9rEr1h8kmmLEBVmKigOlaxqAn1
7A9scizvjND628Y5Ht/C3cD59CebVkiM6b87KqVeOBrlUmaw11UyCsk/VvBeJ7nYmL842bZRBtSw
ahDYi+OuoII7EYEZQPI95YxtnGFq/KbBBMZHMIqb/oR1DfDwc05yPxu7SRQbh6GWjewcf16qUxDK
wKBAueHhPrVejJn8o5kzZqpO+VAVObkm7RrQwu5BEeOXNuohxGaMdq0ZF3n3Ywav8fnRyQgDPGIU
bw8veJJd3P5hfTPVIcK3DBngJQ06Be27s8BImpDQN1dzipO2gPOfbUsX/GIsZLCd90RZwBXEx64z
WWvT5hbZANe8/VGHGKiLX+ZOmckapvPxww5CrSpWLp0A+z+aCoTiWfgHsLdMszAwAqMiSgp2QpCW
yuUwwzh1uoxVDWOABVB4eA2byO6VA+yGkLKPhM3mDdY5IU3/bi2ICKY9AQsQRCkv556yioCPCxjH
P9AVfyq2N0nsMwNa91VxT6VLpkyUW8p5dnhxMqvd/JCByumwGy7zn7JsKjm+lQAqHv9lnV04FStF
VAs8A7t9sUFX760li1/Ia5fJcNqWvYP1QKM1pCFnX/YtJjOOHrZ736ou9epKcv5DckXfD09aMBI0
pe74eeHUNtSTx4bLpqorb7daWRPws3o1EZWRo9cgbDteBdmRWeC71fM6iu56hslhCu2/pAyUFawP
Q5zZGs5M5fpFqADg4uaJCgEWfJ/P8ZqTtKzLWQAaU/J5azJ215ndFzEtDEyCze60nWk/ejEQkTRf
sWrU+pTjP5eknBOo2ze7T2/w6Hp+psE92fpD4D0IJS81YhMDcr8q17NhXF83vyDtuf+i9JNI+nEn
wOFe26KFHA4tGso7prpMUmBXWkpOzA4lS4UI2kY2faXj8+7Rk1IGMaHxlDY2bmzKNvbAsqULkpNQ
NE/Q8HQIkcWql+amfA2K8Zr8A4znDJcY9aTjbBr+J+eEaDVdNaLINdqqylU7Oz/N2xXQ8lVSuCRK
jAIeYJfqASwUh5NqpjdLx9UC0A1aetaimsJ9ZWN84idtvg5bBAZD4dXNaPWyJ9I/U7utLGbyjmE+
z4QXF8+vbpZYXVhL1nxV60WyNlvEZieKgIkKAOtqcNEcrgFMeeEyhNKCpgLsEHhdN6REjmg572gq
x196UcrJyxgNIawtM7YLt/wtmoviAmAkq12BSpD2ta2xDtFbYJCZ4KfhYKDk8zZCsAJrZaYYsxKM
ZddGAzg18VHdGnDPvLC1xIpRyWljL8EIkLthq0zYe38SWVY9YTiSK3Vq6OXNh7vxPv6o4NnferEp
p0ytSWyAGuhtMQnnbH2vCdwtSXz7hp66BkvnM5oT/naFdMbFcubB73FeM1REG+ErrtQ+VR1MbDD+
81x+6640v16qorh6YI7Sm+AbzXFk1r6o2iYSdkCnPP7K8ltiK4AVjbplFdYeL7H0k8GXRZcFRvJ+
ZP3jlLtGC8NUsixGEzk4tLd5/HUm9yjARKWnGa2CSZdUr/JhY7Aw3f2D1yr/jqK0KNj4Po54WBXD
fS/SIox95W5dvu6v4vIhPpqBOB0UNPztIgU0s9bz4XgI528aWwbE/bmmI1OiKk06ZCp0aJeZWw/5
QbDduU9bbHBNUcAwJD7TddKGP4jdEzVGbv0wKS/gbEjGHUTR6otFx8IeX1fHae2m5Aeg15twddXE
s+2r79Ggq3rOzgPMnF1A7athbWV/PuugHHtnclljZe4qBU9pZNfpykeDwA1QkNreF/i9EcWIz0fw
ksNZ3EZPu28oEPMpi9iUjFGXUbqiPsV03smuno++aS2SJbS5Y0n5mgZ7+krg7Pzh5zBcYIgvdsyT
TxWLw+yF/SIhpWGO0fJ/o3ZqtxLvChAp9va/h/eUoNCku3EFxJPhj+1r9jKCSEHpJXz1Toev6sP9
yWCukdUB7FWjEwpd0Der0yFn1DrlCSIdR58uFL1vSKERLtyS6SD1lnH6jC4796BRN1TX9MDkEz1R
ORbfyPBxQwZUNG7h0Z6/5R3igXdKq+w+YxqavbLDMOH3ChcrW+VIlTbftzlaqnAsfczF6r/fG5mh
Z7MJjSOLW9ouyHYKDfdxxgqqRu+slYpkGNU+NudrIAwEOoMqbK4G6KzYvsOMCAWovTrZzJm3e6+3
l3KdgL6l7hAGdB51n+vRDleieIjM8SOb6gU3nUE/Ktve46DG53aHOj0kDCxVWJ3WwwDC6WxmRnxi
0S7PMZBtaO+W3sLiTxsiOr71aih8HXSZ92SrtBmeFcinZZSwOy0Lmuygj9ErFjs8Rs+Eh/vnxKGH
K3u4IlywoQNiTcF37ogg2iYyjWUwMzzz1d2Yybs28wz593oobEuyESnSb0b85pt/Y6M9jLCHNxbT
KsUlV4I1Tc9j3fdwPV1mD+K7Bfg1lImEAs4QHAe45LVD20ABhWx4HYIrjCIh9CoHOXPbkqQdfRk3
DL6tC9XprtAYQXZbI/QNHQCoTkMT5OiwuP9oRtpGg2afH0ess9XzRk6YK/NxwKpk7fvk3eQ9yr6o
eW5CvPcdB3Y70OjUARa9zBh9m7fv0te/fBvOZ/XCyO/9lHZgqqwv+mRuLuWjSATyo0PmwnDtnAnu
XTeoHLF3iO8mRjuSgUulk5EkD/vwtdz5RtFRWnrXuKo048OzSgesk0Y+5uCrXcqbzpuh/PhbkBtu
Bry3AHX9/5VLAsjHZtxBN+AibRhyOLi2xX5c9XPBgR903KsKIY5RNp2iib2uWGXVxOuoyswJODPC
eLPVBM9WQFZLXHQt4H7GUPuF+tN+sOXwdeMxmhupv1YQe+18t8BLeqcUf7HaTaj99cFv539nQSGu
74rckvLSFCzfznX6XIwBp3f3MT00DvEYG0Oyof4LCE4TVUP0O8QKXm4YQ3zJzhBbngGIAFyGPMTS
ES9ba3UOTWxveZi4h0SAdxm0IboUEf0jMjh5ORIp12i6gbDSM3pHKxFPmPebP7T9ymQAfzgzhwkl
Umzn9bz0u70Kb5wDvgVdguvPSxHNeVzGvOTaTvAfNkJpV/tsYxs63MXIA/ZhDW4U1q99X0Dofv7C
U+2vONANzPooJDgsSR+9RhAF+Trx51fElcAb1Y0l7kmoiidxXo/BFoPX32k3j0TVOuFdz8X6Ox0E
VCWP39GpvuANfy2a8jy5dXvpqSC/NmCACVRSf2eLcPxP1qNtnqXR2qvWFdExkUBqOqyy+lKIzKoI
cJ+8XwPVfjwpsigwwk3gjFS/IPbfgROq4VqXI8f7cPufxi3hmooy0KS05yD67cHS8AJEwRl3vuAA
0wLxAJDsPADYMcLRf81Kw9koG9jJ0C5zxJ2URiHL0yKIIyC7V/nAlxZZhdOTHI5AJ+S/4LllcfT5
EZeVfQdQtNoJ+6EbQb3aS0wtwy+tslztdaB/4MzqaTOdaFDctga/XLCE3gyQV24EZWw5muNOV9+n
KWkUTn5ACw+B7xYSn3IOYS8bqdFUcHBzxehnsupZxRPPH8OKs2oo9Xu5E95D0q2Zf6MjXgHcfBLx
mQuJa0IIuNpFdsu822coxj+tncwdWgVRzoiA3xuvGsfxk1W7hJO2TfuJFyPoZjm/tfYSIJbIrB5R
CR/nfsXjD1Zt2J74uKSQPmbycfaQka1XnLf2kjTA8wbdGXueW7Lc+AMsaaOn0HrkTLWm0+qY2gWp
SxVi5rFNaDckU6pcOU2Zqqgi+5POB4RvWWLJ7RoWj29pEoLULnvpyeC1G0MtboWx9lQt+Lq0pLfI
lOlMsZtJYhjfRQKIINehB4xvAxaZCDtFhoCQWoQEirkDSwEZwdNKuVrj4fMCCe1SWI0JP2Rc0Jm9
gkFNpHjHqQlx8k9M3s6qhoZLuBkJDqSjmeAIXEzrJ28MNJvA47Z0/gdQwnhSmCfbUk/xMEAsannt
wxqdCBB8GP4H2VZDjRcnCUbO1IPCYHAnAkF0Gyh4XaGYvug7yas08H9vYuTrMzwDJ22KbmdJBB3y
D3RmpL9od/bfOybnBdKPFcpEgy0tskAy3hnM1hz2DbZr35PE9aj2ctRhzmrUYNOl3JF8wQLhLEKF
UqNQ5CxDbxi+7BIq9s5uNp6IUK/A48LIv7ClbfmL1cqPcTx+I5Crptck/OF9N1/G4pu810x8JkNV
x/7b0JyHMZxjJ28QZSBNnLM48BDCHPPumkoPx001BZeQ/D8w7a952FqlNuNJd9RcAB/K8AtCqcme
/XjwCXF1UlpoJvK5fvkD69SRR6/Biz1qKp2DL7RlfRxOCRt3qe+tN2LI0fBqJ9xpwdD2rfhrPRDc
910DMNb6QMuP3pbGWbymrFNPjUqhGfqvoYbqVJkS8KBtI/29OkcnWo6yTcNbvcFZnMDCJDX7r1pd
mSsvgnUGcwFz4cnFYjWMIwlCjdiqhycAjPoJ1/8q9F737ySeWzE/D330e254kLj2U+q2bBKpObeM
+T26fNRB+lpbl3vjEOfvEXA1vjZ9S7//p7jg5N0Yi2JNljaEi2AGrTcwdkyEibuQOct2cKqyuEUB
P0v9bHuJu03lXTSNAk9PQTRrmlbzK4YoJs88r6P/366CTbAnJw/VCEJXsJ0OPoq4tdfvwqRBXvy0
obSJESfWq87RkPzM9fOMH22HsQ3imd+INaEBH+9UG9KTA0ozSmHgVJ/E6myMbe7JQLYC66Mfukug
zQBPOqxbVse5Rc7j2XgLKjb5+g892fgqvFg5QSF3xV9oppTBdl+JGHG6flTGG691XzIS11zjveFi
xarFpUUtV2UqQrRRSIQRJega+IKZg91BNNBZbRcro7HMFQ8iN7s8fEk1sbsui76sWEi/kwwZFLTa
Ql4wqFl9vzPf3g/aLo4LM+/akmTJSpyUQ4si8fRRWX32ZkUv5jx7AgOjuonynBIOR8OCl8FTAE3V
arCYwJVEoF2PB155L59dNcKoVDKbUwZOWMADXlihroPpvjo59ty84HB9k6uGvXipjPNY3lz5s/2+
vf+3Fkq4V4owjBUxgWmgnGlQE8OhgtKHyIYL3onMBYEz4X8B6nldz+zEW5XB9zzqQr+CpwuxMeM3
TFZtl7NuTY/HBBIBC/uBpLPCFVi7LUarV0Ae5l5ZO+5x7fU3cJpreioM4Q3FmXTnRvBfvrqVK/y2
wrtCxfYmxteuX/nxjdOQPiMpfgCZw1d28FIuKPCjtzwW2F8pkuGP/cQvQ0XvhRZA+p4Eb6/3Ov67
wDeI92LpL1n0UK58UHR8gixBH1i2L8xv99MdcBmdmQljUW6p046QHhAsp0e/rA8Rk9DbghW9WEZb
AJ5Wbie4oxNbMJHKTEfDx2ICUo2vXQH67EgNJ4z9PdrcELRILViqHBPDOoDDVL+F5s5MBJeYmYBa
Rv+7d3kgTowS/Xqf/Dg9jAu/0l30T1H2p5qmN0VBD+QUo6zSDtvjBBh6U5scjPpBL/bgpTaGP6WQ
t3DtOZdKmecNmy4FcD+JQB4AYz4u0RbSNfiA1KT9GSrTgH5I73fpPcx7IbotpfVLfg0wlwREK0HL
UKmuHLppbjIgo3JPXTwpHwe6n6t0GvoJDJ/+zlVn/UR/HkEpS9u5lk6k4Z7H0w6bjjqE66VNRbrR
p+KTzJaDmZDmmdaZOeuurTsaWwmXswjjEe8aWS2sy5coYStGoXVF3a6p7MPGa1dVU+nTX9LwD8Xn
JxK+HcsAUWt+O9yRG69YVyqcROpafct6lQjd5j7+K6vfE8+gtrvu9w3oopwuFRuYOG0EydwkH9Ko
ullCypPPLkSPzOKsEkTe22R8pvfQ3cIj85qykfY/ebYpthlL140+mULhTV8DaAdW7njbRtAETDZu
DFBalYQ+sJG14Px7+pgUTgnLxRpxtHYgfDTmgImoIGRdh8Ms8yf0xHKJgzumYdYeyrCaD8LwiDV2
cBQkXh9i/olIAEZ6Mu4Qxqht1DLi+2udAqzmAHW7R1xerJPZhu7tSCBq2OG1ArGjqGYmbqUgs2WF
3fXfUleWeD7os3Zjmyz8Olofd1fIdAdfvOeCiFiGQPUlg3ieMDVCFiO6piXepb5jn6okef9OUmFc
TPCeGI0zBP7Kyz2v3UZwaoKHhY4CcZgUJK24rAtraTMVgpgxm8kfZrLmdZV5PjrYlfjS4OMhGqY4
yc2Dfx3zWy5ohpDzy27WHqQlFoWvpyRffx9ykahd6DZHu4vz59f6o/7WLPo9SWy+rtBXionhPJ6n
exjeRHLzh3kSuIi5VuH8W2Jlt8o0J1CsWt0NlSjfGdshXCDr1U7FlY+b+T+6MCEsC/9M7rpTHM+Q
y+8RGEgU6Tz73oLhFv/bG2XuF0rF6pyfSJi6O9kk8DC0Ebss0ERcZv4AWFDWQ879ep3cuktEzCNC
pk5z+fRSNU/c7aYbkFlXa+8mPEBw5fkIbQ/qKK5g1I5jNhNuaDYwzpV9aV4HazF5Rt8Rpe5JjbMO
cJTKi47wYBNhpvofcD6Vig8KRirr3WQ5ZGjasKlw0CCrEE9JYaifmonZY25sQwApw9PlzH0PWSfL
KdC7ysJ2jm+2gdECaxdZQkv4nmUd0gFDew82WrjdjN+uCD1EUPOvP6tTANPll3mIPOntSjnYTWd0
Ju4xizr44KixPWEDnt5tl6Ej8LzNjaG0IQ3but2ptIrBOzP9FuEtCnjVIZv914eNA0M3AuBbP9gF
OJA+L7pZGJ31CjNlv8cnBnXwEd2mxJxa3WAYZKzOQ705IW4/zhE8IuhvDmrUl+rNP4NQluhUYad7
WeQTc/goHlPhD45xJvwcPQl5O1fx7I4PYqNsG3Cw/3XSQVEtDeuf3QpZ9ExV3dWdnj+2tES8WXpT
Tzi+Q0oec3iIYGIeHvZs3s93atgK42vuMY2ANazBEQwMXJzVGY+zLe67l6haYTtWE1B+RRu/BFRF
xw6ST+nzVsM/79E/pxcTjT+PvRWiA21suJ2Df1O7rh+eqtFiLDrlpic5DqtHAtN1D3VxW0DlkiQD
mXYIoapnumje6w/JKXxFHkxm25Gja0vEzL7utIqSeMx1Z2/CWIlSjSouUGCTdQW1D692Lm8Gf25m
vDqTo8kFBwRJ+RCDMvPaoXsGnTUEWq/RdhHOhWqbwVp8s97+PdEEwvdIjQHqFltYDfjmshwHWZmq
dzOWTrsQ7Obor/hW8riM9048YZ3Yw+/fsoMjV3kwAsMSiyfni41LRknTX3qA4aDWSk98uoTvAiET
v9r+ONOnTVEqNTbOwc5NVtc22m0itOV3cgvdIfNlFzIAm/H2Ce/xmRcCLwHa6EnU2F/m4zGB5qd1
MSY+MouNTcScL4rh2lhCDPvxwnKBJSzxHLTm4U2buea+O72pa66UIjTj7kfrI+L+CoVx1O4ADrcW
g2BhBuRXWPCFoeYvmBHTNZvuxM+qnUJydgSc49gSC00GH3tsqovyJQqmeHs9pTbOTKHLr6QeQhik
IX9Bbt4JrWDeZFSg+ooI+z77Ojzk338jvE/fWIuVGSpV9ZVGSC9ApaZglZ4T4VNtBCOmhI8iXNGm
OFrg/WgrUrBPrT70kxehMdmnjdh+3bo/IelFOdoPHbcxtaw9cUlF8qf7gyhcXMNOtCeZxkhN3CI0
mzE5H6OOh59HtdQ5LLiGQIp2v+mz4Pti0bQ4QFQVz9KL0IvTER74S0rRtHiZFrcBjPtxS6MDPkCz
PiNBMCvubRq/XsyaYNt+yT/fagXtaqPoAW2pRTsxbLO5xw6Dn+fKkDTemnItCRXELE/lL1qBx7Em
wgUSL0Q0BAsYHegYDLvNUT3ZMESByW3yxwc7/ALB4Efqdcmv/D0Xt/sQJWOSy4tjx9swOBm1q8nI
GFD/zyDbYBzcnVbQeIwQ/C4mf1+Joa04BgHUPzIAiIc7n/T4IfF2qXsmgLkALnWTN8VCpacSY0sZ
qONrXJNOvZq7oWI17G5mKBnZdghPqKLPGTx+VpUjAktGFvlBv4Hdg1HoaFBSU9lKXej9D1uUxg71
Q/Rn8kTAY3GPVmx4R1V8F1utgeW6yzNSAxL9ZZjk4D/mjF9a9IgQvzs1ViMw//ZqcZCdcH2ax89y
oASfYfu+KAmbsg+og+Trw1ReP4VL7zWzGwDVaPeVAlG65XhP07+xA02KujG51DmP7GqvY7m+fkwP
MJuCczNt1SF/CLV4FWpcDEGrUFOxcPoo4Ci8dI2Cm4jHOc6kFRmutOMpcPPMYBpV2JvdgWovPtx5
MhtH2NPRrphwfuiMywXWSYDQzpHVGPDi9VjbkGX9mALowBPtW45nYgNjNtcdNY8Xsr+8QHANImMP
qiRYndK0Wwns//NL6qiEOiv/3dK5kFddC84L1SQjcmS16gqphwbe6l9VxVj/hll4/InbuEivnt48
DJQtHuteDH0TKG1ETBHbtud8kaEDW6zGzurnIcw8VHjqGRzD6+z3GJPaGc9QqWsq8lcqyc0Nu7yL
B6JyEXf3gosL42Xun/E5QggwitvxhqP0jfTFEIGBgHTtgIzUJzqGd5CoPyaxP6zx0dsAHaGxOX/X
aAyE7OIPI1PryXwQGmIo/Rjw++S6PqEulZ+zEVuz2GzljsJga73p2ox7eDayV3lyk++WRSZ8PUwX
JpY9Yp3XAbWdfrOnEvZAsMBpaopvkCjpXz4APoVneHDxgcjwet8pQ7V90m3dk4TDDmbgGz4Vt/rt
3O8vbuKnYNU6cTcefyBrnLSxq2uWgQK9N4WivfYOtU6pBuaf740BruS5vyyD7jRDbiA9WZGX+xmQ
WkQt5OWYvrZzHmIZ3vPW+lnroLZQKvpnnm9EEB4HK2F2Y+55QRszCIaPhV5PRoZdAwPGt8LISroB
EfyN05vffggsRghg2fN7ZeNp/2OFsA8mb2rnY74wDmEVjmhiKZkW/pSsF6emEZdqbQfwcRXqG0DI
NHLACsNOx5oEEW7s1gxnYVK7tZ2MXpNiGJM/eiERhxDlmqOCvYL2Qip4/b2jF9A2W2snyyRY5Yy4
/XvfNCgbL2LYsjmhPN3lkyHEXdvbv0YU4iWz7YIj+bqR4Q8WB1JlZ7vBaJYY4EGPpDlBW8S2xQvJ
7sr7Kv7zNbUqivM7idIAerfUBCWXvHHUOjCi41dtVdfTXoLW+tI9k9pQyPzn8V+01VaZYLq1ukiO
GuAB8SdSArINyvt5/B+8lQwETyb3rSYXbyrD3D6z/rGplTsM7Ppiu8WD/R6eKpwGbV+CISSF/c2M
YAoFQGmMRHiVqoAHJEoN/p8yWs3SL2YgSCZb9XkDYKv/9fAq3d692BN0LeJ15innqlog2x3NZNTi
+mWEo+3xaDoWLSs200okFI295lZGxFfgW+SW2rOYZbc4y8pxwmLkkdCkV4NcHVtSHhIfxGYGRUpe
CZRF0lUPWyC9VJ/93cJFnJ74EDjWFN9mlEdNYukH54KMoV7ltuUil3Z6Up7i/RB5mFx5xFyBN/UU
09p7taGRqsLkm40iK9aW/ekvcGxeGw03CjvAfw5DySSOUtS7GSXUE1A2tSwIorTK/TXfQY6s7DsO
BAihY0Kgkd8zLE76VVQQyAbpR+BhxTMLeKg4WuqjgvOeBJI1oZike63Zv/lY0m9Qp02SSqqPl8vR
x7X5fXHi9lVaEOBqpRFz7Y13tN+GRPcrshBgNDPY3pi2FgkRGIGtRUCPot32yQItWs3d8DU203gJ
Iq65i47zs35rpN5jW1mJhv4eBvgmpCqCXD2nPdXqjnZ4b4mbMf1mIt/kvmsHUDIeD5s+T8uhHQQO
YIBJVcmLXEMoPMoDafCMjuVElEAFT6MmfMqNu1TbpgEnNRuuKX+0VUpWmW7pdrjfNWMwfUYQCecq
ytsFcP+GSh/EkW1qvhamWCacJJcuYEwR3w3ujLY29I2amvyDEhPj2asuXNHWXucEYTIQrocb9G0p
nvhmXlRohtpKPynErATedcZQ1X9iaqYRG//IYXHWQ0kgwXYrooM7rczGJ+luPzasosr1nkfa7v3u
lKifcmUn1B4gyD6EB4fgYgew6ZPXK5eXv66VMhrZvgSEIJv/C0OEBRkhFqNJgzgN5ZU0FMorpRsg
2X0Br00qNA6dKC/lv30A+HhIk/EnB6ShkwNykjdoC+lSJvEJnrZchTzrJxiM6lEOsz7qoQHE/JNm
yGuM2rCIvq+GT6uJ6NhDyeN7PkylwfSSuI1cUraQed6LyNr5BrRzLYl5PTWaSMLa9qe3F5Jb4Fmq
FVmnUurFEUda9RG4YZfYtvHnEdnOgcllY4qHIlSPhHe8gtKmKj69cC3Pz5f+r5FnMwlmWzcBUOD0
PNrnxC9wP7c9oTLC4XSQdptNqN+P4RxzL8LzP/2+5rxc4bMtVnBVFxHl/vZfUDeDom5apDP/3SBl
yuCV1pg3BdA+MHLsgMUocgkHuvNyLfbK4a0S/mijmKQZUiHDgUqeoCcOP462EgRguIjFCRmJyYSE
EAkhKQtHy97sTD5btidTZGZNWQpITFouE4qyT4uXe7zl5NVldPjikWblTQLedTaJc1dpQUeTgf/0
VtcyOMrOasLVwZgRE4Dg0xpXg4d7+nQVn3o8HBPaf07jEcP3MPpu5co3VwnY6zEOA5JUPDznIW8H
uHOWcdhD1Qmr63omrC67ieDNKd4zCBbENLxP/uYLikdYNHkPFkmFpBy3ATVpKReBBDWJPZpAWfJ8
3Samz8hwlTBk21NB816Rf8THs6nj+3QNaBlhubhN4SZdRPMx7pSX7Gdpw7N40n6WiGW7h4rtZQxc
sWsc6f+8NpzrVRcsi2/E8Plv08KGYxelbfMM3RMH58Yvee3aWmQeJTTjjYuKSuSqta8KafX25q1+
qPk8aYrrUszKDkDY6AFD514RBHJ1TfuxOpYQxmTON9lHfICJzLaj9zDtSHGkxin6feZpiej65Q3E
nJFNcV53FkW0ZxvEz/K00u6gMb4hNnbO9yLpP86RVbtkkKRGlQ2tMBT3x45GeLL/po8H1JZRDtC4
qN/bTpN92fJ2q79e7+jBi5eXTYpsFNgtO47t6vL+YJOaltDVrPj92cZbhLTmaLkPq9jykV6SMq5H
ARy56hmDZ/gTtQjLjCUQcSYakH34ay/HTHuBZsoIS5MCCQWiDJ0VpMBt2BURudtMIyO/XZe0SsgJ
eMrwvGBdx5pOjxfBD+ve5hjSEHEwQzrjov/2T+9pJj1psWKhhlCNvghf8omRFZB7QEtMpB+Z+2JC
Am74hFA9u6t6TB4XtfrigyR6XTWD03hol6mKvaKXbbYcDfntFqt9p5ok1RvWy6Xn6b3e+h+9AFl+
CynbGcVVUDgqBzZFr7f9IcejEH9GzNRU32y0xaBjOy899rZV8iupfhdwG/LGIk/Uf+aAjcXOKq16
lw9CE3O1KLsKOdQQZib3x95c1caMsOjWvndKSzyapECFTVQPiBrFYHubijlRUOuykAe3aha8IG1m
shWimbvqHwk5gJEE9Vc1iwObOH6K2wKsPANbpj3oidhRoXInEtueL4563C0D9zCfjumNWKiZ9/WO
9krE9tw3JpCbx2zN53lqhuJvakTQGdxtUdFb33ogSkpiqjz5vtxc2YQWoiW5ifpkRcklMxcV4Tyc
blycl0GvypBhK0CLGR0VKa5pxnhuL2dTTmevod7sJZr0l4StgFSQ8FEz0UqvUOdcn+iLtzWod3OF
yU92V604dUPV2H8B9CQn+l8w/AsTeh1lcCFnZYg70cn86ewkIs/vygktVsODVeRmn558CMfhYCwj
e3oVgW5QNd3W5RRjWobHAqpPLvl/ZwDNYSt4lGcf56ZDaoND9MnWxCJiYnZNJCP36i0GSzu6YQwW
udOFIEniHo2MIurz5spghShxzyLtMAsqqh9Lkap3E8WNbVAv9L/+Dr7NsxTJRoggsk7STNY2Mg1f
Gr8s0Coe4aSqcQn7jxsUe8+KisAOd0XfHb7QERvsF9ZlLH9rrrgHbjFIrNdVZCJYm19XKhPt64VS
uaZVC1MaM2oHYGZQ7w6Cn/bRLGjO7/rxH4Wck9oMNZBN/a4/N6giLWuPK9X5EFTN8ksIkn2Xusfu
wh0ZDBG2opDNn+qVsa8ucqNC4g03/b4NFWmRXgSYLU2yv3hVhjhfzpRWxB+9HX3DdGElF5MtK36q
Fu3ovOmQFAjtKHqHG/8eenuOZeFKZWnrIXYHrSEkKlToz3DX1qgaks2LA0vDAlsHJnbZi2lW1vzK
UW42n+rPf1HvYkjgxG6JyACRYLXKkgGc7uIrjR+mf0Ysn4zPGo0fpCuCaXh0W0CQORF3STyiQI/L
lD2x97Lhwqg4KAMLnBBUbJcRPuKNWG8oSWRuMLY70FOfFjwy60QCD2Sj31yES57RY3z8cj+KQ3tA
etnO1rdcQHmEdHKrIcybkfu05UdIVYwKei1B0R3te/7tZPMMZhVPVYpcLBJtJ6HsRCAojxJiQqUO
uVQfZiTACluLHq2F9va3MPHne+HvtFHGg1uzkz63WNH0It/GUAlaKap+e74sNW3dP4gvpfZ7sY54
ZYhya4G+IOTIgDVRvfS85mV9qOXvPQSHj6vxUBc9tiKI92nWPU6JdV6yyUi6W4v3r8zMUmayEB83
g/uTUDWvGRV8XQk0jUdwDpvvuppnzHK8ZelZuo+FExdjQPmdaI+xaMAfbzwC1MUqSW2qsiQt4oCu
z4HStzplY/lfaIFTn3NfktVKpn75vQUzRe7lFagPAA3roFfTOkXgQ6ZB2296NQaNA2knUl/bqnHu
GPvHxsvPvXMpZPmcCvNwAYPMrP3dleDT5903cLDFIwI14A4QLpQOyWfywDYnameC4fdc572ojgDe
B2744yxUwjU8U7jeoH9e9fZ77wxV3V7HY6TRyx5UaozywYCIql6YSTWhTx3zCFOCrij34Rl5VU3U
r5M7QMhd1rqW38TJFyellHijRFm20Ay3rbvLc4ZDRQ41YNvmevhdqyAsLqjyM29yxbSGhdcPBHDH
Vtu/GKHcWMdfn0nUArbaBLHmZj5MutuBdQDEPU7qfBd2tw56Y7NB6BTjRtaEYd6rAvdJVvnFaPcD
x0ShZrTyhx9qJtRlxGfkNmMmz5RFTMkZcGHSsy++Xv9898GGlRT0aYjLjwgbbZQoCRm4jqTcIoHR
wG0KKkioAjYj9RBVE+nOAdaUkjaxBNPC0pdFbPhYew1RwCZnUgut/8NxjkfE/pNauQuFDShErKyK
fK7pkEaIDubP1QMQKR9H8A36acaiR+9k/fp+bMXQ+Dm2HrO0ltfBJ5HdfaCEi7n8yPv5BktNCoG/
i2KeB0cWR5S3vUrVSxVXKqP0pJYsIiDmyAu2W4an35Ub18FTS09LjzJuXd2KizfjJYfDMzvxIT1E
n10yXokVf3tT2kuth2yqAgomzQgGOZ3xJNKaJumbMpZH5aBzK/dfuVVeGIs9k7Wboe50l3DB3OwV
aRgScjTDi2rrWf5fO7VdYrP2KZ+eN3uX9WbCNKlAhyPE8h27j48Uyi0XHj1d+QSfRoHlfRv7k2Om
Ng0Bq+HIFhbptvZxrit/RLfH9n8G+NKsuPFbpF28D2JK5ScquG/4BSFJg/NKqU5fKs3ymo8IaMgX
ftU/cqCyZ95L4T0Oe9ONgZ+Zacl4VJYn8kOqQCFmxvEP8+t0a/UQtWNzYAr4YFWNUvoUs8MGA/Vi
SQny+WA4BzpYZMxOE5cJ7mZf4LaqsTUzCfmiidvebzVvSVrzku+ln9JU5QyQWDJLgyrwSRUnR8Hy
1tR/M+qe/CSKZAB3mjugneGmBivN6yIFyoKbpCkAAK2JSlxqG+j6vMRL3adEEbKFp2YneNCLoCf9
F/SXoPzjkB3bvUM2OhaNFW4YLfnsZVPsWfpgnTBNtAXuJJtS4fMeqv5DLQQTBuWhLyBoMpqQ3TN5
RCk1dtbeubS0HViUt5aCdsdSjoXRPc1A8osFngItIhy3Lh7z7Lzkpx5Pj/kyGYhaSXVFWlxUsOET
DqWEbui0foJYtbfzt/qw3cpqAX79M/6Rb6Te1+Dd7QEb25QeN+OVCob1Vyp2Azc3tbadao2zglMf
DVvknlX1PhrzwMU7v91DK9Lp7XtkStNIisBNafFkYUaqcxVX5SjRDGIti+cCl/bk5qUDSnMFmtFz
Cf6hXB3vDoEg19Fbs+6IGWN+c2YO+D9rWMiCGjOcUCrWivcmgebNXBFCOuaHSta3G0DsvGcmBeqs
y6mbzd4xryBjwoUoCFqsWuD06HORe6WDgZhFG0ysqBqGyxrNA5KR6Sj1z6ixoOxCqmheuiskX8R+
MOl+cS+8OvZJ8cQr3vuey1BZ/sCJfydc+Z1GdRGt44T0LsOqDVYZQTM+hRQc4vE3vkDm3fwGjSq9
/5XuGr6Yg6Zku0+iDJ43ftcPliUT/nXWhzQrV7ME8Xbc4HZQAMGkUJZlLVsxeamCu5MWxhjDdZw9
b3BnLObrAMwzU/YGrEn7dUstLdZqFfYsDGWzPoKZYQQvvHhjfIkHr72sZ5KU/oEmMda5SvyjNn1n
dZ8jBGvzark7Ay5bg+AZ3NavwPGhg9W537pXowi+LmUe2oMTLh7J4esSvTrx702PWpD1tIVt9cn5
bJlCm9biQyjHE6eqndgdEnqA1/cdGf4vmqHE93/G+hD90C2BOJsUeNeJCT4Bj3XR0ZLeyoxSQrnG
hsLNBGfTsPpO22ExvJ5JW9vLdOoTcSkwNZpKfChY2A9nDYb3E88NJ+JXYiWQL7jPl5a50WNAMIqT
+hV0waNp3xxnELxF+GnZ496Vni5CInoHCZUY6XQe603SaCdYITB6CoHVzCXeZ2tS0HFS3BPgnRUv
U2nItoeTUkuojglhFZCgSSeewLrllO2s+BHPC60erqeyLSHPZaomJOaxqOjvtkEDmZ+mVHkVa0Qk
vnfn/4ene2+7RBc8QGW5q7dyPooDTWUpUBDfB7jPaNV8giVFWv1QaUIvBCTPDJE5utfJWaciW29b
+Wli6NQd1TQHvdAvuLaXYpoUnTRjPxwKAH6b3id4WxAGcdz2l8Jq5j9XvYhhL+2AcfjKwdtyl1qn
aAueB+42qXi39edd5fT0Y2fE12lYgMeNCZcRoCb/iab1pk/NDqbhlT0W9nQjP18lWtITNQo0XrUR
kwfVVUxUqjfUrsy1qaPNjTlXFaaLo4sJyOel0ufgmyx0OYbJW6MB9MeMkwBlfC+ag4sWZpVa3sAz
wazi8ynpQA76EcPHfIyjDFHxKLEm8t6bJQWBe3DuiQqJTscwMKVZsnpEBXsraB8gNYo2PzjwikQU
qyv6tQo8uncdCk999WaYiYFNp5MTq6xQhZ8NdTYRtFaKrd5S8FMqzghbJBLt8ET0gdfAAir3OoVB
fQsRT1SVYm4DXsGME5mnFmUiMmelk9l39xj39x5PtMjbo0WVNMQ3NSwaWB4d4nsoD0UzrDwsqPSi
XXOfzdJ0HDbUdgYCoCexH27yt7IOBYpm9Gi4S6dZnb3VjRNbFT2YoC9fNVtIpiC1RzjFBpbDD1i+
2IYes5k6Z65N16bi/7DbMO8Qg8mslOsQxEQas23RPoNCBuO/E2CYfRFjuX+lxsDbE7kLCbtnvw5S
xxNDpyy3SPMyB3BLWtf/G52wTYARL/rYXFNmUgzBY/cHyAwFy/bLTNDHEj7LADi5qdhyK+66AwWL
qQ7vw/EYn1hz2B6T8MLiRHFEeGSAWJC5Yx0a3F/RZ+mGEDsBk2VCfS9wk41uT415muomNdiZzJld
c4itIrSdNMDNG5WWnBJeFLF8oksoPZcDtlCxseItYwxahP1vijwwBUtNRcSiLmHuuvRyhVzhnZXn
t5edzcrFsJqdzYoZkJJtWaFrC41AjvzvouWYXqDAN6qjQ9FPih1mmYoY2XkFMJWp2Q48LHPo/Q+1
qsLfjd39nHDM/A9xKBF5JCoByEShwLa4f2RzPhl80yWfayjbLD6G3DpldyRHsuN25XcqZF1xnhaV
k7LUEKjbzB3qaaZDQ3WvD6TbxOfPuhaFtGML9vzSirRl18vRiGQFMMXsnusgY6k1ak/CNYLzCq9n
aPVPE17rNazIeRJ2cDu1P8L7ss2tFqHtTHXYowRsi8AY4v1wyczdK7JMfGFHMYfhQcJPV5NOScmU
3l109zVEA9HfbiDKXpcd0wvgasjNXdN0i02mL5uWIV6VpsDT0V3wBKTT9s3jD2Kj2j6DkyL1RyeF
vURLSSe+RZTprqGersICsZAeekFYDebZw+ShxipYO94bIpU/sC68j8U953YroW/JYUQDjvBTbeLS
wIkQfWIge/4/FktUVE3njWwvk7qSlA0cPeRj9N19qSThkiyeuhsnWtdOdDjIU948cgdGUBKwBVTB
tMtDkL1KML8UD3odsoib1aEBWP/mssY8cgZMNxzDJpE0YTj4qW1QfP9+4JKSD2RJMlne23uQS/cA
vz8p0jjh1pr6YGpZl8BvK4WoUErKgYGwU676eWwH5pmwGrOFDoHasd0zcDM+YQ4iY0kCkxurBgo1
lX6Odku1CUMAkpuHe/gqm9LaPxPb6u3lOmMSfz2+MQH3ddIamOnAjYa5F8kgJaPeDMv3pqAt+Nvr
GjaZOsqjkWauCiWd9x7b6tDoHhOIMUHhPstvz3/BdkXp22lwloFWt6SsBCeHqwrQPZ8ep7dESl43
JSeQXPodgCpWhcxX3EnLl+wu1Jhklny0baL9+PQtAYYWigqn9RRJljqLxaFcW4oeu6L20K9dHtYJ
AMF2d5YlaYGJehLfsOt3zkQL2fJEl3Vldo9B6fYhcSLVK0O6UKzky8J2VOeY72FpVZL3xdOt1yLL
tpmL+7JyyUcrqM3uSuKMBudeYCPMcKEvOq22IJj4td4VTvYWnaF/+HbQgx5nUR6vV0qhGbAuZ+YW
ih1MY112stf7VmOPzR6FcLKm11rHjFra07yNGn5VOuL8rCjyIZqGuG2THSZLAg21r0bvtta+sX/I
r7EA32M7AtyaymgI50sMt5mzCuKaqpx449SPhjYI2dq5NUOKkB19kuijrmV4czKHq6gxRyCMDS5b
AUoflAjQHKUVKYm5px2g29HbR5TYdXTLf9FW7eU5gWA9aOHFVG0FjsCkf44e9MS7eJiDkKLCxf9b
XFp3qNLBIYu038oQodxvuuWzCQCVMFZDR+YfRgVqczrtwKBl/C8XmKsVwRH8z24KPovSKuJInnam
M/MOuKzBi85Y7LGJcsyM6p8z8IurU6X9dOP30+zcG0t0g1RPtW3KPAc3pF0673X7Lhd++kB0Hxi7
coWRjAtD/bbc1z1emWP+3NZeDelYowCK4qwGxtHE2xyS7IfC8ejRdm/LbPi12R0IuVYodyfc5W8y
MFmbeRGe0U/AuBM9NKTRJf+ar7dzCTZDSLoV7wCcKe9+6Y9IA219b1XGqRAgL6juXaRp+9yXao6R
Dgu4eVDpQ5wkfDnaCm4m5WD/R857J4Mr3qcg2HHC0jL+T6YLlMZhu0ZxfbRNj9I5W6Eoo7TGC0HJ
vXEx5/UU0SI+wgCqZCOrwicj2MjBlyFKOOX12OkGhrH9P9F+jSB5Nj8fQSCVx9S9Yk/FAXGve86q
32BL52R4QR1ycXr5XEmeu7dqYCaMlObZjGkEkh8P2sM22ibSpZM2ex+fIBGjrSKP7oY+WhsBhg6X
KYs6332090Z3Xl1nLnoV4dRg7LSbVU0MYm73UTB0bmUcZ7KufnZN/k0vd7WNUprAOjEkmiUS841S
dwHjnkLwVTetsv2xGvMsqlfsxI6c9N634GPt9rZLYSgFN4AS1qYXrYRp0kNdo8j06Al5a4kjbjwj
npCYScnkAo48Vj8WwbJQKzV66G2EEidgtyZouLricx4/eJJDDw/EPcBI9+dBYPGMe8UCtkm2Rlwh
zdKj6HjciOcmrzRrIJ5iS4KO3i6fV+PPj8vFbZLBfRBpBbbSh331L3xJD7kl32/jqvJCV6FMWlLz
/11ulj2pGKH7n8uHLNsrNupYfDC4s2Nlc11dCiZdkH2xsTDhFuWV9cvI7MXHlQcU0k2imZd67c6P
aMFA8E80aTXWSRw3N1d9hV1se8YtqD7RjJoFiuI6jPRg+G9lXQamBePxpBwSTlTGuCYWyfWKMOJy
E4OHtSit5LiaV6nvFCXac5ZDs3SqfNW034IrvATzG8Cw1KXp6a7Y9lDAVRueHDv25Fqd5eB9o4Sb
lbi5evEvCuV7aAJ7/zDga4XUxJcT5WZ9OqTjBtt+o02PpNLuRXtO9mYOX12LTEhEv2H1ZCRZuE58
BOdOVuOIOkJqUcwal+Hq06c286GZyzGqWdT6TFdRHXqoTC+fn8WUVg6c2AVLxiovH0HemWqySmyB
ShOEVdQfx3SQDHbGH/5ZLV4eIE4K6Ja0/hpk6naO8cHgIPI6jYbpUOv9vWYXTXITjcG9dnqLRVlq
+VBgd9b5CRF4YOdeDJJySVaw1nHZmlgX
`protect end_protected
