`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
HJMgbjKZihIF5CQQ1gbVDN0wBA+aYxLl4VFMYwuOkTneSXwepar16bNlWEeh9JrvehYveVlFq4z8
ItQU85EsI2ahptCqiw7L5x6XDmaQ3k+70j5LNYV0iuW0ejBJqjEf7XYw3h2icJq1/DucFMakB5/y
aiRnlmVzV6vBasjjcs3g2xRUCBtHX4U7slNWUWyj1cVBuYc8PeO4HfQHqmZi6z/Wlp8p5G1uI0wj
yqs7OCj2K380/mxPuNs1szzXSTToaWotjFJFbLCEwedaz/Q8qKRTySRpEz0D+vbqUmKYPx4K5Zg1
Etho4ePvLWbrb0/4YXOAVOT9YTrOdvbDYjNTAA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="FaGFjwjCQVQ7qmx+x0C9AhjiDMums7hBz8sNNfx2VK8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4928)
`protect data_block
eL7QtuiGjuRhIUpD7UgzJFiS7l+sfFPyRuRs4ISRZ8q6YsLGTeMoVF9lEsBcZ6Jo4GgWrDcKnsHh
Ios9BZ3i2TWiJM2ACMj8kHEo4nHdDGHDe2qwKY1FHBq8T7Jsp7opcai1T2WRFfXkzsh24QSxuCci
ebSJuBbDsdTieuwekdyPRbgP42xWC6S/nEoY25eLuznxiA18ghV2XjRIljeb+4ipJ1ODp16x6VFs
4VSGQWNP8mmRVsgsX6CCI/X09/bB9BsGMRntoVMTTR2lxxLPkAkVzsRgq0iFsaILGNmooZRQRyIk
eGQFikktdAkF0GvbhdbvDHETZ3yiHE/N9zX3GWHHPAUNHaRnPw7ONjRFt2z9PoAqeR27vvYUo2yo
tbsrcY4EjkPPn9xuuPFHyKIdTsNwUfBI5Gc5FE3FxDP/5/KsFiaWmMDdDLAuc0ygi8SRAa88I8bw
onWsW199W6LFtmlV1aIxSr8ujpxH9HdLC1A1eXZzOCJXhrowdHnbCuud1ew7WC1W/GEFO8AyxFiK
7Mlsp8GIMSSPdsEjFPlGeUOLIUYgPC/ipZnYD4D2DQF6YBByqDlYH5SJhuZzl+R7/WxKLzc3RpC7
NhIryRT86OAsWmitCc+b5hUDVGlT9ZFHbal/XCcnn+cVhLmtgbusC4y6tTTnfhoQas7vMQjnsVwk
ieSprC1fGD032GV7E2xodfShVpR0lj7E5j0oTu7gLxH8Cf0xKU1ao7RbpHytWSr+oX4ArHiWpsbK
+Ubvp53P6Sck99iLdOxXKDtR2adNOL+AK0nxoQ96+5GwrNfPDxdoy1Wrd+R6ndyXmLarXgkbaO0x
1Y40uhraPUPSNjZAuRLVqcfxcvw+9EcnW+hU1IrYKWdsIsGI8U9q0B1OJ3Zo0VLWGXKnFBEGp9E2
p8fR+A8VUt0Hgn44NvULxYj9hOet36yarmA4HHAkjW5Wi2BZKvLtWTg/hutfubsRpSPZ1xe5dka9
eaRiGpCS3+vcQeBkKa0OezhdprMWAcNYuYF0SMlteeMGlM71mvaAfkSC65xkoxZXNx7D//WUQiHp
pFTNme7UpfZAJo6qvRIXDDAoiZppEwqcOnychn3uXTxYmrWJkMzUOVgFtgBQDIG8UP3uwnLsKUA3
uTqZhz6aMS/QqK9VY7stXSkXu3ai18sDQ+fvjrhh8pYEpJ0kA2G7LcJ+gbCzYwbOCNzm1rP08Uxq
XLmPypkWWLwWebqxnourRqpzd51e5/D0t9VkeNe4DclQqlAa9RXTVFieTi0SNAgjIdYNd5rA9Z18
EJlNbJr5WTEdFLi+/YdeSuNXbuyPKXBKmPzU2MMUosxh+FFMPWPAZopvRAhrPpI5cAFvWzVK47mp
Uq3K4ZnOe9ZQgrC6gdLJ1P0fjiYHDkhBC2idPsJcb3uZoy4g4ZriZd5ORfmabB0twxMWtvY/2j2B
pyynRwfoQ1IOeZy5v0ReZCwZZxQ91vr9NhEs3IHak3K/XyXalQ8WViJzmLDFL0HfoM/QBHIVxFSg
9gc7Ghp7u14M//Jm9zzASvqpr46LC7Q9gXnL1wAlM5Q/zsOrBVEYynEBz56nRTQ8rTHq4yRVg2Z0
AIokdY9dzCcUR3exs+GeUg/BSytHrlo+e7b+m/tb5Yybunxygv/lX5+q3gAxWHVuDItSdGa2+pv+
LuVruprqRPSsOKO9swo9AlE0B7ROqNueiiPtD6VEaYqJQeffXalndFSsC4iHUieuWdn/lnaPirM9
lsJo43T4qWTC6YPvljQnhpD2fL9KaP/LT5G0JZixiLySJmnA+qbBUFZz3De/x1mgCNbnIJSsb/1s
YC1WGwqMCDQPMY/6dvJ76LXpIAz7xyxeYFzztcSbyd7/OJCU3BA6sY8gU3zC7Uu4go+RhPWViaRs
WKn7PhORBLUyn/PApf4s5vICbCMgMzYDjAEbCH6SNNp6t0uD9US+2nzxvR2j3SCjlZaJrlQKzmjv
x71OGs1yc/kBippySkTuQ+L18BYT6LDD+lKpdxPOs1Unizu/Tib7HsmSPegr/VlUnFDhzOGsA1CG
cpLQqgsb/eLCTmlIfdjCle0IEHn7rXaFmtR+efPBwLiF5MqzG8G5Ct5a7etYqoLT0DR+opeXY4ot
Gy5Hw5d4jPjWaRYhExNxYIoy7XPErS8FM/2vCxlEGUET8pTursCfQkZSDvwE2J2m98613z3jKmQS
fLKh3q8s8oJnBHMuxrS9tbzf84XwTtKvoiapXLt0DlmAnkEjMWzDvQIVVV5uUcprPUqXp/sRbshY
1JN7sDWUOvVXDu+Wv4g9BjRNvveuo7KLOiWiZtWMVGSrAoI7wIuQVwtmBfsbBuOIGznYPHBg1Ey8
otC/uA5C0/DE6kVIYfpKnMhPFsmxISQUmihct9QDshNhul+lghXZlhIQbeBS3kZbLMCoUdg04bMR
GguKPsil3SKmQSgRmAEwtt2nOzPcMGj4iW6ASEgSOtUin5QMUURSkLKPdNoWE943uJyxsYbGfjAx
sxS71iT0PkXxQ18wI6khRUhUKv342k6zYdGhddssu/+RqRPyMBUdENxanZNAL68AXza3KG4R0EQD
B+GtHj7wYnmV1DinIAkOC+t9W5BgUu1gEdzJc+iNqAug1EuseqVWaY4ln8cLuS/CPFZjelo9N405
hjyAB+anfPGewNVszNOGLifIsmTCrhgB79vVuJ0U+bwd2MR078PBX6DVvq0sR7lM1jf1jImKxfRI
IumAAJY/45Vcz0bDiXGJ+2OSHvXults3eHJIiayHsHb0dqzOVb2Jn8Zk7iAnwkKmvpGVqCab0cn8
yoFm9n4D8ndMT0eS33HurIticv+ydIA+lm/rFb+N/o/xmRRmClDbWYsui0qCO30euYStO3ndUzGr
C/YVTB9+F1jHFLpb0KXckIZJyWGmdXpn2anHd5RP5nT0EHEK70fZpG3PNnYWn0A8e1Amo6B4DiZP
ibsiHVjIuFeKBjbfbGH17sYMUEw6bXZP+v3qdR8jTzcaMdfOBBJjY487RSh0lpaRgujqWAQi9hrU
dgf4jOw1sijF56yd1JicjbqnUlnh1CcE4vebKHQU6atz4oqgCedrdcZQXSAI/L6CFHViI8up1E6e
g+ttnUMwCLiFn84MDJJUyth1zN3acP2y0NaF7Jlj18KbpleBUZMurLxXKfMYt8hNDH4wCDeDOB3z
pWJ4JIfYBFgjRLHjz5V9DbVVfnR8TrnqMWkGVeFGW5hbeI87IYc0TpzsYEfk0igJFt8MVNP041G2
nIcUMPwO84QTbvjMdbCGZWqx5iJ7I0E7O+a9GepLpjCHI9Bv6PeE/lJB6NEB4P8At9PB/CHDTr+g
kSKlHuK+grSl2DEz7CrFGYKXL3KodEF14/bIfoL0OnFNdzJqVtwllqHvSRQwI8T72jYyOmssEIl4
P+uNzIr0JCaF1KzWehnQ7XCCHiUgdAfAGAqGcz6zsvGEhYIyLG12xSLON2nPyfjsoBV06LAKqUMh
RDImuFSRS8Hhw1/04Q+Rubu+wqLXgbz+cYCqF/yddJ3XQeL+fy3VKMWyM60qWR1QQFNve/0dE3uJ
U0nNulmGBBq32c1UMFqNzvGVkSDKMEkdGVCcKVHDijobymwBwwIYtcrAbfXiPrgNf0Jqr0T6DuFx
472I2VOITV0fZ+WYeSn8v+EhIBAzOcr1DIbkmL35U3ii2Pm3CvoG+BSbqoa2+MalZurIczRJBL7l
jg/KUseJl5Dyh+quvhPmYFXjOtjxViAu8G+6KAxlH/54m6Bj3zvGy9cyO1MN7Kciv6+ncPkfAhnz
LzCC49cHTGh5j5dnGcXlFV5h8o77LOdFS5RVojpCM10YJJeYMWn5lLWGk7JDsw64YLmYidcDYPT8
CCwIhh8BIjkagmjvHflIxqb93kq1MAdDIQSNIkhjaC7tI5R5ka0O7TAzngIfYjJrbF7mwT4AlTQN
pYbugenuti8AE+9Q/O1Qt3gbae8ml1bOLaM5QbZs8fHq4f7a8LpaQeLdcq/xXSqZCliwMU+21B+k
n/rJjlNHNNdZmV0inJDf0bzlui9z356O8ZWRrz6BAaP5Ny3sQNkAPK57EldjKL8f089rfQOb1+md
3Df+7BtHCjUeVu5EA1SuUkfMuK1fmKq1fd+VVQoQYeqa1vj6fe/BvO/EzrVMsohroHf1uCDVwDgg
eFVGAoHqWJ5BQlI37KJb51+leFJMD0UHTUNg5pkhNzzHXQJwbL+j5jDfyfSCO4YrJtpqYJh7djON
z5NlcsfNfbChyNoZiu0DdGaarvtDHK+QTuHhgWKtX7KU2/bkOT/VipZCCU9qyBhvRKkcrssZPe1A
LLFPuvN9TN1CeeHGrOsxNVuA671xqkVbJmQcR9vZ15YvPCL1vrOclKMgU3ppb31YhcgN3oLpjwxC
H5J6QfwlLOdtNC6jOAN2cVY5W+CHI70l9Bih1FqrBnMjTaxb+I0v5tvGhbgEW7bV8JcyVgm+1/qP
Zj43Ucft95lpdFDJWM0MDZPCKOGMP05GWnYH5WVHIGzM0ye/5Xdxcp5oGGjbkr80RgP4eMUprhLI
Nx2wEjCbFPIbRINhq0XvcgEAZ4Vsyfuscl4soXVu1cbtZ/zWnad5QhM5/rBRH8xuN5ii2I/x56YX
RTLRKVS6qYO0jECAanOecSjTMXtpNXgJJDUmUR1/Z7IOXtsHcvZTZLmGkNWA2gs39/d1r3oEdrlg
lZVtGWPYIJGO47gh8LcX7NDvkbv/WAIp0F0R9bQvPwNSLT8KaN1dpG/Dl3oMQ8ySKfplssW+Y88J
yHe4llGhnWqs11oOvz5XC71qbt4cAqxJGRVFGzjUGKpxx1hTa2Jwzh+9AhljJLcP9/k1zDNVnKnk
vIlYO22XfrHJ14xsbVHptt0p5zvwvvuj3W0EPZN5BiVkuesEuop5TngREsWnzEa14baSrV4xdp/l
Ep4TWvSKMWJpTH1gUEJUYAbYRgw0HXG4VWKnV/MSSncIwX53CnUx0F/egLySqVrCMLG7JccwRrzq
5PONcJbZ0rAuifxkW9T0EvZrlYMDFEaANU1KgObBjp0riaym2gATFQXIeyMpBwKMVVgi2Wr7HmQM
h9cZNnUFaazLWZop8NclOT8FowMSkjmMo4iPQZWOqao8Ly0G9M5XGh1rgH8SDKZpV0tyUc+xbIh+
xgNsHXs9hqLjB6bDUuEdPpg7AJ9F9YUIh/AI4p2gGN3pU7D530T6hdMa4KAvmPOd+WXp1E3sOdfu
nPiFPa1CHEfnWQVLVLKI84j59Pvvu+PY5iNKJOxdm7dDhZn2BvgCMe9KP/UhLeOoqJkFB1UkV+m3
31j75zBJSvSFzbfxMFHmsfwtL5WHxguSA2KC6jUCdBl9qho3rI4ach8j/vSt9m8KBQhIpsSo8g2q
lCseSzKfjSlm2TESy8hRYq4+wTrvnokkfHVcZXJZ3Mn16HPzFLs7D1gJrGY6lhV4QjsRhGLtUQ9T
QWkP+ygwyvFbJ0wc0DHjcbwunqegFw+oo1j3fMceaKB6qHYWLx6HCBQASdVlYIJZ6bwIPexCVpCa
i6aIkXBksDTJnxeOTHrXzNBZ5E26OamXYPQbVCdnvqvEZ5LOYUC+2dxknALXzt/MnURhgPcI2iZ4
CEZEiTMbCxA8qAhzV976FW42XfYQa8vCprR3AIBTzRDCtW251Y+aRijt0XuwhmvbGSXte+SCqyzm
fDl+6/mVUwjCXvxShd+3R58Vs5s7/zsPTTwmvW3xy1oUuIo2JsBY+WYZgKrBeoq/4Rl4gTDvxyLy
/AdYAGAn+l5vbYOhBlMeo4btXJT2l4iKpbYzmP6diub8fVcDL8qJirLwvj2BFq16qHuvXbVZUKu7
xJKlbYqv4S34oE35j4tKnS9ODpdPz+aeMbWCOjq4VPkrwNM3Fts9ZdcHy+tbhiSLK3u+6s61BcST
8lK5d+MqHQ/qWTx1TzriWRJ1pRixvC/TrJvWdbj4lsYQLCQ59QPHvRTQhOFZYQkpSKMDanijuN6j
5rKc+uHKZsnPqNy5GCgfm0rZV0Qmwx/XB1L1T5dRoA1Lh7K4NxEYJ2wcZaEQis52HYxfy2ijyjgC
s6E3yyPJ7CwFz6/lksYUabVFKKRoHk7L4uagHQoIJYwwH4yg3zdkulj5xu3L68jdQCAJ9u3qNLV+
Dtgg8rjrw73vSsmyMftqCnf0OmUzP8OGaNCybjLU02kuJYbXAII+Mf1MMumvvkeRAoL0dkLEqlGB
BFx5mC+0/+RGlolwRufcDiBPlDqXiA0unru/AwjuDaG/6Tfhl6qEuma/Ug/Bx93SrEdNGdt0USb9
zvF24SMSFDy2NEbDBACC67wrOOQaQk1OLWZoDsP5Qthm7sinGbCS7eaS2+0UrENKdnM5P4VArqPh
mmax+K5t9SjdiqMk32QlM/msoWq3RxQDQrNkUTCtfLtK60tj6ocrt1twOT66q5SbJ/eiOqJlaVrr
5QjA9iDZQvDaqA4SZEHBQRSzydG+58oQ2TmjVlMjc+PlT+eP1N7oprhN7jJ0wgR4RnMDhnyoyxX6
+RdUm8PY+xMUiVBy6I1Pxmsuc8GISNp+zFY=
`protect end_protected
