`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
MXGoT0xQIf4q1fdStu7/r7mySjDSgXg+dFdkDelxXLyj/Hp2KjVNH/Cd0JzICYufs/qEtf5GJgpL
DNosu9OGpyo4asm8TV+O5z2w+43/sBsVsrXXSgNH9a7IP9itOOq2Uo9RqCvXZyS/rFRVUC+vWLIx
G7LTCSVR/vXHTMnZKnm45+EVNBAS1zDSoFfJqa/hbkxhK6MF1jpaCyUpUK3ghu3UxRdu6Lwp/0nW
cnkb/lnc+dyc36u7fhSeGI3zbeNheKZRr620VHFuvpuvfP1Y1VLOs62GUXsBs1REO2j4GBleHJ9e
mbT+sNYpgCR+NKa+GYBWANDzc/aVyolJP/ta4A==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="tF6e/f+KTHcuOq9tgpwNyBazp5jr5C+QVT5J4H+ABms="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5472)
`protect data_block
oACLVU9VLPtXsToBX+ntHJblpC9mdlUoEWZAQFNCuDXrzk1mGZPu9/GBT64zay6eXvYNnWwLtWgX
eoxB7bR1K58Gck/jFOX6hmU0Z59IGUazLFBn3ZY0nf2w//k87MNqcfv//29aI5rGkCyDFXiMW9tm
ML2eE7p6Bry43YWZPatHYn1273H4uer8NuoPztLfdBR0KkkBkCCTmxAqGJlFPcLnUmY6Cc2hN+yu
tPZ0FQtyZBvdydmB47ADlQKdsepe6CWc6SKqQRokKVpR5LmgDoyeiIzL5w9KfgitHJX5a1gRKYrK
haGJz7NbGUCzt12gNTLWQjxhcpE9mab19xV48DeEkwusSp6GuoLg2P1BKJ4i7yx8RL2b49Q4Mxen
tKX9rs8KT1MyRRQeURhBpdea1IOGOkIt/f9rY85R8btRhoM3KECztl/CaUgLQpv1QlcHXzjAQqvw
uWkaC8dKf6GCI9wBz1JSGeC2yc6b+V2MguBybZAaZ8YDi+hNtMxXRle+cHnfxa8JWTS8rEj5j79P
EaPQm9EfQjYifsfD8ZPJlFTy7ef/subT1ksJtVlfvUb5Y/DIPQQ3kjb8ZUgFlAdvHmWT2pQiOevf
i5C5nyZ/dfHuf/A4qeZ0JEJ7Joyl8fIre+H8L1DWRL4MsAKXWRhkx6WHabpFBiJaiGmmybjnXVRm
/0ocVD8oZgjEs3buBas/81rT619DA8Xbn+jGPBJvLdbb2ofrZ3qhMJ/xIDizTUERDkNiFyQ45rd2
srUP41Ya40ctceTRgLhzMx1VAu1DMtbGILv1ceZn16QEqyaUv1ghscZPwPnSiLGhrRA6+8HVVtrH
YFwI5UsOskAnRp+U2xVUt9HbEe92nbk34hmsBQW6GKFNWA3jVnvbY8TZ27GCt+d/kbruXysL98gz
IAi+mLgr/YgTiLX3A6KgQzv6Zj235Yql1g+8TuMtsJyfiFEZgc+zuoJYmXHouxj1KitiZI3ZC2md
BOr+arAADt+Fk8cVxOhqixt4DOb6qWHKc++ZibE/gAZzbaHQp9rCoOpStxUczHO61GKjKC1CnH6u
ioXGHfU6YOr9pGoNWUbPVr2tCVXm0PYH+Zsar4KBI+EI84cLcmGR3MIAxri+UNorPzlCmdE9y8nV
mooByMoFXueb5cDbCU2s+QmhssWhM3YNNx7HGsvtzCd8LfuOFRknYlZjqOCUlyUNFNAP6EclCCYC
4HS04Gtt5bF8Hex9xBiPk7/s0qmy9d7Otf2fplBp6eHDpt6bWyLOxzUk2BIltwVeh9xmXO/CQedW
z5tbHexnCQzQFgh4GcJ7Mn/bBtvF9ajygopmNWDWOH+XyUHlywCoEEw0sZimSBTbqPmc5e2r8Cm3
WbCWE41F7hstZZlDntRHbC8xAmGCldNJUDUCVROWPdY3GqVEXBVMzdyHs3ySDKXIq8FXB/TjTcvT
AVSIYP58YzCwthhFr4P1/1b2R+5o6ZnnlCMFqaF0khiyBr24edyz1VnJtXSMEx/CUF/1eEeMbFhq
j8aRfviVFRNATGffLrR7RFC1Nr2v2GDrMHaJEnmadSdtkZujb9VkVcWmvFubobmhTtHpOu2gK6In
23DjTA6JGJJCrTjxOtqUF3Lopy3Ujt1PRX1bPqNkiKgINUJE7xIgo1hqka53rIovN3FqcnZonmfc
jcJaunSbY63G1cFatpad0eE5HWfgUwfQZHvYDkO6as6I9eoFJq9XtGZqD9BvuJQ8Vqd+5s/mzSkd
apEQPEtWV4/jBU80AH+LROTWI/fdDf+nmU4vFVAGeTfYwr7qoQ7yQ8/5IwKGykYGHF2pkFtlRRYi
ZCi3LZ+NUV7Yb5oDqGny3Cc8OyYAyu3xveJplSHdFXCigg1bW8lPttyFad2wUV5F8s+0XQ0DhBAr
29ftTPCWoIl3PqrybxKoJPc1lO/mOqQEoN8OAeRXRwPcuLP9h7HljueREO5+WWGeI7Anili8akqE
cgMzVR6mocT90E8urGh+YR6O0T2MmuRK0qfyKicAAsoBhIdy4b4l0bcniYyWI+z2DcbOvXxB95CA
6XGdjSmYK6+cOJCe5Uhc/yLjfhWscfvRHBhyNhbvI5eKn9tKB+gOd+iqYrg1QQ6JCXAW5mK8W9z4
EHQRIWByGlclN/5f0pOkm7ORJeQ9ZyF9O/H18PR38bRWgusYxRxIRmHxq/skab4VABLHV4JaxVig
NLG+jx0s9YAxHe7ZuVm3suJbiY9d9gQCieosmc35le+e8I6joFf4Tz/fkgla/zONIvzFWCBx6V1i
y3fDMxOIz2dnMqzw34ZD68cOAI3z9Csd/gyT66Ual6akbT+apERGjAv/R3YAPHvwKPT1JPDMHrP2
POr8USDpuXZ0JCDSDfJ3wrw+Wth+yTdYSUJ0jW4iosu50dCqL3nd+2tidZdrc6m/q6lCcoVvFdKj
HjjD6T6R+TbTO+a7pEzkxWpBk8WtaY8DKPZvzp2YM5m2v2PGZo4h1MSZDBvZb7k4iHLkNLzQ/ndx
J2GCV3022kNUYyQHC/aYS/yWZp5AmWq83aRughwrTc8sJv9UtBtCH055UIqeI7ZSpIKKOY+FKyx4
QJp+MgO13Ru6ZYYgWjY3DCXsZI09VTga/2A/O9HQM/fK5g9pRFxjhFYj0C/qxxXTmqNYewnf7DM1
TTNBgz1yoB4oV4jAgBSE9yoGvpubl8JhQfbS2qgI/J4RA1V37PhhkuOGqLDeX6uoVLKOpqOlpwc7
EFWsreWjvCRJbgr/EZaNt+6ZDeQ9HRuRohoKjVH48g/IznnbAIi1/DL3xwXqk3bGhlO7AcmnM6f1
x28fPCzJaMil9UdDk/mnzdaey626WukO4uApQ1TFLJM+fvIC6t3NK5T+PBG165VMDGlYUabGgzRg
VHvoyGiq1mi5GmmR3PM5BH1BAigZTbnGxeVeA2ShCw3gFE99Ko+5E0L1yMw0E/jyL8klbvxCuhrT
1v72arA9cnB2dg6IBHhsA5+9Ng+oqxhHIInB7GqlX958irQvv/f3NrxiTvfv4Zc0OklN8teIUzbg
Di8qeayDNLcVl/dHYo8gD7S8eRlCxi4QZsCiBgLexwrbGXbeDK9LlzMpi22CPA8D/T7skwpEJEEc
hiSAbtu2WvoDsOa/GjAchDdVw/iLtkV6lBH+n0IN9xDCKIQ5C8qGyD3fMq952WmXJ/BEloEKThaH
ukwjHd2A/uGhSxOA73ZsR2CUuPcQtD/E6ejvSgkm2bjpyMRtLlCnwiOBUTft4O/iDLmHpyQoF9aV
EI//b5pQyOKB/CgGjrBDgot+GxwZ1L7njROe5mqAQrSZCD/mglmm0c1ybq4TSj3mET/38JVBp4O7
ByYF1mWDxf4AL/fqytZiPb3GI5/uHLBMLLBkBECntGhtN8qHrUqC4vuM8JVRXbZlaphPzriH3bqf
W9uaYk4q3Xzw3QNJKQDDf/SMtk2WDPUPRpC7GeDjpfSi+1JB/pYub6uz+Nlta9fYeS2yvBewAsxK
8qcVmtr7CzZr4SM4LDLpVEX/VRYbwPVw0G7BBveKPHx7ActE04XOyQ6fKRFBjpnnCaHHE3aatM7m
dxTwuR4PcRwu+d61v2qgK4dXKZWpyO496bvPvXua7tz66iB7fseAQDRlTehjnJnhH+jam7FDhwsX
S69GpvMnis14g17ESLl99+HKlcOB3k6KSIiGmR6cB48z1ByHhtIkd3fqMlfJjbilClre5P6gGTpH
sNB7PXh/wXTfyQUw8MGSB9HTPRP+MiYLVMt9WNImK6XOYHLZR8W0x9VOSZKhXyZBDnpM7h2vBw62
6nOtUsf0o1s0oNkzolos056Gt2G2K3ZPo/SRm9C1PwxpAhfQzJI9yIXLJN852CNFgR9EQuO0l8S6
llV0e7Sh7hVQPYYYtPD09imZ812rpPpcR9GeZDG//v2Iqk9AckddL0KLTLS6wMWtfisROmeKnP3E
0fJjjA9rTbFrSUXwAWx+9EFo8lLuvoea59v4JCOGv26gu9MdPz6BMB6DRb94+VH3S6yiIyLRNgXu
YtwS8spj/BU96/+1tXLzJ3uwajRQUwC0fgpENjoMJ0r4Y2k/8FBzvkYoMtBM4I9qU5qQ6Tv6xRMY
eJsS69PNpQ55zqTAde9eH+o+BvgNc4enyybw0Nci11VJmwBHiV6z9xvTxgKgeaZPfE9rLQUNQQ3c
WR3UmyT3tARjeFNyELigytIkozxlAVzJOAd7X7EB6IEviMRdZTe0yW7uscPvk4UCfSUhr68fitqC
BvMIX962lka5aeajmHdppLIs4ULTzQxC9Zb0mibOJxhcE4o43VtjU71xqagDgkva+XfVZFEM2FFP
bw2b9QOVEQZARm+OetKTlc+jXJhsINCd5tZJ6XYBQoVyOuZU529PaP3rbhX52eK/5rm431KQDO5v
+YwFVnDs64uqErl1DXSRSs1+h6GuE6ralcTZppKIE0aaZ15ahKVAYqeRh6/E/4xquoMSM1KmDo2D
TmsdeWSR2utTUIBZBIdGIcB6JfeUMOz9KjeHxQobo2QRdjXEQ1JCUFtht/HhsyIrnyfoHGL3xjOf
ksiJ2F+BiBnmEBOki1bPhCrUBAl1d9rbkHaNboAdlB3Y4/ak8bhIx+EGJB58lZXgTgcEr6aDl86Z
J4rRyKhJKFalNo+yQAOFcSC+2aamRR0kpgW7GshrEKjHX75RwnCPElYDqqNT/n5NZX4QYToy0eLq
m9LI4eTCvMWpP98TsMnwobsgVO6JR1I+EyOQc1QpRCOctZyBv47PuSKxlQONzPoaZ0wplDSisuVT
/6XO5rFwi25GhnVIYE5fH2Lb3xIEKRCDBB9ObGPG/avq9Wdx9KX7gnd2EocVJfj9F2b9ymnJHno+
dLhcy+sEMvYTZglJrM34Xa/TT9ZqCvEEAGIfqq+j8QKkPOO9lOhvfMNNoRCCBrlaidWKVzdyVfLa
pW6LSrgJ4jKSdVUenHlFkGJZz1iPCMx1Dqlm7pfdfhsybinamFvAAJnoe4jrUdJqEKyKnF3s/5/c
cSjHyTOY2KAFrjhPTqGgkzoPUm1nOrx7SbGPsy5dLBB9bYV/78ce0nOv41VsOful6MlxtDJBdF0K
6jacptq+DlNxL1gtP5qo+kWvxUUDijeUZQc663w5glPlhcM3gcIBm+DHUK5rbF1Y70jHcFPJmh5J
sa+Ui80VEVrnO0J5AWEgchEKk4g/JYSSvYyV2aFZbVwFjwyYVBu9hzPe43v7feDrSa930VYwmsqP
ncRfjETEbiGMATtwavQgmR9EGoP6Lr5Uv+5UEH8gsu/1N+QBFogi7SIk/JgW9hTylAn1zffOBfl4
w9/oq95PQGl9H5Nhn+Cdy47rtBvZpFdx7At/SGyh8ffKH1cVVtXwI6irYm7KEpEDCKvcAGnqzLBc
U0/BAn698F1l8DGQzchtHrU2Er2Km1cCjoCvGnfw/HgNEpk7ZR3QsfjhZJxPptlhCMN5MP86EjXc
mJve2DmYRPjxT9NfvX5nkyHwJsOuTUkc7dkVvZroQn4Nfpr3Gg9C9vGstUMhcQwXJWPUpI9WJth8
mZzdr+2y8qKzSVs34G211FfnNiXhPZQcIYReTvNfCT4W4m+nuUv4cbobjCBiDB8x7uqRZZm4ARx/
R8VYFYkdYij+kzTTortwAWFrb4bIN3XWk0pw7PMP5a/kXS/UTnDzGlER4/NyGWphj8+DyZ1Twv2x
bDOlS/wOn++Xjzt74m0eGb5r8/CQ2sW/3N6m5CIQo/8NsPtHKnZ16LEWv/XMCOABx5THdCzZvhXV
m9JCQzRvYQmOA3HIjvCiyzu5hDDaY+4QHPPJz3De+jVfDgoahTTKxwqEbp13rL3cM/yVpQQB3J+E
OU2fYpZ+FgvIU5HuP7SLMW0YocArp82sldz2IPN5da8WjQeDVw5NvYmS9Sj0zdd5C3QlNAOj9DPR
+oOlPKNqqiE5m8LfNtfv2+i5Ju1yMV3W3z2LVKdGmQko8++Kd/AKOjVIWfDtYiC0XWaXGiXO3XXH
J1qF8pBBi5bZQDsGQ/IKKIVZ5lNXT/hu8OEhvhe7Ytb6D0KgUUXkN6nChpJVsF2s/lAwW5/IQ15K
SuyfGnnml94gpdRZR3+cc6ZNEaoKbZ3ZPcP1SXCeSHENPjxb549Z7+0FHvwIOvFe5e6D0UdKm9Xv
2x0fkF6QSDa8yMbP6MU7WT3QY3FCZ+0NP4znfvP8FABjIBvDFa2vIrfNEs42n5qI3rI+hNY4wefB
+Z2HZ0Z0AIgdbJBFKYelBD51euSfZ08ylcR3HRILQL5EXgbD+e7rKkz4C0L0WyIBuf5OAJvSnUNG
c+LNAG6jjvJMpETlFqaz3zH/1e+ICy8gLlYjpDwpbfkAM7JgvFQhSH5FWqcE1c3Gq/t1FbvcJJ4g
h2+IsJw2ah/KQP8QnyvFR07OieamuUs1ryHPgqttpefF3427ieyHwFo1IbSQvJl2D98qCyOT6XK0
Au4qyBfVwl6UKPjIahJxC/2aqjFu9Ss57x2KIh4rE6YNLKpN4v/yY8Mgate/W15iCSDT9Kq0sHmV
tKaxnIPmKoPOgeO90jeFRaIIYj6qInEZGhWYGey8r3nkaN+IzuwoDRq/CaDzxgwyE3d8Ivz7DE4g
X1YfYICbnOjpO40wufAN7OcFDe9C7oVQ2oNCxTmfTy/PtKqdo5Ci1lJm9Q0yPU3xECSfmmVvSUSw
+lfxT6/mEt3AwHdoHIOWbLySxjsAk9ri/Bb5PQyZmJ4jbtRJrHwVrwLEMMKCrV1PP12DzC3VlLLG
zPa31kL4+bTDdY6hkCCOuy3q0g9XnDnoHfRkB8Txu4Qn+OAFCLtnMtuU/lH6H3/FfYPwoNKBPJyJ
cFmlqcOYtUoWzEUesy3ZEiMMxIvFcIXCjDqbTTzoT4aF7iSMRKYGf1tNf5QN9tCfVClKms/liwzW
SzGfMnN1Wx8hHFkS085e93tQie3k6P9b3ZvuxDrhtZQJG1ahSU7XevhVnX/WA6Sj/XrgU35XpCAg
dLZic9Cxb8qtlnxFMAGVQYY/7fsI6VRiz7Ed3792bGV6cG3/0UqYBA8WI1rMJh3mPvtu04coW3SG
G3MEq/RY2+E2Iw4fdTxHLZGKwzs1GwQgGqVaHDvj/Y1ANLW3PQUiZmerDlXGjCUL2yYI8HrIiOPm
WSGtMD3H1okrgA5vS6mlCrLcGqA/VT7KBfn7I9B7xKP3cf1dOKkmrjkS6X0QN7xlb8BaJp7EJA38
D5dEsIb1v9yBDIZ6SKkMZlDcEkz2Fc4IQR04wvqXJmohN2jJ05824pj2vDcMIroutmZevDm7doRx
`protect end_protected
