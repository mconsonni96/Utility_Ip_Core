`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
YmSZg0BtB1a6T05pQ9edt5wcgZaZGjur8UL3OXkbfRs6xm3q7OnGJLbHR/NntGJ2PAQW/GKllX2t
vfzJ21CNKrdgrVPjyst+aeZiVTYk19sCy7Hr/0Ijh8qFk14H2d9BnXsc+tWWnPo5OJj4r4fqVJPP
58KxdmEHHAitnXqy4eiKmygpLMl97qukvY0DKY3YeZ/AXnVHhetig/ctut6S7bG2ymqEZXVwfo3m
1uBfFq0SU0y5cNNjCQnPvvTpwaRUEAYTjRep68N6iwUi0p3C9u5GY/tLbejlSHyrEcKHkUBKaKWg
ndcwppwM/4BdbTGNtEnHh6s6qyB6K+SV9gnaKA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="UkWHBYlcx8dXLjLMkSzzt3mBOvCNwYADA3uWXcjfNDo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25264)
`protect data_block
8winiPOlPX6G8Cy2QQ2SzBUbQxpfKSG41/lVlXYip1qezq2YaIilHq0xnUT/0PhQNs0kys9tsiRe
UJp3rGK1hPG9TABD3GmVViJFmnCSEE5JfofhjrAMVwOCPZpw2+4ZsvOM4UCmwOxqZYnVQCfYAaHR
C+mLUr4lWuwHLKY+mZtgHxo3obZ/hB30dQ9/xUHdiPPuj7DLrk1ST0R+IEZw1TUtkGUzn5wysk/v
6tBUmEJEIhgYj06aCsp/4B9uQtbriSBNU6JGwuWXAyjxwHRA91uKT9I7vLyrPHhFILUAs4LDgtVo
W/CUD+k/aVDAs4lJxvfFEY97uUx/uv3y0gvxBrdBy3UgYa/6EsT/gAqkzV3bxRTkKsuWYc/Gij5y
z5BpNQcjwmgwJl3tDbzY2A6RtI/i0X448r7cjFstpFk0t6L4gIUjHoGhbmtRBT5FnYJ8JRNgTEGq
l6KlqDBEh4WUzyk+rQuPZfWy3w8hI9z01/bEvPkw3tnVsi7b3G/aSNlRPICUzbgrRLtZAOnrBuSU
kXYVwe4phHa35x+QUD5RxrdYoHFaw9mECr8RiNa4Czhl51amacNHcIwGWgYHRxzsxq7m51/P7veh
OdffCOP2zbjyqqLQQHu5i71HJCcgn3VTd8r1TmqU7UrmtWXqfFoJUCEegaxpuEP431jlzy8oPZyr
xk6aVBA2+JWiUAsr0X54JfZ0SWaS7BTXkma6UGYe0obTKXV2iJW0z96nuf4Ql9bEdqs3wYWnFOiz
lMbLkJIYMr9ipZB3M22WK1N0eNsbcV0eQv/WJVxxrQbypfkwcIylKUplHEtHbgSDAdZFN6lHVdiE
JoZCutcNI8gpjcqt6TH9mmSQ1ZIXq1MjvsRH0qsYONz0N3EI0IKF1K/u/7jfce/G4Cx6dXrcgo4x
PYH/MUUqT99posfCZ31eMemt3qnNbpRQ4bc3nM4xmD2CghN3q4DCCGbtsYWh279vOY0N4UeM9j02
60+czayLcqIvNZwL4m0wYOraia4mcyAdijHONLmeUL/gDPrmwyQwF48n+2tjzBhVGgnfaZUyikMl
AtL8/QfL5yx8WnUJTs9R2BZROxn6BWVtKQ2VrcYMZ79DHJbLiKXHZaI3/5OeodwSxxIjHhw6O7eR
wFJhOLX/MCPRPAMOhnYhOS43EwrNzar736fAQsTdD9BjAISoQFNGaF5UlhZEjNVeFjHN10GSlwFn
+oSWajTvkk0ptq8yfVTq6p8yy58STEfY4Y0SIR7/mrWSbG1nWRgZ3HvUjmY1HZD83X9Mn1etwQSv
der6UfnTX2/Flw3YCSt6CmOGBit3HuP8NSC8h6ACVhJdfunEgrbS5R+N+apDMSFxVJuKYW0OvkBK
qDGngbJ0pnRJN9DLfgxV/kNJ03Ft8YTe6vQlN4X8jTdMyKxsr173Q5nzBQ4P3Ftf9XM+V39w/77T
xCMQzzNt6Ukt0dKQUG+JkMjDlBhDNxP+K4efLhuruACjfMX9oZHeL5ng5Dcv9UuoTCtiPLSIUnug
81kLXFgjUsLAP/A7OjRnVj/e2/qMBi/jkPZ6JYvB1hKCVymmRyLzT0jKp1RXMcv8XTmpTS6Guv2T
uMvutwak64hep1jIy3b7ahA3XWJbjxElIsNGgsDfD/BIn+oRIgRxRDC0jxS8dX4ddt35gIFqQDvt
inxcXwHrIDFq4K1JHfNyZhGpPy5/B1rTJUPiOwZFttyKdPRmozBtbicRSz9HWnwIdqa5nh70ijLM
a99zQ212CQNK1lHLB9T/5GRflw/TJ27PM6klMhxBTvkWDQf6Ca3c9njirdnZb7l870BVs4NXcM3T
iot4wfsynm6t7oe+U0JqR5Eo1XPpX3/3gmR8salJTWcCEF/3pBLbmTESZaF4GGhJ2TzRaOVF9j/l
w94tvAu3aRRguF5NsIkvXamZstMTaRp1pd5AMhO0NSCf2XUnmN/120b5saOQnXQ4NthWjKMxmO3+
ZyIKfnhJGdpSWQ2RDUVhPhV4Tb/09SOrCdGO4vwWmmLEEt3Ug7MQiOX+KFz8TNSxfHSYWvSZX8rz
bYmC8XGMrU+M6878GSVzlBiTUYrv51zcu+knhHY5WBAb7bwTj8vaplks5gKSTZht2vLYzwxk07pM
eQlfWZIxjChoMGJB6Mw+LCR9MLkP9kbNRhzKvvDVVSmgbe0v2jfMthavaAUuzBygdZhYtYIjt+wf
sCi+Tn9tQckch3jeZpYR4JAIX22BMGjmZSsKY21TC7ouSMzJgJqb4XDTqa+BTyHItyV8ZnYkujEC
scugiuy4XoQ2+7OiXoGz0V2F0EYtWWrbZMiSRpRI7JLwWmrPbmLA8MuNq4n906jldrcwyytceywO
PQxhzVExN6hLylagoTowad894T94FwU4tRgRjk4K1s6cJN2AxzHMjZKPBEfb2HwBBeH/4/MZ9sCK
0Y6GNh9RkxjHmRuBXC9xzGUuLyZx/ZytYsQaq4oV7+BmhtKgeR8Yvk4G2N1cK8y5YXOWivG/Rvia
AsQrXyum8KEb4o0IUv6u8iO+lyaz2HYIfTXTopxRKLUTwN+zHYQxl/4kihi6ZdsIEVgaRe1E3Paw
tQJilaePXzXiXadq8qrZJISLo/BMTKb4mhkCftd5GjRdWcmZYNK38dAqVCVxwzBJSChzXaTzDQ0Q
CNH15+Xk1tb9kPrbRp6Fs25+Me0NFcJ2axAsuw52GEG0e5wQ+iITmcYzFIi8yMWG3xCAyCNxLzib
kONtp+HaZlUSmDBYaL0pBifJ4NMbtUF2L6Gkp2UZpJczmzyIcmunZoZOhgFnISo/G/sngv+N10CP
Fdlz+We77RkWfIvhfyQKwWFIUaTz1CMuGd08Yo6VM5Dk8//NGIBD6Ww5QxPc2D/pUyEYEO/ipE6W
xz2hLLBg2cq+gjJ0YytJAUOZh1JUJSGmNt7jc+VyQSJ20h4EOIMtbO3hswUGaWB3hR2OLtgvvdkJ
1vZmDQ6+hcENzrlYR305j5om9+4YJFuBhFVCxnUcuiU0t5MggaH4owGBuFlq2wYuMshBgtAjZeoV
djYSTrCKw+Q21HD0kytmO7NCdecZIafDiAz18Vd9mH56H8l899c4aot20ZEdsg6r1NjhvfilumQi
VNZhIwb2udNCJRDPfCydHafvwfWhZ2o6GmVzkn6XNVRT2ICTBJ+tzRKIEOSGRfB09BoJtiC+rxbm
abOt6YscqicaoWvHGfC9JB82d3CCW4rSuOkMhBxIUA+f/wHfdyyTfmYklE7b5jgP9bYKH9Lby1jC
1Xhemf+DL0x6eFR/whHHiE2dZc4PJ8/KuqtIttdlmcHcUvlf1zBtp2LRKfYGz2TQf83W5rBTKBwh
FvxbYr2i/l4fBFucdnuzpE9Slh2CrvI0546WkHkNGfqHnc6QT7cAfAVpZYtTwDVCt748M7u3GSrc
KVhM3NeVXmcPYPZWyqcmMj3ARQlsJpCN0kWfHsCZO7KsVgXE8cw+iQ6huV2r/xYfryM/MRdmFrJ9
K3e2EBvlk03nkkA2OljLWXH6PLgazDFJ6R311A+IMJ01b/q2mRHZZNvDDVfYxTvGiE2TxmUQcBfD
ELEGjczbjj6VBn9jAuXo2tcwlLhNGtzS7Deoivb7rLIMMwd5GMIscrs/Ui45Tfvur1G2MuFO8OED
IJnkc0aVvLh4GshOj86oUnQpDUAXsG2OvwreHYTA6BmI4baUjGzcmyw8vfhAP2RKU/gcnhhlDq9n
OozwT1gF0BaCNUP2Jf81Cl+Xyx/x4MN6RAqEmXhAHGWbF056Rb+hqLDeaoVqOFZY3EG2twuw3ctW
MomoA15qEydd4+ltQXYEGIbE1T0Yu8zjUPbTHtQFmohTpzFSy5RAE0s8Ojrg1Kf7lNBiI8GF8oMc
opdT9RdHhPxeo9w559R/vpIxL8CBsCCCGFwdwutQX1yeLjesyA+QGl99SX/Nsd5mqrJD/fPC4I20
w0TX3gwK2K60WkF1ApItYt4u+j5VauR77rEZRCdX5p3f7zAMiN6dWNVfMVm6+nbXOoco/jtyzJry
x9ykfIhMEN0p3g1IrTt2biKBVf2ctb3MIJVwk5NOafqY75L9CZuGufeW3xkDrOMJD37EucdZR+te
wG9InfHOhbMLoxDsZX+Rm58rILDGXTf8elYL08xi2v6IslRe2gGtsKys1vQCS4xeOiY5P8/RTKVe
gqtzS+VBhfomIASPxEFEXFMIGkErOCtkj7BiMDlL76RIfzDIK/O7nISxOqZeZln/gNBbEJdLwyHd
yf8aPv//Y+yHGqbhfbmw/FEgjap8wAFRweFsvsnzFrCDBs+gdtLFAevQU/q4qs3JbGpmLVK7qDVP
F0Tja/1mYWtBq3uyRdnRvOmYC88GW/SesvbOLF6XmW5X4caBmw1O4R0XL3dkphC2E96vQTS0xawE
r2Qrx51/u0A53FXfVIH6sKWSKtUJc8qkQXlNYVEhRkKAtoJ8dwD/LlyJvS5Sh88wFKuQOAlaVxgE
jKrfrFWhfucCDaLN7LMyi6NGvCuUPoiS35fcjy1kBtm2kysttiZxpX721CxUSJeDikU9JcNpCV7J
H5Sub9jAHFiLXoP74gMonpEAAVjCP9tRH+Qf6bH5MJ0mUEW/ugnRGTeRQ4YxXerEqQqjynSA47PV
CTfTRCiECirF3XuO5wAZPPvYIntU19BtznlhtCoHrF+kSkwX9TMVjH9axJ0MQmJdfyDf/TG3cSLD
Zk1n8P5Ln8enXxxXHiDaBEG11/FoC9NBNEKxRW2B5nUKB2lR8fFVqRPhvWPQW9HWYrdayFqiRr1H
u34wNkpgBA9ICiSfFhZOt1188C5HsR3RxMpidd7E/IIltijIEgDPJqRaH9hbeksX02CeFsmwfve3
qu16jSzh7Y2/MP2LzLbQFnsb60jn/y0kMSfkqrsK7+hbf+1LKZS1fVTVw4SmJLBiq9NxTlDgDXuW
QND5MoADikPFaK/TcYPH9DsYXpN/SaNGOraT204HViMYYisfpLK5OUJn1qpReDp5e9P3QJL34fTK
ie8yu0RA4QeLzBezsF0mjvtPEpVuqDdPsJcK22IYS8uVLrcpWM5FxMgWbcrXsoKfR5LcHeWjR3s4
9FxInrQvIsZbbsf2YLmA2jpHAdg6Oqr+2acw/XAxd8QElMbeaSVRWBGqW6UdLWhotsZWLyP9DFFw
lLg3GLB411KpP2zVEdxY3bp0VdO71hQm82jTkatPUrmD2c0NtoE5Du1cg8Qyq4M1sFWuXcK4mrHE
EDRZJzxmSNK+2d2p5fu5psmiW9AgMrGHy48Dw0mhSEMny/a+IiPbXmYxD41HBbl8CMlSR4s3N2zO
j1ZlhYMg27BN21aEAK6KvFcFXmcvwwRV2239pYYB7zDx0DeZt8KckvFotIcpNSwF+dfHtyjdNVT8
Dpnm06+ahc38BlwJx0LPf3GU2GB9sHw3KbbGGwD54HnqgDkSBAGIk6eRmPaKtluVx49Mp+e8XBcc
wkm14wYU9BrcdMkVT2aAn1lz0Tll/6v9m69SxW1X+1Fia68RGhlTNK4kejicgKKiZtcvEMzm7UDZ
XH1gmr2nGHEnPyPcnFAzdPPadUtTNWuzO6sT8TWmhO4e/ZfFkZQrluxTxJInKlfTl+Xl582G36+a
ec2rr3YZV1z2kBD+p/F9Vy4YL0UKlmFjrBuZrx11T3gG9F1pN8GcJPx4c51tlAJTt+hq/iJMgMug
QinDvB+4MRv9Sxihvon6RC7mVDdXd7TpT2QOYG2esfNEZI+4N6pHI+a+nBX7WoGOHTS+T2D0JXHl
Rm9YiOUBEgw7jZo39rB+TlQ2q9cvtdHhI5eVBWBz8/RPMOK0fxj3QvyCCQvZ/hirkiFK7js7n3wT
/W6r+pdWpKPbTn2pvyHhT70C0bPn6xu8mT7erTPjBwRORx9Jcqw1SRe4rWJzt0+JqLKvLjRfDO8B
6Apq6albArl7SxDNPRI0pSKIAFlXjGhf/7ZKKWDLtLQ9pqmWsx9CA3hAsmsQV9LNaOVBbzl5Bd/S
wrm9uCmilLMtVPy/s1xGaI+Ecs6iMOkB7c9NFMNstI3NaJYUbcM05aUUYK/r05EYB62PamEkckNC
zH6reQsbsyI1g1q4MfCQbsOSvoglJPsvDEg8TJrzc9k59YTFNTFWbvPnLcEJq1gkjlAsG9r9HvBQ
siS3t6b33Qlye9w4J+MzsQp6WXONAXYcwla4oF1gqz3+RXdDlDs27QgrBPgmDt5+RJOe8YcqLMYH
Ok6JenPO99puTQfgIyjIPyfoUWhr8EIwOHkgb2t7jSnJOcixanjouFXyaGA3q/2qv7TDRmdnzmcc
8oLbcpz2Jy0FdoK3WQm09L1GyiqE/eAC95oSFJ60Ipnvcq815x7Flel5gSbiQpJ1T0q3wrR8qMeF
zOBO1apfObWijxh+CRsQh3a1D4CYtLZCkxs8y2DdfOxZXPgHKL7n3bPHXPcINa0YpC853+tcbKFA
9teXSrTbUbYf30F+HSPipOOCWx7p42Zv8K7j0H6dyrcpYlvLNWaT2jk1rNRgDGxT81pQvBgJStxi
PQs0Xrfb1eChWdDbla2aiySihOC19Y3AseUGwinJ1gvvPbsrhntBrfhho0rBNvyPjskkul/j7u8D
U8IIVP2Z2Ljul5q45/v+LKlB5JrgYwYOITPibiqJKMvrUyvKsZ2+gYNfd9a/GTql3nTgxI32JMpf
uaCDUWXY3xWlzQ3ABxWUHSkiix617DeHhxafwD9XPGscmJWy2SXhKv/R4A5nr2Zu/bXIInlZMCSu
Qy2mNPmuYQm0F7AvlPaDrFKUR58xdzTzIXrTYqj4nQb4Eabi0TrFdlZyZKdoSczjR670cyp20ajk
x+O/QP1mup25C0d9kpIVcgXKI2QlNoWn+xcGXn0CeRoB/QyWLE2f6RrfSyxEI/DJf6bwtX0W0XC9
SLHa4MBUNKl1QAALeWc46dObDPtXESRiV+5w+zjAn0/44cMr/df8v6O2g3itHDd3Xn7G9x2naQFy
ZG8qXx1BIl0hSPMGlikZlgH9KPMNuv0pzhYJj8gq8La6TTuseWa+DrhsDl+c23t2UBqkQ09fvVpD
2c9XY84B8g8PFKcp1jdlUchuBPR9IRfkm1OHnrFb4+0SAIXvuf9iuTbjH9igs5eyLhCbyiqGtbZo
qqSskyG7Sr68d5VipDQd9zvg43V8bwOEOCDTLXUN57Nr9KHLKTfY7f+m+7pan7Yn0awZalJuiQZD
/Uh46D2k8xg6WQRGxqHQoC4Pzd/NnVDrpdL7paU1Eor6L6YHkG1B24TDFWmgk6pAnbYMdWG/vYGQ
kGiZaIAE1lIpD2s3kep3i6MBtkxK6FdCebSqkTyhIDNbbcCxokyUyUXYo7aNoeugacbkkneqcjSC
k6FPd7tE8NJIpqCv8OKl0z2Vn0ZbaO5rvjxUvhx1Z9QtU2pUoKDw3Wsj8ggf+Ofn+IpBKqEYEGRb
WsRDVtBr+e/eWdxYh9AlipFnmCKL6pi/QG/qu7m+9V5bDJ9oActSBGhv3otsRsn+54/v1pMdRD/z
JOIimAff1RhSM7YIuyk9CtwCoKRCwB/VM2zwPf3ouCzXfkPpvryJSlPb7qgIGdxjZEHk2N/19ZUh
ZPuV8hWHcQL2Y4nXJosjbGgq/hLugR8SEP7mgaqyQvPOijHheGma55L4i3j0bvmb+2+VMN+oddu9
3gHbJH7t4lfLgh5mO+oy2tUC2q8tOSxk9mDM38iWeS4bN9/9+GHzc/obTQQ+e3cgFNY8/w3l++iX
yGYSiSqCRoWwFgNg9pszzirFwZU8WJ4elpihn7FhMcmlNkgjcUjldX1oOdehdNADGQirgxmDmGGS
7H80yv+owZSXAqs9aE/MPEGmCocVsDu7tuhwATixvPilNrBMuTe1fCa66uM94x4FuEtTDCeRGn/7
nrfiYDRv1fhfvedpgg7z99ClXDSVGy+xkoMrBSLFVRZjimAHiDRXf112V1xbL5wsXd3Y1YT2Ex17
NrUmRgeFXi02hJHHrTvc+eSAx6uAASSyxEvGx4Zh2eDCHEP72eTAYNwGOON7JYA1yl5tUfulqPf8
Qva3kDpJ0eFH9L5UFMRqtEUEhq7zD7hnMllOy7FTzaOAoGpMWDn1TR7XnkpyyWSbtsmElrzfq5Oi
Rhlj+1CHufJSR/2rb7jYjpehwRCgiD1meG2AghIFhNOwPlBzWKEToVDs0STuw/1YWVC8ZqDZ8XZB
VC8fSAH9bLeAAXFhPUNlLaMh9znvIS4jaOcObO4aNZN7sRw+evgc70bC4GNoiK2JbIAXqGD3wK4y
yW+mm/6HpDVmk7JaS2egIhb34PfbU3LPbsg3sAmafS5ib5Q8QhkGh/3sOeEx4tHli6AhEbfiMpqv
u/AhldvXugKs7Bhxn647be5siwLtfOuihGHV2mzpl8xPj38WNRLi6fqt6PfFwLhkHL6RaRSVc+0S
EShU5rk9vp+XpoUyeTW8u/Q5TPhFcblyld2BxdTNw4CqSIq1EsjhKiy3YL3uTl9OQFM39qgExg7O
ippPAb5Ktz8KfHtW+tb0DmBOX+rSe4hYGCoiXm46P3nZbSe7ugyDP9Q1mDu1/fbAXOiipfJR/yuk
Orc0EXNXi8QP57Mggf9iCRhJ94aLX7an3MlBreTWHkppgYGnd800FM4b+XdaMNC/HGRibciKzOez
PVUF2LNeIemdwYmx+brCnsrNk6BHPpfzFbX/QSxPE70ivTxH1coqaogDtVhr8vbdLqU5xfKzKLvk
5EFmJD/EA88dRKskkttCGGaHsecLxvZTsb4fDxQsd8gvie1V+k4uf34Hr+nxBS+tY18NJ6z1837y
dUPfWEQ8WYlFXZw2L+WHVow+WQhH7n1gRwywsE0YAjdP2H+YtOPt9+UBxFCgCpOlzsNuPHxyADpt
tr/DK3m9yI6fvu5iTsnumZ3KI2mWCT/XWIWXAaeRXxjLk561QX0cv/bSYehHZzRXUquaZPbLlAAW
/kphkfErqyZ7J6Wn8NUbQGHdP5J1h1PRbd9+BJuFqoH0zSEVqP4+ofAhtzl1AtZ4jiN13acCKJUt
QmmZkHPGsYFguvqINHrr4vJXNlDpiiCQBA80CjoauetyyfaCmLJbZZnRCQJMW+P168jYbVdMhtHr
1LmKMRMSxbBj5WmRtG28QkMmLpffv/rSxUd3J8OGZjXAq4XxWGftJpeu4a4H9SiPUmhVfG1YszzO
EgN4AF+/BBDxQ3gYimT8iwdihVliIVFlBjRlV7YR5Td4FIW5NLl8CkcDJ028Ujz/DunIKPGASvya
HV3r5hbhqymklcMYMVlO5tTS1Y9BvEP5d9XyEzfpgaIJi+N8sTVG1bNUu5vZEa5R9FTj0MoOebhl
bmBAowSPVTmFFBTk0jakZwgcEY7O9bo/eFbdhe0pSxY29Q0Gk9fRIaRXSvxGePdLuZXNJIQcs5ym
XTAEvDsjq5HtutrWRrSvrpAFnDMBo20UYptpyPoUz2vrgBktVYWdlNk1WD0cL0MH+wnJTIAOhn9X
btqnpSf0m6/3luyn5olhtT+vL7VnD2IENrNkowzitOzoAXVNzSTWnOd6ahBBuGZITAIe4GkWZLF4
fSGPGx+u+udTP7kpL3N6UnBB7Mm0mlbw9wviIIH/iOkwBufXGrkOkzAct2VPbmO56kXZQhuobfHM
BTc15MbMcfnVZHGp5ZMAEvR9f9Wlkn58qVt2d6sZlKjNL/Qjy7SCF5FJcge2M5/fp1q1HSIqtKpw
sPgIRqUlwQWrVrhUldFiL8N+mSNV8G2hkBG/B/OCUCkNlZ1qGsRLlxhOPUrWMezMKdq3SUuXZFHr
NHi+9GWV1zE9GANajxAS+9sJlNDkkeTntBB7YDbl+X2jpwHueZMFEAuji2G23dRT1EvDewTAYIXP
Pb/fqx+oHynaBmAJX0P5IOS4GO3dTabUeLJU+aQde/hOcE+fp6wBb8poH49LPuA3q1848dEFTnWC
3AX0BQbSixkLmWu9zmu1V3WopvD6IiHcfAiQI8kqdbxECQj7M0QOQRwY9UqB+lOr+BrDcwpGQTYv
+5FB41mqBXij6NLRL9mUABiGJGm8YpzleS/fuhSwanuSaI/LRNOCbtk7gT4vETvWaY0Jvr9Uuxl/
fd88WzzozSCvCVYBhfqRsFMororgatIBKyNLYpmpgmxH+iumKP7jZSu0cmbIMipGJMMfk6b7V9Xz
lSYMp63sU5WlDeKbNTtleckC99/Ip2hxrTcZcOICPuSVc+syp40bhLouvqoX4rPjlvwR3wFEum1n
axWFlKgzugeC/bsgEJqFCGKR3CV7XEH19vSNkaidggy+ZBYf6ZTtxZ1yEjilW2rm29Sc/KBKLrAr
ya2t8Yk28IACzD+Wo6uVUxoKSIOHgeT4/BpVgWzBwGtoN0l81ziBcD3/B5nz453ndFRFl63YMjPh
U4skQdnv8BEldsoVbaG9xD0OwUF5+N8Y8ZxJGorOl8ZAynKyzjp3r+Qtp1GGBIOt7+gNBOYwrFlO
ewTJbl7zNBp5OkZb+aup93Hm18xsqF+QQWjcwMMfc5RwYd9s4QrJ9j+adWZPRNdaeVVjiZqDS1/y
SNtj32ZKN15sB2Qht8A6zP3qqLbx6ZJKPQF4+8mRJyIHU6gAYbuUNdmBVw4n9MtD1IEQhNPFFMAK
PqRjdtRDoGkFGviYo2MOtpQY0UWTBgTQZevLWUhVhBbU/XbNIzd+hBeOLlLZVFFIwotuDxaWspbb
TEDv61Wk/3+8FOS/dhzkyBiklXhUVFAtJmdjHnpIgRISnxZBKw1GLx+kbdMVirbKieibXxFVaRns
3uP0s2MRp6lAidpn1MikfaeuYZgEWPxI6pMshKi2ieFmjvr906rcFiK93HOMQNbaJs+pqo7uz4Q7
95/QLff/tyhBKjUt/aOIUkrIBgM2QUuzvFqAXpzTMi+0cap/W3ZS8rz1oz6jThE6D/NLk98cRi1i
enugEiqya0SUCc2rLZCbAoGTfiAwGxRlbA2PjK6fbXrByDn0VwPtGvSRv58TZjmsC+CeWVV3lE0a
sImIvIEq2uJSTHguGHQ3yvU3ewixqC5YlalzsXXQh2j/E/N+0n5gwjTKCeB5E4LYvrEjuuUxEnWV
2pt5BFTfTDKpt4VwH97m9+tGnmhBopBta50hse3nGeIMjMgGsts7dVJt8rjQNoyFeCVzJP3WH1gk
IZAL9UCwMYQkw22GpULIdHIlwYV1lDkYvleChZfXhtbBizWXRhD4MuSb1oTfjfOUxJTom4/Y83IU
mg9127X/nxbCtRPsH4eZ4+pUiG9YaBbsN7QpAIPlzk25ciUc7ONn1x0lLL2OiEEcS4zxtjIauVbd
tZgG3bXXxt8BhTjss1z6C+BlxFpBp1VRLxU2GZY0OB1wro3lV7sMytAi/PUhoWlD+Ga+/yEHAjEY
yUiHuaoMKfd/WkdsoHSuTFrZ2U9qVNB4AQNdBf2nR5gSGO2TNSby/ig9dGkBDRWM97ndWa48sGPx
FY6FOjJ34RTxv3tggPmv/g4CV5mPygNyeo9ONJm82A04YNKYibAeVhoLYYp5gXSnZm4O8kZjptUg
A+SWzyOk3On1Q1QSA5Ab2kPxnECWDoLeVGOfTgAaOlPiXXGXgQgr5Xqyu4fMIq7C/bLzoYKEJ86W
4o8JUqvbP8iZXEzadrmaPEmEoqla+ekiilW6waobDkFE1lqYmlWBUQfaomil91UyZ1PJg7Jbdq9/
ywGVCt2bRBi26RL4v9yJwyR4a4uzmaaVrTTRbgOmg80ymguYsNfvxIbUKKBmZd1uKwcNvk8d0kzE
KwBl61wQKQwWkiCEHWR4cU5acAGbpok3PlflR2jgrt4v252THj30hVTdWHH9xLNzskXGKaSy3RIx
Uv3Q/DDbbblMvGDoyqfw7SJ/2157XtghN8NycOzHIhKbbjvxKjLj8lPCXO3zr5PDRWIBQ+H2qX4x
UI1U3E6vbK0OH1EhVi1PbUgeWjE1ozgqQ1AQlrW3c3se8tzxw3v/JiO/3mrG1ku/KkmRF1QbWDS8
OzjWbV61m3wP92vW8LfHNcgbJJ3sUE0PRDQlEx+AzTWlhumqapW2iBnbQvO5iV8d641P1FdmbPQT
6tB2oCC3vSKjlrVivYj9t0f21DwpLYHfh7jfuulB/QjvztsFNGIfiyJP2sntUBfv3F23gmAN7BSb
z13qOki/TrKdvDryyxcNurlEk1LSlnyV2rjAzWmx8CnXSpcYRxB4QEzjCwnwqO7Kg+LWATmjF32o
BS/H8JbxmrX1M/GIWPm0I0BVkjfIhtN8bznUL8ciuXPUdevB+WfkfyavWmGyDqFJkSXo28B2dC6n
CGm+9CNvscB5+VTAdSmQmhH1NbMGLkvEyaeE457Y2zZ+ov/ZB/8qQnt6aPtWFamcroaL12Mw/cH3
IfIwOmYdO8pN+MKD+jSBOARF0fd980hS4R8iKl8eUzdbdKTK9iOtg3zh050DoonTJYQkZAatCIN8
WGk/hyXIoTwvcXzXSI5Z6+pSEPsRZawEWMvavwEZsSijb8aqsk65ekOUCTmYENbLuJUy5pxJO4lI
rD1KV5AsIWIHFEilVPLXKxnmXMz3dL8GcR+4IJUSsI57YS7OpAJJyK8V73rA+AddUjGCllr7qhUY
qOMceIe/MHTZ4qwnyewh5HGMINZbXnmqa09Si9M53MEYG/twgHwCP62KpkskVSuIjcTGDeSDbiRI
rxw3hw28ImCucTCaPk3Npdl1ezXWalzLY8GVhXx3XsCWQ2oATembx88pFQVK0eE1OdePePSuSv/t
I41przSgo83oYzODfFE1PVI3HwwVCJ4YjGEsu1hkIfo8YvlWa0ANtJYKFRG4x7S0/0PfoWMTyvPV
HSaDGieJYMswQAHkenr+2AmeLq8rO3cSHm6IGmLZ6bZeCbkoPt+8JJ/5NRbBKpk9mADFen2S83fq
arLp18uZOwx6QWjo1aXmKk5177LgNFRiZQWNQT4bItSO0OW4eila40NoqptfIPG2BPNN2ARvzrdd
Vb3z/k5sNKTGevuQZHfQfgvIIH2T3Y5gj8eZWA5fTXJGRaxQ9VSwZW1vIHgFuIrFn3NGmOXasuNI
jtbXatdY/mvwnNDg6PTSKWBEamhRrmYF3QE5sAAZrv2JjG3u+/LaWio+TJz70duA2pXnIIJtX/ez
/3MbNH/9MAq4HUF92rBbecbR+o6mZj1J/pfwE2n0G8RxdZlBNTJUVYpPZlInj1S+qI+9wYD0iaJd
Of0zajOn/e7yrZPSVxlndqa3vt4G8I1o1WfNyLyg0uslDJ7Oa0GsbDWeguCAl40D53xYmB4nlLkX
qAJbE6tCb03BpNDD+nXtOJupNYitAaOFRbUjfBAn6A0/AJiKYbIKowXWLO0mPUhjByHqL7gqvgfN
67CqIRIrgaLQF6UtHSHH2mNe67rBp+cEkVVzoWOOGwQO3wr+za5B77h0HiszXwUqcOZvRxxwm5BW
Tu6qklq722OUEtHh7Au7ZaSg1WOazB8KJeFiFf3pt9ErEbfZVJl8dyBSu7RqvNtntgCii85jTG/j
yOPvYHWInPTsUmjfhAJlkdw7cFsDFQif/BySjiY5KmRqaieY5gFEkvZCW0f0MdwGIWYWfh+dQawl
0ZJhdUx7eKPuV5phkNwPVfNLTYoXwItJ5XEbZdb/P9w7jiYgWUwplCmI04rHH2KKl2ERaf35W+sI
pTfzCus/xMU1X1bhRMWglv8S1KBWaTEjGCVuBoYNQ+fl4w1mkayRiHtG4VH2zcWLsdjmBPug8ySc
hJKVNN7JHw4C1HonqI6RLbeLedilKJf3xxeuAiNPwDTXAgNK47xRwNuIqP6iDNIbDRz/wz4bDxZK
wovJGisWc8evdggyyqgAGx/ZIzNWXNgb3hRDMYfos2xKtm/slkOmr5qM8g8Y6KXM2kdaMNuigjEs
wXGTa009+KVGYUrku5i0YPPRir8XcKgjoOPZPiM3sfeX2xolS/AcHZJS2iqJpsMsH/42a7ik8lV/
SMF6wYpcgOpuW6foDBzG/PLZxdd7HbuDqQdrdlkOtYSDoT7oaoTnTYPBb7Nn8AqwO3KF5uqevXS2
qoqCN2BToUZFXZ8O8Q8uZkAFu9JYOE7M7teXYyVlgO6bVvTC7+M8Cf7aI35uVzJ/x+WpcZEn2AgP
cQw3oMD7mtjkbT3ADtVs1uTZ9oQ9+UKSAcht0H8/X3ETu6G+EfGw7Koa44zBvCKoz3mkfroKyCyY
BdkjM6W/OsBRGNFUNtOMyPbdhT5Id/PKtCGCdFDcUSGjD0Tzfyeckpp1ilN3Hx/wEY0JkQRbgaps
H7naMHvuzyxOHo/lmAYpi3YTi1osZTBC1NzqUI5iW2RTW+3v4bxLvdT+gBut5iDFHKb7y2AIEPCr
DTdxflTSChPx5uwxwqyessr1Hr1kiBcaRGDNvsrAa6iUBlK3IsbBDONqgbYiHRuacb6WceMTHDh5
O6xbt7x0pfZ/tQTYZylZLU87nC/fwpymm1FfEqK8Ppqkq9aJJ8CmQ00wwLGl5t0PDF9WiGpYRRVA
jD56muZF6s/xsg+ne2+YAGEtPNQ0sH52jRScE454TvgnYZy7ATCk65+dX9uL4Wlmk5ODwClIioBC
wa+AXGib/o2Zkgh1061fL2ONU9ZhbbJH5IkusaZVgAbhKjCo6JMOyDRjN/veN2+m8X1PqqzVqJky
nPI/aYD6ThW/44y5xD1+M+kyrn2uKZPeE6BUQ7SZbEVu4QmtwKbf2cVISGN9vpkYTPGXNcl+Evt+
sF6GfuYGaLbmApnlF1sK+/1aMIBcRg+Werm/BBXbeteT5St9TRbO5oQH2wPimjJqEkzJoSpoeHMH
kU7w2qxvdUgcjrVSuta/ldF+ssltVs1tBtyRWH3tEfb6pC/v3PjJQk6QdWs+DXrf4plSlZUfJULX
F0uZjM/XbsRCZc37Ww85DzolgEQCHCilODMKnCE6cRqWTsEOprETeIU/Rl73cLKTdq3AJPtVKuqH
G/waKZzN+PjrwDmsFd7SCeSP0fXS6kuYMvwdE/mY2I/tnvuTAF2k1IC/vn6HN2yCwNviDBaGodtQ
xVIDjS0KLcHXuFr5zIHZpzJL+WIRgx5BW8stptYVmdig2p8p08rpOjPmTxgtbsuHZKanbWv252F8
ifqoMWY7mWJ8GP4u7WI1Z/uB8KYH0X4Azzpyr0i2FWosNkDzUSyjlolj9DFutfqD7WvVsU+Jo4Hv
201dTt1n2aaWa3//XqG0an1g8du4Leos9H7eaHfK6KznxVG3HO84kGlmgH9zABc01b+mrfGmyUkt
gTVUVdtK/Bq5YmNG6DbKtbHTfAZts8sDp46oiYdsElRK4vh5hutc9p4SvK7l2zaxxRbLEolb2XVD
lJhJmIGMcEDAzQaTbVk2Jb4eHTwcUZ1JrQ9iGFnpCAFoPLR+s1rkT73eN9+bNkD94eVlrEnN/PxJ
dwIfVEHGKhVriDMPmmM6X4B2rgpZlVdDSCC6Nx0yu/O+QEH07k85sHSSFulzMWVtmuk8oNDNGVS7
s5s8M53YmrSwi9gECgk0KE2QhWw02lX9A0Unh53xpJA6gkLlxIAhZFVhdlv7mOkEG71VKYJlCRAN
3lgt1jaBgnfm/WfqwyzOKzf54vKiXePJLkZYCE+XCT5lXKo+6BgTsWjwYtA9RtZtA84ZProk1RyZ
7VWNauH1IECtMP9L11DGyXJ8q6ASiONGhOX+0Zh0EXLBOop+qsvHMwrct9Riy54F/IrbCS9zvquz
5NU3L5NFDeI9Hbmi6DPzS/tFjmzBwN84A5F+Au58ZAqSS443Hbp5ERpTLsinfStqk2zhFG8Jq8Za
NwpLJ0CunI9uvdZYlkymr76FXLesjOc27+zTtp6m7/7J2QgqlNf6iU0/iRvcX6VCafwJNrbY1QCX
VndDIFLNfnb08Lc1EY4pt5NDDBXLebDQ6e08CMG/OBrQNfux8Hu/tsFTtUAj+Q7au2hBwbKdOTsy
TckYspgRMzh+JCoGjn6efHsOleKYhTWBeM7wZqr+ll/uS5k2LpMNGOUkrYY3b0DmXMkE3US7wVKh
XEn2gfh/uRMsWeBMsB2xWCzNgIMYOtvzakSaF/bLkgF6c+J+rqj2icyfJkiehkzfLBRiUaw77G46
OT4MS3Va3m948k+83W4fCF9ks/EkfNeaSS2wtzweev48FMqqnsswr+hCheoNEkmmljTeB6C8ENzS
zTRyVvOU6taDi8oxLhnFfnB/frgzWgGwF6xSjxmxml9Y/eE3pvV7jfLV4C+j5R7L+DILjGTIJAZD
fWSdCjeby9iRBIYuuIDybPpNJ5OiDNtTEq4rMSBdtoKZRnlfedMgUZyTDTfDYsYDLqcKN59FcREf
Rtdd58EILGePAH1Kt8P1lZjU2OvZDWdo5K9NVWle5tOch1eIJdZkgMjxjzSR7xZf95ST0o0d8vLX
Vn9dS0sHCDrDvWvUYlagKaLyakUJB2X07O+ug/EPc8YEkxWVOgXDPaJkk1SvgThBNgIzZ+F903QP
+1Fc5fW0CsTF17SnjUUFolWr+gBK2jYOjXL7QGfEpTM3AnoaDeBxzhLiqLgezWeNUmUyFk2fvuO3
1lWsKYXgH8fb7GUUf2olR1yytWDEehrmr8PFu1rG51mPNLbLnnwPJe3cT0+KE7ouEcfdDhmvStEn
wwUEj4ugBWvrDwAnSP2NgTf4TtoU6mq9JocBh1I6VcFcrvrV/ormgNMznd+JCTHOsziFbp4OJOXf
yrXCqa4FWiGcoNvEc7Ljfh+k6UuHcKZ+6bmBS0GRVCi4XKFZqvGzZE6QU9gKrRN1biyXFwisR4wj
z/HFIbTumKl6mqBr2FvIQdtsz4+HRksABsD6CRTOnUQFPc6m3qJGcRGqIXyky+ml627F7IyUKbSD
ccI3mvsouQ6iqhy0SJadimpLtVTn9Ba3DZpblnY2Z1oRu7OvnnYDcId3Wmp2qBnIiB56vLumj9Ug
UtSuh12zavNAjqcncVUID3i9y10qu4/IYh7/u+fri5VMExn5sjGqP+5nLvvq0zoMLehuKhVxninj
Fk5wt9Jml2gnTbBSdwCTAfFDndN+27aG5SgDMpAg0/W3A2U6ZQcEhwZy880s7hrNQXLaVfRm4jMU
DGtuY3iBARm0jyreKZlV54MR0KxC49UhIx3CqvOBkQ2iZkLrwmhSOCAiaWji2HPTi4UaV8wDLItn
ZOSl3qBAejU140+lPGusJ94z2VWnt6M5ZOso+qAnZdwfTb1+2y3hac+bSsWIlbaqL+EDI4mk53IX
QuNmjl5IcToS1DZanx1Yn8Rf6meADq/+G/gAS8VTnW4Ms2PqEPqSMOdHrraS3F7QXwgtoIFi2a+G
xtoIfekAZRsfitqRTEcDsy6TI5afnvLZfMC96ZoIb2neKcm0kqvJekDxLeKUxd1nbv5cvhxT9lRw
EBZxF6xS3gQFeXiWiurkwahZ44tTF308DsOyoFHmMgMtwdAXDgUtDVZaKzJqPQ/gjFHcLDD5EK21
M0kkUkfvmziDzz1Iy2By9PBJAweajt7nyqGPzQGGG/jCMs1lzSWswqyw1/Pp6VFzhK43mkv9mILv
YRxPHnZ4DuGd0ga8MkI+JTKx1fnNkyGdNAGH8yP0bJ/98Fz+1R6pdq1Cwq51Glylu2JhRgXaEjJO
+BAZgp27QM+cy73QfvCcbn8+e7YdG5+r2klxVy7xOn2amFbWsXJSDDcr/+yBIiV4KWW8eWT4MKh9
b5PpNUyreirs+JTFu0nTLn0jKlb2Y2nIHY9EDuLRHvgIv1VoV63ZDUrDxCBKWyCaf2hqQ/G6C6w7
cmphRgq7u5FCoWuK/gapjv4+YMf2Sky5betfBUIKCqr11JaXxgtsEtWMint7v2Hb+svOa6j0OVqU
KAxr1nwIIb6sayfNhmEdoKV4IvU9DAMMSVWTxiCC/XCb/OIfYyW5RJV9Ma1aNn6q2PVq6uKWikar
a9JexkZQxcibM+oD3RANsQMKHz6Z0Jqg4nDhs0Mm+9Q3s50aB2ydPbTFrZsnzqyR61RmqBG7rnau
E/v7nh5iEKWWPpsjax7cOdtpqi7l8y3KRPjpfzE5iehXLEf3UNlYI/T2bOrZKphphz/cLjbWu5dg
K2B3oeA2w/zLwPn4EMpjTgVte1cHfwxqcwm7GP3g53lIJUSU7gNG4HE1/QTTfUQ2pvUe3qzVNPak
LRc419MnytIRSGheC/cirqKbwFbxpCktpS7UgaA8h6Mw8KvcHKpEotRD1v67TR7A0OIPe2zDBx4X
+4tc11iXYRAGBNN9VaUQIdAxkQKZ3rQck7jcsV17aT/COd7JOWjjE9iyAU89HZ+PxgneLeeIJa+y
JpJjaMyBCXRCSs/V6eUg5gJeb/gnDE7ZLNTgRbwqOeipcjkGb0Kc4msQolS+dXCxmhlDFQn4GZRk
qUURpyvFl2esaYPhfv0jTKSUJ6GIxyIxykVzLLqn7KcnNsAKpC0ZKKrkCA4Kt1ILOmciU+UPtDJS
KyScM1sm2pvGGHwqjbrs9rhupkykHCf6pHUJS+C/2FeRx/E5xgC/VQSKaoe8jP6FKdMXDXe8oE1V
8KR+5y7ivBKA7HZ4BZjhHej1cGNPMZFe0ZwkXjPIPuF818fq5mYYzje0TxeSj/a2/YdglHVX8UAM
lQdgxKVTWnIThAtU5D3p5W5tsYADcRuURCnlluFD4GGZnw9mT5wcaN2ynVMwWw0NKhzuEKlHACqt
2+/2BZOpiYx6XZ6ebZWmNzcYxX9L25BnJhXapR56sByrL3jxEy1Lk6NL4jhFutWz5LuGPd1MKaQy
+hBmVpR08s6GYRKPzzZhZmR42zKj6aEKE+4cHdBE+3zeejBaiDyjgFhFzhGbJcFxJSat4Alp7Ry5
wW3NPvp4hYv8jZtxLneuHF6BRtqvop+0NOA31PQ6bT7Gkpp93npP/KoRcgiuhBXQ5xIspgcXDpYb
AVcQQY6t8KsS0hNJSurJ8quzzpQt/6EtJ9JWOCrG2+eFHhvTbXDDIQ9Qfbmvs8EgdNKNtaZY8cYj
BzbZmQ2owuvkM57kdna5cVoPxq/6qztsttEhTnk17W63cP/dIdvYJRdzNWr/HzP5Ea1qdQ3Fpu08
XrE4x+z+CMPnN29sgw7g5U6jQtMNQ4qdwv3mj6V+a5tfg2WzPn0tjxBtHkImz7TkfhoqSvgabbNs
Vp7bkkS55l3WMd91o0jvVbxFJRV3GGpcTs458gMV2NZHPk0ZjZKB//qKsioNNYtMc0HEcg7IwHHg
Zgw8axPEkQI6NLpv0gWoVHSyBfoYFyhXYAHMqQKE90JV+h8kNXO7w4wD9WSNTEVYBPOMySS83hog
trI8zVk+fPC3CUAgYksDlatAXbtRXzkxY9h7k8A3Dz4/KBE2vP3wHEbj+NvmTOHTx9rQVC3atoEn
snh1qp5z8es67GO13yPJoJ6m1SrOJdGSitY8M/aK/cafZIrFCgPxWETo8Gi/sRMCQrYxt/QSss48
DRDHXbmcEU1wEgx1Caep1/MQl9YjVqPUIRBiDjSqOOXvTBO0Llixfnrk2cs6ZAQGHDrFcoHOVDcf
6YRyTjd5Wpxqx6ZS8dUltHiEldZYiVDjOr7mer0/i+EJsVwIhdlqS2ctX3Vzy2HHjXFT8zImHmYc
OqVsWflMo3UE+rbn7i6eeZBTSFJskJu682ik60LblUQnVmb9xOYYqCgG8oRfhC8a3yEV5E7FF7va
OUlEsfBvi34JXXWl9fFtUrTZGzf8is2N5ZmjVV6Pfd4skCQkl3VtGtfNC81Pd/dhBqla2g4sVDH0
2+afX42XlYVZqNEX/zWy/KuYRv5CbybjhUv2Y5EvQ1xiRgf3hTt89hhJd5EBaYtdWgfCrP8IyKKW
zcnrtZYULVPzIyz6/Hc0TKkw06cedtQYto7hnp2+mY/T9DEK2pgqkDhTqpb0D58Xmao4BptCGrWy
R9zEV0g3zLkqpSEvFs1fwHBIGvYJuzbh9OXFiLoWPHJBMGK+t1Bn9bWce5XmdYVRwX9oyKqSAh4V
U/uR5pjJqQ1GdiiAERutScVqtuD0EvfTD9LeHHqJc0dsEjSZ6FcTNW0BjFYcW3d34+kZiuWQHF8C
4KJ31AtvBY/jha5i/5YdnisKma4JAXe0nOw1Zc3lnN4oP6O6k/plBFuG3ItRO55jGHuzPve4S3DV
nFoCefFKYybOWw1y8AbSLJ9TutFxAl1RdomefdItMYrlbldZcoseNZl4Cx6VMyFwGxPfFE7fezNK
B1iUKDq439CFNAiGbyVYT+TbftKJMeip6R9yRXsnoDdkNRtlPToAfgyD+XZnP6qQIINMbDApPiOj
b7cf3UXbi4EGKCqFtPNu7vYtLuVtuuz0DgQoI3SVbmxV+7t0CcIz1/lLKJkyzhFO/oUYZgCYGiE1
gDtJ0MJHnWXjt5PglttHTcBsP+95EW0PLI6xPe44Y81SwWyipAILg4qFOdnqxWONp+flVR6c2u7Q
rULeSHajsOWV/Gfh3Xzk2GYRZ1BU8jkkNYmS9JhKNBOf/VjAOODtPYhTRgGiKacNW6sZp+gM9At6
h+/qq9leMZv9eViEG1qKSSHdhLxwvsxxO22qWUPGlnswKkOzmF/JdguQCWRcoNf3wyrAj1k8GT5Q
ClZSahp3lRQV52c2vuWv+r3AtSwh3+XLoH0zk/KQbUeM6kuGknz+8/BUZrK+1pzA6l11z14WRPwe
73AQgZ3mtalNhBx93j6Nm4WujgkkHWv/OztUk9efq6kaHkz7kLcH94jdTgsFzZ+4ScaRKXSeH5Z+
3AkZalh2y2HwCi6GRxaHmTpi1Lyp8emwmbCW2+Ijn14Bgxxk6zjf2gZN1YlfbrAj6hw8+pvHgK4+
HSIhL7V9hTDQWrFpSq3yM7uT3kHJTTBz6LH+2Gam5cqolryWefR1jAw87KMEmTk8hTlbmD6i1f9v
erXfzpixLK28skkrnEv28DxgpoT8D66Yr8wLR3Zf3i0W0SlQ/7FJ8sTfLv2MN0JJ4nRSxxUTvkjL
waauQ/CQxes8M7VdySCd4Ft7khyyIL7b6vPO3PwArojIWLH6T3gkCcFKvdpaCNkIGzSRS+gKcK7t
jeJRUhtjbTGA3/HEOWgbqWi1U12a46xGmFKSdKZbYGUlTeRRUvB9hJ59zMt5MsxiENFgXtUiLZ+3
G+E5Upl7PI12BSWqMjWyv8gBJo4AHU6tQc580QpI3EQCIGd+VvU9UnmF04GX7ImXaE52wRqLlp5n
NWcNaK+0ZPezqI/NPulxpeqP3Kjcua0csbO10gzhIeDoYNuVxgZUGkIwPT0QzZ/IYzm1jkYrb/Fj
2+4G88J6e0PkQwRe6kZ64a4SMP1ik0GmHuvJCdUNcyVszrLozEYPufZsQ3zCaaXu7qpWfIRw558r
nx8nqYQ12l7cM8GkDghxFg3PbxfjPpCsr0zh8vX61gp0X6Fb/rQ0Ml25uudC6BDqxVvS8WjkHENb
tT8QatephRGhdvt4EVDC23SMPHg0ecON+WQn7hjI6KYe3Jy1UDCms7pq+exj3XZK27111ruB4TBo
2o/MgMKfEf4VnY9CfCY6iLJ+WP9ReMMup1catqsEcIsJZmYDsay1FEp459U45LqX+783WtsUxyrR
jl0X8ta9djhVKW48StSCGhz98Zl9uqkaBL1+zS7H8KWlkAHd1yQ02XK/pinxs46Kz0V5UxxZlF4/
pEiSe2jVBZsT7bMLxiCKuLY/cXMrz0NNhAGidqItyklxljMVFbjfA5RZnEY1JbVTMHJjJa1OOsYx
m0HUQdc5SRqdU4PG5SJFTvPkLS65vjxHVirylqPWbK4Hfqm1r4fhnbF8umoGJ3gpm4GrBW3Ez2zS
92emFj/ynSiS5qvDGDn5/a671/XhF/zWBQMlWJUb5yURQeJ8gqlb66FstEZ/qViKAThJk8FqsQWz
ZSy4tlVFAJt2tEdflyeVghx439c1iMYagxH99nQs5V3VWfHZdtQ4EXEyEWwpwNlkpz18Uv9NB9EU
7fkepylsxblHm1eVmXJdfJ6Co3KvJ/VLUBR6D0DGKkwQfMXy8y54iz25RLn1/MF+moVtdkbXMJ+a
6SV1H/ivBUpIxFymvsOzGKjUb701Xy3Mw6RnpkNI9c23DSw3Y4rEa9dWvZRZvBlRagB9edhI1S21
E9RwzA/ia9ZWDyTBEifaEKw2xjQ6kagYCQWYsEoDdpPyXqBODOTyKSLqwB+YEHpqItkemZd4YgrL
7mr66hZTgz1JWL0+MRBCiSqN9y/JG8yKBgJEJOGL8grgHK5Mtx8JLj7Uj+6FcNX1BTNagOT+LL1W
uCrwCoQFTz2xqnaCa0jck1+XsavbeLV9O6xEwJKiw5TDDVaRVhFuoRkMyNfAQmF5gGwCIrTaKZHt
LoGvA/l5lwZZ5khrtV8d3mJy9XAEXjNtXL+CnciKHTXvH58O2jbE52teu0AA3K+CzNMlD6GV32DE
uzRgyZte7cpxICHlgdU/lHNUUorJ1Rn4lHoxYifjRFCNXa2Z5L+NjG1fdDUTNG37UMQ/DdyIkWf9
U/EAVLmAvS4e1/bnOW/8ami/q0iOnCEAIknap4UqbaC3doN5mKSbxGd5JOam0WWeI+EoymfJXbfm
qhPu87XrKhkjGAYhyjyWb/P9n3xSrT9toJuCWZbSot5R5RRurfQ016vKPOjhS8wgFUHdc0jcKxpa
8GrEMX4cszLgKjP24x20UutWiK+6ysNAfBd11Mj92Dh4s8wdktfqcarfCgqVzdsUcs5nghGiyeFT
2ekhlTteitsF2Ao0MwZ7Q0Ny4wCapznca8hqbux8tfHnjiLwVoKF1jn3z1ElHbP1P4M9gbWU6s3a
92b5V4jWrAey/ZtgcG1b6xEL5lNp5PQucpdyKVbspfmlQ34qlPUkVqJUK/d7uUM2myWubDDdTJrD
5Ixk6+ZavLzD8Jp8msTICRTsJMDHu7YWx+m5YJGTH2EDmXFIKvQlUfyevQb350Tov67gKcsLtFMV
yOdeLlIgO4mI4IOqR7wvgiwrlppwSmOhg7CZyHlTj95+SlAV8D9OZGBxeNIjKr/f9w5ooNS3AiqU
GoeX5nILsSUD+Xx1poqEuviiA0e892PdrrJIjHtlxS9QM6vekMIrPh8kICDtoblT40TL91ga/qWI
dZa/9m12qZyJnOZdkUKRA5R+c12w8cMPUePnta+AZl03z+bCCgUQOkqXZ455WpugSXB5SBW0STZL
E+9BUvsd4u4j4u5u8rkqzo0Wio6QNefI5pZWZ1+YIfGMOdLTYQY/wxatSEOftxCwAjdLoqCpaG11
KUjDLcQ3f1TJLS0+HgVOBbNq3Vx99dGhgayatNOyTEDGP7Cey6k5I3I06XcakSwq/VUtvE5jBJI8
nOqb8wySAsfCGdM79i/Dl300I/yi9X3ZqlGvm0XeO3Gf8UXyQFh/SoLe3yGnsBd6Jz+2CNHnWdzU
qexnPj0vIyCYMzMdCowyF3MS+44T5fVtgfV43Na9jiBxGJVhvMz2Kl18olrqAhunzVgHBhhTh9VQ
0FM6hTnJ1EKF6j8xHLuOjQuwUNz/WXR8CQ97m31FNrN10Dgs0rjkJW+kd552Rv1LEMgFAt7oxpnU
soDR1/vCdgq7ruqJrEZMDxlQUQIVYK70qteBR488DWqrI9BCHqVoHik2wsLO7S6977ZA6m9D1G6I
PPyerxZPL3P1BWlCLeNdCnv+ppeQMKqT7o5eMqgSK5YFwdiQDep0BZh3h9AwcIcIjgckpJ7OD7/v
UhhgQ/7mmvTQCu2QhUqP0Xqi7KNxej1iwZvm8TX1LFOJZo6s0Zzv/aFYgPp1neb+KVgrNQ2s8IfY
DPIlewPG3tU8zFJzXiasHbjvOSUWkqmlDuWU4qJ6rti0MF07y1k3OTL5vIwDYR+khhoPHbzXtDkf
NvN0hU85HFVtGKre73LNLHe0ze8TZEWIKBzdnq+vIIEvr2A4douRZ60RiS5D5tpLOsXLsf4U4L3m
wjjJds87qAYyR1Ze6/4fO85ZxO8P5l2m3Ry9TBleaGkwqjefUnqqN4NkC4Ycc+osVoAzBo05/5IR
oDZ/Wxk6v8Ki5F1ik03LsFdCOy/fmjYTkts5N5lpLZUAbvO/al9GnTCxZuVOhp4SnvT7epuhWewx
iaDA7lcoRIVBSBrtvKSQQT5MLpU9rq0HnDMCx5fTGzYRr5R+L181StO34MpzI2CI0M9y8db2wc41
k/rXl14HSPpowV4tr046VK1I8HcmvvQkg6VJEjIY8blfKYFghmh/pC8iZrtGyyUa72c2Lxy2slZk
8cfq35KNYpDWEvAhDjHK+7fKi2EeyuDV/zAITop8fOz3j5HCO2eG7XlI7ITp1jrTV/c8l1HCeopU
HrzBX83HNkbDuxOA3IvuquJ4kFkfDGZpMdwh8pRcqo4Cpi4QMr7K5xyBcljLmZlajirUztNDX2Ak
Zvv0R7AvJAeLtfISbq54tzhORU5cGwygkswcE+6uLnEBFLTcGec4dpG9GsRwyCyk9h/3VDNZG1m5
7EtJcLMZofV5Ai5Ewknheqsk6Fublyt2l4TIlHLab8QGJWD9lAhLPMlt/MgywIOWOEqIQpunZD5S
knBJ2mCtvEU295e381j/d9+Cfvf5uB5jf1/FHS7XclrAGkZZswMbPMLtRCEJEgmRUmHD096bHULb
TblEWyjySQjOJleTG65EBu01xiRgxKAep6XLD30S2zvuMPMZf3n1315jwGn0WsmHIZAZY0phKsnY
/zFoImnEMoLXd8q5sNXgP0/u4tbWxmdStV+Q9/fvBOiLWUicGsppBpxrHzEwM+6otPvGpdBncD/J
YVCy9lmUouvcql6RSGSYPfQFFjMzT3kIt1XJEBl9YjiBTaOsLc8zC/+KOZYFrfqc8YxP3crlsUHi
d6tcuWkDCTolgeV5K/XOj/VaY0RzaVRuOxMIEziavqF0gzWH58CUHg1v6imQQ66j3Bdre0FFQijk
zHp1pnwGIP7CXF0atJUu8se4ivcds2icPzH5MsVbqEWdZ27nCNAvj3S6myoP4DuymNQXkzoRiD3+
fO7gr2xOgFKBRA65OsUei6u3gb0/EOYLYF0Av+kt1wo5INmlRr37F+7GXabGmhqkL0JNqabYH/Qg
nK/YmwFGXhPXdSVbJyfLBrhERJ4VWTxjvacF6f6f6T/pYUQQlNpw0u/BeFUMECydq0PVv46ocg3r
PyK3P08ZlTSyhYw6QfWbc4hLQM7QNoUYwij6+SdQepvbt/AKwtNdpfuyBvMJf/dw5XwRNH2L3nce
0YXmreGu++CPE8Ip9WdOrPt6RfymTZ+QLDe7FWHWOVVfk1PaRDuHhmoWhiZ1pqNgKkHmMogxWUiv
TMWNxE1E3TI9TLiyzr3Xt5RkaqJLRIQznuOPRGq5RMwe8jdVeJ8Rid78fUS/watcocaD33W+Rrux
f5ZDWTCAutPIZG+zWlmwofDMxbvPLfsduaadWNXMlflx22jE9+7BOS91R/5/8pxuD3JXzXrBi20J
TZEle18QLo8Uql0KlYPrT0i6Zag49RFDuwZatSD78hWLQakxqY+CrQbMfScRqoAuqZ1pKSjlg6+M
Cj2AAkN5XCPyUeJSfnv/QNIJjHWr03Y2NucxcWtWoCW9zEG9Ah8iGpaRroKjxP2ucrHqFR27BNcq
4vMqXs6VI4X1L2xKetUmFz39ndAq6f8+7bFhuesB5aVPNXp2cfpqbZ8g4rDzD3MhAwZAed0zez1h
GyevQ8ftqid2ChDyJfqlGP0kGjFKemq/iihSj16+Z8gpL/PxtE60apjIhFBMfbhQHl0OGQFnvVlf
7/bK9MdD95fKGL1iYB7sqSgW7NrOVnLPTPwq3PN2rAF/DWMhMco+GzNjR/3i1l8wgYZEjUlKcUHV
ExhX9J1tQD34kj7gJ4tgMIMg7Vst2lvnRpiBm7x+JgebF3v131vMTjT5LZHM/qwz5EjFwduxhG2r
FyYKu56DbQFE8W1pb0a2h5q5wo6dMp+suV410ZFIfXCui59/SRWf1fLaGklSncjXTdjlMQJDc9/h
yN4DTXgAe+e2JTiiVVln7kYDPhx2ewrBri9H1mIJyJ/pkgnLkmSobfkvUzOIqxrXm9V6yBIF7eZG
BlbBn+P6SZhIDb45GXzAM2C31so5uXlPdKXkdRNwziB6l1RH5a/J+i8I7lcTLaqL7B2jhZbc9Iya
4x4FFUw1XAiHbvA1oMSspNwPyl+7jBaf2vnA1awtOjeiJahgY9bmjQZYk7GpS3o0QhOf/TC2BzjF
8l5GTxV1UTaXmDOjsf/r0l8uio+Cmtq1jJPyb8MHQqCU2y4MejoWXwpUKgv+ixiYNITFBd94joFt
ruBR52QVuGNejoLI+Xpizls7txSVi9dRDD5HT18LIyOnjFJVwg59TTZgslzRP+j6NdV8PgLdIm2s
EVp2SqooeQSVU+gEwXMh4T4pLSFWNY1U5KUi7KvTr1PTyystaW5RKBb5fatiYB7Qgdl4aMl1D/Av
MhDidHWcNfAjhrRZ2yPLCglquMaxk2pgjp3/WpqR0ILebkl4wwQVgwO/3J+iv6sQoDV+2JWJgC55
CEfeOR/iRFLnOCP+SfYsekbZEceHtJSjRwl0u/HYu+OGToNb4D1MLNxOYGUu7Kt+gAeFUyQ9L863
rAbm1zzYaA2kks0iAG+wnb2sSNUdRe+phtkybmTadRZHhY3YAW3YdjJCS/lewTVgaN+4LhhJBYsV
pQurVZrWVAFbzJ1mh1hwmbvV5/OcY+0qkG62j/2YZzG6k/UR+Qh0jNOKcbRsRcJMlNU8MTQmQmUx
L3tAUtwHrWfT5VxpTPml7wXwA2roC8F5pFeErYlkQLHCjL3BuplG2vMfbHt8BD9Dao8hOR15orTn
BWEVDj9CSI5pXctldkPPN/fNsLUpnQ+b87isJOL2dSGfRqjSxhOEfP133jjIKPZyZcQpWRa2u7Dy
2C9UroOVkf8CfkS5+HX9biqwfLZX3+5jePYvhxeK5aJkbdQpKtL9GjJFeiPNJFpKM7gdm1Oo9BcV
E3wLErufZZQJCQ7i4ZXRQoLE1cGkIyZMa7FywrMDrritwcSeUbAjTIuZyL28HXTMpID1K8UEchzz
vodE6lv3SZSlKXUumQHeDEUWtdM+yRSGy66tqOuUpCHtVPEhTvRuQTodt0tv6MgFnTFMMq89vFZ7
HMz/XrIcruN9h3Ps91IcYfRzGomh/g3e4vVAJfW6cHlDSbEdOyMjSSICdlT4mXasJF4x06AZZpfy
CJBaTbrkKQjP0vjVzMKc8dPJkv7v5aslkqwJMwZSFfKVtGKhm83/kLB+0iwsI2BomBjmuAtitLV1
4gLpBKumSku3/L0p+2o0txcJFj4JqSfXDq7FBSlNYk1k5vi653qsbqBsLQc+wSEEs/5BYpd8e67P
Ux5l5zYXRoNSltan55uS1pYNPY1O0AvDs/DeEcdoNFxQNkc43xEd7Pywm0BulO3JqeERqorUXIWq
H4wzk+pjoG6WD/aRxo8DCt1P0od6YTu1VS8YHyctYSTKpGoNBN0WFmlkUJluuSWNrqRVmfMIaXf6
h4WCyHsrK+Pv27wZr8kav+FH7RzgjijlzbJCgx/W3oJqIdAVfCTWGPSJ/DmtymYtVfFylCDmgv9Z
dxjsdlrLX11mKQIRJuHr97OsV2O9AYfkHr/Vvw+SPGLWgqZ6F5nd8NvgYIs2iShUuDigfR3X/8Bv
yIhRLpVWSbHxTLv18fsAN/bMyE6kLtzUeYdJTim0ipIOwo6O3UPsFKMRbhysaBdS7nJhXb3Fn5ke
USrvdklgdStaWo74HCfAoR1Oi67AtTU6spKevzD0XhBp2BfrErZV46SeMwmWuIxzGyIMwNvlTdoS
+cjJM1whLRepefj+lWe7ODzGOG9h3llvrXUvEFMxreTYVxENuySVX+MY29BLpmoeMPJl3TkkHScE
QYlwtN34Y83DXKrlSCT1HjjFzxYhkd9v5yJKt+Id2Q8a2cTHU1phPsTKnRpyfm6NhLbXkWV/3je6
4jJ8ZaU4iW0G5Q2MlP4D7LtlfBuQ1SfXUaix4VV3K2r0aDNLVQ03G2Uqj1PlwqKC17qI3MgVdIqc
doklRmL5l0ZUWAar3gCqzzloBZCPq7HbwQWD/G6zZjlZjBzIBRGme7WVcMo2j1CPUDdKhvNTNiRg
cxRuFLegNW/KZKxCQd7b7dnkxqPfRVuLtZxWGVDcB3gJaz/JLXNfo3e+8TjiZuvvt4VFTTffF5mz
YieHiyET/dMnJ8DYyqQ9x0U9CtMzKegBrjiD2TXzZWSKDMAgguHC9gvwvOeuXQeAJWcocEkznaY2
Iit2AlW1QfDWdZYM4iBXwlXWbrVW++aNc7BWtf+DFg0cq1q6inDaSw+DxGPtetXOXp9Hg2NDVY0Q
IqHJ5fiLQsIKlAcvAG2HZ6tVvyqzqEu0m1D4cS1twQeZFeC4/3Zu6UyRYLvQamWlHBt4DH0gvZIL
PmmYJOdrIA5tyVY6PZMb9pIq3GF+dil8x59OvB/SDeo5y07leBsW8gk4idbBvTWHEvrkEqYJNeMp
mP8WvQojw428EkEBx0wZ3gv7kG53vNGaf5lYEYbv4MCkUVwIeC92B4MCP4DdmQeir0V9zUcCQFXQ
8oFwIVeiHhkWnDSl5OHD8jeiE2QENPrC6Jbor5g3c1YEzwwej3To2ZhrYRzGnL9BNmRGDqlVs+nk
vAjD9sn3Zsqfn2b1zu9Sg4g0AKebTeWx8cLETi4UdxqY0N+qOl1laY+08QKkKMeWfSlxO3GgCj9q
jtyFgQw0wGfLQdVRErZ2nhc9icCf4omCLbOzDtYIhIOEsK3IcjAuUYEuX1iYkf+iJ2V6nokEsqRA
g0FTjm3NUvn4VxIKCDbbCJw2rpx7hdlSnrALRHjfjGyp6FV7euyzGzWC2L2PXCa0kPzG/MxHfr33
Zzzt2oK1cK5LJEsn3apZq4mY2ufTRVQl9HJobueFosrz2CAx8d2wi3i/ZOaR/P3mgh120zxhYzS6
QRr96DBz/tw4M1S/B4QHHy8bC9ZQifvgqqOYh41FoOhL2Q5IAnRxuTMBNjNxavnPdk9ZFrd+gLiN
ZfOP/eGXH9mX+joZ3mvJl2ZRxOrg82Bda+P1HqQFzEo8/yMT0C8HoB9XLyknIXLLYGAav2h84AZU
/TqfVq8ivRisRmXKQKAiMjViFe9VuOr6JFpP+JSJUDA0FQraC/4Tv5+yoZMDM4ULi7YMLHIhzXPK
vgMkC7FpN9LfQbsKhnPPUaBpy9+WMRr3vPKen2ZNJbMchKXObPnBOeCqfmLsMIOJC7vfD+EZEmsv
y2O8Nyn6qWv9qIPgQ0i7SKIflFU0wFqfzvsKwG4HvcB0Ib4o6PmC0SPDJd43fFnFDVr35Ey3Zmpn
t4SkQHFRGuFdRUgQ+5pOVZH9O4/ZfdE+b3VDPDzWkCuBRJSdigco/l1yX2sSTucpdDqyuKmDX/Gp
T3Wb7aWBZIiKisacj9+quCo8yEB3ji7mb7SAJ0bvx24DcVrMv6fJS/u0sEzUV3sWD+qit5Ytu4Ao
ntFXtNITnjfu9pIvHU2vXQKbf7XLdzPNn0lA8othffkZURGtSFJAa/EtwGFy0iJQHg2CpD/Dn6kO
wP3wLqVwgFQlbCUAsCqw1R3b+hgtmoMcpFfuPYXW9t7bvuHAoHyTd1JYfkxDecaXMwK/rRieCQ/y
MYop0XPGceOYnTplreHPH5wHPOS7xMsmPOrg2SnyZZ/6NVKF93aDIboSgegR1FbhIAy8tgIR8lhd
kNmczQVJMV9gWUbk278LuqByPp+V0eEvPGq1K2orjsaDo1olFBaswj1FP65rX2qeUqANC/sPh0S4
vqfZgpTAImtrHVsiTly7QykJkOpHJDbh/zznkcEogL3rHSZkRfZQqTq+kjPnTQa7T2yVmIjnQJYo
3wio3Br47zZYAowFoEWL50aw2EKctrVQFBwRfVNonlCdR6QXCj99Ax9SkE4WrceNXL26dsuV6myp
Yqq/PdRsswH3zv6LQ3GgANtZrW0GUdxd0CQR+S1vmvPxMQKL747Rfi05INqUPOz7cPFHC/UYJTbj
7nuLQ86nErCabBwMwaQVNw1KM3QNaVCL0crS/j+04+r8iZ1XQWg3sJIyDiz+7kx2va9oMb6YPGe4
YoT/0PeaIERnJVMiP95poFKwEsVzdaduDkF825w29eIsS2j5H2qn3PRscwe2tDO7oWO4WwvDM0dc
IdrC9tlxhLCf4iHnLrwCeviAFk7YkMGRe01sumnROvuLZFPzCfwTRVvraaf4Ecb55hURZqo3SYCC
O7kJt1Esmj2KL/SbSG/w+HI2BMvZm21UWXouiPa6EUi4xqrG3YvkJa/L++8BUkBTcOFoGeJ1Hdxm
FmWic9P01z+E4TK/vkZvfR+z/OMaIN4friHYulhPTy/hDv6hWl9n/e1l/hgFYZou69pmZ7MdjlUq
xsckB+IfLXnESdgGUebhK4vyoWzF6z+YV3KZgsXRFshY0EQiCcix4qPlwLkvjIi80qT0jrmX+Q20
D3AB4c5UE0njpz+7yA+JMZE0BYIWlGjsCccRqDWnEBemjoExoD37009JPjXDrRUmiSrU8ctVoAuv
4RbSS+IDRarx5f52HQqsdbp/r1UAJY6bZBMG1lxMVwsWx3+fLYkGJHl7KzFPfPoOvk8mU0FzlPrX
7gYtKla5XTnrhWuxhTcp6KLIA3Disg78SBNFfqQ+/4Xo1Lm+UAKghZCNQ7jwo8hFvgOUpNqYDniF
4OWPJ6J5Oj2Q/vnHBxs/bCbhkKEttlBXSpANl7DNQX0tRtVdz/nR9eK8cnvKftIaeVx5mwU3sYvY
yx+qnmROijv9sdBfhQ43FMkGdiUAGNgrGwor0Lu0NGZGk5Ox2/0S4GQtLMSHj3nN9kSh4AINuhlI
QXJ1j1YYPaRLpXSY0QZMMnUIp4GaUJ+LIo4ek3MEF62m0v0jqqTvLpOfSKDXJ2CWyFcpq/DoJdJi
XLskANvogiQV5aO18zb9BzxqZwAcXb79eXZ5duoUrQQaUzB/OOqWLEXTqTSHxND0ub8TFVA6cazV
b86GEFNmlUkEERaIJiAqPWQpfSZSVhSE7x+U0hjdx3npFxnHG/ef3cy7KNgo4RHeqmtg7arIv1qm
fp/8aZ2JDtf6qdw6U4Ruj7j2AcgZ4DHhkNiGIJVTaHTVwTvBI33mL81BLSpmq9rNHKXbspAmSiEJ
slFK8/WyNA0f0tb9EL9D+5JF+9Vf/6Efen9rNIhWk3La5LXQ8DwYFB9itTXajBqb5LxsjyanmxPK
gaGrXi4aCmju4ffQROU/YovLrr4hrR1uACX+2jycr6GrgasrHF5MpuGT23O9ieWU4eexQnifrJEf
O05Ki7sJMtb6e3cysimIDactaHfMZ/MHxmYDXC0NCoL6Y8IgDuV5MxYGbiR/pI7ZYzSBPUzBIKvZ
0xxX2zdTlQ8Wz39THerpkGgbpu2LTMmeAGMUHlNVE0gfqnrLlNcgDJ214W4UZVJkBfXNIArvJyDb
CHAVwivTudKutbTW+A0YskanGz4kvYwfJKAEJtmIF+N5LALiRXRPIy3n+BIc9PbsiWzuMQBm53Yi
US0gTJfu3gbwJpev6MWpi87B+e8wu2id4EgRSat9MMdgFwGiI3fsS3z8XdnNqOAxV3N8ECXsIs0S
iUSzN7ARVTgOoBFal9ga5LIo5IPx9fHr/LN1ElcnC8l/HBkF80ueDSlhAx0OcUshbZmTWaBSNtRy
73heVTY1NmQA4v+8KvyL71Ok1VDYkv8fQryZZHNgYPIa1FAAGU0HWYr8wE2wxb9xJbUgNbWg29AV
Gz0jXuufcj9fOT3oi3kjG6bJEiwnssRueSlWYVTF2x4yYCu+By2SoceRMI0jp5ycAC3Xqi9W30IW
jcz3VWdh9POJd4h8Ql7raFEfboZ3AeB5yfP7nLEqlSc958rDwXArpjN+DxFBb/21f7Xr4Tb/Pz8S
/tlECt1yDbdzFwB3ITRjJ9mNTxK88E7zUS3dJC/8OMvBNx1ZN7kCz5cKnWCjWCulIxr3vqqq6thi
PzC/akMWn9XzpwtqfKIh7NPzKZoTiv5Cm/jKrkIw9yxgj4rkEM3wI7qmLHjEn1KaiFXMVbyMwD9n
6BenjjJ1Zie1P5aZaPN7takWmkX51HvbMtSyM9BF1aKdEOFbOZwaIjfIJyhISd2iVw5YKTmaSfCw
O3qrYwbZPyJTxcNPbUv6pChijbRMIilVhcdKsCUimVO+Z4TxXAYvDohcnr6b8GXpvP/iIrXaO3Ax
jwPxKZkR86D8rLvvNMCC8sx5aGJ2mq7w6tneqSqU3WdWh2T0AZRj9iarCOlW3iFF0BHRiCDzE3+t
cBSO+raFkV6osWCFJdUg1aJ195TGzDpPJDxqUxVunWzW6vWXJrq0t+mT+wqTgg+1oOia5J6KF/oy
CfDtY2YVA+h1jYGhGOEvtBeuMMxDCQqB3B+9z1csdIUn1c0oiMNfkUj/vak4nVgmBBKCqn9V1yC4
mWAX9XkEUp8dXySF7YSoQK2rSUofEhOe/I6l9PcjKVf/MbdjwVGle2NdEGvhCAI6WGdvJQk9jSnJ
PSkVjhIra29AHAwtovZhEPVAaIelyGf6plWMC5gQzjBXE+9IgGb+W9iehOnxHyBsG2TssPt0j+FG
bwIkle6CEhwqiQ9FOBbC2t0w6gPMBDFMdMFE587b9b1zuWnFzY0oeb8qM6seAgwfegudfmCIjdQE
bqqnapL3W5VwomK5uxzJpbhC6WposeKXnkGlmpSNzWhDudV2ZmbNvECrF/9Bs7p3c/NwzYyq9UaA
l74xO14IVgE4x3Xm0FrDaoIyUPoIJJgiHmAlXZ8x+7v5FknyWKoKkBBiRycKXvBIa7d/fnlTn2sq
k8DfVAldCPIfDMgoq6yXZ9EBHfUmeidm3LYQv/PqLEMet/2vnz/rIwXkJp83bjVsrRJKEjttsxSC
QWNxPROkb7oa0sMCSPAQGK+1pkUJ2eVuOSH32s01hh9SGaGQYgrsS1bwWwJ4bXFJq7SXRSqyVg4K
TfrJXan7UEZZ5nP48GzJsXf/dm/D/uzcI0lPcP0XP0NilDe+wbV7HpLsl5knv7bAmUr+x/UWCr7A
IZeN+7KDXoWKRFrw5wE1IWy3YbFNLD/535aLTTJ0YFCywZLHakwUeljoyrF/e21d6j24s/uMZ3L3
lZHDGmiVmx0EXCwusTNzKj+82VRwM3yVQvyhHDj6/ZT1AGxqZYZxJI9ogoHzckG0W545VuLWI5qY
cxzerqedxz7CBMIZxXyqO21DFpTeaREjkYs18WG99T/OqvMwGh48UlZzrJ5lT1iidB8ATilW03it
FbkRQkT/tidlWgguTPv2y5jzpWw6lNcN/YZzclG3c73V2Js1jzPt45JQlROpZjMFKvusZXBUvy1Q
gy9rXcab6Ejvec6kBoQzy0lHQYIDwKLtkBRrFloqeh/ZMRtyEJxbmrOi8S6Nxc1n1pCxL3D37gDU
v7eC+mldLhQ8oCCcmzauEuB67c+M2yTPvXYzn7x2SIcPuMm+i+yKWF1Ua6y0aKIT1+Nsgaf4uXvB
rJPjAqevW1O14DvXRZwEL3Bwv5hwd4X7xjIqWYJflrKfHRqjIw64rkrmKibz77d/rdaxbPCQWTGA
ZWwVKh2bWQ3Ko6su7e3oVVhDEqWE1Ur2ZlXYNY+QY4CAhnwV84Sx+kBGuIXbMs8fJ/cD9I/4GMBB
r4BxpGeDEiqWGVgpBw==
`protect end_protected
