`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
jyd2KlKldZVFYWZrjgNpwzcWF0AELVTC8GKKbwBhxyx5v/CHJeDnZSAJEQZ04aa/GrZxQD4uprAT
mZBDuQflW9q7VGciCc/xl4j3Qi5ERtHVpHKoNJ87chbgRDVefGjzFLaI7JxKlNoZGSsU3b+bzI6i
VMlorqEnMwPZVSsjTtAYmNPXL8Ta1Z2+fxfNYp/cNKYIZm/QHJQTEXhrGSjnQ2+lAyAE4lQjRnAI
k0ymDJi+qQpQGQWVjijVKEwXp2F2dYBB0M6xT/GO2TTO+1ZAHKNLDfe+oDypyDmcwsjP7uKT0VYh
Oso87+YXZ89i5N2x1bp7in6xJFyXIRaKtqJvgA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="8OMQvdwp7lt4SU/N3kEbt2D+3+RxdKRdpaSAeq4+hPM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19408)
`protect data_block
AxWoYSGmESm5as4E83bK4FK41vQ+YNrFRUZnIHzwl2ixoCfRyIfly9txfUuIStJdTwWFAme5rPBN
RWCdGzHg95bnh8KG1edQXC8n64UAOMCiplXTbxk7xr0ErozFBVim4hoIc3IZH4sHvOfUuwCQwZDR
j+7pCqNKJtesUf5hvmPn3WicOLre7LPgkzo4Cv1p4tzRdm9NAmMI98JmhgK7ThyzK6alXUBWWGvh
5Te86FFWR+ATKgS/jtI1SQmSLt2qMRsls+3NlV5USkiES0X+3FbETDPwia1dFAeFzAd0/2OZ4LYa
VarCpzq5e96GzaWHGIUDDWPt5lY0ao270hv4j7qbSUDuD6bSR3bbjz1qhm799DACgb+F01dgU2hy
B9jCDn46WsUWDqta0r3bedHFo9+IibCh7sXddKUDfP59WQ71fDS44rU0Sf4Mcc2k/fiZpITFs5mt
/1XpIPakQC02J4m4EgdXVhkT8U87U9C+iou7S4HdylmJT/9bXPkXJVgPIrS977R3Y1/20xVUQnWr
aXAmUPwwlEYAcnCh92bLVj8NToYm94znQyywdX+QsD2jq4tE/4Vkg0V/zIuebOUqCg6bCXAdZeEI
ZTnuFfg3GDFKZgHtDHapuNDGTMDRi9TYKuaYneSSiKam4ZNRjwhBbp+OQa/q0PjDFWrZr6+ZqtmJ
Um4Jqbff0hLE73Cg0oRvyovEkpPTxy7NwaGSu/SobeXX4spG0NOIhwdpxO5Yay/J7f2rs9AXmYxJ
lU2wC0LPyv0BjO5i3CCvQIvaGnq8hAETmdPMG4yjA0AI+PDRQ7p/zfF7ahm2hLdeYSV+e4dn2oWh
CX3HhOYzrz6KRFqUxe5qp9lBVN5AQ9nV/UEa8fI+uF+9kTG+lnGmQjfWvjxElrlBAo3D5ABxt0uc
ykv+4eN8HOWOBzcCgjhxhHpPji1BvWOeCaNo2Nnv7cD6JMAWxQ4SIY370JIGBzL2oX/m69BLRv8U
RRUdGPrWQRFcEOml3W3mk5hX2mnjSycipxXmYo4Gkc3jJap1T+NMHB9FDulCuFaUIbMNuBrfvh6B
8wTT5MTgmefQJKPqbEyxI5CWxDdfwSltd9VTl+tVMW/Za+PRymfZ2/yCNP3ENxphD8FogNNrt3ca
zz727hJ4TcmuZaS/lTmr6zG2R8CWGl4fpsrMzJ6aClyNEmXX/HemhjiCJrShy1XPsTdoYCKhtJJ3
Epn5HRNG1XUafH09zAdQETmmOz+LjqfT7fvIXkUwGfO/hJrSjoP/r8AYnGvtX7MA+lNT43vHXIU9
1Sf/4Kb6s+ycomrvbPwjQCWp2Vd9thaa47E20ZZ/45IBenDLWll3iBhhlaaTVN5A2h5G3wudClrA
UMFVtCzGNMs+7b0B2FcMezwjab8Nn+xheqgClaBuAhtlSthMzDfMxbY3ox6RR+Dc+5q5yj2/aim+
LcsIje6QUQOb2T/qDon8DEsCbhuOoYAL6qToFCg4smhq17Rf/g7S04/adaxcIrljFMxb5zvjZdH1
aWCLggEM2H+Kdm4OZz0kL6aiAGK13njr/XwLf+nkKIhn66+ZrP0jfJmcT3ylMCugAhmdx7dLPIK0
YV31Q7Ea2IQkn/ly1QORSADuRdwjmXKWg9nPGGfN3oooms7MA3LWhRiXVkbSW350HBG1J6Xta7Zz
TyfNujiEhm+wowcT8zw7uBOHLZKAvzKaOp2A+LC8DzZ7SxkWlNiGCb9j4uQjpSkzXNduDlGhUri8
NRqiWqqVYk+3SEcAtwF/qa79k1QIq7RDtrtmWQsxEdDgFQTJADbftz90QJYkTYrZakSXQKrmBQ9t
P1ucf2IxLDsxHGDGS7Pjn1bTYg5F7f3BkTssLETAtLNn8vy6APWWJuaF29CVEsnig4XsQ00QvW4O
v1zAhz3DWX+jW67UDvfPLSAkJ9JyJryqBoKwRVesQAa/GeBp2JWPiYjEPLiiK0R5J2M6D02ptLFD
WWWKmAy6alSDbADcIPuIFSxAKJ+3yZSPNnhncb1rGrJJu/tOdHOn++PmOV9eoS/ZHrwU4/n1+C5X
037SsffYsO1UjgRzpUiSFdwtb0WUTi4kzcV5AbXhAEt2ynTseSHHTxu87Zz5D9UtivvgMq5w3/1E
pDvfvGeU/WNkbnYFDN5c54YCrgGBNlF8i575UU4NWdeUhieQ6Kxfpv3TC9rlo9Q3d8lFUoencDcP
x96NZzPfSngd2+hoHSOW5C72vWfT5WDX5n2wjOIlc9yt5Ob9sPJgnRp1+1aMTPnlHxFyFKdh/raq
qEFrWK5xz1w2uEDjfIHC56sSSWLqMnBZgGqu2RmOnvarnBs7bHHAxlaO6S1O3viL2xRw1acM3N0T
KxsfcBzzF/jA0nwu3pPmm66niWG/A69uD5/V3vI925eL+dRHEt3BzSCVXTjoVfmji3nWt7weUQY/
qiXrGwMy25DY2GN3r+0Q+vksDTJiiuNQcY7AyCIIx2hzKCj7dsmTQWSypJBIoa8KK/OAbcgsnuUR
l4jNf69zg366W5u+sEI9bnucF2tk5OcJId/DY78AZxhiEgRgyfj7THXa1J5jMUIpIZteBrYHN9N8
s44l+WQQei1PyIl6EoQ4ZD4PGTPaPTv54cfBteqQ6PM5akGC6DhTHjRltf1i/d5b6FCj9yVmwG/g
yHpvmbFSm8ISsYnTRXHfUzzYKp3l7ii4NqnB8OxtwkQr74/R4nvOIiEETIJTpA6NxJgj+DanskpS
L0prt0BZsC564qCrKtgi+/TKp1bYd2b1WgiZglp7G8iHc6ZK79P4/9GVKDn+jAKRbofaIje2bnCA
mS6ghpnMZh8gGpLalmEoH6/5qLVCGAKo7+9+1VGFtxkZn2hNoWp6Jwt0J36Ez36JlTMPWYqNkP9e
I33Zg3TlgQwZyou0UKzSTpdnkjicbVZN4w/GI+nghKqrRCfhr6b8j0Texpx7/jieUzTDlshuvhZ6
VG29H0Hvq360HvnrjR75lenLnjhXTDfBwjoovt+ez2CX6FBiNHmyWjWt8kcF37VYv+N864ksk8FB
/CGUHHX2CpspiIyGwnkNwfmmzZIkkOOxlcTx7aQMwK2pKVOJvJlSfEllXDIf7Z8HC6pMJ+tlLnhO
ApNBUK/xAXHdz7BXWgJlRb+NP9ktKEvlOEPUp4kj3NKak0QarqT9BI70iC+G7PAqXZXXwkJtUxWL
LxEkUHtDChU39BQ++Ak/hlOsOFGxM1zgaa/JsG7JeeH8kmyJ9M3giomTleHmyEWlI2OMafK3BzCU
wwjlP4165IXZrg6hRROT4b1Xu9n5nvdhFbi7ttzHuMyiAa5nwuRL4CkvdDmPnKQ6lUlIL03Sw6az
puSm65qkpf/tAEYwgMeNa/eJKF4oQxApq0VFWsuF4x8V5hSs32ko98sJQ96uw1xsBz9o0o6TkrMd
Z1se6f4yaMijlQ96bs4WPRMoy2XNMwkeqJ6nuX0tdTEjTLJu2OTV6pFPIBbzO6Mw4a2py5rqVidt
zpPvJ4Nr5lAunyPl3PoW+1Iw3sxVZY9tJhf7cl8/Hoqt0TL3H1pAlKLytUf3Q2CTUhjKruoJwzzY
VlkOTXR6OUjPUX7+lfkfYMmX1OWm9q3DfTAEBRPyGGKPfoGuklGXCkOUJIUnxsXAv+/LJeALmzj0
rXnoxNDkUzXTaio/jC/Art+r92G8mtX9gfazLXqkxuwRpnOhqD7+0tzFsoUrJqtRtlhqsPssRdyN
LbkFdVSyH/vrslJ2azbu8rUkgt7hu6gPxFsiTl5bZti4OKlXhEdwJqX70ogfkU5UTjSFWRXW5Y1L
rZnLfoRIB8UAsWjCDnhpMH1VFiM/s2RmpGRBbwPwlPUW+hf3XWaeQuIExXr/GJar0w7YGr+t/mP5
j2EQN7ud0JdaUdX3k+5RYJTjR9sdUmKJOANy83BgXgp4rgMXlietaY7f8V+noqgRVII6dQWId2F3
u6hu3SbFZNEtP/wgb0RQD6okKJfbx8UpIkBwJJLsfrGTqM0LBLTdjGlEYrZtdW1trGZZ+Z7BWkak
QQzjMszEpbAgzICog+12DEYssAF3uU8okjlD1M7ntVkErBVFI5TPgzBECJPBwqXIvKK0Ct8x1mfP
OTCcsc62sEWppU28X1JoXgdoY/3ruOpri0e8OIUL/CyQs45o9jWLVdPugdcRlqB/CcLanSS/yH+n
SXwgF8IKz7F2xRql57h4VOX9ddgZbxA3MHr7z3x4cH+lSFiZWjq93srVOvUrusPPX3NfoU3yMNms
GSKaczDHiyhBEWwFUf7Sf5rhQnwvCLBCkUORQ6xzS8iZTBnDPlvkT7QV/0fAkItD5tf4qCUIeT6c
RsSsJNINpoNA2mcfvTnY9F2cP2L2vBaaDZ5YWxBsaawvat72F2XmaeVU1GX2BuPtmS7hmrPoRpao
qEcBWeZP9Qhv5Vq6ClFpy0GiYEJYtf8BJY77IwvYQqY/4ZgCQ3+Z/onhviXn8Z5X0Vp7AqLpRVnD
B1bJf1uVBh3E3ukzyS4alt0oTUOmBnwabpXAKTIfd8JgCXC2iP/7CXuOdxUR0RLCusTT0tZgR6Sm
51PLHC5hU7ilfvzq3U0qY+0dkKiIk+G1B+0t5S3NUkm87eUkn8oc9zEA/ppcYC+uWzbuTEJrz+pd
Ju3Df0KynU+knQnSpXKmtBpAoJOwnv9H+ZqxVEyUeIbFChPUgBvxfEw6d2SCLQoBlGLviIKgv5Rd
QXC/3hf9f6LjPA6Db+mFN2ADXTvCTjkKJA0jeU/7NgVIahd7+G2XjmgkH8QIIUEec0oVaRPbi4nb
iojikLdNCf1MYjnLGBwzqdadBXbpFC2s62kuKaMr7BrIYVAeB/l8lKM61zq+czZSgpuM+tLgPDRB
GiqvQl3fR3LMJdKlpJTmp5V/zJY0FFVl/cjdj8j8qTiVIzQiej1E5dJ7Fk8l80xiUuqL089oA8ax
NrtW77XLXNaVdq9lfyffxFyjQ/Tmq/NmvoNLwu2/Pr2YntEobx56qe3XG8bAE6FgkImRZJ6gF9Fm
lrWNfXkOb4cFBl6tKON4LkCT0o5ki4nXOCqYD6B5DPRHYEb49D5SDo2O4F2SowLL4RxJxA8es8g/
qSP700VWF2QhFsxX4zMx7jQahabyN5vOKFlO9TAJFgtvBSsI1ao4SyMmEg34s8TF+yvVgrxrX9i0
BWYq761hM3yDVV6cYEs00H2mLilRTzlIMw+x951UTDFmkTHVjfLFFVzSeOrRvZicr0Z0DVpyXRdX
I33FSy4DKbrxbLkLs74L/Cd2VvhcR53DHprSKLO+a+CK0Cuu/ko8qWwQyfnG3twduhpm0wwdPnZh
OB4q/rOyzSiqNH0mgq68OLijZ+HlcHY66FDkZSkhaH+P++dTTtJBxHDU7Bxgi6jSQbfO8S6ejXbl
2uA96q5xZs1AF9rtrweVSffKFNJxlrTJ4HaygRP5epFJTdGpmXuWOB6rEVnJgRbsRYTbXroQZP9O
TXHzXgZAwKjFUMIjfStcTUJipPsrdcH0xj7fT8skonkdYUzKth6BBXfmdctDVkbumQ4zZEPiySZ/
yY/4KaG61tlS1kFVgWO4FV0S2Q2t4quL1qUeNU6PXwmLuRHMuPHU34xXxKS0MMlkZpmKx3uodZP/
The4ziLdzsl+MdSp3g0IlGF0XvbDHIYlTAXR+m6Ofw0aDYTklVhIRrFgz6MNd+g+hktcy7QUT14m
faWa5yChhgvPPM6wrdWBcTt7rFB14c4dBTbSnPhjQRBelD3RWOLO8Dn0dIvJjEMtksNT6oEqS1KU
wzaX0GGbA2iS4bJh2ivYpgWdYOFHJxa2034N0Ja0O0Dr5pOvetO45ZlYs/Qwzt79iIJ8k+uPJOZ5
Gkv9ZzECVZIwm9g0dcjZIWvA4DpbSvV2d+deIHHhvlDHvlkCiaAsLz2gI1eg8YcCoKXCmprMFyqq
bgHCbAw3sW5nGUfFjO/IMhPaQlExU1+Rd+LIZsivhPj10dpekT1ncaaDps6ZUWyE2DzO/wPHw2cu
NMli5f/hgHCI4jQir/1m6eDX3Ex1JKieXuEoGL8fZby/IN6ORgs/5Bx28MjcqpdgaGaXxJ8xchK7
POdm05AH1HwSx0HbmHZ+N6j+F08yyFLRuzo3pVPZeBfCY0U/Wq9pNK+CxLG+NZwaNRStX0KORBau
VQOyarFLx4DOJ1++d97Ggi96epcf/5GW5mk4332y96mTrieHzpdvHVXajxcuT37QAaoaBKzaZOgZ
wTpELrou6nEn5m27My2VFCltauz43mdOYqks4wk3GDKc0bSBpSqnslopMc1hMa9OILf/8FYR46u5
4ok435/WJUZJJIyxYG3cgiHy0CUjHi3adRYNecxdGZZE0lI6URFW2lBQ8iKaRHC1ND0UaxdQKzZ8
OAzdJF4Jbqi+vmnhkE4UtZLJ5Vho29HGOj/RPx97OcPmWRIxcE2gfLsmv2Ak+ZFR3/vr+f0QZd4n
oiXJ6ZqwOfdRmdG9JZW/UdA+enr/dehUtgx5c9Ij4Dp121FhQsGOUyjl2aFGwVCl1Pcger+BTCfU
AOQAC3BUfk3OON8p/seURSfZS8szfx1hntSURcWkcHoPGBmIikv2x1vssQlRzEtJZI/p8KzwX4p9
66Cbxni+e7h75C9QWO9x9tOfeQVJG6+w+e1klwQ5vEqm3wwG6cGXNNWLTsOiUXxuQRedjdaeRKNU
jKZHJxjMvYTYAvL+amCCHpqvN4xj5uWUfKqQwEIRZqCY5rHK8+k4xfK3ll3mZidCAL3IHTsKTmmQ
xAh0UZzchGrQp5GZT7iDW8uwWZ74/gNC2o0MfjW4XuiVgZxHckXEf28V162lG7cQOm2/m16NfHmE
8dz8DxFRTr9+8cYjjtUP9yov/bC7cbHn0vzBWe6Ut5PQ25yewKmSUN5BBOEFKNqbIdMhu4CGdV+e
EUx6R85Eyd5fJMBxBVp8bTUVHZ5o5wQ6/WWudkJlOBJZ3lO1W8r8fJ++O/Ul2wy4hjzPWnRaWkB3
stYXgqv6FBPlc1k3qI7YqGUElaGuAyA6r3/Zi/0ikiqp4Vc4ZGZxrm7KUmYB0a6E5w+gebcqlFqa
jYLO5m3Pn8rOjw3w1hbc70z0z0ZAqgk+w5Asx1jDz6YjaFTM+ynBrSyicG8b+awfyhEk8E3StsEf
FShjbxM6D+lZ/zGAEtOKUiGjosXzgSWOpnhEu78H40roynSmw8aAvX4wEnPh6yy85Cdw8oD+st4P
TCYPGyLMErxODhjb8Ua1VbGCN9qIM3c2kxitlQgUOGQrUXsQJuxmrgNr1Vlda63gfCVtBVCO5KwG
Zth9YzkFkr5i0CZiWqmQUf7mj8gF5FAiciOGR3uXBsNM3LmY8I0qv8Ef+CHjAzKVxj64h3tZzbfU
FAJDT3GhDBhHmc8IKvmH/uVfDy9IVYk2RvoWWyi+w3g8OLnr23UwbegA+Y8Hm51EXNUIyRuetpo6
rJBaIEUZwLsng9W/6uu3JNLHk/e9fdHD3/qR+u3XxMsgr6eHhwinYDOavpfcyQH13oq6XVLBWVq4
jtKCmgTUjwSWL5Jll9pD6DKh2MN475wP9AZbgaYHFfVFbC6dsjDs85jNWTNZTeYF9BQZARE9EaR+
bU5K/P8OjaQHPLhfJO53ejagOx4vp4DZsC8FI53S04XCIvMMPut2GhgfVX6Z+saXwQ9z3NMbKj01
rZ8XkUD4YcRtIY1rwR478SkWsfL4k2qKyhqZ8y6dJK/r2T8v2H+af4tX5MuKaQDjEehNO/oMeg09
xMAtX4KI9z9/0QDTZ6HIIIXom7TfA5GgNZXFVFcMXyoEDs7rTIl6Afn4TwgTXEUNZHVafQRUSnJO
fvwh0wb6iodD3AdfykUvKX2gbXfDE4SSuww0vcoiRAPQR79D9y1zEw+gHK9vsUS/876C/k3SPNZE
hZWk3cDVDOMyOYR7NCG2H+qf5atSgIPGhvs2rYJ/WzzyhPJLXz4NG54N8Heb9etOoTka9alKHN7o
vBgM+NMJyVkgCSGXui7nd4CAssNobRDLVeYiUdNxLGLMkP9G0wURcqYdITe+U+3dziWPa0+OzMxp
sod69Wa+BSXayGupvhcSya7zbEuYT/Rk50t64dBDuDbNtFsa1DvSDX2TI+H0n8RLVktvIIGF/cvE
yStHoJIYm0Qs53mU74VU+ZrH0PseqqbfpEK/X4ATkcjF2YVhEnn1L9BpA2k33vKXwGz4PZsHX9Jf
vkJdHuWqu7O07dsuHCfvVmhmCY2HQEZAx9/Ehz7ZwgoLkuP0jrPan7zr3h/j1ehXd1RGgVQBZ/IY
C3ssERvNrSqmsJXlguF+iiNpyCI8/IkTuQScd804Dn6x0jq/9/Ph3GEhZf8HkjLRsPS+Uh8Ci2V1
gF8hl8lRFRxME2Gn0jRHoZRepEAWAYmc8i0A1yFuu0w6lMzUh8UbsULTAF/ZJEMkPCi+a0UboC44
xrDocEGquAN4P1WD7oM7LQdeMFYleS7g6C8+7Wox7SngfLDeLX0ro7x/aOUxYutltagy7oA/zUnu
QPJe5rlw78zV15IgiuJQbVOqFZXb+TNxHXTNmBp4/WuwRISdYuxqlhbMVFPYQO8iIUXXZJAFR/Eo
kfEIj7BGNqe4MGRDHRrLy4N1L2QOIQh8+SkzN72Jisxaz7GBVtSekbYB4878G6zrTMHfZaiLZBKb
bZdo2JjXVSZNpqelnhT1q9YWI/GCofY6GDiW3OxS1Hdcssco8LGcbS99zZyE1MkGu0hhsY5DPtl6
xs/K8K1uyL9C0QQYH6XM+ORKIBOeu3lfaFM5EIHxTwOSjAyHERIG4mwAUORwgGqb9fbMCMRAr/IN
SSH4ojri2+YYGnvcrxxzL9RPy32jfE7B+UGf5knmG9ZBw3o6gXEAqC29m3k4v8bYS/uK8d/Siur4
HkNh8IDujmXp8lmbW7SZXsY5zbblqW3nVlmt9T0a48+ityAZpJP0Hf4IQM+hiidziQKagCDcNhbG
3urHc4Aew3IlZJeQYg2jCP2jZreZzGSlG56QKtcnzvS7BTxZ4lmrLhxDk2sAiKKMo9eIiWQQGSAM
f5Xx/w7g9AQBSYpWhKC84fGdb+73xyMlqe1ZnYXwTSvi7nKN42C3+PEK7DOrsLPP+fRScX+ODVNl
0U6ZZE1mqytIz5m2Gt45j9KI64erqj/HHGiyLyz6RyZZu3iPRlxKYdSa3TpoEsevpDF9p147px5w
55smsvVCAU2NJgnkEV9hms92p2UcDRKWJP7TmpgRYsW9Ih2L8BN+y8XZR3+UQfV4eGmWruCWTuXR
NRhbiJd1WqIthawKeeO6Svh1Zdo5Bo6GnAzGP5WEYLI5wjD+7CZtwpqReu1iQ7Qubo57F/6eZ84f
06qc49xsOgN+G20i7CWdFWw+uJFBuwGhxsZouSmt+E0aBSH4O1yxTwI4tyM7TUTmfD/HZxHqc0Ew
4fYAwzL+c6go/RtXTJPuIdcIQcOF9qwohRSWjLb/FVfVHDdBend5VE0wUAneOhp+WXlTkQjEcq1n
NeoyV6bBeICsw97+uhdV2gTWTAKZHCn5GFgVQ246+w1whzqbdTjzL2VKr/a9zkKQd137MI14H2+2
uG7St/RbCQqBfe/rAK1BpBo1bfJV1ZgFoQtrXWwYZt81lBYGruW5xSEajmatOHX24NJXdCcO7ubS
arRpSQWyQeMR759cH2YAhDxyXsrTIZ8YUEbF2QuBOeDSm6t1M6iJkljYNuGcDchf8XZa++mGiGC9
9ojX0IZzhoi1Vw9ICLpsRUXgKjqz4VYNGNr0Iudjzi5gfpZcEI+6tlSi/d3DM66LwPCtfVhB51D6
a/qOJmMl2AD6PGDoDDYwvu0RRomZalUW6BgOD/zFBD+oMv9LYaDT6ZI1V+JgE5zFH9K1ddT49tuf
vVtfzKHQeZ2Xy0+3i6Q+XqygWpHFIMa/Lu+CLFa8FnDA//ANxgd1aKberLGL9DyU35A/uodH3V8x
ryrjXChO4cr+7cSBJanrG3PzTsHQvpZSIqmhsC3bNhYASnNoUN4I3aMHM0WTJvoItBuYN5svi59o
2cKnaelWOwFUE7RI0TjX9AHLRjrsnjS5PqFsrH0WXyQbDQB0XiaWk4e6FKiekPLN7V23zglBAQrx
8OGwgf5OrkRlJr15E/IAdzaakQLT7GKIE6VOLDj5ajd0a7dFLQ90e6/XmID3Z+lSNF2FV7zD8RtH
PIfrxAFhmBjXSfYDu4urvTlP9n6Pkrey1CZeJQdet899/NRpz5Rt1gcqRwHiuum6qzXkSAY/kADq
RQSf0uym0CwZKOk5256tYJO+lcSzMYq+0VUVtwVPwNRlQUlP3D8es06fOBDxzfPlcXIQ/CST5Rfa
5Ex48Ta0tgP2ABd6wYccuY+H2BOxMQEfpWAkfMbaTxkmXOkhTIXZbBoksFvIDeyu8NEAj5qZKnbT
HHROr5q8ongYTPyH8bZhP/p8z5jJ7zEnc7s798EEFMN/hb9whzX3YUrCOTYsyKRJnPF8LrDePcw5
B0zBfSMiIGjApP3I/0kYl7tkgy2RWfuIuLpJHC8WGfa0ShxIEs45iXHAdi/Chu2VxQ0YeILXQjkY
VSUUzFvaKVCtGSKot9VmsYm4SyLm/cCccA76csIhslsWdGZzuBmo+ATRYfZmuW/1cYPFLEnIuwHw
XP4Cwi7bXxggUuT+bxBEaz2hcfPQSX6+Dz+Xxg9xiw3zmdmqFTjiQ80lU0xYXv4gpj0xqJE3W/Tv
pja4ZF/FXgE+/pNpUmG4G8FepeTsUUFZOfREJ67uPwUr79LT2I8QZ5ehJKtQjDk6VE+AglG95qIm
2lMcRt+XHauWD9uBq19DmNjGtvU0QxO8LoHwDNjsDh08ZThKjH5xqGtNYMM/9o0R8nHJPc9XW1EL
6LLNqtmBOTT1GMegO8Dx7B1udbtsDwYg42nA46oBboqn+GpVyRkSPdkrA/WORkg5XGMzH7Qz62YW
yrjldaKo0ThLAh6q928xVu7fEn0QQeuU/C35v8CpQYcqAXbCnRGxUsFHkAHh390+SWTpBja8eTIM
I96LBqOuX1zJdT/PMurvx0H8CYPG6ReBwjsfGU0c7WS1Ap96y0soGI0UKV0zvh8fC32eJcHBfOYs
RaAMZ91HKslQC0WQwaYFA+GWpIto8hR/43KaG9xL8pvQa6lOZVBqMF6aEXa6ZBm7+NlVgMs52mRB
YrubGqXUC+3JSASC6I5GGOrQ7L/2FItt4HMCjDURXA0FXKGrfWclZt0nFOga7KPiiuaPZMnKt9Fn
M97G8oP/QWkhoJyzL/eMTi0y9Sc/k2aebhP9/2nMAzOQ2pO+O9gwUvpoUpfwlN7IqPmYM4ivkwNb
jiJ0kdbdXsOj/mXYvvRIVR94DH/I+4RCTNVtpSOu033fquVyHYkrUfzGMtE5EMzliwbUu9AuCuPj
3k3IT6XsbFVxHhhvfwmcUdNKZ7Mto7Ln47uABlqQstBoUMiSDfifOrbJp8LZDOwLbk0PwawT72O9
jaV9ka09Hy3mqvXBuMdiQ7urkneLiIHGa7dcMw//l1jtBn+J0lEJ583d00ZMHc9ZLyj1v/Lh5XbO
V5vMCxGKiLC/19Be4tnlLalVMjCFwTxnVQJcrWSuubhk9/OfvMVs0mz7hJSUixD1BnlyRhM2U3XV
U4P6RRoNf4kzM2M3f6URkx6q2q/F9tBCHtZ+t2abxhAIESfaOxq4ov/Da0+tOGBfIeq5iE1bS1Zc
LdmTY6J3KcgsBkYIDRGv7co9fNYJk/HAbbqlrmRFWqG0QVDesdvDNXR81ZpRNoSP1AoTAivbeUcA
UC5K/EBvZ3X9hWJkimIuxB8YoVFsajnCc0PdzAt+egLvLAX9iHFyN+b7RgEKoRLY9G6vGjLyQ9y2
hgKLbeLOhqNramAFjKWbcbjXDSESjT0UXd4scIRSvgO08bF63qnwBhBw7wUmAhORolByv7FQmq1W
AbVjnVttSlwlsOINgKXKfY5rKym75xaitMs6VHZ2e5Uk5UFsJcPrC6HCqmKaUOvsO7CYxbov4rFn
tgsn6NS8h9+RgQBV1rVpPEnd0f4QFCrHHsSX3E0Ly4RSpCHaOrCvL5HM3x8ymhcBhLIvC7MIg5i7
M7kvaTAxOjXw1WSQA/WM1677kWw6fAmA57OHh5Qje5RTSXhEwq430R1QZiqhD+fEi98wAfT4buHH
Jtb7OHaewZJRIOHDRxEPDi3rbn1afwlPpKOWgtqpaemzTbzAREnctP0AOskPIfrw+fhwtybux/OT
ELUH6a7ZhkEn0KoB8pPbnAAwmaNNcplcGeocxu3p2YVu4/ZtAsLg4/wHqAoRKfsHuYqeUAE6cwnY
jQN+RbzEV99WpEezzDmvF+9MY0Zw39qaSg9iwHCpEMHa+pGLu8bztfesEAkN2KDspyEVgoVN3ygV
r3GcBBb7glIM9vDpXCas1/695KIhOWAyC4CLhs963fYLny+iOuG2ROXzsUmNh24RpFAvyzpk+oTz
MzBWBmdula0XZn1qag7lZhHzlZmrdHPejZxsKiw6agVccH5WWzlIZTLfOXAtmH9JVYEt5b+56uyQ
6hy8wvYisutH+848mr77J5oBv+gpIg0COmfEeqoFnkrgF4aWkiEh+Fb2BWPfCgbEVNLMPq3uxWzC
WnuTT7d+T6pgaR7UOBP8afAbvGO8zLBz2luZ49y4CW9Zu4qcXDhvSi+XZsheGA3WnhIUZJD4gD8d
16rhKtxQVyDRbOm6uAbHXGj01y+voHJYE0AAW1ClYLMYIs5lFYFcuik9TZ8LRsCiBuLfK0Ehuel3
gOuf939xz8GZn/obAG/WtPYJGYGVxQsVBNvv724qsU4gLe5SQws2G1YSO0A452S4nnuQMZZbxjwC
LzTRh/NTtQGgauJNrdo0wCWashyAXUV8VAJRJHbt8W76uzS3553NQO5vK6qqffn4TYj2Ew01YwoY
mnbLtxeJKZ33e4zJgOXsCHrmsf7Jq+W3hohWYxmsK5py7IDaFP8+AtTk8v5cGPHGNkaqj0QJAIu6
0R5U/5lRb72rF7CttHd7UzhB6eMQLCWjrrj3ahHZrDVDmL5fvdgQzcijvf3Tx0PtaNX2a5jhhiIn
OGU/Ja72GMwHS5UERDEgVGhi/4ZycpFunfcmWANjhIQPqXeMgQVHs87luJ1zu24TFOF5tOU3kOac
YgvrLqL3RGUZXGYT5Etwfq9KQja5/STf3DGJkA9xwz0w7Lp8Y+WhEYzLM2+eqsPye30XpaHxxDWg
xYqxVr8hZLe6AnCa//oQG5gCSHzFcCgGX19u8DzYxPX66UcTYcf5X+kXXbgbBdiiekDGJNs10UOl
DiXbK/TM4DSBCKpi3wVfEMr72W3htYdo6vgtwWRROukMnb6S4ginq8qi/iqmZTYCfoEWv3JgROpz
o4YBmwHKpOX4DCdGqIHMcW7LGdZOO41xBMN67k/QRDoOGTFwSsHwRqJQSrOhA5pznkbNak4Io4tL
afjNKiKcR4yZ7p4J18b3fxNtays1Fdc4V4//l6MdpPVQBwV738AAJcOTdjz3XZNyBvjyRSpAkqCy
KP34IREtW9ve+VlWh4jgGbeXGyrvRbZkYWAGKoidkr0CSKYkUupP7I9EedQDVat7Uw9G8rp2pXZh
HbqiUK/b5yU20nTWUlLjPe+RiKm7uHgPJcrWvBDaSpWz+i3KaoDrqMguESL61+5rScJJvlg7dxje
BAyIF24X0VFyxVPNATRekKxuGJLkaBajiiMxK0SfvZGh8tUgZxfLoQ9DSzRhX47RG0w9qF7VTe6j
gdRW8elMLh56GabwxcmMRu+UuXSqieShRl11N142Wo1em2LsHANQE+6LyFUjoem+koU/ouYICrEd
tEzpvdZgok9SnOUfFmNCCzOltiwt5L9en10ykdMeJ4yZu4YN8GbSLfajNEUZNfFv/Jyie1hsz+CN
dE8d8AyTNZiTzN0EUS8ziHC+hp426+L0JSQZ6WEJBPUIHfyEyES1NoPTvP6ZqciMjroMh5G/cw2/
gC8nu0wvY3Ee+Q2qW8T+UEd99Ag8zDHqnLKe1MA3AejjxFmdjondGc9MlxnCZ1a3cNl4YcZA9Cho
9Xe3lQH7ByvaD/lBO8ZXIO1LdHc8t0WAj2CSQU5eJgTPAZ3bGYWgeaeFpf5ogT2Itin0GNCUx5zT
8Yp8gHeFfOOQbh2gItoQ2YE2FSk/pbKDUS/t66DptMwVJFJ1C4Mm0D7OywLg04LFDJaZLnY8TY7/
tDD1DcUfjIVzwpDNt05Nurgerzcxg8A3+cUFRA/L5ormVVngMmf0FXMPS9PA8H1dNPBkoBy0Qr29
MavH7FGwZt2mrRzElE80ZsUSra6vVO9fZJTXxFKACQUv038mxltTc8ODveSRsLB6mpsBC3yO2bvx
D2dNZQYgq6ZrotpVtHwbyTtc60IgGmcG1QGJttSTnY2QigWVLljtktgtQ8yxxGAlEfqKqMghQdwu
cY6qDTpT1iHPlbt5Kr+Wsyh5weWF9N8exPswYfVrxQTHUdCEnR0zYyCsgvR2+kyk8c9U0XlY1L6y
/5LXaBmOQr1XIJykHjjIOljUpewTvOS7jgEIOrzPUFlxYa74IuTn3BbAKlKWwNlYMkCyQ4YBGA/n
GrCa1CA50Th3hXN76IaV+XoIgavUXoUUaXdeHNt7HXgcj9zMNtwGOnYHPRubJg5RXIJx7alR8EtH
D8U1nDA0jWcrYRSzaoRjHfGsVe3NuVGwoGvce3tlx6naw9Hg/8tFJHPo/r1I798WtkJns8Sa1sCi
O/eQihvjQAbMvBMDqW+hbf0hwliLt2+9FL/w0irX0+wmaMQrKiYVs9J08pQkhsfUhZNKfjR+OEoH
KOmpOKYCV25JAUljtpVBSR68Oui7Gxn6knNZFY5rmJPLDJy6LtpfiZ/oQMfResgmW6cZx8pfuWX5
wWgH9GiF55Vb8XYHbKBNVqE7DjZEdfhLwn+HeuxBHiq6pjItnbpuCgT3ejj5x7eexTH64OqW9tjt
A2zljDNtW3cF3DwuFiSy9NRqvRCeFsNUKQloZaCOle5CbHvPcucYBJ+WXSqS4chBTDru+SPqhP9F
GQBXcmOd6ice0iYws2HwN4okTVUy4CpZp/5GVh5KbOqty/nz9Yzxmlf6UTBYIFpr9uhoBkVgdFkR
4EWCTf25VNCl2Od7jxDlDXq6h1dh3aBcb1P4SWlTYS3yO7luII05Gbih0mNH+8byV5GM7yUxF5AR
mYGQbsL4h9djCM7pAr+J6yWc9obaIFAzladm2ZMAIGitc5ZwmRMnTyocMwvqYSHYgAhUwiZLXcMQ
VwRxiNS1VMKy3epo4YXMCsFOtskOVT175ol8e+vtnWUZ0uw7eX/B/ni+HH2N2b17OtxxdKRESiYE
7fS+bMS2FcTdTBlHPBXptmZiXpceAeHzAW+0U6vgB/breYDBJ9pf7GKVUV8XDYptK2FkMRfuGOXH
99eYmFnpcuM/omPTH2CVGOvOq9+hedk7w7WI5oBTJCqdNuUo87QhqbZ9VjvvG8BPQA/Cj9MMcpL7
aqrMnJQ3LEJy08uLqGZwKvnZPUGp3bkIUTxnaJ6PfeKkNh0Dy5Xw7dku6/mBLXyp9q0zznVISXj0
vRP7+mas2GOzXgmQeaLoz6HYSW2VplnSs6PiKlfTMQdlc+UOYfbSW6FrQ+fdsSItKpMwLGq42b1P
/6rRBnq+HgLmuBP04epGas3YG49BSXU4AWMYcXQhhHmT10re54pbBlGDhp8OL4JPHJQ6CIGA5qhL
9yljJTjJtgB10+AM0LjYFqt559ez9GoIzMuVeM1+eI2FiYrOus86RFnrHQqto2Hq9V1WX2LrJYAj
aI2sDr943h6WN0JqtTLW0gbj5w94FoXhivAarwNJ+WFBxl7FsJpHmdGbNOcsTczWNo+Qx0kNKZ4f
tql83/kJ/sHszq3NquPeK3ADKYNZjCUtWJXflo7TbwXnhTQnuJOAhY8Qc2BtK0YVLB4+kDaMrSA+
NtY4EZyMYEm0EdUyzzxnenQJ/v1Q4ke/3h/g5wCpWEfCMO3lVCBYus9YA3BNp4CEnP5OUDpxkAAj
4udyVkA2Bg0aS5Gt2aJg1JDPsBxvnzI8ZRPE8o4KlMYjMIIOUfn7n4SkwDJiEEx82agHzXAQQ/Lt
StFKVrBGajhKVCyO/SojDsbGXeiigNbyYiS9HliJrosyIjg1ooq3KLpVc6Lgqu+CWhxPO+SBZeiM
ecRCY7fS/eadMnApp2ZOyWD3jeOtjXkOCnu4P/VBewPfkAchxLmofN6wEgsrtzuNt6nlw5an7ITs
27K0EzxL/7E3cxFEMRKaZlVBgUqvSrISMh7QCewC0G4iy9g2VlXPcQJEtFjaMxJw/Mpa3px771jz
IPNwu7zrMP2DdjArfAV+AAfNwoXqCwYlIndo6fqwyOSbJGCw4SoHlgo4YUuXcB6b9xpr5zxi+9gU
z6/a44ThNNyjZbBj+btbSYH4sutBgPLnzGq0ZADWWLFx79kau6ZJY8dn+ZR/0SuU+9npN/HPZy1M
8A6JYiEA9STO0jz2e6zzEU+wgzQWp1FLGNHdmBbRNNUH+QKaP49LrU7VWVeX8cic2SclH+URD0dD
wGQMu/f3HfN5mbygG9+XaxNqAwtfMxV2vOBgnK5BO/RBAWCBXKhYyo1m/C5yFzkMQskkj4krA/uw
hkAE3UWYiMkbwTe/6GcFMgnOsuk3jGQChggcQuhXLq8x18UlM7X9/dPVwB7MHTtjCvzfn9F4Lj4K
bA0zaYe+fH8Bmq1szHkbw9VYkx46rF0I6VGtwbzbIedgaLZN1lLL6qa8oAWSEYtO7SDMxYG4Nk/q
HFwtXP3OWBnT/7wK+RSDxlClvLBh8ZQWsZnjleFABUSk6ear73oECQuKMkqz6cIK1wjKd7f93zlr
digc0rtbrdZYdck9KLu7MJ3k9x1DVvCy3pfegT9J0LvepooOjZHYGcw92tDExqoWbSWoVzT1r9my
6zFaUG1nwrofe4avJ9BHZqeRdhcISc9feXa4J3246RKX9pVWa/am+aDMSE9X4TyarktKJ/toPr5V
v93PYGVQqmPyZx31isyS5u6/usZPdNgKQ6KP7zLYotq80b0gPIL5QV2kSWEKPSRGZq2qS0ismL2F
Cww7fd5qBL/XrBRSmyAfV733QuS28lk6uBoVT4gszjI/NUfb4WvU5PrUxf5kiHbsWm3km37yG50J
rreeoNJmb3NBeuWgzklAzDYORdiVzP+5bDZt/XaC72PUhTKUxDpIx70Oan9H2Ia7p99rtqTQ7dpc
X1OgPw3ZvhXjPZw4ryxXYO7LFVAGD+f3XaXSmbTw/DgMrro3tzg4NsWWREwvArHnjCLA3lHFfwVA
WO7cQL/myO7cjmA1k+IS1bc6n9Mi9cVb6K1SwbtH/soBRMPAsNAlUth2WFuSg6Ksu6uFavv8u7Ar
5YKeTRCjy6r/FFVbYim+mde8K1ZkHMlJD86pzG2zKpOvud6Xp6iP7cgQwB52ElXH9DirTnXXlVYv
CVXtDb1XcC6LCUecDNDA4FgVN4FiXykX4fovQZ2h1aQkMGCUgS6Ss2R1rLKbq2g1uXwZUZrLwrI8
Kfqkb6VJS3T+sh6YorY1j9izi7mjfgwbcA5A1lAB+45jqNAW5egDquNTPQwOurNqxbAYJydWcjVb
fPod7W8fJzR0cqBtwSZWS7aYWdYdgX1cmsLmP0aF9zPSVi6fj5ZzJ1Cb3k2RogqkCE2kiKE6SO8/
6yL4X37TJTET2uU25ZHOJzVZfqz2wBf7KOM7q18NSX3TitXw0yJDX/3G3CGqtFY2FqVEoMKYx+Sg
Kf1v9xYLBUMGoyfCBDzzilQO39abpTbTKtFH6x9s2HC3Yvs+xw/1xmHmcBhSthX8+iXpKvLLPjvT
5QEsWt9rbYk6zC1sX9o2hz7fn4mvGBIdWqkO95DGJnTf+Wcx5ayPkK0HHQAHxmHKdViV8AuIFsGY
idaqxAuRui+QwIAWbafm2KpgUPNSsa+p0qUaBP5O5DZeF3MK60B9xHEb3XcMILmwbWSRLi8+/Fhv
fo4X/t/ci60Nf62ewaGjva9LMMKDfMLOGnzXfrsfYsOZOeagzjLtw3Tra2TlCG6t9PDMVsxEl1DP
3soOq51T15Oue+HP/wQAeZoZOLzKHRQpZaJC7+M2ojyZMEH5TXoNiTX+JsU0NjQY7FqgAMT5rLzr
MHqt42zDFNmLUul9PYX9RYNSXgkxRtO7I5+YbUAIV0eI6HXNDkt1CUpCaKmztPnCxib4tLCE+ckd
f/bIzcJVgOZUXMcqFSjFCZcsBWjc5zgUhOKbxDGZAWleMrzRnHbI8++FWngDGDDkyrg1G1125utu
4MkHJriIN25xiPqlE82nEjjcGzYCbb5Q+4JaNRdOaSIsyj33Z2RK9wOKFbHarZtTvdeivOynpb1F
pXqpKIKDxvVrF+P/TBlEBydV5oOqEd7rYVFCwljcS1FcaH+71/ucVrJkfhMESUc/03jBmaVAxH3S
2OeEzyfkl1boeZuOT7cXeIHm1IGGG3+DF3pxZybIPoedgvsW6dc7UhPBYSJMWMRVep6f6cxhzBir
XIOVxrYNw8HDhWH5IzSMzFxi7w26M3ECD0LdtfAk65BYJifD8UDw5N4ysDVWleOUwqi1QlTHc+az
tUBvwDeMfbqCz6U3azV5bLt3g/Tiht2C6TFwZgoYN8+1AOOvE8Onk8wuY3nJxC9/avqmrsCOiNhA
zWon4e030dFh+/BSxt77ZtvFljuztMOmI1kpJYQcTS53rYOLqn77Yi5gbce0RdgsNsdiuhenf9A8
0c85aEyzofDDcTmkWdqkkLGfDjGSuBpWuRG+edBQEL61AlxVSLaZGvWy4MZvwbzEMduFgSZulhZC
j8FbVP0IjvkmbNgKcB+rZX7N4/R4LpNh9SBeeB48MFfDCvAYDx9By04SeKgZDjov/OGScNKaFKvc
s5kmCxZJNrgh92JbwK+AMjb1sayQO+4nSuIjxgWJnAvoo2br1UigTF2JKuFAwyCR0R48Z7L/Lyw4
+Sh2bR+A5YKrI7tp/AFBn8BwMNq8+9Fogem6SUQMtHPsfM0FvnyucVZKDRdhAGsPcQSfy5kL4EMi
K3F4cpc7o6HgEMHGT79GMvs1gh553sQ3bDsOpzIiOU1DcUe9UypJob/uo0BkctiJwQFflmZZs25j
Fo31U9P/E8ISfVzz1AYQLTP2Yd3veeoSlGld1+u6IXxndE4PrxTARYER4hgnH3j50XA802r/tMIS
MGg6szgLedxYBdKyYwWjx5hEfe9rA8+QZCQplHeHPqPylP5o/wf/YdY1rHFFynyJbXuw5qut6UrC
qSUTJVJie6lMkbeMl2tGac/M/Jd+k4Tk3Cis4dN7rGN8/HxZxdt90YqvGuG/UeXDjUHZSbclDHNM
EYEpAK3xesxGCU992AAUMAws9v29MfhifA7FiRkOQMvsyipQ+HifXAH60UFkBUC6FPpu0cTpFIEv
3haNCPz1q4H+LKn6OWUy9+upeV9aW3FxcYwXZCTvBDjYT5fV9Q1tkfWm7LXWCNq7DKWPNzc1m1uy
11a4Yc6v2UrXLKe1wQ32Kvdj48CBKn65DbI6r3qFLrFvc3Zny/04xi7/fT0dTMVynhcykzUHmpd3
4Y2e2QtTvG3paXvy+vQIWs0b3YJBIo6whZbj70u/QPtFjDxhMNpuHgcu5RafGb5YSfxdXP6CnCpy
Y2vx1NSomPsnY1gFKbDWUgOciavtQ47W35lb6UtQgZRMtckrjvuIvIxIQmtrlgxLPYF0R3drsVvl
30ZuR7DYIXC4rOSqzX4svJ2Tl2rT19ZTEvWdbUf0+X30bvD4+9JM2fCl5B5BJHWp3CiNPIzJK8W2
s2UoaCYAaE0P52LnMgH73wHE637cLRS9ED3J+dvUAJHqXydV5FFBL/0WFPgDFA+nYBbj7LpgIbZy
pQ8AWNgx0LO8NoXnDoID1g9d/+/5gMphdz5BA/8g7L8MNA6JghsMkuiTyYmY00s84NGSRzOoVXfL
0YcgVEf972PisNLWcM7YQamGMftSC/JdFgGpm6v1I5F8XwKJWy4/lLdzDmfF0CwCMNh0nY4CCoSK
nUm4LQAg7Kz7rQITznYpPcKO7LdwLdI6oSFRaPUJ2BRVraJ027k+2rpEhDkEB2OswYK1Gff4+Vcr
UZPAwIfF9ImFwnufJABl/2sO4uJ7tIslaMloV7WHtRe5qf7MxomMIQ8syAR5YBk+CJsqZzF6p5DI
bd1UmVMBHFOZlXtJM0RZHlOQBrcNYOz3RmYHamYPoCWZfvW6xsILxErmLGgG3HXXdQVK08qBE3bd
a6xZwVQrXSakHBzO1vXINR2NGOISJlQCYMD3kO5KHt28gQ07CA9HW8UUv0opZXQVB7K4HsUlkLtH
WH6ftWPxnqzmWJdVAty8LdgZkKz7vpGYsn+5D4beKohzkFZPEvJ7C+/ba7W9NPOVKYkAzxNysK3F
Vy+pBTa44sCjp30X3YVtS0G6E+VuKfAe9b74YYOWvEtNrQ0DNof6OWPwcKqxyokKVL3kMV0WjE3P
bG70RPR8+AhTHZV13aFIyegh8QgWgZKlry2SbK3eYCY2ZYnufJhiS4AtORDOe/BhJXy/hhW2OI/i
rtsp1TXhn5oLcWWIAT0rmXfoWugBBPsJJ0qdQjLDBAkR1fGS97rboqx0lpLxTIVh5CXQ+iML7VYp
yco2Zg20ZLXR/sdfMXvf5yYZfwxJTX08wRD7ujdSxa7TPTnyUAylnroP5wXJ6rM6kEQ6ubJzfYZm
3Z2zJHjdzsqp6/Yk1HeVI9of4YyLh1rQY+SryzhDHjMDx3nSh0+85EMGOXeE8sr0vgskqnFqELOs
wAbcgmYJ+1O7wAv2GQlTiPFVVOvDZYgpNPf93e9DXBng7u6HgDntHP89jtxCJL5LcAaqeu9t9S+t
bHMi0QBo5qGs7luweEEfRbUr5FqSQ5fGqdwW9REhF+H+dYW7CMSb84FpYYC0pdhXUVLyp6YReDji
6DT64mk1rTmB32gVf0HGbuFZyYixlXH1/6ZudUJN2oU0ZgFv120hhtTustdf9zup9kxpjnf6TLCX
mL4wWlPsLZgoCPaJ02trunlh3A4T19ghmRh+R+EGKLFSY6D8yayVm6FpHECqIJSOWxSneul1jQ5z
WDbEfzWjpgo7UlLqNzPl2GzEUEBz07PM9GvtmPycfUaJE9kZmVFwX7WrQKoJY5WrFi0+rL9DjLrR
Eoiae/+dqX1Sl7AZgDgZT8VTbSoljQ72BJ20+W8Qq3XlyDF0ko8ekw54RZ7QlvP+j03F0xso8Bmj
m7HASe8RRcfUBpevjZaY/LrN05aIsbNQgeYIaJFIkgqYJmNJW+il7tYpedtNYiiC3fuZNYG+/t3v
/HupP4zpaGhbYh87qFVcN8JLprSma0bPumhF0uD5jw3HZfDtpWZoV/ZXoc36rCovf5jcdhL/HY9A
KvyVUe5pvnxdC6bN06MR6YQomiQJH3z3jNfiPzEl5qxPb+wVj9MpqUOc88koBz/DP4zgvc5yXiWS
5uNHW2+M5ahOF/QgvC0Ua+GzK1NVaTFf95lismj/2s26XHm0mldrQ6KznhL4caMnQWB5G7Fnn4Vm
CLtkBZqMJLTWITIFIjqp2ikbZ8sFDaN/F8j7brSdBdU+uQCNvMSjr+kBDlAkMMe+m5v1bpKodUJZ
H8ZK2l/DGz/9tJp5AXTLTL89sB/xhRZPhwnocQZW+n0d7rDSjWz4F4zml2koHRMnq3QebRqSCW69
oMUXo80XkBIxxFU28xmcTXe/ufrDBYY9hUpOJSVFk+O5OosdxZnsU2oZ6cZQsQ31J8M7jtMnVhYC
WxHqQ5BCi2rY6U92vyVPWkTFCrPcYtqv3V5ESUEs1VTeH67OS9tsT7Csh5761byA6bG3O8k4jjA5
0w3i1LKD/dcxNfmRsY82QX/Ko3/A2Bup80KFcyf9Fh1wuRl38Z+mmZzcTyJPjSfFQmZNYFt8bbcD
yn6we6YsvrSpNsTQD+blrZaw8qdVhjjL7u8eIjNNg40TnAb9k1rltbPzI+kdZsVx2zT+cVFM5dRE
jk6H+qMi8CddL9yQG1hjT41SSr7P1FjIv30QIpWLDdnm9Q9SDt/B0DtoN1bcHmg9gEKFIe5f9J57
kSyiKvckZLBylb+ccbxIwuPzC1Y9q7VpaapVKZKqZecvUCeJ9eBdyZW3H3+EMbFDOGVY0cPkdKFY
z7VHkZC1r6PbuPofF8x3XVKInaPEECG6ui1rc9MPDKNzSWhuPzi1/7mikwsZO9bkeR/YECs4t7SR
ZuT1JRBOr7NCW2M/gwrfBcL8qc/H8ibSK0D1yYJydjcjb8s/D1XyUH+Q+RGpj1Yw+/uZ1+9oTYCl
8Xfj3jBCUS1ZHLfwZwGlEHQoZzriVXrgYZNdhegjNXP73TKRLFdWAcl9PBbiGj3fBYq0vUrPizyi
pB/CgNFeJSFMB6wOlYbgXkwRUBSCwB69dxsiKAwn1RcsQq7AIkqTItoMUXFjbTXNxc00y+lRr8DA
eMqCvuh+d1JVuwpdwfy/kaK0meaAJhZI0Y79svbKguwmHuFdk1C84/3g634+0QrqffryUOWSJ4Yz
1L+quLhe/VauhXuV+1O8FDiJoa4Hv3oRXzeUk51y7bL20ZSAosfcea9tPpmvZJ2rLDqpfi2wxxrf
gUn9n2t+ZdDkVEe/WmAZtGj47BcZxvwK6bihgB3vnBSCF6Zfr5jLUbUFjg23Pwo5uviA3OAOkYWe
rSDsrQZF4lsuzZNXXQ6AwNscttFdQ1+Mm0PzDkyOb0HtkI5pyEjeJc53Nqo+KSX+HVS3BudWTfLc
jZv3V6BW+tKbeNL3lja/qlkKAJzCkOqAqleeuSNdorkf9fWB80wkkpxELzIuJvRzfUdxdO5MSkY1
/ZBnjrZlbJcrGrmND7bS6Bj8Rt5tS5thv3EnCbsFXlcWBCv7yTSrlS9//P7VoaimOue+0Lr907dl
VLQ1cJsoGMKTyNpaRpMSIF3B/hrJvPBUrIe17T3sHIrPjbqfOyHWFhB7ZDxAIYhT0oli9INujap/
fjGLyRFPXEny3swZnpXVL/fdYWtqqPGQIe4O124iGqLjOnSIeWgsCCxKHGvf/rXDD2gpHgvyA2m+
TgGhIGfgVNGS6frTdzhSVXvFzS0t6aTgMzQw4uuJZbsnRCkJsMfG1xWzaU7cr+uPkoVHU7ny5ooe
DJj+3Rmg/GtgsU2YGPQjeX1HvLOsWlaRDEwCk91opwVgpBzvYT7QHPSFOdzNCpYcqenEnDuo0dhc
EeWfiA9R0mNoBKil1W0vwOSaGNltSJViNE/Zz8HfmrWiJGgEd3Tcxkls5aUrxOLcMqmugGi88yvc
13UK6020bKC5V2HFzGWGMDko+yBllkixLATuoyvMZfXo83KUCwx4hKH+12OK2ZQWIfiQih1zjzvB
Hu92SIRU4j/jFmvgYFAO/+vAPJXLIjzy7s1mdr8rPyIGew5gDIcRWXUGPKvTipZ2D4a9pOuj82Mr
X9yULroYbV+Um40tWFai4NWbGWB5fIYVxoGo6bcswDy1hT7gDPSHLIFhlta6ZTkt3JyB8xd483Vu
WKaezB7+GnTXL8VlXT/lrL8Vf+7wQ+CYB/NY+AQWCx+l/5RIWYw0uXLkN2xlRYL3AmKH/U5aypmQ
tDz5/9MIEYPK2Ut2XsqNtKNrgzZYkx1mTIQ36iWjS4y4quFoTp1OPTtm0vrwSqAemAKAnCnFWr8O
5akZUq2OKseOaTq0R8QhKwj5wf5HiH7JhO/qtypx5VILTMo+jUElQi2WynpRRFINBfCYgZQqICfz
jnsju5npU2640qmwRwYiJHNGzJ3+kMJKZeQWRnxXMohvZHGw99NcA7HzD2AnfKupQEwXDbGXIcVE
iGhiSijBx89wFBiKOrb5ZTD0wOtRjzWRidaCaZeMAvFnF82ioJu9CvR0BzLp/d4Hy/4vZWAN3Y6l
OIAMqzuFwoBxjm5HuufsQFm7AmmOYlw67eXPrPSvSbWxX465Pl7cx4F2qxeDHIazfQSmhsZfTgNj
NHPyBLYcnUW2rP9s3xOxaTsWzw+E+70iSeAGiG1GUew4iM/UCVg0+V/lqFQEM8FVlZGPKzyYMex9
gkPjZyuaViL5f7VCxlpI4IJJ2gVtc7uFaenRIy63TORGKMdvgjiCg8zx3zt1RS1gNKRivfyW6erV
kjCwKRFyPWRWBvCJDGs2Y4ot7t5zjzPkE58xleZ0WvCas+niAGdIPQriDlRiHn13IP4gx/zHUJir
eYvVDqe+950dFPkMM0AMTcbqjjBg5RXMXIGwIXqW6vTVxhJLHcf3y2WEu6cV1nVqRCn7+xiILNxU
LV5mgcuFvLcI7pWq9BJOKgwfEl03AdksWbqLf8EMQ5HinDaJcF88zgjgQewkbxssCxiva5U1Gbyx
L5YLTYmz06kWghPrXdMscyxK40wU9F2Qmg5IO8QO91+AjaMaVfXJUvIRnaa2G8nP7A29t9PeOrOC
lm/e6BBkW3lMlxhxEuP9JqF9R2UcArSzFUyc/J6P4vJ8uT53+A37FjgA+RY1pp6HhkmVIgFTEc10
B7X2N4iXPer4ae1lA/Jw0RCM4iTTb0//phKQCGNT8mjjUnxrTa+r0vig+qXTbDWNajOv3u2+XyPc
12AjFDUL+Fi8VTXpkMAbLojSb9JQ/uzDcsikkTOjjwNZTKuB/6t/G/KbtPJXbpY0Fk2Zr9XL6ytP
gWJjJOdFkWnmQ+FBUdFRiipv2UAsPDkk+AMVqgSVPX4TCZQHl8XBWs6MPuN0qtP+telBmG4f29fc
JlapDB+dEr2zCCXDPkY8ESKFIKy3z9G51YMT/3FBbKCQGOSJMoPPpCTXTIuRvXkmnMX8sU4VmT04
BOpU6qDxHUpL2u9cN22Qb3NAlioSzMEb2klKkwE6eMtWGTvkBPrqZ/B0FToaKblvrKP7F3JFHQec
BiuncCsmHbJstEujmdvd8nEu2rKRkGeBXTwks9XukEVbZZoRzqMRYQXAxEkh+Nw93xGaCPGFlaqY
lldYlYqtPDS91TfLcAlr1RVKZhfQhFCa809RMJWiSxEXedH78YF44y12fL184UTLPMKbps+GSf5z
qcdeNC0jv/wI6/qW4KjCYsJzgmubexAdtDFRH8BsQoqZQfz0+i2jJOErTGQWFhVawXCZ/pLWhllj
yfweCFNgtzpAwgxZOytOXbhuhqRFa4Qkzw0Cc1362UJAqfjTmOAVdKYk6L9hCd9c01DJoyMjQLS8
O5s2X/xNr2mLYUextJmK/VlXqdcimPQyCdtfTOHoj5GD3uOrxA3cH9yXHK2AH1wmMSRwpk1SAvcx
runqZpaoy1YQKkP3xVgyVfM8hDoHrboORc9aSPN/w4J5pQvUOhHuHihvesGG7w/Oq6rRQ/lr2KCB
AF/2zD91mhn8P37mO60ZDBpRERJMzhAmwOJjX3dUwJtWFLa2g5xiCNtzeMCgHJePfaVzn6WtzHqK
A1qfik43R9xFt2UVOG+PpSD1ZzC9C1F959tuJxVnYypnlgX3KgRVeF1+aUNoEAMUlwBHe2p/4kqG
6jy7urUkLG7rKh7QL7aP9IlbbEzYQIz9vGt/XrtfgD9zCrrSlEr5oWY6hnP7HDY6GI3M6VuyqlI+
L6wEPBcg1YpW+Yyu2Sn5lxBcUxqPXtJfvoIb/B54Z6mrWBb3U+MiO4pxN5EsWklCv89Qt07bF5qD
n1VRlUgiwALDPWLEf7E9iM+oOan/xJ8OpmDkixHRhWwuVXjQ0cfnzOEJax6KUy0xZPZAmlU973+a
ALkWICC0cBZ3YNOYumw3tAV/RyzgskFbtD1On02xZw9XP+FLls1JRHyI7ICucBvQVk1MgtNqF2JE
f0fuXI5hSP5fOsHQJUvp9rUvjr9kU0gtwGhTrQ==
`protect end_protected
