`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
aNCWchz8pKjOFLO+GQ1jCi+nlKIe1FO7ADaXcJrtJuxYD606zITAWA3cC066sq92lf7DPxEskRts
3IMoy2VlGAxpPXp7aJRiheEfwPDgOH8SN8fjBNgjwyseEgp2a0bgx4G0cAF4Bcbc/AllBs7BcIbM
GbnCrL1V64qtGQakQa+d46RoI//TBPQ9zwubRQo6Y8VlDGwerU8sKqB+q9Rjg9rNqFO2l40fu51H
n4hrmActzzI4iFr/hEJt4DKLfUiSp2GhJystv0cmN9VF0k/YsAIO0EP7Z1LnZKMe2doZsNZk6vd+
Tr4Np3Ad0qjRAlF9WzU/xkXBR3j2uhn48OFcnA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="du+9l2aXG9f3mL8+mE3tMRAXvNBU11k8f77yPp7ojCA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5168)
`protect data_block
ABO3NVCC0P5+k8EOuY67mr/i9TYt2AiwYZvBPxoOgwYMSdl4yiUQhbH67yMMljmQqVsXBe6kSZOL
gbdbPyumxucHoAkUGtYSuw+l55MzXz8ZrMfVu2JgnpK1+Iv9NfyhUTNt2xM2LuAM9FBfO3SXE5/W
GX9QqZw2uvZaRy00NF1PIXxFqhfDAf9OLVVYDbExqgOX2hwR1Y6nkZbU3Tc+DmhyNliShIUDCTQT
nesYaak2eRZe0Hnc+jYIelukSUMnFxUEA2JaraV5g0PoHvtGsfOqobsRhm2A/2ByKSINjLTIJg2H
C5FnKQv4h756Re0nia5kgWY0WtNKYJo79++YGVRjhUKJlqGdExtfslAzSe2CbuI7KRcWf7tYyLmO
U5yVQxuNQHLCZIyp72PMOTB7zZimJr6ksSky8b1x3UsaBvfsd3uLi6kqXuHokJHJalu9L26YyZ3B
kyKzrcIt2up/YZ13Yeq3M60R2QgRVYW6wD0u1HS+7WLAVZZKugTiKrLZHUQngqwoKLYPkhfYjHZy
esT/POV4YbEajDOh/q1OEGhCj25fVWUj1Fh+4M5B6euq3yl8C0G0KvPzMSsMR2zztcl0kcV+30sL
6pynntzCfuc69/41BVjyd2KULt6dOtVuvcUK5xp1tckhPNzPSWyiI0SxXV52xwkLNZYB98neq+cP
/MhKtO6wCOS/lQS9G+Za0g3ObwsNFh/RofpbyOkhgswxcKJn4GcXF/PElG0n4OqsDFY4iko5KfrC
QwCpuVW4y2yuBjY5ay02NgF86pCeHrETjMDIyvjxXErTMCx5vqIcwqnB5hKx99iUUDyH0zyV7oPg
Wt/WRME6Tv5YQYtztlhINr4TUwyJXVZp/OyiSrxKqG2kTapDUVmbgV8d3sZE06gApAYj+QG6UUBV
CJ0JL/ifodvsgdjFgIPAcHg6tEGgrxfiaI+kOxPwP4JMJNNuUhqzfNUyhzYwhdbyVqC5jtCFCZr/
nq4gtf+ckANCd5fJb9ZCor+3QtAqBm9E5jOCmEPQ7GX9Rq75xBYMEysr8WQ5GlNJ+VTe06NkAW2Q
/qS7LdF61P7DoGUEE2RzUpnMVQimTbCXlaKBPbd6xfgp6W5Mqwnpy1+xa84F1vQma3vbapl7uAKM
uKT1FiXm6PYTXm//scuE7k8OARIOhWIjr9OePzGqV1yXEnDLrK4ecvoyBLCc/yGVemtnbL9wxqXU
vDxvqjIekZyfxUjSh8rDowH34SkctEnCzk42Boo2WNHBrld4nqZd7w/N55gJyWJYMFQH4cEZ7XK/
NTOosrLrGtNVtiQbWMoQXuT9c3YrVrRTUEKhx1Mt8bJk7+u6PwC+4nvnhHvJOxbTWgCaz3BLkZTo
QYf4ONxxvikdkNZnade9QIHR1AJKveJOE4TBq1ieksT9XOshk+BjJPDCJp1nAuxqx/VHvdHKoPBN
KwT4pPo8bypK0890ziu8DNY+Vp3G5xVb/OjH8ECIsnb3X2kqegsfFJ7EdLW5/4JL2WKfDfS7HsS0
KJg/bDwBAAA1QBPSvUTwNpQI/+s4OcfMZ+ujCGB8kheF7HdceiJs8zahPyFnwLmiMGBQbIUNZtQ4
USCW/gwCqPgIdCZFQ64oASL4CbUnBm0ElQp1mJOcFheUqVn/lVK8O1sAvNy0XMkNQVl/myzjVP9p
bsh1cqkWmiKtiibAxjegDnoCWkSRwehCCXIvIiHsh+XZSxIzz7M/MsyloIPG5D0Dw1E7fG+BeDCJ
6NUYI3dIx3swElLr+QLa/S2Imk1AlIvQtUaHjglKPvzr+60MtpYoluutd+Jy9jfNCKpJ4o2uYMtm
Ed2v7yDrbbZ+h4IJOTdOlDzI8fLgtmuBcnlfXiavkQ+LW8QGY3ItgO1cdLJBsmMDVAESeQa1JlyC
YnuFO+hzp5pNVVLgXyuvVRZiANt+xwqto3RywZiGWFODXIhLW5cnxNcNyPWfjf0D1nrj0zLbWSFN
BRYb5mLTDZThO3ndKFKXvvR+lNNG7xnRXCObx9+MvkMHWB1tmjNKeKRajU+eTTI5NAUa45tZHpH5
fqMLQIKBX3S81tnHcS+iEj004iQptAw/xZePwBghlC64eryITHuRvFTEAJPMhvP/4Tuqa5YxmMuf
0LIH6W8ltKCjHL7HskYUVwo9SEO4WELlGRaiAgZsCWirm1NLwAM9qxe2qs7L5TCB69ztPpcVttRJ
MbrkUYq43+Hx5WjW6N8r7h7kOePJwhHFpkTOtRLpLjY5KA8+D52gE0ejPxxj65lE5Q29GjuLGkXy
rfSsKcK/zKbUAeY5sQ+6IdK6cT6cI9bUmFYaligTKygaRfMO761ix3B1xS0TBKqrjHMykOBKks+r
wKHeNgOVbGnUTm5hvFvpypSgu5fTQhvCKhwQiPn9B+EwGjb+i9P1P548AWy4N87ScjxnZC32WRg5
BcIP1FsiILGqv4YMdLZ8YeGxQHZF6z2alrG/5cYMxbwVbPeCR/160aCUZVaxBRcvg2a45DG0CXtq
I8Tm1/WZmu55emX+lyJibQptBmvi3S1pJEv3hjOK7X0HRxw39Cs+rJuLdUXitW7tPfn6KWu9YzX9
XomE2N8X8BNVk3rYl1X7yru4fEwEjZPaEal49AMffQ6fiEhdwOCrg+ZjJCAz1ZDMv+I0atFAxzZm
uaaWt07ZXKox/Ffq5HTDDqjKaPrRqUjTVBs5uAZxmkZFXpwqMM9cLIV7M46BH425rFwNpoQ0wCZq
QgOk95UGMpmmgEjhwFeKkFO2ylMj/0sfWlOBquVlWtAW/JJOV90AnlLwgWKjtyGQimTpcCPFKrjq
kxECa2Uo1uYDd5GbwNHW8/PwzPz0pi5FqKV7UTS0tcF1zpBddnbMoKr/5eVQQKu5yAwLNOsKzQ6y
0Q8qdTCh2+VnmbHKLewf+Yj3FbQBF0I0rwLb0fOS4hmLZ2v1hyzQXoBhSTgY885n++Oe8lqEQ+ns
31vdup4pYQ7Hg66FNkdN9e9fTV7G9fhYmTGuNnT2+KJUCZneVIHCVJL6MI1lsZ3fpig11GNFWKhr
O2HhVgnmVc8PDVNyLelwTta+UFh0sxF2eNq31EIcJC0lICCD/ip0+EpXk7CKESJ2c8PK+1kD5Am1
zZjEzZODm/xQXqU2bGmKvcLy3p4+9XSR6pECQoEkqPgtikeE5E+GnqK3QANNVxIneF6kthqYEeQI
eAPTUr79TRsV27ddHBIuskUakqHFNncAWYCznTjmZyUr+mBwxVAwb3AAScOX8EwU4znfKrQIsWYc
Lvz8nswQR7N/hYPzKi1RrfbMAfyWXIg+veGA/WmK1tAqYPOitsxDoVbJUndHSCd/9yGUw/H+6RCO
Ibe0b/sGzOPntRBFiv9gdn6pq1f2fFHUJsiW7a9G6koj51WYD5H8rYqXSG/cXQaOqFTH2jGLk5tm
qnJRxy+CtHulHaI+/FflBKOdPZwb5OMwpDBxntAsquweM1U5e2qcV5tKvB3Fj5lPY/Xcpmf5XXWT
jOKtEsAAs8fAEP5FuuoqLXAzHlQfFIKSxkS2/M4eGd79j/NhMfui49WTo4DY0mGTTC4ofJqnYDJB
OJ7ypI414Orb8fi0WWsBzII5QOMbue9DH8tW1k3Ek6CRUhXQpout3yHoKeU3bNU74Uitp7Brsb0y
4xS630QFAULd2AUs0ced5KGikP04PnvR5WO02RTfIQRdfYn1MgcZlV/IRA/lbhLeBxaHA3aUU68u
/zWLO+lO+KM74pwY2UXfGlX9Mx4iI3zFeqcWg5qJjBGgoF7hGm+MSIQawSwgr7fFhINieABC988I
ew6b/IY2/ilJ4iOv6ibm5aBGciGCcW/IcVWNZdPIxbeMQO0O5W6ptqEo8+aj4iB1TB0Nw1Go7WM5
gFNCQ1TzDTHQ3NzzBQ8QeST1oYGy82sgvOcnjGdyrcsLH4Pket+DqAlMyHcoUvorAU9qsjFv2QXF
IXn7brjUk06z8EWEp/aVulAo8GIXjmYnkrbdAi9KHm0hBNJ1MEQBVktAnrFaml5KdYs8S17welgH
FGdZnSPwa/czaJwxQBRNqkVOQvf6W2rSgIhGWw2UZa//deV9mh4JiCn6BFpjzBq6RIcfUV8a28AN
1hSZmwxPXzRJoFXBNkjsyanozaVXyMIq9N+vgF7lq5rzT1T2KVkkr5MLSHckD57kfeR1kA/G3Qpg
p0RPKvYt1va0ujnTqOQZi1cIHOv1tbn8L8E5zVuRaq1tfwuYZzUAQobrcLtEysrFpTAYE/P1VjZy
VrVnSsD2fmp8V6hnwPxde3/4if3Skx4joKCwtmNExiMVfuse4mUDa6vWhC7iP1TESl0bNy137hBq
pywxrqqOCNeOzX2hUMLbO4WQLHgnDRCTKhk7Uu+gWvLYSUPtrR8WZi3wEwl8F783hYySZtU98jnx
uEtKXSUmeTOiznHb5ORMkxgfrtcEhb7JbhPbVCqpx5sHH+w1RF/XlG9ZgB7Z59IeFVI7uHkIkfyw
FZtdkHPGWZDh3iS0w6wEU5NRxmpUzqr8rncKtMVSb/XkOZ+WAoB6WeeMsRCXUKz3QBrurVdeeULO
a/Or+3f30SzzN/7RfB1t+yh3/hnn48SxS3LgTwMKlnrWZpyvI4Y/qBeS3dH1PXfvSTZttgRUBUKk
64JlHuCGlyMu9WlZ7e4SVStRK0dMcVxPs+Z7elbD9Td2gg5/Yoq5usk0guAuxFpwBDexbGbh8plA
N1Zg424mjZceGoScTpYp/nD8mz9ACfgydEe9hOqCZ53l+WMMApIVV/DzQBJAtba+mhxxcfgNtSYE
TEIoOAWZtVncVyiun5RoIXfTII7AQKuraAywyub/KFtMVTEqONvkKQOWo5vMq7EjpyvyEysrWtSi
puC5fsoU2eXTpLUNtgU5s9uBaATq3vP+QU1Kmu1SSlaFOqt0GnsiXL9utdErNDAGxBKOJ9rseAXj
BTqm6j2f2giuqEqaI+R/ZG11vnzccnDrglS1Ddd+0cPpzwOs9Ocu9bS5ueH8eyP5BQQzeT9DYJ2l
H7Y4UQFI0u9R683KhJunH+3/eTx1OcRGyUcbb4Tck03q7Sg8XFZa7UabQdTGTwU64fQwDlDrI07F
taM/0jWKwf5R865ZOX0iubTYMqZJn6fMdCd3cXCwR7apwcVEKTXHjsaXjashLQ6I8QTSr0yc1uzE
7E+PmWs7pCVI5a8d6RGiMdywywyEeISiMlJwbAXVsXPosr3WZ96u+zFW2EIfc4qfTJqI7+JDHEkF
isShRunS65Mitz2Tom2eAIpRFK1EcF8XJYiiugrFdjthb6TsO+LQo809fbozibzhkIk3WRO05kvi
z+72gdBhAzH1u+frNRWM3yecdIh+yYya+SxL+LxgJePItM0CBWypG0wD5i3mcT0f+de6ByqnjE/U
G6pH/kttHRxuJQvMhVWv3obL5O8kauvHCXtDYuJn71qW6q5t1DV+YBstrRMpbHbLJ63qKxdfxP3Z
TJ0UIqhy01vOxriT0hFkgwPWxJ1bYZJDvPla7wRwF0jItwK6QCip1HzhJET8wA/voRGuS1mCEmxt
+p6i45yHj96XRyNjgvwYtO3YRGiqrTTO8zNZ1jsBWag6dMX4xddqKbGAaqtivCqDTN/pPgfRULiq
7sMaYEs3spaQypq3Wy7qm11AGKw2EsJp+e+xRsJLugU4AM2GAZbR7Bx2/LTAuEaOanSjyVU5VwHX
AS45U9H9byQQVB/ro1NwcQALDoMCMIGn2ovpGaNTHI2CCAkJsMgwfTo3TApqTMSjFjs2idbF2vZp
4SdwWMPmIFxQeGAo8UwyA11umVskjOQW4uBZH41+yLQ5bDSqCjbapeYU5zjslDYCHjh9vQ7LRvCC
MIfaGwju/4q7qiCz7XT78kG+IYfFaHQhkMwXBXn86anNy45CuZeMChEqgn3g14yRBxShl2p2LV5f
b/qaOtXztGe5jI2PgEwcfVDJGf1EQPsTjtxnkVnL9xa2/blzRAiMT65KFa0V7WENtLHNO+ahhWEz
lfuI2fUUjsR3rUKkO0NbAFVHbV8uX9YGm8bdL+BXw1Ivg2ibVZB3jpY7LOWbjrwqknztRsYHoYRg
8DA8m4vGHt+f6l7/CN9H4joedIpqkS3CZLpMiQI7tlJ56Mu5YPr+2pAUTjNpI02hodaVLcE4ZwKc
ePpkDtUqn8Sdn4pfNMjnrsy3E5sGIhC03IXOrk42sRxH+svy47uOqQg1mEjx7BnrOivt9Satxq31
+M6bS35w3k6T65LudvBaE7KlL4iLRXYajOd/4WYcObIvHAZp5dFm7CcvdJeeIBBPE+Nnojk1huZp
5iLuzNAVhHklrp5xfgJRXsq2FIDDz8mdntVXnsF1GyWN3m2UkEvHhlobhUGREU3biQ3mZRfInih4
YNjbQ5ChGo1sjZy9PglF0D8zqRlIDXt9Ydj0yMLmv/0j5mcIwncpXm2/5YMQNpoXX4WTC5XsMOHS
1qVLEdn+0H97oeofw0BxW9F2bGm0wlFNmt5AQgYfkSiH7Sgdmo4lim/bxFRA9HGMR/R21jbT2k79
O959uG+F3N92C16Jnf8u5A+QltH8mFfuE4r3F0lcSGDYRHwX4gWWkx1L5BQ+F+8ubPOQhTEHrxUU
twEeI4J4DkbfIv/GWtywFrai500MA3I9+CN8D+lf2olJYNYdkWWXr8PBQ7TDGmySB2Iq5syDz0CL
S+FWH6IJFNLhrqJnBN5uM6DK7ZYWP79q8yEGwXiMPTPCI7oZ/z38iB06FHzfON7rlS+JRQcndBmG
x9klgOuArgc7BxCcLQsD5HohHs7PE/SDYHZD+U27vdHPxHDGKU9Q5lIH7tDfvzeQr/zVY4CMGB6h
z6eUP9yE2IIM4O8pNx5kElX6JG/i4BPQo0jhd91fcPSMUVFYxpI=
`protect end_protected
