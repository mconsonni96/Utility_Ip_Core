`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
tjxQARN552V491fUuwecYUbcbkjYz/L6Qch+cdOhxpAM1VIcUK/2UtkVDOaYcrGttIE2JTQTwGqL
40oPKJ+a4WSrv9GfsVaPkmXGtusJthFbN6mA8h3YxtjgLRDOqJ3wTQvITGlYX3iofPHnBNfsGEpN
HPQI4rFIra8xfYNi+78slpSdVfjmhEbBTZms0u085wf6Mwxe5Ei1enSMdKYVz+pt6lrfr5J0bbE5
CL0odK/aiV1hJfC1Mb+T+amHnDVOD4ZcjYIb2wvfaIXB9IO+U1ZnaSmPMEiEqiw4vNYJmB64qwr4
il6fErMFOv7tgwAZ4xk6N7okK8llcnMaixhT+w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="nysUjphz2BmEWuPkpbWQ+c9HGi8JEt8fAx0hDkxvRNQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9488)
`protect data_block
Jko3ANoDWmvPRkomQ2+J9RBXIF9MH2MxJ9DRRVBaoXFhkLG1emNMJL7QqBrpK63mm49EZvZoV8Ta
KOqiy5IHUGZWIAFnL1LDyLbjSjSy7ArslRtjBbQ9yL5b4pEeoHyPvAmUlgr+ykNaYIBg7jcxTMMA
89UUx1T5+eTIlaCRQ9fvbBEaQxDcUVU+GUfKXSjGcsyh6MtjB1wBH6hz1RSz8jEohvL/UmOB2Xvh
B9bf+Ed5DZvu8lNeHQCccJSFSWx3a5R7hdYDjJaiF45MwP1Oi6VPhgsMqQgUvmNaDt4oP/whI1Eo
dKUWlFiusxHT8r7yA2EaNwRLebGStbcqpU/6FG4LuEymBv2c+Hs/G8UFz6MxW7XUf4dv6/wlCnol
Q1rJFaUv2pfFQwNEkBLN4fDV7jMBGJkJ8VogUTzT5yuENCCuCDnRGJa1cevkFDCCSKHYOEQBB2oF
578VZ0gS/B05Gh1TZeVeFIdDVaqi/dVJFE28VQP7inDtP0dfHMPx6YBOtkqeLTKtDDFttE4ShDb8
xeHB8Fg4pEWdYrOfxbr8acBAs5NQiS6Y6BRFSB+zQWuyensbe8KmBEej1tGj5YWOzMSZClzvbeMf
AIB/qnxsRCMVIdWV3VPWdsnPDgxrtoqvP+MEuiCFtPzZdR1gJW9draYu4vBrwADSNSnHIxOiiFmm
D8A96O7qUzvwUTN+JM+noGnWl4qJqCj4KDgyI76fSq6Npttm24daoCWodkQ1qGScMznk0mKYKcdr
xeVka1WxYk+Gyb0LVECYp0hZYkpNo1kT0kFAqm2zB9lDl5R1ZexQcLQ+lY0qiUJdF4ZIjMZAYOBE
zZhc+lMkeQx03zs+u6QqCb4AGusQtyCbae92km8LOnjPNlwCMNBdSYJg668vb880uDEHR2iAW5Jh
OSV0wv449YpnfOVBKhi1bsdnAvEKNIniPVoyIYNQxLago6lPpSdHCbDi0h+Y8aGqVU9ma9GiuRhO
7zCY0UzWBxbyw6PopkSvWkIsHwVEShJQQ6ZSv7DpMKGTHsBCIqReCQqD+R6PyyPt9feXxvNOKtWJ
SKlGI/0879B5Z3GZ3jq+c5lk3Rba5cvf0HE3bXHpb9we6H2sc4oHVkMwUTMn9yYEOBReAZ/Fv+4k
6ZgYA6LLH1lpi1AytyVPLUPgOX9Pug0ranEXTl5Pr72yQ6GkFmg6CZKszJKji1lxaJpUP6TDXMxX
uMTJjueyXc+fGx+W93sZC2mvNZirtI8Fm3S3nAkVkvvoMMfq4GOf4JE+cK7oY3xmWqDswAgowFiA
nGzhxdL7zSgJurCsG15I4z27+85w+Js/q6VUFr+SJSq9ESeyKJTWrfE6YyJm+5CiEQvi1+TVSrFQ
eEAF+smQB/qCDkr2dRXOSZBSTu9jFANlfsQfSscTERj7+HfKLsoJwUzkPV3Hh2RQcNlNaUqmf8Me
PbXHGhBEzk9coSl0RXiKvu5dGuXgCVk7pj0Ln8V+TNJnzyXSlWkLwGkqtlUOwX+HAJ0TGSx0MfR9
t50Zd1Uu6JIAWCxTugrHQpwYYw4Sxi2PEPdlY9g4ORs7FYwnsIN9ga0H7ckqax4M8CVOMhisqswK
eLeJynJICBHdH+ENbgtzriUZdbuaYlpJ5/kY3dZDcDWUdxCe89iX+NoGxrAeX5eVnkuv+LHXypyx
NMFGPE+f7v7jxLg1wuaFNWNqyk8VAvySjAxRSqaBjPe3o5B5ZvGpgl5ZPxiBbrZg7FbddQHd5K81
P2BD9WhT/aiJAff/GK7gkovFOSPhH6Quo7eGhhoLkUlscdeV0BVTvjxQxIA9xYnggzUe6H+1DBrb
RMw0WUaERdYq6NKTvJfB2UWrEyl1lMiqkvJCYAQWleeVXg+pF+O1/qZWOIx7tBTOHowkNQmhhTAT
i72PMD8mbmaUxAydmpiVxUMVouTDDyBLP4D7auKwZiTihyWSrtxHG6ASXE55j1U/YYfdR0sfSOml
Cx/l/ErbN5fSBpEDhmfdWXqykzZMW8vK3OiXtQGowwPWTDDwVOWCeeEH0VMRdWGfRJ0zp8FWK2D0
3liRc7unWP1fZi8UavKcHTZCjY/BD/d3rw2eWjHWq8CDiClse0HoTVma9zFbPURRFeAmh+A+ibg1
e86QqdpqMti4f0//atSm7jZsnW67Z0Hm7w40eQH7E5Ca5FW8FVDeA5nvrvy7HelQQGOgcdjbFwZK
tfhfeK+X8evZWepIy4hap8vs8ba2doaBNAzmMYuW8jRdWSHPbcUjx4sCrDKUs/8b1+8vBEWQI5zA
JtYBa8DCFF5t/ulfRBgf1mDQsriK90iLaV4d+B0jiHflYmhyV7wyhV/W6wkN629jrV8FMh6GrNVo
OG0pLlL6qv0Dtu3zAoSdsnCROuMWinZqRdc3+aHf/fShhf2ljyapH1gDdDC2W7oDo3b4hAnoO+2i
sc4MfFv8T1bAby74y5DsTJX/jfaS+3CYF75tBw2PErpoG04s94wgz60wZMTWU/NAScUNe7Ou3iQk
PN7uTO3mg0p7Osw7t3bwzR43I+CfXWs1avhWC3nZ1DgUoxLkzugcSw0RJXwactljmD2T+n3PcOUs
+pHQl8gcbNpsXye/pH8q3Arfj1PF1YQumY7N8Hpgr4+RMC1RVKeW6PttRQDxm3Skl0POqx0pY/t3
zqdifH4RO6MLRPzddEY6K3bSBpv4QYYrrihhiKF1rEJWN89OphI7i0euIl1PCnBdv7bmM1a1C0Ml
I/Qp/AN/80Vq2mvZiZorDtIa04XDnRK9Gtf2gE6OCiVha89DGz4gnOyysPwNIHqBVf/GChSqlJXP
K5jryrcn/Jw9S/C2g5o2IYRz8su3cWYOa8Ngidr6j4uBgw66vTs61jKhHpUiPXQTwik3plyGGCta
FtEa82Uy51Gby87yVFVDOW00LluvuZCrXhaHfIXeDb5sI3cWDPaPUhT1CHKyZT5m+h1IXTnKZQGS
vz/fh9aBDSmqWEKQQjctAgiHKKL+BW/wmdy/gz90iYZC/T6COrRosXGgEtmRpRl4Ckf3FBN1mmM+
1W/6KnQENqXw8eRZVwnfCzBjkkqz2KKA7hH1kY2mksr7Oryf1qbu/IJ0fr4XFFtKtv9uS30afYJJ
tKSE4CI2DxhKKF84h+UI9tjWeB2z5bSG5AGQSbKzPIwC/X7jxXUO+poKddtS6rHBdsbH+5J45l+b
zNIE/dpys8UvTMnqqSa6cfYHd3mray1bmiP4q2kO1xKNhw9QwTaiQzHE2eABPvoarT98nMY0UmK3
VRrfVOb0TqDg5u40Yx4Mwtc7Ild9r160Txi8G3w46b5I5XlacPn5AYWLqPdgfBDVnHFRxJn99vQf
4NqlfV2mZimL+r2ADyKDK9COvcy9bCwhwanevOWmSF0IflRJvpUPmU4BWhSmZUoeGpKEDcPKUN3k
aPJlCnMJntXmjn20M8vvE9ZK9SpbfjivOUp1DiG7efFkGz635wMZq6UlPKSPcUoWRlThhe035UIr
xN9doe/cxQ+gcDNtSdMfyDCgW8yin4uvRaJhAnQ6kA8bCdgp8RDZUm1HCmnOvFAaNtKLtwHcB093
9XlQinY+gRpt/M1ikfiCHVFtVvIRKgh6H84Nfg36xXrD0XiPDbIG2wivEgrekNGA/B20i03qR9k+
ViYsqvOiwjeIKCitSvC0WEcKWWU842fYNwcCjYJgBCSPi1M4FPRNKx+t1cLfsCMkqRf1BVGPZjvz
z80EPCyz6Q/yJrG9chwFBdLl3LKK/aj9QEYnpESBWxqBdLrFhyzzREC49NMbS+Rkt4h3CvRD+A/1
3ESZHCjfVHH/3W0IuyBQANu7mi6FWx8vUVACtIXYEXXP8KEl/nMPkis0fBktLkxMeAELL7nMeKcd
YLsm0V3Zp47RY6PTeEcNjc02/MtVvvE58NRYIic+o5+orFWGSMAnEZXphXQ4fAH5fQ/5ikSlASdF
RCkWDk2OQ2mJhlgVkPOVI2KGwHIZXBKsESDfLa4ZU3RfTUN4OxprWnJBimJdo19Kpsuz4Xe8i/Go
OkQMESqtxsts/8p+bLfiyfSGF9B868sSfCTEXl9SwVxfY8yhN8K+hCEibMtpGa7VWlHm3mNjm3mg
sbzspnToHROzUPpbqUTrujy/46WUAS8lZU6OMolDURbYTaaWAiJh4jHTMEpIrmTlTJS5WEcRlqpv
vaGtFl4kqgXK7EfrVlvFizcNlYyR4VEC2Dlh/w6uq7ZnvXr+6KS0bp+AMxWZVFtuU27PTMtG0tK3
Smx8aRa76xCzeLYhQyt5zzrpIal0nEZlmfyTTaS03+l52RacVI/ImqvsuCpVYIphJHMBqpiq4O6n
wn8VKtX+nuv46JuSQXkUWk67k1d5vOJpD9IvLe6hheMVM0w514D840brl+NILbXPlUThykEqHdYZ
S6bGJ9mu7WYhp3hSh98UBbtSY8e81InR+g46cv+8BBBltkobJUeIHnzIipSsQZA1ktaLa6jFXH3b
p6lYNEheqJs+5rNmaK+9y8QSJ2hOGwzO7djXTff5HzgMQ4J/EktZObK6Bh68Q5FHTXRwEaD/aKX1
wk/5OSw7v8ChSGxWY59P0vUCk9xife/vBZKFnXl1VUhk663Fwq+gMSa+mqwBQdI+GGbEQE53IkM7
rSzt/PzQwgGLWGohEiaq2aonvVIspMsZzMpvIr6BvmHXhC0xLB/uHa06ddNXrf2JrAUsHxclIAuQ
ce2q/TsmuTs4YVMGB436GSJiL2dg0pgAMXATDk32MNZ/vKqZ9uaE0PSm0BOxSKOtuG7E5UvENMTt
W8yYaaBeti8nq4C6TVL1UyEiDunDci5OpLfv0B8Tecqk0BOEnApWILHDuI1ZL6MouwMvPX5R23LT
rv+KJ9Q/WgWbBgg+T9YoytX7qulFfLXuUkmKh/4LR+aFmaGXj8f7vdOauPNuQ8a5RwSgCf45Npl8
kGqSMSOQUu5a0fibt8lkWe1YLn0aZfdIaP17OPxISpp0kuncrdCMT5gz59i5mYq6CjHbJfB8FIQd
AN5br0aOaRfmBGMir9+nWMHEnhHYNks5LzxPkOGNXae9E6MI5CqjE8b+4QzZ9GThMGgIyV1dTfF/
cWsMdt+3rrpdzVFtrqyUkr/cxft2zpKE1zQ0ORO1AxBSux6haFi1WAVBLjlo9rcbCJm7zyhtoM8B
OTCqVE9x5LHYokBqznUwfXrWSTKdRmwP8f3ifKIbHa2DOp1xi8oFZ+cARaJacfikgwLRLuJ12F8O
lhYoZkrQal6E4oy7h7KyHWX8rz8R0M+5t+tsW/jIZBfdun5yXQ8HYsTFKtSj1c/sLV+h7BoWByuS
MvFLZ9klVspz2OPyjOfTJ04IhT3KVRwoS9MqG7PbCavh4zkHmsx9vbvDbSPiiTJrIQlIEADVDwNg
hBGND5Sx0PNvi8UYxUCf+oTBfHI7sDJxVJfGdeYZzAM30rkKEnDLtLVHArBpZNvxGdPaIc7u/1Mz
HiPk5cb7lAdvsmtCg0uIa/mKdJcjzvFdwAH1OIXy+DaY31t310byhKvYPQ1TM10NLG4sc9KgVHAH
7GT7Wb9IP41AlorDPLfCb7+mg9ot106fLYIhc1b15IRuK63wuJBpSzjR5O6ybkIVJD+RdWwkDhaj
hMrjmzUyc2j7ZIxFhS8D0behbkqsctwLdX/SxI0tXHGVEulHGClTfMA+HhIdZVceB3ymJ9QApVLd
mnMTvk3HGU4SutZBK8o1CXW/s6aRQXwYMGdy4rFPrg5Kf1KI8yqc4RPXNjpYoMeslrivcSEFgH2A
bXcYTYeLCELCCKCaz7hdG8gE/or128wrIOiRyf3ET+2BrE1o27R7S/UNHG64eVNdTKJ0MU8YdNbp
ed3ybcmwvTuOq2x9VLrLb9ct+Z0/Kv7dZLcWKrIIdRfLNOoDxRYcxvqYbhEQRO8m8z8XIWS9/2er
V7JLVNO2Pmr5bTwpjrYH3P6wgf9rF+UK5WbipFucTzm5BOG93ciOayJQ3U087JVQ9OBCMqOQjsjd
MCXBYJFMCVg3GFESiQ57KdvGaWXuGqIX/EOj18XGbx3gRJiKXrasg05W8YubLqoexW0BIvcW9e8W
EnhABQUnTpeygfQ7LoQqELb4CYgNdHK/AQ1+cUCdMltut7CQAg0j2n8dRPyGRTGPZsM/NG0FQxHB
rftjiAI/T20mppYPiTbBMJJqqYaon2RpaCa2pWLo3SHVD/S556ij4qOD4xeJYPfHv82qA+0W1AgU
+tkuRt9cFdsTJ4lprR1FE5pFozBZ6pEJPP/R8T5MRnCAa1guAse4RJ/Msu6MwtFhUqbkr7QHiNUS
sOaIXRt0R8Ds8Ze9Yey/HERc1hC7Y+hnlOXA1RGFuqEAZX3fvylSNm50rEmVQy4JI9+vnFqXOdND
p8KFhFYcp2dTsjlbSSeCwyE0zjZOE+FuyAH4GeJ8ceylkrjtgQcbjF3SvYjYjIgPhN1TQ6TNwo6r
9LW07/atIN2GGGQSeKDs34AzsGEm7hwLYd5aN741T/R3oaVPgN1FL6V3gcNRnuEoqMkvVhljSJdN
o5S+Op6aW/UThYlGmG1+elbgCNZm+WMKuxf4rRUBDaQf+RUlRpeYh+RipL8IFS4Xe+0sDH4HMj/0
CCn6Q2pPSTdkisKXBDuMgN2JE4c/FKVqyvOpZuhnvUUz9UH7wyYsRZIKrwy1i5Y4RmDd0H1I2/ZH
PWLsDCQCclxQ9cCbbeblfnj+nTj4fwPUZWThmFoRT37AolBXc6PKb07f9VCQuRdfjdhhEB/yTraP
fBbs3YoiBMpX0jg1x1gxxAE/YOCvXCLzUm5D2LBwnPM8h4rVKCu+LPT/can5iUpu+96D2A+6qQNS
2ikUt/spbJClW89BolqTWlp4JLQ7I11m/SYPHIhdpiEVMHFdYne1qWwkz6+Kaha0VWgBG0s1YmTk
BUF08Mfm7ezu0iniFgUpRCsI5rXlbNnn0Bj2dDvPKW56tnofgTC/DAlUrJogZ36M/j/11hLkFCW9
NCzhL7stpK3p+pbKY5DYdtcksdDiiAMNQ11ozQN9/KeW6Mf7RCyaLopsoL8LV1qBtnt8cNW0REZb
7knYPD7cpKTBWWMYmbiHF0yH9qual/2Igzk6JVGM/MTUE9NS6LQbJlJ3Vhd1GqBUssFX9WK4JtAS
u5pDGECLB8k5nhuXYBAdjKF8OzEi+eZnifH4ItDXSSwPnWIY7kUxJLRZbrFqGnGBs3mSpzUBjyh1
lpkZ+30xF3w35F3iFwhWbeEZjngCfV43mnvE7NHUixF5BW19EMVFWENy4+ZhCngUPHY+NjPS4Kw7
zd3INvMUFAzytFtP8rrE8zH2bB5/0rHKqAM0ShRXUPtKG+lHUAzJEGS/skSFkxRRP9+w4W27sWQ9
SA3xJJiIdbuSIpiI7Z++0cG0HV9V1AbNsSIU/yPEh9ZL0jDPbrbCw7wZx4e3WTp3d6Z/zPO2XPEj
lhWaLNPyH2DC3rxfkgTn1V3DfTzAH/cnpdaBTcVcdaqKcKlAjzr5DS45Oy9bpUl9xxOhc3SeimtC
eRxOT8DH58WDWyTPMGE2Ty2Oa5kVI0JnfJHli5Tjw1isQ9CnP+SDpxEvlppTiN6WzGB0S5j/1ofO
kjeksZzd97mce34iq//nAGNmMUXflUldwGuWMBzsaYz1G/ITN6oC1z/+awALOJVf/cOr0Op3b3/S
yh/v1yiSMzhHms39A4Vfdk3pXgqxO43C5WRCsABZWs17qJIhtuOrYreTJ8AdHBe5v8Igt3wxmrcu
yMC25e7uNTkWMwO5qcEkbmilRJNhyeeAkOJEl/aRYverqXx/t2oK+TkMYy1s3SeNXSEOvyUliQj9
AXxsYrIh6HecqIHAR+KGwfBNf2iAOAH44s/VULwyPGmSIYNjWTC+zFQse2u0Cnd9NImQCdgpo8ah
luek9hijMOr+qpsDiY4Ct+ab5T0kMd6+jESgYR3cTlhb4jMrcxyQqEBkfiZEjJ2S+pYpnAyuW6jN
4guSJWf1BSRwtDyIyUGSab1h1OvSKcPitBr9FtSs3IQkfFKWeEMM62DFV/S3tbxKuCRi53emgJxc
EIcE2R5lHpPc/A7dJYbbXihakPvkTLaY1bHatu6iHHrN0oEHJf0hp/7azThngZnqxUTqWDiDwdyF
7/ADKmRj0UIdz4/eniEcbj+XzQhviCikPbdN6GhIdfwSfQ1h1P24dCkeoJK9JkKDXw/Zl5+VFhk0
RwHI5YzOlO3JnfxiwtY6gsFvPwNlspx3q8KhbTxq950DkyKxdHbNGflj6pa92ZNifywGaOO7EDrY
89eZ0EV8lbDJqmRcc/iyvinY9lRR5UqzMz6u4RqnKQvIkmAoWBH9f0Oi/hULE0010puso2jYLK+d
VJlF4qfum4rfQ5dpGXYfBEptOVC5NP6HcbQ9yySP6Tx/HSkWXf5VoItHi3NOMMfYNQroRB3dQZqp
xHVb5OsffXIfdbgUitwGwsIOyJtAEU4hLasMdJSB4GrgpaYMjPgolKaNMtSSyUWKxJAJ2PgJNBKr
Nq79pvIdKUezXGfn3FFHAn/tSOalVT2sJF6/RxNu0f4r/2XjXJ8roD22AckMKzxBLflJkafJKOcH
GPgi6IvfAFUF9t/lm7b2V9LAGn1uD2PlPkCB0Mv4IphXlsRNkpW7qCqvqIv0zMnyvFYU1rOnZDFm
pFoq7nzsk/Eoy2fnV1uua4XCge847KelXs9RyrC+4jhcGz+Pt4q02SjOS5f4FKMMjBCxXTWUSj/Q
FnH5Q+x5rYyHpK+PQFhYabzh7LPBaqHQJqa2DZ/3z4NEFJY+Ad5Rrn7Nv7w9ipo5R19qRsS8Wr1f
uHqBo34OxFWFor2ERgLev4526pApmKewrOvubo0PZnFoWPcZ62LBwV3j+fKp63PyE0noDazjszKU
euC1gFE+SBQx+g+yFGG06GY5HzwGNG9LYpBy7zkyZoNKt5LzaMCJX0m25Kh/BHUsXYuohqIVPykW
cWEFT1Rbbyy8t6BHetNH/vR7utkyjHHfVia070IaWnG9oZDwSG4QD+5kh0dLIREpQSfD+rKh3Vvm
1ene+Mzgq1ieELTHovLCAmWrW/3bj0wU/RXb6GuVIZL+lEQA0vDPvBeR7QJp0zXw8mt1lANJTTv9
LF1yXxWzr/ztL4Gx5SBe26R1bE+uYRCK89S+QKatEtRKUrwJLBF8cbOmLCh8PdNNZHLvmUYIqbCj
o7nO0weSIiMbCWMJ41qfkLmmdrQfuc1+ibAktEXNXX2vPUJOmEGkSBzkhY7uJYVHg9nmcLzuauTN
3mOUQRz9uWCavAgyL26x9w4prOC/RTAD8sJx4AGuy7rNTE3MLVLzR6e+7gCzFz86UROpoawbIS1e
c+CXnhI+xrPT0DQqofQZxombm3fmTYVhJSkmud3oVgU9q5GRAeia4GYQ+w1Xc7hooRwrcHLn7Uih
jXfV4sqLDWaMK64Iu005kb/Lsfrqa++glghw4f79+t0TtGR0NhWrowhbHvjBfgYbw7N+Quk94TrX
YoEdSZI7o8Hij8qeNesQRspyCldjll+b/YxwIkBIgrsBL1dTXGD71Va1SKX6fZwRI1mb8BCate0J
k0ZKQcOquqScp5fMhr0vBb/wGQnq7KHMH9DB2tNeZHKxOrHC3GgqG0BBdtV5frW3prvGiiGAnGgI
mATq+tORdI8zcbcP57ZsFuEukeGKrIUbTDbGzi24ONCLbyMpNfzaiuReRIkgQ6jD7SEe65gjSUao
t/UILNa5h2Sb7izuCNwInf7iYo16hBatmcLVO0jUyG5S6CQpCl8HQKSC4IVxHoJkObUz1tgjtE7x
1YVCzcr0eMXQtz1lwmNFFneJcmuogS0W4veokwnWAlb4PCY5UtocjYHPjTFTpJ65AzgFGxdPBt67
Lw4t/ilf17R4CB+HSXVYsPhmP9J3ofz27KycDHofV5zu1vaBPsiIxQXf/MnyM81fEMLjsBQhC7BT
sfObBaahTo8Q1ua0GE6l7TVhdHPGBX5JnIWbtMSjDEb8zxELiStpYkk9eMt5iuP6UFOBtYF8o8Ns
F2pKVDetu2bkoZJ96F28Sel8bLD2TozDgtZ1y5AzXf187FEvvk12recil3jWT0smc0+LusTxTrFB
KLr7Op6ay12dkQ6wtJYMKYgtMnyWh0zrdn26gotFs+QIfsTSK55gsL6I2bmCHU9DpAGnkKg6nf22
H2pK7xX4hlyldCbc/SvcMiWgMM1YNXWbZZ9J1rxPF7pPFh3QdwI6f50mAvL0F0Pjwl0X2r/x66bf
HDvnmNJsrot+ph1zDnxYUkNdnYlbbb0TAFkFPlvpicXxZ/ZsvzPctOD4xbPlX9ezrT5wcp5mLjC3
/fHhntnZw8m3bBrgVgcjCNLEs8jYkWy46dxkasYDiyWxKkJH8BT8zsi+h29eIaJiDcNH/zOQmjOC
psY8k+PvZu83LoCaTHBJOBMiNv78vhZHx6b1+hcU+ZfedN1wR9mC+3sv3gB1hoFgphi7OPmVuu7d
+p4St9FY6Rv5n10aKBAtkFyVjTq9F47l1JcNdM8hgHRMQjQ/kNgT1eiH2NiEFOqhaFm2mPzh36tp
Q8djUcnTHCYlSomME8+6qgoXoEqVXDl3onSO1GUVAhdF3Mkihoo1h+X6vuY0InSWNe2hhnpYTvIR
Mm4bbznAYtlhsU/CUiMuuORnTttHXn6KdC2ASe3tlRhgxWbKV91MBce9ef5ty4NOwPjQQBqo0jE4
WCORpz7/ClfANoJxO83f4/F95cV1I/XHEBFX+Kb2SQBnVrI+PNCuZuVijDPPZSbO0oqLvrqZAkeH
Rbp6aZgx9KJy7OWcaKKWJD744RIxXyO69Yo8OiDgVLg4paJ8nhZjFyBwlCeqsV2kJ4fXNvyyJ7RB
gAEflI7dMusgB3MpZaGHQJduJ6xk5jNehC+K0gkWMslJUbnLeqlhpKga02vzPotto8Y45rf3qN64
UzVV1xXMgIi8ooXO4prdqofH9Ae76wChKX4pfCJ0hlJrtYrtTX42PXLpPYnNNg7LGKR5A+RbdE/Z
1qAhnHtzX1q1iJr2jZn93OnZAMgBqUChFRBXIwsQc17zrFyRqBcmRJFX3fD2q/rVJFgwXtnKz5Lh
Bxm/FgdKMnOG+x8pbQgQhOQeq0lhFXrMZG+Gu69TwftqLC3J+TWZbHDDkgm/J2A3ahQB0vAo5W/Q
b77ovyQQDTTxS2t65EkklXJfNtXimrc9LSUgrduuuocJT8lpNPnooqdS/kDwp6/y4scE6HoqYNg6
1ZYH553VeoE1uX1aTE0NvWjTagG4BbiS4nYBm4kjSloYK/koVLZJFNEX4cmHPAR46JBhovzKK8df
zX5hwkvYjqLxR59UovKn/73oWBSZhYpP0I5U9a3gziy19KpJwuq38sqOizTUKuxpEiJsEStwc/Xn
WxNm/zoyfEwVlpGeJtom/ihzM50ixW8gn4Qrz2FF+jZlszRjqeAqNZn5U21gN/hs1v4ltrtyZzwq
bRrFFRyPuEQ7TgjTj3lRzQzDdHNkhgJcUHlSHf4ic29DKBs6OUflfRR+L3lMZdNyHaQS/oURlDTg
RJL2fXAIB3ZVWSciuHuKGrslvvDLfUNNFZdQHsP/vkXnMTUJ31sc8kbBbg6v4MPISQ7uumhJGmcB
zZYei0h5Q5RG4fboFyyaH7/af2eJCnWX++AQ/+ff3vp5U70F5ruyuC8ZzPPafyTmAWHEFitGfZic
Qx/3V776TxBf1R9/Pgt0h2cOflFEIhWnU4q+BlkT4iMgkoPTpADsFTEbnnQywXtUwd48NqRU6W46
Q1rqTu9hzLE55rWqiF7GCF4bRs55MYY+QTumFLSawg382nB/8kHILXF2JTrgLlkzXb2oKIyqLqA2
wc6m/JfDPWcCHdOacNXR4z+/9Fip1ILIQop5QslNAWQT0L+tmknz2fBaMekUswpLsSFe0fvx+dsp
acqWQbb3c80q3gSIQ1jsxX2luUDxcqGLVxXMQxuLavCbT48E71Q+y/9HmvbXdFDs6uyfXpoj9tjU
6vOwaDjuhiyPCJObuIuRp9YtclBQf79KJDnMRzrHjOL+VtHUk2O2IFxUzpnhut7+QZis2XbGj+5e
k28lK+KQzVPEH+Zr6OCO7hzJOSJu9JyAxt7MeqP5WCF0EKY04T+s6SDT67eWJH69DozOpgdiThyJ
Gc2Q+BcDOeImJHXK74yX0i9d00Vr1TLd6a/9/woqZZXWj/G5iZ94Y/MZegl+Hm23cpg2j4bSgRTD
b3N47gCElVl8NitwfWCzm4g3tTAUeT7uxJsv6HRQ3/dZSkkFkYgHzlLjK00oOVpm8CRJcpB581ss
rb6x7IePotFOKHvGvgSNIBcJ31LY9Nmq0fq/VDfAkvx3+nUr9GQU3yG02+ulcKeQGSl5ws30vSVP
tnSOa/yHa+iwEwFnHN3UpA4xbec1MQIXcQR+SOvKqWR0qdW/vBSVseXcISP32Tdf3KKuqhe0m/QU
eO7X2VsuFt4K9xbCbm105V+CEgKdH7X/qPBcjy68uJUT65rDQVqkNZ/cEtOTaR+9y7WkcejQOoZU
duIN52rPiZlCXcJtZtJmgujPrbecTRcrdIx7vxTQ3/GqbDfWSaAsKCYRsRsqwGOA4mGVbGnciKdW
OoBKU5u05IfsezjFdXasbmR5NnCZxuNc1UU=
`protect end_protected
