`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
HqAOlgskHC3C9pZHUzRZxqyYWzJMSCYleFCIFgsDJFD+Ms+N/CwxaCu6ZDJoI/tA+maeWq+9qECH
hKZBsOhLyaFlYxr6La+3k6UlQc7gMJ96ECWPOh9yNk3vgFj31HqGhFekQ2poR0Gy/6NPgfHQ246e
sM6WrFfw5OppKvjf6RK2+ejA27ICbv1eMLTYWBb0Rm//NdCYWfloIJFMNbltMZghpAhVO7HJysTU
8+Jp3g26M07wRGR21CQrpX9RRSPnNMV2ASVb5e+bH7AyfckfdiDl/SRVxrD0Ezda9JdFixiHvqvI
+E20BK9qAPjXkh2kUqMiOnkrjkj64+vgbgtxSw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ZZEn6JT21Ie+mjffMIEpCeKC3wcJyHYg5Cmpp/zT7M4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57552)
`protect data_block
4yzeoxVFtby9q8aeHUY6yu2Tn/aj0qp6s3Wl+P2I5vUqvYCpdM4B9eAKj5Lssv3PVGKnw3hf/64L
3T0IiF/FWwzwas8fp+wyDuJqoEKXKODOSLNdip9LEJT3uoGwX4nNT1pyu5cwdaw/Razgl7h+Le1K
nP3NYv5c4jJdnJp+RU51C3SZsUBdmT26qcqqMiKTpkKjxCme4XWNI7Rl16Up+cVBWjWRtQv3qQIe
XxF/wdoUAMUVACKd/xC8GCCHopXREboCDFXsMOVjyoEmVmT6XatWiHEKxZAsFSrfxmJ809AkBvUq
HPDPrzYo6zGw5vXJO8s0Dos6kNLa6PeJeBLBYBsGaZcu5hP1Xss6TAdBuZ76hMN0CDB+8JO2jbMG
WzShZEZihhtinDXcxccw8GNCTLIX73lLzNsYl7o7xv/uwLRrOXxx1bfaqeer+YKd6kvRq17c/95t
HRsh8i8ZMgDFB/HqXy9Z10mZ0dWD8QqvkOaRhkb9z5sV9R8ZKSs+x5o0FqDu8UP4UGE91Y36mS4W
Z9jccXkcAZ4h3XF9j2ZzrLpMec4A61ZXqfZsQRiExdj4mxZ0AhphE+rYg0SlroOtpN9tHTjsuwGB
uo6KXIefVUd9zh5hmnqTRIrg6jvrK9KsFz0XN8JxpVWtDjr7Mf6I3OtK4VTkLSbA6VCfFOATDzGi
u2rtK72dmPSGD15AJnn6i9uCbOSCY2cuhsMdhYcalguiCA6TqSdvJflzwcvAN+3JZUkbLFg3Twdi
LJrsxXgcbtBY0kLgBFHhfS64Kpo7o8v4qmsJlv0a1T8hbV13HJHzMMRpNVJ6LEUc5AsmnoT/Uocd
yHXtZFu+Egh1PuBRmC+SzkSld8fn+ch0BlDa/ca4gQUZSZkKh9LGh1+uwsdcItNe/OonqaM/CBuj
tDXqUUxOrKQZmiH7Si/88L+H9PwLNx7KMWCCHl/QbIBhCuQxeuK1LCk+TAypUsCugodVHgUmzZZT
Or1w1ORjltlazJEGw90Recvfk+SlKAw1kdfClRI6rPb9R8eQs2MITXQg0krRTAhWhut6k6CcR+nE
ZiBDn1w6gVmdDEBp2IEl8up/JZi8p2t1u4JaMvBKby/Qy5aFY+sSbZJcPE4POPBcZecAnMh+x3mW
1m39gED5ym+/OtEAbEwkCXzq+DrZYKnAsYzC+23a4ThkkS0JC5ny+4pEW+fXWxu+ZAvs/asQQWKq
ovx1olzp8USS0ex2o4r6E02ACHB7H6ODkwXVSLw/P1rR1Zp9WXMtSej114LaYGca55XdI30GFBbo
A9gFVArEUoimTA8QLseLO9q/+n2BLFYqQUAjN4YolNGoH3xWvPOcNnox4H5b00Qj8CjJ0lpEcBW3
2/lL87ABKKXg0Evnv8Vz2gM7W+nUSqk8L9wSn1T1GIurvBUy1mvbChprfvstGpmVeEzAF55ac5FY
4t7NesTdpVHzzd1xlWyfR4dxZepUx5zmQNckn6SlcbE0JSke2I+suo+A8KTsachi7yyRkCra/cFl
wkoSQiJJ8lkP/hwIypUvFpgIXqJmyINmDnyyVwjf+liicu24v0G/Zw8u0kTUbYgoW6hdpxm6gsPW
jI/gSz7f3fAPC0BQfJGHUHd6QpqzX6RQ8BuiyAoRZHtimPBUE3hKScpTmWvL9RDOdMil4N51W/02
VT9PN3MkMuctd5hHPVyP41X2CTQCsHLEEsKD9W7BmTzHIewtqy/5GL4zxd1zKGE8R/NXXYqPyC2e
mt7M2KqFC3Au98Wn0nRlUXmbXRqLxMDByJV9Rwd0ZEVFffLzbHbz4Hj52QU9+KIB07RpUtUUNG0t
m/Ct9IOs4lXExSzAk3hoVXLckv9IrJUm7CimaK51FKZvLaY+OzjwGMOimPDVYSIjUOy9XWJDshE/
lQxQxEHGiIT89F1WAr6RS55Nnjt5llax6uiHmdXaAJWIiFZ2fvf3RZCOLBXH/h+PraaJ4GnewASL
+/D9/eOAR+Q/ENu5VtLhIz+uI7KL9ufkBuePHyrScH6EL1qFC7a2tGZ2CYyxG9bBnDjcITPf2BeZ
tstTq/GqS83pJndJrrQdpduWc51L7DAqUazowVsMMFDD9PuAIygU/T8ZShk8c63tpYl8et+IL7ep
B3aPyHiDn38ayAyB4RVND+xsiSMZiDXNg6N3T++0zOl+HpsPQouh4ZolvBpCkyOZVvsUdrR8upZf
muuxlFacZY5qsJPPV1liEMp9SBz6IU7SvmEbRWSaG2HL9YqnCaiGmRjZjWtKbt481Q3tCJDsDVM2
hSq3E2ky/vWWQx2teSQNNsHPHGaHeuMjdY5rgmL/gcq3zPkZoNpoBbNkBabsfvIuHxsBnD5FlUcz
ggHyVTXS3/dBC1MMGo+k6KrPm+EsZ1CqrHzUVqVdI2ga2ZzedSy3POfEIqLdesKvMvgtX4H17vq7
ursvN3DZNAwdofLWldwP1PR2gYoRazsIgebptQUDggdMo3QOIYDbw68pQmhvhVrJM/DyPysd7FX5
Tj36UJkDq0Fy7bxF4UyR1tU6A68XewIakty8FNj5E4nr1rbpG5Dq9hHqSw/RCDCl9XIAg3ymjC/1
6E5kHKPpWD0jJVudwrWdwticIwfb7pPjrolldYUrM4aQb8GHy44JraKRwDb/Y4J9AdYdBTPmfhGT
6JHv+DbHM2GoLOE9GeiQDlvOXTLXnKYe53U2KKUPULE1ESLJa6z1Sl9prtGNf71cXbGu3nAyGSfx
ae32tZY9TETUX/Y8ZSfUOdmJfYKmAgdQEBWJSXFrHwwBX/wAFi05aMWZAuFGXsgw1fUJ0Iobeszx
2/jBw3nXJCJUiqR4M8xg/wSHPK823Q7mObxopBj/3m60m+9je43tCyhTvRp+jNrRuzohGM0G931H
qZsupU35yPgXi30q5g3C/dW4MqGFWauJ4np/OduDBIR/783KrWui/EW3hIZuyWOJO884R+GEafbg
mk6dHTVSyarcaW0cCb55D0RIY4rSTFUvYkMT6xq80o3i5hSByOl5GGVJEtKunSRvhk2VWvgdlbTA
DpWv4XAA8RasVMMuGCpRG6mQ7jZ+UOF1E/UyOmLl6ru5R6eH5jIowGW5zeS3vZe1jsN3h89+aD95
rizQD5QdN3lAeps8BUcUa24sOqeuJuNEH9pGPCN7ukuEO/rg+uvblOMmfWcrYwMXDrKoJy2C3JPR
zjOYsEhEeyJrZpffkmo2uCOCwy/Cn9+nQp/u8iZ/mBSPdqGx/wX2DV9FVIh9g6lqaVhhiwwt22BX
7uV3yQpmLEmT4OT/srr8a3J/pU3FgQcMYwa1h9449RbpEYS1nOGhV7OMuZnvjr/DW21fCuYhhEFT
34WWPkqgPUkWyFP2ZbtdQ758vHqWi+gF8MD6MYFW2ICK2yyDwGuC3d4WNfFfJ8ldZJf/+6A8ttYU
qMXhpuUiORWF5lL/2mKXVp64iTFNSxOKymRMZHe9dEvU9+PJkBfQnHy7dtrlkbvRScWoGml0wGCk
lNw9WCPcA7ddBzdlG3Ab9eLb1aMOUP9dQWnUsDaWDZXE02UfUgIqlbbnwzW7Z63zl3CtJ/EAjQcq
TqCnmzp6SrTTPDiaR9vdZgoEC44B1ddN88XmLe4mZ1ZyMPqHufrFOxmgOmAeOe719h2viCptfu8q
4m3Y10VUZUbFtmR5u6JxvSaOC7wqDL6fky+ubgcdfi/gHcLzjDBUC+4iZDxMfVVghVmf9ES/5qHj
7v2+vaBAPReVk/DQjNJVqUptnetHsRZ1C+DjkhJS7Hgl6yNN3T2ZJFmBRvZ3Yh/HzWkOTSomMVXw
EHdnt9kJCIrGAfoB1DAasNrAlM1yDgceZw4ehityzad71OTBKd/k/dzZghC1SjvWZ6zAHcnJNLhQ
gNYLmFQASHCyEP9e51rosj92vzyU6sOiGcbJ2XmDZ7VczY1vDEffC+ZZvQOAkMAberFTER3dnOv8
LVPO/IolXnM21HKkiVLdP+76HzxQtpSseRmHebWq1h59giuVTu+X2s9XlYM27j9DZISo24qUGrt2
A4ljdDy6WF8eRS7tvsaXy8AFweqbXIDLBaq6ht2BPYyhpwSZiaJ7Q9UTf6Prq+n7/20h04KTJBWA
fZTGqPfI/y4EI4Aj2jhT26QceLsCdAv3b3qJ7gbfROuyh7chv7Vzr9OXVoqUDZpp9aehXmrr25hR
R/D1mf1XnnuGiENwyD4c5AZc5X4yPzSzKOdEuNJUCBKSaerDmpqq6WZPIgU2hkeCm4SgMSg4YPxr
IgWENrrSucrgJFHzqZTYqTeVCBRSLBd0jy9avhsLw7YgAs/eWag9L2OD5GOmi8y4/RWTqp9BK8KR
sixezCG/nmd460ZXUjQng1dXumtB+Ch0zHr4gZ/pwe7x+TzXvsyJHmX5u/duKzfkAtXAJJ2NWFnA
eDlpqM01BKBXcNV7+oQ3Q4Z48lBTvK3CeYIKGdi2AOwfu3c6XlyV1cuJ8YAr8pNAWIgBxEM+O9q8
CUhb78OaYdd1ohudOV02W+ltonVwHxwUZqruQXfE47ODEX8MTE8ox/uWlnq6ZXIlMJvRJSnax2w/
EeKIlBVXXqDjqlUmvFMUg843mVFzrbnLKfWtlB/sfwdMVH3TCboEGWYfc6Z9DZbtnZHJnFL9kF1B
a/PM+x85FrrhNS44ZQsOvX5FZbPTgo3Q8F44yUy6/AD6nK52XoZpniJgCpWxUzMHOdtM4YkSX2ec
ZXYl2fVK9i/rUOlJ5xca+B06dl7tpes+t6smGThRCbdtmDgT+vqLc0/sY8acju2QiKcy1KTFxj48
N/gEKFZnyyBhMeRUYWoGFfOmjlXBY/cZRbYpUGKz7BV3tGffFDaItny1B3S0Fpqtm1hzlLoLzCTA
Gn7n+Q0NFdq4nqv7IzyqSsbKi2Ml9X88uV8M+NI2+PjKjqTLDCZilkFgdm+e3I2cWj82JwQXdg0/
ZeS3jCXED4OV/ts80YIg4vCXwGDVxDbiVs1IHVS+w+onSb+WhGx+1GR0zFUVCQuqgR69rL8aGGbH
dcrnTvo074lOsxdVm/QMH8nIv2m/6N7fcHffUbQWPeVY9mg2pgEysiAfsmjSzKa7Ay3MEqM9CwUh
J5cBnY/1pvDpX1dCHdFyL6nSdmVAeKFItkreEPi/0xBOZEMbbgvnBTX61Q7KyNqFH3oHAft7WH5+
BD6BiDShvW068H5cRunjiN9Q/K6VdZ0ghZV8UDNHge+Y4HxBhRxDCrpPTuzbWNmbeDtKGmRc0k7Z
G2ubRBSZNxiHwgNgDPK035HPIBr34h8eCJE7QwEJMTbVVa5JJLjlHkOT5kk+SpIulz39GNBCSrQz
BetC48OWuf7SNkyb03VPIX4Iz1WFCF6MG6Q/jZeO4ZD4OxvVhG1f1wBu/TxxMdCL6SY5CLvFtt9/
ObUMhe8CUEaxFPM44VsTWvNNZ9Q6RxO1nMQ1m/QXa987PfnijtbzWjyn5ecsHVODHokfg13NTbvz
Aigja/Lj3TI2LqPefuxc7d51puwsM12QH88FL5sCTQXIcylG16mGHsbMndBSKmsWNIa6BMAaZvJt
KEZjczp1hmk3ikUJzUfEqaYSbTh3YonkWVyOkGh6Pq9X8NU7GyZ4Oj/n18gitIfKLtnCU8Vtki7Y
/kf2j8Izzb2AJEE3O1xpwEOqizTzDH1gq2P9oFYB2hY99P4mMF/ZmjK5k0ryhotm0YMdforBIrK7
WTM7j7xDpvz3+XJT6B8iSL6fxvIV7LUtCO2PLsPixnwHzMpWawpBL6IgB8HT7GiPnh8b5UZk4nbV
6FVU7j7JiOFYdevcsw08PVDzFbTaSREoKud+xl+WQK3bB9NgB17COC1vd2GrWbp6xEv8/vU6YBBi
3nmi76uyLdZQvlzEpMxm6pO3O9oXhSeJs/U1NrCFJovKy1pcSfGU7wCuk1VCBKOq7a7dveXpoQai
XnAhyH+CMdicyOr0OmiqHA2Wp7CLMC0PAfV2tWXzeiuuzpUQG9Ij4jEZFGKXCHt7Lv9ESvLOg4Mf
Ss9bnVJ2073OMBYJ8EfgaRKwtcbr1atHo8/Pc9zSoDLXb7tF0vX7+AZmf7oIgrxKKbQ+xQ+psPFI
kRDoA8UMPdZll0F3W1gW8r01TbI3yCqVQnh+xFzSg8rwW4OsQBBMc0mXm6dEn/3eRVWNjB3axt1y
7fTmZO+9xKhuLOQc99RTdLZkBDgGT9C7lDI0ck0O92eCRkRthppr+GVlxcNjD7BtwEX7SnuqC4A7
3UD1Ook5toIf2zP3pRVuS6l4j1cDBObYrAMfQHLnrrSU28Zjv3xobnu6nZ5DtXWza+umD5CGHt0z
68F4TU12DONW68AJK0UozHCShyZWKnDgargc+v+LVTdRaKeluKJZLCCmyAwfkJYJ1ztg7RFaEWwY
bouHQbYfxnIEwOWQ17ZCG+hAEa9Nd1+doPmsgszUMUiGKXJlC9D0/E9xA6mntqGOFey1oWF5bHzw
GcibMemJ7yHxgEFbF3eMxfoaPKHDSHjiIQu8SPnzTyZSlBPS54Yt1y96PYpKJkGCIqh1GL+GPcZq
M0r1kaNUXD52SU5F7vVhiwL6MMcviK/1G80ORouqIVGmsD2abgNvYmlQDjKZP6Ig/mmzWFp1VH1d
+U7ActrAAcYiZu6iZFEcyhB01DmatP6dcY46ywu6QoowTEcvwwSRUyEDEAu1iQZHwRkzncwS9y57
zn2v1w4vgHVfYmdcHsWqL/63FC8RmEZRX99eS6Mz2RM8TVsvmoxNXhH3KFobW/zUY6jFDuDXGAXK
s5RSYBlcOXxnnazkhNMsfpFRs7YjwaY7WF9f27hh6Oj33fruQVvJ63HN7Za9kwsSSFLOFhaliQSU
QsASB2sV1C+Bg22ySgezqvkv4DLPDQUzKaz/e6nuqgUIAgYu2ek/+wU1qNtPUKBxlbPqsE6pVdiN
XwifMd04snQpu+IgDoScfRoAhSa1UeKApNJuEDx/BUgj8sqPWnmn6l3MfYFyJFpJniKlH2l0bKRq
3niov9GNP00QabHR/URnkRrhZwpaVz7N7MDh5nGk5K1InCo05aqfnRChH46aJ1yyP/uXNTJlkMz2
6Lz9pMJTU6193chmc8MAsLGkL3+X0JFiYDSfd/5LPqyu9OcxIZcBudy3dTNhmGjBHEha5k6RplJz
JGVehv44gGq6HTCb+/g6WHoPw9wkfWsfhy30e5GBGjVIbmPq9vQbKhv8GFlk/WIMIs5aCAoiYG8s
duza9EHwSoW+196aKkXkImyCaCZSYSnfxq8mx43E1YN0vmUam0FME22pSC6KD3NPgNyZgInxwqk9
cz/pA7ncMZKKOJaLFxs6FdXY/V2nWp0MITU4hxfx7+M+dPaZ4UuxpPb5+oGrtwcYZYlg6Z6jQebg
H6bhHBZvh9YS26NsnmM6/4j7tazzsk4YhDCVxuKPHKQkBCnd/8EDp6eycsaMp7ymLxF1u2Zu+geu
jYfz4V22jHVCnplk25TO4Joq2deoloc2snTHmX3YqRgmZ5xV2clkUVn67f7fQu9UIXzxR6Ff9gL8
5qRZiBiv2s+k0ZbHNk+Hc+3f7mX45bRZY9eaJaLZg7jxjnvkSly+wspxL/jeP+cG7BHVYshOulfz
SclsmBil46xF1YT+T9rZs1hXQ5flkIqiIXWCYuD54bCF2LtKlFgwvnhaC8NgTGslWXZ3zbUyx0kE
MaLRDOlSg+1Gs33XgOLo7fcAyP+n6m8/t1J+nzBcu8Dm/kU1tFlBZnqm6/zy3bvBOUIXaxDGKixy
G0O8okynf/38wcZHhRV/frIlYgBHNYjZmFtS2ulaUT632WT+C+5qaGm+NCvdajQ+4amS/Nj5WEsE
fpEIVSQ2tz59rhaKOLoIyzfB759m4JFKexsd/95pQlh6kDqnQjpu06Y+HzyQuvUJFed1wYMV3qw7
YYOyRpHDXm//3lxlp9HUiZGPjAPR9U4h/D4PyCULFoysnmDVfcMK9M6enJqwiOfsucwGIb4urAgh
ygXyjPvDIa+P+axZICD1T9sbI6pV56LxbQNPW50TrQmDj9t+yVxeqzdov5m0YTJpPLmLM43PTgAF
1ygBM5t6tGjqwjQ8yw00u+C7iigRK4mYINU3sorZRZ0Qe6CQ+yo5yaZUh1pTa00XBVt5wxDLSXje
7FB5YU8yzh6J6W4DzY4CTlISpMgfmyja5TEGu1FLHmODyIxD5kLwCylob8lMI354dqnw9L1gp3ao
92MThL7Mye4CmX5ErB18bu9sTG6YpcfzVKIhbmjyYCqNfAUN+f58ld0I/q81cwE5/66bxHxUjwk9
/wYdIbLfZOl+2xIvrCHlVMF3RCdOlV1CO5dh1vLVEzjc9X+NOq/O8QXjWWOZXI/GttRojH1giIl8
2xWbGQC0nBfR7BhoAlmyL3vQNZsuiTi/R3EqtI+U+H512I7c3kjTkKAkdcV4qRHvm0SXxgS7xtVP
0bn0G80vVUeoXA+64LwyHkO2vwx1yeBFubgyP7PRu97YWnOyj2v8wAHD5pE1Zngkp6Dey1gbVLAe
BdjSfL1UoLXVl9tsz9kzJ0JidT9N5nohY/wZaSc6Anv1ehyepP/PGG29aVxfa2NgQFi4Yc+nY8+1
17Gh16thz7OKOEngA2xlCdnndUC8UDMUVvbfytTOYFz0X6N5Jykh2qdY0GTwkkSpGLjjXDCkVtPG
bN6H6thMxFyHzkRSd5dkDfIK1ikpuf5sFwsJ3jstFCiKYDLuLfChjXQWUF/bRLE65+GGBDh2lynq
abw/g5sA+hNmu6P5QuFfo/5kiS9cMc1rhMR16RF/M6SiTAymO/ZOdg2hFghrXC4zvRXVIcDlHvh/
3mBLZm0eD9Ift9IBPsVF1sHA8uS2Q1o+AA1gMUJidKUphc+0rI2O/tjRfKysHe3mcYZ8MrJJQKQo
M1B2+ywDkGGqs7UYR4GflY/wmeJfuZ4QlMoaporc6nDeel3Jmw34f7fcOVoJ3iXPe/lkoiAiiNy6
p31YGiPYXRCjm9k/6dXnBxn7xf+oh0mAwHo5MAoA7r7BEpfbbKOwb4UCzTXC3stftJBYk8jUJx6U
9d7NoEeV8fzOSD+1r1awF4Q1TRmjf+l52usVtGR0yAppU01qjkHEn65JTKZzLHK9mJNi7uagPXA9
dOS+ceoRDrOiVpMLGHPgn9gX9Dydx7L0Sv5xRP//4AIs8YxGFFW5GM0kDPnURD+wJUw/0W8jvvgF
N6Q5qqI3iWnMErxoKjK+taesJgfMt54lr69Ax/ttWzrRKrukwnt8jp+hx/10n/GCatY9vO3C4RHy
dMtsVb7m+vyuMWFNTLjhQFyjA7PY1XqVto3EOSHrJYjtEvlwCRsfZpp6plEGJGsp/WFYUeYoBgxJ
hlu6fiwYVCQLpdi5ELikt3rYniBP3mF2tl3EoerXSutFqyoSWSduNz9WQD6Zklm+jKMl6vpFHLdG
H8d6vZdwNQQm8te4fRmCA/2R3Iz0RsY/WCFgORasu2Pb0GiQ7T1AnwF4BmCrA5XWQxxl0HwZBWrT
8u+6HwDSvWKv22wJUjY4X+mLySP3DI44aHe8+a6EagJSWMva5Qtmw3VlS/M+4VQS/RmFNfMyVOrp
vnBZCGZiMyX528//bmLkFgdCHU01sSHOSGAzirGgGWfA2XxS9iKnePI9PBB+ZT9StoMQLMZ3mvZo
PMO3o/UyvyjMYWqBcvJ2P/tJPdIACp/GtdRuSsZz4SJ/NMBwwK4yQynJWkppxDRNQjzdNj8B6azI
NR2y2ZsKjzZYK9J86p70Ib7qN1yinFA5HF3LAxO7PaUTjeRLLzPXqshk1/EBij/kvOHNVNaNMoyf
2osaOlByFmXCK04NnqbfauG3Hs0eDFeCbgo5mXowleWOOE8PrIYx8RLSttgetZjxvliQQ8ncwKZS
EPDL4iW6Rkrd7tf449Ko1GUOnh9szknnyXS4wmajCHAgz8aEel2lbKQYPJdDXqs+V9GNyNGQKw2/
QoobQfKO6aNb0GkBQEir3dSaCDXBJ5ByyIbOZYGY+yJx3Z681tnTz17r+Paal9u7XNzRuzK5Ao0i
IpUPDhR+3y+CL/1jq0BrBsOiys0MHZLOdd0Gi6Xpj1OOG2aNxFB4nvi5RiELDGr/HbyCvoMVKev3
/3zsaWr4ZRBl311V2692GePgi0Kzt7I02+CYZx+wloHatp5kebENSku6JYsGsM0EtYHmN2CGfZaZ
RZXOeCO489QI0+UulGHyIMkqplNOL0X9ZUrDyUzE41356H26FvfJpm40wONXh0H0KPqJYBPYBykc
x7uD5XDw4SOTr2RXH5YUjGGf+438YgacbgZRVUGDVKYzYZJCaMh5as5XjP+fwA1N4ly4rf70DuoM
IY3YLuyeA/gOGgIRlVf05a/Jh7ynMPBtJDIFlFvOPY2BYleBSx2oNzTXrV8v0jbY5uO6aWypzo9P
GMNS/2IVt9CkA5Jh7rRkv+yoohGrS9Kig11DCDanX3YQ/oXr7jNBXJjugITrMXYwtSEdEVvASvWL
KsgnV46oTH7NaiNEGgnX6AWhfeKXEppHlyStaF/7Zk7YsZWb0ynQnni2vdnqNj4q2kgj7OsdqZhN
e9zoy4Mdp8fBVrHtVscNdbz8R2DZAqHzZ4sfXjbj1oT2dnoe4r20xfxzOKoci1hxehq0Lo5djCnI
2Cy+Qp2yBj8yOiM250zs07PlbMXw7H0W/0nuXvLKuGlDpoKPQXD5IIJSqAqeP/gl/SFQTfb+lreM
wOZPkW18n/Y7TcglPiUo7TIFf9SKRqON/o8cakn3WSTakEq8Ge4euRJNgBVPpgwj5KheRotbYitX
TBHF8mMENHQnTCr9gil+dwfyMIDrnkNjkvIzYmh7XCfx22nj6QHxBJ9Nj7LEofKZMkY5W3zPWBB3
X3IWPW8CItERc4cCmVRGQzRNjxIl+vPgdx/Tx5qi6H8+g0lwsQmRjbXwnjLlI0+h+mWRh07r5XSo
H5vGaU8PE4JJSP7BF4Lezy+O1C/XcqC83MBQ6lZQ63paG8SZeT4u4kNIXgZqai3FMQZvGW4WYUsF
fc8d+ZV3pkfy6CAvwKeL7u8pJH8aJaGqcscqeGmIxdMCZadl2FLA9M63MxuslOJDH4Mx68M/+dLj
y8YPJfbMgCEuAf2yL/0dV3DOJ+FbkMusWxyp84Tik/wQuz43sU7xLF93ofWCDZh9FS3QBobEsRTH
CUrphpO8zrBlbx4VM785C1lipjlg80HtraMqTiON/UJY7FsVgkPe4ANa/2J0M1EJ8UO0c/wptC2n
iLsp+uaigxeG7VKSAbJbVpxVViet1DK4binwIW9gJQsfyXkId49xorwWHL/LKq9/QVyZAQfBzKZi
fp3MUb34EdFUmmo2ehNnyp3d6/CdGou4bpnCt4UlEbW8Eae2jiXL8LubITukHNcbL2zQGaWcEIbb
a579E3HXEbfF2i0apUAMX5KDCPRe2z5USVhoBd2XYKN1suNhlge8RaQ2+ko/mB4Bs1lrqWKrbtQN
8uJI3cbhyCGKlb4z0iNZ1qFZxKwLuCW4rt+d7z+NcWtq56q80LGb2DHYVQ8IB4cZBy7/HLbZEse/
4xrxJ8gU5Zo6xFUE8sKmg2hFPTsGbAv23vWqx14ybBDI8idMUAI/2J0vLaifzE7d8XSMTsvPcRkw
XX5l/a5ADLPsSgeYPsxBYFxatoCc7uWRt1e++9Sre/5ignsQAR3BiYi6JaVnCfbP4lnQNBt4s8zP
rjlmtLOM/ztwx5CoaIhM5JgZSKQ+R+fMW3VqEojE+C+KfXlkh1/xknnnppdtjnPF7wAMeRIKTCeM
sUQQJ/QNAUDtW7S8RjZfRZZ7ThFJMFiJFALygs944CjyVvSZJTKFy/1lfxP69THNbr5o5CY6fL1V
RYFsk0TXL87KKjBnGQIcfZnCZCFZGRtpE28RgjDu9sgORgG/kJp2Cbl6WlZcyDBSB5KJl5+LqMD6
AEYK45455UlF6LiRo7d+onqkkv/tkmgpz1zBTq10g62AkpRfAR+Ajone68fv7VWtlWax7iD1TI9s
JUfyN3u49PxoUKSsXBfu8uPjJckUryKXS96LgXDjCfmFEKoMfR8MEsp1gbQRp2EA5dDsMCcSSd7X
9hmRK7jM+KwqMvahAwpLndBlWDyaGsScc4xp//KVlhkjEXBEB22FdJz2ieDMV3Zu5X5LDlrAWmHK
a06pBeMBVwsLokZuoH26qskJtSYPwhHJ6KGsS/eJjpBGb28vPZRiV192mUFsGUYqw0MHS+Ihhur+
ZPZGJFgt5ue2hTw7HnRQnDjUZgDqVIFY48hB2cKbcH2xQ9b2x7M7v3aawK6chsDciVwKhijLbGhW
aI8Fmc6gb1lTuiOnDmCqOWm6xKc1Zcgi3MNJoGHJ94J4fto8KQu58ha1BgQcaDZe/7i/NmgeGhSB
1C/4jhy84shD1H87+ZjG8DY4zS5VR5+9Falkr1O/GY5nMZF8JPcmxt3sGKjE55+aWiQL01fWl9Ah
0A5Num5hwr3BOFmUB8FgoUD9XHq8BWopjY0I5BPW8HvGKwGA+pGEQrreHU9je2y8GqyE1BLSnE7b
u+Dyk+HMoliLeIkUcYMx66K7z46hlXbpjGgrRt9OAYQIFpKmAMVgfpWDQ7pECxjks5Hbjd7oTm/p
XkmYsoTJ7cty4ERxaahJIm9G920OlZqQdwouK9f/6x3bGdBEcCNVnQdBCF1gz/keFBfT2FMWUIak
WHDvY03ZdjiuiFqSOSMz4RyYlvNirIYYx3nHucjvMwQ4r79MxlN9jv1pKsHpFSPzt1lwzxUNYevH
OXYElglQUDsdn8ZGeMlOfA+gdDJf1faZIDV7SziVgHttkKJ1pLrxPRIodMpsNTZvk67okm9XIdBN
de40/hvkQkhtrwJLpoZV8VQH7zqqfqHKv7EfX7oBBp7Ot9CkjTQqKjjRvs6m0qWyBhqTWfjFIdF7
4bRAcPb7vjMMrUDEM0LemG/iV2KuZVEAGSjFmg2wvgmSrYA18TkfifmTO2Yu1Q3A8akXIzsmw006
ZK2tzYH7dWf/SQmBurjiK/aWaWtLN/s1AQJdZQep1t+flogTTzz8wBMphK9mYGhVrrHCW3O+IBgu
YbgLcrnhY+r4RwbGGDI9gMqgNZ5TAagM5j87S6lskJb72OPTztHSSUBT7L8hHW7Qa+10nNzyba9v
IS6GRLfxpRTmKoggUaR+600qs7SDh5JgoDn7Q0ouJ1P+ioWHi9uTPvbj7UzDtmCniO8Ro1js++Ve
7RQNKcg/aKmJV+mKmxZfEyBMeQFXKMlyj42e9AWQf4hF3/gvwkBsOSen8A3zm9m8lfkGP2dAArLq
IRsSAbrpRATbz1+UY8xsScvBdu70yW8yGVv72HFmus0Yn+cjRdb0zE8eUZsi/STcQVWx89CtRiNN
qWuiiy7p3oD9dfqMiyfGZtrwwxFuZUoXE+yCrFjaVxnSNIwNXTAK5dFtQ+I2Et0098JkU/J2iKXF
zJ3FpKmrqWipMjRrJ/6hqfLiZweGLMEcwuoOHf4GthI5X4TdPyzetVQR3dL5OVFwuPmqltISPRvP
2gYU0KE+22S3ZIwsUjuelV7u2v6odwfNRuEVa2+JR55dqnl4ncWPpJliXR+KU8q7wOILlkIDE3o6
sqYfR7sp/4vg73YBdsOXRcVQVE72Wlx2JFgIY2xMjo0TFYikz4wZCIVxrkML5jGzgSWDRAfPIZ7g
zSrFacPzTlddYyz/TmOrnBdvGlSAPBc1Jga59/e3kRtoACFJbzuyGzBm1Ep31dnJnnHHTJnxyYx7
y3r71uYTxtLrUK2+CpJFD5fTRjW54YhjWGSxa01UvbLyaLObLJNakyK0Dx0ta3gr8RJ7/9Cw/9bG
2KETFbe1DSVkbPdf1erq27WQdYll4cjOSXGSnCIbauAbcWW/KV/l9mremdHQIDmIduONLB/yBzAZ
9ptGV7TV8b2/V2ZsI6dGnSa7/H74v8F1aLh9+VL/RFBRSIxnYvibh7FBC2XEvKk1C1pBR/nXtBut
BUQtCfVxZKfp5QohUM8BvuhOE2rk8NWDLYUm4zrwic0MFg/mdB7SEPxS5s4p4juaFWmB8GGxuTIS
Td5shqPulR3J1kq0JP63xgRsIw6zTWrr/odOLU2DdFCsNn1tycqg6sz+qGlxq4X/jIGGVtlySM3H
apB2ZARfnqi73Bbaqy+nH9zgtVehkBlz+wTTV9OC7b/jiu0qdm01Nr7tif1yX2wOdAotnF28lop4
PPtR+pJ64PiqXDdtaHcUEqSMJweJ8d7I7FRd/ESMaG/cIuGJkG25iSxGF0FXFOOTJC62r6UwuY2K
ImVhsHb0qIJqHltZFWLh+3Ff0vKjM97ioVbxqYl+giZYizyWdxgSNr3WtudRSFb+LFovAvOaikOE
7NnIF8PU23C8QYJ8FfH98GEnd5vL0RSdQ3ldHHmLG2AbIqyovix/rL1YjWJbk2Ph13b+W6AVzN/j
KkUC/SDOCwv55lxA1T/JJpPHrYSvCMwuoCC6FkIz9FC6b7tzp0X6Jy62JR4oMSUvolPqELJO9Nju
SLywRrYAE2F2JeLBWpP3qRlCYX1qEGlkRiDNx/kJOEM53tT8/S+B+Tws0i1g614d6YodazL6V1ko
mQkRoIjkc6bfvKLJreVr+IlbCXNfzAFP8vCWIhBly5yuduAWSY8Xk17Ld0j6dIPVITsUOVkW+5LQ
3jAyhf8fnRrdr/nIdm5LOpqRydPF1oDswFAsOXkgD6OJMhloeMBh0VR0dJQ8MYhEv9JWdNdnCr3G
edApo9H/X2x/ad5TP3ObAiAvPvyhfFscaurRyVJpig5On8t9AHULxmKMOHyxtmU0OkseGJyitnHg
pYZYaGc/+2NXq7HZ8Ts3BVgyWBG8S3YnjZ+0Vdk1wiO8R7p47lPfz3cAUGRfHdyR8UJISPb1T0FD
ZgfaFt8oCIYLPYdvWHVudV7jOWRL/IPAPdZK6gMCDfKmB0iU3JBTK96RdzAgysY+EzmVDq2zg4qu
Rqf6lUDQv7dFtwuMZgIy0AXiccBHVQE5CwZrjyyK4yMDax6f6vqHQLPvbG5CDTpg1lm1DjouJpCs
OOpPknOqwFVf6VLi3W0mdqro/BKBCcytNIjkLSu3if7SJk8Ak8O6pfbkFO1Dbo5M+ftTwdZ52T6Q
w4mKxSmGZiWJ/PgXjXedwXHLYAMAzXqZjCZKa5vXQxp1CvBrpn5dE28FA1fMU4o4bSzcMNT4BJ2/
Jb/w0pss4nTJ0bzRO4bkLdTy1w0Bho6drsxTbk5ecz9IDiYnpEdHlS/ALjTOzj0G5roDROqCnLoL
SRXlrED+QVdWF25aTgeKQSkzXZruz5hGK0r0/5T/P3hjHm2zhxQn8O/vWSRoeS7O6YtPCQIIP8JM
Hmx3J6RyP4c77ei5vQ+byeUOtT1SJfr5C9O7efwgibXvAfwA6VFlmAIBMVakIQMNXc7TQSwR/nbY
TKkn5WOCNJ4FjhUxZmERa5Odl+vI0zuInh3zBLfTgLsuBSD0GoFHsPuRyS3W6GAWf2gOl00moTVp
24EgaIlwq45urZhLHnMbpK3JLgdR2R9+JdVL9qn2G2B8kCSnyhdirfS90DaWNjB/EqZoPQHOj1c9
o6rK6GDsGz9gDnH2mAMrhFhtFxu7Kn/yNGBst4OiWpYay83cJToyNiW4efnxozYVs4ndSLEIaXqE
zOIuMDF01k2zaVuBJwHIo8xQR6xTyRVYTgnxAw7wAxXZnv27MERRqsSAe4aDsh7IH+InmOf5bgF0
xD8HEVY6j8wiCg4DLsmP2HC70kiFQZDBsuWoYKwofY8gode+xQfbt8d6/IVoAPzzs/yX05V1Z4WC
LQAvZrbtjrOpl4HOIs/zV6318BQvVtGjGs/AK+h2nlSAUykPIoyJ/SqdhA1LpqCoV1e/zJz4KZ4z
y2dPLWT194SHMKnyJZmIgfCKuOgoItEvbIZ4piQgc8HHS6l3qXpicAmWjHB/FIOEw/7zRxkLKPto
jRFqDqRzDFrDcF19y+nz2KWG0FE8er/byqDjiTRvBVesKy+rdPW4+scwAVam0+k16YD9wyAfxMNx
rKio1/bd05I00Re8LOI59+XUI+I9p6xcvE7oPjU6/inK9R13VweYaHR6P/AFENyCtrXeMQZMPgri
PhsxG9KSZi36E7g2QUX7X3On6iZjpYTrDXlaj9QBlrDQq/KsGH+aCAQkpWKtK+MIufrMZqAVb8ve
hdujGbavxRaX0drti8EHRtzz9OOQq5qCN8Ed2XPfAJQwvjzE2BDeegmcfDwFD6NtAd2wBV1/MOuT
wgevLhGDi/6spCMi6pQh0fBrONCYLWnLjoufTNIKjjXD74ulkiFiZVEZ1BNi4YdJgiBvEsjYF6Aw
lzlBbhaLaXIJKWdkXOfDyOyKoon5HAVJY+uCWoy9eDLQv4FMfvZC2wosayssoTMT5z53kklnm9rI
nyrOPshdCO0jPP8qWhBuYaIHUYF421Et0+tY2v8nWVwhOfXhbJTHTazcEY9mitvIE0dav0FgKJrF
E44FkC0MeIiGQHxyrUyNQ3wX9lN/f5ivztFcxQkZfCoSIzRZoSJrRR3xe7v9dSod8ulg8FK/A/5m
OizyayLT2gUt4IdXBC+40sPZ1KVUllyoRD+NSMtJRnH0u+ZzhFfh9rxXDXqf7HIKTgbU6QyrcwDi
cgHNF3KnXoUD9YwKM5aHiT+6r/8en1C57m6Di85750gvA5sNj3Jg3w/voezK11YxUIh3wsZlAtDi
p0NXZAsp5C1Fe3waFF6Lq8dhS0ad0ctTkMEdpBwY+O+oZHXRUwCjjyLe0ualZgPodit+J7SsI9xm
24l6pVSqEiWeQsuEtrROaoBQ7+Yro6JezPXdUWAz4+v00mSavLbKWC7Ij1u5zrKiGae3tluNa2uN
bx1QMBjz9JQaFYfC+Jk/PtPaBP7XRa72aUUU+rqqGmV5sjdkNThwxDrpQ29tJ4edNf4MJuGNEy/F
H6iZB5eaHK20ojUGeKHWYb6vcx5SS7G2INekOiSh9mEEGOm8ywG4yGu/PV9PGLWez19M9C8cKon6
axcTEtrNyq2BWLH+qncICZNDcp0gLQqmz4luoSffjoSqqPxtCkVc+mxtjIx82MhAt0ZblgaYTDL3
Uwo1fkLhTIW7SyU+VoJku3Iz4t0Cus6E8LK+05VY4vk+PMcLBJo6OzFwztkQNFQO/G/kGQqZWxPM
oRKyBU5U8n/TaJGtY1/YMoMD4XHQmdU2Kqjje+8Nw3auVYtdP4W3CnCvdJof9sw4mEwVQHsJagTM
Yw2TRtkdsO1cvnlRm6DnRjgDP28nvnWbMfdrxLxnq33CHHUtW9NjfyBEhKW06bi9uh1aSBNJJlqY
QjEoZhhexWMxS83KIdb2+4+sZnGfo0OCEhXSwlJhqAtRIpcMoyjhz3rZNkqu1fGSBva2+zpl2hdi
XIqVUiqsFUhykCxOCoOloYPQuPM4hBhajiYcr91QSthJziWXzWWUQshgX4nRFBokEvWezAwFpXRc
zyNy8Y8n2TkzhUPC3Z2h1uCUQjBI08eWQ0gIpV/6qXdStL3TFES6EQs3ehFvP02ExEE5Jij/iYNP
f6MeuxEmWVNF/NB0pb3zRJAXQLbdlSM08Chwzy71R0OeQrWksuYCPt3XjZKCLXbsz9ZH9OSyAGS9
ojwFbOBHmpcOymsiUT7ls6df5O2dfCQQ3bgdVQKdw+PxU9KHonkWAEEHJoOA+bwjn1V/WmriMRnm
lHoMf+7h4tIEDLZO7Z0s8nzBZfPsOjRN/vtDL6wy85ud7h6PTLZ/93gPeD6M1GlA7+lVQuLDRahj
eVAhcFAADn1cNEL436+HNGPEpgKZyvGGxU2Ke2TN3XN/NvSyZZjxxZOQHbckmzxs/cwG7Xws4e3Q
lZnlulvYCyrG5nzAFtxUjsSBYPIdTvfO/h8kvbu3n0xI1U8MH3E6u90zcoLzNhJ/DQFVbmlK+pON
JqD8XxmBKCIDuUjj1vW2m4jJBKuOyGAzdbLhAwfbnizhwO+pCbcsr2qott2p1akHTCgObO3oHSB1
iDYhdpWnJ3kqWcOlJEwR2vde5QS8uPKYzZCeCsfbZctq0KElZy6U3xt/HcGnjrJ8KOydHVP51cak
j9S1zkk51to6ilPBzykxYZZFWIxE2f4fEviV6bgX0GzsPED5T1H2O1S3UmQW45Iliif0FqtPjjB8
Qum4Wj/FCeyzLYiKG5cqWBK4erKnMga6KxER3KQ/l18dasA84j/6FMMoH7zMT/UyHfMAfEf2tecA
edrLiPgBdyWxBF2T/D06DhFZPo7o2o8kofpQIkzH5zPd77h6IHTX+NFtIGD0q/7u9nHj/ewCed9M
EQ6ulY55QljSfd/XoVcdmdu4DIGj7Pr2NzJxtCYdFwvaIjfhP2WDfzJrsrbYRMaw+lhwj0SVciDr
6S7S6+0KqHxxG+vIQ2kTvswGqXJAfynO2EFSOOpcyuR5IQ0Q6be8MwMK2Nz/iUZdersP07ywGUBK
sMoNBrX5lqMGOmCFVoSAA4KxDOQuNDvwCCD9CyqHrJduKolcIOKmJb2+Yysj0OIcKXWiXmD7234d
QjjxxiuCk+TH+VAykx1Lrc6z0pC5qw2L4TniuohTljA4/f0yRoemUUHEOR+Lsrp/SlvpaqARkXQa
1BezY3zL73mMInoYlaQHh+o8PZq6zw1IGKfJw+ivgek8vIRmMYHygF5CYl4a58yhNwHTmWG1Z3ex
EVArbjeuLqM1nr1MUHOa1IlmsADViQD4hgdsjixtOKd6tB2na3wdEB9BSyYZZV8a8QW5Jg6dBKyl
/1dpzGkWz+CrevOkNgAuYfqaL4+iCYEEJtzpdAWXyU+RBuTu4u/yxARcb7jPNPrM/4UZcONOsZf3
nttNqiPxnmuYyzPDxl/epqETMEfkOrN9BAdHyXW4yFeyYnHRI+GT1FO9HWxi4u7S/4nx0Dv0g/UY
aOq9kCINymNunSgsO6wCyzL+xZg6zzZL/VzwNZthSEOHzkMe+HrqF3cOs1kYxR/XJ0wBVUnxHpe1
V3D+mjcV+ns4qH/iQSfuP8EJ3lICnLZNYx6XEzqUO9pgtw8gUTwHtwW8H8WMeuOlrFA5tFxDGSKw
e5/0E2U8sTyDiu2l7a6G1YSJWkBF7O8vjIK1hgYmWEkdxpHwVVbCuyTGHaJTsGpC3waJMlRHyzKW
RXwwEqKvKvmOEooPJI7LxIV2enfOR9LqOlOs0Llbj+bI4UP2ut0dO6zYP3P37cneYu/0oww9g6ZD
Q69Va6JJ/DripccYFdxQLjsXtDwRFiH5d6+9yqtiyK4sAN3HZ9k5K9bDq6MUy2bCMbpyVBVEqz89
YgYVEtbzBg9tNWcIH4nPu8B8Ed7Sv5E84OYcxEaoOXp9fTyqEncu6Sff1iI2xKItPBdiVsLeHZEu
w2Cd8bBvH12S+VPa6mynPN9yrTuEU/bd9Kb1XUdND5+TnBgEzmbCq/tvKCLasEP6XCCjfkj9m6TP
ewFsfEzHHknqrXj72LkOAQFw2QMscFfZT5l20JTq5YbAaEIxYPGFzEe3gMb1ZVkk4UBcV0g/cYs+
u0BewjUaKN4OXe7HT8DNmM5vM3V6ugwpsjP6q9vgxG0bArrfuO0MAvPjNEx0t0+8LRD50/BeP8Y4
veScwCjIx4LhI80CKlPwmbzrZyiySar2/Ty9Bhuaki9tkN0njyKAb3kMFATCam2oJukYgCydl1Qh
dtBOMlhMx3Ily5oQFINRuFJmYppDXxdCLJBVAZXD7t0rA82a7FRDilkcQvBKHt1MKke9CKGbhTrC
3V6HY899WEqnussMv1k82FtNF+LHzbAOVj09626OApKWmAqrw3L5ydgAitnZd34du7wYFG0xex/C
vETYG7p+H03dgV6oxVc1QVGwHs4t8AgqeClSrsuQV7fUkqOAp3X9o16udRtdVvSPB5x+zN7L8/49
TLAKJ2RHvF+HRugMMgKVh4UdrAMxhMCMRuCNsHS8yoj8aAuSp8UxemrqCakJVO+2RDbg6ZPKP8rp
C2IxTRRtFAW/URCzS8EVqL8wkxS6M3005K2c8piZRvSftLzl5TcMFVEAqJTXpo8CN3+hEgtZQAEA
tgTVgI/h5kurKhYP82AERuqtB4Pj6dNBi9UbFhHJL0kTMRC96E6o6EzNgXXmuBfv6ScH7v7HFRhH
2P4j6WL9eGN/J3siR4tF7M46d8cLc2zGAKGK2TDI/WrDDuF+8yyPAEOMC8LyozpnjIELMczbR07f
HesGLMdMHRWH4ZZ6xmTXQ5qzq7n1Mvrx9wFeyHW6o3Ukc1iO0D6Vv8+rqqzSl+tAjICYflZ+Mkg4
21Gs64Duc18Kiuq/fF/lrM/FQsQZesqd59jcYzI1E8cmbvDEtIZk2/pqmiA84C2ZPRKBWXs9srpJ
XKNbOYYRCqdeAb6cQF3qvofHvPJvJ/rbuYKnpDiA6wXQiciX6hfMBha1IiMqM/MQ/1jTS55VHGDH
Icsajedy2Fi1FPH8u925ej+wCG3TDdbA5ItHFFGV8ybZ3obyuTaJjy/7HZlSJ/AxdjPAMiM9CB3j
W/lqYgiQLZaURI++xfJU5c9NHAnYCGsXFDXPptbKOszQVDVIP493RRVPLBmS1kdA9cKVnozCoRfz
JSiRJ1WIEXBYugKgisIyaaF3Hr7Q5vf6xC6u0g24u8LumEXE8lRzVwAncIi10y1Z5I8EAWWFSMhE
FRSnsFXKyM1DkestCOqFvq5Mt64IHqgaGV7mDGczUA81lN5fj+9BCqCLmaI4GPOJMUISTbG9fG3+
lbHTteFK8PnL97y9J6m4mV/f9+4XvIw894/NGavMRWLBe9Jats16x1AhUHs1lmP/La0BR/D7l+UN
wQR8HpFnxBmQ7NkyDW5TyHPpEbPTusyGOVHrOQOad71uSC1u/ZfjmabP+/oc7XpoJEDdtqF204WW
RGluRVuOGkWzZ8QkQQ+OTVRy43w70i9/wStL5hOae3Vw+n1x5iDbTTAsQCQga1OOgaLWyTQ3y6iT
ANuFw5OB0vsDRnXFOiIXpuGjRF3nSH9GrtXcXSvZu3t6VYXBL3NUe517KlLVq7Nf0QGtklkAPGXm
fF5zpLW9OZPIAzXrJmczBqjO5U4GkAsQmYdz0+9mkZJ1/wIWI3Qo1eKR5TNreLRSJ5kCuyu/F0JY
1fr/nedoZwLenLC1LxusyorLGfblbQiMWj7Sqw/tVzRlJcZIoKi2a47uXDBkvWIOcS4I3enA1xr/
vdnMqNazctcu02WdaEdOZSsutfNsCDG5e6RwglwAKrZwWCYPxsU6XEho4UkMM2SNyI0BnxpGvELJ
UxYCok2EuUIBwZSej2nk/OBQeAQvplZeBfTte0jsY4kBL4vPl0JBUwo7mCjWDvKIPtWYEiq74KPM
o528MUD1eNkZtmyFjNApWy4m9RGME3Q8BesPil2O7WOVApYD44jzZZb2gEph3XAo5+zDghT5k/7I
8pR7aRz6XifNX6L6bNz8DcBYH8Zw0AonE+7hE0wUgTVILZ4Nlovh6FXdSkSqdcx3aZYYUg4pDIFk
JYU3LjGGAqDAKp5iBAb2DahJSzqeb9GSy80h/flQob7ue17HaBrpdwvVY6cOakzRh5e2+MpbR7Ro
I6CZHaX3CHwIhp4TKzSo1i9uWIE1ylAX2z/XaQByI8mhyYk380aZeTfbIeVWJXBITqnOvAUFw6zs
oj1eHJ/wv5+ult1Z1sMupXJ84tQBxI9wJrdhUJ1+TaZq9bUzDQR5y8W6feexwd1+tMBd1EAzA3lJ
gHSLxDG3TI7thGq3N1v4BZfj1M8cSpBjs5TJmmhJ8xJ+drvDYwNRhbZ/u+1o1wx9rySLrTya9/BG
zSuWeu2te09LE6MkuAQvwgQMWqX3385URwhJV7Biu+SD31ofqy6a7mksIRvKpEMrEo0aKMQkOOrN
LzjwPcBaA6UH1x7vCAVUrPbn8Ua5lY/vTjX8jFagZkuG9iqN95b5fwQo7aBmR/JNkp77hnCRKCiF
FCQEYuEkJVzzcPwyje1+aZwjZEydq8hIrW1qNzrH7X83vedSWpgOq0VFiEm4LmP/wYOb/tjErl8c
OelORtCd7ckakkfTWlq3reUNYdwqRG8aK1h70umdfl7hkK1Qi2VYr51gEOqIVw+q6i2sgSHyB7QK
UMvfMbVm/UqJdpeww+xzGKUKH2KxsOfbmrQEuLoxzoFNKSvbN8W4CHyxY3chbJld4Dhgyn7Gc0L8
IEHcidHm5XDbeQvaW4iPKBKBhCAmiFgawXVT8EbiRtgWuEQq/yEyDiealSU3uEr3k+5H8n0VwKzb
no24T2HM76QEumIK3foQ4EKvD/rn0bQUbAhmAb8CUxqbY3QUlgPY9cNjDnT+owIB8/achHrxsZuI
Zp75pNpWRnTTYyXxB3azKp36B9qB4JDxKiyqJLTyTPSAW+JYJ2MO0MF+eOctevTB9826rDoNVxVw
LAHuCsbr50UkX9EVLbDuiMbZEKMW735P2Jt7JGkitrk3UWFD2jAKiCF9sME8U8UtHj9RA/X+mAQF
mShH/DYpCvk5G5vlEoWxVowwcY3Kxs9oHT8fqDFD791+GZVO4yWP4+O5sf1cHS2Q5dJzBzRhjch8
ZYwoQNNOTP5ollzbiZD6arN8zfqI9GO5nDt/Vht3SBL+UfLohx7Va7krfoU3Zzp7fDVh8KkXWYPo
PlyENb4p/bTI9YzqUznypbdMHwFnBYpgobSLOsRqPYChJP4gJGpD0SwXbN3f1VIbzaXiJsNJVi39
e2KNtB/9mnAqc+BoU0d2G07xkMD+yoT1BxnHOdO/o5SQFeRSYMXN4DRkdxaFh5Z9wXhMEHW1rhiT
dfVL/eUzgNzTRO4clZk4z5ai+3f+eYXn0RdLHh9F1HQJgD7CqtPMA1rAUuocIKas5IoBySDN7oct
QRYms5n1N6JbPoPWQSHVSew6kRHY30u9s7A2CXOvLJyyqVxVBN4himG8psqdeYDXMp759xubwAxR
Bb+5y0BOFql0VxPrlPcSAwtLAgF5c2rf5KksySspnqNqW2GEq4E72Ab1NqqkTsPgAX1fTR56ADHT
pHJ2IkbINj9ojAJuIPuXMoukPHKzjzteP5gbuFA2awgchTtcVENSyzEtcZ4CEZD+dYmi0UjqZftI
h+4g6tpwGaNUKZ56pjmO4anVnuTyEe/ohWoqc2X8O40uMNGz3Y1LCow7NzsQ3jtCI8z8ETv6WHHg
viK4k0BQNnFGhkL90QYYbA2eTELHi06KOPXshCrlO3jvVhhd05yA/9whmRnlIdUBvsqZ9t2PJEG6
CLpgkE/lqq2q+2cR24NU7hh0AaS7zVDf0WR2lbgzWGy7e5iEy8VRi5fDKpIB5gTGYgMiGnD6X6S8
tErg2kcVGXDKWmV5f1VPYNNxj1zk9ez1Up+It8p33s2MQg8vzsRNgWThMp3GaSR5X5I0j7/ZggNL
eO33hg2ZVVW+u979VNtNw9qfVJSED2NLrVIclPL+w5wvXalsZOtMqZnf2dUFEvcDTxdhzSRAciQo
82qE5MhHN1IgUioFuxlhkZrF8Gp4Ro5/S5jzRXYcmXOLKykEOIrsY+83sl5GuMg/TG0RDUIdIwAj
nfXVWjn1E3zrHkARqsgOfF1gw8h9xgmyeFWI8+2Wm6iV95a6+5kAgMDqWmbNLfkYZhZ2znbJlf5p
WMzuT8yv6Ok1LbobmqS1su21uo7tMzuuqI52q0I1wWJrrr0T4tJADnPtoZo8Q3wbs7ZTOeJhBoH/
w+q5ip5cHSOFVrDsHBbS5XT92yCAEnLuYW6CF6QOfNpRV7y3nuXNBlUN/Z3EPBt4MZIEkywv8ogY
w0FcqhoPcnh286Ndlll6/g7t/41xGra/DnhEZD/VDbnQY2Kj7k8pTmzUsilAcbptgXz2lhoXcSTF
wiD8azLbTBEQRCB8Iwc3mJA6yXT9LoOHc8lPs/2JqK1PY8yGgKDkVkAAdle7wjhTovktP0yhZQsH
Npuh1mYGwTEw6Y5l0hBAyxd+prCI4NlcEgv7DnuIvBsxyVwCoPEhwwBjyVJoPqZ0w+ma9ZBuoJ2N
LnZoqoikdrF5gJIr9lYp8QENl/iVE2N+bbvsmGw3nfsh5jMI9zceRTPnSzZ90VuNPLh0QD8SJIM3
9yQgLAFCV7bsspk1X0Hlb74UsfYu07cRw7NimpzxRIvGUcYkEVvwnoTPZOfEJ87PviENMKqIivZY
K+xAqlKOAFRWyrSEZnyYUrRf3Vrpe/RrGREayvXdRIpnqr9c8X7jPiDgw++47tzK1fspIHo2wzL6
wzbD+zNz5q6vEQ9TfOdYD7t6vukaYnp41WLKVe/Y79pkq0sCvyoc4uEB/oy4/7LmFKRhgQepl6Ul
vq34dc1VYvfqkh+SKgqHYmRHdCF6rojcBym3UNScwwweSA0FXaGgMPHNsQZW7J2P2JJIG3Fasmos
cOXmPxuzwyN1wKD2ZfRgCEG9hejXD/dIkMZftHFjUKp5f1rMW4uhzCHIZf49g5FTpE6NVn8/F7pd
ih2p+F08qOO+1i5fZrUkk+gy+aO8oCATH8M36Ttfz1VQ1uh0qdP7mV2r3CW3ZQcSG8EgKX9Qncmt
I/C7dS+z+TMKuAr3Jdz3uKE1narT0FNq4VqEPpvYK0gdSlUdWxCsQxP2IUpzw3X/rbI36N2u2mVH
vUo6mtxHwumKhq6AKv9SoE3+0g+15HMCagsf7Hx8aIa2jtEm5byxHqkMilqMCxCtg2iqN3nbvtqG
wV1+ZWiE8ae3HsIEA417ISgnPOVPtFivksRI9m71Yxxh2ZDKgzXGf75ZIIq/ZEuPp9naYK73GiCW
d13RkhNU0EzK9HpZPQvK+L07fFKVl1nX5MTDE2V8CCn290yv+zUnrZ4JAVd/wXyG/j5UtzdTrLND
PnjU8g4f06DMAqtAOLtKTO+G/qYpb4ZRTgW5EmyrXkEA6tmGRSD0DfXbKaFlp6FRkrsVND+uE13U
LmkxgZB9rBg2sBPYq8QmT9B654EUiERIRb2yTX8p2wXKcbi/pPiEp8FuqWvf3hkJ6VnZRCEmLjCe
Ckb0Bl4mLFh55ALPoah9/qOcH8FOVCS9CuY1S3KgUIYZfu3B3nEm8c+bBItLy604s0o7Li2ZgKZd
H8oLF1nh35eVGWJWZ612crFoUog3lQe766kdhPxnS511ZhD0iuywX03bn4qlq2azazpOzKINDfPi
C9QfNRauIfjsHxKngfEnKQIPiVBmwt7SmCKIr3NEQXwYyGdTrMw4bRuZD03Wvw7DRr136QZ0aNVB
Qf7r+FXAyBRDQzv7lY5sZd8hiSZqVMT7pGiAePzP0o9isXAmerqYTcVu4lWun6cHPfiaYctM5Hd5
YMTWu6bHX7MtADH8WljVAgAZEfPnmo365k06RMSNLrPO27i01Tbau0n2tiVQk7SpZYXMwNpiKvVb
L3J41wMa8W0lKNp06h1WwzeDoiZYJ8xJd0s07xMdITrsxoUeblwSdmikzwiwJkr7/wp7cOiH4pMM
KUVMM+gynkBfuYgHRqqitqZIZV38RaX2coepzKSQaTbfZVN50W6vzgtivdVCpOP309qdm4o9VG/f
7DLfBinjGbEHRLNgGwrQZ9/LzOd+nA8GV+9sGGoTE+kjg5qillQuheH3jveWRsYfMC6jndV4Vmfl
PJolBGhgqKMpTjjDdDL96yr7y+tbkPa09idwTI9VqxdAn6qm1/cCiGWnJ+X4ukf2RVeltqAmCtmk
vDKWslUlRWnQ7Kd6vNvs0XmlCzWppbKJALs38N6Ruj76HuRFJ4EGs/3R+1tpi6PJGRv6ep6jRWmG
cWrue27R/d5m7sBD8arMppRE+iJIkL1mlMb8eecb0bbfSE9HG9hSrQPZnYTReyVQ+lL62lP5YIWj
69omL+dBigymUTmpK2nXs6Zw7hGNugVIxfzPHPI4zfaKy8JiyWaqXrfV3PN98D7zMiMy1v6lrO0A
Dg2aMNthiDCiiFth78AYPtrNBEkMoZSgbd8cfzcegULwQG/F5f5Pkjm1v+rIjfg8JFGyYIG2/iME
Ge8wgFJ63gamibPmqKzNrMdYzVHkg7jua8G1x18Ph6rH6xb3+k+aj9n9burwbddJvUNGVJxWV/YJ
eTN9ct3lIysNvC2soVBwhLs53X+Jsqs8WT7By/fg+gZ8o4eJbV29RQGiEadnlf1YyHjKL36LA0fG
6RsVi8Cb5u918Xnnv4KzQdSLEuro/I9v2ia4wHLuUXGq8jr0qilI5GDLMW/4lyRU3cbe/AWZyK6r
cf8nRVi9Z3gAhDWp4LRhcsoMU/6dUsObnA5RqPRkTG6+VmT38WP551cv4/9jgdJkP+/uBruze5Yi
Z0/ER28r6v6iWbYzFG1jN1OixwO8FYtDixc/8cT0iLd80DLYyBh+O7qZOmUcGoU+JubWywtvqTH0
IQYdhtZDo0CMAmnlh3Ig/SVMIEGPgVXYo8GMnEQd2GofuAgSI6KW8hNtA+JYCW6q3wup3i9DsOYv
AN9rUTYUM0ApDev9lxW2ehw02je0LRPxPf3jEqLhfgocnnNCuVWWfBScwfXmYwAompj3j5RpTVvD
zm/SKWH0X6oF7ker3OoVT4jOBeG4RatinRiZWbq+I/ON3D8IK7zrUX4Vn+GMeXvkPD3GoFD+poZX
DoYFJrcPLzDP8uVo64zGfmCw3LhxoyD73jmzgPCYmYk0j6eLgvuOsIRuPFDOL8Kp2SEVktUck8To
cZKIBWBHLUYUqp2QMpgYaP9uaxnoF3LifEDMcl6lKoZKCaJmSyY4F2pEJ0VTn2vLHOCZ+AALmIbK
EVgRLSU+SgzbqxJ1GSUXx7H8UQ7AxINuC6/ub0ANvr/ej+Qt/qV3GY0Z3M2+xOeiIiV1r04NxnNv
0lIj+6YdZRoTIf9Rb1BXb0z2PAXulXvfGkXNtiefD8+aSgB+GfLfZP/a4/B64of0g+QqM2OJhVn8
ne3BK6ffzhEvXS6vcNynymY2XSeYzfT/Bd8H1+bsBXFRFi1/PmL8EVzlOzXTtws4cwE3n7vweOHY
rMIqp9Go2GM7dbQC2sr+nM5z5Ji8lR2kzbOUuvGQG1Q2NIBjc9tnM87PQh5sMzeAPsev9uUXs4+n
fGCHrYvQMhdFvrFCIExZrKjFlUNG/i2SWR2db9GD17Q0vS99n9FPd6FmzbbmonjK16e9/UOe8zNU
AV+67ezM+Tij+K3yjdBd48s1GuQQ0g0GLi/VFVI1aR76uofAEMF4tCdWRoq+aX18o51OlZTueHar
lnsI9h/YpJ0pIs7IA4x6GnZznwC1j3joenA4onveUoJd1yPJHVTT3vu6or0QhmK+7qkGWwrYFFWq
EzccL1tINz0KZDQZY/rYj1SqrBx6p1x7T6DU0DzQkNmllkSBZliJqna3HCbh+JoKzes+VyiIJ2Pm
gwcfdDo4bWEyN9IMxEKH8nGwgwGK7X8t7jl49JcF2GbnB/QN4KYqQDOViJjk3nKJTqfakz/JOxof
lNOt1Ro6+N8M0OG3SmHLArQEXJzEcjTkjHnaXBZl4ZUoRwC3SQt0ytt0PoygIH/RppFaTXwvcw7q
WsDsEn8xNAXktTouGR96A2WBbE8GDQ9EYGf6jMUJbywpJxlXBHtOR/ReVR5f6xOFje7g3M4mtgd+
GCvqFn9C2vL2GubQ3Yb8o4RTJrDTr+kZOh7c7SfQkPt/vhyJds+CvS4WZG6feNJLh0cBIrs6Bx9W
Lcipc4z0D1CqX9Qvj3ED7xetCCUD16t94omOi1ud7OfZHQNBwiMQCGaNaIYOCCG4RjfYPTfRVYF/
mXH1JJEpMlvchiUKhUc2PNzesd3vuNPyBuLI/XvtDtWla1JuSq2pkXHOirFwm6/bAlwkPnF16X9S
ItEWd2+MizMJbvoOK+hlLy6gxaLiWS02W/6ksSKZjwhzihO93t89RKST20au9U9E/MLr2bmC0kUB
HlvAM6CjdAwnO3K/GYHD/kF0AYmP2880vygDirSIs+Ix78I8kObY0YIrnZ280/ruZtimKO2lRRwO
fnW+A9m/5n4p2B+XjZd3pmdAkImkcmCdreFhWwDUmkQMCB6Z5wfE2xykMg6bwKUzJ1UbBcue7AYn
qlQSnpgaDqswoq4dzTfU8Y4kKfAcFj1Stjn3TcWJWJyhZ+i56Y42D+1ZXDaIWaUDJV4NmHUL97e+
KFullC34bRfIpVvoLVCl9eSu9vb6WG+JhqGfZcyWA6AqKN5T4YJrv1QsIwb4+JSvvdsxMiN8K92o
Yfrdrsm+iCWk2kqHpWWrcwW1VoVFvqMJR0Tem/aCJ/zeX0+aEIFqAQ3TdkywXku1MulUzG1W85aP
Bzj4S8mlQvVTYY4BNquY1BiQnYtwBHFt9rYLZ8spKei+5tX8ZLN0y8nVVWQ9xexG9TJSi2rVq+5L
/M9KdYjcM5fZ0kpEQ3jHDjg+B0sRH7wmZeqV4Z0gqBNVb7sKgysuX5vbFQbrZPRHFwFx5R+AXGaV
yXtd23LfmScB6Zk60ynBqtwX8GDw1t33QcM+OAh4dqGZcUYUpYPcPcYaEF6YzB53UNNqNHSyJYWv
RMy0gilnP3zYAcu5PdsLAeGLXwXOAM2LmCRN2y14nsvTp4q2whOobqd9o6Ppzwr10ieGvKxAyJJw
HvT+yF8lo3oZ2ynsM+0IWSQffVqZH2qMPcjfazXORixghifiRWuOaZxTBGofSTdnHlDZtkO67Yuh
1HDvABi9O3mLsNhvmFvkbp2vd3WWasIrV9z9QfX8XfXonKH1cqug2G9RC3meAJDHjt0F9QkHSAjT
neeDKtyuQUTh/4o+GeRuz11on7GHI1fwioIIVmnwBMDn5vO+8Y8Zi4RcVm0yVoEByTP8iFSFyByE
zjX1jEwYPlhLpN5d1a2LTPWtPrhSfyPLXbaJXgVUcPGkjVafKpS8oAIzzjpEp/9FoW2OSanCJyYg
2H6xbvEmLUenmbl9P0bpqac0bS0ZEY2JIGNqKa+LV44PtxzmSscUxVsllF8i76SaaOMRJjxpLMuX
hhYrx/MPTWtIwEDw4HGyvYmVfHDvwpu9w90K8J2fItpE9NHyoKZgzZvU7uMWmYnvEcjfmn9syyAt
3hZhLhk9QEF0DVQQjF4/s9CJibBNzdSayn2gywjK7A8hLTzBkQgks71Z3JZlZ7Cbih/923y/BEh2
LAxuXwKFNikwZ9LjXvrDNheYdbqTQkBclkUmAElfslwH4lKLy2o4EIyahqZUpjQ59iXiDxpGFLmH
XbXAGRpKAD7U34AFebOXhKu9JBvALQvok3pB0yFZfcxeJIFnkDZq/lLoxfd8c3Wc+ezpBBrIbhTh
jn4iNNVqXFlCirloNbDAYnTcqFz1ZpVp75hlR0xtntU7CjBnylXvJMSlDEHE/2teBUt5xZO+8PE9
9gMWic06V4ah9aH7ZROl21cR69KyVna3llbk9pN11t5+jJ+7L5BHFZJEFdcwqhCiIlL4M2qF3SMr
WlVrvrboRKkhIjyTDU5bz060zIUuERob5m3sjvI7rcIHioqYgncKwptKrbCQIAdQ2tucjApgGtuW
V2La96tcLqH8aap6RWCHzCCOy483gtS323zS7PfbsaF6e5vNfpG1WRQCAFAtqzxp6xDqFtnsbIfO
jAOLXRsKGgI40av7ETNbk3uWbNQcJ072WIAKJyEQ6OhLTBUVzFGMH2JULd24taQVYcoldx2mWYPK
RA9hKzeDxXvMaJFpSyhpg6s5BHMWwF8oO41ZzMv/fcFmL+jaJ/q1m+9geWs+vsJnQjyEjhupC/RV
dtX7gibWMbDyr23Q0w0GpBmV47IHob8nT7HvgxqROHGgF//zRmHS+4DYeKL+lVjZS4qfxch5nZrc
MfM8aSkT70gSfLYAduzc97FSWuHlS3opUiA5RhAi6VmKwLvsMBT9szS0DMGBMpDktOcXHXrKSh8r
y9U8XhpGfnRjsC4wBC1Tkas5emQk8gVRUdS1G6xjTLjDs6t6SgvaN/XTymybik5NPNQb8x8gp//V
PNVp7DR3Nk6Dz8H8MkjBpsRwnIAKgSFpZERLJIFWWiQFEA3WuYa1qmI1m2vzzXdB6zOvX7g6AbpM
mgOmMbmYwi5Z1D6F2Ml+7rtteQTVl/LRFmsfmDnZP5O7ve12XapZ77pkjDHkIbKth7cJXm7vXasM
mg/F4WgtLkc1Vdn3VXsRcEd/TedQTqnUgBoB16L8drAkXQ2LxDbvfZdLQyqW0EAFi/HqDLt0Jylq
gX9u+MjiEXqlD1dSKcamrReM1CKxR7m5IvMHG7pEUC7YvUNMiQi71u0WnRJl7qH76Q0qvLDOyQfr
JOTXDJedMtTxru8jXu7rl753ZU+2xRBX/GDUhzBT7DQKoPk9jepZr2NyAY5OZisVJFpHC8fUu9I9
C9iTVCv3osO2zMOZcx/GmQIMBTawPFcVw1GNDGr13d3EkJpz11aKiVh2618eGgsHurGmJi/CclgF
6PTrgRctWGY/5LUlM+uoeTxJPFLtqfGSRnmgz+mD4CADzZNEC9Jgo9wcLac1qfsHXbaWmElX6Ihq
tH7MiaIZ8qzVxnG/PUwcGP+o5wCgymuD5VPUfvQ0SSTpj/anM5N13uZPKeB4LHA8jQLOV5WgDap2
AhNgEC9mOoprjVNzDATvV1+tgdreBQhY0J+VhOr891nZScjaj56myBhb3gXYMRvspz4puCBmtHau
xq4ioF5A5OqwEPxstUwfLTefpoMbJG659ik2esZGHabU+jA6Nd9T9+IK1s6JH0bEOUGg+LvZxAYF
a4fqeLldbbv0RIBF2FDRsKiCRIiw2TixhsxYGx4P3a9m8FpLS1ER+5H3LIlYWnxMxMXHeSvC++IN
+MsjhJfQZP3P7G8tbdSCpwUehetg2pAWqkAEu62WgVhm8oKdwYWCMDov2FKEsbkubXnNQG7rjrsF
cHC83ud9LFWZPtZBQCwAvIVkmNtVMjmJaR7bQwirRHr/ktkTktKV3PtxfQPjzL4PKzV1g+OhPaiP
jnZkmMW91ZG3BZbp22zahS0pErqMwJN0oES4KuRdoh7fZici1bFQEQdqe7AlZNXpAYSYAU402xD3
sm7M7vsMam+7KlvVVD1+cAMNd/HfV/iUtBYWwesk93hYo5QbKhDYKQG9RcdzQIPSYq1FZ5n2yTvq
EQgoup/nR0qRBrAsJqY+tgb6MyyZ39yV6MdDwajIqUr1YTMbAAHMOwHHC+UVp31EGw7sZeiRgcYS
Ik7Znaw67/Jm7qZwfwqfvXGzCKN3cVMDem539sfwdnWi8KPnf6c2yLRsXj3NTdfVyLaba2moqLwB
WB+QHX4o3y1EkY1VZFedcJGzoK45+0BkIYpl+ZZYj8WnlQ64+D2W/B8K2pD1p+q/182VvTPcE44E
0/vH4HA18QQJ/mVmcUiuJqpEvlNOjdoS5T34dmYGueDes92y0r+nSMZmxzQjZVZ1Kz8BQ7WxmFwS
/CMzJjfhlZtO7iQ4A+5EpjoBGROzndBdYThAm9eey2A0hhAxBsNs3n8PlONaEsZy+fM8dBCkfiEp
YCtI3Ofv/ArvjhSVvlJxhZAsMpiI3ommGiZdmTKUNVsqAgHvQnIdflVj/EayZx7RhsABSFwfu+MU
0K9yX/CMX1qi+N/FwdBGowHYL9bcSLdGKGpvHmRHyW63VcTTi4uQ1vcrKPWxduEhTvbvvtRxeHE6
xDtvdyb4E2Ti3LQ0qWjyZ5XRy5DjHzeIvhvEE7z1KVCDtVwusILAavrk7tBlFlkT0zxhwXZcePnu
+uzgue8QcYbUObim4o6YZjX/9Wp0U1xAeIsFLK7qS+u8EAwDZfolXBKEn4YqpS0Yq9WxY03S9Z1Z
T5Pb0O0pE2sG6WN/97B1B8fJ3vPpECCzBnb+dWnL4dT2DAephgn/dxgEZapf/YGZsVf2ug56oPFA
RxGMKk+FAFtUfdfjQa24gedxIgPZLurAKTAjD6KwjAoKTtu4C2w9HxRzEFcTBkkR14sxJTZMID0C
tJSrsXLkQTdM63yLRrKj30VBekTrlzZtiLRd05Z/34arduiT3Rh17iSOG1KXt3YHnaUKGjtcT9D3
jIi9dD9J2XALit5f2CD9DxSoq+T+lPAvCqVqWa5RmqwxIwfa5K+nCIOoQkRgvCP9zh2iqiM/JGbK
mTkxvVExIdQtC6g5a0d2HmSw65XYQnY0l2ze2BsDb53kiE1RBNVoczuNab91fjWtTAVcDjPx0BkN
KdVjqZmpHxqrLFEjPhlZnnOjG/ZwmvQv5IwVe8DIlIKVtE9PL98tvIVPTUl1yyvxSRdybzoPVwnU
qMA83W5VnmfnTrHZpgKEOB/p6F/1tOhZeRaUw/CP4auHT3LCs98sK0FsF7EVzEUellWOmeytk27L
b+NU8NJHXtWz7jOWxwumDQ7d5jRGrBNF6czi2IUXB6le3z63PxdwAJW0747pc9xF8sx3JSF6Ji6k
xM0hb5l4meICu8VVhDrGtDS4NDKDf4HkddbXYr9F6ZeCvR3YUsgyQ2zJjIih4j1TQ7K7uJ3oP77Z
jRvdTQ/vUCVYK/fg+dOLWXVUpBOtFCxfEUKocRHthIvIVC9tIzYoJqPSDAT9FhM5280DVxvkXumP
22p9DwsCdH4By/rNiVGCs3/tPq4p3i7VXD3nKWq9stFXGiliZPjAAZtdlgAij6itSLlCNtLdNvOR
rWlakO/dlQmeg1yPamewMVjYYYpXcI3S0mH58kUnqd0Rto04hedUDc2cECfR5yjgJdphNbpzqDke
QhMDCozygxHFwMoYveD4J5DWiICdLpGZDFyFWi96AoqvS3RzzVoPle75bUu0NfVtNrlttp4VAUmM
i3l/+GJ0n7Fn1I6VwC0YZUMJkop+6ddylBjyHXV8E4k9KwIIRwNlH6bIFhQZ1Taddqxvfq+hAeh1
lg1IQ+Lp49luNEHL8Ab7HRIYrgBTnnJx76MQKQECFTQIpKjtIp+cboHjlQ2JpVo5Ln46ELk6PumL
xWWXeiEddl5n1x5Z8E14hzIJqy4vgqCDkZTxkXmpoyYYwZADjFvpT0MptkRX8yRCvN5nOaNKzY1f
BVBjVGPRbUefBdhxvb6gae/OVJwlvFJK166W7omOc2ohPN30Q9MwzAreJJZFmsuGkhTCeIyWAoBL
fnv6oCODw4FzVhKRlS4bIOUoj0vbDr/9+QMWoUFjh6fQjxgrPy6WP5sOj/6lJ7h4yl8a7/s3W60F
r4jd7WYHjvgCoi4/Dp0JWjnYD+MzBymf59slbLsgchuqK0w0wnbds4KO3nCAGxk7d1nwW7lin/RS
lvfnX1wMcTYIlW+aV9Ub4rk6CIkiDQtSwx5n4UFbGNY/75Qr/HVz0cs7djFeStohBSMrt/Gpz0BY
GKJe8J8px/tTsbUrZfPnZY++L4yMJ65yINW8966KHzUlce/m0BlAvzjYpW8nfNOw+K5RT01ZH/8D
62RVjNvqHpFdZgXQzj+h9kmDL04k9i0DeZUsRExnipSdqnPH9KszWHft8zPh0c6sljWmxyXuJQCu
CzpzfdPJG0xufFWlucZxT6BTrzDey8zZ0UVqnCC/7baqTTJ+qEVNqHQXi3Dr90XqpObJwSxhXp9m
t9vPmH2pGkL6vT35kBZEpYVbHdsd7AILa8McygML5QCE1qNKw/No82s4oVMzkDoVhls3hNvAUwtI
IYtHTnjW8FAU0aS3TbeqODZU8HTHS2T816UfOyQ3OExyXCTolNHq6/P5IALPQCclFUu7ShGy4nYz
vbCM9p/FQ9y0JWlgJqnOEkSwGfIUIGM0awoDzNABROHQV9TEU6V/1HpV5NxNv+oUj1Uso2ucfYsF
5YzTZBV3JKu8HNYWEguzBonvKUp90+wz99vSQq//w1vwutJxQ3URHVOxUI8V+hdCwdqBYnEEGgz0
q+FXXa6+zF2juEaWF5N4bWjNK8mL364ysAApYDiDnwvbrurQba0AFRuXGehq316gWJUaCCZ6IGj3
zsk4x4V19AvPcBcaxbqgT5TOp4Bj+Nh96RUj+hi69pAHAaPvv+COKLdfxRGl3En0mbpgKQLOvIE7
VMIj9mRdeyel+f+4aK/lYRRjJcU5e2xYKCaYMqrpV0Wpzzu7Br8Y6109sl78to+Uc9zhxUjMQ9v8
xGPH5u41HAfzqaZPhNTSJunLTni8bsePkqvDDJsYFEJ6SafF/ZlO+1zvlQisnJJBZJvaFb4rj70U
HVrdJwMjY+SVrFI87/y/QwUHI5sAsbQmIx41Qc6zXf1Kd+pVhzDafYWzAOdtTB2+ucOVkO0CPVLc
LBWi5sekNsPzz707+BcvXHkYtbO+PSLR9E4k2GU1EEmsWjxFhcS1TRiVdroQCrvSTI6HQ9VvA78Q
PPOE4fNC3bR8jNqPKAyCjjOZsxUi+DbGDe5XOpZzoxWQVyleIEu7q+dk/xr4RsQb4Ea9VxehZiPb
eBMb1JEkzsQ394QPen8Ru6UF9UZpUSFHtIqU87oVjHcDH/euMaCad/hjnQdWlyMPChugVqK8OaHK
fLFa6nQ7zPHVxY+/+GvhmyaMdbRzHZIZR39UyaaVyocyGFSh3/74fAyLyscCoeCBIYtR0fKVBHz6
EmGlWAPsGBk1dDrR/R+VGYQdi0GSxv7F6peXCvEU+SNFQC2tU4Pt59T200Rr1Hj9u2yh5FBHk5Vm
+MASUBZMEZVrfe6UKpAyoS1IQMQ/X2cTLjOzfCxo/eC5aFUg+5GxO3J9Nt4saDareMABxX/PDK1E
MeKV3IrCTSYWnXcSb7hUIeo8KnVwk4Kt9gK9X25fbtba6Q6RNtDlRdi3At4JCzop+2QOUuoQ7VQv
Zvjw5PCaS78F53WW1whUas4ROTmGhMd6c2qvby4hi56qSm8GLup9vPExRz/rbTuUy3zO2wDV9k8z
dz2Jzje0cVNWJdODA4O8z96O6UajZHnqYh8VZ0xFgHZerdQc/7STHo80jZ4LrR0DdMllfNZ7xB7D
T8ywX+BYhnU1NAfzRArz0F6zkhWCOt0VdFTEQPDD4luhDDzvzSFU2QMxVL48FgD69AQF65Gccrx8
dqxopdEDjJoHeRxB2gromn9kEY9B2BZARK2zUhNB7ylM9zFuF+F8SB3QjfzmaiVA3kA7KFwRCgGS
BrHcM8VoshVa7gu7obuvXuKBcN1mSZ7ia4WbjsHrsAzwZTXn2I9cpMC2cggGmVqQ5ySHGP7VkdTD
0fx6LnqyUJInRdKwVEdDBQraqXbnPyEWbttMDty1iRtdCPvrZYp6Y38UXyCqvUvAWHrpY9hmDzBq
3d/FuGE3DCtjfEEhAZlThNk3jkL43ctHLYyYfwtAfhgr0wWvTrAOZBcSDyir0JeAcefGV9aJewyq
qzyBuQTnVSBxz9L/9m2FFMJac943aSBYjShnAMGke42ewdAO8DDzFF2OooZs+HB3VCm12zsodhyS
BuhTrWq1c3G077oWhWURqtF3cnaKCeloqeDasNH1rStllciheC9D0OS8B6Mw6/YRFOZu3AR+GBuU
PHIiRa3nFAjFbiEXMR5lIhlGhuKKhJKxbnscnJVlpaP0swPu6Y9sP9+fm74xYYT+6Adwg2eviRrT
5dIUYsztlGFvaSPgqbTT7HKygJIAQCyjC4xLxAfKbq5Lp7oCeg1l7lVxUgOSMpPy0T21hgVsPSNA
OXpweJv5bjxQ+YlsmybgSE4WwVM2+uu+o+bF1Rew0xtwT8sRinUaJubnGfiUKzMUCrCuMUgcu2ML
uqAh4v1pl7tiN4in45ArIYUZpIAak56ERc46smgEUPmymAHsnM1WSF4euAjV9i+tnc4cwIZk3Gi5
DhbnWisBGrtrGpNz9O4+VaD2NSpP9795+knwXidGiG+AVUOfNCFRfPmZoNOP96qY9tYPFM6qhatE
xUlNo+cFuSj1sGQX2r8ZIbVYGs/r8hdHLzwbIqhA26aeg7C1bDCUANaynByvEMlLL1xb8ppYVNen
kts2abPyIQs6RDIVGdGfbDvFwNIr7MBP06qeNgZAaK8pJUNPsoSHz8079FJenCw9RzDWQVLlKCLT
ytktvCDmUa3F5rEUCKwd9QQCBnHqeA/2zFpfoqKgA0jW6xt2+rX4NlgfE5nZE+D20Js6TeHMmTCJ
TKCy5MlEpN8hPUogErzcr2oz/zvWfeg2FJoP6L3P0QULlg64XI9XulftdlzArEyVzGplhS1k4LbB
WoHQE8upMADyRgkHPcDf9CJ8s7tVI6z4USI3Ns0Zn7h8S6upTp96wz3ivUGVr/dX+crEAUndmTS2
aovTIro8nBZLOl1gYh3zy4WH50Uo6VsptY7MF6mRFSxgco43Aw9Y5BImRjHGcMeNZqYl8okDsYqX
WL5amy1lIIj/LGNScEa50hK80NgnzKgrYKqBS0xtoddwXjlWbmyxCOgCNCa+o/+1Qr5XLGi1PUGH
P0RbqqAO/WXIaFEPPQkJK8qXE6wLVwDwOv440IbhEAM+1rVvrAIzRvvSIPcy9QXQc2kzwsaaSaF9
tlnYchRm8P/6azCIQ4bXtVC4OO6//j8lgKS2o2gCNz+QExCWuaEiXOayiIxTcT6ZD/A2aDq5PWkd
xTldN3DMSF+e6pp9VWbJL9Z33EB3B16c7xHtviREIYH3wH4NM/CkfvjWeKukTCOq1pJBE5CfFPYE
/Dq/eKFLWrLxeILtOgEBnibhKOJBRCerRTmql/QeX+VMe0pn4Vxqc7YHzrxvU+UchzhzBFxUgCzN
U7ilr65esJ7xDCFrUa8mdM+Yw6++5Klm8z8GngFis6zDkWT88Y/1BBvf48iou/HVSfU1QFexmkby
5f7NNP7VPPsgkQhZf3ZM4KTqzQM2RpgpBBOsZUQntIz8WvlcL8UyKdDbtJMcXlGIH52s7sSuogW1
VtanGu8fb7ldDzMxRuMqBs1AVnkBXpACKLoov99KzakDHELSFlD40aRzVpKj0502MMNq4HiPdihC
Es2AgSV2tAQ1D9dHQrNwLjv1ybwihqfoaUHDITq5PNGHE4rs46ExDvBVdQ0haTqWWDX82LPq1Kml
APJT5mj0/HtseYK1Wg3juNcWkhexHV7FCX9LbvMnlzOHH8LWVoC1PhIklPrcwAygDmtGR0j7JZBB
GMr/FkrZ0gFfbexeEgeNt5AbNLB9cHnTojW1P/Kk11X5GzLW2PmtUPK66QiJ6lSsx80PvpMUW6Oo
VfKFGK8tLig4JSPSlA8fArU0kSLQloflm7CRZjey9Si29GxzuzgApWjYln8P3aep+ARqOMdSXcrI
pR7rbgvMee0R2VbpzZxg0cgYjx653HkJ9u+ZfeLRin6zD7bP/CekQvLNvWD9Dn+Oy+zyfiG7QtvI
hf+P+AvkNvQEFgfKSQEPiEa5vhBNKmXDq/IuDQXZJaEYorFJZXdjmv84QhaQ+SgQ1EP0ZWcR/Zx0
xKqNIuFl+M1h2jmu7f9n4y+oijcXKR8EeYgrpslopYgsc97QWc63murpWAlQcAuRNvz9qwB0X6RZ
M6UthJh58ZKYsrOkhidXCBx9K13Yz3fy8tGrrTstRLlTvuanLqFyGyh8LJv3ZYHGUQoQ7gAlVrmi
uaCiUg4svc8+Ix/moNQitYimfcjL1ZfK+gC9z1vzVckZLHObXnYgYSlKnROctV3o/84bOusbuF5p
zW0MmsobnN967FApmSdJHG81y3/4d1Y/17edgl+XakquZEbhYubQUN00aYTlTvZbGcFadVf2pZR4
kxHJEYHZHpYAnmUOKN/jL6aZSotyc+7ZX1rpcwEfyizOKV/jtUNzn3IqK9zgS1PFWW8/fPOpjrfq
1XA9B2yXIjyFIWAhTh9gOlwtNQvcKPZWCaPIzSXOz797uiA48PbZ20Gv5P0ADnlZeWDZVlxBm2TI
HrF5SiJPLm/jFS37pHsJjjAeznqS5WfXM4GM7ivc831hMfDxUtPUVjj1paDYoFqWnQVKX/hJEa6H
I6IRZVK2S5ZZWtSutz3zoz+k36ul0t26FjAX6WbqlF5xL57mZAmBIA+RjZ/qVkx48iVvoSpQrvxA
2LH007igo3ra+iQsXV4Gkyr+Xw44PEvV6s0H+sKM9CchRBtBsyAXh9AQkhorC+QGBRvLU8bqf2Fe
0AT7E8enJgeqz22+qX2sEehCN5lSife4HDIGSZCkL8z/Cj/KTyiD3E0o1gnyadKVtbMLo9LdhYHT
v836VqBRUmn5gzEg2XEdhFlwMUYTRvDDOU96+Ta8jdaP4wvLiy99D57UYWzftX68M4udlX4ouqoP
afoaafub0Sd4S9U0E2wAmpuvadsGMVMIS7g1XdagBwZxXzenRrU3VitSvPp9av44b0iKWXMci7l0
J3lxpA2J6tKP+D+9BHdZ7JQjsxMcZxz8ruAjx/Bro0rlKHVNWx8pZUsGiTfkjNymIJeqsRq0D/qW
NSsx4TzKqv5erbdstTu64luCVufN738YU1pnHwKRbWX58GGBs0VbZ8Sq0NBMcVsCHYX93+iLb29j
2ExcfZPLi9ghaRtEFY2flwZhnzB6b2iwyBM1NflWPhfF+8gLoq4I0WKIoJkUC5WPcRjazfYRUFqn
6xEpZlxsgFQC8hd+IY+fKMl8Wv+NwoCzLHK0FneRXHMVVLQvptjraimETK+lEDI9jwqfAsU45ALl
nCyuNCgiL3KTfCw9bbncz7h8Qva+wKpbSfW0FSNirC//foblDSDtUDT675eLH/HbXxROPutitRB7
diLE4XFTnrx6/cVdSgvkyZxREkGg/KyE2oZbRviqkvfOzYfONA9MFAqM57wkTa8/05FGwv2htB5G
5v3k65tbSZ3zUmrpAbU+6TYaLY79/a/IWcGxRw/SK4vQeDbXNmgQD0n/+pddv6WriCZ44sCNmh3X
NYj320Ep3dyd3huT4agzGogNXZEOFGzeyVCbqWH9UlYsVKwFq45nVJk710UuokGcp3s4EWHQ7lwN
0+jCzePAkXvk0q+YD2eCu6HsvbUgewV8LgL7MSKYQ9xEfG+tNBcHC4Y9unfTOU1Zs6AlnLx9ANU6
X4kVjjK7sLiej80thNpIQVfwGT2VwDwBNg2+o9EFwgEI5KZq5j17qI3A0FMOiipYA/LMajLC16Xt
5vFbcrz4ARGzt9jh/3gft5nquOrgGUcTbOINho2qhq+AL73fq71lqGaMoHTTgsQv34b6WcGehau9
ozGNbtox9fkroeLYt2bBepityfEuM3b9CBP9F+9gnF4XY+MrJJQpRvz0M9vrCnYxVKBRaMIJaLgy
cFA7dRQc7mcqMgHelJHsGloiy8b9FtnxJm+RNoqSijPmOydvQ+w5zZoAG2LIxnX8EHbNjExPK6OV
X5r+ndn2oe1CFWYiOky4QwWDblD7/Cun6INN7AIDvUy0iXT/WslPFOS8IbH1LA+YsAly2L9zOsWR
Er+0EDqrtX21KEHuZWEnyqhEq91oLb6uWKgdWaqdrbpntSTF+IhcmdcfgHjNX3uuFVTgSl5ybeb3
Rijxc+jZvcwIZ9vnUwLKlNshlZ/MNyFRWtEvtkyHE90UxkiPYAlaIYGbPPx3ECI2sJvxaWy0DE9B
PplnQFG0eD/yFUl5PJG3dMuQKXSU/jZKuEq27ouE3+AkhTl2uSZoFG9W8n0UU4/4gwUdUwRk4Byf
GAyOn2GAI8M76SdfWlLTr8xKkNIDRbwShifwVJcf2rlOKyby406YFBVoaOWzthzv7g6GHYhH3+64
96XVPi+D/ebQpLwFYUiaT96XU3d3SXHqpb3sGmiQHgcwKPS6/3TRlWoRwZxoy3LatpijRAxWTero
Z/qQIKdimvC76GtB2ldEWQxNonNZdMScETcss7j1qQouyTqUnZDO6No3xsSKIjF+F6b51stpLLXX
AIPMdCSEGVD2QApqNUTZ/FhZYQwmSv7mNM3cIHYXpFHcjZDE8uVxOpEnj86GzZa8J8PMjnRuya9J
xKMI1FT3tJ7MVReJ9Q1n75kzdVSUxSmlZKnROTknjJ0wUTf5pIoV/VAuL4lWkqNmQz3CNm0Zri2w
xBBDplZ+6XhwB4jW2GYyzaJ9tc5HToYwuKiIpb9O6IGWGm/R7ETg/lIRxgT5VlC8CENU87KlLv34
jVtRvr9cPJY3rA2RmjcH5Tt316haEcTAxITRbKQuqoOapC2Xr0qm1GfVhte0yGacLVfbWXJLlfeV
ChoKJwxO9EpW+pcCdy3lutK6N2j6BLQgy4fCrEmRP7QG0+rsTKDmek5w//KKG6E3xxo633T4gS48
ZgeE41WJTwCmYBxJ+42hsBhQIS5VlqWLf/9vg1CCNOMdRtAwn1jDw7JFZVyB6FEykhlJn9gO3gSJ
2o6muLE80u6GZiPXSUgDeFf/adDi5KJdgZlZRZo1VuHMzboRmrUgAzSvz1u7y1MewcH7n8BidJnU
k5NDQiFQKU9ZfN9XBl475UtIGn6EKZ6b/EfBoAZTIREpOnhMsl1l2H7dhkTsDbTbnTi7tK2jjKVo
UgW/MsnUVvVQaDXqpRJy/t4Cs7d49RnA1on4PP4eaBJIE14/xQ9BC2SZZsxWhHzGms+7rwslWjqX
5hUFBGVGzqWSwIaIjI6SNcMIDQO2KYOTdx63qIAvugqoFgHQF4W0vXxDPSqtsgTHjGaAbEp+RNcT
UBljEWZANlcox50LwR034Cmq6IN3/ZiUTDo/3WnvwVIe6LUmgu+zX6ENA1IGw16uSv8RSSFbbXwb
psOH40Vcd9DlAer9N9hIdVo32Bqf6rlI8WD+1AMQ/CcRMf/cTgPiXcZWnLJ7XYYIMb3+cnNSMXTZ
3a968AM5x0YciBWGuFoyy4LCBeNmSVZKiqtuTAh4nlpuz5Wg7RC01zpjT1YpVDweLKjNHq/HRJqy
2ObYPsgDU7poKT/o3JtfMBUB83ucLa7B+L/mh1ouEFHhotX5lr3705LwZj32mrR+L04bGu7OP4pe
c3VaQHVf8Q0nkuRy2BKEa+O4qoEwk2QwUzo5lesRwuXNH5ZFNQbYVOuquT166Arn7x5hkXzOC/vR
iLM11Ved4YN3KcwHl1spbBDLbrXcszWfBncOqz+DGs4rCGOLljqcEfQ9sYYpkZv22CgelX/u5IGo
AqTeEorNoG+OLwQoZRpxeDsO8NSXJmRQxWZUVrtXwZ2OF0zeXq+n3c0yHZC9RSaE1CmX7lP91C1U
5e+rH51w0ZGSwFSIYHqTSZ31IW72DDJV5FEDCvgyP2WeSzvXo4v5kFhvH5+ixtkP0rt3lHta44gK
vkvg0jawBVTJCyjisWfwTcFYzKW3b7/LEFQ9JybcW7L6I/UVmSR+QHed4xeJvuPSG81ygIg80vk7
qFKlx+jC7AP14JzrITZzuOKx6UsYXlHzXu+woAoREW/m3BZPYaSJJG/yT0n2woGTbJngXkuBNP86
wFcQP2oSh4M93ijw8Gr3bZ+TGnGqVL8h3LIz1UjkHPN9y8tLfCoSNIQyFMg8FOk0DEuVo2UKhGTF
GcKtEMAXSPH6OW0u6aRz5fJhOEhghVcCraWPytLaTFir/YKcpYgMBlRpI5leXYUIHBcsKou5oZEy
Y4jFyo8W+HNoVRfDa+dM4tQZQB5Zlvuah9Cbf8pjSCamM4n5qn5BpMlmYB7/J5jyN29DR77yf4TO
LRLaDGuj6cibFTQQNLdVcVb9iAFhXOKjEWgtQQa0HlIbv2P0mDTn3w6a7P6Zn8I/I/lhM4fCohGq
eMhuQn9arLRxPRAlYq574HenCFIUkenr4LtUfSdJtpJ5jQU/UnAssq7wCVAW5HhWtN2W4AW3COLs
tvgELm8DE8eFX7k6yf9IAMMj6PqTgAm4LFnJo1lUVWl1Ri5xDkGy0fgeQ01ckikhU48r6ogs10j6
6QNIgokPYzFfr5mFvBI6a4QBxaOxsixaATTHLOiXgGb5HrzW75f1Vp2+O11KeMD68mnbeexAIUwY
8/jK/fRpuefEXbpYeWDa0MdsQzX2bN0/rELWr2ftHgqK+nWUEwwOjrxBXein060UpZC7+jpR5o3c
4u7YWt7pW7O4OAXVgvtUtENPyUDye5ZnwJifc4+2jrQsMoxteOmmdIVxqoHapXeleRVVUjlSBe1k
8mcxaH2ujofOt+bLLYqRlj8oALSZdM6uzINGqdADLY7YscM6hZ0HCG93FIHOPCOKD3MD39Sfv71S
nbXgwsq/bM253n9aIw68C1XuzOHmEXetwzrXwIlhQ52CiBve7y6R4zjfmcZiXDHL8iRjHjYF0fTJ
6bijMv9PoftnnwmUL+a1m/VKWnv3wmIHOWmKVxSr99sekqbq7BW72YmopeekrDPDfV20qQI/hLyY
+GQOrtFuIZFG23Aa0yeMhkYy3JFtCYsKi0E5riBY0KvLFQruXbETG7klY5he8g8mA1bpG6d5/I0N
tw9axARV8OaubiVBImsquk/SN7XpyV20q6F/IsWBTMpO2S5pDBLEEQ4ANAh1AsU6mSsJ8QZrLNPZ
yCyT9t4YTOiKxlild/wej0hwzt3oU9NBRTbKh7x2Q/b6simThle2l9rMTnUKtKiEMZXc5wrLPS15
3HiFBW4PTmfKypNhmbgFZsBeLpYG2XDbbvBnpbT6vdzigAdC/CGkrfY2z0iGq4JNVnnQCuOtcfnc
zVBIHSOULd0kL2v5ZsqOLQbzkVoXJf/fYUMZ/NTVAuQg4zgPiQK3e/6OTVel3NSJFpkd7/9XKWEe
Oh2REQV/JNKOzWn4mAcxzYcSdgm5bx8AcFVJkRZ2zV2x3TD76FCB7cR3IPMzAORPbOeREoVN+1sK
y+UdfPdbhe3rlERoE+iHHkXuEzC9FrTCZe5DhsN3bdsk9ww6ANaMzWf+nXjo+v2diMF0HXHv6jhN
17Q6NqjhaeEYnjx0v+C569ml8uvkLChFDRczUYXL+xovJ9HqH6ekRPrt5m1bMvzdS2AKZJ18K19F
CtjtIqWh79mQEpAivGKX9W4d+ZcSVBZfLmqSQXYjszQPhO0vyWN9Wq1OEhMESMGBeFgR/rNKhxc2
k/X7HUDRCl0fmgimtm+SERfnHDirUvjwmoNLzsSfSJz8ovbueECLWcra5V1yRU874VQeTFrMZ3rS
LEfpeBDFIJGTDz9fvIobEfIn6PL48iacFln6I2L9tj1y2M0gAjGsMcZ2tvhfqzu0zCMcm8QCx/DH
cpsGTwIAYu6LVvU5nGIkZ2IoxHNOppmuVmHDNpOViGsX4jU3cTii2OuD0ue0QiIKLwIZ7CE+kcwP
QO13R0Tik7Wkg2F2rUzI/q6y6ChI11T8jFz49qq5JF146U8ZVeaP/TZRmH3XEBaWiWJaGBfL6aN8
YIIORpvnumdDQl30S//2w2knGJtwpKum8v8PLzX0yODIjZGN9uVMBwr4B/gx4cXiaoI1KggH4K9N
YXUAaVI/oFxH6Q52mMaEZpz8DzlKE909RrWOl6MXlgco0AIdp4Fy6X0EJmpL07AYAfuqvdPLvSr6
fT+fmQMuxnWWMwylyVsv+1bRBe/DH2gGDA0Hj+xcj/JpBDtSJRZsaWZHR0EiGOB0j6a9xysYguNa
02RE+SWyWlCpYeJiBhOGpkAzm3jpGTLuW5iN/kHFLHkIxZSIm561Q/a/PQfMox4xb3Cp+oVCi2Ym
dVZk85YlAW1QDiaSGcrTYHrkyQnJMZw3boGwXfbWT2wENxRoakqKhB7djmD9H7rb6bVkL14zoT23
e9udijCXvMhGZaCc8Cc1h7pr/wtOJI7OGMsuGV9jZORtdHreQPHJ1KEwPg90vQgWa+3R5Nu2fZWO
eJ+kiXCapY6nUXaz2d9kAsE0zGhf3fkExCcvIa0hqcw1HnAoyUW1WUgR9z62RIL86mQO2vpcNity
Rcmp8eXZyGD14KagwvfL52AwQK7NHI82CBkbB6m2EP/Q1SgHUckMDYc/LDgsxqffdBGrcWU2D3AZ
HKTuzWahyWyMJ33d63ydC/3Fm4z3D+yRr/77DuVfyFni5PREUX7nlxFTBpEAXVMyrkN5Ds5VznaZ
Q8yn4muREHP1CsX6ABSFpeUWDd2Ya2fEC7uf54Kk4JIbPefPZMVZjif3GjJGTXx57FMkScCsfMfG
p20YaJXKcCaZNNCNipZnRgdXYCg1Qx+CYU8lLzUG/XXnjXAdtuQGEvwC8DhRYknmD43XjyYtay8+
Q9NB+sN4W4CL7/+vhsrTRD9yx6ZIU4S6I1wbbSZTw/KR5JNl4G7ApMoZBwI5vBspTYNoYDhGfwFP
Q5SuuIKgEi0jd79E2n77MBVKuY+w3ttE4OKg6xD9ZDMFaa7im7QvdndqzRr+sj4/8eyQykW3fo2D
QiRiBk5vgloSI7vUrxcKsHR4SqRSoZWKDZ75+ejqVcxA6TdtAJc/SmvLrggYIBOuIQ/xwkDQvMYZ
paw34iVFAGh4d4mZo8LoCsa1qawcDnHX4s2TBa3WWBNNywM67f890yB+Mwz6Zq7/pLOX84UXwa64
dHxwdkNFS3ERuH9WVk5+wBWyLl2cuJF0mo47F3Ys28XMWRBjCS7kJNOEh1rrLRVUqmo05ZYLjbEO
QvmcePpVhOuyUqDOiERzbm4zHbBJI9hz9aFqZzVJWD0BIRIhxRiXS5tNuWkl7c/PfzPxHPIKCigk
z7ocFDnGYPzXghmzwRlpFTWsliLF3Tk4/qBs+ZaXH9SU2rGj+z42kcX33cyxoNo7rCmfGcRmeNSE
M1jWxvuCxMp7+L0OG3oTwJ0+lQ5THczflFdBVZf5S3nQDTuypjL/YUbdJvJds7cJBxL2fSrQhbtV
zIth/n1562z0uRl54qMSyedAvRSIYcals78+iGIZoPB07J1JPOyJb4H4u+D1KmW+72G42x9/qZPo
suhS9iMpdnantALxEtxNsB5vgs19ub743lKlDKlqsNWUfTP0XUY7pB+F/Z1EYEPP8d5qd1zA4YdZ
ExkwKvKoYoqo4At458qF1Nkfw5PUxZPKIPKu59dfhj7JfOukigRGT20SB6Hhg0VJuDUjaxnAj2wj
xk7Bf21D/H/dUN7kc6hQTUF4rHHgZqUn7VCIhZfSOPYD3nIMGgcwATWeJX3jG50fM5cIEvGlAKjr
pWIQBW3lYg0GPIB90PcsgsEX40FKZVgGITePj2emrkCTvXDuNLglqdI3dPOSx2Xhlwp8G5orNKR9
BVRcbb4AO8VP1nxJcjRi5B8ONvqWs+2NzluRmjO3UH5MqXW6eDLaAbLeg2Bq3H5BdJce1+CQxFhf
F79gp4qziriXm88rTy9rBsR6OQLzxH4MA9DkHiMXhG/QwWzPysWsZ0ze1cgO0iM93IoWtEMsfQ0R
ZH3ynJXvd9nGiUx0sXhMEUdZoBduZXNjozodDrDgyBdiGuIvQ1Oh1qZLSpw/EkXqVaznOzrI+fhl
XdKxEm/sUnE/cO1ds1MJMS5C8bf5TE4wFyn4xKViQiykGzUB4IL7MZJ3J3TAHbuHMydBv4yVdBTX
1cGPQQldGOqdgDA6n0Hkn1SnS/EIWJzq6f69sUiaXvcAYrMgflluqGMCerPpR5AKDb5DTd/MdAJU
kNAZRPx9AqW0BJ7l2jSuJzHYIZe1GuO1x9dgKxF1LVq6uDLMnRm5lsSRRBDJHGwReGFEm5TWE7sU
ZnOk+w+oZfcUgiCPRKxhK1mSqSwdIs0NmtcNvSnAo+3HvT2yvlvXMKLjo3O21NKWIgcMyGFCRsiE
sSN+HUr6JYCrbAWWxSHjzE/97S+yGzjXpAT6sUCsZdN15zr+ZnO/re+FCUJP8GCwUVf7Fq118iY1
+CVUi9nlbFVllf2J03SzOmo6uD6fVqBEMM+tUINju0V+/eBk4ZRzTgY4fZ3odnHbKow5rFQaUaAp
mwI4WDvbNdPw2WYR+fqg1rWq/sOd/syMjH+pvYI1w9NWHbHeqD4KfUPY4+3eNgsVxm0/R6niNXjm
srSuObey4vNqBB3gPvcZauO80TYxB7mm2OXYHHHXOUn1cJvi8Ko92CHyCyfsdNLTpxzTMwQe/oH9
CP2vlPhBUXyrueggIAWESNT/jbr0pJ036sxlg0fSyKmssVW1aDlqt46LN7wMlEgn2j6RQx1zly8k
8hR10ba0pbybt6vo7BmBZU7uUjyV4IGjJeLT1kY91xYBf6ESpLrCokt5iJWBVP3U17BysJi1PJ33
brb55HIRECeTN9dj3c12IrBhX6owdHVB+MIjEwX+9D0Egv+XYOu5+KqXsOg1GOHWA0msMVZhjGmo
wFyepuF2oMY0i6Pzf+zxa4UyJwc6S1Pp1z90mR2715CBjMGL1A6zNSM+nBfyyvCPlh5wwpuaWjr4
45rZpYwd4pPwcHwBOZFkBTBpmTo9hQhF0J7BD5c+oYGRa+gfd3BkHISryl70axYBoQKyinwFgr43
qO0Pw3PVsJRFCbd91kfteIbQHhCaSCyZbL7t/YQrAPWKKaUCQ5nNzswLfYR14de+rDKn0ZEgaB8x
JrFm5zYcRIYiECe2DgBbjI/7l5dKpM4Xtns7oCuGt4AnjXXAgXvBH8aDQJOzgV2WR2CSANchMWwR
J9lJTf97c0JWO4QB9fWOodiEoGRu/y34bQXnCmjDG9H+U0arGbqPtU38RgVL7DRkuR/QiY4joiux
d5g3zqFsJ0pgSKQYGwTOpCT+/xFofAHup02pzFWXSRIivgGwcWjy/y85Xq8m67jUIBEa2xwoA65j
cZ3myRD3R4gTAWOSTZ8sZs7vPiOI5HD9Qn6K7CVDMc8W+/14dhf/oNs84j5AgpW4LSHulbH+mglW
mrP/ccY1C+R0LoOk1DKuKW0NCN7+eqFDORkvG73XoY+2YhMxwrUK1ZPonZj6xG9QRrf4w8BzrPZq
qsww7roGCH4wLc7tFR5oTyh2xjQkzISKi4yRBuRlUfxUBkXj+FPb5ute+dhEc4Nqb4ZGKSYo8gqU
XMGWaG7gqVKUUj9ZeDViVvmDRNuH4+d7FoXbqKzTocKlLQelxf/hEZuSxWo4vWyCaGrP5jUdCDXg
JBU3QXtzUdxfdcQlnEzPEhtmJOglLt1nG8KKLr/LNAvRw6YFmVDvFc3ZKdccl1vhhQGg+VBIh5YH
+1MF+bEvTpy745/hPB6XNO3LLqgrhrOM02KPwQSC+aXkrXmuU7ST6jt/yVXVIqYQYev9HGbj/iO2
2s4z/b6xVw7Io6rhTKJVtfP3PfH9oW3nLFnFGFoZbwaMjVtaS3ek5jEXg3ap8o66vhtQrCMUvPe1
a28wyKnLLnrBmbPlWJ0ZTL6MJn2+gIk6JLjkydXzjVYqWG3uLNH1LxcaXxTA2FOiF8JfSUN9OFRX
1fkLxeF8fQefeBvRxLNdMNrZnd+6zQihvWuJZ1KRNw/o28jTqvAqFIxbzs2tgjmaovHbYRHe2T4D
UNgr9tKZMWydWytFc3VvbcEVYUgGVZX6eZ6PwQt/65dqV4gDB3KCQBKpBOipIozA+KEdj6tNOquT
NKyei7EBhBl1fphoEaDNyfDvk1CTKpFb2Xw+UKFo0KEVNV9Yp61dXU6k3ZswD3daVowtRRLmiUzW
Bx9ukgR/+JC3IX3NXXK+oChwHTdKtIy7qaYY2mnGPjCYZpNyL572D1rsBTSwP3QRQ3Vr0Sh3ANy7
whUm6NqOzxzIFrOqi1208xGPcUABP8YBB6GfZBXplpGMpe/d14vmd+Kzlm0Jg/SLA8xfTKI36tjo
cwOgNAnb2iqJRR+/GRzcUEWcQ/gTHgRRGMYnQu0XXpOvPAa/JtI2FaTNH9nFN1PmbCSQ2hjIYUeA
gNosqpqly979MkhJkZL0dZzIL4TdjVbkHk0Yd7VqtpAHe98dM4OyFMYi33ussB9JlyR5ajyvwvSY
pL1N5VBNZUmPr/4KEaU/RisgC95ucDZ7QAa0CLuttpgOlN4tELsInLx9A3h/IiNiTw7M4eFav/nr
hD01nQvtZ+u74QkMYntYVpxNE/6BnY6NUfGZ/yfPa5qqLPC/38rfeVMd3ulUdW7/KNFSmRM7qKYc
MKfnfZUHAY0W40jF/cw9SxjF8NbRnRRMMGDgYu+3BIAv87Is3ZKS89gWstm1Qa+O78nLv6vdFlfQ
NfRg7gXVuPb62QjVbfLw39tnWGHarRuK0UuzU6VaPbXtBbGfO3WV0q5TxLlP6Pp+yUYi2PJPFuQX
HUr2kuS6dDmS/IyqpY2xsHVpmgWwzalWRJd6QAQUFmgaSmPjSaC6jGMkXe+LpXjE6fEAq7Num11d
hBBu0O/J0wzruhFO0uIxrxsmpYrqSsR4L0fn42qlLp+KweAe5aMwc426dF5PWn45GdzTmjkbAS5A
TFzMopXGHfmKm8O0eHkPB55/UZRx5pkesYZYSsBuvlps3S+473z0c0uYmbkt9zULygj+jqFe/16M
pEvwmobfHC7SkPZkIV6vsgT7HGSQ5sTZxHamfvvQAn6RuPKtXZ59ugXxHk5Czb2vW8RqxTHGRGaB
KLAXa7jhASopiGprAEl3NVSlU98WocMETeGR+epaaxbz69kMx8qYfMlkDjPN2O43YdYm9WFf7+zv
Jf5ayzMM5z5IydHrBXBsjTJYiTb7DK5RStj8utn8qVHskS9fC811cgW76zPc0hXcmL+voa9Idjtp
eYv1EdGK1cAwEHd9tu8+MbPNJoLY/ZqEGWiNXymWzkxUV2Y5k000BMKtdQ/lyPJBFzbHyZKdPrWp
lw17fImqn8TPFHXeX9lmot/dFBXisXtP0NN8Yhr2c1NKYycXZCENq7XlToHe9jFTzecqbdYSs2s+
TIYbYKxKdnMuySQ9VLTJtwIWoHfk4p1yWvte1hBzDxjXnphIt+kGnNmFbi2B0vp6zzaBRo4PQyKN
MHqUKSC168YEEjVRr5TpsrgOSVVx2icqxG5PJN59IAX4tEJTCrl8hDn1B/aD6NGfMOVvpuJbfU00
yLLe/28hJ72eIPcIMh86V4NJYikP0I7SMA/gZVXMFLKKE1uyQcuDdrWwh2kzUtAMqH04eZuE7cLC
kQ5Z+wicWuJgFnZpV19ESDv2LiK8vS5331wiVJWuaN0H0Lb8TwYRZEvkRFAuttfilywVqg6CrQYJ
RjxfARIZZcjphujfn5PGeDTOyMrYsfpqm7zYn/38SCJPDk0ev9o242WrOAV7wLw7KiT5aHJDh4Bu
UqTzltTHVp+PRfhM3HJQCNTFq3w5b6xNG7mAG9dXc8CpiVRKlTxVDGYYyksWdJqoO9xM4WuyiMMr
OCwS08afaQtS5BzD7xgwWEtF8cLGOOSoLrP8cU+ulua8PDbEBxZyS4C2e6TuEJrz2qbqcb8D7343
6LXyW5eL9XB7pBasScezt+NrryYLzmoD9WJCZwjw43iA0I2q+znfarfGdasn9jyTXRkb8R82AYN1
gOpzA46HdiEslkETS6M5eAIEMkcB38/2yZz1jFYgIDMY41soQM2xqXyR2dXUMskQ2tezktxRQs3F
jl6HhZRBUK+adriKP3tlmusuI6hgI4yitjrqR8QIMj3NtgDOguOo03uLUgdLICm5GCwjNEN9UpTy
4RMqLUYzaquQQzfXjgoqhJmL8Dhz0uOSSgqYtM8clSK6rYZZcYY+ZDlA2IKqiKs12NSl+xYESZAK
9JcnH1pj9TtGil1z0XDoK5SJfHh5G2JegkFA9OsckfODTTzzr1nqzXGp4DnBa5aMS+tMv1UreCP8
7WcgUhSyI18DzH0MbyBCEpIlDBdhx0XoLs4A+i6D+CCG+XYEDyODpSM54ORKpQNZjHqTE0qO38Fn
bc5rb2jekKZV1dYhe9n904PjA2/uIVij0bSIm2WvI3kT+OulOyqkppgkhJ9g15SogTUY+ftvg+E5
sGp+Z0PMbKspOHEeJUmQSIiEOqIvitN7pj+vjXRouD2/jxFhp2VruEMBJM4wSJ2cxLRrhL8ux/mC
dGJ4d5i1RGElOp3QxdIe2d0oF0gLukMSmiKwo2YwUOgvLLcI5snXFfr9ChTKbAEZ6hiEIpnOLR20
w8R+LX4KQfRdrRlRFbN2ljUwYgpUbd84wTJfRV84toJBMgOsB2Y/VHvQFfN8I9ekOrRMdQgpD1Gz
WPqKfCQScNRYCs435T2CPnp/UKqP3PjCC3eAbxEYAqUS7UyRXU9226kETCS9UxbdOijN+TmaIQEi
NrFbdbvF1/mgbRwDR6lrs9e3qoGMF0pA38q460I+r8jABudfk3QIh1N8rcJySTRSN3gVBPzofMgK
AJILMCmd0ny/evYBTv8SygVYaECcfBW9R7hCPOkqR2QqzYP6y03sYlrSbVUodjqBoQVm+VVxPheF
woZNaPDlZ0rVlETKGhk+lH6dTt9XApWN0U5emYl87FfR74Rp42eZ/g3MB0Mz2zFj2kCA/DUV3XRg
RyFFFmsXiduKJImapJzVmHd192fmc82yMxc03gahdnKPSRh0Rt+1GF+rFf5zLltBaqpu2zWueQ9X
2jbfQnaBGaBT0jAJV48H65ijftE+OoQ+HSIvRjTxFUc8XngwnlLQDCS4Qi1JRmfh3u+DyXbK2F31
JasgI3h8fhbfrexs3x3Styekrf0oeGByM0IM0EI77FTYcnPcfr+QNGcaKkU0Z8YXggL/kwypV7uU
5KQad8PTvaQxRDhLg0gbDYZ9ki5WRvXHmMPksbcSUIjmSRYs3pCapOmxoN6AG89vTgBQhqVPExb5
66GxtSOF52fKvjCnfelLHvoXWe8Et9c4C96f+qxDMjFCJYo/VCzBb5fdz9J0+sxI3Y3b+g8JG7Qz
P6CUaaTYK6Dze+ww/6XHSiqluz1Ik93t6tdhBVIF4D4jq9Hko2UcKNvu8arE6gny38Qe+/rgSOXA
LTLcmTI8uVST+rTxq9gp9a8bW7m2HgzybjqNgK4d5NEtNLNIx/Nmfj3FLC84YYNuz4/MW30ps/QO
nUAVqQxXpIYmTTtwalsQHMFK/EI9pjwkuD5x+krirRMZ/9qVrTqHWZDdGdxyNuF3F5Z3P5Qwotnp
z6srD4+7YxbysiqqkeCbm+pq5pw8c8rMyWYZiVbVT83eAvHDG45kEwoIENIX3vYNB8DqdEfpyDhn
1b/aoMEFWEdGZV0DRYdDmaFuthRDQArN6UccUA/yZ3GlnJDJf3slIkOOVIhAtIAIJgBpDIrstAOk
I87Q1BOB5opsd96mr5UL2Bl6nossrv3XYVFrs0lLfcbSLZzGtlfwgJnzhVsA9/D5V6azYv5o7W1G
GQBS/wNKdLHyjiyvQMlC/mhyr0U4SXQnMgbdIR9BAH3aitxEoeSLy/TqvgVNntAxb3c0AYeONV8+
uINnQilnYRIyE7/Eilo1fQNFprxivZi8FFvsjP2Cd+lYJTI6N1eLyP0ZFLe9wY8N1JdZkP6tTKat
1c/HD9RKZRazj5PkX3tp5+bUkknEULXrHR+RBiH7FG873S40340l8jcyCy1tLqpSyS3YFQzlbor/
FMN16wat8oYuSYOf17uifnLYNZaH1F/GpRSXbp8CYdErcx8f9R+WER4OkKCq5xX9p7S5Jhiid5GW
VsmogrPPVfMMhx6XJ2PWKlQLqqwiDo9wcC/jR8TObg+JS1HE6JBdYJvOSn9RNxTrJwqoM2+/Fbr9
Qhcr95agxy7zGwjvpMGnqloWrRcidamzn+aNbBzm48CmyxCVLFNRmAT01VXlA5iX2hZAGRnwKDA/
RdD2vE42yna7k0+V1vks1KzqKNv+W/mxL1bP+Ie44bN1TWUN4Dc785lf6Qlwwo5wtUxIg53KZLdW
viITRje7p14AhNadWIVHDx4A6WW292aCz+qP6cjTmSk3oFNS0+Ds1+vbIH7yFh5fzp9LaljpYSMl
r75itYTjVrlrsOCWhxEo0k5ao9sLONotAin8ldZ/8+3R7amyZDWIpV55iC8UMt8Q1dxA4yKmnzZA
6sqtQpz7PKMm9/pmo/Vfye0qEKY7ZOPnImYVceRqGl7fNH/ISlc+5NdmykQF6Z5AYquOT5FE4bMx
Ddd3b8JKB1GZXyz4AKY441eI967+1PrBbGVBz5fQnWC0wzk4uYxpg/oJtSk096shgdq9QiEj5yYK
ZNJQ/dAFBhNaw2X1ZZ4h0pQqdlYGgv3bxS3XKhmDeuO5uVIoP9jPnLM8+78FR4EF7Fzk9vWfOoCw
YWPLMI8hLXT+4b/QbFJZABFzYr5qj9xA9L2yZPfPBcwWMv8an07zu5c5fR1QWENh2Zelw+w/nOxp
qRKZcsPGU/7uu9PTjHUhisJbBd6sS32f25Vr3jkoOpetXgf6W/qD7hyGkJ5OuAj6XYnNfbk9yuOx
O3ioBOKr3qdAgFLTk8VFSM1gC201nGVEYxujfrVnxParmQJgQFi9IHswECtIG9doRR6stoIWDBxg
ONca6iQrWbX8QOBXg4c5C7Q4Yrdr2YEDTq6DO27M5NXYZHQnGAxAoYI60O6/f1L/Z/QgVxo8Z1oD
P1gGG5gm1aOqjSPXLqkH4M/ZWZ4XlR6W1AR7XqlE/3h1IrA4uFa6DCkjq9Q2KXPESTFRVFTLVnT1
WXCJVQQhVYzmqsSS2oBQcLBiUdYd0fUsIyuuw9lrIUoGIEbbfdPJnh6Q+v9/uwfqNxWOWUt7ceLc
Xgw4ESHNgVQfIjQdc7sJeYxS0IYqmqrQEdBceOG2blOVIr/JSerGsSr9FKaLidJMDIg7mOHyykWr
n1fXGkzRSmfoGxht+rpZeUIkKh8AlPEzli9j/BW4MZdkjEfVlXgsoKYAVCWMu5XzoKYw/o30DHYG
857idDWxuMeTW2GRBWsRUFmezUjFqTk/Ej5qd8DowuNdoDgjNJJumpoS/2XFbwb/ZJZf+cbwp4MS
NCyfDq/2oWd+iQcoaHXMAJWc/ooY1mWw1I7GxP9QgDZEFEWG8k5p4jQTalIVkYAHhP3M3P1itdwY
AvedJz6NTlEu4b21PxrB++VYLPAmlWwotPh+8F5lej0aRhSmiV3QYEq6TbjJiOBZIp57nAYl+Lf0
uaQZejFebCYyXSMZOkfAPqpylNII2LeHVLUBIzlK9YwncX33eSjwt3BEj6WciZqhKsWv8lxpPd/C
7JUcLuvWuF0jfW/WpqTCFEn3Ru6BA1tkNXNkXghd47KryX3GPX2s3vzuK6Y0Mv1e6U++V26jU2FQ
bxv4yKvJD4PREgAcWF/YpzKZJ8yYGNo4FgHMhVTEicnqomKvW72Eigkl0BUFoKDSLfQFnLYpfOF7
spTMfdLFc59tLcSq76cYWcxBURQ1nvyiu0lY12UxdXoN7A0pJUOhEV9kkmtSILBz9xNlMN7qnpjX
uK/S9vzHLSdhrBp2MxSLyzzJ6/tKHZodc2P6Hzycd/DnpN6lypgJNSRJVPRghC0mWefI5/WxJ7Is
yPjUR9AzSAQ4h3AiBxACReLesBhQvn9WdrKpZkSEvf0J4EEM09RBpY6K/Zm/n+KbaoKwRx3DbP+o
rOhCPKVPZO9E0vvsytQH15VDiC2+5iPaZhopvLLJaOj+sSr67i9Woh/NAIc7F5JEudWtyheXMdPh
oENFQ2hh48yjd7PLxAbEtr0NLqkBd46qIsVPu/qGPh+/cxt2TEB/ajQrP03Vh6gaKZl3PTfImikI
WIh63fq1/s57lhMKQmTBE+XUrmSxgsAXtxpG7GZX3kv9iQN9kFswrWuJLAxHPE/S/IYz1EYfeN9G
rkaONeL343u/swbdzKBBDgkvohwqI4eu3ElsiCZJPe+w8ek//WVYXHowdX4tKAxoeUv/VUeilbZe
/5NYN4U1f8ekzGUmBnjgiP/Us9LVmttJFd8OTM0+1JSiLyeJthr2oQcPVwOnI+oWlhbTWv3gDseN
0dBrpWWw9BwGeZHHmNl1Ahl1JY9yvgEKjfARhvp0t32jKcJYgKtJxdtbUmcSutq3hThEr/Tc0Qds
UWUMEXjOJHQI6X5CPCsnYlYCMfywtgWxcGfjL9u5vwMTQkWUn812VvGfi5zL5aAChue8efC53+0L
U6IrhaVhx5cZ3hTVO+HKr9hQFOKFWmDuktg11OniIi8+6Mcl3UvC6dzFdopJmvHgA5T43B+GNIXd
kZNvXeq3X1MOamjqHQnZNKqJ3HwWaSku/FIbCgk9KXoaKyX/dOEH6UYwRvcK1nqEFx0xTKUBHe0x
v1zwSwJsAv/pX4rkAje9J+dZ/26/9rmh/kdyAoGwR3Hv1psur7bvqILtUPLpbfCQJmxzVEZxB9a+
XPOpw7GZSk8bUDg+we7vcJIBn7Fe4Dkk1N5B/g4+QLvjVQnWa196yPH9BY0DbO+EVb+wbZWoBQK2
DNA7vvHFb3V9p57tLGAV607r+EgmxcVVrVoIcQ6m3OTUsqexIxKaXsb/OyoYL30jq86jTw89wZGv
YTpvA/YQS6pjC30ou9GK69BXnvENp4FP2ggeQBoYjpqWfK34edGF1eO+DZf1Sqp3gtBvDwW8lpkT
m5Py4TQGFOtp7xfWIAcJeK65Qn11nI6DihBoFX+KA70NNq3W8h0EfIPOHQ+pANNTCx4OQhkzbOoI
GF3Lz0zb6aIvkhZiAA0iTxuwuxBtX3vzzXYpND6vG3/06cPL+mbLTR3DIdgkkEl0+1FsLo7GmJqD
ATqtetvgDNPDM4eRRXtj4Zp1GXjX/bMfHVAnCvSok0RibyDXpckSmFAYkqm0VxI1JRAwQv5+odCb
n1oFsy+1MnJKD9CtFPuIB2SlB1TT/c6PE8rGtHQCbumwOF6wbP6PvkzRi1g2wdwxNnR1s4Rp+/9A
oR59s5BSU0ha5dFlElUOoCtzQnT7aCN+B+ph3p6WVeWXnTVxnK/fWwrxGV89SHPTDvWQjw7NSfhu
io1NCnGWoCIJ7mu9P2sgwPoYAyTfFHnC8EJn0CmU0FrB9stwA6JR30PchGgirPrGM3WAKcN3U/Ga
bOdk5B7RVAqEECyLlyziQpFdez5jtAWEpBh0z7c07YDCmYlDDmKBlLacYzLIzNqSIPvD8wjNlfFu
u/MMCvDlI2raUoH9UI2MLirHvtiixBEgnR36bDrLOqFQgoS0irwiGLEcZRdLSD1JMylUC2JhWMoU
DCOYOAigZ3/lqrm2NREQ4aJ9gBzOvyWGTfkZZqdQzA9Uky5vGOxamJGaRA7z44nLryHD1vdINGKu
NKdCySXYReGglUwvdAnml/qUW28swWrY0z6qOdrBOeI670sX+aMEOX8AUkpep0x06OLwuYByUmtR
GWxQEjFrcn3DGWjM/IVraSkVQ/U5ZB7p6m8o/fBLQOtO0voHFg/wkoadMgqYYQkCwO6tkSq5zjmf
3dUn6A65r/b2f1BStoyTmmTMdIByV2EUeiRT1xtO6KuMggPtLyqkLeV60vFSKwTF4kvQ5KGd8RXu
2dusxSG+WEyL3ZBrWhChgUg010T9x7h+Zyii8h3sTsW4KiQx6qK2B5wtsJ1NcNNsIuIrG6ocWOvv
c59YWzMVwxFqhYjK0UxJcrkT5YAhIAbJucOkP728GGvKrrnPOiyh/ooYFroCen9A1W2Ipe5jR7bC
mm2Hsu7h1bxsdW51aSkEK4Xt6D/QE8Y7HBq4wkEJNLD/3BETrFWJkI6Z29nf7luT8J2UieeF/3w0
kK4srRycBHJKJG9+1xt6fq6wzZ7uj3LcbHvjQKU1N0l9T5QOxvNDawGslj+qxJPd1z7KPBuidUmt
zCfFwbz6ovgxVFl+u5ZwSXEYw98tlcGidv0AC5kjx5EkDQVQLtGLNkhIH5NE3+XocbXLy7xDB2qj
k5M2KzI4oRIpAcq9P6xq2riPSmHOGq28EMJHFArjFomLp8xfPYW/RUAfAAOuQXGZrjGCg4xmMuY+
mIn0OHgtMnMo27LwQCDpayKtdSV069owR3cmRb6YQZxEoG4IV7VPr+xEr3QvHBTcx6aVSVY/qFBF
eKyA82INCOo1DJYfIhh6bC/NEgzK2ui1ILnbAX2R8qytp7ten/xANc695+dXpN8sIaNICmtuZ/I/
etZLM1bubWFuB7FTP1ohTGyrIngSHRMPD7Ux2TUTXQJOGvz35APjYICdDvnhIhbkGp/aQFgN1KrE
yttmWEi0C/Ed+7dssxa4iyDcrn5NyAwHqMVSYWyz/fgDx3dbNCky8PeVq6JdEleoc9ya82JVu5i/
2mMJyH9rGCPFgc8MCtgstcPTF3Yj3UK8pTM4pPnzaBrhGnnG4sOWnpYs0qfJwloDYanTMk9CBMMj
qbstbZmeB8GmHc19vorh4ZJafKuG8lFlWTuluFDofaTAKNwU1P5FjjMsoVEUuL5AHbu2rKyRy96l
Iu1J5quPPyDrhdEAgW9K2nGXOrVUYjcr8aR+WoHdJMhL+W4DADuFpIuw+JfY2GiH1jyeO5d+HtNE
GKpaRTEje3z83XypSDtJhefWRJIt0qlZIDGAZl3q1w4byGFqgoInbf+hxKIpXkVCMbpawZCqoqar
Iw3+/XkTnPFyEoyyDR5jaUSXPpBjpu0fW5jtOyi7j6z8xEG+sUxhADHShVtTzmvCVJZAroKJdSBR
IjIEKVu/R338UbLrAAW9/+Msu7BCxiZ5WRaXz9jWZdMRlwJqJxTLCnZy9VbYCivYnpGdrUWDyQc6
AlaXnIXiZy1yUerZgwt9lCZFj7xTzsVyrCPHETuN9UUd0wFKSx1k/1E/1gyqUWMJcr4XgVZqMVbC
i1/pWPKTaIIZE9fbO/pymvGaKtUnFuFsKviVPxFdVVaO1UYNE6GId8gtOw4IhuazD9geJWDKqULT
E1hPd9NwXIOCMwM+3CCg2siujaSTP9YDwrK/1IEzoit95Iqyc+1YlHiMAbj6jLi+V3saABzg5aiV
nXucblNWg/ARd7URD/p809wvLBlF0R0KVtb4YP6pLS2FOTAZd06mOq+iMfIje7P/Z2CitRB4fa4s
hR+2JDDxjQl0LKHWyv7/UjoFLNxpg8G9iedhRb3Su7LLFuAM1iFMO7ZlhW9hrKQPuzHez370Dh/X
LI7xjZL2mIXF0frdjNlSofQlmv0/gebHqQQVP4YiexYKrtLxqjRrobzG4JoSSS99FlYKlL5fvJVX
uuv5NOuymbpA3V/NyNvgK0n08FoFannXD4KS3PxRI3Qgd6SBUmYvNzog3YfPPJbo3WAsV2Rj5Wou
OYh+94uL2OCvFb6MpADCGO9IzNLrXT5hZvTIE/rd+ZT0GgomIlDwWcQCve23YiQMHGNRrXVngAC0
XZ1yzxx6lgdxzUdnGBa7pm6BuYFicVKxllXUi1uKnF0HYq6ktSfG7XTS4gSQW39sDLRnavbnis+2
Oj5v/1dYFhTyY7WhHLGE9Ajss0AnnkBe70w1Cie62wRaKJPGJOaSOfwofVBpvOxPODRRt5456D2I
Agw68HTr8tEn79kGFoLMp7GVGanlQjRgTS8yz3kYUdHFc1s03K1I3sfLAhnSPrrZG2sl79nYxnaX
2V790+oIczXVeuf1TnR3gkZRty9IhqTZJXeI5eUBJOqvqGLNQ1JSdtCh4w6pZo7pS5oFnZ3LA5QK
5AxVvpdAdBVSjXFxDqz6lcXdLeC3vOJz4N8XPgX4i9vLOiUmJSGlXd/kNgbvb4zoIzXJMN6Qt1t9
ux22DPyTsEMwczE+UvDKf/9NbWMa0lY9D58NGCC8M9kuOX65MNzY7GUYKHysIZVFbCpED9/I0Kps
t/LDLbE5dlY6mgaxxTArAx2tepDlSpIp/l0NLfBBpF73ty6o2mD9iFJBPPAk8052pAwrQMrkZadT
Ho94F4ruYRMHdJSfpSOTumxvrhL3fISrXzwT/RFz7v0UoXkbgNfov7PjgwkuR+goJQThg6N+d2oX
smm1QvZQuopHbICM9LgtFZ36jlsvRoz06BE14Vktt/E5WVJtanaaRaD2t3WkyKskV9eHbGSMalCl
ro+82EXVdClaGbdvr8fh9HNN4io4LWi3JP7ieOE2o3UDcKdzVW0V4jemnxvOrOl7VZO+z4rJ26rA
rJx0EcNn7vBwnxKMdJe76UtGgqyblQdpyVyyt2x2ufTn2IQf7hbF4vN7mg0SPSkC80S0JauJQQF8
Usqw2rkBBOqQ0Pzf+v8h4H9iPdOOcyMnJ2eC0BQ0d+ZYHLRuIU4xAaP6jRQjwLVF+h80py0GjUJj
2BeWu8pF+yi/daAbqvdOe/WCWTjIstw+Ugw+BXnQGGktRWv9lD7S+euGAC3hxeU0x8E7TQLe18f+
Lm+b2jXaM0D1BJ6p130gzpGqCUl22qb6V8rHAGAF73S1iJxIaPiOVgWUqTCtVKBsPNziDHDE1i/F
FZ61lJrHlcKLnrdjsmAhIXxao0TzpFcr7P5gBoPeDsgTE1nbX+Z1116fGatItdU2bcLgzQZV2A+B
6FD7/h1UAuwspRI/ugsVQ5C9xi8U2/6DnXXNCse2fVWWhe2EaLrslMMSblNF1NQEoqBqRCn25Dou
6ApC2xRhANq6hDFQINCEiIqnxdTwxqcjXRAQoo6Im245Qu8QEzpCV8raqAqruYgzxgRHDuu+3nWf
6KiqShz+jqc4QMlFrRuQxUavLFWiztA/UPq7GnXqYOju02wsyCbZNcKFP44WlkpvcNKickckyKTE
GV2v1nzQOuqyEphtBkVlciOTu+vJQgeZr3GxDO0pLfOGf28W3bE2enH+3lU7+oUsacYsg3w+rb8o
iG1ytiijb/PkPXvWEpRsnQl7+bPJH5LJBkNfOfn5TGbNcK+TeSfa1EPafTKzq4t3Eyj1395bSdYQ
E/P63yW7GhVUVVbHU3Ciq6yWx8x9EE/tqvlkTTjMjeFr+72V1+hc4KEDIZQpEv2Fk7n++jn+j0lh
Ubu4QDjxO/L245jN5T9102AnJxKEc+a+nDoGR3hYDXl/AUkAiMO2ruqtISi5DtMIsEBkeHchxPjc
AQ0UG+Jjzp/M1ru1xA8ssxI4kmtQTaebXRLllAJKv5UGKuMbcoBBJ3RCmWe/+qIe4YlKmzmGhYAk
llYq3SpG/hff6LnZAHWhvfDPgMAWVGNQKB2SH10sUfT18CUx8U3O2/i6cX6s2UrQ52DpApo2rywY
Zx4HUp4YkNxsjaez+CoHs4D3Si3zmrpU/Fbr3jG3UZ0iwhca30xXlEr8EWE7swaeOdoXcmq8D+RM
3iV42QCEDH638k5+qqcq2zfKcTvhlwvfnH82eyjTTWfqnvY858jrUy+k3IA1blKuAe5mcjnh1lgt
Zd9ayYCwVr8vreV3gcZs5uFnWphLDiX3Pf/ecHzvq1LlmbPqdDfuT7emrOvlOc5er9fgGl5jpURz
XHcYl1ry9UacnXkodHgpuhIOdN8u/jbFmFMlsYyYQvrEa9HI1SPaA8tEzZRp5/NpDKxx6vNkDSLw
g1qkGj1ARefo0B12iZ/gWzM9HgzM+nKUBT/k0n8ETOgxmUfZzWFnaiOze8QHij0V5nFGzAYkX20G
SsaYEJT0jKtjcuBr2pLW5e42IivpCoEt2qKjCQvqx+3J0Iow53DEg0L7gAL3tIkzcwdZykZLGNWB
AENrLojWayxQZjR70/2VIgmoOyfG7vhz70z7K3IASMtpElQOQ78ElvvkHeez4TWGeYZqpqQHUNO9
TPfQqwcW5Nl55bydjxVGX7COzlP9Mcf0JPowdEkBgvE3kDBdbYQM+ZZUcjxXgE43bHWzz1dJTJkW
lRz4sfdzfcrKzkMuTHInM2BcsH/jCYWUr61/Or0s81jhcr284xwBlWDf4vIMF6vJGKGQmrUfu5lc
59XCUk0nmNpRQkqgTHBH4N38GjPGGnNnwmXyQZsoUPhv9Ex5hkiLKOXc9x+nY8bRIT/f+vvPdHMV
6VBnzNrL9hzY9WyMr5/tnQHuBNLk4rsNHRhAuKKq6zNViQeX2pudRPHBqgbnwRXT6IzABLu3xcHl
nmnYd6ftSjXyWverglbi7BokHVS81u7s1hTlHxhP5ra2g1gYZbo/JBEeYhdb1n5Es7N4krL3HoGz
KE5mufsutUw4Xo/JTI7rG8pj6uqAJK96TPqllFeYRxhGlDgzOjGsLx6CFH2XyM9DyXwnecelxpWN
pAyUlnvdOUX8WoOLw4FoqJif7SIKUWNx4Ct7XRYwg48o/2pMpNjgg/SHzSC8pVv5pwf3L5GEXifs
ljz+KrqVjDWoogeaclGJOAQc8v4C3hRiKCt1bfqmpHeYJ3gbhDXS44xRAe+IUNYIG4sHSAr90+sB
4pRdCvak5CHH5QsgZ3Fu2zRrrpt3yyhWjTOvIUXg6idVDnb2BS9x4cnLFKhmxpf98NLtjePwji/3
NjPyqQQ7I9mUVtHkE/1fp0MjhNcxqPOZOZakgAnob+LfHz/QMF/heiiq4QLsN/WQToqtuC1Jt3PL
eGNXqRwUbIlOPjBs8dKDHl5aI8HYx0MPFC47LfrNIyRsGsYgiE6Qd8i64AK5FYMjg+z0C9z1S+Rn
SOFfymUAdqUCs1FigWwSPnFFdiun20i1//HAHzRzSMPP+lR3EnJc7+v9K8RrgWZHWBDgPE5TpFpg
IEKnkGFgyrfHEw0fGX0oVt1C59MYUVUo6c1oPTLA56/7XLk+HcZr0Uax8eUKRFlKRsO5eX6WpbRW
EmeA89NSf2aHtSxsxvsG1Moe/BPmQBRMUCPX5rr3YqWJnX2lau2sxEzAT9Fm/e0++ZDJ/RSRx475
ee9Bop5Zd+/jn7r/LcirwCnuVXOaUQdq1a8GjVtTeySpUN5ptESmNwjOox/j3sbOymwKIyCmtOPZ
Z+L+X/EyXVNQVk8y8Ax5psC7XdSRCh64kqiJGdLre72ekvX6lVOFFLp7J7uXrpBmaClC1nzcCrKW
b3blYOR0nYSBWdz3FD4QtE8CrpiG5IV8r2nMfTCF5QAQkrdI6qa4pmChuaWy7xEDdfZ7l6XUUkBD
e1IBPQRS92nZlK3u5HH5UIXHa1KMB2wf92bPWK15xAVGWhL3edqp2H9hb1gS0QN0Aq+j4QgLg2ZF
LqfjRRB/G39iLhFxGf/h4SDyYFIUsdQ4RRE5Dw8PY/+YCpxdFoDTAQe1y5GAPZXga05FTqN6BjHz
k3tAuYKC774i8MD/TYCdO5OtGyk12S5T96odMGDBKtWq4a1LCrJTcck1vYnnl8a1UQMm9F2x6UQ6
5MQ4TFUANWGvxEg1j/zKT7KaCjiojhgx7dPmd3cjKFsV3AzzzSdEhyd2RwGA40yHjZgeRLsh+xF7
yjqfKNoJuxnmj2N+JPd3bTIvnpaeJUpph+BYD9keUx3pXC+s1EOJXam/ZtkOujUEJD5uKgNSCWFk
RQp5QVboFyez4Kq5hZjkWERV5/xyKBP2qv2JEdKhjpu46wjaDV4yp9xUOb+XqicWqZ6L3ELUcuJa
0+MSYaYID6XrILVvtgsloqb2ue1vNyM4qbRaO/n1ZALEy1NxkBgsMsM86RpS6PXVlbKH3dMovR7N
VtB27jJZOvMPkJskhZ1HJ1XUOoFERXmOjHumZwlWzYSHhRpIQ5G5NrZKW4MQymMX/qTtQXIWRrCf
o1AcHVGXb3LrNq85fKWTZ7Bu4XpLhzckD/gQuUbikRQHAC7I2yjUp5ls6QvL6+nVk9+ydyAkOBYa
tBbcNSv1FYgo7FCr3LNri7YF7u3Y05MOX27CvlvchH54sISMSdj8hEjUbcfSeSYcGhgAw4WbESwF
WuqFwNQ6z+nRzicxIW0kPIeT9Iw5AFyecoliN1FdnBnI7anjSf23Ku5Vuxzcno/vcoJMxP8TQ9au
oIL2aPZypKStdMxfcfPw1cMzBj3MTgrCbkkmmrJTD9M3mSr+tjcARbpU5TeT2u7iZs8y7F2PMNWb
sZOe805AW5cPK89KL5jzPJ83wCPTZ3qXC/n2ILA+PP6Hj1XPEBPa6Zi7aW6cIK6b9RnCMW5X/vXI
V3GZXMv5oEDebrX33Jl2gSgxRWHlGt0o9SmyGuJAkLlIhomqhTePBP5m105j8vwad0naqoPFu3y9
UCPY8eTvjMqeCE3BNtn703Czh/9IIdaYu/tIAcyRH8acT7bGrjgIKnfO62rsfTLEcqwcIyjDnNCt
D1iaqYy4ylV37kwYCXgZ8aV28cYLxlhb7rAgwVzdDx1sf7nzpoYBQ0F0troOn32XGGieeAR3trOV
o6hjfwqPAQJY3UX5Ivnd7rdgmgU1J5hy2wRS/0Q9ZCY166kQBLf4c+OalvoHTuVHvrasjtr6nXnT
O6p1OQmOOBuXsv2mEifqBLSbZcZehy37ug/3ejbGO9tSplgnG90NlkcKLCbluAvOIQCYKsEOcgnW
+apDZ3OrR/cmaKhL/g2p0JDALssDovJw5Q7Q9wDNN1zXVNPGwbZwuFy3yp67pcmXA65ap7RkXy1l
iHRJu/u8qCA0MxQvxfentEb9cO58bhovMnu0J5yAwqWGJFu82/EQJTyx25ieRAzZ43V/7DjO0xt5
U6PF+OByVv2FZf+0za7wBojaQEL6mbWLTUBAIGxGuxzNCs6uWb5j1TDGJ6peocgaG6fPIhZhjrz+
XJOuN7QxR+8pEAyQ8+/Sd6F9XziQUozqIXCBp5paEBffpnvn/K9agquF0Sd1lPppRByHR3bvav9O
fE0JDOgZEG6m69S0tGza2hasGZcza4Wasg5TW031rLdyF6+unwEhc6wS6t+Add8qPOP9To1j6+LM
OBQ/uUDOXbpxez7uH9rg3J+BqHw5Kki4i9CtdKZY6LJROu2AewHrwzlTEfL8gujcNr4btv1ErR4R
0idQTwgJ/G9Er/x5ARm62SZXvB1KZ/wNYEWVuTja51jTOw1sA4EoJ7Zpw+mhcBWFHREgbcKC/qdQ
RSMWSCtwFV9Nm4Lp8Dku307qvBJZMBGy1l6J1WuSNnG/2oeEehrlTcyVYdV9YtkJYZtd9HXxxgUZ
it40DaFWdwzf63AumImLDc+EtQ7QZuPntoN25fFuxT5epS5y2rpazy4JL04ikZgC87+XbWAEc4a+
Gdne0M3PxQ7VRgLKHR+ebBLIC1iNInSVtle906T11J440dLphqXTAAAvuF/G6D2db3Kg+VSUav2e
ni/HmeMMvLhqEI6TZRLIPDbm/u+7gbZy77vp6P97rZx708K3lfK2Qil+QUPIYQJO2ix28nArY7gn
K5n28XjgHyszleHe5NMri1VnjGfhj373nV4SQkQfhOaRVzsw636M5prAbWeKciyAkv40v+mAX2IU
9rdZlYJLR86sfd5kCvhxTHxVAG/s4/P5JLwj5jZjux5OFt/kIRhW9Y7ycsPrsYXkA54z1KTnXCJ7
Yq74B2vV7EtCfqauX7RPPVr/AO8p2acd3G9aORHqI0cIRbFggCc8Gd5E0tiL8ngcFdr5AIfNNsZ1
9B4gIt8O/gQaw+gs05q/ycm3sPQBEvfHDJn2vw6Kk0oMJ/LQbiH39eLXqCc4BOX6s9eiTfkJ1dk4
tXi5fCvD6K27jZ8SBZRZp8GqxuQrme+xrsZoxNZirE4e4jj2YBvB5RtvERAP/CkT7Rbdk8Np3+YZ
W7Td+HSNHsTNcG9SnQ0pJO40zrTXTOU06iFmyorjBfNgcJtPCtrIQh40Kcc4M+C4Wwoq1s4LRddx
JUrbO9d2FVm8SiQMhtd86rTKEmUX6OM83NdVypwc+eefijSCQNJgtDyVQP8OQoT7RZGi0SX5dMwk
QJSLv1sxQw5+/GJadb23HmGv5+KCOemD2I/9J6hMAit5yTs4xUKantkq0iI8SrM+xHWvCIduJs5U
QliTA8Uw/CcN9daaRhiqOQ8C/OUg2Jn3/g96Qkt9+UL+s0wLz3/DIF7ezUujXyvpSjFXRU2sZqJI
HnXnsd7YichY/Mt7rto1F0gXNh163jE4VcnHJMPV7uUrYAOQqFA7jIaXoYe3f8CbBBkeXVou0Dt1
NJnN+IpP3Q9HOiOIhj1mEi06GaWIHLZZKTsNghIFE4nUxoaowLxH1VcYo5XSRTTFvKXAjGU2Ed2M
TS0xisyRdxVxVh2Ogiaxy+gr9yQnA83r3ZhtuqOaicCW9oqiQYgx8xvHDLbPdKZp4o1sv404R9Tq
v7MMcoLw0ixXw5amE4EnYU1r0n79lpgsrkJRsppqJDjepeCANVRIZA7g3Nzk+EQaMVhDNtJN12r5
mVmOXYhEgpBQWbFCZapPZi5TEoarhlZiEhoolmRCmo8Fwk9+NjuPRVMCvfmd0fX0AhAsBBBKWhCq
24GYGIhm3WDuTJ0kTXgPIHvMNZt/90Q8at/2JOE+4fgOH25zLgpFamUx4n59ANXWui2UZJNAc8BR
0S1o0EHk9NEMxN0fBV4glz+YXKGyKa9mlQrPtTuHOGCl/0esLoUZq5ti1pwjjdiEHX1hbiEOl7il
Ei19TY43DrI28Kbeu2NqrSChXna5IOKzy3vWHv/YpOjRFdbWvlhyTOqT6t6TUcg9BTT0x6OYx6ku
Ui40BCebut5XFUNkQOimEAZLwAxurx2OyzCvtmYaP1Sdv/QuVuu7wd7B77JrDls5644lF77Lgm12
su9xwLdt5yZeL/CRyAEhGtvQYbeYvMZyyZw6rvRjrMFUDxI7j++laytF1lPMl/0e5FUkc8Ur1pY8
YGdVg5q/XcUjKivSTomXGhha0Qr7whXBa37Z7RLOmXspjI9/2YVeO3+88JbxnNqHJegRtwlu7Gzf
qxfNi4p2bzykUmToAFqsXHUxPNxdKb5h8JEBVhMqz0MGM1FcZ/5YwcSac0P3c0BeYvKe0fM0hq6B
iX2jFj/JsXra4RYvVs5hB7Vp2acrdT0iELl5Px83V12QK9CawjqI6qvXhKTVt8R3Ybb/aOeZ8Oji
7ThOIRGj93pnlXUSxbrw/Jfk2SX+UkqzwGi3RwiWNsL5djuvuSO8JW5EvjXmOW2emqb9TVG3fGL2
F+qWkdmsYiVknwMradwn0JVc/cYVcOIIXDWcRtXeyqIxIozD3sbvAUn7VGhIwdLF6y4CTY77OHpd
isqf9nW+WBEFyvc/FzBrthcrxc/eUgu1n87YT/IoSekf8vnBT5w6qEYChtqiVx0gOz0fTySKWC4U
PhbUdvfBKi0MIfbHL7iNM8no0B07NSPQKPTe3zcvj5D3xq8mNhxPUf0k/npqHHVezsEl9nzyzMy6
ATbKdWGDVu1+t/3c028DrwAnnecS7B9ih4ihOTujmLi8iZvXb61K+o1KQ4dxNESe1Vjyp2VDUUIM
1s8ITbuKTArtdD80wEyLjS82ynW5J0FARQmXXdCoAW18m8hnJVbz+ptSreBREOvWasfJRlkhBHHJ
8UG0ZkHYwxYIxYB/meMSb9qgtfyit/SAZarG0VFHPKKuiU1lSkkJzJvJXn1cULaxrV87vg6G3OaO
0EvgCKccDWFqjMXAg4MJHsM0uzTuylfy1wxjQayRdbCwj8TVz62iCAXNd5152dFrhZPWc47R/hQs
4x67MaO8QxvgBzL+PeP0s7JyKv2cMmtYFZmYOIn5xQgqU8xq5FasTVUm0v51RLk1V1WSEYpmQukt
KGSUx9sCVcmoXBm6Buz4d+MNBOKsnzVnmpiTOIm2+c39Qg5RltdyfTvVrxt3kXcUnr+PKajt5z8J
XSWh4wxl4oehsmED08ZQ9I95S+d3ITQD5B8cRLg87wEdcl6pm4Xm8Sz+/y73o6s2GHYhCK46SxrO
FiqvmckALc1cplsAYmSPBbETD7KcwZ4VbBFQx6M6JcpsJimX10ejlHIGOLbt21B9fEwBzI7I3oEP
AqlEm1mUBCM55HiACPN5g4RJAXhDIu99kg/9VKIXEuDEIDonuisgH4XtHt+WIpb3fHD1cyzyMtlV
ZLYse2m8awWSjRetI/3mwPppo8v7va2nRjSbw7EPkRclINfIiIo5zvLPTy/3xOq7eKQa25BxIUyr
36kpRB7DLuS1fdyaqzgDk2sJkZV+QrGmQN58UYTJM8Z2BVsSKK/GAstYmv0nKpm2b5Fl8Xnr+3fo
3A51ztomYLEFntOrqe28VIc85Pjik0OUZQO5p1Dqq/dq+xdGKBvTp+wSsXCcpZ9OSKBdFSqY4Eke
YXbkufZBGBh+831SjfMXYKYoPo4KMckl8QbHEd1pAPzmWobkrY/jzr98qgI9AAR+XidCMv7VOJ10
9+u/OVteHCY9xZGS4p/EJAZdCyO6Zr2lGDvOU2wHyCmCm5asNley1GD52Q71gauInDJf2s4+lu6M
3tg3IARdakbESqDbYDpxb9pZaO0oShlAQQtb9vDc9BcLgl+FXobh79msIT5I3BBMpsXx0aqqo489
9i6+kq2HDVLPLBRKc7dmfpRNIOd8EyD5f66n11kShLvZ759BP/bjzKf0cUzRCx5M9v+o5wAofR7C
Gq6zesE+iB+e9Bm3QfTBCmZtHQvgpygJiPyif0HYqFPJrcl2fzOHkS5rPe6T2fQsiTwfsWuedQmX
wE3OpMuipScsj5WPjUptac85AsFZU/RxGhzYuz67yVxrsIRwzq2dycSBD9v+afQAcKLesj6Pf9U9
UZ8nPjlWM3XkO/4XLKHhT9D7fT8bPO/4a4YbQzpZlGM0q/cGczibXsoF2tx4efzSOrrw04Hv5f/p
COCrvjBmC31gPQoPS8KACwkNTFTw8HKCO+Du2hOzPEwzVFL74rPu0mpLnTwC7cQxH8kEYwAsF57V
VhvtwHm8xxi2xhGRKIJBhJ/gPefTycnI5nMDXSeHoB298SXgf87ZwUYRSIux2iB9GNyzUIMs4GMh
+epFbhaCsm0lIBE/OlhcUTh4a9jlfH37GZHOMKiGPV2MJ2Z+hsgzzHXct1QrUOmlxM57i/NgPxgy
q+1U4Vc2VFbphKsFKMaEe1Js294lFINKGWJLt3Cy2Eg6CfFK9Q1AVzTZj2/jk92QnmRhHgCAKNpj
Ir3Y2+MtzwQO8wq6TJGEtpY8GV4++KPLKCscO/PjHQ+FwH7WNdlkeqcB7jm1bC57ju3XZ1WP+YsQ
G2t6PwHN6fNd2TJPUvv0PiqENq2NnaGTb4SOrxwRtKLnpvh5fMzL7lzP+XvDcEiwznkSLOx/FQPb
Db1BU5i1dzhJWZnn311jr4LFHqTXazSlICufPpSQqCUidxLUyQXuETFXvBqc1iuEsvZCCOOU5LN5
Pk3l+jY+xTDe5jaKxWyEMbLkEVvTFuBCzo8G+vGIRAS2eToE4xVMnIvvrTw2C6FnVwmncgX/GBvX
Z2cnvsSj+KZjX1eT6lnoziomvT/qgdQoM6cH9z6ltCqkDR09iXqQloEplv3zmtiXK/fFsWgqdyiO
GyAiyhDumXCcIjsYhkOEhZR/wckQTE51c6x0LzqNemxQU9wYKDeNUie3SApV9+cBPXAaFETZS5Aq
REqoS9BLSgzrwJ/sSy7UXWpBoFG1K6Um4T3Y3qCjC83XENx3HWhmwbs/sIVQgy6yfvMhANU2o6Kl
Q4q+az+0FI7ZYgLy8SiNIZqHZZaf8XHvYq7gDsiz4ZSZ8UwB8byU9fmbbxy8X1mjOzRxTYNWQQPn
9tauN+ECm0dR2zd4D75RLNiOwlhDsX1wo6Cw1AKk9jMz04rJeo8ZBLZ7WZ3qzRapFzOYaUzq4B1x
ZScBz0eqQLJQTx7D9U/1ZFOgZdak302U9M8MuXY9vS2mDfo5Dfr/WNrjjl9IlB39xH3OoHKr2Yj2
Q7lQp20wPGihwilmn6ocZtJd9DMqUTjiI1a6swr7256OvkzyOPEpSe3/9nb8gYxxywcj96I1wUSt
kCP/cbjDPHxakkDjsLInX1VOhc6LyxbY2kQUQeqevpAASIC2PnElQ83drjSxxA9U7NdB+UxglYc3
zz3nfXKsV5g171FlIJMLz6o7djW7TUSJMautIXaVZKCNp+FPrIzd9lZ293Cdtlp+UQD5jOo+1F+z
s4DhK05Og+NTkm2Lx0+8u76Mfjy18y3cTVNehbiqg94YsDNXk5+NQKNSuGebvylIRFFU7nZuBOX1
kZshqxIBFQIC+qK4IYqRZk9+gTQ+4bHBzSso5a1wZOSoMDwjaUBQsod5wYnfq6v729EBSdm6qK76
7k49qGhQf2H0r2g5dTXxOUpyw76pI5aQFa3TNHFMH4MjCGL22lA0pJNfv+l+h6pGUP3/tAMCjHvK
b5A7GeBFBaLqX+IyzMt7FXsh2xh8iMbiBirAnmSbd/4ojExIW2iFxQAPjpgP2ybkPzArRx6XLD+w
XhcPbnD2sVKGHEw+v7rD79leWx1ypRQ0rR9nAzpiGe532ZlwkaLNPLfWQ1BKq+bQg0HjfEofIbo3
goxqAK1Bnq/pvb5mw/cqANzmk9STUBY+LkTRtOCDrPiSALik+4Kq8K1jKA+kyXMxf5giZXfAKDLv
DPwh2FllU4IsYQ7iM/L2GaZyZPNx06FOsFr1kbqIkX/BTSVKRIyvXoi28siicn/QmI+Jlmjyfl8h
4c70fBNN++kv+PWy0dciCIvtr0mqa7S2E9TYSbCOG8VPfA5f9j+t5wmU7ZS40Vhta5vdCTXHj3BB
nIEcTVUAkglnGB1MzmIMLEtpLN4uKM+82fjXChHPDP2B0grWZ/c/HTo71ggJyRvrmNXOkMPigWYk
OAkFz+YsmubBu2fR4EWrwjMxf9czvTruxUZiVKVGsOwvFdV9+jKVSQNATZY49FlbSG4PbunvK/Ww
BSh3u1uBgfM8BNZiUGOz71WYjt8EDCBvwYpkVm9hEaz/Wsm7jrTaXlTuD818KBZiaN6LODLnIMb6
1d6Uxayl8QHFHAGrz2ZTFKLGqT0ZJvb8lwtAOEArDRXb6QyNHwAi3Pap5HF0QftlHjeY1eBY/lNH
Vtmgpazo9O+ueQKvzEomuZTvpVTz41qWJrNCB+6Ds8Zg2jCsNv+QgYlJuZpSJ8ueObTzgNtDEd+U
JO9E8IN3XfAbd0WHIsAL4uu8gWuK6l2K2CpV+vjHEpkYBBGbX25FTteNea+WnuYODumAG66NyG9p
8dYGDy1aTT2hHnJUxCkyxj6ZINLlBu1UBEAtoM7xF6JQ3gdCTtuBIfAMrldPpunkLSARE7l10Tmn
Z6WrdI5kQMIuDqmqW9MGYXrLlsJO9mGPH0rwM6UILRIxeTtoh4lazWiICxd46El1TQ7n4RJ6LqmP
+AVpd3B+9u9wAYApzZ5WsHGpq5WC0CB0dBSpAP51U2AIKkhN3yk9127p6nspCJaHinkZzUqZOD+J
G7Q2DYPyE9HrSdYhA5MQl6dkhuwV1cjQu4DbGHmYySc2M68u+Ygw9O8LUv89IJwV4wSQYqgx9V5O
P3bO/N8FcUtvIMfkmNzzUSZ407KIfMGf475ZmOUy22sDdpMgh2de8hmQuOIKV6prW2l3GlEeIZvn
OSzG6reSzNJ3sv2X4mGj/vzT8PQrOGL6NKaprGpAMSGmLzXe+XPZtQAfjD7GY6+L0aSYR/FsRN1y
IdGgIwR1O7ipm5HP+xHr4Q1Op5dbeIQ1Ms21yBhBVRhys4by95nbzNY/UVIYuL8JKYr32VM5UMWH
3fUYOWfXgbEjNfme7vME4FpqhB4P58XCMNZ8QFxcd/yoA1fUBwD509HEU8CMFRzHRnke9K7MSNNP
O/pVns/KkwvOLQQSiFQ2XCrudpu+BtsSKO0UDUIP2a8zaieYj8LsnohuthFqq5E8xy8SXPF1Jp0B
+EkrHmAwu9K522mxdza8rqxsu+4C81oRPrnr7uDVHdnCf1ZiQa3hF8qFbNv6XC/8lLhVKo09VW+f
pdGwQXeUW+6ZYUWuG7P2V2HQsha3TxtXahWU6+HUjWXjaXcpZleE+cT9zj+j04OKTB1NhvqOuOVL
EB/pSdtFAH1VadM30r4+X8dUSocbf+7kA7jn655B+SMcnejn/dWE4W3JYqb3ei8dfvyf9jpBgdlP
+GUb3g7qFG+BpghmSBCmiykKjkeZmhWe0820JkAKlxxuXGydgenTOgD3r1VIYrqaWnnM3VWuOdPw
cT22Zn/q0Ldu20EJkMdVv9Q/bxJMrUTa8esM4B5O+U2wuBISVI40KPrnZ/Dk7ZAXreByFmgjWWoR
kGZt5G36QrJo2jnofMFDsfSk0PFJGWHD9z57k1zlwYWl5yWyQlTLmBDyjgd0TUfgDU3KGa0XoF1H
K5qrxAooRkc2EUC3YgcbeKUD9RXRUarJ7UBjtSvOuSd9lkVyIzCC99GKd1ZVh7s2xL12YA6kMM4O
HgWnTOD7Cpq4PSKGnoy2IHVNCrUg/0rB3kXBB/tSAr3nyOyrjntxIyfi9JhjF7JaNZ3I/MvDW3vu
3LqysFBT04D9ULRGH4kEqx6cyT3le2kXEaQtkiN1LgH3gJJG1NeIuHcX0ayorKH/7wPGxyL6Od1y
O8QsEMKmf/7KBVJMc61wV7LGOH5eJ7fp14TiRh/hw29Ui90CCwUXtDb0pGtTp3ZkeCHzVPNc/KT8
YVrZZqk1DvySJ3t6hadZCc1HJySTK47P9qLpTwGKxmzlecYzvva9yPI2wIGigbtIK6zdDBLuKjuW
PvAnULeaM55SfPWlCb7PE2KrMnaz69leN2TJLt5QEkzYzY/xdirDQ78AvunCVPd2pzEpaLXGdQWH
7UvZijbkI/dPxjELwJSVxuJcbIt+RL5ozeVyqBZzNTrdTHx+89EcQW3GwVE0a5tcEle3lW11zqw1
IkB7n5IyrtKkjBOD3B7QupxsvmSHZY5tTktafDVATYbBcw2XY0mGVXCL5h/h1Z8x03QAwsoRFASs
jiHbZ2KryNlMgv5Ws34aSvg5q9eC7UFwdf2dQ4/36xl+TLoE24w77emIsFE6Y8/I/GLsmNAZ+k4B
AtEawV9FH2CBqyR/vf9hk/C7xiLEurj2leFc8GZPldvZYK83nJw+nb8EkF+L1Fd7PE1UvYwW4v4T
KINd8kUp1nDk61m0NW4GGBItmFUvkqaHb4ZyzWIAF5nwUmGOoDiRN1fVuVE3BPyUkc19Fr0NvbqO
I9FSqfWi9UqzK6MIr2GjzrbMUC7cRSiKlpOvW8PzFHISiBhYEzngQXdVr3iT10rzKSBAsVxR/PRg
X2KOHFgSsD5gfrNksSmzKyZiZxRLryqfLnPOHWC8+JB0I1ZJvs/UQ4V+HAot9XPWxFsWUTNgYKgz
8UC1stNA0nmInfabzHq/fzb+7X2fYzHr9j00XCMHb0RcUOR5xP5q8CNyLcIS9xI4tUvkAMULi9NQ
FS+ESQ0R4NXj6fVQ72TP4xywg9OeocpyVPLzZ151AqlPEjIvn/hksw2eu70w0rxieJMK+soX20qH
qXNuMn6a4rRU1KH9hTHz0AtzS2WQXFvckoRaikDBKuMT0WIC+xDHu2UMPp5O1WkaqVKtFzTLEuu1
bX2nstn5biGEXX04IF+RZCf3MVuP+etHUbJtR7p6N//FaouU1NYRio8FHu/0oXHbM+hrQNroNtJl
6aAEZTcNvwBdEPBmFmDZnzG62I6gWdPF1pefhALirRMzhANcCFAz/H1MMe33BLSY1QzlL4gd60YL
oQyKwSnJO6AbLQBc9d/jmsoMaSIHSZVXukDrqwCN52Mt7yrm9oPgRs3MWl5xdW6jootLOaC0JQ+S
RayznrMpbXRyNFkAQR4ZVKQYZ4Y1/G34DdYek1EiZiiWYOVv8k9+KhjGU/pHPKO4ibQN6d8nTTnT
4LfJSQUu/V7hg21JE3d6UVwTikRJD+luV57sYge0pz7tMHse+sfWiNeHXZM7gBZxaWSpxpOkZNKI
+cUOmGElffsfn74ZhjbwrQaictuxuxLfIYwQLzIvTDFy2xDTlURX0s2cas2G/6XXVtSNK1gFAKoe
IUXsBG4p83IFL0Xn8UmYYcgvW3BUyy8I3FN5cJ+eP9SYqLZNrjcMCCoZ5MCQKPAsStHCAu6Ye/55
aqNjSVAvjgYVyjYuLTYyTNLKHXmVZZNbl2Fto3bURFO9YgrAP9BdPWgQaQVDz7PANVuKwUVmKH1b
lr4WZIaeyWmTbAkQN171O+yLBfmIm+7Ffuc1nleMiUs+VRzEzOVMl+nIdCuoJYJ5xD5lf8fRhMxa
ix4RS4U6qvQ1+pP/h8EduIT8WtlXiVY/tmcE99yGgagX1pHAuCQbeSSXZecqoof0f/K8nK3uBK9u
yBj95DOasTvudOH2YthD8uBN0xDZ7XTjFijMb1mZP96j+xuF9Ak7zzLKFmiwohlTbL54cwH9y8iC
MIfbChIPOpsQvCXHK3Xcx2F5k2/Xt8AsUiNKndUESURFxI4ssCjduvPCfmtJ8Adpsre0HY0S0N5H
5S8TrwTCw0Y82lWnBUNUCofbcTmiEkM+DnB2Z07BjUrLlIfLfbKTndhzKnMfTHGxGqoZr6Eht7rI
F8U6Bo7HPNIAE0dzRTWjV+caNbT+/+Z/FZ7Uhc9AQmek7qP8ytvrP/iBrT8buI8sQcpKCppOGPbF
EJsAyEzP64OvpArSddTAWjV76HrjBdj0bUwWcY+2hYcQIQVuaXegVCOGITlFRVhLzGxARFkiIii2
ppFEN/EJZxHEHo2Nhujp7MKZJs949jWnNwC+X410N8cj/98SQV8U5OW8WSHR02/Ld+dOts/J233m
9h+qdVdDfB+dqkuudrD+pxyVpa8zHajFHAS6CurQndXH4nmpOwW3wAFbinIERg3RFm0rTxmzMgpZ
NfH2GBzvB6bFFAvfOlhbw2mhzstmx1GZiPLiutV7/8C4DF4N2aa3cMKJImBTNoqRrqBxcom0WAGI
At6SK4DF7cFeN7s2ruyuwBGWl6BQtLLNSnQclUMRqou+SFXmpH2Gx/jiuC3fhGFlZYfUP610OAnS
mdzicX0gkGqlMNQy+AHxuZv27Bw2cB07ELodMuBVahZ8T9Jrl2WdyUqODT+1ZIvUD5dIxK0BjrVx
+Rw7T5T+xEUThhpjJAO91Buvbm5Oevtd+qMSe83bbaylPMyxXayZqaSnm3JOAOBblg9Bs9zxqnOU
3seNAoYRidqa7z/WyuF4JvXH4RZ/BDk6M6849wiqAN+QTVrXIm2Ql2xJSQgyGxqj1UY3ArlViHtR
vHze2tCJHMHpz0OfgWhkKMhZWf166AdX0CxCfOhizLHPLdLeg1wBgLo2tmqT8uzSFrSvGEyG0iuq
1KnnBHTCtPanP3o1ZwU1vzMHcQXBDyfPnw2FZf86N5NltkfvMgin9io7WWBbYLA4M41mCvtgBKmO
dsRIX4r5Cd7Qs44iCJSFFqsi4sgI6jGvWTjMzu5HQwu3D6d773dc1OwPblv5eSJwe2TcGO6caUAr
jzqVIZ+cWtyzeh4AmPoMMZpMUE/a/05xsnjmSgK8BVmIWJ3eDi+SntoC3Le6K5HTiNEMAcg8v6FA
GA3BzTAaUc8atoJ1hHBdKWYpo7ZEew90TkZwWJlAwqdBh4h3gxHQguTUcnDmVdMzW7JHYkJxyg8Z
+DNVwUwtbRy//XMICev4m7VX5xA54JTZMugqPVNMSFqwX5ODbjMfNKUMXx2c6oBQkuwKaHB1QHEo
eq2IQO4za2VN82rKab2H37WaL3RUG89lG1vP/A7mxX+UZYr7wUR+iM4WBi0PAdbqBezMfe915xIJ
UlJ7xq69lttCvpVeNW93h/BmN1HSM6+bHvz9zCZlVWo7zj26BOoNe47Frmjg74unaGZf393Gj7cA
JliqAKzWITAyyQ4w5vpZDtjru1+/leZuCeyVYEVW2w9HrMiMykflStsv+ISx+lsjSLPIvT5DPpLi
TMTPf2uPdCP0Lp127neQzA1ceOgDeo6JPpYbi1pWFSql5Y0hc4kROD1wFESsrtIlIY9PBd5KmJPc
R1BZimKMaAVe547n3jcTqS7600FkmENxaXNdxq0li6At3s3s2AY8xxigPBjPN2SCUTyzJDvYZqHH
X1ZSAyvowzRF+pKAKBkuKsXqxH823TlaS7dDcamG76CPsPlA2i4ckLjmUSbWfbKUHTrf9FoVC/m9
swlFeEnndGkcJoJfLSOb2LExk4S2pZ3TuA2FxD47Zuni0bJAjL8REm1j7KLTzyPU229Xz4Po4yvp
w4WbpdHxzuqJFUS7Q8D31hIWldTli4Fn/ce/hhzabV3NeD9TDSwa4LXHlA9/nQ/TjpSzPmDpak+F
acSuE6m1gmyzAIhikK0UBdY2erh53pbh0MPKYTy9eV6Z5Stqw7d31i0lNhJccNdCjPbsLYEVwWoz
hYxLhN9By/r2mG/RFsopGBQTYY3t/n4CVY7CCWvAeFWMn5yO60+EEgU9ymtj2+bTxm89VxV9Hkxm
iuS2B2KKfB8bDE7jma232QktlxwGMD739x4LNC7/4MCJmgpcWFtIEgnViIsw6QYmUp9wRydbRJB9
LPk5Ifjhou56rgUXOBkuEVGBo/Q7xHssdUbNn5z6eDE/ebW0koCZpJAihA+wYQNFBvXyNazCirzF
lWVDGFlC6G1mMqr7kMBOVyOaVrpfF/RUDy8sWlHYvLZ+6dT9JUtRN+FRqin9MmqLmRdSGTSdXkKe
eaF1yaUi2YHBt/j5UXMf1WUhjbdVJ44v3tOKAgRvQOvQposHpAX41yIAo5+2wN7kDJ7889Smr6T9
LuMhzHk2Gry43AdZeSdbjUmtqYMc351gmn/4r8IFuENk1+GzRbVAt7manrV/dgjYXgewwNguCal2
6qhxw3YlPCQ6/382e95hDnNpLlgT3KpgOujID0RDyyP1kZLJ7dloZ2LznCOfWDe+DcjNcJd3DFE2
NXs7CS6HwKfOBgIGykYETBdHy8uzG+dJILzv4QKRSzSxuXjccNFAbrix/sDoOYD2GsdnCo9uI1Nk
KHzjXq3lxKI+5rWNhPWoclEEL9fpNfce7C5iKgr5oL/OFsxuzeKlT/1zHG0JKAGqSFuutcIFq6kT
y9nCJLiG8+4dOlE4L7kd+qtzGyiIiAn93PVp0n5TzJrJTnl/p59vHv39jAQYqsH1OWWeAIBWrZ3a
7O0rEdI7rmCk/+MD1WxMgPx5n4d8bGNzwOgjEcL7XO6Xnj9ysrxeAlQd+qwggxla+wC3Xx8XrEi3
KODM0gl5G0x+wfEE5RyxerE3gc5IJvGgSTljVWA7dqoODufgIYsJdEhWeBILxhtxnUW6/Z/t8q0P
Yk/9oaSOtOwYJOSSl071gaYYJ5iAjQqN7vfzxLj+C5SbX9K6amXmm+m+7VGGs1LSo3JQCSn4ni44
3x+JTvx7StxIBt737QHsCopT4WG8OB4UFakvWSH60p+UVoo5d1P1BaHJ0OMdpXS8NLpN90FrYbEh
AD0eEx3J+PF0Xug5O/0giOsR1NcLRtC009ssfn1dThCqZcDtwBaN5mAxVzL8ckY/0Bfb/QQ2Ad34
89ra9Sy3qpKh3LB23EudzG0ZHfILhkaNKGEuuhxpsDKDNiPrB4uaRt9gGPPJakd9HZA6Ou3KvuML
Gsz5CVE0GSbmbdbD+Yx8WwuijK+3qK66WjE1/msDQPnRcCM5lgUS1Q3C/gBKfIZ/MRD3faouxQsy
ebyzmakmXovzTnPwAw47LIqmUMaegkOb/BbGSDKoh039oH89i1VdMp6yckk91swvTpHGofsLsf3j
/sZTAKzjSFySBXCod8Uie8qtB/zlXcVXzKRz+xSxpULTIOu+9tI+NTa+8tAmeyYCNEiYbIccIzaz
hBLn+h1RwTgr5iOjVBuz8Dws9XeWVaqhcdiylDlFeUEQGhE/sJo0DMifhVFJwZuKcobq3OprLng1
CogrmkKZJgit0dPYqiZlWirwTsFEUb+oGrVi5bMTUL/oiIq2itl6OBR3gPibsbgfRKrzg+utxoZP
P20sn9tLYJfsKxFdgkxKbJc3HCytl7iQWaVXKqhkaQkJyLixnRyIOr3CMOZ65OzVMKq1Vt89aubI
GTOV3FgteweeIHQkpZY/jYXXbi2WfiHBg5Ppc0XrtcslmLAyKc9lbIHfMDxhs8X+G8Lvj13j9CNE
8Z/OsxUrGqU4Bf65UVYrknQ0fbFkOCmBCdsbmVP34Z9/GdpVkdq35JjJ9eZ1uW21v0RHk2ilFvtq
W9/FAImkuCajF+KS2EW+tSEb/SyVuyD1jvyBcRrF8NoSROkD2FpNWVSy3sxB65e/K1HiCyD5I9Fn
vji2vTnDtGkFrFJ6+XOKW14m/n4rt+wk4GYdlc7/RXty7yYvHB54Vj1gC/vjByrk5yJLXlE66jFc
CgXi5qlF06wmKQ0uXB+x1hz9snyXsPx2jNbex1PXjPB5GNocIM+L5wHVa4Vt2Ypzew2gUtAfWU5n
ETkwi9bUCFwcXrJGXg2/0r/GBy5C3ZbzvFO9MH1Xg15Ql5jvRbmUM3qlYoNa+QZEQ7QuZluFZgoD
0Zbca6LuPP92iXDlLgz7C/EaUrlqMtiJmDsR+dEcQkDNj7pq3Nzeaut7z9yxoLzvbsfWQlvsqmfD
5Ahg3+Rn2lwqm42Pijn0CNSnTypKPFLhaWOx36PyTSbunCtPLQ84fDADRYDTP30FE9asKfRtfCEf
JNWaUsD9S2bILAb6IMiG1T2bNQ/h6pJ5JK/492Nc2FOLIhZzM8hXP40FtWI+gU9qUgoO3NPKcNnK
tWmiCpFk2xbWKdGCJPH3SU3Fp4vxPh8WSGOK2PmawY3YI7kVnaf28C9s8CFYgR4fu7S7MejFDJwX
CW4p97HI0eVKzOk6mzScA11SwtMSdA9JoHdTGlIj4TkD7JIU2Y/oBtomoy9rNcrkiem2vzNnL1rN
f2EoF4x7EKBKVmpDeSFHneHx8HcTNHAc1wAe7rzcnDVZfYItzj9IIomM5Ab92bDO0EEab2JaENlc
d+XSUu97MCO3//GHWBnkEeWnZ29L1+J29n3L+ctNPbB81Fu47K/RxLW+J+xU9wTrOejRVtxpDM5H
NW4fzpN0mvZxWlTMaXlpQYf7FJr1HKJy+MdqjNRK8x2eVN7NClTiSRVH8stR3Ll92ntDMlDsBJbw
WwCKQ9fhE8CSe3yEnkg0WzwXZz5ZsKtEudwRN0kiSMF8yqiiL9xUJx2s79lZZEI97ePIVV6Vjiid
c9l8Ohi0fFPtWh9z9rlvDy2IJXlS4shUS8C3z/5YswQKRlNhV3oPINqGIfQPjAcswKvlClsxqq3k
kEWjkLuctfyJSOiD24+nGqKFqRSTpQ68ehrso2kBaTnbwcp4XbNz89mYKQ07Z4MA3ejF55upSQx0
GgvjuOljrLhOh5cGX5vGaPWpisE9Oj6jHiXSXkdRqHdRVQRdfXKR
`protect end_protected
