`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
aFcVoBJ5XQoYi/2dOzRV54UnL4j4QoxER973fHjTgAIHbAOimdGs0qQVbqlc7E9PU8yhxRU86iv0
Pt0dMGpKE8EB9gytsT1rlqp6bchfs9P8b1KGxFRe9EO5bm9RCTvvTYawFZrxqH5XyP1MxG0e0pZr
MswX1lqPdh6676ntictTFQe/PnmNtvb13ZHgP6h7EtH6l2EkJ3KMdlykZQ3NC5UD/+UREa/Lr/MG
a/Md4uQNSi7NQigbcs9fQ/de/34xFw6b0shICc1s6PF1DFlUGhKguXDFxB8G8i7SyXt8woux6vdA
l6M+kTk7UXm8tk94L8z1/s268rAjtWCwzCHOfA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="uGfFcx/SXHgvLX7HZpmySpXFo5MReYkmn0KfJucbPFc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37552)
`protect data_block
zKFBo3C5QUZ3j680ZOvG6TGBeK4QsIKZW8o2U9jKRP8LI3kfScw4RzrZC90afCELmq4JvzNyTW9l
MMgWei7+RMPhIhYOAgtPq/SKc8ETlb7O3NcSFuWLrywfOyEV2BvTwS6WPMGtA3chXoR/OJZ5vI5b
vECWScSVOUj9kHfYHKLnRjcbV7ZhAMIMlA45tQ2fIPFSwu/LnxxA3c04zzjKM65O4RFvkAUFue+z
fIQOtzjM1E9vjm6qR1T+5MJmPHCzyeL5McLQbXmEj3Oq0TCM8jJUhjePHx8bI0NwUyP6ipilEVWt
j8i5tHfkgSF7O7JKbdgg4RuKMLaf0DrZMLQMYGWFAb1tCQaKoRGJ6S42JEko98cpodx2LwxOvSW/
8rpJgEudz9wPNKdR0HbXu9withNh7dMGQDU20Kwr+Y78eIKHgAN/pTMPEaWqxeUkX8yrhM17vLQ8
Y617zduOoCKRNEMo3S2rUN2W+HxpyAAN8cn5Vee8tgf3LM9M0w2LPsLr1gE41ELY5doRWGxINHBt
gemYl+4WSYLGSAI3z2hHeHDRr6HuEax/sSLZSspLDstMPpyXQTB9OKBAJ1WHO4+LS8O9INDTdAtY
eol/BFtCDOJ4uwQsb+x6GWDx5CGkkuLTxAHK9rPAWhtJ5D+URReAhEOcOZsRvJzF1JQnVVjla2Nq
d9mAHnd7lojbzgW5cUHtp0em6SeaqPIik9+NXDNZxmcQhTw+6kMF9GOzezaW7dSK7WL7/OYoq/iW
YO6W5Ergmfmg7oO5bB1gSPcME2DLHpaS7XK9BJCUt7U+bdT2mTe3VgkVRjG46OQzu6bAhFAEIQYv
wrHOWJIrD0shB2iCq9Xy+rL/BVcrmh5XwPNqQy49/8dcwzi1pl3IHTuBmFze6Lgq3PHhVzj4cZ3W
j5uu5DSg/YOHzv/CV18oGbXsG83txLC8DMeVf1+40elvxyPe4Uxm1/+X1mBk4EmrTsrF8z5HS+/F
mMPzPTLceAfhrnHgnGXECbyeZ6XdYAEDhs7zTRC0/FMi0a/FJ40EaUJ2YhHKbsL7jy515AZD5N6a
k0FdcMPz++8pw60kgRob6sBd4frttiDobIa9je5HU4C9CoCzHgpVPM5dZU2DsxnwWl0XxEvemh3+
EaaaBjaqRSqt1MAx35Nk8B/PdEuh2KDeD7EAvP9v9QFP3giml54sm7gPdXkdks3tJV3F6Ne8kd7b
l15B+3SRT1UQ6RmSTthPlpBFUnIjARcnIaRu4UwK89m0B8UEwYOddhnboZdIcV2GLXfQB1bsujzw
j2hv4IuyFoyvZHGAzB0fsRSXszqFirKsVCh7Rj2QKpFQCvsXsV2r2Ro/IIS3di7c7Pyl8AdyciOs
62kQfV5kgA6Lu+e/OepPdgbpSZMHCsCei3xVq/uH9Ahf4FcfZ4znhQ2UqZFC8+UI4GM0KDJS8JQb
I8s9Krd+qr+l/bUOSamx9MDYrAQkIFXwW5vnp/Jci5shVxvBqXEz13/ffj7bbSr5rTn8MgcPmjIo
jYnJqhobxTjR8WFLbQNgWSpfJAwMy/Aupaka5B6BIuKxBF0XIDAyzUmu6dumVtB7vqqlqrVQARrt
up7MnbkgavqcuvSziCM0DVgmu70T+cA7TlVp3KYh5MbFPugBmDdIZQ82OY/K/UEs51r+ZrGZh+8c
MrYOhJB6mzsBEf55tOUAritIVgzat48IvXU8KK0Ese57vyNqC0azk2lNLkDnhivQDQEmRGA9WeWR
fzZQdMrhxavoHdoxRNTVs8u/r3eQMztGdyD7izOVB1gsqJ5J/10k4kypBVog0q8VkV4rf6IL9Rmv
y3UwI57TTIj6jfp4uGVQF+XXWFsx/987likO1Z5llWuOdJhPXmMWHHBj+IQW5KFRBHRQibCzCczn
vmTiRGzNz31YFHZoEmzU3UU1GLbW1TAE8yHzG+WxpIuYFy7eC0WGJgVAnXB870tFHpEgTG0ooP2Q
c42UGBoDJrzoGqOLn33sSgOPqfgSeOGTKs+cZJnm9g4xTLqzt3ptCiDyfPzbs465J5gw6qFOgGXM
CmGRSSgFckvhx0Gu3PFaomAx8WUPSa4GpCdanIuh0YxE7r82IBafKXAHuGDjDZQes3ULov8Nk6XW
RMdaa0v3mT8GZklHeYXAqZo5j9PUP3vESAKTilzEzWhLghr/5BNnWNzKEP2l3JFrZ3zfeoCLRevm
Se0s/EDGdhp7zVluv2Eb0z7YoM8fBq6AnuHtLY8R/jDOa4wJleGsjMy5ISDSvYeX4b7NrZpsVP08
A8XDLdSwosbFd/fM3qu+vCjaNnwvxhlZ04CvBTS9Xp3JBTpdssVi/PHV8sFCuVolkaYsqSYT7cuB
3s8/aZ2iq4uwIZrv+aJKOFqhvvEQPTA/iN54y5pEJOK5NsSqVlkPYC98w9YE7K6hOC/J0xYPJiNi
ZPHmeNWeDeJfBBbq6LdZ+sCdEwsG3rurAA2Inwyvbux8y4mK2axqiz2bxgJlBllcpXQ481opPU/2
/HPoFeincxoiGHVmmSFMa6Cc4ybsnQyRtpcXSQECp6QtCqtdgaj19GUIO2wDBsKWFrxDRya9I1lh
IFQhEHFrypAS+hUaq+/sVOkSA/m4VFYK9ecaZcLqc7bnN/5WsFW7wEFxiqsD09kaMHdkPteY399g
o0CQkCcFgf1hB37bdHP8NSH2k/eh7GsuMBXnsRjH5iF1QbbvYWL4wZ5Ym8o4cCd3le3iW3mD93Ay
OjUbT0x/oBRq/7lDA1awicaIu3tk8Jxpqpzjn1j3iSwTpdXPlE9azhDCxQ7TkqN7vNODAR4zyCp0
H9ruHGrDugCy5HCaSLcRxfFlyl7XaU6R0E0mvVMlWJryKP+aDaDJLymADXqp5u/+pX6X81aaM+57
igLJm00dQ1XMfekL3wiwVTBe+PL/pI1yHcvQ2EcdknfRr/0ONSLKVE3VYnBU/ZcjfUfY26siHNga
8VXLnCTXHIG3x09Tr/RXWrm7yM1PxyVhvlz4TgZMQKteBQPFn4h6xLyMJ2t4ug3WZggY/gOlUdNn
XHyI/ZYr8PYrdFoOkCt90pBgk/Nx66DoJIyLDuCNRUOEmkU8kpXH2aPH8/ssMgukY3wK6RGNYN2s
ZEF93Evaaic9xWqOPYC+YOolK3AyH4ly+g39sHlIaPTiB6HSA2ttzkUzK4ZKNJ8n20GpdtAIt/iA
C7lPz541ZhV83GotvhwOMiAsLw53nAh2SyD2LbhmFD5yvuC7IChyzn9QDxbEnzwmz3GAJzWHXsVM
qRoiAkYzY1qp1dDYrPnRzFiTrNiNEYqRsmh3TnkwhRhjbA3DTAFtBDTQWEP1AljBaWS1uCfoUmmW
UuDdzbIYvJ1LAr27hVtubsH5QdNWQFGGFZea2OZ49zw1sPv+1ndiw8qPB3fHtHberq1RsOZwGwkE
hs4/P5tGa+3GmFHBpb1O68Z5l0Wa2w0zH0LaLlVzQMGxJruHcCbbbDurEpTolxp1PnHvo1XrioOE
e+lrPbEogkNJwoKsx3rWfEPYckqesu5DRMGoVFSmOJx6WHB8kDyu/CHO2mKDZCSEe8qsloIycdaN
XhSE7omdHR7HCt6sMarnKs5pxMipUXxKVEuhgIwkjUHyeZ1zwJh3ut8hjvfNgfVxAWVEoC3uIe9f
/5H6V6Nc3MIZ74HygB8Z6u/OJfML9Gaw9/kRTke3K8iusRMOVQ4rGyqZxheYs/KSXFAYh14rwRnB
cTddV4sn5K16x4r71lRhMr9VhEBamQML4QHqUzm+OfkgtnJ5KaWz8YCCc/k/xiETUnMUxeBEU92l
qPQQhuKo2YyXN79ugpWnuSi5azKQ23msQDJCcZEO7KnVk5FF9LmLIUFmYh/JxFWvgUcUvR0iQ/86
oYN9xbAUr617zdC1KAMILMHRWYxGF38XTZUZv3FM2SnvLRUtZsb/adiFRf/loo5WoyKlZiCVYC4U
gRtJOkRUbVFHHKO6I5np51rlFPDBPw72TcLoB3c3uEORgd8mI2fPq5q7bAIXxyxW/eAunUkKO3de
q81hRKSORhVuoZsW7ykid1o5FceMwykpIyMg+bZMLLhE3cUI+zXjGj0IdDpPsr5Rv3HsPDEceYqk
3gOZQCCtuz6DxysLuS7Jg4qCeWXW4X+o1Slca0qec41rIXRKCwd8Be1skD5tps0iWVYrJOWmXD5c
TK/kkgPHPbjU613zWXEkV6/hTF4j2IOCZYBLi3ESxMlQbDmIGrAc4p7R5dUdWE/jS8BcbvsuwRo/
NyPMvivDW/IFtYujJbyRlOx8VpMysfeO4xS+wPXiq0ywAQ+0kj3k4B0ucG5uJCTiiuYbSKaoKHh1
oyl3SGVTb04O/e/uRyEVTz7AbpFHhYSxOQWGaPlZCcleKdMAopmO85rWJ8Pgj6gknsul+YtkqD9B
ozkKzasoCiMEBeqw4R7I1kMEttVKSLesvlIdx9sLHQ/aIFYUU8cxwQLeaq9zv4wIdjenRz+vQ2Ym
YB6XwKehTke09tP3PIPUYGePH6XbqXuKWTk49nVX5dA5mSdPuUfpQ9vS7TK83R30szOWqTlIzco8
ariEUm+2JfmfPqp5nDe1lHXYMXzecXA/Q8QVSNwOY13aPP/gr9jlEKwDwqUu+ulAE9tX/x7eGA8Z
gxlPD5NhayvhoziJ+OI8u6EywTgJE/nv3dJcsrVcfMupy9N1Bzk7yVSmFbVd7lqR9pe+s1k7Fd0P
PZGNN73XI3LaAHnJzMDD/1NOBdMvHNKufvXT5EO6tIhShQc6dgOfSHyx6fBiXRJfXQwCVusixOhQ
zxi/aprGTQ7vm4r6akzCPerkd+xzPzRtQbp3I9dECHW8zXYm1eyfMXk2i/DxtdBnAtC29XZV4W+U
y+xmUOPMovIxT1pJxoNewF0nAcO/8g4k8HX74BYU7dClyAcQKz//e6jkCsmEU/4NehOKpXSpaAVg
1uzU63BDOl+SMeX4arra9CHbegI2BHyS8aoZ1rNAPzixiMmfYYMhbVpjbMP+fL/dwY8FNw85Sx+3
VlOemd37enCPZLGXuRrppJnaIxd5dfBGJ3mETd+MpXMNhxCPKuapahdhxSTAVHhnH4SpB70Vsu3W
zn5QGuDIkHwc/HQ+lou4t/V3vAGgQ6A4GmOuiHtSOh5tAm6K5DErOfY3Y2e+xvE3uD3WlkGGdOYM
prgme1Pio4ld2HbLUASU63Ku/bwNfaRYMIWuTrTmT5eRNqzfy+EFnoRaLbajA4JhStbRUE97zoB7
DvF3+O/m6L7gl4vs5PaVLWZ6vZf5q0sIYyK7fqo6e4+LcBfL7ktMP7APgdI9086TuILdDJaF7lHw
CbH5d4UjPQILmK6Oi2LbRjIcN8E2VH3MhIr3wjiKts5wCRzEcDvPdesROexiw5SmWEpOlVIP6qq7
Dwa9H3CIWuupYra6y75NBDy2/S8B9hL1i6P67SfW3LF2XtkLHMmaa0p9Wl3hk7PClQw5oum0Bs/n
uhSZAibebpdoFiZrvw2jkKUENiNV6rwo2VqKNuI1dzkfFhpPpumF9VGQFVTgfsPwtjkzripunGOf
0PJXSlzPjDrO3Q+GZR6rCGl2ymaSB9XGKNYPdDQ+Ev3Vt38DbyYT1DLZy8Nt241tvi3WDqPWSdgd
sfT5AXJfnBNuva9n3AweC7ts6rgJmjVU8PCDWd9jvcT4lwYFtwOycOkSGTD+LrRL/xyhBPyWXL2U
JFlEN9Yrw/runFqUoSXcUPFNwy4A4aDgE3NKlYu7YwjHvOG6oFzUMUqKefke4bHhwq8d4hco21eE
4xsjoFsNh9XzWCS38Wx88OFPhCaaY7THFWJHLv+2+t3vaZ4nQDSB4AA91tHtwioP/l/Mn3I1jNti
wIuJ+uhKA9zEmYsGVcSGgM2qTssGV/QRRLgDf9CLNfZAFZCMGz8JOmpNohPqQiTx4rGqfzLZQBKd
cKQ5UN+cgeNvTsPCGzt2WZGtf042y5GmepcPzCm8buAnPjUloHZMh5ue54+lzbEU5aNteWH4zXI3
UUvr+BjD8qm6VF6g3evwR+5dCT+A2aNGMYjK0nIYAYlK7SQv6R1LVr/oqYCe8CbxnddVV5rl1mnO
69VDHwgD1uINxtq4muC+FYIVLA28F+5ySrQofFlpU1XHWc8Z7uGAdvmfe2iCWJeoIDSq7Y3ubUG6
r7cWqXyOx3GCoLT4qSoSKgfdPPHNq6A/Mas73Edx3pu5DEccDT521ztlxmurVTW+zXgLFSQCCWAp
wv/ANO5v160Mg8sImoVVWsLr/Ent5AgwMqSH76C7YCX7RWIvATOd+jTckmFjvdmDOlAG2oXxqb9w
HG4KfTkY6BVY7VBruebk0qgStIXZyYaEFI6nPg7FXSa4xAMK3sNFlKm/L32NWBQN/vrKW3va2iT1
J3qmzZyNzWUdckrjbLz2reG5DPOle/ME6o7EZpZWKSVbi+RUrywa0gAbwX7JSPZDKqfk1k0CPZbn
rVpeokbbAS1aofjsqxCb9g9vQXP42rYjCGBbhJXNjoTcK1fP/0sG43DEGM7DI3LNP8af30u13f3O
AEs4EucIh9SWgnc1EPMN1FQLrgmS1O/yAbZdJxknGd8nhCpDmUxQ3d/y1n8VTSS+SnrTz1v56Wr1
eU23LmcWW0SuBQ1n7jmH+MeMHnd1Pu85PzOeSrLElI+ZRMe4RfPeEAPhgNer851vCdbYy3bVK/oD
qpWmvjyPnv8pEETV3Jf26IhWRHsMCpdnd+vBrurUu9Fv7zGlepv2xNRrtc/TuB9qYLyimIFN1Prz
y/o0Smd49MlhGVLGZYrd7jfz8vZuGYduB/IBTYWescNqqhwQVfekiX/mKmW5VKcogLhbdkswwcvt
wKs0iR2Gu5kNgOZ/vzFgJatTieM6rwh4oHBdrEVB8wg4Z8kgzJdrBki7tAPwXCFvqWgreaAfQ3Lh
hQfgS8IWrUQk455sSe4IpfpBZlidG9tvKi0yOdtbkTEipdMzdmhyIvr3d2Y7nisyzhr33uZd4vk8
3Nyj/pPbAvu4z4zD0d3k2xmHAmuDiXsOIzhi1v9K9YFqzDLb3rSndJGLTx/E8w5S4/t3gZaoh5dl
rxs7jIjv0964IE35Xpe+pV4XCjFEJntS9mezYYfQcYB9zXW3IYys1K51fyj1n4t2/WXjZMVtus2U
j0vORkrbOV+IlZA3DP0id18h4bYYYUJ92u169ZUbon82c6BMK5vfVT+fsaDJlgMaLUnjc/QD0OUk
cVPAl1BgtZw2WdjJkUrm4IGYf6SGrVkC++x3b8Iqi7xTvEUzPvo/bqPRptUKEQuXU2ffEN5IPlFg
3Jakca2k2JUMFO690pdPpGlPTg1+NcD6kRLGQIr7+FEVHcq+WgQxOeLFUitbFztHR0lzaG7YSxb/
ZnAenpQ6XS9iX/ZEowXsjgNre2Ja27JoZb8/qgKsehGUysUCIi5yIb0YEZ6WVNVfaM1Ng73BtJyu
88gYOvRmh5FxsYbFgLtuMu7JDOmmY4bXmv/PbtgwZl1CWf6k3hvaA7ZgGI9rpfAeLnDlR0nXHODK
92MO4BRb0QDesUzlbvvw76XTONHWcZ6iOfl5M6CsX36wvciKMn0/IU9m7JyqtdcV1G0M2038EguE
6h0q9uOShrpG1m65kAthAu6b4i93nny/WzK2tvecdaPWjtxXIFmb205xLQEgRLrDddUZ0dHapWEM
Y6D61LgaqlzStmdPe435+GoTh0N88bI8fJ+hZHo2humXWVAY6UW2MM0CZPZwKGuB4lke+0iLlCdG
kAIgjCB1InPqz/Rl1QZY+X2N7DB4TiVNouL6fQw9rg1Kysnd866p350rveoo511YnqCem2mg73Ex
QATlvMGohcBpyOxZ/IPELHQStdG0naChweVLS5TwqsAI6GPq1kIKQANL3rGqa1UleBKIUbfVSz1k
8oPg8I5rNCzPEawxcDbDQcrMeyjADYinEtuDFJQuKXylsgUXN93KZ/aaQyP3ZWAeOr0C5m3XLG4M
Z62/H8FaV+cRqErQTtP7GfcCwbAEOWn/8LQYCGmm8pAl13REWxFLmuJzUq+GQe6eJNX6yjanZgl8
ilCJTmHjEDs8f8rHxXAtlBfqeVue83wfMlmZZ7X/hKpKiVSrRXz55KwdPHRModS4S8gjTlMjCnrY
FXd66ijE7ApKkuRpLWUj8WDtXYJa0Ha0KslEi+q8xDo2mzWI6aWMDpGJY9C2LZpf7UhyGwO+qkZV
DckDmATQu1uEoSON9BYQMA1+PLYMDLD3ApMImdzeH0ob4lvpGHRqxauwjwZCyHZoKSb5SdZAVKkA
2wlctEYfd87X4sDEXpYrSoVOHgihsSnU68oLVKqjSz4T/LdWaj0bMXrcLYQ4jGA5+pG2qitmkb38
0Lm7bQAWLH7PeXg3EC2YjU5xwWkbdaxCrXEaqsaSqI98bsCBxmHTpL/s4MiSKQc1bXvKtP9R2cC1
WAXrGuKKFQvjE25QvVfy60WBuZMCmmnIzQdrz0pEYkg7oWb1ORjVlF1O99sRnoo2m/tHqovIqu+x
aGlHwmFV1tzHoztG0mtRtig60eeWxwiHSAjZJOUuzRlFTxllDPAVSZQQ7Wg22SzbVHYL4szuNg2T
x4vvXifDqsoXLwRbgo6AE94ubkzdWNQGJlfYZK9lS8NEwXHTdBV5IKVkAJU9VJycmPxy0Vj4y7CO
aFDuJv6CvOGyB5PmQnRzYfJoZS0BptK07it7g5mOag+lpAOd1sTdQuMpeRQbzw5QNN8PgT0GDtqn
uxh/m9mIOGWLOMYj6pVRcPRRDZmmubwbYeJ2GEjq54xPQ+VTkk3o65N+I13gUAcvjwVJngVwlIlu
cmYrtROeYETVAWRJt64Q2ltgjuZoY+eSSxkg+w2BzN0ViFb1sfPu3qoB+WRdiR78AJhJElKMbPmg
UbWHLmbm3Lwh7mYKXC7XwP8Q6pT8E+KG8DLe7e2XPz4Pzo0IvwvsuVYmxuphdgYDOYmqkPuaSnmi
Nq99oe40VG2I8sBqKdNaOe6/Fn3J4/Qib8pajOCWgvEtWLtrQjRokAPIh/HHQ/tyNEpiWbPea7qz
VZUf132q5qNzcmH3gkwlIMzbLGusrYHaWEvA9WhK4rbLJtnz1v9MoK0TCUrFzvO4RheZ4owiR9jd
HQkyUGRXB546ak8rU9hSWYoCTKAdlo/feIUvt91hs67X4ZWatNwSBWJhq8/GJDT7MN1aY4ob6xiu
+NxpdDanSLVNXnHRmGuiWibaegp51iAN1Y1gxOXFCDdHXSOZsemquKr45QeYosKw/ixo2HbnLL4b
JFwvrFb9crV991v197ffr05cs9/XSDnLF/V3yclp0bNs0CpcYH6/BglXXGXfBMc7uf+Ognza1lrK
o7cuNiOUPTwkmnq1/f8Dub1lIVQZluLm+nW2EjUx62FrMxF/ja+sYEnLBl/Ml1lDfbjqC8AOkImu
sA7VRPz/njoOMmuV/nVQtZEKu/mp311DzrQJe2Xy7Ryc3d8U+Llu9ulpXN5K8YF6ITy/3G7hLYOh
ayGm5kzxxQV4y1gHZjzmOW0riehAGzsH4DxmWyrQW8HItItgc60neXyRm/3Zkc1f9RD5p+k+GRV0
sr6X+We+U4inXXk9C53cjknUo8TL4q5OqKf3VY4gE58VcdqC3/CEIEvxcyhiBrTVvRtI27YcRncP
3Fh0XT0KOPg7DwWz3Np+6uuaXd1ZaELhRHeltHqRwGJTklRQpF9rDQygtB7yKPEisqODa3iRRcQW
TxvYabE/Ag8A6bkR2Wc8Pqsl2cbqOWBq3e0GwV07ocPaNKT7qI74p0WzPGuXGHwi2xJ5ple1q746
YhkSP+c8tXWg+pVZx+/+Gwt0N7Yw8Vow2K9WQ9UOu1huA0NP6KDW4/rJjxZYuME13POKiOvPthge
EmGn8rJZJflnxGaNAJF9jt5dC2FX73w88A2w8K4VW5yGD3eHCWF7r5ThcFQVH4CYpM/W1wkqV/hw
JF1Ijf8S2+XzXmxxbj1H//SBuBlnxV7wgpGuhS4Nrv5cdPuw2rcIMDYbO5JrCo524hKe+a3+1uRC
lTpNl57ZCUnYUNUFPEiyPrEy5zqpt4Mdbbs7R4P8kwFzPmhe4TKAk5WDdhj3Iaq0gsL0+gafqmdS
XZLx6UeFPiOW0Ds2f/6GyT9D5hmKAcPMh8zeayw9KuMQkarsHmhuoa1sr2vCs7BNPcLcOroAwmoR
ocZnkFrfAjznpwRFgbgFcHEHkqsYcGFQheX9aq5J9fl3E9S6HJ/EB5Vry0j6b0JtK6o94suzmPrP
9JlVt3XXbWH+PndE/5tRejUo3wg1cupeLligeA0ArY5BcnkNzMknEDbpwxuarlL33BqSNZ8xu0Ut
xix3zPHtI3PHv4pV/ct//mbWclij38c8vxiPuAoEInrESiFzRAZfT2UJCtHBAb7m1i/hsaev/2AL
yCBANr7tr3QuGM6VnCyI73Pcx2EnEStTjV0Okbbasu9aTHO5xe4UOlpeW/z2IJMgUdHOVo9uOx0W
+HlsmNAQ8AzTOxFYkUCEXL3nIOJduNSH+rSA94dAq0uhhvsD7mnsDKJXXO3oGhvjo1zGjjBi+oSV
nQR6RtaKdT3TqOq3ZZkyxqgj0dngsenrmlaOnt0Ca6QCYF0WJorr6Gjkftaxf8sk4x9yKXLyp8A0
Ln+yKtp46/nzWUBnYDaCtm1cv2+IVr1mOPwyZoQsK0wH8Q7eKgXZNCcYvyUjc27/jxYAJ0/y1HoW
3xbhpHp8jo3WcObwYcHSWYfHL7u54LPF2Hf27nR4Bj8FcLd6Dq1uC3UkFPs53A10/WTca1r1ek0a
pO8lN5ADaWPAhN1SyihJpbBNUFLRBTQmYybKtW5sNH/r8cDjGj1GJJos4AXEfgyy3Bf7dooRj13y
T2k/fa/W8dRc49WL++0WjWCqt2/OQDABYK36n4+LrELkosNWpXvU6J3+7+NTTX0fspj3csnntR9R
BcZoaeXVlypv27ddlDgC3W4Sfdkp+E6gFT3v4oD4BXfiVvVb6/67Y4ReRmlyIa6QrqVNapMCLm/g
7n9PT0cS/N+QoreqMNifdpPjzl9MafHW19pTPboVHWhW5oVk7XGQGgbYq5Xmrx7bpmwJOeALenN9
jbRiCgYgENAUQS1rYgt/pO1N9YIYiQlpZWqPlJXpQtLOnBu9887FOt0GqeCHGyoqcjYjjMMUdZh7
V+ofu66EW8Ipx8zCUqjXYvGimgq9IP/f9asGuzxyzDPuAR0NPNL8Q7sMuIhK6Brv9iyimvZnrX1o
K67c0CTlIsOV1e6F2cdDjQdTEHCq5KrH0V/SHZ6jE+Cb3Sl/NIUaGKlpnn4mEsH9K4KCTJ9i6Z+t
yQfpJtlm1iVNJnyUKo67SI4mBGE2Ffhn+C9JTvlzGQJk/D8VmYh7nTXFKRFGruMKlYJ6yGkEAHvA
e8XPiMkGuZ3IIJaA8mOJ9uYPBfY/GLoAT1MMOnTkPkZzWEN5WZKcTkHKUa5uRE+cKQXIDEf9Q/dX
FqdeLOCoP8z+YQKDg3IUygcu6nFAYKgG6vofpPv+hhDP60TxKXyKL3hha+RPD7oEKwuGepSmAQ0X
8LEZCJUt6Yor+0D5AhwCSDiw6wHJbHTOm4CbY4/QkGkKgjroxoO0/csucHZqJWiv+fQiFuzt2YBg
ED+K8zQHl9p5LytsL7Z4iq1gf+uuZ5ORPLVpT/1yUPgKIBYYJss9SE7oqcGPEgGKYBJROZhq9Eeo
npW/Y76WUTA2JhVvyVV5kKLI1CE3tTZT+xJs+Gy4sNYRpVbDun5ZxIY9FAEG6MCpThKsnnz8CYmj
IcghGtH4CtQck0NkkxQyNL3XBR7KBg3YNy0zxGYc3h41sqz2d7IkHjT4WCSqPg/1yBxQMfepL6Yz
jRgiws25Caf6GVSJV8gspjg7C/l5xYTt+sHM+GNo21oDL7/zHWeIjeSOxr3kewt194c8HEaqr8PD
wBibRgsoeVbd13YbdG2/iIqLcgBdbN9i9TVoaTy1qDixkHAxVxNJiFU64UfPOAGqjD1xxz9OSbgW
naZ8ytrcLhP7I1b7HDYjNnqRp260ys3OFuaCcYOo3nY03F3Kioc1boQhrEjT4Fmqj9cqXcTLhA5B
3eBYXsocqbJYkw0LIalgCL16AgvNNbtItiKKneNCHieAJowksoooy1sglbMFFQM9wSBIuC6QmIv3
bcLXUqLm2Kv0OA4KGZvl/en8EDeYJuFyfc9yyWaV8akD2XVBUe/Bw7MQ8rHrVOdSaxvxA9FehGB3
deblDdt59cqw9ljUuqzPeFkz4sHXMifR7F71BBvvAAbabAm+ZhZsHxrUA25QkVC1YuqYJzDt9IJZ
0GoPy55bjyKJYQUejDMrRVCIfWklLLzGtJVb06SmAzU7Zy2DRuC2twxPWpXkhXjhUC3QzbB+EA/u
GasC5vvq/akksJTU6Sbrzfb5IzIvJ6Q4C3Zhrf7lYPmgRmdp0LsAZ8r0D15SsLKfhyiUv/QqHtvc
k1kn1euJkXk0AXbP0eqkITsLekEXDbd8Wgpkq+CkjL9rNZltHP40DugNhNQqX9008fV4OXuNNcSv
aZHV6tELj95NdYtiPoA5mNMtpYf+o/jxjj5uAfRUinlgdyHOssUfPg+6j0+O12AWB1M9b2pCC5fq
TPyVbXVoqXfza8u2NAkn6cZMGBddOlgkTZlCC9htgsgRXqTP+jZgDbk+UevpNEAtHOYN7FDTuz5s
fn5lCCTboTe7KyispewVCisqWfhDmBUnFeEJVJIImocNVSbEEVlcJi5JwUVD8DvMX5oHC6YkfN4X
xVbgUBjuj3zHhl+Ox9j1Abk+3+l6pDfP0PUsGibgfbZMSH3wrImkv5p5iiNRtknxIPNEJB8nJhFh
nS0wd7aoX6iHZHyCCmLCIzDLeftFR5azAtJVT11KnWX6ouS0zT/Cn5q0q+o2B+KTfpACxeP3auDB
vGY3Cw2Cc7kpx39gyUk7idcF8e9H/bL6vCLamUdi+DrjiySgCgXfcSIEWf64mGe3KNwwHTIogfUD
ewRqyjc226UyYkGre0IjRhaJ6aCqrGxBBIlad3Ie2hQiAev7jtMeheRM90qJrKKQF0V7kgfRRYLl
pHvBc9ZIZ5nohubPxWRT7btPFzyTH9zzFUox5DujlVc1tST4c5NMM6IdScMa+mh5Utt+FHQq7Ev4
XhPdYisUxEDqLE1JwyvAGb3NfTtGfcKVznh3b+lQ0RqlAFP3QQYvSozyS7O//nMgZvd1CGtdIkxK
jRWTD/X0b5GPdgbywXiDsk+w/RfPHdM76dJb9pyPAOmsNLf/TnHZ1/7615zgZWqvdTD33QdeXzAY
/7yvCFP/71ejqH42TFnoAHxsvEvrsqc8HLrop+CPSsu2KTa0SCoq9Nc1fziTRmSa4Sk+0CH8sp/R
6ycfff9CEWxkvx3QE2dxC/MWi7Qb659tFOSU+52+FnaLhLeGI+eu7LDtjPswUHGd+bKoBkEMHcyT
DJb5130PZx0HFlmCtp3v3mfqXT0Lg76kHjWnk4dlSn7GXKS9k5nnI1qb7ywPrur2TyD8o4WwP8yX
zA3NMSUphVh/O+wo0VF9ls4/3BhoKKaQYITWdMBxRk8ZdkVyFNG1aAr+zRbY/NsXB+8uwpBhQgMm
WC7oYnIl3udmu7iY4VCKUbjBjo9rlJ4oSYKUy+gjtrltHNc1Yn0z8AXmu/Y1l7Qe4BT6DjV/55qn
OZp2ALJxihB2a9NlTTWIHMsMdg5unm9MToMT+cQCrdqOzrtBKJDD4PHY/BUZfkJDOa/xUYrxL4nE
y1UOqoESkEk2RvZUjqVZ4WuP0xGeSP5zZkf33wH60/8gUg5GMI7BIdw6VYBS9LzqMbnhH/4LbuvB
85Mk0qIx1/GsfAmIdvg6TqVn92qVjvc43PW1Echicf6nU8Kg2POQbW8R+tm9KmcpzdjMuFTqPLjQ
zXy8Lrah11KNW3ikx4sWNi9m6EYO5H7C/4siVFFpYwZKRnIqOY6wkVTCtrEK4ZBVWYv/el/eWVPy
Q2e+EI0A4uLCUeXevZJP22Lvf/37H1xfN0S3IJOf4HmgihRhhomYoBlnD4qlk1Z2sSfNqT4AJuW5
Z01IfJP+yHugcU7taaUe6nf8B0pPlHN3iSh0ecpA+VRyL3SkWY9+jhG0LGt/4AOBMMBXoOQCE7Xi
oBrUYYwqnw/5xPReoqGsh6Is4gRN+nXCPx1hDWnLtupsvPdRsu/CTsDuoL5bDj5NTyxGedwXZz7N
PgC3u2K4cTilxKAdq/TGGabP4v/96OH4cwo/Lbndy+v0cuE4fCqXiEKCWLh9OlKoBiswPPSOrvCe
53/VXr5V7mAp1aZWs9+hCSAF9Sg4erlU97P5Xa4ZXAb6UyLIfwuUtryuuOPjqhJCrCIBuU/HfQxj
qK2Xu2v2tAKYuyEfWC9lynZmQdH94WOIOjnQqYXf9acgHF/KbdRv8KKFXs5V2ydBiLkfB0a+6Q1s
l2QV0jUabsctezuGXLJOpSNHfuC7XWArbX6VCLeagNA5ujR45CGca3V8XDBrhaIlK0P07AWp4m0T
YP0EzuFsio+sfrwmyBz4KN20JLfPjdBtjMjpqsptUZJqJajJ5+kmYjnJpvsRs+DlSe7CBqOWY31F
eDvJx70CCOnXwcKJ5rnDviEgcv3LpAfViVBDLsOzsK05SO9DPBwzAnpw+zgZDngx7aPdXFZa1I3N
Ub83aXISWuG7UosjhdTeZD7qSE7NfbzVqP/CFNwLRG67MPQcKIKg0JtRC03rnTdLGrVRrYbCL7ht
KRrJ2duoyUthnUQARHSZ165Y7xroVG6bVMLIKvs3JgEOkZLm6HU4fvLBQwLh/kNUtqj1zobSwOO/
nBMKFxBMX+SuF7vJQmatim+VmJpxa0FrstUhmjNlYbRKYfINJKTtx9dniPGuqXHI8rB7wBeLP1SV
eo59srGhQjiSET1MZmyq8UUF6/9Ceho5FB3NsoJc5f0b6WTPy4KwmPa5YgmVLhxpyHi+X0dfk6Ve
NUW5VGqsKXQ5AMF9uyj2p54Fqihv+xFkqTe/PjqTwlpCeIsspWceqZSvBe11OcPSvN+EQiAcFXjM
YqnttzKxCcecbOZU1f8zZxh8qbP8wEVDdAmdtBRUuaGLW5wfs6QnxtsBLU7b5VyALfgpF9gObEUw
3ElCxhp3FoYcg8ISRV78DD1eAGNqt+tOoXZRdUtfltaL+/qpp9uMtTjuuLXlYPbljnB4D7E2afmR
Hb8jDquPB9ri1sxt+Bs84DUFSJhoCOq9Ftj5211WUPaHo/bSm9tpa1Cgbs/E2plP6cDxp1106ajI
FhRK6vXmBQObsEXtCZK96unHmFisSZPJcogtDJ2TcPhbWrHq0xMoFMiBqDzv2tH0xPZI4jrNJk10
D0YfAhirKauOSab1Hpa7v0XDG+G2y+NbqV14hGLyfB+I06xcAAzuzAAgEOMCZv2+UJZ8w/rivq0m
UFzv+iw0D8CeS81TR32S/WvvxzOwkGbZdDjvFAvNeiOcuVAttDqUuFp3MbLEhsqFbt7NH6Go426z
PdyyBxGHLZec8gNCSO66qptKWtG/+uOQSnwLBVcGXzpNZnWBnQPsnnJysfTV0zFnWEQaUYrGliT2
GDredTz+lD/5oMwQM8SAqY6Zctpt8SKhQzyBCPs9kVU/60FsvCVMtbeD0tGx1Ysqb/BSJn/E2+Bi
NNWyfAMurvaqtHux22XGgjnNNUoY+HqY50VarwwlqhxLPcy9I+ivmKtPY4nNs/PLtHK+y970A2uh
v/oK1JEc7BodXO2UTSHACjA0L4IDH9CFN30F78jmWoBEzrW1kmD87QxGtZ4QkZXqQ8x5BBrwortq
VH/f5TSAJF6qHZ5Pm0WT/trNTUPouudvD0XaSodGEPqLQUFm4+SuxRm8ILcZmdcyVj1ros5B4QxW
j1d2+9bsLvEJVzKtMENH14p0hscvFu8TcZP45tsoY01nZ+fZn6roLkEE7GdTnDiI+lXOktLHgd13
fflna0VC0y8/mgVbvtig/lgmaJT35WyCdHKrlrUhZqR9dqY5qMsXhhEaT1rULOu2wR9TEDnKYB0k
63oAHdf66PNJHL3SyBVUOtJRBOZ0Jow/MKg+IKktSKujHpH6X+IVyK9NUtXFC/G0pdM9zLHc1xLS
cegOtE3m/37/IJ29d+cH0+TkoKhDDTv+kY5PAZ1C/ZQk04tX1ZxrTnfQSkt1lQFcpdkDyHoDSqWO
IRce8AnmbIyHRCj9J3AF1lOTHmZWgVKuQrfOH2XtWSxM+w7hb+HKE7qjWG9c77prmB2GfRm2K3XU
U7vOEEbFM9lSmeK+ln/3vgzdFM/WZqokT0uofmyB98bVNPyza+aEg8osYA28C5muv3E5D/1PlqS4
l4NRGmZH8At+dMkEJ270oec5weeqWPwmD/P4ttA0Pt6ueA1j6/F6ZoN6KgwO8DqDgRfzSFMQvkqw
m7tRmbVD+OVeCgXozKr/90EKWrAKhndcql3MarLbccvB54lyKbkjVEkDiDv3CloK5Lnbi/kTqVYB
fZjpzGBW8HXlB7IZlz1xw+l06GjMBJzKQ18dNGYolbdT43MoZpKS4vPvOWdjuqi7KNsCT3iLz/3S
aCHadM7aHpQn+4CiGVXch/U16n6fBrP68WURtPrqWXN/mzmcTQEEjgnBC0BtWAZrplrK3g7q5Uzc
YILQWkknN0LA2OxkqAUcFA+aK0MikHH1QfDeEt08M4Lwti2ZatKbqZ9R2YUjiXC0PNzBJMcnsqHV
ixgRDxlvdYYTogoYgCw+dlhliraF61dHhZIBbDyJtS/5rX/GjLpsQ2WginqKYvOuK3mGwxgOPZoD
FrUHNc0hv49J2/c+DRuOJBPe2VQFLYJCxQ4JwadR95LwSORFXGTIoGKSMgBWrFDx3uiI2TdWSH4X
sfGt4gxGoFTmjNg/0BEd61eG/vrypKuSNDEKHJqIXhl6JEcxbQfM+L3QPPqX+5OkS3MOSwAxcu4h
xOCwmzYkonQ3rOMDfAQcZMVnbpF4m1iKqfxWCpAkKE0a4+oEt3T/+gIUw5F6wL1flxTnRY+W/dfX
4VKo0DnmPY8wiq3WQbczp3FxoZ9Nnbg1AchUKeg8BFYwL3T6xgK+LTXnQbzI4OVPA4QC778qOQOT
Ou2k3+i/HEdb72ZcufnYMaUnzuEdAgdQc/oMFsxD2vWodZeNhyKyePFN3j8Kv6d0lBcLr4adZ9wn
egqldRy5/QXQfdMaZZc1IUz6EQGoqZva1PjHS8jRKqPYkwtmsV86yJ1gtdh5oh3CAIKL2NQEFGKw
jWr9Et4H6MY6/9BlzXKh9DlEqXUkHv61cvTDfOYevtG9zWIkBR76afuVzEre6wHWZRsowvI17eoM
k2LIvtfNH2cSJazPA1xcA/vmlCfEmni4S75KXrJWjo3aJTx2yGwn7K1o9My27Xx0/S7SgHGkjSk4
Wjl2HcgXg/Qtrak+OR1N5yPcRxzdiufrx+zzOJlZVTJSa7/qAUP95ZhLGuihEF9UVkmWB5QX+RJ2
qADGXBcA4ypEWrVU44ED4CrxXwNZhw4Zi/eh1Wp3x1pAapuePfXHLfB3tnIaY74WwN5200eWYTO7
KNYQw2XVmXoFFk5dwPSSBnKyClVxJKWvYf7L+wZVgWpbJ4ONs+n2pH5XQL2oLV1kzj2uLylRGbH4
sP+5XIH8i4L/+jpOSPb45zok9saRifZDTTIPcodsVpWe5G3zu+wpVl1bVZh8nbwTCa5C3t+Lx56h
98wgBjGhQ2NW2S5Qp46H8UPX40hW+d60YDjVBY3QXDyntnwaksZFWHuWXwGQShRLUq+tKNVTy5uy
0+rMEXLfcPj2CAXdmr/6RjZuhD5Te6AcL9l6G3vBwxyVx+nt3UtfEBQEmA7MyKrG8aD9ZDxVHf+v
7n4HE78aMdk+eHHhF73LfkbMmLCdVVejGhETRT21YrfB/YANoTGKf+jMquEPEVHYSorntbTeFIFp
2vbsqooxEHEui9Q1cGgj34zww+NwqfYIFC3KqjnRoCCJyhzPlGDWy44Kc0AJ7m8G4nHdVAqBkPDD
XvERam5Su8yui42QMl2/5XnVCGItwp1RePSsPzhbOpuR9U79R4iaDUlLdDAiC5nBaKu8RAA0mg2e
CjyuvDhV2RtUjL3OSta5v1D7ipM+9GyRkNyI0IrMMGCoVEKHZ6ssAnn87w383P6QKm2kWpRVDDnz
hyoljvxvRIgslNilPMav5U60P/Ugj10/bnvgLpLj4HK7GjSYMPqu6gco2Uih2Y/xx4BkanBtZx9v
k+Tkb0soW8OG5GeEwiOyQWOq7dcSkBBSMnleDF7/ftiedx1ZGJ2vxxjNJH5kyo8rNNHvJQzKOt2Q
yPVKKgOSG2sQuoMWRDhPZ4RZrTzOU78gbBlUwplq9UNOTdB1/ZFbix+XKIMlTg2SFM0RhmiaeHdV
sDWDgEqKBGCCMz9NNu+Cd9vIeqBNs1AXLTgnl6li4qUAlMBI9f+fq4/cxv1pjRJanP6RvGCJNaUB
C7txu9imzEE9WdIgSrKr0PuExvWnayaRElSELswuDiPO603DZnrQskY4XdGD4EHdsa1OzCXCrww4
nTB1KkfRNrQFKLdmB3WTx7sYp7oAt5ZevHTmDiFSu9dc1rmxvIPQW/WEr/6rJY7QQeclrRyOs5L+
kjrMyZXktyzTlIbuStRsts10A4hv6V0shO28OL0x9NwNfDsEF4H5EPWxOuJtebrwZwVeCdHW70M3
obnG7QftbgqSXjDiB55fmklSEU2e56o6h+aqF6kqWR+w+pqIMD2+KKyqWeLHuJ8Qh9LjBXU4bhO4
sl/uDUi9XYxPOogFmAqyQIuspddbfubmA4/uywC1P8qYC8AR2MfFQ0bp8QJpN0hm+Vf6KV6zXeDi
6/IOwvwEV8JcjN8JCn1/9Me7pfOjRs27Hhs1QgDe9AffZmQISMJEWG4g5qKLeVVP5LlJNlmFrCCZ
8Rm+C2Nl19s86IIGX/++Og3hN0m3G7uRHWbLlrWAgzH8KkC/+GLauYBOddjhNqzw2NiE8oYf1d3o
FSzhnK5SShXWY+UwwCv+ysxzDIhaFhFL0mIAQjPiFFE125lrOb3S5A0pXE3+aK3SG2mIh7muuSvv
EXWPhve8wVbfcr6/0pDPzO2fwXWTBhM0KK8lIC35LI8fQaNGugTY+aIjT4oOh+G9+jUEJbTfuk49
wmZEwl2EiYMdI/3b+hxkXZS3nBbX17j7chEUMnkaRCZDSaYDuFBjpg4xbq6pOhSEM/CBJwq2j/x1
ymOAAdjvZQC8tqlWuNA/Mg2paZIY6oFsclGlPEepdSW6oWVAvGynIXQyZewLbRqxYm+JC7P5M8ru
oUPVgIxyHB8+GD4Tpnc0FLCsnh+fbqh7kBEyaBCQhOWFp7YNfsOH0gzC84f3SYDkWP4O5EWIwr9U
lcXdXPnRfA8F++82OEL2qQ3968wEDexEPeqqqZ/PxgvmVQIRSxzOipN6DHJRNqbA1UVeMznCJ0HS
bE9bxDVWJGAe0J6N5o+NEjleEzC8uMGvj6M0LRvRjdF3uWuKj9OUH5ZLP0rqEeVqcaRfCj5W9sgb
Uqx97LWSrpZJ2GJHB5MhCUTxDpaX8gmamJ9ilDTCRpMlG03yxrNNVlTKofOGDlpkdVlYPkIVkIw9
sIkVF4XKFTB5YqAKdICCbH1OfQ7ocVeE28LiMDcncwo5kEFEzo6drxisZoAsmBWEaWfpv+JppOo2
ZytZZaR202znAL2T/5LOZRhGggdskCDp3Q5dFVo3yfeE5x3zYdAvNMLEW340LRL4fGdt9SBUcKMV
kCiHsyU2PMSkHFTNzU/vgYo0TNZzwnTosAR0wHLRNmsW2cw6SZRTieaqkGYKgSiTKJZPxaxLbXsE
9Xc84ve9a2gJrKy5LQRhSJwvhJlCIeYjZI5OPNgCGBeDiruLqn88BSiFqeFYZaPLYlUm7t6p3prj
jl1I/OwxqmhTLUdBVfNSCP6qXkUBNjYPLlPF6BtUVie9ORvjT/PL/G25/rauzBIj7j76Nx31cQuy
aKiQfbF8bX+BZzqforfATHU1O2Iw0zyoDyeniZUJXIwpJaqhwYyTPk7qwqH4J+ZPr4Uzv3sNv0Yg
/Qf/eq+d+rFOiJqmGSarXy+H6dpQWxCIlzjPkwQUFAznnpVBDtDKQnbXmo1Vc6FEHvea728xvd2t
pLwdnqsCsouDemnWAzPAII6AQa0Wx3UuX+qUJGlaG5lpyKmyr34q2e1ZImt8cCD4BNel8NzkwJou
T6wwwI/i344ycfugG8AjXop3CBbuE2yA//HUBoWkE4CVNz6HTzj/g4WOgBK0OlIFY8Fr+B2xTjIa
gN2kx0BFOQZO89FDCxQdZsPPy7e2zw4hyZx0HfAt7tOrLtP/gf6uRJ3JsmZ5cHbeQIYkXMiXn5Se
lcok2hga3jOs5ZDkwsfoyEM69dp7OGaTHBKo0M6vwQVLgY+IIOrPvSeEZ5B5g6x0+uUNiXVxnKc3
XATJcH9unmyfWmOct7GH/0Yh6CYIB8/uuQDPKuev0diUfVOCFAWr4CN3Ep0gl7vEecWoC3dSGZPq
TGXY4DcPA9ocbjTr6lAm4qywtfk469pPCMmmfBRdNuBeglERgj5vVHeG37IA6XX3j5IJvPsOzRCU
Cr+5Lz5IGHMJmzIyf5szHK0r/GWmjgleIMPUncy5CHZnMa+flThue4L55k+EyTjKz62jgW9GGft/
2QhpZZDRMWw6CpBB/L7pxwYopELaJGwOV8TWc38NJAES+F8wUj2aQi++fwdGk389lSCfVQs3GvZJ
4sTgaRbYAsfWsHFLHBCIS42KfP+1jAFQgNUQjFi00LaBryyglXxdny50Ek2ZsJfeEzbFNzZ9gvUm
HbC+elpTFuVoXiSMnA1A6T+LISLof2scnCqPPi5SBllHdVLhxzCb10Jo09tJHLL7O81Ld3hnpgjQ
5ZTtaFsjgWHHMTepve+SUQKC/g/syrbn3cMV13Ar6WJhAZMSX/IpQtKC4LCBZPMBG0Go+VlNO9le
ynNwcsttJ0Evw3GNIc3d8901N5YKFl3ixI7Bb6vPzIf8T0AamdD1TGudQbu5Em4mDidWNgaIBSXm
s+dEbcYCTWrCTdCID8xe3aVGIMFWMIBbN8e0mu1pbn9Juvt7+IVNIkIaajF6ASLTzHN5RzjJ5YvY
Jme8CqosFfWXrECyzoB/a6qnZoP2V91CytV6y7ZvE8a46arH/Tb/EOaxSWADWAJopWsFOuEwYsjL
dl6u3Gd+fXEbOlYyij6adMM0my0wmHP3jHDmzl3NEvFSjnwONGQt1YCj7LGb3EAm20uPsJ6S5tTb
JjVPel3u/28vDpkCuRcf+nDFg57H/nLgN8jNvddL6Wr18oK13sSGXtC/AUvIkgKxlWPBlH33iE27
lZt4ykRTHKgNA5JkVCocRX4n17u8gt9V78zAq1vfoO07FLig3yvGhIf8KosNJFFEMofmG9g4GjxC
xcBFlxFVzc38cGnwaXh0mgbdOKUL91uNhVraKGW0fPYwIV/w8TNAPQMJyl98RzXnIGD8XOkwKFsT
ksmGWYeQPgHTdIUkcvnWfDwe/sgPlF5BPy7ob3VxZoU2ofHqhkpehFCSaxcmIiCRDSCR06HSuz2T
CLjk5tLFmJ0E23scHVsZtEBrK1gwA5dA3/AYK0TAHmq7d/ICoj+kLjkckih2IyK2T1fl0dm6i+YX
eG7Dig3wL8cJ+mPG695i3g3sbsD7DF66zRXVt3BAguLVA3I9iwn9tUMfchlyH4EmNsDJMDYG6lpd
Gh2AIHdyfPuv25jeV3ZmTvYz4uebvfJENIm3vagwOJcZpHudX9Od7H1T4KxkU53RbU/ulcxmg0zQ
CHd/afE+95jgv5Vh6anZxgf6BV4FH8hHorAjoqHOJX6eQG7q5d9jkMysTs28VPBCKJA/4Owrqy9O
luKsMUzDY0R0wAHgDsW2/i5wICC3KGIKpJ38ucQj9azLNkvEpVJ6BMS/D0XrUu9+ubkEysqHPpeX
zbBTVVzWtv93lj7Yslv81k92P0d2nJxkdD+PD1aKSAAzT0UXHJtegebmZUuWCcb7MIXAVOd8EwUs
ANn2Z2j0TqJvGhTaCBIIAqBajv3GtfeLh1jUYpoOFHjss22Or++j0yjIvVOGcgDMfQPmYkGqDpxO
XrLvdEIJWLv/a20seVldH6ej7yxnaj2iDvDpoT7dufJVEhyJgi/wf0UqhMibh1emItzYYSeqirdi
Wr77XQpX1KKxGmeO59G5OObFVQFxDkzQFAIH/FxT8StjkmusrgTtmRc+8I+IE9EZmtBMWMC5wTvN
oqEp8H23UxucI2c7C7yA+bX2GYk2/4N4ybXjFsZ2r6QW1xwIaT+g0hbT00gpTz3qPQb6JCIPpqQL
hm62aazop4/dcpZ3ahrXohf/OONhkTgTf9e/Am/nHlxsxAUGx8WKUG2+V9UhDi0roxuR02414cB3
vdO3BchqKLtPY8fqWjsPqcjTvi+XWLAMP2xU2BQawnMRmheRweueg3flysv7T6lGHXw5GRW2RmBR
74jgV1RZ4/QAnPhALyB6+emIdPUXoIE+niTkQln4oeh0l67sRwkMJRj0TTMkSb6ctnhM86286fLq
E5dbIQhMnTYovo5u2kmC2bFS0Fouy98w0N6jcz0J123TeolYJy4cNJe6QYXi0qKR+3jyN7qvrJ9S
Mbsog6W8ESup4+ZNGpjYdLtfDSKeLPJQ8lWf+0FS867c18YoLgTs7J/88Nv516nMJy9IJMkRs3qn
Z67D9GPA/ywyhUYl2tfsmmOYgTMxm7AUKoMQbBb4UKuXaDs0f5lTk7XtmdG2aYyEiVtjGu8iCWeU
dcYf/l4CgFlA2p2oJdq1TjriKrG5aUilj9bddznsLAUBmUcxMJgJeLiArUPNnhmAiTP7k4WwN9wo
6/DxJjFZnQvUiJa/W6HOxb8CeNYQWZ3jOamTA28lZwgxX+7rBIapc+EbvY/TIESY7TQJC6iAhRFE
ZJvW8CUj9c0jAO+yCsvJgH7RLvlxGiPqaloEOBPUdsTO32pdhlFMqkZxlw1HFOKDzRJphjq8xsop
gnHUZ5nICEjEOPJJMTTfH92lUSAZjdh0OnnDoi4hE/QLfUHsZjyMzOWUskI46TziJcC3x1k/I9Gj
Jcrvr3H87oq7gHKx+7bPFkc/J8BuFZEhaK+TwujOm9yK+vCPfC4HoMn3KodVqfSGe7FpEcYoDIi8
QPbVlS8lD7ij9992KSdyXYk0NJr9r3WtIEuT7ZgfYMQHqmITL94fLDQUDF7VQCpt3jsu7hW3ESl1
TkphRZTMtT3f4G2i5AmDCObtQOYaZeBFrTv+A0T3ZAOAX2j7De9Yi4c36aYiJfPIvO8OtMlRJyLv
SfPoiHAa80a8EAO/8yeErCr/vTqo9DGp+4PVCGy7lp/IWzkoGHfu9K5KL+4+GDr2EjSLfpr9+9oZ
0d881t9UnutrWVh2UI3aerSKJ7bumreXugob4hyK5txGhV13IIst8KaOjBWhlWO/aALLtBlrgQvB
zBdIXC8hlaaggBxvRM7CpSlNFzZ9QFGeYXeAYQmm2Cw2NxeirjDJx7qMeMZ++0JllKLWW5l4pt/3
QMJz9zC9T3PtsU0wL8n6AGh0j2z1SBP7QKmSpq1oIiznB3aQyt+UZ0Y4RPL9Q7kdsWSdKv+XhLIh
17MZo2nPCtT55FMLrL9aJPx4zUywxr0iEUQ2lhvG06KSa2hrnveLzHTFrScr/zrSKYa/kLgmkQ1/
d/0ykNJWYfq9QKDqF1EjKeeACn6n9zDM2Ks8bl8GOFBVPEzjPljdueDmpt5Xax9YSHgjfDYTVlbX
qecNOyJIXe+TB9p3ZEx5myoQ2CXy2NP2Qq4DMermS9L710m0IAnw6QIToxIQFqi9dm/Wm7wBwW96
OawzPmRtqFTXGnzXA2LrlQcGApYi9EMZzV0d+iSr0SKRtVqs6HhjSvYv1o8eXGn5vJPi8GX5hOzT
gr0DaxvonY98dfgD/uLycM35BPhyXcQlo4PkeVcK6ay546Zi9sG+Ty1PzBQtog1PdS4K930HMxTh
abCdtBf6xPmHsnWUxxW4KnYfztgaZDzOoReIaRY59vHq3dr5Opzd24DKWnaL3kTYqYaDp3bfWnnW
qrkr9VXc3Z8mM9hhcV/ElTwc2oyN/rUXxzdAy/ONPSdku+WoZmgEPb4OKWt288axqhEdUVVXhufY
UXpro3ixc2/6lmz3U2OT2dTVX/lUaAr/2FJzJuuxzeOdzGFy+y9I6BN4byn9EpUPtI3oOJACwcud
1FSvxv2xgd8V0lodY0EH6lgfAbvLngmTbd8Gn6bcNNSss1TUIoZMkE8OnllIexHhtUtMiZcpisyN
HbSVOeEBFjX7IpYpTt7JODMFk/R/FIVYAcde6mBrUHS3DylEpL0+i2QNg1QxvIUDsOzvFRvOB3Ln
25ezZEfwN8QNpuZto6TFhZQaLSrTACUo+vkYqUi/vmKFple+0SA/N6JaFXMcMBPNVDb54N0aOkum
A4BqAXZFS8cBA6hcUThGAiS9MSAvK2gRG0sscxORIZXJiy26rcgpuR2LaK4M+48RtQxCA66/sBl4
CxdIGG/bsgYp9LO9H8SGM3pz1NVVbw5wJpSTYbNM4S8O89xZxhHR9XHy4+gsnVz9g9tVklXf3q7+
ITNEqhFA2iTmrj3g+J91NR5T2BjEKfBAQIaqtYJwguoeSOi18G4GHVL6h3aZtzEU1MLxGsTqfQCf
nWm4t5ZDoqn5nPT978ZITU4mInyqJjptvymzWmPzPHnFqUtpZiS4I4i+31H+5aiXrd1GUuqzPHAy
y91CsrBAlYUm+LOEFC1lAPkzyjEQIpPGt3LtFssp06vb1NjxIavh6wZRLKR8m+TUviawaO97mlvc
5n6fQSIg5SOfIJcKA6Nt5C4ucLEk0Ev+UGekXROlEccH7jRPss+IKegPyjWXH5EmrJzNFVSsUpBd
yhJPGJbk28qImS1eQqE3CIcjq0YtivvpcxGko6iUxHxotSqDLs2w/+roEMzc1F6nvqv8ya5p2XbO
ox09dMheBS+zZimVizbQCw1gi0Y3qDG00A/VgIaaaSXOVmjvdA3lOgt6lVzMfh1JwsD7UK5cbo3E
LZwmpIJJW5y7+/cEgdv7aOGWc/Uyz3vKa+RHlRCUczdLEyO6h/HzTm+n5NCmBDqpxYxjmmbVxdox
iBFVeTT1pN/xcgLV5/E1tsK1r8qfagNHCfNj7SMmBw/n+ijaWTIz+VX5BQ1LJJbgh+F8pWL7Huul
vfcth/wkQ0Z9VYkT+IqJ2dwkGfInYvF5RPvjuZKCvdMXa87K6UH4UmXMC8NO96oXhuJcA9J6mZWA
W6TkJoaeqYhJbqRz7jyU48keeoyLzX9KUTc444K9rC+wkLcjP8uMOrPnfKd3cVL3cJrw9xt17/p6
8shnm1fTok2722LeZcdz/HHG3sw6Eg31U2PTWq73Ohj+OElH5fYK+rLLARtoifei9smJE6RDFMKD
J/hQ98E0HV8ddke0rZeyKYnGrlx8tXBBUjNR30wRfDfJFqga13OVKCKl2mm8IODZhoaWuBTZSfsh
Gn3nrRxddWsWdzocaJN9RR5r8NJ0Z2rX4IB2muJGfTLIzx9OKRc7x/tkyALTWMNJXCEICBVp0BSn
jlRza6zcUA4XnDbz9lDFmDi+evY0uP4fg0In6Hchl/zQ+np+G5Yq38DyKaxlO9BOKNNOE6H/6vYZ
pG/Cg5LY+yUWh1KMfpZmvVwBtkD/WecxPcTEpqfzQoutLASMBV/RA2HV/BoDCko+ARWrCnZuBY0n
UeH3JJJliyfXbQBdTLf2RDP+l5r1/qEsJMSguXAFYIp0QTyejZ4MglEnV/SN/DnTNEKcLML0xh8F
6gCnO6l7YtS1kuII1WiOMOTqdrp1RjcnogahyuwX+/cQmXyK81uozmoRTKc625fj5xvNLuX4iWnx
ZiXVrHIHxZ48cKHk4tOpkpZdbW1tOXV1DO4qZx4lmTumlJH13Qto5YI/Fx+j/1KuCRpVOVk5PNeE
+9N3y+KQ72QTR/AWI2kdXagPOsQ2BEoLIhy6uel535EfLn3+MyGJsnhyuxFoGeMen94lYNNglO8/
IChWwkWYRzx8HlADG2/9jQoR5jRhEwvPwYWte8fs8y9UCT7WrJJE3+EDKJPExGaYt6eBx2Fkw4u6
6CPGVSNLGHll2v0vsoUEL9v09MyeBHucIU7fA0GhmpMW5VJSrfCHSro4l2ncmBMgNg+VI1YZ0+BF
uUGdIzlB9hXa9LdBXCKebTpZk4/6PwD7DXcUGH58uWpqW6K+d4ovmbbmvxnBRve3w20Ysu9GVYa2
zwXStedAw59WmJunCG48UpAqYdQ+49BWD3edi8jRhIn529giKmw2M/cPN28N4VNwb97z5nkcITct
549dQKYJ23cuFeiXk9X01rAhs/Uheq3WtKgN2THXEmvuVXDWTRfqsrOjf2PoHElLT3KTWeZsbqWX
qqEhAuKODoVpntXr+aMKAs4MzG/SdeHPI8GhydTfvPCXUm5oZUlrKiirZZRR33hNpX/T/oJss6h1
gruoy/I10YHt/gAhnU9wJuejye2Jx8LM5odlwvh7YvjTPoJQXNjvgtW+vM+lHy9dVl3m5RPNtVsn
tx0w5k2uqaMY0ysy3F4RYET7O4rwISu6V2aMQ6dhhIJTrtD0aDBOLvbGIgHZpvjEOY2X58ckkWhp
jPGDkgRXCwRPBJThzWj/V5LhHv46pPtsVdaMOLMuttfOgbopFmIhXvWCymeUB5iWpTrDfaiFIBDu
7Ayo+6obe2Dm8+ANHZ/pyHiIXna+mm9jdQm8WqknGa17Es+FfY+Zde72NXDWnk1funUBJM9rccM9
n1BBMVaKfazKlUyhTmQKvi2fdhVkjcmKFu0uSwM5Q0CMxxTowGQV2yyyim2DmbVyYorM3YBomLhF
wjReF+mxyirc5fbxvNRrbDj4IxmFphn4GmOuUzgP07u+4o0K+2yaf96DXuOmL0LCTXRkkL42+yf5
665QDGzoDgApbQ48PF1hiqu4z/E8rsJ753v58GdzeQRTXL2SbLWGYdrsmJYKaag50hsA1ucdr8px
G24sOQKUmS2xBljERGV8dn9BLXLUVML85GAF3OJJu3o3fIQAMALROMQWM+Z+hPFBRKCC6myUrUGg
E/chLAyePdyOJW4ipPFljMGwPjjQm+5odjd6I0b0j0ocxpzoohue4NqL3nfAr+JxhC0QLk9RZyd9
5+xpmsAsBSh+w+XJbIbv5XOWheBaqwOc4+/JID914Hdf9xU/wLLC9dEabyQ7H5AHg0zdoHknZTuX
vS5fXmz9ehKN419yCrnDaTsrNWFsGL5TvuastZWcar27ABUCGDic68z/h4TwB4QEBCayjiIXaaDW
XoPh/Fb2NRiBHBGl5+05UsBPzwwOqdvlPMYMPXCXxOhfOSil+9ZfJPci9W3lTZwl7Xth/Gx93jrt
HLSyAAUeA/dlulx1YK6JwmLPD1VE11/yORq/WHfQtTbxvZoV+8PY33cw3T0jv0QnVY/GPMHqu83t
gvDiLrFryKBaNcyR+GJnCkNFDzDPO4HeMcY/eH4d1EA6L54w7MKFEnFN0LfGUpG6u6RunfwhpAY/
SsPTfcSTmDIfrWBED+4uVsDW4ikzo10DenKXXrHFnOFHLOxBRJGGsUbDVA5ptPd/gvoXAegvnvey
ND+2hQ3X7HBAXwXwLRcxi8kc5SiUfdHHPK97YKoAPjL6Bb9kT8eNuWzZlZkQ4bFNtZVaPYPY3IgE
6Z8QDo7Uj+nPH+qatlZLIi7DiHocLH4Go1NIw98lhbUWWjOvGMtxBlpiJje/MW+l9CJRZFELr99z
aRlY/OIP+N9WS1XOLgDejPGuvtTftsC/5hALxseGujOmCd5VgLXI1p2DdS1iX76Eic2o56NmS2zL
DN9fOGNs6rxAEKwSOQTQP7vdaOnVr721rY0VKPMDHNqFU1p5tpfvUotlLg3wRffIY5xswcH5Kojj
SqfJOlCxD3fdCG1ytknmscbGZbJ7NgtblY63O0SSJ9KQBbXlChBHLSX55tvP2M9or1TasroMsSev
eTrYjk8JpsDdLoP4P1NVBWdd6u/Y6H5vhfyauuYHzC1FPQWuvskfTNMz8EH9KP+kKiEpJdUCAO56
AAHayhYqFY+X0fiuhxhgDTCC8M4lPa1TN2XK8szUqpznLvtnYR5mZ15/Np8IhGpXOe+QJxxtCJbN
npjEccimAMVOqwfzdfrzoLkVIydLl4GeQIgiufjRzKhcMQBqRfWfyvId6elyh8aDPLyRj6goEsZm
+DkkF3I7Zi7TGvvMVGINaYvd9TKXbxZ8WtfMfgxil/Gx5G5qgbTv5B2sKKnD1Hdx1qru3Bc5xLRO
e2EJNCGxng9IStldz5Bs/XFBW293MI8i2FJLswPNP3D1Ys1JqRTXiHpoqAAhYx4dE7oHeD30szud
c0ZN6L7TZ3qErLpFbZ+8SnNCg88TNkyLYBTwEsGeVMQM2k+4vaA6aPLxAORg0DgHHkaY308zc62a
1KuBBy2Z70hiSx76pvHbsdM87D/bb1ov2spGinCdZOQKGqqjYrFOloPyc4AbO1iQJrdFG1IYoXkj
ksQpI37O8NMbGhzzhADP9vYChIqB8WbvvcfkJVP82Sbe7hkUNfzws9H9M3ZhXMnBRGinJa4H93CB
vU7VwupI0DXhsQ1oD13H2lqZ5622L3iO/XAVynR1oQMxLL4cQMV/+7ppqNGwaMo+8LIv3/iFZz35
zuPNVEhbRin5wWnZ/MAvPJWEjgxxt0f6cMxBdDrkHIZPvRDCKTZ01rOzHMcfHtLYFEQGcr6WlGtE
MOpUSTZvJej505JvuRlnnK8Nd3XA5e+x8e7DYt9qhAvCdBX9TPW2oDXURyjxJ6Ac+Z6r9wzHtEho
CSb6c8OvhAfE5thwqSmH3cLYf4EzL8gjQMi97JcVeP2V9g0yuHvuwDqc0ZEvglnBYD0dEf9/oRW+
rUSqCmOQmkyK3DUJ3IpIdqu/dxaP91A3osUXgMmIcQuP+tvTPw3GdoZLMYH46ptURXUvwQ/tp6A9
GVk4frDiJG/+ZuTawXGReVrs0hJ5w5fSbCkmUNDbrS1DkUGrgXr2CSHX3Y6VwAsxpqr0UlIA9R0Y
VFKaywbeM8u6j6bgxuu1KbA2U283pauoErkxQdAxY+0cT18/u4D27WXx2Li0vXekXwO+xUhiLVSN
51XFibHJj+zhr22UlYaX3/63vL4DBDoZz5ElV+quv7PutxpRvKvoOmyP5aJCYoDvKNEGiH4gnWw1
FfJXwJ3FSEpZwY1z7T/+/FmDjjIjHvittSrrX19Gdyv1o+H1qXVRq/zCJykL4D6wy9vGqhS4w5gJ
YXAJMlEwHRjnxXYf6Xb0H9ghuyp1jvfxLmx49Y060R9pRYpXnL2FQRUj7LAnw2Cybf1K2PyZRRU7
049LTt8A5NHZ/MVMhlWE4nAmok6nsU8iGUBUPocJurOIh32qNJTiHl5WLlDuZDQ7V0IoHpRfj0S4
NEz1IvRALsSpnxUq9cO6eQI0Ce182vHyJ6S+Q6PMyHO/Eep7UWIp9jqKtnvTKzxS4Ug+ttQtriqx
/QklEYkj/dT039/0RJ0wXuYF7ulsiCFTDXUhu7FUE7GUGPJiCAPpeGKkrwEuOlaK3RXX3RnW8gAf
2S34w9qv3Zw6cMlt4DPkv+7OCOPLOilAeqLQAgBwXiUP28/eya1Sg1QywVsgehtsUy8WRpATXJjI
HJvJWYRSMOWBHP0byNka6wd35tM3dHS4xpeGTSR/byYOh9X77/+rrYv38VXTl5mAc6ZgDmnYr2xu
HItPK7fDMi2DroetxameQqXOUd/M8CB2XeeL+NhCrSpoYgnR2GiDZFYQW3Co1TJss1JgbfRHNe6T
GS3FFPUFZTmfiPpEqPWYlwrWHoLbdGRLtZrlOQKdjVXwVJW+gIKRksLSTyjB0KXRz6JIaOXaaaAq
W6mF3c9Z/fR8CsP9RDFd6ho/n7Byz/+9Ira5sjgNstHkOpv2CbxYBJBkR8GqVR6a6/DLC2XmLcOT
2gsJz+fp71c8+UhvjV7K9pFgGAe40ZmqmswArvxYMG3Acmto+BbsVjAX7F37gE7LoBZbSvuvNMgn
rHxEXef/UVKiNC6XMdxH6NH69WNtR4/QWoWE2PR+vdvEXQlwAAkU1btXFVs549Mr38bwJHhAI/hJ
Qr46t5NNclf7G9Bn9llECyvMcU3xOmtbfqQBK3jE+/IOzExHtlw/8iHrd11PnxMGEtZpLPQ7CE2u
mJAlK1AXNZCv53Pl5k2ywl2AKLIhUXMjNoE19aZ5PoN+1cdynfJnI180Dg8F58u0SG5mr8goj6in
GT5Kkdc1B49LM45JfWu4/XSd2MR46NFpauIMwk27p+hc2OkkKoggmovT8r36xj2TCl9tZaLG0Pgu
kIF2IZHLrV7QomRVs+ap0lpg+piSRE3g6HusaAiFl4YqWA0BKIo4O41Nj+d+arDgzNch82UbZlfO
GBxXhL7Nlyr2YTli7J1fHfL697Aeww1SgIjWPPEkhkxD7zM1h8EFWN58P/YryMnr738WdlmaGU0S
N9lEZveCnlfb2dMPaoQl2KiPR+nuOhnJM9bapkRdPyCRJV2w2HMGN3h9osDBX7qbDE4D8oDoAqrL
UZTtvcEPFGgJLi9nN5+rWcZHIj/Taz7ihAcQJJOji6wk+bjrNXkelfl1QbSoC6w0O1cBzoP4uGJ8
W/ypcHFTwj6KXtkn7oCbWjm5ODIwfeprMEGQ8so0PzEHDMIHPV01LALVv5Z8vQWp3trNfU1jr7s9
AoVrok639H/KuVLPHyTRruEXdkaRYtdYM9cNDZi75W7TqiB9Tg4gZn6L6wOerDjPAhIYideDmKyB
YfahzdfW+bjRVtVKLvbZR1nhdwiKjz7p57CuyzP1Y35PpsAW1vxupigefJGbRO3L3faiePhssT+9
mbIwXqI4FwC7VTxRqzn/UKwextngdOADZaTktImOe+6ndZH8vAZUhFHSe70YczLVw/z6NkCupCtA
ew9gSDaaHt11PjP6yamZSD2tlWKKo02UDOKxT3Fka1GaerxU9bePeu31gmmhRnEdoWBflNNfFC+u
JG+i6hQkYAQPP1QKTbVvaee95wweAraCE7nZBVamsLkw/Ies0MQnxlIWmCDml+nCO8HzoKfIGptL
RQVyDlUwac1X/KMlzuut3Ogg9mXGflB6xD+rTrJVUl3rGigRmKa+DRfJpLaQgKUd5n6v1AYm3lIA
JFsOB7/Er+Dxi+MT1Q23VtIeekI0nVHDL7suAuUMuL1oGq74KiaTIo3BtS4Rk8QW9xm+kFZOQfXz
k0g/g33ifs2v1Aipd1O2iiG++j4rQZoulruzBEAhK3aqYXLRhj4f9zwcpUNINVzn96veP11KjJoB
aXn3B+7g9kHmn7MtVekjj21tcU4pIt1+lEOSs/2HbRsdrZc0MkPo7N0hqFKf8CviX/FNkGNSh/Fi
1jFsIEithjz1TQ4ZLVagib58Kjn6isThvaa4BMbRQUQXCqGoNynl7AmXtWCNK0sl9Gp6R/fBFk/A
QJGv83kZl1wFz+dV3FSZJHlfdwy8nJb4dZ5pNgiKOLtyKRq0FQEHa8tcgR0rtU70K4IndnLtmjYv
csBFQ0IJkxXE9WABpI/K6Wr9z43BNsLNmkAoIRESnbQFWXvcVeptsis0PQZ8Orcd1WowPAapi+mI
F2mtfGMpGaeAUJILnQXeLLYdDLi5TZLRrRfWT0EnEbUmeyee/I5QB30cMH2VgAVwQFxgso3ooabv
j1ap0wnRJ6dlrFIkXUuxcHsqSQig2IuNsjhVjtbrDcYeOsL2o1lb9LUBlvPLXT7j+NlKiQBBiMLR
zs5wv9ewpWhP+3z8H0Gel6noYsWILO/B39HeZGYlauyGHb0W23igPt1ffi+0+T+uIAqy9zlnkT2W
cQtKfIgsEHs8lnm8TsagVpz5R/z42+SR58CNuF74s7SpM2ydNVFC8AuqAXXCRXf0Ltr1f06gan7m
73FjClxHimlk5E3Xlg+8pUgP0nykeDIa09VSR4nrQaUE+SnKDaBk9eNJSAuL8q655+76pVYde544
z0hJ3UsHBclzxTFb6nvT/9ogozWYKf/WTbIcvfAn1SFvIRf2A52qXg/aP+xJuEVuQBb3O1RhzQCG
s0PaUogclNtUfctZwLv9avqk5CDvGbDJ5A/YmIkZVJlp0rCBDt9D6a1AtQEJS75eaOSAtQcqMaq4
5pgOyLGaqKM14swn7kApxJhi/WebNO4UKkUKZ/I4XGllCSIXK2ZC/0JirDGRXWi24da54SFb296t
6evJcZLpnhTYoexr/5AofukKIMWz+IDHeCzbVmA648vlB+tjn46Vh473VKjh64jlbvgzcNRoabmX
rnlgzFRrKQfmQoF0OVW+mtck07Bzg489ccdtQ9Vv1kehz4fCTihFYNrRx8r0mFxLa3MxZy5q+DxB
lohpRtjXV/4X2NJod8YqY/h52fgNdIPVV+elIq6mPETKcbP+YJwR7NbCcVMtF+kfump6xZsyvG1m
dJLESViIQ5oZ927dR70hCyafvoJPSGrOzFKiA8ROyA2hVYiyYcmykhXzx/0TM3d3MdgYob7hIcjP
7wRR1X6df7QOrc+nU9Wj0imxWxddnz1U1mVvMhFDjr4ybqthYDRUuVuNh+TmiO4K9UQ5Tdu9FAbk
XZKtKY4kOb8DdZh3cuaGnezz88wWsNVLN3188/5FxmoHlZHAOAKLG1Sk6RQTtuxiVnmoOw0he1xp
2Zz+1y2ANDp26aSFxv51TgAoXj0xoaXoS14Auz6V2HeReTGtLbmVdFAig6GWAyuua7DWfyInAiwz
YMKM+ppMoO5mQQeIWfsM+9BpZCHgymvKOvzbTpllJetksQy4Rrbo44MN6vObUUQucCl1kpMmjg2c
y9FOZk+6yyC+siUgxSERWbQSy7Dj4DTI9gc3ckeuQaoipukfyQnmlyHXD21l5RG3+b07dYZxpmym
VPByDNgd02XqLJCSdd5rPgaSQIY/X0j4eVMuJSvU50MvO3yFwNUAfxmmq6YJ2yE70p9BUXOQmGEg
7NZSo+OYsjTfKiJHO9IvU3uhG1AaGFZDQHFQ9RuGpodqAMTWgT0yHCkBGjguReCjMDKSfF+Qc7HA
v9GUwWuFexG+MyYdLSTfr9HrYYnOAD1XB5ueBUafYl82JSjCMEi5IBOdwlJ95W/cQzjIV9nalFmc
IB/f+91J+KK2ipH0axR7T/M2GeR1vCiuUYA0VlIqkRES/6MdaLK8qfp+DQsGqrVg0eg4wuM1BkJ6
pPEy5lmtOMl+awYec6TNKzfZ2R+vt/1yN8haKRrZpY/5qPZDVV5j5EjbsRh5LXJ/NKQOZ+41Mx0G
ePK48Vxve74SsCw/k6k3uiAwN6Bbif/fjrsPTywohoaBTHr/2xn2FB0rIuKR+eA5K7PHkx5C96Il
N4pH8kOquBev6gnxFex4Dk4Yyp/4hje/PW/mSPtGzMhl7xXS5GcDdUQOsT2Rw7dDo04tu25vzi1s
3c3b5dC+cX9Hfn2jlKJPv2MQK/aIR0Sm1i9CnEF+OrkBzCCJZr8txRXiVZ4zvt9R1W+3xSl+4u8B
rK6hlnZbDlZcxJINDzUzQSp2a8wuuSpMleCdHNA2ZcQOdnegWVWFiSXR9JtMja67akJoU1taJnNA
Bokes3HUUTlqsmvqKaH7CXTteL+RFeEw8sBF9kxa9rKAQ0R/MPl6w0HVuZXs/O+OdnVJESVa28fv
rVbGfmEt4WME4gu1zXKIhD8LbS8n0cqzWdoLiAiEf/jZu21JYleOHjJQkxL1LVVx376noONPt06u
E7mNuyFXGgALFUVX82q+y8kf5cgpJW9uFpQKJVAjZ+oEEk4iIERX/LbbZ593lv4v0qVFDCj47tJw
2W+doRkNY0zD7FqgCekMBa/zEjEvAOuWuNKGHRt3GE89WktjuxOaIE6yXbwMaAzz9ByD8AmltNfz
fwOyw27MI8XR8heWaC9W1upcua4y/yPxsIl3yBnz8AfAn9MyWYH2cMa6cN8tpWwCGVuFD36YMpwj
UmHKkllEv2LfjkFUP9Q+/nXl8I/WSQcFVLeKme+HgDg4hMqx+Jpx+guTVdseQBk94FYCgByIhuj/
2P7LPK58kjLY+TrHbnMUJdo5uI3ag3ex3Rq8D3gcDHDShwSxskb0oPrgjKDmLtr0VL0Bt0Ld2Eeb
37Qfy2d68U+BIUHus00aR4cb3lTa27UUi9xqULNNEx3pAZSNbIX9OjDQ7dj+RvD8Gx7Sns7ecQHk
BXHCd8HLPCAR25+Z5FIc4bkKQOfv+Oe+ubL94tC0SGdAmbsimBPvLWV09v82YVmWvdy34uVsJq5+
OiLNkH6Tkpg0Ktwi33z30IVDpY4ddq/k7A2mFguOJ7zhUmcAi7kNINLDFJR2Mri9aotXFQ45m4tt
5cFowbIE3tzLvY3yMi+nCE2cfbkTjLQwyziW5pKVFLllEeQZ9S7i2PchTr/45JwIinNDRtaUg6Kg
cGlswk/ZPm1XKvUkLe2OtUf6Gtscorok78gW6zjhw4PWx3rG3G1VEnOjcI/xhu48e3+c18ByQ4gK
JoSSbO+xac8LaEwvZPupK0nGE9J5VPwqN/AL456TUSm7MyiIyITIdzPJsk9Lq0BNhEreNMHrWD78
Rbndty3/0py0Yl0l+YuJgK2ftHjKdW8+rovo6FkEJb5O9AqZsafpEjeoQaVm9pDepz4z70JF3O6A
LtnCYw/6VusvIYlMh6EAq8JRxo/8fqAoLR0PdO287Vm5ze5sL4LeU7QWK6ENPNT5iERJmNesiyFp
a9OJlDa8tsuvMDuFEy9dSwzckNd42WFUoN23KZZ4kpY3V+TmwYZ5A959NL1TkmfFLXfPdmWuxRua
K2B6Waxs80RSg1dNH0xOJ+UKRm1lvIZaloiFwLNI9kj5ot/IOAUXYiqyRmGpGhKOFOFJLC0/GvDj
39ymTVeRG6XafRSPiKyOGMKM040oZMjeqcsjmxlAclWmTHF7lTfyJBfI7/50e9MrojIbem/nPmbE
jLGtwCjNgupz771cSXtsV96StLRJ+DT6ZxX41HcwYlWLTRWlwJJS9MgVChmq2ZD7LLGtbmv3C7Bl
TCRD4yhG/A7u4f60HuzxB6/X9Bs6b5rwwILFPtyghRYJdJuDcrqSitWFKj+rvE2H33Pg2lE8zX1j
hARwmmbLNrKU717ER20c6zpeWqoIkYfboIPinLK7MA/JzmY31z2ti5wjbzqBvLD2oLgE5ZIfT+9t
XvjpLga6igsBhdya+/QAygon8sxj13QrxJfbYcUu2HJ58rY3qSN7wxj/cRMT3Z3CHUL2zqBteKdH
+hwcY2UxaOXoG26cDpVn3SmB+IKq5eA/zuAqOUjYsz4lj1GG5ddSkHiNoVyXfjFNKPs0rMGnVN7k
Oy5zUdn6saMKWVpzXo2DLEQ57QX4l8YDVxHBRkPrC9rYpKPygOFnrMvJb1Jm1GiGEp6Ihoh3gLx1
icFrPeFz4A7BVHALm05y24pK5XCfoGYlKgsi5Oo3W0y1evm4DF7J7hj56CYYHyvPkkdpOxJOFE6P
3Zz4pRj5AD2J7KRGKIdIWJFS7PeduR1uAJjEWt4SOj+xIM0F6QeKORZeOSLo+KZgPk2KFUYUX4/N
DWDidq6FhGGxHnJF6sFEltVL2kT3pSH8Io+0gji4cfu5QjOblqyhi+WLH5UzYsiWaD6CtDyZXkyn
iUKVT8BmJHJiM0NqlyoZmvTqBzJRNJIDXJofn94d4alW9T+rjm7QX9OSKl/oS7dMZxRmc3iuTk0H
wIGdFrLrezFY0x+HUqs+Ybo4TGfZCDqo51/atUYMfoR7hRVEgT885NETBkOo/sE88ddNeipI1nR4
x+AYwNYGKWx1XTKuIiEFWkeTq0G6GQuJGctCstuffNZls3JrJV9oWdBb/Yfa4Eo7+6iqWTbVxvCB
9UusK2O2gpcYzDfgmJ+7FnltYVzNS6rie8QHb6rfoiRG8XJIhWRE3AlYsLFIrx5Fwg2gysEB46cl
qZXMe0O6YbWvPpULWvpKN+yYomRUSa0020ZfYiOVoJGAH89qb+lsXIbRU2XVeFwG72eakvV2wEfE
d/+8ZF+BGBbFJfFW9q3d/iNrB/+k8MPnFcpJQwZwtfiAzVT9hJz3rsX68wm/yLhBYbFhG4NGN20s
xZ8DXseyOseR464hR2r07zhuRagEDV/G6J5cXrnXytAjRxIXWB7YJpALi98/xyT36i6nRTtfInFS
X31/8zVt1dCToqZW/PSwR+xggIWNxR98+i88PGTr2JACJ4dcxWXWrCGGKDxySvHMxhxsIOE0FPhQ
yiHjeBz2sF7avsFquTm5t/RLdWd3/a8hL/v6gfa2d5LALcLTmdDQbaqEeUs/UsdQV4qKMGJe+fIo
FrDL2PY9nGUeeuzFL+Cba7U7ZO9+70P1euO8jmFNgOngpkCD1j2K5RL+Esg4gcns6BuJDHkTTeKC
prpUcZQBDsBq2Mtty3LAbIfsdLLPJacqjuLOhwdOIO2j1TZ3aqyuk5D7iyMtLDeVxMtjOEwIgBiG
lkioImXQ+kp/ncxPs/vE1BEkh0PkOmMWVI59GjCqmA4Rfc3D1xGhi88j7yQMZ68o/WWt9aAP82mX
UhiyWiyy9U6Gx5f4SV91A4zgH4nkOC+pUuY6RQrDTYa7JsWeqE+eNK00jA5ksG652+MeALxWY7/J
f1gKzUdH+SQrgf5rbf0PIKzA16sJlwkvhfS+RD7nIhP348jyXkXx7JiNlaF9xtS3hpGr7W+PbIac
K+w9+67Vb35ONa1vgH9mV/6hjGviW61g0bW2A/G+AsiGuFKx0yHFCw07m65RaaqQQJqkFP/SAJnY
uKp73mngx+lHyGkcBMfpQHp0Je8/Y8InegHhfFUDnSe+Z9/fjf8NLHcxEoChmUrY+aXXDUktt1cQ
VLo2TiBp3Rle8YaocIa/D5czmAVq8fZlKVgIwZd3uoqJ405KJ+EOPKINx/M29mUOHGKsVZbEPrTv
edK4/f+9yZvl48uBkYF5tHQXb7iPZ0IgfgP3LRCxDFtsXfl06hUOhxayuz4NFytNyUeBCU0K/D0l
TRNvLJX67VhqAaC91CXEc8MWHllBcnSgkjExFUsGuoqrztpyFcWwpF4XvIg5ixYYdFOB0v3zx9qh
/YZ+2JZuIfh95bGsBnNRWXlSEMWJOphUJ+8PjAIGCfw6Fuq1vPnVJkz6Asa0xgtRpGoonB3b24FU
ZRhu/c7B5Tl3YQDAafCpADPuJHumxeTnpy5zQDQYbGmlfebHKG68t8E0D8n2DUiitFWVtX/HT/Kb
Y2yNWBvK1I/Pw6PDPvYViT15tT9q3WGYAIQnNXtPPpnXFIIKo/8ge9FMoDPiV9M6UStltLYYW3yj
mpy6ZBugcpGL3hsKASNUGApUn8+N67kGs6VelKddZz4MVP5zlRGRbGaUl353UpVXxe5OOn/tsQnm
i2KHJsQHg3YnfEKAWLXim232F+vvovsM1aBYUXVgKftud0w6mE2SYcT4+HaXOmYN2Z8Rz9gjXpaR
x2amFHIOvwxFh7PyHtxnxA7UHp4RPW44ZskkmfwvNyTg1hoszRLe0i6UJrkDrl7Az7KFcMDM0oG9
FqZ+Zq4ER1HSE4N7q4tenMqCjdpxkWKX9/0VSJnkkaEkjA2vvUAahei13GHUoEd9c1W3rwfWn4DT
0hYnZYLtF6JGmTWYMJRUU9CMtHlcPh4Y1K4mZrmxYBy4QkCoZ+5l5KJ+K14JA5IStJ/uw3w512aL
emSBEc57A/BHvnT8K6aOXshlGkudyx7jcuteAWrJD3G9Y/fqdx8hmVohNQzgsivdHBVIaCfARv+G
uTz0gYqHXc1iEFfaRnwn4HwoPcu5aGhG6ApPdYZiN+F+ArFypCIPh1Fh++QX1U/H76kgJNj8rpan
z8n1WCUYSmnKiX/+Ih+g8swiby+BsYsHIx4FRJLsH1xCujl1j/k5B7iljlhMFXRGqcnQx5SSyC/v
UJf0JX1GHjqoLm0C13wnHuUeIr4A3/mc8tir6onORQAfXp6BIYpCYORbeNjqHpCvMv5SzWUG/YDm
Lu3My+OnnAnY0Xpf9rTySMRbQFbOaoPJQkvdMJpyBjmiFx5WIC+7Q072WKLtYZjw43hctn1LWMn/
ra+XVt8Y9p1C4nu0CmsL7RlSv7A4FL97hRZNmhsZEJv7eazMU3BBPWAPdiOLga4WJoES4YfmDOJI
6h5nC/7y4lj2/xiXSBwEpljRNr73vIch6zSFZnv9tcHFdani1PbdBF3/aOJl+1R/Hxr8N1aslfyA
bYu0M21NkOJE6JxYRzt3ocZ9z3/SPRT/RKR0vPtRXdodi1FwcaT4zLkSGayd1B/N3a5fa1LFjYQa
8Q0QBJxCh4obxr0oljP0EZEZtlPbgokr1bgHQ1hWtIebk/d3/aw9e3OvMlsjIHXYntRqtSOR5xAa
Tx26VcgOKB4KwgFqI2Voc6S4Fp7Ii2h0YqV3w0eXvjQuGUFWAq7TmG4FGfkbU54myN+ttSvKHngG
1IsijJMR26aRJ5UBbbo2f0iClxYGY9TLDTWgwiqdMUGIYxzWXQnScnKNPB2BF6CIhtxIHlVazZkR
vX7Cf7Tygc9oFhngn71YaZS2qtkM91IMd8FTDyPFVG9lW89gAlB5g44opiD3xclaP1gR/z7OM6Rl
Rq9uAah1llaZAxQoLI0w4g8OVPdw+sNJHYZCzOQ085vEMv3edMZBFgF1k2PIKuY220U0hHUYVyDQ
uO8VjVnCjWJiClGHyOEqXTXyCHgYvFVVKP1R4dLFOAmW/f7MgCO5wMo89gGU5iviAfcjBOlTAuJS
p4IiEpMqhUkxP7EkOF1qCV/VauEvl41vpYj5wYVtaBeQFujPN54FHktYCudFfQKcdFOzqHCbZKkM
FRbopmV1LP6uRbZBa6HZKAiFXtKCiTZEfg/ytGxwBsSQtdmJXeGPRyW/wSB1+W3oHdHfc5MkuVp8
DI71JBHoFNyQk/Z3VIYdoXS89SANC6Fcv8MqaUbBYSukw+Cko7i/HSzrqkAIAAPjdlxgsclkdh6R
1N/aG0I71py3z52EndaGl8Tv8h5vKzkbvwlfpT8VBGe6/U9dexxsBDqWwDv9CT1jiuVi2Ubiw679
qpFaCUhhSDCWbxv6VkGotv6AcF042TGlWSbc303JaG2D5pEUZlBZOFYXJWVWHxPOWlmisLnHkto5
sg0iYBhYWijlUbqHs2bxTG8QiiAFDfDZj0xZHekLvKJKcPKmTDYdQ4aIFpDhHdO9KgxL3OlwP1UE
jm1NmrA9ZI12fDSx/7n06wmb2zSZHmIjWB78RDRd96Lo9dWa2kLwwBONydjitjtTIc5rj1WmhdHE
qx1oliUEifzpwXECUit5QX1geIuJ1CDRowiviQwVcJTWt0Jo3J0RJz3KgKiqmA8GVwDSo4oIFioO
pfljTbkD36sNh3bIVTvplBmbVwHrlOGjiFM2FpNqaYaRB0Zc9KxcHDNN1BtHtzqumwRw70yoMsWd
7hYwbRK1Nwj71nXdLtIlK4FbXGGwJ575EoJhVBniwhI/ZWpxe9DZrdn3EpO0xAc95BgsVzlAPPSa
WEA7lFETZe+unpNrNHmjmPCOCasZ1FCHMaSOw++ek8jdw71ybE19bNwiyZD0M4n9p3eKa//kskjO
Ms9WxyMWpkYLiLqlSwbQ6rjIyI/zCVQ0u4+Q0Ts6ydQhMEc+iwWkJnfmR3KZpI3komK5bMSUd3xB
iC3N52bmaUykrPFp0OrNs3hga3jIZe0tUn/lzGXfhVOboXq7vUb9RsSSfQpY3ey9rYpyCKHKncfJ
7VSPEd19Q+ptCTVrOmEXbE4Q66DCGXIFBR4P1vCZTLHBYj7DFTr0BFYqxJjSwFeq+UvPxRagoftA
9Dd0krQca+MD0jS391vYfyBEFvU961MotcQPQvRgdld1X7ZAnTyvpvv52NH87qQkfs+d05Jk6cx6
ojfEex5BrSrzNkTq2c+LZXqzkIqpkLGx9XPajBcCCzlThoBc0MjYySwg0wiIodoqjsTQfj69542Y
3HxsqKfHdkyasbDncMQxn52/UZYDwCQfp+PtxEe7hUhfKl4gIlNOeu0EtawBV2Wn25IZNSdpCTf1
i+Hw6EhuNzjf5sfcCNmCRgfXknXST9uOjaRIpsvP24kgFIKaSJOx/5x9WcYUayBAFtg18fPlBMRo
qeG6om2kKVkPAlzuB3d3khPzao5pD2lWxuGvdG5KDSvn6yRiGBYq1qtdGYnnKNoBW91oftKJfsEo
0H9GTHj3jvMDEdE8vOWs/TZErkzfDGs54noq2EKB7Ns9IPpWzJP5yAHiklTLQ8xxlETo4VEePtGO
kJk4PkIE1DQ1/6DKhPoNDJpEuTeJAhcjEaQPvhGn+0yDxaj3e0/phNFZ9H8HgiH7uhUUy0hAxMmJ
Svv9A04/sLyHm9qWi4fV1zkI4hLDdmJeARuik9IPH/U5P+fFt0iCuvnqLenVndyjrlP1+wz32DjD
O7C6pWiWzb9zLUefBAd9Q+ASXNqwwi8XKbaTZb1421MzSSb39F+ZfzTcLPQGGAzY2glfuMA/KFuW
wFtcd3JyilI4xluGopTbfCXhNzDW9jlEHeLRUgjagSEXrGDFvMLbU2NhYkg6NqdZlN+mBnG4oXuz
tV5gtOP9jTitL1esfN+F8GhUHieohmubwl51tJtmgL3MT/5lv6CU6We2w4bwnW969d0YviIr8Hsi
pxD+NlSGBfLsIqFrQm+L6FnwKq3cH3l+YkpS+OAr2ZzTLEUmG10E90Adizy7ImhsGs7f0eiWnqju
1TCBOI/2ufZyDYA1JWmlBn4tI/7X/GmAsWomhEarIqgGJun9CRciCrJ1VrH3J8NamUpgEUgVcCcq
y1L1mDs1R9UTLRMs86dVo+dI0+o1HFi1MaAFxBFRp8tapWT5VXvWmZE5/PDVZ/Gj21VO/6GGS3w7
/3TycC31B4jMlxiSjZqYFUCPtmIO7HNbIFAo7ba9KdXpEqyAjbXYdTR/PgOlgw3WCztl4y99OCHR
IkZqVi4ucY6XalkkCKKZwk9gOZB8QWfZtPQyCTKgE4uPUTmXyhrWcOrq6iuZ77bh9wRstKIzLRtQ
Om+/6GnKKp4c6eUkhFs/Bd1MWcXxrYI0X0UrPhnEfySVtK3+9rta7HfLH1UmXNFOSVv/ATmRbUct
3dhzRat6Xi13zXWzmgAy6lFIW0zXvcIWLTwD79Qgeut6DkmRjnlZcIH7CNSPuHUhtTANzB7rsfYV
+iHyo60Q0pYOmaOOQY4bTTCoS5ed3v9fL5VgiJHvGPqn+AXKerLRtyR8XVUBbAE6DwUgRnw/Ybb+
c+nNYPFfLPnzz76W9TaT7wSJXqhjaQjXawLJVClUyM239GZrpy+iuPHyWqViBLs2ZzM+CzIIDmp7
xl7MoEYD4pKvLHJzC4/z0iiAOW7mhWh4E/5NAOU56P+ECbp0dmMbEEepjW/hprXPPzkwJv19foRK
KorB+vmQ9LqyjtY1XjBOWJ0herYvihSrhA90Z5aE+aYllPX+TqTudpB7usRjGQdCTl9coUPj/FPJ
b0Kj4Fm8J2zIR17bSYM0R3UjI6OQuCLvPLc3BZn6uhmYEmU7eOCbXVMV30gc300gMjl3YvRugZVX
XpSrlPbQqjsZ+s75wvRghb3QDJx1wEDInpsxY+AwhAjVmfP1hPhYtuJTvJf0keqAHaSqKY0BvDKu
Q5C1kO25OKLTNciC0rkRvU0LFbzb24yeJaf20/jtWoEQp1Rqp9jGBQuMz4DDeeGXS4pM9thsHpb7
X5zU/SBNjPvCpeSFGWq7MgC5DRG5kT1155P3UvMM2KvOvdmkHUeriGWQOO3hTdby2uGX4SCq9V13
Z795X71YrPWxBuXsf3cvWm02AScYtZp6Ay+nCXZEkDW4ghXRfduGvrPkZKeyY+nqch/9MLVLvryI
SLX8Trjpw6yh5nP3PvL89RdLHONbY81lEIwPOorcdDpRfuEW67ljeBSeEeE5jByavmIgmaTsS3xG
kZzgIYDL4ifCI2UYCokxc9RwSUI0XuWnHfQu42uDlqfVZ3DOC4M+NZgWbBaEQ6PSHMsroc3u5CqB
ARwk0sHC3wA2qvQxWbOZUhstu6xEAO0tx65dd+a9AgAljltnTAcJTMGFrR5SQbNoB7MPTbvVf5Af
sSrNDQuIDIGnKgB6QiXOwt0enBx6TFOOkzAiE0t4IyGAGUU2tLRvs50OUICOqsWkToQ9oD2BDlT9
UbBw51bNZHFckl1MWF7SJIgS1cPH46185dsRDX8/DOAFv+8DusBmoUzYCOClb9LdEmXNJybFvUto
rdZcF1mkpfQX2Os4z5pfHpgMoTm//eStR480HwGU/Holya94iWACBI57yQHyPB+WOiNZKK9/Slrp
pI27J/2jQd4WSPaDAScRY7ZJXVm+JqNVAKh09QUywAmV6UJa1EuDirUwFpMKFxJtIngBceoMh2L/
7SuooP0Bohk/8lS7l5uwAmd8G9lmL4BB1gzDR8PgWMyCRwzn7HYbkm8EboRSDjOSpoMjDbIcB2l7
4nV0Wla9PlnBT07g8IdgZjLtMYXFPpClGKItw6fPWVV+m/1ijHavB5H5hP0TZuZIk0AmSPTDRTds
FINBfWvawOae+3erWCM3a+IO0LjmHlNyUtjFfnbKWnSXy4HzK1qFG7WmLfOzf+0Y4wssmZHgDofO
cjrVn6hXQjCpw2UlsYzE76e9qa7M842PlT1crFWCIdteVFvSgqvXeXVfvo88qmfHE9nU/vrdHKdS
8AeG+cAfjdSOQP8e0wZyHsHoJtIFCxj/7V11/aHmZrjJ8d/WrhYxEyGAFERQvzdqWoQokDa2vmX6
plqpaMEoSJ5oBpMe2690UdhzIPfNpD6AhCmjUwQT22uE7C/oaeI85YVNSk7dmGqUJxfizj90tgMt
7G7Efa27v9K4hEYVyoyWVl1CfIvRcE4SHkmhZUBll1AcKlNv+h4kbfqzkIW1V+PSnkJAyMxZVJKO
hrKwO2ZQRKtvBhSznVUnL0tQPYFmILLR2/bS7HZLDwqqnq/XdLfHHW8Eg2PX/h67ubnPHa7nyAvV
mrt9skPx5F7TQ4CwLjSK8kBFxV7qNXJkPxMJRbn0nqxESwkS5s0+SMvQoxYyniXFh0Zyr0FPtcnz
cjjRe8tN1hIVgG+ED3sdgQL0FbbtVassGxmpS2xfiVIqh2xOsNcM4JnC7QdKqCZ3ihn3ZOCrcVG7
hy8HqdpkANGB7nizS/GRLZ0AesCqXPsdKN0lV7K+dUG9uCrwzsqVFHQe35NKu7qxKPoGtoWZCYcR
BEnjNQAuroe9Fon3xqseUZrN82vFE56tfSdZ5/6Vjgot+C6ktg31poq+XQoNW9t2uh5F2VKg1UwF
72eIM9rFhNqXbOMRoqOOE7OE0T/FyhLyyyHh2rudhcFefhIaO7kulH57PvpZ9X40BEHIqtNTftUd
QnymzeIEjWcQGp0odcfp8pw3Qy0EA/zSy/OUPL/FycpFWvjwlyZf2wCOk3qc5KPNdHNLSsTSmci1
c3/IwApujGm2uQa3awRYNQ7hLbmG6nXY3/Fsv+t7UiyCkKpMGULkYYrMxQgweKKggaNlXp9KDX8k
1nMXA9GgYzSccXnWcQqGqM4V4hYgyHkwUdB3Rbo2YL3cK6qFlrrSPJ5n/GtH0O99lJoaUwjyO1QR
gKo+fUN7w/t693BZg1uVUzcpT9yMtpJG/VXi2tUNODgtAy4rIaW67ro01LSsCWzG6lG/yWGsNeXN
K6Xvt4sVKCmcK4WZIPx7JkkohPz3OND1kKHnPcGQYuIaSbdJRsgvrnaaJ5//7XeaJB6rf0cZLJJw
1Ahc3ggilqFsaLmD7bunnANgZzdINdY3SIzhEzoSYWscnBpfx4j6x55ejO0bQIWHXxqDFpWwu3og
Sdv6gO4qLSd5xJeNq6vhlaNYV7vsb812zXPGD8OFINec1Ed0zeSA6XG+a4u7NVd7PKfUKjaFhtLG
Vmay5ySZNdWp+7bHwJcZTvF69J75uSXseZ7vh0uk6z7WnNihHO7m+RBKgXCBcQWBlcjBMUN72ata
AELgiq+wzFb9eNu7vgjI7Go4dD186ck+EjovUlYmGHQQo8F++HodJ/zDL+BqBuDtC3PGdx6ioZg1
Ebi3M1efZ2rBIGMUByHJhhBFwCj9zAyonV48qvIT/74eTrMqMpOzOXHXq7mV7+3MNcqokDQZnmFf
bBQRcgP4tx+Z0qHB8VXyo3UCXk8B8D/t95y6oRqH1eAa2425ldIknL03MirMLpI5r7HAC6qGaVXC
ETYbXIvZAULZ1aioy+6uWJIq3dYlts0/QwZ0D8lLVOgW/ZjzawsNcG5chLbGZh4+iN5+fgdx6B9X
nLrQgNhQCx8XwnjubPSNo2TLMRWwSa/9z1gqMB05qqiAGLOn9kG8hTNku8368VnRFRue3o0I55rZ
wJ2TKL6o8mSp/e3qjJr9wK8w3M5i4Ns2M9Zp5evlxmTxci63IsBmpI5JOIXZP1Nr89B1upOzdUqx
RFo4/asQa2KBCvlAJAYcU7sfq6OJftizFK6rwTxst2oZah9K6kaRO2LxUe3gjUr3nF1GG/VG7Ihm
goLaiwbpDFw2bLgXEPfjMeaWcsvKNdAcnxBj2nzHYP4EQW4EVY2fRuyxUoytNN0fHINf2wfapqqe
byg1dSLlwTlZneWukGLL3cSmzLoJO4jPBd5On0vI6sYpmugMzC9QxydUcxWL59WaEsoqRgzHQ3eZ
lrvIbhSqeHqIbNhksmbctc6EzPc4ZVEJ2rqIACiUbOt13qE1APKjCBqKdMljZAcVyWMmZNrkSVkN
Mop26B+/Ks9Xqyc9hB/GlSRywSumN2KtXwCBPQejlJgRVy4kuyxFDEkSADgRFXoWbg1173FwH0lZ
u885+0/n6IukNCO3h+kmAXZuZ+v/VibrpVcGRieT0J8y3kirXypj4WMkzJHyqYaO31Br4tpJ/YJc
AWz8PpYbdRlmsn8+FnZc1jqI7tYIfinEBzeSeYp4Rzpa2yFPM3EE0HSgX1ifoxsg7X8fUdOZOlKB
92IECaEAnibGLl4nutN+04MDyPPE1W1bGAw7UiYY8iHs4T71afA9jlLeU+BDMfEFk2VhuhAmrLB4
G8BlmZLpt2UOJfJTOm7InetpNnHfvFFmfMj4TRWZZAIofj+f3sEJ+QLMDA0WvOumeC/LQMs+Bb1W
Id/gN+k0NczXBP+pGrPzGiuRXaa7ji3TGqTVyWo+4EnctkGRSCq1kIfNlCsJh7W956KnAS9BrUY8
CQv3w/O2j2wj9P4o3MpNey6y7BXkjuGqJqEXhuB+qu3MWQOiuf8XBugSRDHub/VkOWYaK+OMmq6r
4y1GaSsaWYOkfcyIMq2dQF+ESkBRyXddEEbErO29Qf+gZmae+FDGleqrC58FK2mCiRF5Q6lnIVFU
zdOx4c7ionaNJMIS4pgl4Z1/AbGY50xH5CrUOWd4LpZB1rHYKHt3a3ZyIH5h8nbtg+ZMOTfKASJl
FtA4uHf9znyThAv2nhR9d0qIsW/RLieQC5K312BwBTn8mQHEPeZynyeW62MMQzKo3R4WZAmmk3Rg
Nwae9/QH3wnJOeBpMh3x3AQU6w0tmcMe8d/azjMKX3FBuximx5O5VixkJp4snqRS6EGRol6Oq2hV
joLGvl7OKrhGijpAAejjpp8c2ViiFq11DqLAF/4/Pp2VykQhqGrL1SD7TYZCpvOyAy8LzYZ0L8i+
9g/bEV/njhxa9bjLqQbeqDkdZmiKesvkRFqt4JjhO6BWSq1R+ZbjJ1nd//IjJmutN0Thka8OLjLv
DoRxyZ33dnTGXkO8QgL6nUwxXdh2iMY5VV97t7EQPypLy2nVatw9NNznL4EbacgLTNQHplmTkjnC
i0HJ2LGLrm4EPGVDGQf8kGf0pAwOyXK1yq6kGdBHrTGWcLkw0yqYiO7ZfmUjWV76wErEcPmRJMUr
1LuaduwilBJdA+G1TkalkXIU+AFUjeqGNkag/epwUrAiPelN+u72DEAG53y0TSs7//z4AN+XAG7Y
T0BWmKtGxFdbb2rM4cFz1iBH7oJ86+/oDKf8I1qqSEJnEo5RxNDbDx/p31W+lUPxcmfKuY9BoZn6
9oMessBkuCHdOY9Le4JOzpyX6TJbbCMMjvMklXimofdlf0W8qcSTHhfTDYa++J23AxlMHJKoT67c
+dgYHUcggnElihBjQTTIb9DkPLwxrw7GPkO5rwyYOixRFyh54CjuYCDpdZuM8vHOyDygiv8Hq9fq
z6cOv5uh9g7XY3YBFWaP6BAbQACPm9DAPZgJxffqOcY2351Yv6lID8rc3C0EKXyFIksMhEBk1MlV
3Xb9jaoRRVrcLl6ty7cdR6PuFoJLneKv/Twt9KAG7bFPmP3z0LVoIWIaz+Omh/qYj+GvKS3f22MD
zeeBYDN8AqvumaVny5giWuzgd3Q6fgP9cz0bXLeNlwwFaBFIhuN1FL2fH1yBfWBsH27jmGibhYBj
Fi44C9ERbcCYe5tRDQNYW6WJkeE5VxDqFIW8CUCziczgvRlvnzgDT6FvFZoocgJVR/6epDwkveO1
Vu3XdzeKu/HWF4vOC2IrOMyLy1bojvEdXmnyAzB97j6jRhewQ2PuxpMk+SIHy39fXkZwI2irIGMY
tjCPeaZxpD9RF9zsTuKefLOSYIxDLx6HcnVY60S8KcXtvi/ZRzYRjxC0ApMylVd0nylkGDDYg5XV
+cFpmS8wVFf+J6ZoSC8dZqlZt8Oon9DaEPEyN/btRKa8Tkx23w5PhAhc8YyTPZ9wzBjp+f9wPkBL
HC8n9g8+i/x0JyVOaKRttgUOZMz3uMzsYZjGAMYgAPOOYsR4pdTz2UFP/BjGdsb6b/tsLqKLF7fw
YJ71pxZbZs+iXdXoLVQHo3wn9o3jMmceUxNGFD7nh98kZeQkdonsyNxR1JTbnmUFJFtYeSQ1YmVk
OEGNVk/LR+Zknp73tFl06q7IXztCiAeTIQ0wC1X7VAFc+jl+VQKQDFANervkri7LaDYXREuSv4om
7tu+U7tvJcPD3fAaAowJFv1v0IjWMmu8fgNg58uM6GcaqZnrZdwjDuzuEa9ojxIGT9R8bcD7Y77a
v6Jiz3r7mE4oa9ZNOR4EMQn/T+Bo7Bo6kCgj5yfyRWXoOGTpMnm6TpZLJQQOr9oPhiC/5EiZqZbp
OBzOBi3iSFqEGBg8n2OjrZJPjz8SUx1cArTeT4RN0yEkdqBs3uxI1bftw5YiAAKOHanUoBThcKft
K4fQgtZSqfBbAoHCijlHtfpm1SJHq93g/+qCHgQASjHKGHLDiO31zdDPwahfUmL4xq5m4TjcZhpX
apCXRzaR2/ZEjIkCkznFLUXy7cBhtm+7aYPKSj6TbeeaIlUsWYYNDVS9GjaQW1fb5851iIgLQIVY
GtPi1tpdWSTZYoMQbn/R8MvNqZgnbUNPs7Mc5/kvj+mbodGEOCkyUHmesUOVz7Ly9RdD+0Ol8Jk6
jhECwNKIlb9FmCp/Pp4vVVN846es1L5kobtVuVf7JqnIHOTi1QdE4tKmWIR7hvGOdzl7NWO1QXzE
5EB++XPQtli0fAcSojqdyzWYBdXgGyuSPpHYiSLseidIeHtDuujPFojWAd0yMpb8zYmAOCNQIFpM
MrdDpSW38IabmnD9gaawdfOS3FM81sBxg6N3egK3R8FqihriSqXskiYJm31DINgtXqZ9PRn53biV
LO2LQIX0p7e6h14I1t2kn+OQDD2tyYsH3m0h45mwjZTp+jhCX2tS7inPvby3QFFYWXLWFhw3o9Ds
Vp+qPgj64/t11BW2+NC1tLiEO+HjINNNYRc0T/a7yi2SPz4B/9n2zmXHie5H7sDXtHyVJoHR/GwR
KCvLq2IJfbnuXdTkQBqfQhrSQflyqBSzBZ3woI4+AlzaKXS5wTJtUC/xPuQaDOe4Zt9oCoJWLrit
2dCxFzjDZJqCghKpk6emgedRuQIhfoJydDol1MnBtdzesAeM3jtdWiGixPv5r3f1qS/4H4kurFMk
5lX1d24Y4j9TFOGFBgF5JW7K/poxwxbe3fbn1hxAFUV+OAT3woxCZUzQ2q6O113BrCo32kSB7fXH
d1xfqstANPcoH0thNz3AAzv+tnKqM0/nBPhtARWns8o7IosRxhfFfeO6MnXolHOo0HhlVZh2t9nB
QXzd3ucsK8cCeEyTjmcNmRS+P3cr92oqK1nj+fdQhyjP/ql3/WYOqcgpKQ/y08Z3BnP2vhIslf0W
7RjXVPn2sY1whsR7fgxFrxngjZr2x/KrYUuUB+AvHQ8J88dtzspOg3UADAC7lSVkFdVMHlF9r69A
n457fgUfT1j9ccSIafLGJFV6Wv0Xl1UgsaaMJ2UySYlK8WZiYtLfZ0Gq/cckPvepz/gVhwAesG4o
h/URnL6Ja2K9YJG42Bc4rTGEae3mE9fk5DZKVWhPQ0pxRTG+ppe45MQdsoBiXrSqDho5Y/CDUW78
hCLFMON0vOUTFfkFTMwCI5kbIcRc8BJUsoZAIaFK6/ngM7ZeoQ6EKhJ2b6hKf9hiDnTdUchH7tgv
8/yTJX8jIXBvL0KHNyjAP5yQLrSZNRTJxWVfi3QySa1iwcbnP8D+ctFi/0rA7X5f8F/s4obRWFFg
M0ovH06FKo16vMr7bNHucpOhKNfIm/H0oz12CuJ4GH8qOlW89aV5RaNgeDiWU9mXQWbESFLTYbkZ
JImo961n7SYjrHQ45t1wnYxGS0vWaitT2bIJbcnH1pl11DttMxezwDkkBYx1KIr/VM0cDDBuA481
1pg8rEtPqA8xrbeStPrFQ+HcqRU82IwASXvGWF32neNIobGGQKVO0eWW5xMbFBUsLD6mzIl/cznx
ze2V/4YjbOUyuaf1795doEG6FVMfxe13sDS0rzZfijcaD+ORBuFrIoLXoG1/7aOrWH5SiL2Dve91
n90Z02TE5tPLOg214DiwiIVUSi0vEQmDp2enpIdEfDZ5jWwMUZkn8uWOIXauSIGbTUOXauUIJpGp
9Hct7LN7zMtlqP9jN4kOmb1pHCErIpIHqe4nf/HhBoEHfooVeW7ttW1GKw0cwWCwFf6Rp+pySUap
Va6b/VDpnq5N6uAO1nCQqG+H0KpUqkcz/vdzIpE3d8lc1WSA1Ylp1Yr9Bni8d9z+rdVIb4aSI3MK
qXFZindla3h/n7S4xd4LGKMB53FGwJ94PMqUnJyb8bxbLZhQDBaKiaK2sSSPF+rv1AadWnYYyIvH
iRLNmXSYcvRBWh0DP5uHqYJerwu0xQw9942RynQa9LKIXTdXv+aFA0Ub6plSa0AoHZ/wSSz/zTjc
RFp8tLdNR97BMNPUE2VMz7/NAt6JwztD9BsCMFPyYuF4L4H9V1p5kCv6pTObzRFJLUUEQgm6t8Wl
OrJOncSKi1PePK+kFb1NdUEFn+Xy/frJUODSRt1W5bEjr6GuDq9hFyJpk8WDaoTgaPp1Xe8vcC4Q
3P3NjO2xj5cj8ht6mXjfR6gCjj6ae5yxc7JGLIL9QI/4mQo7hTGhd+j3iDBxVZDMW0ybHMON9WFG
eFxdMAynkpmRMasrJcH64OpIPTrSGycgkQHDGJ0fS87OFy/bEWFJr5DmmZAB2QLXr5kt+ZodxtjO
RIeg2+9RkUC93bj4Wx23T6CMNnhDkn1IRrl+s4ocSx45juYkq1CaquajDVaxKdnMKrYlv7X5b0OK
w0v2QEkl+64Wb9rJUYK1OcDfFVfRtTZqp/nW3tmIJxqcGHeQP9V673Z0NpRQbCZa6zeuTArfA/lS
vOL6y1GciJ3Px/sctbGRPNa2pX5CSHoFOTENSy6IWTuMEHO7tJRCxuHmTvST8I6Ttpq+6r0LL45I
PZTUCxhlgdSWMLeOL2TDVM1vNwRhKFODLhhEwDCxzqvJSBhFZRUfDemNAHYTCHEDtgk8txlJq+f3
ygSDzpMbs7EwqUIZrZ96BhBxlvOWqCaqt10JXMJSnLrnwuIltZYU74RhUV2VkQKW7fs7vfE+mNA6
BqUse95eomBCpKp5VFtjLzLM+Ekn3ThbrVkwzicD8ZWDGi7xNCDVnX9iFZ22yg==
`protect end_protected
