`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
JWiNsZQZM3oRdGRQYDXrkS9EenOIiABSTHbuLUzeq9B0+gpki0cAJUh4sFzvqfa9BxgHlR8Mr4M8
ffIhP7Cu0YV3yM69evWBkCiCwRVeHTIcYqN9UaqzgA5EIfm7nZQj4naVG4MN76EAC19FkHUMGKUi
6avivlwJSAiv1SylyU614pLiTD/DJ0CHLq96EDldr4ZB/vsu3esvcZ+EWLKi4jqGqFoD2SdPR8mi
MKvctoDyEzJZHh9aHFksqwLWdWufgTEbQgFmTvmu3ZFT598E9zAJtB74fycdb/xyNZj7ljKGeZxN
P6oFi7bwnq0Dmh7IeeE2amV1dwxlr921/ySpbA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="7uYLjsI7tDuSyFep/0vbKAO+Y0Q+psj6YOaE6eOjjOk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9872)
`protect data_block
8foYIE8qk9VoNJFGu/HiuRgY/tAnpf43l9dWIdb2nawxcY9KklqaigyUcm+8Xq2Z16SiGSJO0uaT
XkBmJPLEm6NJDkpG2iqdlcCyJBZJ8IjX+9owOTSHPc4NCytnGkX+3Bwi00rnDqjrQ6pEigQfqGIO
t+fXAHC9e/zGAh/q9cOaR0Hsr5+yf9/XgvNb0LvRyiMA7VMYi55nffqQa2JJ72FIkqk35VuZ2sid
djtBwAnpiWMamrm1ZT7JQ0zHRS5puiYYVKXKoya8oKbiG8iuf/rRrGlJ/JUDPI5FVZRldjZDfahk
KYQKlZQCmdroBMW+sqBnWDtWHdVCXvSt+nPN0OCqtCsgroMlKVLWEjb72z3WHQi1+3n7jMmLmS98
3hGDv1DIwbUlsNRzRAuhU86DTvm5p1jnH1dhAGAXyuYXT4W4Nj46En6pU3/83SJzP8A4jZ9fw/HA
4t0Dtu4x0P9Ju0XyYV7P3pluHDYAF4vKGG8vNw8DIkMiSem3BtpJfcZxMqlz6bxU77wdoO0Yzes2
vf3WYMQkJoehszRHoZzGt0A3baF8nQklOZuX4pCJ/QReFaEj+oq+3KpwmVatSrEHMubMWDuLTwtw
5jo/zKxCVwkZch5sftoWd2w10f5WQbL0GdKmBSl/t3OHATlAKnqU3C7aN57prF5ShF7UAuDzbfvF
yY95E99mJSL4jrHxVxY2B5Hp3ShVRt7OAzbBHRl5/lI+IBSEopSiewQ/HpQphPyeWaxegWaS5y1N
3sXLO23Hyw+itHCP3pS6otx1WBiFrHqBicWyPUocrt0j9mzkYfjtANDMDN0h0KBmZ3OMsLDmgve6
8YAgz9pi7Rg8PZ8o0PAP0dg+f3D1yFsYyZYNh59l8u72Rt+AtZmDmmVxK2H4F11aFlwX1/em3RWQ
Tv5cPsg19scFDPNl0L83v+5/TBVfFLrHP0ZEGg1MvrgVCVzw2NPhmamu5jJCEBbREn/PWkK1zJIG
n7d2AU7vQ0nh22GFEwiyY8+mcBIBqFzofTkcMFB0WEE4fsAKEFgrB8tdm9FPCtmTDTM0+GrTqKN+
B1DibgbY0kM1oXCbgADIhdakeCLmols7m3vQwb8YnMPUos5bRUZxeNJ/yLsc0q8BB1f5L6zfJG6V
ydABMZWgquSGXlnFy1NUiO1eiId5QX5wnaGiu66WekbC8r+C5VeJ2zEOVFt4KGPNdXDnbSmCpXDj
KmLiHIRZVFslN3aEzeSwFgV4zPr+p3QK17ZETA5qEgQb+2v5iqKYuPik+aQL0HWUM9uUSmZ/CxPx
7dpkquA2WS+mIP41jtMctQVegwepy9BmkKQJESvbZDpmI20YLTgK4JJnr4gFcRpEPp7D4fPPwHGT
44j2E7qnGUVEChDj3IzVj0IcaTFCo676nyVQJOcAEgImC3lunBAePheC6F1SjIEHtDUP9N77Wq3P
FyO+xhF2GfuA/wq4d1yKQtZMZEISNp9Fed/E+Z5NCVWRK7y/yTIK8lAz4G8Q4E6Njqq0ytz6KMWi
rvvnzVReOfGNJetWP3OOevEYUdkMpxVrld94+UnbUIisIMvP3Y1EzPl2ZASybsGxX4WAjITi3MSG
5z+7w2u5gJte7ckcobyXZJXrmUF3B9Ye1kQ9I8mUt70qIgkkG/dmqj9v13JPaYtUM+6ycAfVHID5
Qdh+DwNv/gX3xTxgrv6GrndaLW29I5Zy66AaVKO9jgnhc4/cla5xEQgSi3MlUB6JAzm9FbGJvUVF
Nt0VRBRvXF6bsuxnf3MR2Kb8zYMGYF5DZwHv52gfC7wZM4GNBBp9DYv6JHY5jGlGYbCc6pX71vbF
eUqfpsk3ndhvOUoaoUK7Fafbq0zmUw3Ux09AbwxCVVohljbu67MKVQ7AaWVnKVOiDcCTE2Zt0o1n
DvseIRutuIrDx2a4rYMe7OzXNXMRAuwbAwHLz4YlFcKm5DQZyoSgLo8v3x13Y4OXhwz9ZodzYAVc
CEYvyyUgtGwhN/7VLmU201e/wgodcMcadZDWz2hDH/nlJyrQsQiSTa2c/BN9QkbRPQP+LAQiCbhG
SmGaA5BGCih56CM12Uls3g5eJ3fvCvvSzXYr1MiXPxQ8qAxhof8SdZd3o7m93hNg10FBZSGOrrJE
SyYjq0d1/qjrT/yGeLXY2FN+YnZOQjSsdFio89v01kpn0H6Kz+4GWRJx9I1rvAsjRGBOOn56I7wr
PcjiNt9FhKy5lYvFlNylYaNxK50IYQPAeIQWtgP8tFU6etDh/hI2+ISsXfjbe+UwXDRPYYL8PR7q
VM2fyf2vE7b2UWt8HgWfiljfcFK3RT42MPUOOnr48b6Zw6VRPvRaQSh34Bd3unV9xOxMrXcRy8b3
v+oAfDFFYzpm0/+rNNmg8NNkRJKcNcZeyepuMVxUF2E+biQvIdTqedFrx7/OQRdtQe92qXIHEf9p
81BIvrIidBkSXmmo6125logYOn5WDKJFvQM6JFp3CLWRiqqrhxv0+e8etj50LQliKkd1vOemkf4W
FFygchIifhT3gcqWBAX+v9UrysSsobtEe/xElkT5S/nZD+9UIT1NG1DbFC1etDUxDYrlPf7lUvi0
ICMpBaqnqmrJS91GSno8H8GUOeBi7oGQMvKT77Bw0S8joYQADt8c7MCkIF9aKBK/p5i4cz1DBNBs
0ry9ptJCbJNKgyMhmlZnKmQi7KxMv7uoM8HjuEdwR0f7BVQBWxC1zrRuIFrMHxAp+TlNL1U0mzu4
BVSayYrF9Rob3WRtkiK5f+g8weyH7CT0Zalz0JCE+R+U8Ppqth/8UjKIsl+ftPxrm1aIHiaaeaiv
NcbiE6d5bjP4n1HfGFztpctfiIZ+BUDtXrgQhQSnZEtuObL1B0laIjT1LL8B89QVNyW6pDTeOOMo
QhlOmBI+YERGKZ6rLRUAADyxnsoSIH+x15IC/NAZEA9VetufaF58Fb1of8eBlQvdzOVlH+x2/vMK
79GY0euYcJeyZ9uct3iAUfApCRZ89fOCAttqNpy+wQFRLLMdeAJPHoR2yH/mwkWoH+FahpPqAfCc
7jlDYskEizlQUMwGIxsbn8/0k9wPLWEbhSRY1r3L8o128cM3vgxKKsYoi0GIH5wNx50PbU8F/Esc
p4HfHnpiCbFH0RAue/ibIyOieXC8v2hkDMEgF/WSuGhqcn1Lw4j403eCqo2YUKATdl721x6+0Jj5
d6kP50OBIgCz9oubzfSR772r+ZrkAhZAkLC/p51gnRGo2iYBuE25/ra65qm0Fid134wGKTAVHspG
RDrrbcS7Im6rECrLlBxCtTz8TxEbVtXSSdAxmgRIUNP/Aquxc86FAHDBCko7OLtAll7S/xNKTE5r
mAfD1Ys5r4L6PCqRMSsT+d04KqL69Xa93OruX8+WFJb/h03tzHQK+TjGqGN9eJnbMHxrLS1Tw2Mc
6my0DKFYXRO2oW5K33Wp6KR0qYdKA15YBGkgdSorRsPWF24btUX6p0FwHjuKPRJosjQ1C5T0NeHq
Q1D+FYyWvKF684UWFmLtUhlJ+EKNHjStBzwP22ZWuIGNm23SEXyEkgxHOdv+UZSwhb3rjVflvGXF
8VhHEATbanww8+o6E7cr1XOd8dXuU7mKApdmSURwidB220iRit2305HIdtQHXDuPsZrc008TRdJs
ktSKyieNWwp9XN7gkhe/hFXo++Ap0jjZFzflYnzBwOBwe2R7RNOdjVyGxWYlF8phMvVteNXN+UyU
uUg4cC7un8PZ8uy+HAvOAfwZVf+fF72QJr5vRxOOtb9T7nz1IguSJAmSRAf5oGhooQ8UCOKNtN+8
60tuq25SVIYcd+BH7ipZ78/KlgBzUxY7Mu3PSpXL88GEr3VzEmfXGpCyTvurO64HskD4FHyHRxPE
IAgL/Ywi+WCsRCNpX3HdIec+GyInrdIAEIiIy+JloCbeWE0jMDVZA7E3vnJ7CJlePGjqJN9viSj4
MBfsXMsW2HhI35L9ZI5HgwEv+nrs+Yx7B+sK5KxreSiHxG36qpYG5FPJYbUNd+9ONdvgEq4GOLQ7
oqHRiAXn6jc+sp/BCo3XnkYwpb0OfCwUBs9wy8a7nen9JDUpTuGesOfxPP1NU/qhR4esTtI+EeRf
awr7WUOR6rYQXhlz/q42wJZpbgRQ9s9wAiNLXnMoB6ckKiq/7WaE/3kRYC0tQaJvL3Xc0tmd6gRO
iFzZATVf9R76a75fl+jMtjPNXK/kyGKKR+LJwnv2a2tu+/9IHkxK8u66gBFJs5xhfHLjbsQKSYQ9
M4M8gMhpMhJ+J2FFgdRTVtp3wbb1co/hM5AVMclGhEByf6ehNKNt5zdrkvTSRwGPU+4rIIcxbZ20
pfRPjOnIAIHgDJsRBzElonS60yYfehCJfONupIgkvsPFtxBqUIWIbDhMvdrZXuNOG51onS7zlhXu
FDOeBVJ+7iOl4sw10IQtEympNDtNjes18d7WTwAf3w4kHQqLmL955elVLwiCZ7OcTMGf5UZE4cCH
d9RIiPZFE+QENeLjCdTMhpzBtBv+MuosTUMoVeyir+1V6RdgIkhuxWDYXUTAaqDFLQfGxeCNjxgr
Y9Ml/HPKcuNsKeJ6D3c93W1mRIY0msCnwf73ulyaPots5hlF/qfihnbVTCDlaohQloZ8x4vvlWDm
kmn7iztgk8eFDnAFH6pUpBgUiUqqRLnfmm+6rp9dICgxbgvJJwS3p24d/Eyhr1F3g7anbV2tE+lA
Tb4NZgAlBzoL6FyatJsspFph18k/XgKPUfntnKb70h/LUa8dmY88TfFZuuN/e04YM/IikV1mUWBd
8OUwcDjjigXbEk91ppTDtIT6lAgmFMWiSOsLPF3HJdQ4RyeC09M2MtJJ/t/yvf+ojbQAE+xYtjWT
rkwYF6dSoG/4CSLmK7UhSSRQYVO0pI/5H7kkuG+o9W4z9xXBM4oFJgd7LJbSbgs8K2cG5OTq+W6P
K9m53O/KrkPl9ySdy26pkzRmVLHiPm//KIT3oiItQsRnT/3BSTwvu0jTztMcLzkEUtZ8wUFcas8q
/A1diD1OflsuMSjlkdZoiHpSWfclqcMLmtc0aayq79ZQ139UILSubobYTDp+FGVwiXI7Ql4fvVPk
lsXxPTDh5aoblKlIJP7RNSuOfqJpmPyYF+QM6eHeoS0NqW6g2A5CCIrRR12xWsWfgJxOje7oAr1l
X6mNfUArGjLZS6nVowfNIguaw/mz8VYD6UlwtTyqZKEDUe6iHRTFvHG/loZrh8gKZfbvXEfsGSUy
AAy7oBqJSWnUM8Dw/zjpUZPpziybjivG604EIouiTt3KnTkyZtsGFBFia+r0aIu/QjzHfSqi8be3
jJgH4LWugESXZMehUWRCW5jma+/J4XBX4mAaLuvh90JmMomwx0TXBfXg80J87OuvrqU8Eef21dsx
KSRjGISwOEsdGLrYpq/aF/KvNOMM07YvLp7NIHMGSSdBPS4DRds9YogK4vo9zjTmyPjwlBa3JLtp
/eBXQkiF7+eQDaFX/J+/tRBjoIZaBGl9ILyMmMP45nJu5ALpK7ef29kU+At/ZcwwiznJYFptn26A
9ASU0M3A8wtygTHhIS8ZvsoNkzdlGS/a4JCQnC986Z49XOiyscNO/Fhu8L6DCB7fXueJxs/DeqLz
kFu47aGEaSW71QqHUQDtamOQ4aV2Xwzfhvm9LVw0+pxV2nRhwhKtDjQbbT7XKoiJWjOPNwns8pYi
j9eWgs1Pbis1+Zp1QpV39OZhwz21bWLsto4aXN8Vg3JcPpu9wDpMCzqJd34J8vrSKbGqjaBpjsz4
tQyANh0RxJhJtV8MfYJ+Sdfip1t3X5oNCOPoTG9V7BC6NUsBlXrO2zGbC5bMv4+OsBzHixvl+DQp
qh+tGM9FrV9Wfx21Q8miGDc3rKpcDLSMiocAR9gQO0p2z9gJGm+UCkC99JmKWcCleCLd3YHzYIH2
CFJIi/ymzW5GeCgG44A6xk1pn5wUYhvaEb78cFTf+ulp2ucREiePskK4bjT5NnAnc5pGOCMvNR8W
Xgfn1lJYE7bkKCw8TFEceLZR3dX3ohrb1uOi+GljS8LL6E0ooN6pQ8SF3MrDlJwZ1n6YeRodVu/B
4usy0e6gK8oOmtw9ciOcnvgoAS3WvLhF8bwMK6Odi0MYds7Vv9Q9PtlY6gyCoyAD9ww52Xe2bHJd
wCGZhswxbT8vvSfOjxOCl7A9KBQzgNIcw3ZgRb5bN51OMCjEYaQ+3CvnIM9TVOXMR4M0w0vzJZ/i
dMf1T06QetudlXhq9e2qvy+g2nf648aoia5DFikyaPFL2L8Pn9VF7u9RyWbpH7cDrzWqNobXYA5w
/UvYyefS43RrRh7wopysWdArUyHJ+n5aWuJu53ggjxXp6APpgORBh3493nFx0KCXWNa5XuSnMGE6
nY+fcZX+QO2ay3YFNLkX0hOGHJVH0nGdnGJWODZtx6b4A2tmfOdEmJdmBM8vNdC2kWSMCYXo2mnr
CHp1+Ai08ELGIffwIdigzh+k4cpndcRTl1uyg/QKj7PZmTiLpfcEORViHD+ZxW16+s1DJ8nd/GFG
q9xkAGUfAP3ENmJ0wlQUxMxuHddfHR3Zuufu5chAnA740LC2pJsej98fOneWqfbS31Dx07+Ka01F
o7UPOpAfQUkGT2WvarW4+8QTwrneyaeMSVIccc38vdKYqyfAz1MeEhhqLVj6j0JBzrZnr11J0V0d
G1c+pcdEZD1Bkh967uqyroP/4LEjRvcT5OHF+IarjUJy3l34Tvv3//xjy308y289wl+XmsXnf9/p
YqxxaczH4HFrCx1S9JDWl7c94mXxlI0uQ5aOxcLgYtLaAmpJXR3xjrKvwP8fEG5bz8AjTvqtjJF8
0V0AIfJB107xm9664kqLAEZH8zcSPTR1iNilG2ibgY0UXL1YRKElD3itzfsfKya1889BNEJA1uF8
Ldvm97xxUl9KLEkjY/pjTwR5r+z2t4DJAs8yfIHWQiudAhlE1ULvtMTuX+r3HeuAyKdPhGIzR0p2
O9g1mDvbA/zZ3Hnr8moCfo3VqEmZZzgqvqmkf9J4ISkp2wI/IMFfy8E0+BfzMretu19C5KyaES4o
aIWnph0Lk7kPgXd1bM2cMGynT72UzIQ6t53P0M3lRreboJeVu1MV3ut9hTKi+/GBd8DSiHnfbaSJ
mDbENeShxQABCbz/G6ruAkfPc52MIuNwxcXcXSnE6K+6xt6QQ8/Ug4EdKzDODKAE/h/JMKeBWbLo
8ha0lh+KZvSMA3wqgMB1NXUPE00gBYZ4h7S/zQnJ4ofIqfpnZYC2xENPXcbE3k+PhKUWsw1hv9un
e7EAuN5BB8J3XfBgEKDA7omC5a3MMJy/Yly6YlWE2gjacxgi3rYJxrw/DpuPcHcpy/IabU0eMnuP
pHC4mM5CLIzlt7saxUPmp5RacFc9pRmgjQRWqqUZ6RDEOVaqV82ysRDuKhgFXKSJL6cTwjVZuZlm
yExNoV72wNhMNTKt1FB/QAAOTCbBfFKJQsunH7pzARfQ81SzDl4niNgh7Mr5yzC+XSHHpB8YIlSj
EOCHycdgoqHpUpjeFCPC/8sVUb+xjxkGJ2qVp9pShht8R6wDCpCGysYU+Txe1wEF0PKk1W8/mG0L
+jaB5EX7HkcxtGzBRRNkEiMe+6kLK+BYPqwaj2PRXsE8Hd5jIYW9tEO46wCX4jmllB1v/7ntw78J
JXPhobJwdvxpHhoX5ZoRMSRwcKPABSkc1Ws73OIAXcPSZaeqeFYN7LqitRSux4NAvfLOq2yh0wWs
QdglPGckviLmSFguBYpVF7IxBPdB0uppawSPItYojc1PfzLfKktDD6Z8tag/tHboYIrhl/YQOwIu
My6sMGNAbO3mY9lCwpTWK2k4yR10uiCF8e8Ln+BN4nRcHH+CdPx81QyAfzh+3k1Xqab5V/rfNMVE
w78ZPTudzfHBEMtjJPt8Num4UD4bEZrUCkhcljdmNWWYjh+KMx5KFcLzXZKtTpC3iCiuGFA+V0wz
aT2YdWg9OAmV23PlmzBsYwyl0xFfPNQQKL5lf16kNkSGZWaVzs1KTMM4OTFdpp0vjz5XPVwkureO
J7RVw9SK6iOpfcnZV43cN0MBk1tbH1mysA8KZ15Yj0xXAIbhGw0HV41ZCdbN0uCPVDnTyPeRsmid
rFTpk2IKuSXuzQQ8S0FI9/yZbbHOZzZ8AMLuYM3hdhL/ECSRCdx1gge1wbN2xX2qnMJ25COJBS/F
ET1HIFzFwVnppYHUy7hbduYgSfLcwpVtdnzbKBFtpr4SA9IQVVHC9xmMTLZhgrAmBzRAeE86UKYr
Y14snIodX5K03X2E5xy4H1oSxTvWMWTK1JbnayjZhdQ4OwFVqKw2RZksS6FUndRm4ActkeQD4Wv9
CJEZsrJiUYG43MvULBW/LgS2rwzyoYhlzeQCfrYg2m+rW0jfXKT+qpEwNZKN96m0N50B4T572RjL
FeG/Cim1iKNDh2mbhUgikdoaJzBf9QKpbWN8/tXVIiGyUNWe8QrJ7vnBqlaVygf3nX+4w+V6SGOc
WK8xWhJkkzK+gSSiIFPui6XuRe7/OcGpGspw+L2wDzTr/uNA/JXEaOsktPMKId5yDrdqVYyLMoVs
5Nu6l78lbyQyyQ6Qmx3V9SrQc2/7BN5lzUC0ogBU+JWNvyyvjAVAU5GIseAZbRse6fcONHEkXP+t
4Ou7N93IpbI7P47QsqpBliem8Zdba19pC2OLOEp+o3GArMFddSAzWr10o1dlnO5kuSGnSQZUcI7w
3E/4qGOUNWJ8cNM4imCLFjgO+bF9mpgItEqYNbqCMiXjIpJNUAPUcKO2p1qkC01KvHkEXaj/q2Vn
F7Uhz99kwdCGmcNyPdLNTUcr8oiVUQ7EUbTs99MlGafAjmVVU5lfbRhLBh3+gMtt3EvebPyz+9ti
X/At5vrfSykJbvPWMtgq75oEsIlkXY9EBHurCGZdOi49vsvqUstFe15b4zUmHZPdSPVSTKTag/Gt
QdRo5qKSS4nzo3wPJAIGHVMCLAlwA+V5nH8r+OaBY0gD00nQlajGRgswNjaXx33gqI3xDftqqlr9
M72xzU5b/C7q2uR4dqrutrfPwCzVJQAKKHyfjQH37nV21gWYnDdjDs1Mo8i7E9O2Nv3JEL6kUTiP
iZz5F4OD/Feot9TBs9kcmWW/ogFMNzZ1+xpyuStHT4YgzngaaXELyXcIwk/X2N7t5GY+Wr94Df+2
rDSCcWdUOjI89XqD8kTIFKL4gOMEohvRyEELlSHDjdKh2cbjUVsPoxKeKK9YJtSAX7ocD1H+clej
ow9LlX/o7YoFPwJe7Hh5zm/OCCSAtHzQ9Tp+f9zVHTCg2blUAx+HK3rRlHxyqFgZP4wHL/c0I8E7
gzG2tJxL0AEeLRQFeScXMfMcGBli6MiZ/uHdxygxEMB6rQ8kDvPza1skbefUa3lAu/AS/Xfd6YDr
MWa6mJV+S57quNTIBNmzdZIMnCHZTBH7b5ljkuEBifIQ0IohnGd25qQq0ZaWLdkS9XxYRKaHotiR
4a0HofDyafMguiMs74HteF7ZekGDB0p7TEafjZsUN5FvTrNs2aH+I7MslZPEzs0BQHjvFoqQ5KUc
9pOs6JDtfRqG/lYLVhxB1NPzDSGSIcdhAwf1Y8sWvyZq549eoIL3nCuzUt97RkahvqJa5TktVHe+
ujNMzc03UOO2QJeduqT8Enlyr9Jt6C+TBGstJwRuGbwkU4ykEYt/vavQ4eQ2CKwWQhkH/5btQ6Dm
kbotW3A2KV/L9WpN7VZjTSSpgkdLE+ShZtaDdDNtzdW/HOKBmjcsGHBhy3FYFzqA1hSVCcMLvPPp
BkDu9/Ymf1lTDnJesZc6MlJQpqZknMG4esirY+tsewrOUC5XBz0PRsNOYhmua52xMVmCPDXaD4cY
FixYePlSP+G8Oh2pB2euThfoVDYMT6WivuKcKW7wZ3+DaBvsA5bFHy3xNRhbxmPb+HRPtv2MsMgS
p+kSN2hnHuMoUP6/GMRwDjpMcxRS/Vyn+AAYrQ1QfFfR2ehGYkgHEep3bl4h40eX2ggxh+LdhxEU
qf1G2A35GoCobFHV4RacIphu+4r3g28H3vAOn5oOVNyG1450nxaqyxOVl+y9TwhSUiaL0lGw1jCd
X+RDJzIoSHA6ZHNcp4iDwCtY+nrTudc4LmVlVdb9lFbdzVPrXBoOff7IsWMTUUXk0M3cJI6VAB06
g2/WnpxlVqrUfocj01bWQ77dCceWu3a6t+FIXwsHz4ESkEmxSguLpjj1IhMlEQg/4Cdl3f0uUJI9
667+BeDZsxN83BZNJq3BW2FK2SjOULv3d2zS9b6a4PDo61bJG3QmZO7kaLRXc3mmG82kyoxBUVEj
oA+WBFp7keVQnDMLF7NSub3HHiVcGkH/FppM8j4O2+qj2A+ndgBvizavLU5J3YO4dx3h10+oHYpS
QK1wJQLhM02+HuOA2ASyJZlDg1dGLw0wftwsc9fZJu5tg1OgPWamXRbGBQ9g+4bA5aTi0Mn8O5ud
PzgAu3J4igT27AjN3f1YW6qAwTXxau96M2ScmZw5voPFN1A1ztrznX8SVkJUl9f4km8LDzcVZL0I
nT2CljohycB8APhGuzUtZADMZBwyI6ItOG0hw+DydjsSesMUq9zGrnWotFgxX/a3x/pFziC5iFeM
+SlJ0l0Znwj5q+Qx2m4Zi/VBXyOwtwpRYXmcqMelXuoAWS4PfI8h6eKfPqBccfvm67obrZZdcAXI
0RVW9mGCm59P5J+ai/rFS1Q1j6oew/cCGiZKCt+7pYBWuC9u831k2uuC1gdbPePJu2vEOa7gSKWr
4j8rz0Qrend3SfjbydKbxUFuqltxLyV0JK1lsGIQyf9TqWt5EOk3pWC9IAc4073Jo3JI5MWfPFbu
0qPc52qGLSLp1yIvdoNK6TO5I7z2pL6/FVn7OHS71F2sQI+jo3g4zDoQz9KBtcCrVKb090RoXxA4
ACG+emeLSkcmf1fK6uBZ+E3P0JFR05wffeBigwdXq5Bhq+hfSfIEmBbmm6yWHN7Fva3VCzp3Khzf
k7GO48U5hXo8T2ayexEGrCBP6Srx+GZIbHs77v3gODyvPimSI1svalRElW4V+FUxVwEU8z48xm0s
AfEX0hyTcljNfgo4+Wz4G3bCAdZ6TF2ciquJMpUpftgTcCEvuNkU03wuvIcLq7nGA5qoUW7Zrglx
5zWF1my8AFtgZ3NCc4rNYqDXezbFEy4iDG+RI4D2FPV6D318bKLoB/NZRInbt2jT6akcnEVxpNP4
zuT177q12mDuzfoF8624E0En/26WmzE6KFfasmZfzNrH3yKGwW910M4VZsvofn5I83COOMd2iVsv
fqg1V2j0X2QqkI1hmjPM2sXuQ0XuA724VZKatIHvz80TxkFdbmI8BmncbtRzWUvf/erLyVYN6nXe
/c3kkDAhfMXSU7vp9ZZ4mYBeqKimJiG2LZRJgR7eAG5ZO9Dk+svv8ZDW+kfT8AdCvWgaRsae6kuT
q7w5BasvoVkR1FBUogng7dg30opKuKs79PnDEIIJp1f+bJsUaN2UNGvP3CtAfsfIrm6v8GG6W64b
U6rpjHrmwSg3o96tJunjKLICF+ounf4kEL0HQPyXOD/5J1BcM8hdkrGUedJoyktPP1jGMy8S0SM9
8MyEMhWvCcQdyUp1tZpsK/xm/uRuGmRftZ1fd+Bjf8l8QcjAbwDTRyFjZ+0GoiRTsxqqM4drL/OM
O/KBeklEzoJgp21HSPI2MF44cixRpx0Ds1DAi0tu8izpnnd9+eQWQ9FPqHTCUZUPwOSszvTQ0A7s
+YOYpaZ55IkrxhpkMjylRQkVaabXU9MtdI5nbvMpzIRCZ/3bKrj5mrD6B4ggfvQEL59+BQtFnLLL
hlzijuUZ6ZaBxLHlAkFnU+MLfik+g75k55VzJv/amZc75ZwfMvhWwiC5aFTiZ58fXq4czczLX2Dw
Fukb2u/+Qf1aBp4/cKNO3z2Rf4OyrHznmgBnPj+mL1lXn8I5FKJI8LZPEmRR+LhSTEBuDNMgHChF
is30cT+Mpfu6REVkC/vRyFRQjIV01LgUnO9JVbnC6Fsnv41NeSFGU+NZSHhH//wlH4XsA4PQ4qaV
BpS0gWmu0SfXmRUFQifP8Se/6lxK9NLinsEYsn3ScgI8kHNvaSt96XI+LvWrAvBWK3RqJaidUley
u7QsN7UWfQgTGI7WJxLLjF0166wJL//84E/klT1oHxUDnf8EIV+6tsJBM4/PDtb/0vveaf+kqwxa
P4vnoNNdxpV+qJlyj8l/EjIVJDPzjJX9zV1KXyppltUi/TFdbbh8ZEJHk5DnOMMgMSUASB24+Ceq
688qWwbJe2jpZi5smMuSZAAQDd+FN7SjAa3puQi5pV2SS9lRiVSWlEM2KV93a1NmF/+zv2v3xrS2
qUYem8hFJc3dyQB2Vnu9TUxlzfsWZVYJ8hM4TfP30lEG5IbTSPvKsJKknjVqQcuFzBFC17WkVNoi
T16e+53HfQDeJCg0hi8xLnk/tmN3l+QXLoijXEU4Y0rg6lnQ+mVXrBV9GaXw9vzvQJfzNH4999D4
jt+xHaz2ZYB4gjPwZGVt1poNca05wHpWEN0t74lMWRLF4N3/n4VFqe7qHbgoBkTdRdiu95EOeiDF
VMFAPW1vd5uxx+jft6UjyFCacOxy4xi/VkGtbbYS/32WNlvLk1bE4Cc9Ffw3/nDcGCFLJWA7CLt3
Ds8Pp2TeBEIQMC8ppLDo+ZQHsQZZ1aBb4pWglidsNwLxbaO1XSYeef/MfbXp6MmIr8gMyk4JwS5y
LPIK54Mq8F4Vqnl7ZD2XP05QWDWVsgXocOdv9q+Pg/mNLhrMUEGpeeorzkxmnLOGvEVzQDcLbQNp
vpxzdyCyOwq8DeeiwVrZBcx8OlUnNvEmxeRWL1Se/giaiuo4fqdtlv+tedQbV2A1lst32cQcjD4v
BqUheMhATkxgzfnPm8j3/Amuh43jvhZfFyvXISCzkTn3hoxuJDd4/1Dy/ImwBK/O80/l+pJbHRS7
mtYm5CrqfUHzOvGdW4ZTWzJ5Ds5TboiAVG9eaE0BnTXXcfxWWYsXmR8GFqtl8iK9VxlD2Uu8jHpw
Wqlh3CzUf06LbSsAJil1P8cg4xdrC7mM5eCJ2mXojuS+Vgd7OlANhg4onZyWomANf9XRX5AtIgbq
zEsOw/JtrgGvag0=
`protect end_protected
