`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
YEqOgGSbYpC1Ka0NBGqBGFNOyvAPuG2t95hbwU/u70M2/Ypp13OvmC6Oi1iHsJ7OwtaqhPBxN+VV
mSAg9Kg4g+/u7M3whNLZQmtNWwRJE/vcZUQQYG0RlQENqztm6zPFKlTFj7KG7tGB3MoVlUzeev5H
7TbrNX2EVawu+9UqYcl/YsRAB+yBkH0gUyuNPfysWdqQMmBWbZ/PxSEd5GSQIWkCG1Wm0AHolady
boIYPyveVbHywJ9gW2oAL37mx5ORn9DJw359uTFZV457MxAi1JfT7bvpEGHLRH3+K76ttxH2BIxj
Vk4cEd7XYI5VmBgcrMgwOAGHl/BFWv+UZqj5FA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="9Mi9F4ISeAQfOyMVLU39sUkDDpuGh6/CMO6nsxdcYAc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4928)
`protect data_block
AiZY/4j3QXBeH8o/X7w91gtn4IdjXoEvowRN7xglfyKr1Y5rt+mAR1B0Cl62dMAQLim3CDg9Fbt9
8O51I+xEeHAi5iW4LdCHGJPR645Hgbc4QyvYHlhDbdL/cVxWKVQ7j9Uts8+gbdM/kXgLUgYZcsyb
2YipjTCVC3WEZwBK9YH5GyBS4AjrbztV0Qyzjs2wJK3rtS4JlDJuhrQg2SYukKROgcHPUcIo01gX
zQma1twVXrlx+J4GiafdljSPFSFkDRTYAIvNSa2UXruS8/pNKNPPhkUc7714rK3r/6vkE9cabl2W
s8TelwHShhnOBFx9qXZw6u15fyKCO0TwAky8971nf+41acdpL8fowSKK+aRa/xQP8N1cKpHZMh0k
sgLCjPqhsnA+DcWSJaxpDYF4pQb6ViELYBMChQfkpSZEVFPbP+sJ0AlROLdb4UTAZSI4Q5Hoqy5e
iLqm48cFgBqfLJf+6NnbQU44MbgPfe7y+YXBfs6JvASyrUKhaYOpX//cSEW22rnjGDkEUWjYfpVU
05gCqhHmPyes7V5qhlfYA1YZqBVbaomQOXuRb9OI9urLY69EezMz5GamG+ysimEZaOTMWV7zDDXM
8IAcGuHDfX0goN+pRjLtw7bYIFOBJ/r6KpSXdSzUdAxtkBgLjGcf+MfhzC7tmSqXJER1wGUR13zf
f0LafO/qdi9dwvvyU8RF0JbYMxBTg88ZDKewBUjruMZDn2aNzMAocETKrbXpGZScFTZIFTA2ziQC
IRHnjkKT+AaqNyybcR3KWtt1Oc4eI35ZmROZECQbpUVvX4/dPM+AGoGAhA9p2drPmU6i/wXg+asu
xm+KLUSBAHLZFtNgxd3l7JzVY6ihoYZk5qwqflCXV4s1S6m70AQLvM8453rAa+hGMOW00VmDtOwA
ZQd+yjsDhY5gPyusQXbylHGKvOQFU4H1gNh0vpcJKK5z+jYzBsUwnGlrN082AuhCLPko/0hOkoZp
W+B241i/Y7IPZeHEeImwPHSt19dCF2kubPCyG1Q+K3+M/FJesk1onXo44WC/zlMkC/nyRnVJ8Lxh
Lv7nWboeHdylIzVlrN8tQI8Z5tqNxUsNB0rVIaGjU8DCapXa+mgZMc+OXcDxg7FWmLNFxcC2uKYg
8Em3aFHW5FvLb8NRR0HIWJajEYOsdl1mcKb/AEFJXoQ4ozvMeojrc8Hd8MTKEWC7hJL9NwZbxf6z
xjDCIAKMz9K4dOBZnT8wLPMhOL5HRQrpOI3FKXihy5JisGis2jhiFe0EdQ5kOOsZ0QaYO7vq5nU1
WfjIcicFbXrTxYtOGMxa5UrAeCEYQOS82kAYw/Os0HpHGHJgZMFDwCltRFzJ81KLQEsj/FTjHGXI
bmaShcH+kkMHJ7QJVe7N6Ibbd3vWurpKBenjo2wAIO7CJHJP617tEFNA6RPeskvOjjZVkQfLGZ+C
OrO0JnZMm89D6saLBHmzFaM2ixkBe/HgiSxMxuR7MmIyn73GSvToDTPrEndJVdXLm2+8txptADLk
8WmRPFiRUKfGO8rVGZrLgqxVL2rcP6YtVJUBS1u2+PMNbA2UALq8v//Kt9W+lb3CY6Y0N3OnyrRz
I6Fb3da78MddN+Qhb5xcxr2X6ulTPF1rEhkex+J84Grc1TinA5IlAh34zP2JtmM0KIbIO+IjlCN7
H4RYDVXUdeJjFM1jLOP5pKvIDcelo4iPtCZV8GRMHkWLgkYYAP4yRU6BR/Uni1xFIlZ3Ow36AbkM
YDupIhXEQqitr3di3da7eHxINnHO2vCudg3bEHEeEVEQ9NUHa9ws1WKoe+PNZXG7QvgNUuljFXit
YmMak3fK+0F2zEU3nzUrhPti5a0R1bA56h19govqMEf2SxrOVl3+qtCm/DVjDkZVUxOc+UBP+RrP
N/EmnTWfvcIbNtvyiFQFWRel5B7dgxguUoC7JrPTmPpY+9msFSM/jD630ve7Lt5rxpTxOrDpDBJN
zYSZZUY0KjEedlhi7Xsls+q62ToAmuZyTSCl8En4n6dbrfYX22oslPLPHW0DgpSJSiROmAWOLWuG
Q2Z/4kIc/ALaeoGaruncICGcrSFIdjwPUlzDrpnSzjr6hEbM0kttiWMQte747uzHbctCxfvM7PDj
xajwxpDAUc7ftm+oR/1uwLv99rD8W+nzkCYfnS9W6NniyAUiWXKmeOhAgg8HThQIthdOKZcFIE9X
HiZtXiMI7byqlQ1rbukHx5tmC6twPHE0Vg3sIunxpxuki78AFL3d/Vu1LVh9kHkx48eiyk4sKQGM
TXOFOYGKgcknXzlHQmG3tOHvZCTPK+tiREYxBNAcqBChNZ3ynh6VYyGoBYYRk9YA/DbEs2ueWXrX
j+3WZx+6bis/BQElZfxc04RlB6SPk/d6nunxop0NWRApS138++07pfiRkdv7jAfEE3cYKOC9YXA+
W0KSmvBhlSuDEQtPr6j9DhaeFFkYI/ylKF5e5Yq3jWZJP4xRgQcPDG802hd6cy1+NNciOHvTkITy
uEIak/AW/hb9UB7IcC8fdelwTDsr5VFVYc356Mj2Dt1tgaZCucaLxNMSE8Q+1xq5dL6Gi+r4+7ux
RYTIWV9DCu82/7CUBtw45qxOLGJS+DRh9FNfqy3DH0R8LDDj3btVIeLkxTO0yPdK0qUYaiD3WvSF
e/zXDlNFTnxxxPW09WDKvbG4Ri/6ydGbVMz3IuD4D4hGe497LRApH2F+5ujBCI3v78RmYl2hEdXl
kMRJ0ZrDIWb7GgKCNsq34OofqDu9V+OBhTbiJEFBHmV244tPNA07nUFb41oa1toDsBT0rjnEwYt2
FYkb3AydBmL8es5rp5cR4QdGLCkMxTVGBa86Q1/nPPbd61cN78Oge+3MvKzaVWxf9qYaXNjpJGaq
jSafzoGkxQlxLXZQO31V8+y+I4JfCsclnJqviuLOtdxdX6tIoq9nhkPxOvl7mGBhOP4YPjAl9zUj
W2hDkM22sJ3qMZ6MSQ11/hmwgb6X3dF69zoPvZL32L2x15kbq3pcdgJ0vPQrEdfLIBuVXJYkqhmb
jrBq91WU+FstDVC7oaF2hZPVtsAvgOsvkfzXhDt3SIaAGK7qjTyk5z9k5awxkdwvXmMYG8DaEZUs
qzc3HtSRmbIdOIBKhZaFdlK762xoOINh/Hb2znbFMniLq5USNF+QvioundblTdEB1KKvg+ixxVJQ
bLL/ZuVeCudgr3W310LtCa104fgvOEAo4pGlLG4ekBj0zEIpuUlpQb6W/ZptHOepemODWml/teco
DGikOBkSLkvZJqnWteEjNb5z4Ml4BtO+JTub3aj8j33d0aA37q+BzyRskXfyxpPjzXQ+CnZWcLec
KKOzP6AIsvJijwHBqmpv3leKsUS9KtZMxH9tTzZQblf5NJExayP82Msn1UrhNw/AGmgy63lF1PMZ
xQO8ADPXPFnyCASAqwn97mzOWmlx813jbAqNicBJ9q6qRkkw2AddWSQrWqDt0N+ez7TJ8bzC+ZHD
UuAgF0IrNug6HI2s6nPjYamfwF/PkhhFkWaWQtLTl8t5YrMe3qJUqlH17Q5qk3PFMQdsA8us59Ci
5Bo8jqK+3HvKnPno4cKEvtJAlngpCPVnqfrKQf0D2bOJNJHW+OZEW59MfDuTDUakLQKC7YMnDG1n
SMQLwDNgVxqTTbVnPkMmCBRV5hkmXh1oh7pZ7ecP9B7UQeoBwfpMVWVyzFPk/pjz/KVIEmjXZFhE
I5qzFVUZZ4ThxUe/deQib5itEXverkbrDElWDLVhnO9QhtF2dm5CHLoi1OZaJAWn5zgyh112XMyT
O22sHO2UxQ0ST2HlpsXw8O+4z1gKdmT9IF33lmvvKgZi67qj2BAOhsJFKA/wHwqfp2wai7jZ2R8+
iHbTZ14AlDORfihDxUMXV5EFMhKmYJhby07EYv99iFRME4esORzntcMH6okJ+/AwkADXFyVwlf5Y
x1pcLiRQents4Q1xicBjrSn5+pTuqjXH+Pn8k3AcLNIy8YGq+KHoO4LwzR9E7T0VM0QJWqtTxSj6
7Ler9jyVhZFAMSUGmN8VTNvui0cafo7it9d1iPteEIibCiboFTUheTRIdxRffme7G+9TlYT62xD1
6fMO9u3qBdE+itSdbwPrS8wQwo6wLpx/In5j1y50og4c9kZAs7eUg88jUObCrUFSktZWYym5p7c7
w6I6hjreOCi25G2iX1olZDm/JmxWdxv1NmuZFnG8levQ/6qwoC5+dH3HN2Teyu4EmdNRFP88sDX1
tr5muM6ORvk5xvYaFjFltPlJL7GOJRKiMimzsU+9giAvx8xQp3hX7fNOHXPOQ2QA00/0be3E1lEF
zRPx3sJYDOmibh7ipEvFaICObFzYhHX82Epq/pPmRC9x2vFYmJiRDcEhvbDNuylBilLlpmDj9iuw
RldeZhppDC7XTpbnkJcFxBuQn39bE5Z25mqJBxC/lIw/PDYwJ2EpQWYTBA+RYfWe9cS5R0bv3bbn
9r5chcqY7RLZuKEUxALZ5h94R6R+WViZ4p1S+KCFokCA622+ftpUoV3YvJD7eO6D3ON1WIojVYQj
tByohYQTZ7ZyeZwTW9A6kt9ftxIu+67Y3EKyHzxtjA7k2sxV6btpbZ+zP4dmxtHqG6gAnmaJw8nH
MBTnSfADv313l+y2zx5NKQWWavli6EYp72xN+P5T7uXNvCS/tO04+NrM7xce+ZeNfGwgbR3+mrev
96fdEDF503COdyoc4QwxPi3sCs8YfZ8kVuupveSFqULlELQAi9Nq0j6FS5nYSavNBOPkoMuSPIOd
0qsW59QhAIEEFMYXRvLxsCb1r73yuRdPDTgsft8ZBPIh3H4lGqVFTUZgN5wk/iulnU9h4wqsxJo4
owjstFOfOQ7reh+Taa4S0NKu0Og7uk9o9oNPkHQCTcEseMoP6ML4wMV9cZZ6mB9Ynnxwrrk8W9/7
45NWpk6Vwtu6usZgzafBGAK9ixv4troXjJd1xXegntUAE8rObQgs8xN8HST+5qq0PbJ6Hdsv7+IU
jstBEjWJcPcLLuPeSRw0jLriSHNshazuqeH4vR+/5URvx3Tz24Nf+ifwP9H6fmQOasnoqsTUDxqW
9prlhkAuSN+BzH8mEKoPHttYSQ1tatDsYbyNvYiEGS7chOVMvZcpMLzW+0KYw5EZFL2qU+YAG5nL
8EdiPokBuuSTTyyXhWB1bEXfDTVMQJYsa/ztgc4AVsyJodigwf6bVtwGUdJTzdi9DHbxjV5VQuAU
hRnvpX9VdwPtlkDATi09WiJUMhyed8yN1nB4wHfpUzl0FLE0rLcoixBojAofiVz4Zm083cW05DnM
2eMvb8h2cd3jr2OBlUpKz+uHjzFTEMCvdpkIBtBU8Axb4Oc3DBM5inNatO26BE2CYEqXdDcacHO3
XwVbI3CcUpDSdFloUY8qC4HzLMP/cxYuyLEOXaGUa38eLYjzNCqaYlBZu5USEH2YUJjK0BgxIhhE
u9wFZzvZQ//oOJZOv0MlmT8Iw1XPCK4ttnGjGE1yAewGuafOyZhfDiIViCm2QcKuDn9ryDfaSPvV
ZHi+bcvKHY/v8SFkKwWIEfLvIDyVKr1e9Hr6J+/2EcBH7d3kmcbZg3yOAA3+WR/mPcwHD0rAh4Nk
P+s5K/5rWxHPOwhTkqW4tCZO5sWaS2preMdOpUP+xCEC7BuQ3zriAAJUcy7xTldi2mtw9RxyRBlG
STBSetRMTralgTTI6aI3TG54A8RUlkyDs5BdhkVL3+qvt8juebv3Nd8pQfOgNJvNnGlywGO/WO+A
9+5xt2FyQ27QJCecUc7OZziSd9UuFEwNDW+g6Ov9Bb/fMczEkwz/WRd04Ja5Xjp8L5oXwZLBNiNO
sAymvbBkxUxHP6vT7kLGXzyfd2+yOyxINIOovyqXozo474PRNfpMLWFybmjugIrcaJ9Ix2OOiRYR
RH1M05SUenTeglWVGAtAuJARwkfapANlbvpiIsOw8mxySC3mbIJLjzgTceG8+LgDZmRUrYtK8biZ
TbpTgJ8sOnAL5Z9Pk6i1hD6P6cZYW7P/CiXofoWGpkDD5O9P4Y4KQgLSicAanHrRUrQ8WgTxvzYe
je2cCx3fh1NrYPu+YJjEpLCGn1Mlh0G9b1BXHVotofeLTV9siX28F914wBjEhJ15qltvy/EJo+wh
pm9B/qlpz9qwHN63JZnHiVx7jRuYan4Df5VPIIfpUqhBXNeOrZzgxah5MA06xfoAuH2alOmlCPmV
WGXsutkWVZyQuKe9O23agSNyy1tcAGxMxkDr/rN/Jmy3rPfdfIyhNQ/2hAgt4W1d+saSRzkr1dPq
cCs/utPhVzIW1hYWK6b+Z2gh+U3rjtK9M+5rh8E4EaAWG9d1g5M/t8X6/e9GWTsjxNgPbUs7xt4r
1Abq1hFAtRYG63KXf8A1hG6N4pW9ItkrASEz9R02C4VR4D286H9U3qzU99pEeL5bj051oyLOpfLW
ldjhl8STPMgUBv4e2iwxR8TvZNr98DkiDar9pGoxZW5T2mEzMQ+H7AWGNI8eSN03zlHugTcLXgJh
p94J/DwJYynSAwzLxNVJsMFLUnIrR1gghWg=
`protect end_protected
