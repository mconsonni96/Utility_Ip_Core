`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
CK1TdxqvkEl5Dwbcp0OHrErlCHVuSbAHH04tmucb62417tSYctEFGwMCqBPsluf2UIexHHJlvdxL
67eQIVVMllhY+pWNpPHd3BcTG9OBc0NLPS/qa0+FewQ82XPoMMGWfM5axwOdlrWx2a3xtZk2cyJ7
Jr/f5yp1K9skWhTaeIrS9t9vImRJBcSF2XHBgTW7a9ju27b+Vw5Fapfr7yDbAii9pxF5dq8taDFP
nGAFurtt5uxNxCqXJ7sDmaefCMLcE/h7gS5A+WeKCu+rKit1npkJZKvpntWKAg72A4c+40S8ZqdT
6CUNC60YaJsn4QRIB6tB1B3rlNl5OG7aO24mpA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="nNDmhE301cvvKPFq74X9Hz8KF2g4gV8GuGTXlxJOZDo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11968)
`protect data_block
SUO6RE3zfGKIOc0v4vcnZolfoAsyKtf21COTKjlOUo15N1nxFIB9w7f1dzRkPWmHZRQh8vE4quQA
uS9I6uq2J6/ofruszWJASvje3zUc5KRj/0Q7C8OEkLiLdH9wzyNb73IgTZLizjfLavLMKiRNsw1u
WKKVWbLuRnTeQ/PBz3c1YTNfPTYY/A1HYL+DrfFNCQ8vVJrTOhxJEIJ2rUupoS7NzELmpp1Wx45E
RDHQqPJdSulocnukqmzwyGzzbJ+LCAWgB0gfwG9KTzgxldRsMIsokhpD3yHfn1ynorzFE4bwEcqm
OBM/MNt4QMXTSxG1BRYJBGLfN61yRx3f4SI5PGAtlniyy5tiR3XEC/29axYzIJ43InbHp+wIr3td
T5muyzEpy8mKL7HYnwsAJ3kOQArmZOnjLFEjld4MJyEY4hyLSGKiHdDKyMlQ615mTGA0FOCxeH7f
iIiv1tz7tzbq2Z/DYO3ScESExlPhVET5r8z3VrEMX+UvrkdH4exh5bFw4cgH+oSFPa6jVqgHzSBP
cfDvZd+5OWi+JGEJKXuDRhTjW40HthqO3LQBIl4SbNxuCBIGl/sHtl+dpk0rBJJJt7ymdsgb+6Kg
uw+hi7Bk9swJct9CafIiKE9ViAQUMLKLW5EhZAhshjE46bIHPEh4tq6m1xp9VY4CDm+DTP7rYG4G
ZuZQB/orf+S9Gpdv0KzqNSfds0WaV/qxRq60qB6ITE5Cc6veNChKNg9OC5GujL3/j6O/61XgUnBD
mAnib9/6BjqbvRq1QqImhzh7ejRsOHb+RR4U9J0om998aaHIQpMd2F5ygqyQi5/QqsooJIQysx7L
XQy6+V6GxdTuwHGOGXWXul9+IKsd5Y3mkEXi3/vrM2l6sKNy9We2a7ZblCZujihlTl/QZa9qGIOh
WJlBRsYhZijsOMsbpfsQBEBcOzEn1LBWRhuwk7qSkmnQ2tZM9ufKm5ixptTz+uJ8nV//L1m6IhIp
bQC9obFxsqbc0MrcJtOf6AcQagb3qQCOinNzne4xVIP9GsppjPFeVfKSn6VKUQ5PUEgnUWxhoWkC
IparRQFiDzaP6kt5iguL5eVMaWPYsXJ+CjvrjnmwbVdwjZnKW2ze+RiXPLBw1KyA+1k2gvuqCHaV
rahRmjqfmQB+MaG8pUgbCp3357UMF8h633h2Z+jebt5/MVjFfsXFIjOheY3MoxbpNNgiSHIlNJe8
Da79SRLHgzvr14PXY8kBauoazTXXM7Dwr7P8kuutZvSdKtFWxGX3Jj6sYEwAfBrTeFIY+6vRMhDL
R01w8v3JENGDHDsiR7EM6xDsks6tzL3vgF3/R4TtZ7Sy68q/rkcmBDkTJ/KXpkwMlriowUkJoTOC
Orflweus1m/jJuybRLa3P2B0FW49b/znE9yLDKkUCeP1pMNjtQqBNRCHh+hsya8NhiCDVAKdruzi
yroCkgvaXfznLPoSRnblAH7KZtRfIEXK7MrtN1EmYOKAMU8UJk2K4hkYcqIRKp4+ZWkSEixfiNEX
Jz6jsw6Jne80V+Ce7p0CAml9aUr4oAr8O494ZZevJ/ks5yjTiHfA8h3+NB55ISOqB7cntw4duU5w
NQIVEuuVgjsWb3y/1IVnVCubSSfSV0kO02u+Yb3amvMcuZDaQQ8AHW8TeMpsImddFHESxsGfuPp8
hez07MVpAbrrX4fGDss1Aujk+k+h5SFnqHxlTytKDLcr4fVbe1AJxRRsySlfOjd9NhM2rGq471+O
LGzbZMxE5bq6cWp7JUlfKUEeJKIDHZvD/UKsQn7d0pU0sJhDE1wDhLz5tP+c70r5XPvc+HmsOPoL
Gv+5Koek55+lVki9DI5m2wNiDxH/QWzZfsZUaO89C6IpQfR8t5oflKINso07B0OjRqe34DHw+zlH
g36orRIf4r6AlTNy1saZlui1gcA22ZSIJP2sijnUyQxIq++9mOWCNHITyduiO5WSA7bya3gYLudQ
rmDYuhSswxbUbQ3V+Hl2oOJS5AJZpPwv8Cz5WuGmL7Qvi+CKSx9i5KsVFrZgZKksuVGzGJI8DXup
lmZIT7gItJ2GRCAVGEcWBBvSlrJie+jyvc1gdpmqJUbAabFsZVNmhHoQud/pC2Q4TwNXsc2zgwiF
T71DaL5Ew+2iwaqjEi4FLU/WmXgUI0Sm9buUMFiAj50tetoSOrCk9vD4ltfnLHJAZbk/oThNqi5g
FrNB98A/iDCySHKIq++fWgpInExd+InJOANa2SxLRfKBKSUF3xTi5pbD/uIA2jlB2TtbII9CR52F
0OAY5mhkEedHMn7wZ9nMWiaGJAu6JKVphMkvMjVgKoD4n/Ps83SVfJ3F7ODOowEI3kEJ+10R36sS
H5GdSFlUu8xlKL2h+0KjLURAFIWHs3gXIDFFzqFqjjbjWSuZcoJTTdeGxCPkYDhEUyksGgGVT21h
UrRBJcpCrlRKd2808Eu97sQl3KKpjuZxuPr3za8Oz/RP+NGI56qsFGax4uClfrJIiwbkkhjJEzYd
1xxGuv31/LAoBmOATv+5n0D0eupZNJW9ZZTcGAA8hy2DlcHKIVaVO/WEYBW/I0GqKCUIg3Uotv1h
2bmyC7z7jtQ6mb3vlteeIJubxO1Rg9LPfjqXTDuNUZeImVPSFSFewU1sAU30tKlWMHrNpu76wC6x
rXVA6+OPJE7tV+Bz+0h5oArA0q92qUMhLybfvSdC05zygFmae489lY5N3yA7QG4+DE61zajK537U
ecvVST6Rub5ttPxImYmJHUCCTM7oodjNnKSVIZBBCbqbWubtc5kFWkNl1S4uUoO0OMKgS/EBg6wN
jIOvJngNNq6OpzCrrsoKgqsoN7D+QW5qgfVzmg7bmC322DVI6uUb8vORI+vjXJeAKCYFM7/vtygt
bFTRK1y5Y9hA4O4rKnDZyBYko7vyqIhZjDySftk3lfVaq/XHiH036Mlup9NMQZvJWYQVNdtR2xOZ
OgdEhSzwPMlPFF3X9zWjoMPlrk5o+ewu/ZbkX4yWyZHER2P1PHtuQkO1pt3XQtz0n4lz+2+di97u
AEzc+vv0kwgRlm9ONMJ8NDJGBa0ALriiJNqwvjF2rxzbcy/RobcuttQsbEYW59IcE/edhFa+/uEq
1jEFNfTNwiiZ8shYsBSlEYi+1GEzC0n81BxHueP633rHXhcF0INqrBn8lUSafML1UK3B7OxCF9No
YLHF8XaTyJ9hYDlsqPd9jy2PtOlmkWcdUzvzWieCEae7psq8UHZS+L2IvBHb6NVf0DFrvWsRZ9Ju
dY9iJV1o1K98Obnn9uNLN0lu7/aDKUUE3wF9w7RWwDxEj+pQZLPzP7hsww7+56APFKwHTA3ZKyLf
JFhUPd+vevxmDr1mMKbQzZGOB0sFt/xcK0dzkDBLiIgFCTp96ztGNj+dJaf/2qFDlDoDBS3H0j3S
uW7yLuZ/cmQYcy7b1eh6Bap/xIuCZGYLMRI28ZuBDMa1emFMgBle4MdD2rTSGuK+ocG2hoHMFhdz
d6MhgXQ1S2pQtIi+9cTQdX5nl4XBWR9543OGB04y0SSMJkV4OwInbxm2tuPgSr8XSvGr+/WbIF0N
ySyrRTa7WIJd8KWeEeTRG6bTuX5yu358Kjbnd1mHIZenCgbC74D5Ky+OwZiziKkXvMJgDbCmJEZL
cGLVBbksSQgDPhlcKelRo4pJWeyms5PgLQv9cCa1K8JEziTQ+/jngAKLXxfHXphAzwfGTRM5WU+F
+jZNC5R/SS3qiVK6tV5SF3cwZSLCQwysVWxh8+dhlbz0NtREbrQOsMfYPCmtKQnEx45YAa2fK+I5
O2HKie0mW8aXKFVVR9KngDH/OBDFIP3D3vmZTMEM2uI3KCtxguQ330oECSF9M55tDq7c5Kh5Qd9+
17hBv2hA2hEuVZtRG2d7tD/bu8yoiXoMg3JFI3ryksT45kx7UBldpdFaOV6PGUt5l35IjD9UDAGl
aR5v4sFkVUVVvmjJrJj05NNHTx3nihiJ7T7lBedmp4tRg6OC5m+5ZG+AHytOT8sIrLzEnAYDAOLj
USUNPhdLwcnIlG2wyGhSogeLRDWtZ2IQ0hW7/txbdF1s7z01yEKgU39o5Pl2laonnCzb6brIgqSx
iestMGoWdnCIybpgh5Rul+xcAgtdz/+7WE+il/6RJ+h7KlWpep7x8gGKl6cfC0L28ntle0ilQXlP
NptrFHdI+iOfx3TIQffJrW979YMPw8OxObJJY87OrE4rq9a9HA9imuSNzk55dJdaeS7tbpO8Z8p1
dYGzwia8HRNUln4SDA3WvRcSmv2PljTTdJTMswzoP575oChOH7yZ7MsdXQoN7brR1SgayjnvPv0B
xoMW0TtOyiyiAcNXIMsW4XhZtZx+HLDP8PnBUD3yToSNclf+i/WHWo2jIATohESPjp9Cj4numz3V
CSfRS5jXaidDbKe4By/N8a/AXY+budFYQgKlijEVsdCEWtb7QLHYdxrSnVukbDlhE+bOio1wo0g9
cEWPpfBJ74PtIhZeRjITZsK0b7c3AYIpYtDnmaBrovJG1lCbVjYu0nh/DOGONeet6S9hxh1gl6Vt
ZJVzVShD0osGCA3HEpKcydXx1TQn0xrTqP59JgXX5FkI67gvcY9vai+1KyW5E8WfcSDza0FBwdfK
WByX0PsNRa7AfbZIxUNwroR/Yh8aQb5PL1LzZxdQtECVxqdTdZcjTjnITD/MVezsNAMBFTJPte0f
NnzKvXtSBZah4x1IZoendiuoXVKDdQAPkcaSe5piD0E3M2TuwnMglgf0j+/J3sQv7x3EwfcdGAEv
6cS5btZp9xameewYkOVHm5t7rv7z00iJk06kPd2op2lY7NQsCH6tsJe91CuGv94fWnMxzSo5Nn/L
ELUO8r5fUheFu0owRq3j7BbtpoFIll37nyr+JA1ohrcqHdAIeXRAV3Qp2KcKJpac8TwookydVh6Z
7ZMjabAEnGaAaXq4C/ghxNEi4g9LEMbv4yRJ7sbiOZj+waYS8GV46dzo7IrUIrAslx5qFvXMdIcZ
rHP0jb5r0PiqjTExHBmfUDRoHRkH5eFtec1OFuKZZ2Jh0QeauLmYYfr+2MoqR1MJDWjsbiRsE06r
HRHM9yS5eRBVLXbuGcpQvrNP4KFlkizRm4lznLo3tkKGbSNUds9WIgyxEYwSfq8WDEZonO6Wfsjo
37J/sID2rAZ+7g6o05mG/aCwzWR7In/hafZaaO1jBLgxRY/BWsdl+ZyyPdRywzIMuz4znfgOEudS
L9AhtWOtuv4amwAr6rCjQps7qwRjGcRHN3VZieXihirfM5DyN/BXfW4YMM9O8bSWk3KO21Q+H1vh
KnD98xjj0zYqB5a4iffqxue4pCl8XaveBUoNCu7x6UhKwnfnj8J/fu1eOr86y02D6lEp3dFv5xNc
r29KBeIj0SH46cuZ357Qo34klXoO4Jqpam5UQ7MBKEcfpTI1VKif0hilQKA4mV02jdP/hyNpWT5o
cP/rF9NoPioA94hPYGOXM/+cYqiFRInWO6TV/zrI7VCRX6gH6XbmHdNvREZucSL3jXYzL5hy0gub
XpFLp0UJj1Smn/9ZFjgvqtcq0h6ND3p0QNvC+36HJi/1ZmB/0KkXEYrTQipt7O6nQL7cWO/yldMm
BpxOXljB2hS9G6kZAT8U/89muaGUwhjmdqVHrpMkPAPX6heralHp5xaHTZ8cXwBt5XrfMQkw5tzM
ZVZ6JC5dOdLoDj+bP7lwjjx1DNK8bl0GKwtME6AtOwChGPAXJkaiqK59bvQZHPkN9KliKF33BGbY
U9Kwz63efPInMJRXj56Yd7Bvdd3O1Xz3KkMvFxz0F0mHjc11qHV1bk3sWr0Lt6yzNLXX5cS/QPBS
C9PGC0RHVHFCfte9l52cfP4nXUBud0+bxACdB+J/JevT9OezrSDBgVW9Whz/sQuakR8tMytyCig3
4f1ynyWeWfS1F/UxQ5lk4c0GgPU89dT5nAVgRDE19jFYzvd/t0GDylaXY2DFmPg/QlFGrElPBgFI
iL3jusBu7+ndj03hL5We6CtX1t0YBL2Qr0y2qB8gOVu0Jj9MV1ViINCI1KL9uRoSjtF6/BXp+PQd
jNFnpBp9V19LCoRUzKgx7Yb37EtujSYLcLgayAq7EY/I8XW8InN2J0JnvShavGH+bvsd4QEYFeKc
WXQSWc65mA0Zk3rrBhRHY2rijiWgzJxpM50hRu+qkgpTK8ZV1sYRxLgvBax91XGqC4o3IBRchebZ
3/ByczWhpWuVheraw1V5SWwMIlVmcEYQIk7eFUr7J12dJ758+aygDmWeZsezNAddxh1ssy0NRfFw
d8p3PWo58VBwGUfoRKTblpWrzura9UkawRS/CNHHBHJr8Dcnm4xtiw2lHDphaNuUl7+8zGk0M+yX
qh0CGGCyddcI+d8QUNLUDtPvN1XfE0sMsGIDKi1rABe3HzyVDn+PxtoMhZuYauTZMpzGBC92lGtR
JXnsthehk3UFlKiIxUB3Hro7nNaRVS5NrKUMq8Fh2cvnGTYgLPBOio5e0PtjJpEn+ZvCQD799QzP
cCQtlsXnXcA4PR/obf3+L3NUHX07kO+2O+ERJ5gxVg9RGGD77Jffzfxwybm7GbVptsusia9s2aE8
YsJu+ybQJGi3OgeU6I1Pyty07BspVTebhbDj0ndFVO/AuvTEh7Oj2JbBRhPEcp27NnAMvomVQ9La
bXTUglQip2BsMR6jxtIQnYRIOSuHBh3bdsjUaOzfTfzZveo7ZlYYl6A1IvdJgxgSncEeVBWORc4Q
oo8wJQFeWG2jbmDnO7NKtobzyCMHRbwloO2OYGJz1DtZsxpR+nZaJPSC5fqiqyOR8x9ETc6pBUxx
qO6fPqH/0Pdiq6yE5cwtocgD3s+L7wRAOFvqA8Wk9YrtLCh7hkduUAW7oScSarPC7/K98Ql5ne6G
qh8C1j/6PADINVqDag3jmX3Iu09MVy5rDIlK1w91v9PRPmXPfvkB+56crz/YjM8vlOQ+QQRR3oLw
PPeF0lONeK8IoKrb3qUYJrPxNRYC9akXl4yL3qWMpL2OLTnqd03t8z7d8MX7LW4sqicXKx7UQMy+
J2kkIG2zF8H+ZWH08qVkXU5LHVz10A6DANHQVihUBUoXznyFO+QSWUwe3qyNLth9RgenbN1wfLqs
VDQOeSZXO0PgJ6L0HzMrI/IwJAhRvSzdTiFrna9i59YnLxcYyDFXf6PaNQgXsuj2MXb0ODOPwarG
HVeX1Mrbzah6zZwaDoauQtk9cYOwcgH/jaN+l4z8G6dunTW1+Pi2Z0rQOHkBmZzY14CZb48kd5zn
9/Xy8KuDQiKYuO5Yp8clidvwiyAm8HdGmesGvvP4K4R5NvEe4VZROzeJV3XPoxpy+LQHipBlZ64r
kGcD6dihV1EF6Vh0EXBPyezyGiD7RgNmPXj1PZtyfbslIakf+7B8Lzun+HYBmEioDz0+qWAa/Mv3
RhXCbE69Rlu+9yPw2O6CvwJ10HtVXnfeM/Xh99ZBNGSDiSIWBxzxiUTzxPKKCyZ4mMKGHkbw7KiI
7Io1TM0hVFK6/B1v2glalHrTI9Ydvz7MNW290g6iP/P5IJnIT4S1k/djHxWXUzPTaVzeRmyu5Vje
1i7v4x3kdLrNnigx+RltwTAnv8B/CYrc5zT142sZR0aSVtAoajrJeavez8Dp0rc7w28iJbNxptDA
8K0irf19fU1WOqAcB336hiL3ndEsFyYfUEP5EEByw9wXxdWolgWNbDHedhS1bVIfxKxTdCSDWKFb
VH5liS4MxwfuFLBeg0xFkOmIddf5SwJTpcVq/WwjndE7Xk+gIApn5CzuYqvLLAgFCoptwHb9v9xs
vdt8sWJ3hKXPzXsbM03Emytam3mkOAkxDYOhv0me8sSXfznh9CtbWVpvkSGaKgn/3J3KyKeZlmye
19BCs0MQtrbOHAZFbwOykGK8lWWrBJZq2AeYT/WnUpYdARn6X+Njj2RcRYqMJcc6wONUJLdnjmE2
7KWe56TxTATHypdGoSDQw+hae0gZTN7dEwFad/WqJExx5EMeGJBVUnB0GmZpAXLI8F/qRP+KQTNf
1eRkdytD8AANcxpBbLXQmRI1EGmHEn7xmL7FitGRBM90svB0rdH8k6jdxEZujJoh8a9xj3Pq4RNi
3vTDIZSVIhsLLVjM+FawOdMwNiWQbmeKxFxRFk3RckusLJlYscF5W8M0HwYLYLymNMj4Uld9bK4Y
1zZKRj9QOq/g7TDqX4GlwyYVRy4PnwinsVl1sjcg9PB5RQnoICmyydwdLPIShphbcE0Ede+qEe7Y
Rf+QG0GW2GhGs1l1PhzzzPVbIWQm7nXdy6hVDb5qKbdvGASx9UaGx1VZPoIJRsWvDuEZzXODr4rh
UfZX5blH2NiyICUV7MllM+3nAaPjpy6wSLpmWH3crRVShhjjDUhJw9HzlVqoqTUBohGclHHixA5l
ra1PrG56MG1vnb8Z4jzcKuyBGg5nWa1VWnMkkkpYCjYzUSUJKPoCMp8KvMP4CJc0GfPzQRc1OC8w
ewlQ/KvcSUQySYuChHRXHehlVf9WWclIfbTPwVEAKTcMEk47LVl7xcdMF5AUlfTiUxiz1Nu/zGIB
86UVj6Gud0GIQWRZOY+VYjomsiqZQUzf16KceByC5ILsBU9iRxwFxXUtjDAmamJUbCPzp4bh0+6y
D74rDIpcyPDnVt+im3QZxq5Uvv3m/O6UTBaD6Y+lNrMfckM2LIc0kqkgHclXmJcy/DtFdSwDh9K2
koHiik7Ql0oZ+T9jogLoWGD8hRVzI5Pb23QbcVDgK7zsm69MzqSFumgwFvtrS2LMYHLdttX1XQJg
GF2REQK9SDH/8lXxNCvQ5KXv74oXbvBImyRjI2ymXseFSs6L2V+3XcO+aQ3zQm9EL3L5lNhTfVr0
j8hQ6e4bv/3px5XahEoh/mxohTMBMdXPgfKlRrRgz1Xq2DQ8tGTQdLwOJZYhW4cMkltcIC+54AuM
t2nOW3NBzrPQs4txZGZ+SkosOnyDIt+W3zNHJCWZBhE63iFar4CSzy1TnTsAz1tn1GYXlIuIDxko
s/MgzoID3qEmhWj/k7zAWi6ilDTKtFPRWPkzM6DldBVO2udQhEApCcCMqD628Oo3l34eGkNsWwhr
rKhjxRlYtV4h1I6fqMjejTQg60urNCkxfVky+12WdTDQHbkIuzXwySOkyBI1ae0M31fF79H28c/+
1hyVLFs31X0XK7Agkpm7108tKalktDFTTnMZ30SttiM+wylWwtpLV2b1ub+TyGvpzeEU4tO3Siq+
1uSgGfqX3dib1HqyTcwCk/bW4ScflwARlntLUkiqZDzes5rKCCkPPiOQEI2ktP7arXYpZl4Y/6c/
aUvMj1Dd0Ky95XGvOnF1/6PXxfPoQbo2ETTdImY19H7g/DTfxm7pWu/CdrXgiks6rncBDpgoFVhv
m2X/UTv0ShUpfu1heKgxovao5sDDTrGNK5WqVtqM02JHId0lqqcyjb9dLtzPgO/AN1wO6rEpaWBc
g67N2SXq4OUjN3Lv5UuAai/PA/5IPD0tknGGN27qBLWh8N2nK6UbqHSh8vsm3tQnhmCLt6ruz1xs
QoC8oj53csfTeQMplHeelnuZU4RWNXKq7kLpBmawFhCFjHY16t5fQaS+HCThlX0Q5nPEM9S7hSp5
FMs+qRuW9Zo+Q6QDLWij0Tw7Ol80iQIYHn2NxzGApXe7l7Zo5/IEVWV7KI5W38j4HuG7levR878P
q3miNVcF5ixqn1PGe7ZHdEzKOzQpKM06j1+7ryzNnHwsUyILMOF7ocKuuURwx006omuw8ytvFjAz
llDlD9GnAVJRD9t0v+WiRVdSmLnlTGUslZYGP4uZ1rdezeaTyMKbIJRXrSnljOE77SSjlz4Pb5Pg
x9N649LRnQ6gftLnobHdfmVGRcVQuytNtqSn/yh13dO8L3ULAaCNvyH3IklKRPd3adjcw1iuYlpW
K6PHp1PL9+unVBMBdUZH6Axx0WFmPbz9//jTFwK8B1dEBSnY0YrNLrxlOTPFX3ltP3dCg6xtAPdC
4CLjJY9Q8Ob9Mp9KYoWjbM6qR+BuTRswKx/x8RAyeUPPlCVd+07U+ZUWIF+lQY3aqf2nOJDukbVm
QEOcwWhgMtCg+02aXvNbbCTYqhePOEn+TEwhElgVKc8e/6JLtMSRQAQzl5t7N3nBSfXLijj9ymhY
/zpGK/BNoxLnAuwB6L6UknYWbouzoB7RWXsfFb1vocFi36NWnEIh6IAC19Ymkmxti05g4rgP0e2w
m+8pdjL7kcLqwthJL1jxst0stN2e5wN8/MlB2AYt/mDAwrMN/yiyQOp5qHZsT6Euk9oU6pdWXHaU
hMnu8OO415Kma1TBpprt6DXQOsBiBCRfUY4pgUdooh3gITSwcI5hLpI+CyofpcfUODOXiwWzvOu3
rTOyI5pu+5hdkP8Mn69PbAKphnAfbyUZBZ8fM6l9BX5jn0IIYJ3DzeR4iu0st/r3ZUl0fMy8IQkU
d2fM46XunORnbm6tynbVsCyE682H+6fZWJqpqGgUuHtAMbVyJ1pcS9BJbh9ARY4zNOVh192pEcHf
viLxKGphMrkjhn+SqBRd5W9OHAmapSmVUFOpkJkjN+rZPrOxvnif60tL1OTYypnYY4AvoKlB8tyP
C8cs6cJXROXET4y5hg3SKAaDkYXwslTFZy93AaIt+Xq9CyDR4u63+iaeCWEkgyW3SI4nq+sv97A/
AMBumBbd/IzEkaC9ZJGPKBE1SqCsD3n7ihVPQSrMk7We24fAIOMbGm5xyNrsvebdn70nCwlphlTH
+BnfPootM5AeYQ/fmTavC7eFtGe414yIdkmKeMLNWH5OI2eLV5mDPabg8oqV3DqBy6PWi9S4Jajf
IQKQeC482BPqDgATM0jiGnOdbjOrG9FeM3YCpb3n2aH7tTDY8jzn+Ds+IttdQsSoRYrDQ/7srTgp
o731uWii05ly6B5H7NywlZ6VQHT6yT5qiX5BQOqoTH+eZqnL8gDKLxmvbn1oFDhMKFWG8ABsOK6u
lSpO5JY7LVKMlTws5Or3vDzq4/pwMNwM1rYLnD26k+TEDPUN618jLmZlvh0RPcdv5OYwlI7t4qU3
BCO8e/cA8sxJZ6ng6T/zyqYgJkyOLQBcpHimbG7KVnyGRygT/e/TSFel7zsGpfikBaIo4FXD0uDR
5PWt6V54o3tiGS3Pf4v8L2uqRoXgWVsE3B0eAs7D5rTBNO86AkucMAmWZ9/pchb3/BhVRlcn7Eh3
NOZRCDYOp7vJFcDiKqh96wAADsp8Rej3r95ZqnIhIGDAgITztMzDh/DiXIJaunRy0zaWWoV9aNmc
5whDTXHjeg5rwfc6V7F1RVyLeITTiIWj0Lpd9awf+Xl2hsrjnxRDUgn1iNaq2fqAqASzzcKJwhnU
IaR6XCKRIlqKIuUJmEhW5S+34WpVautzs/bC8GIzmnPHwWo/izvG94LqqV5L0B7F/RbtJmdrXYud
iK6SXGngIVGh611cMrx3we4B2FbvfWl7+fwTF5f9LZFWwfE08u9BVWo71L8izIrhOl3ko9NS1If8
8KBjq+EOrqME5Jagd2Is89FUdawJwsjP/v3XDwQCoFUKw9VVzo2y3P3jMXUT5PraQK0pZqOZOu4w
fRjSr2AG4DAj3HUslsumjHNyXUzm7gq0QOBL+NDj/p2x6XKS2ojjh+pXbD+1kuoH3/VE8bqCwyNr
KzwD4cYPmdSKcIHs1pU4/197qx1fItVvwFvjWYmNUB8esbX6IAjXsNTnEpfnGpfLmpDasIgtBvOu
uL8SnujMsdg8sY57Bqz2cx6Uvui9nvtzepG4AWIwcPprvmsnnadyG/WlG7fNn+c+puXTmzoavHCb
1n0kjw0yiiNVoXBb4FDsEqFLQaXNt6SIXpqxgiGfRwiyKVZsvptDhIJhk7s9/hinAtfUBmiyvYwC
Tpv1ioygDSGnZ1tCFhPwgkFAfMIbxp1A2ZNVnz8W2cTSzBkRzcvdUeT4vCVJjSMzyMXZZEcYhfz/
douIFLEUxVX5r9VrCv9Y3eWTpVndr0qYA2ScxcXNZtY6TCFRYFziH8LtenPvRGxf9BbMp1wqoD5d
0AbZgYyWC3nSsWHUS93bJmZqi6Vdm+QUOl/gye+aBkPT3aJQusm4x66a5m+t+wHN+9DTbEUtnpAq
rfl15QKn86gBkY8HxgY34TUj2oOb0l3umrDD9NqdmK3SufVBQDEoLRqXi0rpa4mC69xuaxCFNhpl
PHskO7/eP5KdU2fop0kzpiAoAWxIKEV6FOGh9WgpbjJ6V6Wr3iEVAtcHUr04oHAKyuXjepdVJUnp
NtKR1GbuPz4N5/JGzmITFphIF2AOV5vY9MZtgHQsqcv0lV0hjguN21J0a2RtLxl9ucwP7cPKAyZj
ms08K6cnmly0qeEwV6b14DhaFGMulQYemPWZaeLU8eqXF5Z0qEimRSNixx7IW/VnS+sj6QUIvX6a
LLAqwd874w4+id+4owCMo9zoc27Ti3q45toP55bp1Rju9A24l1A1X4H1pPPLoW4XD/4E6iU5/4So
BCyYRYxTbI9zSb1UmljDPOoErsjwcMp4VbASQLRg/8ddJmg7qxpCZ5aDWjZ7GT1keZ/pZSzwhfUN
2eb1h7Be2esKqFe+j3zi7lHAMtlMe51sFKfAyB4ZiVdN0kKHUQmjfrk/cLTTC9wGWCuRkbZfKiDU
BduJTUmt7DYSKfM2sVQZLrCeQsyqGufdvZeQcAZg0IhSzHetdMBSVXlsTfUO2zPBj8PBGq7I0sfN
WGZs6j813pqh3Zs+6lNFFhZPuKQkmGWxUKTS75BYbSiLU/H1//GEzLuwsj93RdrtHwqOKvWjPtVk
n6W/0vb9pwCdafTdyxq3hA9Mdgjwxa5CR/2ItDmOmmB8VYQMQSlLgr49fjPdIFZFXM9Zbvdtmo+l
vCh+hSyIhd/e5/lbvIhqJFuN8mIhjYvFuCi3l3NAe7wix4QC9DYoa26TUDViSM0jWna1gWI8SXZI
eawiezFPUuuTLGs/ti70R40+TRyTN91YbDaDJ/1UgaKEAGzzahidS+bvd+Ns8UhX4a5lwISnD2TV
wNfgSu8IYJqLyey4oTRj0TKH+sgcaKHQ/yQhBwdVOzH6uKQULMc32gSVIeZ/+WY2FXkWeq/vHYdF
LxX5jwU4aq0IXWkIeEXG5pSjB7PzTrrteZyqrOD66XlIVPFQlkmUIHY9pRQlrI0LVTCSAM2sSw+w
SzrbxjViFf/qv8ECEXV32SB7MFZsugVv9xMwmpA6nn21G0R82RMNS2BzyyqJrOlwm5sIz09PQS7N
Kko729ZCtn5wFNft+93S4JNRsRgE+YBR89o+mDdgq2jknfSOaK1+mu2oobiIX7p1vNw5BGdDiJ0O
3SB0O9vDTySjjfKbTJB6TzOv26bCyNQhhKnpclwURauYUhn6o3AplJJLisIWHuX7Zw1EppC3eRJs
uzkuCKFYuSy0GyXXbthXncYABpkto706d5t+1UhU1SVO3yhIlGhirlb1jahpEofKCs25p68BnWAZ
EQUG2ls36ACoZMGJUQRRX98jtPh6X3oA3XYuwShPsQ2PgqvEFhfzIx2/HHRFZhnRxps13XFEAEu+
z9xa+avEOeZ3Z62BAUkiE/MeJoSpTMrrDbtBJIWd4g/oHblnFjDIHsjkjOETxLHOlO5kEVWbaKJC
qCMGmY5PQnngqLx12tGIgZ4LinR1Fdt6AWk9ApmTArbKr/FFrftTV2PS9YTj9Yngkw0AdkA69MHe
y81TNQzX7nWJr27ECQuvW7c1Yo9tIUGjJ93FV3lgdG1hRHLT2nHijBPL0OdMx2psbX+cecgYIlXR
8oCNMgyJDrshxyvM2mfyktGXg6zCRV8mk/pgM1aL23drghyieIXv/BwHhTGMVDvwWbOcuTsVSMEx
DwS+ESbfYhnOkqAIWQrKa8rUZu0Ium+4FPguLCcZGI6olL219Q8skIrolYmjk8F3ydLDf1u13T70
jxUVzen4c+fUmAqdghccWjbEFjXebnBXCfwuEW3MMkLfpIqAiWoPasJaZDSdkFc5vH01vpjDK7Xa
tHBzBj3QyzRjg9lbqebkSgPQYPryTt++GZq34O7EuxmZQmUEJAt7/9Hf7iVY5Ew70T2ZZwgbMEZp
3i664ZhlQPIA02wv9S/646vRScVDSin3h+0T/VWO4o9tv0AynCeYixd7/Ns/dfMvDaPSaz9ry+Jh
6jp0Xu0TSxKF6UmbcFozcUhuOtt6J3qQlcvCMgRbUeg1WG5h+lBKNWshFVrrA1rV/45Ie4kB3dR5
3kIM3xnryPlcvsRH55vUBQb8qypCpNWHsO32R5ueYgd2u5wYmOAbDu8exh6Nhxp9bWawRfcKC/64
d+siy4/sUkedmuwvmTMCTrow/x+lu1GkG4S3U0zmIdKBpr9uoEFQ2lnx9JcJO76BDpxf6/5tb3Wj
jerNMyNIRTB1NbjkRC8Mp68QaM24l25iVftlPD9s6AvHhB5DhtTzNCa54xRt83darvkvoZbZWuMJ
Xplibi+9Pa1gZf/SrGA8A9xf7fDS275A8P59NsbHkhBxMARZJVcoblZEaI/3kE49hG166H6GWXdq
Q3RWp1kpItcb3YaTCemd7y7gy/Dv9weaHpAYw4IMXUnkLceQS6awvmZOVaZEO1szKzJpr4LopOXl
EaHaelQcGsu2nAJsa4LCileUvN9wUVkoyvWB5B7FbMK4FZlXSKVi41jMtkjjSYssaOndkjaq80Zd
mNZ48Kn/0ojhBtDU+C3e7BRBr+H8sz/T6+tLTwLdlBcsoyffNqKy++/R7fpnk7Z79opujF2Xshg7
43VLMArMleI5NRBli4UDrc8PJbh1bQFDI6MfyRswHZ1tXY4MGNnWtdC1zkiZ7hp7Q3IO1Kh13m9u
M9oYMR+VdH/095AaFtWZsuf13n8Z1KzaVgAWcy0BtNO3pFnAQn458U9OqL8+cm2q3eN/GdPOdoqu
/vrzPYswb+YndK2jv2jl0vNUgJtaazNKqW/Qess51+Z1nxgDo0ez7GPnhl8vYL+cNeTBVV/cIV/Y
6/Ev+pa+xbWnUWAo/y1G+A77Gec+szibrcQTVEg/YqN2uXouSFemSZ1DlV113BC7mEg3bvhx6rQq
CJkQ8P1Lci5BBmRu0pCj4cREslnNWZwycuDNLkO5A1lkAMugQ2k4dn0qkwIegGi6tA85VXFUmDL0
FXNXcf2qWW6/MwmtujfP0+D2MilxBP8r4+Rdf5YpMsMgSmEeQqK9UOLFUvqBqQkcrC7fENJtq1EP
gmbryPr7oz5xgIazYLOWSEIKUoWSgeG9MuPXmhHB9y1GsgOLO5QDJjFVZqZ06vk8JdKj+0Z+SyLt
RjNlpfqsdMLx3pTlKTentMxPUjNHHgqzHo8JCbBrTwRBGsnafdo+eT02S2KxNhGfGmctSdRP95GX
PAX5Wop5jsiR9hxaBfrP7d4RHs7F316JNsOG+Pu2jrGavTqRavHFbakf2aBU3Mf0LXwGuVBePPt2
9TBbtnf4rYLsT/DsPu5iTVy+J8NCmrV0kB81Jw8x0325zHVBXCa1we+QtCI1Ff2Yd2iXKFE3hPwA
EqTWVet7lCtW3uV6m/VzggTMl9xyaBa7Xuyx5pQJrnrRe2cm91Gj8WC/BB5i76QDaJbw3BZweroh
gFeIWK7O8ZCMZhXhznW3ZlZ3I8j5ria4e6LrDsdHhZlz7sGrgDfrxkSIkVnj9QkcEV6im7ZKdHfC
TDAfAZzIWNSTEOXcBamnik16kKdPYs5DO49VPTMjMOYbksZw89s/aZZiAHLgJOCJGqb3m1azXwJJ
UwofF19wPqFalXFjhZ7+KRYOlxRWYhfzdEUsvMCqRrGopHg+7Kwnj7fzrkZyG8WZOeJrqwaMoOme
0fFrxKfw5fLqfOYOWiNBoLYJkv1YMGiN1XthjfpaxUDAHaw3OySolvCbtlTZw1NII52ZUYhVzg==
`protect end_protected
