`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
rkKiovC4Y1FaNPRRxUtt8UIe250tRkxvPUAYYz4XewVMaXVDIsgXX1ebjTZCjmKlm2Por5n9oqaX
b/8/ZlPzGdh14bQZwJY9li6YJ7yKtYLgy0lteVj1y8Q3QUudpjQcyUUw0LBQnoYkD5G3Iv4aWsGh
G3c7AOeHXQ94joCPE33yOHamGMnUajjyYACEpYFakCQIzNSjrqJDgdaI4VJAteTK5BySwEhIO2dg
VPxGbMIvyKAECKk6wzCQJkOAEDDJI6ITygfHmXObZa8Jp/59MadAmxjyAHDHIptu7K7t+n7SPHdA
owZI0qbePsjhFuXN8pmBU6YjmGdzqU+5B7KoXw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="MCDkgLeN07ofIXBVsEeYsI6dlXesKyHCBQPuskbOFSY="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 73872)
`protect data_block
4XwSeZF6pQWhthNRqP/Kcy87aaOTg2c0OoXsES+uBQMGQJCbEcMfQyWjd2u1MzVeYhddAG5Zb7TH
Ox9lE865x5vt8PHXjQrwwHCuQWy9ko5aSUHGCAr+XGXu6bhfFNVO4J/5NHnPJHEfXYZY/hf6TNWj
UK6CiOI5mA51FCYV+N5w5I/ulVdwuczeQ7OABxSNHG7ElmJwX568cJPv+5famrzlO9zB3xjConG0
kaKY+PJ6eZlJW56/5bKtUKen3RHd2MY65qbHRSfYIsaAzD8Y9KDpwRSKpWxTpjsq+iz7HcL9LPAv
0yDCGvUI8lbDbAyECOgPB+5eqM5QilfKrFzI3fVjyD6QFnnnwBZpLV51H87DFvmQpwahgwhc7j/v
o3V6jstDyLrNvtDefa45/WRYh3rMwYG9sW/Swy/f6A0g7+fB+sEnciVAs5hRnUa/rEzrsXdqy4kK
re1eDmf/urK8+4yQlcVaBcCii8pju4QrOAo65dXSTqNbey4uyl6MMwVTYfboHFQ3l9duRpbah0z7
6pHsqnJyv+zWwjnViq8UT8rEixQ/r94lMc2XvG5SY4l1Ik6M7FPfajq8xcJKUxK44aWPwJ85JCZt
Ud7sEETMNk7nxa8uFa9CpsdtyGkbpCdWsN/RIistxYsaCKB5X8rdzFsYhCPWCCRHZP2vhteQHQaK
qkp+TXomptYlEXbUkHG41RFnb4RK9XZGtxl25twNzFAdiqMiguwaIV4dKZVe3NUYsw0Oj/FfgxCN
bARp8v2LH6FA6IVo10b8tgzyKwOYAwM1IbcN4lvAoa1bsnd2+3V5BbpVS3P6S/IKMGWNiae67iDv
eMFpEhGUoa7vdGih8u+ldXKQyNoF2f4JL7eKfDcqR7msI3jDm4aye4GzE9m33/ELqoYjS4mv8eHk
Ja7rjL07wV1emuXnZ5oom0FQenFhfAr6gxSp3lTEkryD659srN+m/LVch8h/r4YdEPKk7jwosTce
h6mNRxtHdagM+QsSkq0zIYN/kuNNvSaPxOzAOkdXoktdeCl/cnkt1duvuylCtg92HubZx4o6+5WW
6eWGf/DqYEXxCZIRQnC333QfY9Xc1T7FaUtNwC/C0zuieHHxHWGs0ylgTE5XDo9iDNxHbuPZ1psB
HxcAGbzOFSBKvrFeHx86pY5x9omOqrqCVnupJzVjjv75orzMjdGqVnGSbVHZgFocrlceiRXw/eWJ
7DW7cWDYveIJVMabfJ5uJqj+AxybT7ntQm5q2tejaX6mv3wZ6yTOBCWT60j1qGU4sZA/vADgggj9
PIhahhozeFcwaUd/MCbqfenHEUy/RjNnn1j41M6JwFODIHJBl3gYdCmuglBmkhH6VyIuUdmoicAN
/Wbcw5Pnp/qRATye7TbDm6cNzeB6GOjDW0mmWe8YOwTzj7gD3XGckW7qHINs05eCS60DhhmTiHc7
vGA9nJrziYLyK6KskW4udV6bUaeOJldGcN5+2nGBexrx7CtQXsPqbYHPdvVw11cn6bxTvxMtl9gH
X6utdR2KNdidCdQAhs7nd/wDhZNfo5C09cizR4v6CMziOLXBFLD6dIe2JS3bTF6wUgpLXgaKte/z
O0q9ML9W4clghDnFV1Hk63AF4k4ZqoP8P0K4syTbMtHcIeZPowzJ0NUtDHUSL1NVbnvf4cowL0JU
aQaU5GwZZIVIW0pH05f0u1D6Lzl3v+OeQtrN07qofPJvWbc+Urj9VqN9K9FINC0ihv+5S8wbQKLy
QuyLDG3BMuq2k0vR2LoFKD+fX23Dn3q4GCgYAdEFcwqNC4DjWZMCqlBH1HXjndUMpkatZl271Qxj
Ovq+RxLeFQmUIuT6bvDE4mJywM7x1hQCWltmA5XZqIEUUdX1FFh7N50/mlHqnJ/2Ywzh1FUh8mwh
jujv+FkAgF5gOpSFZo6bP7P8bAvcUzEQTGbdDHOj0STbZ8CKSgMikf1+25UHag8ap/JPYESFWaGu
8emhCV8KAdvSFSKoNLhhvtn+veDbszhd6gU4cSCQ6aJKal7N/Oo9uzHwuavLT/cV1tMbWXOhsj9d
bOWuQa8PIxRwr6hw9Ti0UkpqYv1FW1h9t6iWkxpRHYtZO4VWK0hzJ4131dFU6gi/1XBnTBD2lILv
C6nOM6Ew4aaUxTBlDT/zY/meOSlao56nerWA5eb5rCxHB4AMKFX6WBFwVjEI7u/kLhBBWCz2mTkV
Tc5+uJtCUEiX4BgdUw/Ol2UxGeItnQfzLZUXsfAgAoKKIQf5oU4ERVcQbFd+3s7rN33IxmVSdbfF
qa4X4yrTROqdW3Sa6RASy19Qo34LpZPyFc3WIIwlUDKi9TeZQlSMLqNMpzK9sKi9DMHNOFXwFvJa
oeM5FzSo79SRn4GX/bqgnvouSJqBODeuidJ9OED/O0pNSmMpqLSyK5EcN7DEOYGyUtAA60vy7IZA
+rZBR/AHMjAysTt69rSjhveBvyjLRrgrS4q1sjnvs9YTYXjMrA6VDOzQa72MZcUIQTebrg7PlXvn
SR4aL/XZiLEmDzx/qhl9YzKZPkmgQByn6KjIfPRtbZziv+hVjAlnhACRggc3HFLZkHUuRaw3dGvL
Yjwuid8kUpSG3zSR8f2SR0sHxcWvJCfwAqVpHrA2EeSxaJ+feTGgnhDza48dwTM7K6RL9/9PUKt9
aG3I9AtBwJVO9p4z94FnWJIPHXlyNnaVoL0lYg85m2hvhyU6TDpytF24V+V2U3S4ziKDDYLyORzQ
1of6qMc2L+tcf/NEzo0Qb8Tp8R11EuSEEOiSc6Fh6r8FWjcYhj9+jvvfM9dplNFItULr8NzjM5TP
M1NUoOTm18tIE4jzKqpADQLHBigBfl99VLaGaYthsDm6k32bb/LcPr4ACEqzZwtmPbodK0XtHLvF
lLDapTtoass72nHna+OZbeD1DLCq2//ulvfGuBCW8Q3oDrwWnF43bpbIoIgqqSXxDD0LTGDh/6LR
YRzLCfax3GDaq5oJ21/eWYptsVcUQBfA06NNs7FjRMXJSBLCg+pPpUnidKCXz2R0Wb394+opQFHL
CrVOfgAHrPekG/M+2lj4/OR93NH6/fKnEYO5Uw1cP5tM6HZamhx6fERQ67lNYxdmaZ6usS+oW/Co
vNac5+YvY3BFgF03uvf3Ja9ni65qc6vbBxB5oh61RHBQo+KPu7nBeT0gdjwfgIH9FfKbgfCNFv/B
zsk9EHfGWxuDlSPcBB1/gWoZbC9j03POdLD/rz4Cb1MdKXdZu0M78TlAVUorXeCUTE/xa2WAWG9q
KWlR7HfZBrXqH60VQAPqe3fGKuXK5xxQ6InhnYjVkzZZs4gKFH4bXOUz3bE1akfAoKpyHuz6rOEq
p5oL2otpT2qSCvf1h5SV/EQtiG1qYIJ4+CM7Y72tU9k42sa4T4opcAG+U4Z2yLIhko4AYfVzathx
BCLGfZb1dhoKFoIhfroXjSc+geJaYwcCvgQFkm1QYT7ioseYCSMfelrjiH/uVdAU7jPnaJ46emkG
K579cur60aZSyMxKKWJTctEhoQwROwXy3OG4lPNxXiXW7j8mW9hqH1uTCiLYX+qPHI7hFz34mvxO
lW6+1x9Xs69zvCOp11BgRMtf5C4tFBGbZjyQdZ/v/ut48u1qg3OG/63efuR5SExJXSfL1kFVl/tw
clnzAXnQY8gBOmXjX75f5PfXRwcN7jVUr2eTVa4awChKfHBJdMAi3ciF+KmmLUMxgLW2eiNo2w7Y
XTBaYeACB8kZrCmMl75ptoACDjuXml+v+ymivEbk2wc80s4KvPydpED2nBgChMMDWInbGBdJJGpu
cKf0OIqeNxLkfPAVubC/2P0Ot71E46qk/CeUO+1s1BwCLXK2BroC+PUU1swM9SAqPhPCBd5fnFHS
WLs8nTWHveu5X8JEgTguvdWCji/0p+uizW5SiVaLg9AJG1jQkaToH+ulud9nm/Jr7ebNUEFGpCJr
5nXLY+E8CYJqGWWGxYAkrrxsGUqPOg5ZoxB2INoE5oRo8n/mvzdr4NvMnTqqlqdZplnX4RGUCKW3
DpMs7DjrHMb+xLxvxEMrssHq8ocS+1uOPZRrZGzC3tUPTsAPrHx9N4sxB5yw/EZX6ekqYpAOk6N6
jUXQMKvf55Bx0zz25sw3TwB8qaXEgxnOh49BToxUohXlhANA99N2PLAc6b6fAL3JgOPt5vzhDjEc
kQhtfJXVPE43+/es0aQlBwV1Cq5CNA5Abf8L1vgaIPPv48oDhpHP+MqyqpCzk6qUakCuzmRDpToe
kyhPrunToWSOmk4NPau/k6KvkVfTPFnXz0FtuZ8M+ybKcipVvCp18uF1w4feB9XfLzuZ7MYWOr9m
7cAVOCTVTt8ZoA3olvENFKRRH5kWu6AD75h0kA9iiSzNC9/o4ra/XvMRbrnlw6bc6gsEvFYYajNT
QbAL2RxXPrrE9Y2k+kj3+frwFFRZ9PqifpG1OPCD/95kUVw/HvJHWtLJTdL93OFilWaq/lvJLJ9n
hpUCt89mpLxKvssMaT4+0OcBpSOFEtm8yE7HNA2OqzpxavfB37p2NfAg6cYaexRTtmqdM1XEXp6F
mcOJs7vtgD5DW1jIqjICPDNQjQP+VprdbI8Jf6QwGw8W5TGw0nnHX7I9gw9/B/XjV4JDDSenJ2WT
yfXfpGXSHSTvkWYh/qxwgFtUlGAOTchdvHE483nCOu0g7bl0hyPSJccZAzv4eing3C6o6cidrxTR
/OSDrWLpVr9LkQ9h28Xqjsx5TFxGcYiy7DzzSdt16XYXKm08PmZEcSL20TbJYWP2DEHwbvjvYKMF
k5lK5GS0qXgW2ZsMqk8WCdyEo7iRac/gVGXUGHEOts8BQmT4g0CUF+iAOH7f+VPZ1mxQ/Pnz4D6Q
XIxwMmAXRNQeZOsyCCG5WiraGvv5xlavFb7rV97e5DLo6kjRLuZX+dsrQxbzueqReqYZuoUPCZIE
12v98xZ8+MIgTXwvGUKPQQmOP9qoefAB3qrtrFHTjCyT8aMdjYRlZtCiLijSUlEs7FsbIxxVmSmH
x75PlmmEORsmBwywvZOJwRvMvkCGjQo9uQ8PGP+VT2eyyQ0qf2T91yoUIixso6q769lDoirAy46F
NJ9xQqf0m70r75I+qqiN1AEyYQMNdSMNP4PR3/NuZwrIiX7a+4TtdXnDxpJVwr6lQkfPnVZtcAQk
rK870ncK90yDdhdTyBMFvJNCirtDL/GOielFCSWxBDTHGCKMMissHiSfZB9tjLr+LKbxO53iWeKc
9XevZ2j97vUos1XCCCpFTm9J63CZa97SwWnUptWU6l6elxg+Zh8LaIiVrMKxki7/JuSjHQ7L6/Te
oRx09/U4VvWjPEpMzSaHk47a0R9QZq4k+tbvwy3gBhbua4OHDOLmF4dYyUdQM2J7IutdJQ0fy/0g
oDfs51URaVQLOj/qaUBQOQ+aE5T8xmoZnZIsby/xXxiBvWjPKJIkk6o2WWQQnqKIxT595TISOBrs
XbSYuCMa6IIR2VTky7jimO4+ggx7vSl8CBAsF2vG+C3qs7XFFBFtxwDKD48uP1IUDYoJQ915Z26h
wlQP2CMjFJFN/PWcNeepYCfiYvlmNjDlMb9Yfp52o8JnaV2TSMn/OoPeKi3l3WOCTjY0YouGVrkE
ZfhB6A+OMEoUCjize1mCVwTp2BYpmllBWQrqDtgaR7q/0MlmMoP+bA+WBfwpPym5WZilSwUG85zC
wXb49P6qN/NyiANTHif3mYLvbBg34eCO9+/oejSfAXO9LBbAh2Fp6io6xVYiC0Qp6ValkLTathdX
PMeYe5udK7cl/S0S3R8ZUTTzbAalEPJ0Ett3hqs/oIAqw7TF/figsQoYofCNN2cqHQXL7Ex90RDH
SeTfMvvXEpnvETlOAxjZjNIczaV2+GO8CIFYmOyxBOAClKce8BwTl32K9tlr4CT7QcGUtpJRVhYj
53NwrNrZxWyB1dr1hR1cwisz9RF3Vg+OO3wt5U4H/iVO28apXBGteV+nTrSjZK6afk93ZTNkVm1I
vIjCURzotgd7MJNbb4Pu7Cl2L4xrHQvm8jjgnsKwqcmpvPKV1QtwLwMxl2uLMEKus/II0gJuxHgr
aZgBl/o6Zb4mFgo5mzbK6u/UA9CUN2foqFyvmX9xgFAbvemo47gs/bmiDSuqa91yLMhR79NSqMG0
j5VmfDvVUk/NaJu3OTjJAPpAcFzvxl3hcCpQhinoHDdcvYOF5U4C5doZ8uwB6wduVt0ZLaPwbrT2
CYgV8A+KNgmM9dT1p3Ynogi9IBvYxfbUPa2isxyrvy7TZDlbNJP2Zi8JFLI9bxhu0VyEE3Ef2sXS
t0TOaaNLyrRROfcg2G9YBMVdcxSKcGLqvbb4hfmbTAY7wXCcQ7vq20KUVOiqeiHHyzbIEzthFErT
jg4UaE5sPbJ46ptkSZMOMkh8BYobf/ISukSkMEjczBoYA+OoKDmvm9wBJ/gu34DLlh97j2h/yd5S
c7M5kBcPkngMXlpY3Zw4JneJ8nrgccqFEardqnakHAd2KwaEuc90GfppFdgS1WIPn+ViSokQSwSD
LsdLYczt/kt5q+OMCenfhnjq+yga0zXj4XTK0n+DfmPMoefEBXMNdhQoyeXBB4MDcdFBp3HqT4lQ
VynVQOt8cz1JavwzAsgd+bfjC+YXwJm3wowrf+oNnBUKdjAaBL83ayp4rz0FEuTpM8PmcMmW846p
SrGr8GusniprEljadWTcjjpMArsDytxgNuYQGKt0toaVOH05XM/Mxqz/Y3eBla+X6Pwcv75ysi+j
mr9DvGoVnQWopwxHEiTaPWZvUujnh/u2l6bl0jDGWbsB0tMU9vlQJfQDZEw8SfXCM5KFKxo9X/Za
CBSq70TEa0s9GZBzqWAQvl6M7oDngAvcYWwd38ICezGKSsnBg1YLCXzRpK+sVp9I0X3RDCJ7LSeJ
tu7ihdPlOvxX8nkcO+//4XHCz2DllX4szHeIuxgHW0Qej9bzjADGrritDCn4yrUxWWkS1kwR8emq
obn+sipfTD0FtePzH6nsKq1C15slCLp+D7sJ1cAhlNuNhhDNCnMJgvJSzmrZ1eZRuDZCrUAcelbF
o8r45wooaed6b5ShUquy6whcih1V/oQp249u8R/lx56HmHMG+iHrQiesWTBCTPpS3OZB8FKs57k9
Q4M8i6L0WUvI6SJV1UCJ14fP425irGgXYijMCLi+a+kCUI7U/zxSdlld2EwHKbW7sgeNCaPgA1Ai
LMfHLbWZJVybY7JZpoJQmnpjS8VzS97PUGvYyF1slihcL5/z0jwRnucHpEBv7+rx4HyrNgQYiMzo
exqC9CHLB+CdE3cteI7T1g1wdkIiumvD8DJDfHo0fenjF+Pc0+ixHkfeF29WijyIu/itpelSSFsT
+P5R6FdGiey7xtN9p+xaeplSIk9byMELQzdmL9lX3FY3wiSYjOoYRwbBxULxY9RTkQdRsdcJEDzw
h7+kFERjJHaKrAdjOtW4g2KEC13D/PHnVic06Gsv3Al2ZRwc5ffnCkyNp3AhjUe5l8PRi7UjnaNb
1zWwvoXe3WEf6BAps9WQWJaAo7KppuPNaN7zCVUOXT5oIKvSfQHt2neGJqb7jnC8ONDvMxT3o+VC
G3MPc70SgO1nKbLlR39AjfF7uei0O/+ncqqAYlwAYHBVP+hzRvU453Lyv783m8J73ruDfzqQ0FKC
A6RKhi/HCLX87X+HX/o5e78sO/8gTg604lwXgdcGXIPNZ/YJ19AOU069pMLl5jwY8jVKCjOrIkes
2rgrXD182dH4J1N9knv8EEv77HJtJoDf0JwYcyyuwwnvJQJ8LKhY3AuwXCjSkMIkeVXoy26GGEcE
QtS9zEicgncV2K/iujVFW6NfnZJYXOGzss0r2ZJzIFpXk1voL3nEI83iHJvbHg7lmeuLGeZxSJki
qCPqMtx2zgwEvDGINiUKyl6cHpyPNFGAG/F2yzTyadhpRanNToqFwpMh6b1i2gcg2DKcB+NUKagx
FUR/OTrnFQyEKxLl96K5p4xXlMREbL+gPoOruBWrnvVrHoTI2QYB897/XX1wEtnZ61N1BK9WMo6W
mlg+zIwHE0CsnzxWF2D6BHU4AavedIYtIHFIBKV0IZMA1WULuteexuqdKQ87M7+ulNjepx9lXjxj
h6X0tvToAV7R2sb0nKktIPyDb7pnFnnfbAhkCaJ66JMX1OcnXeOTBihOZyWu90Evbr+b3HKo2Fpi
3zBDYYGu0dzsCdZe6wY/x7CzUr9jtQcWOmlGigNxu8h3DEkuAM3q4ETi6eslZwdAazqHCz6rD/Vi
BUXjymia9pF+aertGX3alLlVuuCElLnivITWUOVG0WWbmscCO3Dnzult6uS8Guksbk58ltxlM3jA
xjdBJ/qbUJePbQpej2K7mxeDTukAijiBwwmk8bKIn6PidYvLx4Mi5IjnbnWrzNKjY+NIP740HSQ8
/a97fxJBycUyGYRytp9jl6BYOfLt6ckBDlmFdsjxlfVl5Z4ysQpkcT4YiX12mIrAmRcdtS8Ski3z
xERm/6sKOWdXhMCtTeSU76pBblPu9sac2lXlXL6Vre5upMhmU/jSE9tjn68RAkXM/phbHyz2l76m
G8OzVXaJQmT8hXCQ2KCYlk2SCoJi3Tu7zcT6XE4budyKUoAtsilCeZGxTpkF6LE2f3GvIyWzJB+S
6nJfOOHp5Tao6pPo7RbWJFdRyzJyn8bbJwkzh86w4zRLjgxsT8sdd4pmfRYUbmdGvX/Q54dWnxul
sk+t7fm/b2g9grg/CskTfwkueubgFx4xhQT4vK5zK/mldaOnwEwDrz1QnT8TY6iHm3dEvMSWTPgy
DlucZMMOyoMClZgKjSWj2eHanau1Ir2UfFhDibF3nkJMy7uREB00bUnolp8LgpZCttqIFbmTBPOw
KUQG7I+xFgDU9O10OWy9ioG+98zSJ+gZsk+kyYt1VIDgA5rkWZaElG1X7zL6URJNkG8KKqiK2MqS
1zVchehkHegNHNOsVAOgBG/tV71Z01yE9e3tDrcmJBg3mLZ6/RMxhaygZwLYXnqt9w293m6S9M+m
IwO6wd1PVFd62g2nzNs0wzzDoAc6IjHHEoOxQwJNbnk+2+zN/ZcnqBgNpo2RrRFdlfu5gGEvKzSp
qIrY+e4ZYU0LuWdRfzYvZX6Gs9lufd1LBlcMtvvsj61SR87LV/A9JwaeaYdNyrGCe1C8IXLiAUA6
eVSfj5nqL8PaOK+zkYn4bB+Bzcsv5+vslmwdGKbr7GFgS4Y5ErzVTW2iNpHOeQfaR2bwRoIiXGKs
1fAE1e/C/HYFEx4E5nrKPBkXoXWiB74EDsVOy8QyR5I4p8I/zfO9L3n9ia65mfmmucrYzrRoiQ2o
M8EfE2pqhzlhEWnEuVGBFDfSzuO4XwYNduyl0RWK9JTP+nvu5wbEvkdwe1Q6WkIhezovS2QmvNob
a2mi27tufsh1hrwos0UqWGH1VZKU/DTIoWcE2D5bNPrdE8HAfGxlMSrtU4NyG98WclZu3dVDU2QX
i5JHh89sNmYBSFTLIqOu9PY4yx+QrD36KhI8YIKIwZ/Feu8uz3B5TNXHfAr47GxhtBqJ/dTb+/9w
p6c89jjcZFnVDtuRNwzedN2cNVEFJNASj0jYeXQJRqBOz9tw7/dkb8HiO7q2CbrZKcUiBcpX7iml
a7rhgVfkygQ+pRpRQiobudt01BziPOty2cZrXromshP28QyCFi8b/uDv4+RJwnQI0zguopzhd+Ed
XVMM04bWju4TwCYJPJtzPJe89xXu2I8uP2zjRi3ki9gLq9zWuH2K4HEXQR0LV/W+iYDVIv3QecJd
+G4D0OEuUaK8CYZ/Rnlt8TQoV/6775PkMkg8v96n9C3MweYJXE/uZ7k+OD256AW1x9y+FN+sT77L
IEBiL3oh3fBsnTn9pE9HkJ/Zbn6MfpJZduRnD7oQhqON2zKOSQcOX/oydviABJakXNCNJm4wwDHs
QayjusYPyETnB/1ky9OaV9MzUQXcApXhXvQzJ8vskdYESwSSLjKOEn4KOpzi5cYy4V1/EmyKEJ+N
uKyFytPiCVR8nrk0YKOXQtBTYiNI+0PZxzPB5ihzFm2e+lfqJXPiE/skSCM2WCeg6dWtgerQtEEm
745PZ/ah5HKBulPAw8HZpGRFbioehCk3bA0UP/N7+iVquMitleNA1hAV5wLYsyBiLLCOz+VE8ZFw
rYv6BJo0Mla1kLg8sV7PAs+Yu+PYmnlnUooKdmsjVOx7gwkwb0mD6p9S/ce4T4W9ZB5TJDVYB/9N
uYLcbTgJk7EzKXMTzDd0W3GAfyVrf3chsmhTfGFFUCeOPRARtuK9pqeE5Li+JNEyjpii/ZAIX3vJ
6tNtWipCc8VbcBQ3xBDohw2z5LWu3sFtWMqZWUxByxgESkk5MvTKnjn8YBxbpwrqEErVYd4TKrPd
e4aljj1kc1/Hp77wNDckQk1Qvl+hUk3ND10bsJjvVUEeHMGjlHRjYNA2JFTmso2n0+bSDwGPaGfP
iP5PAGnEx5sQZIgQhd2xfPr3Bov7BzbmmXk3EauIhJc1SHrLuDi42Z4IUlaiwbuA1eji+GFRPsee
BAo/fpOOzfVvN1RWLy+EbF1z9vEpZM6qQwFUiRQ67qgt9TduKvdNsW8Scq+zsKEV6hcYnQld6GLH
MUcG5fj6TXFQI6/6xvk2tHedP4UMo9vcfqZW78Y/N8DWlFDCx40FlWL/4vdMggXQmiAo3WEjkjoJ
dIOiEz+fTBSX251M18LkkmmszwDxai5BvArUb5R+BJYPoXkEwqRnEayZ+Zyp0MRfczDKv8sbYkUE
2XDv1jZ2PuZOcP1C1CLookeZNWt6U/fNMh//bnyvhtrfdeTdyEQka/s4Y7AxCPnP6lTsb9wvOSvs
G8+cY1xQjIdvg1qQ06GMEy69nNIkbk31srlnJFcxSyvUXYqv8GMHmFZ9RwCRUYmLy3MhaPwmJwmV
FyubCzKRidSSKLEC7pC2MgIdujCROGdtjNY2LDnjCuV7nZzksxNF00vJof/T3u+L93B4yIp/ewFY
0c0ZcMoDIXtPDB6upBw6mR9NhfSkMS0uMJCf+TVFljC0nkRPWPOEsOUN3DT02LdCzeKUuj5DFLFu
+VUXbD0GU1GKJDxNRWB+8cQ+vVKyhRBhh4roS0ODZzGS/ejC6+t2qpXhDz2UMJfK3u5grwzm2YIw
xdY7rGxQs1ZI8L1iJQPAbbEUcA+0F1UAcgf2dlS9bkMsZBXuvh4PGHw29YET1IQbKpUi1RIyDdLv
WB081nv4YZAyKPTHgO1OxuwLKUGEwFWchHi+VCVJPg6mnRuF1C4xIuaIYtpod9Wrp4JFPKWyWi3l
RqxsJqV4fkDn4wKRS3df054rzQwYdf7+yPNHLgjckAAHJ97rGtUgGqC+ejGB6MZuwGo2I96XWl9Y
vPQjtH01KvR28QoA1rYZSMFxGyAzKu61hgIFdvWliRP+Qq6YogXiMm/ErT6YpakLhp2tYe4h1jsx
Mo8IfBrrBqm11blCCEytk1Y7kVH96hJymALCJU92emB1weCYjf9QJfEHgFAa7TNmoq1iiI8H+wFu
4gzmBbcc/CuoSAJOsyaHo82n2D3VQI7LGsxnuNZULYkL70DxYyD7slTNxWpSqYIws5WRO+C5kxoF
F7ypKbOAcbCwppqMbcXdyUUCCPcWlXpMoPN6G6qCaOIm2bdaNGRMUwazLWJkFtp57hfw0cuCYwiQ
7L4QI+U/q07Q3z0xkzcizfBCMvIRkGj7d687YZtepLwTiQgZvy5NBh6actMHnK+g29s//1htxeu2
CS2+wKDJh0zrTdKse5VCnolGsdL9kN23RjGmKo4pweYd+AWBy6pQ9FPEQGCqS/qQJ3BU1gVYjAiF
sdc0euQmKX87jb4D5diuF2qwYu1G8iL+QPMI7rXUIQEBvtD/gz0dKtN+WdI+yVTHE0d6ooKYGbGf
KB6zbPd+cFHGW5A5PHiN+CiqCgie2+HdsDELeFHtb6hagsnv9BV3AVPOxfQZSdVXTdMw1tW123SY
RKYA8AH+cd4Y/eV2DeFndJDBM4SbMSbXmgI87lOLK5D8jh1tozI7+ZglJkvuerq7YM8YOvMhEMbT
f0qP/YWWKS26k/Cq3aGHSQC/Iz71n/FU9uqiT9aum5Nr8C7bYrHnDIjO64rENdLl6dczxyNEehc1
yHBA+CWYOfYhiXYZhce9/tuDrwZ7J5oF9iOty2TeGcDPlD0l+Koo15fqFyb8syIx6+BQTxCFvWRt
qw2PBeIRrs3Lf/IpCyp3tzPRZPwZyBS1LzfMCOuCeLSmllAppRehjipl+nlaugrG6Gix5sTGDh8d
ODqP9HlEHywU3bolTx7Z8UHYvBb6FdIpb3mYr5CWuqL3QAvfSEwHYvCbk8YNrMon3HzmKzzEibIJ
vWMEn9YbtIAKHJbVuNqqZmN1x0zKWRInOxxbTPEJ4ORNODl9WN4BxHKIYgFLuGHZF+RLgklesRPr
0bD+1WmB3EGtZlhsH3k5KN4CLYSlRg0VDHDx5L7NExfdAsiZpK++35Uuj5lfHptDg37PhT5XPBWj
tMY8psB8xLjtkjNUinPOhmYrs+L69LhoDZArHHiin1+P1axDqPeAeCQjYFxjxOGWD+Q74Wjb7z0L
7qg6zwBZnaLGQOLiJ4W9sxc3Gq13pD10mnk+UvcUskwjBRdxgwAEtJgAoot9+cQ9I/nnxTxzAkb1
oNC0C56iW5UvXcKp+EyAwoKucIfRDc3hVRSQcOuC0Xx7WBmcg/l/9YiKvpwjnvA5wUKrXmdxYqxk
ihzVkyFp9QfLpnjLgOJmchKd/IRxwc5qlTsH7O1049xcNc3C2n7IOrYUOMkfRgAviQEBDf/9UYe1
u3Tw/Mzh0YAWafbUSvLVWld3CPQVSTlCxM8C5uGbM3NcdAxvKhN1rcjzstTq2uB6fNHdByjSiXjI
UH+CGyybb8nd1PmZKOvNhn7+aDTFHp4priYRGb5yr/3cWdSqSkq0FaHN2DJn2l68loSm/HXAdomF
vcv9YQy3UMOcnkfGbtQhWmJmg4K/lxugOIn1+Coj0pq+8ZenWZ6xSaJw6gt1KzXGtNzH0K9GS1Rz
gTprz29tDJta9UEzasCSQqPgwFluspl+jIv05FZkgpGdkGv5vNjHrFm2yaNHzFrfVOMcgSB9kjnl
RSpDI/N092STOFG8OS9Ly11u7WdAc1sZ+Qaxzc+x+khX03M0fSZs9J92xS2d8dngkhUICQrkzodv
C2RAj3FxWUK3ONHd3zusw6hWCB9WD5Umqs7W+P+6hyYmILh05KmZVLhiptppobom+4sPF4pSFayJ
MhB0xAulzajJA/92YBXQIjCVTEgSVgllPeeDeSIZvhzKmmGSRJSEptbmpz5Hu8ZHyfhurx5joP/k
veyw4V8yB8ix4AzJsObA2UwW3X6k0LCR/4LpptSLc07XjSE1CtP8D1dqE5d2QErqtSBALQXOZQvo
bplVQ9IU28rvVyKJeWHsr5pA+EEYnqhBBDsCqIzrWNnUV3PvmBJwIUCHjTAO9joCWDhUsfQKKaZR
zScf4PKktHk+L9FMyb3wWh3SVbT9iNihcHbnQiVjzCxKPDMGSkGsv+pN7fU0pRSRS+x8iGI61oWw
g4SAWetxKqPtvMCOZuduLWdPqx2OeWRD/wWJglQNI3PhUU491HQmbbcVkTZbSA6KQQUWbfWxJpaO
iJiNj1SGTRbNf1ZAoxJK4HXm59nVWbpJTVjhG1TnoINx7zZV2K4BWM9BXbVrSuveE7Cz59V0NzXh
UxtCJtgYfi82kD2JIe1ktTi7B1OSpH4cdcdQeNRBaly/IWp4l/VWL1Utee2cbQhQH/1VxNUJKCrz
imkt8wxGjQZf9a8pq6ZIqawFBmYjwHFBtEjEbunWiu5bVXYLSAXdWhFA+wVpcLPU4/KQ8yr3F+HB
TNo4AOtDExmphRH4iq5pIAeJZEJKJBMLuj1js9VjcEzWBAWM+EU/b0pGxyHXlaNkA32pHEkI981s
GMfdY/axMoocPx9A5YMWRVNmWodFHj+fPPgxK6j1lPUXzGzDI3+V3TxEDjSA1DOORNMJGoflB0T2
Kq9TrNOOnojC4CbqyF2ouz/65ZAEtT/vNYlnbg3b2AmQ4xemm9ZlnumOGWJQblNLJEVv3RZwwtxV
hJuURonZD+gHcLuADm9TSSgSuwibLuR1CKUgxWLK1rwSK24+ZgjRC0qsM7SHahCJU0DFLLpI9Z21
wDzSLrHpHeMHKLPwwo1LxmMstk4RSA6EF9Frur5x1zI4rqmb6MpXxO2SAGyHWCXhREIRCwSCXSi/
NQVP2DOW4T9ojQWM8iqecw7S6ai0q7PzGs8SQQVT3P1kxmXaA3PNoXHS+pAeh9W5syB9LX3VbocO
hkXIDZ86833Rn3BJOoMoq0QtLwGsyp4XppkNWXMtVyA9yPDfViDaCP+vnwFECs7CHHXRK/Q52nEu
RvTnEpIe/VwxYcaeEkb6P9h8V92721z8ckXCI3FXtKYYUqkM2AbGKe5JZXVgYjwcT3HMDhFIIDpx
IYvnXHWwLcka+I3hj8nsMjrlaFIw1WoAQGk0uzdSovhBcoox9CUoe4xt7bEUkpi1DKfORdbEL825
qR6ZUEgL60cKRVMyPvS9vaebknD1G+na+0dsjIys5Eoi6RxOEQVQ5QmuYRxqRgsV1dOP8UeSWDvo
WZpbqfCXL74tLgx+RSk53KFZEVko8182pRxnNvkdMoeFJlGgm2TeMdVL8XbMwaxA4333PnW7JB0N
WD5aVrKENX84I6Gad3/4h7H/ixlW3F6NOaS9Pya56QZCfEr9sgEtdW5Qib1mvX5vWjPJVxsf3aJc
FdO1uCe+XYSKoRW+gl10LyBv84dR8glfbGArwAQKN5iNWYx9PmUDqh/7IEIiUgsDsIHuARNmvvUW
aFKKELRFIzytGSssRFhx3lKDAKGQzQK6uK0TrKX7XkS4yWDWTYe4KSrrGGAD8FKwE8pLLGTA4P8r
V+mvEobYPWGReH7KtmmKcTvCgnSv03t6oExLV/qlca4okbDXuTUozDsOOUwppwSc3VjadC/Bl+oY
OEZJ0d9auNBP741CzWuEryl6QwfgmjXLK6uQlxxm9iq/otDkPJeTGtXTWW7PRiR5QjQx72X07MtD
jg1Vq2EOywwg/JwmVh15M3qTkHb878PRXAQ+B6QflV8vAPcaFEfq/ze8UxCswA9zRbAbGbf1Yz1V
/36SR14mczYg1QQAncrKvYASlkqjEpcfWMFfEtEoaYErlNyxFAHbCfwsKLW3RRe4Hsv/6IqzsNsi
g8iB2Ia6SxlMfO3Q8sTpfib/4PZiY6UErHpkfs4VMVI2Nj35ol64GXF7+2wzIWBQ8SSsqupVpEId
ep9w8ZmEOdZKP1l7AdOEQL4y+yCIXim1qMw/izzAf84zEm7Cu2t5oNyoQIBkKFmbC672UVfg8cTD
Yw7781vW851jiQfIuIxXFpZJJrHCDykaTFVVUrSxNyJYzo5e41mzi5gOJ9ZoNcdYaevALWJLJgp0
xSl6+0152TLXxKwqS05+PC/cvDB78V2av1cBpgRV1LZEdqoetTqPkOyzwLmudAAkFKQJK43cEFBx
5Cq8N/lYKwghFOj0L9aohKZ/N0IQ10FO4ZiN5wG7OLZ27zm/CIFNqhspq09qhdOFbwiTtRhIlcUC
edneT9WSGf8J4vR8KLwxAiS/9QLnjXvvetYRdXJyuVL4YptHMZMGLBBZ6LVAWuvuJmlkjE07iWPG
cA3EaRnVfc2G0sFNRUSdp/ymSm8jK1IVwuBujkbDlfroals2vRUaN9kaN1vPp5GbqKoNoW9y711S
LMJLJA6ajxEXZJFUblyEMRQbO9KDqV+eNzMhUdQE3wsx0OgiTk/wQP8udQQ3YUxnVrzzAiNCOy4n
QsMWo2MLnwMvhea8z8aic2BEYi3bKiW3OGY7MKzFqzY0UjZgYu5GlZvyIS1nmmHXWeFG1JgJARt2
yvP6cdaz5mPrc5AihusbIBXAXS3GSWz9CLme0w/kYf5ZkhiWHcev5rGCNw5t3A6DFBjBxCJ7OeAE
jcUG/z33acz6YVhU3W4iniA3U08vA7WBcoolwpP2Lk9x2CdY1751bXjy3B8kpWMNZsCg1n5QfB3g
Be2Ir9mNvcjR+mqm9FBmHQ5ctnaFIHyZm+KN25BejsWH7+9CcFwuR4U9gNj7LPXB1kyMxQqU1pw8
PDwIV0Z2Y5Hui/fY+c3jwR2N2F2LPOhFnaL85hYDVE3m6xjQudrTGnU3gq9BtI/9R5hnV3Kz4vZQ
fyPynJxejL0LYLqgYHmyOza/4PD4qMGwJiEBeOnZYzPPvph00z2OZvSiAybYUZ4wzU/HNwBX3F8K
AZOEapVVEsRfZewFdUkYDwmGDcj1rng5ChEcthDvwr7o5e7JVe6q+sa1oG/SWv2uc/PtHVu0vTWA
pRRK1z7EIBgBeLFr51xUKnqgDDGcEVYsGOuArG3vb4UsgEI5A/ZDD63d85kEiMSbzKPmJuEe33Ey
+egyf90rwi/gwE0WSvnNVXlnckYO897bcC8T1kc1YvyDztqL7h0DRY9RC97GZes6RD/39UKZl6Q8
No5ZKvGJLf56egbBgemK92hR0dvu9hKGy8dj6SGE9Tps0UszOJJGnHg9TVe3dr1sphilDqoPLReP
9rd4g5XI40bs73dAlyoy7xHciVVCzP76SSSu1QebWAtxl//Mf1fwvWrXqBnypsn1NEFaeJoYLIeX
jEDxFADaIO5H2lc9EjiibvWGxfCxfR8nbG+vuRb7phxYDXl9U4tlzdEEO0Chb8ttXhwA1wCct6ej
mrWJjYbrd6YDAtFDKdBKT90FYdLdWDYGWa6sav3FYVnkt5yaxeoCLr+gwPmUl/XilRHVWVmLLZw+
GwEp7hUjxGsDVB0phn9m84EX11q/+lf2XWdu2iLBa43WsR1hQnItPRcH20rnRpPjHSKzieWeSkrp
3YldGWcWWU2/XANZQ4qCVTtJvcb42HdjO+cDB1w7BXntiGxrHrDsAZYSwaDA89knP8rdk9yZULAU
GhepsFzvvRNFOYxohz9hKFI5Dhw1TloMmxzDq9Ioykxlb5beZoMWQ41BJQ/HssangZwYHr5h5zUB
CpYSVPeA8b3DScs3HZIuygo7n3Db/FEQ+ePkNmUWaF/2U9+4WlV1YfH9zUO3t2QJwuCelXo6DcuM
YveN8rz8/WMxS40qudBsBwHI2qp2jcofsjfR4IgD99W8M8av7BOGkI8R4EKwJ9YBOPFjuUR64wMk
BYeTIAlolybmnhYJzS9YV38Uflw7AZrpI9bAX3MmWpen8Jg1nA6reQ391LymW7brqAxwpIc042pJ
jjKUFvrabOP4eLUOsrLyBw2c24u35jdvOp6dypuuFE6gLEsaEseDqZmAXkJDfMB6NnLU3QfDm7Zu
hN/FdvLxPKzvSm02iOWHO9oYTQt9JzZDQiF/vSKa3rEIv9MrQ4ewbbcn9/q6vp4z525OdObA2TO8
/mEbfbxrE+nVPiW2hizwDlrgwSoSfSWHN3Y6oSMyyMBdsaXnHe5J2LTFnvGVzrpex8vTOeXf9b5b
NpRY6YWfhtF1mWauj/azA4zhCtgnGqeygPOWaYwxOXWk7gENDKxue1lWAl7+C3CJqW1IRgijB6FE
VkmaZ8SI3AYTQvhF6dmR7/7P6uv66wq0IxXFqwo0d2PXIUIfEg1IVvUTBao4BOgfKUm7T4mb4ICz
a0mF+OcPuHUaMEoF6vNVIznGkzlS4H7ubMrD/M4HeDAnQSb6+b3qp7/d/Hm5W3SBlEhxQBrbOX4k
jQOyacpJepRKQTEoZQLgkR9V5nL+0lTx8H+wRi2Uepmqp4YsCQ3+zgBEhqadT0zk8B/gHB+g3y0U
0YEvLy+6FonRZq/DMupfX2x2LN4yiZXmydQ7UpW0oTgJlLHYYDXLNzrav4PQmUjEF/eHq7bk48sw
h2V84U2vgBB21aU1Flnadfi9yjAc5N+CetUaakDpXuVxjtzQnDXvHepI8kBZtdqb8fd6FetVE7OC
h1Gh1tTIPvbx8AFqcbwQHpy20H00c7/pdhaxB5cevx3lnZvxQ/tXkz5Mt6vbIcRiGKealjzEW0GO
rT9iF8TkyOG2UOYl5gWO77sbEtpJNTg+xk0JzaERxYwW1AxWCEIvND81yfzLd5A75J/EdBjkBje6
Kpy4seNglZeafcjug1wdS9FqdriB61fwj4BhKuYN9oIiZHKFYkEtwCnyJQA8qehVS/3Cw8abPkoy
zVdPlzSIiToI2/QeSX0I3kApSWo30V5dfhAtjRNqRBN+gN4IEMQ1aIoc7rQL8Ztl4CmqYKYQtMTn
XO9yhstFJWQ9PdrjAzsJbir1abhW5fhWpSxfXmcRqDSrtb8mTatcSU15UT4bTuWOki+xT+pjTzeZ
16yaO13sSMveJ4JjODe929Tm0gopS2u+cMvJobQUMgWQQL9FTaf7ElHTPqv+Jhkq/e8pHxuLe7+i
mS416m9chN7l6yWi6LGP0xnOoCtbWHtXVylkItWb/htswLrHVWsEz/kDaqFwXoGVmHn9tZAye++6
Qp+8qpLwnPwh0sP6+cSpo1rs7qP8/nXCqVOILXvjC5yncHdfxbZgjeOdmnRwhydLFV93qC5rqd/0
Yl21CiBIvhqroTOma75t5hroiDPisKyZ5EbyvcHXEqMCUfKxvGiVpg8TZWhrpD2B0OLa6BzEB0Hu
Np0NH++KCqkeRF6iEyKYsA1pQIMjZ+a50f9SOss4cHRliRSA9Ujxncua8W6PgprWv7gVwvIK7VNj
FYU7e4NvEWeDw7Y+0VWubaTP6qhJabUURm+fyoM9dbAleSP9Yw45bVyefL0a7SvlyoSdwd54Gp10
jcTGGKrrQliX6aGV6cIq6trB1uIUUBSUOgMGSaK1Z2kKXLQ1P+sbszgIHRTlncZElGoHH1zzSIPd
hwIldCCT/EjmkBThHCQ12/pkxU7cL4fCmOEFHR+/l/T6kV/RSRNGXKvdKr8L4cSwpoIVNH3ihgZV
l+js4m7qT6gWlLQVAR+P5+IWg55EYvuqTqjwEfL5Eblnoi41iTXtMctrDU4M2J1brqSOYW+ibXDT
AfKYCJMt6WhPDRg3kug3AKe+RKuI9zMjQaA1SuB5k8hMQySpisI9VLykE2dD0cn6LojDJtEHJEhk
UKJOBvIE+86hy0KCeA/S4MaipcHKYRydYqlB3HnXdnj822+xA8K+xVIEYkFKsMaAKx5eAZhHX7NH
ge7mR8KWapzPoe32XHyvIb94DSGV4dgeeXbtLMyA9hn4ah7yarqGViAECCWsabn3zBpGH7OvbfIi
/cvNeza89+0hVzyX9A8KaQwi5grk8IhbgpAMFY9qSfPyw27872vWnrpiK6t+gDchWbZN1dvJrrzT
uzsdpYgPy47v3xZaIyeJVuLcaZW5K/G6XxEhXpDw821J/F5/hk3stPn1mRjOC34OIuIqbw35MMlW
spw0sxExnHpv67OvBMjshlZWyQF2Mskf2SOeJ4s5dfuSOZLZF0VM2piuRVXBWzGIp8TjG2zSpf/3
Q8XgB2dZAf9nZ8nuADbaUSBWakGhk9b82QiSojuP1k5S1TD0omVAj3atsT2/uzR2H9A7rgw8bCAv
DHWvDCGYf66HnRZbZkhG7rnF90k3iDme4DgDuOOzCa7hwYga69noG5Ve23ZmhUHcwgmDwl3FC8Tz
AN0OkRcb3kKMYAmXPmJNoagUORsJoEe29FN1wNWVixCf2CA5koBhR3xFPT/7jgTAotYehDVXyZBc
dxvoItjTasWH5U4XuShDKjNvBGQiIjCApRnzLKWzKusUTAF3ij8j4qK/DMoOwpoVoznvSbsfgj3p
zz2VFw2mv50XrTGlYQOETe+C3J8AaFYVk7noXO/03d1ESPWrnDHo5epD34yi7zpZAzIQmHTSCVG/
b7o72n+lwFVIK/VXSuCIPeJt9apV0JNWJdS2tCpjxRxEOaXIMkSXkGCEoxwvGK81/fJTj6cfJWX/
z6T6gjDRX41CQdKexaKj5m6sCCitkfLI/RB6tklrAUWPQlhIyP3v6dATTMKiGpbonIfh1ymWEtFC
RhNDaAGxV0tLjT8YSOsss5VzCpV5EjC32iRv9b1m5uGzbeypnuNqJVEDj7T+x5sxrjYIjltABPGj
AHzVC2v15Nk5001iYQDn2r+28vIcxpfCugAFMITv9C4/i4EMHeFzIx3CJjglWZaJpjS8aGuTf1Rc
HAH8UDCwU4cgq5a9+Nq4aJGRegrz9Ia6zUCbaqcAZukoZhnLqFJJMidBXy4YJUtKgl6SnnkxEbDF
qdzuKdMxm9dvAAmK7GkzBqPcEZOJ3GyiLJxc18j80TKrMvG812/HtOtP2R/79B9oZaGH9cnywFcm
KeIbQRbnnpL/FGg3quKJb8lbtRo0YOSuyNaZFtTKCHZuA3kYyhOzr6eYR1+2iPBoT/EJagtJOqAv
s3YJ8LH5iGhTYQNytluMiNoW4HbR75qf8GcQdyGMTZOHZL2/mbonumk4YTK5ASvzZ5at406Ax9aS
sfLLYRdEB+4CP5+YWRziF1tY6RTEpDw4T5J8lTm39uuxStbl9Xq8aURgciGFzalzZlAew0FAE5re
Bld+blBxNQOXECWLBnkZ9RL1QiEMrBN3kiofYRTHQ9kZF/JJ4zvotlH78d3zwWC6BLi9lde63GMq
xFT8hdaFDXj55J0T5v5e3DVNQ4RnHJtsxksQd+Gq57TtN2vSN6NdzvUmHa7dw26shjpbJJA6YMv0
D/yJRm/KNKPX4ndSUdoQNqb+T48wmjuz1hoaNfRIVOAgvmp+rwBHAl67qYQ9e5w8CL43dvISV3Wl
i2IBoSZXabvWcMbmuxCnfN6Ne8A496ddY2C8fPkkGjVOP7eZwX+qKk+Z9vHAMlMvJdydyyMycqnz
dWfLg9s8R9Wfq1RCDuyx26PusMK+WxqD99JZwPie6Gyqo2YIeMZNHEhs9d8N8SBTWCYd2l7iyXLl
hShQeeFwtZT2/fFBklw/dQqOQdQD2r8CBCJlotTd5YxIBQ5wIl3WiK69ZSHt3WJ/vlOL+6t8XSch
Vvh8uwIjxxHaGdLHLeTQsGbNSvQ3r3YRVHbkVLJkOpaedx7c5wZi57YwrAgXvJDfOeKYx0XICe5B
3VCtVYUfskLc3HK3kQm2A6rWqCgeCSXcfTulWfnLKs1Acdf9hHcR6mf9N970Ulph9sy9MKeTGgZC
yDnt0fQKl6FJYQWekLfRJxEwggMR5ZnyVdfqYaVnWjcnuiU9PY/En55dVbRSsGr6w22NqqRpkwTm
zl444pPRgCvEtBwJNT7wOFhvHg7o2mfvpmGK5hYeWJdLFFL/3r2k/SWoMnEiIDbLS1jGV0Nv2W3o
5mTuuX1qOngNdWFcb4Do5CFhT3kX4Veijld4mT7m75/X5/zXCLm7VmhfSBP/1LK/agkA5paQe/fp
KQFdH5w0WWsjR1S5r/LlvO8cQErtICDXJ6hzinOPj0X90IPIk9GZDnz/m+ry7wi/+yAatSkzjrYP
tHJVnEWqLKpygGOxuq9Hu5AEjSG8SGtD8PuPLoLNWGJ9yCuzwSdkJZIw+ZTATLPdFC7rtvL+h/dw
s3z/qv2+CsfY5IN0/CJqSI9e0BAwSWMpEVdCwFDqqylqws94BW+3XM1wUI3hH+fA5/Her80e26kj
3Gx2NvlfgCAyPXHdt6mREcOXKGi1zsaNwppfjfnJKtOncqrvSqx2Qv37LqK5mWcEwYDyVo6LaK8l
TKzTB1wS6Xzsvixl+Lx8ocDsoIEfsxdT0wruD0Qv8GlPUSWGCzMd5fHaCWQU024L6CXHoKpngLs5
S67MKnsSduv6UNgqS04jxZdlt4zTJ+Wx6+trxyBKR4oebBWZwQICXVOZHGDMJC6emRMEkmNzk1sX
HkaShJ0+/ZVzMtOROsvpVorGOqAQ3EMl8oN46DQ9Eg3DRQ1BB0j0qwK7MY/0j2xCa0XebvZVfeo/
BBWXidT/3KNVH0621oGsAJcm+9OggSMCBIicq4H18N5XtIdtiwrAbuxrJE7aiobH0l9xaVqLmqsu
A3xbJMVB5ZaChjxtmFd8R0J45an7bYQ8heOwklhFcoPlBcGW6s4zIoo2CZaam3p4I0lJHQFc1eoT
WmVY53XIzQY5j2dHWKwyWQCMjtW5xcaA9HMy/ZWQp6bLkGCXlhcmEgPywt9XS/BxSS3NkpNNp8Lb
B824JppHajRxBAuzr5niNR2Ai0Tkqdug1HUOt1joK6+opFzokgTkoiezLxBWQxEzP7wFwdQK7s8i
GHBajVC46abZZhAB356PmqpvE4dKPWxzJ+LeEI4rpbx/QjpP1T+x9G+DwjgMMDLrFZwYZJ/PMbt2
jHvEBW8K+ZhPXYJutVEWe8A3VhyuMW5GJCodStXTgouEjZvE3er1ArMD//mGzjYKfVNdgOiEgkue
jjLVoBTp23SLb//jl4AFQEJcZP5ubSb8OLdHJwRkTfm5mbi9w9Wq+0W2ptjdSvdxTXkKNUiIx2yO
/JnczBV5G7MGGIym9ilO4wSwXdLQRBJo2aiAcAbCV8dkRJzjKuInTieaUEYNY36na0SWjQckKLMJ
oHefiOCRslh8MJ/xQ5m33PzBjDHnsO3z+5/u8xNHQ/GYx783Jg95ZyaRikVJf8/W+05jQNHupGnm
UFDqPniLf+07Ju43cUGLG6nogrcqXaa18tEzJlZlYZ74chsbog36laq5peQQXLCO2YBkrnO6YjB1
LMQM9/bTx2sMXeuzdENAUIIrBXFTu0g5xi9vPC+LZjMpGjano/dtxBLaJoE4oTP8xA4oCuAEqA7E
kjTCLH8zF5Z0Hfcj2O7k74bfQNSQVwu/GmkY+yPqYLbjKI5N4XNfpD2/CBNFnLhppDaYJoL70IDj
TskL+3v7nyT7i+YFxUUeHwyhJe5j6Uf5viks/m2WaQygXuZLHgq+pLW2pN+BffaIQHLIaN2asiJr
JpqvTIQ1yt/LsehQI9drLf1g+R3hWn3oPcQXCKvfw7n1CZMgTvXG+Mh6UfXwm3GJtZE+nvvtmmSq
KDyh9LgobjCf+kSaxLOP6vM7gVEs9C+IBOOFFGt66jajc7nPDGUQmolIblm3zR9owOdGlDViP+0q
LuoNqOUKUl2QkfkWsh2tFk2FAojUHOiZIKJouEWlN1n944vUwACH3mng9Xb5K3N1xMHuYqBTR4NR
ICpj/omYi/08FGquaHAteYXqI1zghUpRuNBrSW2JOv7cZ4Oc8Br/TVskw62Y3RQ/4DUXBau+bAEu
t9HDx2mL7W0j1sYFzIXiXdfWtactjGN7h185t7ETqCx73JZF8Fpvr74P6NKM3I2C95g158LOk4zQ
38jQIrxS3Oy71f/aGRKEZl4/gFMR23tns40RHhl1kBb0GkojyKbRiRikcyKok5W4HtmOoHAziyjp
5j7OEmf9eLOaOubWIKvpEQasp8AeQrqI2AE6dj4oeIxBzOAz+K/KmgfRFnbz4d/TzJmLx8VInsye
YpXOrl75Mv0H5nuRdDrZid9IAi+SZt5bqyh3IQRlmF3wFzQ7YDrMD7WcIRJpEb4z3BdG06KDbYsS
ESmzWa9w5MDXD2k1HcMto8QVheZIzgbh2y+BN8DK2mJK6m66EfnufdupJk+Di8WgrH9qRJNBKVZZ
fn5v+BvqbOT9hwVVtB+VehUH7sFDp7H/9Iji/NW+65xuDf4YucGj05Ts67BvsYUyJ0/0GWYvfeFm
sECouMhmQp4HwdgFWgBN9hyYcJPHVwOgMTNA5iiEWEwClu3oY0+OIH8OH85qOU7/kCqIPX/ptaCY
/+nTW1NyFwUCXOu+aBs+vbxVLKCVvqfLubYy8PYrUgmHXs+3TqUtA33UHzs6THvum7rYceAiX2Wc
skaIIC/lAyj6eNO5S0DuYdHb6KG2gA6qMOBBh2Qlcwi/9MosIBJhN17iNMM5e930U+Mgwu5W9CkZ
U2d2N35NyShLgKLGQWw+6O4joe1roZ5HtTBy5FYePZ/LoJ0TQPhAhtpe1oLIcUDgloNGgbEdiUzE
Ec/3xgThlLX8b0LbDCt6fGu3szB7YfafXLRS8Eck9hGz3PzeAhfjR+slWEKoWjHNv84A1dVqQ8dt
6r7cFqzRb5Cww+YG5stoYaZUYBo+9iRk69BzJX1ygRjCw2idk9sUA5YFJndzIam8W4b/KdDMm/Lu
vWmJfrl0QXnxDMrv81Fp63Dz1pjXsP5v61A4bgjOtmOF7zbH23MBKNL3DF/+vHzD5D3v9QaresCP
TaceJA9Z62PKwIn9uhtkU7XrUlmY1iVpHLIEAdLaBaiuR6vAGH8qNOCX9hk+/NN/u36Q9FANKngP
djfxFUQqtE72TOKBGdel8LAIwodR8B73E24OHq8BcFd2yJ9g4U9Vb2MS+kiqYpxPp606D23Ju8KR
Z5FZcBTYHKcrM8JVfCoAPvEmbkyP3lLXNcLN5evhsnC8X0l27JmgknSeLTDmjIDRMPc38nUnXoAn
odmSK9HTDU0gIG/QipJgM2m2DZTjcwYyKca6dQIdrPpEO8UMVH/duxOeNvn8Mq8MKIqdSJfNSeQj
McxTZkiSuuK9n9g/33n3OnNFQZ1QKyyNPq7+SNupLfN9An6wXswF2XQzgF9pm8c5tpT2H/cnaSJ3
cv5AnatGe7poUPJVk7tL+VR4THczpXFZdG4++QV9JiZG/fHcFeD8RQEW/0n3xlTJ//hlRLbAb5UR
D/gbf5vjulq9RNCUdqH9JEQyGViGkzJSoX6VAzowgKgbbvLxoO7Th/vEIAFAbP8pPxh2J5cFmTEF
fbgomHmcqAtYl5b3WDcC1fXGL/Rmim/tCb0GKQWJiNT5jEi+JSLJpGpXb+VhZ3ehbIczzKOUAIHi
sKMcfRrv9aRfK6UmsVYHnYrLamXTkkGSoNCZOT1XTKlAlgKBnnDjr1ze0SuXdervwQ1yH3m+4T3x
wfbOK189dCnfBeDCbX0+V8U3xetBVtPXEV1aAEQ8I0wotiW5K7axyImsOee87YjbSauvsnYsPR00
6R6L4IOKnLNjn+1MIs2Zmk3eK/Wv/lLo9Ai8VuQEJhaXqLaSfksmC0TAltWvg//lzkmq+StAlfum
lH+M8JtxyoKaHd7AK5gpYZTOaUhOHcaqcc7GR0UR9SQk/oxKEXDATJdoUe3BDjSfHRd8vUW6DKp9
e9XNt/e4PMCs6HWMTkimPsRRjjJrokfrIYIXeBH5bySFU+m19bhI6vmJvub4L/pMKIvzb99/tQAr
9N5VCKP9wmOoc+hC7ZsShjkvnKz/5fdtw6cWicWeRtvPJFkT5OvkOZcFJ5wNt9PJTSjHuNvcJ36a
QShcAqvBLt0VhD6ttmceGsmfHha15Ksg2Vaqxz8+X9mA16fLUY/s6pmsWL7jEqR6hWPfUH4ZMAr/
vODmqpTJtS+mbSfwHjm0JJkHbJ+OfjXCBZ3YizRJ/Y+OQV/b5PbjR7FpfYg5vb1/yhBWb0lyDokL
+ivQmhBwYHOmCRbWbZoTkP6nzns6otY4IomZMF7YEHfWIdqe0tIUh/uby0P9FQ6wvbrrrr7ENvOr
N2njVBc2oeCh8VL2C+AWU4rGaVaXVxPzFvp5WuEzWDqCk2jJObozwZfOk5+kNxnKXf793kgor07d
fHB46HrQrM+yaJauONk3ghTPy9SxI0Yg55HzS8jCOq52ev4/gvZEtNZogeqUzxT2Gxukxdglee1G
fNdKCLT7akcKSz3uYNOqU6jBH0EpDKjjMqiA5OYPHE/Fi7RKrDgNY8E36Gq6T4//Pb+UBthoVsTZ
t8KcIvsajW5BS6HTWj1i1cw/cNYSnZ1mG4e/NbCJjDeTl9JL3bl4H8q0q+6REWAhdNDS3t0QQwQl
hX7owaMsS41AUsP7/VPG1tUj8A47J00LqaiKEkDKQqFMmR+A3itEqLiuy+FQcuK8qhYkcqBJPP1i
izBcCmb0w/9w/3vlH19X6h9nCgFTwKZYT/6+oElaOrjlFLgYMDh3xsDe+inUJDNPP6pknJek7WFM
EThoUW3u5b+hKOg4Jgf5esVabLRM3l+xaPLzPAnVnBZ1io7EndRmmmsfZpy+No8inBpe/gBvFLxG
fMMOek3cdvgvMw+qhijMlSggT9a1B356S9tqzdI6UkCBAQMj8Oujs+FmMbzoL4fwXQV3mGH76NAs
S2SFv4jiGXXRlZslPCbu8Ev5b+9Zga/QYrVzx8ggBoi6cXO4DjBnksvQHugJUoWLw7AgLpFZiosm
JZFbA1MTEn9en8qJtUPSQyoOzm4afjpAkOFLj3LeK79TJast1UOHEr0dXpPi1UjUEks6NSqA++JT
CrMQxI3IgEyNghZqvU+Qbw8Lew2SaO/LGF9Je3SogTzTsZdknj9sm/rwCRV1mh0uYlBPpXPMp4ap
3OPuJNZFOIu4pgESMxIInnvvxR201GFJe2swN/aCVI0OgSRk1bsvv/JZkQSKdf3DiAy0gWjuQc15
pGpRhFCr9dGEReG0MjFDxsWhCYFSSnkepO4A0CXhzWDTMK00NwqR0Gt05NgHt2hKgKp7erkmevh9
rJbpQrkolcshYfIE6LPIof34EX6Fbw/bOUIezDPMVg5eg4Fms1mh9eKVq5Y//r61b3+q+XOYCiKx
6edFgq8PyQsFjBCOTJOVcLPc47WOVoEUV4JGU7IGPMy4o4HB7W+EQ5shfh0WLC+I6hww9Ym+1fr6
TJK+BRwFVqUOB22Euy614LXiZ/auBn5OO/pdMlA5UCriZO0BeOmArampAkgPYVSsqRz69sF6SDL6
Hiv2awAatN9Wpw1hZcber1hoasztYCbVnefHAi/Vzh7KI2DptpdY0Yk5RJU09i4CU7Gojje9QrIL
4Mx2jK7V1mho7qWvRt49PNY9kSeLfjVfMcM0skq5/VfpTvCcyOJzD8iivkH+8Fb/aiRfZsV8DwWO
tjUwSacgNSq1fe8sAK33mrV3YMuq0Q6FfGt/nmKCH4DntdZX/BTglQQbuEgeJ/H89p8dWngMoVwH
1uyiLE2Gg968/ftwXiWYFkXzO2rrSIE1qHR4gP5veog5l3aBz/OBHjVjayBcGoJwwR8ToIzZmrch
hgrxYTtmYzEwPeNAjKGQigSBfKwngmC4ahHyoDrbkfifbH9jvFJLgJM+SV3Pa7y7InpsLKr08KIY
m1bcAhj8jGOKoRRndZ9NKblLe/ljcBlqAN4Fjn1eUfVQSrSdnBGnLqcrJYlPFCDgXNTAvrW7OIcb
IUd8SVNc4LpmcHIIy9WMpRl2RHRTIltxvg7CKHIL8VHkDDTT3aS8aNwDgydmR1VBYIgwsd8IKBR0
4rC02LEh9v12i37MGwFaTygSNEcFAe0+aCpr0M5UcE/6knIkuucdJPj8PrPd1LBcMenMz5rv+g5x
WMkbFpR4hjvycKw/2C6FJ8t/DyNheFFAQjPguSlnVtvj3dfe2ZUGgs8TXfDB9qE9qBlbaeuNteQp
e5Fliz2dFM5sSPELIW4m9TGerpfZIeYeM0/ffV8R2eH491G55C0AB4ajSOtI2NRknCcBLh4Va2hQ
DBwRAcWixzX+DbNl+4S3Df4j/IAnYRrv0hNdBOKra96JKSi/X3R65al5UQX6ZihCW0Fl2pbstq8V
BAqy/5aL7oFepRj59SkNKaaYzlEv2yDqmQ1YTJfs5/bDYsnDhtxiDRjOVWPIIYqoN0CE/h1uml3X
fUD6xNNWr5rIPYCKoUDMNgSGAeVhyAe3f7gf+z4rgcPukDDdeBo+PHVKAzxGHo0lb8axO7TphDO8
02BG2Qc38QDbWcv+ZZQDKFax3HVU7Q2bQizA82HNQGTd1mQ7gRFN2cuZc7meANP+LonsZLnq+IWq
MO0YyVpO2QfTvDliRseIEBtyNXWA7PlNu2T/qW2G+nlvPmbVmFd/wqCJJFTB+uNDSLVetRYFh62w
WJpYgguSlJSt90N5OA7MTgvXFU4Htry3aZVpmx+szo3rAKwAkwUk+zS0RDcL7MMmud2RhC274jWk
GN8dpXm2JyzEAr3En2tVDhQbUhYOkMFzKVyKetmR6W8C5xatAmgjaSsBAtbJHP9uQODpUdTnt0D8
jQHzInebY4BQmymOiBIIJWOkaZMMjz8X25pRxLlk7qvalxz09XoirUll+Bi3UKQaiWbzAhq20Mr3
c/9TGdd/TzpXPZASvc1jgdw2Si6OD3Fvsqx9kuMkq0Cc98etzuOcRF5YswfKEP28zA6pulvO0BUG
rIv1FTM0uwGUAhYKw6WK9oan8sIQNQ2cuhsh7ZuzRc9Z8MkT/3IAnmdvZ4A3HlzZ9YeVi4eCdxDM
WszsM1Th1qkJ49AlVRrEl/940k0xhAHrBD7X1AECyQi9er/gouMrM1vdJ4561q8Cmw29hyuMoKGP
9AedsmXcyWvpxYkiWJLNNxFeYjjp2y8GHP0RYa43tbkYH5kdPkcSXoru9UYLnReA2ydWAI0KUhQr
UchujE0kFJXcXQV7aC9pL3pjI3I+ZAYFReEqA+y9877wS0mnYxJyGr4YsoPXoZR1n5SovlZNt9fb
ngudpQWxkYXruHh4+cl0o3oNjvGPkfi4R4dLsSF8Mwg3k/SQEmxNREYdbFmhybYzH1IbpkE9UdgT
VJ6UUu4VbVBKafmulF7ti//MlAosfh4Dt43CSBNjThnN5tjgnO0YThQH+WfKzieG0qa8hw7oivFB
L/FasNgx/0rlsfJm2QXow0w4j4xjUbWvs63DBz9hJeiObeggJYkVTfLi4uXsXrv5GuyLVh0qJFWw
FXU8LunYmukmQQ3eW5ZfpkSIJYQ1VuNtptI/ZJtguCcICVWFZIHozp2FAjqaF1OmlFrL0VaDveqL
u9qAzu7xRTOuHDUk+f+I7UJMb3YPAsolzNPmgU8Yij1951JCBh6/tUW45bsHfXtXHtrnyk4rr3t8
ELn2+HuroNX3UJZ5pQSUoOcOmH097S1/0WLUURe1Fxon6BcYCv8tYUIprX1Bqi6fUcMQRh0jOkiJ
hXfJNIxgJv2B0x+zcSNA+9YSCU7eoS3byhj+N2y6McqIUYv1tSReH6ul3Rf8SN3qE91vB9rU2exi
FkgAAlXs+m1yLSDNifDUj2M16GvxYQYbafHZb3nptxyJ5SFKmghojzVl89Kpb9x+EVnU6wXSlORu
EBP4X61lihCkem2psMcjLK8MArdMIIVPyE/dwCzbiXNSLxwA+JpMPvezpk09JU8BFfdSWAzFSTmo
Rdt/LYI5AZhGyO9CwYegj7JOwIC4mMuPilikCwrq/ONy8U3V5UaWl7eJ4paoA3iDESdwcjQ3TFI2
xXFQt5hkk8qMCAFLy0jsQ+1/XmCj6VKpvKySymTxpLweIdbCBb2hc6xUvkZGwOYqnmRNff20glf0
i/6uK2jbIyshzsstxWcRtGZmshHcTWIiq/a73rs7TUR6mVdubo+lC54oxNMwbsBl5x7kg13hgcn9
JwaY0AH4hAZ/PAKZj0kpgMckthBDP4tJog/fY/FzOZIPkukAOFCaun9PctQimiRgYBdCeLqYrktu
WU9RshdgKLYnoRULDfL4wqL1bmR5RibuKa+7ezZsxpYV8d9UAiAK0hsM7+BCTvP+G0Rie5LKXsOp
i8Xgjk3td36peoHhBQTK5hlivMOwNv3oglSpegT79npZnLJg7XBnxhwfQXQez3d2mkFOYyqA9kjJ
buCWb8/GcOHlMSuKuJJufH2h2GgF509OlrhPU8w15JSvc6B70k+kmZ+KjjwnzdMCnGocBEB4SXsy
jE+FBpIZhRnIkkaJ/P1tKcQ9MAWNwUrJAvaGdusBE/3/iyk1lArLPtABjYycFBzKF10EzN80uPEJ
59HAplrl0qOM2XotxYBtVKHeWFG/JJdPINUp8iLGHxD7vYSvV41NDoFw7uhPbE9KdeaRekx/9bvz
MzEG2V6opqxgDtW1sLmUb4AllSrQGKwNl5L9eudSMbbX1SVXL05xLK4TfDvM0TqJmkBnrMr7AOoV
DQHabcVqOiya9m5Qoh08U1ZDnotc4lEht7mgWOi91IZEZCPGpif8VFEWL+pLFtDjiyDvqNOBn34c
UdIhaJrGnD1yoHZk4eV99cLmcXO9aCTwoWUybuLPIwNPEVhDlR0wDcWiFB7TXfN52wJ84adUbO67
ljlbenywT2IFqsPSSJfDfcA/6b9qWgrRH0figpJ/jAt5YPIh2swsllFm3gNyS3Wh9k45d8iMX7qz
VYjQXlgimnEmn+w3Y9y2lPnofpKy8j+cKNa+LgZpvzvPhPodnH7Rb/PkKI6RzyJgUZl064OS9sRd
xk4edZtF8kQJGE0OGSZVMWN0BTqbDjiS8tCXLwywwkuCgIPkbB6+wz4Yju2vTB+d8mP23rFZhlc2
ocb/MmW7iqXS/thLn/O2oT2c+oxAPzFd3GAQe16ndiz63ra6aFc1UdwUoqZUjkDQVD3McD2p/4Um
yN5bIqxYS6LY+Ep4amEIYQG8MIsA0GCTF2lKT/JisnbE4eckIb/ynlIA/xX+8NEcyOIHoNvGm9sU
fTRS9k4YJg+bLErJwQ/dyWtsLG16384ffwtP7ylbgDt/0xF3TXy2WsiV82lrzCvjbPtpkSe/iaPL
NE5hAt9i1w8OxaSHrfGMt1lv5FJRT3BVe8gytL/hFBEAyw4yvTbwdiT1sBca90rhZLydPtzDHprc
gbuXNsU1HhxkQUYtmEHtReFe7D5diyzyd/05E6LDdfJw1FrUbu9PerIm8NuVzTF1hAe5gR2JAB31
EAGYBAzB+VKkZnAttbEh/qlZDiqs5flu0I6aLTuY0HqhGrUqPHXIfEXKa07uDAZ5Hq9UdUVJnVi8
5HGVghVClZc510p/QckU3+xlxvnRdKzvr8V2LbEXL84n4gyxTnzppADQhtXY+asCR+lPhEzwjfmb
P8nXmwg/RODIxyTtSODQGe4JX6766MaOFdrIxVwhqUFfvl2CqRmQvh59dIJqpTqs9DbJAwT7inHx
MkTMveGFL213gGDF5GmEyG/nlYk7R+vvjFGLch7kOKIuqoZ+vW9t9QzjxZmsxWbo+T3l649ZaZTP
58NA2qhuS9TqeJz26WdSGcjBH6goqgOg7rFhVQZXBfWBgGyJSNYUgzZLrxm4/2vrjvV2vtJsxrQZ
Bu69rI7qSm1dhqOwzEVBfzBhcERMSDjD2PmkxsrAd2QdvkHMpV/ktAbTWxB5BcAJy8QmvkMidRAE
6OlR1YGDwyq4uF6DkZUyiXhk/uSTgOe8UWtfHfagHcetO2s6UOFkJHAy0/+PAvFW2OwPcLKTiE4/
ljvHxznxbI04VwFAaYPyQ43kfICfzDF6+bY19VBvPh+cK453CeikVef2M0OWW8266RGEVr7xr7SK
QkQPDw+67RuePMyWvYLykBy5wnE6DWESCYEK0Q0f2CuVfSRbjqSSztM375L+Hil0NYBFZDaxb1ZB
o0hOkbeTKlGcmCouPanLZi2v8aw/M7AgjYTFVto3lbBrLMv1Cy/wzmEza/9tU7yBjypQnpFk3h/o
kzLRiX4JjQEgmBNFr5O7rvtK+6rtGrvOQP7lJPcNsut1ZtHRh/ZKZwRMuMh7bmDrpa/VLq/JvaLe
6vVSW2HOah/FudWwKXWVSSxuoyYv74951x090OUsc/8IkBOFW6ebj4MUdjv9jc+eJQ6vX/4T0oIh
QcafqyAW3GO/vEE+z10h0duOyOYQNGg+xVhsSWlqsGj1YLDaCQvUlGEwEpTloOh+aZ8GuxjyYi6l
EdWPkahKpCfm47lqYc9XvzbdNlPNkR/R+Gifa/5/sCPDi2HhH2fTP51A13nmUUdk3cHuwz5DSPFi
1dTBwGYMK6iDfg5meF3tF6wdyyoIyQKDgBOWU/roHTqxGy8fTz0bFbHVitT55zzQfrU0LY2bf5vJ
e5FmgnDOvO6kO5/4+WpTUIzAoun1U71gbfhaG/NyQorX34Qed4oNHi27ageg4Q4ljmsZdK+Yt/dM
QHOtgcVFti/l7I8TZeVwi1YgR9QMWZi4X+/5auCFK9QZWvYHRoDYTTXlniMO2ilue5VLlYV6BSiI
6eKgQD6JNNge3x63iFQPiLlGi1qzgxd3hGgdEsV4XS8xQdM/72UEzIoLy2SttIvJ+PTpBAMc0yoI
p5B7ZwBqehUXXeFj5KWEoIac4AZ/CYQP7Fxzdgwmveh1GiHeaIl02e2SATJ4AIRQzmDARbvXfUcq
MFneVFUtq6pj5BSYvDxgpqfGeKOIgHuh2Zun/TR8VDaIlLcjz9cceuCJM2TsNBaiKO+D010MzYWv
Mns2YY3NbFr4vAaZnYTVKQAJpjDmv4f/NMwm6TKfeNL4dzzqT3aHbNuLhc13tLwmAjs6DgACxMX0
OHvr8i/d80s2RgdqJUWMmosHkiKH/oh3QrxwRVKa95mzcwo7rwiwz7DDA/Q26V+iXgfdw5Io08L7
5k4Ih4Ejw5WlTMLJiV5lB+3TN+U3eg4m34Y/vvnYIDWbLeiLF+phU7nhsMrp3vwnbxzLre7UlDaK
gVP7Xu9G1/S7EznxZS8eat5ewDtKMWryPtOIDMCdhu9akpu8+LJ12LdTlwJC76VUnCsehx5iOZVz
9AFFUmGUlO5cyEvN+QzS+f7pDDwigIv9rb4A1BJFb4pyRRby/CSRroLKTX+3zbSBOSMCjcX6Bz0G
tCgzVIK8gxi2OKuC1kMrcB5eGIYpeYrZvZcWRvQKkkeJ/+wMJlEyPC727SgdkAWpU8nDuqBS1H2U
zqt0vQm395WzJHzhq9Nu8Pa3Kr+M6IiEurixl334EQwqCOJCSA5oNmp+B+SIbXqJWKl731mqpURV
ha3PxuEuZyy15ODZ1CY6NfCfMHW5fZkE/uu3Op21UC4BWjrlOVnJBZnO0t3X+VABM31tY8rG7SRZ
tsjYB+DvED9FhPMtahrrXAriKbdZMf/HqYQe+DQxG+3oWTLM0ui1i9KMhfOBMGnI8Fchzx693oTW
cZTixWn/dKEMXEfbB9wk2RDN4TqcYDKLc9DJnBL88/ISRWi/919/Kj6j3f/3pql5sX05FvIUVlta
g/l38T+eIbDGXDTSeNXBiivB+TRP3UT/8WPMHrPgLUHtsmx38cihJhRctcfJCHPQe4m+9BwiBEZe
FoU8Z4Ib21e9iXvmA3uGISej/wanDv8p3y2qVcFNmncGd6pEbxAYWdnficyW4TBUrgRQR0wcMQuA
6mU3KQyCHaZP7sn5IMiXu8SzkGqhnYBrYiMFVEfFWivBxRoERPL7e8enejlzEmL2XunLxJhn7yCC
LgqmALScZxMcp7A2MBHWSMWHYMWKwkhfsNLrouObicOXUWxdYl/to3FSoqFoC+nEK3QcMkP6dIPh
t4615e4mXoPCTjMwjmt8yjG1z/a51wJL7jg+x6VeoSz7F8DO37jcF2vSBoscBX+/gIfVIVtnAv0z
EdBe7esyRUxXeJBXgfsXwcHUgfzYTgqi2t3AYzn9Wxtvwtm9rKbuy8ekm1BTBovxakHW49L3LlyM
KDzbYjDNFytRRsxIlQSKtngGTcq+i2tf+bcI5eg95y75Am08k7W0qow49nBQZQbwTmYY0b1anaYg
jUZjHEh2McOlYTXO6c7yCnGANqrJgFIJXuygn0LD4r9hzV/k/trVPpG8aB7T0iaXy6qE6jaN0UGr
FoosdtfysDL+Js4pJP6zNnb9Vp1hLGIJyQG0V3L2SSfoJny4kyFXy8rySxT0LvwK4S/IeGP1vlPm
7Dero1HHNFDhZSRyP+GK7ZU5tiW13T7TZuehGVs3DC9N9Uld4RT+Lfi+LiWPuWu0ISF0i6Sg0Ly1
FlvcRT/VmKqRIlokiL1HsX3+uSwzX1XT48i0O3pd03ohFKQZcl7QLDuLC8t2TvKYxVZVsDUo/HVE
hBY7CKDXrywykZ0oXoT+vlK5dHkT250n7wpaP4Ib75f2xYMvClWtZW4nZX8b7OA9oir4FJ9RTK9x
hmnAdIukji76JBvWrxO572KEvi8lIoyeGBYX1FqcHSuNCHOdtf2jhP5BEhrrBNLCvzsFGUeIsC9A
+qAS/uVXbwSJKFGKof99LAggZEh39JW2/Mu4ArKVGM+W+NEyyIFfUCl2u7/Q5qPf3ZxyD/pPcFWM
SzvsujuCpXsc6VMvuKQesBFiqY7+RYBNb8pHDJApKu2p38eRx1OrUxgEGOqGOfQF7NJAn9oPv8Sx
aTd7/WGeXaySS2wWtFgtmdmmOAmwkUveZuQF/vsvFqKf32YEkb2wvuqe1cvsi7SxIbF0xiRiiBv6
+5FEdVYBBIAANJFxLNjqhEQZGYEu9z4pr/Lbm9u9hJ1qsA+0iJhCc+ulWP0ZMZsNLSTb29FFphFR
/4EXtyu/60RibFVdk4m/HyO6r+/s9FLoX8t2P+5qFEmSsv+2F6WxDOGxQYPtNoSciVVT1hjsy3Iu
Mx3zsKPTegkj5nOzhUvwvmFVDBlEF15znL6PUPEtS7fS+Vbb967I+ZcOe3Ioy7YoOuTxPFHEY+pP
etFIrHyRlqAxR5fp/WH7skUkw+/Q8c0QvVyj7B4FNNHVcJ6ORVxkMRrLJMGhsvdDHzZT1bk0pujO
NCCZ0xMk8TYQWEy0nPN+3CTiCFCI99PsHBXx2oKdr6SmcYTBuyBBCSzH4kyVJWtSilIVmjC4Ch0A
8cCDytUV9o1Px1doqjlFXhWIIm+6rwSFcGwFH1GbfLX1r/2c3AFyfgE6flqJGTVrJSP1DUXFT58F
KZWGGFPOmln4eRvRobikHJvU/spadMUWRslAYjeircNZVR8mJSsmMVKYceqbejb3muAXzCdiLpER
hC25RfIfoodfv3QU9b39PdDkdaAjzU2PiW2lj8dpYX0e5lFSJK6jvooZn86jsPJsfohaXKQMDdRt
uYDgcQn7N380WvB1XiWsqz5BkdMfN49G+unHBqPXbiShXqspluuFyqG+vWCyLJVwRc5E+qBDO2dt
Rzpbs7M3rAt85w3VKU0WLD7HYKY2T5fsQXBk197jYI2vFhpnOYlqElRy5g/feQoFzEm0+ZcJukFB
lUTWzAcSuDR6k5BdFt8gnxQ6ZqX1x2ynjBXPiBWM89dsNEuIA2FNsHbKeIaiV4W6r0A5kBtO1rwN
R7KB+pZFhOlaTOmlaWObX38MlMDaO607d4RiMJ2x/KjlGAwKVc8lnMttn6ZyGl7tW+D7Oecc7+za
r8rkDZ1YV8KElAlgggOvfW9Z9yAjHeNIYX7/eswHxw3NsW6sE6CJh17Rw7s3VRRjwT4gdF/SABNl
zpQF5LJrupVyc1+Z9NwfWyR4u+o6NJRhPD5QbgbXi1tpiJTQ3XeDTI4xLdJDbH6nq734t4cz8v7m
Vyu3CHIOIw/VzW26XPcpBrT6ItO06daRnS2L4ORmZY19/7t7Q03wImSwbVahq0rrhAsicD/YPdMX
YBze+IKUMk1WganOsoGhe0WZHcyyrKtgc17mzxJYl9HPXSFAhH3B8B20SNZYzHnfv1QYUdar6+9B
fC1f6MUePyBJvnwE5y8Y1yX3UiBdl7TyayRVA3/68Alv/Vb+Q4C8OA94dMOeOcXpJ3aV+z4bKKhb
35m8eIRxhQ8GBHSgcKrpY+4DlqCvTmhppqRNnb/skvI3h9Fsa7+w1c1rPxzOwaIy5vLP1z5EMQ0v
qexP+aUwIrSH3jI+2PlWmJo9pJJLLZs7qGkvCw2v69hdzpW54vQTGZchrurkJMfJMoxOPGU6GM38
cY7WhJ5tc4xm1pjhAfWGiprM5fzep1QITmrXmw8RdLGZaXn3A+iP9V1vwenEpaQk37C4wD6xjyma
5SvL/x5jVWxHl0Nd/KEIYLTO+0tNkVCT7zPDDaj6y+g62xThhFe8YzsSHWO4PTtgk2uMyNHkPohT
5wH4s/pSmWH4Cam32UhjnCb5M5CMAadOosfMAh9LNjH3hq3zcZ0+V5oNZeuqUoi+eYMMgYh2yvFQ
0Lpn2dCYDz5K3Bv1fjPuTinNlKATg2L2MUw1zy6T+Yq5+X+mGputu4/5L4bELtLOpAHFcsOMQo48
t9m6EVBN/5yKaofOhvPlSPYF8x7qdBLzKDELuLaCXl8dMndSs2xkLJO7PQg611Ki+A/r2FR0uNKS
Y3wb7gzNN5yGOYQoCIfZULAxIR/o0RwLTmNFS54Wlvqs7ndb1KWdrK8AeqB/deA7/9hmbFi/ZS2z
x8aBC2DubAhlSWMQe1agXrIDwF6skbwb9ZFadg5B+aoiARwu+WjdFPB/Hfjivi5O4KopHO0DmHFs
7vTCQhJjcuCo+jYqNgtaLZri8grLokGUa7h3V0efb8ov7u1tQhdf/RfYYgvjtkuXoA0MsJkIYdZD
ZSIm25V+OTbhncSCrh9N6qbncjeQNtDOPA8t3mwA/wj7vQE7qAAyc3Jxbcf/Uph4ugzMdkmlSSLP
JkTN6n0XLOyBr4zdbmmiX0c3BHWjE6svXz/vrV4AD/lDKXu1IoEU7rz50H3MXv7pldYF1S8mf4jc
Ug8FPpNZKe5mcXssDsNLIpCxOsWRCo/OnOOR6kvZXwU3Q61c9QvmRWMkoXT1tgMqE7jPuLuZtSUa
Us6Ibo7hbhtV6j6YJcUs+SSq6Hei0GjsxA5+/HjYJwW7Hwz8cws0OOnPU6sNsvAx/ERmHIrd5vkP
1+B5/fXgmmtqTcWbZxuvfmaLM0vLaBy+KyPdMq6FIJvclEkYCM1yOnQAICzMxjq6knxdoXtufAzf
Q1g4o6JJmEbVu6Wl0y9gFzdCRe31imV82h4Op/CVUXF1QdT1/4vSdWakktcMk0yjqhCNOv0tigSD
x+5y2PawWUntVBqsWadIIonTj2x1gNocZZir7ATn9I8VRJL/+gh2xdz71VQTHrOXDjF6EjHyleoP
3/fBXtiWbBLHC7T59qIEkWW3K1ozkQ+OAUJQvMxKzRdd8p85hQR83Pc4bZcO3O1HusYzWIHAdBY8
VfpMsUKEjNZZMbn9JFmnUUjoPCqZOp2KJtRqEng77vaC/2YaINOt/niHAb6rjjFsLwcV2+jiwO+W
Gg3ASt8YiOibLejqTKbBOt/5q48oxUb/XBO4Fji2omeQoVh/T6vBqEkK08xbYRIKhpRoMiy4NLd5
KpCUGveAfzsHT4hQoRSX5XWFfFHzBISMSX2kit8NfeUlKjIVkydVXOHgZ2MktiqDV94kyMkzSo3S
h7WPaxaXSmuK1jpU7xYg8i1hppI4DzTbaFNHdrpj6lXxnpbHqBtqbvSCOjGhXbiy6v+AB96rLSaR
4AjtgwS+HbFh88E+QO9EPHcV95I7px7wKQ4p/UXwtWGCxUcdKyl8aYDQZOQqbnQ6TAQOjEwXa80s
HjHTr4NA9IjfUs+2c1htZkEMv3OasAii9KqgAOsHt/EGbsQd6CIwWdlejCmlcb3MEp8Q8l0uVISj
7lOo8ca/2j8DNrkXdTGJZuxr8M0Jr19h27HfApab4YjJQXFrLofifRZYj6jJ5dgahxzAdNtBlI8o
xOcc3YNCh0pzVI8OQV/Dvgzz9z8Y4ip8DSX7Bo4Pn33Gs0kNkbtDjwWIq9rW0jvrIJT34AxqfLlr
QQEFkmO5tCXEwBRK4KCqn77tNfRWp1PyllQwjz1DiDfqWYdN0/yZSnxADMteh8eFnL1HwPze7870
N7wLVVUQXD0pcZfVozJ9GzJGpkziHlokfbIP2AH8nG1O6ztmRj1r7oORb5xnkqngHSusZOyIGE09
ZRtyD5IaIZaP9jdy+pcrVrmilp5DRFHY/GVbiG4+8yBYFU4qES8iGlPKDgu74dHW60wXyguvy/8k
1UZcE4GAqTGW20qxn8DkAxq1k7b4UbgThv1aW5A/Lop7xDkE+SekERC2c8hi03SHUPVi45RcuXTY
f44hdK5bdqXpYaDDQ4ibSu7jBkM0Kkum39LxM5xw/U+288VfDHIoje5ckqlfyDcl3yDk0S763D40
clhpWqGHPTMySD4WT2egCYLxd1UZLN+nBMHcjLtwUTNl5OgkCcmZKMGJLt7J82enfXu0ofFfhKHS
ngmsZsRHTAGp1H6U0+B97dojxWKGeBXfSii2L98EHLz8s8FyO/xHXwaOmaiu3HrN8X7yEbmToeUW
zF6oab/bL98v6R+fp80XmOGaDAfR4xm1CdUa01Bqjt3XjMVjxN5Z9aziMZmbvFDkJccUdXNoCnZI
cncW14c0xfYFlWZosbkxLeArOXeX9au/Kv0PiUZJDtxu7UPJJzKiZqRc/zwHYAtBP0HLxVKg2LNz
kwjmGvCFkOMSO+D1vmmA39hXvp/N11MiG3Rehy3I7vOA5fd8TUD9C+MO1jBUa6PjuJqN1MWRg1+v
XqWeeMCQ1eLBx5SB86ohOoBlPa15vdG6ZjqpKsZ8WtaEGBTF9TQIqGS9SErTYYE5cJx9SryXWwmL
ANe/jpNJs3if31DYXt47sf7oRm2gPhrd3hhS3y9pUbqre9lNl/sNFgd3kOQe7TlLejJJD7EETS4G
rgHotYTNIKNDnT5RXux5CUK6wpi34FW7Zc4RYfoUaRCoUjZgAGHLEqPwihFlQgUhKb3Dv4i+vJdb
i1lpqVGdkqITmHofHBixzMKaxYELizeXch/J9ssgXKSOHXxI5Zs1MdlLvl2ESOdFddZAV/nxJZFO
KclhWbSDI7n9R4Z9WM5+0MZ8ypzt2dhDtXOIoJ4l6nLjUa/ur5lOnFev8OPTDwvahFC5Wgpb6Oi0
Iskw/z4/qh4FBiw19lahR06WAQcMeChOsaTPCNixiq18Y5xyRwZBLvKaatY8P0wSdQryDSf1/zdQ
IvDTo45eo7Y/E1GjKza8aAw2o+Qcb4ApYWQFI7Uh7pycRw1NLmYE+wpO4Rmia6ZBkw18wS2jhzFU
L4ETJiDvGblu/z5jkzm4X8DtFgc72O0BGLV/0nw2yJtabJUeml+cv/i3JHufwdh5GJCi3CN0JSce
5ksI5pV/xN1JgXptwR9IgV2CC6YMmoK5dT8yBM0GlCyMBqSMnrBXZwpoV6Gd3fFRW1XFuzLnalgf
zs6iFyrDkMOCr2PVcyjXNqkcZMXtdnta5cbJWE7oIAU5YStB2tUmjgXdPv76VVCPFjihED98P1Wx
KXV21RyDyByWjSAG+iy5wJLtVVlYhSaf+3iRCLtnHDO58hgJvURnMRywKOAxqT7vAiPjrNJBQjo1
uv93URlpuouRaLG8LJgtJYQjSsmdVIngzP11w0HlBa03X8XTJ589bOKU8TAXcQc8tJ+06sRYGw9x
5z7AmeKYl/wXc8Yqumd4yplIpLP5KsWBgk5yGVI13zecXvpUfGDy3DxrmdsnXBQRNaaszDf06sP5
FPmYzi2/R7L768PChgSz7kGZMcsOvFyTSKJui5aO4t1ppca+6seRiNFoaFPxEgPsGlqF14Nitw7/
nBf7Pyt2JVzzQYg3Eo98lCX7DHw3HzkNbuuaDL0tYBv7+FrU6jYEJ1/WoGEccKcCQsN7GvUzsawG
3yM1astrJPyftxN1io2jA+LRyxXQGA2Gx/mXKDNRaoWgAdRIrC2EAaSFv2aWE5nyNNy2StvuLiVT
55TvOR5yn3+9jQcAuAqAGuI57aH+cOLDXEHo+ocysYlkHxJvvRB9ncM9SKzAk4E/6YAK0x7CLqOj
ChQVYF1wx5ag/ftycMjc9LvYkfn8uKEW5wgrQS9r0eALifxmxmLDUhn0ASTrhBf7sYdETOTfPZQg
ReyXHjfrbUDsww1Q2xhz9G75dM1gx6anveMSaHuKrD0+5vZmAyioCUI3cUi5ik8nNg4SAAu5u3RE
9YdjN1MWLjGE0gdrMwMDa7j6kdnvbkR6d3XPDHqbVXFK3UYcFkAa0LBEi56nVmIuLPKxcYItBHGC
TvhIxnvQQNckmYw93JnouHG+og49MXhJQJeiOurVvxVp/Zco9pGoFUEFCeOLBd2RJpadA45KN/et
6Nry2ojTE9dEI4xoaRyGozYeE2rTearrsSFxCYGqBfvzUA7yF+EKFo0SqD5DWBbQlJg6Me/4V10/
aH6fcSMw7ZT6RwxQb3/rAJNGcgfclzqQ/eE6/FCixKrfZCDkAjM90XrP5pc+sLTDcju4CIB1YaoP
Jbh7s9fqzI5Cnj1Nqa8mcio0QYU2Z0NVEQabohH4sWd5dLwrERTWvfsMFoFHzeY1IVDaWcycipfY
WDdDXMTwG4NqJxv1Bd38nuPSEA0kWINFvSNf6sG23hwBGk/kDdZlnJcPlux3CmMZC0ZWPf01BCcr
SgMQO4rczudN97aGSlCZxsE9xT2+8sNJtVi2TrFgQrMfbdTkpIAdwIPQdNsNTJTsR5T/2/2kDM36
MtSwmMCPn7z2sIrjRewCwSUQjgQyfIwv4TvEdK/0FouSuZE7Ng3OUvpnKhn8QBMR9ieS9NutQyGy
m4Rf+m2/L8elsGzUhuLDDMW00ylIaeqOENln5fyK3hvIOvEy9YyxorfRAAuObbVKruevyYhI6bpV
+PrB7XIqpbiRfQuy970Oh3a+MniaCwE6AHbgMThll7dE9wi+Ws7HtA6H4F9pdZ0T8HeRbahPzKOO
ajYmG6yaS9ooiwVi4dj2wt+xX1J5J5zwNdJgkDBJjUyWd0E2ywGEXZxXgwULa9EGEuNYpvhj7Vu3
QNPE3QGE2qwZhUH1UF3KZUtcEy/4P9oBaYWvdt4AODMCX9SbKXWRzyqxr0vBzrzKQyrbkf8L/CIv
y1H2jGkOZ4oRiqlugH81XuppfZdqIe8VzrRclu6PNVRiG+/SF2nsYk47X6GWKwlHneXlTBaTKqUe
BPLtt5NPOEZxccsyLCuX1NDTHIYFTzsnvtBMAVDqH69B66zT6hE9lkB1TEOfn/noL01SBIBm4S1j
DjZA8RbOD249udAknb/EAUvkDoWooxwYDMifYW0YMktc+0BzJTQEhdlOn5YEK8afad9sw9jrkgqs
azXWj4lMUXhd2f5ddpJxv2USdSmRlZBKrDmqMVd83Z+g4/b3jlo+4pC3/T26/a2AntItKIoZSn6U
X5ffjp0HvtnANHvjF9U08MT7J2Icr7k6FTt0ca7VGyenlnODaG4ESmU+6CttLvxHz87Y7P31chqd
gp7TzYOWNwlJjuRsyi0lMLNRcHjoq8NCKpJYWwxItaLA+F42+wby3oPyO+2e78v+A1KcqbX57LL/
gKBjnpQ24LUNLNGAxwSASVqnhTBE7b08VGaLWVz8jULnKuz1S2Pv30ALA9swxgfo6hdpP9fo8ZzC
2j/nd79K5LWQMedFr9a8ugJP9IcrQFpsP5MNhtjdYK59qx4CGOeJiwSFHLJz7IV60R+zU3DlKqrg
AK2bnlHk6tfVVH6l6b5ZwEI9mqEprqw1/7+QMT8iz+RqS4eLZkKNu7eHyoVMlDXA/nFPro2G8Cls
wk2EIOfj93/ayR5WZkm8zmYad3qubEWfIaUyxG5XAce3HITGj+ddYwGFINP6L19GZXNlzrbzI4I+
deFcseDSJsirT594iu0YChyuKSvaKHjQn1VsE9pdWUqX8Nm891+/aKs7DzchC3FGUprlGPUPLzgw
GQvkTvAqx48/XUZwi0c72vZcwYZdcLF6KHVymlhLfcqyTlJunp3v2VZgVA/btmkjlM+I9VqW1t4s
rJl6KiICZIqkz2H900s8wwGLtNnCsVl4PFQO9Or8sWZzHtVCB/7v+Qmra/4kn5nDN58jxxuIeHmM
uMiQa+2nL2+i6onBMgmNOsX/e2gv8Ex3URs1QfzpdwKZ8DMItHvrmfidbxthN3hRM4PkPccvozWj
0v4B+L/cbGks5n97wQckdXRi4XfhuPq5Yj9ehV4krB+d8JpSX2aYWuJOEGK9WY/Q7V5X5BHEKVKs
fDUjMRGeVRJYEybR52jO8HLbNkyc+wK8p5cxKnVafiKC6B8KL+3sn4NGwm5Dm1jUeuu2nlvUufBP
3kBdi/BUTdlQgb4Yb1nkWbPdaZprYuSVjOxeeVNHongKfrC0R5vRTatWJ45wOMqiKcHeUweIhCLW
J4kXqLEuGfW1pB7EKpho90lNQFVEn2G5R1XvAya2lOhTYoii/unWfsANwLjfenlpVYoS7UjBkpUX
vH+j1rKkRE30qpt6EKK4VI0iJYJAi6TW8QT1BYZGGtpeLd0SoZO7QEwk5jNHBV2aXUu2o9W8LxrQ
i/bx0cgA6MBAF4EshydbyZmY9O6sWtKB3onkoZc6G++yhBAXsJ13kAC00gBwlprYE5sY6W47feDe
WiEHYx/75vvne62tu8AYZ8wLlDX6rXlgT/jlQt3zooQdygo8MytNIAKzt7RCgjxUffdJmoSWrFqJ
6h/mNgc4OpRjutcTcTGAjepBOKMDDKfd0+R+zio+r73o9HyQCA2V0HsIi2/Wdiy3gjD5eO8eeH23
r44jJYOV3zlLrFfwUYlheeyJr+jqSp6VjCEg3aM5P6A73AC0yMrp6LW/WQO26AxhRcwkuGKbhQ7a
BBBQnGPqHy4YnE7WABLA34zK0SASExCEUz6mRBxliHjBTotN9A2RIN/aPWaFynzYNcoZt0tNqUOP
JKhCFSurVZdLZp1htgR6ZbjKvvrXSeAEe/mMJmGSSvtgV0NA7Sh7Do5xIyQY4r2zaHTpwtQIsdxN
nUSXOfumn5Z9YBT3wkcp2X0Em0cn16mj1dylM5NBLkYtIbmUQ0L/A5VCMA2QFVlhX6KastNwAw32
4okhllgs0aZIpLXsBsg8SsENDwaKzCS7oejKW07JAebda5jRrsC5JXewexC2By3lpLeodrgxUAxf
K9AM8OpqpHKtHxrsdkc/hpw39/sKti2MMbSRG3kwmU7hmioSxtlAH/4cvxPsZ+YAt3epBqx7MJIS
rpDnWr+1sDg0gDIbaG/sMqvDxDPJ9njlXC/C+qMrs6rltsrV/6EIqq+1D0xrx1j0N8xQsBJ+Qwan
l7sGgzU7qdrHjePODn7nbxRvItq5JA7yGxPciGAz6XuX1epiVfoNidrN3i+v80msOJlxcaTEM7WP
4VOnJoVW57yahQr0L9W7F7bNZHo1THEaLlqT6GF6dPF/+f3mhgsHlgrW4g5dx/kyG4DThQJq/6hT
NlZS0UGMBKKfkJ1QL97mgWzBtwOis3+aNh0ESt5eBsASJk474SM19UxUfM1kkPT6uUT0FUqu+GT2
g8hhZfcbCY+DKrbLeeNc6oQi4XUAYtimFWe71VeELF7V+0i6djzPmsV1Mujz0SDn3jQrTT7Dkubh
LOc25uqYD4epJAcrNMjKGWmy+ZFrnW9R+e8rAATWgZUIfYpPsz9yET/3dKoGNuBHWaKTCz3UQX08
wtMo1vcfjW+VA7u2jSkMSeoyQCUj3HEeHZXxvlyMxDccBsQwpP6Vz48h8FFaUCS1XP/P/ceRVi3/
W4RT26AE9DkezQIQPObVplz+C3T1gu7vwwpxOBiq/rVOhwAKkKGHBxAkXDkrDATsC+daHZ/C0Sha
KeRYdiRQ9sV1bNFQgLuutKsj+OVaCT2D/KXmAByjbRLAUAfPBArDQVIzZgcMHDSDnYWtxmrf5TVr
iOP+625o2SaceBPWMCs7mvHA6qtUJHA/F3+dCe9bpUiDae2ib2WeXcofM2B7I1b/oROAmo4Uph6j
L7ZV3f03zbzzgZJUi4KB3X6EY2v1AoKMZ0tR3ZIHYpA4jYLAXfAltkqAp39CmT3pnIPyCbLlY+/v
UaD2NCqpeRMXKrHU4Ts+z1boziDjpS+77SNzzwsKe2Mez/D8MgSZXbHUEwr6CSXs43P47yxpR7jo
VgOiX9S3y2Ffzh9sDlzpBMcDXU3qH0kkyNihe9HsTT95Oi716tSSvX69N4YDB6dGlGAA79ElGt6d
rcDAosFmH9TYqjmhRPgCuzvulqGXeLxwv45johMzYsMR6WU3D/0aCZx9Er2Zrb+Y6NSZXQri/uFT
dSCLyWtZXwoCCQMKnQh1jHhfqr0NsVzTijLPM0bwAUvKU5sTG7Y22QZnG9og3iozth4za768QDMd
0drT84n60AvQdvm6oO9IbIyWQliIVXJTsh4eWrJXDllHzXJ3KRwlRMRgyutxoayOADI1XUbDYuMD
jiRLMtIdyTqC2X1SVu8Gnk88K3VHXUzGDERdu1jO3iLMd1TmAwMXUha9beR0Q9aAE5gh1LMe49W1
3D5qmIPOA+deb5ZnLa6yOwnjjoGKS6qO50QIB8o8W+58ljob8Hjs3P+PTvKS1iGhGPb4/kTf1JoA
DwZexIyO3oAskGLvj3cEHTDts3oL9xOiOKE3LZbWH+g/xTVZr+vwFrQabBGwqGJvbF2CkkoJ8W7f
CDo5w1ZmQXVUvtgsNfVlYd6YYKHO9bGjUjMOMaeCXEGzlJluJoPHozi4ef+mr5vgomcS2Xlt1a+c
tPPCDhoH2T9QSVXS/q7VpY4uJoBajXOiOw/yOqnfe0g3xA6EMhp3qiKH7FAtpQyLphsXn6idEWjV
K2sqBFEdLCW9vQzVJcxlzRE39q0K95k1/asmRUf+x2GDKgTrQQt2kzXbAEPXnWF5KDzETYt2Ht8G
ZXUQ1C3bxXzlaM9hp7qkr8bd12UiVzSpAwoEx9aD8oAA/LlVo9fL/6jkL0iM1Hm3OyOYSTWoEdNR
ADEpN2XR+kXsHwN+Zg/zwo6C4RbaTbIepXXKeG68J6zgn0fpBYUhRikl0LuMQhoRSyuWuWKcA3mC
SRw+Pap+Cxnxpwn1B3y+0/Beihk3hMVvSe+ibEDBX0gvrKaRdxDOeU8atyJqny8A1OcySBI4FmPE
dEyOl7bFdU32I5RvRRDINl+HwmE4AWs6mTlEU1OOt3xM0h+0LlSsA7o9sK7E/IGJytK9kavmNW05
QvNNfCRPr4mgcO7cxQGaIN+81M1GLce2WpSPN84Oya7Se1XiH/XSTWSR8oLnFo5siCeV4ll8Mc6N
NTKxe1e14SYEcW3DPZ1855TVGL/pLe3pHEImYrrYUMO3NN7gQIGRBqH6mnFwaoTrXdDLR+OM0Tbq
JXVQKepkiRG2EvxCvPGqz008GeSlhapCzASfRG8eRVKTbSaBXFJ1ZubgXLyTp9FhFPs6BmXhhybY
LfkS3gMlH6Aq8yb33R2RuiII3NQpq25dk+H0p42d38TTmgsJZQXZ63UEEHMMXFTK5DTwR+WIit0N
C65XSpTqPaajLXYmS1yxIEQrS938onR29I46i4F9az6RiGSiB/gT4kRpTjWHOVs+WJPsBc6sAHML
fRWqxpeKf7kaKBEysT89fQaQyIQOLGEUadV5z4V69yWlzBMEhxU80kI9KtdioNkU+eq1HKay2TfY
C6C7zWTSlF1q93po/sTtaT6MJHWktpPKTzf9kTrvQW7SQfJ1NEwhZ15jF5tOmTq5HouKFXN/aalT
DQ0QRBR8x0w/1Suoq7N+3rXduPrt4jPA09dspGyx+PZETOvkARv3EXYuuRIoilIOJHy/9xhZ+tX0
xquB+AoXw2ETyItb+NYSA08eBaCFLTq1SKt7eCOlZQUMIO2gmxvVa393SN92Zix5cphpYKY/zZvD
OJvJq2GODFHqHP4Y1jgREnNfVLOhOOGVVcQRaY4ty8b4V76aG9EClrh3evCmZHbG6vDft2NPJ3XF
faM4zkey4Ws1pEe871NeaacWCGtsc4OGmQHam0GfYPLkDstweUIqe0ShVql9SCaY/B1Ts/cvaygj
31foPZZ6iom9XHPkzc/WUrp+UoFWX30XVTUWPK4y1pkulIa5PDtRzeRCg/j3oxcZAy7M4X1Xf8Z8
dlzwtvLqtklBAgqcxY6iT9COMHtZBPXBjfyiB1sCcFmooBZid2GmwCTCzXA4ghq79EE8Uktk9B+/
kKSCq36qktkWhikEHhv3kkCwMogjWhLw1KHyiJW1mk3x8UMka8QU9qz+cOeSdh9QtpM4/cZidoA2
fquL1Y8YUiaUlf9SO51fZTjSHswFiELQUEhePV/G1+ijxrTKEiA/3kNaVIElgk5GDqK2LPXGMA1p
1OPNw+SmGdDpHnJGydHD9eSSMc3q6OUqa0T246XZItPa2ibOSCzs8hI4rlHuUKHwQW4kchfAdI5D
4uaG7V83JgRki3w3IgsY0eE5AENcaO8qUlwsyhYkdyq0jxD+GHK3Ycw3eiA+cNUALzeXOj7B8jjC
COx/cfFX3KgfbRc25TWQP+3CG6rW+as9Xe+PyLkLhltDpYVrwpW5lWrNzYuBK+voOfnbrzfhi5mR
k7ef+CsBnqgi2WZBQYpmi4vvUM8gXD71em9JUw6YITld3lCXDyXav63Ymuq5UbruubalKA8+kDF+
zx9afVABeA+p2E6VlBS9wMvt+N1t/Gad2npXmggBNbnCMVWLFcZhEdNqmQXxup/HUFKX1ha2EkO7
Cvg/P0Y9FwNeHG5zwwl6Rw1/7Faa1F4LDpPFprxPatK8l3bUIkukcRt5XBOmE1nJhEC1/lWbznVv
fTiX+OvVcrn8krRU8pBIfQCH53cegb+fgAdJSRfgYjlxnukPmCD7c/OZPLHO6llBvwNFav+h2Ya6
w924Zeju8NdBkgdZsx1pW+a+NE4GLCqGri+RIhxbr4aXNhdFf+AdxYTzIz6roALqosDKCHkA3Dkl
hjLcv5fi5RxOpbJC5N1o3FiFCoMtfoMvEir718RX+njfEXdgnGMZm5QTXU79RkZFVK2UnFY9gMxQ
duvqvo+B/8SPqFCgEZc1mDkO9obf2/za3EOjY/FVmWS0djisMFbs6MPSJrFNZY9kpJK2lifiIwtD
YJJLwjXOgwVGnMHOQz51md8POMOvtiC0oqSt9Og/h9OMSEzJ8/F4VV7VTmVTKMZQt28KJ8dYKgCF
YNf8sTF2wTRXgOdPl2SUntHTUkJ6ddPezSEU9N/2tE6OAlrDPTrxkh+X8t6v0xS1zfQpq55ls0Xe
m4lOcpHG104wDUHRkCSo6q8FVmyk0pTCFK7rqn4Exi3uHu+dCy+EuQmVcXEAF167sMnJub+PgQov
/n22upgmQw/7D3NE6Bw8Ma0V4Ujc9onRVStmnPnsRLeWEvaAAb5cmpzfIbivZuJd7gfJBMuiHL+v
AKtsr8o0A8IEjiJIg8G7lCMYAgbhjoqB0qq80azI9PQMBbtADGPOdtRxHnF2jIhi9OR1Dx/zT01u
8xMocc0ZvCqPUyEMGzejLPWmPx0brYwI7+jBo/qHW0grovkWMAbKRTz94rNVYPCrUu7e5gqcM372
haBfwnScZgHckwTrRgMQLTwPBmjjvOirsSlmUxE7Doj6M6FCp4rR0hK/9r+zW4KEDIuGPOt1/+Mr
v/PKkM/eX5+9O0N7UlOR7KnsXRay/gAEK2p8lhooCSkcpbxJF3vNj48R/2Fn3jybHg5fWZIq7NRf
B+enFMXm1sJ+QRqVh+mXRlnoTO5B2oI5dkT2I+JjNZGMi8UkdPI7gucYEgLre+K93EDwPn4SJy9G
FceKAbqfphbQii+++gpbweTrhs/xKOcai0YTTE5KdNpIHfjIczFrB8XNlMC74HoLoGyxlVie/Ws+
aS1ROQbkEN2Avtn9Y0Vo2LszLEg/Uh0FwDKQwKYW8hlHyVqIVD0vH0BdE4UlZjnstjfYGZUKKckg
o9LXpshH2dSbHGfHzNkU6NNfCH1FC7i2+eVVSWEKd+zBneTvpbCH5wm1WCGVxp7zSN0qSkCCP+14
bUiMF+IU9czbjeOfGWKkEsaGl0mYOnuvcf9oMg04MbVAj0Cee42BpWjzrfCv9rH+c/IaIpca0FnT
K00Iy1+KMvPjlbR55jmUQ1tJyaAIH9DF10/2zP+523abQBfhQF37sWNCVO5dia35yk+rnbWxmWyD
NK+iLGcOLzbIUJtDjelsaVav+EAkjbCVq+xWRv90cOSCWMqrqhKiyrdkQNelLMhIUWD0g5bm5JHM
ECSZPeqagAH4s9TU5CRkiHBkdDzZpk/qJaT+8iWqblMtp6R1sYEGW0UyHHVNu9O3lCFThsS+NNCI
lv7NS3HLjk46h2ZOp6sWrFNp06BfGb5HGgWLCUtxCwsd7PMk1FmK4wTCcdrC2Fdfbk3skr6elgBG
h3LS1qvdD+GIXKjS7EWTVkkLqLLxlpQbplr+XUBGZQlrGQI73z/Fa+sreHIKv1tbAas74CtU6261
hLt2mLQG71AVXXFwuXj0QX2j90bhKGwHE4wmCtmzFdrjE0TNGalvULAS1T//HMWWOhtkVj4qzErf
Y72Iqu3Vs7yITTyZzGs0i50K4h66P9Opot+1uqWiFDdbmZrpnQb949gBtJMO0q/S5xXuf6WgBvf3
51zdtjsNPv3HCVBJuU9dZXe+W6o8NNXksGix6vU3ejCXIK1yxqhnfB3f+MPrlFswQYiGft9KHx2x
hHDiyHCFilHpOuglFPcliGTZaa6fT4VgB3swnDeEZKDwNJfKLq9XtJrazVq8Khm28DMZg/6Z+Dfy
Y32ce/pKoZmKtiZjnl8ptNNvr07seSPVGGS2VVRIqVOJNEYuyjkxACQqaomjszAqVxVndSEXb14h
UUDNerpqJ5NFr5EXC1eWdpU6PQSuRTSI7T3yPi4lJ1Q4V5ZVWNrjJwg9t28y6qwK/BK/lTaClfyb
GeP2EjErzKwxTr/Rbeyem4cdGjhDUuPZBAHSt/SQGJpgnaeRHbHmnUaYZ1mHiIPuGEkwXaBcOcM5
Wxdu/46fu3dRNo1x6NvOuop6rVuaIyrnBu1eJrHpsdPCf/IzH06GvgnKHBlsL55R8I4BgZlx4NZI
p6maM1mBypydy67g0w75zLvlBbatWe4J319Lvt2l6AxOmYShHDAsmTvosS1ncE1EQf0t8LOSrHns
uSUkELLcL6Nz04y273yKqQXs8yL/fRE25z0gegh8dDr3dcxuH9KwwQmEw1JhXfNdnnpC0UYRqADc
nAcJbd63MCS1vTENe5UXP232/q679ElzK5/g6KhW68U25cggNmJE3ifsHsaEem9CAq5JozLQPyVr
qGiMNvSVxWEMwO2PirLYGqJME9T+dTN03kgU0Czkjmil5Bm+exdlbL0VqFhjBZ6n68e1MVmQLqSI
wGDNDEw+Kmz/IgPemciUHvcHm7fWWu113+BOhsh0fn9fu10ndTULYpdhUJ18aS+fTPtAIUQpIc+T
6x99Ywb9F63D4WzEYNcJV1lGphW12xI/KqnDMipblW/EOC1WbaSgzOs2wAG+2+ZxcfOpYNrwpF1j
V8GHAQBP0LZhcS2iYOqN8A9LEwkbf+v24mPhTaRkDhG/WWlXWI4xYGiBphoufaHUZa94AP6NHqVh
CqI941iYpB3i9DVwI2ASZMHXlzRTDA9TxpdBnxinIFgmn4v58ITQEWquWmILX7wQOnR32DVe5It/
4mwQBxYG+/6VnQCWBiNKMB2mHi6b95v8ARcp2q54wXdkC9mxBduz0Ka+f6qMvEBxVBHWhsP7S6NK
2ox8hWDM2oFlwf9DeIoIyJG0+KbpQqUOAjWj1QYtN/o7sUpbSb29RAccQtjgN+unUJo8ZcFA1gV2
DjPhjYD/jxhwu5ZY3RNfAGTpv9E0z/pyh35wPMHPUAO8XSvQwgLt3uPe3/ng+ZNqcMFTZIjqS0/9
Bues0Zn/9xDvWFZhhr+XiCTIPw78+0K0riy0bUBTU+C6SRvi1hH15dGUGionigsLBVPZKsRYcugG
pCbJZID94D4y2cK2p9sXsnm0E9gU8MuVabkxCz9Ql06ImOTOR5yXFUloc2euXzdXYRsnpSaFWrHY
+8YEiXJl+ig/6mzJOzx9ru1/nGXBywSnIRcvI20upxtNK5V4Ho+ud4OEab/q3LwToUE6kzc+DytS
PzwAqywjjznrybA76hRIAttdWnANbRMVx4s/Q7/U03euQnE7Aa0p4nar73QKMDRIo5r3j4q8xFjD
zBTTrjYN2ZrdMRT8jBRoO7qzEyqMZ/Zh5xi4x4Tzw3Pvkhj9TIqSPST73+zmCLrCE3Qs0wAmDWeI
kpjY97xN8/Is7kZr8FifBHRpqAMjHKOmGg4q7d+74gAK9upzMJwNXFLC4COMsdFldY1GiKL+E2lu
99XQdx5hPuPptaWzfNDmkoujXENmEgkjFkIZiQWgS93meM8Hdl4Aisx1mCAExCjTceKJYd6bR4jz
My65ppC+5OGX6K8G57A8Lcw8SqC28eBGpS/Eu11grqVnyJP/rZCcYt4QjfuU7YKI6IVBE5bz8GZP
YiSXZ7nlnSmBAxWYBZQWxRau6jEvxl+FHwSvK359iwuMsU5AMDbnRs/dy/a+mUn5LlZWIaP7QLrU
7lv1CdBQbiz3yR4SHCR8U3YbJ6GLlU64wtIolSL6CyT/U57E8ICM6xwNGjeZDD/upKxjKomzYBL1
yOSoig0Ak7WvITAmdD2mBnpouMPzU61+zhAZsRtX6NxDopwX8R9m520XgC+jGCYxily5VrE0R4eQ
FGsijQ23y8TP6GCJ80PqvGjODOu+XGPr0gXeCoPHpkwCbZ+OQHgSxua6sXkBPF776IlkFjM/d8db
7d1LAmO8bLWBEyuHOmAsSIy/P1YoSgrG2TTWYlzdf/K3tWDSyVoLXB24SNTXOlC5THyyMrqE/WlM
0TlC/2mv/w+VveafWcVka1SdjVzuVgjGQd2pbiE3bc7+oO4yKad3eUJAstngcCzJcw0P61YsDXlG
fZhCEXIKF6NWq8Tohe/si4z5ptJwaPuPsOD0vNIKFn8v4Bmt9B7dTUlG3biej5SJ0zSW5lVR/T/T
yI1hYUO26jeuJdzNcDGJfxh7uV5pra3Kq5ah4zUzQQ40XEedrg5+6u1hro/2f9GKtYYFJeqaDIO6
QWwKyNvqWFu0Ojki56qx1/YQskErTrh3zO2KLUofPP7V6cQyTFsLzX76eLwGi0qVpkhL7NSIJFrf
lFpmbE/uF99kJhUgWUf9LjXqX3b4QjwxWUkf0By9MKc1e7Y3SOEjL88f5MwjXrMgm7p6V/BaKWqD
LqE8Tv+pkfd2OnMp+nIaOaMBNUqXjQx+4dkvNf33v52saH3nAr2/8ky60lsa7JK/8P9hE+dHArlE
9LkrsgOt5jyhT//hNyWib/pnTNN3/MY+15tnjBAv4jfQm/OAjJ3S89dMrBFtgpwTNrU3RBhoBGo8
70U/6eX0Z6cC7n+qZ8BQc3FZcyWgD6+r23SD1a2UDaB6OaRbJ12nmFy8Djs4zT5CFd76cGR4n+jI
FSA5azH6oQycPCc3PJy8NWk084ezcyUTnHslCiYBC38X1QOwwFKKTHNw4ELZv/SNOVAxSaJZkWYf
yE6l79d8IKCXAQC5FaroCisj2BgniwisCfO0ni4HGwl1x8QKaPXc4Mcb1jmJv5/jg1ixGtEkcro8
/GIXPk5jsIB+4Tln+viZt1U72NYu2sdNA/lOXenB1MiV1XY9JzplY209XpI4nn+bv3rY2GN9zDuL
gkkMRR4opDq89Zr/b5eYvZHGCuSY0EZ7ngaRVqjOW8TQeOJtvvy5X6w+SUVqcjPVJza5t5zMdfO+
f3lgV11jSaPMarw8MOszh5f4ghv1DieUf9Gm6nJLB871gtCIF9BHDfEb9VvP1X8Fb390ifMXi+6s
fZ3j3eZgzbxA23uOBxUoXNRUVKi5s1SKX58MWZgDRMtcwSTAgOeCDlJVVgMA57AK2bwP5JevfcHq
QlaZMnqUX3KK/UJQq9/bsDCKZIfRCQdc3x+94Tb9vIaDtJUTy/h5LjZnPOAPrvfv0m7D6b8tktGL
loNkzgm6hRq7SLPow9aMVtlDwVP0zD82GcS7Y89tAzbgsvCCe9Z1l0hKetwpEnnLrwAi+5h/+f3x
63Du8IQlGCjNdhcFwEC8BAkyDRflKN1oJPkNvdKvbBkBBLQo5j82wyuqajDoSFJrl6/XzlCZkO+F
T1u9Fv5pcAle0O5xKWkRj2BoFiBd88W32VFQ4NTML0+zOKVnuqp+eAKrh1WhSbIJSxGjQrWVAmsJ
5BvtJJmYhk/+/PbZtZpv9wF5lzYxkazPELr4CnwVsdSLreoH/m2B8al6hDJQAS4oOXZfvwypCc3B
1zIzyoVSehTJO5k1DT+qpUTDNCG52POGFmLCuZKIq417Mg0SneZb41zgiBYJXtFbbkBHv/Iy1hO3
InIPEta5rV7vTK5iNcsVrrbc476gPA58i5GfHHaxqz4ofVrTfhBWC0bJ0xM0M6CkCX5ajBS1RHei
8v7SuR6F9ytFSHKNeBWUx+80XWJ3p0CRfrcRkBFyxelfKIIoVKkAb7Q3U665hNrdjOcMHfOrT8rq
igKlUnicWIxKSmgObSvSpS3qn9OrPGZ+yI9WYHiwVd6tzjviQT83JSLn4HYgFUhK2xoj24biCKFY
gsVw5t3gKdJB/KZnTpJjueC+HwDdnuhHm2DGMO860fOi7Fo3LZMIltaVeyYfLpnmWYxdCc1g1Xhb
rMFvtfXJ6JlUxZ2W6cc5eRM2mMWNIlQVkRPVIpBZjBR9DwQRJ5AdWtEwMONSgFhwevL9I7emGcyZ
kxr9CM5eAfDEWuO1MQbKgSmxRhf724VviDusvILisK2SUe5hlTDPA0ShN84ObubCCZtMEwc20x9S
wdHANZa2eI1uX/9sDKTmrIFbdn2CJksO8llSi+HUDOro5LfW7++wpH2crrNZD1wlderYeHPwfd3R
N0Il6QV8lXJkS30xhQJpBPQjFjxIjC5h+eLbvdHS9xg7NUCHKYR53/P6fq0qBcndTTqWy3IG9LYm
krf2OFt4CryRzcppJpVm4KneX+jAlmT2HeRa+wVXPzTy9lCWTKtb2TeMXSSLOOWoHzDgG4lwuaaH
8FM5JPmsjez9ZyxRkz6tPAfx+QHFgB0k8d4fOfCG3Amx5iGL9lmxTjEGfmCGRwdaEWIy1krEoay4
adxze6QRJqfIvXczYzNGJXc64d/HnwBIvgInZL+JH2455SPwuT0CaWMuE0m6v3iUhqtqZZbCepmG
UH00BDC/GQIbXY8JJJhdBBHGJUreaPVaWtyb3QESLORNzF9aHxnUiaLu7jM0TKBwgWYEz4fIVrnt
CmTEfrGxDqrilXo3e+B+IFDHRqr1sQ05PF5KOAcGuVBDbf1QHnml44Ko08tFFfeakpNwtZ1HfZ/R
5iEspoqpomE6spat2NxXQNkUon8t6xzxS/J53D2iBm+R82krHsEUGfWyvmRP7S5VmhCefaw0LiGP
Dd1g5C7e+xPv+30/2uA2edK1DpBvMZmB5Ihva7R3sq/l2cWK3HteFc14UdTqv999JuQ27yoTSdrg
VYUHcUBWkwsRnRUIDurmB7Ashh1GROGXemz04Q1/Bs88lbtlZK+g1f1zhM6djXpZvVL1TjmUYRxq
y1nekAbXbuw6Jcw4IQJk3r+5OPGtydbJAusKaCXxR5S0V8eUhQAsAA17DP+l6ZOExx4GAxwBAIHI
oAz6c5Ha+TGi3oyEtrlE+0dC/nA68eGL71YDTaJk9Nu9aUngw5eZSroOti3v0iSYk2GjAQdUIe0u
tqRdyO6vqNTR7Dd6RyMlHSxaMyaVgP0Rec9koEHtJNyz2D0ErboZ+0NZ/7RpeooohT1fPX6hT61T
69FBxADxLJrpa630NRDsWvSlpIghx2bdzSzK26Fmhg5scXv7Biy+qlcmtH8TdBRvnucD2P0LI94p
fZ0Pj9PBNRFdgRbI+TCCkDcqK2S+vV1gtdCMFUUg4/pmybqmdhgr1xaCAOGRTUYTRc/5gg1HkvuZ
Yylevp9oAoqWtyAUgGJwcJYxk0CitPnsalOMDksNwWIRDbjNzrBl2l44GxwmNaMMtcqQavSlpZrW
FCcpoDLTkMFep5LmLcWFNvn2MORqIOatElShF5mjvgTn6YKZGwWP+QdYNSKw78jOlrYr5ab9FJQX
1wTahVgjurQsH6bOBevx3wKLaU8UeHM1H0sdWC1Z2QEoYHkL1LwlqvMD59ZRbfU+3xg3mjMf8o9G
481oV6WDWqqxHKee+zxEFkyAojglLCoSN2n+49+j1PQ3G0OoKPhSQzH7kSdal92bcg2XoppWz1Ed
dGqnsYRsYQ5NTDim+z+6CMCjpB/WgX1DG00REfDsXprxTRsrlPQd+kmuRbfIH33DMDNPDBrMXCT0
tHgMRm4zLUt8xJuUFe9pB2qhiPasw+i+IjocWEHNb2LcCcuHd46YrIWzseBwtjjQEl+QPD58Z0Cn
6dIJ8dOgrDZGXwXT3GM0uX+FkXR2dWgOWYVQ2wDVZzV8tVNSdjfGIlo7tkpGi/TFDtrJ9lVKdB3W
ZxbXEK76cr/dUlhfvQc5vE22GmgpI5lBOvQmutYULLBXvdRz+BqXh0Ub6J/5rCJX3az0rLnWQPir
FzRuhDhYNPQIWO71c1LEdAZ9dtQCg4PP7XvrZOxOCez9i2j5aIQ4XAxFpwUQXM2hNGtzq+Gkrf5Z
gfwd4fLgcRYVcBG3vf5BN/zO+akIc0LXDKHdDJC+oi1XlX37AURZgl09naQ9xvk777ClnW3NKQg7
kb7BBPQhHMliU/TFs6olvok5ocXgLLbq40HoQjjh7SzaLLTaIw4YFSXZ8q4Yru/EJG5I2xnUluS3
3BYXA/NKPBpMl/tH4cPG2GM4hxn7AuED5Z8z8ilCR5cnhaD3QOPJOfHhQ2x0J+/oVUfu/Cwgs0Ah
eB8Cw1pqTZSF0WF5uOO1jMsaImuJ8OiYRi6KKneo2aJ19m+JWr0aB3XlH/e8B6KL5SvZYR8MGnTD
CI4qocjlc0JFrbWyURHf8NoaVkNolF3Gg7nSJrUTDZa/vc/orWU8thQMV4yNEZqwoRHMAkNT6zpu
UHFSzfPvKuQDec8k7nPBUEuxdswL8YyNrOgXrKf6Lp+Za+cWxrA98/M30NvASBgNQ74UL81DQLwa
DdY408fGZEBu/b2mY2NtNhm5Ga6/WSGEkL6ZE/r+ImQ00PytJcsZZQELfhuq+RxoUIG2+CPuMpKi
xDInTbwHb++AouZ4JVzMe2YTPO1O1DyEVlY/e2JoPC7OoNOxFF9nyVbtwrNIqiqU2xBzZxA9Nt6C
1GUNPqM4fGZOUohDe0YRm9qaBQ5DxavZ8BZBJZi7tXhBtV1dbszJ3VFALDX7kuhhpwdQu+94BhGH
+I+JYUcgT0WkJp8olnFed24fg5/QfpiQuIUzaqLiRjkTHOQc+sNtqZ9yHYmNtsSdgfBg23/FloeQ
o/6bcelqgk1GFo1LwnyJpaXGsUwoMLKjNblAUTHpu3GFsDoUF1PD59YLyOTyMyRdPuHZ4Dz9ThmJ
70X4omlUKHm9ny/rB7lNsbivBVhpPNuI6V1fhqAnjFLRNSHvvABPuPP9yipSm2HkRRsOwvOVjTOY
GVyNUN1tD193vqFKIX1x94pTA8ijaNiXGeRe66CqXdRpWLrFv5ktdLdTGn/rAbrQtA3hg4TDRV09
m5VgixA6NY772kuVcuzTs7LZ6o+ksCiY7wOcMFxFjeY4xuVfIzKiR58iyGE0oScGLy+lo9u5vbmv
RWX5s5Zc5/VQhStEFLAk2/ARa2I2XIALMOF4zEFHhTmiu2JPkSRg4to7GNXOwFYsAniwU483iSze
it9r+PFVEl7qTexVrcKsnFQlKZFhoj1mAvwert1KL5y7ef4UrBzOuy10nR6NtKoewPB805HUMGuG
fhqzf5FsYl/qP8QD1feDbH5B/KIieg1nHrwIMxtY8XGIr35qEHv14iyhiXkgFkYOQfFVckw4kUFH
SdU9RZwQ+khePnmCQrm31mYT/NoBQCGJcbi7DSoIUlANkJO0tYkRareDZxVb6JBhtf1j3hRTJRVI
fmT6ZbDvdqpgGicuQlZ22CiuudS713LYwLGR+1Y/H5QteG2OJMGaHRBP0Aj4192e9pNqIos72knk
0SDajNtDGU1DMuw3xRbJx+o9hW1NbUyVxQBzE3ejDQ6oeFXaBAEy+pZmzZomg9sAfJNoLfNR/ZFp
/EJ6kNXCWr/Mp1yo2w058ckAE7vuj8aah5m88e88WdanNKnb59sVpD+ydB/sFkz0rft6llhYlprD
fSQnYUjh3vxAZWumb8xiDAexLL1qqBN7yO18jwW52XhSeJAgzY2Vstc7r81rVjvl69ThXVUusnyR
2FD32+1PUd8p3sXpOOhauIDa5XvECpOMs4vjIGof5PZtYZ6WeMTgQ4JfE6WHXaD4ChbNeMWLYhA0
q8kYuzQQt+foqD+M5bmavgOha65hyPNfusgJpzcymbT7SCDn5yZszu/5XKN7maD36jS/6wQkhh3H
hSiR4BIQwqywo1iZ235tP5KPtueFjBvtY1PTlkmEX34kmmMIA0stH77H3CZkHWw4Bvr8nov3NhsX
ZWI58XxeIVru5+pJa5/L3gS+B5IqcuToOoROhwmH+udJGCggqsuZpoy0deY8QgOEpH287ep+y+vW
p7B6casbTHeYi7oHScy2HR/BaztPz0Z2CZmdA+xINr+y7Viq25eur3PXA5fNUbCLmNVAIkLEtw5+
qRhAWjwPefr+/4BYNC+PkRcO0+snClC/lk/CHNyL2RTm9tZ7CNzg0szsP5LfVesh9eOpwJ4pqj1p
ZKlXk+7Yh3eLOBneTHKeXsHBfoRPc+EIWcrVNmlt5l+QM4ZDT1TxAFPKw+IFeAGm2ssdc3ZPRJiU
kI5LxnVg57vW7F7RBf2joL+1LuSEUFuzXP71lbU71svbumibgj1F0P+qQh5Z8Oc1Yb7jBEsFVj+N
BjHRJtcPIWAZB1tNQbwnII64pmOK1hRpapcx43QQHCuLMrt8doGUGFv2iWpGZtgHRh1IlN94sks5
FMNH7ZwLLb0F9Uc7gB/35ql+Kvb3sRHQ+CZ9O/gcUOw1vzaaeIhB9lajK8rDy7NT4i9Y8gKVXUKo
mF/UBTrjSMzFE6LmbBZBBScV2nm2UedLfZ74Euz1bce2ZjdLn+ZGvBvr4Ar/6yi9SF5c/275TTHO
4ljcWZVH4LPUSgs3eOCp5nk3vaOjxEwyjXN3mtIsIU6QhIYKqpDqTg1Zp1kDDcXdq5a6k5krS7SN
EB0pLofoHgk7xtaHwI4tqz32M8V6iqICciTOp+NMOKjCvX+1RgM6snG1omW8pOzlziEZ77nTUCPu
LtOCwi7JPLZ2QwQVzbcwVEiKmICxkyiZeOKhICCuRoOsEsUZqq5ckv346FI96hb8P2WckUBRvGol
ssh6TtUhZc66x4bhY70z+A+2XnBXLset10oOCauUIGVO3cOXW/qriO5PV3h7Cc11HqHOwEnXReIb
ZppZDfL2ZDkRjcFd/WPzxn1aFMR5+7zYEUNYcxPKkqzo4Ku/GO/mMVszTCL15KKlVVgDJgB5WbOy
wSqsfPvTuRgoeawm2Px5T5KlJvnDyekaNcTiEjgSKBkbn9reYsbVxt0KxxP7/xZ9GRSIfyRnjzrt
pc2jfmu1DDHKmg8Z1xAqfE0INwSoHMoPlmC+1l0BvsiuEuuPOG8VMesxtnNxhufjN1l959vMY8oY
tWx7A8GACTzm/3/FSfK5mV3lUXhl49769NyzeUNZY9eGtM//oqhyMP54ZFiNhBx4qAElZO8jPLuD
5jVvvGazcemDb77SaCqsC+kFTUzFcYSrIaiVny0dqqu+Hb/yFOcObMNAdZhUfzS3DkObqcD4t4ZP
FBx1ZcAKSdZul/FfuTlYQXTywO3l7950Hk061INMvjQPBqjZPzKH6MCpUpEaNgwOx1uvmkdbOruT
GJk8VEDj8iCr/cEm8ROswdD6+kP5qyzgd3qRslW+fO5LFp5E7xzH91qiUx7uenRt39FpoBE9t2XN
weHHt5sq0kH1n75iTBk4BZOW+LWKSSQ59kT+x8yhWid/4J/7htRvmVmh+NK47HcfNICQRWmjqiJO
OAsafTFEYgQYyfgoseZMHcNIwwfeJ1iieoQGZUDf6O3GunzlM6MNZZTcseVP1NNosX7ix8okL5uO
rha6sZR534w2T01PS1P+MT/8dzB6LVQR4CJCEB6KBSq9NU6RJc7LWGpbkpApPuScasGKI2bhq5wB
kMCFE+q7pFrqXppvg/LIfpJMaLnfEtJVM1mQ3JGX+2JdPp/7HFg59hyT7NOWCjjzPdshWjdCl9r5
2PHyrrMATA2HIsQlc9mil7oUINSt+TPP5gm9pD84d2+X/gHe3F72Rq2un7yAZHrf7FVjCYlvHMoX
MqYT6s2A7GiNtflJ1qMJQAj0jr6hLD+iKB/UbUFGcWXIymoBYfFMgKEuAeWoyboWOr1LX+lHl7Dm
uQDLO4lWgdfKt4g3SQCfNDn8gxk2gywWOtLVryhgbJn+4QkIBktbt0p/+zIzKF46f4UtSNmPO/ue
T6BRiBs+o1z1/2ateijQi2gfvjnjwLpf0KQsHZ2Tx/gvM1rAHfGDlEPOZZnXeHsYYTwWK+kLJgdg
OqQQAuR6swyrmSEc7lu9wDWdkHyM/FJ2dLSTK7cU1S5B4lfiMOnwJ+jKJDeukRB9tYQFx9uLbIUX
EjFnZRhZIxgYkGGKGw02m18ZO2haIr3shMWs6SNMw5qjusL4LQFZKLEyCwxNPudZPE0MSCicWIZb
r9z/oYZw4N8n45sEqD/U4ofz9+CQ9w223uCCSBnPhdwHrMxQ+Iw4tQVk/I+ZkQxBfhy1Uuw4AhLS
UF/snSw7ziwnrVWlrcGYUwdF/2CoztKa8rqsEPsHzaKCujWMYne3F9tC9GKMt9QmiYcJhYow2VYq
IofuiF+mWxaIhYRxDjnwKGo99K+/6NXZVzMToZbERZ04j4qCF99Qj2upz0DkiI68P/FCctimwJct
YzutlVGkE7D0it4SQAPfsxU+FybLKm0yCkXsSkQbteliqsM8m1Dse2NhueYDz6H22qSIYdp7bXRN
Dc1mnlqQi8w1pWsdF+uz+1c0k0njDHJpe6M+HQQg3sOBl7kCykVEz6ML3kJyL5RocJ+WnGC2Ueah
j92IG07Vz8Po8TdsyVACfTFndItW0KtUIvNI9dR6ODZ8yodW8kV+e0q0WiEFQyrDLSivXD/A1BgA
gGtM6z3JFhMVkg4v47n8Z2ywaTMRgrsE63q6MWJYpjm4sNYqg2BlM0X/engfZeDQO8VqC0VDWMBT
iK2Ha2o9Rzf56/5Ge7+btIavORFIdeqxjjLJtEAXgTBSGJXOlzaxb8Q0bAdBZU9qeuTNyl6HAr5b
dqmd/mhH3A2TBNNK2/ylT5fLeDzzbaiYTW0qm1d9Hk2XYOUUGJijM50YbOi78oyS9gnfish8UbDj
E0RpKiAE7zCfVrPPW46iPzSmWpc3KtTsKncVDAp/lHgbyqepM2lul/Ll9/LIMsSf5sl3OKodCE6Y
Omwe911Q8VcfuwY7d4O2uf9v7qQUPeFLn3qKR0HeVcuwpovbV2NsQPhKYjE0pOxAy59SCj26FuGQ
OD6y4Mm8nIaRtb5hPmIc8Int4+sgN8U43/BXZS1V9splKrVgIdtdww66avZI6lvMwnLQDkcqJaX5
IeGU44B/ih69iwobFs7VaD/AROBej4SN0/m9HMKR5pNsMHdZuUF/ZN6lnqQfSPZUdHiG8IMvezZd
7lCsHkI1OMFa1qqcdiYlY93tDRpU0eLHfl70E/iEtp5dgZjkfUlZJgGj/UAGwuPmnfa92B9A7QV1
lYXoXjhCp5sWKrjnHjmVO2fuTQQFOoV6N/tc9Sf6TVsq1ViBtGA8yIiyW78sh0L+DwTTtBGGWFMb
Ebr2y0h2w/kxK0sti66mOM+bRf+9wg+PTHVgkZM1meprCxspLxQnO7pDHXN9icZh2DoHk4JqXb/l
AIxOueuQ7URdD7w5MWMjw+BUnjT+GiYHlHJE4puL3/1Y0unoBbNu0wBHSH+AYJPzgmvRMor4hzh6
xpYzjR+nKsMcYIePkocHU4Cs8h/quS25p2D0QVhBVu5R8eEpCAR/OeJ/Qp/FxCjvmK/mWagkjqSs
uj1PHsaF8h0Lqs8OWeFKw00zd8DSbOboKHzBdisj64YtXuT7h7DS74Yq3Z4jHMy+tuXUQ4htpkpq
YgIKFMSv8xFhUMs0rqQ3Tw4C0sTABX3GDPh8jGVKeMIO/FJr9rkVmPSDBkJnnkT+jvFQWgQH42mx
MT0YRF1awg/UwU8JlQ0XPumD9PRrKgphLYmG1AUIuVc+BIjFbmUD3aI8Emkp6w5Rq5UYrgZwMx4W
88PDsU08UkWKIkUbVXvW5ZhtiUWMOXi2VJBlluVWgtIA+qnLU+SYY0Q3245xV+59UyMykfBmFaBw
95/dhyo/CcjS9cRQxFENXx62xseg/Hhk6Db4COH3FT2WphmwRc3BAnJcFYDAQyRJz4t1pQjaKz7B
z123Zr5/1Kx0+D3/jo2ZlX/dolxNRRGSXfhYbU+ee53BaR99ZComp9oANrCsn3RF6xeFU+eKmYK4
96IgTWAvzqzZovvu8kx/3fu6HMpe6nvraP/6ncn88gyyr0N7ZKLZ5ct2/rSi0iRqj9n2WQkzUYdW
Dv4zyhEAsWq2rHZYHMeiVhvHMi8Xmd0p32dv3EBIEAgUlQG5zUjF51+3uJhXHt53m2OydCTJDcsF
Wvww2yHnKmPBdusKqMEZdOPQY0vvmNOusBtToAap8CnbjIGkHK+9KeLGweJOlwmgEaSasoNrSq/N
mKIocd6gDXI5481GHMpj3LTYepe+iQgLv1QPEIrtD33vy71EFwB1H8FGkljw7qzH8XoBAmu9HkNb
ff0iAEE4Ff5gXcklzCWZjT/fiM9BBzqQDktmkNjbf3kt8sKWRZzmsLk+cUpOdipEPz9bwynC8Cw/
HUFAToup2DDL6CdQI/vfhjaDHq1m0ldd/SnDBQ2OtcA1ws0FEJb34JNY/bQkT//wzAtiL7SOCkNA
oa59Sm9MABVVU9Tf7lWn8WTvQ1tDcQEA8JhQykTGXiOtBbOjnS6LoxQ0hQ6FMJo33gbetx+Xo7uK
+mnHRqM5kO0JAGDxI/0CBoQ22zB4nlLxb+7BF5wUg/hPg3smA+LULHI+kce3LNkW4MnzzRy4eahE
X3mQfREbe2xzdN5AHlfQyc7b/T8jeFoGLVLfle5J4FxLHWKc3QqbFx8w0gARdO/25+27Glqbha8S
NBSECfPjLOZRuUdbNvUdYp3u7nIZLhusxo2vtVSnhjBkaOkaBQC6BPkj7jpW9fw8RDFkQq3aPsD0
MoKplwEUfgCxQcckyxXm8jVLWUaJnDIGZaGi5IPK2d7af8tE6ZOrVPihQ+hsYAGAy+lc38tLzPsA
fil4CGvGxodlPzrzwZD7RDAGYlD71OlacYcV4gPAJtqB82EOBRyC+dpkMGTBuL0JMVNMzVyhx54g
M6WkfOxgZ06YhAA36MXTHD8mqVoXbfY1xeOJ9OLHmy2FOsUs0dN+Oiko9PK1oFPoKz5v7pVl64CN
VKjtaujZ9UH5v8SbEUG8puEZb94XzulviD1s7Rb+JPlCywAUDK70z5119cU54vq21gLftlnLD19G
WQLY3FZtp3hJ4YacwXC7N9xcfuY7BhKyd8nYQVygjyrbZ/u1Ky50mD9SkB3+T/ZDtqlHeO0xFQHc
bbe3NZi3JrCeW5anbyytjEhchUoP89I0hUyQMRA5+rgBDT7Ol1rd1cEU3WVNM13u6J8rsj48bgeE
/EZuNVDwp47JuHz/KWI4QUnv37DbHVXy/OGl6CKhYhr1nt+WNyi7ZQhBZzF5QPbXICT52OoqLdUf
Pr0BbzgVKvWZK3e12ptGYIjc54CQK78Eo18XamsFvh+zFczcgnXb5s/fHax+zRvE2o5x3SJlXOlb
cUleTHSznGz2baEflnTfSvPLbrFuftiRp1JiGF7IUj7/pM4V9EtCZ7ZdENL6VHvcRrCtM59z4Oxr
UavJ4EnUk0iMEqFq9AeMWfu7wu65+YDb9vLc7YpGak/cmi7y8V7MBunKj5eyYb+a7VO2TNe0g8r0
mb88+6pW1B9jrPDcAkWuCyXynaw0qVf6SOLGUxMmk14awGUJ9SF4zmt/RjAB7lHEjZmCspaZdwHm
hUevSeDdnFGr8KnwjAUOa1uYNfa96+aqtytAQFDFyAd1iGA/EWik+MTIEWkQJ+JD9YSlsGMWqWs1
LgljyIgn40V2kYUDhQ4lCC8xK1gu8fu/dy2XQJamENijj2xdVE2ut2kRkNXGlO0pkhLo7FVGMktp
KEhDypHXSUI5lKpNznk3ejai81RbkTGv2mf5dlBi/H/3yIvsabJV+puiLRP59QHYIprvvERn+Fux
L8vRQ3HqC+v4buftu1t7SucsXfzTfxYOaeuxpPBgWHrCOsHh8gXKHsjOrhVd8A/rT+nZeejv4Ez+
DpwB2c3m9n7upQSV3aoN9LrE2r/p0zNXiURkMZjOYdaiNNBKufLevQLm6rD+pgK1xrPnBUEqMmWz
yg7PcLWalw212EAsBrR296eJGGA67E5g2nTwgY7bjtfqfeXzHq4TjJPuuf/dZLUtHyImtDGSBMiu
ZiIB9Z1Bpzoac0Q376tRs0HvF2mWQ1uANgQ58IS9mSTq0eC9cyHo8XXi7VcVimNoTyXpzwQXCAxq
JVffAAfw9QmWmJht0Zmra8EnP05hHB0odUs50mbI9SbU9BokpSGJaWYQ1YGeVJVUs6ddbpoWgR1h
37z0FfpmrrDEVkAWpAeXXUOA19fBAfQhA/SFbASNOJPlYpEYFXwgT/OLRkUGMVh87iafKbtcB599
jsP05fvDE6HW7a2XDYY0t7P7wxsRx/wgstgfxBWK83D7bYBkIdwRF0ZlizHetM62zNxcWVmA/eiu
tte3nthfIqKldRwOBPdBFUAz66cYe5e9xIJ8azj2hLyE9yTyBGKnfcR+sA6xayetlqlXcmUMteen
LD35Itl6gvsvTdh5cZZlQVZcUKmcdrTlQPDEmNaJaSnUDv/aXs54GRrEt1+T2h8EhIBIrL9MRWTh
GGLatfHdC/Ty465BdFO+PW2geyXuXFUD/8Pe091xjR48ldiHhPnrz+OhAIOhSP3L3i9B4zuO3nmQ
LEjA5g7h7eQWah1AWNvLy1Er6NCxbatgKwVMQTi+/aX6SziLjcM3LzMFpRoCOLQSSLr6vGzAqVx3
pE2GIB5nZrGiHMMvLsMMWz9HF4l8k7QJlVQV+BTHX7qWr0NQ1h06KHZ3OEO+/Z/xRzLUIWkZlAVp
oHiacFdImTuxlSG4T+vD443xiM8gCU7hqvswUYZEB43qAzAiDY+Tn0ih6E9MSfo3dA9SCVYb/Ayf
9If8uN3+TKZaUsGtpoGfZod2jINazVhgOAtO4979hgDAJOYvugaROLasoPFHCEplUv4BC8IgH24Q
Ssz8USfxlBFK1HX4z1RxSmsjTEaq3rLd08vYxN12Tq5tTxAAtALc6z39CGOp9RxxwutI/Pm58lWE
LF+b2etrOZl17qex01P3SK0XHnfttyizSanwItFJQteLvLPHo4nzr5yqIE9kNCt78yIAjOInkbUF
8X+dz96AZFR7I1UqjZb9LB2BWTRQ3a2FyPb4AIDXKE9PazoVzuPhpj5nifzM+geZn60SvAt9Irz5
0NOMxvrAi3vkFc0wpqsOaN1ocKHJGijTpzSwrKurSTUvIM88jcXLH/DjCUMrDDH9D11QdVUREBzd
yxGlzX1tEeS6IMOtjbCXGEIB8y8r+i8/SOc4FT7zaD8QQy3GEVriDQBdXGSQlRMJYeLlaStf6ZOH
0cODBRVekkU9eaER7Eci4xAZPHwvruvAI0z6w1wcGju9qqjSYlr6Ypm/a8eh/HgqK5AdvDWmQXfZ
msKfojbMohoGEwX/i68o1JKAl3rExxWOoziQwgNZyuuHYxy6yKN1KbX9qXAds43uPu0/dzZCelAw
vvMhNrEwhjc9QZg9PsWN4MA3mUjmpo5T4lDPTB5cah/UOeFk2HRI5bfk3G4bOv9/jwJD/77Yb52A
H0gyP7fJKU61ix6XuemTpCU//yD1Q1tbs6GeJZzQSrOivptTPlFkJP6eLKfSTS6girLpptyLoXlu
OIue3+c8k4M+Ts8p5+FIrbNW74+8GIxocfRajWttnrs/c9GHyqnB47YwUMeg8C1en4iAbdNZES7M
hSd4nvLIDxOtJh1/5fL2Vl5e1ct0CI7N0HhhGFyOl1zofN8rUBbVvfQdVgZk90S87vlqUzGz/fWy
jwa+gph0vIL0uFDBmbAHYoS7AIdxVIaaO2vawU5lRJ+pNRUI4WsmV0pxXhMWxLl6AMv9BVlQd7go
22126u5UfwUXQcX9RWXvj+kiZBz0VuMh6qm4W2Pt4opW5cywsXH9C8+IyIFTMMuyI6t6fLtzeSS1
W2M0qpZNJiqk+dJcrfEgDVl4xO834KKedWJj8Sio9DJjpxsebQchw1XPaUoVBUCjpPaXz/A2jCFX
EryFx9T+gllTvv6mhIVtWTY2XX4L+Ls3VQ+JNtFfqMqwqTb7jV5To8ZDzyVYxFxB2MEFw7ybYMaa
sqAJZISJ/yWQrqUj3LrxpGQgRRtEFGvm/06exA06c3NiP5IXLw9Er+tYtGOUnsNHHSzRCJO0v6dY
hGH2SqMyyrnI+03YVd/HGsjRFvmfftdZchDkdz+EXNLnfDnOrwZOko2WfHsYAaWcCSrXpqwNy0Zi
74tB7Q5AoNEPeZrEnurWNyoPfMag+UTkXDC0e7/ucGfTACXykr8yl6EqemTQvexBV6uR0QmwulJg
C9XCEmtrSeTa3LR97eZ9EqfHiIDbc6AMgNwxzOKa/PkJEXrg6fAPA+CYyJT9BafJjzfUs2lq8rKJ
3tKovEIRCxMH9X+XSNccv8KrmiMO2wR2VtzLRazzGrKsY8Eg+cQcbSIoDSmNHllfdIZGXc42oUBV
Ro78Uee1To3JT2KaIOouQtS+zU+UzV5AsEDOWs09aC+d/Zuk4dsEQA9ifD61laUIjfgLLTyEecUY
q0OYD4mmHPyZbB6PXzHb5uPx9tAQ61rHwEtRm6EgG+0ReWhY9oUT/IaG9XqFhC1LMGnz+ODjPjCx
uzifXeUi8n02fjZWYBZd57Yxz3s8SzkD8x0S0yOV9FVtHi0zTWBVtyTLgkS5HKUz/Z64N+1akeYi
y1uRh7XXl/I3osX4UxvRHSXU32S9xgHbFXq/BI4xyu3NTRC7gim9L3oFvb519sjV/Srvgw2FpBVy
Osnb9scQ4JstBxuoOvZjDysm6Lg+2vadij9WlOpT9ccCEDV8wkhUgnbqZIscBe9u+/Q9zXZIKsey
IgQvR7RbnhNUpunSM80Wn1K4D288cITHgXNU4ZtX0BC8rLrEh6/qau6RkfNqYyeHEZ9mRjpLa/tJ
hvk1LlgqlMW6knKq1EUCjTsMDy/YQpX6+JQGFvInOCOvl1HOic6RImEv7agjwhYnQaB7Q9giuOdP
EgYzOriLujUhQiMCWB8a7pt5xPwS8gBPRgy61sPRBmEaVXIuKYUi9CKkgUfxTopxS5v+pqGdrwVs
8VYuUrZRmRDAblgwa01L9Gk5lhYW0lIZon3qn+C7NA8Xlcn1H2Oeyx3iwM6goBqzROnG3Jrt1VQ9
5RU70OZXp67Paaq1QBgmZmV0WQAhrD3eeLaCcGqIPpSMYN9fVSB3VAGK4BI55s8Th6CrnSjOaC0J
io17TQY+lRIxI8r2TKp/SpRhYKtjx0JIMUSbzh+h6IEAGTyGVRdWLlAoWI4IS7n5pmQKP+oMNvTf
03mH1Tabe8JzyRYmNga/HIzw76+hwLivIqluVfrovOK88Ef4jQNKmNA9ATBDTP9GhQaqMctG3o/H
kWcgFWm46v+dgPeyqhRXcJb12Z+M6r+Tc6ACMeGDGsclMPJ8jhVL8UYvGSLO0ftZsX1Pd5gSaud5
NPmH684qzAAO/Ih5yka4tlaEczWT5E0KUKodEqRKbAJW6qrECMtUyo+hS6mmOCtHEAAjKyQsuymn
7xMy18zm4bIlpxhYNFmnAUyFrelQBjfN9kQXyzf8BO64QAkj+6cI+NhJeRnyoD1pWJ/q06UP/nX4
AJMTJ5MOMqZKtrTTTCxrkp3r0FTIgX23MGvxdJ5c2MlWOefswt5WW6X9lf+g1hOxBcNsq2AkR25Z
xJnCSJklB9gxm0pQ0sCpM7nBmms9f/IBw3OxyS0k33yXx5QJNtWMmHUchh3gVzHvq9xuGE5vPGv4
3GmH/lnB1kTPDxii/tcf0qyXQTahNCrA8Prd+Kqs3eDgMpSIVLpNkCBI4KRG/lijfDXIc2jmrWc5
CpetvuGjNIxh0A7HeVIt5n7jjWEbg6RYbfWdG6jWrhhr09QnxbnS7v1NrjRmZIzm7QXTxCPvwDpE
7ERzFbebw8pBQmNEk3YnZ8tPXK43rXzSsk1WQjdj8aHBnqzov4mbkkxVEcsV8yHM7xc4NJS2Lzl8
W3fUtxYi0kvYtkLPu5urK3aU0jBQXTneNKs+qfpa/eN4e8xhCCh11H+WMRCsTQaZT0NVo+aPNsVw
skxjwciARX7karilzEXT1AxMxZ5pO6K6KxE2FT8ihWrKUf1DOqiMpPHCeA3gTfMQmxLluge12Cul
esdJp8vtsPw15UOaD/vm1SmufKPrVpT/2tGSpxGy03FHs95sVCz+lMAX1/O3DS1OEotusaUjnIjA
P9OxWY77ftE/QcOsg1cAaEKep0pnzCg7pWcj6ghm8C8iY29TCDxAkpdBWhdbBTtsqjY9NQOso5Ex
Xf3soolGA+vFW4o+gXhJrrT1DgaSWT+xoP+s7lmE7JITKDhcp4cil3AtxKLIMRHd62btKz9kgFuN
IyUUJs2CBmsuEO5H9Ud7A+O9iCmQ9c/QVkY9LHaIYWpEUXHu7GimjHzM2BGVzLsP2GNLPjEgtlbW
DO/R1iAcB1EMyjidbNHhki1IDgr26sH5HS3650K/Hwupv1Wk3/BResLf9VeuZcUNicU6gdWmH4mb
uc9drjX1wPs/fmDe3KL+CAteg2+CJeY81mSNDTvNGgDTxY929iPYi6Srmuo99mqvfR7rDvwhBIXO
bsa07tuuf40QDsGXKr2Ij4F+qM7P9qr9Z3aorsFUiryMn1QiiwL8xZNVDuc1Iax9E+NONxG5bAKc
DAA4hm2o2FQ3/urU/tHHsu3YAKH3Gz3XybCQAaH15A5OVAAyXw2+uMVU1fpPMh1qcma8Y9EBZMwL
Iugt/YTVmKG9DARupxKUKNkzrtEEddvRE+6pmUk3cQd8NBHdB3FW1PahBeqnnuY2dDAfE55aI0aI
bwa3RSSufNh9yaOmRSWf3Td23hZNH+P84W1HCeocfUYx5B3FzQGEZxjCgqv5EHLK5jX1r/oDtWiw
yt14gVk6bbFnnLBhOnTuG5OZ9VXsI8ufWrhCItgOtBCu/mIUY9wEcID2/YqcuenwxDB0CGGh2nVe
uZx18dMNSveqdielmEReFUAzFtApD6R0Nl8PahDwTTeNpXx+SHe9LxPlYAJzHqFr0UD9qF53qGui
whU+Gur4utR3jIGD7WGxkk0RKbqCMH7iI6o8zaPqzgIRGOJWS3t1McxkXPN75Vnhux5dOm2e5doR
wh39ohJ2l7Mg3qfTeMJe2k1nh23GcYYo+EW+W8NEDolF4MOhkjmvS0dnzQlRaAcAgiT/7bOHUQaH
KijC2tFd52rY1YhSv/NvSPxU270gnT/IeY54TLjnLVlwmF2d/2GLwsOT4LQ+DtqT5OlDMsB2AZbY
leexlwXdQhfRSO8ifipP7mKGETrdIbeIW4ZQQvDgRqnNg/SsffoFlWS7uA9Hpt1zUE9SVuncI8gI
RKZLuNIuPJE6QIowLK1rF6Xzf0WhkuCRLQwcPcxSzwQhFRiwBKTgeAdp+rTCxUAXgCemssEl9wtK
5BYCFpDj5E7WVjEC5tI1xwXUkf6dmfFuUec8W3zh306leoA7j8JQTiKQ/K2S7Dqzn9exBz8KA8Zw
r6nFgh7LHAOs4T7ARNgJdqHbTwTDu25Q5Fxjh+J3ZqfzGZvNDR4I9VEwVYzteEi42jKQBc1CKcjm
6cV0DjqwB8LDEytMVrJ2Ve8nG4Lm51CYFytRxpIWqtieUoDvO/5INOo208iFbMVFc51QZW6keDEQ
FNlJ9dkkwhSjKC8FXLDU7noKz9HRkmBZjHPo6lCJlGuqJh4BWrqPNxORY+QHEEKFYTG8Mrt+TdA9
a0g9BAL5r+L9aKTo/I0X9JWYhmzeUOHymbIb3+hXPaUWuTP6NcGK/tzi2RsIkFJD7NKcs3yJsVNu
Z25ReIn7QmiIrxh6wco97YS9ztfzJku4930mHl+T5Owi6ugQprPKwq1EuW1hLCTNRQMTN2V/TXR0
5Lzqvnhm5/vbzGj0XJa3nsj1HgCNTkQayYD36RypPWFWDVuwI7N/j2LR5ShDC4okB4Vu91Z8gZyf
83i1BBXe6vl0f4IsrGtSWoD7C7qJyV2ac4waZvlDhXM90uv6M9ZLhNCPxweImhkYKB+aJR6LH7MC
rMplD5kGMvS7OATlwa31grXoqxf111s1dU/0q5FScFMM2DQRaDQ6vFVq9/Oumb0unatrA17VoKJD
kKNL/WCP7LrlNqgRfV+UUrmxCr9vrBu6mGn6/Gnjm2A8jreNiauHEJrZYJAGO3LMPg6VZMG5dO1O
ivmpBm+l1nkFWAnwHRM87IRyskGLcn8W+CiKBrdpIDaklwuULbKF/WdAbEV+Rxz8rL3IVDvQnFN1
iXQ5XHf5xmlWXkRkUvPBIpOFqInK7gcOLs2KCndqonE0RNHm4WQ1aTvR3LiASg2Wc6f1PANYzuz5
LPcudouv7ZmdvQR07GFRqLEVvxmOUar0ibGYRCcsO/HDg51UTas5/MPq2FSZPKVyzp/J2donkrwD
KIH1aTjP3uwsADUa1VTch2DMvmRjTKHzpq/W62XRwF2g9EOejxP0hjfekCHPcvmV5wv8lKM9Ss1u
a/R1lYKqytOapMNvCLUppUjBJq+Yey2xvYniL2viyWtBcjRAesGgMN3/XaQbziF6+T+C1U38NUQW
evD+O3PaGtm0OTacXVRZXifdPJsE6Vjv1kFOnSgjR/55XIHstUqO44+14VcRpU/lor7d4Jm/59P/
WsAPK0Qu/Jxdrq3ok0NSxlEyfNAe3op2QQXImeqLm2C01HEfDhVWUtuBpy4k/SApm1h7Jf4eEj40
hAA4tHQx+/uOLy3hOUNPI4Fw271sFK3NBKOwy8r0HMJm9ZlHwJE+NonvI41w9GgnRgz1LtLoaQQj
8HmPFOFS5kWWrag8e0bj/03JNf2e4zC7JD8nKk5GpBOyhLfXVtP/NWaNuIWIeWsr3hNO/owDkcgD
fYkbeVbpwOtNN2UbM9IoO7kTVpY0bKchpPkTWOzr5pg6fFxmWc1YyY2ttKomqMGbJ4Qkm6yoNkkd
tsl45mFTfEsC97ac7IzlpZBGynisWP1ZxQAog0mcz/mDvS440S1EjZ0Zf096AJr2l+6Bd9dPV/Cb
Il8tzj/mWprAHwDYdaHSwb0rzdDcGAqqo38JivAPa+ohnkrAEAIpM+lc37e2GaHvOv/DxeZLVAVf
MagZKZ00QOTQxk+wcnA7/WEG7RC0jhdTaEw/JV3IUid6zstacgvP80C42NDxq9zj5SZpHAxpPY3c
eDokXxFd6cXgJ8lLqX9FgYl0ooLZbMxiCY+UPypfsIUh09B8lUISbOVzawI9TGh2fxxN2aZ1D4v/
pWhWF/mUwwFxjcVWEGboO7he9yFllkzfuZHQJ5yNp/CdD9wNNPq186OTon+fX5vUNfr+eJbbp5QB
hPG8HsacM6RGlSdswaD96/rgcpaa3qRp2cnaitndELEU0VhbIgBWI3X25AsA9f19Qp7Y5K2jzem+
hbOhPGCDyRBuLVj520h4abqEDgQbSMdO+lw/BjA2N3D9Gz6tgAAL49vMOeIGVZw/UOP99R0cub4P
R8yxWHRlBjCE7lS+EZn/rmTphthagOT2QZLcL/2KVT8JpQ592h4OTImb0Osuw23hxUy9visXEe/x
G5zRnMPLk6JsZgpSQaLPOWdbbzsaK/mckcsLDES4tOsXY6HaAp0Iljy4+hL+pdZczWcmkAX/pYpG
uUdoiSZ5pha2IooIKyBdPaxKSExU8eiVmZaniSoudtN8uVMZi1lwsgey8R6JPmVG4XXNCNCqmUN5
hDk4RGz8iN/IbwnRD3iQTeflKqRd/ShnruTUVHoMjSczT2c8NAv1d88hnujgq5656P8rULKUdtRx
95bJmDCz+smU94DldEZZBWgH1olJHfeBYfsmX9F8Wi6uCtf5PrNYaE60Anz1xdk89r+dKECMpaYE
flZZkHuXi51URnlWm2+2Nsvyy3aIcsP4Xyu6Uc571w/X8gFdy0ky/7HPYrXZLQrQ6mOgAbi6gl+e
gjgJ2yBnypJgPevET4KC4I+GmY8Y+tYj7QJ5YlxXrQjcwqnT/6VOZLVGY9oDfUpCvz+8fcY02Ts6
H6L+0vJLZE91bwuLQA/FT1NQcLD/1zTV3ioJNNXe3oqVf8s1hjrh5nibGZ0bGrgcHhPAeeQqFucA
KqsDQcyyjTFBQzqES8yUtxn1iiS/cxJZovtY/Y/owiiQptSHOkiRCcHstd9JWh3ED/tQbqLHDzHc
wv1b4blqkYWkyBzZqHesC364VqxvXcuZ4bCn6zgfcoaLVGCYkXlvIcIWe1U+5XxXZRJAma565/3k
IEXMYnzmt7BOxUp9Drpuq7TSqsDIFQYTSo8t5uVJkKrLlKsIB49xNU3b7GaO7dmQkh6mglnNXeSs
MhVW+IuFk/LdCMFfS/Jj8U0LrAo+cx6EpMECtxiP0oLi4SVX614r6BoqIxCzU0l2aljw2a36fBlV
CtJncMcxuE5wWy1sXwiC9tobbjT060uLN12D6kJoJNV3RNpycx9PNhx4vKMRRhtFFSFqdjpzL46u
OSlCeppl440EcRDN5yE0Aci1gB8MBVsXXrssFxj6rPvnA/iOdaJBMwjlbvy15EXgbiC8D89IhcW0
6wG0PqkLupih4Swom4QvCKeII/VnRsnyooiYaCqdaNqkPuKH71nkZduvgYwwLDufRoW9D5sqTsEq
40+rGPp9uVkeYaob9n91sZt3dPe2xNpZuGaUAXpioikUSPNjQ3hZHHFPZGNAAEYmEyDKJoITlreA
fuWSQeErGXJuHv4t7O09Yyo7wRw8WooLy/UryeMZ/cbx0Hk2JR87OsZh6susgdo0XgKi6zj/z4Qq
hF0Jk6Y07Wr1UPo9aw6mXTZ6/+vr92s/etX5LJEz3ZiGXC0WRAtawWNQSxRdA+WoNhVE8o2U4DEX
fnew4EMdLdeZduKAh0iDBk6ODNlIH+HJrMXFGzT1HaBUQbft0bsZYic9lhzAELTDvWkjoDG+78tQ
kpq2iUT9MHIWnyEEh8mvN5EtnM979JHWhUW+sSf7vgcwlTVtYoOSe5C91IhMiGi/DhMbNKtRzyzM
pevM6qp0heNJb5f7JeMcd/XPxSo2wzCMu/u2bSRH6I6vRZzxanNpw6eIc02PsENPWBK8hnJ/+qrP
/aV/jSQRsdL2au70El016ZLUA2/hc8TpAxNxk8/p+qikwRKyreTuan6avuTdiFHVuayft8z+Y2DI
g7FJjvj3xyCzT+O77yCdTAXMTcyFIgUkx6l860uiLL2+9ASgzqRSWLnLF0+M7kBlqXXyQGKBLaQr
NeBzjWQoIVwMDZ3tmF8eVMFdi03fF4rF6g+d5P/OM6WbCwUnmAh/sZmhlT3RMxjsMuPS/A7AQXJy
bgjNnPTwc+Y+6KeqnogZa7agID6EKXZ8SHEUFGIxCMWK0f9LJBrwhbnjVojQm3igKGzoVWsOpAPi
QtqoSrWxuj02C6e+kJd1DHuXQ6uH6KA0YKneeOozO+vST2E85xX7V+GTofbC90RJXiaWT7MN8kUS
/W/1aU0f0UPkmnvlCi2QCtrBr8QH78HnEI8kBstWC3ZlJt3BbGVDu2ujo6j1XXOncdkZGxvdM8Lf
kNE2Uf2YQlTjJ2sCNJ4f5wEkqMyajDqVb72/mcLYBxWs1sSeo0rgXYr4DhHjmf5MC+0n0Vy9jN6b
+pr7rHyavDzu3QkQnkShyRwfA+40k5jREHQPbVwOdI1VqNZFBPIDqN8jACAqoF7bWfDYmiu6XQop
335v4yCAVXbv5r82rv1UyTbs88GB+lUuf9Gd1CKZScSdf4QUBMhxYTXaRK9NtVbJbKdobqHs+O3M
WOdFE5u1dWyktdSfaDXaUDh3FyzDMj53VBb3gaA1suk3wbk1U38khnKhITFx4vYSEK/ofmis7LJQ
Kxi2tBZhGA5LjCgT0xdeF2hWJemNnxmQPx7irOhmoAJuQNTx64RV3uruagDUPRU2ap3biOx8bgPV
8RRA0c7ivRSo+mVKYGd/lDx7CAxeUd+BN87/jd+es1XqMvYd9jjGuuVrBDNlTBLq2yqtX13z8th6
rMkcolraZ3T46kk/fbeA6vHdUzx2MAOdidNmfUr3gqqgtHwHdf12yQCtG4dRZwXLS6eqiTjeT2F6
ESBsh2denYQ+7o4BwYS3n7e2BnKJAaBGzHM/XIApeDSn2fXaIjOa6EVUGmOEieVTYFJUHGEkeK2/
Rb+Qtb4L7aJY6qVdQI+DRupHPBRCCe9HqOzRrX1EPlZwPtro1KFzUTLT0nypQVud7hkUiYsQtu1g
OrjEXHTXWUi9R2/zma+RZT13CIaon9mwW4oFi8mekgaCKNVUmmBpWFoofH3uqrco/WXHNYPJtaY0
6sZE1JLjHkoc4h3nGyNek3Hiz5q8MWs15HMGbBlnNjjsYosiq3AMnhhCfcMamt2RbrKGbEmmUb/d
qM2+Q6jjBoV/YHy5S1zAzVi0cqcmyKdg+w836Ves1p4AqEvKm8HiO4cLOf60DyExO4EYgzTPxExA
arq0hzX7e7jkgC9quWDW6Wcz4yJl3+LDW9G2U9jdT2Kl0B6Ds5jPZZWHbWteTK5NJFpFrs6npMFs
MyJYx5CVxcOCo3uGpn2o3rCOur29VkbJp80tSr2/rltGf8Z43WbDYCFb4EyaM+Mf8vNr1PM8VjSx
XevVcFIKGMgt6cbvCh8n3JmiwRCpn8dMy0zdRRCmklJ/9hDzKFiF+nwPjk0UinLU+e/BaViqwBPe
jU+cZMEh/o25fGhl9IsSslNf3r2DO+1/tPGYPuB8MwF9UA+OHT6tAQT9WgqLq2/yKUuI5yHqlyix
TJYaRseKzNisZkaKSlDbL8iSoBecHd27Rt2QUwIUZxcWWkam4OUapO6aVLpc27d3x0EFKNkrYddN
HSeVZGvURivmUstUAVgZxPgN4Qkt3LQXqgJl3SyxGq7McgPtAT1X0LtW+WcacO4kTCbmmBslqZu4
AepJaN770oM1vvJc0GlibF07+D8sE8GQ07JvLQcASS1r6tHj4U7BpPmrgZVHZPGU6P+zY7bvAYD0
45JpKmn8MSYWFjZa789Pr5igINoohwHw4egYgU0+gjQB/Cehyv5NWhSsFqKn97WEpErmX9mkZQ6X
2WFf4lg1bx0NgE22eI3sjLthg0BQ+hk3UEK+4iI5ja8A9DeDfRqYkmIuP1OWoYJjgzSckEIrKuXO
hppG67Y627e74gTx/mM2nkH7H2QJEdMWWkU7N62FP+CRV+0v+YRn7FPMJltwELpvbJ8BJDCcjQms
f1pHcRnOEQVVBOXXYR7H/vp6vWUWQRuiNickjl38VFQRGp3mrrz7poGDGHVJSxR6vJZAei4dsHAe
B3+hqfhkNDoz6couwDw2b53wjEdRCPXfVYXxIsKObOys1IpPD6A4TRAx/ls4iPU55fFhI77WG4TQ
AXnsIiWKmCdj+DOflGHhsZx8twARTkvLWqhbkExbdEcCuDCUCBwQ5E7XBOyI9yrmAEwQpn02G31W
k+KqUmr7xmlRKe4C0GlNvKmjvfWJIxzRiEQIUgxm5fJQGy3Nh0dU46Elkbo2xXpk3NtCHeUn/XvZ
JSzmmU1oq71dLGKH47kukbOMrDp28C7RYojBLAjJwew3Y3CtON0Xhgr1Q8+HBrLBhSPPr/n4ljRU
nlNWurqFTmEh5ZseE4b6CRZpOJAZjwo+TKKEU9jRwaYGVz0Tr9uVPprowdsjvpsNDaqW2RWPIDay
Vb6wGhlt4+tUUpbtr3CKHZVzoKpS+2nYhDhPXDUy23JfXPa9qaN/fv8ca+uYRFIZSeiTKNwrjY+F
bmxvto418JQi2popn0VCtC4GkyqwCh0PAQNc3o9IZN9BaBnOjxOMUxJPYg/V4pbvs0S6fMDx8OOu
XWX9zZ4uK3CZXOoOlC9bZwJRZo4k/CfXlWGlGER+mMGMgs6DSv8qmoaiLVM4pji8PhdSxeoR5cP+
zLVbyidpcECZ5TDZ9hJAqvZz4mlhgGUGPKoKh9tB8RAAmjyGBHGZZ1sjn+le4lUtcEt1JpU7K4px
YScKrSeoJtSFoXE2b0vsZf8IwJqpHnsSDh8cIB6NCWc6CVxQ7Zd8iT+2ObRafwA7MaZ0kVvHipha
/clxUfK0BbX/yiE2lsh19ksDpvV6mloN7UQ1ss+pTEla6/++J0ybD47YqNisaE5ok8hLzkJTEjbD
SLKQp5UhTCEdS2audn7fo2HlSZje0Pq9jYfg45q6xQ+ZIkqxdKBEN4rjVExDgcQ8rqPvxSdWYJhI
sLQ3bpWh9w1TK7klQfJrULird/BYma98EXV3vJXz7qeVMCBeaxiLfs3msZGXhoBkRCfgnL65ascb
A3+dOp+cULRfLUR0r5Di4IUjlP/DW8rd+vceUXWzSlm2x4HS308oKwbwGw5GYjHdZC+AhfPNzEQR
fPPxQRZFUws6acqoJstp/mDIVqijwNbQRh69O/oFXHJ120Hxu9CethIk69C6GqvpPPQeDTvZsDQY
xgFotNWDDA4Xb9uc6Mf0pXIQCFmjcINl1wAWRL8jhr2CRj5rxpMnDM9qPxgNGXycsUaNbI5yIhQd
QdPphQJaLAAEMGjShid83jyizrcch/QndBt23hsO1QjFFtUq9GQmhWg7PCl1E8zvoB6r9J2YoKco
qWdP/1odAHM2FvZIE9tHLCpKe21lKn+hReaW3gKqTCcx3z3xqhxmyY7piS9zf/cPNewchdCk7YsI
8ZBtoS4u0e0oCpZP+P7H8bJi6TybcKa74XDCB5od/dPdHCJLnIuYcrJ7lzem8sk3lHORk91bpGWg
uCQsnpglG1uAOaFxpHzXVgXv1X8MOY+3u+iuHtblcob7GTBkevo5Xx1PEkO8e7yQsM6y6yoQWnwD
9Epe2FDnmQm7/j7NNfMrYAQ2cwefE5CfCJFYcJm/DTs2WVLJbbPDHynz/u35lOx7GBYahOVqgd37
zygwR5t/R3xDVYH/2edGq8ibGpep/npgJQlSHq4SwIXh+l1QDJDEXbHXH1ciH5qRA6tG8kamwd5x
udHV58ayLSlkjVmp0WXawBb8RvaYkVsx3i4vkgpfAq+tkBaKYWwoPSFExiKDh21vSwPXkLZrcLZi
egPhCBJ9yDslbF5kElGRt69sYN9OCtO1SlL3QQ/inz5+9NRHae/3aRxCAY+bOpDQcgbGFr6ZT+am
tBmovBi6r6DJ62NcCdVdgdvUeIC+G6HB25657WpTWHlzcorTDQyO0Fzr4TAniWOABpVNJe5BoPTt
i7Dxl2WEJ21LjAFWC4nuy7kF7GmsI9LeW7s7EjooFe+/gbzU+dl1ZkpfM9DGlvPMM7Q2VxJOI0Ow
WFihQDvkK6TE7m8yYapgqm4OX6uERp8Swm3wVV5WEpYFJuh80VcKwBO5IiRaqpJ6HfvsoeDJbNHD
L4fa78ZVhBzJtavxfcrWZxWpZFkvCK6WCZy8sEygtmPrOgYas+lTB5ivfB7lx484RPupCzbVcGdu
dFSbI9MFOpGIMbT7Tx4K2nyNm++oBs7evqUDC7i/drI2feZKfgtJ53/szESnQJedsi0HlUiwAf98
mcpQLnQkhm/E8TbZJHCScJ36AYYI5IpAwKvxLqe7r7VcF3m8MckVOxBZSuKBbuzwS+ln7979ppD/
pZRGDcrN+5diWZWSko5O+/z6pYpri4fNMxn+VT+E4cslMqMcFK4sI7+ysGgc5sct6aDAOyGrxzdz
/xpKTHAfiKaS2zHQjvUnsmcESpaMaZTOl4XJjEj05hXCQtYW2lLZb7eUc+bPEjENxs8fqJWIk4Qb
QWy/6CgzbEet77A85eX8rcaa0OXc3UqzXPzea6TC/X2h5V81x/JrfE4TJR+8DcrypCJ3ocQHsnVi
dsyBrDW69GpmPusIIlPOshHU4G9w3eO5EdhWf5k08+yv5FTSMTVBcIka8QYvhkvHmvqVdnpOX35X
7+U0vyFgRggsvsA1mZV3j4WV0v7HaqT7Ck8nAFXWh0XIJlA5Rgp/UKJ1ZXhyaM8KO2f4o0mwX5h2
DbCwfyd5pTC3n+6eq5kkbXB/nLnNryARt4R/1b8SWdFZbPLOeqWPLRx34pNlZvkp1i6LG+9JqmPt
O/3Ty1N9g5/vH5+49Y37IAF/xb5Yk3eKHOpVqYiOB2mJ1oJyfopauX0C/8QjYdsxFnLIzYtt6m6B
MnPC3GI8z1OrUBxQqRSCIS1cgdFo7VQkJMevpkxG/xYqVOBLinYSd2iSXeewCUFHnJ0tZfiS+MOk
/GBaB4jwo3qWNJvKfZ9KESXnIdJdmumDodWLf7O5W7NIjU60k3VLMJA+lPRcdOuEt6aMP4mxTpdP
WPVG63iXlIiBmA2OjuFSTJUZtVUAS+t/5YlPLY3N6ocsqvVLJZXPuq3xLru+UwXLBervUxmMAX11
h1f+6k0J4FSJVktk1+1HNk2Q8LxHOrf3QdASjGZCiH+t58aKuy0hA+2wM9eTZ2J2zAHr3muRG9mD
i3X6iThx/L9iXZs1gvMyBDzgCkghG/dqNTmTWjAjNnL1093aG7rEX7rYDggpivJX4YWyW6BrPvMQ
e6mGfoiTKdm0C/695Bm3cCzCFsp5VSf7+xRoyFhtMomeAKwx/SP/IV2QvOMIi4rxqGEiwY3mRstV
VTVfIJrxEsp39y7yOO21FTOpZmEifdcdnNEmr2byswC+eXIdQQuh32GXB0U7rgWzhuCR42YczAs1
10/Gu8eAfJRVYxfWtf1rXzKOtti8wateCjKXI9wRwuReRuPEsrFxiiSiMENm/vHZqhQZ/ldb9vw8
qVQapgLrjzKLVjSy75GRAtKUQyr63yIleLRGtuw0GLlSjgW4rHxZz7rEDxeWJ0fLnSY0xF2gWl/Z
x5PWQmznTkaea+ueVp+5+SkZJuoi9WiLrC30cIpI2jrhJqBwOmWH2G0L0kZGbSnLgMgAinBO4a5n
pFO/Har9pwR5xXyQiV87B22m33kBJfL41oKCBL+p4mB7sBqXWC2QcgTx7YZpNezGvVvu0tyXhIN4
jSmO2PHO8dYKahWcxT1f7I1om5tS2Z70MiHfjdF+a5c2e2CSBIGtNngmTjiYW1n6+iiDt3k6XjFT
seQf8Y1wJ9VjS/vFI0iGd87ba8FxaNhJzBWvMLkph0v/+ZzQQnxsQm2x8/l9AZ1JGvImnORDHWS6
Oz2eA5i9z+uRBHcYy/DwNxWk+2oiWF9KX0UOqz5UdW+ozYGjbZ6+qfu3EIoRRZdu4nOgIIKO5FyU
QJSzF/aiPgd6T3doXMIleH13jyCrU4Kbvvh6bp+UtO8a3wEpoQSWWAOjGxCVYuargg/HAWjxX3/f
mI4uuHx8M+u0SIjZWSAEcwr4SkXnXVibeHq5YsB0E0N05gE3Rvluyfj3DrgRAJWTEaPcWxBwkz40
XypV1BZG0DWTXeZJU/OOlg/RHkpP68SMq8b2K7gY9BH3pIWCbKlRp5Jjt6gad3lt3js39bvSDphE
FPls0wfkvhXj7BXOaMnIyAKUmVlJw52kPsMRVzWXY4SZ06vAY9CIB4RjY4j5/2w/FUmB5BsPC5fa
yznJ5/0hZrn1xIcCnQXdYrcdjV+dLhCO/veW3XKhSRlMgn7RXirNEw9ky27NZuCNOraXex1i/mFU
3jLqIhIfW+EWQ8St4htOmFIjByrXNx2K6W9sXvpc5yWlN11k1KEGO6JAwmUlxtvgFN7RR944uZvy
iKSshZxOkw57F+EJQSqNF6a9Q2Th6iu6Da8bez/AmifVGAQXHUrbj0TtDGHXdiPqvKDdh1EMQRGH
U+fVWBSyYW1o8fLQgj3PqF2ZvfBmoJBEbydlnKMESe9DgISDb8yNoNeHjEfSh4N8Ht13vkqDwyUS
cHT70WVy2rEhiFumls/+wV05Y7sHh7T5pqoFbb2t68eXqgSD68xps63XePTPwunsDpYGvhxGy7G8
qVNVg40oQTxfERmvVT0mnxeoKPkE8iFpqDcHw79yMi1vKvkNA+n0LQmOqPAJTwqKSqPtIVF4MNO/
h5EGAV4jzcgw0VfPFiSKwGUAsWr9QEal1Mhi3rnk3hUENB60Uz+umhl25KJrQdVflStmTmgSYveC
EV6sLjLYuect9oVV107j0qU+H21lhmC50RxMREe/01HrhnrfyMRwl914a/Vq5Wh8w6dWlyjYazgw
LdDyuRTvI/mNpBZkRrA0pG9kDmjXPRfJWUQMiyUpc7LH/3YmeieOxWfdR/t9anB1k8NxXhpnr50E
p9YBP8lEqTa4ms5VxmmeOPepPC7lHgKSuNNQu5RQ1Q/mNP68fm3vTnFzI9ZlzD5P1rLxv2250h8g
g4OP8gtNTVrmNARgaX7LE20LL4tFQRwDfCUFrU7i37rkyDyF2YtKoqzq+3LBPy0tMq0YStsqsUn+
9yBX2MVYa9yeKdO5zGr+vPkAh9ZD9i90FEJiGO9BX5UzeRimk0CP/q3K7mxxuqlv45KhOF+2Ug5t
CcvTij3gk615gyqAEAUKWO7GVK9gMz6s+pMn4ZRP8Z6sQo1ti48cfu8CwVEWsHfT37zHh9gsN0r2
v1yH9l6/JZX+AEitHzsWtQjAOAG2X4AFYc5VzRTEQczYTVQwOuOrqWUNKFlSLs8cQ/tpy8qgtnzn
D6sVV9E0uL7evSiyhOQB0Jp9UyoXkRS8czBZbzy3w0qrKQ+ZAMBMRPMJP6PYVuINIrMGHyN2GnaZ
8JfI0k9ngphr80Rno6Rwbn+JevLv8YV30TQk0aqSgN+lg5/xQhbH2jY7E2XOIQuON0NA2j0Os3pV
aadOpGnMv2+aWFaEh6ujE1JeVHx2t0ADbMpE8viP4szbIYYYWMSE/Nck8iXyPfmbMmdtxLY43jCo
bffM5tmrBf6Aya4JAaiXFity4Isv5NsUeYDSyJmvHJ0MoGaxQLZZd0INHvfPEojph4pgfPhgruy7
Bi4GmIExcY5hIWAV0kwnyH1EhAP1YpxCNC2cDFnpgvAYkIngt2TIZSrdLfGXCtgK2Lng5TuZlC9G
o4DsIfh1Ntkh/FTt74E6ylT4rpk4DXIIVyQU8HA6CqkbM7pHhUPsDV9NhUYRslDcNpD0d//rwM1r
dUDQJBfBopaPpeNgZ0AzUl1coEhmiqcNHqH29sNdF1ffvqYJaWOohV9HTnLFuIO3KUh4ewg8Mjt3
TrwyOcUyPHpKb3KlwXNimZPkKChrE2yQV2UvEQfcCLteyoGThNtOIymLle5xP7aDkxvy2D2ELKTG
n28Zuj0iCyqZgWSmA2tthNJ6J/saLUkIs1nD76rMZJ+fjjRxoEkK4cm7m05gXTpb3aj3n3ygDUq6
ixRTh+gSXzFlB6jsmuIFEQFy5mHs4t7o/+Idbmqd1UqJa7Nm0UTiWBUzqd2d5eKfB205efzDJ+DA
vwD+7Qgkv7Rp4vptbylRViC8rxINIsFTpzTaCKYPY9V+9OKH3iegWFizko/ad8WaqQel56v3YTu2
392gq9EzwiImSZgL8iqrDCoFho0EGGWLwSVc8ksBOjutlTyNZYj7PuwDm3TF+BPIlTE1WvCZXtPk
0f+EMCu4MTIDxMnVQZUrPkzt2nzyHhIrDLECD7zvTydZSESTl7+4UnuIDmaXkbIKzOwOaqUrcpa3
NPg4Jnk79+lLWcSYiCvcjxLm26UMmQxYRSdsBPOJc91/YP4Iz/M3FZNFyUVngTJBLjwbqdPM1pSU
uhVRI5v6yWBb9vnGkukUCl16u9p5PhZdKI5RRK73g2dPEZONzUUT14C4Uwvm8lJHQUfH7vIWNBLv
QiCUQTYQLboVTCaSdK7vh22fqlf8nCNPFljMil6LpRhwpStO7riMUrBV05E37zV+NlhmsSQNjc8u
zpAEpFY5g8CNpxwTYcD2anCV7LaQltLZyzR52HM9m7oHV/cvfjETbCOK4TeKgM/tNzr0I25tP6eX
nkhFYMzvDYO36RdNt5+C4j1vRmaeuWKxXQ8MBAtc8n7GTpnJzfAjZcDcE/KzzDu3q29XmRUbSLLN
F/1RU08fuyXfa3BKe6JGcomRG+k+AznUTAdkB9kG7nrysbx+ErYEn9Tt3GM4sZPmL6ua3YgV+i4F
5cpISbgkZ06lInlaGIBAwjsJOPVsfCtEVO8/moPCb8CsXto0vJT+I8NeDLZivnJqzDzNalif+4lK
VU1bOZZ329gQcxzutYCab55tJt276gOV0hRO/TH5n7ouz/zLhClqxBKNUzwX/rZSib9J+olrNSmq
rkwqGAYz4ZcRX/nVtBScIsd4ZrFDINh9QARPcgakkyGszH+bSk8ESA3sz/80T4N9QGoMXre0FKfR
sHeGuLL7/N5X+RkHhI23Gl0nn5x8PoIXceogrzJ05HRmXy9FuwKLX9MTY5odvJYthQP1DaiSGlsR
4pinrz7BbiIxvC++CgF8LXrYeI3MWq2TOFObaSUU0VUZ1uH86imYC6ZPaDWC5BbJIR9nhDHTVGe/
LHOprI62FhBoCTbXzKmSp4KYdS8jq8e4v59hgm1Ss/g2EU8VbetjYThEzrrTLUMV4SQqdAIllIvO
ajSGHwLCpvQ5S0NV/MiDdzVJuNU5OgV32yx95x4RzOwDR3Hy/1XagdP3iSFG9oW3MDG1sbTDbMFR
Xoj1FmaszHBZXvm2iZDNQUasIs/fM4lUHwoEeBrqthJpXS9wOz2pMtVs4aao6W6gx0ZZyc+pRQBb
NXqQzaowVoiOJSqmufOhZ7rSiudgfXnLzbHAx1TYnF59hIiWUzwUNpFn79NaWwwUCW1/SdytVMIz
HrIhGeqx8N7OGV4iwCeCfZh76W0ID574CzUe45qMdG9w/lQvpM8aoLvj3NfHD0L6aT3iQRY4HZe8
FGae+qPkanWeM3O/2wcUYZ0cRmgnhERmfJY/nkIt4k2NgDmzw+IgJIGxPo5+1yS0p45qb2NmK8qs
k40GZwLcZMoevqKMqnl6H8iSmqI4HYPu1Qq4X0IKDQW9/kNvVOr3FAQBqJKFzySKKPCFhXgADgCw
I5lYlE6MZ/ls0OCCQUVOnXmu+d95NZVjc7WQruZzNyEiVn3JUe2L4kzvw+QS7e6pvvTNmaWNRYnG
KURKGzuQtQ20TlolrjFi9yuTP+Ivm1LlCUzAgDFEoHV86fWbLE0bUFMMtpK+uAUtVYHNZ9iyoJla
//CRrNhZHr/OEUs2RRtrWEfyTouqe5vLcMnRaZ2gIpYA5Z5ssVytSTiW4kw3ImiYERdM1l0uP7Ob
kM3v5QsNwdaSs4xjBrOW+zIUEISYiiwZZjjU1Rz51KXUQcIvv7+rg5K2OyMrIFwS662QcQfYT58v
FPvf0IGoIll64Cs+ZaQ+2d+yz7h5qRkobBLE6tirjC169xAg3cYzPFvy/dBV1jfVCNwlgppAgkc6
2D3YNTWeTWynn3Ct0Q57isdCeU7cfV7NYpNqaSbHQY3UOwOOhPIu7Qcq353RP72Z0S3KQ0DVbC75
I3ZrmBQYXeGhR21/ZI+jqqaaEdwpkZVfwlzOgVd2eSvHRxLeNuESfYf1IvVLey/e88K95MDyc/UT
7wVJaniwzTsUSMHhEDdEezY4YdNKQlCFQdRxqRkSYPi1DbaGcqelKg4nhKPmbnBT13sdQX6ZO2iT
8n/PUiibIfkJq92reoqt6WuiR1tf/1pVn3KqiNhHJp2SUrb5DUcgZSptqte0ptHFI55URVRJa5G3
jPGfz+5sLV3wxAz8pVb3F5Rf4LTohl+LSyxT17MfcZmRK5WnPegA0xb7G8RNtNr3JSqZJ7MIc6HK
GjeFcujT5CpoaFckUahbytLishaWEEyhrkvW+ha4XaJioeAOjHdxwATd/u+JZroVRLsCwOw1SYlo
dFkvb3aVl/Pc2Ezm4C/rJW68AEvNcLMic23nX4fGgiABqK80Tg33EPBeprwj/Zt2g3J0z08i6f8U
+fKKQbvMy7VHYGcHiMktG1qzdKon7itknOUhtoMDBQqeY99xgQMldO0+w5ZGFXuKk61CYc0ewfp0
nK9YEaEWvRJDcg5Ob6icZ8cgvYkmLw77KVc9jNREtA14MmX3mOyEqTPcYSPlU+yM2wdlycupWuwK
j0Bo9K8yzhfxo4o/ANmfnAXXMwiJOMn8W9flcgZMbVHFhRzsu6KKNEnTCybXw1niMavu5jnWv3wh
FfdE0T4a2o6d0OUBuesWy/cKq5Rvb5rCl7ldrRGLLVJTQ9PT87TtHwXiF/B/cXRNKOWERcDbpdIu
P5NREokgSJHjlUZtVuELWZdf9EOxEYUjF+toPmV3rUoCq/i+NbsesXgqNO7otHOJ+2y+ks9f3pi4
zoo//IOzHR+BC+nhS7+GqONKOiH3aAeLwnAYXGmPtrT2AkapEiNYcjsSlbizfeW6aBUCXZvKpk5Z
aiAZ5yiLowx6at/otDl9NP3hiu/SB84/maIeK2P5oq5dyeSH7s9egwvu1c2atyTffzpT+DR6+pDy
udierx789GuR5TZ2a/6QVxD0v2v3zazJT3GIYTxOYerJRJarljAE47jAfHmJTF1aj9bhw1CSB4Yg
Is+OwlJ+KAAhAGv9bwyOHvI+qazWA+voGdDx/1vHQRJY/2ZIjl8gf1b+jDUn6i+tCCdvGoD53mQm
7WV6jn8Bkc4DGwoddnYXRNJMYfOHm0dpa7Vx9cp58Hn9jiB5VJwloAbnYUrlfXm64qW3l1cdwUnt
4bCXEbVHbtM6KUMDDDRpdHlkZTKj1fbpAxpPcSqprzUult2jr4v4kIIstrdSKg9gqdBwaySLIYOb
SknQoug4mhIronLm8yPoVDRBJtWJ88tg/YjVYasA/22aiAmvWzoiS4dx0E3acNt5Bj288ytf6Mlq
rakbs2BVjZm2xzezyK1CnEZDa2yLycQU8uOzDahY4YNs7nwH+ynV6KMYwj1VWFve532piKbY5Sqi
1zXCPp0oc2k06SJdMqopQb1iGcKrii8cYAeeushwQxmT953gD0q4HlGwYxI/Vnwy9nR2DRrFYePP
50eaNq+wdZyk5j1m2MoHLZLSOWSRm2g3/4SiyPEzM0f8l9BVqkH1SCjS1MLEdmcizj9tPXB4Y6fq
jVboJIAvyNgDXjJQND107uGnMNg7qzCFVDbbBKpY3ENs/WhsYRd4w0MNZi0Bmeh8v/HmciifTrFp
T63FMViEVx1JkVPKyAFIJfeVlNRAnbV3GDrlE527Snn3DqVnN9DIoFI4JCEWniD7lzsUBDSvVuRh
z92daquTcUyxqiKBFmkc2H/u1uP8AHsAQSUeyTj2xJUNADwuc32ja0oZTHOFgA5eRm3Z3adK8Yci
qTsrejPXjB+oyjCq+qXwlT0YpeS3fGkkecJwlbmnfs+nFcl2aJri1KiNTkJ2CRrwpCJ+CLnsQZsR
0FV4rXUgA214aL84QDkRB1JYkLBv0H+E+LfYauMJOJ0PBQGV8fwulmAkalJnRU8XqOFO/BFmZCFB
YT4ORmv4MWVrEZNbw20rb9VKxzYMDvjuERCb3b/N2EPSNxu2gZuLMAI3cwergMxkNd/cMuBP1HmY
fqGqBE5YF6uVCgfqVHt3lTH7KoTi6CRVF1rEjMmn5DFVlBPi7glDUugSlAOIMLwU2XYDiKla7AuA
e3QlNxtgWwAuCeqcuvcXi2iwQBqmNsnqy9dtTzf+YInaV7zzGDxqKsFQDvLX14h00pPAQBMgygaT
704CiAuDpU+Zb/qdOUSZXeh6oy0/LqfB6vHcv9XXtnK/983473RxwiHzGsLC/e1ZukLzhMEY83k6
sxtyOPLI9ZGzhf2N/3ck1tmBMqqrUS2z23zo2PHv3OZzOIv0aS29N4/GcwW55TCpIaBzaLwJQs90
rf7t633uWHtl7u/nDzXo4kTLqHD+kOAFLXbHioU24zp7r5NbzyXgdlKBVfMBSdyO5e1TANYZ34yB
ay1qGxfZ/SZnIKCiBDc2xgVwcy1TkZQEryNG4PQkxFlXJi7LaW8JihpgVvcn/ZqFQ5x3vM3NmaXl
H/K9Yrc1JetMgzcc5NAGZhlaJtNh/1Cq1XOlTwhyRJmiG9NFUpxnpDg1GhvXT3pR+Hj5Jc20i9R7
FuOC7BAIMsAIGGsDzFS4MsQ2+aTVYJUsSjb4zPWiedQpDL5izzhC7r0G6ZG7S/4SqdL0W4j49Xfh
IFMPTE55dT8Xq2aE10ynCcE4tV1sufa/6bUy2o1m2D9USjhte+jJeQUUrY5J3vRx72+WLfxJbukn
ohNrNkzODDukPQcD+8i++EDotX1EKpUN9OToaofBYixdLgFUY0ihH7mZqGHyikZQYgbwWryTXVYm
KXAhHwYBlkDlCCNb+1i50EcZkQ67AweHllhXKLp6O7sIoh1NgVsgDqDjV6bbQKk8iBIDnC4A1hT8
UTrkxSa/XYNrV6rlfg3Vsmg7ea/zpqRKB5343ZVqfw8G80ESPjNy59PzgHuvXsFygO3sGGEms4KR
2w8WZLYR1/oo1uEK2826wOFt5BsRF9LW0axVcbdvVhkq4Sf10S09sBloyxgRwtcdEaViwwODQhxP
43qx3XADAh76BxgCBL49LL+Pz5UgUO2k97kx/WrBC93fFjvcOVjsym3qZBZCwXFLDJVcmBgB7IYG
yNdhLaX2sEI62wp/aaMHVVNLzY6LvGLWx+nn5NscQXc7GecfcQQ3B0tC/Gs0zxn2MAPmNat1BWDM
cEgZyGoizMUEHFCeUZJw58EmnQFs3zy0Idy/zgFPL83QrH8rePS1F9av8LLER5rk/evZ64LecxBj
kn0Amj+YuaEXwpmsAVGeIiCtyBZyIfl2ojQ3LI+Ce084mrXQR/293f5+oo5IEBiFtccMTEITx+gX
LrXNi7A9+XWYHaLSQ96M8N3T+aE2j6hTRIWWIjCO7B4aeZJV2JBLaaxrFPS9Vo13pOImx6YQfXK+
tuXOIC9J4nBTzv/sWCjzuOq7O1GQ3dEAN+KXAhelaB0vXdnrqymqObUI32OUO8xRC2eme3KBAP9P
OXuj1LlZgP4o4H0HQYk1fH0Lb2quH/hyS6aX/yRcK3iDND+RompJh8rrxEseZ/vIdueAlqBqxReW
rcUnGB6CzMcqLVCdaxn+8reMExwPvosM7Nhawjq1VWJ5n/v1xT1h5j+i02D9XwP8Zdt/mtE5OiHc
ag5jnKoc/vF1fAxL7EWBbctMd4ELpgsIOqwq/ByU8oVFQrACaud+Xg0/YfWUROZk6O5CVG6tK5Bz
DMGGOYbt6hGDt7bGfD6V+bqOxc5pia7kBHDECiPdzhc70pa4W6hxw+piKe53XV9Y6J5qk9qET65r
yb7n0iCEmVFeHVugYNwySNfsNRGi+Abzwo4Rf/uoT5P8sHm3MLYIaLV2P+Wr9VHmsDK6JGHdU7v4
Z5/T68zcAmWMcZbthqwhtzwsM+1+Sk9YHGGLfk+wPpg2dJqCa+sJX8Dy1wX7EMqDutK6tRbFgztp
r9rrhlTHV9bV/oNIghNklMg0gth+ITqBeXrtz8C8sV0qM6MfCDik4nTYnbILrdJ5VkMYhkBM8BDa
9AsNHdR15CqqatYaeEedffqKIeIM7ceCUZfaapEORq23mTo0XCiLQNK01a1Ja+iE6mZOwhIDPKoY
bxKvQXzf/vpy8mYCDAZ9OjjH96bg0Nd7sBfEP3P2rAUqO2w7fKhrKvR+aYsol7sqP8DKoovVF018
0VVfPDiNCthF2hHjaDntr24L/VZvXLqbUM4mybTvp1WEWx/0aBEWfBKZAt9mIlRaw7TpBK5S0b0W
uHoe5cjQLgmjERhv5cTzZjEmI4pHgVCDzSTWFTQcQOZMFmTzZWp7pZblK4kxEDsY6YIgQUeaRQlg
vvc/NPOdUWp0JQ1ucfIzF9zXtNmnpwRnTQzmSV7w0BDLVHITUmP4ot9mNfTJgrtsHPfHiuO7f/w/
Ad1NGvatxc+3Ka66e63x5KU7Tz6AuTECXNLGJ468yuqt1mbeHKgbvXEtLsIesVieY9jDHmDz20pT
Jihef8Q+W+Et3QN+0FyldjkbDx6t2Cl53g0rE/eY6dSABDHFlgIGLNJMQ7zEOlczJzqXCteYMNEV
e/M0PcBtNZX67NR/SPsoV71mNIcUVJBSBhQ1Moc6z3NbrGne9DaSGmwNPdFbAEyTQZQaBowzoOqN
KxzkWJfrGV5g6FlWBjjrPlGA+hZHf+ysyUkDaJS6A/ylGo4Fu/d2ZYVtxhcWPI0Kc1+VvwjJCVSH
B+rQ3rZqaZl4JRo1tZa9NPbK7mO7VpNpseWHyHeUES/WEiuGA2kg5fIw59aS6oZQNxvnU3EFse+Z
p98jqpivyDapXwpU4HfkPZ3GnEM+DcKYwwXnBQrJ2ys7T/8GEOJMqEC9Q7qcvS1Xu3Pa/2roEUl2
vm8ugeNBYxlAEEv0Yc+q4cOMsa9V8nrY3Vg/NqlYyOTTXvBhtwVo0Aoq8rcf/6pQPq2WC8lGrxhX
spAdOMhRfTeU8v1iLTCM7mq0pJY6092WiI5rWJpF9kKKhDLjPm6Yu8nFXCgBr8pBSw60kuVc0/I5
PuD/5ewwaf1OeT4FDeJyDif1rRJPfQvVJv44bTNRsz6sVytYX/yFP3yMbQvJnBSO5eVkiMYkWHD4
IxfrQOmVOzev+LzLnI9l0+Vj/e0uiW8UXB2btvOh08qIaIzg4ZoD/sKNT9fqHDYhFNLT2ZAkG3oC
SznhqEKOsagD1YHKq7sfGLjynA6q5xcpACmt6KTgdpNz9y3ovR9pxsariUwT70GLUhUDJRgY9Fj0
tDUt0YSLBj2iy10iolPGyV3ck2uJUvfZkJ+mBLWvANmf+1I0omc2xQrj04jSMMs0+mnIqQYKVGhC
4C2k9JyG6/vNZMTxKAO5LnAoZQUAmVeZy4T697A6vlJ5iJthZI6dXMojT75fDZ3hK/afIRRvJHd7
W1jqc/hNqiZBqjkhO3Cwrn9nuj3Z9undM9avwjSkzul/oM8pRtiMut8FfXzSrrO5pwoQabmKRRgp
zTFTZ6tEN3Qb/xGJGdca9IbIcVnJ4BKH5MLNaAlY26lctjZ4dNEW49O0LHKcgxNrkTPBi1kAPEuO
mE9uYaV3uMs3cfyCNcmAGxeCvACpSG9OLzLbAKjN4SoCRPTjoco5JM3BxzeB0vRXvsen+/cb/kyL
PO3SZSaPcw7bwHfQhhufJlOUP1MUEYUGt2SdreZ+VJa5/txpegKMYpVIEJ++VrYCH+fgMzNRT8X/
HUukf3GYSfHU8E9XHGVTHpWGVXNOhXNGxol+Xlbpni2bhURPDfUxAMl8yq9M7Quuk8SBYY98qzzS
Se9A/ZAD3a3vY4rYQ2IxjYt8op3KsvdQ2NMGyzNa40UpVPbroioeXOFPUbcsV9s30Rs4Ogmhw/Pu
N9KkT+5MSw2LFOVCIs78UWcqcurtVM/pjRCeRcjhcSak2MomJWK/iT7AUGNGa6LBaI2LSm1iU0Eb
6A6nitFkegOJ3TXHBYthggecL8sMOM9A7ItYlwbv866AHnL+BewCUx6YM/BVctJYF+y1I+9r2EfR
Z8xzxb+PNBjh+kcyrvknMS/n5xQK1hkACGFBQQDvJPVLIpfQrbBoUHBPAOyNjGwHKXS1xW88Hu6t
7XaaRUjcG3qXzN2XYU3/YLSZjpJUeuCT65KxTcaKx/9bD55U7UPQQSpgQ38klPFwxAC3o4Ty/V02
7PvtslFPHqENNPXCjg22TlEPuTnyNtTgP6k+i9/+OA2G1S/1WKLxIu/+43i+jNbnLqqnD4CYp+Av
YjmLXnvbuSp3q7a5dLe20xZqWcM5xmrHGfE1hrXJIQJVDXxmbDDBKA785gFgMYfZ98kE0hClk/Hr
RLaWB+OO++frovfyn1HMBGL9/AFarbEV/WG/tOZYW/yKSsT6KTtMMD2k+Da1chwVO+Sb6Mghkplt
fUk2gw/aOKwKd+pMBI884FW4OchW+6ewXSodMVLl/yybTCTosbK0DWP7wp5sH/9KwzEMc4yMKAqz
xDpbOGKcjL/5Ft2/NIuZsPSD8kDS3suXA/1l3u5SFUcFwojyAZBbZ+sIyeWmqHrd3neTnheD9w4w
MgT5ixBa40kO0oGpnNWNguYjQ3b5wrZhdjmd1YL5kEyAqFAJK91dFHBV0t+WaEo2fGYNyi2tqS/T
J++QFg+cjANIGdUskC2J0OTwOUA1B6EzxxUOCjBSPrLSk5dcDrmP9h9fOha4EC742ubdzkrySE8k
JVYp0qPsYksdHVdTAblL7uaEQJBDGEO1OiCGXe01cyd+LRsCpncVCwM8zt1gTzNR2hUGL/kW+F+Z
QFFRQACROdOPvimlRB/SqOHpBWxXEdK3N9oTpBv0lfvyz+K59M/iAzdguM6RVpaFC78b2ai7QauB
yIy05dzgIpLY0cEqwo5pobtJWzLt82FcK7RfcS8JBNEq12IVz+xXa5r8PrnJoeK88BEiD1A4Ahsd
fu6BUxsbYTIytkCjbmZa/VnNgcPp40kr3PHLrSuYK5ueUThZm1e+7zdcg6q7e2W1QdJ12UTvhEtg
xqR8Saebl9nY2kLfQKLjBjsL0Ey+LLivOd1GzNdB4FsH4xTx4VrerI7C2hnz4cciYkWJhTZBrC9G
T75KhvXfmaCKPNgMQdZK3vj9mImQzps6f5AIvBjTfTAEo1igvzVDY7seMzWzdD3eXsBMtxjmNeif
JGj95Dqm0eBEo0GDQ7QOvoIQ/965gQa6WtJTNGp0Sj9qKTFH8bMkVv1nXprNUY8489iPIJB1WXoD
01KhJQPe6evsWwrIAf0W5J1BvAYojC4+RXysb7QYwWtvF9Ff9JT9ZwzVGuCvRpcTCUAvayhKhrwV
vkX0wy9ZDWI4lhN2LHfwcpy2oFsvCZt4hHWAB2RpMJ+vBSzS46MPOCnpXzdr5ebU6kkjbiY66Q2Y
I4kYj0r/rj6UR0DUPmB1Zx7Ledqwg1TPlY+grZ6/DLHJR2Pii3lMoDsajm53XwHYCYpnCqOK3JPv
nJCb4zz+flHroPCL/suAgCUyaSXhmZof2OadLx3xlMdkW5bJIiQSUZ8ynfPv4STpmg9U6j656rON
50EIqM2wPXZVJ+MQzd+L842k4lhJlVzbTy7wv+RyLODE0B0FcRBEejvhVL7RAeVxszEpmW81g4uG
pJod8YA00nO70DH/DKze7U3UvPoaLG23tlNXKnxGp6+MGJOoVp59BsL9rZm5uw4k55Mz9borDpgb
7du/sWDu53GSgfYa52f+Jnr5GXrXOKkAMuScAtpwka4Em12AM7SDhhhTNt3r9SsUTeb0nCJuNV64
g0mrxDPsWfpZL5Y61s0ywBuVReShgCYAiI2lcEg2IE+A2/vfSBlqmztvm1enSubPx/Dy0O26YchQ
Ww6ORlkVrGPHqfSs6Xf8kcELqPs+BDf7nc/lwblFlr3CihCsYGMkLLA3XdIzNsJKXhF4uyAautVw
dEmTgVhSUoeDk9PYKhnITsgaTRgHHh2Cdcw1HyEOgVEsEeTN/AOPioqnUzb1yDX3kvXA29BzjbrK
U4ps4vFGcT9261BVXWHInIe+bdf9gQsa3WBx2S1p765BkgLVM7teUlyLlHtSR9UyIpTMPhogQfX9
kd0IqVUiEo8CigQ2boj0XnldkE2grn1XVfryLt/3PuCBrAh6gagyfEtUXvTom2exZZKbaNxGIwuq
SNwWT3P0zNCpx5TbsKN30kzov6IfF2CJ1YVz2k5T/wI4K+eE0O9wiRTKA6+NnWM1uI4w0hE1cAAO
7XUN6pJeZHTVx8xqUgcvcktsyyIudDS1DmD7aiBNPmTtASr45ramlD/VcdDGZWBfuZKNQsmr/xzX
J8F93jrsAgL9lkrZ8lkOaM0mrDq/UKdvlhp8JvcQBP4eQosbz6FWMhKpSvi1CQNSD6UmCzTya8xn
8bHjh/Vls5M896axror3KTKDFbM6rblOvB+Uato8O1oCmMiHQr0T2LlGMNhSLY+CRARw0WtgOWa3
4Vh5QC1JUm/FU6JMtpwCxbRZ/U3bWT9mubyIVnEHa46wUtWs/VSO0pyEheLlFl63uRSg1nsz4fWN
EpSSDURnIGK8SK+Ct8S8A7mze2cd9YdvXVSFY7A2Z79JKfiMIjq+lJ4ccG2P90IIPy6r0Bsp8CRN
iq+cOxnQOpTmSN0+YFM7uVdMcOtaPb4RXAWyd1FPdfuChMT9xVWfwuRVfQbvJNQbNJNU9he+MSnF
C26BYBX4a1bue6ALDukgicfGQmVd78hp56qJsMYu8j783SOHaRfwXPu1u8zYBc8up2lkwPFAmeHn
sqQkpVQ6OeoBBbvM4NOOxLWMfqOQVPfmfGx5mSFQ4AlBBDv+bYG0TodLkEa0RsCIjSC6GTF5+ztW
yVQ7a6GZnnF1j8styX9n0gYxPkm5MzYwtyj8F1raWE9dSlrzBSJ7eJWTOZ+YweQjlVHBF8r26jhc
d9c3s72cK0uv+S2Ga6a6ue2PktOCEzQgYdFG1ZHmFEoXAT9tcbgy+TD8fa2cFyb9c5mWpITx5Pxn
E6MMgloNJ6zr9XUv8o104TcHHTobwi5nNsmjxkJhkWpUZvHvK9uYGJE79Ux7ThI8hoc71vyB6htF
BTA2IrwL2TmO3SfE0PSp9SKPSbxEBvTiuzvPzEQkpfWH2LvZcuxDfiJETZ1q1mF5gdqC63RiApuv
vPUTJ70KdbbxWgpY4zbf6nNUwXx7LQrb4lpISvsM8XZRPR/JPTe9Z34sJLfrjk69gEtcT/tdgUQg
aCMKLbAfJ12IPiX50ysLoaeHU0qy7+Ypkgao1X/ENPjnhGr18UMoex0PyVF8dLfVpke4M0Wj436w
wQhu9Xd80JOcHmgTCMRx7i9FyZFjhLP5ZhGqbFnplOHy1hyP7hB6cYev7UjNxYcavNujbv20OjMF
UIlne5HZ1z8KNiJYRjLh9AOOZ/B+brxxC/Li9PIVGgsy++tJgsPV3Ft7JW0/p0ppz9iGKvNu0h33
4/5EGHNbrvB+l8URCzMhL5moMw+pCtDJ0T4xJzPw+XcoRI/B9988MPXRvSB7zHyBGjVv5YsyPmvj
n+ADZ2Zwd1AP31735UPnjVd8ZeHWQr+DylmO7AsUTtoKsYQ3mc9IPlEhEAC7DSB9OYNgG+5BAEgU
QSTLFH09DvrXVsaGbDhtP/UzkvoovN74WA89qZooCWXpIlmbIdB0v+eWUv/LDc8IUQfCNgPAh+qf
cGGOXkJ66opRhCYqDI1yQf7QycVlnyY1YoaMxVgATbZo4AwHX7Hj5WAbvNZNOsCoktk2u2gwsNaE
GT/PmekHb3eA77TRdydUoYAxQbb23CDdWJC2zrPxe61F8Q2hOahDJ2sAcow16zoHu8gb5SrRMUH8
tjR2X3JJXY24CWhvQsAEbFvCaNZpgKKfnW5oucJZWjCJV7bni2BE9XikPM2FjQFZxgiN8FmJnIas
zzsC0TkjBgPtGr4KRySHMKA/p41k5RSTRHUNbIGNf09vorplZYebBuJ1EyQ0ay84YRCGcN2PicFX
P4mYTAnSm+UQSm1YsQAIW7lD09RdU9zgSBkXh1AV2enlD6AOzn8h9yzDp+WxA2+lPg/GgW/Q6rN4
+qlbR9fLTDUUtUerERl35kZ1F8uhYlfc9U0QbUIZDL14Bfler9yGzs14wH8fyauQspp2KTvTUu24
eP6azpIeDu0FYV8NC+eNz8NxejbAuyp+6Zj28wSMxeDRW/UmYF5cnh2dYc96egXxmQMfuWridKLZ
uSUqPfsafenXSnvNpkGd0oIUeCGv/8+yoRE0JkVhiYgOdDIH/Dh+sgwYp71IzUGseCph0LzGgh3A
s7gM1wdF3kXzKsY4aanhWCaRxePwq18/nhKXdvCX5pcoN3ZMYN09Z9rai1P+DXt5IDJ5yZqwT9mh
RdbeaXb2En/cMAxXXJJACOG4etiKh89jRkBdgGulec5ofFYFEANPJQqcALoSrApuVnLZpg8x6UDt
zT8esZqwpiiCBZcnItCJilgAluKA2LPtA5EqCW7PZ1PFkUafTBmQ5kNAAPQY9JbjLI7hkr295tI1
W9XNTOk/xWLK3+AR8fxRtjPVsj3IzDpHNJrYXwGbMEsQ3bnQUGiMJL0+ci01VN0MPMhK1zJMz74c
NaLFbi5J2FOu/zqBqKdAfRqdsMbyx/ydVfPvpDKSJxTi/Ax99HNIx3CC5xb6TgzM40P5Mr/5gXzu
ajVoV2EnCSgYomNts7NZGgl6ywIp8jeuxuvFrXDKKYGkElSrSetjcAbVFZrk1NXeg06XhFjjXLM2
5hLh1TdaFURnxSjDY0wMf3vJu/bS9HDR9ZU4jUMVIeDdP1tE0NHvrbv5BREcEGmIhkhdoW5n0wcb
Ox6/iMhhWcc5eAf4cxiNqD8hZTt+E+15DUv5jHVKjjApLPnGkurbjxqruXCG9AawJ59o2VTEu6LY
qdA4B6xG4SMNf5pMQrrh8ssjycakUafLnF2iwFrDB9thFoqYITBPr3tIJ+O7aY2JpwvJ4QyZcZkE
7t1jSv9o7CrDyIVXvNGfpGx3tbGL9RFmnHk5e8uw3c2Of4rGMKiCRDiVP03vffo5bJ+wcqg+3kJU
dTIZ9Rnwi+IQoFq6QQbNxg6y6j+oP7GMN8DVVovaLlePkChIcw6+xjPc+8TF4g9YVfUpXsft23sT
AWHVI7a3/IA6vxgv0L8fvK0f5+hODWbZ7mbwnBOvnHtJNu//nHl1DOIrnz0ecRk/jr71aSYnrBE1
CZcWKAdYf8MOxPvVUiKonizYJAqnTuzo/ciqmicmKCWn9dHJNoZTnAN3t7mQU29aEZJXKiV0rCfL
wZdKL02u3ZSawmRWY2ee2qPHJvUHzRvnnDvKDT8WursnDfFizI0IRrouX04Wx3S3T6Lh5UNHQjO1
aMMdfZkz3ApE4wLCVw3oMNZStGhqirAW4oAREKo4Bf56HpEHcws+jUdLdITO0K6GYDh5TYfVVqse
5sYCoss13OfcKxvkH9eVLcJvnZrUibEtgPzgf0+dDunipZwKEyYaEicttl/hY7LPHECbV3+XcGYL
SHVJG6IzWpih1VMfjkRAjiMFrHfjk/e+2sJ15ef61zrAf6V5ViLMHycrSktnEtLsuBxnfyrKiA1j
rI1dZE+m22Dto2f4/2oeAPYJJye64/LFirKIPTTcFevljZX64PpKk2PdwuVN+de7aRuf5hXm472S
29v1YtaXQSzbiE6VbDxo4KGxqWHTNbkhtyI6J6sUPuDxWGyl+/zU1rG2NF/hZ8qRfrfEfkUk3wnX
WH9pUQ5jpcbhzTUj49A9WQzWkTDDgGdPScvAGjWtUPYAniEf4aC6PwqjK6KQOf34BVheZtI+9euJ
PybUoKha23XhazTVwiNxKOkB0sUyBjzCRAIXn1qPkhwJwLWfEZdYVZMoWI/WeCcGHC6erttIpyxU
3m70D3I93EgkLSTob9Cj6XDpq9qszDAjyYYiLuDa6W6fPf9cm5bDFn+A4H68NGn6UIksZgiyOzx3
Bd4uhfoavw4bzxjumRS7DEHOqC9NRcClhJCwB3bTPr5q63QHusnBwxivbvnCvPdRuJlB0nY0iUDl
KlXbz6dWtiQivs4xOFJYwiLmnvXZ+IkRR2Ew6PC9c8FmL/ZTHmWAR/FqMCHvJQqkYZjUli9MD3+V
s5X8cIIfpHxYcbdVz0lyGQMaQNKBQuYu6E5ffPHUPkDZsB+U7je8dWYUggZAHmpyFR8T0DLhJS2Z
aYAkYdZ2JmGcsecBD0v1C6wqeAvSK6z8V2Veph6njaKqsiNRDREIdn9lAXmzz+E21AhHth2n2/h/
YHhma/L1EYN5LWO4/HPjT4qZsXMlh3QIP28uj1n5biZYlLum7DV1VojOhLAMozx1PYCzE7EJzaPz
Cd2mx5VsiPTR/tMblyeveYdxybJhp/8RHLvTpczCuESsmC6DmTZ7+VFL9MHYODKqAqaFuoTaHkgY
80hQqQ7fUAjgo+/Shh8i5Zi99U9rPc9jHqE3cOBf8BbER2Y6ukyfiZ7ymEc5AETMUPk9U/htYJnB
GdJdbGhvs+NUMyrJYThpH2zdWlcRlPE+TbgjqER3l7sYfXlaQ5S+9H3soXWLWfxjDrxowlhVnpoT
+2zdC3bI4fX1EL9lS1pGt7Wrd6kd7kmt09h47VTogl3+XSRvUMpA+dXehgzF/DvUUHpfjSPjDnIU
334Id76OTrZpo3YgHkWIalPCYHS2aB/d4/BI37RjFIIPj2IycotM9arSVrWXG9H+zcs0rTpeWTK1
7k/8WnoTjOcL/TY/YCbGr1ZzTdqVaKWPQyVFZnlx/vO5LUbBbHixarqdPItvik5OWVGwS119BgFS
KWVLmbr1Hn/Q4zDrHKal90q1MvUJTTHJBGoXGB+Vto7EIrzmXwr2G/2DHHoY+FAc/GXgVuOzhKze
B6pXzD/85FxD+YzEgSzt90oxxPbmESjCKowR0NUYfUrTyy1wPmMgQqVwfOlU7OX4rLSD6j2gIvWG
g+C0C3XDy/lUYWpsC2S+D0PJvoYABoZuATb/+Bap+UTNGbicnaaSIfytZ4xMAapGyQLSl+Y2JQnf
eB0rRrdDSVl015RjFVHUon3LR4o3GvuBdZi/sL65HzjblhgR+8tTS1NbENXsDYAbGGk/+Qnme/Co
Va3ZParqlA0jSDKXe0vbHNk8K8P4mKBYoId3r76dUBuIimsnZwmIUSzn47Oj3lhJyqTnH8yqGakC
wKd1dvrNW3uI05/CRioY+dnREAZN8+5hxe26xcidMgWwvsbXgMnAWXfvLF9rtLra9EW83R0OLv2e
hqy89Ez/PfZAfwscCMiETDdK0fLgXSOFuOprjgBO/VXbVkJiuKadOfb6wRW5Rd3bDDWZrkVzVbCY
JOnxYzIhw8cRSDbQS/Wcdjgsk4fNFtWYwyzqzZItyzFJAT67HN+ollvldLZ+BmKt6kCBahwh2RfL
kLF88q/L4j2QM3xRgRUaarAe1TMPcrTx+BJSFJBcGX2ACzZI/MAfH9AFIwA6ADSA8/zJ0L9Vuh1I
XMSNu/3NVDRgFGWTRZ2LkChtJ3PJhpo5V5mlr6f8PBfM2cJAqS80Se4mLTM9X3/qQNH7VFSc6cGS
qjszxHzfdBSl/A1L1u1R6Imh0IHjNOU9PzNwTWzecYmmTORMgWeiaj4yqgD/erSDhIWTZfrK1Szo
aRxnn+l+hTVhlKvwfYCsYXvbZgNhjTu9L3lN/3i732RQOXy1cbMz5ptpwlXr9yJ3hsX7nLH0AxFL
UW46UKFvXbGW6I6nLq9U6Ba1gY3jnDiz3tIQirbfBWp6cqFLeOz9ViHIn9zHWNcYFh6+69Xrki5n
11PKOo1XRgLIVm1QoHjH02fUR2Kkaikw5lXfonl/coWe15k31pzr/PV9rFIzSIhYu4OCToqyL/zH
OWDml9PqeqFJjtm3lGn0oaVhAQqruj9qONOcuY5GALfkxneaHAdpEMFI1o41NId7woiwsEzHcGGT
HCwesYdX8dIPhrFm3nik+NL7Ks+n+pZRfdoTJDvrLRxl6GihPTUs5NNJMlWwEKCLkAnc4sQeO/Mn
P5FXfrfMmdNmYpw4wMuYOab9BlzJKYx2x583EUU86iSTcqL/Y/YlHHO3RceYkp5y803nsfSkTvrK
C8eCERfXVYY//VIepJp64WoFGG1s1XmqdQl2tkix4dHDPJtrBUdVdxUKVeFmJu61/+loNF2rUv+w
+oxD/aTi2t06II0IbeyQ/Te+CKJlvQREIik9LiCp57NANzVIw6znYN87kNP4NAHJPW+d5YikhZJ4
9iwAdKIpKAGDVqG/paxm+fp7CW2OA3YPfo6y8f//UI1YedDFFGWj1LLRyPV9KoWH/1PrMz91Mbwf
zcDJ4YAzdyKhqHOo93m+WXwoUNjRiFNpx2QUBy0a+fURefaYT+6B8KQiW6iIi6ucALsLRwiIYTBe
hKqxrATRO3iawU8ZMEq403isG7Ls2i9WRj6M/jfEtRQwSYnUJbp3mGms6gyiOedv0vxG33AeuTJT
ClJTYO0Jr2P3aPl0Vps8eWF9EoAgcXGMW995nVhGzwMoKTBgJN2WKNx6KWeV7kAsWHUMzmvKHwDY
5uM87YVDh2pCyvTAnE08YqWZjClO2Dc4rcF8IS4jRiAVQd9QHSkFvkw9QNruB5bKAq4Dv70dR6g9
HvCkg79FAj/1Pk4sDAF1CWyrOWJlCRVzzJtiRqRquY3xdThTPX1NaNGQgpIAi0WLhA7hUA4NQhCK
WLmCWHM81iZUZLDAph0DxplXC20cqvS5OzY9w+LwC9kIACrzM/NrUhGdHuT2Xh6RJpYfx0LZiprY
0bir14dBlUkt7GiabYU0nZhdadwPOHutSZdePQjWR1O6n43ZQBPSlZ6Unri70ynEZA7oMxDR8QIg
mV6xePgdrwDk6AqHO/jLBB+MclTUz+ad10iPnuh3fg4e11aA6dwm4ZJGMH011y1ieSfSmSwykrd7
1WJ6EEvBB/h7ME7WQrSYbvpYlBF3JspTBENqJotkgmudp5e08uPtWX6jGn1yuzXs7AShUQlEtUX6
bxiXi3kbpoW4pR9/sT9UbT6YlnM6J5Av/g+ZvhiQghDPuDqjGo//aEV3EBOdQDOiqTfGJQm0veIb
YIEos+yhCvzJAp5QGcj58GSQegR6KbGeq3n3pKF6o6mwT/URtTmKlh13oYRIROAHh4whXFBg0vqb
hBoNnE5AnLOWhgTfKNhHxl67XM34gl2j49taxJdBgA2tPSPErJtIz1WuWeKyLGJR3mxNbHASNV42
KPzMnWyi3klOThW0NorX85FgvTUZY/vFPK5jYDp+58rckD2632hYGgw+7fpYL3Hho/TzQGcE8/Fh
27L8swTJt0X+L6PGygXfcynpju9x7ZyHON0N6muH6qxunXA3zy72/PxKp4x/c7G3SirmQMqjW3Bd
A6VIQpImKQL02MGjWKaQlTh+Ojs/s3QfDBsSdtFib0875RShRPwsD0ebndcUf8RUdggVxx/3qE8W
pPR65iJZA5r9y5jpq7KQJ2tG4LNgh+Kx05WFVM+hK+TwUiWqCh8/OcOsPLbF48icbToeo5yBvn2Y
ulTcEQ9ykIT36E+TFTKdqztof5VC0/Mu6QkpQrQILFSpwGq3+3vrfpKtTZ7lbe9VxgRWCRlr/YwT
Q5mKY65V/K5m/s/L5gJ/F4ZJvzICSEDArzK6RM1gi4Q+He2XoTN/cbzU50qJeXVELJQ3lqgLKDzR
iWTBTbZm6EarH7zjwQ9ii6wSL1+7OinEZfaJ/WXkdIV+LJW3cimtpbWjxDDuJv8DDOUoR7KfydE1
sPGmX3+I2OT/IyLHm4wHrEnRtpeB8PUZLPNqukrOgQjuaDz1AYCxQezcmQXyftG/10lbiHmbcRPz
CfuYKhTN5ChGcnXX+Ox6/lmVLydnRaLAnsSi1dUIZZl5qsdCCfef6MnGJo/I8bSngb+u7dPKzF+f
B8/ZLuUWezUf9ZEobWJL3/z6Igus867uIJrlcFHJUU6wph72JiYbKyEAuQ1EAQ4iiXL+ZV7hAJUR
mu/hWTTrNOWMhg5LNg6z6bPR3ZBqqTA7KTMoyqOiE32XHFTm+4gaaVw/IBrFKgMetC01Bxn7Fwc5
JqLIS7fx63kdjidCVVczEDivcGiogdfaxjygC4if3R3WciWrlYfOpp28reB9oJhq1VVXqmyRD1eH
0caAdXTUWkfCZtpF0dME8sPn85p/JFx8hhizDbCEUXVLu8uTdjKBDiaCydNI2an4V8gIK72Ke/qb
gF2E4Ptf228XmEOX6YwCbz62SVTOGn3Ujq9uQFjpEf3lWG/47Q1gMxff2hPdrC9p0doj/CE6+JjI
grd6oanmiuGdzZHLHQrBFdsvfnVTSddAPKsQDjCXAAcF+zWgSBuIJbbi1W806/JDMyhhTs4Q8Qxp
6pabW0bHW25/IvFNwHrHgqsgFnCJDhrBbVux+AgSfsBUqHWkwK3hRyDOcEo2hkpQRdfsdZWD0Kdi
xYi6fwhHXvWLylT7Xs1DBJVesY5+bQOCNi6tINoQHEp1lfVcTpvcFcw1/qFSHLN+WrIHjI2WJEUj
yZeRpW3O5Y2EHTabFqIIDJNbnNoWv9KYRRgmghJ6nbPnYH9DB9E+Q+36kKGBocv2XfcmL7mtiWMH
ApRNVvDg8GwdbNvz2xD2aiZ7czaIh51dRNf3oZCg5cV8M4Y9KBD2W4oOfHlolfm0POycoPAQ+Ybu
JiF1sO05lqiwclHGSJFVwCP/hkp1+Zh6vpF3Wun1Wgo0JUGBj7dITfrEdfD9g82se3+9nffvzvc0
IK8Uj+1Lk7h3G5smZOpDOJ9K+FQaex5L6rYpZIwHascTOP0bRSsXRjuJ+9P50vIC3uW/QrDXeYiy
JJzq5OGdygwDKHObkjy4xV/pPnE+yCM4iqPNXjUM9CRFeysg6IhdPoXL72uSQ+ZzvBtYvmUxIMqW
2+1Ou6WccQL9TpcRXNhLjVhe7ovfZS5opQTueT+g2fWtp/3GchAhH4HNSJfNwZs9K/GyMdSgIji2
spy/Z97QWaOj+qFavECIhnDdfkkcqMUGd5VO3/NDg3E7+MFi3unAZNx3CF217+UZnIKaNxJj5Xzi
NjIcDrhIlq59fLknyzsyvkK8ssGDgZ7DATQ1vgCyyM2VCwAA0uZS/kXRNjfIzu/ppD/SS9sKoQc6
`protect end_protected
