`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
RXH2OYSS6rA1a1hsDIgIgCN0wsjVaWjeqZ3M+t2dEhliPKSa+u2rCZ9kcrXN/RwMOSZASz/F4GVG
CTGoso1EEWL+ikm6+Yd0UuLbmgjGxIIqzVc1D41Td84gdTLVoeSu2KhbEbz2IROwM2m9z/ScpVn8
roBmOcDpC/DiftslX8Fpo7i3k3JbUY0wLPorjDKK6SZa9B7cWIcMzX1d4Mw4MKtKwJBV84+hxqN9
AgT8Bei67tcDI+EAyo+hRNJI/PSAO/jPJdU/ZRQyi3IabX8R7ofZ7rlXlbAd+s6FvMR2FEm/FaA2
wYEcMrAvZLzMCx/S8HavKjvbj57kGzv4cF7I4g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="cIzB2k58g0+dDnhE/Okxp1Zl81pdNsL00clvewUUkO4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 70544)
`protect data_block
GZZXXasCXTMldRQ1mBNG+ZS6YtqO5/r3ZSAPnIOypVhLRcFcRq7vVd0hgKMwR9C6/c6mvRZJLOjl
gl12Ql8jElcqHILmELehuLKz747GgOzr79CEkRcZD8sBnzAOp2LVxwuPC7bmMmmcJOS0sTitUZuK
J6qM9nGvTg4afV0f0lF6MFX+op87hmqm4llOlhgrcOOIRqjclLs9lPkymsdrrVs3evwyhqbjxLMF
AtdzfK91dUvKtqsqW5EjAYMz0tOlqw1Hy987VLf2N8C6O5ygj6OJVwm3Frgy96VrRsGwlAlTyWka
VTZ9JJJ9nx4BK9LSpryqtQczyS8Ks1s18yQgbzPNwW9TJnRiABSml1MO54TRZUMnwYxx6oXtLkw0
MVTqYH1O9j9/Xl7WiKwRgRktsTyozHLjI3kd6ZiVZQprz4JpuzBgM6Xb7lA+11s7D8oluTzxtOg0
ML4kfiD9DdWiFQS0aUATkCAEcJMtHF8rz2IAcoBXBt+Kc0LyRk2BypoZe0KTL/x71jWOMvX958ZO
XSzBweDT+7cnBsMte40mzVUFgWsYl2Aied7SNJBNdky370eqqYgWzce7w7/NUsJ6WuxoeHUUnvqD
P96AM62MnJ4wFEJB6Tawp7C7vRq87/MwT5utnktKqcGZgffzjXlnq+DFX0yQ8wYWuclHwtXYMXQO
tKRKg2cyHsPihcXQpkCgXbgrWog/bb+2fzOdlBZdw8pQnlM3I9eTi/Bt4+4Zjk+Sy/KAfcM9t4OI
IVpM9nKF7yM1zSfmnXeqwB8J7ubR/t3eRqtm2seqYLGdzR8jkStOGM+0jvG0bpdxKrbtXSqi1brs
LokORILnjymlt8tH6eQyHpVbQwLmD6hjNIZ8WLQ5BJgn8sJzrR9LVdBArT9yrtFTDGibqgKOigza
IiBz+LSLQqRaSxj8A08k7scC60ivURR55AzO15lGps6yHFR9F299ZlCh/vG+UuDZLzWNCIbP+5+G
ivft1B+zKNLh5rLP52z4ZsWiIF4bpxNYy4BJHS/JD/cMkrP14NzQ3gSvC6yKNtis3PCKJJUAT9Ta
/tjOB45Q+SBqYnUnvCtTUsCQdagsXRZUbAU4rp3p7SFPMXh9ZzipDreGdKSstqIX82BeJFRQn0B9
DqZmkSDopvcMuQfPPsiTsIvYHg2jfiPs64X8RW+tlkuoA4XAuLfASBxNwA0odWYC7+iW3l8UFe2k
kEnl+8pG2J2WoaaY+A+gJG1r1y6TQWuNN6l+ctF1Q8ag5Fv+36BBUn9wkZSbmRiQRw7odI4W+QqY
gN+OaqkQdPXnJf2xJLNHO8ALdacHMTXPYrd4ifmLx2kALeUF6nbgX5653b/K0LNG81QKazf05cwn
M7cJuxWHxBauIc84PkoMunvOlN+Ui02j3Q43v+nqHsAdeEfXoiYQsiSDAonQG7ZKF4AjUkQ0bzUS
iZUqyOfDAAQO9eW6KAp1OAMOsLivXs7W3qv79Vf/PpOsj/ciH96Gx7EnsSu5Ab4YlN3nqoX36QoL
Gf86XS81StphDqZ7qHSTzsdILdTkNKWuvJk5I2falQRE3A3DlXWN/K02j2yod8CbjfGUFt45H0F3
VsSa4w1VKgEAwhneqBHo21H7TFrHKNj/GoOixPvtyZq61sG3RGF3G5rnbIkqvpxGe9afabYxAYfs
X5P1gHEEuGRqMYFM+davoHU1diOo3/1o8z4Kn01EEkISRpkeRIRqmv2baEs1ByQ8oWd3RuESbmEI
XxJPA9h12e8e/oh4qc/Cut9+oIQRGi4L+TICO4jRR/gG+IRIu9Wzi+9JVnPdqvB8LzYOWuujZJ/x
Y3mVuTfAJgLlstZw7WYYcXcl6+tjMASfjsDX0qcM96Fi7ctBeX3uTF1m9WxPKfj/L/Myfkz8ySaA
woSrUxfLqFl4HhcDEbe08GB6FPdmJY83KkJ3qTYvb8v7o/c/2v6+3I8aZKn2BnD7dMrumrj99kQR
BuqQbRHld+2F+EeEUL/TuUxsnQrWTLr9S0eRQ9/ExPBq/aXx3WaB5f1XeqqECjHOcfMMV5Sg15KB
L0WWwBMNOf5AcFX7sGOUz94Y+TnThC0NA2AJbkaNtK2lkGdU3fDJcqSTEwaNZfLBcrGZYfThsnKP
+2s6cwVjSCQar5xq4psXXlRmPsqBursmcTWcvpVY9iPSRS05nwXzbNQET7Rj4zTcRYFrIBwXG/1e
fuCJySrxM3XXXgM2ataAEwJGuBC6n4jGQEnMwM+432o6CcgIZ8xwmjZplVBQH+V/30Cta4vWRy6V
jdQwEIXUy3E86Eiqzy4Zk0tOiEXgBARiCxBTcJtNRiaYJcMV+msjxnA20JIkAOWdkasTkOmIN25T
SZjCmBA7pGiM4BF5zpHsl46gd0N4dzgLZGkPIRX3xXZDXKbHRzWW5IEiR6frm2jAwwMr1he05woE
ylktEExWYTLRGyy0wB8JbnaRJ/fraC12u29pofphPRAytcRHKUppGjGiVmCu3MzrWFCq4CP42yFf
0z/9hWJL97Z/4KrcrEc3f0B1IcRsy8l1HQYB6PkSUQC2FRsO+KRxEHyJzBCcxMGpiy1vidfpuBLN
OK1pzLywR2sgozFFE/w/wTmNQajVdrChzZFeEJh42cf03HTnAnc42/LWeg4GlFSFa/7SIb7NtpOU
S2KiP6Mg/5UtRl0QJrK/vmqPmHcOnIIQPgiYDrj+zS4pRMUsdNEiLQf2KhkXESWOB/xlc9L7hG/8
k8w7qdCCs9WkIopgtFNo75mw9HLmv4cRTOJNo2B3JLaGfNwaiSJy4pnc5560S6prIR3c2v/n39Gd
HxqEF3VCiGozA0N10mCs/A7012hjOnV+xY6JEaH64GVUyK7cMfjVlolO4zVl893LnRJ0aIt94pVs
vti2goI9XJP6oafrGC3UrsIlQ6rMUoTLAn8ccDIqA2JMb4qneX9kgM+KoO3+fdQNF7wWjjSYYEMb
iOM6tkKbn7YFfwQfsOgB9HnC7fK3YN80C1pvZVYFxa1pT5xv1HS1a8R/quS1EM7wfC6/HJpsqeUG
4TGqDpo1yhRqkTPc89yrwIGIptxhzGihfdSTbgIw/NYocIYoX7m0u1Qwev/WjFJNTpd33WaxpFmA
KNTy9IFvOZi9v1hjq312E5/MqSoGpZX9sRsY3cI+o4fBSMUrHHmO9qhluuTA40gpLRsP3YWi6ibE
cRa8gmhD92XM5zsx24cA/7mLN1BTRirSvQ5Z/IYZ3dvQN8aOAlSyzIGjrUoVOInV4Ts4dF8iMICS
fpxTUDt2vaMhKXSEYNimYw/s++oc7Mzxwg05DGJek5bjyYVlTGIocnwY7hjxh3Vho53PQW5DYRjN
Az2puDJbSouaiGronih1rJhWWaCm+9M427q3Ac4RkND/viE96V0PxMaHcaI7FhzhpD5M0DbAvL2X
v8zRlZyOWaxhswSHjeJ8iloIPEapfTOwgO59kLptdRQ9tW2fNiLyh9/l6i2n8IBM9JtdXMBluyjA
tgdx6+xBMGc8fnpc9IHm4lq3ctSsWC1CZpQRNs1BnPeLZFKZs0sJThVhxh7yHFUhZmpywHZQAcqR
K7m8p18q14u8hQhOXJv7UjGbOzxvoUaWSnpxpFviMDrEMo0CXWBfCJH3wxjDueY7uMzAniWTHbE8
47QY6jrHrR4bJH3tfgtBNH7LaR9VtkI1we+bKAnB0ah2KKSl6OXni6Na5NAa41b+AZUfIrwXlGQH
qYtMy4tjc5orcas5RqNPlfx/ymX/g3NllS5OQ9+427fLRW+DjocVZ5dBWeOwUG5Au9GSk74FkymG
PUKPbdW2oEdJZjbenu3y74453NKoHxjaBYgGgkIjnIu0Mo7YludP9Bj4ZpaC6imDngNWXCXQXh5Q
z5+348a/VQq+EpnU0eCEYgi7PRKre7DDq/JnnNQbFx/euldfDQ+zAjIdN+HZPv6sEM5d9RKPO3Rx
bS/KwjREftLuoSRhh1zPV84RLSQHQGSRiN88Bc4MRvrD5upOtCJUzfoLFS+MFrMI/l5iMhGMbHpW
huoZ7bzn+RZZsuGHWRPsrrOrS3NK7gcstt0EdtPYz2hzxQN14ATUTkItjKoFTHpUilDihWfy8yme
hc4BHJeo/kWc8+LLdrAcMu1jxyvUzsRG+y+hdbzI292G9aVKsqabRgVZ2obL2HZT3928WOVnVyA2
tpAgXsOl8HAoWbomr9k5OurGdWB4y0zmrySUwgZ9bTbZdklETg35CHVWpwAZBZEn82Pc8qX6hPz4
UuOxvk+8ly/2chN0rP+OvJ8QHZ3ac6X7BDHyWZOTEK5ROXnVaD+c3EI/V3MSuSPsdpkqhmoLsuuv
r17NCZww+oBD9kNoBeV/8yLWIe1JUQZpF8Tr50OczBheE/7IatGXRByf3HJCN146UNpP1cSjHRt3
9xLRvo5L01sqNFqHqh7zsQaqFB6X0o5nQAOevnEDNwcra2YKCdHaQBtDmp0ugcPH0oVJDc5qc86R
2hPkkE+eEgxKhAy7VO3ZtygTifVO32fjVPxGX7vtmDutDWPApt+cNxXSOi23Vy83C3NT+XzxXoBv
1HOTqnTb+WZCZaeFBS6AeJYm19eYalofGUslPNONSrZFJZhO4uS1YKCLdrTdYODzTqfNT2JIcPno
RQMov+mYADIEBTqXUyiZFN6Wm4t/14qlwNuKxQDOexbNTmaRQAyUCylSWyxdAiyHZ04g1Ranmp1K
KbgP2khbA8I0m/yvOkLisy37bH70bouDvSyjj71O9+8a+9TdRiwaHRvAGKV8tmOYDQQDBOvcPnB5
P3hyOtAkoEQ+DsR1+dpvV4UJkw8noya8Pyx6oY3+ft1Ga+AB10YbBTd62y18uB62wj68LhHdHrN/
YykxmZArq0wkaf9rb+D4REFMLXguqXPNOuuc3xdJpVbO9Nb6B5bT81gSnVgThRQXOnSu72p6jswm
y5C1wYST1y1xJBWfPgh6uUXOV/4eki7or01TF0q+sJ6S0Y5PEVtY/Rq7p8AYslmNrNtGLjq9G1qJ
MHaBTA8/jdBvmGVxqNNu9hgGfC6870RD/xDXsCytekvEdty1v8GTWcgQ5zjKaco4h5bHGkAnuSPz
HUAOOpmfanx84G1mmtOjLgiyT3gSZoocjmW7/f7YSPVG6757TILPNwXNn840ixyLwCCvbN03Ld7X
MuVyzfTsOx1lHNycEbe3kxq8SISeLDDLOUpJRSlB3pV6VoJi7S//rGKxNTRFjoxtuC20sYTaHrNu
dbTjlRXqfCWSABNr1o04cFm7HMQ9aqoB96wlbwgbqSt9RvMBS0UApZs/AuypJuuFk4PC4ut4jymY
2KId/5SdjBFaRyNTEg0Qhou7mhICXG4F2s8qt+isK+bopUVgaxYPRJObf9q5UyqBZfaSfYJk+/SK
GOyRkAVKt0v+054r0V57dVF2SdfWo136KhM2P2SXX+HMdg3Em3enrE5q2489Pa4H9ZtS5du9UDFX
GJLaBmr5izrcUUzO9E/f+fm/B1DRk9T2ePcCSE4QJ0Ylhctzs8C/o5u9RpNngGLh8P2FFb/3VrgE
+dnWBMccWi+5JbxqynZr08h2g47MROaLVsIg8wYLBn/OPrEgcAO8FYA3biOFM/Fio36aEwSqYG06
vP85rXA4p3XrrI57GV7r3RZgUxyLtN3QjM9RXlw0NeoOmZht5YnaDasUt6iyzDyz+mv4HVMHbvAV
mTJTPo8HQsz0TSnM8BCZvmprNmUM6aWvX9tnH+1bwXMNCImcWm5dkAwUTv98pf4bJ/YUtlf5RJWS
AWFVgkBbJeFCRBdlBVI1WjZKDwTZz1pRtLrdycLIrr9qFIaUTX0WpoQR3rqUUGeXjOHDtQRzlfDc
CFePEvl9/jmgY1sWf8fVOsdYJ3zkP3xMjB0T88XhYtxJ9O4fNztUSN1NqDtv2atrgRZ1nxovjkP9
4Rz0X0eYTULwhZ2P1obDNO17yHeGdpVp58o7CTIg4AuqKIoC2nwA4mqSn+suAQMOK96+rU9t1KSA
cW8qDSJv57+4Za9mHN3NW2eg/AieAoAuCTjL5WlU56ZvJg0DvibQzfQ3wOk1NgAK1Vrc0DBvmLje
kb4mEaSDFUJZH5i3eXc15Nn+vFWZ8InCtGEBsMpkBpYewzUJ6OpcL649gQoON/2mddjm3GBGD3yA
PFlprKT8Uhp4hrZsMxwcJR9Vdr9cRz4SqcUVWkU6cMG3EjRtHopNfHBrXOaSp0nA2TrDlOCnsmAu
3N5eEXQFmre8Xx8pOYgafWuAtnr5LuZGnj0XmqtTe4x9LALSXuf7Kzqc3bcvHYW2Zmyh/yGxkV/M
1NlyOK103AtPQHmzWXO2JZaKPWjU/1LtN09Sfghv2XENHWuLbBd2wRgjDXMRYWLO77LAmF77feZr
sz+8f3XGnjguzTNqt0C8hO8ZG0wlbBWK4KNEWVUW3zuBJ3GpXuao5TV/hc095fuY5TtDK2IwfnLA
kkuG4ZNN98CHGQxC2YMIGi9+IilfvzSkLx83w1tkw5iPKw6itxMjS66c9uSrHb2lRVv4+qb7y6gK
/TpFRDw1sMLYqwzF0G2C34TEtwfIedUyMrHoZd+UgLUVenewdQDB5ROW72gx644IOyvkLnf+1eEi
422Nrc/dIXsDGB/Np2Xj5pXBifWd2rgxnIaU4ChhfYR+Lal8hQUYA5BQsU1qCvu3rNe0082eUpsZ
Zvho2l6fo88DS9iJSQS2hYtqMxTtR21EoGlcyKGDj7VqoWNNG0nszqBgy1UX3+FM06AEu28R8Mrp
fFBtxwlRCaBNNC1n+x3dmzUUhnnUlNTX4FUnbLjyQNAKWWFc2fGVygMzYSkYyugCEt3YRBeygJKb
+QvnhmLEcyRgqoDjm0+NTX2Uw67jkkAVI2cGeMaXTc0NjKgJbRHmJrXRMV44Au8b7iWQRlS8hgSW
wPMx36/kOBIkPAyg4cIC5UrB35jx+fLVC63JWs8/zjx0gz8FU9i2oqWS+h3elb/IhDm86LEDiE4Y
Q+I5/XPyc0RUPKlP7CW42cQgxBASzznEB0h0qOmzv3fphqeck16sOlbDS5mpMkJzxLzc83I8BzSs
zarwlhhJJbbImKuC6oTrA44OEpuxnIpqrl/XN1BIRSTbpM7UcBaa3HTWthJo5E/Z0OK5XKbkQkdB
VtT2FQbCaCOc8EZeu/yTQR+in7/idcM4RMNCbU3XrCGVdzDi7ZnEhsDHehTX9yqwZl/VHTC03T4p
vn7OQFBc4P3L8cT+mnn1dmw0smKrR38VLZqN5js2w6APNyvl8IX1YX04ygx9pWqz80T2uRcYKacs
wYiib/UTjvmsxKsF3CyKxiSZJHC4OY2K78dw44wQ01y93wXeL+wy+wpg1qcpEGT3O4DbXgNrRNcJ
CkjQZ4XnzkwMEudxkVZPUC4Wkyz4DYZxPoNxPDZeFT2PjL+0+3pg6KjzOQc6mVTSdddem4oSlrV5
2+PIiC+leWg37PU97AroYjlQUraV+vF4WQdRTmYBMsimGWbNVp3hMqIX6uqthJgQ+u9UunbZxTNo
9JuVsLcKNPK3zBPYLk2LmdpvW0A/vYKdWogOsYOge6H1UxDdooUK+BBGfaYm66easrWh+dRuUbvP
B1by0fv2kdTCDGZNd36pWMZar62og1BGTZt1k5rZrD0R1CF4oslS9NdxhEAwlcGln4CVuwCxyp3X
+2W6c48O4tbKt1IUz8VqO+3L2dQQz3dXY6V0g2/cjuHA8sGm3UP57FbWBu1v+ZuQRxGhI6eZ0eIz
N7igbAE0+oPiVEno1LCp3ifdU/QrrEXACHir2JzVLh6/Kpfjq4ySI8Pi5D43cnoR1cIvf/WemN61
70ZZV6+LvdcEmMKsQvFCGDapktEEIoBTfF8KJLzwxCwZNdefdt4JC/2iCNu9vxlSvrMo1wanv0wJ
W3eoZc32c6BKeUyvHnZ6FcN05SP+IbllqGMA8JIyDEnZROXg5Ww3mNPCCzKzth2sQ26pG4gV9U0Z
3xm/QbatM/TInkg5EpSij128C82t+1tdza6jomVaYM39H8vjetMOmoziXeygZmT2p9RbY321yhfo
USFImHb5kWGD3h86Io5wFtOICYXdA1R0d/5kmYLUo5xKer8B6n6S4y6OAHC8CmFMTA/VPycBO0ZJ
rAfcbCiDyWh2HAHeHG/4njqstk+PFOK/EIMQLAh/2ua2EmL6RyPAP0aE7Oc6aADPHg0L9jw4Y7OK
3WQMzGOJBh0zEAWEQRSSytl/IEJBDHRonMhDSc/oZWfZ+B6Cq0DHb7SqKBIl4FPkGzlR97i+icCT
lZoFmaxsqd0nu38q2sKhrHTDvVKTJs0cc3AG0IY/GsnnG3o0LrK/mvnNEJ/frgr095N60SWuSiG9
v1krHkIOTGAclM4/SKnidQ6Yat5RqC3lY2In59nHL3yts48YeQDg74KpwL0rqTNxucXvrh/pduLu
RL6qfbbFe3+2OBY1wgTOB7fctzLC9aGiC/DAiVYMxJ8PnZOIaaOAVTLV8D6V3v4DAgR4JJJgXIsU
3Rq2nu5Bp+6qy1XhUHr0bmyzyihSclkCqO9TYnD3SunYfI9aUc/qthfx8svLoHLqmGiL7NZOZZxv
hC+Hzh10+F5+Roel32vc4U1dsaGSjhPX+GTLJ3boyg12VHTMHUtEHPg9VNySsH4lIHydzAMTW3lh
INEA48I/8LQFVfx5CExO5sVESz+WMvGoSq10cD1HItWWEqQJDSuyVp4t2KEgG+n7OzjrWZagj/Ff
Gu7y1OYgzJVSeAxK17Xcpa0Hpk/DYYBblSugjxAXMmryM/gKvdv3k57zQ96N5mBZyNEMzqfoaWW/
Sg0VuPtQgkOJhRLyECq1wAT4XZ12bYqHn98VcFrh5PhIC0wF8JODjqlOw2FgixfIwjHdQduTG72R
O8t937q3O8CD5MMZJS1uZJg+DkA2zf4UR8xJIUm6GXs00D0iM/FVlRDyWGwHJ1XygZ2XnicRj2xX
y9gvmCh9pj7+4kYzUQfOiQGhlnyo/F+7Xym1deYlUtSDI0VltuEOB5LbEpfzgMg60uNezwohMNkm
n4of34ec2tH7FBp33T8Vn0aVlSMq/88/LyqnPIoSoHSPuoZtTPDBdo2S7J5mtbWaoMXjt6MeG0qW
Hl7RErFdUpOPoakw0YRAIVxxoZaF5Bgv3vAW/QtZw1IW6CeUqaS0JYqnUBputcOtf4nxJ+zhTV24
hHAHRyeGRgoxLvfnO3EdtPKVlZfQ+BP6LSB3AegGwNmgsLdI0QyHEjMlUQ6THpizznXB2tTiyiLO
lzrVKYmChgUGRTDPoIzL0gXmcTgJcd7COqPLPTl2IMd6u1OKdx7V9NDa/RFlq5Nq8dZduK3cff9g
oTg95wSe56rLkielqhSVE0c+Z53NWB1GW56RB7MBjumRR0DYNFQ7LMIB3ZqxDi3Blx51xsp9+JRd
HRh3LKZjxglg7Ef5jztG7McpXFgYGwBMSXWRDTTrs8Q2cgP6zo8FFt0bYWf0xIf5KiFxM7N+m2wE
e0OG/vUEqRYxHwhDlGLnK+3DUv7AaThhvIEd7bfOIZirAjg2v1LNR/Tf7NpqIws6XyPe8ISL4oRD
hvbgzORdo1JeA50nl+cYCWvuCpjlDJhMRNfmf9jwK/oxN26nTgfCZt6M4Pg4dnWTodRA+EGAmk63
NT4Hkepgub8raKS93I7U2SbCerr8z2KjTfwN5FEdLuhGCaTXQRitomkVUeGBMukNF2t0A6mAmZB8
+JYvob6hBu0bbGi6tXdMVNYSnkBl6R2bhZLpWikGrh0n4LpMVQRhGYFUq8+Sb7j9pPrKzDFXoR06
+NKgSt8DTxuJejW11kppqsrXevbvVrWpCAfhIrmLHJRExES8/G7ae81cGGGSrTGw5ihoI48+HmU0
Dx1ByrdjFKW+gZa4pMIYA0YA3cMYnMba+dLtdZzNhVCBGubdf+G7tPEttj9NvCD4+N+tG6DY4A3o
8Qs7wg9Ca3QBIJPVxpNENtmExebQww6eIImQj99NCCp3GQHShDVAIPzQZtlxPH9oAFQHY4oR49Jc
rggS7ZhxoDFR9EpQWEZedJ4cL7V5WwbPppY2MlXyh3IDq9UuoxQifXBINxZcoKDTk/et6rXt3ecK
2XIMFWbDfTMhvAlgSIi7xoGkFhZOHJRWeoRwnB6SAvrLVgmOMSVhYDvbyN55BwGwkbMz34rnB2n5
RU23FViCSrQq9JNtgBf4a3Es91itc+oPVbCBElWrRPRGfpxgskZDXxulbKmUD4/zybIY/dMJwQZy
EiO6mxjcBBoiyz7qu3Fpe/crGPw+sQkEWMVtOl/zmwe4pJV3LIRkT2dRaRusmMaGvmZK20/0Ur+F
UWDT0AT3f0DEihKllRi46bJQsDExZ4F8Rnky8YWSgvixVLAOxf3oGSJcc9pnyUpv+ae5HeG11uLY
oyuasAZlv85PgtHNmlMt9HYno7Jwm2LitTRc1rAfKdmq6mqC/Kp5h/IVLBWygQmL17vWrXmTJHjw
yaD9nsrtF49FNIL3ElSVs/cVVOlKDPxnd7V73abXA3k3stUzg9IeYHMD3d6LcaWWlek0V8mm0+MQ
X/EB59uzmhUsaH7CeTM5rwqr/X+1YJv0tPXNBxt3FGxd015zTMyrAoSHUizSvmnRYUMve543L4KS
onMpZ9ZH0uKS07uLaWZYxBz93jNz2+7HEhWwmE8Jxl5VTkH/IzkGyVtcFvIC2WTSnlluve0vWw53
rCASDY49brIbE5aftC8F1GpGffJ3KQBMK8zr3B7PZkAJ9ZYVrstbeN7DnyIoADNV1SuLpT2FRZFd
6kAjHVgBP5m8rVPYWLLeZ9xjUhLJWEGBQwGRkvD7nt1VZLdbykO8IwkOe1zbM1fvlsons7K3b0M8
UActnKBg1BPDaKeWiIGsjmp3zeWQH7VkfyvmwzLucEq7Yy+X/3ba5QKzjEPrVpFHfLOzgLFOv1/e
quxNpS858WkJTzIshL/OJUUwKZp9DLV9eng5uSWCEbLf/9NhBF/OIk+O952TgzgQLG96jUC26xLv
DVn21EdTIrFy4c42K11zMwZC21JgruyO51fLYP+oVp3hTykYpdrT2UOU6OBzNXNtxfqTkYnTHuDi
yKXazbsxkDLiUa5S06Q0D3Z1v3BPauP0o4AWnBnLpwrzbXjNK6E0Hyh0IC2bxLUnVLX5K42jR2qJ
qxzHPII7P51LSCZX/xKate8g7S9Bhj6fEo0GnKrOwyRNSCkq1s7QaFgxncNT2rtx+I41mECx5fCf
NZN+pew/PWRDXI6/PbPz4w55u8kcFYTNuGPJrd05Gmv0fOKk1xue76JO67mfJqgd5TxDOL6Tn948
oztZDJYN0FV2WvU2ADjvyJVwXEKRsGD+2SqA1+a2ySZvxV744HlT75Q4KoQWIhjRKRH2KMCOltER
Y1gsPa89lETxeT9OhC3n5C0YyAhTnkRpsjs90pz0943XHHJEP8Xu7walcwvSFVigH5DLlWKeBMu+
xcsJzWvuCfIBihuqoYspdRj4tIgudAphqxkRS9Lozg4cJS07lPwrMw38xCkO2H2+mUTGAacfRUR3
NM3f8RjHUTW10uW5fMiVeQlllMVXd/5IwAeakJI6QzH9cTa39s/SNLK5bbfuzrKJQblpvGP0W1wh
7gj4ec5fzgjNLp7tPCC2cexX5B8Wmbd5U0z9ScoDXUTa00Y771x/JXr6nx3SxLbUdICAn0A7UhuD
mjL2gchyL4bLVB7MBQPwtndLUulcdbo7f8qhK/VcTA3/57GYn2Qilu1jTkZrCZluAHbgf1qBV0Ri
MixMGX1lc/MkeQSyFW4ulnpLE//xEcf7zIu+q37bT9nFg9AXTArXZ6OOrNW2hHgZKZpblaheZjGn
dMGhLItcJ/mwwWNSJlnw51Sm8gNmiw9TCT80ELLyTXgNDuNyDURN+aRRt2JWHssLf3OiW5hpE5Da
ZoycvuXh43S1QQjx8OUkN8nuOIFMjQ4kCUJqQkHF8kAfG9sZ0tx6EoPkDdUWd9AgUmx+9W8SYC71
gf3mwUc/1n0v/x5zdHiMoqvLfx+Ap4AXPlDFVHtBGnJfUq7vjsiKR+WsMAA65CisO5t2TSVuc36K
dt1NjSTVcf2PyABbDpa7k7k+PBNz6uDv4I7NZRXdpTPihd2y/gWGQ8HVxhmnnBrq8RsDIOLg8Aok
9CXjI4suBc6t0PTJilRpkBLMdjZOoKOSGHq4P0TiVaSBVAAsh/Lf7MwaeoI20wLR4LoUO7Nrrj0w
TkDf6eo7AXtkbWOv409c38HriwZG7c8uIGSGplMUNCUqsgDFVRqb/NGAVsClfPElJomSwJM4QvwW
roTPFBS6BOLlyJL+f+73rOb0jqgAVUTu8bkc+j8dDNKSu4Hr9mkOnWbRZe0R6QLUdE278C6ZeR+z
xbIBbgwATzjxarkPjAu6aD7VWf81NtG9MXWYX2bpDpTMF8nqTTEFL7s0yASv9/hvLI+PXt4f5t9V
UVN78qSxJAW7JliQvXmiG1hv5GozyPVGRdmT8MaaFqXRttpcFRTommbU3CLZoCPFCXfRF+/6pdmY
pp8vDwyygbFGgp4ZUXGGDm00H8jAwiyODq3bfw0BA0gIKCkbhjWv1NyRQ0g8eInJILY9jHwcwuKB
V1lBXOIpuJpBtf3I44krg0+VO6KpXnlhooNzpEYBQGY6At/UAyVRXzSRNCVMHrh+Soie4VwDPp8j
EOoOtkmoRylfAvNHCmug8J99k40iXka5wsQl6eh+fMZckrQ0zQib+yoIyr7ud3zi6GyRXCKL6kz3
mUP7Wv8sPJ7IzuKBxfja40c8Q8KtwK3QWLETb2LqKb8MDqhjHHFPupCPOr0rDbJtw/dvWzeuNR25
0e156zYDhIrv9Wmfh8dWTZjxvX2W3bc63lOuKUHR8TAV1pq6ISfsyOQK8RjGnrScacEu3xS58xma
VxvbI3NorSkSYWY2GVwx6yDDX9v/15T4sg6EEtNkfgOfVVVGiJpfDZ+XdyUntTCKJmHLxKG2u2dp
AE85qmztwHt6Gd3JzBHIdjYy6Po81jEAYkszxz/QLm9DduYV+XSrDJPBSrH/dIhb0b9Uh1MFiFqJ
+6e0ka3v9IoPwuQXyc1iUFT4/XLzqS6JXxZcApt2LCOyENwnrcB0GNeuYwTd7Gl+uBhX98fIgL/y
kh+AVbJ41UoYL4GIU4cBxz80NKOUB1Ta5Bv4pgVOXYDwytm9pFRaV7CVbE9eXcircN+KUNvAxYYE
bHbk4fpg6vnC3sUWdhF7/R5Ty6KY8o1WWSryO8+12GYLGQuQ+Z7Z1vuwa9Jfd5w9RFmXmMpRvT/3
rhBvM+ACCGifzIp5XX5EpNkmNdGErFlEdRkmJwU3tfJ5qS2+Hslowpq1fcTYJeK8klONSTWda5XL
WYHGxIfquqS5RbGRr8RUkyvBmvMgQQyMTwTVdV8//1s8SS15ngePVrPR7AberOzMrULcpbxOY3Z1
C1/x99NkeBKitWvbspw7NXsEF286ti2ovtkJZUvZykAvmJLHFiKMc5pPw7QVpuJMjI0Y2pjdnxfw
DLkVwiueSFZi+FYl3uWpwjHBaFL2k5HFm7kJnO0JAI9hhJ+jF080VIjon6L5EYUwLuLJosjNgi4s
oXGO1n/iSkitf3/vroi5JPc9oxng8FkwjsXwOuFvo8GWtrekpL9pGw0iZO5vYJm4+cw8O+A9pACZ
KYhRQ29X9ZEXtzfj/JJ4wVBQu/3BR4iVUWo/O5hL6ah3TJyu+WtTZGOyhqgVC8nDJEbw8lBy2u6E
MNhJCV8cQ7pukFCrPEWsuUzmvNA7z4arKYujLQI6GiAaECYnwcoNhW5HULHsEYJ91tCUfD94yKsF
0P31VPDupLwuBU44gt57CWqJAIeXIDm6MSAOiVq605d6ofSGvr9dLxD4jEsi9C+CUZyY1GAkD63Y
judvF+qk5cfrBmcyHz4c4oaGBadQptrIZMUGCHMiNTfXXEkMHrvMzXaZOJc/kTYo+VJZ2nPwsJ3L
5IGtwuVcFYASveNye7+b0NU6jsiQnVq/H4/xU+Ej7Iw7cQkxrtycokC7gWZWM7mjhmAOro9mzZAb
KD+FqW5v/MQtcQDojH/gmOGN9kwJ/7tLq2qeyeoD3M+d/LW5HNE/ULiuCjhX7SVIYeS4Ye2za803
NyPxpWZxGkdy+PRiH77fzjZx699ODLRLRMcMz7IppZ3Z/uFnqO6QmSl8bRZk6TDzcWk9UqGoILZW
5NzE19N35oBAptj1UMlBY6dqt0AdLgg7MKygefBiIwMCa/g1c7ACb6H3c/HIHcQ9uGUWvZJfhlaF
xQ+ZSrsqCGgLdrx18iWzN2G9TolO7frskCDDcqWIpmWfTzALeS9KIF8X/YKPMibWGV704mbusSOp
WVbePhCMz6/49Xl7WXn9SfPxbMpan7c7JqJ3U/EDwBTxczB9CPXuTAyGlKwFADJbgijcqx7m+3ti
cOlAv6jHU8YzusO6PUzckmOKUyzStDmMH3DIamUV1bxUv6Dt7/tAkjlJVw1o8vrxKQy3A/L5mRUB
uiH6s7JulEwspekSbQ3Nwq8UpXl4swN1ZiXnbG0DIfrC9biCoCXEH3UDKoUJqvJjEjkGV9XGnIDW
rfi6JRQICCzu3ch//7nW+oPtGYkybPAfiXs6rW15SB+esHQ+tS0OYdBq2FBSk/jWyLrGRPnr+Nke
PRUllQs55/sHFAQF6BS/bPPIK0sxKYJvHhGZxrZeyclFxBaLH2aOgucu9BMCLIp84YfA+ZNhg4q3
o5YT67ZCe7TiZmYfVA+1SHMKCY7CEseINNsSV68g2io96oM0drEPI0NyCoYTFpXtjhZBiX8xRbCZ
GjaAewX0t66mfWYUiAPEbCspTZtlsynE0XcQT4zb9FuNaRLWUvfXu9A0WSkA4kyjM2gC+VONtWIh
nrkjQxpJHyOnKQpZ5d+9eUpI0S3Fjpal2DnHUBen3KjGWl3jnRLHaeGsf3elIoLlVxvejKTt8G9T
316CId9T9LMghxTe8iLlPZbMIj1UDIwbl1CHgivx3MZjhcR+sGoY+HJNDvErdaGJ6JYA1e618wtO
PCMfL77jO6zdt1olFEGbqGO9kt55Tphm0OfLp8HcXhIhPYSKa9EglJkkfzIzx3Q3CEFUDw4v/cfx
M+fJUvyT7Ty9b6TTMTkGd4rI2B/1LgsiT4ZBI7bV1La3K0mYPewpmYWRhXcvNN3xhDxmbUmfP8qx
TgSsXYdQiF9jdjtZCu21ptxDSQC6wF+Ojj07Xuoc6jNftBGana7RTEB96z4xVXFNTaNz7UdbPKMI
iknn8XXH8ZoFA73RgOdUF2jgpAchYox4CwgE7AKC55XmPwGNnxrH5VOJb+jtIONhMm85ydxRCfct
pGsc6QWy0YZvYz49ZhdOycCNWmlkuBytGKxOAZ9zjk0dK+N4l1Mcz8iGAD/+UPsf51gsG6nttNrG
5u+rM/v4wioP/a1h/kv4gA6D3/mEerZHR7jntxDClOGLgdgo0tsOJhFZBLArq0CgkPdOHI9zsYJQ
/tBzP7X2n93+F1HnSH6VIQ/O56VO+jJUykcuEU22MsaqXo8ILvcPRVYCr9xzuUSs8NiYVoxhO299
ApwgHldvy0SKYOWvYxidA5FI9n70VSjVl6Ngj7TWB7T3goeh1aO3FGJ/hNFwzk+99cY7DeBhJcoB
xiz1cF8ZQeKgIikAy7dh3YyrVy8jF2BOCpzlVIcz7xQpbb8DHoRCmQQwIRoFLbaDTMu0kch2FETC
Ppnf55fb5VjD3kHvC0Yxr1rM1BQmOH9k9NuMe1gcOfIoVLsW3UnrhQVHHU1eIcZVKbjn0dXN9Seu
AHbntC0rCkoDgO2AecitoYPCaVtQ37hG3NQ2rnqgFFO5+MDBmPJikRl31CcZcFfeZ3If+j2jIpsr
X+ZRZbaAjUzz0Kn2rs+i786575PeJZIkzaK/yTcbGNyFsZRu0GuTMlWihhw0GO7tKdWE2sX6kcJV
Sdj6lwhEByRJnx35GfPpRtpW9lxCv53ITDOQLyM3MdeG4Fps77J5MPXUf3Gr7i9wOlBrqcXYngMY
pezBNbvrwOO+rX4Qp2fFZKtTmTEr/pzIx8PL7laYTl4F7x5+LhJ3kDCXy2GeLxPiJgsgqZI+gOf1
xIfx5VSxQje/mTWBTfI55sUVjjrmhgtURvQGItQ2K9kKPz7UJrzDqi4MBdqy+rpjLOXUbdwQIYuw
0FRpw2r55nJaJxlhIoQ0F3dW/6YG6lsqBgX6FS+2oMndOjYDUSKHkqfCkk3tM+80giYHS6TrY/rR
12/iN/N/7Mz/lIyAPb9RDRxe9lvUCcQNw7pmYfVjdi0zDDEuIXJ7BRLVlzx968E5x3eMPTVMwW/3
bf1RqzVSStsAPZdjV2nFokoNXmPifqBDXFRLChoDh+y2UlpoxX96CtjU5XWLbUevdy96xDctqiSi
yEN2KlB2fM1iEJyokg0M3xef8iXya+1qnIWcQ3YqJTR4L+zbN/zbywn7RRK9Rs9Jh7ariFM3WTay
/O/S4rVSLLtj7tRiLiHLM6wWVkoH9znVkK6krQNrXoyqtwHzG4ZeWyLDsmQMAQTpJcN79PU/Ds4l
9GkNf7PlTaheV8pH6ZMkil8SG2kMaiMXyAG2JLGfsQQR5x40tPYTJOFnEfcv/gJEtblBmVycDige
zeuZlKFqWFscfH1GgLBr8bRSOJxhpGB0qlBNDYdNNiuoT1Fil3Y/XZyAgFEQZkMIsn2bUCuHKaWq
HEmLIgpOfqVG99wG7nEkJKlay72yCGFrTwub/4uDqinDUZRqIz5+wze9G1ta5B2K5VrOWKOXTjWo
GBPOV0nUnzmkYF66v80rD5hY5nvB8rWlhlI6ibxcEs0Rysy1DzWPdbKCoYDOV9j2WXNcpt4r3/p9
wtiKcsA3RR6o5xGT8U/TJZeoNU6axR5wH2d3bhodWijgUc6V7mXkKX4IV02M7DOHIgaljhB90fiS
9KWXuKWMvPQwDXLGk9DlGDPm+ha/PzFI8HF8VlkvpJEGdUDtTdBwfodxcXGgN4k7hOpTlfGG44VX
JBRaCDPjF7WzHlBd7JjJ9vCxaky5TZeFPyRTxcpYzzGRCpSR5RXle2T6D2kx/klekadcnAhmXO4z
FoFF464Arccd93gFHxCKjMJwFGERWLewn5x027qSSNHMiyltwZ5MBY9JUyPjw9y2v4vloVQRq+sY
ka90t2ZdyDI7vjoZnzdiAWKPf9lvTvxp72oyANPAC+SMU/i2ouaT+6+aNrS1BtdOBCktznXHi/Bu
dQWJAjIewM6tRDKo9zI2Z+5FJQjEKz0PNWpTQT0locCxf4CTwTxnuuhIKTHT7WfKWDerjAXe+Cgl
7bYfg2ik7z4pBsJUMRCdinFiOoyLer5zvx09lT7l7xvuMmj+u+/gSM5B8ELZ6BlmekqaV+uAiHuP
KJsbRA+Y5gK6YeSj2suhSonNxuFCpk/rT8Nd8L7DuK13SHsnFC4/Kc1tUjt9RSbjgXEI7uzUZyxz
k9hCuBRXxJQs2IZO9thUGPzfpKnBLrDmG3jWKU6+7+9RMbokfDEbgjFdGNzBy9r5V8yhxGbKWpL8
OUwpTs5xUO5jN1nmzakLUL3L4OVFqofwW8Ieno6LnPggxCNj6zZi67/dsHONOUbR7sEkotCDLkx+
OCN/QcosmGqik52ImrvThBPUGSR159Ggk7uG2pmSoEhXCyit+UsJFd8u1bqM5TnZzBQb8Ki4luQ3
ZxIJmRr9eOspjrkw+qgpLUdL91/O6/3eo5/qfzb48n0Xf/ZIL/fDjIYO+904lbmysZCU1fXxIErz
QNHchzT3s7iylOtylk1lM7wzQ17MuMguHiS2IwTSfI0ZW6fejK1a46yFdkXJVl6hbVY3zwwcFeol
Fos7loADX0g7HzzEt0AHXrvslHHEYxo/j07490T4eQAY6H3onepAFesDPWA4KYQlxpAUYNm1m3ch
7xBj1jBK2edzDvLxbttc6RF4tyDyYtHdcmgdtFkQ1bU9oZCk1HNLTq33VPlK/I4qbzjNX+ZPGVqg
k7kbaLiikjbQ0/iv4DZjX6MEtWYo+O6wahHXjey7EQaymL3miAymU7eqURGojMySM/xg0DuD54qP
cM8vCTMef+E2EEZvH3qwL/VRGK3lYgCH+ZiAxJS0zmfU63Qo/rgMzZ9YbgyrHmXNOX0p/gjsqCYH
epyitRT8UUPzGX31xmXUxHZcpzzAk01Z8hp79Mg+2Nh6GsQyasBO3fZ7B9EBkNFaNbj5OhGY9dg0
szBKVzaF6n/fE6uqFNzV2lsjfVarE5PVqAekj56lQlPS51m8SEeZ7uzZjQwEsG7zVv6u0q/5E/oG
8kkJKlxLpTdzsIE+XRDXgzFt3dLJ2aai1awQtZAwxIonKZ2K8Vg/0L5pqcjIm6sXS/d51dMifF0x
0HyuioY4kF1u353T1UuUMQe/MsZUCeWv67+SC+iaXiihA+RuVA2CtYQJvc5tGegFVc3YpSALvSbW
W4LoB5Xvz8L3zrO7a0KoAxbUUr/DY57E/C0lVsJkgkTLdUHjsxxo+ezp9I9TUide2cEjoii+xizG
l3Bu/ClM9+74E2CDn1UBSC/C8Pfoj4bl52ERQBdhrCN9p8dTnjQrOQmXF/ezCTGP0IdkjNvIPf6O
4RfSS2Mm3kOySlxi47sLoy+3gNY/HmMFlyxXwG8Is2ETeJlNfiQaaRNyfox+XNi7HPtagdE4UlgK
FNpm39dnopMEHmxNghEJ6EmRT1ylsbq63nbK8iKUTCiA/JZGBjEfynyouIlP+kiz5/bSMIVplgdG
AXbEN1R6I3qTlOala5j6NccgXZvUyeP+b5wvNgLQYDOo2fvoZcZsYKWVxXhqHOQPJUkude7X6llN
BKczeDhn+1GIEjXKSbRsUlbHnFxfu5QBRU2oFACXoNAL/wE2NE6VVEUXcn8myyAn+c6F9xCKIKFN
fttbPOz68q8/bBuBOFY0BN9wYpHYWQKnMYuRm5F0QBLBSwTN2mmv0hVKppsTlup4vuUYs4KlftYH
mhAvkNuI8Hnq/Xbxe9TBP7XsO+h9qSKvFD3vIZL4b9gvQ3L8/PcC4pgxN8GuIX3v5BJIS7hwq2aO
/iPCW8hx/LeqbvnozcW2f4P0hMqElfYhz3djXIkWo4RNBkjA9eCX7losWOZPTkfa+K+ogW9BiLIb
xQ5RfCl7cNHx1jExv+G0+mbYCRwVLoLz2Y1TVewMFapg+3207uoljy5uFOiPcti8AZC47YQou/9N
5+gPSI1+gemOWIpKaryJ0tesJW82con7pGk0DUWKIkkOKOe10zK8dmPYwuZwmv3/zB/Oi2HGd/hT
dWROJCtyMf8nCgOmJo9E3BaV7tYDA/5QS8MXxPwSgFXzy5AEcD7eh1ZiC4aBTkdahWFZxW+JsECO
Apx6lclHmxQvY8PvjIyTw4d2JBPubAt1miqQhX4Q2og760lTUX6ezrhMGAYQGoJEFovmGNkPEk1p
9MsKaTTM/pOX9071ken7uqIq0GqHKEfvrHJKWEgh+0WZq52aZqzNv6Q+0efRV18wDSnKl72LX7Yp
0OJvwQfg8E56/8vwySapBVAxh1xylyF5ffFyJ/LUMFWLyhxl5lzh5v1y3g/rj3UeoUU7+wnCOnYa
PaUFp1BSvfZYwj3PuqimgwiPX654LGzRgXp8tO4AU3CB67yCPeTFxI11nM2nqo6hvnKBBYQxzCv3
lNd+V98fcMT7+vpZPPdLmHbpP+jXRj6ik5ptqmlyg7hN1nO1YzJmlwiuXGisl3NDnNUe7biGV6qY
L0HndvPyXxCYq4DHg+z0OnB7XcruOUO+zcZEECCvxd3F3ANDCuiSMVGKxGmdzn1kcQDfheqfueDg
r+WtXOw6/sIECaaEBUVR3xbFgxXo0ceouqQOfrC5aGnDAZuuoR1C0/x8sJO+niXDzJTLItDI46bf
6LyEJtZ08nnZFz0S4K1x7VbMUuvSnZ96Nz80FHQMJaev5alED7sTp3dT8uZR5dNicjJK/GJ2DIv2
jRRdMVNGDTQqOSz2Ox94jqUBlW9btMF/BBra+Q1YWYdvWR4F8YijYINBnK0BAtwVHs7d5N08ZPlv
2mwGX9DNj2WBd7EhDRl3IUqFSZVE8rsmvv5ky9D+Urlx3j17018GxR0+Hu0Jn5KgTlNiLLxxEtn/
UPn9RcNFn/Ypx6p9T3yhyVotkdg27X719avqW21WvaGcKXN3JF6mKXFWtxEDiaetz34OAKRqMVYU
7BHo1GHj+PYpjLk6DK/fpIxw3TNGEDAMXeUmiEZxLjQzRKqHskygxOCgqNE4iLrN7kPzbNkIAU98
Se3ewH5vfn/82aHpcfHY8Gcu+t+ageLO6v9LEM5Ndy/JVfU69Uk+/pfkSup9hSwJcbF4tjWsz1Wb
rUO1MXrILGA1FSV1kRdXIQsRo7mWP1aKydlJRdZ/GPJ7/hfQhK/bvbl2V8j0LhxG4o995UtWAEji
fm83ciGZH0kEA9y6/YQfrbsr6pSJuQ3duWcExfGeBI+8zYsghLkRTeeLQceZFr0v7Dv9gUZKxPLf
ykTcWTi90TKRH/OxyBxUu2+q22XEVwwa2o0JRnMl7bhgEDActNIdlfsnFnIZwJILZWdIzge/KDGB
JH7hF6jnA2dVXsv+nhbTHF8SKXLDyP8OLB3X0tDNQrrLTizLj0a67IejMMerBoMspJo0lflDwowJ
zKtzLXapneL1Mrze8WtWIScFWos6kI6+b31Yphj10fVl+IpFIdZnuBqNfXYDYrIyRXm4Qi9YrgJI
LtsCc3/quL3jRLBF5Nk2qkxKGxcnU9YD4YWMYhAYcJ627X1nnsIqUVoFRJM7fxU6Usa/+mHPHwvW
he0FWeJrH2xdIL/ZUy+o0YTvSAi8KpftggjftZI+RQLuawB1KhIQIPXrslfGg8VxM2xtFFJ0pCYI
Baeh7qY35vwiRIKimTbxF7Bk2zx25VqDy1q9YMvVkujJrnUNUyXW5oITb4OO2MLoJBARtP05x7r4
jYDUnJfoaYUgsCB7Q6oGq47k4tz+JzmZLvO5A//oRQhIcxga69Ec3VFPCUwC3Dd8z1AujHF3fCqC
xCKo9Yy0waJODvg7pSWaJUkyiSXXiiYpe64qzGIIRdUvr0M7LSRLnnjL9dlS+DPV0PIvsga1LvSE
1Kq2zeBl7x3Y1aUcKQVWF46voFLEeS7WKJAtOhdUMl9LGYRaf1/6La5cZ0s3ZPUMMEvmE6ztODMD
Tv9TmRmsucF6kim044Uq+ZSya3oyJ9uKqZytYkLr23wQgMRewO/x2VPg/AvgcYOeTfzBw8S4MMXI
0bGccgaGZsbG0RWRhCJsx6qdVQ4ssumDwxWn4UgyvrMabzpmVKz2uP0O0VOPhqeHnakpB4w09gMC
xuBSRSTDwGIlsVmHjNKZo+Xv2ZLew3sjdxj1fNIjIIAyyjiyhjrUW6x0g0KpA6H0mSzFACtQ0IfH
O2SjOJ4M3AN3UyZDyq5Ae3ldsctZHd6JLWJP2cXU489wUXQy4aw4sMSgkXZ9ilukLpuIajqXV6BP
NKBUXwo0fbyd3a/DQZGi716UyeoVsmcarbfpWjhpkT/zS3geA+DcdwdA14tKcBu2//fw2DJJ0COv
uYfZZp5dId25Sqld49s5zUANPetoQ0OZt+tZd/qo/c8T5IIY+Sbufqp+acFSBNjU4TVpaYFtAHIq
jjh88xyQgTwTEyshYx5GLi4EeoOEYEzPQFT0GXaAfF8AYRqHnPPkj9mb3r8GvZOi7M4JGYps1Zls
D1S8aiDtkHtwjIdD8mji8lgNfIWTwTMSK5VFYQlSu7RZ0k1k7Iknu3NCJAopKGS/MWEq9tfA64K7
yzQ+FfJ5c7acVEVwBaD6Igbl5Pe4E8H6leslJBjDbrLZNhSptwf/zcU3aYmmeQoUivH3vub3z73V
qQzbuXVS+BdAlBMrv+AcHkux99X04cZJG2OSHRFF32dh4NMX15UMIVqaYDw5bqx1J/1VW8LpRyls
+sCNOKQvvco7N3BlPGQ4MX/3X3E/O8WKAXV8Ctv8qWB+GV0cq8OfBAKw9Q30t26zBJNV0EaDg/Lc
a0hsfnGsq/jczsUK2Q8QuUqFXSYTQPsie0eX3YcN+dVixWM5dGT73Qfb2OtApdn0qabQ6QtOgJig
bbZpjWPB30TUMqqxYEeHwXPMBlARXn85AS/giwCrBJcufFOZ6bO36nw/b9mUqQgXBJSc1V68AXnx
ZBoaohSxqVW8jLjKfcUlmB6JbLXLf6AQ7VgVbnV+1CE/TUvI3YLDzw4hPNAq21Y332XZcBIooVFe
dOrl7oXo0W0VXQmSQny2TwNEHxEptGSJpYMYzDvfpUsJnTsMIyv/YmI1gc8yUnl4vQLowuCwAdJa
wugEf9UHqjivCgIA7nh8cWESnI/QXeIWF+tQ2swvbytJobmpBh2k2H3LV1jgjoZTJBh4Y2YcWgDe
hbDn6AfZX72jB36ayMYmGMFZsHIPP5tZ/Kb7czSLlLge0S5cP7AZFnSeIuAZGmgFi3HO5UUH7rmo
NFLBw+ZS6fpWgIqCVUg7cotSJGGpymOnnxP0LCIJo+pDVyH65TbFLluTH1EF7zytWp2yi2oNaLnh
DtzOW/n049uVZZskuWVFqF5uEAZLZo5sxYo2IGcROpqkiEBaTq2Z7EBp3UWV+zMHvFr9zkDMHHOg
P1j5Ea1cozLQUkcrJuTy1IZ70Zwnd4fu+UcD+p41jOMyo+WF39WZwSnKBmuqgu4WcEGLIdwdzWHV
HI0hB4YKJeXc71QCMtkSCVqkNVPVpiD6eC14q+DrgnjYgyq1Z7OCY5nEzO+1GwnYGkSx6lb/E7om
1YkMr9wDWH9tRS7kG75SLbOYF7p3nKz+ODdll3Y+E7kpH8hzDnz4ax993xfj8XvLjki1cXTFJSv7
LO+T5nemF29eldNNfC51uRKFLHu9uk1LtPrpBQBhxox7jr3Z/RFNLCFh3Pjq1FKQ6BKv0OkQ2hWJ
fjTDgzIcLREY0VIqQotHyzhTLC2dzSn1RiCz93weCI56wRPkTt87twqGJz/QsVZMzvchX9v6GvRa
I45VIXu8CgcZ+xI4rtYAxMOAVs0rnJccOmqcBz6Tm4SEH3S/AwAuYfjtMG8iQCUElUJsh5Q3kcxV
qWliGKb0yJQC3Gp36Jr7lr/Bkr1z3x5PoR6hNZekQj7LbxUlsZ27tNJHNl57Ev2G/wZXa5HaYune
8FZl/gNpySlBA2AApaWwdAUQnYGpL0mwL0d13wKjJPl0DSrPjoF01RMqRam5WO2XE14/SoTW07Hs
riora2e1ypLl4BISQhsRP+cmhQosFF7ElhvRcfyQc0iZ67kRIdt99Elc8YJDsD9XeQ2/CTe/xQWW
f07qos+ipYVSIbH9uaQhpljWOXGEB49ZEnq63xRSbOCgdN2aRKeDZ7oyfTdw736+LX+MUmEuEJeD
jmC84VdPtJAC+iGp4ddmYqfkG8pzBz61TBcLvn2R1ZaWr9/aoCl5Vog1t7xdMcICqlogZIn4hnMV
8MxHerOOwbGMoboK1d3eKIGmrDX0qrC7QaxMdIuWIH9gsnXaDx0pB/qryoX+acLYhGPCTCfEDuEe
vgFUkXVShH8VthFL4KxsiUw31joAFDWVEOrclZHHIUaKdrsDxXDLW/njLdnusW8reoRcoYWtJVSF
ovP5X8S5vqYHw4NP9xvkToik6Y2WIqwlPbTs+3y71D7F7804nHTWSHq9H4R/l+Ne95O4ZpHl/d9e
gRRS/yaN5py4kKkxG+jdvNWPWiGrvAWy5yii07U7LiNuryCQG0/Z59u5f82+4ScM1+ZW1nhOHEVx
waxU1A0i1rRl+3JhsgR468wRHIMpez1+rNLRPEAj37CntbiLP4AD9q3quRnQ6sAD/jvc4YjS9xbc
hqSuz7dp0/o3P8uK0/uCZ3cj023RfoJalq9x+4YoJgvAFdKw5UajpqZsWF58M7YoL6qpqj9AbJgW
o1mYAVa13J/2bwIHiLH3atUq/UGWtkVB0Gu/HIqhbZefUQud2+z1YMIyjg4jjEu7zXuqB6RtJpH3
kVynICj7tIcuY2UhMu2dp/iBJd82MTQ6TPp4QBFK1tUUyjntwygb5mCrIh/X4Z7HdRNvNrWc6zlS
ICfeq/9qUs/4SOZvUxN8B6VUMmE1R3HZuR94oK92U/5HnyEz/FLzTxEdCsoKUgFnp22YeFnPaA6j
unG90fA385uRzqu+UrSLwwGuWibQWcUaXbki6ryobJYPyxGIH5+oa47fAftaN/DpyCBYsnqtxzn7
2sdEeH5oWuVZEoUEJceRvEXyWm2Vp0w35W2NNhB48eXw5Pb3JL7w/FiWOw1ULMl4a+JlipTTHVpQ
zGkdyiautgKj2IiuHJxnUGTcj28LC5CI22W1u5SYJ4CUZk6uoOcZqhFbUTntp5wO83yoeGgQTqOL
mFYt1vq5wolhF3jwT5mGv0ShLLKLhQUhcqljk9Bt1HJJ+NpvZZZj3ptrVUDyPAreMbEfT4qRgZGh
xedyisiuDRX/7q87WaSyskRtZrB8M++ejlol+joOJABcFd1kx/M8A3aBBAVXzseGrJp8GnS0cnXO
C26SmtlzKqx1U1nkDLkTNaBCZRLKwXLUNSWGwR500c1T1jQ6TCxfBVpxxgAd6tqH23rUqDRV8iU/
GgDwjveeQrFSRS8nKxXLq3mGQusUKlcwJriWRy703ZMdknwIKzC/JJpHvmMK6F5pbtDqc+AUl1zu
yPPuFS3eeaFrhDcL780+b6Ol3L0y5kdk1Qpl8WcZAX0JyajyL1g3AoambDxqpHgddF7v1HBCclGT
bgfX+Nbr8heYRdh2ElkiTQLM/KtEUZATiWOZ6myd0x404C4C/0h50aY5l6Ytc0Oth+brwMH6RV3c
c0wtefrDscOao8IoWzVmIqhiApe/ax+kGn1x/CFB/Eayzg6gM+kInKRYi9luNOziaBAaIAwm8K+l
55+xL570vm9DmC4S5Ukq9T1hTDVOAQDkK0QYHUWW5dFshuKwfrReAFy5SJYauOcmlvLRJD7NqbZj
TVTCGwY2JpXZ8lP+CKEq4I3n2US8ZJJAagqyTLBBbFEGFz4oGjG/yoroXxe21okMoTJVEY/vzN2q
6lDPvLTXqyuh6dorjKiIKJ/lhDuIG5uyzHz1du8ipxquLhdD5r9kIitTJOHwQDGZsK+Hn3nQpEFu
N5Y/ubNZR1qEjhB6BD+6feUdgggzJ2eeZsxe0BPpPkTA+nfPPt3OvoncqQUZ70bvgW+aTKDBDyiK
Wxx4CQVUpV5AGo8a9pyckCnLI8VebMnBfdCC8GSPPWTRgyamkWjixzN40XNOmUD8s+IM/fQCXKd5
8tK1hz2HKhwuVHPbcVrZ3EVtE86aOa8lNYUGInpkLCkAPasOq9XlYDUcBndLMBMKerihMq/ghrNY
XLTKXTV+B9S8W7mfwHVGFRWpFr/nEpKL+aykGlGgNH7eTmoZFeLfQvr7PynT7hqTnxX6kpJpHiSX
eNjOVrhC8SrxmObgGHHeiynUIEqWWkUHVg61R0k0u4sNxzhE4HNSPXJnhQOIybai8aWyfAhQhVA2
cZvIEyUeLgvdIm2yYLe49DqKHpV8x57gkG+5MTFGxLIQn/T17igdcuk02YfgI+w5h+3kh590AF8V
qd4lD9pp6vuopN3nlmUVKfb+wsTkpPeL2Ae9ZgWlOOioQ3Aphsx7dzLe+Hpy9xYTaL+b5PxPaIeF
2ZY0OYlg++nn/YIm0PQ9VE/sZP/IfajEXNF1YcN8LfrPC/ZFRIVDAk8+4lB4Ia5TmMhf4uJkvEhP
PmqraQ5F1XFT5KWfsFi0mITLnpQpLogWviSWRMhQNnZySqjIP7d3IIXLIYU2RH2ZN1xH74/H2Yg5
67/3JugOa+ypbtdytwPt7qoXxomV9f1WDmmX5X++/fXFWRsPZJJaHF7V7gIK9GzA7PSfKVXeS2uD
irx5gIizvEUDT0ffI0RcUaysEBrzruxGxzq6JXPKa0PGPu+ZLmDRLYDHqIQQ+pAFYeAOImcTf35N
TUzir2MavsMjRof5vPKgwRgClzJmAivsUYpcH3wsKRR4oVn31K67nYGd/MPL+eWsxl8qs+wdM/Xk
VrrgI2w/xVgtw9G0DCun8TmogsUt6Q+tYLuSW2pB+PXOwSoGQ4PYJxWWCvnNrvyCIy4t++Ox48Pl
UUoMXp8/Lw26lD8RkNdAWTek4akRMdSPRjPiKAzHc5fnT73MWoRC8Mhkdq7JFRGspPZs+9AGeqtt
9oOyKjQQrW7czGb8XPgNdqzexPnXxiGTuFCeY11LivOTOebeuwud6pkDn7bgtdJDlkBP64fHuSVi
OQZ6jrvA73r5GncY5yluyzOYFEIwjAVJq6OfBw2RnPpbUCCG+soRzVrYeB2UKNAgE9k0DQiIDHUy
33cyj/C6jxLLZX7ldEnH0/RpN+8eBKmoxrt0FMTSTE+kAG/kAGvYIbcz2QkTR0H5fC4ShIPtZ/wf
JjmOmfHmlJADESBG4MOMAvRBLOOjDkU6FNwT8+VmhHybLbmjovyLrQV68PhMKY7e6TuJUisF+6aD
ILREYObpSmjNjg7RXOMJV4TLceoUsipHX79UzlDeyjoPtEzmHjaQ4WCLtGprGRHCxJ/dEKNnp2Ya
HFVGBtXkvbVsRBQQA75RFfk/FPR2XQXV2l2f39sNsuZXA270K0cpPL4Oc36bl35loDNO1mqUNxqg
d0Clxw21Hh4Verk2G9mmJCgKyS2DfkW/EEYNrilz+kJOThPnalJC00tupTHP2179QmuLgpQesXQb
Z/1kkWyBqd8Hb0UG16Spez2L737b8gcKb6Sae2OAT9T2MuXTWWKX77jtehHz8QCXz7HLZIi4LqGJ
Vgs/5QaWzA2QslAffXr+/Zjq38ZX3ActljyqmO6bxR8gpd3YBW6RQGGcQgwlANqvkCM7W4eBuVV+
5UGkeZtN1rOshwFYGYvwPHiozgp8v9UTBw9h43PQfItL2p2LWezkpNvqLvFzQwXCiucfxym2GBe6
XqUd5mUkd7gFXYoRVNaMebuuQxAIrmvDpbM5QRDOEq3hVAxv/2jxqJL0L6ZRyUZWuGTXCMYTtfhw
6ninMA9QR9dNRzPvsI+ox1MGWJsLWbR2l1QNIAxz0BEvw5o1mBc1wMFE6obm+ZGaMe46MxTtKalE
665NS0SapnI47/5Sc2WMlmKUg0RmnwsyAW+nVlhW4zgwXbqCKGzU6hk0n5k/68OefRwzniAeZUdV
O9uq9kUos6YX+d9esv7dYJM0MpxeAgbJuFxLFOKYC2iffy4I4WSEjUGZtGCt4EtCK6anNG6L6ayR
VBzvil7cIDxRyFeMjSFDWR+E8sXIVJj/DFtuAtlPRjDpLGNgg3xm5lgbnNpTZ6i+mR8+NDrYwe/d
pB7Gvqcl8ynxdoSj1izPQTq0xZbHp8IhRj1RXpJ+IHctzsp8/Wcg7t+8RDU4680FOofpvsphuy0j
H3ghIEETUHc+DGz6bUDAVqtzUsYadOSejmFlYKIbTNL0/X8U6LdpVXOkhrWTdbm0uAPyB35rIaQe
M1vMvHRtT1cP4kVv5SZLoyFq/TCtYYn6dC4oNU062r/Fd0J/BJ3AUi6wQACkzRKf4HEz+Lv3gXgU
PsnHDdYMKd5xSNJaX7N0pqP8Y0AKmTMCyaILST149cnCYXr+Cci5yiYJUVwJMdr4GZXdbtyYQZh1
GzAM60e5QSxv3JpWvuuYjIguldRHbgZrQDoFveaJUau07AU365qZoIZRTvyqz0z/jdPrEn5Ys4Uj
0LtQxuXW/w0MkKYdSil8zGR4H9g7LuhFdgCxPebnFTGjEerIRZ8wWLarr7ypUqGG6ym7KwFWS572
re8gtdBaELJG+Ma8m+WqC7AMmG9PJ7v4dSps4x9JRBj1ig9IdWkehyZ0PfutF4uAhgHv8BuKDJo2
nEOU0BvSw0bd6S26UV4UlPYauczUtiddMLhKznSAWvBC0IpM/SyWHI1qK+FsasQamYXl0QQOL7tt
6zeZf571Ebo8omJsIVhFLIgeNILyWBdy+N929Y1/7iormFbzjTk7Jw9DK0mab/lsAWxHSGYWI9lZ
aFiwfOgg9pBwjJ500VoirLXaP254UUjt4KuR28iuLA17NS2sdpDrX6UMfHOi++wItPgYCNAFMMwV
bbHVTNZEKK6pa2PQ1l8WFJKJZgXPnlkIRWTZu2aYwt/IlXtgEHsFgEWDpOMrhwWB2SwEF/quKsGd
bin5Xv6tRcBJwih1WQKBTq0V1u/gsvDPBcndNA6p1MwD8EHzJUlnICOnZNEoybU8tLw97vix6PPv
jS8c4S39MMplorWGK+QyJklImrSnSkfRT0wkfF71rUbR8jAOVXfm/eaBKgF16fLV8sv2C6CAV11H
iaEinztCu7B2kzhEUCLu+ZX4FCbInq5nNiiLvI2XOIZjzldFC5hX7daXPRz53phb7FubP9AGVv1F
RDqsTp7lqAidn7nkLBxsmf78RB+6Mmk9aVfcj15TV5Osz2p44tcviFUrx/p++RulIbN92hhgpNSP
z03fqPvmf2g4YAcfYC1pdlfMAvpL4Dt25CVj5o0hlzJUciCmdBEgkhLSNR2PQN3yxyiZXTIhK4yI
ve9bs9Sznf3cpGrjKI9Z+6pWpFgNwtS6iqwYPpgCqhK/gtLMLFdqHtcEvuN6dRaZ8LlTZ2DIuJ5B
gPAs36VjUpN/rC37w9fXqsCOBPgwZzEDJYGeR1NKgphPUslNp5HsLuc5iiny9J08DpUpuUs6LtXm
5FsWlb6Bh0gwvDwroKFj5FbThr7H0Uth/d9bCvqICftpOKUn71+nhyvXes6/FZVR6Ga0ILyeV/8y
cPuxQVDZQ1/PqeuYorWYdCNWHJOohvWapldYC8qIjqWC08p2C75sqhT7fE/8zPLyA2cfiPsuOgYw
ObVLsInL/j2JkLe3lAnZZnvvcsW/xePBHQTWG0RAoFJkdnoRkPmY/G1pav6rPIg6hNtyMeqKFZbl
DyokDJYp5p4RvUM+HesxTFEU8Ner7jWaGUPV5XbmMqv3YqLHY2G8HXyYypBJBETKqYIolVfHsDo4
BW+uEbv+d8dpd683pORO4dYNpb5OkhQCa6m5eDXQ0F5HIsaRRgVBSwtd3+SZJXwK0t1rIWPK2hrq
Zc5HBt9UmDy6zDbHAwDoZH3p0AMNdTwiXvEmcDEW8KzIY5/gxHvxMIXa2J8+/Yrp99yIRS3ybmd2
OaEc5kdEWjLCjQx4muxVNCTCUx/+k+nHbWtD2fv0wj1o3ge+gLJKikNoXKFq0J3IUgA0oSvceumY
3fwOKNsh+SPhayqlNfhPUciNzNiHIMJAIXsTFqLQwlRPORkLplgYPMevMzp9j7fNCcj19Fvj2d+n
xamj4b83ShlTfhh7Dw2MZTrH8n7QFKEDCTT5yoa//wqGa6uTY/p/MGbIeaQbqULketxKY5rksNKz
b00djHuMvLTsAht7s/h+ed4Fzm//HK5HMulKeQ6gNTdmqm2Q9AeEywCW4EyGFZx2p4Q+tBsnG/Mv
kZZDF+UZt3RGw1UZsUTKpZ+o7j0EsroEMhEIV7U/lsEth5nByMq3G7HhMTRIGO8D8mZYoXA3DVs7
BaTHnqwZ4tUJLMW/BS34sjGC5AVvEgTJMqg7NDlNBUR2WM7BGU9AFAe1AQnPj0pM1z9Yd+5HSZfC
OIyOXS2T3riq/beQY0q/ncfaMsa2TelgzvGJ7dHY3eN7Pw/fgpoADyoG7kRIOFZwYl6j4Zmaa/Gh
/O0M+3ApmDVoJZAea5SmS/6cZtgc9oGD3YXOuP7/zSNqNZuu6yb90DF90QJNmfci5BPd5Oe8wx7v
GTYyb9ZFpftSocWNCtvmYw14fmOS427yhrZs4RG2w7TmI9nI4nIKVf//dsEyqZdC91GK46+lFQ82
76GMiIH7qS3Str0FmAa2I9UvvfCFef98pdZXDpBnjLEoTY1oLXORMMglSDaiasn0XorZJ7uVySYW
vT28sxRXnCYhRP6lUaqGI7bKRd66u30rUl5a3nCzPtkub3M5Otqlf1wxyEgGo19+QlptbVeJUKfO
nP/xDO/8kSsULLr65icrD1MtuZy4sbXpTFFKehux2LFsMsJ0ONWqGVoxcztECqRC20cxmCXePR9k
mEstH38Dk8kOOgme9GJX4WRDtAllZg8b+anh97ExNUctAvOTvN5XOOQjPc6eIIPUUAKm5c88Y7ia
EIoN0hE3F8i/U1/BJRtXaV34tGenFH8B5jX1QGMuhQAVqYt3aLI6zy20aZpBrhkLhov4mIaqUfNB
7G435PT+gyK6Z3MUrjj7qYj/yLl/2tpbMbAzuENmzl8Qy6sGjnDdY6l9SBBKHsS2HL7RBVUdwkRb
mkidcBQXb9h+YAP+yuXu2QVTLYDT98JDZyApufhtgyPD1EXmrUnWNYtMWjtfBenOyYVibFs+KSU5
KVOHaojwUap6ENnXsqbSj84hsoO6Cdi6h0e2HA5p77OapcIVGbJ7V+0kPutDGQZFgVHJFGcJAelz
G20s1ozsjp5kLdUse6LJDGXhsG1PoLJxXV1Vo91yttIS4TtMtutKlMSTjMPGEDkYhwHJuNvFa1K4
7DQjdcv14craEftT8bfZBsVRaNfJo2HJXgZZesu1QNvgkXOC31AFDpBqb8AsqTU6uqh0/j7E9iY7
nj7BeS9GHHXYjK1+7lJ5I/PnKLxdfrZHxtPWmDwnfQ8J/GLTxiXxpyUdpi3KpUT8rvh5MPkHH2p6
w7kc4gOXwPL2ywQn7ix+JFzG6SqzqJb1sIfSQ6D7vb9FQD7nYOUOKKJlfbAJv5zVCX/ZKua/GL7l
7IF9Ep47nMzZTGy7sOrV4ekcsJ1KXTWgoX3coFxIU7G6Gszve3adVVgSdMOGGEXq/zYTq21ACib7
1NyEJFAsjDTAJvj+Xiik4qK45yKUm1h/I/ataj4exWVbJiXee2qQWXcnV4hSc7x4TQfmAbctA6oO
wbwB2Lu/f+SoMDzwnpMHqdNT6vF1kKuXKOnTa9AeZV5cvbYyw/OlICcGQ+bQdSAL5HGHbQiNDcpT
QGtP5+89GckFcO8YY5UiNCx7lTu+cnAmtLTZ2R/+q1K9unQys7BQu6XUl8+3nAvdJEWbxdUgpUpq
a1Gug5VOT+JB6hDN2sZBXvo5cn4VKsk3lydFBQndiPJOqPBy+B/DosG5657eNrNoZBAtwa8klqrd
/JTX34BFU9/tFmL0sjMkIwZ+57aegFf92R64zYbFfBh59yRnJIDWWjjsJii82MfEvEfKxZAV+Uuo
oHcy9qJ5p8Y494I8YcIdgwnlSVh9LnGq9OPfXUViw1vmIPlfoNRPd/NUv7lt/IjFaZhcB5O77r9d
zE4crurFajWTbxKOWz4LY9x877Eb00kyEqsoQlqKeMFjYjJTPeATuL/3qV/n4W4vayklyun9mua3
wFswGTiApZIT4/8G9k8dBrRsyhQYiE9ko6HgSzK1+OmpzQlu4RttPIEq+d6APo9OPghW/dMpJO7B
N2flnftOsK2K6LMQlAP9rRg9DpKn9hMgOVFwFuL1M4p1F7B0TEePwxSHqpbFprSfEGmPo0oQboVB
IuXrJtpqM6P9MjQrd2v0zD1z1Sgrrfcqb0Fa1uDlwUK3jmnLKK33UPMpZaKJv4ebKZLbQL6abrLu
Qe1MzrIAUUoBTBViBQpriVQIDeVbgBl2WaK4TS6bg0gZRsknqtnfkdltcq2A+ZyfSF6bswxZ2WZ/
oS7jegKJgISc0QrLoNIxIxvuutLmrVniusHdahb/ZN+iDNXgFvbp/3SqrlmXjfI0pxZ18U+0OF9W
9jZlWCeCmVwdkqmtBz9Kwfzgpb9nbppDIzrYHd6emeavW4zOY2DpJV/qEELCOGXSfZvEiPztXJoZ
1th12C3Jb0gvb4UMeLokFp/pwJJxvhdBlkdUjb0AAhC+qyAs/BYYfkS/qxbincx2drdsrmM0HIwS
KP+VvQkFbRVfb5onPr6q3bcKxqp0PHvJerk2KLyo3fbnN6BSq1a9skGPDwhJ/6iz71H8is9N07q5
nyXGoOvSRd6+RPgEVFXbbRJIYDxnmgHurmTxHgSrM3Tv8izrReKX3s2T5jekc7BeZd994DDc8ZYe
anL7QkhFrScekeARIzvfh+nIyEpkDbLP6VxX2Qt2qRlGneUUBsgEraI6/RM+SPSrfAjlO2PbimMR
apNynIUOYhhKqPzFFjjK2eWMsdAEik/aTXUvpnLRGa4b5S13KRYnhVGnVmrNklclmO+n1oau+ewq
V9SkXuu2VwkuS1VtNgZSk/w5lLn2qAEB5S4eV95hNqksd9bNgr/SADsmi+Ak1GquiD8Gp3S8pQBJ
iq91CliRLocoQ4AXzAt+i2ssyfputKaVHIIMizQph1ItrCbF86UMDGyo85tECxIq7LsTl5nz05r7
pee4koZ2DL6TFkwAZpghJzh0p6Zc2+HCey45nydtjesLDa07RnDwsQgO3+DMLjQDE4+kjTVLTM5X
wyFVkKIHUBeZRK32fAxN1vCogzIfrhYQkJKS1eOuKyHBW3jHH6YuUaZFSuA8ChC3vcogG1umknNd
jHo4yjmB5WOe+RhXs5sFP7zaFAwFpm6JtpOTGJwHu9J+v8iWLRnizfcI+WEf0hFMvojTVqclrBJh
AHi5Nsw+A5YK0/ma+YE2EIvvwjLRxYQ4XxrtrL3V0H/i3k7pCRx6lydohs6ONc0Mvfcuk2i/AETl
HfOHL0gtssx4fC4xtBMX4ImSOkcMkC25DfnBvn0+cWvEsKlMYo5GtblRWI9b64fb9jq++XIxyiWA
u/1niVgFiPkC58Lx8VSJ7bY+l9RCdj0QlC/O+vcDuzl7m45r+ZCqRWbfN0X8xPQsHyfDNJe++MzS
PyBscZ0hK1rbmJRi1iJIjeMkvBr4ecu0xI48gLqKY5x48Xj4vJb5qJQPBETvnxK0fc9Wg6/2adiV
0rmE44fc+tG6OMyQh+2+3vDJT0yFpx/8aPKv08u5vIepB9mIS3b3X5DvQndGtm6gdfbyIogSaQS7
wsY8EVLtTqa6Dwx1DnZZb555HYRjlyiHRO9AZlSuE7kH+w9ADvq/iM4Ur3GptLR8FyrX6Qtqmt+Q
K852boUW950CxC6W+Ab10NoWLgUfDVw+5OSgUfUJFBMMMBAtmF3z1SkwcPlPB6SV/LnBj6RZPq/q
Nk9gem2k0xXMH0sf0udjOQ5VizTXoyCFRzjTRqaMDWXFw0aWRIUA68bV0nZTxs7lz3YzOR6aV0Fx
p5zWKcDuAji32mumkO9bfIQ80dqUmZrds4sCc6xvJMmQvhv18EWD7AgrUDpHkfXKY93UngFbzFIJ
liHwwMOY+NT8n7nNh89jm+8ZRR0DRfUFl3vNabt2/zeT1txO+Hz5zBc2DCoQVLLNzVyeYi4LMWxE
jveTLF+NCt+bktKaBQrMsuOhJERWlQWbyEeaFnO7b9ei7TUMeY9Pp9WHAhtYa9jspG8keUGFhgfE
44VPIl8XiXhK6LTUSbZe4f3xaS2gBBQYn1A75vnCFMM+JFecJ3GKGnhkKC1e9LC11JRgpY2QY+5X
Jyh42ZsMyaScokdO8nhVhEdaIk8v/AQSFms+RieiR2lcse2rwGySm7zUSRUVF69/mfmllK7rBqmt
jrQOVAvwGom00w2i1fC7iJSMx2glQLkXBDVb3j1w+nPa8Std2Wwi9nrtbFL1FDM8a80PY4g0Xtcv
j/XlxErFfqnqCeitotqzHAz5+V60rGnz4OwT1UZQgm2jFA1fkBD4JvjNYROLGBJXH9ciTZkSwKnE
PZCvvZ3MebLGDkLoYF74lND0h23U/dvcqYAtfOdSyxyQxP0foYtRye0vucIfbOpVEslU4Jr6p9/3
/FFLYnmd3fiUaw/c7r7RAyoaq+nSM6Gs24y6VIZLibXsWOTxBoWW+8Kjxn2IhMu2K5160q9VxEDn
x3DyAU8H85quBTnycVqY50/YSP6U/8Pw0l7wllbmxxXUF6yWYhHr2AkCDo421qirf2pAznqPp3jr
jC8X/mkOCOIZGEtIcZXLX+cU99UlHp2aW2oqC77xUyN2gG4VXm+6U+XQ2nveXe9NaAwGY2argiNb
z/rddRd7cf0jPUQ4lt3W9mUPA/KKkbvLv7cb2pc789MOygQ+CRoBkJ5/kqSngNsHRthdLCo0N2hq
gu3ongfTQVaEXaKuVWPXf9wcfjmTp6BfNOcdcFZAhhCZtTpcHJyWc6NQwAl3EuVAEbWKwquAALKs
nHXSLeegXExoDpbnUtnjaIxQADqH33TUe2aF25OHz38IYN8G2+dxttg+Ml+NzEjdadVv/XT7cWvG
sbKRh9uIeXW4poj4e/hhBJ8VBjvxC3jnKubtSFNFc11x++pmBshM+f55rSMKYMzLVjYEHqlEzCYa
isDzlr4WCE3Enk/7xsZGgnVh5pgiRLM/ppNK+QnYVBUSaoXolQnYtbj8iASbuk2bU9/ZDUYFprlw
6yrRTJq79LsPhrZdVhwZkGYJwne0FdtwNNpfiFDPxawXVVyEptXp/mwxzyYqS5mhOLc/hOrKvjU/
WecVQZD4jrQKoK7H28FLIG6Th65gNpOZO7KGQ0/AEY18iIk4EM3UpzG/ofX0KzbGBohgyvGSKg9T
aghbExvPLzsOQq2SnlmiOx5k+NQj+mmEBWX0jEv1w4/+Ul7xzAM+GBBZkC8AlQ74WhN5/D6zpXMs
88/KZY5DkX5VnfZQ0JfyZasFM+8aasS8TgAIu5ac2t9iqQ+GzpeNy41AjyntHrWOZjSrwhFL8dux
VoNqGJYUdED/NWWBSLMdc1c4IaUp5ORK8a5lcoCJRNXEjgyj6+nmLKTCJwVBTR7aWiCqhM2hN/KJ
YAyfwT+Z+l8lV3HIltDIIlkoQXipp3o2asQHZeu9vQxQzsWU/0fTK7jN7NnOsbuYLjFrhl3bKYsE
WcumswscvRYngxmNpRpouKFf/uWXI3BG1ROA0EzGXSNvqvhpwF7B0DlDXT4t3o+LwJLRh4WvwARg
fd+cMCMcdEdYqppHtKfIpymYDw+O728Wpg9gb78py/oTgAcjqvTPKOwt54KTD0JJGzsm+loa2pqR
TP8/Q0D239KVzS8BT4cWzGl/XvmSO8LvYBeJ+idxLUDdNa/auTZeZJ1OCN+XZmNUbyuGNZ36NH06
LzwQ5i7+ShW5HDWbX07wIBBuiLIiA45kAT+HKwks015HJj3cWstIMkdoETBFf0ipe5/eDlcPO/Lh
rt8oKsLoFY0TAx1B1v37F5dDAuQRALlST1zGZk4EtTzc5nkNWVlRhay0Ib0jKIx9+Yw6wagWFDKf
nEn1TWeYttSkiLKxkXpGl9eFnypkc8dWPN+lLsIhPWLNb85PYP9+nDLVO4pnipSF2LxCqbRQEVHn
ommhxgZIItf38SMxk2Eaj+k/xNG+C7Up/1Egv6ZckuPjMqYAOCGOd0V7r8tNGG7CEuLeSp07lZ6N
IiJ+OvPKCfy0uP69J9UY1tzrRxZt5EWpmWcc5mk/OxLG60wM6v8mXmOtIu9Vjze3tz/BOHfk8LmX
U2sz+cIedQ0BVw1/xbDnHp0JliklEFSSBaW3xxm2yBR1MG7kMf+Ptzig2iOwMAaqMa4ZwUa9GS4X
+NDmsQzTB4Shb3LDx9LOcHdTgeuVBs86VW5fRDP7C9Rn7pVuU/aB92qsTrIPpHatxuOmbwR3N7p9
DwIzXj6uJlaenFRe+gMMh+Y7gXfqA2TVBoJgBBdxnbGhagUJB9m0N0NskOVI7fxfxKKJYYE1xYmO
B82Xm1bQ/x4M7P1tvJb9IUpmJID823E96GTFh1Jg4feboMGxR4G2CS6M0MHmhU3zb5e5Gq2D2J7Q
odxU6TgtmZlJERaZgAlKmtG3ksuMKXpsxT4H0aKPjm1JWGF0H/5gVYKWvkpmHrhkQml26VzVjHLW
rvEUR89p8d8WQBDhF2QfDDDtd5+wMAefawZXfwqPwUHdK0nNyustrMTwuv9+CTA1JXy97/uEmckL
LnMAlzGnbUuDziLHLg6l/+OPFKk480YTbwW6fIcr+ITAfAVh+kcEH8xos65ztW5ROuHRncPf61mp
gh3aMaeLdgYmFSfoaR7zJhOKJvvEbjM5VKs/SB1wOjSx/9CvWo4/JqanEEWsWSkZRGsmXT3cXF0z
hIjW7HmSk8VgosRmiyZRjBPoMQSmPU1rVkUpfAFqUWBKp64/QrUdBXVcQtZLu8wFiLMZBZMNko8o
aDhAz6u59/+ETdHRWY5NPWJQ7TSqMDm+72Nd9gau1O22te796pmX3btAwFokbnrgyb2AmCE4N/s8
PsPLuBCLU+C7PoGZ5QRwSehF1F1OZh5FA29DS2OmtaXn8YCXMBeu4IoMNLJ+hm0gHxjcrBCG3oqp
03DOqo7YPSdXXmfaKb2DWyfNxwCKJyrF6qm2XKm4ORwpHbJPWZ0I0sLUUnAQCIubTbFoq9GZGdmc
8uoh+hghOMQrilP1n51EPk32ygSNLpA4EzycaTXVJrkTJ2R7oMkqObJYPcdfDQ4VOoXR6tTBQVIg
UoQPGeT/RRAYI/Db4nXVtPChWEvMWfouZK6puWOlHV00Z5Yq1x1UH7XulYAkC2rhwzCiMwRJw8GX
WBJR7pR1YupX8MYlOgrf2cbvp2Wjz+9+K//VxMcnSn2wHg0MfVNBWAIpt0cWf1Zb96uhj+UcefRB
efIqDG4SgAIRzmx3Ycv5a+YfZ1mu5cyZTr6ssxQ0/PrDH+keOEuM4A51R9jcLa143Lv3ivBQmYVt
IJNYWWqQD8cnlib89Nr9tjMPCNPxL5/ryKXPLYqG+4rEm0nprWbVb9E+wFgLT1VmI25iyL/UZ4Wf
62uc/ctRyXYpLcpcb7zmrYdXrcNroY9mnWFgM9a9/33LFCPPTPDAz3cLx8N4PxnQQChk0kN+7Nk7
IMoXLu68sVFz+emoDYM2gEPO1qToYcrhTmaS8KeyD6Hr8LAaeTOeYmzPsbPn+AuEYIPO/635fvIw
T/jWIbNGk22vVgz8MuEDdpNunC0JtX8JVb0GQ5LoWa9b7RG5ZX6COt7tUb04QHhAJ4hIIKcTfrRS
lexcs2z0Jw+ttS1lNjCv5BBNJQa0v26aA9Rvbznr2o++Wn2+4dvdXk2EUKconSmgbwcDNL+hF/sh
UgZ0Pbj/7FjgxMbPtICmHFrbaRtoRJAtdYkLFtOquZ1G7uvq+C0eCYy+19etrWe7iTrPnjCEfclJ
rvI0isAqzhBx2GeRS+B+z7j+FEy35efurbFdI5r0sodGtOgcihocuEQvPUe2vsBx7Fg4PWvvQxlT
TuU5dtXrC+t+/qJbZuFaZEEbdKjYoLqNLcv5ZISs4VPSg5K9e5l6ia4h7rQcaT3l0/RUlPu5bmB9
pd/9ucWRLKJmLHHNkNx6pxzRc7bXqHIRmNY2Or1kqnnOfsAaO1L6qNI9Kf7dN6bXZ08uJ+ohHH0f
LYSe7kKKWI5ASmAlIQxaUx+QXzCoMat8tJL5fdPWE6DSIM/uCcyGNn1a4xfDUaxq166E1GCwX0mi
qk4tZAKAYVdBodk586GaZZhr8mStpc1RgvUI+SlXx4/5VUcAykAN1ZfzEZ0+wZIkwrmmSNV4N5TF
AICa09ltdkEsIlFIcDqLUnLZYFLSX4WgZOJE5WjFyWQZFuPOIbiG0m6xhRgbPTqndvmNdC1shbB0
rPUiZBwrpg3TvNWf7pZQanaeCm1U6b6sLMfTb3C359mrPtzqLHaJiHv9+j0u9fLW2xk19MhsEcH4
tBckPDbhhH6eHy8ywTTCdWYj5t7JQGeFRo6C1+Vlk4K1/9JSq8Wb5nT0FWTEeI2cIE2WfoITOMni
9CGNW9Z9bko/IY5yC3/ZRzCgI2XtrrgpexCuRNt2dUlO+i5OipGj+KeYs917JkVfstJnIFy1SiuB
AyjKpD4o7eEYHCodcdwIYO/HgIwCBWDYvQnYwZlGBq6BU1ITupRIN1C2Pwo2fKYx4633tEHtv01c
M87z+Th6jBLjmj/rg+vOw6WZ52fsrN8oNBrWhF3AZ4L/diYQtiS/TONVkU4wRv/ZCDWO659+fhLZ
jQhHhrbteAdSA3VuDI7BkVzkNKaqD3mjovf9qdCt4ULsdYjmMLDOh63rdhLTF/f9LwCFobA/x3vM
xEN4To03lUrpuD/ooqVjR3sumpl5hHtJZLVaeYz1OBMbl/l3Naoy/lCpSycpyPgHlIxzX5Zw7Afe
btwRVlseL7V2DY/+hB/cRKsiSBDV4mW/lg0b0SzWwfWt7RrdKUvUFst4lcJDeaD6fMssPg/WduWB
6I58ZLxCeYo3Wg3qhQzqDc3vMmElzL8unq+gxJp9p0lnZtn5IptGNae7dOpvBs9f2i3Zd9kPQoki
AitZHP1ldXm803PT+WmjwbRzs9ncDeTHGslXDWwbQSYRo6f5ia+rX5s9Jnki569k+SByvgDKp/vj
zmyPzDv7pLo4rUu8zEEkAINvWnGfQ9wH++qxPVhUYMBp1DOf3xXLUPudV6ZQj2Z2SkMB6XJoyrQD
77vsKqgKOcqfXw/7OIiuJ9d4m1Izrq77biKlssDjM/0SY3J6TGOofPlkOaeGkL6jocpMQVa7S+Jh
U0ypv27qYpAzogpcWMVeiIlaLhF+yTef3cX1FbjyO+zHXho/BaxYVDBxwHW6xfPYDV7oi7Kw1Gkc
iGix/d2lFbixADG0ZxDAkQBYmEUDbng6OSL14fgSlYRxkU4TyhyFVMfGWGJGOpgGdnTDliB7chZ6
RxZrX6wGlrK5wWhnKRrqji2L6OAyJL/jlkCjO/bdI8JQiKtfoMmeEW8brtRdUqDU1lyntm7HxjkA
3UPk/ONHa0YhdNdIvAP6JXt15rRYaOQpnE5c5temRjgt8oKaPCA4z7rdiW4XxYoC/+m22hbinQvK
vK2xNhMHnsbkmUtZ7C2OiHYabRbxh7ZAN80TiMKFNdl25OnD4kKtAX5+DgU/ALROJ94BcvAtaboR
m0Rg3TNtlAlegY1e/U+2FZfvmKwm3+VOfs6vRBRCYVXU78ZHZ3iyF2KDjZ8CE0QN4KiAuN990i4c
zITM/cjMEHVdos4jGyQWlhAGkC7xZFwFe9upHxL9+CKsHb3PUAI4/7feMZBWRIPQ5563Sg5staIi
8D9qihkSp8ZvhbfVt1AC2lc0JXDwe5I/OpfA7AjOCji7T5XajbQ0dl2SWDwVRKifoeHjCrDGBgBP
i9wiws0V2OP0e9E/zTUaI/PTZ5sveJ1KiJO9t+nI5tJ7+6udhLHTEhfq096MGA9tIbJHDXzu+ga/
wPEdzyP4RBa+Bv2SE//zx+cMGXAYzNZ3wZZ+AwW09kvPLnAKxgrOUdou+quzy9IyvPopvKR6DalW
ryYYLhOjibb5GN2mKf5Iq3mWAIEWDUbqoW8RPD73jjOUbGrF7a9uCj9nY4b07xBgzZ9Aa8wTkBOg
UUm8/7E/IRCB84udTkZnlYSpwoINGmX2AIHUFqSxm3g4G2d9vbS9T8hKevfrxlkR5G9/36cxQxXx
j8ulCpNqqX6JfIC39HQijr7/cWyzlVrqwYhguBI0A/tOdohFb2VznJUSrfN4PG+SaiII1T5Utzo5
VVMtM4vLbl/JrYDckfKKWIMw8WEYQuC4//0OP4ju3pEad0KEK7XdKR58xjlAgw+WdpRn6BnwwiBR
19wjiDI+lNfdzDeSAYUw4ZP4FyEW+U42JrfNMlRdT9KVqumZlyRTEGgs2xMkU67W8EmsgnLKN1Yh
nYh9w5FYFKXwA2H0TVEx5EHPstCRUSrUuqJB7hvsnWCSMQ7CqplyO22avO+6iMRJCliZ/89CGytq
qlqrL7kri+nCiY0YEkdOyMWTm1OYdu/XlrkW1p4KaeyvRj0gT0VvnvkfOgII8TRsP8i4/YCAwnHR
brifimFmyP6wuaCAUnV7uxOrG5MyrNYI50JXaWXyI7k03hXmUcuft3R//yP3MRtrqaNx1zKU9Oe8
Rwow03T8xIUqMbOqOUj3AdjH17UyF5O1UAg4vtOPu3gtz2XzBabFhT+7WzQ6XmCpRu+oBKyhP4PA
2gddkRtAKD12PaILC721HYnZVwFcOW+HK0eGMpuxeOaRiQpUxaLJRdBqsOfdEcRMMQ7tfueRbCk0
TFQFmjkxzwJM4WrFvml4RO6slEkq8MoOZpNxsIboFnS6MR82V1lXT4He/x6GIrjWvtW2R0jcwSrY
/EmLuZzToMg0fnz/QR9eou/5tCLZ5eHo2EwWrniz/j4tKoY2cMzOFS/hvCctMAJiA0A2XoWv6DRr
aLz0TS5mt+/20Jw6uLMBNyV18J20awTvCnrPCQWNs926XjTZSxGAyMO3H4wqGbfYEmoKNl+InoFN
yT0DUJ4jzqTW9uRsu5j4InB3eYgGtZiMOejflGNAwmCr9NtQHhBOOMOezBgo5/7izBnDE+6oT5Tg
5GQEA/gaA4hxks9lguL5pRHGP22wVjAYYpQvD+/G/+Ha/BrIG8DqrtscurvEAlAw2zV7kgRP7Jvu
d7lqNUSTzf6aWtpjszMK/G1DTVWoHanac9lINb40QqQjv1lrNA09PayiRJ+iqGdU4sVWq0xSZMoB
51gls+TcbcyWo0wE2APkE0IcIV96atgDFnbRyNq+VqJiUnF7NP7ueP7eZ50pI6mxZEb6uBK/TusT
vOxiEKC5xWYvb922GNbV213srPjDb8YnmA83whRKxEg5zwVrzkHoYoNo9MyZKUbxbgD6jSWnhSWZ
TmBlyP8KIVVDMkJfHrTTVZt02YrGWBjep+lhjOtyfLdCq/tvURhdfCd5gMn4rec4Bva/0vRinVfO
M2K8k7CL0j90ePqUqkA2kEgTNOxD9kTn7J5f9TzEOkgWX1bLlC0L46xibDztRyLxCWiy8XDlOMQd
SF3247kR9cM54hFIng6AP+T4E09tYW6ROyh31rvxQ2Vy0L9v+8Uwk72dCTjfUfn4A2pbWKflxwG6
7uai6IxIGCg+loWOua/JAU3lreVPL1m0ql9fqloLvMXqtWOLUV5NXaDjuaNXcgDaDN1KN+nlZA0V
kyVBgYG3gEFjFv3SH0fLaY0cKcIui52bcj1cu1DHWyLZ7HCK8gEeB7wct4sOn4C/4AentNhppLRN
qKErF7HPwDM701k+tTDGPsdw2vtf3BnxemdW67WOjyOFDYnT3RUk7logHUMh0frpgM96YoMFBgS7
RAxVYpS40CvFh1p8alAM8n3dLOxrYaC91/KLi6wqZrK5fSOj+FLFajKlZWWytXxME6q8SzVqPAm0
62Y+BzaC/E65MCPKpH0N7S4Hizubzf+5nAjq7LQlpEv2AMco7a2XFG2A9CXpxk4EjuxfVnuCWodH
kDBUrlFaXX1lAwC1RiwF/ySNKUaZNB4TMFY2ndx5RaowXYh20gZxXeOW9Zbw6WUC5pyC6vyU7na5
+oZYvr7SM9Vw5VctWUFqEGnckyMMVJzutNtMw1QO97HGJllhwJCGjKDHtFOiRGeK8k7FsEDNlCI/
wDBfxExtXaGbh9XdVyJmli9p7rkEMJwcxAERoBl9u0LwXeOzEnedIoyJyxMX2vhmYDTfAdeWab2+
LW57G+HvvfJKvAvEzxCe9czxHaafeB88MLq8qoGN0MAulmBcNGcBzEq9xUdMa3CkSavTEFUduPxg
knTA0ETnGztoCRG+TCvFehCDvLl6M4zDhA4nNftV6aRypXSbNqi+kBRg8INVdOihxH1Lg8Pz81HB
Nn3oSO6kXTBuxm8T3+W0fZOKy0zPcHW5ktcrOeG3VovMjlHN4t+SDbTxiyHdRG5AVtkHtC9Smjok
vLkDyYxgxKA/csg2B2FlIdTd8eN2Hxs89hnZGNRjIzMe2JxOLFXKh3N+UcaOX4i+qcTnKuXkXHvL
HN2Z+Wzp3FVUpV5W6TwVwJUfjvovGGg7mSw8z47lWZHUsQPxAbcNhlIXAfQcNQN9Pg+n29kRWpFx
U+ZozPxz4ZwW2bPtZ/mF1EblOcAt//+HX51ETRAJ5ofIJXNYOvD24E1u02fJDmmQ348ePd3Suxf2
MxGusSULu7JHHaFs0KRsRyx5Tzl4f97lI7LhbmAdRNtnuTp7XbTmvPEskSdY9RfHw52P2u0ifV3S
FNAiQY/ezOSqcHP/7NbmfBmmJihdQ5zM+mfyYKZwgAYi8jU80lTv1DEfL2TkPH8vCakwOusvSP+i
nK1afzdA82zXXkXQW1SkMpwyGiRiP4OlfvXtfC+NjqRFTeVh2leJfwywzsTQk7ogvv4X68VXVoa1
gb+FVdecQBN6Z+4pSCrhR3Rqq0O+6Km9q0mv+UfljeW/vr3/0Hz1dUFWyZ2TOMAN+5ja5DPJ0yZT
A4jeIhuO1modbFdEGvakorxebA7jHAJYpWjfbJ4uob8txrio3+/u2vlbJQKzfrRArnbRwEweTH1H
IVy33dSiaE8HOlea9Yi7mzzLJWoVXPqgWYrui/mkOBZg/OZDS2EkDJEXaJw8sLDs9R/i+zw66hd8
ZKagG860k2SiNZqm4VNKHLBm/8a8B7EP5Dsc0MHlIf8lmxjlgKmu0xLJo+clG3YWqJVVzRK+epBE
hwzdPmYUyFMI775PIxgZX2ZSwNTAURy3XQYX5gplqedvxpymSJ9s/lXObYcNem6cOFvuG7rcfteq
iuWaBSu07ELxXJfPpNOEkyvAAJa7EDjD4THq30eHKqI3JA/h+xDxlh3hv/850DrqwTswwvcKAOTp
2l/bpYtc5SB79kjoAD6Q/BnxxXKd84q2kTAMOS7LNWgeGpfNZchpzpBc5EIwoRdoFHz5W0hOf/OV
QFXeM645pqpBwFWLh1MnCnXa/ADCzaxP9o0jCbQvDVkUFSDxPnnOrL+w3o20P9oYUmHPwxz7yknr
8RBeZJB71Nx7uK79XxdLceMwEZVR5wBqfeCEEJFXI8DMpxPxZXub8Qbxk1vcVC8oM1G6vAiCbRbr
n0xpmALBGVGcUpsBsk5njwN3s/sd5b179X1kUJgWG9rsqzma2M9XhBUO694VF9rgnjHYTCmD1AUw
Dg0MfK9O4tgpC6dBfhgK+6dKiMDSxoP1mvZ42X7VNKniVvuIDRiM37K9enQcjWbedwQ18h1X75z/
axMZJWeAVIvLqRwpTOmay4+JdAzS5Olsazzlk5cN7uJ2I38c/WIRZ74xtvT6AZg4+tgxzY3ncTiI
qOGJjUo2BsSpWr/L53sbqYSHFMVAZDPiJ6BvgZgV3P3weyhhS5U+BLriNLa2t7sk7IPwXLH+s8wh
iBO9qnfOXq5Sp0n2jSaeSZHEIovSh+9g7ClrzsWAVqLuvNlkmAzZcIEq5Hey7wenQmQWeTadPhkP
2MA2K8YoSRn7i7ifW5cfLlXsvEKW/Lf8J/f1WLa4rNkLNTQPsr/vCsdFMYOIVHEkywSaGw4jEp5i
yXoMDeBRZXZIZy+Yfs29dCyBFC6onzK4oB49pwF+fnIalic9J91Wihy0JmdEDFvwhyJx9uzJFNsk
JxSFKfvtZQ75TWhJqiQbYGyKLjMV1R/39lM9hwzvr9f00lo5tGalQisaxcWs0LBvORuGbJ1HUw3D
wqXzT+j1KomwHMf+8YAYQljjgt/ExK2PF+heWJYTZwbpZf0HrSqNoN4bei2QKsxyt6LUsEpxCyY3
wDZGzSzgRpj663Nzntmhu8X8bxbdie3aTirWznYUM8Sw5nrLJh0/9pJYnuh200tETEhmljncJjOW
1FgtHmFCRrNVCj7J78LwZxHeORLQOqyw6kx6+RO9zsPCdwyLLvV1EfV3g4tYu3Q6s6re8x4k5L+C
qQq3YCnv8kfWLSgvO9XfZB6PXZI0CFIJPR9d9e8I9uujuM4r9aobQyPnCiiIjFt0SXLu4NSzWVBi
TsGI9a+kBCPGswvrMJFvpdWcB5IUIUUyXu/VyErvswpoGryAijK72pJlzea5SGx2aFH0VdWH9hOv
+nuLfFOt4LtOAgM07Lu9heUEi4E426iNUGraKQ32UEwpkObfPXCXW5zPRBHqAkLOV6xP/JFqeHGm
foaUxjAdUpBKO+eB5EkK/G3MhRMNAI9nKvxTf7wV0/HxyZapJNy7Ex6eNVJY5tsYSue01TzZCMJ/
o9xQXq/tuCsvA3ADwqWXDOQWlllpczAhAQA/MNxiwN8vYfLR1i26MoMJkVMGn6BNrq/g2v7f68m8
oTCCS9ZjMY+PBFPlrjteQxkX1ggVltVy9sV5dEON0Mv2pBjdrnnXuWtmhPXyWeLOVR7wYr5HP8i9
uWSHD12ARYda/ccKPrAXBm8KGn62GeRIblptlELcQ2WNeqlvANBQA55pTO4/liKBpZkzdvyxXmal
VbOj9zQ9FszQsV0qA93219jHaFkQ/16dnvlL90K5TkMnSZ/WY455z/UkwTfh7Pkr0PIWwYjIHsNg
NCuz/RpJifqdeSiOCnoqZhQYSTSBKVviKAFSq6Z3U8jAHieZoo5FduwHsn67DaY3wHkj3bCVkMON
ZB2Iym9ONZjy0tQJwhQlfM84bAuecdEVc+GYhIpaGoNrmkKBbCXa9rhe7ZntChiUpRFUgqOkHZ1w
akvmpS/qQb5Jk1Y7BnQYki4FnnRsWEzAY6yeAFncyFQepDq/4fD3ksgHappEV0pbnLQdDtJa0x4w
pzHDvbWuz2y6L8LmPYr/vZV7nsMsAiVFhOBFiiO2PFr+r+4x67epHc63oj/LCduyva+pashgfxPN
zSEdJYDyYiVgZE1keUIADSi71M3suhwxAcJ5UxptGEQKEVPaLk+FvHo8F8jFTwLHNNaG1Wv7bD+r
k8sd+TN3po0i5dyQ0h/G1cQ/yE3ChcquC8XsCwH+BMu0FgrEuAxdChlDuYtyPPJ6SUKc7HOeVy+n
PN63T0OVwHK19m9ytZXLZWM4EQiSQLt7tUmOQYsPd7YB5wTEMPp8sTQDfY2qzCjhNPd5qyWpxaF5
/1SdCoZH03A70Tl0KTKc4hinJz9ELqxlkaBHJW+7lZ2DQWm0qGN+rx6lZEbypJRlDYf0YZri+tlk
574b2oTtDgoYLAdWjHs5KYkG9Yk9+GpH+46gfhyJGSkWdgstKu01cnmRovxe3O/cNybMtetbtp82
YJ9SfK6aIL9mYpeCAmuO88RfRCdxGf9crcpFqstAQ4EVo+KJJZKtaZufXmJ6suhdlAQzkk+cOmZL
Jq0Jy1ljtWY603CMSPx9A+LikF2StBLdflt2as2FtgQzgWHEvwTVAF2XLFJYz40HHgXSVnK1FWtz
1u+KwuIFvZubOzP2dAh6zrDPIS7KVEGQELa5jvqJM+GDAzK0Bia3fYQsviAymG3yWhwZOHv8xCht
dPVB2d6pdgbRpHvMZU7SSktOPZg1rvR24HH4Bo4jBhEzhb8hUf86ayCy/Nmi43ktc/rJO74iEoPY
a2OsWpOaHNL02L9xwTES+1CvCRs+r2676kYU7JNAiNRY+1fYD4/lJi9YqUagjWP2VOvMqxUa0R87
yuX5/RAP4m/bGIowSlutGGzUfK8q4itUXdDl+ufYBmbVWsPbKo8dmkEAexGZiV3HGqOeH8+8N1Ep
627DxoIfALvrHpK1yu5yiFoGq0RHqcCXNLZ4vzPgGxGkJhZWOuGiEE9sl18h6Bu2CJ9CZPyM7Ste
Uo74NB/1HzFuWj/7JPLj11MeFVYSHjhp0zRFbl3GkT71McG3Sw+hs3LPsQxN4P4JnxFIM/Z6D3lH
tzGueGmpYZ+2RFJ/eJfQinzVWIs7oPAT/b1Bat6N86eUj9LgiuUsrcyXGA8Tk6YtJ4MVpIsTV8xZ
hCRfvXqq1k1txb9ytf9FtTGUIkXIeILc9FN5Q8L81AbmnPJV/G6bxn1kO6nNDFCJvGFkORpD9mRx
fFuKRpZhulrS+W+XUAOvJxZYwg2FjDvHi8/2GWh0z1gyyK2mFbS7Qe0dZTJ7Ckoiq6AayarvQsPk
bNtZqolNZ7RbM1DPnyccdgiWY3+nmv/BmVB1Ev79h8yk+kEIzk1/lRbFmiNJPPROChy8Wk009JBz
F/DojLaQEDRPaKmos62WeqwxErDkasTfn465EzQfpxB4hJIPzJRHrhkQaucB/T2S291kVhqeeNxr
wxRwp+N2LQIy5mQjiXRZbHsi8JF3+rgSplj3bd0hVFDdhu9NtpcQWYpJIFtV17UKTa0tlGVEQp89
j/RAs7cl2r58E4j8zrBH5NWDHm+wrSW3R3KjOEpQu3wBfmUjK15XZKsIlLr98udZRusm5qwJYmw+
I4LxqfICN+swqMrscmzYvuZeoAJSav0aY+dGkDBV0EJkCSGFei4oANrB1zKQXGoia45lGa6nzMdK
PjyTOFklopYolzbjEM6goOBPmSyOHfFC4kDbbMm/MVyytEtg+dcUfSPJu7dScnHesxja2tuPhhH4
Rb1icAgkG+zn7EnuYvWXK4f7m57SBzSr+CY5fpbTZ5Kfr8k6Kc/JKwKp5zKb7VwfJYIIRjzrt4jZ
t0HT2G8E2tldsYhCJPxvGwTxne6nyukHXNbLA3ut+2x+TFpzU+Sbmdg2KC2BZkMSxPjL6QLQLLXi
Q2yH+GQkyS9Q6p3/0dInU7by4jY4LIOvBFqiPtOBZ/zdyjyw3lFe7hnj9PNE/0LbLIO+/OgevfeM
IRbuP7hNxRz4ep7PS6Q1CIY62ptWwNBuAmhbaVuld8k9J+0+68/QSKo83pGEe47Cmz+H2hsdqZ2R
4ITkENB5VrnxPZTgl5hCRitx67Jxe185e1Pv4zASIj74qmwKHp4PJrjQo6MECWrP9L8IL8L1iOtR
6SbvjAaA2MS8FRddjMVhmJqoFtHk8zpQMxmrCn8ZYi5eB8OkcEY8/G15AVBbs0iVBXoOxe6hL/KC
zQVh7fAL186ex/YyFOaMOCzdV/HiZ2xm82926v38ioKjFZwMMbv26+k8T0D7dZLBPBlrVUy3MdlJ
5JEXUfDEWDT30oHaRjIX5aWF48+lR8pz7Cjrd2T5tbdOc8XiwMC8kCD4LXrXdGNsAD1WZ7V51was
A6HMhCLQ4JmJpdWfk/xyCODZXg7LpQTp1p0a2FDnsWyfcfE4GIeOnyuIY6zleeEagO6mhsci0BB3
fRYbxpiA1gM53iPXZex958qkaTM66tc9pSTrRBaBq+JRmVk5HOte1vHL8AbQ++WlULfZsMl4UXNY
rlwUAwIGxOVPK/rkRmhlQ0mKUQHAW/iGqgesD6K+4Jf3EPugF8OuAq5sj9m0wuf07YrLX8jnu6JY
j7DAnZblVZf3MUFOfsduyScB6o7KSkJfUDN6oM8gNnQjz+wK/l7lVWyL4XEGjSATzyS/gX1K6pj2
hdDWkNq5CK6US+HL1RKlJ7VK8u0zTR8TnxVXz7hVw1xg+Mw6vSmWXL/je80tG7yhnb0bwNRORmcP
dsyUBs9x9LVoYGikaBkFYSBOyHm6AC7w+kIDlF7pitTW/20vijChUyoi/iywxTOXZduSkIDZWqlI
0QX0axrVDneHpoWu7q74xuMzDcoQa0vL2kU25btEyV7IE372lsYG4jnyyRRNy+pzy+vrZ+Yv48Je
QIWvHlILlRtEUBD3oEUVOmh0mKyqLhtXtdp6tI4x3LxnN9fD+TgXvKMaATIUD6qh31q4a1kjK1/9
cJ0C9D9jtKJuGlCE8yoaHR+nhETMBXoJW96cia8PNPRqFgmhDQGgaL/JuOosBc8UCkqaPhEdxzPo
t8t4Ag8tLC8qyTllIpguyQsEOl/FrfG8SqfaHvuff/xtRBwKRPB3sSN9squU/rHShpNQ6dhwvW3F
cU+iKJUCpu4sCSIKpCPESXDsVQe1RMjzwUU4n7OjAafeRmMzYXZ62rUYDuzKv2PvrSjR46gZwMwk
3ce86xDoSFZmz+/uD6smXS/IKJsyf7ylAJM8HK3z3zX1Zv5US9rc3J4FouVjSSJPpvUCKjG9nNg2
iTxFRE9lHO7rbWh1R6FuKIsKK5igVfrZOXPPwxwurHyXOgwUPANlpsP/AjgVNJlcfbVJ8qOnU9pG
ZnUfBS2Nq+ESrI2qP5XlucWlZXiZpSr8zbSpYQycrDGVdHoQmgHrjo2uelkmwWE2Gkm90RENyqKm
XUBlrrNzcxJ5Le2mOu7/r6ELylAAVIpInHAy9/FIQ2WD+9xzotIfFhNWiKrIMGn0ieWQv/WMCSen
KQWtgUmE2TG64ioiW147Iu9Is1HVA+abnnAxJh4oxc374yrnlor5xmxLwxm90XSoGVBJ6DJmH/xW
7invfjjiErJ0sXswcAS76YbB0QXJJrNxVX9lFiLw/MefrmCMpBr2oylFW1wGebWYIaFXQU2XGYVn
7AymgJ/Nx7I0aORGzL/8+sQXPqB81fsYY0wRZoqT6/qRkL7S3622DV+H0vE2JBPt2o0CnsKYMu2A
GVb4kYeoQiCxMor/g8C23pH3WIA/Mo1M7+lctZQiAjvmiNhrDVwouW+b0AnMZ0BZKOwY8C7j77tl
H/ydj/BP63uZ7rnUEqktOSw22T9syei7l97D2LyG4+yxV6OuiEvnYI/w5sepqJvwnS1giN43yf6s
k4j5Azql5coIcO07PSp6Welsts4/weChZ89WHwWlpqfbOk7oGOELtkxKXnWnGOxgRGkb84qcQ/Wz
zFtRe+TWTnsy76hwnw42F40+j8oT/oBv3TC0WzNh2Y8Eb58sEqrYL2AexS+kmI3froVhKWTXasyw
XZNxKLmXDwqpXJ85mycAPKvPXV+Baof0FHW98rYCTNmrd1/ZKWNFU3/2FGE0aGH2QU5qptWHsGIU
0GlhJ9WRwRwPmHM/VSPAoasUuW4q6mpTbYtIR6timW2xWzifkWjSCPt//tugfoOGjLHgJ7K3PjHP
5zCFIZkYHL3qkTgHOxp3vKx6QHsUeFqIUx2reiMSXZCXWCMh44GLv+LHRqY8+HPXoZkdReiNkmpD
+Wee6RXs2gvb/Fd/d5eixVCIj8N9reHiEBihLfxZUFunv3BHBvZJLWPkx12h1sJm6JzsSWN3lbe8
mLPxuJEye7Cr0rODwgTWChy6uy8z1HhysKpR8EJLYuVi+ZPu2ziy/vw2I8odJtk2dxLolKXnhqqx
6qkF9zrgkq84uL5yusErVrKU9RtqkCjKenUjMC2NBlrlZaR9gVhmgTMTwByCcBa5KUU2fwIdfJUW
JffqED73fWbJdUjs/Ud3w0Pqvz6dxFAV/G6ePMVPqRmy0iqcIu+jPeE3ffMYqr6bmpvE6JdPzmE+
uYNtq2RVaD/4R3dcgoTe/9NlhMZ6FFXbo06b3sx9CbjHDsR4v+R5ln+eDouvWUzmvR6altMgud3d
Gkd4QWhV8+i5oyYKylDigFLjPqgqUiJWzfdkraR61K4d+3T2Dpshb9D0O4LKkzo4R5ZAt1AYAnqd
a5Yl34Sb1cqsYF+y4fZ6FOn67ICqPijEAalGY8ZZny+XyJTBLWncUhV6ATOf172eKVLKDhRpjjcm
la6igW1wbotNq+dxuecppjWFAo6/wrNZX3oNlQJaafOvG2uV6IdPNGGuLCIO9cjNutxPq2vMoZL8
2ZhPsC3fPlo2E5fqYaJ44z5F+HHj1LRu6kJlL2IBIOlB/VZlHdTtUMabwFCPAa6AGKVhmnYtszoM
Aam3i+A33NxZK66jk+kYmFryKnQ1UCRzNF4vApy7LAJJy79UNodXUz2uiXT/HKucJRIoPq1sK8NB
NraihtKcUkJFQGTIdXeQ7GctHerY3TUyCIKS2RPJdmQkrLExY42tdARAyceirFvPD5eggQvpDw1y
3gfim+EbCKWjn3eKzBzsvcfzEQNwnph8xd5lv9RUMAQZroMssyAtjs3PIZ0NZfMVYuwwdpfXTZlu
3FDv0ZS5ywEDl+iWuO84wSv7MA7X7ny5hbcpjEU9BRhqhReuHYyYwnkhMz50WrYH7O9CtP4/1pdU
2nnOyMOc4IqCWIUGAWsBVEO8zF/4ShnwzzWpLLvirUNyqyReF96BP9dmwx/SRWG7lzU1DNwWwo0v
DqoFdC+aDh7JfJlQ1vioX56OtCG8hynoOZ/I6bD+bSYDat9QkLnGkodDs0ltlLmM/kOFoYdK1VXe
6Bea9WFAARZzjsec7nzQIOQEvzaCiApHyA2r6mnmWgsVRIF2Z2iR2G0lcheh7zn6/QoYZURDNlCA
2z8eGOGfh7OMZ/nEIjMnyAHuArG82jJPduQQeOei+T3iq+0PKq5/7ai/qhcJfvvrt+8ZHwxokly5
g5p+juEWm9YZ1R+58qdj4rAZGZEEm/B8PiBkCG0Cd0OYbz2kUd8NLkj9hK8pLMVuXHYGvj2/DBCO
i0X0gXQMCFL4SA7cfg0mnakA0xEPXnIrrp0LnXlPCFIopb2B69HInx9QNHRES4Yp0uz0fXrZUQFW
7NVm+nRHvXaK5BzjkG6B+FT4i8JWwzsrALJCj0Sv+DY8KPP4UKMSwxIWlaS0OBkj9apCJXGEZEwB
27Ij/2+mzfiCYrE8uXhM86ml3AMnA5pga8euZQGBOTGJbs+ZwjZqNZLPeip4OtKFkutsxbKjf+16
qH7T9+z3BuA+saV/ZeZCuw+TfsrOk45RmJgvSz+CFwbU3HDSYK603ZXOFLeD1+SZQGr6ug5AbCnF
vqq/xz7yerJKBMB/zSQbjL3AFGy+QSczI974I2CB1XehpKQO0+gJHx0eZLtxsqSH1sIYNniVG0Mp
dcY057ON/oMcU7Ll+lFCbiL3gBKyfKdBQ1gGqnN5MUUeoU5TwtWsMFjQoFuebaWeTA99aAsKaR3P
6Wf/OFvxh1fcRAgbUf/byefYMY+JUVhIasU5sDWhSdLa0emjs8siV6tMqDqv75JaLL23Iioug43J
a9S/ovLH1O+TYHO9Y4CfJ5A8OtYm4qQrOh9zEWQYOBpcTBTKnWCpgK5lReoHXABIfYU2sDDe48UQ
6Hh/qNyxVhEqm7ur+YVgUGAUf/GT+v/ZQkfvD5vBpjfBGC1tyTszUgnWxyTqpCcpOvbKY8EOsloD
x8l01pR59gckhbi3PI81QqHYORNoG+Em5tXOGLiG/Sznd999nudcT0vCcm4XwY4kpfjAUAEGOhRT
tg9LD6MfHwnSbxJq7a7ORmCWGxBg1rv78NuA49NibXuLCTiZxgmNj5O8Xs5FbVmMjzPH73o5WFzs
lZGK+VZpVyz4i74N92SvwnU1k5mrdbmmVPvjOMufVz0FXv+hahKO25SyGjfM06pwoRh0XwsVybrI
baxVvkeShFvCU6ab6HQbINKOSc8Ddkj/YnbGjdbBAkjJGYUtTy5RMQlzt2LEOI561p5GcOlpU+po
SoSMiSKgq4rvOTAQzgzOg663lm/nD8vLFsO/dWonjCHvDqX4KU7AOP+uyJckysPvH9fNa7cIxi02
5LPS/kX4jjCCDb0zKEBBqyCVbQfZlokH+k12V/L8PfhfiDHOjykfnVqU0pNI8m8PA6q0eXHtYfuu
qzzd/Js1ZZN4VcHFcq6thXxexYOYVCr6LKY0DIGJOpYo2ixcrEFauIcglAafbTFcj96W+ZOQChFU
RwEwF8Zf0Y+xGXejF1EQQj5OpvS5r3ZdO4KNsFE3ZRMwEKVs717E7x5le7HCeLTwGVUP7IjpjeKS
q//wNlYDUIdVOSLVA8li6Oc9hZ3hge3halU+Kt69Dw/YtfUbgPt3do2JMwm1cknMXBHKTop/D/5+
UMJtZpPoz0ejBlJLzxhpYerGaVq2xH8wfr4nyAe/GlOMhYXR3H5C/iJx7CQI++lqvTx22hJ3EVcO
6OMqQXvul4J7BkJZm35zU2MxrF5hhkBKjESaIiZu9/CgKnylAyI/vAKS2R09hy5QXjAllLZU5iwC
sPHYCAVDFsipGclhDi91R5Y35cirJinbEP4VJlwH3eHQBLrwOLogqVQ3LrbxJFYZVfVEr/c8qt/a
DiGk6irIHOkAfagUOmsjCZDbnATxLnoxjJKQGzo2+9+SYTrn2NkvqnYb975zMLgNqb1qPqZNsjR8
hDp5yJMbZiunAVu0m0iFA+rbeQIxQDGuO9eZqwvgpzQpIhjkfJ5k599oaIhHXAYANFSTM9bweRih
VjOIEybtQ8WeY8mdi3L9Y3Tj0pT4E0spwzQV8nBAvuymU2NNJfgj2xgVvjIOSMs1S5ZF2wYpF2sQ
S5Yaz56lh9yezJ8RDOM87r/anc2DtDq78OtXvkFE+hZcw6tcdMziQQzLs6ED3LfLC8k9oO1gkKUU
/HUKBHEd8a4X9we3zutSaBUx7nvVQOfvkIdun2m0jrF1rQ3nEQhKKLnnpl+kZc6f8NTOfEnpMf5w
zDjNmI88kOlddfGFdgFzErZxOGMtq+UFr0uiUkLzXS/KRk8E63n80DBtvcR3vEoebv7Nr+JEdnhM
D8YOcGdniEdjTSDuw9YKxNR6dEM758VL5fqAnGLswO3Jvg8XxlKCTct9v5UYDbgyb1+7hbk88atz
r4bZiYQFMbKyta4eMZxtvvaE0ExtTWCc/jtu+91aLvpo2OYa+BvHqE3QUyj2NhzCJHEDY9Ctz6yj
lCzGv/J1MTI0/V/fqeEZ9wNjxPcPkZntAE90mXP9IWXOMmIQYQlCL3I3cKRnJhLMat+f89XbfmHp
uZ3DN80zOSOFpNEyT3dzB2irO0rLTi28Ct5ZVPnlxuNaHDhVH3SRjTrHYCZbJwbpEepYqzkwAVdD
XAYsB2ESGzznx2UlJYa9BOtkiFVGqwoghof+xpDhqsdmCcKZwwuM1SKXQx5480i4Rn40mKVwKhlb
APyy95Kx0ADbWWMbOtY4B2xr+o8JExdLQS6bvlocsk5SKoF6mhgFIh8xhgq3xK6za7kznSkMWWRx
NrL1btCIBB3avUVFX9VHUcqodPipjBGruuniKl7EHVJgZkB197mgWohZQM2Kaqmg+nq3d7cPZl1c
rMBytu5V5A2VDxcLeiS9sy4LPm1p9WjKTVpg208/KfEPOpwfvUJuY6eEOSRnRJ4hmHCcenbLvMVl
TvlXMLb8W+ISiSbV39IByS+dN5AVQ0My29bTbeNOBhc25ou90LkU3rm41D9UL9nr3jEfxl0Nfqbj
nQiQYcLfWjoaHax/n742aZ1BWBHiXZK/LrRlz/nvj6tdMKDNIsizJbv0tNHnNe/3xs7qvfSw0Y/a
llyKFgTF//BZ6U+Xui0DzHzoYwBA46JLp5N3EM9KBBw5cKfJz0J0SlCqYBbd6LyS4JNZ18vKGA0P
zmp/8mosIJ7yUrpg+hIGiHVihBWm/Quf4SwceSY3gpjeTviL5p4oO2VXkSBoGQW9BFPK6SWFdlAe
cK9RMT842XVxsqykm3rameFHC/CENBvD+OyRsVcdcQ8jp0YXCTAjRJ551b+MLr9XrDG9uMrSm+pf
TX3a1BsCucAmSjbMKR4A9rm+6PWuoJuDbkV1MEdRHP8SDpi6L0mfbcMGyfxdJZIApUqfJNfvHoQE
5qzkt5inZ9BJEuN/AZhLoox3wc2wDKKszfxQNQJx58Y9Ht4ajhHBXYzweIpmsOczWr11h9IiF+Er
lVbF9cABQhvhjFvhMwj/pMXHo0Xv479awX8sABJhaRe+Tq2CyBm1WLz2188dytAmfIdoH8wRI3r7
HduooGMDYTgt0wElyXFyBIs/wVb1Bqw+eflXNAsGcrQBAauZ3DTltRJcLVuZAkp9H73easIP73Y4
3GL1WL+QD6BqCa8ax2JYXoYDtCHVREFK3YduC/WMXlc1VvkyXOBu+fybWZWia7Oukx01n0EY5Bar
EeAVzsUCeB5RZiwI0RemkSpfVwj8UtueGHAWBFBirehE5Nq8WmuhbSmCY8YPfv+nx9TYT58+saei
ndiLhac7oSmElkWwmAO7USJldrJxcEO+DO2cHqNyo1PqxTN1IQlbnJ1eRDIxw5B8bD0U2BdOhFCO
eckOkouEmJx/nGfWXmK3b89TrWUMIo8EJArjhXOoQdU2YYTvuPbCMzfb0lRgSvBgMZBwEWzaakZf
xTsQ0RemXn0WG75TOf9OXoJlwDji0J0C+YqIE3ch6kfFsQpzn6VV8LhaxnSGC+vwCHLfJ4Jr9iDz
Krhd2KoETeFCWGOtr7+iNpS6ZfK7bvvjbklJ6b9k+KiDtSE/KW+yUUNgvc2jpyIUI4jGw5V9iDjf
EpUeB8eXUdHR+SBkg2HoWISsIFqjP98SmcJ59sR+VEy8GRGR/G5tmQRFn0ww7GmFq/xplX19tm6J
fshYVflc/nStk1VAFqq/nxmEzh1edstRd6RbNlepo4wtWqJIVKDlbY6dxqu/YGUbD+pfuv9J7fNp
SmNxu9X3ETjSCQ+R8wOwPBhlwixCrVHs3QSGvm3P075TGt3eBO4HuL7NSzN7wLn3PGQ2PVilPp8d
qQxNtaNVdQYCmmm/paLKMv8eCNryQWV57mMo582ylU3S3x8Nax3Vj9sXiKRqlRFEo1hrnJ8EcKs4
KcMVa+ZDWJEEn6bh7Lr4AF5DrYQNYmMXCcNPKMEam1faRD8ZiUU/ANIYQLSI5Iyhiu5cOUFDmXOv
Cp7OjRhVfP+VOoJDg32wGJ0nd514npbQGguydxLrSlSUBzF9U77q0CWpOqB5Y70abEBx2CXEfn17
zUOExUjq9JISXMd1xbpFgITAF8xm8q7M0icgTNZ6KarEyfM/tECapq46RY6AKrpwXIGbFnMvQ18N
EA9irvCQborBjO8PjcEF5merq/qK1QQAyQ1Tr7dNyJUVQb5Uco7qtGMUoGtOtpJZ8Y2v/bzx2DCf
Q74hBdTTiZ7xtjf0HeyhrRTwwTrdREROSl3SHeNV9D30RTXVxe/Gh0blhM3iXVJ0JoefVNyL3Rs4
/hK062RjQlASDIXiQIk80i3frQkhXPABY5WFkiiyG4x9E48h/YkzIYLoY7g4wCn00iuzZzC193qQ
M8ZKv7+nxfFnJ2eoTvnR0F6fjA4/uYaMME0xFlvtgC0mWA0XhPSQxspO66hFBcwq+5c6gKRMCgs4
eDCfnI4SNMZNqHZe/5ii+8ZhxYd3SPdL+Y9JrY40Y0pfUTph4ATUhO5QEq5vURNXODnvVqKBXs8w
YGMhjEEUHlCkVolaeMbr7q5bBAFxfhdLy0waSllpRq6beYCkp9cke9Xqq0rFsSs4pPcuy6+A8oCV
iH2qmly7HQhqOAZhMaVfEdpzCRpjU1CRL9ZSpbFEI8Mq1XIoTbhD1O98JDB6E/k6KUyt8v544esO
CUFcKzM+THR8t/j2hFdBDIA98wdZU6FOKkhrcSVutn5WBDe9Jop+9GBRGZZOUKOmgqiKU0+LqtZK
gOEBW++w0uxhBlAMCfosP9W7BgSKopxaZaDbrxShIg5q2dVDoeeBV9oZ9fs3uG9gknmR2tePzCzY
SJQGWDSgOT9uOM2mKkTirwe8PiyKGRrohraM1thmcDWnxlUa6SQdhO7QJxRbbpq/gW5OvGuuJCci
06YwfadkVjNZ3MoEySM2JPAUYOffNBHybumbmkWlvpTXoRHJHkcCsc6H/IvO5f0m9oTnaIm8/wf6
ZCCryIyr84AvQd6Bul+Y6ug/lC/TuUmrVNR9mh3GbCNwYWnspvyUrtoHxXy3DAIWPJYsTWM4CfLX
9QNnNaMtD9rPnYgDBWaHyK7sQMhKLSyuIEtBjWrA6bah+yEz4aY8okgwudU72flDXDzRpUBkXdXy
9UANu0CMEN5ViU/h2tF8LjVx01QE+FjgetQFIjlLW6GsAeFW/X7U7m3bLxdM0sH349317dDdOTec
nvKcZQaK92xlFyWmVwSK5QT/GvFU8QWPhMou7eq4B6XEo0Jhi0NXFDjpuOquwB2B+RxNofiAjGKU
H97WrJFS3pxoHh2x5z+w+iXy0TcCuMT252F0AbgxIdFUT5tv483KPwuvKrRguhbHeuevrAUzCiTY
wiPkjxHUzwmwZc8BTx4ZA1dTwJbQeIKBSAYpLXrM8ZC7K2Xnf/yZMGG8gkwChr5NoAG1itXeCeOF
4xAxN35OZt/pl/CywlMN77eE+e60xzMnwpDUdtzTinXc11SD4w5Q//agulORuBlKRkJAu/GqicY0
N+KgRGEP4AZ6kEpyPuaSOxPVi0atkzYZZKZYZE2UnO5qRqmDzgGlS4i+3tTfNZRG5MvxEUAFWfic
VouYToJluS96cg1NeRAH6WyHED1OWPMWKQv0/oFAs3rMOXo4p6A0PcxxwsyfkHY8M+r+7cf1Jz3x
Xe1gbmi/Qzj+/dsP4bG/ZitVnrVpsKnf6wO2N1Aftb1ckk2Iv3GDuXiC/yKS21vFAyIe28KxBjqK
lxFz8SqEGLIHB9g5orXr5/j6yonXaIiGCQ2QCvVPYVrvEooW0PudCfIRaKiUh4+0YJW6LjQ/f6H+
MW92mcWlGgWrxzK/qYME0zMLThXBbbsDvuAlHpSb07fu4whL7pu9/1w0vku/eg/+jqotgYwxCo2v
8KhJPFwQt2y5+EPh9CSiTnyDT6lfSUDowN/4BmocBJ58oUj78RO/PVIUkRruoG0lWa6XH1HCDHjr
WKv+8seYc9Hkq3s3o1Yvrdr8TRFXQMk6xDNLlPQUA+G7NZxUUJD1jLzb//lTiwhb9LBCZkQyj8L3
/LDWyr/R60pCQkUVruwcihJrIUcILxrlez1NlwBQFtyxYbTQmDCSr8e6V6Gew6rvIqgczrtzy0mk
Q2Fo8/20AvB4sUtklw3xV3SxMRxlJusMUxkSUqkOml8NiKhi+L8Nhxiu+wzTiw5G/LZkK7atfbMw
bvXU29303Qtxh0e1sw3Q95vV6LpBg1CdHcWTFW0xfymsHzV6T9jLHB1nJ5l94IhHwAdbi0mVSfPL
WdqKkULJuactKD3cYel1Wpft5WW3YGHV9pJJVtJZtf4n4wS/I9W07GDFWVQgWj1TQFmIZSgoyIJl
hTPgLey9QJtgIaKu02GNzM3odWka/AOW/fxy8tyDxSxu6LltjOIwwFSL4vnP7hxYlJzY5BzHJ5MX
rhax+Q3DwLg621h2C1fJ61brfQEluFwtnlDTEoKmojau+X3w+xuSRDKxwFgB5ZY8Pkwyry5jSTIZ
YV3yzW5+6I3k4RxWT3VDc8PNdcGp5EviYTBCYzneGqRj/gl+Ro1S5mD7b/Bn8sReyK2LoHqOFG0k
5Ioo5Qf3aaM1+UAk8cHNjR+ECYmEM9O/LqMS3Rw1Vp8Z/CY6dKCIWrMokG0VBG4wcLm1X6AOWU+M
JUg1S20LYm1nv5X685jivYB7maugUDX5iPvVS0ox8mXhiyo44E7ar3t305Nks+TPBD4HTx/P0KVk
VTag4MWy2xFEJ3c9DAEt/7IeGFIj2zmOoIac5Yg/OiDMAeBW90/6rqK6xgEvGGKfzcNmROYhNEpF
Tv1vz7GK4ABLEUdJgaJXkbdrAi6yYtJaSkYze3rP/UToQpOy4pI1lMAsCRCOVPLPpuvTb9zxfqu+
tO2Ow0yQzxUObq49t7kIMbIQNhCmH2FsejGvIrpG/XclRSQgOIPc1wUI3xw9ZNZ9/jYeYAHUfUol
NCcDcVPIF/UoWW6sTt9w+Jig/sOHM/2iGHPw9j1EU+j9f5lCT2KSv5aZjlnBd93UncyPbbK+tLv7
CNpwhqOecdYV37aLANe8LxFXEoi1mbIi7mtGro83fqP0FQlBLOdspZ14Swuv8X3kL5fmwEXfOs40
EJy3kq1y5BW1CsQxMMwBXf5iMsppUB+5MJ4i7b0GSZK0KVrsH57cvxEvjlQEl788JhU6HBXFdNXV
qTRrGV6xVI9pNh2c1FscA3WWk3ByuqlHmcYIcc55kjLzyvL8S4Uct3c0QlRiyYYAoNbFSKv/cXXe
62Ztik4vZiJOEHwlxUxPH0Zwz8GFsnI/L3a9mjeB099iMbaqhKEI/pjBsocZ5AFLLkzfjzgn7JpZ
SZ40Sg5EpE0KRI4MmFodFQ49JSB3GfJx0zinN3lwwm+X3HEmQToOQhK1lZaxVVq5mI5uxEoXJEdV
IxAAszufMkdd+LrazggXyubYTw+nGbcMFr5QQZy/9wNJ9qSoWZgb+31LvG9IXF6AcVzaaw18Jhd5
+HxRcA7nsIpXogtUl4viuJhZhahzW/kFDT0mUWojBv+m8gzRz0pgbEUZKXo+zNvyI8OKRWzQBDuP
ROxlgUiqawGRfR+f7S/tuW53TqUJsNT+FLBYpdhxLJUjEXrQIMQUu0vbuQvw5vnZt38zoxj6na9T
5VUbUH9oTsWlSSVn7Ry8dVdwg3/ulp+rIwyk79xSjTzTqb6mBpmYbRH9M+TTjPZHGUreyzgdPVp0
GPim17g0lgQhxVa73qEnjzoPSOQnjN/SiLgsOKpNSuxx3JIap6t+ku3own+W2v26p47fglolGwoZ
gxPupx2r7daH9efAD4KzMHlo3cxe1iiisuAYtutcrcir4h38siLeC+tiDMc4hWu+tZX0OYgsBvY7
Kr7yHnqRfu261Jq9R71afgqIvtTNz7fVxuVsGhT0+2qpS8hPyQuys6/ug7Zd6gYmm7BNla/+t+dI
hGDEQZ0BLMbtT9f+MeTakSPBgXuZVefMiFAQMyTqfGg5RbXuTgpnGmYHjVC/Zn8W6be2197/TVHd
rn+NUc976NydnxFZdZ0RxdI4FkGQHsKWI9jSR6hpRQUlCcXkxeX452Fw6Qwwt0BfrczkI+O0tE7B
1FYzQHWg/EdpNPxFhcaUxC057p2Q+34V76+Xhv2aer5lp+S3ADFtavr0XyfXQ82qvIlff7R3LFT7
C+D3AYQ1zCDWsMb8SLyF8wYtkk0/mCop2D4Zt641I6ctGsNEApRjUKdsZVm0Z73B8t0+NGdncpf0
E1f1Fbug8Yh0V51fvcGRGC3r8KhtR8AirhyyFv5m7UfiwW0IinVNZzqvqF+sZ7/np/z/2RadzVZv
NgLj1H36zuJpy9H9ti2htL0QQluuEdIhAE2eZA4k8g7sERE+cwKdusY6spH3UYX5g3wURXjLJDmX
OoALY9elq9pyxoGd4GoTn36+sQZOa16SXkJfSy5xIcs0tHr70W/qDRNMxftc8PL0plB6c0f336qv
MVdDYVisCdf3G9aARJw1sfmOFt3Dt7ac75SPAshpodiTBufvhM/GcXfJdToDS3o8OmG0BwQWs524
XkGHGFXdOqq+SiejmCON3hn9+wQY0D9m5XFVo400QcuPjIKoVuO1qQ/pz/Sn/XrT5FFE6ChjFGBd
mFOKQtYWdX1rjrslihKemPXt09X0qR/57LERLiLGyDDviGnXd67H7/vyPTxNNIbPZddxF2AU3dDu
NDAQdVAP+epipD8QbD046Ivj37960yrV6w0z9YnSYvG0RKDDDVV4LO+smT5HRru3j0EcN0rCY7Vb
7ThfdZobJ9ism0GNG4KhFga757j2/SOe7wTXMxlOmqZbfWiLCW951XZNf1jdN+831JgeohPzi54V
6fvMW8bey8pNnpTNg56dB06j0e+NE6gishkeKwFlcKExT6Qz1ofncdAfMCp7+UV6CsFA/dhetLuF
nys35sWP1u7K4uTpEFwnK40dUHtgRAYarmCtc5pqnekK3htnN5/9z2UD9C7n9f5ASH4GhIC93Rpj
WOqaNM2srqA7OJf82sA+NRd9gwBXdDk5UC0FFlNryMlbqbEjceY81q4lPjjWgDB3pL4hAiBMbjYP
H6Mq97iEGwjgEcyx7yXnkpyifWKax9TX/il1u5IDmaTfHWQ++mzO/BAarjGS5g0n9rQvB5eLUd/7
7jGqW06NWX04GOjRGwJWXdT2Akv2Hh+SJynRDor4ASn0KMR7rbhEbbi2iJ7MBXy1ZOz68vv3nx9w
KLWmG6uLjG60nJV/Z3ABRNWycYm4a/d5NaKT2LN7Xw9IOaIGrIQSD5CjXb8BjLHYSN+EjQmAQvhQ
WBQLDts83RYe0tVUwLV+FQsGayy7QqNOmIy4jEkxfX5Cko9xFoQzKdSs3LDmcG3EBmezfbjZa7YT
NiDSwEOIVX0bWXw17HSTfyt3dIvbQg9sUNA66WN2jlz+lLtLGdZFeQAFaqOFXfjuxARUvCM3Y51y
dJ09PS2N9kziLfXyzfq0gW3CMLcP0f80KS9j3p2A77mVydwh3j+GBHim5ynbbKHIsUPOl3wFsqqy
/q9CAlpu847zXYP9Sufj2rN3e7osxdE4tBNobzci/pVSrk24dlxNCxJeQ0dEubLgUOYtD2xfDo/s
X2PgzC7tS8ETkT3YbYRBAxApzsVhdDoM+pFlqiQrT5x2Mhc4UgTGq5Vwo9eE0adzUoyRtIC8OH8o
ToTsJ0YslKJBp2kHNlT7spmKrbukYlzWH7rF9+F7SbEAM0/HNpw79ZUuibLK9oGS4Ztwo5B42et7
MVK4EaNlws7tEBHNpca/poJ58PM5iWgy54hoLh36jpk30BDFja+Ll0yHIX/Ynr5x2prTGRXea1u9
hcM/7jBSftNFqaLKoA1/PdTLyYRB/aZdaKfUwyHr6deebvDx7SF9I/W29NyNLAivtQ6ZalyEMnr6
uBvSM/Votyc6hkawRgkBCBxGHGEArlGa6yQAr2zyED69XgwxrZD6gGshiFZn7563KpidEvH/f9og
Hc9LC08AOtDYFdy6VgAcm5gBOlL5XXbjqPqp+QpuvM/2vI2+j5TvY+1JjroSnezxZAZ3YgrCtyoT
8NtAdadMLbi8lWRVY3aE3jLFTjHEwPSVllo0YKW2yB/6QS+TQLzWESCoW8rPWSJlj847xUJr4IV2
rbOWYbDsnI4lMIhs1xfVIZCDeM834a5jIL7QcCscCWkrbh9Slc2wdpBslpLUosrvpeiey/1RlfmX
jzNtbQerwRQwj8dLDWo0SQGAIPvt0BT2qKrBnNVWzLjBvGPTh9Yxrg+3uIOBptKktNcAAXBqs2d9
ssErxrhJxxg9zqS4sHxdcuClAsDDfpOZe0xVH4rPNR3s2YjMEsdH3B9ObHWrDICuaUHvDApTSYc4
+C+VnScXlS284jNYV8O6PeUt2gqb49csXuq2I0erifA5jY58YQyycZXTjYEvST5rVvwTBPkmEgEX
sPA4HZFIleq8GEu0Ax5o1mP89xuv6dZ9J84PQKHQTGhGYykIxufKDAVSy9kpt94ft0pa122Q1ZO2
LatgzDpbg+uW8Hw6obcxqMHYNOy09MfXXTqser7aEhT7kx4Su4syKBw2UhYM+zOcI3Ap9dKAw/fL
IQr9yY4D/IoO+K+dm5sOpBfUfZrVms/J4v+PGUrKU64yXOF2dft5S4EcQwHayzOR9FOAG3u3MTGo
7NRCy3k273BGRvZs8DWdqSzk7rI04tK3FcQZhyC55Ic7jd9iOduH8z7dV2HoPlLk6NLDAtJDaXwl
eLoT7dWP1UV7NpILgaptHz/zc4zmf4Vq4YY0065s0F8gXJ1sGd6a9tn1GKc1NYTLSbirn4sv4+6F
cWOm91MiZ0vx47mOlE01YC/fKJRQ7e+259WY4/5nhogMwpWegAZXsdnrmHTgcSzBWQo5C4fEYGZv
6tDBreHPpbFZkSTzn8/3UPPXu4hPTUXOZUSyLJfo2hqoZwveEPOYODpKxUMmYjX0YlK1iQHKP2L0
nZ2rGBdaH4gz+hciEoYApkFuA1vz+Q96KxCCtj3yq/QYY9i6N9rj3/9HXZzxU+RydjeTGrtRhRIa
q2LeDV6mEz9Im3KOUCu/WVrRm2cvgo71tW3tql/DViPGzYf2Y7+UTSh14sleYtXtrX0mIuj/TkRt
k9PUdjgQ0b7/0qazEVeFRmXRu/UuAZdplBZDAfD9lTxGxzC3HcEn4NThLOsJO5TghsoBk80l/8pQ
Le639kPP5N60v0HmOOlomX/xY67TloXjNKWGujEqOzR0LynNU+RBoSDdrj+olqn9ABW1Co5h/XrC
C+mBAEVRO5r20SmXE2TcIOwAB4CdYwHYguzR/96pvvJH9hg0yRg7VECIYK2VXDovhloSSDVS2L2S
f0ir8FGleqEo1xAXgVIWMz7DqFvK3/Dwq7psrVm2MVPHiciZNLS/Jx+e2nXVap94i/Kwc6B5nG3H
9IbE21FpLHXrkGl2A12mFrqX6DahZ9dCINpWh7Ny19aAMj3ZoG2LlDf65GGua0NpGPkAgcE8g+sU
m4QLIE+DyRe7+u7KuNg4dGcN3ma7KXyctOUhiQl5IoxIhV9d518NELx/3GQADz8yFqRlFZV6k3w8
8Vi5+snpw0gZiP2OkzaYBOwX7JZkTgR1ql9lDhpVY7r7htLwDZksxF/mrur0LOR3PU79qkITXO7p
ImIdCKUu3cFPSg4UpdiglSg/SUQw5skOwPzvcm7itHm3Gvib6WOe+zQYGC8rceMqR6K7BOgWNvXq
CTKF2x7jlQfaU4UccVW6SfEzA8Du1mnQokijoqCXxsMKrYuZ4mkzme0lJ7GHSl/j7q/R2sHAfnr1
iDi7Y9CsvhlwgIKCtB8WzpJfQjcika/vaafL0DWJXmzIHwTzSvhT17kSY7t5vnYIjLMTlXtDDJoy
8zlzVhMP+6Np7JYCVa+ZgsyG0DvsftsZyF4lnvtr11O3mCi/TmwboUvbefrFn8xd7ozGCOmhm9mO
2v84SxmwjLW5EyYLfJLld0U08y9KLio12zPMrVaW7PnOtOQ6O0c3iS5AJEgMAZ/ZHg6dlWPUB0Sc
LLpwT/IGfRul2CXA0yKrWmQoRDBv23dtyvLD9GGfWiZqQUgQXO7HHLI0LtqNWduvCHy9H9z8KQbG
VyxbGEy+2N9wDIzsnvZdskilGZrXqKhoil6INWpIanYW/n4bNMMK4Ok3A/AOGS1ETtaI085tCRSx
vXNgkCnkvQo8P16cDCd6akuSVJgT3Qp06HHX+foVGLD/5kcsXsq2UnnrNZliwy+6n4MuATYLfPwK
sk2jBL9/QCxhV4ELojmSZ146mQxu12ta3hZloaJYE9L5wv8k6rUfgi47VhE+1BX7ce4xeFVO/waq
jjs3XOmKyNIRIoozFccpBBOySL68lbfVwNIquaaN6hYkKhlxt8lxt4KlXQOXJeFekdDDwzzzbZ7P
XVM1r6klRjGuJW9bK9TS8dfrkm/M5p9MUfKWpA6ynmPyzXSfyk6W1pqZGiVntRgxT0e33v1NeFrS
mAfWRj1q/G77dYVwvP+seH4RtaKmO6hmsN9Mq/6dt8gwSBqBngLPNGlHcFi0YatkjBNqMQNEbJSA
CVJJQDDSA8IsH094kIt/JaJ4YZ1rviz/SoEK1YDV01FtroolyHp3cPNK+u7/5ho5BkgCZCK8uBQq
i24708Y6uYb0bkikNAPHOcwvvygAWdd+yLNUFczHkxgJQ0O472di8BvkIiGo5C4Pkh3kCeNh6Zhj
62dmP7MYg5FgmWFoSiCcZ3fsl33V/O10Kn0DPQfTymX1WXyORkbAu0skIEgcw4iyh/u4jc/s/SjC
2KPSbO8kTAKwAidB6baZ7x+UlsF90rEMpEzOjfPC3wjIQpibt6mUkRYT4mGZysn5Vd4OnQiCwVwC
2VdPbCcPGy56hOGj4JinY1Ml4nDCEe2Dqb+2aHj7xvu254GQczxozpRhLTNbZuAD8JEGKX/WCMx7
s+dcUM1M7bwzQRgSeI3PnvdwVTM+iE1dT42bUf2D6+QVkZBex8MutSR+mQjHfNDQQVVwTHoeR3mF
zKsLodCffO5GW+1yqY3b0iSKV8EerNyBEm2Gy56b63TEmnLyRP1PkLXrVf5tO+S1g+er3jmxvTX3
Hk0w5lPzhL7D6IafkX0bMcRb+WafmDYndCguqM2GFvYRnItO44aKb79LJr7F3oytgolXOkTjZOQG
4nAT4+ugeRxq8kJGEem6wIzcV6HvbKwvjIF8XtkX4H0+W01UjvPKbAr081J1OgVfT1zFArqsQTYY
4J7sM37xptGr//srzvr8f4x9yUiMDr8Xkfyl4bTTZb/oHkQtNcVKeaea+sp8t3J9LHn0hgRdEkbK
W1Z69r1ELoWWuyy+KA4yhMxigSO6nL6AW4bLLkA9k+YrutiYOw5fWTfNFEvLLEg0FlEANfrGGJa2
52gc3nZ6ZbvIS5msm/0qLoGN4P+qIPNhAxL5LeNJUNgWZrDkp0xBCvsUVES6g98k3KJGO3rdA4aQ
+KnMp9G+h65mvYOJJTTNMY520kVco4Y5d6fCqpc/hxxtQiYDRTjUtJCcLFVwZLtCyVu6TSqaesHs
EguFgCDgUtYV6TULU5FmRIu4aNNVbjXZ525verx4xjx3RIDFbjt2FPXZ9yuuqMHrV3SfIe42xH5G
ACsAawSq0FaImSGL8jeALIbWsjGUW701dyN8yrDajuM336QBGlVsbCuiaYF+Q1wkRoQhenReNEWl
cwMwOuJ5C0p68ShyI1TPj/+pMNDyu9Nq+sWRwjS6UIEOMlzdUNWG+TAqvEDp5LNi1v7aRll5Wl2z
xT3sDgnkJihg9JG/nEMkSTsoKmWSYT6p6B2/kzc2oVPG63t7bn8Lc6y0qaTu/RbKGtY+/2QzQE41
TApL26p84V/c6b29N4PPX0FUSQriJ/flvv0f9o0cnbctxnT5HNHSdD7YSKURwgAL7ucSZqHED3NK
2Rt2H1DtxS19UXDH4V9NPGl27WhpvAmHXyfZXgS95QNGnLhkaKy28ZunVejjqWE1Sue/kChnTKoT
1Wvs5J12GMvcTroqHBOx6Uwk+TwDtk3lesxkBgD6EestE6SzF7p+2kDcmKtcYmflklpFD9BWcRWW
MXHFbdoOq02vhjII9S6cUdWtGh8Ev6gzKTcD/ai3IwhuIrI/yvv2ABqbcw7jP14d6fTUZ7XTEDlP
FnANbfGAyYDAIK6SVWoJ55eG+wAVpDE1gyD5qqg6uf/w3UI64mL7PKraxbabpLz/2rGvzoFGIZnV
12pGATUskoqhufQvSitmTSemudtj1lNGuLge6cwVlvjpaSKHdCL26SwbbQyzO4wYXW679gK/aLSJ
auXywyEkBg5vXh1U+opEQ2XKko1TMC29jV3tOB8ZbIsnxP1HXgph+E8Qd/h80KW0midG/+AN3UYq
idh+lNC3gZN2j5VVcRtzNxhjx83T+6Xlp0i7IjZ1qCRqCVjpWo0O4U+8J2pnR3zfY5sHgH7LhmlH
sZ2Qoz92UK7RnChv32m0ipIFp0J3W15H1EabXDP9dcfrJGgee0HLqTLtUYmFE5jdfXfzI8PRlxA6
FuIDSlY/Mq9Dqwx8QrpcCnEOor+lXh0PWEWlNfmr8eRwbGzLifGrjz3d8V9ioobIafscn4LlUb6v
dVQdnOHEZtdXqWxOOYySmkZjnRptlWxmOTEpIyGDfI/WQIZ0gg8yNyOPveLeU41d2lZ8KzWxBOgb
dxqJUEz0s4yaG8l/tuSbIH6tvkBE2jtMzi6Ake6iT3dLFpIodjlWOnzYh//5JEmuTdsjvFS7cr9o
kGO9QKaKF/sw6S5XhEiJUCErhlsABSmtSLzJFbRM5i+xKYIGNgbbdyjCfaTgK5biWwtOWgEV6AJS
kjw9rmWYj1KWRstc1U1B2rgCCBeUcTQZiUznB2byD5p9WZ8nJ/ZXgdqPIz2s8412rkrExuBKoMmQ
oo5PttFYv2kr39biDiRpeSGkEpooOixvItOPttkNvBdKlxYHCQGWxw8Vd156RsC/aqUiAAndTRFI
xxc617o+dKVESNrhHD4l1xywtKUP9NLAUoR/DtvEC/NJAJaHJUGP2/a01idb546Eyh6uFAQxZj4i
rbN/604ppNQ5MqSqYuQY8Xo+J7JxMFGi/3sbhbyYPYI9rO1wc2Z2ETmxwtzXDHu+V2uC7wUNYFX/
5QLCodY00hG6VedY7BdxRlM8VviHwrfaPnqJK8VxdLqrO9BPss3SFENcXpNlfRMY0IiWb9jvpVtQ
LjsHK8lEpdycDGEUrZOKtcp8LYK8+4fKUs9NTVN2qphXTK8g9Dw53rLW8RKcad6wLnssRZJU1L2L
rfDUHUm5kb2l2gd8adcAheTCfGq3hhGxSx2w+m1GmLFW/Y3aOItDXWDkJSzdBQkBASR91D20538n
jWGNNtHebm/+pE12hLDZCgQhYZpfPtbcVkjyyCrWLEVYopiptakPp1VbMfZCQRtWQXjWuPFzVCZT
KxAGAsU8xQTIem/qiliCXQOgjEWRCuPAxltUB4ogmQzwVvJJ9KKLYjSVlG/YYykUjmBHpeVb9puC
FLZ0Cyir7ujfvzPIuRUG6GFRjQQBEYMNGMm15jQCmFw2dKroVRpf/XEynawPy1tw3pmWrjk7KE0h
mQxCsEB/TYnN9z91MlsYFk+lrE85AE0D/NdN9Atd7/JXIuUJpHQn77QYH0UhqEGjU2ycrv7EbJKB
F2eMyKchQmxV26ccWkVtxE0ZKeiNCH7rx48YwXCBX6wW5SKdGpb4bot/3ALT8fDkkc9lr3pIQ17O
6avyr1kZmRsnoAWbTgL2GYmEjmIM1KCJyV/fOgOs9WqFIxhDGI4quXsP2ht9QgyZjBOD6Z3KYgLv
kJu5E0aZNaZaBkPyPVWimSxuKt/DR39+0aZgqrftf7DouboB/Bd0pYV+eIbmlPjEEV2UiG1gFOVu
uwhkFTAIS+7EFNLQocKsZLBXDPqb6Unya0jQqReWvsec0Bcug7Nzgf1NEal1yecDEg+Y1TJZq9xM
OH1MPzEQvTiqmJlbXRdIHBfdQBaaTGWpbKNQ+T6/KxPy70Bu+PCYWTAJ4KlT+zCnX4bCJN+91vxm
oDlSVDhFgl3UG2/0rZ6OZuifGMxdEi7FGTmMVCpD0PWUJ8nB2H6m/Rn47eJsVA058v41l36xqfhc
iR12K4soUEuGfKLu8xYaTiJYD2ynNNvduEJrdrDVaQ+Petxjl+aAHs0dKKXQREvtfYWuumVZG6GP
rH0ysbrtMCW5hcGLiZLL+qHsDLDiTOvKpYUKLEN+WJMLFWVr+XGy/J7fkLy6gcJLbZuKnDCUsbqd
1km3ho7+UJkHVK8+gfGJhBARZ/fX/738KnFtn9u7u2robXVGFyQ7BqKBjYwNdLH6HIZ7vMiaGpIG
reNQCymzuZfrakZ6zcjAu8gzACW2Qpd4TBXJvtNwJMieJCUqr3OtEf27BJONELrOi4GK1ddX4/PN
tTPYZtVq1YaJ/GeqNvs75Bfd862LfK3utANcM8Ein+/8e3xqJWjyZp1h/qhGhtrZ/ZxgdCi6ZrsQ
A4XG8FCyG/bwwsO8Xd7ERkyC/anYEdb0UYmrDtsQfMLHf/AtDXi7slYP9l7am6vH2Mk3nSPFleQ1
0GwezY1fgSNaPktaRrFNBUbicBT3j/UncZyjJJQK4seKxCXKWEARRSAinXQ3S1ge+r0wNdhdBXKT
uBlvHprBy92s5ekqia7HVyv/zSWhYVJgt5kM2QWbZDihd3HvhNhANYwHg/Nvk7lyl/anrKEsc73O
SYie0HuZ3Hi36Jy2kpMru9KIwl2k0GLXi6s+ZIf8hYZcYz3SAEr8yS1MI5VfnM4BsiccVd4wvPsd
RV8uWJ0ay2ib0DgmGFyPBV6uX0GtvlsqSQ6npngcWVqeWU3+UfBqHXqAH4ZrIJrK5R9OXsUo03po
rc/ZstwD5ISVPd63/jT24NOsTPg8TExQB3bR7jecCOQuGgLaepIeiOZAs1W5sIUtZKHe0xpElf7t
cq/rAhJsjj3tZTKiBpmT/rlYqwz9y8GqUX6eWqzx4WNw5gd7c3t7vqjHMp7naxnhOPmmwlVVP8r+
60awPqHOgXEWkVv73KvQrNI93CP9wD8Q7BMMzkVLMDS3TeqAg00sQkvhh1cnYLvN0vqxL0yU+6FO
0tbCEaoKGyQAiniBgYj164XoE62BT8PMn73INT3rEwcpc5Rr6QyTOcPhk8A2W7nDwK9qm2zVW81y
z7j9+acVM2YShh3LP8ag9SfJkEVSpVLDGNGcZdr0cH2Buv3cjjaT6dMP6oDwrc/HCbUOS+WG2KlI
A+1EZMpmN/OYd7+4WCypUF26sMofRnglngDqUuKJkBGCgnZfHB4hPpKm6D3oUgamT8n+B2/xjYK6
NRLHgJRwYSlPd9m50JfRjv2y6yuU7Q9DEI6Na34838yFXuBh16hHcfllE/lTxmz0Z3COt0YAVhp5
3vtWfPJmpNI2gQgVQlnphfy6ukQHfX8kcKAh0BKunun0UsKKzOqbswMXYZLnDtjKR2QIw3zOIaqG
eW8nc+vI5WFMxxXQ6O2AErYwWrVQBFQgwobZ5uVqT2fB7uRdMfYDBScI5np1LjCzXZKJC1XQUNIz
pc9bQwlF/Drrk9qduFSgPzuvfo7RmdQd5d1b9MQ9tgGedh+AvAXBi9CyGB/qDXdY7zEUwoF34YD3
cHMskfhb3TDUDDsIbeUelyR17U7f7tyZdFwTEjxRV0IocUmk8DLrU3Z1YratVSUTaWksy7vVwmTz
tf3dsYHbX1kGpovii54gXpM5V+GkXLEWPAdQ8kVlVHBA/bbgNFGwuAcNZdCY3BrYX+dljva+AP2/
GcYwRntlyGcYWQmjWRSPFEXxKazL8FxOE01kuVWPP6TseV8Q+0g9lbcb2Ctx+DOn2xd5FrcHd4kL
GFfWsO62m4OuSJ3Dp0mQBwfxWLPVpubzRAkCXfqqPsp/BaybSZP9eFW3hi2Z3e/tIyFK+GBUpOLz
YRGSEF6C6w8s/vV6B94pcSga1yYVJsSXJQYBzAQl8Z/7k6eE9Sx/UftpP2HzJ3bp5FL09Eawa2dR
OLpa7puosjWtBT+vqHGEl3cKELGSWUQdX8Msx5V8ZD8SZMEacJfDuv4zOyTquZa+r9LEIYxZOv7m
Th5Vy+puPTDJYYz8LuEC1FTY1+2Tssfl0zNrPUXvtQVf/rKR9NSoRiW5lRCrRgdZoN6DASDZD81l
IzereTvAnVrE80rDi0sxEBpsbgBbGKMzFZ5GTDxcNYxf2tgrkfiCnFmWE4bfSTo/F+LpCZfA1asn
PHhqtULUBVC4eXn1xCAJM8HbGiENgUdGGc5bKT5C8XivYEkr0i4qHFHIexg2sWBHnJPWpcaHS/ep
VAl8bD4H2vQLsH+EiBB+hDZKVSp3YnFol2zsVjd/XoY5Dmjke2TtBX2AMeOD5/wj54/YBQKj+NTm
InUZ5NLF+9jxWAFn2IKqNL9WwsHA7DrfVmfpb6gNsIgz4ypNMTraV/Z5Vgfzg+eEBsNWqMsCfzBq
oleSrP4v7Rzn/dUHNPWb7oBzSKeb36hCDdIVbD717pTlvUc24Z5r4/P/NdMPHWvx0dvrwBRs3d/c
RAHg2+xsl+fcJdWlHIitPB8pWbEeFc3V32cxYEfTpsMPGqA7qEBCI1h53kMyuxyFQhBrla/68x/K
O1YpPddyGHfI72ELtSKcJfXQgRwmqL59mP+ZmvmFNyFis1eXElTV6Blp4jJy8tGEsIaOXnbmh+sZ
Z/J9cMnNAD+bXBZu1W++W+TgWBw76Q97VzNqsLAZh+Xwmf9POqbxkA2rZigzb96r9arLWu3BTvbw
nYfpQslCl5GP1kIeqME4417Pffe5Y6OZ5iUUmvfMOilGLptTPqvGItWMdyQTBvAXiZY+7yBAwAz4
3CLPQlGXqCytqwc04EVbaOFyKsx1ancMwm1153R69wuw6IbtqgdDdm+sZDAfu8l74hdNi/y/JNgK
mGT99j8YSXR69LoWXJ4sJo8H4+UO88sCeaZbaFg7zPA9JRAusox5WKEc2up+hy9nSPTn8Wnqpbwh
tNYeGDihe6n/89s6bEtVA+AFPhtB9ONRxSxLOHD8azAJ+36WlSW7HpaoERjyK5GUSNKpXO5X2Sbh
4Fnh3uz4OtLcI6saVnekaoCGjn+Ylv3prQnFuUzq6rqVxyByuN88/Obk+hdBCr/1I1l20whTiyge
MrOOtRnG3WkPPG9Av0jY0O+jP/M/Wla0MT/rxH3Y6f8xY+MGL7IBBcGkQYeF5i14J7NvfvyleEjR
X/9eDXtiuyYxWy7bVJeoksckEpRYS2U9mCMy87rON/cL3ytzPFcheB9wLDmk1sFYJYDFuKDlxRC4
Ve0amWfaC923ONUIC1cSkPjmPDDlatPCgXU1Kh5tY5hYTTwa0XIrtPjZDPCWMt8PK4J6ge+EhoJ1
FA7YKjXM6RTpBCTjU/CSoR2D5wy0zxXM4c982Neo3CgtGDSGqLVxCrUm2RPQHpapbVc1H8j4C12n
HpXMrLrhFT2e53gWXS8u8AlnUhtrKM7culgUNHPvWl0Fm3N7/mdlF4elf5ylJbLEhHQoaOamdDg0
h2JSlMfbxdpypWwHtUa+HX/CAdKnjdmATQd7aKIrEiBaSd+RaMPF5HDnljT3WqYLT6LaJE2HImqi
dL8zMI1rVIr5wM5WBkjdteFdHQlLCZUzVY3Tstnlor5G3mUuKQGmPXUm2VUnplZw0yvYSeJuZDXE
06q5WtrCx7usPQCK1Pu9j5YLfoRolJ2SREOKc+J36bpUMvwndyX5B/ASWhvYrqcu+yuIALJ2X1SU
GrTTCdwrLfaA6okb3buCEhcjLyR9PszHPAWWq+u3Q123fhyK7m8I3D0KoWmJPFDsrrA5dRyGKof2
10Z7ufbxEJUfQDU+0JtV9bpeyJmSiErnteyDasGhHH27kSlc4gmKjbfFsxHJTpb0y/esqTR4pBny
timRcJLKxW//2zbo7EZjXn2F0nFDWozLgj6diOM/R7g1vczkN49htYni8zt/S/ZCS3qFE6V5F+Fn
iIhpSkPtuvPIMd74VQDnEwWSA+IKVakTZxytL4pyvb9DB6YmoskPA/M0TNRsKaCiLqoaEt/hOs0e
dxfqq9lPCaOnWLHaLPhYr2tJJ6Cn0k9ZNcX74aDcIXbwjdn9WdnBhui5eV3sLPLhUKSGnqjZkLsl
zzL8qku8miAb9AlDb70nx6YOUrv1PNEseCD7xnJnwYkJMA89RaGgqFHBWljcOduSZU5rgF/HnJEL
I5pgIcQ/Pv7ZSba+va1qUvnIEsC5p3Gng7TeA2dPqHdpPWxEpvgxZ6oWt/3/8S8ZvFl8cH7NfrnJ
CRg6hjqebx+u7ma3K6S9wGWE9fsGfPSZrfQy9+/FIL3f3fAOCt9G4KQ3L8unCRaC0NxDn5FcpSF7
FZ6tTdYG8bi0VcwLjYtLV3XZ/mSchXfGz5dBjQ90fpL2/teZapJGLj2O5ieCALJj1hQEGT8lZ3ON
zxP4Jkaqlh3i3KhzFQgYJ2N2RPl3biL0eXAORhctrwUierFP0G344HGyO5lhUN8t/W0iV/aTMQVY
8qKBrqrS5Srsa+tyixxV+I2qHrhKzCHI6ClJ/VCyUKA7W2QgT75sKTFquXQVeOmSdM0KAYYpRCEV
BrCO2BLgzWecs3T4AVZ4d1yYD3NdQbFKfsEdqU3tixkAXdrBkcCdi/fySTEj+ZdHlLYCd1zj2JcX
PF4o58bYTkRRq2RsqHlfBsc5hlKoIJP5AjOKkkqYNZsT/+RBwX3XxcaDpUTUX+sUvxe+7WTaJ0bl
7jedxCa9VpPQWWkXyUROBzE825CX8HabeTLoPzLbqo1+/umUkkM9uZE5i9/FgPXU7HOIJM/ZAEnY
KGTA6o8LKCntDr0fHWu03MCwu8yyx91jFET20sgunr1hyzfaAAAIfemmPEIGbMKlpxxam/Rn8wMM
w0E7JvCLax5SZti5xTk9aLKBpxYN0Qzrd1bQp5zats0g2SdGkW+5HxBgVhG/+6zwDHEs4NVRHuEg
Ufg5oE7qPwTMaAn1z6R0M5W3yhs/lgnbqy3qpoUpAPq68c7O02+SnS6SKFpW7kKPDQtGHjrg5HpB
WkHl4115mKvj45+7AYl4tNRfJukUBGx3YWez3WkZfjrt6Zml8iFlBc0ci2zoDjW49xiyWUiJrJMG
BaFeIX24EAXw+8unydaI0IyxxyJO/CM8zDylkgRx0OFkMWnc5yZmkf+AQkpp1gWRovgI8Sc+AiUP
+Jgyy5S+Z2am33tiCk2Gk0FqrW7IUv2jBLtJguNwjLbcy3OOTuwvRdwA5d0D1RtwO/prXz+ojWg7
Fe/cE2DiJbjgSNTqvERXTMX8aD6LvlNHRjcDak5x4r/txWnxRGlC1gskFeu64+2+LFl3kqNx2Y3m
0N1XdgPqENJ3jqmv9wse64A+E374Lwv3PAQe3l3UdMEDNRm6m0aJDb95KCQbpyKMnmvSTId8kY7c
IO2Pylgf5W7BlkcAE/1YHdLtPD7Vs9jd7h0TQqZlOPaRELMET5GmF7ndXAhr0TPtrpV0Ir05iR7V
XXTmfUVFj9D93OlrS4lZ8NB3L02UcF9x/2j9ilVPBNpeYL3bq12aIAjm3wmxYkr8Y79uj5ioo+DS
s8AmgD0xpBSbkmW77AJ9klLhMR4h19hfP5uSyx0k0+cLVIwcn3wkjBUwcAMngWx9O0h0yLQ9X27O
UhjFXY4N5xMrwavuO1GlQUt8I4Axyfv7Ul9+QMLJ7GC0Bl1TOAfCC3469uCO1s2KEEUyyjzn3JK2
Lv0x4NUlIynRf34bI1KvQsVfCv4YapjY/wO/0aXWeO2HqLc5ocfMeX2htp1t5hvZedbTDuljEKor
qlCEylIufvfNxoFxAf/ONYkLJqAt0zce9agr9oCNQmIV8D3EcFE3qkMjMQUVisILG5FHP7UkreBZ
mCgLz6p4l3Qee9gZ29otfD6xruqYvrLEHDg/lb6Qx4Ybo4dqaNi7pSZ8zBvcGTHCdH25ZuxyOeJ5
5/dynuA5ioPfCHal+aWaL7gZCrOOqN+hfcLmoZHewr7VX5H4QkY5UnifKRmE9k7ZjwS4sPmRKEnh
U8Tx41UL75adwOQlFdlnSu1qrK84uX20e8ONrt1SPWgGyzDkI1/MXxrKBanxtLLFSkMN5BIkMlLv
8Mr1/jGznnAOe7oQsEkG7eMURzSIYmO6UxjAugDPeiN+jgRARl0XFjG44yqZI1LId+keRTuFyy1f
cTzNWXyI905kDFSXq3t/7ggNI+rbVIZBo1LQhc4tesaD3CDBpW3tfQE2NVyUpDrjy8V+6W1YsMwy
st7z5RGK/Xadf9Yj8o64+v1NHJd3P6EZErlID+z2HntWaWHAUoFQQmdTov8tGvP+nT+NUkmeaZ0S
LP3qAFOA+VRKZrM4OD1DCJUXMPJOh1a3lgmbXcCnNxKzRSMrRVGoOFJ6BnxzUD4Ssm2jfDa/7doY
ACX4IMZSxcuSqttwTYRdGd9kQOgmZZ0fgFkrCc+i/Np9iczbIkOBOf0KopUixF+CDKLObtYCuiaE
t1legFY0vvc1C24NJihpTRdjBlK49Fhhe4gfK9hDHS9Cb6mBWDyeml/dPUPXxfSxh2EWJ+L9OiB3
eTgGZTirkaOFu6nhJl8SLzd88oE2tdqaZ9DbwpUdvOEghDI8rpM7XYF1T9DdhYlbQ46k1YuVsbOu
6/4Q29JVodo8vHdUE34sBaGUvv1l5AS60k4CUQ0KkgfJnabuGvYENjq5CmM/PSRXTXcZmuIyBPlW
obsNMcU0oiNU6Wm5oxSwnWp6NzX8dnF/wQy1nPHtnkvcFMMhw8fa5HHVQ7P0S89ulFpj2uPW4Bbz
yBcJynU1KcUYYDREGkE/3XLeqtBO4in5fI21T4TPZpes0Jh/o+L/KjdIcqV95YRbrk7vv7jH51+H
MpMFshr3+beWXX8s4jR8isv5NMz8boTiGbKodRIi9xaM1vOprfjflMnjGAYXMPcNVnA8uKGHxEaS
1XPBTh/L/4cm/7H7plUBdjN3qEv211bLYV6euUOhIFSe3+2PBivusfqrice35quM0Cramhk35owW
wyDy5F6/Z4kjBrBhsBpZgDEin5e/NDdt5vaRv6EJnikvlVNbaYwSNAQY9GN8TkuVxK83d3EKorx2
5YNKi2UdBJDHJvLtNTqxQtIOeWa7MLlZcG+yDDlWukl8YIbuDM8jCORmbTyemGiaDLo+OiXouNiz
AdTwa/p09T4RuCkMCVgRPVpDD0XomI3gRjtSBk5riH/swDPac68GpkQtIAJYMTyE9E27n2aZpypd
O2UH2cOelubtc1tkQeiQsig9jpMDIVbTru7+xKGtLb/SpOFlJ9fzBgGA8G4zm/zQc37G1mulcB09
uyTtcMoVVjjFXM+ZlH89o9ostGWs34KGLS6ua94KhX1HFDmoLbIUOQDQ4poRyCmsdzlhws4N/pFv
syEfaGi7r/A5Ssr+O++rvyggjyG9xGRrjGoSSCSyg5KCaBEMvVe3VoRXCx94BVqpSF6qWDESPb8L
M6zR5dQ1afJZ4Ad/9AU9R+etOLCTblC2Qa9mqQxDCXIsf96rt+4LDf0PRszHVPSviSN4kfTZ0C/A
aJ75fD+Uy1nC0aHMv1/3R75wm4uscmbF57/jOh46Qo8QoEGrHhGPr5fKG1J01besmktnwyIu3fem
ZrXh0r7ly3ivJzN3QAMRa/6905ZAZxxQ7XLHZML0ijC20kxmonq3gMML2rEFq8rWQDiVLg9jqGPn
yMmVajz+5//S/tw/VnpByq8o9oQHJ1R9kMOb/WJrGe5+At9gMORDYZs6PpdxnJWcY6+A4wWRaPFR
DAUobze0OxGIKGC6GFgGEMyEs3uSxtXsT57r5mlv/0ldssYl8qoB6TydpHMUYhcvlmqu4J5tG5LM
26+zBbOLjSxfZDFZhPcD+3WyRYNVpq+nGsOBzhzBqy8LLuzKdRPkBLDqpgI+D75jy6DiD1BZbMb8
JQ56AerjQaQAGXqPUy8K+CyiuSURrIa3pvkZlbhjXU7S235PIyzv/Pi3M7/XmVQSRypSM9ECWhnZ
xCrbkFl0s2od7fY7zvObnKoUIkloFJlxlUF1m/dKJPGOI5J8cb7P9/I1nUprAtbM2nsKrXj5Qmzt
xlE4J/5zBEM1Xt6aviTszY3XQrIhj41N1Kgu53s6qjkbOWJBlfuNKwmUnQjwbIIuK9wzmznlHIfp
qfAm9CKiPmPsP9xqlx+YCKDdExGCKKxttD8fLh4sXZ1GfhpeckB2RFc9A9egqiYnc/law9Jk4JoZ
gAzn2dTgnum4rLVFraOJH36wTSWJ0Ierg5BjpyL3S30CeEco10AcpH3Kug9I0S8yXcfn4JS3fBZ2
sA23ZUprzqghhcgu9VhThmLl8m9Jq2Z2Ixn+S2BRCxpF59aJI/7fCB+S1w1i78zj9YMMcrqFXRaB
uo16vmRpOEkXn5V92/rLF7p+Fy2+TjGWy7+g+Q/s8QOEoyVLrddjaC8J1smfJWdsySIpPuTiHWLa
zzo7FIPYNIQ9MLoheugCQFzV86hMDL+IsKw7+jmXIZLyiyC6+kW6sroD8C1n3l2g6Hlu0IbCyi9s
lp3YrkjxygiH6/d6mEtnEe3Tvp6+Ey6KysUn4+npEgnyumHF2eMc7XJFob0m2nZUnh3tlW/dLW1h
KDZ/IfKhoirxPrn5ta3BvvhP9Lkr0/fbOgcjbFSBekk1k1MqO+BrH2zLtReINXtX4+Jbkk1XGNHq
kA4VBBOHtDx3h1ua9WES51Y/3IkrIRGxVhtw7kKSJyGi0miaunDoXZetA3T8Vh7X/JfQQ9OxDn8y
Giuvnxt8UwS4ZRwqAKIbeUAzub9g/QOdbxvoYwi+8q0XPD+4WlK9nIwrBw9AslkWmR34sWEcG/An
6Jum/+zn0hypNS11eheIz3kSlgHle0WctPLkHmFSKGALi/ltMuPCpqQCGJs8bGclwPx96O9599JS
jOT10vXxVt6Rpv5hygj31Jeifc2CJfNUhrGOgIk4T0Bxd520Ml6roo7lLjmftuQkYUyRahBO/CRN
xT21MOiNIcN1y5uP0pxRgn1X9hB9yMZmcHZp//Go3ET+yIqBM0rbmGeHroQcatAK2pBiDmGU5JO8
Rxim9DyUeuNQB6LAUBz4CCnLSeSKMo3dLSjsj2FkLm4BUVV/umagKZ0T3MP/veEecMggq6bbNsvM
OLjHW0IE+KFY+buGLGsOvYBTJdPOu3dY3sSzGxh2xE6+JYnO5tSbRU0hS63/rLTqNiohQAaM5zog
OIra+TRiwVI2Go9oM8zYG8wLJMGi5OEXJS8SJyUlN1AC7vggdOkK22Rrhazc4l/KP/XIBO0n1v+n
YzBqZLLGhsi99+xfGvBcj4vL570eP8yJ6LM29ULE8ML+BA6j7rOBcq/Rrtt5xgv0kYuyRzjiQspz
1DG/HEtJzEcH8Ttn2xFxvtZjAYpIF/2WbKgNUU6kkZ/tbre2lbUNLL0GuL7rTMWTRQ/UvhUaxG43
RbAvh234tuU7fqVG/59whlNoAJGLBwJxFsSux82P9JM9XDXm3/g3mBY/tgdt4U0/95A9tsybJ8Fq
vvgDqgPnCoLdZFBELQ87p7CPjG+CzidGgQHlPGpboY241x2OqNBONH76lBxnrDGfWP0i6jCUGf8x
9zFG6sVe18JWW4PODYJbnLgmte1AmxRSnpLTRYDj2hLsFQsz0465Po494Ib/Vnl3I9I7QG0/DnCX
Ine40Ki3ax33usfZylJ2l0pe7Xhv57yaIUo1iMJ2pOVyvZH7jf5FwwjzLR97/VoibVnOCYvnfBcN
Dgl0WZJXAWB6u7fmBEOSts1rFK4gqKO2QjYHTQRntkWaJ4tkcbR1pi+yPmnl6xJ1zYI2XbJFVP/+
/MTiIJtbDGGNhFTfS9FOf+/lxq30aZAwcyUK6TI4asUpP796YDRQ/uyIz/E0BnTzAL+eeKcmFP+b
ArBE+BsBRD4YDavOOSETcrzdPfpFJ294fB9vXDkAvvCs/xFa8n4M5m5vmA9o6T3bqOspSK657MYr
dpiwt0E2OdE7BsAc8d9vV0a6csAU8Ed75hLK8ta24zOcM/fh5Sz/oBAqSKirGcGi35b5xQ6qlASV
mjS+Zhe5Z8e8JBT7kQzlOmbstQYcr6zmArcY5p8felyu/O+VdbzeQ/CB9OUToT05tH6FmjpP6n9h
pXohvP45ht55mx4SAsVn9oyh4ySn4RNKJ+RzNz61VCDQIGWPk0NYjsys4WXJX8iF5bT8HQGCuZfl
oPkQO0hJ2Wt7Y5B377skMo07T2HkpAU0eNAI7+jZHCJrdKJN0tYywJD9DRPIlWs7UWXLM3waCVgs
/yztV7OFhKCd4mDUY0ZxArymelH4fQeMxP1ceT8Z751eMIuSycyNTU0bv/nVJemUDCJUCDS5ZKDr
+WvlLsTWWjJxVb/cfiIfVdvgRyTtibwHuD0iGiW0C6wNcLrOwMTQOp9Yy29BAxda+Co5i78Z5h/U
clw5NPzYO2DtllQQ7eT5CYfeO1g8Sa/zDI3O0H0+J60pagyTHrnRwsurUz8PI44/Jm+VmJX4qONl
ewmBdMTdtN0k2K2Qut+ATpUhiXoZEiks/yVoz6BsRwvVDgs99KbSYdlykVtZmcyekC32w0L1EHrp
lD3B8S9zA5iKF37L1q78Io5TFUHJjYdV1DkbR7gF953EZhHJVCPFzgoHPDpTGvoLNTWXQvYoGwwd
9srqKi2rxc782Rvd56/b2yUIEQX4d6VJwcD/LoQqanKOA7QAXBPxJs7wjkNAAWj8QZbJRADpVkQx
kmXsOAmHNMTCGjzBVoymBhfrb6kbPHDzAzXurpAuwIZyvxixBRxBr6UaIkbEvujySEvARIrjnE3q
4sdRx/AJYIuNQBOLeQq815EcJEvjCE5EwhN18ZzRgBMIli3AtpQggWz/r1z1/A3+UwbyumMJr72M
gIYPZQW3un4pJkUjEG8UXt7ru3DeteMQuxsXcTyT9/UlIel8/mvgDTKnjYL3AKpa92fMtnSzd+27
EK69+Ol3dudee2L2qTPSXokNvaOSN4AYLIZoRS5+1k0TcbyAJtb19A9zWHXAVrJRSz1XdUko2y33
ZZQwURafNvaOmgYNbd1VyW6sRvAaC/2S4mrIqVsGiTvePZG7I8VimMKERfp2uuPWYPHBXy51irWn
c7xfubSP8RS9Zeeeo6gTpE9NOkux/1u/VekMcGJT0iIyr1LpaGh6ufx+/CFewzWViWt25F6R2PZa
te3C9W+1+1kiQLaBtDHTaypZgDpMCNOiAVzwKZiVcWWQItc+ayWUtdwB/g2D+wZt7dwcVyWC3GJ5
AcORQ1te+Sca6+NnEraozLV/CXLZbVgoIn0ChBI89c9bMBWnA47IEopLUmIekeCbO9tjBw4baSHt
DiBvlA/pZqBI9ZZ2A9YxDZx/8Q0R+YIqf+NpwYW4YmDBsxSwrC0adoHTFhSydJ4/iTe5Yh7GiUW6
P/OGG1I9QyWVSwrDHMDlyFTJFqy2Nu/dJ6ffGpr6fMWl/5+5iE6+AZn9vhOvLtrTAc1iQjhc7zxp
fVuWvDjl6X/C3S8YZS9f5TZoJhKpApdI8PLDYPdpBPZe39uBo2BM8cirzWwFPeR5eCGbbp7/XmI0
+MsTjOGO0WKXfwaxFwg9Iz9b7KOrxbbf58zR25+jbCNggPhj17+kk3lzrPMz4hKomSMUgHoWIl3K
tCZQiWxhvz3Iz5mc4UqSJ0yql7leR/fCakdNvaURxkamy3La6AdcdbgBRQEbvj//bCO7SnV9cbp0
yFTXhEaU3dV1bqoO1xhZWulxPD7ptx5iPASiMBb4BWSpgCuMeXZ3nXb/zOUDKA/WV8HOq1GvKVbI
hIIOTtdfJ9m0icuTGsf4+klhG+eTogWZRD4AlA0i59LAaJlzguI7tDZ0H5oKwBaxDTX2xAOGdJ23
roytVk5ckC3vbvuNsIHsP13O666CcJh6uaHFAEJsgb75JTGX0CGiLGRIobMxzrdWliDcjvxYhnYF
OCX4sH9jgwzXTLw/7iJwHxp+KtPLDLFe2eZQiRWFfjvc0hKlaxgf8nhT3F9c+yjGxk6jiWKGfm21
L9hH8i90e11uSOFYKKkdeLYVgFCsPJT8pi1Q1vDVLQ7Aw5V0Vj+e+XOoSHEo9IwhY0ZkJVZCKF2m
0d7QjWwF1pmx7W8KVtIhRu9rmEQg+DuiLRtvvJGON1f+sYa0jeiCHo6y4Tj2ADrCkAMX2QqdCq0Z
9Aq4FMYdRf7UkGe89gauADgJnKeaCT68EkIbBg6oGVKPN18eNuLzV6ovdCoHB8oAIDH2wk9Kqmdy
sEqSJrVtcSfONv7TZzntMh64ViMZjoF5Iqx+fGW1NzbewzJTiYStcwe3aP59StkAystGhv1+n+hO
2ase2ofnG4Qf6Wz4MLq/PxlFGzDRbulQCU+x4PpZ5xT7vZ7WO0KTCBl2pw9VuTA3VMCv9DKq3U0k
z/wtfwwNuKcav07+VNOdVs4MUOZoK4+Zh0adGSU+T0Gs80h49A49tZoCjNEroQ/lMYq3SMkpd2X6
bpildyXZhchjrpRr/Lla84qb0GZ7tz74WN9dWXzKe4fex2j7Ecz9N9TCcdezbM/7PpRknQvcIzwO
0ZDKECG82ufZsbBgB2LZOR3Q1nqRYwbkPIEfUuX5hDeHMjqekQpEXkhGeLtrtBMIX5OFmObvbm7L
1HJlcps61iKFOGPtXFScFLH7+Fa5rKrgcm2+DbBZGo2ms538iI4q3yDA95aXjvhXipIW5yCiuY2c
3yyuUDiuHrTX3SXGdpNgMGspi7VbN/YnwDLQ6A5NhG8wkFkhwJElNzmD28hSY9tLEJZqSOftC4qa
kbtCfO2SkSzqejFK+rJZYyC7nrXC8UHMz4Kvkm2bxA0BW/d4snVUPdRwZwuuClSNrcLiDGosdKlD
+YlmlZlTGJM+m7Pnj0Yz8Ja18EXwXbw6iWsFQud89FNZIwh5qJKEMNaK875HgRH9MPpH16iAE5hl
5jKeZUHklbrf5HbNPJuofBhrCD72CZqZybDNuC7nyNMiSk7FlwEbQnnox+QMj+ea8sezvDFqkNpv
y/SirMhJHTWzK4rMRl9UbTSiWcONj5FhzH0ppVuytLSVrx5KU7XfiilTtKYkXq2N9qsIMNAyhcwT
PUdGxHmPf1r0ES56rtSTmx+/Cs2DrP1KqrYjIt9gGKQaXshsLFItv1B0nj24Xf6tH6sXgF63lhtd
E0F13bW9nlU08DcVERplaUGZbnuj5rmwgNnGRXzYfWf2VvhC5WodutQaMQ+B9EoclS8/i9cr4Wz3
78vDbT74PvNvVvjXe/yrD9jIU60xyAg4IJPXoPw12ODLoZy503+9XqXufkxKarzaAJNJWQgzcU+0
weFMGLJCjqZNHRUuZhghjGxjPKBzu1abZTLDCwXPuxpumdclBBrAupsUB7EZEF9CBmUC2LJxuwwP
PptPcMOoYJ0HOAW/yN3mpiJc9Xm+jstOZ2mlTI138oLQWIGhH7txU1y67n2r8me8vfy3Syfz+Rd0
GkxZMFgM53MkJ/eaxr96ly6x2VLyWhWD1wNWBffl2tP3qscIoqnk8w5/lmSv8lpNGDm8Hu5aFvna
8QuVYU6rwh5ZdV0/SItxMGSuoy1sbhsWPRcgGX9QKIpqDXLHWO68CQpfQY3XqeStakZj3FJpHWuE
TKtkDiOnnQeXMAKhQuNFlgw9bNPwSNULrd9IoQfpVH58dVH1Q3UWhiqyoabkJ/VG0/qvoDt3svi4
m1YdntCYRMxTMi7D6jd/zSre/VWyMQTZxLjOVyN5QsZZ+yNR1enAG3ir/qCP7RMVMnnQhKUKpVLK
VjlOgm7tQE4NevhlCWMofaZw2yR/sWF7Vhe9hMKvYCEJwJCu3L0EsdhGJqUrLTQkJ5tu6dJ4Fl+p
MAKzvm1CcbXOIhVWmRsoJlJaM9wSDe3509wV5gQM3bt/ZhERJkkWnYPVQMXIe0RPBwNPTW/agkKH
+KXNIAwG2S/1IhxCV4tD41NVFuZsk+eHCx0dorUviL9Cb/C+/GrV9jXExauATMLm2za8vtYXcexN
5CFdUgwlJfdtEP2a7JNO0RWEJ5P0q5eJNbDMR6MKOiFYzlzdQuWBhWFCg8cW2A6+DdB3Xmxw2rBj
SIR4nuQjk8ncXr913panSvZVPWksjTgMyN8KUxZ0mFnPFKcSS4iCBAGann3HOqNKBydVFU7TYG0v
RH76jIyYAZNG0q745PrQjvXjJAfZRNbWsOjR8YvCPBncgDNBHygUP9V1ukbn6x6WB9tf0dtADEKA
vVUcNe/e3JkdYosjLdKuGw7R2Z91dPRT1BX/rNVj+CiSgqvPyZ1yHbE87vrQeRgztJgzvY1IWl3z
nEzpydNdqbjfMpTvZf2Vus1ftgzs6s5fqbgvrDPlMdjMiA/yvOwAAzj1vnHPzo+URshgXpJQIQoV
0Yhb73qyMGTK1dEmTes+Ajjq4iJ0F4ivQQ5lOeqcEcj/5FE1itQ2VPVn9bO/j/MTJStf9/Va57FW
jFx8wDxv/Wxj8RNsbq/ddqdW4sylD2vAkHx067LBDQC64SJTQ69sGQic2dIdVlBa3PoIyuqsQ4Np
UOTNv6JVfwvU8SxrCvRm183jCZae/Sqyg6b2kAndMIqb65h0kH2UqWN/CrxA7Ta9+ZYxDtuuTRSg
qGszs1Rk316KsYoNBjX+jquLxVBBvlOydzSd+iNf54cp1Cd2pMGlyE7aTeiQRPy7o7j/WQ0HqjuY
UaZSLCGu8VQbYR8KIdFm3ftyIChUFNv8IWmeOOFHAk8uF1FHoKzs9Rfw3S+w2Rhs/IljTTEcXYM9
A9Yuil/qcWXaQoedxZvCuj5WOyU6HDIebB730DawhNAg6bPo02H4b4ApvGQO9utqlRty0uR2bpbW
rXE0kibJ4CyGgjzHdHFTM+Rdk6W6BGxgy6Xf9qC/Kup0LqlBGfHeV8KGgiguodUxSeo9D7z5cIgn
qw+P5AfZRlIrnBtUwPSyBFP/N9Gd9S9pHdZ0RAl6yA7lpBnYHCoK2ta0jJ4++A+9PbySeW2LoUtG
VS7kVxmKgyVq4C7N8nhY9uIa/i0xTClDc+/tN+wCzgMLuKHiDWPv9JXHJIpNtVP5oan+RzeaoYNJ
+u6k4VK+IEvD5CMUxn/ZlIYOmFvY+JeB9rT0vmYT9ncq6mI2TezZeneIXR2Qk6QqigS6Dk+IgydT
JIhcr8rBhhAgU6AG3lMydbgeZGo/1F0eUtS3nggGr+HCJRfqLxCg00XB1j5/jKMuBqqL5Oktzj9N
cofDWO/B4khTdy+6JEIzFjuDrFzwvKW+FaT6ClyTPJRoC1JKpl2GwlxIgfConlJQfDpk63CY+UvW
3BrojUH54qQWDpJBpozv04DpLHpeeMse9yIlK8Kla6x0ZhQiyCYHnMewPB3/1u8jt2sfTNNO/FFX
a/WSDVye3FtDe+UeIfBt47Q8imzYPPBZahxJLjJzkORWzmUXiMWJUNfVRIlJrTdamyQeyGz/UlhJ
i3LA7GBW2NWe1Qf+15GdrgrKFiEOwze/d5tc4kkEP1GLV0AAe3i88N+KvpmL/KAxMM+DQhVQXupW
K58uNMv0mlYpc3J1bELqD5t5L/aog68SMKRIjLK367wEZF4jHxKZpjAoRNGzmffNh9U/t8ucH8lP
LV0RKC2w3N6pAncBq7H00+p4WnKhI+PVujkhn4DdA0Tuw3a2mUDXadlBeX4FETIN5gNeeswPaBwx
CWSxFkGJzSop04nfLEc8oUAAUqLG6N3nJhzKNcnL4v3DwKZ9qfNUK6h9yRPbRu1SVJeEPdxfjJqg
JFLJ4/igpQUa70hRt4eSrSAN2iZxpmHoygDrG2ahzcVTP0q32c8+fCC2uIVaT71LuII7AAc7Et+6
g5EXuYR3lii8GqacZGIOpV21oo1682rt8N2z2Bq+CT4/eXKctsEJLfi64kXSo7G09C8eihSr4fW4
966BLHiYSGKB83EWYiQLxGinwjnSE00paozgeZyTIrJe5bBhAZiEYvYMLwn49p8GZ9I500XsSxh+
tdBfnadvX+OdpeVz9x3jvoyJ7Vwohhw52A0ksFMgGnD3d13tUU8PWL3EOiA+Io7gxz+k7j+slUY3
rTrakyaxka0ELpZ8YnXjwwDA7uVlL2qEvhm+S5XMZ/pqn4aQwhEvgRQxPMxJsUR2mMRHapOqNVlM
D7POGPQUblowQTj15EfRU8+Y+usgfbP4qW7nljUolFV/LOnqy4/qalUxJJLHHNKi6wQY4VIdFCem
0KCnWSnRyOj2sYOPyvt9cReOfW6vpGfE8ZKbn/TQaS/RIXkMM43FDDO/Ynt8nMtAYCqf1yOsGyYo
OiX7PXVrcNV/KspS2wXlaMFr8rttEPLYrE1U/QpxZ86QeiAQpJ/njyA6k+JmCV+4XDijZTvcJ/CH
c6X0nUlsiIwIFQlIyWzmijWQEIZAE/sozDp8jljdMYSOJkd1AH4YHh824WGE20kMuLXmM0w+wUzF
heifii54SAXOyvatc9o/5P2ot3tKoP2SkcvRejHgcdb08ie/IjON41S7QxVfkh5vpAdUeFulashx
2Ci0C2St8zfN9+vXf5ow13m3WZETcpFTuBr54HhTdorFCFoTSg17yFwtc1OylqFEMvgSWRxrVls9
Q6B6X25rQ5KLpa4Cucxozu3kyry3Cz22TE6l1wKaGKodbEsIUzCk7TDPgEciKqX3JFXA5FWEK1Zh
e6gYEZiHO/nAaKOUNUxeUUx4GlANay/Q4pmXKahKf7Bf7Xy4+wIC1q5tBzO9T7TTbXaz1DjLBtlD
rcupN0b5Y2mT0qMuKiJMQ53rZiJigbzyBhUAs+sk+eUqI3b4B9LS/WXJmEAURIsSYH/xS1MvmZ4p
PTzLQg78Qe7YnNIqmlK1RswEI7ouzKOuvYVzMTmyUo8EhHX911t988yzfVJJ5Tik9XaeOAD/rCTH
HXVUnDsdcozri8cY/BcU2uv7La1RBKXbQZIgynXSC0Nve2mAUXN19+25Th0d4D+V0r66Sn6oaGnG
fix2ye8j0uJ3JLwlXlow4OT0/vcEqwthqlM71/URf0G0CTH+lX2VbznipuMQ3RC+1fdwoMoKptQ8
/QhPirCWH2NxpkestzwjdymtPrEFXaSQQROGqnCd7Jt9pqvmu957JEavkFtaggZeeSYsNgG8VKLA
V2G8Lm1DHJq3JY+87LvnjOcIANWgH8edrUNpwU6on8fsBsL4MqHKgifymBq5VN/sjwefJ/t81gCj
ZrtbLyX0KAWjSUXLdUWKzJdRBV9PQ1R2yOHf7CR4DZzb5GIND6YkGjqyOb8uGXdhrZH+pmKT357B
1/PEJH4vxLjXEsXJ+8O6POMxk7V/ri3bcOzsH33qP/ENJTkxCLRn7o9Ghm4pZG7bCaiflmIxDFa3
YLXWREvrgZQarHP3Jmm2lTEKaTSD5DgG7qNnKXWhLyoawK/5C1bDf32iE+Xk3UK+QEP1Y+u+2rA0
10PQhfjsnsO918AWkpV3xDx482MYMJM2zjdPa60nLu0rW563/bMc5M8u5ym9RhOjbonBSEeAViS3
Yppr00PmpgNQiHNrAWa0Exyv2hJ+gnLaUqmqL9AuRbE3DHUHy7g37tNk3KiUBAS8iZTNpyGqUjsM
TRFqdeaWwMesKU6JkLWM8/nxjFoeS0L1InakmLLhnXq7FOMVIxXM6DlnWkoQs6/YU+cg1T8y6iIP
OpT4MLxXCwLmLG3VS5m6Q87m0FHNy9HM2/2VkDhGSEntIZEm6Uq8zgy24K9Ny0Nxk/k6Gew2kCqb
NzHW88Qwd+PbLSW4XaLhRTxbeLhAPqz2/Z27ffu6bvmiHSsEjLYZll4WViNyK/ldKTR1b1oeZsFY
oIcjCsvfJzXqPZPuOg0scSxtgCRyfKUN2tKujA3q3iX0qt8/+VQGvgzK9z7Tm9t9osa8lpEKy1yB
xIUTT0Fd+h1EguVEth3ggpHrZJAFeD9vcJDrAnF1z+CvBKqYGkWjEn6Ar7YG2k3mt5qm5qWIyOhZ
Q/s0cMvpg5YnudoTChTYeMAvnpaLH6bcLFZ7xQP6Z1RsY6o2xpyqqYFJS5DADeyrVAAmkEFkj/r7
NO8HFpAZNiGXT2NYiQ/nRzMWQgcznfHQMsLTl6WFsYE+X+qeZVXIgwV7iVc+/nSh82KlVp1kE9gZ
mDDfzPEpjeVQ/juTKtb5+OqLGlJTKhp66bTQuieshpLxSO0UcnjRF4TRejQ/Jm/cKNoS/Dk9f13n
uMVFCo1tXxl2/0EIbyIMIqW9vieohjA4sPqIbA5LJniAhJ3RuWdjA/+Gg/gFs2jLry8DjgqNG6Lr
Z3AFUSwhNKXHFdGrXkMmMbCvzUzkQQ48+Z6pgqNi4bndM+8l6TVfNw2C++oMCRykOooqrrzwhwB/
Hh219jgLwSLYH6V7C1pSAds42jzJPhoXt1B30ZKgYXB8EnoVJmlbbqeRsszQe92k0pbpoT/rB4Dm
yi1azjTNw+aFxNvgb+Gnm92sfzgftNmmWlsYS5nHyArQRSgwni1kbsXUCz8ZwJAm1o3w36sg79OC
Ebc8IzpDdFrMCr0QpVY2/JUf8qEqm/bCln1HIcJlP4fL2KIBLSmlZDbLINRNtTIav17w84wkTwlH
P3O5IFs+zMeZCTDEZ9+o+nTVhuQiotFytX13SGpCvkPue3Ygk452jrJLBqu1c70hVH0xnmNX8Cgc
srUWmHsH36c97cT667P012S2WeBMmQo8Em/78wZSO+IPkNdAOpIZQpxWyFuP9owbt7yPzGS3Ol32
d/r/lkn8ez5PjnhPfYbdLuC0gksqLjVGfcPIPRBHwBoC4LzaNEq1alWvEcQmR2ahBIZ4OzZ0GdGk
le6fo/XVLH72XjAT5YgazP1lPHW0gNF2C062Veyi0OBAMN+DSlSs0HuC3015a1h3HzimIWXNzKaK
Nf9XAjXoe0jRmGpdyZK0hU1PNtWeopSO7XJ9wHmr1pfSJyIiEU9Yj2WdFCWxhPohIUg4C6LKFg1L
PoBWZhiVyRY3P1k9WWRsGZTq+9tNVA118avQA8yInkq6A6f8aWw3Hxzyp75v/urK+DY1CitttWxR
IgyM7wlMv1IUL6/j5XcFEprCJKW4LWucNvG8xzbKyNRO1x2OG00dfvdpShk+O20XfLOvMu7A6BfM
LO/+uDoi7pQ3Ye46vyjMrfO0YN5llvZF+qL8sK7Ne5TLw/0S1I28Z9EWQWsvJsmz/tsUtbxfsF4O
f8r1d7Z4XCfugHZZHSmrYhxZVhG00iL2v/NkRpe5N6Y1zfTrhp0UyOfUxS66f4Hg+xC+pzf46PCt
lCPpFtB5hEPQvSFF5dl4rIw/Kuv8R54n82IpPEQvqS0+SpVXOx+ss7aO9Dyn9N4DvYKZqqS5Ub68
gWE5aC5I1WXWKBVrGYnUJJjbNS0CoBNI1sGgzahHuxWhxbO02+7xNUzO2U//mnNOEyQTVLhpo6hw
4wilmqCKcls/JX2NsVQEDtrNCLg0Q2PrCmL86+7G9U50eoLL2EDG8nb7Mj6c4MpkgHksUN7jgOWl
YGPw8tzuWvcrmMs4UOtLn8P4Pm+BQM8IzQFUe3abt0pno8a+LOypYPIpVLDh07unFYeYZAg8ZsRh
aWzmVb4EawXi7XgdcJc9OjIQc4Fq0aJM4ps5z6TlURdftZvipz/z99UhczCg0HOh15a0GOUF6dRZ
l7qkdNd8qAZVOT+d087Dl/JJQwSMcIFiWyicIGNZnFC7W9OAMSGvpd/oYPM6kSQ3wKAP+FEccxkG
XwoohADnn/rG4kjQkBIuU2EuWwi3gyxL17n5vkGshA6HG6sNSNd91p5e49BbsrxA2VHwtsIkkiqu
3djeD3JXrUfzHY7LSF87fYk6JftY6ZeSOuJOyZUoXlAU83lv/QLmj0Y/5eyOuxdXqfJvNgtQ2VK2
8JEjcuWBHex79Uac1+QVqLfJwykUEZG98UF8j0NE+L8EKUS3FuI00TQxwFsvSskiG5oCNu01n/W4
F/plfDJZqpg6xE5hnbmLYG272joRGZfO7G5U/QcqFmWzbVhORWg7orVuB12EBSqQfC20vtrMhh2t
lw8zVxPTRrtt5msarho1CDm/3gsxuCY8GJOyPOC5SZ8w7fQIkqnM0rsm+qpczOfSrXS/H8VC76KO
ScsUVxo9VyfbaGYpXGA9Ak2ZHI7S889FpaktvBSveBNlvFXIKTuopZncRdNozoIIBli78LJIjY/x
I1BBV9NoMjwPSTyMMsSR8D0XEErA27CJ9oQ8Gef9NDUWwP0c9kUdwjMGbIU3seei7G90vdUGM7Pv
84sYYINAiN8dRxon61Dlt8q0ggGtcY+dnhStXspPZ5UBLiomBPtOsAif1k4iFSPDz3uI1VFpTJmW
NSdrun/lo3ZWbb5nv6ihbSCtzOjhov59h76wvpV7YoUVbmiokqG2qkEjZsN69oz7VvWaiS4Klgsn
gDMKcG1EYGd4ZLw59n1UEuS/RmUlJf87NvsAVqgah0AoIGDCSPmcn8HY4ZWQtU4YE7i/DKytOBGj
yvI2NTn8cvLbMl+jWRWNC5vo/ad9/dI1F3h02OUtDqBsLyPmivQT2vsbhIygambpvWKBLS2p2w8s
W4BLBugYrYe1hBC6xVQfhYwFiU2C+Av3IKpBhz8kjVOUgONF3xBu2i/ty39tJ6veiXfXNMXAvELh
jE1g0rUwVgUbq9lId2mTHFTGWBjHcRgpw3QK7LIxEAWM5azf6DqW53TMtRPZbKULA12ugP/WN0f+
FNbIfzTmCKrlpg3UN6Mp1NSk/e0GlJLsoC8MdrwMyXG8z+M8qwOEbUBI4rSQ++5ck6gYOIjjd/xk
c4blUMZ5yGZONwIJTUwO59DPbOwhveC+fVVEAYszWPKsjkFlDwXGiwutWJp6PP3btMY4tUZAHsms
aKnUtgqSOoCzdQAk3vZEBcqG4JrxN/VRvlEJU7WMQjmpWT1nithdW3Rx0x2Hx7ValTRA7PHri8/j
lIqmXWvtWKOv7HjcK1/MEpHGLTpCyUGOsEf5ymbGqyGemM5kHR1s3I/rQNlzYwjvLwA+b5DmL8Ao
0ozd5m+DSMvHhcsen1pU3so/tzMPSGINVV7OZJawgUFMawVntHg4MBhKnm0den9a8OsaMib7Wbl+
x/8NZ5WgolJMykKQH0KCLrfSsPaS9QR6eaDN1h2/XrPETqxhzcF7nhKBT1lunqZ4FBmKxzkDs6no
d04UhlaR9uUqPpBh3RI32kGaXoRhnArYrJKGj+wHbbZ9ZoRwG2cOqZ/ugRL8u2NlYWZTit3xi2Fs
er7KTJc065LvF15VxwP6ws8XqvG0zqeQhBCWe49rTo5zcd7+iM4/z6ejBJK1Fp/stBoSG1XJt/TL
DEzV1zdnUh5NtVGZl3JLHiMA8yOu6SeS8Gl5bRnfjooN5YFm7MQs8Cjlpq+shIJWW/2eVOUT+mZq
QW6pARe2s5rRGgyNBiLsblcSzSnp09OPkK5NReUSn4njf44B40W3Whxmn+jHpcpGFubqTfZdvIvT
ABWwNlVlk7qEOgNo2SZE7APt7JAmFcvECQXYMdt5tP56ryunGjEOdxJDpq19We3trI8pjOeWQ3To
kTZoJrvTDdjrUaJhjZ+wPQqOQO/+e6E7Ru3kV+aW5+JZYr8bnu/jjzHM11cJPYWD9mpuWuN61Pf3
ilDb+cB9n8Hn18VHQh+5RN7nnOeDXNqnjDu18qr+vx/ovghiWMQfPS1yqPNi6mf7k/Q+KH/HacF2
oDwVzacKXub135S7huyJmq6eYdyZSbDxj5h0ApImZF4T5g6iPgfv90HNE38vmQEYPfF5Z/TRCoqW
KsGebKaCdzYgA3uXiGrG2v3HyAah+djx/k635mCq8K6xOqqcIvHyJczO3AUa3NOhaKRBhBgG5v/f
XtAQOWb7F0NmESJGZFsssOK/qqzSNV/mGFhZaC6c11uspIZ0bI9FfNUKGYdRmFfLG3mvQ2dqH5+F
8rgA2doAxfrmDoO8DB2N7ivWZWUT6tALDgWX5r888mxx4ojqo2lSIHWVd9ioEpZEO++1LfNxzMRe
zKC0ImrvDO3yqDHjEQGD+6p2ukkwAayZNgusk8C+/jAvExFGQ/RWZFs5Zf/keOiT26WcwME1pRrn
+h/MlD3QfJf2rAGZ7HOvQpQEjaFz5WvRFRlYRsfJXKaY13J6SLWNZ7Z3Rd8XjgQ0jqTHJmEOrnb5
J78OT+Rkq3lpb1wYjCcdEv0oThqqVJ+DVdExS0VQb+KY4P2usShy+Lgw2imUxBXdbsofIEFLeBE9
1nLpMpfdLV9aQtDtrdV5g0foOFFBanQ31Cc6rVrseER/XeYBE6f2inGiEm0wXKwjWRXCw0WAKsaz
eE0FBG07ixE75RPnIyQK7WKBDgJEBOOCxdnpRSL9zERbOmR9MQb66tjM6UtZJAW1OBdZm/EJ+X3Y
ew09RrWr8oAO4cZ3QRtdF0ASI6szVlb2nzv3InyAldGxKM6lxu30Jkf1CI+2KjdCiwT0Ibo9pFzE
rbW84cBXyUa9b6U3U/SFJGESlhSREdiSifbgip3/EGlsBdM37OehoZvCNatlTZXudQfUh4OuxpO3
ewoTwgY+DuRcZUJ64Z7OEjsO6b6Vk/V7lA509avOgJgWDvWgWOSDZi9oY0bATMb5IgYN5zTvKfsQ
oFcEO245YkyUYGz+MNSoJHMeEw73MjfA6aI4SOo+atzdd98CntlxvLsc+Woe+MboXV8IGrrz1KAk
gSymm8Qe5iQ16EikjA9N7Wd8M8xDAqCDMxmspXrrfvMA8XSFMHXYnjurvGydsCTVjZwRkrGpUJg3
BjILmtskZtWC5S8cFt563LYbC+MVV6nED+5sndvbBufThoVeiiHrBj+NJ6c6TgtZGKxNbfbVxvxj
frkuLAFGAMfF3IO96mhHLWEw15C7revwgaFkyqmpIyzYTNi18wFeLtOAM46RSIqfa71hiYUqV8yM
7jZO92V0lunsoG8j4/GO6CjbB38tBlNDg0JxdR//95eJoSgF4w0oQ7QOe4vfpUriqtlOy8a9O13A
1Ofiru9qTj/11DY5BmmRn0rxscCkvhPkawwG+E1EIFDMc5WLwxzaJPb8eYjxHQUvqb8ye5v+XW7t
yZfmAyv8ihmk7FlhyTaUzs9Vd5zzYnwqGtEqhBoJMnoa4a8Qiv6YhnEivycvgFgCqrc2RaFWo3j+
QOtGkYRdynfx2kiObmLF5pVkrlMa/4ZolyKbFk1Fj9lPjcdQ2QBEO9YIOSzoasPYAaDdtzanRrem
JefG+hiBth6clQEujngCcmAJJp93H7pARglDg0t46M+JZcjxhk1fL9BHC5yTL1WLzEiCaySPVTJE
uWfBhuxs+P9UA9tYOb0NVxF9jxBj8uJjgzx9/eubHFFtfUf6hNZI/lNkZnjeCmwEBhdIxnw0Oyoc
JCd+Fg/27zOQlXCdwdXNsHDD9HPPvVfTVDNAPoouX/s8i3gv27XMv6nWJPfjYvT8biSjdNsmf8H8
HDJwM/oC7rJVRZyUVadCgrGgNXlxFYLzuWoiIN4Zp/sgTES3zSCGm4rLbmQbP0xw5Yw3nCm/g/JH
/GEdsXkjKsjjB4iMdofmVweL/Kq+22QrOllwS5XmgKGU9eNd5zM6GRj5bV7z8sGBIrNBiDHSfGZG
FSDO9rhxv8Z/omvqrguzTDd+X0NSFmRPC3WgFRnUoGUI6GZFUT5Szpg7tZMUEZ+A1NcaH1EdrmND
sSJL4Qh2s6DkhS+eApedKG4zT7T/P2pPdXdYcMg4r6gzEn+1L8tgx881ddserYNIQmkPjmdw6/xr
LPwCE/vIrZHVOxqTFYojcUKg3I1wrBzUojQ/G3bKzGPr3QGgzzhIGetqFu2dZmLTGcHujqdJEwtF
yymH4AbeAGewtm/OBJ1Q5hij5D1CpW0XB+YLfQ15bCZfU6b57RdQpSzYGg2PVjx6lifxjB2MApSk
M77nSvx1YzFYxZ7yLEm31tKjbpWg6jT1MtiW2Yhm7eVvlhhiJGRs9YGVATXW4jDc+ZgeNskjPpuQ
zFKuiCAD9jbpxH47XXpl9iJu8LK9QmGsHzEbFt49gJNZTcU5UYb7h+Cj43i8UUgkoeeK/BC/FCGw
h7bbA2VnZLUD7g8lGstVrGAwhGcEAHwtmPHCuXA4F7k/xU/KZS9+U6158B2bFS1XaGAeeW4ULviQ
Rraei139GCy5u5DizGL7ydPuWr5hYCnvgFoTDBqJT0a6Ftqrylx89eUpTBGDuhMfosOSGvOQykWc
H/lI3sO1neFCBZw8aD+0UuMrTVl9Rhq3fSNMx+l+MUNCtx7OxrRJtkySCg3K0EHGweudGc7eQpuL
1q53gLrKo348cdoZ6BPkl0KY+S+PU/3YXn5smy0LcifcPHB4KsoT/AKr3UguVuDrTDZGq7dQ3OHx
xGWNnyvgR9v1PLEzMUsZ4Tguyvm2veJCdJ+LXxjX98r3DDrr3A69fACenEKA+hgTKjUWrqNqI7Qi
U4WrQdFI3gfo7jZOt7LY+p1/yIu7Oq7n1jJmtoVJk4NQp/ZykW1ZEWJ7ce0hnc97t/uFDyhQrYrm
bCnm0fZ564gKe01DitBlTmPNAxALXqaseIFI1F6qwAPgv2aWNzgBJH0vXS5i+CJHvKJmc83o8d3u
nX0VZDWjV0HUOgYFgDfIRpfKhMFCHa/ueeaWa9cd9gjRRTbOv9eRNM0bUSeKmO29/tbF7glN4SFa
zuRkOSSCv5f/LSt3gO+RO/RTKdRKL4LqZEZx4lHQsqDkqi4jT0a2ZIy8bLtg3fReU0XzLrq//h/1
zncrbQ7Z2DtMJQjOtSyLPsFnpNMmdFpOv2Izx3k3CrNFFYr8J7/OW9o53uD0rEoeqJbaSdbolQ1Y
lIBpU83Ev6T10FF5Wm6qvL3sdb3/gAg/RAilmJ/91c6t2EeHH+zf3rGWRSN3FNre5kNPHA2aPrl2
M2mVTs9vbVvocNHh2ta6TecXNA74Z6i7c7m1Nvl++r10j0ARVD/09Zmc6zTQCYI+9wSVFLIg8n7W
1P1BirHFsrUewKEzZ+nMpv2oZC2Zb9WxIsvykfGcrgyw3p5D/iXCmncpMO0k3qeXnU3D9Kh6OMVm
hi0lohH4eZLlQ1pR19MLsaadwHNcV/NeMKQEugOdgTZ4UcdxMYAlBUw8QolaIhWd0I6A+7QnelEi
QK6VOdBv+0ywaf1p2KlrBH24IBhD6m41lZoqrBQFFsN+QeHw5fBOW7dJL2AnelHzli632O7qlZvg
UQk6PDuQuektzXuj5R+wH0jzAiCORQwNXLZu1GzxVo/LlRioGkWtd7jcsgilmCM52jGdJhuBQ2k7
ZvNmpeCzGWEd3YGkkuGjQX/M12iRxawQ+XTX/TJyTuVy5Zee6ZVQ9QDTrma5W/hQ/UC+Ll5D7Ycp
cSHIpQWMxSEB+Wob6HczuwNgtdBuOcF4Wik6GM+2WUT1MmzRJj/FGwBii8RmGqfURBB15vybZ1+N
T2drMzNoMofVTWtCLNPGnzo/SakEcXRzBcozlm2yp9FCPhGXiXXwgnfy8XN+Z0lFld8vFXr7ZSV3
L8gDO4z0dC2oEPP78xAT6AJm3tIUeZbC3Lh3izHOUqVXR7WFp75MiuIxPUPXQcyaHsxwQezKElft
ydV5eSHBNiuAM2b0fTKdzMz5dYPIuDp5AKWVrOEEakKMQh+f0oq9As+QuaYaLMO5gDSgFC7RAQMU
yMUZzEaqEM9+0Fm6dWnJbLkbz2EGJcp5JW7YFwuqYe5E7BTkGb2jdeP+upylTzdHFFDBS1pwMu/B
0kL5MjTnSrfTtEp0YpxCMoF68qVAF81UfIfkrQX45Ozp+rCD3MZN+JKJbHUDp6wWemhZHdDO4T+u
YnqCUWn1y6+wjipkYzNymQFnZDzBoSiZDserYCV9UCbSIuJGV6OPtqH5cCWOvq+YMhRvbwuZF3ah
AFWphwrsZTd/CJCvTP04lOLh5C8HWSk8CO3T4bTTS8cWIJxDYjtJo709XQrYfQma5c8ZXYeUuwCf
2+D/DIpK0eo2Hi6y4f4jWKax09IG5XdSAqFIF+EviMYh2tJd0jiCe56acVdYSudpbUPVDb+CDumg
k8kGvSYnyxdaDelbxHyK04sXOm0VGsqPStTxJGc4N5RxNaqws2nukFHTGh86fWQzQF/JQd2FMFxX
3I3u5g+7QRiZUmeSHcAw+WLJZR+4MhjA31d6MunmMG34zqFTEyrTmwH+mnib/okeZNgu51z6u/28
82whGX8P3p6tavsbx9LpTuYIcaXgQ+tD9xXFpnvr08jasI4XaOxI13HgYQRVA/k3EiO3SWvuUynx
V9CD8APx9kxI893RtgoGDcsTgE9NvRrNqmd7JPkrBvgcR/ErFI2IMCNKfNdVKIOCNDGlgR6XMmh5
AQnS9AaXZ4ObVevxFd9yVF88QmEnZfZmnsSKObmsPhOjKMWGGlXoUOrWvke3spGm60IoV5MKzZlK
h6LF+jrcMWU3MCTUKznw0zUFrANS3TugRxJSETEcEm7QjUFFOT8cMmM7hlG65ooP3sMRRROpHid7
hUySMqwVSHmPsvrcmkevZcabDdmBKpvOAbq8aO3WYP5qg2y4w77anr9lIAULkxZPAjrWhrQTO/Nr
XVVDTNMfVRR8Njd8mjcompiITbJgxZuBj8vlM99txYvckIagjtALc7EPSQiXlkiBKarm2v4VyYE3
PeSFjGmAFHQtXso0sTCfnjrmbj3jDVk8o3owApzwqk7I2YywlINyncbg8eWJGqW6L7cel+zVAJEy
5wMi4Gt8KV5UNJQ80U5J0Tw0TDAN6+ABvLl7uzGOVd7Hln/PwD1g1COCKU+FCYTmFUKIWHYGMoDU
guJgut/FbDCboOvS++Tea/vb/9a4C727r5pq8iyqHBooCRqrCkIlIp6M55C9FHFYnmwkARI5aSkM
Kyu4KY3M4bnudMh7sozUxVUdYsXgnS3eh4G9PFHUQNs5oBma3Bg3p+o3xwqMnCNERZjOZnuomBci
W3Hc3YQcc/EQNTvT7QlNA77A1u5LCDQuOaE5VvdZXrfHrACeyBshQB68iBPQOAosmGceflP3cudY
HnvYR8GTo7Hh+Ymd96IPKbfgKms8ZQnwHK3lN6I6UjD7KjluBnVTgqRtvXpv5ISnvxol4SxORMvf
vrH9Ewh08fU82hsE3uxAwh1LOLbFXbkwJKh9G8sEtZCZQXC6V94UlBdcmYLPj8ED3FaAN4kPHI4w
xzKLHDEBsDpr6RM7x9EZGOHpFtsY5gvzzcba0qPm5e/xYNbscrdbR/98+jCmosV9eLNA4vjS6TF8
4U+QrYksEap/K8OLoJH3XhVjv3V2Vrsz90QXXBievPCFfoR8rE0s0q5IwT4NlOBVHSNRHYr+oCZU
ppAbz+VvZMubY5vrLBiSN5AukwqXO1tYpbfOLHa/KJxhwYIC7HA5HufwVwc7gDCRqv2FcYi738tR
abj2vQVWB6rPyakM1SMtKXQO4zVi8JDa+Et2QCOcEc0DM750FlRoai3a9QsnxCkZziwvF3k0hOAJ
oORvCkjfpAM4hW4SGiqn82ju6KWPq4e6EgkqJlttfjHbqwyvcbTGDKzbJmOPN7p61Y8wqfJUaDF9
obobvyufoYHGuo2hBBa3FFG+x8Ls1JSPPlHcHME/IWT1uXHYOsADxNCQVm6eWdt+l9TMqc5R2reM
xcZrxFVhOJ9ADHYRKcSQ+p5Z+zXsAog/z1iJVLB+6TA2eFM=
`protect end_protected
