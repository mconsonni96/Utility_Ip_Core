`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Oi6WJU6F52LjeoEGMLmiM5TqRN3vwljPgJFa7bW85nKRixzGEkMZctckbXPnF4uVa6/VSXfWaMaq
uFKaNurUrKSnp4XkR26XByc7VqYEv/N57fphGS2SDBZysbP674kHWW1ZJdAdX4G6/Tub88/WRvB+
/l9k4IbRMuAKUGxf808p01Q8v3aMrtGwqbLOaCHq8Tb83S+23Cxr7Bs8hXjMjqvacVLwdGHChWz6
ygcaJk0rYq+MLgyyug/vh0GccIujnVnGigKQwRCrajaVz37BVpnyYabyitrM2MLydD7Rt7e7Evbs
/6taneArYNYXk6u3tklIyGY+ezrbO2xxYJuGTw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="7eldWm+U6/GiWZZsNkwyIli+kbW2TyK2wQrEibbdipc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 130800)
`protect data_block
o5EfzS56l+UFo0Y1iFYCVJhptzn2Tqvm7lGY2czr6LB4npRVvPJIIEUm7Pi9rfSbm5ocK434toMg
ZzSqOFOyljCwpKBcJ12/uf6L4HLQchteHiNDI49rLEPHxpREt+J7iY276+KtVxkPS4zIhea6lylI
TzhsRrwD6DJ2nPqtlTXeUVy/uwvircZqhR83mBufvCgGAZM0QkVpSHXb+HZYUosX8QvwIqd9oi8p
khVyle6TgzrJUNkoIu0cyx4gyzcEzGwlm+2GjLDRdMkegOzv3jJGKE6K2c/xJqFIF0QiyWTPYMBV
Nu5U/h72mR4oLX4PE3i4gsHKRrz9arI26vnNqnU7AybOiNOAsAZtE6SEPcKRboMDEtNGJVOLOXrB
KY8tisXMZZpIsbsKlzGZhxY7MWn4cn7MkQxgZmLYuE0oUDFmRitP2XBSy4jR3EhTCJ+lRyOb5QW5
Wza7buEQdavZAXwKCeRQDRmxPnlMLVYyZkTECKAfYNGV/MeCBDO3M5yRzlTVXd9jhSKXfn9owit8
81S8VBSu6EueOX7oNSTL//S82wD4GeLZnpaq49cO5afshPxRrXh0QdnrmtzXM2n8GM/+bMrR8upQ
GbKF6UK5/x+Pj3W7NKnowSdAzgB2ZOArvWrOEra9u8jaQw71U+SyblhJ+2IrGhjvOK/dA8cc6TAi
3SmBYLN3XAIj8FI9SvRGz7RkKCDjL8qFFYXKjNDJMADC8RKaqpQGzvJJGnG8cxYeStGz6qhubi5L
ZNyyxE0VBtZYL52BIyv/Mz7tdvR3QDUkSF51IClNjG+nraUlakoSGxklEk8LHRt2ftV4Qy+F8UeR
wvdxVJDyZEVbD4JH0+7eSXuMCyMfNnNkD0cZ5zu2oBxFr7VWd75CjGi6Ybhc0RN+ajLp3Yra7L3R
LZxaT6rV34aThARkDbVADjbV0RkSwreiHMcl5IfgafrTdnjafn65IMLEmVclDg2A6c7SgSH49kie
3Tk/kxEQ63cLB8vdSYMx5Xm+JVqZFLdqCYcPl8P5BOA8iPsXz36w4tyH0FCmPcjicVtYGKC+rnhb
WR68MIBGW22+xPahi/wORtH6JxKeT7R0uTkbVCpEpqXKIyVMOPOJgnTMKAnWgcRrBYwdYrMWpG//
WS/0iD5DYYEfH2wK2/aj5LxwqmVoQrkUaPeibE/kT6tTIJSGSSgO9nz4CgB/5ywxiFHOIQrhAZxP
xRjjmjH0rxjkzTNtqcQjHA0UhML4V4anzxFETJsJu4EnZLhMJIEfums2+3sLQtIRxEAZpw6GxihT
FMySe8gPO9kYhrxTjBdDrmOgxzA5Lhh/TXcp0stHmjPv3hmq3r54fPCAAZ8AZSbHtJGOtk6duPUK
MkOmzcQhOGkIWe6uu7inpH/sunkBRRPSD7yZqgrfd64ZGcpF/WxbJx6frWs4ApkhQqStTtgCm9da
h9pjmWR51R3OD+ydx+cTPfFu1dEtjn5mvL9Q0W8TuzxZdj0jdfY47YmoWg+pfK/aicW/2rKzH4vP
nWFcaCThM8PMofdqP4ooNBthiu0vAP/MXcYc+oozkJHNRAM5fGByMVuHpWAtPdnhbWee1bq8bFWr
LQ9aL2oEezoEvlxGChlBcSsnmo5t/KDpe1N8VM6QpfsMq9gQvm+t4llc48x7krk13EfyUNu6TATb
rXAp5uoUdpWgfIVnX3GUSjGPGv2Zy+gbzY/4Y1MKdsG2dygT+jKH78AgzU+rt4Uv+9Io93l2G4em
IKfMpSswTSevPHyCjRs1/MhXm6O+UChdjZi4JhFtvvFBZvO1UeKKCIdlvere0PQ/nIUVPTn8ifzN
4hOzLagdvvZ3N0aHLz/USOWyQ0087RzCWyk8PjRbuDb6MMFcAeFaIWDmvPQLPQ+uQwdtE8TsGIUo
rveoDX40IuF9AhhBgGOMvB5JIWA0+q9v8cAUsNR567KyQbrCyEJYOc/bZyasxfUlC4NwmL2N7FT1
l7uTJNr3P2WvoHRrHSQtnkWQFAMCX4Q4YMmG+9DBpVZwWy5P0bWvgPa32eYWVwLSaDUF6XbL2pF0
fjGsW2fg7jvVdGzGDrnlsaGGJCv6v4kbhTWvzGdOxWoFo/2LHJX3f7v2KyJWqHtWnAH8Gi14Hsed
W0jkln0QUgkYHUHZSJqjNd2E5eeNuWkOA7ewtRoWnGkwT+wcxx7LuXoHbKBzZZF/ZkHAuWuQ3XEc
RlUhnxw+PBHeMTArYN69QuI4RxZVVuJ9aeyr/mJCKJwCLRjETPaJBn5W6rXksNV3gtjqhaRqm4BL
HErZDP0qPhaox//lfQoRRJUUaQD1cOA7MvNDWE35CXLR4uiHSQ9fbofR43dChkrtJu6dy1I6kA0S
g+PAoLc0M5L0EUp8y9Uy5XWY7xxtzrFueo/xEhZs/A9c16aznTWbGH9YHCmmPlEUl+GeFZEs8xd0
Zsee+8+2SBzJk0XRCcTU3DmBSxQwSHHbO+koUOItWQYm56LWv46Pq1fBSAhExEfRVl0FL2n45PKo
CEIyPlqIbOwfcG1NHDUSrtxP7O9Z2Vo5SrERfRX67jeRQd3dLQbS3vQdd8r//zihbEpPzUtWzzMZ
3yEhzK/ZBd6hY8rXO04cSEbXka7FND2bps6nyb0AMnLKDMViZkUqtMVGcAqz90SyBw3v6efmqkNg
K4hk79sm3to4a5eq1dI8V79HfZQQ9TbnQC469biXvQXiAGUZMHgY9V3SGSQfOXcmii7aoQYkwOFF
CKVe/4KCaXxQbTJDMLUczecgqOj+4iMv+wXIsyArO4mJGXXvQ8WwfwvqKSXj+uReWn8Okk+yhd9i
yLmrARi8bX7ihog1lbU2UG1W0JCnAML8Xlpu+2Mo+Ojnzjudzjj4+6/E8UAzxEcMcPWXP+6ziPKt
MUa4rOqahtFfsT4cDjNs/6WypH3VJsZQMCrXvZoCq942OV7TfaEGi8Xi1CbucfVOuuGCZ0LDF+OB
xrUfbWqOLRJXej+WmYYBot6v/7YaxYYrgXiaL/8i7XsGpD3DfR40vRg3NHusQgZ2YYvVv9ZXiDVG
WaZQgnlcM6xnAQYfcjrMFIRpcFIiXyJgjXhtXjCVArDGZZ80JepmKO7kEiJrsnfE8IeKbcQZyoeR
GZOKDUdukZAvdqZQJw7IPQNbGfoUpa6QwA8+Yumo0rgx3bXUQGaeGAaR6pBwCk+Sb0l5llMpzq2d
1NZUZqwbpeIAT22Rz4OB6E0lx4OLucTkuUkecEr1lcOjbYEc9gIzVlCEyQj7UwKDv/FjFWdNHZj1
09ysqKWoSz64fuPfoqzRPl2brLSRxHKmcxCKSveOYBcC8RTkUWaFeRRew9D27eIrz56+ZGiW+wal
ULLddSK9R1I8xNa0ZM8KEtJtRoTOhAXgA5En7syiIV4KS/UrGwwTXSHIEqTkenuLo2url/z+RQJ0
ZJgEwSMYhe5t99ibsngMFjoAfs2CDmHPrm19DGaOK6SXIiT6bNBh2jvFG/+0xdXlw+LeaqL93mAY
mir5FbmA2yy+uB3knKHOXkhkn8SoK5quFYVarf8oglW9G01s7IFuka3N8kOdc+YgoL2BBBZl1saw
VEfvbiSVGtSaFCvyKlmA9IrXKKCs8LGpbVET6Y+UlZ6EGqYLM8ltj0tRtBb86WndfeqJk7k7eZuL
qlqynQjVRY50bzPDvETBnWFvrv2MlQcSE8xkShqhy1wYMai35FO5hHehGvpRVZyqOuYSjkaIOcho
pp7Rak6W3+ZePgZVav7J49F61x0pCwQ4cWL2yJ/sr7nRFqomRz6mrXU+g7GfXC4OYsOUSWLDAeVp
pfdcTnxInY3ZUaPwwoqp8uLpnMImPkiU3reIVnyiwxzDLoKjXAnPzvL1X0+0KOMp/iKjAFpTLWWG
IlLLSj9EhNAybRcuOy7PQCnmkCg46l2c4B4LCVAIy2OapCFVaoUMQ17jGI34OGvOIg+KO1Ru0r6n
I3Po14Nf30683oBMwQAptMwv/yU0lwQ2unDdgSEGuJ/dqz5qaqFCjQM/GtW3xmB035BRb3dYy7ID
1FS3Auuhg7O1/I/rA2r28BudW0IPtvA4D5otb1FoxMkKULAseKSsJHrVj9aEWDKzIu2YlelsdKCt
UQS8lE5HH4Bqzd4M1aYQatspgFdaiXuFp7RDob/dWBPftQ7c/4jSQ+UtQEl9qI9UprVclUTku7FS
tC8gMccm23Kn9j83zMXiHfWHvWqxvUtRkf3ITR922if+yz9J00Z9zqLBxADIOWuVzJ+YluNS7jcT
jG6t1xBhp5FoxKyORo2xbRIT3LbSYPWQtM67Tvite3t+EN7Zl+6DzXuWYhuTq4+gmboDeejTzLd2
zQA2YzfRv+Rj/FFyDmVyZZInhOoSNSR46lX6XuZTmYdNnCfbLmBntCWfZbxIRMjKq6iy6CngYAuP
vdElhtXQV60FAHl9flrOYBWNgE/EDFejjGy5bVQv5wMr5Xn7RwAskCVxjS5ZzdsDvdUauNQnmxLh
XTkSKkr25XBJIRFKBRdCpZMVwQpJq6C6jg8FiJqKPurDjFBZZKugaobhyHR6iGtMT/cGVhx52703
P2/ONFMgirkUCisaHr/Wpx38Wzse9S0II0CaHWUqKO1DtRpTSajp75DpI/0eVdZQhAFgmFMzEfoj
sroSBELg3ME74yIdv/qWfxpxHqzRQ8yV2uw1V1sfCwLhTGhoxka1zZCa1gtOUFB6s/MaOgq+NxuH
Fu7WFTuw7DWLPDXGRN84NyEESGgFkHKW+j+crobGSFoOdYZr+grbcH0FUk7vYRj1wdrh0fPQXqvz
l179QKceKaf1By1RBsRY9B93jm2sGJJUJACdauschkM18tgKtopP8vuz1rz4w7s3c2tk0b/za18l
VpLmFcZpiIvUosT0n8mqHiPTsf0WXPqFmeq2rUIdUmFPuxTfx6Z/2f36WjM8r8GL1Vfsv4Zw841j
r6gbOAtx7ITE/r9j78ruz4PdV+v3FkyzuTb+jxDs7tavdei4C1L8z+jHSOhav0DPHek7Nc0P6KHG
F/SRNhZ6CwPdmwZ3T0fdR6B8w43Do7g6sQUKPwJDUBTkGZgh98hucRD4QsTnNfKwY9n50Ja3Sjg9
bO90tp/JAn4Mb74wC+ekQqvjEzlgBLG35l61I4ddxWJ4UP7IRDLe/DEhnk95kxojQMLmhSjo5uYS
JjGRHyVj9jRidK1KyqAM5utS5/ZaaYiLiQmHhzXqIC1AAry3WEUthNabNcSyXnVm4of93c8eaJ4l
/gsTmR5Uh6TMecTtiVKNANaC4QiKUYl8QuinaaBAG+SL7inGVyx68GdFiN5amFWMIbMySIp8T1/U
EzqJXhweEmRS4+ZN6rpNtZYnrfDiQ8RKfJoQ0o2ByBOMLZkfJFUJzdIO8O2F2hTZnKDSirikl1YT
3mwDQUgVeGuUXSG/BPpwzVMehj+uE8ne2mA+Dq2jhiN3Uc5qamcgjY/N1Yy6dZLZquR41L5Lv0Yk
oMRA4VyM48rhT6EbaYSExlrybRGcsLuN/gObSX9y287CQl4LgXdX+LPl7qMfBRELwgpuxcLWLlUq
LXApIRTSjemHONE2omc0E8g4IimMkegFSDdL1BsZhwMK8fTwf/dbgLSGjZx6tqvnkh6duMImv+9i
snQKAHr9IxqaiLtPz+2TGACb/koafZbcq/gziBWk/RC/9kG33Hy9xxz5LWiO4CdltJZOVtfE9lba
0bI3xtmD5OHkDGKXOthmZ/Sb7dkT1C2ZzEpHX06yZasPLcmeWj8oAFYrr+MNV5ANT/DU8shK2zk1
toT6O2l/YXcKykmVr1Sf51PbUsbpJisXrK14P3RwGxU8obXM+Kf5Z8d15kvn/pZbSihVuTSHjyw2
8QOFQT68W/7rANmrC1r41NRVoKvsdsuXx0cVZr10WL85KwtcNl3pAgnGsBRZ1V061AoPdluppwwL
XOGk4IWSBNOuG7wVcWOL9PNAChvUkFPbbdljjuOz8JGeiVHEn0ONyZDJsgLY2DzRcbyRxl5Ldhls
oij+PYNjkRvnA1zOLnlrUKeUqi7kzOOcEej5+BltvfkTH9Et+BS/ll2g8XSZ5kjrLl0/9F9oH6tx
59Plhy46my57AAg0yWU+/L0O0CoXOsA85xaJ7/RKYyUT4bhJFnH33qoJ3EjdOa5OHqQtVxFxdne6
yfQC00rfm7+0Im6nwaseQT6lXcl/4T4mLhKFTb1kYyqLfTXMoo3odLFjLJ21pU37XVsQiQjkroDJ
8obLDyJgDIpFOQ81hQ7Z7uJA8sOLsaFK0mBoIeU0mlq1TJB6rhKKnLlQvpWsb8Yhd1+T25Di7R+6
d04rbxKOcvjtOO7P8YNNUvG23hwTBKX3JGxrHfvFuDBV4zphTcZKISDMh1pt7QeX46zR8IumFwLf
59v1OiRvBYUU6KV9+OurpcGwrNel7OekHYr57S20SoKMchipQGErq74Az5QRwEibO/NMBvNeT6CW
hUiaHjSUX6g4XKBaabV9x5He+snghCuij8zkHEXN/NYqnbZhK3tVHet1ebdtJpW2eVsBVe4LaNDM
e7X5cqOy0OvDd/vI9VjJDME52nS0bITccXxGi1Z9X4R6WKphT45QuSfpnkMGtxUu72FBOKIAucAm
PsyQTckfI56wWoIM8mU8VHn6tDyuQ8ZCGGrfI6TErvjimFm/XMqLxW1t1hyB25Khj2zSiOMkWF80
5nmMLuKG/sGM/+PHqhhGKq3azoWd3OmDl6r2ai2xrcz/XnyHkjjiQXG4uSwKtfUAmykvCxTJQxZc
6KlUO7p4i33vJqt5TxgHCWYmk1PVM7QKP3DvWqXSnfyLLD6uNctKi8RHum5iidNjTx/zjfx/EMbu
P3afWj029jSw9rxcW4pKLRZXKzxJq5xixQ1vRtRV1JscPR7o/lm8stxr35B9BNqdzZJdoY7R0sfU
WfveNNdV7/mzP/K0vxZKBME0UcYNIfEZzUtWgN3evlkkUYabGPDWYaBHqxAeix7nHSX0sUMrMQGa
aiZFuj1rpyOoKMuZjpVsQx2RbMX2kJPJAayEDSRgGbpGpqQo1y4Sa4lw0oZbvZlzsuwIF0k01HOC
/X3fGYgFu0EjhGlMhU6XwoKdxzoiXP6l/7YxfiTMf/RWbcVuKC1gGLkT7gi0Hjp4LCmgcPkfYZ2O
fuLECNR9Ihed4ARR1NUcImHoW2l6kzNjpwQWZxRfH5DOlOFNKvF2corg6woIdnIXIKu+sId8vAng
2q1hfXPbL88MBEhGSsDmodvLBL6+bZJoweBIuvWaKKhD1l84+zVECVe4gnRvClX4ZSgc+AblJQid
dp6OphY1G4vCsFcdyz52fuu9Pw2BwUxARZhzzd6RrUVRLa0V4087KtRQlE3Egluaes8D7cjDU/Ls
j6F6pouYkZOaT4SYDtVemA/Ysox1vVgRWPkbV8k9qsrmNr8EuONPzT/FSya6S9hmGvJoZHprNP3U
51qowDJebPeIdAwKw6b8DPOuwA79ByMuJ4ENCswrBtTg70hFaTdeqkzN3cm0gtY0/kJP3rZIhDmW
7IpRFVBW0UZeEQeLT2hGv7rY3lTIB/BAvFvkUsZih8YjDyvd5aial+hXhH7Wh0rDTCujQimCFk5w
j+ONM0fQ6B6xnfBtfX9T2m6g65IL2fcvK6/jqpEn6gIKJrO7X8B0nPcZj21U6D24N5cfjJO50LP9
/DX1AX1ZoAJR2FfDTu2VvSuSb58bTjolGlgJoz9SVFa7VNMb2AXYZcHQ0cbeBtqVnpMsD2StfpYX
uhr0GJlplSTnU1xkiaCpgP6dYNKQQDLQ1Il9NXOlts7lUt7eLd9Rhu2w6xSEGZm0cVwRAqLIakjV
x1THJHL5Pq1ztOvAh5CORP/xihGV0Kcr4ZQs8o99rEwf0KyrWtR3mdxI6PmefyiQyRTTbr+C3Lao
fhob7fzYdQAcygK83rXu9n95fY7wgkSOZ7bHokitQhHGcHrj8SArmfL1xS0c7kYJ24M758Rss5Sd
BZhff7vfUZO2QsGvN6afKC3ehMC/GG6E08/LNMOfejTs3aoSmNM9qyqrFrXmuTdavKjyPIFrDn8w
Sw5sStaYbsMbMdtKmCPuXGawS/TKmrxoS10FjVaydZcKYTrze5wKMdaFQZggl9LtDxQKVoKvsU6/
hzxfRPtGVRRzKnWN8KGE/yCBZckh+9Rv4Lyhk407BdqluU02OZII2k3C+lZVt8CCQk77k47VreI5
jzXkLmYtJDio1xa4x2bQ9/Sjs5rVMkdFNk+TFJG36ruV9a6/io/O3grksF05VyB5Zgmb4wFkUEgh
lpIV4C6oN4NZqh1y4X3zUN/UfgdpIQQa9AxDRzWZokUQS8bq/CzRWvoF/pJn9fCSK5x3JL0/U7rj
jCe3iQOdP9J3B/aEtOl+eHD83H+j5m+RwUnUCk2/87/TMvjA/Q0dirvXsMWNdzLP66dSuklMXd40
5kMVP276CBM92i3+Wvv4jPyZkmjWwoz6u6gfbA71B1hStAo2ZdQY5+delNl8JuWVbc1zHdSvtAUa
hVN6FUc6/IjNKAdoYCcifSP50r6BvK4N7Zf9ondPaNY5justVQVP1LL5g123ECpaQVBMfyh0QxlH
0UCFnn7J0OoxK/fslyEJdilpb+kk7yNpl9AkO8foTctxk6ZiV6b9pJzZ+4D2qrVQAnAYgqFCeJsV
0cQcRtNbm2jaMbCDaFkFvAecBN82AgwMJx75Ned9aszSA3M7ZXHoxgM1kp/uJegq91TYmfeuwfAQ
dJHs1UlAzoC9LVyCzgIVMsac2KQPxQs7jX72HSDBpAJbpkkOV68Wl+RmUvkCDM4PHj6uWzE7OTqv
rf2tu8lMyvQnyHGu87cRUO+PHylLBrB2XgvXkHhK9VxrjDUPs31DYY0jWiYUVs1skNJkNk81kw1Y
H9WwGvJP9KRJ76swJPMCzMHL13raCGaLmAcjl1ZWWsybwJAaMHo8BmFc++OU+Xj9oX4/QopBQ31Y
FDorDV7G7IXqqR/OrNdia8vTlCljX2kdsgxHc1mx204PQ6UDtGytJAZ+iOfteS8Py6clN3J437+k
6v9C/u/nDob4ywgVMIB9S5Z/JiAIcw1ExwRSzLfzGX51ulgeNTM/SSoptVov4gFJGS0kM0a1Ob0d
zNiWAXyPOBSvdnLl13jhC0OUnp6ZY44N8HHBXjn5SFnOL5gLMj7mqJ3W2qHmCe6nU6+WEnScmi+E
DFDVJtxDwifBzao+Grcu7eM8GPIgffrFVL2XiLH+GnzDuceDfk9kMgiwfQgSJHajxIra5GJXbFh3
WzlpjwS13FqXqQiIz45+3QMu9NejLH1Gc0Tra/rilZo1UGcFCeG0c8n6OVExKstkdem/7wBYlVQy
5+oOYU67q6QNKKruqlZQC4iXGbE8XVgK0YhE80TheMmBPTzYc57hUvPVgewD+BCyKY0hvSqEmDP3
C87eEoKokTbx685jacsQfHgiXnYj5E7KmuDP8zUEEj/8w/X57ALKm6pU6hzJNlU3Ac6zmYO6CEXI
jNtGE774oEoQW552QsNmmJZxs72SsW30q7URSHfPpi0P8SwAkkb3Ru47MhZbaeQ5aRhT8xNBxeX8
dYiiaDxGebqe4DQIgwJ4vJHwX3bgzyKK5YwCRLGyTRP4dpenTGboYJDEwQ+jcDmW+iNI9AmmRgSe
GxrQm7oIQfEmRjURY0KPmNvrosaZlctU0txih1ooNvuIhAaWS09rTexV+XiZGIpmb6lT4rLxqAvW
7vnBlJiN6MAkMRd9nOxAcXkedAD1vzbNDkYbDzvZQdXDa44ZZsVeCwy5hAqt8qJgVWm6WtTphJqE
kWWcacO084HQl7HC9viu5Y3C+gLbvVD8PxxF/VXc9NhBOXFeNTLWeBA0mWCXQTKb4kRgcqjv5yN1
JbnXefMVTgMibvq390D06n38xtQ0eaoXS1r/4vyfJ+lW2bGiTrxVhWySKnTeUhYH8iZT92ftCisp
d0pOJwmrbNw8CKU/8fTj0/UMA+xMOKboI8GaEsbOTtT1ZFuQX59CnjxbrKR7wpAORhz1cEzFOzly
6gU9XWMyFjxPTJPtJqNwaEH8Hi8U48G6ecp+h0PwC4aqiwiSFEvYkZMQAaP+AUTPxJObN44BSHvP
Xa+psG+DaqqxY9+HYu0AQSbsWkD3dcc+vC/NnB1aDoHPMfiuX7Q7wGLjHEPRDZiQ9X4dVWLGmeLf
i3mUQ7djoY0wXbULsfArmOyanT2wO9dRGestjEaU/AdPBA6ydR1KVgkWCCXhhh0S5GZ5aMHpAjWn
6Igbf37LBlL3iFoNBEJeoLgFonmuKzc7kJW4cjsh8Ner3idN32UAGSqfiD2ZzgE1ssf8j/Pw5WH+
ODVflsiS7/A6LmDuL8rVFSmBh3VJAnp5q7SXOVeybnx8FRmspuDHWC0bQ3duwn3PH+jV6Tzi14IG
dYDuaPMxJ9XP2rVCZxtphnd4CqgxJLtuD0wuFIlOGYxWuNk22UgJzkzvYDpnc1Ka4H846zK/Roqi
6mdA1qOy1/0nHr12tbb9VyqtA2SffsTLe0GY6tD8et+aOxvdwhzP8JcHZuht7jM6Xa/dk5PwoQDY
kb70852zstRLbmQBchKxXwi9ed1/465Kl6cbU27+kObRnFiX63nDLL+g64gFueWu3kiLIRYs8Yjp
QTLCdtkF67lUvZ1fxqsGcb9U8+eWvTrA97pDVRdkobbNUHpphEwtWn28KAdmHLaJSsLMtoT1CGkS
OdaaVhS+jj9O4RdcL3hpiCxNuLGHhbVW1A9YsRqB6aVNpKat4lfM3OoyvCm6NjHBNcLSyBJQfmhZ
dY+W94tFVqtnKsBVtDT7EMjHBX3dNGZukLbJNc6knlBfPma5/lqY9R6+r9RHPG37gEmnaINkYp15
yH+qgMmVN0zH2W/lc7wbDarDbtldZwUSycCnXkgKgJbIBCadrdfg350mKR6fv4nATwZxy+4UbCEP
beTW4dBu4o/r1GK1EQ1unmo9LTtD53obzxPoFVQM8kC0c7r+osSUOr830Oo3dgL7QldE69+m1Jp9
4vAt0MAmpazWPPhNny53XIYRFHJlWBN9qjET+be5TYDSYg/kRjgbgKRDlqXcZZLtTA7v6TqeuwUQ
UZ1Q7giNOF3e0zP9CvzlIwJYfQ6ZZSZ6PmLJJfNT1VZCgeJSzC3C9yDbxHb7z4/py5ZK9eqJL2Ow
4a/yq6dEleso0YyTKBBAI7fwfyhdtwB6dBQnoKXnFUOT+cnmD+gtsQbNunA+FwCBo5sL+kxWCamF
qzZzSbBqVJwf2cLgOZhvjINp3mlHxSIpp9GaaZg+SQk+AAcgspUQaA4NelGj63SNtl36Ulme8RQg
ahzFxqdzjpGOwXF+fyhCTmupHfNSGRbIDzlL5Zc8vUKw1Qe/R1EA0vbGQNjwk6aAnbiDnk/slHbI
gnI+J1TMZrG8oomK9URAO+3RATYpfQ8AdDmEsrlUNerd2swzzDb2L7MxdSBrYe2cbSoLAWkQz2Ts
rv+mijNoWidie/m0aV0awMPF7OLCQfL82dN3+kR0ANsfwAFmh7sn2oMEig/mSM6sMua8ge5w/j3k
Xqx+SiE4b0RP8V4csYj8hJO6g2Zrz/8Z0DCGV6gpia+piMeKZSMPrWKZXEA4LsYdDLhWf2PJy7rh
Gf2yL3XITmqyZ+XJM1yU+fslikw8aE2twWUPAxFs1miKnZEjE2e2Koz8+45ewf9HkutgiTHJHRZo
kIziCSIrozYUgegrEdZCZRtnSZwhGs+Mw7W0l5aDFYYcHzoUYS8E3IPNNGHl8TFiGFBb0FPs5/FB
Kva9ih3sUriLSAPJEQ+aHpCh9hrOS0SCGfEZCGIoABTrLy+0Y2UwmZoOIU/L6YozNVEWgf96s3um
e7c4a9Bu9ICIQzR/1FPzE+WfGY6btsUQttt+pHzNY8VI0FTonr2ugAfqcc3MEcI7+oZmqPDp9tpx
ghWsOmdivIAPKGLiuRZCiFL+DNWSlIAe7msAGB0vnleBTzzK48uAsw1VgwKxm/SM+BNhh08goZhj
e8y/B/rgXCQ35OSr28IyqGQSHSTNP4AKhD4aagVjqDWXF/CXuhGIMKszV1wSOrXNwh7M/Xgsbzbe
u5eAX++W3oWU9m50A+atZY9Dd7cld2rGhGNm34yN4bAHZDsuNmyLXVZmoOAr5MRujywE2I24P+6v
4C1ZSRCzVRaHOwqis4CImwjwPef2SXxp9jKnvTiRisjBsNwtch3YxZx3dTQVvdJiCWXfn9QMjQp9
pW6rh6/nf0neBZ5pAjVRMKhPAeAu4V5UDmNZmwbw2KC4gYMHhQJ6++8dYl9HdhJPwMk3yezA+Omz
zz3oftnsP5bBKGo7aNPLlssoAMVkEi/QujkBCXD/aIznJgprY9sgaIiYFa+GXyMZcO1bGeRD4JGR
EE4zvT+L58bpxSMHvfdUxJsDchzQ2iBGkxKKIcI8lhfLcPfv+EI+E5ZB+r6x2GWBJbOLcqrIudAu
r2ZxKgnN0WDC3LUoLBYx2Yv6ZGbkT9PcttxI6ZYI5yrXqPKqrH/a1aP5zFbV7NkMm8hCFaIRn3mB
e5Ju6pCGRM4do1+50KcMaRsgE76hZs/KEwRIx4y6dYIxawCud5PB7ztQc/DyKVtPfsGu+sbi7XQE
7ZEL8bUeamEUTDFitMl4C/BgCw8LSvQCG13lfmrzo9hpkClXVLwjSgegRrARd86garVyNsCecmM0
QQQMI5iOsM78ZHqssQh40UtlDzGu0cdpM094I6upO/wH5uFmzPnQZCSz5Crob8S55pz3xnR4e9Me
zKs8PQqbIQN6IwSwORBO+E3XcjxrWzxqEts/TThKo4btGUlthRohAArc6BYqdqWLnkTGfCqf1NlO
lZ1V8qbKB0VyciY1XaNsPrGCBfQun3Sxqu2Gb8xA5e7zZjxna36yMVHXSeQPDSgaKfhpYUlqVd/G
JoHkRUpMr0q9wtjMU1xkK4dtEyraQn1IzWccjjJlpsXUwSrhCBUoL1bqsJWGgIe2erR0IrSJxMSe
OrOtq5o2p8pIsPfhEcH6M45RYwz5arDFFl/826NyaK915Xnyd+5NcN7YffkTzbI36P7gWZgIuzw1
bUDteQ4SpNbnQnx5P4n8fcHCcjMtIeJaRzwkLXY6L+Ys2wX+g6sELxhTVgp31dxlVdNR3LKhlyNr
xXKuiSrxMyHZV6GA4Jq3r+/zguOsdAAyKzD+M2cJ69RCaqn4Gcvmatc7LowdEFyPDVLtIR+l3K5M
HZrduEAQcCs+uVz1jgI56n9kIM+PEXTGZCca0weMnhuleQumW0ZJmXRSqQG5si/7HRzmFAyMQym2
RmGOjWXv27gdflmsK4DVHVljgmEHLNnmqmFyVcotPbK4tXSl+HXFGG5M2nsTjpyQSQFwtuwxKiu+
8wMCOdcOsboYjp+i7jQGlaBWVCdDk0/GWXatGX3nudzG3x3BHIkSoBe7pPVURNZhHz10i6G05whM
Ie8XK9UNK7OdYNt/w3jJhbP9Kg7cuNBeGVjG+YHejp2yRcufxDUTXYSVzUV//QG3sOJXwHqsq0nd
SULlyLAOFHYil5l8N8ExVYPP+hkPTw2J8tKCXX50DJWXXix92eSyewuylvwdHXz9mcWM+++nkgcZ
KIJ4NkVH2rEfIvkByN/kLaxsb0V9ZZCk30R3W3CQjTl0S7iKlw4IrVpNzmftBMMI1f/jcFUhSASi
yHciZlX1xxuRLH2uuVsjuBxzQrog+foFCIgtCkeRvu2nO3T82JlBxxd/lPreKZvSg67rzYl0zUKO
BavdnfR60V3poQfDzqs6Xz1NGgbZwbMkBOvHxePNZ00bbrwsvFJ9GXHGqbrBkO+MwIBunlrEoZbA
DurUTZFFFEbvoZ1CV9av9L9D5TGLodljUVMinB8fI3ouw+Ui05GfhDR4SfMQl6XJ5LQ363OPP/SI
Z+OKTfgDg8NA9WBB+gBzmdTr20OHcJeLHujYSECdJzK6boIQxvGavlQqEwTZfSk9AsLaTZJKJYIJ
SfS3dpIvPRWYcA47ykpvKw/yjdNiGgQLNxricKsolxIRu8iOH4zivnwFrhJDjiTv6KgnEAkhUDyw
B7mYG7zxgBC87sZ8MBJLMh+L3xPmTHMo02Db/28zhZUd6xWnecdQ77qAWim1SRGW0nCd7R1Y1poP
f8ZivraCZ2LMmP94t/+pnBHdxxfLTVSb3fAeukhZTFil3lY7c6obFVIbxEP7YCxIl9jN2m0VOMDz
w/8NQ3oHkspAFbJ8I33am8pJLbYt6raQXLnS24a2X6sCiP4i4lbwKXybRvaUxFiFEwwVmkudh5c6
BfH4djdBSVEL4Cs3v78KFVx9eMJBI50eyuh31FiVpOkOOOf7ZLRFwQNImyZ5Hf9UcRqnfh7PyuqB
O3+1+LxYBARrVavL7844J4ZoLCVXiJwKS8oY8tJ/T94ZsRscVw80rnM5RiLN7AJQZtjmkBrjIU9c
FtP1jF+zS2sI5S3dEtuoOyM+GzMlZ5FwCIDZkX3hjAqiQdBWjrKL8XaUQx1Btc2CiA1fGtn5M6xg
5hx9DkoxU9DQw9CXmBcko2bobTodjBAWr/xjIl3+3t3tdGoh+/mqxrIKd1mP1aVSTdDIEvjZn5F1
K+2CY+ZqAT0S2XIQgcJYeITf/zThmMcnRrC4El72qk3sEZ098egfj8/nMza7KYOWyyQ0qToqx1/i
8xEZJFQQsugg5xyOIsxxFrkbggJ2eDRGfGM+0PnD9DyeZqFABJgfT9nXWQ/EJkQH3uOgbmFEfaPX
5r7kORSMs8XqEAyb44okykursa+f5amahUPGPrgQVkw3ANzHGsnW8bQXSTUOKCEV2jvnRP7rXhhX
SayZD8LwHSwesLOIZwri7D4oZC9soyVUq3yIKf/DGdIF+mKYKVccKzF+V4eCwJP1n4CvJ+G7KR5r
qfAo6sEOUgdtZb1UImMjvgKl0m2nqVyM14BdWpMC8vPy8Ds9dtvdumVJMn78oyye/TRXm0UZzaxY
NDzcJ+sLZUZ5PSbexfOFVuBF9jvYnSBxU10F7e4PQWl5mka63uvKv5Llvq+FrhpmCU8vPCJyK8IP
zn23kTBgwUSay2jowWyDGGvlJW2tivZOBoPo2TYgMLyjuwMgyluY5aJZoYovsNC65LOyVegvSA4i
MloJSrvcpm4WCOwgZ5sZHxVMOLl1MnNkhBqSPuazEWUHN50Q6n5/UiCN4RnEG0V+iC3mZGMMWyRA
QBw6WZyINj1lsmIolsiP1WgfxlkHeYcrI1YPCynQyhiKnC9tPDk38ksbLiCThNJJbPwRqO1NTtQZ
8y90/JlSUaGdfyeWUXT/85VZVN7grr7E584SIDdVhwzlHy5s1bSjhgfGK8V/yRzPUlIosmF7mXbX
uUtyrChq+opBbof2J2a1QWsEgAnmHu+VQtly/EeS6mDKsPHrsJuxAipvo+rIzmiQzh6lUa4aL9w2
J2ZQgMq9XSWrCFfeEge3czeNLghh6pzI1A/2gPDNLwY93uRMFIC7lvQGJlVJX53tkY4UjCDo0fcy
kkNHP27Hl+crteRhPDFiafgMla8HdhsyD1tonD1ozZ/X6xmduQ/QeORll8Wr54erSbNq9p9NXeS+
OkZcStxiw+SUosDbKEYS8qEzhMH6ZNO2Z2pLFBEthHcZaeXkG0BfmCIMFLqi2oMH9BCaGIsIQ0Sb
BVZw4nzE9gY+QUCiKUGBNyaD/+oxNSPvlA9H+6CMAuwmbCqenQ3mH3tIdpAiW6xacirA2wfsO/oJ
GLta7GgQnbvBn1fbowggU46/MkW89oCNn7cFVCZqutt9KuvoeUKGZn7D0pUKGeeYJFWwE4c6TB1d
oyWguE9Ji3ZBNHEKGUkxfON/uA9h2kT/WqVCv5Ty9s4ST9W9WZllp9DXw6IUhoGtrjzsElECmyEV
8oIL/sBJiDUKJcy/mQJmiLeM0uWv7/Szic+QCr44SNAyUZ/lmMGF5wGa1LVmznwgI/vz2QyC7cDc
GQH+k5QSgHiGubjNBb3mY1eKzXXejSmgRr0Hr7bd0PK+ozXZ6AhNY64G/Ah5q5SPq/PxAzD/anDu
4YSLSxua3ffDZ/saSWfBoWxm0zVy1AfWe6QWzQiMTZMD2jrwV364CahTbSadulrb5kukpL3DVK4n
blOnDHQEabwDg0202YDtryB+ywC28Vqmqxyo49U4hDjvoJQ3UWfn9uZHeOaaM1eK47+97AWz1oa+
CejdzjdOgRYLfkuHtuakzfJKvX+1fjvUgQBCcWilr3hdLSYeiJoM2/XJdZNE+LnszsxSL1LTs5RM
EYOTY1/TBMcZyjrd02m32wV37j0R4eOGZ5kdWpIiU52UOcVi51IqJvuGO36p8B1WcHNjKT40dsBa
aJB1Ewo07S+8xJCqce/59SRJpzVgih1Jy9s/bqxQ5dSS9F/M3is/27ROKtL4W8ERSc/C4IoQsgn+
7WzL6YNciUQTyw3MgiKIQP1BiJYnRPANB+zHop8AbmziyOnGTjnTqqhr07yPP5/FyIPCnhHsn/oC
ik77tOALFMvxy1vDLYZSp8VcdvW+9EMka3+P8Mx0oBGuC5mKjS8JEJlu71h3+lH3Py/Tabhzj673
dcdCs6vf9KyBgR7LJoa1orFIzuWUlLpl+oJYSaOkzh/q0w7vBFy4zz6khCgwIb7DQhWIXptN+vbM
H0YfeBR5XVRq5/FoFJ0dcdnD8Ks5q1l3HNNvJ3FG6Bl3LxwPiHJ0XAUAU3Fp6qQ/Fp/UB7IOLy2S
ChV+0GgCVDQa5r7inXNLzZPeCoYMLi2dz46rbN6CWUeBY/mcy4wX9J/iIUCfdUAB3lKc+2v3vowb
r2M6pM8uPrGdyg8ib/zp84EjLpXb2ur7fz9iFa+4zXvMmjgcZkIVzIMMhM9pLN8yDvgEteR4VCrm
weduljats36HlNAwszDkFIh+2rHdgdrct9WiprMbfSKtfJ0YkVCNZstHcoBigA4caEG0AxLLEoIL
77ICm8+7vC9cWp6ygBTW5lzcL8Jq1iU++3/GVcuv0gayPXQ6YQfID+BLMFSrjoS72nTjL+AYMu63
fmR+9HyDSsQSl+Xc8TAoyd3zMDhY8SDSv+nJPnLkp/uie6WBmToeQ12AYi+6e/LNCJWxnrC889CX
3lr9N6O2V0sgxNL8mWV6ww4mx6bG6ExPwHP7nSdORbklYt6LTmRCR21XhBTjiojqYpMG4mahHUj0
u6G31nkzlbqRrm6nd+z8y1N2bvSMpDlm7u5l8+41oj1Ey1QdDiBs4XxV4193wHekX9NDanpG9PIF
bgvZaNQsQVKLJI4hbG7+LwGjaM9ZX2QZ+Yty0uJSOWK4cMwCsjbGGE3wnOyzmgD8zhqCwkScYwSv
0Y9TTzTFBFjV+/w/mYs470Xzgvxp3lpXvnY2C5u0Y7S+GF1NH4UIcfwjKIbeDJ4uB128wSVHPdj5
GTZK3Nkqss4OwOD9laQJ2cyu9nCJ51DuPJ21PmPykOD/JPHu+vZzuSkNlhOnaxlfU0+TfDWrdVmd
KlLuicrOs/tt1Yn2HBqq7eB4K7JghEt0Dm4t0Cfj7Ef4UHXp9TuXqx0yxMrzBe/hXNPLMk4HMeO+
4OLvv2oVnQyx6XUCMgEZ2BKfye+IzMMc1D6fsYx17Z9NVftbUMm4/luN5g0iHVsoBEzQKDKkp+7B
aMtospunGPsc1CSeD0gmX4KFclGtc1BeaCh9YDvJ6+CZedippw1mTL0XPepdDmPNVCNL8TRf79fD
SQv1xSfoGdoX+QzX/9SH1FDFZReplMJ2GT1JsK/8ugg9QmnoMSPV1oBkS5OknLKlIuuGExbzOILy
RGXt9nuS03hRPtFUAzLrTBkW0xabi6vJHgAAa2AueFxINXQZbgCz74PZcBnWKTZX9Y1cz/R0CQM0
hPOH4E/myfVnOFpcLJROrbYgnruKDBG1yb/94pgw1PDaU3DtFRPv34goL/GC2r1zTp8gZSriyRBS
4i5V+u+ZYS88/bBx0vxh3Iw/nlw/3Z+R4Z01sbLZhzsQ6CFVLDoP6g0At8lxoYA5tcz0kWFuuaYm
hM8Sa8SymTaiIHOz5Y9mnQgnajkLilIjVeY/S2nMbnVSv49Xk4XooYCbabz7Pauodwhbvg9VrS6q
hhpHdYx+8pW2atEC1YYv5LUxd6F2rSotxWH7E9owue39Wm6rNQG0I/GRXVUuN0btlzSconAa6waf
44wsb2XedoKsO0Y7AgOGHJtoPrORSjUk9WWLjkPA5FNyu1EhFOTfWmPTpCgAFSEWFY+7FEtRE1H9
iSPWF/pN2ZYpoaw64FcHrk4Novj+1ul/Pygi0r6VVsPTeBcTgwpdR9QLbVsI10+Rd96oMT4GR+j3
OS/P6iW5HcNncU4bzg3lbQSs7J/nym5yOrTfYY/WfjJZMyrmi0OkP1U8QYrcxMsM73pIluRhD8cw
eP+gYK2S9+CW9NbRkLtTp1ABiz4KMNwVvI0I7ag191BimF+P0lVCMGbFHxwx96mYBbL6hSsrtyej
GJeR9//Y6CHj8VwaralXzahYGNzlo+Zp0sRMfWdx4tHzTseGoNDi3ixJgssqEd114XXplhcr2tvK
9D6IaMwUKmGwSjJAfA3O+soYl5niK+xwHfYVAD3583K0ZQx1JIPCDzkuoMMY43uNDYWhuFm4lVPa
ee+L9igHa9A9liuF4OUpS2D2FKSMnp+6WdWCNE4WtkD0drLppJTNhe6hU4SK42flSZd1xhHo1rKI
daARi4SkWUGOYOnmdX9Y3o7kQRBlIH8dzCw8EY4QkW2UXKndsYlTVs1Gwcs0g8jxbgYjTcpwNb/O
fy79BhU42vxct5+7ziJAvsq6Q4srq/HpxbGYYT2G0GoPsEcnQUqI5lOjrrJjWz9OL01wTuMWoqYG
e4TIENd1IMRJ3seyMDvauwjQI/fdD9wHzyf6y7SFVRrTLyBJ6necF5v/GROVDCOMl6G+i4W1reuA
5z3gLFu4rWUWWbUi9FMin2ncin8Z1FXiFINFiYZeSgtlaTkVWfRtWgGeRl5wavoVPfT5UNltsmGe
9+5AFyg3XNGsgJTsBOjWkiStV3hK85WIPx9O7PWvM7WHMBMhX9D99maU7XuFjXl672vq65pIPqO0
oeRwnnIJ5NHxLWq5kW7A03oaARQrVUKAZi2TbAJ8edUdwuddDTYQNjYNx1rqbH0RpZMuwKz86M5T
4Vm6gih1u0sIoDLtnHJNvzpcHU81kXLzn2lz6WnsF5BPlB0MEMkCl1NnpR+Uw4kx+DJJ8anm7cTQ
GmZ98IEQc/tlOvmCAzDTN/8wiAbQBkRJR6OY/PN+J6UUDysUbxeVsB/ePjLc7FqIvfKdA/EMGELE
SCYmXk/TZFKGLZA2b9IirUHVVyfppg2TNewneo8Bms9BXLEMJ+/n9Xnu1afX2fafNPftiOe1EWa8
mlmVyA0lJz8JYe9Vx5Be0EwSrL3LOtnE9XWNJZWFXs1YaQDj/8NqU2GbKsTLIOO/cCYH8rxGOxZO
YlAFbpY/63uGK7/7lHE1SQdYtLDhYUGiuqF/XEpal3yj4S5ogSSkFmF/3J4ZugdafxNZOzUhZNfu
k1FUkwItOfkTU+wu1k1DglTnLeoIG142JX14mXIsyDjh5YfSsL3fNbWfJO7bzDxikj21WtY18cIg
Kv6Xtw+FWi2rmqtsHLcTO7fbG9Gx7qzqqr+IOWtCI5ocKb10DmCKBdpTTMuobg3IWFgmzWBuKpSS
nobWH5fczrHbJGni8QyDHOl+/NTHRaPyITvlgbOVgJURixZBsQdjaqUItw5byWQyAy4/znWmGZeX
Q4Qu53gATINpUH4LYgAqwNRGiTF9JMPlo8i0juNHippyXPVGCADEiVzE+/vBhjUBpKFyLBDL5cuY
hflUw9wCm2upD9UHxw9Xh6g7Kp84yzN+CH1lRmt6S9l07tMilTRizbWzJ/q9JwIKzmvzhknJRJ3t
7M2b4iwprMI+fFrkSpcw1p4ythjap3dtUNFoOn70waiFlJXr995sWoBwpEuJRtwlYzgqVppH/gKr
/Z+9jT5LBIbiFS0HVxVMtFi8dzmtK1pqmtTFmynL/8KadNnt14ux5fgBZdUFMmP6/2P/K1lF7uGS
n5QE86WYKg0wKkQeABcDljrThD/TBjDr1RzH4nVUw6u3eomTkJO+cLswEzJxOJYUobC5LI0sftJW
JqT1zZbBz4vRFua0beoJ4sz9qtLwurM9w/LsRHw2rmThL7p4gIXzEraThMPeHtxs5EO7WejUu7M8
bzYuhbeXwjHhFNYJmx+Jk/V2Wbq0pzWGZa3FFnmzDk2Ec/qcn7Tsu0u3JzUO8kUlJTmlkfTSS90H
Au3fMQ/L4IZkFITkCILWWT2wd+/WQoBj717oPINz9yg5z0QWEun6B5Bd0+oS+XQ9HZP54iKge0T3
UB98pn2/OBz9j4OxSnscxhDaxJAzaDpbwa6471v3AtjiqAQ8tWAz2b4lkvJEx2cc8UyjSFCCCi8s
p9kBvuygMF9t/hh+vjMz8h9g7Jr5SUDDwt8VTpTZqYI7R4iB+SsErKCdjaBuCNnCyzZq42hU4Myj
pLbA52ActC5NpONkezO4H6jVd6To6S2vvckZ+3wBUlwHqAt8qqfwpXoNP4fJTy+k1R4mv7LVlnLe
Sb8EXu7aWexp9TyUYmFV62dFSO9RxdL0t/cx+GKU71Hjywas6dBrRpQ3WdWHssNOAXLTY/Gyb8ea
fobBVcx/Mlp8rWIBBPZbQnJx4r9TD+G62H9+tNbLCpn/CLkqUb6RY+c7eB/VWj6Q9dYNbTRYQoaE
NNeIQb9cg3P47OMJfvz53vqFi6cwL/iBdoDePBYCQERoFBsOJUP+h9ZDsWIiqERBpIgeNGEThEgB
WKs66ajGuU30SomYeLgXSP1I48cFzl+kU3FvA2/pIpIHKBLDgiAnYL5vct6GfuWkZJ4jMgzWPLA/
iUrQbr3QNKwgtKrkrBIAMv0wWBQMd8yBkgj/yS4lr+noiTOLLpHT+VKbI3K/QuBswI/iC7xrCYKb
jUStiOP3CvGeIRucDR2UKW2IhQizETEztQZ84hYsrMNyK3+dKuIqduoAZXjAFjYr6zwjUnBTYAzZ
hrNrr00G46DdTJOgfIgGrFVMUzXIvbT7suJrBZ2u5eEmAC9ZB1Agg7iy4tZ2WKlKHdZAf15Ysnyj
bZiV1NzLSV23N4HyiQBvoR/jYQ8ni05zMNI1Q4MZGcno0Vti/UlgBPlBVZ9dVig8P8MqKlrS+iPs
aXqmlqNVqsK9J/Khy0+3caMml5M1Gbbf9NE0Cs7w7O/PkQ1Byv3DwIDSwTxY32xRMyXoN143uGw8
5qJksryIvoQfZj1D6e/SmSPuAvOfjJ689Vt7EMkUFUhWgKR3CmreYX+cOqIgritv5DhdXStN6oSA
uRYSg0fmyR81FRzQOMiTW5DXv5lglnZcxFFV8bUqi7sXuV43//2Vcfwhhgl1sozK4G5BLRvRupz5
DMDGoz/joskD65jy4NCDaHRq5tb+QO4s5VNbh3KMtPGofN+CBqfCe10M5TRhtnH05YnPFV2UkCqy
kaCFAIxznhGEuGpKb4gb3VmppVm9Gma0UlXvYUugehP6TgQijFPTwIF43h1IC3FpU62e4CBneBan
Vpt/w/sxbXHPz8DGrAEmN1u8o4Yx4/u1uEKg6LXz6C3jFxVvxtKSRxI08pmR3UBbruMy6hN4sH7/
1EFZJ2jRURJ15be+r54jvnTUVLqk0q3rCDNUEw8NNip4f0OG1QFOn3A3V7n1K5a4erUXm5wwMX9l
XzYjYWytF2w8YODvb7IPPmklCaLK7g1L8S6KulEg1agKGdmQ5G+Xtj5H3BkEqsLH9ZbNxrj2LJzW
1bsxPJpdl3UaMcaNpDVbJaBGIvjouNFaFaf9EXKserhlFnx7dlmEhQCeI/CW7C1k5b3pcNL7wBpX
Mv4rgq0XZL/7eDQ+G6Zl2iohk+Ed+v2UNA6wYOHOmdzfpjikFKY+EweH8G8hrPLA1Qjs1xkFlxIY
JsDdNCNLbH0vPHW8i39D0iizVnLA5T3YU3h7Qj/VW8Iean4duTW/S5HyjPtPIhK5ExSK6NsuuQqX
TJWATO/JdVWV9+59DAzBmPR0AHjR3PNcacHh/vsOSxta7QIyJKPHmUIMja//SLFoEBeDZ3KKK4w9
u8xZCl4kQEySrnFmlfCsoYllePnFjI3Nb1X3KkcY+KjfCAYm9xCzHQlI9OgWexyxRC9KL6W9JJ8n
ROI2b2urSUjpxuekjlDSJmpyqZcNQO12yGmvBbs9OBOjWxCi4UKzBBlleqKaqqJnqVKuCJjnvdOA
EIcMQ7I+FUl+9f44aKV8R8fZm6IyajqPsebXJ2KNvfsOSSeP+3ICDUpggQq+cnnMFrlJDAiV/+C9
UJlNOe7wwZIofKN2qIBYgrX3rlPvbs7pu4xyQiwsRWh0fmge7bxiJ5QmuHPYX4AIqLbugf1cwx8z
U0UB5XVWVKa/991+k2mHMxPmr3UfYKCBdPaLYlvfT3B03l45vWDYDF/mkkafz3TbI2Qu1vS2GUXD
lnqjGrInLqI5SPfSFqo+Nmo3GZxQr44yQrA/7mijdHXzRDcz9+SkL0oOfu5FUDKAqZYvESmhBCgJ
Jdr85rHPdlpkcGVH9GuTQYP7sN3p3SeBWdW7qiftF9gKVHambAUmMsQamB7mfO0rGdPt4tps3Vzu
TKZD5wJ0QPezl50K+ry5wV394D2OY1zUN/VTrtkl3ZsBeod3ZFhpxe45KIatu1Y05J150thRymWB
X5k1WWgUm4gvecvLPdJVXMi/mkZk3uP1lNTk63I+fBA/VVXZXtgcRTYtc7IhG3H+V0WKeOHXBb+r
eVIaPsldl2vDmFZ6h2izR2HH/LxOQ7x3EeTJ3UXYlpY9fNz2zcByjLxbaLAynMcqwj8YvGIVF+hy
BDTBHlTU8V1Ht0pskcl1NOIMSQ4Db6zbDgS1FLzLyV6LQ5fADdg0j6AnUKkiYSBy4eikIqevl7Nw
Ps+aXPer3okgwqWavLHXoNkTstSeoaiYlSBtXZFKO3H2R8D2WlIl6W7SBywiQKq4dCbwAN6xmgdh
JJMAL8hg131jGaJfysK169rB+cUnm+1ny1M923p3YiYNU1mM9QSNEIwTk8keExq0sImNduCAXT7r
MVTsBErDTOp4EQEVm5VfZ731EbnFECl+kxIPEFFCW7NHc5UbMzhnsKrQS07dGWR/mhR8eyfHQObg
HtfwPcgBkqDcMasvqDZG+WrgYXJwFDUZV/bda9YhPB9c8XMerrJ8hJS48loYoNYl1Cpk3PvXUdyH
lZd05Ew28VHXgY0nkLzyW5LgYcPXsckQlgsRgkGadBdizYuWLw+kGiPC9zyxFEWtzYMU/pfrV/9s
iK9AjJdZ6kjQWauKgtVuZQDsjdYFhMc3Mzb940TbHPF+qB1CZmQSn5AVptjZofc5tiWFVqaLsMOJ
cxMJkAeeAv7VzzXAt8y5eX+oxBv9ykGnXD8LvVVwZmt4kbhDDp80BIB+tzk2Rl+wevU3bC7CNi1u
FVvm4PwP19oIUjqD+z7W08gycMK9hUoaj32n59qLzIfbQnL+LVZLAGhkuzwlfHhcR901qS0nT2WX
On0cTTIPlqtLRc4vM+Bjy/uEk1vo6leZeV1w4N9fb02clDHHS3s3KOOO6vUuLTXqOcYFYeuQdAxe
im2c08LdyPb4NCc+LiAnPyZ1AIJxB2QsyU1mi020W64ypEsFoG1yMhOInabJBBcmwmEhVRc5dNvJ
/IMcCe8Ivspys8cFuGK8g8lrJDRX+0AwGUfJyJiqpXlm514PQNNc9sO6At/VWxYWpDI1Q5et1Wza
nUDyaMtXbQmy5Tmfvhd7idHUIRR5Kgjp+bgYSFZAeOJQD8lVQv8OHWXjDAwokp0sgPySzSXr+YFk
7dgJEIDa5XujqFXrWbG/NthOJmqD1BxZV+tHNzS4WWXFeSoe/0fp7R8jbMZbrcGoRbZafEhkqg8O
sGOc3slcC52lle0rKtr4FC+it1NO1+Ysi/kTbe0cE/zzHn64pbNzO0S+WB+0vkteUzs7RLHgzWGf
W3XhsEXfCjv+7rUlojAmX8o189v17lyxo/hZxwa0ilyjVZqkMcvq/Y0hlfrs9W9/Q7jZPQUlXlre
4ixt/H2SYhJrKJyLNx6nq2Up2vpzu7aGsWkuP9Vz8B7lASVY1FS3NbXCaSUKPakBS+kKaSbE6w7O
2GzLNxETxDhqX1m9QGk1y8kjQ40u2wfXl1NNzcZdvrwDjiBxow4GhGW1/kA/Xw7W75Zui4tz6hnL
bJbWsiiMs/DJ7Efk58bkCo41PKsMJvnCu97JxYdwVvvBVfsK595ngzkDbAp2SRl6TwLvUknQuwHa
erTr1ZNz8/B9vJZKz+qS70vh58CMUXLkH0+q0gaWByhkoItkHT0P9+LYNaSAV2STCqLFk3l06uHb
Lw+IZJ7qMrp3acuX56pYJIYjpo0k+17HYEIMm7D+4t9OC1WDMAezvCNfpknxLJiKU5BD2R2dxMpJ
UvAPezmilG7xhmyjhwg+mj9v9G5hzrmL8hjTgzqrgHsqEnmYE5ZR1t1XN4Slmj2AMLfdl35NwiHv
epjrVBtsE3mPTtvb/8zPk2TZxz/7AeGipcHrR5T1q0ECcdrKkwViJJSKQy2UQGjHRfP9YkeCPAhl
Kha9MuQFidPfTsyWHjbrddKpe/E42WRi/57o3HIYPXIRHskvKwXzX9izGQHcLGTj/7MdndzXqqma
RPZLbd5P67oLnikLQSqMUjRVPlwj9ilx084qelcjhJhC0Gn+fOp5YymWwBxVFR5iiMDh8wmUPQzt
KIAION2bDte3ZGV9IvrYoJnoLjd/5bvWcRwzv3brgjCKWo36gDnsWoldgJO9zr3W+DbEl0xN3eDZ
N9Dhrl0Yng/olLiXH8RWJBi6uTYcXcekSP0jic4ocQbW64cQffnhmWMdCY2MY7PbcsAaDsQZlxlt
RPXW/Du64MfkMzLyRNBz9Sow7jyJnlHNFaKsG8T5U4kKgONeQOdTfw2x2MNzFKYuWpjQViApXDJ2
OTSt/zcOMGTBbS3aYtlSaLDgBIhpr0JkMzO1tudeqsUHNZDrmiOe8rmVUvL3zkPwT0tgfX/TAF1d
t40hVZKmopi12xgvd4JUCRiO4jA4X1DudFkI8sXXj5Woar8g3r8vSfWWqFgAiTHrREIRscv2JZZ2
4nl3oeVFGL6tXO1ElBrCqFs9SldsvwX5nqFtwOHhduwZGdy5wYM7ksOEwEWNVOUEuHaqwgum/79/
VZTZZ2OWzrtdetODqk/KeTc1goHmk3erjU+cualVtndfYoQfubXMYCOWPAOZgzA7MK4bA0OK7ser
rr+r3DRWiRF8ESnYAFHDIiFgGtnHpiKQyYNoP5kbuqo2JMl68GPVwrGA+xvKJ4pqDwTAx1TiMwBp
1TUd+IGHKw0gq9cerIg5uKzQImsoR4cFuBSDaI/hztCxTEEd1s88VA9cTOZqfDCgGA7aZQBwWu7Y
LgPknJ06e9NKAwQaYTeKGVbGVM5HrveB1eDCBfl6Uy2OxjTbQNOpvDsPJtXy0wtP5ZvzdrN0dcMo
lPsmKYyU1O7gMbMahW8pmDWveqM5SRIKGYwt5qIfDb8fgqUh7nUYLqTnHBil3bdndA/D4L+Pz33i
8BvEG4D8j8Uw850RgrdfjKNYwj1X9TVLyWFOKWRlXAMot1ya/k26lmr8dLRqBI4KSzUGoDYQKuxf
x9OtpkdBefFDnu88Z1Ra3KjskyQqkga/c2Eu2Dfl4kZlEzz67HBYyzYQmQ1RKqrzG5wxFv1XvCpu
xQ0Jxwr2l+Bu8IBIfZAzmsMetDJYA/VDQ4/tQURXT4unHGPtvDLIIu56osJ7MwtMxmH8jaxVbbfB
51KiTUHdNSJH2Ige2YUY1CRI1STwldpAWRPbPW7qcBA6MuIBRB2yydB+MdCr5/gYp1/Up9YBIwWW
EStc3UkFIwAFIW/7aqMCDT59wsUpcNrTjuy3kpdBVnhHo3c4/mqPRcsKXoJv73wORIg9N48UNh1B
/CXLeTOFLhYqI1WDuZ6Ry+WKfMlcOo7dfL7SJlxcLfhGw6JpbQXGRDieHzZDyes14rime3L6GvoS
CLMMRS2rDhLwj5trYxqP20YepxUUDhxLkH10i8bLV4wVhJlsKDzd3895kcPlnCtOmg68kAvXrxOB
GzgNz7zKLQoVoiYTNqVsypMz86reLhI+iakzmf3/dR3Fy9+yhfkDYDz0o1WJVGg9UU+9erkd3rtI
YHY1gst88H8KkyXcXH5xkIKfBzXELRi00Ozwy1aukAoxIQzI7XId9ONCDhsodr57zx2Xh47TrNYY
2lNIcNMGcwYqz6ercqJvu/nVu6KMPTyPDO0ed08qtjOzUrqmvVDls/BBituDPmU4q8ZoBPzg5zK0
GiEBr+dkCZEqIF95zVZbODdjMU6dtqV4QizTKBptGjHaejOL9wBY2R8h1QrA0Q1eRezyXOMtJmok
P6n1nalBpJHolNHdkHwAcwIXQBrS2wsAiYK4LqESKxPmX2Z7xZa/YQJqTmn4hpXai9eRbklEyot9
oJUcWItGLrcb/OJ+Nxzr1hin5Wtb5Y04D94wLke3H8PhtS4OjIdPXsCqA1EA6MYW3lancX6yLGpE
kNSLmmso147RbuxjdFTmX7cB6WZFA7RV97nVMlspLxWDc3u9nQpvNY5VwF2HJ6Z4376aRo654q/A
GFpI3TWaPPMJZiUyl/CPqAwmIpJ8hm32gEMFSPCXH/rhEQ4Vr3YZxSKoKv4pOjTZcezU1rmU5hgJ
QPewRZeDOZfWM7YQUDK3vYdWOjSMxdwuqteMO7n6VnlchUbMBsoHOWMEBBoP3Kf/K+3VjQ5qc/J3
Q6v3IIPf8Mklpctlxmio0CbpVyvmytL9bc1KaDT6sbf2VXbyYVihP4PC2czL7346ViJ7VQANlosZ
IPEIelZEuQnB6TWbspSAFYnmi+7SWLy90FBlWWXDNh1yDPqVEyJARYkwv9KQgkjtlUcTO0HyHhbD
6Ynbuel7+YesS1k/xjPvS3txPG0vPI4ykTdjkkCEwOlEPF5qTIfYsM3Lp6sGy/U+xMjXzoxRMYOF
uY7w3dKuDvi2iG0gNTBBUIJaosjPf+QH/LzPI7uduCqZTxDvcPQbK2bsJPJs5E8on4xcG8FRNlA1
Yo/+D4sW95wCnQIyj/oMMTBX71VvkVBP9R6c0Vh3wJWzbvhG0s7d69nQjCBVM1mvYqI0nWH4Ph1y
gva9f+WutRmPvdsFgevR1v6PvubkZSwyCCx24Vv4r5xkNWnB+yGM2Jp/rTGOjxneBXVXr/TBGYNp
m3P0c6pAbY+0+x81U+hrOAtO6m5OqwlOw1zTMBcwqo1EMgRajTCYS9w9LNwUPPz2Do6fqpQYnB2u
fv5sZataFbAgJTid01qZZbZZeEG2mDbvI1KwpA0R9fABZ7OAk4J6mZgYKdpDgUwAqMBTjU/IFjd1
FzswyMKUaMGQ9mEHuLqPEYzWbJ/mCyoHRn/DdZn/eBBhDSCSXb4RfvtOAstyq065TIEZyfBzFWyV
VyXbfW/FxK9dB8J9aTBNAUoFTA/3TVbWQwZewUBheOC+7+Xpt1zkX2hnTuFDx7oeODjajxIHuraL
rSrMsiVnPP7ooQ0Tmrs9eYxbntWm/Gc7/D0/CC5w7g+/680yGTrGI4CkSPWdFOaMqVZUfKsW3Kk0
2muJ0PmjSNUiOuYk8SV0iCBV0iA6vX9PrmoX6oVy8sfKJ7nZ7RGmwoqjv8nm9DD/ZkFgFaw+mGCq
csWGobvTUnJDwR97plT4/9nDyrqvCWWWfD2q0cQB+8QmveA/MhSy8ZBFccFB9o1yBqO2G33ZhGss
0h8SM6yZs2w7azNVDJ9C+D/iP6P17MnC/RKxWjRPjLHxjtcdZ5Diq4FeSezSVOD23xD3uwODbn02
XtyhdCPHTOMfYr/gcA8vPSAPb5LWd8ylZvVcJ0qk5HoLR6oWoAGaqAwQCRE0WJoffPGGFqsrhW/V
EC7vHRxQ3clzGDCiC/x0VADS8+zapbSIfvp0PzsaL4MFfbvIIYOcEv8mZDAuhFoS4rSt8BHUJbSg
czbl4SH5TuvsKVJM6ShfbTndv8zTkWgfvUQmlB0M9DCN6HZVXpNXVPsmIod3bQEOw5AVdv0uWGQq
Mk5J1CRBnyxlcjwpSh1ITE4mAeSnFSPwmnpQE3PNlOJcSJS+9t8dUQPvNZjXNY6177f/ohN7T+th
JvSUhodEJKwQcFBkxp8iqgt5K/bU5Yuqw4Xr7AxnLq1lwxDqe3fiyWNa71ceyXvUzS5+FNTsb/uL
yC31ruxSMjaCM4ZaDnZORVtQvJJZDpbtvSqHPvcz2buC4gZssesEVlueGgvyJbXS8CptYK3wu3eR
ONk8UuZxM1LCRCD5j8yB20tzxwOZYBbuP1m9nMT59WmFXIwO3+10U7U4vF2n5AdgSocBp4gFn7ok
IY3jIBcgaHAwlCESx8/fMr6Noqy/08Pt49O9ukyKwS6lvvkIlI1fJGnNa/3ToGW4BvG1T47MLv/w
rO5tIuT8Xd4xD00xHYxDSskIhL4H9oy3h0Xxpit5N0XS4Ts+hq8Ema+vRSzOrDct278dOJ3Tvk/0
fZLyhhDa/ooI59nVFov1qivlmHn3q7ff/AcG14PdYLriAddEv/Kb/7veWhdBzJjg++slm+dcqDs0
UoGUJUVBpG8ueamSsZwiycG8IVYINhm0LvohxnjO6loH1Ajw+XiggB1kuPhDsQ7DZdJ6yVWy4Pow
eTbUgnsntpGnhy1p+uzYkV/yav6PiNCNSY9Kp/5mAWpDoPFILVZe6Pln5bmASBK5WLwFmCRXaNNz
igRovRaXkiQbbzEi93K13J8WTOFIqVHlbnMxfffKvLY4QRZeMOVuT4aLhghJ6iEr/kWLeNpLuXJW
bXjmpMWau2ze4lxe3dgAGfu4bt942M+VHnaHGumjEbVB2EAgEbRb0BNpmVH+qeFgrRbFtWtO9Gis
UgwIpMxDzQCdrQPsxbECn4EdjU3ph7T0tR2SsxdHeIZRA2SQR59oRy/veSfTyRn1CGBrYPnVWhTg
JGFAGtUuRtvzmYE6HWehxgMtR8wD5I5GbeeP6NCjyZWDXM1y5DhQhSrJBkUVsYsglhJ9dFGQHVaO
IXXqMkbHrYmTCGX0lxHPbCqYoeYLeyLXc856RuxCUBv9MXemlLueamLO1FvlR8kUfFfS6efDQwGm
nRqTXstloQtijIUHbfBnaka0iJ3jvSYe6/pKfIKScepYvmSNQr2iW7d/VssZXcpHa01lScBESc3a
NxLBBOWCkopNAfGRGjA5FdlZt3JvYy4ES9ZpTKW5bjzZvShG+rl1dymkyu0t9K9/WOrLQZ/MITNA
uc6S91GM8aQmAqMjIhstHiEYdsgIYIIfe3HWvQkdKYWXqWda5s69wtccprTb1gyA6ItZE+guBcGM
+F2C1CLkDVw6fIGDz3Y6+0niQS0NYaByR7cl/iupfNdF7wAGc8BqfBc+6QK/nB0mVXvCQ5RcbES7
l1mERd/ezdnwHyeepUK5+nlKVKYAf4pRW64BqYFLns+13AdcBcsMgPCtBMzSt4zbY4PzyRXMu0jy
tEhENt7dOGr/DMeXLLtZ6WoO8FhR5Aywn9vgFq3qg3rZlxxNCOFAVfaYWRyTUURQdmtWpiljlRX6
QEuCoeXy811lJp1mDQdJF9Yc1LHyDIkOD4HlpcLin8S38nqef3tK284t5mdNwroPESANAv5OaaZb
ETd8Xmfz63jA78FLEIa+zQf2tP9EbERVo01gJm/MssoeKTEsRGVDotm3HDVCFN4soGGEFdKzDvH5
G+q6x4o6Aurr0siG1npYlYURDApee/HMBxyqbNMd/vAN625gIG92lS4XdJjHOZA6bfjXqXWbYnj8
vEJavXa2YDuzASjgDiuo74IO/Z8C7372YQbjHkkIzyDNhRFFeW45s5AcjbXXb0wA6UKovoe/VkKb
ZbpL+RMPkNgG8t3IVGZRocoxNW8n+fwx9BhxelP+RR6cjGn+doR5KNKXzImPJ9oMKNQ6aE0Z+YXd
Acz2vTYSEUgERBDDUhUYMZrx+kTDzt3mKliC5L9Q9D8uvG1jDTfX4PZ3k89G11PX412kDWMJ7riM
J1N3J4bYSqyt9yZA6e4uSCxPpfbozYwyBRHvs6+FF/Dlpzg1Yi3yM9MaCsVRvHTSENdps4Pjj90r
cSjB4HLS/JdDjAii99PkT6ejMJ8CrPe0HgiG9RWjuoGdmFv5HEk4npkg+LqYzYhXjFTh4lPjx+62
AwydEiv3sX0dcPhHPNob1fOR3MEMVi4Myi6o9k9Qso4mUQH36OPc0zivgFFx2ukO8V1NDHJ9bc3V
Ef7m29w1Wm06zWcQn35E0EMEzjrX2e2Pu2jtGLmbGH9ewP6fTks0zN0fyWLT57LKGepUHedRHXXU
9zMboYDT7d3v6C+P50bOyJBQvgG7usO5J8GxSD7So/Rh5EDzLy7ATWHrIpxiWf0H9sGIigFE/n5l
7FLPfz60ZYDESJ+iHBJRmYxJRev2tKNEzR8AnTJsRDo7klzxNrmJ1Vgs19voZPt6aLU5WNUtqPCE
ax6otkMrd+tHFFIEGT4nIToXU9aAnZAUJLSc+Z1jVnqkAyfm7CV+nuLVjodo7tsIptQQ1WDDBvE8
4y1pIZvQMZG0kz9tURejs+g1bnSKaDb1UWlvRxtcmxR+Aw5+FH6shF65r8wx8aZ7UVy4vUMLE/Dd
+laKU/Wp6aaEKWKBD5T8IdTP/p78UqiqBe1LUHDuJAvbiSaFsG/dtTWgTowvxxk6d79EMASzjh8y
yIb5CnhvLvggGXoRjE6eA7pWMLzSARZBrWvxfGZ0MoTkRxKK+wb7Y1Ffyuz3SwZaufwMZjsirg9v
bqPXKib2EFHeeCCjZPZTjLSoqlqJwRt+jmYvLIspwf7vXZCvYN2gtkgkgDuS0F0elPqL039IplQj
TdTUW2Q2Se02DtpJfBr/LGTgR1zX8AEwFNScJxNdoWvMl2FEEzD/LYTBaS3OqCcWZq1Q9q+Ka12c
0E05KHHo+Ygy5xN5DTIUaFbaX8ierb3uj3n6AuNwFFaoINqOBBwosq8ONRcRikwwJ6Rd0y+g48GC
vOz/KpmEgfgNFr+aE4lt5sqGiCFu2AgTVRoBEv98BZd+wJCkUBBn/Xl6fqsskNVyKexuJn15jkeg
ROJd6PN8QnICcvmXLzHLPale9dUZTsiG0U0YxspOUImr0U1ARPtVN3MvnvT7Xarb1koAu9GIM/eL
Ct5tnjlms0hxVuYsKMgHpfZqaXATrmHnwMQZ+nt3d6OC44B8/9p0KYIbvVYdgnQIn9Czsi9YfHhI
VCfcqSbTcmuHMyy75wwS1Prv4u9Sm1+V0Xuc8OsvCAjmOaq3TUAYiPG3OeMVTkxk2HZIzMHzQuHa
XXIm/3+x9Z2DR06PUd1ScUr+rNvu2c7QUX5qY2hKqif1kTcXUneiasoiPsAoRhD30W58zNpNKrMX
A0mHf6SvL8LYC+lmBUhSHPNPNsbcBGZukgXIURKXRce+x1v/jh0EsHPObzgCKr/zVbJhnfiG3Pe8
DAjOwnK/8Ilr3CiKqpvftweHdW2nGgxCCQ1cFhZZNGSGj1uok9rwrlgaERm+nrnzrlVPA+jY3FpE
hUivCF7vQ9QOTqGxH8S2DKRbLT69W63j29G8Jaq3f/g9JYJFdY13oyTD881gMNYLw7YuD4RTWcPL
mT9BzZVqI1Tr38EjfQ0wsFA59IBUPM48ibFsaLk5bJIe+aw03NhdCRS/bEUqPgxlXrWEk0bmaUuf
E3z2paKbPTBCAcufIAgNoMNYezn/35D68g2K8a6Oi8ywJXa0I8T3bk2e2Ej8k7ISLDkWJlPh2b3X
fIAjeVqvU2p6v2oqbVMrQtGsmuE1k+ovX/x/4IR15fPAFZhru4TaWsvnM4EPClCFjAgTe2NZHc3w
F7oJ61k+T+lVMugW5XU9WhfutqvnshzDvTVS0qy+P4BlObAGzhkfgBnCjx1XNeDotZPa97aeqfXE
DwLUypNrDY3fgX2hZvu1aP7yS8n63MVtNApmdX3Akh5mV21TznLq/MMWgVnyIzwZazGnjRpTNlyx
yzQh4IJHzhgpAgpyxlMxWNVYfTCnRLrV0aLoWDElfFBh/q29lZ9YZZcJKNR7wNkhd/YQXAQ9j6Fh
dpMDtKK9xk1tdMitUTX4OSPrg/qOcyyIw9zq4mjCK43Gwuoaohzi+Zz+y8SmYH/CyYVny4+8UKyq
JKz/dUVBth8fjeIftH/49Em2E7T5mJeDTGC2SOPMySQINb1m0n0DTSBem8sCdFeO/QooSLFNDZOc
y8511A51j+pu8VGkjMq0WCKDlZtIbZc2sHjhkUKxa0YLrFy9itmtkrV8nIc8T62picWCGzCi9RM5
4h++dWsRFFDktAsxLJbz0QkZ9OxWlHNNgfu8MKvjqC9EuIVxQx9ArwcTE7y6z4vXbi2yHJYQvgH7
misFQjLxWVamt5U1pWtY+2iNL120w5zLcIBM/R1Arvxc/kKjWUtw5z9o3s1iUgMcxrQS9zLkXAJy
7zAhEStziuMKWcc9LW5eU/h+8F+YL3XOydIok2fkamTdq/g+bkLhPDkgAtsVRTkt/cYx46JYBAlw
iIjkxk67UKcJxvPnCc5fKX3zzZV+0nA5QKkk8XbfiRXhJIidGazDccVtFdrryQdmlViJMtnq+xe2
XmN9Vn8jBqO4w/pqNX89bu6SxVC2kC/rUCsKD/ulwBH9dHFhjLKDaXJq1YbjB0/YgJiEjhQr+UZI
29KZdsX9MRod9ZmI1sXbCpnj3l15IBLqsuJ98fjvJkjlNovFI/gSyqqYaP4CIsINDnOyJVRPHW0N
Bp0J7IK0cgfEIxgeZu0iTQDbkFT94u4AS/08k1ZWm0faGCnilDiG9XdkK3oD0CS62k96zdBty7RF
OHY0z52ylRoXPMVl81Eko/AUq+C8cTMrheBEsaA5AWxEsO6FxuuJuivUalVyL8Ke06sppG6kkbg+
6nogbc0KtpWJt9biTHzwR9xJyu1pQr7h3MbT7Rhw3RUWc3AOuoWIt17779amgvpnSBUa117X7POM
oMzZsr78en8w2CKSL2+IdDqJAkaxGjd8Ck+JsHL9Tl6tmp5SWBElCHe48l3QHs9Z+xyTeiARvpE6
T8jkhhqIG8aOBd3KaFG+fd91fwwF3lCs2XTgRFA+m/280lG0qKR3jITr4lVZQQ9nhx8JniRhl/Ff
FY6i819rA3Lu96i0kqr4q7Yrjkf7b9s0PecLS/Zsc27YVLjBj72kVja8u5ibuCOYHQhk16lpAjmP
O05mr6JdRj70xi0cCD0TBQTIStWm6KRQYXPppY8f9Vr+AGYLBzXC/BiVi4IQWPq1kXE9c12u/umL
1Js9TdVYiPd7uqGm5Erpeg1YmkezqS3mFl9Dl+Al8I5H6wxfb8BpxWxwr3C4TUSkNzMv6sJE6t0x
3ZxgwCSd2HRWCSPZzFdqfLoPnlrRiGPspHNgYk9vULXGCabYF918/7QyA3lZvfuuRBYr/HvIpr5P
/cGVF2g6BjXBng9TBB5GH5p+IlMeoSvYV8FS4gArUazuqnT0xNFuhA6bYqOlGaG6nkb/PPgSrIzP
tmBbb5n1/hciHhA3EHZYez8ipaPeUOpQcjbSoMybHVf/4S6oqwY4vQwacXYzZgXkqgDE+ielkyu7
LUQFyl2ljaBtZ2jjKghEo9UTNN5ivch6JUSE86B5xOL6Z/IZlTDRj7Px72fNPF2bGrURTXhWQdEZ
ssGyZYXVvge9cbpF1xvsssP1WFAxji1USQQK99McMrjC+FiNcBdVwRDT17HXcczcX5tFyUo3tQNj
77ZPicrPxqkb3fRCiGFViG5zBofyhbYA2Lz+FagKNn2prcNthsx3qmTCkkoMVcQWqvPzmLDWY4uc
+6j8N8Uoo2Mt35/xrza5s2injboe0dDOkIwpBTx7j7jHqme4URE3zSx/EtdAd36MDWYhPSZeVV2G
HJ/liRXgqs11JdVpS6WCHcdYFPHU6h4KJ8/7WysXOEFX9qfY+GKW3xG6/Le3D8UUx/WHA6Ac51d3
Ga5aK7pqFgMnwgvE5cgX+JyAMxOnw49zHcmMLfPGTB57piHtDqBSlXci5JkM1GkUhFAN5v+fazQM
c5jHMPehyj+Hx8un4X7izE/SXkkw8sOdXMGE1zfVTfaHpv3RbZi5/Vm8qp/OlXOWQ9S1zvfdb0RV
Y6R2/zOixJiabjrp+0M2x00sYJyU4TjbmW82poK9Buntj10sGkhqcPkiVUaAHYE5deQSLEsqhIN5
XzjyYhMIagUbz1t90NmdpEPCyaZX6PS0zt7Q28uYewZ4wuAY/8caPCDw4DXve7OdHyEOGSbm0zAt
JGevBRYvOYAuZbgC+RUbz7DHgopogQL8fZvbFU7H1KKRElxpba13lM0/DZhGRbsXOp0HgweO5zDA
U9jOnNpE9O5WxcGDSE1a0ZU8qzEFJga7HxtnMVIF2+TZog6Ts1lVKmrEgSmY6vvWSWGwNV79Remv
nHaEVRgHHanFBDmr37mXXqUBOkt5sHGigsvvy8DjD8yNehb9ARx1kDR1OIgUfCf+iZc8gpTqR6Kx
VxVw5NSOO1rlBM4JrnTCF+SMUAH6howIja2yVQQJTClSCidof4xmVGO/OoEOxWx5vxR7nB+Q0BU/
I5RcjGZFcUwkFiS11pgWABonuryg7LwrTRRwxrwIt9IR7SgInUnSZGqXVI3towUY7RokAs+lfKiF
j3YkyqBG0FT0tTWNLrOemAxzPJGeiDAQYdaXOtClhu6oaLOSRt16RxEK4qmNgPNDkvEMvWEHjraj
qAaBcmRogzbY8lnHVh2JqwR+W0GjLgCqX56z03fyft+/ub6u9uFQPWwDtN37EzF+vwf5h8pWwM7J
i86Ym6b7LwmjtZQUDkB5U8fwDPyYSIoiZ6e0GbKpUutjsKDxR75YqptD0eo0bvQCGtHqCBU15i14
dTObVnFqOL1ZeLaUM/W3HczctfzikH37sWSZ6aCsXgbuY2r4nMemSUbdDAzxKsH6VxL7csUx5s1i
gTJzinsr3q07rjACuJ9LfN3OYfzfxQ6mj0g1fgtzqcePF3QywAruB30c0F2Mje0vj4ake6A4yqd6
XSF0Y/jrL/lX0oR4nPOIaurdlkoG2+ecwKrkj63T6eEORJ4O3C9QVOVPDqo05xO8mXTZsrNT2BXg
7B8Fyotgpt3reTYJ38xPW0LrQHMBWHdmtG8K7Ev/Ddy7ZLEMQhl9s9FxGlN89Kj+gP68r6IE0kuC
JUzjDM2ep3G04AKIz5WqKBdXa86mjmPF9M9IL3HRgvEaA9mR3UVoJ60zav7+4h5+t4QMZ1T7cemK
9WUnUSoHzqH+ZaSshuKUxcQHxDZXqVE0hyRTaGH6kO01m9176pFv+D4T++VfsvtmnR0yew39pf98
XsGCdUqvmlYBUeEkBuuYL+meFu9XfwnDEP27nkeGYQ2mYM9Wc36c7v0xPddqfvAgq6CvM5yFpnB2
TfPTH7rrQuCZx4JZws2DPPr5pfSwONmbLTB60eaP1PJ1oMpo0gWsqvdfIHZMd4O92976yB5T2OkO
fs6lJRbvBvWnLUnqy4xkOqY0Ivo/p/+rSCi+tMW33SYkVp8dRIyxPjME0XzUqvn/zRdjQGzILOgY
mac1zqNvLI0NvGA8C/TD68CHYjv2XtJmAsCUAHeT4ZHnDoWZBuKlWGqNh4Tckjv+Mp6hf43nQZ/U
5AR+pZLOTHrNmSBATLkXOJ5GyKh204DWty6fdyBR8BwOBo+/uXCzv5pWelvp8CQuqK/hVe8PJMNw
zjhQDffIh2QBAeWGOCkS+5u7thX9NsGHaYQhCiLqO7ejPxYxbmohkAlwGbMMRlt9iBzHeMkrKDGi
6tOVtFkBb+7wN3Snyf+Z7S4b0nLZCEomFGLSCub8HScgJ0MN0+9SOIF4c1CDCU+aB5Rw/KYvrMto
Rr2DlrPF9CZge3SH970Meu4fTofA0IeeOuXEqmtaISjnDrYx9lFYAalEVmcogUocyFv4H9GJ8L1n
JUKaUgpKIbT2ozvpn/4uxXg/1rk+ClQJLPFuC5Tpk7XmqRjknFHk4Cechc0zu6PQXyvrd00D6ABG
SEkZ8WjD1CKkZMMbY1eaHHGWkGIyLrsOvRqvjYi0Jw5kJvUsNvh9lIQOm6IjeNGdmDcNFrQaLaql
n30kjA8GxuVwXbGgCQRjDsESKGwiRZpUt80uMd+5xVmskPpDZ62bPseGAgOmSVt4mX8TRIfRzcrK
J0r90YnBtvWxEM/AUdBnT5FRVtiWRm712JFuczRxczo5u9MPqzjqVjKGIjJYIBcX4JV035WBu55H
rZzfwt9bLoFfIWDMrnLedBUMCx+ubsMr2kF1+/oBgVgSyw2hnWOjCIC4JOWJUdQ6jxuxDeMCMuvY
jSIhIER2XwqVxG9jR1eLFxORqQBtvCWBxRfH0FChyIoTwXWgaMTIqD2vZ2Ehl7Tr5ZAwRsNToBu7
swdpyiuQ2S7ttJ5uGBUje5JKFcJKpxroacO2/Wdz30+USdE2OHc6MaUvcO20tAfyxFIDlS/SuPq7
AO4SdhdHOS7TG5rV8lHzthHr1MW8ARY+6/9FJACmM0VK41PohE5DEKgGkCWSSJ18tc49Zs/L0hqa
pdP+JrRTWENwDGssnIlYeNw9DTV6diSD83ChZBEtoWvJS+q/AcquRGnzgRcoIAvnk/YlU4sB9dlR
HaZ1EJ0LT1xHfadW8R/FRuYuH2b+tqos/GpnqVcr0kr5qypDbla0dSbFCkPAJFZm1El8AQ0fgPjU
JhhLbd5JTTcePlnEkTbTWSOXq7MrTruuIBOwH9uVzyGx3iEK7a3igU7Z4jYvnpu32Epzn+wg2v6D
KPPyVKspdJJKRz7bSmyri6EJ2xq0jEQXbh86TujHDDEoAK6T93MGAU3Kq8+4X5u2kjOPWQn+FpV2
CNXYlkhNB04EJ1LlkEXVIoAH7MRQlrO23CcYvrWtLASNKutHuh9v7+Dg3Ykd3ks4xKnFbfkG1NIq
eygn2WnROo6vwbS/1uosVCVeTwAAEv57VGU/JXRQluiHwrc6Kg1E4tS+IQ7/51/u0vurke9EuZBF
7R27ux6/rJB6Q+qPxVqrV1O3w7WUEFpZtXBpEXc1eDY+Y59a+8ftcggqiIE6p8H7veXhLw1gS1Gn
+L7qrTdRnk6AP37MCRG/Zx/wDuALBIuH5g/pZAQ3nMpPGFAGU2Q0C3kqab/DYeT2HE11og4jg9u1
1A1NDMp2uf9T3wvrKcljxwwCGfSqDl+gL0rnO4tjjAu9IlG/2ips3akVon742PuXoNVpYBIKG5G0
hWL7ilUW284Balzak6LBiDVbSIrfX2naGJiqEDhEfj5K2sBFjnJMBYnZY1qdOP8J5JXFfEgQKVrC
tat9FfGTr+KYNzCepEAmdte9wHTRsDfOvD7CoKi/nrXT4DiD40q9LH7gXzGv2Hsl9XCwqGMsBWCM
bIGFo+DxXfQAvU7+dxTlebe2dPrzzhiFBby54kvyBohpuKVrQQCrLqsZeupRgsG6JrpXV9jNCw9D
hkP/WtsZ3LENFv4+Ouc08koljifeSMDsey/4ofJBED/suDVUh+/bV1I112NDpt35y5FFUTEjg/a/
PSsm9cP5l54BNbRDHJWoA2cDinhhXTMyC7puq3VRCtu8NxyO2ib2dvA9pDhPZjZU+pKjCOnIoiVQ
Uvu0mDoNxFk0A8q4/2XoxmdN4H47pjIF/s8RcAqAW22gbh00eGfYTgKSRl65zj6bZvMBPS7Ypyuo
eiW6YBQuEfDiXy7OI7lSzphZX4qrJITNn71vPZ2pD9MC2fAkOKjbRqoWI4iiXjPmU1fK+EFDk8qF
cQiLntgM/Ed7+md+ngqwDQ2qWYKnPwYyt8sDL6GdUVHiKjNomODeaA+RYyD+TpLjac+97mCaqt1/
R5ux8VIYC0wx9UK+7hGkYDBs9LqFyZ4LSy+IRE3db2ddMCeFQwHfKG2SO+cexlY9WoPajMe+QS8m
AbeD38BBLSlBvBYxmkIkkexJGV1FcP5nRAs+Rgv+vejKpUHVz+868FhEoKnp9Slox/FKgJHYRqz2
jBLcWoiq1DXuT+SeAk6Y/oEHptwv32Q0TJEL2dErUXHNqvxHLfTFYFEHfwoKu2hhrYjJ3vq44vkr
wbeGABJ6Y0m4+M1XHlrrNup94/3CWvSNY7cjKsra0eY6aqxil9bMLZ737xMBXqC4yX7K214r7jiP
DXWSpvNSaPz0nn/AVhaQC7NgFi9SKDsznQCN/hZyRfGMS4KI06DzpXAkCJQSrK6k2DOJ7G/Om7fb
KX+mLCMz9XNYfvvAELe5czpYbz8e4W+BW/hVxExCqhEPL6uo+iNbpAjBz6/Gh3cFb3JSU7n2a8AX
XIhHv1XD2FxBPW5ad3OYHv9wclELH/TLG2iGV1ospypm2oKQuPG87agHszBhlyWTAeniIzmyLumM
rTywqmVUs1xJZAz82TxMs/fIhqJmGkvUTrNqcQVdGMux3u1wrjCI8bye4Wdwztd+u3A8EYmBYFsd
5/rNdyiy6JjEgPS/pKe+ZDTcIHSSqm8pdAdyuMMqanby1BIERc8jG3mahGfZL6o7XJiUzwSTX7aj
jDRnghZgX0uoawoX1SGNm5Mi/qO1v5EddDbiWMaYmBI65MjpNdZXH0cNwOhtEtSSE4jhMjCVqgMi
HRIoKZNXHDGJsvDettW7WRSY0s6RRMuNECWcnHRdf0WvdWdCj+WIDxkKVlM6A/9YukPtMJJZenaJ
WkRB3Aein1iDIGeAj311b9YjkchdEQm5aOoUfdSo4BMB4tY7NWIahp7YgDlnNRxzN3gLETxun0qL
qyIyz572QvtGy+QF/AaXxrSR6Ge5ldGdKbqvzWtm6GS7WngaU1a379hVEIkJFeUvGAN+azqys1eG
UB+C194GGINg4P8CKjD+4fN1Dvq5d1Rm3Xv/rFOLo3B8Zz+ZOED4MVGx2oDEiY2KZ0XUwuuDQCsu
pPx9CNr75fOiXhbb0svMo8cL30d2bRiR62wuOsglnfFKgS6tA46my8ISORXujQlefK7oE4+iS4J0
Pttk31dIvaYeB2b/bv81262AQfhYxcLFVPFciTfiz4CIw1zWkiA08NDDnf9Z3HZbpgThjlEelq4h
xIdMXHyX7QPkIwV7b0x6gJDYtNQAjMeyf8hC/VZTZakkJoyFR807DMlXx56ziSb+MlGG3WqnEDeL
IOPADCFHmYWRfEUzSQvH6+FqgfVXClSbtbZoywrS1FM/Y16ROiCJOBvUSOHqmG8ke9057jJ6p3yi
slv5l5Ff3t5AMYPb6cUA0wWhvyzS3w8XdWH+PcYPXndxO7FpbkbDhw/9WK+JryVlCFA9wmgWHLOn
Hi7ALv3JZwyBT/fbTHW5IPWVe7Fl3+xF1n7weLFhFwKaqA4PZ8fmGDjEMl4e2QBzLqucjbE3qQeO
7+0eKJ68NKPumDUpD/EBaQ6Bu1oFLWvTRmONAQosH3pV4etYAx+Px4ARAxe9hknEstobablnil2r
MyytnSD3n5AuPjD1TTy3VEhF51DKDShsG4fXEDVT4mA+4ZBYYhE8hf4ZJYu2iv6D6rXysiuW0SAH
dPXkchFREk0FVkjxza44VFCaOZdahgk2y1D9UDjZUEumH4BWgUAA0NSmpKMx8wtWrA4CT9ZThUWe
sjRJ2o+iu/4h5pRyQeBGR6vKCHyFZDEhG8Bd4Mh6ghcW16H+EIw9xfieNc/LkAVqtOgvAMYS+xGA
JH/xtQhlOzT0kCsPyfO29pN6vcHtaF+rq6vVZee/agGRXnQUm9OHpm3uj3+7nnuDeIhjDHSm99qA
Xsqk2DoSwgYscsq46iljXvZ0HIRFCrvBB7EaZ1XU2QShCJJHzKli0hWbeHROa3ah0Y3WO5MvIGhg
C5xaKG5HziXgUGH5mhkiTkJqmPjA3344PTPwCToiiKIFdCpZFCEh9J5qSeidvotu/KCVoqajxxf/
HKhLBP6M7CSzOJS3xcgcye3O2Ygs0Z9zLUv23u0Zt9prgGgwUJJ2f8/K7ObIAZspfO/wx7z60yno
ta1B+WUvyzDwAoxJ3K2Te9u4EhAk0WoOqDf8++Bi4XD5xhNUGStHrddHllGD4Uci9f1Qwku5UWGY
FuNSj6SUDHzbYoom+UMEOirkTe6TkCtRAQDz14WvfGFWWySO4hczb6sfWDAin/PJsgOCdDlY0evA
OobOWHUIlGdS4h6GmvaQHbm045+SCgH5qBE8UiweEhpyVzorCSjEhs/sNA2K/PPI94FCwpAqQV/F
3t0dZMtmXiZOMrCHqpOgUwVWtULThkg3CadFgq/FWdv8okGvsTo35x8l+/WrNQpa14K0dGfp78qm
HW9fM62dhtlHyk6e2aguTfNoeuXRYdcJoZsJwZ9hZd05er16kTNOPRajJ6Hvz1eTUQXZ69K/vmSg
uRPtXedX+eiHijtSolSE8Yxk5tDnkwPhBEku7HuYdw/0s95snze+6I7iXJZIjjoMjcTBrqvyBNdG
IL4Vm3NEudj3sZqvaMlEZeLSNU53T27pzpGhlWwKrNzIKhSMxlFVWvU/L/SoaaHO3mDM7OPF0232
xRsAL9OW7Fz0Oci24vwWincRGs94ofe6FXiK5f2QpFEeAOCvan3yeu4NjlTdqSBea9e34avizHuG
K0JaMkVU09nF1nKRkDd7MDWVP5XWTfqWOHSE0qhWKbi4uf/TEm6G02NeVWFtWgm0OJRqGmCFPyuS
zzZ0tFZvnV7Jdqa05WVfFfUthw/C9IAYEO38HxwJdQAIDB5qvRS0Ni1cHROPJV3RSi+RcYlk9pG/
j1whVanL2yng3EoAMDwFwQ5ne/bu/OsUysbJjlFHaQvllNKgXrJuQCh37fUOlnB/O6HTj3ipH32M
HFFhwxJC8zqOwxTYSZEJTa6LSc8RhyBd+D6E/AyregSbY5J8l8XeQRrDu8sg2SBPsMLR531pAiJN
sC18oN6McI2cYc83Q1CNzpDyuRiP0HhKYctPnjf9jGtnwn5n5EEaAgwMIJlfDCMthtYy/XtTDU4X
gv3w4G+iIfmYib4Eh5iKoeHA//DW8z/hcOzRYc0oIrmNUpEZpkBs06BfxJqNhx7wwcGQKKe5iv6m
95icivoI4qKVtneKx9F1KraTnTpYqe3yWMCLn0/L+5lOFFYFlwoENePPhvpk1nFD7cmGYaanoxDn
8vPrjeov4qEN4+pTH+6MTS/qxxoszWjNkxFArLbMzsfu+hQvjtdOgtillbPsR1jfsbPb3vo+Svoe
g8hoy61huvp+6Gg/y1dgWVZe9YL0LVkHcvu8lyoxVfZdIyFiEUN2JgMwG89Ect+yFUiE6PKJvqQB
uqT07UW3kP4qfLPN9vARGKghs3ztumZBm9tG+Hv5SksDCtJ1+1F/bMNRuB3vZ59lNiwoiVcXfSoL
twp3IqQ5ieYK0uye3rnbqTXv3Zk/V0THmBcBlhl61WhELe3P57ZnMFI8KA1pDy+0tjIM0zGoVDwb
2T4bPlJZtfCMRJsu/cUFmocfnuAHmXyo7yHWivLN15lEVnv2UMTJWXLbRk2PQw2J3BWNJR+2tB1l
dkUsT/vaYXqaRm35rqpM2LPAM9aWDxBo1Nb0QR58tm8tEtbH0MoFaMyTGPJvPS+feAyii+kpIG51
sqi6HEa/Dhz0gv3q2qPEKHwI1V8wG2ji9cbFTQYvshaG4SSLgaOPWEPOhS9zPEDQLJuceGAzYSrG
V6c4YEWqXckh4EZX4pl2yl1fE6Xy0ePRi72NbYRJ5vX68BJUddX8nDbP8mVO/yuG2HLMOViz/H2H
bnZf/j6IRQETWRtlUVoldQhBmiXF5KXFiCTSBqjdsp7adUp947ay8rTSlnzOa0K81jCwxNajoyRS
udSD8S96Mn3W7xOraE7tvDZPSgh6Jx3g7rwHZCWr1V3E8Fe3Yi+/rJqEqQkdD6iNFCq2niV3iPY4
SkGwXFj0TMNHKtGjwhfJ5pVLrHY0SgwgVprr39wgbnLoWD4U26Sx9zYguF4kSIJf7QF3nTvwZQde
hixxdV6IpanH5W68MO7rLNdePlgOX8z2IiIsKd8HOh/vtukR7eOTM3m5LpYTzqpem8rGwodJYAWY
mOCgziJYzPFBB2SID7j+4xzUwndXHirrzI0NmY7Q+/1nfo03lnbKbpm0dR89ECC/2y4m55mlBaZb
wNNAECilFY4OiqMDcNNfu4IbhVL/TaMiGql6SqYIBIFptiRh6VFhRVm9tC6vBWjIuaAIxuffElIG
pg1almy7w23ANmYI+BZEcMn1jP0eWEVBzuOtwsLMPKda2+8NR7R3gMJI4s9y2Vd9zt4h2boYz2/D
0aFQ4+vgNbM3KPvyYklyHfjsqWuwE5J3+PRQlHCUMsTwB2WY/04QVWNsFqeCZo3TtiJQvyNg/vm9
3dFNW5iTlC/3luAXU5fsWhog0XSnPL+0XubOlopEUlOC/qjvBS2ANxNOL8KTYIFENciw1xwR+vlS
ezj5ncnsGAUOBKEOrd7zaK6zYUqoGn4vUY7HZkTIq/KCYx97QA6U4Z4dGyQqyz9pmxY2hnk9Zjh0
9AePgZUi9TxvA3UR7FYiQakPS/uLWTtnG/RE3+/PMRtcsrbHYoMtvepRxaKPnoOk05Itp4zh27dN
xXiqEcZ/dQmpanbwyBiSQPvnmKhb/RQOAV7/GaGnJidl0sdRr1edFJnkinWzUD/rUKfilWd/MZ8q
LhcLcEcSXt4OuteeGnXoIcjGyg3gKOBheCiZASjqJXpBuV6soZxoIQPl3DymBrqBQzydaJV8ARAw
ZUKiR/eNQJTYH7Th27Ls8My0sOHf0GUlkpuMT4qoWp8+qVjA/RXqwMVsnGGy08snokbseHz32bBX
AbnA8YLUW4jrufLdCibsAEVVzGJself5Nc0O6PgP4OFRy4MA7l0GsZMbZc4RHQ4MbNLri6bY/8PU
Yts+9a84ceFtNNwCyOpqpfwMX917keR7vH9PkcUMiZbZhB9y5It71BV3hEtQklw7XDyxHqwVP+hX
yUNJjAkIK06iHWlrTYHM5BJKiTpwcxZvKXOakQYVPVBwuZl+DvL0OjHeK2WSwZpO56bMXKkhSxpT
XEFtPsdCHePAFK2N+EwU1XEDTAuoVxcglyWDi6rr9eGMWeP4ywmGL5WUaw/BH4iFFvG2pUxzEWLQ
myL1FT2NeDGLThtvrRmks87df0bmAmgrc0ORGqTES5Wdy9MH8iJu3HoANX/ABNhwGDSt1Dvji6yg
dnvRH+hg4zDfKK3eSScR1NUvwKpZJ/zoJvleXuo2MZdIshVQEDv5Ixm8MHDs0buxXYrk9yXd8Zgw
STaShFBEGTSJsyajAEwj73oTJzEOexN83uYnBlOHJr8goEDG1EdQEOvgPN1XepkV/al9fdarmpXP
hZZBxb/Vliew+Qt1GHIa1jScYDhNOCKmw6rcO5spgXZp3TV7ISrRZqb2hrS73JhgGu27XjVfb83j
iA+iQFJRreJt1XnDVsjuqawizgk56FlK8iEDAb3pyhdcHgzi+sbVrTogaP7F4XuX2WmQFON+UViu
Wg6dWCkZgO2oiRygNSCKWNx4bFOrgIXSvC+306esrQR8pydacBj3GFzgh5nG/Swf617fOFkUGW5n
oFaZD7nu444lh3pQgie16NmrExg9cPQN2oaiPQ9SpHQeMmGbGNQe7gRl9m6ATwSe0Jei82DdBTv0
SDS7Ec+pEXtGrdd0BDBgiDaTp0uP1Rcr1HTUBswWUYBVt44VRxIErweCLTa2jfM2tMu7NOmKj85g
wfMNR8jasKGhNZuSS81X6G9Bxxmdqdi62hmzTNawlgM3ul+Wx6UCckmRS+5B92cFZe/Io9pY1oTv
aX3ovmcIWDyYX+H2vIM63LuhZtiUZNxKYjskZ3oKPpVYoTzSmBlwz0tKRylAR5Uly4MwPGIfiKzW
Up2K6B4vZ11JjGxWC7IMJaU8+BPEf3B/s3gJC5DGfMK4R1CgToQXgkHMO1y8KQm0Nc9TgnBdFXHz
dusIsldIHUWbtbSi9yLU85eezrQAPxnLOiTuVGSqJwfgU7sp31w5vsBIgFDSECd/F8fv+8JXKD8T
LE1QiBTuYdA2yQ8LCiKvcPHkIEInxwn5/ULl3TKJBiaIyFzqDFyyWX2TR2GwpkKbxroa4k997ThS
0H5qwJrzlgXtBcmq2vdL7zEjRwzfKAfGEcrvs0UHxRfSVLHqZiiWDMEZBCDGQ8d2g/c0/wj/KsxC
iPEj1RhD/4XxJVvwDRoGYiArcCpUG0xEuk4Er5raEuOe7PyOY18LYk/3BEb73gwj6JA1q9eIU0YW
CH9t+Sqp14zo1Vn5XDbBa4ubVIx4CEIFsTDMdpducFBQwh0QUUpJ5ei8vW2Ibzf9GXAwzdyRjbVo
0fraJlyR6by08nKjK/vjZh640Ul6sFgFHtbFun+xtruNuhts9gYStuFfdrxFKBZ156SaywwB3XG2
dJD3BEa6WCs5gge9LGIV0eE79wRzjJKp7g9/QdXxyezFXp3KSDc/Iacpu9sXeBYh/wlsBNlmYaiS
Be++pmDytZ+4R9kpbUjsbAuqZGdLN9Z5Ri+syYAAPFgL7HVC4Bzgj01FESM4uV4zjWU2I/snowB3
SG5cO6c5MJtQ2L9qtYJlupmWHd/n6XTktpyHf7cgE5kBsEimcpdEJukF4lUBScFPEuvxHO21ZyxJ
L5jHP/ll2XBDQRY725hN1hujjLrva7yCqd+tJnVALMe5fQgWsMVQspeggw3+faBpLdWIsoPFqkRD
XPm13/I4VpyHBV3GKsBeRsPl8Eb8lCPhRSDysjz/CABEGJ3vKAdqQFSbEOCJ00NYfkH9LBQZBShA
AL6gPr/Du2A1gj8ylxRg3EwCZAntXiuRJoHXs4x3Bu7gt0/1pnLELxnScSG3XkHcmYW0BLMwb/8b
t+fPx3aW11IjNhJmiO8NeKov3QuqZ/ljwwsDvcFRt60WZSUrgT/HdKyYAcNieT9PlmCdS6OWhkrG
+w7DB7V7QKIjxl3pkHZt6AoiGSOMICqqgw4sORbCJrNInXknsLk8VZDo3PkrxKuRqNu0G9Bg8Nwm
MiALeiqJCQwtrDoxGSDQlJLC1VBN/Y2OBtQjR8POnyVxjC0IMBvnh61qBQrWkNb30uD5qEZdTB7S
gDGyJv7RmHvjhFfvk80wZPNMzSJ/drnw56BCL6KExxGY2ZP0pL/G2WHIPMJgzdbC3uXEgXtGrxxi
LhqrMPHS8+tq3n0lY8jnzWR5HJOG8Z2OXoVMhQ7K4YJO64DM1/hURm/+9qNlRN5TJgSwPwbK7058
2GIhBqc7U7jAvjIEYN+YuFjS7GUKPXCLVJLFFIzv+LUQtr8C45om9euuoiruW5AqHkgZdBHzS/Dh
GBD8Oaz3RYS0afzfuLJZP9Giuysg17AXQpzNR+gSmcR3E6Ak6CgIebKvp97hCtcXwzF89PDeQl7O
rtMjgKvY3L5opskAwEH0Ot6BKfqWfPfAoLxEHdE000rizbMdaRD9uugRSffVuphEmd6IEsptbWPi
G2nUuSfQ4nJLIUZvV9pjpUaRSJ/QhRQeE2zapQpFwQYFd10s7sjSiCo+IUsQ5mqxsJCUtBdL7Q3n
t7m7ijUKNoIxP4ROEObGuNl/XF6QyxEukd4toRrhw1Z1EmfrqXrt22tnA2zu/nAk8QUaemzSUbb7
8OUelYSMmss3E7jeiR+azfetP/fqypWj5izZTwtUxA0/+i40LwXUWMDkihXxL2/2l2KGd0jjIJDX
mrrz/FoIbzol0btMrfi3Z9MyGVz/IL21DnljRNK3o8sOx+UY5NPCBVZVdM3NaY0F8579I8zqhx2O
294wLztfK/GmW6k15+FhIuZOkn2T48ksfXEumar7dLfevAzfLzvjEmNQPVKOHMJGWZbFHOJsiu98
Ag3Xb0/ukwLL9LuF9OU6avA6pkyuw0XyJDexzKM+bhoes2/RED2coDDuZK46hze3I/SP7mQ9XTlu
LTXdIkIC715S1w3l83ca/0B9vCA3zOPXCL0leo81TSUalXAIHdNpvoyTsAtH0HHtFsMu6LqZExOo
0gFdJZwnGuakBPAQqJsxF0oxnl9RoZ5d2B96/glRFkedHaE3ts16Y+krLM90BPQ6q+kwq+bazcAV
Gx8jfxTAqGq4qmdvp0fuuusRsdbEFLNC6hBQqjo4/syzDmo2qbNGrzaUd9J8tPC4Fxty6/SGjFwQ
v/ei7pqUwTnLjx0L+BcmwTp8zU90z7Eiu4BkJAaHixN3j+L8Tbtg7subHVlEnXxzN35G72jz0KZn
j6aJkqPM/bvwZRaSGXazHupjMUj7IEWlXxcdvuDU9i/pqEbw1By1Z+wCnIPFUqN+V2MrSHP72jVT
A+pwt+PYZSpoEkRRWtfxqwa2B8cHfVi1FJIaEdxaKkfWIxhj0FqWlNPVzvGYSJ7ksaELEf3fbYRK
u6zdI6e02ISix6CrYR0ZP1sOPg2jS0/6yorpRacRoQ/ZktBturh3zY5r1czfCudRXBM93J9IArYh
X/D712s+D5Xjc5eNAJGPGNNd//LeMgCTYz2sRRH+JJwtjAIF2R1flysvGPIYi+tx1wSf6fxrAOuK
C+M1Hvvga3ZRxvzopJRCARFLL6gzDv2LxqXPcRuuq7HWwroMQeIpcRHxkTjBBwWtcsJ1eZWJ2Sin
93mgsUWLfoluWYhrnq4dhisEGd1ZuV52QW2LS08R6gXdRX3IU1NcXbCE3xtPAg8JUoioRALOHc8G
x102fVt0UICB5wZ9g15qoyV0QElOsu55ud07F9c/EFvjVPaD0ri+HXs/2wn4sVayAcqXLUkNzfdr
KOVfraWY9vVcp7lkLh26Wm+lxbEghiE8dWQer/cGT6Zo6Geb1U8cb/NtCURR4HCAeYjiusUpgiOA
uztj9trABn7GO0gH25IWeHHSjRupO2D/inKz9e33bVr5l/jpPn2xKrU2WnVPNMuH32ExQB+WHbno
UaWC87myiU9Zo5AEX6wu/p2E9U6TAqgY+jhoyzUjx6PEn2ELX8RQHxMoRWaE/hvDqQyyaYZAa5Fe
1MZ5j4pnCVhgqpwp0pJ+9gSGVQvTCRa42/e1hwjiu96jACeS058mWP+IXGRtqLCbmN+DTkA92E4P
yxjNt7BwnQpeYeaDLe30heBwhrUipRCZMdrOGq+L7qjNruENlfVpTOAD7A1vQrR2PbnHB4enO1oD
PvVgV1Lw78JHieTFz6bifTAI8D7/Hzt1aUC9ocRGvj6CbJfxSYGJXz3F9INNIim9j2YnpytDJHFr
QOhHIfefM3YpQtgWSlNmooGvag6GPQpRANhL3hOY65jr1M4KmpSEldOARJ/HQzCTEGrhTs6AM3Jr
kGRWIfZ95T1t7AQ7APMu5//DyP35hBdmlAKNyCC7qL2Oiu3CsQOrgGay3EYL3Bo1w+3b0iLxTxHe
5kk+9Lz4cAvSIuLqZjQrzVDv9ZedKj4/cjhgYWngnkNra26iBWFTiIuT+CcH9lRuuRQvdG19tLRX
1IVOmhFzVjPrwNG6FL3OeFRox/vMt6TMPc36zfBl7NI+HD30YGvmkjhmrHm9EzAYNkemWmg9kJYQ
wFu+PVzk8Ss6tXgsz6H5YoYCDU8Vrsvw/iXKR+a137TLY4u2P9QFcAIJspmOBeLq7PU83wV7EB5y
dEllJOxtbmVXT6pP2th03dzEqKB5ii6sp8nZll8xFsk5LAE4mg7cSdEP2UJmBumSIRHA/6xmM8Aq
XCM+oZTlGydgMV9RDf1cd6o9QyGrMUTzODx/lcIW1r6ee6Ro9RyPVxFKwRzZQI70PSrNbNBxwXuT
BZ8y+81pP1ReDjxGcca4fms0GsQ7c1ruge846cjzgtCeq/FmMuqMDGXTw/ldhZFMvjL1AVNDuNON
v3ZxghmLdg8zx0plvt5oI2N73Lo2uvB20joR72vYNFazGjy/fOa0WHbxkOtrBA8OnSvEnRglh/Dz
uii20P6vxHs6quuiMXrvYiF0Z1u27QnxrX5AEacBM/934JRJr18BPoNMKX62yBDPuV+qVnzz9Z8w
yqa0eAbP5J1MGlQ9+CuN6/KjjszLSibIuDJ6Sfv2w9nYPn3F+SoT/5HDEUs0hza93HgjLxvyJEur
QMQG3YfLYE4VL0jQaboRmsQ8Rcy4/5tvBlm84jTRBhE0gm1lnebOuF6lE26gu5XY+84Zcvaj08bQ
dgkqculMDSzoETCqVTszauf+EEBJhRM/2VJi0ATOhGrt1ZSxDzHLNkdj6ApXomjNKGImMIak3NR6
JD6EhyKET4KVMQ3chu2l7+JkLkleEVMFZW/71rnfq9KAvO6xMuCwn+W58rHfEzwvs3OFljgIYvQn
tw+wdhksa60jsXxuGnK4/fPAOoZliXV1xqoYFwBOG0fejuKbhKfpxvvl8FzQeiUT5PRNDqWNbsv5
FwxBspaP4m4684Pm831f2tjdAQ2AhRbERhJSFhKECoo7Ryyp4g88+7tIr5iYw9L015IRBsYzpTa8
XUwaQicDzSBcnWww4XxzH23w2L4kqJAYSm08rQdbVglBsXjz5ft1va9SsUNWTQ18uI/RcHyJfT2m
d0L59+JI9bwKoq/fg5UNA6ADTMU+KX/bPQbcOn74JYTLel+wJgbyKCnSjDan9DWuGQ1y7FZr0dw5
t7SZRfTdX9TKWKw6zUgl6f7npt9uX1eJsT76l9JEnArpuAkw+o0XOzwHBXbnII7/zd659upkXYeM
tKnv5szvjX7MGyFo3dO65zk2FZ31DfNdeTWc+E6jrMsBmChxyXq0ZVtjZb4j+zMQdr6ePiFV7Weo
7Pq1J1Ta53OjMukH9lnTLcogzoTuEwOk4grqHvAI+9xnepT7pwG86JtC5HdVoeSQer0tiZ4Ndobh
ufVZE3ASocR/vgqWnJTMsz4j8iHRBadANUPxR7FqwRboGXf+zDO3zojIeggUvakKcjJN+A7hV7PM
OeB5QpO4Zgrt4MgFNcFLwom8V2FW07O8nuGcmggYR5bLufw5uXEooW23LtOG1cPeADkAylbAhRJq
fh8vODCrSHz9NAKVr3enOdfzMqhyd4iMP4FZkMeMUZ5fmknGhSozpRtmIgXEXGRk+LEBwLRi6cJg
nRhNl5+I07+wsrSPEL+8trIw5F27uNF1iMt75m8ixX/OSTKyqE6gPkN8JI58ZCzDIoaRWod6IkFj
p1/ASLVsRqqDYkLKw2/6RT/M2iI5H7GLllcJYj0/hTBRSszChWUpZw4wVsGt0TzVxUhuiYTxkgE9
OJZ0Xnaj5wIIpo4Rkw8rA/9RdoHYbMmWplbipWvRk6ZDYOPVjFKs64AkiuMFI7ETmVzktMhpIcXL
QAQWxzl40hY5HYkRuWLtWMUZkNZob5K58CJGib7GQk36JGeetiEu7L11KaKSngZ4ot4KhTqzOYw3
aH+swsjL3k3vreQEDarSdyLJSAl+Y5b+0+L2WxAUkNpwTNBDH6XqmqMroUX1/CtktID2VyxW8SFL
P9iFpW/auDABLBGMD+v5/Y8pbF2/JbwhGrGO/VdV5CYHIeA18dSwhlvoFLP4CYaSEKuaTtViXsPa
Jn2/CychBirmi7seqruj2+5yO5gIwZHdvJg+ge3LUUHSobxHEQUk895GtzSUjlWNq5gIplH38YgM
JNNZJC4HSqFo6jhwZ+7T1Tuc6kzH/S2DhE6r2zOJy0WUthbL0UTMq2ra3T/LwbeuXx0hPh/gBvC3
KwLu7Lkdm1hV8HksdiO//vycpfYJ4LdZary+GEQ0RTlFMqctQd3yQyc9/OjqjS3sTWI0vNf8vDz3
S582toU0b6GBXPBESGDkO3s/9Ce93cP58vG7EENgf1ssXPYpAJi6kGhNLPV7Yf99xf0NtMef/hK5
0b11bnwtLhidI1QMYSJGfwWPlZA972QxcGxtRPPTE1A+myZ8+8Qf28k02xTZn8g2kuEitEtBlS0I
UwP4xENew0YmpkIfI0gVphLGKp81cltwVzCXPn1NZ+frdrgasTZo8suuGzYiYTm5xZVwZS1EFc+w
2r5U/0VwkuNBiRCtgGH5qwiZqxmLVvI1cZwB3umwXBPFpW5A42B/g91MpRWPFGE0QQpMW+RBRZju
qOvZ7sedTl80ivitm24zjVgRV0UOqGuUbvA/rqV4wc+RvT38lmCpt5cbDQhCEObW9dBH9hfv0h9x
9CdoYQLtK+Takgr10Ponxjh+YPtn64lQji3tFt/rLTeycKSc4jkw/f9PJpdPmja0Fh6jwZyrEw9r
EUbyH67Rk+8N3W9D5EY0whxRVD2/ctd4o6/BJMpYJbGAs24C7ojVm222gnie3pnVP6Fx6rBa7E+B
DtkH6HSQ6bQuxvrukftpfclX4k+Q6drVQTmCiZnQ6JX8+g6v5gGAee7wZOkRKZtiUUoonG/oy6vX
GGqKlZ6S2rcZgjcta9icEm0FoSU5wACAKS/kknZAGXL+G3WdqRFwHMv9/7X0LAfhcfTkSWX37qfp
86UtCJ6HGDjqraERvfY5Y21gSSoLqD0WOuzizfBuwyNOZU2eKQ+Z8bP5avXkFQWSUfc2tHBAmTzo
ISQdtWIo5aEn/q5kSZa2MesxR5cJaeWhEPiqaHbSrZjk83FL3H4O65JAg5LhHYxlMIbWyWF+VX+6
VGjDvC5Y1qy74dQiIA9PQbxBRcJbaVR4qISXMY774h0+VCqFDt1yrivyZmVhtS0vZZJwSW2kjiRV
g0AuoovDp69iSjylBPaN1xehUEqdKsZKngyITHQruKmoQoE14BYwOfhDPQs+m5Jn82+HQYbmtlPV
JJvMUmo9FaEUY0FWyiHt7QnJ9Euyn7jsFMbek/wC4cMYA13wy3cEm6mi5bEDb/SEwKt8v+NY67hG
kXU5miq6mu28onoVtc8IZXYL9W/ozum1yZW7lpzNEjZqCbs17ETQcjiXYyXX/WDLnbbRNMSzDAEZ
dTcjKb72clSaSR5Mu8KXYWqjTU5UZHLLvKsj+81F1oKHi+bFLto2eBS84d+Y+FYpsGXmJ9IlERFs
+DjFTYOHudFqgVZyhGuIV2I0lwsJRpiwSncimoH8iHNCcoZtCPxP6BeYd1Nqxmk/hZxCc4sZt5ie
hvNCY3nnCKJnjUNAD3yq7iMI3z8miNEoTt35pYxKDBa34vFP0OjLsndF0FiwH+3HtPZKAF2YYSgr
uCOhBnIEv8a4T2ZjFwFAp20vUHZk1TXPVzSxuRz2fSDFr0tjIkSIoekfhdfxbg5L/DSpSt8SYPpb
gtzxWjnP/a2qZXdUgLjJ08thfcV5iqE0TUK0DV6y0GeBzS02my3HS9tUKl4Z+LxTKsxcOd26ogAw
mg99Pns1/BjDpHxfQ9ggjqA979s34rZdJpjkr9H/RhG1EKvriKP2V3JficAPMVAl+V03uOuIzTlU
3zgnuS6kxW7N2eE5JFAUnS6+VuhADNXMcg+7DuFyYBhqA08EvLPuTbG8IdcwsC/cSb5i3NDlshS3
hJFD06hqQU0iU7md4UU//WgHnt6mjcqLnROqNP6bdigcC0BF/YrpI7pT/NuLYfqv8pC8TEJvIEfF
4JBOBCDIbSLT1WF+FY5XShqB6vfvbNPP1avOj5PE41SHqFFRhmNzdU7u5trCN48lCDLWKUNJMJ3R
uSnFSiCS2LDIQUOnSr1+2+eAzvotBpJadxir8U5Kv8GBmW5cXa7GTRXALUR4UT48uYzwNeRCNjOi
+U2rdr5b/4nuu626grVC4gSLIyzXQOeZTVWCUGpm4ucUdyZwQfqe8Csz5Z78IP2adjMYMIdtG5HD
COBl+SOKom5IBvYSW06/XscjhbiunqEFOosvcbWfHcdYuzlzD+uJPjI70NrRnoEqAHlYHrxpSbU2
flNe6wL36Q7glplJFu+hkb5l5AIXsDQrxzSIPFJbFz5JY/A9Wuoz9xR7x6GC1hZfVV3aW3yh6wce
tdBayXa5a6ITAfpZJcdLdR9nJKgaJngWEws1mx713g9XcR+0LhDFF5eCDv0HWrR2cdjhlReza/T+
LCueoSt9PLhLQ26hWVCBI1yLDj5847B1/VNLvF+Uj1+HckkxNzSn/hLN6MNWR3uyigfyUWj863I6
akt1e9kiVo3SrSoLW21xk/HfPpB+FXJ+Msv8aZlt7Kcet2cXw6BxZt68iqjynKf1a+013QwBOCxG
94dgCEMY6YH5BdUHIzY7hyWk7afJoBqBGLmKuC+KKb5yAf/Ztjg16JFDcQFD6zWEk5N6ip0FBwYU
EEWDUgrxSoMtw2R8AQQ9OlfkWxvlsCZKA94YGbd9dNo9nMfNzlKhEfi4UavAUA2HVeoSRAq+QMeQ
cgPvXgSsLK9EwbtSOyFjihcJR95U3lSDy6cPVSYdnMiMo+7zaBqmtZsZU5n8CWPkSq6fl2EHuUeu
vKpwOcsZBtX3/ISexJy+Sv+wGtS+O2xRGfq4TNXmn8hAnHtVOIfs7hNEAk9V7fNxfikhkuOTQBGx
aLEYzQbv2Duk+HlKr88MN9F+H8Be5dlAMMqYQ0O2MJJrOLhnpkEUYdF4onI4qe8UaL+i+pIKzAqt
20Rvhy+rSwa+HRxnQ6SziJOv3xySDBRPlX5tRtNR77ZRGG0vzdre8R3SklPfC3NFBT4zkFiB9C7g
QWq6IiMbF2ltEZiPs2g7G6J2f1qDnn7FqjBjS2tBdGWIAcIcF5PNLxxDYh4h4LSLuKDRfFDz1qpJ
vSRQJXWubtkTqunvDjqBUEUiMH7oD93my2sx8lYEK44dqSgo2Y4waJ5Q/I5/9xi3he8SMc+t8y0n
0lUCErtSp7hRfPyhlz/i+0uf3NC2hB5JDzG8kCYZR7YLvlLsDg2gd3YgCoJaaBA5JQA+QVx0nmjZ
uOirqEAZsfqZjAMBSHwt0o+GS8IaSWnLCdzNmo3Ev51YPL2NoYsmQhsfXnzq+wnrAbklHFeb84Fe
84iV7Zxu7xFMM5AR3e83t2mzLwDCUb6fCZEt/MMqy9mkwXg/bFWpJiXo0e52dYEma+bMHlODENjO
HGcfD7UBNTncVuhMJnIOrNIOx9Ja2+KY9LGhABuHSWV0LiVMChV0J4tgam6pognZRASpqfdzhN80
hP5BiYdhOxRuOBqLuVII0r/YfpjRc175YjYrA/atU41/IB24HKm+QN60/8LZkMiDJySe9WKHXAsx
R1qdswYoOxroxhY8toi9A8Hp5/zfc6rYn4mhu6P34bcnvR7tDbsp5zHFocFzSEjQ0vGS+A8Mw9Yu
sa/9ihHMWXN3QVxEFQ7O7lTRTrJ00ixMJ0OCmMmB1n/aXNrnAwxbJC2vU49TtJriITJSqIZhSYhK
bmhy0COY6VvEdeJ6CB0amihCN0ixJnwgW9UFDnKmZUB5sUdop1QEp06Kqz7m0W+4PLWcu4i31bpu
Zl+IEThsNHaKeEgq07MSY5v83sOZ7cWkah5zciVL/hZtPKbNiK9lMON2Zcj6USNcab2nIm0yyhTE
lB/uTvW19oRDbrQ84FxV2L3bqpS4A28kGgClqLGbhaLz36WslNrop8CK5mIbuN5CKrZFiHbjusLv
fchT7mN/Kup+VGULDXeQdL4nukN6TS8hXPcoUz/u2waTseQANhv+ZLYQCEGhYHaVdSsiEdltTxvX
7EM5fLB+SEkylcqOvhcgRXaDctUTRpeNGO9Hs94Z9ul+UUoOn/BGjkaShaDjyuGd4AfvV+VKBZAb
i9fmr2JmyeW109LOdmpDmyKpepGqojJpAtJ79JlHCrHuj7gjKBIRMIH+W5MLDSY5HZlet21F/xKs
n7iJSXRIO5pMBEqOqTF9HXexi9j7HIjy5FhnXw6lL3BxPJbbCL7mcTr1KAxJxnhJun3JFyIDTD4d
HAXtCgPnNTab88ibjMMiiV8aO+VpTWFDH9v9x8WDKGdZuhqMfvYFtdCYkBfTcQvEAhtfUIAaEmQj
9uG8QJIxhKUDs3iwFtOHbNC8oUkmm2PnFOJ21eFZYOLJq7OI8othd22dyE4bbJQDnJIsCFe5VYYt
4MJiwGsu4xV7TLdckAgzYAMQbdLr1gXg1oWl2j9/xDxfO0ssjIcveFMJcuaPf8Tr1+yADSlAYvSW
FfYPaQngKkUbSliYpwWHXFObkkQstFyq6jocTxG+KA3jXMnKYcPA9h107Q0nNRR5icwCuYWsAsHS
sHSXgq4fSZIMaa6aQXN0mqFApfQNgSVXsF1o2q/Fw2oUvNdMEgw7bEMYNxru8E3F5SQSHmiGuO7h
kIsNmXQ7HYO2Rul5Lyw5fIQ/6hC0MyOk0vIaif6SBISu/UQcnKJVErMb00yDXqqZy8DcN3xchtcc
pdVKjTKeVdZR99BA6oKUXJ8NpVj0wYeq2MojuIzrLLBd11INvG2ewNxlF9iFb3ivmXBH+ZhEH+0j
5w9/t1lYXo2zRZbAj+kgPDMDIO8x6PQwp/BZbC3PQBDkb6nvY7jXZksYe1aZWEghMGXhZsFSDKe7
usXR9eTRPF1+H6GweXaHQe7p4APa/n77qp1J85sdvv7n7fCjctapI2z0Yx29+qys2qLwKwla6zk6
tJL1k4RdPvQobgxvUlbp5u+asgwrboglzZE1I7Jyr8XrcIQbUXS4AvtTERnMv4zzthi6Qn+Z0AZN
WfIllSiQaE084Pgc4PfFu6bqn6/YFcrCtRSoh69K43vaQPpBXQSSdxaJk0MNh7r+yzUd/uUHVpvm
tCrCFR4nCB1tkTROT3sn4E/BtWzLZtDJEJQci9tQSGOP/joGx6vT8Dse+XTBefXtiiDR7SQ17knP
nD8vuGWKh/2fkP/PAh1XVyDZc4MrjyrYgK/fRNOZDSArD2YKAMaxaIOX/a9jEnbMIdCnJz8YZKOB
mMFzu1FFnXpqvGhcyebThJq0hETD237WTyp11rf1f3gmZPjuvphmSYRBCSTfuWBku7p49/3GNGDx
WUhc4DZvsgIDJUsG744I+ZHWmu7oqXQA7ClWtl4b2o9da/xWsXiOqtxXumhr3AbKujKNspFDhQU5
w/zsIYdFz75vlHNjVpwnDECud5wgoO1XN5ICOopIRIxyoCRDRqEG6MDOQy8ZiEP+nlxhG6DmMYIT
uwcXdG2r2VdvN3AqmUmOeBdu6XIhinTxYuXyPGOM6VPjm/8rpKMv/363LmgiXTmk5XnId9TMKFSr
sW2kqn64WHXB205spF85paksPCmEqOJaZ2VToLfuRYPM19yfdGz6usA4jzaojlvTJ5ikM8FSjQhP
uT6piD8Vjzx0bEwLmkXzWsbUbXhVSsW9FhnNGynbmLe0dQYFgLMb4mkCv5F0YnoGzYIOnj2Meeyo
sAWMS3E+vvpI5G/FfAGDA+GAYnq4GfxV7HaSCAA71PM8qs4Hoe3dlF1tcEV74NiOnU0nLl7kb1OT
m8bYpo/k88mB0zhyTpm5levbS01fEbjrjIOvgSBDG99bwJ2/I6zj9XTnmNWqcERV9TDN56Jt7DZa
hgBq5AfrI7iysaQCUelgABV0xmhXiFi19UgN7LQZ8daIqR7rQa5x8UE4y8tngiBpMK6veaeTvjBs
ORU37RHGZyVQxG/k8pOunMXSF47DEdmGTA91sIA+SM1XhAxcCxeCaljpC+zz9rPZ/AK9F0Vyg9Cq
td+S0a8XjZ65kyUdRTnNjcXHulO+LLfrbHaV4lI7z+YL5o/TQY5BnySnNy41SyKhperoByJK8xtd
v2Gj9Usr2yAumHZHGFFB/1MMB42aFF2vFkzi1Ij4PGq2afkO8mYRYBLo0bdTvSyqgFnzNX/KTEmf
2IFDByJHy6mF55IaXkjRb4gQ7zJdWq4+82/5u9Y4Ddnue3NUD0EQ07A1Wb7tCj3KVeiRe5KGnweE
IYpQ0MMSD0IR8ITIdfv0NtoraE5AMDKrsgJnWzZoGg/fwqPt6O4ywq6LZDYq0pVSHh/bmfOX4en1
hytM6TsTSWZlkGFHdPrKwgtEmiAVSVY7HdfZtzb7i00IyRcHpFzn+MvDu/2PGWvgAOBtuhwOBtmn
LG/+QfQmUqF578rOjMtYKekbkyFt/c9Yn6r5poRV/o0f85CTxz0EEo9ngJkwg4PxA4BYFwehQ4q1
+rkXGlHBsa+/6YdSDXr9oBPIeu0yQTvJcsd+xizeQja0X8zAz5R/mRqh34FMMZ/Jun2INg2m5bE0
oQrWjluGHKvLQ0lqWyut9mLsCVbZYLDdKCmbIqwz1z8mY0XxldAz43qoBKTLWe4IeDQDJg0qoJcj
+BgZEhZ40GxV/K+ROcsx7bWfbxm/Be1oi8z2eYsd1Yxrwj1bQTDAjekcnOTCbhK6haUaioxPYTQN
xn+091KaUoUYt8KEEYGzpGTcyzMRKPFzlRwhfXcnBXPbvgmlNnsC1CbnMXS5c4KHmX8iw20HxX/B
a35+lX1gE7dQSdPn6VnQXP1W+3KlVNdEfBqIdR+qxL1V7sFHBtCaqM/Cpy7OhGuoplH32zFLLDMN
uYJ32c+lWRIkEkOXd+VPDv92pEsdVdWXlkVWZHgqMWXDCT/A8daZWUh2gHMSEP9bl73oO/NCaV8w
FNuUi8A6RatcqMF7srwTh2BIXXxSQrROlNXnUmEhq2u2zlCvmtercZ6PEp1V90Lz7UqpFJaH4Tn9
yQ1Ql7Hd9pvC9sZ3arODEqBBF4SBO+qRZmoOSyu+LneI9iyTOkwNsGNq2bh9E0Z0UibIUbJw1jpg
1JAGDO5GwcNo96fo9NaHvQn7U9ARYQjWEaCb621xxPYmycvaFzrXadrKT/EItnjGtnRMfGiUJ5GS
gNVLU2GwSOQ+hiCV0GZt2ApG2+I+8R6mjZfjSGFqmg2Rs59cUSKEcB9uKTYtTCnZsF/o1q/a/KcQ
ZUCr4znnFt5HSxau7KMdu3O+w6qqO4X5CxkXXHLagOaQL323Yy9TmAXmrHWVVUKcIeruGqxmHxwe
+JJrvbV0MMoS5mKxkf+T1R03x9jPdg0ROW5Rj6us0odwSwwKd5I51THY3DENbEea74/raCjC23mt
uqa+CdfHLphAxUu5VSl5dPFw/YZEgLD3AglI73syXgRhZaR5kvZXZbRdQo1ZWCmcP/jEwD969vGe
34KiIixK0LQTLafKKMoUNFYPAMMKBgHemAN7YZkGwqmrsmdKuMTwNFnM48C2k0gIS1oN3T2r6Jo0
cCdhZ3Fx5taJNeqI3S7nxaAcvI3nws6LAc7sYyGx5X+awziwM+K2y4vZ1jkCLjS196bd8kGKVMC8
JnGHeBO9vTV0bLQDQQynnquoNrLlMKhMmlTFG6tvEinOv4iQAORLliSLTxP7TrlBV65nl0oh7aFw
7XEd98JCAX9+tKBLxlS8lAKRByq/0noJtB8N7ljLL/LZmlOi5e0KW9jesZSRTpynH5U1O3CgOlEH
u/BSSMBDBv28SA1kutLXhnp2p00kMY5Eac7HVL19BXT0/jj8WOQbtaQAvDaG6sQxA34wlecUpHZs
DBYu2Ra7FCZqdNdCF84/DGcUE0oXyMlyMHHUBVRnzlPNNRDOYcE9871jvOnkibYqflyZkkCDlEe0
aMurAgS/vEh4KBsv3wQI0HxSwuPcv/kZ3Oav3eO33OuwgAQk/Bqgl4nUfZk+UWzhM9kTbwyjGDNW
OVo7hEiOzTdtoZ1aakWcjM/6rb2fFNdg9vdkjednzd7hsSM1/AqpUNzOLrUqvyV5zkAyX/2v/f+R
WWs4yrgu2csqUBFZ8do6Warpb/EKGYUSPL7FMyobzTewDV14C2IbC0xjqoarh9iU2yxuDaix6JhE
y9SQEaie0MJ+Y+crq8PVsI5uUzXoTxMZY+Z3vMusPS3f58WlODHANCEwlHvFwgun/lSoG01Wm/Jk
zXFdPzbBiFghRb6wIxH5Rce+QiOn5Vu6vYgaFjPgo6NHd2lRh5iQSB6qXE7D99hVr1i81yDlV5+c
7g9TdZMt5CERHWDVfkcVpirVAzZ4DEIONba1OJ+8DNUVqifoXKHR5XYdN1bfOFykrHJc7QJai5eP
HC+hzHix81tamN1v8WXy+Qv0yxEOq4jF/UfxFCIGfmux2J4ADn7Kn12MWIwvTdyHVP92YDDqltRc
kQSEu92nHGYF5/temC5TKnHvxk8LAdvaQmCjTYzFxkuQPhEpawpSTc0uS3lraJDb5Ag4VSf6IgDk
JCLRYQLfFudKE6W8SodQc+Q234RiLXpWypnbTsEc67DPyA08EJ3AF+qP0jslDGzlQgag9QMbmvk4
IrsiksZAQydAw825YVkUUlY4zsZsR8wGU0yy0pr0gnWaZy2U+p7O/g9Q29IPXZuV7/B0zyRwpkdz
VMIToPqLdjcKH2mIgw5XxMjUww4J5lwVSvArxv7j3AwyqBug95+olf89KyP0Lai+mH6qMfXWc5u/
c+ar9fXJiqBXPUI6/W272PI8UUadbaAJzdmAOfUMYfT9peInnnqb3xaVx+O0E+yFeJc+AEPc7IWd
UKIrZxqa6eGdcPviOmO26DLzcS/BTS6swKIEev7Y6bS76tXvTx81WARNPzm4Hcfug6DIt4igYubv
PDtSHYa6aJ6vaqSgra99IhTLBJJ7iGv9a8VloUACFAMkfpWZdqT8hnppFF40pf+T2UIax0k0EMam
FlFfNFIhLl31ierRD+lw8v8g4sW1E93qJQtT+X7whkLOE11cmXA7xMJWnMAfoVpR8br0DhAgr2nh
6q/fJ7lDdtP2ZEOYHGaJ1nGMiwaXL1gAn3Dlr/qr6VZqz205xCpwFO1Ncc6ngXHYFA6x9Qt1FbMi
lqy8OTUPyU1GvWhQ1/tXLd8M70w0z3YPNTLZv9IWWf7JKsZoTOp6NBL455gMIO4t66UF/RygXdoa
SFWpgtOoRDa93iEcvBnQvdK+97Y1VsJsI1KiYtJn/a6H4gKs65NOmqTCFax09nssF9mWNcrxLVzn
0yZ7sCSODY2LJlPc/SIWPOiCrKtTsSN4dM1+mTunrvtq1oSdVADUEVKNC3XC+xXN8I2LnfnO4QRT
GqR6rf21w5/zpgHYAQWLRj64meGKRB2nGvA4RLkVJxLkkCrtXDx4aLunISsA8pue3iRX0clJiX/u
9y9xopsSN1VwDlXNh3yYZfj+xvOBDN08jAjG6P6l4A33EZhjP6eDCImhlgEyePAtbkuAxrv8lGzx
MhsXaJYDmQjck5SJJCBgDxDYfE9MorSniyXyvJSGSYUMweQHHzkAQq6ENFkv2fUTIoInyQ433Ae/
d+II2SQ/dYF5yF5iJE8Sy6jTPrENbWOmWt7g0gfvGGbQ5h+lPdW6b4d166BBKCLyisgnrjHRcXOO
MJIusk83J0I/rdLp2zbto0CZfeTxHIJ9GcwZCQhI4XXKMU9sSLioVD2GxA8CDm1RXNqOnERgry0B
jXARbp4G0NXIqc+XbeYoMT5gEtWtKUUm7xn9AncHG42e60DDmkJRzTUxuWCihUdvkJ2SfyRuuRwL
HUvQLlArf3Rb45/csdNDZ57vfS9tMltqLTkzICGtmkqPOaMJgu2X3Rm2EXDmQ+k7Ey07k7Pb+LLd
8a4SLjeuDsBjR2Ijo6oYXjj9EoJzzlwEG9DDMaZrxzYULN+NQVjO6p/va/449ORCd8iroASCck/t
dY6bluFlORR2J+ocdTyyPzzOs0Dsix6rSQxmyP9TkdrRR1p1j0IoUhLbKpeTsnJnJuDCvidbt2Bn
etnt6tBYDg6AR7jUMNT7hgu2XyOxo/ikBtMF0EeWb5qRY4XTW5hgOVg8QoA11yfs1Yguug6qB8fH
FTs30okbQMDP/r9EEaav8xUU15/TdXlnJfeN2puQlntE8vFlSWPkN7fbQR+HRF81Qnf1MUzK3P9j
8+zCUFmXzscWA3bXCs8V/coWdcndFmKd+3fUTolsjLlOwTuEtHpkD4o5/eJuTrIbv8KYDyD3AxQe
F8A21JVc/DpyW+p3s68u9A+y447+D+n83OXWzsF35oV4GKREZct55n2mv4nhAt2jV/QKimajc+xh
LbDqXAOr6q8JaZN7rko7bAVHKt+Rwy/gnnuMFqFslGWJFuN0XOuBQCpwRdee1zO+W+K8z7QtyWlg
AfV6CDtkw4uNB/xFDatgGi/dKXe3Y+wh5MvctyilIVMRRxiwbtmysscYOEXXF4WSJWi56Kqbpbd7
0N2TB9HLHD8L7qepZHH3k9Qsy2YEb5aueh7Sie3+sEwmR4D8K2bwxaVbI5dE/kxkdjF5T/mSj1P3
72tj7VPDKJ0fh+Wt6TdbKEbCJFwWoBD4d9C8jp83loKF6s9zxHiY1OCbWw2j5/xSQ36y1a3KRBAM
ilzOPnxFtFDD3ejt4SCcIYpwIoWffnLhLVvibbHVqvrnrZVQQPhkcvxduHiH/WAtgiMPIMzgS1oW
nInTvWaQS/9u8/J1OcHZaVP6wWLhJNBoS6ScDaHw047gpsEB83uOlIqSZKhbQffbvCqiN3XSXW0/
SheusjzIDJ6J/DM6uQYLrpE9hocBPRdrpzs+V3/JXH7smb4Ea4O0rXeGLmpk+1oTXGK3iUNjB+Dq
tbYi59PZfhItLtpCVtVcS7lwbDwPrArdQQn+r471nywUMDR2COyJU+chq4R+ohGmXfvNjLbS+4bT
EWSUnL9irYw4W6JiTzO9Zr9Zmo1xy0OZtHo4276jf7Y6tu+3BBcyFnkFIWX0eCHDYJt5FzL7Ushb
V2Rb3430XYR0Nb7Hj24swIhZpytCddPA1R7JfaB9I77fyT5dI0FpKNnrKhYbW68LRQ+ADuyTuvdU
lQtQu4bfHWgo9n/Vph+NIvXw3JP2B/CPAcTpSYqaaFJVPckAVt+ztlHSvrKiwc3f7PqRSr48iHeN
PMcp108mr9dTZbS4iCyHCd8nKXhZGYitdq7uFgt95YWStctCTKrInNa+k0UiyD4XjgQX9ccee4LY
Rs4JFgIz72G8Da+8/aJRNhpVWVojmrGV+O432t6cCNVfepuN0CvzBR+p5116k6KqXf911btomu5n
s9fg0juNCKBPH5pzraDb/eRv3cYOUG6/cGiN0+bMcmvFDcOG9oT6ANDIPg5ZtSFpUG0KkFhic5Jn
1iEzMgNZg63+/uMzp0RddRL0VaKKBkfdXrae8f+sUu7BQvivHjrZHyTH1zdEY0qo2VX/+lV1d4N3
1+IrF4NFmQsIbbDh+B8WImliS2jZ/Ne4tEt2BC6CkB64UYZpcWwxCXo4STzNhIjYAG2bCXbtDlzc
iTdOK04fjWv16nbWIOR2gRc7x2XiRVRuwagrdZeowwDwYZkNJtvhRaiIZw/OPdHIJ8NZK26deqOZ
F+L2nwQ0MYIVu+L0QjyzbcfuMt+KxpulYsABnBnyDVjrbwhZH4is/iwP17nrsCntaZCGVnL3KWxB
FkJ0Vb/20bbWDA8i3RYoT0EwTtLpgi4jEib9UoEW+hkgZqpF2sPpaWQdqeVSxC9lmKhexr/cjiFJ
P1Zs79bFuS6cHEpQAldmB0Mvi+xcLpB8ueX7mLO8YUX0rxnLpYVdZLT2xmwoFOeNw6LkZh9+VSfi
rD43ZUF6JYKNZxE1x7Aw4UAWihOBOYumcs/dKZE99q7owf+LvG+HLzvRRol8e/pgQHmFMo2AtZY2
D477ymDHcnNhDbS5mm3HJBnxI93439E/z4RItxseJacxXWTpEONhm+oDci08gYN1gkQNvpQ8rR6O
dRQJ7+EeQoNKC/E36O2WmfmJj+/Q9S70qJuRduTi/eVa8l55bDCVeIVW4VoPGLMch1RxOKbIgOZl
KKy1wKonLWp76H2Ox80dICoh/krGn5sNswBQwDkmOl2HWl2ondH72yiFRiNu+iUKT3V7nwgGtsaO
Iy+wEvbaa/hCuztcejDyVq3Q/G2L837IF2nVWZoVYVNiA2yUstj8v1MTXx3I7xb082KylvUxcCwn
tplos0uaOaOh1GdjMLk9WRuCVs+0K/7+7J/7uTQs0tvN9ZeL6ktLeiYEte6hTuqlg2g1S2sQdls/
97f5QtyKdtvcmOViSn1TwOu/2rgSzLWGaWcu/RRoyhJtWq38Giwp5wzanI5RCen2TY/gT/SPPZv5
nCvlTTxCQgQen1Mou+hJcukgkDR0gvbFvoufRvqiQ1B3ZnEeuyGKUYS2JFKnm/e/OBVURv2Cdx3x
ZZnKmOy9bg1BjoEuKfNIQPvzVUTNdNNHqvEl1+duRZFT7yBMN4cWHeebHeK5jfZRkqlKLnCjYqaA
Vz8/aFkiDLMKZrqagLTFvuwCbnCiJYytCoJQB6CYhp20oVKjy2YbWa3Ou/xmQWExfNeo4vPO4gjH
Ct1f13dKJUWTnUinik+hZg9ips5VTooXGXoGnZr3aPA08CP7zuldpGXWXhoyJr6pM4cm3ovmMT3d
auAJp3IrNK5qZ8+Xasr+sIzqyYTuSOOZgdZy0Tdw5o8QZeH7++r31agutXjcBvM54fqIDZjtfb9x
yBqOcT7Ns1Ci/5BYjVvIF0MgU09GAMZKWpcazVMqj1KDrxKfBr84GTGGlo0C2u5X8pZjeSmWbZ3I
5qfalwUhhwO2+yqYdBszA476ynvXWNyObu7A9uszUBliiZF4q9piY+gezlLXcs/P6z+6tWMj6gif
CHhCinCkQeeG9u4Kp2D/4go2qqGbU9VTSBWNixPHI5ef7wrGzYmbhVXOZ0s+zd5FF5sXkkfXzXji
gwaoJAGIT7EC+JrVmDLBPOcpjsgwEWT0sWIheMiWk4sEMLBD6YhyIWcOgnJueXMWTCEJAe65NtRV
7c5Yad/Y5PK7iav+JUE93/cMd+8pVLv2s2k6uX6V65QKKqmuRdcH9MEj3QpxE5BGqEXxdhoTtn5p
VI1DMS6lrFVC9VFVzwuKy2ZBdfEcuYB2QQE8NngnHj3AhSwX4fvRm3oyZLAz0Dnqjfo4HR8Nn5Pu
rQjyNwf0Lxb7iIV1CtzaNC0qgarJ+Ern/i450FTLLQvbNIRDOVViArHPjjfDiHpojo340qRVn83p
V80MiOg1sm8a+KtXw98nKSEquPtzokwQUiWOb6hA+byougI01qHSsbMxQt7Akmc8VWkciqccczGh
3TC3yJMUmH4vuXWMOc0TvAESn0N3iNo5sv6+UGD3kzZ3nK7wXsxNeXZNdAKOyUiTtrvQR6uIwakn
xQ8wwn+2ax0r5cto3sCAR0o4uBRVAckKvtO0GeMPhoy8kGb88NRuUGVWDHA4ke4lAp3oWIdDYry/
GYT7NTo4SEs9EGVSADW6gHG+OX0gK0LN4eHDVitYN+y3vHs65bpWrE/s0S84UyLpiXgpkvs0H97x
YimE7Ip9ZxPGdV7q4OwHx9Q5/k/QLI0PszZ+XbUf0LOZnnF18KM9ohBkzAVyl3jq1BEE5ESYLq05
IPobxRJnP8OWG/mELmAPQHEgizv4zhdW6iS3nuBCLvcziFbtZ0mndx0YhXoUo7AEen84IQLP8T18
tdNaYps0tDulK231SRSIsMdk8zilj5BDuu9QInpBEKUx+4yey6g0qLOcKTkO8bFQ7wjplY3ZDW52
8upuEoz+b3l9oZqBAg5/Nf7FlpVwGfW+SUXMARAitwzOzn7vKplo0t6QFvSIOD9cI1az4oPcvIx/
9Q7ryGQmxHMqZa30OAXmSwNwHTngYk+BkJJGxytVhTNaKwD7OlV0MqF7zQ10WmXbVGMSkxYtbCP3
Kuh3Pp6lFxIljbp7uJ1iDxnY2NXov5OYPkAzTYbbRH56s24o6Ih4HX+LKXHh620izdh75nKK359K
8kgZC/56NvL8AobpMYbRTT1ZVX+SWJoUBvOjcCm2+IknZCUW4f3NnLaE4yysXeRLNNiW/Y4WXZJt
e2in0OB1dYl1RVdgD/5Wrz7+EUCI7QyVn2xWwal/JsnwWVMDdKlh63kwb0k/tB62f5X37r7AHcWn
upAFSHGS7levdcHu140Lss2fs/cGq14JrvD3Swaw2Am4RQdyfdCkKVkO2pHYA7YxFvXXlo0j7gWi
k4Tijw3Uvvje6ATCkCyw74JoGGg0Nnqz8WpISkV6FC0A1BP0QzGArM8lXhH0mI99eVkfz6jdifVb
82cxPw7oq5wacPRzO/dRrXxaVbaHAOr4LQcuORrKyLNkAYuKZDKcYmm3KVwN5XwwwyMLQqhD8TTT
RniR1OlP8t/1VANnAqdGviFCjlqjq6BntjpG68Rp8CYpbOUF4JZJqUPjhSXaQhSSwFkUEDmg+dj9
5yfu4GHY6ICaS/o46nTCDPvF+pq84vnRqMMrJppFPgGUFQHkn125GnhP+WpoSr+xJWgj1LpXGYqd
qZH//9qIV4SeB7B5Wh7lzNIpOe3JwS+BmpRJzegjCF5yRjnrS97jQ2cnh7yUaAA4xIMX3BWWn+tR
pVcU4nu1xznWYzRv6Znsvm/DZgsD9m2FeROPJVstDlz4v8LUuUiKklGhDQK8PS4cqFSq+JkuPKUF
uPdBuh7VCfE/6xIQulODx2cy4kC1o+VLMiZjB5pnqo6JIdrjA5MlUHLOhOhvLRX1MLvYM1FZ6IDQ
DfTuuHSHhYkwHoCiAwj2TmL48fuj58pdcAciX4Tx3nIl8ZxkBNkdh2vWB4xDG0rsTYVhHAl+1lWK
sIZrQBNfXFynusSRD9/w1bu7HfdcOVfL2jQcsXJdMLHof6C1pITAAJeh7u7ehOCSyb1X9fuHnPjw
7oPrR/tSt0xed0itUOAsfCwuCl7obpGGSowBO5Nl9z4KC6rtxHSVglUfEmtSOjf9+R60EQm5Uw4D
EKZDDgv5keAUSGKK27k6e8VM8CcVM4hk97B50AOM5DI3z8grbQ2TeFtsJYPNAONJOoQDVFPjPQdF
l6kQ+gSdWGFHIQuIXPHUz+wzfdSfBODONBfN4zpor1nE3YI89N95tOswJtHWeHPAUtE72gKFwPnX
c4FaKeTZGE+H4qKi4X81Zm0FMw70df823gQ1PJi9oI37cwobXg0m2ZvErkWQUlhiOlEz1kkDVVbM
8wjG4dmXUhIpUnwAOs1E988HqDmFDvYGDn7SXebLbFEftU+RX7DLxGmMR2Pp4wZROyL7Nas/DLYT
QhpIuLYPiZ7+SI090Cv6LuvVdy3yycKXmwfJyP691jFKLE8oO+9OJKGC7G8yowltSHs0wQ/1o0UN
aQ7LiZVb8aIXJX0VRfz368gZxLCTKJO25xhauWV4Cu98R/w1UDqGckHGmYWtkB0Dl+uJWfuF7Jii
yzLgE2Iw/EIYJo9AykRr4gvPM/oJIosfBT72eVY07Cgj/vS99hAKzrphOQP7twa/e+FUy8Zw2goL
ATWZEHxUM90Rq/qIfodtSUMck9s83ZriXW5PdmcJxT5YYDBBQH/ADjtXg/uP96BIV5LEoGPi8NED
C4hvVNjW3CjxI1bOYCRHBLtnjIcW42LiFd+J6A5Ibqvtf7TFd20gUxKdpHBLDyLUr1/1uDfpiwMV
PO9rOlEWBEgiu87dxOofmXMjqr3antE6TNG6NAlt2Z+xs6YgBgxOVabMA751j2nqrL6CerQxbe9L
5Stk2sg4wsL1DfBZzJb/YHL+r9+DxNrmz5wBc+G2HIukjKU/fJwoEBflPEPRjfrnAYEubpcP05EE
VYkG18mSMbJrxNMWt2MRgawixf4k6ZZNNVwSHutcgDNiHpc0u3njfc+JoGtv5iNvvCVxSH6bVpIm
t9X9V8aQa4SMEt7y3VEU81mNmUzltDe8bCT1kAtWmHyNSTsgsg7c9qrz5IGXDYamikeFGji2zPot
wVbWpf5NJy2QnviNuYvCu45snTnQ+2SvtqgACgkKoeoP7IKCu5Ue79s2+vIHc8mHJ9wdtIHGOxIF
UouYNH2C3BSjOjtl8Ym++SYTzbfu2XgBk4m1giedkkh0pUm43Q1/N7Jvh3XpVKfmqxxxMasALZae
jSfpPl8NyGECS+2oIWW3Sk9Nry8zUWQIH7PQeRa46EwvuF/XUqxAZK6dFTwYEjkbM5hEmXpAD3JW
rap98J0pTkYl+cbEfQLZbPzyWXlCS7QWnC0l/5z2iiRXrlbE3kntO8s6AIXwHYBxcJE9l/chT0gM
5N3wafIEKBygsci82WhykK8ONMiKXpoJjX9o/jqTQSXlxcsojapQ65/Y+ITsrn0+o0LgvNAgo0v+
/RHTVn0at1nojabMF5cDx96RLEzbjtrGD2B+0tfZswLJSRzBayB0jD6EzOqQ4LvG2MZHecqYAOAW
YSLisAFE0dlQG1miPcKV5DgByXE790GRs6BJcXNtbG2fJEI7Jo3EhODrWFKnPaIdE4rwwbO6mg1B
9bxoe+4jZwPxKZUnxR+lR6/fAIR5NRFvVUu/cD3+L3mEBrO+epLaZJJ/bAw9EJ1lC+LnERlg0Cto
kUfYI3Lq93MhiL2N9SI+csIWdPLvvxSFl32bbv0Fw9bn+FH/fbYE+jOveFiIsyq/m999qAwTnz9b
LtIOaPCEe5J7D/WW4cHIcKkdsWnk686MLHHiH1QzouLwQFyq4RiJjPHBO/z7SbugDY4kuFXXWSox
RODOkOprSfKh/+ZNM2IpMNMLbK72l9RdzWZaUE/fUv7o5f7S6etmin0VqSlPcyjPWb+IyjRHVESn
5fFyqQUnbehDQoo4u5Q1UrIlROegbvH0Of7xV8Y/V75WagkjWcYf5gE84nzmoHW79Rg3SsdD0cfN
RTqsD9sjRE3ryg37v5a7y4OvZMxUkKxunU8pib4mJgXH6bwwiHZhU5k4ULrrEwb/u8rb6uEZw2jN
rYgAew5P6Q6cZ2F2dOOslTQb+0E9rqADN2CaxyXNCgT07dy/B0Rir3PAQ/wKNAdQuhmLyPN9Poo2
hgQhO3nnsKY0DfPck9HHKNAm7UmNJic3d6rawDIbs9mZvHBG+r8tUAAerfWlQ8U/xGzj8gSjjBgu
6eEa3KRJRPwIsLN2Q+AsULMALRRtM5KgnHLq68RYT2w7WV0azwMBD/V/hV0gRhr1BCzbvm8rHqOR
/glISuaVoDTk/OFZlMIaJBNv0mFqPHzUjQCAF5T6oZjLzbbw6TNdtLnAEGzr57nkIbR8UCX4Uw5q
lbvsRm3gq5KKsn7aP7/L0zqItTdViceBhV0CmjIpH5wq/Iz8NFOFoozb0CXnyC+br/jUM+waFbaF
XjtOk49+O1TIQzSDuOpT6GCWNmwKWrHZyZTMQG0l/GzKnj429JRjO46ZVBtAbklMYgspejBgJtew
Qt4gjuE3qoSkt4OrnzpF5uz49dA0cM2uj5ubMA4CJDxr3F+08bRum1U3pXSZnjgMVq7SRri18trB
XbF+iLF6EBMguUQ0/deCobPbyJlJEO6nxITilfLRB6YtwZs7T9qD8UyAmLlAuFHsT+LJQciNpn8L
hS0A+Bv8r1dhaQBASvj8J8zDNdAnGI4xMqaa1eAzO6G0vYOW/WsPMEsQyX9S6h38ST+l/FEMRVxi
oDO18bIp9mJk2axB9GyPae8jiZqh8H9gp50uU1XHEbL4pVF4jW90ZkxFxBUWaKIKJ9WHY7ddrpnN
G6f+O/HbDYSrWNPwQVFzSU3DIQsO7Qhf55PuWb1KtKvcaw8cGBp2MG16byPLCpNxqyoCRi4azWxA
qSq0N4r4Rf7WpzrK53EFDm7JK8TeqVg7RLlj7fCyUWKaEy9LLUCYcc8zEupL+cUmAUkUJiEMS3Qp
O+0+b/JTp6MN7OeF5TvUxpk6b2Mm6xqC/24TN2WRcV0IfGY2HFs9nxG4F7zod7vIsN2zJjFNhnnG
wigLM7QgsK9tdI+ZB5Pz6y4soK6g5H3V0/oeNp/uYxgzpmtN7pDcMB5OrGaNu7hiYuxTTDNoPRgT
6FPdF7g3DSyWUPjKApsb/61AtQHJROuOE0arQSEtUPQp7n2wX9AXSZv8ugqtBH/mAri/HQsVkmUv
DbP4Q/H7F3wO6J+NDrWam/x2Ae3xtPPMT/S3qgERU6tFfUdw5AIVYahzkU/pvkZj99UxGGXl8L+B
D7hRMZ3Pl61jkYbjtLnOFGcZ2cEP83u+bQhAXuj6QXwu1UJxKkhBcz55rTxr4OxQFy+bzyJ7SLhx
4L8NvpvspCclG/lOgqSlniWvtMIILDacjFgB7FvJtkyMAd+pGS/wDgw0xQ27vDicfw3euozP25eG
ZlYzQxlDf62NBuZsSnJIQxjuk0KphFig8OApKRrFiIKOF831belmwYVEGw9ZbvTCFOL2jz8apGGh
5RpcqbPH85bMkxY6CmsWi+P5hdwJiFqpy2DS06vtkPzYvzENGDEeD6o0cGZMnOuPr8Kp5nPqPLaC
7iYqDrPx0IlFpT1S5ByARHQ9ZsaMKyYxZtozNDYdfuCiQ75327v8Xga5ldZfCxE7uLRAgpWoq750
xtmPSmN0/Dh65jRPbS7QIxe3uJHmwLj2KtPonG8JmpPGtfj3GRhsv/wLi9+kKxrb8+hA3YAIdFFi
BxqVeXklkPCTqGWEzTjag3vanpLu907ljt828+DKvZLZXKXDpmuN7LFlFLIoGxybHJna8ei8sbgB
DmoSqiQsOe+PUkFsYhcEy+uWNlpd8gv+Sg9vzq94y2RKxBBOOIAc44l/woXEpEVhK881YV/uA2/U
YvAcqA32aA8ro+Fjl1qxOFY6NXkgUyTCPQbU41Z/xDzi77AFpITzQSUNBeraSpUCPydA0i+vYIcT
2mtcopAO6tcbV36ZOEFxfngTsQ0FsM7fII0uBFmZm73zlgaEc8jKZufduz260Emag7F8Tc/iKaCi
pO/LhhwEAMgZOt0CLzxskRWWDbdWvbhut5ZI+fITER5exLuPE+7LOo33AoKJy7GvjTIJskKvNOCe
MqQCC2EUHFKPXeuEfavD614mOrCwQrqbFS87+RnR4UrEe7AIkVgkSnt7uF9tdyxMhtJWpUo6y/nS
5DvaIYi3vtAeGk5ATlCzCUmwp/SLf9QlbIs9mbI02s26dDTMslmdp6KiTizFhnjHIy01ITQvwBka
DGIvM2jkim6HuONbXUENYGFNqppmxVj5P4jL6xRbFK3CEqIO5FHYaE4LXlN+rpGi5Je78UGP6JJu
jPhS1wFmn+R6KJc4Ov8jKnSGJHkdavFwGjNz4dHzXfVlZo9zzuuT42fZuR+wC+Oo676gh4vEMi5V
EaApTiX2H4cE5dcCsot3z2dDTugvzyEwMxwGvLmd3hgKTj5qC8NvuaNAlwlyupErDPT/hLEUktTS
45f//R50O/OdM0J3rIM2wF2F7gOVxz2dCn4dWtfDpbEfaS2djyVwLKVXwVRZMt7EMe5Qn7iv34DR
74h/4M7sEtsYiuX5B3I+gxk+sGV4duOzlbu8rrCTmk/fQMNzXZH+Tog7wcff+sCd8p7Kn3VXfPli
VUa8fa3LyTsGprIONl66sqPGeMw+j3t98NwnpRZMnF/dT/VxIFh/hsTFvEGXi39xNC2zPsEaEjdL
IWmSAKD5pL0FqbnCMoV1jZ1QMl/JFFgKlwAkeosQShcPT02IpHxM1iyobiDlahJMNHrYVWdQGMlM
iOo75VbX+JhqtYIeCsUw+C58QHY+xx5YI5bV7t4bXco5VHEmgZViwlKTt1s8e314zYe1xEhFrnJ0
VSjkIzZItJ/3EoZ8gmHbfWEIo7VPrHvAaO0O/xKqT/Y9qjO1L8LNhWW+B0vnvjQrpUSLX0ZPmJEE
OFFn8Etwea3T+bPqtXpRuN+mPXdfB6BJeDgXBceVserDaj6Yjuc/byYBnjqd5t29rGYJAXIRUYz2
qdDaRhPvsMAJZ6zT4r/mnAWSmah+KBcUjpnZTqKrRkUwfK+ZRYC8qARhO0nIkq1gXde5cj/iyihj
Ag84WyC9f1wjvd+GiEmTm0puT089ttCG0SOLZ5seE55fvWtu5Qs9iIIkdB+946FkvMJrRvEkEJP4
UYbkjdc1c4ri5aC+v9fC0WNaDPmkfYxTGkJVD5sj69GMLJYVdQlWx5ogxdrXop3z1+0uv9v/qPxC
o765OiLB2eblCjnf7Ao3xIJQkjeG5BchUXVtg7tfVGhW0MStq7SccC0MBAeHFKflMjV8tSRFeiMn
yTk9dOeLmDidnS1+hIeRcWGT7gj/aZoe02RKwET5gDqO9KW8jIJQpSIotTpmWNlA8LvaoGC/+YXA
E0oikCUSJKFS30ITNT1LdZQd0xuVa5SS06ykIR1wgAnXq+t2QU6VvpnJKcojRF0mw2W2cUfQDwQU
Ek/E72tEnvyF/WCs47dV4gkbDje84KoeZVgJCsDWxhw/DkbQj7eSlufTa31kdWVKNlKn3uuHEYUY
ieohFl/iCrnSbSG2QwrpzqkzEFdQhSs85wpxM+yz3yKVPOw7HmPsscFuHLMccsfQYYbgsTAKJhtn
w2pKZlQ8rFawpyXHmwX9RzjnrRiaJil5zYoq7JxZb7AElezo0z372b03s8ULkDfEdFfXjgl+7nm2
Tx78sgJUuDxcFVE5aK7vjko1wsSuARPAXEI9wVFESVIM4VU1bpBe4w/xyQdDXfFl9l8U/u/9NjL6
diEnG/87Py+7qw+Z+MZxE7UxXP7h/uAGDxOFvL5vBkEMGXnbnSM5tCOEpgZSZ7XROQ5GcQgnFv8U
YgKIp0+GmGLSTAWlrUL6XM8jQ2p0p6taP9xERyPykgXVf3MIDfqhV7Zc5eN+5z+ITBU30Mr4fjVs
VEeScb2nIwxaBOXAZ4ZDCVoU4fgVn/mbV4Bfh7gSDxn3HC7yLtP/8KGXEiewlEBSX70QR92RRF2b
kzOw2i4SoPdVfbB/sLWPx6dnnjIlfxik4GD/B2aRHjX21lymx0aQZQbLt5+BcajB5seXLWD7dwfj
Dca/53l2yD9lGcltgXW1PIOr79Pheo7gvxlLHO7lzCWffYQWasCJb0fL1BLXWKXAi06b4Jh3lJ4G
vQMa7mobqAB0fz2lRgBohWbM8zROL/51x78io7w7BahZKg6GFNbQTMy3VRctyJMKCyASMsAK0out
3z2Q4+XkuQGcMw3j2BRnYZ9zEpKnZQJlvhiNV+EOpYQnl2k/dOeAnGge0ixeQKFromCiRc4Oh3P3
vqrUVD/4rfOPxozl6kp4dJ+IsCF6Qr9FPK4afr4zDfVSNKMzbMe6bfhkiWrpMk2i/Y5Pe4OnwPz6
gm3W8pKZUe/mxPYKesT7kk0s3sW+XHeo4+PPzt+mXKNjXIU0UKSa8j1zd01RPOeepETzJt1uXaiS
a85+rm/noYcpubSTBUvXKp24/kxmnLoSDKH0HvqgE13qk+NHwLef4u61H4kkdxW8HxJpCTRfuOhE
qp+z2mYs/XNbpSPYXwd7d7G2AfYR76YtFi/gy0n6V30bnx6lXXQuZW5BklyrNHKrXUtxcqAzRl/y
Wf42NbyyX1buiNY+FIpj0S6+4XN5HP1rgdPj1u5rkAEerjPXzx2PQxTZ9jMd3hJ4T3kCA0J8JOh7
HcwbSiVpr06CMiqAHvpHlwN1j/UUBsWNAfoIvSolRwQb40DFqH2JoeFZugF3x1sUtSW6oEYLXvMq
Wk2upHXSBOVfurG60ZqOy8RBycSGRfZ1AjOaQMTwhAfiR/azO9XiWQySWHbTdDkXNESmKz6sfKl0
DqiL/WqS/ZtZYjrf2Rhzf9GOIXXqsOLqBNPYBnQHbQCHBBk3W1zW1hRUA3d5InefzhyHURITZpGO
gt7t9DhBqh6K9YBrzSWz50krq1SGFCav1qTgilyNPgLlysFy1Eud/JqqAFjjgKpvDm24xKl8DjOl
lVgvEiYkvX0aoHxGW4eB2XFwiI6cAZldnCl1DwOoLOt8M7o+GT+ykE8u9CnCnkLrfZc90YqN717y
7VVfqWtE+LR0xHMVXSeQfNP6YcXXZ/cmTqVVL9lUsP4GawNjvFOVlSxJ8+8exz0y68wF+gDgNJa0
fvUTYRPoZsypnSG7Z7kR3xpBk5KY29Uc5gGibz4mMBS/l2qJ3yCDpb++RXCmQ1ABuKBMbD5sSoTY
G+sBe65+taYXvz5EMJJDTRC44OOvk/E/cIzDsglOlQXrLGjxF5aSKtjJR7T8ETrIWWPZSbeteiWg
HUIaTvz+YIVnCkFnXL3dNhmBesZbrceJZPxKUhdAVLZcYTelilvoZRmzToTjtMib+9C7cJYdajql
DCS5cQ7RjBrguLVoblRreYj+2cKg8bZ/HmUwXPU6x3wS/312J+nTmTj7/so5O5iKSlGgATJifPjm
f+u8TliHJYaj/uZc90WugDWxJBmn8TeW8dLcepTnZmZbEgbHa1KpyDdl1Jjh7d7fczPjjKR0yQq+
+UoF9aH/5Y3rbMyeMk3T9U24GQVcd+WVyGNeG+iLJGE6et2wL2CsqEiJ+Hdjf9gfQOr7tO/YmFOe
MVB3FBP3qixQl0vGmxTbdOaGzaPdCJf1Z2uKTxnrP3xDybvBDA8ab0FrbY+TmUQlhF69tv/kdouf
flrU/OcWrcuR/38L/d3uuQmkTqlEy8NpyaX3lQV4FkmOXhW/dHLtu88Hpx8LFn+aZ0ZqVlqW0El7
LiYv/ApefMRpC/nl6MVYXvg7P9Udk4/m/iCI8VMAsvYtLj7r7bV9lSMpdvuolDy/KLIZzLujKWqv
juUlY5gDrVNjJxjsgGg3wY621zioSaLmdxOYDvxiUvhjphQ63S9enYCIyHLPRpC9ety+Rj/xBkPS
QmWFIdJLm9nl3vPu41cDjNE3CcaKq1bkGGBKFPG31R6MHCM+ZnFGiUHaUHzTUWGMZcSN1+cTEoMX
/hj4RGazYI/5KBdUFrtJ9dAT3Grd+s7uY1cgLgKbLUWoJgaaa3WmVNJN+prY3SGQ9AKEWJldabfz
SsE29XD9gzW3i6yWmW0Nupp/CsLAGwTkAV7a77lz4anqzTrp/egUVGQPg/lKkGlHAJau253IjLou
eEHbv293mq1ueVdEVhPfi2FpKXprWVdA72AdE0L+pji3JA5RLN5PCVHooPPmlPfUvoyI93hzsBbd
QQ9yTkA1IfFNT8/85PN/sQfm5hnhN4gsK4nGAOEAb8ERQ43vFy1AbTXiFOdXfJQPO+sFQwd0D3XQ
6GSrjnzRCFkacNOGf022OmCNVquemjckDxshfXMw6d3v0vb+t6rsE4rqX1DmYtu3NQzZ9u2z6kFA
TY71lYBuxqesKLKC+gTgtlq/8baga4VeFNqbu8wBe5dvbhYGYB671w7JaRks5NFWO1eWgJARfRyg
PGFM+pkLmZcfytPTV3XEaPYCPGwuG6umSJILkeLQIAA+j2PtCZiGUJEkT0BnXG7rOayAcImQt1ug
cks9S9twawsOhENeeXmDinCs2hGr7TGhsv4XJxvIKCb3hYEUKNmwMbxYLuX9+3Np7VFQd7PRS/44
l2l1jYQkMcp/3JJWPosqS20N6MgPILqQWtIF5F9gswt+KXXVYAh+TyQ+T38BeT7vY8/FguyEOJHO
iyJeKYKzdc4wCSF7FX3QXF/3gyOfE/CbIBLO0swY7i+ESqQx0GfelGR1VaeZfyWa6iZU5zM05hsV
3S8EanDObWtrrGNZ4O0OkLXBjgtUMXgIDygtGGGz0UeTP/vjUuCgYgpmGXnPs6+VJXQbrvwychIr
G5YJgofOUugLmMfoEgY2DsFezjmfXNAcU/3RSY2HoUfuQCu2M5GJULIDHq3CeWXmUknzolhRR+2u
wZ+k00V36WRHDGyFIQEvU9evKGiAYReHHSCm4qW+HZmwsXF1+AbHOeWQurOyZjbRVaoNCBgzN+X5
VdlyuXCTPqPszuInEcXjBoSDBYdVTnMOkqbR6aX6tADqCiGaOvX/5Rey30JaVVBev8DZ78N8gvyD
xLUPZgEmmVEh/YJhBaNVVR4d/lR2LE2Xc4f5lzfFSHd0+KCHPknxTaDT6GG480NzC2XmdG/fpicz
vw40wLlP/KQukvL5ElFnlvLCc90BQN1p9KaCqNgipMeKgAWqI2yYoY1vDA83UWOy01ZQwFNmViOD
Mkf3ZgIWJQDhaV57D92eFWKSX/GN38XMNn+rrcKBnjcmKkXRQuyJhu3COsZi4O41DsRDAaO9jpFY
XD1bmn9pR+PAxlIbrk5RJUBKVIYiRJ9dI+m5GfI4lHcA/yGn36Zc1Bl3SHXYeBKSYv7sjuj1YO0W
sB1BBi6YgXCzi3sFn9RN0E5NBv7aLCWTers5IHoWg7iS8xlsNkaFxMZLLwygOLAjBu+TWLZ2PpmZ
G0QaKTgIPGyXphiM69tXGubUWTIX3+71aoTUjDTbSR1EGQDNrZpxuUFkEhyPUC9TXKx0utTKfi8/
0m91CgK/LLQ+ixTw0ccyCf8nvRcek11ha7iLgWVp3QzVS3Go4nWJpuXPdJ8PXJ01Kaw+8pIpBRqS
Hj77yYtEtFy2qvMyXuE2Ai+qSO4vASgbuaF5PaABTbvbOmLz6wIXoNFDCW3CJEBgzmgHuCg/o25N
3EeQkVIsV8Vz7stPBmg1F0tAM2cFnAYV+ZaJ2icW6HdMR15lIpUg/iSacipt+BX6xkoNuToQCt+Y
kbwMKB407+g1oBsI1xDhUbbhSPLBqGAtqZ7t71uGXW76QV42LGqRF5KOUfrfJFww5YKOHrI4qMYe
z6AWJh1AA6eAxjNeX8o+C/CDdZKEFeBJAUvMB1sS21VScSNyXv8vELQ6chCY4mk2vY15O03udVDM
tPCmccWXEPTFRL+lsv0FYF1U+Lpk6J/DQBumjIKOc4B9HmTNs6B6aHFtuztm0aZoporBeDCqBnt+
CV5jecY8jyiXp6O098IyEiwsSByv6MyAdIwWClFZccH32cRwHUrANdSR75ezLS6xDcdTnTAmwm3X
oCwfuNFYhJLquJXRf2z0ZLiQIth5D/rI/eQV+I7xrjQVxcdUex78jrieYUIFstbJKOJLGK6chuVZ
rQjrQCqJpw+cycd11P0toYvsfYrb4dcA5Aj1GE2den8OcQTADfWwMvZT55vT60jyIPXjaTZBYbK3
wmiHv7TLRRDdhPlhdaTHit7gx1PaC6j4QJMMl689RhyEHyKUshhuCjAdfBccMCczhHv+kvS0qs6R
XRzlSTes6cJU17jNaRV+UtfysblVG0ACHcUMs8FRkR/rkrrD3xU2ZPSl7RSWao5HXfVxYB/Tt35V
aR09kyzMbDSfLM91ei+Zo5NRrMRVuGoXPpUAnc+p4Ly0frZb0hfcm02PBlgat+I7QyMvywnUr/z8
gAkIgV59m7ANQeK8bc+BDws8w1GKbQIZJhp9I+Wy2PNBexR5BGPfxONn4/VfLYtT43OCG0i236dG
Cabkee1VX4mGnl4zIUX7JCSIrY4eCx+6MmRhx8r4apc0QDAnxVkOzbyPdVNf+jZFywxF6K6k//dO
8/vdSfKSJHbHGteCWOtBe9js9n9AAGgRtadoIov64xQikklN5jS8HF6Wh1iF1DzT7ECvTl/YfQs0
5e+f2/+TmI+rwCCEXtzIa1QxEF0ukNCsJ/4hHm/8lMgLhJ2WHoJLBveB0l2AjUBK8TH8JL9kSslO
2HH040djc3IJLH8ZIWw6mtk2Jj+NmHIhTlyupzsIMPf+5eiS6/lA2re6Okreemlc5XFeG/qtpnyK
7q9MRiMF/u5n1goV/RfH+mUnBhMOZCUUP0WbIc4zrTrlemldiy/6eH1ThHxZ70gqtjoLcNj5pNpI
J+9Gc7fx2H7Vj12WWg1+r5blTrlzV9o+UqMOy52O+8dnmEgBmuQSMuJ+tZ7XvcrEOQHxgrg4TNqb
IVqKG+VTTGbrZXby3m/nNiUwjm1ynD4xkG//WaPVuhLBwQ5zolxBaeWWdEKK+yosGSSTnKk8cZAy
ZziECofqoglKjr8yrZvqgIwLe7YC3fomlwbD+kyn85gAMlxlkW/a2vP4zDBNeJNIDeD/hmKVaStw
5FMx/XO2gBYmxKPWccEnN1Ra78PuHXoClmge+TfaFuxjfgmIeV9GS9RE8UHgh9ob80PblOwfzRxs
3PZSlAyT+hkoGoGIKcz/YK81y8wmsteKuII67RM0dgeOlDJBbI7pL3af+9kiv23+v9SKFPmGKriW
nwdqdY76ZF5qP+51zhCgJz2lPfeOVgCGzVQHzEAo1DRXpuE0Y/Q2Z/BzXeFM2DhDBOMkY3+vRWbz
Z6EI6aqMiuV0IWDc5dWYuZq/uKYkZZIUAPaA6ERd9k81YNA/dun8a5KB5RjCFITHJ9kZNv85rqHb
GNBsJr3bpfJvbBDPggknKvxxHU/406DCBaAUAUwty5F2poOc/8gVR2iGcMYnoES1ieU3zesjTlpR
Y+pzyf2phiblm2l3DSKWfbY/J7qigqcabkM34/6jtFvOwNCjhYTk2X5Ed+WOFiXH9fz5PcIO83AU
6XgTdKQlms5SMSIa3aREZ+TX3/aO84aE0N4CtZ56OWgh1Ad10MlXcKClvRFaFjOKgMidjQlsrhdS
gitQmqRM8elaF0zsce3EX5bV4rf4UpDQkHLD6Gf3a5i5HDZkkg7wx5QmzTbTDGpybqj7mKAvmXmd
7kdEeTWrWIVMncasVSC4bcJE/281Qg+s4KFOwbTQNMYvpQNYS2I937uNKQi5kzkm8Jn/RilkfSz3
QU98HZLIcRbgrK8Xo017bNNlxwcF9M8c6bGstEsUdl3co8aT1oMj3yd+uw6phTgaEHsuDi+ipgN4
4dwdaIVsYk9YYiz7yQ6guz6dZVazT5OxBYI62WIYGVhTx0BOOFW7gRMaGP7HvOfudKsO8ZU4mBHc
mHvD0Y9aSvd81QzullSTMcDR/WgimhOtfNCs/7GPx2/2CwHUtVJVTbeXpGtI9Ij0VuqdmuBjykMG
cyAFDDTplQRle+PmgTNGZwuP4tn2kIOpnCqfMcc6iL0CUZ/Qu+0JiIJWrWqF/s24wti/AyEaxkMP
bfSw9b21dYBZtOW2159B5gtOZqLVVejoOH20S3dXFG59PDSxWRZl52S0P/3HazF9ZfDGkf+4dvUU
jy4nedYCOwIFQTZtERUyGfN3ke3+8WZgKO//p2WX7LTexGYhkQ627DzwW4YwvL2uI+it4pv4JgzM
O6ugBC6MtJdEnHFmiEIQaMoXs5NatRmGf1PoPjqtS07QOscB/6eMMjHXGO/FFka7RRj98inlCgJ1
VZEKgRJqL90+sX5fwLiy4rfPKpsjMse+xBUEPLGq7FVdDw2pzLi2aggl2f9miBod2tV18VqOvib0
pA6/M8GeqVKTq2Q7z5NfkDLsOQxjz5ACJczIuTzlpX6Benp7GfIqmJcqrGS7wo4uDyXaaryNjQSm
oIo6pmeB44rYkdVr3S13Ap5laEXFFcNAHOXe1cJWx0Yue1DWzs7UFp+ylR/9fnh8qW9gRiaHY7K6
FQYErfXR0Tk5st4EQBKYcNKNAxApDeHLw6onbo1MUex6OodRZI5mTl1lQ0hpn1ZqWaFh3B+OzQew
N89js5eqms1QVIZ6qR9favVs+xleLIi+IfTqkZ28/BAjcV7rySz9TU6+aq2b4Fiqp4GhfYC3NiRz
6zG550wssPEn2VMa+evNj7HagyUDRuWKkie5rxxQo2j+mZn+ts2NpfX6hARQzK+sFKkuEW7JzP32
tvifM9VuU+LKh0heAzz9NoGSC5cjAPudaAbf9BeD6CZfR5bDEBGsDsNycuqSfOQMuqMfvP/sc7aX
I7AMo533fn+z12Sc9mg5cDIyzyT7Or1bIGuAixk/xmgy4kMryJ030SE/LM38qBvANJRH+tts/3Mg
3og6pj0GNez2ta+Gf0mtbRMaYvbca7jvnPEDvzrdX6XHt/JI0nx2nd7iA0n2FxQ8ERBfTj8HTL+f
u3l6afTgKrLZjezDRrLEGQGX+yL6GzJUGLwKF5+Qubqf9mrqDqV4OmyHZEQasBMLUyp5S41HVV4x
WDTqPRQNI5C5p8yB16s0DrsaCH56kTSxCVvu1I2eyCjaA3ZI40s8PHRTMcUjZiKr78YP+wa9vkRz
Z60ABNliaX8kExrYOGvXIYlR1v6pnvcUBvtaKNlJ4dHK7IdQkPX/dFfEv8wZ8K1H2Xr2qCC8AlJJ
UJX5CeRn1HJw4UMyQ0QLz1EoD9Rcy+Hs0SJk9YEuxFEJbGOBr6O8kwbqk6LVnkOHVFXzNTRTtCop
DbwV4l/2L4ifAuNrdlME0VxnWsTH1X2CzVrg/b2fEXk82EEtQus280s2cW9EtNGzYMVOD4tB4b+m
f2X6eo4H7pZKKl2YeMU8wQ5PLhSJKHVtPW2Ho2gRQAo2uwiNOHOAcSy9lCsHgk3mdB3xpwTF6lAF
EFc4gDl3oNaXH86ED9CKSaILBv4o43gGSC+3ebIsJmX7EsS/aEEJruahBy0+bOL6HMxo83JY/7D4
SAkhpnsxRiKdIJj9Zi79e2mrrIUAJRsmlk9ld0DCvzCmn7C9oUmmBY43ym01VF+lRrj0qPWo1Aec
PPkvnWm9BaROuTyuLSy3sHh4dHFOZj7NmzXZsFZdAgOc8LWJtYawaD0dAjhY89DEJj0C1HMxUq4D
/mt+zjg1cbHolPpsiMOR8zLmvPrin9CODzre29JkmZ6iV7db8yml3r7C0yVln/MpQuLguuR1CGJR
gwuwOMunXlk7EgXzG0nArDxl7r0cDYCdidN6oMRFqSVQVN7qoeTWSecILvSo3LceXdkRd3MEJ2Px
4UuzgjC20jTqFwx1yD6xlL9LVW9UKp9h3vM589mN9LKylQ65MvoubEfo0GbIXjtH3YYw1ukqO5ha
x1vWWA+EPbmfmQHvYDVDuPddNLbrY95D4p3A0RVujeILzAQZ7z7h+5871kfbpaCv6x0CZDAJsjXQ
bSwckWXQ0d/Vk/cmNUrlUKB6eXmDRcQG+cFKfWifkWd7A0bpu2fO8C8fVvjZpAr0aTjmRN/GGYYY
5YoWD0juPvgfUj9Orfij20xCx91grVk3lmPXBT/w4OtlrgSuxGRYyyUhlggd9vagoe72+YAn9EHa
vKrGdGI2DpvBJd7FAlsc690bX6RUZPadSKIbTXyNcPW+q2chSdk/8VAXQy/NwhAmZDSEoVcjLoXx
1X3QcX5x+b2i/b/rfIBRcxC1+7w5vYbVfOgnzQT//mLu8UbuY0IjOeqFNLHGd55j6bzaqI17KETv
LkfAUdKrRvdM/JvtmhzomhQk59u0bUxoYn9bdxsLhZIiiFE+4c7GWvfhJaWqT/FMLby/K0SKdhwS
oQV+JRtxEmShRiUMthgRZOBpdXH8CzdOJD4eGh4T5KkF0Lkl3Q9fy++TCiFDG+41ccTFkMufI/+1
85tbYjw+nGNU1jhqnyF0Y6Q8uYotaDcBl75uzjrOX9cy5nMGIT9X0kH8QniTxE02XUwDZdYg9PB3
JLxdcBmlBSeciLO21QlEFQM+nmckHI+f6lXQ1OhzRn4u3y9NJuCZ8rSFIw9lvGvF8S+ryaXBhogV
y2goveRHLCZSiNyQWoxgbr9wkKaLhhbG8NwoY1iPJwjohcWtl6ake1OPsY+a+3R2WtiLvGzATi++
EUY4wImYo9LRiRG/WpJGjeGdZxQXwcHfnkWEjvUyARRUmK+8NzYRATivpLVsm+AHLAmadVVF0ptN
iWuUhSfQvZ/SBGtklcYB9y2BM0GlMOhdxbjDtow/ZEcFEOLBBRn2F4rPbY2jdLYtxFkZN0YgmNtU
H8e9WvBc//PHXv0jWEBkXstV1Pf+jJ/sHi2hrDaREtO/04ZguDz1060nTnjqABNrIehbcCMLJ1gP
9JshyNeGPs8QlvaZDUK0rtKCxFgRyawjg9R6sYXVF78HQzm3db0Bk/w9F9AdJD3DD6hJWZkiRRDF
A7evf4BW0m6KbfeI55s+kfppL5W9F7G2PwSSDkuFN9OtgqK3zVWKZpDEvLbMsPjPghnrzL5tjBx3
JC2qMOhvCtFQqxTcj9ns13CAw+QTQz2byyHHysxwF0SdjnlbEpS9IiF+LOtwfkS0TljK54z7AgFh
T16xEuo0tErdaUu9JGf22g3H6mJPqX9b1rbL2058I+vp5A/8cgGD55sA+wBTDkK2UZB7N24/OK4B
ayz2V7paOskQSE0N2rDLSuYALBmluw8zzEdz+Uw+rUkBOAWXJhMGY0yJLKF+bxpOMX4YE5n915/0
IEh0bCeQebeFIulm0b04pnae29j9urIpdBJIasqTjNTTrq8DWZlWP85oOmJFNuWHaNi6qvqtfHgB
B2H5UQC3RgUImpL1FDCBMASYLopPmgQtSdDlfs2O/6Mw1JhQwB+VqhF8oVrhWQzrVuJKHr3sH82f
XTT/VkqUopRN07OgDsIbt4luFdELp27hQxLG5AyGZ6rzXbLYfeI/WO0oJFHsg4eQ4pWRFSFWoVGZ
GFfILnf0xNGnRNGH87IInE8ym6wnqANLEWKmrlx89pIQtxqpLjY2zA84J6ciYsLlbHSaSib1hw3r
iICMKTJH2hj1PTAa6BmGbnMJBs9q9Q9t1YCrWjYcwlhaXBhd9+QmMzDeCyX4AeY0mY8PFHWjOiBl
2cYU76qBRZkY4qx2rZblvA49w0U/mlu4Ycbl124/j/vGIRe8UdQqF/9GNzIvDt6aOnkmxWDiglfL
IqOIDxeKiXsJRntN7Le9kDuk7sQjlv7piZJXr+3wOngSLTYb/oFXi9GiSNFhiQ0hqk38GeVafisV
dPkb10qTylFAw0zwlkO1RPG5a78pN7M8zTxJGSDW2mz8u9+2rx27mHRBQSCACoJMCoD4ImIvQE/J
3Hh/ddjYAKoFdQLqLpTqG9uZpET0YebkJXS1FMHqud1Pf7uaGBX3gAjU7Dp9bISiWOL071C/g7Iq
HBq+5O81fkgvfZ1WhHKzQDx0phoPt9tFv1z3ICIZHDFd50o1q5pEPXwqg6dF2GnEuUe0ZvjSAGwa
SIM3p7zZlDkK4R6zqrqiani5u9L8mtr96mvtZWZS6HkudoJ3VwnNo9rkuwLDs7Cgelq4mojBfzoj
PpJVVpDIWRAsg48YghzWE/AGta2bS4iOEU9z6dz7JIb+TLy8QfZMr8A/gBUabAOc15z2iAC57DXd
vhs8MaOcNeGx9I0rCYYfvZm71nxdZXge22S25zWDueKjxzSlo5gcN5ONpC0L/D4VMTCV00aJboxd
VB2O072WqPYd99DOyEJa9MAsRc+ujj1oGQjgl7QN4FJOPLodBSNtD83CbVr9wRAfg2H6Dbhr/xFo
xbHzsz2K5AeHtABhqClx6ey7hbZ5afd2mTXXvH4eTDwDKo7iJ0PwL0jHfg8E/CCozrKMAQlA9ZO2
A9QIafa6hTtVZHTtrTcF7H8M9lhwFr5m+AUEcVQzFmtKCPHMxnnqIJvjGYwDRSff3khFjLjhjneP
vvwDyNDDzOrkLui2t/7b0+2tBcSxzedxjYHyUNp63cUvwWEMPCsKBO5Z4q/7/rTey1fQPEmhUYgt
uWZzpwT57T+qoCCbb4gP5SEsWorGmxUJi7zFjG4s1ENEk0FtuQPtu4n9U4ZXN4bkX14HHU1iXRg8
YKFS85s2RsmsmYdB+ZYdjsvdYdcVTeQuTKdUV1aHc7N6sDm4XVB4jzk+cdCRB2/xKXLQZRQ2BxEw
sfM2NyGETwVsMDSqAqYt4JJnP6FUXBVZrweRZkaagCvQFt9dpgBf/yxxRQBWkC0FnwCZ7/O9znV7
463u/3GQRNRiznh/UOWolOtOv8EddUs/t5s8Jju+3Ezch6HMVeumUr6nqd+/RSVJkJHU2Lz/iLGM
ovmPYEU4IX8lk0prqOcYxi8j5Q2uiOacqLZWz2a7DB8zHnGWagN8X4oiK7hWe1MVCL33KCL9AaHS
X/ZLWhgABkUnbU08ne+6JAe71j20vHOzEuH3PDWzb3T8GrXVNmlfJQg9l1YyFa7zwljgc9GfxjqT
IlG22MvIwMatfAZ80rOFKsyQRdNceSZODoIGwD5QDFBNZAKeSWwYy0e5tZjwaKMtDGL9dPLroKsN
V0UXDcyJ8J8Wvfko2A1QYTgEXIzstNc2Q6WC7Ep+vEFsgXAkcz4VwxLQuNn8ZW+OaECIwlUdqcg3
mnEHBGsqV7tsO31w4dc0Ee8WDUG/knPqXB8dIuQPP3QawsIIgIj/NWLF8ah9DwA2zXliZEyJUJp0
2rlMilTL8FS0QtO9kUn29p5qngOBRzPI6YR3pCm2hMmGXIYaKPPT09NiLrWsh1oO1hJt0YWX+EPO
XUkmKwagHwGgLqQfUJqxob3fOTwumhJp3PJgwSoNzXSz/NmVlxsGPOwopAvEGDY8GqQaam1p0Kn1
c6qSkyQClz+rjihUv2TvaZsP5YfP0yKzygZnvZNVkYQqNwfzhmGK3TQXNtWFyDWes81ritOZ88+s
RIIDVWBifZPSM36OQViY98wQm2RjzJU6xC/fx8ZdbcV+UrKqns8ic+VoiO7N+1jaikiY7gxGqayQ
dOv4No5LzmLJ1qCmIFVn76dA2jOmfiaqW/BgHjaWVvJVdncwlz00YBwsGqRIp6/JmUZCKBdx7GlF
+rm7Vg5aKeKvZjGSMrvns081BNt5RUuI5gWtCoI/KghADwcKg7mLNjNvCGDuBJ5tAnXcgtty3ocD
yKaOxWNAEnHZE3dBRqzOYECscKWhLTBTx3UQsGG5cS+d3fx1j1u0DoiV9MHCYd7ZCfOZo7HhT5Ho
PjneZFXs1S+uk9gvqK31DwIv++/lnvqrlezl/lv8rzzewqSuP5sUdO/JucmCAJ+8Qg2MsI6bBgUo
gHkso9DYedUzBWREcg8F08iny4lA1SD4niI3NhENvVaJ8U9esxnyl+g9pRrWFlUapt4CAWON3znS
jFU4h8twJdm3suJKzDLzbHDXAYopXfcD1CbryOEyNqR8Qv3raUjTg3s5SXjK7UUDaD0CgiiZW9HY
dvnwyhQx71UzzzFipa7VYBQFqKrNBGjW72GTY0jXTh7vnKs/sLsZYXlbMADibMgp6nvoShuPDcfK
PPj/c5VHliVcvHM6WCBFjSPsXE57g8wpu2Btl/KTGTsk2i8DPlge8bEqWbaDF59YRFBOb7meAm4A
KI13TYm4XgW/Xxl4ejeh+UEEA0nyw9rjFmB13xDHOKHMdgQCcOo92zmNKSkgtnweNvluvOVt01Q5
tmatcR6OEaXySP5NPyXEXbMjVAlXM1t9Bv6qjxaWGCmYEeAKc8MPiHpzCFdmK2GlDBzaB3BitTlW
UdjTquLzq6KrJoNGEWafxrxIjPrDPdtNy51+2e9YSPbo+q94w6umikkbKUGhLOroFuWoqnlso14/
7D4X4e8EQQILMN+kAjrfzC0W4dkHN7vObQsV6yQpgNrPv90eEZfCFM5gmtxmUKw5uFnUEB2GDI2P
cz+oToVEJdEG2jbaGC5DFX+AnsobOpT2BmkyxmPE1/UVzovPJCP/bq6MuiCOc00pBSMfNZzxMnKP
K4I+57+FFUly1673BOMnntX+Pjzkr+Rx3MzJYEvsJxvBOiQo7l8wplv7aIDnXL0eZbnVpt+V1svD
8tckjEU3MoRixLU109fE0Ni7QlkbbDcebxU+7m0UwjtQ2dG6oZ3Ni1DGNB1sP05ebWOe6U6Ak1Md
hQTjQ/ISdgSXJpXe8iFWAAASse6rVd41EAgNVkczILN6+nsuOYnIX4oIQHrQxwV//om1d7gtMesl
J28jRIjg9DYfh+6HLzzhxhVG+3X33ee2Ekl6EzKBeHB7clapnC0PRX1wwzGXrQsgIZjBx4ZPyKI6
0L3w2J/XHuIGLbF1eAbKM3XLv5TVCgimjxrb98UhGrmXsZ7DV+BW5lIK1UwkUkxGGdGtYtHvvXHE
LsxsR04QHHK88S6/MqbqgyGeJD+bWx5ABz5j7+ecmXq+U6fg/neBNCRorNlbRvyqYfWYEkjsExO5
Pq8TDmS/XdKF20dcIkFFq+XzCmyTu2Q/aP8g9idVaOzOTMnXD5yAx5SFY76n9lnmz3Gdk/ej8+Xf
jY/wAjkTvrGLlHSgoegc6yk9YuHGCvjChGSTSniwYQpwit/UqNj2WQO3R1So/qnX1qbkInRGM0aI
iaLB+IYWsx+z9TlnHG66JBevuMjwU01INgYXrTjJoy0Ywc8mfbJTN4uL7Qb+NB5a0db1UjYfEfk7
cEvw4i/kE/YZSCARlumwiCSLfnF+vtG6uyXasgm/TZlagAVhs9SDB7KD2zP3H1QyBPvvdQva6Tjp
qstmYjXQmNgQZaxPNGcGmUEyj6XgMZ9x9ViMS8HH6f/ZM/GFIeXots73QKxC5K+DEJwcBbUcRX+X
PCuwTVP4Voq0NjFluDMjQO09f+H18HI2rtOPYgmBZ2O6ElmSDSoEj3bYxhmPOFNGiYXxkOlpq+gv
6s/biJTq/EDeHD2/SjRSlQTo8fE/BLCXkSdIMQR6mzSQ1FOqV6JBA+x4j4CHWq1YSrPOWG9Xk0kn
yNVy6yn/RHUgBI7mfIf/Ac3IP8A7wzr3PSCJ3HH7APefh0rFZAnMMWaq6lxR7O2Jt8NrFC3P8OuP
4wkPZYbyyrVn/jH9Ta4/wjputVaO4Vp3jd8OYE0PvGeWbHrcBhoH5EyM+S6V0EHiQFlD5dPIAdn+
YOYcrqhykGuTyitd7JCl6fAeZJ6kKGzOywPhVpSF7FexekWPD4AoYbVgj0PYkVhhkpbMY5VQDq0Q
Fkw3+XlbVdm6LG1MY3GjoQor1pIZkxe70I5YOZGdTuUSooWSZgbCNme9hhOneAq+8zpcAiFr4JCd
ycsryML1est0qcY8/oXw4mS3UsYS9orSIUjnftOURDHJYUld//Ev8CHl31eq+JZiClu6NAuijoeZ
ECqFvQHAEeIuK1JxWxFgr73E4JmrXVu/6zWjqFGqnDbmEONdotfaDsF3KJFlW+jNdK/RVaw2+0CU
sXWvwJS9/ui8+W3dvgrwRvRzyINZFjLDlepIf7mSKhi35+XZb0vfahFa1cc2l4qx6lJOObrSSKL0
0/kS+8m2ADt/QNxXVQk4um94uItfU3theONlskw8UAUxRtnGagxBO1ZMeKp67BwjyiGqw9SSoktd
gaO4Tfl5y3wPbtvfs/jN4HdRHaiMIzEK4zF5j1sJKNPi4H6n5LxuuVoLPCM8iOfy/f8s8TlIe/SM
taUBO7Mr3BVlcmJ5xj3llYllq3Lw61/Ul0+gUoNe6Waagg6La7CQbIo31fg4dd28Om3qwKmWvl5J
26wlQrVoNPoMJ+rPjNOQV6u2leRtSo9yLl5CDfv2+XBuEiYPnM8oGYsKytyvnnwlbUxXcMXE/8V/
EhScUcexkd6kGpu7Bu6bTgvkbeCBRWy1o9DSg1U3okUKVHEodYXRXgV4v/4tZlT9vIBSsPF1+PsE
pzM8bAmAA2wlZb6VOaqZdMDB0k2VKpA1l+797rz5x16ST3S8hXnkBpttUyV8FxuBFAELzbWqTKi+
h4LyH0HT9LIldKQRPSRAM3xWoDl54Lrenv8WR7V/K0UXm6Qcjr5fR0THzhstH+IKmWJbPNu9AU9L
FyJ72zoV74sVy8i7OjMouKUfuTwc2vv/6bvNZz5qtMog+6fb68qIpzlOt7WCgvAjbwrXspZJr3w1
iKKydHxSag8hC6Kp05fpSCZ2S80+RV7W8VyB1/8h+ya4LI5nEvZyYa0jwG+GqOL9fw3chlvldjFd
kzbVHUzHUfwhnqfy26AB0K+2O7IfGCawsHR7CRBcTKzfu5OKeNsaELWO/2Y9XwPUM9B82uMi8PNG
Z9bdF8vQNy46h0JipLGsPOI7QH0VYcV+sNP6bxwNGl5sqTixypDd5vkvCcdZLFO9b52UTV+QYtnf
URRubqjnVAxwVqlWqZb0nXBXGHoBirkAL+zMkPDmsfXFogAgWOslZyKQ9EJijIh/ciXe5QWL798e
7/nZfqvFH5AS2SwN4igUVV22FRzrZ0TzU7DtNlDFhZy2BW7Rd8BnP00cQ7x6VQDFykUKeH6w04XI
+qPuOz9900C/45CzA0bborYkuA+e4OTUHvdLywqTc3AYCfQ9jODeg/r6ASwIyC3esCkIw01MUh7t
Py3NedFV0S4GJNKFAkWOp+NCy4kTn5O9OLP1SSPLNik6OtAF/+Aw0FW5djRoHMazix9D95oKCSEH
w2USKEA8IsbsOuVDCioF3zojTGZxpAIqXcJCBxZxBtKQ48+N2GBKp4ZtMGthU/XxmarXEHIIqryQ
kJlmEjkNhKhb62xRfb5ytRqyWyvvZma1vYBXwoawhxDsLUOSsioCBbMAAND+HZgQQkn/UcdjxOZ9
Xp8AS+Dylhb1nxOwxl3l5uMoYvfQAE6DJOeDDz/zLeF5Id1zKCRuanEpw8qAw0Aztwzqld94VZ7N
bOvGS4JkK+uPIwFwgeajhtVhXc0FU/x1HADk4o81YFFc4gLMmWk8+4odmQrWi1+xBkXaitk3wNw4
ylRcXPW3lkFXBJM+jrnE5E2IgxCcD/fvEq7Qt/BTM4a1OmOi2fOLNdrtB/wztD0W1ggMKbVRVhWe
3fKG41UoGTcEh8LsuKzBaVWQLKgYaDkpnzOaj5aKbHeOJ0oU/DRnUS4MS/PZBTJT9Yat+w52dPMP
BPcMyjJdg1P2IWVtSZUVFEd+aoBxGjGYds3p6FA4Z1xXNu7KVNg9aB3IdG1ihN1ju0b0tOe+bb4A
mmmmSbJS6EsP53BXDiVDJq9Sxf1pzh+jum9JB58A7KrvryurdWj+BE7kkN3F8DR4wVNGGJJKb2L4
Wyio6d5DyW1O3icagAukNGm6aGkCeHuHGvlThhf32Eebxx25IfoOoItzvoEwEZ2wgkC7snLNZpCp
EUDlBKb7hHDFFqYSZzq0mAdxbU5OryKqtpG6pkTQk6oBQAurhSPLnE8KFCdlSdjRC+F+PPnG+0+d
0odWZdIuDv/AaW/aEfq7j1LZXjcGUAjXVLTpP5uEL/91LMF4nT0NQbVtVkTq5bbcbxV7kXHaAFgo
6m6T5uinhPIKW+dkRxIz4BYdyfVL9tpWWRW/TvgH6QYhKY+VYZMFI00rlLAsBr3SG77AjAX3Hwe+
HGcfJegCqCllazOJPJHw0YQLrGlz2XeCV6whW9E8FjYTo5Bl4EdIG4e2pU0F2IT4OL3T3YPlCaJL
kJge3Le9+Eexm1qGcFafk1toaQohM7nUo6Fakg0ut3O+j/E/fgAa18yVhwLbPJ1h/k08oU5yMoN9
cPhLkDJx5WZ4Z2jkEroRZR02YDMbZwNfZcJYE1F3aVjTX8ZLa2kuQ6glCzelnaK4b/I796Fg2h5R
a1nOv/q34wM5tbzXB0tjDjuGoX1FDBtq8INv2UOWQBXcvXHkfob45fHwWj74lQJ+7/3c3LhiKsvO
2Jg7oRNWLkgax6mTDfNLxlqOD0zdbpUazpvsTaTFpOvVsrQPWXIJJ8S3s1xIwEXNoTyjrQr3nC7t
KgJLnQen0+KNaOg4+exzgytMoaOz7BfQh7M7L6cpHzGulqtHBFQ87cIV6hV4mNY6I1TiYeA+5b8g
z21FgjC0RJAA3MzzcW4K6upKbPeFbZ38xzz3d3b0bXPZreiDZMyRb52uPmNoPQs38ZGVJpGVWBAa
YsY2DHQIAunODaCs+9MTxTEnvcRO8dm8OWjExrHsapK5Iz4i+dZcSuSq4zZa4ROneqhh+sjCgyqW
e8IhanJcv9O6wd1Y+aP5zTnPlxy4c1L+pPqt1Q07+s2Wd9Dza1O8Tmfoh7NvokAJf1CA4OggkD56
36+GrbkMcA8NcBQ12AqWYhGZunvzbrGA/RfUTTdFemaFX/dIEoMLGqGMfQm/cizcRYxEpxg0VVSo
sXLuXW0P08uuVX55O3QPBz6FEGMd/cGL6KDpNLBcYewDQFUQ7ECKQ5gLbcaaQCQqAKpxWvfxBgMW
Xqfr+m1JwLgOePeR6/YWJke2cyK/Gd0cUlNNLwCUUsec8obrrwNCQ7JHk5ypOVMZYUkyMt9aon13
4nuKf9abpWYggGsIi0zy09nDgq00hUgq/0Y5yBokJAkbtPHf4l8p1KE9XtzEfNFR2vaFaKCXSYoZ
CJxwK1EFOSU6HGOPOvw7Y3hNEEK4aELaZXlr8esFXXdfDStkmnDwJxKcp+V7EytVA9DYmaYUcuAA
7N5M/gHwU1ZVuOJvdZmS4fJ5ZvBgayVmjTS1hNZaJX0Nk+9k+TyxN5g91NUFGkQ1OD5SR1sjwimX
VyU3BkaEvw8Ym3XO5qy1lRpCSgp3RDA1aqx8AGCBszc+xmhXovFmNKZgUnxVzxGyCi9ZR8XavSV6
oWU4MgJIR7ag+/sVSsJ7XDc24xiYtl/ohHtLANbKt7JYLzr5SEQHlWSLpBqTPk82Iz2XrjCmIcJ9
WdDegL80VzIyHx/JrH5jyhL7jHbj/N05fPBiOfK5cqpN0P4XFMRfN6Iozr0E0FdrL71SqaAtAnvR
X2dSX5iCiErKaEssgT8pk8Mvr8eDBNG6f1gpFjY6LK7MwJTDan4tzy+hzJ+pe38mqM11xviPrKi9
46o+27ATND6yRoPGsRLASzUyULUyrduK4Q7xMDhwoAmxIz/JyOgEjpLL6D8wNB0HpoMPpxzD2Pc3
m8RTJTrvE5jrj0smxh4VOugEKsl/2DV0L6IGJojjcylIBqwLQSbExEeZn3QNx44gLM0kh0bATEsY
5GdB+b8Zw1lG1+xBeOJa8eHsZP0QTV7HSaJJah7j04OTln9I89n7dQqR+zaeYq5m0Ke+IrYT6JhC
a1U3HcxzjCy3XYfeCj43+cHbfUxcozSPVIsGu9ejbjU/uXDLdOLU9cr/ST9hInfaXEa/ARtI7Q1Z
5tLAbIfNz3VR5RiORHkH/Y6PoX5jH1lXdXFH7dRjUYbd7Hd7UzEBeiQcyDPGHIlGTdF0V/stCuVY
+F7LxGMYJDQ81pTXZ1VFRtCHAA+ny82UhaIcIacTdDxld9sNVjY1u2P5AAIDVnnKjyCv5eadFvdV
VZktRWLOc9NKDNhhEhRbnK2AkzJGy+bQClGYcyLqs53g8cdLhLUdgV0caNdZ+/3BUpPyYd/2qn0K
BzK2zmbGSdM0Nc5//CdxgxLFMxz1gZWmV2xnxfY7anvOXs/LgrYzUsuM8ARJmGzRVGI9ngWbQfp/
yHbeC8cEagtWWLxVI3UHGntjNYrgqH+D5n9aIPfQweVvXw1NBUctwfaQTUQix3pjYBpvwz7EWUj4
VQynTl2fwhMgYY5iZ9lvtLO6FBU3+x3G1n6fSosA+0B5F97zbSiIRu1Av8jRbNmmzTtcsrUF/m5o
WE5lVSLjKwtUgQA0R+9hHdkC0JcFbyL+6DU/SxKoLfBmwKGqj53xBi8KrMYVOxG38b0QsobG4lGl
+NS79qsoRnTdMApb/M7XVpj0BCijJTsI5W7tH6GmCC8UPJV0GHF0xB8mRSkaKhpIewBeUHpqMpFu
tpgOjoU40kTXSpOusCVVRki41KPk+UnJ47z+V0yolhJ3ESFTJ2zVCHrV/wwAqE9OA2dr349acr2a
mD4VouR8djxyN64nC669ds7AKPdEbe0u36eLfFdUIUh4Q0FobQs2g5h1Tuf7UGj755NOw33WfCS6
wHavp9f1jYDJRs583nf9pP+gpLsEvjqgFQBB24K3VrRsyyBqFdj5d8H9VcF60XHebfyMXREzr+el
AKdOxTCQXviTEBKL4dP6GD5ofZR6zUlMFAZTJkow+F1Nk9SvgrlG8mJmApDlhwwzfCIOA00VGOYF
ec3VB1aqwYpaJwkelXec1sZE7JzAQaHKSqJ6JgtEa/iRlE/7curd4YYVb8zG/Pn6xwevA1hsVaFH
PaNS0GFwSAjmZJb8tJzjvWPGCf0OaA/iACiRumMEpXiPc33Mos7CSlCovak0mZMg/LPsraxnMdol
H/Yg77GymmmNUznFW7BKQzvA5HZvYXs9k+1H13ypgL2I8Eb4IJBQTA3/wg2th94e+fkQjGrZQnu4
WBbIi/7U6Fdcpe1pGhm92b5Pxf+f+FiP1ZeRZ8etgxFJKBMZygiBcmwQ5FArAda1jFxW68xTJ2pb
DzaL3FpnvxCA8lmvfQe+WsbY1RCsbXqmZ1O/YzCjS0GcwPmXpfxAqieUdQE6dK/Xe918hisHMnW3
jsb65dewKt3gRWiYIMfItQ8cE8m290qrPlzM++dmGV88/QeZEniNVL8u3VeRtAr3+AyUEPG083TQ
lOlrK4skS07Cswt+ovyCJv4rZBDS26IbzlHcQay+8/dm0VQsVyvnTeKMxNQ9SoRBB3NXTrzM+VV4
sgStIkpP3Gm5HGEc0fbbAPYariDCoMTg+1DruEI7XOMjT38McADnTCaFlxyfr2E1da3Zv+auqbh9
WMuVViGf/QD+PKLSHzh5iZEr4LOIoqSpljCLLqprnUQamFF05oFN304ehDLtLGm1v4Clq+kJTJVK
UBXLDJXnyw0kCpGHZW6sIVJTKo7Cl3eCwPXQgwdu4NgeOuHmN6tsp7aGFzcWJHta+SkMugCTXeKf
OMShb+Z/KMUCvNLlCKOjbOSS8ZjIoITGYcaWNl82m5mr87M8ZvQYkiZqhMisYMKKG8WjcTC+8DqC
cPdi3b8ztQ2QZ5LHgi26N97VoMJR4tralCY+HvpR6l1hZVXU/fhsPJFbOVQMFQD2D9TIbQy0TrbD
b8boi01gvy3X8hvbq1wsEYnOT6L7szeZe861KkTPDZtSAbkcGg1DBlmzq3G21z2wRCsfrHzFAyBD
iXDZoYFcLadXmsFRWIYdJNCOhcm4TT3L7SEV2nejPeCgACT3Skyivjn4dtVBxtuZTngs97HxEqa1
P1InNJ6aIw9HJUfbFFflYdl+ul2ZBeP+oLfGP4pHvtxXcn2qHMzBfZKpuV/RRuSET4yGXKVnB88F
dfvSsTmUxfXhznlzi3EXzxzJUjGQRNJRJEpE5mDk4LdGW1dTsmENr7YrqzaChS+Qh1EJ1jttRhs0
Zouc4UXdYUCrDNptcjdruTHUN/HQGkecyM42NcvJrXP9W/+rPSlHOSX6TDfKy7E4DgMfeZ8zbGv9
JgAw2KaoUuNS+F3EePOk5rTSNDdbF0r+6LYIgR75riyG5NAZEnrE1pI264wZO1PL6g87kIIdZun6
dxG+44fttrNVzjbDbZ03zDI/+AzDJ3r6GK+NWpWqHEt7G9rtg7snmEgg9NC6X/OW6rrjr9aylIL1
U22tLzfOtB0bkN7bafwdigHaiE49dS+5mgSi7/huVOPINyCKgiLQCPRkpCGkr+2JeJoC7LNYHYnH
lZLx3tHYb5JH3L9YdLGvROMXSl1QV7HisvcT9ukSqGrAQo3+dFZfwqCXjS4FdalRO1b2s4DaTx4U
9zV1HEeIj85GMqB6MzU0IudRRYWHIn3nLjDy+5k2VqoCrR2o2LDAdhu2vfrVO12my7AgPudctAyA
miIWFxzONktIWOEArsscFSqux7OJBuETL9gsoeqEkSRHwnevLIXSiYlfOvJySUz7m41HSqqQsGlF
uiKbELaGlDiaDkuHfCe8VetYflz3Z0Ftf4P7J+mpv/xDRf6kZo903PRE2PBIOZwWiPq5qq5CIY0R
XaNBaRfFOiOY9q/LxWOX59oZiSQXfOdTWfYdx8dCdgP9yBSH9Xw/Wfe7LxknTbOnQMNxhVYibon1
0IbhjHdoe6COuHdRv14F4XxxB+/I5StEE4UFv8fUrhxWgNUcNNXXAAx4L1+Fu/VqJd8GIW7SKGz9
1fv/dJO416JwC5UsmvSK6eM3W+aoJlFaJ1joZ8gmMWHmWoEl4QnL7dMInXZQf0meQYR8/vGYzBrN
TPzx9VgmW7IEU4Kl7Jzi8p0QPxbAmhABsq8xjmE9vndeBM6krcxo3irxdngpR93PhnUOFV9ev23T
juQBbpmUg5Fl0RRBg2agsaYUNoHQkf+cEAHMWgXJPC8FZXIVTzMUCOZPlbYtm5Sr1wjFSErMaVXH
VMnd/XNgN1M3tNqm3DfHSraofHXpg19W4wIOAyjSmIPZIjo+2cSFitIuiTbn52JJauFjPfmx9+GL
VoQtMDj7UxGP5refivu5S0PAT9Tpwr/+W5RUSklk//n7zgR1t5CglIm6pE2G8IVvK1wejEtI84ZX
UwHSswAZnlUxX0Hr77Y6iHrqRN6WlEZg+xnfKk5HuH1+ggM4WYg9g83erjUG4qSqWuKTT9shsg5h
vrpz/aAky77Vmq3c6cqWn8V4f4HuArYEEPMUyYpZHg8d7OhIVmiaIU7bdR7+iPZV75WBB6JutA3M
QhTT+sTsdBRRT3KATkTToWTg9iZB7He14fXUap7i2w1j2zDTDjqloDsf6LCrmkIAvPmNStBft6wQ
wrnclDhW34dthRge6OaAHFutgec73i00Swlndx0wXhPCTUGEsI/5GwXZQn+zxMh1P2R6NJo82Ro0
aSlQfhIDUNMe7eY8XCaI9QZrOXJ+fNvA/1kJKbDzxgmEbGRjXS9XlF5TLoseaCl+7md2Y7znj/e0
fc0CINPBAIENwcmx8Ze2tBMWUwkvrCBe1TVfzuZ7TFO2JTX73iJaSu5wMkKdBeyiUCv6Jg9JzoPI
Fm/6upDqF2NiJ1a9CSqBy6n6Wd8TWI6x1VpfmBKsodQhKYd+/53tKKNO1oaRuWg0TZ1pwwHg+qOm
CVBnWJoxU6tbWURSNlpuklr+Pf9p0DPfbNnCJTNTaaSX76gPxLzsDuiN0vT9UmlDX7ANUSmgU7gH
5sgs5GDv38BbLqjoBVgq1X9CzwBmpowhE6c0CWXH8Fle3UIXsDkrZ+eb0YvUqunyjUTGhY7Tws3M
wpdKAALSQKXLAKgzqQGkN3pYhbyFkbje02h3/DUUg+PN65wtDEn7cyvmduRK6KTt3Ocsgq0N+OHe
jeFD3jHgYo1ikpStStKmgy8dQbz47doZz6YgLXd3AjHKWFlY2o813eRUdz0UQsJNAI4ijGAlOH4W
goXT9TAWINAGf7xMKfTpim8YUf+hgdw1p5vLYlK24DdVziZpWGClDQgZx2zOgw59po8ze0NSRRcK
bKwQhZimYoIVAmKVEYbTchaZQTorw9oyeE/yYmd7uvw19Pprl7pErtHfErW8QOIX7X12fneM3uYu
LsmhMSKuMeqW4CIpDlgNu4VolLz+qT0cOwcFz0KZcT34l45Pf/LV1X0cVsA1MKOmCoiTr0SMs/7P
rhdGwA6H7i6HaIueYv6UeNdGhj9i7Qq488mY2mMnCyfdXnQ9G3bAtcufW10PTNcIriolpfKvcbM7
icxb2ePWTaoOugXkU8DrrE7Sa0xH5c0/7W8dczf5B8s/+yXxS294anfluRE4E8yaAlCMVt7iX2dB
ojFYyuqcepPlhQSgR+kxudpUIamRfhZtXeNl3l7M1+J2xTqe6ZbMH0kRUClXha+iIqXlx432ONI/
BOiJ6ADZOSnsngl1EhbwwZkbePZ7+SoW1K9LYIdFrbyXDwHuSPHT5Bi5PDb+Y2TSzbduh2dqn2UA
3uZ634Czio2jfpA0fmn7plHDHOZzQ94wC+jE9h2oOUNIwRI5ErjYRlLP2yi4pO1I4IgIDfnyILv+
ZJGuZTQDW1BKsW25gfFSv8VFfxpWNjR3kLRcJrgrVyAUolmfZYXu7vxIPDS4/jtsK4eTbKEiPIAr
vzMi4A+lxFb8E14/lzGg2Yvdavr8qhOJ+dL/mRwS7ZrARidAvGB8dzmh93Z+kEPe0qpOALYYj2NO
jhSlVCCi+Vekflcqz1TVpqh3ybtb5p4L89Q61Cj4yUNCqv3/jAmIQtfm4TtywItHQse18voFtUoY
3PS8pmOHczpYQAco9usyFYsPYAhjWUy8f4ydwnlej6aZbNMOOCL3oGPhGwDlSwpML29G6UnOQ2Qp
rcaWzWL4o8ffAsQ68jNw8q3V8w0vkMq8LQrFCct6GpQAOAfxZa4Igo4Vhdo4eZxnZ5QItvcLDQH/
kfNkbU7Qc9Mx3mCfJTDo6fBA7YicDWTZzOqLmmT/0F+epYo8+Nh4OYIVBbOeds9udoLn4pQ7o9Ca
R5rT+bwbjC3poC3tjB7c8oyC8XED4GueOCdeHGsOagoHZpWjbZD0ehK0FS9VQ2TzEmwSPfTpmy0f
jgWrsu7xZoEJPy4O9pR+IHi16FKzlCq/5PnKXoMD3Ju6eB2aiiO574FGbZAeWjXzru24GzU1Jyjh
WE8p/NG0G/MXttFIDFCZDCscEh5hpiWb8+9O57PZWkG29j9G/SMuziUGnpLakXRIrvvjU4PfhEYi
OFJ2n/CYcXQPnI0eV9usb3JJoKFQePw0EHeayE/bnCGFL5uDmsRccBwYG+BaDTn0pRuB9ggibSGw
wJPjyJVpMljlpbeerX+OlEPQY+gB9ejhKUWYunQpcLqJ3OjVhKT0UJJ248cXz2B0iuYBf2dVjqTq
zZ2MsawwoOqt6qx85ytDaWRnlAxSey6WkHcOAdBTpc1YSMVUCwlGpU7TmCe+gghrcEIXkZPqo0Sv
R5c+zHjaqGVXZ9BwVHSozHRdwRR6Q/PZJbEF8cfvLW5DHPGFZsr44tjrQqE9vh2+4tb57GReSARb
BaNEC1IHuDs0J2xXX6EPqG9J1KgYNrrc3myvAD7p2ZkuJHp2yLtfwpy8wqR4WDZYkcFXvifZ8/f/
oRi8wJODu83+BZ36/PZQIR+UBuz8sJyc5o97lXgOemZOrFGkK9WolaiG+ifNYFD4rflpuXSKTAqW
5s9D8bIeMoUC+GwdoI1YA72vrnkVKh7Nq710uzNPBlapT1HN72QHw1yh9xbs9Zv7Pgw4cb6b/wGt
shUgYz7qBJpdMdvE1x9/fWPL+rkHv7Mj+tU956EPVKl06uxjM4vENPxm1sTU6lgKb77AscsMnNAe
n+6zbVSONKHNvP9QPYLct79AtXfBwKYBjjhx/9D6vOf5hoihBCdXDLa/PoKRuTjqW0bf+hICmeBr
cZUI/4FhMoKuCsdMYBP0f6cxcoMHcSsZpu3cLRthAkr0ul2jxo36v97VjRp7gD8np21Odf9hvi+Z
Y+mXVjjvHpo5xIEed5BGeE3YhOp+H8r2xkGlrc9Tr1g40G279g3v2+tIXjhOsH5WPwoxoojGEkm8
YGYUMHkrCPW0HPBQVb2+W4pDhfsf87vxoxFvHf3TIEzxH7oRc7na/V7BRAdriXD+Dhf/zEPy1H4N
1Qydu4CmPGhiwetCyI/XDsXouq3/I8Qmaw7FUTo4nywv73mXERYmTnisVKX8WTLYHNGwnGOuyOtz
SfMSmVcJMIxnzW0GmCdyPMBPbjpt3R18WZaUZlhnsS5xvPv0041WTWf+uDi4eO39y9dR2rsJqsss
MxNJChCznB+DqBT7AMbfHCW2fed4U799tMKsMDHqZdYAbheyE/veyW6tWP/rk3pPhnPCELSC7Pr2
80q0nTttlN0KzpHXueeukUuqxosM/fK+l1nFhWRh1EeR9iLTaRnDyxUkDUfmZDmfnshUT8JQkU4x
7wm/VVdya7ZO/TVimiKS0anFrjTP8Wu1Gv+6S5Kqx/KOMFaj7KX34ymGudaHvS3t9wDOznXzg0jp
Hof35F/2bKVlvzPvoGqnaz525GxEln4DvF8+XF3v4rcdfy9FThcjGjYFL86ObXZTbmBpkQgMTLEK
s2ODJ0Pk0dscgZNsS3llQe8e8kfpv40MzhHDS61JcwzTinAiT/eGfHtexx+mjI6ufW+6M4ibXq8I
aYVvKPyUfeDTX4cu6KgRid8JsHe5tLCLMPwzgO+UBv/F5A04qBbcTRAKsNVZ/ib26/aXUWDIkyAO
PG1LWkxuwTpJe4wshe9wr0oCYLffNq/TnMENJrsbSaH/lfFhQsyIFGXCsbRy793wWy05kDXePSIf
Td9ew+g1N4ifdZLzOW9o79zJZcO4iGCas/SwUBjxfebpYzj0Hz9mmrdFQxFIXJjF6NQbjQqCoxEH
fyJUVbZMnCbeek6o5ArgllW062fqLWbD39yhuVTOWrw51vRDzkyxgzXnedHn1Z4SE6oUiE8RCLw8
TVA8igLzC8Lh+kCD6ptiwYDlVEniM9mWJuBooC4LyaI4N5lTIR/aNoJVIurETpV633l0o1sWidq7
kHMPAzUixv8wXPfHDjIPCKd62SWKF8J58ZV4DNcl5NDLi1DuU5ijj/WLvfU6T+pd0UzqVXZ6i/S5
rI559AHPy2eg45c3MMvwjQXv7htpYrpahP8J8j0BYZzOipc4Ke9YfWeSnCndOoTNektALzRNa5eQ
fDEc4ZJyg2Uzp5natEgcIH3pB60a00eFW12ZZMwfd1lFuVsp1GjsLJfu0qK7fyT6rEe+x/7hHcsT
NzKISNzTWTpELF+qCWsu4B+oYtvwU5B1GqugySGobqSEMACYqfsTNjt2MR972uEKV8FBD0bLNLVn
lAZLCtfw0gwm69GvoO11Ear3seOH282fG20k9GevPA7FQxvP78gIIQepeQM+SI2tyoE8tSEHRWs/
aIrVdKoAZqGOeiDkxywGSCjMs+WnWkQpCJ6lCT1VVPBI4cHBywktILq7Kt+PH7CJSmtoJz+aj9J+
JZvr+kIuvMtFCxqpioeWFBjkevHvuC2EjaaxgX9Sd90oFbxSIyfzYOycAo7HMahtM0YgA4C1sI6x
8yozGlYJz/zTB6j4OkAUKyfvb4P4BaDfctF0KrxFC8NmEiCHUTgFcbL7lDWkj57aIwJ80aCkalLO
EpbfEB63pwiQbWlACdTSFU7I8f4D02gGSLY3xkSwb3soZH+wAjQBBxE3T4ihvu78FR/9i/PhPHdr
lDkBtCy6hRNDnbbCD5zFBPtyVmAIAUN1a32MYen1+jT7uyDp+d2IQIP9szgiKk1/FgnOBRfoPjjl
0u/weZ6W7MWzUP7+zXkKwSuBE+6pyv42qnhpPHY0IdJC6BUI0I7uyT9393KIg29H7UFDfM/XNJl8
pbr5FlE3fuQLIzhDXJZymqDtZAUH4cXv17zjMrj/UcFtSm6JA4a9VxyXRoxy07v0YtQNQR1uhe6h
rhDegBRY1jiokh96cnoylf6bYASsgA9pmezqQlVDWI6gOvKM38hOGY9KhRdG59yXiAo8kwbq9VlK
TQXPx/VQAA95cNgVWfwYW2IvlE/QIm4cRb7o6t563DjZTs3+QWvVsiEAh2d5vzOOweJHcdHqOAPM
bxv8w09bzPqoPTgvRHcQohhF8N4+g9R3qKqRZ6A1Y7GeYob7i/laWijp5n4lMtbyKy9sFdD0FuZY
uqo6arnhOroguKMH0Eiifab5hJoEsLEUQqm2P4lqaGES1BCvX+QY4jXUeME9XQfcNzP/4icrEc5I
aRG9+Lil8qTbj1Rbeit1MWxjF1WtdGlp3uhDmFQZbWrsnqghnfVeq5VVhAGOqzX8uBm0/OIzri9g
6rPjrLBls6AtD97EFBmoUXHT8U3zBnmI8alA1uWXvrePaxYINO4MpoVCQGFot2mLFRh6WlX39OPq
+6oCOXOKTUcP5odJuaed7EZIOLfdhzk24dxQpZurLTFzFrvBNhsbDsMxo9VSyRioRobczq80KvgG
JFBw0Cfi0BfJ5nkbrpfH4gSneIP2qaM2TSC7zyyKknaMI1+c9v0VyeGPL1vO+FQC9HDPyb3OwFNc
9zzuNMb1RfDnoCLSTCfTOUjcOLtoQcf3l0MCttYhzJ1TXvOPVQ6e/Gz4eEyOTWWflnasmF0gyfns
uuuYqiyf7h5p5Isn4YwJFbyosATUdMIybK1J+ZZ4G331+i9pFg1CKdWBYi1LgxdW2SIQI27ktbtG
KrZW1BuMcA5iIqtwSQ6GgOlI8ugMU0g2qNUcRBgdjcrS0gFZ6hV3dLgGKi+NSjK0TWzvtDh63HiR
sdwOwCSHtVdZY1E34p5zR70tdAxh0hOBQ/EbfV11gvUx6U2VadRMGSCSx/zZsMfh9IaLpe0rElL4
3lZ1ID7tD3vqpxv6a6BZSt9wyLJhtEQ0+UliABlB6gJ6jMN/DdAnFyTt6869je3OW2P1HtfvkHP4
jjXCUwS06CQDdEZDJxLQsYjwe9KWt149H18uluYJrDGERRkQ+jdzm0766wlgb+niUi/LN6CuiBiB
QuZeTvz+ELOWTKpEo7NWq9PAtgV64/R0HDvqjDUlhhWXlZeqN+s8fJ/Q0nroerUFSmLt10b9f+Km
m5R3/pVzIwNeVaorOAVUal+qC+GdwCwvaRY3BalnTUnFVzhLUAfga8XE1P8suaM2NC1ym7CEr7D1
jHiifsS7woMR0GrJ/LEsWUFoUNqJUu8xxBZ8L2wOlkFoQebM+4oUrsUZvOH/ysh/tOInKJQvEcBz
kwke9gdZ7FycpRD1shNaBQR36DHjp46Ye+H+R2irSg0vHQWiaUGPrGr+7rGVbGxIw4aoNq83Dhwk
EvbRlNUNwsnHeYgmfTMS3jA9jXvGo59bLZSDEBQ2Sked5BKMFny8Zll2a761VX1kkqe7USlZXaDd
qUV/VAjKWzowENigszHdZ8Fho90XcbUwnRMi19XVy/wbZVNuB49rXVDD3uwW2KGbYuYqL5S6iQMB
uI5SO+ZTJshPnE7Gv8e6hjcKjkTGYuQ0VIM1Lg9avc3pg6+Z5wlqy7OCVMkmQHg17YoHuuKKTPcq
ZRtkldZHoGxCbpSc614DcTBXCiutlT87sTi79DOJ3hXXHvFJaLmY+skYp4TE1uXpEkw3xZuBd1tx
8uHhX1f9dY6O50lGu+JIxR0sn3iza/kddJyPfYY48rRdYmiygz5RA9lW3oslqjjKniz0X3IUKnfd
L9EKvgRweDVixh8sUTmLI13bIyMYqkcgjgCXWSbkKAWJiw3oInc1EjPbuSjHVkFhu0stwpm7nT64
g3sMfdByJFOG55JHz/1AHh54krplTfurLHt7JAFFlr9Gi5HKwcQ6h7TLwfa5NRBSyB64Qls71TkU
lGzDTwxAA0ewn9orHVdq+hpSkLddGhPOlD5HeucC6Xlyp9erShZ2f53aSIngFlOFDQ/hYD6BcMqE
rEfz8joNo1V/jMDyOv/+GlhB6N6TwfUqPsdNs0ocaTygFegLPOaUnBZ2AC9jUzyCAwP4zYur5Y0W
EVa+zSD0vukL/ZiayIjMy+RKZ+8xfCGnShC/wevszql+1tr07zFwCft+RNeuG5VISYrYHIhcNpjy
W2LIlxvf5+AiDZhJjSwGKR/0Zfo4lV1qgnqYukunhvK2sHnLa12bYKY1azq2yGkyAcYg/VqOdTuU
AXxdjxHWVtCD9eWsR9AJo9EpXF+EvDwS4zTTuAWuzK0xmSYGipiVCG0DT/XzMb7n/U2uLFumNYM5
mwaMKMxzICzKmcyUGW5vq1luzXSTrJ0wXH20n0/Vi/O6yI7bS8i7edcgQ7Blm48WpBzexHX/76ie
Hj2894mXyuZ2V3GIlRwNPra++cGNshgu7fT+/6tpHOhDQSDqUwAaeWfd36BAeeuSpJiH7cuLBTdm
DUgfZY/l0x3q625t5is1rKbI/VoykvC+vGbSsoiEZs4ydOKmzoCzmpOadqIjtzxTyFzcnhiFWa6o
ngEHdW7bigcYoIBpcKFFu7Ma2Io+1V4mZlIxLK3l1ddH84t69E699HAVRu7L4ErhldAZsX5eLU8t
/cioZ2l1zpGBPOIl5sOFCBLTgOrNcWUcsT80VXsrt0OF231Z544i/GZ2APItzitL+jo+Epg6+RtB
3VaSHBBgsrhPs9sstEKWfXAWWvW9XRZZMh++Xbaa3YXn9yqJAelyydi0kmS1TPMwsMBIlBLnugzs
aLq0ImwI1yw1yQ+iDzrhEsQ/fNYIn8SzWOHOWN3Y/gqkPnN8jLYyGx42gN3gBC8NBQ6cwIcPqeJq
b2MFM95MzfmUpS9TJ7/Mul4ONrNjuLRNOCFNbsm3nxo+GyG72Ud1rKTStS60jOlrxcAZJSF47FwU
FLyQhoj6MtCuLKoszidcBhE2wH1qZzTtKV7zLbeRqNSZgQz4bCi5oiON7swswF6NC9ey72Mc1pwe
w0HUj0KljLTmztA0/mIAh70xhFUXvLmRcXwAJPEtZ43i5ugm6PcxfpL3HoJC8y+bMssLq1UPl8f9
YcdUWsLVKHOjaA5Y72Zfv7XdGZYsN7YRlVIPPDyJzo5nmsaFoNCZZe6TBzXX3w17H7sxLd7vwsn/
bDF2h5XA0Lq4Y5KHMbDeyVbL1gDWcRcB6SKiCmSin2hGQokVJNDOOVBqoAgjTVSoycdWQUn1Wji7
DZym9rUgIXrx05ieCKk5Iqd7yHt4NxjvcfD9ogs9kZXMQoHeEzaiTxx3S8AMlI/EjJ2j8uhQPbEO
fs7XjsPrVpQ02iKEx6pLktaT6/W/hMIY4sCoFGCB7xChhkLnQkqmOBbEaJyq3U4fOusZl+Jv287E
LwF2YkrmL26vcjgasYRgtIhfjCoqMCyAtynbwOIeDvnTlakU1hCn8zHTm6dAQw4XrQaseRLG12EQ
qeGjsIZymwBeTbQsywyMLswmoLpJNjUW5vffJs8L8w+KJBYF5VK5eg/iIM6UhRHMYNruJ7/dIR++
H/SnXeQ6sGBWo4u8srihjoVwGX/vMe7A2JjeYEfeClKou49k59HjYD9WldGjWRfsPN6xEFtmO7cO
34nJbiTZcQh/CA5e42ws5m29cwwaSzHGBzoAJpwT0LrEFrxcv1NorA2GQRdu4vbDamVy9waZKxws
3r2pSghq0C7XBCjjPrielkkKoMBTVwsUxnPpf3eMV3QDOag+6aScj1A2x7RVrLkINxyPJTre/mkR
yLhh8E+lctWD6FrzLR3td3KkmyU6QPbU0AoDTt1+jtqS12YJ5jblCtvul/Bl0ouJ7ZP8gDJdDv4i
/gISE8OQqR8sEp9wnTCu4CtI/tGs9h4RwLlA1w8mAW4BdE6tykOzEeEdsczsuI91aGaFe22lwsCh
5ytALRM47aT6x1x0Wb+MqAnYzOEpdkigPPOLIJA2UN4Ye0IiCaAr+Kqu7rJHD+qzrry5wtsPXxd9
hCt6b+iv5gsPaXAlqspGX909rp3fmaiKDXyc5JKBF+wyZeCkI2RAa1mY9MSISlyZffsWlDLjT6Qs
teqZaJRoN3nJRxa1glukozqqLpp5uPNiKLwXOMl4JWBP5GLTAwz2bh3yhtWJ2Y42bE+jpLHNQL5m
kSSKMS+TyKvx99M1XxxPjcE3zKmGql/srpLEAZ0DZXrQj2Qr76dZ/VmJtJb7B2P33uzU6yowLeoA
mTwQMw/u7gQHxyzEypHZpu+cL04gzpmmMXr+m7GgJuEhQRiPvS7iCmHQbeksNY0EZp1zjVFcLubT
WBwcJChf+ZDbyV/tH01Eb+Kpe34YI+K87DbXUqlD1kXwdSr0wsqMeyeITBm+3bwwBFPaJ6Y4ZKJU
6+xge1cwBBA6wCEARRjygYXkNpwqQ9cWstp3ehDR/iV8RWhTMb36qh1Ign9CLthFKEFOcvLKC5O5
y1MVioIs9+zEc25u4QpW3BIS2Bf5QXLiBTDHtBE1huT98qB/VxzWnjHnRra5CxbEjfvtXRbIaGmp
5l1QXytUgMSpR3lUVuHbr6UtT+rQjPjcJgw+xQUxpRTH2X+gZ9UPzXIQ7iE2xriTxD3l2L/2Yp+V
+x9URNwL/Lj3u9UfXsj4B2vrsm3csz0Dk3WCdrE2wQneiN6BtAftlGnOoCaPE+3uwBt8EcKKh6Gq
TilJLMpIqJ9AQD85/A7et9fAqwpZ3XJh0w3Tw+Vjgh1jiGxJqUUZfB1/xYAKRRxp5alQ7FRFoUTE
ACIcT1sA80hXq6VcxbpwiZjROgok6q9macrUN19fyeB/RDrYqFyRUhov2p4FqwbXvq+R8i9nOmCi
K77A9uIV5wTrHC040C9SReE5C8W3LtVjETuHRRH60/DPYzvNie8bwCU6ScsOkOccr8whDWSs32X3
q+Dowu+6GotiR8Nl7vNItluSrL6kDMj1WS6XpN7s+ohN/UBsAa3WjLTFiCItRbo2eZjndHJLVwTJ
TYPoinAZ9LFK99YYAU/4NaiwycRhl0ciQK3q9Bxz8S2fgUMw5jHCUVVthZY1ZUzf3aj2sdqiqV2x
/WlObvt6EA8nE6A4Or70mZ1BVcvrqm/z23nc1ca+1ulA//8GyVanamx5Loap5BqjL32nzoLfysPh
M4imAJ6M/7rO2jUWkeDlXsgt/YAHRqKAiV+2EqlG70hXLp5Vqi4oPVKx0et8KcguWAq/CEMGfcVk
OGiXtLUrI+lgPeQAEvNK1CdQbwO8I5njfOAqCM/VjQS3GsUDLjy4ZfdHK/oSJc198jZoESRhvdA0
6XByIVC1F3Z0bkdYjpsjpKHe7bLS9TozTRvDqmjHdOVbHhiY1irDc5zZOTHG492z5Vp4rf2+olH2
J/6uxz/3fsZmOYh0o3LTbUOB4pC8aF/wxIdVi/g3I98ChnER6uCYQDGmIA46h0LkeyN88H6l2Svf
ssP9YcN8Klz8tXmKIWrup9wQN7PCTrYnQEQQop3bGYxbO1DaJ6AhS6i0nJvkks/ScocTcdMgx9fr
2cL+qaFVt70YcPkRCZ2wC3lWxtgGfBsrFlKAV5TlotilJUOIU2QuVJt7NF/RIa0EK9oUgjSJ1Tyx
THYp+lhmZ4iTzzLjW5Rj8hDkn4SuVE9rwzS4e2AA4MzDHLpF74mBXPa4q+pk/NyZcINkooMHx9+L
jsj39BAugon3DUR+00KnpFxOCVtMMd+2b5jilSrMP+zM7/cW+r34yGUqis+noFcMJ6ZxeulAS8BN
SwPkHvlnnEFZLtN88ysw4Tobax2WYOnb4IBOBBGYIlh/mAp1++xoRCfICZnrIIW/wRPh8tYF9tp6
jBcD5UVWaNdXGDwiKc1Az+RNYBXIxhBP7bV2Cmv/UjjYZSfNdMH4RL9bs2sywm/2m9pw+soNBrZn
IPNlc//koLKMtUaqVzY3dffno17mAWvHwMDhupMLFZ8QReNZlpuGatdiAz3buKTVAMEp4T5E2uOW
x5h2M+EniEW1nW1V507lJJGAi7uITzlRMKdzR6dGRSl+DXV6MpdDsbRcQIIZFNbFUpicgpx2KYKM
gSmG+vmr75BnSY0R/9sJ5LPNNp6vFq1MNN4LaFRsFraSzvVPXlke7lFZD9UKlF+W2yHpQZkzTaB+
hns8zlMeELlPKfp787L2sHjgTdlFUzk4XsgruP6cYsgrn8Mw3TG6J3XVQRye0bO3nHOUrWugxX/3
990hqy7UmkX9YIEWjdBxucEF1Rz6bBrqL2g9/ifI8yEGdK6Yh3ekEQux27x1Ymwj3wwbUdfHnfG1
yl8l/S5+Pff34/1p9PNyO4tJ0ve0hvnvB+639FQB3byF0KPsm1WFPRPPRjs9Rty01ytDF0ZgeH4g
dFNNx/teANO4fYMPXaY6bBnto3F/d0L+wmLdfjd5j1+dkvzmfgdIo313LUV0iUG9te6cJe9F/mrL
te9Y3Qg/a3W2Hyj7bmNaiS7zTaE6yCYBH7NjYyXY57g3MoUl9XpaAnzMfYLt5hUo9yC7u+ZKH0Sm
RMX4sZqg2/G+W2lF0zRSGjtoI5OZI8jR72RuWVkQ1ECMAHyysvNNwRSClr890S+C983qIKtzO2D/
ab5e5hKTuRiLDh+vAbM/bt+ZfFE2KKGgbRiaZuR73OF3WXQVlrWeY1hqVXG0phWXixnRqM5r+EiZ
2lma3NLdZ2ZvWb/emlEZiEv8bjq1dA3TX88uJjYW9stWdziFD3ERMV6gFH5QdlV3P6P4gY33JV1U
bqoTxx5cPrAQwsqzHln6n4yR1lacocmwDtAOXZYkgoqE5MwwwTszPc1S91A0D4nY5lqZDLRPubNj
8C6RXLu1TwRRMusdWcutm7ZBWFz63P8GjEN+NCfBxlJi87B0OWAPQ6uuaK4QpA07eDwao42jShVt
PPx61kmXmuwA81JFuwTorTofqWtun3d/Z6+xkoJpg8iVFdURT+nKQwi1ZvmKAZzY0aRYLTVQO57e
IyvaecSbaI6pyXC1asPKwTStjmwMDU/TsU5sSgoxdltHSuxQfDCExn+2jMMCI6xtPGKcrJHqMRPX
BBtWATyxkFDv8CqnZc+mS8n9lBupaepldiNiL39GA8dUOufXyekIJ6sBFmnY+JJYztUfbpVk5ssc
uNOd7R/1ygITDeVG8cOvW7ptyJMKbunCPfbL+api8Rq5aIr/bxDqYrlUwUvMR7nw7Qjrr4xLuui9
AWKqk31Of9yqf6ukOzlA4jXv0pHGMHFyKquVGZ70kr7Dnt/ExmiR4qOahyYkT22l7CFnOX9PQ3hM
DLmxysUMn8+fBsd03u0WgzHfvh5CtCwcuj8L1OKDBaJPDEiDqYlBarG/RWQr+OI2K/+L0g9c9l2A
gxmFd1ASF8rC3omSmfOuKtKJRDqIPbyYIVNeaaUREFayGpt5B5ElsQQYBh1RWEEh9N5b7DRzd4jV
G20ZVQHpvAQ5m/p+U/PUf+U7J8MCP2QEs1kdvIk55uIjWVDjJC0RIY8uYulxRgVSFUlnpUMxExlm
zfifzNrwQlPDPKfiAvbP+tFwHGKcMpXFEt4FYu9nPV01fQa1GGf33uZ3fQ2VhueIeEVUKvzoiS2b
N7Q1sNaI8OksSxwnCivh7erfNM+i5m+90e8NI/0iZUQTVLoQrLNwPI+kKD5IBYvkSovpnZ58Fd2/
/jJVk+2VHhJLRR2Gn78pGsava11nWdemMIknIGgh3U2+bDcUjk55Ws8vPbhwGyKnXXzBt9MYyLFC
0SH1LNVHLWK5au5gK6paNbI1Roh3tuDSMgnWEdObTnVCbD3SRC2rDlhQqBOT6+FR67E6bv2m/+Ac
sZM3hQdNvFTDVnXTCL0eWLzcuQWUi25/eC5xO3kDneSD55h3XI+ZHir7Txb2/aPlz6tsG+7qVbx0
cZ1/u6bnBtFnFQoR7PpxoKNP1OrmrJFBK2+VECQ2jfASdDNam5rXEsMWT39wq2X7NIF1/v9dgXAA
sjMj2hjxZUS8uqNz7WTVbiLt9Ev5HWSuMd6NdkAxrfpNbokkSyA72NXJxXTHFTo9LZ9no1qUy7a6
HB6gC8TOBSKIzR7cs4lVzuuLsGydI3bjDKdYhpKf1EM558UugC5hjkWqfh2MifW6vD8v/5hsaDr1
angsH6+0xW7DGtQpwMr6G2TzkJ/VQWuUKwo6/czvQiKJ8Dq25qQyFYmB8kflTmwxKipOv7WR0cZX
tYzvgMYAhAHH+OPOWxWkhrPMt4E1rhu5k4Bhg2VOBVOmN8SQ3ZhtFXj/btGQEphsPnW7axVdzBzt
mIxW+diMiplcbyAAaIoSTSJnLqVbP/sEHvuuZH4FHvRJcA9VZB0vaItA8wxDgmlePIkWXURn85qY
cj4DccjewK0jjyQIJUK/YQ4fwJiLXKRKC5I2aj0tXOzPItFQw7EyyRVnyDyH6GRiX1grxWPf787Z
jM5i1ku4TnZLc9OnjSBq/9J3Imco8TuFclQ6gAAreUrhai6rf4+FGDlOvSZPOaem6XnyODIpaa50
4l8tzCcXMtwSByX0Ae5MqjIqqNVDrAUhC9hcemWj/KAkgI6GVMBAEukh2Qp2AHIvJtlwxh72sAZI
hQ66Su++0M0IDtdLUP7T4fxu4BB7AUS48pRD+N+TvLHmAz846CjgSnukBvnFsW1hC3axDiFHeUv0
BCK9B6oXdV1lJZdu7s5u3y8V1vRzxWNyhi7jQBSV5CybAsmd6nO6ej4QRkTmd46tmVXco/9zbwM1
qhtGMmDBFROXQNaEoqykxK0KgOnll6V5VavnEacVKVtztERwD8Wqd7xWN+PhDc4JiQJhgDZ/9sh+
NP1vxiDU6IticwbOWKh+WriZpfVyd9LX/UrzNbPfQ45rAMr1s0htq/I5nm7viwrT0uA+86T0urGm
BJ2+VHG/k+Re8pBg4ZGw61I6gFPMiVNGZIv1Niidybj7AaRm44q5RfkLW7iRWUY4W/RuQCs633BK
eFzU4HNTRSdYz6Wk+7xi0mOkrEwaCrcoRCWC0++k9Wq3vHR4RqwMyJGfih11JayOmiOcoO4EERCr
mNInKVWO2ZpWNJaUhzv7HSaoftgm4/tWiw5Lotw0Z6AgcJ5p4lFAtHZpBSoaqwkjA8cDEmhPS37J
ghYuUDXjkoz9IkoCyssfGKuA0nhgFybG0NGcbBKiuIIYvWltrYTiHhEbkfckmMS774X5JecV06ys
uoH7uFL6HGRq902QTBAGtsKbt5h9tKGCDut0A0m9hQWt2W8mYh7TlZflVYPtOFJFTPPdzy9CRQXX
GVFcCuIxY7rzkObUNjW7rwZdyWe7v18A6ek+vk9VyVbN7zQVafivF44XXZTzuDPxnAem9a/mo+4N
+t6e4/EewXsDT0gXtJlJXo5zEjiQkDDsIYYEb6ODa/H1nA5mPgrIUFn+kNesO6Cfr+JFJBXGUDZ9
JizXnOlfRQsvTAKPzkcUJ7AQo9Mx9GEBcwISHXXUDzK4huhILs0jTtJrZ33Y1B9hEeWrLieaitm2
rHH17toh9epQpoRj7PRMOgTMuBSmpMsWfE6DZz2ifnOav3Qa1Sd7r6jh0XC99xMDzvDTnPpdzcUU
m1EyVgKS8kAUXkKB9FWHQpiWSJl5iDHhm8KEsI7OLoYv5QtVy4NB6FRffd7P1lfU6rdyeP2cIeFi
smzDesXxnjz5Wu8qKuXsph6KetCcuHBTBrjnxOUP9qyVLIGH+dETZE17krqcj/2jcA5AnigPcEkw
CZXP6xs8k5oTHzLgueXefxVRxJ6Xrm1tuGKDpcol07AywpkCzAze7Tby/PdLE+GLNKRwrKdjdwcu
V0FsVFO6KnvTpP5CJl6beoUzk5e/Lt2Dme/b5fk40VMNgLTpiAqwdj7tXwN0GmHvR0oEzDQiTCzf
dXBwcgWMNlYZIncWiXerAPfwQ5Q732RAgZaRwUIlPk+r7MTv6hM9acFb/Gl8iZ5VsXXBvX5sVwJC
GsfGc6e7mN6fpa4kGwm2Tbgu3neS2si2B8WQGJFOuecXZMZeLaIHPSmeZEPGzz8qA9DYirx6LVut
dbi9E7Ta6ZWpiTIiSaXH6SuWDcs4VEApKl+LPn5PWKvpyovCjZBaiQfWEYFKmC4pFNFWaywCSgky
xPfP22gVt4KbR5DR6is/nCDLIRDlh8bDr6dufxK5C/oc+2eILeqgs9YBT34OCAmdpKCD/DpHLQrl
An/hptrY4PrqLxnFCjpPIrT4PPnM514iWg8QIfadfGwMtWMwbu1ZkMR0xuuA1e7AT26o5L2ldN8e
3eCuJBlSbTlPGZzZBBV3/Zix1pXaxM15EMKfLf/MR0GrJHX+U+NEfWnC3OL7S9tcQMdvToxTfdy0
lCM4tzWAWgYdMAoH4tSU+SQ/+/+bpxsGBFeSkOTtghk3N1GAtsnfJnfebY+nfEkeLdQFHwC7U6bH
iuUI9NFmLreZ4XRrvXT5A7nivy2slYwAk7dW6kx5HdpBRYb70VpZLrh/87ZK5V4B0P9BpjG70LJ1
OznCKMHbQAqIx9vItH3VmYi+uX+iXV/ITHTOKpEfzFPdWWKD8JJR0WyoQWPjHVJC2RZtlJ82YETr
CYpW8ZYUoiOgiXXILtpkUApFY6pxcXFv0GvZBxAJ3Ch3wcHbmIhV7w5BKPOAnU3hfpxylh1f3tx7
sgaavQPcJ7+Iyw3rxH5JBM1BlKDkte11of+cUKaehs+mZV4nXMGFZMhZdoU6+U4VUNTX5GlD7ReF
0eG7TBg1XfXXdLRzlRNCgzrEuTrX+QXekLnqM6BULAcM4jdJ1LWmY2nT9F+BOPGc6B/nBiYBqgfX
/XECTkxsCNgMlR2IMuG3VKNJVcTZjeecW2JnKpLHp8Z+H08gCJmY1b+3Ucf89+NW6jmi5YuJuQgd
T84jhaSEJdQrxgWmoBK9UgBWlF0jJckRLwdjkv0yE4EKQ5a7MHCGMuBnyd4g8UKy1+kVuCHruFZX
pkkhntD1cjwlvh/2qT9DDegqmVEtq6np1BUk5RT4T5B2kFy1v8B7nn7x9OIu/8no5SRcOTKpi9OM
2PZNmbhSts6YdOQuFKi+3/S8AxggwfHlN8kffxPZ5iZ1IfdXocmozACVamxcI3Kp5pn+KgcLjoE6
rWTLCsJVdYcxMMSVBp8rSjSXiICd5F987MkYyBq/TprjZ9cSLhfX/e2C9Ucl6n5oKN/w11Kzktgw
1Yv9Cg5k3wA5n8rgaErw8X9Q2NNi0y9fW2l9ldMTUsG+yEiQQ2yDXyQk4aDkZQRHDBtK5D+KJ7jE
M5HobVa0U/XagoUxWBgW+EdcborvZE9ZA1lfE8cYOsshv5v5WiG1U8Xu94IpBvrULYJM5zk4et1C
tl8psthOopZXd6/PdWDWFCAitbE9CHBjUQxD5azGW2zTqVAwBOvIoptVzhoDULe+oYf7o+Qj7H+g
f+r/+kkzeuXdFSjsjYBOjAE5s0SK5MznzFU7cNZeSMFbKlKPy9ErrTap6NcOCicPQXcpdcnigDXi
Um31XkDfoI3eCjyliToweAgFAmTBESvmGVbA3FdmnM2Yf0+XbbVplpampLRhpBT7e0/+b6UWtLAi
6HYjdi0WgZ4LlQPN3UjSULBC0htWn3lzLjrggn4ONXbovMxs6hTMJYKD7KagDFBs1MSbh4T0Zp+P
ucPVtmvjYKpQ++rBwR5N0ArI804MJpW3UADhCyqJ7fSopHdykIUBBtnGBzIueJUKoRfBLEZThfsl
wTTn5yy9CY3UNcqouJF8T0WFgnV+L0PpgrOZzYMf4YaNADL15JH6wocwAuPlFnyIpVNSUFAXaMyy
P6LJFauq+nU6xZau3MSg35B0mo5/39hualGDWYMq8WiVRv7GFbGKdmpg3RVxy9URjfq2Ws8ole4a
4BhTTywM7dos9CQz81/B2W/MnsJtLHChyNuFzEqeavhEBXysf+/SI0maPfGXlX+3ib19zpgvE6DR
7qjbAeKkxhKRJJ8HqQqBjz4mgxtdBbTfbQxW1nUXADHSshV2MgoHnYnMjdgZLsPhlxvGk6ks18sK
pmKnbrrQgFnpbqcicL1m7uTwXplN7VNXE1cpH1r4vBtRvEgHS7PXx9Q+wVXzOW4Z/x3RieB2ozJ9
cXtALQTVFCDaZDn+qCDzzsNZ6Jp1DXSrjmIko7+dd9EoLwTwP8euhFCNRoaxrYXTV/1Usp3TBquu
zoej3WCUA/ukYm/YyUsg/HMLJSWgV60t1br/1iqJYPLaXeRH6d7LMxrjcIEkEsfBGZDOAF4r8hXB
kvuPtENwVmamjj+C9J6ZZFzPdiQ+0OIZTKqe74Syiu3k+B16d1tGUwmItEN5GTfeRC/AyVbrLiV3
+58D95amqgUOVMN9I3YFFmYzrV1uypQUYTZkM1FbLKjmeyZrEfJG7s4Vy//NF/ZU59fk2Z+tWiVO
cPJQpNqIoxbCiPtK3GR3mg5e3wenAgS8z8jyXplBt+DAEdiwiO5bOVj7SThl1C1xbnUnHbovIUw7
EZVBnKTmkqAQDrLbcERNX094hUwB3GzeEBhw4zB7iEq4yGktlCQhZG7CpCLxLnK7SOBCqMOkly9M
jjS3Z4unvUsLz/7m/5vD7CAQt/pdjweeItb1BgUzhgOQI63NJ6MkFwZkQoVoiCQr2MpfGfAm3bL0
EEspa2v3pMeAK/mBWFmNZmpWsWGKRhhfwBNMEIVIiGgzlnNSSzNLI655QP+iihLDkr4vC92s+LJs
3ZFitK47ejKB00YeiucAunNos8oM5VXD4A7CdVSu4m3L90oMlyOJ5Ftq7YnYg++lWFpf3pNd94A/
cjE/rBfAUOGdp+oW79txbi/aliQNkzSt6zf/BeYNnMiWKibnr/TZGvzALpXiP/Ol9HF/u9cZgGpg
sfO2dNPw5htLdBHceB4UNW2otNxg6IyD9/fltbnCimrX4iFQbd8hgnU74LwUQXZ6VVaSY8D70c+v
U3tf0UewLhps+pHdLjsID+D/uJ28aF1eh8iVJXOaOM3vFj+Q3zqZolwFvFAs/nDov7T5DxJG+YES
CiMW6DzA6zAo0Xv6Exy3cPCJe4uvul6gKKve/TN7AFc/2AadvighY/VQWsdr7S1bBn5daWQCoLfj
VwoznE7mTeFAW+L2jqt42uz7tkSsDdMsKm/KVU2FDJStn5C3OTuwKj4SE8eDM2a4ZfWu4RYeecBn
OIB9GYu7WBdWqJXKclhjVkRnb2/lJHOqg4Mt1BMAsLukz9xNFnHjGQW7Nuvo286WenBYLnW2RaTo
L1u6uDaTG/5Epil7dEaLCa2xJxpIBqid0bjr+FCWubh+pofNrdWasIJNQGLduRN+02Q2fHcyY4d1
ZMyGvQQZrzQAib6apQjAY5q7xDLXb9W+MK8ospXiM8uyxd+CBCFRZneMPDPvRzCBajorAojlVX7w
iqphpAr3rcbzl8mruD30C0oanfBUO+4/+2mQpND6IZpOjNWBxAkAljFrBCUzc1zAi11aarux3Sul
tMW6eSOdDYTfkwPvpIxjNOcHh23NWiCBkmY65D6Oh26pOrPefY1F63ETh7fiNHZwLe0UZysAtp/k
2Z+uh4UR52aHp2FdShIxknBbaMNZl1cKfzZBcu6PW8jlNun1apYRA6uKS99K1vwY9DNTfoEX+jEo
U9RVurctBq7P7RldTAnWXUlz7TTFPnR+csxLnKe8aai0jNUOrre7Ca6IxpXea+lXtPl8fGNZj+69
VUIL9E/J1aqMkfTqDggYrtnelHqU9FW9unO25ZdITn76/UO/l28zUj8EjKtWOH4Edqu569mMV2wb
zkejVSPCd4cEH8+0R2dol98FlH9apH9vNiqCs5uxp0VYg5lelNnxjRKd2ZBvACkno8t+nDAq4FS7
dx06XZLuGjAbLMkIDeI4EcHxUagiAmTtpuS/chFbp4AU1oPa6/U4zDW0JNlLXb8QIyxYxFMCWUr+
s6NdPHjiS8tpRn7RFIBoxHEAqFqIGjmxcHzdHi99Pecjx0I9hqEd+XwOy+PeVXRZbq9rMm0vYoEQ
YZNcncjX1Q15BFnq0HlZj+pTgap4kaLW/6KUtLTKWDHcIvAYbjHpznjRXXlpqJFZeNwygumMeC+i
pOJhFaTlP71WMr3NuwyAu1/VQdypspbxmMe8w9Zw/ct4svCRLimgZLhqyHJYf85CDtgx1x/tdP21
prkg+t6Rom6B4qSAsR8hOdJUn7i4jAK/16pnKzYm9devgQiQnYgbEYrmkxPb1sfVv3Ct1uonFjlF
Cs723QZ0HDULsLyoOS/tokNcFnn2uXYtjeaa2Y9eWo348z7DaNFact1IuMpTqimFCl1BbH7Dm7Ub
3iJcNpUcaaJ118FtmbDNXb3UXVCFKgW+7mf69aFOfzpz3TadexsqJgx6M+RuQmd/KUSpYrvoZpcK
H9vISnXkYaNgvoh27a5j6ef6h5bl89QSZn9sKq9idZ2OYByirOdI0lYbyY9wzRt/lUzYVFUyTSbN
WeLk1Q9x+tdr2kJT0odEIBsM/zs+EvZZLEk/uj+fhfZBc0dgZ8bOYLf/Tf47+iZ67e0jBnGHlQNq
l9asPXCi+yCDukXrk1fxS8T8Scxw/FRzDq4SXjAXbCybGE5RrtlUCt3DrVIhJuOlyypb1c6ZrBJi
KVfLecg1M1B1AC92nk3Jp8r+3TzL2myPHQukSx+ZEF7XUGbMUm2Ju/1TeTpTATZMr4HQFZA5hJ2l
elHj/ACsBeufS0SO8fxwGfl4jv3AtJW+V+15cB08/VTKH6Y0NPrMUf4XL2l0YNI/rRiZIxbtkG4Z
WEYG11hPMl9HA7VeNtiANaaN3ZRME5Xj+ePvOm6u1YvbLrMCNhsK9P3bxKOgTYXVkgasv8yacKYg
nHD10jIaOoFHV2ckyTUFutTo9s6zO+/HLfHOMe2UPy0PhkHYzRC35NRR3tjMbHIZTC+hTaGrK3i9
LUEe9hM17C8itcgxvr04v23rDNgLXEAXjzC+CVcdl0qSiWmZjRxWszWt/XhFt8e1N5vuD3mtpXrk
DflmoBYJuhyE/dm+Y0NE7hf/Ysqv6Ca8dq2ZYB5fiS0jvjPW+hf8v6rszlBmJe2Vcf3IPNVpgohn
IdtV0o8HBJCnzOcOIM+EOr7u1jLwnof5t7yGqy68dwCE6AGAr5RF9+XMe3tr94p/1R34Dtr/Tphc
GmxubODTYC7PbIIPyl2XJGXjk0zNKC83PPeggQf7oF5tHbcqe8DSqO3jgOAmFregdLyU8xt6qZq7
sC7XtsPOVM8BseU4Ult5FGOYudYghSUIh7nb70AGAyiSNQZ/6tI+xKRFJXjQDnLyLDoHaD5bnFBa
UB6ZsDeXg11ynXz/JhuAI4PebknQnP+TJp/hshvojV3V2R9C9qvAyrJ3akqtNjVpTU0SzFDk6aNt
vYHtGA+/j5GB6q4YsYmJ/p/1JX3kaCNkppZiAHJnN6M48NLHB50ml5SBOPtJzoBKNGbuQNOMmcOG
dSLGhcU7ONN6YbUdoANTUVmQaAWLxPSJi864xIAz0h0msrrR/e0Xy5ppgVmgfajuALRqKGpz7CXc
LfBwhkgM/BLfad81OGedafoYnKArOWuCPUNPpF44TnCsRerD2H9zz/3h58f3LpfQ/zTVkl3hwJWJ
MNmRnCf8o5yxew4KLoQov6z6REZq4TQ8kTvGJvbWuKD5A8QnMigedD+VBG87xSFScC7cNNk9HZhj
5Pq+Bgqh3oFtO6vrYzPfGpCnazQrHDI4I9Zblk330cZRc1VIici9W2pZCNBSZduskAo9DYEqHef+
HE4tp+1vmmvi9qqHmNjsIdPbVqZGmxvR24Ppp1QYOHIBzWOntonCQXZVxqE9AuXC6tOKqcpL3Bw5
ZGGb3fRUDPaRbrqpaJircD3otdEwOR16Om3kURQc/VHaQeq1M8X/11I8UVR9C275rN49OFbKtcYx
fvwkdY8IWUzbqJ0J08t9DSodQdixSGIucefgX4ppRZ8kb5mmZURksjrVWfKmopj3/2aR0BpqVyAE
qC3EUsCPhBSSax/mFYtn1rmL3VZ2LucxL0mByJNrQlQUEx1tU2tBP/TTfOByMIq7QW102JwnLgmY
tpWyifgfNY23zGTdtSb2a60mjUvT6pvtIpCC5iungDRoKXEOpYtDoP77mgW2ykInMABEx+OiNEQ1
gsdhu558fLx4jX9Ok60hNwXQ6H2I1IPXXKyCi6847krPgUXRKDT1AcurehShBtYfkRQiz7XgQyl8
Pi3cETVB5NyMFIUe1xTNVnjm0v6oopQoQaCTadR6Kl/unRTA4AVBLAtXpT3POulHjoN2wGEiQMfG
tvCkJJnPXXgGnEkAZ8pxveJgBuSvVanBmG7OLCgC41S6LPM6iXhIJfcqH2RlnUFo72zRvHHd+uHy
oUbGsSEcpH72apqw0IVcmRQlrLTo+JXxvRkeJLBkO35KwYAssASc/WB1SmUvygBOp8AHr2a6wlv3
TRY5x8LUOB5JYw5F6wxrFe3rCnKPWVuYnv5rysD+VbxpKRdFK3xrYL2j6cug4WAam35SArB/jnL7
ztkaaEZto+V57yyKG7JOiKRto2UTHlPmvwAlvYZXWIGj0uH/biZgyxSKf/vSWW9lXjGfpj95uApI
NM/1sL8mimoZ49nzoUssAvZMxx5QqwshXwOGq7jaSgi0uKQA+89zlv1vctxFiuno6/WV9s0+X7Xw
mb/U/ekgG2kLXAp+lPMdrJnkM5FsBl97Ejv8awUpXjGV5LPCGaHcBJO5KAWz/coWS+4GWWSj3EXu
Ozb5JSUy9FcYJwCsD59P4G3W5DDZpzr3n7dSRYhTH0IZK/9gu5oowaHB5DGMbBuM2uh1CE3hQzpZ
FHKAaZm6l7GnLbwYLryyAglb0qDInfH7gHMZCei3V5LSheCSGV0qZvE+713C95eiVLq709W5mvxM
zdYu3z7XJ5XSVjr8p/DvD36WM2o+Ba3qwxcno9r5jq1QW6o7VOui11YCthYI6iSvTGgXWksUH75O
2ADlBgPUqOmYU3ha56yOKgwn9thbej5TUbVmwYnFGw3pN2iHadD2WiN8ntNdAqc+f+xEHGQnQKpq
6bwrTCfGFDa0UKmi0iSPcPcqubnHYi128zNbsfmd8dG0yNdbmWqcflCDimmFGyEgAAYZeeJsN6lM
/N6AzlLVtDDMLpUtS1HFFeT4OWGojSNaEpzGiznYvKAqkv+U+Dx01A/hesFZjuvnAvNIs0Do3v4c
3RDfa6IQqHfjAzH3r2Bjq9kXpcdMakJZuK0YZIn6fc132huklZ9YjajPg6Anny8Gdu96L8HY/cAU
BldX2Y5czrUd6LiPRxEZqMiDtXJgQ9Nf2hyLV23CdZfDb7vOe9fuAul6UJsehN6DQ2nxycsb/LiU
IWtn1q8PdpWaqBwLf4N4ViNr5KVeC4MYYhr5viNFF34U+MtU39d/NZuu5PV95UinLEDZkzTbshig
NkBNckA4MZRxtEdoH1klpLNQAaKYQfo+NRe9OTUo5rdmUeqdCS/uVzLkU8cDbbTt/t0ioWIPDtMW
JFpUIWddYJEbdhEA7n3mzDqput2Hdn+R3B8RvMiGcgmHgCqntH+xQ9cFN5IqCF2J+Cnz12pZjNYP
FifHw0vzYzGE0P1C41o37gMTJ6+LRROS5dlnTdMc+dITR/1Pj2P/8Y2pqVH8dztcWqJBCxNlvhuU
iWV1wXNaWKEVQwoIaMt5u2J/yeSa0df3KiAiNenDT7qzFNWAEk43LcuiN6LSfHtygLcDC52qYczq
Umf69adIAQ6fbB0XC9GxEdO+oxB0myeZuBYvZC0tiSu3/7BSdmYXFnFFiNDftBhcN/O51Q6G1mVU
PZbknP9XFNYldlbfhpXLogJj7ZrTfHcnf6TLqiewnfnzl6jJ82NLJ7hLSK8dz6rQG1f2b5FdAf/t
gf8Bd5Nbn9dy6L/gbS7uyFYtn55LTUoc7Qj7UiI+60a569ZApi1vl163DMYgW19qXnVAUUfPXOJo
pObadHtPHAjQKHe2q0dtCXgtzEyq2EDypYa3mUNceOwEZIALBy8oBQ3Yld2aG7WJNKpAszSEgnp7
mWq2vwCzm58TGUpb89LiXYhokVLj5OtlzxSP03vvUuohWroKNuGk/o/MiumOs3SAwVMzDRLABia8
pG7z3CL6QBv/qoda4WWIpGsYLMRUUdFci70XT7+XA0kCy6e1t/Nnx2OzzDK1SxtqxsOL/4wFepKp
wPIz79SzTBlw5FJ84pi4ycoE3jzpQRqSUojB3qzlZT8o2Cet223wQnvtVR/cFrkxNEPkmhamHE5I
Lhi9GSUPNVbhVDUWgdWDfCoSI1xRo/9iGsJwUm5/cfl78Wcf9AbO3VxoyFatlK8VBXcvgZ3r8z9N
bqFzysuTqQxf2gI/LXx9txjLkN3Vi6RKEXsjPvpHPpP6eOTCxe6oH/JvsFjmz5uew9REeqsQemRy
8rFK1tu+Y3ME4K7251i/Wcl/u+Yrg9+ueynotZ9e+EuJBPk0AUOsvo5CDXzE9GgL/BQ7kYTEmqiX
5CCrwMp9KRvj/kqUfvuJ+gshZczyLEdT+F/ec6H2HlElGpFFtLjvviUJddJpSnyNlt4p4cJ2W9ca
InxhRpEkr4rZ4C1q3gEhdxD2WzhzuVGk34tBupOMeQtXGkPJesNQkUDBFQqWakCnAIjSdvm+lo9m
pSpRyiLuSws/wQfkCkAI1A2UmM0IVKWYwsx+Uid+Yd1jZx85SJ4XhPISlkNTsr1+FML2qiBeEFAd
zczOEgKCpV1rTa5v65fJCQAT1ev235sB0o6asDwgUt1eilJrpycXJXut5eFpBspezf5nmMqUkLI3
hKHBxyMNB4OimMl3t7TLh+4SWjqGYX0MSkRl89Z1yN2MF8fLmoWJfT1XRafH+Zfs4iC+NFrzmcZ3
mg+RumbWi5UWl917CVxtWBU0DXuji8QHuKRTTeAJcnqeX/RsnxqkZmydsrj7HkilMAGCed/XjiqO
PS9FuMWEc/mkFJVBR8dRU/szFDoOX/l9CiexuOIm0xQrVxOSTB5E16/x1iiJkj4RA2qwJUq/xK+Z
2GfI8Uq+lBVyrW0jzg/OIz/LZXd2B9BjeX9gVK7SXWFUBBopKE9DyWQCrCePUMMNal8WYEVPMyg8
FFOySu4g7K+Ya0SBNwMSkU1Jemh9948PC6q97oGZS9uKj7rpMR0MKzwGudkHWl3RQxDUIP84sAw/
V/Rz8X18zG4Czfc7jZXkreEXRHdeROktDqpInzhi7n8MEIB5Pf29esLrxH6y2BN4xhVuvZN4F3py
6ux42Owi7ZsE7M0IPztzC711JnqfrEdjZFrr03IEqtI6P7HuJD09vY40WxZYY0U/YMSz0LYj7jRw
8nhVMsD5fa0tcctov+Eb9Upa7zEY3yapOa0vjJokN87OZSHMF1ijkMQzicalZ1b3UF+I4CCu6Hvf
LrGq/36vOB1LtuRZbEvAHR+LHt8QsnJN7xtXpGNP8U1EuOOLP3dDqfP3O1CWduAjPQPnRMcsP0Ak
XxF40Fqq4RJpLAbG+zxwDvZIVl5aBY8pWveBJgH92Y3uN8OsrHNUuf3jsdt8NHiisFkwLkFEUkBj
OJdYUMkQBlQ3jKvxIz6xXKrNIlJPZ0P0ATtmP+sHuXmAiA3IsJIU0z7r/FFV3Hn3/tv96TzKLoKX
7QZpAAwc6AHcWmJd7mrU8CXoiaUOl7ia9B+pKygE9we8PKkgx1VoYrfVxYmZfBQKw/xLZ79Dbk3W
slWSF+im3V37seWoqO2LPYJVZSh7DsEaumG6Ji7Z8ag9CNQgh+sqcrWgg5MeonGHGVpx/NaTJqwe
aoox5v9gtSMG+ioTafMQQmlLjUZfuaNIfKsU7SJAhyK8BUzyw5XKVXbExr8FmPkLOdBep92Hchge
LUfqMzW4GLt0XfWiso5LIKBMDMsju+/luxCOJsNY7jUzsHiM3fhfQl/PSbyZzAtOEQEuHbASwYwF
qsxr9YwRsPmkkewcVitzU64XS+V5PIpTPiYrBXU2kqu1XU7Ynx03tCfDsH+KViKrlK5R93yVFubB
z3vWOlNRuvSu6lQfRbumcTlejAcmJKyKHUCkW2bsqR+YTEaS21B0Enc+7lqL/MyOoYmwEUQ223vr
pFsPUKtAYEJcPWj6lyBkXCuHsY6oI+/Xz9GC8sfQSZtCcNbpTU3yL8PVsBduthbIdjnJAoZodisp
4YVlrMlyBVDsbLv3IURFvWrOGdhu7g4DOE3y3vpZxNv6iUeHS9vRgSsaVeTtRSE/F8miE88cSA5H
v+tE7MwhtiiYtsyK/uP3IlLxkCLyv9b09+rKb/c5XHRxwejN4OWKQC/yF/S3xCdVhdi6B+7ddqpR
+2oywUDKe+QKzXNcQavkZWT9tALe5ufF/TqzVDUDYNi83V+VSngKxP+6UnVd8mmZxMxbJPpizJQ3
0Ep1sSXLaX+FBgI8sa5weNic2vF9a+KWYdO1z85KEuEZiGCLedej08Q8GBsEzM+WOm3KNwJBED93
fhfD4FYLUVVj96V6o0vuAZ4Sr2VpucavIvyLdEShzsjIUUm5s951lzum7xShgsYVIWFScAG7O2qA
tTqzddB393KB27fSRzdF0KO2aCj7lLFtNH//uYZQGiQD3ddR4sMcfIiFRndZCp/suJYGz3EYs4yz
Q+wFIbHrkuqHQB2gsD1JI8374eDtGOg9S59ULA5ZpSsiy6+pGabEZNUf3pw64XiwEwa5nVxYRN5z
paPT28LcuNV4uzjp71T3qSy98Eiv+GhzMp1BD0pdrXIM7QMWQkoXCSxxyv5pd0ACHTok/8pexafi
XYZo0TWfUONss696wLqTi1lmsPX38RB9IE1h/a/xB067DIHvJPuhdhvRYlDfqqFpvRP/2JHmVXeC
mwn5J0JUjCMIoySeoAWIGxzFwy70ikyBMrcFAUPE89ltLhlJXMPEFIUhwIJB0caIOpRDYdXOfaxj
8YRcHEpCC36pZQ2hnSvS2hm7oE5DYTAmnl+SJhiPvxNLglQgi6AsNIvvTZ7SmxDaJHQfPtMnjZlr
AGtPiX6Tij9oCUiQGEDzLo0RXGWqGS3j/vETCrgGQyfP0vm77owdVUaYofHOBwaUdYP5VCqm0/+Q
1H6zQUiPXS4tDWTwQDx7UwzBrcDiSr8qFbzefsjVZaN4KhqvzoevzfoOMmbpkq0eDvRMAUSrm2cM
evPQX3z2OTPuW8PhIhB6RgCVcCC0vIll+KgM/lvxgztum7ImhKNtjuRyYfjr4ACFc3IZYsPCOCT1
GFjp9D26MK0Tczy925ZEn7E8iuEAmQFBWwC+t62yVV6fMlC5URiok6o7iUEpALTWKqWKmw5DI0EG
UFjOEoqdpOVLYZzeySKkIkyBI5PcypnpTXh2l2CbPOQ0SvuW1id1K5PVZoFIcsbardScPGGHqCFZ
dpGNSknhi3DaLkXCjjTmXL5CoPUWvqHS1ACYhYEPuKFnRkKQN5tRVyZPWFv/rFlR2Gu8kGGfCcYh
bxCmv1yVAczbRNEKuVDBCzCPyQfG5elbuRWOoAcJYnCm0BoNorCa0IpF5kFwQFZmKWZUmsfYXAgv
QtvOQ/Q2GmSEeZh6N1dAma3GzMHyW4GvlAfhyJgpPSTTPrgnXXy5ZFv9Lvn/2m7GuNiWN/7OObyk
NbXmX3dnd9bc8klW5Ce8BjWUWjBGF6dBefnvM5EFytOk4rlCz4l7JNNiK7ep/g05fZ4mZbN4PnRR
1F2yrjk1yrb0V1eETr8l/kRiP/UIyqmVkykQo2svWw6LXFUI7mkIwowd6Z2rlUuRkoAA1CwpV0Lm
1So5Dsp+1X2UstWKYZ2aqSe1ORZPvd53IbV4tZCDSKsbcm8c70LpHx88sFbCPxSXDmKgjth+m4KZ
JL70I+TZFQ+/nYwDO6zU2khJiAqe0IED149R0Qhix/lziD9GLQRcOaUo8FEKN5tmgzuLtFpfYXuu
xyCrfHqYTRrl5tB7+n8jn/m0THHrifBM15whmCJDIYbaU8rBY/S3FEQlTU/cZgBCNlP5a+JbYMW5
gJtOarbm3vM4vMKgpSCKW1L6PKjUsNlHldBqmf3cidyWfnA1tqStNFmKn4gjuzCKgKPDfNocSOqz
dY9XvfozBH5eByXxVixqcgwxxlXTrLTmTDHay1nZE63Eg2ARm6xgyuAYYFB7DrkT5MM/F6zDBxPU
l4xtSkE0b5hhZlkoEaG+DcSISmTEvEz9DulUZG+PttI7dZHmdEaD8pyyliBCRVTlIizezwHLODdq
AYZn1HYdTW3Z82jk1PiMkK4b+R+PdP4Z5X9Y15UGKhzxcSmpRT+TIXw1s8RQMeFnMvQX/SLgm6YB
kGSIdHpnw31LRR160CgwUXYLRaSxBQ240kCVeZpsUNQ/MeEmfZP2qCAVqHulP0TqkoKPO8dFFNPv
q7RZ95D+gK6NFfrYgzgMdE6TOdEQfcEI3CcPLdJoMbMNfDkERQObjbiQkPQk8H1usCNArmoabb/W
VsZD1T3KzAPDA1OUSiDNpshH7NU1kVi7IrAn8JFBSQNEUo5AK4FpARqQ20O1zh+c5QqPmmBXDFHu
Bab/7bbikkwo3djnj1EOXa5oZFtW3kSFB4ovE5F4afLrg5n3ksIzx0ihr17kLl3dAOxG9pbPDf7a
M4MbXLVoGil248ckwAlNTAxofNbTDqihd4Orjt5IWnrFry4nUBSE8wDvtp84YYeASbOMsl3Xjd8l
TaZw/3UVXCTQuiYHewL8ghyyW1CX+AtAvfMCegcpIahhq9by18aZ6ssN3uU1YjCZ5UB0OkM+EJMU
nSWlEgukuqn2zgINTtv0iVv4l6eMh/5E1ULCoSTbJhntYjgVQvaCByYSALX1+MdSJ93b2+mdl9FP
K/E97Js0oVtX0hgk13uW8eVT4nEOMGq6N/8u/fDu6J7RPVFCAj17Nue53Ujo59LYNW17/IZ0Lcwr
/POz61YxbYLM09VFweIvjhCXrG3bB4fHbRpRi87hpX1jhN37WPD1pV5q061NV+9ARv7m0IWmUXHZ
QTczBpLAKpzV07uPlzvyS56+Yvj8DGMAFVlbpd87iPUt51EQ0b3xSyRv3lax1ICodDxRJbilVGCJ
99r81pAA7DQ3P+An5EdACbPt+vqF2baMeNXygJORMy3acdXrL065ZNpamXSz7oiQQXKGRMhajZSM
T4I/X3yitGlDXUhlullDb54wPa2FXGH82KUVyTSTr4RMvgU4nhW2VtLdx2rnS9njuwMn+PzQoJtT
j7qBHGuDod7xUnm+LiBVefXh0CTr9hzzCfJe9Wmfmlo1fskNdEVfIF9NgYpgd+oZKrqnAu+wacvB
yNsVZyQSNxWestlKeUBJl8WEcvFuz06/v7QWnSh3VomkgX68yrDUmmPkmuZyWpQOi1HudmOeB01d
ObNQzdyoTDaZJ61xWIEOl6xfbl5G6aMvlaWGQNVlVGpGhoy/m8oGrMRPUyRbWMdbWWnqbuTWtABY
656V/n5/3ijlMg2adJr2WgiKuBbEYfBo8Bf9l8SZ4toU59EJuTPrHTRVR9qWZW2i5wtItnpRFNk7
jBuWlK/yuqQ7Kl5VaynvQ0fXKfKoVfba2DE0RLFeCZeBko0Uvv9viUTveGyHw0KYkcCoTPZyWAgL
b7RMoX47LajLwGXl1EyjbWGObWy8tI0HyHum//mk/NpOUeet8BU8WRX06nbtnzGL2pVH8eGvpZp7
RCIVGtG1ffFM0DLK2Tz/6Pnf2WOkT+wS9yz4WhCJxEYBcov5bYQPTOa5WfpdoYqUyCa4Gloi/9Pi
vNhmZy11mKFqrQKB1Ghnoxq9BLKDSK75HTPgVMQEiseVzIKaVyEFMAj34c6f4XHnpoptiAJWNOAs
KBknoOeVURV8dVeT3k311ymbjit3EX8aL4UmMwsQFwJ29aTsKiLiuzkg9xwupYvcTMbZYNbflPdI
q1ejsypkew9lieGpp3PfDTq8KzUtEDfyX/kqHq4gQ++80r7fs4rkcl1ZdW2i5kZFeOutIhcePEWO
mXV8BJ2SSiB9RisqIAoc2QxtIyHROLFtScHh+tfyYi7VZUqMp5q1bg0IFIVIOBZXSiY49QGRVJrt
VpjmCH4IgHBXnNpKdGvMYVd3BXAzLoaqdIqpjmq3rn7vyNCBz9byz1IJUnx92Z3KdMF/DHFCugPr
NiOHNuHyqagAqCQNRq9vOXs5amDPpgSb30W7I2DjXogQ+VmLkMvRbS2Mdu3BbAgPqRY/NwNJnvsn
vcvMjn8sxdM57gb0AmccfdlhuGUSjzThlZfwIO8qfSwu/Ig9Ps1ASOVdDrIE7T/WNdCQqAiL4+HE
Lmq0y9UeqyJb3jQqaMV14N3NWwowHI/ZFI1Uafr24ImtxEtGB/Q7VhUV5CGCZeHvdfeCCv/iu+32
gEmoWRJKjexi9G8eywtsa0tEkcOfGDiOnG8Qmm9wZg6UKKn/acBl5SOH5yNvcovS8Q3wxu0nzPnB
AsiFrB3YPK/QRrnpvCTducwy9WIqcca3FRdHk58YOnKUH31gr5qN4IqDh7JRbApz44K78Zi7HpiH
uTRzj7WK87OUarWTHQyj/AsA4lLVuhvg2voQk6fnnSBFgpQj5f2y+L9KuhCUCbuncTn+gYJdLjZG
fwcR/fcwyBdiVcLzWJtCgw3IWw+G8cvh6VKOTK4a74+1J68Dz5UJsMhZQdTAcVCS4NYw5G9ostb/
Tm6HBIh9q+p0sYWHnQr2r9T2oVsyBUCTXu7wKjPScvjlfqccyC0HDcBIDAfGXXw2KJcErubABdIp
OyyPzHOrh8abDxPVnAkHjmYU35r5T39MOrSJF08PPASAxbkmd9yKiK64eFp5dTfWpsOIwSar9KbJ
4DhMFt4FE+7LIEeUWWvX0XynSH7/izZ77FUaTWG+lhXKGc5aflP8ikYK7G7RXSxaH37OAu9DsLhE
0/6auNSN/IIULOnB3kpUwFKvEwaNIILn8gLslWahN1CKPLsb0yDVYsw451XiuSjzDWc1gxvoBSi7
lym5+GJreuOpB+01R2aTqZFxb/8RDTXh/71i+vA1ls2GhiU6oLnVm3iBapkaRdNK1NFHx9qk5FAx
e3Y7SqfANRwLTBJckqTAa58fqat9ty1mKsWVfAYz16zg5AFfOAX8/UMP188SOlH3qN49Fr56VKUI
La6MV45GLuCk4w5G7Ln2ziGXF6AN97tpq1eai4vPnM5ZSZJA8oWElnE+T55jiOi0H7l5XPtCmj7b
MRP+HrtC6eLEUSRxf3IYic10QqhivM27R4FTbe8ANh/q3sjG8QlRslU2wHhH9QLilUZ6IhuPLEUM
nELue3MnzXRbdt/mVIKN54OsW9NbQ2yonhD+mGGJQSdoUhmeqzEFKY+MIBMRBbfScBZx10XQBgI/
zzZivQjCZYj9YOaif2YBtsvZBuJea/BQVXkUMsJQkYMvtcEX8A41pvh6NTgyjpl8IS6sSaq4SOcp
dTw26j02812uhgSOMhxO8TOoFugPL6Zq/GXeISPc3yuqUiGgX9Meh4qX3yPqPUGJoMAsb/V0gx4P
bTxqWia3eFVqbRKH5gIQsWwsjTZiTHHjK4G3ZpLTq2DNQmUv7jPJO4reVJ3bpq5+jC81MFtPMzOs
07lrnXadxVNftRt9dwFeWx84Db5qqZ81GWlGzQFT9Dv3wcKnIrmrMgrT/T9HItTv2OSde1U0Gt2/
y8cK8pi+sGsaLLBl+g2BIJQEr06NpA1PgpYxrS3+S5Q7kfhxgXpYhsXTjvEUDEjMci16xhkINupt
TqcEaLDnPNItdGuC/nH6pXRmDZOyw2GkmrSslCmWS/4weVoCi5WIlGHxdLkJ7oqTZpW1COL+EsWh
Gnw2Iau9jYJm5N+IeSymYlMJ4zDP2vV3Rjak9D6RYsdaHcTZpAEcJMofYktLCWbZOjYTOPUXAVMW
aLTKTHPvakDjBGnVz8oLsbEDOeIkYipykwuMqHjLN5dg3cwUO/Yg7MMvotYBNHe1UqY7BBMje4Dz
/JJRmKccyIlX95FsAKKWEciZaLhxkCm0eEySdnsGoNKtt1oP8qe7lNctYCfl6NrdrdR/Z3/Yv3Lm
YGSSnoVeqqeG9Ht4yyIEGlFV0ucKFfTWIyXz9BwJj8HK2BViVcxmCmdSJh4MLOoRe75Xznd3O9wR
hr4VjAiMzYizlio9un7SWg64mSayB/oAW3IZ/kmteAHm/ijT5QLqcSQXzPFISJ3s2UvWavA+5mtM
DVRrg5z8EKADAabpEQz9lX0OTQgHNm8ZDfq+scVWgv/dMc6p81ATReveDpkKE9K97Y73hTm6sCm0
ta5876RGSwn0NTPvxerRuN8oyjVjEG50+lKxAg3NbZ56xYxi14L1UQOH59BzC6HE92RPHK9Sb2/F
93TdoSUG+uJ8R6D3pBK7DpQRW3jMZOeazUUr28WSZvJYMXfqRRescB/9NhNn5eg1vNyNF88J+dTs
r9pLwILA5ohj6YiBt89gY2fNFIxKJl4Yn2w7++2IR1H8LvpMMlWmyYjuq2N3OgmGqCZWkl5UxO6A
ICv/jcPcnndbpeXuKwImWLo5xorfQdA/ntnsiOKIP1EAV5BhUtovoK0OIAW1QmdGoHwhWx0SzlPD
zYMOfDEknAVdbI9nD0bnr349fImaVTT7SMXx4MRLGScRAb9ghPu/mIye+ESxB1qZrWd4erc6MOso
L8T2Pbs1ubP426AuN8XY/pTRnCFpjdGHOmM6bJiN14ydJxxtl0IyDp7u1y9wjjav4OzLT5OU1ulj
k97sBhfnXL1x6Kp82fFnPqHOiQ6x3nRvbBl0rctHhxSfGUMCs2DKAbDA4XKty71G6e4oiug39ZYp
9N3c+hrzt7PIu14eyBjMKMXqN5R13cbCqsEFFzDzA8fQFh2qfzzU5Mm+b9hl32f7X6Tk6sEecHKt
KDIR+0V0P9NFJKoutnqvka3FRzS40IZhfJs10Q02Kcfjsnx0xX9FImd/FH1uG3ETgTNUAvyALTs9
A2xkYZE170gGErxefg6zTGvUsQYh67oHKAscuqbIkdK7me+Xir9+8Y9/VYxFxhHHQPA7QkqcgydS
mS4dvN7tRg9DTBEv+nfo2msAklPFgjr9ZasSThsCa5Ty9Uro/aM8AITjY4ENwjNNBQZgsbuiQJ61
gN/LuoStxTJRg4w8qIfQDiFULRePrFSjIp3XyVWbxY3FRrDekejeIUgYu8H9vEQeMdo9W6a/7SYa
IweIbrNDktqiFa95+nNSQtVjQpoe+QEJdbCABEw5S6PqKWgqg+1g3DBhgnf7QjeXrgz+X6Ra07YS
e1MYFb2w3vwXl3+E2WERyePNiI5mMToVbUw2o/buZDkEVkq1fcLaacDdebTK01xO4QaYnV8omuDt
uWu5f0uZDzTaKQ95Lu4fbb8aZr77TGKPyJbrV6wDVELBQRyNZjbn567LRFFJS5IkBuCHY8m/2z2B
dhqR4R3uyXXYGEZ5+/iU3fqXC3UJbX7aXDS8EeP8cTsaxti8FJhnJJf+lrdHhHFTVzBbZnzcCqzQ
oS6zzXApYb1tuQOCiEHnrKcIRdBPiBcg61RY5h3zWeWuguNHz5K3zuqkGE+tABmIXK3/ZmiMDOEE
ppzcKjyV1b5x7BF11xGjq+aY8ycug/HW5jh8W6yODp4t7/3NDDo1sALbBKQ24pimc4+9t/0lAWr/
ezXtp8XpG1UmPt4+8cznX72zgt5z2crO7AAGg5v67Iu4PPkwlRQuIpAZ4lvz0iVb2RMpnm6cmNTI
e9v9TQ1c7n77adyOlYuGU6dgGr7asD8yf/eylFNSYQoI05pfbqwSriLwmMhoFHNxZ7M5NaKulYJF
mcojCGSI43PkyILjFtQ2+9aQupGFAy1mUeVlVUgiXaxJBVFltK+gkKBbR2bpEF6UkdV1QOHn6g+f
bv0bRpof/LpJVFQkn4bi91DxBfWmcItsCdXkI9ULA42qfu7XEMI5uIKqHCTwOu4WnYB2+WqEfxin
8CGhNWP45O7l7eK9rPTT6Lvq9s8+R6W9x4Dy5ILhjps8yveXaW7djcfPnML5/waNyaY5WnLfmV3S
BvKsLOtQezZPEoognyV76i1K4WIoaIUeRd/VnUsV7sPAb8IJk9CUqWu1nvqtOZRh8QncI3BTVm+u
q7ySQinS68K79XxbevDRHGICi8x4H7oqHIA1quPdWputapXNQabgi+3jNYF39AMEdcIOcTKnKjXc
Pgou7+WsmlEQu2wKivYdRIND3kl3QCT7Tnk3Bfbmgn3jycWMiCiL3QxvuBSQ6FihZ6uzb+RDzX6M
zCLP7gyZGTxbNAf6oO1g3gMhSS+c4GxfP6wvnmFomv4W5MP7FzdHVbbfytFi1H8m53UiYTy9eYYb
cV8gq9krR6Y/h2cXB750H4z6bSx0scrHnkKe5pHD6B82x89Mym7BEzYOVW4x2DsYvLMwD8udfn6T
85x5IaJ+LKAGw/ASpBhIAtyTIuiArhK8WmKqplI4kc3gTupNBBd/WKlV0oSr3hwFwh+63qDqFSx6
+smYXi+oCHCWmFTw9bKpYW70/2l3xgIdnXawAOs6sWCpgNCc7zkO46bHdBZhDZCFYH1OSk0ob0Ga
PR287I2xgibuNgM5j1UabONeF+qpwHZM8RgbpDJ1fTiPBaVdc0eU2C/8ihDVn+DXZ16rVdSBv8hK
VK2LBBoonHAc2/gZtv46D4G53s/HM05WQuE7tHU1Qwqbi0Lv2tlb1KFKd7ieyVzNzrww7zV/lPLq
YVRWoK2D6QAlUhBEudTxnl1LoNaBryaqgtloSkectkvmw83o8uJmJzNgAt5IXVFsCkzTSUr0rFYe
ALzn07RKJ6ic56PuOlB674BFGCNhTtg2B2h0qTgIyN/3gXcRIaD9++bhc+FnNKiT9iuAm0zY2dPq
BxQR/xf/ZDMgFuAFEGl3r4cxxRl53J0NkdV9JxP0oFGVZZbV66xcFvdT+1fMJA3GdTcPuNM50nxY
A6DKAMMPGBZlwl3dX/Ne0iRQCXGohcOFJtjBowpV2Tis5ecKUXaVE6US/xQ7amoYymSLbpwH2t+Z
kFx4MOocwrsrxm8Sflr1+2U22EStEVPH+50tUEhS5FgbkcB4mH0rX3HV5vibdknmYLiTo1a1YqHh
MZjpCQGUyiIvnxnaXYav2YNl8rnUsPQ7VQXIL2Y1/dHE59/H9kaSMoMgPaqbm29RaxGIUBYESxsI
Z76x2oU0e5zi3N04SHK891JBOM0gcZJz+9Bnus2gcEJk4sX40ctXNUwod8Kuhm6VjOoL435xZiBi
3mrIB/OWgBVwscE983jBfW1NldjZ3rxoWpw/DahlybLSasSWbXSRH7kb2TwS1pEB/Zk9E8Yc4H9b
iW8/tDo9dRfxNbfIEJNc/xWwtwwcNdn70Uj7wFldooquZmqddQqf9utHH3l4R8CNl1hizpQXFUQX
1rJwk/yeqsriwQtSG2BgWDxXGwgRVN+s7G4kFDa7r3uGuJMZaKnduPUhtSXmqCf5sZHgHRmtus4B
F44e2QAaO1pHNOVa+ncCESMrlKflIZDiPmuMy4yZDGA6n6dzwXy0zsavzNaINiGJpH8b5OOenvPS
ozX7JGUYh7rOCVmlhkCI2LlGxVFM+LkTMVyRpY2SPFWJtnReR+tEtwkZ9nWL10sQX2tjbZstOSAa
d9aoEdXgy0+3INS2pXpdY0jXhtB2gBVzozu/B3plP3bnmrjPb0t2pkJUiXHGgK3GioelSlbL3SEZ
NCU7sYJW5sNjfWLePNovTltkH9ZIR3dnvXQEYkVdGjdo2f57KgM6PkummBpzWybcfUIX5CzAX48+
Ui0kWi28aszQs0msw7hyQpm/+NaC4d4ANaeOvLMLNQPb4am8e4smHvvkwgoBP7PzMFQOHNWzkB3K
/uyarHHnYys/l+NqdZ3HSJxSW+I+86oiiWTiYXRxZ2GpC6BTxHP4sylT84SuO6eqG27RsRSs/SNH
GTYqmhyB6JZpC0u1eRdvcA0ymNVG4qaju7f86TVwwKarZZPXd6KY9RmF4KqIO6MSvWMVVu9vl9To
3P50qBI2eW+s7yuI2VnARWWSLjXRJVrwHgn7TEtHLElueWh+teNrwjFLPjdJDNMffI+eWnrfX6nR
+vEbEnAdTufpkFWQt8rUyBwc1mGmTSsUXn3stHqHvn8/ER7hXgMAO04A0BqVTa6i5a41ENbbwkzI
q5xVJfBo3mOik+IZJg77zYMfN9kDwAR4Eyl7eH+5zzFzXMo0h05RvpKX/ULq+m6YBrgjQObWt70A
CkI7q1QSRbBojZYnCk37/An/pIVaVcFzhM64z63h7HCw91S6gIiS5CdUAfcqRbVmpIlodvoeK0Qg
bsebLGBXZDFgTajgcn2LrJIQ4LXsP8oIk6vwt4L/Cph5BdSm0V1CtMB4PjI/IS3IfcHGR7Gfq9Vp
nVGulbFSajsAyXTRS7lIN1imX/atBEwmphmKlZQAl67FGd2OuYhaTurCr4TJp81Lly91kBitPLNP
QN0+wejcKUskaBM03piX5UoxHbMBiInXid7SISxSyyjPd5jQzGcx6pypV2tpezXhquLlEsjYL/FK
9DTN64syxQbhPtwYubH6W/1FNFkpKrrwXLuu5FQAVTU9hacsbNpk71VS2d6RrxB+1M7/yBwVXfnZ
BxJ2W2D7XlC2r4o9Jp575kScv2BKO3r5WmPPjrdyEoQQQpes2KrOcR5oKSfRG1QeeRCXwI3SRNS4
G5xR9XpvURfqY7aNcGiL6iNHR+OgJXiSe8jf7G0K2z5PQEKUh8dmTvuywaON2I7Fw8h9sW/3HtLa
a7D0D/XO7XwCO4h+iqY0H0aBjfe50wUper5MBpWRDUoTHlohVLhWssuEKqG2hX2uyS725Ij6IGXe
G+4W6VYe1a3DNiqTDHbLFDljXS+JlVceQtxHj6KMXL+8wQ5I4Z4WkEGEQaO8N+RKH/kYQ1EeGRdO
3jW02oOGVPNEjOAB/C59neFiYOk1oyW1bG6wvyr1tn09Cb+YEvXmgHUJsBAV9/0sU8ZbfILF7qH1
2gIpGHSWEtYfKpJRyULNVNwZDZ4rBA65tF23v1nzJiIbJnn1NYCe3u6D38ko2p/sjWg+J+vvVBLJ
Z5cMkoPv3sEz2+EXFJMZgY8IO0qdLoaY+m8bGEiiDwABQVkjKQ5730RQfZiHFAOItYKHYp4uu5Bl
72ber5Xoa+QCtXOCbQnqiIIW6jCY1S1RcM9CImJBr5JTwfhO286kmRT+Tmy6tle4wkrCHdjUyz78
FAkN/4sBfQVqOxytBmCmTA79fN3oxCQ91BYu0pYP4iRWCUH32i3OZLh8KllsdD36KPz9F6a8x0ro
1HxDTtUmRCZvCpZuGFOlauVDwSs2hqhu06kpS3GNJW8aHwhmK4pd7f+GkaLrWI4Hn0d1v8LVQQUf
CGS8esZMtNsyKeILYcFqsljcD0dlFuOzow3v1Q/8hwUX4hwkYlkSu0i3TCbl6iK0wWPdGvuJ/txF
+CtqSZEnyziGt3Iy5AJE5/HzaRNjnNzu2ke218JLSvGJhdkfrVAA8QzBAbp3Epb4pkEObiRHdrgG
uGibh+t4Tm5lapZqH4yJblS1z4U2P9ENYEN8sw3UIpsGO5GuqB3yw0Dp9U/qP63RP0oqaV44HC+R
SwB3edmSFksn4oabCKcgfFVIORAc+v5gkbeIUA4lOKaYEjsvXpQ09Ed1AKPKDyY99Z7rrcHrr8AL
hkQ6cSaCEn+iH/P/dkzxxYCIRYZnvB2iF+D3W7wsqO2gCRIPimjjgNgoBFfT6t0xPw8YGH1QNS/T
aEVhZbDXPY0Sqz1Jk0NDLoAUkTaA3HBFCKwI3hFnaHjxbAV/AMgHCKrFgSRDFezzOtAS1I4gyLP7
oPsmjMFprsthf4iM4kbv9xMOC/ML89qfFyK+21wAPqqE6sGVM1TsWPuYoBUC3RmgJ3CHQZq8XybL
KU1+i93ZVDHrJYfi3yevQ4P2uRZ03YaPoa3JGsdPSKlCHWFy8HeU6ms2fUYkPhXiVamAUs4lTM4N
UXe2wzxj7tUxZv0lGc1i+1SQCWa+eEsh97R6EgkIixRCEfwZpVvMaS93hKsImd2MW4fOtGTyTiqY
yfdjfHMdoL+BlTC800FDRTJ4mnF/tK9dCEcCGkMUZcjQv8sVcGvn+fEPv32MTn1Sp42FhNi2URPq
YThYPeqtglj0hWGWw46VgQHZ7BsuLeGgB67VIfsOJjYoKBJErjA8wGjYoy+4Q19rDXTk4nX06nJA
fUT2ZIhHUj6zLVlEI3V7X5s1IellMPvOXsJ4pH2lxfKufp7zBlPG2C2lhHqOBdWVceILxgtxXQVn
wrnQl5DiqUZHCCT51RLA5yv+zpb3Qyn8zdW3OTgiZgYZf7jpi6WZvBc4cWG7Zp14L9h7JL8MrD2y
LNtUX7DDTkKAid+ipukrRzInsifebKgtsPQJw55nXD+dce60vKbL1fTuGlbib0HhemQ2OT4rfJlS
xeIYT+umaOv6BIS7wfOJt7+yq+TAD/xrk0fN9h03YJT0XaDy2WXmOEiBv0mc/n2ZxkzjSPc5ws3a
gso7L84t1yNmtot8roIaEf+kvVcaH9U0nnsORhaiv45oDPj35CxS8Wzq167uGIUP3w2m//qT5UuP
eqBk8d28hgcemQlImgJW8gZ/QMTAKYGm9aI6cPMeNs8gQ1WZd0uUKX/V5BwxBmMr42vXsxyep600
GPjuk1XoTS7WhIkf8LTza4cjzoBTj9wlWs9kzQbdN2OgubRE3qemAaCFO2Yk8SYnF5m0Jc/9cmHi
AAqF+M1NK59vgN7xbyhnC7RpAl1T6FFh+WuREsSaf3kU9Frz0fveXy1Su8lkI226G7vvClnONOtl
xBK454qdJ0ygS33nhYFvggvCsioTdizaKVuLKEaEecKaxw8ECxkswKyllK5ltNrJeeFRHXgZODaq
rXisD0IydizPKJAHXc7mLNSjk90aPzO2Z0eMEfDhGPA3b5KKMa8ve5OyFAm9d/mZsrzdb820g/yj
q5R9WMMKcsmSoX+F+8mF0DHPHnqz/Y4/nIHd4BKAL+6lihCScZw+OiXtdRYxNIRju6Hp3iJeKYyP
wV8n2/6SD++ziBTJzaaqgoQuvJBBFiV0QcoSift0tzU5xbXZEb2eRIPogAu6+undJL0v3rr1Npvc
/5SR52DmrYInB4lrlgF+S2B/g3h2ia8GO4YJAenpa644eyQA6z0sRSPZ2PsU9CbwhEgwhmbQLut5
EcOwFli49IL5hTG95oMT2gqEFy2me2YSGUfQeDycIl8irgTn7r3WPdzBXnxlbowR7cLb1U3+I0Dz
nYsAPMuX2HCik1N8pPSRc+pn/lbfc+0VzMQxry+bXeLEHS0dZh/yhRfoyqU3HQ16RObQBb3wnGW0
L9ofKs9stAmKwh8UURJiWO2zAtIZe2YzrsWFKUDB42wp5n4V/fE5skQMLw3GO28wovp8mnyqv/TX
fbpWxdPm2c7aQXWl/2BQhWIuDf8d9N3QK4Xy97QNtwU6OXS+QQyjz0vEGEQ84camfhtSeIZ/t4tU
nSncs8ffxJPtMjIXYOWQ6kAg/tLL6d6dYJz8GcTvJciQrBGPPmujlGPeOprIqzT/7TeZs8ySBa5U
IJKRHhh5iOEjKaMAaFYdk8rZSZ8STaIQANS6IIKrWgmx9IwW++nwACf692EJb9Qwrn2UoRB++nZK
ZFljHHHHJ0sofWqX2KGESzt0SJnBF51pIGc0lsPFvmIZeKZm9c/D1oNxcEF55lfGMBO/gQl8Rlb7
lw+GN9vjkzWG43XRVKfSOI1NghBqszTfgEd3SaIjDkz9GHt2zxYiVxrfSDzxrhrpNgQgRcZcsP3q
z4jEy9/tmUjXU+VdnSJwkxaXTTaXnF8geMfjTiAS7WIwJ/p7+JEdFllfslkOXJiLzgCPfjwxU61A
7vQXu97sXbq/bytCgF/4Xjd9zvleYiMP1OkhlFcfEw1bsySNUtiG5hs3AHI9GrdHzmm+1a4BzWiu
JVj5+CPmxzE6JsRxT1KXx5ZsBA61T8FjMW2R6f4Tko+WDf6iM4jboov7OESAhYTUkdtBvfbqr9Ex
7zjKY7u1nVFiVLbyl+VOo4y+2VdWvpaGM2/3/wFDmuFMJrvcca5kRl2ZupzU/nz9BIKxSqAuyEKc
QpG0EO3nA/NQ0s5hpSCdWpSnAaHhOxcvFk8mknBnN7WsCbgRjKwkH49Gcdu12VXSuCrlQ4iwd6eL
byu3er0cQvGzH+ALMqopJgDWF0CFtmXwMBPjV9sLGFw/jgdkHKBWQPq/jIzhYmeM7UAZySftsxaC
+ysTLpIz/e5DaNBkxyT9vFBI2ZHxra+yarzUrCJyf+DYX588b5uuW3H9JUX3xmJltLFOuyYrRpN9
xWQYHy49lYIush5V6gmAg7SLKo8QPvPprPPryJkLbZVHxtVYUj8UXiQio9P4l8d5pqXba5fVP+/m
NHRp5Jjbswq5GjRF9nBurRcsruj5S1+7CtbfhxCXIIyWOTCbBOhsNQQBqcTZ80HToQPHqOlV6f0M
J1PmrxCky0VYY0058CP7icR55aFV9h5SGdAVzcukxVASCHHKUwPeKmp/iF0aS9uwi8z/Gm3vhJDl
eJaueKyc9J6KWJnkvjDPgHPUZGNBuiOvlWOMQooKeR1yfFlxJvayRVJhnxDijGe1Bt5sG28LTSiU
suj21xzjfqduCrLd+Y69PI44RA6c7gLMi7OQLOpDPruyfpaIUi065n2zE3u/d2MWRnsWgl6bap7p
MEwTZfZF6m8ln15V3H2sO+f49fjLU/sxq2CAJSAneSV3OFEnP69xBad0gH5KfdSJf5hNuKGtkr/o
K0UttFZsJskCQ4Qy9RqyMvtS/5tLyh4KjfXPSfTmdmqHJmxjN01XJ8K2GmG/NmEcy6csCKDnxM1U
SiqfJsvcregnN6619JTK3ZCMLmjDiSVqEmx/+YC6F/AfCL9YoWNub1JvE378sHDwmoEm0hNgjbay
FZ2mmL3IF7Jdr2LDbvthHHEzQkpiv98qKrf100Eft3emLgaoR7w/lCcu/Ytx7TbobiH38JKdH6Kg
zb30qg4EkywvgnuY9TjPMDUPkkdvD9aFvxAz/L0WQsafSQkUTF5iGEwzc/hKxal04yd7PTc+jyVg
P6QjvIYn/c161EIx8O8DUKO7wfXVYhA+ILvdBRGLQIfg9wxLMVksh1FYNiKwey8NmTxycwr2LtbB
7esoMxmGbNgB2N1MPgfrFJcOLe23clp2dIr+UfTqI6wX9JBRRZUqbj202DRK4lz2BuGT9lQPkh7Y
0VLQtgi26q23CZlxQRiZj88E1gXR/Tb0b+23AIK2nZJczM8lEDVXm1MaoxmBc7hYjAsdTUOt1eSG
OBrDsO5466Q+TwwwRQbtiSjiBvSbrV/U1r++mxCImnhJ7o1iPL5x9FLs4wU/yOGsGHF8akMf+VeZ
+boLfHZphQfBfkj9eCoNSP82NhwuS0DtyPr+7tYYyqfz2i/lPUgapC27UfWGnLurdc223hIyKcx/
gtah2Dz108e4VNNjb/df2oxSL0Wf9mTdq9/JCwWJk7GKWFUa5E+2eng7UVX8rRUW9wS0ADGsQslw
hkLplNGSPg4O8X/pZLbvngxpEMSKRTPEM1NLomczQkqK894d2D5D/0zQIt5W/NyZYRlmTCaMiFtJ
SIU79naNJN6xv3lZxoEjM8c9BBcD7W6Ln/cCUTeZ43ARqGDB5vG/Wq/OgY5h736LBzJBfMidy3vC
tK7mBxjBSpflKOM4byXYai16o4ZS3ysAjdwzeCC0VUlLbqjiE4cPSSB5ORBwtJkfE2uEdS7bMsAp
PgSVAgFIO/fE0oaaaeyEfg5ngqxaEwgSo81G2mb/EmfTxr16hWtzwCL0+T0v0SZUIR8gNGuahOzX
VZFxn9LsuJX8Mz7cAibwWoE5PMiGhdT70nDGS198M5xjnHUVq/GMthWyAUySED38WNu6a1OVJqUN
wQzeiL4RadMEyneQIEwwQD0fHCwxewQbmObkzP2y1R2UhqoLn8XXS0X3McRPLoFYxrBriGJLeB7a
eNXTQfjx0iiiRoTsM32iW4IR5OBbDW7RKtboev96cGNgrL5YC88i/jnZFPsRHjCyrVF/T15XAOSm
qUHw8crAAdbXNJkpLpyJuXurwCOMQGKuUV7B+aqorgOpRj5sv6lgX9i/Gv9+jJw2bNXw0ygs7DBt
AVmHehTZG7iXNVCpLtjBRRTBqyFRz427eXGdDcJvaKuDPIdxiSXibLKaqKnoM+ILNe57VLgwfK87
hpH2xE/eXbhxoyyoiIUFwVrTU2HnL5KkBF+e8zWqfUb1c1bXZ/VmfX615/QJUtO2adTo17lvpXom
/G2XzzCP1t17HMqIaigk1OYKpcf5LSfG59NCPChBFAg3GWcnX+Wvq0iiyIvomsAfN7Of1ya6wnTg
9ftKK8McAi9qKaxbBemw/mtzz36GYYah2C9bk/gKov+pzBBIJYtCGAAzi5tO/4H53q+LPU/UCG5X
iF34ZPq7/gQXm++U0fSb1/k0mhZ9aKcWlE438b9kbZK4WIY6/8f04q1lYm+2KqIxuXYK4Rl83tMq
5N5sia5YkNQXEQWWqU9QNIrNEeYiC5FnyszSzjz7W43+W8cPr0KGrfqFShIhoZwPoDNknkdDdxZn
42bHg65nVx2lpDzog/FNM2c6tUXDorLCCk+/2lAnaYEtP8cjk4IPUt2DlHJn4s1jzMB9nUvrm8+8
dqtC2yenwd1PAOKKvJf8KVYqzl4eTPAq3GwANOc5KXnS29gJxEEunUw/m4Uyqy7gQjVClP3esDPO
sPZ+Enme+RR2A8OCXVnqzseZKd51SarG87gkrhleLQHeuaTNG9e7VqyYZhicgVY+hhEzvQXy8/wI
qghMf1olw1EIR7B8SFrXTBzpdoH531/HKgfD8NTu3nCW2pg9eKHfAl/vMeN8BmowIaYv5GdebzX2
E5N70P206tKs7St94Oxm0d9QdclmVDNx84Fdva43+YjvoCl/ykLdzV3Bt863brcYZ3xdzuwRntgb
klLg5Da+NNdyTYQ0BICUxPGL7gwFsDuuiSseGtA9vdlfPQoe4kXGlxgXnMUIa0rjL7HcLs3yy4Jj
eZnOUM5iLIuUCLS0iLzoP8BNOijF8sGq6XlYoiXyz44f+/EAmNm7xZgkfFMlfMv1Jc7ihdIDulkl
+DWt6jHay8gteA9vACBbG5ZBI7CIZYLOvK/XdMa+TWFi4i9pzfQo0w4iUrqa8Ab8ORzuv1uIS/ya
bF9ssfAz4xSnjVQuxQwj4K77Ox62YeAt88MP3iMsFACHcHF4P5ufzucxh9ytux/i2HO9GKt14HL4
z9UdPKuLJr+FjIUwzMONrahm7TetHkKnEfFaUa/7l0WFb2RxkiBbRHqauBi+NerSOB0kW2CJ421X
EBuM0jgk2gNvbA2GgS6mN24oESMnx2u4N/OcWj3AGrqfyPYQCcl6jNmQ/OlnrW3KJz41EBBEi7e/
wF6IvxcsSYP0bt1AYQjbTPKKsqyVDy9x5iGKtyvz040ltXndBdlSevfe58FZn0D+vk0vqiFfSXri
gvwNpo9sZspr0Ew/bsECWnkXK9gnM+SkYvJUecezNIXujUQk4tbSLJg5hlTY+UABYFtc0XZO9aYZ
TTatUjJt9R2K7mtdGuTDICHrzwFO/9VJ58DeY+7USnfmtBlEONnM5nvJS5qVyNZbJ6DIjOBI5AK/
6VRDRyqU91NsfiA7hVrgH46vIeMdiDXc+XDgHnYNPJjGKrHVK2UsV/K9NJPQzdbqo72nyZEqFl1f
pOjX2sAa04hj9D3buv4W9Oh1XyArUQ8WMyPo/WOB3138DIDag8VRDG862T/uJCf0EiTZE0Bkm37a
uvaz23YZazVXzK1OrHJYHkE3HWVOD8Cy/hX7bkHZ3RswOu2TIJbW7iczfWOE8A5YuCBL+9SQaR4U
iV5yhEsAGkqNkLP9aAWNVIbBQYMPdXU8AqaeTbtYtZtWq+mewT8jGvYOUoNPszmAf9ixrtSOcZYe
1tPm+94bMY+udUNmMEb5FWubs8PJvCoiFfnJalbo7eTOYV+ZlJgLYEmEaeHXxYrL3O7FtgFDheCc
kyLnYEFhu0ybvlyhEo2rKWyHg+xsct3vYzjADWcqOzH18XnFq1Zf9lI8qENx2Sobhfk0w3xZZAxw
u6RLbVAzcHtOflgvGwhHkdQFFHK0vrMjo0XdMHDtDoceWgszOo7/7VOIH54Aq7qOgMuQQOMlelEW
Of1GN+vmrdlVvngRQyLMBNMQsfN3aSR3oDoTqf49w/CcshfkjgKeBkGAUAmLJmOOmkae4z977c/j
VuDJHAuIPPXr3MysEjBI6aKnL15XlflWnVJSYRz9W0ERGV6pPxVO8GeEnK5VwzMyiJvI/cWUSLq2
YonajU9910hpTmzMeIBDYbPG5QRE+Jw1JEc8n5bR/lVOEq278YE+GcUdw6zZe5qU8gdO8unM43Jz
Zs4er52/iRNkIMjfG8d3tLMBQ5MC0Y9RS9OF42FpTC6NoShSWwIhl0IvON1Q7IPHN8y+/hZQirG2
H6f7xcKXVzWqxGW7i42bZXBFxzLx+8+KNtc7ptNUC2Tq9KW8IlTRvuV18ekt6abTL7fH2/aO14bs
hRqMD1XwxFed86i1S0c4xPSQ0PdA1UkQmcFXLlAXA1ND+YvW1dYqPDolvri6FfdAke8J3pdYTOWC
awCCJeLbB2FNMwfR1oSIABCbcvqID868b7TRbxpFjO4323vdKCjApGAtdT3tzk7jD50p1qS4G4Sa
eiTX+vqLzWXgzntbYnJVfPoBrc78bnqiu6QVTUy1xqh3KN2vtxwCQmifp/nTtVt6gHse6zqVugfS
Cnmj1yZ+xU36PBW4rQ2fr3z2EnwhXeLSeSD+OzU7wQYn+uFLeyKtdDSgtUItDos6TCVP2Xawuu8c
iifKKFlCvvePEfbari1g5Izhj0YtgOYKSiFhxa8vhkiCs2O5CvU0C6Gzae9Dyx3PxFBx2BIYub4o
d2xt4VzEQQ+DnrdcMo0V+gY0nR4HpH6wqxg33dIHQsj+NrqiJgdB3euRnEO2K1LZHrqQRB3otDZ4
GcEqxzFtuN8F1eGGaj0hlJnQ1x70COyRDxVWSgJMpa57OYafoFGlKr3aeCyrCDZshXpxLFZwT3f+
LXFhfMx+37e1Dykx57JeIvlcRt7qNq+sEMICd/bp75oC5IbcVGOsJ+ypcyqTqn61aqZpUnkKlkvq
17lVwzCLVpq/dwXjhCV5cYeBIiEUt9A96bWeoKardElurgGOgpbVUE5ggFST0ouLk04uweX+mweH
DokSnp6BegCGBON6raFhBucoR/pcenLLkrZp0t9MBhum4m3ytQkB2uvTBHcS6ouU6iEfVvsAZ4px
gc/yz5rQMblOWbp5cUWcntKtG6HFfBkPHg+n3bacw4MeRr9yHNCPabiFxstuA430A6lXrI08EHxn
MRxT34IaQ8YHqQzv0iVLemBB2gKdLvOc4Aw95gLrECeCmUxnZvKx+4ISDH4xh/SwTyz7RGtYNjEQ
lMrckUPfugspIysXzi8zTYj67keHV4X4lrhBvqPPDyZehbX0V9ASPHeFPoEmJXPAr4CJtpEQEGJ3
eFPzVXNzMAED3O5o6sKnSXtcRO35ewZyZMxlpHewm86c/o3two3p+WEX4P9Lh2hvsUex6bFMHXj9
Yfj7VYAa1HBlmS1UnQkfNuWZFv8UAzinI6coMRbDjlDqZWrrCpDbdSlOKrtqFKRebcd5iAyRuMPd
WfS5fRAI4b44+OvJuyahZy6eYtDL45Tvu1aPCPrGmwIKzXQ6ElqSW0KI0NDsSBONDftVxaEqo7Hk
Q8Kibwk7T9S7Ph2YpE1J06QXFcQNG+42OUhBrvBW47HrzZv619vz6JfKHDVAWComuO9YNmHIKRgb
a5liaIkoB/ARCSB+6P5v3LH5ZYb6PRE8LbW2zXRaqycVsHaU5OfVQxoiS6W1vFTJ0ldRGJzQVxV1
2khipTkNlqcEUxGHGZ3YyEBwqs7THtpXt+JsN/xannoY54k26Ea/2CvxSTtGX2xOXYsyZ2eVrz7n
9S5AO4F0f7Z8c+m7R364DaWvvM8I1NgdvQz+OpiamcaNYYYBuCv6zFMUwjAAGSL1KJyncg7Unh0g
0VQ1e+OPDiDW7+GhD27VbYMMxyrr0Z8jNflw5GvGeQsbHptEGcyZHhKPmwXA0IGKHZ7uzJjJYYNy
Unvq4OXH11prD2Mqq0//TSrp/91dTEI6jAysOWI8NvKbwNOH0hzCneYh386VayFVHrt1ymSrWCbr
98FuhYIC1eqo8WJvKLXdSDGdJKtmem5kZclcN2Um7KZDv99xZCzrds5rs/hxuujm4Wj8eJElz83h
7c4nn6SkCQDUobR51cZdj2Nj2PZIQcXVSdazl3cB8x6CgJrMaievSo4YKg3C8ElyCpArwZ97gKvG
P5nKqNesgetUa66lK6zxTCzZ4rDXCoH7PTjzwgYhUGhlygxPe3wrtVVaxKybwpBQgWE1q66rH5H+
BUucFmPV1xC/C44xB9CLgCm8+VJ1BoJZ2rncnFeZ+FTsgbtPDSL49jTueMq1b+Nqc5XY77j6a92v
GWk6hgUgxckSo6L+q7t9tcRSyrZ8q2hIXnUkGdiuOinDWyUloJ0egAtUdt/K4HI+DdfLdPAsThG/
OSqg40beLmfOt3K5c/c9hZmxsmV3MkdEqCL8BAkPDZLtj4wfaQTRzCg935ed9EEZK8jetEeZEIF4
1UVG1QfhA09ygW9yqWaJsqMQUgB3ZOk3G1P9RiMiGSu9krHieHLJKAnRfAjSAN6iZEI8sWH35qUX
1lPi7inlNT88yIiJgpjbo6gdw4/Oaaiw6yg5RkbFL4ScY50becYyE83O83t/0TfzrDdTrZAo1RIZ
SvxHFDyfNxxnXRxIgYVaCeLn+b2wxR0cwYo+lMH8or3E2FP9vX7YkgvXCVPTmJe4NRFak4LVWBFv
swiYxnPsrgz+B/nAssX64/YikKUCArEeoRMnkvzx1kjzpTgfvmNlPuZzrW9/gto7ATdAACYGylqD
K8/SeYm78MbmWOUFXwHZXfHT++IUsx/sbu8f5B2yKf9d5mfN88KjbD8at7XgjlA3EbYSjR3kuKgV
XRUIlWFssvbwPlbex94SKRz9wOW4dCGOEdUYBc2cIfrwLWqEirqftNcKdByxG2UxbQQ5dFB8zyr0
nVFxaqjJioG4lNFIVnHGy5gTuup6wsW+mvgej1NFpkicu5Jy1q+LGfDEmeVXTg9I+zmOH87LwRYO
50IsXa6PmLbnqnlS2UQKTPu+AjIkBs4ETk2NQjW1aFYLZg8H249GJEr3GfiGKXFvebtaHOioTquX
uxg12wfPOkzIlmbb2KJ/VhORXrKhfPvKQkrdS+6utAe8815HSG9CI/B2bP8ySZrOAcN8v68SJsWS
q9OT0scVDYy2TYHyNJWemQYjduMs5dv9vPTz6Ttr8xTLnL8mR21ONcVubt7EFD8w6JjQH8oI4+fY
hnkQVw+0PWnA+qXPUSIP5vvEWswXprIGD9PjmFQ8jew0kIfJjEP9F+VcPJdxB235Wo/4iAzuwidZ
d3BFJxWkZHgF5bJIwHNwnrdxQXFwdtEymQyo+gLrk0dG0XZW0R8yI100w/AaB+5oWRbz0abOwCOK
D/k+brnSEJUNG8i3A8RPaf7oPvdzyzhnQGto+k0/Nx9uJANGA1ZEHhFb21tIFYhYpKbN7pgEYFme
JRKoIkvf6oWNFOWMacsGwTKfOjW91IpVt1Ds3Uzu0HbsNjYZD830coL6ndhBn7TeRu4QpDo4LCyv
qt+wetXJ2lQVLqez8XKPqhgG+FREqizbzwoRVJg65qbEQw9mWZs2UZPz138SUBweBvaJgbHvIgec
prtvJ36nYVijZsMQKt7ewit+XXlci5nS41/8we24xV0p5/7eZfRBzvwM3Qv7iaViOeV14AtgnZzV
XOW4zysUvl6bTi9VkSCl9LOZf1B65uIMvZcgCKI/sw4jnulG3a1/M1Vz/FryxG6XVx38QqvbnJR0
cn5011OInsAg/Tsy6mqF3fh+poNxqPbyCQ0kqCvGi3y3qfVhUnOPcbBEqJMtFgoWDiWI+vDFrH6u
WZpMDe/vi9HRINGlviWYoxib9LFVB+dRr9VR7tMZAhkxbdvAl7JSbO9pwQRTV2bPC5FY4GmJh5Qr
x6Ie49o1XdgTUgKSZJ7b33fSIRm4juXq6K1WNdHkdd7+mgKXvyvcFyAUiN2+1l5bVLMfHZePxm+U
lXmaQheUgXT6aWhaSNpUoAOmLcVFJP10KNq8zGdqAUrRpyYrjqpU51h2OWKsZxn9FJZrl+zBv97O
2wRt40br2OK5NFuM3gFrKliwb/OP8SvtVEGQW4/isQ1nhHsAbxARXtw0L1UdquMeQcGyMw3KvN5Z
9f1iXNLkGd+vBYtXHecQsvxpd7SwEehOUHFFxIjH+ggVUJUnr+Oa82YUvmdR/qwvfm94fyXtr9qS
zl7X4Xt0u0w6FBYHNzzSW/fpu3Bx6IcYfismv/2bMsJ34lMRToTKNgH77P5U9NYp9mc80f/+hE9L
TD+CgV6Rxm81ydMEQeVP8NZxPHYeab952/K2Cxb50wsdSB1NrkjPodKtXjFs4x9gC8jhnI2YJT4w
oYoSVMPBsgJyGkVO7SvLlyCLXVCSkWB9V5QEEJHylNEc4bkOgc9NhIeYGWsls3VHw+xoRODkd9Yn
HAD+h2SQGuWIjPr9nRbBe2b9tj1upmaVhXUXG21MmTXtcWxIo9Bt6dtAAgxHnGSOtxS5tyhk0yu4
LJ016B+PiuefMtrke7+PXUNGy4S2f4slEisKY3VdGJCKeoFSx7BKq4D7v9qO4Syw6naJttgv9y2J
oCLXlw5e2yWY6DStZCEzD7ARGp47Fnb9VvZtln1ymykOfS727algB2pT9ZJI+RDUJvvWr052N+gt
3c2WmOjJXwyY+ERslSlTGwEA2Nx/vNoNRc3iwGH9STv9VD1qAKsiDTjt0UGsXTkQ2a4J0USBTAji
blZyfA4TpC+LKMdGWlBk++dchAZUzM+SKyYgdho4sqVm1Yss1GAOL73oBqgGH0KE33LyX+0W8jAK
+FnuCa61weQCY0pAyFxFBvM3yGc3bwd3OIQPT/6n5R/+mAHX4svVN1UhDvYog3cUiOo76KweXkTy
FMGRjzsYFqiyOu4aRe9EdcZjU8eFe0s7TvDaMcgHVEDaX3hNI+NRxflMS3lKdfYlE8+q8dw0cdFi
ZWAe2upaoVyjs9v+qol5sliMFXaQwCNps9Gnd4LXEo0fYn17OKTqBl9ptwjaip4nqhloB3shguG1
ikSyddpWdygiVfxDPPj0kD6g0902yzy1tKhu0HdZ6/HIUhCDFG0YgcLydNbaZBbFJxEP8HugFsBK
Z2C/SDVgcjb4ShjD2FBdF2ynK1d0q6XcSFPFqZzVBsG5kNu5rN1YyOW93zlKG/es2iDB8yfm1PoN
MNTe/paKVVFDuk7BRuWbzvxCO6cVQYl+2whETL2p/A4mnQWbA9nuAmec1vfgBKm0svH6Ck6xQDxx
JxsDFk7HkoMUXemqsOvBdrYYWiUQL7KNt9XA3CcfjslpRmoyUfxgD4S/ufisy9gkAFHOSeD9lFip
BpigXzrQyD+HpqjUOYrsmWnBCbKTyEMQI/YnfwSRGRapWdbLn4OpouDmBdviNkvxprUgHrQqtikI
AF1D9yn5Ill1ej0WTAeQz17zfMztZSaaJie83Vc8b+FY+CcQ7BEaD20MbWgbmAbcR3+WAWm7CZgi
vLvRGUTSg4yDQTGyTmahAdHvttRiB3SILDoyv1sXidJ7Nijk639TYp13XE4qd0tgXONxmNL9o1vG
hplHuXdFkLVHYFY6ahlTU4VPpP9bMdtGs+kr0XNInqBJAsBAlUp2nzm4vbM4CCVVG7A++PfZI3Kw
m+ORsOtiuVNjSjgm+Sv1UYdwul7vArrodnImsGpvioOZMRZNDomD1vSKQv5B79X/xEkv5z+f3whB
dTLNQSHsOr0WhY45lA2be6rMjZXC91H65+Er2GNk50f/0HF6eaEAr8YhCWedzsrFNSfB+MLLdh8W
zEmRgUv+O+CMhBF2T8/JiJA09oN2Arbc4TWiS9ildxp+nUmOvDfMDZSQmnCpsKOcEVDwfJXmW+zM
Z+k6o9A3df5IippOVnInt1/tTb+4YPfpv2/Pwvhf4266MKao0E3vAcnzK+ZRQD+jNUA2YNhTPzwj
fHgODjA5cwwORVIQlB8OMAMfZAZsB/OQryi4AyuHgq7SqjcmFZwvKEh6wLSBL61Qa9P5Y1IaGMGN
ok6L3TnXUoXzD2tVSCuxu2nkieU2VNxyLd8k9ftzrCHHAK6qo319PNIks4I4Vto4omXoBaHagXrP
raiNwDevZxhGQYunNwpncgh36a0uWd2wnIw9Uwk03lCeiaDMRUMtCNMvSP8ToBklkvR7OzHLZ0YT
MQwQyFi5xSmSI0SsZJ8/VZ1GjrongALzSwlw4Z6E2s59UoZnqjOQNd/bjBOSpHHlXfog09x5VzKQ
j6Q9XOSMSzlpLqFHSIZ0sEpNs0q9O/qdBJYTtrcT5zIVDKz5wEVq0w/ieiEwmpYyaq+wPpaqPVvm
Y+kWEHZfZD8O5xY4WoMMoOssP8tW4Mx3PtyCaHTSYwbGL/kPCOl6lTFDdQdmmYIoCArvfoH6Xfxc
EcEDQuJzHfHF8zdGyc3pnqiRVDNFRGA2Fi9qpLiAfqhwR1fm0L16vu4isFKoR+S8U2Qd2wbCEbH9
vXlyYYHuUFpEEkJZK3W5l7Llj1CdgBbphuOVc9iFiAscspW6NQAeASMJCl3KoDCL1siOF1y4lqo9
cqDAc5QFuk+8a862X9E9qIiU7T2Z8WgyW4xhJ6SbsFcKUbV8O1yO8VgCkJ5qdbomye+Bx9esUuYN
9FEseMkR9oZ4laztMb3YSY7rlgqp5TD70vc8Oz9uZn8S/DzEmw2QgzdlXQamXgc231qbbxcrBhpC
znAat0HPKD39LVxmS6RYZgQgSsAL9QCaV+AksnOHkaDNH5ZIi6mLSu8NdSxiiJWIYv1c8CVyHulr
hQbqrOu/53MrkcBGmYjO2W7DpaEhnZjbHOy0vQR2ZJmi+YW8U7ucj/JrftvZioNL2B87INYY+PRN
KVR45kbe0VoqORJ4syKP18SO2EC/aVv/eM6whMWcyXkiUZa/EOsaYddcOSJo9TAAMvia5CkfLRvk
zyQLnIksDytooTTKMmlR+iiE3B+4w2Sf3Q1yj4LFSXCnCsp/gK8fRRV4U114H38acpY0HMPW90wI
fmUwimuyMf9xPcOb2mQrYNVOdh6twXar3kq1P9D28dD7KJ0wwOAJ7XRAlmJRTmvYQU57JNe+9z0r
Eo7F0ni5bfrFHpnV0OqHTC3PR7WUfS86aZLnyYxddLlFUiCrdBnw49vkc2YFNxiRZFiWrc4KMZdU
TUn14x+Ll/ynliaAF/FoQE4wvUPgeQXjzNC4nOZU1v7OTzfZZnCVVg7KO1xj9fsCJqkuxnOz6zcZ
jppWc2ZF3M1A837EzI7HwtPlG9az1k1RSZ2i7VK8EBD8Ty/P3+EqqR50yFROGCxi4f1k1FTwywIH
vO+3oUhUE/tcS78XZ+I4sZDH1WS4leEUMoxCyIVHTCt4RE6ctPwLmzX7A+etwXSGSOJ5OIPOS22u
QRvTsKDfEYY6I9rp0K4r+9f0gioCM4jo7rgUiNzIi/AudFXHeryaQJ9kEn9lASi6KPMeV3vsFk1Y
n+uBd7nfUb9160HJYYrjBXpQF65G6cTsvnokhS25Trjlvyp1PC9Gl7iJ2i418PlQ2B3lSLDFp9xc
Azw8IvFEYqMXIkFs5raGQ0+6XNj5kxw422yEw79k/ZOQwnkGlgW/bp2LzRu+95IAlT7Ug4ugw/V1
Bql12+mvYEQlxqVLryEEvkhwWCBbSp6YXwMgs3IAk2eoHa8vmDnrMtVdguPZ4AvTBYI+QdLBpYIU
kFBt1HVvLqeSzjEGr1ZILlsHFBonGXoRxBB0ZsWgs8M1wAH5KMzthEe0ajLxlWL6vwSY5n8y++FG
z5mJRES9LAMHQFcsgRMpGvQM7ZkZCBy7CJnK6ZhljTMwXpi5dox7QkAv1yxzdVgoGhPYZ+ns5x6s
Q1ASb305m/0EiA7vonpJM8aGLf6ADIDX0eS2eyCB6FIPUw3p4XTWjYRGT4LHTpU0XAs1IdgQyEL2
zI1sarfSHnc9F6jc3XOBR4zYLipCynITyuFkR1mX0MOVdDzonm+VIy1rnCJODryxJAgcRouxqQq8
l4/DyDU6tlbthyRxtSXJmmjZmyu5Twzq4nobU8dG5k92tZ40nAu2WIE0L/u1/mHQn4BMzvucff4Z
azR2XFELz2Cd2cQ7Sfzk8tEfui/VebV2FHM0/ewT139raihTWV1RSKcUPTaOnvHIrWlSCt2rLj2r
wvRxC6nXaQj0mfjKlZ4EMJERlI/VUKyMonaeVSs5r5UqyT+De/OcwT1a6RpIuVFZjAkNJg0fHba3
Dm1bPUBPo6CP6JA69lprwPbEXOiFtumHPwt7daBlJo1h8UJVmelyzyrXwH/FONzkT5kIyLa9FK02
NRizpdEm/bCPmPJFpQw6Yplgey8ErXcAWirSiIwmCum5tU2Vn3K+PFoh5wwJOpduNbyTaex/N2w6
APDfcf/CR8ulsQXcJl316pDHkZ+sRiGY9ld2ZwxptUissGP+tbs3xaDYRVAbsuCUDrjyPgG9iROZ
UJEbKq+47Me3MBBq4f3VtQaWnpj4xO1j26TmprFdTvGysbjqHNy/grbiv/NLqIWO7cwyz3jQMw82
hv/pfolYE0jQvryVrKXQGnLRJOhO4RBstqmzueQ1dwcAxIa4OYJUPDZxJY5hggTHjREy9yuTf9wP
tT1ExSOpcVXHRoM/daTxs60xB660gVxMDq+924mt8c5t2/06YNC3q6RggNoVBhYl1sHZAzvS2LHA
B4a9anASVGG61yEjLSclLm9wVgv3FYy2OZiA0g+VscrEJYFkgUsjEemWSHbrgKbwpylaw0m+Na5k
cEFeQqxQEf8OkxMknzM1UwAjuqX4iP3fle9uZgCxNxc8uIpqFTkzkANjUmUx3agztYFU20acJAZY
GM/8tVzmGfOkjGQ480S46vxY/gvfPUaTdooip+/VGlknjJ6tyPf6q4UedNwKz4JOiQ7Ly1jeS+jW
6yPnIOzr5YZ9pcbbdNusdFm682MVtbvqBVg6ru40xvz8WplQ7RUhLvgfDVxV2A9XQjULhajtrQCU
GfDvlm1pNzpxxnJlgXkWb1d9wvakbVX5FDsMDm1L/odJ0Jxd8xkkLzcaCWHSLWbVjcGH9/mnQ6cT
q5JKYC5UYxE3tEGyVP3y/iaD6Tx0ucBWahbhodscAmWcTywR18Nzuk3XDBKLvc8SBiOky4UjBWkf
W5b8ssSo9DkdsFM4jATqyv0i0h0+5hNsykxpnvlPSVEAL6txfQduLXbowkPbTyqsuu+2ZHoNJVjo
EyfY3xJ1jAMGMzI97jIVNlV3HzEvch+t428OC2afVHD6vCCPFVQ8hM7rwVEF8FrNdHPQG7E4L5fM
OR1YIBDqbOfRE2jVKBQ3FVjIOeGCP7owiRHGCHNyhzNuANQi5nv7eg0dafIjDxey+E9pfYnFid+K
RYAHt9NXqj5HrfsZrboempq+fy3O/CqDUJzEFKx9DwujnE5ki6xKTdAZpkUNkaQ52qxp7PiT2BQc
K7US80KWFy/wOxmtOp3lymPwGSpje5Tfke528oUNcq7LogCx1Xo+915oITjheIqvoBTFxIiTgLQi
wt72zz7r23EaJrpU0bCDf+yRVF5ZqTZSrLl+jgTyBKIsld5s3fA4wLCRtW+eEvmsIv126UEbx65u
TWXVNAcd4+Nm8wP/ySInijCLqp9SYLHwKDkegkfeRq8vzO6dc9dlLgREBiZunb31JhZkei3NmYbl
AjmWOZ95Po7OeygvxJkPX8C2KY4enF3rkr0RMSI7IAc/acMW6W8Zt5VGMH4uUksWE643VmPs2F+Z
xELUbB9zqNF/VdNta0CYKJJFE29v/Qns6Yx71iMu7siBuwFekT1d+PD87fa32xigm7g9Nd3oJPpp
SqqihyjoCewdsQPyuQVQGGqLonsBAxVWvk/1tne42eYXY5Cm9540vsJOn4LUbfLCRHfa58blbkhb
5yr96Wxoy75Z6Mgm7vw4+XLfKDPMcgh1NAcrDnU9lwRi2kkgIzh7ms3hxFxSsRNYxXi3bbBtTTKN
qEX2PquV5AbsoL15eQgcOZ/BhaZRwo/H4Iz94O2593dtTqlkDrneynbmNwUN4xgcjFvD9OAaQWA7
tmdT5IjhVeZRcWxhl9GUxuqqQxklduj7a5ipPhQMtIbNwmUqaXPSATCK4gie5IxXi9E6yJ3yshXN
sEAlieJYcLFK+T6hdLG7W09hZs9aDXkKeTkxVQtrKOtCMxnDapWDMuySI2AbFnrloyBCWpOOf4zO
GHts8IHwRf9iUivEWr9YOYoBfzbnWJVc5EfbQTsTmAzeXEOd0SWwSW49x1Bs30iYxO5UaEW9C6tk
Dchm5htQxazVeOfBA/m2RbFcN2dEENMhwKkmzEzN+qf5/UXbgVb1RgU6u45/R/oX9B5EaEGrAmJR
jLbhFgWQYn+v+O6SveANNYmuOOosEzxVYI+bdgDGX6P11XWrCRw970Ky/FTSVakbNpJA7M5FYWyu
usRDntYieNwWn9dOH2WIbla+ycouY04PKMMVYKf7Fk3tAXCfHQ+szsQmRgUhJPIcWrB1fcdw6AeT
/KdZervYSiwBeCi/+Aiy0ulMccFN62XPKOkjwi6I25HNv/+1QQRkk1BJ4XrjyUzSUIEXx/V31LI5
zkejklas/Y1w4v/Ju0NUmBgDED68xtXSKHu+3X1rzjlBGpSgW/HkkN2ksn3rOlVf5CLXlyAzj7nF
Gp96Ur3vhBjQ7H24MsiGnklG8uxocnpw5mVybqg7VfQBDWKSkL9mqEIMwiVfKoC+0bhyMlMEnNRC
TK1Euo0zb7wCydbxMeym6Jb+HSQv3vDxLFF5kl1wYruEyzaDcxZYwdSpHQTIrGbWVKSDLqB8mnC1
9i7RX6l7k5isSvHIFGEFxAGmBiKMzrOgo32wrxh8NR1PUHmyqpM3maD9roWlJbuK7+OATlWYNMCM
sMoBkiHatuOzQQC5oi8gyOXS0IVbyXwFU1kRnN1YYffUI0KUY0I+CpN+7lFSMOgKV0BdqwtI5Uxm
dsV5VUtV4dK16J8HX8LvvWMchugIX7JibCqXoK4dWSovRBXyRk+r0iukh/sJ9It9hI9WPHr5CKWL
rsxBOzir1Q/kP+9ezDD9Md5EpvpUa8Pk3Ta89A29HkS14IymOJ81m2efMfIThne7AjlSe+HWEn6T
fkcUk29QK1axqNg2MDRc7FN1ppmexiD4XGlwbUgq3SGMMPbSWYkBRwiilfUaNKcGb3iDNstLGYtL
BEW92hJRO74QPA6DVPaFeKj4xa0T69iq8vvA/yxX53KGoKDSAGM0yWEDDE7m8SZHbFqscbXCKBl/
yac0K5AOJyBqQuAWMM56EwM2syeAf+3TodIfBTqYA71R8a9cIeS68m6CBbubG7va1mTIhLT5JEbz
vJZchGXH62ACdUb+ZG9C3wr3ih0gkzt5zeVv9GX7fWULSFy69uRV7Ujz9jT1jT65wClFnPoZ0ezu
u6ana1j0lA4ec9p98UsS8/ZSEW7szUdfS3kgoVkWId+ofYsCMUx8GXY3qqfnpz4xYA1wgkGX4uPd
Jk5j+azux27h2WuVo12GbgDjNsFkHXzCI0ko9C2Gmy/h/4R1nQQoSSqBsrL57hXqtowISFCb9lH6
xPJtdi4MT1mZUJvGwq97m9O90iEpABSprHZpjHCm63Brt/3tHHnc6Fea74QgFPtbCYs0Iz0x99Pu
azMg/6CB/+By1kqsOAM0E97iz96piiGQj6R4RnZ4LIRVb9KSiHIspw2XuTmFsa/HlVQYohBw5N/X
hFSDtgIz79Cr0D4K2XfO+GE4duBzBR32hNiiCcrq0mV2fgvrVraiy60nNxmT84ncsFlIc5vk7k7A
u30H+myKn0UTLDs8sJjjdg6ltLkMCcXW+NMN3mP1tuGEGT19edx14IyLFS7wNdhi+RwTHQWbSCWV
CrFEZ/W4DE6YjsO/AdA41ub41cBb4VKCJ1ycIVhmexbKwaMLlYjzmLsfVkiTz57iaOtYuEb1v8lF
NbzJuCbzroMUf3eK1Hsn/nLLAJwCWZtJZ+qrL96+DUmaFVvREbX2c/IDp0smoQLHQ6zpmSvLg6Be
qWkQK0WxtTYyMcDUru9LGzDGlA4b9q2O7PTxzKXywW7B94KjoFc0XpjjCshViPm5fJDLppHkB/Rq
KOZI+37Nd61+gOOusCTnu9pY1yNUZovSh71i1OZiRzEZWioEdwuy/5JUS8HjSCMyYuDCO8pVL002
EhdpXCQMynitKZZytqmKszGCte579CLyoN3vkVW68w/jUnKtxluc893zHaVGuo+x0UlFXTablIDK
1kj9hvglo7XnKlF32N/0vsz6klHjQ9gsB66TQGSNPZwVz38qENAlMOHWzaFyZAEaaj2dJkO1iTFp
swj2A1hm5wqoloDlQizTMO7Tjhy8sbmySucOEMaWosDryT+kKIxSTdoaClrZWa4YhY6lix8mJhv2
BjbCwJzKuzT3HveM5YSMPZR08kLck+8eke3d0obd+XBhfOXT/7aKI82kULhhLpw6QSOvGnKsXoEh
HKQwK2Zm5vIlnFtJ6vloe8DvUTfX5/DVTCRrCC4UC2DQiLYm/39ZQ8shqU1psXceHU27zXl8acvi
liS7adU9eLKr/XhJTFaImgdE2M4+WYHg/+Vnt3b3ftnO5Pyy7WtjQHMVXM1PKyeMVtfVm9LF9HLz
90VWsjwA08RF+GBQIzS5eMiOiUgOsdubHeU9DOA3Fh1wU8YFw+T7Uh9eM2orXPQ8+mA6/VhS4i5I
P3WFoFaspgesPopSzAu7ojLQffSvWPTP/5tpMCEEvvHRy6mJgJR/Hodgda1EamhZIa8SF3ODjcJp
JUGmGdut72jRzWi3YdI1wIw96f2C+UKRd1PFlYHQzyoHLKi5VPEjbjSJlK0kusiHAKGfwYTP7v1d
8EOHjwCW68MiHTDgJVirlbkC7FJdY6Ed8LEAtqtQRMZz1+a8O3KndQZiTwL+oZBsj7HK0WlFQKR8
jcZaXjPUPazjqD5Su6tBrKTs6HiU84wMpX6wgZ3D7V0xoPjbZ9+yie2zR+RXqT1G7D7sW7WIDG8P
sUD4jA2QAEkEailc/zTej61PTY6hw2edIZYm3dCyO9Ib7eQwxIH+sXT6MUijM9DgIXwI2C6VyKXm
+CJ7bscUEiYavO8ROYtB/FxWK+keyxDlRCP7Lx8K1I9dYq88QUsGg/gNjgL+5mmCgDPoUIqipguV
S8xPiHtGXQkc7Igv5B5FYnqGQIOsp+nIOZ2/cXvpnbBH8O7OPW91Nm8rUMYNBkqRjraOY+6Bma7X
tyWC8fa4TewjgHEQzmuJ4IRiUd4tzhgSW7L+uTlD/UAMAb3yMdjTzar7S7IqZdK9/Qk38/c4ewf/
ltZhqTsjHj/QsQSIrEM55ssEpTwvg66riXJE8JNOO/YVNp2w1+bNK5KU5o41xClQdrqFgZ6moesA
Z0eK5cIj5DrDxr9lAOuBTweWN3dUHZgytCe6H6hhkfZpRFT43bN7sRpJJxNy6COSe/JHkKYxnKJr
tsF55DRgX0SFI5cg8AjYwQIewhGmbDdPDK8jovoR50XCrkS9IlP0t2JEpPLn5lhYIV/v9ZCUvBY2
erFlA08O4GD2MhrhfnlAJYamz0I83QVwwEoqjskzT5py7/rU0toAVL8FXp2WKD7tliZAF9pXJkvg
aCICsxlCRCvuo2EItGRjWH0ZwIOt9G29gGhAKH1Cz/O7yIGRSR+aVJ5jue4z2TOJtbLWcGsNUwnW
oT9c19O98ya5PBjR+mjFlgPFP/Bz1P89yyJQlyjF+Kr/4hA2idan/IdVKP5EuIZN5KZ3jMoJSX7U
ME1iWMEkVcsjDkii+yENgePUn/WUoGIX4l/9f0UBILtAYZWp4/ul6Pk3LVU1swmNwEZS3xIu/Sfn
Hajaw738Nlsyqrjh4WTLGK6iTS/6tihmzcYdXk99k8n4dQLgRWcTrknSZtpJbFaTbZqhSr2iWafE
OmCtHup0gTJsh9zVTuBw4Klmd3JJLL5tZFhwSt+x/mh/uORT84lLmeqeBjSVYrhz2xKdQzqI1agF
FUil82fCmEu0CUgrxVnnLdj99ifQoMpk5wXyx9oTYKuWO0TRKqPajFMUmVc9/aOLmAGemdsF2bB5
Bh1Uiyb9QoAL8inKJZTpMVqkRrG7u/9FQMK+85HgdxbqtMCJeXDLJudNBRNbp7cYaE9GyhOMJZgv
ASvV91ISGhZuRQ8Wd4Snxtew69m/Qxmc/fS7px9rqe0DWNFTv6qy4f3mOQNAb/tA5RfkIDc0Y92B
ylpV3U4PUgKMQ2dAbm1VGLWHEVzC/ja/8odAXsvfoMhQOXskBLdPewd9LICUx3Gw2rO+BFgTa07U
GR42G2x9BqUtYrvBW71Vlajg6x3l53mpGwYxGU3x7Y4jlGz+Gxo0/ug2KRsPoNqzhmgxApaptIcD
mzsfGW4Co3fsp26AEHqUGPZibFsy2F5C+XGGzV3H3zPqLWY3zmEFIyESYEK17mCWAQ3hmTmfE3y8
9kb4CkY+G/pDSE31XtZLEOPeQ2iFPsGwGcAlZdaS0EHyPBdGoDXFvujajFDvGArtvP1xRaPaZIzg
+v3mGNPb0pcKkZ62Z8iQBvPFXdFTCU65hYI114WCtaFlDJpZ5gjzHgoQP3UNoycYEXe92TZIm4T8
GzX+AMk+IxDhJA/KVv3S9acMv3XIRvN8NNz96xswXqUw+gw4RswaSanUfCuAVhHDNZ14xvdvcYNY
2PZJ1tRUeC8pR9HtW5VzaROV4zi1HoQj3HM1+MisjRyFrcoryNe39yIeQCsyeYW4ziYsov4x+jos
VvDSDs/UTecze85/vbG0PusAjy9alV4IBDSusVtjvPx99SJFamxhVJqeB+xGSICLldILRwfpsWfd
XRZUUXRyPx56gBdh5OW4qLqQZEh7mGHWd6LZlMiuHa+DPQGVtBux8SeEf7x5qQkxe1xc4biK37bn
5BdgMxMsEhpLhLmjW+B4nGMl96t/faSnMToni4uv8pvjPfkxv9phgZe3eTrfisG9A61GecJhsxD0
nmg57WW0UhI1cBYzFioufA90nYuWb87OkPRyqT5i9Tuxhy8yvErPOVjv7uksi325bXruXLZ5R1TT
yn1eX562fV77gGQAFNGzBsgQhBeB51ein6Dd5qCe0ARAmEXHnNM1Y6prTPKqwG8FE6mYWDba5k64
CVmoth1l+LMfWIhN25m+R9KBUal48xeYrlSHE10CqeM+FJtXYambMIAFXp5iR6n+T+3exsRMwiYR
obB1Aulcs3Jv64BQSvBh4X6FUtlF4UAt0WeqpctbQuh2ZR4r5H8K+3xs9phkh+LOEM15Rzp8sOjU
mbdaRLrH0yH/to/axS0VIN/9iXaRDoupVGGdgQkDUanRz0M5vxYdJHiNqzQp1DfZho5277/W/ynz
9/WMi/VaddVxa6KGET70XlB6eThehocYtYxl4QbhRTLzjZwjBSl92v2GMXFT7GAXYaAL9jB71Pcf
mr7pNRFyxBrxmiUFAs8mHMuTRknU+7llxcvndnxNlraDEpTdSDhx16jUGKKQIhw67YlyGFDN17cL
n8eE//gw+yJKRMQjc+psW7eLZt8tcjXwudX7zL8wfAIfrcjgSD2b8GmMxr5EG1lT0euJEhj7TFlG
/h1jNYswIHnyofLs5ngltW0UmzYN8CdF2ip6JXuuz8299lZqm/DnvLVkpVq5HMY+Eu35NHlUK1f0
/BuipMsISxF+R8m8zcvCrqGCVyK1xBjXNzcN/qr3o8v544Pjq3rjL5WFfF1Zue6k7dXmCtfsbJxl
atGnUlxIfJuD8jpg8UWS0TJGB3Z9CAyvjWRDW8h0ljQ5F7CV7jSYhWBQaV+9iHBOXhGhQo87JLAK
f8oilraG4724CI2vdlQKjnEr2XsOuf1Gi9jVpWFlpGlK3FELsiuJsi6/D8nPZZP3Rscl9coAmv64
2Pb0+C1hdHDYQF5XetrhO9VFTlLRlS4awtYP0wwFxxPXsr3UdqmT5+EJJgYc08Qxfa8NO81YmDK4
YY/r8ROKmdshOVpFv2FmJEwrtoF6SLUp0TRCSnk2cNyK9PAmeb4U2lVC07HGXeApd6pw3rtv2/RR
pyjRkt4SHqEPbBu6pOYN6FKHxU3Us3OsAcnKdvL658nAHBdWyNgvsIxfMFz9oRs8wEmF2RWIhx0h
h2+OxW9C2xKArWhZu81wF96uvlxyDDx/BSfJ3yQQkmi5jH+gzv9Ng0MU5Z3grHnM8EbWtgmWZm0z
9k13K0uE4cbgNI1Zh6tYu1M85w4cbp3OcrLkvRRFKLnHnpYylIoPOipyyxZJc1P7V/nzblBtvZij
5yorYsoylklvNMz7WUUDREDV7TYgDnZfGHWUwd+MmaCxTNv7eIJ+SeMOTjEEzi6aoFEXQCAu9elb
TuxEIOS680Pi0gNxUqLjXnhgXsDBRZkoiIIK/fd2lb8tvHqXC1WqL26tQI8plp94ul14PVSv+n7q
oQA3B5WfJgMvQL3wvebz+fe6UH3YXfQ6WIHDvyVUcDp9YLuSkORWXT3FigMxofwQOW/skyS+jY0X
yCGqC4J6j2Ljv53Av08Wr7PZzHv3ucPVzaZVbCC+VXYT2TYOOIpMd4K3B3APKDGV7b0MuAA3U7k3
BXZXGOZ7Xi4w+PQRn6P10Cgxb06jOb0KVsuusxttmXUAsezf8bcSuyXIzAidj4BkCQbfhY7xGaJO
h5XLiuO0TAQSCUFf9iD5NyUqYtIHTjt0p6oYWBixrMbQXPbB+5xHkCUCmUTRJeM18b0EBS24y0Dy
X7aP+yYrOfbVGJkn10shkjnHXKMZpM6Ss+RS+AwHjk2EBVs6VefDdKeBNfsQV4DyGM2rF6JMWEEn
uZtslX6kPFlMS6sdNpIuCKO5ASdPoAJPvdKTG0oMGrokvLp5z/T9Qyt8i/EZNb4ps4LmG1kQFUBi
BXUUcf/SkxrPRf8uVUFk5CxUkJNzeAd+/B5i2tK/SrQ1PCYMO2ol/MzOnX40d7n7Nt2WVpxqlvbu
y9nJOTj45BlmsxxLuWI16rcaV4StAjZZ82vmYnLilkJdBUQgB0mZYTinpOqAtQz6szvZC0zA9aAb
55Qr1DzTqttjcIfmp3I+jt0oRXT7T87MgIk7LmNmN2t4mmJdvXa1x0YJBZKeKuop1rBIrruPhMmN
Y/PNcTNwn2TCaKlMfrSw9FRjRlWaIMipvlxVz/KOVAkZ16gistdZHHC5PeiJMNkcZOJyJJKPhJty
aTzw/si6ydfOb+TtWPFD7yzJABH8/ZlhKxn0ZBv6kk+oww44+NxMBHuPaqPAfxVbAObGnpk9p6/N
Es2MeGC9UeTfJre9qa+cZLQdR0Gr7zCTThtWqijKVXUT3ykpOAQXvZj0yV3t0iv/O2kN9iWFUuOz
WNuUyL38WxcUaMt255NLzvzt7w3fECCNTiGXy0PJ1Pcx+VlXQ+/Xd74deN7dSpWGT3WsGpm5oWEG
BH37TrsgSetfcyPwk8/OmgnZNFfD8+v6gx24rIkgktIVTzcubGdIJ6MsFfWFWFE2ZK2EQRvvqg0M
Q64Eoo7Jh84D3ThVbgkI4laNpWrwIqjg3s+GcsiF4HZQlotvyiZt6Uwg52RhPOtQGxIB5DVdMjJH
7HBS0MhqpsAJnoLFlYRgpp8IgUBap2WIZYwlP+I6kaH6qZQYwZZvaR5NPmN8FCKO3rRR7g6PjpFk
6mARRZWKBq9H+/L/+/mOREv/V4ygzMGWlR2x9gjm+K1VDh4qdr6awuz3duO9f1TIuBFETleSexqo
ZQoUgJn4hPYxdRTNGmDUxOvfKc9eAJNsDyPI0xkP03jeCKwA0KKAVQ9iQ9eraYHdkxxfJB9gGN/2
1A+GHAZWSCqGpx/0buUkxrPdECbYwbOreOJHDgi45LQqTU6hdmLDqkPmrBx4yAB3Iap5FGUWj2Xc
/S7RgraGBSbCWW1lVXlFX+S+XKESVuWbXumia9D7elMBkMqDDtRs3ITruZr9QleSogJgrstqm5w/
gucUe8soqw0/qmUXtyoIOeex5QIUdCno8n0xB0PkRZWLs48hjCzSIDrVXUTgPwyA0l5/nbsT6Mp8
UXg1SXeMbl19LwaOPLJKMo6YANJmhIMNIbb10EI1GxFes7pg1DWVr69ieEKaimoagib5SGKBXCYJ
r5q+no4lGMV8jIuvTkGKEw+cx/k3cqcAXyfMvnlNOI55niOFCoULGKPAvyaC49qo/nn9pkLePfBy
dAYnpqt7+dExrbPPsWy/C5WBlfjria1NLVBMB+I7Rb+fcbLZfP5b4K3cx1ZLhMpQ/g8/XRGna+V/
R105c5z6EL6qC32NlC38QPYjkKbB67xs8ZxSB1OHjEQaCuvJF01dWt50XuzxpBsfLmXBGsYQiOwx
xOtJdR1YuwqwLIdge7//XWKYp0GO7jaSbjI04lHiG+GAqlIpOXUphBF3rz65oW3k1Al31awBHtm0
dveTQ+wJoI6dB22VisVykXr8tQ1XnbiaVWjvtYuU25kOlDneaVhlWSnRILWynBV5g6fU4Iji2YWG
ZcAlIRs2VwaTXHO96ePDszaRCdkE6pRIyEdVacV92mfSORNAOewo0/a0GM9PHHsqL7cM/r1RaiHB
NmZFBcKqVjVStbT7Q/M+eCiIQ92PBG8v8zgKMWIbgipGLLcsqSIwg/6mYKVAd88etplzCCZ/T02X
fxmCc6aCjHJjpXTR2jVzpUXqxCUI3nMb6oiE6EIkpBCCk6YstFCBa7jt+VgX8z3dgLWicUmgHuiP
a8q9uqIGuV4L6cTvjiVeyLSG9MGQl3DIQCy8PSg/szXM0diZ9vPY8AmUfKkqTKo+rPgapD2ej6jf
KsdCT1WhauNouwqUIjRQYCdDHp8//0S6Lsc/IW/01qRPtK2kIP0Ns0gbN9WiUIzyoB0QQhQuMlfX
/DQm5voFJeNwmCW9kJruOHveoS/X68oQOuKe9U4BbsrR6Ev2I2DL6mJ/JS2EhDLzi05mjBntaY2h
UX/6ndxrmtAWazZ8fuoaOs1gaEA0i0vJVGN28TmMPdc7s/BEy5NowNyu36jzdOySl6x8fMrhePQh
PW/bwS91bmyU2PKbBsqEXWxkfVr1DfQkXtp+zPmrNO4M62IxUTGjkQas7ZupUYxhQ+7ItuO4runo
WFWfT/JWgisdJQRNOPptR9ddQ8nWHgL6alKyYVg/WsVmditmGOJpCKBWNX30TbIJgzPF0QkQHh8S
ay9wPb4Wb5JBynKIjfn6kxHI2bBBCVOSJo+TZjJDLfF9vTOpxubJkUK1WLBD4hPYxK7hSEE7TPlE
WoLwI2jHTZ9F4HMIZh0YfLCZRr4flJzL9Z9+DX0IPG2kuYwR06ym4fyzxKTe7Yrep0ZH62KYEJvz
CcyqRaIGt01hT0Jig1kIBcuOSLduggYUu2qdQAzazoLTQ4P/OhctFWdDSfYEEGOhkPXPd9eBV6wv
4V5Idr/Y2WfFpS1G5PF5by9rJcm8WnWGzLVXnkpZ2KOx4xBe82fizD0zJU4V7zkpYlLk/hLlUMmC
YTpzp3iDs1VHSeMojj/2LfoqIHlN+w9ozDLqeJgbh0X3dfIlBhXE5OHloNXr1gwe4laGPloxXsDW
QCpkJb8JO2uCezXZvb2MQwGSV1LVWWcZ5Q3yrJo9yoaGXWoGpiDqSLZFo4bSZgitqz2CmT0acCM3
WpGyikgBklWCkQfWNb7SUfjaI0kRvaK0AxJ6NGBxumwvF0JRMXdwm5vhhKt7wHknB3jcTNRBkjgB
6KJV+0h6HUyNTX6q8jdoie7k9u0xXCz9Q5+A71yW6MFZy6ttGYTnU/Gxdef21UuCenH8suDhA96l
qPHpUX/j9+A1Z80dpttBYSIregjU04Zc332NZHBVh8lG1mktrRWAHj2EKHXxoVOmY503iOjSp/rc
PliJWndnQSEMk2U3OM0BQKp8nmQzcbJYllSbKLOuP8nS60V31k0NOOLfiUKTegB5EWbeqRXcMSU4
H6lkrFSXEL+mAze9J5EAzUEqf/xDhVmCPWlmmt4HREeRyyaZSE1RLkdaeiHRxHeOl+PdfG7JPfQl
BX4ZhmU/8AFeO/0cFOdrjlxm+Dd/eZTraC1qcCnhdD/42pAoRP/NZyekZ82Fqox6EMOYGhKSru3m
liCTm/55CO5pCP8cyBEKa/KI/blsmgA4O4albPP+xLgry9XUyTx1DUpvqhdVkiJTfzcXEGSPqs53
KYuex64ttG0GwRO3wu6teiBXMTxJUYLj0Zff4H3NhhHH6b0v+RlcKv5mUonlAbyhdpnXWqGmDTih
wD+7vrbTn41UGYmBTiHBCKDfTyHETw9jOTgb7P/qeSuwgJAWowXx+YKBrLLla8vnWbEdUdTV+y/X
SBcBr2aYMAoD/YsoiqhE31we9hnAu38f2ghd5+ktLBdL1a07/GL06K98cWPcZSJfsp+tSQgfHpo9
Sdkvy1sqhjLUWiqJCb0ZvosdDRRRGDzaOoeqhFX6R8hS2ymcN0OJw7Usx3U5Qy/MmzAGMf0zWViB
ffrcP+X+HSPx223/iW9j5enBlq+n2VphWhMypySTycifPMHUCS/qvv2eZ2HZDPPE8gSBZZURcZxq
50evzWQTlnczMmAjqIR+1f0MTdHidhBCxCSjpWY+45aTSe+rgGrQCv+Hnvm6Wer2gMj9bPy8Jegi
Vtje8wurvFZaR/g9EUp03JBv1GowyOjvSpaS3cvTTac+t9HthphCpgE0PJKm2Fvke3xhylezFW7S
Ca8C5UkELtaMp+qH6n8f8+P3hlsMczu8a7wfLrCUsIHet94MQAR86JbpA1U1kHeCttsxf8mdUi+C
kww91v4Z8BXnaAneDnpTu5H1WIVXWIpEcRtdmxnQaucNryTfdeqF5Otm6wIHIsoCjKwhxuc4dzPf
40nZ4Dbfqn5bF3qGiDuIfsW8QDMpr5k2gmmF9fDID+FwGO1KqYXmMw2yfAViCPHFZ56LBmInSaHn
H5TTvdzjPyD+/92W89+52i0txYqP3WWhGw2ZbmbpxU7ZwDMNEWq/f5fHMeoEgg10Hv7h+7goAHYj
8E0eiZ0IVw7T+lfuj5HTc2EgcWEu4x10oCKUw4f71PIpxzkB3bi9PxYwRFlKeCQm+dnA8GAhXRc+
3tJiND8YI9feszZAg7666NbTe0HLesdsUssw1BkofBOLD7VzZA0fKoU+w5h/nCmY6cElVZfPrvsF
hAnEwzdgatm7deLA2OrjqLnuCxdltonr2Eoz+CpdQ5r1kS1rZuESjRRZwlcallWdi3HB3mtdo7J+
QEJnA6lCNsklbfdlXCJxwVx349unCnZglcMBR+FbFK/j4cmksCV7Y3EF+fynMaPzsP9ECDmxdGXu
ADjeprgSkZ0KIKrsj/exmxBjUTXjc9rdtJlFS9x52IQLObKjAx9+JsajD13YuuwfxVEIwG8JakJX
3lM+aHSQ+NsgfFmhHk0V2u0FDpQ3/XP1/wY9zVE8kLUcEVL8kBxWIo6LxtnwotXDPKqzm6RUiavr
u950RxXvqNAdWl3srpOrtDi55fjqK7PcEPvk2puk9gwQOGxyDIQoshiVGCuNc07xqr6K9oe/ycbv
urcQ1BzcCuOlaa9SG9i8Xqjo7oENV3ICuU3uqbweQYQoeeqShIARux0hakGrKwEGL0eWA8+TQNA4
M0yV5oiMk2Unz9U/k6YR0QHHtOlkB9Xi7hx9zEut6Jq9z9vzoWSDeu2oKSbXX+AYSBvkATAh/gIU
19KchoJbuM0xPPdP8x813ndiS+GLjh2Rd+2YzantzyPGP3X3fiY5dnNjKWRNE/a5up65GhXccgV0
4ZN+RGqcaf29KZX4siK+UkBMCrkaAF+3Lpj38zont9MOuaJi4+Okl6z1OHtjohjX1p6j4BN/ofim
VSP+tuxTUVDCxgnun0FIDF2LHbVXGHnBimsCbidEVMIS8bD6kIwNu2NQLv9WQnQsZ9fbJOpOzFMJ
rO/LveqLjJ9Vhc4fU1U44reRHfDwmnLZVIVVMyW18IC4/6CNxuVwVQmsXwFQXTrbekbDzdywivGw
9AmwetjzCKl2z4egoNfMxIoKvWnxlP8QTLT9I1S9HIXhTjWc+3R3P03H9RiXtiyZP+IaJai0JglP
bdQhWKm04r99ue4i+C5MkjZ8pGzKip7eTGVaKQ6dyvceXhZP9Xp8w/O83zkh6c6MNLClx5e0WzbV
Stf3x14UEK5qWROekZjfAM4I4IptrJbYiO0YLbOB7mMvBCQe+qLyu8FOJAu+EpcdB+YzmG09dKNo
S5W0uFLybZewWNquIWB1gbfIH3qeHevaxwfOlJ3ja2/PRrgk+1ihB2GK353cLof0bH4TGFVrzQ99
GzpyGr5Jml4upB/IBIs9OSy5adr21uxdHJbs4YJxPIUtd8STfSZI1yepneeu1ucilxD07cVPl0xj
JqtefaWMKjAqq5oNo3mMnB6ucYfxLbF5q8NhCVNiOBldgILV+GV2PBKGHKpzSDFEky7CvmP5RWha
+S1qWm1WMqx9ZmWSYauQ8xV1kfqSpTa9vX8v/xsy7F5+jiyFY1o/mAx1py/49HasgO9TMHGkYEOz
TNc7OYI/h38UquE2UowUACHNzD+HVQvv7JCEQE9PMrcQ1VFCNKmx5s/K6qfCq3OLZVQX6svVcPx9
2G2IbNK6m204h0cJ7GFOAcce7AXD40bzTJKlEwI5i1Zz1EPHTRsP+QmBp13Y6hTUlA//Pu4fkjqQ
ej9mNGOsfp7VjZbyfSGOhPv8QRbf3qDlHo9pQIjEnyM0st9dOAOBkLR79H+DuhRgIuIz0eGlUx9Y
OMvMq6fLVCWL3NIN1Nzk+9jY0dhquEL2EYjEJKF2eYtLy4aGXFJaWEzyUUhemllWaLtk/SrzPm77
IvpIIBtzczoQOVZiMT+36/0WbOXsGDr6Rut98cSFT9YRpy9Ob9ZaNJny+jHtK933gim96yx2XzeH
W4WriMK+/57V5VYQav5qqwJmDuycQ3x3kkW9r9mR9Z4JWTJa5NFXFB6va7zC13VMaQ6MHXpJX347
c0l5YkQk2LRzjazdMGMJGyOI7M3XcB8LbSphtOdfAoTczY6Jbt4vHA+i0V7ecgamhaX/Mq93QF/R
Z+mN+3ET52uoWjoliqcevvpmeFr3cjbmp7VYc5719KNkTSh1dOSFP6P9334OSVGWq9DK1fVpJRzv
knUdNIDtFJDgiuQJUocb+Kq6SnBssY54i9bONyZ3DjtWu555MHhm+6YLq5IdiO8UB0YCsDDRpdFT
Fct6dPV5ihwATJXw08aOuX369AzJ1WEH0BdjmGNSKINfgNLRP5GyQD7dUuVzH/STe7XASoSN2Tou
ywZF8jcb+nNW+M9mu1FZkRzuCRL8XPPt/I80IDjrSFFiQYiEtgQaTWnRNmkV/EB9kxfNOx5+/f+v
qGXFozqm7RH7F1RHbhwkJ9KIrLjW091PYnCs56ihnD4cgfMTpkl8gz5fihMCNi15zmurxOktfsln
ue3kjkS2wKZQ371YddVDQ0pjFQxiiw2O19MaiP/tUCvvUfYYUB/ZDVouf6L1vvpBgZtJy6xmPFqM
y6wbnod2mn19Ty90ysfLZhto3MCjqz2nuBa96hOfRMpLD/Umf7Cw/xc12e4i0PVgiYv38Rp3muo1
JzzA22oOOWXkOApFHgasURacAx1Lg3ZEujoOy1ZJeOTN5adcgKw8zy7fdygL68Ij9V9al/uf8Vfe
glVm+DJhg4Jrs43m/o2EyHBbLXTSkleiKwpxkddfd0B0a/Mr4eYFLE+0XFdp0lAACV4CeP3/WBeK
VY9TDDOXfvq3xQ9SQDNfOKw3SydLVoTc5wpEUhhV03KkNkCGPBkDAvLpyNMyVLnr7fC8Fzfs0rEv
kIC8bVA32llwlMjENS4iHvMG8y8MtD6drIhYI3xQ/Wro64PK79z4yITj3eQRWsBYLURs3jLjYHTn
6JjlSA3SPBl1HPUI44O0E9mVRnJUSGP0TZuzjiMpKyp+jKJgNW/LKiEGBswQiI2CA5Ul8Ue3wlyf
JUlG/Mk1RkfXSJlL3F+UC0Cz707WWLPC7DAUxxjqZeEIX33NmCzg4sO/9WLuIele0NcvOJCE3s0m
JA19XCczVzjiOMtAKlx+DYcDAwda8euqsCSj9FCQNMj9Wn/lEiaeZTRvcvsSVd6QJhUNn6Q2VpSO
0zpk4ZwDjRveRfV/L2cmeaq6PwBiyYNYQ2hrRPIN4RnD/5iwIWYFvADLi+8Afhf0fPuCopeUTcJu
/6njINI6ykXIot1dNL+rgt2kEGUIl49d8DWayCW3xZ3fDCgTNQ51TMdqSNq7dNfJdoz4kDT9s4lK
BkNtylrisBYtu0JLfBYss5YCzm9ttXWOwVIQut/y3lCrpttd5ptiNsONxwIlH+/OuDc7UpBDUr8x
mbriN3u2qKIJVZSDSbucWfUpCeBfZ03vR5CeKSiCiJ4xaZJ3EYBtOWlCoutEwOoHHIxbvLiiTPVN
4xLi7Rb4o6Cfkry6uKnVrMJJJF2OLNTEofLW3elV/T/mHkETkPHuXsiOCTgnrAfLc1sJ4jtNKPQB
Hv5aYhfZFux3f37niVeUtTqM0oQGowicuzV1/4AM7QxhHF+IklMc2tmEY8eooidIt3ITloVZ9DSu
/t8DmlB1zIFhH/plQQpfQlDBC2/1l4NO2dQnLU+w1ijrMwlh4IxU7+bxhxwim4Uz2oOIdwOB1KLK
8H50hI7cy7tAq6S8KSok+TYfJVHMuuh33qrfV6fhdvLQ8pCqDpfx+SUKBS0u9CrW+b/Wc581ciWj
W6/HZKEvmZo+cavcBzkFd+0Sotq0mU9qdNcxOv01LW9qkSvr0tew3Yl96x/7ZWcyFdaWITz1zLJW
/J1K3icbjOAufkQW12fag+gfzhC83Llh2QAjA7w7oIBlqpmOBVLh3nppbFIlU1kTg8a6qv/jnqcX
NeMiYa2PcjVkTm0YPO0KtDZNTSM1J6ToVuSYAK9xBkfNzWiQx+ZTx6+3o5czz8QHbZbe2/9FkBcI
gnWWiOXcyHooEB1BsQWsNAG+f9cXZp3J1lzSKdjK1uY3N9BuqRgGqS703PgLRD94EjfjjpRSAOYs
rLBcpiOcjOAgmKyikATuNB66ubT3vNRhggNDCkysHlpT4wetmviKhFiXOjd7wPRKymlYcRAR566U
Rpf0DumlVJasl3v9YCb3lyCL90hRRiM1HdO5Rv/kZe2v6ESxXuqn/3Rod0PpnCDj3PL+p9qlB1er
A2tJAWVvs4T+kSD9Nds5auvT7tfpTQORc1r1vLyekr+kZNJ6KLRUlN9yY+Ec0uR0Bb95kOh5dkWJ
+lZFwardxU3vOaebidUbcZ4aM/jRXFYJ5U+8q9fY6zOVFGcSKsKmSM3b2kChgt4FdiB0+jHHFPMQ
WwynGocsy+bVCDXdW36PvzbLXIg3QJSUx+infkleTNsV/qAenVkiSuz1F4o1j54uDcRvxvgOjLp6
C5z3LrPTdZNg6SAYv2JAmeaCPmWOLcQdviUQ8I0Ed7pYANDdVLT7259HP/q5RVueIPt760tAdHZW
JjYvxZMGBpa7FIAMzA2pBEP0iDzslYLrD+fgXNy22WT/k5cLq12q+BTWE+iL4vTlOz8pvsBFKumL
PvU5PKVczQzwp3qYHZIrcVNw/+9GeD82T6S/4oguOJOBXNuHFU/8Kth0LWBn/9luFB8HadXSnAxs
qtba1D/OmVnQ+evBmCCF6f8P2NMSNnRW/NKIBFjMcmUOpGBa1/wNTiQiT830Z794M7/T83dUgTS2
WFCQ3v+rFewLGBLB/6qubjNZzQbVbWOjY/5HHgzt9P54/M30Aa37rKLQucNEj3rfmAS5r3A3NQXc
wZc4EHyr1JzZub3rmED2UnWWVpJhjybNW2Zc45l44DDDIHsT5khDNcvCOwLgGJpPlkb65unB3r7U
c5/bKqmtxuVRoNGdHBZSFTcNxi3ufaDdwNbZRel1DfZtSWys65d1XMog4u463306btcF4Q2glGRn
PdFX4z0bJdAdQxVdT8TzVP8Yg3OgNnKEbWftQQeC4fa6DXSEncONiKDo4NAQoR/OpWUfdW/lH9Il
EZ1opvMpJoZ2dAZ6DXd5N4j/ZtFl2tzaK9f5DPiWXwi7EDWAYmeGPApT5y+rxOzc5EFFKwm5eDsQ
5N2EIglDfnaPYSUQ18qR2Jy8tDTUHfp1stQDIjfLsRaxP1mkOsheUP4moatNBvoIaw2bUD2I/F1j
zjkAmOCToZCRzlRdi0gvkCYtYy126yaQDp1wFiv2WrV0+gXFRArSN22tpHAvaAV73gTZz6f9/L/9
N/laFCnOUdTSclXXhxQryKDJjxDUzn6z0OjSBMW5r+qi9j/39XL+ROgN0Nu4cqUdqer5YoFmoX8V
Z43v/Mlxcp6ki7ZqH0OpXf5sWincnchbfsrYEM3R2agskIy96y4i7q3OhRquEVTu8pKvPDrSsLYY
fCAUYdWC3e1AkQQ4g7J/cUB9aTM3c6IxLDrc/+0M62MwIxUOB0ZlZc4T5/uinQuP4a9QDcUeX8NL
8hh88Hwolsb+2v8NXtGCTQu7zvxxgmorLjlQY9bWIv7dLJk3HndEk0lLpZzLfbQDKzbV4WWEYzUh
1OTrV1eGM78PBdH2yZvTaaFCDLjfWkuuRsA8CJxJ4WsCopI4xMY8T2HcSEnzW+yMb06Ac9whKN3A
dRM1ubGILDIJBItfctbjEXFjhsZd0yHW+CnZZMAPuhCkswIm3rlaloR7QKBVlG0+0/kNb/H5Dlnn
OjpflGMsxkDaQf94guzwiRUjGjxlUojWHdTLtuGJ4mdhQX2FCrtEZQkwvviuq3wsDIaN08omqzC/
QDLuynvxulUnOZTTRXowEKbMR6Z+qfXE2lRhULjjNDl0mPnaYdzQjvLdsoLliT6dbzo3/i3zdbjt
WTruEre1GAOma0sUkIozrhnUUbL3VLeIBvbN6S5jJB24hwTLIPWxm0fGigUxnR6Sj3OjsTEBu4Js
j7FDSZGGULWLgtos+Dl6osLDssle7o3Rn76gOvyxp9OR4duq0p2Kbl5ZBYp0iIEM3oTyjArwCwMn
vXMgCUMI7iDEGbD0Bj2U+IyDnl226yYQuVxtj9n/aw0Xv7TRzpmk1Gi4tRWAWSs6uD+YAFOKtlJ7
pZRckhkJ6JEnL7dL/fba+BBsrVWZfz6WliTY59bLHrf6sz38osQ1TqjQHiu6/TAZRF74Ykgj9vXX
v6OtJ0ZUKrgz5KWroKjhrfiVjIqYqHzzFLOhf/ZyZcJhWRbpbbwnPAdimdgmEuwJbwpo3n+2N6Xk
Arll7HeVkQsFm5zV8PU+mrlO9+0Ebx5cpGBG68feOAckUnXnUmpBlbxXADlrRjUWZoDOXlD03pY2
pyWIM7W+MBO3ImbSG4trOdKppqjfETb8coRASoUqF/Acx8HDDs9OkoiCwhi/EaRirHbKH9ue2lU1
K7bAN09u6Gr7pQx0ZXqlhgR0jtbXF4sbOekozL2qEiY/uDMI91zzH7wonnU6qtWNNmG3MUyPhFh0
tJ3Na5lynWPRf8xpfyXKpzOMcXOls3SJzg5Ghwwr3ezc9gyLMXaPiDpAcCgz3S1zMMKp9+uGwkAH
JK7rPhKTU2mzLW9txi7EK0do1JQ/LX3cXOoyL2G5NdhPKBmSzDs7yf2UP3h+pmKYIn7oe/aORrZU
TajO/iiDKKcCwWBRHoHlnmwoj6svJlCDHFKrp5k/GGO5mEGjcjTbkdRGOh/NDn8JvVIg5KuSuFsj
km5iOqwVMs3pb1kCr8WZ/o2qxEd7kVGdMNb7FpwtcGHoCnK2J7Py+kj8jv6ShmHNLDbmaq1zfHj+
4yeUuZzFuQ8vTZnS/NPuaSf/ddG42Lr+qIpVNDVqHOK4YSrVN6getz8zR6hntdt13DqKh2s+MgLY
SLlzvq4nJcNEQTyLvqnsqohgcwN1SH2Y49vGAWuALdstoJqyCTGqVvhdV1LLJr5TIRbizvR02w/F
b0ZbF/8ME7UuyBxBWfhqboQDcCpgJ+8QkEmjQNs9CzlbgaqO9+e2o39UA0X0pMQNH3N5l+nQhxmm
yHGeCDxXQj+MQ/oOOIs/Wtj/zCcNHeRwMvFvVSjESmUBt3YfeEc1FggrgNS202IirQsgl4FTslDs
ha+vISFqFfcVDWnYTK+KSg6djZk0iHnH/23u0SeSS9IkFy4B7iJ580vwh4zMQQu1PQB5zLE3HYCp
XkzJoMuVPlbw1sIeJVdt97x1jugFdLp4aSIcJNPH+gAhd9iaPdhxjOLw1mL9POuBBUoz4HbHHXF7
qmv+WIu/RkbENaJVeNP4EL+jvvYbP6T5BnZo4RAlOMBWomoOSKpHPI1Ep9qIDf1TnyHIuMUXDN4D
EMY/V+kvAWDCnURAT5VR/i8XEScniqmtb+c5rhdmI9By/FEXUeg9kUx6LKgMQJbhIOtLZZBKGjXp
fTGCcMQLsPohOuHlXaTc7YxKoPEH8FQ5gzFDkzxgCoaHaOKl203A5dbCBnNq1+p1/oSbuXa/36FT
mDSe5CAJzp7uaLXpeK/70KKyR/yru6D9jq9oH3U6YmnTRFpURjjt9dTgAU2Zpt46kmHDU4SvVjOb
6OIScos1+DtmCiimMOj2FOoIuTUgp81mAnh/s+Omf560qUXapqOAQ1cAZExoRUOWStGlq5rfxGaN
N2RlNn1epe4JCyIeRmhhfCFd6ZHLb2JpNFRHiq9yP4nh2dBAVnrnckCNPcd1dzhyI4pC3S9K8lZS
/ch1zCD2xpv2N4i/u17mMcS3n10k0jM8c1tu2zSVMiVjOwxUVEsqZg3c5k8dlhomTPmtDy5ZL7eI
FPUeatBYWzc9KotWkNWMKbrKiUP4IaykqBCNd6Q7G8BXHoCOU2jJrzizZObxT/3x46ZQ2LS6CZgS
m6Z9mJdMjO0L4IrpNlDJEQ/r8taOBZ5myIFTAictG1eS2oKJcEduN1RAuN0YMX+11JrDfp0Fdep7
rejWBB23wU59Ri4j5o4tychJJcPwNG17MutRNTbNxD+ncIfjkzjE7iYXTz8s9fKZ44s/kIn83Ghc
NqACAugBj46ZIkTODRZnNUvyb7wJGVN35yTmAS2mQunCEDGzOKxVpBzs9WvJ6pOBk1FYkVto0Czh
2xZ+XBnl8AI6YrPCa5H54iXSVhFXXboc30setA0VOqF3lnV9AeVItx3iCUGhp7CJMHvTXtplQuWM
f3pHEaWfPJ2KcYABTBlRw6fikbvaKxJkV+Ao6TWBIjACOgjJ5gQl2xDsNINzrbeRt9ez84J6vLXe
XZiG5ha4uWyqP+dgeSp/P9MfTnDBuRhgS3KCEEmnwzU44IM8Bob5DrrASOv2GglPkDTIdjqRufUF
q8/sadFpwKUbFgfWLnBgk7IIDgwInW/37QMnfMDS3jBOTLO6GAf2wZjVjlRXd02Vb1NWx0SLgF36
Aln4xrQwc35uRo2KdJC2Wu4osM1fQOUf5/ZdUTjzIqNBM0w+AFcKJgneafaqQ4ksC8Oy8poGfWZY
KZ+bSA4QWm+pG7ieHYuTksdwO3r8u1M2S5p/A7c46Rb/VLm8267yPNfiEPodB86nict32Fpsg7dm
xZ8ItczkNna8xpj4Pmc1kPoA1nBaVHrYRefGkRmaZGtiJts0T4F/TCkaoLXH2XMUtW02UlZ++oqw
RcsWWavwe3H23CNOLKnH1eWU3+3rTrHsnFmuxJDrT8E0jgcqY1vW+GCOk2UDLN7Pw77Ij0gE6ksI
pu5yrcOnNgkfCCPaiY1b/6jxS1Ghyq9wGyjq0vw4CTBKtnMKBBD3bo036WaXLYiZURTHbc3OwJkx
jVUsJ4UwccoxFKWj/CjItZs47oY4uKDOqC7+j5U+BXeh7iNiw76dtq9fOAztyNbY3FfboAuzeChL
UrMDTRR/nZYEyPiKY6Za+GmTSR8tVyFnBo9+5x34wjeRroA6U8rIpoxk0WZsAd44gMe419Ca/A+/
i/0t7RKopAclDGjCKOmG6iUNf4Osxtx/NXdHkSPFrWdu7GyJW0IAgxG9NyCLY0TNNtv5WzPmpVFO
c6dqC+W21Mq6E6WQU63nx0/d41f9tOsqgal32GNTPeyZIDSR9dplBr+pRzBWb+Tk6BNnLRd2MIem
MPFtmkvtNR+PjganDxy1/6jGKH2h4bVLT/YqsdAW2G66HD9xda/zxbildepREPqdQMRKpvDfRnhB
h3d/u0CixGqrPHWjPLXzj/m2DW5Qyomva/Jpfj4S4rJVqRn8fN6arln/vEJKxvZSxy+qdTt54Rd6
vyRZhO/Zlp/bIIdarDeh/emP5kcbt3MuxejE4hTx32OLRAFgiyy2LuOam/cWxEhAgD2T+ENhUi+5
Rb98CAwq87A1/ulCe6pA8ZRVmsyPEGvBJ1cXYvc2OYRX+gizQ1uG5u8YZ99EGHxnwxYDWYbMsPKt
zCTxAad6CgB66l/mhBgHUGT5JKzEr5JgU4Vc0GCcMIfOHWPbLnRa9UeSpmXWsHdIlE0oNnyo2b1h
/QsnmpQGADSncYCLWHyyaLh22WdWj872XJqtGeZ9ZEVZgi6gAFdTzr0G4RUrqfTEPNtmZkGYuYuB
HhG7HYrx5+eiecffEWdjAZVEtOcDf6dWPu98DP3ceExt5JRke0k2ZDgypfNceFO6d8hhLoBuVlcq
y55hFnp4b/sBtJAH68BJGd+zg+QrgV8YZyjiVdKn+Lbvl8np/kPyBbY8d7vPNY5TqhH83rKWj7bd
B3OweRxO8mgFm/wBhHH3bflaCaFc+uYuPlJC9kZGolJppoEGI6c+TXdlyiEVOWpsZEtvmNrQBt5z
HOyIW/k4l8egvTJhu3zNDNmllGQ1W5picOVQwvMuLtLeiNAV4D6Q1sQe0d3K5FwgpVbPOyx0Lk/v
Sql10lsKrjD3EO2baKur+IzWXL5divfIga4fE2fp11rFJij72cVRF7tLLRxPzr3LeaexxqZjbIQI
T1MS0riDJiOWCHuEvb4zYxpV9CMfJ/ydL/KxjrLF/GXprrU9s+6iKQQg6IiFiHXkgbMFr9U84BdD
7yNItrTMduNe3GhFpNsFrkAU4VL/oF+7GA9eKY66HqWzwHbAn6Agt/1OS2YyfKu70eUAUYeJIIy9
NXV4cmVdQ3FdJq/HmVCF5PKcsjCrXd9X4NoSk93GX8q1WZ3BgG0fn6Q642A6koPVx6DXejeyckXQ
61jXE98XSKmI6p3Wd9Y62uX30MVzrWftSwEFZEhOgwmXOV1VfJp9EilvR+5Ck2eL1zwXhFPRRijZ
Er+kUUqhoddweXff2B7h0wRy11bdndhi+d7f+PCC24oC7S6tar+KQ+4Xx9MJ366YE/hct428VUM4
wXUSPBfgcQSqCTrdq6cgqxlIJQbTanSc3qj8JKuPnoqfbR7wWiKnjTPOlamyB7GJsKeKX9LE1J8z
y46AN2yzDSFzwiyBjT1wVogqWVdCVXzUOmDVOumouJw3XKAWx7/u0BxAijvGpzROYaJQ1RrDURwd
zxzgvQSG5zpRxuZqrfe9rey4MeQsQnkvDwale2/Iwiss9KzS4bOH3S7sBbD9h+vBiFYmvIk32m4Y
L55y3cO9li3eTjvZR3ztnsCuGC/ih4ZmH0elCYOgILwXNMYK6Eiuc0LTy6VJF4iyeeeya57COIB+
wcWP4cythQQhfXJVgml9ZlgGt4kxUfeZCOKVQ46HjOqTi0Tfly15aGb+JhopL+ebh1bj6RDEylt5
/Zz7Ug2iYZ7dVaFnjhsoTWvsuGR52TlRsn7TiNDB1fWKy1I9ab7OFYlutaaI1b2zzQP8OpgQrE9o
+8fiVeiTZzckbYQDgG8Hd5/X1QxkcxkYyv4wdrDG7VJakl25MPx4PHqdugzyvxozZB+Jlcx1pk7P
UgvNHRE2QQG+ik2MGYBaWoI3wP5GLTWyc/PQ4ntK77ChelfaszZYEyX2QTJI8kpXo1HSeRn/lVYe
xEfAImWWL0RyB10hq46P6TJiMh4r03oz8Qdl0HCrgspAPqqEt6U4hMN/kfCKcnI/j2IQ4qE7+gRg
Fsvoh0Y7w4vg2rEweulqLlpGdv3m4FdB+GJEWJ8DxqzU11YofHnkT2VLfIfZgtt2bGi5MV3eLH9d
caqG/LLA3CYXjHZyUoqUt45fRvxeTX1Ah+ZL62ZmL5M8k9/dQQAnISilO+FjQaGfz023ct+nWe3m
3e3IKjGCuh3wHflVIIe+NI8MmX1PQ1nEbLDGrcuaQ/0wzKp19meITfVT4wtU0e+1JcpKViaHnW9J
l2uE5YnsAaKyaeGtEvu0mWW8R1OsLKmoO97Rk8a9bK+zNd+fcjFpZbYt8fnOiW2JeD7WjRgZsizG
08adM4dm+KAokkHWAEOA1c3GGOIfEMCJtkef7fFaIPkIxUC6kYlq3ThVXoUfI5u3BjdlSjo4QW6C
xHs333gWBAtdrxAwkW04+sEwEPCmAmvqreCj6ZxKMLT9F8m47B8C9erlir5yHxYxFMjG9ZbFpOPp
oM2aR1h+7q3rJ6sapY+FaEH04a+rpN75ukt7qmzf0u7QDblA+hns7lheLyw+mi3Lzkx+hECIy/35
z9pwh32nd1Gp1r1DSgSwTSIhy4KKAlu0LOGVgrgzo78UOITY8M3rsQaLsis28Y9+KSbNHtTVnnQo
WtAU9eus7R4hkZ3r9ao1WencJ59+fF9dWG0Kz80VVYaEuiy74+xy6V/CtLfd7hEYyxSjsT3BVwKz
LaQHT7EpynvqrOp9/GjQaZdj9woFf0OQc2D+EeYZ+96PqsNLSc9XDmDwSHayGb9xXRDTt9vCyswV
xGwfqxVBAA0fnRA7kdoHAbX46MRUvFNP+RJ7WVfevTCxA/FjHVzGd3NyG75zMQb/U1XbkFjzfT8p
exoRaQDEx/h4zsMo1dRFnZjoXLAlZY9fg0ODVBrTSv+UL3hrcama3t9nm2413neSgKGTzY+gDk3V
fCzlQssYNglRigMIOL594Zf+gvR6N0jqJK90up1w1Wwk4HcHS3STDsss4U8KR/5dS7Eajo+5+NB3
3IqOXAYMrNXV6J7onKtCZWVyN+3vKotgw648htulSBg0QtJDfyeoJPqXbD7YU5DZQ5Nt9vDnfXsq
yz44ArzrqAhrYwRP7auRXQAaiLkeh8PuHEQutaNhd7eXAVz5YO+POqJzUS1as1knKCX6XHdp2aS+
slp1VsylbWG9F+7QsofyqaOUZJvlISY9O17G7PjnhAiLPQAd7XuZN+j3GX4kn6jOBGPD7jkbgGuK
Qb7TsG1ejQ+UahAGVL7wugeToYB/3ov1S8EK+Ho6/Bkz57gPj77yscSpA9fEgrqYnuiEKDmX3jDn
2AdMwRSWLZeyo9/OCYQPm7iWMv/IhE+qXMVCR/JOtUJfZQNmouuKchssnaKLVjV0JG1B6t81Kr0t
yz/Py1w8V1Sz/Tjz9pNc/4S1CVkdjfFmLUz3RGheoUlCbRnjbSW79PAhQcbbyEAWHoAnGQ0Opqyu
qzt0UJWpIn8LwWQhSorH4L19XLEKRB/4I2H++hbBF6hN17aKDzpsVWA6V58lbXr75vpBHypwRErs
SHrAj6kNCKaS8C5PQQbRMPuN2prYXSm4D6C7kgvJdkyqsE+moDeL8jFq4JguxwRhimjcftX/eLOJ
O+hHwC2J/fJT0RvctkMUXJjAKurGnhQ3s7tbM71nxRpjARvuhN8G6MUqb3Tv6NTPCnAaFIcnzTQG
KJx9aoqz93Vn9aH97ipKS1r6981+3oJGI9BfTTNFC1os7BhAGAzxPiuUkL86O1I1moV00gc1YfIm
Qaf/PdmdMwhZ06xVCIleDfYIUjIiP/rYdw7z3cw+f+4o4XCwrsAe5A5MaMPuU7zEr6t8VQyZzMOb
L54X92qGR2NQouRl8m5adqw8JflG0WpAjfRbIxAGZSmiHaOhOTvv3Py5d1dxjSaE+4XdamKxFIOM
e4gTtz00uStNry+Q1/VVHoS6nTurPsu3194RaRvVkdYUyE6HpfjSGEM4O4Nx0jq8JT6+eBSaKhYX
3sAdDiwEJaJx2i3mPbkJ1No2cp3tiiiSwbxrchbvP5j6QIeUlIN/IZB6+Ge/9Nr6bYH4bZ0iAszf
ssF2mTtgLH4re9Posi/XoU+453ecMzr3CdOlCwluhVDUTO03JHvh3ZXF3KNcE9RflgPUrU3aRKt3
iJ7h56Ll9zEtYyy4CjFdots2ykFFwBbC18FZVEYMXTDBd4fp9nkGb4/i2lxujvPOmrrsERYTdq3A
u5Hnh4mdkJxEu6JcGu6mk4gtyAh/QUkncB2jTjMgnaNQGOsqiP2bEqDsb9+kzv+kckXY5NPDwD85
4mHnVWwwnWdS7D3LtaG1gotXeCbSHkGMhAAkR/edWLWpunkKOrncZoOGykQiFaZkkdB78jC/I/Rr
1lpKUe7Ii2ZOyP5LfJeoJhsMrWYdBtmNvSG1sjHKBZzmHIfsRrRmzQgyat/WzQdEzn0CKHlc5yQa
gSe2xSbwE9G1Ok5R+F3MNdvdQ7MNZ/ZnFrZrO5VXhvX+PgM7VCBkbnHgLNmNq5fqTqTN+lHnaKF4
FpoYrOxTdnpXHpAXCxbfLBBA+a1ikoMmm3TVAN3/gh4dkzereamvbSLOmPSVkZFnDv5+hOMv7iFM
zMcJaMQHUBfSjE3FqB2XKIcwK424iP6KOdnGTgHTlvXHgZEW8fg4DiQ7nT8/uw9G2GbjfcEmfN/A
0TOM4Vml61OGY1Ns3QkUaa5vBJREn//w+tVuz+SZ+XsHOMAycOikZ5A12km3cWkWXL4RW6R8GryW
2EmDosZN3ebGDoK6nSstabf41a2s7bA+KMSHbwzVRHomW2uRCUW2Hfruf+mSDHeYVbAAmmPD/rnj
0Rf5U/CGMinB99vAIESkQvMHHzJoK0p8KEwNU5V6Tls2Fh/7xZyuzIEqHTAQW/Gfml7hOnBE9kL2
ku8q6JT2/XJR0c16Ikla6lQVm5FYWeYr2ZTuvwznAL/hKbJ4lDYz70Yshy+SAgyYAwIn3T1E4j12
8RJ5ZsWf4i1qxFamkfUIMBBwKgi8c/TpliqvnDGNQyUEa3vToBs0fE8LsgKzIwoouuG8k2rtKDQN
KgGQUvGndZp3BcBwpAsXZ0Nxz+pr/+sKdttMDTaYdDbDbE/LgjGOScZOnVugevezJJJU3GidoqNC
AG2T2SFiYyWIB6GaSpPAZt21YbySf41A9VEc2LFw7h9VMGkizvgbkUKTrDuguhOuYamIK4WYyec3
03AovwKYlWbceQOG/sC3Aq6/608mfDoz3R5AgwUR9F8FXSYU3qFEJu//JFzWFIh8g4BfPcZf8sGf
g4BuczxEMqZ9bAb+0r4mVcw6CH9oLp0/PA2y+BgjaSf1xLaEwco4sxWFJjplI9Zmx5gXnZg+hi85
l7ERFC8Q0y0Z0Ba3E8tpUqKk1tzfn6lKR2Mz+Ha6u404QJyCwVYimxHwTD7rmRph2ldwyjGzX0kh
zhtg+Py6iTaWlp/Ir25pzDnEqnMiuOgukCRsoI68wp6GAqyk6DGbkvwC96Xazqlxmqvit6zfLQg1
0ZQNLJR8wHrlSrWAUroQzx2OZ6zH9X0kxs7SF2Xhguu/e4pGLURi9VxSiVMAfz4NbcpjUITIyg18
aYVMWLFPYn0fc9vKEnTOUrurXNvaMJ+qN2ScckDiPSUsvtE+ZJJtdszedf81pLB2vFGiYlbMJZHU
YLIBs3nRluPnEAtSTpGCHKaHy27zXQDzbO/jgzFLO73+lG79Ti8qdPCp9F9Kqu186w1eng3MV6y8
ZIiGcI4/qjdVAOHVdmnorsHYIy5tQvjBymCu7cvXHuJegD01kjNOwVOV7Q0EZYdnbO6E8gx88SDx
Myckz4V780u/W33d+LyLnXFir+Tftg4LuY4d9gLFUcAL7sm/2C2urgM8Y6G6wAuyOZrDjs35ThTs
V9qgCpz1Q2Y245EpDPSjLYy/xsHl16OInTrD+jJ2mJRubvDcGbKyOsHPS8zyHIoBLomwQdklp+Cj
phrHPm6S0iQp+DRTsa4lELU4sh8ess1i6OI9e+xcRP+imsND2facra+9Dk/pax0qc3Vy6sO3495p
lNEY2daJySQY0ejkyLLSHEqnsY2ntYrPoJDz0InPpMdLq/pg9bRgAvlKYy+I1fuxbZYSdq83Y4CT
SWdCFP/7adpEIU4oV97sKhyOW81WBn0GsdL8NvB4hiApaSK5I8qezLduGT+Q2GZKOECcPeL8IwrA
co+HjBsVsLRePLEtvK7loF4qJKY46wumuSItcDfWD+NqLJO3Dtb8+qkmpJmXblmABQOXOH+Qb2pO
8Gn10Sw++cn7fZV7SOfh4lQLSCr76nXkjBnEEIOG4dAA+BGpS+PQMGgC3GCcZ0KX413+NVYsFpqr
6jiE2kwQDCigEPrgS8mX00HiYoy0VW/tbN1W865QmrRWxHICHhtHqVGybVi02ke1G0BkbXuAWhTH
seExlshKHluGLsfbhKY49cK/o69BVgzKLYLtSRx8fyLq9LergNjg53zOKESLa6IsDJvpIbooyPd4
pdsHmauRM3gbW/eZat8ySNy4GdK8pwy+BQeWfi1XBypY0BET8SNskp4THLsRx/48nejf0jHhc4ib
aLQ57K/f48pB0gwUZHlSxcCWyCR7MOkk2cqnhfGQSEDMCwJJsCUre3neRFa2iiSkvu434h/ArlYz
tHpuz84QdWEuXklBqdTFha4yKIkEfgP7sxBbPlg3kJEmrc2ZgC2QpBvgFNTuV/wXB6uWdBSGGycy
MmPeJJthbnULYlyiX3yAitkHotLzmlqypigt+CSnL7LpShi3G59PU98jwO8i2jtgjTHsHRSgNdFc
lv/pPGYaihP/Gw3aFmbfcbncKuTN8/lVfRG0noFVha3FhGf8oNeYISQ3Q6QYPFOIBRmnLXy3ZI0U
GemsfZnZ6/MsAuN7k8dSdWhMVKZh9E1FBUkmPJJrx3s62OU/cW5TLF+dXnJCnUKj5VuYVWyd5IGn
q0gBFrkpcLl3f/221sCLYG1FwnLhhs3xev22N7hA5bHUXErPCmEr9Pq+1/GYHL0CLUkeOjS17NwC
zhUELQkKkFrUK8Rrdo7Zwl/RWWZB9aotSTsrD+WBgYxWwipFwlRP2FLMka3KNB0lEJX44kNJ1OIr
4FMX0mHFVA+E5s2lbmnuV60x+BSQv+Bb0pmd3UDjap/4P/U4d+FCzYLGHP5GQjQI5FO9C5j/LvjR
sdfkbjAKLpQPgRyBQDtHfx/vdrEWE8ZM0rRgntBY3HzVkld8ZKPpJaZWVKWGx+JOAR5stjUy2Qig
53XptiXw69mSzoWQBD3+Y2lwwihZuVMpzdjlJ1t2I36H1rqDUZVdO/QwzFLPnuyxsUDb4C9bzy6V
U9xkKR+JlWu9OIu1Iw8mje8wjkX8ZVQYCjQqcDB+tdcdP20SpkwoHx82CHI8prbCJJjwIK4fT1Dk
2knkqpD1M6gAdj1Fa5dtKbz1jGC/XVanpOQb+Q079F57utbvsCmhBfMYpwmBRL9gy/1PKrdXnXxI
38n79BIB0g8Ycysxip3AQRcS0jtFizvxpGbtOZRlocT9BFNOYYpc0+QyRVkELmJ5y4UhCsb9xe/8
rWq6SVOZFdVUqbZfPweYTN3dI+u8ZRadoq5MS57h41F5iO59TschSn7fPs0SS4ONvaqPd7HxFOZs
FdTn+PHK3GkS/w6h3wFx0tCYnniOZAqTyljoYW9hnAbhb3gf9tKLRCPmc6SlK9LByp6hkvwCER3j
l9hx9xIemz25EVBw71xn2nHpPoYEycLuEzhrMiYIIddYTXv6ncw4h1dyizu0koGMijePMOT/V7eh
dPcNGV6rt8FORdNZBcHqYRK2M+hN23/ApSpCZ02L7qKdm+fidIEnJOiuPxqzpZx9uQUo0GPbNLJR
u4thzDAGszJDz0JfUopwOla0vQJ65guVyIfuog7MN8YtzDwaXMB5c0Wh6na8ft/aQem7zIY4wdh7
ggu2jGpFc+LpNBX79rOxsQtb49j2MpDbhvDTbRRTPeUYCzWUDsT1VNgACzqabHqkGdm/aZrsEYOI
29fe6C9kM3gGFO3zQIJ+n7sldJzzUNyKZNWmn+5Sgu2YlPRU0Lgvapj3s/vtWUOPaqi0zIZxLOxl
WvdfeURmxOdNWMXQIXxMoDzvnCizOcF+vzpDThW5NR2pHAs2eIz1HyhN7g3SkcbYmHZ2haPoIX2n
tK1rwyFmZ1Pt1ZTpLSS9hVRq5vtbOKaLlnJzcoYB38bAaoJKaEorI5RrFh3bFEjK4MW/j0Gj5hm3
OKFbvByX7FHhz4wR03QaCUblc6ewqa+m55ew4h78XLguf0Q4Q8GfQV0VL0IA+dUwge1coX+J1gZe
kX2EgzA/LC0n0yHyEEDHS6srS+7JhiuOYRjkM08FgV0ZMLC+ptSm2TyuvJz3sMlTyd7KXHG6Wiou
4XGB75V6j0l3iUEsPPmHzc07IOT7W+/xaLEfxJOHjbA11m1fdPHH+KYsCuaL/ai9ajl/poqYjcdz
kom5VpprGQfUqOMnTWAaiuM1JIPgj+Z00pDAkKj4K0nRyXZVGuRzXAyTlA1OY5p8rpD0eXmuCDUo
M6jdaQmA+DuFVCYFVP1Mj8Vn3QdMa5dEf4kycShNfXwRFaDVN0ffqCg7Rr1Csj2ZzxgEF2wxLuDa
c4f0/I+hT+5Eq8163ANEpkDTDGgMQtoZ+OqPKepkPKwAtMaWielkaOPZTeHPXxkbIMj2A29WtbEu
BGdw6comevagzJHt1TNq5Qvi+ypR+wMIcaAHppKwiX5qwNg1sF/wG/ZxyXxKV3GEEdKUe3QC0RRJ
ng2XnsoRkLd+ZtMtkkoSC9qUipzUqj2TnkDyujvAZ6mvB3ClrS0VyahFnEugCpkHGsnLY/NcwEQf
UTjGfl+BnsdHBNSXIBLyDBoXGxJYAP2fJ0bppKtLf4qR5e9JCxFdBs2zY2Lyf8541CQo26zQFO5D
7R9YpGvckMYxUeAbh/ign9un5ABC2Jt6AoULfgXmFIOcuRHr0LyQIumVspWNS3v0OOsN4dGETnkQ
NZuK8Ve5dtIk0BY6nImuGMvValWwjRN+tfblqHRpilHWl5yTl5DIk6WHtjRTLOOBiKA2PaLpcztO
QdU0NHFXtIq9oDuTBIh+0/9QifFTkorzB/LaZI9mL/q2u7jexwDqtoRNUTAwJH5yeaJb/0CznKHm
qJO45tV/i4akFFYIcfQ8UiVT6fOshb/86EEgdhkHof52CXiq2XmVmw5pMwcviTmJGGi1kqYwAbjN
V34ZzvVqAGb6ErHgvtFCV7ESGrgFr17cp3WyBnQeZQR1nLJL6uSrdWGcDC/lp7ZCqm0c0BKDXNbL
FNYpW8yHJQICaCvzUNyDroqoaq1m+s0E6x19LiQuAKbxEPrLvFw5xhF0pt8MXRPE7JIwElOecBuN
T+ULhYQc099fEMPTB26CEm+L8t7o0RhuRXvzvVwMXl/vWsA5N3Ucv7yzp6s6xRmx3oZROJJmsnhy
ADtxdgwSHSUQjyFDjXu8nwTQnFFnbm55PAGnPgTgpKaEutszTG6eWwfiQO1syIwjjIteHxJ0tuRH
5B5JQGZjypV3dXymcxHLRTk/vEb/7PL4p3+wF8j4Q8aSFczNZCN1bw6h/a9mD1YT7+XZuth6DXgk
jU3JRtMVnkcv2DeN3RJ6psxFm0h8c6uHsKXDTbfxOSv2KQNcQSP7PYdOSG2fabfzZKBPcbDYYgBX
W3k0qBaGogwjt8XWLCWWYthkZkpkzB4F/PGrjyH1tUq8Go1Bw9jRKnAdwK9w/zI2IjODKkV2Pl7U
/Ue2N8yXuu7OSn5E2ll6PD0kUad4ILdPqZTh/T7V+DsltPJQ1VSA7qDU
`protect end_protected
