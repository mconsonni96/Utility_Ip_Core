`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
RFNWQ3O9brqj72Wegk+N5dzgRf8TbaatmAcfOKtUFPU+tjSpdDZR0CXGs++uI3stUTCF55LPqXbo
FGeHkGeW2b49CQni0xoDH4g3hHTr/G7WttFqfMUD7OuR+JD2hJ1KYblQWSGSg9U/ScvId6qWF5ya
k2zcthiqCenCJpJzwRk5FN/cryj4e9HuiKZ87fp0mu10BPzmVQcVw6mrkWspPLHHmcXcj91uxOjw
iYOXIybW0YM9C8uEoTVNmSJLiIO5e0bkOAH/WA/xrxa2IG7faOhQdeeJCX7DYK3X8zCnweDZkc9D
e/ZHBv/rSsJ1NjwuYmpt89sKyJ0FbAbT7RR5Nw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="iTCoY9IR/2liliDmmZ8UoeSuh3PrHBLiDRyxG1TUpHc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 385344)
`protect data_block
u8mxi7twYh2OH1Cclt9D5Y1QZ32yWjwzDlBJNeYhSfE33yRONfTK/501s3o5gpIPtvJoS4mLO8uB
mHn6Zbs1C2b148OJdUEPiKwVRNWqCeM0dq2QjbkRKK7s9w0f80aSRbrWRWZ5wFfEaGLYWEYhwsTM
hgDAELFgkHtNshvXHKo0fZMPkwPuTnrmmGH9JLj3AruZXVGEjRrXwHx/mOXCptgHchGJ4nDGDV6a
0Wf9RnZswSl8R2c1He/xvWN/sI87GBjlxUOu4ReOMKRlCV1cnsjotYTP+uSpSEnr0Ox13P/bEELA
Vn3srQfmOYRjBoDLXDxNm6fiHgSKGhnEjzjkJ5hRHPb2i7T1bBFXmAJSgftYbUng7aMOHHW5zzik
G/18rlPEraILYHMh00bNtvG9b6JzZssvlabI+FyGEMbUfRgFflzKEQkTvYbVFdpXh/QcgbByaD9B
wLRq+NbgFkXa4m/aqV6wVCzWpPFAR+BMD9J56LUENUx8xpdQDlaQ2o7Y0hoLmy9wKGMCoucaKckG
E+zAduYyTg+Kso6uLvvEnc9JQNEeFHdGydemfwqpcgfjiZiEgyzTxVRxJ9UE/TvO1VT9ek5liKwM
LD8OMMUYCmEY6q7TLJjlZlNbVrd/ky4x1s+iwiJXoq+SWAGL3pLu3NyG4BEPSkogXdAWol3nH/lC
QhC9wdJxuBFbDXx+ek9BHjxKT1XrKND4yZPtWtw2skEmdNjSUSWJ5t4Smn7/uqJlR+gjh9BLC0tR
/qINZ0s4mBAjZfJwqSCCeCAOsZAbyOM6b7yN5Ef4gv4r7jjJbhJ8lDP8EFDC4Feln3D4PicU9v9h
q7FjrkBqnxFDDj1uv6XOUm2gQ7JQd0yoC2M4JFmtvZ3PkVt0nWlG7qmLm/967lYnhvx5MpdGrOWA
jxFTMQcWAj0N1BZl+IG6yLcEqYeRF4Xhd470yT59bvBeyjt5OAssneNns4GkxK1QQztx4bTqBa52
Y8ElpJYUoX948uJfi7ZwPnTMrTfNZEiqyKYDQYOKOYwejPQ11UmNGs8f/Eoaoma1HvD51vW7Z7EI
j5DlgY19Cu0LtWDTebnujAa8mDhk4x9fpKbng9iOT7UuqIBTHpcyaTVzPl9UeoR7Gfj7G+wvvWjZ
/SbOmdDiFgh8BmiUbtkQOUGsptl0MvrW1DuVHQia7zF8Qj5VsyDkKEpkUs5zmT70b7Z5Myxzenbb
cW/s5ZdTuzUHvAW8RRkeDhRwSUAsH8znyOCbHzq8aSFmjGXo29dcEtrbNOzow6mHCdZ0qtVplYnU
qGwsDeNwt+f6W5ZZOtrGyNOhL7Yjvwg+vRXk+Kp6fXmSv8M/4e0Wdc6oKHXUr5hz+b0tRK3ulY6J
mN5n0ujbeCGBIJGrUEVVZUA9yYYpUiXFUTR6/Ocl6z86cGsOPToxd8KK+yvjsDvEH5hMKYEBZHzd
LQDnm2ZPJRWz5xDDlW7QJsebtzmRL/sHldp6fn369S4NvOHHsgXl+tcCdywE6LWSpxzEqq8DQqKd
gmN4FfIoLC3fjbstROJcfFNjFtgU3YsMdYoUcPHNsZYFkn//mheJez+p1oGsaAhzlSXPT0AxwaCh
SJrY/wTBK6E0BmFzg0J9jaMmzoWm2RxN39oBY31lYrtDMmWr7zmvVFIIpXnksNiglhgZ5EUgq9ds
JMYD1aamlaSHJBLLEaeDmn+aqyx7yx/y01lCbBCYa0mqz1LxnCcoeDDB/m3UQEQdeaLd8VOLXDOW
iG1ejq4WoxK7ObDPmse1tCnuvbIuTAUCmzlFoI94Cbqcbdx3KoV590ZkfJ+pfPZ5rkSsaeyuntFz
q+HtxRvhqsp5sjvayZuvkdA8jBIrT3HrllS6sOdOK+ocQRKRQXLKALiX3IxMIfZYIhObe8dEI4sn
gUc8bn6nUzuv67b+yDyWgUejV9+joh7jj/6zRQlzh7ZGL9nqd9ydtc6pAfyoVnRxfEHcJZHjjDOm
S/d6/0umdK0XQsNCHKCixk5PyJU3M6sLLWTFc7FuEmW9m6gPj4AHJK7Amo8WLTHvcJIA/pz/kxcW
SEcClzQ6um22GCdgs9JcGz4WerCP3K6Gux81sf3m/lAfndWyi9LuvocqWeDwpGIH6Dd8RUOUiuoc
4CEFjKUHjYYSBu/OE/druT9jmT97r87SbqgAcjOfFxkGiqEcdSjdSYbOF8B1EVbjK0q6izcbpWl8
9VGgo0BaxihHmWq1nfADf6xEXkXY6X+Qw0DJbd7s9samF7d1O4Ueo1ZOiFNuiyHlkl56qtmkTCyH
heKCIO+7i4ruqBM5zDS6gNduHyRhjHfaQQoNsDfKeq9VEJjp8LomvVGYTkcncEpgiwPwR7gcPNSI
1UOuNqVJTr1cQcPjvUakWsWlZExvS209nwLJ/OLSYUFKxPRfAveb+FzBhG+qSDh3TEcuI5CGE0IJ
fI3uPeCj8tWH1ChHdGGpqCbovElhP+b1HZ2VZXU8Uj0nPBtEio+KNFSB4m93kw/6tMz1oT9F1HVy
q0D8LTlUJ5IEGHXjxjPwRkSZxlhSbquu4tEKCwY4k2UhWdcQky9sqP4IMnslAvxR8guhdejeHVxY
IZi+O2jon7rMmshcLDUi82jZCu26a7r/GMlq8OKeynZdf/njJZpDZawW4wfli3dzlxP4HcRfup5q
Chi1YcbGDZN+ZwBhPRIfapsMMlzxkCm52dogSDbVGZ71e3MaWlIGatRJBnr0/MXu96L7LiIXddvp
eJhfx6MjS2vkb4KDQR7vu1StMbJcmOrbVYvk2QeclqiLOUByiJvIt9O+gV9xzW4pzh4Zbt0b0TcF
nBeoJmItfPsfonkaFdbQuko+ic/Mj+WHV52UbRiTKfI4fsqWpUjo0PqRgKovxdZxv5Z39iTu3fx3
WfJx0g8+B5PQ5Ata6HgI/XSQgefUzAEvcAbXr+kkOIJNZaS5QPZ1IgmR6ZKRdy08OCnz7DNQTRPC
KDFPR66Yty1wJa98jU6tAPDO3hzvODiIbxY1XFwfJRYCUg2Hw9KhyXUX4mbIQwSM5RS0BcTCqzaU
Nuyyulgy4XpoL7rTrQISy+jH2sv9jL8030IVmddZdUf2GGYqFo4qK4GG3TLk3gy/id0STWekBKor
rN2756EpglVNVEc/3+CYhU9agcJnPfExnWjVOTWvxRKbQiGf9h5X/cc8SKq/9kEScw8NNqY0bMqc
uuzP7LWc5MM+jArSiyQWFiyZmMZyIjtfBs6UiiP+faIkKje1/nm3wx2EZ/BioEEbOlPISotx5Tmf
5EIQV5epCSaynKsbNRwhaDJIdAhcGOC0aGKMrPYXz5Pcw8NITaw3qMS3jvIEg4E1sDDjATUg1Xt6
aMOsmnyq6dyaUXbiH6z/X6RSE+o8SfXSSAsTweIaqf+RDZXGvqQHwEnWPc3XnODbhH5+ahHyj+Je
xfBrkcHrqdUKGvVRiSJVCryEp/iph3f7fXepOrhN96W49FcwnbSYdSZS6JodlBlfeo/jsDZMxAPT
BZ3fcAWhvvcTLmo0Mst+HpMopUVUpEvFykvMiMt9bHez+WNPsFH4Vx87bx7oVpnhAqKaTMcC1kMs
Ujf1MZTuYlFBeadFoR2exyqThlQUtDlRo0M9mSNd+2M50rvYbuH+jSXX0MpnIPhTERmPNs6f8OCf
igRARIxd1jmlYEqBkyV48SCT8nxG391dqC55K7XvB/7HXmiXEZm+g8wLqO0XpJEJLyUg4hydnHg0
By9hudx+wmI3SmGk+3y0dbk/zcWRho5fNWzX7wjPO7W7B3WkJOexPDuqnSdDSvurdgfdhblddyvr
BL+Jb04bQ4Oq08BH05wcTkSKwkpCdo2+OVz+h67sbr1lbMfKNolvR3a3yZe8mMgeVt0GSnKqfWBZ
33hgHyAqYxbRjVhCrSRUvi2LzZo4HGnvFaq4oyDWXJwJAjjYmArtoJyD4Gb9zhsq9XJ059GSxKZ7
+ec/O0YMuh2kfadnf0lhh4jbMyYu+/VmBwMBNjMHh1xXj405cjl44ND11Yf6I5GSgrfIhPWnvqZp
eYx5XW0GzDXL0QZ2WQNwTEEH4cybfz7IQDfQ8ovGxyY00a/sxOOrodAq9B4QyOXrreP/btmbhu3q
Ku9AO7OzJmqhnfhWyqfDCmMRBgvYI5NEyYq2lLpC+/2IP82xfRLFNYY/eSIQiV0N8z1jwgNXWH52
mtwL9IVZgwTkrwlEowyZbVLA6pYksoUS7YlnqSqsHxbDg+u/L8jFZlgWF/Ilg8EO31CrSSiHsc/O
GODe4pANesy0nzsfGCfJ/uc2eSfX0GHj3WSgU3UJQZroqpqTfcxuuoyxIz4xM+C3hsr49QM3N0wu
HIC334rWdX8vGPTODczzQprx6svDm9/VledDmD870rS+h36dmsOi3E7M6g8+d8g0DWc/OTKBtDeN
QKwLDn2/JUoybO0bjjVHF9rIWJzkvJwZECvy1GlCP+T/gisCm7YcXtThdug8Pox/H8q/h6jDvKnb
kTLngVpKdqWRYWa9K4E/kzVcqgpKdJeExn8jRtQxhMBoYoNTlgSiKNYWTlzOx6CWe0VIoKgBz076
Iea4SN0R806/qiGhICsZFgDIswFppyR8ivvnvyLTHHSWcP7NLXbn2YgbjIo7gbiT4uw8RvsfXByB
AhV8IbTJnXyjwne9ffryKJ+QlBtckMFmUSWFwefFuFjEG3a60Bga19J62eNxEW/VtXsonz1r6HJp
OPwMJg2srAgTbsVRoNZR6UOo7hzq+E+fcDM3l8FMCD+uX72wqhuAn7F+w70qX6i6R+2Tum64Vesc
rqn9nNf7e+dFl80DFRbAMYtgK148Q2qHp5xKHYVg0LiwgC5EEfBgV1c9ZZxFohCl5sqxj9CSlBzj
QnSaspmk4+C0FZLvYUcNgSaCYgHEeClsdBznNK7ptOk8ft+f27uSD7Uvm+iqFmeUV11TN4iOGACv
atKEBRTsv9GU1vheF3xQHAEt5iyuIDhCznQpyNfgu6+96SfGO1AYzrhhSGfPSFw1RyaCWKFSblCF
42Dvm/yEMSmiv9yH6CYMpctgnhpYZe4GeT7WpwdK2gV96ER0ZpmVWaLCQ8qx3U42NPNNQNj9sojl
I427+yUtU0rqYN5KIFL3j/8sYXSrEcI68PXykgy9ld4Ap4l6Iek6zP19ojFV7mV1pg/0Z+Kn4h3P
0ry14aW2FWcIK69B5r3n1pmXI01110DGvg9N2eSbXjrSuAjwklWAME/mtSfYN4TpsO9o5wN34UDM
eoUSI45ftSBT5NJdbSm3jiss5Vf+N7AlCwwyTbWc8wTVhZzMI4a4yZ8ZhAqMaJ4ZkNdSO/TRi/iu
MIok4rGU0jodU4hnYpT11wuVWZ5qLuy/hEfN7gy1/8r/CcM3RLTbJ1IV1XLW314S7lWn+yucgFPW
24OaX8gSJtmPG98RMTXoDUqLm38yDCEucIh99drnmIGPPPvLULuljYo7L29XPUqzNTyqCk0DHq2Y
+CQ4OzU6AEAqjsCOHx1XEmRS/2jXw7NUBD8KK1iVxxNeMRQm5ZpRjqPkzNqHYbBaeZwtsd8XBavF
DNVxtJ5hUVcDdV7kF9z2+ptdsDBIh6D2NE6SbQ8oAXg/c/Em6UPEsdLCkJIZEtueVCjSoL7xgAb+
YxB+e3y7tE9m8NP4WhgPEYIs9PvIa8uQxKWd0CCy9BMYzwZ6zAa07I2svx5FXF4dvI3AWAdT3HUG
UO+yVqbrbXPZRbxO5cdl/CgmfRthXxWJ9hVinPDDxIjDCjVtYpSBE+wL9zmqg/zoOgmy8eqESvRP
84GO5m8exQM7KmXSj1jTp699KBeTvbQA8ZSq7gJAJiSJ/Vfv2FoR7onxa01c7NTZ0nyiOb/UeP7E
T3OFsO2wFxjif8a1nBjo19SeWQAuVGCIFUbChsr6KAkSggVfn/eZZR5+jl+M6HTtg32QcEeg+OA7
tY34YLKXmujN9X3gqeVIfJprwuRkk0zK1o2TU7rfYYWQ+mMF09RD5H+j1TMSFyGvs8qGM3rlQxQY
c8GowRh3jzjPUVSel6/JtJSD5qbhzEeINR5OuCT+lTSwFGno1LJjw32npsiwnUoyx1g2Uhv1aFDl
q/REM4L5FF1SqZ+v2mES3VLfsTWNtOzj8nENA5pXsVcgCU/OaBZx8DJOjL1KphU2z1Y/HE7902PO
S8hPJKGp9GULdMQn1uvOcT/uSxyhw9kj4bZzk6U8h07ybPxyo7nNL9tUDgQ04tymBRvBUvBxz1/w
BfQRyj/rXlBMvoqzGqjJcABko3R4V9T8ieWssu6jJHEtbv57f8K4kDnyjhmgVq6Ncl36quFLSLSd
Xm5UZUHkWquFEv6LID80fdkNBWsDg1ynbIKM8Vn7rOXIZ1iXRztCuS9bGSYtU8knzIFyRveM0rIH
KTzmC3niWWMTqFyZrp5kfql/5w5iOQsF1T9DSZyropxQCMBJyX3c1DfFtJ0DPVAtJ3l6rLtiM2dq
px7kDOVKtl4pzjxrW+7Mf+Y/V4M5NjPuAtQMFNx8GKYVX6BdvpZJSBYkNvqay5SsiAmZIWq05dD5
3bdO+dsYBQwsM57nej91HHSf7ZDgyKV5WhkBwRV8A/0orgRUKpmC3OJRc1uHyTxD2tYhdQF5C23V
mZ22rE+PVpV3fkEsoVxkX0VzZRJAHGCSk2DqXZX9ihGViT6AHRIwa6NAjnhq3V/DxMoHNtlzuZbO
KQEF8u3X4mT0JceArnAeg2CbjKtqJYEKEuCr6Zk70QV+8sVVQLj5jsHAL9aLtHhQCp+tRXU6vKXw
fwn1Du9SS/US89S59e7yZWSrv3giXLGlC2S4cWvr2CWrNEoamjwTNnpJDam4U2L23pKSICZQhGw1
/35EWN84UPkyh4BAVzlkv5gP9shTbUTGhWmL5q5tiggB6t8zSJZuXUnjRyFkGxXnvgR4MSr1VIly
9jYVjif8vTaPngLJZqM8JBqwpwuep/XvpyVhJJdClrbqJcakzPyHOVxULqQeaDZHAI1obGJEP3SJ
42gSOHyTTVZvEGjek4ulRsuA0+brcaJpUeYr1mLYe+8EQiNMFQ8QdnL2aKdA6SyJP2pRdykZ8oFG
X3lByhtqlOEplLjS3weiR/aRGuTSjMneQYVPVk3qeQwDh0FH/lyvGwJD7yWOowbxPylDafw0RrNH
R/dh7HjURkB0gb2q0MPl+SlJUDH5TxjjGgrCvpHG1Iu2etg5TjGb7i7ivXRDJDvR69B6QitiVRVW
sQl4roc86K0pdKWMxph1sMcfcvrPFfC/YJJKx3TWl3e6pyMWViz5Om4wn8MHPa3lMPDeG6zqOOmh
yMEfdDHp3HQBvcAgPy7fUXqMmau1yU0I+ogDmj+6ESPQ+WP6LQ0p0FRbYChO3lRfq+anzpUvtm2l
Ylub82HIWInRhBCMCQ6AoIs5wGg15FroIuT/mYjR2mLgmozzZM0Pntx0wWPL6DiTpH/M5qsNNR3z
bQWrk4sc9NaQgOccd4g6gKFjf76quBh3y7WGCev+SpMt82+7wmmvA2k21WZhb6dQ9Vw7F7KoChlf
WRk7NW1oTfX+uvNM3rV27NFnco2ChWI/NDQQXeeSsD+XXDcoDxQqpFOm1gTtHfupOPGtViNlmV5E
Fo9YhXPHpOMBk+KHcGbUzYONJftHlmPHfc3gzgUvvkCrJa4o9OhDrgLTfgIqQJkLXuXO4uO88PrY
YRuOFpRKCoJMvYMOJbVlulgAnTjl6o6l0mSnsPc/3LREzGFGCrSDgukxoSZDeugzyVmEf9AdZZcC
kfaqkj2FEX1Hm5NQTgFj9JXzMSrzWLEtLkEONK0iQ5XONFvDpp/a4SVcfIA320RzKwKU/upXnPO/
7RfoTKrWN6/dIjdRjzoJk33OF6i05W8tPpVXoFykAqA6Msc01RRui5Hq5YjyJqNM6uFeNW/A8edU
2LOTNZu/1Zucicxq1RRFPeWpCJpUr8la4ELIUwDwsXLA0bfhq3v6ZpwrzprlPQ8wqXACOUr6Crih
6d0vk596U0nyXzHXY+g/FdZ1+GpE9muGMDpT7eqMCnPZ3gNmgQGeI/4L8nr0nlVgKTpIA8LRfH7A
ySmjbFy8CVX04T0F1E3SM7VTSvWDct2fXOYTyxI+ExduwUiHNIt2evhOQlBhH/VyGnIj2YHP+Btz
TyrSZw4do5/0+5MyH5BRvisg4KKEYdrAYQf3OS6s77lIj906OsCrz+ZB+GQb9+R2WU/s1ezT5MQJ
ecppmrEiAnhOvrEFa7eRLLDEwl8GBJ/5xb29jNKOha56n3Q6YeqwADv7KiJb9rVsQmljbIoFbHMf
g5oZkcGXqfaTHyI7uHgw5FuZm0ElglEu5bG6s3o5NdclYqTLtE3319RaKjmOEqWa9C0Ai9ZQt5vE
IGSINviqkFVZbco2/1wDlov5Nu/fRrm3YoUdjg5H3XlNNCBLCtrfvE4FnFCtE4+j1XKiwr1zN7di
m6kDti01HXgSEWziWffFrgZep8Gw/1Lq9JwuY+BRn4JdtEwdgJYVFkAo5JOZ1w5b+4gD1jaE162A
BHdGekFevb/p5Ifr065yP6RC/B55+bHkPOaA/iDNWSHvEisTt6LjzCB5tisb/1+ds3HbrNZvpZrm
pUDMGq1OL3dUhU92oGZPIaZTh8Y/eHunnwiRGgGMGUNgCFnPtaOPlSMleztS1Bv5I2aa47zDpxVV
HwiVnUfCFn5wkcvkRJUzAubBscJio2edBYiEiubG5CWnzXWBUiI0WUQCh/m/qtIEoMFef2sGR2sS
+rnm8/qT7QYXgxkWq24kPvL28obf9hlo6Ngp4T+LZunrTlUsJG+qgYGwoB339VjyvM4zdeq5TNnB
p9Cfir6TUflu3mBTuBkC3QTQ2mKq9vyW2Kh+1YnCKemLX7cNhW8tGlTaPVgP+XqN9AKedoG05A7L
TmgoiOralWZ8GfrrSoLv0TCsByZigxKkMC3B6gOS1MbFGTdnSaMsFgyUoLtTG7eDsdDdxDMnjY36
Kx43A3eVKidXRRXmutSwdUv66ioXhk+oVeDFWdenyY6/CVFk4jM0L364uSLxo+ZUKn6cUFPXfc3J
tG3g5e0pDpzx84noPuHacD95nsXw2SdsiEF/IXjTWOrGluowSWJanXd3tYgGg3dpk8utxsb7bJ8C
rlUsX96uyP8Ljyw0ZapQPDsi2D2tEh4RTJaLiRlRDDzXHu0ts/AnJd0ycMa1mVzBRsxafsJl1+sY
G9T/xl9qKUcy8tV1NJaund6qGFuUL2zjqg8v/9C3CfPSLdMu5sSBuZiH/MvB5N4iP7ddGG7svkoj
ALJNVgyf1YNyNC3IsW6LE72Kcvw/tX5QQk8SH+RZjGJ/MSxzV256e1znvcGaDAcMDsLfnB0lo6ol
L8K4SVmTjyz18+g58KmCAo80xKuWxA4PyPydsdZvSz1aq+O9ylrLjMRt7tL0NQlq9XOJ5+5Nc6fl
+1/76V0UxzRqFyH19RuQy5AdJagkN7y/bWPoia+Lpdxq28GsGBWhVYfx1nJjH9jrvyLDq6HrHy9v
m8k6DVXRui9xgrxAias7z3zHcuBBVtcvX16ySPMymh29x0AIKmRThAvhYyuZw1J3kiCtHevMn4jO
OkQz1sLWlAv92trPJTYA4JB7EPzhij7ANphwVVK1xRGcGsPf52Mt6xVllEu7vPu/Buz65KUkzi/k
VUbBbYKQZD8NqyxwU+JHLscr7l3vZtnj3QN0YVHcOitGlxXvghJRy8hwtID1g5FrntJ+6TQ8ghKV
lfM/uQYeNuJ7VMM6XEj9fRjB+HkRcnUezjcdcLEzGt1p/2h2NwTlXoJIdtfYR795GBVI7SSfSNie
XwjX73u7qqXRd9wo9Eg4WqhM9BZH0lFqR9mrV/xFXA+LWYfDDo13hfroqrWilS5A8vGG/abUZXKk
VqwGYIeqNpZTKkqg3yQfKQKVPjAUy9fCGzK6OGNOruPk9rmm05d7fLyguSiac3DbPTxTEVwuoN3J
TouLrQ+2Fo9dxRitYY4j1+Q7roxO132RGnXWp4BGYW3V0rX2aIBrUo2bXgzyNARs2i0/8xlUKv3e
w6tVfYMDzyhz2+kVFfMy+Jf8afOaQ++YXnau8vp/JXmQ8qVcgEeaIVRBrv+0XDkY6gvltVAL9VFV
ZXLCVadJ1LrizJV5+jN7e3/haK+EB9iQbBm6Vpuq/ERxexdw/AxMHSjXv2jQJGX2qKuEY9jDAAx7
WLHicIg74IWcLvKXdd1ikhGso5WqsL4j5CV1YdZi8Siwqu6sstQSOnjfXCbMgxllsB3TRVSrkc3B
rWzq+RAqQc+GkP72Tj48q4DLJyITfW6LP+im8NrXWAmXJKDlGgdIhRpthEesRiaNBlO18qvWfzGQ
pc68VGFOGW2CpS+oOXcjBsXBP9UcxgGWmcROKwKEjh87tG+ezjmUVsfmncmXxAHeEbdPLZp8skXW
scybt9llCiIwB9fy8L5U9LfYg0CmlPNdUQZtwkB1hSLJ4GfIz5OTdZP1xDCNCc6WlKJGcSquk/d1
pljxp1j0kNSNfC1ONaYr4903joUlwFSQ3WwBThau8Q45NdXAmqoeI+7fPOLhM0KqLTyyWotvrFd5
NpnHtoherjMRT+lWVLGEPNhIHm1Md6LfyiR6l1/b/AFNv4efwyPmWqRIvS8s/U5UAPMNqY0H6lWt
N2C0cFj1pF4O3/il/qG9HvA9H/LKIuwaPn6dZm+tQxPK9Lw3V35MzBMySOfP/+DIb1vpIZXTQB9I
R8sT4eIznddHbW/2QGZZvGbaoVGCDTgRTPNIFRgCsZk34I0XmgJSeULgxvkBRGWqRP+lKRcKnVLc
1LB0P7x/bGRX5yGtIXhB/2kbv1dUxHF1Y/g2GTrZDYinvLRBipOKG8luoKonGp05D9RPe9ljUSuC
CjrDi3xQSOZ6GKCjNlNP/67pT3NifFP5usisYHzlKflFH1FRr3FwZvzF/m68vP8v/sUC+eUD6Wvy
nVcR2sJYpZ7dgP2cRSei2taBnwXeXMoy3Qw297DeQhyquvL9/MtLqFHHg8l9bWLdgFKUzY53msT1
lKVYrkd92md1cDHftyYDk9whzXW5MyorK7KdMi7rkAImWieM7FtJSPKq1u4E6fJ5n6lOogm+DmUj
CXLL2T8e/RtcQzha0YnuahO1v5cJAbVPbTcc9Q1v5LVOdwoZ0JE1LIqBZae2TzyT/ee/SKTfYsav
8LeKqxe4R/A7qfNvZxmqEe7jcFVQlcDuDSwww7np0zseishOcQ5jbQsTFEHW7SzLgf7Z4yIdMmsM
zdOjaXzTavgS0Lze8FmnqnnqdfwZY3iyqtiAoiKGfpICQAUyxnJt5pqPqSFr3QMHaKR988F7FmaD
kO36PpB3u3mmfgYL3TWUdXol2WhWDUYbr7KobVQwU9twrV5MYOW5OEvEK0p8CJqjVoraEHwL4o1K
DmcrpcaLa0xQBjAfcLxaEGDJuDzCJzOxssodJkMtl379fC7drIsQQoO8qmc9TE+Fc5E9LGAQe+Ij
LYNqVVOb8uqOfACAYJX6dlX6WsEriHARsQ1+FsHsMqQ98uffO6keZ30nHlQf2Vtp8aKly6PjHtzy
adLR2cmlnYCw5p4yVMir4g9y+d6XLABxMm46R81/7iNZeboRipuY2K0zTu5hpaVBzVm8OqF38UnA
5KGaq35dhVHyyKIJrdTT/aq26SnqFbFOE+rGFZRmDnbTGwN9Kgbe8fD9R1vmAw6h2cMLZNtnqVZb
wu9Mxylg7IcsVvwVi7byI23cm+YBBb5WOI2gDJjgcLRhstupWjZGYBrjBClBmux2DYsS7Qzh1dta
aog1sJA1v0QfUoFNtV5QZ8vZHkWvuqPLte2NW7Z2fxxh6Fz7RXadK4TGnziNTLp03b9V3Xmw0Ksd
o6qORcM2uQ17PH5vw4QEeTH1789EtxHpFzUNr6FfxFZo8gXe95Ym8TUypnPDPHvUrScKdnWpRmrm
8XQVUKisuaJaST493Nqbni42Bmwl6hQWJ71vKOMLZr+FQcvLrikOnxyvVrdAfjC7XGJ74ymZ9Oj4
JOiUJIFsv5vGrdCTgPKUMoQu+/v0YKD3g7DfWLJCNQEk+BGbeO04CHnlKr8ror8NV5U5kz4tkJj4
Fu8zqo4JutzE/DtYz3MmoLy1aYay3aburqT9yMLjdO5gC7jZuxyhCg7HAIDfy62UPujK8w75Cj8o
A48vXbt3zakLcO1+sHYvTo8sLhoWNAhJlJOCh/dnyplIj9wm3JErzd4iZhDcLG9t81KEFeTfXmjW
Y1Jh0JrDxZ5eCAPTxi36h0B0xM5RF0KYKZfD3lWepeWfzfLPZEISES5M90uU0bzzOBQIPAsfbGYD
lW31T0adscLuSEUb83v97HzCEjbpnGM1HiUV26TXlLROUzkZxcXnX7tEkEKj/KWTNrZnH+cVHzEd
j41mVPIEYlTsHGRwLUW0Z97WGRsojTHcHMqEFjZLcEr5ju/74wRXLAKDHFqzI3Lu0JZg1e0hFXqz
7ZmctM6i7kGnE4qy3JW5dPHA9wOO8Gsd3GDo3HWJabDMuRMBjaa430suCXPtAU3pegAavEzdwyjC
+QoPQyBHabc2xgHAKhRnGHgQoGXtgh/+LWs8SlNpfyXEQIXJP6Ftx/jl5xyn4qYFT+9GbQIBTBHP
dCQcfch9UOrjfaE8tvmB7f0rQJybd1r6vq8N5D1mdcQVZxxCCsrrKhhoJXmeioJvr9NTJcv5nc8o
YehLSEV5ttmu26MqTBUrSfzF1UWrOEpZJaTF4gzbJFOh9D8AlmVGKumEmdK7a7Pq56Y5ZJq1KWNK
oy8dvd/nemLuSyKR6c2kdslz6B+xgWolzjEL3X/LehNg5AFCNzx0S/2PseK5BzWgN/JgA3sXh+QI
5bsV3CIFBDsGL8MLUYHqXHQqh9FH4q+cSASr+LSbcmKst+jotFNe9pJeFSDgLqWKtYdVuBRQ2ton
JhV044maEGR3j12+E+I2hzTC5QUiatJfzZUDbtzSHPotYql9SZtXo4KhP00a3u+ddPJOTQ7upYi1
PLR02O26/jMlw69Bti1j63fUEEHy7ugtqIfOH1YQ67Mw5rPIuTS4Z3Q3k8HbR5159HZbMjrQbpqv
iyCEQNjlJdtclKYtJ1rOVFnILckqvaHlSrKlrhWyByqP2QzNjm1kC1PcpccY+GaSg8TWrCSLAmJi
Bmh28DywjKy9akve3d5r05ExWxnZsOQkl4uwvLRdCa/qZoaaZS89E+WxmktClDrwJtj3yeHO4Gsw
0a2ZTE5fJJZZJ4fpbgR2yhSVlcQt3GnMh1a4DQwmqZle6zN5mty3fhu5vzYrog3VgGvF0lgPUhLW
Io0Vq8XI6SF8xOiyBoFwuRqStYoveID1qyID8yS2yqkoVcJv8s1aEmgi4S6R00vf6wPwlMNKNz8P
u7/FQfji9C7v4CcXb1/RGphsp8gPSAqmnvD0PZ2vdt89iMA9yfCe2tagcumNg6Mq2l2lnlOmwTdO
OMgnc62QV9G6cBobHj4nlhYOSCajz+bAHz6cy4K6Pyrh0xOiv2fddP66tO00/zsCIyo9sh4SB36x
pdIKLsToI6rJNNJthiPAI1ZfkjG3e4NAO0Acuzpg71/AZoLAXJ3DexjF2vWnXoOse4nmPzYsOrUO
x77bK1Y558uyqofICffrPm0qq6th/bFuZzIjFMyZBS+SnE4oKx7CvohVV4NDIGqLOBhahRTn3hdS
XWx5atWu7POvEgTz28U+cCvPZUW50zm9ChcfPs/bQGjGMJsAyDT/DGPlefmYjs/Q664ulQ1dKPGN
mKH+F22GiH3X4DDeNC07AxFVcnFx4kY2X0ungK19+z4D9KRW03xS84/B/XBCAnMxySm3vmSTQdmT
zNlYRjL460Co8ZKqXEHOK5MTL9LmOJWr5KfbzxQVDdujksSn05lNQHoI7is5ubMSsVHs8zz8nl18
hRwF0RHF+Xn+64fcJvKTcxDMFUOBDUNdA9nPzZhJZDZT+k8cDFaZ0zerXmvmt+ELN3yeGrBeH2ar
VJO1bpXY4mHp/ndCnS630yNhLlqDJFcOump4FokAA6+N7nUvzcSDIyMJcFjQLd87pJ98+kHs+WWc
rIq3SDRoWJRZ1ZksnC94TaFCCoY6Oo4AtD9Aivr/NUTvNemPMGVy+k+xvkwe67UE/kSuTuOWSUOu
jPkL6RgROAeAsVNKdeaNVH41BoApHKlTgvkSJ1rffhMuAp4ghER9/XMEnw+gsXZ8JkOkmuxbY/gE
uFFl0On5JywxZDyp2abywhWkkpg8d4zxv20kFZKS+gsJ8vrmigJhFgbTLJJ4JK0iIOiqzSZi42Wl
btC0DJyJttPwsif8i3/36jhv5EAvC+SCx+ChFZdKgdbKEtbVxKOIK0Y+1m/MLFjup6Jcic0jEmzI
Xw+k/sKmmUMIsH2aLjv0QyY4DZPnx0GbjCsyhrRNmWEEy45NldODH7/DUQyi0OKM7J940oepTC+v
Le/3zAqGjmxNjl/TgMduju/o7E0Zz5QltvsWlK6caj4eJc5f3hdzM3UP/meKWirQ4bCLCawsX0kD
iO/NrP8APSZE3Xvn1NRjAj87Uu9ievC4GF+BfZCBi4UUCU0ww27eZ5d2mUTUUiKrK7dnTEMrMzRX
qY+NYq1Yic8Y/4BFkWVo81+2skTKfIK8tlRLtSYX/0g55+wMabpSCjlaw76vVmVXWuOzk4qBP9+5
NFtluNQZUfa5fRjqclGEA6Rg5kWIF5qIlmRRjVX47yvignpWruS1JkWzPIx5x/UYXSa4RL2w55/Y
BtoJBW1Er4bztOVkEGx6I0VfBUUBQqquF+aVbBFR40doJYzYznLrkeznWsmlHUijNBuTKN6HY5Dd
sOWNAyoiGfs/ysQJbird31SHcACkOcz8rUy1avdQwrFmU4Q7Yo4sYBm7LaJOBJSFrpM+RH+ex3id
shXdfau6OoiNpikzqc6AiTX/tKDWBtO5zn/+brfTazUY/cxgd2WcVDNKEGjPIJ5ud1Pd9MDGyfR4
Iq0zZi5aT7Tqm2XQDOaPddFVWrW+Zkk2789TpO/gBSziIWYkb0aCydoJ8iLkbw80nhiXm25On4qG
iSyrxFkdF5AD/CFH5dmhQ3yhvHxuyKDeoaCosaG3oNki33bT6j2XOYkfpakB68zTJNYKSAY6TpCw
Q2s5Qwm+fqfqrghxnNzIhQzktNxXYi8uQuhYP4Jiw28OVx/i5oKbya34BgUgHrhTob43hAOXQvJr
z8R7LuQcW8cv7K5xvMkBRb5/8FW81nmsZegTkFvmNHWmxG0PxHLsJnznEn6ckylpsuZi4EJiVKHF
yHC9qmuWl+lk3nvuLFqfpkJxDWueLSKDtsbGW5eul61s+R9kVuCWFTE7ST7L/RICg3AKXJm30L2v
gQTJLr2Gxf2OU4rgT+iQcsUlYH2lcnZ1O+XLYfQjmCJkUJSRY6kilELqpFC6hjPD7I+Wklk/5efB
/nO4CI9jhWp1+meAgkfa76v8gY74SQ435GGzKugua0KYUphV08KBV2ETlwjtbdqHTTG3eLmsGkXY
/MwUCSn+UqwDGbFuBc3tGP0IrmXriJ6fiHk6c7tiBkp88zQGP2kKD3sHiP3GAWdzOfMOVi8UiUzr
KvJRbqS+ywHNnrlasnrZzLeP86zphJAwxiSEpfkcHDZomTdlYwy2tA0t3jxpbVA5j0vOIK+yKJbM
gvi10GFGkEjX7w61uATceFqme6PgE1/CSNE9yfyKnMK60BMfZ21WDwTjdGN/NnIzCr8DDdEhlf6E
izyTY1mLKLfeyMF30Vb//o60+qMe+zxWAISGmDvQuDKO9SpUbYXLxxYpPJE9uqYOK3xoE2RxDjZ2
D7kbZIcsELjb38O0HG2RbnvPcwznxbVUuL/MV3tQPOxa7NauBYsPs3fwQhxRlW68GtfAgacUgyNa
eh+4A76RGsbCF/pqcX1ciktfI6GU9pKoGDA1fuw/s9GuxJ/R1UyvdCFtHHhDnmd23ulQa9AaWT66
JT+dDEYDbB0lG30nHxm9tLQ5W994f3wC3DqtYYrT4BtrO0l7jcuarnbpYmyf3No42/kQCwXN+/ue
2zt0sbll0PAih3rKJxOrxMyrEx1m/s1Gnsx9Lo6F7W/dQyo/w+r5HfsGUYBZb7uXAthbefD+aB5R
/0mBKXflWz+S/p0/x2JdSM+QnLGUIANNmMDomZcBSkN9DGkmqeS+Neye725w7hgJY1soNLffYVm3
9nkF9TeavUUggR8lPwu/v+ahRKdnoy1iXgsJ7URbHt7QdJY3fRkicnSwONGyn6b5yvZJJWzIHog3
u5pBg3ByUKPcRkH47+dxv4mhXC10wEuQ7R6sSloVFQnNioZZsIL75lLuvJfgMnGj244CWrKcDLlg
vEm7MnBvP2Tp1mHmeHAyTkEMKAb8IU3Ho3xj3xk/yOQYu6vTT+YacYvSQTlVpmEQLAebI60i/gm0
EKI40UluEctcOJf2g9NexeBBCELtbCnvZw6crzpVX1jMPm0UyUAHABCiql/WbeZNzYcz7/U33NGL
ETE8yvX47f5aOLwNymi5mMQP6faJ7RJMUSlf5bVGCCwki4qw6ptOaDtgEc+Bx+I9Sk8IBNpiYmzW
QJtaJlHiVjukOs8zgqtjDoOIPNXGVHaU8/XcsM8a4LgzYhxr479oHRoiyGmzOcHDIxEcMIhxJ/fy
b2nM9WtGiHfzOvjhf9aSCUBmOkJpyJvAZJiuPIfVaGdAwFmnDQjuI8zlszrpVzC/ulPw84CosAhD
AVNaGrUe4+4WFvHpZ54ZyMAFbKxDP8XuWHADpbegm2azH56rMM91pajftqFf0o6zKITMfxO02YZP
Nk14lG/2YdA6ZcpxRbmwN5sO8z2xhRarX199sXoXq52XHPn4ikDsH0aYF7fhW0wskstXt1deHavx
Aa0mnOBnhn+RsQTnAb4OD7d2q1PbXS33Zc6XbbUwOMmCX22L22iF7CTI8sx6oAMfNFJVbySc6SDs
2B6gRvjNnWrUTJEEis5ooZsskbv/532NOG1szhJeUfKbHDl5BvQ2Jzly537bcUP7UrHoKwkMUoSN
eSwZD0sg3y5jI3Rz7pua9OmwqKMr1s551GIaazzr5US+X9rbIFrnizv17kUHkUfK4hAxjmIE5p5e
w/W9UFn90r3w3Fde+hFMo4EWCW4gEEefJU3Ew5ls4KJ7cFQEM1wwJj2S2zFoHcWVlhbRacj6H3Tt
jkmCnzYeZxpe+otP2A8YdWY+B1BxgkboOUUE7DSqp9kl6NDa7m/0LjbGsI1+bukcBa6HUWkD7rYU
Uusv2am0jQHQ5+vLcQC/WdpWXUa+ITDnoPvd1kcr58g/B6NBC8I4IQPH1Jjy2C4j5AdhIyoe10xa
VUWDyPwAFE6eNdkBKCbiXkOMJ3sSPwDPF4Vow5kkX4vmoAkHyenUS1enRrRmuuqUf93cwGwK2q+j
2X91bHUMsf5UuHzZ2QpM0RmOCAEKZsiEcwAGuJVmMeoIudiz4sBivJnGonQXwDeOGArGl9k6uTWX
zMqiCd4qzlsZ6XhTQS6wRlcEhHMm0zdWud1/M+cUMC5JCXQ+c1yjFO08/K6UJFx0vrQmboN+IHoR
pMZvSVjUOrmDpayQNjlKcitLTTUBjQIoOCSWBU1zwL4Jlg4Yopo05HH3bOjjzWSKN2yWURxFQjMU
4+Zmy82A9JjtZ9159GEzvpld4USoSE+EUDdVcdBQOJG43P55drUCYJpWFaprIWB1IgU7AznGohpC
VWq1+UvdQuWm2Bk8lVMqThxkeLqk4eq+fw2UT/5BEBGqo49fz9WzKTHoYuENdzO23AK6QJMGyaRd
YcJtnmuQaVxWulKZ0eScJZT964GdKctoYqBO19z1271UuxJbI+ppCOgm30BSJrxs8obfI/rLoT0l
bSgyolYfEwpoDxE81OW2MSYr/N6TBhu9Hfz6XDHN9dWjtkf3euuau3RLidDFAZgGkEkdivss9JRI
Abm/qYk6odzuCjZir1Jqp/ho65d9DX15HZw687n3x84Pt6hUx8HOPo2yyocxW8CSYqZOty33CaZL
yoxNosNSZIUPF7o5fAFwhUCeBRFHg/m1lGI4lresN0T7DLxHroXph5wFrbGs0gIbdbpl3eGTQ56G
/mnnLQW2wwVfiuA50490sBjBSay7iwfavNpxkwf3Yq815wFdwa6Fk6zbHb7wZBP9UmXbywtvSZN3
7lcvUERT16B7iwp5sgAqmGg3dnSiDzvmnpEjG3WnW2ihvCtcLN7TYgFjusZMEWkjHNzHNZqw0TTZ
dkRo3mTBZQMQjX/P1SnOwVboxUMRwUOHWMhnxiOEKiIvwi8b+hXJXH+YqwkIpod1MdcDl2HG6/2I
G8Akl/vBbMw0g/xsBFATF/YtUAKoR0tYffENSTg7poPYXHUwZL3FL6A9PZvPT+Alcqo/LyC+923s
TUWCeTRzByleeYHZZBWf7Mq3kuNSLQdUAnjXp/BLu4fqK6BAbuTXAmR+KIaBAkQ/6Y9hFHd8Aq0R
H/ZkCF7EsdMA1oP08ePydLv8xGfVuIMnNqAvHHxrNe3G77dZctQTIYqqe/fl7SOezQyupU811+o+
bqb7kccMXBjd5a14JaCrDgaMaPBluKrKtoT9skIF2IeYlw+sKhSFvP8karyDLBHRuAx2DODCoN3H
Fs0TgtTuJnvH9yqSM/L0taQ45Ra/0OWDQXJ1lfaWU/X70dWfH8tUNv4EeSLKjdOR0Qj9G9WiMwxK
neJA53Hhc9wcll1TWm+ST6rACaCge6OLE3iUVAaca2vG1ZXJotMaIAL0hk9TGZTmNuxkRZRyBWam
ducBHxyw6TmWOVg6leNIq/aWCe5VFXkBfUpfh0kjDIkGIfqTG2AjMuwU+QTtZ/Q0TSd3W+0t6fn6
DR0tU4OAV1GxaCvnCbIfEeMDoWuhDO+kvdm0R+SqIMDBil61BWC/sDFxgD/1JELyuJpXRiJpCBSW
59fwn0QJn8qe+7oYH3+nLroaoTcbkBxnmmwYzCN8g+DAx2bETk+tdeHeLbwdFtotkeCdVJpzNhfQ
aeA+6BfVIxbFYq/psJ/izgb86YBSp+7g1XYo328DKsoB8hTsYNpPnuPqvufZ6194ehRCHkw0QenF
8T8lMugb+0TUysKdkVPInDdm42BjGJAS2GtMK5RkaqTWvXU4Z9qZ62pAryN8MMhXCbVlCEqqGbLA
iiZ33femYOkLLX6QWabiQ612rfMuQNbWJTcTZWtkgIEVgyZy5/k7ivaM+YLsfEznQ3JMV1oN1iGn
rgMHde1PBZt3jEWIvT9f98iusuM8y17NGh73THfaIEj+TQVBteyM+c7QGWzXeRH/lH49vd4xRqQo
BoW5+PDlYlDiKi09WRmvdHTUTM111sVQr2bTvUs9xfd6mT6axkuUBaw0IqxDFamM7Fz+fNZUBv5T
qYIK6GXeu+hUfw8KhomDY7Tqm+yH/thv7POvxICBjSM0hGEz4SHOWEu+hRTysRq8ET4/GuyvZbHb
wT2SFHq8J5EsCsbE3jNfe8I91+OgIMNm3Ws57SCAvXixQV0d50+/Nnm3z5SFSgRJs6VFIWEsS0yz
o4qf38omw8R0Ch35ZjE6gDYxaSUm5b2AdItCGnTHXS10uDzNrOFod1b/q7S6J6OWbTUGKycQwHHO
D52Tra728gJ9j4H+Hci0N8bYirymmpuTfFy//G/bvDJw2mTLfGHXBS0HzOE9uvX337v/9YOiTj09
DaMqmevrHjjzFPlpBwFy6ybP0O3DkRvlzaV7HVP5HkPXPuX0MAL5FIE4YGRGt8/+m9d67LIIob7t
OAqoaaV6fPHRfKuHwFrpu4hIlgbbb/gwvrCcvxpM4vPQ4ZHCmRyok7Yw1GyACSbtZ9iKGu9CFPS5
MTcSFJUnN7iT7VaKskzHiDkp0whgW5uW7WJGCL+JIFD5cq/zfCYOI72tLy2nuxtA+3UqRwg37HXC
gxNwZC3h80npu/oFeZlhd+mGTwuW6jSKw3Z2gftUciEFm4AaaKA1Uq+OV4priX1VmXWww9o2mzka
yIXpSWpJeN8OCiQyRzAZeRxJz0XLvI/S2/wxznjZZOhq6pgluayJvTI/OZIjIBcy78Nq+CwggVkA
ZMaEHL0sgTlvJvEb2Gm/JH+udZKWf7NtHLWJ+NQ3FncBswmLHBNHiCUe+aNsUBLo+GNLzeD1JOpQ
7Ocw2okKhFTIE6ZvSndayQgA7c+4NyisPbaoKpC3qrXRS1lEXGQrjSWq5f6on1o/DCCXQYz+Fgf2
HbUuo1wrHk3GBlmeWLe2imgV9l9NBWfKS3g/rbMrieY1LH+SUMQGvFgHVaOnfHYo6BqZx7I53Lrj
E4dNwExKxL2yQQr1j5AQy18WRyIVvvGxpdlTznmdK1wC4N4V9Bk+IvUWzf1nvIQ1YqYyCVdXbIab
63SVHmyPc0ABZygsxQj8AjeEmBBBezmDa2AonjVgteVLOAoMJUpk0gVBN708/EDH4ruem9p6ptZL
xcWsvOxksiy1DJQLaMnVzfzDQBBzW8BPH5RXr0kYzLxB0Xs1YiOQxMwa0SsrapjoqWv1/pgO411H
LTQlM2O85gL2A6XvGHbLEwD1o7IHUQykl124d1GGAIafWFe5EE48kt0TeN5ndCIsJaNaVqBfyoXH
G+RTGI6MBYwPBhA5tw8Qsi6Fv5zVXjkJ06YdBOop+9KV6DFkpW8IRYr1UWsToEw14dQ0wkktUbXt
QMI+fxwr/joxktm8xrwJhPM3oXhMwPFQqxHl/3XAQ4+gHixf4VpsQZZ7KHS2QEilJyJiV5eXiu4S
uIPKiujmqe+MjEdxtjGqss21MvasXHLuP0iq8RIkvWuxE72nwdsma7v7b0c4rhaXn5xnCKM53P29
Ib+SN48jHGSe5Tt74sCrF5tawHQMLQYvlSGB28VI9U9UuBuqyV8bhlz/rHmRE9bZFVnKlqBs90cO
7d7q9qcxi8S7QtznM84BjKI2iZ0Yn85y+o6vZpXZFOoVSunVbuLSYg/VyG7EsshNEg4CABJOJHvA
K+j1t+ZX6dO3VjLo4IVs+sZeKvIWw136PFXQbzzeEd00q2trn83IgE0XBvUlEm/hJ205jfMDV49s
q26/yYdiFfHUAC0OiEymgrMt9CGOBTFfr1MiiKro1ON14q239hEvz8K+8VNU078vSdrBIoawl2ce
drR/6rTUKpnnw3MpWDLSG89b8xU+l+Q4J+aiqvt2Fho7GnAr1w6O3mK/UkaE0mUJ4xFUxZPpa5gk
/SGCe5al7lg/TGYeFANazSt3uz2haC7rEhlN77VVVNLS0HHJr3M8D00L4kg1hbox2ykou3SmoKoC
da2Wi5iXI0xjp58EaKhabOvKJAfXdP+2qckO/NHfVDLeq5yjf5NmPEqYWaL/ezfnsrmutoM4EHKl
o8X6yUDwbzRgFvYWBkFx+g31frGd5etyO1uTyY22NavnL5w6zGTQFY9zQV8l5cvgl4LoQPK2vG7k
4Ol7WybO0g11bx2MSiKbzg/z154Xf6jJEG4m94RaI6S97PwE8eYg35T2v9bjxhZQJQ9V6LMcUJbT
6kiIBDwo5JgkW1Ax5s7fwpaPA8pvRkCV8c7EXTGSfwMQvlgmwzDoVxI1kqY7WKuObelR/A+warE5
G88a7Tp2rTk2uErHPow8wx/e5Jiv9ERNCS7XhRL5MztzQt5R5KcXf1wa14D6OH9eCAvG1l+p9H5O
jkhDhYgN/7cfr8l5iK8RJvL7hJ2Pgutr6CEKjICGp1NpjvfbWBykDZ7B0IHZwrIRVolb9NcyLejc
0BeaFcvA6HiCmrX5DRJzuYgEDLQkxYsU+FVCxMDAtUPURZeUAskqhq9vLwet2hvrLAHsQApXY15Y
ILDKzhzxhK3U9YSLDQ9NFsI0s6XegPeZnsgKFRZeWlN4ZuZ6t1A23eCksJtBSgeTLrsLfgA5f27N
1VSQzf9D2E2A3DHdEsXmekj1lmMMtK5+jMAk/Da8u8HQptgjfJmzgcc6nDvR9w4/+Z7p04op18a8
dPr1wgn5dLO/1vlCvTxV4kyYwho18blAZZvCW32e9lcTUO5w4mUhjYnpAfIP7+KDfFRi69adzYNf
3HxlrX1avbNHnXSF4ZUPIl4QmGy+z3k77ED2a8QHMt/y9OX0mZ510cBYI6IbDHECLt0nTQ9Z+mYD
O7iHfZH98ZkZonqTx+bhMhiS5rHlCHC66DAdIT4itgKLMZEnk/JJ6OHCYNuluwdtElikMqIEXMLm
pC+l3HfBb67F1IZT7YTDaxbIw3ato4mxA7HkyDpQ8KsvFX/iXBnwjpOVLzqDgylV8m86gZUE+NZv
kbUcIJHkBfzYGgUTYKidqjQ1xjbD2gu/K3LqUWVqIgApTROXy8avh322kQRn8qXktdFYWPbalmle
kiHJ09OghUVV9pzUYCLDXFsHoaN0GPqqwR3mB+Dbt8SZ6Es5SfU/YI+j4xtBFZ5K2D+vSPc2nDJ3
N/Aj1tZQqZcnyT/xTwlUzSOzJyTJv0j01O999ILDMNhJvfpVehn7t+cQcp76wg/9u7w/nxzu4mFX
7edDvfZepgzDi6JcCSsCxtxgsCGKhhJi4UV6Brlce4z8p3DJ80RKn+vTFD2sT2wdEZE6/3p9Q3/K
1DssABvlUGKEhb/GFz0RTDbU3TcRv5ZjuS5X/WMbJ//gV2BjYfCtma13JcJzNR7TDNFtH+T/xW+9
kq1LcYnbtwyfLTVnIHMtmEr2YFFsLoK6kTDY/CohcFYSxRt+BBTBIVmby+DK6GdawpT48QeBHw39
4fUE8fjBm9YjeeZXKubwI64yAPFL9lGQ82OIjzKnm8bacdbPv0Qr68RTv2tw/CN2xrY0ecvJCpoi
6tY1g6+1t4lT6A1rF5Mm6lfVw7jkk5zV6h8SfIWo0ZBcpV6Ndqoj4Tt9F12nqWQA0x8xjcfoyyUG
APzolwGh7+lCaDfHtmzWM5FPpgWGmmS0tIzo2L5FEj8xhWYD2SOEblBrmr/bZH6g57BqykBQ0I9q
+FMMltMO6rRQ17iBUG6IfdUjgyLB9PPvY3ylv7U6MI6JV5T9R0vF+ukBsIUwKTgcMV45jTMPdGLl
Q9wvlGfOHHRJWl69MvyTz1kmSXAxz5M67bnD/bD9VtgHfigK8CG3tE21iOs1QGefjBbFgEsPrWem
/Z4JSxi9xD/G5Spjws3Tf3vm6No30ISX2cuq4qAYoBc1e3ksTFWeJq6WfA1DcM7LEJgd7aiNa24a
S8X9AZF7JW1OXowBpBXnS8l2zBwAKmSDfQmOKhN3IK+VJpOo75tVRJluabWJ4L+1xdlBG1KJ0O29
MLY9Mwtfq3VVeRfpI4gckH+h5H3Ckvl7BC8PLUkbNSJB7zxsZNcAUzPXpv9QMtCNPVspeAvpVq7V
QkbqjVPYcmMJduXJWu+EbFv9+w3dZCcpVeQVzRqVvgDj6zPJyGDdg23kwUZR2keyq01zPZRvTX6B
YKSk8TFXahqKRdvRlFTv+8zkmF4CEVeL7xgvOetv847+40wet4ZwA2sbWOVdJrLzKVOSLnjkbMNs
wQ4suJw5+ddvXP66MotwRfc9aJWkqm37aQL2Z0hr01YUqIheO5Ytg13HeLPkLiY2DNNPIAvwRbkA
DI/T5qOSLwqWUZ7RKbGmqwddNpFchbkVNH0pAyUyItdZaSgMp3jCNx3P0pDg0/eXvEEtnpRxlMwu
ZFMgPOnq4tCghSTCXmHFPDLSJVH2daUR5dQtJbPJye8DszcvUFoW+4tJFjDUYKqsbCum9KrpuKDk
rsZKznmoINhe8megfYXsN1TnramBcOS4xzBKh+GvB6kyjH4VDJgO69ot4SC3LQK8bVXhF5dJjRwz
6931nH2ODkQivmtDCXRq2i8S+7CdlV/HxlaB22SDuMKAd60A/rvUsFk8nZng0z+dATp9jrdaFKYN
k16dcal2YD1ADxy4APQSt9539CQNoTjwofNuAwhqKLjltxSCYCZapd6xVWn7vy4JkKtLbZ60GUn+
YFpWjEe2pLyAQRMksE+SDzcp4lPIKcrnU6HQdUAB3f7wvfJGQO0qpDY5YcpmKpaXJfNrsNoD+Q7l
4Dq5zn1ua66NwdGLEs9LZv92Y5+0/Erdlpjd7iSLNtSq7dEELF5v3P+8975u7Ka0zQauij3QJkW/
uqzk8JCAI4GSRaEXKPNmWanMdJQ0JsMkswI33dWQtYheS2r8st3C4ft/srKDhj7O0t6DRv2SYVoU
ssc6pFwmKrcZ5Lv1WgpzsbwKzzf2sOaQ4iU/Wp5EJZlZ290OqUnczjfupXAso0G/dsSKS6GD71LP
VeGGQSF5zcaa1kiLmUs13DkqVOdoIVMHLJFaO13/GRMkG3TWGsZA1o7+W4V58fyWdGNFCRwXvrz4
e96g2u5RuJTmn9ozn31vqe7t7EI2mlWzLGiUyGJFb3l3v1C5tHD+RsRSE1zXmSxI2j54a3O2j6si
usn07UfaRSGzKl4oaGAHT7oimwqo99JRCy6HIRkRS40KExo69vbQVSj+NKkxGlFToNvzau/t6etJ
m40lWExyZNlgzS0vu7TMFcGc1GmeYc4kfmXuuvLXImHiQB/uSA+abywt3YuzL7wldqUj1u82bV8I
F4JkNkvv5nY6GdgnKUfO77hS3Y0Cn7OMhzAUHzRACw7UBeZIjHpWvVCgwhfH3orcTxee9w2UPehh
jbDgd/iDtEl8EpPd/dd7vY0hSFEoN+tVeXx5TU56e/8uZSl8gPng/i51c6nUsAvqhnzKLvdm5+9L
Z4yB1jARrm0oL2mmWbiqhz9vf29x/X9hE6XiaNwU43nmvPMypOCqgqC3w/PMAfOPPySXUIh30iZz
FD+fndbUXgcgwnJU5EfhhMg+2ZUGxiSN2O0ulRCu/7hyFkdVU5tbR0POsANEe/pS9dA6RX6Lf7Ya
6gS6vj1sU3gn2g7JQxQfSvB1xQYtc6IBm8EAnQrMKJry9Xt97fmD0yF4rQvPANhRvU7HheM/JccO
U6mgJMLVcKM9ZGQeJGPUus9D9wLRjJvWNr4rQPOhtiqNWWKSz4ZDIba8KdCsGqV2WPuLyuDffg+f
4jJoNdGhQhtLqAiDeDzYHpr4GOb6KKoCs5wxrRCv6aQ1qw5OVxMBDFIeL8oAtLThloWU1PX7hBfh
UyNiFQwDkueT/rDYchDP+NkS2JwFqCEYyT//Hej9xC/+s+PtGX96BmU534P7ug6xJBsgl4GCU0qP
0rLPzRz4nD3NwzI9JpZHPiRiGFGSzq0aws1EmdUSZAOHHYQI878PyfvPvLfptuO+AH8aQYeUNSXL
ff/3fDinGrNSie8chPA6Jw335y+fLkX8VzF1qCRbk+emkVrf2w2rFnLg2MS+oZWgAHrUUiR5sdZE
N3qpxXRywPJ9fdIpW+2SvmK6KyafsX38smC3kzAXNpYHS8+IjXKwIdSWyBXFYu0nrdHSjDBygUUz
szsE+4VbVYCNtLFiD3UD8EuH1mmvsnQliykZKr9h+lqFc5tNJ+/q6Ka9JA1A4+/8yiloafjDRS48
zMP63IZ2erzY6ElhMI6gHIYZ2yFwR7EOe+LflhTZ6PKyXwFx5xuSjQgYdIRBZdPe0yQ+4o1ZNjgu
RLO2eL+CwU3GLA/TCIlOUoU6x4XOVbkiLvix4vBdFS5D9ZP0u/VkFp2Tb2WN2xqovO6XuxcOEEVC
n6uX9cQQUpEZYhySARYNpU81HlpxlJMdI4NKy9SigvbwvhCJa7QPm4a5zKxgwCFsHzfUi2B7A8BS
wOw4n28oPBa3ilj+Vjt9KwoNBEyd890pRD1NmurKwtVrqmF/LnihHUdk06mDmcLwko5hA5fD+9zX
WIRooa9Rs1jQibECAoRqbMc44iDlE5wRCg/VJ/haeGUuUwA+rthrILnFNO+UNcftD1ut3eLCdr+F
FBwKhLm+aQ2ktfHW9BBbOqbgQDVdXz/+AIwCBr1kBlb8LPH3MTCHwC0zpNI549XyzIabgfwFblTq
FkQOWIqSioVlUy8NDbtb6u2coOuGO0vhyOu0HcJV5HWC3W2NEBVR3vUHEDcwxloxjDPrJ1mSm5/5
T/yby3sO3nzYXkMjGTudE9C5CT1jNGA85B9XEUrfI67p2Nr2cYZtOCuvpOkCHqoWGLURMi3jvhGZ
UXl8Cm3W8G5slmzQg8C0wkn8e61uBL8LiBdEHpJ0NRhK4+MSy3Eo1Hwy7lsbHzX+gimdUZj53i73
rCiwJwjNguInLCICFwJhTB8d4ozz1kofy+DnaIDz91dbh7eDzAOOXCkpvCc93WRhLJvQ/Pc/L922
bnLF35ZZ6qkQLrDJsKil43IBlEmG/H0OLYlES8MKRaAxOkgZmhyE5fQb8T+hQqWZl/VxsW9Vj1RL
K+fJ0GVxDI+Y0VkeYLdx3Z3ipSV0SeXl9HQsiQGx3sqSXtWonfF9Z6y+XWJ/dyvK9v7XbiaxsZwy
FwzpwX6obuGSC9iT0evL/kDNh61nwbwL0S0hjEVqfxuLaYkIPjpWEqauBBSgCGcp6sOUYudDXO6g
EiRvaIexqI3UvkeV3Tr9ChweTBbdJvvDFuCUoazbFUzr5odXiin6sZJlDGkzn5x9/NVVLeOxEMAJ
XLQaOhgPZKRDPinl8rMg3p80HQyqwsBE1/ry91JF3JQZJFqe4TZ/XzjEjx9dM9EhJ5mKv9DhCJDw
0DAM2fsx2XbNPODHqjtBQnlzGgsMeaprI6aWGGdwrSc+iFg6BWYZGJZiEoW2Qe7bN1+qnjym+NqJ
6HSBps+R8FOsMFbvhD4uR7aK9PXrFiDD4BuiUwMNYF9cc1+N4Qgilasr5iV3/hCXFs6lfnJkSvhL
wq0HsEoy1BKEJbSEvCRlZCiwmNMewUj2RFfxFITTtEq7o2D8T4BLy+svnvGlmLqEYpPTV0erAfua
eym4VbrqJea7BalkkrawWe3DBhgyG+AQC/gp4UOQ4dYnskqrEYzK7Y+YQEmXU97tf1yawlMYukND
jEW+xsJlfqkb3GX2QhISZYRM+NSg93M1CNLuduYMT8ORv81aYR5FzrU9uTTFixwv896HUI2ahbOt
8JlFyc54dGVBkbhWev0Q5qYpdG9NgBElrsTRXIUTSK7P4K0oZygvfHnOnkTmxJx+8tvkTe3yK7xh
CxzYeizZJoVQIDdDzLWIQwYgxGFHd50HW69tesiiSzjk6dpekHcKQOX9GsDTli9uddlK9i1Vy8xd
+y8tlQyDt0xvQuJ7omrMSkwlu8a5nX9xShafwndXo5aXeyVx2/6bVD/87OWW2o2MmbbvsHrp1Tme
pSVMYhZPiAI7IW1JzsGvuB5JC6wxLGiL7Cm2vMD0DbbU6fvFsCIV9YRAZrtUcHuDnI4LOxrlLI5R
eg4s+DpTBBZbIWH0heJtQOgwWol4YBLMrwtNOZOWJWHSvQSigGpVr6kht+zAKwXkpj3YhaTS9OJM
D9nfms4HEk2sSUaHE8fIO6ZzQn0N0fD+krRiFY+/noB3Y361f6Hys+MbdibB08BxambWsJFi536r
ew+0tASb9S2I+n7T8/Vpa3hnPfOlk8ESbmC2B/985JzMVMbTU83uNd6epBT6k2br3pw+nSRtm96+
GOa8MLsJn1PccwF/ZHv0qd8AK4vn0d+hQs+XgkAN9L3ncLNo5Wn7ZjX4JPdJ3tM0AIfOi8RRJN1m
9dfGKJ/wZFdeet8MtiULQpvwAvzlp/gJyGhb9na7pl5s7NtFrVyYCSM6uu0T34XmvnyOEU0C/kX0
t+WIRoCuRqUTcrfVzOM7Sc88WPUVAC8ajyfYZYs0VuLkTjg4ZL6XDDneq5Y4TfGAC6tWjqwQtyUv
gD/gxKFe4Mnhym42DccFGKwzNuugKq6SeGGBcVEWoE9JwyMTHdSHXnlu1JoH7dzLOsKeM/FIsnw5
uo96EvBcEUQB946pJVSKcMbhEBnSOhF9gmlkfbzfY7N8fYE4MnBE6enrn5qxbgqtUUihIV3epsDm
xjPb56WFCD3OTXMOM7zISf0iuvdKmG1LOS+J7XRDMgUTh4VIjXoad0daenLWNDyvWNxLsebSsFHh
v46p/tTWDG4DGkysmE5zdG8OhzhHlqs6a2bXiSAnYan6wUOsA6cPOTEuaMtatSbu0k4ZjrFdLhvo
WLaDEo3teNJO/QtJoBYMbK5kG33phtCQI+FoYOY+j//UhQv5tyehQXkw0G00ZVGBITRwn1GdWnUW
hh1Cigu+6PMwRqtwhOx9BO3XlUU8y5SIXQSPfRdJ1QAfhyLCxXfwScEVq07BBUr2u1W1umBM+cf9
+MuX+eJI1JBl4Qvda+t8U/E3dxRywUqoM+rv9caORJJ+BtfqedZUvMmHyyn2HIpXGUEDtQEgEbVy
3UaQaIzcPrYwgrPipTUrVz16xVKLH8a5dtqCJJFDs506MxaRoqXxtzjaPfIPPoNyFERSTjvDjCYi
Thihsncpr7OUvrqyZp0ZA6uQt7G88cS0Xz4hzu7bYfrR2e2qBKBsRWATqVonq7/Ejru25SkzvGz3
EGwQ8XWhnF8B5GZat1AIlqGDGzNBmsJCNk1bqswu1VaVGLT1duOrvVOAtIJNfUJ2iL0bZCB1eCBO
7qb1Aoh2ZivGm8IosCnlxKKEeZ/AItXPYT/STjSt4Lb4DYEnmeD258zEZkxOXmNfoiEHPVB92LvD
v7iT6XsLL/etcTnOVI2zDunct3lSPdK2Bg5Hzzydmx7IGl8pk/jBa+NHFsdFht8nBbo2A/UWcCYd
UXXRi/8VFlTGXDPXXd4/gms6K4oBauzhc8kgYCyCz98mVbnaS/9Eu5MKOBkSzlFk7CMTrn8GEZEa
RHStdAR9CXXKXRG4/6cCCpy3FW/NDIWvUGPyTYXRQQe3yT7iP/bZ4GxkfFOAJ6je93Hzf8XH1no8
q4TE1WXkWKSvu0P1X3CQ1IR6qJbXwxAX+nCzQEfQw7l7gpqa0BaVwJ3NqG201qaFdYNAbyR1Z8tT
9Z5DiHHjrYdUCppv++0YO11uGcssUnP+nxpV6MPYEpznKhxfYAsc+UwfC7jBeB8e2D88rOnEuiNM
a8jgTOJKCW6toJcnHZ7dGRKbwhWYf0R3TFMURYks9KQIOH8SnfT1GHhj2ZjmULOoVf9IpEeFr2yH
FleEPNveABtdcuVaSqsfxr21sMc2hu2JX0a8TIG5BG79QflfkKg2MIohT3gFlGwwdhujWzT9EN2g
5v1pLSpymotJpPZlsA2HIq5HirJKNXZFdlP1H+MTxY9RjxOnLa0MJQhrqe32OmqFHRBl50AtOnPt
MQiQtBT+btPkT/OknI/EH5/bgxyI/x/Y7pjdOh98Bp5GdesQ2+DyOZPFjszL5aZ2ZPlWlw7FH/7u
nMZRQknkgKoln2bemCn9Ot86CxMSmO0fmARkUganJ37kQ2sckbj0B8CalYlI6b40p5VLJ8KhG6AX
3lRIlP7UBxXsXwdzRgDcPb37rb5v2MFMqDCdNDW4ku1vgp+GWrbLyVqGs0by3GUbKKHEmg4d9wW5
gb3G6YvKg12y7w3jywsNJd/k7al5KPeE2mtLkIj2CuDI7+Vbpxv0+SA/WUH2Y8F4fN1aR+maxjaU
4POLvsUWtxRRi/L+p0ejl6BSR69Mdh4XgPU6EYK8Lr5eB1SMNBGg7w9ExLEYmt8UBxSCFqEdQJTs
zQ6mPfNj2NoS4jqNfHDTSatX5lzvtLYgkzdA4QUlFydTq9lCscK/8twmyLIAhj4KBMtc3VgxGofd
g27zyRCWEXiM/A1Hk6Fpbd3T62gREZr2nO1Fs7ZSEAhNbJlxTXbOy439Rg0GeG97/83wxD3fkJnR
vrJl0EVhkAJBSPLeVCrROx2UysJxkFu1vJO/0oxvyWct9c6qStIrMCQKGzKnvV4ZiIS5GAZKSV9U
HII3dU9ZYoqCKMVYUnVm+bDFkju8blCwZRrHZicR/jBRAPMr8Z4S9CdMBn3R2S861ZumVHoS9qAL
2G1J0pzSAvubiY4WfvaR90Oam9rsam4olm+qIiBddwGCsJoDPvqTOIo8t3zKKLSrxs1UBiySjs+c
lf40Wt0eYZY7lks+axPOQfSH8Xe2vpe296nipJKv82P9KpOKpanc0ST55fbJfqIfVWqu4Z11pzna
Z9LgKuZczPBj+OKCnaOkVfqrdVHTVFZ/GE3kr3YA3L8626Q9C1fjP34Mov+KGDQORMBcYRCmXtK/
hsUzxTPTz5UB6Xhp8EQHCOcuJrLghZMkDskG0RebdkBqM1OIZypxuxQ5G5sacOZds6r0CkU3sg6L
9TmZ5oymYNLRiJkQqVJhwGZQj6q3X8j1AsrATkcrB9HdgNNutkjq+cB5h1vPITsyhH9W+irBvlTQ
bjU9vowCcz3eEcU0orUONX/KeYcbQBoYwiK3T/a5aQxCPOqflxVpikfA3K05OQ3Sj45usp9E9SIc
HcGeB5IhbH0z4v/UDHqvzm7CYOQNlxuVoD0ngTZ0ER+njiosmruIl/3VoxJYzIWa730e5OTwTjeR
/BzGRfoGPkFdAVg6jVVJpJvkLCRNfTGJrsomN2rcMCVqdEWw3YHEHgp3DIu5erVjMxdBnwzS4wUm
huXvC/fIUZr4L3Kq3dybaq9w7abzWcslgBP2tHnPENkY63X6dzRo7GXdwCm4wVmjub3XGo0MXusN
niKz65sORvcRYmlZ7HZO5ffRgApZwGw0B8wWzkd55qZ0qcXCsYDaSVyT+RCbPCKVKAqyVeA9s3on
3W0l0xFhufTQ2VCeI9v9paIPkc2ykte2JqJaq8A6Ez6oRqTwshH2BivKW3f1+H9rmjn4X498sAHT
XKl4vC8zs2/KkQ3ENbDb3z9NsBsIhUpT6cGWyvcxOlPdYcJu/cYTLU5RdH1iFeMT84tdrubR24H8
TyTaXfYjqbJtYNRjAkkUCNWD7BozMimSPls52ynnzoprsCVBjjG6vsYdyf5ZsojhNygAkfdpS2Hg
NgDrZLA41cOjaFtvx8DI87iUyW/VmqseV7Am1lAYqoaGQK4T5YUbKr3zu3s9j4MQO1lTUnn0TLLr
ZWRbCvX7Xqt/8RQ5GHC03iTUxWYb3D9DTCgwsci3Yz7JqLcQN+u1eJyySD0KEB+3Sq20Muyy6U4X
5Xvkqys5MD7/3JaW6TGXFEUXSGQp7JK6ppHBb84sTZEUESXxDsr23MX0wVJRWR871IZocIbGBEK2
Nh4YGcziriZRupgmC6585B4/ToEKTqBm7Qw6GYsGtzxsHYHcNgwqv0u8X9tgbCbpUNZ1m1IsepKS
ZwFj96nhZpRg6lzu7hPPwBxOT4+7lHfnjijKrfJjAyMXYpDiWsq/bQMEo3q68znSITlF4pEHeLU3
BiTADFK1a5I/RKi2relIVxIgDiQfMn1hQ52yhVXPSzfgIpI2aVJ+k6OeKIe/lxi0zmS4vr6OwaR+
AQLKjEjSZLfj5ha/uMz318WOheZUiINBQoIsewaQWlS4n3D0RevM8oLMaBRwtNrM7n5w7as+q5dX
vQf2HQCBJ+evKBm1ryUdk7F/etPXyzND/bhaoCViyU/kAYtI9TeouR08LsVb3gA+rvQ/1nZp0z7J
OnUhpRaMiqjZlGtdyqa6tlp9GMJ1dFYC3tpi6vC/nwO1izqj2/Ekd8Cbiy4oSFuFr+XrcoDH1PlU
7jkTSaE4c4p9qrQ+MMWS28YKMX1KqG4Jmt+ZZ1MnOcP3U/8hbl9DJyB3p/oGgKhXirzj+ZC9tCrd
yg++VMDSU02Suem5IqZIisQXTSaiybFQGNY5MFRx1OiKAYST5E5nCVrcMWpsFzGY3WToNqqP8vvJ
gxuUZ7lYjvgAa4CV/jaseyU7z8wE80c74Ik6Cz7D0qYMe4aVR720nrEPjPL1DZaQ6Mn0Rg3J2/Od
8zBQXRhvf1g0MIMn55QswVRqvOPrZ4EAeLJKE8cepHaAnLow1AwTfOGqK8zJmtQnc9x9+Ow0oEhN
7mBunki8Dx44ugK5x53GkVxXj4uJYG17ciPe5B1NOmQ9fy+tWwNyjbaGOTSZvcj38rFPdLDLeGUj
NImHMDf4+yiBMe9iEu5qYYixfNrYvlNVRJg6j2iQc4RyLcEdmGGxXMubqfCXQzWzzOgh/6EZC78Z
vo0gL3WIVivNl33YXyqekmiarIhuEq5MZSG+dIMJVwsEE4JO4Z2MbXsn6kU4qgK+7eARJU6hSgJp
W2EkfJUOLJ0CDnvZGd2JDgaA9vVI3hiVwinJcWz6d1TBxkrVG1/E/WWNu5nKbYA4a3nU6xEZhBzK
gi6UnUpyRXdzAH5pW0qK0pqrAJpd3cxSS7pBPau1+zm9fqJf02Eexf9sjfLOV4L4kPAz4u5nAwKh
zSPfrtD0J+7tUoAEQkP9rcQdKUCDTXLy7eG9nF2g9kLPUi7W2o9pKscsikSznCUxdxGTSKsRUQG8
C39RwXO7keQw63IkjTSFLlbh7oE8/a0yuKmENGx/upT+GVIMbQz9M3BWG/5TLbeTrcMerXsWmiEe
2H5jHjFYJrSXIfuxyhm1Tlx11I8lS2fm2aFEA810l0Z3OzpDRwDvSNn7CCet5T/ntJ5cw97sd2/0
pitPBHOU1d8M84ehN6salR2CjklYs5Vh9YVrjLGH+r/CtEQQZKP4aMj1PIij2Cz/jnksRPQTdizk
cQAQ+9qdWDT5YYd10nZqBU7SHCzopShGqZ3Yz0MSGqLPHpbDwZGRbtGeWtZSLZZ25IIi8yAmzXQH
GwY86zvHX3Z8UKV7w43/iqxWJhXK/WBA59lgHY92kqGwJNi0uggJA252YM5XpUMpWP2eRewA9ZuK
5bXiRyDj36DOXRFPf+n95zHCQWaT9gwaeZKCRLDPsD01eC4TC3PDlY9qPVCBsL9cawu557HX0lCr
weRywuQn3mjIdB++QMQ+sW6UaRYz8+dzwDJUVzEqNsmb+O9HFm3hvbR/lXrueLwLNkov5hZai4vz
8SW2oBQdatBh/80EGEqmjgIEEXNrSzRgBY/C89jUU/tufBI+KQiQ1p40GoafYR6FEZV8/xF49xr3
MZrx5A/zPeGEMErXH7PBN54yikU7bVzihF5TWmCvD8pc5s56lMX3SEsNmmNxFQ5g6gUvfZALJ89x
CxWYf5XgKnCd+/U35S/cBQ3uPZ2vcdS0xfyl2kk9IEre/tdkg6MQ6pyOaUtpbh5LkCssWL7LzbKY
WtelKR/lKzEhWhx+undulI3t5nx+LnAUMn2aXLpUwK7xxWN8FpExCxbo7ZJR/N9aOQtT7dTRtxZn
OinKsU7s9PWx7+wMRpsV96/0IqVZsuq+1khohFZC/bSsSr+AmH1jxBI9mC4StS+ljYKEbGnTh3Ui
fIor8DP8YwrmC0B6nMoHmMRtAvYiLNoCMzq78iNkQpuJ7k/T0rjgDCG0PGxIPQJYqBbHLev1ess5
pX/Heh3NHlI8JfbOMv1cOgUY4EepLU4ZIFYFV3eDaHg3omleqRFdyV+5CB21BExwvuaPrduDca0T
Wwq3nLXS3Y6Xd7I8Mia50DPO9BcinNb1E5eoYm4LCxks14PizYp6Sxgo5qYfTd/gmEdDZLVWr0JI
EogZ64bHVieHYcHOCXULSW7PZzcwCsgWTA3Kkk1hAi16GqMMeeFLActvACUliVToKHezhusxWDan
gknH/XKSNNfT6yW44SXqy0j4yRvIwXfRHh/rBwi97+gkqTee/6FInEx5KsCbMaORuyuaIHy0nhYh
xBRsmHxgH3XzeSK8pLM8SeXiy4UwE17H6U5hQACC0V1+on6FDjRFyz+Ofj9+olzs0LMMCVT9kxp2
pp6kV83b9V2eTMrml33gSGlBzkvqOQNfOhfjaAtwCaR3b8yPbYPaAnuIWtEG8ZbbVQbRGiD1jLqP
wYFbjkD+K5WEFuLYFsGnlExlm9+K7zk8Ow/H9r8JOtFB6uZw5CJLbqdv7QW9SoasOaJ8nw00IvAF
cnTEhC1kuraynd7q6e5Jt1ieZWvXu4z/2JROEbcbd+3fqsr2fL2ftZwD4VL3yn68DIPs0AqPJ2v7
Hagrk/qFpSZatWB7W/cdcswUzhaxFjbNXYx6Phzn6sc5paLL3Xg+SY7Uz/HqhQ9/c9GpEFjRW4JA
Tt5akPZ+h9fdF24lt/m0zWGM57/NdvBsA176BpVj8o8g5Y5jYFzCq9uBs5wcMN1AmC0PYZrQz3Xd
+JT67zjl80PIJdpkOQJTrpQprWgjAFDN4MVNKnh8I//wwLN2T9i7Bcllc59sCnCQwNbvc263dQkF
mgyG8BWw5pbrPZ5K3P+HVTw6TDbych55/7KP/c1CXsiqv1gn0Z6VRsaOe0RJIxeUq6i+vXndFOni
TpyEScjCc+HTSxrximrmnFurIbt3nzsV5+EPHEdiMOJByTYOxXI3+P+hcsi1tCaSeA9tceCP1M+P
rNfFeQsL+0Cy1baEfGsAoDl1xrgtj/z0qGNtV61mZauh4fPySiOo7brrn6v0F5GpsBbBMUCw/BhC
wCiBJbirip++2RyNkqBe5DNOc0csYat7ln2NclJNwbcCtI6IYuiwCjZ+s2BnXLwbammtw7uy0YqI
xYJTkTnQtFDDxmYtEFk4X86Pq4IplqmxvIIDQyuYU4m2xmTHAJPnvsFMFlg/i6TnfB0NYOQaM5zP
+qajmm9UnRYK7efvIubn+7mkTDs8jbOAxOd+BnjGIKjYsazHCk3vXoggwy/xNlaV5oj+LRZRfAZb
/4WvPJf3dTzz5vf/kyKSC4LYeNiMpRCkGVYsIRLUk/HoBqWBmRF4f46y0c5hLqsh/HknrK56ieMU
CLZiVJrAeUOthcbJW9DegI7Oe8IsyblUx5rKvCKOX6rdvht+PDfj23efcHYEqX9UzCGoX9uvf1zR
bQ+08skm92TEgUy23zPcQc/Bhkluijml+oJtjyF/Bii9CgtsD8ZjIWfEiEpuwodxuAKjvQICdonM
rg+g6bo32+Z8HVsQWqxQl20bKfRJQagpbMIUiYoosGntCLgfXcieeVfV+FiEIblqCS+buyzNKAD6
YolaLmIkj6YQp7f3NCXwz8uml2pH2KXe7hQKlxmfnrOg0UyRyksyRnG5FvzmPTPQV7UCl9QOkPt+
rwuuFoDKviTctrECBoXleJhN8cBzngDDFdrwI2rzMa3apFU1cEulWyaJXoZWusF7lBSpX4CCu7mL
SogrXxNOYrMXKYlCu1131VjXZbW1rWWIcgl4ln6QtzKxaWntU2qhYKe0cVKX8AOOD1LvnjDFuppI
yS9E33cqXAuML7mZwKXo8w87RpYq6l1RpuRz1Z1vUOnK8bOqRpPdN+n010rZfVskIdfgV9l3vlk5
3qJYNAtXJUAf/eHIzzgerP2thdUtezf99sHNY+u55Td3WdE/QQdM3BuGAdaiuRFHyPEF9BpA/2Nu
yklheSUtu2/qMYg5Up7cbJrofU13yRpt37+qvH3xM4CmcSYGLvRpoX8h5GrOqt7sMAX/byGxkc1M
xkc4LB3q4Bt07QQERxPIsL3WWnDrJvwPBuDsvCA55QH9Lk12EyJkx8taQ3KNrMoS0JRJH9QwT5Uo
8yWGk1W0rcW3hT2sxBTTiKeqftuFAokVpsGI+fY0hECxrcgPqJ9HSnpwamz3MuSjFhC5YbXxNY5o
7IqICALCdhKWJgV60SU8XwaUV5uVA0yei/u2zSFx+rIqC5VjgIlY4ea9Fu71n0CupS4MS7uJSbnl
xQFcaHuO12vTmrfC2KCYa7kblPDAGGuYYIvbCHr4psExGoXlg0p3WE2fTgh81S+OBN6SCAKlj9hG
XWyoT+lUXVyZL3kqm+/ERdIjVSn1ornjzHAemxRWra0yEmTs7hEfF0pAOrbHRQ+41wDqlee0PgUq
nGVqVi0ZdEoW+0rwudlkrG3jgAnw5zxIHJnJk72GuFk8Gszttrqt3NFz41zz2s/7+l6nAvHrsohv
a9M1fZ2wK636ROWoowid8w2amORJ7YiVCSryAF3tvbVaDegaHKoPxjQztjO9Tw03RsdtQkOvGa7t
iLUqAkMkHrNtZaugAOiBRwi/qjKHtnUQZUTQuUj5VmpzpFW/gJVV5RRM7v72pz7Q7dLDAntfu3zq
JTsEj+HeFVPDlRntOmZ3Gn4LCjpvl2qv/IYy2Bedb+CFX7/MchFFsbmUeuwqSEfeIoU72Hj8yEXa
kzVBrG1AftNXDydx8PcCvUjjFOvQZAfzrXQJVZqBqPyzOYl5PFH9LxRlNGVCR6ehgmQOOk3RXlWO
xnDXFWpH1Vou8CQQMNV6tZTRuc6sdIzz99fl52nlnfcYSfOHUUS2Tf2p23w+a46I6BUpqIdHdH4H
PIbDPj4AvLBfkBpDL1JlVcMeG3pc/z/rJ1h/AUcyHRhfsT6exJkEwWv8HssPnJdtQd66RfrTKawB
pVSbMoeAzx3xFlkMqCrivu/+5RrG6k9Q/AjO2TdUA6ERnKZeunxZgmT0xyfmdQI8ZsEg0fJF1sU+
OYmJXiEiMvA4TjhPxoB7aw1ahphDddzqN1RmejIiLryXjGyRGmZDc8nc9Uw970Pv6AzpEAlpFMvj
5uOJr0qfT6hG3qjvJBEdJ8jSW5DB9Lmy35hVwyqYA1EM1SpBEduuDUV0Wa+FMgzfbBLOYC7hufpH
FaxVgt8qGLwO7stIf1ZVOm+LNsc/9rLiUQtLzE+7y1fpxjnfmAS8eXXvxFRj7g+CWin3I4bCnUf/
RRgQaF+wmuiO+BcICcuU2kGJUEwn1kpXgeIVlD1kXs8j2DDDAswUBRPB/67yBhL+1USxBsYjgNo8
0SioX6i5mqoCi3KbXCaCQ3rMm6/dMbnaKdhBK/kbIL/OfBJ1kKRUEptPUgujRWCHs0co3ha83JvS
mhiD/aKv35w0Wr9D6TVzfmU9anQTIGCDUcW4PEatxNTLu1UYndvGBVFkgzvBU/A0ro/hIrFa4Cug
xnxAebx7WogYXLt0TQtycpFTL6cohyvebgoQ9XlEDXOvKHF9VyqA79qrg9nRT0Nsl8R7VA8Jiqbe
PpwmuVnwFPkgE4tRviJ0gPFEi1UhqblwFsuDQGJa4rmoPfbXha3NHF9MpStfngmZ+81CZl+MkUg5
AfemLUoGIBCETMoHzO97zySq/9ZehgwJgVu3wFIcRLglS0RNbSPyeNoG61XwdivzApWxUsBJVLiC
gFSLnBh5t+9R5cFg4AKy7S/ceHDOvhIF4H33/Swzv185FI1RLOUiCAuFUY7I2Z/iP4G7NSNscW3E
fpcqc2xopm+2Hpo8uf6eV/Lxd0j+xjbNz87/sv/nHqIOxk0xZoIGLAHJfTHaXjUt+hQ8V7MjzHti
KCDB+/UDTks26Glrbdy9FrMrtrTuaER4qb1ZjG8bnOCFzy8OXI7beSqWf31lzXTttQ6yc74FzMpN
v/94xqzIaWKqStn92GN4aCJdoJfuCBIQji20X5cUJGfJyvVjYEmLq9o/NkK0Qmbuz3LkjN8fX4kE
VfuzDyQNfO2RXj5zCdMm6l760EIIp6pcIOBX3WKznm84cQrYG8bWKdmMyeGnznw2ZUhYnLFLF1qV
IyetmcInqLyL3F48FXD5/UVQBRFN68afNaGmejpVonpfSLbvCxyERQdWTNmSPOPE2HPoOZERub6r
9Todz2S/4ctU9R84+LqN3kTd8ANO3EVBt7W3MhLI7LJTxuiZPOgB9b/L1HUrQ7fPLVhHoNwsIrxq
FSlNzc9fxTuVymkDJarKVRj1NtgbV5nqkJscycUDSxc03aGoSx91DvwHnPN+FXq/bks7ShALLucn
UuAg/W3VvXeQhBxgggV+uM3+gkcn6lPE21D6nJ2Bfv3ofQ9tkS/Cv0UMBTNg8SFl8LFvATMAB3CM
tz1K7/wPbXr5CVUUYUZ6Cm/bTyC01uQ03/1nSR0IodM7vWuufQtoX4/4zY4HWsJJTxL9XaLM6gSq
VcLxl84XzKt+Ip2UVGoM48W4A40VaCxML3lQsMNU77oaWcXzs+0qg9GbU01sUiUqbCaNAmX01Qwn
Npul+oGZ2VFwzba61Ax32P0m92WfwOyiBhwap88AEyAMZdPEjED+xw8s2Ntu13xFHnh4MF2SiUPZ
yHAsRkTvpMmS0n+cqrW//rTQSHfbxsmVYX3hbh/61GzW5ffAQI8x7AbumcoBInGIBbJ+e8cd/VWw
b0eB6jMVUCzrNf2Qum9L5Q2XjxFNYTHN211eEPxjO1mX77K983Ho2+XzlobBaDuXNMWxvZuE0iIT
uejnX93dK5Y9V55PIPGLlaWcUODlOKJOB3LL/1SKB6yRbvFzBn/psy99wRZHBSE8db6RxGDP9bf8
ED88XjrpFbDPpFTIlDM57o4cNgpndDK7iRJdGS7ZQBEPqmVMAS7KzA+o+veqqbvKykuEj34aVM60
wHwpDFZSz8aU+3eLWfi4FLsK1AI6rPZAAqFHL79PH0LG1SBfwa4PBN6/F2l4PbUy9i4JG21MFSC3
H2VpiyLr42BWwj+nXFokBDF/Yhma6lVtZ6346qx3xCpO4akXHc+oRk2+Hi68sL7N3hye5dpAg+eq
FB6Wz7S3R8yA4prvq/ZvcwPbNc9a9ctxtcI3/gYWLpBcvLmR4CCPjoicQOZEIeF6kXIYlPrh8Tcz
SQ9KuJodR5LuET29XmbCDezUD4joF83TvvpVpSXGRuemrlPf/gwnlR6CUu4WysbBoMBEcMyXk/yP
CmtIDqKjdU+Sv5Nu9jLNbBsA9L/bM7G5Lnz7lpi1x1GNJIrnoRTNxWAk0PlH2yRkZ8+P5bvC01fM
gWvJW4QrQ54qEO8eljVZ0bpx3Hr3CPiwxRZCiXQo5NHPVpN1DGVacIKI5rjXmDiqT7LNCnPnshTV
Yc3U6SghqetTlEnIq2P7eusDqaZvofPmAXqIyYkOIk1wTgTk29cflH9p+bvzZNShuKlRKLopuGEG
z9/Mi+syr49GF6IZxnqb9iMFPN00IfZG63ct/oNeOEemJOgBwlpJ2cq1rRuHIhX8o/HqW8JJ8Zlu
1svrLVM6qbUkEnNs3rqXPxs93Cz2YfCp9+Lh8tPgWxGuWwt4COmEtjI5MUuJZTsY6YDf+RZtJh6+
Abtr/dW+W1/zhWA8Qnw9yZbE882cUaXWDo9Qh0Wp9etoeL+L04OX/wRdXGGnz7VN2bumw/C+5BvV
W0gbxLBhQnCHfCLJQjWD/zwIvx5GtOh9U1Fw6dSRBN9P7bnHI5WU7Vx+RZcgbtrOwm0iidzsWfer
vzE+aN7nCFnygNzijfBbmVzObnsYD3RHbd0N9mXXqq0baa2RSdqab1EAiwfOlFgkMshXZ3xDp0Z9
475HyWbIe/9nwLinvxaQzFPPxTF0hIIXozUploVcF1LWX7O5UbAtQlKer6VTV5YC72acckPMCuF6
9OelHlBxF/THF6uoJFC4gM4TZEaRHHLuhFCMcntInPVYf0fV5KY5Nq/mhOzwdWQ+vACcOZU644dE
fwFUID8KcOS0xxIUfLy9g6ABedPe80Oq2kutDLEXaVnJ5ZkbyFPLaAp/PQbPE5WouAJ/JvSU8/Ca
8zx8c5kjia7sLQei7GNcPuwT4LiCZ+xrjTc1o4PwDVIYdTOFCp+OMr9unq4rRAYv0MpZjnsqSJC9
i4JCtMsxtET/NW05Dv2mXIEmzZTurn7nTfJtGK8qxkn58nLz3WvgqOiKOuuZBoTA7dH9OS4/F1k6
UXpKFZ6Z/RR7mngiwwgIR6W0Qzb3F7BO5H98djbhz9j3OoQO9/exAz9/9BkV5h3o9TcGuSOjLf9w
ekQIlfDD/yQBz/4eD6hzyX1e18RfG8RQPOQl+5b3gbpFjO0aPDCPU2722PodeDtd0lK3z7dWh1O0
WffLVFErh3nPWEo1TgtFrxx37Krp+xjGF2S3x1iLZWGvwNlFUbi1aXCLRJuXRFnGymfNS65KX9no
tcaJ9jGCF85v1tp13AyGnbgCRKQ1n6zCFmbb9Da7NLxcrJa2iET6W1/YOarubYRZKw2zBLS934uy
2Zy3YJtNJBw03g85BKfqfPMRYwbsa1sDHU4v/aJuAjTQvEpfrJiAnoWhuYWoyA4GpR2ay/nzxcno
megmf1RuDbUskUe1+Um2UU6LtPHH2q/w0ThkIQxQbAhOuNq/gDqBXpitsjL+Kg6WsaDRTJdYJihx
pMMyQSBdTQljbXsZ6ltHA9Fl0RzOQLLT5XuMa29u9cOVefDjNryGqQ0+XXqb+IgBXNs5oHfUtT68
0yQ4eRIRvp5pkwDhpLUU+dx9cv4rK5TAvOk3RRK/pvo84a5UNNNsWV4M4e0IGyBoEPYXG43qIU3u
q4LglF43j3W6mYTdPFZZ5MC1FVwcHl6gt6wIo2qw/4El74pANtW9mHAkJcMgIJf3AyL4hXLZiDnU
t1fm1hiJsj4kmCaTsYiMBrXirvSdoqsPVE6dy5FJ6cQL38+ho3WvN3lI3urOFlme8hTf7jDzI8uN
6rWWq5q8OseobdGO6HGM2/E+1EprESuNyV5IWSDwcqvquxcTSJU7KPh5DEZNmG3TyaA7b4QW3UqF
g7Z9iwmcv4+ZC6yZcaur5h8s7RvaaLRZpZ9IUQnBtztKTRnQQ21p4cJKR3wmGmsDcjjMKmR/TpLG
Io1eXATqfZX7JxYrm5METuQybT4apXRCTD/J4ZO7hzjjnPmrSUw4Xk+jMvIRFAJXeEjhTlCZJ2/t
kZ7v8hhpNf7OWJPyRD6w31wNmczpdDMWcv6fO61Nto2wpxyV0ji+QEc1X0G0dfSw0nfb4ujzKrwT
f7oKIoy9XPDdlmuWY5RXxNWl7JbbULjRC5UVrwBlgDBjd6ffRnS8nmTF3SiXMWc3m/cbSsYOa7A1
Vm5Y1p6jPjaHTaLa6HbL3uSZmtYECteJh2AljJPUQPljM56XUHT2Qz6eJZ12x8c/yF9NSEyi99p9
90KRfrSH2X2/YY7SVMqizPZRh4BIm/iv0e5RUI13kUNqqWBL3bMZr1LtnioLNtdLY/hk7bKL+4e7
ieYU3Uj5FEV1Bet0+EbgkuFnOJqD15Aypsxp/JEVv4ZX1T8AdGhoVrd5WnvkNf3SBzuWUSRdJl53
C3v2JdlJX02BlNvraajHa+7a1nZBG93bqsBqHKEYQvQGQmoeto6szszZWZzQD/ia72QjaKBtsyzi
zU81SPl8rnvCHDBoOto5EXFrudrOO+h8VviU3IFgRnq0TSrZgVm3CkySgsYrMyBJQmHJdUvAWQke
LrWrIR1m7nMD1QEkNCXV4Ud/X4lEL58eu6rimTiE1RhBGUP0DZmoQRsGSRHrcj10Tqc0rCps4L4I
fubwYJWD4xI1TM1m0UI2DO2PYdDTdYFCHRAdgTJSbc4gTN7ww7D9hKTQggAnZoaXYXbvGgFJ88B1
EXNOGdGmzzoZbDiXaGEOx0f4F3v1+X9LbyCd2iKBGruB7aCJb+Fv9K1lXG9VjQtiysEfgSeLoHmu
vaWZS0KeyuG/h4uJxfoZwznVm1jN8MWeG0TLoGNjeE1B6kmZA54VDnpmvIBV/Evm6/zf5JlH4sEH
d4gAXEC+AC4kEbK42wffsTcf4522pXmWcl0Z/c+2oRSDBNLfo2EFYBVAXcKREIBkjAR1LmXG7Qv+
JsI7e6O1GsEaVk7dIaORKx/2IX5+sqg9b65bZMQH+dPWLj+OjhR7m1Kezjx7JDMwBc0bcW63VhXw
sMTdENLv80avb129tZsW5ZBTbsFAoFLJIhj3W2I+rnhm25ZG4a7ErZWDtzQCeeMH/eSgv4acO+Yp
8btZFYlJpkludEWXCRiZRlHlypv9g7/pIqt3osjw9liUOLv9poPvkTup5LTL2t5X32DYqhlPbjwv
N9FVL30r5b2jdoiVH3eZylpPTONhwQKJfGoiErOIYPqn+GpfaEoPdo8PRIZ8M06H46u8d4iuv+bU
LeECzmLPbI/EGQHUGAAmYyNnpENVJkc3cBUOViq06OGCQrgGXUDzZ85R5MC4PFnBXhtEFIDGa22T
Z1VgM2ul87hROgt0tR3NFzfk2G1pIcNOOuqhRfE2gTjgy4yUPvw19vT4aw8g+k+mB9lQUjfA49su
Kh8Gci1qyIyvEyocdJCqkC0MCt3Sx5rtuDK9rFzek3y1HGbAy00JbClWSJhhSQUVqj2TGSeiX9Zy
UlEUg4jPzMyPM6ypEBtnV44aQWxI4Om8KnWpGVEJ36RK7AI0hJ2tJZSMmrcW7AZ9576boEy0oSo1
U7vnkK5xGfWqU/UwpiRnMA5tbLLk1zRtZCpaLl7/Vzto7NRuddiHSpB7oYMB9r94BPpBGh/0PC1b
VwsiZCz41w9tGDvf4sGEEzM+99G3FtzcRkh26pUjr90c6qlOg0f/1Mo0s5heZYdIihXUl/5TBRzk
ulBjTtwgQovyXNu0kENZq2nrh450JZNGBqoyHYzQFZMur9DglEOm2crT0LKtDF9ZZbxcNpKtDrBA
PYqPzo/xYA/ZwDQPaZBqvgMqbP0VDbicRW6lyQTfhrmxQ8al23y8Efkk1mWY9OGtf3o+gxub1mFE
yASDL+mu5Cjsz0Y6T/bXcBlq0PURFvlvZtpSk/KXJRixCtTa6HmLZGYlU7TOywswsj5zTBeeKXS+
fHZmHW2kMr9oqV7vmpoTRUZlUJifJpZQyx/RT3m+F1QiovNmHnuLl6pTdOlWvFjxwnxJRm7afoAn
v7kxcKaE18Kz+KgLlZgD1S4g2h7j8GT1+401UmjLwFW2Gl/9cXqweY092blLFmnxFjvgSiRqJKM3
hglEUDBDuAUs/d0w1iUGHBVpt9c1SQruhuxewczoY78ft0S+KLhCvaRuyuIYusAifXv/MvhYkgrP
KU+fYxKy7XylRbaTVr8mrlQs666YjzdPXlGu16MidXuvS8/xzXMCVN/+wNVz/sAIyenQ4TfcsOOY
L6FkgZ0cIL3N8qfnmYtBxTVkdXK5Pfy6HU8wbxWlGFQyqTaMVDD3UtJxEp7hkC1nlCBlvaE5EXFb
gw3nXC+WG/T33a3AAoBal2YH5whyWicrbyOwLHpTETBHdjcEyRhneF0AJxjwTwNeYWNUbzOdWrmn
q1t68OeRJgzjwjGjYEAPzhPfsaIkrqfZlV5VamF3Fb22xyx4FDOuu58MDXIcX9xu0nOFKvKiktbZ
5TrKQVnznmhGqDJfo1RDSLYaAKROAbY6Sphuwsc+3sbHCc09txBv3pjFtd4e793yrIzuV+pg3WI5
wKexzuyAnXohzzTH0P1WTcDJH+fIMWawh9ZwFnSMDJCiqJfikwr3CZ3opri2BPzYCAvOINLYbkKD
4VGegMPzdWVfpuU5xgThQxYCDrXHJgDntCyLBby7b4PrqP0HILeMC0T2yNNzAMR+x2pWR6joViDT
bJ+F+dJM8xDHwsuyKR9CA5QowmSox5M/hlt0CKh7VMjbM0odFXRQ4+J+r6tjkO/ihzUXmySzqL9I
Cmy/QHv5Bi3wIiqbzXi70an4djEW8I1VWYOvbCf0fUV/rLVQ1o61K8oPn9VG5cLAvf4TW2yNGtQN
cuwq+egVT003KFIYKD0+IyCWxED/QZgyZyBHes/BkV9pF/rCfQ34b1B7eSIbQbBiUZnDLWdnrdFd
rDLjIZpYDQBaXotgt85NBDaIhF2wEl31+qYkjUbGhLrkaoFHNqRWv5K8sLKDcO6d/bzue4kp1Wcn
AQb0CU3xJxpPRXFvuJg2+R4CZO9e/+QYVFm9inewg58hwnqcvFsrcxi9ikDaO1lVey4kP2Ph8Px5
WhgwTyjC0k6sfGJD65b4uHf5BJO7h1K14HZt92yOBLc8RWdzu/of3Z7GiBxHou32PRImiF+muN5X
KQOEpOWrbUMA+8wC0EGiWlaXW//ulaH9u0tuM+K58lvbruITi7t0RTZjydN6POWyV7X7bFP2b7Ye
/1THH6tpiUFmeibECw8SNDYoTfvCyMe1i3Ft6tg80Qhv/zNx0rfBAsXRIycJqr6Xt6kvg3KCxlKn
Fa/yxnYyz4OLEyQj+EKpuc0WPbju8z3WHo28MhLJszjM4845Gec97b1Xsxty71cr34apYfQDu6BY
bJRF00lI5gf9FzK4IF6Tba55MLfublHHOlk6ETBIj47YlCooTCFIwItKq4sIPaYVcDU58VWG5nH6
IkJ57+h0mS8uwyCz23FumvCY04ussIUV17sdh35GoQp9Q+65m+eLKa249CZS+0fPPfKYQcKW8+G8
Smz1VwEYKu2QvgCg6qJxJvSgSjWlxnBXRcCqKt3a342qeK+GSF9a0tO+q8M/vQvb59dp7avEa0X+
sYdL8dSe29sQdmvDCuPF4kvg91I9vVUBvOQiWlCRzCJOvkZUOgq3s0XyvVpQ6u4ikGZR3lbHAYBB
bYKB47PlhSNi78XQQD5UcIKPtA2WrivczgTvFKW8jtNHm5WmfjIhQY6l74B9dPue51Yx9K1c5dHt
pqO9BCHVuwKObf9/fxIdiQtuuO2zoe7n34EBeRM9h+JNVbMFl6cw2j3AVmHDUWUNLwoGiW8uGju7
N38zqt6uNi4dZdsMe3gd3k5RQxH1BBQDyI2oDVctvA9BSf3gCDexhcziCj8UI5mZyZD+VG3vE4zB
f+mEQEFiQiqWofcn4BbQbtBwhEmgiuxRbzFHnsumedt1Liyb4Aq3smYMmnLbt3ofE+rY7+sYnO3f
I/decyiJeJ9aJ/BLMdG/1CEc6MzD6OMRou1g7Xuqa4TpiIkx1lJEhoII8JQWRmMavafs9d9wGpAT
tKyAK6yhuSAL6cijZRDmmcfiEUyVKFbiAZ/SzgT4DtsiEfPmuKzBT4fDmvwpwDELE21LfYWDZVJV
pf+kv3fOIO4JQBLP7xKXFzZ3AitKX39hrRb30daxYkBE4tybIQX0EovO34aaNoZCcOHbZ/wGjvoY
o2qcpfXCQL0EgZqYX8A5imXQfT5X/YKRs/aKh/xyErDsC9/pm0If3yEbB/PbswoNjQUU9hNPrlJ+
pMQTpYylwnE8LTI+5uzZ/NgUXbCpSIIqdr5IC4VkEubYM36AUGMrZTQujkS48UK81L4/abMU2gqa
5Sx0S27SBUPOvtevXnsEsNN85y8Wyv+K+XwiZpiiGff+AZtFxwbzj4SK7rX0QfMLsi23VwJ16ido
cpc7NV4WMZ/r/jibpbxjDoA/p8pycc1VSMoDjNQEXqPfjblNENHYqpOwrEGZvUFvDb1wj8Txkl87
RErMv4DEROH/flE05+GyaeHc1+US/KRKXWJ9gXMhHNTBXuyG1Ujzho1K4AiOJk66/xMvc84zH37g
5agZPgOnnR7Q1uvAhuxbTciaj3OsVn0Hfa0vz7swFDJ1FgLU3iylrxfggarCI/GyAHRYiYH0MrIH
0mFDPiMub01kOH0AR+M9r+8X5lucVzcyAJim+XaOeORrOUtxE7+vxAFBnjYD0VB/W2Cs+KFS33sP
mNHDNeyhCLkgNGn2Brw/H66GOeQXDCVDTwY93m4Kif7miTFmHCEZw8gArMIDyHpg2q1OPdEZTiBj
ZZkRPVVlP91saMsVzT7e5fwZBuV0V95JvaAKR9+8BezRBUducOxypDshRNBqMy7b6p/cns5FsvL5
oJYQSQMNiWOeei/J7RzHoVBSK2zIfHxZKnq5Wrl01G/uT23xvit+cPrH9aczKVzsL6j6ER+WmJDx
uLl4hRsuJ+SnRpVwJeoOiuBhHSSYLVmzWuGRNopWX78pAk6lJV1Y+8B1ij0aErtdwojqy8GwgE2a
YXszdQ1emuDSeuPKMZGApPEOOhZGGMMaO07SsLZptzUxmYZY6dq5emCKOlDdIiwplzaRF3NKoQGG
VN3VWg2hVLE16J7iAcTwBRzYRtnY4tFj7ISLqdk3K8TRQV18HKMOLF5Gy3ro/SP+tA8fGSzH8Zgz
KiHfFud+dibRq4WlO8cI9ah0D4mWMDLqyGdLGIdPNQOPyQYDy8LQrdvPuooNRx7kA+TIKvtDGMla
BjbS3bA0zpo+D/WD8rS4VKpU5eVC9GvWIGdhSJuy53DGfdSbW9p37gsJu/GXNl0g9AEnKKWTXp9O
9zeJNzkc6Xs2sv40HLRP+U5n23p71gps0I18nOg3H6CWrDKmwp27qnux/EWHS3+483lYcNKQuFEo
2BGbtBYZLEhNkbpDN4RbeaEoOhqziGRxCEKupxpBb+/KC1Y62c30vFdwzZC+uLUQBqF0xr47oWyb
n1G+ak2Aoqr+t1Q+uXuGE7zzHe/Rv22rfvVedum0lqIq3oMUt+w4SVnnWx41p0CgXhzpocq9sT3t
DacUVQSFoAmTq23mkW8nraUt7wIaQbW0yb+jdIAgVr5NqxinSlJhQNLyNDFou4ULWZTySgK2HZ7R
gvqZFrtdEh//ig/r6LgbybexDTH+6TtFIOAct+Cf3vMsxTOQ57724Pq+ZBFOTMmcsJ7jWDXiYFAe
sVFWruixcO1cJKz3iVGrjKLEMeo2jKMj1/+v2F76fSofe44ru8d8UGFS7ZnZNNieemfTOEeKZs/M
5tdWTI4QDBRhHFVvq9n0GKvd5BGGJtxrxAUqiNj9xP4lc69jWfXvnedNFIOXa0/3M6bxSyVDu+sP
aryza0bQj5ks8Dd4jdm6sZFSsF4U5ywJcomIhbWojMBwHBpCb1HCbUphmCOjykgYE31d8JRBvtpy
jJkIW2W9RINKQd9QBJiIPGHJBXAuY2cSzy95Tp4tggzoAnoKBKwQVq8+jRb9iJkzW41nvMBnqqpP
FD/Ir1DLoDZFZIlFI+ngFC2mFwd8F77jwWl6eUUu6PdRqXKc7dMM/17vW2Ib8LgPN1CJEU3GhHLK
V5eIFBB2fgDAO+VIeegyiMqyBNdEbITbqcnLxLAdNERuD7KC+L20+M1Uc1dr4bhdYef/ibMffngw
1C/iYOcx1M91mVBcENVhSMJ7Tlin8T9X67ksKQsfXr9hkAvKs6+VknnX4PiOxAIOFxmUlrQoy++i
CBJQr6iOgnsG05k9oUhqaAHGoQ75QvONKgtY2RzRP2qSswgnAE7VfTBz5CmTNDHifN65hxQiStCc
ReHKWFazE3ynyHeOk9P+kHPV85HaJ8gHZjZ31kOJYdxgTUV6iHG5ZQ0vydt8KgH9dBfm6KlQBKkJ
jg9Ghp7qrSHV0k5A/XJlU3gptpHsamdMwQmmjaLs3efjBTtfFKM6V6ajYVVasEtYFB3LBrs7s9Ej
mODYjJxPznqcS9fekj9F+O9tKPgL7OIO7jfwbqiDoWIzxUHqPtIjE9KdoDpf0sPaxuKzw9u5/rP7
KjXlwjvSqzH5JvJB0I/AnfWqJhG59jaY2ZHKyqsrK2VV3XMbd34cssF9iRACoyiUihm6wVJ5gqkM
/e0ZcwcxsL5mN2rvB3DnY6kb3xgZJvbg4vCcgbv3YrHaYzC6erZR1hQPqAiy41jMp7ZXPElnMe/a
wnKt7ihcgbvLNMvl1gmvOCGOiDfI8/WQes4c+JaZg3n5I4mob8Haeqe3NrzCEMcIHzJixlQeGoyt
A0JPKeUjQIPS6VM+AZ/Xh5C4KrapAIaEni2v4GmcQ/Iz+s1EeNT9IaZbxMo9t0IZtFW4JzsNYFUq
mGONb7jsRjxyOVP10AXJ1Vr50V9fc+j8OSSmNeDtvzUWdM45rNQuhn8yf5KqlIX6eglhWb/gM7lJ
htoD3TP5w8YAAP5sHWly/AHR1ibuFdDuRcLDbrUEQ3Qj+ITaBhONYeMzNP836AdtZcYTEvjqthzn
dGPiZ7egIGL3VwXxQEUBWHRC7zljF42Ti06VioRtysDaNKAW9DFdMT6LDr+c3dG/2ZP4A+vxlisO
Acz04PodBg4j1mxgcDcaa8fvoRb5BN/DTfJ33pjk9kRnYVeOniiZUe7fgKxeyFDY13Q5vfDARAJO
Sbs74g6ngSCTHfjByWAsAbJdyjYu4l9av1MfX3IzB/fyk/9HPh1K758rOhHhNUjXt5TXuOzSb5GG
bKRXaPBIXwTUpuz25Ei6MrXmoEMemdhXNWFKnw44SiN1Ps0+v+hG0dFyNIrBferZsVlIagkM+hXl
zj+xdBKGS3b5GuKGndg1nAfXIsfFlWIfadPBCnuLc07xf7GoGb0EjPVEBl8HDGcsk1aIVYDPj9Ih
FdQAO7I+1sFGE0nDQIKGeJ4r/6j7o2PHuTMMt/RZRGJWTUjW7KOoREDTvAo8QluSt4QwGlibzHr/
UzNK6c66K/VfcdD6ctCqs5J03tpCH3kvoGo/DMjogk80L5KqMrIyOva4RIiZOYf0NjsBccSpadXt
YDZL9k2+A/hM1aF/WpMiHAcAAAl7BYq8oVqtfGU9uSLnAXJmkQZCMZcg0G7V1beWsO2872bD6mb5
QaYwd3STJLI5/lDgnoHXXNBfoAvM2ahbQh8gfcldepHOc5Deif/xrQsZy+7hRMqqhOIyy812pzcW
QpX0dWpF2mqjJPb8rGS5cZLz6tCz63U0Gfn8N6h+RIMHMQ7kdw1e5EhjzpgHTtc9K+o3rgDeb6zb
fd+cUNRMRhWngbctGKllj+ekm6xXqYjuzV/u5BMcl8xNqX697IPhHnEIrPu8jGTg+T0FkCUVNxqb
U2denm4b+jus/X79ZQTS0U4ndltouG1+IWmAi8biv4UGzqa7UGnEf4rl+ioEjmrDPcrYn+9tI3AR
QlgAmH1wixrphjncWgIkqUo2qWLyCq0wPDttDbJgbenXV1uWi8zu0kUN6wjG4Oa74ch4iIxq4NYf
10Uogy34rAxFcMa/AnsIKP7sdI4gSLTqaridX2nZJ/ia9w1TeasUDtjxgBgWI3qZvCvmC/UOYaRr
AAwWWE8bIENlgLM6WNpe74LQq03RrOUezqS+JxmFSV9lqZLAAPmWTzpMVAc/i5eFHxExazt5jXlx
wW7mXeKT/y1gL15tQrrLTLvKrvTfj6KzrSFE29AUHxIRC/GjvZb/VKEpuVtENdErHn+GJcZwdZVX
QCI4wIAt9DnDHwnnBOUrzBj9+aUhOPz3Pr8MBdSFvmFd6+r93tKBzPgdehmHeNgbbsSQmykXOq+Y
ljp9LlfSgKfnAgKV4nNWIV5f5GGGVAssBcsnF46q9S4z5d1o1sAcZXuJBXUVXcW6UByoHYyw4Hej
aL6vUAjq2zRxyicZ6bd+XT1zzmiZWZ87XSAtS71fscrqXa5PQnjYpFW5JIQjrlcJZMpj++7SVJup
uQBDz/NYjg6eyZHIuf5NSdACcy3ETLjIkrZmdB3Nij67pNhmToHRpVcfDB8HxtQ8cIPRYoLlPG5A
nQfyTpJ0NuO0XzmG2q2UXdOeTdOSxFLZ5Arl4TKMwDU3LE2gPvWKAsBrRUaYh914RYwFbSbR6jFZ
jTXgDkPC2SlmY0MtU9Wb1uI1WpzOkzlIz23N0Th+OW8h/X5IqkqYLtVGzeqKpebF89Cohi7p3BbK
cJhkYeKQd7R+AO2GlSrVYsPuTBJBB0N0+g6/l8Yekq5sXsexpcATnuGbOpUHcrYLt646nIU2RJpy
Yv4KMBn6iB5lQ0vOY4tNEXfELOlZ7wGGi/ffVVVth5JhL0FTGgFDclqgH7aqCr7ajk4ZqG8q/cjQ
KlbDOHi0P2SJf4fb+i1y+VwMddpYJ8aEDRgdFcD7E/4OAqx5ccQ7GnYH4/u1RjL8p3tyHeiZDDpe
58FCGyo/TdkWKf4UoQZbRJRsvuA7rd9G74eXrAep9zbtb702cNrgsVJnzSVOA8sVrEYkpTmeK9ip
nhB1o4Ad2v3nJ9hFZmPjbooa7oCcJKsZqHYMjQvuyj0nPFdcAF1QY+f/AF4YrtL8e8pJb/vWq7Bs
/1VDNs3d4wyqJVsEdSKofAPoMfPpzeF9kRNrWcRNzAkUFsPcVikXvTm7HW8MNhvOYsrVgSiw7F6a
Kx8+MRyV90OuGkz+QCU+b2UoMo8ZSkbn7T8qz3hWBuRwx6FKuhZtFhZ1AS6+sc9DGqj5nFjsGbyM
GLX3CNBQzbV7b0eq5wK5hfynsb3izB2pqmF0sBqfRVC3faIob4pAQ1vFAgLh83mD+pGNU7HRIxGu
seB+jnGsBOuUSb8SmDOcIRM/ZOfq8+z7ivf3pfcY8NZU+vmL+TiXu4WAk2tWti8LHaVgEiyejcFd
dwtonuyBFK2EO7I16i+nghbqC/eHn2Vdfr3CPW84D9CKh9Sc3j6nMKzr9V8/ylRAycybwfn6eIpu
eNim0H8qSNV/c6G00bJbWp1SB/hT76xLUWY3oy4VPotZS0vMfJ/fRQ8JD5jmX2K+GqhvKnFx7oOR
ymXSGxyaIg9IqYUknf7+QTuvpVpoGosk4gnENNe3B7NjCmLCN6LutQqk3A8oAiKm6ehoF0Sd/xP3
RQxDmLEEZRfnjP7+uTXUCAY3MFkqKcLCB1kodV2pIVz7LNtebI5Y1LVHHjDLGm6T+1c1npSwD8ry
ZZs3i8+/DOeXrfmnoTPBQeqGAojquJ7CacZhH3HDbjRCtybsW8TY3ahlM1fFHsEjDfg9eozH1BGi
bFRoy78v5jTNMIFuho1gN4oBMzObnoCQYmC18XhmuXRbPHCWKd63jXjnv2f+OyXPXwi4vs9i7tdt
0QkIG6kTWhDzY48fHRKdyF+joBvJ66uB6i3/xi0Xrqg+oe+CGaV657IiElns/FAJKTtlveAIaHGm
7Asm5Pw5yv96YLMGjYYTUsMZVSYMVFuUPxun4mwvG3WcLbJqJzFCDU+zpKszDhJ1r/ZvpInoWkmG
LhuC/kl3b0u+j49lT4D8Z1eTYYcvj/MKF2uU5pxvBSpK+AaeOJbGXMsBkhQgcbo5ar2w4Sk751v7
xW2T3w1L51jXoubhF3zdd66R6lpmRaLJIi2AFK0aVDsIgdV8+yPeF9IEOaVPUd1+aoQ7Sm77jXjz
d1pjuYVHuo2vzjzihdrkwoAwpO3hCuulpcaN5gxNI2t6M+fuXd55UvfWacuvBMYsObTM69dq7ZzG
9xdJRJXKLvnvuEJ/SKIlXPoPyo2nksA8+2VwGgeafFddviMCB5s273dxeu8b8j3p1qwO9ocV6wqt
5+BXJ1TXgqseWwtjTJYGm4oPk+Afu8sFeIKB02eBlbVCxo+EvNlP07u+NGvA0nSnGOfhCDmiPrqo
X+N5ZVV++bSdCiWgfjtk6PzYB95lACFOcEQXpE0ikNMDePM7RqA+MNsy/Ns/IDMzpbxECvOyzTtl
AFPmTOnp/u29FYrB1lGWqcqMHjSa3MUq6vJW1Zd+hsm/9ScuwhOV+Tt6aBkh2ko6q74YN4PfOsJ5
3DDnP0qyyiJ9OPZRhGL9Hz3LnJj3qKkKq2QVRlWx8FPuoWvn06+QIFkjIYqPjrHLnHbE/yf4t9ed
eY8KNnzRePG0xBLPFZKUMu15/mSPjI/lnGOpc42SHYDsRE10+5s4dQds8SBfgvoUoDP8diQzCf4E
j6qnbBIbFcYUhsknbaBkSbpqamkx+M4MRmq70GNesT92t0JSg2ZY66zzMNLF3CN2eQmR0s6fgnX0
NSryGQt7c0UJpX16ypF1C+SZHbB/thFdcYjUXYRIIoKHVWOkl6Z700vjfv+BeTxdR/NIYoMOMhxq
GghQhBrNd+N9i3lVAlhW1gDzzTygEjdMw8IHO7hO9ExLNq0kVJnHhWpH3RV3+V1co1P74hZ+WWy/
rBIMW9gqDkG5QwCWzZgWH2APC4mifWSL5tDDkVVX+0q+J2xHueKc+g0SfCiccuOkajmSerKHJQdp
/fJmVXaDC83IytdlGX8Xj9tTPKv1nygVQQy0xO/P1OrPBdKkjGTfa1Sn1aOIrWhvMjaxKBWcyx45
NoOW81LMPdmWGr5fy82v2GENIZAYVMsE/DtR6Q9sLU/A7qLTrgC2WVS2IWqQ92Kt6krT2zAMdE6e
wFUaM5jdX5uojRM3+j5SMQoKxBac1sxNX3evhVTVxFosjjfM/Zzzla9D+ThAQ8wwol/09tpWZEWt
82mt2UqPsOVmrC8+nU33DLe3kkQL87x5W7F5AbRhZ6O6+pV6zveIjzwsIijni8diUbCDh/8rnapR
jI1A0k9DrCPTf2hqgd/JCaiHCAIoj4htKn+YiSAVCLckPdtPeRWzk/Gr2dlB5gIfDN43/nmNnMCx
ZJGF0r/n90T2ediZacsOPfzW6h6uJWKiv7558rSqk7G6WM1QEUCcgJF/U9J+6l4/+hSSNkyMYmCz
j1Edt6I5AAUzc3CIExgWe+rCUfFAyd3+BPf6eia46lKHWis33eiDGhrTmcUM6UOt68NwLhHH/ztL
1N+RxnWKzmcM49pYxLtDLIs3IoVJRlyFe2rWHmiKiCKR1az5uvXPCZmFv16ZRrmpFVZD451eTl8I
YZw/OuRbR198yYxyXu6pNrYvXThN8WqEfllYp3vYAtxi+Fn1Z9eb0ektsNzJYQeovpBMqEpHWBht
bWqGESzP+EtIgbnZEgnTBxLCGfc/ksoXwQ93Gc+0HzX94gFSnuj6UODwnIVNQtH6ga5/36AnboX+
GsPzJaykQlybM8zuG95JhWwBSYSoF1LfJ03FQHte2lvVQLuisfUMLupChu8tltsxwLOMMQMh1OVJ
8PgjG/PKqrVndBtprCjT4HCgtsK8Sn3ZGVOpMRJ2viWazad5408h2uzpUAyYguTse/Uy3ppS9h1a
M7wKsI/S7Zn8isqqqlT8t40kItuGcskmo/U2omy+JDa26kDY5ooJNmA8dZAOPSyUqEpDvObCHfPg
J1pN+F2DxLpcWdKiAsd+tOOS2Xnb6ELvZ0z5G6aZ7JtHFIyB0zNcUPc7hbd/+ruhXKmn8KMy1eOG
8WNW7hnicUGjTMrHWV49U2M6FLCL219KvmhjMf8iogay2RonfoVs1jnJNJH/hE41TDGCCZOG7sYS
WtNDKJp1NOv98l/Ufjfik14AmdMsY0a61zPnxEY3o5tWQ65zGG+QA/zvemnMEl1CPqmGWa+cDZC7
bDUnOdveFy9eovVAyhJ3Xgt68F9ahYNLEw6ChoJ4zn13hi+e9VhNQv2OZlBSplgPY83o3wlxBw41
3hKwPOGcbijDbSpXUCOVWeba+hpRcCSTov6iwK76k/mM51xCLRCEEVhBG10ofVqpC3n0lfCrgOaI
gwAFWFz+fFVDZBLka9rddTfo50/uqtJsVLzDpL0ojdH7zBsf2hOnOzNovI1ZqRAHI8XIL/+4fHv1
1shq6z6e/bgnUwd4HBSmNuPjhcueGj/dz1I6GEVfBXoFn3ORfspE44js38Kchg3OmYRUYck4sHFF
lkZ1mjm9K1nHu0IDT6vpDIoFr1gbHvd1WNZwvJn0AihH81Yjtf7RhFdCs88Rx7iL81/3sdhtUvmu
LoyUm6uGsY+bAyqKr1/darDw8w9B5KUAppoSuy2aiSSgMsyyq/r94tL/vPAi6gMk1yM+jnPRiTpz
ZkN2SIdXyrxrHaq36vLkfdZzJACH238othM0FVEX8MDGaSN3wSTwR7UqAyqP/v68D0Y3XWZwAYYw
tlpsBrJXvgsizhinYqx99jyp/yKA7MJmrBEKKCcpN/MOB37bujHXQkFyIaf+CuIRBK2jN6Xjh2S8
VrtzfMx39lUaNGp9jCeLJLm4wQWKSdbTe61UmL98g/dKxzLpfr8Nii9jyBdo3F4+vJdHdoR3VGGb
qBbtvMn2biKS+AN+nlCbo+RRdQZi2+3mGwVSC9e8zZD3R7Htzm/Ec+EqeRbOaw46hK8sTfU412mt
ErFe99s3VDH385T4y7ZdOl+t+USElyG0JdItmq2ABWxTHJbWTHrQQBLcLhSUAlmzbkw/q0+IRFG6
VpCmDDCGQrqpr/US1rYT9ByZ4Mef56dEeW6j+piEwmY+ien5XvuK7rPZg2dbfez4vIPE29qOKOBR
WSbhNa4bQKuAi8tm4AkNkahDYCt+SARZpgQnD950johPbY1GX7g4AszKmfskxZXK+r40HorBe0mi
ao/KWNdFtXnh0fRzzkN4K+wftwNVxBLxWAX+qN2HWeJ1/dW6UfTpLBF6757kifCB6oEOdfRQvAAw
jm0b//puKDzEbkicGLpj/nndvXg6aWPmhdjgf16QN3e/K4wFgSWxr1uX0cd3rIxyl3zB0I+At9OJ
JhP8J7qGyPZyxGVsXYSSjdg4JqXvUrbZd4MYvazOwKq7PTGRMl+GFJq+uJHtaALNAMf/KSlgnhwQ
Ba8H1KRcRrhLuoERbq5ey938BiKvek9wa3t+iRNOuF9pZxzYRBqq2XC5V/NxYUYmIIUwoED2piSG
vGmHq/693nP3Q2f50FbGyvWEctp4hsGvYjqPnzUnIniTjcQ/IiJbP5DaCIR8ZhfKYRjte9RSdg7R
WYBcx99/mUjuhlf5+ESRZnHiSvPTSB5rSwwo+8apbCg0n8w3RWcKCBZZAy9RcvIPJK/lxjfmPPA3
bPWKTIMr+IDzP6OTq3yBYM9loXdUBTdfnJKOakT/6XgsGgJz0jbu1DsmM3hw7CscFIRqBKnVz8nJ
D0V4kGCBlrQbcc8ulVcAuTaLtjKLf/CxEdRu9SFPRDMO3yf01SiQPUZaTfyF1b2DWgeqkZfwZmKp
Ftih1mB5i+uoaDVF0QmIcTUKjUI2rRiZ2z4Mpbr/7fOCuwhRbzvHoHoAnlcQKsss6i6PPlfQc3s8
pKHGS6Ocjh767OJgajdl+KYl24WwMgVz6m5gyOKTzWbXnZxqYoQAe4zu36itskH+fwP2P66pr1ab
hOA67cm2xrXjt0bZnJMxINqAS7keQ1P3q6U8kZljk96smod7h0ojLbGq0tTJARogKvELM/zEF8bn
j/Zr+zpSCxQFUwz33gOtexQJJyycIS49+NMtd9o1u7D0ghnFQOt8TmfNRyu9XV5es6wgk+hqe5Dn
T2V/NtNTBH0GTnjlgVhuBeB1YdRmdiMZ/1DspcJC6bT2VFocurGjOcguzkzIULrNTd3NvSVZZwJ9
N5etBzHcJKPiJg19Y2ke6iXMp7HPXQFkvof7nhy6Ug4cQScRET4vJB+pkxcPujIP+xMp4ZlmTmYW
zlJt48Sn0p03G+T61yEHg8EF4A2Yiv50Pkx9jz40kLGdqx4ampCNE0e+4K0rEU3DYDv6/PEjHNVJ
1Tabmu7vF97maZak55kZFxyRneR62XYmWDyXxKP4v7e2+47D9QgtXknlWwI9N25Y2CwkI4vh4cqJ
JjK8wtVlTNUprzolhU93VgZ5ut/FvXHG/9wmKz+vORNHhHbOiF/znq10ePfjAf7SnRFiW+UUx671
Ru4KxqqG+0gjxQc98c+LpzRJoX8+qco1xpUk8yEQ8xxtuoPf2REgVqDMSEHZUg3XKxOXJ4mJX+bG
bhQ7JmCjruJxglPqMHWNdHgwIFgwda5fiTCFn9fhEda6R0l23NEj8K7/XSF/HC4gDVLtPOcq1+mm
M+alFotspHLYqjCtJe7hietJmabKCF0V0kGlpZqfP2Te+cEOUl0WmKzgyhXUT/IVnNcSjOE4wV7i
E/scBJ1SJAVQ+lusiu+IL1bZeGDUZ932muKAyKY8hGz9RiCfwYHPh6Xa1/udGVybDt9NJXP9FLLF
yjTJq5poF0iiXBRR/giEw5YJICOmjC8qapx8hwATkGMoH91KTD926h8ONAjk5yrTvZoYLhY6PhKm
S/6/XoCucW4MS/Fe+sSI5L+X8zj3qV+eeEoxZVGUq+UMjpGXGn0wSTu579UHLnRQyqO6xqhvkXt8
lw4X7wpN6OTkte0awV08X3VV6g1ZwRzEoqSH/h0cJWH8zE3cFuTd6g8fqkfDA5WlvH+Yd8BuFEFp
Dnd3kR5KrgQqjD/yAoSz2sWYsI/tMGSt55JLHhZglF5471Si331BFKv9KKThfOVlzxbxHj8bUbKC
PmJbcTs8+4WQsYVdtrBiefY/cFk4dga/j5TmcRwX2P/llV4FALwdSMiaouR8VuLMIqGDX2hm0XuN
4O1WsDPdugxOAFJhwW8mt5HltI93H5RLbbZAr+b3sAflkeOp9pLwOztvGn5VsGioIyJwSusiROLu
ITbJSfVD0idZyzx65ojjvCyjO/fG73X3K2NilhuDHa/9ZH1nc2vflGpM0MjVRcjjeILz2L+vE5B2
yc5HEmFWLGPKJkn39mXZwiHrbrsK6Xhjl+88aQ43W5NQGfezhdyUl3+SGLk96Q1FSj5WQK86VR4p
akjI4YT0ZGtQxy7QJJ7gyC/ohvJn8eYfkoWWwRDb82BfEDpm1JyEEvVjRmvwVCTIPpxAyey5nbe3
j6nOga14X3AZXqSCRO3lbqXjhCOU3JP2AlKQ/LImpRQIjZXZoNwmJozLml1F69AMSlOGQYl2COdN
6DmhaCFV3F1JFRUkNJoVY49Eu9yVRKLKKrhY36SgpoH+563B8Utwe7Hr6Z4h7I/g5O+kMZ+ND+S3
/HMfsSKFz1mhXnb6QgjcFZht63qwlpkhGA/G9Az8GbjF7Ssix5/KHRilbSFPzNlFNbBMlFujlQPQ
0bTq+5tf4ScFOcBWMqXi6YatYmjxNar6CexIqVlHVVv7rm7QBZGpBq65rlR8I/uoThszcGeZJpjr
YOg2NvURMJE8QNQuIGsZAdIZ5DQ6RFBgdk+nVcmQ9029B/J7LgK2l40TW6IHbbTl2/cCNiH/jf30
UOTALEkMLBB2lJM92A4UQDuwj1ONI3EvecZQL/HIDPXPQaR/A8MCWstC/2E2/8l30mQ2Pt7VUJUe
F+j9+D695eomPWcrtYw7b64xAQ9YCundpWHu1OpykM/8iN+NQwdGDfgqJ8ey4Sex/f0lhGasexTC
2EHtWbLBmabcEc0NxO83nWNfWOU/93tS5rlgjc4pa+8fko0R8cN9DAIkg7ABIYN3Im9aaMQ9H3rL
TkfvPNDeUCXNz7+cQRrB1XfGBIgt8Fn1+v+ygsjwFNMlZ0v49W0OIta6XjHmpblWynNOfqQa+f2L
xYN/KNxsp9crKusx3jsFBfHrigiyPP8/GT0B1CizyJuzOC7vSTPYxg6RrZufbPUcjs6BGrhErNzB
Xu5leihGExaGE5bqddsRNSERTPxJmHoDFYCqCSxukkfagxA9yy+OzFTnFBQoCwLxNlGH1XusM8kT
mwUZPtsM8Jgjc462gjAGkJHGfS6KcNoGNlcXDCqppv5yFDD2YZoZ/GF838frLciFDqIEhAK0WL5c
QoEC1UWxiRl8tgCz/Vx7R8yM92pDueNqMIpxXz4qkDIHErZEHjFndUyAl1L1CtAxaK3W651vVd/q
rQQUotxVRjFSHW16He9uV1UQnmXsK6a8G7bAaruRkfvhxJMJbEG6o01J4votKiab9FSBXw88WFFV
LOHZx0Jdks19Fl17hxG249IpjRnyf6YKs1FAv2BHLDEhK447PVfMW2bhSG9F5p4dUFUakCA5S6I5
3bzQUHwPEcJ4dFym69x+9UyzAGiLXGcr9rv8BYIpgMb3aJ/p9dMnsvxtJ+e/xsXUVlW9XJKVLBKS
XZSssx/WQyGY5yOswZyfVmHI/UarBIqqIkF+wBSj2RTUIXjd1jomcZA2g18BbSNQgyjgmIAw/jW7
WBICFvpLzyvUIz8ojlyETp3QbyyNRu3/mD/k4ZgfHxpr6TKnr9POaI0g9LduzxOICLfVprG8E/7V
6hO0QFGpHSsrkGzqiePBkYcp5SNjVwkuzMLV9iSK/kdlBbp+ufBkDkOoyor+dIdQsEJXNsvtVCcg
D8NML2+PPIceVjFRrSNQU6RvrKQSMLfOZ+0navbCeY2gWgQeF+PD3kRGdl99rC8Kq8cDkSVx73p+
5A+kkh0Lzihy7o+nsiPX2EKPshh/xpHmEvdQWOm7vHLDAZOlNAuYKjcoxXKWZ7BLagJkie3ppQ6J
LZH1BAbTjaL/10dlMbqZTCAvTbGay8M/ru6f08RCBpe7+GIQn02HT4IY+VSXPh1M/PVi3G6PKJuZ
cRuWH/fJDeDkx7CQabvzYJDwm7anpZ5GEtDtRQlE6QaIDE4B9meTbrsiYEUUKX7JjZx5gvz3GErl
TTVDZdbncs3ANbmHMWMpsZgOvPU0l3W4bQzbeUWgLPAT1yxEST7H0y+PEgXp7zT5X0wStn4IIl7b
9apttiZyWNTfqav4rBglwSLAfwaJYEYB8lHjV0z82A37gifsTfl08WAQDHvdGTI078sUv6LzTU2j
C6mD7gmWvfknmaPDYTalvYxy4Z6PkOC04w96uSi0sQc4M7+AvUs5czoz/cn6zwV4dLxzfBx1K7my
kv5Scw1vkNZpkfGXkCDg+2WycHd3M2B8imNBCzoIeJMRUFrHtua24RCHG9yGfqNGMA2NUMGsskzF
li4iTOch/Mp30N378lMghO+CZvQqylNPzK301/DmTgsQDRAIzsBiSm4uyUC1ELmAJmGesN0SI2le
LvUXy0TzWBA83y1a6zl975pZGEYrJe1OFlGpf3EmKK39ed+eNFiHrGnmcPETQ3sIgNe0oiLakfxV
OHhPB5p8pU9G/lNtJi+7ou5TTnvuxiWMPLXNA+S2EE4z0WFXdTQFjdbIKgtq5lo2tUx6gY/g+U5i
RT1KsN+wU6I12zVTKg8bXXW357HpdLZ3XzaPYp8yKU1WIMWtT4YpQ00930AB1tqE6Qkrm/Ru7MMh
EaaGUjU5+f+7fBfQetVn/iUxSTB3GGsalJWbwHeB/i9H+EB/Mh9Q0dlkW4OsUziamNj5iT8kDM/n
+r+M/q/l/a6NjgcNSvT0FSSN9V0re2AXr0fb35Q0MBV6kWHn5uN1C/C9ct9Zl6+ZQMrQs2SX7vUd
fkv8ox9t8Jupn/D1TEMGN79H4v01TRced1izp2jXbvmbjZQiLQ4v6BUwgz2/3jNrWlA/oNo1ZmFG
vpV2CFMm7Kg3rpJfOVKvtXPDfxdebew8uJoMNIiG51rQz8XNo7i3B1kHPBDixxUt0BaNkpt57PPa
HvZGp8HuPZVCSSguuBzvDj5sY/7rwMymCadHpwsrPMF2z6k3YVbmIQWgL3cGbPZA8a87gLKCZdAf
EH4xCXuwbKVAq18q8SPX0JaZDdsg+wFWyLSRpLM4NQlp5doZfCwqSRwY+BXmFKiHiJf3s+we4pTb
ga6Ql5FXwr1JUZ5nfsdTKTrI2O4I1Kz/L3cXDJ+YkkEhBg+vM5iQqe1Hdo/1D7X74rb0OWRrFLXf
SpXcexDmufzUpgp+Q/aKytcCe5j2R1Xul4JxlTsNzsIy5lXMgkafCd/+efDiA/OPMnpX3UUuz64X
zYtRVbQ/DsPVl1qIo3/sxKK7maPp35/PEtqYGx+KVWN4u3QhosrWP5mc2QXmQey1WKmMNJ86523C
q7e4Uri99czJ2nMOMEF740bmST2czKLfiHnwannt/mwa8ta/rgg65+C8ZmCUSu6cHRvegaR7Jy3U
aUEQ/KijvA19SfWUTjL5nFM9T4MBMAcP4z/80MD2uNKJRfp7l934FliAhbQuD7yA+Z+CSAyLLH9j
PUDZSnl7vtEgcEcvd5kFEfDVSdY2TfimdsfqcrirNCSoGkUICl+bWhCqlgffqTzSGGHgoRC6/xge
qOwel5Fg6+cNffs+ZG9xUqkk02syglKkbxu1wcNBUwGo5jjBRWNkQbobWu27pm1123hNgtlWR5ke
00aeOcuo3AM3sGBO3DFc7USrPA7tq5rdaFf6Gn1Tyj18/fEMODfv977pKMLWmKAvIbA80t91hlWg
2/Lfov+Ruy2jIu5N3OKYjovJaTktx2tIO26pBEEifxfQcuYKAw6ApebCjLs4DBkCBk44jLB8IrUs
LjNj14kVEgL0q9gJgsWfvHihg7T/DKfhTwgNIBt9PS7erqn2M7lJPTw0xOGTxP4EFzgyZeb9Alof
7W+TTcROnBGhIyaPdasrQKcOwbjUNBiekS3l6NqkjdvjrIbBaibMTDvK6il9Fbj2lfvbReVW/1IF
fX2FazmLEDZPEbbQY39lQrkFLuSsC5M3Ers5u2iqA71tQTvXrTB3IRgM2dIX6be155xtIrUNgfQ8
ci+Sppo/7PDfp+TMmBJjHIKZdHJSdC1KcvD0ZP2ui1Av0tdykKPALGy4WyqW5XaYH63ThcYmDOvR
13ZYHVffDk0spUFgq5fa1M4WzXhi4JvQApsxfwOn9C1j+hQEZA4j246S4idh0E0qPQ+TOXuo3ego
4PjxEhvNDKpbjMLHllrkLDiR1EEqNT+xTVxnj1u5BF0jbfJUEkRBNQZyU6uspmNg7M6wF9kUoko4
XZbrvaG92qvvtQH/7k/kMgaWA8qyQUUgCiKZ2EDKPgfv+NIUEAvZv3I1GfDmaBhsbuO6v1S9Juxg
CgYHyeyTAtJd/C/NAiycrofQxaX6YLovsmJ1vrMNWOxg4InjOUap5da7G4UfZt6seu3VZdGoRyb7
oBbTm/NMyFhdTHiTCy4x+JeFhj9rlqXoxmjrOpkPYDd7Piy7GVejFAqLdgHbYSqS1ab9V+duPg6x
urTuCxZExjXayCbsCUTfhm4kBbeQQJ8hICkxgeNuJNXVxYPCtYD9Rw35bJLqy8bY70Ubp+EvR1lO
c0hC+Cgu2yb8A84/QoCXHztZueSISvLDYL4cZI2HHGekH9C+Ti7YoSKjhVxtigFtR0zp5ib3Q49I
uHYb9A60N1+uBMhunK6S8HsHnxB5bsiToYCyIP06B30A4M6Tt9l3xTG0XJTgcCHsFS4egHrf/yFG
R3hep0OpA8UouohWB/sOaF703wpqLLfHaDtXD3Di4udnONsCJOpa9QxXPo5qLH3ms+mxAW6slIFy
6NrdZ3K1xcCM0tuxfqduWPjvu/xKZvextRpO1U/g2EqBbI6x4/7/HaaD4rxhpEAgSBvH3tbYoxEL
AwqgIyWKAWcFFnI5msDylNRIzd28OpD//wUYelPqLTR3SsngO4XJJH+T43oY+EpfFpKAZZOzfM6u
Vv/fNb9ELkL/N6KVZtQTwpuskz/Q//cRRGBaCOCUxLc5uhV/jyNLXqy4SodlTTH6Wnpk70ZQtxnA
00+IoK/+pMoqTF4AH00qwXCJyxTnXj3mNk6WICFgOxqBDMy88a6N0hbYvmjT+iUZWZu0qSw3Frk7
hknVGRqWTvILM/Hu81KNF0O9y7U0vJh4lLKTXGrE7N+H8SeGAdMyN5u/+QFK8mG5tTf5Hcg3Al7S
XJvr/Lrd7KB3yKV09I5M4x/vu0LcFkR8uQfRaG1XXBTs+OG5vRmKVbhaYidhLl1dNF10rusYjgM4
yrNlPzMJrKpIkbibq/wkiDg/bEQHz9TaFJ+lEVmx6ktm4VY6Z3uZ3CpbWHzCU4jnpGy9SsLkhGfH
FhLdH7xYrOo4jOwiDh7fz9CaGfrPEZFuOmQcSlfwu3rtqWfCqZToZT0Tf672TiaQWOrTN0s9n7YJ
LlmMYDRNf/sWfH0M5WozBK1H2cHVFGswQMdjoDKmwWHHv08Yo8e+ij9nmwT7sKaQaPm5EN32zqwo
JL6O35Js2Lii7H7ttHePyGDvdRKVRqxPU2AV29S4Y+4yVJNIP6Tn9w3vTkWr34UiRcniNWRklE2p
aKL/ublFd8I84oTACqKNrV3lJPe47niKbeHs0m/5DovIEEEGGRwcwpYgXLPmPzuR7gIkI/zKewYH
Gv1XBOiY4pc/gYhgpaDVpuokxW2arNXpJUfT8dL+LPNSBquK1QLX/i4FK4u5SLFfzQ8DCtfsGsRx
UG60GV8ia9mGN1iqvLBU3TTdEKFPirqIFVWc/pDgPr+IDksGLXpvFK2R2uZ+ktU00aGes8A1GfWJ
Mz+MUBbcez44+ewRR416EZJ7xIMyT8ZYI5gBDnf9KPCqCiLQ52R8fNANRr1DzTZhGEmnGDqjDexT
WXj2iNT1DcYmjREnvq/ivjohpx9Hmlc3LcFKd+OtFFhNAAtS9gPI86Gvtv/r1JMPGiFOAJuAW//8
yYGa0EXn2N8mzirf5ivz3hln1mpA/p691TNabW9jqSo8p4No3CiGzXFjf3KY+SGSRLAh0IZbv1cH
4G8jeHoPCDMgsXtcw8F7ZzW1qmL5QMRaTolws1VuTum7qzGvsEP0XiJtMlMFVdoM6QsdHZT/39Jb
VVlXiNyAsh9P8DJ0ZnCCv/uohYj7fDOFwNz5QQKpdLcZW2DjfAUuAGm1WWq3rZlxprh1pYlTKoNH
AmY4ToDaQLsoINqfwj66KD+8xMDVHVwMLf7oCTn8TLBTTUHA7xM7nItcuwsxj/f/wZUGmw40gP4v
l4L4M2LKT4L8v55zAr0ur81+9ifdHHh1ZDgS55ydeDcDXsMgjpNrsonsBd5ey6WlOARHLXmGN/2x
AQkvGZO0dOOlCEyAetMVzSjb5DxjUYE4fsOK2TW2ZDBcGpTnTOiYWBLMfL6h7vGPjNSAPXL2yxil
DkKs+aDcjZlEa1SSdAM135UYwhICz3ig/2+UhCRo+dHKu0Za3YDa5Glyu8eK8sfQQ49QEShIRq44
bHc/jpcUukb8bgfEFRRVmSTTICckWptbs75YeieLI4U9zU6IYqjN5OjyOyqVQowUyZoxG1fI2uim
DnmgK+L8S6u/DZGZXpX9dt+aRUsK2phR0RwUgAflFes6aYVUaA45GTHkcD26SYQMRsQLdqOHjRH9
Z5GIo6fFbU+/q5wcUeP8104R6x0gPeVJTr6FIRx+9aQEEOYqL0+GEEVnFmlNOvh4tU0eHpG5xkAs
l4j3iLuhlponoVxH1EEu7wNTI7E7z3QSsLmxCpkOtZjjL0M586Ou1AURUbZx9Wtj+qJmZCEK6pHH
8waxr4wKTZhwKtRbVDLDP3qdUy9yosBEPLGpf9Z1As1ccEMSNrQwOEcspvEyDpzTF3cCV7moOmF8
sUgM19WW/XbokzFn8d83mdHt0zpEChi/d4nC1ukwUtiBfRlFJH5JfrPLIAFjl0+utqFLq2x4ch2/
3qudcOIjPF7XqLrTDjnsXu4cvW1Qj1D4QuoVvf7doNcZ8RIMQLRAPhXhM5GHrUXR40fXnaRdZSFm
ncm3eyCV/fdP6VTi/wx//LY2G6W37MlEPoZD8dcEx0tdvaxcD5o6jIAD7cbITUoeDYV3Z2dwTfak
MeLDEDvSA0txFvMrD4AO4M5+TaVykyAQPPwnYYU0Iuhpcf6skhm842efH4NMVJqjMEDVcrmOV0C6
AZZBocCGrEbVWR2WhLvQjGquOgwK2cYDukCXhPdboQNOYJQNuHBoxOQfSRHL95uYIQj29Sum7nCj
mKCq3N2rrkpHF+1zHuD53ABU1IrWset+E8VfNiCEkiNqSQQHtp09Fmw3VUm/bXHzD43UdULl3fXu
JAJJ6eJyBY4Vbd+3x2ihj5UfipWFOWoUgr9VyU5lC2YcUoT56QNctdtF4cICB7RbDIXQ15d9Nzin
1jRUJWsIQj6OZ/nZ6sPP7DNMcSFGt6HpUabZ6P2+L8xzTaGqJ+j6+s0/k5d+C/iKwpxMy2tLelsW
GfHUwgRvko6E+ST5OIUSYJdq+0Dr+cIc7iUIF85+3KiobJFilcScy0JPpSHpl3jyZ58ieRlz/xNo
9O/ZmHAUuLlfjjV0NDcNKU8/EiZpL3yLP9nihfrImc72piLx7W78GUswIVUziUFgjJ1pybNUtEZ3
SkHSSDapRZdJ0IQwC2S4PHiYz4RLf4Rt4/lev+H6eZvG8ZzKKGj1io3idBdLRVj94X0SSblty6an
mgkAGo6NnGAMWEec+ZroybMS85lwuNso8zmsAWTgkN/umYwFAbFxHac478beRejOUcePz+QqgDeb
YltLi16hkRg4vKSKsnpgyTvvkD57cRoe8CF8vnzxG6qPJCh+mPgxbpcp5Uc5E1tf3aVz0NQJWhoe
ynU8ek4eben/ktn4Wesxk54UsH0D/HXwh8/44TELGVVspETIg2xbO4I0D/7IK4A6C1NrSVJebjl1
fwuzd57kwQEW28l4hJyXjL6VAAVrily1ZNXDDJPDPuDEXxsLhjWpxnBG+QCyCv6C1pYx5m1pntDV
gI1motBoTkM0ZfYkjdE4op5Jq2LUM4Nsh0cH59Wbkjc+qr5O8ctXiituauORJ+A75Gh7GZbrsAjv
dYFbovSoNjxK7MBUariwUpYSBcBl98+DLMHAhMkl04P1HU5x5nRgkiIGSB5Gl9KgHrECkldojcGA
yS5heH+7I1yIktJsXl226SI7a00CSJXZfOB+USUbbg04vP8bg6ZRRUZVs+4tAb45IRLClUWeojRB
67PmmCsM9/gnpek2i5QYKh55gftcXIPq57k4FfPlEomJqhKDyDu4kHAQIC3Lp2OA2V/chU6g1Eki
hkAGSN3xzkR7avPjtfb2kL3hCPye2URJJ0o9bP5Yo4b7zlWnQf85RppiN+ypUF/k6uhI88GRz9wO
7O3ficE6GCZgdQHyBgiMdZyUovLgPNxFCIRqdou5GzjbY2Q4236jy1izxzv2zApF/O1Ew5EX16vb
AGzupasw90wE8JihvLXZq5nhKdZl524Fz2n3JtVSvj2OPbM5AoaVGcnO+FG3uoWc9QLYF+sK2Ofn
BAizgBF49Uk5CNNbgrMBl7qPXxmvj0+ZDwjKiHfPus0/bgFJGyO18yxg2GJYMUFD52jkLJsbv9Yy
j/O9fv1lu5N7WzkTnb6INZuguUNqlA7xo9FPSiM9k7MGik59Tw/69+nbvCUV58iQqos2X07ZgthJ
gT1LJW/I/UiYl01GWv+0EMlqyQ9G3DSqpI3rxzsuYdQBoY9G0I3gq7hb0Z7JGT7fCMNzj4fJUqBo
9NzIf4yRiVyFwzAl5X3q/Kxoh9UJrfTPN7Kr5KFtKsNPpf57N3Pq6b+nMvVgRGFfpHhEgu68OmNG
H7pfhp3tN1OiYPptkCrr10TrQafOtop37OP9K1ocm70PHawkhzmkXP25phDC25+FZphx9VWOmVjW
u+yIV+FHgEPy7YanqR+L3xztnfRHE0F5HBETI4FISkb/ZruS4YVeeBxcshuEgGf7fO64vIkRlMbA
LWGbYPREE42+GhqpsP+uaS+hCpV7AyMz/lLH1G7FQctJe8IWVbykMp0oObJ+JZwo198YioAiA8l1
N2wlyLT+uqCshO+9q5nFs9otHmxrYsmYiljF/vNSAJtusvnWkxhah9lJJdWD8118XQdoDQ99uVwN
Q8rWWrikH36NqZlJ4czOUKC3WN8T1sxy3K9g5yVfNfqaPFJF4lUP9tHX5CDwVqOaFHNskb0iDe5z
hro6SAWEH9OyyeU1wEn7kzyvl1Zaa7C0uz4KP/7mbSFOQlmDCiLEszrK6XIvKFB2rMB7RISN9KVp
e1EufHM38RNq9MPal/VeSdiqkCWHVPoYM3UG2CfbCnagmFA+8Xx1OVJXR36eZZgroSZ/BFp2dz6P
anpz3/BnNxd16HjYQYUBOQO0kivIpkAHbuM94X9N3debH3dDHFzAMLBjEBR9etC8d4+tt+4RvrgV
kBec9gmKtSSicxxoXtgYYG92Ubz7GtMo1LthU4Rn8HfiY+weqQiTpRST5hTyTSD5FRBmBQ/RK7Us
4ZgMqs0bdlEVrsK+loxCvhmKWnIsyTkvUTDpuPDqdRgOL2CtlVP+O0HVwGBzPq5+xuv0ZPFCzZ7E
1TVlVBoQe3M23m6Gg3DzgekpL6uP+EAjKeJI77qgj2V0V5Yu1ELeY1FAaY60TFvrie2f0At3ExB6
+o4Pz5p1yx3r44Lg1JDxdFErOjVpV4QzRpWbiqRalbiP+9sueSKtusPIRluYSkIkZg55kMR7Ex6C
2HMRWOAukEr4Opv2zSUOL0qyBkhoTF/YnCj05TbWTBtHFlSCK7Q5zqU7F1mcRkjkcAZT1tln6txS
GCWyW2HWwkkLpICDHrjc+tE7uwvH6j7Q8RYkZ+vNEltloHgT6Ri/9tpTrEDOXTl8u8dVGiD/yMDY
ybw+Z26ou3cqvjS5uGzGVlm5bRETPhKQrxXD6lb6GyUyzRcyJbbNXY3hHfaoqkdlxu9ep0nP9jCV
MQVz5mmJ+77NeEGgW8ohxSVGynn1f5WVZeUwScUdC5q5IJe0mMqQbKJHdt59cIHYfH/Z5usCxclf
ZSqoaC5WliTRgWN0MlxIdr6zHFovOhS8fl71zskWpDD4dcV0wcJcr8f3RgLp8OL5wguyD7dY4XES
VEZjxE4o7R+29ELEcbpOZxNBRPprv0OjcIzBk8qlwzuJbrlXtVXy6hiZ88aaPP74759AJjwDKwCV
LMMgCPE9ecjqyvSS6qJhd24hFycPP4fPeJ30RsQh5q+1EeeMFGAmJ2J+GoL7EKNik/zz7fzpRyIz
tyisQAHf7pecvYLnoCNno/UmgwnHaRpXke9DS8xVfFm/OXsxL42NQ9Cnp9RDZTgxJ1ctMfC9eIw5
VZYGMjreUz3X4As/bURrWSnQUqlve57mFY+l9H+qJ5Jvhd23U54qtjQgAsLeF17qOpiyoUEBW3oy
ORaDGEm43jRz+52ZqqhQ/bM/bSnIymwdbpf9wzcuJbnUTjSxlPPvuD1KHDhD2SviH5dIRVwr+aP9
sWK9lBUNH64FngvsBrfMQnlhmqUU3CWsVFI+fnmxZI3IgteZw7Ih3WLK79AnbCkG5irV9fiyCKSk
Nqi7Bd9axstW8cmzYYP78141LxivRgCZOLpkJUZk4kiPbjV1l41A4PIl0AqrStWx3MIgYUYzGZLV
/fN4PLAB8Dh5BrwNrAMmkO6/sky2GDeZw4RS0HFeE9nA5/5o2ElgvcLlXgARTd2VK6XX2iTZ/VbX
uS8j589a7PBoXh6J/FFPsHbxkF7HP3nHz9oziA2zHv7P67zUH98XzQwXjv3GxJpE5kttqeKWWZ4N
PZVpcYsJ8O97BB9shgBPGiUDaItyc69uJht8xC07LsfVLswY9+4PTkEymLO5pWX3UgF7uYKLPf8K
nlfJWLG49x6/Db2Gbe3DKOnlRHQclVBvzRhkJO7UodKnvYtm+czWXdPedKJAsYSKQXo6g3BnriUd
G1TosRffSRn3raSuH9wk4PO99kfHXRsu29DZn9Jip83tnJrMAVR0x6HevxCWQSShgKj5OzLzyl9U
yx2vHl8MDxgVD97DZ8UMDnTOBt+LYytsKYnSklyTQfG+SY/lweOBmcbUyhvvsUsUpMG+0TYnOBW2
tmPf/NFio6CnD6lOKqFPEqWoMYLCIdIwaAGMnKkSCt+ggcDQVYsGoEB1IwKcziWBXx88J/MICOrO
FQjF3LP2lAI82A9xCyttp63Ee35GCOuLTW02DBZ6QlPk9nzpeBdJD7fJGLaUvwQKAiM4AdnEeF/c
j7dv+q3r1H3AECI6M1sX2h0LyVJYoXS3dxvU6KpA5udyEAcaeWXeNLFOXe8XIXpW26hY8zwBzsmJ
AZsufrEDLLakhDAmN+WlIF9sUMssehh/67zuufcjRC73SO26IewzKXLEvrBF82NX9NDOv2FGzWoB
LwU2GnwSadKz04Dg4STyRUdoDgn4WU0C8P5jvmVVvCy6+kM1wY2hVbbomTYuNoyFhN26YnS7s3BE
bs1tnqMyT6f2S/3FIY70O7hZYNfVWl3z5kaEyTof+fTys5t5aFfSWJrwOooUxiHVaw1f/PbUbmtb
68UHdMOcql3WWh5NiWKf3OG0jl3Po6KsyITC2GVbwiQmr1c+Ru5GQFukj3E0RXJTGM9a5eOkojyf
7jHQfnXZvuDid3delX/mmOir4XwdvCN7tr+glgaukIOkRbopYjfPOb1cuzTzPA5YO1ldZWn1a7Pw
2Qxn+C0cKUkDC0NlTJkUJT9ZDw0TNxyPQuTW6K4pybqfiX2eWIqUBQj+WGByPquOR40PYB6kQzl7
t7j+JWc2pkWpJmyX4P3wdql0Oa9FRRnNOPjdlcMt6uVAtGkrNKwKuXfrXahU7huca/swmRfBHu4Y
tqoSHPYivIpdjkvxV3mV/gLVmkszJFq0IQ6J63Bnu6GkmqTr+Hqresam8ukMKDi3HUXgkfx3na0S
9/IBeqGcf8x0xD0SQu/KitXEzVeLM0loKi1XDQyWlnpZS9dDRFLuui0b125dEdOv4vCuBU9G/rG7
xq8Vh1Ar3tU090RID8WecQyo5W73f3xRdsUdLNGaSi+2DE9jYqldui93MwiJ2iRCpyPVO3ut3lN1
KfsH6Seh4jgaLrKncb8TUVmpu8jV78XCJ6zgm/WjRYTmn53gE1Y1ngIy3yEhQFU/sI7WiEhXM8Yr
VQz0/ZCCiSeplswziY5LPyrYa1wIOO91qQQQeyHNJ2LyUkmODFKItluT5Cl448xaa2RFjv7HSdbk
I/2o/P4emUX7m4kg9tmX8J8Ofj10ineUFG4Laq7Z9O9X3bGt/qwbP8AiyOwJ4vYU+ds/icM85K3A
tass6xVPJLsIGgxcgX1g13cX353HZzJS6fZ99WCGw2JO2fE2nK9ENrXXrUsy5eL5a/H+AoU8dBpC
ItNG3quOJPsznmF36+1kfciMQgHZ0RrKPuuIccEz32ypHGHeGWv8fgyCjg/LLmaoeb7Y8rekALsr
YvaQIr0NQKfrBz7UaBGFUlGsM4efaAbb6/PX7c8ZBWrGcGkohWJ/Tv6C7ofngxUPX5xRU7NXIcml
RaHzGANw1y0v726E8gHS68D+zeAS1jK4D1+MPyUW/vbEEguGGhHih1K95G/a4Y0idjq04cdVOL2E
JLnUkcobDPokpZ1pQ0O97zUKgyXUH8s1ytIrmT7U7IPLRHtUiaW2nYizd5tp6hEzkSIRaVAGq1rB
qU/fExnBXN9cffFu8mg/I1rPvJOC4mzBskPNh4xv70piWxV7JsHI078WTgfzRhSceUJtbgps8xcE
iqOj1bVvyEeVXIfw9LmGpHGiXannycIgptgiB8lL1L4lTlvQ+vV1PXgivSfxC75tblm8rCF0XMQb
ZeCkN1TKHCuLWGiLLkRZE3B1vGpsTEbahk8TfchA3g9mNYT6uWItlez1CrjYR3pOw4K6bR2N5KuI
+hH2Bf4pj4JGzBQpXDGwCfd2uIHLqSTsfz7Zf3tJznR29cLmYUhbvnCGwIHd76ol6tUBuCKUQRRM
tOdLxi8SxIs8zgkn8aipfL3cqUJbO0WIh5fzNIk24bHiNXZX7iZwHWsuFSbkR0PqRk0EekwiLmI8
K5HrUD19J/QOn47sw+ofL4tEdTIpcOJsuF1zZKIipQgvOPvqiu2rzQR8DbpD/VC1BOkeAB9IltgC
t3NtwrWZ8iHkrF1xNZW7U34+02zVHjLy/O9LWJFMFXMR/a5XZOXVH3qA35wpsG4p6WTFmOuCzKj/
9464yWGq7vMYylis3mYO/ITFDaFfjZ5Z4qunVzGcdRGWjIGNASV6t6E/8Ae/1bVTVTOTQ6HQTcq+
VFy5EmTF99D2v4m3iIKTE1bRHqIGLsQ53wA0lA0A9NbaUGPqR+OKb7TtyEDS+1XEph1AH2J2i1qy
Xq5P3Sbbxz1dOnYEwfMjIMNhAM88ESlsLgElz5o2ulhVvafPXesws3Y2TdssxRXLH/QDmQ3cv+qS
g+LPg4I6ZWpjfVZv3BLYlJJzt4oq0dVj4eHetImrJ9XHbuhSXS4l7P2IRQdAsMitFPzrsFmsDaBm
pSheSbO6M4Ghxl1tDYz1rpIW4hpeSvPOo0tqZ+8QYanDvEYuKz4X3i5ILtS82bFs5XXcYFkJYe4s
dzNQtmRR244QZPBKTUWfZUF29Fk0Uyt1ezY7zNgxXaTlA4AXc2eZ86bJHogfC6vvwBrEInfl1jf+
VrMVFMgZZzmJ4Cpxr/XpFpnFezqsBW+ZPKk1NKWR31f/rWjqYF26OCZAQ8n/rJ3ulnSBjbUNBCdp
YVkYysAaTC7ziDMne03jtAF7HwNMPWHEA+LWhUjRoO2bVugpXlZy2So0+DMkgjj2YSQ04ozvTrRB
krpQIJu/lO7UBVagy058B46xj+EAOsudYFZ3hVL4PVkDiAgFmZxvo+OPfW+himHFi+X1VvOjdnFf
LPcJh3lkGkdHBKmiic6eOJHuIhny10y3HBFzVujyuNwRGlkr57cUgggC6IQhgPNdZR4ZKvwEXoT1
QNgia/JWs1jYLjz3qr8GV1dCEt5nBfBQSls0JLPYSlA5lm4NW/Y0d/XbJJ2dM5XK8mYNvW670uHr
RApHlO4Fazi+L8mcBdB00bsUhbYmtwVtziK2s+oJWoTtxOc7tSHjpXFCriAnIsANlJOv2JG98W/j
sCScecHjntcoEyEmR1p1nxcSjhYKfgg7fK4qQGfuYnWcnXJ4G0fTTndlUBDjFcOaXOVX7D/nB8aI
b5JlT24VEpSOK31s9A6cQcVLLD/kwsjbx6gvyBczzZvWkOZ+a3WSMKK3avEUqSshUb+M8TbS4W7+
iWfGCFNcaBaIkE7u8yLJxvqyPtqOHnpzMFocj3irCb+9yi4+DNcEgpDWkx0wUwVw+T7hhCJe/Hv3
qDWhXXdzqwb+38HWJiOwHVRxgfej7G9kVe5bEKFJionGVdTo7L3zYzT1L1h/UlppgBVERnzboia1
PtQ8Uom3U8Bcmmrlp/wSmF3nRjT1MpA8eUie5YveaBFt//B5zbDe6DMwi393RmgYcCvXJzo/mEh0
2yCK7NV4sV8mRHLD+L8KRXE9BuzqU3hPdO/oTglKlHgmBpLD8ciur/kOPhqqBYeDbtqpnix2tTWj
dyjH1+pvzdvGatrRf7zTJ0ZTQkj3ALBtkqkrruxWcebMsX+XkNp6SMizGvrBBGoKZjdYdcEvpqf7
gl30iEPkukX6BO8ZaFQOxFEZkZ+8dEzyF7Ea4N8A9I9O0kqtIRiZyjNXa2PivsdI5goUmNmfjg0y
w+vEoW5L+gd5QxlymM+BzsTcVnU+/52Zg4a4E+rVYYsJxp/g50IcZ6W+JtscyVwy+kFwSCrTJKDB
Jr5rRiekUWzm6b7e23nub5F+k0TAytwfE1G66H0Sm+HVnkJmXUeKKxPKqnc1A66ejOjX7j8L9Xxi
VKMt3RkWmxQRZeSrpoMC7njJTShZCbou/yi+OJKVPW75BBWDNsQLvw0CGYOisYiuDNJBFA0qJrTU
dZh1ZRmHEh4iRF4QTThtn9uj22HfITPyFcobiK8Zq4JH5ZXDrKM5wsJZbs7Vl2hP/qWyYXeKKtXQ
0QB3Uw6QqvC3OgzAvycJl7QqvR0ZTXClgDza7fn/ElzOSbOkbMCIHdzPmNY7Mm8JMx4FiXYRjGZZ
GXaVav14IgZc8k4i6M1m7w+QaWL7eqCeghpds/kQDWqhwooHcdQjaY+p1E/N8iNzI7Lhem2fjhXF
XoOD0zeGeCJq2IZSMBghDqzp15iXeTG3raLi1Sy6/thiSIcrOzcAldwfGM5+bgreh1eReTSmd/TS
T5JhRoq8gLsHQjw2TGzVDbibPxPBrG0Cj2XqgpGgn2HXxYJEx0dsgfpSW/b/0R5VVQv0waWWQDY1
IAmngF/fa0kryJayN1luNuDTaGyAFEMtyWoBUSI4MNoh0TE2K0dwiL19BWSgqVKDeEeTSAbu2XC7
zm6R65N25fMi/86Ip997atOtISNILwoIqEMh6YmWZPI4fnGtjMviiQEDDZl2EIXnS9g86lLdnaeP
0yYz5/UsAxVkrnO7pfpm7tDx2+bz61kJ81eEPwPnGMYT21mnzK6QIz39SEPB4YE9wFRNc78l5ZJu
XZVGunoob4z3QpV369g4YmIOnpJrAYhjB3VHGSOU+03JLE9x9xZm3vfaI7RW4I8LU3Yf3S3KIc8M
MuWeIcqweeqS/v9+JZvizcdp4nKT6NYVZz3tt/Y5h0/s1ac4KP5KDI97u2C7WM8H+29x2r/6hhZx
LGfTh/ZA1rCt6H7voZhKqvjpeKBZQY3sBo56x+MrXsVHxizbl34VcErkI2mD/Vd3hKJpxk98Nu2V
Ad3m+p2KZsuzv5/alu2hMbU9Dbu6DX4vxs+xkZxuiWXJMCMb8yyUkMfQ2x8OR7gge49l4zcddhxD
M7QzDavrfUehfTwgvmNRRM1CvsKzjr3Y+XghF069J7AtWPP0rG8v0OLlZEl8IkNRp6K1vIsHPC6O
0O27w8G7Um7yJnOYDFGSH5WvgsTtvI8kVakVjoFsCJrGG5mCmwn5LfIC1AA3f2UBmLU7LOefejnS
734Aabg2j26phDoaJ7IlPQRE1SycAGkEkFnfHdGCB3UFEFyU7pbws4eL6AHeIeWKIlDbfWI1Ldf8
dCDMTMhmo+EA4IZ5FqlMopJXMEYlAh5O5Wmr8Cx1T1i5H0ANptnKVuDIdEfiXyUppfT4CKIHYlzM
kQLioN8vdsSaD1j0J8EStY7rULo9w4hLCPo64ZJk/ruzEjcM+d5q8NaQseoTcOhdTYjUo87zmWQd
BCbk0Cnxia8Q4uzhxT9CDfZv1X8xTl44UvZFn+P2b1D4P+EiXijA9/7JfP/OFpxN74DeSN4NtSKI
o0moHclDB0o4RmvkVyYERdHHe0aeplIaYMaULfLOwKDH+tAEn9Z98ZRY4wNTc5j7MSsUAHjAZIit
qi3fHniC7XcMbYnPWv5KhTG+w6Kf5E1l8mtADqv4/QJftvQgp8iQI9UJMf9BNgk11OQ1IOc06xDu
5PiXgJDQ4jNVZ7XSwRD7XxMnQCoecg7wMgoewX0+2kst07rIklrUGD486iq3+aSNr8xRVfD7jX8O
5Ywb1W8HRGxV+iBrGPE5PAA/CDkvfPsxcwostf6XNVqyu2QW+q4QroQImz3wciPFFhBbQrOaRlLJ
EWNQ6aVSG5Zr3vlB8gO0GuqEaYbwnRiURpQSRvpXsKInTV16SNVKSiborJXdG2kWN8gaHk2NlzBg
6/xgT4oxN9qr6fVoYg6FVi2XhB11MOk/9KRmCqKtiUrGVvX7mH1VtbrjtgiFLHuEo9+ooVF1EF06
ORcFzcm/4UNPcm0ptXfuNf+ftsbj7zbJjwBIPyzUmmWbDtlSTMOlZscH1wkfKmmCps05wBi0zcgF
KmKCdoY65oztceaZ/bbxYkIXc8OutRmMPS5zB1zWCV2t/xWJWCyxmenz7Zj9TJwZ5+25l1i/9Ngj
ZcnZMaIF4+4Y0CyvY/TP+etUCcod9rQB+9c6ph69vjN2Q9NoG0O3i3FWhPPehlur1lvyCLZBC+M1
X9D7eA9fLR1g3/fWtZJddTpGQ9gxAJhBLHTtt+sHZX+emWsTgxC1ZuZil4KibFqSyS2Ve9C3Ctti
4d1f4Nm+HyGGT9sf/PAuBdKbXl12YPPyd7DYbjES1uFY8/71K648geKNcmvv8Kbfd/NgwqgNIPHc
nKCjtm4HL6GRF0EaFH1TJ9qc26mIUwEqcstqMNrrw/SNRuXJ9x/jn2tf2+KEaRQiUPTDI0kCn0T8
Sjw7d7n6c/TQacdjnu8dvVZs7ApaOd0jnbVbVUPJXdM81GJt+esw9b16TbYlt4VYrEQnotBFLiSc
fDa6B+xZBlXxZWiLJdaZDC9NfMINJwwJhWVUKjrB9gC2IjR9FegsbSlKV2trWrOzvDCnn5xDZtYI
d+71eRKwe4iEjVDcSESaQI1CbfHGiXGtz2CQRUfrJ4pePGIjx6j9MCzUC+KsX5mcVLepOBKYbOk6
SFsuJaTvcpA1LNoRFE0WwCH1iYB/1+unj31bd5s87a9uu5NxJvo1pm14sWP+v8ViYGrNU48tgZZG
Oy2p3PoBjHiLIGv5X3ayD/vrq7xQqIBdyMn7NaHnT/MESzgDgIhhXoBnUxgyCYT3tsbRYSRBGLLQ
lAaRpQzbne/YtH+eY0Z540Uv0Jp7rCfQkccIfUZBEfPKeeCJxKorimlZRORkR33iAPk/WNI78Wv0
NFLnglzqeXVNhQhsYfXaO0brgRMm1odRuBKocHahtLFMBYoLnBL2UEoaonzUuDuN2QVk0Eligvr/
oqhG338bNwigHwiVJGoWgaTiOLGAD++oA7XpTSh+e//1K6mso16oTXWOn3SrmUwBoutDZCYfaQuc
Z4dSTxIK/tpDnArSZiHiToFNhB5aElaVj2mfNGahFpQH+1r9rg+wIwD67HMUebQzFEUBXgztcMnI
khBjn/Uog9Yn9On46HlDFwVCDDyakWWbN6kFKlqWusiMQ4oR8D9rel77KjTE7oaUhikeX0B0//2F
hBk0sLwrppzkY5GZ9EG7fzXT0IPyTfNRdDxlVaQ8QXt+TPAKg37MuuIRVrWAM1KozEMX2gS2LDsh
tg1ygp6fWTTHMDc9/9x0IBgc3F6upQKrQYeAQWGUBtzpkEO0H0h1z7tGFlw4BVO9T4HI1vkzKPH5
L0LEAe3sqsI1whDTETraw2EPt/3LITtrM7I/KN4Vxo6GYhwBuifMn2nkPDFsmSqmuyqznhpn2Svu
QoF9zB0qePo8wfcFZIYw/JYTU7FszcD6GqTuMGG+GBi+ZNCQ9V76FZ3iYhnWMvGmeEdUtqVQ1LMx
fqiIg2WNFFrtqq51mHzEOv1XtMHh+lpiG/I6eW82Y5s3plN7qyq4teOVIcK2XtUwCS1YK8QhgWkc
nef/wOhVelNpOj6C7vOJCDhIr6lZQqB535BdRos5g1ZF1dxZeAX2ErTEYAbUcb2iaxkuTyyYQqni
0PRx1BaKskQdua5cZwIycT/F+jTmgrOykufOMTVX05PvZmp9HUiVHQxogJbcF/d5Jh7DNWvDghBJ
OSMe9XZwJzHsdimDBs1mIQKVdH3YieUi8Bp7YBDGCs1SJbTXotcv7Wg42XYFWin76xtVhwpq4v5C
H0VPkFguXrYvWhhyuV3zmEXjD6gSb8Hzf2ZKb8DOFlpFWfmR4Q833Xp4u+f14SDAOF2A7/1v2g0k
6GYn+/bB1mZT1ZUa32oCMQaFJwbTQgZTWrhB19ZZcbaCfQRjH/jWivVvwYBECuo8Iz7ODSaZMMi+
q0q5L32/k6rbxxYEeO9k/KN6+XkaUnJS8nrh+4LpKcK0PlNjDfxcUU4G0SJ5k4bUfJS9R8lhl7AJ
Rm6MxeNzHFIpY74XsFhZ/mhNfoPkoDzFNSA+OjzxeLsUkufcpkdsm0lztHxfGbskb47FJIQsyjMF
x6yK64ZyyEFhKnfqGYfrWxEa0ZTY2ObP/JhFe6Zhf7lO2hp6J2CqP0Xj1hOeInV56i6WN5PFo4F4
iMql2SN9feNCWNYk2Q0SQ7hI2Pnlx9E0/qzWTvRc6kDr6OrQEwBjNLM4tKQNDcf2y5DTKfqTdGR6
cNWQA/sZQMXBC3ZXbQdxoAfElZYrz1Iu6WIU7oaqF2WPw7U6w3feSFXfy5fQs/0ARuegrJGJ1bEs
2oIhYEwPCt89FdAjslMS9EsvEUQn+/8cRSnka1aeiPqlA6mopW7/4SKo+YdO6Gt6Enn7CeT1L2pR
zCSyzlvRRWyfqAvbxTHa0A/rC0C5Un3txQUh48J29FspQT5pOgRtEGuTokvyBknWjqXfUQi34wrS
i4PaVi3zk0WlomEiHN6hHBoJkmi6A+sh8hofJGKwbCxj7lRo8MCnjMYzKQeCbdeWe3mGU5eue6o0
cznFjVRp4DH/8b/v0Dl/jKPce9ZvPvwJozd9er4gILLF3o/Ii5vtEltcdyIjGlfDS9cnGCCCmiIe
xLMMY+WC6ycPS5vL1/qw0tunDnp/XDGATLzR+LiqBYXI9wOy7SPl/udUSHj0R98N/dnnWv0fkjjd
in9otn8xK0OovdnlLnugUl4wcTFNECLFmUEJq7EnEDgxuhk/VGqU7m14+KhL2Q2O+QIb+pi3QZFk
9pnptidtJqGIMp9ZcDMG6KPilxaiJHnJJ6uXvYb61DRgyxdL+pQWT76TSoBON5hG5jSXUjqADBPk
jcRYAGu4tyYcpqyZk80urLY8nExqZ1okw9VZ08sibpjayl5TMW1HmPXqBn/y2bsZ/9FcSKcXxqZy
qK5hdC/EQRsv51skurU8wpQfEWERLtXjHTcMumMuB/zlP447VCYELIzQwjUpAOTqYAgxGOoCw1Rb
m3WuERmIAQFa9NEO/i4m/II+I7vZADn5u1wBgXTQzW22r1N4abSECI2AQ5lMFf1aYbdsTts3HFQo
ftXiD0DTpf0JHfUCYtAw9DmijeFp8rBSZPhZt38IIbF4vEUT4y6SPItwP8T7mkHJD5QqNWmk7n9c
vigoARzIRBL+VlOpIrnD+ACeSyrDp8R7UE0mot4hxqtmmxoeEh9Z5oSN7ska/HYFK0tKWFjFbSz7
KuHK93QS3nwzgVqMCXw6/7+a+FK/pu0BM0HzoJSVO99Z4dlV66HGwyUyTwl/QkUgpM/XHYlVjZ2j
F5TYtHGQMG/CW/vzeiXmoZrWwfOo/GKVf47OZJwszwSuktc7eixDMuQWjiGepQReDkRZyUxIiKOu
r86gkeMT9eS6JypZs0COQiRVlLptkKuI8mJt/e9QzFfqNrFBaUydQc9WcfZRwCE3+hXzofYiiQLf
Fj2f8bbUiUlB6feMkYBqssuod8txV+jbVAuvBKjMMuqyqkzSs+1Nob8EAi1MbIBizfqn1oi8xCH2
sIIfnJ/nGjA+etEBfrktUaHq1jt89c5OcgugOkryeCf/DkbRC6TK6zzLlIPX9i6yNWO6k3cs9o7y
zIEpLFP8RJHfyxDWLgVUkdRSZj6NdBvPz/h2ipejE5J9WUM85852CwBEOCizaUDw3uqNTCg/Sxaj
gQDKpB7Of4kXYlZ0hLM68t3YeXApoZx7MxtpiASBL+TGiChc4TLxs8MIRaddzs3Pji23oJX6RcFq
jBvtWxDXOXCUyOMaDpxbHdFhNJOef+jc0P34ACz9dOVLowEnSuuspRm1VweDiOC4+wyJ4ZKHfrDE
PAwFG0tHNE090TK12u5t7buh0IiRmmNoB0VVYA+Be0VD5SudxQcpMwuHhxdY9wExHsKsvLUKBYXP
HeVvGYOpbA1ETKYQK8+CxP8j/+7DzZhJuJDexKnONUsAramx+UYgwY/NAC8dXAd37lHk8cyFwSzo
ioD3E3ryjD7khmjS2H+pbsHJM02WY6jIR5Ci4sPeqs4559Lif87MfNT+61Orb44xAL9hK4Zur3Ts
PGNLTsm4ffdgjZm8k4anjcAvpwcKvWfq/PnSFBqvDABElZ2aZPPe3mvEeut6Xk7XZWIaShjrgtv4
+jp9yYmfq8dUJxu4JaqWnO1xNR4ELNHwZjZpGGlH7jUMXi8GynL7LKxCqEj+gacTOl9/MHa16tmh
19W9/qG7pgr14Z+rG5ov600CaP4VCA1JVSwkzFbjBZkdrrVGdV7+SSOOkNQgjmEXsgi9Hgd6Kd1O
VnShsZF6qIAJAU/924DypVvXXgYO1q4Ne4SMgL2PhiGQvws+kYbKcrNc8iJM/yZq31XOfZs5ygrl
wx6+LITV8otelkBNYvF571tDeV1tai5vQvq1nR/simjKjbyhUJTA4KUBC9TEtUJpr3MYHAB7o1FA
4HHOAoGXRVzzayb+bTt38apuXAidQmZHqcpJ3su7he7MKJJ4WVH5hRAPq1GRGBjEanWgORcRU+vD
tz+UPGLl2N+YIC57zkDMzevImEU30H3lPWO+cKZc4oatvZ58PirD2jq69uVsp8tLrQP+mdyMMXE3
4lwaoPsi8IzoU/w2ZYxgzMm6zlPJU6G//jAfwzUEt+99bywmUcZ+gv2TzpTfkrtCqkbR9rvBm/6P
brCb79SW45AxX+4VsskDGCvHbRY5vqw0uf50HC6rWfOlqPz2uUHIyiqGcOGqz0LFNTTvSFZY4dsq
fmwitZhpqdoeqcU4SCLaHRHd/zZ95hLbQjY4kgyqNFO7o4C8dpoJrO108T+VkXiyxzRfN6s9FVPW
LxTMoJhPOM/MqIbK2rbDM4XHoqMMN1QFyrBiGbM0XiqBbRnV78MoMbo8347JiCqD4vKNhYVWTS53
p894c9Cc/o2nduk+GyQH+GbBsz6OrRYsu9dHpg21SLPfv4O4pyZ4HGkK+J9mPWvWCM5DbWx4t7wI
qc3hNeLs9dCRWdJT/bR4wtABJR82YtstySQU5XKEpiR/xSZUxJpUEKZO0AirKyvzIgbNxqCJqQb+
GNU5vZPCczvpYEQJUeZkLLZ2QLSTMIpdTBFBvljdylVwgyRPZ/YgJOvDBaH4EbXXxHXZwA87fCoQ
MmweQ22ypGJqxlptTG3aLR4HI5V1iW8o1NSO1+7tw5e/j4uddltR61oaXNa8XEVd7sOf4Sv3RSj+
gMdiusGw3FrbyOWIB+dhiusqI8siKrzqoED9h8k+8IDHCd1Un3rn/sijWq66yfzF2dzOOgR8/rrV
52OdKK5Z9Gsr2gEBIIrokCzGksiKzNlBnwC9qFIfXY3eD9MAJliirQ8Vty1CLxoMLUdcsey212dw
/WQDqTrvhkEJvz6TBb6OX9FwFkq/hFRzsWBoe8M5lDh14qRdnGNyTj3XSwCOg+wwwi6fO2eMFCbp
imN1a0Ou0pEXGgn4XyHvH9r8fh5tbUEI9sJRMsNYbzGzIdABIV2Ud+tsz4hxH+vi4CPSZLdZ2lWP
nYaJmBJuQbhsTtg5n9t5/1CduW3fCTUWpaUvGLJ69X7dnHuS/LHMsqCKztL2lkbvLpqTbVgyFcsm
a+bnz8ECCGCttKqz13tBaKDeJwKRd8TbBJh/udE7wp979eMK0uELMz0RscdZwhdBDRyg09vVSJvY
0wICRQoI7s/KUpZkeKhOeJ940bW5jo80uVDh+zjbrHb7RS60hnQP+OdiJk56vuSCPGqdZVig6Mqr
nQcAVHM/6bRklftQYG3Vn4gsDzPmUjF+ZG5LQdqvsQSFJurr18W23py4psTuOmFfyy2jSk7JIEfx
2GnzAERysgMnFAX5HDuK0//j6dxNTsDhXCsUfEPdlRyNmq/bMOLAtVvIObLOnyk3akhbEyOm4jl8
0me6N/ovpal/069kNlskpk1pOh9lnse43mTSF2OKdNVknHn87viNy8y+wokyNwxMhxOUbCMcWBEK
nbm+7BOpZskmQ5mydR949wSobwG7Ws4B4RB4+qlsB3a1RuyKVxLnNU1oCvnp6BN43PdSOIaJZwbf
gjH1dduNPVyvHLhqt57fyrOgyk+gGUTTQKH/f638TWmne7Xw/8yk9gw9Rj8gBU+g2psasmz03j7O
O2Sp0Dh3tKSUprp4iHYmxy7lfX0VAjfoebLsyVJJI3R37wdAEaWBqK6mrQYsSNvZ+F5tqZNd7SfI
Wz828k6gCsOguY6uVdCHNZ8Fqra+2cI5Ta7ZkRqJ734tEBjx1srq6SbabRWcPIDS8XNyEqHJP5JU
ONT/byFCD6X4Y7FEyPQjnx+5Q+m77kNnylk/ha1IjjrAX0mPtRj2aPJRb7mld8dT8Hq+U1ggkvBK
rDsGRPVIlwlNmgsGsLCekzP332MrXuWb0SqBxa4WJlzKHC0QRNCvwL+NsE0OEq+n62J+PsrcUtMY
OKVFSQo5Wivg/VgxuIoWhCDdtR9imMsuAOs/85XFA6S/cr1ZVJw8LWIRH7vqcr4LERHxC1KVRk+M
pF2C1CP9IG/DEYdHWVWtycUEzu+LDM0ahdDwNH1CTyZMCQOwG/wR4Ay/7DlY7M/bHbe6WxxYH0gF
Kk7oezJe7AgT9AKO4npuADs/oqZWmRVPDRD4MQHNo6I1dXpurGz+4z7xAJA3PQDe4DMWfgZ0Z1R+
mthWB5CfCKfeUfcF80Awlxn1uyoNbYgpSJu7E746HNtHdjq34YeYx53fT/x9bc9MfCEyOJsFrnpJ
ozPe6WLj2QmiMlvQtn6OxrT+0jFx6b0TLBlsDcVwXqhoKbEjyAHIDHefRA9Qd5xUfAGqPUcv3YPK
rauxii8r++sMP73E+2zTFfiEZJRPCtrPyOOq5z4z2pLF1xvafH46Q631QUAjhJoqmTfLuu/h+xKi
jWlCJtMud8HX2w+uCS6F/whPI1ewxvf0ldXhrzBWF6GYJPm6b/jkqW01xZgXD4fxY9MSqKyb/N8C
AgHg0yi8ESWaWWhd+h6gDCpojUEP8sfsaMunVLBRU3oepbg71MWud8Rdte+Q4F5OLxQm4A7waaYs
ajvBUJTzvsg0NpzcD5y0R5BVlwkiUxK2g7XyO0z5Kr6zqpbLwCL32X4W5qQpsDf/VNt3sTZT8XIB
Wc5JNFHxkpfWJ8eCrQvpkph5/tWiOKkQrars20rzHENYx/e3cQrb33+pVfMILtklCPt/AzRGr5fy
9gEi3sIsuaf4bQxuXmEn/d5XA5nYF0s5xzXS1wxEJ058y/QTyjxnrGybihAnShwGElUMvsiGwTgt
tmmFRpM626qbqoOO4vkaDjhSZspPMEReYQiyy4214I8neXJjP+WkpsN79Ps+WYW/J2/s+MgrTepG
K/YJGP/h3ApSRUlAK7sIuDuIk0y4T/3I+ht78g7rSKHUVoFHtimzXUwQ41z4KCDuv3WqW6IAFuua
X941Bu3OD0SmjT/w9Q5Aamc0PpKf6+eNOiuSuItusqyoOurEg6ckmPc43gNDlJkCF1fMdH8rACw8
263RnprrnLP3eo0OOztbYDW70UbmAax8cCqhMx66NZ4uWsLLN8Oof7TzZeRRvqh7Z43XS7Y/k+NY
OARp0HL+eYU88fiDAuE/J0Ji6pGjf+bPmBRbISxS2qb83S9YagtuWT3/Iduclds8flJP7o32aTD8
6imUO0INRMLAYGToFnJMejuq1F/afZKPpuF6+7m2K+vnCj/E+OV+U7jTn4UPkRQkHEXZjP+cCK9s
9YdqRx7tso9Z3LnufzpUdEDv27mm+/3KkVHNqecxTZX/SFzUpLO4N1YYIEPuQPuqFDfAtaU2rdG6
9kLx6wbVcOaU/axy16F+SlC7OwzPLGPLlODH8pD4ltW/GBoOJWS7+pBqOwawWUyTxHP86jW6wJA8
SwO9peJICdnLMazw/LfdoJitzjslbF6hOOKjSP461BWHmyaCG57fzgl3sQFt8bvGomX+wkuqm/UV
uWHVvW6eJm8hH8KfQ6U1WSD6CbY3NSkh7ZcpR9YvjkUuI/zZ0bfiYAbKLkUaX5VV3/HGWdeC/sD5
hFcgYhZzdIjgWgCjL5tqAldxm9s+HNtN5V9FbGtzGIMdqrBJJSI28qnoY+sWpKeWSBrS6x1Ojt1s
H9yi/UhHOC57g4J7n6LQwqt69KtVRW6j7bneTOnRazim9EFSyu1DyqiDeObISmixbpHsjO2RhkvQ
B2qPyKBXNArk/KJnYXqqOnLCemp6fIbdO6e6HzswvojoISqGhnDxzBB0GfDeqHvW3M6TPMHJNpEU
tYq6ApQxqbuEWdwwFYT2dssTDA2EPRKm5+fqXObHNywsD1L2XeheyRRrMx01P5KXdj6WbaR57BRk
8ndLi25bFHzTxMS9ltw4rXfKiveu4GKEnZacdMfUfDXAYMe+EqTsOzIjIiizFcQAyK0kiIHJ5zoB
zc9qQt59Yfl8QlaWOlkJhRUbgkjvz66nIzVvTMYfIedDfsJ+BSq/wKEBUeovqbM2uSu6OmIs4O3r
t2WGfMBqyUfXpolfb2+dndODI1y97D1+CCMdvVIlW/9DxAfIQ/RRLNI9kWy/2sUlG9D85+1CytCl
mF5SuP4m9tb7QPh6+P+anWhL3OXQyVl6rk7Vg3XQNwUbSH125M+f1SbIu8JDeUsV+iUGi6fBbhzb
GgtkoL7owTTUMTD4SWugHAdYR+j5Op/ycBhzQ7mH8xmA7TE5jLp61942j19ciMgpy+ZIzd9CPWIS
21VjSTutNRN30JW0Q1EgXRd0NRtJayX0lKP6GNIlhPhUVJ7rqXIVw3Z40lqP/igC3LWpjF8ESTGB
nb11JV5qc9Ra96h6Hl4TALJI6NAVs8wVkNKtWdcvO448IOPLECh0WvfPBE+01dps9gzrjYmnyYus
TeXhXmSwF1RiRYF4XB2Lgeuoq3gxZTC6OUa+MuU2QOz3Rhkn6ibr/mMZ4t60zSSYbhbPLuaizzmg
0YkWEhZA5NiSpMSxfVrTgOWgpmI08l2SCX1X3ano5b0fUEV8nwDVaSGaqdT8xhtOoyg7CAj4tpzi
XbBUEYio0UToaPv4cPRkQfZXfwtbj0XFV+cemoyzLJxxx9aNXA4OmEMxZrdIh0l+HW6R+Ht3jUYU
vI1iMfQ+clfk+KXcVUpUkfRz8d/Uaoy4IEpJF9ZPdShbfrZPrq7hX8kJ9IrujNGnMB+PdNllgWH3
BxOK6LIt++gPn2eHOr8aZNbqj0kuVgOKTv/yNYDfBx8Ml2+yffRu66kvydFX9ZCB5FDReqIHdkda
MgtL/RWRgaqwx8E79qUd7QegZ3+I3cmS/utvzEAy8IveN+wOtnxrvG/sfx34l6njf48OlwPh04u+
IQstOwp0alT5AtW+lGKr3U+kcUO7Uf3TZNNR7MtMfKVh91SIKz/9TZTPyLCmfZtu6sT5m+yXUuYt
VtPyU+p7NiEX/g1z8U83gI+8CJHsEQW139UpIM28ms/YAO0eMOyzyuIo79H1khYOlBUFAqE6KtL+
1PHVxfCpG2fEveH14N+QtNynv0okzUcWDGYG7I2eIuS/JmvAvWE54+enHN30LH38L3cTH86JLOKh
1vTR0DuPxqiEGESJ0rn6JXyrwLTCSj1ErCwMZUfDfbN8Os9g84xjgs7uUCcdhAHHA/lkksK/UUW9
0PkabIcjzlCuhRJXqR4/Pt5jNxEuEWp8UAaVTMWt7LiaYIevVmAtV8wJ1iVRnr9x4q4w828yULbN
368l9OMzrfwCJdwSVUuu4SaWHICtlrEklVdralrybhRsKfgnq1O1mbJLSDG0iZmrmrBT3WoYcVWq
8uSS77O4tNhCzk76lFQPrHcnvlCEzM0+9fJtZ5MNwbeJVlF66w6/mdECWVhPiuorcIfCGrV6utKO
QmEkpd21n9H+oXluiq41Ac6WofQsDyQ8oy+bmaKu6CcmUbzjWniQCDTkj/o6/MTrec4amoQceF0h
m0V+HNJNJJNVYrGHmcigVL6hAgIAF1ClQ9sKHgTdaFjC5YtJY7OTUEbdDHLfeJslnPfP2SIQJsTc
xaHD8NAJmqfBpWcvqNZzi+fwOFXCFMJ769yihPABC6dTaYG41qIsUfXjDpzUg+LQsB5l0APu1WW6
Yq4048ipjszeX4bZuG/gY41BUbLIzM7Jd39xARyXV7cMaxg4aW4XtCeEGqknKGTC1z9rcgaYmxBx
fzY2ZrIVdfBNfl8UzHJHN6tAbSLwQuAEmWXORn4XaWeycStslhYqesAF6XnFeS6udYh/PcDiCm3f
LwWeuCIkLfGwx9WBpy7m0ZC8qQaRPlDSxxWEDWpv20+IRKAhabKY1DCpK8zV4Qz2m0KgOLlYOkHP
2htwJ2d8dMnCB6vze0MSmKybeAMzUaWVtotmaJcCo1w4jZLHA8chhTvGTFBw8e/BY+GLUKmsHtKK
jypQ5YJ/DwQiJwh+FxKeYslNMsrG6lHQ5IEE9iz27tIO+SrmVaFIerb43AT6KcDCvZXARVU/b5Z/
Y2JBdIFUSFFcT4Mc9wHlq9oeNPW1JCJqanjQKAqVTwtMr7QEcOrThB3y1OVhQsWV6CiVMZIYrhXo
fdztEJpysWtUhC1gKx0zqO6i2/ZR2tBWOroZXoScixy+iv5MpCmM12bwUlQAUiX3e38y9wINZcRz
kW08+QjxH/JFf3ZGl9rCmnVukKq+w5vD28+DPPLyitX+iIdX+gPCmTxJtZ0tdTIqaU0vBIjmcZQ5
gXuyhHcYxpxoNUM0bQ2ym5sxZStJaCtaaVNyYePPU1hfzm1MJna2fLD8bUNccXLd6Z8qNrhpKPYw
k3NerFnJkCeoANPpmdHFWY5Xt2wOY5QDzCA6KYd2WmS3vQlVLWrKDnAocH4GmmuC9/j0cAQbkc5M
+06/WDxSqfheduBa09D4muPXYTQLtGRY/gXCsPYxcvt5LEd59pyur8vhrhjb1MKqasGmFFov+O01
4mHlGfTqniVfIUl8fO3Afx/AQtN1YIxL5kUdqxWXnV9yrPcTjArDGL4jpZFRCQAurn0cu8t/nH0r
9nA6IGixAMxSKMTHovbr78tIZd6/KUz+JqaCw2NOff3zCTfmHYjn+iFml8zL+/Y3Pyfh9nrGlRYI
yeIxmXZfooWmL8SpVkG3vNV5KmWkQcD2gsIegv6UZsvMGaPrH2GVlBFcj4Runij7QDu++MmVz7SW
iiwzkNUfWTuhfLDrejlj4K7kYfgXLdVjeQyfuUwX6uca7QCTIzpVky70rKW68XPo1DQD2y36KApE
wmmI/H2E4U8wVC9BESOjltQuMLEkAkba1OpmtVrbDIqdjt6BPpl2IfKhUOOISq03cQg6aVsiIhf3
PdqZ2tnEwARdId1432uA2a6huGiPuQ17RoAO/HUSmZKu8TwNlyUPtOATgIbeaJNsSUEu2E4qmIfM
TTMmYhLrQh/d3GU2cMkVkfDQa/eCV83NuhTWi1W0S+WSXczxOHJ3ggVMyzJNo+c9dPTZJIV7nEco
qBJHUYrwXZABZrm1EmiUPdeCH414fSClXembZ0TZreuwDDlVk8CylZFEnbccY208mjmf+T042UNj
B/O5Wvw9KS8bPxbYg0x1WRCnF1fv2nhQYmgNOiyagRjVCrGOuD+FiJw4C+oSwwiFC9SxksxiYtrN
MN45aoF61/Tytmj2VEDOaxyYqVmvf8nPXX9Ycj/0hm0sQce5QdAfbhoocs5h+TSw+Ki1XjezSWVQ
UkDV62NMfEEY3JInnIBzOWhSbNgl7N2aQYLqHkkfV/qOeIiCHcs/SNc6zUjtTobZ0qHahpkvCqjk
nd0AA0icswsh5h852tRZxVowZ4PLzRDk+nwR3Wc4sBtiI61l6yahj/XRR/UwWHEksJRVkwGWVgef
8FSu1elLltZy6p9YNZDsSPMfJfMxgcVf1OZhqC/+YetVpspPsEFriskc+HZ9wWcrymlWS2Qx5FLd
5WP1IsR8UaOezhrsEsvsGLHKsDF8ho85Oy7pz8vxgIm5oiTtt+JrWuC7O93xItxaCBf4xUU/VYJS
ybZ86JgGxXSv4zs2mk1N+BPge1g95TCZC0GCOpvPFf6J0jyS6c7qI8LoSPBgsBvp2M66DVCIQOOX
veEDksLYbiNLikUzODsI9lXM8Wc7vL5B4I2VUFkpAL4p+vfrKx7iNHw4xzPz1QLwU5KtG59Rr9QH
Uj2yaMOILcb3riZJ2KEmjL5O92M7YFcimjkqphDsuKio0KmcZHvFIc5w5ANcrxN/GNOIU9J/PrEY
7Def2PVQnYEfMYudarHMvrevkdmYDS9t9ULAFjLtmL8/uxDamLC0Y+vJusjJve+Wtd6w6lMKue2z
NaFcLAeywQmV4dp4ZRFrVQk0H7FToRHrZDBmp6IBu2MJX6dVzp36q6cTzEu/69E9CBMT6oOR0s+s
lEO1WN/wl0mhtoFCQnWMGiCirgcZUXbwieaZswm2gqN/0BlITelyEQUoNnv3MhJojqO3SGo/fDcG
mFkPUaZXpgaa/f0Iyh0FND60SXS6CMIZY7xnJPqNkweOORisZiM7BMfNY/QIzhJHWjecVtuCWG2o
X3UgaUiX1CFGO+l2/2t0jxkRAXg1wNgqLiwTqI3wLAgx0CrW/fDHabXuKl+vkgq5Gg9lSF71VZZt
/SnF2pc3BM4uZpYsUIAS1I85WltC3bOeSQaBHRJC7NEZr2Vw7Fy5794SMbm7Tfd/bETo3gPtFSXd
KDghqcIgwtmeTZNh9bKN+aEb9fnx5fDK3nqE7o7fqaUv2OCWd5n0jAv+wXqT0uJGS/kvXWTtD3LV
byXBiavFhnhm/40KWmSATA6y6+006IZ8ohXJtztk/pyb6ET7N+MWCNn5m/g+r3wLFfmlhkVSKE2Q
SSxpU+bR+EQPQapw9ZRGNSzf+PuUWLpp+gKWIDWkoU3/TkXTERZr4Pqtz37t55TEiFAPyLykW5Kz
V2UZaYfdi8L54aa7TZY4c55WMtLRP4ViwF+x0pn3tPBWDEW3xbqmp8sLWJWJ/1bzAiZG3Zz7tXJU
nrC4LT2eImDqoyYYpYLX0kVRtYKsXE5UOxaPSwn95pg4c94INZGfG0o7JQqFk4l3W6Vj29B+iyf0
GsYbwBXLBRNr6jg28wuyIuw+Tsaa9yyAvX/v4l5KbL+sRgO0jNhkG+iYjKXN+vBNcbS1c8adheKR
STfRvfhIZx/GFDrF6nZJpR8OH8HsWbcsb3c7KGpMggKHdanqHwBOfvXmWad6p+VJ+N4Gwxa4HbnO
UICeP6y96xZTiV7u2KttfpF+/mGFfcbSwbyHE4y7iflbzvslETqw5HjLBM2LBqHvedpT84wbZsim
XoZoAMkYnPsr7G67VUar5KnHFdr26/9vZV6TeKKpIZi8bpG4XrTELGVOKkZSpumsgxTNsXzL1N6r
9yydxwYgRDooO13sdF+BqFBo0Uu2ZNO9BGYJH1osahOu1uLvLYMDZ6AhZU90SsvUWdgRU0aGGX31
52RpdGbEOnQxBwuIpn3z8PszMVjeaNE+H2CsWCR32oxns5oylnd9O5CoKEAliGuDDHZuLy+KnBdY
o8qACYWwzZSrG/oYK/dnuR50gZf+pISIJ2yJt5p7QeqA/XVZRmF2DiXVycLKmSaS5xfusROf1yyB
sUSXJ2sLUI21VbQuvIiKg2vExXxgTWxwDjMkRLGYV0xIYNVR3y8YWTXcOw35p9LqbeLV9XeDR1db
hHxIE0wuwaOEIj5Vadb/wAEqYBVplRhXyRr5rY5NlxhTgYWjG6H3r3Ht6fn+qDIRoLdoOwYkdiRC
Os65UI9vznS0jYBR3eAGAz1fF6JcHTDrD0qdC+H1fxSyZzPhAPmELoiNgNPAN0W39kl45OZAKXMG
pCEQbIboOiL7zsjuUXKg6zG4Nu86V3jH6mTYkHrKvj1nAiRmq9ILsJGHhMLhTifw23cUciZYb8d7
xrzQW17HunKh/7+uKbpu1m7wOFxL7xoSw2pVAseFrdJp/ibBGG2e1jj5qnCu9HKPDW6HCQIk/Y44
LYD7Hhq16pSBSqpNoomFKPXmVJ80bdsJBM4t/C+q/zIKarUbA/Ts9Y4DGoyRNPwVrcY3R7Fx4b09
FYX+va5zWZ/bJJtz5owFzSSKDaNW/5+eaAGE+RGjJtasNJb3PBReZOX3qH68St5R9vLNuscCOC+w
bFjZ3isWuOaKj1m/ZJaLejOGq8Adc7k/NuzFHbw2g2T7qyiJoFr3zCioUnPryUo7Ve1u7Kt5h1qC
iCRum8GdwXZfik3G6d6eLvSAwzbCNubCzojL/BxLjKqZgEiUcxP+i+T/sinPwkOYjDzj4YbMpEoI
TfIifbYsCVRHWMUKaxOFNqX+/Ux3PamSkYp0FQmObuz7q+vpzpnBp8AEzx54GCrkygHTc3NRpEJQ
GwG0+IuxTM4x8pF2xt9QRMUVf/LzVMREG64zhh6qgpMkFrrrOY6xNM3wp+CwalrHy36oH5egOwge
zYytimByL8KoNeroK7zaXFfCNtBEbpzESEFKvT3ai2j2CiZqCQAmOoqQn5BujRho0g0czv7Ry7bU
7/3Dcj674i163wkmRSRtUvm1Y5H8Rc9XI3yiWe7bvG+v+u4pfPBph2NtvvYJwGg/Vqxr9fZuoRN/
nOHRvaNa+yd65NwBHB9iIxPgpgQQVFm9YyFS3z690vsVGhChAEcWDXGcrT0yIZKFi4kurJ007+Iq
Xf6KK1s6YrCvNQ1D2IlDvuXF2ej+bd8LtxBZLn9iGmAhaaPnV/deYN4T26aLmxo/VUAclJxon3B2
LF5JuW2VXy/Ouvn1zZ3bH4T7bnOTD/YWRNR6JpIhXe+rhMLp/7o+Z6GMrCgkWytM6id6NbMZc9m7
r5nv+lrOB9dK3U3yFSRh06XvgvewDtnnLQLjALzehjLUtA709wLn/b5paBEqQUOLaMNlIuO8d50Y
g7IIRgLY+Mc1C/7ahIottpBDVqyDLkpk1T/QYILx2uhq0K9yHbvgsrXrUreUNjGhdGpiTPnbCk4L
SwInOPc1VbqT99kMoGYaqpdMwLoAB9vh+6/Dm6+7d23xzOz1oaT6W4WFeDYLhOzCAg4C732bXhKt
8znvtppvOUDA0tdY4ZWgSV5FUomtgNs4gsy222zfc2jyI1FN3Mjr9GhkV0hQNXlIw2x3OoTrRzMk
vvyTqg4yKl0zXjSQQl5AX76k17NqgJKhb3Z/AwPcZPy5bnU/vhd45/k5cXFP2jXCAuZ4nKPIYytl
X2uq0HBm2PCp3kEnXcvvJFLUSnjQ56I2ro0bHUdt0r4nRyru+8hLK8583jVuOlWy9mHbMJL9F1et
LskfaYiJ1CMScyV4MiculUw3GueaQCa8UHzc2UNLch8mJVSUjb1f0jBHzjjgq4eRBhyNGqEvr14o
V5oQ2ytQfsIDtImdk05VPoD+U5t/CeBnK3xfEPu0NosQwBg6MqUt+EbVWkCsCScB76Dy7dX5TVcU
L4UK4smK9did45ZK/yL8BpeUkomJiDYVnNpOZzZ2JmRp0RcfDRqbp3C05xLR7e3CFPYueYLyPkQZ
PG7GO3858TT3g71xn6FNq1TojSMeTcXaAHKLmV9Cox/Rz1OC7YMoi6fFv8ih07UG1U4waZ/4OY6b
mmxpIQzWBwuOfnp17MClPpoXIxpLWg4SNXk/MvgrwRF70TGs8qJbHh3B+GeI1jthx06aXbARWXCP
S4WTH+G2VcgjiyKjeSZf5xd/3tlp8hsGAwuxBcQzCc76o+KCMsYeVt3hcZPyTi3q70+ACyaOSzZp
FwURUGs9ti3HNRafu2Tmn9MxvTJjDrqrjXK8iDcvyi930/moOblycyCDCPkpD46dleYN7FEs54t4
HlGtVFdxEgjbNIOM4YSUiJO87H1nw94rPIF2EWcqwFrH4amdH8/0WLt7++tnbPCNVAgNwlkWn/Ab
vMfGtDWxvNrqPSjzVW2Ya8CQytlHWACild9RZxGlYhBsZTFXIIOHpUSD0Gu6jEvHJ63SsoaU7G7D
UWJx1vkEEt4J6X5I92ERqOI2PT4qfcZ1BvJT3PBswNy4Mu4VxHdHgBWige3efFt87JsT/mKMOBGG
K45F/7LcbRowYv1B34PKBBSAoVPLt1gN5AhNkrfKIEHbJU/L9uFSFd6qchxCSfWZ2wymRoXpiAfy
ITJKbYO/lPqTixiTq2JZ7B6KTE+/0HSDgRi7kxq/QVZ05Cl1uPOJIqvLroVAaURdtsXgGdxH+RMJ
3aRZlxUB93+6pwF4vLGGhHs1ny/RnMA/7xkMVnlg88aFavPn9k7fWk3gf3fHeM2w1nE2ngofqJLg
UsL/hfmr82MvH8f1MbQB/bI5eqOBQsveE8nD5/Gon/yhRfD5VQyX1Pl0stIVslTVcf3GNV16QijX
g9JbC5d/MWC8jJE5CC56XF0tyDYWvVTCleIeVb5fSOx7MLcA+g8ACTTffeh+kC2bf+tW8OrO3ePp
4vVLqTS3Oza2rHQbG+MQ2ADQPeJXVrdSKfJ6vWVNGEGZXvWV5GfhkF7HAheiyhZA0NTXpA9d1Rsr
WAL3oKUsNdKIpMjyCt0vZ2nFuxNomF1f9isVv7VqTVP0MJRdXZ62XjT3wWyuO7P2C3H/dXfVbDRi
wO089mcpbxIilOH2NVUHlJre0++EM+SCmAwC3XUcrlyreF4urzh/K1KVosMwMLewrU3Uy5YwO7OX
AuFhbjVP3toDajAuEmwoJPaDBZvshFeex8rElZCf+aU2SbzZvKVVWs7F6QrzZe0YwlUM8Np/ZmYN
xBUKDm3rRktTRhYx1OWWc6fWf42iKOlUy748dq810xH5f+xt2ne2NQ4AonNkruUrcTQ71l+tQNET
IRab06Qsm0vYTFaXzEjlfYMajS9PT1Gg/S5Ealea0lAP2Bsrp97mGIMDGI4PqTa0ZJW8PAbzNdzh
9lp6OSNetl5qc8c0OmCAytVDk2Zmqr3ZBt6uIs9DVt3hoUQdX0ZwEUbH6osqYrshL2iS01IJGvMJ
SB3TJRu0GWiO1ydg34oxFDw9VP7u9ETsCBHuDNCBPkSrJqE9wIaYRd5PX8+VvVE+OPcL6V4TIM2V
5Z8R040aEvWP7ymBUzYq3KYiEtIUq0N7CNVq2wm70kZGG4cfzuzJNLmG3vLs55TLxyFz+yIa7QTm
HaTHR5hHZikqDex/KMY2xnfoCX4ekuB7LockwUdVrR1JQA9Yz8idq44+1OWtgBObhPR/uqca2VLw
LaTog0MI3YPQ8a6PzL0s8q4zhqPi7J4zkxGvuU3XgTgt8PXditLy1OFf23h1JJemtPmQVCXc0YAB
+TVWaYuJheG1e1imX52aiXUros20XFTeUs/XDYweDan9L5IeQ4zpBY7dWA+kGdM5T/nHr4gMzSsn
1jqp8pbiCwdhJ715iLhdLCOYNQpayN61PyKeXmtMRRNPXSkj+Gn7gz2EvGjt3F4UC+c2xXkLG4EU
ZSl6LXKLKzg/K29FnN2Cj3tdcvZyLBVV64ukM1/U7p7mw+NWBbhQ2fP4drz3AIuqlviXGZYjY01N
AoeOwejDqW4iO7SUX3kvdnlkz2YS1iZX/KbdNvrLwSFJs4mrEBde8p5uToK+wT1/XOC8yuZSDRp/
XbSsmz1HQ2M7UNJcvXwah22Ys6ucJ4sRiKcihn2rnlmdkzYwF+QDaA61NHFv9AdCfsMEiMqsUnru
PZiSVcKEx65Xhjmx5Xz8EAkTODl6mrZXm07JqXOTIQxhIBqhDQJU2LfpVbtl8pN6iBIV2VoVbsVg
Xc+28p3BP+vV4aq6xELWYlV509vyvefWdWZ2FB951b3b2s7+NR73mxOSO4lUhqWse2gRpmpClon1
iek5lNvNW+ZvfXH0jB4cRVdH1x+rclLEy6z7hzluA2Z80+Kcw6s7DaWhpxWXq6sZ/BYhtcz4YwtW
XwCqXqLFPYYvNXP7d9+Kod5wVp1m1fRcSaX6sDN+W+Rc+UZsxXiOuUaRlq63lDUBwEUTuPIpmSBH
y04uP5SDpk3NTT2/5obioVHuBNykUAFYd41Lh2rUapzhi/cEzrJIKQU4wFeBYBZJyv0KVJ01PPqg
RWDDLj8VvYfeMED5icSE5U/hiQxW9b0LCukcrg8ZRuiWoHJyOoaSSunw+reHZWi7yAFmgSw/BiVA
OqmkNmIQxqnM7P6XVSv87SpQuBPRDxgqL1BZ9+ZB3Z4PvfEDdl8Y1bFmAqcS9X0livuJKZzulDzK
cvOYNnfsO8HrPjKXKbM/4A4HblSHHukKHMjCEkyEJWO1R1cA63v+gMTutHaX+Yrn/zo2qQNrGz2N
5k0E4K1Mp2lzU+w3Uz0XQ/Dxmv9gD8NZ2kQs71KV9KsCMai1SPky5I0DJ9xFI3V0oHvo5XW6nHMm
3m9jkT0jJNhrQyKiJezG4wBmjqYY1qHRMIL2ANyDtzyeJ6L34dvk3ysoExK/8rqAI3q83WMCl7re
QwqJPYFBnbKVw96VFSPH+Y0Mqxmwx3IV2tV98mLp1auVQ5PFW7xv0djK6wtdk+RCauyTdNw3HjYY
ci/8mYR7O2xHBMY0hVVmlk+LYY60h8CWfgxvrF93vH1XHM2NTS5qQx1EtTIRn7dSCg1vPQNQQrAd
r0AU7qBkY/BVK7q3ywBBNUuDpsfwgDO/FVWn+oQiHLPHkrSmOwt+FOFXfzNhqSQ9cGiJ5rrXweXX
bvWgBehMtQ5+RWGRNP6MLiHgmnXm+66Osto314Affgq8ioWKSKaxnTAlsM3Hp6xQiAa5/qqzuN49
o7eW7NezCnHlMVg8oVMwOFhYwMvvjvCk/gb7hlJyV9kRJrEqUAqC7ptmUQoq4fzkFA3K8y0/wE1h
yTOHqXMWgFf0P3YTfMtwtiRYLiy4hWYaO7NezAblKKZiMvy1zcLm4MmZrStl2ilKmOhCoevzu2+p
mu1gjDgq9f6YEf6q0s6qXagNEFWpB0ksHQMk4YdyLPeOZ2IhbpRSnJn3EexxQD6MYu9/T+JBIzPR
tpDGuqZsTHl5ejMza+EB5RRpC+MYgVfoUcFxDTepuA5YUs6CJY0vnYSlwfAHaQ4BCaNe+dDzquZt
HN9cdLLazpXwZlte34rRF6m32nyKnB4rpT+Rsr8VpkISfkE1PX5okESc+T2p0Vtk/ZE/AJmSzq9b
Bv9Qd7wCT8sTNbj3Fa0ZfqyEP0PAVrhihVEVEDfy5ViO9aTgbDGpZYhxfDxC1qEnuxmGkBISY5ip
Lxvy1P7UYwQgzRoB4g4zkqxQkP8ObR67X3ZOV+Y+iVHyNxh6wtru9jAqtRpzMXn1u8g/rwZ/EcAw
TmPz6Oiure/tyuBb19H624Pik9qBZsC77U4KPWc3si8VB1tOpk7Y7xfRY8tdNHC//qxVFtTU8/e2
CmXemxaMFc5gmuJIkQqXAoRCVq6IpbEMcIsXZpbuee2OUgYoHHrQq2dM/9bAHu2GsvPBp+Fz5thg
JZ4eNkNrc8KOSUTLFw7ch3cwr8iIrn5kj82ISp837g/ph4c5Vue3JbbqfH5ePO/SSonf5WWM63pX
OGxNM/gmmTkzB/Kjb8c9DBNx7fbeD1MalnWiSk6wjhOpMIlB/LGarIJ8wzXmn9Rhq/+4g4ANVNHe
HtTGDo0ZwkgPzShfeSGVd8ztoA4Ja7lNuZ4B9TJY3fRJwZ+9H/BcGZlgMzvjPcuWcfApM4fpEZXk
SHQsZdpUaNbVUiksQYTVPMmT0+Fi1RB+8p8D83Xo8fZJq8I1tWyrKRpCKoz9pStyupfkfYP2+b5I
PZznXQRbmuJJOKBO6EljXm1hK6QbeOCQYZPzIPyZDiT0bz34wq6AEcTVs4y9J7vLSf/mC6SBNo1R
J82GdLQcojc5EW/tLj+85kP3jfcqBGb00YJRjtspf5pzlhBXarRJv9J1H6sz7ZDZ2TkfhR4oaHka
hJFaBlpxtPh3iesOxXUKD9Mf1m0nToZ5WaMphF1t79m0ez1sFKin1PNh7WgwWhpDErauI+wtKYt4
tyPOrT/tW6QsQDL9IjTTr7bLzPGQZeoiza6VoyW5KqIkVvVs+KIVrZYRVWA0cH/zyqlnTmNdLX/z
Y5ihecYEqJ9mKaD8bErJ4aY+rxp5jTeQYQYJn7hlRQF7bUQHa/WIFrRyTfy85tnxnBlRhwm3YehS
wbfjfqFJMWCSpR/i06z7hAjpwGj++TutXLpMj3nM5/EDElWlkWaLALsDnGhtwIgPX4Y7FLykOJsw
8ve+9WKjcVBdJJW6Fum5b3h0A9jsUHm1wQ08P9RBCxyJYs8KbIBbcgvgLkrI2zreqTZzU0C4Shyx
GxFWCksNYjc7s17/S8LzLRpWtY16NSULL1eeXuXq5e/ipQgRk3AMZ+6jnRTKY4cnaRf78jmJeqKr
j068EETAGouVPEEz4zl7g61JaYTy6pNfm7sYmuiY1Hky5oa6bY55qu6kc8ZHw4mz9LFWmFfkv0fJ
44ARvDr6XMX4w3pVQP+BmGbC45aPBpZLG9Sr8Mf1B+UzyVmAX3b8Efx9ruSNf2tUVxFwtJlpzWkU
zUF73rdw0b2EnPNFtDrS8D1WCh4NPgnbQP7D1xLcaAHI6dHi2Y0ag83zWrHKezNiM2IEn1SIDWTl
aAGQR3m0q8NKfn7P6LhiPT5cXrulEuzTtt8lgzti6feDjtKlsw3glhjXkUy/fBVzk/YZ47QnvkX8
O6kdR2EikEyP8ZVJGzX5p7cwXqV2pzr4yoSBUVDsNgFs0NWtNoiSbxV/k7Y0PhRKLFMIvb3x6lwh
9rCsFQm2p9xfpqmyyBz4OoOspPE1nKbBVmwpdMxs3Jeu8VKPQxymz8vATf4Yun6k128dE+js64he
AsPJpUodzPLvPBGEHP2ceDJBcjx7CpYny85w3Tz2/+QMHCeDttPtpkn+em7zmiO/35bvOmC5KVFq
t4bR/3Y9FQ7kvPXGApwuOpCNm+y/zW/sYN3CKwejfhgTWCGe4xi7LT51qknPjfTPGWvm/JrKOCfB
klanY36uMsx3IbkZhPQ1sN3IDOX5DJ2ZVmhOq/2IE8N9alk4k4i5/GGiaNYXis4GyLM3DAaDntbM
6YcsW8fiTpzGPnFu8LxCj9Lkv6KTSZL50uzsIxCsDttdzGamQgZyzWVugEQlN5078MeS1XRGwIxL
vsYQ6/7BhCcmjT7RR4bOwAsfGJ8moiq5uFKDxLT7o+B84Y7T3n8m8wtBZcgEAV5T6wRHQjUJKKPr
WplKcnaJcGu4wqjVtGuOtaSy1tqsg3i0IV7C7aBqrBysJ0lE/IufrVj+SLcs8/qKviAgnMG/qA2H
Cyjr7jCL7dodwN6zzLAAJlMKULVGkvI2xsIsTP2Ji/xU9Po9WABklhE4rb3wC4/NXnDsERbJgXQD
tCNxDGlQKQyHkg6tOJPJsOnU7MGZ4u3VecIDxBfzLISEEi1h4Ry23Eza9WCRHaM//pwjoD5E0I9F
L1EvSSEWofDVNDdmHm3PuB2xwPC1UXK8S6+eFV0MTMCmycUdvycgg7fkRQi550e4kcRkIW+Dwh6F
1WO/9SIlM+WssePk4jQznl5cVaPN67LVl/dq75nLQ0qsne1I2UMznGc5E/yRcnZsAk+JarU0Il68
VPTYCspyJBGDmWqWrdGSlLf+m0mGvMCwfryOJIJKNs8rLvmEc98DIljVrY0MGai6lwkPhiF4e8Jo
4SH7n1pKGaFiFdASWU8JtQJ8JDwb+Q+iTG6BcK99jowPef3NgjsT7aUAMGWyWeS3z6ibCPsxdemF
3L9McWmtTLxyTQ6YdYcAjBo3S+mBiNU7yQgVRwSatXrJjuhpKpDXtKBoQyIahijcz2iaX2gU6seS
yeSIAEyF3l2MhuL3JBzots3MS9DSVIiOcpBwBCg2mmt3APeomQAWo4iorcwJnw3ndJta3kdNwXdX
ygN431sVehKVW1DFgH4qOzfNngyEXbOfJKalNmXnM1xongVHjMJZgGCHerOm7xM5v+yFy+PDR0Ed
7DzoenExDX+DeSmqXaI31kCMr8CxDYPcFxcj8M/IkQqdLg2noGLJ80EGt1EGtYFp0QL0vaaFByeU
FBJSZ4/w0ffIjD8MLyb98Jw0Q63qnw3SZnF4Ca7n9BWs4jmCn0p6CiEmGN/i2eDmuqcGY3R2oTQ/
eOnj2thOzGnSNAF64jsuSYsJ6OrIliCzwEp2RRS66/z3MVvOnIqNd+eLFmG2aH30poS9jOQXEIL5
MMPNFXW6rNPaYLtrRggWMhviYnXJfsW26ugfHGlyWhDko9x6DvyYLYlO3Slr8aiXhOe0H4jZ3wCh
nDQshLANfURVdXea/UeLlIQbAmj/4/hB09HPBGUtlVfmq4L27zi64gyVDwM19Tcz8QH8+HXHcb2W
gKfmpEBS0EvyAFoIMhwLiWYbv1ULuMYeVWryXUD2lSnEUxIh1T3k8+zcs4DkmOSuA6bCYcKLq2gy
03BKnZThIU5WRWZO1ckfXfI+dXYjWzY9zbNlQJKXFXFBs+oVbKi9+zuIK2BEK6XOu5SQey1xjY8Q
NW7UPt8NBhRwWWChZdv1xAnlD+gshFnnPhVu/SzPhE33c06kXKdH7R+4QMcsAYuai07Fzhk/l+EA
YXOjPb1KAPEU5EDBMvnDCyBoT/ehNDGlkGhxVS+e4EDi7AA0RkMUyGgzuVPdbMBlsFdArkaqm2jO
By4LrGitiXiH9fjdc9PpL2Oqn+AtG5eDubFUUO9Fyy2dPc3tk4POJDBCszJN2+uwtzTxdUeXdH6H
nZLq7XiEeUwZpyAs1S0L4M+nNkuEusKHqyP33yiBiG4Vz0G1dWwZ5klsGpS1tLzRvLKGguUWUKEl
xFgTAfjA+a24FakKNFQ+1eQnh3ez7flh5RNb7bXLmGVP9TFg7dD8l3g5lqAndsrUzimHBm2NTDqo
83RZbNKN7269f7vkNAc43mXCsM6B2QMSQSprogR73OxJno4Zbfjn63SX1q5R82GVIUiASk4eRfrb
eqJx4O3zDCmAHk9gYMfaSHEQO2o1YlMH/uhDNbJ/jQQyL7MPoVMmaJJ8chUaRbFPzfJfj4/i6DmZ
yt2qEvYj/GL7ZpmEErPLw8zGGMstnTi6U4+GVup3ftFU1SUHXmQj1XH9UL6ELRsgfvIQDoJhbcVW
jSBc3qNeHEMxMyprk29reITksSu6sMcnW0nmSnIizCjeuSiyBVPoSLZTY6DdHBZsuLelihrycxAk
V7H8K/WXvsoCs05K7eOoQD6iPJMDEnT5VXzXYvxfCLQu7ACsuJuvW+E/PeLGKMJY7NeS7sploXSi
FplS3vGMZRb0s55doyss+Fs20DnfPDSWGAY3PywMhrysUS1GL750fLHzz3buG+YQr4Vpm5CpdQNe
mL4jFiYxsODuPjuLFAbB5dGb1v/A0zZTaexo9RF2+atP0q1ZX9EamerbjKU7QKruEsvDlYZqXfCn
xizG3bBtQ/xQ1mlJZaOQsPO7eJZB8dq8lBUnw09GMJABGtG8D7eQR++wUvu5g556zlsH7Hcq5fT2
JY6aFPdt0Y63EO/NwUjC9hEGv/ZFYALnA52ryReUN5uzVRXzsKbZQpNEKbmqjasCQY96aVg6zvdo
m7LioYkJa3qguwZVVmm+3re+eSKNyXeLqSDnFayQr4PzQ3tDXF/x0JhQ2Lglo0w3rfr65a7lXvM5
oasm/+dSxGNgyQSIlHjgf8t27fymc6fuo9bbXaEVJVH5OEBDjFNp9ztvj3dtB8UKKjoS76RXf+dr
Jx6xJH/KkH0eIEliaKBcf7bBrnRTRJ5Yt69Kixax197b26tzEH3VIK8gWvziX6y6mP997rzENIEh
3jRBcEb8A603TuX//noKK8vtGy/YCv8TOkjqPef2haLSnZxdYIm6gXkuLmIzTI5C9TuOPXiMnALK
J808Y7F0/eayrXStXIglgV6qiQOCb1yD/EofkM9XDTsGG4ABrm6y3x4JqOuGHeHoSxMH1VnJzv4R
hLgGehV32MHBT8WyLv8hnrSfwaGs4dCdshs3keqHpO+9OmC321+4VDnGIEGdJIfkf19QcGwnQFiM
QR6TnMAbV06PZ438BDb7M3uaNl/fqLBCc4itfmCogmJ8LuDD3jW6dB+zm3ui6dtxXGl/AoXCfYgu
yoKHmSL6aMkPH4z+yu1n6mWGVWbYAhyjvj3hh/eJAc7g8FYlajWhTH6iX/e/f7sLKLySeAnRPcko
Y49MWuHalhq6Jwow120/ZrcN+jyV0lDOMy0mnlUWFOQNDDIyDmJI/Sl97PpwB7jBoLd85oUNPpst
70jNjOYUymcKvrIEn6sTDnJx9/RHgkvulqyBGUhUrEGcOEYM/coCyQiFkH89f/yEnTJBzrW8XX9B
tCDrzEHeJMV0dlwoANkj0FabYKITNwt734txYlZlYVs9sZ2vaxNUORlCPKaeQuM6bSi2ZPZSWhcI
0TeQtM8Cx44xqmmU4dFvvupDaLF4y9D7vznIeQM2HFDwr9yzuEfPTp352j/7aUlVXQWCtOHWyAKN
PlcfpR7T8FfY4e+8ly8grC4ShwQSe5t2clui7Os/RXW6OHoA/Smv8JjFwMCnshuZFZz66FHonjrK
RM/qt6600XPK3m9/e7KylNLALFyhb05rHbDzwqZ3OYIag43YRkKIyzshQKZkoBlitjNk39qNWUan
vvmgjoBehdOMf5vSE5Sa/iQJM5I0n+ahVNwqnspTgz4TgrhrsxL6UHgRV98aSRv07P56pGdn4Xro
fMknzzyCKu5S+2vd7bRXBMVq4DTMVZ0C5EhuweA1ygSwnqPaTi4nabe7a0k3FaFlqTR1qC/+PixG
BbJPpUJnaMs4c1p31euwlZnBei0ZyvTOavwwm4lhaO1lgAO76xalweHJW4U2tJBNbU8ORVXyt2H/
8iaAARbbFyEJRAwRjDlG/wDWV/lqRkqfgjSRaZrMAP4Qs6r3+FttF4ogc+LTlpZbyuSfJrLYot0B
uM7Fn2nKzTPlMXxOe0253ea/2+jqkgqv6yeMlCK+JygxYpdBrMvCESYIUhLrezoQWCPgNsYXbwNr
ml0lCX3UjHjFafpnZoth6RPk//RW3QG6v6BHAv6ziX3G1TxsQw7z4VRiVblBo8M16yfaBUBXEEN+
3zUfXJTMAla3AW7872UwbKrpZykcno/eMn3hcXQjokXTT400sAgdEfVavLZA3f8LWs7dZ10iJW7K
OaMgT4lm0/RNLLk/+evSGDX3yG97kfvRB+nhQo6/iSbeIV39h8b78I3aBkiWKYH75zQUDzEeHsGm
MskgsPW7Omf4Yxn6siPxF9cYDxc3kz2JttnKx9oRm1QXNmLy9QdhiWJDxwR35HQq+oqRJPDODTsJ
/2+cNWdjLHtUpFTFDAkJGrGQyXke1CbFTGdrMda75/rCVixX5vqgtxnRamOQWwq9HYiSYZCHt/pa
06yZUCm0qtew+kUUYi2eHoTAP0oAaeCc5Gj0Mb26IfCZMap9Xxyo8AQAINdtuCVpkUU2UIzgukwS
J93sbLuoILkVxY9JBZsRMAQEfBd1/YmpGGckC9yPSX3eDL50Hon5QoMH47kqt8HnP6lGC6RFy8ET
KCUbrx68bFxEOXMBVezYJAGxxlM/xXyR6JVudGg4+7J110FDgK47r8PXZZzm2Kt62r6Ngyn7sP9z
IpeXFV3/ObA0H+pW2AligUwGoEIMHwHik7rVRILW9vWGbS3Kb+dMmidmzcbCCKugQQnfFz9Z7/si
yAK5Y1fYrz9eBCp3HX5tqK5oSCWlr//IhMsoAqHstkIHfiEsq5AL0kzxWCI9vjcUdNVyEZwYX8Cl
vbIFTY3hnEr6qVgepETo+J4dY3dypwE5YaDNiRi1bWFIEyajmlYSGarn+jysjr8xi5o61FTjNKYj
oXO5RJh730FBPsgFI5PPUzAqxdaMHdT4dvGKQwcrz99codgrzcppddW58CSIal/88giOILH9MHfc
tAtD9XmlOgVdY+tVTLNpkaMQuVi5xKUTm3N/om15YKbHUlhsoDK0ho8Ww3cCFOiSFnoTdIqfM7Dl
KqX+SQyaUEqbuRxBQ5CTXz73wdfVJuokTm6SCPBEvV3945yAW4ByIGjwjWo+gNMhj2kkIax0VEMa
4lu0ULmbUCWjb+CuKV1Qt0g2CVIBSFmueaF6fYMLtQuzGtQGjoKoRpkIxKcn0n2j6eEAT9vhl5kl
ewmZPPENe3nzpbaQy18P+YENX87mx5tb4ToD+KJddqTHDVgYxkgWB8eFpzWw0IzGgk2UdsaXEwF8
A9vSRkamsoC3+4V+Ju1wTg9fq9w1ftdO6HO/pynoyWSm+HRi1J+OCNx+bQYxLa1ZSZ1B9u8ha5JX
21qjUlMRJYks7Zv/WhZfkUeAfgEFYnRtdsQOAOdhktvq/XJFKetU497OupQJO7luAvbmmSvNgUFU
qNeo+4IZc5kZ3dc/TA5OBpcKQqqqeGjlryoRPl4MRBUbj6OiIQmYLiEyAFXjAq9EtrC4x9ir0/YS
SOTi3jfCyYSBKOTsxTP2f4v+m6litgILISEJTVaGEvxPll99n9oTi/7LkA9BHXEMsGx7R04PDhk4
MnZzv5QT22fhEAq3aQwj1IVcqB7cSLFVkAVwTdbgPtDSlftJ0NobcZNCyTW5lLOUmRQI5RKAtTxb
ocHg/pbGqDIiNmlKR+7xr7DEW/enJ4pglsKPIjSYwp6VpCo1gSttsiQXACftgIvo6AIbFvDzVG+W
ScjzcQ36Oe4sdRkE8lkj8NHZa9P7K672cRJBO05nBMnymIjZR9jCmfGBllJJRgx4pEMEhvDtgUiw
fanl8kLAtSx2kM4fWBEFSNk0DovSefY6YVl9D+r0SLahXhxCaDkxPAuhMY9Dq+WnjY41Cosx/j4n
AdJXONE8VYjjebVOIEet3xBPkbhuzDmFyaZLnSuws+B33dYWUKSCPNYsTnFZYkI3NnSM1BZnTHpK
0ZnZxzM7GDCL4DRzfSmvF8I/GkvYPkq2x7Hs9v/VVN99KLMKHsmoVUl7DldMz1X2i40xq7/TEgu9
T1YK+YKbZ/tnFeHxaZx47BHUnwRWw9e+oHKb91Zl2K9c19z/9lQMQwJ4fsstbtXYUeUgKSkdRbjx
44qWTLzT4q7y2+ZZSoqFP2We6zX6QlyCAmel7c175iVdCsGDIAXbmwh46ib0ZKbNCll/FWmkFqLG
wIafaycGW9TMIJS4Di7WgNkJQRD0Yx8nxBghGaMMAjDXOhR3Yagrs3HcUg51j101l7UsNYr25W6p
N1U+A3LbfMQsnDHth5bny45oIEwA+2OZvzr+NbLeICvFEmNFgrtHiADp374n0HVCeNixWX6mPSxR
TFymxxFC1Q727Hl/APahHJX4TbKdwkiDe40u06NKbesw96A42QqR1q+ZPRSmkaq+3QAyAWNH3LSZ
l/CEU7ALLMfOyQBJ8f0D0L82nh2VPfrpChrYFfY37aOE4XHFAST5Q1UhrVm1i/xtgZZNXsV/VDYi
533KhoBZfK9+QWkMWn4mH+v/yVYGMsNBV/1vIfIKKaYCs3xHqj92sbf40LDNcZW1n1EZ7wPuX+mc
EAg60ppcx6o3X1hnUZTRk5Aq3T/ZBTldP+Snav8Z0MH6BDK5vPrFltZSt1mQzhKRfBVVWdaGWtmf
/HLbJRPhUR7gVpfzwhOOFYCPfaipvq48tNiecIyD/l0aVSsPzBh3xwp1xjnDAxjYkRfPuudTULwa
LkTjmL5roI66RRjW5+xwOyQuBDKn7tvpMuVsmD1WXLSOlpZJhnUwCYOGajz5rBF+aiQgljFS6ZsZ
1jYDkHx8TRVb7teMdBITWcLdcLZkUhgGRkVZF4RgfcxiJek1ToekEgNfTKCTfNitJA0ATfE6JVTZ
9UmYu/NQf9G6UD/neD74z5B32AvZGez4Qob5CSLpkrLBXNoRX6h0ctsCVStSBMVvegctmAm8afY5
yUAjXkiG8/Xs0NjJ7ef9+pw5YX38jmW0ihqEZxUSdvODQYuJCNL+ToLNqXYyR9letxeIY0DvsKSP
5y0nSN80Yc4aapdTrgT82gQ/rmLWcCelcyPEImn45re/Dd4u/2Z5cLDipDX854L0rLdZp8IOs40U
4WjHlvNxB3XCooYF9MoBAq4TtGwh9cRT5ciDryp3JIsIl3uZyCby68BFjzigGHqDBu8p4UGxCYNa
NARX+b2SSQGkFUtRdATrmE45xMzFWK+I28UkHxFmyFXfww2nMYSUmoEGcQGMDMLrlsLbg7MAxeOU
AYD1U3fJep1dGv63fry7+XbhsxcOUB1TDauxoZP6K+eQD0Ax1foZWf0ChIkuauAr2D0SOKo7PeA2
0l25y4lTGcDCakxDr7VyIg3Zr6jrSxijaNgW6tGoewMQ9tV5y1Mpxf+Xrbman8BRtgB7ufP5qnjn
s+97qg2wiFkwSNhitFoTCwRpAVs2ud+TAFCTy3tAqnHba+VZQBFFaF6AwFgkOrhsR2mwCadVWyIe
Og1BWNHAKC/QKB3sY91d90KzSBgMk7XpbLdp3Qa523KxoEEqJTV6CM0g6Mw0bG7sMlyt3XgIAdzC
M8XnhRv23u5Ufro9b+qrb1mPJ0mvZP/khMCNe2b9HJnzaf7Ta/ZfL4ejyl7zl1ITIf0XA62blI63
ffbEb6KprVNnt4eW62ch9KcWn8PN7vdRvNxKtDzmOR+xgZQrIBMVZRJouXBaB3CoBuYaKPYxUps5
KIGxruv7W/0GWUcyuOgXRQCNiTbh10zXCe+N+Rd4kF4Lj/x9qDrAMEo+DKVClO/L5dkX1/L5Ibrm
LceX+DJuEgwfyPW9Z+NknAzx4BhCAkwgAjH3pgQWUgu6T3gB4U/dFgorUUrpuLFSXouSBdc/w3vG
VXOdXlnGDTVuo0hZi4sYCwWMsmNU8Or7cZO67NiRvUsCcJoedLfeQF1q1AqEsGnmgOkjd2wNVZFA
LI05aI93Zw0MHX6Wido09VcN9WgKF4OEkr3EV3rhzs77S+MNIw+xIMpIWXvBgib4T7FAV+HghNYd
+CMZp7T0dL70NmPVJNgnhEeKYVTns+rC9C3LmMMNyfzDtwyF1QNKckKELjOv2pJTvNfN3OGqer9t
/+hN117fTYEd5Gqf6r8Fud21JLLaInghaitDbq5Cr5znXXPJqM/HRg++jHwPRCZkdQZAA9vl9q06
gNo5esHQSxL3++bkyS7PicNME427lLTiz618DKISOouPdAEss0jySr+KtP/3yH5s80W5bcrEslrC
1Jd0RM9w9LVqIzTipJ4hqvK+1t4tQD/uOo/epPgXNYhFV4NlfHzGDO8Jl2v6ZtVDy7m29bCsR5H+
RWjRUa86Pz2kVinrvwRvkBcuOp0N8nz0msXqQLMn3eoo4+c28zgkMKW7E5wY1eO2p9w+yZaUZY/F
NkwWSMJnP8yIgjrsD6O+0GcvEwhG0sLZCewCr/wvKdLVyY0rRDv8QXzzWBcQaQ+2O07+VWBjD5jR
IGr+/u6nykRE2xEpRRKwar5Ev3m91Ll+sBa7M58MDnyGJqGG2fz7JxMW1o9SKE3c/e5qgfiW7ZU6
uTyWSV3ZQY9SldvDGP5Xj0CPChA+GBI6TDsb1Mu4tPxcy5PSQ1qnXmYKBsaGMJHn1MxCptoxMqTM
nLpkelDoO7Tj43JBXVQsvj9+4dCss+I1eZTcUN+mxI8UFt0p9AG30l1ua5wJ9MaD3j2+H7UElvo0
qom886+mB7lcw8E/N+AVenPMfF0MLDwD8/v5bDI+Ri5ghC+1ADT7iJsK+2UZxQ71BQ/Hhm68BwDF
Cqk+UcxInqMC4CHpsYX+iIaO2CLWXNrq22819mrj+yscf6fGCSZGvzSDpbfws5cPqn0IvpdlA1e8
jTQEfXZfIMPeaa55446eRxFKtCCQWz/EywRcij+3kq3TRrEFQDzqVmyYEdVIBmGh8b/xqe/CgCt3
CosUWi9bDK1crYtARG97W4Db1aUeRavY6g2fDR8BYLt2ohOQIw9qLanqiTdGmPUvEb1jCaVaMVU6
AKfXaiTtehAe018gsxBIYJ2WukaVNGupXPBxC35s08hnwFeg5TZwxQIe7qB3zxy7apYwHNL+ULqJ
1OXSwf+mLqFqRpunbPD5nVLPOCY3Q1j7iYU9GFDelGLs0WT2COhuprq+kkBZfgsr7/UHepBj+2C2
jT6R4DSo9RjZrrOY34z71ZRG3yOe3pvQdj35rYIorRY0Ks8rWHhkVYTmuL/qqBGEL72jfIke6SeC
5qdNKlUE6JOl+HYpEjsY1KPFw2uI3aSxNTFSKLrHWEYM6EPPoqe13M+kLAuledr3SZAjKOZUCXp6
ua/FC4il0OePVXR4Ur5lg4gDR504bQgKlm3mDlueqmxE+4tdUsY36GCn7U6nqrEgEV58nUylFUZR
GGqAWv+8KsCFisedf0h/dkVKRTxQiWHVhGEf/jsPsJxUcBDWx0X/fHdgOyvby7GPiY5fKec5rBH9
GXPzMA9WeoPU19wP+pUDsvphSmGbsaoQk5NKkeM4XpQrkDyoudCTOZ+rCbtTSbDs6KNMxXq6x204
ncX0uaGTsEIPMK4iWzWlNqvOrzh7T9l1UIdGd+iZ4a6HuOgGfh5xTa3DWKjonoZcEByl/Mtf32Bw
J/va3DHkJifSXYt7Fm1dFryDPm/x4Z40GxkihQoSrPKLGTaizD+YlQM3G8XrjLXyIlvNwzSlsydW
ZGOuM4wobWGVhH3LVZChJVMknZYSTjn7C79QkrFNC6nI3W8HnyBXXJ17KcOMij46DKqfJ6BU4/9u
jJhXSi25F6n1yxZ8a8h/W6s7t1uZPSne84jELEWfEdc2jWMbp4bwa03ShQrhTKO54jAL7nZegioJ
h6yL5XWji3s7Txus48Q5GY/AjJVh6azuuxhvKDu7a6V4Z5vT9M6wkwAifRte4wTubQcYTgwwjt8D
aTXVuEZk44Fkmg/SdDD3JjE18Wcbe2Zm5pczvEPS3ez+l8tsuYP0bd/iXiMHeF0jUHEuMXeFhVTG
Dl4G2X+0INxNhh9G+PmYhqfvtFp4Q7eDQqkpO1/BBVUsxwsMFgzDkFaKbmBc3pJ7UBH7gAUPE7Kx
idgWiPWXWEQQreaqRtj6ZBv9ybXFeKfC0LWZsMg3+6PdLNydpOIuuFOOkBrJTdTCmYAe872StF3f
sQERtDaFbHr6dfIHU+XVlisTJCI4H60ybZn0NO4gK4V/qez4glqwyNJZ0JcNh1rrkz0r8ff7JHe5
uwaVYDZymU468+NOkWOBvCBT5c1bSw4ymeBYwGX3f3cU13GtRjUlUYXnqcMM3MQmarDmlFjZJh8q
KPsL9DLuvVAjNbkwTBGae8bQ3R1k3QOuPUsFofOLqmiH2eqvattYFm8zxlaByaIvIE+LIYFnRc5T
lDZHiQZpCVSMyHt4Zo2J2dXg0kXe7zt9F1SW44IhHgh5zl62HOqoiGjVPy+Z63/uWdHeskKSleri
JlkcxQPkJLQ/uAkC6sGpuvnVlPBEFKkANQq7JutsnxLRtPz7cmGuozDvkssQss1k5N2cSeMcOgTo
xd3/Cxhg68k0DlvsHNxagjR2WHDby+2fsrBNX1+MBpn71D1Y/2br9mVo5YBVGldJsDcGEHBQdOVV
HgLS8DUv4fAqVgD2htGo1/4dNIlLbU5zYDEltcdiENui6vgs+QqtUs4T9LXRq4RxGIOheQeg9lDR
r/ODVj/NNPDCCTfagVmE7Q6d0wqJx1nsFcbGERTwvo0bRjHaOBUHgq8daPrWYXsduA0+AQnRyc3Z
b0JCTXUk0niGgDVcjGu0Y54JAD7Io/kwTkY6xn8mhUalJIV7Kg0L64GtxYuxQ/piB5yfvbQ+jg9O
wkeb3rnwAtAGgOsRYpeh3FwvrxRpjD98UgI9aUMkFu8d7JL3zwROyJfKpTWOuVEXSrYcbcSg7Grh
ewJL3h6WxppB9I2bv+/4f6iG/+loCu8kfXHHCdiyHG4rdl+0evSEMyj4aKWTBy07Klkg8cc7521q
yCsHoNFoWe/xxI1bR1fVYqNKey0oRd4p9LPzHVG8efmHPGsXSVFK0Fm/7JP2wtufIs+ZI3mNYqay
cbHUZ6sXBU4FxkReMCTp5LQGbFHHMGHkPkOrHWd2dE+ICer+h68vUFfYhAax00iIJGE8FL9FnYTD
d2kaMIs5j95rnFGEb9gNk46Y+se++cdPIT+2xHXiWCtM8O9ZQk4d9fbNyI+FZNnvtttcPYmEiLl+
pRiHIie62MWI7whRN+IfJZ3vnV0ATONgQ8YEqPLhKQetd/YA1Kc37iqsW8MLmWkPGV0IaUMubU6S
emTvbUtAZPtSkGmL/EhPwtDyEkvwPKsJOJjzaPrgV5V/VWfD3+/jpCBQETTqpJTFK7S+1OD9xMXj
7tUxpNDakUZrcwg/2H23Y63x2/MM+AykmltWuKQLFC7nx2Mo7N4AY5iPfVXr/iWIkrfcVKlNL/lR
PPy9/9Fj+4D/u/cjAulYeMtDkVZff9skp17UW+/90hYdeoYK1veWR1OIzzYmQDOyzwfyrlJNC5Ot
bV0WopHlUaAV4TmdOKz0EOSAq8glLNqt9yDNrB79QWSKVEU9KU8rkzDpP/9/kxqZBJQSBlZty9o0
YW4za6QFZqicdKLQAzr8OBpXe35srfW4n0ugUS8zia8h7BbkG8h4aNFHZryUwKyISH9fgZqfZzlW
OMOer4byAZvETV9m1bk8oRjRX4IbhpBi5wGCPqwoqnQp6OsIdKkF0BHJDrc46P258AUtNFsr+U8q
YRJm0ZAy0+R2o8niGC3LBQLQoOUUn1ECqWn+g6S2qLHoazBqitxD9jaOIrGi4EeIQdTAPB9hk7QB
NAwH7W/INTVRO7KeMGZ2WuJ484vBYGvR1Xmj5DLrDi+K3Nf7bwT60JqV0Pwlf82uv1O4OkbsKGQJ
cjJaXfV+ROIuasTGE5hSLuX9/zZoYQQ6zfQQyuNNDS1i1ae81ro+Qhq1lqCVpqvjlaU/yNWPxPBh
2P41zNfI2vgklny0ISYKmmkZYPyCF6DCapfwzmxEkJ7FlTTNMloulm+fBH8T5I7jTaO7Z7ntC+u7
t0TfYeKug2/rXx1XEGa4YG0vT0pxLZ7GeRpwJnQPu7Q38NjuVkoMK0k0BS+s98VodFrPGsGPub/u
h32jhpoO64U1E0B3nGCmO+u0ytukxnPJA3D6JXnWearuAG4HCc2NmpiK/W0maeqpQNrSB5fQN+Iw
zIlwp8svVSEo4gSGb3f8Kli3n10gyb1fUVbR2kPZQNrhcWGz0UITiY9oarsYEw9awk2fjPGBp/0i
QEJWYISesP798M7Aq60kZ3HUSBVedcQptJUjTegrrmY4ftjXpqmdD6xsLcF8PaD6w1RBcC/Ru+6f
ISEWvFvVCqTcZZlWguLDvv0DWBKXCc+KcocDeAbLS01WDRDIWiK5SxzIFmoYg9801fKoDMEVjSqH
k0cx/uzi4tN6H6G6RmDuYIjR8HttEzH4rXPo8upJKgP4klDsf7s8l2gU/O4jD4ZjjHlVNAXIh5W/
trce7LVWBeCiybOnIIS7FWVodecxI5cRRff0oBHG4J9Ya77NTw55HWoNoFzbHOvDMOuQdEv2x/TN
mk227lXxSSeA/y6Zb1fyIsr0qvQOpc4HqvzwA/zxc6ttwDfj5hwEefJMY44Ul22nJbieV2T1Vqj5
u2DoQ6o0Xe7tZvVaklPMy6gFf1s25uMWEDZD+qZtfJtCLsFxXKinTb1hVeh+K7DH79wsCUVU5pCD
RlmotVeUZs3BYDMHim9A/Uu93RvDC3AUs5j1hAOotjF36tzzToyXXsiUbCj6LvB8zwaSPsSIVrZn
qbvpoaCBFPotCCku8iitAjw+lKCCH9KEhUdMLGtNRIpxBFUAD8biVHstM8JA2BSeNmxNFP50WvoW
UhRCSHx20O+JbNdzO+yPkc0Wgbb7nOyuUl7+FgNi2YI3Vzd/P25S8AC+6qCK2WwsiXxxO92FNdSP
68JRwJ9XLVXDT+xl/BSkuZ+53xH2QHR0u+rp8F/GHuuV9V4HrpC0ZPa/pUTalIW4nOPtQOGCGd2T
dN6ZlXpGgFPPQ7hycteXvnaemQnIYT/QtZlX0uWKcckN1jyRNFn7yBOxMMPYCsEBKY0CUhqYrsqT
fZezLu5WXrsT9C65AOm0sVrXRfgOMQAPHVJZ2UhR7Tq4JAxkGIdmZi4xdfKymcJqJUJbcsXjdHTb
2R+zZm2MPMo3pG5m+IyAG7RCLGe96v3gXke6NOMepve3iCfuPJidpq9BWokboNzcs/daB2fEnJZA
/8AvDCJ0QtVh19MpODn1Rc4mJoeiGDWM9e2KbM27m+q+2nHN0u9G+HUkz2y8SZH3i1GnJlXeWrMc
U81FZtEWpbvBqRpkhYcpzXtgl/3JQLxrC+zXg+8JiPeZ4gKMgiLSZqabs/K4PBfHS9I0GvMBcBFA
qRVOk7i5WpaFsyw9bbd0gHzY2NfA5GgOLjt2E/++Sru8w+fnyT+zuoxHf4q2i8vHh0qBegwwNnBz
0p/o6AAT/SJ/i92WYWHvqzpBRlO3CLbk04eLA+qH82AgUAIx5DztqUr+5mfjLS6PtMfERLmGReZQ
6bSirmOBAxt8e0cQzeUxozpCorUYIIhtkECb3eNZOzMkU034s5EI9A5enqX7Q1R6rI8u6WIoFM9v
VKRCGhTrv6OK5OLlrQLsfBVT8PsUOreM68VSQNSkgF+vH1QoWJNPxcC9+2FLhcq55lMtrmWrgugG
QRiZFUPOZANoJiTN1q810v0DElZp/Kf/Oqv0SNm0rfv4KPsjd9Hd+QSOXJS6k8ZgutKXSsYlO29M
s1WOq2i2ZqdqmyNLQOiZ3nuBAUHie8L824o6+JkhuQ0VRWk8WE8OBHPjcVMKcN/05MqX/FhExu6C
xG41qxtu3jWExfYnueh4uMePS4rDp1cd+BZ3MvckhaktLF5TeWmr2S6LER6CDiwDzQI+FniujlmT
abjbXmMlIyHb9xkrtESshyODeJH0YCYv/nUuQV3esqmAkk2DamdwPBsp5PxPT155c+9ERnvG9G4Y
sQfFhsA+fecT28yJGSDkbpKzGDctaRBySc5RLHEQOlRM7cNbAxB0Lzhde9h72jC47pcvfK/yf0sT
UmkSRKNef3jrdTxJiZjq/sdciOywedM32BMxT0be6j1auO/lKB1sce+ulilztlg2JawrEW8K74lw
h9V9yo7AcZoFkOVMrgutWHOyTSvdrbxLJGmTN5a2RoR6XTycqX+iJRNN0hqJ4h1fPGoEsJxzebuO
+EDhaerRGnhnBhTR/ySDajVPvnBLiIHVeCmj6XWDTvroxV4JkUI8UGEv0K3NBYolir3X/v5XOscP
dYwwcdL38w75/7W+O/emVCmmnmKPv6deF65bGnvYev9ClHjT+MFFzAuyTlehe7GiXl0wV+eaCkzQ
X+AFEIRlqZeLZF0uXuLiKuqRxM6JrgyC4AASyU2WByEr5EZsO5pEEOjC8GRUmsmK77x/PgIW0Qlj
ZKccz8TAIfE3lfgnQz9G+yfW9NAutSBl097on9tfz/GxsG/Ugj6hsJH81PccXiwMgfhEw1TcxY0m
ZV0MUplVqkTo7RoIlInd+9/sk1rchZZ4gb/xaSmJmPCnmaeDfmQmAhXDg3ThvpAPudWCLDpNNM2v
A4ZKlIC5di1nTrUXX65UTJKshqPBuyaQhGJV/BDg7yXZ7zQ2H2zCuEd//lzY6df/GAh61QdyD58z
uFz8YJh0esDaom2h6DzEYKfuP0qAc8V9SQfbg6qYuOHQEx43WOerbpaVRLhv/YKC8UM8PrOrjrE2
CwQF3tSb/2cFsZXEBpzOWGpUeLA+jsNyXZN2sez8TNdfI4BD8daQ41yI5r2Ue6iYFKk5Sc42Kqqc
87ugds8erfpPUQAiXdTJMrgg7yj2Vk3rxhDuoFm8dAFdOV4ed1lyYGG1/2ZMhJUi7lwkzOAW6HE8
Lcgx2c/PFB596TIoPyNfTTlOE9GReLbYnZVSHa5jVZjHcxobyY0bdmHm0RJR2qJ8CZbN9zlJdmdN
4/nP8h2Am5Ql25AxsMdLTX8/dVIwfKfhjKN23HerxuGk2lHZ1sOkeYU9gSmfFLA3krKPcUMt5sLu
XVq7z8HyNpE3FiC4691BEgrsIxPEfPRgliedhvX2JupUZdLlP6mR41a48CONMTn6Y3+6S0u4F0up
e7yig2mWu+TwCwqv7jQMLG5PYicEQlz3uHfpEPhruU1f1ojv9Ecmz8BjJZJgO5MSvh5blkPoL63l
3tzuqnXTlENYdBF+RQzlU7nC46ILWwACZ30vLPvA6X6wQfpE/A3zYPKRYdNO+3Fy530GUy83lbYz
cIVt4EKJ9+18TwVB5w4x1P61seycXs55ykj5u9udJEmU95dbhknvb14y5/hEClMP4zzAQeZfVTul
rX3SnLS3FCkK3Fztp6qHU3tczACpltd8MCkVjFUlm/Wg3+ghfDouo3VehoOPADsF9vdjCxWThIxL
uR436C6nG81qZ5BA3Q4WQi7I+ZQfnrKytiBG+OaWqteKEdLOkt8RdDXFh76LK/ae9TA+pjWcHIXq
fwTWm3AKTbRNchQTtYSp7Y3Jy6UsWsu50nsX8sAVjvKNlI0jJR7UT4rjivh43mDAyZ0lJ9XFII6a
hNBQetmVN6MIYaZGWE8YKDNyPHkdXzdHDwNNgA4Isvu4wP1SE1bNaemTTXPYj/Lob+96K6lmGExb
kHmIab18sVLQSJLORP9HGUtjNeHk9wCZtSouf4bZl7OEqJzH2YzXYSZQgpElYdWhhN7D5gKir8Fb
sTa9Eso3u9EZKJ7wOOV+oM3edOq7uq51oBY3X4aa2dtEBJzL0QEmEIbw41VRA4rpkd7V1UysT9p7
Rlmm3By5JnGesVfIKCgCuV+bZRayd0tsgyhDq26xAZj/d7XjVL4PX10/lX72KU4/3rvkVMM9NpON
ff5jfV/Q36XytTt/6vL+T+yA2fnYNmK9aZ1UYvYNcARCqiQgxjIfNM5Hf3cGwIUejjwEL7xqOeu7
0WwJjKvsmxzs/xS3IKqISKAYjjPtlokqmskJ84/vqg5SA2Xyo+MD6obwEuQeHoY/IcPGWWuyEGL5
Zb8c/mGxNjiNt867IL3vzUVSC9pXpPdvHc6SM/jFh+7UCD4HzN39vZSjz0cqfQIEy3wmhW9nBYuw
zb2bb0luVbsYbqXesDehpRG4HhuoABLdE7cIhGxmvPb2eCIdh9vxh5HSBNaD/ZPOCbFgNq74lfg3
ILJtc0Ti5GnpjPzZVzRMQBWWbDc/gl5n37MiMul5VmEXrSW4/OVBDsbPb3v6P0YM4pKVwas4Qviq
KzfkSW7JzkNXsgnbDfUyCgfdRNVK3JeOySBset0vLaXbR0D+KfFdmlfjn+CjGjT2NKSDE4PACjzz
nMSY7p3O18Q68ZvjGKQQpWLdAWqDtgEuaEHzwwet59cb5MKKGKG9GNAF2qociLQhBaCQo3ZY3Pmh
vO4y9rM3Cv+31Yxovcsn5RxBwpIp/zqyJO0E0j6WfrJOH2lqH6dgd9wvjvNJRRtkknJ57eUEILZB
iyJFzcy3QdlR06dOPAb1p7NvbY/iC3LDZktc9g6alTcEqpZqPxv/qIOPsaDPr/pdP3HP8N7kr7rO
c8TzZ7OVeR5xlKtTWvuw+0gA7KhowSgtYsHHgWeZohr+iI6AIF0vXP//p0/ly4uDtG2W8l3DuXDA
+FXnhL5DPyxrosIFmoRJtMI51oAGiVRpTAs3Fn1VGaMwCYkcemgAnYLy4ETIfsjog37KtAAi7fVO
du0RfJ55K3CdgVxZ7JfS4NRu4IPsXFWXI27V21rWomMUX3adtv2qelEPHzRhc2yzjxme0KVDreoC
4LzA0hUOxCDsAQn93i7baffZiOKFhu1SZjhHqTPnb7qI6Cw8yQYRofMyKbK9sepKoa8iranUcN5T
vZ1L50xt6uoqaU+DlRDDju3F5/6Ibmga137DCk2iMTwT+lEQeXO1zFeoXj01cJ2YAYrADPEAOOpU
SB2GcY/DUag72sEa+UvZitLPwr7LX2bD/K90Lqre2/AhsuXbY5Bg4dVa7Fefc44Mg9vRuPGicoGD
lj5zOpKBBvAaVz3sveYxafygQpkiLijUhApIPU7GKcNxggmiGKrvvHv8WYjNEuf2neYtp3xUOc2+
/DVCxm8kv2STtpJ6n+5/qgB0Nva3Y4Pvhqx+BbA4QOdSbEJFrKXVSjAWITw6MdD+Ayg6W+8IbOeh
913oVCFl7e21y/2D2+nPDyJIpIPCx13/cl3bI8pi07uua/VkFtG02IoMk35X+6ukbmb4eyFhVO5g
KdO5LfE3kr2k2iA5J8zaaR+MkykqG+eUeTVxDepyjYdoGyBAOeZG4rAELlgmkwgptk9kLvjUf858
r0CpunPo30vYHf1GBrKrLbRo8M1uWrqrOtAFc8FCF0HpRmuWzWCzhpGD+xYo5OZM3XoizCU1Ncd1
Xj1f2qTslBaSSHo3tIpZDSVgpPeUwvlv/Gy9jDarMGDfNUESyfoQaKu/1m4wb0oasfFS2NOoRA+3
QWj4cClNlAbL17FJfOBi9LI1rI62E6tLrOumuD8zh2OwdXnozaUCEfUxU1bd/pYkOinVaHZoX3E9
e9Y2FxmXGVEVxAC+BSvuojndoqoxrk4yosFfsUU8szhOCZjtjUzJhzYWqpxJs8F0URuq6V24sI+h
DcG4MMfrNamGs4tpJXroD2drR39kKo6AADLpyJmHz+4vZp9F4xYuhKhuecUTzFC2aM89kAbBcBTC
lfILNzrVVQQ7E0xO6EKytDg4E1J1ox3tuO2A+JXkCe1VI3bvyRtUdJY6nWxvlVcnUqpCPL9tzN1X
PaN3VUDHRY4q+5UVnhgREw/2hhmFh+f7wd+wwYvFTyRwt52iHjkcw8OWkn+I7VkBe2zpJvVdKiiC
KWXdo0KwFBAdvhkPvQOnwuyvXPw1mdTx8O5viC2okyRUI5/drHOCjktKd4GaazHGXzp79YAdUp9a
nQ23aApadHKFJwFFAEytnDKrYJomAwC+KYs4d75cFZPsJvNhyHu4LapIfsDfBmjMs4SBn/QQ4gXa
LSEyMRTcSxEmEkt2zqOhCHWL3C74NnVm87j0pNbo4IpRMquLLj7oFB4HMIfybxjT1810S3HjUrmz
TmxgWeVmVtQ8o1j373p/8WM17lr64JQm8VtuJ4yBXOGkj2tPbCFKSbqSHnCuUhigzX3DCL12GR01
9OukswTMABkO8h7Ixc0m70TMz2OlPPhLyRB3imVEMI6nmuLPU/3gt42J3Hurqh4zi0rakta7bqGG
4a1W4zGjeGwHx+44+QvgUjF6OSh1QhnVVwRi2mrsqnIVNAvZrIuTPyKRMzeEfXjRkCyFv4+YsP+b
nLL1lRzmwqrU+hvV+gmPWiEtEKz5V3CKMPKdHsmeZ2PL6gcMZvTcfwLBQCTeaodnx6RQBKfzoSNa
bNMT1l5LWWbogwjL/ho8F5FtYNa0/Fg4Fqj1PzAgKoV+VKQKwkbj0kKHnrKF8xrMqcWq50Dg5RAk
OTJTm/uYqV817g3k+iPbgyWx30ebXZ+IPti3z1MGh80QDdJ82nSDoHktW4R1H1UUuJu7H2oZ5RP5
2V5wn/C9Fbk04TVrlH7VDEI1d5mGix+RvyEL8QioAAd7yA6oBvCwdfRDfo7SMEg70g0U19As3q9L
PeHWcNYypBBYHLZKJa1kOKfipHREAZ70WBd7FJvRQaPoNWkmmuP7HY7LhtfYpGTyM/09saDGCfPQ
84bx9sGOdxXO5bNcmSEyr3f0fERNYcC4wVMTrCrvgDApkOSdwnjz+9m0nxecQekzL9xVKSDH0Ufh
Zr4MgNRBFq8HYNhfpcfpu8m0iE3bjmKnJcwxw2g+lS+7wGGRNDbCP/qVsY08MJtWwwNqdlPbhdQD
jjN8mC4+xvP7o6wmeTFVlwyvZjnWa43a0piPE4TcopuK+fg819PgmrohKjUojE5ML6a5nkAyQUFz
bWIPtuPQn+yLNFYwu+b/B6/si39MxegmZMU/DT/svVNGM85viTl81wBLrN1QwWqdkTeKTa+7IUPq
3ep/uCb/5N8mbYN3uQpTxLVWNlHJMs+dm9K7lihHwrAvJeiq9lFF63NyQhUaEAXhBeGD7WCAcajZ
d29UWjM5KlUaebIXgSOdczB0t8KwKfHHOrnooP6eNdsFSyD+UwC0Ncj3BYkmom8QMvqD7AV9tO+C
CysGF5tbNodcTrcO/8UteVx2BfUVgwSWmbxzswwSKCIGwIm59uQA0FduUSeeR1iwl2pTtabWlpK6
XYhMMlueo4wm0abnZRGLp7zE92zp+HS6wNh7eWnpjiKJbJBvY4Vw5xT9ErXPQIh/HH8g7itutSBG
w3Ef6EBx8j+IwJhJU5gdwiBeLduzgTrAAhqb0PKHxiscaN496vAYkQF6Jxvh0tPRDoFZMZWE6QNn
WJPI7HpmrOhylW9jhOT0BK2kS4w1kuJaoqhGWbSujN+zN1pGvIISpdLH9m3pYU5CsJROHlyXLS6t
WiJG/hIYFKXtRO6ExodsQJ6+r3Gyo2H7wM88y97Va5jXxeIHAweQ4HrDG9YdYQhLYQHQmYT21gaf
8K1uYffZrNNfmIuCbfOniy+KVouyfgnDmeolRAMJNdJZQbe393MJCwbIDJag2CmTsZHSoH+3W8ry
Fe35Om71341h7JAat1G12lfaRu58nNZhA0YffTRrl1XJ4isYMf2JQ0KQ1KFO2ypa6iCEV9rOwyuv
EsqICuZQFPn5bz8KgWSKqlT9YlGQf6Xgg8HHBH/E6B5DmlEYFHAs28MJCmOJgEMODlgN+W4/tIIA
AmZ47TSmbGxb2aDO2ds3q5Eg1d7Y5XaiAn9y7atp4tKb+1YHetqcXwUm8/bH+jw+XIT9nJulRa8J
HtZL1HqevrRUq1wZC4iTxuJyKRj2TeuCgNiVuvH8jxtcP9P0sYjts5RIo8IMHPSF8rpMKPcvCM//
kahI9CG1XyUYPOYdeYbFTVyO/0jJCD55oT3F9Wc6xxg7Vk7CWzCKjvezRVUkIA0ECsbqyxUbcXoQ
c92Le0OL8actjTJzZr8lf+tRTxxMu4ROzLmZNLnfItCMzXDKrGoFswd5ODLwtFFnZqqFO03zPxqX
tQjB8/omOb723F9H8iDrl7o5tBL295/yRXsnDTIj0+ziVwZkhjeh4MPDc8MwMFiQgwI2Esc9gRbC
mnkf9Z9R6gaxwpVPlrA6fAHRwEk/MzbYyXAEE4qLBdsAOxpvMRGgRhNgEB1lsS4kv1q1C/1N87sM
+IIehw7qghSKNnmbGIalc4BqmOo1MIyLnPs3QyHapq9+1hfrJNPlYZbHGP2/2MsqpLwpN5FjSuRr
PBkXu92LT4DV2uGDqSDMaNqAJO0/ExvQ/c8TVpu1aeCGqlCZ6UFtuoOr003CeFDHTUTAF+8eEg5f
vKVFC/+rPrzq/c8LBh8exOq/MoyQhVMe35X1W4ury6ZjA6nzjNvWcW/aY/EovA4BqmjO8jsZ46m1
1VKXzjTfkuj91ZgoayAh5vkuGOMpU6XEuRlK6cUbiW8tOvXp7sNmltRxu3zBolJpxmCV8Tq+Dud6
9luFfNs9VYCdrlKjQ9hzygS1M+v1wUN9AqHpEgZWrCScDwPUYdVQ3cT0103hYrL8vO7SkDN288rC
d7+EO75eWssKx5SCz4DpTzAY5jGEcNHr2q+y7S1xM5QWI6lJ5bGjdJi38zJNWcZRSnKd2q2jPKq1
9UEvDY3wWCMjq0seFdhI2tWaqJXcw+M6vafmoaphlvnSty2MmXUrb8nt5lnGpMoYaa+GAIXPgf4l
cBxhwCClmttG8fdsgjzpcIDwVmJyiPmP92t5//5iLc0iLNKguSekaRUYwGAIvgkNlFMceZY9XqFx
zzP/I0dc9B4j5IdDssNqsAOE+E/E8hJMeToK3EM/znwsTpRiT5X8j/1CG5HblxAHBIkIupllVF/e
9DnLvbLu33NnvpDNLci/Q/ET3mGRmoqpKAiWju8isAK4Fju85LQjSVnDe5UKHA4D8uggO0cobA7Y
4kmVQBFfHoPQ/NiG1DDQreZ/PLO7ehIXDm/At9ulLafpN5+UG2hwD8oZSwFGT2S+Y8Mw/W1WZW0+
cEAMDIBdQLkh/HOSYpWkvy0T8W5A/RhHg6v2OscVSh/FUZTjXlvy37bywN4b/hKdcqjrgOI9nF7T
7tuwFVtM0s1O4jhMuq4YpCityfM8kwLpS3wEfQZANazQFEyVm4zXCM3qCAh81saL7yTGI0L2J+Qu
jmRmC02+AeQQm/5hmKhdlQuDAdP7nFv4sCZ+zq7RYHE5ysU2ePXLa6mPm0infBO+c2bLB9GdKm7E
0TJtz/vM9CLXir9TokkmM65xMkz2V1oyn54CB2yAYvzUFrz6ytgHL2baU1qeec1HnIHfcf9v4DAF
CFEJmj7KU3mCA7iTACIsa4GNQx15nPQXnU4ogGwOTy/OJYW2yvRLuvE5zkOA0I/zoFXkADmjtCHy
M+N/VvaDNx3mN4DC/ahILNIbFstizUblJGuP4FSfqc+BVgllcx4bFm+zCYl65qux0LbpXXEhH4ar
fVTBf0uohFCRcLjbWl78b+LsLFBNMXVUWuofZ3hfLCvkaZyaBEqqcfeLhrT2XGE9doEfR2RRSt7X
pmecc6/c50vfHSsNX0z8dYcGWPUDZdMTvstlqlIHW29cHxEa8DMqVA2pssbOnVlyMZF03cFyO2YI
ds08VXlgtLVCADVlhLGlL5FaiOGqlxUtplcGapA+vojXKeWvf1Zu6XInj75KCZVNebQObNzf5jGJ
IATmMlCWPyjSUiiGhzmYxPX8Zm3STj17zpi2Akt7vDZQJTsAohzpOIADhR7CpaFzICD+2IntIiM0
zxMjJbsKWkhztk2aDODP816IqE1V4Oh+lw3GilVD/a+aJ+Bwl7C8ffKxTfRpuDHqOVOMSDwq0jWQ
MY7ylT0++d5DjlHqVMz0rhLQv7YJijL4gJ+rOehfPARU5do++/0qeiIM+jEFFc68In4W+J+vKONE
jOLKeSLqMnZjQTMTt43J5GeetzSXTbZeJFSdwoEQ+8zFBThDonRZn0XKdbMLQJbWarZZc/HKY92F
k7IBqNroos6Nan5mlkkAQpQUJ00OioF7hTv9uETvgb6ApHioTJZgbjbAANnpVa8yYkigUdJ2sL9d
EO/uLGCw23UVqFci1H4gYUxdAOXCzcTcn60CbrPvsgW2qL/o1r3JQitLUc8HsVfmYncma422AzzQ
2sc5wFmaJEDiiyP3knMsigP8jQRfuImvuRgNwhnqqRZe/K6vmQS1fZHICb4+iZPTcEVbtIapFIKQ
0bcJjrEhU2Gi1whJndTUAf40GVTf89l62/1Bh7WEojsgvVlndJWQulsJxlSxshhyWZj/GIxL7aDT
+Ne+ziO9Bw5JOnlXrgsFDD0qiMRjstcl+Bosv8DWpscGUGpKMigDfOsxQxrybydXfEQLoHSxf/+q
y7Lyx1nTib7HTxHxYoD3vOiYgSNDUHdgQKT5hCq5szIGeAEcROKfb9QfhNBVMbNyXTISfLrWleYo
D3giRzLK1a9DPrcPZ20q5kwiCH82aq6LApuaElW8P6tArwv+CUKKAWQ5TeIBf3WqDBvx8R6/EcBL
Q/ZQm50WbzoZLE5zy0zWXZykyf4gwGFgrBacvfRo85Oi2RXZmYIbqPIF9xMPgB0QiCWgVdQLhtmB
xBHnbxqisDkcTYkPxDMdZE6+D3gNlzaCMiju0JX2ne3mriGbhjUvqQeY+2OMd4XN1fDakttGwu88
v1XRS1QSQ3CM0mtsyDmjHCmeZFnQX3LmGtgwGkeXdeVKX7EaWw11yqPf8OYYgW0OKkFOkgvpUw7f
JUASGPjs42Goze91/1p4iJsFGsK5gBD3LMQASkOvTBL9LbxwR0dLkPtQ5Na/pHPHl4q4vJ9L5Tme
uvW2XjCvKr6BpJ9NrT/wF1bEnMK77A2kDBw8LmRBtaX7yH5l8hN0e0vkIOhEmsjKNdFsUGbcrqTI
c2qcilUzEqJ9KR1F0YCD+SZeu18cLYJmNk0OC2A97SjkIRwgBgJRm0lirnwh/XLwMS2gJHtjpEG8
pjhSv7Qwv9fEWQT9+uooytAS1Y54i5xJ0GucjW2mvqYD27L37ifqZZt3fWFKsB8teo4L7ux8EQkA
14+0jEn6NKFESLZ1FvQCKxS8wcbUXvlNga6NCRXRN9r9mdJEkwk4HFFADcg8NNAv/uX08h3nYUCl
1VihrFmj9dL+cbe9kc4q2C1L3i/XTDOpiNc31S0gTtqGwYSl/ieCQAY3Lge1ZHvn13WLfSAOuvFz
Hbu3Lf7ZBIsjmoj6YzQEbDpm1NlrTFcQ6Ti1jPrKIreR6BlEdJZh0Dm9Hbb+ycEdkbDHbRGDPJLr
W02dRveIN34b+ADgBbzu7AGb9oUiKcvqzCSRbmP4XiFvQ1ZTu+Oqc//NV7WFGtowt4xWdHk2nBtT
yNPfhb6b76E3I+Msg+VHCzrTybvFxlfmYokH/vqUzrEbUr1aWFRyrWWLous9pZDAVkIvqtIaLYmi
rkCtcMDIXDcweoyZA+hb1C0DJybWT8Iggua0bn5LA+6wHgDC0K+9oCUwEuawOBsRw7S6365Jj323
pBdZmnC5TLdhzF7SLnJkKDvM/OtRYGPfsPCIiKUugM7w2XHA6m2jfQFLj5by4TxqbAcw/sjXPeAF
x7RYEp7MMngGDhyQAx37/K2du5ZcLm+jV1v3TfH6UFDUhAzJCdkR6QwqFroOr6kCE8K+W02+zWx4
KVwlk8TiHVIzswe14FAtuuMTqea2rW+HCjZl9w1uDHCoaOCz3cMl6dOa4cR94y2ZypKcKAvY2pbI
Xmpvkzrs93dpCq1dsoI2qDm6QyOEUlhSDYUpfZmXkJ3Pkj47TuwZRpNfnixAszDJaXpaEn85e+Io
Kcnponc1lUoD2lTSOdGxz8iyqPxwWW8dWZc3DQhyGIMPwzkP3zd+DiRWDyQno77rpbefT518rcQs
W/9iyDaukYQ//weI1tUdZfQtFWnO4SFFdlWEMVdyzGEz4JEix3mMCCRKWvRsgZckIZgQ03hocJC4
R6m9UW/Vuq2IRCiYKuBYk8D+n3/sySN/x50BtznCsar53nduBKY/s5sldhKDd3dwYxLIKMkj7MUW
moFRs91h62RoP4eoomvqxQhR6C0gCHihRZQK2pY6Wijuc7dgDuM9rspfFy8oAhu9fnrK6Ako/5vb
3T4C5MxSCzsZ8EGDFXDQLKvG9uUPOfq1vFE/yI8HqVV+YEftj0HwHL9xypOzPg7U8J5RycsMSLYi
e/sy9C6bfzA5F0NMFMWvYl0PViXPFgLRGmd2PBov9j0K9SLlcsnGoBoFmS/62v/ydfmD6ayeRs1t
8ikbL8oMFWA77CdyVDIRfjiTg65p/ozoUVbHw6X3fEz2sDwiov3M9Wq51hziFmRKeVol+kKmUzu0
Tq41ty2YS6yN8mVX6UdMnZOpEv+MXTGZLM9zIi6HOk615AxNKttN2itoqYE/Lm8iwj11rBlOUYZB
5pGaIl6ItBebuNZmYk+SBP/FS6MgzNIy4sKt29skI1qnILkTHs6wbdH2lqdvNhAwcQvQzTObPhjP
/jxrelc9pLgbPR6B/IFf8eoxADQD1zshjeCXpZM3Jf0ag79U3WB2ewm6pgjKhJiK6Izdv5hqB7Lt
dTANZQRiHQ4+uYMXJvIDiKdNZaSUwECc4k9PCUc/v4esBBRrONdR6ZDvM4faE9EX8YYwU1DAC1iA
wg+5MTsUiX1CaOvToXHjI9SbRozDqYKPdkZh4h/r5yw3WC3XsHQuu34l2qxGKIdoGtNjXb5AmE9P
Z1FnsVEZi19h0i/p33HJynupJMCjBDFTEBFN9kgnU+OQjMmSHZZ24daYJbFRWnHTsqx7juFSI41I
+wFuYmiwI9DDTNvpQM1mLEWTqob0bA4ax1ggrdJpOrYT9JA1tHHYQZGOtDmO0C2DsBiiS63BUm0c
2esQZP09jRdg0Rl5IGqQ93wcRjM+khdFwXSXYirl+9oETx7U8fqJc9fG8rUEv38Ea0MH6Yfygc88
XZ86lg/Fyr2z642E/8af6qSO365CovJUH3tfarYcGC33W2P5vIEXTuaYEmohilcAgNBLnIUrhLb0
OX20FoTraLoG7ILiFMAzX3+cSTCxw8j6P5FFpEoZfGlau79BzqHMA/mL2WNhxPeP08gEg4DQj4Gi
Sey7ofFaNFvWWFbe/9nHl4El7ff2U17MvkXuF1cYlIN1u6G1M0HxNydhwr9oG8AD93LhP0YbkKjs
71IXfZSPTs+TWmvjwAr/m8khjpcn480PxOgNBepUF1UbJ5VNa8r6mVmBqmokCyPS0bvNmK6RUkeX
6mmThuISFY893p7RLMul66c1HteLO444i4GbAvWhLtD5M9AXMfUZLgr+oSSoXn2Yg6ZNbn7AUcrH
YQrYl9pALAtn+nNu9MjYr+X+ZQ/XTaabDs2OWztv7nh47pxbnZb2b+YM5hqS6Ux0991wHfle3zaJ
R0UsKyb7+OpX9hpbR2ToNJdCDUYkqbiIMFWZMj5dhOr/q+2w2Fcj37fKIIbRTDMzWu5bmvdVLVB3
eAWDFFPUXt8KTS71wkfrKylq03Ckyzqx0MjCim/3fEDkxuRG0ms1rga2Sc/tN4yo3nY2qyHnLog0
AsnYdaupaSBw+JFknP0PmFUBdsPR8w0EKp8BhaR1y8djXkKpsTrVAI4L2P3szBiqZyMwz/yvyUT8
B9XOeYPfjKsRrLbPmxvV4Iti+hXTLmnWjeOff58VaxhESidiBUXifPf24I/mJhsGxHdv3u9ZDOpP
kqf9yzWhGwvlwpY5sUxvVNECGs7OOnNG4KqIEiN6hM1ogSXg8ncjvAIf6JUGFY+PCZMf9IQdwCCd
JV+HU+SE8hFZS1DhdnjtiEpLGRSqSLP9jx9jqcnZUkh2lfmax/bg/gcDFNFPuRUds/z/0L7n9uYL
fT/GG9luIU3x88I5jxidFNhRhX9gkXfIL3/xDiOmFibCG7wDfJyF2uKwHMsrCdq4xXhD0kWMMk95
hpyYhzJ5NGJ9VszJI5r8UbOI9bOKbxTvx9giO0V8hbUifD1uzQAFJux+q5+y2afXlDDNGPwHFugn
7iAY7XDwP06mOx0YTMxmC6oiuXAR06wmVyuBlXNkBunZtt/ms+D6bOw6LMKXyE68c1AQlxeko61G
cLaQaR8FYBFbzNpBZxb7iHx3vVgYqw68RLaaRJstYcT34j84OXHNxLqS0yrooLJVh+M20uJL/UJa
iy5l7RMsS4zNYq4rAq7AXw03py3uw02Qain0r/rABAxSgu3Ez+0o5mce8s+FLT6QFnHO1E/OYEYx
IorJNUDa3/cETGVrNxNJz/mM1nzCRslzfwueAR2rYDVrgydsIkJuPCKi77i5S1Bq5FQbm9Z8PQUJ
rqyAQLnh5pWv5hpap8U3vnUbvNm/0RI5WjXGVoedLfomhe3PVIFcl56fznHbvf8Q+PxcVdYCQJks
lMzk0UgfAgtFY2jxhUxP5IvPLPO4Ga23kS29RfXIwGdiPDsnTfjRZkNp5twefUlCPWR4/2r7Q1jG
hlcQxN/D/WEC8D1+6WUza6WK8+cmymF4K4oAECfMKobImr9zSEnropnjLNmZFzdKbrYGa7ZIQYJp
jZSEqpQiHhGLmfTqUaqq61/brwS54+K38YgOUcMMnV7avE8pzUXFMKg60zPGyNmIiaZCaH3KVYxa
lDOhMZIcIQghLf1OYxfJALRpDgRjt2by2rk4/8LjwGTDCsukEJwOnWnYanWTsRSbxJysXMFqAaBt
3/7hEiV/x4mQh8lZHQYuuAUlK7HtPbepmzh7ywNBcBDz8IJcXRmqNzi+Nw2XxfJhp3vg82I9WBlR
0hDJnsUD4qF/y5V6GFUnTmDpgGJDI3hcO9kfpHL8CgUZj1PwAnCuGUWRKtHP3q81CUcBqga68Y9G
ZMMARx9Hy2yxoQr/3fau1H+Jn3Tf7ba3bZXPbZywI2iTD+dO+odUvacNt8jyKsIJWLW1jvhOwThU
k5RzqMii81Z3eT8finSc9kVZnLv/MvEul8u0XMT1jPgHUu5ciMqz2Fhh1+Zk1JDoee2ii6hpMPC4
P1jgeZnowbKhejMKS/7Q/gmGYZoaqoYGQPMvRd3vxnoAmyfO3onmaYV6zK02D4nYemn/SjaA19m+
mraaJWr1mTEQLiI/A1A/5R0ueydxK8HAx5HCoGncOwcP/vDA7BovbjttBCd4TMhMKL9mXvma5yGE
6jTBBy0z/xEJqZJ9EYZ39HlfyV6tBDeLMfSrzu+p5O5g8CG05qie7J72h96SFyb/D1CKgpxD58oj
nWQlFpnS13YWD86Bwe1DFifpz9DTuSDyUnVUzN4P9mbyekg6rTBnLamAnVJwP+60KQMUTv7pJC4V
CLQ3+cb1IpdYebTqEk/V3yUpg3FZB7ganL/Sp+J9pzvAKWnZE5PaUGjBYZi3MY7XaLjFgh1EXBHt
Sy+Yvgoa4lALfkzRnZPqN2cyXLtZzSDbf4+gAN++aUeUKgFHwwkWbm4aBTfFJs09xsCs3fOtszc4
010/SuvO9at+647nODiKjhA9Ffb7qgq8J0RR9eD/c2oY3wPmJEt/FBYAwfkRpkMIqy0sQ9rDOd5Y
+FAb6XwPYUjq80iSeIuAn4WeIB7/GzA/eIPQaO7GULHirgy+n63eUjgEVuJaNMyoKiE1QsUGfs9b
29aijipAhdKZox+kxXyqpTuHdjW1ok6Bgk374Ur1ACLJCYeigokudtzpzwS1xyc9Rm9mF2k6XX5a
yJTsAgdo9DgGh+wFVfu2fHsMJbgeDc0WidRtZ+ka/W3M0fI3EtXoVQZqM/5sqhNUYzX8LbofDsU9
nG6hv++r/Q38GUj5f6CLg3WIbIRuHzGOEhQlKNF65Kbi/Ds5+Hzm3rImUG8qsnpGybwPDleuotgA
Lnz6d3VEnRd244JYsEn92po9B9pyLGUKSVJ2jVHJY8Sm+4WzwFtcTuJNe0OKtQVqLrMJ3UMTagNQ
BhIKu7EtvuYtWO48a76Kn55dU+Re4LGu5DhPZ8fFKDQSPaOTMkafAPA9CuHUQd0Ga/sgmYnv+Wzb
cA3gihg2j81CnszCgzI9xveQUwIS1EegDipSYGaxArlh+26qDd2m9E5gVWuAbLvB0TNYPLDyB2L+
yRfXLirxHoRSPeoMHmhmZjNh/Y1aXgu+slEMHjVDaaeaVH3qH7BWBE0vtH9xMcWsu47p52uU3gs1
qsKfwXgq+9vhBSoKIr8nbGhlPLj3jJSdAUFKXON/k07NVFsaRDZPuJiFGO3UCgM62luUSYJ9LI/u
yaciEnEMAc7Udfn06njcPZVnYxCVu+AOpFcKPG/0g7HbionLUTXauBM5zpxHLL0543gorb0UP6JW
Ay5M9GNGWVFbYCoXwNpeegZzYesrQfWKjh5X7EXW73S+TubaMDF3TxO/XLYSIB6Z5tPjEzPPRokK
kr1+ZxlfBydX8SgUMfOcuw0Jzh8wo2OdgPnAhX9WzkmF1Ax9zYRuuwIc8DmBfH/6VOXMz4vMCzcO
panOEol4f3eyXcBlto9mfOmXptNDE6K5R2lc+gKKEUSwBg/98ieKBRmlTQ4z56my4c53CLKmm5gQ
HgpvOIRoDcSbsqHkJkc1z88gQAD6p/zEHFH4BWlSKXS7PDvTJgQAP86QlRqERd0S4DwfY3L8D81f
/I/eERis9aByDzraEqyi6kuCggXtOuH+qiljcPkMyhHf5inVBjtgvAHdBaO0LCuWTNk9adEY5f90
cgPuwFX8KGfnbqwFs8/3zs1rG2DxKqTYxIe9vzemhu5Dswmt2RSt19T+BC/sxBPsmMZxySt6X975
VaAsH6EY8peZpR6PWnltvzgkFbQQWlOk9r1/LI7s7U0HpfNpUH+MtjKWHoKDUT+VftFOqW/V0iLQ
0VmVN6Y+Xt0Ia2JQfBIdVXEcKy2CtKGE1BotexE48ueJX3PX5w3IgVTJe1pnh8seNft/YA+ZdXHj
qBt506Ijtbb+yM9t/NgUAM3hHmb31ftCfYSGOctfPXWoLDOoQoRIIxrmjH2RdhMNg4UblIgLodtX
fIcSXu8p+10PFFlbKJjQeBpkivxH4wrykP0sFEIjlntjdaYcmr4HMVlhM77M7kiOw8eRlMM8CoAw
XWMl03YZDmyaAIEA9cis1ssjQun97My10ENkX8Y/9h2zW5q3ynnnuhRV/Ab6g7GKnnQQD7bx8Oeb
oUZ6DiuU/McIU5Hkd/byX+w9dGbRQhJwVxLwOs/t4Oo1rZ6Nx632WoEhTE31MQ1xlrMrRdGeeA0F
Qhr980ZZSZb5dvA0rgR+bw8AuiNf2qknANat1dKQtRxJRpTFsumHkaaug6X6FYpxCfH4t/X5bv//
hLw5fZIJCqBDTySZ8nl4FLUO5Bpyptl0ZRBd32SBSr+e+c5tYlO0Id7JooK/fVYzZQNdng0E6+az
kz2fbkZLWcpvUJuF4+OmKgti4nL65W3euYepwu9nvR4RpNnR0XwqIZfuNIiXsgcgzY6ZRB+BpeFg
LlQyaQ95njOrxsSBe6vuzuy5YOt66SHYFqmpokHkddolFuAjZQuwSJEQNwsWEXAlsuNF8yaA/Kaf
2UjUcy6cVYs/Bq80Dcu2VqpMceXXUcUzjeHrjm633xQ28DPERWwHf1So7Bn9g+7sPhBSe5rKVWla
gSptR1aaLW+RJUbwUm4VWMh7FciyE+4IivBjHHkLbIl+DOL6ykRLlzUaqlnLKS3E5mLc0roQ6x8z
EkUjHfdHi73zQYmYTzsMPUx2sqivbej+V6e1FA1Dm/DxyE2OvkDyjSVwZdQUTd/1RkSA60luZ0nw
lP1XxjTwbh4iy0yOMKbH0N2MiY29vFFxZkT2ni8YctE5cS+A9JwcXnV0IXxIu7L3tOdcrhhl0Cq5
Tc9ulpqONlQvbQHnYjMK1MDpoNnLFVbysW0/h1vmNtYeGCrjzchtkQ+5nX3MJETvw42+e2760F4n
0bmKZH7ZBCdepUqEM+01x5SPwSJnrMthMDBSPDiZftdnlrh/3sefFpHmg97LaIgSzyS84ZksuF60
SWfpdn5y65OaovPR76+RiuloO4RNsTj5MQMvBljjc8aQJYx8Vx4NxdYFHEXvGfUf0BmXS57eeOjQ
sPBuHeoNlVwhtAOevWKEUWlufZKHTLlFnP0cdhJxGG6JsskH7YyaU52jVZQ1SK+UQaZSeq4mvW6X
ZYb4GTfWwG0UwrE3Cq4Ah29231WiHWSe1aIwsNNIm5ftQuRSFaw0RoduQ7n4hBlZEFaDae2VLTza
N8yEM2SSyXuKe38VwH9QuX4F05DZ39B8Alf6CspifUS1dkEljuInEGnS0XKjZn7N8h608CQ0JzrC
lRCarhbmSugnzkduqC4yz7FaWTB4MVeAiJOPN5JMPZffhatpRNsTQWgLotZBZbMyhGh8ezIz/s+o
+AEsCS51ZAzjnW2krcFGdXJIV19bVZf0a9hU9rCdr+AdktfOGQuGb/OBlvICsTnJT51wdLK53Vn3
MQvJVDZha8XlfSl5vv8rbApdMKzVQBXIbx59Cd0qgu1LCwr+Iz/A9P5wimbR9vilvsWWXbfkhZ0d
Vu1P54zFRcZf49UIy1WBtbMcwQ/QjPe3QGGbcfrwOAGR0DrNlUNFLl7xzcOLOQEEkfoTP+VjH4lx
eoD4nL/p/NExubIzFxBq4+gfC7spUr0qRDqZZqIsyiYywR7VtoVzlA53jO4ZHFQIbW+SXwbzfmVF
Sl1pKj/xTWgDdV0v6zZvGTX8zE9QBlUeIA+kK1w4GdGcxVjDcgrOPLhKQNVnnimmn1uU72aN7K61
/WoZeD6GyMt8mdd/JZcSqhoRss90CLsVxP5C7CIFWpaHLwfbKbKoR7wP6YjPZme6NcEvZbe3qkBV
PI532pPJ/N+Fv5RIv8Ixu/aKdfkCXvXpzRGoFHFB1QnDNX60VIVmbJlUJtN6OHdhXhNa7sB8loqG
7YvfEDc+kUe7PTeKaatRZxlIs9slKUHSdWQNr0uAm5MkdSZcHqOW1czHQtIEpZBxnzNJyDpRgZPp
9E100hDevNlE70coAFsfy02g1Pbj9TNJRh3lM8y4hg6UG6KQduzyYIVmqTqpHmQmo/2Bwb5Y21Fq
BCjKt0TREWsXJJgwkuc1fkgQns/XF7OWrCTFtJwUIJJnSr32LWTSoZGrw0pxGN78J8k4U+ifAHa2
Mqbfs1zJ3uc7AR2Tmd/ByucuCaJjZqZTSEqvFHMmr+EDMITkgD+jGJH9v9pKf8n0ifPVekIMBAue
AAGhLLp6cmVmyuhl6xJZTCnyJhNCYsR+I+rzkmZ+qTTd15AGkE3F2TYjj7Z44PSYtOB96QecNmyd
HACVgav7aaZ4/LzpdhkPs0urASoiKcEAIdXV9otkCnfMKF8sCuTzUhphP777p4bZKgKSAGxPv7ND
O5AIAAvXADGFQQiOLDlznCjKCBcwjNcV3K6Vxs84qAfv7sj1fMNqhzOwas9e7ExkI/lumuSkdxkx
AwGi8Y3Xvaiuo6GAjN2ID08M8t4312zsrrDnZGiDdrZu5AYpsRUmXSHU4JJ/iK9myV53NF4dKiZS
5Nuriy17hGx+ymyktGRyQHhp/EMqYidGua12xaRmAjlr65Rsl7MXp5V2UkXY2cdEZL28ETtsHTfJ
+nEI9cFsMDRFv/MDoRZ45Z6vR1qCyXu20Es9rxcUAzMI8GJclMrW2xGFHdo50FqusQv+nNPdmOpL
F2oRL/k7zrphrtOZfXxAVMa7PctfyHpKwaORlqRsvpvAcjq7yksWW+Gz2Rb8k1Y7Nbrszhv9NWxG
YiMYmM1jbcTlLQ83IdLZLghb1VSzI1Ji11QMKFFBinvb409F5KhmhVgmfAn2g0cM9hMODYty85l+
vugIcIDHWx+/Q2e2Tcn0MVl3iiHwim5x4Rm01Y51hxBzs+6ZqG4A1HHukWxPxdv+Ma29IcGTK4cP
0dBEKCcvle7lRDSofpjAIr+e8mcmeDrBQIuG1gdALmz2e4e871Bg9facUicjM4vSSLDzL30gkjZj
DS/h6++JKKE6Q9bB4ivABAmhv9GvL0eHp2toLCzyoHVIRki0sFz921ej+V573HCRQwFrYRXt8Bb3
M7A8fj/zgCLIv+xIC4BDT7HjxWc0zWUf4C1nU5FLK6X9cV03cv6GR0Jk+J/1QW1O5N8eayiD+mkw
2sw1ZRPfNPGpU2v+MyylwX79OF1Js18vGBcTISziPXr9NZ/Qjl0S0IiS/6Yr7qvYnE0WKTXjwA9q
3hEvS8JRYEOJHCxCQDFSu+pZ/m0pOeaDMJbpEnsA/ze5heWxBzCgpRuD/2wK5SVT5bG9mpgTMTfm
OKhB2huF2V2rXNx2bFiauXvZdvbZUolb2260B5FnZTorFmywNZZA9uJayB7ieV9Zvs02MGWvmbZD
kfqUmduyvsNhXav1t6gG77OKhns2WjDxuKPszNFQjdyfesQfwdjXekpb/PaNCBwwNfYa8qNlOnGH
8/2T9CWVQpFsT8IS0UhFH5DZXOkteWBBY1hvOs+AQIytxuep/3M8Pww+dpIGupPlqkqUA26DdntW
P4tfYeRUt7mj7MgP2zbYpJY1u5u7x4sUN98etMD3l/vThzrtO5j+7Cgr/AuQh9WloisTDr0jjL98
gNQg1AB4EKmM36oQmP7xs6VFnN7H5LCdKfNVMi0aQGtl7JrmnhOaSo7gkDu5OTRtLHLJ5yQAJp3E
5XSZ8EV6K30VIkBPE9Q3mwG5l48A3QRTptXRkwQRUPT11i0hYy+Gpj8L0wZS5sl4dqd8WArDqQV5
fsxCOSUwsfDb1NW1hMBQYB7HADxbJRmN7rwl5UozN/C2WSTceNFJfvJaLnbwS1otroEUAGAsH73J
5y56GO6orfdI2P6rchWVJtJQHwQcuhXHJQjYyg+q0RJTi0Ez8oGcvlIwcBCyADWxPDIJJM44gSbO
sriN9QjO16vZsVBOsWiXZgYwbcnvcA0Lm9hXlD6xAsUgwJSnxSk+vilIUCLQjtiOFeW3oxrRs98g
4A7eGDcHyezNqBQ+3anUFVNt1oXLqba3AATEGlEpe0QAlPgI9OrqxVb7wrs7s6uGT8YqTjpsx+gn
Ie0DbCyEG5ZJmNH2g6wUiFSzUlM03FLgJnn4w/TAt9mLeWnnvDXZD/O6tPhlVpm+anFU5THU6x+2
lK0aK09qEP6CM4JhmjMTesSjSIZV4iZVWxsJuYb1evbJQUxjym7jwC8SLv1O9WKPPnn+94C8qWjf
VFQI7+j941HivpULuQh5a/+V0ur2ZBwAG7jdPk2GVsgRcMtCWmA5qfeLq6Uj5S5ZMImOEfXjsqdl
EKyBCCwJBldtVrR2QGEzM5j4w86PjNBRfKE9o5OIyKgWZPtmLDzmC4cImm9rK2DKYE4kumrqE9VX
xAwcaeCVZ5T66Zth53ibEbrJyhApMat+mTK1zIR4pZU0JAWBqgtAnYeGOVhGMkIs0nBQxOK43DzB
sfwtnZGDS0Pq//vacvteCX9DaZ7PMdw6KBjv1sPHvKPjrItiXr0UXF32Nh0RftRAjdTLzqlEOugL
rk1BpHqQglM2axs8oF+8ThlNMCtKb80MUauEBP4mB2HNuC4w9DCR5/kG9OZBsF+SdVpdWk0aY8oZ
55WAwIqIn1ZV9309L2XposThqOh5S446FamHNEj/wR5jCZ+ba3zuf8GVhrSg9jaYmG8186Te/UzI
8KsxMSsvKnTvJ+1cdqxGX+2poI8zE1UB82wOfcvmZAo38tH/41ME/3xgbr3UIobUlxgLIXWD8Ke1
xk1RIPgxSG/FOMqQtKlLZgfrwSuclmN048yfrWNnyE85QoOQ+RRifLdJRkfd6LCtcET+sG5XAk8Y
D5q7kZozxDuE8iDlpCy1PXGXRWerNbMs+HXsJGFIh7QmCKSmnGQsbWyjdydIcAjhzRceiw5tQ3vo
oG9vXFGBnWkbuHtVDpXTzbkjXA0P4ew2z1ZcsUyhRYCfLwaYg+lhkDTSqXwvOPwO6YbddNRqZu+r
Ti3mBtoIZ4/g4z3/LP0teiUPcSg1etaQ1po2jv+vu4pP5nrRZXZogyVTMNG/6U6S/n5yhULa5K/U
UrVgoeaMPvuRWL4Bj4SIYK/rkOqKiZB2n9TUt2OjA4r2tSLOkwsG6IjXFkUFoMBVV52riR39/nvh
YeJ/shgBGUU3KEijOpA+Zp9T/oLO+RmghPeGJieWDiohRvIAEQwiDKMo0btqbiQFgFzfo6/TXTgU
RiUHNVQ1fOaLQTtfVGJIOzeYtaFunZxGFoROmeT3AD6uvAaDzH1W+ZQXRluI1XyPFBHxpBBhuFRn
WxG/QOMiuJK6IB0BYrO6LX+Wn2Bhs+tJFqChF/TuV2dCprxtLa0ZjNP8s7UTmtVVOt46zOqUa0Hz
IlSCa9kW3nbkkSbyJTsTyaG4ATxmfTF0VaUjw6vdXFRPhi2FAcC+MyUViDFKkTeiRraawJr0HIVI
mPXIVSQW2JJZ/gIryoARjr9+8dOOwWl+HEbdj+1QazDigSzktqp/HjUDOsPXnGSmNf1+zN68rsh3
DMlcwczWAbGCNGLyDGVqjeq+05x2BDZh4O3F/cRKNwMDs7+a0WRiv8+l6Y/i1LzopvKQcHJizxN1
C9iO8xsd0L2eVSAQXNyJOs990vL91+HsAc07z3XjiRfH6OBdE02aGr3A3TJzp18Fc1M1HtBwAnUg
SE3OPdQI0OX2lz84EevXMlyxNRO3nAowYyzJqGl6sfY8fj8PwcOkFMSAdNEXEDr4GXQryY9mD+Jb
MiG5wfTzWR/7c7i4LQMvy+SQ+BgqLKGG+tgEjriStWJyYG7EWFR4e9vfleHpGQWHLOe2rkOCFpC2
u66TcXJMA6vk0SYPxkxZaH87WaoOlRVuDdxRsJMAqQCme0q6Wd7GtsNiJVAhFBxxysbtouhs9CHt
huQh+tx+/mwGJPumSDTEp5GJYkLfpgJvjz4G1WnhbKggCUTYUZ0z1Lezpe8KgJSQhZfsvEMQ8hzb
mWoLwUa/LvAe4RMQ1/Bs83nE8nmvCsxbMqXemSNPn1aFihNEgWMuLESgjMX2NGEindNRoyJPi6D6
swUabs9ykfG1ZyvDR8sjZup+iylCFQEs+OpeIoDI7zCc+/smmlmgexnd5UfLLjcdDUte62TBeSCd
h+D9VJ9b1SKsjo21auRLZdNKNMUCm/wYsK7ZbYhDCyf+7LESDpSj+KGZ53KnIZu/DQ+FR8hqrn0i
pr5Un+fMGYKEeETquC38Krkhm2G5OBd+AvCoL7X8251qqrEIdpDOZW5F1eLfdCRKaSbjigBfsqxl
UxhXrzrZR3QLztT69rmzOUNyXsjkD4PdLL2RkttcErkfz+tVf2AYfVMAdcFFRBvUNiuz3Cb/NB9p
c3Qv3mPbzXrWKk+BuUn6OtP62opglAJam0FfQRVYKD/yAQxI7JhSkRPdEHHK3XUuYLl43AWadqsx
JU2ok308shU5igWGucCVRfYxdA0lm7JcsVLdXpwSDJyAU7sPnih+R+Om76FCMLTTW1rEJvW9a5WV
PVHxTV1qrMGzfP7a6i7x8JDl/R/5Z3QuR175u6l3WPxvg3Nb8cxBVrkn+xy6Ev+UUW/T6knYpdDu
8nYVF4momya1/rY5AMDt1M9BqOAe9hmqg3l+RZr5wMTWLnAX9WZmMzapuvN7HxfM3xfEWSf70nOA
HQkKT8ThVFi0J4VSCWkwy8tn6k9Y3La/JbGIbxgvDSACqmbqQRLa03mzs5uW2JM9pZxa6hK/zgfL
ZWIUUIkiqV1flB9VXy/CQ/Eo8qKy6DP6ZHtQJPmzgtO6XixYLCiH+ccn+2p43LAWXMfgEO3XNSS0
7R0/ImitFdJH3s+P0yP993J3+ojnLBSzzPxN/LCGVlkrQgJc+ZcWH3T65/pAeAlT1ZqRmTSdCuq9
4AfMsbUqMtGHG+QeDwmTGrMmlpxoNK2/Y5P1yxgJlWCmTgPvthrjXWNHsH7hge24dNkOZILJf9vK
Bd86CyZJuW8yT0jFSpfaBnmY6GiqCKguzuZr4kIJ2ouCpsBq48sisppbeulQO79K/YEjBSy8bbEr
qnIGEnOIeW2kEuIiOwkxJmiNtKzfVXkAMR3wOwtgJ5q8Hc4joPrjXKASizEQgtJ4qKFvgiAcy6Xd
YF/pOEIdCFVVk6uMwvwc1eiH5B068cNMHg/z6XCOhCGcb+TCr1yhRl5XuF7BnRrHpROi4C1qiuVi
Ma+pxWNGHW+YmAGrzAht2NSc09/7ADiZqnHNYuiKPcp4VLgjMis0ynqfmYhHWgQIsV/5CGEcX24j
JVhQn7kGdvUWNiMWR762Mk6eivhzFtqZSPUSDjlBqHgxY+EYsoRc4+vHJCMIlRapqN7quogX3qvS
iCuWvLXRIWV7hzrbH47ajdhaso4UyVX8HfNK1m+X9CkpVbtde1EaqyoikPqW4q3BsmxxIO1xR/JD
3R47O5IPVC79YEk1E+mnE0PLPNJOTF4hzHC3b83BYH+8nInGD2cVcfSZkOnayZ4wBBlru/yx1gbg
pPBRNBCRZIVwbu+vYlgsy/5sb4AwK4OOyjItV2yq8P1nJoTbhwVYRsoYw1VkXL+O9PJUELXkC4sy
axR1bGV9auHatfefSgdVFSDgmR5W/B3VUa+Kvy01YZa0bU72HbUOMt6v3V6eqRcrTodqYtka5+Im
c5zpzc2UvvNWaGmJ+jqhBg18r7R/hPVkjcSRjElflVzfrBmLwraRRIQtHRhlmpHBEAeiqeXGJ9pF
yfZ7msID6vFvLrba1prZJYBLq2+nkasq8dm+ZNw9d/l88+zDDeM+Mh7JUnSNr0hADQYR1baXs3Gb
lU+V6vgoM4f4faChoKe1bIDhRo1aY4R0y2D5lLcKPRTPCRuArUO5uWGpsSn04ejFCu3gnw8Yxtfo
Q7c4gSHaJnsyby++Mf7Jnqb1y80qjhTOeIRv4CEGnyY/eGUVZxAInZ1tulZBulwSnPK8iKCMnoDe
Z3CzwxX132fLr35tzdzkcJ3bMnc+boaDJk0cuYezUuSMHdf5VG7kauY8qG0W9D6Sn6DH5ovJgThb
+t0de09APwQ56sMN647qfajM8nQHmUj8Qfoj7Tv8bkI1JaRf3P56m4UhqFiyXjSkJ7nOfZYe2faY
2yMqyTx3bJMD64XHKW3Zv0sTGZNcumtBBFMhoho+/7P/27taQ+AS0U9aRxILBlQsSqvHp3jxmH5+
w7xXrJYlakUIZQK0HZXTgFietovXvVBx4TaExvzvpuqut7Bz6Ur0T+fkAIzy83mLY+HHiUkDzkmC
V1beO2MSUvLrfCspAf9eTTibMw/nQUubn9OUShFdtDWGqsFhNMs24kORaHEuy1hUV8XX8SqZtSKF
vFpWI7BnEgOLQYmz7pW1v73yl47Z4UPorD/BCPZXFhUKdaZK5sESVIOcgTESDn7Ys7U9mWTO8q+o
QB9J3mWCj8eWw0IoPqLgDI04aLJnYm2sAus8zQCPTbVAuR53qw/hm1896EDlbBlh+IdAa9BwJIGe
VtekIt5IVxPaVs5ZZGwFdAdexs8sfBLvEMFxH3OaX9f3+8BbCvp7GqpcYQ1yNljlPVxh5/jM0nGS
UiLIXi+vh/RnLZg/33Ea6whhg4IxwaXlpldbCf/dp5qcshSEfvJVJMnnjpvA7oTH+nUS/PcF6Y9U
or7qGV3ZujU00QXr/1YPMfBxCutFMtCYV7YkU9kqB2r8Zc954C68xUftFz6iePgAZqINjIFHrvjF
G6oN4qIYahl/iDioN4pOpSSLTZbtYfdpwskM28FSbX2gCGBUxFRjBOcV1tZFr44oxfJc0nApfZaA
e7MI/4ca9usts/S9H3qzOjIa0ttgJW7lBAUYRBTqxxVDGmCEnQiY5Dv6tSXKEa+oYR+N+vIZBefi
dESx9z7f3CC54nzHwSoDkJ+8VE1JxsMrQNGMpQlIyefaUdFpIkkmx/sfsKfkILnRpe1oqVt/YCeK
lVpEkOtt5knOmwH1SGeX124pAY5Lq7TAeugO4qC8J5gat4AoJ4r+srtEsss2OaqUQmpGriz1ztPh
etD5W5NH5OlRe25XKReRa1OY4F3bPscrsrXIVRjrsH2m3dCnim8UKZI41j7wTVx2tGLM85e0w92G
VfcP52QhhjRxvQmSU6rsQ19d2tovvYN01SQIfqddSn+yn1lFH5eDdgn9DRAoHrxgqFzPpq4WSEkJ
HiB05jfuyw9txLXRgEONgCNYkJDRew4zrVUro89BunFWNTH1f8kyLh3HqqsEAPk0/5kbuEOqqwx7
k2FmkPsBiKxr6wvCL6swRMr9gc1f0+ZBtavLLDwQ2LhDlGDIrf9debihmekYajbPeixjhDpYHJUv
yNh+gRH2QrLPFRB/gRyoThjePm0KC1El3XFELwj7c48b6aFFu0kQbSlWxNGdWkApYyegQwFXlNYP
OHWrnujF9l9U1jCDjMW3rny7VF4l6VfAXEMgOeskFz1ET3rUbXH0RVuE3Zj91jbAcxpXA/hweRle
A0raReIr+Xc5tosJmnw6Ap6bgKGvQqt0nj92g3GnNO7WVE/aLmWaTX2KkgrvNkE4huyo+uShSwDb
UPSBW4PRshCcMalcWBRm9rfFSWFxmX2YmvwCe2S/5wMsXrGaOijpmfBJE5R0Xt3tJN5xWBJRj9G9
f0kRYIdrkjZoEMihzIQUcbWmZrFDPN+ahiy7M+DnQUeItyvVshiefAX0nh9aW9eC1aKvwO5AoQ6x
yDRryuuxNLgkHICd+rpzee88ezV9pDVWppJP+fnBBryBQacIxBIPpWjkyF2kAWIwJtbh0O9QXc/A
89sPyy5qTKzSPbDNvCiZ+LJ1AZ1+3TPFlJfMYnymaNEvMVqhj0tIOHgCsinSHmRgv4/Cqr1iIrXE
Jy/zqzNw9/ZoByJLevzrO7BZXIBf0VxhJRv5p/XCugcaAmZNtZgTkp+mrV9nWkUNL78Kr4NYgoDi
GqH7ndHFU/zCAHrTWUYhfyuXnqQB2Wk7XzNOTjUz4QPFkcI/7noHB005X0JBdjhofEdMI0+oDcTW
ZsJ1GpIaDmRBqgjukib6gUKK9l+E24ALZcNgQtUTuh63K4dYwio4FwwmfbUU83KbiZncVdA7o7xL
YDFxuf7k8Bc+k4gNPz9gY+OblfZ3SYmUC1tICJVFhHDa27NBDwjmp8mVz9nc6qeU6vBPdm3DPmWu
Q7UzVEnYthPHuP/t6xyEO9UDpL8Eyzki8ZG9cnKh65BYkpg88kne+B+9ZbgWrb6q9htTlQEXTRNJ
vr1BPyrsXeW60HRWzEEhrIprLsxuKUAWAbcQt9AF3m3AgiwM3PStvxQ0XY3i2pd2dBePKhIUORbP
dOyAWN8js08ZxGOywOL/Cn4UeR7KUXn1gF3UrG5AKvOlSaU7yQoDZjkg7DHGAX6C918Oa688HaEo
rFcUZikBUp8dlA3U4M4iUXn7zIIf4fOrukVV7s/BD+C8JfTJjK/LKKxVdmkUbtyvTvZosfFyJOMj
xDnZrAPww12qKuXLlQ/UNg/ptrFLxCF3G0TmTxhmJfE2cFIfbOkRE1104Vtd0FSYQUuqf6zmApCA
cvN6iW1u61yjBc3LN6tTN6L7YD3kzNEucO89xTYZodkvJHG+Y7KwlnzcmwPMKuINpl7BCC67FJEh
owCn77AXA0oSoiO3pc2DJ/59iZPVHRiC67XNQHAB27ojV1tE5Sfpo7gvKnkLdf0otNrDFFkgV7b1
auDhysxJBaisaa8vHU5aqKjNSrrypjUtO5yt0GDcf47ARdGc0likL/QJkRG9vMvC/dVqEp9qAXJr
hE0xW1F4FstFysxoiQ/P1oG0HxIgEtb3wz49jPponUZicFEcrTb9Mkiyoi+vXESVe7LkyR7bvc6C
qIbA+8xOnVEaIkO3a210xu+Y2CoN0aX6BD2T/zOcAzfFn5s5A2SssdDtPxB/KHiw7k0tSa+XqpdJ
ytU9w17JHfa4fCLp/7fXn1ecZHzKA2r26YUDURCC2anRLGuTU6Ir5cWi/QKhjKFW8EpHC+gcmumE
CVMWtoQCU+kx5G/jnf25g6PLO3lygLVbxvbP4DLbpPCmWHGxVArlUo9sHtQtlmTt7zs2TpvBKGtW
5y3FRmNgD6PRKQ5Fr8FWo5HMoixclS9RxP0iARXhB90YxGl7QobfoCCklcxUUJMgAJ7+QBk+can6
8THCMmiwHVmUGg+rtXLhB/yvwCoXGhVdpxhLbzvc0DSTCOlXgn6yISf5ad4Rn40Wltk2VcplRHXJ
r4jyz8RdkFMKcvs9uEDA/+LSf9R2tqcyKTomum6eNYKIhMSJr8ohMpTz6qb2pe7qpDfL/zD352uf
EscGDsLXtXku3zJM2LydFc5fU7hZCv99pyc0LfWUcSY2rGmbIQutW5QlMCxrns7xJI8v4Dr8zcJN
cJkpGQTBUHSFpT2UlfT85I7fQCoLn5HFb0TQZMXemQ+bXJe+mbbAKR4A7YE9xXBcCSN0VFgXNE9b
oB6UCp4VsjA9lg//rkw4uxdOjePqyOcE8Qd3ZKiMQAiy2CAOgVxDmCpNu5Yheq1vBEnKpxBSaUjm
aQFLvJasgHmZZyqCveH9HOu1dbrLBZWNIazwBaAXLYvga5fGxgE2P/e6Y5zI1LdFvv/w1C/D0xK5
bCJmTKfzsA/1HHoft8iG9A8dMurxSLum1e5nho8hiUcmqJkNaOx30L4jq4JSOg5ItyVunooE3B5h
MY5zAeAaAPgJRo2QLkQaj0Cbm3j0MX5aKxK1bM0uXPYoTV9LasnL0pJuTrerFCoBDBTFRG9BD71Y
qvFtEyCdTXGPIGc71y7R6N2DLostA8JUcIBdopFh9NyiHOIrc12h4BzLI9PJqeVhoSoOOtlxOnOz
bCSX6WW++D3wEG5XlFeuEizE/bvAitBBxGjS/IUNKLOnqVI4Y6U2clWbi80Bjtn9GumbtcHuN8YM
vcyqvNLe4H/CLLCArK6x++TZlQJZyWyJ2HCp3NY/R9FEfKQ6iGabz5zKu/BNpnXWbSoSH5vzrcvG
yr2JnbHvAyp2iced73kOpb1ngqgxVJchEfSBQZcwRHnjZ1lF6yt1QKTweUjUgFgCdGYgYUpjfY8N
jVMNkWNrooI5hzUHBEOgIJaQagvKG+8tBee/tcEelO2zMnw8BMaVCNkfzRErO8BqGiLhM0cJcb+H
wQ5b4yAW/lBmeW/Lpijin0DNwRlnobJCXPLsyW7PRLZhXG9rZCugzP8wAJgaj07LMoqutlJVJF8p
SsUppaXZyQJ0AuhVKb01txDTb4Xzn1PXFwEvUiLV2uHyr+Al0Q3yGeULwUpfocHdPhCAIPo+cwUn
ppZuflCr5MOjfial15v2SK6REPla+2fOknZTdW4oM47Nqsu94PNTS2y2TDWSpM+grpiGEploGoYM
vhl3vDkhHmVxLeJjEij2V2DhSuWHdnydyAjY2nNZAMY5kSES8R0Dhl3fU/20UX+8m4fkothnq3SO
3MW6AqdgOeeBn0KDbyrF1o47hylLHannfHANZk3WIvyr86pCzSwdv/2HEbmL69kEdjFwQ54unOGF
o/R1zCHsDOLw0PdZT8ekg5kcgwykNqw+lTFCCC6Y4yw04q+Nj1oiQNid6UI7ANltlWxSaPyyHxLo
ri3mwAGRsv8Rmy3KPMAtkttoV6Qvaa9JUUE7Zue3mq4MMByPcLWoaS9KU4DoJQi25xHKExCCEyeu
FAuCCxwe/33Y8ZmPbYLCpRysO0t64xZnxKSmlOpnWVySO8idQakAlmmDnaMlmR6OE33tTJU99YDq
wS+B/o+W1BlyyJ97D3AMw8RbPY9bzvMhu8+XCM2hf7gTQI6JLzBv5KuZykHEAUf5DSctpPxeRZ2c
HRq3JuBoWKiqFE18PSaWyd4P+k9zjs74Fqjn+FlJKDUuL4ltZjNRV2ye+bKusLoUfzRw668CyVBu
R1035jdV3y7e2k/1EKoeTrVwQDu2KXp2pXlpUs6EssOCrCMcEhVHHIUZKc2bdxFskX1dxDigRo+X
dZO8ZmNoOnsaldKw1+HIgbkCjc9fHt4PT/AhsVSQafRzFjpJF4ZJyaRo8ObCeBDyi3j3Ws7hfMzD
U7Tkaw77exlrBdotHpWpYBfmrSIulCyT0Z9Vro8wUGAdkfuTCnZdvKX0OQ62DEvX8tmfqnk3ELxx
jL6XjM7Oh/ekdtiAcXIWOS21DP7ZpYyFSS07P1QeA7B5bs6+zcrv+Geip2LXBOc53rhOn5Rb9NcK
4mu+8etQWQ3eJdhJtL0G+psfUUedJZPTC2FLl6SefrwX8dENssdlHtSP2XR+uQRbqLTUk74wmSrw
7X8pYwNKBCyrWM5gspCnyrYF2OUmg3Db82nbBuXVSNb27vt5xxEjEzZk8QKwvwWtkbvycip7nNiD
+zLD4iUQvHq7vzGFN5YIKQmIoWYr5NblOpph2Xe3foZ2b2XJzMEX3bi1KaneZc6Q48SNPamGg9rY
sOYcFZMQF3/8y9N7KGMCa/VvR+EhcqnLwYYrEZ35ruENbon48he/RLBomG72PU4TTiUjYxLwTWor
qBMAACsE/qJ4HFEFOgRitGKOczW3KYjo5k4kjAhSQUHoqnfbWwtRQG0l1q+PUZh73dV93mINIKnh
Cr0kYd+VAzgbMQCSVD+cZZF1SgL70cUYiNsUcbcvm2wt7LauvrSKeAZ1CHPbXNqjLC9X4F0woBEP
Ziu6LnHDLTaevaNIE1zNfeTh56X4BkdzQb/LMy9xfTVdp7IuvpFEKn+hlrSbC6hcGq003MLoxbC5
CrEF2xzt9WmtHWoeqOrrvFxWy8sTtb+iCjiKeIovAHw3w1MgGo/Ee8GX5XFpLIDrHVy1b19PsUFL
K0NcsRg0HuzRlbu7EkNfzioGHPSPblFt9T0b+ai/KfzHrlCBQs25KfygaMD4aEtX5SD5RtvRzkiX
Op2jP1Epfa1SJjpJKW1c+yzApeAmojl10tXTmR9rTtO421w8+p7qQbn3/2OzwtdTl554B+lk32fb
ZhIynHPM5V6Wyq9R7Wa3s8DzZEf9Z1kYuzlpu6+oUYmob2pYx1oYqELy//h4yVBgRaC3svijyIbs
FC1OVQsdTRexlbTsG0yXtl7HkMqvn6CZ8/l5yotERu8pZ7stb+gLuHNjpGZRq/Cc3RU3OJBC8pnW
YLO6CK2bcFrVj7JVaeGTlGuxJzrtU7uA4g7p5/lcYU8Gind3qVfxlfdJJY639auC0Vz+Pr9RPyrL
CzoN9W7wt/aCx1f63+09sasPcEeNUXPMyrKtNhxQW9B7Nqjp226ys4RqCZmr47lYRLplSzJy5Al2
n/zmSl+mbSb6utZJV+202uSRHYRD7a3Ledpy3nx9xEJ0rMQn+BcUfXlnhIrI3DAdIbmr2y2MW++B
Sb/wXAxNqkmpK1j0HWXOK67hCdh9Sao9My7jRkTXFIVTM3hYEg8L5hZY+1ES0O24UKP2XhRDPtRo
VRke5mF15jVLpV6tXw+RpiKa28MiIdZ2QNyvVStG9EAS/nAxeiDbbnzebvBEAj9I4ArpZTpqsKWK
qU1QIvpKmY/ZLAKGcB/DlgZfCOKKbst/T69SYtEh3BgpKyZovacmB7Vp9aqGYr/FA7sXkwQaswLu
HUA55Bq2UNjdHX9pdHhLHwKrQ+Fuzii/NJyo+mTN2Vg9spgoAdIGpchptnb0tTO1uNgNkNIKLUCZ
QQC1Sin7AxDZM2SmuRuOg9c07Anv1X9SwyN30LUYc0MhKF/b3o1I9Yn2j8bRMjl5ZUI1BDfX28ey
iZPFa3MyFWxePhXCsc+5GsseSiFEmn9khUEl1Aeqt8d5QFzZSedwstK3fYMj0cVKDrT8QRNxJMKz
BkfwMk1eEiojeFn/VFDGzLKxL8BdGm0WsImjPfpnHoDYIkCEVE9uTekP2sfKkjxd/vMjDeS7Iwis
OiY7HR+7ohp1PjBkIbjmGEENgEoHvzXholXIraTBm4nbdj3Mj+EV5sRYvizgmGk+OX7IBTckWWR8
4T3eAr9AfrHd2RXxP/Nx99a2tNVhsYbEL+urNKNyvqmfCgMXCBGRm1T/19r8OeAXzWuW8GfjsMMr
2apidtQs8pKFHRqY+jb4cTSe8vjq8QDGK6YL0fEqjBH0pzl3CyDOUWxLfXXOirLUZRg3OtJJEiLl
v9iSJWGmqu+6yG+tuLNYFi4X5agEc/tB4uzktAvsdWtM+tqxy2mPzrTdoi0z+6nUVgBxRFg0Qji7
/6G9e06i+ytAQ3teHxe628zHpoFwT1tU3vO0kVWcvViY/OFLQ1WamoAmJZEEf4G9759IUUBdoNFT
hRQI5MinD6XeWSJUIVHrQtUtSi1zu/pX9hOOh5hZJAGIdlj5GQqU2XtyraKRKVmP/KEjb4Xp/wRA
BSDnVkS+wE/o44TXG162979mN7+GoHvPEHTBYq496PVcbCct1liVqSkMWkFjK08B57BJQLJu09Qu
IJuqLmsKyIMxd+WPkfyvWPT59GA4wMabVRucNtwwTkK25RgGIYsWki8kNQC8jSYAB48nCTnZs59A
W/oWV/qxY+tLxYkJn9oalQmFygDVR/EnoN0iY1RNqYeBTukEGdc+YYpkCKGveYBPXByUm/B2KQGc
Mka/b6DI5ilvrvr8AuUiiIA0WoM69TdelgVirjddWyTJH1m81pX0T/J6JIGsJgL7A+6Paob4VQG7
sEymv9sHYR4L8n/IeGg11m3pxE93uwYtVysjUQRPJTY4yYO1rR+6jjfuwJLZiPwq0zcXLfTTveiM
dxVcYvyDHW4qO03qM099RvY8jwBAVUvWJLkBq5sB8dyCxtRBXI1r8a8uG/aCjrpuluJSprOf5zWt
szTpqJCV5fUUpflvNhRVDm3FVcnZVWx/n/acGuONrDIxADWVz1rgPrv7l/0vEmRrvEb4g6ZngghK
MyGKvVjbwXdqB79cu9ExuvfASqZOFAH1UzDB1phLe7B1Y2P4mjgsMWDBkH+Yy2BkTh00o4J3V833
RcDRDPYIG0GmfFYpGBbRaHWGeCiLA3/wPwRsJb1clN25ZqVwL+yb0I2LGPFTeZlcN5ty0D7N3dJK
PE6rnBX1oe0cz98bJvupZ3oovrMZrjSvNUCO1p8oiDDXcDtF4Njjk+LXC7Eytap4XTTJ9yQ64xdJ
jjK6tpbdYgIT7iBLVBPDBwSW1nTO2InyeW6Ns5VTTw9LUl3q0WL4+19+vcmQWvV5ckK3eMFbs8oP
S4LI2Ea8I3gImAjYG7OdkKlAPC56E0N3wh/dTQ6niqa+hws4K7WwmimST/56+zSrfS8UbxfSq47E
V/M3RueJHc+tF2Pe05gcIVvQknb0zdXZ5mBUnFqO6AoS45ncz9tzU8ZMxQhB34O9dLTxV0K56D/A
c/wxYtBJws1A4O79vybA9Xpnt+sQ/XOXsZMmrmDZ+VuNpug9ZvgqnDw7UL1xB7CBFBR3UyqzMo4X
5RVHe/SSH5oxsOZ5oTgAd3wjdkWu3wPYnXYgc9SCJEqhQzxHJt4fj1xPccOdaFg9Lj8h9wLdNUgH
YG49M1cv12fW5/5G3qfz7zHJDSQB6BCzDRqE5WsC41a8w8y7C33JNPcjYOifBca+4AfWVme0l8rb
2yYfQE/dj3J+gA70blF1en27j+vnsLXbmLP5Fi5zhpi/K8z5KzYy3fnfoGlZdoJcs/+wuREj7XE4
iMubU9wLFh7h/yr+W8+1cRlxGp2YBKIRngL7e8RH46A7YoOtoXbLrAWaauSPBCG2IETwp0O4yNKi
wMVw6qGRlTvcDeRs/GNKsYCLUXg2ewY0twoqMN2Py1Fea+oYaCYIgtvjTYGPUtL/YVjRtxQjEyz7
P5k6uaUWy+mo8pOMQEgY4E9vuZxty/0zRMxOJvm7AzogzeQWMotthH6dPSfuIxb7xlSNyOhoryGR
xaCe9dEfq1QFKYeou1BpGpMjzpBH5h4NGglnvTmKrdFolPZMoXS88IabSYILR1EJujGSCY1Hgym0
fX4wc87WbySXAePz01fqu7cskrX58cPZKlF8SMouTpYjGkXsTTzuYKC0ufAJmkc50zsW9MSMl6SW
3CuJWjepzSP8MnStV5llmyk+/Tgw22I6UlG/Jz3AiAOq45IjckWck5kPw12oPpOPqBxFELK7jsgX
0jXbhzEedS1Ahl0A0HmRuAMinpAMOwf0v753wwtJxlY4qLgjlC0/7BHRzM+e0MWxopMAYpG4CpfU
etKAynIvIWsZjAh0CT3glta9k7O0ZbWhQcqjCrsKL4ntWcd8HuAfjuAA7VRdhYck3J3j1TjSNfIY
vtwZJNJMoNSrk15h7hBj2928cGPMc9FfkaYkwyIAS7rKoiav/6CrndidlRflk3o79ts3FI3OkM3i
mt3n65BNUwG9RIG5J1zEl6OFClMFbMAL7rWvZnGSfL4HcTJGjxkF8quizkojuS+QJBPuQEgkyRAv
AyzT6KV44RtzjmLKoBluHkDlCqtlRYNKSCPNiJpK5zQXrmT6QDNaJaYhoj/8oS71vfqGgaGeN2oY
PbRcxGY33kYjKKdX4eFmmAexu8Dild5x2QFpst4U8W6Sp/erMpkqilaMXQcJaguY1AElWYI8IEqL
4NveIRETnuJgc9F4k/LnoY8hFvAjp7uN9Jn2QzGsrmGiPethMHoekso/O8RbgAmFaE5alEE+7Gzs
eAvXaM7bu1kdAWk7K7sqttXIeYrF6dmXwXsVQRjRt1fcmKVjS5zyg7YSw9Oe+/6OXRBwiZhT3MiI
kVg+KFMBXfodjvLCBeMbEyhcv7bGNx6UcIT7nGA4eF76ciosUKmpdcPw8kwfIsvuz215aMIeGczc
tA8Py5f2JUzMKayR3EjmMa7BIopMr5K6QiI20DvfPQqswRluI2bwgNqMw3mKU2iCK+c6gO3jlvJR
s+HhZYlxFl4v/rKg1U5SmvuMPjzbPGHuh+G9rQZxjxhskhfPCFXyYt8nOOIfbR9Hp/eIYIFfj+kn
qwhNLhKJpdbX6vO+06/9SsE5xiO9UkLfVBV3qQl2tJCdzMGs8OiArZUbajSx58UtHdvUdD0j6T+f
3mXS0++7zwjXQ3Zn8/KNrWH+64k94I2DhyXdWGXbdY4fnvty2eX8sNIjS4y5zzqqh7MLv/CBW7nx
BsIKj49Nxuu0kk/hPhKlJDktDQ2jY3Gk0hmKw0WY6SNKv4Qh7cbVkQs8RUmObPA1yQ7LFdX6wsyC
cUxy5ysnlUtDeLOiVmCDO3aCILDxud19Pm9Q665IVEklrsHjNKsB6WqRrXYpRhU9Ja1j5jiMIreG
i+hvkYx7euX3/t/yh3SFMaaajhRcy7b7AWiUhJyg/CXQP03Dp78Aj4wwwdP91EcBNVLPGXD3yarX
jcpRLe/s0g/WQ1TQlgHGcx3Pjn2aPs0zgQPgpTAhcc2p4AU0PP7MSQOkhg7whnLdTUfbhg7lFpzY
w6ip38IT+fVpBmKPmW6YJha+Pv6DO8neUerHu+h8dPs9w4t6mu+4xwT8b8fNejAlNxzm62aTfwtk
NnMXFbKoQKPRD+fPS1TqeoeqDHtjujTY4c3/zEUHSBAkuQO8kgVKFFMHs4d77mV9U0jazFaMeIqi
RcM6PpKcH5mu5oD0zN5GZP9WMhnKcCzhUDxciRm30vQdRYLpofglfYT+lLr/LTbW1AJ5MTzW83zo
yxS1uDiUa4z4SVLyfyG0PaFKCe0zZ/uL7Ef6OIIbPzj0j7pDPZaRmMp0B3TlaSRR3CS7Y3eRDdFv
9q02oVqpytegNNhnEEXJ0sHILjL6JQMzVxW0WVuNFVamD0kh6f9u+NwucOA4+RmTrZ9uybT6kQhn
3nuAjebVslK/xdVv10ABRsNwGknYP0D6j1VC0Oevl70AbDSAsN/Hcg4sbPBwGqWa2xZXQAEWfEr+
DCTx3NOp2NdCjfvNScL+fKDRbKNbsVooJoV1m3jyrt6MGUJsOJ2Tin1TzjFxiaAnb8WFZIihacgW
ZfAvdtNKQKggH3+NyD6jqIWnNyb7k2kjLqrqeGTfSADYagFk2tcx3EgJj2Gyz+sop3hQEaRdpKU0
yi0IwfjG2Weh4Bz/btsvWnYVjSKUYZZian2wkfGL+6QDqQNmEuZtqOGMRx18FAwI0iykkp3ch+wX
C9D+kHPtoWHRTSSGZwoey/WJ5JhPFBgMDZyrV4Bi1ITDCZ93ph3xEI/xLLUn/Ig/zGjMhBLojQQO
moB9byk7LQQrJRiyrzWZB1urE22KHmCGSH2be4x3lYTnQKw/NUzoLOx6M7UQrT4urHHOyxlIc0D4
h44nB5q0ECxHPKh+fwdv2AvPRiDHTXiodB5WutiO4P+PDpowrVL8mk6ojtChc81DEIakstRv9H3K
HynhzC5RcYWjyj6/oNrA4SSelnUGL3g3c91Q3ejuzO3DJ5AgtMtxZrjY1KLRGx075LiAspQJ1kuW
vJm1fM5R8mlJXb2YeANa+/arf6qx/9w2y5T/Z6/TBZ2LHD99VPVwbK/vGK0cU3fclhytHw8moKq3
eYQlguSf+t5o6IbNTQfjS0ltRGdeH4zs5zYgWPNwA9kBvOI0MGe+Vfbtta98arSa/nkSphdvpEJ1
qCR8OLIeJZk0hLWL8Adpu80X5UHZpLip6Hup1tD4LdTo11InOTbLASu3bHamnN8NV23gk4xA/1g1
cGsqIkX7Q7DJViXebusXOMb5ps/Ayxg1wgUYS50UprYxGqLafDemBO9gy6V36bgJo0LpqMaMn4Nd
pm6ID1e2GYIO0KT7WzYq9WxbaU7SkDeAwuTRXvRNp9PJ049SHih1Pm/iAMit1vWm86TO896ikjut
TP4lMu6JuoSMxl0UZO7zAD6E2R30OnBoyCNAR6h8AEZ59//uZcGBnep2z0kH179NcLzC3TKGw9t2
zZJqyBf9n4ewV6XZ7wfOiXH4wWk85ErxRcMYS8phEfuuy08p8mtXQZomXBX3ffHuwAkmLxjWwdhF
x5zRDMktlbOeDAu4mH6dGU7I3E6STwwqwa4mVwAKaaTpOYOTbL/G1MCsDcD9Jado5zJrjGxx1xHV
8NZ4FFwX/zPKg69wOSdPfFhXFxjcprOcvU387Df8aC18vP2H/rEOUOn4KwxbNgIh7JwIk2pKLOnc
YEjUngPm7/2sFrxcAjok6jj2V5JjTX5gVveAEnmmbbJoAp/YqEWAAyQ+d1x40s4p7j8XkRD0r3Aj
a+MnSsTqspuPaIOEsR20i5uZYVDFzGt/g9oA16aY+FwzEnD14vOLmmkmmqt8655czud1pOf3Wtdi
d+YHK/rvZwkqzfdZ1jhluWJCe44WuCy/kzjy+5fc8agx3otx/4jR4/Xo5UlH0q53N2PmC8skCNC6
f4+ouyt5zSAYBp4hi/HplA2SjE+U8KqBsM6vqkBlCwjHxyiB22ZvrixcEar2L25PzYLpnpEP7wlN
fN0P8qd9LOgIB3QD6LX5o2TBha0DX3a+EFGTVMC3ZUphBjAXcZILfpPfWIaKHc0CGe7ttTS8mONr
BZBAhvih5AbVi/NH9L9o2/+Ob8A97jthhP+tvjlzCpz0uItnDnRx+9jRWrc0laMHnQ4NiaJ/J06w
u5qYuYzI+/F3rMKPLGhmrQqkVqVvBa1BflVJ4g+1UboU1NjtFovoFxeMDQSWwfJY7cm9Si9uIyHy
LPnAA3wKkW4j/QzJjsYOSZPJkf2VU82BUscOceMvnZ8s6aWxqhS8573Kewz9UC1pORWG+DBaDraD
NCtiOLnCojdLOGXun9BZqUfOk0M7XBPh9ez5uK7VbLP5zZs4cAGLXXMnLfffmpfYwGPlhk2qi6Gs
mjpkaxfOZlFt4hJ5E0f1LAfm6hBlmTA3GtEoBkc1voDSkbr0hZHDT2wyx0di6E3+utdnNIORkKYC
j6zMxyy1jyfSZ+pvzvFomLoAWtcmzFPvFrLYvUToxtb1LFmWC5H/NHDmH+yizm1iXqPaHfeXwlTD
yTkZM+jflV/85y6Lyoj8Fy4qKgfELke8tW988T6eWv9dn7LMyqhtWWimyJQ2EL1fIVurTuoYHALh
XBrNjjaDNX1kVg9supRkr+XU4ISMyMkP2tiLfZZD6EgWsHP7jKHo6YxsgJW2iaY7luV8E4w7bnKO
bwqp4s8FpWsWorsTkvIG6Ysq/gxsff3XKQ5DIXDvDwEveUmAbG2N+wFgokI3YvDbaSd8NJUDuZ85
DawOA7zmTXhSR4VHPBjYpqziAVJ8UjfOjlrp5ZOv5gEKf9HL/jCDFPJbAkkTl84nMezok6iyuE43
LxaCT6YMp+dbgOcXS2FcLXtUPxKE5h7YjwzURHsOivn8gxcu8BtxY5YTAgFDQiFpaYqAZku9/d5n
UEgybxsX/KBbnYz6NRhpsviKrgSjgBD9jOiRQ0mYDrfnaIZ9q/J4kEsbWxbLR9A5ul9R/GJQE+Qk
URezRlRdbhyR7ImxwXUsFnmmb0dH0LuzUmCQbT9OhuhH+jpBZBB0bqL52Z7huQ2lDx8WZxZzz0Yj
/UM1qIQuePTsL+yGMPlwSq9WZc+2KhrBeqaidTphZRPFEd8FyyfmljaQMb1+45b+XYrJeyGs+NVX
C4UyluAkIm7oT+qf/MQRHNUzQOPwC6P0c8A8btx0+bLV1+SCYnGyjg773ruHQXqcJzSg3FgWlkv9
N0i7qvKRYXTSnM4Ea0ffpgd+9t6ko2Kr3qcdF/fkDsQG3Xs/FIsoR3T88VdwjLaIJ3t+umPGmf7Y
I8DYZ5Ajj1EyAWKAkvpD6JDOZ/ijuFzunZJLz/htLQ7xNmInB4OKKJPmh1x2ZnbwOY5QNCaxZ1jQ
tS8iHY+8srax1yB0VabEiCP9t+XbL95c1AET5bjAP6scus4vTj0/IENU17LwGo3e2/rSX7RE7RQz
nmyGR/M0gIeRgrOLfL5PeKIOosSkRCs+l4aKOfqdqwyV643Uj/q2ETkNFIbDL6WrCnXUNEdrB40e
3D4NbsrIhxVxLfiqwqdtBeNxERW3Mw/YGCL9hCnfw3+aurE//0NTb6cyAqboXsGJxbT/lbUv3AuG
OjpBTwupl9vlydwMEvBHu7LQr5FWuCzVvK6P8ZtuYvY6RVeA4+8qETE+qwbmfVM3SXXPDvgWKSjI
kVDITmJC0c/FwihVPk4AaVUgaUKgh2TluvYRdvghDPwrGoDtTJyHekNZi5e6Pz4z7HY+4wQx9Mz2
KK0naTYfdHSBOJl1UDeKm9s4BZigukTG+sbgYMdguvWY+xoDS05lyE4KhGmfek/MJbodkaFexYNF
owcPb5HpYjlcDxH+o+K3r98dIISjVbvqb+QNsGM4OLbj+9V67TWOLcFU6ZlVTp9FyKWVQZvAxLw6
QgAs3LcHaV2cRPPqL4zv4/l1AyShuxskCcyBG17pqXZDKV47Dhk8eVpyP3Ps4IaLi84Y1aiv/pxa
g56rpjrh23nJuMgiTyZnKaFOv7ygk+HYWf8pRmiytJkE66iaDiNs+H9d1nM6mJJJFUpVYHkqo11D
88feV2Q4fEueK58c/UbfjAhRc/POa0VrFGh8RbEk+7kL6w11m+Ov8h3TBGV+o8WNY05wLxhBqQk5
/Go6sWpLg2EL1o2efzy81/8fnYsBHRk/7kgb5P2dzKPhfAoJWf/3L73DabaDhU6gDuEqukpe5PyL
OdZcZbRKGW9aLCab4seLSN3OH9Jc0Fz3Qt7gjAozD4Fd1dAzTCt7Cmmgmld87jCHWnR4Xv8bfIfp
2RbEz7+O8edXe9kXjPEGi1QBKYYgyQLcCT+Sz+sXXGtAF8Sfpg576ZVQP26PsKveL5iKeJdddmj2
HIRbmqoVPgFvwCSZV5NcRFs1A9edt1F+qQODxUh7QWLeWB7EXYlxGKaNllY6CalI/j3shUy98GjS
VIGTlMB9gdNSCE1AybjZKbCxPlAqOsyzpWKMSxuCwoKNfH//MMmmEn2nobTJer+AtXIQUZzz7ZG/
hEVv31ZZCfpJhJrwSdS1XM4vj9MnjPSyX9q5OlS62hY6uG/G+BfrXCrW9K175nGjubfMDod0ziPC
UwLkE+XXBbXPT5qz3pW6XqNUsH5q02B6RLvkoseRzbnqelhH/HXPvvM39Be4Pj8Hs5et7yfuxn1T
aFNRXYfjGvVuoXTe+zMTUXUM5LDX2S4RlIIZt75w0msqWjn5/T2yyP6gccXW1kiBg1TSFYUrdhjd
WQX18ZetthtayOVqxOOSrcwDJZePxJL7tIqUzSu7betuSUqI2e7+/vys7N7VWAnSpi6q/oyKO/Cx
h/WfEg4AA7+L8fQrKrYjslYf85qX69gJdXgh67PVl2UaaA9Vi2R7Id1f3wR/n+Y6QmSOqBd0J8TG
wT+nH00KSpPPndiUZm/1PK2JToIHZ51uA+9cYTQ7RtcMLkubJxgDbUr5oErlKIqF00CbUHsp1nZy
eBU+ustzAugL5lbn98M25eGdKu3sXeVgKrKSkx4kBbJ7s041YrGufdnidxzMyaQ3JvQljcOW3vuV
9zOz+BvXSyWLkHGR/aL/UQetXpnSZafQ8LM8ZDR/eQaWSQJ+wCeDTlJtYaJ7CQ//3Aggbup1W7P8
q8VKEYdtOetEBHfkhYEbK9QfnLjGEK2oJtwSFKqA4iVxLENR/IZSgzqccLSlbK0j3jayRROKCOlh
MufJehdyg3MvO+7O01JPhUPKDHg6zXYyy031t1ONdNuVTr9Z+LYFSNZ0JcFLK+YK5bW+vVg8Eodz
4U0Hj6jSw9/fusboQ8MfrnocIEiYKuPlVCu1mrkN41ZVLx7yrYlPS5NFbThwsgd4WLLe3XV12sYD
AzeKw0Fa+zSFAcb/pjotys1829AxDQxvqZle0ibBnXvtNiiSz6xs6bFYA637+T/r+sRG9R+lEE4k
T4CFlCc2wJ+HzdBGJYdPDLms1fxeC5nwFx+phCFp7OZOnjgv/BM+MCIQNk066JAfNZVnnFfyGl4W
b7pNw6T+ndwDd+16Zn1qztQv7iaGM11WtMdTC37+Ke/l+G+L6aNB4u/vATazKpDHQ6lYUmQdQAbl
MDZZJo3c6Q8lfXUZjgX1qSzPnsVuqFVplgz/PoW2Z3JMiLdJ/1Q139moOGxVHZsDurOj7VjBZmYt
ZjwZvpjhgzyNqHtvLWRijy8/nS2df6zbAB6bvEioSOEWvgaEtjAnRhgfsdu31t9t7PJdUsorWT5R
2MMYN3wBhRlj2zX+OKTUe3FIXDNTiqwoYAewVg1865fkRQcPVf584Kc4A0BgVbEeoFsv75vVGDLW
wdrFHI3lkH9NcAsmgQalXg4ha+rHtJozZ2TB0I+5vSjJZy12pbzHnZdbo7SPBvdQypRb9QaQM+jR
RXM1K4Dvtbqu5vvYWipJ2gtNUYr9WNYkHL/bFh4aQO+fWMnOYoj/M+McjkpjhXhhfaS/vn5PwUV3
a3obzHPywq7OcI4bmjgHpY0WI/9CRIsGHMNuhiYVW6eN+CA+yTVFPOfpJw3p/4cpSVUXRWL2NP/C
g5jYigzTrMjIL56fLN6qU9NBR5lT5BEQizmG3kagHN/7FDXGlsAMfZ+5OmGi7cNvPeaHRILY6m74
8EkxJKnJgYs5B+u61stjQ3nEwORRIDCrtCtB5X/lk6OdXVrnpmfhbKlprUdxW/2KpHjHajO9E+lb
fJ/WVwhckdMjmVH4rMy8IYuslRixw1THIY1iHGkfSAO9PGTsXeMtncBNs8bHOReMMeQOLbqWO5C+
wa+SB+Txz3pOn5tU7BGRK/RJbABQB+8ELfbcohkm76i+uAqm3hqmGFfpyK4LJ2bp189BFrV9JbKU
kq4R5CatjrPti5NpLIJvLb41AdN3ADuhIIXqgeIrii04LPPTvaE+fjIlgxzknm7cn8rVVyg1Wvxq
ZZsYiNDs3mkoS+pCacbXJKdgyTG6/46HeYDZkpeN1VzEyRsAcOSOEcGVSXFc8a6VL2zxmiG9Lxpy
Vkj4k5V0eGzlPmXsPqxbgIFHAYEWj+Lu4pt+GLNgu6zra4pWldZVfVMnD6ItLtnK7vc6EN1B6Wrj
OZ8LVOwSA8IM6hbpKV788DdveLvl5abJhz2TduuPGZwRu1fpxFx93uLHNNgT/M+KolwFT02sFodx
6Hc4aGCW38SKfSfwxU66zHA1ILZrxGVqocO3XSzBaNx+AUCEjCnYTAKERo4pSb3nPDNfoaIa3Vf+
MaKykkM6lV/FiKgQczJzCAJ9BvSYEU+oSvxzEfu+x5lKdq3h/JmvlaAXlea9JB/4wizavfadAecZ
GZsAzMJzrmEQpXVPoQcyPSYjGSWO2xXpgTK4X/imhUqs/Huy2XnbzrWFck70+26s5V5GL14Ciz+j
nq5DT1OP2EcTfMN/xzGMWr2ieHTAUNYH6VjC5YlLMN+69zHJ1t/cWFlbFCW7WGh+tldwfQdVzEhG
2muUBAeOrd0A3LyyLh/8XIdbPLcGlgVN+5Ot1J8g8WfRb+R6CrahKHL03Lx/EBjaiQ1Wv5pBIVbv
k21r9+pjbw2LKter2mby6+IEDQE+2jxiiOhMYhFn4MjkRXKPs/y+5t0WDFO/k/fgLxkoLc+ygmCB
iqoLiB8DGk3obMuSJqeLxUo0eHoCgbdk31LlsXfliuedFAuzMna8ldV0u92T3p0ugHFx8SN5QoWQ
PPLeRTS9I23v2kCfJ5KmN1JfaTMuleU83r9fhK03iNk+EVCeVGSJIr9XDEhg3l45UUtJwyF89C1+
gy5iFurc9wH5xW1TJLmYr/cn5r07aDIBTMHoHKaPbzJTakHKUAy4EL1SxCtP+7dSoz9P1rQjp3ju
IgU+6VNxWvaLdDCW8pH9QAIkyEb8i67Gk79PWgExvVTJDU4XQqq0D5aeeTEQJWZDnymt0+RcT0tB
5qif62dqGJL9HO/nQH5Ik5Z+0jQxc6Eh+jKn/2SQCJR9XvIuSyMDXdn5xVue4BZhDHVb81VozYU+
o+c0/N7DKpwmj3W/nVBd/yjLHc5wsjIgcBnCul23iZX35F9bodkQZUfgxw4J986HHGSN0E+Hmi1p
D9RnepYS6ISUnBBYC0gxZPO22N4+XYlsSQAuoO0oENawqkPGGICzFYtAIOmXyQTTPeOFff8shWUi
JvvkMdsRI5ejVfgkcj5buu9epp96ANjjjOzwJ9ghqA3tIv0oAS7wnPb9YxQmBlCbJ+yVIuLSc/z1
1FHCMLtCZ21F4bPwOZO2cY5sXAB+yXu9GMN+rN6nMN7VzpoMxz3F90RRt3x1cRMJxSkRIp2kRnkd
3ZvXJNCEYohKCD5GNQxx/X+JHQpMWzStCis09VJWTJaq2IUDcEeKR+zQytJEvXS1olg7bINGdesu
B2OPb/mGwJhQIx8QvnJoW9SQz+Hu+1HIHcOdmhPmIrV/2FdkYkgrZ3McGm9iHOU9WRRHpLmhsWya
WkL1aArBZ7cdFTuLoA7esJefEtC7FdHuA72Zq9LxI0fLEccjJarRYsSvxsNuxDufu7Wa8VshQbXW
tEXSIEXJ9q+1Y0L4h/nNMGxSwVKNY7dICmDXxwIdxYocixdAXSsh1uzYob1EgbcrwMpV0xvIYea9
raK543JfYDjUERRRFhgVyZccJa6dWs7y68wKu0N8KZ7ATrbWABAehT8hZOdU9PerOWl3A3nVZc01
txJD+j+4USEVjDjDl+ZVl7dGI3j3faH1WJCmGkkla4f3UWQfTkGu9lq1Lut3sMyOnRgmDXg0+njo
NLiqLj6So84XjGJl3DQitxgrMgcc86jwsKWFVTri5RYeRr/51Snbx5t5wAcZKLaFeN1bK2VMbNZC
VYsvqhKojhPXXxxjDJgyWhKL3lIjMO+X4qXcPxsV1mdI/unqwq1rGEeuWuMQWEM3P06o7qJCYNTj
30uPaEEjZFJ6RN2fWGAtnSXJvGPUqD1yROmU3Q2J4QChvmhSunp8hB6V0PG4s2k2LQy1goScincH
WtEjIaPWCK9JqerRGfRrC5ziow1lSA+KNd8a4QjprAoy4C04I3rP+Yt5ZlvZ9fky5gon5YX07TRW
8L68PWgTEJquz7LQxvIXfyHyj3aQylz88FVFX2l9+ll26ACpo4iMV19zKtF8LEOPPOd4UhAG/oSI
X3UBCKLXloYfCWpZLH238Rm6SwDY+6dtYvlkxYlAO8u1SI6A23P4wqypk3acQyUJ9K4azLVI0GUi
QiMxTUVdbwy8Cpf0S8Y6xZ9RlX+x4FTNFTNzxNc7BqqSKwWo/zUOjmp93KN6U2rwPZ3QmIoWggMx
Rw8uHjmMav6CoO8XjQyvoXhueJZxSIzF1CGIulLdl6LrJjlQqlcp2XWeg5GUe6GPNeJjqpMqmBfx
LeS2kD7iKxpiJq5KxfZnzlPCciahO7oAUEco4ffEjcX/aLbIOjz43xMcEvX+2W3fQLLcmhidc05v
7JnU9QsiCQjE7ZTKeP3z+I6nzOMdXrZCzAvrKxrHWc32iseZA9cyI0P/FFg8AeS3U21UUq364rB0
x5vJp2D7r01VdWZsVSgtJ1kv/M19xZx1GxTp6iKMeD82dOs8bNc7l5yFGzz53TLDiD+phgSE8GWs
pcAYXaYE5/6P4/5DQxDKYly/BYRVdtq7oUVm6LlY0w8H83VZM7xoMRyMq6CEt7tUBScHQhbtPyME
qU2SB0NNHe7xiPBxMPELZW3PJu7pytXhvDMoBhl8yoE2csdXuDcPHzYMTWXsaBuIXKEJpggf083E
c3NGetuxi8u3SqijOyWLn42dcUBQWLb+Zp+6NsiBlqZCJh1rkge8mKBecOBPF3QlyE5BN1eYtwSq
xjqjqaymeC9noTJwigIIunTO+QFbXTKWYSkeTGrVCzJSj4tlFtcXZSbzrF0bzehibROrbhywU/5z
tAErREBDlXbia2l28p41Dg42BQQtZjWOTkAJZYLv/JJ071pg/UvccDGOqzfsVfaYiWOSzQq+e/4N
1Vyh94DC2X43/jkOHimu2xW6pnrj4iUuNE+oX56fmieWEoHlZM0jGyt1dTRu23y/xOeL7fV25ZK8
+ax+3oKiY1YWZHy9Cmd8+mGLXzoSJwiSGiVTZZoXjzludaXL0fL1lQkHrHKavg6qIIC2PPCoZM2e
EMFUPMAuVJbtyVFzKutbhw7oRDrwnauxMD+WnSJsg46iwnmcqbjoYwV6hSo944rbbV0/StQ+ukN9
IUaGKHwb+al/22iPiTd8rGnAgoeD3P704ikmfFy59qfe1uGhc9pZ+Dvza2PQtv0uJfMybNUS5weN
rZTHowBsJwSgiaSmvzdjMgQKve+Ye6UdQi31VDLJaTUTnglXI9Fdb4TFtYhr796+VJKmsY2CcgZQ
Yh9Otfr9IiGfxuxbL8r8T9xAJkO2jA5DLmml4uvnnIWmRKy9xYBl8gGBJgdLA5OgUwvtgi7BZexq
5uCiyTlXxXMTSNzhNagDsl38iiEmV7R31XqpqCGfSl79qz/gO9qFCjvdVKv2sEj2jWA2LNVvippO
Z8iehVUeF1IGA2kJYMWQ6zRVRsfnZioMMB75uXGMblkhAliLaJ200kWh8FnAMnNnLYAkoaFdA/79
51QxaJ7fCXJOU0sleq9gvQFA4H20jxPPE2BaABipasBNU5Rz0GYYInK4hOxbgxltPNuXWPu5Ff9Q
1wXnUaCXz2NG/T5PT2+JcXz56P55EFp2jJRP7fz4jtn4aWamfkYV/sThqw6xlP/8lLj3jV2/ODOb
7gLze+EgEm3Vn7HymiSo5GuWew/I436WECbHQIG9stjKAoC7H4ix/To0LA/T4QcfPLw9bVoeZ56w
FzypZrhmKC2ZOnh8nFuornohXmYpgpfTILOD2iZquUkHRjpIgRl5jnUGFoqYL8t7/RqwOM4QblhJ
los9c1meYgaVDmi0IFuZ/xi0w5vXMPWGxcnvIZSBlmposdX8s/oQXNFAZ/bprkpPiTP3qFYhqpvM
xONfV/M6/7k+Jjbs+tsY/4ZtfneZeF1P+KoFHvonSOlkQLuBRHO4UxphPePGZAfxfRUMspSxQoYg
X1WJCqmVRv1TzyrOTmftEGMW05AY0vcT8wOsS5UN/76Z0bEXDxmxTLBSnYCWOsSDMQdnax8NPjP8
2XReWI5a/+d12Zl07Sg/CLkEpbA1t/z78OTABFWBQ0/VG0nLv631zitvEu8mt991SXV5aQVrT6Z8
Wudo6Pg4v7E90dZ28+1hpaDk/2arTVGofTgrfBnKEhWQ7WtWX2sxESdWpW+KCHbuCamphs0kcTvo
EBoNJbo7mW57uXiIaG/YljAy+M9ycdTh3GL14RGdLZ9EY2wC+bRVauHn/srXsSjLMyatvvPBLgjx
Fm+xcaGK/S8eD/KIJey0E2HXGUD7Wv0QQwBXHpQxCfePf+5Ogx1x6si9+7uPO3BN3kJ4mIZwBFyi
0GwdeKi8zhCyMTOCyy+yKC0z8Epe0So3x9b9HNhOXnEHUDkMC1ihyye2WOltKvsaXv7Ge5jH1lhG
VbnNHX9wY7DGxWMWOlRXVnXeL4fya62nNZumCBpVDBn6k+z25aSYKcmqxi354OT37kOC1DXusbDB
6O1xRdn2gNz6Pijef07L6zWBCqMdMTtFkVc7Of0sMbRMN++yFkVDAiUcxs9qQ0Y+9RUM7QnZ05o3
QGU4zItHRc+fXdH/xchXx/yypto7hux5eBfrBaAjzsZ6FecEAqPsQztjlQoPEGQOOYB6CJ0nG/F4
5ICHnlJzmqVWnCWbI+XfBjCgsjoSvcC/OvFBmQRXusPG1fNQxj4nan1HoRwEXKoWCo0hjykG2gTE
1BW2oLh7fnbR4E0QI0g30JYsbhzxrRG21xoMGoa52+RfVOiP62LHP4Whv9S7RADsYmQA28ZrlH2j
Q1SIQ6DDfUWg+6Q7ycS9ta0OqHVVzfk4aos8cxjZS4qZLJ+fswMBcPMokepwdi76/8bCx9NIHKTH
5Q1SCLHc04g3A/9+gAVOMmkJfc2k5x967Ekhd9MsTzCgwyant8XopVU9OyQKNczxUzqJbwRH+9U4
knMUSWcWbFagc1wXM1mw9KNc9iisoDd1H82Da0xePqLKYf1roN4N2BECGDMxdKFdJxFTbAkZnB77
TNTaNsucfYFHiRsBP5pQo3grijSU7727OmlwoJm0Lhlt8/gQh3VSuQ2N4dDPQ9sTmSJrfsN+IemN
qwvbSsnJKlG6zeDt9HqaR7VbSoQ1d4h6OOPZQBDldFq1CVbVHncx73jbn8q7zMiIVyq423BtSPBu
nDXAa/7mmi07TB4xA5B8+AxAQacxU0KwGDsHNhQmKo7ZhJP3ixRwR+/AeUewBMTkLadj04BCTlVG
ahP3t/Jbx2ml1JVUI9Xeb5PRDz7QAsi11fCR3qTTN4VUxLVSWhfTzUjj6EnKyGbxL4FTirPqT4La
eos5CbBsjc2F39pxDuWfexb0PEZ7Fxz0al0tXtn9CJnqwYXJSbFrMmN5D7kDHDBE6Dzg6dV7WEG9
0GmL8w/zekfCLkDg9zz4Wh6YlvJ3v8nbg2A9NlQJvTR/dkanWrK6LG9+T5cAxhpILMpMa44QpSSe
6wFbaUA7SVyfALYBT0v2W7DJ+RoBch105huPZosX61m+cn1h7ef5AMnOSkbWM6+6l6/z9y2wpoJ7
l/8ItHGm+plPEekE2Ggu9fonvRqngI5wbfe5jZ8elXzX2+0Bv0RDEfSNt3f+6BaF6oPehIq7FYEZ
t7JpoNob+muuoc/B9HWp8HLHQdlX3zt3k2ufw5fZPsQw173ZbGbgXnxF9+75cl876qMCWj41GSpn
3OjR0OTRXxGqyoQ4gnA1heTY7Q34chFLYbSMPr7jZvqTsypZAZ+/EmaKuRvJYthEg5Mp1CeQceng
LyqJ80J2eL7koZ5wQn9OWKbuA3SwN3Oynag8jib9hh20eCXKXS0TMOoc2Px+p10elD9ESRTEhctK
Jerij6iT6mdAIHz0auToFssSd+RFO0FbStSa4fLnqEEM2nfSAGa7vAnY9wghGz/2spfas4WqSxMy
a6DKhUwPF5rea1Uf/u3XsxKwKwIWPpE5l8U+vQRTUk5hh5nm6OJfm/CydP9oTfNjdKhksZyjcz4C
kg4VdJBheLtQujrE0UolXTZHq12l+7fYG6h7U+ut1g2P8gRU8j4Js1Yzyo30Ej7bYDdxl2kyhmIR
GHVzwMpDwq/RFPp1vucCzFgXHfsiWPv2LpdKSKMIYajHijof2W03qgVjfIHoYqqmXrnHq9ceZuRQ
iiemjvgfVWu5QrrzOd8nEfSosQW926Qcc9JiEzfI5jiAUZp47dzLPGw8dOIE+Z+bJK5ycb7S6ZlS
83TVeRXZMYlgqjor51Uxf8v5jzfghtKjmCmddsKh8FRD5f9U7ECRtp7waTUNFqsAvsYOlQOgRQ4r
hbOL9056EbtTGi8MNTV+OKSx7x8vZ7fNroqHCaJO8L+pN5gCi19f0hL8o3ViWdMlhhxOjLTzZg/x
1YrzK1DAVwQ+XU7F8sRcbiSU6mOxwmN7Rrd+ZkYW0X3bl58iNY9bx/d/41DROgQMMgRNC47A458f
43rXiDhGwNLyOSo3LgtenhyqN+0u7Rwmai3FpIQviEYpyBEgx0KvlWMhKfL5QsvpgcbpJC3dAzP3
a+KfzkT+wrAjUGEG3qvlmzjyUGfZAZuxZ49GT/sI3GsnWmH9xMRHxZKm01lzR6wQzSCFsM8+HfrH
4UxWxtXIWtT74wPzcAnK8cjAAPdeekCXm5dwYHAih6lv1LJ5TOO6U8lEmMtW8RnkE7lDk2QpmPoK
9rcMQPPj2KNg1I4bSLzAziz9v8zrsvhKLHKJL0jRPbOxaEfc8XR/p6t90c934EiYxPRj+iEanpVW
Zji4d/OUZf6qdkrVUSkFXWkVg94DVH94Q5uuXgOdlvOYYfHBeRfCuP/owMmEoKK12j1WVj8lx7g2
5D6xuQKub/gb/7gOWAhnVpx4BYSByuSn0lnHl7ma/kVVbP4nXnbmSRnomghp5ULD7KV4UZrA5GzC
3BPFlneu5LEpW4KUOJqFaIbFebmAYr69WZK0wA6BMJ8hJC6ktYxVNUqjVZ78PNIxSwmYrykRVmDI
OUdUCMmk9psteVciSbADLJiiIH7ThL3NHkAKaPojce4nj+BAScHtcnhFsxo/qDviMIYqug5whOEJ
Bied71Dn5kJvBa4Bz6eB/r0WgRlbCAVE8FmKKMq3EJwzRB8zniTy55jYFAN7jodt95eQno2K751o
nPHPEAonxPf2NF7Ru8m2XiiL/ngBXjmfyDdeBCrwX6TcW1x5VY5azRifdIWfMijgweoIB7YlDs/u
GAUHK1fGG0sZTXSY9hPxY8sl6DX+xs2EiERO0R6EEIiFjN7MCWWL5RBmAdOhxz/dDOwqwSya2Way
9+zpfaXtIBv8lGqSKWToSjDkCChaggrDLfT/3Zu853pRkyO6EnH+P54XpYUpV59TLR9g2vS+sAhL
R4oEnbWIUNuj41GmC/7lJom3e2XoNG+nI/GuXEQeuFc3gjZHE6vv1HFRnKdKfPeL5n6qe+KDMPTh
EQdu8kQHaJtXgGX4Sa4r5bc8lW8VD69TNBP8AJcwfouxIrXS29tbX1G2NrkY6hbfQwncXPHC0QAV
dGxs64Nfl/ffMEWnnk4jCT87PJGeeIb9zaUZqoQ+5YLXszvaRxgsXBgpuHaXCA1bpThwvOKZFGSw
n6O5kp5B0354yjwiyw6r+EBI+557MvTzkjeQg7dRm6OmP9/uvUPdOm/25QvgbTzN74Bl41mSEBHB
ls8eTE5mHPSbBVIs7QMHAFSiSjJnotpQiANscVHDidiBYp7rMxaZ18rIpfleTQFFZTWa5HImwh9d
I5wnugLDI413XmTOltr50KTqAI9eEWyXKhLfZCHbHt6u9dxxEqtL6WKLTZbDeIKq/3Pyg5Ab6Miy
lp7V1uIrKWIs7d+mSfe/2OFu1rR1Gov9PAx3ajYHuqPli80myatWmeGfulwoCZ6kDH3nlmEVBVz/
WtC/4c0OkQKPYkGSyOlpd0fFsVII8CkGiM1XKlah4Zl1YMdQbHYs4K+GvDOt/grS+viCtfzVv++B
UPh/JBDB+VK4VKi1qM463298ZMLbpFtCq4++IKNa5EEPLaIihA9y/ZRrNzNWVkQsLcDIOzspxJ2+
naIuA9aqlTwHradR4zq4Tug0WQGMjwYsGnTxq1MfjYw2nUL0Yjh0pq1ra1V9k6HcjDWvJPuDac9k
CROPcZXPjk35S1GNPcRAMjIr4kLyGQQg2pHPWzTWOeY3CTmC5OrmWIdJvXaWveWROFIZM886YI6F
FLO5KHOvHC6RUdYc52hWASXyxKsjmyxSwhOsuZJ77pZjqaGiWcEJ/f8gcm31D/uTyNkhxiM30pyh
c098cQQGtqG/cxcmCInBM4MUUan8+hnmwtolcL1yX8wF17Yzr7RU+Zc3OVr1WWdENP1rWdn+CAA5
C9wCNhaYWI5roudmx4CVvDqoHWFYi0pS9qs23JIvzXFT9jU8Whl16zg7a8CNKwAB4d9Q2hofFx+M
0Ce7CCzA6t+qxBMj1i+BrTd2KWrttR2PzC4M2Ueb3ARewwbPySeEIDV1RdLbQLfY+sFHal1XBwG0
wTJVEZnThQdm21C4xCDlrNbK9qD4EA/jTRynFu/fMGPoWVELnSMWTGDW3/LphrghdOKs/gLkcxJj
VCWWUJ5EDG8zg/VmzPWXVrbZcsKETs7Qbbl2HDuQCQS6BmtjyRpDz60tO8RSK7ZZxSuQKWlDOsrN
dtOWkjfuhtz3VLAqRwZWNH3XRXkuc/AEoLtXiGxA62HOBrNDq7m8EwpbfauvoxHQcpdEkzy3QXH1
dvx6HzXfcGZaWWDJ1kVvU7hxNaRRDUuHqDvRw8WRlZtC2NddJY2Q4YlEcPEjRLWj4CtAzYki+EXs
CNVMGFybBwbkmCqmjOeRS40xSYrk27eim9/C5JbEWS5YMgbgS73RU2XWhY4wEWnlWWwFDht3orGt
T6iw9KkubbqSXwEzmWnZnttrMBppFI04PV6cc0gZ4NTMB9vqW7vY9X6diCjEaqXfchhTBBG+OCig
JVGkSCPSmXCP0RfT3qgo1XZK/YE0YcRFzOfo2ASih/ggTScAxSrKoHklHXObd064kUwfGSVzqmMM
3tWHxA5tJFoK149ux7OrFS6L7B+G76qyzggZx8MQAjnIHcGeirUd64HajRJXRNZwXBbZGHQNhacE
WjLqNryQy7IZkbO9qHQY5buNZgucgN695cuk8BSeeOTrs8zKiX6+gKO0FTXjsbFtfCRjt0B0f64Y
Em1i0PcjDX43HUsTmXRUmo5Gfq8I+kR+ZZaeyWf7tdxW/zFVaAoIPMRmrZqahBZssSvgIML9pdGN
ltfSqh83b8R+o4Rx3vCTj2TzZ4DsvXJ5fUsw8mYpwu6YKabYzUIM5kiIdI4ueUYKy0tGDxehp87M
qe7ZcpDp/SrwgT86gMWxxJbS1xRLfJWfhbhQL46FYVNGW7OoceTaRc7J5bfsXnu1V6WJV8mPO/BP
whhka/g424TYjs2LH+x/E8fOY+RJXIq5UB47yHwKyutddhf2EDJavENF7kmum/4cd4lxGIDa/7qB
Y3t/TuFrupCrrJt16E7WPcK+Ars2z0AwC0sIZDhIdw5wBg+LtwUoi0OsmWrrYQgUH++d8vZ/MDEN
SgmA9/V5TyHMEcl/xgptmQYNaq04DMwYexx6S75RrNnh9esKu+T0+XzhL5FjSRMS3JElthxdn5Bd
C8Fjsi+RHHnUqPYRCa9IqOjSGCW1EnTEZI9zw6fsez0CLvfsW/VFi+YzMQfIyvMFkc9r1GQDq8I3
gX0S1JDmI+lKgf/9lW+PAkL/W3sP3smBacId5PVZ71DVO44fJg3KlunjHZHHg18YgXNAe+pVHEZp
4FGuf9wlWqTxu2kVOPJDFQVSJuOoroF8r3WpWmc9yHS1GpNKlA3rQUvGjLTM36TOsC6Qtr+0c8VS
by2Mv6d+Z6ocoAySNsDyO2L/USgzdgDMyKzFi6tvHGu64viz7mjbpYS1iyiocusNFcXurgPpJelp
Rm+pYupUs35D2ifxTuP7wam81zRxxVJRkVtm89cmL3o1aLB2ZfUyrKAFie2JkMzqdU8+fJcBZcIw
pQgsWeJWXHuCzj7CI8Pm53KKpxaVizjmtM1BBTlABomhSGmYtQ3hqNsfX4xV9iGNs2IkIuliCmYF
68mhFv2Dc3uBwzrlXv0bznM2+40k2yH36ghYi8Heh25K3u2S0nYtEm+Bdg9X9xgdee5soN03AKfb
efl7LZQHSf1rLYL+24MQoWrOZ/Cg22+l8TfV71gGl8xHMzES2kcoj9ZAA+S22vMmBiGmpqdGPZ4S
Z6caS8AB1+A8ejFMGhE6Jxsoq8gUUaPzia9xplBqcDJWqp5ADSKo6ke+iFdTXDTuAi0nxWrgdAmT
bgXOroZDzhmlk7LekIxPAub1bLUybvY+9lbsJcGgODPgarfjr082oY9MyQkVBab53zIcP006/5CF
DWIu64VBR+BfA5u5MW9gPfisjjpXzn03Wh9S7qHHYFglaI5v4TJRtDFRuZxRzPHX68nrSNa55QNt
GEC5nHesWO3KMCxGw6qhuYm7O66LVmChs+v6gt6PneXk1l2EQQjatJtJLswkY//fwZIFWh0hCmIH
5swKHg8rmpMEsEXrGfMvjzrq0NoMH8xZuggroPrfmXJoAQyZ/7Q7JWPR3aU4D22AiMITTsxI7x1j
GLdDJtKeTKbS8YTbfFSeuvlGZMTFQZB9NQ8nemYlHWO29ugIFGI0BWRfvnhplCREgvl+Xm0mPGGr
B1m13A1AGjhE1+WZXzCLfOpEo3rYYp3SKl1xCeWa5mB5OePrxhsoimSeJUO2iV61Q/rCPdYnqsHQ
MVZA9IKcaJUZASHYbRPQCs0rdXWDyqReu/z1KHRKe1g+JMisf2RQyS6LKbNyDPyvX+yrLKCj3+BL
3hW7pc7qW2TEI+EzDmtTjc2vwTI0HP33Qn2YH8tPJu9TpYP15PaHHfTAHoSm/SifxkHNeUXaH0q6
91KANB9QZ6fVznSkMRQsIyYIFshFnjKcXXtZB2qlZ7bl5nosHKh1M2WGiS6sPlLkwlxrKV/ZXInv
rxLQ0Yb9jHcNjUSjsboON1BEuDr7wpUAxkme8yfKEyP/I3J5NwqnT7qCueYUsrX+cduxU+ZoOp3j
z2xXbbUQZD1hFA2fBHIY5QIyRiBykiD0P3G7uVhhBjP/0zQsOPdnyj/q7S/xc8sFs3RCgGZNo0Tx
HQHEiezmxzqWkJmKXH3FbsyidWwMsFxZW/XJWW7h35puT3Apdej4541+6rKVyIel4jrl0o+jUS6l
IiEsAui5mnsgxITOoI9IBXjIKN94qA3z+QPavPH2V/FMdJrWcvQUPHlMfbJnHeqmGH8RDDkEFgJ0
lhGw1rVnV0zZ07yErBmtlkwY8ytiEnQ7uhyhmCPQvX5MzhZxabT2PV/rcxXSo6xWfDmifkPQ2Um2
b7W99ci2smanAkV5wXo50VeQubgQdxt2keV8nUkqz0xqTl3/6Qvcl/IjNgFdOvssG/cosP5cBfMd
f32kbbl/opwePBeQO+uNfc+7UQocsqB1B1krP+BCCCzAf7wD7RaJLlsakVbNirwpCucHmp6w6/WI
IhvX+HNleG97mYIQUuMoxp64TUbUXv3jfhUO5o4Zw+PdxlExzWlKC72V54YpqObCUfnSOs7A3ofr
OruBlGYKeWrxh8/LKHOo7Iin0QPfa7AmtmBzwavnVShCxX9OZGSbpdQAlC53d1tKl/kphug1t13p
HqOaibaG9zMzTLSvg8U0o3XlqmtmYrkTmOZG7cmcuJHHym1orIusNoycR9stRm03wc4RUn0LHL/b
yrKsMWaG04fTggp5e5kMPLhSUHMOLkLUE3xyqVlI6cK2cCij0DFZmfPaTT+LhLwvjfqz23CV7Y54
j7K2V1IzimERRx/9e5Ngl4LIj5YQ+uUn28wBcXKMdMbk1w8bLNzaNIbOEvTSzvXgQ0147eB3axei
yKgs+thgc3mnd1m22Ixka94M7MqHShRd4iZ2q1BbrvKyInyC3CFvjp8pDO5V6BvlyF5BMExQoiCP
y0cTZVYaSt7yKl7zygE73YjpA7ZiiOYNLt+HgMFMF86VyMMpsw2ZGL0nmSaPF44vPaDXIKLdisYG
/3H+AUh0HT0bTMP/su9HofWxhevkJNjpah0K3uDiN9pjL5hGT7BQK/VJ+SLoWYeqgG3levmNlPfZ
h61+5vek9f0LBgzNYOckbZOC2KF8Tx7yBXQzU80DHqec1vBjxl/oPXGwpC7wJuFq9aabx7qk6/QQ
gYe/rXIk3i40qUj01jgIaSv+7VwSPQExZY2NgXrCIW+bJ2xYH43x540y+FeEw1iJJYQ7f4rDNHl2
k1Rpyq5OtSQEtj/lsbReGRhA+12eZLfqbj4I8GpHx1SH/ACwUJrFcR2pwXs+2hY8dPGbXS1MQomX
+q+jcqnRVz1XyA+Q4zRIZkzpTwl3CjQIcAgUc3/9UdJHu3UW5EVTe3fBKaWkSAx3+ay6G5n/Fwkj
8dnub6f7kGKmByZBng3knLNyiokesVvORl8B9RqQI0lcSSfc1HSojsj7zJIG8Eu/aw0LECNvMqGY
yjSQ+OHLAbfV8VL2C/puWcPvSbyDLc5gmcbPNMqEdkalArwwSyyXwkEd30Le3AFvUMA+CSe3bAXd
H3xXMncdRvdzJ8M0jKMB+wCUeycgdSFLnvn/Pa6aYXLpsxyh66t2uLZHDwqpNqsSHCVx0RlW70lN
RV2l07e1ZSqLTfuon77o3mExd6RS3m8BMX9Vlvr3eFZKOvcGUXX7dLPw06BHTTlo5W5QkLGZV/Nj
0CoY3uZJw8RZ0gOsIlVyzmj4Sgr+dRoYY8dDxL3WqOGM5hpuaRsfc2d+KQVi/Z3WFSbS2jLIEkjl
va0Pgk1C8/o8uJXq/wVUR3gquF23rISMOHKG7mkYzmmfmegpr8VFwuAKIDBVYsL/CBPXemNFEkL3
o5CCGb1gn4MCheaNrzANrfX9W/xsVpp8+vyZ2XfZQBefCnsm/cKgqfu/zHtf/VTJbVN3eP68krZF
v6z6qzsans9Y7fUdjl0MorYwptRm3ClZLz0OSqhbmx12tUGXv81CXTIJm/Hq/QQ0ELtnop549pJ7
5CP/YXinRV4pU0OpzyuA0q2BolxBPzK0GuXLTv5pPI25LgJFOVK5VHDgBYFAeACwEkeMoHWGQhCM
DZDQ/9WOLEwUWw4AeT26SGPVT7AC/sqT0k35k/OtvZ2mkHZ6vyGEQMBSeXEPkiPPjbNK1yAmCqZh
3eqh8QswaFGYan0peqaq0UzrX89Hvs7nQ60zsAEEjAc1hPp3JdxKv+13vrv0Vbj2nrehObT6p3c/
2KJsu9T6gKDPTtx33jY/Tk7txpJhtmu7bYejDrK7R7FsEKyMD+RBRf2QpochZEXpzxDLLoSUpCop
Y7kocJew57yndE7dBOFhzAt1LNOK+RKrCGQjZ2185GqC3tUFnJdAGokIPo7uKOi/wZzjy46V+1pw
gKlDA/xLD2+5pQxdoh9oS5BcLga0rddDppo3ytmRUiGT632zrLTaTetn/p+xiwUNlkuY6d0HKw0G
x1zDvyJpVQrqttRUKO3cWVQRZxrFMxgXk91afK2SOxteM7vkBnGPhGOkVNedxoKq129JdQt//Kbv
IQ96cS+nCOOzGRl6dIpikaaJzL/5zsinkbVTzGVBEQurg8d89Whqg3ZAsBrtyR3OZ5lJwZ3RtUqV
fzJNkh7Tdi78HqdB3j/oHto+o4jpxtaCA0zRdD44vMoWCbz9aGa+PJ8uvk6gYIDFfTxq4RWvY/k4
eYRFCmeNqXIJkg3WrwATV/2xb+jiiWLVEySKk7ssUUMdr3TNYJblV66nxf/Dz6HOJiYaKkiQGS1x
qjRQebHRdyB8WQKShWndy9dKy5OevJzsn7Ekme/EdwgA4KQXqWZKFA9E1RjSt7ocUUjP8/yJK6du
+866TLc10NMCNeXZ9Qp545HvM5RnFVKjB3uKk/NjhRNR2T3bRMVIn8gWvrLzDfpyyK2hwMTUWCB2
GcB7XZOsUsCnD3jtYXwtF2xmQ3X+NGvJ+eau5jxFCDQzqY0tvRm/EPkWR9bgJsPSkP9zLy0j8PZP
/vUGXuoutw0XsZdt2p98ewn5u2EzDRPHOWvA5UvsBuDcHbCO4jYQSSf+ZW/NKWP6c3FFNXpsP6ha
ASsJqSpgOtPQoOYjmvNup/NjvAi/DafY1dqmSCRqBnHk4nU8rq0bI8CRqRd1UHYDJyqWlfAlv2wK
MWW0s1ufgPv9QruzsgypCs5gO4/hIne0hTGoncIc4/aM59LPykJU5cm3mCjlOn+yMe0fURHLcc75
ueHPOB1xir5AwlsO9xbUOgGhWIt3EQWJPLjPQxGfiHBhij4ijsU1/Jv05WVroHQ6Y0HX9XCDI2LF
8Gd+7Gwj94LyOFohXetBBsQc6Ke+jzx0H9PlBEO7meAP6WlxsGoR5P3yeO4Odzw/XkpglJGD1QL7
LShE1Hu7HtW6GbZsqBzy5hn8is0OTiPLgITvPeR1KM5wr7glhp7ofwXunxkf30cddQv5pa1Sta9p
NkFLuRGcZRSzE7PanaJubstqrdLsdzbrrbR/O97rIAsg3oR1BJ2BKRs4NLf3FZ0i3zyP8811TXw0
xtRGg53/E1aMLwxqG4KcoHfH3LHeO+rJw+simtkNeRcEWS4kbt0XNU73Q78hbkFwqcKoPuHD1uvc
4OMZZUWV6HdYv11mqLef/VBBfUYmvOekCZFwRpl7NgEk4/NN+xQw3RXBfUK3StekhQgSjHgbY6Ji
geIoUT2H81VWVlxLAlHUOJuBdCHHdIhqln4RpZbLPL3Kqsn0q0QbpY6j3qeVLb10XL3HrrZ2CKWc
OeiFDxsyi+fKLlcqPxpRTfKCUlf7O++DLQfaV1Ya//VCyQl8jMEyo1k58Fue8Ee+XVDvRk8hhH65
GeRVVO8wpWFjCGropOzsBCHH59UQhiKzFQjwzVkfEMxDBH8BSm0GDzHlhMaxU9Htp9OMuSc7LHM0
Avv9uv1x3OavIPYXUD2DOrGvQWy/xAZIOCcQp9KLxmS5pxnFYIBw4knzOJk/NtT5yL3Snyh+QzGl
wlyyiuTL4Dl0dEiS8HfQKp8ITSnyKLK5g6LOoLrGo56rjCuhCptNG/EkALoTu+bl54xk7tmy+7wp
k5voIwYm0/P5qV7ZziUQsI02FKoo85nvMLUT4hOsuCnB/PWWc1p4vYm/8FZZnd+M2bU4xzdXJeSc
eDBSMlJ/r917+Pwf9fUmWGtC++od3NVXakkvjMmLuF3BH1VIyDJbBqZ54CrzRu9h8OCcfPQkzBcU
m8EFT2lj0XpB5mnJrpry0J4GrUYrBce7VIetSPMi3t9xNaD/a8MGc9qUjPgHLiH5HypM8X/Z0hJD
VlZ1xBgkMKJLNmHdpeueGbehwN75XG8soQ9GRIuCO4JLFh06yWOoRak643uoNPP1T0C8R3+m/ukY
vI9iCNAZViVp4H8mBIIxCMhx3cj7S0ID+cfVlpWrNNAQiY13ESzGoWLkL754NiTsHFV7HHE2oZuT
FaBwEc8Z1X5pWnl4y9TR3QhJQFcfMtpW8FUjz53m1SUoA8eaSTfgAZmEAun4ArDMAkrhZ3f0wslm
ArzjgnSExORKiS/qR1OxGLVFr+lF5tRRke6dydaeB9jRWTD1s1NOV3YFsTNwAZketT7xtfMrS7wO
eDAfd2FG8gQsa+uPUMnrNbAXMoA0LJsW3+qDpEwE0d/DpYzsyBv2syWrm4mAILTg0iAb8OyLO0Xg
JkDjd68mNBqoHQbRDCcuekxAG4o6VdkutDbP97OIr6Nr+98y9DjgP8zgufLy6E2vGRM/QIAW8s52
D0W3ixYGGbs3uXoPuDK6grQl4ZHT8hSjcpfcW0Dk0+2nKdoN+eBKO8Nha33diypMxcHfqjnUqwpY
IeOa4rL/KvnYlMakcB+UZzGrynWPMfowR2Sw/j6eVvT6Xe27TBcU+poaOHHPE7BwG0fpoMfElVBH
7jCptjaAsav1+HvI7Q027UWBq9NK7SJbKmMmYR6iVjF5tgdPYKqEXtwgN5gCzYiAmTtWm1HTFX26
DYKYIJeUZRP4p627n5UnPA/ufjrstEPcGRae0DeGEY4BMSu75eolSnn+BjtSbw2xk5OYQnszKUww
UhQRe/ZZlkuxq7dSmToaR/LUfadRy50xkkSCA6WLwmiyIsAGXChkMtNzMo/ftb0HVBr6jr81lf6+
6jeOP/x+uwS2XKLbvB9fWw77IZJgJ2ObQT+rUveqF1i1K0ha4kY41jOfiz0SKgr+kCEP85RxZNpo
L56MXtfXTs1idYdyHGkyKiKe4EoBrO9z/NIrssM31B00mplC/M7KznXblR6RPoLFkFBbF73g0RnV
c3KYuGciyMnxUdthi/k0PBqFHzCwedc+H1qu9nhVpt3zt7/+Ruep+QmYJtWSp697KXoEXVXsZr97
PflyMzIEqmQYlwFTtvp7sK/YoYpe1Tc/6vtyevFborfrGfcC75PArDxxOLAVTRYZ8CfMNNJRDnjG
MBhgKikewZ9d973m5GJLDNEkLSsXAKgG7Ym30du8GJ9qgC57tErMnyvJzkhChMI19DGzGQyASHUb
2XbkjoUu5VLoGTNtK53HrDtFLJv08kKpasp85bGeAh0CfOmduQsmqLb3dqbqye0vmEjJtsJkwDQm
Le68drQ3GF1Fd4tK2MD9so1VgNKOQ+kVnnggzG8RUUs/SPmMJJjY4UYpbnXx0x23IWNNig8DFEPO
aE0fUAk2jag9/8+jKEZRFKE6jjJ1KsU+FJjvofaJ2yCdSM3ese9tNKBuxawixI/Q/Omhgj6ypjpH
mOnOO+Y4nGnFmYWNc6hsvgNCeiR2eNZcSlkd4bmeqa9KTVJC3N44lh5VQBtaJh3IWxwrutaLT7tn
w4etNrR/NogPWKh2ZQiBH7UEsZmTVVd4y98na9E2zOX2KBWqlW0CkGsm+wH6kPnxuLgKVP4jZptj
7n1ExWXZadKRd29+nmHNbb6Mev4K1f49Maaf1NrHBjoJdeUtuGlyNnDclj5N5PxEyeT9AYoT/1PM
eKwzMnsu51WT8DwumQVFktkd3JzdX0uiDP4E+LuVoLutX2FU+CA7JzOTq77SXkxl4B5tXKACY+gx
ouPEccJtCLru5vFQrnKpgN/HnDSBwxFiFU6R/sQXHWpCmhFq+vHBMBkaUv7yyrc81UoGo6F4tQKJ
iOPNZ5FFvO2AnwCCkPiZiaiFV7k91dOFZsytMxVPUN5p0jiDUOJHq5Ap8BPGWvwRF5O1c/ximfgh
XASBoQvBgd93Sds8xvrIw8NKeWDfEKK5rxvVAnMTUq6O162rmRgXy0btey6wRPPWTSJ85hJCSRCJ
NisK/m4LLhSpd3AQjXUXevxBEpL1H07YfsnsEB++3g6s7WX8hw0NCpcHmR444wvZ1Siq8wac7hWT
bzH9QIYsQWXAWeX/qJxRRoZ7C/UC/SMsqCaJje4gz5m0zOqS8N2Dw1DikjUiSA/a8erpIOcL877j
SBNh5e5h7ru1CpzQvK7q6QuTBKexIivmI3zJnxTCHmcDZWb3r9zYJ+V9ycAlOHkfGX9UMQOL+507
z0NydoTi1gxPMVsRHqUvrDZkfz91bHTBEQ95IHbCKfknBWIldmq1yr2yXLnQwloMgZoem70nXnWe
1Q/glgR1yIqzvBXJHxqq0Z5CmKoVBKqbSFa1ToXYQeZE4tYY58HMnW0Qiv6JlNC/rm8bLuh1kMyI
jAzHKFlGuHjonynLJ36LFnD4pcwHyaCuo9Ecufk5NllNtUsjbzLc7UcDSkE2H2RD/gpGuWjQs9WQ
q3eC49q3nvpw1PBVLI2N9vCiwfOXnUpJUHRf/lbTXJZfCftvGdPrebiuWwps2aEdVHr8Kyc27t+Z
N0Wr1AMhDqrPa5p9fTxLOpItvWRtNAsPTcjHWnxzf66d5CYA9g6/4sOyOp7w4N+yRQEM+ZBIv8kK
IA/f3yU1gmc6ek5xJq2N1tVVanLw8yetyqEg5WNKtilE3/kR1kE+bD12mMDzt+ysmeffKhhGMI4g
TdkYII2F0rjmjnufe5/7xuNGCdnqb/LJiHoq24/f+GB2HI1TpCu0O9sDRd0KZ0whu7Pc7ARuQofJ
YQ2AQsFU6BbUhyual550HRtZ+9aBx+VNpWlqJTc16ADM1EQ2v/DNXDxEd9nbKzeujfN2+13mgSY+
Qf0fxpx+i8HPp4U6pmg600VDqaN7KmrMBuV/ltgT9vFOrAsEKUvCIFcVMUGYDSJGRwB0QnDkpf2u
3eukNB/amBZ3ONKL+NoB5b9Az6h5X4Xb3TrVA5njA7JQeQuvglc8fd8d5YHq4ecPYQDaRmNfVFN/
vdgO6gJmt+SI8uaNl0THEIggR8RMSrX0fozY0LegHXnhNAaunoxmjquid7fQ60Rym6sy1DoZQ/uJ
nCaTxCZWFi/0RvFIQqafcLZblzEKpIGVA+eKY5mrxJj+zOToYpjdc/Q2X9in+dMktoNpYgJh08Mu
UeF3bc3Eyg8gsjubPbPkGq0yJ1eajZXAmz2EX8aqV1r2mGnks8qFUFwgwhnx4vdg/oz+Dq5w///k
K+Y0dAnUVEGvuuMslsaD5j4Wnq1AntgB/nNfxgty1A7qAQK++2JZfEARwDYV7yXn0BRvGDnQNw69
Ymm3N82b/yutSrNQOAhFlFPJxP2wc7IacXS7Osn3IN9gjaiH3y7VNNrPRyZYkuXqGgoUcw1st65y
RV00jkT39jz3C1kaGFDTfgTEXThT9KDQfUBvtXLiEdQBbg4zUKuLGnrtIOB5ZqbU9SN9Nlpk3La5
qDhJGuhHzlvsKx9oS+suIKvXuo9gqwN2bLWYuKN4XV24Kan2+Uud1wZkGi73P6QFN9LbQGX8HbxJ
bFFUmZDj5yGYrd5+ZZC9nc7LfkRL0VySkPxSv/8HGPZNMm1XsZOYqun7dsimv8SouEGU97rEGYJC
PjedOERoHp69nYzfIVtALmfr+kbpj7431pfytBefIR+VCG2im09FTeYEKws5gVi8JMNiMzrdGiom
k3Gw1Q90leo89xBpmHQBwmOvuAU+S6M9bVkikDDXhPGCF0751UUR91SlSnUJMaXYbqwJ5arJO7qH
synT9+Wi9ydDmbNP7iXvYXZX7i1tzz2yRVvUJKq8lanvDL4TM52YPtgyAvnXvrpCCVLBzVX1z01Z
iGwf6WZNY3mQIInaeknAPnaLkvRCUPnBo3H+Fd6umxeGO+amn3qhOicus3aPbUYkivNR/OCQmftm
rvJ7uu8pf25jkPhFB96nV+dBz71YDwJfJ0JLqFI3+ZrbM9HFEqGtwnSMPRmmtv4o++a17A8VGnhS
Y7NdxTarytstX3qw5QGB3mJ+KbYpB7R4qG7Xh9ltuIvvCuzbtyfR4g15DRgGk3I5EELTw7alMaFS
N1kjVYi/7fiKaiWCBrmkhfT8mL+xbclHV+U/V/mUXEDAoi/PEdxkRRGCquJbRy42LUuH1knw/kN+
2bHuc3HyH3yze8jyu6m5xXRfHvRVlSfvIUq2Act/YHabJgVEM0n5yXUD/83EtW6vqp+GL+2SeE7d
Ae+Xr6mA0OVsGkwoqWjjUo8HdmevWngoU8BEvF3slcCbZH1VMbNn5k+xhvgCas38olLbU5Dxo4oL
g7+EF3irhF/QLRWZHOpqLVdxR1AyPQCJxMZCWDh0OOkFafjQCNGBtx3VWVNv9nOvNki7bOVaE2Wl
33A8AhyCuqN0nAj2CHgNe4XQWWcJ/Twa7j28qGlOeX+WXdtukm3I51eqzXUCNDyarCKW2g9V9zhC
hRksQPyB90Lt9MKn66SpTdMhaqzjWzRdyCw+NEEhLl3iHN+vU+HJEqsJiBJ7RzNqPTXMdqneeh0K
O/uEqE3p/wD5j0aAqJmhu4btPZjnX726QJbdPTF0g/Uu4mV6n+EUbk3OZhBbQ5VZquKwAI/lAcCV
DJgY882004smR1ZHCONd+kRRyiLTUktVNc8axsNjmIaQ96RDqLsY+grWyD3ULOBk5XB/Z6CHa0ja
KG7GiKvUnuWrgc4xoMM+AOAJsr2wxxXppBjtKf4CzcSOrK9AEXxaUNUB/JwgjwSctApisPDLYP7m
88D0wmtukA6paQzmTGQpOAvhjzEViEq3uyz9tFToRKHJSsDgO+W1Zbpndtwn5AJcwSa2WtCuuVCw
8Lofcz1gv6X4Zs/3LchdF9+SJv0NvTTq06ex5GCGXj7XPglSA+wcg4jaQBk/u0v5EvJiNwmdgDny
4isqaVTMaDoaeIs8snAlQr9Pm3bV3ycr2g8AyIKX2tGQY8YkeQuvXFUnn6Kry11jY1GSyMpKcsfp
g3orB/whqZIgpBu8i5zfhHbI8OuthgTqOl77/K4Pti89qS9lwLxP6dJnqDuH6OtoIHj0rzdqP2Eb
9KBIYoLDuohhA5cr/vo+iqi1UXVW9KB71dTpbl5jm2ZnY6GtMVP9GUjBq51soiNvWRL3eTQ1pYiB
lu45fRVABdTp3krJvlf9ZWYvcwEMKNDmJdG0nzj48eTDZkFmeHHrn+iUJxT0+s9aGxWbCtn75Xff
fJErXiNYFBAfr8l9S1NjPVge7HtZfYi+EUWvRnnB+JkhtPoBWRMElG2Ti4CboGJVzj1+97ZgP+3c
GEJ4KG30sclGkS/yZjv5Zr3MFIxPvFvB+pgZ+WeF17IAfnJZLIschV/dJFG/b8sMr77EPC/2C7rP
6RR8CxciZnbCNFMyFiqe+21Yj/XTPuqyINAlOjttfu6x3j1FEcNij8SJfwFHnWB4eTDiHUsGJ6YH
KKlNYuGq4si+uAgUddEHY9DReX/GcHhZm/F3iv5SfOeipqlXgkCWulDqUNqsSJ90n9NYxbfDY80C
B0y6/bQw2gD5qbyMSXpMyfT0i3cQwQyZYfUCo6hFQUPOJMxbcfq1YiTkV9Rw3PvZDEvp/DZdC22+
I6vRzMURAj/a1yNENGSdpeDbguoPicEcZoL0oacmMi83eJc2h/GkW+t8TG8+z52s0oW8tg00xOeT
5fClugVXR7XyzREBRu/Fh5aeb1v6FIB6uAT93iC9Gr7t9sLOvW9kokx1kyR/B85ieGQtWre1l9yO
w5k0GlhtZa4QFbE6g88MVfvrbV/uXQDZUpXjMzOTfSu8bDKCQckagojP8ofJFQ9mmVyrYtvfirCD
50JMxwjY9dwufc4PuxHYz1DHETyo7sWQUXAmHx81VRw1GM/wxA35czcCWBoX79JvDkozK5bKS6aI
lQUJ7WUc4+1gQyHoP2Pi9PVvTtQwE1L4Dy5C8NrTA/XZkkzGpjyxY/019JAhXkvO6qSwf3UYZ274
GpB8lJXmW1Nju45EAU6fvBGaVYfGK2/Jn8UQfA7yOjMZs1IYEo2ZrT13sF8Hsgp1O7qT0SzKv+Hh
ECwLoVLr8578UdVxCi/twe++DfPQGuCY9mBFmwJfCM/OPqm9E2CaoY1TtVbmdTR1FO/0hv+LOe/6
91u2eCoWkW8LDv73tGu/Yf9xuf6BVXjKKXGWjb5rlzgIxeaB1Ewi7Az4ZfOfpDtlELyth1KOrpnx
IorbZWLZ38JWAm/QPoR/BxzZKszxNVtCfUsoLpWEJ6Z+Ja1W7YCvStLYYdymdc4sxNFcLteqqN9v
R+WHYngebMc9rJpQLd5qRbgL50bF9N9uTfuLQoQbA21838QYGvwPzWPbHePcM57rz/9GC4GZLaxo
U1NrmnsDTYRVUBSj5w3klr99tRE+2zIvQFVCUmSgYjl2J8lIFBzfeCqBh/G7F7hXOEr/S44piQtr
OhDbCH/b0geKjtTO9ICPETOrJ/q1uXpJBUocV7svC2lUrc6Lv7QrDBIr5CVvb4KDKXYczMFcXeLn
0WUZgaTL5rHWPKMPPSt4HZh2MYUMt9hjKVJr33ONdmx3FjvFTe/jmvqmMr7c4TsWIJJNPGzfIOgz
GBYQHsEC13M4WRmtki3kXEQQHrlkdjqqVDYI4zlGe4CZwXE+sF74R8zosl4BBRcQ8O8ZuAiEfAul
w0hA5gwqn3+sDxeRFNJohfGWQNC2szhEfHzvoUg6RVWQcsnFKva2oHPDjpsnwi4M8MDfVbwxKcuY
gWGIirQMJtpDaC6oWOXr2YBnp1shjhUAmQ0zY55oM8QPyo7vFa44pZQ4fdXt92f8QMbcxDlUx2Mq
nPC+sv0k3qNuUKzbw5bZC70eoclDrJic94yPvlUgtrWCQWSolJcc0E0mI9GY7J5RrMRa4EihrvtA
xB7wrpmQX+sHvRdL1m4FFPpj27Nsu4yX1Y4nvfU+H3uenBxrG9yGH4OmuThiMEnPC0C6nuHLbZDU
EDyIhO1PG3kZXOxN+6iHG2Aggh4o9WkZUhpY+0nDMjn+JAQs74jxNBOqiXZ1fNQyC8lgKQgWLfgo
bleo1iA+yc670WsSAuZf1dTgXEo46tV0BWdRBALOQBJWlilYyxQr/PGhlDH04RlmNBDKIpb7DXWD
5ZT7Ds7WxTI7X6Vn98o7utmsuTba0rYSUaKNSzoL9BM+I8fw6EL/EYV6pbvMhb1QZj6/xQX0lYJ6
W/EbN06xTJEmf1aLWAAsrRDe/920bTiu2Irf91tlguf+kLsb4YAwMveIW1NbnoUjF4dOQj2cshRG
yP83k3M7dg9GfkO+KDsyQ/koMOlA0iIE5PIX24f/c1vjUB5uQuKL0vI/hrmYnDeRKuKxjumkGVzA
g/9bC9OCP8OxHo6XKRtU6Z3zLsFbUmZofH904nXi3y2kLz0VIzydqT/s7RtopOBzG+1tSZ6bEg3w
Xvgt41cyDEzlW/N9GrYioR20XY/2uqdoRue2cag/jDjaiZ85z2IzfL8EJjp4jpGAVwkuFq8dHoNT
KtR47yh+ltCFrlvjBhCA96IsaPw8kk4GL851uLTYn2GCMom83kENkbdBia6227Zhhpn+r7Rdg88l
Zj1UqCyeVwEorjs4PfX45uICBfCl1Eht4oHdYlEGKSVFLmVI9FsPapeonABKuB6209SmVIzoGCyO
p/2vbXFFfnW0kDfMsBQxz32gYmmyQnk0N0SpzL2JZsp3p/+5riXsAK0H/GN8LoIXuRlMeg7GNOHJ
MsXPNN7qiAz8Lz4V/5XbF8j16Pm8B1CfDsUf66hF6IZH7WQSxAYqkC1eT/IrZ62jHa9vVKDpCqyC
PwKd0IhgETpoGLulictPIxRy4ToTJA6cpXM71c4OLmh6UYN2GBry56P76Q46R38t+zet+t51Ij8L
dyy6kl03EGKiOPB8a1xT7CvaVQra2qR/xOXhYMaMIH71UyWukZWdPDOhvknRA2jqkVPx06+HgMu5
CcBO+Tsidj6bISogxoM3/qIX12RLaS272Pi4NKVcsAg7NW7CH3prQKbt2Wk79Pgmgx37Z+eejHoV
PkJYls8t+A60FZjBBsEn486lPz2dlM3ecQ9RnlSXT3S5K4VUP9+8WDUeg5Bba2HmGZp7vnfPy27u
a4OuekCAAzYxXMMLr4pYBLc85gWGx+vFgR4OvGzoxpBFFNXYYgd7XMrPHGVXKONiTaD5MoSCU3T3
FLT3KHkYvbiydo+LxWq9DtBIeRYEGpFwgMLbYApAkLWUGDcGdshUucWyThB5PiyIsIBqGHmaFbd6
60rD/A3qTtQuc8JMQANpeibx2ylypEq9hD4SPFYexmZHXBLH8WrhDPF7yZPzfYnjVXklpPvU7lZx
dxum1FpH0p4Z/m8qnbz+MP9O3x1aXZ828JY4NaJdbg/UXnkZnRuG51vXVV90VqC40nOj5jnEbCR3
nxX798fH8ScEoYtMER96v/tfuXnWKsEEyBOOX6pEGTvlkAhrvwvYNoUo8+ks05kGOScjeLiSPvPH
GypF3ER3aqJ+GqahX9TiCo+ODktbpkUldCRtk6IFBs4OAGtzEqmTG3wIO6MBNh3SyWPNlbhjZ/cZ
afgWKIvlBnPT1yBNsmFt1honegm/TE7QE/6/sUjclY4iqMoFBsGEybBMSrn6pHT0hUCcQNdN/dzp
FBC+OVFgkkRKJXHqshVbXfL4VJOmNg1moJhKTCalDuRDWsSqgB8TDoKQFqbpgTsv4Mbs7znzRXp9
BfIn7IqeILFJ/xbrbDOE1KDULmoNTVTMBP9/BQ4UpQd0iPGz1JoV4buB/7dZ8LY3JogqEos0X/15
T7qFrxhlMYZQUnZ2pYo1lFFLTYxrWqfqXglkYuPszZP/33/IApOPC4yIQcn4i6L/tgCFMaVrrsAU
N2TgmRm74paVu91vByPBiqR1afx1PJ3DmtlDHcDAsuNbcawdGAdjOt5W8JEtdboQyZe6qcuwHbqC
Ix2w4JzZ3XjLQHvgjxeRrY4oXlnAG3wZrslvJYn9uZVU1BL0U789ebR9snJT3pIW07Gi5vOk5EID
4S7gsfaAyYowftkGnRQIc2jByloO7eMr9J9hINcbVT1ohkbnYGcf4ougebhd1HnbT7Cn0cs8g+6L
x2fq+buvGgi1lren14S5lKlQDEZDNfrcSJdIhj/IqWP1NmoVx0srNRfirTQaNNDCtIGnpwn/ONjU
9vHVIWf8/yWTs8jYvZvhLKkq6ntb0r+njZTkaE86/K/oo+b7p9DEF1B19rzZ3kDxI/wGK/DAebXd
lR3TSO5ExY3o7Kxy58BArIz/4I3i5DnGzmAu9V/ugLroPaVZRMjqwD6oSBkf2HnNZA0cuEMJ0cC0
vjDDra15gcPNgIBOWcUebdKusDwFtRj3+QxpvgrUZG7gMZraAFXXcJb0Wm8FulqIlGpkiD6LxIY1
CjDLUGcnsGlin5T4HD5oUDqAdNHMwNNKf45fHR863WzxUgUiaRgQrLXFecQFWC0cx2dmOWjZ/9Pr
bqU7rxAO35Gpu2JJtPzv2WB2h6n0n1LOz8zZfKl/uC+zBOxJ7IT3rg1sgnCOWUZiJSxy7/PpzQqY
Dc3V9J2Bhsr+6ciS/ivKrGXNDhya3ul2N4XKlUNwF9nuNr/lCg0X1KWWnPPX4Vme/W+W1VcpSViS
6pYELAjPjw4z7DkM05ouXH+b9EwhjAPoTLXM1VoUu9GYmKeyZ2YPrhxYBz0f8r8EHOKuT8YNg487
TwwLc/uLCasqRz8XoQNxOrBd6KubMlfYmOplP+oR4z3YminooVuvaW9EkExnsOcnQ4Gk+/ts2YQP
d8pK5/nc0968MZzujN4iRaXtFQGelb3Drc0oVkbhz/s+WJ3iK4idsSwSt3wSNggc1umZ6lA0JWyB
nsKH3XF3Dz/gBYGfDNQphusApccdqweP5yG7plRGnzgAPCvaLlY7SHpnLUZ9dJrBoQPI3FnxPQIn
IuSlZgDPW/NMX6VVcOEdqrmWOjwJEzN7CRamSYz6eBRg3xuyJL1YlLVANFmR3V53UQ7eJTtMuRPM
3TGdGSB2RDPanpudngl5usSwNITPICZ7p80HjQfizzVoK8CN/zG6BPY7aJBRu0FZGsn/FQPOYZw+
5dkMMcNCLIX6KeblJQySnETf1FyVA/iwNNuKULBE/ek/uXQ6Mm9UYS0IXxLDpXEMegz4cEz1M2wZ
hsm9GUUpHBxZSeZLFZLw/QFFubgRYi6B4/OQkv4za+fxsAvQPSMVOyoblqc2+QxW+q74iPZw864f
YMFJKfgRM8ZEBc1+m0q3+iSIFbG8U0bTBfSo8pirbSOMS77jJHfCC0Y9rH5Ck5FHaDp7Mphy/7hl
4oZJ3EWP9ClSsYF3hZSEz76bwpaLLC1cGoQRMO+QbpGbbxY+rX73G1ZJUcYrxshfT1WMfMqHRscd
0mflTnUy/R5MN0LHzG/RJ6WYmedC9uXvscBPIIvLVmgESXQymYR7Gc9dOiAflYxcP4BZqiuRspDn
7SfQeMrJ5WyZiU7Qm2MHHCBkNDOo0mATcTId7QtB2S05bMZER5ssnwPqQQveYKZiEylkNfZG6gpf
KIrSdFDWoXMGrMt6FJoTNq2XAw7jDy/gnn6jaZOI9LuQhcYid7T7gE4dWLObumLdjbFaqng66mrr
fmprgUXSiBensZWBpdjU8XGcsz1Xxf1qg8cP/c/H2W41AsldrAWTb/CyLiwwVoT0Pl/65LaP5k4T
p/KFOYXclCa8d+5SBrQmXFup5220Df55X4iLw9QaQa+MFoM/8wPj5Lh1PCqQeq5WTddNWNJkLR7O
KcvJ7vm7F5lGUyI1CaA9Hb1ungMU6mZlBg0aZ7naWGnpei5WbETeT6dXkHdx4H0edSFliOukDj05
aNlnrFWMnfWXD95uXrAeJbGJWwhPbDs/WxHEnLSnwKgfAJZPXTkvmduSWelw+ToKiNF6Z8Y4ijXl
iOcql1DzKOHcb36ZJd/2lMOnogcr4ckUwR4hlPAivhkAD2gE89GX5z6aSbBB02BOef5hCEWKpLAV
bb7JqJToqx6Nhr9RP4E7wSb9wlkeYvEP8kjkHKXIBjGw75iCih8KOpaaN5Vs9S1jSLrZHx90MYvr
Lk7q6UW9B9SZttXvczs3pEr781NYNg3eL2YGEAUCJS5dDu1Ypn5DHEGMY+kvf6lbMRkLWPLh2m77
Vd1W5+JbhBnBbvzm+QyUla0VF4wyA2xEHCti9HVvgr93n3x3MWi1sOe2eYXEbf6kTo8gPUr4aauz
ILaSXyOjhssp5oyu5GecGsofKoQbVzT+8FeygnVtNNxGBEHcuK7uc3Mp2UbKlE5YcZZfodzh8Cf6
jAIZCtznvs1R8xWG2eVYjUr+4t0O4Qnxs9GL+0SPGaBEh+j/vW7H2LfXiVk2qC5/JGasguKDyhNF
eVcX2UvKYgLw0N5ZB5jDm1nAHb9pMj0jwKEt13U+tcp4wb8aoBML+vhjB/JgNPk8KdyiQj86VvvK
jeFosxmjaHelq1Y3pqwR7to3fSfXD74/H6RaAlQkiHAGkuv8genLM9xuqTAezoDEXdwuE24qzffc
qe958d9yUOwwD0sgXhzLorcIJd4ioTF7RdtJDHYPBrF32L+iyNlfVEsIBjIrk9j2103v7PUvfvUD
COZUIqYImLuG9Qi11draMjSIA8wKR3q5gBKrflbk3AabMNy1Gc3pzHlOx2lKOHxj3Be7qAhqSV2d
21gPlw40g57+3iBZAZumbciuhJOlvHFkFlqaDWm9dySfY9nGBF0vZmDtirrJSQ9udLONX7/dewEr
oE9gFqfGOtnkcZuTBWklH37fkGxXqxrBiJgUGGQMq4Wlu6mVXMPk0zjEurO2cCuCtyaYu7UtmH/N
PqEf8ex6UWew1yyGGYrNuIFN04uzymjqVMxzQorsAlEEt+Z/fN0mcvfJ0hRf8e2wtRuYih4YH0W8
CQ4DusxeqsGp7YsWNxdOC4bM6E8xQ0hQBA70nY/YP9QHA4fU3edHYQn7uGQclAF52IehlZgUhxCD
K5KrFFZa9EpdRQQD6dY0T4GifPKqi66lzudpH4gQeVkRAkSQJhrAKcNLPD3VETVE5e3AEkdRT1S0
MxNf1pEFjqlyNrsdLQMIFEYToGu1Y0/hKpxjTk2RlaJDb648FxHOpt1mtw+pfy3qoh8Y1IxeHgY0
FBCWSU3yaL7FdLbyFNnBVp/U9yuucR8Q7dNu+QU7+RLWT1MmlWcknsarBW85XeoETc8bE9mJq8fx
YF5T1RyeecwhmEkjzajm6JUKRw+KIaMAj1XkIZUfrngVBILmExY2mwP1qXwWS4ywO8PKO1zV6TWU
S1fXlBdthzFQ1XVHjIunl4Zqj2WgUXpxEuB6RWr7xGuNumi0W7/AQh/+uL7SuOuN5j4BMSfItCbd
5eOcpZmi195qIZXVens1DCcaxwz4hj6bqOzc9F78Vx/zW8uGVnqLj1PqcYpiCUvkSII25wCF1VuD
FyO641McqlIz93axaMPbPQiNUvVE7Aos9i1teGVg+gwN0ai146qDQl2CZBGBE+RTxXsxPaTMNUc+
jjWEhArhrzg8KRgMb4ndYt9uRyVkD7JUM7xL9hM0RV+OEAhMqzIU56de1F5DTjh42UQnbiALtZ5z
jrrrLRzNS63/YFxX1bY4fL6I9k6d8ntTLLFA74agKjI5kn2QN6ImeMKz8eAiJLNSK/ZUqoPXnVFz
LUZg+yS83Zud4wZKbCbo5K8HBpsjktGZ/JiWgGsBtztFMrld8KjumArMoogF3RSXuEUCx6+wT5w3
S9P2lBqT5GHbiWvp6xFoziXTTsLJaBxud1vPeouCsAh9WdDcMkh9857eI1jAVpSnLmlAaj8xoVez
CPp2daMmJj5EFcKBIJZkhpIkkSCqcvlHGBkXdMxnjzGRmj7J3TI/ohji2dHglZ6uVEerorF8Mqc2
e5UbemLEpQkIUUugIikUs7jVX5I7VdqYKEwXosk8EPTY8P9f6QRQMpPkPB3VJ7F1iSU/7jKT4zF8
y3s2tkar1KblNe+vKTWz9QGBUiHxCUUKe6pxWEuyXYrirErB6AYxsIbSvPFFi1yRCgYihhZGrZMq
+Zk19mhLWO/TIuQirBmqpabbPQ6Lt5Tgbu8a0sKn6fW5nU9cHkFFlvOYmjz4d4HIm1Iq+US5S5Ct
Ux7INHLcbibOLY8tPwsuKwDWL+qp4E4ji67SRqOMJdTz1QgBw9cvUwIruQ8q7OtI0sR8wHQFp3zH
BEz/5LunVXAYhajGq7p55u/iR6S2T5CqTdPgECyhZulkB8zQEKLOQmhY3UOM0ghrBLHDn/SH4S1z
u2T+qf0Y8tRU85rx5CH/lWj4h4wmDs7SZqa9kD5b9yN/C19JbannAmdwuRTJadxAk+hUBg+etNJc
LPsuLZnh4ovoT17or3vbUvYKJTY6kKqwz+zD2+7Rd36zcUiHSBEDSsQNXJVBa0u/kD1MPGQM7+cp
FyL0i3QOLlwO81/6LJFz1ZybI29UCzEMLM4uZqiqEBXU9YbaVu+/pRpkFiww9lbLXWfrTSSm5vS6
kltqyVowakHcBZd2H3zRCp4XdHBW0bwXCJjqjlzqkLGHhg/vYAtu28f6hqhQ1S+IIEpC4jTwFQ1P
CXw4973qFCl5xbItTEMgZYQAmCp+GJjT7aQTmS65qfCTs0pQJNaYQUwApNS6tsBQL0ld+kM4z5Vz
dJpHaLqDltnTKb5Y29zYY4YY6wjoOIYmhnq9VZKcgjhboe/6yQk7JQARUwHvOiWDFxJds280HYpK
YAaxYBCM/kGvXi5fCZTllbN2K8aYu0tVyhtJpIA0MdpGY/f1FsshFOfRrGTXJ/TkUSWDUM7/huwD
cZTvu85Xc+/w5k9KZQ0jME3Z4xorHSKEGuvbkwSnEeozjWuLJr9vUNageyyoM+q+q1i2Q6XHEcf2
2NvojqiPz5Iw/iVsXWHlYy4D4iwtWbvaCLb4uvrkuePN7n9yndufhir8J8iGEG3S6IPR31GKeQPq
C2TX8KWaxA1M+45glSljR5VPhsqRA0zVRL5bWzNcD/WcbWdyuw16YVO66OkVrpi327e41BlQvhTl
7cd/ZPrCJd+0tFTt0cqP0teT/hG+R82APLyXAqInbA7/xMggHgqkBXj/MZNymzH0j/cToBSJUyzA
X9C0/TdM6Ii5TKGItPSrD1lIp4/WpIqiJipEb3uDjEwAJpUpgJGYzJY9qp/gNkbC+5CV+MaHNgZ7
G9ZXWPKh9AHBcfesMUOMOyQ1GpSF/4MYb6I7IIxKxc8n+1fsIO8Y8n+c9BgDaVK086GmTN2dxaq6
tT1d5mwKFAEYgKZFau8ecbRnKmCAuc+c+If3YCcHOvAzFdTjsbNZ3TLeAG60clUlIqVGcDB/qYr6
bf/sQx8/Ifp3FTl5+rbAUQmcJi9wjuy0kmnO08A8Yo2EaRC0Tp5q+OfTh3N+2xLYAqqX8ZrJCSdu
BDkW8OSw2Y19+gOVW9OytZrhQoE/QF6L7oETSA8upTd12F9AqhpKSMhzICbazM3pbSLUiS3kSyLJ
8l2szJ+LSu2MwuLzSSBzG4QPq2QrIRcnZXhGsmxjN4DqUOoAQPPANVni16L2j9DTh/+dKSRbX8Ch
lIsWbdtuAOSr3epzlxnxTFMGqGiAMHoZkDb0qWCFIEbzICh3SpD+6jibcRjvJueDGMCZHAWJw5gJ
0YVmZaO0iJiQP7pyePN7c+fcikLIMrnalvvikckbyESD/5FDv87Z1XGhnCulHkXGhJeyZmSlcakN
Gr36eqRYUtacPomn0K//nmfDesAZcezX6FsL/5XoQbTwOL4DJI2j1ACbFvc+FRceDwmNCXnNUnIe
j5PVQ1SAzWlihfLEMdIs65IIw7FHNXtjLmUs3Kn4M2B8ZGYttjhwr/KrQtk6eMOGmrg2ckGvdYwW
0LxQG1gq6xPeSoRHnqAyaLAVETzMtgkK79Y8BEqSQK4Pc607Ruo4rg8J4K4GTm9ma+QZmBgRYtvh
NwOtdDMK6nrUgc4kaCWhSxDdvluIDIVDd3RAb7TT6LqV55J9yhgLN3cZKC8OwOONf44AeyEdgPIY
2fkcUysmMQtEKVPtP9wh2NgtdZLBbO04pAnsuvkbgSvvg/9kZRZQ9AoSZvi59e8Txw4vxkimqTGW
9P/qDCDlbJ9SMyglt+mNKA023n3DPgUnvmnYlTgtR56TdvmEufLhM31okgZDZmzzeB46yRfaZsCe
wk0tnXah9Blq2XTErTCFlWaDjR6ihao27H5TRwtYZWfo4bAUJPBSy+bV/jiM72u5tNvbO9PRtZJq
ZPZ5YH4OpQZz0TET586I+D+3vqAQqb0KZE1Yt+0uNWldjSO8CLwnq8NDl92oUhELuEqPrfX9x580
ZdtjLNm6CgM8DAOAKHueSzUVA69tsWoe0jzlXOjZKwq47rVuKOXUYmP6ySHT8NOFk9kDY8qX033J
NvVH+LxxjKxQv4RRdFPiGqsdIjchE0OmcgxeQX0AElJBjuq1ncFbuNuyDqizrZnnqEEnwQT0y8TF
7ryDPZjJ3bqkLVb3nXTMJ+9UlaC8ZPPAcVZqgtgfynDpxlxAZtSy0JB93CmkHRSObdWt7Sts+tA8
AKexWhMOB4Sax1KGKC9R07g6PqtzDP8X5vUHDqp+bvtO3hne/ppJUikY1SMihHClT8kNFJbkf7Ec
zrJHHeoid1DRq4NABI2VoS4h+NzydBl/dn3nyMhs2omONGXujoWuvuxSH9ddQnjKLhSuEXutatSS
5ijXC+jihaI0iPFAuomnFbnYStDGtf4ZloF5KqcTzqacE793T0AALiF0h2+b8DRVSCx+JEP6ELjF
PD4qNqsKAjDGHf9dDq+cWJRzCYUIZZXMNcAOUH0xfdloHaHwF6x/dYAZdGpuBplNOQvvES73UNVP
3PzTUkvvw+nOH71kohY+feOF5QcpVGxvN/Yujks8ocaSrk+wL0R89dhIV79k3uzmNIFWxFfsi4Et
E+d4eRHGBC4O8UpU/8Ir2isLxlUeWD+hUh2nOqjfk22MtK45Lmx1qYBT3JFVPh/6Jw9L1Wn45cZd
ie5/a2sjtapjD3NxeUOYqmVBIrp1UJZyAY3DHWIk3kbpUaDMGnMTJYK8F99Ox23XJyq0RqCHZaSo
a/fyTRQYGB+Sho3fMI6I0U0Df9bjUloPvER4KsEOdDMRO0kl7vfX+2QmYe2vtQ5zH+Z92MDJbTRI
q9HEsC/blZniOV7IwKsSi6dYCGNe6m4fvyrplPgUBpge6IGdtFOWP4lDJOXZL5npMqCunVu9j5vY
yRtvDgXhOyASasv800ZiIvwoqyObkyz5kuKPU3xwdd96B+3c5DfzesUs+TmN6XCnips0UKW7kcg4
FRl8PV2P09JvYtxmh9ukgzbCbameMB905Ba/OLdNLqyisKW6Xgnbjf8lKV9OjTUMxkwmFlXGdMvD
lMfF1Op0r2k73/q1TzfKgtjO73/MKLwEpU1IiE1vSwEB0zRfZmEPMtSuu9/VWNWSRchFnBRRXtZ+
N+EEyF+j78lgODAsK8BHvyqdv/CGNBkgEhsB9q1S8ohJN7Jc33SLeGuV3QZk3JZhRLs7gb5nnJ/I
tHW/CA1TFVeDAUVfOV1Za9jBgVDmBPvWwsxj7cAaBxOSOUnSNhvyYPUbuuK8qHDY0CJQ7J3dxX5j
8mRYRcAG+Yb4p5pGrQvP0JJPen4DbtxiqNSL+rAX6ktBJ/9mPiYD5wReiPBgvx8YmrYQHMTza1Lw
r79wfMxs9rNnj+nILQWNkcXM1t3noSfY8zQyQsm0Xkne9qB0YjnaE8DoKc3xVXB3twrqVxdT8UEt
m6RzDKsHqT3O0ghpu3z9FmoQPzcc69+JM0doj4OMYqdM9XQTCmt9xKTCUTXZpvglTcIuZGv2oI75
P9ig36zDl8xBZz+bLaWj1rluXCOyheGXkUB4QIizjtaB7zfaxS9rlO+eA+6VIrZExI9LiwhWvgYD
SH+ZGoVrvKDCK+cFdTCnBfvDxH/j3pGDUsQfOgQcbm+WVdVBTbU4geEnvKxZ3A5RLLRe5l3VyTNM
k1amCxVidXoRj/itZE4f5C7Lo+FGXcA38TBdvv03QdKaZ+dNdyoczrqn2Ug1hRo8LUIsABP42iWb
oAaevhjNrvQpa4fi7SdXhHHMwX5E0+0dJUA4ulZr7Em/8sFZWIPfvX50KYWqVVOz+2rImcNdRWY4
jTSDiRwerJDYFTBj5ri1a0OmI9Du11K34as3Xwj/+rjfEjFbvDHBF1Qt09q1VyBVnNoha2sc046b
MHHp67+KBiOkbL5w6fO9lI67iYyuEL3Zn5EHdb3dzOwy/SyluOTCizC9EsVty2D7OlEENDkWGDnm
ed7pPK0fqPLB+8Z/yFlZZa5ukXBsRshiiew/9Tin8+i18H4/rGLNPp5LDfi5kA8TTnehrVIyRNE/
zNj9fY/FI27fm1+8sOXPSDgzjN4WPUUZgdNz5i6kNR1xvm77FnokmNcDurC3VRDDUfih+03kGYwF
AARzII6qHiR6GrB8yhNlmkBVxZ6ue1rKEO/WGaWidqtiOF8+lYthZ9ZUw+rZP6Lhf4jqiaNj/GiE
Rqcmwl9iiTfwGS7Ob18j/OmzFGR4BDSEJlim83sU5rvzgXsRf1mfm8MC/o/XWLnWir5XthCrAia+
4CzmlQEynw8jJljKpqHNA1xmu2xC4e+IzUmB14TL7E6qr+rZTUfR21p5YItzTt8p8sgNcF/p1b8/
mHjVOhr8zlTiqmWHlXtm7z9cQAjWswdvgsztc40etAUI+2J5MZer7Xg4KszUdBtpHGPm8++oL1Be
Us2T14oWOpQfN98SR0uCCvJdmF8OQxeOmwhIykmusQAbJOe0QxPsjOeo55SRRQANfCKu+BgAcuT1
xVw5YTTU/OkR50VpphCO3y5v3gECWv0xBfyu3ZEB0TunJmCYUBeWJKkwpZtu22u742PRVXRaw9M2
iSL//azEKoXN7SESAXMJqJOm4z9s7a73xjLvY+USxyuPUJilkJBbAiCdb5huPV4N1NDMucpkAOTO
yeCuF8lIzZmou1GTrB1q7odyOdlXMrMhCmIB2D+Xuqi63u3kY0V4cb7YZmnFaGnQ+FQTO5L6FucA
/NE0JTBj8mUAr1BrzCRlneVIBkullNY+JdBGww+1CHGrOi2gludpVK7DvtsGZq+ChopBb7Duhw4d
7PWot9NAIQ083jhN863Z1IKB0189dPZQbgBxO5fiXqVMwBmvLDpHUpWtNL24vkrbWc6MvmrjqE9U
H/jwhGGyO0TXGc8+vtv0/JyNpjnG80ypJ/9bRXLa/RstAHBGxCh0wFDuE08KTqxzIWKYu9Y93+Rk
TWBrbfzl6OGiFZRD645Abru1T4xPbtoD/A+/88viMni11jh8ltfO52ukaYwu25+ldphVd9VPE94D
iYDcaeHadQCyunNjS39HKT/yw39X01rXr1/BCtuVx+9yOs3b/B2Xqy+hwU+kE1RC1+xLO3+StnPP
0n9mQjBRt2bICZwAFXP+GvO6888Viy+o1u6BcR+XVXv/qIXKZN0kRWvL+ZvCXkgHYh8RBEhdV4+f
gtFO/zh/YUsU5JofSB/GSMIX9YBWa/i+H+JoVtu8kqEwhaktY9HXDtxcrYHwnPCH8gd47AtE0n9L
6wvw9u6x47ObRcqvG6eaVO1f9tHiJQmdQregIZTK55Mv13GfTYEnNorpuQRt7nhWluAll1xbooX9
kGJ0rJqxUEMPyPNIoBgjjJIsmgc+s3zoDlkPkIll7Uv9DpIoT0ps0eqtcagKszmS98eE2Lp1kHVZ
xwb8K1g5NF1vmU060BUv9Vla9erjQHMgDem9GiNRecUT+AE/pIeptKhIJ9F0Gax8gWu/dv0kTPLq
rqWjAuJmAIrp9KIMscrhW5+dFLeHo8xl9aXdCS95mTDGWwW+NtuncZB1UijFlLvLMkNv7JGxun4g
ugs5ZJzekTMahYg/ztbxjLVq8QV02gUFezN5SK02rjZMGY4AuAB0mUIC+f0hFHJyP8T3nKQC4m3g
rTOKVZHglM2N66kj7s8oMWmqDq3p9mPEU5jVkzphjC0THvSBEq6ul7Yw4El+1eP4kXxLju9wMwpF
x0pjIoD24ESY3SDq3tkdt4g5ZrMfFL0ukaJak6uwu/zHU8UKLBoSuoGQTLZJH+wkwKrbagWYPxxm
s+NZVJBV7FSbNwXeazfZ+2iR1FhrysJAtzzFIIb4BjcBBQHslM88KV8oM+EZnAIwiqaKHzp84Bsk
ZqAq5gChewbNOLrZ+OhrrZ9ai2yi8+1ByeUhz/DnRInTouUFF2LNvXL2XVM/MqNT29DNJZqiKCsO
2AYy3LhwcrYgGBDwn/El+Q6NgF52Wc9gdQan1xfmkCWCit1WhKQJmU1VNQo9YRn6vSLkicgRGe5P
FJj8tQ6eW8MCzgLoidc01R+BnENtkIUwn5I0Q52a8/6UhGk5zCfmLt7U5dCO4pci4vsBKx3dw4tZ
2ednCT2++jF4XWJ0o5MxKhgF+ctA8TH0rpxEGJoydkkduQ2zQAQdI65ovT7nutwDbz7gpq4ikKV2
9lYdO6QlT86nV8lKUAi806VUiJMniGVssQbAsLCyP92kKJNwNfERlsl5jbbuN3FPmXjeD2TAe9LY
/6D4y5pTu1EcIsobiOziWxE9XeI5rne+uEYXL0xV1IjNIiJ0WApAue70vwOPoMq3ZM4J3pn2M8px
PJb8g2+riijreSmJof8OB+Q1Gc9DKhoUakYvIlU7Agncj4ui4hhtUA4BEy8S6HOMIabklAFa7izN
k5r07rjxUpiQDqfT7+d9Caq7I2oeYZzWEfhIu6lKIBudYbvBesFu+XEOujVZAHpmnwESaTrMz6iP
FNQFCFR9DVwZfPtYkB2aBAY3ndOAsU3R+fHOuYobUpJn1TF1kK6MS88MYEfv6pDYgu6gZxl1J1oz
6SrU8v060I+oOm0vLQIeXlhRiBbrzxczs9U/7+yTzUqFhMuHctN05pYhbmKlmksiGpAkylW1OgkS
JpC0wB7/JHmFv8VORAtPUztib7Awy4wtnkohyS6/KSEx1dFqEDdYYXIvWMj5Omtq7OtqJ+smqwrm
nuqbgFIlQ8Qlgf+KIB2U0Oqn5Pq9dXtpZ6AP28Lst8sNr79Z8OMU5C8HIq75huZjzYKj5Y+M8jxh
L4QRYaI54NmJkjUCg2zCwdceIrBmnT8mWI/mWRwrPcFs+GEyXoIYGZxfuZWE0zHQUSDSozjg9yco
1hG1tweg8Z3deC1bwtnIelOP+1c84QjBr8RHXXPuhD9xwjbe03ST03TydPgZCeRZkklLzJ9ufyvg
YHhe8l59jZLw8vOHOWH/jvq97AwGlwVkS+dDM2d1MmnsG5s6rPvfJe2aamPtgg0/vm+oD96f7laq
lkT3/la6CkrktXP1JUQuBWhEln3bt960pU2+d7S+BZ+XQxLcLuaVtejxbJNf86LWw7KiYygXQMeJ
q72jNUCaW3F7220hiAEZqpd2qN16UApHl6hiWljoJCZ8Ko4nbjCj0xw3G33j6chBNMFFx0/COuMZ
i4ibbEuUC/2LqxDfexK4I4hw1Xuq5R1oHQdU+kmSIhvrX4ONIcMsjuX96Hc5XIZ2qR2YHcz7SbTA
ZjqXFQyL5huGYKh3tRzRSCEY0M05g+J6GYc05RIkrC2DxzROtxuuWaI6y75giokRBt5FJm1aSf/g
NKcc8HekTjYUi3rh67BdJ4tmgGt1AixPRfhxYm6ti684OgR2CC4FjcjBEoT4ZlwJJTMTNfKa1iSG
8TJT6iWS6GsKGxP3hME5qcqVUSsXR3Z2k/j/vmQjW86JYJGGZpBlNPp4oMOmyNHG2mUVFLHfFlvK
jdcwVqg9o79zYEgfFNB70ki+veg9fZ0ZYGduFg3TJVX7B0flqTJc6SI1cQ7pbudCNotvPyJFjBLj
7neOkfPejaVp4Vl5f1w9IflQ/m2+Tvf3fcpfjXFlg2bsotNZaztkEAq3+E3tAgAy32OFTp7ebeUT
vz5b2fqdJfQwFOo+Vhl9DzDPChDvu310WZt8ktX164NFXTzP6vsIPwHOFQsKxT3GuuxWyc1iuxjJ
cgWhL3CJ1n3JgTAMphDqMqnVzT/fyoqZWZuRiSh7KpfVB1c71SvyA8zLT7udyT+Hioi+G8tjxV/M
T16CAuwi4jj/I17mPnBiQXqmhONSfsVTYBTk6r1yNJvnAAHcZcVE9qtKjf5GlOhMHySNtfvdwu7O
qzklFx4T11zcVR+HmqFqQvP5rSATK67S7Y8z1ZQkXfiVctAt27zpoR0WpQSr6ByH8KaRGWarS9wq
cXLhffMH2KJKiISPOnzqLUiByqtKKud+mJo0bV4XXuK/HQynPkxSXktxxHQseZoKELT/KcboL3mo
dxBQUkYyMjA6QiAE1yNe9c5wJHHyLTj3gpaKyASbwv/OkM9uNwuQsYZntbLcdpg796OEHxZjCe/D
w17JWCd/RQ3o0u0B23zJULu/uN9bI1mRRXD7jqw/1QIT4HfjmtuPWchE1qFlLwvAMt6AuIAmkIQy
2dTUw2w8Xopa9D206UozRiquilScotENw820oLqmh1vkKqONfLQTYA/YDZr7ZPIDaQLE3m9yGxZg
loJQwACfdE8F48xefw/ONz1ccrPTCFjvJp7bB11bxydNWy8lFBRMBpHbDy0DG+/s82bPFmh18MDq
Ys8Ptm8bn4OgfI1rGuF0zG9bYmNXB2l25q/pXPfMqrlf7K33bqDZihbNfE46NM/fYOBrLXfp9uhU
vrQVngetQrVy8OSoLlQrXDYqPn4OWly+vksje1zWFbnQZOu7uczCqpeqc6gsEwRDNPgoi1O1tLWn
2+GLCiYCtKSKmI2u3/rTHooAo3kpBPJxfN1n7ZBMky3vnRgNUf7AMLL8E1oGkfB2c8NIgPf7c+Cp
Pr7SUWteNwPgw9+eyJlxdBAi3vZI1040FHBlE2aypzjT1jlXi0Sho4ymFKNEiJZ78Q/Ro+nWj/MG
zl7hJLRlKm1sh+3stFnCD2jPraTzY0dPcsfRC+SjGzMBhx/BYw/f3ahW6AhsK49pvAFxND+TNjWS
VLK+CKPelg18CDxkuXh+KOi+dt1WyUEjBchgjydIulbEnVqTDEREZS/26wFc5Cy2bVKvznPXbMbb
MtZfSc7Rza5x8QqbtwPXSersKVeOli/eerJYxkwQM4ean9hFR2/UYkzYdIXd8LSoy4OqQqxe+Bzz
LRjvxABgPjmDzYtcM2O8punCZMiOJcjPiI0KP6uT24qExd0gk5Fi0jIRL4bpXW6U05cVYGHUmu7K
pdZY54HhpQSdyuavZS7eux5FkDw1jDC0ME/HIINJpEhAa8vsaDaFi5MdFEd9/YwloUcF769rOgIn
hJy3+g0mf5Kj6ofZVPB5t46jlFBCfP/lBzLHnV0VBxhvgNNpNuTS1YPxAzx5Vr8oV3oTwsK+eLQu
kE7s1iptz4LFl4GURKJFVqWE6n9scuQKEQTi5TcZJH1WpCx4FNXPev7Q1PCD2uXIAtElp6kqCjWC
tJCUyscPmC28LG0zx1uoa942hyX4SqkqtHUU1hM4Mw90fSfzhScfJgNmNak5+UYvb0xHsj1rlOCS
sHgIZ2+4Z6EhPpelXcJ/ukRErN3l+Lt78DlIKKJjE4y6/h0GurIWZiZfAnhS66++SvQVLA9U5HXp
xCiidD5w4PSnXWCs94UpyFBDjeDWmxgS2IUV2OXC/hbcN7YFP6/x0YdBHX75ZO6J9GxdDIEWOQJ5
/gE7pK8K6vvoUspUXTJIEcvWB7BVMsMkS6+wHdL0aqgu9kjVNsyUcT+ZV+wEpbIRD4TjwsHbPPSv
Zev0lzk1SZQ0TIXhjFngi5J4DD0MU3S4BgVTQGYuKgYucQiN3L7aOVVRHYmzRyXy2az7xOWshWqt
Z6LqSKjuhBw0MUDSAFSdLnh1gg40qJmNr/LhGmubp2ushb4+CqnhdbIAxEHUGsszJOarz8zBWuQN
SDKHSYM58ZMuKI3hhrgDSbTUvn3AgOVFt90pGFwcldILlYjpyZiG46yw6MQKLhDR0tnxx1EPgjow
+kv2bSYlUtJlh9Ivv0zyRB8IFN3kFF6etzS4NovR46J6bi9JJD2IUl9oliojSVXdg+VxC+y3246h
K/nSc50PNnv6TCsoDKaphixr1LU7Sf8wHk1BbqycBAe/2qVZpY9Ilz7lhVhC4Ksz+8NAG9gMhYpQ
ZoBMBv94MZ1TmCsLawq3m4EyfwoigRhJwdp2j/5xsDOuCMUF0qnspZe/iHwyTePp/rxIOHL5g90+
SkbGoa9ih5gmfrdYR9jcbEDgBzyCRr27mas86XkT3pRtj2ZhMuofQxeap0z+zsQuwcBeacZfvyL3
t8EbbtlX0xcLdcaBN30w9eRaiwe1sV5eLHTbAoZXsFBC03VxR7+Vql/R9xoFfmKnBW5oPee+q8vS
LWgwsKxpDYKhqv8UDhwQVo4tVMzepcxiuAExbH3euA+a6gRyql0yjBcoiEV2qg2yCZFEkvy4Vkld
gotJ1CAgt3iWRi6uX5Kk+vzZdUODPo0YEFRaXYOlCvPA8bxDczJROa3aF4CCYw4FIRhasDZTwesW
9Xf32TbbzBU2Pv8Ezl9YpxEc5SsqZRf7sIAj4HMhqpq6fn7y6QqGSSGF0JBvNtHM8HOSnsAkeffj
SWuDFUBWFhAuCBGANmvE91m5wVJMNrMRPqmHnobzjDbmlOxvZZjJ3h1A9JMCXRDUFOh2Ht82+VGd
08y4LWLuon3blUpnivmhZUK/gSYmO4NxMlY9Ih0bNtCuMEHnuE84SCKvLLqhXL1HmFMeN7feuN8H
s4NK93kceRNT4kFr6ZOOhOCFBcLsaX4PaZhWPijiFI4ARN1jFctK1dau7zS1F+tFnmeI+20cv5y+
nqIOutlmjaOMANishF5/RZlH78l07zqlHwEcS9svohv70QLDy3yl5InOAaI4BQttzGQt8yXycLTx
vtr0eyuo9GaIcJuIVXcTvS4CDAAWMmIRwd0SDauB3ePhXYmlJxQgu/myz7tbUwk8K9tW1Fz9TX0+
BgZ93Gt0htSJ7a8Jji/Erzxrru4urMM3cZ+PM0A2KCUvGYP+GjTMWySZZymYmOm+Il4I2iYVp+4V
xSnsE4xi5Tgs93xAaA3T5cjqgke1atrGCvcKeAcK+UC1Aw/k39H3mnDzzgX7abs8p6yejW1OmIps
0o347YsdwY+GDHZ8gUPTDjbamiIlpePzq4rRO0vwlCsYHH5lgfl59czTMj04tHNUBHp4//jT1YF+
BesGr9xqx8bwo7jo9wskNJNouufkqQZvmhlv8K1mIFY1bqGXsw0yINDUBI6xOfwacU05RpLkQscy
bQa27Y+2Ulx1kFcyf0FG+ku7ISQuX1BM8PBoLO1o4c7rhWLVPNgD1I7oTh+DjNQm8O+qMZv+trBk
1X07m4U4ts7Q9A9zi/wKJi7D1X22EVO+uiTQVeMokoJGLBrpCOHYtnHCfwJ47mGu1QSdI5A+h9Wr
FK47FQTJtugb+a1kuLshpY+C1TovTeL4NpCPMCLS44t2AEbglpi0SYz7k0WQQQaT9xzs1S9KCpgD
447mOWPVqXVz0IGbmSvHj1/hYCze6h6WmE3ZcMiehOYrV/5eDDz6j7emgX8qKlL6N0d/6TQgMW01
uvKG1Jd56xLoKv21AnJMfgz3488+7j+w901FNDD+uPeYVImfqEZfRd4kDhJQaJpVc+CH0GMk1+Z2
/UOq9iVJribTLiQtLN91RW26jKn3AATzU/ANc0nRCvYtWq92JxkvebUruU6GwY3LxIIz6w0jlF8F
U9HLqRXjUmHSTG/kzhnj9oahUJ8E8X96Ks4xvNX2ErkwfkPw4Ctr52sOdLFz8zDv0SCqklx6iCiU
LP9KupbFG9KDdYNcJ9by7TQfa+pC4HuaU8qZL3wDaFZaUTaZh5Hm11ZJpFYa90GiuDgRWhDxBG13
7FUPxDi3mHwkXi4vQNNsqZ3Pxo5EUCLOrdNwlZC86gLfxVeGTF4KWSqD/x7huXnFhROU1Njv5PRJ
PvoSZsgi0vrrR61JNMHK6UCF9hUZMOScsG3uiey2+7OGALhh2ulcTkmtoiLJRXfqgUrIf17z2ieV
g7gUJCai+hR1NZEVnfFATNSs7N/6nLrKZQwIal6P8cibhmh97ph59Qanwin+UIuvM+fIJ7xvJFK6
B+wRFA5L4B8f/v5S7xquR6q7zALCbV8D9CpkwNtfhALVSvL5yJwRwksRwEgl7tsfqBd+Pb9kLfwc
21yaiJL3kxdPaMu9OH4AJm6RlvKj/SJOpIctAvluNC7laa3Ckx01OHalav0fzkedwghwqbWbjFW7
VJs7lsTp5gT7fy3HXhOPUDnDdrGOJUKBHezMp0lI4ijJ0defSvemtL9nRApkqU43jGfXsnfB/y81
5GLYAqHEBjxyf+v4N8kA9F4LD3Bg5p7ie8nhUxHJKzb+ACMiJLNhT7GqOPNiPGHsDlcnJa3a8qKm
5Qu1KW6IIDNOfMtTwhI6akWZyiXQYUnVb0CLNECvxAdUmoau9ZDravFdKCtqgZcu6I9NauFURJ4Y
ommGDqkJMHu6CvaNH0HeGZLq9r9U98Nm+6t5X9gIyaZDx+0gfPwt0Hv2GUFSFXHsKFB5Vj/K67SB
uKhzLgFvttcWHkfLPFHq81lWuxFar4CwtQeJqrENlQnyzxSlwahMjxNdJjOVggBffZfZ64G00L9c
gElqZ9cTCufBnGucxiFCwfe202+XRy4so9uWif+2ih67D5nmTZxFTAqyQm5LsgbuJ/9xCuiPg6Sn
acplrp3L0sjOFpG7tQw1QWfeooc4JNn0ZFxqtKIkpUWa/dmoCJ4IYbsITFcFFR+oxo7b0HpfO6xH
kF84mx3wgOenDp3TndkQv54fEJwV5qYMmQdnWS8oThzgbGDKmPvQuAnlbY0nyt7G+jlzANk/w/Ap
+foCyWYWjLdi1TeSHVkPAZZCj/+bwkyag63QObB/TKQXm1iDwwFBr/NG4j9GbFfGhq9RlwKqXspV
Ju7XJf4dh752zYPVQhKfezoUlekniot7ueOzE+lrg2r44KYLekK1r/HMH/ylryMLBEVyYqiKp/Ax
16OSnT5rGxhUDRJZtm4qVJg2kU1qndVoKA/hh2pdupWhDldiRp5p7J/SA2diyj3dYF18tJCusx3t
lq/bZ4rUbTe+IuJ3ESKTQVfgPkDVPoJkH3EiWpyuP4qpDWT+5Y96MSjePjzBa2CBxbR9PpXTxPoz
a97fobsQgdHaXL5wXzVoL0hrBjGLrn8GVCo2GoTmqjtaCmxFtvRuKD6h+UaxA2VAVV/EceY2EBIx
opwX/KXjA5GM0XqbeC63IiSj2o3coxKgQyy8sT43sQuLgKjvvzCWIHFB4ayxoix8eJzfFkb2siUX
HGPc8GZN6vCiRStUk4qRa5er7sVLA9/YGCu0kxeRi1Rw72G+S+yxs99VDptzQQ6Lda+n5L3R/SGO
1KayPBqGx+KFmcIHE6m3ZFGwKjHPXRjvvl7Ct/QPOwvNROmnAoe9FknJ5y//uuw9q14dabn4XMcF
hDjMQlzEMhdlYNq7gcB4QXZ6tGwtkvwhG7e8tmochZozKrVILBubsmyBG83/4vxcdW0nr3pl2x6Y
NwP2XcQsohQKIo3vci/ESwSvqybWEBHhvc1L/jglKr4ZOOteVMC9CL6dQJs+f/lRvDKDdA8Tu5Mm
0APFEN42AlTeSS8/fuZg3pWPy3qtsBzf7Iuqef47DtXXwuxZ5M26esHTBrRt1l6f5h5GOqBcGQAx
jWY0tABIWkJj+bGNK0uw42Fi9qOg3trse77rJLIdaRGGl0c2KhpDuFYl7rm7FAHI/2VNYzK7vpZ5
gs9YiyHhauSoxbc43pXWRh5fax+WlaIezSNEdbAZ0MfH9h7aAFym3OjDpHwYq1wBiaSxW0E77ouH
Kj3h/skeVhbNXgT8bWqQBjQ9gZR0F3JTFj5ROidkXBe06jlt7nr2eI2G9q1nb4jXB5ECXXnuVfyM
oI4FlclGsBYq1FZUEAC73IaBMfMEXpzjUWvVHA9/UrO60vuwIbmtofIOsmwcnp+M6te9X4EPz8nw
kxYiHEE2h7aMVlz0yxFWuekQP455iEqQ6xZfVM2MvXo3IzOfyunkK2KIGoMmxE9Gj2OC8XcE29FG
2TBk944jA+OzDpwpffCKgdgGey5kajsrEIFZ9WcprUKZzryN0bpfjmw+1d+9TrAKCRKL8ZU8Ozau
NG3DkAhFjM1tXCRbuDCgTcYfs/b9R00P/+p6vlo1GvyUOPh6WjGQAB1xYsnVATCrQwhfNSuQOcBd
RFbCYh7BIpbtSrSzy3/oP9iJlCjscNgZJJ75fWNj8ne/Ls4yl0tIZP8CW3xjrTfdY8JobOYp8gd3
a/OIiES3fsd6aRkiqyOW9/G9HKgoi1uQ3R6AaeGEn5RLdtmm29fqern9prqtDNFshEk2T+ikcb21
gRbWjDv+CzAvd2py9E0dMkLr0U0giWlc68g7QphjYHtYPqYPtkEoaftcz+REHaVXWovQwEufgzQi
SivP0zySXRMJTGaLwKRRPQFSQJlqoozobr2yZASEXLaLkHrw/vuxkcsptydtzCWN+aKd6HDvBokR
rdjDF/sTQj/F+U4fVjxFEejXskxKkmGWx/uvuU7RaaEwZmZuRwOeMmn2gtsAzoSvAquQpKbexFuk
jBt8zLqUOFj6GqlaINQxlQWbvpeA/D9stw/pm3Eq5XiTvfPmmbqD6iVF0HN2ko1lNj+5Kc4c+qTv
5EezKsaDaverP7DfRWv+9gsVkQ7gzNBB7AQPRU91d1Uo269GWEkBOeA4SIWMwH03KPwpJmo3AX2Q
hE+OIvqleE9vPvnIfpock0sknAER9lBgpJGBE2q/lem/aDANHKVOKAAwaS5tHmEfihzPybyAWCsV
Dr9hoBxn/6xUBL3BvC9MZ32cUej1l3UbDhd6e90UssS1K2O9YJoKbsypq9wQ8DB7z5oJHx75Vtrh
qA2/1Tejg/SxBqVNOrzzirvAazCzC5cbRvd/XuMb0xugrjVmFitjNum4VGMF9HSrwbpXZ64NPFM6
cBTa2W2VAc4vpScftseID2VjAmX27fimGh6062PtEDDUgNvNxK36HYOf582o08nXbv7C3blCfRyc
9ztqx6hZTAOHtfgvW/jrbDUE9pzaoDM4cK1zlV6VAHXjVTnQB5d+wfvnjPTx3zLltEKHaes2UcNC
xtKgq1YTNWqpoZNmr83tHyXpeKyH6LDMXJdbFITfMjpZXqQ+F6eh8Ib7UVLjCJi8Uf52WbZTMA1b
3mR3R+AVwiZ4jok4ONsoLdAObsvQh/ijVe1QJiGYElSdHc7V2c5FhQUqV+HLUIAUzWqcIifzyImO
wQ2zHzbFU0RM9bl45lca700dit5VixN4roeqak3aU8bXUIga5O1c3QCsKTlTa/hFH9DdaZgntX7V
nie5bt0WI/awdaNELwGMvLBxbnh3ri/v0L0zoMB9wWC+dKQobJJGlhd5mzRN3RQh+u5L+ntVCjuO
K1Qm/DNYHjGfOVCmLka0TC8oqbPsi0JOgyPg9lrmUPwls/6NmwZPOFENbaeWSyRACux97V81vM72
iVMTNm2TaMX8aA5YNU1uhTZozdZo/uHxbq1hJnBYrqlzyt5slIvvsioJ5wxRbHMS2CXC0xGAfkY7
HgmdfHxI+V7yWOSM79naugrgdgwZDa+rPMgbVc7fxRQitmkbynOAFgVz+B5GktRXAWqrraEgW9SM
Cv7Z59SUiwwPg9BkCSxFGQuKA26HeAt21COPixjwonpD0iWPlOYR/2cnGUbuIDaj4q1vKx36TroN
zdKW9fMZGP9tNQ9qwE8WYYpnrmgX9K1mLBjD8l4hmOhhz5fV0V+rFpsLOljqa3/h6bskTV0tlJfF
IDl105xTLW2HDbPIb0r8NDu9EeZADY0C9EGcl9iW4/M4EqRHKH3+1AWi96As8eFApJx2tmEy3ei8
rm9ATk0wTyx6I2NZjqwO8mUnRIyH8IyUIVDrVCdj4RuMhKNvSRM2kI0nDHUaUReQmZoM7Kz70Hff
+V75E7b4KhrYjXHz9LurDhGg3YIdGiadaa0V7lP6nFycFi5dx4BreWVwqscCYvXHpZPRP0YmHnEy
3TMWmso6M0kDvXWzfMohKv0jQSQGEGyw3illKbIRClVVIbizgeo7SlK4t2oKWm/S7X4JV9HqDDZH
NojYaq6d3MELMUdEaWQU/4cQz8EiaNIUwBW+Wfq6+rJoqoC2Yfu87eUC2fLj0OM0uD/UgAwDxO6O
0xj+3R8nDPbBEnryflO/5aSTzz1wAVA/Bz2X5oFtfKUowYiKho7l1Pw61oAsRjRrG3qpE6LGXeZ+
jomddC+h1nXVO05cdyuw8DysRNSC+G798cPHUrxFC1PzR3uW6BwAEdB6i910N2oaXmNL4SBvEGha
OHHqYL19gTGVfoyahwMvuKUY4iI4WBZeW5DX/vlUO5zYVbpQzBSPhuaqYww9xOLeGmV9Q/GqHk23
cZebKiF0uxsIdCj+j4qA8DYvSsmqzpPNLbp2HxM0evmFytw6VNF7/hNxMLuF9o/6w1BUIj/TAUvY
oe/qe4zw8CiRZINjpQrPcGAMtrZUl6Wc3VeKQ3PBzgn7hPO9c5m6EIOOVVvpEF3OD/jMSzqFCJb1
hUH3aYX4Sx+bcCJBmCBcj4Csgdrq/9PHTKg8rXd8YXD371NjDnr70WKniAalHY58+KxA3ZaT/Ls2
BXfZB0XvXISpS7KkX79iNyD9Db3wXM9aQ98JYUxujZFzEGfioW0yNmIv0kiVj6z1rF8LMJ+f6g9W
Bakn+8aIhQLApeMogfDZeUaRdtfYf1CYgbJUUS4xpfceBH/Dwsx6HiVjDKlD1hru9f93bZs92rUe
BO5w2w9wbDf1hpFN5a2aCpLMFO2CLQ00brVY02FMUt3TKVi+KPEgPsPqnb5h6AJGPmV1OkLLNPNm
krhBwXTB/Reiw920MX7xzVIASExrTTt3mynb0njjH7KDLL7SUkYsmOHBiyAsebn1EjokvsT/0oNK
7ZkzwpioEonLSaNH0/Zfnan7EImPGVUDrK/tU0CnaqdI9O2pV+xZLVtKCIHF6eXFwzMWeTIpRQyU
CwKLAuXO64b3eFnR5aAc0qMvNpEDb++7qeKQxQ7wpu4YsgPypTdWMiOZqZ1ugOtPXf8SSIdMUfaK
+JIwU66WdvNHDTL19F68HNAQWyNUq/qLTUDNIigehunhxoK/7Fb7UZ3M4+1pewXdlpSNL7auoPsa
eM/LAcyecPI191GaihCWY/ehN8WTIExMZOFWLU/WgEGf8SCSOmnFQ30GENf1/xB9a0yMNOgL7cgu
or3Sh3eZXIekYQeExguUF/gtqVDrG0P6p/2XMnst4UNHHGP+kskSLJcCNJWifjocK15VBI9fQW/t
7meT+cfF1mg5o8CEUCxBiAxBHpOKMH9lCny6+7nTKR2S4vhIrNs8N04O/bzpFv7xZ9Hu5Met+37L
CAkX2N1bsVHVmR5XARiEDOFYGvAzpRmPBYvSfd98SWYS7nrIemaCdn4GYqbhZAqsq2xu2zBakI0L
4RuSclC5gWuimTBR8IanIT5V8Tb31pBZwxpiIanTh4fuRwNAkn95y1hNOvkaZEEGqVtrR2oGXY8k
dfNTANfTkzc6FYDVy0/UBCP6g+5Yl8NWtX2EJBTwBSRMpas39k4GoHSzm8GCqfyaH6VtVyy5RWrY
cQSADKoM3W/u0Dx5cd+5jRwmVHpG2mj8wAdgVUVME5ClLVqkCK55ll3K6KYgYviEUp/BelEru9md
9Yw5Ew1YNOlos+5Sk99M/HzGAn8n/rbsEJaMN1bmBGBfeuu7YbQRPBVZT/+c32Wm0k/QGiYy13Fm
c+lGciGQ30Em88a92asmcM1T4kfxg0WVj0pnRaKedBEFeBQ/SOcBG98L9NC7ObWsW8ymAEA0FamA
9htkQkLagklQolsCo/UFm9GS2fZNG+TsAkmTtBzo0Tyyv6YCd2nwHxtAgOstxhepWRUKsq4w5geL
cis2JPHvC8w/k8teI4W2O6LE2yw0KH5kfIZOUMzD+xgdw/ygXh1UY8AN41dvTbJI222Kf8eA373m
SumvBTvXyENEgRyFa1iro9H38CDiJjBBJuLhXWC7bAfKzkFIGBOkMTBEjCXL9ff/LOLc3tVE90tf
93DqOoC3X9egpex+BCAc8hzUCUry2j7Pez7vkfyoRGDtSuOLeupwKR7PwIC2wmJR5Kos+7+wMJsh
8XwDAuOJDKWZYPXTWYU3Xu9NYVdnkh3ovy0E35y2M9p6dsIUVIiVJMm2Sma0QCmGBkGgD8mfW52k
jGsXz/YbFn0dlLPzCFMXLkBsK7Pv32SgEO7qw7acR8N6nYhJg0iyYQB4keXlpO6dYEeqhtO+dJQY
GMA9DStHyxXrAjAyAUU0zxhHaqozCeDgPVeq0gpOxHi/HGRCspTxOGuZY46dNQ2rZgsYWfMFbrHl
SPtsi+qHb/6rUEFB3QBgDi0e+VloVFaeZK5l3fO3TJoBvt5SuGhqoZSY1GNUj4LLRBFM9iDuYLv1
uME2AOL0cY4IOpPz6NVjQiTHQU9VbzNEIRQfPxDcl7Bk1WUcUci3NDE570YDCU3Vc+ZzWJzdFL64
Mws8cCGXoqXhMEU1HGsYyMheki/W0cAyFaq3GCFFIIKDkYEFjGMZnIc/yJxU7ji4zUD1hzF/QpR4
bS/6E+1sJeqGNmvvoZt8VweJo0VZgGZOlQbIum4zAJVep/vYEBUhr/ghzcJnp0p3jhia7z4qJbL8
I8ugjCLHVLLXG6Ch2l8cVl/iL5isLUOtviaLN2jXZDaN8y4PbLvWZFRh57aB+ve5GdUO3thU0QGJ
l27Xt5aRLYj/9EsjCzG29q86Wjc6liewmR6U37kiISdIDADoPSVSV8lFGeTdvUo8l2/DyPQoi27V
AKcSCHeBK4hp88hadZZeMU5QZlhMLguAFRzihP0TABicKyEcj1r8Va1ZOLoMOUHp08zZ4quhFSGL
6cO3ZUWlWn3+PtwvIcM1msL9EJGtVu3bPQq+3xWZlkd2JcA8wr5PDLtZlxRTsN+kmgCjL0fLX6Pv
aKIgamm1277jpQc1MLjASBXLmesHVJOQl9Xo0rgUMOnQUy5BT0iFHjireDy3Oi4NkSjCvO21p4R8
Plqxsfg2GaZRmB5FLK0alcvmdetRbwPoIZYv/knuww7lea7j/+0dJ/afK0L1dJwwMDiITPhe9Q05
rnbb+jcpZHwGGGJNvYccmdyXLnqd64mw6C2wjFiTBgkFghsGiGTuKNnh0DF7VzMdfcTGr6IrgTtj
997x0vgft56HusiHrVDOfAEwClwNV+QwVqrq+XG++vCYYYL3GFhq7IDnV2eabDoX9j9BJQn3UH8u
Jzz92B/d/stlbg3wOXiVqVaIr1ss6j4nu7I+TleHCZwa83ay/TuVpUeQw0AyXZHMoHiSR9YeXlGN
T+tYeCwumN3cB4V4x83cS1moMs12Efu0J7elRROwVajxAUs0JjOIix4KgX2urqLdcSL7ZyE9lQAL
LO6mWt3a88IacLg2F2MEY/SnkfTLLiHcAUvx9BFW6/zDa1bGrXVhm+EI1C/6MSioyW2sf36zmn/f
WFx7Ou2oNbfXCImjT2OU8d9qUo6lCgq2PzBfiAM/pyevm3oeB/co0Z9Zg2G68QRSU9asVIgS7PoI
j2OkWuBX5hfddUonuro7EWRVq1b5B94bbylWPy32jUkFqgJKC6i+OmxmamCiwRh3gAmnmJV6sbZj
pKeQXLgcDB2X8PB2cPpfPzuczqVE5xBlxjYSGXIDAl7nZe4YgkEJrT+S+BSthlw0rVUmmkxfqRfr
MK2/Jc7Ew5BJlUhdNlRNAUilZuQ1GhcXUs2f88SIUAvIokHrXvuOWfSe70LB8KEBad++qLzYY9DX
oPqiiSlwda9DyUb8Cd5PPSXH/4RtOzniE741FDa4sgkphc2REZ9byMypA2KhqLKtrTS2DppmjBXf
QcFtALu7sdpw84i4Q8SseYQNGPFUI0bOo7GNBDcGTyU9VDpzOQ4fcEUZ9w2ifH5YshznWtbgsrKy
rYKm4BEGgrdhFslHt5jlJE9gKl5QETuSImCUvGN1kja3kUWxTJy7RtOXrU73FGAVwVTQXwd0Ew+u
zDq3stqdQsulsX6nl6SIUbEz6YnOYhT8Olgoo/iRqCad3qLBoUAoof5XwtCu0iq6z2DCKUrBjUL+
xherd9g4JPlB8rG+xrs7rEs1Qd3DOcut4/rNljDhY58REMIbGfFYEkZ/mym+DJ7QwLTwvREvgtgE
IxCoFlqovIwdAx4m0ddkS8LVGAdMI+rS1xJ9VYbiQ1n6ku+Qn6BGybzKKinnMU5urK6W6IRVS1IL
k2R7DNeuwp0EGtmXTCaZpazP8LgUM+dL5JLAsmNeBC1ov4R34TH2MgNsvUfoIDzaCht10VpIOb+z
oAQbFUIH+GkJqGDfh0UNb3mu5j2s22v8/XUOCFKgr1MD25VqyjvO+xzSoYtX+nxC9maFQxUlKjOH
BpXeJe8X3f9/asAuOH6x4fG+kFEFX5zpt4Z2ioM+Ux7o2BVb1rVBwiw9PkbjHR9dFnjWee4uoWLb
VbPduN9SZaLy5w7m3XxsxJlvFPaQv9OlbIu9ZfJLqdBMSAjB+1LFIllrBrSU6ej+r5nchD5LYkAD
BSVmrjcVt7WGO6ptJImtJkdkqlNEdGXM7c4pC3bnzgQ0RdoAKOgXlfeSk91fqA5sjwAIHbsZs/Ay
KhypIbe5VOlprA6ef3Qva/FcGTwSVHlGetsZ99cv7wOlGdE7b6MnUMVEYJt1dngUJ1+Um4AhGUoQ
i5ZJP3cD9ksY+v80PcFatkJ3EzT+S9sbPqjhw5dySHgatcRC3pj11iI4LEImb6ybdNyqpwr64lcA
uhYbj+FbNnBx7dVkTcsUIJj++Y/1NnsjjNmMlyBFqYWwGawuc1dGT0umJ2hfFJo0niT0wjJMJ880
iFYrmF9+wqKwZ/m3Yc90MzmcZfLnPsQEdhcTYG3ux1Xw2dBbV5vxrtyvTBBcca8/aQnayeqAS+Zz
VUENEIs/DjyjVQV9BCvDWgxG+kHui5+xYrx8RuG7mQ88QrHQVxDN8H1z2ZGlE8o/XCBktbnKSQyG
TiFr0T/srN9FuF52cBJRXzTPGFN5bAdrOVc3gVQeb47tAwc53jCHK/E9w4QLO73vsKPoGUlWDoYT
YOsqD+lOFlg7wFKhwiHVLcHbOkbWnZrV97RmT87su4nbTr7SEhmB9yUlbuaY6R5LgF+WgYd9GScG
9Qh9Oc/2bd3KIDFe8AA/E0AscEF23hf2pFx+dYr4ZMCQGxpAtXLHsZyou+xH/f8+3CzKLH+GxiZp
ZUlXLjhfcysymGwAF8+cdzPGE5jZe3CKRlzq9it0GPEcc0UeCd7iHs3EWpm97XOP5zphWcjOhidM
oEAXTuhAo23GG16/gDc7bJa7CflVpWmEfdSV3dGXEE20mnAMYkEh67qbBP35vtoNhY57Gaowf90w
45fzKmh8D3ny2GtxBqASSGjGdoE15A+WYa+prymXyYRN3pqjfYVEZy4Qx9HZ6dUY0nXtz6WkzDf8
GQTpEK9u8yZn8Ne/YdXXcDbZRdF7lSMFhUWiTuj0dMlI+pd5gxRwnfLF2Gsk7fVhSzoXzKxHnlLE
BEOXdyNR0kYWoODMSMumU1hmRirHDYUZYbFec+2auUxzww1DMbx+O1RjHUQgzTRbDdsAu26ol7uO
LBjNcFOQJYguF6tsrNwrXJfNbCjgyI2UIvRRMvwVmzKnYHMFfJXtjWeo1G8MYkDD2Rb5Zl4FtrgQ
MDOYMgiEk3X1d7UeKRAandJqz1j6xmyPf8rS3V4Pku4BNwSBtNqWwwuXKc5npRRhXL48J9TzdgdY
mR8gLQDMRC1ScW7J9IbaznvazM/bCXLSwgSCXRUu4bIma3+5SUrZIb0ciR0y4VUQPgWO1sa8o9i4
DA82fHyWgaXEHGeWTgb5bceohY50Lfwk8E6y+SAIFnxKk9tVjyRLjf5ElklWkoVI5UbacFtgEOnM
uUtO0TNaNAoEnRnz9xgaKuek917yPcjoVtrxwEf7hgLFa28cEl2WD7GrK8hc4O72pmA62KAPLd1H
z0Bl1cAp6a0dVIPswTELZLBIDTsM7HabLRZy7D3SRq7L0rlQm/bZ1bVzOR67BYGOVE8zmma7gC/4
tk4cSAQx/6Lxnwc2ABdOhv/3Gd/YYJcEYGPXP+nuI5nhIpr+aB+NWizTEz17Ggbna5coznXvi7tI
r3Tn6bfV15wr8qkjTzVSjL5XhM+zzrCf/SeoZ9sNdhg7dvkrJZaxadQOUmVLsGZD4x5zyiiabHB5
zpWUqj0JJRwmxdKq4V10BrNHSdRP8/hQlO/CfB653ouLOSChJuXgy3QPf9u+80rms78P1ljdHU9y
4YPWsB4VZ+s7Ai7GDMwDOkFANiLjdPwIX3JBNHomJG/OFWTUf8lDaGc1KAPQgwwahlLFKOwz9FYM
tYP3V1gwsi8b8VVKsWwPitJ2dAceaqxCGx5Tf0fQq02lTmRoYJS4/H9DF2f5By1fAWLTz3PdxfFE
36+KCUgui5pt/ETq6d4IlCkXkgM/Ef1eoV5hLFtw7HbOxYD2gv3tCT5is8JSxqUUjIKju8z1klNe
JMjNvG74hqcPrnfshCRifX5lWU7/JxC5FP3DJ6ZC6aIwSqW6n3qXYuSR2JqGjJnv7l4aYOtKCN4l
GxQaHSonftznvzcurTQxrbVO9w4zzS6O3FSmv9ZRIyR7AI/s1eHAAE8CqjcSDoW6DwrDGe5utPrm
IfSAjo1geW1hCNv6UCs4QrjodZkPOtZfIgQERaE4ovAVrcfpjT1NNNPHMjgkn8XxmTbsGg+gb7vF
9V1mWZ8LZvxZmpnHbSaREUkbUn7YYd+4ijViCMFtiLUqs1EGZLRjyO0dfmzx1RnnX1/JJ8BtDMJm
2b5566YFo5T9ByY5Hm3AessvmLSnjNaDsF5l0mFV5jdBj2RdN9IcYr5GXNFHJ+1MMauI5QnKka+M
wLJNecDtaF+d0B1gbCGR0ECfGpzJvW3k8P857IOF9I68iF1DUnp00I1Y2DyBz5eStkkT7p0L0I4/
nEf6Ew3MHAHAHMc8gwizHhXIfq0IPLFU7axGEfxvyEr0S+Ov5UPTh9AuV1lc3GjNE6QuujKdi13I
CRAzlauT4WpcHOE8KtAIO7vQelW+zjbNTvTyvY7JYuxnt+mc174xPcs0O0b7izHk4iRez11FUPfn
t+CGHqB0HgjJXzbxTlLBzaGhcX+Et/b0h1Wi4R5prsKA8IqdS6xOXd+kRBaJyqdpM/HLWtsbHq/e
m+uzTI0ZwBFvA5FJu8jfScE8c1uqtBDo/zRdZAbV7KI+9npt4Nw7eT4NiAaV9WJtmclnouR2FyCD
xWTmkLe/qt40DQQayjb914niRMPjjVeeyFgZlI4KBlzf0kH9Y9ECPGhF9EevfuLvwqR4O0T172fI
UAlXWSGuWpe7PracmI6eRjHp+nXpfA0c+7EI5z3dXMjEDmrHA0/7x8B4jiq+NcWDWNuwvMHsNo4p
yyszEc1ZiXmyZHwhu3XAPle6gHeXvbNZAZZRDGmhYZJmnqnZVV4jMsuaM8ei8NCH2UaEYGvQ6igZ
HHUx3ZYdtxqf7cCuUU20i5qjcHGdtGLXmC84OCbH9uz7PsadG9MFCx3ZdCsgn646Ww6srV8PR9VN
xRsCY/gNSUu3Fufhu5gUtvYbaxyX5KxV7Ajedhgto/LO3Qs4rpi5Ps3dfDv2faUuRwp91wi9Ap3L
rXU6HGHbt9XRPWztXAyq62vSIdUgM7KAxd/2OTSeoVDsXIJsBUv8fTnyQj5yH4rCaj4FBuNopkbI
vf5Au5KENfacoIB4+eMymLQMAOjuAZ3YZ3XF6YD2aF4e5zyB8n4KGaBjd4ut7h2iY2GeJLwWtfjg
XF/6QHFjD4DH/0b07jbuBAP3e932bbygW9Wvmq6VIlWkNfBu1dqQYiRlRWHq5y5NHpxJ0qBOR1IX
jEV1DSOJ5ZpcjBPNRP0rQ6phwSDpTxA1L3pirND8TJft+sHg50DCKubEwnGgDJGmQfogZ7tr45GA
ludwhzv6w1GE/SxCKSsJfYGTx9SuDQqne2w7Bs6JyIXc96GsWkJHNScvtOMgX5wWMuLbyXJ5SwZN
Scon4Dmg9eaJa592OZb32Tkpqz91oFAbilEu3muYUrzy9goxLI5/alr7r95sQGRgz0BQX03hddhe
F/hVlcbGQsYf3vqC8+nWEQiTt3GYk+wnI+CptPY9osNSJNnLeXjSyQBOs0WLT2TBkNlXqaJwewzW
0Zh6y5Hz7iTnjNrJdJnOr1JJf4UMht8egMD7B+nfo/JS3ljejSx/3OG0LqtWYbumuts4/RxfpAtS
I/sDpreoaYqmdQ+4G3uxBJDoXkZvB8I4bOYC79tVDpYYfPbFsenkAZtNIayCu0aG5cdjkc30z+bf
y/Cdb5kGZ5n83if70HJYurbpZshwNwdoty9AZiqnkdw7ayuRSEGYZirh+SH7mPv42/lIbu4d2fXl
K5SvWdYUnr1zKc3jRd5ub8PwmTVMplj13IQXFsWvKDDGRHm71XLOg6j0Tq1gE1YjZeuLjSSHV6DI
RS2hg5mW7jSVU5CsBVdYXWczliFIi8IXlaZT7yzYO6R56b5ForB0rmM4rVpJhnARWQaKUHbEUMdy
AvQLQIoiGH9AW0uT4zd7LkRdhTy9O09d5TZ4TPOWgLDO/FDVUaPpoBVrpqoDGewFm3D4AlxSjEgV
1f3qSnVGlUsacYTfQQDMycvqAWVbUs6jG7IBMWTVhgrjQpfjwd+kFgNwOcz9mpa16Cd8dA67uc/2
GlHuliwROAtQXiHrQK0jAJXzgU5cSpYhwjc4fMWqu/e7Ncxdded6+ej/pPY0bGtfYHHEY7kO0VBf
HENVsuKy+Feee/ZHWNa+gEbKM/93ZcwGyxIoI9iRIsbu2b+ocw55gAskAyTbNqypE/zLhNDY/Acn
p6/aLSsikCiQ01QNCbp483faWBS0P9wCoRwGy1R6XMD7xPrBMufUFHh/HZJkobqmX4PE2/t9Lw23
uSfhbKVWbC0Y9b2BgbSvTROZCsz5t1FIiM18oBaVIt/i3V7igOLOwkuxW0jOIJezVGQcdg/LZ/oL
qeXTyeqZbwd/zaxGShMWO5S/YFSga4mULocVNw05g25LWqnwbuKcLfwuWEnj7lpOJooKQBQPkulI
OSGhch04Dh8YQwPPi0S/ZmTQ0XgnGbKWzC7/V0edbQd9mT7tm2KjfGoHgm5drfXv5y2aRty1SE/g
kCETVVD5CSuSb4WSy/dkS1kAEGp57g/zYnzKbooS6j7YL+M5zNJdbNxcvwAK6ghYu+fDjvqAvb5b
0ffgU818+bMAOgds69IozJWglJgIt1pM5Uu/EvKjdIhYRJQvFuC+9Z4fI5r0ZoBBxH210NS8rv0x
yZXN7EHqbGeyJzACLXrYSm3XXy/sq1P2j4mgd2XJqgCjqcc1SPX8g0J17UuDm8KV4Oh6NJlYj+BJ
bz+/6btLDapD6PEv9o8/dkEyOXcNBiABAG9jUTJR2BhsotlKQzfejqeXMU+UpedoAUU8y3KuEdyl
Xf3C0pwdSw6euJiiuDmsc38x1+mfyBjqwti2buQnIfdSP+LFr90ko9XP406qhk23LevJ/9mzRIrp
NlX0TXBhbqOqmdhSwcSLIhBRlDkM781lq44/6bqNGS+GhT6jF8I72qo6cFLgT8PAW63dckLINhG5
pcB8mfgDK2W6D92G4lkx1vdeU3j8GmSNmdhwY3k12AJfMwyqkdpWqIS6LzCO641DCWZOshNoldC+
YW/xHYVyCE8h2CRY1DAIonrFGjZLye6cmlfGooQfiEcmb3lbX7QQBzd57/sho1kq6BHpKk+8QtYe
aZgD0PgqFF/bNeC/QwvzbAn01NEE+qXkpl6AePJqbrvznkFLhvJOJtqdNB9dUQbi8BoXBi9R/pHg
mTopLTVWAHGf9NI6FWi7D8dX6n/ty6ewfOQHVKdohQEi9Zp8RMUPKo0OuMYZjrd6zOlofzl+Lexo
nStCCnoexfRAGiNBMrzLCTC9tDNYM/ttlihRteFKOZVAXb+fXFDUMxtYcQwuwzHpY5ZSfGpzXKUQ
inFrnru1EeBRd22wIlTHO4Kml/4Qil1MpcZWgXSvIyzXRm1EP/Zo+5cRW5HDGOJfD8bUxXHQnbS9
0awA8ov2SS0G8KR0Y4X3xuP2TPc3XKTw/gghiyY3z4zbLcOtGCJoQocP3jdLR8dxLs5g5deNndKX
ngKI3NW92q/nb9riApNW9NyfodZJcb2pH1UL36uzC1jVQIQeLbh1lZ+Yl+eo0wzzlBJLxozGkDLC
ZfsxpIdGHByD1Wzgu0jP5JpoVNAXJcxLJmFqu0OK7QchvhCzLs+PaNN2Pp7DB0ER3ANjJkAJRl2m
soRy++vVXjuMQumNXbBvs+hkmUbqEaPvMBFgzIDUIueBtYm1XL7hxns4U8Nekz+nSit8jYGEvU+a
VMFCcPY5aq4PWLd3FDt9SLpLNXapalgXX7ZwhHSmrY4nVdotqq5lDCB60t7z82ksbRQUJV2eGQCt
01UZkNfnKff+DP6cN4DFsp4IscTsNsZtZ0HMRFQpPOM4/uBeEOCw3jPTWDMQsd/UksX2FyxjruxD
5JrMxFQKZMofRT43GIgQyChjvfRrl1HW9Pxiz3jqOwPXrMwwiRM0+uRu2LrmoLPUxARDOR/6WHrk
C49gghLi7sj5xs6geCwRbQ1Qs8mgdPh5uRSpxwYva3eSzU28SdkLV9v7h2vopTscMzwTuQKXHWwe
x7phqH2UJm+/W2DebssPa0jtvEGVG/LjB2le+Tzf6HPUECfGCiaOWPqL5WjELjhR52mGJ/G1Lq9Q
Fhd+pCrjz5YATPOifBbxIAYmlqyF1poxqqZNLGyw3SYpwGXi95rP9YOm5mGnVKtRXNG3IccnzR/l
GhyLUlNPv8eNrreSxOTrunZGw11Nhrnnub9YNHsfeujEup2URBA6YFpRIn6vHLnDMWhfvtQbXV1Y
DP21z8SdEj47qXw0d83l/8P20GA1kzwrKU7Vyje6GHLSkIDe+xuuOdfj+OSO9rCbLKR6x5k8U1+j
J/SC2s9t4AQjRofwG9EJvHVJVLCMlUXwSDc9BEhG/cAatB66rlhVbht+J8Yk0tcX0rPv6RLl6JTs
u8PaFoyyBAQV/rvIbGKfDVZ4Q94oSKLsDz36NwxEnMYUMkH5ku3HF4MqXfrFDyCOQRLb41RpS/3z
Fyhu9kxiFjcCdikA6N/aqV4dhVqdoPamob1ZL/WNbSJLo6aRfLltWMNva/4/tqXFG9h+uxNyEfLn
+sfn+hbwoORe4KZpDNamdp/yW7FjEaL2+9ETbSH0fi17Mkj0+G8TdPmi4uC3BbVHVDFz+tJqjAZ0
fcoQ8g6gwez00LRYOjnp3ouKHAsLXupWQcux3hFaufhID3GRwH42RGli3SSn/+ixkbKXlLpEtxdD
bLFE3ykKRZSwT2hGxjTfbyd2jHdCvt+In4LBxylBa1IoMoN492b9D4d3Ii2kOKt6bdJ6oNZrxDl8
W9IHswwR//n1NDdnotINRX7GInVW3M4emym8zh3E1jjlcYp/m5aE7o8AJQpKUGgmZH/NlTjfPN6x
F66Ar5L/nHFkWsSPCiQgnj4vC3CmJT261gC/Vbdv6sd9Qq64lJsuT287C3B3DwaVDv0i9auItN4X
OldLCLCEp9iGT6alRXXEKXtPPlUs8HwKqwjfm89pQkIfDDIbs0Jd5Ch5LzWyb2OxnqpleqesrX6X
/1cLUDNQXR1IAvzwy3+v1UiB7eVmZFvj2/0HkN2Oy40ny7sVMpydyy56fuCIj5tDQCW3etUl1Hg6
zPasdnwc7QK+roge6jwXWfsfwNLl29twGPM0LwRKhcQBZq/FgtJRZTI6c+Lq23YoO+5NJxE1wedv
K76WUH6ZJRuRCIjkmd8HBXL0QEOxpMcXYcBacmUxNnMf71gzvNWu52cOVF8HgtTrXx6PQK/BagmO
hhhvD68sz/ycB6Ic/OD/QmoRmvCduQFtZ/gyi2uxOcUx/bCf9tJxmW5WDKEMPb7eAzSkLTKKFb/8
ILrk8OgfxbCaEiu7SaRhHh7PBJYQjBnJ1N9eii+aWYBSTSFuqJ3OxNbuMXEqWDbeYi4UAbeUw2Uc
jRRM7Ro3dEXQU8SJjdYCPOm9+Mzy9MZ2KUFqKAGvx+76ZFHYHfiUx7oBrVJHS/SqlvkKIco8nUyj
XusYr6/hSUmeqmoDR8eMe10VjCaYo/OAdpCxK+o742OJX5gsqJN283FuSmLBPk3GLEaQDRoogT5G
hlo7G/psBO4uxT+2yBBEAgedO+eU8CsaDzYj8dwFBoqwiARATLMVf67mhz4VtBDmOevg1H84dkPV
7qLcMqaWgHWXupWLWpYbvvyJ93KUlaxPRX8a7yJs3O1ucEbal8UHajtkn8I6C/crCO+5Ury6Bb0n
Uvcix5wWXYY5pC4+UhI/FpobtfixaXgpUDonRqnkJl9TP8tDy3uyJqW6KFtyKLUIeUf1f3WWcqCD
d1BcEZ4hT3V+TT0cB5Crip5NkEaRUMqlgGf87PWgF+dtGLgMJMg5pmQaNxx4wSaRgEOgQ0rb1AwR
kLdEgtqQ3TkaXRi/BDRx5oZd2Pbf5c6qjYT592uNzlIY8QE/PrPX0NlV338pDI7TvwhEW1lA2jTa
0q62tYfPXLLqtb1wIdQGNnZB59EioqVO02fkkX7bvMK8LY2rgVXcO1OSYzfmHSIqx21w3FjIrbYq
XEjXdiI5beU9B+Hwck9d6voCoNIPtiNX+aa/cLR9yAdWRCa9TGBkkHGipFJN4Md8r+k2B2pmoj2t
R/5DY49MvlAP33C3OyZG6XJgEODiBiR/PdP5+ajNVNr5XWHm8W4SMNz28TQi9vamqQfzW43cjauV
0DAPQrcTsGIaeFwuOir21APM9miMIPTK1M1gWaZx2BJJRzApb9yxTwqRhKALsLUMefEgOi5hZ2s6
IO7i/VG08LmTMaTgVpAojIE0SOAXjSEcmAZZCrB0gEuE/cYB8iqsb7YXMwAIUrhfLDZywuPfN0FM
vLjsQsTDr06ImPIp6LtUcOpR1IpAI4PT/6DWBrlExK/qdh0NsZqU5HpjM3RGutTcZXAn/POHQL/z
1o2EeMMAqwT4oKVJHuyRfxdo7+L5JKKv3y3nZeBe7VGVUSvmHbKVLgc2goJIEy8H07vuwtTJp44C
XNCpVAVAFd7/Jq5RY7Uxt5mejslSOkMgOvA+Yl/EGqKjrJqpOPd2hKe+G3YXcpQERdEysdWVjq9p
WEJtrs4+kZGndL1Z8WGOdDROkMUkpJ5KY7xjGXmDQimLLv5FWRiRcYx2M7+F2jKyiF6elexqtExm
0n0VUrR76p70mgHC07fgBndLXfaALB9EmHQY+TKrXqZI7UaNq1c2028OTONJ4zQAeqqd81uUtLwP
Xp53TBQNmYfLm8FEgBUOk1hARxa4Y/3D2TOBP42EbUWQ9Fhs3BC1pc3WVjU5cR+PJjyGtXLpAEmX
6h4CgNLzYCKW2lmQq04Mci4OPiOpfj3LQOkH2vTJjBz1xSUS7hi66OqixYYFZVDhD3W3jeDvlHPi
HwDVNHKI1A0cw24vMkeIfWrVRBTyV/exuBE/ZC96IG2Bj7hI+qIgkTCs2cSVt/9/dKAHPmQAXK+N
2MnFl4so6JVf2FAay5NocRSP1j3DaQhvUtAWrO2WDpF8a5bOyHf8CEDHKvAQHX4lwO+9CTYI4Nu+
Ti+TAOt6APLEhALrdG9QWY/zLfz+H1bjmvC4N2+aEWszUSgTGlRqYzMxLy3wDR7bAMBxuBfXpvcB
jeac9ZkoqNbS7r4g2iQRLtBQWMRiKGFATVDH1KuIuglLPO5L4xLsqyPSkuYfMKh05Ov1MAluumks
cqGEk1a1Qr4Glh/8igyv4J9ZUUMo+qD/nTzLiarv6GC/elY5NdU7yfeJ04UxiNo6c0qs6E0ow7hk
adApdhzpekthrGgdXehVdS2MvcSMKGTfRW29J4KI3w2xz0frzFM52PCud5m/UvyJUJt473m25tA2
UzeV5Vg3KPW6HIZfLSwzkcg3Gm//PGMUgTava9pnscGJGT8jp4fsCZmz5xjZb+8+CFRYJZ2v7ZQB
iLyvja0t8iyUqPWrX8l1+GKdKC8qJu8CF8oa9GSffx1tHnuy1yb8vhcUgWzjTJy9UHrsgNnR0t+m
AvyAyiGs58EqRl6jZh+jeuYFkpZN23PXxSHyi+rO9nu6o14/kzmO7WSnF4xm6L00CAYwtCRxlpef
S7RWqVRDNICsOu9e+ZHEmorys0ihTHaiDpvDfVf7260UoeM3atbnLDNp8GirJOwsa452FaUjY+1c
OsrHuvdVzvLH3kegSHMCylwUQVz3Gazt1NQHbw3gWab5K/hLwdLc+B9OFcVRhNuygXrfDxC+5qlL
TolGKzL9feIyw+EeGwfBUZ+MjxcU7teEk21eqdozo4MD73fZZUJpch+2hvAAIOIFahuxaHxqASjo
TfwyPt+/3ing360qHvcsSzow118rA441suUkJBaSKukzKMV5u94ZvfQUMimjYj0i4O9Y83LpcEE9
X43DeGVzhDAFCR1HV7HaeNyLOwebGkTbE1D3hM07SQhbKhQ5FAigQbnz1iLwIMQ02F3cNjHjJIOf
pGfPPIC7wx3GYqfRAM8Kd8Aemgy4uQtDMC2dys1zatp0NKNsmOBF2iYwIiG5l8HOTNNVH3KxrLO/
QTAUShIn40PX3rn+Ew0cYT0CyrhAAYbKTUeK/k3vBblO0OEwOrWIagqdzRd/8Av4ZJBt7Dq6nU6Z
xcdfxnY/UrLHhU5XCvsGeyVr2S4j0w6SWnARU8naYb/MvYq8N5XQBToNgsPV4dSN9uHF9iPURcxB
m7HIrLa3AB3CRrYRXz/OmE9ayrGrDJyF/wgezuq5/Hj00pGtlxffpvhY4JnZts3vu+ORe7nv6pZ7
vX+wX4+0HunpHzE4Qs9Zxuz/5EmSWf55HRqHa0CjBZxBUEYEM2U4P25SZWWYO+OPiBSKoYmJXKwo
jpDl2xY15LePM+hEP4Z8wyg9SddTd6c9mofQ7Jqay7oh9YwIR3aOP3yXDVVqwcw9caIzlFGCfVpR
sVydRYgYSHza/0HQXPdeXBxXOVO3qssM0cOjbhM/xodLWYOJpFpUDQeFrru0FCmgEhqrVCThT4TQ
98M3fhuXH5qbU3ox8L0mdbIZwQHM1AEz8iuTsAa4eqileQlpuMbwFcs9p3B0eTHQPmj7kyzAViHZ
cYM5ZKIob8v2E+2mFkta2hA0cQjQ59Q0aVKt8ReIFIKZLwnL3JVoj8OTYUjMPdotzolCPa/1NiTy
aR0RWFM8x1qdoTy+24Qgy9g5XJivD2AhZfTD7iEXtr8cnhRb+PvjBCb5QlpWEHJKy0bzAKm9C6m3
ee4AmKELPDJFEGoI9t3nJqGsVhu8jg96jB8WeYWLke+M2hjtpJOacCLFUhvYyWYtGbhxXkFxtO6s
MQ1JV2O/4wBD0kq9Rr41vd8P0+JG5Saa6Bynh/qBTRUnEfWDGMolXGP2ccYdJMwWii/o/kN/XhdL
/mXDZZFOSskKURyKpFx7vKNiGanZxtZZF98E36bhnULB+bYes8+cdermIEMYTzmI8LpXitgcY8Ld
kn2+pYhCDfvpv9Q38oLNqLY/BpYI9mNms0yF1Fl//rYfF3r81vrFXsP24zJzINs5Kk4eh381X39k
V937ReIMFbCcDGZVJLDoD9haVsnDb7/W/tyq0Z6N1qmF7uHcniJO0P6CFAIh4rwN99VKmFTeA87h
UfE9On0bqXy9GQSSvnOW4u/gxE5DtaXyBSPHBc60WZAnghR1gi7iKvZBCTQGaiV6xMCgTMvcZToT
7owi/0WMXajdBNJU/MsxVSX1Dgc20A5jb88UkkWrlJSAEmsbGcska9eeA12aqwN1MP/FsCVvt5uz
5Yg4lfm7w+/o2CbjuTxTa51D/0FsxcuzgmDcQIjgR3KTTNW67dj1m/n3/4M3lPocjaNSMVMw+q0e
s7ZVGIdV5//YHBNhttTqCsl2VVPFVhXe83OSm7cdNrdgWPNKIGivPDueuXLrQeu0Mu/iGrOAQWTY
nRnhEWWaxHMMIfmZHjdgpm8gg0ydaaeURSkt7g5GuFMqjy8pWyU9J2Ypj2Z3ADvv3GUWJpfAiUaV
u3xXZHHfh6vVOCOANNRpZ0x5LGQhO//PJ6ppCaFPviROYYOpFEGOU0PCpNO8sKPhl0N0sF7Db3BB
9dTGK9nyJozagAmFxfSXp3eSw4Y73GjFZn1pDPol5fWq/aPvozGtVvyguNCVYdNc+gMpi9Kbjkrt
fl0/hobfTyQxMxyleS7eCTQKeTDOSVkENOLCxR0Hs1e3OrxSBhLLPMaf4heLPcAHiYM40aesyraf
y4imOCEay8C3brCqoAeSbHiE1lzAdLeOF37yAncAvZUSaXyFlJeBdTpkqcCbWfu41rS3tzxuacuf
KSRFRgP4v5xzkdjbfFXgnxdnw01q1YFBx4D2DfohZ4CUPjCXkN7Zyql5e0CzMVtLMI8ECUqLAE3p
kbEIB+F6QsUq0oCnvWp2+lygsSTYJK/fXVIrhlIaYW222ZJoOdJmboHX7jtqp7aWjievjLCjFlYL
DFpkA3Wmc2sU/43YZJMPLumPO/62E5NX8Ew4uRAWdavCXY4prwtNBmmav+nfCoRD0zpkpE07ozKq
C1XP+PzWgDiNMVR8e8m1ctxjQmHaid5gk1AYOEOFEYRuISxPl1M4C1au/v8WNhW0rpFu726oq3G5
51IsH1f5x7ywrjNUMDF6gdFye6WpndfIwfuYcmlpc6WT2LR9e9XdxAivI1sLvczbZ54DKiEBkSRb
DB738Xl5tP+wNpBYAohdS6K5FB5wQM++u+FF/kc6e+uJDxzLxT5iSEuOKEeVowiobVc4tfcE36H9
AVT+8hV/C1+VJMZplK62YIKsNMZJ03P48dhLE2E+K8y9691pkiV01YhOFJwiLncBqlRXP/q2rhQ0
BaUFtofbr9ycXQVYqXVP7Af/745OGcwYa5eal9tXQyzyasEld6pQ4XW+ejHVEXGUSm2uMoAlLE1D
rUofcUMeCmD30H09nWBklHCPUKcdLrzVHYwXw4Q+QF6d9Ebh270ypGinwbACpm2DYLZywhca1bQs
bGfbJ06N6ce6XV62BqBiIQpTmaLTWBybSQg+eVllmnmLCTtrRFxAtC7DOmVXOMRWulexz6KjN17U
dBYv24bM015sNWFoH3huDt/VxRHlNXoQZd3cSHpZn+AebD679c/vTMRn/+ksPJnpd+oKKlDy33MA
S0ShqhJ8MNXxlyL6K4TQqjLIa3vN6zez9kTMbmimcBb8OoXUwTErm+tH1paolnnktXIb2KdighIQ
9wTJUttU1UVXNrlfsqg/CFz3MBkzPWOVG8TjH1pwcZ01RMTd27LcwV12xZoA6fEpt13ZC7xLVKLi
qTLtwk3Dquy7QdgcJTkq3Ri2Kd20Js50g/6bRth0Mw833ts6hpnoOWhhkV5PoI05N9nUCBmnggAG
fbIA5JW+XnsjmWf+B2ESKiPLdQvfnR32VPGTUhBIDWliDNokojDo1Z5MlCBTL6H2tig4Ez9PsBaG
95pDgkRxsptHwHiAmXSuKSfiRak2wssktY11Q8ZVREMBNF+i6TrjJys/hj5FgwnVI1zlVeIJg93x
faISjB6n/1HtJq2VyMsOyOe/F8Mbs+xbRDjnKC8uu1FC7L1GqH2F4S478iG+Veh0URmHSymRcUtw
R6Gf+Zc3YcHj9TMErMANfzrlMa+mV3Z5wV2HFYt+Px76o9w9ycwwi2BagvCwHin8XRxhhb9x1+qh
0lRjfVKChuFuNVdYwvwZQCcmhOD7wwBqRrc/zFhXIzqLq9wO+TNECstq0tSaYXtTyMz1PG+2wHq1
TM3zdLW088kN0T5/+V15vh0QzAS1qF7G8I9qO/beYoqyBLp2wMNmJWEuKT3wvpC71FHagEYCt/Lp
LRIBoQDX9YnkXeiVAvlTm+IcAO1ccgu1xnxnebQ3v0Rp+1rae22EomvcZ2c1GsEYZ/TC4oucuOXq
sxC665VJyA9Gq7/5u2Pi98sA/A7eI2lSHzl+w5mu+ixDiG9xXXrTR4LWvRakFipYbqXhFZR57vVi
4JKUn7QpELfFNpQcmj3GpjeTrYrnPJVxoqUPV6K2OwgDVaGW5jFmkg0XWjNlwXaMPC2edrVezp6M
140LNyer13fZ+GuxHkBfdDCHyQ4ts8uyeURIcR26bKKy/2q89xP8CLSonZqFQOLjhy3dI7iOOvFd
X/zzF3xzOOc3pSGL8Y8HRtQ4mkV1+M9oF5/bvfJzyCunsurca7Md2ErsVdGM+4Pwnahw7WD0kQQ9
8mhyTExDsA2m/JgsLmFRtTWKijGqZQvhXqL/lllTE6B1B1GVKZVYY8OqhbUQbqt8lBuktEvlv3gW
+sNHFTg8nGAl7+LZPTHtAyd+GujK6h11PlfaD70HI/5mSJHvPX3sJwUJNC+3j9HaIsCIW2HH0mL8
3vhSwgk2q5uxow/Apc+sUqiW4TMyJb7DK1wu3VYGeFJrajb6tw6ObUFQMCR8CWMzwQ24Jq7LWoIE
OvaZHuRPL5lJavlgMy5bh3S4ZULV9k0D5vBeQUK+jkv3CEsu93cHQa3Sf20p9W0UMNqESd0A8yGa
j2PEgv7Vr+31JBDIcPHBAvTnXqsnvTYRu+WHSDkm05O3dX4tNXaePA9iZEsBBYQytQjBnZIAOWv4
MXe1Xft3cQxaX3mUFTb8qLMHjrRo6Yj7TuWRDDkn2Zk+OLoU38s3o9WgaiR6mjpCfCP/akKmQP62
VduEAr2+KhRp1XNIPMZR2l2f48KMiEJw+hS1ROLo47PMf+xCwzozrJQMXoeRJXgaROzChER3iUTt
S1JmfNveSuzSiIRh51zSkQsDXhoxRfelA2qc6Y3Lshsr5uY3+Cx+iZEFXy3fSYzM8VuPMYR8u0zt
ZtT1wXvIo2C6rbgaHDyy5ENE2lwBlIaae8XiNkz7DdPm4GCU8AUAEwTeUYAgKhDP5mV/QhIx+deB
6jJn09vORpzLYhrvc6fOgwQSQ9Ih8GuwEmVhcXXJG736mF9UoRIHEWsgvHqDRrKQj+Ul1pXNgRU2
IO+V5br2/UJQMHkR+jGYqyWFRzUrtr3q6Cjr5YmYIB6/4F+Ygr3yDSuEEVuRF/rZCiOKDJHkR2vb
C42udfQ3YOVJgzayJfL0VrY33jiZXuB/fJB9U7TBf+U3CqKetFhoB1XwfgdXnhJcs6C787XbdCQt
p1s28r5w8KTKPB+/3IUiFMg5QmqsPTtuKeCve2uwQF2c+8T3GWlUOf0u40WG7le9BjuQQVWTHhDC
ljdHT/exaZK4dXkcndW+TrejV18S7IU6qYobFuDx+fNsy9r/1SW5Xyi7AjocwMQY/nt3aRXdF6QV
WUYTVIr/2cPVPYXmXByVyxOQ39/845CBrMmqJaSFLmNUX9JD1zZ0ntCGjNfRVyBbn9bTBmbSsvSY
U97EZyRUwH2XKemnhYcAETRLMjoA6cyBRX/LIgVTzAYP/6vitYcou4C+FsXp5c7sFnTYmmUHvQtU
XejZs2DJKievNG45LwqUk4iA82qTOm+lr4nWlu/V5JxMDgro2S0SinBaU5+IUmPbQLgSDX053ENy
nmN/tmA6AgfCh/UQK/ylaxF5YmiKxRy4CmhOmNRXuV1wrayrlvSOuKSwdkfgvJPi/uSXMr3gW6t5
UPEdoBXay5f9GnyNAWsyU9M/RPeB/m+wXNU/oUJDCArgaGC8tik+OapFRSBBKh5MgyZIihB3/d4W
Esrivg9tuLL6eCn3HOgabMekS1pMPfHjuYGhOcJc/UJAMVTXzb0R/l7F8et2ArkPE1K0ufltcUHV
2U+WvblMVfJ6Y98FE5wekjEzqIXhRSPBbYGNzyc+BK4qsCID6etBWJ0BaSHzAK+lPlol9Cz7GEn6
GveC6yyZ8Qp84Ma9E7nSCyPNg/D1Hjg+gJnZGa0VSvKGYVrZ2XoLf95HFnwf4ABNNIEdEAv5iyz9
OQqj9yYOr24HTkmw1iE2fKS9ESGxtuMNBEbTtS+N3aZwc1v3HACQ5OxcT4TSvDHUcaSE82XkXsT0
myxyoduaIkAEMKAeFp2M/XOQON9krDW6ES5hzJ9ghec+NUSdt/e5S+RtpLkaJ/DZFPVNkoGEGJmk
xlf2W8n9LcOlqY+EI4t+j8385c0MTt6Z3mgGVwhFljfoTILC6g05SXs+155ien2lSaB3+VXt+lOV
AQyQ9SQenugehHygGEMd81OMSxgXSRQ6kZ71ulxCm2nfGuQK/R9NGhA2BLSNy+p6ehuuhfdaOtw6
FFfklHJmcXthvcZd0sReVmCQUQOdlW9S9glNfddUH/mKNkjGalIVcLAvT5NkbVHWeUzu2JWsK/Lu
LisrWLoBJ8HFqrtwGKMAkEW455z78lK7AOk5xScs6Kla1wW+1tfU34mGe/LTeN8vIJvlqJDhU+np
7JUPJ3LfoRDZPn8UFGALXZNwv/o4BNckh/laHZdAtYtfWoA3AvmnluqvKgIDxXXGYnS2Jucc/JGk
X2LUiKxTelDBWOznKWVJTJuIM3e2fz8myoa5l84453jUVMp/MfnPD6qVEl75/FNzpxjHRW5CqT6S
ggIWlAXsIQEisVEI9sxAN9IW9/IaYGUnAHa8TwhjLzNCfejMOO0EITmsioknyXdAnEO3GWhpBSR5
Tde/taCXsQ4L1c8qL0xEVXXJvL0i2/e/gq253b8tRFK0PaSHQ2k6mmJjHzwW714r1IX0FkKGrL+3
NSuEYPY24fmw92MSQmHZshbNJuVu5TgzBwSydui7fy3+HW5EF45xw6EOghNf122uqiKxJd7Eh+4v
VoH6BUzwipvVUSDschYJaDDJ11zPKSzBqxZur73kY9UHlYoJLaXr6OvaijdrrgM2wxEClfhB4C9k
/tuAOKqC5d4MMpip1MnJkbOnDHG45A5+hgE/RWc0p++XaZSmA6V32H+6IAs+Twe1gYXjWyk+IPgP
nOuOzgLGBUxBZfg/BKtWNixUb4IhuDKTW8unHZSWA5DVIDtOXJLnb5OGnEvqhnwlDNE7+V5w2BoY
s8Sq2MaOHkgwQkPvl6A0NltrvAVPwNO7yuAjrybfGyY/Y8UyQ3mdEqmFT9JWyMx9etN4vbXnoovU
j/jNX7gODSh2DC67+vLYoRXtpr/2p++L2fHdC478bHdofkB6PouUA9cxaZUNztBAgzjRAdIHcOaR
uXnAL/dEjmMHF3WMn1266LWYb0h4VSB4T5l8Hz+RcBLH8KbyRT5i2IV6dwYJOqj7qwnDPLv1c1MM
GZWKNOcb6IiX6b5dtZ+h/mMdjH/HV1ehUlmB4TropeuRLHdvH7HB8+RdkXM5nsg1Zf94l6I9ETDZ
/j29BQAMLAnm+bxZsdHo6ME3UDxC4BTJkKOBYEDyL5arcU+BxhKRnQRYG3ehz0tgENR7wj+xTzSG
f94nlxpi0jbeQ2CKsAts+8GqbmGdRiEn+1jITrfUEcW9y1rz1kNEwwNur7JSB4l+UQU/ewZbrBAH
pDdTjS5EgIMBuEZ0rxn58O60KtQKfWXlIkWudoJP3N39wwsxav/lN5PrIlorV/ROnR+VHlzQrgoS
j96RIM8dzuBuERT5le6Gb/zHjhmzCRkKuCImEsyyfS7nm65g7XCl137Yp15qaeC4O+rYNO9NqL0O
4Web1S3wK9pSq7aH8ZeaSay6rvWcHZdKiTHSOHaz/LCKqeSQAymDRWHUMPvyijfSl4xoxAD4q+Sj
0VhYeETeOYMv7Lew+2G+FBIy8j9RuzI1BKxd0zIsln5cRUwtxf+Paw7ja5lgNXLvFZBzd9N19yCS
unGzHAWAhSjQAPloudosAmNPMBHepEcxctbfj7mk3s7un5gickBn/m2zVX7ttxGxkD0V3XIXnSd8
o7m4lIvGn8COvfmgcHpvg6LjE366edQzHfCuCs2TVd1s3ujuHMD5XP9VL2IXVGk7TZcXAw1BWqYD
jlIJ1ntthtOZMXs0OL+egSLgk8nH7GN4H7GCU+NnHBpU4iXWbe8dAqmlZbUFpTkKFhnfN+syPsUC
jXAsJbEF0xAbLWGgWi+TCd9HEPJH4Gt6aN/av3pQUOtW6PPtrpP/ZvewGvOk9fHrTWE3J5TxkFtd
Lch/islW+PCuMVQ7zfValPwryex29EiAB1lzg+d/ywHktC2tA3+LZ5vSKv5vh53hwPcpC9+f2leT
asiTbthI82S8jkSqLNiBHRI7rx1WUxv8dmPUnitLT774KlewNlnbzStCkcVdDvPUY9ctbI/+r7Af
J5x72lnqlK2vbbJ2P7BACOUMtknwHyJrochNoue//uYmUicYUqgZnA281M/ZTQSA9CpshPd8c9ZC
wNHqoUShNxAp/cHn/whn380JvSjLGZIOq6H9I/9yHP+ZwRL+qXqegbV2Dk0JRUScAM7tIjVMPA5J
rQM+xG6/Ld18fQ9nbmKS6Du02w71W/6vSCRzKndENT7oGW5qS3ptxQmX8VDCf493ZOzxRz2M7LWy
cBowM23Evvp39bqU0MWS2SbM8ifWESP38duZ3Vukj4P0IiOVdq6e+lmBToi+a7euLpnBEtRM8xgV
lRa8RS8I5QyD7rY9Vbe6Nv5ua1Z+FTdOcR6Y2sSwfFNWpNnbpAw7aguMlbouSCZ/L0YK4ix9Smhu
VwnozW1rnsldW/6wn28YtLOh/K1pghW1d/nxW4635zjnbkhT97NPsw4A9vvAwNEiGAZURpem6SQM
2YZe98jxfnHzBhBYDv62Hsuqk/Ahc3ozQmukr5V1gUO8vnv+VBW/zmdskJkLYKr/CI3KX7mPfP9G
QQlnIFHZZpENB3SqlkVrTU04guMRP8xgZf5UmrqAMryLassinaG6RN4aScQA+pTVjlDMcHp+OXJs
wVMUgIjZ85Xaoa+wO9hn2RuxlYJwfTlcnMurWHMPZ3BwxbGvxLZjkAsEWlAT/lGPERYlCwZQOr36
uruMk60xw6FvGAkPwydAyO4nICY8ah3Td1baXS/aIm7cxlEU1ZlLzvP1r/kWaBSEk6bVmf8cBtDm
2Slx2949P7BlMntLgJs4jbuYF2LhkeZTuzTvQ+hAxbvKJ3NYTTxjL4zythAeaFSWp7TQWlLdC9ia
BXpf3hYS9oHysFYze+zbd5bbobBKDa+o68nKubg/huP+pAbxxyz2OOJwcOda3hz+6AuQHmar+4/I
7oJEyP9iRcZEm9c4JcJP31BkV6wYLTCd5QHoGgoLp0tvywnKhlsOMBP+z/PzoC/cKZdWFA+14WkB
ZKoaxqEx2YvenglOP05XWQaUJm96xE7bPhHp8YSbgdcq0tHkePgeYrXIT8sCUqrCmXgF8ASjfByw
by88RnQT19oVKN1VRiHdud57wXzweGv6dq3NtV+TZKhRQGpZvgHT4Mg0i02U17HsACnmjPD1Kyur
eSQ/PaV9vXhIjfugEP1BpORPOmFYz4YCVO0WdIHr+GSR/QIZ1WuGJRU7c/0HMtvqvKdul7ni+0gU
RPV7BXfyOyx4Zs1OZsWcT6Epj1KHsWr3eOwpaLRQeMjME6NuM6SAt0rzIRXno7Xm4Lr0/bmy07Ah
4DfPPv1bPEKbaynU5OXa/liLEeebeW2XgzpKK6XaRGSlx0VSWXGOVuM/NRtNonHxnYRo8O+qtEfM
dOccwc70+mlsqO17NQhf/IZHHra7EW0LUqPX8BJe4mKA3QMV9xR/YfkCoUD7r7sZxLmdYfQIW1b1
LXIZ6IMdIVVkGaooGxCV9gmqINLOTCP/MOFklLR1WVIYAvO7/IcWNet+CRfKC5HKL4uF1E+OlzNy
TkO62G4aHRod3rlwrzCe2PZbvm4WSE6idA8OXCTPrv2pT65cDNLO+a5Q4Oyq96T0nS6mqq80AIIX
MO1oLLl3t1/pLMF6K7yfq/Hi/7CEHOeWR1+YmBaULCSzS2aN9ehuxbgewOVDdaGS6Ak7hKlbYAam
LiePJo2s1fvHM2QccHWK3fWZGcKBCwoTazhrr6lUUz7yxWbHy3minsH3Z2nC0G7W/+7ma0vA4g9o
sJeCNmIfvH64dQa5Is7lpQJoor+H3jxGq8Ayfd2GLekuVVPKG1lFuhtd+THsGsZUEWCN34dffEux
7Yhs7O4yXKZ6d8w81KSELYBM7sGADyYaHAKSji3yzhh7N6+e0xLwSdm8SOFYoykzm3qed5efh31F
8HAMtotErWAwXM6FZT2c49WKoROpsvMiRijEfFewi87ZobGOKiLOGAckhrPqjEe6vazAs7XsWYk2
XLQYIDu+uocW9Mri7cHmZSXeBe46fVM+TsJFNyXht8l/6uzcDkInluzr1YGAsIvMTd5XBuvMEg+Z
Jj5cyAZeBsdt/WWv60qPoO2GQx3k28aLJN4LwPmmSvPFzFuHU2zsic6iDdljn5DkblrGWagp0Nij
mg85lxuFkKXGTw0eHjgQkNVwsan6XiNem/MZkBepBlVbXkjBGOG3oSw30OalqsLAufI0AH5IaXCf
Mqg8be1qpOlGCbNaT7YzwNnni3c5xrYT/aYEBUzhfQ2H0K9Nj2lpssgHPvGCLpaYVWf0Yg6MZgPb
iu2IlN+XFKPzFJi+A9u0H/H31b85IlMkoGhW/+PlhnEgwAWZs7iCYEq7qc0rcAuQwo6mE/xmnFdQ
Dn36/wyU+lEGrfSuNyKqN86aFEmRpAQi3GrPHPVPxSscRJ1mwh794NLqRrtOmddyahvXh66tteAy
TYKdMBIDiftk9xztm76tz/EkfIei/DCJu3m/eiurC5UPxNRgbg7jP/rYj1XcqbChVJzixc2TTKK3
Q7eOUiQLPFxgBzMknCEDUmGfMoB2ainWoO9dRVgMH966aWyrtMsXZOzVa8RFJQKlIbZ3Q48YInRV
D9N7LgQQ57oTKBoKYM27TPZr5fl79nHqbgxMtGhRGPVwpRSKLDu3d4hqWnYkO8VrTAWsFYEvZVhQ
fQ2PuiicjFFqE7ue2JXJAjmatW05aB+6I3dR4fcaDCu2/+XERhg6rK8weN3KJfA1N18EW9b/bQQy
rq2/7l6jegInAdH0T2T1DNWCorc42/uLf5y0Tu5nhJeUgtYW1IQ9Fg5skn1sQg8u6CJLo0a5sC9u
3M7emr79cNQStS2YIdoNW1WgTUa+hvAlqMB1NtZIrmR3pTeUghLHgo0YCAbdAyvROTKUEQYjT33A
Md+pp/6qdtSVbhU9wYs74AL/YkrLOzjHGWrNc8cuWl0YzKFtjLrArr2RAs1Wa8NKCdnGTHT5sfzO
Ck1VkmxWwO0NZUKdfqeOf8UyDPahv8n8nlGHbBcz+WXG4YFSmCLukD4eWrWs7pNVYZtYTth/5OPO
dsggpbrCiTzm6D8msGRBwYexrhWm7HHwB3sGeEJoHTYEbFXeHE4WhbIR92e2xVpUcSmKbmbiKYbc
frAw5cm41hoSUGyECsmdh1Ty2O3cn8tyQgSbO1hZihp7m0J+3rA6BvzcqNfdME//P0OqVdXv8WTF
aFHfoXguQu0WkMIyB5IWlXkYzxumA+0HCDCNfMRkYY4QhSv7YrEikBPBkugMaLv9V7fKnBfKVLSs
tFGiy4WNjUStYNNlqGJDcIic4tKPiEFkDojiF4wmHCjtj/sPzeEwGIbV4KwEPPKQmLW+wzhNwRg3
prxGyuJ3DlHPCIipLJ8MBKkG96ORo/9zXSRwYvc6nCU16HdKeCGggUP+E6mOHgF12KSSHLVYCXaa
Ftk5BcWxsoVUZyPNGodXOSp+g6aldQhZk0iMxAAlLlOlHa/AyZIJB0AFIzOkI7bj5XfzIzsDLOZ6
EpKSJv8oQZoLeLNXpeCiMZBCpPSskwp+2G+cT5R04p5SokGv+AMN47iCtSP1h5hy8cCFIpUmjdrz
rTDqAlMAKUJ7OSIophBq9TBoiuvwJTfVSIAGTMdiC16b1jcD0YMpw85QRm3RLAoKV82T+WWuY0Gx
hyF8kpQrJJHg+nWD+blOZLmeyRqqpMt49iejtB45/CUySjYJ8O8e8m9sqfU9uwMssjHNYC9oNHnC
aSZs+JFIOLnFQuoOR6/1mZsQNpUEzapx3jBnwMtVcBdbZyc7LrwZQLb2BT5VtMUDhLUQL0/r0E3U
DVp4gM8Dr/6XE/pDL57KU+Qh2lTO26tZmIRJ3HfFd/o4B42KkCgMaI9MI9y0FmZvtsHXjQLRgYJ8
FA3xWT04ZQntBBTMGnQq5kPnLRknXa4T+M9/HcWOaYAVy19FoqfB5+iPQ7rmCsyy/LvGRhYM3RzD
I9eN5lE4Oe2j2gmz+WBqAIi6yP0jm4LCyrLLrrc3wcD7eO8jTO0ShTOO/Q4dDIJq/KqiGKh5njKr
NWCOtRPefVRUqTLxI9q6bhttjAZUGaY2u8bF/N+S/qSueZcgFfD8aMi03wXzUYtFRfGJ+oXKcogk
BfUj2Dr778DvuMoNeY+QnYkjJYWv9bGQaFal/gc3pWwn4VdN6VEk4eU2UjWRiR/Vk/mZ3vWZJ1Kn
soygLVe+8rjccETktqzgskFwCO2//rl5dT+paK3oB7d/e2DJntj5CxjBuj/W2yUTMOSBfadt3rQN
/O8e4r8AhNvpaJPiLf2LooV3WJrWXTTefUKuFeps9wLP+1mIpYPhskHYpFpFsHSR5dRzA/WT3l0W
B3GcvNtGOUi4NdQo+biQGBIynFbV8iMPboQER8HTvs9T/wRRzc1NBhDJRqc7le69EWir+Pp6p0X2
YpBPvYBsl2TGa3S/EeSLipFyo59o0zqZGaUY3r2pRO/QTCpbm6YhMxx2/I67d+cX0Gr8NpdKcA2G
NwXEDCilMggoimFHPl8eh7RHwaVrxB00XDF+1FunJi0zbDN8QtGXyA93Uqql4CDWJN04MatpH/I+
qJeSaDVA/liHfY7pVnsPBI2QCSINd1EBM8ncuVlI51nuFf+t2bTMHEgacT7J6GDkj0965HAhHsON
dAqgPScsI7NncNgHEPLVw1pjbPCdFiZ0V/uPCzC8PLMje98Ya6oXniuYYpaQE5CuGNGla+VMj0xL
UDkSzVKT1RCPUXnVs3PoR4bFro93Sbkjbp1c2pCfi15L1v5UqLSkI7ZVSy/5Xr7cXsf7Dw1exWKJ
Mrse3a+3AKc0DrC2ry+IDBCH5qMGioo6Z7qjTlwutkhGKqx1I4MCXKcfKxYtuv2VcpmIhFiGuvAS
aEIzxlXCW32zWar7BMOQ4ehRtwnL4XSo+02xVNqxIdMu9e9L4uxqKEaPpYKlVmzUDoMLTLZoA9lD
9rWnWzopmln7jYZqrXmnq6gr47fDWykh7gsCKQd1/Qi4VOIO5PUimqwd0PuY1BQoihyQ0HvxKM01
wTJLapvJ/gTJHtLziN2Cj6YON0p4N/MFTo/ou9r2GVIOux918Pw0vedMI73xKayUiobx+USTpurA
kQbqINSCRMZooxd86/9oPDpdfD+ZTSnSBtF/ZOKD3/BGGdLbysaYUMy7S8hLU73m2praWFQfOekz
Psa2cJZGguY4k9WOu9R5D1mabTEjDnXFqBzzDXoVK7Faeq6qFuWnb3IQu/2xQR0h+8o5QtVlCw+h
kUJxoUs41zamQRqblYLPiuO9bl2GeoGTuHQUUSjwVO2lj4yHyx5NEpNg/OSi4cflYL2+3hUcWuZi
ZYDyu/87ralnV0ePEcK3Q0Z/hqzHFeuuKVBZshOL/Onq9QfZIlLNcdJuCEVFTwLnyFee8WAeachb
3km104f7hEyea8naK5Iix4J1DOrZazy7A8YD2FFvhzpBKY89cabJEpoCV/zPD84tqLjk98f0g0ch
4vNybKiK8kHyXJ1d7tXzHFefqH3fRNvew3TwLm5+cYqdCCyNn9Mj7wSoZUf49Dgz7RVyy/XVsTPL
YXlyyjnMQ9tdJQoG+olA0WtlWTZmHoUQvUvmEhYxDt76PlGRoI02RtIy0UxeV1ZcCqC6HpD62j/k
Nph4XxfNCaUTuClTQV1iZp2LTL+KlADwISr8ND2TF+/+CEM7uwZjoSZP3ygzYes/nJlGUFnYR6tg
SPbOxTAV4r9085joU27v8F8p1PpsHj6wvgfpTmq4sgvh231qw2fQm17iT9yyzy92oZDH+c65ZuRZ
58YawSTc364o11vGfOL8qzUQnbe929QXXT3g50r0qkW5A4KdQXDrlRf6gJ56ug8f5/keSDIUwaBk
eAKNKYIu4IH7ipIov6LXjgimxBIO6Hf8fxlMRpk4Sw5N4w+8gyruorJpzYBU8vgihnZcldal6cbc
CZJUyIV6LWDkuIgiDKmwX5ht5aBsKoBwMNfa7/4CRyVI8eoZJOSu1tyHDPvG+mVtt96Iyr3J2Eq2
EDEM9hSNmScRATTrVCyHN3pjFmXOIJC0pOdAZq2UP1miSZdvPRRA9s3IF9GAr+b3N5LLZbFGiWy9
q/l5s12RCfHFgT+vUrKM6X8L4N+OmsoqDfr4tVMNfklochZe5c6clI2KM3x6aFvVK+ZffI7W6TtA
9hFW/SZK4csvVWDcfE4M4xyi38m6LVAJaC1jwX0eqPFYyjF/rrorPyxNTa082WzjD1GQI7EhAq9r
FjqVjITg9p+WxxQNVks0+UYsCv2UQEfnwwuMFTMvHImlIaMyIaDYSjnNnyePw0tbXp9/62eUkgXX
dDn34HS638uYPjA2O6HZtI3EJB8kgJBiZsrW+sn+n4amMfuL3vRAzwvKl74RX3aFqzXvYVRpVW8r
Hh/LpKoQUGnaDNrnFIgauzVp77cQ/YAPF+XLc6vmErLPxxdUHcfef17w83iadhrGKsLZdS8c8fqw
Qv3KYW6MCset0Wtd/RqOHta1NMAjGm/wDrSHnfPhOAIj1WBWvaoer7vEWC0Zb2iYr5i+8YhINSES
pMFh7V3X0cGcANizbo8+1IqErAVAjLqZ8Nx8gvWjxnBBwHJvibsfcwWfXoCJMkBPH/WRNseJPaPh
pcoU2r8JNCiD+e+UZI28VQ122bksczoFAyq/N41x/a67m+KTPJBevTZSbZ4yqdIsLBzL5JGDWWkg
ZRpe3M1TIyheYZLn6v64v9TXq8rMIYt58uY17/CNMgNBRpInaD66vXTGW7ExiBRLNxhLMuXI1swf
IIqg77jHmsNzjF2/ecV+Wx2Zmjp1xwTQQtc3tbo/rshXawR6DDwdbkcoW5Qi4kIGyBFiHaVDu39s
Iwl1Uhs8v8H3hzp+71Ak0Pqxm3+kenyfaxp4wOiLLospyF8UlvTxVId2A468bmf2w8KaBC9C3co7
N3tLVxiKn6rGdo0pBS0JAATKLY2PfYfIx9tKQyDv/hPWKRPyMmnNdJ8vH4FDupsonF9X6TZPn+vF
uPhhURxkBBfmnj8xIwL0rlXfxD3Lo28252/7bHN06XK21w5ZO5XEF1hrtRuQ3m+pHxlsaElfHaLe
g6qP2i9XSTowYRs9d308isPDtvIJ52kRL0AI1+UXLHrxtQqW5yuVyljWiJc6kX5Kb5Qw8cwfKZAD
3JBFWSSg/ktB0oL3W4tSa9RijDOs87GOPo2brBnS1/4lYY6jBRsze4TVJpMEmpdFQU3xWZLumEJo
OrMgHXENiXnW7D+DgvcKdDFr1p/1fTGTNuZxIVNYcE3Xx/nZU1ReV5nL2wBei5aiflsm8X0D8Tcg
+z5Ee8VuWtDSqJs8TSHRrvLmzGZyV50WGDj4VzuDfQNqWcjKQZV2HUTanHh//ZTH2p59Ke4ShxRd
XZSzX+NCTJHc1mxiudtKaZOdJz0dZxb/R6Tc2yWuT0A6kZmboB7EwgqgRgv6h82PTJFKCsI7LMZN
ikx7Zs0M+0Sv15Z3IG4zgQtPks/NkicOZq7f8iUWLTRzsHuH+YaXADBeq+bb2FdPtk4K3ZvL7j2R
5pGtYmZUz4gJ7+t2S+eaHWMdqfUUBGfbFLezlQhdQnQuRCjP+s5mSYMmY2m69TSkBDJvQHa1B+lZ
ikLZQ57OwkuMiuXpexXEMpzPWrVVtKZjvmpir1C/0cf1z0NS+1FYIHDPichDbysgdgxJBiy3PNJH
/y9xdof0VpTZA0XqvvKg3PMdIk1tRhPniC4EfdVWMwRbHOZPOX7k87wTymXt6B1hX+ZKFAIguYC+
Z+LyTlBXnk2AgCZUYuWjJQgyhjDRnXolOmwRTB01Z58j8r+PpkQeMP+43LJQLM+DOaEur+yQHAiA
9xeLLar0tzEHkBr+CcyFxEXb4UWXBdEByVzjF07uYdZvFPxpJJzZlolBhW6EcSgGtm7QySNiT6iR
i60KbbR2vfjXyx+QtvEr+k4oOYgVt1gXZK7cQEtVrgj8CP8dS9a5ixJdiIX40Kpfa0VDwcQsQEN3
J/7WXGLmupBcoprqxXETFVgpg2P6CYkrOAiWna8lc+EM2cvhWBhZX+BQn3pGQRQXcqez1y938pEy
FjrWAY6xtqjOEtOUkW+Ht/yr+gmN6SOB2Tpw9ZimXsmc6Idp+FnIBWYCK9m43WFwEptlMKpE4j2x
fwxj3DdzkMl2oMyJ/+QiMiZC//lajYgwikD9RZHEWzIJVRG1KRxiSfaKP6uvEOdMeV3roYQi+a7y
3mI/RU1Kkw2F10HLfkCK0YzVBUXqMxAPW/hNyEvg6AoLGKTpjLrR6EQDx2jVkvr5334oz4R5pjbz
jAJbGbIqjnUNv5w27JR+DJTiR0W1AsPrTSo0VRllJbqFnIddv+SIVhOrcB2iNlxH41grAksYrdvx
FKqbMQ+WhswnshGa98to+0Scyl239CewzMqxALKE3M0hbwcPTU47pPQZTABYrkR2ySNO79DhBv3M
fzCEw2XCcpGVJv1/lVTtADYd0vJlkdzWZcuzbCcOYEg0Prij9M/ZGAC9tSxyP5w5kxpGg0x066g1
K7nOwrh4UVvGSlGxC93uIxDTmaivPDB1SF8+8K4bBEzaSU97WBN/gbPnRFHlP/ejZJ3dDd0fooey
L/MNLwc1JTDT3i2o9jB6Wuh+9O+oAAfk3mE06TcW62YqVQTUy8tn/+oKNFM5enEzKSq5qMLQS1tI
jEhH4ZKolHXjiLO9IJ3Zwx3VHrv8CChHU4Wpw+6Lwlxz62gaJndoCl4Yr67Es9wKhLOvp2aWkCZP
oshNxoLTas9fvG34J0X38ffxeMMFzb5FtL3P5swfMPY41RtJVz4XyAaVf60e0u1zvnsvGE6w4EEw
tcpMZmkvNqyoTpDRXHUNZuMgGsn7uaWQb+fG+qlmajnb8m+6amQG12L5OWgxgZoOG73q1w+SDQZg
ZDHDqpOdmvB1SAN5MA1622g3anpUkeD3XuGz/rMlKsEuAzAiwn4L6kWJc/oZ0Ug1qod0OAGuDXZ+
XM/u+WeS9VIpHDJvzwHYAQakMdQ8miSQodiOa9fXa3Hc+0jfHXsDvXEYxj0dZyu8jmOcfOC5UHsY
/v816aEGzIDOaPJMVbCNxT2D6gZfZ/OblNahPesB6E5EPByFIwrsE+xoCcVFabLCLngLspP7T/FF
1i0ceaX0Jwks0iyXfyaCUiOJVdF3LK6QD0Eax0k5OLWOYkfn1h7a+Uob0cl8/VeC3J411mDbfU/S
FJSKEjTy4ynvPKSpsju/sEnFQKLZN0odJZDMNZRE82Kquw3FqYYZhzGR/qw+0/pQQFMVnmmvC0B8
C4NNmgo0ru2WhAnRAbAEJGntfpck6Q9abKTnJBQ5+0utsmDOh+h34GaMy0DdnJO17JaIip83DRT2
0pm96uTxZfMNgx1S3Wr7M8WRu2q+4DkwOmVCP4dVmetBkgdaBLH20xQ4B/ro5A0nrctNad9+zuU2
AIvQBwQXJaJGGQ4ZmBgFTVPkYETXOZE7eJYYhr755N30O9ABDVj4U4lnuQW7eezsXxEk4Rm7TQ4n
DpBKYWmDyZNPPsbiK5lVrNpTtfDPnU2K17vmKslmR3jMl5aJzEJNybSjLQQj3zy4Yla7wXObb9XC
pYUov52sh+FYBOyx59sTRAHY0Y2BwZ661NipUtes8i+yFr0mQLfjDWpnjJwiDDqO/bnwi3QPGQTS
LkxEFXUyR9ltyA/yUXOXY0+hrP7pTWMs7pTKDEe5eU/aHe1Is1+JzPesvZikVaNMa+WwowWCOYra
uAP4Y5EoB+EpUd7wjxe3vTHR3be1LaLIDOXxwCSrcqmF+NRBhi3EFXild83iOpNrV9PUs8+DWMEC
2e8Vcrdab/oQDGQfolBZsNZpEk1cEpBUS345nG36eqtgcirBcMMGc3+spluygk7ywOpFVgmhbrii
eKvEx2g8o2TuJY+wUHYBIlMaFGKYZptI2W4TLx4EpV9XFxSy4wXht67csKpmMItwsQbHZNt5vqox
hMWGWm8VZhwZi0gcmwFQNLMyBZC9v/4HcPmaDGchT6CCEbuPGVrTuE5hK0tW85yt6EEO1j3BQomr
y1M09otWf0v5M7mMdGN5FQm6tFLAS/CXcXSlZ4b45tEIp0ybFeOrayQ15oNJUs9mFAmcwGVrX+PQ
AzeqD0/oocZS4OBaeKhThqbGqVO5NhRnhQAlOnR302//TwgOgjDYXTtc6jZZXD5N/xJEwG9tnb+S
gkL+Q78kwkYlspImBek54//HuyV/CHohie301Rt8pG8AZZf5qw4bQVTGnWUQXU6pxcA+6doJTo9G
GwOmBiK8EJaKL0WbBUdYje3pPYXD164B776MA/YW4d6Q/2L13g4PKvzmesT9OQ2byfWPpxO6R2z/
3+U93mZNPn+qLI1bIJ7mPB6/jH7HzDh3uKozvTGR68a4UXNDSk0g9F4P3o/iZjdBFYXgBOeMUfnH
vCj58HHYsm164djBTQLMrjnXinitj3HIg5QWEnY1amHw/rjpYYtuoy6Mi+NBTGLQ1B0/VLGdjWXs
lnTBMuoDhtLzO/7IuCCCwlX/G+fwA35RBgcC6PZkvEg4FFRHZX98FcWcmzvLBG5ZRbt8ebtFQ6Qh
COZ0RKfkkd7Hed/RqkJ440FdLuceJdHKVI8oJUhg2LxPHDABik9OVdK8neb4vMK/3Qy5ityZS7e+
Ezv4aeZ5FY1myR6hityWcUYhRTst3pxkynCC7aqGuJxmrw/lRFdlZ81mNzYsHE3SEOwlteCBfJV+
9UIwSWloOeBB0uQOFqK09Ww99jaMcKuM6pbU/i7PbRKre1IR7vZ0muA2Zj8ddV9jSLQg9KR8M9fU
yrJm+CcsVsdsoi/8C2/s2wtB0GrS/WbJI6xQhoHMgLSYgu+1aBsFeD4Cuqjz8FcYS6v+LqwnhqMd
hjMaadQk0OPJYoRt0eJzp7g2YlSHVHgWpjuDvy4Y9sxLr6NtN0/IZduH501Ve4ET+LgwcyE+zGTx
cCjS64ljhHAI9ZO4StJsyzVQVx3U8hcED49El05sUxYL5RLpMJEJJBHrq9jXW7myM7nBJu3yvRsT
0Se3FcHoFLyGPD5PT1xqfgI9+CIsJteYblXSZUAiO+/ie7En2FcE9YCcttS6Kr6I8CXfS15Ch1eJ
jOZXUSGMuO/Jd0V8IsBKfBdMxqRYyOEz9VAkgTCVQBsXpzpqZjf9QONr3VYjMb83kSZIOebdzr8r
C5J3H3DikGTjQ/6TlqLgLjD0FDskCxqpN87hJwLPMpplyT/FmlyqiL1yGrk1yvsoNTXnmOT84tFD
EAiQKCCP5PwOflm7au+Q4I1cfYIdUOaecuB0Zg5DDgK9DR8EJ5J16J9IgKY2SR0FHYbdMbxaNfxT
OoYuDy0cGFrRplMH6q7mfaG8/xsWiuYmkvHFiTC46G/Dk6u8dcWt6ooFOqNBBsdVAG3xckQoARdv
b59+NUQVGMTe5/qvP0pW+e1byGqqXU6WagQE3xLHl2k7A97rwzkJa2AReA82taJDZpHFQKUpI7En
WYSFF20hNF5E4lCWQfHRv2bdAIQcULljVZ3vGtzMJQforaqL+drjoICmwfs3xiNb0KfM9YiqnfNO
XqOpBysKN5axi8z9nTyCUpCTCn9V06XcTttC0W4vrZuvuq2cEXWOGXUM2GVbDIfD+v91tRP2TOt/
TCEOWs0PG9quRE8iH5PXVlJdZtQQf6vu7JjtRhcsJ4qFl/iTzeQqKZH4vdLsvAkcg7WBUiBDXmiJ
T0lnzHDMAu83yXiJ/lqj8nkJOxNIau9GZJSAi1ESirdVZF3PRoBvGFvNPL8+32UofvxzjWHJph1n
d9GguD16H0ASiz0Yb1ndBy+YWFIXlIaZzvStEGYYvuw8WD9v0zxZnCFT8SaDwpJuZDLNmJ9/Aaj+
LOoj8kI2BOAft80BWc4a4/RBtnejbKvRD7IvCLiMBZl0K/BadKQxYL2+tzPgYSU03ds9t54ALmQD
bt6OT5EQSPX5H/yfriNro+78QD/JUz5+iHtL9SlmYKNa5iEEGrt2LfgYJfz5r2/kSRBBgk5qF//q
wHUDnEsbR3bGFoD57bXiF+KkLQwt7Cg4ZLYbtmkR+QNezYDadxy4CR1P0AXaJkUndgCXU2w10xde
7ZQ8pPrFCwJKSxLits+zOm3Vi1OBUULRO7pAa4gjPOKaujSIM3pmDyoIpXJZtwJYqzkNvsUO1bBV
OPZ5bV1PhPrRyN3YCN9hDra+B4tmxHl0lnj1aWPfJ8FKfBnNX1zC/uGvaaIHGriS3Z2QRYnyvpi/
WqifNjSk4tfZmQuqW/DSeFOvThSZmH2n1hVf5AIOiVRU057A77eEzQ1Ucf4gAoQqK4NroJBQ/ph5
yw494UeOD+QQWI4QSekfkN/aUAJJ93Nl3HYpHU+WjI03MCVYab4SPIe/b2obRoeQCsWs+331zPer
05XtNldHa4WfbJsaQ0sqkm/XxPY4+cUwXeK7MdvsnDSJzPAB+Izzq1V7+tSqugm+YexfZXk/zPMv
g8sREbkOMakGEZMWID5Ig+kib6krqgOO6tImClfqb7GLVDfFFCIOyCIDX9qR2Jlq7qOXgIx198q1
kqBo0Lfr/v720pqBXS424J8ESZfDo2Y7tJdh1Q6yBVaAaAUOnC166lyK1uLEVRyJ9KqWl1LSK97L
Uq7GSXdBaCpQtuFw0rXDDZzhreVEyb3ygjWNPIIYnzfJ4o+ZjvZKjU/tkWqyg4CNg3gTjs2Ss6Mq
idqK089cGNL8JEmmFBCWrtOsH/CmrVNpV6O9OUFuVhaNYgBkoo7uyFBtV2G+8E4r/2kOnby1/vm4
KzORWklfb21Sbw6Is9AldshTod1y2TBOpnTYFeh5dtgktJFOWf2bIB0fm6krRpD5+U2o8/8Oa6na
lEtHmiXlvcKx1PvIKzDa06VK3cyqbYZSbyozDaTuc5bAL5MKTVVe73g/fvJxAjG/PJ+DCxyLnTc2
6HwAMtUU/Z9Vp+F8qvGXV7J4e1GtnIPmGpHumNV+3MPSWo9d4qqqKENlOMzbCG9Wv9szJzqRHRLP
HOQx8jlNYqJb6+J5Ko7V/TaDw/1WEKpNJhhzMQ8DPThCL3U/rIbFX+wk8KgDTDWZfBQMf3NMRiw0
l/RHuOuZgD6tiswIvsubxTQpTpsrTotyLI+lYBuKTsnKydq1qEkaFqjpo+ScPWEjDgHWKabElXwI
uAWC459qC8EirfEUYLqWJ9kTAc9P17XVYFYjeyk1zz4sF14CQWeoUCtsyKIoIy9humP7EsJvLSFq
SheaXZXA+R5Gh0UpAOWQoof/LPOFyzJtjvD/E6AegMT1CKuUFiQ8T1RWxkTRCe9St881QwG9PJRa
DuxKbE6QmLGEPGowSEV1iz/YToYEtv3/RpplEmM1qkdUFqRPo6Eb7LTTWSRmI8lMYjBqFOE1iNvc
CDswkUb7g67JDJNLBe1892xK4gitdFMtBDhmf4bT87v1ZgjyAIvEKgd2aSP7dlH/VofKu8FYIZ5l
ge1Ueig6oAECbcb5zyC9eUJa0aEUdEyebpClJ6s9R5oLRkYwP5lcb+93Mlj3uAULvkue8Tw9pIqv
F2bhy4pMWq3nlOtoT6adbdsi+2ZUHVH1QtXL2hSMx5KTwvPzLxROGnpix5UziTuWAFdQcvhQar/c
WhT6SMG1CZzHYEpIAQAGTFR9weGlzCJNgYMweVxf527Gz5qOkJF3krSuCFOGjQBR/fR9b/vErVhy
j+QrBbp3YvtoLlZtOYIs/ESx4wzXcRDNMEG14aTdvh6NhiqDXBc7nL6r4FT4Das0MDYOGLE4MofO
7Lx6b7f2JCI+QU9Uo3pUJkQvoy3NZDAdUnHbgCYwUCDuZhQ52uS6ZB1U5BGcWarlO7+gqlaitMv/
qSjpDBO/H3BJ6ZMVTToIq+FnO0cz1bKlwxKeD0IOcgk2AFY93wHELcbbQPqaKCs9SUlmuxnfLfKq
q4APIZInnduJ5JWVX+cWK67BOVxfBuNNw2OKH0MAz0aig0S5JxwXe6HQmHZ5KEsLiP0cH5DSn699
wk1AwVj6IvmFjLN2MFu1aGYVH+mpTklKIRNnXeq3p/XNY0Pg0UOr0Qy1/pi/ZWbgCfYY7Y3zlXGK
MrbDXSW4ecaq/2yQpMzhY6uYYMBSGPRSEuzGZXirCeAFFFJ/ydsEy87a+S14Npc7Js+JNsA8cJfj
ZBIj8xvWG/rcLX//huVxtJ5+2YMS4LLFqR8qxYG73iyx5rxQUdgAWGY7K+rq8MpNquMOgxKwF8xO
MYfQ0VXuKQZCBnaT1u5bMisU0qMdCzrenqKWntPx5oveAwWabmVr+EFUTXkNsLuCO3QFnBZUq+Dy
PbJ3JqpAIjuB4CiPNTl3tm6yPW8FmyAoc7b73WQAO7KclWnczcI16bxoQ6ScfjaJwtP7sJOWylFo
QMGu3VwwhQCY0+lG79D1kAUWQpxOV6RfztlX6cDBUSZaV2G0IjKXAmpNUDJHYZRf7Xy9hjVIGt+7
VrLFl7FEPWaMEHS1nuzKmGSqjc/jFvXmKbhMHJXKYPI5bHnPUvmidcRgEGprb/7fMch6wFJ8V8le
RseC/gB78oOvVWgDMnzYF61UiXHgkA2lE6yliC2RGCROGvkzRCG5aqiRtg+2Q9j173ZHs0OFmObk
OkTiRfZo/JcRyose4Qm+UXd81pFAeoDF7gDlh/h0gcEdgx260dSS4sv3/t/UJjmFT6mh7aDE0tUo
vGfajejVSYdKdFkeqfQsmaWX9F+KW8hgYl4u3Fj849+yGAnMKgKT+qdwOQeIM+HHNGUItBbEG+pa
nbYWDW09VKOFbhTtAjHhRfwTMcgp9esrt6O5W2dTegsjOAA2361TmCYVCXeErVEP1w0k0SW3ld9Z
h0S/DQnpYxKQOTvzFxYouhz3/J0eftg5eeOVJk6hpdsHFqtDgZJw/k2YeDkoh+62EUMWD2lvUo/k
b9bQFEaB20bcjw/egAKDjW4k+T/gK3HwtJB4f8sUljMy2IfulFz7CtlSzTgdNuzJ8vHrSmt/tq18
lY1HVGXujFGe5PiktAler7PsT9j/9LwNuLKk8otUlKzryyxWDjAbjbU5PrEp4aYVCiDNViV9RZwj
++AhaFBVhHRl2H3/nmJYZKXyeiyMS4uQNmfWB1SyT0NCK4MSfqbjrtxHMb0vBxjvShQIKtJKbsTM
8vn4IdJkeBMTlUe3jRRpLrcgzJccabx//9DPfRRHV6F64iM4Y54csA5QNdWwGoGfZsz9b9PnRtTw
trBTze1FCEXBGy7wfnT7pogasY7XT2inX+MHM4GVVQTSgyBRKsnWu1Kn3hM+wSCf4agIKDBQfNip
zHmo/cLx/45DMeQh6rACDalQQ0PwHMCL2ofcB3K7cMTvY6g0ugriCjpxQFFeOjqZlqXSIFVuYRnZ
HqnpLdkfvm1dVdbJTKW7aCf/KQNDc7oyp63joH28vsK0l6Oogn5JONBXgxxcnMVelK7/SwVPukd0
ypgYaTj26NQFE3zA5JX5PN39L4RAN7Ngg9GWKcs+53tri/Fsdt/+d1FopNJSSvQmYSmY9gLo/lpc
zxtknMf0uhoSH5GzSpKYQrQ7gpm8xHqYQAT2EWXwqLnJWBGws9NC9HKJN/rQMdQJmt5a70utRNFv
a6HLkZGwxdKmHfzMJfnkvimlWTQQUA8MdSJ/JRBOB1rwdkLsIlCAEn6tx8BbsIZESvtwTuzSzHLn
V0L0CPLJgZ3Fq/QNm771mEoxnnNeMOSDlyAC+7P1e0hEyurRma95fPSHFkufFRNeHmPoNI8S3il8
xTf7UtYHuS44Q2oEzMn58HQD4U4YCc/e8GYM/Jcbu0+MckXnm7t6fRRFwj19sl5ifxXE5URQM5Lv
VvqbwV7VOdj5S1+kHVLQgUt32SVKMJvfBa44GnpwiwUi5Rocm0ACdNLpJjPjL+M1kLM+FCRqQN2V
bY7oB1ZrZ3T7BrIJGFVI2/dEFWNbg/+dkgySxacotfqqmP33+vA5Q4SWBe04nIjB2/Eo2B9QtPN4
PredCtiZCaod93W2YOTXc8nIuo0Y+46sFyNDBk277fesULzM6sruKZwrcZn2sGdOgz40aztyDEzz
sul2loc0/Q0Tc1oAe4CjULHZpJiPIoB1CqCZpKqwTJSW1OoqMpPpvzmbIPSLAH+LEahtRxOXzqBg
2gCYEODHz67SmatIj4isZWA6f64eNDhuzIWJ8YYtxBLnqQ3vHSu47GE0bR/bNKKrJBI86XoGO8wW
TF9qC9vuMyJfTEUNc5U3UolmDZbS9+KsUrLn6bA6v/ujVpR8dYzjZyVOkk4eP3j1J3WfKE9tf4XW
LZNVBobBGsdLb1YnYpaiw+uDDP5H6k7WqyWvG4tYFapHhq9ADw+BRKbb4T3mnHqNPMKnRQ8YRjk/
Doio7qMtjVsRV9zpqK0gUf6wbI8NU/Ah42wBJGNR6I/sFQpcsMInT5l08AZ/GXy8TI8CefOPf8uI
J1xiOhCF0pf8AnIaEISf3LqvDq7N1vR9CDrSRARfv8kdb8C+oPZ5uHg+IXmnl2K7WMECxEUdKOs+
3oT9BRMGKErslNdbKfwWQDClZbcFy8PWZQWqZILXPeU+gapjefPmvZruNFnEZP8ntQcEBbF3TnA8
b/7Gws2rkO9dv4DhTJ3pXM16vdyFG9jvetLeT1abOwdkg6J74p4NjPK6nAqfCAvwmMMAVsyMv5yB
KNKtkiiqqFLJR6ThxUXcKPeNTAdeaW+fu8I/BEXA92Em/YZjIaDLOfUqchSQz0nZDM/2Ol59bBQM
jqBgNOEPGJwW7bc8ZJNIiYiWaVkYQvADkhmMbgdYIOmaovVG4REHl5VyQQJSSB96bjzNETMX6kj6
5QU2d1tv3G/xO9k2rtEbFsdvvQabAaXvyyWiZezTa/xzvd3bhoKlJIAyNUggt9TdyEfhfH4RWI2B
uQKUI4n/KhkIgaF0emrbMT+TdutgrXl5TPMzWjgLT8ODmbj97VNRjQcSOip5XvZE/65UnHZ8tn5V
JN9yQ4wax7MrMoAFldf5/LEuLcV0eLcYye1ZYSEpgJuQHJyE68es1OtFBMu6t1K/xN6wc9zFv+Bm
7ESXwr9sMkTLIC3xBmwgKZO+DywDft+ri+XtlusRZMDB6DhsHGVarWf7Iqk3bQv2TtMuFbFnuMEd
wYkJ5emuVcABHt50xkPHooqyEe4FtLziPNmSaHHMYQvzvSSEKfQqBsDE3bm4TTKXMkGQqBemRmzq
goKC3zXpF/Mk4NduLFAgq9/nyuXm70dboyjbFOR9FWICt/sDkyeKbjy1b9ihmISVAnpnshYPsIoH
957+Za+2n9dcz8JetZ185l1HRxOeexuBajMgltVc77XZgVlwkVM+C0yh8o/+Pxt47LipFeFZmk9q
hiezjXtTOj2KSoLS8+ux8VYKV7B8ze3XOBroqzy5iPUl9U5yzjPB9eXb1fLdSInIDDLhnDMhaIwn
ho1VfPOmc1//c6ks1IsQteBVkXyDt4aLocxNiWmVtWH5GaZRsbBJVy2Q6zWiKJS1WNWPUSO8W7Ge
EeAzHOfdNH4dwYit5vm4vBx0e+rCyDz+IEXwcLCwn1Cb0NDU4TvhlZzTHYitkpiiaMizXKeL9Iam
U/THEJhUD7210gpwirZpCARX6qyLZ9X5McZzj0Huz/yFz4XrCOyV30uQkgGIoMUZxPi4waO9tdD8
AZWClsBoG5nYn8c39RvQdurVkVA1cSz2TKTjv3ay1gOzlKicum2Mc/n7F0jfYmJzZ6N7eM18D1vg
Mp/fTQ/WJ3hnem9Vu4sq5In/OT/kDgXib8YMOxFLaQMB4HPMtBjPRq2CrpVpwkxpAzL0aFoUW4kk
HlzfO4Y+1Tjnqoc/W36rzNMSLnMYvFXtV5spqKSmsRjOTAqkTGbjNiuHxC9vTd/1Rx9v/bSk+Vsw
YryEH4tHL1iWAwroSmpK66eyB3m2H6JzgeBRrwAlRQSGAMrHZmobI+RZPVf2lj0nWyAYHP+TVNEQ
szgU0bxhraMzz1NvvdEMg3zQXV6lvJznIhGSV4qsnz0iSHTSeCz+FjMrnOgIfjf3lU0uMQs01Fz9
YjIy62sRMnwI+eZhunHDQSY7P9Q+lbABYxVv1Nea25FtzvFZwONJv3sxI7kv0Q1LIKWBRQnwPapi
hybj+7aXI4MEtfrxs7X+pBD1D4FSZHdl5FzOy/ny5V+QF0X06diCL+XEksUKkCyBb7/XSFBu66ZB
1X/PsmF5lCmpIS/RwyOCKfepi5RESOQur38sHAVaYHPrGqfx+PR9C9p13ZuyApxPPC0DCjktZf3D
Lg05U+4VRXkiaB3DvUhAh/FwDx0cZY8UWy5sQJFhYSLIF0a0xv1w5Pxr7i8Dj2Om1rtoFZoK1aZG
+n1I4dfMwwfIE/FJy6IAjRUSJosg5vpA3skSZh4CEhal39A3JEbkosbAt5AZPnBq32EJHXQoIyKE
OwocEiH1xsd4NZ+DRxCOE3ojBFhOl8Dt2uZ2y/nh9s2tiROEY5XST79Z173kd98+opuWsgqOiyxd
OWNvkD9N3/WddDclOm7/ck4y9FDnfKn9KU7Z2T/lHj7K1zxDvLsx+6n1Auw98CqWe1yKYof+jUJm
meb4ANidzxtCiYKGH7jU8F4UKvBXjBsysiH+pUcrdVgVVdi0rs3tga83eWnfxjlwMLn6IvimD0bg
/Z2eDtMhuDPBzVBbJFrG5X4PqdnEies2TZMaw+p45prXORmfM3ils1AT9j45n8aQmfW2njMMWWOh
3mHVdi/aygqo+OjhCKdRB5VH0w1FujZsQmUs7svYg1MHmi1sFf52otRX3qhnaGMuGBoYIb5f1Kvu
F1A+ZvdRKyzJeaZXHPrWsaero4QiG8Dnnx9TuhLyVDIXqL5Y6TW6oagNuN2PfDMTEEWczcJ9gKoF
nfcK2EWPSp3z+vopensKQ3uKzLy5LPWsUNpo+qjKlgn9cPnuaFh5hECVWkoFaMygpRxuE4yaagMz
QbJleZy8T/L76w2VkcHJz6DBvRfuao3A6I6mUeMFz+tbRn4BhpgyLCD+DWqsr4nuuO7JIGyVRJDR
+mqk8AiT9Hz1Bjf8RnDWnm0eM2RT7bNLNStgMWx78kLNOci8rRyJhoIFWmF6cgn2kO1PALILZ/Ck
o+b1fvhgGnpKKBSgayX+Nu1XOhdolgiI6JNHUCRVODV4Kw+Y1NJ6zTiYjUL2xfY3oXYUBgVahsIV
E/QEKkjSCrfYDeaefeeTSTF58ptJN8Px7f5xwOhY7M8d9WhkihxNP9ynsTY5FQclRPuCHEt4rrpY
pYt5Jge73/INUOSisNWo+dUOpqTWIUEzaYWbXBSeRaA1Hb2VTgCR2pSFq5NPw0OkFQ1LyzjBM4Cf
ABPqn3CyQ+dYO1XPjjK9+gCMsPJ/7zHARudHcO3yu4iNkIy05c96kTgWa6IAd16nD9r7HCczx6bM
jNc1jlGU4nnj/Fb4aTFlEHmMlAaaQ/S7/SSJLOO2wil7s6szwRCLEGeKcCbfn25jBJ4B7EuofR5C
UNimI4cdlHgPxWsLvFQKyYIB/Whe1zLE4oiUUh9978iwmb5PFhawwWan1tfKB0UGeDjX4SEIxagJ
zc6uylMiaphDzrTyWxzXNC4vwHEJQJMyUt3Qu8NHFvT9G+Cy9bQ+R0qk85tFfHwlItDruaRDZaEr
kBIl/dLDOYD47GX3UjXgf1qj+UI2tl/v1vj3BALSHa6cu2bghqR6wE399Jipuc3VX9rHx3+p9Y14
smH4+/KePHgu1DgjomJoOb2Ot4tyWUewkIvuNpnK4MMiFxQ8ZUyRZ7hkH3tNY/o5FpaiMJMX9Efa
eb6bOakUDQZ5mUajsiH2ZrrO3zFfEoRurudFj6t4WebyLg35eiTkiYmyQrSaAVoN1trQE1ED/449
4twD0ZZYJrqbFa2IwTAO3RHyIteqxj2U2RnRHBduAzs+M2WdK74RXshNZ/eGVzfdJehCpo9LgLRv
G5bueDXxEqjvDRyZq9QBrr9wpEvtP0yNT+kehiSdYS2X1gQTgK3tb6icE+Vsck1znu6OWOjQ9D6t
lT3Gp56U/hifdruGWMp/NLpNmMCwtK6B8XT4XJ9bZFzkPpCLcpuHojONA/XhxHA9pqQBKgFDrdGw
L+hLsLNkilmBqW27TtuW+x2NRv78TMCqJrVm3eCWNhHMQRKDFXrEH/aFiG4D4VsTaQP8K5541cN2
CNqXOl5Nk5XY5bxSXqDA954TP42ZxewSJp/XQH/NX62/LI1dNxXwMiKXIUnOZRA/X5tEncvLFH4r
5RvwqizaPJlzsRnoNNdMWKYWrSW0rFHXTs7JPBGTSzEt7WXm3nIEPGeTuNmd/ya/t85CrJrf6Yn7
OhS3NdBjSIOo0fIwXIg42iZPR2LajPTooGQmvbuMhggSMyRXuu0bhzZ5jjEHATniOdJGzJDKB/z8
IJsiP4oBdH1Yd6RENdtof98/5WquzhDs5MS3v1kDlJCnmUfl7X2MXq/V+0LbpXUplooABYaQeERs
LQli5Eokd71OqH09k50AaPkfV4hEdbFS6tEDnSI4+Emhwu+87XiXYwAo1mnST5TzMi+zoDNHrjbK
0rICC4HXVFAiW9M2oIk9GXQihDBwAkB3T+GKg9xCelPefhmyzHrJxjJxutiw+i6dFaghD+6A4kaE
H7KsVavygNJirB8oMQZP26+m3+evOInvkXtqg3HPMCiDVpHki37pAStI7ihTJF4UkDWEdSlbEqea
Up0IzL116PNmd7oeGscwKwaYR2xxmrkc75AbyH0Oi8zXaDUIG/M3xhTQ34gZi5H+wdBN7ALr4F4y
zVXNZgz8iqd50+lCJnZCD5WUAwV5Dob1gLeKXwvMHPd8n2FGXMhVCyatDpFrj75XC50S1XLU0UEr
+YbRYwLTwEY6rHfM1mqsVinn6uuZ6aTZeA4vkmy80ecEoMtwHRVOKlEaVoQVyCnIALlpMjtNuVVi
6ooxbFhXqXnPna4rBumv3Du24IJxVVIJD2uozq7/fq8AnqqOuQW5OCLvwG4oTjuD6ukcMmx2CnPX
ISVDk/gjVASfXByT6dbrDgFPGKrx7EKB3/lfm5UM7rAgj8C3I4WcsHl0qmwW9yk5WgQMG2cm7xxp
XnIYfN5QzRHMMGnPw29pvo3Y4yVDhTdXwciK6ajjzj/cYloUhBke7JfhbkRRR+uYzBjdnAVSmnQQ
aJ/K88amWHixIYGS+reCXmxersGanRG99Dn4ic+NQfb0z9tRFvyMRPXfXgLEfw2z4RbHH2OtFqYD
aoVAT9Y7XC30E6rtrfKs8zDi0BqKSKqHMlvPP4lHLA6HCkd2lyj+Yi+XHHPElSNOB9pVYIrY+Fbf
wSsvZGXotBdFzvyg97I+KGvh4zRT/xEBIAHiXD2RdjJA1dLF9nfn6Anxa21h+6NWSNizM3PozMq8
DJ7z3Lu3NfR+/Ec6w38eo7FCUWDWQ+l2682XrufykndZCdmR9+KlTKq3PvSeYuGVszOjurGFOGFL
70IAdN2UdTfCVrtNQpkZ//RTzWtxvSCt0Hel2EFqnbPqe3ozy8tQgLeKtZjG6MzUmDWA7hPILNxX
HXPqmURElV0BWPlYUwIz4piOMo71WEHcisXJ8stRWuDNPnd9CqWUxA7kTJmv5vTb4uW15EACHU0I
iDgPXSCXyY6TBNFcWkLnO3d2Kb4xPn7GSIT2Jqyc2KXumBd0uxupqKr1Hp2iUn545LQWuR7raOxD
4nf364tXgGkOOBZUo5F/6L29g5pwSYbw+8w0+W+jjqW8neAVHs/yvXUIgjPJsFfhPz2d3nDsnP3T
SOpStyA5ivTHNqcUU8I/pRwdsQoY2vAkAt04hkqeYiblCgtSW6yoCOdJ9LHRUY0eODtOsWhrZy/8
qvnq3tmx14Qtq+DefODjiG2VkXJa/cQXr6bHJ2NUfnMjMFbq/Ds9eOfKhWzoJR9+2N/izQy2nn7+
IuKAKJZPxpmceoUqqUGm/cS7KG3pLzej4aenBGNihPmhlorqzmB9LlZL5NHjsoXtew/1WbpI7GNV
Sog67ZsUhyF2KNjgwdDjNzILaJMRYkpWojYVWY5fdQYi3KzmRGxAwbTXwIZJ87kr/amx9Foc1rKY
dWKkbMw59lfClwmQ3Yj0Jevqc1Pg+Pd5F3NKaJEHMt2bAIJpjnPOgtu8OvTV05YEgsjfF8+lOtNH
bYM5bOqmJVQW3XZW/6VqUlWBy+HmYUwtRLbZG2zwuSaM+A32rJ2JQKKaPDZvjWZE7uYXfJX4pSUn
ccQ6kQqBrWLez2p62NiNpOSj7EYyy4RmUn9dtSJQYKOz4fIhXAXj0lbCHGI0WxU2g95FTXlaTElt
GZpJzZK8ObtSsqDfJ3C7ev7z281sLuWi356OW++1s0gipqWkB5w72JZD6RNWn7uoWzt657W+UA2t
tFHmFcq7DG8vJghgpWMINA4MMZsEtWBIPsI1w2XRnsaksu4mp3dfRSEWPfM+duZNSp2myaUBCWLE
A8VLD1yLdx8P/ikiYl27bGBlf9wkVajkIw7V5CidKmdJHOI4WxKPjGC7FCFopDhKIFpEhK8pT4Qm
CxlZM6yIcG0VrqX0u/YqouNK8cP8d1nddLukt8vOyMNxe3T9S6YlS1E/DwSDc+TCzBqWdruCDWPW
BA6ISJ3I4fvxO042Qv48c/zJVlYtbh82SwHSy4PrYOSKpWtwBMsxn3bwL9L3FuLqDhiSMSFLeiZR
XnWHBx5Qg5PLN5xltxf1pwmmd332ul/MwGlt4FzXmA+emvIaVMlGHggO01WkpsbculdvYkSYAjnX
y2AZ29m1KS7SrdwMcCQ/TR9z3Meo5xkrCg0j+ZdsIkmwLVY6Gfsmx4e1n1zctPxhe3EZT642Imr4
9FsGlTjShdk+vS8TX3TY2Vce3j1U26Zyj/OKl6U2FPia+1+nwe9zZ51p5QbSKKDDSlTadc+hx12p
+IYDjEITpxLJGPy4snIAmLx0sPAMyHxkZvJnyysKvTQlHS0M64SzJ8BRNw5KoNZAbWMiVSKcHIoX
BdjDk57OSsBoa+AsXjZSNSLcbVnbm7H0atcPhV3UT1EXktfLz5TMLXjwFr6BTwfCaoqQeto5EVtr
OAjkF9qxEyAHzTQzPtWeVNr/a1A+cUFOgezKmQ7L5OtdmH+LfqI7dBb4TNpQ5EbzBzl/pO/Fo5UE
ieEGM4eiUqJtko/yJZ8KmB2f7mNnPODtrBV8LiJ8tSLzox2ZqxWaf4k2ifVcN0zCdMLM2cBXC3Z9
AkhivFtITcxmtQd/47lo7YF7lTUeUig4xlwSqzuhf+EgN4M5zRm9uNRqHUk+/8larvmhg2LqUbdj
XM+lbXsNEnbI12jzjhQhuUo7scIvkqJzDlO+7JZRt5pL64XPu5wkPrcU0HZUqoJPbI17mcsosRBe
NbvdMmMqJVj730jynItoJPI+Jz56cIDqy4fJtIQcMoZkmJfWBaMHxZ9vwh5uGTdFvQV5htlsoFKP
gnOAoXnWeiq9iUaodnRnKmFGzRlxpdAS3Ds9ncgQZOsNZXKUcbJCnBnYSBc0j3NyChskW6qTSHPu
xfUk4KUDYRCfSb3WjJFEIaZVhAFGhiKIczE+0tzwxYU4XmrC/+78cazopzsJmzFwnqFKwuuQcWJG
FSzZzFaL4raJ9ZYLZ2J5KBdM4m2yGA6iB5O4aQyFAQGygrolwj2vHret+zErECqlQNTKcMuDLYhr
IsB3/dkVcTbSGzFcNEoPos3Lvc3Z7mhQfxdt7+58MdGvHoCy0YxLZ/npdi5Nim2P8zJf3lLnBiXO
vR8TedjhRoV6JtN7zIy8rs4CHtzU6TC5WgpE4kKGTIr2zIh4hy8YrgMCUwiNo2fadqnTklQnyG+E
eGuaRWYC8F+TM2yGP0S3lFp2nKxPFfgOa54ZVV9Oek56lMITkNKBJRuDNG+k04V4noNHCwclXwcI
pccjKqLq2q/6lBG3GcYVT4TjgjWHBvaCI5of5U65dJ1dN2j9HWUEM1krNUYTqROZWypDI7dFGzZm
Le5Z5kQnCCZ5Chkjwhdw50q26D5ketLG+7zrFArNv40D+gUddF6wKaTPeBht6vkxEvmdG7SZS4Ay
HX25XLDnd/r4kg+N9/RmNZjfxy2bc+PxNi8DwROTsex+Xrwmx9R+wLZYJxgHFhN6OhBFk6D/G5/J
y8ZPFYh0gdpK++2bAodJraA3EXLcmU90pRw+W361VAQBPkdoPsWaQCm6m7ulkG5DPh+okTZ7f5ft
kN4K/AG8K79h9N1/ID+8vaXQ0MNBuzbI/2R1blj6cBgMXGOfriqsyHfnnIxV5ozhrZaxXDun1wUi
4o48vCzBSVveVLT1hWnRjqq/J7IgbR01vg9kWcv2F9c8L/psJ7fQadrBu6iWsdsmKTVXYLsk6+xA
pM39Nschw01ZoawEIFMjqps0AkJ7jjCSCbodt14Nx+YCGPw5Wm8AD58GcKFJ170ZZSXx6eEBYb2x
L2gXOEKULIEWN+H1jHfA/KbPWKcT4GAvERrezhntQ3yesLApytinOhZ09rejYvwzxz4HBl3BkBel
qnrv5X0fhWLBZJSHZv9Fl87dZ9tooWnFmUX7wuqgOtP9jV1DQ6CAgy8wClTv2kvNW6EaAfCv8sO3
ZIpqa6BINM8YL8TNahtSFRTD8SozGlRZc1HP8FKJRDskLTAU5a5HP9Ok+k35GiCk7imuMA4g3ouh
WCquwppfFthZ65nNhFW2WomdpUQQcVWLNb3gwLBc9h8MjHdmcEkEnmVF22e1yQP5BrkObnUkBWik
KUzAaNJtrr1C9YHLE8l/QjPXrkBRORRf88p+uHJk6vTseYwpsZ8dER5GZ1bpmNm07h8nfxT0An9L
c/49udcb2kt4jsMI/t4bCUx2XlkwrBy5+D/h43DqoIZqeKQ7Jf5g0YaKC4NCq+WnmBlPLYTBaH39
TNmoFGE0hOf2Ba1SngUy7YBWfPpaZG4u3DQAafZsV3fkzvfi0eX6cq77HwUxOCqolLTH6xP1lAt2
IIQRnCNJRWeYFYlyBr48Wj6svGdD5Sh5aFgYHOlvZ2zq6qJGynqO6PJKsN0oYRtj1M/HrxnFcYka
ZtIwiXbinXWZZHtS5Y6wyF5BsZ5J80e8gSF8hAFHag8uyRwWNaexbwOqmuO2wApcKdtsuI52kUUj
wL1njqGKjU7JEgylfgHNvvJLqBCxSFw8KJfWuTkaZnXh1g8WnpcdYZz7AKhUQWBX5iyEyXaJ36Cs
1gTt65cBpEyLfKaC8KkZcgPYycOP7bXlXoe03RXmSwfsMvQkYsqbJIU19TmfQr8e6XCoVGeZ2w6q
fkq0ki/qCqZyECWAvid5FgJssQvo/SE+Sm0L/Vs884zUmosBfDUs1coLkjUzyGEkG97WzvIqEnQm
vF9Lb3EwgreyQNT+upyb1oKftsEdfCkYG38u5yBwagwjTa1UMtE2T7JJg/pYEsUkwPoYixDR1IfW
8eiDThYhwp6kuxhz4AsRKsMzMkdyH0qjS49A8Fezbvpqk/gdsFYRqXordUEtrlK22+m6kGgbKLWb
NXhlkhrgJZdpgQw1wMWCu9Dw3Dmpet0lcouvdL/L9cWdpEXxujDnWbPMNsYZ71ULvbrp1P9rx5fN
fXmEl4rXjR0nb0kn3BIfNI9ut5bDz31EvguxEo5/P5KlarpKmTR1fUWfPh5PyoGOPz9rRsDBKTC8
TBGK//CrWcN8+LMKkrIPAZ3E6+376QbLLdyr0NSwu0LcuzzjcE+H5JDTZykFUzHUYEw0MbMgTDri
0CAXXeGbs7eRDoJnDO7vSOs+rfTQI3ZtpcmoiMvpY01Pa2N1qYuJjOXCyuMaGhcGBbtBKzQVLR5S
GNiREiHtY1rpu4n06bGv11zHtz+4jsl6VZoGo8Zjsu5FM1hgoQVnHqwnJ/VcVAfDMIONdinB2oXv
cT2SnN/B90AlT77q8a1TjueruRFgVeTJ8prUrABKvaq48WbdhD+spKUrzfmEWKpMFJz3J5dqj9Rg
zOeUdCnAqN7ShLcFeR8hXnGMp5FLk2zCyqhIFtQY8cBDiyRwkg+fNABRVDObTC9rkkxfCi1KJnC0
fNA89ReKhuFiFk6UinRdebFs16mJEz5E4OJ0y1vPw8LpPTAVc1K5zSwwzWv+r91RB827Ch3dOeUb
5uhcR9OB0CEVmbDOliiuE3Y1NvehiwG4UsTYHTLD035vq3yuohdHOj987p/cSIF+UFRqiyOi6byl
yKxbZTDQVui1RPF1ewptRcO8cjKLP49b2Egq23X7LU5HnYRIhLjWFx/De9+iwNKxR4S76GSwl8j7
CUi0SRCWYx5p95raMI36q6PBp+gVD3MomD8yTJPuNyu6Gi8Iea0A0TgAEbmoB84fYRBN4ygHllSr
/Z4lhxruspk5/YCmnzLAR7zs/hZmzOfmhmePthd/Ddehgykkg2rKEbWKM+VLT1ceMtQoPpP/U9+l
4LYEI19w759UvkHO/FvvKmPlPrS1rOA4J4hFbM6aMyrIT5/qYk1+SXgT2rGeIKKjm87DPPv6xZVF
DzOIoajaxFzxzqFs/9xtisWKud4+Q+i1+vBHaJ1KiEjsvRAikiYVyY5Qc3ZdpOaU17NM+SZweQsw
lFfWtIb2yO9qBOzmsdrNWI4rYz6DEfgQHPuWKpvzorxwCpCCNEIxkhQEg1GT7ZZZq6779Fn52jZg
RU+HwVIakXg4yJWV6kTuKeeVOGJysxluXQlgAZ78NicQ0fj5O/pFET1FFPaNvJOxVrgqrbXAnHdK
3UveUvdExQ4NXFgoE7BIAZKMSUqJpiRAeE27Xkao0aPkRbQGmEWaxobTh9WXH+Drf16hqOhOFdVL
JjqD+zVEmbcx8MjdPxYAEpMbJBnmM8oeJy5/BZ+mqzlwW3iBeEdiEW4ORCWgNshPx0wq3kUBjS+l
Z/mn1/AKb0zo2YpwxHQLb7RrE/U44Rjj9uwohZu0Cg7vm6yc6/soHwRJh52ebzV0KiFgGW+qPoyd
2ACJCey7y2NL4MLXxd0WjLX1t93xR+E8+kpcmJMfPP03EIoAhStLHFCrYsnY2F6YN6HGAb7kqLef
7jvuVNAx1acip+HAmDGpVtyjJnvLTkCshTtFAw7ebJV3asp6WQXFiHMBi4nZJqqrO7jHkLrYmzR1
xs+wfwsCKx8i2K9vzlpEjrzq9NFD+/ivne82T5OEgg6QEUmT6kwpKnl/sRFuQ4p+ft+bO4mYq/E+
wj8rtjOVPBlYk5JTSkukrJJJ1UUMkVvNlKaXnQ+SVLXDw4kJ9jHY5HnpNCLru3QAn+gIUY926pCB
x1auOF6MvgW5WtRFd7+I7dz/RubceYVOUylJNiNQgwdEvN1q1I8qcY15rK0dfKQ8yKIPd4LPEI9C
6A862fIVzMk+LNJvQtfAuG//8DbwIgnZNuz1/CBW9z1YjWzuLyK6Lru9RsKxbpwrnQl9eHhn6xwc
buurkGeFlVMNr8VqOjN9iqYwQB4mVUPzdshnpUp00X/ZrOOIJ2Uxg8KirsIbIjgkPjjuWJhfYeY5
G03NOVPS87y5vmjtEOxSTwretBhoFBg0bF4EDIhr9AEifn4TZVyiAh0v7hJfGhFN3shGYvHlYgnB
CUW6rMIkGiNstqHdfYDAzlfaG0dwTlV8QC3kivVbS0W8jEoaB2F4u0iu1c/t6YEF6F0f647yO1rL
HTpXeMmFQZMvE2kLCi/5IA+1RUBrmtrIyKEyNYaswZy/wCjmPs1RtJtU5mNfB1psgq1eWP/ObEWw
hHm/J9hSdxa6OAe9vVagogcmW9SDr8uhlfMJsN/+wg0G86zRfNgjFWbkNdikMijw2EpR91j+wOeH
BdnGYOVL9Ob7Vcq9eYvcUVVSm7dZVA3h0ilIhYQTDome1DDlA115Y1xTExl2MpMAyKN+EhO/0iTk
zxa9pYoPS7r0AbE5uH8veeSw0/XklMZ6k5NoReKeVBoFYNUhsDpxF5MeyoF6Z4oCbALSuqqbwoFA
hNYQhTpivqxL0KDj4FJCc8FP8JRSZaTyvgEVyn5hk5m9KSo68T9Kdfx/78O7hZg7LYerWsHy2tqU
tieqHEHpaAuVdlLhi8TXFCp+JG60XuJU+OhW1ItVW+FfCr2LG0fUNdc6CHjxeh9EHUSVUOaJsnoE
aFkVEaVRdNEKawkeXLfbyx6QHeY4ZC9p/PbgALmMntXa1sEpa4Got6Z9wA33j1e3HcC4fNeTZ8lu
mdxXIyO9MkaZVMUx+iaWRRM1p+7iuAPhgc6jmN/sMRO9Ew/zPj9LRXzPfIAxYMCuEwSq4Pv3DXi6
VSYCaBv50Q3OqHeI1RiGmFSzqooVrqpWL+hEj1Ay7AVUPxooYIfGCBvPHffJf2ESLTfRCFL6WH5t
G2qdVVSz5QWu52tpCRRMqzc7zIXsUMhAtYG+d4BThC9176bPOLCiLGBty0SLtIb+UFYWWfG15nyc
AqqE2v5Qe8nSCdHPOLLwjZFOdnOnSBtBldRfNYpEI4pfivRNDGNU0xMxssXyRaYcv7PxHd+pMzuo
LyYjG20Ek6HHB0TpEY+YPrIlcga0Ydyu2u6bB3CVbTEQMa558d6vS4QxCqJ+n1nSg8ocGCaTbYVN
5z4u5fCEJmagxOIQRQiupQbZ3aX819vyIzTzpDQ6cTVC3FyhiiXpRLfrtztqpcqcblcOsUhbzf9/
oZraPfwdOJSemxXjqjgkh9KP6VR8mISA1LIjU9WiRUR4YcaKJpM6ZQioEbeK9fWeHb6uxyTWPqtk
8k7JNHvQxWss94eQ40z5PQPCfi7fYuQTEhl8nKx8X/+dFDYRbcPONZUncokAjuN9v9Oh4djR4O6n
BIzy9+x6bPsXH9XoSDuo0jt0/Pc8tNRb5jRI/9m5lFn8gClW9qu7kTj+6ob2OFzCgHyh7i8xkshg
Woa1z2u6B0niA4wHOnKa+BUi/iWM9dO4N2RupYaFHOOL/vGWagZzOVd1hwK0/Ofcxmgb2TUTrhAT
+Lj8q6ORG91/9DktsXK2Z/7BdatKdLqOgEF1xn4V+0HpJ9jXS+TgYeaTCu+9KE0Z5mtsm2vuvpX+
Ulbuwf55DuelEojnIvjriI84MfmgGWQc4Y1Tq/iy5L1FAzk7ENtObntmifvEFnD9Dvor5na2JGap
PHCrdwnFw7Fvw/ypsaHfx4gyhahrEt0c5H2Ip1w1v4u/alXtWUvspH/jBBljACQBpLKhnU+g20jg
IXCKW6cdurG0ATsGozkGKb7Sn/VHpq/X2BrxGxG4/zFHkwYzdF8stlkjgCdmmU23owsTqtq8+OFK
CAKql//YEo6Evgb1uS44Ex/5zthzLcOfC2jC1mF4CvJ3eQrJdBqezC5AAjSHC5oeOdFU+KPgMRSr
JaBjodB47lX2KdUHc8Sm3OckO3+JQkACssLflpnFg1D48EfBLABSTpvtIOxBbF6Bt/ujW/G56ere
FgAmfFSYr5IE6YkMZ8tmlmfbnNHx2oAPlwch9CLpMF+A2vLjBeUtufxYKl2e1FKsEpurD+rFa4bo
RdMUJOcgg3Lhz8sT7YRhVqRqZXfOWwExEMhNV+uQ7RmuUhB/Vdr0802ox3SmzO5dZTrFTD0h9E1e
KzgBmbYng7hLp76AUN4Y85e8tzs0A5s93TMCZe2hAsd3Sf3xE/eeRvnKryI2wdV1NNcOMzjYF2A4
3oOuV7I0bfOzTTs1WnusbTQwKDPjwdEdYQ42pwBzvlseCKwdXMCe58K0B4+Q3Y6aowIKhJfEYUez
hcDZIXkd8h+5CT9RBG2uVzlxuNRgNpw6IBwzs0LQGA/eNQ7o/TQXRKTbHh/mS5d9FzmOTa8eThjh
5Ws78WoUjK5VFCVluUBONhtNdmAg9f7rMqeeL5gbxJjy7EVBYlVhf+BEd5NzZsNgy3iNqrQmHomp
bL7LTSfilPmNzSBq/PiKyXbxiJdw1JMBWRzHrOkD6id9HAvkY4OOUL9el7pKV6peQ6ELIC/yyeLl
jAD+rGLUQ+xWzLNDelBFwOtB0zRCTKCWt303vIEdiq+vp1VBQpFY3QzeIy1Dqzu8+YM30TL4DGCg
6SSu2xrwwNtj9C+mR0UySesjXn7W4MvBP9cVSuqDb2SlFO6LnRhN4ZHyhYcoBS+35gv7kpSC+1tq
yBCbDqnyMZ/FAvv28gYQv7IVLyw/q0x4dIROLh0Vu71/vUkN2uC8KNBkwBvimNPom+AExEfpAOSk
w4W4OhIhjIUswsPbihtwGNwd47e27tNZBvl56hhaV52MahCVtSXVFUfVspgfXGAaxmV7Zr4iYvnT
Si/eiNKk+lA0rTyX/ZQaVX3aBePtl5IzDNCVFY+XgReG5cfW9xf5T59p/1Zi7YwqI2IT5hRlS0JD
rQ989T4S5FaR07PpROcA38oKWdtQS9pZ8BBaPCRpRECFNwdF6zFLL2HCT3ebaG3rqdanlJB33ygP
zzNT2JnHe/wX9/cRvW+OZ6s9jXpPOhMYSrOT6PP0qVsL7UDJmpFAU+TMNb/QvxrniQferpGnw0o9
Q+b1yrcLrn+3U9MmCE2xoMavhNQBbr0d1xV+ohkgc49kKfL+MToi25cpUJ+Auze7Xx0C9FbvR+9G
hPu668QjawHFdiHzPR1fODamcvRKFWdhJL4nTXqFzU1mbvQqPpYIBMl840flLnGknnvsRNoc7X1T
WXQjB5fC9eq11JIrLh5wqejxwIx+hUX4ukoypKCcw1AgBMDmjMBZLY4yXPfQ7oycKxaUypXG2bSj
B3nb33mRd0SZ0rBFCqDbrzmgp6iFBm0SkADqUjXrf0e3EkZd+MRoKLX703eO0jr7xY+FnMTIRCtB
i0OV/4kkX1JStZfupdQ9uFlca6cfMfTZGLcXdbfizxSV2UOvOiAPyamIwTnSEgx4IxyXk4JxRM6i
ENTMphx9ovUKfTIeXss0rs7kl922AcmOc5ZyHMnHClShWw/nv+0Y6BAGq1UIpXQP0HllC5QTxT47
kmofCip7WALGPzpkylnUMpdkF0iqxvF16idKnlYDhKqNrdH1VnmeQYLq5t9MKG+LbFkPNY3kTud4
nEHBsqTqlC4tjBy8WnZabT+GWqMZ8dSnthP+uFqZPtMt29xrDMIEawFriNNJXtE2Tt6nthcBWp+i
/n9o5C2od0nY9AQZ95/nihvpEBI8iJBNH4a3Pn5yXqZ7DxAbUZYAO/Z0EmAQC6eCluBT2pCdBJKv
3jJViROArmTqKfvr7LBiKgyk7rs1r9nDLDRFxavdt16Jq2/Q7LYHl5HMC4CBj801hTRLBvcX9Bu3
eQE6sXnua/7DnKFbvyliRWaU7n6ypXg8GT6Er+H30wEOcBc4jcSJfxMlTvHpxtVmRHsHzOEEtfZo
t15gG61QDgG3FxHDI06d+DKMfSlCOawREd9dnmQ3wg/39U/CwOxP+O2GkSidgu/Du6/idjpFgvN4
4DdGgW9JX7Kyg1PnlQ8bUFBXZaeJ++Ow63lYwtlon4zt6TC/e4a3LoITddRCbD6GVPAYz6t5F+1s
J9wB8wtW02hu40RnzdUDPVrzP0oSbsfTnUNw+XL9cGUOZT1SQQJIy/zkac3a7B3E9Y03pkWWzbNG
YT3/DNEHDX9q02lbm25CAivWm5pHttgE4KoBf4GyYg3qyx+WDR5D1IPDqRGEo3fPT+TQVv/oIgrA
Eh4WjshXJ/5nNb0v24ixYyluHrcIFaUcbnULk4l+CutHA3XKb1udNMWtm9FbXbxMrBojVf7srMQ4
NYuJq4pgcKrSjsF3WjJP/4UoGptHvwAYDfChQ4+6dd57EqQpu2nTLzHWPK5ChQ9SXAeKCLSxB5RN
mjFoxE5MZjB42YVxcE82MA8g9FzlE39QxCoQnFLU5QXpQ7u59cAjvYo/rVsm4Wzx+OHE4uFFgzY0
tZamzwwwG9CA0sl44iGpppOLZO8eudwsidEya+x4jq7Mko3n4WVVG2yuWNKCnytv9gcvWdnPhJqp
m8AkXVPmOEBQhkCW8yHl1fEmRtHRRTg6+ZlEIZRe2MkdAeE31P65lD0Huil4XNokqK1r0nmzYJT3
HfPxBcduXZNyukNi/A9EBV9T6NrP/W0TRKjYyjqbV6zHzdbgBGOBkDhs5F28HIJfWkFWwcAlDEcz
YNrHezPuEAnaz+3QgsgPw3s2E6N489wjs3J6TYLQIFLfpGsEm5cEVEOmowJJxs223yE+IobiKhD2
32cHHgWw2TM+iEA7Yz1BwmBcyLS0oBJZ+H9scwHoTkRrB3+2ySA606EGcD8floRJmsagQaB99V5v
+g+Xp2nxWnf+n8XviFNgpQPsFQxWOoQ5RZ9QWOrfuM/IaR8ThPRr2EnV5e6YOqQK7H79X7bZXAfC
nq7vzSSX5AlSvYI2Y5kyuycbbHQFzu+cPTyykgpF127dS+FRjcqd13KN1sU9n/uxTzhncrcItP1R
h4cvXWHbzNXHOBT/ip0VwL6ZyAoZbhKfHukGnQ7xqsE1KC/Q6bKG1iDbCnHLvTfIIbmkhamHbNTP
I3+1MLtVR+/HSI0G/1c9TLhqDK8I6x/hYDT15k4lawKTHgwcaBzGrdgaB4utsbAK60yHiXk9UPG7
HZeO+FKrvBSYM3ZiJ8bXD90BuqPygQ89Qr6r43Z8HT59X7Cu80ahMV22E9eBgcyBDlbZh9MT7r7z
byTFslI3wrRbS3OPzrdKH3lzUV7yl5/qpmRDhNtMP+QDmRUm3r3QB4qlaPRm7ZlLRV2BbvLxgtj6
LNcKzc9R1+Yc+YHmX2kvc43xgFaVEmsFVYCsOA6ij+rlQggPcYFTpWLI9wh4PBQL5gmVRfBLcHrT
Zzs7xtFeTEjv88gThO9csxo8x6SVyVP/GNX66PWB7SyOQIBGJ7ZMkWG9b4MKjr0gwtXjmg/c6ssM
ar6O2K+kAS+EaQd2kfdMg8C2vVVOTglkC18n7fjZqxM1xqNIYkQsNzF/tAK2e/pNxZWKNI1DcZtC
FGccDJDowVfB0YX9eAKdMUTww2T+SRQvhbKEk45Rmx0i0Q1TuCWSUv+iRjEoh2qX9KVeFp+bepHZ
nF/l7hhnmFOamS6zQQpZi8rmX+owLZtfonBDfbB45N/ptubZZ0HMiCa2X8cnjGNicrsHrvb3FK5A
3+C7a0nku68ZrlyCj7ZXwCIlpLZyRsgLynrP7Siyz2bO7YHan5DtLrNXWa/a9V1qoKeGwKnYGEBf
opNMih39QafJJDiC35vcpCrz3UPkXs5izmZ2WpwYNnh23Fw5BJuNoe2dQPmL2B9Q9sRl5zgesPbs
8Wb8DXJo3Hdd1sTY+6Ph0VnBEteglJmmJ65SAm50jrxcOoQwHoytCAdJNN6wK1Zayvxwz14OIGTu
O/ZBVEZ3cM10mGHYyZ3iRFUV3xdDmCYEOj0G8cdq9SHbauiNlaOGLFJ2KcZ6D8eFYrAN40Qk3K4M
MtLwpOpQJCE1od2tYy9agxL66wBw0D5BbUhbneP9XUMpeit54ssMa+ZCARBkXCvtpm19MeZxr6Ay
6RYaWal57x/YOO+Fbtt1GJcuZvSWm4z48ATvJQX8z31YJDzBXZ5ApFqDgss0MMYOcTjv2SV1nC3l
TnxX1udlUOjxL/u1Fe+dzUHcePzxUzEE+7QnyGoFzSR8flENrRIhQvI2O3OBf77Kj3cMFyYWXrF3
BQfveLE1JTk+6MlSr6RJa59R7v+zIJUiiKRd20meZiLLTeizRZcNUcwMZ1FKgOoyGJC1a+iGkyYy
eU8yKBUzpgRr4pF9cNUrrStGGzWJj3sM6PXKJOqZIpWl0adTJbHJ+hohWVAsMt6ncqMY0dEFrc6u
qmwWQcDLFRyyuA4AG+4B0BY9PRVUBeWa9MTHSE72DRXUBF+qTB2NE7cYLln+vw8SxFDuZeQ2OrjN
B/1SUuRPJDfFLzN6CwcCiYt1oH1Hk9eniMW86Mjw69zhFlH+O2D0hJ9js0I9gWXUm+gIb9ZyRlsc
F9zNmsp766AJxiG9Zatevj6Bj8CdPQxquiZyZWM1lC6zVlcgc1q4nmssGt3XwJTrBNyn0D4D8rdz
CHcCYdT9MZLT4fopqay2IYNZnrFCpfQ/hCNJL/XgN94zDgrCHweb0NVwyaD1hBi6D6xGXwTCE/jm
NtEsVNXnRtaVkyyErI4csdbRyAbffvL6Mvf7Pdb4wn/+QO0oFVAN29ZwuIseBP8K8iZTMJpC9cZf
BMzTED4EDi2PXRjDBAmbsQRgvmRPVOaI73b9vADntkPHqq6AhuZJ/KtZoUzHgKDBQrpkvx72vpjA
vJqY8X37o0Gus0gAIObw3+BIQ+yVSNmXxpxLEBMpZsvuHhZNIrS02AM6p3Tu/UgJAH7ehpFoPr6x
dCYbLCiVELGKd9oz+7KgqnDcs0xDUaxXV+Gviu96z1Eq6MkFjA5EQd8G+1IjKURXpGIoRZVLyE6U
yBsxCfidqfPiw5MA4sLxXkarGUTuOkrlWSJ3vJikKQk85fxSSqsOnajBbE6rYZUaBEh8t4YiA5yc
5gRxOBRTywwm9Ajw/ii3UdrIFzQtOcYVELWT3Ke9ymKmYIiD5oDwFsyi4fk+0zRVXgrvyk3zm4FW
xGbNZLvSxYqzlcaRETNLjB1uOzd9e00nrUJQPGaw5lyHG0GkOjgQuK/e/8B3I0l9CZogghRMk2q3
11+lrHyhADYbfT7B7dVG/u2zXFnVbCr4mUkkCpPkdkm5XFc+MXh7zttdrjO+t3pgKVsEYlRmoCEb
Zx3582Gdlv/xPuuVj2cA/+u1Xnx5ISWkA6NuY/3f50mfQMJePQe0x2Az0kmulFXqnMTgwi+JcjhO
FBDuaZeS4zaw+AnLKMZzc1xrsrDmoV5FDIcgkF9gh+eqFhPN7B16ciHqCoXydl9xA14q4hboad89
nqgqd2y1noAUTgs+1OPOYeLD9B0XgLCqB9LvYdrzDhWczKFovraDMCbK//miBh2lKIxGm+MieKME
sjdUtBdPdQOeoiWyZFtbWPvDIG7QFWpxw89R104oqEIczQOAVgCSlB0zR6f2+kZ//SVz1sA4QcX8
iIQEEQLDFVr+MelaWtYfYWU54xZqO0kkl9d1we1HAtsyyuVtrraBMcqqt5NQO9gMbnRn81KEqbRc
uYh+WFy2fZE5TNnOHCVGcis45kxYRhVpq5eRcxw2PkzpevZbrUo5/A6MV8X7VuGQqRzcfc+Bwn7e
5i1Z9IwYa3RQGS/fOI0qIZyOeBngCD2ij+Mq9y5Ib3iniRiUtz58DW+Tckr461LRpG2porea/65K
a3q9LLCsuV/umW/wyuAuu+3QhvOTSVQaSoLmffPB+/gMPTbOFdOlGK5dLWKHsSQObzKILRkvhrIg
ia1mg665vX+q5IkiUbOx5ef2/ZIq9nozpejYf1/qmt6d9/kWycVUM4m2qbqXeiRj4HGzXGkikjgT
vQY3oLmqCwbuJcG8mysG1qFepykO6C7o33SAwg/d9J78UW/c2w2e5+VE1zaS43KYAovWokm7wPqj
e0UFm1mtcuxMZ0Qt91jo/qDQXPqJdBHB3D5J2dIUkUgKAyHYTsaGh8e/izdxF8eDKnIO/p87mnhL
XTjd2jQ0A1WCgA2ZVmS+FZ6dMXharUun5CGi1ZcFemhHfmIrTfRcrev+ctmeJhCnJC9kZTf3sTs/
3/1u1GwofEknddjUgdOJTxaaKgwdGHOj0k7OsQLOTDeORhy4+W49QAs2MbZ/glyUym6YxHVIKZKr
7YRQii5WGWIOEw6kc2n2I2C7Jf4/Ick6usQaqHTFI7cD/1XfFGxAk0dNvACHIdQ1PUf30axdZSL4
2+Tn/ts+JecS7s9mv4jx8ZVThZ0NeNVXzimPXPboIqcU3WdNdQZbEsmDofqcAsi21J84brC8Rik7
7ZKV6vdhvgByII9WbBjAmGG/ShKwnnfBQyRS+pLAuEVi8ngy3HhWpcaEGTekOrSY26Umwe/90eP5
p8W6GiqLE2PCSls/zeIFIbvIVtuH9aDZKNgJbzGsdZHbg2a0j06XfyjgFnOv0iyGjcbQ94N08NXr
OdHqBz/VNbh5oCsgNAWuGFwKj90VCMmT8ExULWAWlS1I9Dbg4X9fANAAlz1klmQxS/Sv8qAnlm7s
FiSNoyHQMF3vc0HC+j0s7emPkihBhgzLgghpe7i0zfSy63U9rz8Zm5DwD9Lt8yXqGlzM/a1ri8WL
siA0vafRBCfCwm8TtQlg8wSADpoK8KYdyLFY5gOtugJnX/juw77L1RYp40LYTLnjSOVzTAGzcot0
5j0JJsXPC4rKBP6kQqWpyPdssNZB2JzkImZg8qUNsStsv908hrFLzmH1fu819iwxWD4ohGpnfo22
x0Kw+83snqceo0IcpkZz/jAwx8h0Bqs1t/pCNFAO1rPDlk/Q8j1KkJeGbIXXWIDJBoejLiTLdSCm
MpHeDeIzvWcjLjOlzt062/853TStpADcxcLCDEWe0OLRlU6wtwePA7CS5cC0Wo8ChMmEaEKzdE1t
36d6ri8gxCkfrEwjZxVN1APudF3Db3HxAlQkvs6XWMGZ/j6cv4OlsWovgZKqtEIEIq7izkur6pEf
9SBkHXIECbYpfCgsrfoizAkL4+T2rL0xOWcPy/J2FULaJiT7DrpqcMueqO6Dk7p0StcrkaT97RRc
0ccabKW+l62am3TJVBsEKYI6YRelA+/DRQDyE6tgS9ZYjM3mrCzUrkbwNroVfGZfWREVTuGTe+l+
UeSvo4l9GKtKO57LQjLglsW5giBaiZbx7BEzaB4EbOI/UAHScm3ADCK8KvqVQT2xQtZjxqr4HHI+
SV4SfHxPJwWOkcDJeKlerDIzKxyOcHBt92eZE38UFG17k2guKn5E1wp5M2BNsvVvge9yXfHzv5KY
Tu4Wx6UJLR6XhyZEJ2oiDw5mLmF3A/oSRlUG6DPJBNHUkVptkLykTWJn5VGILGIiB3sytl/87xqR
tCF5MvWbIbXTFrgPYC1a6UlWAIaxCgSPRCVdwhBrCJt9P8tPC41LxUM5FVS8z5RS5u7xlrAn99EU
th2ZrqdKFhO01xU9Cnf6uFPVxuqVId6p7xH/bS7yoxCfiWO9bSRSehk6qyGy+9uQlBvV6riRiv0S
QgEVrRR4u6LajDZ4eswYv3LAlW8+QqMcMzj4gIH8AP0Q9JWocq23uRHcpnle+JTG3qPmKpx1d8L5
/Jx+x+G4ZRcWu7Twk6c/MZJv2JC0cQNfw/xLuN3OR7S4EbkmzussknibK+/X+lGANQfdeNTywLZF
HOOMxsY1ygUJCZzsm98IOuARmQ3mmbmNiikOrbU+dcu920xpYGZZJCtH5gEPHG9AIn8dXhAzHl/S
2F4t1zXvnLMgct1wQFewun0orEGY+ihvCApBs1uYfTt/snrKzO6mczIPS2Oup22tb9iaa3kjzQR5
R9JmBGAKgpC/YRYNsFvHAJn4JeWvoBVAP0cq3tdmF6pwSIzkvTUc2MRcTvX6N1EI5IaAjz3xjMP6
Nk97lLRY9E3fHNCoCFOhkb92meJKbXcG7unNNFPAFs0dQpamyXohHpo++al2NlDZY9BmyKxAKkVY
151P+epRwBAPfFqDBWJFw7FUo4TvPHerhEWIQl68d/damsQFJ9CS4fqvEL1IB9UCE6xm5p7a1M1v
hnZuuBh5D2AW3RBzBtgOfAah4Z8tGXgi4ig9eQtqHtuKZugz1MlN4eQa1DzeYIrSW0m+crXGVe7K
stbNYLrhyHrSzE07k+MDngc2f0ZwMe1XD1KW5u1XukNT6rwTKOCwgyZk96JDADPz41BJbpjIO8va
1+LXb4az30Ido4oeQNjnY7NR3TDq2ZY2HNwNeQ2lwmi3STtYhwNfdXrkcKjCyL3ECnPb7WC72wZl
2JFzRSduWIkSWRwWvOGRj/vHJIfke6ugnE+98h00uvWsz/rCGMAqTY+YKNRTaP3oi6WyzDxEhdab
3ASdOuAt/xgBfO+bjTcV5n5D9+NW62DWNEPIwLDCNx0i2D3un/UhSoJPhTOnWoykRnppZoXRJK8m
srmcSR4rgBYN3UcaN7nRw7scqxfzBORYgM0F56qba1ZB2ritbPyKwD3Ag8RYVBo0D9jfP6jsVoL3
Kg91pHl/zOajirSYsIPCsfLosVtltLelWnHQB7YjHoCtnFM1X77ULTgDZY29eE/nF/aKg678WI7r
f/M0C1H7GP/KxhJK56lTB8m7od1jly2skPeCAkbVNzJKZ0A7a89spBf5NfBwjsLplUUjuWG3Nofc
bgVvWBD+1QXpI0HWwnTmNBA0eLQPf2sUCFmxPJr1/7pwGu3fAT5iY9KEReLNqV/EBmisxgMfUmTS
mE8yzzaio8i6qus3HusEk8Qrzx0qruxy8b5xFCQYa9kTlmIOCG3VlX3eSXcHCDX6cQfgai6W8dNk
eJEQNSwxEtd+cRV+7xqH9yb6n7GygM/2e+j1eg9KeU3duDrhlO1q2rcEoZxcq/cDzQdsQt1XHou5
cqLmgmy1iRn4gLzfBgHXqv5N+Zk3teCIE+T6z4lpPlNYu7eMaua895av3Iyk2Lbk2AUjuMgFizFi
bZYuGOrRX1E3GQ3pzSKPjduLiZfSRklMZZg/x1aeu6H6ix5GhXzC7GBhjb+WZn2d4Ggjj5rI5X2v
lj0WzUmtmTjPXsLYZNqyQBLC6gtlFMGEBou55U5geUwU5XSHx/W48cEkOK1/FqWWgxDECfXgFf0y
diFWXXinE0O8YQzlI6pv1tV7PtHbCP8M1v3h4p2/9eIIi/r2OF7v8929t7lPqAsgEY95LY5KFs0e
FkesY5xy7XVjiBJn7nmhsRH73FtaJfSeEL+oEyxvYd4Jvy77WwoXZ6oIzgAr3i/RkkwW48kecDKk
zPPolS+HYh+Rz1zq3FG0JLcKLOCg+d79CDOEAr0OXEBCRF0s9gbuAoqU0h5bsbC8ZjUhrM0Nu5fC
EwtxfIFuZWuZPpMtXbG9YvMB4mdHaYkcnFE1P2tVD+3TYRlHKJs0RsyfbOc2UREg/slNXa/Gh8uT
LbCqua/bbThsgL3oSpKIuj6xKc/CgxlmzhDG7bHkYF75+M4VVF6r9euCRP8ztuFi9yD3Sd5zXSm9
41HfnzPTYWgbXhEVoAr5W2Qlv9ACFkLDI5wp9dDbFHsEw1zgtIGk6W/H+DQvQoKIG9h36CS4X92T
GjA3qrYGmpi9D6h49k5ASViR+V3S5DZAD+jTcNDmna68xekhNeevIqMoSjv6NnBBTrnQTXU0KPFL
B+v0YcC8byAQWiRGlpxnX9gwmMx9MdgUo7Efvgkass66lrbAQwqPgAeWRGok/4Ff4ekrJ7miVRCc
LoZqF1HoFlD4tc3fnIWkOnSf6OuMRf1pXstG3/+h+UOJXwRnxsmJRmXdrwTqAM+x+lXH+mMCYI4k
qRmNdEf2E9ZJ11kshMxMcdKs61YFZbmysdMZVA7nNI7h+g+/jaL1VMzzXC9q0NCN8xcnPHeZbn6D
v63Wq70zFyZxbYpvhEvLBXc7QBN12fHDJGmb4UhCj8+4ppGavMXcsvKHNOywD67IBGTu0mywyaNg
bqYuJyNzHDUi4pkbD5rDb7s8lgSKM83EYQaNzPiQIH3lNezivn1RGbK7Bbsi1VozcqeZC4kTKhGX
a8iqPIFLf3UcKAmSjgFYYZ48/jYbsOQc7HfzpYEBhE9LeNT5tQj+zSiITjSNnZCI1psr4hqbg7yG
HhXe0H28D4DfWovqTnUtsF9zBn0loHO7kvFrBt68LcoOrS1/lVGKmEaqhAHGCP/h9v5KfEVrkhI5
G6+K7zXEzBiTo2JjGkQPVtszp+f7pahyS0VrF0LA8IXmPpDY2Yx/qtnw4ZXADpXJhzYqYE4WqGPB
Rh9fseGS1cn7po/3L+IqlISqICVoHnRgAG0hMVy2ShjPmwOXbCJ9wnb14VYi2j5PPKny/kUgzD8k
X9WMi8Zl0jvZc3tAUx1Dwkd1TJsAGLBIC3r76EVd8ACjETMhpmi7m6M2scWNRxQRoknstSAP+oV9
h28OB1hzMUuzg7AvqQnCpIDEke6TUb3FfeOxbPO1AYO0pCRdWDD1JxDRf4wovTfqBPGcjeu1tGf0
xRdTa6DugdCQ81G7sbULZdAIpuEiNqk07fEdilfPkfdZJf4xXQUxnVXolTkPEHVS601e2ZK9VLQ+
Ya1KH5evZmxangdChfFSmx9vrPevhn7gyZAjsyj/2PsN1VN3EOruoWiBPIqVv9NDl252/Gejyiaa
XQsNm2JIv9/BFeNllLX85Z7GAF7NCnc2ZUxE/9ojW9HThpk9u6Wk85vjo+q/nT09J1lG/scTrNvj
Vm2yiXmMPg4/IwfkI+gbO/jum8aYIa29ciPQKWUB3zCx7r+K8fRAeNLKVUegSoLJauEovIQCXt7t
7EaqhhU4CgLwELusieKNKTU3cR7GFME93iiNObgNT3Wzi5CHv98s5ba5wOPG/iyrIsDKHeXTLStl
bmAjB8KiBMMFktG2fM0t4relnTZnZRiPyw7SJonNRco/VmmUlvauYN62tTS65cSi9cdDmqTmjt15
Ms0u9pZz3jcK+Su378yTARoitq+mCHM9vfLjhPZZKdHwILRT50Vd5gwuU2B3AYFm9LruCa7j3aGj
xnX/Bt60mCj58TO2MMJsF57+wPmaZ3RCXKSApXWel6bV3v1VGJitpgPgDZWNEmwB7uWt+gWNUKcj
HkEWZI+x2vkebRHIPYy/LWvYzKefr0kjOsk9yym4y2+KaqPDuxVFyQVjBipol6uGpvRijmVbEm/B
Vw42f1KrHBuf/d4PnJa2OfuWP499cfeoB8SPbz8G9U3FmSqIPgt0UqnT5dM1SQfhaIRK2n9tfiL/
N+RaGREAlU5qaTT/E2cT69Fq22kieNxXAp0ObB4rapArNBwbIuJP4gGWmrzU1R7anh4EWQHClFwH
ypa0cPA2tR/QbnLsmzx4bBGScra3G9nMusHWEZ9IsGX9I/SWAsKzHyUv0ju8LRqwwgTf/kWBlbB8
hft3OaILq85qij/vBR/Y0XHGieFWTuPdYzA1IpET8nunihk3IeaiSzlUIpD4SFfi11YebUH728dU
IQpP7JKU+XJ7r5dEcw0/G5HPikoTg7sV+FOh0k+WbJNoikG+VBxZQqfTpGC5vVWYEv0zXP19RF2E
4/jf3N6pWaYOKrUPDe4mEA4P4bhyF00jUDW4cyqz5ZQa4jO7PyXg3f6DalZu5+wbBBxbfLw5vv8M
VWtwB9WKk4uJLMWpXlgBhUYfTR6C32T6KGRL0N99SPt7oGqoBMTJjD37RkLz+IPjamhhG1/uqaA6
3WKwmPgVJcrgjj7A+an7bhtEeVPyOg8qoe+MOdEFTJPgA/HzhzKmco2YiSsB/mK3MGQz/dvH/Vst
UfJjqaPiOOsH5A8PaUuXd0gOYZMU9I5xy8YR66y71p1nd8JtsF+ETGylkgRaZ6Tl1p/lUgqc1Gy8
HGVLYH2SeHDsDanKp4GyxykHArtnEyRrDw5Y5WlZpGvVHulbfR4xeg5N5+HUevQKnF4t5+IPUdyf
LX0c1HG2zzXIFqNeunVuEuOKTxjVxoBpWVJgHVTMcfzGnQQqfEwyycsbzQOtTxPy+PfD69wzvyla
p4+w7vfG3HAMTFp2JDMqwHi+G6MCwyeCxkHuR04R1oEQJCfA5sVewhz0izpXD83E23bwtBg2MAvd
ufeLoOgb/G37ALdN6+9UybCqagzeOUU2mGuMOARTxUH2o7Jjug46ZkWFIDM4KE94apbOJfWE7uoR
jWxPvdOTzvcmDxoEi8f6I/n1+u5xasBIt3B9jzqvC0HVn9t3UOEtzKDa29+7azDsLzgBN0QNnMFI
CjQugTeapHW133C5q8fshNj5ulHAcfRBAYSzJpFkUA2P9an4tV0emMRX22JMfsmH7/sepi49QQfm
yGhWwA+UyfkjyKyRv+k8LQCJGiYabxaFtjim++MH7Bgb2+biLTUhC2QnQVE2tsEQ4L6l6l3tAqBv
G0h7FAjQ9hvZ2Yt/phu83oLIPe+FUxYHEN99oMjmC+TegDCMtwkJLjFw0SwtvHer/tyGsuAR0YI4
U1R8S7N7hAb14gIg0vqAgv0wRXu4OkJBL+f86TcjYqMduitF6Vgt2f1+f0dTvdT6qot80lQbQtjw
J2Bd5Okairs8pzWKZWMRQgwzV7JJRPIDh5mhPVwp08lpjxsxN0/mftS2D7dkbuO3h36t1jeHCRy/
I5XmgeRIETFxsDQ89MopOGLyqWs0zqygE9rjMnDF/67lopoy9KJP0gUL26NfLtI7lDmfEncDvuNQ
9mwMnfl7BjL1V4yskfvIx9uquQ2qs6hwWRdsM9q1gXzZyYT5pc8zhgxWdK6em3Ksn36yhfYPOk6c
zBucZOIoWIf8YQ+5lSFR7Gqvur6U5jjl8tnFA86zSPFhZKEJIXapSOQefPsxQcgLf0hRfATNIQnI
tVSjbSRelAXq5NFEPPR+OVpz8x2xvh90IQYgijuIVaJS2KxLZ2QzudClxycey75yUbPI5DpETHjt
9IGW/YuiWvl+aXIgQEUUjW11Zn4tn51JWtWUnAXLXla3pwqS+FhA0NqoudLL7KMRQrf/Pfj4AN3G
52WsAxUQ7HfxCzd/IJrhYP8aUCyNuTdAMMcyBVR3xHafYSNz9Js69K+APK6hPzlYtIUVv2iFl8jN
VZdZbSMYjKtpHZuCjYRhnLSfkL9dGXw6vpKxyjzR83MGD2FPEfRI/10Wg2nvkkh8P366u/NoyEe0
Gc5WxEx4YlM1EF2gmdW/3tfsP1yVZ+OWgbXqSGwKLQCrBrNnkJrqApJwoM+zaofxZBXSYmLyAYp1
Nzi0Q+KTwY6y1eWdu1kUVtf+N29qiw1vhS0/aa9VyDbpMDhXq4wkR/2gnI3hDJ+LSpL5Nq+6rkth
daAMad0wrYWk8g5Mv5X7gDeAANW/lloyKAgH/vGoCXz+umz31ilCC7imY3hh7m4DPh/H1uyN0GGg
INpzPw+eFDKQCOCgm8NpRJMzvVa+DTNAdTyFg8GA5dGry8G30nZQkD5ajRscdIW8NRLE5ZQ/xwS5
bHYytQCdTRXws1uX3bpYj4SKBCP8cq01cpS4ueojeAaMtJnxQwVP1nn9Kam0WTdw96p9D3YZ9bK0
ox4fsg9DooRWEVyvha5AtvCajVbBFSdkLVVQAaqsseazwNTCOslxLuKCwMsJWRQN9yPsnLjcStWP
4HQwDmI73Tne+s061QjQuto+X1LTQp2Leppde+ION2Zmr4RU47IFW95pZ2fW5Q5QSkH0hECujVhi
4oTU01fWI77Uyh/GfsYmKJtuzFy4aIMUvkPqiW413abCkarv1SvfLhZvom3WsVsdRkmdYEPTJCYM
lzxAx8JfSPzXruuT6AJ1ka0V9eIZ53PMkEDZDEkUqdo0aZ+mhTnui9zsgITmHQRVkCg0BOL7qwP0
p8d8HvIb8BOiLyFZQYW0KOxolvGYsm6szfJ7kSDBxeWuPOuxKODYkLMdfMexU1WJy/9CUgjzIe/U
YaD7Af61XBsxv8Fy9tcvHMwa+fABHr3eYNbXniuxStGKtJ1eQTFqq6xmcNGwMVAmu4MT7c1zfVUT
7v++yhh2Yh+3W1ylfLtvyT15EHPbef+UyIRCaZBJu0ZuUkvg2GhxiuckDqWIu5+MVZgLxPNs2lM1
egB74WCGw6gSGSiCY4ZQKtkwvSXwap7klP9t+dta6fxBgK70WHClxIyeHZWMwoZmA9lBQFf+9nvD
fqb+yVpS5IWe4Lon3KQeNxri5DZrUddmqG6gmniA4OHIclgvOgq+zN/6AC+/YjoZxffPiJVhxTil
aROlYKrw0cYZl6IbG7uRPs8wbE9l9eYbbt1Cl73owKh6tm8cmL0sfJ54jf//1SrqfsXb8mM/j1As
S7u45eEq3YNutevVAWyxhLQjYttHIVHgMXog7zVO/rBMPjOTCE7PZqmPv2eYulpDQwOOnxYsG/1J
9NUgkj53UvKyGZjMHla/FCr0O6diVRCqFMWw9WS+D6AMbmn+Kf3t9wNDl3JH9Esq0Z4hVnwfAji0
wsFwiuL7TYH5W6Z+965Nwgq5pEjSx9B8yFk8OnJRMJDqpWKgkNzuuL1qOkDTafH56PCRsk0jnoCn
cCSW5MvXlicuJFbBrd4MdnQZmbwN5IQ+VSsxIlJZE5lEdwNI4XzFtPMk5AfCy62VAQvp68ph87Bj
eN/F/oGxuiMjHZLYgXnEzoTuaijqHBZ5325OR4RaUAmQAOOao+qPJ0CSaK7XJY/WYtRJUeVAnrd2
zfPOqP5GdrRBsKw6roaVyrZxoW+8UEpID2VHvg+xe/OIQ0jDEIOhdn5IAsS75OoWvsbrUHFpduIu
7+zMrmn90GYZOe917yYLQiFCuqVxHPvRELXv1SrsAsONfayHuGMtoYufc4Ll5FoR3LDlbybxta4h
cMGcFF/8nuk7Q9ZGnSk8nukU5U+LDrrYwY2jBnNXhCn7+mEW+s8EJdnXDSmmr4/U5iZ9JPB3w37d
ELOpuuobRJ5stGAEknI+phLUigD9Whv6BNw8hT9Lzre8Tc2JXsVeUCtDdQeY8NXyRK9EPdn1it3c
AH4/veOZ3INm0SdZ5P9KV0U0iM2rRTulqIakzaYk5SiBvdmzmKOg+16Y7NNHv+g57zifEhlK1zq+
JIOJI70ipMwMR2rW0fEjLGF0H0B1+OXAGD5eOTYZ5CFf86sqbxMHlRjQj//d4+gtoBJsH2TmI1Vh
QkCmGpxcZ6Q+wm5bDw9Ac+53ya9ydbx4kqJDawHYnmC5pKyFHDlleNaZ5BbvKspajKu+Gv/0Gf2D
HZLFvPY/FjMy0fuHo1Y4T1jo5zZYOG59ew5TOqQBRnEKKeCzQxxoagNPw5FXXUh49Tp8QRg/izEh
BtiLbVQt4rZWdiLtfkCLf6U8PyoqTiV95eLCMn5R2StcK5lU/4+Q8obsdJpA2T5whAiOKs5TdlpE
/SZqdjBiYLrcM//oz++er8bH3LIUmxXSPeJWcxdQ6Mg3ZDMGqwGMh6F7h6M4rAhLvatpxvZ7xQmG
tt3sf9aiDyn70vIIQCwsb/TyYK/82pasUcu13JMKX3zxWW0fvCbHkV1tcPTCQ1xTx/PIXFdFinbP
NhasjJhNlCBqOyiOwcZlY2RfZOq9u602udNO9ZIAYnJ0qSbkh7GJPKA+UNj48xA6Yhd511HuKg7+
U/kgQk3HC1E0SXT6hb7i89f/LOsI4/074ZcIVf8ovg3AEOOnylTVNDDyQHCpByuTGvP3f8n/l/L/
hcg8jg7ZiPvsKY9xC9ZsDw/5w7DfEd5Aw/yW+6gr3UYGZzOsJMknPaHgIEcmO7lXVPD66Q5zGlqo
LywYtjEPG7wae9ricp63kxk2lBiMMaS/bC9Uf7hCdZFUmN6lFPfNaGmyN1i5+e9iGwDjXWphlaUD
fLbCCMd0Cr+q3msE+mwdU3JPG9LY+hyubHHSyC/bakLWEcS48XmRfIJjyw9rGQS2f62kgwjnuXHB
1pAeB0G3sP6mcrf2WcALu5VAG9SNOGCpRgIj+RIZ4Tk6rly+dypYgbdRHXe3lb9kWLz+w4QYj5+E
L8jQf7WMZn/V5v1NwHSsGw+uDQ9p5VCw3StVk8Kizm4ZsT81F4RT+WPlpSHA3rBArND4cbkj2HOR
JApmlswzOWdi7PUjfgenTx299jsIdT/L+zgzLXC9fyIzWA/YyBJ5kzKF/UrNAEoVO37Qsaa9EDQQ
x9Nfxqod1iN9H4aVBEFiQ+vJmU+kLHp3QWCgUXgQRFAteu/iJ1AoV2fLN8uxN97mUa2BY97kRuKa
GSPg821tsCNQy9izafXBIgZnfhT22Tu1r8/hcx5qxN4/aZ+gSmjFYhqugDkwf8w7aYFxPAMg9SZu
nfjv+l3oRPrjP2cNxIOdeyySV0R133luW/0MuuLdgSzQp4RGxdKJyWB+4e0BdnBbxfwElAYqxgbX
KYuej0WfbrSmP0knabwky+6Ws8OAmF7hql0TeE8MnPSWJ25q86OgE2iL5o5BBXTtEgYdFODVfuLO
HzO6Jg6I9rV1Kh43LM9u28bNStj6VDfp4cVtBFQdvLlOGqxexaODslcfH3T9yp2CSaJREGW9U+RM
HypktDQ2qMFqCkeK1DM2QPq6GqsRzgIQiqbubDhUs+o1fVJ82jpaagC7VSzQTe8Oe+rl75Nzlt3k
ZqAtCtdr29b0YOhk3tssU/siA9iDFpyB32ItL4gmM9XqK+305aInXIWN5NKQlITK/3aEXo6Z5kMw
C15TiCKehvW/1VGz4Ug9K0pvdvPdjo3WiTL7eMb24DYcELSoO9Pvtg0Yk8prFTpf+P4AFLc+3D4t
UJErfVpXd03AWb7WXpXmpXw6qjfugS57MwLKvLofG7fP4xgRYev5IHq7Y6sKRSOTso362r4swjyA
sTvS7lRxIRe61AoCCZ0INfQSjsCd/aZ9d5+BwhelqlgkTtTaMbszqgIst9lwz+idnRYDcnd8ZgxS
dKJevyT8eOpLFSRFQEUJWMh2pEGgAXzsxVpJE/GWQ1DQtE7ERqgDPOYT7THD6PTwT6SIpZVr7GaW
gZVXHKdShTWlYcDOcElHOAS4Kxio9gSflA8R+5LhmsGNyH8D0tbniFYjVF3kcPDC6IttNiPyNEM3
FufyvXsnp0X9qUbLYqgp1mpv2RJ+R0seAyJTAF0YkGaSsezUbiFcuLhvflDSY5hqyzKzKNMR7Tow
A1X++x7IX53dBJdbSOgk9gCxboVajjcd6ZnYVY/qBvK3pCcwjVjHKktXQo7vv6O6GtRz+gnuPZVo
dzb9R021duD0BznLBr9ZSbxKbkFfRKGwOetzpWD/cL0qn3ICSAJkpQTplVX/7q/GFqw55RawWwXT
jNYVgyqENwY2AUqCJJFNsShTUQObACY9kKLlmUBIYfxnyAMLA6JePSV61AOfsGrPCl2L5+HSZuCV
KJRAX9vm84evQZFlz0z71z48hvtCe4wczlQcbOSC6pyNMdmbZpiviRGmOS44uRY0TU3T/duW0+Pb
7Fby+7PrFuECS8XX00Zhu13uD4rR+SLC3swYT9SBewRCqVXOIl5sB2Qkb1Scx29/DQN+vT8FlL2m
IK+nJvDMjJOGPhA38JqBUGcykm0YbMeHdeiU82X7isXTgXswmyHf3YSwAHRWvoQgJxEawAD/tuCJ
9iL5ECnL3HVr9OJ/spOlpVJvdIxcYBnrISd4npMtj040QDMI+c8T3JODdRB8484D26NbbhKC5KOw
nSs3Ew88ttydPp/qMILQA65VFQcumkHRc+eQpPgi3PKIdEDh3rrOSCxsxpFfvQX/vAUAJfM3nesc
tQydIGghEC8U1M++/pdVHxPOWot7ShP4M8jHmEphjzCKQr8reEJGVBBO4QL3y/b//eayqyvcOn07
eRMqnHtEhdNtyvubgoSqdIZyR/cV2mHQTZehsowwPf4xTgN+nvkroHjG1Zw31ZjBX8pFooVxi2fI
s8JZ7AMOxyNxZIBRhQ1hlSKSS4ExnjewnV2kYTfRcR0m+dPnq0VxjJP4fZGwNVUcUPDPfeoRf2K5
aSehEUU2H0y02hYbMb2z9pVuUrERoHhN6Po/0no6VMENzwk6V7xqKSpiSF5z5sCaps+hohWAgnfd
vYA6ISY6v1Ocjgk3v5vi/lAANKbGqaeFht6+48H9cNaBdTFrpnnrTufzh/Ym8t8tlrQ/3kZvjeL1
5ZItVnNfR/QD/4B7rzyl1l4BQP/bY2/7vse7IRmE76caTekp6ZWa/rKtsBKx6FyTfBDo3vASLX0L
rLIKigog0/tu+KFAYw0TysdlDEAi+FmyN6Hh86USozgv2ej0shUBx8M3ViywINqnkc/86neJVYSo
4V4jgOfuWSRdeF6FFkKoctyFzej64u0hSnjp2KEQ0VnU0zFE4J7b+v1EkHy4H/Ws7ZBOMfgCTBdd
2mQCGoLDp+cJ1IyWQOCuntG40MqEh/8WAHlyJbAqR3phwbJu1Vx4gn7EPEOmcNCaScmydMHR+P4B
90fxvgZAXkcKizxQKcmM6f40pplphUPbQlXLqyxGFQnsbcvFnPxCHn51xbN0OPz3Yg4nSs4qGpfV
agIDKQWVYP4yIJm0Mak0alO+Sg1FefHHO3yB5O1yFzqQBrx+bQcATh3NJGgUOwN6Rv91sQBA2K55
n8JJbXvcXkYLiIByyYtOC/UZ9H2AopyDST/xtTMJ2RM9IrqKKKS1PTaGlru3sy1zuhp35i2qZc/Z
HlFWe40Rs1B2tDc5/NLDuBP9MG81DlPXn5UFufZe9dM4+c0XQiWVxy0quOnXFYnxfQ79N2PhtJCt
XulT3w73TVWRYvGp5uZT/U/M52mlOlZ0AMr/VS13ddfXyrsAVoBOtDdJH4Ap/EsxkI4Zcy8JJDe3
ZDycxXT++G5T3M49E0zb04MEddVOLaHZzw19F+WWq4w+iSkedewjrP37xEuJPNSoTdKFic7vHB3k
ccvwp9XaSqfM6XwVNAz0pFpPjGUZ/o+A3+S6tuoN5twUBD/EzLdpZiFhLveaM7VU/ec7811KggqL
pN/K1mInS1TrzdPTraXHnEZN7NilC0BQn1Ru7Xa7FwYqcXgYDBwfpoXkixKgFjxSLcxU2ydZz5PT
U+dRI5Ek/k9cBHAD0z+tVlQW/coCDm6jouehAW78LktTVSn9hqx8V2uIxPH9V3dxosT7e/KBlNQj
JNp8mcELaR1uaVyGshOsv0fgFXvrxOjo+nSw50o05m9rDgmG6JFXdHn235eia76MUpQAIS/lV1AX
rnWWl9ZOffpDcoWFURHvxi3Hlq89LlgD/kgfQjapAmzm/tj6Roz6iWDlm+cmdPOCoGFa6pNwyvG8
adAElwWEAHOlo9jIph/eZQ1FT82LvztrxNWszLl0HiTi9tfasAXKeEm75lNCK4YMNRmFk1jvThyM
lhRa/ss7j3deZNqjP8bMf3YR4pYwaHCewFhcuJGsaScc5mKgz1Ade6lLKlKFazTt3Jpr8nF7nPDB
BqD5t9frv1D5YKqo6hGKkZMD8p8l8Okp8LnhuabcSQDdZp2/veWFLHuIavxmm41OY4Qr17mNfmsX
WuaqeWLWqyzG3/kODCo/qq9xY5dTEBFNNmqCO0zaEkZOjLVR6nXJzWrl9eE2WE3ZJpTRTJ86RzRb
xLOCouSXHznI69WJN0+GLfsYaSrb/I/ZzXmyDbo8d9kPdDagRochtJwfhl60GQ6/aG7OtvhBLg+U
CDogTiPR1/gIuM1Q68ZqPiwUf8l/MBzp6xOqCqwu8bQcBuUIYc5sKoa8iohwaqx4eJ5i/+Pu9Scl
6E2VYyE3j2IjHDyQYDtANLgqLh3/SYwEqpzfCY+dryZZiZEZzESRk8Y1okVtGzSljQstrgmfmXXf
rMnm5t/4GuYbntnaXSpPUdKMKbCklqMnMMqLbtzG+6mmdGi44QWOTXOlRVr31PIqqwnjuDKC9+vq
v0C7HYNa6lT4UHNe5p9gpvLJLkpp+RF7E5HtG03jJrvENmXysMW3ZTptGVjX7v0MYVH9VWofSn8I
i/ZBSWVoAFo94uk1cDlvBhrrRdAckU+lMa4KQF9dKo8WQE6CZXKjHl49Wpkn2Ywta+7DuUFLb88r
Hy9cHv6O8ClFevsBY9UF6C8oZmLQu1sfsyU9oPu8OaEcVyA5S0cTcGUwMMq2AfMFzLcGKhWjTHEU
4WktWxQKGS6eMgQQJvj1sHYJavSCghvI3USQqMGIPeaJeb4qROFjltzIcIxf8kErviEZ27iCzN82
hnTZZALHAFBWScsWY98VgfMBDBFmvacCxOR0X6EBggMAlyV0PLFvrMaLKaQXsC6EkWzX+JGGGVpS
+soVk7z+cg7pBfqDP/Hd04t8Nben686Jc5fL78sJzDzv6z11lVGncy42koIoF26gcWjk8FFKHpvS
MJgJ7ug2UNH9+SQs3TIx93k6k6ZcilrsnsuAZettq4La2cPTb6OefDVhqUoRp/gUCuK7+z8zDB2B
X5jxOmetVqSh6HNDP+rRWW56/lkfYUJGNgTXkiacdaoEPwwKnsgQOGc/ttitHwh5Nz/OjK91i6J6
gKGaAfgejImkhAH6cs80MxDydlH0ZCDhSBLRXAVcUNS2aYJJD+wolz/dXngvQn9qvOI7O0kpZSzX
zJHU8h0o8v/Q5x6BZxIGM/GQc4FU8/dms1CI0phfcKWTefzLqxqDc+6IDkgQ6w8u+SJzVcLW22jE
gi108sN/13OeIO8E+GsuRNISN2IjDskmDVswuFgG4dGtSNi0pr5pKG5F92xPnAHYwmO/80uiUNgR
u3v/kjKfyoIhWlgVpGd/5WgAx9vc5OgnCMEwkhsl0668uYhJ+CmjLyPWesOtmgne929NB0/OLbHS
Mv3jLIFkICzCZya1ii6Mpffeyipru8AOedvA9JxkAs2PbPDrATyCYQM4mSEmVhfaqd7GGL9L4bYx
l9ZkEBK+dJ+MTtNrGd4NmInjCbJgoIWGP5z38CtG7vSCDnCw5LwSOx/QkkP1zWdv9tpIH/pRg5qo
S3TuDQ+M2H58Il12XYkBIxUFm0uqi0HmVLWJ7P9FEpUB3Lc+MExOAMkICxgjpk3314y+s0vYjjXD
XEz8QpRq9G9cPPpDOG/GzBOix34BbG+W1xhfKiwrdC86yNJqNAIHanjayd68sbxeXwlNfewGPHuf
hBORldN1K1ItU4TFVi0YEMrEZkyR/tEy3KkfpzurC1ztbqPXATskW950HEgIApPHOObp25PLW84L
i9B+oG1iitC29Bz6eAp7PbcT4c7aPRM+SJ8gatOHQeynK92hivqH7tS4Nk/xpTEAqPAPmGwHrO38
CebXfSpkkTKBCnl6jCv78zGu5z/In7rLRrczQuwrLOl13OjCmvoPK4ZUUBrmWUs2vBPOF20Cx2vp
eL05Nm5Z120vO0NJylU3ZCGiIfe96xr3WTuoG5mMopH5Tn1+73+d/1Npm7GvCu5Ty9yziGOG+4YF
fzACgWx++JW/XxAF86C9K261QSQ/IXdh+iZHvmwn30jsc1QTi5UaecKA9Z1AN3OZJVqNLP7CKYc+
f2FRUDxT3QKnABhzkSOARixn6QJM0kRCzYEijw8DduH5gB8kGarcDSqmOGYtQdiMjhX8DzYev+A5
lURuqOFACSra38nww9y2TzFl2ggxth60Yw/bbc4InuqJ0KoU6Ud85IqNuJulJlS9iTHxJAga9H1U
HZLza5d/w2uFvZCISVeVHsDW6XMDyYw3VGMGNdnwd5P5kHZ8GroIOjLKfoN0B6GJk8/HtgxjmJfV
LX+emdis5MJkwNzhiAbXHRjx+c7bFRpsBNe9JSa24uWJ1bBqdH/rcUZmls+QRlz9fCa4H4/pA4c1
Tx+wEXRSjKK2XLzLPp+uhNeYIcd5Y57JKzjXWO0mb/sIMEoUq3JGPIbdukGfbt6FKUWuELvvUJfd
u7XwJkvPEKyP5P3zYXtXYe1zZBnGAkpjhHI0r8yLxxfvFs//QD+uUXwjTMdONn+7PARnihmWdBF/
aSk2GDDzNeLycbUZc+ilfaH+Ll48pUhIsQeFN6Q9euHMGLhHB8P/02A93NVDwGwCAQmTEUs12JNA
VK9SfoPfnyZV/vPGV8ZVc4kGc+MHLOYrkHVWiMKCnT4Mk2ySeZf6bW8CSaHy4wqIgXIIlNtfaHd6
FFFjWNBW/CudjJpaYJIzPpMyPrsz5Q5bR4QiCJbAAwawTMls8hu5qJCRET9/lKjEQDPclWQRhDWG
zk1fUZNCjmOFuckWKZE9xbPbpUnOsbuUIqdsru9Sgdxy4Rrl8RdS6WSX64xcn5YwG2BBIh5Ocdal
uhSvcoug5VvnR4aGTP1prdwX43GnIXRXJzsn377L3CBuLOGsYt6bKaCwICpLWeqMfvHJ7o8BUVn/
YBKLGygwVMVc/QTMX4MzwN8fqya8dE4cqh0N/VXcIuUnVmr/IqfFI8abjGLvDr9BTt3jR6wMIdTT
PW8X7Gie9QpVhGK6BDX+H9aXHdy0eZSFcaMxpKf7EHm7jPZsMhMuNLIoGpbAljWfnVQMpHPwXPhD
S3McbXwOaQ3G8S0vz4H1GX8TUNW5+70tTON2+hUQB+SvpreCYqizy0pnxZOcPj0ZXym9im7pHyS/
/OSi1J37wZY6dGZRDcE4VQ2wH2zVQ1y9d/YbZZLXzliTWaW9aF4rAy48/X2UlCoVJ7W7iN3q0dWI
w3IoQ11qvOKLZAVnGEnZo/zRH+aVotLGMNTt2j6Wxiz4/n65v8WqVYNVHrm0jF7zLP8Tmq9llTGl
BOAiy+Fjf9Npup8jgRlbWTJhWpBbVI4iOA/ussPOhND0Hvqz8WCvrUOGGU1hQVywXBktKUtMsjKK
l90hbGUosKnv3/6OIIkcXhZNdpZtP8zPIcGXGTWvEHBioWaWIKTMHRF1Ln0yJbD+rYa+jJ9Zcc0c
/BfitueZtfAms9Y/3kfRixTHPByTTzxrgCJq4NmqUfQQixhtZlQgVbjByh1MiCE2lklr/A1uA2WU
VoTgjQ5r5x2v5FAw9cd2gh/BBVVc5KC2pCedyi7YP7JAKv9clzjqsMhdcK1UDBdb1AbJvepPdqJR
T3EvyDhNDjjpEvBANribQNUte2eDLyk+Pf39d3TU8zo+rCK61rO+yDeNaKrOXgtV4S6ZbWuwyX2N
bybVqGjJdtr0FzUbyk46qqEueJXVSuFadQPJWNmpbMfFWHO1Pr2C4k+1JI+LTRgN46E3AZpJXtvk
1otncb08il3em7weezgVQnaSDOJJBf5Jy8OKiWzTBN2R1BuTchekXMHc095bSOdi2WvxEC8hFjU3
imr2PkJmqmKVC2bbWR0kqlhkD5bNnQ0AYlxnsJi6ZfWIKnY+4oAuw4nv2wjB9zHGoMXxB2dOQ1M3
tPfz82g088n/VTotR6JR2lqA6gephAqFJ7RdSQ3Z+5Tq4x1SpgAKCGdSVI55PZndFc5qKV5aAPqn
P52IkgBkmnW/kAvACJ6np7qX60n+VQluTftUVR5IH75ZlpBz1dK5DoOxz6mNYnfaZznQwi0xEtnR
P6wTKr9Dxfdpb8xqHbFBvCrt17x4O3+1XiDzuMt04dLUOEe4Gdbl4wHcF/S2L1d4KezdRhFe7agH
wdemtBG/w7F15JjJgCadSMz/mdtoNUtBxYDFWvsAs2rEpRStSGcqbRP5m1F/o1OlNyD+vaqODRvv
0rQf7ymj16hUAIa5gOCmk83oRimw1koY8gpoEBRA11r2wb/e33VrT4KtwfFTBELVOuoCI5f5k4gi
MYPLd9tmb9+iC4tOeHtzX5RscLMyfIFLar/PJyBT8mPTHBi/tjctibea7o4+gll5zThnj9yTVJIJ
skIG9pdniE6wwJ0ESCIdjpcnsHhBRXS4729LTr0PRRXRKTsEm6ec0QXbPi+9171wpQqVkKwFyAiS
RAQYVHQsItFXjGj5Q3Tfd0x9uRotEFm7A4XPqh0sogXEdpSsrFsoDalBuX9mVWf1Nd8+X6OmREeq
Vz1t6bnfwpsK0tv4TBaLPv40xitcBnHK7/nrJc17tShYyxAMvQ4n6FjHXwRh5wwlkkDsuG7QK+82
L5gQWzF3YotOQtVfxK3nlIRMvzjxJ2cEWtR6lcH5AjsduyegEum6+Gj/iLfnuCQbSaS0IKIQrC08
QtKVyayqFhaw0IGKhaTBAL1O+MHytQ2ocROFAInEFuC2ebms1ltm6Es94SmAFTi523frfkru82Pm
ItdhOipUZmzM5p6YCiiyv5l6/EN0vm3ycwSfrrGZbOiKyLh4MI159/ibpOStbfBmHp8ojJdvBawx
3KoVmNN0CL8up2URra+fniYzbVGHqTa7vGVM2IsYwdPJpbqIzhaKsWn8EkYsXTAfVLe6SLjVdJtR
RfL9TL7z5FUXzvgi0K+a8nEYzrwHZZwPoht3xKgVK4NjwXduUJffI0IC1y7THc0FS8Z88T+3fgqY
0ihPDSMTf5pBcVMxAtq9p6QOC8IHIeRz777KCX+bu65wf2MIjwGCvmwpfAzWVaF9X/Q6OozJ9/kf
uOC6G5+zKrSRmAtIZfZ7ZrBsQnfzlw6ivdIrkRobS0w1jKzutEBUvmOzjYwgy2gzoRv2AmwK00CX
ulK7/LqEHz7xMUd8Jma706j0kMljhgHCOr+f8g5qTfuEDD5AdG4eRDXq/s9XpvWYbFnmpH6j8fcx
g09YlPDIT0gX2CjVwUke5ZmOxg/UYcPiRMXvoNtrQkzuBe1AlbWJS3lT+hyzo+yCCFtQcOjeki9L
xO0IWnA3m5SKsuOB9gsmQTNsiAvNermKzuPNXNtQWF1Wst4mmNFJykBT8r053qVRlSvjU1eNGSfH
CasM9azs/LjBsIo2iJD0HFGsVrlaieOMdwJfuhj+al9atnxEJ1EksGJoX+knerjf/92JPV+UFSHk
vSA1o1LQoLKusEY9EsyszJS+L5WyMi0Xi7jwt6KhFtlKKjLc5jgAwJmJM1r2P4EdsYpHhJIGfgnb
0cYi23qpRxCBjlrBNBZQQR59b8yTHt7Zk1yGPvTSO1tB/WaDNHWFajvM17MBwwZr1AvJZtJlRyeu
PHBhmtuuSDT0T84bMURUikWWcCYfFdpeci6hdLRi5SIGtzbo1cbNtVl14Hbn1+pj5Vc1X7u+XMfE
hM0CuGk8P7/dk3cihyTn9ZvtqcRy2Ql/q1zLuamFHGtFYVB3GWuw6CnC7NEmwiAYK5bJemLzPn+J
GQC70DtiSTuOvB1MmpMcPQWB5xc9okynfYr+k/Y5d774o9tcGHjWQbacSiC+aPMWGGDYS1QUW0uJ
tR33cIscrrdiVva3kFYfCuIR1aJLbnwX/qnEpUl13twbPBFI1a3vRBCrfDwWdoydpPBFEhThGX4/
6V9DtcZj4dmAKbG5jhr+DGB6LjSUp6To9MUp3C4sGdSD7NSK0LcdAl7w8uMCzYogCYoBEmgsCE3O
A55OT17gb3AMWQWbGTPbufIhGk2xFifR8Ykoa0jJgebffMlNRcvv/9VRPmMdgrHrwbKGfAsPr6eg
4KqW3y91qR0b6kwQPOuH+Q622pCJPO7+GGhYdLNEtCdY6glmjpC1fxKR761sAR1MVTmgAldgmOLi
+Qfhqp84G2aevLvOB6eqvWIKQ5siDAU8vXV0xbKvGu4nfC0sFip1CRkHWJwtKld4kDF5FsUWz+17
bFob6yOtnAEcIlp6cb1+7GeyCdYI86h9xyfxtMC1nWrLcilgdIOje6tNzmXh+9Tt8+EY8PpXiWpo
NrIlefJHK2RRdDG7tqjK45NPiWB3F+2mlsxI8L4y0cxGlQV4sN4JGkPHNiwAOXssVe1k1VbUxfy/
mBcQAoaeq52XHawz3lxvqo9Y9QEe1scsyhAJ59csX8UJlwn8jO4GUOyyyP/oqUGWvJt+O9qNOr6F
bOFs7j2GPX6ywHKNUSbNuuKHoUtlfidp3IBDxih07UsRLI2+KVsneOQkUf85tIiCib6jhE+OJGXz
VT1W+qRaOxybToIUosfhxlPDaK9JbQtqBk+M0NBKD4AGWemCLJEGRvN8zbHeBoqiJsFaNbJpSdsW
BSmvhvr8JX+U1Nt8P3W0JA14GiFbCgrdkjSf7ES4AYQFOcgCupZZMc45pW4FP8OneFXLbSI/GWrq
VrfP/4PmCV2spEGulQ9SXOawHaAvxY1xxRVCnlmZyC9OHgexsfuAOafBu4I8xGh1EhIgnWZrJIYh
R15HaHuKMqgh+q+bP4SuzRMCGqH6f2744CTwYfz7bQzYzigU1b9ORWCoPSLle0YNwkQ+IwrX3RXA
vhHIAprLFikd3VrIl4piEKhSsSDAVIIJDBCoJ/Rm72hfq7MBcd5FlYWD58EK89GBXwaP3rNi/4x8
LPMqcK4cylhs0/COrvuIRTWoOHtO1TKIL3g9+E0KJL2QmwbT41xPEv+sZupiZj62dxyNpP08FSNo
7wncmQjfgnlxEZYHVhybBa3J/ldecyrjLSbr8hWvXAp/EoCG2e3C0gXb9t/DsC6l2fjtr1/3L4Tj
U0lYgJjJR3bQjPIEX00ne8skB/PpMGOfBtSet5ZLP15OVsGnds+RL7lk8vG3LMJkhNArTvPCR9d/
DP0+HBexhN5GZ7AJ0wRD/1MGeEmhpW1m8ZAKRGa/fXcBz+OBal8B3bIRKgyw9j0VP6q18G9jRBdF
ONgSwKheFQXTBW9MWgqzcuIFKgQiuNa1suJD0Oi5zpECHKjL/INKzqbtuqGPzlHZTCYdMIAqpq0t
zjsL4cJjoQpipx5oLIkRt8fnd96NwkpHRr0eyh7JC/M9jJLIYtRxjnRpST/j3htsMnBkgy51xEUQ
+AGgOwX22EUPKqEB+wR0t1jVW3bHf8CsdzVa5gthq/CFm7e3dLLYhAFha7LRUhZv2hRwqdTbXCuB
FAQJNvb8S8zRD4r7gvlWjwBjICW9Ju8+uDJhKKuXBslHdXQGbB3vh+Zxwk8E3031wndzCUrzRlDM
rk9jgBwjrzgf7g1ioQTlxDz8lEK6pU9Uf4XaIMAShk1jqdPoBiA9QV4cYTy1EuqkOGaaDtwRyhAo
OfSHeHH7/GhE3cO4zZ0wI0Wb2bCuY0r5PgooWaxBSVnJssFkb0q5aNBf9LZRb0B34XOtfaClpoQE
T9ZdA20sUlAWAX5aXbkMhVzmBBd+AWQhw6PZXOJtE1szcqYUKZtCRP5cGMrOTz53afX092pPNVw9
kSfY2Yc7PqrgIpt/CPPW3r4WUjmPu/h1RfxmJDaDUP9L2zO/CSM1l2L6xnQBsVt5v4T32Oz7NGtY
Z0wk2HZwfGFRrO3xguV+uqEal1e1JSbf36dcrau98Uh5Hf2bODtpGQTQpT0TPdybl3Dle1/FGjxV
BXsrvahpVow0Z+nLzzLiYzEzoRn3ws9fCRE2vBzi/xO+wvIeQROstHbipCrFoZMourx7t4ljASIw
eM4W38LAfW8IV2u2zpeyeXxUwQDUeHiXgKAl/S5wmHcc2ttjsS20lOeIJ7TcGe/3ZjxYjSXSdC6Q
o8hdvqRsCN4EgWWXz6FZuNUtipF1ovhlj51SmvWkMRAUXGJhfiwl5E1YzpzpXhqBlqHxUeRYWQNh
xk8SCQXmdtvNzvrtDpmW22chNdAjonx5sR2oEw1Hm+fqdp700fm19dOf+2RJz5tFuDEEySE0TNDH
c4iykfoPdZCkf/8sjhm7Of47uEPD01VWFFxLPCkJ8zw75J83zdpZAve/6DqKBRqEzCQXsw2GKStI
kyUePxzwN3qv3YDk0f5g8kkro1Veh1KnGtdxb9SCb95h5AGedIkZ+0Ff+SYUfhJJnEhZbYB2uLCs
xhL1qlNOnv5DlcY2IQQ1OTpkPQJKXgmCjs1I6PiYVde7IpP5AVw4wYphSFEsr1QVL63QPbjvRYQ9
48SQWBHEegEoB2al2U029jv0IpoOvmRqxAxcK56BrteiaST3wKW0UWA75ampg0VpdUPaEzqgYLQ0
6EHd+jK4/5cvzFKGP1TKvDXRQYlX137q0ylMnX0HLo3EeVeedZ7UiqVnRv2T8HzDDuQSSPg7Z6rY
msl5GDqyIWYK3y23uIyjU8OH5JoJOKjJkKunSErx0EV1Z2M6/t5r8Gp1qFCivz1QiF4cANW26LOW
8Ylw+QxYG48sThqC6gBTsbFa896biuxxBU66RtdROCSLmTm9HdS3NHfw+hMlp4DMOJVVSt51w/N0
jRhC11NLtx3fRroYMSeuoxC1XxS95vaWub1SY6d5jBAIhVtYGU3d4fQQ5LN75PSHQWwBxcPZ6FdU
8LFJmcTZe41C8X6sajCbhanONAJTPQrCeVsF/dZkAz/jHaEbNYIfsHN4nTw9kgR2daeVkvuJbUT7
KstlZwqa5MW5fHFAUhZjXVlgLKXymVLGQHQOWxnyyqM4aETg6lsHEqWFqGtxQjmP7UkytPHGMHvM
/sU2g4Rh62+VlTHh5kveYpfQCZZ47lU0+YZ5MTkGW0ypJNetLlW3+40GWn/pbkBFdjdKQMVm3W7a
L5IxNjvSDYAgLLn8cUFHVxbKUE8fAeMPflB9q70YcZhTegF5tm9+AH5+ZYXxOebf4qmgS7NnJWjB
MgQD9p60pk7XB6ZBajcf5vQz9Ax/gYlHPN0l2UW6l2L/34WkCHKDd4UGqwXWS/NIdZzSD02rhjoz
nYMVdbP6aHGPw7zEeVz8jtm5sS2qVAqKrdxTMmDQFGlp8Y077nWz1xdhTCoqeN2TwnVcAqTP9OcT
ezNGsNWHi3yNAl9eQaEKzmW2H/4XPNIZWSa7w1FlRZBNAvMs13snKJx54yC9jzN2I5+g/gPM1ROk
5kq3M3py/zWgJ2+O8Yuhi6FYPxo5lXyRsTJpIahEKDHmPUzOzZ65qScD+vw52TPjD8OBB9175ME6
OPJrhSkPEbsQxVcdvlglCAvwBX4rgFSKf9vztw4n/HcozyLIjKYAqk60yhtmwmkNROV9npVYqLZs
Vh5UtqgHfN9IsmU4INo066wruoCn9ksEzFb0Z3PZHTgcg8MeEYMXHKwEE5QMYDNa/EZXUQbnSB0e
tQDlMzPUyN+tr4qL5TLmUURCzPt2ULGExp7rdCP6Ju4UUSYQ5D2Gr4K1Bk4b4zO0sDrgGJfk5v6H
vUWKpGT7TbRRlKey82rPdNONeOzZVP2r3iTrjF45fkndDH4V1pagWWz4Cpsj+GoTXT8UKX6AWRZd
Cc7ZbzxIVVDoKZRBgSYGu3DbWOLbgm5UAsdESwFfF5W0XO1upJWWd/DEdyJBeXXFHsWcDB9aioY4
FitAy4tRH/slSROlAWlIf/xAD3E6e/oNxIN3CAge10xFhQn/xEmxWu0kqWtlypOni2ZNbvPOUHzR
747D8lJFEwUYIoRsWAG6Db37yj4DT1hF3cJQLexk9PlpFWTceCvlhfHQ5zBJehM1tir/WJrr9dCr
F/CIet7HlBxn2BKMx40+tudzP+1nf+UBk+A8Z8OJjWJj22ObZlSzwK42yU+NZSEavbx//VzUE1Cl
BLQrR/W0ifjYr80VaCJ3/wvmtgQYQrBpYDrpjyGkrINo5YRWpd8UabNASOrLPSZMXV6FXKj1KO0N
KlKmwT7nD2FH8aKDO83km3h0X2NPHWH5vFAg1H3tBzGyEc2Go4lNf7utILnurNnyoXjL9ra7DYts
l7iY+oMj4iBzaPssGSHd5S7s00UsaMhIyh30mWmMCbu3tNsxjtLiqAKwVThY5Sc1DvlXrCoHKe98
SroH3Q0Gy+DWs2Es7WZ1k4sd5aR6+M1DiKg1HdgFQysodJqRdOpPALXH9Gr6bM6jGTwaFRm9jaZv
fKrpRXcclY+80m1VUNObUxlTK9arjPysR50VpC0nLi+ADrhD4zuo1XcP47jgNU39LnbJnUi+CfP8
O/c/NImAhxpxc3/za363CZlZY/OCXvuXto/L3za1BwWiH7ITAI0eMUo/erGixTqcHgaDAE7lRqJs
8qbAIxBdP0KijmuskORq7p+zKr51P8j3NdxlVIPasVo3HFK2D3LjMSGrdoKXi65oVyzZhLWPMxKW
RzWQgdSETWcN9406NHiOb/5D4tdvO16IXu08r8T4ng9AhJND284Lgw2Yhmj/UwjB2tuN57Dp9nV9
kCBIclk6AJbpP0gKQ5jJeZKP0FQlepKzNWxQWgWUL9eYDt7d197+RYSHhiHlbQJKZULxiKPeAuG9
35aLr7RyPlm+Dc3py96B+xAVVYgNF4vpbpLFCSgNtZjASoBGvOAOhUVTSPlwMZNNhDWDZdTOW/jy
Ee78ZPU+pRrIX3OuHlSwMQwoFLFTR8jyIaNSRLAg+17ek1rtfdL7uTHXBK4T11e/QK8+g19qPIZW
ELx2GXyIlyb2zyPMnGBpvFrwNwKlJIe3KzQFNzPeIsvMH10Bf5hCyfYWCDMj2gr2HlvpUamFEZTa
SjFdT8qsDp6iyZ5h6xigyeteRS/wqcebGYYEkd/enqUOc0ToxsR3YF5esX+xnOhJIql8rsO2wGIi
G4HdYwtFT3vp5TmQkWOuHD+wfaMF81UcAl/BoTEmSUwmm4LUEiub9b4OdOUXV+IFa75TVkYsKqn9
Iai9ZY6A0yNa5M9Ddcie8ePY9PsMkExARPtG5tmOrLdPACLtPHMjBrbiqJpERJZDjNeFa6kq65vu
gmkEhOMnjrt+nJ/ETfOkRZTYT9SqlprSTOz1C7pHEJQBaiQCxWwqLWTNVBZzx8HFs49p5Twpjc2I
se8H+F8djP+HV2tOCWmrcgbzcVTyb0FvhzMPcbaFPvednjcfZWM/rEHmDBbOWTesiFAuLo9v8kFw
SHnLFxKh3AX//0P+wMkZH1JKZ5kl/7Zh/Y7E/uiU9vCRjP0GGUNJ9L/4U802Irc7lH/08bXk3reg
sJ4H/WoqTz3OYXojL2jgYNAT76APOmVbvQx34dTZmeuh+GVavc2fjyHhHWi0EJCV5q8iIx1KYL5V
hyzPb3bbeB7jop8mJIM8RWHRfQr5YsOLKcjbbBpGY+k2DQs/oxYTwW2wmv6wfi6GGpIscFAcvEm0
8TSy5OYKjDcCMz0+c8MTDmAPNRnWXSC1YPZ260aznfuUdRQOaPYMrCy5vOCKGIOI6t1FsA+TQOwA
w2UuBl2zVftul3KJFII4WbXmLkDPeKATCoCjfrRZqerfR94wjFXTgaCjEeG7KnEL0k8Uk+A4SGWn
7PBOuIBl3GF/wEaR1VhI+gyGSV2t2tPSpwHfnKpwmAG3/ccFql10M2MqI1TY0fTBQQcA72ZEr3HC
8LPHyKvF6YPop7RyHMTNdjPHGQzf0EMJAToVhjKtsqZWMiHdDNGlUBuBqGpEGXGr0rPK7U9KF6SL
ryaLtpgm+CimyMV9yqxRA/giO0IaYN5yv6sfJsLGWhmk0+zIBHwEmrlpUlpSSzS/F4ffOWyeTMzc
HDcnssFSEyW95wIfe2td8Adt9dyIyf9SJjsaKeyL+j+Q6wMNEN+JBy3GQxU3/V0kfP03BzgczL8N
F+QvwNzmpIecmy0oSb5eRgR/vpjQxIzijm7Jnf6siqg5KV+4I+UkDIWArBZ1CBC46tG3nVbrQJQF
qBdS6dadItvWZwqzBPI5qQg5Qp8n3bc+P2r+jmraciMLWwACLeSWcrdKbYUt9SLREYhV10po0gfq
KtU4hJnnOCI9Wx/L/SZQRY88OAljQ2QPy5wJzScyQubqRQt7Lv5J0QhFJvLF0Ivuq47S/kKQj062
Y2PXIwKoysy6Rg6htO/16XyPHPr1opIqevZGk1Fgkzy8+vUTpVyUWneGIbtpHBpnHQEJ3CA4ezLA
VIRCa0apRbB8jxUPgmVCUrEsSo+UQTkKDierlQgwhVpiDoqr1gTW06ZDZhu60qr4fr/3n04qjwyX
0zmRcuVk7phq9dE7JtMU8bHVtxqSRui5fZPTZsvY8eJKGDu0WxNrcBZXtubBwyBTLV08YUzoot8k
+uJ7ApMlr/hix1j7Q6r3yO7Oo2qmhQd239DEass9l0i4r2Yna9lgq2psf+cP5KfxWdnR9PzYUqno
cU8TFhRmG9/rp5zDGIstlZ6q5Z4qzhT86nfCY0dCVjPevrcD3JSU8C3F71MERklJ13BvANPrpJXz
DECB6WPO54jOD30i66v1ZF3tGy7EFGTvQYB/D4eqhrZnBLIyy/gX3Qy2ojb8f+FoZu7HnU36Bqd4
8crP1vvDjBWUl9sstucuEqVJ08fv9iMGV3wsf0RCOSLDyao/4R2TQMCtxf36Uv+m1fIg7wCp8ewt
RKqxbqkJ19+9Vp7i0UF1iiV/eyqYy6okH8ctklVE9EVblTmy59PPAJDh/hHt73wL5b/0s1pvh+Ie
VelRuWrIFX33QSyIIVgk+sDShPKr9Lj5g4DhPpn962xOiOzcAyOEzFdi46x1PTYxy81PNydEHo5V
BjtRALEMhnBV8YpUe4gtEeIX0v8j7/aHfnaZ9t+DNhyyiNsfRJWKVxWqu3nrRPa6VyJDPtpmqhxY
LlwygAnP9n4nxb3ZbUWLjrVmLkL97wM38ikWx5KL5tFWe1LXlVzik4SJq34Xss7/0QG+etaNGWYz
DoMyiiwbC5YFKWbLolBn/JhXFOjj+FGJvfEHuxp/ot1tN84EXwOa893P4YoIJBS7tOUc1SeAqmsu
s/COQKiABYbwXdnKRxQigaHNgs2HqIJgAErLNeChws39h5LVGFvydzfNVAwL2taOLCtrUsX+OGct
ppPlwuYBGMCZpPzyuqOvLYpRuaLV+W/Nx3bKGhSwwLY1dY73a4gJlibPHP7q+KPBhZuaAbYdfAC3
y9QBG4Df+TUUuQmLRRPbAOWXvk+WifOUHNe6gXL/VY9vN0J4AVaceI13RjQgS7qF1krINqE2bRUv
LO+NE0gKF/V4/21xDMPbAgpYtnq3GZ6b2njeRb5Mle0Xca+P9nKfppP6+gbOXW/UxmX95SS8+aW2
DTsGu7V2r0ZSNUXT1zuxjFbMCDxpKkD4Rws2BeyyuPpWkXdzt7cHGGBt0kFLPJAZYXFJ+niyTu8V
HmeVOMxx9KDY2BjJDfwHV+OtFN06ZL36asECJ02AB2XymWJTWDrezOMd1sG0tPdF8AB3XVtiKLU8
XVyWpsm/3sylivM4hbhBTP875wlLKMikI41PQfMtfwALxSzxGtb2qYW3T8A3cGGZFXcsRxk5QmYe
BeFA1DFp97oAvyREpWqV1V974/B0lMsWEeTiVX+oKKhQ1wXj/f+aO5/v9zDVAaOCNfyRBqcrwzC8
zzLd2wnhiC4SOp5Kp4wDwaDCxU+QUPMFh7ahiblR5RcnZZUhCFOOj2/6jM6aXCrzDaNYEba7qQcl
ZE8PIiQxHblfzIHsCONDKtEbB/J9W/m7v6iTeNy6o9iv8FhvbMd/DY0iFVYUiieioVaQgZyybPT2
bnwF3Zto1V9MGl+eSHZ8RvBIyX0Mf1kzAXF17XZpDV5N6Kbn3Y20Jcdn8l9v5AkU8lwrHM9qMOQj
5LlZeC4QArXNVhxGM3RZI/ZPSEeYh/RV/vB/m2bNwEbkNI5ic5dn7hus3uEjpgxcEzolmE53+L2+
p+RrSvHEzdWc5n/8zJAt/hffiHp2+aEH7UH7K6upBV9Wm+/7peN4+hcnOyfwXb7NceWpXIYDVm2T
XruMpcw+ZmK2Q6NHpPeQv+Dorqhl21TUZeYJpvyci3P4c6T6GqWHM7s+13LzvbUU/vtsZnegVFfh
kNEAVzZo8RS3euOoQNVk3BWYx8Rof/EizP8Barpq2KfNzGhYC+NlquUx8S1zd/wZ7bufG5I4gTKd
CLoZoJ4vc6R+T/+LreURLIGNLzLhOoSzNMpQXTLSNrAxsQyjrFoVyHOSPOtsrxyAKIgI0/mCbX5X
OMhHXlJEhFZMDKNXgXoH4yFCSSSKrEE1ijFSi02YuVgUh5qgUwx/VZFAiP+yOjGlbAbBb2Wt9CiJ
H1R8p/rmRB6Lfx3gv2bzw8FcQWnczHFdcRuVXFADnvku3MFPe8Zw95a0exJM+3b9UEQmXTtYgIif
ArJhmeuZLSXqDO5NbHxDbUlCb7snNOeB0y7zOMTaBeFsL+aEDxl889A2vcbYK4auxga7EaSoHRai
gPL1LAE1p6P2re4tT1E1vVgY4BuOgooNpUaQQ9+aGEyONckwA4S9Coe/eF5fJu0YfOwVPgxlwNG/
Stt4UeUJ5On9zm+9M++Bqhw1k8OYSN+zV3/UAbbJk9fwIMWr2e+77v68QiL2JnXqOuv+y0JOVkho
FIUMFoJAo/cVO52C1T0M3l4R29IEeYQHmuex7cWcxUz4yJKFyE+QgS+kCw9ftQ9USfaac2XtGXSF
3+5Y4DO1hUdOrArnl5FDaf3iWRVDEDITHnk6Fph+mPUAn7ZJQlmsCNpXQpOd8/npYNZC5Ay3jLqv
0Cmy4M7eX5mGjVU6/Hb6Pr2Exb1OdQYprtxtYCzVYBvInkpU1k5z76LDTE4Bbmt7DsMHl0FgPJ7N
bRtKWv9UOcC12xfMgFqDnBpr2dA3FGTeDYjK3Q9dSXE26Ah5FeevJCx+Udl2mH0kJ5cNC8tttRiS
JO6DOqaMvVxYbGcXNtnKwYAzSLlZ1r2KWWmN0B/f3fb9CflPbOQ37q2a49mqXUTW+Lc9q7v1HYPb
/sJiIegbfzMHK/I8ai8yAQXDGMEDr88YYj4kRIih2VFqyahLsdDzj0hqy95dzRd1OzpRU6ofwVb5
PkvZedB3xFPAOhyltfi4A+DoXW7zeJy6I5KKWuYPE3p1GbjoVMbFhArxfdaKRtyRUacLpLEZ//ej
Ulwp1UksE9DUh3l827ewJvsAo2Mu9v/xu4dj/ErlqzxWWOPazHvp0g2a9tAOEox/+q4rHdiiVPG7
wtsvuHz/5DiPoSTqNRtuBTiMLib7DC5t/AggGBWZxfwGCEpZwM3uXdB+H9qcsPmkbrGJIW3w3xlx
YyE64mAoQAiPzKPu3sj7JU5byqGji9Gni2T/OcwmxIuFndSvyAZ3GSjZFqlZGd1GFKaZUdpSqivX
3Qp7vcAZrbe2scU0Yx3Qi930Rl3oroblijm2/N2cRnHjbcx/kiEaFC/BXB4L7b+U9K6q5gYQipWo
I/zniQstOFkd9vXXg40LTCXKTWevMf0vHeo0tcqvwSsCbjFyUguH1OdoVcxG7nzwd8vND8ztYEM7
Xqx3xK46AKeq3zGoRNUrdwbXw0JxuHdLsw/0G0/7sPpxoeYOHs2vMM0StFOsg5Vzreb5/VKqkphn
xhYXkykPVQKM93J6wAlHShxiV38EQMVK3pj/poFHu44XNeoqVmOlcHeHp3MY7RFtIkW9Gj4KpHQ3
N1RAbnKIEavFv5pA5hvaPT+fhaQhES/xBwwQi1XCmUeWzenvJdindyFslP4q9kgy3ha3d5etImqG
RJ/tIRV89ZKdPTgFFZ9rtFyagvyv+yzSB8vAairasTBLkRZlCF5YdcWDfGi+roHMPBJcVKkTu8t1
YEjMsTr+xg+d9fZuZQrlXMB9PxtAtxgkzUvRLUr1hDjRnm5h1HpcRGHSQmL1F425JeNDF6vTQQD8
5U0uMiH+TJ3m0/9wIz45EPxqv9YU/0YXr0zMnWbI0cGe0TxI6RVoXutcxed6jwqNyDW6eN5hF1rM
3FlETREdIpUC2ucyyP1jSw6BVtF/uzKMnH9Xbd3FXsz/PSE3ZPpmAMYP7x6AG/7aHb5ornzxQOuQ
8j+DRxKWXt06E3JPJhS+4c7i3ZkCM4LjcXXo6TncOYObJMWMbwBULN+hZBfuncJrAPyJXTNNRoAy
nSDD2LklthGBVwXPTDGCmauJdAnq7q6BmUxSvS81EvzCgE/Jfr4SndzTrJUQY4ZUDl2z3r2VwaB5
QhqPBRx12ds6bwt0L3mj5syMX+hnRuav8VBz/yTER0kF1qToyamU8hFdB+NwYSGsfSUdkDQsPTTT
BXk3sHzLUbRy44wEqRLGaHfc0x6bac2JApJJzatQPaXfE2jceD4MMsTVBx65K1S9PffzhlG26pLd
/jtqN7oRUQAQutgOQaPqU9K6sx5a/Q5C7PatzTDUyuD5R7dI2S+N9M+GO16sas2fQqmeGDyVb68j
IFBRqKFXd/mIt6FSZ/XGqWtrbEdH8A3Ou5AnYne6rcFgKH98T5HcWX2ZfRn1ArXV31nGJUq8HnoI
uIl0th1C0ZiwyZqTzkWmoUZWG211KYOHP9t6b4Db0lIkw1t2x8Gpr4A8rqjl7JRwmmUe3ijIsCdf
HQbW4sYsDNIOS1735t9I0b45ICD31njch+5iVeV0gtUk4bkv8NCwfunJ4VJAkFnW+Zg3cYT4rlhN
4uJSVuBZokpnvyN3UFoyfk98dZyCIDR6XcudH6nIQlcrEk1dvNiNfGi8N+cxzUqrp42T1KGL/2Qk
Kl1vNu8NVWX9DFJaiUOEylikiqItw7HAYZam1VzwasLomHVJDo0mgc925yayTzvhKYfoRvVGCCRF
LVwBVP7/NsQ7uQqOmFxDb0kX8QVHKGCk1bdTyGk+OmYz032EB2fCyY1/qDi4Vq44idmL9RbLoKPy
24QOPa2fU4vEIA5Vs9Q7Ys7x99DufYrVbhr5/V9+ozO83zOVF1zgBlMjmGjLpd3pLrR4L8VfiVGD
2vPFVoq4RnrQW4fjwZcB8Xh/nP/huzn79tKXVl/4dKrXbz5ss4S+eOKiJnFE/2Y7o31Hy0BbkR+B
DuIEkLEnDHHr6XYN86fkLaJr1H+VDRoQEdhfzFHyIU0/SxjOk+yqKZM+MbrJNUKqcV+mZxmdB9Mu
sPdRD5RnAq/AGe2wEpoSzjAeslvtIYU3COIHZndl7xeN4yFpljAd6QAAbNX1EpIcbJJ6kuARR63F
GelnM6x1a7f1a3QYV7m3Bpi5uGIHkSPhBKAXE2xRNAENMlFIhJjTnm0L0Yfg3+7suHLNfPotDj5N
IHnXmwvE/frWeG4ZuYX4Nf9/qs7EgRnNdFVA286EvFWQfosGfuMneh9jALnNDgaTeSrp5vQUi35G
MKOgPWf9hOPThfSiKPV+SVjlheSZ+Y5AoxvB1OHQn6c/RvQd4jmnsTI41rjeqdj4zyTF3NdmbDkH
Cw7RumeOep40zFaEXqgHznVQg4u6bOAWaR3/EMkY1jbC9Q9AVFCAE2Bt4BOzc/3J34botLtqEvmg
516SMpZksrDN8IXLaP69Meihl6low4HGpOnPGxieS/ovSkDVyfmi4/OTksGNVCUj9QMZp1QW/hwP
xRCWLscze3z+G/4SPELu/xrInvZBaAKY+dOlHrfOMfI6fSz6CSi9ErcVMs3gFUqxw3tVQR3XW8CS
zD8VN5ujERQ4gb5l+WPHqbIoIXX2LRWIFnmQx31aQ+NqjvnzeFKtug9xkMUhWLXTni9qgcU9Nl8Q
5j1QX/5t5Ck14OyhkHPfeGVBSfVLfeKhvik4n++Tu2ID01FwJiM2kRpEM1ZMoRg68aR/RSb1H87b
1zoaMrlHXaLc92kSSJy9NL3odf3VGgs6gxuct6OHQ4OxOukkIk4aIxcTzsyX477fw46GZCLOV0EQ
J9xquZhAibZzZyLs+8GGuT0Z5S3bbiDnoY5qBXviKeYC7MjlFFg63OS0UknhUQD/7/Hb2CsiFDj8
GPBfol0rEdG2QtyWambC7/u85iUqBckoTBVpqZ4d3ERNEawDN1jKsnelJ3hxELq3/WSHyDPrw38J
1wtH015PEz/kIogQLiPJMfZHMu/yn6FomAM26dC4D5Y3mHTcj+TqBKyrg6sOXzPTB/nqCIjgkhwV
coMWGbRB8RlWNFyj4IzZCWEH4iGnsehKt4kR1iIx4EY8MW0VBless7V8oTb9QTddL50WmcJPPcCW
8p5gflCPBqsPGzP5fbWcgoSQUT/Els119M/NKFvk77gtXNph8IZgbNuDiwNxQGVbiq3Q3jtw2nLW
9Kr9mJ6qTCH9YUn1T8198DeUeQ70/KBoeixyrfJN9ctMZei3075QqMj+meXxeg5VcSD++6E5loQt
V1X/gIUdVenuyViJwfqfM6U5baZeXl6HtrtgjH0QCBYWF6wS9NacoVgqh6CeL4IVJGtv5rQnWtPw
PjC8L4NsphvdJbIufgUCbASCb8Ir8Loly1PgllnbiXDgIu+d2sdXSdzyHOnKUVovllsbe2CJvqFt
ckAhYqszvq7r8DLlurgeIyadkG6Ueb2Hln68Lr1wnRbaj3ylE6yV8NfSKmL9YIcXJ0aPLW0jTWP1
OMOou27VoQOuoj+5i1/GPWkndg8QeqgRQG2rAOzo5UtnC95h1hjnSB3RSKpqHG7x5K8Pfv8gKRsD
ijaz174Cma9gmJsFTzSmMLFBTdZqln3qsNEBekVmoW9vxBMF8PJjQgadO5o6zNBm1GwhnzZBpbjQ
jIK4fkJ6ZflPNgtO0sbSg/rGnQBsf90B22SWFHQJhEt2Tu9s9o//PgWLn5pwVoDfsrf5PCO+oTfC
hU21wQqYGSNUvqSdegN+seKgK+QbReMykRD0TEFzBAi7m7c/zVYVovTNeVOXecxpidmssNeEgC2E
RlQpuxPEh7PdccvtlskiDm2c0NnOCqrd1ZqcQfqAHTm3HewGqcNs8AGh7vLnvXjiDrn7snUrXqOU
6O14RbXv7Zhg3bYQqmIKzw2OwdJ0rj38HDfBMMLxkmNhLkS6bPn5mskXv4KH6lK7EmrD4nFWSBdK
8QZyJokjs/xqL4cWCsXRjAK7G2eCvCnv1FQeGxNnpt1hbyiJhQswYLgsiNKSITALtKXmFTnbpbXx
Gp7nM4AXHKYFWcvMmTK68bybTdUkK4kfuo+Tdq06AZdh+hdAizvWlViih5Nom5CuJUUgEcfH3H66
gWR+EsPa8LYLI4SFqVtF0hba4oM92lui3GDeu+b3Sdba920QdOeMZ4NpwZEjEYxNIqC8eHrAoVAz
g6wRr3bCT6aGYpqu0aSBJ4v86fX2f9U1c2kSQoJHyWaUb+Vcqpal6cAFjQW/6AjaIFo741jK99oP
qYMTGWdXEG+ZAJvj0WO7O2vXE3fHbWEUoQ6QKuozmYV8OZUVRGApHdK+57Lw45ripvfR9k98zrqp
CcizQtAuTuC+5O26ZCdRIEplK8TCHsTlz82zcIvRhnRtmYUxYE5bfQxvQJd5LApakBGEiV2d5y7c
I5RL9c8Pe8ZDYF+ZCQnzjIqVxZYQIHzrgL6pR2hZo27gfqox3siQNUqT3T0IKbzMIIkXWuR7CM6R
sN27H8QXJ1f2/958JDIDdsN8UoV4Yz0dkczLl9o7QJXlFEwXvOt2pmJegKPkGBRkIm9785bElqv0
JoSxuxPCjnr/mETk9sTMXRgB62rUarqYQPcUbHssoFwgjq4qzfmeVmwtUbIm/ZtByI62nw/AjEYN
xoM55+VO3aVfLCeDXjLQfGPQTevEOBCpIh9HSEAC9eHS4Utm7m9rDyby8FmQdIRHz/yRlIS+I28a
nYYAdO3dIuH3INm/5Hfy6hAaezgpnkGTevFfitRCIPlxHxhqCKX28Xc6XraRhmsFO+mxNSawgpoC
XXtDT83Ys/CdzEA7q7gOSuCZOxzXbyeD1LEMjb90BbAfhUKSOis2vq2fsJajCldvzwq6l1zxELHT
9Dt962499QXPi6y5T9kxI0Byp/JJ3f5iCaHI7ij0n9qqJRGl0wfTw3SMQPRWwq35UpG806PW34vU
SHPFxB+vSOp1AWQT1nHLeOh8xqQU5FYnEtjT7Lqi8MndKpO/iuOfgeiEHucWWG6RpyDbQoTeE2gb
I+GRJU6bAlMk4BoKeMtRZe8m2s8pFKwx4hUO1acXwB8yf8Q02AxYxik7SBDibwFvxAqLJJEJt1YN
d06uPnsRFlYH/cI0bbEOP3FS4pPCcuE5r6mYfEL9Llc3rc+fhZWTRNU67EJXxPT9+Znb+h6GpzHj
iAory4DXBpk5otVyl7U6H3ynApgETupcIYoGqxCbfzBpnkY0NT3bRBN//miLhfy8WdgAVMQwLNvy
5WiHbRKyRpURaGLZjpOPBijJ/GbE/4hlwTClsfdVzIOesXDF9J9Eyiez42BhJ6AOr2oVDjR+RJEA
4ezixJouhYqPo6hrggk5kkqEpYuaySJLSjjXbLmJCoa/NArnteQmT2VzghX3ZgeUHrLCuI+kbal7
rLfGLowQQmWDCE/lijt/gPxuzmhCuAnd50iCbgE0PACv2D/FB3XSp6j/b6YLXfvZsXY/2enZRhLR
+obrVi1jCg9cE+sk/LAQZjqiwr0z1I/NOajMIrMZsSIxaXeU9YJ/itrem1vt6kZEJXbcxn3eTzQd
OrB3obksp13meMxsA/nRuwviw9/CC5Fg1q4eHPayXwqkmoxQtGo+bwjaxmCeb77eNrIHjGODtQaH
xw+2Rxs1eXUwHB/h3pUvw2VwOyQJlbrODCED1ScLuRaPFBDNthYwNuW/x/rfg1HYSYXptKW81r/o
ftThm7HWOJQXhcuALNM/QRP4YXOhLUFUoPR/oT+0M+fAXu2wMtU+th6CMYnSqZO1ChO8xuZPvYOe
ahcNPFvW/NMlnFaPCSbTlOaae4CZlO+YZyHLwgIJVUl0to50MpALNfwaGPGB4XN/CGRWSx+fyz9x
5byf0NA0YNmeP4UH3bq99iRjaj511s3RqxhNDc9vkO22E8Xc3sAqV+LIhtfYgFlpXJ75PirvJjdT
YbsUKwJGRxRvA7BF8nvvO5aYbz7aaR2OSEjaRIRsJNDvM3QQWxWdvEwTiMUF+YSZD1csw9+T7bx2
wYk7B5fdR0S3PlU567TQG0fdcQdETn0VOhaEz41qgLvqehp1h3DlXcC73pzcKVKfFeq5i2NjpIfe
/pM4dTu3WlFIpX8OmkGcm7P6A3HPyRDYJsRUrCLtPa/BPicrCvadiFe0E7TkqOvyFH58LW+pxzYi
zBiIc4HCIH/7g+Vt7p5PT+6TdkRwzamcYXgEeJ4evbKizJ+mr0EOWQljMGFgHScE/yZ4vohAjXDr
ld9XLFxnFsA7Qwn/QpyGezw39mgIoapI6d010Khtuzn39v9I5ykg6NvFvirpL83G24tG1AEM/S58
CTSvWayJCugVsIGSYFsO8WLqnInYTN6Umt3tRJEybxUu3efgm1JOanGwIBpHWgIwJTkRupYsuqgt
FjXaxP9T5qkdL4RelSXn+NzOxGG4plCM22D+oAwz2/WzCu5Kdam5m1Za98FBZmc1ETcZCH1Wl+tS
o3ysFiWCDltZUxzFePhJYbkBYkjkP41DCkB3sB/g8Rcj2BfFIgtW+AUxmiuPuh/iQEuQjGMz7IDV
g/BxRkCGy74Did1H560qYs2KBBOuPRDr4AGPvIr3zcvFR9xOKMyt8aiPBn1U/JbYOg3sbyq88Lxv
dnkP4sIQTyJ4QmqIc1w7cdRt8pymHhZS3SA+i2HnxgiMYb+cGtKHcTa0cArSgZsRsYL2en2id0VZ
ZcjgKWi1crnQTptTz7uX+lhejPe6LWz+/Go0Sld2i+3+LD9FuBZUqqhBKNbzqphPazlOMK0aA97H
SKzG6wsWXrNIcPdOKs03vQUT4VJm4SuSVfai851NEgu2vsjAnI5oQEdU6tkwAdqMjiPbg0nRFBSB
ur/4wxTGeXumqKkoZjFQ9HqLKyuENPbsfUMkfAtfe22xj2LQhiZwq+elXXq92qoDEqvkiU24pMIy
wIW21U0/7fxRJDecU6QAPlqYF7i3tR2rCZbn1aWL7VI/xeWF/MYlcWXxa6ISVXsp2Yv8PbNS01uj
ZMAsR/oIY/wZBzi+ZxIs4Cxc5SKPP+nH1+JruU0RCbZHSRmzqsV2truzyZ+J0QJcqHckg52AoyPo
mzscb6RBNnGU1BPTdHjGQm53cj3Y3zssoep13LwVBpgDGOKbSLxhEwmINE35NA/nRdPJnc4NpPpH
qg5x8fQrcDpKIbboe7u4Q65+eY7nF/NjnppJ5Xd1Kisbqil4SkK/D7pAJLTpkelIL7/k7m5fqAar
tYLbSvF10NX8gPS89zEI0ZrC5Af0IgWClg/AHpkGsqIQsNyySYqEDI9PmrxF41uCtf0px9Dide7h
DakRQl/fVAqm9KlvWJfonJffMuEdfLRQ/XhjMtcpu3gPrksLSUOqutRg8PqzVPBAuKxGa+z+AqgW
GiXqgjBH0Y7eqmOoPM1lEPiLvp0PdO8jqqvN0FPQYeN6ZrnNKYlmeBumSdsEVtY0ZSOuFmBeFtmF
85f2lDjKEZ15oGAVCvTj4z+XcEl6cdgvLDDw3dQMXI844xG+b4pAKrCj3/czaMyTDT4nKlm8Q287
F9ztxus66yODdg2l6dZB+p43UxxpFO7/l0sv7MH6tj8jfmde2Zrd+qk55Qrbr18YWWzuISwcF/Mq
BY/y/l7Je4YS2J7trilLDPaY5Rjbl4vmZqwZ04QEu5oV46re7dFrGJxaqingm6kNgTg1pHidy0VR
5QbZVhMPaE4n7s/zAC4lDHrGd5Sk5MpmrGhUM93phHGPCt5a4xZWQp5NVzuHSY9oXxnwgBXNgsdv
totjS+EyOmrZoM2u73YLCS3N4pN+o/srsz71+8CsDYrENFh0CfUGZeHwp7VKK2DzKC5Gkr3ZNwVR
stJRPsRH27OsqX8dPIf0K5huBiYujQazry17Le2p8HZTLSBf2wJ3o00rl147TIHxVBThRJIHoX+x
VRbPuJ2uiY08nh4NMkWRvgMjhESK/S8qgUySFQ8OLVcn5CnQnNvQW7kM0wUptrIiZ0sTOtpNivgz
AlynkNW7zxmqEhHUWng9YAwfwbj3G0Cw/Rmu4FEFQkNPw1krbFTx9qvu10Mk+MCYPhaP3JbwQTlF
tmpbkdhD753E3fyo9MxgupXfrBODmXuHndw20jzilV7aew0IDpNrXfwAnn0FHtbdnlUMl+yo2ubo
xLEB7y543GYROlW2xmaAMDLyoRCPVG1TISGn3QQDppnzMTxazDh9PjtpAtxWuV+JzmdBgKMoQ9bj
k4hqnKcrVHXCe0SUHgddW7RzxxaL6YyguLULP51CotWvy/9TdFde5hrGocbXRS0rry7+92o8GcLP
NBPiqJurIbTtbfxlFFdM1b9/At18dZLyHgOZ7O0Znzv5Wbq7VdZeNdUDy1/OoDdD+oAVTYdfLrTB
J1u2E6eWrCl0URVWH/J5C420nHZeRVv5BHS8Z2nhuAkmS8oBHAH300ZATepGt3Flp5RftjCwjMJN
QXJU6s6nEaikaUkJ9719Km4SdrB/M7RdEzTzM5jcskOwdrZgjT6llYk3Q0MYhemfYM43u3hsOQ4J
2ur5Hkd5NBxIn4+UUIz9AsFZA7WwdtHuQjJKl6udrazNBv/50EfHuoVNe/P5a5CD5wPU54T5e8qV
3PlEtt6wYFL4+Vp7Mk4dc0o5zfYoQ2rsKgUXzB9QKoYBkr9QiVRBzo2d/in+u09cFsjAwk2zBcQ1
xtUq1oc6OvgKxM6Z/7AKDI/XXABNpxjJmpglvhv2S7ufRRar2XMdfufcOE8fg/ZldfjsYMLjzuoI
P6TtquoEJYRFzRusVuHvx0WRwx2lGDRcTBH8Xkr7YiY6+jphJdft/qyidpVmLzxDIOzN1qZWCqM5
fQsAuxkfTtTpUQSf6qFMiFxBgXBh4fVpHKUoEgSEn8UYNsEEsdIBDmYiwdaHeYeQ9ivbqASa50q9
wPCDrA52ITUHO96WMukhfBLbwRApw35uVRLaDO8+w/85wWFXmPgzR+Zpwvb8Bh0/JotVCvZyIUw7
ZAl4Mh1zhR7KtDMbCotzUtB6ggzC78nfqIHALXDsTgnaEIdfwgN3e7GWXBWtUSSmE22wluE/4KAq
UeiPrR7LUkio/0w5/R2m1yK71UizbNsU4sZRlb+oc/8Dak4xtx/6Youzmmuw89F7351AUE8Eu87C
kwpy8bfGY79kjGIemuOgAHAspvuXv0Fpwx+SxrT3cXSIz3yYhr00FgwFgM2rRNhzeiipupVNif7s
F6fGGTErSOPok/4HHpjf27FytjiOEt0pv7qH/y1teky7UvICrkOZODDXHHRInFY8TpQ4HuOwuLye
nXChkEqufbBzxTKmKHR8sgD3V9XfUpaUa0MEyxmKbgAVM3dTFAtyt36khWwY8E1YgtwW44RXbJ7c
jiEt9VNa3/WpAJ3rUMFKg/zgyV0E4+KjPwny5enEDxLWtFDGCwBIgMVuv9we1UKND7/u4WQLAfuc
AwOdY/wrugXDSOloO/WnCnAJyz9cvh/YFw6FQaHSxatvV1YNiVUfuAitnQXK8LudQNiCaHP5RuDd
yx3hI6LWD6msMkamtf4yPu7s6MV3vJXTVcEO+kGCq1r7ZvujI8mYn9M/hEcwuNgvUz3GOwkb1a4s
F8Fc3m1kydHuy/Q2dHoDmo+Z1XkKhUg5WXhgt5NxzRTKfdMsBjNrT3CR9MBFWO5mxgT7jd2igwSl
vFnXvSaiCJ52bR3x/+fjwFDxn50YabvHrkBJtXkJQ0BMj8fDXvPeuZSk3pIzLKB9mYn4CB/DA8uF
ketW9vQu7HLSNLswn9uUSbZ+yC1w4H1zZ9sFOv+jo5drpCB1WsNkx7o9VQn4Hihd8yUoVs+CEAdk
pJZXgsTcAyhmVZb10NbYL2amX5M06pU+Fpyyr/iRB8siye3FMQnknI6xrcppDHB9R12CWqUmw00f
NwyJ9ZC88MdM4a3c66ZGqp6xUqIpDSR07/PLy+4bSmWmhkw+xD0dr2lN2qLPZa8gAPKUu+nIr7fl
iqAlvtdV6fUiWCz0QZw7+HdXgssOR+c7yZKuLEI+5GjeElWA+N34G98UqtxX5+WsSzx0VRLta+Cj
+ft6IIQ7nsxNArq2BsvN7R2l2krXKpSSfrejTx60Reo6RsfsYVhSj8wf+BHuYBr4T9odgxqPKPxb
8a0WfNwVgKZXxv6aCcuXSNFW2UbAuDlL43BPLmJaFF//qw9oxx7jXkIMJdYL8AujDwHHnlJ1Uekm
Yl0XvPsvmWeE6iqgfdzXdp/Npg3lbqfTTbkUKTtN/jqLtqvIbGCSAKYqamw16mrePG29MA73E7Y1
1KgGoZjozXNixVF4BLnkbFUrKhaXm0TXDLDydcWCOw0Ak27zgE4PS/rGfsRIUTN+jWrrNWorVUkh
Asxvr3NG7IOKzYVOyo5NxHSJddo4S1PjmumMUeBY9Y3osbQh4id3+o/9K2rbwxdI02/ULK67kIET
7xE5/apVyRMQH3Mlm59Cx0Z/tsQyUOi39gDoPL2bpNPsg9bl4KhavfEfNWlpSEHF/9dO6oEREnCZ
aQkWE7pEjsQpbFxNDr75lQPRr+9SEwejW8PP9ruJyPuVMvTokXqZrWti4MzUpRwWpQnRsJdAJuq2
u2LY7c4ToH5YfqG2HAqu6FSNobUzXPNsbbluQ5VLaigwiCVeK4B4eus7/cqkQH3ZRKTykhR9hb/R
YF1XJHj/b90rhxLvQ9WpkihBGfprVi/AbFECKKOZaZyAUXXz8Xdr+8xeH1JCv1I4MYQE0PxFsJ6m
YTRtb9oaQt0bdrdrdvpKoYcpMuPdX+mzb8sxZZd1xzWXpk8yGFpEyrWfEhsqalzaVBflfLP+bRoM
zTG7ZKJ5y3vufoQEolovLU78sQyWSNQhndl0kMPB5ntVv2SkOul5SLYefS3uVNDjB+jkwwfu74wq
Y+T20jrKWS39ZhNipGz30r5Sn9ZPnrm+HgGAiBrRMdpfWQ6lPQmjkSIW8OibY8t8YHyyfLEG0p64
hcRUDSxjPfSB94slkohSUTXVV+q4fJIjR+NREBjKYJjAtquyP8/2R32dbAKYpvbvgE+/e3qvTCFz
DNpMug29MSVV15tVcgZa1rZ8ZTYWoJoqwbScWqmq/an1MTykFHfHAgFxtePqkQGLC0kY9Zy0045o
ba3gbDos9bGByNYsQOYmYAtrLpp0mD8wnXZ2e38XFWbap15MFfY/ZFFH2THv22vUnBdgXIkjtK42
IsfrVes0y84Y6JoaPjKqospW8bB4Hm7i6vSEiNPXlG6IuJ8+HIBBU0cVDAacuc1tLOIgZ2i1hslD
KxOh1vPYT+yJfkzaT759bdcIH6Ta7xom4FhRPjaPkZfd5SHfmnEGU1KxZTvXiBj6SD/1v00Q0NGd
2li6vGukeyp5nD4pfVGmZhPY8N6R+ZNpJVX1/RVkGhEp0jialK6NIKat0JZLjnOuinhY2nlGsCDo
jl9Z2Mac8/26LTAmcrgau3fDNFXG6/fpUITx9Z3PXd0cNJaV9Xexy3hH2S2r2nKlLxLkJZ8G9ZnD
2ZvJpYkDZrTdNUqOcH305m43DjnQ6teFpoEOX2o8nT/SLjxCaLt+zCsQIOjlNkptdDXT19uC8Egp
OPEQDNasrIVNQs/0PwIhMAeOCOZeHKrbKK8CNoCv6NoLHzmbC9ZJk/2zTD1GQWVVTL/3rA5CJ+jj
V5pEAUm3/5GsqPAIlPHsEOEIyIQ7UOLCttdRxhVH3uvzHL2scZAmpwoWqu8UBWm222VEi5y7vTsf
VpPvQy1tdY3q9Q7HIiwjHmOc6TwhkkSqikLQQXECghPG9P7BDNSy9VyRyfnNsDgDEKoRyplxysMr
YB6jsyMZonrBeMBwXN52ltFV6hKeMEFzfxdJDPkovjJPdCuVA4PqWeWfCE4pFPHHQMTaNf0Josk3
kid1dh+/pouDbkuKyrtikp7Rahs+6HAPs2YW8O8SVqIM2SsRYLu70SOFvJBq6nFzvaMBKEEeau6T
wey9RtjuJFddnUw0PnycApGTm/KLxtLMGXKaQEpfVbUv2DS6W/Vh4nPhRhmwYZulAHXZqy/AkG8L
xPkqhsWb1S+LFpHcLyPDo1s00u7W/ZqKvxchlNSWt9u3eIzxm49VkV61Lsd+kv/f001t4+q1uF6c
eWHYuw4erCybhmFRiK885BDGEW0IsDik0dlq+IUo+9i+kaHpEPb8CIelv0SjE8nUNu+R8N8NXEeT
vcQpTbKvoVo5S6YtPl9bGbQSEQoCIYSOvq0y1emZKu5h8GwPwWCFiVnzN+WWpnyuT8NLg5RQHlRV
qubXeYkPNhn5yTFqIlG3CQoYhoBzre69t5UXPnvMLMmyG0SNPEqpwnktfUicrF7FudTwXigSWq19
VDY7BmB8NYRlQHQD9RUFhw79MsDpCp71gODe19acxDjXHOnQlcLZQW49Wz3ZMNzaOPUt51K96mZf
Adbf4PPJsasChKuoQ+U2vYH3H+8QVBc9QIrdWLHfehnpamOazZDIsGtdzfJvMtf7Ul+BEtkSQ9vy
FlolQp2cakR2aTNpW1kOqFogO+2TRTRAMbupedScGD47Nn7aUlc0cJivALAIoZSjqxTGsarAcrdE
1chL2sRbl7VKXYMbkQDmOnCPFuZjrWknwidZ5W1poGabnM7Tz2R8L+3hPoCZgia1tZ9M98r/uelK
3iJ1cx5WJPsrleVeqb7eIaQpBDz/u0iuA8GCyan/N27/VEt0XHwWamSkzqlJNVZftiEtoIkORqv7
RSPwvY82hmM1uIQA4xVH6yeoY5T0rB/W22z8Ll5/ias1GhKkozD1ForZxmWq8hu8QBh6G4O3RQ+d
nRe5byjEW4+uLsa0dlVV9r89BlX9+fmvPRGLnCxavleBMe6GceYKd+RKYo/GRmjhyZjuW1M6Q5zW
ZJpy80WXRS1cznnj6dI4KFLym5airyU4r5MkF2kyOJUbWMJZwYi1hgfG41gfCQTi/3xO/dCXtuL5
D5npT6wJr2Zf36/eVVmj2nLQAsbC4d3o52l3qjFuhvQj4Q2Kwp6Q9YvW8Ixr7yFnRVtw048irNT6
MHRnThE1khKLQ6bZGMjhdKdEsZi6exhyCfBxA1aXF9SXAKJ96jC2ucN/yPgz3dpr/v4bXCBvbwqJ
gWnte5Z67e3lFKME8AgAv8/sl/t7pjtAX1cWChpQBbiOExtvOlWBOAJJs2YgH+HkRkGvlCXVTYL9
ZZbmaua9mkcKcEJ2eaaUqs79Ks51R4I98aJYBY72325R+gCEtZHxkOKXMQLi5FafS+sMuilSacZ1
+mY0i+ull0bkd96uERmKxinInamhYe82Vj91r3NLCaSMMihNVHJxGx2PXE2GOwFXgNcNoAc2Yp4U
wSF5XvtYbCugq+JwPgF63THk6JfioZVRG5O27MvcbKJ19CrKL7JeZYkdjBgzPHFH5JxGr9nk+cBd
QYzHul3AJz6LAGT9mg20QZcYh8STnJOCRkudDy2psph0fftQEG4bVeHvktjEF2PcjTNdK++rGAQ+
3FIlZT6Z+Q4yOYCNC51AdfLRJLExV6L/mRCwarPxtJ7DWe/f028luw1UaxfQvkm9xXIvkM3dWnh4
A2aw3SGr0ADh2dyXjr6GOjM+pkkEcxpnr7JRwgCEkDhwpcF06oWQs0gkBi5tlqxBClSPPO/gCy2Z
09h4c24TMK9AZfeo7jXfXYTmoCxVPI2O0OiDvN2QEN8w66ZvU5WJteXikME+RMjQncApAZKtfR+q
CwtmqShEuHBjmgkdsTmJ5fNrxmeiR/D89RrH6AaSKXy6EUxI23Heq7Yvq7li3YtKf5LjdtUU3HkE
lWfOZxBZiP6r7iPUSekbuHktBUg/0pe2RJPqJxIgaVHxzFSFvprYzBk1z4uFu/sje2RJilhZPqp+
OZbQYPDfCpenpksStAtZb0fahaJR9uPSnTXX+Wyb/g8RdDS7kP7l+/0STGLe18XpbO8SxGcguYO8
w22TiZbGhbn2CRxHxzB+svVFqWmUtlm3EPPeW4ITuBngrJOdgcygz5Zkyk/yjwEO1Fwnr8KjbSiW
Ro0GAt7xATFrga1OxyaGHssR2Qh9D/3IIjG/7xDXoney+ju/NlF9+F1jC4N3tz4KREuoFQ5An5Zw
mXL3LLZd51zWs7N4jYCgVkt1Rf/3IOEjMwVHHgAVoakOjGDTb1dhMdKKjP6kS6nK76SqioiCWw2A
AMH2osIXhGWIvF8+o05bDcpvte/MIpdt+XFuQsUX7+PYqCbP7PlfLrXbIpT3q8f8gPyxZzL46qUl
VBwA3erGDMg+XIp8zjUlnzBfm4cM7sF+Xta14vqHtD1j4/Q+A4hi/B0oWt9J64lS/+vbRrh2LtKm
65t2AxuUIRjZP/D9SGcs+V/Je3uM3SyTfjip5TgTRo4sh5j3HVcCgTK/NvrVItDa0cnpCtvAYLSe
pmr7LmYHJSi5T9YirgUUbbhHEflUBTxmM4bukR8VwJiFNKlIlhmhpZz6G7czeBl1ciBBSjo+JUoG
W8IFwZfyRFv+G4HUfELGHg7C0Pyv/zcspanZ5N1lzXJeILnKe43AfnaNgzxmpRMWpI2Ed4wMuIxX
E4bNvCER7klaBIdrb0JJ3UWB6f+A6zEL6Wu0mHf0HC3BfBow/0UR/Z99tWRGE1HC3a4jcFQw8AgR
ZShXvigSzvDnq+EI8o8Og8Xsav/LmldWGgYA6lnAJ+Kqe/CugWke2PGeMnv6JrXfKUj9osKgRzea
+McmXfZLaU0FwRjBiybB5JUWr1NQl1jAQytGBHPgU+NkK91e2ZYEBOnv6tdaGy/FgSuvfh/ZSMrC
H9UOXm89Dd3qPqsjJfnSUZamXtKXhwt0AbMiC5hvuKN1ZXyZWiDtydVaFvb0X6H27DquM9f8fosd
6ZFyWpKBSFIClZD/kzXidPxZV+SIUEFbYQ0fwHzM5Ne3hjclXTmEaHSuMjXKClGdG9Okrws8O7DO
BwbpXQ7SkWbA36yIOQie3SJwLJG2HF5O955JKQkOGC9v/+NWWRFOE+xRnrNoH8A1IpxwlhIMr8bZ
6gbMthdkBdvvE3oLhV4rHSMK1gRQskknkOoLcx7o/g49uJ/bowCP5I4PGNNtxIfyN6StjQEP8Ohx
ESND4tNJRyY4rdl9w0vAO7IBMElBz8XN4UotqvX/cIqZurNWRQruf6raVSJs/W3UHgCCGOPEWxZr
Qy2Oz4I9JMU0OLnxAZZfzYbMengu8+81J/rc6AQRlq/jgCDRogT7VpXetXCeqdjj+6LDbP03l8JH
1VEMcXAGahI46MhCfhsppwVCzHc659bImd3hcj81syK5U3H/7nkvCOj0ZpQlDMW54l/h5zXaWiKM
HeBFZuvJ+XWzTwe3cL2qeehQnAZXnCKy+WaEf6Vx5A0TFnVIXemwdsG3TiLBVHV9Vf8zYByHmeFk
2nLzF3xt8Im19xgPhTO9vrP3ZXXlp8YtbTKm2bPQ/a3KMcJ1tJytbwot1XDVN0C4iX2QT/KLHq3x
qc0LTzAYB1jgqnBYOuLi8tV13p1fKYuyFLCWmLIu5g2QzExgNwYXNJwdhyIXBxM0tim3fO1zPAut
K88M8l1/4qukC9Rlt8AkKNaRu5D9IBcPMVhSkvY7ZHKm7QyF4292/ojZxaFIZ3oj287XvNKMPwaO
wp7MUyIg5x6DYmjRU/5Un8tmxNF0gUBHtQjiMsQRLnoDXSxGkupADE6ApzLSDq+JGQ8GmXS/VQuG
LC7WGX+PaE3XGZszn5EwVriyWCtEJqRY2P/mwUh3ORu1xtPTFRcoDhCVFF6p0jEF4sPDhjfF/CYu
AcR6MOVaxHGNDw3FcD+3BAErKnmgNeprAm/domWgjMOgMobPKAjQMCI9F3AGqkulWfjUcaQnuBQp
+53A6veRR4VZGC22eWFZKDpv6Q+Hq8oLG297Big01l3PtixwVacUPvQoc0tAuZHl2SiZ75aq7d8M
KW61hhnKnBI5DjPY8CH9hD25d6AtIns3hpsZWl+GnHCSAF3uj5v7G6pPCqCLLSxnTF4lFngG3UXk
SKDcS9LsoRPliTiOBFuW8BAZ/gFl/XKnMdNH3rdhlS4NHIhks3JEDx60IqXwB9BUZ3elETHI2a9n
iWNv1RXNqkaCMQ51zeAfO1w4y14nkwL5N9hwyYLFvbiFlYcoC2fgJMJaHXnVvXwO0X91gaXJF2dY
DTvz8LiGX2kK+LCkbBiWC2QAOdsMUJoHRxBdN+atxUcRJaBIxKHq/8LkoFh65ralEElgfC4VAwpP
XRsz5evJSDArgdrZhhXhSrCkJ6b/bSEr9WS+0k74gHuVOKMYsSG9CXNLUT6ZS6vh8k+rqFoSgfjR
p0xKEbiDpEocHmUIAZ81kRynWOMdXqKI28xDoYPaTpbJcyL3YcT+L8+GyNehLqNym8IPUp8u0Pyk
s57sC5K4NLhh5OL/0IvZxXIe6rWxRuCT5fTu32Ezsq/bxYtJf1BmBvGqRX5Gs18bdcuNLtrSuB6w
0jlAXgS3PyCc2uSYrTk+cCkSOtmgcPAmaULPmonYmJu8DjwJP2b2154x4X2FJe7ItTfOYYX7leEe
ggyeH65qe6cc3ONcIgFJMDNFcop8e3s+2kWkPWuCH36lDH7PMBrM5myAtxM7Pan2ixmLqCG/7Gi1
7fFFX9r8e7VSpbyIByyMpCBQLRvH5rquGWj4FIme5IrthPCDaNQLwM+gnd5D7bnmdmre30DrRxIp
Y3eukZ8J2OI4U4ORje6mUlNicP3gpkrnzLwyFcq4de5j1ngh//bSPVRCS6iRT2npzrRsJJy7uB8K
gVj0SwvYi+XrJaafaMgVoFN3+BqnA5jLuOo4a/Ty5cuNDiskh5yhOzN0cCc3TdelWxJ+l9X3bRpO
o9zoq12OE7AXyEKEa7weTHu/5DYBlggDRUnGYxucN3CdXFYn/9hkj3tbW4DjOWzEB24eMke+p0DI
CKlTAC5NFsJwjuIK3hrQ3rL+y4ugDCJyQ6cnWF2PJkGA/21nl9keUrm+pH/Z0OpfabGYAXuj1yfZ
PscvyA5Up9OLH4Q8s6UNMQjjQFhAnu3j4OMwj8X3OzEq6UHoo6MIs2Db7uLF4q+x6/y0OEJYtT8p
YOVh+6VucEeeea5sbA9XLsJojpiC1r/eRcfERnh0C4B+loHyCUQR69utpOX3pZ7dZUHytqFVWxEB
IuihWVuKs0jm8mqn9JKSzOaEe7q/z7SuWwW7gy5x0dfIhQaKDxONEJW+fus/IMlaOnuBIIH+bTHc
NdUgEjdmQKBlx8UtKPG9DBJYU5KI1ZNQZtb/z3oNxrDVdzmkavvCM/oeE3McL3Z/vV3URs4t6Apv
2b41ngxGMbFbxm6i4esidnZdr4kY+wRAJKhBDl7N+R8iEegLEsP4vFYnT0R1B3T/bEwGeiSplFEM
LNUv4O128l1O4r+1FRkwHxBDuhKDfNHDkrYiGu1fDn6+WMpTQpWiudXBDFgG+SX4pqxMmInUv8iR
ATm5HaROsVVhFvTBL1r1A2PyLXD7ga5zARxe+PJSeN7+STo3M+c/xnsZPrB9smWh9KSt1ORaIuVe
1ssOnORyDtyDVTL0MiF1O3qIAvidTXn1ucGTi17MIA7h4rNyr7Z1Zir7cCkalVNWTnYZIyeO6xsv
U+3qKt4syU6PwISq2BumVVjo96d0aX+2nb7ie1BUwBASV7gIJOMq2DXhN/azL/XyZU/Mcd0ZLUdg
EEQB654lt9pXLi80vmwHbCXBiiPefOJjUX8QhHrID4N+xRZwDD4kdfiG+3UKV9Wpv6AH42IOmD6L
CCq0y4quNBQh4+BGguKMqip1UQHdwuGpfusJghVlKSyS/77HP+NwSj1s5TVToeGi/btkWzUOuVe0
CKAv1G5ubtZPYmH6l7M+gWiFqs7V6oQ7a6dFntSm2OTYWzefSGlxSDt0Oq7ojEOQcauYCkqWlzid
ACBHODhal/lXf7OHX6KOw64I6i8PshYQfHZS9dPPc7LfdHaTh5kbj8fK5+iJxBTH0yFw74d8Cfnc
LyDtQuNF5Ph8syOUN/MUHCvXxh9qsFsuCxUbPIgzbs85ubohg87gJoz7EnUEK5szFLjVPaVMTdgK
RYzGkwk/8oaqFaV77d31slKX6hStDGLUS4qMcUSmGnXAwHWQaRrzj+dY2f+HZnkweOybx2KF8j4R
p9Wv3p7gmDrpuluQmFRQav9cO3lqpD8RwNTmJ4nfEsTQ7ib3NEcGIIrgCbDzthrmdjnb8a32+2OT
OzsaiiWYaaXsBNFT8rbNRTAi/PdE0qniPHgWZ+W3nebupMZOgjcgMp8W3ms1/UBOwaX5AdC4kPtw
fopKxKmFun83XLoHG63yYf+hUySZtfmwkQM6fJiZ3UaTT5Zls/5eg5pulB9SJUd+ql66UBCylDTl
JdjJtS8ROYlCYUCWXSWVomscYmBa3M9ecbJHR3QhdTzkN883fTW/vM2PABW13MjRK5oT+wtW+dc6
WfAWbqiY86w3a/F1SyCSTd7JZdM2pDojSPseoh+wek78QIc/8z7eYlLkHGGVyvdAOpxk9JSM1Vi5
Fa7glr16sOJKIJ8BNxU7pqMSbNUadQfS/RSfGZjrMfXNMeiWacvZ81eonQgrTMk70EOiVXbYP6mO
oLvNwNDdwgfLezD84FHJs076glHSx5Y+B7c0DdDKvEzGpAxgrv5V8m06jcOiSTGTtc2j4dDw/zQW
DyUTsEO3zdQQ5IiwLNxnM+rAoplH+/sjwQFVLDOZZUuSEhYiSgX0nulXSU246+pjgTjYrcicgbrp
LoSR0fpv5OYZMDZHRLin6/L0RZ2nJf57yvE7vTjyHVBEbjjdaQMU9TDrHMLQD6z9w2kLAq2R/JCb
Zk4tIBn3iOEP2jhml0jqXbnY3BNkiOVIVd23BA9JhS3S4nuntspnLG2o5Fg5qI6H9gEXjlofe7C+
rAn1OkzyRWf4SEfsiL9vE0TCskmreuJopK4EItBMfPXZ98RcyZgGf4UTSoRUqE4z0TquPq+RgwlZ
L01436yTRQn4qFVp1P/4ti1eCU2UyW2WNW4gn9GVZp8bzM5rhvhlQNuQ3CDttaC4osUaVLLdBist
kpkqMQORYdhAnKVHyPVl3PS4ZtyQgvd1xbaDuC3YUl0Q2OoFloXfzViVHVIwwUiDC/3Rdy0HgKPN
C/l9S3hH0rLo1Su19LgqkrHz56psJ7V87qlz7GF+24FvG5RcvHL2kq/jhWAi2ToqP8FTSP+jCV7T
mcLUEeI3wH5Sz37/OrgaVI8GsYQ27hhKBAdMujQbJF0AuUQ3B0YDdrWUGJnJf2+wVRTaVwuNInwD
oIlL3kVqTwAJyJZRMVWg55hUoN7cXe5PaBqyt+Qimct0Uc3EL4z07P4ovilCiKAUVhXCMup/kpyd
m4NElRH9qGa0kfdgaOL8l5pBZflDoP/oveIAfPHTit7CqQzT0RgCYzZjjq/eEEogpKi8oN0nO/6z
j9z+XLGWPs1hflCtSz5IgRZSnv6q7nx2laXZG/GyqwQ94LibuBJJaK4nW7Efh6EbGYEaZnkm+RXx
Ykgt82KuIMv72nP58koONJRhNVGyzbOPIuvIcbnfQvJUfq3OBjIsblh8ENvfk0km7R/N7NIcRuwN
N96phG6LVvUS8drVcOIdZYwBgKLrFq3f0Ot7IMh5Zetst0PxFMxOeWfyOqiWGUaGEc0MPZo2Ux50
Yw2ZcqUIO9YUOjkpGJ9vOpgBgWTqu9Su9wABWfFmrUNm7j5cX2PxvFXWUtgYh2kYsI4XpO6D2l80
9g0vSxapD9uevYPBCt5XyyOVC5WX6e+FxADON5RobiToGfgKz9AgoQSWgfkvKTfcuXQFDxo6704P
3hZBl31xOBWJawfryPpPrP2zn3qKkMu28jOcqDf4ad6Jr7TABI9Figjy2CuTI0Zp0ssdSK5lzyT4
wngyLE5eWZ5enSGGXI4rqeMOrs45MwrD7Py11boS6JEf9uBKtV42b3e/O5Irl5g4wiDqJm6u5QqD
3UFCgg4t6AtNG5ppPtj/vBxndWFuG5kIzcRNQeCIzg9ASj2Didnj31oNf5tx6DuFO5vgLmuN9Z+z
jhZFSbtfPBA7zosnmt9nt1HWWjPwemQDfR/znFoIRjq8CA+P/ZFAxOovpas8qbdwij/pgsC7XFo0
mUSnXaaC431pVrTzMCedNi1AyVQnk+Vuq2BVuZnnN0Ubw7oUcu2AXuDr05jzi4cbuqxyEMkWF6HD
MDj2t2bRvLiIN99PRuA70nSfvftySmYbgwrBUSJvsqXqjNHoIbcvZpsepC7jvrEvqhY2CRgRk3zA
0vqkGmBPiq4hEdxXgz6VAVt79KkYLTXij/CwENkXSQuXPHgJITsQ/ETPzxMkSe811bX6mIy4B2oy
p/tOdLhJrMnGddzIGxygm3I+EHYVQKxTjawBuXWDzdl4G0kA78orZR6MP4Q6UDgWCdSkuXLWnxII
on8cWOft+ec5yJ1/562XqVVlNgMREZg9pbhz+ZIKP7nzcReZzHCQJfL/eiKoJoMY5eQNKcv7v7gH
sukSuE+BAU0D8A2u2gmtmOOIrm72g52UjahWbQHh9HDPvWFDE/4eUz+C9p7L2oVbtRw1WcIvU6a6
+gWWmM8nmvg2TLHxk2tsgHqBUcMkbZPfDnAdRqzqHSEGNvt4LAFoYI+jqqnxtLwamvTHjwhZFkWq
DYulkfw3JT30XIo8iTioPUs//NgpCDsoZWVo/qb8BkUQzDoqFsdDFi64CavjqWoMLActJ72mvBz2
xMsyd2HL5xX12c1iP+L210WnA7hllLTUFlGsb3R8eWs1B54C0hrKq+YGuwcUtf6x0SZcsQVUlRj7
oRag5ex7dK7b/qci5tSnrI0LyAsqr2pfftPGc3ZfKYbEzFjM+kexEp9FZo+B2hg49nN2eir81bB/
XqeviG+hGA0h/TN757s/t7ThFnEQ0p7KbiavCQIeLpZocc91ASxoh9YyJN+4FQofLyEeJXI3qrPO
oO3BIkLNIvJRbU+mwhLyvZ3JdMC28ic6DrKVDgXAEtDbBKwSdAaqKGd0/KCSGGfX3EUQitWQN39f
K3U4bhozNkCZ+xmcEu9dABumNyVr6oFSSDnlDvXF+5rTs1Z3oaQfClDUy2IFJMDxtJLxpS1Pit2y
kfXjEqerhTOR96bDHI8wUN0bQPf0y53Vcrv0iPYNb6L19zkeFG42g4uwZKqbuySyPhQ7sOH2mu2l
KAW6jnyogxTvmz04FlldUUpWmnrHPjyOxYa6cQyvdJH7Eh/vLOArUrOEu5BS4b425lp1K3M++Kes
+wJ+7IBMbYAXK6RVMYuSFKLGABdDbdjaJLl/FtR9uIWp6zPkVRvG5lIfms98HiwHRcTHzkGrtGlX
9peQdqP4n7wMVB0jEIhinyEjpV5hpRc9eH/7ZR7St5fCU8JX4ARYTupVfxNPXPhSfPEsx6j63uKj
knE//AKE0TV9zW7/0EfHe4MAPGB0i2LGAFwObOR0VgZ6fdXKkFKvHqxYpcpYjiUoKMN6AvFtEoDl
LEnw+cq9wloyd9+g9c/lRbFrZIRgDng0kgcUdeTBLaeizI87lwnKpBJrqnvI6Bz2LKvidin+EwN+
cNgIGmd0TaIR9luZ9Pfk1PIS2MrJjqHHhhKywDS5YAJtIUDFzHBCPH0i1RwgKVcWa2J4OFG8PTlK
sJ/VbvbdDhSP63YMXvyRu2g50keqGhjpFTwE1RE7Q2aZuQcmAl9EuAEJOck/FZfOD14vPZEvYVCP
XlDmWJRdAUJjVN0kw3nJ2Yk04bLmItBndOdR62LNqj/hkRLd09obLBWLHytCGp7giGKizZfDY2ko
eLdJ2Il/ZgcbbcUL+WqV8JQ+QdFLhA7pu2zG58K1dRE0oSIu5zpGRWbGyfQ1/dOC+N3vbRYb/yz4
BS0n0rFdlhUyH/OH/uqr9Mq9RGE/d0eA0xmunNESXeiiJLMWsCp7cXhGeGcIniGZQu1EuZuXq0ws
++G6Zon46TnIogSdTSd3dLJcZMVbty+nL8NHSaTYpJjFYEsnlEaIPiY9m94nK5+SBfU8TM4wAbxX
dokwNZ65eggyck6zRKr3+F2e44wofnh7p0bak90kd+Vgypkm2K0bhkpAlp2rqsooayBmHQuyPTWG
PuHzsnha6E9cR7Ji7I89a2UYVqRQnSvjlDk3JMg+a10AaCOdpCWCl3ZnBIo5G9cbWHdC2NAG66s5
0zJckahzaQ0z2wKycBhKPAG5jWHVe+Rnrg2daJQTIK7oGzExmHHEP2+cHXlE5q4k2beq/YoEMWDQ
7fGreRRgG0eh7hd4aWiTAIcIORn0G69dxvB4gv74aWTEJK2p8MPq4Kg/Hbgw9+fS/CRuQP/oaj2b
1fkTlVlgASkViGuGtLd2xlhF/4+Oiz7fPVBmWnU6It7WD/fxxvVc5fcpvI7JlgXhvNK8/Xi4CJ6a
+4nm/Z1AvodfKrbYcbrd9qsf6KppMNqjiwwPyCg5a3DyyN95Wl7cUs7SjgkUULhG8nB1vZ+ChJBr
1CqIY7J4nLr9qurM7BEmYolnhACOgCZEn+jfEvstka8XKvRdFYdrtkw41DwoU9SPaxNhXPKc9FKj
UdxPGJe69yfu3T9a6vuEe8VnZ59V5abJa5tdhjCIh1POBsJ97S7/WLBXOD/r7Sv7G0YSXKMwGNQl
kypEKAKRJVVLUV231vtfU24qey7dMi1oM7qRd8PgxZ8lrAyOXeDlXVnm8bgkZRirrXoFpsg6CMbA
z7nbt3yr1cUYZiDCAaicLzfx75uHiVWVucCMJChEp4vogY0kV1q3slKhGhJWRkFT9dtXbffK7mF/
PS9ZSLXnKz+k0FQfD0vvDWWNBHAPocGF9mDghJpYTdh5AS5dwCRqiRH67mqfyjn3Giwu6FBa2bBJ
JrPRfGAU2ViAofAW01vst3ZA/GjTzKQ4gg2vkYyIsIaFj/O1+SSYC+cH+2cgU3u+pvFS5KVKMqdr
Ht/Di4LQla5vKvLobAvI5psFZPske4+guEKDETHThkHHHY/rfGdcUFmwuylmswiFsRKEVadxLhfo
eGS/2T9HrHOGuTojZoXSlkKN2PCeiiuWwcUvWF+1xDz70+lDSq14SW34wkK1JNYYdspxXrgqxt5s
xWXc020BaBdhG2sXgABdCsV0mFTX2q26QB3TuZ/nHuJWyeI56mFVvZvq18lC84GUkp8oOh0o3nMt
9KGoHpp0YRyRfYDwwx5o0Ex+peJzh3OrX7D8ySqjB7XhNWNCm7tqGNxPT7QQY5E5Pclemt/hPdBH
K67JwwdmtKpJu1q5K9dSdqaGen29L1Vh9DCRyNsUThz18L/jdKFX4rSiwIkHkMsVNuYH86UybYir
Pfzoe4A1c0geZ0SnFQkzaBobT910r+69nyauxybFkNwLGdOloYl/intw3kc2xb4VA+vO2Y+SypSE
E5m3iEvEk8aL9b5dQmUKtMCgwYCYmqYW7h+5jIvx6uMs/7d+LwziBhf5PnMW+0sHxWlSVhnf2Fji
UI6y80xw5dr8o2+42WBiZxeivCP+WHwdA3PjDpkrOCk0HO+4YCPXWENek5CXcv6yzm1nw4uYQAlA
60Ok8yOnyA6W11c8E2hj4G1/IyhaHXrZKZe0qBZsn96aJ8inpCDzxxhbMH1miAUnbicveQaEZmOF
byho+Ak2PnQw0zUU6X1TK7IL3IZS8psggdW39B30gkl2kvOB2+I+f299B5YdEADC6aWKdfp5hUQ8
3bUuVzLKrzHvVQFojTtriHZJleK2uLre9IRGZX0GAy2b42HaUNWKBVpDCHEIxhhavRIO69I3WAHU
FlqS/nHAmIdso3Pquipo2lPKGx9ihTU6eR8L3hloyuDUEDRzkoZOjx4h8DYezc3ivOYGR9nZErSM
RVn0twe914X8f4vQKHr7R27y6FRYRzsQmMOrzBYNN9whtWXsstALwldaGaa0GmEba9MMR96psztF
FWLZ5u+kNJKAWlRpBX8p35wtMzswFU0Vw7/z8RzyjM6H5o6P3pwRFgVbuF+r1Rua5lbNzk77hhI6
sFRjZjlYv5xhpAQ2kSbPM4DuhdMyQTR3W0YGeQ5f2iT6+jumHTLsu7sn1st9WcDlM53awNoUpbSI
tGSrhI8n6w9LWCW7xBfE8u+PJxuoVTMkIZ+OYEsCJbOzzvtshjzECG66ROZw/bmS4iIvzmO4+f5D
W0Hy9CgKReE3wAHi0zUKhRo/jPKA5T5njE9PqJKjSa0sUC2CW9+mWRt07eBsxS6Y06QOl52Oo+id
W1txNolUkXLjHOuabV3e1Gm5P0j+Cx0dfUpET8jkUAxOYErjB9LUgTGZyud9nHFhOKOOWfFMep1b
Vih5fpSNW4F12OvItLWbkWhkTbzECrbin6fOKOPualLuXlsgawoOHa4aaGLXSTbg4C48gNdh4Jre
u6QQqB3gHy8o+UY3Xy2cx5aLuH/BGhIyhdkP+g6UI+9gp7l2sFvFlyLv7IRHn+XRjU4cLv4ZBrVi
bCkE2HUhtBq90ofrTNsrexXrS7LFsReUuYBpZMbzEXW6G1cv1ujYcWhyPwjo+xkB7Y9XDyjDIEVp
wtDlbaHU32F/zgTV+/Q4iHelb7GtYZYs04zXsw0hsstKPEgwSbciRNpoue0Qp9/eO9a5QJkB0PLb
zKhhbZP0Tc30zmsUjzqpErQqkuuPjO0X/woUJSsh8O9ahZjHiljB0Zr/qdq7At3En3EzaO4pQ2bv
dzy48Ft67j6YaNV7dbVJx8XjuzKpub0Sipd5UVDeqBFHrflWqg2DPJY7BAxkKhO3//rnxQZwOUX8
OwtI8LlyqQCk+zl35WzMjH66rm2hB7VrZgzFSlXHipb0Gh3bisOAQJdgG5izc50CSdxN7a6WbBxK
x7tGcGTfbaiFZ7ARPkBg/qlUfywXCR3Mqp63rthu21k4C9vHh84+0gp+owiNKtKKfEB3JRxM/Pj4
wVaUYtXIbAFSkj+CEZ7HvTGM9J8o2JgDYhU/vwC6KUjKTSKa5wtPdFyrh+5LLGb3kiFKPJOr1yyU
vjkVuF7CP0hC3tQIk/pVXvlsPjZkp9k+/DhydAlDtQOCmMSQozosjESTlf5+s1tTqhuCJBMHrv22
ff1ysmkjfean2xT1bcMX/xOYLX5a4sI+NaZWrVrLcrA9feJeZgDv5G4aAfkOGHk5l93dGiWh0G/j
nBP2nar8ntU/621sUUheb/6/vC2RQW7FYSPOeErDt4FfiKUaCjpFOPoMNf7RUx0ggE2wHlXjkhE0
DhZpEZXdJIQo0PJhRJB9fCnBmLO+nJAVHZtvATNVDv0LDD0dFhGeUF84U7XYWxwLCzFGGHvf5qkK
p0fUnhHAZOjaBRmV7PTa++kbsuLCkibG1e6H3ciGSzwZKELDoQam6vuCYdPtLu2LW+Wi4dv7FobR
J+TurtSFZYbQzm5bfuigf3W3A+Z3j1JM+jn+iE2w0sQ4AG+Lwzn4ISmW796mbqe0NbLLjOzMnYT+
+/kosHMKizko7AKAELkEjtaQGGuIrSGugZCeQliPU5V1hxkpE+wUfTDHyksw2k/kIaImjTHPS01+
naY4RY57F/k7mxvaP6RgG/pxVcLFn78/Xk3VT/+ig7++CYtSAZIUNVzdod/xTqypMpQSADxQcnER
u3oY1NI/8DGMRphsE+JocsfREYEDFCkSNlbA8kBKmRS0lyI7F8IZYH3U/K3CLS9XV6UG5h0JDtbD
W6jdq9IGcuAAlHP1enTBZtoAmbDef04OwEI6OV782Nn8NWSzViKYE/HZHJonSEz5vjOceejH16qT
ZCmrQYyiZC3XNdB/Wc2RbQ0ODp701+J6/G1/cFIYWb9f2otbop9Q5HpWATHV0X8TINI4yJisF69J
R5A2vvmg6IObsVY6ltxKEDDiCoOU2CIxM3G4AxZpgNcOhT0K9ip0AFWdE/gQa7p8yDWmQmjjMeZ8
g34CbZJemn05S7c+2Glsvz6p0sKeoMgDkI5ViGdlI0XnPxjtoxm/O86zZUixbIrzzzevOwiYP9jg
r2nJEJBev+ghXWKEI8fsbisg4c/g8uVoaWhB7Cf5fPdRK4FAmCBxTf2W+BrFpkdVYt6UjzN4LQKh
9ePVu3KFJzf9tspbjycl/7W24RFt1LN2ghkW9RFJrKavIObEtDIz8rcZXtUiD7tAPbaFkKa61UdE
Hq026ufyTfLjblIFDKdxL2t0zxsukVfSBS9QWJTCMVyWZ/IQVHABWc1LNr8QfvVkWxwkNPdjB1m2
FG47ASV3LPoaGa9TGUoKOikU/1rlW4d1cfGWhhmlfPCsT5skhu22WXcU+uE6AwR+53OnECwR0gey
iWUmJSZl6u54OegZdFbXCZifV65cE9qfuYWrDwEXC58To/rvB16EEDxsZAkSTWXrejnmLFBebzkd
UDiWTSJqC3BxThBDo4Gg7qSXKmVM6ElYLjZjpHVeJHC/GtWtybZAUOWQB6+q1Uhtg6pbeARzDHWg
eXMWLMVtpZULwoEwZEQ3REOBXaeRXOWOoCs0Rla0+YHc+C3qYxgB2boZKzlUFy1IhGDIZxk1av+1
twMow7q6feusetRQajAfQ7kSNIXxP1DdCS0W/q8xZP4HDE0y5lNMHvDhwQ4zzvFfCuD7fN4fXtJ5
9aG9t7nGMoRtWmqqQk+9IoQg18+VtkElLV/8WOr1YANSFHm2wrl/qZzjep439NKdEN8tWkqZOwmq
BeD/CYl9YAH69ekEtBF/+hqpNHjuKNL3/VZoSqhzgVx4S9Zuob2wzIj7I79qDLBjVXBCngkgr25U
opKS/BmAeTQJFbqNxRnyO4Xmw/ruCcsV5gfhOKieTPEVXp6Fgh0PRYIQo+flathMpFO/8eHrSd3W
NejcYvpRgQ12vESZrFLBEI2B9NMhPn6F8Spz6+2+P7X1NxnwTO29K7irPFJ1sxvbo2WkCkMZvziZ
3R74veaBHikxjbeCD2lF6UBgYWe8o+SNdyM7Xa8z/aLzIN5jHzLNPf/+3+kn6cjmmZJ/Ex3KytzU
IBSWyHkzCxfSdzA4Em1xTva8w2HD+pKSbil6OGyYBDI9LA4E1YJSt+N0LuId+xUg5DoIPZDC2EFL
BRmz+LLGXlXhMjkflYaXcQmXEUhZojRKRSIiYuJt7pWDaP1Zs15GZU1glytxwAqABbIjgPOAu7II
sAc69Bs0hUgkwaNsETta6msCl7O9ja7fwOT8pnB5qNF1h/DrZtSFOTER7HL5S8MUExRVDjaqfr5T
YFep/wDOZy2njgrEuJVbVYzCU9VOzDRFhDUl7D0d5v09SLIRA48RgNeBsqQrvuLnAOMr6fxlcC/l
GzDlTykApWFB1QZBTVFa2uPZZk5VP4+WvEc1Vth+u39Cu54T3vP9Ju/3wQ9eZDcyVRxob6Ng/7cD
8IlliB9j0PwYwaZO65SNRg3halABjVFX8/+Nijuhb8OCxeosI0XuZLcCui+22S69yxuEK2CTYPO4
GYs8Fwi9qmX7KCJfvcg8LpGoX9igJOyFUT0RvxS8vWnt6RTnAk1nqJr95iQBcq1UEIjFkN0kpYmi
LL/EUmg++cMeXPAljwg2GkJMCpM7/zGFhjNCdDxGbybGu6sLOxzMD70DNPP2cZl6gn7hzp710vI6
D5eRHo8fvcVMgKDyFfe9G1Z3c7+pq3QCG44iQ8Bc1A0kvcriILOB7IhHNe4+Htbl5bxSAncOEsQ9
g1QOMXo0LS68yLjwEkk91Sbe5KtEg3+/4GeZsLbyRQzZShckhKI3mJrciQiA9kOhdHdjxUE2kwQB
qRRSFyBGFh35PUgTTMMzm4KfUlpjVqCw4InBezCiIf97OjASOHM37vCOhPm2WSfDrbIHD2gGjjwq
TuyycjbjstHqt5QD2HxblRe4HG3eqSNb0b5jr+3rdkqp2e07IDm725oCuA/dm1ZNcyPGvv2l0Wwy
VI2+Uz3Gslnv7mIRgUSIEZ0TIj8CV/A0/dfPScE03l4Yb0ARja4Hss4lcu7UmBZTlYD80i0cZmff
JMMNPiB/fGtFGlt0E06Bkbk0pTOKW6zbClgTDeW/nAsCrtx+ETdW8V73LsL0FvcynL6sbHHvrmpS
9y13fuSQitN3b6duRb31qYVYwZf0a4Xl4tYnms9V83W0XkGmcMRESo3+6B9K+JZ3Z2ZyN8DKGamK
CTFVA0FJ+cjYaH9IjbGuoSe1uUGlZOTXwV9sWAt80oN2v3n5yLLD5mlfZ5fqlrATHjyB4C9theo4
tkrlnccMQfsHXL3ybaESra0R6f6GHuQfyT97Uh6IRVFW7+WVzMPfXFNWoT5ZYIT9LE0ixgA2Xat6
VPeDrf/Pz2JnSriu42wDGI+diC3AYpiiZnCE3D2RoPvdjOYls8M3Rqqb3zu1gZtXlqDUeb+YxgpI
oFXsOEMZ0h/2d1StKxHxHKF6M1GQLRkptZpqgwq8yeI4XT3Z5E66w1ki9bVsRCVovjNjG1FBwJxg
7JbQ68jxkCrFSivQv7NWDYKAM/gwP3KOfY7KBIxn8wtBTSgTdz3mCmz5lyFVnbfmn/aDuVNEoqtA
FKMOcefjlMtv+WVdVUJc+ejtAMZJRYWet/Sh2JCd5t60E9VAEFFs/tW8NM+7iOphrZg92VjhlSdk
2+4yVL8nzDo5myfBvY2vt5uz5VHHEAkKRozkbHRGHUGsib84mARyU/9LDTjDaT4PQ449LQACWRqM
sTnmKPzjWq8/BHaVZgS7iozp/T2GhU0gby47or9lYVgsHnUN/0JCRNmmqsVbaPruZTT0qjbRTL8a
g3+dKwe9DdAyqEj/vw/5SH6rqtBMoGg7h0hzNvII9qy1qzPRaFMctlbyGW/HcSNQSQCbnXxIuHUJ
yvIdJ1QSFmzNiZkYWljtrtNwo9UZ4LYYI9CbWTrZoGTsdpAi53KJx3xDf5r3oky3yx3kauEmeDyF
NTd17Fxl7iz1PGSkt86OR2arLBPCxMm8PnrK3Vu2DucWA56FLCV3SOpeKY9df47J+CFxRm4i/mTq
L3RoeMMfHxKgFMSpSK6ja2cdFDzGNi7TCLks3MFqXB8Pta7Sqb4TXoRwOMxNJ2JboJPu6Jx0oAYd
BuJmMLViqx5qeL2UWPbPoI73dzTpJ7TFJTVyFDlVWrhWrw4J2Klzx/n5TGI+yFTX+xeBg7ps4NlZ
nfSxgVXJwgbi2VvOMT4c6tDOl4JmIHPQdnxgUzmVw9DrrnanGt4ypsJzwjyaAUEADnv8Di25DLb6
7wI3XK+a4ai/XUJ+z1Mrd17HtDuZiAdng/pFbCinDfNWhNgD6oJRtCxnwo5AIFAE06kAkNECR1eK
tmSZqkqjOGzzNn3kw2ed4oW3a88UYfwOQZa0hbI1gwNbmHjc8SKvVp2jB/44/I4x8/vHzHY27t6u
avuNWjCvYcJB/hD06nUToJIlQ9NFw2erqcqSmxuNuKmYPo8TUO3+hZO+ml8agzGHFI5uE9BB9TFu
YSfmg7UonV8Inb8OjWUl/+HFZnMUBvWJyDOosih0qG2vI4tmpyOmEyBelNboDR20rVyQPSuwP3IB
/RHex+/XcQKTYCVNts0Oc/uMK22Yhz0v9GpM69fOVcCeB6Em7hVPgi1ePcgIr+9vym6T8WcrsGzX
2qJ4R5oLmzzVAytm4W6dHNEMvUmZFhOL9KNNSgaOIJxe1cj0pLL19dvfKTvx9hKelG5fuoWEdMjY
ro+Oavd8dWSBnB+Mn0AvXnMcjqaVIA1dUe5rYc0evGUTwTOq4OtkjT7fa0Ryeaq/2WOlQfvVhvsU
RZw6hRCMzJR8E/RzXmDkgcybsZZqRnYbZCxCO3zP4rhfeAR0rXQlRUDW8sMc4k+hHiObyJA7syYw
unzBjU0pNHYXyFsmAN7V1t7DVzQpIWQ8sST0Aq4FdLGMDQw+hc3YQF9w9YEkOkV3CRRxIwcLJj81
bXSsYuICWTncQQlecWdqBO26uSNr339IC3gKMeOXio8Pnt+9xq5PbId7t2zu4gWVWA1hMxaCTh+H
qZERITl3l5ZORoTWuvwsO7Z4ePuQGNV5NwETy7Lfr9SKlXpo0IFVZNdbqnyFbWCD+IVGTXJ7iPne
NegSGiY0cxE4axi/iXRRZgRw87ACFdDttIi6aX+BJgBlo0jH/G97rSc61CO/mZ3EEIdwEnR6qEAw
Bd8YlsLqoRAlo+Xkc40D8GogJ/aST6itJhxIDnDqMhdt/exTt4vwgKPPZPz4BQP8dfTuL+hFouW0
ee+k8KtUthJbKlhtlDa1ki2i3BMwdsx5LXR5xxHK/VAOw8DgSs9L6aNlCEL9Uo599z5xBZguFQLQ
Rv/dj5NRfM1Pdj8nFEonMDB1R6Fll+Nf4BaDFht7o1Vs3vYLvBXfMfoS4Q/va5WPQa/bDqlUJlOF
L0RksN82+inQmEu0ciug/OQTtv6npg9bh5SpGDKxlNiwuxnx3Drlq3/pxYXCpbDFq+FVxXfdkZgR
pOnRq0GpAR4IAv4fl0PAA2Mr57tUotthFLszY/9iDlKvSXZ4oATDETwODZlPspNJfNjmINqLRFmK
nNuoE6LkY6LeOg8XZXv4En9o7nRKj+4PDkw9A+H9vYHkZWwbVRtz4Q+AeWjk8tUGfob8Hex8m3OD
dFnWfHur69DhlZlE/a8QmfBcvNwz6bEsmmdOKsuU3ezAb6x1VhkFulNDMbxcRjzkKF7XpVtdh2/N
Pkr2GuwNhoXGUZmQ8Z7pKa8aTn8mtGlQY+8HSof94bTzlVsRfWVm1GCIjOuBBfe24kzr1+D10sRD
obgqvHGOJk0gKh6vYodct7yX54W/F7jiXH8rRP43v8PBXEYSiI9MXajolmoax+RamPhHH2wd8l0P
MOIMepk+Bk5WCqBamfybOxTAB4sGSZ6NAc7lbE3fqoOEmfigu7s/lrNfPwj36/12L+StSoXc9/6e
XRB8DUUYJPt3fAeYSL7wnfEdEhqHXRsv3gCZJ+eBs61giSp0RATyENQErJHEU01i4iWbZ/SW9hn4
AAOenIW/zG+pr+PqzmJ8/0qt7hMkfO/pKE5D1BnJwO52mcxhP0CIRkk+IHS8HmgR8S130o3/dGOe
kF3qdifUYdRoyxmnCUF+XGdy87VuWaEaL5IPDqjqRi5aoM3dKmklDJBMaPGgvZQ2+g4RHsFCxhbe
G02JCX9w4rxHqAbCjE5MTAI5rEwtDcc/4/jw6NZ9ySQi8Ss5wFgaTQ/Gpnx54n0JWUo2+CWQlOU8
2zDLq1+9X12fWtsUDfsBMR+CyUrP6ObkLQjwvGTpiAr0K0YlWyhdCSP5uKlVdudaotALQvudkBH8
ZvXTDa7RIi0S2QycOP8gttP1SH7tQTQOnCfGn9IpWFfDz28QlSp2QfyvSUwnDpdYISFH2ddaFSAs
LaEf4YaUauLo+FxdfLUMoBcgRjxrXihoy4pQznaup2jfKycga5/uYUHyk1XKq3dBDoxL/yy+Y710
XmBFwSyTBQJk4ZPtYiUwkbu/Fzenln2TDbVcUkWG3acyjA6mneT1I22sG4sRlAb0W0QFo+JHl81W
V6uTY4A/faAmjksB7EvyUfuJcO3hoDAdN56XweZv/nQSVVcPZFMT/Zu7M9CCA9iBu7GYj/ro9xph
M7A7eadQVL5b024FX+t+4P0sa58ZQ6xNMChJ7a34Eivt0m1d2SXHgdPxgZhrAzOuibClPxaszSrl
QgGUkloXMk/Be3vwPfrG/h6MPUZomAfzU7v40qUDXaIqnvZ35eMBVK/yXJWyxRRij6/VT+CkwhPu
actRpuqJ2Kd9q7O4W5Ay43h/ek3/1Dd1oEER3/5bXvxXvd3sZnuZvSTx6VTr5W5Q+2JSx92eZeJS
nSrYYBrt8f+j04Y/6NXe8ZR04C+z8+9Ty0BgsOa+20QsvMzFdVzCy9lF6GSLIEqHrOL0Vb0zc3eX
ACPN2qrIkT0zsAQk/Wwot2fZ5YbuXuac6kcslP5aBSWyiSH3wpCUb3nd08k2rnze0LEO8f1vFkH4
Zu6eM4GqBrJjNoOPQhD2EHN0zMKCTicO7eAy8MgV6SWT3x9e8MSdaBtdjCltpZgb2hYaKh9Dx+de
fEBvZD8v1GfxulA3WTfZaFFzAFRqAfHbuexosGCeiaIZCahZoOQG+7Z+qkHCBAbKCD4Zj+OzNw5g
FVgjKejkQ/PTZJQM+UVZHgNzIoKbvo1wC+XvHyAujgW7jPXjo8qSLR99PwWQzVfMYSz/VSVP3zPS
V/pBJS2hlkYh49sqbiWqH6utnbknvkocl7LKIy/zg/pAKrWVQqnb6DiObWSpolxLHp5KOHYChPh+
NEIkCHE6LyACCbRuVwwge9o/Hg7eAKowZS8TPMGG8PbEDtSD/z8NZwAM7oZrv6UA0j8VL9sUr/jB
YQKJtDUaYGvxWHGu3mi1hH0NGUaugayjjilLtRhXJS4aCrltjhhdfHiixaQO9WDxfFeszfKAE2hN
fVZbnCFS0djxj2fUVJBT4qSDG7t0/5Ybg4iVFjHSrxnIHJhpVOVe9pkwMsiyWHnDNzZ7J+ofEx6Z
jZZDW5AjdfLbD122z6kcFQhsDTZOKMg61BrdLqVKB8xT+h0AaQ9U2fS7Tsn+kCBDTlpKrANbtz55
HBIztczqkT3rBkHwHEZ9ufbVrDwDm2jurogtbUSw+c1nt7wpcYvvf7pagWjfA8YISgiekfrSRuts
yWtJeK0622Cidt8+moDwnfUALaENjR9blO/hTtrQ/VDB6IO2wGPwX/keBmqUTdqTRqff1UhIyABY
40gnSRJHf2JTybHFiARI4FhBw95chhoGaKZC/dwojzj0yf0j8hJh9JLtJUdH0tYNvUPuvSNqKW6y
4PP4hN1Vermr+OgSHAGjrsBkvUfUlwVymhLeahIVW7KK4XtDWpjw8+iEPPonaFulWV7jqpoiVW5V
7CmrlvfOLiU9vr31rn7AFcQ9E00D+Zf1UrqJ3+fciigDEYDahi7MG8eBFOQCxJAElcaLyeTjAVC1
PP0HV5WH29ImQnGbdiKLF5xLDhr63PBmEGUDBCIlCp6BpxyGmzvPTOD6yDhGZV7ZYvpWYIP8/ZGd
7I6CeruD4QQMTXIy+57BUbp59uIztjCT7/q/6e3P9u+1x5Hdu6jZ8PgWFPpwFOa4MUcYhFsvETFE
a2Kpe+V68TRuI2Ggr2/LTn0KgjO2H9uRxvfzZWbbulnFcyGKzM6k2hTU38lWRWN9J5q9zuxgLyn7
BgbUYQWk4ODPlRD2EDWj1XYKukNjDcV8hnOUQyw+gRrq4lne6Dig7dZ/d4WZefaqFrCBzDC7PzT0
re5JjullBvDRDR6cHiFXgDDVnSePuwLVOZbsgSpaimNAFlilpqS2Tp1H5Z7nPeceKA7fwSC5AHBf
D3iFVPMzmhmOJbEXwm8QvreIbO0nNeztBFubZ62iodgpIeMnKRFXvInqKNjkjf2QqQ1rE3Hw3eJ7
cUMvweQAY/9aqGJBBqx+EvdVsoGNLTcb9xVFx7w9yxdSIhwo9YOBSj0IyKW3k2/yQxrhFtOr4ESP
GEBjFUWwiANQp/mw8lwv3DKQn8srWNYOe8+JTs6Hky6AapSVuUyZzKIrI49oNOk6A3A7kFGRCza4
ynKJoWmLqpy58uLEO7R41QcHrfxkGKS39q0LoGrcJk+Su5vE5abrdLaJlQh1BW7+IdB/XBuNA8jd
M+eBabSb1YRUWjqs9ck+m5yuYxyps2/twJ37aHXqDMWmZXUwJ13m8zmLlwDq3XlvnYZCV7cmvICr
0xbzQJZhSAIYBXmJB+e+5rMo/AM57heK3qtabLEHY69qUHTZ7iMXYssUocRAqfVb+ILMpRr9e+GD
i8HHG2lZ88CwN6AjasSopon8Vvl/h1hhuT+2ypH3V89Km2ID3vVbGm6d88Tg+Mb+m8cNhC5Uf2QW
tRnmaUXGeMrsZRkvt96nE/+K3KQlWuG3NNbWYXbXpHIbQyCCjnT37mi2Ne0WVBiSAeGLPuAGcWpm
dPalqZbkgow2JUZHbLUem1jM/U+eh388DpQj+so2ncIvmWt+K2rJi/GcDGRWvmlyfLOefABN/XT0
3pRt/9pC71ZDRuFLQin0J8DGRPgqqOvI17Hr44Ms8h1oPbUHbjLtyr1xtzkxAX1G8vEOCsofA6nD
4uu855BgGrXOjrJWM2EmE6BACMSfzuWv20zMyoVPyy9clUDZwgodeY3S2NhaeB9L7AxszQBhT/uN
rACJTUvYs50cqQcmGhcgxqlVJ4rJc/Q6YQszuhKrA7ujrcY3YlXtHWD2cj4P3Du6L9bZpXnzA3u8
UNzBWazMoGd5qqHbvdID/yNN8SfBGO77A/vtdRUdqBB2aMF2X3KCyOJbOqK2CL4o/rtP4wJJB/Co
erQZ6Rzp/dys41XE7By+A5NTCZDKCdbd/smCdtLNu4qwj99u1TeRUSB6QAroYVxnMWPt03ZgTEIy
yTSyUQpOdxXosVbnKLfj9jPKUH9YCzya8agSk2Cu8ukFx1IVEfXbgaNqHiZpy34IFWmAliItcY8s
h65Pb/g9ILfM7orK8ET+Kz9T+TT3W2KDEoEgNMOIN3H6zX/gFAg3+A2gk5W4y7mJilpqKNIHagDT
xlrUCsRBy23gvn6wL2BhNsCtG2+CSLIpJo77tebCG7xMpFe0/GYZlg2276bECiqw8paxrCUqra8p
Ccv1kwfwdIVkU0tA/rLztCvYpoqBUFxIvCgZqjAUo365kXNofjEiTIw7AkQJMkptMQM1PTF/2SyK
miLjkKbyOEutMcZ274Qgv7966aR4gz22xeBYWxfLjtBNhOO0lvdXHXDje2LCfqgBvI2pEyCsKrZR
pu1XjCxNCKWL7SOKzVdZSM07PIyFW0LDh0NgjqcC9yFhWwARTSKRrWB5r2yOJ3u4xH3UWC2+aHZu
9k41+kER9U+tZgsjbwDB1y/Ce1Nl6WnfzhQE95QwHqUhVEmviAhnOLoJOnvPNLGxiuhUoTE0EPgS
0TCmCPBj7Kcqm6ROqFNmiJK+xWqz/oL7kRHYsEh7xnsi0p2R8LVhgubIVb4/gm+TjBaLqUvEYEND
INMmSO6h1S/Rl4zd7I18GI/ocwRIjUvoSbV0jnMh++9xCYyCCHfc+ckHhlzmF6LUTjFR6mAl7foj
+d+IDgxLp0fQFMLORrOBvsFipPM52Dpzo9N8C4rZ7Ev7zHxhZWevYjiyYepzbcyDnYfonwlNRuXd
nP4zrB5qSJcbH0pbxnlXKB8zJGQUhoPQBVMYtIEGj/j1pdjJzW0aBkn+8fTNrmlveVhnexIrYBS9
b75QhYckVxg3mxekcAx0I3f5AfBxcP/eMAdLaqenrLSf4AiRSGykHSC4EyG+59tPmBVLuFeAiXTR
lEdJsGLm2ZQuFtyFtD3xpqiPnxvMMr2ld54BrPsvzmkjhzMpd/RaM0AjnL4VX0OPt5V9a2g8J+Wo
wUglT0mqe3KnezsRffi1562C5gstpc2dnaMmmKcy7lQhqmMIb/Wz09qOZ0yz8phHqdo1z1lFpndC
S99de8omkgqHfDBqL9qXjKnwhtscfE4LFlbVXbvFxHZP4Yqr3pYVZkti09E/BjpocqgzTYhe90Nl
TYyxzKnC0KXoB0dozTaWpmjOSZYWCPOSdw/zoZmIJWj/2LoEruwHI9Mg9dFO/GKHgcCCxSUcsDng
hYiIPn2blMx2QbtaEcMVxDvSyt985+BqyTrFOjp0DyBjxLM7OGXT8bP8cH0s6bZ7Aev8V78Zmw4a
OnbuHkqNPXandjFIphi78CkUy6uSQn+paCaSkt6+Be5OtgG6Z/7D+EjKLRvR2aVyX3fWgSTp9XVG
0mCJ+HMtEyPCUX74BxBCm8vTI7y4nQHwQ3TSlW6848VmYoSVZXiVWjS3x+qzjHXIDJKWSE5Pnijo
jc++FWKWoT7bVeBSN5XuQCFh/tv1JP50ueFcIpsqVp/pUCo2utBLbK396VR8Ue+Zw5ZTG9MUMBpU
5cS8cf6QRQQc4JK6DPK1xzbXE/gpV7xUFIqItwiozqH64kDqqOXVwhpkjwAMg7qDe11OWLJX1cgR
Wyds2KOig2xlqt0WaHx3K+hNDFF/QNi+T+xvaU47Qr2K0Rs8vUcSlIevtpnPdFp5Z9O36DS3VrNZ
S45C98TXHEqoTXyTrunkUoNH2k5dMs196Eg5pDRWMktxuejsIEuweTr7JG37fnyZd/TBLyvWta+Y
ltZgC3X+BvSBj/GgUkxHAQOAtt41ToCfvpLDFQj55wA3MrmQFlQQ19qsAwhxMQJVFLlDPS8ud2PD
0No6r4BHrhjG9f64XT5qM/FBhoP5atjX3Ya87ZqWBxAIeE/ZclEuWwVGCYM1xWRcTy3PvcDPBS4E
4rbuBdNEOz4G3ub39JMbMNtjniyyX68T6DoXXf9NPp+NJ1bZesKGj5pdI41v7hhDJxC6mWZascJi
Lf06m8qCyqs7asic7tRzfqkCe6+udr7n1oxC5uuiUT7xbMSw+ZcrLBa5XTY+8p1zNuqO73vsWm/w
15wrNaMiuSaTdzEXA43XB5N0WdFuUuvGi3LJKRz/Ii8Au3KNb2vAAWabgHFFBO1+DOYc/jyqAOba
c7y9QszjXW4998F9yVuci8P5iMN5yxEH7IBLbujDt95z7vmS//Uomiv8FrQq+yXfN6PncNtGtaSI
nQYHvJXQXsCjyWMIMUB7kn5cV2RB/zeq2q+8UB6QxbcsP/MhqIUY02f7aMJgrLh5HJ1eqX45EdIY
MDXDOlAgzVUJ091rtQF2Q9L8g6KX9jalfpNxF5Td/NyxYNObR4JLTtKydxAE17VjcuMcpQdyole4
gBO2VBANG9RRbhL39Szv6ELjm4WVXdZ6lIu8aHNLVBpLY4LhSYK24zcsdTm9mYkgeWy0tpp8Up83
AYySAV5jA6A0IIiuPwiZg9ccEDMT1gmBgLFwZWDOs5DKdaQPWhSe2kLcOZqOEmSvnWQTuWzxZWKJ
j77WVXaltEyQKKC2gNJ/u5XyNIL1yCHmhVCQsI6w5copXFpREH852aJ3VI+95eB6Fv0zGNnfgJrP
FDGeMOLzbhJrymwXFik30QL7YH6Fi2w8OzTJAU75/7LZV66KGPzaZ5kHMIrMuWGzkcrBjCWbNvuS
MNKTtjS6cIp5KXQ2zEeG3j80T5AUbzfDC4f3JpKpOmDOVDM6lbIQX/MKn4qwO+WYZKTStLzxfNTt
eyEmmyj5zqUMADvZleZ3vXvEB0mCMgtsWArcmN8Lm7b5pD0do/cl3o81oa4eq5m2yuO+P/um29Zl
nxXj0VC9GBCJs1rv7DdfEbzTfE4C0KLAaXvxQ7pVbQz4deGDrmHfWga/1SCWPXFBzZ60JQXbPFmQ
C5CCepAUy3ZWHdBcQgG2z9PnGcro+J/zRAe3zQGaiUhcFP2GdsXwUOy5bsORJ5xlsvkVIzEB9uJV
a5r57/ubDSGXjDwxicnYQGrJCJuKV+pS9MKNnXEKtOM+a+d6ipmRw7V+e+nflMAD46Jp/nOsSHUd
iCMwaQE5ydLlYzCwO8EemiaxqKb0HLjBwC9XtIp3S+Y40N2yLz3DBKPG5xETbPI/JVNWe8l/04xD
FmuQAxoNKpcXj7WQmS+g7RurC55fJbSlyEUDCk6j+ExxQgD5duJRG9ocQ3wWy6ZLpdTDEazj+mBP
c81wanaaILkcK9vcT/4JyE/gBvLeCgLzywqVYdVHKZKjrbBnCfzNsp34UM/5K/FxHKRfzdUB9dEt
flUXmWh7ftCBNGnmLzzJVSaf9G2YqaP+srkpmsx3vK3LN5hYnk41F2K9m6hYPgRWRSVvGW2LNLSa
LDQEQO3LqhcWT2ed3OdaibF5742tLLK8PMeUjtSQbvLatydvoIccSnL0h+ir+4DmSLJB9KqfwJSS
EExiMlgUwnJDSfIvuLQkicLX13COZ2qUI7PBXnktyYWAtqasDxhVsTmY6BjhQZ+YzrEWTlWxPnx8
5lo3ESng5NImpq9ClRgT9fWh55h4f7IR4hVAPdaVGZ7bR9ElyD91/OMBEWHgRPrdFNwcW7bm3pRI
wwUXUo/UC3clYo+YSjQpP/dEkxmssB/RtcOE7dvy/kqUVdVn1ghppoiu2N/lZ20Y0Lga1hmLF8b1
NsRDFpoZ2kvCPW5xqJMS7CadQIFS7VjZ8Ey5OQvsz9Y1Pm3B86clhN8uGRT5XvAOrxKX6WzWtXk2
XevQeZSF2Efdmbl0HErELqHEk2YFyspc9Zq+SIKZOvrNV6uAUAD8yAPlVBSnvaj3Th8gYryX8bGA
6878FQXiRBEMwcIasrJXPA/s2fM6Ukk9NGMY6Dkc0rI9V2Qn5+qie66Iid0yiWXZtXCf6dHGRWAb
Y9kgcnx1/2A1kSZECA0JTsr3b5q/ub9Z+urAoieHQ9oT4yaU229ImrKIInR337mn1eDXe7JnNBr6
+usVHUy0M8d2dw0p4Rz/vYUOAFDemm3HEZPfKehr8olXesy38T1SIbb3SlOU5QPlkOAwTBdhzh+C
GnDwlhti+mQO9qB3om++zmF4z2pX1UHhr+JBhczyvFyoNS6EQTylUlfi+GkyxksY0k+dqzzyrFlX
oR7RL2uOf3yjwIsa0xONchn6UAUdhFsyGAf+YAasTA1FGHJ/sARIRdpENEGRxBD/jmmFZSqXxFoR
qNjy1cwRgmz/Xvkg24h68Kr9NhOaqfVdgPJsb9NvKBqRhxPCHkkRa8wQtnuDtUGLFWg4JefqmqRH
AcpDekY2bU0N5Xu8xfFUSCZoXCs4A5rA1NK0Hu0KtfQ3opyfRik2G7HXLMQTM72RIffV861VAl6d
WRkErrJx/uR0hAiMGqCD617Yvlt/YEdSr4DHmwuTgQkFxgy8AgDbImcRHhujbdxrxKD3CRo/mvzH
dA1c6nvCx7ZK3el8s/3EXNfF2GMV7EMWnyzXKokkyNPNZMISpKo/4khPOZYQGDoRhGK73VQ/Seub
gUmNpU1hg+skKc4hx5iEqps9TS4/kAEREnCCUBPBTzlJ9qAhfYw0CrQLNAx+f9LXLzvh96P/O8wC
5+tQZUU+Uq2Ati+IT6w/bn2bMMS23RgS6ca9hz2L7XbCFhl2OYuvAI7xryTwOXxlJMCZmUEBqZV9
iqL5zUmU18VjqX5lLjZItOXIkoxRRXe8QvHiYBJEWHTvm7levlpZBXQR0RmPHYVIitA8otiZKE8k
IL13IFM0LwCuHtsCudmg3qQArnNQjjmAQCgT9jZi0nSgFSilTlbOAtsGJ5sr2967I075S3Mc+G0q
Taq/9DZ+7ncdaS49mtq1pKeWKyRZNpSRM28S9MMDtXnGe8WwDOfBBg57ZGTfsf1f++OoX7SaGXuW
fBgORlDDAGXktYekW0FlVNgpU6UXqoy/BEqFK71YjoJpFQzx6Hs/rDHtrQ+Jue2WxMLHcTGg9Bm9
0xT4na/4zUzAs/6aIfJIgqPLfXuppWrF40OSZOwTU5A27V9n06MfqmVX/R4UkDNA+ChN7EFt87ur
hTe1VnYCPi4wC9mHnpJG5msUn4Gt3ZytHvhIK+QoVGOApnWvR41IqvzElliR27h83vWdBtACNASH
kzpQ/IpA29RFa3rmFSyC03MprZSQ/uiX8dHnZRDwTDkRsWf5R1WTusvYE21h7xCcXkDplYel1ykA
lZUBciYx3tphwrAY+Diq6+pvH/zeXqABDjitATOUNwgD48mPZv8e6WHcMLB4752Zwou22pChDo3I
z2HLhynd1nOrUWUpQL5yW0aYBkjD113Jlw/sb117qMDMjYPdb6ndMvnAokr7M2+Em+R22o7bmk9w
+R7pM6fXZ9QE79i10lg+xb7z1tfR0MSSLi+kUb/TVTN9cm9kuPyvdrDaAHu7aF5p434/76lYVr3n
qBkkp9v3tj6xbjUlaKRoB+IpVd5s5yaV++4BZXLqfXeAuam5N1m4JSwz9qcIBYiWkdT9QJZEUJhP
KFBPpK7cowzOhTvkF4x37ldCIy2gAB1ouLPUiD36r0uL5qzFQhwfP5Zsw/mJ+ldrZigxRPApkcvO
BY/KeFnzC98eR3kaMcCY8/+PWdANW5zhOH2xG4xu8LLUQWt+c4BOPwjDYtJy+UpICkmSeZsm5sns
A+NlmhIUqrmEITyitnJn6CbH0DbvSG57dxcZ8uvT+dKo4DnFuMFrq9GOAg870bAfPoGTYNXz1hn1
rjcmcPKHclPxfpZCrf+wQODyD7jbF+sweNTAqCxp2nJIi0YX/15pey4kvgcgefJRPrUJJ961CAb0
A5OXy2rcyUkHOd3e0+ob5JjDJsjrDeIkaUBkdQb5mGaPuFA601xP+U3I8BDMzwfpuMKkPs49vSz/
FCyOqlVV4pZa56jO6YV8IcrKTdU7lxUbNF5V/DlkC2V4kidEnRW/Os8GP20lDO5UUeP+SCWdjT3O
5J+ytj0ntnRZi8H2NYqxk05pKg5PxAWjfdEr5f6GAuGSiAPxqoH7vZqVVM8ZCLv+k0KCEAVzEI8i
e12b43DOhBI3xGf786tLxF/0i/JKkC45ibDKtCmq2JUC24HiXxeaPNw/xb9jOZKoLa+4v1DAVgzb
v1Y+h71fRjP7jo553JfdjAiUsq+EoW4inDkRkuHDjn3y/tG3LHwuIM7kWQryMBt65w8GwEK8Dmxt
P3dB4W+w3Qu8Wefdw/GYxShkgU9Qlvd05Ic8YQa5jEyegWUJeiuMdkXB9lIE77QJiVfjI2XIuDoO
u6rXZd3Jn+vbcWlXCzNcGEwsIkctC0gekd4iz8oaa8wTcS0tR6Rd9Tggr5/P7j4sNQukKq5dNOVq
LAUjUAFMK1QLmxS6wb6nRTcxi5fv1l7TQB8J0WpkDh60w8Cz+JWek3GlEKj0VXA7Hv8wg7dd378x
LdbwV98cLB49EwomgnurY5Ilyz1ej08kUAq/qxBwsUmxbt6ruUBJ5hUxwi/dC+XlVlMETgvDoMGH
mkRk15SjPtY12Yz7PBFoZ91w90xK7fxoK2he72D7CSWRfis2dqyJ4JHDfmeLPqhfoGl8MURLoTZ8
KTJcGs+s3t3MdzgkfRe5EQ/y+WYkVBbbc38QlRQNXfX9NREGmn7SfyNBRUJURscM/hALAu10idYl
y2SzFirTewRZ4CWywjrKqBR75wTzpvghwk1Zvi14bHmQb1uShUbiuiZVmrfm3bPGsoFDGIaZGcKv
rSYvBoRrBg5VyZ/Yuck5xqGLnRaD9PC+28dpf3HU8ROS4maJagBvqPmjtfHJPoCHsji9RCt5ecfN
+l//JA0kdDURmVdxs8vUV49GE9XF1vePEuco2tWKjGuW3HMWYvMzhffjm/pG965i4owOQtHXJ6+a
lsFrH+/X2MTBjUIGlsNOJwPKNEtPj5zlomPpZl07iR36Mbrpq5pNQvLF59GRW3XUZTxaI19XdWcw
+t7ucYdt3yLT/1dLq9MZBE0DDj1NQ52bS/Too2+6RuNL/9GRQz0bMJZXZNENpuUQs86Z/JIXrnFi
kVk54mot5qEFtoCegzKhcxbzfpri/EU8Sf56mdYzNp6NzoeionDyU5qfmju0w2tmNKu8Mez5NizU
KIwyuiA7Bhuwl5ThU5iy+foCB1EBDDAtxx9GaC8Sn5xLyy+peXuBqwcddYLUY6Bs0j0efdLfCYOY
ZuiKoGgyvM0czPdfP6zK4PksIoTjmwK0jjB+riK+gvP4hjr0WMtZSYHaCEWF/Q3gt9rs3cO11vnh
s0929XeBOepnZCZYHOwq307WnBztWH1N7Zgkv8qQrm0mMgcJlcKSG8RGNZef5LXA+BV52GtLTvlS
/E3U71u7G6WM5K7ESOVzj2FXlwHCICnXAblegyhAxFtjitx72OX1sEmiwGdhHbvaZa5dqPq3L/Ba
vfbhXPa6x8CGpc+B+NEXaQYVo0gaFdKt1BGmwbJgECK6yPn20lwTysLzIVBD0dFoUgppiIxrhB33
fbIH+fXCNaxWjnNQthzzagJcI5hpzz+Y5FMNphx/Ijflza2zXBJYKCIQfY8nY9wLQx/kVlOMMbcx
2xJ/2vCN0JqoLdJ1k2ejl6Bg8EL1CHze41MHP8LO5QooREQ7nQUnkdwJQiNrJV1n77ZUfXRYmjj2
tUk4bVEDK6jvqeOfZdZHFzm4aWib2JtBz/9RbqR1fK4ODhJZbdEHvtcZ1Uc+lnNu8PSHFM0r6bTA
rzk3mQi1qrbfnfhWdRFhU5XmCX/FEmJy6HVac3b8uRdhDqxutBZ/SXa3z6Y9MZlqs3miRkaBQgw6
yVbHzc2OJtnQN1ho5cPJmR6dW9Y+lcfoyc16fqxjKN/YlI6so2e65YQBQkYWurNrG9QcfA/8op01
gZWBFs7+3goRmn29aY4HuPodNZZhqFosF8SYUxaVsImE5TRbgHAYlSA1kCNm6Xq9BmWt7w3e+I0F
OC9gUGHCAMgllxQ+vkc5Kgy5b1gUYGev14xe7dfdKJ9tEOloxvXqEDyEl6BP9EHTUSerIqvpF5Lw
d7AHp2Kndp/GwKqQz6VFpMoj1rbXtGoaHjiSQEFPi2H0C4GHbSbsI1AqwlbSOS3k0kxGM7hy0KuI
0b3+IOi0s0wug6GSNR92zq+/aXHWRsAekldbdzvBr4EDOMy652/wex30y6eOgp6dvJxb1D55VOfL
Rt3HfSsm4ROxg2/4AAoPYJpOjHOGm2ofawd5kL2XVtkzbqEXOaFAKV1flxUkZdLonOwg5pmYiSMD
FBO2O0fB2Nbi1WvFxwlgiodGJSTg5p58xIPP39nJK4m06SCM7xPw9PUEV1OXU5UrvHXSBHjRDMtL
LceG1P7YTiFz6/suBQnZBN4k/rRvrOa8T7hgvjtV3NkEZC2xQmFTGZL5Aq2Ku7OIATLRC+Rh9fEt
TYHOp5NhP/Og6ky4xa6FNRtxqgjmjRnoQ4hnTR/3fVdnDf9qVbRUh0Vr1A9lliSRxTnH/DW4red9
cG6kYju0sMjgpww88SOPO+iVknFjtB1CF6lbcb3F/oTR+ym3aHvyUucargEhQ2rUSxJ45ZSeN4AT
VNwmBwZPdZI1Wx9ywoSVNOcRPZYd+x+cj8ICAPZ9yFel3DYe6VcrWgw15P67jWg9ra8uf6Rs3k01
GxMt9dt/NPkFxznQ9kDHDVnhouXRVNz1Po7Y3evCh6551TPX9h3htswcpNJC9x7jk5KO4x7XGa2P
mtfvHiMw/CT+fqVsWbNxpJJNmna63LoZPRi3ODZfU1e537mytTN28SOG1E2rR0LmDRZK3D7KnygA
jCPeJrtQ5ycLzUkwNZEzR1J3ZuWwylawbLk/wPoDSsDlpSPC9TIwZmx9dTsDq5V3NttTNPQyet5q
b2vyjs5gEEaeznlhCsgJwjJa1pgNtBPYejJYJNsexchXoh0gNCaxHK534IfeBrMIUd8kHBbofMmq
maoMkX4BmyBQqcFRUSo6H1OOFNLvoT8pLtYe7Prf1xTbV2PiBMUdAPU+xc05WQS/4jAOu6wIMUBh
JOp9lE8Ei5tFUiE12nVOkhkFgQjkb1pESY+/N1hnC+BRn13htFEVcwnj051QGvBIUQLfDz+WVZqY
K2Hr35w0LvFwosTpIHx6PxbP+TCjnxsN4sqe4tob7XCkvNHu7kWaeFUr4o+J56xP6XEzFNy2Lkx/
1BWIuQyOqSJA/851hyCLFG7bs5+56IsUYatk5rvwVhR9K0ntSx3j0GMAn8vA4KkquLV85Rj9cF0v
pg0QIuF681qCMX+0IbEk4NVypuAiJGC6Rd6r167oNKn8ZCatAn4Gk01h7nUfP/l0V0qAxMJjKsAZ
dMSOeuI059PKVC9cTNoSbXgEw1oGm3aROOU2mb5iXOZjeRDEqBza4agmyx6NYiIzNw9TBDr6Jvca
Y+CGUTL/Si7obJmiKd1Daj8+YGPjQIC58z3MX75uOTiXl6wk4pTa2Ug/QK2N4zeuIu+jYwe1fEkV
bgW0VKkMpMlxiFs02uhGzHHJiI8ElFaaz7H9CmJ00BE9n9nTg4Jmtv7v6DOcCQYSUVmfaBK5lx/j
p/7FopxwT+xZBC8RwLNOXGTOuVnkfCrLd8cVEXPe+Y0yq+bY9r2q7JuggdbVYJ4mhGmLFFwhahIv
oB62HXtbtn0oBdYqp91pvZkvgcb1ukg5rWIHZVGW/1HUPh+s9I6GDeIUYMDOZZQ32HixyppcSMaQ
5u72AS+q/rhZsinp5MHEKuECWxVl8NQ6jKPC9Z9U8oG1fpYdzEWxgBNd1xORTsOCL8+xum2oKV9M
46chv49LdpavZXTUHU5nhFrXJC5doq+1fd+moo9sU+iu9NSNeUP4t9zFqUdjiT9KJyf6mCArNgzN
OZgB3AMpl0Wc7LJ0hkUdtl1PlQJQNlYLize1p5XIOuU34Hbn8vXA7Q55twe+1+ZZXegdOXDA5ZjT
vYuz+d9IgHS0NltyVyOAm4uGowCweG+9pKAfAJtr6owji+G8+CsKjJ8lUugaUEcZ4Z766EiIuZGI
TFl4Xyk7oef5rg4RRunLNBAfRRzKG1Ytdnj8/IT5oDO9NbpUQ9m6KHdC7hGyeAmKFRG/bJZs5ICT
8DMBczMy4lIgTwfMlTNQcQzs63NBfkP9wcrk8h9/b4ASiDVEJMJ6Od8XzyeGg0FaQjns1nCXBTu5
6HRvBy8WepKYOboEoTLEkhqT27VJHax/jWl0zN8seZUicPh4IV4tXBj+Hr4bGgyuFqka8r1AtgrY
1FsXEuaoODJSQj5TS3p/9uWflzn+E80ZQmfs76/qKpLtT9qkgW3+MRZOPGF3FscE48Z6kl89Jgl0
5UNK3aJ1pZmJ5Sj5iwgaA1nkYf0HbnU1b0V7s9nNdoHXBwhwmfBE4mocMqHx1GFauVG0Q36DqiYD
d90CdrMH3o4ppOgEbLTVL7NXzh1fgk5/yjRAOOA/uGjmT9Lspi6lE42rpWBbFxZeQk3OaIPLruqn
G3VVgbTOwCwxbvMRag4AmW3S4KtS4KyNuU1MaNaaj+yF0zw8diSdOUDZnGegT/ZNOSuSaj67QaBi
GKaI9p3aulyZgp/s6Gt4R80VYBG/D2tAAgijVDxJhwa/LCUuHAcphnRtGxFUxZrfON0mHGDBYmLs
lzteZRprLNZlZI0IpJ3RFzpFvq2SU6KKae2QB9bsFDK3T/fMkv/AL2EJXKgRvltYlIqvmSt5sqJK
U6Ykd7utLkWqgqIUmUIxAPnp05nOUfeORJeH+M1sKgyYzX9QG9IQWiOupCOVtWiKt1Tll44tjxp7
hXgp512BGRYSqUuz940ZlgnvgM0OvJ4+xDW+D1enjx71xEQlHPxnIIEyD48JaOrYLAIJVIkM18J0
3VC0HuRTduFIfVF2f6+/M3A2MOyWaQ4Y8C87wutnisTieCc4+iomd7A3/GKG4fy1p/8nOeCc4AY3
XCfb+ewHNNoF1OnuByt+tkybJvZ+LUfRa4awsd019AlJ2ih2qiq4+zYH56rRDrZmIt5onwOKXU1R
xVS1ORsCRl6+8MRZkwr5HyR8WDLzI8pSaNmdgk/joSqGlXkNih3MZID8YgQ8Tf2THdceY8Q7tmgJ
ZxUXd2LlvtjkFhG+Kt/cPLNaabOqAkqRvyFkzLRufZTo9N3BqoggUG9ePiGh3iPiwxCgN95c36B9
Kra8nG9h/0tvACPkRVfso8darg0VIyGwa34dJZFxiLx3fiigjY/KzCYAQznFVY0t2bAZiKoI1BWv
xMZZqTjr6cUOkJtqJUaf+xq6hA8LuhDlgsqtdAOuMt6D+ee+/yT/w+GiQoac7muUlPaf507kU2WK
qLsoylNHxnMRuFomuXG1djmUSPaFZFGUdFZWJVSTw5KXFYjKwWbhjxL7eYZrAwK5wfXSB+vXblQQ
sBINpWbqSU8oFdNINejjGdA4pG4Xh5+7qFnCv7W7Lg4DnhiN9dc+wrvPi31cYHyMtixEU+9hCs/4
aYkKrDETClJgIF/2U4UAStC0eV9WwOP2a65WTFNhJsoDhW+p5+nq+jF8qPFHLoqYLiZHvj+n/CXH
HGfo+fcyY7hvChCmByxPx1EABwOmIuudAoOL2yNTATDL2feCK4vGbBSPypUSUJEfPzZ49dLJ9Jtt
rUxfYr2laf2dxfP9v5C97soedSwi8w2dHqQrZ1nRHuAGkiAso2Rr5yzIB5x+U4yH+bmO+0j3x/Ck
eNAnKhH2DKbosvWIABNBtr+hEyH0sRk1EU9kjW7NP11BgwQZiqBsC67m4LZ3W84NC6IJmMeZqdXe
1lCUtJUZkACjJV2yW5hMQGn5tXTUeW+kPempQV7wBEdusYWvCPvOOH+G1lp7Ko2K+kQMkW9Q4jHX
R6Ux0z6YQ7PyGbJCaxpJAZCcGrWu7Qkr+1tgEKXpuKlZEH0qZ+pMrjY58bnH+rsDajpyjyXKPAib
xx/jFlkeME4SzgPg9SibwfVWWjUOqPvlZN4WBU+mbwKTxdgILe6ej9U6yWPKG3sy0/4sk5gLpDPW
dkehujpIE8H8wgEBSOmIM0jc0fwZMivPHv3+uDifkeY1YnK83p1O/Ji+wU04F+Pj/0oPBS0HIQMc
3wj4058JwmnjNc4wNUTUH68AZLUlNCIN/3aE5OvEw8/ijU5c4KNbg4Yl6sNvXg5lUI6dq6SwqR2F
DcqI83wW5yREUJp9h3PQxSOA0lGgIDfBnKlMohDPwi3EvMuv2PYvJ1fuy+bOKjZ6KWULqEjq8zsd
PsXqXOitdJ9vrnIjy5H9ezI76rmT4ePlf6Tfo23UqsJ0k68l5mcvmv22reAqAguIXnZIapfKvTX3
hTY/JFNA+VGo0n0KKjRGKvpH+uG284G5UOyIZBZcFVux07FY87y3JVK2aZIqF18j8O0ZSCTC8ap9
TGWoYpCgYRBYx74rWhYlrPfgEkC1X28UjHj+PuO2FzW+yFvMRQ8kg180quoiOf5UY4m6WzA39miD
A0m9Z6MUxMgqHitvrGVbWMq5F1WOcPUuWdQffumxUGJpPbGrDnQ6TdlV4mqxEenzFb92AusMTmyc
ZvTeWnuzIQB0e5WT0qIUNLEm+2+wMsIAiZVcfyNKt96TCRIAo/TsQ+2DtdQI06YwPhdN7NwqvSy4
JRPqPBkNJxmcMj0TR6Aqr72SjRRhbvlx3acx+nDWe30mGBPUVi/n/Vl+fElmAiHH77yXDXXIF5yW
X/UbFezr2l579528fCk6AL7WW25YQa1e4UI4o06MWjSPu0NFGqf5+DL1o5AQsf3cO/IURQ4UrQ6F
97bcDjhW+EZ5XhQPxipTHvtW63rK/tTz6CsHQnvn4V4os/GPmHTkQD6IzmOeIC4llL7dvuosq4cM
2hSlaII47wlunQNXQI9DHWSTj3WQIRxW0IA92wE5eoEx5PoUF9lNqNvJpt5zAhqviSZhnBTgwwjw
zkxPqKXbFl+0iTLZ7nJRIz35i7fxonyVd4nlEpiT4hTHw5KZw2cU2QH2XSYp87f8ynshgMEXEQ46
1BkiCC+8y3hiDuhaqsLosGdWOWSKU7USIDiUE11IWL2syJduFQRbYmmDjmtAXeHD3WYJqsXTi2S5
SiW3z4e4Bx1vYyTI0XJK4N6uNoH+iyB4cDWp4T3V2uxlXxbuRhNq1osyA4K08ZfUHZhZYdAwWQy5
EvL7wMg0yHMpHeF2NfkNTMbFziSj6aHLiQFod6hYnEMXFFZdj0dPIKqt+J2KeMslG6H2S4MbleS8
PTgqdswdn2+q04059uN6+o5p8bnU1roKY2fempts8gy2P5taxMytFuZngLtgeAj8YI51yF3idOiL
SYBj55eBXUur+EVU/EiMHUystz9xv8qZKiDcg09z42hkIruXXnA8xa7W52lS+4Z+KlVYyfTcLpvj
nCqe1xT38KXqNi+6CHzys/W9bf0TC+KB0D36pmdWuFyhmhlPRRkyEoNel5bu3hJjlShvT5GWFlXs
8AqMUGrXQjASiEQR1MfP2LpE2qJWfhWYz2qGv+IGW2XHvgmIPPHbOiIxWmkDtr2xejhgJVjqbtnY
ibChpNAWef7jLmgJTePEdL7+bnsqwct/9sv9veQ4fxHECU95qDRUJCPq3xDg24MrTzd6ANFhjovA
yIQxuGvDrEsmuNc5WkowYBG9WP2OaCCWc5OfGNnkqURCrsTWn5D1iDa/BjeU8rg2YOqkYjXCZjuH
0juhK8TaYzuqKOtyYbdWGONwvCtBMekQx4aChl838PKNHzMsCVo1eRPdb6vBSN/Q3cHcKn5n0S+U
hswfMyGmIkcdkvKBOke8kdDN8QyXwrYd8Vla75URMsdCeStGkt1QJk54xXJQs+47KgJ3VZEo4uad
QZvp5QDw7/U+dvy2ArLt1NN4YwOQ3IX2RoWD7P02corNnKY3JlVIclX+kKQD/945KnblBY/nVOIx
KA1wxqQ2rFMfFlxyEbMFytuP5T/gthoO1P1NBVPhIC1CUsHF+h5KHqWjxXYdu6HhrWrTWKKN3oH+
VUDxiwjV9D236sKMlNtCjiuM8Y2eZea5uXwYAxgn6JZGA51tCcFcXGfmzAD59Ziat4lTZWVz1vMe
AXKH3XyHllMtAcutKo7PknVy5xbw52o114bFNt33wFTObg7II8YkiCASbvWVriZyAbL/takeNznu
vsgLsW6uinN2Zek/Lj5kgxewowVhcUn2jjXhcXd8PPLsF7dRYaiZ4JevKTKOB/y+KHGwrABtUrZw
TPk1pLbOCFTVa/dU5da1ub486hxoTT6w2TPFCeHd5ILQzgkBP/p3TufUNyui6brSjmNUrL/qSNop
p0yi0sGu1RuNVEgAwaLVYUdnBeP+3hi+cwliW4MQ6QEIhyrYpyFCHhPR/+w5pA5FZI83DFQt359R
25Kp/0x6ZVYNhwvRdQWpe/mkOYpdC1FE4vU+14O2gjHD8FauAwMHPOtATSuYNK1dA4qsw7iP2Rmk
zT3VRnz7R6y/3hQn1PGml+wUtEM2z4RtoiGxc7qDBWXrDOLrXgjTR+fE/qIDimj2pPiiAAO9bsi3
n2UvwAYXRUBBsFlS1m13ydg4a7udQqCdTzHC9DpUCxhSXw298omh65NbMOYQC9jb+VpgFa+ZGFBH
4IUBvBTltx4J/FCzNIeRZVQwl7vejFBNPipOEPOvNbsj16VR5VzVq74IWw+7FeZQt5ENjJXVbO1a
pu0uftEHQslLiFk3g0Znapso6FsCkWxupgBw0s1/3UdHTcno82+Q9RSj14EdVZkEKZ1kYKWvy1nm
r3X2hw/F9HpbLk5WK60guvbISd5KGmuxhavdDFoFjgTsYADQxfYdM/6hB1Ctp7mIwbCTPefMRShd
hT/rWefF2Jbp4s1zBsLLMDDJV4deppFdW4X/zn+7Jj48Vr2fRoob5jbsu/fhiR/6itQs6V/9W8w/
y0m2SJ5Cog6lvz/nhkBS6oi2hIjVOAY11M/b3Pz1949OsjdkilJEbWf2VASG76cghB/aIlb+zTJg
qfYQ4uT8lRe3W5y1mq1owK6Sps8bk3EMmJpWUhr3uQDhIHiORSrAYoDI2tDUQT15JRsuNznK0PdB
vyDupmlUhMtqrf7xclOAh8c5/sX8jEe9/ntZx5KKuS9Gxj3q7G216QWxQDGMAeOfnZD/RFbWeANv
ohWHwU3tWE5DGedHwq3JakDPPbyeTX1x5LoTKzYFhXCw87+cLXdqr31L5gDsoRUv8PzX+0q7j0T6
eQVAIC2xNCSA7AiZZ6vx2B45uOydVqi183H4ZS48JzgxDlPYmY0qWB6wTOCnAKJ+36it2EPyCV7v
zMTxLiOs6dgVbwRndgrdA8pY29kXYoutnw9L2thkkPnGRMTb/j14XXUnCtvJ87M/WW/4LcWh4NTi
8cAtJXvlJ2GzHlN6XdxaM1q7xbFMqdmSlAWITtVkbRGHwKT59Mal/Srie1ApOhDKrIg9w3xK4bEV
lO8ZSyvjWYUCqBsCFbiQ7w0baL+BTD6lmopWCIASPpBtMkOIwOTvHQi/qABC3UnQyn4/i8SIZYDu
jZ0XmR/PIwuezWSo1OFB+qXB+ZWyvNjGYycS3xfupbKatDPhfg8OI9Gr4fdIClj9c1JXzHI8QiVs
vri55c8iUAk8q74lJjeX8PHoNLztvtJjEj/GfQbne2UfweiVy/HuYe8w91WwmbsfBDXoagqoRVRD
Qu6rtSZk9uSLmU28ZDcn/sK1/ezk0Rtl2/gPq6rPNyZ68h+bNPrYV2FCoHoIkwttIK8iQ9OEMcSr
xIWOgbsDPfBaR7Q57osh7829906H45ECv6Eyujo+eqxWZAK3S494b0EXVWJgW0iWGwus0Z2pJb8v
NfrtHFIFWX3p37ve1anlk03mItDiN7+Ih1CXKWQfqrAeJK9DOnY6wD19ykgKWDOzbSvW+g04J/08
72IHjOgMCXXuzc373Pql/uYFUSS1E+JauSaRp12uS1I5/ePLf8APEFUdrgO8lHF1eOQyXCUb4Oot
A4rnK/AV0hnIYfyW5rWX9n0gE8/1PVMulRGQGQVqlUFuj4RgI1fEm/gcfF4veEy3LbiNasALFitL
XdMgAUsMgoyItHwBrbsZNoUq1Pmg0e+FZuKWZiACeeqpjnwPw883N0ru/Xa5B46r1A9LYTLRp5NZ
KdtL2UbQBwyzmSeyQh+w2SK0u/rehPQIqwtI9I+29uQasnB6ekS/AtfUBjfT8OeFOUGgmHilMSGN
xyOeQhUPZyIrV//gxHPKgAOGmhzYcYntcgSWoxKtktXdTxwod9dmWljHMjwGMA7VfG5SylSRTpxy
DxXvOKcnRg1W4SXtInsZnRw4edLiNZ33Bi9mPqwYxhHAycEMZEo9jJKkfu/AVkfcX6/7TSSxueiY
lZwI/m40GthdAEZMcnK9oJlmpVQdkJCbm8fJlw03Lq+Ot1HF95oApkLC5//YxvUiEx4JWUKlV+oQ
ekIsc5KcrzzVs2IwAWBIl5HMc0JJKgqIYonqAeW+Qy8Pq5ziZyI56a0xk6BGgt9HgIFm9Hm+OPsf
AbrnwP3dIlPaD39L2kxb53bx+J6q2GGs36jjCOna/7rjIVkevrx9q4x37sa0iqlSaAOuEMvZYuUU
3kPWLtLBwCnqmmit+i99/N78EqqU4Xq6jSZtZQNSk9i7Zbv0EGOt2k0PZYMduwU3g+lFLcx1HfvZ
hUFMp3Gs+YEe4mNT3l+Doe7ahJju2Z2DL2MYBmMh8SuQLINaV7rQxjsT+FjBxQTnAUREXuyOyy5S
Pr7WUgVZweVj6mup/2LCUwYM6TYL5g1Fh0X0sdjnJfkBxt++BxlQq0JHPo6hmSHO/R+PGljjUEuL
xOtTgimQtOCCFMr4Vbg5GZDxoWHRRqlAtcoDeldHMKuxAx8sDUsMQJC9vmstiE8DQxsFH+Q8OSiD
rLoM1rOgUkdJoliMZ/MyE+hUwOdsf0IefioyvT7aoHBcx8OfVdx4NTN4zSPnD/Wlx3AhZQiKikqE
JxQIMaNbbv80RS9mQYv4Wjf6V6KJfJWJNFLmvctvMEwHRX7vEsyaGDQzQ8X27KlSHER2WRHV49M7
x7wpKaRpbdLhMOADtuReui0vy3QFx/I/HdwOoICApKAnbhuXk3g3K8HWG6Cw7ZJPVkXRy7l+BUJb
qr1gH9MTFlNT3CKhBM3sR0wR0JqD3ClmLQlJ1RM6E/d0de2Lf2em+fM91RqCJ7ffR2vOWaN50TLe
3J2ctZFjiUo9OMRzUUVfe8wwnOtfLKyt/lPJ+734D3k+vQK2aj8T1RQmu91sh+keDgm/ETqQTl3x
z9F03jFhHHhinvhzVmj5G7IFH4SdDPhHfJVMVXkIEERP1xtTXgObqSrrO0ussPO0Fwb3b5BkAF5r
gKN4WJ9wdfd7dWpX6OkjuLSpB2euDD/DxxrLFVaqwYKDk/voGpp/+jluXl54YZT0wwZgtaEe8jNB
QprFe6QayG2zy1RjwcIV7P/XENGFsRYN+ds5gc3//D36Mr7CyK33tAWVJo5/TzcmUsnb2xlvB2sR
55wqomA+hhXRzE5AwDmCxbvWDpE0rcNNWUXpOdTkCR1ba7/dY5mnMfCYpOnx9zO1IvoxuiV+BkQP
iNxDAkt3cychcbMqcImPoJLzotHzUIuYxO1aTwYnUO0rFaTosO5fNvZxzA3Rxvexw10vUwlCzRJT
kaYJdhwwpivjd9QAsQbfpeAS2hfPFXDehanwqNo9gXFZzaZO7Z0WBNFbeNQKVVrguPLBGFOEtLuU
zdqKSjd9EmK6UBcRhmjwia28e581t/DQemTR/UFCfEIjLy7Bmf0dzGm1o9KJKFW6wsFhVHX14IWs
Yl6/l12fhuYgdoHKfzptUYprMmctgXKUhraF+ptZvA5V+ZJvVUQIHeIWxFwXOeo8cXKYz1IaBPNH
nsSKH7R+w+Ns9npIuo0mcuyMYDZJELiqeYJ1go76KmzCZD6LpIAZxtMuBj6fFeQ5XIBwMJaPwQMm
DF6PSY4zEHpQW19m9N6mDewCnpe6W2J0/Cm0cSYr6mzBAYnavG+nRw/3bs4t4KnjH9KmCBqOkEQ2
/xNSatZ50s+Ka+HiMM0HKT8qfJxsMNjH85Hw/arZ05064tvEPep3wgQPFAStS+UQw4t4Y8yV1cPk
1s/xSM2IHhH9m97C9OK/n3Y3+XmpNxahBLWDvz4EMY4PHzAZ1uBjAlP5lhWcljSYtq4Ce81ma6SZ
sUwOEmKE0BPOtWXiwppD+hn2IDjwP+VQ1n/e0Qms5xP8nWe0aZsrePbqFardWyxP2D7zBB71H3kC
MCYFkdxa7UT/5yPfFpvX8KPbfFIeiK3CHltW8emacApnXEIxsne46wgaTbJj13Ol/udS8Xsemy91
wvqO0QtvwRQuJXJHBTnLaiiin3LasN8KddUUzvHtOOGZukFWiBjXnnvikm/MN2U/gE5Ku30JTjl4
mQlSFKWmqTPi6Xz3WiUvjBOGvxCbBdtTUJYCJHl03mkAHOvBFpCPJrW+ePjhDswh8mRgqwxmays8
SYOpUu9eqBser1fgzs2R1P1mdRBp2jCbwK3lWo0L49kPFdEgTTglBl46MnfN9ur5Mb7mDlgwfe71
JZC9cGBuhm7IqYetF9zHq7WP5eC1yHhUlxAhE3LDKbaV0txdiXYvtX994JEQjhcVVE8kfC3ZP92k
MblSjXf/IndmWm0mxuEIDIvciIHjmd3FCB4e/bvzyBCDkvcMtzj6Sin6DjA5yMChGwDqcpN/hu8v
tD0u6xZsuge/w6Dfb/8xwla9yjmFqRYdUQWkRsrUBUppBvFlQGykaY2Jozc+hLvYTAnGD25j38Va
dprVjqIq3exx23Cq1jYO98njpIwpkcsmsOhVoeGLZ/yj3wpmmqriwMdnmcdM8h9Q2zYo4JHZT+H2
JW046URjODwpjeFnxC7SLja+NgM2kMfE2UObUG+QimmR9rt5sDDVbgyZr9ptz7H1wy0zhR/Gb4Sg
b6XWooIk5N9dSSxNR7QjT8cBkHq1dOrzKz2l+3AOuIs8ZTHcpSbwK4VG4Vif4doIR4yDuK3pkBw1
eG/FWyxiSvnqWjptJye5eKbShonVE54hByqINKyZ8nogHVA4NxitkjLumSrLudERidyuya2q9yMt
rgyfsHMn5PuLFlhpPV9LUz5b6maqb26QNjbmQWCdkItyPMMYtgSBysMIVuTjbYtbCQH0Ld1gggbB
g5z0TAxBqcVev+Ikl1JunIHCLzywRGApLqpIWAh12xEy+5Q0uK1gOzLbYypvDTMaSDhb6Te+hQKi
bjd8QxYjGzVuLUv2/TFZJOO1x0aKDq7bzqVj62utVKLi5hlbpdE/tb7r4astgbOrDUb1MbYqDvxh
K2GcpMFH/qRZsq6PvCNm1I9zKw7ykW8Ca8s9w4dJvj9F9gSuZ+H5AoUQIEWAaC/1G1bwXyyUh+nW
xcxJSa3lw2Ao+kQ3g9yJkovSIBgi7OX78ot1Q3l2z6+2nm993NSzRwX0yaXant1kZ8kiwbec90Pa
H9xkijDGcCEgzfy41VCgTDIZDTyUJJrFCtNQHgabfsa+1KK0xo5VQOvLotuWKujLDj5kM1su/TQG
yzFxv8co63s5CCpr0GnkcUX89nahqv2bshN2/J5RCItlSUulAIAThgukCHrNgkVoDELZsNf9zIwN
Y1rmW7ON1GD/OGKJFVRzSLtJE+ITb9AAU56+0wmS2l3EDHe7MEbINQpBMFPmCnInOtYIE6sWylb3
qKTl/AJ/otcPs3GkxxMwUunPnaSZEB8Uxq80wjSJdPco7x5boDow9Ut/ZUN5X/98DrW9rzqUkQAY
54zVSd+JvCsBidk5ztablBS0KvJSOsfxpzETG/noZfDrDnczBse0u93t4Wpc5s7wu8KD/8SzUSxU
gO+arJUhiGPi+7Ca9JkclAUfgEJejqh5VWOtEZcNZMSn5CwCzkcYOfuUugfQXMs3iU3dWt/56ZpG
18Z7wXJVRvft8zSnCw77KhfYbkLu8bmUCk+6e9avkV2GDhO+Zgh5McfVxJw7jh1koCi7/C2p/HXY
fnu5RTa6BR+dylz0RWxCy+ZTrPzIOpooLXJrp7M2CPceodyxCUWlurRkK+UkPgi0U/L6cUGstO3T
wmve8AGxQjGQZF02FtYt5epR1CXmeWs/UByqueFx+yA3LwgXxJ7+FL35+GvOQWPp0a5F3rnSJhVH
HQde3/ee9KoN84Jz4KsLvM10c4muGFW0oZxRPS/C6bnwHKK3OSoJCh3KxdasL2IFlqnYQlIPq9hj
aNbhMp7wqTn22gHFHx59Kr34zFq+vv+87jtxQC8ntawGSzA9v1ShskxoW3yZs9umcv4FWEAO0tmE
WfGIzO5pBTLStobgevEyu0SIjsFmHwrQyGBkE8eJ03PLrn+vIM4/8SfIwAI0GETE5UTnJoJm1xca
JVFPAc9jkSw9A7MfL97Z6cWkVF37F6t7MiOfP2QU2N9SndDRqXtcfZ7F/EOwNgguimctJ8vRdWip
f+2FddYcy8lfj3h7mqCaQpI7WUXArb+wBYgy/LQgwU4i1X/Vq9pqr6EqCYHckeGKVAhMnNV5dQrs
jH0uzBzRG7BVZbUHtTvkSE+GeJoLzq5i6jfuSWomfBB6ONebJwZVi6qA1vuKQkCJb4yUizfMn24g
lwHmNaHVUyj+9vmvViZLTaCxIbaCsLT85WhAmp8GyGVcQJPgvlnllxrjuwTJGGmimvVkfIBv1G/S
nXMSI82aWcDiQPrVMGWw4Jr70NH4YeQ5QRqB7Jpgma4ekCXPflf2Kx8BbKNBUp5s1j52eI4CMBsq
6rVIIOIBzLvYbEMKUiyMhke8K9HjJOekw41yUcxCFMpP10yMtine12ssbBpY90SLEYzNy588ge4y
iIa5QxMzIxMLkveLPD2rs1piM0ZDqMwWWOmHF3sJOczbBEQMVr1wGfxRgS5nbn4d8oqIH6ah6dP+
9VoiL01klWj7V6IMvn3MCP7CD7UjA17uvuaOHn2asIvFebQvqAOgBuiT37BKIIQCn6aO9Q9TZ3I2
vK+AVOVdzCZH4ZEtAl2grbl38ckbcMXAUUa8ngTZiaqY+yDv0lPNzZKQL5INPvFlerB4YK6uXsjX
LD5D/Rv9pSF4EayVEQisXt2v+ov3lfRmdbhfEw8yzZxscSqWhWZN4g3AQdGkUIqZZSIyNuBXnnoi
m1fw/noKoQ4mUZvvtV/YfAEx9R3dG9pcJYvrNkI6OM1ns1fjb6PaFpKiLkos9VoYpaKf2K5v8gES
oQ37PTDrDPovgCm4MGjgLBzBP9InJvlkxRsU3agWkYXsY61dNrwtYmnhHFq+p/AMIwCDhMmbmOgB
ES5+M9GlUiWIIzXfi782sD9mnEn3mcclM8J5AFqox12tM2Whun/in8YPcv8xb1x/iIs+kdni9TbV
CH60wQek3ZIguDOSzseXHyKlyk+x2f9NnhNRKAej9S4UCI+ffIYqOGHFNXR085H3VMJBn5hspeYK
CXwhKFXi/4LS7tuahUcX50LSbMtv0+DGwR596Km0ksI8AxRXLWF8zy6erRCdXFk7EHjz0HPMHnO/
sGdAyEGKlqw2IxyWYmjVvD1v7+fulAWCV5i0iK8TpjvZauCeJlTONTWfr/0gEVuYX8fMXpU7UOfr
YAE+5da95M2j2+CswyFyaaUxjNxXTG/waq+qA5EWdES+rKoQb9oBuNYgRnAPm/mKuW6AIbPwC94W
4zZOept54akSR1hGxx1FnIPhlkn/5HchXHRMrfWuDdXRVMQZjgSBcsWLsyzuT443xYeFI1Aq1C88
3jFVZwm3su+wtfWrM+h273FMSHCGb7aFrA+VPmjqYDr8PaB2bRKVYMPqYULAlvq1LlHnJQk31Gr/
mjBbU6sW9gZZwhvUwWsoA26Pa7PbrxcunbjLNncn2B2Tb0cXmRyCeo8K0kGImzejat2OxH+Wk9jA
d+GmN5eNE0pvvG2aax2xH2ol/q54le+xvtwpbpXQXmCtaehvWYtN2NXzr/PneZYvn5nbfSv+wAz+
hx15ZMImPDk4Vqk8ZFd8/vw5nLgk61Z4B9Ge/AT8VaKl0LhL0tUWCxf+iCrBaoLCX9+dSJ0chUAE
7uMr3Nk1j27Tu+8pwZOPFOt62DQnGWH8e3OFWxSwImuTQBNfap+RJ8P3UwQ1Q/SqcpUvFwEiXaI3
sc9VSQHZxmy2LSPhdrzKLDuZAdTYw7jjZbHVfUZdbawKmkb57g9LjfU6WbAWVzgwc6jVXivUedfG
Tal5PDn0ecCyPpbmsmdtggS212FEBha1NEM4d5ZEIkQhUreZqaf30uHT9QdTNyMkZ5KGY7NsSqs4
ZWRNBY+E0v4ehrYaG5/mFidHv8B3Eif1pkesUArMi6DBLUY95XLbl3GHPcuoMh+8rcmNO1q6pmjX
nUcj2izDsZRpH8xpjSJ3gVMG/8iO9KiHDlwhplA2Ejte3o+UR0g5mLpa1xcUpVF/mBVs5VXWbOTD
qHvct3E+Ro2oRz2UkAtJf91yKTBfzHcym4nh75GeauGu9Frw3CwchFVBEahPfHGX7y+0ie7tMU/B
nt/aJoooaaR6tibh+C8LNPZ/YoWlQtmYQFgaZbIzWxswtXDvI84tlLIxKuEbiCC6D8rAPV39j9uP
u/hdwyrZl1cfqiC/VXcWsspCflTViDM+5GZx4CF31TOlvizZvhZeEJmr9D+Dl9frIxIuvKLO4kJl
9NEwEonMLEfKIFEY1FCIcuSYGI02KldSuaTCAf2MVlUnzVwF2+bfWmImsPJgqg1wxsVoeTO/ST1g
HO9uc25l9D3VHceubYNChedJqF088SyyYaPp/EyOPfh3xgzCakKE9oi4i0XJSBWigNj0Y3J1WVfy
wQNr5LZu7vCgxLfGxPmpAik6sbAJiPiyRnOboPGRlftufjlr7a/uiiPDz2LpvUp6p+bCaX+v31Vr
2sBNVmGJPznz43c7OY/C1sMtdJdR1FBAQrs/G0N99rYEG/9/KxYPLByjBLZy2U0hkvWsgCSVAznL
4+GGKBeqSWXNuhJ40Om6rnDt76AlLtCGAbITev5NV0LU4SnkGcRSZdt7pOaBy8CPoeOe/YCp8D3x
uFlGkpWxKpBWoxPc5wGx+I0m5aqI9Dw4lOfE+qp2Y9j3Mm1ao+nhDCy7VLjwZtvZXsxbmE8N3NGA
OC2bnWGH8R69qUIWMobFcH7HEp/GCN5sE+1pO52eUKWlsmMzRUJt6gAotq6iDoMPxfmbN0fjVu1Z
Jh0QC10r+g0EF+tI2vg/+Nn+NRN76Wm6XOasNSRF+PmJsMx0kGlo3eXp51JUvhjBhScXTmu4ZEI9
uhHTbXr3Z+GC6MW6phF+LZeH80bVh0fY6ajCb1vL5tklAE/7OWlwPxDJU8LbfE/kWU8K4bNLwYir
/8SMjYKjMpNq58Vvtuw7aT1nKSPlxKz9IVtABOgS0oUw/VgTYK2r8X08xbU3XH05xXUOuP7/YdgF
Cvf7Pe1mynH+vNLTjmcQpu/xLy1j4tBbA6h8EiTIRlwy9maisudBflDJo3baMHpvcLQSX/Uftw4P
5N4rPU37UQjfP2ordHA5QPuLpHXpMvgM+AQ/s5NuZvdy7FGf4PGvhYhPL7+65s57mJ9JCP/bawOW
wJvbSBPywNRmuzni/UUIB2uIB93IlcHYzdrz7M5feAQKIgHRtxkUNLR+F5exF+fsliXbwo6l+5M4
9mMRjf+XXaNqCbp1D53+NSi4UkYyS0KcYwjQTUzV4JCjnHRpQ+qczCpo0cN7aYg0jbomfEyst9uy
9o8I4aSrjE4qM7s/U34AyqPaaZNzujjUlpUFUDPdoo8DFeedmI30FllEKlAMxfdFFDl37lowv+iD
PC99Wyo8jVc26s7OZgQo5HCxRHqVfrkoJr7dupeOfzKDuaugHRN3XIyWZoQ9NB2a7SmmW9kQRHSn
YG1sUs2C5AE7kAJ2ZVDbl0OAWu57T+EJdMRQr2a4Aq6e48cVOt0zTOYpeCnHyIj97ugdFeHksDLq
M5L/xSq78erCWyH/WVqgMSPBMEvCcmxCVrMszrT2n6a/9lf8YNog+e5KJbcfA1PTfICXRBdHDz0E
u0j7b9h0qdemBZI0qmwxk9T8hNpsS1p/HcdLpJaRWUt1vWaZFyk2NfapLjyB0VT2xTOAyeIuCr9X
NCtX03ctFN/lKM57Qqy8HIAQWF3nAJhBp5WZBfl0kyWDUplQaySqs/Vn2gzxT4hntIcxznSUm41Q
kOp9NVshbsTbDw+30pZ+hl6iB9GtHzh4aKzstqqnO3y01v2UhDkOUWX0PxdMyn5ESjpKzbnRNK/P
MuZJeApgki3nevN3TKlfBJMr7K7IbISRfxOZ+GNzPQ92LpW2Vrz9Ok+N/4Pa+CNlI0foSp8KrabG
AckjrrJTnjB0SBP5vEBZlnahRcz1V/lpj9mvUDLQT0Kvbu+dNO4ZQdo8nwfDZNS0hOoSjStf0DHq
KCAx0cO8dhvXjBF0Nz81DzvrlgamlNDZ5PsP2GsLU/z0XKylYCzE8jciVM6cPzAdJVexXGcXWjzl
D7bQwsVtWUh7GrXWygtrhbTdMgDqQtHVWh1ENQMikz/AeUq85qvcqboNA+AnXEfmE+IsY0NrIhcz
SKt+5XR9MZVOWw/HxlzL8ABulh6V0qzjhLp/NBRR/lmXCMFjGg72uIlXX46rK1bqbJLamXT1LpIx
v3YnOWVlZLwIQy4e/m5HfG80ddvJcMnihzgfiteRG2mBQykjON427DGRHiKmeZubTyAfha6w8WZt
jDP13RKtVQGJyk+BHvCOK3iQpULrvT56/k0L2IPSgxUEZLLYh3o61xapMpzX/7zMAKlUfmL2Xc9M
FolgxSGUcz5feRMpzrC9dyiq5AZwoY9puCqmoBmQ905Jcvuex8x8AHXbOrfLvp881bIGiQIU1BW4
d4dsBljXl1dx6/MKgIq486P1ZFvt040Xw25iJmXfPnEpSmILMTWdL39O4muhkTvDnnfhLBuAbdMe
pnW0i2/HxkqfOwyIki+ajMM1iI+Qj4gIHJJqzSWRYGlJuSW4nRuE4bvTLuZHJ8KZ36BKBI4sx3i1
qQrZBttzUM2llAt11fWRxt0K3cW0PXSP8ilNlP+6GRgdyAqlOF1qeJEm74oaRh4+5TygNgxAfMnM
qJwKcEMD+zuOB9fteY85LhmYP8dQMSZ4ME4mcHBDQ7eWsnol87ht6lcyD9EyUkp07wOh9/f6UjKd
8gwyrMZAy2Acz6OWfZ4fuYK1JfyFScdugwc7gOECODWRO/fKXfcTEFMSEl8BrCD3xFCUaGay54Q3
5eDbGIz8ykJTLeXvw2e92+DjEJWIyisvWx2KlIc4drFB1c65tEMOyh3sXhvBkoflzFlJWFLZJR30
q+kwTaVAmOYtlz0s02rWb7L8fbXHF9pdNgcX1SZQ/dqwWBzqvD/8H142z2ltZkWU40SH6fB1XY00
I/NiIwyyy1nS5s1ktRuNja3hFLSu3SFV32nodghxfEYskOfqWC/+vi3eUsU80Ln5O+mTvJf9URrz
7XPgjlJFF2MEVSNb6lCT0ZWcTx+7mcgT3dwwzzpwMJCivyyn8XnK1F6fKp7ntxCXkU85rCqL8dfV
4lEmD+RPRCfgthoeg1kfVN7QmqoYe/nCGObrNb53vjXi803QPgb3aiz0ZUzEHnizp4KkpUc+pDAi
DuhiyPU3lDyNGhksq6hY4dUYJZ1kPc/njSCKOo9t6am5CjkAUB4D2a2hU8Aqgt4uLocHhvSngZME
8BVqG34eZY7dq+ODJRIq7hCEDY+66MmQ82qyjE8Zlk7OZu2yPac9BSTeVF/xhAUPAmFtB86c8Kgr
6WfM30Z11kPhZEzderoNA0gmnqw0Fx+jkguCxBIs09fHwtRHyfOEKFtlNf+bdAkE4KnQK646cy0p
ltb9YdyXGBKP4/a5xWAmfji39zJRPx+n5BhyW5JcF0r6BjZjzrYVJDRoKOkYkCS0N6F8rAT0ANtZ
OjS9FeYAQ6ZfaS+V1X0VpXD0YHmbGPSVqC/nEyHIelMHn24E0nKSlES49+4U9Xu+TAixQocVyL0N
SfuD7TqeOcsXWJdrqso7XKYJwNClZ6pvdHEYmjtd8yHUcwJdivH4Hp8WXzKL+wYZdZ8m5QCtP6uk
RSJR1m+qkp9uTYfVyLvEXdZB2bRXsAMrB9iwcF6EZWfIrGU53dmqEpnRVbqcMhRfoWF0zuYPHD1h
6Cfxoko30+4JNyQ4dXdpAkUDwjzyMiwp1ANkuKYum+LQFrJKt6ArelThg6X9r3YfuITsXbvcIUFd
SLBltnvAiH0SA95GDYmwEb4VqN9cYc//nLlq7pXy1Cw9B2VnYaeE+xL52wn3k9JCKQveOl8KRVno
gLeg9H25bcoott6dtE+e8ZZ5GDvaABoJei3GB6KW9YrQRvblz4WclJ0zLUR9v+xOHlXBfgUAgyyV
5eLQfxzaU61sfbZO0KDlOToMTxN7qvD5KR+XL8il0s72wYGdp003rH95w7QN0dUNckramVDTHnfu
ovKDrWwIwV1aBFYPI5gU6a1LVjsxRKHE5av9W85pshkFNEvz/8Y8YX+ABntbblO1F/wZwrYgcM/U
CZM/a+prO20oBv00Dw8AZ7JjcKYbKu2hun29/1CAwsl5z1GAYEHjnSfjipzBisjd1YLDVkEMvX/A
h1MtAxUXeO/saM+fozMmHrm0vJtp2SxPe9RoqEkT+x/ron4cvWItW0AQGqeEbic7UqD8fSd8zT5+
/EVtVrvEs9upAiDXDzjFnIpxUBO/SeavVfOUmFjncBZLZaQTgzeW04rRZ4+oLhSh2r4+2sI+3WgP
Tzeaa28UJNmnHi+HofE11dfGNrmWBHjiyYlaTIYjMG25QPS5oRBOjC/1YqtDq0PyzqHAFz2P/3qS
NTLFkJeTBn2DiqZV5Xe7IHbRhVDPfSIHwIAlZKCc/xuHDTZ8wDPl1Zkh34/kitUKyoP46FjYcnGj
QGouimQtjrU8YfSjaB5igglRJp2srzEnDQcXM62r5vQnUETi+JeA/74+m+uGnSAE0GhcmsR/S+cu
Gtq2zuuWm461CfOwE8rhxOgO6GTTzYMx90o9aYv+Net0XE/AW/Mj/AeIBgFROvkaCXKAXhxSSIDD
QkCzqJaGycK1Gp64unVjCbwR0DN1fcvgGPAFfcU1Rs3Es3nQ7gGpWrNHaNQPWtwOfnpJkOpri1M4
97pruPMeqNpSJl6XmxsEZufuPU+Dn6IpjgmsWAE6sbHRWGEOFohGh+ihANHzvAQ9HVhMJxmAeqxb
TBwdlIPi8yyXqxG0qi5ve0asWZJ6ATd1mN+CRoBsIX6jiRrQoYmKdDvpgZRniTT5t93lVuGRoSv2
jA5dw96wvAnfshQtrqltaSHOSqcK/GIFZ5al4K+dGu8RqAIPBiLqqXGMRWFm3rP/Dannq5NWOP+Q
zELig43cLp9EGtPmVDMfmCwLSzyYa3M3QrOsX2pZd9WHE6DWD33G3LY9K7vdkMCE6+HjIBSkbUuJ
JHgcqTk7KAb3J7PsM3gyseOsOBBMPCwQJVkck1Q1IuXCJgAsb/79IBJgzdc76zg8SQR0LJgiOZIc
RkhoEGEv2asxKfbtf+Gd+gQHw4zeOoFmhbwBDu/7RcSqBXsg+jyjeCwA1MGctIs6rwjrRRP8B0oM
kYPQTm5ydIeEy7df04X+MCmmDbAxdjccXxLS7oX579uzATslrm3fuTJ4KeI+TxDP8ny8sLe4LNHe
rqV3Xsmt8TW+xriAUqBCpc6BziVAGxK8K0HXtFmRo+2oRWzrmSL84Vfr50PAcD+gzOByOvQNk32G
NX6DWO4ZSPebY2EqCh/yK5e9x7CwmZAEHQL9B6eZzuMR52GxC2o9cXiwQRitF/NCmC9c6JdLhiNZ
BtwYGQYNVDO/Js7M/fPZGVXIT2iTfrxnS6EXkv+fkSns7SvhKd/OiUivz3G0sv2tBOIZJ5A4rcNX
sBxJ9j3bkAxfiSaBJkRBLi1D67R4edEYJoGyUcODBb8ZlboyEQJ+INdJ+/kxTuoNiOeJ6ePMZ9V1
3nzQcMJPS+seo6W2hT6ghng2lNBKlK//KpTCecuJUoV3nbF+B/lKBM71w6PgjBbTieK/Tl96ueHi
bZAGaKqxOG7mYblWa/t2vtKcg3zRX/AXImJzIz04NKQ7Q17rOFg36yvzFn2DLybXSr3UaC+vIN+c
VqfckgPwda/woOyu7HafhM9a6TySEFc9dK3v5D9W+QEw3wyHSZe3wzx0SUdSiqUqlfRENChzKZZq
a/ZrnwbAAGPSUjF6LhoElUNA/PAY9wzkootxKAZavG641hHWOMjD5LKybDS5lS1OOSTKj/WdJdsG
Pu6WiVvOVXkxqjSce00DgvHiB6AHbpYd9WBQVRriulTyF6ZwzUm1czMyfjzRbyJU7BlDhU8Mk5w0
sMGusX54lSvTp90vAKp1XnHuKjPYtaBt3LIuf2JfaWUBVemoiL4iFTtD5Wt0hU099o/RYSan5JRY
e6Iy+CjKvJfV+xCE5WxK5jQv4hrYOhkhTCTM0p+lFZnIWeHlpOx8SnCP0OpBnDySeyDNnyaAOEuK
4bupu4lQXpAHVZxEZM3RVzoNg4RXp6x4JiD0pIRXaJP1S/8Kn9T5/gbjIXzZLQQibQf6i19IZ60y
vkkyJizV7Owe4B53XQ14hBbo2Tj/h59zEPXA4Fh7ATDnf/8iYHDC6Uv5RJbDw1OFBmbu40qX8p/G
VBXdGlB0YKdVWdmUTrB2TZLCLBYCcVmtdW7rcaVHeBI1DjnhHoMG2iK+uyXiT3G1spbAqEapUWqg
zKe2ak1IYBNrtef3Xjz5HeVNZiaJuYaLwv5LeJig/BeqsE5Hotes/MEIZQ2Qq+iceWRZNq9dhz5l
ErR3sHO/CCkBWQlug6ayxW5qkmo5jHIsW/9b1jE0Z0uET3XSeUgNCPbguGUZEQ2ojgVU6s1RdbW5
b7OMDzJK1+0bKD1jdBIoS1Mw3hsGiytU5bJ8PaSZburC52G8eJiHH5Ccx/bc+wgDyCQoUyXMOffZ
kbGoQ+IujhSKot59DpTHM0rTKbz0Y/DfEhshnj3+FpqEeY7zK9oyyOw/UX7/LfrtOnPn8iFzzBxN
v1jEbyXvpD6+SruFbVVKggY7FMkTcOdTpnKyQObHrZVxfRtSeMrXkA/ZJWpTOIsPwH6vjSLm/tgK
fvTAsxQCCGaIIiRu2X634LjOwDou+sBmLi+HhD/51Tq9tNxLxhJYDB1MAxHF6j7Id5aVQ6Cr8Vx0
aVm4eXFEAB6NRin89PJf04dFQwlHE+5SKPjoV8oKnkXbpopvwQAIzQB5r6yLWpfXIVRObZZAAsPD
wyEf6JQ9mRgvwpwkwSTdv66bKenhJWwzYhdpU5r3uv6s2B9ENlzfgRNeDCq9HAelE6MP17S4f8/o
VdHwGOtWJ3IZ6C7S++RyonTyi6H/ZzT5ZHl0cdRxJCIwtIZz4Xh9wTjHYkFrrCflI3cSOvn5iXMQ
LNXICElr9I8Fivr+ohkZfI0pS1dfnMdRIN4pdFYwCDfU/5GXehEiVeqE1kZskLvJLeDmB/5bFubc
ZyZbJKniI8m6byKJDEg2SOo8b77b5x3/qygIoc0BbymOIVia4q5KOdqlMlHnLOZCylZfgT3+4MFA
wmKKmych9chH80f55DU+nItlV2xQzKKpUxC/RgR2xDHhzcTQGHKJcY5j3wbe1HNEdkZLG3CuCPqj
XtdmHRNVNlN1+K7x3fXfGNWGxBLfo1fk7ceMY3FDFgmniKypu16jJmbkGUQivXaAHP41bqrc6ZJq
9eHuyQQPJucQF5tUFgqd6DRs7t6tDLNRRMmMci6rYJa/ufM76YpFBP85K61zWND0c6OddCf8vzii
1J1DH7fSI/avusZA6nYAl68WaOzmbcDrMqtqsQkpHU5SvTPZuOz8o9NOfAuHopNA0M/nSRDVNVcQ
XDClOLHFIhjKquHi0lO7YofPU5AbIFZ4WGbwtfYvW2xBsQgV8USU3MDqv6LSNAK3cNt9gomO7VvM
xId3aMOc9cy8i2guhlbyABOezevRrmVogqjUswlMImnmcKbFGBvAhNeZMrdD6RlWoskymhZScDmF
QOUAbjVt82p6Hew9TVrGkAI9tNzTgOgc8ut3kEen0Fyoce12K00+ivU+eZUQPf+9fqgxj4sp3M24
lGYK69uzwdocjU4nbkDOo80Aa6UU+UowLmFodqUvQ7OYh8/gXOnCD7QPxLbkRpuB3hdyyWZm5p+Y
B9g2KcWSp8qr+8EhvPdz1XapEh6KCAL0+EiZ/CsDsB0YiuDCgytWAGd2q/7w3sYeLhGfGlvoCC1E
wQgbD0Gj40MbmIaAkYRAQsZJUGccB12joOGVM6NkLMCvTbGWxn6p6xzwjVtqca7LwHHntMdJEyG9
dlQVGdjM/sfNEhiHwbQkhRYJS0WWrWjSWUU4J0wUm3X97Z+Q9Nz2qQUqWweXShW8FSs2R3AWOv9I
vMSyYYmsuAHnQZEu8zFfYAMZR23WTLzeDXg6jsoAasCLJ+KMHuXzDy6Og7+Yy79KI5fNXEH0UPzJ
O++dmfHiNbiUOHcOrrXFIwo6KymBYlrZFTiBxn6/dTetw8Q/OziIH/0h+bLrBGWeRlvCJwUAg1Ww
ZJxXv9ph8EzhxwBdjA3Jn5rIkXgKB7wynzG0qk9/mUXd6bG6ps39kqhvF4DqC4GRaxzy1Fwpynzq
SU7bdEZnnJUz5SKp9djdbM0h4o+05LvqEakCRt4TUiJ6x3G+5HzswZeWNtNftEuxkH4UgHotJWKr
U0ecnEm+oYAgTfcaSXEKcqWnjDPZLtPUuEfBTnmGushYrGv5xWGicomBWus7HPRm7uJRd3hX4sHV
Q0a2aI3Ca+4+wfgwBsdzubC7NNFTehFGY3WO+8YpWHKicj3CbJOJyhUpefMrhnVOMLNkZAU6KE1n
4SuRQ0QgCaCsjgHfv4qRNQSIwmY4OPOKgwONopzhsbmvLhTTAFm2Y8hOOjvmaHD22/P3xYC8UKhJ
y9j6dq42xoJzEhlC1qLBD7I0qX8hE/EBARz0QMOJ2IT5qwPu+B1kZ3HRa5n7SVuzUt02zvTrJQkz
Crcrbc1p1+b35JWnTZP5UapFs1ToHftnd708Mo18C7S3XcVYVdjtiSZ1hmjKZT8G9MtERYfZ0gbU
FM5uG+LAC+pbzosxD0wBW6crdnbzNe4q7LMYIZtEohqcsG6xfRNUI/GrzcZQR/hX6XtoTM8cmIQ3
r6TICD1IztXInO5lflAHAH0v9ziRJAEXac1mc/YWtMF1LZ3+pKZtVLbdNiaiJ8RtNNNw+lduMC5b
/Qx7R1crtjlwAA2eLCaKBOtP2pvp7dY+upgVSbRzxfFpZAVp1ot34a7LDJogyY1zoTDsWxF9xl4Q
5tTIlkDL7WUUCdQv+pWEEMQXpgiCPcyjlCdfR7+5w1stSuj9fl+0GfSsgUmoSuiv/TY/dMSOfXA0
OWZvTSJeNdUNYQcN7XezwweQjf3gMeb88ODtmoUFHdeMtgM5fwVSiVJu8mUyzNwGdh8q9D3Ugj+y
dciPWY8DGp+voqm9LxNQ642P/IQ4ett1C3eQY3ngzbskIL6stXbX0H5xKgnz9Z6m0QIlBgsskPm/
NsiOOBfvwXR7aI8LgiUJg2TPD6pFp9Xo7z9YedJAiUx8HLZUPxiEZIWCLPTOPAPXRS4IzxjdudNQ
zuhdBJ1XsP1LE624VjPlIwdNRBdE1Rl/lt+AQm3IcvZwdYNMsofWFZPu17OtWgwy3RHidNC/zBDh
vEm0wbEwyFZ8+oLgRqYkXjCrvcidX/7WtkKLHEcdDuSBCEOqO27kJ+qSuv/o2db6ZQNTFx8aLmeI
enm1hnXys2DC3z7NG9pfuqkSekqeYXGXUO3TJ+6ZVOwW4jEJOQUfJWBJpfyKa9wugkaEPw7hf9vN
rONCaQj5eC+WYgG0Fif4q4oUABp355HqTiQcTQVm6VA1YNKsuUAUlvZ1G8juvq5pLl4F4KRzdyL3
sFVnjdmUiURz0VmMx/htqOcvCEsqM9EfSCzJ34YBetCDvIETJwzGcPm6wY0xfyBvlrfQiUwiC70g
SbasXX17NvbxL7GH3dUMea0NLEn8gH4ALzwUVCQi9J0fcFVQMu3pwjPcTx0FRvNvnHxVmdBHhkDW
OkJulus6DjytkowXtWM3CZkU7RhrOrUc5na5l36yTyJXTXxUeUtRhItJSSi8TSxSDj3ouJHNzFmj
6ue3uzQKZCNXFIoGAw0giDWeAFy2JFeYKT094NEzuyg3XkI7LNBu5l3OJPwuaPc83SLRvjMoiDQp
7UYwU9VjKz4VbiDab1dg2Gzat+yQDYieP61IKzkwa1CEUkNgSfd4SRGmAFMJQWDxEnnneWgXOF2u
kkxfo3Dzr7BcDCtbwNMDZs3zGy+tI781tpuyQP+45vx+8KjtC6wGIcoeuahzF9kp/CHXNyXhvZVW
oxpzjtWw8r1qIMHTJsSHqxjyUkQmEWE/Rm0q8nKAKOjUMfR0s3vE0QaaESFd9cCEmvAHKa6o3c7a
3/nm2Xp/ppKYZCA31j+SJ9CluMeUJV2dsTqkCLcMi6I3SwBfwp3wkYxTDWcE1qzQGpDm9OU7Uw0w
09zrGzA2KBlcu7bLcgLqHo0sf4i5HdsDaTAL7EOiqpnJ2qLyJWSIpTJMxs5gYyXZkefsiBl7/Rmu
ergloE6/FltYtX/iNCo+mYUJMoof6RK2bHJlLDKSU6kU4fbsN/WiwiBB2YiaiLvHCaWD01rPWFbp
L9v83ohhxLVElDQM771mYofkfvKzhNpLl0vCkQJgnaUWf+boleBnIWk7YqqQ2ptxNlAZ7jrgTdN5
iXMlJqQdR0v/b/sOmE6lnIrcOFJaSqrjmbV1aYMnocjY2ESnpAHXYC8Y2FWEjmj/0/FNiICNOkqK
L5I/Yjtkb4B62RZ54+UBZ1xP7bMGzplTx5yAzDLvYfQT2pqJb6DK+EkUVo28gWMvGCxcKbs4NUZ3
xwt06QxrgxZVHctjFExJEB/hRpSbO9BPsgr3mKSHYfzK4a9SP19AinLcfqxsv9/Oh5f23YtNKHEM
KLMb4+TSAMPzXWQ5elaVannk5TrPc8MFiSRF/FEU+XZNvTfB1TFAIItq3Lc2WiGyIqtKyZvxF+I3
Kve2ZKUjYgFwMrFL5+Qx3k5Lor6Z66786md0uIo+T1Jv13A0N6Dv+dtUxiX64XY+xAZGLQ+517Ml
tX7BgIpgxHahkthuYCWrgJaAqhMh8H4JBIbx/sE7iqYjPmSdPrsc8LijDPTE/gUVZqjWDFG6tyMh
FNwh+Yvwx1HbyZciIyi1y72bxuYWcsdAV5Pv7UlmH4LmvGPGRutEqCefQaBaaMsF+ES/Qn6MIjTu
Lzv0XbHpddG8qY8w26KyQ1P9E8jd6wB34GVzFr6VTxyjelp/0bSccoHgqqKmFEK6e7hi1k2b/nev
oF/ztnSXfpQ/OFUl8bNAvkV2UEzmoU4Lu1c5Noy7O/2YXWvkVu/xgi0KYbB5rWPdSug3a+CamAsG
F8ntfaP/nFNSwpfojpw5Uvl+giTzFOpUiMRi2LK4kGTDVvgAElZlCrbMfJ8vnIbc/cS0A9Gqmfew
IjiZb7GwH80E6Ias24dNLOTm77AKJcEdFmNr6ogDFlfwWVZn4HjaXKPl+JbTpCECMZuFGFewBtC8
WQfNgQ8doSn6DZLpIOgwL3qtvoRDUaT77tdHtlUivbeWrtl59DB568D4WrvpHFtUPmfo4yrBk5R9
hD6u2+zBoONG+K7uIDw4LNP4/pHcgPC1kUlNcM7p3kEMb+qpmlrWFjGsTEP6YbuKayqn2ZX7bG8d
pUmv7e3/3Z+weYGR7ffdHMfFHIQzKXBdMRUkcPkCLTOuV/QInZYA4YKAQEJgpcG/k5ineGZhDvsf
sAfu17oGpz5megHFgBSgwSI0UIOSjKjZXoPPXlUf33ZmTFW84Lp3wvsZYNsBe5lM0pAi11aOFQoV
jSqUsgC/9iQNYuX/kYpDwDd/yqPlMGfzysv5/0mF7tOeatLefR4RF98XaoYaRblj6LMgJDJZbyQy
zyFUGBvPWqjCwwEL6I9g4fFaUdUAOxv9ubaI6eXZLGu4y8YGTzqoj8Xzzl8FMpXbvB+7/Sdiaw0f
BTaBERbVYuR6t6artYzH66bGnugJRLHCY+TPsIbjdTdDBjj4iEqUjj2wozADcWxCwNxBAbLrC2D4
4ftVKVGbf9//1qQg29cPjoaEr4cxWiOi/nsqz4Oc4g9I5KhI/RB835YD09BTf9aMfl7vzy53dLNu
8Rx7bA6xiWhHML46frgF9aLSX4RypgU4kSyiPTKhzCmyloBQ/TF4mZyqZAXoN+VNR2HnwenP6LdI
rX39sUzUlQHtbnh0ZTrwXjM6FN2TybS3AS8W36y+Jdhdn9eKGstDu1G18qBKHaIAgF1sDelYmgdD
vMy9afbR11+GkrasvQgQ/Ot/lTK/oOLT4aCXM/s1ImwIAGMQESW5Cl0LJk/QdMUaLFFRWw6nnJab
L7QW2RWI7a6aropKaKm7HqvMPlolu6xLuloE2SSYlRXgKmzW1ldWUjukErbHX6gGqCI1ZLCPJrzx
IVuoEdJ3/HAoF8heKnU/VQv+tM7UrCGktUZAWDTAGQbVIjj0y7QjZOuY/JjiJVSzYexZUE+z1ES8
BR/lwgnnQOTVsahXYetrv68nR5fOC4SL8EXedbJwkw8kIPjQ4YK5uYP0GwLJ2v1Iy3pbiyIRnWrU
WJVg0Eyi1fCrSqgp6qxi1apuOprZ7wh+UCaVFXOPPbqgJ/mlG6E/3prUpED1PG/EqE9CTw6j6deF
iu3f2Q2Hr3gbcGC4IzbA6di141QMlT7p8cTiqJzMoOrqOh+h3SCSWSv6bVcJwp1FGIP3FrMK605I
ta48dJgI+21P1b5qZarqfD9Nk2mqCmS+CsFuJqQTlByb9aoynuGRtIB1D8pnGhh4qb/vRAdUlcEY
8wCVPUjXWK9qkqO30L0NEBBYPAT6KQrOGys6O3s8lCnGR+T8OXgSiYx0g2Uxk/Ko8IMhqBwEe6m8
ifzthAOq39YDvNfgbD0nuLD0MwL0G/PwMXfONJMrtTkozFJsqZBPqlI3FFRYDj4c6OmoZjnUMrPm
I2QrbEhgB0u5IlYnpzRXtE4kpXovce7+Hcyl4sp87ukag5fMHcs+j47shlrRCxd/wv4AR+kPX3QG
CLns3SSETuE9ZYrtM2Bl4IPCHh7fxoNRjlB/s88fZdrupO+vgw5O3TejYq7HCqUIp2D280GmjBXv
uX759mq0JC7pAniO2yJkedo+aH7VU7lMQEVinIKwJwXzvVeMopZdakLdrTdSV805MOmGxyJ7X1KX
lwn6UzBaSzPnPWE3P4RzviGaX26dboim05INQxiyvFPXyNpqi4dFrp/elB0V5nTSI6a7T7C5EpEY
c+mzd1XlKaxXnQcDjp2theCXFoN8ZgrsMuS0DuMlI0UYmQcRCJfocX5DDq70m8dHK4YUTY2HvOkR
s741//QaIPeApz7V5tRS/QD2upxmQ9uzXKAYd5LGDXVcXM7RSHV9TFQK9g4ooWvaQtOry0T/E/ut
aNNMNFK1QSgKRh6wdREVjHxFlCZ9C64ObMBZykxDvIvrp8fNxERsgOsSxRB3+s716Ew2O98O5Blq
d55/UjIQsVvUZ8O3HUB/A2ee2Pzo4IMxPBthN7wEL3xqgACPGnD58gAUP1uc9oxiacA55G28heRF
3L/3hW+fduxUAuN602HDfsQgBE/diLv/c/D8zyDSi/tw4srFQmmgb/ua3zbQWoUy4NgPXgXLZa9+
fBr7S+70QStwsmXVbDiHYUz14kSvhRiilXgtxq20JRXR12zxoNGvqeCgv521+b+vtLs42yTCQkDG
mLvV488Z5z0dzHj4kyYoOUH+3iB1qrX7IP1BHAvy7JA1GOEvvGp7Tw129etwO358LLP5Vw6vTxN6
rkR8p3Upok8Vf+NHWBcOk3Uvo1ntHEHERZ3/iy7of/Iq4zS0nYxcUAaN16jNa5wXNGJKZsHiya5E
cDsRjv4eOaZ7e4jlmI7uJzsBZ7JYNfiDhU0MJjUGdn9mSiqg6FOZ5MZVWPSVw8inNU2g2xmKViz8
lD6rp3Fsui9YvizPWpxUuP0N4LDMjz7hjcz0uUgXAXvFWKAVVBuEdJXBj0bTr5kmjtGR49tZBYW8
j8iSUSH6fMH0XZ484u9OaOFgtjT+8Fuq8JBDZERlf21fropF7cLlQngs/dVUbn586slf8ooNc/fE
lHQ7wNy+uMXaoDoWTN7biyihTFlI331bge32105EZ/sQFs0SpRiMFYL+XVeIFkfVAPY87O2ZFaS4
dJvszPbcsRTh46v9dz3TM5dqOswC7eCBVwMYX8/RH7kBFDLWzTfNYabr2D+8TqNryjDmmLAdK9qN
NguPBrWzfXQjkbT7JSuXeRIj6aOp15m7LufN/e/CMxK/NogVrpI7VYZQBKY70//UApKix9E5xdLQ
2WU8kor/i48WS5xqQ3NNYKMltni0ldhSHuW+Q4Vyy7wrjyxg6UxL+rU//kGUdi0G3Zb5OCE5UVIu
2Jonv0hunXgx0Gz10wPZpLpQaW/Gyhpz6SgXl9txcLm+kl3T9e8pM19nL35IgWfzYrmcw/XJ3dzK
4x+c8+L5UzV9CHzO/FN6uRCCtd2IB4ZgGq9BchbG47sDCiyz2Hwgv/l0DDX1YULGIb6TwkCl55lc
u6+BaIut+5dynb51fkBj7rhJRnnEzGXE1XI7UupdWXTgseIUqR57H0u93ZqMjHYZsRcFC83Y6HeD
5fqrxFMhaQoIStt//TDF8mvFUjPay3wEcDm/QZfEPQK2Dr6ytCCCqSLPT/Ru5EIqxFdeKIeH9Tvw
oGXqxxJBvrNwWPBrk/ZuT5pVo1b3lvdiK5nO5hBTWPDK56DXfJzuVmQ44M+Nt3HDhJn0ZosTzs9D
yGogLVkDqmV31+9PKFng9Xq1PDlhNm4LUtel2w5a6v814XFPabz+eLQlEepuanBIbSYfkM0CVnsF
FT/UEo2qVLizyWl2AJKtO/EEmW/R4jylDgF7dseBH5hLYa+/Y101abeNwaibB3euNPuOI0/a1F4y
fcUBIbpz5Xq1y9PNWb15Vzf75h+vP5QwiG6ryzvVVMeEfP26JzLqE8qPCijiUUeLV+OlpZCIK8Cd
IFBG88BD8LXo6OJa2RiaZ9Qj81UUiR936LKwlfBpkz8iYca8sDYNL2RgufI7e875ilI7u605B3Y9
JNwDgiFBJGGq/xDOWYvlqoyPsg3QECNpUV3BLcWuxeFvGHis8QI+DRQYhk4n5SxdqddA2tT9uVSC
zHC5poQ3L7FO/0vTcj+MBnrtxmmohnL3p34XY/90hURjD18wPwfr0g3rcn/ThZ7ceyFt+9ASIsr8
WMIDmasc6cmPyMFx713pbWTGrk0QxnEpd1JHIBvy0qNUc7943eWvTqbWGoPD0PGCHlxstaAoL4kc
3m5fLA/gNBEj+bSQJhpW+ADsceJKrdrhvU73ZqPCAKJoVaOoKXeQmeeK5VrNbuTJHsDol5GgouRY
bGaoBJ0T2VxvHKHY9Nuo1m2gUAspIxbkuC22+HtXgSAb/62Ug0O4GDImsBPMvf8oZPw1aqGkQkDl
eumvvyB8qB1p8mFhEkARGQ8Stn6mU8ZxkOwBtsn3QZfn2+C1/JV1iy9nOg/M/O0aqPUW1g4QbgCp
pBuzG08Wa7nCagCXFE8rWqg0Awx/OHjftvm1/Gb/95+VdNyPU5Gj64i3YHrGS3iQZMLYzyvKLm9e
qEmDkqJUBZQMw6N9sluogKkf7OKfpRV00bro30L3ghDZm75fSDzDxNqLOZYvwNHvI9/z3sbMieEe
Bd8gFc8wvhbRembJdK4Y+ozcLTDO2m9rt89hNhuuETvp7iS+fKNuWVDd30l6aesaR/QDDlwPotaM
djzIZT5leqfuD4/+TRC3DVJc40T5h0wG34+ja0ViWKZZ5rvyfyxIBqDqz8PDVKtZoqGNKy/AVu6a
DMXBpDMUc/gCggK7gIAi5rVlisqN83MeQ4IEv9m/Vv6MuEO/tsizGKBbgaKKuLPph1CxnwOIqbFe
9E4qq9nkJvos6p3/pUsI0fRHsFwKOQoCCyGRI9Gt8yG9gaWUytrwr/oflz2odq5NmXuYqJC2Vchi
sXskgq7vaIsMvUu/m/zC5D3/IZ/48kzczQ8fxkgc6LA9tVjXqh3C7PEXO455j0bSUl9CdmhnPc6v
GSM5WjLGPOW1OhhRW/siqljH8He2GADpUGy3EHiSOHYogtkhLZ/QWMcq8M2I+L4doXIWUxGH7MYv
A0GWTyr/MBwEsaU3qwFmy+9oeOyrORKcRXQ97Gr6g765bJV4GUxHJggrOFtDdI83sJ99ozDcMtG0
JMrL+4SQfYM6FYnj3Y02D/uZKNWUfxbULC6KKT8pHFi2ZTJtVoAuWkFIyrBY2ev9xhDv/nCzb7lN
OVVvXg4EDltd7SdoMLgx53sAzGkHaCeZaq5U5xLAhzmixfhAzrLTtYqV8GJfu3f3dIKj21mqXjAZ
dRnIBy3lSBa5Z4u9RtpYBdzfQYVTnmDWOvPkTxXttuV3dUdlb8FyWo5jn818DmcyxusJjXVYWCe0
dd0WzfsfzHbHSVLogaENDh4QTwKO7s3mGxayIebqQTWH2RjfQK8jVhtf8AZSRbOTNs8SVhkQAcDz
5Okyhthmf+kgWvj9BLQF9+0LV3KJViK+cm7Eyn/Fy+K7HoAYIuBR9e8u2R//M6j4NOe3ePxCaP6N
GmwoiXVqNqMxDvIvs+zqIbNXbpa53oABa+jb2OGI3wxVmC936RevFLgTL/vAUGUbNSA0j1PzGwtB
d8chKG77Go4n8Ey1xWTPg08iF1Svh7KMYn8KM8M8sa7N//77dy2xyQEZYN25Pw6zMZYSaEtHw2hv
n0EN0fV1VaxyW++lRC83NfiaINF2zFemJHPvPZPCcP90FVckpaBs40D33L7NK9SlKhfoe+FedwT3
4y7ZMfLhXtqSC+2RzW32+vmL9Oo2ABbYlw8S54VMUP8ucqqsNl18FtkpY8xCkuh5t7hUIm8TQeFG
YBZU2BXbqT7v4jkta+vdOa6Kdcphbm+M9mfM9Gej/iWduHjb7TsP2nZlW/D4HmGiRedtjKdwAfvp
k0f3fYvi18N8PEwMzytCgtn5/a6i7ZrIugUnhL6HifOhORDvJNzd5hWn9+LMAB7jpDeAJHFoTOkX
LYGaqhu9PMtSVGqdvUAGGtzI6J7ICJSlnIxXn7wcwmF5wPUN8sTAYlZC4lecaWTn5mtmSRAISP25
NUzS2f0NGpp145LMdQKZMTQzJwDeAgnVx7D6Mmh6eCPVxjKiqz1UpxT1SmYxntYdq0kpYYr1lvJ/
eBGzLnwxrwx1Tkk40OgLJCYc6gb87MoXRuvdVAALSrva/69MP4Icb38VO3GXoPaNpCGWYekJtUG1
wbt7354NkDqR1s6G5vXMgihjhAO00uDTIgz9vDweflijnFW29ANEh2V2p6kXIeegTqrRCuWJsPak
PWJ/yyTIBNtU5WZ1tRCsv5sHlcLZAkmkySAI19R85n2rJPE79xBBYNM5v50vaMAD89oWicCv6YIj
o5ieFWgBxWOmv0/OWiPu8+GdFNc3OaeUFEQAPs5NZcd6bpgNZ2zX9G46gXdxCRBLGyv6dphRvsS3
3vALXjfaHOqy6UwCHxJA/oaKIEFWNc4qb8h5Du3PtYev8WKn3FOuDQOmwMEULqdK6BF3auGeKK0R
T6pA+ZyO+zGX0KiCO1BXMdm917A3alnoXUdPByZOH3zni1u9pPAVYJVd1FFH36GiZKtizn57dLt6
5yEmiKfF2n5xVLzmxXG7F+CLK3/28bMEFDuAqpPi00Wr1Nn1i7a2gkTdu81wMVVnRN0v6PA2yI4S
YMpK2Z2KrCBuj8aBhhQXS4tNiFVgJaroWgWIzMR+CYOanFL3WYj1WRjH+1IMAD5zWmTlR3XnVZI9
v29sXetUS/DxuKYoe9zB4DU5csyxt3SKOoRLvwZb3D2uB5+LZ97DiawHvGRnv2Ux8IVICpljFa4F
cNzRDO55WPIzWfnc/84ED1nAxi12r5YVTYMuwY+wVac1CddXcBuCjxKqj1wUgvIWqSQ8zgY02zuf
YlL07+COjaX5cjftxEV4sKjrfWKEVenuU6f2PEjxU9T4+FgTy7pu5XHOfD46InwMaWnwXNh56L0o
ji/0zp9gODkl1KIAy90H/bsIvrFm5pz8J0ua1X+ALAyw5se4iaWYBT0R9E3JyQWBcveKsq+WzFbL
0XyIzmk1LkIx0nfSBoyHepPReqCT6hkLDx+N/pb+b2ILocPlhCfROnD9wdo67DOCxevamR3zRmjs
5Jzy/bk5RLP/h9l4UZm9PRSxIX1JIYDCezI8jZrEbFiWVuch6EGZV0ZkB0JOCOXzNf+qYvF4xsOa
yotg75FEE/feqfwnGGen9U7idAVSQzze0O5p7X3Zh4XlY+Kv2VY3ja3CyR2+pb7IMZ+fbbwYju5s
WO3z/WBztzvc03Zr1ciWT2oAJ/Sgc92/GJNSqevrjv0MYcsgIAfkuYqPBlP1aOPDxsCQXI3/7C6O
hpbthn2ON4ELAtEBx7VrDqf0FGWKV2YYnGWYSd9Zob0aqMnyeXDvbEFRRmnfiIsU9D9BRBQ7MaYa
F2tvrsawqveIkM2FuDzbwCcnKP6xbSvuygpDjLnttkD4xNAVsi/i9AcIWQpbDMSk84ktlzdU8S5N
qR2RupkgRNCfnjvGQY53Q+sFFMT0vmgZJMxMNhz1pmOXMp1wwgmfAkBVDemdrLs2P3d04+9oVYZe
D8jq70PB7d18K0qgGTuCcbodNypu1d4zsw1fFQDFFCg8AdxitJ6PUs7V8kYF2OJV7NqMNIUUmDWk
PmHLhhLMRE2bjgU1/Wy2ZIFomnLqEudF5auHzeiMwvZpE8VkKhmNfscmmvGeT+cz3AMzf5vg62oG
WN6zUGhmDct6DjclfnANirVOE4tkgdCDdx/TbG+bi6wBz6zn1TkrCWB3KaAfrhjkvItgneVJFoaj
CyYJlTPH+qmLoZxyEFc/WB39ec1XvzR7ML/7TYtf12XU9GmQZOJKk7kiIpYCgnEe05QDqik+Uosi
jRdMQeGaaeXKWKJYu/f+pyXNbXYpB/K9LiaKHhGYR4GauqfajNNpG53RRBzlnK/2nhCg0+EcK5Q5
mWR2F2/TDgn1eDT7u3kcbae2OTiYh7ry95R/5IICLnMfVvLTzpMtjyrj5VumxKiW62T6AzwbrpLF
1izRRyWoW15nHl95bAycZGl/tDtN+oDCI0nEALzrrZJIzny3nidn0ctUc5WptOl7vWB8NWdNngXK
CTXL66B2F6K9tum9yea0etDOv3zll8vI2RA7jt68QM4UIWYmbnC/PGoTA+wCkkbBgOXJhDIiqGlq
LfmDmvn9XwkRmClJReekXcaI3E7Z1Lx7HvLmLjouvyTGijxxYSmSojXJbhTo70jyxEZhqjix3XGS
f58AHlyeDgrH8nd7BMekEh8Wgxj58vposnxYCmKS0IuQfbtkahrEN5dAUu1w1wlRYAM2Tw5DLw/2
oeFsGN0LdVo7+WE+E6QdJPvXkWU3cTfwaRLBq7W63kyRWt3zXJgRXBjTi8PzUzguxLYyRfs8GeH0
TiYujkm9UzIUbYTwgXOCiyPNPReTcTMUZHqNP8zpMemp/BKxCEwspeQUj7dJ4ebzfJRHJ91TL3LP
GIpyQtfdTBD7wadlR8XFfYirFCw9uGvlZRezM23Rygvelmpq2jIR/wsX5yAvN6+di/yemqCVS1I1
19B1mTDzicO+tFJGkbTrpKcpiQt7oKOtrO5xyVdPI95+io78vaGRFTHJErbcBQ2ttX8hhmg0efT5
Wjx5sF4o4TQxxRuRbnFbt4nIconkARczglDn3cFIAv/a5CNi8AwXtGbchbn8a9W55fJ0G9UutNM+
WeK+pzMcb+X97RrB6mM/6Vuj9tF/r3IZYWCwu3swQ0Uf40PO5FzBXGVJs2PsBdWjEayGyab0q197
jp89B84ocZLWl30pomVismecHM+fmsfDjoqYtdRrqCGNk3mw9qiq1JHstd9YxO/q3W+UhGigcdsa
V2sufgl+KaI4y6MJWSWr1lfAY0x3Gawxx4Er2vKV8CODiqa9u6S7Lp/QsvqW2rBcZ0FPaIi7hl3r
UH0uZBg+o6qO8jTp/azV5ifcB4LQnjvagUwAYD495N/Zqlpth0ql/baaBN9mgW1GDB63X5Bzhk9n
jkkbQBEEisbWnCZC0xdU4f8peuzLGZWbiuq4Aqroc0/pGfH0jOlPpyLYJsgmD7GKMZR5AWMD9buK
3dwIJLOSV+b5GIGVa3J2SusrJb6yv/FdvShbR6K6WwxZUQyweWHSBoPkBUAV2Y4gOSEM9WOWigtB
ir9DIkzOpjdtM6KPMmR8GWb5T0wVhWZWJfRVMyVqgtQsTSu2JX7t/X1XIVMsIeVcCSa5CeINgfAY
JnYQalnK8q2lYXg3z8a9kJOG0avcq5UnAr2HhCgu7ujXXPBZQtVQEirSDSyzYLtg4q6yX8LB2Ow+
G9UgQtjNWXqsvQv0uDep92R0M7+GlJyGLtJsMl6iluYEw5V17XEpt53Z0xmVz4Nm9WCsu+3qtoEK
WHW+jd3q8wK4cW0EnTGjNwOHVXxYQEFSBV1ABR8Id2E8HdpzgKPlO8HfXuo+28tx0snAIfdCkOt6
YuhHMBPEPygNBJJgrwSqRD+gEvvzTKB+fN9+YnKzmsnpTdvx+yehpbAANOox/nI2AZi/0zGVDqZ3
N774eNzGQCg6Kq3ySFWNrYQA5ChWrhtLZ0D8Sl13Qx/AMCL0Wob9ikFT97nus/mtjslohWq8PqhB
5xJL9klg7/9ZFHpj7h1gmQgZY9wbNYPVsy2AtJqHyu0fxnfl5QPi4mou0gooxAMzKa59Qbt6jc7C
R57Nt7fPunEBZJ0w3+DU6taJlHZmLstT1XeSuw+HI6VgUiKkAhVNy3kx2FtUT4O8toNjWlTW5Lc9
FTh2vDk07kWNlaUTc/759PUAUhBwgbRNaHt9Gg9wxHDGCcWJu5bwCHnq3rlPOi1BtiOtY1SHUqzI
1k8CCEVFNxKrYqZ2vPTTB2tSEX91qefP0upC9CpmTGd3y9m3UoS+jwOw8EAcx0JVUcg2WsoJ0TtQ
RY7XgNqys1iwgGbTV2Jv6cxUY1sw8mJ8yEBzn/GngmZL6eejwtaRetht6DE7G905H5hzI9tOEKBm
RAwHWrjCoqqymL9+M60Rn2LNbO5m8Z8GWntQI1CiABv172dWmd/jUs1yzTwEibSlwgTvicYKXmOc
Qsk033JUHqf0ep40b+J508EtPjGXyI3jroeziTx1tdGWmFjTNumHiyYXZogUJzty4Tu9YKjDYJu7
uCvnWsA0ZPuOePLO1hM5BNK6n2oexZIuPUJpgkVAu4jwxOBu839uoeuBkindR1mTCUUFJQPrgvVp
zmtL+SMBNmqhjaQ6jdqoVznvglo8BbhQl3nkV3RkDHR2cEUa7uE2ukflUFfLyF5TOPQ7Fj4t1vSE
IpAd8YzpeF1SSS9j+V7ymiBlR1HU/EE4L0liK64FLcSDtg/Z3mSiw4bKvuzCf0tfPcnvwApSjVTS
DA8RAuh+rbgSubGpTtIxO90teUC+vexqTAqUHQI6P9VI6Ocvr5ZHKolYE5o1UvXt2S1NVPdd0xxe
KUsvZ978sA9iUqW5umyzuv6Krl9JD15kkbqBNV0Bh5bSG6bCukK1PCNmFn/PLszjUvPU6nBRNzoY
vNmMoglHwxFHawsrv3/uLvKXu7dpYXbr6I+c9EJ4LbSu1Dam6plBR/214fWHodVqyukxwYYVSoHn
fg2ujttbXg46hmbDNjYs8GKqlZA5PmtifMMzSIpwZNmJ+fRs+16Yyvu9yYOJudyiD5BoNEtaGSML
e4aX22+eicGm8d9C3WfhgRKdkon5pSMwAHIy5MnUMxvbd3qhGM8M8+m95Qa7xaGAmLNDA+zU6Rb8
u80RMCoBdJJ1QeQAljcvoxFhLpabI4kL+gGoY7KgiHgTOT3fa8f23deSHUww1Nr8S8XowqrJP17z
UMdQnuIkz2pvpTrbx6g1tyInwQvvocx1dgHw7InZPEvsrXAVGGga5+oi6bQDs+tKg6nbwoBphNpS
an2OXRpF61ChHpMh+gwgYqCsh/TLJ0ySDaYhgLF8+FHDl7S5L/m/x367VSkavPHBjOS9U9CXByPx
fJCQA1Q/GF18GuMl5wtUPQ7OKqNqwAEaZaXHxHQ2EVlBhOIA+xy5apuJEVxDug44RoRgvLwAs40y
sg52qwAeMbCTlBwAqceXZdVZjNlIj6Yo0dW3yplxJELDso9AkCihjrXRa8McK/cU0Y1d77oAdXZv
gOl2z/hnpMMpz+V+3jXWn9Gmp3udXV50tUETlzq3hYo8H6yLo7yCzwS0NmcrqFs5Wjor+lZAh1B4
opmpWOPaJ1/oHZrpnw2oChBMD9jqdaJRlAoE/wUduNna3WfrgtZx6mfKSLCDJ46hYcCVsdARLEZW
bHRQwHSTW966it2bOEeoM9+BJs8QA0R1LS5JnYKWtrmFAf+ZOXXf93wn2Cj1d5W6ZxGehWTQJ2O1
UQLhhP7SHXga0LkLgtgTCQGbPEM7uBD3dzk/mK95W9Ga/FWuZRbyNph4LvnfwrBE6G4h2DDi0tQa
1vJUbvUKPL9WIK8/zENRbhzmjwqStLnaO/StAo2q/ge+BusJm4+qLhbo+CViQ7YomdI92M4mwnZm
E5s2eVmhaC0NxnNdtYYGT/1Mk+Oa1xHQIUzqE6t5Xw2aizTgn5xYXlv4rb8H7QyVsCC1RUaGM2+Z
VxNbVBV3rnvZ0dnMtyp3csuPeRFH+VeymaqQlPyb4xswtnK6q4+sE7BfVPLY8W9D7+2tOoxDqXyV
/El4mL0UGK7eWI6Sdm4qbccChTJInoFQpvT0DL5Lbekw98q0JM15XoL3iOeqqKspfc5WFMtGnx+b
s+xE8PnvROmG94QqAbiQfYYQTS+z7anKki7EP9y78h+QJRSQiaMrAhAEyZMJNziWaPWltlx+UeE1
U2HIaxwBOt9ZrffQdsU9htPM7vtYo6IBkqh6pinQCqh5DMT3OlYh6ojvvezCSCWkqp9FBds2/6E5
5lznJBVjE5LjiPInloePcleO+vPRlwNBuwX9dETY3Szqw/znCJiKRJZs80tQrUoPctq5KIZLTm6f
r94yzHalxtkcGHGsebBVs/me4buQxfIECzlc5nPIs8INdAxkfpWD/mjX6HjrBJ3dVBM3Fb5p2R9G
A4KmaK2oclwQ0Eb7iU+fBOrLvZEzs98o4ozam+AMXfe28rF1uemqX4LKqZEH1zCBPF12TBN1T9oF
U2+u8k91iBc5tVoXbEkepfoR8Q1/UT6YzJqyjRIw1WYp0pKKl08c573S8Ibqf8zZdqBV9g9773mP
rkuV1iOzEi3UbffkVxjsmQlVjSnxa+nxkT67wiisoTGyh6CvPUx5O9WhWbK98fldpKKJpxBSTvJA
EX1vAJIlHPl3OxXU2AmkXFYReI3nO9AYEEGRiwDH7zvl3ImKJOz/hwJuGdCgqKSNwqqydQaBp6YA
ZLy7xopAc2rBs9qC5+SGXwDqiJ8r1x4EqM9kRabBZmd4bhJWiMbNo+Dlq41VWVC8W5xzqMP9Od0Y
sTxCnZ3qtIrO2EGwL9AHyR4S/91AbboZQOsiM0vbx1ks62t5URR4LdbKL8QmNPPDJFJHeZyeiAvN
O1H67iTmiFfrwrLmHj94ksi05pQM6K+jNcS3wBATWNasK5ytWSvG/2/L8TFXMq2aAa005h5ta8tP
Rtt15Kkx/g02CDCEoyuNDt1tgH/AK1+0a3nk5+SDK7bENoPbAwGyIsHWimaKJWMrgnn1aiH9HILu
ATAQY98TDBX0H33IYvVPxmexcCSP4iBnLOI7U4fvwPcmR+t9h+Ip3lm2CoDptcbjUjzjt3UMfgxP
xtwuQ1GAlqaW9NY9B3sWIGzTruIGuJFUfj0omKFMDb+YHDDxe939/rgIccIBTKn2mZbmGhZb5/uG
C11fi0lfpDrYo89FYz+/wU5EaxrdXRzZ4XfqwoqS5iRg75OeWGFk9bj/vPdu8KRab95D1JsTS7Ch
eCwjCBRK3gDcxbGdKmuMcblnEtZyiuDEbSlG0fdpHufstBY1/45CeOKNWTlGrOeN6+WUENMSSRCq
rXI/YyG51z+gUQjtPumYw6JhH3AtpoVoSLqCH2pEpLUN9V4yb6IIdw73111gE2q0/hGJTu0twX1K
VsIn9pid+CuNrgW42FSsmIPrtWTgh3vnr0PAhDtlGc4y4gXkxKKkNEKGrdzpLCf3/yYLNeIiEY3U
L+PaStVNqXDf0L2Crne7/lgCV25hm4eubKX34c0bfIwqo5Eg+FniiOL4Lp8UocA6cyp5jK0E7BsK
XNUpsw4hhybLQkBo+Sh9CEBcJW6N8B8DsECGP3OxXEMOYhjTf3BXvoTo5jxGYmnfnbnRl+3ARdAY
2ICogPBAliWy99TSHBB4Tvfbwx9g+WANNaZamek8xp5YOaVdJS3S9yaYp/4kmYdiHijkFqrs6quR
qrlrY3Sjm7XoX0c2ZqbFiFJ5ay3H7B097Z1ASTHGP+aAnth1FDuwm08D8gNKmAgA9ci3t/HXUsP2
V00EF1ttYILRraZja/+rMlKJE7EYrncqYu1tl5Lkfctpg2V8v9fhpGXjeFV+pyO9xJoyMZETqhd5
7il4792nvYk9FtlufKlzFDDHzmfZIMbDgBRyK8eYDGK0Y8oTukys7xCBByR3MjVhTQ/E1OQPmaea
LVzdBH9qCzQu+sDD8rJMMeOiSlm2/6yxhMw5KKeQwyNOHVn8IZTlzotp8JM9fngQieTu1HEEsOMQ
EQwm/qI+Id42O7M8hlee6h2lZGY9sRqAKXuqumkKAlizkW/EBJJ0g5l+9946NZAXzM8yOWCHQZ4r
mIW1jkG4gCXDpEi39JDgmiBZevHPKAR9sOTAXMKvUiQkQYjVRSLL/sZPuXyxtB1RUegQrob10Otl
U7E5GPXhiFdKA+P1rSxcV7FRJPTXD0OfQeYH73vfqevvdNu5ySrsFiSi1yvJDF2LuPppGy6acnDc
CT6iuvNKajRfRkZVw3Mu++uGLL3fpT40EC6IiUWzUWjSbsOnC3VfQn9VrDs3jLeIt+yPXVvgLbH3
w6o5+cJKS+TXwkGZNAMYZWZN/bfGn6bNkNldxtqapMUkp9Hq0cjBDe6X6skx72jadz1xNG2E2M5T
uP52Q1DMDoyjrvqbBadKUZNasvkiWvLIZ+HhIn3knDC49rYUeOqVd8qRQ487xVwxHlWsjpN/tMiY
9Sa34OJsrQkNzOjT9+5wGbyIQv4iVxYKvYk7G//rqwaiF5BgoG8oEEE7jttpscwBq2bmxPJMjtzB
LHDWf8J3QOCIOgD1FuTlD3KjWiP89b3p3wrC97PVK1twlPvD4/hNhkH458IewL3QojoJZ4BG5YBM
1Snb/kVq2iRGq1PlTN9uRE+aVZJs5g/HuEW5BZL49tyLOrfxk+rYHdFVPnk6j8UF7z4fhUq0IiMV
6uJE9aWQ6FkO/5RiSLPUgoYY7F9U8EqGgyv3ru83Ez6NolGy08vgNvqAVOWWRSyROkHOhvbfIlxl
6DZAcQgpANg0By5Pw7sbcOhVgBCMpHDVh0ETcl/YrvcRSdV0t1d1NBKL1VrDciBovnhJR4r33DeR
HhudIA+xeZaILiMjpMPiceozWU5FNgyVit9L13TaW7/5EKhCmhYymfziTIhuX98IKZbPUsFweqlj
aXmYzIX/Dib+x1Eg0xfvibJ00alTyd2eY+85f2l7djSUnTj+BXeP5jlIUo4pDEXXUPCweQRTTNSs
Ai0yfYm+jM1MW6yghKAVBHzyHTTPat6LGz7FX1wP06yHAv2AQZ7grcs1a1wzbOQR1rKBEuGPEhpG
kWf4+TdDRV3r4FInQN+015Ip377XX1Rm/PQ9pNQA5nYWp5ZEiE7NSEbNMUPX9XHO6YrgylgLInrG
GfeWQgQxpm1ldN0NmWfaQJoq4q7noG9DxzUlwC2NV3q1g87IFkuEmUX7qRxAYdqnRQA9AAs7locg
5RSac63+rOArbIOjZAZhy2U5CT798MTbiLBob2dN5FbKBJbmiPm3X5Jgkhrx5aaD1hkycujEtqrM
65fwEX3yIuEyrBfQOaqYNvMgR1u6lwAXgYeh7gSKQSod400i0ZYu22fo506FbhmHmM3O3mG6cYP5
Fflz9lF4Ob7OuJ9SkF321nBo2DS4DNIHJjrTy4FF4cEvTHtoPfxuRZgLvZuG1myqXT9K1N8t1Ea6
HQOkJcDPmzrOyHpA981T7dSlmAMlBSU5nrhaJQSvK8xeHC3kFerW96abltkXFSOvhY93Gh5vZq0p
skZHjq8K8nR0BUydQXMawoFQYdQfVhxBWsWeUFf+WzeDf2tqN7DWllIv6YrT8N+IaZodwLhVSNF0
cRESBkLp1teui1BIgKrdMzGRY+1dPzOyBaH9KioQ0iOVo+7sib43vjTcjdwq2ePp8AP8Zw4hv9Ux
q9P0ybixpbnkKdgSDZ1ytkCRTWI8rXMji2tOzxAdj+59JXkAJ5zJSQQxyqHl4ARDBMDkbWQv0uuW
pDAw6Xd/94KAGrKAGO4Zpnv0Vkp2scqkEYXc3fHULUYpIeA6mf3GBi02B/Qo8ZIUn9PddHJo1el/
Rd456ddCpXUKpgkGNEmkjXoj+6YSBROVz6AtE+MQ7tSmS/MsS4NCpKxQpsWaMM9aqohXqj8/mexn
o7h5ZlRO35Za/+W5njfeAHGShjyukNRQ1XgBWv7HGRttfZjkeR8UCOv5CRf8y+TFvV+NFRUDbrnC
o2clgkpDi4CPpqP56YvEkxeP2ulP8V52MLvDW2s4A1WNuyCiGQvSF8lfhcsjdCF+sYF6XYWpaE25
h2S0uflEXxlAkCFA2VjG3+IpjDbi9hljInbSGwXTD5AUlPnxKEEVr0UjOUqNpnVtG+Puq7GmREZm
puCTQNEm7U2u8/mD6w0xMkcYiY4/1JMa3+kwKZ/qRksj/gBYeRjCOxMLFr/D/QjTb40eI3vpsZqf
mgZdMc8wVcoHds9OOGsA/cIg/QuMD8RPgwtI5Q3xhFkhYxpia0VBkMeAUC6IBq8HV7HXG2j+KAAf
BhGFCpwWNJFp3UnMQC4uq0y4d9EJ65JT9Q61naLjeF9yd1pO4SMQd0qM9OtiImEk0th8FhW6c386
mfMqOcDRANM1n5IvRO+cXfhUYgMdDuwJey8VeV8OjM5KvMaElu9KGJOioicD8Yc6IlfWOSOXJdVw
hxUEYRFnufseBlDWKu3Ay6aelsSpaM+9v+dfJ2HoXyFc+rPBZw1sscoqc5xVEPtK24vFwmogrFSC
PLsH2uP51MGub06qGf8bHWLQCVkT/qNLNNHuvhYw0PcQUWPrIKMr33gZ6S53NUvCSc4aJ3Cl1jzE
/na6bNI8i/TN9yqsg40CbPwdtw5s725UxEM/cqE3iHGM38y816GkcE2Hrmy1UniHD0wCJSQjUs4d
zAHTzuSK9O43qsDYTQ161b5O17wmQFCfYAweJatJZOjJiVg19EjF5470XU2iToQ5fefsVsb0rMob
qkMSyfFAdDUeQeOehlCB7b1ehHE1h3zbOCESmGX6GGHgKxZZeFzGUnZXYnWMdmmRL0M6yHe9Q9Mc
wrW0KBeymCGsn77FO3Xg6jiLdA3wE9/asCKFzlnU+ityb5y1tySVwLBTpk/xdFfZCJfHkl3YvH2J
8Om6ZPypr76b1nmRr6Y1f+Myb1yXFUveUjcEpggfd/c/p5QSZIGSrr0lMEMTe6ebn0vN0LxrdZr+
tyKVaj12ZGuAPqMQ7ddeJ2WuLpjyiVT4nGyeh8fST+sqbMW5ctgQ87kS74L//IY/fzCn/qGAklX2
6ZGgz1wmKZxGlG5Ujju6l6sU8BEECL7tMNJ37BPhsWDMgPgUAmek6R6kMrGSLQ31JipR44KTTqHR
xU/V3ctPTfPzY94H7f46eUcP6G5QbrvUjRfSuo+/p4h77HbycikoVh2AqonpGrGEFZILKfYhF2gt
dwjV08L4qecmf4ZakBTO8Kh0Subsxm3mOvDR1MhXraHNv5Y8NnCDOfv+dxlvNOAVCDxO4Zm6nyqF
IFixM0Po6mF6zQMKUc53FNemwejyuz9Vmi2qa3yLPiuh7ZnYBzkXh2goOlzDb+wHUp1Dx3t44Cdm
aTxBJdLlgCcuB4bm98xTzPCf/smCc5m8c7p3lzNg45bTJglphYTqecoqA++KXx7VFQlAAz86ZK52
qr/dIaOvUQcDUQI39H2X+9AoC/Y7hgfRME9PFNw2m7yHc6Gp0SK30LF/gFm3O42KtKTHwxKOHAi8
tV1/EwiqLkKqsS4rlfhEHSiATGja3VGRMgb5ZeBI6cuoWq5l6Iwemi6ePQKpyB6jIBP+iE8Kw2iz
1XUpqj63N/4Gu74KIrLwlsHmTEyQdCfbIxGOUb3NysGafKI25HLhjlrDQ033KaGL3VJ9jRiLuier
EjepviCcl+Brf+iy0Ihx9u05enh4igj8z4s8KOxCoIxALk+rIY5Hjh87LAOC5B53O3hf4wLIwpVG
FuJuPuTmhN+oGuhj5mo82SpSfE9m1ijtznXYu3d1vpCRMGpR2Tt+MYLOYhtE+Ip+eeKY7c8SPDi/
wb6I6qRxbZRjMbR4DJpDh7dDaZeVsqVsd7vOMNy0gbFD9VelpY6RCncy2wKGm66AeKbw7TZedUkT
ts2v91xTNp4Jo1pCr6tavwji19HOv10tGYJTJqTtpuXyxaXC2Hq6t0ch1WubgiItApgU9tziwzNM
6HAPioAsvTPPhDGJ20HLMYs1ntZv3VfO7QmAMgArC4sdzhmsb6Qb3yVMV30mRdn2MbJi6MY168P5
bjf+OCviKGM03HA03CRHveunlf/6qLSuUccmZRuZvo8GVmL9V4aj8bU3t0eoxFcEVnvVcYEyQUZm
K4d6YxINEkZjKDe4QY2ZYY5lvyqESup/z1vVRGLNTjhHPCX482iPuV3Yghsh4+H2sVJIhJ8c2gHc
tZ+47mV/NXf2ryU36NXqKzxB91fukfLiS4g2zQeJB9uOuHI3Y6QF+qFXzg5s2MNTocLB88HhQ4+b
l3/q8DciJhO0yirqnSKyc55q/x4FQUk5bKjP3OiF12LJeGcIgxrfBnIdxs+91RcK6wMJAED3yPHE
BNT1zEHHRtwkaHSKywwj4SQz+Qj5XH+nTzyzwqOIeb5xTNoiDuL9R7OYb6aJh8sSlIGahSos9Dtu
uZKxmFb3dbG3XZoD/5tA7HVvjCtrXzzRam+7DXppGEcZgstgzyfrGhlivqsS/S7gR5TVJYFz1ILk
bP93ZKqq/te6/05HK/375Yf1nWhsT8kHM1ZXWMKbxabk/O/1MnL1dbawKAG8kk7NHOJ8xb5kNGQu
BRYPcQer6k8BHgADcv2aMZIqoYyY0b4rXY98M74biH41FrRweZ3ChhESPu5PbQpFvGUsphen7WR3
wFI/pZ9CruDvzvmtJiBaTGx26hP+LOYaPD+PC77fEn9GxRS43CCKPdK+K85CBFb/Mtmq9heWEzm0
jT0DGMEI7neajGukPeWIw1alhmTfOXlF7KPQMVqaM7G/Sc4FdhLia6sLA1oEGf0MT+RzoM+hu2fI
sZuYTLQ9ykI+Y8zODXCVik9WL47Z+vSGIqA7qjXlgSMbE58WfkH4NfSDY3I8wm3X/bnKQyFIaIQ3
O/jlmAtocjM5h/PJM/plMFQXdU7vdHBeoKP5iiM8Qm2HBpQ0bGPiN8I93k83A4nG1xqrytIm7oGP
kbwVD1gteD+q1l4hrnmMRO2QmXYt35qA1teohv4c1iHBdTCYx3hwKGLaPDYd80mM/yM4eyEqWHJo
tmli1pr9EvQ2w4c+SpivCyHbJ2EVwe0RPmyjGYfn2aQy0jXXjYGoRn1OScHSqZNWaijBgBN8oPgi
0GMyEbqKIPgvOGSMNfK7EpDCL/7ZE7HWAB5Rwkpk61OcKlyvfR0hsmHSmdpOVj+TF/KLWIjx9iSW
hUSv2mhAaEF82TQuY0Nfjdt8Uae1NvVN9SISRZfCaFjgeot3Rrn+USsRTl7MX+WvF6Y0NPN6Q9KR
KwmLp652VeCb55Cxo7UhPUp2DTkJq7kf9JkRJjP+XngNAXHUA+16UXHxj8QqBU7Yt0aHkPijFZEp
tX/N6YJtUXmamYHRVDoHZAy1LQHL9VDCqNnDrRlk1agMbV8X/0d1saxe3y6aFrt5M/sKyLuRfVVs
Y0gTnvwcXv5bH/DxLHg9aUQrduY5bajYZPXuXfgEbLMLw124xa88Du77aibNGQDUeNx7Mc8VVe+x
ERTYJPz0xZ63p1jqyvIU1mQpqmCTCfVcYHPDE6MCu5lW8+4gvOWuOVRzKwivNghoPj6KfbAMKFaQ
Dw1b/oRgHLe4DxFty2Q7gJ4297CPreBpPMYXnNHqS7Achd+7HOQGS973/aEO555sjG5TU/Jv5YBa
63PyGqnfPGnIodrLwZ0ybxnuFeZA7wNXy9tnXvi26bbaKcr0AKcWniU3qKO6ep7aUI3VgTZfU0cW
eifOgU0R3hVh/QBZNIMLXyuIaYxQvL91ObfiCJXzbrzZkIMClS52Aw1DyL5tyJsHUPZ6ATU2XJY1
fzrIGD/iXMUgyAz1KKc57tfB1Cz012aDD5JkPJwGz/y/Wt8QRe+2H3klu3AsbXwMvWQoS9Ro/1Zl
2Dq/dazNM6M6txGO33GO3o1tXFpfwAUvMsXpRJ+tloiGLZYrJ0JUbjLjzfdQvo1tRtaBzMhmYHKg
kxmSbL3OMiG2e0H4p+mZtnf+zp3a3Dp48Rpa/8XRR3dPknMx8FvoEm22JTZuCEqSmY+FOuLdnvA7
rNWeSolj49482DYgfXDcPZmnnqHupKtVxPLfKc9093YbQCz+fo4RrsBue3DZqHq6/M7YMEHUDD21
hyINh5MBR74ZH1JgkpTx2gkTczzTsmdaCGPut8er8ExfspnczuLRARBxPIkXo2jy8YVAiaVy2u2z
6LxdX6y3BfMMmipxydoH8VbL86t61oMLU1LsVExl0Cf2zTuVi/t1c+dj269rM/GlE33Ta6Cet1Uq
MLCd2JCiLcfarJWmDcy51hxuG6dwVJ/a5NwH2iKbwxHWB7cuWNKqfHzGGYYNqF7p0R0KVH887AU3
n3hgfnjzNyiVLxmY8W6GgP/qmMIk0WRm+tzP50kMYDkcs0dID1tXV4vc0uvWiXYS/9Uhse+WKq0W
jvMfNTOzxoDacaLlrtDgT9tm/7VF3Nksh0wB7JDkGvqM8txuFiR5Rd9z9CQDHzyAigMxUWjxZo/O
GIXOCYocEpo0KkGwIfGj7He3ETSJz0SKCBrlQHEAiAU9FAo/6tU2DNEGawbX6VOXNcPwIrdRxzYO
Zi40KVBlSrVEGH9goxKUzZ9dwh/4BpgFoRwqwa+cqs98rtMfwktlOPjaocdS3gdThytGJgeMcW7k
kSIOr2m+QyA/zNt0B1YL4JdQqXC3VQiLLmLaL9kI1o3SAXQYdbtv0aj9ArJGaocVH+7zaAGGf+8+
J/EuXWwAtwNMpLpQQZaxZ5wM3YOdEGGD1V6Khkp7ApixrxXKsW8RPUqHkx2q2SKFgKjuIqlNl0Nr
/3aPrN5tGHJgnjI5GHRG3M0UCdJdnFEzbnVigTSr14SQwm0KDvPe18KrO0Lc3i1PQ9cqwNe5hFf3
pfZO2lqr522rt9vbtYBTJmrBPpNxD6zY0+E2myip8/PPUY/w31AoPKWmqKr6f/HMJKOqQdhz8Qs/
WY2X9ee0qXIaB6YYf5ygWoLep0DCwfXj4Tyl5ddecVWKaFLDT9WoywQ57CvoBn1ZPW3djpJNJJdk
8EYeQdDoGO/jDiBHp3oBLwQcLcfuv7wGgVKyfYwoHQHqsRdKnTtNZoniVXt4u2F5Yj2o+GBit1sB
SVr6KYmKYi720mZW13IIa1B6RfK3FGOeuhWv9rHFPv3PcLkRcfwacaTpVTfHpHyoMUfTnN/kzJF+
hW6A4tnuOd3Gg25Bn2mJpQj9BAOqk1pnEKqZpG7W95IHCIfT4PAPB+2FONP5sQo9W/Ys2pi4AaTw
rf6sRSFKdUSd2SRkA3c4v2uqfQvpOgfOodVDv0uAxIAAclQqNA3NehQ1nxzVEZmwvzww0WyQXMwk
zT6t/Il8azR4ZpsNuAikRvQGa/KYlOOLQmfZrxhUiJYSTQsAmeqRt91Xji3ome8gfjf6c8FLZYqy
7SsDrAz7s14EfYTSC0mlC8Tc6C+A/sRRYuhIUbnbSwp3WgJPtjlXKOUiwvAAOI3rPzaXqMetcNlJ
SooOWx30u3xhi+izSbddpUnvtBNotDwivukQAC0oCqYa1zkBhheIHujym1MyYMgrXMiZhgQHj0si
cY+JlG4xeCsew6+uEVbenEsjg7VSPHtqe0Hui1kcdsQAJVPvogtQaOh+3jpGi6i02GeiGY8zjzou
AedkYGGq1UbPhY3HQ362u/3SOqX0+zoCwTajM2SSc8Sj8+Z9Zs/JHt3xLKF83qAq8fxN4tm/BYvM
3FoEZrRmgFfuNQYOFNDCYiKTkf9Vgf/FJ98euzLC9Ma7sMtoKeVa6bJW1Rq/IpVtiVLaXokZxPSE
i2Jll0F5dpHF14bbcMZ6PgpnQno+w5j1UdWGlbbq166nx5xuMkAZyFoExYM90QQmB7ktKai6bbnX
wA1Ga63nuMboqhE40eaaoPcbdDCgaXnPDfO20VFcJgjd/f2GvQ/zMgPt8jhkc0N69dlc/V4PP3TP
s732hjiEid5RbCxVaDzlfXA1Wbvw5P7xuZwuluA4AUEYnVZyZsZuMPvqfCFn9my00UVqzY/fFPa1
SqvesAhkDjcNwSCwFtRbTWpA56mckG9Py8jFmLn8z3iUxszu5TGdwjZMEDrpwcZIJps+lWBel+/F
0RZNqHSxcPflqVz+680ISuD1NQbBnNzmPmJ10oNFEfev0JHZs4PvRbDHF9ALnBg0YvNczK3LWDRK
yAb022YyKoc8Dg4MOc4hHEEMe16aWaEH5coFWXTbp8mHGhdLEXAq81sRUxLpvLNlwmeayMqxjxsc
ur1We52ZTVY0yhFcawTmsWESL8U1racET9dKj9UA6ctl3IRyrLOOcHgOZ4Zem8fImp0j6mHjoiNY
bbgjQaTaLBVzqX48sc4l7Ud0908F938KP+LSstm5wMJXZ0e1aR8dNpEYZpjTPYRijX2xpJhVMhXU
AFG2M5QJ4xI+1xkSASGOk8NyDzx46SQrnzOHqFHsxAZoqp2/uNdLM0r7AoxORmaNT9aQzqxLwQ8Q
HmifVWR16NAw5TsdNCZ2D4/7ER9ZYUmC54L08kR6aD9D7QVzhPjahT3dOAsZy4x3x88/WejXQ1aL
BvXHI9F+RtxBLGBfvC9TS2EotF97YvnMT5VAAo24C/bIWIkoGrSseMbVnjuD1aSeIijT624iJNWA
rIkOSyzZh1JqwaEYRbL3DtoZFLufeDwIFhbXe+OtBWQoqE0mHssBCeLxKVgTy2WpAcNY6CZDCax6
po/e0w87oOC1KIzeQBZ/18YMb3KBHBA9MnpPg1OysVH+s0XPyou9nQpukI1ZMre7kLOEgl6rrpfT
41IEIlmJyXbli5S7y9ZfZ0FOI+S8yNN6rg95XPzB3y3LfcVNdDy5lY6+2TDKK/o7DhPKgWx6MwkS
DLr/QQ9T9BcREbLht4ZF7kGK/BM5vxV173sVy5uFDxNiDwvyqv9rbomm/oG8LAIPwxZzdzh3Pt9p
wtjck2Jr0z2pi5yILs5dS/E7Oh9yfJh859jP83rRWbU7xGAYBMpv0zMzwIdSFUIwxjH8dJj7fziL
3uSHJQhhFgSi4IBINGz3+UH2EqIv14p1ZsAJHkBkaW5IX4QBeoiHVZKzD9GNkjvwpJMNq3Gdoi2r
4th575DIu1DVPp8TSYT4uby10fKX+IoUiiIM0xC5uSU+uWbdK06j2Yw7UbdgOuhyBq8VmhYMIbmP
oCKdGO0dSqa0Oh1AVNnJyznCxle2p1G9bMfvom3gbH0MphmE7YW8Ej85cSMkJxUbN0ubkf3aX6f0
9PRW62xbTQegTHSZoQI86p6EBWqj99yi0/vajBk8f4c4t5DA41u0OsIcAJOZ1DmvyTANov5sxokx
/98myP9KsxGiGFRLpyKBFlxZS0yBLEoxTaiYP3FChm03kL0joPqQd/EzcVCYGUGElCW8PgmXwcIj
ezOXs8h7UFeMrS2HdwlHVttOAIEVr5okIlDdIoHzIYoo22ChKrcn2XIsWEcK7wh/4WLKf/BoIEKF
zxuC3QGLKH5XOAQ6rotlihPGW8S9sIbhoEJ6h0VA1CT566DKqkBVFsfEfCaPg3vXzc9/G9pUar+k
goH7Z66A9MwE3mUSIyhWjImvv14G+D8KjO4CSJuoc4wOEj1M53KyXnbvRvdAd6FXJTzt0mJbHtMC
CzZQ1hfHaWIYUhC/zBYr2hMMxMvMiiO95zg646BhGlBJaRZDj7sAgGcjgmIIpXjWY09uzAHvq83m
HVUtv06uKis+u8crLqTUvB77lpEQ7cv4PCgNsG1gxMvbBENNDyJMZQ8zi7d49C2J0OeRel+U6hh+
s8T8j+XhWUu/YOscDkWQuXki4mED+pbcL+hZFUuH3Q1LpMtC6UoaeSQ2MSs8ecgsGK6foltgRaY0
WEuL9/Ls3L984VIw4uSAJSyRA8Rw7+r7ZsGoLT9CPlVhEsHykiP8m0eadOzwiqQPuNTy/q2c6Iqj
XzKAqO0PbSLSAwiGk+FFGjvJH5bZce8zaLhAW48L9nzHJeNiTq/znd4GizTfiFU64WgpT7A47lMD
r8upMGPYnzyV1AR/XxyfOAsFVT6Lx6Q5xybowz8ujLSc6CG63eUHXoBMCaKhbmk0GqNtAIM/yEeM
mFHiuVAB5nmncCu4TzFYkrgggFxZegwj4mqRC5n5c6E3kYyuJ/K+VLweiMR5L2ogo9URbuenBBFf
X1r+Pv2KEEviyf8v50L0p0RO3Z9nPbNmeWjUZ4zlpXLsnb9FXIFg56JBFEPEAGbR1h/rNRlxdsBI
sgWwFq6n0AKVvmXPvKjLzCvMY7uR+XSDY0X/8Aunrph/nDAZ0JvB+88FRU3mpuCFx6/HtAb87Cjh
F/EZ45xOdUX4khGnKYnPUcly9D69+9w5XcdHTThLbMhnYLzhhXPsjV1lwCFXj2iIbtYH2Ft+e/NB
EmZ4wDTvsTgphXnDVWCfZf9S6PD2978ZP5tCdRwxlQo+KIPwKw1cN+wnFgAqRsbyEFEhr164W0Dw
fy1NDBtm1DNhlZIc+ZBmhFpmINQ4pDXA0/urIhbyW45kNxkk2nmbhu0GI0E+rPc3iOwVNEJ23/b1
Z9pzRU8NCh9iEKenFwRAjVIZNE9jIHjI6byUpYJ5T3NQcFyacYW1aXXZqYUqouu2ekar3PLbkEUV
JHaQuhBzsoA5OwdKaqjx+Q1KHozj3j8cIrlEAygVmDTGieZAkQgHd6PrDHuqmPibmGBmFwo15BCY
AhAcirrLI/PApC0zNF4HHeeiCVYBtzlIHUDzNVuuQVEOsUfaQXIo+R01DAVsS3l6AVfyvuNQgsSq
IeYS4Z417Q+8VwFW3rospQW1jdU/MLPs49MPAMHDVv/JXYbGDbOnwpOgjQJUpCJcePVDEFh50LTj
j/8AsGA8zsh7yV2JRCv9lsSQY+l49XWN6HljMPgIYOTCPYYcIjbFAZUnn5ff2z4bxA1/Sdfnduj1
GwDAP/SwPmtzf0aoFO9Ncrg8ANzyDVkL0Kiuq+lzVNy4LUHFlVroVETpe9NleICTEV1Bbvr9+s1D
d0jMtuNKbP1Ik3IZ8iB5+KD9w95dB3M470ECDv2/s8yaAlTF6kK8bolUPQV71BT9NAZJsMaddPCD
hpJbCSrUZfWQUO2QmF2RmFLBwfy8y0sM0IVcSq7ZxNOavWMUdbbgoq2XruPDzGUFTya+VkX9gwdg
YFqRTHXREUkU3RP2y84rUUHMjUFYe/lNrjzSjDlFKrYXBYYy7SHiypO6vwQ68IYRNwrCZch54px+
FMz2V4yU0VQfa+ieeAaSrYQE6K8F7o5F3G37ynn+kzkg9woa2JlyGx67XdH8amFolC3ThAkkyab2
8gZnNKRznt/Toqo1W/NQogTtHfQBLEOaES0YoBNtyB2m/1HhCsDv8sfAtpIMBeSOEt05kHOIkAMx
nRC+5v2w6a/hvTcQHv/mjdtiI8DnzQiJk8OtgEJPh5iOieJdZUp7fm36Zfuzm+IAG+lnDU9fN1bd
Bug0rHbUWLVvIGi4RYUSJecIqQjg88wMZ7kRNkoKb/LkBo53Em7dgSj4ALF8BuxWQ6VyB9V/U3Sn
ad+v0YRxOGid6CJw9MxZg6Xlr7cYodGH/h/VJCKMjrJLS9DtjvtvBTkDU9T40pmvKBlHzFitzzcX
LKiOLeqRZUi5kgpOOtTnHc4J5lopaPhiYM5cV872eY7L9QHNbx+srzBOP7PePtuumgfjL9udxL5z
Go0FS4NDKZtJ7QhjwgaDFj2hAZqyyPmoAW/OoF5Hs0OdwcF8bq3Fu6ozppaigJ8T7Flf5MP3cKrf
0PUrJarrOhPQzxX/x/PNvoORkWNcJ35a4yqVeVP1s3AWHVPusldzbREZMQCAwazn5TeDQPoub9ez
vSldXBA9PbzzmkeEXN4Zml8AKt0i1ZTAgzGOxx5RmlclKhkqKcdyhb1vaFi9HAWhux2S6+yYchwg
pKgv8IEpkVbjQc58ZAy2jGy4XTgV3jhodmP6xU84AjKvexlZr8fCyD9iWKfwMmhn/jxsweJnlgPG
igmxA0y57qs1IanBwICD/0oawqfA9E4q40+UMlJkrGsz6/8UGwvLSBqTBra/A3XpuvBxNXcnvvMB
dKFX5LyFFg2EntrFo4egp2d2GZRSEBeLyD8NJll5UiimqX9JhYeuJE75jhTu4mY6qCTi6Vrdyv+A
adgPKbe3Drpdy0TgPCLQq2nj9cCA2ZoV9y5Uw2iW8Z1QHxlbiQgta/h89UIcDlqE9e8lmJqmhK8/
PvUhMYAG74wlZXeapm/blFfHHv0HePz+sebCCFEK7LK6psOr209zoDoswwvHzkx9GOcnXBRvshxp
UEAUHXuetQn+Hz2207BDgIDH7CYEz43NCmylS32ImKdzqmeq9ONIGCvTMrXxRtttoKPbwh+c1ePq
76sHNiUO4RJAac7sNrq7+p3OUBXZhJuCUTE1XSzS0n5bNaRXxknv/sz6/dbihvQtW0aZIhQ0PwOv
7z2GrU50/ng+ND65AZpCgKYLhUJvYhnRZf76VG4LkysYhfX2fhC9w7kR7Xv0YZMTGH8pDE0Jzixn
WSoCFDUFjwpfkz+Eb42fWh/ytU7Ihs/mzqrkPwzD2O5rTmt1mHEehlUlXRs2YkqxBJ1YUddUlFQ+
TF4sGZzXknm/JV3GVQif7d5l3tKIPHMbcGyYbDK9WrbzDo4qHHtsblGD72KGHvBLxZmYOdpiBJXy
YoGLoPVVpvNRqQ8Gw3IxK6YLQg7sp8N+Da6TLWaaJOjHuXohrpAvEpZ/Ve0kEwYgjAPALnnKfpyT
8crmJPssPanmCLq5LhKUR996BckdrYZuxPQyeZBhKuATgFH6v6h2qDxBCjSDgj6bRjorYhVvhHPY
MLDhBbb8+yX4le42NJZKl9+p7QxAVlNXsDFMg2xA8Hgb9KcBY0fpBkCnNy97syrpzW35BDUsNfm6
KzU3W3iPMwZUwGVEroofVbWf6tb+KmWzKz3TZ/PK0hYuh8Hrc1q1vjanpbEwTbr9/quADls07TgA
KwWMgGkzJuJu7q3cP7eP7j3/GZV93vwI4ywZHxz5ddn9pUDeWV+nYmjllmLfP8c/eKDhIQsvnDEM
pVY15I7K51npMnppWkL9YR18BbFlv6UURY+m8l9d2+WHr3+OWVNncivhA8IUzoVoWZrmgr4loS9A
yGiZ/s2fOW6N7dzM0d6Qg2QDPJ4ItyOpejqdSmH+VZZ9tpG9yGSOc/I8DCSAIStLQ/SmvjkNIZFR
b1S+U9t1JpFKjkvF3TidLisUlz3+UV4oNvPj6ueKgk+hxVM1IoMhAZ3uYvSgy5r5usG+rCodlkky
eU3fXaLz4LWw3F1/9DEhtdETLKl3DEZmce+waDTvWcnTSR/xN3vNApzbAaw7jZu//16eOI5+RIky
HsT100geehtpgoZqeA5BoFdTSbo8mHKnd7Q9vZ5T4AmcCUcafssmimyBRBpOd219Ev6X5Gs4NjF+
fKHIuylwcQOKeqv+8TEevn40R0E/uRUs1GoopCjPCU85/d0sh15daWKUJ5XoESj6Ql6oClb+/x4G
dzw3HqUZyK7zT4nK+rhN74r2S+ngrYBL4NMvzp+1OERjFV1i7kh8uqN4N/sC1pb6Qhhk0tvEqSiG
KpkcwxJ4IK6SUF/ds2+lTdDz2fM7wG5n1rvyG3706mciOoFO9rxt5t/NzZpTUg/1sC3QSLHM44DV
QJKdnR7el25oxs9gjZrUsLAL+LpmIDu5ySRinK2LswcZfTzssrRCHR1C4RMeLODhxBhLD7DoO3Vg
u84LDJA0HphpOS2W6I/X1eJtAgkFaPClDMMF/o9pNO4+uoptxqR3TLtFaYK9J4wvW0bhyjcs+ydu
6QmUn5eEo2uG5tUI/WHQgMyR84LAFIb42+ircvnn3M7SQ4/uV2oP9zNrSJw/IiDeJmzLjqyJ9OXU
wiPWydIZgaBShuF8UEruqO7mXNtVHnF41e2xAfQbioSBjrSNlDH5eFDSI/1uHw3NES7wfyAYcW/6
IXmsG0rpJBIA09WIwZBf89Ehml3ncW266QDaIWAY6B7Du5Mgai7p/EJZ7V05huW4XK0j7wm/cQG3
cGHjTY0ilmShk78CNwefA/yEtwqo6wQ43+zBGxwsFngyDnBJhb3FmeINlHRTK2JGoys6nPCqIWJ3
+gNYu7ZMyZ5bzoFN7X842F0hqPbRHEyXGTigyJDrQBp8xcSu0XqRt7ap3OG0GjLAXtAxyYyPD17A
EpGbnXSpx6FvtvGkfBbSlsBCPbPL7/2xTl1IWQe62XXModIdJPoTqUxvIbYsrea+jYcyIV6jW28p
Qqqzhp4MIU2dNdOiCUDeD+aRwQaAoBpm6nPJn+mzp89j8xXF0KL+ZqrJ0YC6jRSSkr/RjtdbaByD
LkZ20XSasBraDf8sPyL2kckYbw12Ef+SPxVKBHeXbjE/GkB/9Lcwq24lmZAJns8cFRSGJYCg2RVT
80iFQuQP7nAbHQ8iA/TI9AYqrcX0Xl5AtFWRZr7//OOLiX5P2QVRR8dKgY87d/NW/RNtAc5guC8a
Bdt+iLbpOStOwfRlFj/YsUCJ/Xlui5orD7A6NdDhrZsnodja8AxGwkxp7pZwq9mFSHwxqm8ufs5f
MG2r3H9No6q5ssPHtwVfwk2GCJtgIBj8aUZf6KGQIHIA5b37M7/2k4w6WA2x945oVzf5nJ7q6e8N
flEp8qkvaoFtKIAactD00bcC3VuxOAx+nIXMIr0yLyd6KdAjLa/Ewb0WVXhAQN/xRxSd04D581uA
LfMkhJLfHcsUUg845Cg+PKLB/sA0WTWk9vdOpzgN0hbDHbisDMnuc+vB9ThrEYPKVl2lqEj/BFPl
RLBOiWwrDDdwjsvcBzG3b0y3v0T1NL2Hj5aHtqqH4tM74aBFBc3mvMmEuNOyxCFus8BUAzZsftCm
H3gZ7sr5nbtC0pM/kpXtx7EER9NkikWK//CMRjCwIjEFniNZP5Zq1BQKDJWERh+688HsCegpP4J1
VtrQ18UcDe+z8F33XnN1YlvBMalojUvwQP8nH5bCuui+trOsd2OqHlKHNjco66fiL0dQSLdxj8tj
Z022LtaAp3Xv9rv9jvnGuRGYwbjG/WnQR5NY1JUCGyyBENiNZf94wBBLL96HsL9hz2FWqW1cgZZ2
KmEWHoDSBQrJioULt51FCoyWF5yNaXzsjvZjOs0TeYo+sAWbI/7RnuxU0HlwMsMbEfoNqdQRisHr
jSUqpPKKBXh3/ILwZlwcNutyVAzDZp0FVo5pgymSb5xze7RCK2g0V+NNiWSs75KIHB1MoAdm66nq
oKj5MdJNLluUjD+Z9gE8uAj6lrXy72pun+kItjMgM2ZDnwL2fN1nbSpkXVPk2LaDA/ce8wqb2wNO
sO39Opr3pX9kzhRpi6rLC5/6mDk4D8KIZyR1HhQLMK+Y7k4+9rjLPP/0ua7xnslBOiRpptGhiDhP
AUTbnqh6polVVJOP1/RIhOKmDE8cOKDa49sGJezqzB6W14qzjXGxKguQZKIkNp+FvsSAHj2MlzPg
dI6Smhi0SKpJNQWTyHXjrwIuarCwxFqOWPaAChozFtE3oqc7YNCdEGxlO9+O0CNL+4Z6u5TY9oCY
VovjBQ77kajjGeCWnWUcscvPs+XLIPwGc+Vw4bS1coG5+ull0j46HaGExjF7d/Y44fe3prHBLQys
dpIVbepAcwKlyiNnJuifoiht+HXDL5eRSR73VrRmS/CRoptO6MKuAw/i4AQtf714vtIT/mQZuVjH
ffFv6OzbtGbIeGJaUdYXJ9p7cHFlKJEETTmAWTj2bTzvkIqTy3Zno53GYlVqBG+hhj8wal0Zy4Ub
KDbt9MCq1eMXYQtXqeg++m1lGZ96D8WY4OUtM2bZj4YHDS4ziP3N8SV4Bh+S49MH4KzPg9gAG2ui
VPgHPtjC1ljJ+CMUIhMlguQ5DZBqS7LAj/b5zm9uY6ov/G6Rswo1O+excWTrzQpKk1DK/eYuoAYf
9/uMuEFQTtI1m/l+/9oYisa03m7KMkFquAnLhS2gaxSfamBfNUX4Wa7SifFSi/nbI67r70k8N/iI
UerJSeoImF9HXjEf1qNyq9HCGWKsacBS53Cqs8Uql2vZjfDGFsNtuKBjdeTIG/ZBjf9nFYmK+6Cn
d3d7YSzsnJJODkKI3drgCj1EP1eSRIEz7bHDrz6FFyB8yHaj2cA7I9I08Za11plmm74YJ9GOpjGW
HFbjC9dFkYAfqvze333sv4kpdXctgz2m71hcKFTHB6VNhO+Y+HvpGonH2CCWhQz8/p7ivgEjLb78
wo0U1y221hMmsJoQGzgCoD7uf0aI74BEI8AqVPDWXzpG1SHjmi7dyMdo/nub92Wk4G3Jhhda+mn9
unk+oKtKbT7yLJMLWjzXRIF9pD6AmcLN3B6OCV0cLmil9+YCnIOdEY/xPBab7i9GT5JdOlCRlzQo
Ub5E1gekKcVfrmJO33OwiMroZBfqdEmOEiG1ui9nU2mKjU2wJjZXiJvtQLEi3zEa6jEnQTESGKHb
VXJGKexyVmcJ71NrFe4H0AbDZLHjYREcdekPpsWJhDt14RGmgIoA+gV4ZHEnGLOTymtN9tGd/Y2j
A+IfIv4U4J0USTRBNUZk+re0uA6dZrjrM8iFomh6wRhAMGRAswn6P7okRM2ZmYJSSgDHXsYZ5Jjz
Q//Tgl8oiKcAGUjhSBStYOIL/wyeIiqsMq9uZaUJT8AnQiDAWZlikB/UlKL6e0I75e2z1ze5sR49
71s4rkLx+zhwVelZoZ2+Zh0ZL4GJUUlv4GW/VD/wJBlTnU5k0Om9A0h6ol6FDTsIaYvpuxEQFb6o
32eiiwQU0fqYoo/IvgPhy6S6jkcjJ1bRb6GycPT67d8MUk0zCWYRX3tYc1oUgr2yPW9+NFJvnQbC
040a6XTujZPXgV98aw0FzCOVpAWOzN2hp+fo3nODjsT2AirYM9lTdYhWt9EGvPdJvHb5kNBCQseU
MqHC8/1sv+kvaddLJPF7Iwz1UHg89Xk2XhkeAC6GsiEKScg1JDoJd4jz6L/O+6x7cxZFVfBqdMBK
EbCCC79VocJAQ78R6Ee1fP/uRlFeewPMS6+qcXi2cemdWy7ChRTC/SMYaUfhbGq75M8HAhcDUQlZ
i5WbXxK7Xb+XRqw11bp/Nj78WwvsPFaAtGFUxhzIgofGpV3tOr9Kh5/tYBU+we8tX5rJzvxIXcKJ
3RLRHv6JQmJA8u6cBZx4ZSbZS18BxnA0S7SOzNfw1yyuxLN6zpQxEYgT462iOD81gdkMyatiJ5I1
NwOz0WenvfjZFtFkFKR6nyNqLCHZ5mTD1wlcUMD6BX88h/pBhN7vWifjluqkG2oXNbsqCM5KGDUR
AJvfLCzmaHQk/QYIQ4IrDBONVsM1Bgwi9ztfXcCDs5BffFiQpxTrd4qGKuQZTFEPmh+8WMR0Dn+O
Ld0OxJLpEvbsQHZRIE5hhzGz6dR8AyofGQp/l9KePkwXll7f2rpiDhFwRHvLv7VhJ2C70MfPeIYN
nnEg9RCF7WuvKooHgnRy6FHdjXd40rrftZ1daL2k+e6oV/a8EVQsQY2jmjD0SSaMubg6OfopfqPC
cv+rzVjgMiuhRyOdI0C+CZa75ARXzxKCbUesdXwjNoR/dDYYIxYBuijDmbFcb/8QXZm3VdQ1ouGP
0FX/b7Apxg5N6Qu8yNg1OUlIq4W6rSJQT4Apr4R0eQRUVEUer9Z1fTXYi12YS4lECbMegu3sRVoW
CmKrjPFIilzbjZj14B5rmuIogFLCmI2BQ+ZS0Fb7F7or+1Z3R7uwLNeMKol372Gfaz+i4jGu5C23
VbJzVGbE9T4beKzf2ooaKZdTegM2efGTh0EWgqiBfMv/MuItc9TQg3T2ZA264yvlbsIPWNkJbGV0
5eFnUOemB0bILX9UhdPbHVukObDLhI6vqMHpJuPGbgjCCq4XUaJqImOPFnwCKg1SiW/s0waJc+pp
QEpGgnnFQ8OiZzw5M0B1KqCGHUzXzaQKPhtxzXtRkky4TWv361Kela90IT1qN8DmeNg3RHli1IWR
jOhTZMLx+L1OZXdCbCPJf54oXD/23cEeMTntyOYaQIIj559ApgZ2ZVR1J55UL7YDDZMuuH6QZ1BS
J4MaxQz13ZHZ54Oo9rxxcOIsV7m7aEg1+rstBKZjXs2ZF9/UE0mWWIG6VndUfS2k0/TxQTFSG1L1
SYgV5CA7BrZxeSeYvRGWTUzx52NRjM3WG2N+58TL8Zh/0g8BFVVntKO3yTkOvkldVQaV3egJGz/O
l5FLQwa1+Ph5ErwdepPvHlAnCEZcutsYUOmbajRd/C/vB9lJjArCR4pGLbju3XPAL5xinSxqRSQe
H7VBdvzjNKeePkNk0qKskXzfIYhUd0VXKfaGk35n4Sf6vUmKONWQOAc9lbPPgVFmf9Y2kEMNvbth
v+qtfaJrb0ukpIVKIr0vvHUb9Vca8KHUNj7SjkAPhECWACUGAKySU7VCJP1pEtkP3vsqXOvfmzKI
jOR0tMlcta/jiydAf1CxPn241CBTAuALXto6yl1bix+G6lfYYt3hD8Ry8khg2IBUhsZ0RDjOVxMR
hJ14Ls2liCPhRT9Q729UgHm+aeTvbebscnl+mwjKz9xuWT3ZQpU2sMMGKjvIUvNKmHThfxCvyUA1
PxXOH7FwmU5+gDXu+dMrRBs2LcvClFMTzaMJRoOLSLqpSHROdWxnu1QGTIEg7tHOdbcnYrSJVAx/
BWL/SEjaDs/kZJQgEVE8YGG+c7mYA8vZO/HuoGR2bljSDy7V27+7uBuOJT1cOliNbPLcFC8lgQsM
Cl8a4P6CbXykPMc+Fxr1Upd7M/jW6LULY9LajkNL7VpZ2oZR8plQVAMcgJjQo/nWDuO667/HevnE
7ihJLgru885AmpYW7AJN16yPZC5+9+YSQBXiBYSbkZk+OdV4vHlQa5zqzNb6EaSJ7oG0zFifHRQE
QGLdzMiikO2BRDzW0fmDsuVyPhoO1O1s06ltzrflGnGnYjygq42RMMuCvUFlXYyO23xiSoMz+lR4
yRaxICQdX4TqLgcM4CLqrwPls4mHSiczkEiQew/ic5/h2wLuEAjE0dCkXnskHkA4RFYeahmhJGIT
XO1tTIAOam/Ep3O0g2wIM5BtZlniH9JXDuH2qBEmDInXRdJkK8knzObQHAo/IjwDBVqqrmcxHJi7
GXVuKa4yJMIGr3VtgEDswWB7N53j85ioa1oat9fT090dNJyoTBTsf1RsPK/+3b5/1g+jpwyH8Bee
0pshUE2HrhtyhnHpyC0e4UuCOWQ49qG3A6QMRdGgjtY0WaNhB9LrWcj0bt1x1BuaSCt1GoUnN2A3
TejnNbxLMhOMLGZuKwh0Hkj2jL1O1BrrC5ZtbdWNmAkOf8q219OeIwKsnDZL5027R2yzt/pXI08b
apFvHW4FqGE5blZtcK1IpWJ+UDVgNvzI19svqZz0ZWbx9I542oWEg4DVVfAb8NP6mR9DfnMLEDg7
r+ak7WjvRGK4WWRY8zo/eA+cIUy6ZywZ4wXcwduSnA4nEBgvDi71Rh++CAAtZMMvFkkHkI4BjovW
5b7wxhqk9kpj5z7h3g//cU7A21G/oLtVvceSJD2JgyIOmZ4xiafC+arTJN75IApGyC27/GEJgckJ
EB1VBwXLCfqX3afbFA0UR/L+34XVwe+QOZy9iTqwHJLXUd4ZdMgdc+L28nMRTdImQ/riQFTkftuX
m7OdmetMfhQyYjJ9shjPv+3q+r20FYQ7AG7Nj4U2/8G5lpEk+Hm/XmDKX73jUKBWwl9UuyERl6y2
eMnc3EkOCAELEXSOm43BPwtwjc8WqQf415v3M27xwLTJ1QQ1XkBBnSGwqHFXZbM4ZozNDWaQVmok
/HhoIzx5rC7Fz7zAYwq6GAPxv9wb38MTL0nUugxBuAB5CxswXvzsyLl6XiDlZWpyFNZ75QUDl1or
t30p7f6kJqH6S9SZm3KPtr4AmFq+gajXB9nXSc9xyrjw/a/265HI2M/xvR6Vo6jpNS3w33/WXS4/
a/YYxh/LfU59isaYkdImLDmYDkX05pj9ozdUAfLKMSIE1Y5eFKTs87C8iKqGlYrTRc5zLy4yDimc
3D2Wsl6OUY7iwgByX0KMTLXgCoPxcDk6rnrz1eVjw/xQvvlDDwfc4G7abfGQX19qMoPzSwsL4g6i
knuMqPMXL08o2VmqVgQMXLc/lPxAPAf9SkuV2qcnssbvjmsmpQ4hr5nRtgZPXIr9GDSOEdRrrAig
eljpFqQUYiqFuIo19xVwkYetOTag9IcU1cvwEeI889vFrRdHHZMV3mrENCshmEQB5Xa+I6zSPqvt
JYuWRcMK6jEg4Xl/ETI+udhiKqoqq9zZIqoSVdkiag84pIyLTw7Lzxi+O+Lf4v2dJVNB6xQjYm4r
OWvyZiCb3atbj1NOuPUcAUHi94EF8bSbdd6NkHGjwTF9b/hf0jZn0AqvKnzAqF+fz0PFiB1PxMB9
QYvS/DUtcWryrhb4qvfrWANp9ozfc+IK0uFl3MpXYcW9anA1f8J+JlQvtJEcLihhaw2JoVUH4NYm
1Dx1Zk53X5b0+RF5Bl46ZAbptefgPnef/YICN6BmXAeKPX7uqpXSp9pwtzGZDEnrukPYPY1gsLhH
E84wmGPdUfYSupWPh+n57HGDGjRA/ugX2FB7Zh4PPw1nzm3m+39lUNiZiSHWIkZJgUO4TCDmD5C2
dfAcBIp7CXTvP4I41kqwa/wZUIGp9Ik0zRF51f36GYZKVxaiKXKD9rp4dRFFoMRx3DjV0Anojzxd
0zFD2BfW9lg5wzT7PwPmgan8epeNFuWt5GKO1x2MVeuWYvm7161EYOqJi372j93AkaOOQIKq3zc6
csq0Hcly9Ce7ulxFSYau05W6ifnsW9SBo+3IzfiqLKjbe1Pa0Drt/wyeH+OGvyRD3BIEKvKVPoJR
8sTyw7gdC18WIPQ9b56OIzBa62us+hK/yqZjKpum1Du2wuomPwfzdsCe036wst5w+jOtvN/37eiR
U6fp5Zl9R8LJLsJEGMWzO+phRDPe1A53gbrS1IW8sBNqdcpkc6X5TzIv9dor3xMmJr4fmZb+CtDs
NGCfpgMMYzEdBqjP1UCf+qWoWMVadGQqDmVlr1VKjul9tILZEU63dC0SPtUhrLDCNw+r6fJhIdeO
HIkbknjuhOg135weA9WCYogNnYYpxLubuBRPIVRIT/rb6Px0zUHzhWgpkbS8cTWsus5kJueIuXAQ
jQ1FLq0S9FG9Z+79fcrTwJQ9k2bXAH7MxtdwEBkPlXsmsmFYMxtXqQTSboSCpeGS+8+xghE/AS8g
LgJWGvlSN90HKkBt32MPZY2OOJuk7SC4Dlftiuu2MAw/vd71KLMN9Y0Tn5ZxWSnGSrSNb4sKd6AN
ah0buDdknsg9kG9ecsNbW3EdY8pb67CgsQMWbxj8E8VHraSIaWfv/+ZyqcJpPul+svr1Be4cjMRg
b1FpfswQi/yDHZ59M/Zr9DLAdBbdMh/zevusipCJJMRsI7a1RpHg1HFVFWqzHu66I49bVvS46Sqa
OI5WZLt5io/69XfpqXB21A7PufKERwrvGOts7szq+AgdhK0SDvVeBgOQjWV+O5r+jIPE7pSTdgfl
TMfDA5k8KJUYF1RPAxaeX9jp97mtu3ucLlx1s+BAqV9EyRNErfv1ZNIyLS3JbWGRn640pQ8f1vBB
8JdDLJHjUwGusEpEmqc9BtTT1Lby/k+lxTbCqebSp2qRT5Oy4/hO25R//KGhp14n0KXhSS1QPmUU
gz11/4Neykucjd/kPBSEwRGH26jrTAmpKxfuI8TjgeaPsMvytfMT9yJVy0+eIYBEOnlaszSuPuZe
P2/Z+VRABe6lbPRCKEyvz3cd3eE6bpSUBM89xjtOCQ3VTYXwaNQ86/uaSkZO7eh978+Y9fO0w3Ev
WwQObN6YCbowhTvU39HAy8f+RwEMQQ3ghbCz6ST+eT7SOU0R9PiKCraTThGVFy0SqfmnTZxrmbxK
aS/j5k8ELs5NCvHWoPqA9IhihpqI4gpnkCplCgjQ2b0jHKr4f5zD+gkmJi5Qg5ZS3aM20Z6iVu3h
neo/5O71Fb4nZDmqjLLiC9T9SQsCNjIvLQwP67ptay5BOPpEZKQDP2MBsnRgAreI1CZc/Nm83+qO
9IbAVi05V0g89rbsZjXVThSzXwtu71HJk+15T579jX1a5uapfWku82QsyfKq7GQ7PmBeDg0xKcwN
mqBLMDm65Xg+2LoLUP/tDRTaybdr7dZJnU0LevSu3Emtny15oMcXFuUxYB81AbBmNza9kuLY6Vn4
j7J44Fjcaa7maphq6tz6l+VqFcPaorBMvrjU1AjpBnXtDeqq6MANrB9AYjm3QWyGTGfk3pw4qEMG
EPAes2h3MuPLKbD6IszNuqrxoBnYNpWOjOyO85zVj9qYXhK+pkNUjH/MOe4VGxD+MBPi4gTg8/32
JzdezVJ264El8fFVhiUPwYwApQ/Uw13HvSHN0VCFq6jCJCWWdFEWrLpV6xoX+5wIcZwMZGcIxCkT
jJpI3ZrVq3g/E1yRE0aCRGoIsMgWWWvjUkiJm/AWbJYC6TEOYtazqlaB7Ljzf/5/bJQ+zV7h8XBr
Dz24aK7k4ghGaipfA6J413rGu4PZ77PSSd33ZCFXZ8rAUJqGq9wOHGl4z88eUs1jfDNoqMbttXzN
DVghDCevo0Yma3u9P+vOEN53rrRBkTrLkCfeckqiB8HbDjcwqPgfCMSpVUGRpTXLTj0jlzTrQjGA
LAdbSY5iw7WmZB/qFL7L0w9jBtb2PVifYTXMUOr5HUHb0cNDckjT8uCprc+U4uw4KODFb7FLGr1W
JZk7cg5zcO/a408Ir7THaMYNAEgQmAjhy5B/Pda7QzkUEkZerAWOWdtq3qjI9jFWXqLq7I07twpG
OYpbPFqI+1Y+XYTP0AZ8o8e4F0qgg20/ZQ79Bmuq+QS8ERc0FpDqDCWNzQFAN9Nh8zrF0RYXkXun
hppL/Rk5HgGry8uzaKHyv6HcwN+PjCFTBEYxbmkqauQeVDPgkavl5mXY9Dgo3ClPZUHCi00n8WuV
39Lrlr4/Wf/biBxczm8R1cVrZwL45b1YpAoPr3RDu5EplfMezmhwewNcjTfWCMWZFDI0gGqT3op9
LwCqvUSfmUMgpmmCrBo+oNBzk3NyDBq9YiVYyh6s+aTl7Oyb/4bRnCEAecUpZHc0xA2pGZ0qfvr1
HvQwOkndYPgP1DjNa2S72JB3gBCgECnCKu45QhOnPLYqMAZnE2FXdwwKl0wI0a23gp6qCNNQiUnR
Ne33lh2LXsgl4oYuAcEIPfqd5GeS0c9dabI4hXjRVEJoSJvMu8/zdWQdTVyQfPHiLak6aSs3DP97
Ie1qhK609uT6n6a2fnOhWoV6LQdLw+1ZQDvutaAd2VZx+bKJ44MDdwqwPjIW4llBnV9kYhG0KbVs
DvG/7RlVSF+zHAcVVZuT3GJdDql9CU1lPhFZlborc0uapbF6OLZrzhvbMYZbRQmONElVwx+lKTdP
i1q6KahPem7pVrKawlZJUay/6zuTfrhbX7Ejr4vumGvbN14AHjHRq6GVrHvvQRJxIO4vIdhNFxeK
ox8tM48EmKneywKTq34wHzDpqMacPsdiju/nmqg7KtA+i5UCutOaGOZLJNOB730g8ioQbc4N44ar
sqFW3V1DakXGoqNtpqLbkslnswBMGHYmjq+wAiHqXFuMIlOFXnij78C2l7+RVRcgHjVAmD9D5X47
VcKwIkXxuRD9G9U7dr83XghuGdipliQ018H2jqpx287i9iJrAtmi03s4Hj6S0iL5M20dKjehCVw8
VW9/H3HhqvsOCdqNh4qNzu3ZwNP/B6od1ZxPOQI3lGhovaD8dLpkrmBxD6hp0E9+6bgZ+eLBOHIM
Kf0esYAyVBTZKKVw5MeCxNIt3NzLEEAf5hvQ14cptgjKjSUC4cw+FEiervMfkhLbRfHJaL0ksy3r
WYU084cu5aNppQ1uUAl2FacztEt/XTZuDx/t/hGkW/9CXngBBkGjPnug1cs1BCEZ1GaK9EjVOvuk
sTykBd/QTv70kafyjo8S31wIolar9HFa4gD0HyRN3t5h6XhweRRWQWhepq5ubTD3Jv3o0N9j6oOc
oVdbcxOUAn1v569wEtfL8Z6j8USs09r7AqcvlhUvb5PYudJJNdXtyB6d6UKgu2pchvhCFDdcEfqH
WXKIOhimR2NB3XHrtHN0TeQ6zTWASoz55WOCrZ9KKFciJQ6ZDh17tl5/YMLXtAcl23Km4Z02ATVl
8/Ot6fbwuze4zpcFjrlPxXfv1/5cy1ZA2HLZpXexnSwPFvpTz1l8xV8Nwqv/RKxWNUf1CrzTOY8C
9NJ13kmvZBl0kaOoj6+a5cHXqzw1A1rhH/AsOq+M7j+fS1QOnlZpX727sTAzy69lamVnohLyxZb2
s5rykR2US+rLoQZtswjMQl9xk6wTQ/XZ50g8Jvlq9g6krYpUexwHB1KRHM7p6DimkwXSL9zmJF+3
mIvO+gYxcWVIOdcMnPAu2imLbKWqf31p6BoaMVmiOgEFTHzGqM/lfCtgZLPmqvO5sFjQX7azR30Q
5f8AftxTSjkrwEL+V3XiSDLW3/KGCG4hkeTJMVR6g+YtDvEUYq6P3CQE74B06uzQkJmvp3xavcYh
wuEm0TqcVIOfsCB5xKaLFaLZErCHFJFwU0kFC5j4ejTUd2xyBA6hHZ9ep4YxsxuwifmUCmvy3iG7
R/PjCEaHGz2nUCPgx9VyGm5kqwnwFnJsN4DIFDiwpDVjROBylW41pH1o9ciEZCec1ryUKuujfgtz
S/A1U++kM0te099kDML4mfoliqb2IM9aNBI4qGPMApcdC84uHeJJdNndAW0ESAiUwJma5vtTuOLs
2Ov1YXuBQHmEaKOy+3CYsvfxVsvoovq4rHS5PtiIdWzu6SQN8MuhDFE/l/PZu8iA/w2leJKnA2ce
RFuYucJTeQ3EM+BUsMv8KwEEutxibRu3TOjO3t/o3wnqV3TNado9ukAzaQw38c+rUoQz6KPYGGIV
UHiTiN+9XXNK61/UPA3A0lnqi9B6rKU2QMJPLwL+K9dhFhYcdmzr/pQ16d0Hn8Gh3vgaP42e9Yrz
g91CzqyNskV/oQVbjl5mlyryPSoUVfrNUKyR/FPm5GVSM3nu+gkCxem19cbiuLv3o8tVC8KE6jQy
uK4aEevVfkP1A/CG8HJrN+omqCoFmnPqlhPoNd+31LDfkfGACbVCZJwRXuRBDqDukaVpzQ2l/fea
27uanH+cer/HjKlyLYHXiDCgOAYCG5mGycXrAjnuFIh7tGYNQksz6+fY/dDh8ihgcr3OP8l16bRp
5762bnACZ31jTh+xqhIRLosJL3P8lx/y4dUfZavoDxaM1bdVLf6p5IeSDJcZLrBIvuaexB/Bs+VB
C7IEO0//3OShxlCnqgaQomO6AMvpnbXEbFXLQEcaNQQ08BePAn+rjGeC7a1/L4DOnYpmslTUxZDH
WcW8x1MdWailVoGzbR5472F8+cPkNIX2TrQgV8lSGiMbFuH2+4zD4A7jv21/1KsaZnUmzaEe2vlA
wzjZ7IrNW7hNBNLPZQ0Qr1NHtufBYQ96zOjaEwvA+TJI7MOp8RzZAQRUj0Gym8tMn6/A+Tssy0mB
siBneYqqdYGIBBXj6/q26nFKPgNIswnfR4tT6s8RTRvQJ/i6K32ly0q3TqXeKlOTUcpSu9AO/WOH
bBUjBEuknM84ZVA3+9BIIOCqGN6aGbWlO1OrbYK3CJYhPL9Qr786IOsKwQlG4btpLRllvXPyxVnI
GHVItgMYyv4LGLCsFdvyRDZb+XeI57qcD8DxDlpA4tAvLiK5RGTB7Tzv9/LHiLmMLTaCELk1PtST
eWxczVCv863elORzoG4ayx7xsMZU8EKDRAFD1UkUJwHgDeCZAZ3vEN0p3y2vy1AeeTbdsVj5Uz53
Rb4WbF0MBClPFxuxqMPtfWoeyHyHVHX/zukKymQGkgnoSi7CjeIXgaYKGdNhf/ApUK736E5fOmiZ
35ux5p1rrjVf4dkJK3CdcZ9htEy7ZC8+fml7w+refR1sAiMrn4/jsmJ+RSc2QIMeaFlN5XEclR6y
NzGtg6SBThIQeHO41Dvrhhx01/R5we5hkmp+gGXh8a1klg521iTK2LyTMz3Cp77bM+hbLBIdUs1x
4hOQUT33D+wXk0YO6dnj0dcSNJ8o2fB6A1mvbDO7VdNrKBilVOInbg3U6aabcyK182/CiTpV6iY+
zJiEQ9vC2KXdZ4J8XmngdA3X311Rt6e4761MEktYQOZUGJ4JuFXwh7kV0/Rv8hipdM+1a0ERrHOi
g4xQUeD+iiXKW0JeefoNNc/2CmaolpvA/8e5HpKRaV9OEq9M5J+1evB+Tka2QdBLgNn55aANAM9a
mOMuUJnxBas2SzG0rUmedenFXXdYHzoiumrFT0W2/jblZT0j4lbNonK9ICa17eO3wk+7+cTVSk4P
mxVph9izhwCvrxXntQhd01VxKu8gqLuJUMzylojmVLif28usXN8RnhUOjUINJM8W7N8830kA9SZ3
hiivtVaDNnuiyBmyRgioqKm1vpWGTqlUriX4FLoEA2o3EkrTEarCwOGbZ2p7GgoQNHzsAZPVHIu8
spTbNdPjWIAUcKHTqdXMy409pAQn8NUFkNQ85WK+OCrNWe0/7eWkBqJaw0vPC70SRb5BRVvJqaX5
K3b1rXOtK9HZMQAeUvefMcEjEPERwTnSecQbLDg2VNmThR40fRUV9mABsZcCwY0m3LBJGMSyeUlV
JFnRMgTDGE+oa61/EJ4aBFlWl2ExTeLyEP56yr2pFBEV3H9zDL5sGaXUchrG7tR5MeqLYmL009fI
Ynlo6P/OmaKxgDSH+nnitv0OHddWtS3R95Sbw7eGDxb75OoDbARgx201tP4n1ngl09vZZtCtz29s
p4YKsi0fGOeS70EWubDg240earUp05gqAbjpVvMlBeJ5m6dCJjWzCxvjXI+VtcHgeyyYagHseEbX
ZfTlofqaL6VUlOY7EE9UK4O3xI0hmc7bF33c9jxz5DNBvk8JCfKHzsiDYea22AOYJ8hyTYrPudW4
JuhvJ2iB0AONNbo+rPwE6qCwgBijRQFjxrLQ/I1bn7YwajA+g4u2sfqFkpCpam5HLtHZFrD9vGc7
q2l5zfVIW0O0xB0zbwBxe3XI10wmpZkj64fkdJL0WKoGioyOlGQAI1H8OfLbp9swEr+1ExkU9J69
UgxIJAvdeaumLpwGJN4UThTrethEWFQbORehZWRQxYBvEefmkjEkbPxrCAL+D2qI3x7RoV4Pssjk
suBBaZ0w4yNhL01ih1zMyJ+/d8gPP1PnSG8+h2j588okdiOANNdPjVjsMXR/AW5Bpt8wsE21lRsj
VRuzMuWlimq00zPPqFbf7b9zAzrH3a9SSKIg2v6u1IvouAj0dYSZqZ10ldOxPUZI1FzM1b7IvKnq
0178vCraFMQO7uYUDD06vindyPquDgKQUvT7CsGmwuASni++9r+hW2Udgv5QkfKe9ZOz3W6SL1nI
LV9W1P2QbMWT7mCZPpYNrBC5g8GPwBfy+Fn0IXkr7wGW88Njpzbo9g+Ku+qTdeRkpDvFlisrbQSJ
+wuWTGTkb4dvwNqmh8/FT4uxeFuPd7pgmW4ldqTYJT9TICW8Qzes/Z5OVvex21rD3P1yaAEL1/Yx
/ulRCt7VUauEsrjRM5iPyViAQV+vJTMH3ht4rcd7xCUVTYv2twK0a4yPOYc0+E/d9LBPNs+NqjZZ
KxkfCl3IHeXSNVooM9IGMiywijF5PhjBCxL9qlUgN8zm0cNzH69/9g2OcMcvAcn63e26wApv1hNJ
tD/tAR8+nvqiccfo0sYRFYVv4CKJzTM9sbpCfJ1JFCQDIObCSkiQLlXAvK/SUjjfVfWKoei1/jrn
DfzuVFvt5i386RcjZZh07ZlUuom0GCtAK+5GHK9ZrxaJMlFQ03iZnB6bg8/OJ4gZSXsF2HW9m8fc
032rNcd3ekav0zXwCm6EWqQP8AIEXW2kOxEDbt62XYQpQpAJE/uZNNSwLneNJzudchJikI/IxFrY
mulWrsDSPnml5mBIzcW0APfk6DrGsUjED0GIa5DU3xK6CbCue/K66X5TmGa0bO29XJ63M9p2QBTb
LB4ruqXuH0TPub4ZsXGtxUNKFEY0WzsxzSFekLgtljRuZR9tr2pL1sSrO1RpyRyJWhFtvc9jfuTn
wvTt6EWaSJoqfEa9B2Sv44VAaTl+lYxc8ncJPbER+6GZv88mwI7gUNVGH+7Qfk9kgp0X3kk/Zbjj
90UeizDU/xg+FFov72GCmXuUwLyAeqA6cbqhKqsuCTxczHmy3mCsU8itm1ZxM908Q4nz98r9Xqcy
dmHRlFIv4FpwHc0D1U3DqZWCApsCd2chwgmXQKZjnoDQeskCl0DmSt+ikeAPHo+FXz9qodOD3U1E
Yxhnpv1cu+c1mGzIZ9JSFzfpKGoKlO08ZAH/P20j04MdYBdTyqDrpmHpNxp0kcgcepj39zsAbROn
W059zPWODpJqlzjpgOtOp/jELgNM25/Fon0SRyYMdaUY8asjwmotD9ZtnW0aM+yYfHdfF1nlDtH9
1mXuF9OA2iZYO0Or7qcaEK1ZaDYroBSIiH5z+vhGnrzUQ1IsvnqocR7j+Y9ufXT08deWpjl2djJv
68kCr81vNpAJ5gXTxEdfSVs0RZPkL7Pu+aeImEnMHqfhx+JVoNpohDVwsnEAFeAReDBTreVNMShf
lYauYWFj9ZPgX75LE5HJ6sJTsBa1l+J5UnbNBEJ5IN2SEFhGxARBVeqmfcSktSmI/n5h2hj91hxY
eNmHwvRbhyLIiOHs0K4lpasEKbSNJFXUmDEMgFKmZR4d7JLlYc0IHMZZ60ke5huN8zQZTRPYqbsr
Qj80xNIRkwxFo5Jp5fYM1wM3VA9di8edUB7AUa2CIM/wUYB7jH6ukTz1G2Dpu8dD+Wq9DTy/yVXV
TlA5Q7LP51AE++a6V/WAHsnZrj/50Q2va7jLvDvqZHrCw5HVHQ8y6JMsN2YUX/Rl0jDzmwx1nzNT
8bmutHkPgO0zMIz8c9pLAe1JUrkQ7+NeB8LJjcBXf7W3gFfyPYcyLzkeVST+eZMM2ZC2h24+/z4k
7w3/RYLwmYeG1c306NQESChabd7Tf/tjwy9Xrm1175h7ihyP3SPG2Y60bvJZI07E0X817C6MaiLD
wVUKTAix1XUfmTRjtIOIWWlCG3rC3pkmHFC4XjR6FPxTE51czxi7psReqKkZV0752+KMxtFgYU9M
M0Zvs4oWJTz6xOAeXHRbJRA777qmM87qfZAzO0/TAPiQBafPWuUntZiGQGV4Ts/CnRHFdRNbzXak
+VSGgTr9OHCLr6OMlI8HZTWrMR+VbS9pDTpAh/42JEhnj7Il8gAgMlnUIjhwVZFr0GGLmmIjMBgI
NapQHUid449NV5nqgWPoqEeboO1Gsz3fiKDshlucUa4fpkEeVyUqxPvnoM3m0utiQCKA6wyYaDli
yuZ1vFjagSb22ZRzFgo7+w0Vz5uJ7iq/luQx1DvvE+bjQcMw2tAD0bCIxnUk5A0nuVTSfpvf83Uc
r/4lvUzkGsOLHzrHqzNHcIiX0sopBAJEj1ZoDlzXLtcozogT2YTXthRcIeEzGqP6757M/dDSDvlX
FJIqmvCKgIp2yqSvnB5TuZjuf1oYQNwFtRW0axvFLKwZsI7kSKkCOj69NlRsNdpi4MhTeBDgPEFh
ZSrYgeKjSA3kBfhShAptXDtPdsOLfXfZh5S6Vq7L7qOoAv3DBeE9DXNdkaToLDzRFGxHBW5XGHUf
4cKk75dDrGCsdKBo2WA62ozFEcNDrEjLEK6/ka3TmGA+UIjjmlVPnl/AwgOAids15BVyrajUpJYR
iSI4SIuJJQv9JLGjtsIASrcPvgV96pl2uPhjsHRNpMl8EOMJn5cd9tHUgb7WKrHiuQkQq7e20t/A
rNhLvz28I0ivkSrYg+WywaJVvy6nJCJPNy2oyBkMWFnnG4i9PSa6Lbo5jEgskHdQMUmYxqUR/2Ni
4BIdlUSTNaRNhpMYzQZCBY/mc4ljCRFWcbgdvQ5Rv8GBP+wBJn9BE8CfoFJEC3BTNhthA/KA7CuJ
DudVhqwAAvGi5dut3PlpUNIrbSE73tItbsXyoJGp+JiZZ/BmW5FOWMZ7LWziA6W6uOhqMKalWWaq
9F8WbXXkpfKCHhT6Y+4tbwgnS0F4XKYJBH1tu7kf/vT/IULD8zD6gOTwYb8dBfzVt+Yp1SZQGdJ7
xqG3VulFCoApuyDXCWfadAK2lXXeGxiIUMvFzDxJkdoOWRXi1VdtaIak65rS9Zu8mhsv64wBBRcU
eMIg/9CghC1OT6FEYX88EOXi709Amr0rUh2hAKXPERiv1TuZbx436vql8kO52/Cur6ozc1eR3crp
b9eviWHARIvMTZMSAdAHJn47i5QSgavbLw6LJUvJb/eg4uUqyuaLNqoTGXjtEyIGvZtguFV1O2H6
IZ08wmwrqKkNXIU/4IeZN02EsyWk0u4ulP5rkkM7pFueUHVpxHngRgJftbFCJsa55ptnIlTxkY9d
kb1qtDvb4rsF5+BFWhJRQqqaaTqx5e4ErjcCyKCxLVg16GjLAmpXH60wUuA8tqwXwCEKXDD8ECvS
BC3vcrVBQgiHa3LIJYdxh2+r4wV90fB5Sb5v7zICzW0T/H7FfOJLy7hG/xtfDBcst0GMfijbwcgh
wCuif1tn5zXrpTi331n5oW+la0u0VfFfrMrYEEaVqKIRO/FGlhKTkweLZ5skNyKUddeiUdHQPmFD
eeHRxIqWXbMfJs6BSPoxjWHG0fE7orWu2U2v3N2aQF5ZHFpN61ylo9aHBCziMs5humKskuWXzvCo
UlfcUOqiH7U3oFPvyXxHsbBXk/n5VrflJYLBgutQ1VU51g1iFkbtlQABy9sA4WpRZ7YGvEG1zS6q
cUX8R7/yP6sXGbzp9PA5T3iD1BogxVLO2fiexbXtbuEUpBC7yttALDOdF/iIVXVZitdbSKyvT0wS
ly+YiqaI7W1BkiHaos7KhQL/ohmI5iZOfsq52DlmprqgymG+FuzWvDxESY29np8UpUIm05MIfXHk
+MLrJ6P5/pAJJKCtvU+fq1ixa74yZgsHThjImXj+x09KexjzKTFnNIy3gtIlwWyT4rjt8sO8WIFj
VHEavPigwbtP+ShYAAv3tIduP8tU58psS91xeSY7jBZWT3JxZMUkA16eUCC78upMYApxigQAXbve
2Awz1SqQsl9/ufob0dN6+TjymP8TOJsLQLTq3g3d/xxiFyTYMGEXymMVSOZqRhbS6JUgY3WgbP35
W/kjFND2QQ7cFk8ZrQ4eMM7PK4Hoy6fITDjQWTJRyWlsYES0BEWbVodt55YbiRfrYaVJ+yspLegs
qvN9utL57RgirtD2napOSLEjgRxsc/EuSmsvtsNsLklKDKitfdJxJ4gRVgRaRhN0/2HlW3YDIDh8
bI6wpyZp1K1WkNbBCvyokBgIhxbYccbT1pcQc+iY3FMvaUXQ9fID+P/9rCJ8AEjrq6dCkPUbeicK
1J9LpzxWv18qpAWjYN+HMMwn2AnPFk+Bp13hgfY5qJttPgo4OEqoUIM8fM3jyvbGpj40MxfzSIYQ
tWAcoz3KiN9GaNhxGk3s6hszG/uWOUrWSbkGD7aixze2vMBw2WeGtM+pcYKcLzc5ubHp99KKuDA/
In7tXogZopC1FJv6DJ28AMbTdxOG2c2TPLIQvFZde849goFMhjEAF5BImSJeix5f5eG/h6R+gjvc
PiiNo5rNyxrjGZce2WWhsH2ZvNIMeQWLqDniCUiQTiWY44dYum2UU0CK5J7Ib4BubIkdJ3d8xv3D
eKDQ3D4MfMbtZMvilDvkGEDo7+zGuGBTn3r8Ac4i/0aqauJZyIfJldeHNl0U4YIcaIO+FzPgkI2p
MAXuK16Sjj41e8T+eMEHtk3fTBBAoiUCiTM7NaN9kccGdCRxyuzQ2rXs3B7Pc7xqB1oj8OMgKYAn
IhNs+F48jRj9FJvUAv3CiqNsVrl7u3mjY6+xdZtCmn/mlmLT1fzj39Ww+/TK30e9bANj0YvOu8W3
59GWOmY8ke2crE4pUHgYMd+bVfR//pJDa/BCPyfZq5fVvzgpI53w5ZW/22TB/4J3zT2zpf9doAXF
RZOwjLIJx52k1sq3YDtDi2mfbYSoNjvA84Zk6NdzrkvjizWRuFtE+YrIpebxKuXOyvg9YQbKeB3I
D9iaZ1dP8QHdhlK7pT1s1VZWg5fO0aS+K22uMvq79aQANqLTNI3FohmYkrrb7YsGxE/X2JNnZhAd
UA935/LPKqhJ9CQ7IroE5UZE3223FuTXL5QsVEAc6iRTUKCGz2iZUc5wKJnpsnA/kjLdjbDgjOyj
gelhsOYqd8yLZID8KMXxfBT/vyOBYS02qfAK6LwfvPuiP7svji+ER4R/cw840m6RRuUN/1V06/dV
7n/tBn+DKynMmLKs6lvzjQUVcWVfMWoiID37I8t9SYB2+puvkI1mdrVlIH1outXCQYUbs2sBS+XX
Opl1UMpuHjwzvXtTh8uw62PabZhQOQDmLGFmLl3BBuIR4b4sny2j3/lj9VlITlY86M3ZnMK0awxF
SQhSMzpt0OxPvV1fsyHFa9IJ59fBDkRD6Ig6BMPCeaSdYiew4bh7pSX3m4v81Ra2F/55FubOJSI/
wR5teIbz/e5B5r3TDUerfDwNtfJnGwXI3F0AtScKErRvR6zEWPJlAYqmaVP022jlYoKHobJdDvN3
6yNcFgzDBMHsHO+Ir9C8nd0eqlRtS/JIDci3EIN/5eXAqhYvgLM0rOC1z0cRY5bAgRaaE2BTFeIK
RaFRE04TorNthmW6CMLp9voR7vK/MBt2PkAmlfdr/Wl0Nt4jZU7NYrTAnxhlL1x3Oaj5gVmi2S7G
p1nyodc5rOk7Ry1Jg4cKT9nTxSDmIG8tG5xo/z+e5wHK+qSESDO9Rx6EzP8khO+0tV8ZVa7chrp5
fwBOtcXrt9BmikF9Gh1I1YZ69a3Oa0Mmn1p+Win+rXeFmn3YyJHsmSvWAUqESfvsDpVBzCrH7SGQ
dtWPpsN9kFwK26n6MYRRzb/z+5Q2SjKpCVoHSbnE9GnsVTMPKbH5/hiJ9nBMq4h6GzVw0EJT63NQ
mZA3BMbMa9Wy58xRJnAp9G1bvgGUbEEIGJZU6IczKVVYj3cTxMI7Jf8V+EFHEqNFEzqXG+CLupb8
bR9hAmP4cM6wJpR0eiSXoGBsbxDiFoFo7CVkXLdNqPrQ0HRxeAwjnekzI/U9PABOSf3DPRfjmK8c
z3fB2CdWHCVXsJf9KAC1KI3IId/Y4uSUlI1Y/j/GE/4I5iqhMp2WVsOmYVDsjyYXpmLTiG4T8gaa
CLUU0YYaMgFGtH/LYKelvTSQTn9r2UaXNwBaxP3Q6Qpd+DdKh/tayvjqGE6AEWMjz2uioRgE1ZwP
gasKwUJhaANXoOEnJdoLYgF7tkN5q1435kP+Dsy6USYS8EdlE8wV6zbyeV8rlHy8Xjl7+yXzXdpv
HfUDo+wRiXbkVUw9ioOkCbrQlyopUoewcM+SNtdplkFTwxGK/aTViz6vI9+L68EbSOZFhujVTGTj
3OVkEmxEHcdRy6xxIq+sUhhtTZ8P8AhS8EbJdlt9zmGYWHJLL9UkI/w+LhUdHe4b4e+Tm2wQRn/9
mNLAik/IA1RkfQNjufyRV8pccdHA3JbIazbagUxdix8NY/EujbS+9xow/B4hlU+bNqSq8JTeWRw0
wVWSaWBV0LfSakOlFG+1bv9GdzD8o+l5pmtwWZtb9dcLfiL5llyA+IGXoFIEi7OAFbTIuti5DdXA
GIAeWwBRR2eW+VJTOojJt1blKIPcubMY0bqc6p8/TxpyyhGwukJJCeSvVjauJR4cg3gMx2f41fXI
A8GP1Xw0nSBWw7PHoKvEAmqZjo0LZFw4vc80c9IzehBEFBVH8UiwshqI+1ZhyRgejKVilWSs9GUN
uldP8zP0o7VY7FtScrJWQl1128K7BqLpueJsnVnuwP13qW62SN+cZTTj1Z+Glq8zjMATHzuCVMlj
U67iWadUMW2HRolRmBI6ubiIED+osk0hNybT1RB7zKDPG1deI4LTZr3VJ4SqrDHTO0LJ6rKUgCgi
8ioHt7BNJkbZtjDqOjplT9nWs5YsW+Tdsrnnw1rKn7PZs6ULYt6b4+RGHf+uvbRIpbX9FbTwdWcD
RBb8Ko+wGdjDM4feMeac1U5O68/UYsI1vsJoIo8K1sE1WqCpAaLAU5KYn/E3wUWcs8VFd5QKijG6
o0pYVR8FJGbSeW2Y5GTLdbl9nSKWruKx3nYwOAb0NPFsfdAmGko8mVtRMHMSp71wrdvt84eh643B
eMB5Wn1B/pCEU51hPb5ZOjHk9B9FMfRJmEaMbY40ivHTqX0UoSG9r5boBrM16ngxOLbTgOeXfAJ/
ywunjH8Y395uaW/VchVmn0eQYCmHjiSICwzBPK5SOIPI92zorhjhOO+krm2RdbnqupbTSqEvdzH/
x8iwaq1q6eR/e7/DTwzIM+UsIdua0ogmpWQkq+JwH4NOyxP8V2rxGwm31xC6nRzVZgsHwAY32vO0
rX0VQKl+XjVeca22VzDFxYwL3U5nGRI6u1y4g5YigmClNaaD8h9gL4hwp6AcA3iHQkGgMSjTJkJT
q8yEsNI4JcSkYD7M8uuCFfQEjWFqt+Q/smRN0SwoK7sDuqTioEUr6iLrbPcZMrB3+NHFUAaLBMwn
wA1POkOd8ujHBTLqnkCzb8eYstu2QHAuK1ZWP0p7ISZgUjzLbK9M3TMjUZ+rLgBp8EWxr73WLN27
ln+rSlbBXRdm+bMaHBzywOjg8A7ZUXRSfrqGo7nrQcXxTOEBqT1Wn0ut67hMi1kEd/ANU81gnwB0
vh4cdXUxOgCUWGCbywVVCJh1vOm3ua2de8qfEU9cLqcyEY97G5iy1kxeuNKVFbtJ77Lz+ux8sCpJ
BRb+8YmfRljaJFXIATwNM477UskkfBeZLIb2+egWqPabB/v5ZFyb0ye5Cb+kaC3LHxfOYS+7PcuR
3IBJBVxuH5gb1g+eZq/3Q5M4XQ8f+ti9c5a5OOW8uNeGIvBECN+BP1BG1R52l+NNMwC7TBLRZhej
orfsUZcoea8nI2yDYoB6e8LVfbcFl7mbo9Zq9LmacTwyOgIhSqe8EDhyqrI6l3MpgP8DJx3PFWgh
u4tORz8J5p4EktbYad5FunQjN2bBaR4Dl4M0i8Dbrbmu2I3lpggd4rLg9/H2A3HkIp5HJx+38pTX
1q6w9S72xQm4IeFU196zu0u+JyBLtYbuZpvptv1XFFyYobVVlaQ5YXauHKmBlfX5oyHAjoAR0Ouu
nUUIUws2KlavZ93ihuCXF/6PUHI5WNf4K7HlM3t2aT7Dknmar81GP+FecSlPsF8UbI92FhgyHdDl
3WoFkf/viEm11trwBfMwXpmKps9KTWvQKniWiqPdJ843RYzBq0/UJ/LClQZgU/AASaaHylbf48ta
23iuSh2PKIC+YTldePoFwgcUNFuWNp/uisCghGvBXdnv+F4j/pM1tJjhZ+1bYOnANZsG45N+NQdf
Aiod5wNbpwNxrgkzS/CT0jQ/QN/J7ZC8tNJR0Bf5/WwLg8l8j0iE8E1kNd5yJouyrAaGIXEAmUXn
KTeBY8VUk2jbY1Qm/U8VFOKhj6LE+Adkx/gF0QTwN0sB2TkEgp9ZEiNq4JpHiWYOBgXjb2KUElwk
7xKggpcKd4YdIHDy5n0mOvnRT6DaAJoZCLnV0l9i2Td0oyI2NjPTVATuChigLTjrS1KhsG5xCf8x
qZTHDgXWF7qzu14L5YnVVzJ01AUhga0bfFIjZ3Tq8l1Y12pw3bL7bCi2ZU8XGhJZazldYrLYd8qI
8Y/BFFOZ1gm1k4y9m3ssfbd3vRreZpEQD0gGKfxBVjGeGtq4FudGF01TO99p/2qYvkx4465iC1s4
4xMAui2Mf/gCIFmpBLTF8NgCxMN3abIVQp82Y9Wsdgt7EjX1VUN+M7YkuqS9FOP6aiy4ZwcJNP0k
Z0HgTwlFa/QF6m/teA9So7gX0iQ6QyU/wmBco61F7ohufIVXObKF1k/1b3Y7Noz0SitZ578hQ4fy
gfBtp67ah0Msxwe76uGEsV1HlmWweN2mgcG19A/sj2HF5zzQ0SRkaoUtRTJ/fM9a3/D8l4d8Qe5K
aVXQS3VmSb0shzL8+B16+6kXhwLX0m6anygpcYl0Ud4tR0AmP+g4ORPQNGdXAGiRM6VcHZ3PoHWt
2FGTWo4vssbVBkSAj3gb+E60MqHdC6nl9Bw3DcLFzRHCTPQviZ+H1eQpKvbLNui7uPRJvoQH29fM
/07C1/P2d7jlqi4wB/UBGoEGiA5P41RlYYqqEAB7C7gLzAAK3inpg+UPxWJk6vrwyBXojUitqXwU
KhE+rPD5tZ755swI2510XT1CEMerhwuWhtv+jDEUgzFfCFzaE37EgFahZc14JUZP8/PE/v+vWqUE
Rrcn6ZbJZp8Cmz0ZNFal2B7yDGpH85VBFp9MylYlOwQMPpuih9/EcCz30vV4MXRRAaKl+AQzkytl
txs6i3TA52eetqdoM1bXgAMjxoP1XghkGagNunPZ+BmSETY9/dFanqQ6tZlrM7Cfqy69SwA3c1jg
hJxvRXx5a9JXVXmJyUhUk3WA8UKTXfwPDLg4UJ9B1LhDWhJFJWaYiiUWiqpkoZ415bU7PZvCF3nB
IsC7x3FnwHJep0iBO+p1AbhRA9+8neUNpsTeThp5ptKO42/ewXMmTaB7Sx8A4vE4nd+JEZjQaO60
ADogHWColBlGudMV8PV5omRQho/zVo+1zFkR0twcyU4vWSUZvVfly8InvuBGzIoaGtlMNkZcUG/t
wWD1kicrRJq7YXVDWorTmECaCvH8W3Xb33UaLeD3c0qt9UFGcYpL2RA2d2874InQwZq9kkswj14E
ql0HjW1ikxoOFyJ22RNOOeUgKqoMsKzOrDReOWeCa53FWju9haCPQASWV3EqIKcu838/lmJl3LHt
No2f14P88CAymGSekISZroZnf7N7amGBQCec8xw9IA3HzeHeCNDOjrn+w0k7fn/XGLHf/hhjMsfF
bFFzFsITY+/7tPgHdx6CTCyjt7ku5BfaFv3EFetuoHGRbQb90ijG2inW3sNJsMum0i+H4PRUvuns
+F5D7w6OBaP80XAQVheXm6GHWY+l2YXy/Zr6wtRG9NXwhk3UzV3LDJxHSawz6QylYTQBG41lMrXL
5E1UW3VQst0Hf8os0fAaEOaG8S2VQs+r3JzoWcPzP6YPTMZ/VFjUftZyJwEzD8bMHNscmdmCWqxk
e6zLnWgkfhACH6RF2pZxz9rQAA3bIYgHwvipufEhYPAxHFXZcTElIuhj/Sb4/bscglbLRxC4ZLxm
/Zx575hyxCKFZK/LR/AzGD2AaGqfVIOAAP8AaMjUfYB6ZHGjcdxKyDTaZYFkZDTfDWPp4WZsuGFK
6BasYSwFzh+GgD3VnY0lPnqFibeQZmYPGoMY3z8Q1QCk8erqbug1aYqcZFkd+ty+1HDWCp4bdTwG
ntSYEmdBoPamEyWWUXDuZ9s3nwnj6PajvtCljz1Q+eFq4f01AOODPWi6qboIia4cZGxyptAI09xi
usKokAM8esI0dOQdJI3aN5lEVXSaXqkRZ7gwak5YcGsHyuQ+tnP4qgmS6uw4eEgkdhLiggvmI7Lk
PoSI+PN3eYwUDwLq9JRtWunpECRrbecYokg+69wNxRJ4SlHZc6o0sTPxNDtjYE8SiedEThAkJYbE
1eXSHQxUsru8omrTgyaysNNjlz1VjJNfqmZSsv0DiaYE5Jd1o7T7H8iJ/UnyHEeCGWxkgESmLmni
QoUMIYsC9HJ1xUM7rC/Eo+ykRuzYbquba5aFxBZlg+s9zm1hcV2rlIovlRRurYGGNqjPzrXBu2Zs
dP7IYPo/7CcXgEhPvubSiLYnYDdkC4ezTCCrk45PEhLU8fww4Xtw3krtROuH8AmPcWn4J+9SJGmm
lSJwKCp8jLxLtmp92YnJPqIX5vSAd3DbkwQVsdNvLcMSujbZ3UJF1Q6iqluLVRB1x6nvsHwW99pB
dI/Y6/wTgo8ZoRns6E0uaBBR3WTz90ehnaN+C5WAdqQhgf9DQuq9FtUcrGo5U0iKO/E5qJ62VmG8
9GegpMTA4ndDejL0bmzGJMO+rR11rgLujL7Y5Csgbzz0gIsfyaFM0vX/kZWDjF1unFOFEPrG/CUx
32MnU/wSR2bVCDxqoP3MATXqvO/22pxYb5ExbyyPSysQgLhqs+CHGrJyYTggNaHplgzkUJKDBSXV
tDtbVuBA5Q7A5qfGOW5x8INFf6GbzwIoZh2w99zTAHEEeGeBpQ0vMMUNS+Od7onncc82rqxIcLnt
cb0JTEMEde5hW0ZnWV0hE+XxnT4vIzQvrBrwWn5MWv9GO04QM1M79VO3vNJqo6dIdZgx0oNxZ4Oj
9TA7L2Rq4AK5nUjcoI7rHrAVkRk12Nl+EMdZAhTYRQFrN2nD4p5HYlCh/cdhB7DnDa6VXTrm+Isu
LKc0Lv9GSneTrIvQcgKRjSSjWwZd8WC1IJH9tam+ojrF78JvQjPzEwFN7MvYtES162TuLQwkjW1w
0zlcOlmDJ0SPdrXcvqx9sRvy/G36RlKIhzFu6z6sCK3lVmsEPOXLsrmXMYpIyrUMd+vdaPzsupVC
BvvEGODT4fBQ/sYPLsFZKSO9ryYyqlnqeQkhsdw0XGZvlwJCc9YhGUoAuZBheRYFlNgQtFXGwWkf
uBTNMG6EmlAoqS0WlghKQ15FNmI7XUOvBhLALgJXx8mX4ERUGU0vMgGAsOJP7FfMl4oVCLIPVtnz
HhnDBFKYPxPqkf0N5QPWL/ymRTSsZZHiE0ph1sp3hi7X0AWKrNOYPOwVTaONNoHVNcFm/VnJLZ6P
bXOVrFctqgPNU6FlVPfiJrVqpytpngIi2zbuDAeuMnThcko7y1cY17+1kl2JwF1R37dDQLPq3Aeb
7/4vHcRytvOiE2sV5fH3OnoiNUkK5uDJhNamW01rHo3zLl72BGjBVmQg1IH0RpvrRPhzHjfIVcHB
T5jbxOOVfxKxxOX0aHeY1dHFDEvTDFkh6pRGX49Ad3wlO9GJM3hCQURWId+PBgKuE9nHrDO8tSZq
Eap1bBI09uDAzzrPYLeHaveo7PkEQOAOqEDODXvZVYjpGcU77XaYZ7zP0GEYvdajGbelFc+2pnD2
jg2QTa3fi/25GX9fHhme2k8zw23UTnK/wMPgSINxlF3uJCvUic3Q2jNj2DZ+Flq9hCX+DupLhRQ/
tG7327vg7hFJ9MdzmAKWMIuKorg3CbAw2FCA28+3ATVbphbOByEnB6yfI61ocfU/ppmxPFm852o/
Q71lXHSySJ1q8nzuXlu0WzGsCNVR93ywGlTmwFYfh4vrPUlo+EYUHehqdOt9UFhxp9FyfpwFEtPN
K/qyjCWwESP1JSrA2dC+Yvk2X1eiPkTRCGcY2JHlQdlbmEj9PQ/gtZMarHSTeQClzXtcAukBTrua
LJf4bvZ9PJg0TrjnhbGXLWB6rn/RDA06c9yBXbNw2dbzRU3cQUT1Nvrlvlj1v+PnJD+HQX8dz8SI
IaEOSUSkm9utpTQ3oMBhLR94JhDxQrOeVt/AZnd1UumAkhWq0laDrrCsOo7CEOEpv0UYWpHJaTIM
37rSignzgIMih/IE84OtGfr42VlPRLjXIEMK9qwFZk76wSyQVz3ulafNEVbfo7OSgzheLJDMM4XP
a9PO0s9DM21XlEWpAWTNiFrLMNYONE6IuA4+7+mR5Tuwog81XlkMAwWd8GiKv/x5N+FBb/owyXEy
c0o9aPZVU4s9xHzWTZBu/KB62CWuJ8EXCv4kb4y35yf4MwXQFfFm8m510izTFQxrX3TuKDd6JMIw
KeC5/ofPXkFiKnipxAISXXBwJxoI89FJnSWx29c0S8M3aJaMqSHRvqmkIUAOd07v1OwJ57YeSSej
mDBJ6g4lq75NdOYgPEfqriTFw8Z1xmCeuC4R/8OnN1MQz5j1Yi4wkyxqZTIzeZg+bh7fCaNcBxgY
MVuoRx9yKMKwZYCdcfx5dHMOO1xbQ5mInkZFRHvQyBcIZYGzauvVklSCeP1yGmfbHrnGozfuXDV4
7lguovG4afae7TCwLVThfrkfz6cd1WbNDcloKKIbM7ee6/CPVIbIAWHTovvZHMgM2NmGqpA/n3Mg
6dyDEjQfktrS0JJ3FPFM8u0DAXPGCXjLh1u5zRW8DUyPA/HEMq7XY4AiTiGcz90dVN1EC696L/17
DzsKqus1YtYrDBraS9vUqHC65e4V0DIl500O4dFF8TRVYfyMug4181o4WQDQuDDl+Kcj6/A4jbqB
tB2VBnP4Ftu6i8sMlVrvyTdCmgRpuEvTdTgmfPG7bUR4y5e++UwGuSZRQ49VKBxN3E8TwSscZCD6
jNo9kCzioEoikzd0od9dQA0Q47qtCpQi/SZuthbVTCK7s1Pm4GvgeZIfPnbHuzyng2xF1Xfn4YUC
Y5MAUJFCP//WyRwGSh/0WAG6rUZeLOYXtPlaIGpOc07uMy+Xea5fqFDk2/6+Ry4MUNefm7RTu+rt
9CRgcBrXSv4DoRxqISr3qHC5qRuGUm1VqZTTia2CvmU5f9LB9aZwtARhel35jM9C6pvx/mmE02xk
liD7Zu6keydi+R1AXvFQEIrtxlXyC7Zm6vBxzn8TAfyOUsodoHZdHSVbKAdWQTNC8kT3k2dUBe14
5wCf+vHNn212coUM+KwBBEmSb4v6isFXB6wYzfrAxmiGZ9TNESKRYqSqY/7QQF4Nf1TUjbaLLzsr
XZR48TG9GfFoTKdu0Ri41M1LR9OE74gVPxAhLtb0cwow++2vr1sartL189XqhWD/Gi6i6EryTT4x
1S+oNpbp0DocXVIsMS2kaMYfbsmOyfLI7zqSVHWcvnjiEpRpKXMMuz9heXK73omgveZJ5v5vvzY0
WmA266CSfzSxO4IuO4sVTu34HLvYhaN+gm8NuMMueYeg6H4z0JTgEFI9t8eAnTE9TDJnU5gAvpWv
Xper+LFqVAHSvcXLbfr24LLzOngGVXJDQNJTI8UoVH4DMC22NcoJMynIICto438h2zRcdbNt8+y1
kEFuM9aQMbFWRLGcxcDyk9CU77tIlBkZb4gJ7ObfbC+R6BB5sIMjFyBYDU9rvEc5+zghkPTGgFuL
zx8I/AOX+0cuXiHjPU2lRI4BeXvjSXYAxWq5z5eKXfL/zVvoWpsyjAy+e4owga70wvud7FTidE5M
RbPWGGIh/XcP/RrPxOdSovOCES6b0a77LJjfGG1HlyHrn61AhqM0ukLuqhtwu7yXWUnBycir6ilQ
AvA7sZ2A70bIRDvmKVcrEclaQ5WXvByy+qGjrstTVbMtAn7oTj31LvsvfmvwvoLKgeSKDLXvJnPk
dZR8tknH7+QqqOqe3dyfR5fvOMAdPhoSVCX48jj+QZ38YTbfhl+mISdbVcw9OC/VWuRwxyBIbBM2
sRPBwu9ATSrjY17aHatxoDk04nes4lSqRN1DQ2Qq9UhQnJELCuMX3NUwC+wLLarMiLSeQSbCAIIm
BrlqzC7MrbpyzfAUYgTGWJje+WUY/M9fYSZz1usrfaTFjqJ8Ecuq4tXTvSOMzy58KlajmVM4qyEL
WHw9suunUUKgCfsyuEPkqC0UVH9P47y3jWYaEOv0FyAyXIpxtmm6NsnXwzCKywNcRI1vpGWosiEk
S5C6bGibkq56dC1haGne8RokKQfe8eAvB94D8gbqWmdMB0+dP5/jktY68tLly4In0Tj+Et7m/Tt9
SCSbm9gk/OXWZWr9LJW8zawgiPq2eb3YfDnQphTmxAd2eadrbijdRQ7pFdhkr2FZsuWQ1VeIgoFl
jn+RsYK+VFpAtV4PuTtVKisy5Y18Hwdn7IiT05CJCy/fvnlBR9rq7iBAQZvKg7zJH7h2RrNj0yrD
aYMm7GbCflJ0LTY7SbFmOQFiBcLjZVbVya3EUoDQOLZWIU/wM6LKLb6Dzo5hbdKyhKkan+cM0prZ
rXS2Z5Atu2SlCTJMJ/D3mu13948WpNiKRi1q+1tj3bf9MOOJBBsa9TNCiRydt1FnUTGFuOsbPy05
AK7m6+twdBCTYHO/UalyX9A1jRRZ4wudWkqOTrSvURFBX5Q48+YvzRG2KhdmJ5iJLTclo+I29NS/
BQGK5Ha29GKeYanhqfmDdXtAc7JOqhGPb1ZCtM8gXk7iY3qbYw0LDUKp7v7pK49CRXA52aFr/fiU
2++nHuiFywdsdImA3Qoc3yy2sWGw+xaS5lQZ5sd2+luPOfiYmiBU3JLLQDUkGhp7jyW1omL3llYd
IgMQX62fDWdeNJpbifMXhodcLcLO4hTMV95KddMzwmoKS8iv1JJlVYkiFQi1ZzuQ9ArtMYEBP/8u
w9s309uYlw/0BPUAaEe1mD2sCTtX+sgnrAGGup5zRSH81z1wLoQj8NSPmaZdAJR+fb/1519U47mR
bXolgca4Ti/mG45pXeqH3BY2CVBTjtKlWekVq6fm64cfAMmGl5R3lg9Vu27UOb89AA73517m3d4e
tcu72d5YXQrdsZn+vPSGc/DwDZfm6ZrVRK5crc7dzNn5jLIYwL/ImZKx5MAc+gieWvnLypumMi3E
nspvck+A8p3Pl3VNU2WHJz6v2xwdGTiFrpYdqTBJlmHyPlh3ouOgaHEmImdOqsPDFOyrrJj1xEMB
qhHuHtUkuB5e3k4BgrJwvO8zWTrMlGFpgqW+C/m5KXQd/Mrmgr/XBVTe8ESNH7QPiZIZAQk2QAjo
Ve05u3faYPK96G4LUR1Y523WqWMnClXjZ64lJ0CKkyakjh1uQfNqlBqj+EFypNsYu/Ciz3jh8E7W
iy1T802c9CPQRHMJ95yhqv5rxaKISTbCdHgjX6cw17CxrMrKwnp0NsdNhG8zs3pYij9Let1CyLCI
T0rRE3dz0/PFQiztgovVEXOSmZfq5tkfQ69tZvguEKTyG3J1R6PnnCQ26tO0branzQ8YumbridaO
k1eI19SdpudZkAb8lKBAUmXmxgvtljkMHIR5hJ0lL1ED3QaxgddPI9s0wTMXEFOk0Dn+EZ5uIx5N
+Yjd2cEtgTTUagQGL9ciGc6d2DR2Ajk8kLgJZAr73bVScjOui+uQIxzQ9+EicMsUnkvX0xxI9MwG
O2ftJXBuCoH0yrKVcig0XXbnExYGhKZtugGw7jxBwbn6HrS15fceRFNHm32zlVUnMIws6JaOOSGE
rddmZ5u3G4FbWCveqkR1Ga8IEam2GOfRio6LqDSnEos7AOIuzpZvrPONILbjUnEqChR5PsJGJk/K
nwulinVuheIuLOU3MZxX+XGnmcs9Q4Fho7hdANK7LjwgdxbadXI1bVC/Oc3GNsDHXWtp+ILOdbei
tPL9ymCu43ALqzYyxNaRSqlLyR9g089LJus99FLbMcgmcXdW1TEVSpT6dCbpmB6LnY98HWYNJ9Ap
dl5reaf419dnfP7wwYw4X5uTUKzawcZVbSUOxgeaJxiGC1/1mLviAysvrc0RU1P8ttrZHvneSPyU
Tl5SbAMx/ps22MwpiHHFQOgexwQ90yP56m7flprga7++yz3h660EJLc+ANHtYEMPz7ufcOmOmo6E
+FPamoksQNmNFNBG2nNEQZEYLyzT7897X0ot7hWi6gyDMBarZYYnxP4XtqpbbLQJEAPNt7oGWsgd
1GGR5M9bb4HHjK+9QlZ2eD/T6x0N0WHAbaxwuVQbI0HHvjL7fUrjxTOBjmZod3hgim/w3O0SJOur
ieH08CHh5Fvq8aAFPKrktAS5A7yt2QFkRvI94vfOpmM87uwD8iLS7VO1Af5N31kwE2o7WHuwj4Ck
wXcrHaWJYhO8qN0C7+Omoi1Jiq9EmDJaPTNS4FmbODC5Uy3GkXPBS0md3KBYZXTaW2Yi5VAOxDm3
OmOzD/CC7sDYlY24hw9pBz1AamG4ucdCge28VBoYr08nbwEHL+rKb1nN2q/eJi3PcvE5jjNDaxAi
rVwRX/+T6QtLG2RZ36uJqmYGdNlTScHTwMqsG0HcJlooD2GcPrz6LYqoJKmMc9fbCAYPkhqXVamz
LkfkvzSJDOZtRnX23dl2c+iuS/9aFbh1j9Vno8gTn4Vsb9GJnYIkCIsIbnTrJ46pY2ECBMu6HecU
7mtErdGXdUrd3PCx931jqBM6EnOvJvuSfn61raLel2Xfc9XeOAvrypgwBHp4IKiKMP+ARCKUn0WC
zr0MpQFCRUmDrTrllEEzMRffLGey/uaP8CuvzartumDReYduYS+mdD6WWn1neLCXh4M4HuCfgLWx
KNRecq0wver5SqMx1IRHqzU84FihsWhEn4SGpHtPjaX85fwpbb0u1BRS9DIIVqCrmpfaZZixEjVd
KqjZ+Gwjel/4yvZKkZkahVu4uVVRnWOZwPQG2erfsEFyRhUA9rl058d+2c8pTYFstkvtEF59Z9gb
jUU1th+QGX44kFx0PnIiecNQYiadk9LzC6KVLoCqubk1K4XHQ4GJg1S0KF2Vh149FaCysosdZNbg
hDJ6vqFbE2JtUl3vlTBe4fPpBBoYAHyFbd6aZrhJ8iTrkR+lYwbCswWa5kH27ztsefV2Hi5uoyIX
vjD0njfdcEKPvK0aA9JUOA83trShRUhAX2R4fAYRPEsylR6ene/0ECtic0N2apwGsqtkwrDSEeSM
pGL3oMfblrE4jS6kIpgypjfX/NJWD5PMJXhNXWmCCkNutwNQ+Ok8gIeFOFZgSbnJUhEGRlcpxurg
6k6Kcw/FoswvkpzTV/OU/0ylvi8/IjCNEziOd5NZ+NLsUt919YsrZE7xmsyqExKxaDK4iAcUv9HF
2k6O15svk6kNuti5MhYOnyNOIId4tCusHkz8BgliifwewuXSjdM+0c9slgUUTEXTbVHq5Ve6iWKt
eRO9IYJTLXoavWxLIuPuZ8S3w/+NCw/VBZ92MUwmYG8f1wNznOK3mMS7EIZfEjHA1P+SfAgf90ns
6XtGV4gWUqMlERrYG2ePzLBKPAHhvJAhjcTYkVyr7nL9V61kRMsP7PcIxQlKrc/oFMfHFBx/pJtR
jfAjghnXR4V6EkK/amRed+0e+kOcF5k+NQg7UKRr7wskEBCPB9+UTVk8YQa6k1ZLcOSVo88NWMgX
jNAfB+Ljll6njB3w6jWprAbQb7GmaXQCYTlBJ28vbQM23y6U3zZM/+Skcvod4gMM/pd12jdaQW5a
Lmi2/JVMYOj9N+8lcABdDhcQD6g+OldxcvweSrFOKg4QjXaFNmMkqL1jryikrwwys6I58PKpHr1z
lcqo/0hCf2bzZJWFBS0w4kmubW11v7ClXLM2TGsQimoCsLzLApp8RVtwuMaiQ4eP2BdXqlRyOZBw
eMNZhczrEFkHyEFU4NEjJQqbQfGzkbf+QvR+RF+4cL3No0P3cIUcPQnSxBPASpBFaAEt5cfHdi5t
L8MbPTqECW2rII+ibBXK+Xi5Cg4JrRu9i/mYTjX5Sdi6TYLjlS7Bxc0OSWvI3CV8g+8m9THQ8MNs
vLJujDhI4+oAtpwORLFWM3yxUAAgjMXVCEnXQjoqn1dywN1Ef//8dXflu3b5b2n0GJbz+Ekat++h
ARKqJVbmeB3SALjB7JHX4HI6/SRHjRjp8OuYYrIdiaAjqEYWBK+T10js48yAaq86cm4OjJsKTL4n
71pJ2t36veVUKo6vSzCfyqy26mcoOszz13sWHB+3y8lhwrkuApdSKeCWvm3uheLDXbzjtu4gqrKb
rjHpF6CKoaLu5UVuYyxZ+9F1Enhlm2YfaSarVaMVSY6qz7SCLDUgWWboBFTqeozmRO4Kxfbo2XZJ
kSxvIFcwI5YYqw8Zrwzs3HTwzXFFaucOjlrB9gZHussh8QZm96FJ5U7WP+K9hvOlLFzHc1gDstFz
dJhjmjGaxbJ+bFqyOC9OeiD9BXuYQ0zm8S5xLFixAkhRPs0Cp9wwf/wIHHYdVdEV3dPYt0ymmHBF
s5j7WRNRn2isIVD5oG/ccF6+aXipJuan/PFj0vA1JyE+2nMOLGGp4h34OdEu4VNvn/QfufxmwTCo
890CF1Bs6JOz/w8KXSJu3eLZ2AQqBaMB8Dq3yNl8GJh/2WchKdenH2FfZbcOON6z0s9H/Fra0iAy
yiSyEU+BZ/Hj3lpqcOR32a0w8VJY5MzRhdUGOkml+YcsCor8AtJmRZF5rUZ7r7r+fE2db1Gjl4M5
QqYN99dVGLyC2cIZxI5rxrvLxjQiONha3pVosMv031LO+jBbJsUTkMVI5KoHVixxzS3DHk6gwoJE
LBDdEsU/JcShMATaOAE6nxuYDgrPh3X8eGDZLmBpq2lJrza4uJgU9VTHIfWwspfP7Iq1EHtUea8O
dfDPt6fD146xYtw5aia788zGS64r7NXknsWCdIhkYzW/ZqQKBP/NOEjE8dCoMzEwu2tx6pSetHek
mgyjvjeAO0TLEeCcV0S916WmUAvbgqi0Bje/qN8Qov+cw/Rg2LofKgEJ7UGZ7dCzOaqSutnQCcm2
t02qZgVkModsiacThLU20e4/PJKRrZVD4uaeMU6rRgOYLaRa0A9zjBTMQnUvN6BS+A/Fi7mlQN28
x7u2wX4ZJO+VpkEVS769B+aZCIZfh7q5dYHxitshR38LH60y0mjsgiKE1xgbPBCbEYPsy/cFt1vw
hdtJ47+UOCmKQtNQaZqkxo0EDhghozqMJiBQAPIwuRb5oNVwF/XzUL/33Tav7qr7RWPlxdp/8l0D
cqPK2e2JTPyU9DTph4WD5p7CVa8a/1YCEO4mMl7/7jmUo+AnYrEfNDX+lXEnbRi1Cpp42k4qxAdR
A4QD+EohH1Rw36HqrNjw6U+K4kdOnn/brfLzFTTA9a+ckpAEaZhnjpxqaUxkbBRCInBTCqMQektF
osBGMem1EfKhC2dbBvO4MCOAYPA6UUtjh1DLcENIkDN1tWYSo2bdLGlEWg/ddpPqpCK8Qd8lKOaz
9xAJ5MAjunYMR/4YJdW6urELCucBQDKfKQ1jVPj/bM/ygXdoVwvr4wbLxi/GGeYf0XrccpPqVXHz
A0uolWj9q/229nBFH0F7Yo+krTV6rig0fxR5vEFPISzt63VqFE/74DvTAwMPW6HaTz4bA+vvaza/
gGgRFqZr0/PZ6aYEn4joXZwdq7VsR21rZJ9x55JBkB9UMobRwsfs/Nia+k8TrUnL+Kb2Dm/Gk3F3
LFRdWk/vtBrWDk5GPpz9sgYCypJru5rQYnGNluNltK8hdYjG74S74B8buykqvonLrTHglIYmrRw+
oWeO5vAk5+M793Bo+fob49VLwY7WXxKPoT/H+SQ6pxmAl4r3NuhRC5uhqkimtl3FvdON7LL4a44D
R96HgpE5W32/FALBH1S1ORBYrZv9KBqgNzPKYtfE2gJBQdsIOG8vIF8bSeErJSw82WIGIp/9XZ0a
AOlv78fqpDGcAynDAdHUnbTjTQNu5j48k5LlvbhKpbbcvAYi9Qd5YK9uM9q6iVR4J0YE6GXQhCeg
5+g34djigdZUi9TETVxBVx2vCgXY5L+IbaCwffxycmLtTX9Q2xn2uZtRgmZhzEx1HRUi+04bV4Zt
Ku3zPdyyX1sa0ijKVYTLO2vzwXsBkXsqwSoFWYKIrOMFv8tkamxnmR5Brz5D2R4U8qe9E10Lqywy
3emW/Qp/r/c7mwp08riCRXB0Hxj+4ayLNbbSUofNoEr9X/fO6qmMMfaZCA3QewzHM5Upm1KXwQhA
irHbWl6YaXJ9/ccLSBnmEhHNqtpkpu1xu6G43tA1S1D1hI7d03rLKw7cKRJek++4kFi+ihTXpxYe
ExRnjJSTYCD931ljtd161YYot70iW9G1wxTTWIkKlII9EfLaZAq01GE5/YnCUU59CraZacHChUus
69TogU4uMzPfhnuJVHTO2HIvabtIgCFcJ4UiNc8tR5nJrda0eKbeEWfPd6GrYTuK/rjMkqm7Tgey
7K7Aoj7xa5Oj2L0AtagLCKJ/B6xjvYg2IKcJHlRANNb6Vljdqsb8SYDCJkd9OE8IbIwZO8swcqs/
+UNB1fLBErECVeOLz69buIEE4uTgkY0jxbqz7iII8tPr0tgYA6ozBo+WoSzAw+TbH8HGKUwSgrat
ckuPjDYyBPf0f6Fs2M7c3MG/lc11OhutJToLCWjgsjWwgqpeF8ZyMgG0MtkeE3V6kDzlToGFa4ZY
Ha0SYlu37o8YWhrm7Qz6i0yIhtK1w1goHYYlKjBfX1Rc9v7PpNouen8IjuBCbcIVRN9I1LDms3WN
V2pDQ6sAHGi+TQtVZlht8C6mpjUpSu6wfSCOPsjLJQ0R+Env55rSWB5ZhyofxOSKbzceYS9g3IyD
ihmCFFMzPxC1/7KQmzTLa2d6Fr2CHi97Wa6auQdXOGu34FYqgZEPP23BsHuHxhM7oQ/XD/zLmXLy
nBtEn+zd7ahIwe6Rn3oTICJksc2mlzbweu1Vtvl4rMbKCzZD7NS8/BUcw1H7gVaU/ETGvWHIffaw
YDFlADO29/yuugWh3RIDm0pm8bOsxkc7eib1qET7fr+T10FkF2Iljzk5HbVM3GQ/OiO4Xj/ZUYmn
vjRnhlAELQX8hV6NenRc0rTN0HSjZpEAlrOpNX+1FSTGVi3z1h7puQXjREXxQh46roysZY0bZqVF
AiboctLXPw0BPoeP5igzfdrFaFWNgXxavl0B57CuzlNEi2EHsjAMcHCnLReigG3xpFGcCPs4ldtA
fF4RQLGpscGJi6k+3XGlWVOOFJYiSvzgiXF4rHNEN0avKfw1rKvHGhP1M/VI7Uqh2+HKiZbqSbGA
sa+259cbxXqYfu4ChWx1yjH7riwcDbieLEgok6rkYgul4KmQGkO7/5lRxEBt0uuRsOMMSW8fzK3w
YNC/Syv7ZQPivyuyzENh6A1VfgpULDl7aXgRb4jR4qEJvutgZnFwXmuoUf0HZf40ifqYp+ITpjiS
6A2HDdweuENF98qnJxehUn5k9BnxW6kNlaK0n0oQvQNbpYDDYZDrWrqpSP3jC9qWXx92248KemDe
gaXYmuWCdPu8tKdNyNKXKDIUaDqt7GrPLxFL+NP5A9mbmjV3xw7RU35oiCRo+dwZxFxiYF7fWe/L
K00LeKPRgCeEWvfv4JQodCyg5t5mLDOMSuUIoR3oEDR6W3PBVzLKlWXaTGhXTnaEXBzpbXx9Y5z3
LyKwwSGMWgMC0tQYyVoDibHq+c/9AsnAGhXmUzbm9C3OW5XVcK6L62dygQdqgfR6S/FXKsIyRQNC
C8+kjyFdUwo2/r8skj44jPlI553KdscS4/yf0Xf+IIxZpfGmOUhckKUIu/2jTzdav353lF44A408
WIfHINFyDaRI2KzjNez5bYkdqaNiT8+oXEuj8015P7wUusxZ2aYC3KImP+kZgTS+B5Il05YZiFVE
5NgdSd4UXVReFM3j2H0nXcQNcddWVUR0//xcUv3PuIwIPpKv80uJil1cFe75HEECyItB91q7vk9R
2Yr31vYhuI2ghzOieujRjBUzpN+TklT52ajoJqoLC1NYzwt9/zZEaEAVJkdR9AAIa+slQYG9d6ng
yCogP9KliNHClj3yWoKdS3POwYika53gyBxYdIbF+qCZFSH+KluXHUqRJ6iLqiocOjo8Ppr00teV
IiLZ4AP9eL8tJ42lDin0wfmxhPegO5Kc+e1OeV6SHEV7vRtqeL67Fy7GrgNtxLAqRHF7hFz1GNpq
phcTwjcutwLTfN66JBbjqsuRckpnKqxQX8zttqAo94UcOgYtKGEwVx7M0guhADm5YV3dVnONJExC
CtaKs04LL1Zt3dCCpBWG/fdJmx38SbRs2wZfWIjk7CefZMNHSWLS/pSTmRKD1nDykfVwHt6QgOI5
5D97nWDuqLisktMz9eQnQ9fM+80x7JHvsPtR9OJpntcSzqoqypyGnFL20K3IRixPDTnXmNZ5uZ8S
v21KVyN51kPLa/aJTWG84v+4ZN59Hif8aa2ev3EM82AmoX4ftwLGGGxUU+OHye7phySGhW2S8Wtm
DjbhJf0o9Nv4AfniOuno5HFSJs5D0pTD430buW7QdH14SmPZVQqnYZPCMRhwbAWOCa8RfO0Vslee
BrZi2LplC6Vo5KqR8iWDsDcVeLXoqsNTwd1qevto5XKgDh358aUKsr9B22xeZ4nsmuvtH4yZd2X3
y/SSVTprtwzQDF3OSU1DGUl5LGruHuGUvaPZ7ETzdWEvHZ4pDC9E28rPkog7nyQZtPA1GmpcN8HJ
j8/2rc/K3oZ0LXJwzFRhagGGV20GldKIx1Rw//5lThBXILmjp/aOzwsOpz3UTEGwBxNchAPn8nj0
GWRHbpA2LlkxDZ4GSjMfOzDZqSObLq0bLpvZGqebJEhQespd2RcgwWTOzPvQK1D1M2K1V3UmMYyI
DwyCg0jrUx+fHZb/MjfLAtw+YdTwTqdKmqfVUoxV0te/msAXHkusAMeEZ1Cmsb4h55eFG6kQHUv6
AorZGXTK17a/Apqw6gpTd5exiUeQwmjyhJpGbz9aBfwaMg7IJCgAkbXqdm23W74C6oj4aBxeRQau
/vBnAWqaVBP9p7pAuxEZZozu4RgujYuHcDHiLHDmcaEjQxYVOetGuf31lIYQo7tuhCLQGvOh3vcx
589jjbIFPRutcOZ05MPPQGWi4f8jgZrzK5lmYjIxh+mkSojSZoGjATvSrVTc8LgYFArzaifiK4WN
sVq/CAOwGuDUCcN6B/w3Mgjnt3PZINFRCqLzSrxgvJpWYFPZw2w9Lftb4c4lnOewjB4vvXVfaYHc
VUGULdWjbsmCJ1/FGSbsuc+OamsFibzh/0r2H3xWKrmlHDy2jn6PohKDxVmAYsXfs+DimwQvw4yZ
1PjRYjW2U6PtNvehcZ82jMGvYG1+aA4OffaqOhXSxqbKcmYHYZlbQ4PV+DNjRa7xiiWR7/mNj6c3
1GT94t6Klj0BmbWbD7QXlUV/FoPhckvkj0MLeX/n+HIddMJtU8jYlOxg/DSBIkYOMIuEh38VmNjr
93fS73Rat/HlsPdsWlI6wfI6XFSTSStiauC9NJWG0D3NDevBSxgDvZofAs8Ocrxw9Fy/21+ht4S+
d1EbMqZFYDzh1ZZpKTVJX5Cbt8HxleNqC9JwGDDyBJWRc8WEbNyAb7o17kJ/3tZDFt9Mia4AKs3E
VBCSGc43sIkXhJc3XZ+SLDp16dLV/Ef/kEQSvR6FX4fpkds4kSATfWjI19axch9Le5BqnpVoCuxa
cjNk0K+Y7kyom53d2WAlmGxFCDVnnwqt3TqOlJKq+CH/L+OZwHXK6aJzYX1JDqbWJgAgcWOL2InW
H9VeQNjqoB6lHFe/AG2A3PYxB+SUaLrB1wbMZiycXPMJ7XkPUCbLdDJxibmqcUeLAED7443OAzQH
0wR3v3WAVpwMNcCrEmSeoQAwuK/6MvzJxOV+VDmXJql8adhmqYxddXdZnAyxD23wLRlWEzpCOznF
JjIvTxJd1jOufXqgTzf/ce0iJwI/STTHn8xet+GjyVt67sunC89sRxlqhUTTGf9nvLQkOhKBdXKN
+B6NuW8NSaMI/f5IcBYGbd3CEseVRJFa4Z3fkX2CBWLGQqRCpq4SqTuzR+qj3BqhTCigqlKdDQpH
QFUq0RwnG+ls/VnqtYFaRTwpj9qz/SPBlhol92hQT0A3FmlqSnM2ldMaQGL9Eqb+wGIjVX7cgS6n
/HLVmhaekVUny+C0/8u8It8tRqcGTMDDG1xANpXcjU1Et4G3zK4kVhlIsRe9p9k0Fus0obMIA7PD
laElFamBXgV42LPmflCeXiBaEBReUyDZqq33BgyBVh0Ev1GGug4n4e82ZaACxGGVHF7ntkETVclo
9qLbm8DAUkwO1Ao9+8/3ZdGu2qam+pO3jIlWmwdsvboLFLNXRi+V9WlcyRF/E0fzJVFkWMBSKcpp
K8xKf16M36U5TzrCAiSxCPLGLtpbDUPokAUKDdKY2za0AJlQeiSFDSVjdz6gRwo2ZK9KhOlU9Av2
zpxiC/2au91ogJdHW1yTpiCd3u6+UYNKBvdg/gT4Bxke1+IFBjrFG5EZZKTZ/M6+iF9v9Y5xoyrL
KVfivpAVH2LF+YVSbUGcOwMSpXcJfq8dRceJk/qy2BeaIkEK4CwAPONWGJeehaakk7XAKqWbaZbZ
FVH6sjFrKrf9Jt4IhtkRN7zydljAkUqvmpNNSJpmyQNb8omQaP9cib37oPxn1KhndRWsN3mb/0EO
tw+bqS6A8vqHj9Av+NdEAX50aM6556qMaT7V1dp1emt0gHk2HRi7NgBc8D6DnelZM22PQt+RuWrR
Dfea2PNkBNn2UHJOQQoJkqC8JiUHKV4t5UQ9Xd2CC6sWGAUFU1w4M+7CIDohlY3HIH6baotEJU8g
xufLFVTvMAzoH+cyb6uHiHd7NLUt4j69BsvZBdahM6+7na0lIlGkhrghbF6d/BGPTJmemuSRLfEo
2+3wgRNOKbe82xNBCgE/wkBgVECFH1ZDtMWoe9dnG0kaws2+VvY6LnExONLjHor3ghaKLt1vrjqU
GnfmlP0OF4PJ2IriZvGY4PwYGwTKVl9sda3N0J6yTCARjBUEsvcRaogUnIAMqECQkR0RJl0rPCx3
g5uvc6/NRHPz7VRYJRSdgNjkHQ7tJ2D2pBDyiv9Xip4m42hNgPwVDJgevZHDjizTILH+r8ci+4Qp
gnQQSEjux3DKSIqHP2im6OnolKAfclz5NG/S/HWJZZTIpz/bmuYR3k1aHmDEfuNEmsykKVQ8ARIs
Dmu2QQUr5PBM0+VYAub/4/5UDZXlLk4HGWB0FuIwhcv8AQq7H2jtnxkynbqqoMO+nu5mob7fMcVF
ntdRgCqh43FNYmJEmZeLOLR56edHgo5ee1gch0qmCfx/eK/MOQlTVDcuywPmG088b/WLJiGpJ7lv
a/Q5k4+RLPT5lirdeD5SYUJrsnvB5fPe7yzPDYvFFEFGXVURB5AnDOA1RZumrHPG7RYvUUcHUka3
igmawwyB1JQ/W10FCFB9iWv4mznjtdF5oidaDwPZDviFr2e+YYgWdoVPd9HWCp2Yt4XbA2nCYoJ4
560+FrIGvepAePCCdySAiVpegtnHVsGk2vXmbuf8PFTSOsEpfsHAtrNppwBQrT3/0eBf7EkUMe2s
abJq6hTaFayqTp2DKme0I4I4rLSwWssOeH0ESeLIjWpow+JtlLXCmUIH0mLt82fO9SebL3lXwhUM
Gg8uDIVCxU5VKkAJeEBkwnx5vwNfHUQOxbTckOJc2XKM/cC3rC5v9LK4189mSJIUWtbroIs1urY/
qOts+mWVkLYY8sPsE5ub9UN6T0QISSOgRPKKStLTTWbRCqz0OrMK231lZUU1PKyhKCARPNK/8izF
HZr9tHZ2vwm0oZ7wcMqujKopImCtE5T5TX0wXI1nzmCvmbAq+JMMGvmPUeqZPtSQOG9FqETzx/sK
WbRt+20q/hkq9AjagXJrwH48L1J1k/3jLmyzFfj0eM9T+ABWvGHegDmjg1wu3kU0RQZ/7Kk9I8mA
Kt8eq1c4zQE2pFbkYNftVPam7oLQ9uq5twWdsACIoyydSxwApp3wUxx3M9gMfdpPPpFP2g+B5fEs
L65kBfGgNx2wx5eEAGFmus2ejtRm0cNBTRwko/iNm/x0XILtShRqhglx1OvVF/boGUoAbUu+rVie
jlEWO5a9j4Gb9L5sVmxK+fSVztUrX6526nKKFXr3X0lMeE/u/YHhARgZ1llBJBLtMHVZFOvYh7wK
3cCySDrHwhoftK4TE5NlwCPcsMzqAo5kuUtP4cpiq/1bhmEzI8o2VI+qZzQbZ796jTLkxWrvFkOk
+0J35WIfmx20V5tb/q8nxP8rV65esHnBplU8039utCDdFCPS6/+ZH/X0yycwkOf4Qngx42l/jTb0
HkiiLF7iLZgc+ppMUfGP3M/vKNbRIMZ3kZSkgZnPnxHBj1C4apoTecT3NL+Yl/sU+VX9r7LJUlxy
43lblj8uzkOwcNYlYg7ltBVQKRlzsUYBq4R//xDx+Pq1GPcDKPHPspL/aO165StVT9SWTPUaaSu6
lrTNeXxaCVOWRJjJMMFoW9UC7iaqHSdJIuTHdRbZC8gdrd2wP/MpiJG5gLWZk/lB9z5T95cqinyi
LqP9oFlJitjis3kPcq+SnI5L2t8IhOwX3nX1TjovIxcXy37EEj1B7+zY1dp4e9i8k2o2rXU1dwIV
WtUIP6ByqT/itzn2mISmptj9JHKwLZlQ4itA2QyNUmwNvLfFv+RLb02BkEwnryHpRce2MV57uUK2
YOJiJM/rSYmhWzN3i7x1SFPVv5MwrYDENsySpEvdjxOXdS1HMqjnuJf/+pPYTmeSINOQFgEothgD
kJs+6GJlJ60oJRQ+0ZRvIOwcxaSi/NWhuLt9rOEcEwbx/7UMfZpkYlIe5F4ebOTskUuNWoJMFGIl
BUo8j8zhG6FkhnKXjNDuyoFF4QipJJSucHDvBBzYXP4TAp4ieD1xn3b2kQaGUCQZTB1+8ClUnjow
4nE5ZbX3g/65RWJ5orqS065LCP1ueN7REvKmThxrmT5QG2f9A+k8q1OuQAOu2xQbvQ1HwSbtHCt7
MjPuonUIS5udByAVi52HPmM8xCrUmUbiuQzJelUvsOPWeb3XBUi98+gewu3o8H4PC13kYrWUThEJ
i44GyY3tDpt2jdQc/+mS7yLXnSzhw1Jmcdk8aj+s/896Eg1qbx8U2lyS2wy5nmWMG2HqvHOpzxHF
nvV/Hzu05EgHY7bYMdGWmwgTwiMYr1VHaEDCGR7o1aCHsthRPVWekIBVtZ4Avv2SF8eCyGam+v89
3JJRENYBrW8A+xGE/2pMaNqWPeQB747T3gnyOJgn/XVdxMzFt3ubXAz1Xq/blz1KDFFEJx+j5Rlt
G89QM8FKe6/Zv4ibw/miI7Ipz7pk61qeHJAzhgkceO92Uk/11+T/MIsXUQ9z2QL69k7VMjitgvph
9TdhYxNnTJuFfqV9h0pwiKS2pyw9bpe+v1EaUZKypnh3UbI1bIBwClRdgsCYqNQZxp4uTVxNA/XT
T++l7GIngZmDkbJsX0XtQz2aGn3S+EeF3yVnrcy/iKBX/Xo3yHZAW2oUqhVbI5yhZ+Zo5O4jsrdi
YLOI3tuJl1A+CAeo+0wo+iHAa/13Ap0fywS15I/LY2S9NrFDNv5/6ljXlHB1onxILqH0iBbLjDca
hXrIrFWG3bUhQw2wYmr69p2eXMdRT+I0AXkMFjlXlWfo9O5UcM/tPv5xgm1jyFs7ARq3OzazI5Ho
xeug7Oicl4FtnGvqAZoEEksGjjsjZMNEG5I/d9QplqnVSMTs0mTp6ej4XNYFge4KZ/TKufwu5cdZ
HNNg5kBTN2e695/xPhdUG/G8s5giQ/gcr7EfNsY3283n6rY2rr7VfQesNrPxfJp3pF97Bq+7/HkN
JdPXfflKNVdggYyszcR1tquGuU6m0a2Rszt8RpKQt6n2o1UNhQPFYlQFN59uxQPvla4IR2LTeArX
XvrXjiCPl0HZCNS5vAK80ddxz9lCYvEMfB1wfD0JIgYL/ugEJU3iaf7mn3SrGy+QRfGIWSq+U0bZ
lKooweipwSIioLR1SiVB6vr/gP5YiHPwFQeZqmO5/ijGhIrYbAU/6hEwyDHaq0625u439w1SZqxd
by73FgQmrN70xPM5EYxoI7AcO3l2O3H5WEG38oZpHjgjVGUyt8ZZNd1E8cRybNX3R72jnVb3Wsdl
W0r9R9otZdmkAXg5yD2DAKs/9cxPG8odlZJC9aamTdy7KeWABrLLmLD/P7UDwbdO62fyPbLjQuXh
xAtCei1mbiMxTsbreiMyPwzez0YorfpAS5RPqtjfE8A5GX1+ZL3eAxbFNLEJ5tADDxKJ7by3I2x0
wm/fz8Js649X21vJlv4Zls+cb/3m+dxyksG3kh6Tp2+/DsOkExhMdwXL32LTskIzwMbe7yr8IxB0
c4g2TSV8UaAPNTkH5hVXjxYetWF4jHvL7LC+9bDL6Tx7oNHXhWn3lEH5bwlAU5+gJUcu5zlcCAgI
Tax1bA8rP8jNra764G1ITBH5xgoIa9Io3/r+EyfaRYi8uX1NYKyhQz5F74v8GRwrCJN33geLtX0R
5LDjhqB2yxSs3KBPFL43gr/NWat8VpS2Z42sL5Lsp5MmzCyrON3UtHw7FNoLl+/lIOCRBAlqGpD5
+SMUg8nEYJsJMhPJ6ThlTu2riq7s82ghZCsmTecf1XdTUnQ+JVhzATCMZzu+aaBGmx3dQcpn9WQE
LR9FYraJM+SrQOY07vrqj4xUAhFfmyYez5zhO6rIB1y10+0S9sqXyG/g/X4aI8xo4JK29fkE2b8G
7HTiN9Vb3/EdlKU1OgeELEHv/Mjuj5SjALbvkhXxF0pGPl9/Riueur9typoUm8eDjyZ0S27DNGK5
yrLNjSBVedcYxpsz9py/7IxBIexa3pJ9K8M+CcCoNj6vpNJ7QSXs+shRg9CvJt7uzmy0QuU81qwj
bO2OWzw0w8+iu0uzDjFSNSNdQOePwP4B1Gt0e+0S4oCA2LgN/GV6Erla9RWypE621UZpYWP/T1Mi
WwgOuaVXCVWRZoCZivM546b6oFysYrTTJNpSrcNpyPZFWU4q2fJME/Tr1MC5f11bE9gEteVT5jEf
FO6YS2RGF7O2pDDAI4w388PvvSOmFVb7v//HSJVjyFGnzpZ1rVkMsVFtR7LyZiJtv6OnOSRk3vSW
TAi1p6bo4kGY3Zy3MSD0vMPWuqK135/1EkyY6kW2ksXsIxaGZU14DR+pPHOI8BouM1lGSSkwCpZh
7rrGfEhopVvdy4TDjNxqpKR5icKHe+dweAtz0ORaySuyuzwN8RJYcACysfTt5SoKqg5sNYpFFVMz
YAP3sJKf4gu0FPyPdcNhDXhNjYsGIHk3Oy44s9mhnhQMLK2K8/D8JgE/9taD74Ocds6QT/fg/PU7
xDFEqRsLTVkxLPb/Dyb7O9OlsDvp5q/n7z84M1bcCGKFA4LGLXg8P7Bmfm47XKwl/CFXo28WS1vt
jHErgaQF8OgsUuNBBRUKocXeqREDeHl9BkLU2OrVt1yLThBm2fI7haUzx5aHtosrUHOUO8yp9Ijc
4wKkK7ADVHy2sU/vvDkkvDOVaSWCwkcOajGfwBIdM/M0kwhHQLVKvB1j4RyH+7ssSixk3x0szRgp
Un8/2nuAX4vZzF0RtSju012W6oJFKi0xJdrnOtBv2oDSBvcDyXQml7Zew625lKnPLb5g0OK00+h0
BIhGiRc8EQDAtBqyO6kYvGU5o3t+DUbhYnHCYYkPB1oho+kQkehb7+4p0OG9jxWVm32xV/Y2aJKQ
vpzX2WACtqFWk45Kw//m1Il2GGiY8CAauXfQkxjvOQ5/vdGv9QhoZAMpKp/Ktd+jOQIgElfGBBEJ
0E2JQmqezrhwYCZcCdd7524N/GzFdw0ackcSukIt7BM7KmYvEMe/pq92Bblle4hREKhGbf691RqN
JLiCyUhTxHMmnkNynj6UEvFb476pxPUXk8BXXW0Mz+mlnKHFDSBctXcwTo05PSu3ojtPB4LQcQ3z
xQ4Be+OyKsq4HkO1bEXikR11nQmebLxprZKdzfXnZgUdIpeAqRx5uTYewj6spJN8E+IcSQkToZJ7
vCP/gvYZSQzLfsCQhs2HAdpgi7cTrBRntUE+qh1KWjfs6pQfJlTCzAgsuhx7MW/vbQxb7jbpak2I
5DyO8BoqkWG/4fVuRu/AFEaj0aAYA6GNuKJ0GluX1ePJWCX69Rikydwy69zYpJ0cWBe9CmEiRdD5
JpCvRr9zLNxeGcmCmUnrPjQDN3FHgSXXyrgsu2L9rjOA8mvnkhlEfD40WaXj6yNgdQU76KPSW503
kMA/9cgaQMcgwHSr2wtSjZBhn7TEoNgWB1SjJZOX6L/J0qBfrhBNhRE+Ki41U5LsmbSkarYsqXh4
Vy+6fR52njE1YBXQVUJ3qq31gMrtF3uAtJ26dmGY3G/cXmrCxo/vvY1etXkqHlV1qbbDqReNCGkU
lzQP73lIjEhxROm2yxJuWc6GvPf34hMyvcsUFc28n/ID88L0jt6DApD2odaLHCwV146i1CGUC6dJ
SKOPLJRTzc4+i6Fz/HrmNP2e4aaTV8TEfdFgH7kdyMq2kcEtnk8wwpzvEcPnFCuuivpWoq6t7Txw
Wh/hgvD233HMheEpj1ZTDXWH/ks2y66oaoZpEHCmd0xRK/aTPcy1G9ycv/wkg1wpREs8fBFecK15
Qvsx56GaxIzKeEPAARvqN3piTVGWTViBnd1/E0R9zDS8vmScKGgkMyjbxxbgv+PjNg7/j09bJJLT
bwwmVuZKkaDLQLbdyiDXtnidQysZ/3ljDVl9sOXMEuqfIQ8x9v6ygK8g68kvOLAhRbsLwqsBvovS
mB+AZwF/2isxGHeSZ5gvycIU8WHV3aYSHJAvr0DYJplD9c/FCtmeAbBxZKIw/jlmqF/Dce9MOODk
tC/UgOmtAnn0d4A/d6+ZJ/d575eflAEyyLPrAaoT07zaGz6e22wo1IP4kzalAPqt61HG65aZeqS8
nvTLdRRF2obbtiKbt4b9A2+bH2OUkAlpTAhcEnsPNZJK4pO/VXmoUZkQB//cXNIQKNNlkacb04hg
caF/tDdW/ESut6zWeVTe7sefBVFV+RZxV8242J5RteZ/RyVoZcC3GNoNUjixhztWSVn6q6bK8QE4
qrchyqfmFV1F+lDtdaQfSC/kdMoJARav0KoPajyvhHLKnxCiR6zxDOH0UEKrH+kSM5Lp47XrU+5S
doc+MGuJx4Rfni2k9nnngn7/2xcKyL9jQuZ8u5AYn+5MGOSrUjVut6wrAv8v+MFxoprd8Y3n+jIg
cL/N++XLcrLsMKTT2JSfUqq1WBxeiOTVlqnii1dDFwsdV1rARzQK3rdosUiAtCXu8537vqsgYBV6
I1JfHmGyF0o+KjoAMxLw/Kkk7JrEG21TBpW7mx2kfrSJjZ3p+HSCid+06Vrcjx24ffUphL3SbmH5
9MLdBAAey4OHMhbOSbrD5xgBwoMLpphA51jyfk/f03DpzU5yrKW/avsldfjl5n1jU5dYPnO3RkEW
MZtSDLYbhJYnTJmCCCGoEcwyJcZ+Mel4LWPl4f1yCgnNe8c8lV3MAmOfgijlKddPsVxtQo+H1G4a
bOYEVaNY5yb2ZeGASvsZkSE+JdacxrnfmpxBWwSaiv3fl6cfKdzaM6n4JZwF9M7Toeor74xTMYxF
TnG2BVomngHbZvl4bUx+0MgGIhaDn4RHOczN0RlRxddURORZBaVpWfi0KeWKXGxae1bWxnbBrc7F
QcPWIHvufS6gZHBA/OBxjLbYb716wg99TjxXwtMXo4MIcGfZlfezb40RH34OFip9ncnqvHdA2/ev
J7Zm3sKz0ZGPunTDEhIrk97tG+9DTD62HjAo8tHXmt7WYgaYt1lplvswyVWkhMo6nF3sZkH06Doa
Iu1H840r1e737nH3iQdL2byLUU/mTKhLwK611IT2tJMLLHc71QfYwCy2ERJ/BEPXcCalT9nNpeau
+MNCCu/Uu3IZ5brPquY7GJdJcR9jBulZK/GB9c7tTP61+naafIe/FU9HqgrtbtD0pK6uJQ2ALrIC
0ETAZSHBGpmcoeLhD0jAwbYAUZVRHZI9fBWVtfrtLxcRR5QfaLYjKBrij+RBPx7ym16/2CmLzxc3
IFGM/Q0t/uFC16iMvJVguKdUT7HYiIQ1iKit6nnyHYdxCrizGdN2LcxMS3d1FSzxAAxF4Nfzy8Do
up4bytGO2SdgNYAe9XWiyw4KTV/VNvtEVE3iLELr/TjGg6k1G/6WoBZSxfknakZtJf74SEL1MIQT
frIEIlDxSjb9h68bPPY2zhOA4OTdTCsVo5bLuWVUW/RfPrIumrvVFP40CevpPBzCIudPPihqdoXL
p64EWLp5Me1NIEQ2d05EQ3mgfXEBfvsTXn5RQ3Ps9xbnM6MQIU9IHJc/A0S6VEwSyiEJrk/ZyZwg
dn81uo+ibzKxPnRsiRJRM/1EuSQOaRSQc6x45ywnOZ2xw9b1mM7eNJsx3if0Io2f5ZBVmRFfPSkD
5ZuwdSjU7dfWXLJefhgHAKMnYE6JqJdTthqJkpRc6wppT2r5I8iBgRjMBB5qTUIWSwKtVFLk85VY
kVrexNoy2UFvu+erW0Mh91XD1OkSr8K4v73OUPdnhYFJa93GtRZ65MECIHBNgdtTK05KJ65kLyoU
PU8roKcE49VAnykjkK6HEqxCC48qRQGuYmrrTo+FVH6Cs4Zjj9HKWcA3o84R54WzoTrAGQ16/OM+
NzjoXfXvlth7EW6P6Zmv5HIHoW0glzt/Klm6O0EJ+zdR2OSPc9lf7AX+brDBPu+8IderxA4B432/
sgTwkpTl29kkUxSU8DwqVorxDeQhBusMv1sRJf0HdSgIAN2lXFAtSrVSrPmDrQN/mSHbswa8joNZ
yVwgPo0db+Rdu7ar1WFb+9ujcxNMB8a/5uxMa1RNLzjEXYwsjUxr7hnYI71x0QURTk+99nijSPdN
yG80RgRtUzmEHf6/hLesNsfhLLJxxemxvYh/nEfvptb2u2C+HegsWkWG2qf6zYcxDHmSwgsKEw2X
PLIssUCx21aQU8EjoMyw1s1lb1mY1SBClGFZMEA9FjALPO6gUFgqc/Q4LThR+r5CiyySO7AmSjiR
PVOfNLqnGGouxn/YSlT34FeRICs2gsOJI3hAevTfbqsaeAXDxg/42eGNksMEoj9ZOun0n33wQKam
hiT2owyWUPyAbl+BBrZR0jmHN0Ke9yAT8tEjwCt/qs8UDS4bJGZIrn4pDBb+WOUZ1N1pNM9scqw/
m9d1saE3A/chsnQ1uOLlRiyOCUAPfigSN8gUxa4nmt/OWOsEEpS9lunb+HqRs84FXgN5GPNVhSKa
aak0AW3nhnZvMe4+mY0UZ1V50fu77a9YjDV2K1Xn2BnlIXVYGBty6Tgq3Mk9FYGMhiP68Rt83Dkc
8OcTGGR/lARJQU8Didygv9D9xeyAXek4AoPzM1MCsAphIAyU8f3jTrY0HWfOhQkz4+07DpVmpHu/
4RzOczNKrMQqLOie5BgWpdpeFQ9H7UXbsGwYm25JtIpj7HeMwBweupcAGpWoFp6t5r6kXDmRaDVl
7htq0kSy3CIwiAPdjJqtsobNfiGyI4lYuX9dx8DH/+jxni9YhewlKa8otjiAQukU1imjrIfLn/A0
59rgJ/7t1iYXU3YbwUHOnOCfulTC7FJvE7Z084QsDY6QQqaumQdV32GOLnUdpxgugZtY2v/Mdou5
y3ytY709Q0pTPl4Q33mq7XZ7BE7/M8vb2TLayZ195nwdGukkrMEmOA/IQxrUCoeQ0HpwwIa9MWAi
oxPiyB8NXJUNNDrJrrQ+BCNJiQV3GuztkhJZyHBpV91Qewl1d3e0tAKoYiA+iAKQm8UIE0hg7/Vc
P+hPtXA4QgigqKj4eHd62b/sWPp3FVl4HmW/ZwHF0GdH55tVr0gTOfy7PqWfQXP1LA9NYUqT7VHE
HxVKrFHv8rIKMXdaDh0pKaRzG52Abfvr51foEO6SPWXwSoGARr+MMb0fmuPD/sppPabhzvyi+r1t
nkggMRjjRUu7wLFGtklZ9a6y8Py/ujg1BqBc0sTMavuiIDGGbQ1ZCidKQ77xHfZTTaE8e8j6vkaG
qXkgNtSM1ZUoLOlbrvYCnMuxpnthB7tyNU8+mLEdVGPBjabmNkR0+MU/m4/botv20s7rWZzTnH5Q
YikeOMNuRPwaiaaBajgxGhQWpSQ8Kyt7DHbbW2bPX/Oz+oal9bGqHbTF5cfD3VUZfsTmszgRU410
c/lY5Lt5UEYoQdADySQJoHe0RZSuLxllpJ8lwSH6f+cwtZ9AM/nEn880XaYQlMTtF112QeiLFUH1
bu5wc7+e448uxlgKDYX15dLyFE/Pkch00uEIXhWIN+AnBsNQrTascTFgW1maXb5PbgANvpY+Qiqc
bCy9Sqa9cH/q1/sZnwTeRlFDUmihtDzErDUJdopuyzxARQySZlhmkwUij353HGZCzn18gg3ssT85
0PTmKR3uG4D/dznNpNfpsbJ5Xu4ccFup0zoAGQd92Dr/p1o1AI+8MWEVPe7m1mTwvNlpux83M0dU
9+D5D2O46T/e+MR90DdeKvS8yhavo0RxfLRozbEtDURHpT1heA2OkAB7WRxzQDu33ifcvkhJNTqp
kTB92jOSl60HvOlgJU9YGKc2f4BuZ3GOAoWUpbDG8j8U6xkwU4738ccIqH2K2gO77Z1LW/bfFTU4
PQyZ9g6iMHTZQj7ypLkup18Z0QTXjp5EgXgMIDYwZHH7m6csVBSmlRE8yQ7g2ASqOwkj0GpRBmLV
Ya/dTz3CKb64IVplQPw/7oHEheSgWgawyPuQoDbJJ1DDtTxyUt26aXRb4OchiE8lYndgPW/kXhmI
Fzdg2QBG1y1TGDUuacqMpD2zRuv4bV4DCK6zaQqtf20aj03KUL6W+WkQMTX1pbNWP62bns8ZiS9f
4VU56D3aHU+daoU+fg+44LHFqr92lM2AW5V25zJSTbu3GUg8znX7zxJmqIAiJXhzIGtpSNa3xUL9
AYn14R+eLy0BwzLtxcKOyzLwwf3jW2cLsMY1uIaqBjOVZHUtoy0tkW/CqiepT2JwP6tOTFi8n/yZ
cxXjl77KX9Fh+4MGRtuuXVU/rZvBy6woLSeZZS9J2ud4wC4+0R5EvAjjlBxlSsbyRhmPtAmum6aF
aGqLbO/hs409aSQE8bQaCyx2U0tlzUKsWfRIc0HjWFI1L0BcPVT7IKFPLfOEw3ojmYOvlcaC+qAI
mRVuDkXyswxwPOUsxxK6g2IBk6mK7PplcGf5scjIGDZiAO4oDhBp6qf//pgYNTMKRaMRUOa1ykhO
xs5cMRGDt49KxVx9RIqKNDfKwpohthQ5+4mOnad0wcSsfwWNre0lV8KeaEJMc7OzQJCzJFKLJe9L
GYIEjIgHY3V4QmakMAbnyfgLPQ6VXGiFy+XRBA2mjoa7wbPMczY+XgzOCMIER7Z8vPpgws3ARNcO
rwT3Uaqr1lHeWl3DLV8bdy3tG3gLOttBbBjPXY5mTnXXOA1B8icsGHSX8rkm28RRaU4HRrG3dBDo
taZgd5ehEhtIZm95ZVGJla86tAaxP51RXHLdrCjBh3xRWcjpMMEuawfnCeQjsoU3Mgf/afXfh9se
NAp5EUkwVm+y1jC+uleXIjgwoQUNR3BNcXkURf6rk2d3JHonpSM8S41AhgHvnIFoFaucCp4z2HsC
djPUL3HEN0cO4P2JwTmXB2t9Oa6MAO4MmMGo2RXpNZ1GIcDOSCt/Olv9Y0MplOuABUCq54eq4qQb
qL45/UDdHGkezB4crXTU1t8xiG/f8reeL3oLlw3j6Zg2wsIAu1STyYVGEmShDsAkQ06tZA3PND3P
AdtCBPZ510EcuHfm8PgfVu2HxPhmgGU/SoyuW/WoEhLyGyhk7eYOt3WYIFSmTk0RegLoHYhJsVfE
AzkdSEmZBdeMUMBST7ssbu3bJQMETdsnbuZOzulRYFSIjWi1xjZ8fvRENXSti1qXSUaMVmzNTlOU
OJi11nhmJ7TZTbss2gWkoOO7Ujb5khEcxx8XuBgWuHImNchcqH2/EczLk98j9pvS2AzmHHhF30Ud
ABoHQIiy1vTyHaLm0Oj67DL/xUvGPl4urvuUNNI7UdRUxJ2EBhptfXvMQIom24Z3wIf5dgELyzne
Jn/ARGAmnvRlQY8pQZYGSffp7fI7s+6aXMY2H9TeTZczttM2WSKQ8yd3Qsye/z6ZWd8H1Kj6Q0Lp
xaNr5JKYYPRrys4POWeV4zjUtD4Vp761C9FlJwuAw9GZx6Nl8ugGTJyb+dQ9svEX43vq/p5Qi88O
zo71dIrws/a8OcNi6L/P3iXzgDN/8+92Zea1B79FNtmbNgwWxwbtxr/VAqxXkxI3kcHlXsAVZx9U
W86MKBJxv81lmw9/kGShR0CDBlNcgUiFeWC67omRYqHFet6aFWNX3OP3eVlQWHD0AwomqpanHkTP
Bg16QU900j3vESgg6cxUBmRg8GCqvY89sy3FaVuCCet1Y4FpnSRTkc4Bz8/bxn0zRQcaKYKQbhbe
g7F9o2UmNHsJJkhiuDDT/flbrrnMtPPC78XKf4wefJr1SaCM06carADUfyzCZA5fzqDlqROLYuYV
E9q8t4cLnF+u7xUA0rKfbkZf56g5YvL339U2lnKrEYJQkf8HXCI68bImDvarUjh6BCdwvAxpEcuR
F04Ukv87unlFVrEToIWoyoWUkN4yVxz5JK4e1HzQli7oxOcAattkEuyr9J3Mzu/5gqmetCxhCDXm
8Q3PjaEHNeBvDOm5bPB3+4B7AetSExsR/vRgaGP7lQqyUgZFZ0uwY5V0TAbDk3LXwezM2YG30iOe
jloZ1gzY5YJHdtKX88s/7Yf5fK61FqCo0qAkoQo7DdQiMs0d+J6F6gENW5yIHIgAZl6ZLXs2MTtM
4rdvZPAUtw9NoVzBb6bxkF5okDx8kK+2HaOyTCpIuttyMh/TQvK9F/WiEd/YHQiWZ7KtG41CDuHx
Zir2fVPp/w/E6NUMH7yiAnFWFKEPPFRqVqG7Hu5Cl1LOoE3ygCm474gzutVGiTQA+A/zHwHV9OhC
nVhKpfDPNTy/U4JNG9nEEO+qX1rGYl4BEfpJI/6+4LlcGCXpHsn68hOroDem8zYUata9evo7x1aj
2KcDddYOEe9VIzta48KdWqR8Jr9S7fTjRCeBTYlUVu1eFMQtpMU/yI/tJ9NqNmbd0LELg6WKCzCM
rA8M77O3GNJOQacUBFtOhUo/fqvjrTnzKr92aL4YF1IiU8iS/cU4dAPE4oxomBBRhM3hdZexu9ie
JgBEMWwT66rUiwRaTHIFnY+UZI24S9LP++4owvzTBJu6ctwEbFwOiN57ufU3pVUt+v5I/zQD1Cts
ho3O3aAgxVDhbLNrJX4Ao9/OgaNJKw3QR4VXBHcGo7Dyy+edy+bnHCDIKtmDsytB3Q8yKEd+q7rx
a2g+BPUslt/5YpWCIEYSbK78bAS+831hktol+hAbcmaUVWoJaPt7OwucwL1TkwQgpWGDROcj1vlG
b3kdUsYo0huAfMP11Rzsrdy/WFCcD0oCC9jL+dspRdJCISH3HSkFAh437unmH1UToje5F4nRjSxg
OUuAIYfzC2VcxmmUYDYxIeNuUsuyy75ENfs5eN3jvI/08Nxhs8iZcCEeseH0eIpFAsoqmbayjf9R
EgjAroBEUvOijXFp/ZEdCTp5c7O98Zgimy7TpEFMIPNO1M4G9fAUJZu4L6LyrvPgTXnJx85AhG0U
pwBQvQ0DrUx5AwlSgRj+AmV2HGaYi9q6XeGR2Pwy8l/LLU/n/MXEyfyVUKaY4ijZGzG5tAHF0K3D
ioIqSHzWCXv1t56MekFk6nB9NGg3Lx8sSer5kyOOPR9DgMj7H5ViooJlUHiT+E6NcgO7UsAWagBX
y680x+UuGhxueSo2TpDikTB70yNJ3mApSonSPZk4SEpeYIRCAc7sTptQNcffc7pqfb/pJNY8L2jZ
3Wctw837g2WVL4mA+5g/SfaVp00jv2ngQsF35p8KbWCiuOXeYNyATo54QnzCf3wrRlBVC4y+Q3Eg
SCeZc7mx2HC36zxa4mYIpbOsltXIpvTbq6NWdzenVFfCPsA+A8wXtri/zRabvROUUOJdntU97Yvn
sAU0BJGwQgLF1sBHpvK8ZWZEYAQfloh9/3oNv0QhLp2SFYp1cMECBElzzZm2dUec43fQlKvBbTk3
NW+xlNHGvvcaeVzFoEowAAk2uHgnqPUThjR+ESL8ku/1X6oGhm7oGcKRU9LZflOshNVGPrNWqRYW
Ft6VP1rgKbvON9FeH21cDlZhdXfTrWmROJyND7jpeiuXodKRTVDX3ZOhAXdyQM1zoJR/OIqzQaml
pQ09fwVuVxgXZqCtS8ClgkJW85OnBniD+KdpcTgKqBdvgLNgZG8zJEjidiyfZVa7rbUsbBuAhvtm
ZDq3AnE40aDeM8zTymg/fY0hf5F9EwXsyGP4Zfo6oGiO6Y0R1Me52LWURprWihe3zGyU6rhJbFAi
pY/IsXs260XqcM0Db4R20VgzDt2MD15KCjzTPs0Jdh0KdXc2yc3j6ii2dDqY8A3lVuJdgNLlU5TP
SnPg70saoQ8ZW5J9hJ42vK+9uwxsXq3rst9JrvYxereifxFheevkMk13YsRyFrknF1q6auLaa050
kdXGtH30oUvGulhK9lG5DiH2Gw6FyXqD7u8doyTa/3u2CrwlIgsHDv/ig8XVdfU8VYItC9ASlIBb
V/h9mjHCMZOEzJlLqVGeoBKi2pMIvMaiDQZbBp7RKoDRkz9TXRspjeTWF90VV8Epx2gqpp6hvc9k
EQCg7lFah+WJs2zsfGxBsuwz3SQz0r9567TuBo/I67+6D8XoYIoxXrj9bf639Xr/97NQ/rqMapOz
eSEfJJwU3g7doo5aj6rlD4mBwXcYSlap8lCl81MUV/eXiHkwdT8KLmtOP26iBDmVLucVc7h4nKT6
d1Ju79ctu675CXhTHWknKTMY4NqezNxDqkv56tThpxsHpmiBPWC/IAy3C6V0AlA9rmlFv7tYCsFt
XxDk5vksRNemN/Lmu2Tr4eLkDz4Le2xvkSDIr/kLiVm2XGT+vsh9MyBJbRAeUjtRmrvt/U5VBzAN
hIDOfDz8srJiPX82nQysQ4+wVF4zhnvC1UR/UTLAN851xMeELg0sSvnP3qc1kK/o5QjRM7NDhzQs
vWTHL1TALx3tJ4OJFQLu3p5+wF3CX4F4EziwqGZF9Z/XE8i7k+fyFQh1rcMzp3Eiz5Tb8AMJkixS
QZ6dlqjEGmDJOXtiiLYYK4M+L5P9i7wrbqZJFBLzaFPxeDTxfYb0WhQs/vcCI6phSRZjpb4CHtJG
OUY4a49Fryown88Y23pbM1Z9vzBUi0Xkn7PaNfs9twnqv/UfOEZARY+GlbPTQ2b6lh1ipzaoD6kr
JPfuUBgb5IBPdfbyV0qsAkfhuSQBfy/hO8jDq+CmX7bE/m2HZ05RLqQmOmPmJkaIJKz5tFqNRj2y
ESQz46k4kDbYVvfKjBOuAe9vGKKq6flLgqj6hfX35VYmEQGJiQxMSHkEPjol0Slp/okPRxCN3OU8
R5HsnJduFKTcaSBAJL0oKvfNKdbgvv+om+Dqn+mkcoxK5O7A4C1L8ICu8fDoThPQuSwyc+D8q53O
HXKMQUm2YeKigbBppVCKRH37jVRBNEvzodBHbwTDd0zbb60i/bWP2R3MW+3yoAwryw68fvZ9NlKf
LLHwZzk4iziTChNZBS4Fic8BNcYZCn5AXkQyxIkmcRHctP9FlwqhFRlUrX0C3jVklVcbmuVV0qrc
rz/hHylMOC+nAzTqIutmq8oyaBD9jGJE5/91SvV5J/mCX/RjvoJS0PvkwDlQmwkgja+1qhz4V/kR
dKntGgU/CVdZW7WtGNBk/1+wtqDWCXUdtQHz4K9A87fjS4h/K5gNL7RkezA7lwksyse1nATyT/ME
rHf6VHWSDQzsg3yApPd89L7gck9+Ily3OR1XSGimmQvHsKWfE8KIX/ozKZOXixcWLJ2Rn29rcWdP
/hdmh0JEHldgPLxDXbaqPPs1xaxPtCJ1jVus2Zdmbgn7JcOMSa+yvLC0fKmGCPrTP1j19OD0x5Jz
FxWwW1un9Qq+nKNhvaoARxLkZPVlz3n+nU8U7PkxVVqjQAI0BcMFjod1vj8GkAhab2jk8KI1dHJq
w+L4WEi5UBh8IQ5VerpOUQj1HfD6H23OtdsW0bQY1+Q8vbRJLfKLwnoLw38F8vwErpz3/kji6UEx
hM+BM36Wh2Vwyyfyvu94YCk82VDd2trppku4TaS8xdkA4fFDag/NK0Y6oa68PRFW8w3JjS1gUpng
Dp6RBoGWy1+tReVAx+8kf0L2x2XlHuTtzKJnIB7DOCVhQPxMCYubk15sj+YvSSXuxb1eynK6pTAs
aywkUBVIlacWw/7+5GXgfUz1gdwcux8OXYaNMnjgHrIkOc25HyP8XsHndFtChku1PmUpxPlaXfpG
8+7gRUMcAx3xS2wp5W/Jz/3cwKKYPrOMqE9lPdAWdSB7MqdRB9YuNVcTRCOoLiD5jM0O5Zl+Ybri
swlIrovlIAD4izIprUpy54hhBJmdLS3xDSGvkuJ1EcrZU4+sepTHv8zEDhqMjHoX7xoOGwRVlRzX
vmEMMDlm32VH6xb668eRZ0YRqZmameIcD/jWkQsCWn0vgJCd7YrP2Ux8RBAbtNn7Y+uqgMRlJDYy
QR3+6kxcjts2n2BOzmGMWnVtr0N6gQP/DDhfWceSmhm3nOdTZDVmjVc/bTFlZy3hlfiQ/5MZtWV3
0xfhsopl7dDjeu6icG7vo9YkxN1vWb5ssUknuEFh8BN/dbvSnwPL2i1tgbSPynhOODQ2vBRf6Vkm
5nq4mBsSRC5Wl3NUhZJX159CyNM5w4D8GDQHQk4Ip6JU+GwpC3m8WKou/QZpzSFRVA45AFck5PFP
07mIxmFFL/p1IN895YRXVC5k1jVUvxdUcwll4JlG1HXHXqG/aq8RIA3R8qcVUNj6GDbloCq3Oh+/
S9V2MBJNwF+oMDRBaC6/1i73gvwg7bqdYNAa9PsEwj1bewKD/m0D79zwcU6qbIhdQj8FzcB5Xt5d
GlIBoyCUPGolebOIzGvddrcCJpRFOFn6Jd9Sz87g/jPw5aU55INcw7W04uKjV4dWYfeQja3RjDj5
s26WXrbj6drPdMeQAPZeqoOXUmFp/Bnn37aT0nIjb8RwJ8zrz2yZQ388btMeAvAuBNJ9HuQVbK6P
rlgtdUcvg5IL4n22Opxz0ZmnkoNS1Mw6TFvvJMJp+qIQnUo7rZyEHwSXrRd3EheDjr+4jrmg4p0b
w3LJ4t1ra4qL8tWpmfrBdXpLJEo9Swz8zKbYK+S+A737OilCMrMoLK/InDkpta337Ed9AxiL4rgt
+HkuoZ7bGuTXX70tyRJBwfcEsAZAkeTR2HXqKXg8XIXglNgtNNs20GIVbR7ohobzXX5+BQ2qz6Id
PutDyMpQZcKSkU8ZJS9J8cNqQZkY6YhH9k8ujy2iLyB9kcRI+nVd4109znhs3dW8n/ktEwH6aI8c
6WCxIa0y1WX2FBqq7bbSsTwiWnhVpkSzDDNL9isvsVXNotcoQfEAt0YNXannXEcPeaJ9lH7I9CUq
joMbo9h7rjbxnZ0N+T96h3SFXGvrUDvolwtRfVMXOOWogGNluFIPZ0KX0lHwGQeUoUjgs2MZYBTo
nLn0CZqgoahcrkONLKE3uESDrrVqyyg0Wl3nir1WZ300B7Q5Oodrc12SP+v31J6g6dOoHtC9Mpdk
Zm0fe+SHuO3+1xsd/79NuuLWIAAOg0f5dTZCbLJh/bMNnxXes2FAImU50HFTnBS49GbgFolQ/Yke
nPX1yysDu0zqeiTDhP/dh8b419QyFv5ZRtpq5h58bcmkosvh2rUy08qIy0INED4zV8y7ocuoLTN7
UZ2FkKxAFZ45zJrUjZIsgvYwboEM6SaFkgA1dy1/OkyQSyaff7vMyWOIdVfMb7V9NFrv+LjegW+E
Cq9dNY/dK2MUXvR9jY+l1N/7svJCRQxDxXFm7e85RqNndakOocHHRA8wxILoSmxDVW5i1eauCmt7
G2iMA4qHEqOAEMKeoagEVMn7q4VZC0w/aVNB1GlAOY8VmPtjwEVIEc3RU3j5EYMKpDPlxAVo+dY5
VGmsLh61oi7zv/GgymfbbWc2bjwzRfSMvCwPl+t+a/UBpVKYNZoVgJntaM66ahGl/HT83epqkC6r
pQWT7l7bhPXtU5KANQ+Yc+O0xbkKz0r3Lw8wK8YCa8KhNVFpWMKP9/KR/pvLgiZK4dWT+A9uLm6S
GWf/8LvHx1yGiUkpdDbGJztnvs+1kX8a3zT7T66fr3JX7PcRhqYSXHhDBQA9v8cve0NGr8PILYl1
PbYoB/EdyKLmlPAmA56Tv/leycZBQj2GAbf2lTSCckfGASteSutW4XPReWWQelxYayIHCWjNK1XJ
8U/hBarVacXIJfdIPbm1AJRPXlof/3ypAvKUjIyfXCsHftm3TB5nBquuA+IzNQVPCmRqIYuDfRCF
QgX0dKjUnVoLsNIEZLo+1QFchPvq++ruIEQtQvC/StIv+Ygmvs/hZwHgXtt0hFEM/FOLNmdupBGx
DQYmDohKV3k787aKs0M3i4FzplQIQQ0qgYvAjnZQVKA5bMOEOcv3bfc9+YN6QvIqiiNVhD9xUxTy
nmSTohldCZJqIIvPARVW6oZDcbfbpX/6TkyXnZ2OtfEKr1p+I7BWydZa174NwgreuK3gIVgHj085
b6y8BuIjLZLKJl/35r/0XNKquullAsNANpL+FgTBlKbuw6+QXSofVWPj0DfGmajPHOHlFk775088
zlEatOZVbbZ1yF/JYiF4oUYn+hFUkwHzncrOzqmkdqX2ieVEhFOe5SsHHoBdUWSMcIjj66DIaDbp
2wHZXJgqM8Of/jLjYd6tTRg6OuOUtYrLScKou2/hFwiUuucW1rcDIfQkYeYnKrs5bx05NCD6/QX4
d/UXv93z0ljXLcdt9gFy83QrcOJLb4ioWAy2acntzgYQAQcWCLrA2Kd0JqEzzO5oSX0E8fxuER8F
rXytwv3qzxHwiuldu7UePf6HyXNzmDNXx477vJpfJl7OlRHdc1IwhDHC9P1kQ02fqO/pmSEigNQO
RR94sJ3SaxTY39650Kzm8M7JGmoXoJo/xMLfmLMe6vHwwW1m1qMjgN1PaFQ+AIMg+MJSFV6vIjM3
XgYV5iUYoluqBRjr2n4aIojRRUAma793HhHZoWCwdiJLMP0AJ5A7512XnRZOq3M6HrhT2UJarq4P
Cym9YDCMCSUoPgc7W8OpaJhP5KA23Sy+n3DkHU8pQfeHmpbjM1mtrC/Dh6lhlALDL/mmNIBrS+xP
F3MsQRedZJb3ZQCdbFh2yg1d0kBC6diVS/apyX0LIf2gGl0Fp4cxdlTTn+nElUx/xYeQxp23gAES
XWQUfD5DdL+81FFBos3gBy+AcOU+xdseQ5O0Xf92LDrnpHVbS7kFBB5P6ziWS9f+3cCUnaBzl8CW
jQ/D7Ez1FpsxwSD9rxfSbNCYUPZnttrbNeeRMMZmwTBBBs8Tcl5s8BWD+Zz/cVTc8Y0eZ1d/fhqG
CMazV6UkpxUQ/dI8QyYxYJlsHXR/VsOEb8i8VxQdB0swtZpb5cQQghn5LXacCxLiwJFbT6iREdgh
meM/HA/AOp83HaAL1Cvgu5G8YrDs5Q7mzPdB1V72Po9yCgtPppeIKqK1Vq4IGC1ywDPVf6ivpbVj
sCbxYygsHQUsTo25v0amNSZCabDvho9l6zHwxcPqrjJYWNS0CnO9By7m+fGJrTyS49401UBEqyDV
DlYmNuZj+qHUaEeSWVHmvNGalZYZeF3ob6fqF7hgS1JiRemHvLxDvOD/IwBurUMJ5ze7IHXNT2A6
e4oCjhsgdnMeTetka4/TeUshNJhKqNKRQLDN8qSlYJN0OGxm5aL6NM8QiefRrtVU0T6qx1l+xtR0
UztiBX7fumjYptogVmdghNyDeERc5m2nC/Sa8SG9HHXVTq3CsO21E/cFL1U09NfoxA+WfEHEnvd2
Z7WgvCl18G5QvW+6n+Vtrwm/DJETISsm47Hw5kuI9V5m+nli7ISPR+3CPpIYVJBRhFtisiF5HScg
M8BBXcCWVNVhoeSEXpU5Xg4Gb+tyqHgnU1sOTrHpu1aCeTfIHQUQVDpxHRvtqKGHeFBYrENaTjcx
ZFwrmkB8mQOuZ1fyZNnvTS4eCQ+eh/c+mH4vp/KsXcGEdWw3YL/clAWiSlvbfcKXq5tyaUeiUYHx
rJ7ELBNtKfTAHn/6FQoIlCD8vkozKCEVDRROIqx2O8tZg5luzoWiC8NJFTAH1vSdSn7XuWSTly2o
SKPMe9uqvM5GFExoUxJoNTQayV0xthET7nI/i2vsOFbK4Ac7L0VIyzjYUFzOqTNWt4TX6x7VMzAe
LdtpPbhPWhfCv4Sd2hJNS+C+PENOnul01N82YbbKYKw2OozYlYPKBzbGyHO5Jd2iODgwaUhj5nsE
Vxgi8pvxq2YTCB94rIHBBFk3SVmQtakvXTECjRZ3LCh8mZcfnhmloAaKplvikfiKBL2HO3YrstqU
O/ins9HpgWKWdJ3GXOHoDuxo3q1USgn5D5O2fv0SYoRSdXN3R94NJkNg0caI8ZJHN/YsOy9rgmI+
n0Z18C++SnC7H+ZP77MuuFC1Wjf+clW8kEsV9WAoYQvqUzr+6kzy9RQxaEq/ujTt2x1tXe3yjtn+
8sN0Uuji1oCLvZX8Cg9pGoBTwDyFZ5veUrTrpqmx/BiLupBKFfczyKc/MHo8K4iYxa1khu+wkAPz
szBFCHwd3ryg5RLwjA1dDuVnubFF2EosjQMVqeifV4H2GkCSt1lRnwyatuFnOVvBhAHJJrQIFdGy
b111pESo+ADn8xSZNqli1vcAVyZPHEu9DM1JBEJXUm9oainpoteKHsDpnzmaP2lRhXGCe+U5vTlF
mMlqywxhO+EZUDcRsAeJ7GXkvmleNEfJOXuicLEQ8SvydT7IRGCXH1qyNPobEbxsoKj1ov/eokDk
GRL3+Fx50upP4VhFIwfkKq25It27Q3fE3vZM7wC4jum8OUBffTu1ze/qJQX6elLVL0ZOm0AMRvFZ
e6ilcGSfaCm442D5bZXmZqcY9g5ZelAjIgDrQS9ilvFwLz+UoVWdW0xVlGXa3/KY3pTg6Nfnp6fm
NeGy7XnPTyOAP8jpDtzPxw4h/lNhMTo++XRqPMB+6sOldS0DYhdhFJQZwzlKb2fTHW26t5VQ7oss
Q4W8L2wHFKNrCF/dchFU7t9ZpQN+J0/D/AFgOCvwj08A//WoM3x7egIG3+GFoe2njqLRFwN9kSZ8
/pvViJ8u+AzcUopxRstT/kEQDHqUj0+ukmxMG9uRiM/JKvToHOyUWt5bAutUnYKFak+6LQxChD0a
Ero0fWwhWqtoh5drJeb4BTkQYDVLAqVVqLmFvqOViqjBmtgEGseM/5uD25zpuTYGrP3zWKT5FKTU
85fd9Zt623gnxL6915YLfETZiZk6oNjSu9mnT8p1m674y/dH9Qd2xA78KyAq1ENKxXLyY3WfiDKO
FicvU6uljeT8ixV5AjxnxWKHoeWdlSSfRKWi0zSor2nxKaWOhSGe9VKjsX8WA3oqDPibMWm5jbxW
1asrfVt5UY6cBlzPG9tw8mzrBBdGKAVisCxsbmRiZ7dz8o9gdDCIim/saA/SYkcr9PUxFSi9lEhb
tttB8AGvypPPwMsA4Y3rPMEKwHEPjC5WsOvRzoLMnlkC929Hbid9+W12e/TDyvuEIQIWL++sHG6t
HHlFPHjy+JpMvMsRxg64NjztXXuTACyur31ePLEkQnYX/m0ltyOvDz7GAgCCzQB4QBqobPUBKY+V
IiZdA4yku1ViwZv4yoN7cXdmxR3sCXaM2+6HYHUB8aSJg+VrDJDOZHHaCQwEACNWBNAQUNAghprS
B21+ZLqKUFCisBf8pKmBEs0Z7dF6mhzEr+vizN4uFR7xp6mOeyHSbRjssn44qyEXkRyt5rCa1D99
SRVfCBWKagews1OCFopB/va43dDpcEO+V+wnboOPwC9Ut5clwpiw7SWnFc41FKMY3grXbxoUMPGC
tZ21JLEViOXkCWYCpnru4IVwyf2xLGfWT5WWMgZ1hlkpdbr0qsJpfSJHNxqQ2+HFvSH0P06kuFKt
4zLX+J9hTKISd5J9vceV6jwjyt6wb+HCC+vnAAqLWqcI6u+R7SrNqOxrqD+QnCU0EwVNskJiQiD6
rOy8DLIGPJNuJwejAbPFA4oFkLzvNwXHD03QoQrbGR1DN2jlEQUA4dz3abrzl3NJpYH+tllWqdnm
29soCSEcsmwvS6XEeYi4HKiG3TD9aMoLu4naUwhLRuhpT7kD7dofhpEBxMyJ4BEcpXSSS2Q95NkI
sTuEN+1gHzN/VA3nhcsnC8ISbmC7pQ6iF2UuwroxjH+VQW2d84W1MuUlU7wreQTYZyt2ykR6pBN2
uTvy12Azst4V9/xh+u1xJanwQJvVf+msHxvq07wPwHOR5G8KabfbZHzLJPJ2QGx+fShZcPvYnbVt
t660pm7R9yxpwiW0tp++lC+iMOi7mW4BRbJL15FZYNMRn02UxXgT59FU2c0gZz2VGvPQqibix77Q
fdE8xunYmQJ00sw8+pGPeEmu0o+yYjgdeUWS2zeA/qFfT56PW2RKm2/5vKMoOlf8Wyzozb6sosiV
ZWetadfdTffLmy2+6oi7XuWjjsw2ByFJgQ1o1U4WzxuEADg0jakhi4uOLNumpwMF25JwKhM7azEB
AvQnlOg0iHmG+dfLAGF6QIzsM5wefltvrxIK+spikjc3Og6EcYCdtnGDqJ3CKH7lIYjyYLu+rZrO
/2dI24UP0hJ0FYhIxV9ZBXsclX/WAY0AA4dnC+XUeZg9c8vePREtGuzLV2TJt0DL316N8ukFTMBz
UIiw3zyIv8/WZUVVmEMVPeJhUIRqY6i5599sylpHgTU3GVykeC3VxqbnE682Fki3tiupaxV6Nw1s
bJk6PwY3AlJmmeAMIV08Wm/aKsmJT7rVZu+R4PGbvOQq73yp32CxUnhhjUqlEXvVgsBHc3rZ5N82
OsWDFZcvR7KeC1broHXTQUJDyLQpxMNA1ziRxu+u7lqco8mwFdmLRHfphkrM1iMEs3w7Afh3y34S
OvCNk6aBWI8iCV08kgOZmYneWOl50iSvQdNXIktCD36B2TeBdJzF2vbvGOdCkhALJkcT27gCyr7/
qf/HLh0jps0IDKCKPNZKiYua1jAQJYiaQbFfaOQF3fYk+1zldBJkKLrve7c3YmTqVFyBJmDWFRVg
S9PipoqkjC7pe3C1WJnRUAfHtXb6YbL+nyK+JIEGzsiu3G2/VWck0rh6CvEBPy2U2mp6KqSYBhTC
bLH3zzspfu3r3XFf9ZRhip9warLEMmPAnxy8U6sa8LUlMpQcrhwhoCX5XeSbKwr2ee0U0Pccc/tg
U150DdBSORvVU18ChGcddsDBIv24spf0mPcnHAh4blwKRQeqlBeLqr9eD3sr5xdh9IrcXkWl3kFU
YiYgJ3ltLqYiCUKFZA4zjWeAFiuBkokYUAr9ZahmIODFTMoTkneRjoFA8EMCo9pJLZftu+je3Lyp
8kaaoYhCjk7xmdPnGTM8k/SvsccjkBtDhJeiNezLvZaoaqv6TwI3XULqXE220G9S2vjsonTotMkb
TnBfBzIVlpHxZCJw+WvdEsBUs+QubxE7BakyOGyguTTkqftcOrtGTl9i2eTM1VoxQaOOzzekKVkQ
pFGIh0exmwxVK2OTei8Y174hYixXaRbffGYZ0oFxgsIiQvNhSXj8Zy5jpzU5NSYg1+zNhgnQIln6
jq4WWVD6C5hulRNpGJgSC0gsQ9UF0g0ikyHmRK8RzH5xBlqFU4a7ZZGvAySMZD4gcE1BwBgaAZkV
JcD3XDO3vbl5RaOgi0U3C3n/PXkynq8g1WNiKlDwkR1SDXOpT8rZDxXdeOFNIw3KffzMcdIC4l+2
K8J9iiGACw/OV3/DEm6i+W7pGMInND7XUsxOhPVIuwp27EU6gk4ZZP7DPMhYIUr6ME+a5QBSWJbx
ijQDRXviJ8i08ybPTDBNpSLC0/AZzpDNkwBet6WkKdqZmd2TCemQlixXqY5bhV9h808MWOLVk/Lj
D/EO6W5pVSyxguJtZ7PZYdpjxqlZ7nYeO5GPIh98WiDbFuDY+6JrnYQmVBOvHJWZAGBZvxW5xQGo
YPpRp9IaSSu7Av2GruCnlMRO5f/7XazudtFmQ+zH+aTXCMTkkXb2bU0KZRNEab6sKFr/CY9MUNaT
jYSTFKEE1ZHqFEy+gdUxtAwDiofmg+gbvf037XkMAUzGFDh3gJ7XkYcLl6a6ToBM81K15DpTKjzj
nzWq6VUycCMM06kKdQpZKYHmMNhP5GGVBrxo8/KvFoAnQh6IpuUaOV1k1ILwGBGYzJZ2Eyzn6/Cv
TfcrY8wPTszegfh/PkPsXI9ztERg0NpYsFnfkZvDYSB7HcvQq1Zke6U7vWBCHDfA3ZzDLcR5eBdH
ANpgwtEaGMLe45v1C59tVTMJW04H/E0MRiaW1laNW0VuwjX2F8NJow2ACNzkW1W6Jwu4WCIHQ133
ucP6f0xa3txW67qpU+f4Sbwgo9NmHnfZw4DiqKcbi9JTjjNuErrXsVTBmbpfrFiDrT93KEnyPYbU
4Ljpha1/K1sLTjDtu04FG7+3w1CRMYnCp9ycE1kP2WP9Yj73r723XwLnuTsplS8ZfdmTprATRtsJ
6Ohd1R+XVntHQ0o8Qyqb+VQI/1pdEPoMuFtvRsQ8Mk6ai5epU02xDfO9cAyA+ZxX9xIMnd+LpJ7K
AWkgGgdp0aYkc7u+EPSB2PiLgb5Ey9jAc2q2N61l5fCpOlzh2zCjjjR0ho3zNMGcxmk4WxT3VbYZ
76diquNFxgMgqErdRvmE4sf6roJZiSriexsT0AP8XV83mVc3VqP4L1c38HxijsAiVc2HJxL3rvFI
eNVCsbwPuZTLZk1Q+JRK4crMEG0zgIWaTRma/aTXqCOQY6scCMHeFMzvFx1mv9ftmLQXwtE+aA6e
9DnhZ/9w+SWRKcNifxwWCFHDS0iomSQnH0Nqk4IH+njY3tVHI9pye+Z3uvSUWjFPVBy2FCtw+/Lw
7h6wBjI3E8aYGFph/V+VpG5udV2XyaTQthLLP6W6/Qia2/w3VbHgdB2sUxODd7h92/6VfJ2QaRLS
WNRAOst+GAuPo5jUi63CrY70crz0s/QGPhuYwoaxL/8ocs4C46+hijHBQuzAQKH8pQJDmH+TTIkf
JEklhZRr9EqYLexvl1Mg9d48kqv/Hez/tZEePAPDfd79sWMwRm1BFdcOTXglpwkSv538z7mvPCve
JcankjnqjB9Gc9ng0skso1WcWmU6RjFUjjonzfQuauJCZY/+wJTgfqA1ngwe2Ic4zmgpBnPSBjxX
Ouv2zAejXi4g/Hpya1A8AKBTIqKE1+KUvMrwa63gmMVCwf9p/jrjoAiOwHhjeelSFafDqI+OTTyP
U9bw+S72ID6XSI9f/a8nVO9uZ1xsrP3X7qZeIRjLlDvCpY6kUToXq4f2963ZCZl7qvCrbzJRzb/n
CHAUyTcA9Y+TI0SJkSJRsUTHgj+W85VYGO58ZaYox4wJFFERcJ7S49/XqDTRLU9CaV6/L9Yb5WRm
KfTI40Qp7eEyUTGNpe3VoDOaOcrd0i3565NAVXxQQ5PIh9hAraM9iuPlfM6Dk0kfgeAnPMcCMEe6
pjCpBCHwhqYvk3BAMokr42JLFRHshbJRa91OpnkaGUbyfaA3QLOYD+lhirdObuGtQqa3r68OU/oN
QUqnmBe7zz5NbrdjnVEw+mD+gAWldPqS+zDOf3kNHmJEqR+1Xba/Mlpo35Cp+NviIaqTrsOAotxn
xXGmq2KvxavUXfyFudHdFd+t27afJ9L0zFy2M5V+n1VxTTsdv5f18olN2RqetuIJ+O6SOAPPJr/p
GVSIykqQyFUf3F4N4MAg5DDzEs95U2n35+ZU7CHWGGrqnJxmpg4k9jXeROAPvpb/p7gUUS0B8lXN
zaevnRZFxbx2+5B2WlKuCnP1qQgraJ1wiF6Oj212NvKLShsuFrMPwBxIPi3J4JfUow8VhifQzQs+
aUqvjt9XwAqpS+dpbbjYCAYoucdvvEYdjpw9s9qGT4CPYjcRgUOhvxylD74iuyTrEp6m6mOrMw/N
QmOTxRWWaOsIkXanBB+AKEiOBDkPCanN1G6FglmqbH24MBY14DWOgPk3lfzp8RsU2X0wxDJZ5rsd
9v/eetWNjLmCxsyeCSgBL0/sZ9/078yaLxZfdwnMkHCQNYuuFgySXTfqodbPwJC4Gko12YX5MiIv
5hxL0aoFu7mkgDSFLL+4QGKu/HnnY1OjODeGsHI1kD+2Zd8YjeivB5VEh7C7by5dZGfkf+aJpaQZ
MtDMS8GGCwn6uTua+PfIbGU0+V9soXCvapY/k2ifj+8eBKf9KTQHqI7Q0U//+hPA4GlKD1L6GWFy
r2lbcQ4uDuZBba3/hXkctp3/SWJnSy+dUYED44mTslp80O2kA3KUlf+tlCxd5BC/yr/0ragxVd+J
KeM9apsBU/D2FlHaBoit8ZJyZGOShUIym3J2XZ6Oi5Z/rywOlHXGSzFIpQyENJilVKX/ymravzsz
FIe/FctZQ4CBj5f4VHR60nSJGDCJp9DSVUMo5toR/mVDuqIEzVdR17cmCmsc1ldMi+LaRvIaYTNW
pmk5zSVCYCiPKCK7C6Fi+nkGhSVBD2kn0tZmxkuuJGtU2rUc/4sCj286THLMDHi+MLOnom77jg3H
9b9Bk2b2fHLCu3OaYxUkokyCMSubusTTj/XfVqvDNYVOVJLRlQpNEy0Ae/OmNhHfsujyKWvYcM/U
NX2MSc8SNQcAEcB1lIl24WmokXGdnTLA7Su8tCpbhJZmGrB5S8gpfrqC3/p9EMxjfCqS+o5tnu9g
FzqzSbK1o70sQxZDjWqIjrRLpjl1+fkub1+ks36ausZhF8xEge7mJ69iY26Dsxbs3HGefEiqfv9a
FQ+kN1W+Pdc6Aa3hVFjFh0JlCsPSfgnc7WPGEgC1UG8yky3a8ee2sAhluMnW6Ci5/zlI/86FToG/
joqizaeUnBpqlFYjOSVc0VZ3a+muIhCfPCXElUQIosmNHGkOj2lEhox0T9YmqBlbNVvCeXMQJimr
3QBiyt+fT8EuVZZnL2i7qbQE6qSIIfbJD6vol1uKhE9qkfPcSEKzulqhHZ9Q8ruzAknl/693AEdU
hx7FW25RXJizQdiXC3oa405KHO+QCkNxa4YqMTPmO1amz21/VxhUiaOSGPy0l8EWz5wzA4dg6RfT
nUbKJF8x5NLtLEQ458nWxh5MfwRB1nN4ASV5JBOBG8nps9iTzOGlzQ3SWtGuf+EbVdZl+7zKP+pm
9WLPNG1MfKwIdJAzYqpifjyU4TIvxi5zq2SQTJMdJjfHk9g6FhGSfBU5UzKy/rH1sljjY+aaibbI
jzQbPyZnuqa2dH2QXBQxoqS0Bx3md9JWontrnM/rz4rjA80lesd3Kg7GgTNSTxts+H6Yx6I/+pjm
7JkM5OMfpo/KArqgQbaqeivuYv+g/QACLTQWEtNFov33GjXv33l7RDHWvEj70Fb7RjAJxVcQvInu
r67aTx0bZWlnhlg5WOVxRdkyEsb5T7jiKtVj7DFrOfUYkhEoR5w/0Ji9nxBCqDFVAvVHmgrayqlq
Pb9eotH75mMH3/LGxasf2WzhpVxWnJ5HKNun9JWXzjC5/fMe28UHqglSkINkg4zD1GEpJGjwiw1l
3TRLd0MABIqAK64//K/UKBuaaut+LmVM9lRS/x9aI0IJX2h+i2zWSMbtLOMjlRrPzipUx2BXiBf0
srt7IZA0j+iax7Qu9g5I0VxMDsTcoqZGirTEHXQeWpol2peMihVCxckJOSEAIUEwhqk9P3tIDt5c
sBwqkTfEk27iWlnqhrN+oRil9P6vrq5JiC9WcfrEnxX044NOcohhz7DT7uyp0IoFxuB2agQmJ91g
aGdd3hZWql/h80VP4/U9+S5qTWwQDf4Zjbj1pd6M3gzPXjCL9WZU9EgFALrst7ddz6yDkoB43JI1
jXepGPs2RVZOATqEMKnCDaKlv62KHgmknQ0ZVjA8dytJZv5Mg9i7MVv/jlgMyCaHkuLVfhhJqNU6
MHSIeEqQrsovVQYDENETqF3PD5CzcpIfhBwXAI8p96oHxprs67WCoWF5AEaTaZZfYf/1yvB9vVTp
BHlLq0pj6dh9dz0yq1Zwk/RZXOPvxSP7kx0HaQq1kV9zF5H1Z/xvRXrxr4a89Dt80wC4m/h8fIXc
2mXJTLpqMHDF1YrkXRfosauyHFZPzKc6wmD6gNhLZwFUQY9pfwQhpkbH8SwEM3exRegmRAV6EejK
LL/aVZPV+aNy0u9gB5s1KiiAHD/GPGPb64dbVePE9kL2a7qCuwnwyuiRoFnb51Siuzc8hyPsz6OX
H/krY+RcEeWt92c/CxlN3I2na0I0dau2cB9dA8IRJp1WcXPijee8XBxzme1O0fgf0DJoycRIj/6D
oNW7uTcvz2mBXA/cR3UOKgF29weld8v/Qi2fhqKJOszyHSq09PBfCM1W60D4CqZ2QBWMUvOPOvma
A+vPgwlcyjleg1MfDs6LLyQukqJM3Pqh5UiZR7LbdWPWM14tei1F6AhP5gRqsyIUNgiKtZ4Bwk6C
6h/VLcSnpPHT12qUyrOAF3QAuTpQIoMLStiCypMhE1+k8hF2jdlV4khROzzR/yaQYCjQ1yqQSZjW
mlM5vLOTU55vsdWoiePIuAvdm8bHlgCbyMea9neC1Rni+cfgFM8QGVhske0N/sGdlnexHuxwuRpm
LKkLT3y7qwp/pG5QETNANdw7cO62RzuRZZ1CukC3+EBemCJzRdpgKEzczSJGdYnqn4ZxlLyIQC7I
ZHhx16/A4D8r8kcyW+b06gZzEFilv7mU/Keci8rBGalhqWxgJesPYcXSlAQws2lDOAaSL1YDgm64
p90fYvNIMrTTxjKutIV0mGaZJZmQM6wVIl6GaHJQXsT+2HRc7saaLOdxfMwr8vC4ZGNPvfTDMORk
/hJ60nkTLwWe1siK9zQ4wJnT0ZtaqcqFbUuOJBPVTpcx8n/gj6ljvGiLzGb7Bbha02OYHWqu2VZQ
ETXnAzkQxHs8Dvy1UMNS4LVpE8UH7rOjr2wOoPj0WfoKUS3me0VZvAHBHmOcJLtcoDDGzY9oXUCt
iPnZnRoXj/8GzvR8Z16AO2QR1zV3C94tOLb8tWanA210Q4ANr3Ymm6PmazOOmiRAICifU6i2BIIz
ajRM3MSUp3m+CUSeeFYp2ThMgGWBCNI6z/XzlMaoBZtTDd1RsoZb3Q/bVs2LkY7dGWE4YbjUNqp9
Kz9NVuF+xoKR53T/dVMQrkWSBGbdmiRARPOCYqM5hHSoUpLRGmlWIwhlvVVaKqc3SS2XdCIzKxCD
v44D0G6pXg5vBC27xUhs3Lqk8duZfY/CB+/40wo4B09Tbf+KhuzK6prdIj0sCUwVv6Wv74NKuncr
ZLSXAjkxrR19Arkm4QvzN8g9UlNZjonyQnDR62m7vDrh3VsizGlxZREMTuhwj5P2qZ22Sbas5H8k
BMaRrMcL5Zxg2qeX+Tr6Cst8bxuG24h+sYkNqciJAbaF0TtcUQsUbE+F3l/qATFlQBEha/Apf6Wi
LfCyHcbkAdKheJRQm0hClTFi5gMDVoaYTWkEeh7LlBFx4O0lN5d2caJDjVOObypD1NsZy2J0jOr8
5OeCGHcnK9S5OwjDIZS7H2wgnTVePiBsAeeXlTkTc2jcc9PYpcwQ739HJHVJ04hAxsMG4vt8zDue
shze0rON6MPKdDyr6gKNRfxnIATUPFE1uzUUYMEg3h6oWlJXMA1Pztqb3R8YzSV6QKFQWI0U3Sfs
Y2KoEhZGOfd/qkt04Hfv39tiImZKpyZyjlCACdfNJxOVg7MUShLSJ7pOldvFzXmHVn3U8ynwtXdb
ulTxWAL+tm203oZcp1kUoyG5DaF3zeL3RNKVccp16ycx8tcEDqamW9JaJUqZNlB9aiwqdz1N3nBJ
xRjKZH2CjWRiS0EWuG2TzHtz1wLHZTtAt+At7RVNBh+YwIP0pzS5IZXyb3rpL/qh232WBu3395Bh
C886Av9/qhvOMbyeYrgp9DIDPwxrH5TakbwlvHlMppUc2iqSzBHC+2nB6ygDodzcaA2zmc/3UU54
CZB44KWSqJN8Ze6Op/oULxzlQ9hFUfIHp88YUR10KE6U7XUTsTCCCWrj88v+bDxDIqf2Ao6tdL9l
pzEVXdSeRBVzD2dZLRIGv0Daut8AG53VW8VZ5aEU+Y/aFAPDWJ7NO63Erg4SP9wPP+CjYDgzhhdj
VXQ5ufPAHpIhT+eFqCh2mxTEu/F4HEF5/fQ1R6rqOaZa4R4I85xVJ2mBm/JCKZYT+1JfnI7jIYX8
hXmGRQ9vZHmBznKuDC2pBMHVwHWXbnPLp8m3z6fwTv/kFpqL3kBwj9q9bDW2jWM+VwzgJFQmuJOH
gbIjXLlv0AFqagELTVXI7CdjMrUWgo+fsbLULy3C3NVXA8qkkCIjxztZ8lgXaraCy/B2/jjfVCJ7
OJHzP86ygDdYIZQrJ4wpPOrHdZmPxyS5GdsWzNDlPHHtl1jTBDTqz9aHuUK88c3SxK+iIjphtquU
PpA5uhNFHQSM1Tj6hIzeFus3aIQRsTJ/EzjOak8I7UhjBITtTPfyFN7vAhu5ebHcg0UJ/Qb8sNPI
BIeUexdgW0+jUMLVaO/l01iZ4wzuxzoshy6WfwcVMdbvvkhI3WG4hYNX467MuXLySHqo8zYpGhru
PCWGD4BiKo37V+7afwR8V9C3r5nRuihapJiB8TzqMW+LhmSEVnPRpVgPPmDcban3UaoRQivcDTAs
ecr1695SEUnKBtAhuXMnvi3md8sIR0qg77+4cCXpKiHtBQwR8qjC4Doai9Vg8O+fPjim2jfyG+Pf
xk2j4YwweX+PAem0HaqYo3xcUSHcOP0ivN9Jg1vrN2LdOrQa+Jan+G43OQfR9XB5fnv1M+D3daL8
EIxZY4EejNpq3ONpMQdw4NxAr8huhWpLKdIBNTPYnnCxgYW4tOFtQD6nfOhYw3h24xpd2+lon3vI
CedHRnrv7qHvYUAsiK3aPzUtwYC4TyhGjeT7n3RKzKproALfMlNTBjuiBqD14w9odD6Dvl7y61QW
vAh2GJBinTH9+heqsFFFmdLMqhnYngyCL0ypVnSPo/r13cI7x5USnzDFYoKk+0jVNWiv99+v2H5f
Tw51p0Uy4epokeXhjD0GpPPK+Nwr1vdhBNvrRnzGrPXcdarggpvLJhW0ZduaDGMIDIPpwon3/ItC
w0YgffUC+H6IosRMxiWFIBagUb0ewc5eJPP9czi16eLywFpwRN2Nq75387BE5wwF8g11byVnbFVN
hSLo/QxjWHnwBnZ17ltW/KUy/eRpZ8KT7P6qeCrep6xfLZFIbhL10Fc0uJpceY2taR7cH1ChLNFP
NLnuWaCxlKtGEqgwDQg708b/OcanO9AscaGAOwziMo4HrQsaqlD+tqo6vfedSXoCxMS8eTbPDf/m
wEcvGe4+n3ejMYRUR3Fxxx1OndPIV8oqRTXN4moxOB3Jq8pMmxVdlYjSal1uCawNGIbm0auxuhaN
ydAGYzrWUR6sPgT2vdh2l806qCF9Z6it8lk6aFxMGSRwa/uonfMSdlpGaPQsgGAZwgsY9u952rQl
SmI4q5FhbV/G4DIszj9zB9Be42mQAPwrQDF8gZcsiCf8XiVkZZmU+fXwd6b0NKBlfVKRUYmR73Nx
Yt8Y4F8Aia4NZFlK7Ykg2GBT4layUs+bdMu2Xh0ILzu++JxKzh0eZK7cynEKFlShDqsJAnenvpb9
Q452ZuedIRkbuIRPRL4qpVML7HOZkZJXGl9jloqt7VbMh8CW4qzG0teZV+DbCjNZ5duPQDNP982k
xPwa1Pdh7mW++qDOp83bO2HYmHRoE0huDl1Ym1wjF3ejQ4i+CmZJ4aVGpWZsuxZPXak+AqoZk3N6
vM+0q4JKC1RagVZT8+9VGdFOcgzk91N3wDpr9dpjLPkGq5xsYLdj4Up3np5IDrUAlZXk4P4kij25
KQm3BaZoN94NFfD5N335TWhgBx57kB5/IKQeTXBaRed9/f37TtrDECCrumGpruEkumRK79XqMcwl
2Pqvm4jLxUssSApiU2VfG5g8Uuf5rz3UYUMF6J3gkJfkdm0r7hXU2xdFFzlJFRsKQO1r05HrQn2E
1UD5p/jrw/epOd7SbAYw2oE+wEdIq9XKfqpbOU97JgNksyw9V8/pEOc2FXAARQ+jAaHjSIPMb+mr
1hkVsxU/7NDJafxqQypsBfjI6aMu6B71zdAIezVqtDrwgiN7g2yveyUg3LJ0tqNvHGnqlm236FI3
fEkQZ6VYZOgGiqRbQuvqJbTLUlFY7MZFdMKFmZ8Shug7E9daQSnqaVTluiQGrXfUWdKmyZ1C5vGw
zbKy9pt3V4qbyOMgZp6QHbSB4tvaBObtRX+zDNzlw93qbAfTuXoaC520qUh+m8XOXQYY9ygaCh7s
nr1Kd8/C3Fb/WSG55zHctT7AbOd1X9k6pZ/ALzDYWq1CkppPyrf2g70GZNAbHP+K4G8q3TcGt9XG
0Iz9rbpqa11tLOYTyonRoQfIf0a0fhyv+WtnZ4HrW7MjR/M5oxXCgm0b6DIxSpHCf63hc3M8WYZW
zHIqsod4Ll2SbwqDoH8s0upQvSyuA/Bg1MT9N+Z/BBgTrBVikk490FJC0B3NzY2zMaH5iI9dIWwY
dFzoa070Fmb6WxleS/rj9Grzo7ohHQMG+qRtxXwOX0aE+BdAN62WVxobcGRf3dBROmWS5sJt2jP2
mNW4I3zhyt+T/Od3ZSOJKEKBQiU6vN3P3lm6LgeIg2TLK80+fEQJDW0vFyNVc4P4qyooGMtBLPbx
fb5LXeB/yxcSlsf+qVYw5OvHl90W3K6teiIf3EyD7uFBiHIhh+ECeRlo77yT1dtGLFc4jn1v46uj
MbOS9rsEsQl96K6c3TFBXopAj1qF7XJx5lONXJN+nWMn9a1gcnQtVy1575tkoNvC0H8Z7D6FETBk
biafc86RbJRbxH2cH+CYzdkM8WAvevRhf8pEuRS86aK+OOG2V1bSu4NjUuYlkafc1F6jYg9nWman
r9lWP1K2QDy+iYtpv7KvlkX6RpLOy1z9HZ5ViARIEtsjplDcDgUFkFuMGkFR34ir2dazM6uZanmJ
C+FAvuXs1ez3WU6pow3xzeQyg09fS7Y5hOd8yRLPirbe1s1AlpIhZtDVZ/CqmpKButi8aZTQaGfS
/wc3nrbu8mZPZSTsx9MV6nSY7org5SvkzE8iRCu2xZ99zWvh3/IHQhDSGp8Nd2ZeJi1xEIHqMfs8
i7j/bdNIH8kMaIhFkpaKhftHJCCHIp+MsfaAFaa0Fq0l26n2mr7qSimcNY/Z8fbPUICgbe0mE4bl
3VTi3VBdgZvWq4LCiEI/ZkWlrW2eZiBDjDjPx8escyUwESStf2O2TXPpIbIZrBlvfnTYhozHAqtP
CBrPq4SzcuMQYIlt2mbvPJNlt7mpteaHwtCTRDrHQOpXtkUTP8XtQR3zFae8hDEiBUin+S96JN2h
N6dEnKZdR4/p0UP6wZ6NiyCPS6G7M0IOSDn3keG8QTVTm8TiKKwcsojMOeTBr8RgKWvZtbtt6g8d
6625KEkWcCvPN8RjtmUVLLIrBIEwHYaPCfaPR8F4EtAge/udr7lMhh47tXFx4XrU+e+hwntvSHAc
i+5XLeYK1IcYW2BXOtQ6KKUXgbHz8Av1EQjYoNFksHPD4B0XiovC/7jd51AcUccjQIu6wUfRs2mx
QRkDxexCx2kTnvPW1yqu7jCUet+6wUJEiyfeWchMimwlnIaPU01NeaNW10VrX8e63Lv/BCx5m0Hg
Z38AK+JObgwPSN+rteo1ijL9ZioFVUv2hSmippfqZ6C+ddFZ5blZMn0XhtIQMwxMyr3Z1zywGS9b
0ybbkuhC/7C4InsfrUr0glQ2vLzLf/Qe8ZC4AylGehNZSFyEyQLsnLvEm9FDnPe/J3s5hsn+icn2
RcQvafOsCtCb6rwHT/nIx77vpAsm54CG41ZADuYEbZNoR1i/vvzs+0qMKj0FY08z4uPbb7TmLYHR
auojlKZOXjwUed7jKy0D42NCnNGY7J0R4AB+b0XbuLKZFJ8eiDASuk15ec0NbpL3lAS0LSYGvOVp
xWvx6xshOeqq/8w4e2qdnscBxO38Svz8sHhVKcpZw1n/tp3J99VtVFBWyk+FvmdzLzL3BQTJ3nQ+
ESY9xba9zGqlklR1rLBFllT1V3CgdwlwUls/d0sEencpk4+HiRN/gcuDDwhKqlinjcdhD4cFbkEC
mUe6kwvK1g1XEotjyRU940rL09QPodl6ZHYzhCS9KtwFZ0IDc5BiXzUYHQP8v5F+fhUPWWY2xlIA
itSArc/wWfgU1tzq7Rhv/7oDWr27LStFJ2h0aIo+7fly787PITw54zuUstUKXuLgDNWglNHw+2VY
38iBnrbx5YiZvPBAErh6I7fG565d1NLAeFeX2EZ7PN90QXx+SPGs11rJaYYhxo+pzpVw1yppbYz2
t/3V2M50jJE2GV+jOnE6Hm4dIlIC4Ciq4p+dHP4LI5ufgB0pNjS8QyB7jgLo/f5rV11lPztQdWfk
Ol3oMubqtDZp2k7XIjE6ayfWVSGssB5CMrd6msqef6dVvDgnwSyvFmBBFXfZVCcPBO9mKDXEM5rN
eAm+D3CybOXgc+q+Hrvs1FAQbsf3CcNqATPdMUWYrAGxyLQnd6fRfE0slkc2I6DNXPZ512zf6nh5
pSGsxGQ67ILZw58zJdzbZdDL1lzxsdE0ZiXqzupZYxksdAJDGfmYIv2jH3Zke29ytaubYbWL667h
Mnrgg0Uvqbyim6Dtpg4Lg1gn3RoKlKJ0lewyUyqAhs36Ru43DpX0ezYN/p53vomoHSafjngG6Ime
PKAcnKU+ByFJKTEaUOB3nTLEX0PAYqDTLTLIGke7qPYuSM39v2Fp2EokTOgu6K3NDUx/ps25ycxA
vrLwf/ymi0kuAF0xAkuQ6lnqytNhaktRGZlgvi9rUvGUwzbKRW8lYtLOrU3MOHut3fvcvvPJeWjI
mMhR1pei39KsWLs1nXcAKfQGPUGP4pvc60M7DzacM+tBopzqT6g7SnTX35OfG07gos0WkI3ISDSd
cDI/cLlo7DBoa/1UAoSzDGTLULFhK4zLWCW1dQ8eyuUNGKEcUBFtrJHdwS+8OZwDtaRZZ9ISrLSJ
GUwm57cw59QC8NhDNN40/2+122El05yEiHSor4fZQtG1Y3DgdgRbjhxwITPdV8iWfEQlYLWkJHP+
DXBMcLRGCY0TE28b2CS3vITf0N0UIA+X4BDu+QPA+e86O3LMV/ThAz5yco6irTe7RHoIEBHGNM9B
/irw7o7H8Dk+JtSHuLNUvTwCzaIpN4FcmKi+ZAbHpP7wJu6dKy5wywCp+3/2U7NmP1HCnNfkFPKD
V2Rrub6tbkMA9A7ggWItdDoUrZ6lF8kYDm61c5yowD8IuO4stXwc0RX/yOQjX4s4VLPuEY4aNhkK
XWY/RrQycpql3GaMHBkkOK62Y7Gy2pToNYLHABS6jAmh1SZCk1YsZmpWYpEtaYWTZtOQQxDnz9Nc
SfTXMYOZ5wjpWcmMWYlG2b12qB3TuKVTEFE+VyzaRYhJTq+Mc2YggWJA+nYbJzHzzOh/+JuE1tbF
I89Ymd6df6sCv5AHiQtKLOUabfys0WlDqhTfWkTqDCQBmfGZlb6IgmNT0x7G44aReYKQf4C9D1f3
OlcUguq7IYHTI7Hs3h3zg/D3xQ/gop2mynyRNHpkpHwMHEFCoh415Yjk72wErPCZyQmbUTfZ4Vpp
1BlXSUf+2WzryvnsL3Mqa6KqjD/rJ5XMyhKq8cTgnQ6k5JoJh3EtYQFKLAnXwn5KFIuAP9hInWaS
hXC2Y+Z6M0dfpwgVfwGQVRuG3MOItmu89q6KDIK2Mo/9dxD2aNgbjqLj5303c7eIV6zZbEjeH3y/
VazipZqg47Sd0KLEmTargATZU3du+buw9YESaHA5IcEZ8L+6DhGXrLy213kyXoqiHzHZkqgBkz92
UEyn2krUgBbHCGTrtECGXbTLnE6WNQ7lBtyUZ9qeEk2XZNgPSTWCTiQxfDtMaCrMaAhX/d5CDrVj
X6UPriBBx0wQ746N9+kz7ILkxPXKA43HmAf5J+wukDaYNvgCqDnBHFiOsRm5pIBbri5PKsAqwow8
2grhuezMnbw7NoXSwRMCL3JXI3J0ws4JFkLhsm30Wdj9I4ir+nB0AU6flRHWQEawmD+Om6LkwY+9
gNK3+oaOJoG48lSnVXb3mk3LMDpBRycoGL8TT++5DdquXhnK0je0xTSfGM6LiYo7SLtbgJlpv0yZ
039QvhdSjJvr1eHFBCNGYk8zIWM6b0XGlHexYmlO+pYMz15sd+LiFGvwoGKGz0y1JlXBLRHwoq6w
MLOZ9DBohTDuc8TaNQf1nYGFiFrVQPC5v/a79niMc68HS/ut7MgWLSmRu/xOMWOHjcucELA85Emh
POfMTh1DUlYMI0Q4S8qXUwzNz4U5GWH3P8bC5t+vafmhslHdvC3oGVRuSwovbCXbYKE0eqYs3cOF
q9f0CR1o+OBMh+HS5NSwfyj0U71LOyj02MZUwL7Eh20F/bN7TEJ/yAPnOB0WB9PCOGgzKwOVNReE
mLnpjfu7jyol5OT6qgTQnRC/suYIYG7dOkAWpUbmtiAq/6Zu4Zay2Boqew92cfdAh9u8KRZ5njVR
EvV7Ka1q62Ek8Qxum6CViqIve2ja6dQaVh5GRYxoa1NEJZSdJ7o8YvlwkAjgAXbpFwhNdH4yERjt
mS9IFwBG+IuE1fbpOT9cF5n0kRkWLOgwaojYL1XQXcw8ti8iBa3UuyfvFdcuJa8Ad+VxuncGBUrB
g61gFMuFZvbxAA8f1TDKQKHSQuB/QwESjv4YAZdHtxyD+RUcxqH4jf1cOKFvqLuPEaQc/qvH1ZqV
TuoCATneZ9VJMJsBH3y4aqi3P99j3v7/fAVGr2jqZaS3LrMyeWNvHx9HgVbjxwfh/WMWx80IPWHd
9VV8G+y6zlUqjnxjEHBe+r5PhsYKt4Br8g+XpJeBR9ilyBNCnxhe520cC1GukxQ2EfpzjrR79T59
GQQG0JTDAG3WZTDqToTfGeScXy8ydsfqZ7N5NEyet0O8jfRlcRwfa+jtBoODuCGT6p0KvJWJLnpM
Pe4XFR7GLEKWX57SCykpZo8y9Wew8oScUCcD5JmP09HbXv57PhftcvJIOOJa992TSykm3xV04DdF
BXiqmQto0GCEm+FM3cy2Db3PsoFVFleatWHgBRZ75Rbgz2fK5yTI64G/p7HppmWsH44HnR62Z+r0
0sObb7Ao16HdmEVEeQ+ZdbVW83NDJcojZUt0yG+299KLFN2XBeUTrIDaKp9KUzF4YehV+yv+b15X
oWghVHVnHYTKIUrK8bPfzNLVTaCwVtR7NWROROdkzIj+dlyuuWNP4mjYlT3+v3UA9A5TvP5vH78y
YmXFHglPNRMVhHd3e66Szi+d5uNzOgUOXxAziipuRWE76gFwD9yvgSmi/pYvY1e03N7+14A59FjO
Ga5ZaF6aiubKYfGYrLtHdKqvhyjc7TWmWd6wuUrVoBig9yFRtvup0KAseAosRGHPT6qwdmEmAU0m
j1hFLiQbxS9aA00gaArHnOgiOzEKkUJrwZ/dn9jN8DzEUXVMhyEbA2QpsFpDMBdsKQxttPiGqyGV
Wbkr8oY7jx2Npv+2QNIGNNxhMHMagLcJKy9dUEwefG8yft+TFSRHJx5xhVmBgPennyGTYTQ9EII5
FtKjyuPFkh0lgnx8QZfV4RlSSY408ZeIOcfa8lRGoExE+4vboe+X5W9ydGc7u7ygYIHcbqoElvn8
GO1ByOiCSCFi7J4RyGBd4APIOieETceWeFIlxFZj5jcSPnHLLnElnZQg3pSkUUD2R6gSzY9XVZKJ
gqRMBD7NgJReP6dh6rLesSdVTWxISv5g8yLRV8Sq/FZZvftgdjrHlMyATFeDkb9D7YRR7RuU9HqY
VZftt/al//0Zg4/Pm6W+sDMUcVJot7+T7k/V9OknSatNgMpe0eQPAMkZselFJkJ3/F8YWvbCekB6
0flhSyNqHmE8QoUkjQYXQuGOuQusiRVE/FQzMStcpVNQ9dvSJvyt0KhwGMuTwByOP87eSgNLJdYm
ykOoFBGtHyCOSe6fOeCtnp29ENOA/oXd6qyaW/BD1mpTK2zvNBNC27kef2IOCHzveCHMy3M0wXI4
mFZ81DFQDxXXLzfwmuIHqPfB3IUkS3m8y3SXqd28bUtLQlGPhqLgw60wUSeAyGIwR+j9F6w0w8HG
WMcbtEHU5ELsb6U+yG3Ml090S5q4Bb/bG5gs+XLsW2+HFZ8gdZANc6J7xeIWlCn9hS3eJhm2z2XA
PkWTDVx/FIoDvXLsO8jLHkJDWdnX3NjDoTlLudN3iyifBYy3H7wxKN2tG2anXwpzqcUh2hNnj99u
aNt+oTfbtKw8qpRLFABRVHAEEWXNBqoHzTENn1CUNFAkntZLP0pLT4trKTKBCD9qpJE0zg7OWqVO
K6r2y6Lffk1kesA71jvSWqJtz+/Q1qJ5WLDR5ckYYRTxkEQ0vfL5VSdPwgl77j1Adp+hAU3iSGse
GdukA9Hyew814fOaUe4RqD997+vCYZ4xmWO9nKaUKzsWPCKzzA1iotjKpRcVejCao6/KOSnBq+9P
o+Q15/PY4IaaspOALf3HuY2hSW7KdIhj/fKiHtLcFG7O69njF2eiWFvdoGyWTNJymsqOWzXX63jG
pKCn2yqzCIZprHN/l40Jgm2CghvwZsvw7mFOsxZnk3WN24SpUuTdBetfGM/qEDmKB+4/6GIjRWjU
xVGCbhk+SJ+2cC5uxWZdlw1sHxShJ2dEzw0tIEc3zTtE5cKfBrzkpJOMjtIQTKB17BH2Dg1pkhgs
IcfKhqj4xAomJXnROxZ96WmmAoGyDM2ukLlwzqaiNhUBUCIoOJz7sCA+4Qm3Od+5tqn/puUnAnHp
mVtTIdeOoYktAHokAI7yz77nALcSuoCUKlP+L1YlW7NR4L3Vw2JMNuQQO1MF+bhVkF8I9Cjec2XQ
tNwEac/y5Hjiew0csKGhtg6GdHP3h2FqUltbwhwiAaZ2yz7KvA8s7PvXHxggZZ99IVVkGUF0lbcK
BeByqi5/7RqV+aNW5vjnZrJtvLKE3vYwvVWqPTbBGfKhxXCqZiwvjO1WanMsKlfTry+6ybhIXY3R
mq+FTh85/Cs8Wr9WeqRvQL+9DOivrhPhvUKEcwqzRcHX4ZyCWEl2LhiJykJk5COax8g6OBsglgen
cBDDA/6Ca/Qs2QlFqN+YD13P/ztoWslgbMwNh+jMkzIla4xcd0IsLhQfpUlJu0yyfDUrBYyGCnn8
tobKvcMi6vQK+CYIplFSZv9OhJmpi4mu3SY8Wj8KPdgNwZSpUWUei29G6mykGjQMIm4hmY5I1NWd
cYUA2AvJFtCWTi0cs7JYm0qQNaLoYtgG+ANsfYChDAEzwirnh6nD+MzvTMEQw2SCV5wNdoJTnlC8
yqpcJTjvB7N9Ik0wLmg8jlJsnbvphXArK40pEQEGZgo8FjiBQ5ZdoZMg+/wGtwemc51H3uBpSTwj
UAi+MkUCN7Nndao4reuCb/k2zoxzCE5A/RLCAUIm/POFgWRsZWCfxcc4a4ADk0KjlRIeonDieKrF
rU7q3Req3S6RuMsO7i0XHN0t/YLxeaGNZtvmTe9cNrVlEQXoEBWw+nIAvBTXwDiIRVxeWgA1WGSc
UhMxCxxj1dUzpQSmxUJf25fiRle+AeucP868dxIwfKcMAT3YQo3K6QDJayDCAp4hNgKZ+MEMSgjO
zFhCFALEVraDiIdZ5Nrs9jTEzc0LYLzff3mf+x1UgeWl0pQRWoxJEMR9S1vFStKdCKEFyxLjblCd
XoBEXn8nBAgAqhGCa++10Wx2ddH3yn1UFs1ikbEQcsOYG7VgZ6Xw2wagqaHe1lNfcP+JactQlJ++
AA2QqCv6tcDTpApOMB2OkKX65yJnjf8HSgrarDQVRzK34+HRLJXKL3kiMEeRHnjVtSbmg4zx/oQ2
iJLNMxYBX8jDIfWBxgo1zrxcs7oJpkK41m0SVdfLHTHHFE8IoMO8J+DmhhNGFb0XFsJxLns/eGUk
Elpz0PEcNlQalMd+8jiDKCrK8+iv6SNgrb5LJygRfL9HZ+awYn8MkApqyUTFlxZQBRxoc7j5oZHK
Kvnpg2Umk+gF78EsB56oaGmKpu+QJ4WrqeWyzcWZxtRaxHsNLDheO3vc3jqvg7BwbifO9cgaDmv1
RShRFIxXTmQdOfuNA6wiJv0k+XPgibWjodq5PEddqz0Hs8DEpPLwGeVNZroGK3f1r3YyjTE8Qyla
vQmVoRJ4h/vXbTFuiprKZ0AEqr5So93uUEQAQRCwkFWIafQul/8B4OrYXCJLNDYCvJSJwUfEJ7VW
ioyZxOG7FUmbTuvfYqeRUYc0NeP+km63LkUKgjiyfWl+QWwa4UPQGWuM7p3xomSJ9dWUH6y+194Z
lmG1Il4OTndRSaGTfdid704h3SRtyKBxDrZpN628JJzOICpVIh3qhDeINJ+iIumywGHsh3gMiy7a
p4ApL1xeLQQyWwEJ2/JQ699MH8caeTXNk0cDFDhqiQVGQqaYuvjAaiAd+xSrBnP1XlMUEGoOxx8E
ebAp0vkvSlDwmbmnFOodWz4I3VKMeb4/4I8cZDxB7SRdYg253APhw6NfEc6i2PBjmMF9PmLo7k3I
+ZHQvu3khPcFKp0jlXmp9Mstm0pX0OfoYLz2LFUXz0+WOhe3T5XV/9aV+7voggrH35ScTVsaAE1Y
nJEvdQGBsc3wR0jCh/2qwyvO1qhft9/eQ2jFkGTLFWxnuHlpZaaoQLXmt23lGn99rNTXzIPHHsHD
YsPNR6BPBPGW7o0swKBs4Ikv35DuO4SlRs8W8iItZEafVpXYWVO55rvvta21XjFOr9l9aUZdN8d4
CxcDsNHE1ibCx9dX8qz+3dQJaDhjfzEcFrV5Y43OasJIYK2HSWyjzsuaw+Rlg7p69ONtR7D5RhnS
dm5FbyyH45JuLkWZFZ9fenj2eqpJNkfwW32V2hrwZsxtRgz+eITif8K4zPFyj2N+N4nRCwQqpnta
6QNyDpi6wucLFHJBuRVZyWX1eq8PTSwKXAAjoSh+Y1IMUXtL31eB4KDD3x+RoR2bXxNYLzeqUK4j
dpalRyzwhGujSOMefsFrCYq22m7cXQSm0O3AbUwK2zLLVQl+vcsBGpEZs97hEAmyTQ83HswJa2/d
WzNUjbtdZRWdOdV+Xz+tq576kPKTazk77kZ8TMn61uGIQBDBldNU4mvyEfQbu40SpIbulBhwnBzZ
7+YmidgM1mHnQ1/MDKBTauXcEXvtTGpBD0bjsSw2jiRdjBnZTkpkUIhAG3Xlrn/WKRYzvoFxAvlD
X2hVdaxS+yY2pOZ+n6hWXuGqf6j1HX2c3WcJbg1xgfrvYnugpQmgOlvQ5Tf1MLQKwAZ30JA4MXkK
EIU7neeoIgune+FRZOFQZedaXm4zokjUtW+TBvQQbDgBtKzQgq7nufET9+3r+OLYcumRdGmYAv1B
YW2TVFlMkVbUmJf32PuaOY/wHrKlMHdQx8oUjnmnZdECJG++qMOObfmIaJiXBFwUm2wLOPUmQnsX
uKTEHo1ksBNvQOMly2emF5kuEAdBsBu8qJVGG4wqES9eV2sak0j69+RKWGdKA+H/kTOj4R+yKAfF
dbjRcUyP1NYhstMU+AcKulFZr1UFiGH6TlfMSEeINc0Xt0VvB1rqHKYsIXEcvyQEn+E2HIrH64D7
PwrQ9xa5NSUPXX2IuvF9/faJ8pvAaaSSmxE37gHVtXlSlz6iNnoqH3lUwrRQgvj6/uqpXLIXVrgT
u/MKjnakqKEHToEyjW+bTQ/YSUP1EMKm/PRYBg8H60PvYDDEgsEGpaGsf05PchKsQx8KynnhEn/9
c4o+j1ZSNl6rSuibINAKrr5gwun8Zu7fLip0nxGNkzbrHA6V8xMellat1zEFhD5GVuOdxjzSUzr5
IHk1vGMqtku7hIwaW9apgCcyH28iQQ2V6d1+OXGwEFXgZJG/cBw6j86cro1xYXQcqvlQ2AiV2YzD
YCO/9qt1wYdptLJ6RglYsQSDl0QUG02D5mxMCBFLZY6k7ppIrumJGfGDkFXM9lwith9ue+cc2WF4
m3dmsRYoL2VDS8ceIjJDTWBR5y1XX2EVJ1SDnT3W95scpE/Kqd6yHpNC6l0SF4d9NCj3iwacxfEp
Zcpwcy96GoAdfpsrH0D9/jgU/pMiuU2+T9nR+uGwH7E7bKMacPtNStgUesb+Mc7NtR8dJv23pnUb
uGw4cWUeLv1oP7s3HU1ETyA43v9GZDktgtej9YYKc4LpO9btbss0NKPdIJGlErc7ZdERat9Q/IUy
K5B95NeEOWsbyGgatftZktfB75yT4zVxBZKF+1GCKAOQnNflaZaOJpCSlYVCdy2lSDdLGFb3H04D
v27ztURU/9nIUqmcRGOq2alLa+MAXTh4kAVnYF2DisWqpallstb2T8XnWAxiV4owz9jEmg5rglBb
IE84TnLmEQ9Mte5LUQSHz9xcmewgJAvYksj+bj1KMQCa/Mm+qJ7vLEsKyFtCeMj1zAUJm4ABe9AH
kNtnA9FrxHRYc11AVHPMb7QYKT+zFur7MSdafkn9H/aZ3sYJArHd3jj4Xsc4JxXciu5Asiw5f/U+
8Td1t05CSRgtWMhJ0eMM7g1G2gSnzCa3aU0Uu36lO8188pUSFlXZ1w2Rf+mV7uBoHr6gSsmsWelX
1+e1nUvpEqAiRW79Y4N5Q696cF0RFmB68GDkIqQGBoWt1x6Ut/+MjZOANK8YhcSUmzJ8msAkXRLM
09jnxnm4hSFox4EyA3Rpca31JrtUVZrAU57wJWll63Konxh1KTRMXMKjgJGZHPkc0m4drRwLkunB
p/fK0mwkvHTtkWglVxPo/Lq3hP7x9PGjnburZdoNBWifkdXOwRDtwdID/l2M6c+SDc3K7olWDC/B
qVoPsDvktMnmoCvQ+RUQaTYTdnVodOcAK4iJ97DEjtb/BZ+PMmTLb3aMNj+a8bMTQqMYjtwwpq+W
4HI8k0jCKeV1h6MQxq++ZNLvmXXNg+XUYJlR98wM6k46vWEQDLRzOpDYU937t72lYZFhMtKWQ1zj
9GfftZ+k2Qle3XQ3V55bbOlFOjzo+S5ta4xvhhbrr1Vge4+MoQIYdCd/YargpuFJvmpa6Esk9LvE
Lrh0eIAIPvZtoYwl2RrkoRe+wWh89QroNnOChFwVYoMFMD1tEJN5yxY0eN6EnV9wwOinbRxAFvWa
al09ArHnfQ91ON5gW+y4pm7+EXFgrWZl2vUCQ96Tvue/q/yljHBDVDBIC4n0o7DdseSLyFOHQU4O
HwzwIO2jzCyzB+ZLgLgbLTcaShsIgXfuu1HqKirj+BZFeIxxKO5Dbtw/8wvdQdiyW+iEwpKahy+k
ymWn19BaJp/+2XMZIry++AuteDHmQwXGnd8I3Rma0r9zMqpg55lApHGQQqAvBZnenMnE3an9Wi+1
cbAGVMC5RMCv1d5ourL7rw9A5CMvEKRw56P80uiR6KPxbdmZYb1w7g7kLYdwaHQKQjCVnBqmYNiF
6wxPYUlnefF/yKObjMS7JbYcpoxAwLh5UUMZ7dWcXUrLF9adlHJ6XIvzDsgDslx2QBxNZVaNgFhu
792iS7wK5fceV6NGL0DZvVrGwfxLt6Gkb0jn9e1kDTgIaocl7oQQIQVt1NruZhGlGg+ohmzvyIoi
UTVYlDYeraukt3EinZYYYSLh3o9bsexet2RulB4KRR2KJOyaeJfZQGSr3mVb92QL/T9AoM3xMoFW
CNE7B/MuJsnyg6zGB+XBOF8iC8/KCdS955hvkcSmco1TndCJwwMTyaTfRjQKSr9nNdMVQ+S5CCcK
30O4AVqNRpX7ht2uCEswbeioHDnIH0zI18swI8fm0QiGQKSdCTETfqD3DGNPrum9n1iljm0O/kSE
MNm0BkwOdcG50DFEHqhtcmPQ0tEt7MkXB0pB0BetbAbKvbFPWp6lXM3r9wsagUyCOPWMliFHUBZs
wrqqwsS/19SdiKT6hHkyFVrN9ahv28NM3pclZv3eh3uRnFjhM0xkZdeAmeTQBsbVU+73W6eFSn7O
K9MHlU7u3z9ttqth7TbY//Dpxzr5mHUY+jh7hPP/oLMmjLlia7b4wt/5Fr5C+LMCh+QYkl29L9g0
d3vzrNi7x4pnPWIRZ/ywIyMinOk6WiBFLmeYARkOWSxx9X62Rcdvl7vnf4+o8J/A9cu/UhjQYaDB
VIbxTFgorfacQ0MFnP4NS4pnPNNk4xcSAuRIw4JIkW2vcF3u9a77MFno1gMESjAqiZB/iHe2/Yuo
H+I8aCGBxdLZYydZNMabGLQzu26mAZ4hch7UiCWrbSu5XzPp1tBvujJJ8SzjZpZ4gPRorb393003
Z/A3FUHeCmfwIgm1Arrjp4WGcCB2dkn1VHGuxiU/AEcS+WWgRjZlD1k57nJvPui9u7lRDiAwnM91
mz/Lq1f1KO87TNDFxZsP3IPgInwVs91EtWUaaWk9Cxl3Ci3ygPPSSOe533oWSevHI/X+0XJ9dffk
VH17dlDH5SQ+dBJ6me4OIpvFetWLs8HbPdxvPUkp4BgvinPAcEfJpTbVUoIIktTW/IqraGedx8mf
VnlWo9pDEg3iklSwgrPvrX1+p7Cc9QfNVXI2QNBVLVWc0yQ/mg9mOT76MskHZTbbJphAif+KO3IL
VIdCtI4an3Rjdv/JB0GivjvpzFlZMfJzQ+TqX5k//79GCnMgkqjzAoDnauDGYcQzxKwCgkSaMR0U
VDeF9MubgtEnidPkJs9KdhjRaN4R7cvbd/NbfODYGl7k3Fmokkaj5dteIPWqO3+2YRMtZwEB6MU8
uWDESikCZuJ7MIkEsp4kx1xHRb+N0TyREkwDnLiM8nCxlYQd4OBHi21RPWk+CZBOCBqNFeF0RT2f
j/98+ScwYXTvJ5QerIb5Jsak+Vv+wyGk8eQcHCyVKP11zgYwzCMFPEK+BzPbOkyj2uj1IAFJpBmq
lReHOHGI/f3XHGjJSrJGoWxgBi5S5kaxBMkThgAf76dtB54dnIDwbj33y4yvbj2H/nEk6wwVY0+U
gdePlHU0JGbO4hFCVc2P12seZdR6LMbcXSjpegtiopSKUgf5NMJnMDb88oeJ/0Is7Xanbn2VtLMz
0un/pZa8op5lHVrLlEEcYgyaehcGLvb5uLoHtBymuomzkCiLC/lgnB8z9OqT7Ya9EueSyyYxRG7k
tnloL0vznK5VoZYYy3bxk2yO7IpHQCmDAg4OyTVFgoWa5OYio8PMJxrvoTl7Ip0nbnmQB/qhpRiU
PEvmhRdGNX3gOcuFyeLDau08nfLCH/jRvKEiSwA9QXZ6FF1GXd7eKmmqmFxpDZZWmpkUP5/8BKz+
aR64z6N6MPiYsxsMH8WQsPtO6j8YTkSSLFzquwLCLMnHr6lz2Pvsb2vkrn0nvkotIgd9TdSI7koa
4inTnpoCnG6y8uLD+H64gsnaSuz3qtd45TtsQlvbfGS6n+CODT2ImYlQ7VVDT29jzmYETaPmePtN
YZLpgFJJQtE7QGAawdPEuuGAO2LauqbDFhiHnOIarFqjD1g7tjgm7nIihKbMrS25QromputP8GO5
sFBrgwFU0stTYLOHyGbGyZsfm3FZV7gDSGvBX9hvdv7WdKYZsXS+vzKdCU9VaH86PNHBIU+3buNf
QyzBdv5Nfw+UkxVN1/JAA9Pkk7RtlKCj/QgeUFy/Q+KVrHdekidydHxzedLw7zbSbxP30rtHGH7m
meUDlpVUoqq9TPUn0Me/hWZGZT5XkhlsukY+emUOyi9UGrjt36ENmDE0RV19cc8Jg9oQAbV1Wxuc
xpZnnzCsUYHFnu1nqnE1pPzSQq1Fi7yw/GU1eJHYaxW/FhfySERvuM+Tutfmn1GaPadr6r+q35yS
FRtLEtVHtgcM4j+vj2BNhzUBqqmXOl7M6jKBwfuAQbWCkKIKkRWIdz/U4YS/JdnOjvOiT6td5qML
gfe/U+wEWSPUYJzQYceg7K1YQ2ZejEE/+iBUVvAwdcfBWS5kuFbFsnSNhJAUcKWslgZahPcNBsgQ
lon6CeUoinQRQODUKySwkc49nERqRTCPW6XdvTW4+rbNLt54HU7tyBcUxi+iPKHLbokhITW5ge02
PLVgLfXm2f+OmvOxcmiIw6t90DpBxyhUmNf8G6spKHZ6Dri1Pohl7yFycNsSjzJRqqH6MJDHIgsc
Ai7wu3GtoJ4WluaLI7kvqE2wmXGBn0wvJlW7ey3Z6+MSyuNDXaGE48FBt0pEJj/ysUyG4GzESXQ4
LaTF0lau159R1DsZv8cXpLlhwLgMxEi3FOMIDD2wKqH1LwtgguaWzyK4eHgDH+kg0XQSfHnIoYZB
WySyWQBfubyu/3Pk+gB8d8h5/ogKRrnD9GrcIAxlK5xYk29XWgUFdEot8iy1wYjY8qBCBcdx5ywo
Gje3WH55XclCOgEAXrp5vn5xLdFoFb/y9hFSecUuRHisftw1MTGfUOB3G8QtCoGQecSGcLmL7UnU
Ztw+PWJaMlgr0F4ILIuIxRO9bA6JkiNYdLrMhhV4h3+K6rShkbosYy9RdU4azo5bPdII2FtWO91R
7osgLnSaaJmoJqYMHwXtsiKa2REn0sP5N4LU3eulqWo5nhajODBLguo3S7e3m1rkXp21IfnIT4ZM
J608TrBibrtDjwXQga2pySMpAepIxjM1qsyvNtE26iwLc8/ojHpXDYTpL4xUgtfckk6/Syi70C/7
iD+tMdeoxlrJBkEOskECkYyXZR8U9BZJsOq0W9yA4jRoTTcATVp2hwd8EqXUUHqVc26JwsTX+hL2
rdctv8A7CWhL9sIljqxYTm4X0+1LqSF6hRKR5Czo3cwlMyCC56m81I9Yemed5hwMyS8FrZBV1bSi
9K0lE43x0YJIXgVlyGYRMN5UbEUUWnEoqR/2jfiMenJn2UXWz/TRsD1afHQNNje9mUPzrsu4XlR7
DwIgAoxAQLRsZZ3qpunGihl58l77X1MKEyB9SnRoarE8YP9s5FbM9eTn/LHfBxju4FWS11zUpLQC
LezQT9iHB0tof6FhId4Rbn+8NDHUGmWck9pqO6cTwp4H8nG/VT2dhZIDyLY1kfN/g0l4Ov/3/gQV
1UozTsX5ka/W25IpVkB50E0EI2YLZX6OJd2GklLZZlBy+w5xRI38s2K02rxjz2V9rAHCwV/Cv2AF
BfXnPe83co3kzTiW3nxe13WowAauKo0RFLzul/EDv6W9SuCVc3gzxssguMz/ADHYgiM9m++qG7vF
JxCrUdP7SV13/HFsE72cktVq9FsOjOHiGK8vTQXHr9Pp1mVi9IZRh9Ycm2g1ai3HJJoBdHsNCVMw
UH2rgkc4fSUtbp6rEAN+yH48XbOiVdjUfnrc4nznoFTwDc0osPWLJ3HZbDUEw2mCMFs6mlpSXfhz
8ayCG3T4bnD3eLlvnQTwlKmsaRpT0mUoQr17PcFQMjp8vxAGsrv5v9cU0K7aBaCwL/AOelCIacNu
BFOGKC2r2YYjL5CEslgRUet+6bYf+4B2tFPNwO35WQpHQgxULOPhQjE5YUKfKJnjLP2A2N5hHlOU
cc59WmE0fHNQ25zZFnXjRu1Ppdl6a0P41UFHeZQngQWGOGsKB4tRZe+FQS8l6EK1nDqbWAlNJfEn
tWqOWsbQ1qQf/xF6Sfa8iEaBdKbAKxCO4NDJtO5iPAU1i4458Qa2+bq1KH4JFtc/ntfTgKoBl8C8
9nwtE9uqpZGJAi2JxFBa01vYOxHqm61EUy/zIGXvf0wz3wFCCnGy3svjzsbLMk9ZH3vmAviiRpUi
KTCaQ7LlCzkyPTpHNELRwOtRA1Co+vOpAX89dtxzXeu3mzZVCQI09inEuh2pP7vXczBVIWZMKjAD
rN+c2awoZe4C0Uh1roh0mwyCZDyhyGmcGr+wC6clcIieBHel7NxqkF1jOwULyi4cTwG9k0bAUpVK
vDB3avEKTb9wjdwYGQms0Va79wNPSZiZIGu6dSSQznVYqLYuZ5D2IOYKT1JzMm18b71QpVp1V770
8y1WbQmVk4ADdFsXuSiyOrFrVj6ewYeqagXlWF4APUA+QWSSr7GQJysxEvANr62xKe0fEjXpWtFg
YtTU4M/QV1AAWyNR8txy9FtFTWGKhdtBIzWmINO8Ss6oiDw3nk1hq7a4tPRyr8Xpl0qPCZAXg3zr
coCmBVV6AFbOIjS0TACTMcmmwODq9SvPgcP4ugPehvG5v6RvMV0kIYfav+ILfxth0z5P76Eo6b/a
rTg5cuoYeO9xpH2vG19KNBwnMrYVjy28Q35Z/vnTcyM+glcSdP8nTClD3NnkBvLJVKYmZqocRWN6
RNfy7up4rTUBn/yi0N1c6hdiNSaqyJcHEg4Sqom4DAu3zrg3fEWlUiVunhWRjrWcR1qSeHkxArHX
dPtmJbvQ3QnGjX0Y/YMar+1PxkdSuMfBQl9hZMO0xoGt7eNfYmCisveyBIQpK1bXnXlDmIyy0hn0
2rxXyh5tQYVP0vHaRRvIPY8sRS0Bp/jnOx9MNxVdg6BxihDDzU+SJf8U4ga4P9hbEBUEvuj2nlOb
oX8xkFcsWZn5J5sXVy4w6tKtqcexOOpzQYADIuInqEK6ojGEIheNoef0SlYQYXrziFXVdWYKa2KA
IVCHmn7AZJERpZW1RhmIhgKo9QcjL9xKT6O84cBIRLj9duz5f8FIySXccHmHMzFfPSs1SHhlSPrR
lcXi8gTZs7lvsHBou1fKVY1xw5itBzLENMN8qSann0j9u3HHrHlBXhPrdkm55wiHihVeeDByAIPY
3lpv0UYexvq2dBbMOAI0c8u93CykvCC7PkrBh8FKuXRPw8bvLZ8eJZh/xeowNz/QwwPQ/Mn9vvMI
2ddLeM6ztlKWx87T9dBWqrfFejN1aWiEHaOJnwN6Q+rIkv3kkCt+zcQwb04Sw6ZcO29HA3GJG3F8
iia4r4mCh8+61/ncDQUrsYQZPzUuo0igha++Rh86oFKcYd0axEpeARS/E80X30bi3QrtUs1Mjv9Q
w6chDakXtpIeDEd8FwvBwEiVxDf7G5teRwdpEh88xjp57v/emoq1YljL5bPbv1ldWYmvubV7CUDM
RHKYqJL4UHmwqi8S4Kvrugo/hydKOCMRr6iPQy8GTnJstxD7w5iqgIDof6dJoW/kwjszWT0it+PY
uPEtoyLcSe+VqKwlD5SbMVaGecwcrYmuOnR08r+ENYmfe36MkRTVoSlTxuR6FmG/IAfaix/4kYXe
1t5gvHC373da9eGMSP7r/AypMb6He/jCPwrpaJfPyhkXq4v5txLFa0P6vMNLaZNiOJMP2D0qWKNa
GTONEeSenahijSc26UufioH4PoFxuxgTb/JQpnEJU3LU9fXf6r70lwqwJokR15rTcn3GIlraj25g
I3tOBbtmklPecRaItKavZzbPu9eLlrZWqy8K1wvLuLWUD23oAPmUWfmySB1aGQETFoZmXKEIffvX
YQ+CqWqLU7iICCybNWPPS0JbgVe+2NdVMEAKfOQAjH1JjWOhpBMnoG4dP5d6pYghGkqdvTy3hCi0
NY0emD+sH3UePwZFWbZtPVscmRYvpq1vnHRCg3oy0lEg0kTt6FDaXHXx9o1ME1eCFTwDzCtThjfZ
Q9/vkEdFRdU7XFk3kYtvJqoejrZJ3CircI6XSVfhMoGBcJBSgQEf112YXNUhdjLPtxRxn/G9iwV2
LwDrUTHJgClC+KgmqX3WtHLRzkulxKocID4h4c7bZbXNs3jdf0+4EphbADc3mmIAbC+2sUmwY5Q3
5YbCfBcBJgJOTf4zeEAXJD6LbrxO2V5tgaF55Iukc10OWA3lpZDuLXCcwzl0DXZZzoPb/UOcDXzD
cBDZC/8V8gX7PEohB5r2gFQRqcVvCHUiWPAZRS5ekX/9XagBLFdApx5/2lipSfVvQe8Lhr5p3pBU
+xn3Yzt6jiJkSDjgq74rK7ztbQqcZvb6FkmvA7X2KHGmNcUdEGc+s/Ib86c3zTngkjABWWRPeEV/
kCxtpgCYUS/+GWxUsVUwk9be/oF4IkWk5MdXfD4b6ST7oIyEExGojWcLAXshFBmfcCiTSkpHmsye
6c2UTbSIEoybkXoGtAUop1VeNKnA3Kd5ogBb352ae/S4swMI0H0QDdYc32pz3GC/HbyXuWVklYGv
M9pVIarTwsXctzNk3/Vbu9xDFQuOL0TwT7PcSWz433jjHLynwpghqcBrY/X//Xlj/VTijdO7j2m0
dm7Cn2eJoA/4K4mzGRGVMhU4W6zgOI+qJV4KmcW4Bc/VpOuOZPeOBs7AX6ORqvi5r9umUlwO0uGd
EPUfIezMlJxV6+6oMrrn3nJ2j3ADb6ioZlpyHmXCL1+OKNcbEOiXgvK7tt6eEU/SEjGkPHxjCrtK
5i3pVE7fqalf+d9mGbDxhOAh2N57j/7qxF/7moccgglfN+5lGjSFtyAiXFe1ti4kYFg0ltpzeKHD
WU0k9R/ZKyvm+z0ybwPgy+FIzX+hDD3WwRBq+kKT+NnCMpcn0nv2m2SfyAcNGJGPDbCOFai0ZcwR
hqwXIMGyJx15/Ey7etJb0nXmrFCqX96iLhRRu/b4zc91K2PVCva81UNlDin+FlnkngISc+dK43D8
kw+GZD0n2Z3qizwzAyxuFgG3QbqpDYsOoYs/l9k+SoDzG2PIihyf749LN61lQVZyLr+Frzt7nOq8
yr9xyMC2rFBpRNsNsOMMwql7mT2UK90CBPJhra1N7p8JxljMi6DZTw5T+TVEbx3Xx6zrl8Bm87ZD
FFaPujyL/+stILGdYTK5EgL8+Vlnxj+EOUAX/bc7IoAcl+yL6VWaClnYSlxCjcGcpRajtiExPsZB
WwCFGFb1uNaTs75dPJtu6pQF0B7GAZMHy4uT/fEMLFL2H7H31jPnFR4aUW/n39uzab9qoJ1w4OCq
/lCuawM5PgIU8S0OeP3kDsVL2T3wx2xr+LrtEJu00R2uhEKChkPqWkn1N+04EKb6Pi63Dos3Rku1
BOFVOclRdVk4/E+KVcNvs8EmEK7Ljd0k71VWGBdGaO1cBroMIkUUzW9/uqn6AZTM7JEPt3FG8/kq
W8QFmKbLPD7RCdpcR11oCqS5eXs9Zm5bKqoNwVli+Yjs7+MMFjf3nAt0watNNlWb6fVZ7QHLDFv3
+kpMS8GezQs/neNkfOt61wjkGWDX9toihqjd2PDmvSv/uzNOuqrfCT31wLxD/UANUPbb/3+EZ7w2
9BNd4raIUYGTvBkbQBpwkHgLs9cxTJ0G9y4Z8tQfp5u8hP4yWtMUkXd6jKfQ01MeBLvOJyNAp7AM
c6Kv82gk1p53PFcysi+FHuVwJ4Nn9EwDiDhsd2vWg3uPV0ARRVA+l5DttionOdVAP7N3cdwRJZqY
lCFWfysTsGLrG99yebxndqsEM5Gky/jS4jR0MKLJ2Fl24nvLm46isBa0vD+4re2pAUEbduoQ8PJy
BUq4o7jYbx1tFfQf2OFCi+SmiVK+PNn0hmKntZx0fs34JyCXji2JrZ6OkmY1+x4s8wya/W42aGtB
orkc7TKHzl9TXwRWdoN2wtu87Hw9KvL+W1d3jglM/999jjcaGI518Fq3beuzOVp82zmSQ93LZ2Yo
vIkR61XCxiUDs0WebThJ0r+HOsguwllDP8Lif65A4dGYL6ZG/tPEVVn3niqi9yKr0d28AOTReetV
RMkEpzxLUn9nJXGlxAKdV4moBwiBHt4CYFQ1WMsjBrjmACGc4OwOSLsMqvPRTnsxAW1Kmg1eRBx1
kLD7pqNkotlfjixi1GmzYRwF+GT+HpBLy3EbM9B0Z4Ympbm8Htage6bYzVtNe+nDM0IghzG+jGFx
R25WtpSTgMsDQbWcudthwT7SDgU5wIbNnZL9P176IhTT7ZOGN5yGtplbj2FqVydCgyYvx6LIgp2a
ExJGYsInMx+gQOyLGyhPrl4fORlE5nVIRHlLK6N9JzgN56LULs28C/+r/teQrpZ/ECO0RbuUfPQg
sCnIfQfsJHwWq3lysV4Mccqv728g94mY6W1sIzy3W5OkjxoOf2j7f7hfWSTpBLlhYd7+bXWjVnvh
KCe0kD51aXYZHeCxx1Vim0qwHx3QJTEPcR7nj0Oof8oyi7Uohr9AFTS+QXq+waarNl70VsqVKjWM
f4/VARf+mKqOdUultDJcUCFLlGhMBOpndBu7e5zyTr1dlm5udRya2ZqzvA/oc7T2jxT3JgAMk0c5
/gH2Y7uyfopSgJVpuuHJqzRFdnk8BQhtEtr8sNt1pScWWrlNPVnUckzyYt3A7Ws0MsVxPm3/k4tp
+EYf8HF72GGj9V3lf10auTpWwdxtwIVkunMcoph654f+8Gsb5JBVyYgjy+DMalzZA3vrNdpqY+9r
0P6yWVF/VWBTal9i21ejHKfzGpIvcSO12R/KeOjtpR630fLBi7KsGDLC0wQi9ue7DL0lLlJ7kOZj
Z56TROGYvFbji0PaY+v4jmP8eeiu6ZdO7J9fQ4jt+gGwab/NrNZXlAqa3MBmJZKA18xdXh96g+78
EACAGOpKYBqTm8JQpMcb8VBCVX6THVeFlsBdzIk6eOe+W89cJG3W02rp8Nyh17pwn7sXs3x4g3lv
QD2LQojQAkGdVlq8AePhAQQHh+cEcJYWLcFcBsuTxsfmy2HQ+1vK6rBQm4ELqFpT18migxvkT1K3
jzUD+RPhRXHm6YTemCn+r+s6O7DTUtPKJubbh4FXd2pd6FB12c2MTxaDIGgxrzmRm8Ji6/9jAm+S
EQLxpvnwx5h1IqiV0u0YNVVXPvree1WgkHCxbT0q+UKN47OM7HDdU1ehEIDHv/xyx9dHpHNn5Vav
m9G3ksry59sE/+BJAFKdBiNq9tu3x7vLSrzI9viByozmBNoJAO7ler9xLsLY3a4iP4+WdarUJhWb
uUJ0CW1/wq38qQIqwu3ZGWXuUblMt29owo6bBTU84AKMuxa7r+lltjhMAiC6zRo3/k33awTXc/G+
Eos9Mpn7Hje/DoEMCIWgQLx6IK6cyrCRewAJ6ZmX/lqYGRvpSskmAo9tfalL0Y38UoWELYrxgkk2
1gblE7kJHueCA6BI6qlNOclOPUO7RVbMQhP8cSN4ByFW4RCaIzLCoj6g7DaBpzFKlnZsPyNNlfxU
9tTNqx+4KpbWawI/25rmslHOcCecv0bkuSwaG4OotkPp+s2VoVFnmHd24XtGxM9qDwVdMhaUW15R
zLxG60D6KkwDauD1+ExEIw9phpaTttFgKsRJ61TJI+N7R/F3sdxhNRZrQhkIm1YvMe3wOz2x5Nla
oi6T2rI8pQn4oND/ip+B6p3U4AlTvkAv52zJy/r86IYkwv4fDjCh/sbDxwqHDtMY5wDogmwmE5GS
9FS5q02ylbaj+bREt3Yqos6rOVlIxiPMlQaGTnZ4fhMqDZww00rfvclywsE1f34Lyf2zjCCSIgyD
1hDluImO79Q8L43X8lNgNY9zxBewcPSjQpid7Dp4TBjiHFrjsutqUMpaZY/jqWNyv3DyzXpaqtJy
jGdnwaX0MTUK7BquDzNdSUS1IBgAscb+l0eXgeU5UbGDAR+NM7qCcZd7Ng7nRacHt+RbAdC6IJgv
FIL8skVA+gvmJCO3o/Sja1QxYXb+sPo/0YcM9sJlA8n5sC68vZ2WfRlwtN7z5XG9d9kGHQouGKeD
5G8Vp7fxSrghhgcAOkM6Igv3ILhz9LKOeLz83Fjd5ETq9INkWe6o4z4SYt0CKdEqVMpncsPf3bfu
7aQOWrh38nIcYn46JLHM5+k+ZKIJaCPQEKdN7eyaSeEAf2VIxLeg0/E1LnAMP36h/AOS1C7sBPZ9
vS3Ixemcd3zpDL7aEOP24KXhVADSVnCcGIju6oNFjySodbpDL44wOSmZ8GCKgiIvUaoT0MPjUFyp
0SrtV6lyZz+ySEX4thk2Zu79kQygWB68J3ZfavZtf3uAwvo6h3uGILD3lRnQPCjURfkfV5DtHXTq
MT0Y+WKbwX+GRP3IVy5nLd/+SJDXypuV/7HcUc/4/2KtaowIBQfkCmhu8Vg+HHhQHOOqO/mKGEuz
jIYHFhuMwU+gA3PrqGrZta7/NxbHni8UJXkczo6xW2z3NuufQ+h1fvYBA9tW4CZZ3gTIQdTZeNBT
753iQNq4hbDYKg66JFITE3FvGjqR9DAhVrvXawq+6qazrTN/R7gJs5hZCfHsCuOupJ1vqhair8io
qST/T2VXKHwxXocoIg8YimgPpwrQELVl0j4CnnjLzKPCjGfE2wUaiqyvEBAwU57cb5cRzhWt+j/7
AQivjhDigjbfvfuY5b1xpIM/M/mxkr3Hu4IMPx60bU/OWicqNdARIh5ScOMKtAnu+qv1hHxZnP//
6jALywZSbyj43AciJhynhMRKeaPXW68bh7yyJu6VPrfiesLAEmxXicE+pkym1cQd0HsxMHbQ+QCE
ku/gCBHOsnOf7jQ0j8BaNSeZe8O41ux0RPW6BMGo5+Rq8VJO8oBMkv2B1vMhjcKEgDqs7pxcqPSk
+CLThXwz255njFadJ8+kgG/Xlx4FpGridyKHIS2BEyExKH4+Tqh9ZCH2bBwQLM/E4qY6a1sOHyqV
FJabnTliOS+mWG7ZwHkU4LmnGCqMdt+X1Q/pYyZ7F/IgO+0gClE9CLaXffjoXpIIkYzaXKyPdsES
caJcx4LFjFKFP2T9WWUd5oLdNFUiB0+9tUoNTIKBE3TVKwTBYP4Uk2Fh1OEfX056D+YmK+M//wr3
IwAPWT4CSuIci0gU11B6vmLmAn7aZ7Cg6x9VPC8tn0FqAzdIE5FaUG2lbb2CsiJzfwQr4kVUBbat
cLFiQEMtAikGeiJ7uzj5Mfj10DCedhO7nn8x3GoBE/JyHRInmh7H32wCRYLoalg7ioX+DtDgZ+NN
fgBmmDzRgqo2wtRbftI/1ZmuHb5eWNGrpo2K0TXDjS5MjD+6MCBXiEOUsIk6psBw8I0+Dbk26JyM
rkNI8vQ2LFweUbHdvm52IzG79G9czzxiOfr7MheBiaKVBFZ6ldw+FONkSvO/ZcKuQiIOYiyZM5LI
Cuk9JZxmLMSlJC+55KJ2ruu7Im/zSwvMYo5FWAgSE7CH3/jqlm7lhOyG+PyLSy22eCggUt/+sXG1
1u/yxKmFyfWkHOjDYzGD6gdEzPkQrFV+T6Fvznbje8yYaaa6CtD+ThbXHN1Pv1CE2wqUo1lUnWSU
qUFdRy6qM5veeeWQT3zYTGJV8pAU+Ior0d/6hpo0HvvNa+GomjEtW3/E/Mu3G/klnTpEBOI3hyhV
4qQx/m2W3ohaazAUYjo6CDQxyzuWGnKH0LREyt0wdpvPqn2Y0zG7UF4XfG+ybTOFnhEIVqtKYC3Q
2oA/WqsIqI0tflt1TcqFLPSafysefJdsGVlmfJ7jx2E58TIk0yQjQ5pZteF6MdGHD5Z2EAjgKpJd
+n6lJUIbHIaqFZephNwOJLb4vDw4IBCWmKkEDw4kN81OqH7qWxRuJneCRHsDu6vu16kOA0isLeio
+G2+2y8fJTf8vom2KCms2HsKwfGUVeAk7KmFw8lQvCeyJTvHKX/ba5Eqcj8E10uPN8Bb4NkWjui7
E24euQdzgnoXlvvgI6n+pXMVBrDwVEZsn32CYo1H0B9y6yjypVoECUtqnzIgUDEoiMbsUUkDBP9J
WPsE/vbpcM5yAPV7bfqSHPGaWH9YiOXfkeHUWsHbuTn1dELySH0mqWFj/tmxgKrQyWiKfsvBQ8Wy
4Ehis3eKAB4QIyMr9WgQXGqjiVr9iL1bJwe3zFH0wwWKLwQb2H7ssrlgT+m5sNEHtlASZ4melvXf
Beq+uNnXXYB/U3VGn6WSWLKbmyjWMh/V8CnMwU6VBL+7W1nCwFJk9B4b8EgVP+q4QLVHcfEKZ8ha
lJHz/qaNWzMDBPSP2bjLU/YDnUF552oJVlHGXDorCRE7udbjx9ZnrvYcxkZbBQ4EoKZQt+hAwFcI
HdGjSMFZaekuzzthmOztH5aAif7xfydKnR7l6C9h6u0Q/VNeBwW+y6GyVbMKnIkw+8sMj6T/zGaq
YsZHDEvS1ZIolcVAacDhJ1vJ2fRpgKfXLYWc3DgSVPJ41kp4j8jTW7s6+I2bmeiKENe36iqEXeqX
jL8oZTHNeoCB86+scOUshLPUVJY9amyIkR+O7b+tGa470tAbDxPX559TZBisNgsvQ93iIdVGXQB6
8qutCuP3a1gK2JDk8xHkL8JzTM7MOb/qr05EHb10FJN2zhbp47fP921Lme2dIjzwa9NZhaD1gJfJ
B1J33zRB6Oa3YwMUZHf0gv7yJz1xwwGsW0FrIs8zo1sJR0ghpcHqDCqrXsGv5dNrfdIebJscZ660
xq14xMvpHxoSzivr2JaWjxjzMDGzV50FeqR1k/wzoBYJvtVpGZsbe9LlYaEZO1z1DxVH35lPWiPI
s0PFlbfPNxI3uVM5Vf1G6ihGhF2k30Sx8u4pfTNb9QA2BzUw9FAVv0sJes7Usgs6MrlCQw5QXQ7d
XWWYL6cLGKyQDr5R02fG6MA930oNBH1EhQX0Te4hR6P0JAF2Ql3WJ6EnA4zgmskpisz7IaGv3/pO
K14wp7SuLr3WuTjaatgM05LVojnj2oB/ldBflrhG+GNBixILWgTdcYwhQIIRvah7AtWlIMkWBhvN
ojTvHDrkgmw9/PtTpqDnW7t6u07dQbNxVCWojkO21Etgpkg/KK4a4wG57nJp0ZWg3za4hyMDyAFG
YK0tqgRs6rmn9k5jLB1ZEM/pjxVjhQqQtpIZcAkM8VpwoCyrmKr7D2WvrNdVLQQEFrfxtufUdqz2
Jdl4HCBMZ/XrvvPwUee3c8sWD+RnuU/sxeaXSsQUeb1MB3p/NGKNDCTOjjMvADoMm/eIsBssu4z5
Tt9pj7yY+oU8v9x4So5yPSgtkKXSC3OsyvYzIijFA3u1gJgA85MsVXtJCDf6LDz8SyXOftuKKhIB
IgkfJQBYLaSJrfppdDfXlvgOUrhtylYoVB2rcl3L6dG2/3ZcrQR7gmWi1+0T9FpXZ63/jBwYE6We
g3YropBfNxgGJxetcBWDlZQ4zBQ1JzcA1tQm2idqGLHOjCUnz4T9sbRio49G5ZxgUCvk4nnaoJ9f
srsGKl84665HncdPD/oP7Ac8dwHXvXpuR2Y6C77d3eGLhM1lkjZt3+4wifsL3NFoUk4WnQjzT4yF
CpOwooHopEHOExZX5bFujs7+OKTT0QLDGRUoIV0b/1+AATeUCXydJBAcgrtSJPzgVThwRIArHZLo
1ByikF2MuUNj28tjIL+7M1ns/1cJA3l7SUTdEeDCHvog3KVl8fHp2+yfpbvGTNz8yrijJKqtgS/H
K93nGpk0NHXaAluQyvfRWaSd5IxunThmSbw6ajjzY29H9XHe/JFEFkC/cg8j73CbMikIb5IXfqqI
fa7YNDIsBKbyIt1xlq49b1M8DMmhbjyzg0H72oKJoGPW+dZhvhadBbJbR6UjLlVLbJVwmtZVxv/W
Mbm5mQLsiljDAt6lZWyTTn3o+VvsdlM/tj6rus/zfiRVbusBYbpnwUmtNxQzrOoEwXSj7eLecQ8y
LaF5hicEZSfrN4sv/ZLqJIt2coRCIihtgU2gOOjJmTbazkPB7g/qg1dK+UpCPWsKUWK1KLOahZ9a
fhM3lgQ8Qz9eEMPcQrVwu6FUWOa96ZPHFTN7HP6GlRf0TzkdXUFCP+vNePMzws6w5ASOu+mNmSwi
4xME7jASrbHQf+5zzR6JgBVUwHlhAXMbslDRXWM0OXGWtoSuDof/LeCX691jRCEzO8C6JW859jiJ
3m/j6YDmVBUT7fx8Y9B0iQWLzehF5HUIfxYUP48i+MmR8xUDRf3QAnN+TMMsu/63hatQ/VB5Nl9z
44zEU1tQr/75JxSqJre1d71Aupkn6Vhh+LJ7MyF1IL9vQVr+sqFRLeojhHibh2TuDYEgGBDR1+cK
ZdmyGt2Fj44N/vEiU9n8QyovCzF2qaN38prbPl7fq0hkkQdkmueB/1fBMA8BP/RO3uprGjpZ2jxa
GpJMjf420u8knXZbI3PdBShee3Qc+sXdnZNqU9eiOFkxPRop2AJqPQiZRGjRv3TRAXKnEynH4whc
zX8pENQ7s8s4QxxmYEwy+iaZLbkGr/dwVLbfwNklpkAKQ67lFjpJaTzc6AY9ZlbyXSqW79iuPP0J
gvESwRSD5HATNTsj5MmR/r+YaAoxNE3YW+vBe79hHCLkOU3chRzqsgyJaB4ykiud1rJSJ913jeNo
mqCLihGzaiPgkEnx5z3L2NA4k2z6XsxgEAGa3FkyF4EkMN80lpMpc1UhKybcuyBsvct09MMrnZBG
F+SHTMoGcjeWZbLMlMNLHxVdu5yGKKVmXL2uMQpIgZs+FgX/4e5ZwrLf8aYSU9fI5mZT03qAXysT
mONtEbqoTF7LPuFmS/e9GkFb05FGA1jFNvbZ/i3Kjqc5sxszKD8MUVU/F1pQWantoeJJRbZsNiUv
vVPq6E0R0W3N+2dgHQZ7An5PNqrCVIh+hE6MFCv1zqIDD2X34BkvlFHoG6itcqvqF1xGhKbdxbRi
3WPSPbzF2PPGV8GNSSqVdV5Km9bvyxi8AE85dfkWIalukothVT5kHguM1QX2IxZDj85EmL+Ea7Pi
oH0LYbFhfrbs7CW+ckB/6SgKaonHclEKoIjPzUxi3FEqkOfAFbWBBG/YGEkfN6HB/8X5tdX09F/E
nqQJoqzP5KTlgyEGW63SX03z5uAssEfwTFX6R8nOrB162zBJ9T7/Pob8VdB89cdiJCTYe0+t/fw1
ft6/GVzEhqQ0l0wV/44uxDxxa8SMl0L+vt/kHKesMENmabxVOAGyo+FVT2ZqF7/O7BvlWALV8m5d
APeXIcz0Zp1qL9s6SSSjI73I4i6pyV1Hr/TKmUz9qAuB7+x8oufFcD4YcObS09X88Y/mN+6d7bJw
vaAODngfZimglCzqKTXoFxbEkr8GugSUYHSgiFoDrXB5AjBqbEGOJ/8h7bGuFoP1wHErpFeR8OtJ
MDyJ803VnuiuCikYWcdbHbEiLmNaQK0+HNF1ORh8LdTLXRkFbXv2Fpyx7VHbVgkQ5uttrS7Osy7q
dN+ggsTDJGp7w/ci5H+jypq+ewaAVR+oh/7fhYRxnbk5ISMaOUgJIgLP1feEPmKKPQvSmoJQJMNR
LiJQ4HF9F7jiEK4BMPS/nl+WpbmmQ9IoETWTc6c+UCllf62FwI4WPrCxMEEPwnhsM6k70jC1toGi
XTklfOPKWmY5N2fdDk4K3+Wsc9jpVeRs1nLfl2Wyk/9aYfdHFnz8+nFrM+0pQhQDkoq9vLT4b8Kg
4sUPsk4pbo+3VFuCGeQW7u33JieVi1vBqqTWsQdro9tPSpS6wv7fOC8ix4lGZ+k/xATRucf4jT1U
8pMSXCVFFtZv/oZCA20sDqrRb4rm9nu0zckFyhM5+kK1fn2Ezf8NeJSb7htmrOtFoxM9iZRn6zBZ
Bs1G3ZqVcAFshYPPzX9nOuCL7wGM6e3MjUQTcO378BF/BjV7FNwrIvHtxuF0CMfwPruewSigHqNr
56iw/4QyXOZ5gzUkV8K3OJkgvV7Vv3hazFjKNFkopeCERuVVJEZkWWmkd2Fcv/1edOFrecOhHepl
Lju4lXhPiuYq6K+yCIdnGBTeUbBtHQJKs1Wa6s+4reZ1FQWK1CHYrijWgYClGiAL1W7OZlINIWvq
Jm+CBY+Mt7E+hXDU9fGNv9bV2N/omAz4MB8w50Ya+9pvI4KMxVrdIBLgzdQ4gKopBp0qbV0hZ4ww
84/9nLrSOPXQQOh1Z4+a01AN9iLFIwPKBAKf9jNzo54THFxb0goLxVTwIcBAAez1DBPPYVDgqsYv
ez/f9Se7Smdc7JmZdwDCazmW5j3Xat4AavFU3ImsHZxa0A4j9BSp967dfpGsIUpxdu3BKfuWWgzx
x6SwTaqXSLfuBQbeSjSk/ZPj5AT/PviL6CrTDonZi19iQW5AfbognjkujGSRg1qOAMilzoADS7Vi
bHZT9YcPqKj4/+j+HVi/ncmlYyx44C57rYkvGkB3oz4CxzFQFnykOZIq/3AUqHtffuyd/UBvGiSv
MLOpBRHYjUp3NnxDsafJ8LcfLyNia81KfT8bYIm0guHIe+UvV2ER0MuwtpsX/w8NXivY9R3CVW6c
eE6ktakOfLA+91qYO+9LuiC+akzJyapUg+11seiXu8y1/d11mHViLSYN7uRhyyRa2WriHEuARNGK
DIHeh+7kd/iWKaPIZy4UK3ZFEDO2PdYb22ivCkr9+otZK52dUDH+DSKGUstF5UnOU630D6k49j3P
N/bR63Y7gy8wxqNWIYwYPgfugOzDu9zjNJ6781gQ/B6Vy8cOVEuTQd9nXtbWGX1/Bo8wu3FE8r9/
3y5LebONdO6pSSIoSAd0V827I7evzdvCpjsU/iJyDC6gdg7WeL7Vlj4cu4pNLPLpfjivEFSEirkm
OdllzqL8MYE6ippFWvRe7xIn9Kro9AL609qNXIbIhnesql2X2pgbox/jeV3Dt1BP7CIn2SpEKrlK
yPsZs4Z3dR9cNlaVykNKmnW+sc/FXR0dyiNV/ze/f7WyrxA23gVPGCFJL3k0IrN0Wfp3v2cvj6wq
YjOF0jCKTNpj/67zshYQP28LIL2+9n/GVztz7F7zHmlkJvDPnJiAqqr+uK8PkdMLeSCC15wJSTqf
eEqTQgyS6/XbHwJorwiB48TuMNAzmOdSv6GBxJGASHHM7exEN5jFJRJCp6HpCxTDDbngpljnCoMp
iW/mzFEK4b/ZH+ePuTku7WXNFuL7nye0aLjjkK84NcXOUS0Oyp91COwfLjFjMXOcIprVoa1Pow2p
bjNMX7XfZL0TQY3ts4KiN/qVSvIYV54Q1Hnh0w5I0sJOmGuryLTIPAUt+YVtUOOcflX3MHNPUjop
/EMhSUTXYmUHEUWmaR2+ec49HFn8cikF+okVoKhiMrJRpHd0OmwX+fbUU50/ZT/4LUObSulRejQX
R3pd6l/1mW0BLnfmGfnYwKDVUGF+mEnySVSM7kI5j7lKtSVSKTiwN8U4q8npb+RbIiiaBPEFhSNw
AtrCNZf9WaSdgPxlZcZCwj9PHjJrpMSGyaMGIkOfAIudqwqgQGyhC2etXhGxpp14CSKiJ3wq8ZTq
+AgxxCa2J/QDjgnH/OprIUwseOWUoswx0mwMso09SxL4zl3WSwQfWHjwQHjQvK4A+O4PCRphyYIB
Mhmo1TS9pLv9QDEzf3PltipAm5zlHWa8ifME9h2XEROnvb6rkcdHOjvpihGMur888TuvUr9Di4Et
3GT6D6KuwmwpMAw/lW3OW/7y5RimEBCObNaXEk/0jWge4JL7PHjZ9SYI3HvIDEG0A4hPDzCiWQby
WHYLLGw9WsRbrqC24d2ocZoLqsqujSTnhf917b3KwV3rnhrNLPGquBhv+0jubyJhAYlhymqCLOgP
nKDkwfXBuIbpmIbxqIXGVAJBUvnxcC3+JsDe5H6dSGkXjgXplXTa7grW436ejOBHAY7W1F/pDBlY
ElOnhtNTdV02bNcO7RMdgrHlfb4XgzuV9sv0EmMW6bTrTZbmi9k8YJVNMX/pn4x7c2WkpowOfdtB
5fZ5B8ELTgJf7mIEmTsa/kuQdAhMfKLwydwr6gaAQM+zrc5Y0cswbKMM781Q7Jevd6aTpDJ+B8/b
kblKRE7SFLTTWuBbZBsGNaWvGxCBenZmXndr5gRtyD0FQ1LHzzs+YRcQv3mku2bcaDzVVvUCTTzY
MXxsVZrugSM9xAlspRhmC+VDCc2OS0gOXp5KAWSApVdrW4ojUEw0Lj9EFA0unOrU3bgZd07xHGZw
wjJlJ2iZ1GDZuLWYTF7d6ntw8gr8LL7IOdJf2s4L100ayMWVuvP5ZD+19gwT/Y0aDDh76jHeJjEF
IZ7WbVsR3vO7uO0Eb7uGQK+r6t2nYCjOY9lecof6JzyHrZUvLqgXWZD8zDoFBdSWuOn1wvrbCo5U
ZC/xdB7X5Hh6mftOny80A8odSxCPq6qu8Op0/8LRjwt6UDxQ1yEpfIPCJT58OHUfiC6qf50neoKx
I7HzyfQ87TjrUP38AfhAjKc1M2hMrAsm6MjB3+kcsyTfoU8x2T189LBDAkky5GCtnweKLFOa0Bvz
nq2sv+wKjR6IkwCO5/M/p1J8QZy8SLTZB0+qu8PuT5ImJ9vdlR/j8ffjheTt7s3vQRxWJQUrqgEN
yc8e+ZnI/TCzkVUDVeWsXW9AB2jQJNUoOX/3qfCsx+Uz3ooRPkCs3VvyedkNq34ap8TzA0qk2oTG
092rSVhuMqblWX64AzvslMr637sFxyBHVZn0WagPLRpU0MAOYas19FLpAxSl5++xxxF+WhOfXGai
aTcDt2OAgR8ZwYbtUPOZ/tqaN1bvs8B/wk0P0d4VhYFCU+v3uGPtYkyT+rGXZs8r+6eSvFeHnsmQ
1D4wGzerOLjzqwJVDZ5B9HJiAgCXKpJYm4WPSAR9SBQKWpPIdXM1cXtC8zT0/V/Ti0h7jPc8SGqb
inzoOpnOPkf1NhIamHcCCgGq64dgXadMO9ikJ0Zry9Z38FMpKJGrPWM2owFeHpeQjnf5DJd0AAXo
IZ4lPzqwN2fZA/rZ1APLAE8MbpIsGoOb8xe3bUNoQ3lh6LkggGs8Mm24+aLndYuAIyTryPG7mVSx
vNZw/ZYdeYVM2/XCBqCpwjTXzcu7FPLuoNOJT4ej1DEleZljCIrf6gpUgAEl40ShWB3663Sgnd7D
M80ZRmdc+qB6oa+jEqkyIL46ApMH2j0aXqVQ3DXMCNG+U08q3nGKpK/Zb+h4dps/UVwoOMRYamci
nSqTZ4E6/TVzeDCE/QgMuO6wIZdI1EGpfI3AtkJfw9sXh+sk85Azscf3vA79sUrzH7tKdu7S0Cyp
LBx5ZIHnrHj7TUTvQJ4i5rEV1If4tTO097tHxmMbRnob2DwCvqmmPI0Qs0VYCXvdXrF5xCf3oXQp
uC7QcdAt3iXGOLQZA0aPUyrj61nfHM74HO++WQv5AnlfEos/b9QBhbvWtX2FFBvEcSKEQ8oGKtMQ
Hi8oS2KtA6OtalG/phXjtu91cOE2EIVncoIDRztsLq29wxzP0lhvqi99NIddwpuoxunQvpx7rIN7
oSYFJpFLFSEnZpQHJKIWL04iNqfAbWJNauLy3tQPZ4e/3hvKngPJpqVXrpzAqUlx9H0StRCNJxMp
jtPURBDSb+nnu/PUPTI7Q76EucUEYTp/3LlIccg4ONWYbQy+eLbNAas53BY5RP9GpnGM2vzahEn3
kGYoMCSoDqW4ahRAexJ/MgBKn1ZgWX0NeNjwGZpL0hDRm4Q4xp35EWpjOI+2cFnU0LJ0MuxMBC1t
eytp1r0U9FwKQebRaZeGH8h4C8GKpn5J5QuBNU1HMDYXcRhKjxVDIatew7buoA4CHspwTENw6Jfn
+o0/nL+FdJI00+GI17chWa8jfj1pfxQpM3Hj9NlNWa7RdfsfCAGTe4KQUHVKbUyz8rE8wukx7WLy
KCMHDlSKMMjav0N0McLjyK556D6TUcIydRfBfEc9fOiliS5jEj1lyVQUFQd/G0ll5ZRlhKm/whMD
MmPfgV7W9YIrDSIIESSovXNGQOO6WxAefQQVFD3lgvEuFxKzM1XhVfRuTlFNtSXCYAROSl3fmRUA
agLLAo4yfTFnv+LPjvfkHnaT2OWzCRLZLEC93XOd2E1sHslZ6JLr7Gz+fyhMUjXTOmYLh/MfAJnp
K8BrA3X9puI2LmRFj+dGTMlsFP9AeyaZ8mElB2ff52lZOslcjGemVj2dNZiZtY6i+9dug4jGAZdY
+PyjfTc4quEu9ZYBS+2EIIfWg5n+r5OAKis11CBOy/OrBwphxGdfsFA5wR4uFFlXRHrDkkoyf6p/
L9MfjWBtjweYzaH+wmQJ+CFqDkq/8UVpNuPLTh1+CcAb0NimIkdzRP5KbzbfHu4gMwcjRrTYGiXm
rG1MQmu/A+SGmeuzGoFW05WYKGkSOZDuTJcriCCd+Pj8q9HwbwafF+ABiSbNtHooR/uKw7HB/b5H
c4HClhJSw94Vcx64Y09pVwNTrTUYAMaFjMcgua/BhD85y86OfsaSU8n7SP/q5hw8bG+dHDjVj9fP
0znJrISvZ8jbAjPUdIJ3S12wf+VELhRhaIaCzM8ZyVEHlxVcrhXDYY3FmQKtEbDIrjxKhhQjoNG9
f7kdBcJ1TlGOjvcf/3YZ82OT2MvKMVtkI1DsDUM3OWHZny6cakRb1cUq/FjrriJO452vQbH9k5c0
CbOre5Ow6niIJsw7opztaesg9l9omSjsQNcwWTT5io6DckAXlzL0HluaEU0WKQOSNiV9E8hN6ksf
A5wiYeIdj2YijjuZmSjLFKmxcwDkocVYWmjdlhm7PptXQOAXRa5k3m7k/jPTO31BUtZkRTML3ssG
TDO0Szt+UYK0rbce31kJ5SDm/FWh8BF/tu/9XJGt/gvbtOeiKpKfe/OfYuNrNaR7/c71j17iHsty
EkuPJlE6iP+RTfEon/+145oJUHgZuiaVbOAGlUDUCn9JKGPbidvQF61+OUEv7BPiqYWIuX2KLOYk
gzFOl+pEJbpFQ7y2U2kVCUTiU4VFn46v+ZoWsGHX5M6xI74GQG8JebGBxzrKIpQiX0vUF55HVTPm
mU/yJ+CwbPpVfePeJFWWww5S8ysKNoU9yeDbN1G9/pf0jpyT9asw/5GGoWmhr/uJX3jYVFyGVMT7
wsiiSuXAFT/Odvl8NvaL8kK3GvJCl1do9CAU8gMF4+eFGXyAzt5uLQ6r1r+Ds8mcOQokhSvu/MQT
th4hlFxwuC6Z06l2rDiW5nbPCiD8Wn7uQEpgcgz0+zy0nEqgEH4KQKlTOV7fHOk5vjuXFLQFkCFq
6WNpSkbM4s3bHRMFAQRBtBcs6fZ6r9Fa+QQBW1JH4Icp/vQyJyCxZg4S9BATb6uoZNQaO9OEqNx5
pgyCp4bvlzHy568WfzPEJxq2mXPKEw9vEFQHRvei8HRYKOLTgsKBKHyJOFzQQCZ9cNyLhBfADKXj
TN7/bTLYxyWcu8Czau6vfu5WtdhS3l9cc4t9C/dINq9Gw0rFj1r4sYSJ8i11HDkQtJhWnqPUGxJH
NpTu0kiKyd+awLNIhSYXmRijz5HFs5sHLgTdoL+8q8oqNSEGPG+snqFY8lfb//PVN4HS4ae0dOwI
CFZ7Iu8Z9aaC44RjplpAMH3NQ+71WGBfYTEWQDzOQ/8czj3gJm5LUVvQknzycVVOqX4gDFxwL37C
/hRUg7Bnl9LIB9Gekl4SlkkHj3g5T0NfMJYMccedHyMwTVB+RFQX3SY7b7IcTCD9Upt51PF3cH/+
Svm+pg1yuEhQF3aXT4m3IaJbV9btAJgl5CI8rfJyDjaKDrKYhVKcm4+msycirsAxRzjnTWX/PNe+
wDMK6uotT8IBvVGgkHo89DIilVnV67xXTWkZt0qv/MuENT9e0yqlAg7fD7I0XZulFLPf9dPI+3b+
QQBKgDCZmDt6TedPaou+ebQva6OgCKMy9dlzmy3fDQ5ZapM1t7qZiNKDn5BmyOvhihMA2Xlmhoks
+ozQIhbOp//E0/hOjc+VH01IkWVoxWPnMwY2izK3MQfScssZlzS3yWBMGP636WcOe688jZ5kixL/
F6V7tUaCkE6IGYvCHEfElYZ3gauyIQfXIsgbY665y8R4byU3F6RuCmEXPAl6lJRifhcG1EdgA7uz
JdsU/pS1uCA3sA+TlwBo8r7Rawaf2Bbfqe4kP/RWgZcFqNdxoNtFGY5tj5Gw8U4CHWed8IfLNRzt
RjL14AtyO39p7bjZYnZbjLEAn7vtEA5gObaKx8ozvG4Dd9wk6xaNu6vNq0iC9g3FwSjL9gx09qVL
lF9/q7ojUBV6QvVb/nqHX4BPTA7r2vkzHeJKStmNQuHuXAtJA9286+yB9nI3gbrAlTNlNh1RB51w
zvg0VaRKbZLVD7EefXsfecqwa+GZc8OCgYlPuAerRxR4J9cwK7efeTOu9UFtW36KRosJSxLP72kh
MXLB0vTWLQGsXK6xjdn2hv0WWbDcWKO5bGNwiVIkCXCsWD+jCBBaQI/neklcNuFF0qe3XSh5gfjZ
KWh0bc27aYM11Kjk0Pasqu3+LbHMGUYhEEMRl7vYbSKqecyf3i/9cW7jSX7m4n2RfrFeGaMRyPZq
GzKet/2gf4rCqQ+S3h9LWPkgiHr4c9dkjqBRdIl3UXiUsm0PzvWDRqjXBjTf3MPZchgjnoY/rVh2
cHCRSR5s2nZuvkKULEHV5trk3vBBq8YRKS9bff6wmaIQwSPcvq7MiQRfQBmmH5qqXnqMf7oTOZO1
s2xH53xB9UxS6U+N5c2GVf2MX93/tsuJ/t/8oKEwXkBYiGry6MevtruNvo1Dh7EAdGBOugnQRHy2
ymOwMHZgY8IRe2OYeu+mvqd6QN2j38BBaDToadG0lhyvCxvb7bd0Ep202cAqfo9FwBU4HO0FerGS
sJKRKErHZBpf944/h0oUFmPW+xEe8Jlgrn4lhWutXAvQAooY65duMHtEN8st9C32hkqemmQtPGPz
mYmg0vCSE65QhlG6xJxBeP0JrTbDrPT/QSoxtqK/VxVc1vTFdBKmcILCyfNdg/waoSfM0GFtLHVX
466rgbbd+cmSwniqoTC+hI+qRn/fU4M584z4qGR8hoNaw0hsgJaW21jPlBQT7qjfi8jFvPmxTrGd
OY1T1imOM3zqZXOmVrFp2rkgL4P+5Afg5z/8chGSuoL5uzsNIY4I8TZGZDCcDLUAjZ/c8L8TtZL4
fttWEdgS49U53hWZhX5kevk8pwFCVBgx5oS6DnXUX3eKsj4Z1RAy0lvfL+ZxgRkbEAfAi5WXjhy2
s5OWoPV28yD4u3Z3wLyZvRFvm/8RM/A/KdcJrAldiU8sVGukwFO8yNDggjMgGJksG+XHUjn2jTT5
hXVGdk9hWhdzAHI+Tjo6F6RQy9OPTfcMlzGlONJl4HjBUC/1cSNEZIFfHqtQeZTZbLqzl9rDVGHQ
SLWlAWYDj8kfO+BS/GfdEFxuCA38uVjH1zwxUWdvXvre9bGp3OKf8ApWvaKHk/akYcN6hvYiorCT
Of1KE8XEat5XKX7IBmDpvAPVkmgcNH10jr1vbkGI1vvT2a85pi4hU/pyu/pii+UIBNsLQeFK3gD9
SznyV67LqEwgWgUmbeG1/uPypdrGbOEMrLiGpg+q81/3POyd3gSHxxh93nqxvSat57GBkvGU0tyE
AqGnGNaf2u9oisIjWYwSr2hLgRmfqfmHo9UZb6+qWHIYFuOdfTz11eHJbwP2DjxYXqdV5W3R8rPP
dCZuREWWv22DShpwyRleqD1S+MGKhHs856eQzSXLC7NVYiSgrkqPwrQv1aeeJVvshvKOGUIVyfsO
snBZJDzYkOjCU9EL6bcvR8R4XRlueeBccczB1RA+WM+xGIrW8iWVykUGEHV0W4nM/FAkMaUIE2M9
6AN0Q9+fQzZ7Fe/rDzNxf9Cq6FCclR4VoMrDyVhK65RtzXEjU6b7Ab1itO2yQ1q4fy01hofHKdJG
KwmRLdEHP84YDcW40/Rqz/Td90r47meVScCMujet9WO4/DRxReQ/Q2B3Reab7kFpVpSvtEg42tcc
Qme2hW70xBJo2MUtd+58a64MRWqbQ9R5Jtd5xjUjDI9rempCh0jnF53sOphGJ5AgYOJLCtRQLyrb
EF7MYnlv1TcJ2P6O2NKEm2TsQun7IVOQibez13/KZA/O+v2wSnwV5vG2YU10L8ZHa4F4qzehkKO2
dVvKafjk7s+ZmtT7LwVJZHLGlXqeFhMR0o9Y3cNEvb7uZQmoOfVaJDtH72hyOC/TBgnXPJQAQz/z
hz+QkVYTibQeKavcuEk/CLRE6ZaI0137PyctuVnagAnC9Y0W1HlyYVUIw6R0XR7zGhhY5vp5UvPP
PV3YUdzJ0TAOWxNFGquKffXWUuvu/dsrHeptd1yjBin16N0kQrGEk+jZ5LBIxawR6BSVNFMWpRTX
tyg+5pDS6ydH7g9B7dUJuYnRSKvpD7y2bmPOO+ywn5/e6qdtq2o9d8imak9ndIXmPtYxLbJMSUn3
KRF76Byz1tLzr4/oCqmWZHRzNdeUC6mVNJcHsYNIFMh7MKIFxe17biIeUapBXswsGSr8TWxheGHM
NQ7fwV3ogQAc6k1w+gMglnu1tCpcxMuveWjzjcW9r9RO8fTa5Tc2nKIhKxmWVQt8fsFCIcNOEs6g
stBDy3zDsx9qZFmHRl6wy0c3FHdAmRtAh0nG9uxXYwMBEoWTY55Qp/iVVCgpvV4PI/atsHB8AMau
n/FgnLQPcWMuRJmJ0p53tEKi09YYfHVkqRczcJmy+8p6IeJ4VaLagtf+NZiX1KIuAPbUb2BIgDyW
dFdsWKKOH4rjt97Bh3PP4Zxa4Jx2tacIy6ksXwOH/bzLQzFs+wMIs2tqvrIITkzBF/7H+fvanMrX
4X/8t9mvMLpvQcbJDe0ztfh3hHtVWtmWKSa0mhLybXHUFsP1R8oU6cOZjRCgGpCJolg3Q1dUIBdh
LWjJSBimOFm0vfQFxEhgEegTJ1HGi7wg6B3bMw66ufRDRzRSeBhLxA7ZFQt4ZJqlyxwVbATGSmex
9uf0G+7LkUepq1s/6XjukgCFvdLX8CSz18jD3rZEPTTkjotpow3ypNCLJl/zv1wzrfkzTWdVkn/G
DnigHTKbDbKi5QBAQ9LupREHCJqj7sPKYCsQtQph5LRB+HOeQJ35oQRXIOIf148V8mZkcQyk/ZMp
CyGCGYv/Qx9SLFJCSyd8UOMK9QtGl5xOMqeHWvl6YWgcXaB1cSYFtH8YyjqclBgQvHDytEQ8Ukbt
AUsRgxmFhwlg8Alr2XetDt3yc17Ihqy1SBUZyRs4kcT7xcWxwvg9hHAyUdK31v3Y2mri4znURHgS
Wt0HfjlN8xSHuFdoaj4DQw/urdBZa+uE2L3SzVt7b+PejLRXS6eCpUwEPvDajZphAtfBZCnuCSmf
E2Iv1GmsWVaux4nXhNBuP2xuBSlhWKUK7bgTPs1q5lUrmzqWkH25Pxp1Hr4gUvXeQm5gH5/2dYaK
8L6mGOp4UKEe++L3SJ7EoMGzUDAuEThe0GTAmhI2k7sHjskhenzpUDN1v0eOIePLzBwGgebLx2nn
k+tEhKcw4wDW9/0Dthw+DLTpFZey7cG/5jocAVRCsQkScf/V5fv5jcKdGhuCt4+mipv7+U4nn1b8
T+DBpWdREyx+A7VDzb4umfi0aa5qiQoNbG9vMBYb7SOHl+fH49JrtP0SbV7/AY6c/3BglK5o7Y7/
RDk4L1qh7hUDCsGYFrtLD+blcT4dCPoN+TtvaP0GjJxDCFBYzlk4eIBr1PFjMFwXl9Czwb+r6gcP
HB/Ay36rDfUWfBQnLZ1lrqhBBdyd+f9EFxU4FJcjT3Sz0omicnB+n3ZN066HGSYdFE8KcJoJMhei
mk86pmf7pI0aCHauPBfNZVNJtlnNRmsUXZs9sTLa3M5KBIYa7/ZbEF/Hi2iGqMQhQTRlVinhR3cx
puuyL7R0/n2h6TKsxIe2zZn/XZuAWIjYodOhQsMl8Fvr1ywcPuws1pt+7IEB9JNu85LgOrUbY1Bo
Hpd2ERMS2N/QEALWAbMnOkzhqFpdIx36enjfyhS8S/TxywVPgeeUxQ//wxuBBq7/CR7r+Tvelmyw
Mm/Df9eVNFvCsY8a0ypvygPlOGwaPNNlX/hb21jx3OxNHb19rviTgbdVWmDgwpqCm1je0WHpb/+g
pmyYkYlc56HaYkqk0Sy5c3YevXR+8W7cB1On+KBRB1l3Os9OLeseK2q2sddKWkdkeBCi+qVsLbIw
KLnq7J3Nh/1XCNgjsMWzcwMy9PtKN4iXcXLRpkTRPL1YqYEfXbYbndOoIkPB5lEOykEMuwY4Ju4n
LzaW87igg5a5qLI+0MTqawLsWzyhjmJgWbHUJlh+4wY622cW1d2v30cSKU5gGq1nBNzv3G7QRIQ1
7lr5YhbM3M+pyMH0pZq4UaxhhHuEvAy+VMF6WiZTH6iM/TZloDzVY3jEYGSSuTIFD+0wW63ZCKON
Yyc2PJ9YrbIcq4HALrK5NydhYqmiPlIywC7hxL2Dg//rNm1VIghgxi0wH16XLKXX/17dsg1JxLMn
2gFkDh2xJvzdi/yiTCa7Aky5yj/DSPbVKaFe4/hHQyIPfrYTtKH4nQNZ1TbEUsnfSowFtFHIXQGz
j8hxaJZx7ce/vMNXDWT2mPFRzKkIEz8yDqckjbCkZ7gxzRpnxMzyXYKCDH7IE5zY7v3Sv5AofIja
+0fA7I9XDqQjLR8q7OW7QODR396D4bdZKcIMiMLG88p42K0pKUsFS2FVkeq28VWSwrmnJIZDfG9Z
W38ZJjF3o7z1b/Ut1v0QEsmalZas1/VaetNAu6jeCpnvvCoxCeltBPskCWcGc0gBPvfNcMq2hQVS
CvQIdGT86bLq6qiB3Jf6+655O1UGiEnbRB/buG5OdoB2tK1BkZla8KKa45f94Bn+Nh46UB7p3S1s
GW7gQR6hLMnHANm8n4Xb7DMPb8tcl3vTlFrBw5EoHT3ppLaQciLyoG1BqJZXugQnqSs7MlQCKbs0
THiEf7WglNpCFOuOQkqXDIrLb2lGI6r0uTRIQtrdSXNMIMFZ4bJM8yyZErSLegyHOp3hNva/VT6S
C+xCdeIArbn8c5yTxKVnXOdtp4ZBuRjNfhdPpxKni5ZbTwfF/WZ69+GKGq5MNbawQeDZ/DUo1+dL
a4tBH+0f8RJyIYiX/hJi1VTsqT9rs7yiwNU9gIIQChHy1u9wbPR8HpZz/yHo9RYlO2exAo8kzZMa
3hFPahSa1OkJTXo73iiJf3CM37KfJyeU6R8k71/nnYqB6bQhUFvWqFdr6BDdpXZF4bVhke5ssH91
1hK64/cxoy7SKR64UF/9dK5FayNdQ2fdV0mRXYKOEguhjm1yVOFeVWpdVtkEqWeZJ2dui4SeCvLy
fk3VflLrsDZCy2nFol+EN81lLDksk6jbifscOGvVeixLaNDDAZ/2pBwkRkM3fYDZcwYBFZVmo0DJ
ST8WZ+P0YS5Im6fZ1mYetnimGkzvJlOHgPSBRorYpP+t0bH9fkSQ4RMQk9akJegn72I5vv9bmF3m
x2g1bL35Q5l+ZLIzEw34phEDtK5qRJwvAvGyMp72/6JjxsV5DWLIgQy0ug+AaTj2ZYnYe5pTFMP2
a0ZJxnS4ENS5kiQhPa43wtfIQ0J6E5IBMcQ566/Ghf/BP2F915LQXbOTg6aaX5D935G8IEKO0DUr
nEae9uZoALi5IuJ6ZHvLCO6guCBdowd00oObmTtsw1DtMdSjFu2A4g6Q3Qu/Igp8yhCoOSPpXHDY
4qEIuTmifriy++bKJT9sZD7+V6HBM4A88m77bU8IOAnu/INrXikmIhe3zUAopXotzDamCe33orsy
2xkGYTXe8u5JLEec6Z67vBxXCG2D5n9k17J2qqkcB6xIgT7OZPybFXNH2DK7+6j7K3uhDlAvfP1a
HQLFlVjLThOeLeHtfZQul+BQi/0vSZImRSborvOjC/7xZ/vJsyzNd/ZHBA+t1vI9wLMFSRviC+On
EtbVc30VDsEA95lLO2djGgz5RWLeR7ZTWGdhQ088FJMXSRKzir6FJhQBV5XYt0rx/r0eSPB0k2j8
hdnuxjCICkXDmgm2El/+3JOS7Ez8/MlJnYRklda7rBsDXnc9/D/Vq919raAivS2kKfZ2xuF5ElbX
A66yCHYdquDFZxSExEiStTB+sPAOpD0NPK+jM1UJYI4VKbELOuSGlyjbolXYgfizHZbCmIszbAWI
7rwPocUQppbKgO3+6+4AIQoDA4ZA2zeo7qrAno8jMOnucb0UlwQWG1waYmiK8nlp+W2NH1ZTCAWP
mcAY4oOqDQusrSwZSFCPMtWkgklscbW0xdkHh7D62LKH0sXkJN1jTQoa3X03ZTRaAXHl8JZasFe2
QMWXWSpz121HvGmw6tY7eO9LNQkDUo0EcyIMCNUDXD2Xjcs2LYF1NxAasHLjBHce4X6uXZ10I59u
yidnrAV46HLdHe8QbunEv0spyxFAeDuBFDzgRqgH2YgX+Bwb+CJaILGtjql6SRJQCwCooOhh4cfY
Jlrc2C6IS0oqMkb0z6J//BvNzoQWKo8K7e3KdLZIeJjtjjkhsNR1zE7l0u3N/csDaaiyzafD+AIR
acAs4O5YDqmTIA9S/5IyBRF5OC6I3LGXtb6liv2mBnnGqyo5T0Ot30DUWuep1HtX+pN8pW/7RGml
Hs8iKWQ2B/g0xOYaeMUre337LAsl/MUE0h8hfb6IfkscS3FzkbL6goKgQtPREJkN9bYHxx/eIget
S9lbg+fwEshm5mimkQyoLrv2Vh2gQ589FFGp5JHUm2c14RD5lAJ2URlJ6vFpsofWy7ofFUhm2Mv+
6shyjcqbdpioW6Bwf7eVZzb28TC9Vi07Npq9SLsq0Ul7a74mDw8EeErh4z2DT0WWDsrRAyuy5vAD
AKkvIByb4I4N5m8IhkXIFVQ3Qhy1wjHFYTjk49m+rlmFtrlxL0a0XOTaAW+OYe1DJJaJSDe7wztY
4/cREqzU9yffWpNOSaSPXee2HIUqyWqUTwMNGav0eYdGJ8uGeGyYEQDkU1BaE7RoUU0LGefiqTrC
s+Yy12Bv2Ftav63NjOd4dBsU9vsO28le4SuWxn3mz8084wk7ZuioitmO9ZHphi3ofCLWhpoGH52Y
OKxCewt9gtUa0OiylYVjDDBeUF6mfTUKXIsURUT8oYWkmUZVYToZReLt4heTiaQQDoaihkkdJ/Uv
nSqef8Pkk7cpNYAbutwPK80awSWwQLilG0WnP/BUls6LMJ5vq8Cqbsm/bTsMV3rxLkAB9B6Y5tLG
Qfub9vjgwn7sgApgFIxtKaYWgFZav8yeVxaWaOexjD92sGQDFVMWT8xiwm7MkJcdTUDlArnfMuoA
OHQrV1b/SDGWRvzIlHJNYt50GDOEwfUKDB7nQBLXeIZkpr2Cnn35u/PS82fnOEYvTGCwQLaaAr8a
yx+gbRjgUDcFlYo34DlxEODe2CTujjI0bSo/dJIYvfJABwMixueYsdlAHQ0wwauyyz3CH4fHXr0n
q45O9wbs0ofDXLW1Pen4JA4rDSDW1KZH8Rusy0XuTVSiQ7c022/vfBm6wQxxfpuAOeeiD7tU+IRZ
jfsbZJeMX+67MeqaZH9TxNCyy/Z73BdoUU/pXQNraFj+EazB7IKh6aK5mfkyHSZy5FwkzGaRTCj/
2wJCymuaByxNsKTQBHHizX9sNzSxzO2k8Sh6r/qfxyU/KB7GpAIZpKpYHuSOMbAC8uC0P8llohaJ
r03sa3qjh7B/F/5XaWT7c3VsmMXs1BsnIGfGYLq6vCGNLpJ98vVNHvLlM1gya0u4mThrUTxQ5U6R
dd5WTpe5zpP7B8w2R3ZC8bJOsoAT9cxTSfB8MvkA3B/1eQTS3jLU4/xs/DgYoEzJ2Ry9PHM2KJtS
q830FcKL7Ex0LU5/sVEEjBAvaYaestry//+q655Oo3n682UapIcg3RpCXoGEbo+CmG88tEBHAxwY
qWW009MiRN/KWE9MF+vgBqymF6FKq+ryM9Z4aOpTLmZvECV8tPdaWXHwtKRrov9FIQLNVkiwsRvH
E9sAd90Onh4wSwyQ4FOUEAosm1SPdJ6TrXUN++7NB14WuS9Djviqjiow5Mxqbi485YwwhLWfg7mL
SuNikvS5t2AfkNuSiyiAbq3puj8Vhee/OLxrSQozGncWOAYzSyqTdEb2GyMfYsZyHx6qhPVLtK41
t7Ep4UbNnLhNIWybGaot3z1LjPv9unxU3PiNji43fhgJc3H3P8V5sAiBLeVLreCHIABMXINiTi4T
q9G6E/loOVbgvwkjGg6lv4F9CfYdHkxzoEqBBVw0YsKYzDd2Qui76NKarUUO6B7HynQHKMtdAE+J
vWFzKrzaKEpCN1q6wvixh2cgzRfjiC1sVvmccberMYoWhIW8f0hpFAHo/32eIwWyUzwfGQJd7esH
Wqq0Sp9ywq3G6FHit9cdo1LisBykguUyWjKC6N12PtoE6Om93vxDQIJjkK1uhiljJAKV8tek+jS/
mQVvVNTF2fIdXQLN+gb2vHNde/OYwD/NPE/PStBgKQwIR2hCzcAfBia8v590nBPhzpyUDPQ8rV4d
wsq0o2+gxuw76mX8sBVqOLjykBsZrG4ZktuEazfxqzL81xiN9v0BXNGNQ2oZpDWtzmW02WE+tbUv
Qvb18qospWo0itv0u6t0v7AwwKZDugB6DDLHbuvORGt/cKss2q0MFxk5VqqbGJENQMqXpfvSD1i/
kQ3pCWusFQrKj+qp+Nhzct22mj0AlSJZDBwb+JHeJek5WQZz9JDcYp55aWGlAa3KkWGCuAneSI0c
koDzpDMQEzr0RjCNdZFcMQD3O8EXvBsWSgmRLCKTaJhc4u8xXl0WvztTwwBzxQgAA9wgm9gbhptD
QEqP1PZYvmZO3ScAFZn8Yp2aMJxBd0O4XGY9aMxvr7AG3aihaulOFhPU7oDSWQaRdhFnueH3/RjC
UWqz9iTdMCSwkc4mbOVxUS7Xax5m6e6H/+6KlnfV1yKO3Z+fgID2AZVVDbFIZojeO1/Pp5/Ao63C
h/Ze9FoDxYZHiH+ITICHlxjzyetq4OM9nf5UvJehiC9OyjBvfvbid5R0tnsPCetTSESUx0pIPTTY
5FuloFdtKPiVOkj71vgBMC7Afu4AR5LLNHNTTk3pxE8aN5tcW5+CaBaNoLpe+2c7d7rXTCudXf8w
W8MgyDQxWpwQUWQ80ELkSHrRSwsQS16fkjs6AHzERGX3+U7D8K/Nhm+5OSof7ZiEjcXsQ9mx2Qbo
+XCnSDk/eOWTH/r6h5hJyVLZo3mvb6tXOJVfu0cuLdCUlvHDTiAhvmBtfYaVmsJ87tYl/CJE6o0v
EQQHptGTKlzReMYlX13f92owVSEy7PcpKZHpCQpMm+f05Ev+Mn8hT2AmzrFHCXJKNffcUevHymgt
JXOArwct81DCiPAWpGyWlWKjGTnJgMlC4pSnq+0fitHl3BCNkJiUfMivQp7pa8I7hE6YiDWVLEDc
i5Hom+uZFhsyYlj6hQ24UvuV9oalAKBOMeCodsZnrInijuFXfGqh9pr9GEuchh3D8se7QwbUOn3b
iq7DquVtmegBDmOpUpddqGF7cdJYjAyh9v3oV5vH4hqOQFA1/r4/EkhJBmA9GtiVnuo5n/an0bhf
1/9qXD8BMuqIwwlZP7XVUXyE4EughaK8yu3QLPjE0AFUvOf4tm6ZBG3dFJ4jhdoS5x/c7cqtsOCQ
n6/kd510O4xFGCa63+1ZEC5zDhCIiX7XsQB0HvjLA8h0zgCfSev1viSCAJGFPSIrq2+p9i/cuvpP
3HMobYXmu73RQjTWiX/34p1HJhzHgXe3wsSMEWnRj+euII8lmFTsUl1xTZeCKow1wmGLla4We7KE
udJF3v6HIXhCe8lfT7dwmubj6nCpBvymJogZFOTl1+o1uEDETwQbIk3IKGqJ06P3LMGTIjTnRJyQ
nepFUcXZNoDrqGF1sXPnICMaiJ6u8wKU3Zrgb0pcC8Mecgz3EQNiJj7k22IWUqRyZA34ZccnybS0
TGer9GP3RJ52g8wR9S5NRrVJcYYWj6Bn4mKBdPu8luzJ9Bh9ftJFc7/bQrZWdOoIsbMmxlLdy2+1
GWx3QEwJOxbl+soO16sKkM2OSo6VfIa+urESGq3Efu2m/dZFkfy6XE/fY0KbV1eio1WN82tRHYvw
/SpJ/QqKIfL/g3b7OYeYbIFF6TbEsUFu/6YqHb01GiC3urTXRayVuZqcTTg+3qMGfTUOAeAk5MFG
3+gzxE79KD57XQ42Mdk1pS8ThoIxRzz4YqKed3rXILC7JyOLbB2ZbFux7WO8z2r4AXrt36+0qdXd
VM2gbvmq9OaS60rlmXN/24Bvuq2o+GHnpg6l6AjOZKM8x+FEBqtH8SVUtvmAetp/wwcQGPNt/A8L
wNwtN0Uc7sAzba9GJfGDyFpkQhKRa1zFQFRS3zi9O1IoqrsYC4enWg3a8jE5kArxixK6FVyhY6bg
Bm7xzb78dxgSTyPw3br2vV76krDMthBzh7l7tiot0BUw8sRJ1F0hm/D/nxFAtCyc4nKrrRgWMeUG
1+FqbD//Rtzbo5y16sKXUJ1LvE87L/GkpblZoQkKyNc1oOYqjx7y5Qrz+8ObYxiBU1Xzb+JwxtGO
LTXg5rjHn9n3TUT71v9DF7VVW2itSgacUH7En/L0dtHZZoCU/A0APGAB3bf4wOynaThedNqQzhfs
CUU+ERX1fVyXbdqIs7IR+I+EBRvu5TV1mpguHFEciIwhE+TKskO6dRMetoLAsGAKtopg/YAG6ihG
IS+KuszJOqFjLbr8T6gtrrrIfJSWoro84j0+CisLy/MCc7O2+1QN/OwAD1Pc70nkcnycJDVzMnGx
cWfoFrz4XIP8oRu/yOSIYKiQH+bcHmYTJ3oaXfzyw5J3aWI4+evejpDxyvIl6yZ6UKIfN7V5BT2K
emSg8iDNY6M/KuERPPef0IqxdvYratPVADD2FywMFDgud+YiDuQ6CiplTYTwGeRCdAQdhSGG0Cgi
Ui4A0noe30jiZf33e8CjDQO4BjO/sJAJfhNrppVeXyFJxBjgnAI3v4/Su8MtcN108ZYvxrx2/OO6
2txuhL4WFOXq6fGPsr1xMfptue0C0dy08NQwAuR9csxBf5qfyD1U2KfAcEWxM28UhIt23JrTQvUz
j6tayyyQVfEuunByhnfJx+zAoMT3tD8uiGsgy3xzEwKJADHVKDTXnHteSBi8AlVSQEaQXDC/lOHg
7HJpODcGGK/jcWIdITUENnOaC/VGEH0R3qtaLpvCqIV6FKTNs8AFFRQ19XDxovI8Fg3PUW3wNYNF
Oj/FEOcQ/Yy2ITurEBWeX5oV7TH/f8yOlX4Su1c1d+IsgbhDjEZVOqCFrNDATEbAHQoPfLPDXaWI
02V7CXgH2yBKyYntRvNV2bL0nhwJ0cgbm+WJPRedAodU4x+Leie9QJYjSkO00G62b+hTXcZg0wHK
h5FB3hLzfSxqmjGVvLXQ7TAeBKhhdq9u9Vn1qZjVpFTRQllQ2foGZt3dShX/g0Xi1OUUZiLOTNt6
zi87AvDJaxSiBokmEykKrVwWx/MV+oBchLb4Yb/F2Pb5d0Z50CkpZpm9maPk1dRB/KHD/SD/7jeS
4GN6LJ5s/QlYdiTLa1YdWBnhVQj1m07fb/Oq+rTwEH8WNtEbIZR2VVVuDnml0+aoQgDqesz3cYNK
21WWTqb2BMbSy73O7qgGePYJQhfwpgEZJPZ9VV7gCdMHTjJq4ksNMbc5Cs5clqrx5AQAojffwXcO
OVBLYSh8Fj8jt0QDMZ4HxAxo1DlRkoN+5w9sJZt/0Tj9yyjhNt61JC7Ce+hoUJ5F07GrjKz4KtGP
5nLcgpJ/L9lzHoGQbQdncFuuETnfDDtZJQgWPEZ3dAIbwtuOjcaUemCiMM17Qqi5NcPqnCa7iFJ7
B+7/mg71xEOjZQLOMEa5GZ3jvOp/jV0FYQpf5frOskc3PypLUCauDjxQlmhEF2S6ZIC/7KTBJkDU
/RMZF1Jvuzrd1co1EzS7zW0B1oih9Ujjo7KA1x4LS6uOCTH7KQGBbmwSGofVQ8Q9DGqwHfirofEe
txAQZ0ggBjfDuOmnkKNFOImJrDYX2ycECm1dw4llGcAn2DXBe0rpilQVHGrnh0OewDhVt8mxl0gy
D6lZG/EVnjmIFNORbNyckmFZM1bPT6Fp+F0AvM5I4h37UZRsWS0SkN9VrsKhT/Om3taqDPcjVufD
frLa8S2FecWw8o3cvobdLKLPCeJ018kvEnlD5SJFQO3+8dKUr9701b59x/HHupddiWMhM2Nyy+qe
brffeHn4W7kpjWjtrHBZPkZoi5qIqWccAu9ON8W6vcy9S9f0K/N5FFjOAuYVLcmtWej0bqsAoxK4
e/QwEDOElzReFhk4Auj80a7D2AoMH998FZdl8pyIG4JF3hOIs7X7L7fB8qUkFL0autgy6++IW9jM
ChWafpzKa79H9tf8y4j2kcn+BS6p9iqyLGJWN/5Ek7qgSg4vOsIkgq36FJDLW05GOOK6UGVLJOyZ
m7JrAdPd1i1hYknPmtBezuWZM3P2eTjGVnz8S0RWWQPs95LGrcURC4UX1q9xUomdTwU2g9jLyZUZ
yiGUKN2ns0zsnpgAtagqG0Bcnh6XFlfwy8Ca5tlRAEQD9iZUz0cTJ4m5nnoZMFBELI9ilC45dz5Y
Qka446Bu/w5yHj8UN1YEh05zub4WCiu5hz0x9/k/r41At+eTMSELzcpoifLmZvX5xyxW6U0LXBah
EZu1fI9OfGDr1AYF8NUp/drTTYIyi2s7FA4unamDesTE+5ehMkHSTXP2P7dzczFcyhpAwTbbsA/G
0IujDUOhXbbfBKwls4f7LEUcK9tdiczybVjrsYH4YoFbX/q27Ez5YVn/BLC+xAbiXXDUtS2xgG+2
jh1gnwNI0ktb7dNqpgZrExiHKo00mra1dn1Z5Up3FM4opL6ZqSrGWXFEczZP9Fs13ZbR1rDqxBQG
yx2l1ieM1aHprVn7GhOCc9Lfd58ZhWMH1okzIDDADUMByKD5aPCMe0S+KwEsOIJwASlFQBv/tcg8
UwvvH+cnWHk8x/4skgltcflPDhx1KY8O8Y9Y3dLBw61SWGayENfyYZB5qteHLWpIKBJx6UOSofbf
oZJoz1a6/dvMFDqhowbT07F9r+iU5RGSv7pS5236X4wk6INNF1qccoOo3URfDRMSIoMHZZY37zcQ
GwxfoIQx6/YaQO4r4KkLUk2Ycket+3SBBDYrrW0yXyae/0gUFC90g9EnXyLFPUhlUZMrbSZI+EXU
YlUIkbsOAIurL/BlfXP2MaPu9Ktz/6VU7a0Yz59c2VIJLMrQAotHF0d1PsWeyxnIdpiNJ1xMzz2u
cKLkzrkFm5lo/q2wa1pgUa/BFSVcWXUDAYPk4BjiBZpMc6a6tjHlORKuV18lesNaFkvMeal0VDVM
+5F4kPiwmprTgwi6oTjSPmWxKygE4y3ID40/E4Gnc/TFL0wWdQMdi9npFXLmcpXuULM8ADpTKu+l
92FpVdcykNPXH/daHO3CTvrOZogYV6G/Q9a5jB190MaSyqbEIboHyN6k+gjr3rUfkjTJtMpFNoyg
cjDK9f5RfMYUQe6hwQnI3y4dyP5hWHb+NbulvxCyHfPnZLIGqdHreLnY3ec7K0ERmFsxY8IRh8qX
aE0UEKvUI8pSTR0zRMSi7VL/gZc5A4zmpbodB7gE3oFyy+QaiJpRmxcxg5dunJg5gKSh/PEsuxmN
H7kRcy2YzncSAhturh3Przw3+jEpqOEj2L/hjkCC7sbBvQ9jyN5TqtKLazoHJcErLBvVBznElkCw
UxvpIf0JPpOzqywV+76mLaiH977L57wcIuruRyq7V8OQjzbkHehYXilP1PCTHSQHff+UcaxdcvSt
1vhAg44JYE7x4laJRGmLxN87Av4ouzJxBcM6byG5OW0EzJ3iCUG5vcUGxnO3GzEcqdjXkwCZmRCr
sIxYciBQCvjOmZ1otv3yRWIY/3V5rG0b64txV3ZwUeNlEdwc2Gi/HJZqpQ+/OX66BfjGTraO7xpd
vDwQNFM+ruJEI4PBjSeIUI2sR6dQyiyuvtahQIMOgnY+tyd08fMsLfrK9oDa7SqaDUbl9EWICdMh
LgKoLfsI1dEmVyC0RRZsBPR9GJS6t8jOR+LgrXV7/gpkLUZ/k4OJ/fetF1dtlCxED4cCxcQLAc2N
68VwbqFhxGfT2diM9yTD/7Sc5eXSdTPsRs9I5DM5g2cMkMHbs3Iv71xF6Xbv7NB2tSyDlBNHDey0
N99h1G2UsLsda+UT9LG81+PyS02ar0Nc9fPb4d3aaLLaL/SCIU12ZsVDCQSbn4P4Dp9XYxracgSh
rUuFDECnBNxK6Vmx02wM1kMNX/YKNSnrzBTLbfp89WKbopWseiIS5sJDIGe6NHaU0F/UQxA+3z6m
rWoBpymLOZ96I9pwXYEustEmTzh8QSWPB3xRj80HE5BWC2VgZt//KN4YcEbbyEUGfPljPxSQjbjw
FULacXFqaQO0ngPNGefRTCMdmGMwO5xp35ivtCNlf69C8CpFZdTfrKMuU2QeKNFKAWW46RXLrIcZ
oSCafcuIan/TH7bkZCTPn265PmaocvoHh8X0ZxncPEXP9QYgUehU/g862h7jc/S/caStmev+dMJx
wWZmL/9QIwZQ6bsosyBaRkXQnRydxQIfGUKIucP95PdEuT/7zQrZ95jFag8XafMoB96+GiOzjXRT
7jgQJKZf5K5m1i0ULj1QoZQgmguz52cQ+yC63kLVhIMbdyChgEcXaxsi1UfVZP/3aGpJG1n9+mhs
tX/WW6K9WIViB+8eYhwqyP5RxNKccNrMd9PqcIXNZozusz0HL0bgYnDmxjd8JtG2+2sxBgSs3gaG
f3ynRTXk74SzdXmO1BhV6Iz4ldADo1BkJYNwCcaxGyM2Z/NfFJHkEjq7+rMHmetHFUYC0Ak6KlXh
xeBJ3fsTN+mLYMv31sQStSPlXlUjXHBSiaKNmfL0HVXGG3d5JCkfjj/WPvWGyDBAiiD75Vcp5EHQ
w2Eo+shdCxA0EDzrhFPx/3pTGpP87Hv7RsJ3b9MHUqIletwDk6c7Ny6pLMKKRpxo3/SYEJCkFf5T
A/GQsuhJhuQOTgwk4/y7ATGxTjdgrjmqXdx8VFUcsic4jQnk9wndkbYkoVX1DWG2/BXuAYrqXm9w
cE/WAt7z/8PSSCnmzzm5p+imteOi0dCNiXYUqUGARUddzT8vQsBDm6fvdt7kpEABebkKw0Qq9sRZ
ni6oL9is1JHM8R5HdMCnWBpoEI2TOiOsIrHtjEtKEWLb5diWvZPbc35uBm3inyCMhguYDgPeFGIr
Yq4XmXMj3p4a/dGXHAwBacznyF6pvrPq3kZgDFVhoTzLItdEwYqfUc44aWKdLwF6JKD+jcrAFAWk
5cJrkHYUjHld/M9TzlIbZ3D2FwybA0bGu6Y961CTe+67QlGiYGB2UbEhRHDjuGPTx1dQMu1FVcyw
ahK9nb01hCPzf4hazPBotSEMiBzycEGovkIm0/7zuH39X9TAu+kSSgt7EfBlt5ij5//hIlLF7vff
9BKdMdnzeDIWFyZRAs/VT501GXEWN0Zw/Jhv49YarP6BUATdkJITeaqPJdbyGHkt802SJ9hUKdi7
lHVh6SZqWaTY1igmdmcyOG+wVz929f3aYeNi545BCfm6X0suxL6IOz2XPXW4esyBkQc4TZi+Zjpc
LkYnSdAHWwu35m96b3N8pOJo8vGkSfTNObbo8n0vgNXkuWV/bH1jAG8RhHA/OWHdtCozvWsnt+FF
GTSw5T8Lg2ykDYuNl1jGjnIFyVaWPLuhqoEAyyylcj5COUKhCsGlBYUB9HPavaZZKoBRUCZkXQYX
pV7SuMfObpTy4LkJDQv9u4qxtn2ei3NC+yCcSsr5/HHJ0E3Ms+t8Pfl4uZwW5pCuZpFXjobLUgNx
Rtn0ZDemoPAsWiSyFVXpOCKgmmQICkURxkeIOBBXr6+bhTZbX5Fi93U0fmpDYlQgwRBabtYZFDLP
rUSlAAlXplCLQLRs+ynV+swbPvQVC3ZBJeYv/6SiWHsKN9amaiD6z1PlG893e8GR4cZg3bb02u2I
uONRs48yoRPgbM5bUImzsaV8nY1yGT7BeBH1PMqcbBq4j5RCPFQlSV2xAh3frNjRntyqOCH27iDp
7W2bF100YfaLzGYYKG9zGbtbKFrO0E8rHlgilrrYaa8h4+/3VEqsQtRQ+JxvGq6Dg8gVPeR+WTzS
u9hUIiDAFFwuUdqBjElrLVpNmsCcwfvMynNUAmjBfaTK/0A+oAH7mZ6NVdcv4iXZfvd5WB2N9v/e
Fw94sOa3RX5baE9FKRMQAp+v+JdT5dn6ThFvjl4tdSzl5Jy8THE0gPwvBVAvAOUOzuXr/ZFvwWk8
msbDPxjwdZ1N9PSINEefSwlWJP8Dw1a7mMa8SoBObEseie4WD4IyIjNLEIkcO5AcM+Z7Qs31jYz6
miW1YClg3TsLD0idzJ0KqOiLyY3AMd4PmW0KsqemiE7l8QAaiJeDFhHDP2IIUHsh1DGxkTW26/lo
CFRG32UMtVjwptyOlAKomuPul5dgsLivZ4Jzk3LFBgeOWEuUR1PhqRSV4fSHwuJJt6DUpRddABlO
Zezfrn1/ZUb31KV0yrdLfKhdsSZwWiJlEGh+h91Po18GuWNlm+c05VL2QG0KLP5Q4yQH5MCDJjev
oeoRrpDmtlpEFKxbGSZVsvHHUZP/GbPgtUnWrvP8bIbLzy0hfDKxGeQKO8Xh2K2Bqd2i44fNL6ZL
jF96lJXiRARnpzN58jtnyUbJZvYVbOv44ARF/jEeNBoL5l63nxG390QYvkoJyYrbeB5u3U51nqlA
Wse2xVkDae4x8Qbs5fEZ8HiqSkZb/XZBoeAJNfjEtl0yo09uBlFpt+OE2PKQ+0bJtrk1GSIClQ00
vlVmINuBSZzA/qbL4ta62jIhieqy2Rv1OKwcEvE7MgzzyxaqrDe4cb+Z2FoKVFz1ABmEajjXkXN+
fCQaGw2M2UrEzN03i4zoicmYB7rfxypojYdhRj03Ct6iuDiQHovC9+ogScu/mam1qvqsMPDXQLPy
4dkDa7ZZYevMKHgbRPVbtLdL6SzZUzmMpmF+GTOB6zBZ6aUtm6xbV/ecwL89i0ugy4Ce8nuMOuPo
pqUPiRFF/po8wY382uzBGXZHj39lC5WzkKmbuYajJePjjT0RlYqIErMcoc8d/SpNi3yJ+Lp3Rw3s
BiUOUzk0TBL7DNl5PcMpt5aFde38uIT68/NTiWLC6//OBc+by0L98QS87yt9uRZiAHIhLiz6Gaph
NCY4q/3ERKxPK9HbvSpIO9p5PFy1Sp2f5G1XtSHc4UJfAM/CexwXirWEHIsDUyQr7j9pZXXZNBxY
nZIvKlUHeeXN+lT4w241SfetlfeqSh3+YrwGoOQZ07y3ZqW9YZGqOv1xet2ddKczjj/DCTr1NaoU
nBfoD+d6B1gaMFsrJntc1hm3EE9O+XOowsvLHRnMuaY30g8vrD3ekXxwwW+8f3CRXiQu5bLyYcOA
HUxrwjxR8iUbjqnAAKKS38pWtWVrigE5A2bpqgy1yc2Pp+BfO8VOwmd5dX5Sr12PD6SSNAI0fefq
cte2McfTDSTJtKC4LsPl0ODoJdgqnZq2O11XVassvHhfpZbs3qRk3m1VgH5iVHBqqs9KPNYnkjNp
9L3Wv0pUtU+wpGzOeg4pCUeo51yiOvEYsuREbo/z4xe4DivvHehIQrESbKRkhbUiPXpndXBax37+
Id0zk1olLUV3xQDNV2L6hKb+n6AXfp14mFMdIgDZ0tT6DGQz0QJ2SRlbDplHOmIthgIz2xkGS50O
li9q9XWxCkBXgwOjDX0ff/JoB9afvZoHE3D3IKI8dYx0ypJSGbYTPTahZZ3gWHhtE3iZUa3QgZA1
kxNKDSoDo0tq+FjQu9IJ4TZ9/dxsjBlvwXgDibmNLAnhKGopYQQ1mLo6xvbbJWYpObtnDy5mPWJR
yAuqv0XOlpKNE8qknM4SbKo9M9OrtvRQztyx7+nNuTiE8nkjZmvLAsPNflV8qHV0DOYpj+ZmcM8L
Ka3xN8w9PqIDdPzuQKldRX/LQF9PefX61AWz0nN3rgGHqhhTeYzj/58k3HNSTk6Tn2pIF3i+vPA0
vASJbwwteorWqXzVGbOq5RuGIsbivJA8SOK3GkZFlhqMFPD0qisUWcV7/AT92BaJYImNKNZ+mwxE
LXK3gSO31YcnH+aCJC6vfiBs0O3VX+zj/uM1brvMWTMkozO2R1uCMczAiUmEcJLlHkhrCkUp0q7N
u1k9WzIerLXEmnxH60gvvKWYT4Ybwgo83ru7h9wQzJf2Pz/NQ8rMThxVflP1FiW1aj0Hfri/6F51
FhY/4noCIPnEyB+rAOnIUKFXSurTBoHaTyviKtBQE2EyF7eOO1FUFw9asOnAmkrNx9jsaxbjYoKX
m7D9EyHkHIk06LywG9EJwjGGTdTIvBB7hhkVooT2bmaxKjemk/SmJdJEBQawWZgbgpUBIOjGQV9J
UQIGHr7M/WNAQFDBFG7j8I7mL4B1J8AUsjsS2gD5sLRvYhPPxVrOY/C+E91CNn63W9XML6I5bhCr
A/fcezR0tHILEZUx2MkHIZyQSmQ/r0XV3yCf/42t9huAMlrLTqIdf/6t3SNMgnhiKBu2N4DZakPu
x4s0ZSQZyAX0oG5YRTWGy+fQ3hhDdlN0NW2kFol2pDkMLIT9prSKgutQq/MLS67hsXAjBl5AFqhI
s6vpNw+UV6rTf7b4rbaIxRxkXj7CrSkBFYFPmfCivH6NFo71Thfg6k0M1i+H9WTmPhD47Z8HDicU
MPUGRscus4Rj9ZmsrIYxOTC4oHY/lR+2EFTx9io/5WkftZad0ja9/SjcN8p+oSlm98LJKkFJTZ2x
M27U/EEhgYoPncNIXPt0grSIMBAf76tB1MrqSXWBzpJ5H9h17yxD7xtdgR0GAFpFjf3UgF+mgcqH
XSHXfnD3Xv/z8xVOO37n+YVzWRmaJb9lL4iTWsCr3OcBhlfPlbsUo+ZNGLJdGEgcSjNxgY8qSI2N
3vpRP6jSgsbTQq+jCN+O3Y3T0SP5q4q1X47lE7YsqIlJMNftqO7PALxgTNIi7bI7OLrv7ej2U5Tt
fGREvrsl3bmZRtRkYJTdhQp891LQJ/2WuZhdBqoYyP3sUYg8CSyGdtEc/krTrlTPyHiqR8KyH7Lz
RpAthOSS2t+vxWzyt7N0TMRFnaoB33OiMMIwcmr2xGPGeR5dw0n1IVFAjMlQxD+yadhRTUMq2hHq
Wk0dyPCW0z2Uz7cyHeZBeXzb//2uk9EBjxVCQ/o4hEOWA2yvnEnnO8i9aSnAVhDt285fBsam0iOj
Atyp/kJtLRUMI/yUZpcAGSVah6BVoQzUmfNsEI6U09Rfo5mCMxZPoGCIWA3CUteyJfsS4/Cov6cX
0o79Pzv/TExyTnzDs310A3BSW608GpcTzTRrt8bn+lKsuhdBdopVoxV+sKw2QOuoPyd/NQ9+DVlY
SN+wgOjw0cH5D+QHdKsQiv8M7pAmTl2OLUvt8tj4arsFjNAfgNai8xJb9pog8hNjlml+5zK60Gi5
uLZ1ZnasvKFSAY2PIzPEqtXtUtJWXKzUBmFlkY6i/JPikrM0oD8To+G+LX96IfZfPDsLMVzzG5sX
Lwvl7q53xmt3ocNLtvywFMmt3dPEBKDa7ANfK7Dtqp5KHzlnxSVtbgwl/GZnDgk3SUE/WDIi5wnG
0e0VY1tBuoPbGp5Q1UPqlJPT1OkWQh52kAyx8VQZPPW0+bZZhfhq46TPI9oJzE5LQM/30IPhSMCH
A42RtghqMPqFdQI5Wi6xBTJ/xAgevKQulLulA7srctU3oKbpmC6hMct5BM46IL1cOQ6rsBiFAD9O
Hur3T/JZtiOQ9okJDUX09My/O/MwFfpP6ABgDB82u+Qhc+Wv9pGATJgv+eM+3fCPvUO+gDIe92+I
sNYnt2ffQ9iooOfLZykR7CyI68k+o4j0W249ySp+u35Z4UhCkzOkTegpWkuG86M0acZttXwHK5Kf
j3csJSkuRxYjhkFZE8UamswSZVEXgi5Zoqps6pbBsAvsRJyibTdzoSGubKg7ujAe2uVEbIJG4oRU
J+CpkgNQuaOXedYH+SWKeM6QuZ0FAwNt5kaE88iNUdNCXfOaZhpXkuOLsmq6c7jHFoY6/YRO9CZ+
mz29EeFYeuvvf4EaYgdVZmPC45TTVoaocsGDTR7Xhl30bIbdmMQZqXtuLnnZ2cSRhi2hz14ozoMS
1WBbC6L7rwk/jgN01crKDZc3b8voPi87QDqNzl130NopL6+Vm/fhZEUldcEQzcsw7HgiBZ3EGA9e
+3A6H7vqHQ8fKjH6B9J+DjZKY+jo0k1mhQCydspVGrzy9l8LzYU4NQggEVAmnXQkSDb6E15JuA6Z
MCms8xzeo1EaOQMzNoaSaWihzYsv1iKQzVXLhFJuhHGKP0YUXwF8ImqABzcz7f/uv0r80hK/m6nH
4VK/HF2TvuLSssi/Ksy4tef8hfhbdRnBShuzgR+Tc69PN+dvM2sIJl/N692rgaI+yqG3NXb+S0+W
M+vdwJCpQAGqCPqarfvi6RtqxQFYb7lRx7jsy6KqYB1iTes4E1F4vo7Y3kdp0nRZ8UxVnDHB16e4
GeiJsnrh1ZolaNK0QAj2tWSMPKAbI3SFwyLS/OO7k73RKZ/xsnLsflKqEdbjoYuPrsNl5+U9c8HT
O6llbbdOK7EKcjC1pXIMOe8AkjNOSifSOzRdy4FzM51NVRNLTl2im3a5BZB7N9BNDfBOPIaWLOxm
BpCc1XUbBXvNWr2qqzXCadwesYnM9xV+gPM0IhbBlAUnHFGMPVPp1W/sqd+V4hR5U66pQOHN2qHy
pMobGhNfO9k66rI+tm+o6IEGQtmjsSs6L+UMLcI9Ry511tWGzIVmo6aMWjAJAwGiJh3Lzqai/NQT
ySSDLkJ5gO45WxZErnU4z18YKUN1Rn9hinTDlrQnndpGBcH0bGpmW/AAnYgGWPzpCDflH33AgH33
nApQxCx3KQZBGnhJTHnhoyMxCRgYQsl4VWsoEcOpEWzpzplqIFDG85LHxxfgA9BRtHrL+QIMdUHD
8GdbjDkipNxq92Np9MaRF0FbbvmVkuLVyzM1NoRd+aMnqiLcXl0DyUCQyUvW8qt2bhUx3+5r4jbi
Jcf1p0+0NMdrfP6eIVEv+HpHNAhChqMguxQHqGsdy8wj2DJHMLxtWIcMrxCMLqJm8Bk/gxFhjqu3
v4tX4TMtu2pHLXsfWjFZhOYiRUxL98jtcSZzt+/8H2MM4fIyQIWPkKxehQr1IS60fIheLs/PA8hA
+YrkLQbH6K13q5lWScKq0k7gQHHAVh9bLoaq5LP2MRiLKQ/BNiC6QuYrPWkl3oxyRByJlT/V9VN2
IJzCFLXg+tEcn+fgHD8CyL9s7Oy+ct0w3UCXB8P6TQ9RFNh0tQkmQC5HoqXmLUSuAx+q3HFosnNH
SLYhuRsSVWgZ3nHQBfTlXSqhRaXHk1OMSwVJThRo7b60HHfIygc6AIuJWqLYXEPWdS6xpmxpI1UB
3yIo7I5d25zrJ64i04K0hrjhM/kRqwR0yKUwodYTWUgC1hneQWnydHuzOsSrvZBmBi1MHVfkBVmx
2Vlxqd6AmNvp6HjetxVxT77WgzGjBj2uyxkzOS9uxUrmfwMHMvdlM89etZ9BBZwN1jU1Ccp/R0Fc
qjrw8Li1ne276HZzOt4cpY+VFnBANJN9EX4qZwq5vldsYYxVYQExg/G/w5nn02Pf40PqUVFFdiPV
OZEoL2EMmfWEDMdChpkpbL/typSIbSDnR5iMfBHTf1+fBeWmlFgnuyyeJfApUeT9EjsoEfse7i/x
hRaEVk2HenMVQNBx9uwfgvMcAYK4CGZh7KNXIVmhfpLRcG8DxChNF1DbLPdEyOoc1TqpHBNhGVqX
HsraWiE6cc18DME3KHRGrSsT8wlD8J6IcSvA7W8ngpTNLQvZx8F+D12Wg45hvfYQ5tJmTeCLiY7R
+Q/4qfEdLETRAsxtE/Ygh5w0I7GrUSczzBspOPHFQdgExSYkBPDIApDXDaPInYSShCsXFFmJAr2v
gS38+IUgmK1Sguy3b2FFvP7ViE5bTUFhric+dTP6SjibQZxhewKNBwftp/8v73s6ITWhXVSwkQNW
V8o9a2OlJOmEmJqfDEnPZQV/R6M1Alp3tUk5O9jIBAJ3jtFOIWMJn7kCPxq2VODTa/+h99gu5Jn2
zao64/P3hed4erzkFHEY3lpXJTZdbIOdGN4mcchoJuX0UgHUI9GT5XsR4L9S5JW9QYF6cp2MMTVY
raHNPOJCt60Ly7hXXj9XIsp7FczVPsWkBXQgnI9U09oKL/YyxUdUisnFeikDQGqHAitD16SNp0LL
AGoFACt5Ksdb4j+/G8QuPk29fkuv/pyJWw/MbRQTi1VhrVTzpFS4ftU5ja3hFOWjRqmue/e9QxJ6
MPJmVWttXnV+O8m1eWJDgj0cVqq5OxRVBJMKU4M1HtwKY7dy9n2zmzoS3f+kB2RYi92Ignf4DVAY
I3v/vtC42lO2l2nsKBhvXQNxjPMnPnJTJZCbQqny0NtKF4EyeJC/OEA63mVdsUscTK2mBfjfUhfP
/Oy/odgGh7HpBpX3YK6pDWhgFJSXG/Z6/mDekG3Dw1y33vGWgqSY5rvON5+gwVciIqs3NpbunoKQ
EhT0uKuNluar0TI7DnKLyJy0z6W4goqDZhHIr+eUTZk1yNyomgo8yExrfDQWoF4oqd0au2GshO+z
V4MxFhzu96TBM824MvkMkYbf3+2vC8ABzj3zl37o1tV4RWrBaYSkHR6X2P3MKAlt7UnTjbA6Buw9
u0Y7R5kUZuSZ8Zw+5CnHNykswx9jEEtRM3qsmgYsRRhjd76G5UgBbWDaeNSjK2z5qAB4/C5zOE0P
V7n8pWFUIfXR7ZH1x43mheSKDCWTZdjpuGmN6LeugJQF9vwlBTLHtVPqU2zu0k03Yf6EBhmXtHJU
F418AYq8b5XGNJEDpxQf9wOVNMOxH4/6ZzkLZAyES+HVXAWxJ6XSQrdRTXavVJLaQRjURTT6JfdN
haJaIg+k5KA6VSHO8lXfjUWfPrmAf+BTblGdad5D/hc5w2/imq8g87wHLqLyDoZSzfegiIuWmpDA
mTpBG9ZzfHLEYujcSsda2b8SDWc0DDrUfWBrpam/5ygUube+q9iDt/ECUOkg1sPBSyAv1DfiQDc7
cWdEQozJGuPH6WHXUnUl85WHxfLnI4t9DUBsY88PE0ukwsqz6YvMEYCPetcI/Dl8ovExyyOaoRNo
jBK7sYxTuu5K3KBroPVRzYujpSiheDhiOz4ruCNQOumj7CbD6qXmASm877IED9jd48WcLI7Fzo9o
ec8G6XKM1dkL/LrlRopKXOts+9cVokaFk2bVFq+ziZ+yAsYKS82GaZi/E+pa4PusMybiP8gln0iO
tOD+axBeehF8sWWMPvGW5qY3wo0w2P0sYhHVk6vHfN+TQNHiLr7NG9RUeXWmHrw5r3Gz8gEohLDd
lFnoO3cd1YAIdjhfuj9JXF2ImSnQPAQEC6EDT3jiHU83TCLw9legJR55Je0ozlGir7UK6bpp1CJm
zE0N3pQ4yvh8Jod0KF6NRLnH7F7XS6fs/uQ7TThATHoCYkSp2htKxlzB/Cn5SDWBrqaYtAAT9dEq
BJdQyv4gWMWUTFtX/xTH/Y6BF0/X/X49888shq6ei7wC94UAISjMI6/6BaIuuK7QePPwW2ho3GkR
y41EfZ5jBFZhUlU3nAjOUBVVGM5F0ho3PtfSWclQ/7q9gs978uilZkEawsl0lMU69OOCKGoVhcxZ
l9ouOsY7edCY1fEY3n2nzqiPBok8njdLM9a1g4xn196QkC28HdGEUCTYDnSqnuvL03OQO/2y9YF4
7jF56I6FFTQpkrT0YlUX8bnKslW5rf9N/wx35aV6uEKF4Mx+NtUALqMQh3Q8rbvOG95oO49jvY+o
9x7czmGrwSW6cet4X1ugUmrac9mD+Wbtkl/6/WzamMTzR8eKfI47nJ2bm0e4uyVHdeR9iM6ZTcQm
NOVDx22CSCY0c8G1fIDllmzHc3Ab1yFr9pAd/KeTb7Y9VRTi5A4cUUoIUGt17y5Uhsghf2lx1T7A
aXjIG+40QGsMsZtxh/KXZnjZM4KW6b4c9TKt32kN6U6HntWaexbT66YfZsCokEUSTWKMYPqsTNM1
Py7D4vSTF+m9tTlUyNpuuXDsPITk7Nokhwrj3IcyNteAzbJ6sU14zo81ba80IwKzd0b3hgA+E503
LWi4gbdbK6a4kVChLks4ATIW6lTjfeCdC6XU8cdl2Dpiyo0kzKnu50UIvmQX67vNV1yo/y0LswcF
d0DMN0nFySyetHQ0V7mMEMldt7dlNf68OYnQz48De1fL69r/d7i3il3ywc8+lsWE1DR8R+VDYlbK
SRG7w6IuV1Ofq2BU7rjATM/qbSrRCInViR/mbc1ecdAJhxgGpqCY61ZOzRy2uFwiDyHIWN2LUv/M
AFbCEZDj5UCSaQe9ol82j1nT71+EU8VWaMyf9MWNJ9JuecelCavTPtE5CmPiAjLNZBAwCX52GMMh
PSLeWhzmywAGsqNBcAgJkvVKR8QAHxsJUBsnuPATb0huvcO97O/4V6KHaG308RJoPuWLhx41Cpss
lCzPZeZ6oANg7IITmSoiSWlOWj5kH+iDjL0flEZOq83Twq7lsh4fLaeOkhnln43b4WAXnQxcBKYC
j1zGeOvBH7uEN8bptlqOGE7LGyMSNf4/ftmXBpyvnJ/OfxUtesZtwi/qMZmrdtx2y8vWA12o5J4o
atBOBXOeZxQLlDk2sJE2vP0TQ+FRpHnUesf+w8ok2/IG9GFKo5kbD87X8Y4RXMV0XKAn6fhYr4CL
QJocqAgxqhzrmhXQK/ZRWEX02l8abOvyr+J5kgCgg7flhDGOX7C1cnYQZ5kRPSPjyWj/T/Ezn6p5
3z8cogvXGm4CaUMdD54LvRFmnzsGUVIfrUFP7KPjl1gc2Z8xw4OaDsbSK8fO0nyA+BKXnoguk4A6
JsoHUw7la0X6S79YyInGcmK/aX/+dHzV81P6ASvaSr2JiLrEBeawLGG43/tD4zhebepX0MDXPhWM
e7IcjYip0FnDbKN7/o8/BN56riW6kvCsTdacccwKXFojFzM/3TFWWXc70mua0QZhw6vk2+FiNdO9
Al4d09cyl+mKDFgsfnRD5ZO6VAasDScXXSRzQNyJLIRy9HKqjgmHEQ+N7rXjrJS8pBQqF/Asrn80
YXQsWdu7VzSAd4ciXE6hCxFA9gilfujrjaSGFMwzytgexuZpknIJc5Jjr7L5twklqgSNJSqNv1/w
iwgULTlTLmVLcVj8+6tibax43mIqAYsEUXO/rhxDXP0UOOKucDDWqMcjMcsdwdOuNifHkZTrCAOb
haZpMDuz3aLnQCOEAgUB8ZbsPINYbnwQmowOGrcetgnk4gZqfdBoBrhAo8TE8LyNkhmdR4HHnrSH
uiUGrp1FH8dy0L3Z+C01+NmH2YxERYvlKfP4Yo8ir/j8lA1PRmv0Og36sIiLLiIJyuR11ECYLziF
rCgMjFrLy+0S23QrD8/4v+oL74eUkj1kAPQ0qppcXu7m/qMpPG9xaZXfnYUB3Q/FWfexNSpAc37S
OWMH1uZx/hPgpEqSH5lyorwVLspFq0/SUlH2EFw/udW6SQT3U/Z/no3T295fmYRJm0Qyva4sSs8Y
GoKsJVjK1JMIwEGmBLPzuXLXy/Hn6HnyPIij+fXy/HdD/sTDsuEpl/UDGOym0/IBKc0VrTUYtg0z
pkQt1ZgXzVSn90AGGUuL3YNvRwEZlGDf0/CjdRWfsTUlby+C1U6paO0ujQkruRprvzJnZ7ovFOjr
i4qpmAr3OklyJBwldQbgc0N6XgqZyUMQO513aft8le5iZwPfJSC2LdNV+9sCHER4pv9dDGsThOd7
bHIhsgPNqOynVCVgbxpyT5bKY9ggvB89zeKf/S9RiaewHu9UFhK23R76efWg2Zyso9QeqybPCjeX
lONnx9ZDJ8eR6vkXs/vIS2d5VgWSUYeSxp3/wFunQJH2kxG/RFmEo/wEPCJQOQzVBAUtpyc4vNEb
U1nn9+BnNnfQUAqc7f8RADyMMSfyclNVl+1b9Jag50Qv4w746IDRR+rhLm6a8NDa3DRLqTWnryNE
s2Lis4n9tPoV2XzP3OEoAUrojV/xo6ANVNXvBXjAHKfp4gJze/gC2pvOMCgUWCK0PiFOpKV8nIbv
+ZgEkQhpTbI5tOJK/Flg8oGvMu6u/6argYWQTxRqUHP6EWW4U+/lu5L+/gslzwxNWIino+J2lnT/
6Ob+gnk9/J0o7Q11eXfFElSFLk9I92S9CbNmUM9faeB27xFbgp445ygu92IU18wu1rEuWjtXXhhS
4HsVIrNGJ7XvOrNLI8Wbpfr2yhX1Nlc3z+nDLNxZsuoYCw3YESTxKgDY3PsQrqXDvvME3r9oD+Jf
3VFMkZk1Lc8NekonL0jQlezUQhpzoS7+72olmGJfZdeLRjtIuFaeO5OS0YdmjAEHvz6vKVeZz2jv
4WWoXvpY+VPpPz5rrVJOtN+jWhehS7uMMjD/8mLfXDF+eelxdyi0IiGJEEBDAcLNSBjNXHn5z3MR
FLWH6yPdQ1xNdvrr48i2G+2xLHlwwt4Tdbwdn6Y/IVpHT3dL7r2zdNBlD5yKzLq2u1+3k7nAqZjr
ulYLxub0Tb4doCcV7dellozFUvs+Y6bcsvIYiOC5ZoTy0ZDyLjCRHtaaoq01xGnjYbNDt88ZXaoh
7tBVp5RSl5uaGPJ2r97en2DRxiJqWUVKkpaFAJu+oCtQ78dmIzJe+jsZBXmQya1JqlRM2aYb+4LV
9WHsokYIB7/hQ9dGD2x+wNdTNBAGP9jO1KTpQ1Pikk9M6H36mnuOB77PxxsdbnrYgi/3vP0FTcom
o/JUl12vZhnT77/UdFrloQPf7Rb5LmtS2VwTULqN03+Fil5s2EwhLE6KDZHuBv+CdE+V0ny82nNP
M2mvHgyO4E8HjXJPDtK5NXKJtKQYw/KFdWPRoL5ALjd4rmiGhbJBJIMQR7ACKwcnbYWLDBggepVr
s/bPolMgvNdU1JdZDzWO7HBpfQecFHfFiBSXy1OOmjhXnpGmBypK0r7VvoxPvTwQn0FALRfcj40Q
9Cm2DQjcWJ42qSl0bMBSuH4Xu1iR09uAiY3YfOHwjyLw0us/lWn0FaOWX3SSIChMKLIPTk0KO8uL
tsd8YcK3wfBFB2mCQaeeMnNx9DSkuT4RAlxKHKKPOZHPLQ6bNOUZq9Q+qS7p7VylVHX75MLQXBZq
VFtaHFoD/BFAIVxRnxYsLlFCoEnINeUY+Hz+PPo8hQygmNxy9Dzl8M7MWm2a41YmGuBXacNlJ64c
CTusbMa2tttQHy7K7CcykTcyufifSthS9OOtTopHrvY1jQpvA8M0NPoHMqLNIge0Msz30+YC7/LZ
ZggpSe9pxGqn7niCI20ry9mLbcmOwHAXwWeCtAjizJPnHBd7/rJzTkfBBy3N0ks2QRBCU/lUMomx
fANB9MBZSVIgx3xy0clKEH4Fc7Rnn93IUeV9HjxUq0F7jyj3xXIwfQJK97f+nZd+LG3llYvPuhbY
ZkKrwa2hX5QYYsWF1IlLkR0RLiS+xBZ/Uw2QiVRDJAAUzLcvIP+HIEh2KpWfg7xHPmdk3XxSE+h2
ySYTYiVoIqacepF0bsmh5ZDSRS9Xjx8s3FLuEGzE9Q4l9p63xdofxlpUUe9CGhub+EvhesQjJKtJ
HoafTajrfLXQBwIy94X4/joeWXP0pOrr9qMpRnal0riaE/XQYnqqW5eYEW4tmg/v3N0QdTr8eymY
6Nr+RmqwNWWDW78A61YWq7uXsh7bYjgt55qE9tv1QywMjZFVX+NDMea1nS7MHM+C/dHkEotl6ojf
cmLz8eIPbAAt+iGNHZ+I7IO/00ff5I24vCZngtNKkpsBBKBihGRzYRPX8mk3UXo2G190vT2gdhEd
KjER9th5hHSXD//vPuYavWjNvtMVdjf2qWeLLbD1PRcsOk/V8mXlGRBo7kzsLdQ+iorYfVNK1tNS
Mf8Y7b8axxT6C+sjGn6j9gpmDl+31OBgrTwZrCZKi6qoekG3GCdT4EvjrFpAPXPaxYRjKps2DAHs
nzvwkPvNDjB0GA7YlaKbMStLJ5fbWfeQJiC50KPl2pEw82uJGYqvXbbHMa5J+JQ+X3waIsiqALzh
iGbaHreuL1ESKc9NDJt6+MlxLu5Z6C7FhxjCNX3+PVTzolzmNc1MNtrE+CQPNr9UIRDlFP/3+0yh
lJ/W3z6rB6cJWQsVUjRBaBGUx1bsh/UFnsy9opZ3sRXcghv1+FKYbNYDkZXCb16yC8uz0gktFmMe
BJKA4uhzXUuwtU8W33USncdTaqrUvCMt2b6aMXJHMAHZtFbkzbE1He4aN6Kt5gtZtseBMM4fLoau
iGKexM4Yi4qwBS3xZCXG1O5BFdPFAHp1fVNwIKX8tVv1ZJAJLR4tp8BMswuJrP3Yl5+MyoYfmX7i
mKloaXMZunBkA8F83hnVS0qAf91Xbv4vQbe/EzJAraAkOPd3QwIjiQcOI26NDuT000Xfgg0ItNHV
LCHJwMYBxn1xHRPWUPoz9w5DyUEvuG+yKVcCJdA1XRclLGQkK7999AKeGPeWa012R1NrTdGarV/J
vBTPxeFY6mkwEjMLaQCkqy3TlcZudMSSjRFJooxbZElaTvDHRlDH1TsJ4epYJTE0VYjVsgLIIHo4
bnTHNaQvR0CpgnZVLDJjhEWd63lpgbz3TdvRDiOCQsDBQdR58WLrRdpJTpR3/xPzwywZHrMu/VCn
KaN+mcz4nIXUeYROiZDLfjcEIQ1IxxhFXmMO91yPkJADdZWkU0ceNDlPh1c65mInul2QqmokbrMr
hPDijXT3IwLYySutaRDHudq1RiZEItlGjHq8YfkEiwKxhc0p8mSH1ewMHkS/wHeklivdKblCTKj2
oU/1SHe+saevSpZ3BGjmPEPSbOOiUHT604GlCcFoO1TvuDINnHso8b/xAvFMcvqRpznQvzpNx2xP
T8QUH2Dr/inXg+q+gJOwUbbLZ5dQ6VNydbxlSPG5lx7yhRZcb2PvyuBu2H/Jgnu9lPZ4GkYfnAAF
lQ+APyuIc+ghraG3mJgv28xIH7YNvKA0K4dm9Ggn8s679Df3ISg9uZvPkdBT+EpJuGJAprIf+/r7
Pmn89/EthgSNupbQBV8ky07RI7XIBdHDY1WLgu4q9hJBftUQrbFg4Es2dEulLMzwYXr9K5AcqtXZ
jYahn4sIr3FLdWIyGjb+qp0EMkGEu8/L2gw7WB3tLkEViRshOfd9W4S2xD5VE8JXg2boYJIEXoNW
Tv08Li/UnFkL2IW51uHbQof0B/H6FRaLzqrkn2IPwHtQUXKYEbBjVzcpVQcUjD/6bRhJoFdrkm66
KVlCQ6+HEmxN9A0qpgIkS0Qw2TMPqKy6MMT4mZp538dWJGVI3Kf4crciJhW7aZktshIU6FyjvH4f
6+atpuo78I/dlsd9Q9D0920vT4mQMuFc65YNj40AL/l20lDlzuv7tcTJ0aVKaFTBIXuJunbVEbf0
48UH1rmWhDugLelLAdVQkWiif+AlV0WXgnp8b9pZg6nSf+mo2LaYt7wDZNTl6XbZh0SPpbetoYqJ
QqALZ8/YjmdWnEva/o0DKFykhcCezgqUtc0Wz8bLL/X/j2PgyOXrjei14KTpeAO3OLb5s6bvZoqM
Ilt3ZZ6Q5FjDpvHG7bwXhiE8eVm7Y597K7UygGc0daYGacYwHAkpmS/VQ05mmgkArkekGdnlovXt
2+qw2ZZfvSTycAtekDoG+fqzlqlhhduC19POnzUWcedvfL0Qb4pdGjiTF2yFfJKUi6MfkFKFVSdg
So9lnvY2UzNQFpnFqxIOYg0U2N8yXNuTQV8ew5VOmliktw0AWZSJVpJfW6/xevckT8m2weSF2Zyb
ZloNpfh5cLOHNOAwjTZ0wnv26NX7kAzcnPRVJe54Quw3FoUATBF82B/L7zzUPObE3nl9iklWOWsy
UOtHOeB2yWSaSFSvM7AXbMJZrDOjkX719zWfQwWh3UWcAaUoK9qXmvCq7fCROx5xbSGsB6YqdjSm
HJ0+dDoDK9xKZW5quQldblDGCGLAjofih8+JLWM+d2vw9AG+bkd69Igej91jNXhVotufs0trZiv7
gdeYYSOJQWN3NsLrY08XTZlFSm45l+WJcH1DFHIIBRL4StZKGyQE0Nn8FTpgbYWUm1c/YhZbuOZp
7WzW+BqKpf25I3G9PdOhSqg3dHjxb37spjniYo8kOaTzpE6TbipO8PHsy2DtEbLo0lVydYSp6Aq9
0Lab28OIFbb60VXA6OF1pDatwfVAURwF4PKrzftqoBzOAzwVfeYZECr+TWSQXdnDBKIrxM5NqYXG
9nDSyIN+ZxzxEbjBQri5KC3NRXEAbncCQyh2uHlN4h4BeZuot2Gh+ugBVT8riRwxWbnupVkUkuR1
G5UQkO2iDKLy5roqTKrNiNVU4Hx4Og7DysUkZPgmqKwSGBy4UCmCOfItlrl/XhYiWO2RVmtp78Mn
OWsdPQ3uEAwoIhp/NYFZeFdo1Bh0de+JPIJwXZsldh6Uh0XwH6z5RgByrvkwzICkHt8MldV8Fntt
LCpUP3qwui9D/MKPFoHdkVi8cEUrLiDlMG10NB9wTTsXENbUCI50deG3fmGSCCzIEnnZX5B4iO6i
ek/swZvyagKCJNQ6xlVcVEA99mAdDY5GBMc4Qncd1SYsnew/zQL2s121+eoKacnqVdQloZoeGP8g
ZF3Xuv2HY1vgF/9su0l/QebCcveTkLnKJrmvMEqj7avssbehN5EaJ3L4BhdLMVnAgTp2kxMIIaLO
l0TCcdLPwxrh6kvfkyK+jFIDqSLnSpocUZG8hkMsjIChia9kNheG1agGwqZrrg+pMoRMsIdgT+3o
OW14A2UPDVG5OUyU9SWq/AUq+XAvYdMvFM0nq4iZkiifJ7gtBtly5PATaFTwkWCmoLrCjW5tUJXI
8RlgHH1eWfk7agCpuc0lauaxJ6nN5Q6OYT/GPqK0M0iyz56hDU3NWxl5fz9o94r+l8VmS4u4l0+/
OjQSPEEvHf5vwsTrzg1Cpi+ER6gdji8KNBYq23v3sCW8xCA6o+RneyulgLLlMuHvZ18ZocQgvLb5
3IDFzOcKcGsUVkUwjI5lopyAvOoIgWHqnCb7uynpQQZgp6CEKv31eE8PQjYccbtT88deSQHYoB4T
jpHefS+B6ARTA5OWuQDnPS+zXsj7Ami55UzY4TcK+QP04PWjpwJ/3AfPyjmpH5guxW5TIYmkGq79
Ss45uJCLfsK9eIiZs0zoLLH1B0bXyEg0IORDLGC+KSZ9YbwMA44BR4TRnPeWgDIn4phH5T3jIf4S
gSeWAc+mR9aU0ACfOzZ4pSRgJrXAVfcxLDFzoVQwwWZCV7KTcasLL22Dw4VGGnTfR6+JQXnQ8fKU
vNXaMkBnSGiZWAZyI1PGeDZ/enk2RXE2prhwEw+J16grGQzD9SlCxcnh3YZI3HARaFE+g7bTJu2w
Du0dEJ1Oj9Do+ButhrMzfHwz8AoKOh7hATgh9NnhDVcboWHbISCvzYPNGT6RSI8CuZVIRNaRgaDg
MftY+fD1f3XCMgv+hHPyTi0ucZbTydNPzE54yhp8axu/RgWxBCyZSDZbctG4EX9qEad8TaEo+8zf
avB2JIotfHbHe9mbo9jcLQgM2fxLZie17OSkGzUnZWC6aD0/4gWsoGNmNGwdqv1/1ZRHsX8Mx3t+
luRZhe9M78CmZwE8ZVXmpA0lkUcZ1IUVQvo+YOPajnMOLOWxwhYvMmRsrnPo7Mr/qR1XxqtZSYlk
RyESzdQaC5yaGgNQUjwZN31ox9ILRopcSXbJ21zOc3Lu/gwo+H1L678ddJzYhAQfCFtlv01bqqrh
KktRsk2+8KjnVXnG+fIRFaovozRc2eYZ5L9kfkZtRBu02EbQv3Pmxw/tCrWPM8RSWhAeyQRE1GFr
OH+mVr1W+lPgdX7yUatzMRATKNAXAy5Iglsk9w2cvdqz+q/EWGailh4QunD9FcTmU682enjiyOu2
Mq/52we56lbeAQFOSmZNi0nyMfr6tn54FoYCBXL0exoxhAVijAE41PGIrYuzfl92/MP64R8k8jMK
wZMu4aNYp0oM8kTkCpNi5h8Vcdb0g4rKdBirsElZRth0nx/bLKXkpd9lgKW14uiZyJfj8pRwZMv7
5swQYOqhYa6lGdhbaUkLS4cG1Ct0nmV/tua6MWbem8BGZcCCcLUmRDdrBtKcqeghRbg9oz8lQnRJ
gSP+Jz+n2OMotRg3K432ZZ9vkx6hLQWkGHRjhmCohXWRAE3jqrefMM3NZFvbav9/rA+5TqBYuBbG
cLon/db8aXnspd9oYF14cXsboFPgyn88YaZC8almYECu/M4oB8RZ3A4buLWKT9tHa/p4VGykPgAg
405wG+Ck40XO5e0Kh4TKARQXFHSWCfKioAgADzXd9mXu6ZgIVeijl5JKJwwUAupHqoUk1b/mvuPb
fhPdy4DsLrfLWHTjJxDFZ5BiJCwAa8vHkozqLAHgRcuUfnJXdzgAKdmDxbORxqV+gi8xUZne3Fed
Tv2n9iA4N6xwdfv2Vv6VAiNDSMAQsZ86cZ2+GjPTRMOitv2drAwcV1QGcfxe10KF8PxGJV5xmXKh
mvie0Dek/QYBi4htKGM2YnQeSDCc0t8ZSGnBFWh04UsdPDS2fnh58jd2Q7FUNMch13BuqHWxg0oR
0u44KVvifR8yhp20QfdjOKKk+0L8W1NoBX9uxMwtBGaeFdwa/5PtnEnl/zxTd5JPXGKQ3qsTc5aK
U2sl/pNcYQlQc2elVkvOKpU2qxAEOW55XtugNxEgJUyerG/gWHlXg3BWNGJJuy7dvXCm3iJguds1
O8IiDrViN98U+6XGnM2Gtxo/1eORam4eRZ13dI4vo2FkhbOFkKSFfpmsFIC8HWczFVNjRd3s6ZCL
p6ZPp5eFvfEb+HuEvpEBj3V7EAhBEgF1gEZAlsdSdzgaKbVE6YhLDswYYtEr1lIPGku9UvBVxbfe
JwrOLNbonfUn1N1mZJvNXUgUoLG5wxNN910aYmivFzXgcYECHhCbVHFGJyT5T9FOHmTp6A6mXE+0
ujTTRWwKleLRHaUUYivHaok+/IVQlwSEkcGu6k5oDwHEo+WFb+dc3zikFOdHbwLO9I8lShjLvgeK
oQk92P5cUE4FFVasf5BcP95f+7dXhTiN2IGFFLP67UIZWb1/gW8fIVcgfZlgYEXe+YLc7hvOl6Un
I4fIDvoDWUFJWuZB0U7m+A5M0uZIVt6ovT5GV769CtN+bJiqPiVm86T2RmPW2bG+3pZPTpVjFXtl
0TsRQbhPaE6HRUKwXdI2SfNJu3dLU1zEY2LY9EEGEjnjWDIBuXZXHeawyROy1QpNPq5AQIZyl78j
zC2x7f3lACKlp8QDixtG+UbkXPLH036D5DsETov19DNqfRzLxQulw+vDWxNLW4vX7qPGixD/pGX+
PB9HRvbm0QkycH7pJAj2W/iEgZ0QRZUmvPUAyHL/qZPROVIAWnGjOn9uBPbK9sT9vzUMgE0vO+9n
blWI89LwOBSf3Rpl13LsgHFzMq6j43CKD/2HSjNsCZ+Xv6QKI3cQ179l6tRjtXX/P1v3te9ZJctG
F2/BPKU7VjQWxnnp8qNgkErxkrY03ZoWjDQnv6//Cg6PJFGf3po+zzy/FhdkHJfgoxZYv5CTGeEt
3oQlsdL1JHwaYW1KTE2FrDBzcvjiqoJlA/inwthWj7Orbbp9Nb1MiqKlHJtW3P5DdBvByXb+ncEo
IHnsVpry1d/X58IoVqp3Qw/kSIGSb37Klg61G0Pm/q20PNK2uoNIPhlOtvxqrhCzwxG87H0k24Ed
jlPZudnkv0Mt2AIbFvyTi5JaoGw49bUuH31B4gtnHdVic8hYst9qkHOQ81n+NJYEYuH9ozlqlOHI
6YVJnzyWwmjZSDgxbEA4gA7x36HyvQ2rEKTaBluOpZfDxoZl+4fHcro7Mxgjjcfkopk+LFlpt+Tm
68lJL6vjO6Zreh9KTHEindmG4HCkrTKqUNfcKT9/wK/7kQa6xPeZB1RNrSBRXv7Gi6Qcw5sI5Tp+
KydA/iHq2RjwMuyT3oogsuYbpiT1UZcidVny1y/SLPjObgLslbeacWrqKmK7JnzIQxOyqioc2J3l
YbFHgocXNua8axEAbjDCZJSYlD60grVwW9yaxnXRjzEf0PqPljpqjHlcwUV8zIq2P/DOd768cxQA
I37NNm50pb2CyK+asSOjRjOjGO0sBYpbnK/75/G4zrxESWakkrMfY2zW4FgttzwPSxXeufOE7OVS
NHOoZViHPZngVLcKq9f2KWYg70UMEKsKh0wyNVJBwz7kfsXGT7JXj6Nbsu1x3R4Z0jFmJgHE83tJ
mjlINpRw3N5NhC3nX3gKnz5eEqF/hKq4n5i0PGnBMuM59ad8LPYkZZaGkjwTTIKN61Bl/9TqyaI5
xY1Fh6ZnwRjN0wpsuCl9l3VXyxPRcLQl0zBwHqaZWVXV72aIjFDCNB0cxcCFZLUiL5ZrvBNOpCBG
GPfnpJkuT7PfbnjFhY0zh+vsLTT4dChKXLkCdrCkRf8CW0YNdmu/rVsRls29jPxbYogXXKV87TcC
KmI8ia/djBdis19y1e3k7VhosMQK9A8lDA3p0Jnk5rE3HWn00vac/Cfe4uvxCaMOEG/qFkJ4I4zL
JfnWR/lDqxMHEFuQu5+9xMMLFDUHIXRklKIW8IvGvpOviJO1qUKCuBXv0kFNSifJ8/JGpqI8f/NZ
lFOrww+JeYMh2r+ZvBPJZUOeLgCGHxweqX+7GVjlWy3qVUzqfQ6iGA+JEpWtigIfOfC9BaJQZS5k
1TiEbgtEsIGS1Z0W7du70wR4cmALqlGxD4HXjQqQgFERP8ZCIdFbgpQhowthwBRQ58fMsW44gV3E
rFXkvx8C0rs2SZf806tYaj4mDDnJh9ZRm06Hka/gbq5ASdEQoyjA46UFUWT1JbAAQknd9fTiM/rT
6OCtimjNzVrgb7XifacrnmvFAXcAeAstZpBQMYFwoJ1/Ob7bu2lNcRYm9uY+l+w44ZeQ8oKheAlU
OLmxSr2RlT664n9hZqBfg0RO5dGw3QuA4O6mwzFmpiHYCQ5TECl9qT6aGH+A89tFojXKv8ro5APP
/D+S8RVNqrsmPcwVNP405NoPmpnLGI8o+ER9fBgp6aHL8iwwibe5GfyHgaqp1AV5zVlYPfL2lstR
KWj4ZxreU89bz8HBfRAtjSbC9q1mIE+BcK9FEsaLpVscUf2nkgnhRuDSgLuvPuDLYjxUUfevpL7t
hYm4m8W0tp5ubWlzUS2IQHoSN2s1KcLMRRC//OAH6dRbgBn36rij2nLdhnm9+jhXnlTExAtWeihN
I9iN2yydW+EDMuqutmZIo9TBm4HmWvAGT6syhCC+IckvHWMv3iOp7IGIabGbbXnu13Ha+NcTlJFd
ntZedI+ACjOLVdo5Ga0G0ak5ahNWoGqxbyxG6xZkQau7CknjLHxnRBrr7vv71YMXHHm63uIpKLXu
CrXwS0+lgmyBn1SOkmwcqvX74L2E7Iu619LhTklsKeKMP7zYnjVKSVVOe35SE1K/yfcI02wwBHiv
NBsbC3BYX1OnTYl5vnaHqYFfeaKCTQgRbyJH3T2pk2J4/Yu7ioQ2uwvzc7QJQ8YLry+x8b2zo4r8
BGfzyIukTwYD/Mqcf2J6ZG2Z1saaeDU664t3+awIkWCMVbDQZAvHCnhu8oPSP9j8Erh7dAwmbWoE
S6MhbGpJH3WDelCLa8JS9S8nQDHi/6b61d9glYnAuMhVv8yWwBjt1n06gtk1h034F84twZU55CXb
eVcuqDXvNdnTug//UdXSXppMCy169xjk3LVR3qc9UrtsC/CF3RFmg98FLODKaQLPuTrxNXABCxMm
vDGMQkHd5TcWZJ6omNg4NIvAJ5k3RQAR/BjnJnjgHpeEbQdNgj8EZyVqDLD+Vq0WIOjIAzmgHl5I
92aP2xynyBpZCnSGKGppr9v+8yVZ215hNw3wRuhLADloIefSMvoxEY77EuPSCPAKq99Cd4g58uHQ
Uxr8O1r1gQsN+TZ27VU/hRGHbYJ+b637eB81IK003wjp34a8z6/fDNbfzFSTPUCKelbCd/+vXpdt
ekp09MbiiKLx5F6siAku/kIYX676yzTnc9ymOdYZw+BJ7zg2xGuDPF10w0F/h+h2Vk24IRKpajbf
YqKdyGyNYFbqUa5KD6NRmPSOzBcWoompTbKuIbdWyKJa5xCWtFHla2J0iH2O+zU8k+3pqtX/R5VY
fT+77sZz7hDMEau5UG2sIYJ550a6vhZ1leGzxYlkc6xcweWJYiu3/Cf2VywNqdJ9tTCo9d7qV14L
+OdTEKXkzOIxqCB+GivEVr0mb7n+GqijZqw8DExviy+/MgPMe3MZh8jLOuGkedTy3vLidHvGAskt
H8cXiHsnMRmWdgJDRACn+iJlygtJvCgaw92ItxeA3L1J9M0newHjiZsZlI1WSOW7USlwNoh5BAbW
PnZR9WPmsC2yLRIKIFP+Ij4oMETa9b0SkW8GUP0xdiNv+JD89XB5fqM9VBOSIYLGmsYl0voNuiHw
49UXzSDdgpAW76G9CTUP0H3N0EqXwbci5/CaByCUn4M2KeU/+Usk5cJZUi0jTe/U5bCteBTHL3X9
Mf4W7nSmShXDqFSp3O/EKckitLRpsSh2XnAPtyb3cNfvzHKP/KaB4TuzHa1+Jxmh/5Yen8b6h9Xl
/+vUsKGQijXXiWcFBElafpHkCXR8n8jkXkFuBUW9WpKkOvO42DFaYi/lPOlDsDYBhFexauqk8J3o
wO+CuHEWcgr6tGJckTNnftYA11ukVF+FGt7MDWlGL9YMC1I/fHHRszg+OwbQk6sRf6/h7l0FVSOD
vgFMaJqv4H2Ee87RZUpXVkQf1qbI54G5UkAnhyA1Sr51iLsMkuLhgAGL7fIPe0pjNboJDOJzjZYs
k6ynkbVmVi1gtnKm66hvlpcK3XAbjUzZD4uBTJTuXB0A1AshVz+W5VmgsHHGwAD/w2fDxjXuktIP
DbTBiMpZCAQK2nRO9fRX0YljH4efvm6f7H9M0cTFzjYFO1n5y0oHh2o3TZ4huDnb99UJmqokI4az
1Ulo22hqh/x85el4ujDgt2ZtkyVGMo5tOxTtXNdiv3Gb6P7zRgE+2/0Cbtk01pbtD6fMyZA+EmID
lJ+89YVQHXT6zZOWeFmAoTDbl1vM+xIvUi4JVyc949GR4cqIn9SrZOQCUPxg4HyDxOKKK8viVMNi
aiWweEeyTz/U4pFqkIOpR3RHbZu7Zya7SbazwyM8mSo/4cdg7NHlHGoJndJ9+ZGtnmVp5/RGeTar
rQRIDX9PN4tZ9hIFUCg9tmWwdbIknuKihUu70IzqryqHVn2Lo1zqE0BKpWVJO7LHQZP2lgoO6Uq0
h5UUFV5G42t+U4iv/E6NaEUFODeyiR6nJTano1XoN0MxGZMAPbo0BFuV2s7eEPvtiWbHwCi5Al29
8ixDX+EaIFRlTJV5ViJ7wiQhwCnSI7cRJGDP9tsKcAad6Vaqu/Nqd3xW36dfqlMS9wTBT3+lmsrz
Cwm9rqI/QGQoPDO3erPrmZbrh7hLS8LkxyPNEiVRF0extGeeX/U83dRIWoAgf/aTjvc7/Nc/e3Lt
U+hOcrzX+9wpOICyhBJM6ami7bBSkwRA
`protect end_protected
