`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
r0PjKNZwkpAarwvm4jTas4qSepqQWk5z6JKqAzK0ed2izYUSokQgN6Af9NeiqbZcxrx0nLdYwfyG
+0ZOf8VxLeX/Tl80Suc9W3IxexiekmxATQfeOtQk8If8hJTC9Q2HNJrjHSKPPwIEJiJKLoqbUKZO
xO96odui6lygNVoYEDRZJE1WUbRbW1OxLPKyY9Rq/iULtouuibxdpieCuy9JrCayfWpPF1xFbaAh
e93F/qIGJ3D3Owto6zgOmX29mwFBYDrGHXwFwTfpEUZ/PRhs9Hc3c8WV+FXFYQx9Wzof3DXFFxWs
EuPMSwtStTbaa/UhNYWlZTR7aY3It1+6q/aMdg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="4CdmwnwXEj0kfO0PDOM90KHqVIbqosNwWoaLgVMJkqI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22880)
`protect data_block
IBUIeh141Jpq5cSSrrnJX46RKNHQTWhJ8JpFAPCAL28tFrdPfhMf24hAIzB2Ro6SbUUIxOkyc0gz
jj3aLGjYGOXKKfA291Xtq3ADf/VUnxlUGrTyk2xe9PYw1/GHWP99w+clV3XjjlV+KYl8lC9314YA
+JAtIfVKpnjL7KBt8jYpcov5XAsSZqyZ9TRXj/3gnUu9/d5JrNQYf7XKL85AYZQisw1DcKIvf/ON
oXIGaI7RAggYki0DbyomL7QkUOTHH9jOwtcPbtM86QK03I+cNuEWr/NqJWpoISqyRt3IHj6rVH8J
BVerjm3vLalgPaZXFn8F0T1gZTqOT4pclEhQZ2Y6ZVaMmWjEm019LopKruojBsxvrZU99jAQGcy1
h8vaXEx4g5+OAenLHsyt/sbsu+E0BtNTyJqf0t4aUyDSFX25rffSLmnrw+IhLJRLdmxnaNiQw8Mp
DQIAO7RVBGjf/4vuMCh3DCV/zTrf3q1CIGZ6BDpOLZ6TUyIV81NzLSi9OlaC5XSjtHiO2QiRcoZT
JCPOpIgnPsIBZCxNZrPxsdHBgRYuRoyJaPcBVxYvf6FwbAJFS7EwfGs4QjO1rXe0KJ6yh13M2lEu
f+5jE0Hrb/svB7drNUHJoO585KszVkzZ/oyV4/yM42WjUAt8xKCIJ+xFXYeBXC/KmEfA2EAc7szE
FuH0ojpN76uS+4mGVrcC0UmGvKJMXhYEjTpjbXeGslFaHKe8wyhq12vePtfMvfajHZyPCNwD8wXB
5owbbvBCutFd9Rg01W9dfw9t9c/A2nhwL/HidRBsa71hWsdvIttoryuBTa9gkSamuJkX9Qp9AEUn
xsYMH0nzzTvsi3gKNL8tgwFCnP7djyOxITIHAQZD95sY6+YZSehrlNMm4wIT8PjDrtVTrkWUQKOT
ZQ3+tS1o3spZv8CSkY11sB9bCLt6K2RzeMv1HzRJCZWQcyG4f474T58MlkJNQrKgOYJrQmXnXBXh
/8nss0JVEaPI5RdraC9hbWCJ/XpMWHQW00NEMANVkLlhQ4Nfc6EJDn75v5YyDAn/gEJWF8LXXM0z
VNzJlnxHMnwmKLRw58QtN60atz8W09N0FWMADtesZ3zYsg0/ysg3taD7Q0heuacOeM+208IK9IW0
8cSxty2EMhvALJJwjeM/MUuVg9GLwRzguUwmWzUjts/RSv/LTPCGTBPjspBqfNLFtalsgvWC3iFs
0/BtSnNj65rHQ6ZKbqHgXuiS1jRQpRO5XdY74a0bybc8AzNd36BjVTJZQuPmpV82P6OGoQTsYqfS
NSb2yTHqor0bzMG8AvrHSX98u/tvToDPgMtBXjWR1sLcXY6KVChd+I/HqiMR07mrzSxI6CzKBpKG
W6Ortg4wX4ubbDb6HP7qt7KbsviCWzaJDRctH6eaevf3MudlPu4BnJwnmvNqI/+RQxxFL8KYPCkm
pLFedsA/KO5ivcPDggN6PPdXkoeHlzIMx7FK/5y9t4U9MBb4jiTvULTY12n+7lRDLYej7usSoysF
iSahGq2lGxYUF/COuip7GvVTqOgN37DJZtJGp7/XQoROtS/YLJnhnYa0d+G51VwmB98FRmMF3if5
vCs4KXgiwWB8/dY59I69T/40vy178cx+WZutVx5m+6x4xOXl072V1PRtQSXRpZYVzvgrPnxS/Pes
1b3T/HC2qDkFj0egP+01pKSU5IdrhrITReUEfXCwGdQ42PGgwZG3VRox7P8C6+znddkgcialsri0
CfjzCTRlgWl1itO4ldocVtY03M1dClVXUSRZhHwXjytcGX1f6GubPCqUMk+LLf/oJXoqD37K8POd
kasfbCxwRPTLkG++Beca/f6bFXDb15J5mFQgRxiaz7955qkNxEYVKlfTq4de54ODeWSpi69Qov6S
k5E/OGIy9MhnpHkZuMhC8QdiRK47kdYaSVd5pRyCALuXy+2RCgWy+6lFTaTOxyx7rsq/1V77J2Bu
N1dUPJ0+/Fa5F3j9b1kmzNDlT67sue1Mzx3vLhEpCKirP8SJmyh91PpRby1dH1/CI3QS0YtOIQDN
+iLXlBd3qfbdg+K4GvJrejXdiBswzCOCi9s7BGu6HyJojiKr1y3S1MKWO6JRh59rwwepSRO1+jbJ
mykUwt3r7zi3khs39y1kjubEKmsOjK91G702KwN5LK6xA9KymKgGRntXos/myubaUh+UFDPTzYLh
PGydAMoNKVGFeUVJ/bFbuyJP0FfxeYLWzUmh8IPKloFkOoiM1a76uSZFwoKuHCrhu8SWbPBEo23I
uXRfOT+K/sWiaLF4lrNDfSPdVuOtJP8TPFOi+Mhwssj702PBIqUfoHwRHYtGmwXLHSTYrKJjv3vX
y7vhxL5a7jFgzK/8D6K9hICrrXv0MrOVL5DO1k+llVayCJCCIVwHjdrpnCI4OvH94ew4oTiJTosO
pTuIdUZKrD2vc8qEm6WN9vom3zEo4J0Y7VfgACWC0ZVLWdwW+i1uXtD8TnrlR6dgCfvxHgVOkfNJ
gUhGN4+YDHupoDTZFLrkORBcZgtAO/V1xWbBMBFCJ6oJ7HpJqa2OzBv8b/Xgb/2eIcTCTMwjo+uI
iyDYpQPmYVlCVOK3nNVp/f+b7gr3vJLwxU+UYYDEK84ZkA45dvhEF/JRZXrnbkkzv0UexIQpkHDS
1xE0qK3TOa6IZLALHHJ0UGveFaLBm4nycv1bIHDpT9ZKbIDcm8gPQs3cWWPiU6198dwkYsoNKlSn
1oT5cSKF3OuaMDsB7HUpD1YZOns8pM3C4dl+LeaDK+XDP5QBj2ILrE0lorwhFgXmDj5Nj/QznAYj
xkQInk72wzmd2lFSkagOQmx5mi18EMIMh8ksV9WVn/S+S9iIHOOeWeeGXX2OMFr/neBtqeOmQjXG
99roNvIlDeyomer7h8/6qQT9L0VJ43QYwKmnjSyaHjIiYpMNrtXLxBrhKKYlNBd3RH8BfgLSjPAf
+FSL7S6HcoahP+roAjS3n/FS9xaOjI/uHIu4oT4KrwXbkEOOLKrCWJU2mqhVQYyU7d7yfJW9dybm
oCHG7LiNUWWoSnSihf/IuDMl1hqdegsaYZ+XC4ZoPMX//SsT7x3F6bYojAXeFuQyqaqvzVOxdojH
1FcoqW4Zcs+oZB/l4Sq6FjovU2n9jyQs+ZJrBZkvcyMNnLCB+TZpxns5eeXV34k/Sa30+6+ayRK3
pScnSw89evDKdZNjtPtlVZ22sT84D2dSkJ8ALEgvrT1w1dO7a8yltbh+QAGbs8b9EdQ7iEA1EorK
NIdmEaHx9x4PNdNoR4rrUJSOD/fXb0RRgsPWjiKheY5aMLKVxFKG4DbqA7N0HH7+KdAgHf2j5tI/
caR+9YrU6QDrcOW56sF+nQ3QkfImczjJ7gCbgd5FHmIKAeL/u6YV3BQQtzwL1T0p9ZbYA8NE/qJp
xypI7my00qsj+Wdyq9TDM7mOaLvJjA1dQOEV2tx6Hg2F40TpylE8N8XUaOYlRP0B1BaK+g3RFh6a
4nF8wGnzx6PHcEJjsRL46ZNl9SK5vc3FCqTPDLHIcsKA4toZGT5mpQQJIU6zH8cc25cu8KVeI1ZY
PxaT3euNBd96aZgzifj8yJB93BMkl7hnLYHiRtzGv+RVtQWCCsaM4MewCQ+alXmRD9Vdn5cF7ko8
I9PGK8ZM1+vNhoU/v4WRx862wA9/dQZea1AfNmQdtnFN+L8+hEcgiNl/Nvgw+PRMqc+2aavQ6iGT
wZEKhCvIMB4Hnqth+/Ad+u/c69PpmUOVdW1TQHSEExs8BgVh/DszqTerODjPbZUJ8z+EA4Ami4Nw
bsG9ybM03gwm4g99pCnkChP5xXzG6nkehaVdGvs+wbHXvrZOSm+jDMhyzXaacW2GzZbedwqT/bXc
9CGMIzddVthIUzcvFRc3dznXA2fACKIxRIsit0Qs7WBYTFHbkc5NVytDXtnTjWFKpkgPSnigM5lQ
GOCz/MxGibm08FZdAhbz32ylkNZIGTZ0TMJRx8WlU53mIP5QOLF4kLEcfY6tXBHKmENSRVza28Nf
/YigQ4C1JuEsmSilGehtmS8trweINJEskApETp4GfcbAhKJAFa9YhdlgGt3W819k9s7/Xqgjylz3
CrBwp2S3ZPw4wgCoxGoraY/awV1Kn7SSXoWU3qMD1HazxZ33g17x01Yi7nBh4pufWwDQv0k5/+jO
aTpVFupK4dQtOIGmZBfXXVSSmpNVHukRSvvhgjK8frr+FXE9GZik29Oc4fQW39dvr5Zx0u1+gFvA
VNYvVQXt3wuM7PuaJCb5YDnw1x+zqwdFHXiL43PnsuvFerfectkzU8SVbr0UjcxGBysf4SSPbjIl
5sEhtTu/c1szNhU7zIeKdB+MLwHxt4FFhPuqeyhf8a7ufkk7HNvNTc7G8Q11DMgcSAgyrds3Jcnw
tbXL6Vza283G1zjpTVGB/9vI7DhGCW2ePxz/HWppBiPQ6HlDYanHO1q5yCdZgU9jBG3XQNmNcGRt
FYB71ajz/yQc8ajD99JjX2yjBE1V2aDyJ1eETxurYWi4kDibkzHY4avwshW6zTZ3f08wFaGvTYnK
v9alAVc2awGeHPQyMINTpakX79xAdYd1ga/Wdh36NUgtGukye10+ATXW45lcj+f+aPAOLmsmdjCB
bjeDQl0HWc4S/JPlivscbJg7qdFIcn/a9sEiV9/q+ma6nN/Zczr+J6eqHEUECL0gAsjjaCJXhX1h
V3mshcpEgWcUBjuPoBuZfcCuH2d0KPfH05G647ul8l4jOR5skW5ndXrmNls/xyE7HCuccqaS+jlX
jd03QCBzhOv1JgZEAVmlVuJZBZBcVPzpQLd6xqYwduUEfwg3wVF//CXdCPwCNog1QSjutiQpnxGx
yBjLZBVEGhsApBSHrK5dZ7CTa1VnCSsl8MDxFGjQv/ATlwDOhFil05M15igSTX6gx2Zw+ss8NjYz
HEWu8kN5dUTq1CwSJjN8Oro0a1faNa05KuuwSbR0NWR32YYztw40HxkgNOxf1p1EBCmMqxl/V8pp
p3tuGXX5mxsi+6LgfNi1p6JFKs+Zko4/Ya5soYPksajEOZSO68qk4jKIThBC6RA7hK/wfgdYYbpe
najUz1/bEsLdgBxJ2iRHfWm17nWXSqco4lyodr3BnD+rkuUkimp6rndiMb1yvIjy+KlVqVefr7/E
iSC7X4oECGqiYoP6hI6pDSIxN1sfIlTpGW3vKW6sxeGjctx22L9mWRyDkAs5mS/2cyM2s59/q4la
LEJjbCz9F5R36MhaRrCGOwjHVYI4LOqmHQGQvLht0cDdZ5UiJAzDmwZXKHnNAi3RRKqkOXgrGQcx
M95aLqQx3CHFNQWU1520RJXvCo55+mTfBwYKWNHXoaIW7h4waMAEdQKKcqyfvNjKsVGGFF9/cJRr
Ht9u9yhaVJe55G2mu81CyjVotd3L6yYzkX5HpDZ0lV4mxEQLH5CQFvgZLX+FSdosyf5r/ma6h19Y
zOK6+28cQ1od/MM4ITHoCqmECmdtx+u0/SaM4nseBfOtu4bfHDWOF8nQqyZ1p1XeJ/nsy1ICVorp
hoB3UfYuvI0VXUJsP+Klk0xZRdFLYqyC7paqdDJYxl14cUyqxtCQBMOOEDlg2Dp0VSyYaEEKPDql
yVBOY9V/AEe3vJ/MTkXrv2+mHVpVF+5sb8VFMfAPPxEcJpc3OxXyEU8P3MTfewSZ9FlYQY79qmm9
X58E7tF/ZsZF9rPgnDgvh9HQuBP9tL7LI16KnXSCHRz9clrgO3QruILLiIyfgoC7S98NRiCKLpy+
m8JinBQTdhsOcwFVnyraeBEZZr1upMN4o0QkYhB83Hy+Pz6bFmD0kNScbS6H6Mcl/Jy4ImtjYzaH
V392qnopaPusLy2oouvWRpMfwWKnYziAOumiiHQLKU+TU5VN8m9AFJ0BkVGHRq3qI0mlJBBU55jt
Vmlj+COb9+fRjwjpAv77Dsqx8ONCHTHsPDKPwNrRcuMBPwA82utPlBlJDN8Nmp7oeaY99pWHwoWB
8VTPSll4J6fgRklrLsrtL8YjSKnGk3pfA92K5psW6xoS4sg+NJiunoEBiEYcQ/iljocmvakLUdY5
4XBMroa9303NX5PJfshcMYgdmJpYkjod20y6oPYw9YVhqRhF+FT0nIhA0z8yWnJ1/Yo969YeU3DY
NzSEThCU9Grrz7GQliaWhHhtDejvO48M8L78gm+OjVQEFesrqpcy72vOz7UzuSZ10G7/wsIQEGTP
FJWOrZ+IEATFRyLN8H4GKxX4sU7KQEZ4T9TnHNgcRC5r6+pIW33Ju8FfdTogSfBYaWH8E+/Q0hFi
ynbNGHrMG2LYuTtx3F0pY/sY7PFV7Qlq0a16XPn/eRPO18t39sgVrtK/rSDYP9qPKfHuDJyqQivz
/FNSsX+JtE1xIjO+3YIVHkJs9NSa1sC+kiNcmyHBLi05M948kO0Oc17Y2WjZBNERK8+UBbC5Fw/k
Qyi/uPc0nWdcp22YBXU20HOfaEzNeBFigYiCM3erTxji9cJwJoqLbkZs6VFylWOSNg1EH1mPjNzT
uKSdHc5Wd2LBMXCcsQHlE3ZmGWH19Zm2v6m3ANo2Tr97bKLYGrsatthVEzY5tECp7fXqxLHHBxLK
eKGGz+0i3HPI+cfJUEelq/wy/UQtXwBwHU620AofDDDlO+KCj0lI9xo3+FWnrYYX5zpT6j3WyFYc
MZAFbm3IGlADhiXyK2HEYGQUqS3e9H/ndKnSbvmvy1i0DPo4t6V3clcNSKZU29V5KsXh96hrubgm
iqDjeWm0oYC96zjy94ffjvQ6eHIybG09WfsRAynDnXUbrH3PCNX8p1ZW3eiAzpBZiYZpOOBXjhI1
iOkR/zQzASYwqrgUNpaZU33bpVoFtlktZUr12pEL9hdhhKuUvc+WNOoztic93SkwiTMQHXhcC/zh
TG1Uo8fRaa6CI0OSClwMZM5VQeLvI25kfC/nZbmP+KmcrrX0s/7LMtsVC6BwDkMm5lshnOeEknFT
IFsNu9iKhkClyBWPm0bmML95jauORAEO3tEioOf1HUG4Imb3cexdnmDuQH6Ti862RLkUyYHsRUIk
JOT5ouhjqEtn58L5/enJABWEcbNyX1jFHDFCzjzpbz+jv6rdwQdXqm4e/1s4jmjHadfGLcy9FXtn
/wC9YCQDCagongmz96G//z0JLuX/6lk/yT357OxPo+M357OJ63YWDsP4ajVM8DX40P9pDw0a8YRV
ZqY3ZAn/j8rUBrJ7O84gvqpk9tUOhb+DCRnpAcw8EdEttKvW1AHJl2NN8FSBj3izenIQebfzHJMP
8GLOsyql07AWeYYW1fl/2HMsCDH7sBfd8vmhj5K0cw8dy12SxpKnhGkfILHenKIRb14JosBtZcMO
/u1UsRxam0xo0uamdk+1xceaorkU/m5RDIN9SBUfR8MncVxaaOYZZs8k9Ycb4HxYDy6aw3ld4QiG
Uurpbon7RDIR0zbH9wGtsNqLy7elUBxUkZvaims0HflXyaidgKpoDIMAZJ9EitnThY/EaeuBjzTB
coP2eSw+POP5bK59JTKI0ppdKK1RK9RgfB2IbBXn1dKas3cSfmBxjYHMraHLEjNBvvAgbbtlVEzX
FIeyncJaskvcy7yYJo0F3pb99HITWy9dx62FDMcuN1Hd27YC9zqW8wRSRRsSIOgyvTl0fsOXLV4/
ngWokhU4ywDDtVLmHTUCi3PCLE0TekPssgwHRWnMG9OjzqpXYT+NJixTeK77orL/UwV8+OfppZvu
n5Eu+LkkrOz8N++bnT8Mqki3QTmlOmF3r4V6+1tt/7tMlhMhYnP/T+vSuIMCDY3IOz0Q6bxWYCBS
p9zOJpeiGaO1craOEF2csHBTTltPOs6xZBC2640f9BMKVWZ7aeX3ABdZEeCKOhhyILx0xfbNlNun
XQLD5/Sz8HbOln8Jz24Mm7AbTs77Ela1CYxMoQVAHIcYfyIRa9FYnY6FgvIs2sARFhUlAKRKxJyx
AIIuhCR5wV6h5ZNOlUtad3JA3SD5+dAeLqqia5MCnZtmH4AZx4VrBOhW2XRGJ7ShpyIHxND54Lh5
1YF1EZeZ5mLdl96bw/8iJC+9U+jqhWuH9QX3aZ3c9+GPgK8IMkmPOywm9GNvAdgtLq6ueZqF0ZFr
HpJXAPRQg770wj4D7WTKZqMG2duTUJePQkxHeUsYI7BWTMXMtYZlL/SJmfNJKQHnvE7GoeXl8FPY
W0+XANjnL0zivr+TvZWyuNXhqHHPxl9tdKC4YRbjVMgvtZ4UYDfuQ6m+XHBywOhEcLmTPwTFjXjg
Vpq9KLWd4kH1pkJIBClCWQx6SqDWOAA/FYrY6skfijBSVOJjeH3ln9KE9eSkhxK+s4p4zkyYg16u
Bc9TneErr26vfFNLYAtbDh0tcCqwZtzi+Qjpk8W4LOC7QxtlX8Bl/kXXp/Jwo2JtenO3RepMjb7w
IctDSVGOO4tz2Log/KWCC+bCWamGFoTVqwPK02if8apdqqI33Svcr7tELhYc3s8zoJ8BIppOUYBf
roR1ASkqs2Sb+WwBmh4u/hFoZTqsBvOP6AUbk4jlAiXpdd6jDEiYCITPJauRKIGeroHsFHwSvUIs
wXbVGa4LsIylp+62ssfzwHkqz6zjtKW6HGjyJwIwkfC0HNLFrkUmDxvBIW2JsQpR5yQ+qED2c6ZC
DzxVvkfyCIqraefNxCDqLhm3yEGNXh/XFpth73cZKNeo8FiIBKaJp3nGVxsESMpEBUYT92cdmgp3
inpv84vx7IZbCYjVepiJwq8tejl+gVnlJdzhCwPM1WUYakWkwVLTsO12bZI+cQoYT3Zu+DiTdIdW
JCdibJrkBxYWgh0b75NUaTjhgAoYCA7g8Xu87DzTHFLjt58lhjAYEkxC639JFOCJWZAqFuR/vqtu
SelijWWSyikuHYJs7e2cQ5h8kym+YlUhPgRhE98PkXoj+83hehm7s4n8VpMH12WmBugrEXc8UFF4
O1Xg+QRztBPyW3j1vVopZY2TKjRviPhPUiEOk0GGrtnd7oFIn3hDstZSSyPEy0YavjY55qt3oAWk
1+1EBzZKWSuV3FWLzUXv46KgQ9buNpN3pBoW+wHn4UCFfz0CHvrEIT+PBPUKOLpfIsxgeW+GSIGF
ZW1dNeWaa9+wUdj4NyU28H7XYvgwdLYFaihUbrFTecMn5gkxAlDfuZ6HgNwDCvlDto/OAJPx/uc+
jyYdkellH/s2VFgoHyM9y/5Bz53YAAR6e+Y123sKrV9PB3G60O6/ofWY2qtjyaiDaf6GxDfxC1Bc
WC5x8FQ9NSKCh2Jy+ZKkPqdsB9K4ddTCSqyga2NA6AsgJsSXBWvaXoj+YaxrRMc1o5zlSyqStj3x
KeGsG/tkxvBfwuxFCM/GChRO0is8l+UK8k8TswbE7QVDeW3F0+D1C6fglZQbzGC9JY9RBeu04dVy
+36xKDinh2+uJOm9vF/k77CgTiTELJN5B11IzXFR0gcjj+J62nzqq6uNr8HXZyuLCtdUpsQa0K91
Rw/uXS74pAVhqfKFKNIvYX8jJeNuWNUMjbpvnrzNm9YkS9MQ0tZGPRqmX/zYLzGCpDb9vDl00nUv
uXd+wG+ZPpcoxo+y8RxOssP/k3iRtSGbkvuNrgcp38NOTt9buHjnm57hLAQbMrTWAhaJe4epZBHi
Zk3qHzLBqCNGWkKncCSlz4hKnAIHTI+t5WT2FdEd1YP10u0hl0nX5xtsufg4YnqlfGlF7A0PBwbM
JQ9OyoSPmhlbO5FCHcz9dj38yjWmxVRmAyb6UYwJuslCYhSu4ra6ikxGuxh8lALjbsAbN5i7dDBs
qeZY1ndfIGOREMYWDVcCeuQwdkVG89pDutSCHqZ+jsTO0Ipg71Is9B+lPMYKcwFlZ0gdt0deJlmJ
mrHk+jbT5Xy3vUOSIPqKAaPzTH137DRy5WlWiqfZY8uz7kZbhFA/ZDfJRJJdMfMzuYiiwV2NJ+ZO
KzhyQLQYpcoSZkS0JtlLX/jYbD6P/6Ll7Hnb9r8Cw7uJcT9/jrCER8leOgRMvvZe/BvAZQnZLA3u
c8vw+DvMi0zEqb0msCiMJrRAdZIX4tzt3AzsMzDrOSEqK4gJlvNvDLX/eqYyY0l3U7ad0pGBBS1W
TIsYWZ3ZuBd9ZOqJwVh4A4AF3kKsHbiNRAp8E7ILN8Y1YTo5VnpTW728xvVtDp9mhGaWKtnVB1j+
zUuVwmt/jzn0/1sTTcUxTdpBpaE1o88xzIWdwdInChHd/YYU8la9nEgfvk0Wh3aRDL/Mh8r5xE5j
SCI5+fM/JmaWhwuNdN4YvWPkpvJ6DZjraqmrn9ef9GrBfQPiyzGiSZw9WG0XhGadlgB3yjwik9ZZ
Aj1UHBtM9upCSf3aSo3W0WC1doo2ouZjXpvghRK791aaBEMXTv8wM++jzqaHZBTV+rXy8ZQb7Nqt
KxSKrYepYi9gtypnuj9aqjDAeEFEyGdhLjTcDnB94ZOGqw2UGuXdxoW1LcDghJeXuNr7D3vf0hev
rXEf2aOKH4g+thBBo3PiLRakC/hw1A4L8p3XhJErpZRmgdGEZYwr2XF3i0aDNciS1ybVPs3bMTeT
joqSMCaxBg1EFzr+ar7B2Dm63iw89mgLGgw5pIHvlMAloTNBvvtD5Puu3EVtJwhzSQ5ugwKDYSm1
7Brj2kxsxHQFb0rXIC/cownEBRNRHu13TFGCb5WBFevvHVkgkv2ikezLCWh+Be5QGEBwB9fTokrX
CqK6DIWZFqqCfEbC2x0t8tepBfLsf1OEEORSjEqhhztYFN/H3amyjrHrf0xP0bBN/j6e5N25MlxX
/ft7dENaDAiyoX/zEkhi5n31osFc1wt10F3Jv5SM1MJ4J+VoxjVDucA3o3rIUL+ZpJSHBX4J8eaJ
hDQwAEEiVFfYRWoNXWLweBp1UahjnbSVzitNs1LuAFlatDxMu+hTT5WORrlMWk2Yh3MWzrfBnzLb
RHdYapSCg0HQBN59WKuG7CwNZRuJqBpBF7L5E1zkp/onYMeWv2Q3UKK1K24B+L78O9ZDVscCR36T
jiXwBK4eJo9LDLRBMam/OhrvuqD9SSb2711gj7VrjWihOviF+AUnUIWqP+JiygGmcdrap8gU5f7B
jnHkQEliuMUNgMC/iZTEMoFsBKKyFz57YK7Jm5tZTv7hCLtNnHOq4WI1uHfPOwcz2dxxFl768yNY
K8/p9/pAwjfSbaBuZx6uob+5m9g9ipUc70rOh436qLcVK8pIcuwL58jYCIYGLSTHACiMWPzL13EQ
g6WeBBbwpC5y7SMAORXLK50+ImUPml/AA9551ZmDFuWDEEmo57b9ukYsA4C9Bpa9PJ5iyILv7ZPc
LsurXWkg6zF4joKJQeK6etVYIhMB0VOn2IKbjPeWGTmLHH6LS9nNhAbLQ3/No9ujdhwi6tZWI2M1
Y72mpbNeMOPqoC6S6ypwpCg1xTixH/slLi+sRRqH9ynxZzcT3GArlcUvSY79msfqGpLkuZwxU5UN
RjkuX4qmIVvRdP3grOzoU2WIEDgQFaRV7VmbojmMnV1AUqK0q4tLyxqv3FkGz4zb2BH3NPEWBbT6
cQtZ0ywWnbdaBAsc/2a/+C0ErWjxqjMPsZZHwCr8rhxSflFnyY5kGLZYgaTIYHRe2ckL8JOJaVID
ozQVItppcB/NUq3nn014LHfLh6uBpbxo2XAkJK2YOg+Et5EwNeKnR6QYfaSG1ktVXnRA9i3NsOAm
ArA/LvkczzDGOSEfSN0GQAXj3DiYfRa6ErvSFs5pdUcjhagvUCbA/jwAmaKP1gpqkroQOpjYVuHl
Az8yKyghXmIpa+2M0WieKu8pP4qKNY8wpS7YHsK1os0+HfNz7Ql3D/d9Q3tRjc522LYy1dnwbkiu
3KWxcR+pgAINj7cnKd6LiIGu2/SqiOcTGiYjnyWfxcN7fR5ZsZ5wOrzpDDsvtfJr1M4QEJt7vyAj
e1E/974e9YBdvRMWvBsD2hZZ/EwpVw05gZSGjAeYGABMi2dFwqqvHQkfR0zGVPVEXhL6Ne6zZZuk
6U74+z31O88ODcY9ZCbtaMurq0crUIGAwKL/rqJ9GlMkihYMRWratRzPvyoaHHTJvGFQghiW5EMv
rjHQ03cTJOVRyjgvrCVSBht5ZZNGSkt91hZePzAHK9JIG6ZAbCV1okHEDWbY2hDvneR+jCOz1qf0
SvuKtqXI2l5U/MdLG2An5uSk131HAlVmPx5wWsby78eVuqhSwO0wNMpxH5EJaB0CClLMzOSSysge
PKPgd0IQW8T21Zv3xW3Y9UEgftfgCcoWQGq3dYiJSjDebiyOeJt05FcdVElvRGLNZUnhDOXLXkzh
E22GaneIBydu1nByRnMt5Wu5hjguBeziRgW7GAeTRtG0DM5gwrckdYg4XDmDK/02bjIL1LAomObT
UqYOO2WJ2mco03uS0iCzUfil3texz2DnHTsBj4juj61sfYP08FnqQMKMZOGC9hyJQRmR9JaJrRao
bZktmJFJ1ExeJZaiGr6+2XM3CECETvnIAbh6YFRbRM6V4JptWMcL1MGceXl1cVucFBmGK03upplT
/N+rs3feXlR67Pih/hkiwtGVtCgJ8bB6ArnsOb5lNRL9bTxl4MeX5d/YZUw3mSV2Uzkq5oO+miL0
ZBhgu8umcbmxImk9UkMsMPkdUZ5c/AVJUt2ArlyroXeZyoEMVrSuakSSDdPw52/N9DNajSXSQztX
qQ6yYpNKW9MHA5/IFwomI5M1i1QMuQRaE1qO/dEQOXGNeDaMOq5BEXwMZnFStSGeN8OEDaevoLWC
jFw0qN6TRlrlzgTCaM13VP1p7zWhdHbjsjR1+Kt7fMtjCTJCrNjT2viiFgsyEe7TLqSjFLypNUdj
LlUSpp+DouRQvcGoXLtD7ma562c0Wga6qjotSp8LAEED042dOUo5H653GkF9ET1FeKu+cd/jGXK9
1vH5M+qXLk6MHErtcBMAdriCu6GBfMvgiOQXQUdnu/rYaYavtL/oiRF4TkHsYBxc7gMpp8jQ6Mmc
x4ssUP3dqclHK6aMhIAUcu5zbRKmBF7pZ4MltBmci6L1w13+xqxzzJi9gu5GS5oFTXOIoA1XPzS0
O7EYADZo9jpO3iZzjbbDNozLZeLOwRaN/ZNMyzKttwIMQWQLh0rvvkumJmGP9neoEYlU4IcTPxl8
XI151+ApMsalliuTR29ylEaOB89PMvqAGzGl+oKoS33JUopbzbvaB+urLrjsdzKEKAFZ6fp2OUhs
etzszyDCTn53Iw1ASuh3ZbwAxMeRapnG0iIjpjZ5G+JsjH6ZgpK66VeWc5wKUrq+FkhGg+wOWSed
J44Re/cSVzNcgFThowbtZqLoRpXcTYdRnBvpE3W9/Kddq3vHJfGYt3qze44I59TQealPxp5cKSXo
6kMmEmSyDHSVLYLSv6+CCzj4PxImLrCuiALVtUa3YBaCMQyFX4K37gWLWjh92G/esbKN5e0n90aJ
pjXEDpcQe4+hFSZsnb3Y+Lm17FBA2pfiiNbSsbRlu3Q3l13Ucvm95L17zhsdNkLEhDDaI9enHdWs
E/ML1y7n5+xvRykrOfMBBuY4AkC/aL/IufDoH0h4OwMwtabGIjzph8rnADSAW7gC0D/zEFNcYMbv
Hl5peW4GPVSfMib5qx67V6nwTqGOqMVc1P+Wb5p4kTylnFNvs9a0MggNQywOndynw8BOj9JVq7dr
ldOYSUt30s341pIu3VWq7HS4Btm+1GwCb62Y4pNctp94WIBshC9FbCNPHDDWMHXX0+dkHp7F/j6u
st5HTJmocyLv38EdClqYo6QRlkdrCmYixT3iTBmz8oRdWZY2ZWBBfeJuz15zsNMlUlYmdkHRIV0n
Gehj0/KJj4+x1i6vT5dCPvJMRq6nO7AqJrJQiY7Mil3vresi/dpfRwgREd3BohNBOLHW8OMer+9s
MHIud6rYnM8D1c/8ekSJEI8i4W9U2s0MEvp8Liaq7MZnYlxOlMCWUttdqbxaU5uHt6Qp4e7sAGg2
qcy+rMEBqY8UkrARBAApxo4V0LKTslg7yybPtoqBAszyuX8oViJTsdXllEUbXL2713be1GChznSe
V5IprQDnfGa5sXGFSztuIG/u604hNitjCQ5RwWVIlea6+GynN/dr+/+Jf8ltgVE8fJW+tZQLzNIg
ZXIdNS72R9/8l9gNMKOLm3JO/N3E5BQsNQcklLbPVvTnbR3zBNR0M4iaxC17sFUwFVCYHOf8UFC1
RqU6A3i96u9AdR1D7BFIJ/ekBL/Rj3iqY/sGFifTYwUyilmXRm/moWIs7OuNHowA8a9YPURTa7NC
nvIVTc2pW57cDWfH3EjLKGFaQfR+6B4Xtrq/VIe9Ckf2S9TQXv2ftg8FktPj8D3EGEJOkN06kYn7
5ay1tPQYXXKuu1I2IWYdT3+Orrb+E27D99572H/Rez/sc8Ekd2hPiAw9fnDP3SoPs7G6fRsftRs9
2Ijl64BpXoj+NqFAwTyjJpUdwIMuwjCnSVdGmYyclU8vL679Gr6yjhnb17Dr/QLSbraCgjoT+8bE
gMpE5MVa94aH8kYYgy6E+L5mukupV8+ZvOVoYeJLC+AAC5hAfnifJMHqibtQGukg/r44ALQsArrQ
taXFldTPmABe0nxDhxnWGNvC7BsJPLGDJExZcFy5uXzYlzvgeEAXqFVIFzzEcZBPv6XAPeI50vPu
KDwqZPlto7JJZ5/8OAUuPygMlR8KEJle1AWmtSlp3VfyDfb4nYP9lbkE/3VT1YdqL2UjjSZhqpJ2
35YWyjfBByUtIP0bl5FRwSw3TPUijyp/xqGwBAGPrtyNZs3/V6ywOL1o+4y72dvHkyboaz1PBkP7
nfgvSnu7rEMeh2gDniLTy2duIU7QJ0soRS0IVFKIp+BeVvWqxeEJDzzvlTASOSmIEQoQJONSsCez
aLzo0gsT1cg9hQ4BTt5ckCAgbTs8VTsuGNPaen0w/Db+NEs0nrb0SgjT0CB0gKCi0eWZMM91GCRS
YnyrYD5Mv6hCETQ5nWppNUQpfEE3GPRh/OATXbbG4/xn5mQM26h78UNazfalcrdvjC3eT5wu1Zyp
U9BeDP7ECRIlSWegJ3oWBPM1FyaddYrgXs5furKrNOoIZ/6ktT8FahOXQnDNQxHKc6t8y47gmpy2
UFeuKPAU5l8tokQZVt+rAj5SeMjv713yIV/LaVxkYLSsVVQfw3fEDG97v59ZRnQ2kJxx1zQ7Gfb1
M965Gw0mn80eoTKDkL6HQEBdBT4v+/TliZTVloOW4WlVXlazoak+J2QWh2LphuByNRgH0hGspCPr
z+9WCLZAhU2o0Qv5vNT0DK1cwI9Q5Ber2HKkhLHdmvEhNvVg1k+tc1nIZATpdrLtmPosBnWgadQX
DTBpSLs1G8W+rbTmmOJBFcwQ6VXK04P1cT6X/ocBtPgCzHEVWRk5YAVTGwvv8rSJ8i4BMwmaU796
oNTYws1psO01O63nqhcLawOgwtKvB5tnEmJiThhupqnk7zty+g8XFgFlzJCBC/2HXc50runXzu6U
rECFxweAI1MO4SG1fjp6JrqX83fTgcM5bh9/FuoT0tP0Wn0Ec7aJuTHGuem0JSQqPUQ6HxrD4uvx
Y8FnlrFaaXghkatuaYiVLuj+cDSlnbeFohFy4orHVmO1bPMID0cQpeuRVE7MCZw4lJQGMxMO/jPi
X1OenkJpT/G5fkybYQ6dQcOJvP8hflggRQnmaBubHPzjb4MMIlLIxo2/jcLetb1vecjqn1IbGTSV
idwP8ew4gpG3jTm+roKzfqiuM6po9moUv8X5yDEQKWqDhfFj2oFr9XlOKIUb54Duj06x/Phzc5ia
Axbka83IGb0HLc2vc8X3e1h3/qATXKG5almW7Gq7T3byNVVgE5Z7KMi56jjamT5OsNr1NJX4cpWZ
QeA1FEGsxViaf4xG2vU11wyYyHHAMXQAect49LbzwgOI4JHHg3YL8/i8EZas08WVM7KAzaOjsoUh
36N0z4bhhIs+NEa7/Qii2NhdclDi4TyqLo/AV2qy5s4zTiKC2mKZrzPwl+3zkceRvgUXxmet9Hru
f8RA5UJF326IEyQdx7waUbL8dh43o1PYsT2a5H6VmgUOfW5iscVHCVhVUhqBlsN7OJY93Xnl7PRp
hERLoel96SFkM2wFeWFJC1zMatWFmo0n13NZxxaMcGN8ijypzx+cItouJVm2qdfm5LyYYgI7cMiY
OIBeCfTFyzu1HeFdu46kMmYw0mWp2R3Lgx2Knbs5GWMD40LK6VJ8meOnScNyRIKVLSX9Jo429tG/
f1S5QxnDoKHPVoSvctIcE4h6fVwDVwTKiICbjrsolgdNJec0K8gKY2CM7pAp04Ceu9BUh7qDTggu
7F4VzxYN6uzxE/5xP44G46Kmig7O1f7IJW0oAWMyjmy9OXph+eJp0Jy3OcNGzfo2nQZT3fma50HH
ejfFUZsIq83/qQkTv9+XMSzrRQpZNtYyrc2GZoTyiMaQ8K1daYQ+7ThAIUSkKOEpNntNFSpXa2cH
BAOm41sUoZ4yw2WU20nIAAoifTuZa2Reftdg7UhSKOAX29xmxFcTUp2anf4tkW9/F6I3eqwceP08
l+EWUR8vJvDoFMgyz0fJZozEspo1vCk/MIBo2NtLePYdziMxzP1nw62d/54bkxr5BIg0qIWgE2/X
BhoReil19hAvryEihE4g88pd7JlWDEI7f/NwZg36dRUEm5DvM9kIbqUXNTnU3f24lVfP7h8NJeq3
HYWo3ys2KGLpUkivjYWwRfP2BBaJmv/B+kdg6TyZzOF+18xCumHqjVlNL4H61fckEbuc0amuh3tA
d/p658+MNMyC50iINmV3DTlm1/jasNCxJYzWD6KYIQRBwO7CD6VenvHP5Cz5l4IQBF8dBwcl1e3Z
dbfb2rBkMLYwrVXEZJuY7EPEy30ghzYukhQ9afY4NMTmrgRjVch2dDjE+C79fSJSFpkyCCmnxsgS
DMNFSl1zmhj9n9jDuAGRyDGkPk/9C5e1R5CqYyRMPwEh9cAWIfIWM0rTMYQnHzu7uoeK1DYtxEfi
lal2mVUaT2j1AYgG5qyHmum5ttgGZxzz8yx21HAGr71dPPUQew6INY98VeQA+BEIkpxwQIUaFDx9
uIRitZ4Rt/1ybCbcezBoQhzkIi4FjhbBJSeznGZxPcS67m3kkNNDQGPA4Y0FqIWqgfDYx0C/1T1i
w+HfJzLxA2jS8pf7MnjPRM+hgrAnW/Wq/e/ALV4vPSU+vL16GgKSAexU/wPZzfCu/m3f23bFmVg6
MGxWBdSli+5lXClNB/qmtbQZ6aeAREp9MV5tQZtn45x2U8WLXf/6rNmXJfOR0MppXHH7vpgE2duW
RAbUJANnEZ/iJXN9EZIa97Y9MhcPLlD2tQxLhWo1JuTo+bYsSy6WA784XFZi9jdjy515vmIGQi/E
mEeKAZFr0MGC2NDtWCrkUKDu850KivVYebW4LfFJNNeus1hmzZSaBiUInnulZNidLcad/gjKM/A0
jzzP8vYIJ6nNbLeCsGFAOCZkHuFyMTzA8kEt0JM4TGr7wQp+SYVjrmPCb9k/jy79raEuabMqWZmd
IZq0ZYv441dtnCjD6mPl3Exbpwey25e4LuzcYbUx076s0siD5Jyfyslrd2zcFPLNBMRWfKx0xjne
ZS9qZRYFOxWENgPv+taeuSszO3JqRT2pxwwBmB87I2sAGQyGOLB6/Ah2LSSNDwGZnHg2ZU07VC6d
A6t4dSqShYUcsyKmX2NtP4zO1Z7LXU4304afgZCKht6VLoNxpkVT4W0lAkDsPDLr1hVLdWVWAlU7
hQ5ebRnffERljuk+KkWrN1e1alG4WHh8k7eGWg3URtjWDmJsjB61rosaYHEZERsXXfseRU3Fyf1/
+fbODzUDOqERcLUPFJ6ySvli66lBD60Fck+gCqfePlRJjZjAhcTTe+/aWZ6qLm/cUW1T7QTAwwFC
P+nOHAMfhgI+CA6oTl0gR0/mkiGcM1UY2VfET2Ess6Nbz2YFOKKNgohY1zTO5UpCu6ReciCVuIQp
SQan+MM0+pcakjV/whtiEI+rALRvzfDfRiEBF8qSb6KoSYA06PBLQxs/DuojAQIndNIcJ6PvtkCU
FfSILlpNQhZE753ifhNsgLsPPjV8g8pSQHz3iULeNTEeLZpTiRcoROMKZAXtlRtgFiywpd0Yb7ji
Z/Stis/Govdj9i821jcqDM8yFLTejfWjbeHUOCOZPe65bohsFkGtvKjnNpV1fF+TslLxXOUKcDYq
UPESj11pNC70d0OObGMiLN4rRus3KjO4Xy740uOEXRlTONtbaCqd73+Zp6oC1ZH57w2s9GU3ax1N
onCGip4HnwY8tQkzkVviM8/82ZwNcFtY3ffbfTtTQgo/7nOwT05h9Jhx/J8i5mr0XapYn+0u7oU5
zG85MAXl6qwHO1iupOXEP3bm+XqSgleyp37bmco1pXWed+fi1M1jKsy3kGD7doANXjgOz2ykGP//
La/fL7G4vIvw0Hf5o3M/5IABFr1jzAhqvagP85YZXiubG+XaZRWh3nM3D7XmAQOnQUSXC5kQGgnW
EviSIbzh4vP8AtWsyWvSO2no2ZGjAL/+1gQUwMMAvUJizvRn3HgRq5aiayl4IHgcuyTylPeeke8r
D50bIleHCQYEn4WsMyRqJjt9z9cxVIR/UB+zIrUVD5guY9+08abjiw2kjJz6ZstRYdqjHXggPpmw
xoDyF5Cj8lFge065bq5OJ6Hl+YlMA5/8O4mnsrW24JJfIPQ/kBOyoq76ffcgpbGfUwkerYytgDte
IilR1wURx2tFDeNFcIBwWGMK2JHE+aPbIVFkorltIwJwQmH+1GhfdTKcPUKpMC6fu6TdgaJcjqfi
NRwbzm50v/wF1UC0mJh+BnpNkVd/rS9uBu1jGTVZ3LJcIXu4uHLq+sG+0J5NR2kFM8ma4Ng/rQZo
Wyeo2kBr9RrtxGPOvTj1s5eUIbMjA7CC+sYH274FRlZaACJ96ezkkpgdMsftqtivaLI0xnqdN9O1
Fh45NaQMM3gRiN4PelmX8VNNxE0/X2b8a9u45Fjg3+EE+BV0Cx0wWlWMNzfVHaLTloZf6RXeR4ux
NEMX8Y8Nr45z89Oa1JBca1TvqtAmxzc2qFUZfKSpuzauR6F9lzGqEnbO6yI5+yn2fAkdzPSbMAtG
5Pfacv3U7HCfh3fs+5FEVwr5hWP8BmZ6QywrxVtDOPhnfNwjsqO4bhxGfoE5cylZqlGurxlcPpqN
xNDBqZAnsWxCC7cMIKgZXHgapORakc6a7fT1PwVr5++QBni1bcchkj3OCoDJQNpoQe5G9iNdAZ6L
PHysJxzv44MLdL7DJaz+FpoNPPFcnnYMkNXvZ7x8NuLFt3IUsTalGlAeONPh7ipetOW0wtSOJbP6
dGwaE5JulAXFKTd7LJ+IYC6FQqzTsiniHQpsVUS6b+4/HBHwh1AGFIeKHA6kmskeELFiCSR0Xa5j
BGhCYKhL8MdMQ0q17PE4m9umjcXy9EuRmj3jI2LsMXnBVs9C3j2Rn+JwBRkusykRKKjB9lCb/JQn
VNUIeKzucZIaTSd5g2PTUtX4FT5Gl8kJWPspAsUknoijKOl+/natx/4hY8QNIoWYhUTrEMk6fFgE
a+tRMfSWBV2ZALoPcxLvVOp1O8SuD2VaJ3xZCZ1fZVdiwBVeQe2Yzthw0cY2h7t/CT3+IOig2+Xe
JR7tjIbPBHgu9XRPtTEm0bcjL3uw5LzUJLKbyYJYk2wkRrR/L6v3Zu3cxoRWJOfsbz00A0wXcV00
OnhmaFIwPoTBo5aMyPlzaWIgERW9PevxsqYksqti1pse6YC4811pZGJzWiXt25tU8gb+lCUKE2kO
vCPLN//hKByae8nJUH3BUDm2LTZBm6QM+70e+QJrHZ7bEqtfivgWgaUKHzXvx/Rg0Mzx3Cl8KVDj
Dz8flmZCCpRJM9v1qV+SVUaRpCla4TdAXZWdWLzAzJQN8lsb27mHXbrX4H8CgCpbC2XlAsOHAqFE
JPSsz0/jKlUOHmKGrE43aPkVCvcIq9QKNdU9xHwYxRYzT9uqXaayjag1Bh7PjmdG/HiTOxM4ozQU
Gun51Y0nSV4HQlMYAmNND0zg2vvJJvWY88INyEkRrVhvnJ6siBR7hmn2B2oNWZuIhO1e6ZcsQcfY
6okN6ucQIFE8c9UpvkZp6KIIV7mxS48cmN2M9834qEpsjvN162AV6t9kvZrOPuUQECpH/ykXcFhh
DxFG5uJP5MFTjA4Nt8eWSo8UrgkeJ/mMsEpGCIKFqYWiQFphfacdVTDb/J4eOQRlLA1JjNugqsol
fgVrSst/PfHjM5EKznU9Okzl4WF40pJGgfoZ+AJDdbwDdxC4Fv7nvli3A1Pc6xsiAuMpu1a4/Sxi
fOPBpeGe3OwxVv/avK9u6Syhokjz3dYLKfSSxprS6CvSPeYX7QB34UOczryn5AuSxIyC7xGY65St
QDkSGIrUxiwc+Ii9dqSENWNWu8x1acwTPeHzayQz1QtaiSBFkZ/7TVi4Ag1HbJmzl3ikaazufVEa
gVaqIvFq6W1+FvOlw/CP5mRyGlFMQDQt852cCvRYMXSw7JlM6pKKalB3nRY1/K6nyTbi6qq6Ub5N
EqkNL14ttovSB9G/heedm6dpxgjnEz8LvWDM9RXcQfh0byrlW2aJCTL/jOE77lWREFVd556Z2LoN
ZZTTZ+4UcdrpjY8Cy/0VNAGTuhuFUqN5Ew5VydAelJOaUaDY8Fh690trd3BJWZhAg9Je1lcHyeTE
PVSQjBWpqZRj+yZ12MYzV4toHHiYmmN0rhDzvRDN6fuw6juc6ISPEDk8cPgmfuQP1o49R+WgGvnW
n/onTmINiSpPUwI7XA2wCkrEoTGFXJTO768acV/cjdcgkKe2nR5BbF2T2xDvxR29C2q97OTZbeJy
eeiyr5zDeHCSnnz08bdTnxc15asbrBO1SiA18v3wWdVhQvLR/w8+7X7LQrx1JQAqWjxOJ0dLLRQF
BI3CkvWYFvlEb+a+6gSrRszGEszLCDILXn8P2Aa/b2IaJTw6Fd30VqU6bLLjbgCHlZ1gsTBH5kxo
P6yHctO4mkg8Bhi5gDUVASxPuOUd7Rhrmiat2rKsUlbTuVM2/6S/uoABFcjNP98r1vQYOom42njc
L0wuJKCJtjaPgZTxiGF3xJF4b61zE3oqY7noV53v8sGba0AMao6xO1jf8ZbV3QzL9xCyvoV7g+8w
gu8Vw1RTutZ3DhVj8NwsDHn1H5sZdOnvz901pabWoR9AaVz6hdXRMl258KnwheoTKYyThzMTznL9
EoecB2RyLJal6k1ONzYPjtIFrki9JlHcoe1l6dIoCKnecJSffEkMQ7BKFadEvdtgkO/xbRJ8Ge8v
1Zjrka3Umpt0g6vQXsZ8F94xyy1cBqV8pFXeS6lHfCWEFpHAqcV2/E7YYe8thghCnvxsqNcRranY
Q5nimiG7k0+XAXHoCQ7NvaMw3zVZQK5WqLs4RqXeVFGTtkBdKGog1NwaQMTKUuJ0RdbGNIAesQAo
5KIlwSdJpTHIJeL1B9ZKyLKlliEK3YeDab5RqrHwqnjHO3nFaRjknRKJg1U1pVIB9wYJFpqdTVI6
DOOD7Hbf4Ab8V8xMmPQO6E6GfJcT4QYv6L/lZDJBamJHrAC4dz0qAj9WUxPZ3CfTQuNO4vruVfNU
xzeYlBrtih3oXyOzWiVg2FO56GVb52txjBkXAeD7jJms8Wc6sTU8+hftyV0MpqNsjdZByRZoY6bw
QW1/r4wg3ANS/Bi8TxTzjK30Y1QDcmkp031NyLNwstjUFLI3Xdv3986eNPbLJqAoHjziKwxfdydd
gHK7BD68c9eER93RNvRV3Oz0+xROxK35nehTDO2P6qgO7Olng6wL5k1V1NT5vXLb9EmN6hs7/Vio
DtXv+FPQbuYPn7XVcMYtKs5U2o06MkD68BznfDI71Gc7ide45GbpSJVw6gzUUs82CixtVB4Uzt+b
9DhjdJHvcbahsBJ5hK7/uJe/zHz7U+/mhWHZiua3HnUlbFQoZ+aDp5NnP4G1Wh9nibYraiXcdQSd
mskml4L28KzxbrbMVCFBpZaDLKUKdXGUTStuZ0lByT8lHp4ERzzSBE2YwoCq5L0CpV+IQzigq1ge
944WigsSX+YKKJzJjmYCixWAFaSmkPdZJ8Kp5vQqu8rp5pIXKG4imiK5laeKWhj5+P/+J0xLuo23
1Z1YoPZg5Vcz9G7vYANSBIjmpx7ME/Z4C6eZHqcccwDCnZlqvrGZeZxd2k1poxcIXuRPn6kCFhn8
W1YmvUfwhBJPhXHSQccZhOyTjPnUhU1O7R31iallAkWc/0PeD4c762Q9ZA9xGbz91Yvc+q6k7aIu
Tyn/1GhmB9cx8Kbg5DfLOSLc2Tg0e8BVEUPauLm8sVoET+kYqcJQe0+HLx6R/YOTtVFxPpSiMV0V
+d8YjUiqgZFxbUNOmq11/uuyT+jrTOtfPQ8xGSTs6//Kh+Z0SuAFq2RLpBdrxuyIis5uZroLk1zo
FQVrOIDXj7Gq/m+DfrnGUX4DZE3/3TCcQhK1bHjULFdMC7zMISQX0b8Ud97lGVXBwvksIlGzj5lo
9KvOYkgElX5n82eDT3K68jBPFdz3+2kSMuHGvSoTQOeXLv8PQsT5Y5Mm/pHhGzLLhwX5X1DbKLzC
QwGGg4s0h8iNfs/Llqt29hVQrAHDDqbd6nV1Hv3ke1Er24OpVM/0a0va+urMrvjfRnte3r5FlDFg
2MD1tvBa/bXRUtV5YsKxZGfxBMhrUF8XBGRKdUbuHdD/DMpjNFecBM89j7gBLshNcy+XseC1mOaV
qLZZ7zF5gyuUtTTmbS/Fislhe26M31Z4arKkXYP1Bzfzn8TjWkEy2pdSRMVWiVxepckRePfAOXBz
ApVfBI3V/1H6ubLM//caRirBSuP8HsiqhvcZEcX3a6ribDYF7UGd+DmTV/58bFXg5cdmQABP/wAX
VDl2fpSLByveMRbkKRvopqmjCNcNzhWtz2cxE7nt15OFKWfju4e1m0loO98/Wz8YmaCFWYsBiQrk
UGlYBxKCbmHKyZrw8gXepiyLf+MOXT87zKnLtUslK5Z4qP8Pr1ZbHm5/ogyEfXJeqmSw8k8j4ish
76MJDEkZCz0lR6l0E6C+qJsUBpgD1LgEhGtTGlSlvM4Jg8eLeLGbMH8pfbNMGcfQwqGOH6zgOWuF
LKLjkMVG1wFb8exQcRbUmDYbmQmk0Q55DW2qR5EbC9ka8fvGkGE/su+Z5e2ALMTxijEAtKtrfB5v
YtK5YuIPlzQ1y7aWLYG/zwYkIhjb75mRAUJdOHpR9BiOdZ0fn4T9mtzL0dlDbE9SJkBiSFmWv3Vo
VhFL2kWRddnqe/dkNI97LDXw7A3UVZhRy9W12hiFzh9PEM+w41t2Z+YT/7ay0o51F9FiX9ZSk0+P
5lJ7mwFybFp9420YGcc6QAZoGPymiPGiK05XysdjC0o/9nyqUn/ZlH89DnFtOnBF6SWKIEnaaoh6
111smRapQiCcH5r5g0TYhyzAm0+CdyrQTCLUsHOWWd2CJt5MR/fWdvy2m8Cj8rHLPq2kXl488BRf
PqEYTEJjN5oxA0bFdt+bVZxy8BWK4RvnEwXCpB9ck7aqTns1WUGXcXvdYqpbMrksWleuL0eBQMe+
o2+kV1i2Fv5mIQB10iaH+cSjV38wMSKum5uqHYRAyzSENFofk32n5b9XQMbzxw/NdYjKRdGq7Weo
w4T37leRIuuMYz4qIlD5EBextYgUPQYXGReWpeI1Huw72Mrmavg347LylKa9L6oBJJBsuTeLSJ8T
SUyXxSXitdvku4jdLcmIUFkR7KYwbAs6Nvy/m1TQNA88WcLgMMoFe1JTRrEZCp+22lr/b9oWKhsw
gUWmQmLrghGWq4msIcqplDZVfWDBPNoRG9LJjYz+oiEJ9yrGH7ErjajPemCEJyg+x6+jKLWQYocZ
IYMFqbmuTumKi7SoZkXH+3WIsdN7pdqEW1T7DflD3J2dSs/e45X0zmnVf0qNeOJ1n85zVVq/hCEE
oDafUtsUiIQcDP3/3xI+Cjl+G9ozhSXDLo5Kd0ZbY7oaBJdmi2klJq5O1XvuAgB+i7YUTB+jty0b
9FA4E4yCevO2anwEIJWidn/I8Bh0oDnzdRFlEZ+5tEyip0JTCnXk/L5NlQ7Cwu3OM42YdHpwKn3S
e+HYNDUWYAgJTOFooxdQcVznrxdidt0q6Bp18Yw1zt/kbJd+actlvByBZuB3tmnOWbh/RQ6ZXika
nRqr7/y7a3Ua5JMdQXju9Hka1ydOJdeOJycZBUUXVEBfNIU9AydsUNTnEIuI+rVeaoTJu60SPAHp
53unHywjoxr/pfsrA5s11aNwwIdD/QMulKjqdJX9lKlcetqe5H7wIStcmqNlIIjtc1NE+sHiCCkx
qR+zqRYqR6vRUPTvmbkpvUiD6nuJDExLKD3nefnRMgOPw0biDoDz2Ox1ZXY3ugM9od+/TAHqWuat
/cAyrDH/hnL2ammnMAtx62NEpAE4hsYLrowXJs0aqoQ5IyuApbI+qNXd4OijIAxB6l6XltWPROIV
K9Ha8zMlU9IqD6nSOi4gBYZ+9TVCVp1zkdwadZkEyh/lVhMITbiD7FnVcniloJGvXFx8ff5y6PZ+
bw3FwI0JSD4kMLNYeyYorDF21NtCnsb0o67dni0t2mEvpoTxVg3hSAfgFjjNXBA2T6uOr1qwO+OE
hxvqgvNT9zrvGg7zO8SI0wxVrVnAbOm2hBcTqkCesd4OMJtGfEXq8XPTutDPHTjhMyrDriloCZeM
mZ7dCpyL+hctIY79pB5Mgk2YYXKLsqVRjPGmNkw/gTLV4cPgdq4xX/F5+5MjxRxw4cEHVwAmmUKX
dL7VmP5GEwoVLEZgN6vOO+X/+eaPb5G4YHlJGaPsXgGowsTFgGE9CLCpMtI8thuCO1M0ESo0IO5c
pajVQOKX5i+pKPK9PyBSzjDpTYtiLt2hSMb2yII8QSHuEjP1hp7GOQXEbxZIRtnDJaHAB5u4X6YD
4LbnDY/gMLkDqqhC/WYcyPkqjxYAFvI4G3T0g9H4HOqUq+zwYhn3TJrywVDMLw7QpYVnO2q0D7CI
WM90F850FbGQ/C14EalIdRJ9ZETI5RJNMHpZ4vAusPEmS1w4LHanlJXNgyY7hvd1rvcCQui65Atw
xNUJ/UL3FXanAV8wA91ZGGJfP6Us/Sp1fikQySm+ggn0ygcGFLAeFNuujo04fekJPIbZz+qIBfOB
m9LPR741LjhR24d8pFKnRAYekk7y4MNUAZdcx64oaV5S8HRi+oEa0MgG6p0JUuVBWzV9EVGhiv+B
KTLQwhSrcybXUeiOUokYzpygdDIbYpkEyLj2GlwYKKhz3Rg3gO5/oVysIOLJ1M6tJK4yCHCk2uBn
pFp1Vm7VVVfidmXn4jcuflMy3f0TTvbfmMzCDyMnrVtwan5y49r7e3ybpUo0wHFJtWFo9gmE0jpI
4wddmc0LKQEzvN0bnQWPsvg18op7Dpnq0mMNtmJ+8MgNwyfYrY5yAuKHk2zwhZiBm6RwhG10esUc
L78Vtc6LgFPH7ihNyHk85/aAvKNr9cur/HRuGVpISDr7Zmer47eK9N/54eBmFBkFLuCew3YVgrlo
I9Bcr/5gg1SU2cOMk00DaxcTNDShHFO/M0rcYjoKMzSWHO5ETH8PJHqF7ArsvWLZjFVgVaIYKx6o
eGu5U9NShOA2EsRQV1PgsRzJb10oR1aRkWZcu8Y7PzEpahOMXoV4oPBNJ7zSB5by6ctsYNy9TjhO
VjtBCjz2sCxpVkpXoc1MpF0c+yXxP14OsrfWMnexaz17OhcHyyzXJGnN353ryxNR5icHPx/48HG7
PfH8car3MC2woxgF8FLsWUAyZ0injynHzvEGaRBQ0xVJw88iqtvF6FCfjxRpaMoMM9qPil0Uqkd5
Da1KDNSBsZm3DI/O3Zae7BjmR6tm7SJngRwWpH2VIME62YW+mKbsRbrmcQDcrALZJKnZFK/mU2xP
kYhzHdMXemzTeAp5Bw9fNp2Gkm42ydtvzmhTJLuKSeBNbdUZs9iZ1QFGedbNe49g+4KUdKcyhVpp
MrZsmojG0mWReb8idHB1D7Wmsyo6mxOBP0W57gXZB/aXDieT3xYP/35/gU49+X8O5v6eUfjm9UJF
EKNKnI/AJiPa0mQKlECAG8W2bQ4FFCAaUIoakAA+d7icNN2aNDw5lC/hj9FrOUWaHsvVHlKFkBAS
BbOiw+E6CJd8FXTYJbvyuPuSBIncs9MDB4vYwBzDuuGLm9Ec6LjEXXx+kemk7i9AL4utaA+XFoU0
ks6DZROFF0ylhNpqSuauswwf2IfmKgl9VGa6MYK5eMXuJoLxY2xh0bevdBHaXeHA1qg25e+pJkHk
+0NYC76HxG1IgHNyXel9Ttl0KDV++gDJUmEXF0sKTnObbKWhddOnmgt13qhSMJXIrSWKJ5IxkxTn
7hZL8AU2et5pZ+zwb61712b++Xv7e7IxVEMpSSINKp7OchP8ftJk95a3vgzirGsxW6daWQ8LdfEr
5IOYRr19/UiNG+m4ANG6yeumOw8mNXZVEfWuxllZrVG1qfH8a5uBEDJWVSg1RAYqwTBnppyNF6g8
NMZEmrMQRP+cdzyLMYhF56mWVbYSzQO4jXN+Wx/Bg8CXMYWhUNhHWS1GlCCoWn4jwpAkMmL7XKSh
3S52RdwZFnnDluk5tLCSpWEuDw7bl31KaiDHqKJitADXqH9CyEYYsDm9wP2286lNuV7bQvSgV05K
wQkUelx/VQ5gqaG+URG5Fc3lywWI4comSb8bSWkwwysMhmpmZljcKH2iAPl5O3cdSRPIljj0b5l0
NSaH4sgaYT1zuEj+mITerzX8Hnl6YSiFplkhMoWiQ14DQLeKrQ8aFl+fbnNYeMThcCG6ABBXBIBc
VfgWPkSTmzI2qQvy7AzQ0U/pbWDBDGSxO2XuT6yYnTiKa/KLXUfdxqaX1lDCI9T8aGQdhL8oXlul
dZvpmSfBvQRuL81A/gPhfg/NQ8zKotGayEq7zGtZCwVdEDx5Ia63gK2xnQiLcyIP57YtIPPrKrtz
+OEZMuSPe5oFwG0S4rVpyVrryl989hBzKQK/v94JS1grIo67TEoiEyd/AkUwO+xLvIspWXVrkXHK
1sP+hVOzjryib9XWPmgR/5rWLqcUOTm0TQjYehvdsvqUPor1v2y5plZsSyerITMZDkFiQGfilIQ1
CpfQFmAcWThCYhgFdf2AvCqx3CklDLvLY6zHDAFjp+FPnAELFdUkqvUlWVgVY9+cQjuEufeJnL2f
kPZEBeN5zxWLHY9qITSgcQNun2rcyO68oThwHeLfpvptKUnTK4NL75TheMRM6VTqDodBpYypawBp
DG7yKi1ghc3LmPCCt3LR4upDEOF/8OcV56bfKD8xiDqOWFuN+9i4gU7DrxnHf0KCNzkokPKTlm1M
wG5mQFmoeu1DI+LXtw0JvY6VH96tkWDIRWj64XRGLtN1DobDRqzNkeMqJ+PYlfWdBYnLazm5UTmh
7WndnuL+5C/Oa4S3RC/2SAeltZSv3EAS4QwP2nWtso3FEI3Vqs+9hB9Ja4ywImcYPOq2YrT10TLA
rgAtpi/6htkeM4ADzI/vkWlrQugf37Zo/lQh51QV7SVB3OenEeg2ihGC7Zf+m1b26VRJ4Br0yN5R
hrVV8T7PjvAGzt2Tle6zORh+O1hrQt5Z1/w/olCMELKa2cuUtdP2rRWhNWwZ12DPgyOexJ3xVSzs
45v9W/WWmDG+ufwfSJfan5AkpNBNkKrzsWpUvzjifNoPIY5tN51sWoKI1vMZqqGThGmQ9V11jolO
jfRpcFLAgi+Ryc+FrfK+8wpnbi1yMkQHbxh2+sQWZSuguRTU76TxGvVb3GR227ksl/bV4FBulcei
RmyV7p/OMDIYmTP06k5WsrFcqQ8Jg6RKN4CNagVUaKMWPathH8rkp7p2SsamFN9gQ1ISZCcjFMao
yuKxGH56GTlSt8MeUsGada9M/JqhedlYQ7SdcbgbQb954wjyVK+6aCvOqnkiYtYZ5temF+8sxt3N
jIKnLr/bTkiPQKLlq9aKVu/gZv4z23aTCzn3XNrKQtED7H29xMjMriEB5oTG/QOAwHrIsF47heRo
wKLRv37QqqdO5jTPAnPgc8ZHuZ1mDKzbu2CC6KLj3mY5gy+GP2RQb2hnkFaLtQr3iT+5Bk73AZOi
JEyZiUwOlFNOdgCTFc27pG7UF2pyA5Y5rTGXCdW76yYGz6fWmMB6sGFjP2cnjxRiyAw5IjxWkpPo
jlu3c1LKHDWqYEY/mZCSzUFBWSAMRyrPJN18DhCAJKv7t/yMDtLYwaUXqRaYxFhc8iCyQfzJdjsf
8URHxHcY7NuMdG9tyNs9olyF4+QYrwxh0+CwnZX+VyReC4daCGMMjuGbimztifkr6jHsUWy1s/Um
GPhvs5NedkpFTGavJOp6Ia60OG8TD5SuEdZVKiXsKwL8IWVbjA7RgsToAxO+n972iBVvCCP4ivCr
e+aIumjEgsKgTcYFvJd9zzNvAJGMuZscw7+o6dNiGZN/3rD/C9xt/xuI7gDU6Da5Gjecgr/iZbda
Mtib989EI69UjTsBzv4OUm23dyTo6sPoLhyEu4b79xbqH9jskJtHxqkNOH2cCyuvB04MXHbu8B36
oUWr1a7SiRPxOAO7VMTVSKsTzNGy04s+s/c7s/lBO5xGsckcZDOQ/uNxVSBoRRql1CO5Lii4M4CY
5mGnln4rvaMzDqyIdd8xpsiFBxQRhhbFfliUdSjz4DYuOU9CaoT4FRENtXYMvUrpIDfqh8O5BNUu
JXbFO2lxseAyzU1u6ArjmZokDd5EpYgOVWomSIZ6fg+HNbywSrYgRZT5S9fYisDAoropRB15lQgU
0afXhf3fOUfTyClqWkvV4CVZtQR0kzIgAB8PWxn0zDtEzPW8rDgHDgyBQGENFAZ3EWofeGZDRAvI
C+DSLvacIF41qVXZYHF7rB4/1xa5CBBQkQNsp/wKMOoOwBFYmhyB4UqBAPhbL3GtAjz7cQzz39dX
FnC482pgydTSIDzrM/rJ5KIB72N9V7tKX+VM7L0vuWhwNMAh1PpAoxK7oALlTZ7+QSPbcimkZX9Y
gnPNAEya5YvBh+vkokQ0MswhopeblrSKXAmPhroG6R/6Su8k4Qmf15lPXzmEqAi+HRzFbaZkhbyo
NtI2R0NUBZefQF9ZMkt26TMa7Xf2MK1zO77OJ2r3VziIEsMZnDXxEH+KePlvW0TnXCsrlZ5F584F
N35Bfj3YsdW9G3RnJA6lbWS38h0lPd6k/93ma1n/mAy4dRWhnN2erIcrkRNPdMdAe9pSF/zQ0vs5
Xo6RSiYPxy1v+YF5l8bi3lLQOMrExGYWQF521HkKMvsHdzfxCu+Kpn20djdkX+XNFTSa4uNPK9Mn
akUlBXeSCdOtah7RaN8lRelvrm6hpwChU5LX3qomvPaRYRKBIyglq0/NPNkerYRro4F8hn/1bVob
gvLQYJImP6dn1SJod6wmcQW8ItJCdYi1RdBadK21d3eXzYa9D00Zi9IHA/nFsiiMiQQtHlGVXEeV
w0EAT6sBTUSdVCmwP6qncZ+U6OAhijex1MW/kj/+GDCdsoPt79SU5wZLIbUR8kAWzsuSJWPO0coo
l9GYtGqrqAhyDgV0dyrJ5qgQ3cZ5/bBhfEI3isgTP1dAGZDG/NCJxXsxN3UpEaccWZk0w+V7VA5P
krA8c/0ucMHnEkEysc1o6vR+Hr9fUWbUxHGiJGrrTgWGhJu1ILsbFGUUPet/Od0L73ODx+LkK/gk
y1NHAqEWFLOxns30x6gLVWwXWjqaHBSiE00iN0cUQf1Bv3hIIjZoj/2n48jsfcYXm4RhFXnWXTr8
1vmWFpRJDayR+fqSARrRDcSTnfED7WnAomcLEej7IoPhqB4jsU/zxWtzZ1YN4O4xQ2drMf1sHUSE
wpRW82JGKPF2NL4SKTbmGvFevC2yH6zeHgSiTXAWdHBgs76ZZ5mCYMALj6Qekw1TEQ52LAcVh8h8
oDcAwLTjUGqssarVChh1PG7KsHtk87uvinO74Q2pITB8C94zFBNWDI9ZoM3kRT2+TAuo2N+xxegd
55NwoAMsbuJJ9zgeOUWVolxb55dIj0prpV7G1P1jEn1Xrbz9aWY1ochBDSl0VSbgaVvq4NikzELB
PmcXaWTbM/ZRkgtijQ8HbRbx4C/mMLk27LpsNj01LOqz8BU/nwq9TORuq7woY91Gan1/2S9WsxiS
8LODbob/cMtk7zykoRR3FwatWeI7zxPl1TmUuQIQYdFED0d0fNxF+Kvp7WqJJD/+W9z4dAsZ5sMk
ZgRFtNPcE/KegzNNqA2njUMvbKuKnQPBB3Sz1gzp1e9CJHuchueCB6k35rNEsIVcpnQnedTl2nfW
tPeI5IMQJczQ8aTrbQOb99YipOpDpNzZ6aDU9wGnqF3pMur0HsqlxQUR6YitVWZivL7jlRCrEXSt
danTr6hCr+eRyv5lHnhmEu7Bn9dZZxU=
`protect end_protected
