`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Ygz+5i4GtnsfewHUftwgzW1ws/nOQwNWDn5SBMtBThP+Dwbg9K7NyUsChvG8Rx+qTZXVyqlZPs9I
9nVG2ljk7mS/B4Gj5drqhZG7hbgavIxa6wUMAVCHbgIw27mCrpsWTDMQhma2VEql/QtfBBALLURG
3qC3+scS53jmByIICyoZ/Gvd2POrSEz8PuuDso2I+xEln6MwnjP/fFigxnglKZyX6NE7yqrZUC/k
jEsjpcHHwKACAFzvbt8Pz02v5iWI5AWX2OiLkEV/NvqlNrXlS+TC9c/+6nnZOtlfXQaX5E9Kd2CN
pOjm0I7Vc2ZDWTTMy3lKIPrbfN+USen1eESWnA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="AY4uR/IWotB/DE4iEqrqGOXjco5mc91eOeEdd/nHhTA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37200)
`protect data_block
UIQFI83oeCQ+w5qFR7m5vXuPkVj3v24WOPlDPr9V93x7ZZN0whi43w/RzMwy2pfIejaUwWOxt68U
D1denIMnBucquryWpoS1HAgzbky3L6DkMrpe69GcsI6Zy4ecKQZaXmsXt55dzY4EIM030HDtmKlM
/kwICXYoFPUPcygQ9eQucbdYXLlacEB+l1qejaYRY2RtMKdP+yvann69BbXZFhwfC154quxm1mOl
9f2ApV6UVhS+mgGdE6nCgLssbSeoHtZb0+fwgpI3Qpa35TC6lXArzcoepUm0oi20ySR+w3MEmsse
ZiKCkinsYUQmowewSkOofkxPXWr9jZC/6KFIGrmfa/ZXmVf/cufylHQDl+EIZty7XJcNlneLRWA8
VogdVkIhPHkkW+PZw0LnSOZLNypkRAoFfJSyJWgABSvTqwJY0D60wWzdYKHYtbjpFS9eyb9G6fay
4psqVIc7xE6fl0K+zyD4cj/qRQmlsfLq5Zwr1qhf2dZzG336C9CZr6P3+IPlE/CbZtbuOuPCuO5Q
wX4O3I7fK9qdfcm4xZRhJkXKH1TXXMC/qknIYYY3MHw/8kdSVLBbyhpksEGfaSp0kGlPi/NELZZO
+GUtRYvK3rQUcSLAxnMyXw6BOhjgmhZTK3pPAF433Ax31TqrG5vSidIZ/qIUdPk0zrOl5NXFgCDe
cH5vWnEMZO0ShxRVlyh+8DAoyNiN0OGvmmTBl/POslHb5M+5b03KnyJ0U/LMkUE74bFVXq51TpwS
a2gi/MCZWHyKKKiS2TF/6DYGjDG+D9L8TwNA61Pj1N+UDDV627bHEuLEL+OKu7MofxChL45E3FN8
tJwgcR52zwDa/5FEdzcmAPv6rXqHOIhMJEYUemukAXxQECaPTeNzkXMwr7/8DdrOFbZkruXj7YaI
mP/4N1vCJ1u7tK/oaRdxlketYt0lJuiapXZE5LI+fTpg4rzWEQtTWoEVToue9ZuIJp0zbsRrIMj6
vF7hW6X80Gg9fZAHt3wAj0GRTGF6qt9XZrI2fwtdkohj9WEH3olywOpX70Q08KhMI9YpiqWAvACQ
XVYV4o6p3uY6zquyhxH3cJ37QB0UJv7nlh6WNvzcW02aio8I+cIKozV6kdld21QGwwiDchbgBTOi
ruhRGaqimTXFuf9ojDXSr1r99MYloSCfzfyE6G8sMWoeRMtDZLIOBGMrLMthTYHvbOXk2KquSIL9
0ByL+CthKDfxobIpE2OP+VzWn1PSsRU5wwiUwQgXwWDjRDoEa41p21MiLWgz8tIYIQFewCVuzqO5
NquRYIf2BF9L/0V9zJEm9eiYHs1hv8BNeWJ90/JcH51kKH/ApoF93v2ErfWwmnqWEwGRZw8HZ0xB
3nwS2ifISjuvkKOqYdwd4Bv7tMzSrUFqD4CyOkKraKQnmY9LdGv0qJN4Mqbh4tKBLRgQJC0xjmqt
gb4sIDXW3mrrbKfte30uGtBI30mO50zCoS+nI2oU0TNT8Ctws1PPz1653DGBkQewTrnAIzZoFQwr
t1/DXbBSE77ncEDvHGmS1EZQJiv0d4hRIR7vxO9hfnv/GcxUoR5i4mpomZ7eUqCndo/UfxbiEktS
QnW7hFZiAlFA5grbGOkf+6pUgmLquvJ5x7QUdxQxwEL4x03frmE/cSal3XDx1+Fd0s/4kUIfLgwM
UisNTnNHSq7SFFMo3SWY/YtZeQgpB8BrkLqTraaCkPprO2sMWw3XVh/rM5wM5HLiq/5NsHxbTDV4
1HumAAdeyi9hGF6pXo51iQUjYL9iAcXR5lHTkfRku4PGclhgamr02mrkmYdlCLm7pdTrbuuZnNS9
7szv/FyRus0CAsaQJwsStZlD7ts+L0MtSutvBNfnMuID13lC4rlpImm7V9KlePVhU36P+28pmqO1
Yfh3aNVDYvGJUyvLfG/VFCJ8TQ5lL8jN7DCxyUK+y49Gs08lAcPQS7U7l8Jai23rbm4KETJcItMS
Y1WzfBIGlj1WNwXOADfBsOxdJIRpkFWzcxAmdoaqZSUSV3GAN4vwcrgHU+C+Pv6C28jCqNQn3In8
W93UKcvTKkE+6pwwXU94T8yIOhraWqtBIY0MfJX3fyP/zTUM/VHopE4RseM/4K7szjXGarGbrHOJ
wxSQ2RpoEruXLoZo6ESNzLAj+jhnRICqQz/08VQ5JFju3/a6fsQz+M+IXqWX7kqxGrTw1X4QIYgh
15CmmsOvhfwBqwVNW93UWH/BEFz2JgcYbpNQNK3L+X1jGc0nfsWpprxjGqCOfNGR66c6PndFLoxD
31v37e9jahsAu+Rc94pY1rq/ItxkaK/K4aqp8JUTA7Y4VJC7/9vHuWHIwFWr2/7OVnw5nL80CPBE
wCJZWthJLhyEHgMCTd648pNwTvVFO0t/8C3rZgn0zYK76n1VoeEPPAvgS1zcLXE138Noy1liyTBl
9eGvz+WZpIQoPL8nEzaPtkJK/PdG3G3G6MNTKd9+c+LWoKyXeGlVbgHpKAlUeRECnSGwrMlNIkyS
kqvA3OXaj3B6z7Y6TkzRpnCNaOTKgiihlU0Bt2gguiqbVZR3VgE3wjDQOLqns9bgLJjSv4bfvRrO
zDocnx/K0syPyY2lhwiceGNiCc7uDsDbrpWsEIHB/0EcFsYe+gemB7upE/0QMOms0drrrnzPSCxm
PuNk+szLO6IXwZ++Vh5grDgW1QYl3x1DuucVy6u+AFdont3ZA9WVFtlbeaqXRcl3zakpbzzzfgV9
hhx+bem/wOTGgcvyxKV81TKVzOpnXW7Cyo+dCrumUmVsRu9hac0WeFYgd4vtWWSgW5YliSl9Tlqe
yCLraMW8ERsmG/kQMcZdjV2uUru8CkP1EEjN6hITgruPCAuUWOh9HHu+hMmoLyh3jw394PghVrW3
P0Oqjdmlupf7BBDYi5XqN3xQnF60ctCC4Sh4EZv3H8iSe6zejzrApd+hir881R6Q/+dB2WZE+980
8WbW2VIkrHF0NayVge5aI4uvxCfHAtdFAYW191GHR/lpPXhd0+YhZs8ydmkW9fnxWIufIA6fkWfN
J0BWIhBMS89P5M5TYfBTPLgN+6ft8ysaf1/3mwwwW1++eZy8YG0kiaPJWUTubhDx89AQquhmCLqb
sd4IuzGn7OcpMLcT4DXPeQrR0GAXzeFHjjkPkZinpg5qg8K8yNVdLQJSjj9Dr5dBx3abSirvpAf0
xT/r/muPpn9DkIFq1uNUsMOl7pM46Hgm9HlrAmSh8Nq8NAU70B//2ydK8DaM/aWuGGUCTEM0Mo4K
5JZgoJex6sQIxJCeqdV1qnhLxRgzvgjX57tGsLbBQkbTwKlq2mDuczqCUsJsfKRJHhZHtFtLeVgx
iyLcJxj9pWx6hmKKWZ7RkSFMhMA+GaQktMlI1KVq26mAYkptejpk1poXlrvVP7dG5FyObJPszpLI
TrYCc/JQdiQRqkSnfHpYOxS8m3uUfD2sX2Mrt9nbHXZjghAdABBjhF/gFX1U/8efZS9Z2I+WlJ2O
g7xxqibZWfO4VagDKBLnRaitbgbImNqCguJF/hwySj3CZhGLJ/qCBzteXDjwOMU6PQI8Soe8wmZ3
jFH3D8zfkAO9EVR/HcdU08m5PIqU3dtLVHa/6+m4XWKHHBjTKy2RPt37jiYHKN9Izsdw/nnTCM4u
lpiEX0Cwxk3gSIm8WpnqLixecD/geXWoo51KFqkRgxDawH9Gsj1fKaFCTG0GvZg/Bj1z2XeDYkl5
5NHcgI6lJuCFirPBCUlj+3yg+zsDQsG85uHyANNrHQTyfu+FrYWL4JH0zsG5xOkkydVirnDPMKBT
h6pt/+YB5KhKg4Xem6eU071TKA/Jvrmjk7DHhQrdQxyvw8PB945a1jqKcpULautwZjsMs4ckLdBp
hjZ+eM+y47hVYTjHBukrgHNT9Ey8nVZSgNg5c7IPFLe0+yszTl6DVPomNuskGpvDQ2AeMhmjJqcM
IsErpA8CoL95edGYP+ipMBNccFn38PmEU/qvRBeXO0q0bJFdX1yXw0xEY1pG/2xxHmj0kEXskjVR
BD50iJh6ET0DveQD8gwSUjcqlRBHoHIK/2OmP6pf/6odVKZ0Z5aUt/BLwNOJOfpUvI+wmRVkWgVp
6g8SFxqZiWoJoQhCPEun+oyLvbiQ51PdQs6xh1tvVwABItU0HFfl+4akCB60vsSmev+YdqQVtxuq
EMDeb0qsnsoHJkgl94XWHFOdqUklnZuZsu3/OKtgyEx43Zd+SqYcotT6IZco6kqDSjEGGH0AEBRR
14mNez3H3sG0gVXL8mva2HYnKOPbcHqNz6nzpPeFmVU/ngg+z2z0JCH3P4hTD1afSCblrIHRPeXl
9A72nz5mA4XViuuy9fr2f1wwryjiumZ4Byd86wHBx3k8OLoRPmiyQRwRr+vyWiqZtobg450YX58F
mtFPjT3d6zrtt9wrqMYyMdl8fPmpoliPbpTtTXMMXBLII1EAPRBqg13fl3E3yFdkiBZlsdD73dd8
mnEb5oKJlbYucmNvZixDKubmw0mZHz9PKDFaI8DpoBfTyevromlCcmGrRjMfEOsDlBEg4u9fIa3q
j+3zduiPWFRr5m/LOxNjtPVbeLCuXowd7F+iNqo+hPXNecNDSKBr7yWdZkS5j4pwDxUKGOTaTHdW
GVq3tu1fC5+IpRDS8dNakeZ4qDczAnjvLsJ5GCPsgMypgdSbnXel0P8nn62ZF2vMp87KBbSF7Ec8
Q2M7HN+QBs7LHznFIP4O+mHnyIkQorXY+fhJDehLV35Y7sYnGgUSwDM888NK42r98I4q/fyRvkql
tbLaZ566h72dSVfbeM9DwfSktwj2q4yEJZZKZAtGo1GFD1oB0EPm5eN9ka2DWV1xjBiBBt7f6HP2
0vh3oITUDDgWWWV8ev8L7Fe7QsW5BoXaKOfCeURoZ3eZNv5j8BVs8Q2q0AMNoHrkCKbXliHRyng/
Lb+H9PWloMKJ9VSwL3Om/7uHRiz4ggeBjH6j/qWEMqJzGzNhOb8JVsiFPy6Pdt67m5BNBn0ds9+f
06AVrztMOhCflWqGPlKER1n7Ny3KaqpaCdGRoM+wLqL/HxoJF+VaRkgol3ihtUDIcyaa2nqB8i0D
FgCbDYrW9q143wFaN7cSkPIOdO2BUF+ZcNdGVFxC9nj64NdFAOqXwFl9v+wlaOPDY7ADBvb6GgFp
0g/SifoBYGhDT1zNto1HoqKZhp3Z8AvM4K+GmCAV0OBII9N7FkmAXEtYSxDhzWSDSFwYVHhOaBaN
Ohuw+TSOBy39+r+d2BQwxNTU+LPDqrJQY2gjaYx+vFt7f5vg7ZNlAAQkkmYCylcJ4bSOUuNpbBWq
yEOMe91nYap7klKBPgAB+mddGkkCtlLHz4sAKVR8rFgEbelXcDTasQdMenc3t/gBPaXlqt7rnGp5
8XTk7+oRVVW47E0GEwamuy7wOo3lLTXUZSMi1pZMLThlV5qILQHimOFjzUS4dhdA8raE3Srzhl/S
cXupunG3QrPldwI1mw+Nb9oRY7NwC3MaogioBbKV2L46zStkq/VQrz5IT+ib5Wh3+dqAmTbTwz2L
TiTNwBEIrO1X6jODVGNiAtmLOBCqjuJqqy/Oup20Ihgmeb7nKXw5DYlJcI594noHdldvhFhzx1W9
JxdiEggjc3iAxy1QUiRi90HotTjxwi7lY144P8GGizos4PYeuVNPn6M8h0CqLo2I802YmPD/STrb
Mb0ViLBLMmlnI3bU/GXdKHSIWzHl5obMGXZM0b7d3vd+8b8hu911MancqYY9O7y1eiIZOkJ0+X99
KcEFnxZJA53oSIdvl1MKf+LuRWlr1kxD11xD7fy2WbyVG0FytdvSYtP5Y1fcvNTBUs4mdmqOCSMZ
haK99Aot6UC4CwiofxSjek/0hl24MlCrMqH/Wv8LGnf0PVES9pd00tVcDx136SgzakQtghM4gtw6
Gbqi0BnDt1cZdpXxFlv8/tqtAqdgfvNkBzqaqWMukBadIeKIsXKrfJOV0vZNX3YE9ZVWY9JWiPoX
nwcO2okRHOrYdJa+nhIDZfFiIHSkXhlAmLuUC6G9GCxSHmiZCrVRR/T6k7rvWbvBnuYT6oKg6xkj
bpj8hZQroBqo5h2NR6zwycNIthFYGgCSVRzfpT5jCY09suaP/Q5nGx2fQZZVb/+Jz4p1oIwuB8Iq
DPCYHHcPhr8DdR/2+Oe6flH9IjYnG8IIbyM+GGRyyJeWKGHXI2iJr/Rq7kD906SMxf2PpcEvNftq
U8dZHwK7YKnPCb8VOy/HPpFnOu5+Jl9wKYhG3FjXwJ8M5csZasmqDkTxVXbcVW5tm9Z0LvFgLAeI
3uuoKNvRxND2Gwl1FzBR3IcKjEEKsOHXVfxMc6Q+EQT/cC4wOoJCSMkgu0Ph2QVhZmKf4OuMdy2T
QQHbZXZYItKTw8+/pjZwRAxIAYFQ6WHfr+lHl34gDnbu6OqUrDI567FL8B//SoPIIKfri5Fm71+k
PlaXYWLsSvwC/ePK+HmVZuItjLwEGFAvGAtP8hZh1BXOszNPTWG7WzQXOwWNwm+WE+R+NmxK+7eK
ppzTkRZqIs1fycS+hcr9925tzCbFzJweWSyTvewFw1YoJkvsD94srqb0YdSzWvLNfaZjQDGUQz0v
eF8vpnK5TZs4zEZxEYgx6Gli/cJobWhvHeBCYhj6MKs/9rv4eHP6hmchPJEB2WmVfY7pRvpunQHy
0Jes/EWaewyDHFCm4pEmsSQuC6WLEgypXd0d+LmiR4xqvTDYsyszXJXx2sFoWNjKCxx+n0jQdnwA
f2PLlSmLjiC4MyeZ7clDVByvPxBCu+IcBqOmoK31NamZ/LPim91JhufKVS/aGJfNdI5Rbm5sE/tg
SGkOtFoYaZoo4UBEMAKZaqKjDPCppIfy0XHW0ysGrVZEQiDuXim4dVkAv2WAUkd/ghAEN4e094C5
bV/5ihRE+sWkfjNIpKeGSGHxbWXF2AzmxvPLZhbqk5gQqD7q4ILD0EnHR+7FHyVgcU4FlC6Uh7r1
zdIHbDi3jAXnD+jAx/afBKBqT2y6iu7oudhibYxCm1ldkADuh090x+J1mSc3JxrHEtPxJid15DL5
/dQ3IfyLzhbJVCw1/gcr7YsHQB9T2pp4AKPc2kMFrlC9QYnzzT05YRarb+q38RcS5OhxnoioVDia
YZsi3t1mU0SxBfZj7lBjxGy1w1CKrYcWEApCDCR2zFsbngFpDo/mZWTp2+DDEQHuRZuyNxc9Dl3R
tU1Wx9ok3cB+C32fa83ZmqvN7klTSoko6ESWmRWQYGLa2/FxzrknEwIax45lWl0BvJ3SXeQMHOm3
x6JMo4b5a2U2xxhhDO4K9kG1g1FentzYDWbtORLDYvjRxOmpohIvL3/8cXQkyhkjQRhLvXn1uCYI
cbf9wj8+OXOpeaVTymTdNQlKQbH7W83IDRfyO+P2/RTTzMAczWkHMqJtZ6/q6eMnXbKdd89Dtcw7
jP7DbfZRN9+DVMG+pKjQS79HRUhQ3DrMNY92GRxq35/BsOxYprHpNTlwCt2yC5ghXBDCX9hHt39I
taOkGSQ6Mw0T++W1f9a75ZmnyXua4DDG9GZAxyR08KNYpDJ97jS7V4EM/5z5tG5IuVVoUNL5hEem
uVpkp5Mf8hr//CX88U0yXEDDYmDbPCLu0KiVsDxwcYb3Xkf8bT8aSPym9MO3BiiSRONr6ZuRVA9o
ljtkq8pkMi44RMHIo9Q6BymcowwmSNU8iwKSSbvXKTJb1dy1ttmrZMKr/JBbfOYV7Lq3UtESz8KZ
oZD+lZBw5wVS4SfhGYjPsn0m6S7A90yWV6htvmVprTIzjpxfZDh+0S7EqOwfjMZao0xDUXGYf5m/
wra26pFbMFAFU4lpm+cautMxm42z8PimXHSirjIJmSKDFg54q1zh8ioJ3wR6Ecso37XakE+yB0T0
RPjT5aGITawm+bbSjn26lCdJJ0dTqWM53/Zo27i24/owWBN+TQSnlzzI+UiLxDQ3S0gbfRXxMRGE
9E4dHLPgkDv37dOboWTBBU1tS7lEVUKxzHCCdwZa0tqAwAKrYRmsVcme1yn+Zzq/VTfL0lmo+Xpg
15wgu49hDi9cugmnXf2+gHUT4EFzQnN6Me8mZP9JMlPTJsUxzotNDlYRlo+b0Y1lTZUwwogcZk/k
SNxNmA43o3vJUCrjxUYjxTYoowG9bj6izZEn3xuSJKeCRFhxY5CTlqf4gjM1eIgTl2Kc38JZVvOf
GXcvXoxcLbzK5WuAMIF/Xn+WuMK1W3WdJ1TOpqmPFgQ7yd+QbZvqZ7XFBxQEr72qpCIlkNhJk8Qu
2303E6taggDibv2IZbRTCXtlwIzoJNO+SaCV9pxRd/1Dg0wyaodsl7Ahvk9N0MBkCAUN08X+5HR0
teWo35iM9OOFnbikjqbqXiGTD9veW+/2W9FhIPmND1G/cmf2hzSEClXJztg+JGUwHkFzJsPN4xVb
m7uaywo0GRevjnzq/LQXZV70PZUtni4r/flde+Z3tLfG8jEkxMmc6uw3boHpPlwRIKLuu3YucOxx
uWcoPGRpeetf5SrfmmpafzjOe81qBcNJmCdVLLDCln2s0W5O74EgoQNoH34MOidtd10Ujk145UkA
P2JzFru4mv/VII5IOZpl4k38GhxgrXFLUNZ/n4ZqRaBjKs4MA13mL4OtXPD9uL+NbgWEjWclhqe9
WKcQmrawNJuRl/Ry41DiPXMOi7em4GH2fHFcVS4OOdpLflTyalwGg82HqARd891zoxfjz7Q2/1wZ
YEcFdXQmj8kYqrm+G4fHdZxnRjUzCD2F5vrgVO3KZRs4FWbO+9n3cFWZHZcMSEgR4wnYsn3eu+Al
wF66kKkRDp1is9nqnLJG13jIO9Ao4cuLnVNpRgHCfvn0I64iDJGHTNDhE4ILWn3rZYYu11bddiKO
WGLfqKZ3OxL+2gB0qztTUlwp8uE0TIUnLFroe2xz5Nc/IwulZk2Joi+P3IkFcAa/Myu7oOve/Z3B
Ke74I0kuX7TCkNyD5vgF2uSKBzAv37iTJMIUZdtaU5s2rJWe4ujWwISH6bex1F/wRWkVea1tG3Mp
crxkLdnAm3n6X6sOvkQ3KG5NjJle5bwB18U6JvTQQgucGKwBAbNk1XgUgELzQmjAAnuPpMLcM6ja
iS0d272mbBV9lzZISpta2XM7tO70+B3FuxTXDiPTkNX6xOtM57Z5IrHPra8GMZYtUq/wzEjzlgnv
6kpl+Vd5ktsbTI0XkVg2Bg9i44bFYLcxl5kNrA/+4Aam+8B1iXrrPzRODshBTptcaegK/IVGXbod
4ICT4gCboFTaGsXm7LeQfeYaXbsdHI5ZiPULfxwdLmOFgOesRiNkg0jsp9CRfRhv+j4kGBJMC7nk
60oKzmrTYfnoJTkN5vn2OjOFbk10wHEYi06emqscinyZ8Z9fnQyvHWt62IfYb2FP1l/O3QwCKeWT
SOtNg660wUxeATWeANKPnAxPjBP4/n+NQCYuZj54NGnf52nFwlV0l0AxUQldp+DTyI+mpTQ8mA+W
OTthtGABbEMMdS12w959w/Gbc2m4zo0agPqrBXg/PXBk28SyhZo1ZzNDq24AoJqDq413bebexkWg
lgb3ttUyd6JI76WF1ESV8daHst1GZxd0xc8YCccxAXi727n6w8Kd81gx6m9aEkSdf+cHrxcJ30jX
QpnlrosEalu/nBzss8jj+BVqJpSer5yBi0ynbyaJwUN7GEpbjs8hojsZGpKoIxmrQp79sfcQfezf
PT5zSvrMyM5uh87XVFzGbLxLsaONEpwGge3jsG20Pa+zKkAvy0NKEqmlBlHHvyIZBZiJl40c3Esk
LQgqXXhfdOt4eh8uf3dRBTgLg2ERCn7W5CxUEtsdXWe95Z5tXOcI7n6WE8NcdQu95zwNBhueys+a
iAyOs/E+S30Mf8WhluobK+EYnM8zav/XLfs9bMitILNrcIzm0Fh6E+6lGAU0p1uA83CtbN3ggR5L
bhl/97LV26SU4Z+EEwTrSDfypkMqLPbKIjXdWfnybof2+medykhwiySFYVcVBntvYqq3WVKp2M1B
a6QYORpCQnl91BfQAbZp5XGcd0iAECCtfDItnROI0drQc/5MPhZda9JX084srzJV6H8W/KPgHqQY
nh1xQhia3W0QeBrox5EMR5B4lK25b/wzEBiEHw8YMrmMwplUNPW3kWDiJmkIZcWDaibEHWc6NDdN
P76MGqorkBXnafeHk+EC7k3tlg+5B/WYzQYS4kgzo1SpuAXOQdLZ0jL2CsS5iUMzEnMCYZaLee7l
gQ6Z6de2MfK0okLm/U+uFwWnr1FQnm99EBkaq3MwbaIKa1Yju3QBeDZ3uvu2u7vQqXbqXW6Aa9qM
2YbW6taJpprd4xfYYnNhtQdlyVe03sR1L3HMNC+oT/SllYH3X8HRzHYwDQZHYIVweeFoyD94GNE2
7Y16To28Gkhy2oSE2jA9n2gmMxCvaXV03wHXF4lJm9dvna6pOzb14lHoUWvReNndz7x1HJQU1/KI
2oU84fGi99RELiN5BJRXXfdx1XZVj0Ct1tcevipiwG4jhwetmeooeQwO9fW/0uu69JCDHOAVgmn9
mrb4e1+zLR7PWhpKwni3GNoHjJO0qnV3OPDhgEUgIe1bVZNoj1F/rH1ncWRKnL1JMZK/0muxj8g0
5Ys7Iz2GRsWYAeyxgqr+IV7Y6jFINDKTBM9Kg907TxYrJIWFdh+G+w6dFN0f/zhCrZpgicRhTGDH
aullWk9h+1Gd69+k3ZWp75JCQ9RPzS6nygzfCbPyrwoXfT3xav2qtxLsa+1jA04+7AOwAQwHcARq
kayBQeok1VvxSLb50fnsLXfDNnGLxnAIjCJoSDmKxrXBx5dVg0MKpQDSKlR/mLH9/CTrlJ2uvnfV
DL9TBe4Z2yUBVYJTBXEc5gTAHSmM0cv7728mjiLVA3ZxVZUjQvEdoeCMUIO/t1cb122onS9z1Qq4
/tdWnzxiuw8EUV6/c4EleIt/6y/I+jwlHjimKnK9u6xpG0QZ6Dv6guoMsDQ9bnGnKWN2f9MHsKSx
SedpHLKu7WRWiawWFyK/+PQ9+l/NAEEJs8q7Nyu5Mq/reqdudrZnezXGZB1wjrptaCVZ6GiwhG9n
hR+lqtYKGp/1URlDmUmifU540kL2RWyOtkYW0+iXPMeRd64DAnKqOEC49NHLyBe5RAVo0QAxeTgp
O0PbPyZN1RYDYdvojNY05bHZaoHFbX2y4WOBjW3EEOA9HGhOR/W6txis/YYZjaI3ef/qT/tPoa9z
u1n37D+2McaPmxNVCFMpJgLh0SpjJKnZPtpfOZSlnjiEmc2WjaKAxbVGBnsZZdEj1bU3e2O8858F
a9VgzOWEh+V5B5DJtAUTSgDa9O3KK+UMMuuqxnGqO+Mqdos4s5Q32dvVdtm32D0M5mSdL/Dxgw6B
6/76RfqFtUDqHo3JMiGVJgch3j/Inu5UlglNRtah/hcMCn4qTRwj5C2SWp4KgMvwcHjIVm7eh+3s
DLZE7Um52QiEYsLANT4F/HCk3CbMbkslVCHFNsJ1TiPd5iUGvJYHhL7fD+P0iPT25JDH5OZEEWbE
J3hY6wemwUtu+23m6eto2WWp8u+OX12IJ3I8DgAbikHKUrBUckHN6uVap/5Umx3MUXxtdW3/Kkfr
/OeO+O14Oah1cUyNwIvwl9MxBil/ZgrEO/hwQkI3XbaHT7LB7+5Pw8ABVcl/v2zd7/ZbvEuFhJVq
BgrZySWFDqq1lJMglCh1HFkaNYfEfJ+O1JxwuFnsFWpSme+brXJSq3+zQKq6FUoM9J1JksD0WMTt
KwsGLSUHeJGK85cEETX8x10bWDeqh7zzapxikIodvO+nd7pMqXRWfVp6CqrfiSXSzgSM30XOhxz3
K5n0uJ0mkqz0AOuLeEC8INz+Zt4mo/u75TkuMdb6YbBR28gVAVezI7ozIq7Wp2T+nSYYHaH736nC
9NwGAN/Gq+dwvb/pQwBIWW6ZhRAszWQV6OM44H1pi4kG/lPyKyZ2hwq1MXi07Z3i5FXoZa/p2ts3
P3b881Nnwvgzrwe+qMM1eJilERM4Glef3iBGV9dqNxdwjhMqvI0DH8HbVNZgJ1c0GCQ6kFsU8FfO
dtOSTYd27LKg9t6nH7JuORzbuqB+YsOAvyCCRjwKjXbawlOHbkx6Jhb4O2/lXb7wDMGvmXkDUxjH
wg8fubdkFmBKVAbO9OxrGv1owCCxIe/sgJDWmCdomrPz9wMvF+M5j8zFCy2FNgl1oHkA+sjrxmJ1
oJwE3UGaFE4hs6Q1YXJtL2zORU6bgtA98HIUR9xQWHv0SarFiIyiGUEz5fsD9NoixnyCNjtS87HZ
tWJyQjWcY+jWt3rW0wU/voA7HNB+Ev2bPD4MXBg3IhjLXcsw95MJa8nXtSlQbiubDFBQ77okV5ob
O8mmp84Op8asXZrHxhm+usZuV+7HDACtl2erSMcOXkFK9VMM2wD3hsSFijvf6w+i6ypudqIftz9Q
cLo1EvmgGTd1XQAKdIe2BPQ2yc8WWxH64UdtV9zXwrB3WBj2Qj1WV6P/zw36LiNAyL0hVc/Hm73Y
9hp2AwjOR+/iO6zZj3swmf/iBEFK1AhBLq0a0zZLgyrA7Nk8eO9kmbHk5BXaViECaCgTM9k5ubTg
FSWE4aYtuCVC8x6Z/t6IaOKVS5y5Ozr0jU09ZU2AtC95RN204gNWOo/doqBljtM4piwF9pg6HSU0
f6/gSURz3akUPT4dwkFA+81aMuvhAcmu9rtsiSMYvzMZiug4KffPg58EA2otHLIpJ5ZSELpMWG5i
Dh85cXjTP2lv55uKB3uG6VBTNWMxG0NcjyDf9Z3XBeV9dYh/Co3zc7dhfVmjmTpw8AVui4jYR3Bo
/M3PFC+auTeGejhnvNsic/9geyhqe6Yp0IQGOapa+fpQYEqIPArwbjIi+pU0CmD7UmeVqEfwtqLI
gapNjondfXc1pKHrHq/3s2pY8gLF2tJxMb/xO9f6IZCxah8wGJnH7WMO2PgK01FtrLkjV2r9RDwi
pUAgeBqndegExSjMYeuGt+yTJYACjn7glLL9pte4BGIdD+K3NtKCF8bWDxXzC0D+UEpgb2jycSE/
ZG9DL25R+fgNGwgyelmx3SfXcYu8N41A9yxGsQuPLxeJaoLcogPNLgJRQpaRUDTDb2UZdFCt4OTH
Htf1OPKqSAPT4iJBFxvO+elg4iSFfVYew0tbNqwINGa470uEfoZ/KuoIATtK4Ix2dnQHMyTuzhbm
2xZsb3uy6JNljyZkG5qfUYuX1WtuLJc48tw73XIoTaFlJFOjVE/MD13ccAcPjEootLNvk79nQd1U
vuCOmcLT/EMWOHcFH3raZRUcd7bBmXbrz+VlHEBSM/IA9ITJ8eZDoo3a8otp3nqNzOtAUQDQDf4h
dtwsM+Lmz7DjcT/JL0Q4eylobQo+L39Y+EcVvxU1txpZ54WFeIsc7IfrX9fexGrorMT6/63e7c+F
RAoao42HwMUnFHjkEb5DSCnJb8ruldWtAbq06emt0IZyETXWTqbmNhIsZ/mKRtcf0ODdc50AdLzw
oxrwF2gXysJBW9jfyV8Wyadlrpbghd7DZhaWB+CKfhfyLgfkEZPYbWblBdMJFSywrJEHk3N02NEs
Fb2hfQHPmH7Kms/ry3gjsVqiNvk28xImp44uquFWg2VuS/Br8gWv1RD2VUUmoegsA7+CvyEThocR
AnNfNXeW2hSQnwveCq7D1ttfjrqKyYgpp/aSM4BdnD3LyEVk0LlqK6hNYdQVADigoUTNmRgnSEx3
ryj41COpNUNm0fpixl071UIwi1YEhbLsNSonbe1PWwMf19BR7KzZUE2weulY+7LM2ZKeYrUrqKVu
/SlHcwo18r+cyKTKC4O0ERjssUrqLKxQq88U//kpnwdUEp+2zpiFPrUrsy8Rw3fG4nMOuPoSpBGB
toOqW1al17An5jnIdnG0Wc9/yPxUEf5jgg8mM858Jbvt534Im0enjeVhU2Q86ysRTDmmHve35DHS
dCdbN6dwpqwKWW+j8/01g7zDdmKhGVl1GGziFZ2od2RaEcKXYeYAcL3xEiVw5e2STWOjQCF0kGLy
7E10gDgSgulPXTBJDPjKs3896g5fx0d50w5Eyc+KujyydsM5f9mA/FKT58zW4rlDUo47nmS4CJRE
2feKq/RaO8m2D+hpCXuIa6WJjRBB0D3knesbng2EcN/xP38yYAkGIbUfwMkY7tgE/goqVdUVEgbz
oxuOLJ3602TDIex1Rx0Fl/b5Ld5ERPNJFFnx3ZdPVv5prJAX9k/uFDFLzC9OEl+tucyEWl9pwKen
D1eOsjsp4+v/izU/Mq80Nub/UN3C35K1s8ppytg6ZlCuTbH1OgbWqSP7wNrFm74jEgIB3AqbThV4
UoDonTXSq3/7wRFnJIl3PUvSBYvi9NjJ2ZxV3+v6FOYxh6eHIU09gIDn3sx25gesiVitX5YhGdZX
lUxRXuNdRRXUMoxsE/OWgnktdGd2PYSYE6S3RtV17wlF9AUQlfnp0u4256i96U+sM3yjIkhuMYVD
pw34k6q4o60cDbGB0PJ7K0rxOzvdKqNedg6OApp9Z10aMtaa3HDT8B40c5fiq+FwpWio5aHaxqZp
tVb/HXUVZxmWeUYiisXSl9zb0mwac2R4R2bIyKMWSyv7FSZXBRvuLnMFCtOy6A+N2hIgUojl/ZTu
WOCvWY8gRXg4bXeg/n7LMVd5mpt3y9e1mLe0e5nQOYDIjex8kmIIlpqzKahWFUeMDOeJlPXJSVit
nTk+mLqdd8cTQfVweRsKb2SRG6OQOxvUalvwusXrKweLpYx7/hhecWlffbqvCKYFj7wRkWol2mmf
yA16WZQbfRILrZDy+5KqSvUmGURDL3czNkvGcRljY/c4axIFhFID7jKJVPEepujGxvHw0tV5PHc7
rzxjv37meFXDyV1ZI8O5P4tJh1fwB9p38awbiE6xmmOqbCJi0BtNuPfDLSJkbO0yPqu4MSSkzQqr
UtFQ7EwyXqbDN7h4el4+czHHgIa/XbZCTFwtKhNo05VPGiBynCVHadIiL2V9BzM9QlMRS2SV3wk1
iG2hTz6fq3M09UjptnWlBn5qcQ5eoQBS2/K/tfMPuc0hFffG4vJbJl6FrIPtnb9jqy5qQsyx1Eam
ihY0zHov61VD8zEWiZkG5Y4N5QF+5vBQgjtmqkjLEox8GJ4CU+PCAHhBIEi+BeyrCiTH9vCKlH1k
aYlCFsXgyJkGpZRIwHtKKhwswL17e0m8gZ3i6po2HXprL5VNQqQRdTZaDLJnjYhNATRFVULKwI3/
HCORf6N+B2eRXfDDCSamQjmikNmMVQh1wfyDHq3y+Yc3OpGCyijNOvJp0xGZ0y4SkjfqGn8hMnQG
fgGndjfw4mYVXXp2EH5azKwD1bc8rT89KsY7MRzUzwoWNr7FbH84taMwsTzVzhYcONAvAjbOVbiO
1Qng6STlw8a2jVT44lcRnKR/1PDP+G81Jm1BilXiWoYj0LhKGD2/sVygcOUBUP9Ty03kL+ycdFqk
JJ5lzhiJn/oePoxnpJaYWN/xwnJURO1Bz08i+F2krZqxeEJlzqw3yu45vr4aC9v478DJejEyloy6
gEvAYwMo50SDVfwR0rL3kSMjSY+SNIXjV4zugrvmtVYwARKcZpyLj+05tDgPeYEgwKg/7GrQgmWo
VgI1k+g+C+zzs5Az0TkF0euSDIS7mFEorMKnSx6IDHtPpiubVrd7frx0JOeX+SUTFNYYHm3Ue9HA
Gz1iRZvdeIPgw6KkizlSrnatwcOLOO2re17evaa6/vU+ogXMR71wDn+OaYLq5yJAtJpEIX+yxqiQ
gIxe+lq45qzdOxuZRxJa9+mqZjPn7IWCe0drJAhiIGdKE2t2TKzXr/MXcrvo7I7Rqp4VDlNsBZP+
t99XBhoDKBzGLj0Z5WbYLMd9qxteuuaHv8K+m7dSj5zNi8MZx6PbM0lczMYzCMnbsNNJ/zk9oATI
re7/WPJsdQvi/e+6Jdvt3xsZkqDZ9elDH68iUwFf7eHp1al+0F5g/ojx64Z0XMw3UahUPyBOYuNt
Y8DojQ2Gqf7VZxTiZ7TXKtk8ZTDejA8Q3hODTFdq9/9LD36qvd6CQLCQm0kEmijVsX0xaJSqsL19
NOzK3OHZ3Ie0y9PiywyNfRmG/bOmZmB7/FlBkJsOLNNs0fE7L2d+G5/LvtB/3poaUFNrt+6Ncw+B
a4tx1PDz9OeYeZM61/E72gpZjwnlR0EcvqlN18TaS8gjEMzUad8gcD+82cIyx2ppLseUTdfTS/r2
NJl/w2HhIEPr/xn7RedOO/A7NnkITDRp8omQUJl0TqettucEN19MK1ZXxg6iCJeDFleGLU7y9eNn
q//r5DBelszK12/IDppPdGzb7noCVIlGs7rrZoME8euT/EgSUhbViwZ0J/RdvfInCCu9iJsV/Cqs
ogkgl3UQ4CoBFgflaSfxG77OTS3SR/YMoCgZ+CWDYd01zCVWwGehTKFeUkg3js/8MI6cl+3GObGN
ca1FqK2wyJx0CX6ZM2Tbx4qPxiiLbanoBMPICjVLgSTItci0eiED+hoxEsku1viNQGqcx94eVTu5
ZszzTVAiLu4O0hHyYweg9OlMh+ofvDmyL9MlU+9qhZIaSurRE+GZ5S5QCN3RjPCJ1nRr7xNYGc/t
+NJJ/+VfJXmU0HHETvldAViLH1YGZbUPQFg2wxdvrJiEm7Rm61i9ey3MPYR+dO+zNy5Ok/PbTq5q
MVRCBN8zYbmqBNBbRQ8WHzJs/hiU1A+5A6Gg1e1jptuw0U9/X/SkhbDUx/jjBkX8yRpTl0bg4m1G
43nKOUarRUWmOtcTrPJ72CvbJYmhTCJ5MFayVvVAwU7jdmgjIc0kz+ippJmQXi4hZHE9u7OT/eTh
nKsP2c8k3dc9cpgOYIhdY4tYIOLjzDSPxPYKdMc9Hkr/d5Q/M50NeX9PYnKaaVQtFiG1Ys31p6gu
6Qx9Vft/CfJrMz7WTm1hLRiBq2Z6tgd10gAIaf7aU3lAIc9W1AlxPcdAy18RQFmAjogi44NXWG7+
dt4d+x8/qyZmeI7+MbXgYIhW6Hk5z2UTWmX8z5+NM/zJ7Ki7SKXLLJBaUkdTa1aaA4cB0CQB/NfF
7WI6MfUzRRduTNp06ww75y2BwU2DeL/Y2pJBJ5jucUpFMP1E3sxbiC1C8QnNbsF8Y7UNBluTCCnI
U1v0GyIfEg2CbEY9AOhGbpy6FETXat5cu7N1mm0xZFmJbWkH985ElNtFZYTPswbedaD+tMCi7jeW
xb78sfWTN9h6IN9yRwacqwlcRKD4LGO/Ou/cblxwL9H76wIXsli5YnZAeG5D1atQCU7CCtn3igcL
IwhQO1uv9mF9bGE94gHaYBYNW75kknvknm4oF5LrGQuYX6o7DCDwIlHvUt5cw2nOKOb8pNfkaSNL
nO/tEMgyGeuGTA9yNP6SjO86Vp6VaGAXXnZUZuZWGxntH2Ujmu3F/5sx9fzwQ64M8t291Ctx6eV0
5y76jjhDadXBl2Tn95fU9ldR6m7VMOL32TnJ5bkmBiIQDbniGS8a5YfYfhynkQNajBVUbFjYoerQ
AvpCnpZRujdt0Y/xGjMzmBD4TTR3S7zNq6ofa0z+IHljJ1MPYS41AFYTUWkMjeYnlHB0FTVIoBvc
nWV/8/UAKS0a2sk9P+Kntomo8LLB6s0P3oSM06eiLatf9T81V3UF6P5D9BhYiNXfB3Nb1q7yqzWq
YzJItdl/hFVIH+sMDY0jpg1AWd//4AKISJDXyXKcrmTfN+fFPrSHTk90NJIE7vtlzdpNhjvklSAt
cFaMIqoI9Gh5u1sfdUrPqpwTbg6nntHq/H5B7qmw5ccbTH/ygy4wdQNefU6cFdMbvAiM2Mn5uEaH
aUywpPwJJ40YSYJZnJDFxZxVaRd/7d1vZdG26RvH5VpqArpD1x6CRLJriCE8VJKUTwjTLmUSs4u5
Q2jHS1Jo8AsWUyZ2DYKdg+LIjxq4Vg4ycKRx8TMibihVKBe7VvquKbqh9QJduXC49cETkJU4RkRe
vKQwkh78TYDPmNQWzrHC2bEFfPchf//VkBgKRPGP8X/h4MjnCwlo/K+V5cWKur4YKT3qQVUoQx6G
okFB5QFegw7wFqLxk9Nw8ZF0ZsPOrP+HEg9d9hbgzRSe2Rj/9cIpwqtmJmiotav90jtgDUtEsJd9
2yFZ6pux9oIL3lOK8EJZodDbJ+pDqj7dklSMSHmzmebFF2e+uA3XFzcplsG8+PSpSPa52NGA0WTa
hhplcvBJq72lkZcxO2KUq6F91IdQKPpRSp5ABdtdRd9QXAV8+4CWaSPn/JSYYV6r9uLa75Qe+ksv
ZNfHdVMZyStZx7rf1SN5sNMD0D4om3hlO8qIKX5fa1J/ALJSpoQIZKtYPVlW4Z1atQBurV7OMDfO
IeLA56d5TWU3hCZiLKifI5c6H4956O8LpMaNaCBmNZxOegUjORfQ1/4B0cTb6gk4TYsj9srVQcht
LpcS/aj3iCKHjPfSuDvykwzVKGgQwmfHbEkLk/W8HycBAVUdSYchfhyKFjsDYFDxZ3oSSJmsG5L/
f89vLDIpGY7+dvQxS/6Vl6GN1tTKbzz7gIs56+6rKakuUCQDKFHZd58PTduywY9GYfuyb7TRR58O
V/cuABMw5lOHzbPy1oXD7HDTAG4uJrqjrz3vPhkMfB/iNUrWnbkliBLNuomLO678yKsvP4nvdSbk
jU4O9zUQYJpyAuunJlk0wFxWkIKeOlwGHVJnZ44NGtJ2ZUT6tCRo91sHBEVQwFyfgagLCjPIeitN
McmTRP8YHJ6RjZC3FVyiQ7c5Ej51RlPDNWY9cpITFJ7yCjBfiAf6JatWBhZxNouZQrkXJeZMmklV
etZk4873/IUppX7GokMu1ydpOVdw2OmU1AQ9x5Kd1UXcidVbGCE8t2FEKm7YAZMsatTuT3VpEzfS
r1tFLGcbjaWF2ta2UvhtuAetjEeKqFr/kR3b0uY4nuplHyPA4WQBa51x824RX+07Jon0zGSzqWq/
Yu/JB6TUTBHU8I4pVxzwkkFpe6FkhUmrkm8eYBPWmHoLh5iMh4Tgjf9Ve+V2mP5hSyE3iIMacxmN
OzYTYUnOTta2a7jAHX7+r8dzxxYTtAfmmZcZlGFtp5xxGp8JyWU2yC2Fo3f9oX1CJkhO9xRkz9yH
BW5xFs4T2IptY/xRh/D1NkYY4M44/XbQ9jyEiTnHYdWC+B06mAe+Bbf51l857xtAyfyYwylSayPO
jltzf2n9pvjfv3iXMIS+4NPefAeytiozgi7zalDAzCdUyhK8xt/JvKprNbCSxqmGvorGAd7MJAfd
JLuChFts65e6xNOfH1wZeb0VmBM1ruijynQfF4baBtJn35qzdWLdupLpJiZbiyXHZpI4Cr9EY1l6
HkppQmB7wvuoxBL6dbcFn+kesou53cpz/eYldx/xnpLW6Eqm7XPCkCX4ekY7H71qVCiK0Z43JupV
e1QVh138Ycs0n/rsGonbISIKDeO6VBxNNxcBfrpMCBVfPmNZkXIpFmRI9gLntK4DJlOUqVEjuAeP
5O2Xkm+mVrGxg7URvrwSRRtWUOVoQ/hwzIlJBKGuKH2phgo2F4n4odQQ5NI/EZnTQoUPQgSkW/9j
gYF8qVmOoZKPciwo7KTzQMdIdCsROrRxw4CQAfSesBZT8vUgjSId1d0isUDyG+GHyVtJjd24ehya
t4Z2vLhloJ4Gbo8ijYzNkOmjCGq3RW2Kg4v73kEzsFUTXV4W5/xS1wW2CBQ4q0+SbEels+lw2NK/
hRk/ir90OiDsIHKK7GDjbqhUMpweW0QxF1BJ5PuUKshzzwFVEUWMs5SGsHNxgMI+T3GwGf1az5cK
LBj1iMoTV4XdsjGLQ/xNqwbUZVl0bjwP1gu3+Ed1c0LqAxjVZcyvM4Dy47Ei+uQ5dN570DIhlK5M
JD8nRh7j/n2AIi2im3L7UZwi2Qvm6JEKs75NtAY165p0FIME+fctUvjkCt08yB5SXUDP8+PSSXXG
QPZZ0T19TGzlwDpRJxM/8vC1cVWj/Lc10yW37ILNlxTns580qxcXiWj7KNzBdsW4DeEjEAnbe7DK
YNW9TNaeaOEHH+WEaBpcNZkH6OeadLWMKWWnv3TtYJnwbeO2ITq7IZTYXjzIyoePrntH14HrvCN/
R2NODpSTjG1MAQyb1oAn/T+Ad8eS1N2bQG4KUvDnKC6rKrL9CkvA5FVQPUk7BIjasGkwqfAe/HHJ
4P1Ii996Q+qQgaxXTdnOqZYpTD7wSwe2jDaD1sXcaRaMSPsiM5zQSV6jgyaLPKeKsiwmcA/96em6
flIVVxqJL2ld78CdIuQSmml1OShE0SizA3OFuAVR10oHeK3g4zagM0dQp0d8ik4eMeE05xBopKWI
hXzKFi1hD8im/GaP+6ZXIXAN/C8RRShctMxUX3qzF5HKHNa14ytEC8BhgLz8Dt92mUD3FbkneINv
YTf5Hh6iPlvR3Y0CUG6IW7id4OoTnPilZ1HgJfbhrQ4NaU6iNmlQe9+ZqVZqN40KY3Mwh37YJGoX
hhdve3zVWcFR7l56n6HfzHgWXmLLc1R6B+LyZdoACPh2UO6+NoQsdszQ6DX8Ns9Gd+Tkg79XM6Gl
UBscwOKGMcZZppJABAk0nn03sCp1DjKnjeja8EnXO3lhPRlmtB2L6ZfY0XYvOIZfZVJS3X6H83v6
bjo1Df/mytw1PMsjIx34RYGF4hR905r2+zY31hUr2GP5EOLm+wTKnezHjd29Mv7KB+mHjUMH13Uw
dB1XILXzkKY1wwP1w1nuO2qvjwjgVZtSNNUJXb1ePYP7SD+O0WYAvBRATFI2rb8GOLOtjrI5VVPS
OIJqNfw8TGgPGUGJX3A5fsiYJe/0UElPLZ6ytqLlk2c9EuVAG30ABC41Z10VRahFSGp94A61o8Xo
fwIOUBbfLrC2b3Y3VjO+rxov2JpBWLyrspoSCo6e2UrMwjm/nS5Iegg3m/xmqkPfG+7H2fp6bmf8
jSxrdVvZRuG1Gb51uHQbJijicU+9lfjoiu0Z7zxrEuDxNiYUU58OY+Zj5dhmrcdgVUgT3nDmJ8By
jqOqJ6EnwIhPuCXkf+PlVoscqFF+mdyXH2BDNcpkc4WvBVV2EESb93czJORfafnoldGKNOTk39Jo
Me0cx0AIjT1FqyFy1ysVhu7qzj3LWRaPVEqXaE3E3EQ4LMGQjjnD78kLKtJQ4xwkfaJRkE5EXwal
mbxWAdzKBxZBViWeO1de7Fqrw5XjP+I1Y/xdai4YM08UJTO5nK/m5yCph+RldYxq7e7bkXEXqNlI
q1UISy9bJJJo1jp3i9CohD8/luwH920nr9xUMkonZKQSUCTaSZwTpGAW3wG5ghFvtCXnxlOCYydR
XhvT6AsX2A0SguCcvRhbQGWgUWvqZjMMufPkFcoM7xPiQb1SLVtpx+ygWc0gtIitennQ4s9M2PaL
I3eIrJSvE2oA9dul8BD2ELSyQh5UHXVQ1/gJ/wtmLPmcXDlzUF+CSXJuOn1hxvzLQ3YLp3Gr8THk
kZxsaxESVht0rNi8yLwrHtp9/Vr30CU5XFC2m6J2LAyhpDIsdecvrhGOLjXojmhhc2Rw3wwIxJ1h
EcQt69zlXzv5zKZKtJtfNy/Ds21GWRjxg3jiL5Fkq8meKX/+0ZZ/y14NVJ7RNIfPfA4r2cXWzx1F
I6jcv7x3hNSh1Jpc/Gm05LiLcA8lFcIw/tqU/sDWkU9wEc4AmKViZ2RVFoRiJV5uEAI9R3EeChxy
a8GmlnpqFH91w3Cyae9qzQ6LdwtQfYhiHtjmYyCTxtcoEWMEZ8EHwfVw1if46bYea+SVWo2VBkHX
BCknH8nhXJuZOqMAcAwna6qbU/kxciPKA1V4zyrpz3zzERHP4OKf9o3gUxoIWiwYjDVf4J2nqyLb
fT8QPi0ppfgzvzk4SAf1KkyykQMLdzYs8EbRQHRfgFQ3Hb9Cw3PRVjx7KHAWWCU9sh4+gJ4D4kc1
ZrZme7lMdzUv34mHkGCbEvh9fA2HILS1xtlJveu6rrO9wyanD5MMwVKP+VJEgEdPkgZRa6MPogh0
1o9AAeqSwihze5jkmqJfyvfLHwlFRBItBdsRO3t0PdrJlQlHYYk+NVPg6qTfDYiSsAtn2pD+c9H1
z8TINl8AZXICILu8Le+CraX6qP42YNpaNQglv8MoQL3XjXykQIPrc4v2ncN/7sk9RprIZTuWxaZx
4iD1uCZq9KcMvsyP5lew/rN1VBzsZadvxiqUkRb3SPGBw83+ctjygZt+oRDSWzFPwT7XEIpLisVo
amifu1bMWEiXaR2NtfK82OIJ/HkFQtJLD3ZahofoJl5TVL46uWEznuhuLRjFb2ZpYURPS6fTmRzs
fmCryJA9jvUyXphZNI4B36DT0TrRUFVMaXa8aWvbL5Mg1p7giZV4LtwVH1jmn0/cEOzL9bUSc5LU
xwDN15AJRb6h+pLef8ByY48g7+AcLN5DeJ2rxX3G/H3NrlHSoU6cZtQpf65wYyCZd0FA5ypeXGzS
H2SaSUIPQ3YrDq4EdYugnrHycQq/6xxkCsiL9a+YT5E5CfH0pYoP2EGX0SEgzU7l6ROqhKVxG/PL
iIymD5+u+LigTUdUPkpeHBHvczXsbp1k66tqJfAinYdA/W9feo5wVVMjSKRUuZ4v33fuG7qYspvx
dNhPznCVlgR7x3iftgQdQKAHZWN1iTphX6DNZZ97EZPlEIQJHYzz3GUp2i+dEOODTtaNSA+/TcnI
pSs0AZdtMxQ5kBgP0j+w+tdfes87pjiqYLZQtogphYh13+BeDnXXFmOIkzWoTCB13FnmIEh4mKxa
UJaB0FLinL+P+ZwJB5/AjvpuFoY3YjLLYE5Fje+3h1wmZWpyST9q3rpHxN9FXqR7/K3hNjVCvbdz
zBx92ObOmtER31SBKmH8kPKVGpkw2o4lUbX5Us5vZ3PFp4YRL624wgGbpylf15EncOiPOQsW0Ngw
x+0naK8QZiGgSvDiCfs8C43DhNDtbhjhn8b0Fke6YfcUCpbRikGhv/nvg8ssplPVQX9sbtQ+7XDB
GGiDUvU09AVbvbsgoOtN19HPpiIlZLAjRvW3KQKZYjWY+KSJdgl3uh1fHQjYOrF6rY+WGhGE11aB
Wa1Qimc+HB2WgrhfAtJtxZjkqSAykpKSNvMpv9g6jyJnXUcnh10QNaaHF0uAv1d6JmhDlnWF6xzU
oLYvgZnPgJbMpIsXihEIp8+JzwYJzN8xFBBjTr+nMt5ygyYkisYu7u3rr3V2MjfKzNuvuHA04xmf
YPCjB0hS8ehXxoUY4NvvPqmGJBM4Ri6NYLy2GzFAd2+OZj4XwtbUMkyjO3TI8/LXm+Vrbg7G7CTl
zQ1mI/BJy4JcucUcaXOhj+ikkDduLBUFzmWMBnso3Bkvyt0b1IqAXywxHz8zokGNknouIjyEg5v4
+ihX7T2oQzCPFhm69QYaN9zcXED0MsXVGT5FOaKwW4deXxcnO7+Q5/ivihhdkEbIR/Ch5iGzF67v
2L7wCz4pJwe/aYYP0edIieyhYUIhc42IyfVoiyUK8r0hwvzsa5XMenmazYm6HMBj0RN0uu1Ec3s1
+CwP5eSQIQ6v3fD1Zl07lB10QLqm6DEP+JDGWqpBj5+T3lOiDSbJ7YymbDgqNGC2dveeUrivJZIk
99JVXSorHmRdGtsFBi6Y73elWmTIvOHHWZowdwDEd/NVdBDvC8m5pxRLSALfU5CNujHH9yUSsFUC
dTBMqCC1MIGD123/ZF3k0+IVI2SCc42wRZ+gt+CDvp1LsSfAxvavBDOrC37HOHjAcOnWvDL9xhfM
sMon8obS176RV5TMnj6M/GV7ZQyHB1teZ4jg1ufEfQp5xgRBBUleoSmVwLxFc0TUgz85OcAeHOj/
YSJwFP2Sb7uMD+Rl/gTDD88XZbLfTLRp9yeOadFqFRbKtMRp9e3SiKpBxFCpOZvTE80zgrQFY+LP
driRwX1Furcx7f527Wv3azqYYC152pSLyTGgOttGoVuRgQsRd2SZLEWZtPFDEdgJOigOyX7c0g5J
1DaaOLeBwRgQ/K1YVTt5YGdX2unZZiDc3UmKLvCktoHKQ3z3GYtDsPb6Wa65lKtpaOsYZz46ZRqR
H5n5DmTOTVDDGshwdOVsb+gzgq6qlItqr/x1IlQC/+BZsGkXznVyX6B41zLcgHVjMrSmyP6XQbAJ
sBO7jtCM3k1QQ5bPEPUK/hEBGUp34P/U9d723S/BRIFjdwuqO4AeTlxyknF+pl5U8IzgOurjbKoZ
gDC4bcO1F/vndeaKviIobYAK4m3RujEAX124BCwbvvE7Rngkusshs+KdAUr0TSJqqmaXiQ6Grihn
Kut4JuOWGTMHYpdnTXGeOMxibXr99b7nGu3kahFgN/OtNSiEuNJCxLO2X65jpRMYf3Fif7n4VHDu
piJJKznii+h6iMIVgFGJCL869A4NSlt5iSxQPDXllrD6RfqTDUhtwlm5g7zcCHEvX+c70yiLjcXA
P4mt+8CSjTIhTrbwWQiGk8DCLVwzzg+4v58InLyx6YoVvLzs56H23FjnudcfG/E60k8O916VfOc/
4b2OD58mq8dYEN0CODuFO02f2ysSQARHUiOWBaLqZR21IaB4Raj2C7n+q8vgTvDFFosuR9fj9xub
fwVQxRASzaghXn3lNNRwercHguNNwbZDLFmU/tK8UV71PuCiaKuQzpIQXMHddZYuzD/gyj1hpQtj
7aAdQU8mSbMBUFqaFUco3Jc2qU1CNX+F/gKJxx97qQTzg+ULteZ8XimDkq0HMd1hidyQZPt8/Igz
6OdBPZ7xf8pWax2k7+cwV94H1XJJgnL+HflHhw/L/v0sLEsluGI4M9w/EzJud24MGeIQBGqvFDO7
HB7xXn5186Yj7y5eGcR5EDA8d9ziB3VdNTZjJp5AK5lSvmI5GbIok9+cGMN/MDHR+Ke1LgIguQgr
ITie6ZAw63bpGuWmghXDxR2O4P3FoqRzU3G/Y104Lynf/n3sZxAGqJhOuiFSvB7/tY8dw+HhCdMx
rpzHpRxbQ5LKDrB2qbZQfemW8Wo2/uy+Dqu5W6zqk95QGvj7jCYv9oh5ujvB1/Or5EUljz5lfrxc
x4Dm3Hsi4xvSQQTc98BBci+E5EyZsZQCIpqd9RjR3Y5sWOYECxbwmLW1apkJc478/XcNS16GOg5a
Mje8vDmb7jhCDgXuCqT77a/FuEx8xGKLrtHGgFxePPocCooYDZ+1V2ydzjNDNobwQl7DtoLq7fww
0D/+x8R8j1zZZRX8933dVYoMERSSa6AEd3CEcKodLl2Z/Tj/UA4Fq+USJeNJetdH25Fz6yUIOWI+
0F2JXVTUKjsPXVFQuvVAXp1+RSTcFEF4gf5TkhJN5/tiqBBShl9PTc9QAXrdVayQ+FO9E/GUwBLv
xQm6JAQEsR3Ra9F8+89hKpmXL8Zc3/496jDmYIIYl/qpempIb/tsm1EQGCtlCo8x7TasnzLkM0hJ
iAJeSNJJ9yLAiudOnVQFHkQm+Fd3XWcv46UXp6/5K6Z83pQo7/bluNTU9PfM/x79cnkCUK9GbCJr
4pHVnMCP9ZDkMTJuqDfbEkkebLnz02R440TM8CNfcbK0apI1rkvuXstbkXU/vwRUKqHLXw40FlvS
iAP11s1FudqXrdCxoYkY+YtMF94bnZnhQ2mhLQk7isRR15NPpc1CM57r//r76aZ3fFj9gx1qifDq
N1YwUkP2D8omAtc6hMi8AmhiADd5dCjNuW16IJe1JkOdl1Dw6BDaXwWZ72++U0eFZkO4uZSgxtZK
91bWKbhGabO6p8HU4a04X5NgR701j8eEYVf9ZvJJpaYQxjMcK3h3GeY051MSxYnCfEea6hG75LBL
eL0cavr//9U/udLJ4Qa09+Nr/SdmO51G1qTSiYvYpr8Bw/D6NLsdQpvpwVXCTzdh1vQnvE3huuDB
BnOzbsy/jw2kNBBWAOQnZQmikz/8gWNB4ZMdx0+FDJTrL4h9E//6kJmLBjk+AWpGBGBlZbln8SEu
NYi0zk6v9Ji4H56Hus6pX/EyGs//Cbl+Tcx0Pb9eNSTBya4+nZyBgE9VIHrhLJ75pHVj/5F+Kldw
aqquy6Xxogt7CVfPGBt4mXbKYe47Kmi6Lkq6gr8qncaw6ugDL1HK1pacCqo1pt5umt4VhB7yVutJ
IyUV6NOsNXATbB6Uii2cOS7mUArRiNpDh90YoZ+Wkdpi4fYLh3BwgykKjc6Lj1TfkNPg15LreXsE
hYGurW2cWttzkzeKk/M1L0jYWxWpxTkFEa9T/lBgOdb4muDy22lnjPXEPFdE5fHjEn8SfgjaQbfR
POEdU250vEPVCL3VZOD12VuPNp+05w6q+w1S+RBn7mDoLY9ra4UphxQ8ECTVD8cxi1VESXHa4WUV
DlBeHcWwF19BivrpdQ6X05TXgeFo/ZtmxAdbEmX8XjpkNS3LtRhG1bneGuwihMD1z0dtnPQT5BEI
xAM8LDxHd+o/tJwCiGdu5aR9wkEQDSuZkQRQtk28ySIRjPPdRNbKIvaKiX2RaaNFjyHc912BNdlT
lWfjlI26n+7NZ3sxExLdAgAjEl5dL1JW0lX1ehFZkdrhN/rAGC2nky5Z5K2D8jWL6TZd7r/4x1Bp
QJrD47r1eQfCo4wudXIaiMd7VZmmMT9mu/YKBuBIBiupOaL2+0o9adWaal9D4QZQdb0volm3jusi
SOUxZvLcW94/4MRKu1tzQ1klx7TbhuDAyBDRvjxzD2kuFJI24H9qBKW+Q9Qvx/hpTMapnNrMgB1I
CWRFyMt172svbTTFomH7JFIYSzKiIzMyqbRv8J6K6EzD0YnLZ1r0fzgJkWUnJpJ2PN2Y8SB+wDhI
gR38WAhXpcOjKFHcHSLKxTrInXdRZr3GT6vH1bktJZvGObACH4zasIXGXUkWP+ltvJ4y1gyzIXwP
lLT4cGMkRiyV/wMrmnO6dblN/ZPlOGGqhKLzZRxzOcISQWUWJxoZl01ycGNOvZ6CoG22AFnDjnTA
8z0zVyzBDb7bOtVPSnq/6xRV2FK+26aVLWt3lLWIUjtqWr7HiB/W3kzxmthxnngbuSpRWtkHjwe2
BwWwSIeb54Ad+BJpQuoWkSDcymAEcEVtuHbvHVzkou2ADZ42qpN+GmpSOUblWw9/LJLtO3jfMw55
JN5PRI0hak+qdMRRYsKKPG1T5rYq2x9LRjhcwxPBSjhLDwjAQ1bQqidxfsJ/obucReBx9Fp/5x6n
nl15PUjjeE6EtHvAawN8xRbfx2wGo+n+TiVv82TmRz9AU5pexoSc91ADr46tq/jdGNyxqs5Z7mm1
DX++5pMjPxxCjJAD+WRjWr/gqXB7h9pnKmmgrwP+PvxzIUsqHHHwRlxuTk/EecIR4DH1oaGt7jdi
/EoFPfFoJXOD1UCrwpvnQ/nyq3bQhpPuq0u0OuD4r5bUcrphF+mx1E4mvKygAzSJU9kjibIZwN6P
C1weBAqbUHaXdN7AnlbbYOaQ72uGsaZYA5ENihm+Br5oZSL7e/68bp0o3zY+dcB2J3wMX/IZTXul
wdRZbTqwrPM3EzPOSIIlkajpiaNJXfuKxZu70d7Z+0MSVoUD2j925cj0hghydJiQGq5gIMRgN3qM
6bZu/tKck/FZtNLiid8+zdgcv4YkgqfmBKzrKDdjkbmWIVOqx6CNv99nfVCvlXBNj3URmHHqB3/y
+ZwaSgtYqgBM/BpW9apSYW2Tb4rQFwnxJXQV3qh0QAxIdz4lFOuNxp7Fee+1/YV5yOlgsuQJGBHx
rZtvaFM6Hgn+7Xn0lZ0Y7jKFaB4qeK7byDUZ2P54hLpyHfzXE410AxriLZFPP0fkL+ClMksCXISh
cFURWejzoAqw7ZE9sg+OZ2AUC/x0oEWw/1hNSCQyVANWxA42FW39J8mCIgHAqUONiA2JvJP1OdEZ
l4Xpyma6cdLwtaBSQZOcasnXynO97dmwXKrf14m6kguFKwX0J/zECwXGic2l5FB+xdEcjlo6vTUh
UKPOsff1a7bYT+kELV322s5PzBSk8IA/emjm5rmBebZe7kuAo/BQfgyOqoMYItkcrvU50j9DiQ4g
Dx9LkvpSGft5nRHm8k79jg2T57VNoF4Kp34xQ+D4yVLBXs9bNGKxgOa1g6+WsSF0v/EVparC1phF
rGXSzSrdisqLVADg51MLVuSpu5rls5zUOjDmoyxByynVbcj4Zhs6nhdlLgULDKKVL7u1VSCxEn3w
jsqOc9ZiAPV08VjLLncKOcvsgG0rnQgAb130G44/gWNFWIQdoJZzeRUjpoPlyaYYpGyP3EmaSJCM
5H41DE0W+clZUQQA89ZmHBcaaOCabo8+63EwNqJo8h3IcNKDgzb7UD8ill3jNbOgLerWotMpgzD6
G4BLe7xBHUYpuHceojdZsjaBD8P2Yf79EEB48H0Ox7FO9re0nLKlhZylkN4ZBqO+Tciy2IXs0iJ2
mqLZSx2UOcXK0Oa1MbZRsgr+OLqC0UtOn69ZMxCjKvTgyCq+YKNwVHDK3u3ksADGcbgRd0173bDu
pnHFftWMGdmuzPIi3w4r9yrX555KjM7eHK4KBML69ToN95Ln3UpbmBRKTvz9fa62yEhvhbHs4FFu
700Z5W99RNy7nd9f7PDbmG+IDcCpzwj1T4dDE0CZEMNhWyDO3pqDpyBDr63R7qTL86Cpa9ybet7w
EaSxs7ER74wwEE8p6+2RwbQes0H+Mrih9IRyavl0QGfR2opCTO6ZKSDMvV18aNCcygrSPApyO7+b
RxedM+hUEzsZQha5XjKYNWxmSTXuCP3MGPVSa9WYck0J+GQKlvkmESU/YUYuLjvbOzBqmJFDNzkd
PeGq6VLO9hjYMEzpMT8hTuuJhQK1O2M/GxXR6BbLToyQjlp6QtblJRJiL2953Q7WzFn3ZM6+8OaP
NSnf/1tv2aZkHnVzGrvhojFOX899dVWVnJwl/nZdLEKcy0jh9eGDD60jmzNUPKq0FJzqePv1MzLn
bJCgm0toMDSgxJ206hMQVvjaYEPKFgGiYUzZ+xGysuvNzmQLJR2U8HkBAxtT1xd0mc56xP1RUcQv
m/1aIlxB+2vjIcbOgS9+6m/Bqls9Z3B2xSy6kbHXOa96C0QxSCGxVxvAdm4ixS/aOgJ6yCb0olAA
NalwlCbh3cBMRXB2lAjtjCp/a/2cYaEfx4Ch+qll5m6svGModU1GDiEftm7XZz2nMOKfYym/ngkK
O7+l2g7/JhHgClAFm/9YL1Pd932FGlwJeQwV/9fbQrxiSJQlpWM1lMpO3VmQz4nWJRmFJJmJsTE8
pba8d8NOixMidcW99HxXALKhmo3niR7fSYsfO8vDV3OEfN0ZBP2zdKhDR6dt+m0OSl4Arn7JLwwX
olJRzmwBNOjH5qTcSkFK5MQ8woWfW41o7xLVulsgdzdG3izVGBRPqBahAeQB1AahPRs6DXatp69H
DWFu3dSdLQXF8zUA17nT3+AZFDhZREcNu5l9snnJeaue+JBqCNeU6TYSP2bXuwuScQkliwLdWmRZ
vdK3vS6hztAQ4GKgg8rNz4RBK7O3d5XbGHu1iruPbxbTNCO1R+QMEWMLY9V4vTYf+oqreVgRywPX
VJMLt1EMrlEwZbNnxMTJVin8mUkHItThtElVUGZXylWnrlqvao20FdZJyCV19wUVb75b9T/DYJb7
9Mc5dkrXfJ3Q2BiI095FS/+4jFRtFaoafnzdumrXRJ6eyovm/cg4PKcS+jD0IsIB/8MCLRy9boox
+iNPuG0LE37zlW0ZbU5tKng5Xq1VqMqrnnPPQqMzvBWMC3d93jD6de06pxJ2/1/0ThO8X4wuqKms
1nCn5L5NBy7GCch3URPTrBip7QqOQ2wdQQ0Ed9n5fhxefxFmI8AKzY5kphpHbDatAyVVUhFJvjxT
fCGdXIHmy/CottUaR5g2DXd9yAIqxi9pmttmttCHgj2hK+3fu6ThmEJdbWdBix7s/NPQbvexifoC
AjdtsbUDntrGdn5LySc2AZbs9kaZTn4WrmLckwefDxDekEBz1PwnpkZ4/iyZwWPry2qV6rtFy8Y2
E+ujV7cKkrifH4FZ2d8O3jEKQ3CHQTp7HlO8wtXK/+Y3uMjCPxTGfssLi3gV5jRGH3HioMYSRwi0
4sBIqhq29wvarLyXU0CJNKvH0tyhfzY1Svgfhak2sfyDmjZXBQLHMn/Ypktr0ASP/mJCHxwMW4sf
HHq4N//vDfuPkpTL+RdrkItRRr8lZc1HXpURWL0d/BrFSTcHmjPa1Ko1jt+Gx0/y2TurJNPcfMA8
GSOooEIQUxacd36UVFNPtkJModK2bL3sPvPHWqsVW5TuYSA4IIZPTcpNcykULehIIUDxI6fWmps+
CTsUJM+W9StDuu2RBdd28UVTqiX9YbrfTB4hHjvXsX6VK0P+jqwjz+r1LLM9MMSOxQV/njOcaZqp
IPKxwN7zMDlpl/gyQ2/6Xfivm2Iu09EJUAOncFBXbqWg7c4u+JRkPTmi96L3gmcQN/it4LoixQ9A
WSpKyIX8Zh8Fsz+XR42B4T1fFkNBf3pW+ZIAdoxfHtuT7LLEjJ7TSx3OjIE95B5FPYLpAJx8PYKS
+o7e/yvdOg2eWGaGDBHV59kxF75zIvpeRM3Vbb2FxNRfSeGJGP/XW7S54SL9NUB/G3ujllhaJel9
SfLTv5llGDNRxNz2ZfsxVELlVUllUhzdBfc91GBln/M4pLULN4WEvOYS5iLIWw58N/e3Fp+t4v6w
IhOD/ydHseyajkNY+ZDwm6OCQGqzN4AhbuMO0gkzniRqqh0L/+WarnadklQWeo05wrNJ/RI9wysk
BGU4xu0sRC7tgKGXVMQaHmjG555jXZPnh1XGWeBwGy2eHK9PzclDNWs7qS95RW+IY4+rHkxsBUmA
hAtHmV3IEAkz3Ionq/CA+EBMhgnpZgU8F/dcxcq7Ty82TQNziO94sGOv9qIVgQlbAveqMoA0k7Eb
cYYk6yr7mU8Z5ukBddCIigACB0/Pgu3yDKWl41n/qZAbEDWNkkTFpX7iXGXKuJw6UnrigNusDXOI
KY2NLNBjIRhON0BtXJFYpTYp4YVb0BUyA5LzYS40+iJlMw1T+uZ1x5+rc/WR6qi+UpN0jN8+f/Cp
PrprRNzprSv4lMegDDF3EW7/WYpava5QlKPMt/ybo+qwEgKRinRHm1cwaTSZv9KdnleK3n9015zl
47KAL/IPik6z3ZcSQaz+zywhba6OejxT6mQXKwFmJMP+YPXl+zxiy1k6ewI135Ux4m9uzF8i+yMw
zMWFVunOd8Y/uxFh0VEfhR+RHXF6l9IJki/MOfcG0JGXqi+ixqEGdMssbaPwKJTtPprmKN5pCVgr
SDifUdgEUp8o66w1NXXYJgoGTqHqcKOPT1Wv9sn//CysYkflhd45bEqRQANgs3Knp+VYZQRmdwld
mW0ZGT7mOF5Zox2pK8e4b3LbZ6icPnq2SGZhgzLzePvC22aTpBiEQQbg+/G9O5HoL3/UaKRcGF5c
qR7YXzfThHOA26sM+cSc16xy2mAwll8fkyNW0qUWN+eAbe6kNn4outbdXm67MKzSClXJwbTtOwDJ
ZnIAXLfJs3S6YA5/ixqMFRXJ5kINDH5k09fm6i5FMpuVJ3BaZfG13NItANRIvRxngVYo+QPLF3+X
dm5234uOpaSM3iJmAfX3OKI08OvvefpFrmJUknp8gGG8u/wqN9KYnj6hBJ76ZA58KqgNaLvDWizP
hOHIG9eP19dfV4p2Fp49yM8AHp58mnrSA4zKGtt5dHQshhHNsvIQryW1tNz+TwUrDXnqLm8Hba8t
6cSZ+huqbqE+GphFkMI1MJkjp7U9v59mMn6rh4UtUH9KbeYy6gbmDJqMrzbDy5L3dzi5+P/fxvDX
5aJXB10HN4AcostGLe4NTgUxh8dIIfdYJhg+eBh/V47KhvGeNH1lY0SAEwzaoAi/G/yjSDH66RH1
5jdFGxV4qxP0TrdxW22kr2byYy1J4wXxU8z6AhvjoPxu8q7ElSTruQfMwF+bOl0DVJfeqSegsw7C
0E/AwJkpTajeBpIdIas8jEgoPJSm409Vst2CYn0u9edDxoPGwtDd76fpRvHxK2RwoAANRLruPRaz
MsosuG8AC5ZrbLw0KHeihrlrEun0ZfMbPSKJ2ZYt8CrGHLmmVJXpXZ2Y6tzCBIXWpVQcTPx6foLk
B5qdVgZaoDG4FNAKA+e1SeXO4I0FHhFKjPy1Ldpd2BMlVZkWpC05mhq5SxWGIqXxWsV/emRcvnhh
whd0JDHBKEm08OvavNl0+6WaZjUQ8Gi6kkEQQgHXI1I5Ymi05vChcZDEhM84WM8Sx8Av2NpIJQY/
ptQp1Ji363+2+uXEI2ewvFJ4aB6D1Wl1sUdaQi2Jvp5K/nc2B4pqcvLatrpfpTypv97XYjntzZLg
WahyUuX0d1yCIv+gOuDZGrLSJgQeY3N/QO0NkHHwrUj36pZXF25AFg0iCbjMWb0VaAtlt04MB3Yl
PHuWwH6+BFwMZDCqYMG9jiTGK7I9BX6T0LXbcLfhZ0PS3RFZCA2C4+0ytDILabgkP5bZ+TEfTLLd
7IerCCQPCpW0DS+fExHhMjnD22vA5e/+rveeLyyQaHvK1yWXcIWLQouiglF93DPQ0ZVZ7ZoZqiKg
ditB0bK3z/18e3e4DFbus6oJw1gd5P4IWQWAvfu94+ci4DN6MPOCxfhf4Lxcyak2ezRDxTfkhAoM
oWtxbiouOWXBkx0VzJRGyPUV+h7Vkz2IWbLuN6v6gP38Fn3QH45IPOvzHlYQb9V0/LwmnFODr+/E
wN1q7T4qbPPhXy0Gg5Hfp7ciXtYdOb3eYCN4PDhg4geDtIlSnk83kbgjxZYtZ8Uvcwhw1Hu7i9fe
NEm9F3gSczYc1tJWJ9EXuAhegn/WK871ClmCW88J/3/UbfjyOWa0sSuTf42mCORk4FaIa1+X0BWm
tkDhrbODt4S4ih+a3oxa5zg9Vb8bf9nkJemFBw+ET3fctYK4dOVE5qVztjloobRCk+qEeLMIW5dD
Yx9gCXmahTsHB0uAkSoakOkr1Y7nXPB+x9FApo8yhyhpOxhD3O6bwSIBZUFzQvIV+iGymG+91xl5
C6v63Dw9zJJNF3HeFnrH2Ri6kyKscvFZAlCSi1Ni8gL+zbZ+AptgGAsZQvj1TpnmKf7cQPmDeGxP
B3/BOzr10TgjrZgCj1vp+ovWmqB7DGbNQiTesHfx3OuFx4T0oGS+azBjAcRc2Xo7n3ZGDG4PmgLw
rfFPMwAz+HqN4VATLXGcNRMed+QjttFyXdKJVsaA8m7VGz3YZAGv62gas1RnleXIVs9D8xNMUF6x
SziCfyXGihAa1SG+Ju1biEYfiiPczvCtPuTYzp4FAf6Ddxam9wFzuhER45plBVxO+3Ofrfj+bQcV
8nM477Vd5qaeeLZUS3GitGvAMXWHwjglLj9J4eAkeiQ6EFh04JyDwrYqPuMl7S3WRIU2WnLz7LAs
973M+ZP25Z9tY25EzAo4y/JK7VkrE6XW9vFBFqe9aFORam5Xq6LLKOwU4kqR91TOkDniksx0rVhp
+LhqUQNP3bceyAmG5SnSZLECIXeLv2FfLd0vTwg1/jcc7U/e7g7Gd4RahfRdd4y8HIvCsvDp+kMj
q1kma45TGHOQ4ar/zOG0BnAFoD8URjJ1vxQ2scpmrQrz1Vf/ys5lDBcm3fk+b7hWkZkwlKkEHc44
8Mw17o7F3mF10B56w9oo7SOx+o0zN96lT7nMQ1ddAvSj4i4LUjxmQlnetlzMCAvANI8WUue6+wK5
Bd0ayQBScrxpS3cM/Oo+TunhrwWi9tR7X/UqbR4MtuzQfKCh2fGGQLJoVrZ77EPxkNNztqNvzDK1
G9B0qPCSh2Q0beLXGBmx6hYKdAzCE1K7i4XvvwgCSLHpViXiXDIbEKJP+FndgypEv/EQD1EglwKQ
0/XxwV7XR6Rsjt/piejGHcoaNGKwCLNdCcgmmm7Er4CUIC2Ms8p/B+p7RN6+lY1fGvbDMbhOfdpt
DwiquSSgQBFuOhqbkD2meZ+B8VObQY11ZEoucPNTkPt3vY/64wevLm8uWQwYrpFXbeG5RDQlrrrC
Msj8d09OU/p0wsAzppQNcEK9iaBh15ErUDn8JlNMSB+D+ni7QLV/m+8JBJ7GDX/ccQ8CN28Ez8D3
qYYuTveb1C3yaQa8YXqfHOrDVbtI+6OOdGsv3zUr3v6xZXnOQkpHIdvOP6ke0ynMWB5sujEA39cD
jQuJeqze9QIxQg3jZaag2ew9h3N0k9DDnbSEe+tU8uDCQh3f0Yhvbjgnv9clVsK4Wu1AKACf8GrC
+tErDHDn9OoyYBmVF3Z7SXwr+woZhBe9/qXhtotSMrMAST2T634+oTXJrkTVhM2iMMiuL5YzL5AS
rNfvCMNiN1iUCd65g7Qg2Ya1SLDmd0d8dM4DEyijUHb9PdiMirMA8XMdos8LQTzPb9zgyT+RRKe/
NHvEOmmm8gja9Et4ixJkytkXhqVEKbkiDw3E94bsAqcqaPi+5qbE20pvyZd2iAR+k4w0l1rdwGfB
tEz0k+/o/FkG/arCUhkTUKi29aVmLZTCAxMVQ9jNZImE3eCBB4tR6bNL9iNHunHsPXVoVDjzbSvj
f+3EadfNAAovA3GdC7fo9HjBvtLvudx3q0+Rxh8dIF9JcrisA+Bd1efkbeLNV1288NAETcxrk3ui
WABuWtV1axpZE9aJ0HAUMZPWpCmO3UGkdnsiDPc4KXOi1KtKSNQdokY5bF3sqLhwVXCp29lyOq5N
Oq06Jw581nhEdYabpFqTqmlsSpF5NmDDQ9hJ/xD85ZSRRENQz8KnrqQWqycDadX7cJF3UQe/hUlJ
hqeXEPSN2Mt1c0+hUunVXFKvs/XJdAHw2C/fWxUlE64QzVTaE3Yj7WBBLVEEVeYfn6qdprZE1QA8
Q0a/YvXeAYbH67nTFkae+11WReUArgXgQb4xrlc44Av7z7DzP/WL/UeiD7N8UMPaG87LaYx8MZB0
KCbVs7sexKGL86CUoqzzCqA90QZ/t37HagnHHbq56gye6qIIWuhvGbPMdrdHeDfdUGZebnXnFkXo
NbZxTeUAjIhzAHaKPdkez+z+ljVC5J7+F77hEgUXwU9i1+oJAntR2yR5qguK6kd62/rjRqoqtjDO
cjvjRcGgebNzu+6quZqVxu7+MNs2FU0owHj/TWgCiMNcjhG4R38rvY4YuovuEymlA+jDmwj0SxC+
vLj+C0A0FBoAo25qVdF9WTlZj+TEDavRI/TIV5gzjqr+zCr1IwTG1CJc+LXBOTrbKoTpMWv6W9Y0
sKRhKyH/WN20uFZhq27jKfDQl6yNLRDCArTSAat8okF+NJALXBuGWhUFfYP/diwLIc/6ESCY9sm2
H6+1RtU4gMukquLpVIIvYU5M0FF0zrNlFRG16+FyHRz+6ljXxiaLilqH8Z3mQCuCriYElnPIom2n
HJoasCBFxSmw3J0wS4BaepokbtjL9HAtvnvCEqSJrGxYSLFFr9P8u3ul50HtyRuO5F3eZr2DJdKy
wGjEyj3J55mGi7N4P8ui2wrxUnOiC2lG1f/eI6SOnTY3KpYJQRGRlQmbYtcAAhASmS5jY7sn1C3+
5YWAwl+HZOXwnCO9VI6hD9+cTKtBcdyZ7V+2z+2N0s8CeXlfm74VH5QhYaQxc0m2ptTMkSrrg7Lp
hB11ltWwWU2fCpmjhKpIp291bQWxtrVSXtuReci58wHYVHHbH+3G5gh62MOSpzuGtnDdCltePcQO
z2vAgDDQsYYjUmMCI2EXk1mtf2Ky/YQ2taf6JXVNq35UNzJI338lpj5LSYolXRPrgMngBAa2kq6b
CwvF1fakr2wdKcu6uF1D5zBnZhHcZvk7OBDvUWD/sd8Uicj1inU4SuXhQ0lcH+cHc8BBPGPyJAhv
MxyucMotfnPj9nktMNmkbPxjGi6uGyi7Hq+8osm1AcJRDfeR06nILlSD592INFx+kZkWs+0td9Nw
hEK70WN3vPINRGQH25mhTBTEruLtYh5oqdlaCj4JSqnNJGTNAzVzp4zN3I0GdkCdcoGtYvXYAZIM
ohzX1fYqCYi5MtF55n+xXw3DrH+rCfkNxyfBpgBvVEQMTlB4a+yMyfUI9MP3HeHbmAIgtbUi+XJv
N7jVXyXU2cS5IGeOEMqzw+Pmge+K3EDt/9OcMPKHiCHntsJFHV1MMjFE1Emp3w9lms+0wYZNDUV/
Jz7WH3BnPKjJ0cO3n1xiJNlfrScPazz0rPYkL/FXKb+O9OfGT5A+sgpK5Wlq/UkUiQsp2L7zZYKO
+B4nZqM3CWEkl0ZJczodaSaYOsQawVD04vfWlSjpByJdFfFkmeN9m7fg87+Ze0xZ10PngP6lPHza
u8Wb0K7kwj3UMb/Naus0wBEZ7ZKaNyGXK8rd3NYFIsFgFbgpFa31IgdJ6EJG1iyAh1nHHR15TvCc
kaT0HshKmzQPtb4IRVNNfD3MFdOOFTCKwtUvQnU9W0yDPG6jUwjcbEeblqxeQ6Hzzso4LgqUhfi2
R6x9nqqNcEvc7SubnBPwnI7hHvuZbreK90e9Pn667X9jEm0yZCKm+e0rBTgVh9RYeGah36HlJiTK
7v9wbU39SeBesseEZe75RSjzufDp0NleOh2Do2IISxMKW+Awth1vKeeJDJAIxhxYVBOBXVpEmQ+z
l6ds9ns8SnB4hueqJgELDWCfrWwRWloQy8v0Xa4D2I2EcuAIYf2nW/mHlpOyqJVzWxdeIJPp0ywt
nLzVthxkPkZOGj3xk72O7IhJD+vz/EDfEMHExNTGnyjIBQxjmYaJy2q3w/jpSPH4bexfP2/UjoBb
EEeliw6Ya8NKDoEQkmxHPkS9OMPRQS2RIMHAS7va0mHxZ3+sCnGmsce7hNnBErzcr60zzymzKi/v
KBXp+8qtOCoAYt6FBhFTZWHTjFwtNkVExRC9L5QS7G/O0yoJ/GEdE76+oMP6G+JR6ULxPSw2r2OP
TnoTV7oNAQzTDcS8A5AidMRaWVETyGPkF/53xC+dyP1M9RNMgr3Zc82joOh2FWaQBgF0o99mPb41
xcuFouNoPLMuoSUpclUPTVMTwc/t5sVviCdfYiK0wJi03U2AYZyaupuR04pecHds5HLe9zZjnpbO
yNgtwgxgAE6Ei5bZkDCK9TnlzvrwALQ7h/wpT7O7OmqxRcCMBXmHx1RvvYkGy8Me/GFpkajcsFrd
tqVeDFXQzY7MgQXEj78fFW8NbWWOL7TeFfChprhhkGWJoegI/Zv509YstSHmXwP4yZzJePBQy6nH
lJJxs7cuAwx/SjTJk54EA4EojiiSS6hT6twMIYrdn/ykfUB2y254qnxMwOpw66fXtxSNpBmDaIdu
UANRJQ3zFI9bksrdHDAbQXhQ3iETVx0c9kT1v8+jOTn/80jr5KVj9LqU4znXesLJ/ZwMW4wi44u5
mqeyr3IEEtilb49tZYVnRKRC4053Sk012wQrKL/Wbx7mfAduCQH0P3+1kVPDVS3AzUDMBLRDusFk
h/lRFjBrCm9J/5ZYriCeDpTergBvgdQ1eeZoYaqT08qvc973VE5j9IlC7wxfrA1Q0iUgr9leJVoD
G4uehlyJekoW4u302ZT0AI+RmEKIZKIl0BHwupJpzUg/bQ7idbE1/4hUIwxrvz6D0L75XAsrMMvm
j8B1cAJDqmQH/7yXp5nWRQ8LB2chWoy4b+7QN5syhtNMp7w4nFx0+TAkRfRf5Z71YZhfEQ+7PgY4
8sbnFdicAVDLCTedJera5xU5hHwX3TMX/VfWQ9LHdk3jQw3NfTh0FRcwPKbLqXexqV1alOoa7Er4
xIoOs5AAGzoOtW+LGr3F66sP/elxXOjkvCcAnbo+hiJ9H1mVgyPT1b0DaIZkLwI7VM9JXp6bYCyf
O091INibbC7VK0jkDOdsNK1InYTnLJlQyDL6a4ccrQH1NGO+OOiHS5dcmhrPjQmpGA5osiDJQgtc
z5jSHQhebhJi1aoSlAvlfEoQ9kT9Y6fK/AnZVOHnhcxzMvqfwkHiTWkuiJtvM3hfMgsVqtRXDOVM
z8F7ZiMokXQbAUkrKrsKvZZ7lWSK/INAfIa0sv8t0J7jFlvBpnZXkAYUjUBECHE9z6uo14WBwwqJ
TWI0lf/3Tw2ebL3+UXWBw0R2cEjgRi1zZwo1Qt9FoYvwsclS74pzhiFRYxfQufDbBgci1d/cj9UR
QQVsjFeu90lq4dODR1Npy6KPHuDLuvZGOcMN0eITpvwNyPkZ4DXKACo7eg/O+XjA+wkrFCKGpE9f
NT/e2zDxVVlqnSIqDbzuoBYprycASdan8XvXvUcEQOWOOayjofqFkJTfwaXKrGtNfifaCR9LuDS5
uOLiJXtiIGNdIW9gdWhyN4Hd4IAyVTEhTs5TYxu7V7ilZgdqzKXAiFxuByxeJnhC6g6EFSvKk8lM
JB0vzRpb53+VZW7iPEGttxq9XH/JCAATr+0ztgU+3Qz3YcCDUtH0qd+bqpNy4otwLlLt+301KUhz
PDb+Vbr21RPL2XgrZQkoHCM64bOICrwZrxDBwnFecB/oOw9eDrfpJxB4GgGvtenhqI5BflbUxcTh
tqaYLE6PSXX2VyNA1KCNjcyiK7FgerpIwoxOgKkN/iDaZb3gyv9EnVeEOJruKJSRXNO4wcDN+xrq
w4auJgu8lONxQBYfyvQkYPVWSWWknUQUeX7GOw80jt/or/dur5g9OWObjIGwV0LX7y3WTuxGj4dw
SoOSIP6TAvOmQR5zZCNgZl60+Jw9kcKxwIb6hvIsW6HZnGJb/072hTw1XMm/oKQWf5grKtvCFfoQ
Jswf4cN00gQVARs73W+2ixUNCWn6dRk5ui1fXlHkjBngXnhwGHJrqfVq1AY6DZOUpnWQAbzz0fGc
nx9McCPByt9O0wautgdatdDovw8YaDul7WEDCuCmg2Et4Np1zz9PodaF1kE5B3fOoKPbbzLULzRy
XYBk0Y1KNLSg0pS394JdWnLwxh+K2MXz+WKPKwU9hADECRHWuUVokMro4xznlNc/srEDtUcE4hj1
lqgCRj+faDbCV+ylEdRINLuznKoh/I7YHDIxUMUdws3uL6Hi2ayOi6C+mSmb+cSZkp14lX04ffYO
E1kl3jA4uQh5QadBK7EbXn5HjI0hH8tC/b3qgc/z5ib2dYI5PdESGahKJwt3cUlfCujRtVhJKUFZ
FeB6Jfegi2Etgj6ALDErdH7rC47nUlByPUKp//wYgJHfOcOXf146Zl7GqH/BTAgTpUJkTYBtRGMy
5UiuW1NVZ4SESNfmXW/S5aJDsNCBNtgzU1yAfBboGN6bRz/xtlGQUwNpjRZX1LVgWKNQpBZChlGX
pmKWuP7+bPry8k48Pq/L3GibDBR3B36e7g5uhrQ7Zahn2ic5v8dUl4/iwMDrro6wLN3u5HiWIOGa
xO0HBvV9od31TLGOAWXjJuytKC9WB18o6UDunCS8NBsXhAJiLyfq09/95L+PNmk6iInV1Xczetbx
RjFQJvzwqU+Mh7d9dzwTBLWwR8ShEBCibeDM1Ejz2P206q1bJkou1R9bk4gs2lKhWXVELqQR6CGZ
JtI2RwP0dbBubPMqAXCEv55w40payMyrO1pCt2se2odXqtIhl2WAQKlSfNm96ifhLmdyCBhVby/p
zTiTHPTRWfl+NyYG/xDiYCtd6yS98+Poj/xjUdzfpE7gOtSZQmyQdqgmlAEyuyvI6y5UuZGIvF/D
qQcXmBDfHTHwVe8HqU9fK9cGRoET+K+8rnD586ZCbtKPtiBVgerujw5ydE8tAN0yHh2MB8Tmq0B0
evh2gJp7GjxLmSYTqJZ3PwELaQm1UkLtGWyZh+/rUSnovuxvKNxSR2IjdmPjATlGj1Ht5LMdt7B/
8RoDjeEmwNSCIbqRmZdLAc214J6IYTr/csEUQGSdLqyfZx5M9oC9Iv7Rvq56t5L9gmJKzuo/26Oo
PXbJg1nAi6INBvUzmLV8ggyroQtEMzJnBucoPowWzghjVu0jj8a7P3hxxLmiNefz+6OnmXfdhvKT
cl0ckwv4BCm+cLGI310Bt8qtUuBX1ftN5VtqjjsL4PesCH6C0+fC4UIn63ai51l8y7PI+1iWf6eC
CRHfcT54NU80+XoQT+bunK3xw0vbqQSAnhNfAAzyFvb6DGKP2he6D/QdKAXgMuVCjMH/4a2n29Du
j6cscqay+TdGzOYnXmCu4L8ylaTUyT8TARSG0xTzivfpJmfesxW/XCTXbpkkG4mASu2lvIhr1XC0
D4aLrBqh8Oo/3OSOMJ7r4ipIZV92mU4FvEwq+eFJT/YN9Z0vmgGCCY8rrC5++9T+yJQJhmngWKNv
/NZ9anjxEbWiNuKpQWdW7igfuITMfleFKYABoAbef/4dvu+jnrI9dZNYoE7pfQe3WW4Zpn+t86Dq
xWMA+inHkJf8vDbOjaJifftH2fXQ1oC/DKU41PDDb27DHGkpE/RGQZAI89lVEnoo5kvm9EfRZ9dT
3r1p0VBKRmakrGEw6l3OJUo42iWwyoyZVZUFf6/yGFDP/nlJByhWj2UWNQVLIC41MmtbFukuUw5o
NmjqaAb6mUf2g3vi79pTkFL4wRN+cecpIHn23rr3xAc1n63zn5JIoTWMtUk4hEaesjD+JVo1ZywS
4OrwVAnY/Zhj0tzLxJd6faMXgmfCJ7b/JjBIDetzlGNIVJqPefHUlqu0Tl2QHWjVNtE7wJTNPYLd
+ziwO/DgOg8qLnYXUGgKkCwarEORpvwglYFxQzWsMS5QS7MCEPf8Qfk+SPhoyxJbp9WCMCpzQV2V
vEA9jhKdgX+Hu+vpSwBGkF+J16ungaghJpR+HthK3dETvFNtbmXFizUwhTcZ3SLAqsT5q12KsCi6
OKxwKKx1+PMttoDSx+KoSYIibb06UsEfwUyVKUieVJVYN/VuLKFTs10GGdWSFbqeCgBUPVEgm0mM
op7PyyDjYChfyjbuqw3/acQFIMD6q2eQy0Ed8OwAtokbcDwHlR1MShubqWchZvvaeHqtRz1YySv2
wQrRLga8VH0QA6efGF1AP5I/kBQfQD+gB0SILoHuADT0QgmhCN+lgODhw7otdo/UBf/MShRP3N5A
IyO3fnFjM2wwkjE9Dgsd297xbiibMQegqhmLiKnJg3e7m7fo+CsePNGmoTPCQ/RH1jbjhQ8YGIBw
NflnSgoTGRZi4BeHYIkrYlMhNzwcKqEWF8fcFCoXDo32wE5+jTWwNNzK1BDwGEd47uMh8HrhgO4r
xVN/LQzGk4h4x2C3Cp3ys0hZ1rSGWQ6pCCvkNJ+3IHRUccaNssL70FkELxZ0hj4zbrGflEImMpBU
FberGpVZUxomaE+l1f5RMZOULKuN3/EWPAOaVxSDuMan8m2+ZhFX0rRujt1o9gNsI08jEPz23yJJ
nlLXp4oYsnJ2+CipHt29Jc+3hfJHXsUQjJIOM1Ad96rI8FNPkR4OsY6jHMCxB3rfeh32TaNUNV7t
RAAyH2asoU/pzsMhGD7ZniJPnBr4LXyTXnWjMg8fqemZePfdoBVJFgpoBm/MAfsfC1ZLHGujKwSb
pUVjWIuxZgOVrAevnkTamcWCB+XtB5hj6V0OyG/ooHpCbZC5+zCH5ijzw34esP4M9kPBAPxqq3W3
lPe/rfOqz7HxqBVpqNjooIFl5wMDkA5+0wVVOqhxnLG8V4BL3/NbmCsXa2a/npfLwUdjnbslW49v
xCCI1EeuAINU4ZzS2rCuyapFW9uKV8AClyq91/+Vw8UJc/3te/imyqvseeaHvGCPOp75jUXgqN7a
ypinyv/ErQZ/yqd5JamN4og+zeZB6aaaUqRubNQE87wdz3kSn1WwO8VZpN3S++5wgtMuOhxVX4Vg
l1934ATP8+3LOIebABBY9ynViARW3L3MkWnX7A5R+0Jw6BQRhXyoVj7PnTnSxaWw6EKtatzwWk3T
MBJHTJI66sfJNhmCBn2c7ttpxJrfohBKCc3ijON6uc9nmhg3z8ajPS91SjuOSy3rcHuNi21yqeG0
u8nEDme5my40A8a5gYzqudIeMT4O1NvIHakZAqhSW0R1AxtowBppYLAoJD55KxhxxGuN8VrZRK8e
ZC1+hx/WGkc9CX/owo2oibt5ap7kDFQVdQaByGLLxNjczz622e0bHXp5nmmfQxaDgupvSazwDjg0
rELBnB8wtZweBO8RoHdTXIR9A9fAxs5GVIxDYs9DkxvsHV0+cTDv/jnjXZhGkPQEZiquLyHCDlV+
2PkBiPcTRYiAcesmXKS0JO224JRwdLqLtga58J/FAw9+FxjkuaaJQNdFk2zmhw+868BIQ6kmvK1g
ScGU37c4EOqR3PW5qxtDdKRQZQsHV0bMeJN7MBpURT7xzIs8pBn6dg4MMZVitzpgi2clLXEWq0c8
B2DX87jf+5tyhCwwhVkbAaKXIY673N3diFHFXI/z3HMpouEEBj8ZXcywDSntuUCrCOnqeUhjiTs0
1Wfm1JBEXkwrguSmuLMieS+G/UnaTU1ZFWDdTsSmQfpI/prABkEbDJz+iMl+fCC3Yl7l6CqG6plZ
JfMOmJypdmQN9+o88fcscFKfI8icK/Td619DrasOuLamCd20b8wNezS9l8vrNMiglLBUWMEx0sWl
X/Jql1JVYF7tFDGhO4BFERCPIKFk3b5xnsEda66zop1qNNyOi/rK3p6Yn7glRdyhgVnVt2Lnqf4o
bLpAQ0YmJwjZInu+lSg8VqxzcrOrcGaeX1HW9/QIW7Qa1ghQHfeywRh2qWCuPk4Ki3u2KP1LckbC
sm5U0RtLkr6G6JoE6XumyUN+cJVAHWDegoOBUNQ/JOOwwaExr3noJeSZurmJqhHzMOqkobH9dwf9
1klLug5usEJvTfGlQmNy5fmMK0ThHrUuOQLqQvv7uJeUHB2EvCZkTKp3h6m/ApOUha1nrT+AqAMm
RGd36YtxKyOHOnlbG40VYfbb8xmAjrNqaHy6P8IQ70u3Nljt1D0af+rWt2wmVA6Kl/UTJapbzAnr
ymVqzBR6I91aYQnXXwyefuyDlNshpO/3PvqskvFnvXdfs2SxvsShp3NrVbZNXKGbocJzUacDKtc3
VqZaL3JwC8FAIHqn+q4idpSY0soypMkJXhAgh9ZtlSC32S/E/tnOEErGaqT4DKPOdFxejBNeCrDq
hV+RmO7emCO9JXglvPf1wouwWJeDWQ2rIbddlXczvY+luEJyaCsUpZN3CM2oXX0OhSSzqIrWVqrv
sCm3es+oUvBIY7DYhAcfcSgvz7VbUla6R3oMrRzCJb5GgyOluOz+Zgh05Z/+Kb9is88L7nSsnSZP
2TrmrAOWQ/zibNt5g+runfcUshDzTNXYosWCWVCdOnmwTHN11XkqdAd0oybgey6P3EQLABb9YUhL
cyl5CXqCu0zHJ5/91JhLcGukxmucA4BackKWKNvqQT/l+va5PQ96bjAiJvUUzoEXcbH6J6jGVaOy
uQrO3qx/KyBQLR15AAg+OHrnGFOTtS539pom3haOB6p+N1icFRXYj28AlyuY+2GP3VJJulEZfLbS
q7SuTzvho3HbLhmj5B8nFdN92/N/Hix06oagCzGHbMwN0DbyHsZx1dURGvCPwusBTHf27ZoA8cuk
leo9qZd7h++l0JBbjS7MoJ4Uz69vJ/NuzgxjwLJXfLniSDJ3fAbjMRMP4eireFeu4gIQlPl2cxBE
TW/KEnspQT3uQZ5/Hb2vKiWnYTvXDtIdg0LQ7nKCTVcuIHnWjod0T8KYmg1GN9F9DqE7SzkECvHC
ZJJdL26C8zJHzelLnPYyYo/KFSPcnQIvQs2UWPc7cO//FFaciTUf6o085j7S4HBkSgNo0Z1RX2Su
pi/ZjZ4Q2RlmDBmWHUGlvDWFQgfkktkAnL720cVbFx/9kcIpeVC/NoK8IjrlOvx7H+ELyLmjsY4/
1y3sH28NLwYeIEvhcfQ5KWgGjHGLqDGfIaxS09lhP7uh4Ng82RnTjjXV/MU5GtrmrTscqp838MzF
9MCSzZ8BBtliDitxeYDgRsPZ5TOxfUdZEq/uQI3USls1ouCo/7UOk8ZSnsECP8Kp4IXsYVz28wMh
dsKqZiXcoF7L8+RGrT6qfjOrT4ZgQUfIyi/HtLq6jy1vCTdd2+tD6Q8N9ZAYd5cMv1hunUzU1Tov
ZL/8lIDEfhhiK2f1EJzONSPnWQtg2QxyihYpoGu6gpIPPZ+QiUx1cFCzdu3LSwH8ZygfsCwrTPGA
RhuAAFZM4W5X/LuL5e8vfyy18KtBE9C1H5rZgPNJJNLpSU+6NxGwGsn6IULnazoAcqpeaCxwlSs3
hwExByQ6nkRBaXAsRn5tG53NujJHD6wndFngghY4ufJKJ7y3M+igWyhUgRBlRp1scR56jfoDA0Z9
N2I92kL+vKK41yhOZ5tZ4WvSJcWr7qqse49lZYedHTOh20TuYTQaMjfy8tZRWnuLTv1p8br6XrLQ
+WEE5fpWewurzMHiAVj1EsAkUeqDuEjPobRXSRg+SR6JsKCh16aY6/p29ZEBjJVIBarF0X1GfSZ+
BmSICR9YPIhtoY0pTQNf2om4gEdd0FvalZiUCTwDOeqYOsTyZ0FsnXcBmewii2BVmj7rR8xtFCLL
uNDFinp1bBRB75Hjh6nw7a+xt08l3oNbWx5XSvLcuRINQfe1mDp6xjOaF91DpuPz6RZusOEsZk8n
cRWKqjVSb3ViDpuweIC3g+lVEwK8gX9Lmsp2+p0SxiYzHCTMBFyKMUBunE89yH448IpBiiGxMtKq
m2bD9eBnMFo5WYUjpGpWPNKfQOrnOmGDqkLdSBQNaIP+2oFrsBXwn5UbnewJ4K4KSFD+aD2a5snV
P3VysXb4LTvRDBWXRD3YEzamDTa5vPXySJHEg81LesQ7o8ngTmS/8HPuSundaqTo+Zq4nWQLMV/s
4FTLGkv5j5gvzjmayh7Q8ZGOrk2ZW4pEI35fvHTUi2FC4q18zHtJhwGKIIxAARLX5khUIHTaMfx1
3HEvYOu280Yc2+H8Lq0JmO8QxtG5YFWK+d0LKnczmjDls/SmI31piwbGK1SFknSILVC5l2iQnop6
r6kNIISmbDHv74njBQaIQo5pLWeomMOJ92KpxUMrV0t7auzDQ0jSXQsM+xgPLt9OoZKqArhS896C
wOEJ4EOrB5Dm8ouqdGQmLKs2SktbHaM+/r4/PqY63DAHpaIDjCuHfldiSGMl6mmCqtWRLQuqsNAo
FzL7XDVmim4DajKUxtKXK5BBYcNcgCDpTR18Jisf69kUogMj4gpQV2fAi+u0cM3xAGgS73mQ3Dpl
IJgkmzeYcv2bdR1j9HK73gYcS7AkqPPSsi2+ydeBcnyWOxgJmd5TEtECA8xkCvIpFoglmCbQFngY
MMNIccX1hoQdoQfqaDQLthJpW5IWI1P4E1lBWO9qIGVTqwQmH9C8QJNkCoRbJdGLlE2X+hN7t9vJ
FpTGJpqqe5d2rY2lXOZvdBRpIXRK7fTpZZAChJZLi68+g1E9c+UuWoOdy49fcNAF6Ostl1NHekr0
aMFZPlh9Dyz3KpZc8CjKb3nwhRfBhrJ40Gyr74dKDnNRAli01Pxs2AVjcVLh0XdDY37vnMZHLyD9
PbyzvFboKS3Yb/Zp4/ERKdKlTr6jVhCfxhhPrJx0ESzOKeAFiQGqs40AnXZN1/VbqgAQTa6VfU/o
ONeuUqaWxxg58Bm7SGknMOTY8zas7mM7vBD70DNSOMyXkQ1sZ25e30xmiQk3xyjGKHkjTnrhI7ph
ouCQNgLMhG3FIfJPNBwSDExBRCf0zXgY2CaB7I4DnOuj0/7MI2Zw867Kgpr7PTkru+C0spQ+TtAH
hflRJwpSduUafvBn5KeOLHvb7QDe1/23y0Kid5hUMUsB7vN1G4qXBuQIl9THl+CuLkhKlwmOnZBJ
9t7ds6mwhpgSn/XchjT8zhzECM2kQdQZc8o+quYEFRwOsC/MnjQSvJwTYa9GUYAHfLKlC1D5QVRG
kelQ6WhmrjiMSAHbwSTAi3UOaDFPu0XN+J2FjdhgVi4WKSyqzw+B8Vdg2RUOC33XgrAn91KqBSG7
095tVz8i+pWvs5dhzi+d0sNavXjE/TQna6UFsskNWsxHFWYj6OKkYRm1NR94uzninXfceT8OAo3O
PJ1S1rS1ldn5ZUu6G+3tgjrEMZkLC7yWxsWZ1va1FTbCs6iU/4g+oyZ6M4lxg9yxsi1qpt/7UeT5
lwlT7EMNbcJ14lYWFXZN3xlALQ1WYb4SuIDV8Bb9zVF+65iBNGe/I65oU1lHz5lSreCn4+RXp+18
RWcNiS2gT5/yHGHCCHUUCEheT5yEzL+urjOLsUzHOhuyYXpWhOzyESHm78FfYJiBXghjxwTWPks1
gi5EEMZNeQRrqcFEBNxRs6V7vorNeLYXvvvgsom6IDFhfipsHxIGztvFzAbD8MJimAh4AY7F0HdH
iqP23GCcbA0UC+jNRbXXDgpA1Exry1r5FTP+2pir3w/THhdcsEuawl/+Mtpqka51Uyyhttw2Hu9I
Cfw76i45hRjm9tD9xBxC0aJr5J4pD/lU28ybHy635tEsoKA+7MOykZV1TMTWLY6BqKf4ILstkLLe
UPmXeOpaXUPjg1lovaIJjM8LgtR+TSAAWxRVkkcPkUw5RBU3/QIgf+e0FORovLHxFhTYYbDm0zCU
whms/d2HWikScWYf+YpKuwQuS8SXmQpCKzvc4z+Shd+WNUYBhz2gwWr/Uz9I2gKkcI2Imw5aYpH4
8awPE65MOkKCh9Ee2uYqmbZB57NzfyCHMm9ZIEaMrf4qltor9ZSHB6yJeKwiDHRf6gMWtHC0FCWO
Iwx9O9XOq4oq87rb/MuEGQ/bhe8jvdvzWTiMZswnIgiRnADH0BBoIdsuhnXrbm8plx7sY5s5/TJD
wU1A2o4Ure1W+uQOJGvdWX4MsoxJnB7T6YrO8r6Yk3cs918pNEc08Cdj9QTYr9bTuetNiKE7L1D9
7G7ILRLvy6TSxwf9rKMQKqSRmYG+cH2/GKN3TPSUwk63rKR9LCAfdZhDtR6Kb/epu8ivBUc0/Y+F
QxCj0rLmZBy+1qqVYy0C4RvzG6OiSxfNC7SVTLUVhQvh8DhISX/lOVy1j9qgkajAoSc1c9mtUDvS
RvV6qPpo3KN2ZKT4ABM6k6uFf0lwuHRys3jiQPXU3dLdAvU8hWW6d+kgQVeCmRgbvVg6m4SYvfK7
A50esvrbVg6ELogTRe3NNUR4VhtCipwxBeMzsYJIBTPRAMPG7Nbo2/lxc2uxHPeKAgcL8xejp0Hz
45rOn6TNO3www33cNIN6nWEnZRHYt36Q/TWfIQ6T6LrsbRauxxyjdEquszJzKNeMWAOffRfNtkCJ
Cpgm4uzFo+35VWEBHTvYCIzbQIOtUPNUt5hJM08JF1l9/OzfYS6Ws/uEeb5zzCgk+M8WeJTVUvQ6
lhjDmkbk1Qnx7mz/Tthoh6beCm4KajwicwX1HHoEAFp3/K7c9Avl4eEBQXVUwZFOu3X37t5lbrwq
afJyI0YSLTt/AtwzBpi1+Nr6B0Iwr48BftBjbB7H0Y+NsjEYkQpTDkryAN1QWxBFvcEZJhHBBSFm
A7dTtMuOSRdH/Vpu9xVZrgxErqNqa9OpJohV/9/kyeiieBDeBbfWOhiPt/KtjQDD1iuZJxUG3LDz
aFZOK/OG1LklqQXrsb/eoSALzzjzdnfBWv+s9OKs5qFnAFCsi4UAm5vsAlUot8WC13LPU1Z84nVD
qI5srlpnG7eyhVRlVlAaISoKF+ixf1e+Fac8iTn7Ibcu9nhL4J3SJ04MieDBnWGoU8pJlat9+0im
omJDyu9hcS2Cr6CxicXrASql+yE9ZyZx7fCkb48BFBuGXqg8I2NNSnK7MJkuu61dAhnDwqazhvqs
Z8yLx3hRH8wofuD9tda3aSrW2TW+ClL7JlWOPkhbGny9ZL0ca8G+Ij8RfqdG0orBy0zafrfnNuax
ArMRlSri6aeyGF7C4dofhPnQ12QEmf7U8WzcBBkgT5XR0GpGFvkrvt6nDwKrX6qLXWjd5sXbMhvH
dtQluwBtQt2XjHZRi7U0Svzk8kNBjUHMukIjfTwFi0b/h8+Z2Xm9I67Z6iu7eH6PLQZl9bQCGtdx
ZXD9D0EsMd518kwVEKgFd8hWERGfvnK12uj1dw74hUem5kzbbcNIGcTkl+qoLuBfoUDmDJTuJsXQ
HufYX/DBUpHzIXXE8ElDGIMNylyd25sWDcPjrhhdf4xGGv4I9u2LNvf9RzcBnkdbAbB82EPsXeMx
nf/wJqvYj5wL9VZxNMl7fSjN1sLRAWEYobI/YEJvxSt2TQ7kMatr8kjies6YeQT2AsFNBeSEBhdw
SHV896HmJwV/vWc+Vxvh0G0UqKPLIfJ1g4teXFiB9HecsxqwzLwA8U0AtCpUFbsH8geUJaRRA4cL
Xg31Eh+gA9x+lHGNjGzkcjXAtsPg33SLFGtVljQ5HjPYGolHyIehCL3qNQtASC2ka9Zh27hOgDk4
1u0XMNAMGxK9XkKUE8rclS+PN+UV6io2+uSDEzMburhQlFEuDKJ/bi3wY2k2hcqiNpQpk9EYl/03
OjfFAgtQh630zzopoGLTrq+yCn2spAyvGIpziCkCrIH82lly3o5Y4mkLf7+NRHOlzwd/G67dE2IL
/Y3FNDWLjWKJSBFqTAy9gOrNgJK09M18UFVv/07xT6/B1/xWu7q2vbN1vxge6+k/c8SYWZuY6LCc
EX/Vjx3wblb4a5c28KUlqGlapY695zQTpm1DKUvgHN0dXRAECbwvDlIx+e3vdSsEqpl4ZiEsXCIW
RHhn9TXFv7TM+mhWGlfyUUSSs0uyUd+FcMzNcm2Y0eQ+LFqn6zoW6pmFGf38d3TVApGD8USapb03
jX94K/uvgE4JG6MDlpD+AU2o8us2FnUPiWqzJgFEQczouzm8XGsofeVxJTd1KQECsn23CqBa5g0P
Zo/aRsO7Rnjv8HZCYHDepbKwUmopWEjrDEAfVaFTVmHL+XluEUpM86sKZUz1Xic/49sWxmzZ/gyG
eF9/AAtO5z0ZG4h98QG3ImJy+ue5l9v97oYvXrXV2WGNpMZm4BeGhceTAZGfqn9FDShIXM1kloCZ
qEZhgPnxzcEsX2EykuscrCgnjfTJYc7faKR+9xGImlIUT3NQGfWUmhDr9Z1OTtzTotksNefHVaPf
c5YWhTtAO1sLlX9cnaeAqRCfNjMEmkqMBjS2mpMl6Apf7axeggqytfQliDf15s+I23H7FGPS6ZCL
zeWTI204QJiOkpYNNEraFtS0CTVXyC4tbAwsor7+omY5myFAYqqRNYZsHhFW6BVvlItwYrL4k8IV
9xOBgoOhNXCmpUcwiKOJ+jhYOgEEOYWLGyHQ1aWH5iK3+WO2Z+tO/JLnBsKsQsRnhQypiRExcgMn
b/8FUFfy8DG5CBAkORlJETlJF18ybwCpmaUnGVJe8iV25VqW4E78ZXHgzdCG1q3krzpJdEsmv+No
9QTKYIeCBd7seJOHvTgOiF+ZuzmLmeQINjY6TfrOXG0zfOpyskBRN+r4kxPiKbiPmdjvypl7m7dt
qO93HrKZEW/djnY0uURGOs4+s83nOIbxRvFAvHkFw7lVYBikbUJsDUWJRaqzaQLtTFsB5tePM8r5
81LdhgJ5wFF6iJkchaHLaKFM3utmqHs9hHRFhFzR8wI8o1GE
`protect end_protected
