`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
WFww0Nub0VyU9R/TPiMWDmzq4wYMmtU3revpm9Tsh4nxCKDTvGnIBYtUklxNwqxTtePTTS+ukj1W
mV44KIDWPOaKnmGG/1EesJQcuXWhwLBKcA/PHnrPrmsUQPD69asqXRWQBHLbA0/0CgwJGnVrayaR
v0g+VDyjrt4Yk/HoTw5rsfj2OnXS+yoCArXX6mwWHOTNTrkYoYI6K3NE12JTRYtchexWBpbWpzSD
/J7LeLoEX16kbBI22tw9HCgEJbgt0yx2EBv6Vgj1bsRu4VFs+9c5bmzhBscCmNN4SME/DYhY8BbK
rVqnMAivka84uU4E0E1kbuitG5KT3oegN0d1sg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="OwDkCTRGx7xS8IZyfogpi+GRIeOOccRJOrbzQoMEqXA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19344)
`protect data_block
bARuKIkMH+9jPb7t/p+iJDo2Xj2c3n8y7F0fHf1U38THjvtme336YK12Qj6nwwcHzFJu6b4ihT8h
UTqcuK9ym4jV93YkjWWz9StyX3G2MRM6LEc24xJVRKzBJc1VvQkTaNrHgzourMkwGvQ3aGqDr009
jbjnV7Gaah6/eYncrs87w4B86zNBzGdEVZeg64Cf+Wa7OuyJxzfD+hbOUJCzerYo7+dEOlXQ5WPh
hyyHGO5vWgcPb7oNAD/ij1yLXZtoYbzaJsNdWAACF2E8UwrW3feB5gTdwmKzkwCTNIB1U9+ke6st
cny/ZZF0FSRWN+eze91pElqlj82Z4FgQ5GFQKXHTPv+LoI0aTm7WhrYG0Reul8buzrRV7mWrLY7i
DywANwaylhCska/9fwCw1UFccxXLp9U4Nyzy1eRHheMxGc/Q+WSYYtmo6cdeyGwzJTfn9tT2SFAg
5HQl16/iW4Kgzd9fWqq+btlGbd1YdK5ynCKClP+W7VjkFe4ZBmZgWmuFKGaqFX0CEvhseiTF8B0x
KTmdJ01cr/irkzLUXZQhHwM6sZ2CGtpIe9VmaDevwJTv7CqnxzBtJ7Eq8PHXOxeRL1hr3rLoDqny
Mbn5320XnxFe8HCYgR55QSxunJ1VfxF0BOaXxw4uE8K8uGbUupQaQdDySQ6dAyGJOs4VrEeHfwSH
ArMqwHzrWIWxg8Xbied2I7OjU4oiRxk+G1H4iQHw2+AnaoUQqhl6RgDdI5pN37M3ZITbi72hz396
Hf5C0yTXdxWh+jlYuxtnbeI+k6z/XVJVhSho6SAmyh82klP9RIKOu2HSq5Zm+LLcagKuc7tKsAI8
B0LgB8megz6TndiSVUtflfDRyx1EGgdTaCIw9U5tLu7J9fatfeo4fn5VpXEns1MGuvHTjfrMnhRU
+gfSdWij+ng6AIuda4OdZNLuc7nPqixPuLotdPuzixkcrmGV9+f/N7AM7+6U9UujNEEFs7PAHcMg
7ayde+ejqHwdsNto4gLcXPTPdN+/2zN3MKHWALYbLMMemR3U11JxoIUef56d3h+gn82872q5ZGGN
Xcjf/ED4TtLJUbF9/7xe3DeYyPfc6HKLMr2ffgcSqHG3kfNk5BzHGqaKzEuVMOesT7m4i96+q5ML
5MpYEaPlY99k8tNa1nIxCe12uVe9j1Q5djoaLe3gZDkHkSLcaUbuJ0SbmJ6QmSBvGiyf5saTkYGI
X4Bk4pw3gRtCZrJx1/7mYrYCYORSk2YA+C7iGscJVDEZg0yXeuMMZ8k6N3LAAfJKFrP1B8kjxhsa
noUPDzeizXtCuOS9s4W7InjXvQKxxi1Ix7+oVLvNbpnkvRsitUEXrUmarnFiqdzIlkHzH8f+V7YC
FCu+cNMyhKLjcdAFNQSfeinsTqmqrQNqSv51DHySrwlNSQBGBvd4Viln9LWYnC4GEsVRWao3wIkU
5PK1jGQHXj9G0WPZvvzT6Q1GO96D2MiMuWHDIiO+B+xW5uDk9+0y28qCwie1P24rUTgI9dlk7Cd7
2M6MPVfFFjHsoaDVfT3qSawkUNRUk4ELBA7LPNhi/CSxyOGtpoAIQ4E8RmXsukHzTdcoFKl6+Tgd
aFf1YlKKlaytbUW5+QvXTdc+Mnz3E1nt24O3b8RFWvAyEznRMPY8ToIvqewU7fa6TDorkWphxeua
xrzJh9FJJQx56r5qVqpcZqP/l0MxSF3nPy51uJtnIL1hJmFBZazyvjnK4PqMainVLsdzwmGripNI
PTtDDNPaJK0ijCyyw/mRSuNlMzZI+BW6iZZCEnlSiecBBQCO/i6+VMd89HjPqxywmR8aT4Lqk+XO
CDwYXD0UB9X76tJgwkNuD29SDWEVQBxqV+NbMSkhTYUOngGP8rEvQN0OTsYrp8Kv2b0fUpcFPnjZ
d4OLswzpgXlod90w+VnzKsBzAL8XpsHfXvlU9xhmKVxYkDeaxNtaaid2KOrH8Q8err4lJwZ7jT3b
0COVy4b093ZP/5Af5FRvLy66ZSY/xpk5njlM08kH2npDKUgaWqyG1uDS7kWwtD4Ks64z80oFk6dW
jguwwsKBKhQNuU7bp625FgfmnSy8LBUwX9yGoIvBvh51ZELGb9G3TPhFZ4sMUZll0bbyTsdbYBL+
qtnLxanhlmyIDO8pcXmejY9AWVcEhrXcnRstqZBHsn9/e+SUwEMfVhGFy2SbC4XBKq1eHa+lNo4n
j+GP71fHIWozd8INQIEQnoG45FkncJR3mOq8kAD862i5DSSUNQD99f2d9jRs0Xwaq/FY2tlxntzv
geKzTAiwXt78ByDqwOcoGz+gFX4DocE4WK+4/XkecoGmFr8PG+t0zoYsmGUgpIs8kIK+Eo2Olzr2
qrOSjzNlIQ+yVrbitfi8J/X8ZSg2Ajn9d7cd5S1KI9ue5CS7+K+Lw8ifv3V6iWhYPYamtqChMLST
bZikBvBtQIQmuk1l+wot07NSa4FrPkUf2MdJBsKxw8qFgJRk/Q62mEUcDBzxqp9Fm5BGhgTAYJjb
KQQC6NlffjExt7xv9kok8ETf3yiqUNMFgEXUT7aCAKRaI0JucI8Z96rLEipiUJc63S6Wle4veq19
ggrfiselHJDf7Eu7I0zgfQ6VNZkMrAvxpkpnljcNIo3aKUHSQgQx7tCVJ5ycuHTFZh+zEY1fFpmC
Xn7LGNtAlhQTaSIriJ8hUl1KuHpFDK2GvmCCkZOslCwkIq9fa8TnnjIiDQoYM9Jy2nM1FngM1VkT
zUev3QiLliZwhxgXTydT37MhhZLrF5dDFPFB4OEgxU2GrxP1+HECWQKNtWKC1K1pjDUi+nuZNpSh
BDOPPYNxh6meEuJMPMG9cLisKcNLVzOPmeunL/UmjqJuIeLIJyd/DXfsq1pLyVUJEpgobJdwK0oJ
1aRnj8L2LV5ELdveuGiSTI8UizgX0F23mh5w2imc7jlf5jDIROo/7akf7lNREHkr1xkhyry35wLu
aZW+x35OCnIFT/ebx038nEU2MuiRtzCCsXYh4EbtZnJVFjdY1MvlqTsXqJye7LRfLrjg0HpUzP6/
bqfILLimC1u/b+DQfkSVXVp/75SK4M0+lSfitbFrTCoP4V4gRvcKYQZX+weTjMsFWU2rRSix44yD
e6LL3y0dgXdQ5RCgLmL3nKkroNEAzZm587xa+gnByifzDTKUnTDkrzvFrgNwwgdYYv6YBMmVVx0Z
bZ3N//xdfh0C+6gxA1N6obdZKAI8HuaqI3R1trhrt2mxCRvBTLEOkhmjwelUgwxPGcarOwqlXDoH
nI8p6BIbpL6CHzIeMtleiBgybIzjSYszyLqRZbsyrg+UCQmyQuwEEq+9Yjyt0IymuRSuiFBFVKyv
eFPs07P6KDZIGkSCGsT7ejyyjV8GkHX1bPVmqu9VBtzDxegS6uggYQz/MjQPJMPWuymIiKea62Fk
uxuJ9xT8ZdY1KHkoyvyOE3bMMgsEeegvkAT2aVFVkdVn+EMWH+QpJA7z+LBxuYcqOojfJZGrqEqn
Yr71iEBGF2Ow5xvYAwsOsy8WXDA9f1G8NJJiHHNle/yGSiZtoCFfc6AESaY4v9QMAd1+sSooEGbC
QxX+Wb3qQtmx8sPpF2TiRFxU5aTsP2aVUqveYZt/OBd/DuMn04mj8I+78ctIETX9+HKXaZPF9S8L
eu010g4cSDE8aUGH1RNJRMtFSPOcbaSwd3bca8tyfHDhRznUvYjbsuPq9/eB+S4In8Hx8vKgUHiN
Vq3Ygffz5cN7ZVDEYPYzbn///2ekGilvRKaBLb9lefpxJCpKej0Iq6P02OZWYDmhjJs/9JBoFMRu
/kZQwWNIQZ5pza7YkehkZhiALT/vVsautqHu7Ane86qII7CZJE4/7Q99sAgMz4we9NqlpXD+6Z10
0v2YuIttvAPnuvLokh2IWmJ2+A2BnSU2zDgLtSIUUMYU9ONXzlcPAsOAxgiG7qWtctuuyzdYkSky
V6TyhVbIi+b8gDiLAx3ulA25glKdn9UrNL1LHkQCeMuQoB75sMDSuOeJv80SAb8nU5nOtOJzeX4T
5w7L+LIeaXZXthbtPsOqcNWms/iLo1KBqmovck1aB++xPMo9+hV2JDhl/wCqrTE/VBPq734GM254
YV74VVrEhhUhRFTssZvymczzy6i1O2b8k6mXiUxdF2XdHgq6AaKYVlgNCRFzMwgADom3v54uRqan
/myhZzSveSrNCVVi4uCZpQNLMc1K62DzSIV4/45EB7MO56undzlvR8QSLGdqByg8dQU6skLrMoCr
mw8wWDXs4t/MZCs6sphXNmAAAHOkYKjTH08cxSI+D/SEPtWfTFKd5URAZ9vNmRlVRBCOJSuxeU06
k0uvr7iD/9Hnm8HUN10OhlLlR9rSl6jB8caIewqJ235YjnvAeWM0E3n6ukKICrQROI6YaMF0jWIo
j/xOFvsuIKhNIZfvXyi/C4oArMEUh85J0uRWdRnRtzUN/AdFBejzNvOVOecwIzKWmXFnr43B7+wF
4CTh9+b0HPsXc2XU8TdrhORJRsqE89fqgwjTYw+dnhtnboPXL0DzcJ6z7tKWljsK7RRg3ROBEfEh
TPAG1EqaI6QQp+KrHVr2mBtZEToALEtSNFN+2iA1TH4SHhv0obBaqV2Fqf6W09SV6CUWUCKvmwDj
Ro9D13bkJeOOW6p+deMbpsksGAA1R9hSSWwXEcVoIFFyhdb8wHcpQ0ohVrEd0fUhfV4333lIpZuE
l1am6OPm/wFBmIKNh/L2og5rVmINsoE4r4sGXMupm5xLcVDEFPdqxevbxet6dPKGWZAVdVt+xHZg
w3jgqtzRFJtXKRQUG/09Al4JbYzOLeuxbnd+0fSdhzKX/1l6SZ7s1IK0NWJhrLswcT+m/boU0mLm
l+toMWRVM3toLzsd6kLEjTxFdzBNDm1WxIeBPK1depImougWPChuj1kChwHybz7DjpDm+mkqCT+Q
zdtRjc+Upd47t8JBepkAygUFDRVBhob+gJS8xWVrXzz4o9AcmjaqOzV4/Eiq9U/xU5CWLjTfgen2
h1hlWwpQgwIQAS7p4B6hIHZPIu4YfwZ27Yjo7T2fe2ABkqF4VqNcmetFXN2R8QsPKdM7JNzJ1lnd
nDOM2J2WeoKyyptEPl+vn0KvCw80UvJ+nGRCpuVWEw6cao87St5LxdJj10KU2jv6lUjTnocpftZy
DLKAAVpTdemJuYqLE12KdrsFbCxKWsiTGEfb9ev6v/vs++aO8Wf1T+Lf9BKfoEdMxJQjbbw5NxMF
HBZte4lhGlnb+KIBqEOPMQxqmjY37U4IwH/H7cHzPiHJGxOWirXagLT+Gb1RcSS+70hROnDY9Dgy
v6pHqSDfK2yuEhBWXlebxHS8NOrPYvPqvRM8BS1XG1N5TlNGpqcC4yyEeSO4o75R3OLQfc60w2ul
T58kZcUQz+NvJngZX6LCjg9np+r2G+9hLgZF/fOUSqWYzjhxNOxf2TGLxy+V9V6P+nrN97FbG02G
VtV1vjabFPTjKU1GWt5rmr6g6J/UPfgcLDz7+6+UD832cm3vTHCz+FQZ7JKX5pr5nQZbAom2fZBz
AnRPL1Ek5wZvktewADPeo/eq3Grn9DtmixFm1Krkcd+W/yPqXkqJ9P3GFIAs8cpbIpcu+yeniY91
QACxKFNNjkqcZmtvGNWSnq8HDZiFKUPJn6SIC6yQ+ZJUSw8urkxnrUrFG20PJGwPU37r4RA5lUfj
LgHkhojt9QvmBORpSNpoNExWoBRfIqAK8ZJE8ryyFXcFBTKsGocD529LRfGRUvy9L+yOxQtkUEvo
a6EQQwXV/iq0nu9CTa+tpXiAf+bnMzwRDWPs5IBwByuDpwKapmUA1nGuoh+g+7xF28EOk4l1rx84
xWllyUdde5diSZtDKWsMv+nqsbqRCGSbNBBsl6nDp5wGMqqejmKEhfwKK+33xXpinY+Vs0azXlQQ
FI+Ryq7vzwKmEc35s9QH7ikj7+WnQvz3TMUyF9q3UwYm4Znc9NWgj9l1oX9XhIvq3N9AqOfKGSIC
PtEQR5A5O5qWJCKB8gsK2eZxUwxBs8Mcts0n4q/TbGf3MjMih3gpAabiMwPUSezziBImTbWSrkM/
j0UD6BgBT1GvRI6EdxH3Fptb2keNEgCWy0UbvjvHpicDQJGt1y4GaldMEZ4wjg+6SUg7mjzucMvt
JEuFI9esJ/wsIWJZJKkXluQQYwqbNLW3xkrYNG10MKZa7+h/vPKAxOX2yzVrnp2Vf1bGgsNzi1Ty
zGhMtNn9M+mQLB/rd8OM5pMYYJB6aw4kFSc+Lbv3yKnUi/Oryl80/MT8/q+sqm7ydQok1rB/d2IW
iEy8mVhECnzP7YwDFI60IlydfHAhqMOJvwdnEqQdlXg/230HLa6/6kIJZGy2hdvu32ot1uSCk6Vb
nzV1yKlZdhSKLzTfiOF7miVCAaSzdsd6hp3wc4OZ3NDCNmNgo9b/9D8bziZ0K39qcpVZm3zMCVb5
uLYlSEu4xuTldj/jRsQwQKEb/fW0Ljpsky3/5wAS1MQnSmB49EfcBiUTZQa1sIzp+mbrr3qRZn4o
v2tJg+QMUoWh5vxnntXzwB9gZGKUV51bfIgpjHs/DOxwGIyqvKSZ74RgwojXZMLJAe9cTAdz8Tlw
z+lsZH60s0c9DHayNKoxYe18AazpMFC5RkpwWHRqguZ98B1pBI3LqNHjmFAQykDTK2r7/wsXiIOH
uLkzTQ62g6g07yyKBasEaomwY/44P+B/PKpFvhy0h4/mcYtZyGupSaZHhUNXhg1nd89TUGy59c8X
5jOj7VCCq1Lt1zreCxEynOLrFqNgN2T8YXoFc7gmerg2lP2ksimLOLVg1jx3cyluqwaiEfYzAkCR
KuCM6O6Ol3Ig7UWaWdB78wcmPd8r3NDuRQCkHBEhiXc6wkWQky3fuGCzGBRTTM/acSmndRm9bjCA
rcxFqXu6pXRY/4Jae+aumRyN6ZQiABKxsrbyhOB5agmKqehz3J9HsQbj7sQBiFJgCT3GhdeiF9OU
t+ZkE6V8lZWgItGpfOCu8BABU1zTajA2f5WetdIenYuuLH7GPX9n8khTkKoy22ztk0iMB+uHvUTA
wkVKoDHgYm3i0TYZoIy1Egzp7OfDYQ4OQJhHCog2KCRghLxDsH20URSwSipEaPsGg129F8KiYrqs
WErS1b7B2cXKD8PlEONo9AOD+WpztoE+ifdpZ2a5Qr9VM1yORAj7bsq9RPwY8ke5ExU+pLyui9Bd
p6qFq2iGIPaOhUvWbRSyrcoMKBwvEKsAp1KQT1sCEkMo1b63HrQISBZ7bW2+kisScOGFichz4K/v
yQCRVml0LlsLuM/zfxaeFpPta2w01prd2uUoQFW5MnF8rH8JD8Hf6QnmGWL+a0/dL66CJ4s7yrSf
0p++KhrTk1OBfs/wGwDXPTfLvh01blThByhuKvtiyym8rUZjSunUlXP3NfqmRwMSXhTNA+XHHD1E
zrWG+WoXhmSVvUuFNzdQ6W283xyKwREEbGoS8YovbVWmgcr4LT085VMNL5EEGYkg4OP8AAzLWbRP
g/g+6f6mGKTX7Jc9l/GOSG+r7fPa3nX/sPeAgc6UKbte/zLCXOU4RknOXeaUymhva5w33kDpwfd7
deQGMwLVDO5cpEvPmY1sjoVLzioANNr/4xKctWFS1DTVRYAlXQk/6dHEOfSKLDeKEWSyvZB9a8WX
CjPVmdiCSEcACmgTbOR5fOVixN8vwA2GTS7YrEIkwe95dysnT+wKWyM7glOztTinbpb9wMGQqr+H
r4Mi7qR/msdhjCR2ec7amr2yfZ+AZgScQ0zt7lVcsKTgEaRrIL8pFdrdo9Kajd/Q6seSfk1rB/J3
sJTz9CCJwvbrfyvGRg3zn3bh7KozsF1F/IzHKYhwTg4fA5aIyDsHkuLvFSg7ie5YRG9kI132EQ0d
7Ys1YWHwbM87n25dr9fL+Z+gCfYGLiJahnuSXrGwdmhkbYWbVLaNiK6sAF9LK/8R/tIM9GScjqEq
4s+QECvQqI/miFVLP/bE0jmY/Hv4KpjskhI9GwMpEzm+yN8dNqWCHoin/15bApHxnvxGZ1w91Zym
BJLqtkEHnHa2DMDBRNbwX39JpRfJBtC2nZ4EwCv8cvfScrRIvmBxkZGh8CXoHVcmzKVZSXhGfTOW
7dWVI9zTRyD/CAQGqA/XrFKpGfhZRBuz79mG1pqRExCIRrCgaq77rghpRWdM1IK+ugz+dP1X6OP+
UgwmxNDuNdpgPbjF7ZgwFQv41OQilnq/BMrz0aYdp+NNg/TutOtT6TVJi5dO0I/BaCfrlNw6KIBR
SbnB786qcWSK4saUFm/mYS6TB51EaWgB1A6/59DuYQLVmcf4SxVPem8gEF8b42wtVkDRCmajrFKA
zGfBlBU/moYPEHXI3jPcoOOROpRXBp122orYWXZ/0tCO2n/cM6VBcAfsDaZ9rMN4ii8oX5FKCILw
OdA4NAggwOe4m7QUt8n4JKVc2IYnb7jUPDVOVgRLkczJS09h7Drc5DqT8neJHOkm6YC86vlV+Alb
pOpnncMVdo2pwNxeRMcI9m5DbeizY3nqRMhxcu1X2vnnOowePyeEpCp+q5rWYTnzsz8kdZHl7bFX
6EkrHE/LdFYNige2OeyqIrKt6SLf8cJxRJNhDL6+AyyX+qKgQ3UcXKeOIDh6Tb+JXiSsEt5rXE0S
+xtBh0wQ9WTyuFiQs/597y4czTXhlmlmyP2A6EANWAkZ8EZlS7I2y+s64zpGj1JMZmqB1ifDnGMv
zAF8k/6f54ELb8j4i/+4emoQ+0dy4wa2wnxC4goOGHKaf7TNjq3rbWNBECcZ9c1B5fajaMP1RyRm
3O8GjsnHgMkAur70kpmFyIcQR/TCsBqwN0aeGwB3fkm5XJg8rClV0sWwJwgYpyzDM6+Dv0fJE2pv
mzVTuHezniyM0sqkT1jSPw72fxQOfchar9uKW1F9N4GCZYmlFC7T6vm/JGorLLil95ErK+581eNj
sdAId160XiRMJFu8gT7LVWHiCEOcUF1sd82rRwWUb14ZI4mkIpdPfdbJLm0eveSSZ9MgBxY7Aur3
0dQyiItcf0qA81viwY+JKWYk2fIMFh+tbkZ0K/pLL9zVn61lmean+EXHaVCPSB6rq3gKtOgRXeKh
nqT8wOF0n58OSrxQCWDuYN+9fxnrjgaLhiNJ98+QgR3O12VHw9oFbAFgV+wuRfrkdDWnBf99bwGn
2aeiiBmQSkgyFKUbGPp3q5E35oV+w/76G8jil7eZpcIXKbcvoknVx0m6wu4eJGTxpB7cZfi5Jchj
ZI+9mg9xZabdImhuNJkAgfrpad/GWACipVIL5vn4zcnlHt67T6xBaa6O+keA2ErnioVV0fWtlYAm
RRqTSfwSK3KjgdXbYWuL+pI8mpdsdcZeox4j3i9kB5uCyG4zOHiHCijBzyghpZ5Xlsky1Anf46Q2
WeFQPzOx8PDcdoICfUO2Y+17Z/KqfhwPeIwEe2BRzsPDT6HL0a60brxvBsLzckk3sNqPni+EHu0l
kaItVbAo0dMBesYnTEr2iWfvyF9Ry4r6iDXprGFG35o9HFT/CYDfvO+HUUQ0jXgPPZtS9SAy4wY+
rca1pg/pFR8OAA6HaJm+k73kGaYquLtc8skJt8BzOrNVOg8flRAXLS/K6ayfYpbt0if8RBtMKeQP
Ms+Kzdl1G1tuW+uiwfdEzJX9XUhzQv2Y4EnJ//md5mfd7iBQM8obI7XVfRoO8vQ/p9Kz0K+zaRXe
vjneb0+/hsZUlft4b5gakfw9ITZP5a2zvJX2bpIQXWwDGiHs4Sxk7MnWxf51sKjDNriAMjw4CQaR
CobnSYac1hQmomy9lz1NuXOEc1IuEKgJjr/6QULzSfytlI5OaO/fdJ+x2uUpMuHbiu9mPTwV6jOa
XJRc675L4SpFuCK2OmR6MXcqC/xQNxLxvcIqlD6al2PFzvtgJi1E4FWrb6A3fg8q2Eef2QLn1wJu
8/ze7dBqNWdpVlRY6yQGhBaK5NyWMvBi6d3CT8avvcPb/MYRFtOCR2qkq/4dimJsbCdxKqMcGO/c
mpdxfAsua+tHyNk7vJ4QYuU2UkAXLCK/rX5H81VEL3gXIx+Gknm6K2JNC72znlRcQrqPa77fDirh
cLLEGmSQRL/m8yPoeM92MeSmaJqF1MT4y2EGmK5lLSEX6OCVPWAaadZDqRv1z4cqtgZp1QjxBlwP
HWMQG+VUK7aaSfMJpTEIwn8xYe7h1p7QAEi0L52wj13E7nek+yv0J+KKtaDzIUZq6UZl+3monMzd
9w1nCPkUy6FjihXzAZO0Edm3ScQnVIzVgXWb/boGBnbxZI5icpQVt6cU99eITuctnV3kvRsmr6G/
qlK51kJVKGAtP0/eaE9zRcNLrZB+z+5EF69eIXDWaezCCI4NomSN19CjrPzny044xDr8xEYg6lRc
++m9+vviRCEWnQsMFS4MveetymJtT2Xpj0KidqFOoh345nW2/2mVuAKB2MtRktpaFt2Es+r3xMbu
S3tvO0uwhZpx+BjEj4PgZv4pyJiY185IXytk4T0JeO+3Sda+/GXbPHT5B0ap7ymvGLG69l4fUoQW
nH2qfBDwZYJGHMWV9IqFQ6p7o8bkkpl8gzXVectG1CbRSQ2iTVXb3adkgJj5ylDVW+dXmv1vMnfp
Mu+pIp4Vsose0sgaVyPxJMTUMgZLomC6k9O1N6HHuIehupK6bNDxbrDSfCV9zI2Bjm1X4BdD/lFl
qnEC3up//9k6LlMnUxlUNwsdMIUoX+u41UPM7EvFX5rlSELx98VLGwdmuribcN12qoW4ahg6rk74
kG37wf7wV246M/urvFpd03eVxi/AoPypvr4WEScJXuSlNVoMDKWRZNGrxeD4lw3DIe48jLDV0pwK
/BEuhH3/PIdBQyHaN0SL60WWGOR4LgTdGR6RcB9oPoDDetG3WWoacywM96luVxc/5pBu1W4Zpg5S
VWlAULMvqOFPjl0wuIRbFDhSN6ELWcimljSCjNe9nPnO8FVXlIdF664dRhUtK4M2d5PoUjn3FDqC
w8ZW636L+1WjshTdOkiseL2hdM3i6lCMMpljSj8nnKYuHxRnAB/wuirlXzXnQoZVMqm5GKOt5V9d
9VOe2ejosJBFtYlVn2kkkWpJgeokldYNgvslat15UV0J+XaM2iDQpHhuMhwOccxu38u9xnpcnB6R
3kqSYweTHEqJo/3KFkfa+oUb1vmD7H4LG+NDCvil25EKkkdSGADU/mh3kWmSbItqRihARVo0hMVy
aP8XHZ0vtHI00WOPym7M2kapB3K0653E5/dHtIrb7coZeveJt0JxAl84S3KB4DLONXKdzJ1Crvx6
u+RGXE1f/7hMfGMV6RuViiwMJ4hT5AG1D2hofESb3ArrvAJrYVG0SW6EC1V6BPJHA8O42QFylNS8
yBREgkQpD59Oj4jdI72QXN5JnF9SZIeNYXAn++zW2Trkyte89wrOUbJB2mazLPPkWrNtqJryEjHM
8wT0H2hIaydlZskMf+dLkD8OXlm/GCDIRf+QE4H/CJdDKiiPjmGRLWC+QWpmfU2wkV+JVCjLWA/7
Tyi4OyOZW4oBOYa3SzEHHpDR6d9ncJ8nuCXvDEhJNBcSkXSxzUztz6RPOHeXw6HKzfj21NDmhJgE
IF/sw7MKeRIue08DOdigXJ5gEWVVsBNTWaqGkHAxPn/wpEs3LFZDznXntZ0nNJkALGN6WbIO2ojb
O9PWd8J316iPwNPWV7oZMcQYkJXZfsWxeQHuV2BY9Y/a99Y8XEqljH38FPJHa0jX/0qZhTgZEXy7
8HRwsIG4xJQ+e8Xrl7ym+piA3bztOCuD3x8bXzDw6ge9fsWBKN+RT1NAAgpHBpUzdJYFHT3gfnMf
G1kthBa8JdBv+dVjejoX/E8PDK+/zbVUgtkg9ZMbqYaj0fVOM1czOLGbhQ+qqbqnqlByAgkzCZQj
mKtS5U2N9lA6l3D8fq4PLdthUWNhhsjxo9PfaIg9A0LxGqIcWU2l7CP7Lo/pDi0ueFgmXcNq/s7J
nx8z2FKhjKjjIpa5/t9PFN0JvJAirk4XeYgGUd2m6Y9MO3bQZMhaDJEqJQTe2cSk27ahnHI+3Lxq
wmBcCfmggavrqBZ8KVVFTS3WHiTBxLPKZEamTGpj9H4KYIaSYuBVVnzUxgaHejI4/V3ycmtyNO8q
IPbHv9F8NjtwoctJX2BgV72cyj1wwSrM2dqDzjRb5+g+r5h2xZI4ecpk0jC9IfMmwzEVSR3DiRGy
rOeqYUm+tr6Rzqr0uMpO/d09OvAe1fo9wry59ENcQuu147iLv65//imjzg3g6vB426ut6cHz0tmL
/Xe+anN8LPuS16i1DFnOLHYzJSC2YPlpKFs4PXW2zgKL68fqkPguXGvz9JA1zPpBaxJo7NMEepJw
yvdHNUgzaGiI1gmoi74twDW7aSr3OLVAEJK3wIXSHyHzcbdE5eRErIljt4ncagBrzz7Cm2Tgbi9c
n9ky4HiND0FcFQrBiGAIBiwhpr4Laafn9OKVQuS00X0E3EGDKePpfO+vPZFcG2yaqD3hQUv9nTvP
D3H1Z0KpN9AqYucWwYS57zbho9dcHOXzHE95lbV0x1XTpoIFtSDActHZv4/Jno3j7wLORSR18IYQ
dQyuARnkhQQLOgzduoMm3Q0EMamAK63uOk3Ql3ErLdls1IBJxCNTZyhCo/MlBmL3EoL6E7OiL2q/
3mXjZSyWfzd9H0aSSS8b1aQ5QOqyqrcC2rTsETX5j+ESZmk4ItsyIkoqFitYMiendK+cKtXjO8VD
8JqMWe/5JrYJlTG7lVRqwskPu4I0OgUoXNpsKc5wsvJiZqRnRHQu6aLG3LighwrHoqyPWLTKDzgn
qdjkf+M1QnwEHSCoyHDA0zkdrh+so1yV7GIttS4x2zKaiAxSF52usWze2RfsseGSudMcCz3CXblQ
ugp+w7CAMxbFGU4rzl0JotJZj34JkqYmR1ILaomcR6A7nzRtX9WfjegNtxw62NOScQxseGnVfbT7
S61rrAR7tR2Vz4Sghd3d0GHk8DP6K9BPFD56XkRUpB+LGE64GZa+LQ6b1DxQLIZK9XYLiUF6Og98
2V+tAfpouP9VJ9a3fqk9Pdq/42QnhLdDBGV9/AsG0+0gUiPu4SZWUIlsw8JuOKScJtyHhzj0GLEI
tEZknZIKI1cfvtVXglyQIKxt/4Uab6gm+FZC9Ije9EASmDpAKsddskGDIhO02OYhlHcy4y3EYpEx
kzb8IJ1em8rfbiuqU7jOPF8sfkcmZ3fahqzVAXeDPv6x3o5T7M7aUqjRnb1emVtaljPzxHDkwn3c
efKdOESpF0XyLuML52REOn84FN8+Cki8SqpCEjjPw+NPkA/9aMY9wp0H0WAsZqhXhXJg/qbPd4Oo
+ZvcDVAXmB1gd3diQ6csjnWQpj3IMqQQuz7W+dLxC2C5iNLypxj2ilJyR6Rln2aSgnnQcUAr0VBB
Y6cmYGE2sEq7um89mJ1qg+cD8ScEaCom0mrAen9dFCGGTFG3x9YrFiqQkzf0M1guljlGMFNWybpb
qo6dZJMcUokU3dfBFSjXrC5vYuFXrXR9UipHc3cwm6OgZ88ITAWBGBFppQfI9EI+USs/fJrhJCaz
kM8yW8y3icrTLfp53EiAkLI9s3fd/7vP34g05J1IwO38iPZU6fTRp0BKy0lLRkAvaWS0C6fuoBW6
pB1TGRC/eASsTbV2VSAn6rBu2u7GEVHcK9fq/5WyigCQan7JWecgDc/NmZXuriKL25FCjk2LuddX
6wLsQ2PKK+GklEf/Tfx2nsJ7J9EBy2HmWdDxkHyVEWF0gTIUillk1Ue9455vVLx3mCEiX1Aj//pG
Dzq8yz1570oBEAiLkeJNrv/SNLK0NNN+MlMy9oqrkD7TMTAbLB04aqbRas0ggZSyX8xX81J92rmx
bHodc/epm8w/hvJVqhCn9sA2E6t2sFIMCX7Q7zZcFP0g0dycdm2c1Ud1rj+qoWQzVZGH5H3MFDNw
+TH5ZOhTCJVBuQwWgoqOKOJyJA/ghd/UsxJJMarlHbpHhc0nEUJ/1BohJoFlB5PizuIWC8jqPSni
tNDQT/bdo0gr7vm+p6ZIfPkr4foyOvOgeUT3O26faZPM0ucD1RBr2V5JvxfL+uzytg5ZnL9EJ8QS
XmD3gbeU17w0KJpvw6Ow0fUC1Hq0AFeyPQrOphe/zw+vhvbBrNftjfw/wxCO6t5cTVFXDUdAtINp
vM2yOxD7BIMqjJx6QgFVrEgttsmCDM6hk5/BkXjYwzFhJNHIJDKC3q/E1FZfWJJrsuIsVVVbLJir
y43O2vNvhCGBo+sTn/MTWEV7KQU/xe68eXfzEjEBtNCaJUB+3jhPZtPW/zyYhwmjbbdZKM5FuvNz
QF8Sj4J5JWTE/JnML2xpTvaT6SQrgEhgQt0KgXgZk3nEOEGuZjMuJQzqbKxNx3J1iDBEqaVNOzZe
UGN4IhNBaDoqo0WX4WPuQNNZOYYNrc4jSNYd0cqSsvI2ZZgMzKypw1wkG15+s9+/qPc0+1U1O8f+
OwAQpfDXb7FORXAb9XXnos4kwGaeAx1aEeO13fQWyk8pUAceu48AE0XEweJ9W4kr3vnJ3AN/cGbd
016T8WQKpW7vsZayO8/t45w60kxhqeDLPAo87iUNV5al+zPCX5QcsjXEaKDNIrf2fSSC9do+tpJQ
japvQ8G9BdxZNqy9kgWkAXmRKSvrktIWAuZUEp8CPxQ6U3GOzIktHqlcKN/WUqrWVoF2r3KxqIdm
egpECPj2JdWZSQJNGt4MiLgj0EmMDyX6CLhEap7QquSdpDjLBxHAR13a/lKUvUbx7fL9RY+epBOS
CKSWDZcCUDYJISQOPNVu46lOhohxVTjSDWxJscJGmfGmcYl6qARADH0ZVSJ6M0fP7hnExyU4y76X
muBB2VyI0QXmj0vOmDhcyRvC6px+6KBQkfhrUZnkKGPVMji3/j954PY1s96R3t/La5f1PRSmdvtC
dC+vjAJFihEpr0i+JNGDdlry6jJWFhaTw+ibOcXUM9aKrXFkUT+3zEXP+WxuOvIXrm21c0qXb1dD
yDgcXX8WTQ3hI9sEgVPoH6SpIQEvDJaODfJtFr17shNUc24O9pMXI1O5OCwv+IHulcE9sbitzOpT
B+PgdAK7lv45OhUuSlbmTyUoOG9SCjjXGxF5fUfxw/SFjzQ315+FPSNnDNp+ucO3SZUaFDN8QKVa
ZcDZVxbUcwCKYLY2CpDzUYhykIa6qr8D30th2jQtGbsGP9xeEr+3cTDt1IJJN3yjeW4m3PdtIAqy
bxp1+T9AHpNVyIbWY/pamO2Vd2QWjOkzocwzynwJO4DV/Vr78O7E4o2Mrw44DYAL/q4M0Krqpvem
xWI/JXUjtKpv6ylop2wDbD6tA8/5g9yFQuxaDUrzOW0QzuLkXwF/dQ7BRBBlR6oj/+7itz/pMycq
7GmxL5J5GPtPZMGEiZmdvPyr1KzOXZMhIdh6EiF/bgnIrcLq1hOHt4kXhfQm5BEVRY2ObkE3wzS/
f63naQchajRX1zrruuOc+xEFgtGOmFtGoui/qkzXLZzk1HaVibjUEGSj9PTrL3KMWB295ulnHVqh
oMww4fI2FY3xCnR80jhNpivxXwj4cOYyC/VlTd5X8rNJtE+R9kE/c+oogSrMJfvnE0FM9/Yfa2z/
LZ2lQafipBJHVm+LajLgSi0+PKW0qJHcOpHYeeJUoa4jc2KU076ca9BTi7fNQUx6k4P8vQMU+pxK
AZyOZlL1j8p1LPUwp1FkRXWixQIys4ew2pQXVrO0oJRFLto3ZGBrr5lgjDknopYr2S4mUbnzehYm
OMoIf50LEze3bq1M1GTAZEzO3SRIECbv48cSBW0cMvktCO/56Wj7pvdBb70Nr434fy7Nh/Qv1OUl
3X0RqMMGYwvvLUHEYYzyaPqCDOvqJ4yfWXoSinqUKkyzOu66mQyqVeFMdhb1HNBqPLBIBZdVnzMy
1rgVqcGlLjv/Ngk110aC6T7FNtKl9REVih9AnPfx5kwJ78I+B7+naiIJ5XtfkkNLrrJRGJA3lNC2
zscwsNXFEBjytZ/S03NCx5hGYqOjz1vufa+zVt13CvW9uWUk+TXG7EfY6EsGzYhEDzSgU56tqHA5
jPlgbznnVdIHloDnWWTjm/0KX6RkkFNx31KeRGFP8mSC2GyHwuwtn16oUH7SGROjQl9dzvJiD2dT
CCnHO0hGd3wOoAvdey7i+armfqDbMwpew5wb571RQkFoEnfzNBJXpmT/HnJhBpiNXv3xcYUjRvZT
ZKAFgQ6rYV/YD0EsDkEn4Mwt3HzxiCUweyRt+urub64lIUEmZNBN5qsBvUrHvMKCAStDxg9CSqEH
bmVTzOuZ8qrh3PIF9XgkHV/3OXQtAVyHPonVhr38QkD7pOBQlkQkgekacuOzYgow989yIEhQ2xA5
wD0rVJaqgq3gQ0sv78Hi5hy7wW5TB7clFNcn2su8XxM3i4KLg1RY1lI0hwYTheCMAvXdUbuD5HP4
t1Wxhu36Jh2hPGCtP6nsKRqrcSJYnqAIk3I3rQmYOVYgp2UPfKDR1q2ubkoDi8VJUr+6hJ3lSi3B
XC79+LGtGs+vj4gs7UKvsiWdgS7uw39mNUPsguqhBne3Hx+mvRuDYlL8Rq9bWnJUZo3tnhCNaCG/
tP69qxxcTB3dpA3Hd2MEppZs5iyVH8FszPyKiD/IpnRHtKvhC3xBlPv0hNkEu0/vCEQFXQb+/iII
hNgiLIBs7l855ZjGMk/rVVoq6XpqlGASyRuNjUlF+hRNUfb5aBh5/zLUXK+T9s5rvyd7svlPUFli
TJ/yBUymy5UMgh8Pl3GN3mU4Vt7zefRAwxvL5kE19bnwsvAKUnoDNOCwU4/xFwyzEg75h7/mT3ey
N8vzHFOcavicBqGAzvJnKebYNQKjKspbV1Cl6MYhxeD27HSzBc37XTsRlbgXxkg8Ca3toHGktpNN
vL7HIonL1LMBcXM0RlHFISLA76Ziv2Fc4lnpZOZssCBUvU20fWpCro93QYkGwF4nhs4wraKXdSz7
KuuH+UOO4CgXt5M6cpo2yqsGItKe7xYdFxiHIlwmPD5hMu9Br1ZcVMliS6LMvJVwn5A3+pFODIYk
9McHtdodbnwhXzY9P0JjiFGYEWbrGJD2AbBCqehJc7pwoeEvOjVA5ckuXDPEemCQQgVwOnp0nBdu
kXyyHTFKVJc0K1mG6S2qiq1vLgo8eyiUGew/uuMPdnLbVh5yY27I9vcrP4fH+ZC6nZgjZLXGgmJt
XqHsqwffWgJyyybAfDJc04Uqz6IKnTa7ACHH/I9aP5si8fza1l0S3YlE1DE/tz3mK4qhGR8zLQP/
cMW2rvJ2xCaEnB6CYAR8P8aZEjAzo9jL8M5I06CAfQiE68Xk+vhB539N/lWK+ZCRAoWqL8InBhZJ
PUp60vzFRlK9v7N5cXfQEm9o0quzXwNFhEZAKrGQ4NacT8XFLPA1DQ/lCHilnWT7EQgfNs8RXzdn
LsvLPmVjRQMadi2Olt9kI/pWd1eOAdkIYl+3QrYe18XLx3067U79RMF5v+BdFuICYH0P/d9sT8kk
uzpbiQgTL+BmNBy6n1I3wE5Ct83Y+V8rKFeYMxoOvEfVbMV6n8jlvHixoEJvVfuMj0tEGBF2jitm
az3hnrApnKQZvF4JOfOn6oLW8GkjfSjIo9aM7Op+oxTj2DF7CpyksfdgGhJnIBjmTqO+U0a8Qqol
ADXHoewgBzexNbcRIc09cRdPFmtYGyqGNK1g04n1dGNwCv1kRKhjFo7MKLeWIrvRlhipUuyG8fdC
/mCIpECgYJGz80Lhwe0kdxB5POb0LCNTuLjllSCUED4pOYQxR5B1+qQxycvz+5xjhm137iyaAfr2
PP922j07cr5Kwd27IAgWWW+4frS693Fslq4N6iVc2wyWYq+SZWT0aoEV0Lwaywr3khLfRR7TNrmU
ZVV9hm7MR4v8UqLBlgxsF9jGe+3+qwp6SS043i3/40+Ag7SqfzDNkj9BJ87iS1jYhmh6aFK3z6Vw
Z/Ubch1s/GqgmIL3IZ3efsmqixHfTYkE7Hi76Ou0Afxrg5EY6cQdsWUkn1iCalCLrUvXELGYvjj0
8evBzbCbyh7iQfqpLi94exo2kQyAAcozxIXYBTzk8xvI8+NqKVFGa5k3GxRw4xwKuglp1DVfYDqw
nrL5ER7w1tFp3+iBKWH7fU+JlUMdx2FISV1v6HH/EiIwUOFh/FABnMVbnO7dcRzqHPCz6tS5ClXU
AXgS2WnzAmQxRuIXLQcr2NO4+t39Coiy4QkUQh4KuvPb/SleENkL88seMKLLZL8zRlirXsgdIK6y
3sS+V+36DtlOlmaR5bx2mN6X08kGR2ht2cZOL02byW8XG0VlUplwNswnOHFJ2k9BaOfz85jYEYy8
DfohW/ou+JXc11ymA7zk2FdKOPnCEdNCueYbCS0I8T1hkU4PJ7QoZkuhy+A8JiTFy00vIXLjjHXi
Puqx8mkOyzdY6aykRf8Q8P9zYc4MtO/cqZqzl1uXvx4Wc6fT+fGItMRyCnhw4+cabvmwL90LSOTR
qvxOosjwpSUJngQX6SCQ+NdWV48aSXmyTIIRYVZr73faIZPD1t1rDXEPLHnLiI26HX5pQ86He3P7
CIN9efBEQN4XVwOKwxG+cALgJe8/nmPtik7TJ0tVyPY0FynPRSNRmtkTtT8rpLL43PHgYKAusnH8
K1emAkeYlbqWhuN558f7gLBalSvfkI75lQjfDy9jXnB0E7TCyGmW1EkvVW8KXz7obAC9fBPJ+4OZ
oUasdr/J8D30Goo2imanJgxoUGly6H/yWcbDlQcp5zD5lkZCJZRFV2EEwLhvb1k07xkGkyanNy2Z
uW4Q0cia1eisBucCQrzZlw32Ra5Zvl13Egbd5IBUDtTELtYqM8m7NOM0oHRxjrGgk7fBXtGbBNzU
R1G/2+f3ExDPLYNtwBaq4B8aAeNnPKq5hPry4c2gGgXS3cD1ey4wF9nxxXIF79hPElpY8a95IGzU
QoJkqJq5mbYJqngwI8QDg9hCWeVi+xCDhtQynlrff2KlIMGdYeSDmCzjAAU9wPzxvZINYeqm4rEB
/5m1CL/mb9mSk4ud84YNDytZTNV0U4hVZey4yTyXOVwMi9DS/S41geq1YgJXFdpLPMF04iD9mdS0
PxcZbB5yVA3hy2k2yg1iGJaFKHM5cnJk7yeYHaqVOtxfNEMF2rpWlAzpTMI9/ADkNoxrVeDzvUa7
slPPZJBf3WSe8X0zFvkf1thjSjzEH2XZ+vvy2qW5bWRzu2sNssLlfAcg0nZc2GKvPGe1xOLktokJ
73QQnRCakumKDYlhL78c2MojNqoMLW7zJSadsHXcsU0BtxTh8u45W1VYTSJYdBvnQeeo8wcAFwWv
O6V3En6c8xFaZqrM4/fgebws9C6H+E0pC5Pepx2WF0a6TeaparnZDG1Qelp36x9bAjHr+1ifQSQL
ce/V3q+tdPdDAPhQ/x/ETOZ/tE1XKgQvP7KAyYxBOiqL90mooBtUec1e8NQDgbSFNmZtF7xsZynY
9GP5ME/OZulj3RXpZUUBr5/sagNbtDlCWpDgClrFJlG3dG4ANyXaBd0J7zhidKmsQqjrOZR2Xy4B
SRBQ2+yQ8XyqA06FdD56NnIMyKCGulW+FiCyetfUqja4774lsv0OP+cgz8KDLrMTCh4lnHIBTfGz
8Egwxn19aHad49fnojB98MZhjHirAGSpwuSulPbfSb+bORY3Q0QztdTMa3bkKFqOK9JWtUq7nMGo
ISs94tzrYfSx6Ry/JddHZ2JNQz/QRzME9UhzMwV89N+nVB7P9Oh/0dAJ95VKJXy9ONmaU2/ERWvh
jKnxGI9tcVrwayBx7kG6ZjFQyTlQxXeDXJHMikJtkR32SaHdIjaN5/Mupqp5fXgdcDBsKCeH1IYZ
sM4uFWH1DLezonL4yO4WE711h92WGo3xlBXrGKHvzPlfcqlzTmln0Yyv4aOiManWDJQXxvpOI89i
ndo67y0nsPf5m2vt0+ZXZl0kSCWO4+4cpoO2rFhYZP2CluAkx1aPKHhRDMCA7ri0EBMAHxiXn5wt
0cCRhU6CiDhna+Zn66ak76BWcCdw5Y++nxdMq8f/N1qNTAvIAadl2Ay0pXukfJOxS3ffsc3sbBNv
RTtOx4y76jCRcxTlgnpPCKkzlqUpMe138sW+GCbwPHKDVWngkErNxFZU7Ez0NvRn684Eh4cDlb6b
UpYlL/fHMuyGdEmsXMParU8OjoYYFtG6MQ+Y9UhONhaN6yM51u+20nrcawmt31T7aXk557HVaMkk
9M8QgOVn4gFLK7kkejM/UA79V5AtI7t1XQ7UbUuT8h4wuL0XUxW8PVp0ZzZtOmbR32TnWKcyjzNK
/LkouV4qhossuQ3cOtDBiK3te6z1hOq2DWUkYXWAufKkxW25/1ByH4oE6nTCww0jdYYOkvLlJ9MC
20xmU1Nf7xqV0nTNUiYCOL8/bphFHKpjXkvOGY2WvMa3Vqb0QBHBM5hPhNgkugNOyIZwPAyBTWZH
yRBv+O4UBlCdKyBUlXPoBreCAvb1elkHNFwDeSEPE3qK80nF9M7MnA4uLNe+ghbrBu5k6P8Os2Li
hiBWqJH93X4l86u5HpQQrt3lt3TEQCVuQIb9MsP+vwkRsgLX03tUagFOg4URwthX5TpZhkx8ESfm
PnREUGBxt0zfQ0q2Pm4KMGe0YOLcQIIgebmcUrcZcAhgn3Y1BpHhecIAzuh/D4eZ4dJC8dToj5AT
62nfMcza13+x16+OzZKoyyAhbFqkGVw2ZG4ViRg6xmtQN7xwOVywzq8SYBKaSqwMW8bIalALoCdO
DPXpTi2x5mZ3G419dMgXTzMd0EIMx9M9UCcz5Dbh5FXBW4qmAfOv4quHxAZQkrf32GmYJwhDe1tT
rdbvvuPpeRWCrdQw3TzY+lrK70p9CiQLhZxDfymweGMzN15SmluxL9UR1UAqln7rKfdgqKUmhVg8
Lf/AmwhgpsCx7zudoeYKqm19c85QgGQqj6HQ1As5ngt3cFiUBeqjV/IMeUrsTnrSVY7FYpXUxc/7
uWKb8k5x/Ay9/tbwVoQS8LiUiQYyisw4Hcq9qftCws0dF6bJeGVGguPgsUDDXFzEcQeyvJO6LpAy
9nUUtKGPovEcvziG4WfYy9Oq7R7pGeH0PwZw7y61czyXLvpO6iRkIUMqi+aTbPp4+cyspjSye9gI
7Dz0Uw9ZojJmvpD+L7cBB80Hl9VrvJ+xWGSJgxhD3J7pwxlCIpt54Gp7X9gdDXnzSzhHMgnSiYo5
Klvre8Glqiz2hTOZQ8JerytunZT/MaMKrx5l1e34HkWcseo/gGwVE+0fYhLove/7Uf+wom5SyET5
t/ZrANmFGqcPahE2kTCS1OwNIJF4rBeEY71dpSPlg2yL/p4KGjuaLuAlL+kAa8QlXkR0Wv6UUjD9
wx17I+9QzCxw91xW00BYgZn9zLqVY4bdnPaIEJfHMsLSuuUbLafiZEyjEDLwlMGavKiwkaV3Zq3c
d0Zd+1JNcG/gC+4HvNom2ilH+P11W/pJDZ3CTd6HQE0XeU8zyQy+6fjVXlNHSCnok+OiaydNrXiX
yzItUvkkAZZx4w2MAPQxSEghSkmxj3Gkrpa3JCAt0PlRttrDDzcdRTvbOEz13j93bDx/uHnbiZRP
DE52b22qLBqGu0/DetvtIaaHrHgWEbXH+My5uHqmByt/+qWqoYILqaA948UEAM+gYaMA7JyWMTZX
pkXfJHdc1VSre8wmafTwr5ZcYE5aiTKFJ3gNTH/QzobQrkVt0dgzo1cT4PfBBuW/7uxXltZGMOz+
0fdyHxX4GeNB5cmuzj1vnQcuoQ6xFZPXJeNPngXsHFXFqOYZnvAf0emne8r2e3s6jI2jrRF0y7Jp
u7In2ISqHlPfv2AYlnD/o/CLGvjUw9Uphy4fZsVUUh+TvNimPR7S+Ju2CElSD9YXvSowauh+MTdu
xxmK5NHNKfRYPyvCl+dRIUwjOQxYR+EefNV57tmKiY2Hr0guNCUaFgM9/Oa2FX42MDLixpBVGX0K
kAOyR3G8GpPpUGu8tUhcVmqcm8Xk3Yfqjv2HnOXbxUuIdm/iX7kEVq/jTM/y/iqSDvFHpnWUkerK
0wqYjos/FbAt/QlwwDzfk5zjumGPPFcCl67EVVp6cSfyRMTvBBV+jNBEVhjbddPJ8mh+R31kE+bN
0SWjObHVJ0D9Ep8QE6Iwn7tnJllveZaBndfIPVSI/TGTPzomUJAhIS6wFq1Mfzpx9yIWhBXrXoRP
ZifGf/R385FO2JggcYkSi8XrhNFT2ZXblLwUwI4JGEtH3YGzR7qit6vh2KgdCvHfHgdkTyR9G9QI
pxM0YB2Y9livDYWsZAvvxzShOQqN9s0u38inZNvwUijkvzIfD9h+J6/Q7722DdNEVDx6CyK3qjyR
ZX5Ekkduz9QCtYVVhSWErMv/KGhnF+NwJCR4tTaqHpSYS2qgRmzDn2pYki4YomTrtndtDHbbE6sN
Z2DBgG3j17aANKffkoFpGseBjV2iuGfLJV5dpGJ+D7L3UQAQTsvNUGrpy+o75aEkbEwanMypu6dY
pYvaRtBWSPsiX9CstuYrhTF6X5x9OJJfeN+RVmpN25MkXMgtQ57TEqBbrT915iPcatkbEsBfhQoW
IZNc50lrXvjBDUTUG596xISztmpO2sMdO0ovKaNhkMJBvJSGRpusX4FI4Klq4p7aB8q4eL2QdN6l
1cN3fOXPCIYMMFSGsWm1bbsri6vcetNnf8t8v9cCHXKUNYOBz95NpIYpZ0XdwzUDEBkcODZqoCLY
YpAUl/gF5Xu63WZt4hmtgAN6vuNwlmFT/cAA6jxqScmajYJpGcjDEsSS4dA763AfKu3srwigmxS7
cZ7RBGcpwfTUdPJMbjBnU/KgxJoTZoLnrjX2cz9+UIjRcUTbBim2c4P1GagFKKwRJ2nrO+zkBcaE
0wCdG2QENj+HtEI89+Y4c2cOvU0ODR474QllXdwgeDgWklIIOwN9Fi2iJU9k4xeKCndVoVwDA/Dp
V9Gaa86aKq2bfylFkjv2Sk2iDW5IdQag0cUUCCFTTkbtoVVBA0Fquqs22rvyR1N6uZFfdipQXnOm
3lgyHwxt6vB66Y5daDACdkpFn8p0nwwVZi4X7kKmg39wQkGcjf7H4kY3eoxLKcBqwEo/pD8sha58
T9F6livtdWzKFLi71tpHI/++NtMHvR9zAE3CxWvUF3f/FqlITIDAyQwLOCaId6GUCjGmOV8raGpE
08HX/AmwNwVZiATvuoz3s4thWtQRhUpYOQ4i8vHSnVK8y5HytTD1hwtaCLQd1QXg2CZKB2KLCOZy
05pINALVZyRin6t2ssIZRATPrYgjYtQIUirhhf2FPMrNxXkOW73FebXfmqGDelThtoEXEvguzUn9
6xrC8w9nul91CCWHr7+0Bmg2GVpaZ7ZB1uGV6iPPswoHMHTHCWnhYkhW20bmbg1fedJ1jYMIjwi3
mXn/oiQj+K/K6sj1WlhpA40rGW7BRU/BNa83W0/2BFA6K/1MKBibm1TKD3mj8OrywsM3HmQyIrIN
nEILfKp+jSIulP5fFFxFa0lytbVfh4EtmE1H2e5gw+UykeluaBZxwn8mfMG9S1NhIeIz7xKt2SDL
GUTjc4JoKiIUxyw8sbOmZ/eNXtxRlRSrbZ64szswAVep3eDeLG4mqnuFgqBipWe6RQZx2e6EqqVF
piK7xJovjIW9OF29clepyO5M8yXE+OneXuCRFmkecIpnU+bwvoIG/YwgLsCNNin1cL8YpUCmCboj
9jEx5a78SkGVWizA1BdEl2WAKeEuMeulpzrAAUkJYAkowI3S8DZG3WumCyHS3H/3Q5uuGuu8/y39
NEPCoi1pFbiz29VIvQOnXZQmhHVIaSSKBKyCTY9d3vrzHXfrU72e/fIdQUWShBD/Z0TYXI/4Fp2m
w6v0NQui/SOwVS8dKOZw7TTN3rrOBScQowF0ZCKMka2DvtFliE+GHh2pYISDrsacTVeg5KsQv3om
u9t+9Bq4MWlsxB9DADI79VZH8DNeU4m/+/iJVMm68gy95mEVDt3GGh1SuehtvaZGXmyG/oMV/GaG
B4pvnACFXmwLrbgccJcjwn3IwuKCEW4DveXPR1qeZWp8QHNuycllqQod2VlQl/9/wMrZkzLj76hq
6reUZd+GTA2sUpI+GyUstpHL0RiPZlKFRMOT9erZP5sBkFHQJxo5P4U7L6P+UvOXbNw+ctU1LxA0
JfYUsVyEgDhM5PryP5ji14FVCqD+2lPgWDR/T6BGASVFvmf4aSPW+W5NOXm05IT3D53mPBCw5iom
4d+oWf/WMFXGvuBo69XIqeZujiMorIwSqhohZpSQ3b2xjgF7LYw+kvu71bTTPUBq36v8TE8j3Fgz
knX0FvrnNjfJy3d6VTi9oJVztMYAj7C447CmsMcV4OXig4NOrQ9Y3F01XgUc6ZTuNUa0l3hlrK3d
nijpdSMZX1SFqxxjvqzHEO3Z+9WdUaaigVR89/QaCJWe0kzgKpA0d5jTrHlp3G6LuctGNg3VUMJk
N+uHupDLVy1nk/xmsH3TuTWVUP4oR7x88BwKnryADiFvJsFOF5X/oS6LHb8Im3/IVJ8ekhJ/3l+n
umThjx9XWUH8W/t8B/zF2eRORRWUbzXIeXxnzTPy3awe536qkPhLHAYIZets2lvqAEqKuULldUZO
LgeNQVfbxZkf8YsNPJW53L/TE+PytBcdKemW0kekcjXdZIHPwvc+ivmcmVq4Ixj/3iyaYai0Jll1
6x4FiZq3cZhv8TdDC0wKhSPZ3X8c0x27KCgNvie+5D9N+Z3PdgsluA0P+tHVyW0zk8YuD7bximKp
yPyGA9FgbnGh3W9u4w4i9Dk+uWwGXd0+EoexTQPTaGMdxAsXa/8PherzxPpWKh439+Cp78MWOYTP
nzWoNDrkKMsZ4wEQrE26lDjU6/h8WI7tPn+RqXrOWoA6Nat+dzxfEiFIAPAoRopiunuNC/ifB3mS
b3mPmEKikJLKd2AWy/cltPrmupv2WzKbiBgTHYhWawqBkt23a+q0WRbbo/+mz+u62sdtwaYDnJ7B
V/qL7u0tqNuoyY0IjISrvPCBCZ7ooJ/RofrzatuUUbJm5voHVkToUPrRj3bwwJOoDFFUaXn61iqV
n9bXdkpyC7s1bi56HYA0IdF4kqUrz4Cst4q/Hx8hzHKvIkTVG3txs0ftLNgrDznJKlFDfbbjglJs
F3rpWp30gZVLTHh6aSsfcaAXODYGRn2ViiqjZ7Z0py297AcfK7fyq521j6dOQYdtcNtVrG9Xfb7Y
EB3LXo2193Ew0rWIgfqOVERyfiwjhLRe7DSII7qVu9xiDUM+rp35KCPTG8k8BtQqbFaX72yjJJn9
A4ENEZQPtO4YYM+SI+5EXjCcujV+VCo3Xnt/IGnBXi0Pt+ld3QsmczxsIEnHw77OQkzq8uBMZ0PZ
7lm8QE6G+IaI+tF2SxLbHX4CvCpr3gjMJ5g3g8sstTUnKy1RMeDPaHgIrlLCBgXQiSYp3Kzs1png
3lZHybpbei7Wp9vIJamy+XXfo6Dp2POWGnZrklPyu94jJoy9IdDI1q2CityC4ocIFXlf0HpWT8/k
OtAjZs0V3iKQlIkJLNDgwlGwSUjNHXvcqqB5qCPMY+6R4DJNbUEEi/Ny5xfzaS8dFNbd3QhMi6WS
b4FAb3tJmez60Gi51591M5c2r3MzPcH5byeUMMsjf0wt/Xg8NpCih3E29seRevYfg2jDKtoHQU/J
mBRTzv0llUDwY64KN21zXyxbS+l9
`protect end_protected
