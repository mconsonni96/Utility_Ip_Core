`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
rNHAMRKcGCI1VrTmYvUsFXOyfJUcJ8vRhfrzWpAisIiixww7OwPe/5Y21eGi8AAfUd2F0XXUjbzO
E2jH8rY2iBPB9P4iyF/PxxqlvQoCvy8jj27dVU00BGt78v5dt12ZE2gBJ0V6kaG2D53wsA+AK7gN
jFkVLfWmQHH+vyvJK30507m647rHNCzozUixGBJCJayQvzHiVgI8y4pHUY7asEK5808LuxJyhkp9
yaF7dba/P5sdxu6mx2L1d+xeINJjJ+doszG/Bu+vTrP5kdiHujP+BF0m2eBNWsPtrnMkbqDB2KMM
I+Dhw9vKjNnZHUCBhdHBoQ/7mOGuM11RbGbcBg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="FmZtJ3iXyc+oWt3M2N8xWG36c7rQEZMa1nkwuySV7c8="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33552)
`protect data_block
NI3us8mHIajp/+cMQckJKNImiO1vMUhdTwdrUFl0nOFz9h/QcNODkd4GolnHEfzDQl8OLitnQat1
9Sp2dQL/pq4YgcB05G0IzUoXIcdEF5x1AiKePSILQHky7ykIzCe6OGMyhhMWl1Uz36V788USvw/T
SJ2weZ77tsV2e08tVzN8PnzcqQ/ZoZ/yz60RZAz14UggiUAUb4HFnRPbcH0yPwl3ewFySUvEfxrs
kvgQYLlHeJPkasE4TsLqnFQpZA18XT78SjfbjRYxf+n77CLX/LFzxm1llC2c0jjhf/lkQepgmJQo
td3KWR7XWzu5Nwmx8YoerYf9ZmTgR0rE1Yhvr0Id6jMuH8InvD2ysM68jlDRiiQUUNzVwFsvgXEB
wAIvPZxnOjFdOcWS/akzdhuzCC+Fes/NWkl5F52VJr3OleOfMRMO8M17L3SDEomK74StPTBglo01
fsUjwx1ggYXXgKV3W3SmTnYcdSYTLaeJ8bNLb58zgdjWr5fPbOUw3PVTcAH1XPnu8zvYYKkwjxtz
noZyvNx8+3ws0DItCLmo9Y6ul3tQw143QoJEjGs2eJvSQ+RJfedlSsW2Et/BC+GwKiUFrlduJT3L
bJoTXHxbAnj7baE795KMmwyPA8nH7vAF9iVpqlHE4Ewt+qxdZ5LGYVyhYmSGadgo2kWtMB/Tbvhy
kkf8JUTnkvvthlrPVc8yv7lIvBNvfQw8g9XhMuN3nXCP3v3br0lW/p0gut7vW/iXpYEKURqybocE
Z2rcFTqnYfHXSVHb/fpp06or4F3mIUypSeWHFLpYe6iO2ZR6RqQObrd6GKQ///AmDQ5Fjr42Duku
pg64kJbSeRU8UZYQTM+snGqmS42IhaQNjrRzsLuJpmtqC+LMrgR/9AnUAvG0ZzikFEOn5vKIJa+8
WnS8omegH6sQEgynuJ1u7HqLSC5/d1jaavb9FkufBi0Qsp15tisaHi7K1LDDs527SUKr1y3Wmy+L
ei27FHqfniBFSo0UFEOk6IOv3+GqgLYdQ8+3zPmcJGmZxRxzn3vq5x5HPJ4GmMFMNmNzZ1T1RgTP
ov+T/FZUwDt7gXKY9nORqGBjEMpeuJhTqXrdCMrUS1UVTyS4hzWGzz7B9+YoPRqW/zIkIpLrpDP9
bqgcdEvl8+g2rWLCm/fVv0n/TalKxjboz+HUikmdpTN5FmGwQkS0pA0/dFiyDIRSnyXYoNq1mwwO
TPDHGY1GXauXXvK+gSEG4Ps3dZsd0bO/jIwghXceikcHdDy7p4+v2eg2SBEbZWG3RJ0qsdm2/fdC
+qQAJwNgwVyznCF07O5PPJEJQ8Ag+yIbPFkDUxMTF+Zj0n/byDhk2xz2n1tgtiC554nmcgB/9Leq
e6Rmg3dh6Ontqve+aanlOc+nxoR/gzwTlE8ODA/FJtii+3suAbbTlVgux0FXUciqRLcDjDBKDFp7
fSKSEyMav5DAbSTSQPhjaOtc/oDuKFU3Br1aw66JA0FlsDok6bmQ7mhxCy74InrXikCtRNvELe1u
gHkqp+twOXozeNZP2GaHgKGj6zxtHpRQaxgNBsp4Tvf6to7r6tEIj4NkSa3eJ1k15a2XxED/Z+Fd
tFZsk5eqUIJ+OhFfhSiM8FWYbI7Pe8eLIirZBm56LPsRqaVaYF1OvH4namF+qdge/XQ/uI9NjMX2
7Clo5wUW4I7sXL1O9bvd6RUTxOnp7RWGt68d+pV38DCQnPPiqPid4IgzeeH4WfnhkAxhNLbjkUHF
60RrmouUE3Y2MTnP+ePrQ9Pu7HACMfuvOSZt+wG/QsNOcLvJM0pXmEbNZev/0PZvi7fZu0gsf5rL
5K5+F40CNEc45Jz52DOoaUuc7ftk6k1YQ7zK/Y8BGMrjRY4aSa7N/YWBSEQwcaz6rwvAZGTrHxeb
9n2wrPKJL2hCx1bnNtf38U0HoyALC8uxggVQsc/RmMpH4xBUEN2dPY9q5L/ujEefEt+CwuPYHxcU
Tut51fA9sq6TaTOKPqnamxWxWUMtVBmXaWDQLTlAvLeHGErbkopRV8Ms5m49I4ggyjdtSN0f36D/
ioeurbCTKyFQMfGqCJ4g0z9lWmpYoSgLjjpKOYb3sILACgjAV+kQDTiKljApXJ36NBUv1YJtyuIL
wnRbz2rab9QMEwbdlLRzbUVHVpDzbjTzdAC71I/0m2cW7S+SZ+XbStPBc95LR47CdHYJCKyI8nzp
+b1enXCJAkPjnqCy6RdYQgqANNUiAaMwhLztG+qv/88bD1Lb/TSiHfiPoO17ie7esFKf+cajcQVE
4eeU/2jSxYtbvakEOuo3+jkfxMqkszVR+NAx3fDqkJ8ay1zVNwlkknHxCUWNXGLRpfQg/4AUVxWe
VUPo2s/I6ZSYpdQx9xaOICs6Gfn9f3pS+pXNes7HzpBe5Z9qOPjguLwYA+KngidfZrR2XftXbsyj
IZeczO8Bl17keNXXe899I+NQqLdFbIbbsP7YerNhlvIpcvGIj02g2dhx9u4hAiJwVnL3KVdgHcLo
wAJ9xdWi5wlaejqy91QNK4y+Ioym3dvVjR9kpCifV86O0MqYCvm0/GddwblIrIv5+J5e6DayCIDM
TKDgxKgth0g+MRgG1RcLo0NbcGWv5jrr+wZc2DHourdnoztNH11Le63d8gp5tftEKnDPXQoTL1o2
687FMIBhnpuGEz+qM/b/q/ThZNmIL+5gz6lBzp17F8S/LcMEI1t/RlaD2rQtai+0oTfLuS2k4f9x
8gLYIAddtUfoLBdrBRweDOzAsdQfRDJ+GF8IjzZQuf5CZsxNFcYivLwQVkwl+BO99eVV6fC5MTuG
PBGlYEXOCaswAYbrUu7IR8TJKmxtk6JIxBYa75JzkjNMUVoJUOFmEbokFQ6yPQMliEqFxp7GK/Fa
6b8wWmFvdc5GrakQeiBZU0z5Ydu9clKYXjAsAVQCgl4CRJBzF7uZv+43g1fdaYOttkiXn7faFLjD
53q+lSraFIrnWw55/z9j4fPiygQ8OuexwlMIYXbq7EOYc0c8JckohTjRX5rBuRSlm00V5CVilj67
nwJHRaGDlaXnONlQJRUSbuomqsssn2hcF7JEtS/NxzceJ5mbuDypYbedJfoKr4mVNsTGiBrwo0KY
Tmw3SFqfRrs+WM6qmPhA5Qb138i3Aizj/7W6IfuuAodPdfnDrjGLnb2Y2n9oehrypzo63q4vol+u
rcbMYP8KtxL4M+3J9nZQM6+ybZLOzrNbdeNIYu6HEu58e9RnDKwEPhJ8hIizlnmHHxiuk2qpuIgX
DYhP3DH5tTwJZXV9UTc621+LZ1BISL3RLyyfQ4iQ6tvgeHAZi3kO5sxLdWvftmeww4S2CXsRRhQB
SzfMvZbH3EGVYSORw0Y+1XLu6nDrvI0cBvAWrrFYtzEWRNF/igy5FPgBLP/PaToWEYDPnfeACkZp
J9Vg49o2xKp4f3temp/WNAa/5EAWSNCzrED5tF77PGIZcvAKaGqbU0KkeSgJjgo54V/4x/nnnvUt
692odGz/AJqRWqQ2nce0AkqVUA14NrKXOQb9Dc0iATbYUrmJSsK6DqEGbddHTstpuf6t0+67axbH
nK0G1+JbaJmlckM7jiALK3lcEBb7+tzQFp52Gj0qALE/SEdvZlTZPChY1TLjDAhVgyulmExoEpX+
X5TqmrwGAE1vAqaCH/U9YjuXPMMv4qoDRWbtJ36MrJTXurQezSthsMwcnSm/qwlen8mS9W0pFrOY
e15BDgwebTfSvuh+y0Flkg1WyZixJrbIzh8mP2XXexNDHwT5Zgddvt/0w69cnQ+KyjhxTeKWCd4b
uPVQVpCOCrhmsXrEwt7CifDZ/DPm/hYSX+1lDW1/o6T1PkrTY3NTc9hm0vjTvOhR/yQa++JoEScH
iE/Yn7KdFxcXfPDVu2Zc0NXNVAoS8t8wSEiZYR5SQl/mlgAmQj2vyX2kaVcvg63qHh8j9ivIcE1s
I3EZ9IExQbY9A1jqyqK0xp3Is/im3LU22nxs4Aj2QR8JpPpRR2pPDbQYtiUO7MvPI4jcDmhHmIj2
Bu3Gn/tmghPTq8sL9b9K6UuzUyUYLL4rhOvV2O/vMRqoiGB4ExzKdI5WjFWldo1o7h2Me9EFN8be
AeoYisn7bIXdQC9ZYqTwDmfQtR98nsqMNTRTd02Eq54v8MWFH6YGBIFTE6kqmHFUJEtMkNuxm93s
UB7R839hPOg0MMFL+2jjng+CdOfNe4KQ/wOO8s26AiMzCTsGdFebk2EUVf6GBWeazAhFbxOGSq+L
FEpOH6iCX0F929vtsMX4jB8V/uKkDq2WpSgdXp5y7ABmndAQqRCw7jVnGd2dj2F6amTqLFLSR736
Ym6vhcCzGML1lArlYOXrO9GAc1zq2q5GLkJACGcwuUVF1Xb56d7eSpqT+8RNKv/cUXVObl0YR1o4
oF1uMrsD7dW4N6TxUESVDJD6yviiGmFzhGlTT8dWTyIkFDPoXR9uAJ1+BF+oUSz+SOG8urUKn51b
SEaaQzOm8IJHRze/vzNaJVyZf8itTD9rhlqLrLsPo46YssRMWgi9eFdgt0MxpW+dW14ZpFNqb2Yb
2Z1fA7vascGrePYfrcicQyuoh9PFJ4nPH2/1XxcAEV9SfBfxp68BCWpVpsePWtw4MzYnI9Bg1utF
DwCUYcqcw64O+eXhY/g0cq70H6VTN3l0PZc98SKFkZJAJ2E0POwnjP5J4DFfNwBncnKLXTNVyQDk
7siWmLm0phnO8lfQYi915MuG6WuL18AGrmxH0qPwDBrV6J+x50nzrH5BdfZ0I+JRllCV+LGr6twl
Eo91fARiK89WQQaUhB3GicbNqULkQY0pw3CwUUFkPfgmTcjKZMkW0jqWnIualfS2S7bgjbvPJxha
Mo6BwaxiOjwfLA11I14PlvKKDdWw9PjdbZy16RJZjAt+dUvjc1E8hc3sUD278VErdFxJp6vvRo5L
iKSLplF0ZmzSz5FVy05rEXAOQOA/E4TnkR0Nl1Pzh3RSQnS9Hs584qEPFlXCB7E4itMeFtfR/cVH
xbcFdfMMHpoFiDXQnokhU89GcwB7b9K2gvlERZ6eSpuwE3veZq1NOyPhnTBBlqdS9VMt8K2onq+I
zusU4AVpdQg7gV1x+hmjuLGtXK5JpNIT8od9Km6D9aATKKQhD74W1Y2P+7JLBkIQkPqa12IkysV3
iDpUIIh6WIuw7Lc3FZihbYFObQmXg4ERyCa05gR2xJvYnG5uKXs3VCcn099OkETj1ImyzoUJsv55
UV1hxy8EBD3BuHIFoepA7sCpNMYlwiUNaV3TBC+16vdszK/V4u6ZNuJZZ/SZtKHX4zV+sYn7LqQK
ZO0rlG8T2GuUig5g+qXAZLA2021A/IJR7GAdmG01NU883d8N5+JNjS9belsxXf0RejIr1Acgc0lJ
F7v9zGqvZcHoJMzs3rUTja6TLi/kzn+jPav3kzH+wx8+s8WfRV6tibgCwss/h1bszinLBY1SDgb+
bvVsycU4+3/GWQqt8x6PM8VI6ysqWopKIUkoMxN5+4Bw8yyc0Cu1kvGUK9kHnVLKzmL/hY77myK6
x5mK3A0j0ZhOfr37PwUlUb+xGVuzCuOB3M4LIIVmHN8HRN87WPlbjFpa1C32JyeN747Z1OJnXbyj
eld6p52rOu78AnByIwHeTqmrwcj56xN9deR07nNwLuwNPO5OF8JCBL3TsvWDVaZMoIKw9YV4eTNo
M0bCUXvmtkKpOGL61uVMfGe7iOHc9kQsOadx+rzP5c8jDr7t/XYiAOlLoclzzqkSY9mG27nmI6jX
GjyECO642OrBHejtv1gX8hEjcN4mxEgC3B1oMND8Wp4wqm6/9ntErwSjakZacOXhZcQv9XDPYogz
fWjbNGqFOe4AOIjPTl+QD/jnS8YVltyrLL1NvfjsaOnKhte23PWKor8Xo/PG/CWOcT46EhG4R4A9
r+sGxDvvLSwr+Fbr73+U5s9WPG7OCVRypHhwov6l9Yhjn9jkdgV93M8m8EienKITxFNKZZV4//oE
+Ig2LkTB7DgT+t9ioceNsSOPFq0F/jRO9fzx7LnHHDhrXKC18NNKlJQ72Agi+qFp/iy5YZY8HT8W
aNQ9HSY2l8NJva2xgdYaUbcUYHRZIOZ2SA+8DI2t/vd1q8FfdxD5NggQ0s4ogmZDLj2EXH9rvwqi
Y7OjzxyGk4Io8vM3sof2BclpXfpnxuo5SKmFexATPvyh7dgSKr+EkCHM2yrlWRDPwuaDBMspYHz/
0PBOiXpdNBcwiqGZ+9I9l1w90OjFjQPlRSOvBKjnW6OHKmwimYm3QACdzUPQ8n9PLeKyni2CX5Xn
g3PW6/2zl14h07dAYvI9q/gdz/vUzFgUlYOL+L3DJVciwLe0MY1Yhr2NMzVwFZU0fd5wmXnTm3lr
f93LwlOyLjg8dOtTsAiy50knkNYA1Th8MNkOL6Sp+FEPHhRrLE6Ts985c2EPQkC4Ralj2cgJ5mFz
yP24SMLOCIBxPUqbP5BMlpg1KfOeJ52j2o8uxH9f7C0txv/bpbyZ4XHaYrm4tNj5i1MrDa9CsH/x
uv4Lv5xMyiqSawByZAnHofvuWgWL/fBo201ktiVQnHr5lHSLuC5GFkbPs6tzWP7qEeUELkXqYx8q
70lG2+GiS0SkzTEN5lB26en5DwT7dpWgMjIHcGtO4Yh+TMqAvESz1QCGK2Sg7cigIeTdg18tuQ4m
swN9wgVfEn3at0vbxOteDmix5ghEhMiJWNGLxM9i4rcb2FQCuuxaxkXFVG7abDcD7ncAI7igW/Vy
26lAXKPpQ7IVNOdBAq69HX5Dml8H5ME4cADvsrSSTVtdTIRbCU4IWLWkpk1hdAsQG5YWwTWIqTkU
jaltqrDG5ZAw349Vn/E8LDbZF92dlteuLAFLE/QjAGCnCH1lCS8g3QJh3IEzXnpWqn0zzlcQNfNI
zhxtcXlEedj0Y2aQR2qi6Uy4WQsgFzenz8Vf771LjHN1OUOyQgOliVFK08WFq8nbxlfEtnBVJUPZ
hF+r60bn40ZIU49IEeQzH8bVf3+rHT5dWY4CQAtq6xzowfxJ9DuU/sRg5Vi+kwmhtaIHROJHpBjK
YfzmJWJ/pknZka9eUzLCmFii0Bo0oZHCMsY6HOTjNCjoSM0rCdwGyZ04vJwm72C2j/Objnl3CgRg
oDe0vjHP50wZhVXV+bVqtTh3aQs2Hw6jS9F1muLPZG5HXNhsAc0spDrpZbFFXnbLEdUPzyGGGQdS
wLD+Z4n5alQQ75gAa/ge6y1ApK0zUB2hbCeyWoxkPIgnXpfI19U7ZqpsccEpDzyLZvMheRgKAVbL
Mb0hhBagfX7xkK2goIUhedSLozwt0HObr0rdr/2caUY5kY5Fd79udPCo/HJ4tkQdy/Y0yWjoiFi7
FJrNLGBemwzfRWYxd8Gd3+Zvax9FY3t30UkcDMHjcnxqVfrcjozfCHQPzdlEfY8yzHbSfJ9o+FGD
SaUv/oTDPRSL6oNb/Hq+Us55AJgYBqZZM3zLeLsRfOCfbsKzk8R86t5xwQbxQ0ZcYOr1SQE9NKtb
ToRcG4ptEJkBD0WiHuNs+bjHSOufcJ393HW7jzqFBLVCjbTaBJ713Kj7uVEirgHxYnsv21rDgBng
1cxCJBNwHrOaswHtITqjwzmaNgs8o/SEoHB4NLNh3TfTnUkW2c3xP8XZzzefQEScrCRwl6ddg0e+
0u+yiohYMFPrODE0D2PHlCRSMTaAtWt1plmh+COWO/Lr8Ne62rL4xarmLc18Pb2sogrQmFjXwwe+
qgYykJbIEy259vDdcg9P7645JTdiqNGG4ntEENVRg2CGtSV7LLc2+7chZFRLsgzlIke5+/pKKU9S
6RCxOYfy22jw4SLYdRFysjJz2A9bvnyhkTkXi5EPAdwjLff6s1oboo3hsJBf/MfanbDhXq9TaFQ3
vtzHmsx1Ee0qt8CHrYUbssIvH5dUsPMMpSbSzcmTK9k8R6HGm2pMstKmnIapftpeWnKm9MOl6588
7SHA8O1pjtehAWwvQIKybZFpUgs3sOWyWGv/XHEfIdLHOM2F0BcYdEHPFxQ692/iTd3Sf3gyG2VD
cvp9bxybxBFgu7cr/XJd05xkPPjfPG11UswOMfoIcv7Fqfsf1hkkT5IPMsBjDMZVHa/uh7T2lulj
l9bNRmmZdL7HL+sa622bumibKbIPSYMpq3d8xmriTwxlBnSF0R7Dh7tdxWX4utDCnl5gBQmApCaf
Y9xkvqSO02o2TMZvDep3pFozG0kuT4mnEOlBjzDAmdL4nuW1MSjmO6StXTSbUtW6w4sG46de9ae2
VsUKOcBmQHdwOoqFpUbypjmxK7+EjQmTqAsxFnO1l+S5+QikmpH878flbiueFRU5S7BMSFCNgVYM
oRTVpifzPyM8dC+Rz1pOtZzUHEQltmUTS4skkmVSQJspYTcCyCK8L1OT6ffOlfl3JHOwzG+R6cAh
0GB4AInOELONnx5Gq7RJ+Jx9cM2djM1XS5d5YphKVgxS4sZqfek42BCt4jEVyrAH06p5qfflipWh
NvN0eOWbO/IatmFBR4eAyRmpJz7eFPjgbcjfeuC4wCjMaQt63nXiblLikzbSlkaNWlI0UeSP9B8l
LLvPLAWxZCm90qvDz25hktktictbmMXwPfyRUsaSzRY1M9dLaiqux0E0qsyC25vwsAyCUtrLoCca
QLZIgfxVUKTsj0TKNzTe9ZqOWK4AEsZkNJZieQQBQgD55PcQ0Cr6FE9tj5bdM9HKngF+jDCU+6+h
GTLKjNhmyp/xj72l5Xr9HD4o5pi1L+8d2wSoSZ1EhVOiTO7aG8p2smXxDR5mP0fxT71LfDQZOJf5
AaQLruXu1ze9EE1BgrcM9W6GfL5r6NHj19KGNeiXfWyM+tMjAP0a/1qvo2z9qDaVrvXIMqfzMyoQ
1IgAw+0HGN2voR9xF/Xbqv2tkrYO83ZXbNOO22L1SVFmEKRNoKkACF3K4DGSXvBRc0IzvN2wG9ip
fSMzClgrb/eGjPfFkmEcaztGq/ycYzs0NscDP5pRfWcyhacl1p1ckCXczSAjfhff30GnNjCEldwb
lj1fgEDOq/TEu+IBUJe07Lo7Ha4XbdkeSJs/4D1zBRhOr8Tc4p7SvrlIKMwB4cvJqInAyAadYqET
GaY12wOWf/H1vp7/JcxMzMr+UyOYvk5KEh8PjBAQYNXv3tfilTH/KZr1rfyR5nWaLMsQimVx5Gxi
1jYhf3siHm2SXQREt4wIJ62CM0pooZ0SbXO4EBpcXfnK/W3A6sluTFDW+Cq6+yJE2gp3BiKHzyNW
4lFwlPlKuErsTAKXutEKRU38OTOAbCVCcse5BvwZATU6zon3RhyxA5Dr/eTys4otg7XNVs3IT7dp
EGfI92MbtrB1JPgb+ZnONV5RVQ2j87gOxm2Z+euOFOuKZV2OpVUVkWH7VYCwrxpvsbayYJKTZjVq
P381b2snGTgjVxim42K8N7b7vRtCisdLZwB4f65wWh1bOU/bAtt++uMt5FjuNVcsZaxGJLZo5XMI
QsMCE2niDLIY0eSe8sPP5EI+iZCeOCicMPPpz668g5W/fj5/OZ/Dl1/PFRNmiNPZVnYcFNGsVYj7
7wj/mF542zzNQ8DDH9WqdySxbVEnUMLN01JvhQx3CW18BVVmeyoU0Rqq+3gcGO1yw0QOHBAU+VPx
GxijdbVnPUvpvFeIXG6B/wSO3fHv0l5js/VdJhirNxxMOubOWHcEb5Vhhh6tOUn7umd0GTd+0z7Y
x4OgKMOHF1wf0sr0XVbIIn4sIdlFzWs6oahnuEXFQAlHhYcIqEPjxUm7d5xH46O48S9LjgkrHgiz
wY+Ck/DTFWfHS3AoyAzPpZ7wDf4pnXRSuiB0nh/itbBuQ4TX959mMVEHBbNUPDkq76xX+JDOO0R1
zEVcSByshqhT/A3CH99dsZs8QUcrFf4wbvOMaZvLTR774fk0ltVA8/WXIuVYWZf9/43+wbQ9gpwH
deCg0O7s54fUtAltiL2UxQjslmfG1jEWtsRmfVVe1P7XP11wKUxExqN8GcBSvEqAFouhA3HiGEqn
Ts2oFO+YG0IkP9ybIq8LwK4/ag/GYG53KyQaDrnPPEC7C5qk2BWWQ141A8l8LC5gHcJIXkd1CtVg
OnXbuJGcZ1/pH9CfppHknH8adI7R1DjVt6bFOWPnwXLMlQbUjSZ/5+9WGIo5GvI/Z5vp4ecbMSWq
yjPeJaAFzxWgIjCC0AXrPmZ/a9uHT9O8rbZFo06N7LIpLTXOBfx1bdeG9QTVcYK0VbduNnVYmkYH
zFj4MLD/CSJOJjyR6xmGW33CHdWAHMsR3mmWc6RqPsuBsaXj6c1ATLuSTM/LfoaHyD417snECM5w
C0Tdz2SQdbRNwMqiazDoQg1CHs0vscpXcjbz5GYoaOEDyyiJfZawmbD88xjMp1LDDYEAND+5zeri
RA2IPg9E0cz3mhI1RzpIS1jKhNUsp+pVmtc7Wz7J+CJ77MxuM2BaR7QT9ttSSO6kcycsu51D9v/w
M7bOD6agCn9UrPyKXWUm2z1MHXTZiBekzPbQT94X6DsydRPl/dRZJttmta98QBPgz9rQe6qGdH8b
KBX5GBaVA5ragbHBSA+6e6z2VDmeZSRY0CHVmbQi4tt//S7hYyPFsP7T2+bzcQTIclAS9Bmox+CT
YtxKe872nnhgGUxMxTRGl3LMu6r+oKJY8vCit6sEArtpuBuNmsJpm7LziCA9FDA0t5lcDNjXTpU+
GMb/MzpMbLzwkJTYWMFxah2zU7n+sqrq+xNiLyAFNtr5bSEhTymhuAxPpPikU1zQkqp7BnNL40T2
SnmVRqnitmrcnmxcjAfoxGLYCDZKhn8C09QIjbckYAOspCFmBAbO3s6A5Rzg/LCX4hI4pJK6dKtR
iW/WOxa2NxV580EEBTjHOR9qfkFieILqma5a16SX6/LQsDNWtT9k52HLwYWIYWqqKNiMdxvANlMQ
OUBslaS+v+vCJlnO6L/MANu1S9jrVomdpAC3Hm/CU6TlYqxhrnSZDi+O1YFLUQJNazcTJ99peC5B
r7F4GjlRAi99Jvgi++YSCY27AAoa0LSZwIuruoGwiavWN21z2z87gwb5Y/w7NwYHrsx/hUsd7dS3
98cs7+PmIYER5ejkJa/v4jsTUCwE45MKbPr9dvZ7261R8Yjswnl45HgeTqAg8NhFgW+ZtMAWM6AJ
/tePpFPxqlSpWEiKtiBK/FqkqmfAsMDBLC6e2hvObKpWi99oPCYA5vAmMoNsNrqKFk/qs+9V9HNW
d4ISDgliAgG0VsK5kwq1XojN/+CPAmYTue1+HuuaUk+bwvRRgQiU6FK+jgHTiaEvbuJB9XEX/KDm
clHhR8+En14RTne130ZuJ8e56gikGxlgkCMMZCy2lIGQ8PBTDBtrTKVbvJ//cX8mcCZlBR2MIhj9
plnJbCTH4RuC92ryK2g6fmRN404gfMz44t8srzlKreTLYMR9TYGSmZJvFuFbCvME3sSgQiP5ulB3
FYRC/8iOvvyn46zJh07Yg/W2xI77KoOiJobW/y8Fvl5T4nnLB7M7woI6BHS0o2B1eTkK62kfFLyR
XmW1Ao0LuIKkhTzyBK/cuQqTZ5JHcrfvI5hW+u9JkWnPvXRUo6dqa1t7a014VywsJ9rt9JxyDpuO
Zt13GH39+tFpodpN5BOPfSKa/V4fR26qtfg4Dpg27l41qYbKVIunL7rB79zCBIpRT6aNWhz+vNcx
aBjhIsyzxLsSEQm41dPk4kcUi+3uztMOs8h7wrzzKfQlH85fyjXOW3fEGKoB2y3WuXDf4CzA3rQB
y24nM2TWJmLUqbPkxBymqFCqXKTgZ7cT0buocZo3XSRJBTHElZ204mw+thqPfKMwtNt8kr7fDl1Z
YSQzqk2UJ1BcOkZZPGNn60+OJ4tW9jdMvgmjNWbn00Pt57brCrg6P9rUyH1YKsWlVSlL+SgX2fwu
1YgKxEJhlLlIoFikjNxoCMsxVTO4OZ5mJyyRwn/iGkvEGJ0Xn7muVG7kg+sbbx5VW68b4SvqALXg
Dzho5qsD6cWzXP6x3vQQej8++c9ujyGvFBoOw4iF9yzSBZ0HBk8YguVF01pJVHv2lLwZKBq8EkCn
J5VNQhGDkRe51cQuz7arh50n7DcWiAoRiAoty66Jel/tkRr2tRpo6CviMYLM2S+o3IYGz84dQFez
g8fXvLZQIjtNkJeX8tB7Wxry38fk4qdnNqRLw7aPTGP4W6HC/eIn8k1SVHYDhoo4shUZRlfZjMYK
qiqMZbVb7Wot8tttH6kF3aT/HbvHZmnKWHCh0b4WiD/lNukyp3CJBk6qUVNmX9yulkOymG5y8yPu
9GICuS6gyTx+Bi/t2dvyFibRUJFWUMCeNZJHXQc2/nNiuNVOvAaWCBnXPvys8OjDNg8iEP3Az/HG
gZdKxTgBOTs3kZp4dU4DZ8YV0cM8eEflsVeCKplEFWeJRDprUHmDZqJjEgUcafZjgCZTdRj8dXTi
27BxtySGyTRgzHJ+ouiGZdDWS5GSrYsMvvNPXoRifAVc8e4PbNbUjYEY4DbzjBR/lhYAfCxy5+x5
L1wUkN6tQnDTovXxQYtFWfkZt4ZLkQm+bQ22Cxp/UgJKIGJhjXAZqBdazYmHH4mOEienq3l0+w/R
FPpOeEDhkl4s0numlT3VFiU3SQij07BkLUlk9apGb8Kf2dHNX1JXokfBufzN4cX7fPKbgvBs6BcV
XRLLE0fTFUoXcYurF7nS8/RclCdwePL3ztxnf4eLXmJWXFQhGqlGACN9AFhd112x9RyX+s+bIxrD
VoJ7YukMXOTGrYZDTYVUfyDi6TRlNNdVIg4q9Q8paZxuEraD1YJlM7hxLTSKlft4iWnxD2OnZVMQ
U5EP92vHzV9l1wa08DpmEQSS1y1u8NzKKgL7PspQyjNTgj2eWOCD6U3D5TNMGtoAsH0jHJqFIrND
3ZgIEtuPMGtXJiYqPTCRsOxBZ3pIn8Ori0iVoc/Li6YkSBzGPERR7MWvoc+X52ZhOjTtaFk1tLUT
AuxRlKo+MHF7nfO5xChcDZ6obrTnTSO7rYQqp1dyuwLDgHOFllvHoEmZGBqx0xnwhnJqyUJdZelS
0+wKtpdNyMP6KFPSHZypP4HXhD9GjdcXKHquxw8wgzhg+1tqSMboBsIc1as9BJ3CnvRgpujG1sE1
HBNyA6xz9/n0bOvMXOj1gDjTeoIZZ2M71BCvpyrjxlkkTDcDhrQxJy5RDd1NPO9uMv2qLolqW/Ef
fkduP2pmJiwKJfWMQbgm4Aazq7hRpEdCSiTTjFt3ihUg7FTxCTVPaej1p+d/H7is2KHliQaOCu0l
1WdyLmsJBsE7DbEeUjunKXqVoCAfBff/lyMuRj+LnAKc1QzMhaxWq57REDdLWJKEemEGWLL0bn9y
m8AD9PKpGeOANOAVgOT4jvMhG+jrWcCze8VyZQi9VnpUjM7kb3LURbIZ+6t+B1n2wx5uQgZykXfo
r5tWNmIzIWHN6KKHG7wHXEaXYnDlPZKii75ldM2cnm/xk0AJUf5kUxnxVJ+5H2UdK3JGwbRULlxX
v93RrwxAZKaihxJMu0l7wToc/CRxgZUKOQuhlGD2EbvPVAXqZlm+2hdkbN1TsjdWvq4j6rqztzWY
z4LLwWkFAVBg4cnd5xm9MoW82XgFlKWCgbIW4HWhjq+UjetjzQ3OQEvxyRYR0eWcbeRDFML/yAAw
6VmvICMxO7hNGK3PTwwdnr0KP7VCr9kFeGU4q+lHJEARZnzpjK8UAatP+5SJEDzaVYQzggedjctz
ytYjbUKYId93CBq7VXscEthFaMdKXe7jXHZPlGRdaPs1h42AIPzDxTn3Jr+vuMh+QY+/SWnq8jVb
1/vWWksXp3/dehh/EjL+lfW4/CYQaha7U0aAdwNP6HS6oXpL1LfXz4uXQDtuRp0FAHszRl+tKwEP
jFt8txc++lD4RFvfa7VOlRmmNHvXsL+WwMz35mcfOuUDYDfEPKWpphpUpufnTZteTVPFqiKJUFQ7
GGr60jzKJNVAMOiOQYgq2eY6+aY4iY/ZzaPxGOQR2PXGdBChPaB3VUje9UAPoQCxV7DCAKznfUPu
EawZvQWidEYunzlN6Bs8jLEw7EeaIScBlbdCqA8LNlJ1BhZkLaA1P/8pkTwX+rh9XuE+YREhhlw5
akNHnT8jtpOWODSvE7fg/gqiV9k1PceQiwcLoEIC+nzcLORkGTSiane15gF0LAKIyNWQLl/PD1Ux
CHiEuJJat8OXMoWPx8/100oTHFVaIFG84zsFcp7nfzdu6MhyocZNuVklaVM4QBnqTHZglQYnd10u
QIYJIHWUeEf/02PlwHgmtTbXmLfaBq5Nt3RLq1BChln5mxSG8vUj75M3gE7y98Ey8AZzV3jbgEsZ
t8lX6JfHLvNXbUAxeCvbukR9NpNKxnUkkJqarpP7Xp2vEsh67VE8KLXrvnw7/B/YdcihhGUxLwW0
8d9kaBXu/o7vi541wUSP2ndW8sMVpFrkt+0VjWt+izXrZk6Y09VqyNYy5HbXvsiU12wDYo2F7824
G69SZb1dRPkuvgxsqabI5wbcwl3zMy6v6u7pQXElUghhYx+z046HwWADvg556i4kK82Zpk6y8K7N
/KdWvL9tgkTDQr/JD6Yyv6vyPdpbz0uVIdqLa23hz52xYkwSx1fHVevxzRCVy86+njO8pDqXgDQh
a6MAikgZwiqZeMTSXGuHUYrKXB+8Q4DJ1PEZn034qtVC778hnVr2iVsDMIQ2Nk3Sm825J0f8LJ7f
Oc9OTia/D7nz/wKKSZ//A4OWbYr58LLjVjn2PYX4LNRXHyKl7SCPaTI1R8Do0IzovLlPLSI8RMqe
U3h1mFEQn5N/TO3o4Tuq4WNC3ZeyxPqua5jkfcpv0wkC4bUEqws2npHMh1ceIa9zZdSa13ELfHa+
BnzNz2MDeqhsA7vgyjeWaI0bae/j7+tU5pjfg4BHCeQM1/PfefPpSVvW2FK4pQdwI3r7XNzNs+Gu
Uidbuv6QfGBAE0C1BdCu+RRLgGBV+ERVDTnDA5MIjRT2aogqjoj7DBblGWbCruTOYHCljuqoUpp5
nPqiAsm2V5jl4zxYW1iMmAqOkE3tbYX1WjuElATUcZBsVwZFC/He/TGjwqFJJWDKMF3SGNheGsHZ
XO5vq2LfCPP7It/BZf34HrxG0XmaTjTgSsr6+BYq7cbC3ggfPl5dwlcX0WtVQGhNsARB02kdMLpP
HPNm8thmaWpOFEqZFbtEdX818XuRwhJeQ/3DSv5tkaLJFdIL+7v0Msi9xVoPhVHBzDxr/8F1SJ+/
h3xmhILdGGPBMB21Wcx4GOxUoMiepwxSxZk93Dnq9ntbdESd08FOyPzQ7bk46h9SRM/i8eI9V3OK
B7mIZqN2a25+VsgzqeLOvcYBcqYfinYwieVwzSnIjmRt+5VbOTLIzgcR0rRQOEZ2wZZkr//eKJTe
IqN5ITafKFehtTWllY55Otf6F3vBGGmtjKdoco3Oi6wSG1KaYXiVGL71mxSQd7XiNJnuBGBApj17
pvAjev3SuDCKOzX/tB9w1KEajgqA1vXkMIN+rF26g2UO5/wUWovw0lnsKI0sDpY/sQXFDbMeL8l2
8OTuGWA334J/ttrAicLscFcs9cUGDtuChZM243d9wSkVLgu6/rE7PFHWt1dpw2XORWJMA8tFIIOR
y1pCuCpU8kEFGYulROiETEr5Drer1JRYHXFo376wTKmFDzytmpBdHoacDqRZMLr9XK7ks1qN1l5+
NoavHjzzIjCxYamzVtvxc9ZXyQNrmaocywkBVvOD+/LgE0eKGgsAaVBr0loEn0EBkS4VC+Nju///
S6SUcDEeFd86L2GYAT+I8xysVlsj5h4SiY7uh3dCxOgpft8S/5do+ZK3Z3TF6e6RqG6SjDoVvLey
4KaB2acE5z1TRx75ZMGUqVGobtGa5KVsJmwSQoLWAceDAnG99Z/FzD113Xiyx7GTwkbOILvl9ZSj
xjgHqirX1d0zt3vNSPk8dBpJi1ZGCOz5nkTlU2rlJOeyfjNlI3ov6H9wpJMCCbakypW0/if5z2ii
zMQWDbmNFpM/1+bB7I6miApvfUBkKE7isf0zRKlKuUiSHDg5jGeUQHmT5vRjJqeCN31O4t6CLojK
rMzob3Z0p5w/3dJSdFoiRrnooeaSqBWCDuIbc07uXePx6IttJGbinadu1s0HTTkIqleVBlbmtbFO
Txs9IDwoc8fOaS2HBDmt4nqa/NOzzkZLWkYy+MvQBE1MmHUW9okAWqe7vroPBjQsXsuKPJ1GLRHp
Ic6OSraGDZ7X452lIRargCrJuuwCAaIWKoSMv9e9rk9W0ryuMtiK76eFR/5C1zULr6zlVTg750Gi
28uaHRUksSU9Kmdg7IR1bzHGDUCAnHTuECHfK38h1fOVUw/QVuTWzSDy9790kD8BtxGoK/aTSHbO
kZki+W4NbS5DV6o0I2xSI/9YXmTx3UTAkOnG/v4uePXUVhVqeNlPzXLXOlUCtz/6LBbmv3Hv5Uf4
1vuNmWXSUoOzKB7dRgT0jKvGjWjZfelYM3DEdHzZe6r6lPd/0V2c0HxO46yhFgWV3SLLcwIaknRa
JNUw0xbW7r7iVtN6IguzqVRSsDbTvsItmC10Y+40UYJ54bR0HOaodoHVw4ZstMx9cNdkzr7Sn6/h
HpckC6OvWurbgASF3Pbn1o+RCFoDyJa0b6Vekwpp9V9v7kv3AVFUvpcANViGKbBb1JavJxoN1kl0
Y6Vp5lytB2gMfWxJvcHcxARlkDgAUZwuFcRVsEjJsxHy5RV1SLp85H40GdLML/jSr5EmuBVRbXB2
ReiM0Y3R+387v89+B6o569qkLwtPM8qx/5KFqXRu83eDhYCE+olyqB0btpzZiSDziF/OLO0ENu2q
L5s1SXJJMpkWrRrbV+eOUSv+VgrNdUtLUZtWXFNcf9rikOw9CH06004USfvy5CQVyNORdXcorckP
XQ/95NnPuoehpbQgzhI0aCVepYp9/Bmzb5D0ws4qRVhMvNERMXjuX1EAiQ+ibA21DGaKsmW+0WR1
f8QzXQ3SNYNAHMsWDI2CXHdNQ0QX/uFVYL/hbWy7gw3X98LWuROsP5RKP1EiukUtiY2E5nHjhD9f
shMGMriv8BSf0LNBVUcnqaR4xedYz8j31t32dev1qYdHhjtuxBcpc3yDqKo7jkZ2LQ9RQlAkz62m
GLFs/iw8RgCIi/dF+hy8M29ZaAN8VxxoWUWBDFgtkKN1f8d6kJVQdszOkeMAq+mvBx0EvnvM3oP3
p4We/DkkhiuP4YtgUyyHeJaCRntxe+6kgZHAFDiR38H52xr+i/ag+o7s32KYq48xW02EKf7OguKG
N2Xg9MEGSWeAS5NvuLGeFXbHejuPdDizBDN3aajGLdXSe2E1lCY2C2OWpyIjKDRN8PuaSAca5Df3
nqI+5jTPJNNzjiPM8pW2dnGqqKPvbZ4f2scypK2f5OBhpgC7U9i939CxOt+A8fl56BAE91J20+1k
7MVCb77V5QC9l0HXFSXx6hb2lDO+2GhS658QU/QsmaonfGFmnrPoJpDg0qrYQX1bG0tvlLEIbknk
mIBdh4VVPDUYtC+ZITkWYK9TRe/b2H6OBjQvpstoQmrx9ZL6FGfgcsS/qkIZ7W26aavPVVk3Io0L
rBz2bfbX83cW2ofYoJUShl7G6qbNzVo+pU+v3biRP3pw8/Koodoi29DuPWpxAVUJFsmLrer3SqiN
oH3wibv7IPVbmo6YMOKHOTCuhWi+LUvVmbqhNAkehUFi8HzFQr71AIRxS5r3alJJ31SIygfKT9qH
Zciu2bxjvgPAs9WEOlPYk29l6/3iUTQOim+GRnAFq+zZGlL8/DHZMsndqMA6iQrLuRwK+cKN5iFw
5pjwoPHuBulRh5WfO3p8jkkPZZblERW7qiJNG5Vz8Cz71r2X/qKDuHnKH594Gv+Hvd4Aqk2UorUb
Kq9cEsykBbIWCPefgTR/KXRGJv8EpU01QUuydw9QXbGpkaG78YyIJ9aJW0W5O3rfsJZipRV8pQkW
lGBetPiMHagbO+wDzf0PPjsA2fO8x2z/SF0kvaAVwuQdTB34E6aegm88MT0NTYyaYJILRkzdvMIA
wFtxUiD+3824QDZyP/qlWEhlUCNhoc/g+lv01m1ugUjwaoZ1JXiliGAtYADQxS7lMOsD4dYSv4Ud
ZkSt6EiST4wDQQeoGMFEvgnlJgmmrw8Px4pP0DWf1kDt9zcx1SnFIqfRDcG7QZVrRHQZZ6zC4WM0
4p86o6tH2BWPefc5sephjGA7qj2i9uw6NkdxpsUVZiTWsUcbIZ2LQaUovNy9Fu6tYbK3qJsSaPzA
ojZ4kRv36b3gRpGVg2IMDHy5jc9k7s1h0nJkpIj/BnRGZh912ufL2V9G3Gie8GLWNbnlVS/VsA4R
9eIyoVyAZdUFWfqMz1zV9vjh6e+kcFkCGfNnNubeWbv5RlZ9APdcQQfoylXVLOZXaiQUs3u2IUBs
fXQ2RaWkCZnvagly/UM2WUqnShD5EquU+7AHxKuNq/wFrnIvttZ30x7R+zztHPaNhpqKWJNXNuyj
gJiFiuyvItkA9q3a6reO5CuRwGFLDqApxcRrVwNp84QAsDhc99uneMp0UTUcv7e5v2PfmLo11lR5
8JagVWSfAMjQ3MGz7BIBjd2vfdV6dqIyYL7O0eU0fRBEcI0NYcPRcKRYw9yCflqUK/qpIADlYNST
TizMdRujZSPlK6SSiRQMbCQceD/ZAMqwtPIWBT5BzzUqPm4W7x0HLeQx/LoFTG+fceG2Dgv0pwhP
mYSR3m/dEyb5sUya6Ln5bhpSzNaATsU+b7Sa2wYjkkVN5CiL5iO8iOK/Jk4boO4DgJsXAEYjeoGd
81EXOl8o2/bHqEUcVJfnBFdqg/GnjILwc4TNFdKHOzSNw2OFY9V8EDExHgXXJLen8K28MQqzzw24
D/XxlHSd78zUm//DqbemQuIJhETtJcbADHeV9aYbGK7NoBkp09ILJvDuSwwE+pqy918FnG553ryl
Nm2B8N7ETkSodq6XB3xRKylIBx3z8zNbV4Z6HHQ5syA/9eUiIMnBSxXMbGHhxU7tgHRBInPELGOQ
NQ5THALUynDNvotkXCXOTLvFNhhf6FmemQbVCFarwRMaUbQE8ov+dqNd/FyRYCnfYHWsI1GbCbRY
vjeix0F+dmP3W0rIsDwX5kl2Ke+rKMqWxheVwpcXURXmOoAArlgUc/cRmPzyBWe2l+ZqPCJr0RGO
pX8VzUmGFIm0TVUL01Tkbqi3bLql8zJQ0978cSokp+M5Qwoe9u9voHVRjkhEE1IdSIMizT3EpX83
ZicxfZiAzhLswTuvBn3vDkfHneQzPTrPKUOJXx3kx6Ubl3ku6h5aLiENARuGfVFJ2ZvIxIsAMmam
U/xcnvFsIuTcUCT4jSVMoGbcBD2oNRto7YPUKwEWpmNn4dlXGS1/xYaF1wcX3GnO3yoe+w056yr0
kLw253OuqGBJGivvT0w807iYX38IyURNn1BpNH/k6CU/bloKLf9lEq/2PLGm9ddqkaG5YLAaXlRM
uiFhJ3Ruo36WgDkZEnuHEn1+yCXlrFkgvZ1le47YczgrU8hgVi8fnGEIEP2iV3yhDx4ayYlZqA9M
/XL+9JjOszOXHZ8pFPrjc9ulGXcQt6PbVzoYfQ33EVrnQsrUwayWdM/shpkso6SqO4EdnJBrbMG0
FD+2hzspYqCQ3YNR3MVb20Yv/IFjG6/fN3u7MiPRwlFS8JSIIXGXDUdbfU+zIMFDbem1c0hfBaf9
2JQNSe6V8qR71Z8A2EOavNYqzVIIcagEMmPYkYSe+9SAtHmkAw8dzONyyQ8UaKQxRmtQ07nWnol8
tMOxXKr0jQEJO/A4JvnaS2dAstSyXQcMwJbcnJrYn6B9s9ZtT/CfUB9zJzW0IbN41jswBbkCW6eI
uydpfzQ2CexImuyZrRHoZEaVl00BlzJ1+cc5Q3nX4iBTXIWBAdCT71kZ98g9yjtHYJenoNGY55gP
VLkERtuVjcj+roNmPwJu4Ih3ccRmndFdJ2uXU6dV4m7JMwyFcnoNeACYfx9ET+ckcAPolFRh0JI7
8pN1mHdVaXcb0U2npiGh2XpoteBJJC38OPdn94VMQMJWdZrKPSTI2sX4gIMg4NahVKb0WIO19Z4i
Et2bbtlqI7GgEQs/hwiJmWun0dz6JeFiENZSjvHixSD4he3MLfoUhTas+xhKprSg2qMCBGYlBro9
g/86KoZQDfEP3pLnLAqfxxxinfAiLGLFUiy3n44SYtJ7gu4mXrlnxzYKGZ7/5obtKwy5pAgOsNnd
4wYBo9BtuHVUFaqUOW34LO17pKwoCEDS2qtOWfy+dy5P2wT3U4x8jtSx3Ht7L8+a4kwKROdJ2Ml2
fByfysevSk02RTyGdk2Kx9L6SkENzLuPEPZ1QZydGkn0GOzzBbhpNj6156MRDLsGDSPcgSVWy8nP
blYkEjv7llcPiV5/x3C9VJeDfdLHY7MAW9HR0YCdcjBY6ynIqLJG/uB2Wk82g93Gus0wjGSTSaS5
nypnmTPKnL9hMV9xjbp9Le3wo8HHybz/i8N2C8BD18awcnyAxWADjDZNWrpkcYeXDXp95ALRkT/d
diNHvkk7hqIvbzxlQkH77wWH38KI5pG5pzD2lubZsW/R5sOkOGVwej7Gmo287t+lk3RGZdnhhySJ
xWr7DPtj+eWixl3u5B8y74KscfCN4p+aBAaSSPyPWi19qDGv7CdM0NszSAQOUSNEyOYE97NtGZfd
qmEGFNjSFjsXpyShDPqSYVZFSHqUwA5i3GmflS/RsIxxr/iUtrrNStZoeSLeWFI9qvQrNxcfI0Oz
F/wF32d3AuEnaJRWM9/+HFIMO9lF1aHH3yR5JxfRB1VPKj3qxYri5HtR2sOLkz3u5mFyuTl9e6xj
hfX5OQCMy23rcHHrbEJagX9LjVTQ/GWoZu08O5Tv3/qKj1AxYPlTXxolKlfUNEsFC0aRTQAA7EsS
bW/9xBA4Wozdr8Y74eK9ZFRX7LND8RRjxj/fv8RNm3oZG5yxk3+k/QoS7WofCxS/7L0uWW/CfOsq
vY5/JbSMEjyCTBp+BN4hqwWK4vcPbO9TAEpXw5Wva2eF0vozaxyiFGaeQz9OTkJcoEq+rACJV3HW
i9UOu2aVDEHTUnil3t/jUid13FY503snOq97tDG45qTpGtJ1YB7IU48wo5wXY5mtp5KhrCWcKckG
Mwi9VHHAZPmaH3Svp51PkjuPRCjWeCjRf87uxgmBmIfpt9gFLQ8tNd54cm5xbMJNW7PMzF2dcQMO
XTQtFvacXVThB4lbBWxrov1E2Vl3wojsE/m/zeWOM1jwuQl4YaVwpoLpaERY+wilA7H71ie1Y59U
V438Ez5j0UAY74bo6O8nSwWxYd+y+/giI7I4YRCtQrsiCeE//HkIuhLFgz7MOx0B6iT27j5WLwfF
ZWnhtZedbcHmSJh51hwQ5cPbkpEC0gT0Qf1uc0w27kvAAbnEFMR1wrcEWDICs/Rb29Jx7+WnuOnx
nkNoQpR1IZOrQcoD6c+AZfotGgU9XWfu0ScHqUFfEPVnt46/x4uS/ipIucp7QM4Bh4hkFfskLRFa
jJF9QnxQV5XLnufi77oSkGs+puGXcvrKheRD4Jw/nvfYvvzRn3QCc+1k5OwcXyKliB6sZHv7m7sZ
UrHAuhwH7BKzI/0Q4tON958TUiGW555n7v60ZPfy3FAr0HWtXNJAKdk7siFT0aGCfwXio8moirJO
jSBNc5NjNZBXbSMxahMnpMKP3IHH8VHsMNnbxPwvBI4v1tsSWXKgWUc3/uNr0yPbHvniSFTq2TYL
f2Qd8QICdUy3Qkvx7wCWTF6DXG/S4rE/FyUBg/e40hgwlaErJs8qPSDwAPAZjFJf2uHiXx+WalRb
XkBHB6pPAhzw8juOixB92xZ37sN0MbgB40ofRuHtDkUJsfjovbShhXTvxV/7MhXe2+X0qtRCioof
pFk1C7nccZAU3TNRyc29XSoPjXkZtE5WbzyVlRoKSbwSUJoM8fr7BJQo8GhyAHU4Vq4koDX2ujnl
AnS04N5ml+HWuyJOEVrerq1yBQFhAeoWxCDNLD1C110BNubgnR8IchBy2BUXUgx29ZahVyI+juwb
u1CgmLSrJ4jUp7u5OvniIzDwkBlTvpzyvoRcLiEgIsGkirAbq9mNk5cJ0f7pc/tWdctyOVzfVNef
uUe1G7V1YUK58xBH7XWFtnB8XC9xgJ8kp2FZeKrjkElBLpg72qDXqDc79yTl/MXLYyunqqxyO0J+
i1BsG0JXnPKyxN0vjr9i0MViA6Y4bJiwZBhvFpU4b+u5tN8i58sHjzmU6eSpDYqwRxikwV+UQC47
4jOkyHC8Oej0ecgUGl/oHy+JkUrFCjg/gU9sFoCzNdhaoqMNOeXWKaxvG9zBidwl5lODjs2NzRKd
Qr95OFSMtZghppjPtAoqTINfw0j18DVuryv3XKGoIQBd5r7L1c2Hrd0CqMwrwzSL6QwQW4/tsBfp
M6U3/zP1LQNbPHAeeES/63WAnzCjV2MLkY4vHugCzwRctMccx2d5R6oaz9zQq56JhpdlLn+X3K6J
eCmAs7livDQfiJVmfhF5SzImQ1actXUaS4PiEj0H8Tdxtq2jV3P4SjRXr/vGMtdoSeFhO+Vymw6S
DzUf/Lr7xSgHiHNAh9CdURf7rBbeq9Xz8j9HHz2sr5U8hQMRlGjt7PaR0+nFz5vHM+ggFKYSTKjs
bhHBrnC6oU3A2tD5u2C93ZQEb6LIVEGaWVANuJyp5eGjLm6MlaQp5av/wPG+mn3dW5nAy4jBvYCv
Ibf49gAIb6qbgrfBVVa5UnH2HOR6Wmo4aEossSEkU2eqivbBPa4h5cqyweijf+H+bHeJBt1BIkc3
YBIxLBOmdPlvCeAxFjF59rkmHvyeHCvAJewih2c4qtuIwK059m9BsclIDoi2rLazySuGhRf5/1g9
kn3fdxLG+BvsIEkhwF0Ev+EacTwULp7OTj3mo2HzLA0mijsZarKWmcM96RxH3mjLtQ1Ib9sozX3b
IcDwUl4cG5qlcwwMnsvp/2qvOEW+HByYaxMJio4YsGD3f1JmRtaV34u4JE9II6V7ubCSpVFlTnk2
AdILgmWieH62Q7OqlrLtziE6Vlm0/nb3wbJPV+g5Vda9ai8lm1a1wd06K+lsKWNyKxZVNP6JQmys
EnCvkwJgMyuFnxNRhj1HvRH4m8LyvH/q2EAg8saKz4maxl54kuNAxC5tXGaMottlNg7hW967axgg
2pPEj3d4FPPWpGM6/ciqRGdjaTXAt2o7Fjh6xWZYslvuhiPdXgLRw0RLjhtFzmW772zHsKwJf3vJ
ACyijqWN4Js8DRVWSMOSO4GyaGSfd1O34dyjGk10EN6KOdxbTlUNxerYRL/VZPqgo75Tme1u+NP2
HbXBHxS9AfeVF05pDGtFl/PmzZa1GSBguZMY0/VNl0pQE1OTd9JtOgJImX6hopz1VAg+qYwX3W3n
YMXIURShYgb5B96IUL0T6VCj7IX+GYowLnSvxR87UFmVzMUcjtZQ5Eb1Wxe6GB/tNw1XuWFluuIX
E+dj4MxzOFsoFKEEsrzCdxmwQVdyV39FCP/Jhtg++QQttWyiNLXhJfv8LuLuVF2VAjUb6rnISSuK
d+uTVLsf4NFgYzXGSCJrRtbeBpFz65oxqL0/rilpFBF6dAfJd5xJszZUCu6b5Qf98VbrGXSGhF1E
eU6FQRXRELIpqo9GnZKFMux2o2f7c6b+TWE++TT8hPGyXEdry5niKvYAgxdj7QKTfzII79sFiZZz
vjAjZzGqETrgRe7U54fTIU95c1a6u9F4F84eEpRbjAkvzs7QoQXAStodUTZGilCCxIMnKRSKmvQg
ijj7QGw1Xt5T+IYiQ5uw6dUtBQvPNyBAyZggm+SD+4roYkwaXlnJFMOh3pAbDCVK6e4A1r42oHTz
mx2VPLEXOpG0FVHBvBdsRAuYg/nO7mna1gNLusROWWjVZ87q7vhayY2UVhVXM3K1+KvM6e/DMl3I
d9uzbaqXWPdGzbEXAWFv8Cn1IVZeW+be9mQnTF8hEI6Z6Fy0WM6+K6mK9WHjT9erz/3kJhXUa0p5
Duy+c5pn3CPJ1+ngPKzvYXl36Sp2icje3LiAG+v2mSgC8xqdr7Smgm1WeCQjKRSkl5ZI7Rqd5cve
iDvNTbbY5eeeYNs7iJGt3DiDUBQT+N1gY/TROWf7Y9n6rjUFMIukiwBb265eA6UKFwI/J6JvrO+K
yHsKDQq49BXdtF3ZafYpEeQIzE9MkRRSqi0M2kGulEl46uYxow9JZbMRzEUY87nCiDuJj9jAoHdY
KPs0X59Ift+ilJJeDtSIItnM+yRr04YveqCXvrFaylB57pvtkvE/ttvA5a5yg9zJGipjBYBjbjgT
gA1UuNyLaA8g7gSJQtjFXfVx+i/IPRi/qttzW6hIBROD5zJPR5/VBgIZIjlZ3Rj9l9x5q33x7Ddv
QIPeO0Wd7x+sc1fp26vC4A7YuGTiilo5OKX9EZgYf5ykRg4BBK1DTLMBoRM90HZVFi83wbI7ydxi
C3q8lEpbJ657h0AP0FymEXyGjvTn2YF9KlazFCGRfKZfLDs96CMvHwR8lLjV+GxgRp9AF7J0gCZL
f93Kxv65/HdCsjR/NgeC/cqj25ODmL33aiYpo65kehRHKvgu6GO9bCzsESrYsLD5vYdInJkFFgTC
kEh4BiVj0WnyhRwHuke9XEgQ9sHGyDoRYPoEA6w3Z5fTrQV+z0WqmF01G3OE7Z1Gkm3F3pEByAOY
Nn94K9QLaCGVqMnGlyX0yBn0wo1u8998I4dBrIfGjEjcteErgKMFCQd6aAazSTlsS2OOxrR1KDsH
dOMPy8YyaBgdx6q+SJPhc/4AxL/PrrAZukAGJgNTBg9/ZghvO+KvccDvI8KY+bHtYv54gW51uvwy
62GYW5dVOi8fcepueIItx/XFJsppfQ7nmJnYQdzcUIepbhLrh3T12iuBTTOO9nnJh5LOuGOkmLpe
O2xej0uK6UD2pF+7Bw/WLFutjUslyIyhCfMCzxGoCB35hnNjOyf9P+ohOBA+xWqKR3dCzcoemPYE
rLj4nWCaA+KOVfIMvo0ZdzMUpdp0wkeFtDqyN5CngiO7mdeAwsuZ4QGX7ONPULO/t9QyPR53Etyz
Kuei/j55nMbyY0NT8LRlA0+ZOAxn866vou7Nc0bBb5OsWR+S/nM5dvhy6A0Osviy1NP7BeYhKIgI
WRJ7sUyMrtFyBBgdEF0isojWq4CrOYc6LJGor/2ot5HB5KZnd9X5h6wzmLpflmezzhoe6frFuXZc
6EyDnMfqrrYPwyY/BGoX27e4RsA9y4Q3sdoEq3uxM2y78439URmNJZRPNEMx5uj2gEvEnEkACh/y
KmI6qaVLVL6jiHkx2J6LJaE5C1ZiHCbkZEqKWxCVsanoWKK2uOfqOuNdqhzZW3kAiPfMJ5a0HHAw
7NgIGG8WCWkhxIZ0X/MsaKb7NOX5g19SWKKElgcydZGia7Di/RvXo9XZ5t+mP7Wxt+j8rZH2VqKa
wJL1pPiP7P/M4d2Nh0n3tD0WujgeV3dKDs6lvDa5Qs2SKyNQWQLSSCHR8wXuOQCgpp2eRrcckKfM
021yCZ/8wLEO2LL1Od12ElgBx1tBJwfX4hAeimaqZT2RTNezBhox3N4f6QhmSAcLoSBx9+CrzMko
z9JLNS7mMQ/ggJ+TlZmugUA7Ta1DDkGKJ3B4CxcWAFg6h+Cu496qXRnkrBj+h5RrtJPn5QZ+Ggi1
huLu1xzmf5zxO7EWEVTsfMEwB/QkIYSLwnxnwFo4UK2ZAmwvvPkrAFTNCZLfS0Unu26AAh8DGkEr
QKweHjHzJIa4gMaxixkuAik33d4Pq+TwTJm8c4NI290ZYfPg2u16QVun0y7af33XbHNwZ8i/OVr3
AzfyyyBYyk7FiiiRZtVdZ8L8IWxfWx8kB5Z2xGoWm0hT0uKQntdOSeWK6vi3XE5NTE/h+qUB3HJf
trsbJIWdo1cfyiXUva8VO3cFSkqC9Fc8UZWz7mgKn15EXxosI8w/le5D50QJurcRe6rLq0OqsIFA
CZX5dpTkBUukalH3TUQ9nZpYbqXvkWH5YzkDpndX3mhAUggtmHs71n3257DBzcNI5gIC7ek+Vicy
5DvmhoHWhHOu37+0tzCjEHs+ucbJjqMEmZIkomtn1F8SlzDnfludpmOoz6W6S2gZ52mZ7hEB91yT
cDzjN5TZcTQg3v4YwGcV6BZPEUv6UTUB4AV84iigCkrGroBvFM6RzLLAfsgOUvPMUs2Di8lf5fMu
nO061ItGjKeQSMHrzjFoBqAYIEeakWzKdkhsQ5zqQnuhIcjk054gknNXsjtrqUgG4lUPFUtMtAXS
sRDQsmEvUoHH/RVvhZvwvz+zM21ZgEeBaq7dKQQsEUT8xWFPI8dRj6t1ShxsNYGiZOa20a3PLRjs
S4ZAGwv5gYr3pTDePmSY4Vw2MT+d6VTkivxjqamSNyalfDGX7y4Mi112pzHfTKSBCFh10CcY4/Z2
m6ZrSJLu9cbMm11p6hpFowriNGC+xrz/4IJe5bJiwaQvx21Z7awFO0TSnKAE9ovLyMS7a8DO0alj
WVkFUd/RGAuuJ2xLzK+of5wStBzXn+GXys+ZIvWr4fAbgs8jAq4+DOm/vwNaabAfPKkAzil7QnzV
MrvLXNEVkDIvftcXjUXb5JQqD+OQoDpYcsZyX2hoV3eyYS6lIkKk37coXqzS9YCbbMNOoAE1Rvdk
9jkN4BzBP8VW4BQhQqtaeIYIwvmyxYHyAiGelWeC1SVtSObtS7gE6ZEEz/maRgjh1ZU376gOL3lg
uVYrIZ9FYu6Yy6hzM6krCtVsRcfM/2udnnWjkdmulBr5U0vb9fdVYcpUZdMt8P92z0aseS8QwXUW
3+nG5aR1QLFgDnk+0sNr5SHoTfxWbscGzpcr+JujMD6rObKNkgW1wHuRSm4M0DLOUP9Ybkwl0WTI
+y6EfeGBAQZY5YhObB3ElszOdZnJHMrc6vRV+DvojZNIB2H+4+p4bcG8uNSUtU1gHFh7i6cAxqSz
nTHarRZadomH49PLs+/O1R/038P98OO+zBqmaSVhDN9KyLyuLNH7EoYzMCJXb9wnXHpxecHh9uA0
DxMsLRI/FCde+yR2//U3e1aVyWtuEyGlVQECADB4DJGvGi/TPaALhV54Nbq18HEKVu563gK8SpNG
I2v/uB54JOOpuiRCzX3wsyIgST2mIecIl20jfhik69qap4Zoe1BRDdqPu0TwtY05meb3R+EsBgmL
llLBRU+WtWWALoqingC7dOSsNKpmVbihgzqOzRzxwbOExQdLvPWEgeXeSp4lrQbeEHDtnQX2Cpb/
lLw0Z1Lvb7F60xM3odG8fTik1kPI4xJ/DKaglqsWequzBoHypAOllnPxCT3odDNWZ1B1tXCFoXiD
mWLVDQwJsY+ZEFcgXMrXiLq9s5oQFekgEgF1f5XBbS7+wDvQyEVjz7bsLTFFaDvAPNN5Btaa5giV
pQRJ1uc0tzrQRRTInIno53kMuLY60esVDaMsDponyCGbl1jtxdWslplXfhv88tEHmheeVPuFKq4y
tWFMDSQanLWRXKfnY6nY53Sg+Dc84KcWLfw1smEwRVnnOErUtqmo9n1PqeMrPqzHz1zQaSo9uHDM
vuyg0SaU+PymRUGodQvWXbkrFuY6Zw0ymVQF6IpzrzTi3PsZAMAPmSlE75l7cvczH8yVidLJipps
KoGZqnhXxEquGNnq3JbWNrrer5hEUHi/UcFcs+t+anvIZu6+8cM3eTBdLwzWv40wJ2dRqZC7TWB+
97NLqvGuUFttkPxhshCko+V/+U+EqETtS1b+exg/w2xsaY+PuOvRV9LHVnipv3m9zpipUIdGPgCd
lALw2gXsYdwn8HSytT9eglHKz3BKEZTE78dwTQTRKsKdKGtwJcMsz0ukzMjhf5m6Y7F4MTrq9Il0
KGXWUQy8gZ+oh0hBxZodHDt6U7FGIJoUX1EH26HN3fq/y4k42hBlAvHEAjCGOIZTwg+YHaMpAfk4
W7rAZVhxB/JSa2fOmhjyFhQkQtpV8CsPnm6goqalmeUVkksRjyzxCYwwsFEK6Sf9Tb3sNVbPc2GM
z7Js2TmFgQ2csYD1Iwv4OqATG2ra0UTcJfWR7fKn6V5GHO0goeOoZ+QLtGr9XAvIsVtI6hzo+JhC
8xh4Y/rE4gNr5Sv7jCwi3b6yhbFd1MK1EqGpLCO4fHECX8vLs0lbDuubQuQLWiB966a3gEnBvt4z
ehuILAkMnQEl0A4YP4ns8Gw/GUUffUjQLrOD7q8eRcuHNm64buvknv8Dhz81jI4ZFVdyaojfqadi
E4qoxFP+zTyMWYkzWMo60jtKXGzcykMXaXP21pA3TScGJqGn/YdwICyol/VFV31qRdbSe7UsiYAL
QiGIt5odW7qCIte9EmBGv0hDymEpDRQeEpp5D4YQxdo5BuVJKLy3VSvN9h4S+yJSxYCPXh8s+lvW
OVbRVB7UDhh1IxcHfSMdiJ+V+VIr/wx513jYtROlr/WoAtCdhuVcgkJZmy6KyAGPWAWjF9IJJ4sY
VQGqDApKVpfflwcTQ1kfbVYnAwwA0/gvui4O5NrBZ1wnEOa7SVpw254fC6zGYu7gXyVB4f8uRBnM
YreFTNG2PpXyw98M8L0rMZ3E5iNw7oA7yDUPg4IFKS4T4s1dzhOJ6PalwN5vP6BjFbhtTj1D7w0S
kkpajBV4+psmBia3GlKTDVpxBcjt61bv/pTxPni38TB2UXXfkiHykbck0H5Qxwf6PLgmN//tmjXP
8yermD3BCRggC4cjkCstdVqrSjsU7HeQkoo9lxEk/DTyXJu2CYJ5wbUsDxZTlSScJ1krNcNcEWH/
eBvZERH0PmUKdDte4Mnd/eokFnArHkW5cXJCHWvNJ2ykz/eQQjz/ULP3eZ1SNIVaH2zoUoEOjDdc
LyRGS1yc/WU5709ysZv6GBkDyuQoWAJFm7GmlxuIR4WTm83sAAXSLnHg1URUSObB2tDUCqzI0+Hh
NVaZ3wHzKLHczFomM+KdqN6BrTOSdPb0TvTOOUAGycrYfMFph+Syg3hZFmiE7vwzMzgKAOzrJ++e
BHRnU6NZQG2D8OI4SIkZJb6lx8THBIp6+XO8Kcl/GYKFj0ccgc+lYBkugadavhecQJi7xIiJUF/Y
0Yf2aZZhKrJa7NKOxF+zbzRkpt0Bry3YJUtcT8+pe8RVXslYTE3H/SegK2jKnHe9RV25u+0bcq6U
Cs6wU1d488rt0AbrrrBJpARoP+zjhOeaCsdU4nonwjskTeD8/T4EiYjW2ZDaLDTkSxVyQfgApb/l
RSIUhC4kn+ggoKRBlv75vHyArVm5gUTp1aqHhBFYsT+qASdygL7yFWFLhfhLg9NCLrxV8/ZQjSxi
UKoHS9dQ5ZP8r7SHJxpQgSHBQB3OpPKPnHc290Dl1C4kOhFlkuONLVy++Us5/hELhYLhSDBPN3El
XyiAW5npTYf3CfWG288DjvQfspH18A0nRFGPQkm70eNIG/sMzQ33VpFCn/2fWWfFPcjf3TAHwRQr
726L4UDWD+fGJVLOVsTzTkZ7JWnkyyJ8cOPyOMwQEc6qyW2HEUdGoOnwKUW56lOmEWoPo46A6fEc
bUvjoo6S4tU4ktSxiuTYxaIelbmrKR1iSVFHVJ1WAJpQWcTxtdgcYc1aHbnSkIe1pY25Ny3nOHWR
T24jO/gTKzhPpu+wVH9VwQCVLkEfqPFJ0YNAoZK/bGk1DOPa6b7JZujHT0pbnMfmgRalCNTnMeFW
Hs6D46XTOqKBLGGToJ8j4WO8f87vlsGdid6gqvfkTebStGlDrVUfuoRvNftTXwTOZydFmEcwLURa
c3IYN3BykDpO4KTh0FAcoyRxsp6wnDInw22ESw6ytbUjHKAgYdc1roSkyh1/RRy87hsDzHvb3Qcj
fJV+anodQOhzBaHP6fkvJUL+3iuRFCIyYaMW3IasvcsKg0jvPAj4dZ2e2o8ryBNXbtUJfvWoAvRO
sFieHqLsuVhNYn07PCd4UC1eMzF9eXNsrMVbu5aeyGYdGKctum6rRDf1krkdd8Ug9ep6PeslYnRa
d/gXVa1LY8hBAySda9MyAn8FsYLXWJ+mVeWOxwO8kAhpTJ6cL+f7Kp+E64YEsUqszvXn7uJ2BZCE
xfsNTgCJ9lkpE3s0Tz458fZ6wdHb2dKTI0b/I9Cj00+ZdyAEiGuOkhrqDtjk6XdXqWWiNLuB7tjV
lBONZsrfJJT/rHyywvfb5+vziohokUY/JlgRukGjhcNxlvF3+2CvYrka63QUNJGfCsrhn5FcWTM3
XDEL3ZFjOrZjAeS2pBYOd9cNA0x1tDvS7JwZX1Gvqvi1fiUxE7QEas8jBkWWQo1Qr59Dvh0hZ/5t
gR3gf7fWMa39BCezpBim1Osp2gf1QVV9e+F/gcdBRAfZG6DRVansHHCaxn0SJcPzqPIIaje7Jan8
8LACQrJj9XYtho7sujkt5AFx48Yrrf7S7ju8FAhkVNGPGm05CMEZd35b+cUizztBYWQDvdfybLuO
FtDF44j42rW0/VNgJdEVxDVy3VN/NkdwdWG1BNqcOrHN2IplmGxRtWlV+2q7qEyApyVJiPVYJGKE
HD5Uto8yRLLyeWOBASHEGoVz6cMyGrBQ6KzCwjIyVck3fCHSEhRixF3ry7eoCcnTu0g8TtFtj4Ov
/FIbqeKUvFBeju78QaZQZ5PoF3dWIF/P2L+gOnoeAjuXW0nTOtrpriujo7ALwi2/C6wh8XLjABIW
8jzkGVhjwo2AnZna1M5dJwPB8dpigytFqme194ZyPxpk5OC/sxD0yW71g2peYJj8ICT5fDDVQADX
9IJ9LiYXUkTqL4jJCzi8P7oZ98tlIwR6eutKHDnZDDPsimA0iLJ1qARTTqojJekd2BA/hPemPvKL
WEZLuG+rPndZqiS4A3ThjRthY5eoee2NgJ7XrJaa2HdlMPax8Nv4g1ETl4eQncSgAIlB757fkDBh
P+HImfHLmKeT/8Hqq0705Wj+6w8Z7bzoN9fcXnYv0TnmDDesaLTN6lDyrpBHKCTii82VKIKjFBrU
OgrP+gcj1xIp4FwVEcHMeXWs+fIJAqrS33C1GuvLJ0dyHtTcijjnMhBUZhfR3rBIG5eDWl8mx8ma
QvdS3DTW5RpByM0sqv1hSi+s3dpUmPRx4eC/Y3zRLpweDif2vybPoA9Y1wP8UFnNtcYsHPGlzgM9
UTnbMV6GAgLwzQiItEGEmmAO918pEsc9ZqFX9cD5XcJcOBAYlmbx5JJdXB2UgvGXIaFIqUhqdq7q
myvM+7MtSI7l/xZPs52sOZCuLTlG6z6sFOL77wvlOSMvGbso+e/2wWFTo2Utp2oSczXvKcX2l9m9
Et/yK+AFbmeaoCh80OOIoke3cvy51cAs4jHxdAqTrllEtK1RI5IPq+jXcSt+gkU9gv35HJvh1AfX
Ll7liQ3rrA26g9HmyPPUrW+J1H7hl0wuBlkWeSC4/jLGt/bGnuh0INKO6GOC3fV82h22nzY8rlOx
1pXzMvd8vKszN6zqZGknpYsPwvKgsmP3MW3vKQU0110aWmqQKD6unsvoHDTDNEZB55PpsU4kq8B7
c0Lct1gfX1Ds4mbeyFjoQmfKdq+EVDPnCM36fdJwj8bzkFZEiiHxEDhibcrgGJRHhKaM+gOYKeVf
ol5PQcfsA835znX9TsAN+v+UUHnHLb8qo6buRkojXmbs7I1ExsFgvtEqlcgpdP1sw6RiYkITRVtV
6S7lS+8D7b3/Y2g2jvIGdnR4JLR3dzpWm5y8b60reTgmtmLeuFUv0wa99Ya7/1UnvZ9bPZMyJsAh
mrvE3iG8YgLQ/S17IK9/jdFKt5f+CVpHjTNqMskeAuutJqVUqyk1t3dtASuHpqb2rr5DZXEwcWSX
MwPph1tYw3dTWF5lxj7cexNq4EzCori4QjGqDP6RgyhGzVPVmHIGnPCI06iTwjeZfr6jA1HHB54b
YPQpZe7vPMYK86pIrY7912pBgof3rgwWqcdghLQvf2DfU9G/By/U7a9cmx6Dr2/lxbgBOBSdKvZE
bx7dMav3LUVd6jZMviaKSfQVEwBNPzIp1OmZo5ttJwG0tNlMMT5aVyl3Viif754aQ9ikJIHOodw2
7KjWGvhF6wxdIiUEpPOs2Zd/W6+oj4mFhCubwG5VF3gIdd9pHZ47YLOZwgXp/ISJGZlt7jfWmOPt
G8k+BkASMwuH2AIxl4yiAq9WXmrt0ORzW7WQk5OxAs/XyYmR471ehy3mhdhb2D3qAYv/TEHmInxW
PCbPe+AUgYXYrDOERIOO3kzFNns3GVJO043vv1I1U8F3eLCji6hOInjjoYVzn4VjD7eb8TJhZSze
pDbX70CXLTMjn3rMG1xnwCGC+3Hf7tBqSPfMQS/4YCC2TO1rCA3+E27IcKNr9ATLi3jin5T9/nF+
fDKraVALDqsx2DhYhKFQcz4//FRl24Hxrvcdp08wYYlMaJI2RPWzdpfd9KPEhErn6Zg9rxKnCOfV
mT/cYhXha53JJ2wJfkNYgSGr0dHXFyd5SiQZuYh3E22DYerVKoWV1NWxnFi7JR0BEtAumJOVzuSf
V16gabpHkHCE2KJcRpB8iycsoEtWGEavli5G/t/Amkq1ayotmtYBVbWYWtdhNNvA4kWh3srEG7WL
MjYxyFHAhSdSlyCLUKmmiOj/zFWdvi783TadFrbfn8oli+6OHRUy+3V/84ofIgKZk3sroBxSibXa
cdqDfvA2Kv4wVw0wRSjEl2K2tLV74A0sUPui/JjPWPwdXQNFeBuCcExuqAxWTSyqIxyuGknWRL1U
8C+VQtV7ef0AXmvlTLwjsiywxBuohHI+XB1bTqa2KQIYTj/s2uIri+SaGgauIk5sTsTkX0YuhLnf
BJJmvlFODkEG88nlkJ/MlnqeqI0WYO4Qt+S1smqCoo2v66Gb3zktQjUGu3t5jawFFNfiZGMHHmDG
ilVPGIOyoUCw2oc1tyI1qjdadlh9YVVqIvR3iCsY6luspWMyeyXAvS0LNa76956ckmYnJwiAfSRZ
BW0jbFrPzPM3KnHFFFJ0D/EEZtZM5bGKHXUrG+Xp5nkUwWYHzcStUjMgtZisnxx/6tfGiYp0OKfK
Bl1Gsu/6okUc5We3qFILjZWauDc77hdkx6Jhsj0Y0iu+ZbDnk+Hj0xE/IVrfz8wQNPN6AaFybMkg
z72aYFFLpE82UO9C5qYsA216tRrg4bHnj//pA9mTU8JPnF127aBe1ME2PudquWGqSrL7KAm1gI+d
ehweodiFDWp9fHH1EzpLpD0a/Ayq1XM4kzYNjXJduunoj+e0DthjSPo0tk6bsmVs5Vwoaw9/87+H
iuvowRwNHg2NNw+xtSLm7mdV212QSZfKd8990ICu2Eyd5cFHBXY6GU5qdVoMDawoSHYJEjce9AoH
//tDU2Sa+zqd6iOLNZ154jtenLYbjNrXvusITObf7ujyr1r4qILPAWwkeV6JdZdnCc8PcyLKltfH
tIVnnFOrSumuMijdV7jb2amfW9Lk8lEvMVsM91x9iWzMxdgADRtQqgsM3F98KHX705A1abKKaiVp
VZYIYq/++GZWy8gcklYnM5ooZoGIWZ73MMPJ0X6Fiqqt83BfyBfl/9asAHnnnaC4Y2+DYlYUKlpw
Cl1L6v/JevDmbnPrUeAjpGttLzNjm/Ld01y1Na/Vwu/IOoSIe7iy158/kMeEAJUKCIfmHWVkcBXJ
tVR7tVG/sGg0EEYAsJ3gBdlyg6etvASAkKW2/7bYJEImmwvXlgOO/8XuYezyrat516aQzXeiINqD
KjOMbLOuMvFNGx5r0Dse8WQA3SbNcYTKpjUzTNRgkkwQhD22iQL2oxcQPeLudablB4snw+eFwon1
sxXnFK7DtpKEDx5WveflgWkhJpZpu1tTKd9mCa8+mL7Cr4vul+uWB9s8RzDeaDz6fWTacU8r6HE/
e6PLallCTsS3KuM0LfzlN5oqEZSm8hGW+QYvO/HO1iQCHCOPEvEX7RHgUg5gHjJcRy1r8VSk9ExB
TUt8YOr0YHxueseCAbqBVBq9foL0IRW4mL4+pkA7QkWvlj5PsOICismbVznQJqjWc6odjmamFCvA
uiPI/pEQAJ2PAA9Q99BcXanQ+DX1VqRUyGWklP5WXaARbXvjlvYJDtK3xF0DK9AxAlfziDq2LCeC
Sevyqhm0vhD0GTIrQNWWeYWiSVCSPJx8VA/e/1/zubUuWg6vaoK4duyqh5rqpJRwJF7TK6Yx2txB
R21AHyadyirGxY6g/nLqTO47dcBkY8UU6Y/u71vqoEdlUaFkoqBV/E2qzwc+chOnsU0qSDA5dlZk
/DvET2/eWQIQDlutYU9R1RKzU+qs0VQAkkH20k2dqaXjYj1X6Ny8ZybZDbVm68GYeLMVi8Wr6Z5H
vxDpkhT3K7qCoOIW/lqfM4+lQ5IvaE/oyM3jAgEjshL5fB+9u/BFl7a/eopF+dUB/GHxq+r5SKlr
dwA/rBtlZSQSJAmvYJPmdgxQ17EP+GezxIoopuac7QZSVAMELDDKj5+tAIdNNGYFqqq9qoOZJbhV
66M/Go66ARXEIQl1aWB/gLkg/KGEpILMLn020Clnl1YvqEOpfvjGpAQHrI0G8HhnYFBM9yeg+FPK
CMCl7YH9HtyCpWMdq9yzcvhU4FQIpMGsHtxu226UUPlATuf73o3qF8xMNLi9fCQtEr0yC7dBwnDR
oGy2+dl9SC7Nb5kV57WV1RHW8Ie5rFys+vnKSiPeLfmfC1MHtOHpvN3TAC3tFduxSe6pmh6LNWjo
ZabXEx6uF1BaSRUCQz29vES2F1z0XMW5vwnHukhUg2IAx6L7BsJtu/KCSdhr1qYzVV3UZYwnTqaX
Cs1m+eHjqWVz0LQw2S0vJ9zyHi47ScpkDolF9bwIdE5H8fBoohAaeAaoyzJOLwQCmKFHKe/Vnr8K
k+YSaKDXIX64rBUKFP3wY34GbA6oUM1dcOQlW7oSeBpwAYz33TtukBJRlCJ0atg0Ei4KTlvyFgro
w8rVP6RyFUn78ivfo/3yv4V8TUSS2ibp2G4SI559TojGAp8RtKWIYCdB7bPaUv3EUcpAwEYANlT3
j78S5FjToAL2hLE2y/WYR0sMZ40rS86Tcx7KQYG6r1d179LxKuZh89ySjTnK21cA7d5Kn+lBBIiy
sLGzbRv1iF7JVml7rx1l7pS0hcgFrqaJ4SPxMJ/MR4I87M7akNt2UxSuubOuP3DloIfRW6PUdMeH
boYMulxCvz8dijKYuEG+BRdCAJGLSdyssju8XqH7qd4RyvTXHm2rwDV0epgiVq4Vei06Ppw6u73J
e5k+64tqKEXhKaH7upZL6WawtK10yL4vqMpG8oRbu/53efPD4DOsf6UGNQWeeZDm4UPTpVbIWDBh
dIX+CppMcz8BhUUxeWpzDYQIYFaiqaxB1OI2aCL7RTC6kTGgIV6mh/t0B90mGCLyMAkR5PIC1B6m
nrb6wxxdUtLjd8ZqLWxgd/u9ayaZeEwScoL9Mu1kkPyWVaUN16kqOjfAprduOrWh5KrabRz+rsTI
z9yYxn9wLU5r0RtSEL7UrK53DxeGRR9UwqMde414poo6w8qhZzHRweoui/B+OIGSrUkha6WSHkpA
Wa6K5LvzioN4fngp3C02CbBUr60/4VaONn0cm6/43ttqgXJ1dx+1SGFjhwmgKyii/asJsWCRiJXh
QEh0owYEjFnoSgZ9W2afowqwyyA3KjGiioSdwzdbnij5tWrT39qiubzbVoU0l0PB/AoPvZb9dkWP
f7p2uTiV7pgWdddpmTVDJ1dlEkvrDRmrGE4WBt7jO388FPj2Nm0YO8qxZJoXgRBjkVIDc7VASVEg
laq4LztdbxX4miwKm8MiziF8axOujonScYdHAlajNl5xuiJWnBwc2niIZ2fwokSW1enrhMjxV50e
vE+r8UlHcGfqCwO6p++2cnloFU1n5qM0tg5OQkDdWyYW8pA/gNKVp/mzVmcV/NdmRPXW5ADvc7SC
1WZm0wPTOq+U4ChzxHV4wd09PGVMvk79H16a6VE7z0UVR5DApVTQ7K44m1xb0t/0FSYidbGJc3V4
xLKQQyS5cHbeleEphDEVqK/iMvERpVng9DdniY0t6r6lUrKZoDVtUyJI9L/M1P+wHStgBz6RPEbm
VChfC7pEy0isugh3Jqb+tWvn+exlv1/tKRpom/C9ixGXglCnGD0mMCcr0bLvchtwExlFNT2uoxr7
z7aPRP4z3IhSm7anr5aCqMJ4ZOSvfa90QuJWRsmuusDFyuM6qGgRJX9ZHp9OgRzxEmCoMU0VJP9F
XM82Mo6GDvVoKTmkqJykEQPKZ4HoPLoNDwCYP2EfErko5QqZ8/x5wYnKMjH6coXR7kW/7B/HWzqL
jfMtEhjls21cBhJrLPaBblLoNiv1+lCaryk7uRLvB7ThSGrDp5+UEfni55l2OS94DaeFsekzTW+c
76K/GhMBpYf3yOm3y8RnZuuYsK4ImLLQkH1Tz7u691LHrDuY5zTjM/Cdq1WfU45Jf6YYpXSM/tVw
bqnTfQtWbQjS8bQ/HSpjbYh5jhb3W5yI2AFC8QR4ATtiYf8LbU7/+RcFkuZ3vYewRaB0y/itlwu+
8qHhKkf8iWySTCg7AuMOqF2fIUO8/50GHxqN0YmjXpPHr0kVUM+8Lxb/V2BeALj+KRyvluEgRMoc
XKbjwYZoF5zeBIshbEbDsQIe4dHDOYx304VcmmftpBLQ4eEKws2nWp0FJb45Sdzd+wscTbkrrr4V
OJMU6cdB5uWuUi/0Nh2rH0axhCZVfUfjQ5M39x4bUXRuRM/vzGwRrhKgVn1axpLRaDWj7AhhbQiU
NtLj/+Gy7okdi2C0VP/eTLq9pQYK+dKN92svxJjbTapFynsOhXmuCfpbbOBSmVuvpkMnmVf7Vatu
Jxl5E3bnqOjL3RNVStnx505W3EgHKhuBf009EaWXeoJ7z5R1oEZEwHrX0iawqiAO07Wp9chbGi2/
uoFEvQ4TMhNqExZTQaMLmRWTukOavK1qjRp4Rriu+lyIB/rF1fkUsUBoheai2QuUsEdHJsSSUSA+
3TFAQGB0pHj8Yp2aK4JSUfydXnnQvOUC6FvZESn4OsWMWnraq5YQBMzNWQVxvdtwYGqFBP9dzCjs
Io+WR/fUMuhbI3x7QFYDup2rQ5VuWQHGoMpGY4VkP45K9yAHTcgDqxdkwSdu3CPpGzE8Yp12Tqbx
pBnSwdPCIQ4s0rQQh93QH2ofkaQbl+IqKuwhvi9IpLz9KksKj45HKfxyNFVzCdf7YU4znqgWDurk
8cjUpZQqRexPEpyvv7CTSGS3DWXcGeucv0V99UBSbH/+kxPRGvZrfdveuxOb6Sx5vUDzH93sKCze
dWiehYLkXcAGnmd2z+yKmCRxYz+wi/Av42qr9kiD6gOD33/rWmFDw1BdEjxxfYS/YBnIoCQOJ1pN
G9zPQgiVZatHmCKpbPO/37ZKBZWyMmDoMEe74aAnNTjvjQF/uJQLUTIR9KuQf4OTQZs2XWxph60a
19yOB4KrZTiU+CnOvXnSCbBA6HsP4D72sKfcJoA2eB+mYYLjVoGLmd7DdcA4pEttsmI+KkmBj25/
Mm6OCZbfIka1nIz23RHMEPFtKWWc2dgQl+LCkbC6LUOrHFG9BKr6pdt2XmXyQxVQOiiiik3x1G+v
4lXG0IdkXygSmBcSFZegkGOqruqyfxHR9z41FFuhZ69LOZgmA25ju/S1BoqMGHuwEnDk/z4Ng2Nc
YjMTgz+pzMmn6FjmGvXrqOE/oYr+GV6AR/mqihya97h4zcqB+ID/6Eo+q7jUvP14g9NsFLXlMzUF
9aqMMUoT12MxVfMBcW8uXPM6cMSYdXb1WDQgRn+bWmVWmxVdLkMTTODshxblhp5Ot2RxWaGZjbQU
e9QUwcv+h31YICD/zggtx+4vZ1KKM+vlBLKmeirq4rrXxuh83zB+Ls8kohv1MqfOu+4LsNrqglbv
PS5HLu0F3FGQ0QKJsbT7KphbsP6vb/nwy4H6YlTn2ki/iSHE124whC+8k83jFNFQz1N1OO24WPZ1
Irafl8TEcFPJxt6UCWL/6j7UuWSIeQmSZs7GaQ2j0APi8aOqazcRDbtItEy8l25kvz6OCal8Fnnn
XnrVTxIk+0rANiMEOQhpK2QcYi3aF+WTv0vpjKSdeVtqJjhfz0DI48MUTaUGyVKfrVzVq7EhFNVT
CdMdAi0xZ7rQUtQiqBPeCMjK0vB8hCaWKCYOju/lWi9rPlxuMfGL5RzOdwvXbECJqp19e2Vkw76H
J0mzu2KOt3yRAUmBFJNs1P0nn6EUh3KWfrBNcnNQojRKuWhpXWgnXJR5VdwYsjb74Xp2I9jPJORH
OWUqOVdqIwOXGPR8iOjdErHGbEmXUn45MO+WX6oeY+kz6Y5PMrHAugYjEXGSg6fIkDmx1k0ZaIXZ
s/LjvL4cYj4pGEQX/1A55upNCCacKbLS0Y+pKqpe5IcNCqyuLgAxLrWM+J1M+vARqXW2pkjKWYEV
LfHukX6Z31+Y7eWAwaiAocNqG2fdd+6dChieoN/JPWC/HTPTi5/FtA6WsRLCiGnMlQFZ7weMh4ae
K2tcg+DansMQ8m0KCn1o2r/6cBZIf4gL+18M3eCGjOkjAEtQiTcIyIIokv9+4d3qwuHNsV6XN0X0
tJNUNxJP9nvMhAPWfsOsW/u9wOw97IGe/cbMaC6eOYpDg3afPTfU51gzXBHqic8U+VRf9KjGPmZ/
DNETecWhL9Q0iLo+KsZ3DjBceLzQUneAl+AVt5V4dkGQ9kH7HsQoGzjXMzxEd5gua6Owj44R8/x3
6fBCIAjIdAFPxs9ruFs7QmpXzV9/aH7ETOG7kR94dYaf+n2f3YINRp+X2ZhMfuCIoB9Zoit53ah1
9xNTtQ3f8qhUmOUGNh3wQzzz/BjqjMqnXbN11bP3zNapxSQow9aky8Yw+JsFVO6PEK8N0AO0Tck0
RQm1ocgTtViaaPiiQlDCsq1/0Nao48HBrsHTe9kwAM2ciCiZJYN6E+IWHbap77TLegCBw1Ai0seU
jIG3ktahJCPnPhgbaEVaQaG0jb6KeiCzHLEKNi75EKEGK3d7zOKp2hn5qKxhejM5eA7tLPbK4MCL
HLB59T2S4Jhz2WioaKfySMMmI7o7ZrvbsgeQ9Os9ih41gxMz4gugmwg+aj3YWB6tX5tIl47gl6AF
2CIMNudSeJjzP8M570fWhpNnhJRWsJOiUr//km4I6J77Nv7LOoSjHwkM7sErlN0DoLNReD5YS/5F
PWvwMerhuRPB7qn1IQXFwXMxoGV/2Q4XymxushuxhkZpcSs/VzExSsQr/qIpGThrxJv81b0iA0ay
SX5lHlhIPmzQszrXMipj36tgzAyFm2It5Y6PleXmXER3qiRimpYFSr1BTqwnDergv4kkX2jnF2VI
HbCocOQURk135yI6/F9e/NxvPkHkAc/0ZRSJ9BKO/985yvUg4LYMfgUrNnITC9hlzQBErofMSdir
tDohGNo7yk4jJhjtVonsqBeOQLK5+gELqRKVSTlco9XJ1RsdtDtXNobu0x8QtGmnn1mtdTwOX0tr
jBpdpSTcH5OVhEIKStWARVR2Xrjv8219BwsyBt7b27GTapQhVa9csGSKy0IxVCj3+ERgzIYr+2Gw
wlQZrxhHmsR/mwBOKGI1ouzxHJvE3vegZBq4pwkRh6//hyDK+tuCpd83M9O5cL3un6Js6DS+seEj
Y91NP0fUWhLpcK8HHF89JiLI3T4IthFa87dLNoQmyj0XdDbFD4Tzi3vmh+J4jX0nQ1xMzvk8J3n+
UDWUhrBmLyOAIKSiNEwr5Tg8DtBEAbJSWVsZaMdenFGt3SUr3yeJAXrx8zWd+WMXA2Xkj+FAQFuB
V767JNl2FNQ/asuutAJAerkz8kIZJBxtPDPcfeDhtbj7zpDSSZpHWRRLQ6uqpHGS7itQBV7fb0rs
CyM3+ajLqA1WwzDq/nV6MS1rFbRwGR1spUp2APM4GuKKifr3njDEilg1IlkyqtCPW3SPK4ZN8Yyd
51K3+U1m80eo3J/BIzhCVLHIkNdMgqC+vAQ2uODIDPJr9bQeS9R7kTmI/prrGF8qpdm+e9XRR81r
ch/DFMrigLwUnNy8ei81LRN7/RWj7+jeY9bBUTXlw19pBEcoFoE7hdU2A+26XzyPXSnDaxGiXbgQ
vkqXNHAFC7cVSvV4js2KFX9Y9QAvTBfw1CqpsGoFnJX8iisC+ISoNEFwwwkeUDdUdFAOt/R8eKeP
nThhQzED4EOV9JFBg2ligCGqz+ApWKYKO7pv9Z68uWjLJxK9bPDbDhX7PEg5TqyznS9ES1Yt7wrA
uxx0HpPWyE/cE+CJpWg9HPXjN+dMipFGJteRsJsQD3dehHTrg5M38tk3YCfN6ZJZ+sHKaB69nSuK
3/7x5ooSWkouZgZxKgZt38bKPXK1gQVIPDX0FrZW12XEehGlnP66J3Zrlnj45x2n1f9jJ7qN+fvt
FAVMZeMN05kyLLG5728nSJGNtfim0tTJA7fMkPew+VsKCiIDjwaAjrbLZnirE5RBUmjOtBoUmHOm
OBv7vwTrMpYJpjgjNSNOG7LkIz29xhwWwX+F0XfbISW0M4NZOCe+4vOxwq70rNF2gLFbakCU0HNH
xWRGtZEiL9MoH4Nkj3jaOVdcl8qtSW8ZD+//l4Fi56ahtPiQwC6+fPjb9nDad7Qgk68G28SAYZCZ
vF8seGeZxXHJsB3PU2bzBVAx/7FSjWa9z3GvF4Z3iUj9noUu1ZvEo/WMAOP0AxMW5xNJ8obN53n7
KiksCs5gz8BYdOz9mcyxqzxYxChyR/2Ywy89hLhQ521BJaElfcIF0tHAycnDykOQMIm4QGreKsdT
7gmYycECTYQ07WBLUmXrkGwAYLfLtg1nnHvjPTH+1sjpWOZLsNYtWjPv10zSs2ZiXvZJ8qWBkszJ
PpMmic6Fbes83qWoYk0DB4F4FOSRbQsy3mIPwsS76LK88dgvEzNxivmzuMLllH0/oHpNQE0cjpLi
QF5TCHRJE6ciLYod9G2kvA9tSb0MkLXbllrYIEDHT405de21tu27y4f2psBSEco9inGDzTsxAj7U
F0+5p/AbC3GpnknaD77Rv/WXaPilQLh1ByN0Kk34LNJ3eqfUKz5YFMARTS2U7HAZjtnEDxevGgaO
0Z5mCSlIKiEY1LveHccPzLlk225A7Bw4dJMOXIjj5ZsXrSrQH+iiQslWG0nTbQup6mOYdvm9r2zB
9WZf2JLyHD/Nx4imjiS+gsp1pND3nlOSvVgX4PiE29nbpK7aKB5mVcy7ZULXwrPzm6nAIRSFQNpy
ZhzcefWWbRG/MO33R3hJ6JVWBHND/uTehWF7XaA/E7qVe1Anb/XsV30Sv0ZHSaPSuoJ1GfRy6jlv
sHR32LTmBwg1lR57FOX7VJCAitbfKcy1+mMrckaBw6EaAbgmXzp26dX227hO8NW11TaTEoGKJPu0
bdt4d9/ifJWtagMDGxqbIE9zk8gAV+bG7U9NrRH0ICB2AQEwEixqx+X7e2C8QIiH2qiBtbqs8HlY
XJiqs1tCponEJyIXu7Cs0auDBy6Fk3K6wYhEjVCjJEXdFu6EP9Fmfl8nFoWzz1IqrCTUl5pQcW1x
zMPMct8M5rDN1c3O7aTTdugVAcJeMZ3WSnMrmdMe6XBFWsAALhhgfPja4vPNndc93s/aCDpwAsH2
q5AqFWZmTueKvFw2DJVvZD61ZlmUcq3kHRdgZXotqoEBYOgk4+wBMMwkPb71ycTksuAcGM4zIC/c
SZXuohXkolAIgigCYtpZ/sXiJtINmG1zDL2I6l/uMK5yeE5srnrDEQjD+WVxQ6/YCjY3qKjoVVGw
w9YrJgRolOxKVrQhoHMHYGiKjYghQb40LD8VV/6plDPdxPatvMSQcfxWdmJTbh2v73pDwvbdcDg4
puJr1lIUNKuda2dKTQ7+LEI0xaqMXwCb/IRqFUIOd95KLEIWaPGjMz4Tjg+H6G0n1UHej2jHQtjE
fVgnQqUC/oDdDldKkkr5zXZU6Ah+mM6DaX7N31pslOhVHVeajL2vNU6KMgd9M0gpiCuu/8fHcN4T
4k6kh4I69IXs/a/7MAvlACwpNx2eFbAlHIrJPaq5q+y9Xu8FMNps3gC7vbcXArhrU37jXXt7gfO5
ipMNkB3ED5kWfz6bwJJfRZYnPS8NrAkSgSr+kAjdzWKHV8E1nJmlbg0R1d+CeAcbduWJFnAUNKec
sYoYXNEobJ640tiuP3EMgq8U7kd377xPlTIvbrEqlJYd1uNpX0VVI0Vw464dpuuVlfVTB2YrsnKC
rSvscNLEZwlLTUakSlxoSIPqlCv2E1v4nMlGk8zhC3/cfwB7e3fRNBvNp6KGAIWxwHIYptX66USh
lX44EfECWFqBXahEhhTHX4qZZXhCzyavXATQRwiYqZ4u5eFRCLOEX3JNDTajgp7yEH9xXZ75pU4Z
fuoEsITzRv5PkK8CT7NaK0Z+LbAzdOs6cP3jumGP7H0zKR1+fQNsDPqAO5A9h4ClxYmqH66RTPBz
qQi3fDR9N55n1mDgq+HWpv2sE5RQzWz11JqJ1CX4v4ctywDxKKc/rQUqmOGbLDLmJ+OAONmGWNDA
W3OWfyXrIyrHsXBi4XOCg4/aw2T4iX7hKX7ln5MwDvcNt325UemRquUHU7EjPsGL4qCsit9I4kkp
D6nT+CxYzVeq5s2gYOm0UmqvSc3Qcu0fksDRD/IJk1oE6gFRR1AMhQiPcHGNGKUJts5EGV5nY8J0
P6gGQjzuEg5WavCkzl0R25Pu73pyn0LtA4yCEQXbgyMhFeGMaif/YSRPmUKLKt7+pNBI4sOEnAcU
wsDRts2sWw6Nku9X5Do3lXghlg6zmnyDwLt6PB5YzOpHf/E21V3XG3oQaLvckIoWLyTKUFHOVdLx
jNVi3cx0rAuAu9wq48a0VvHyOTckuA94+Xil/Ags3w65YlIcVC7Dpdr4+5BSaxQE8Ku2aPj+9mzW
Lf8av/uIU5kPsslBra7gpIGFGrsIxglozI4j31C4MAgfW0uJFwueaHbRA7sosseMvxndPK7BhokC
2brsgkMgBi1NmKT+vDEcEkigkF072xr8Wb9oZi6iiGQhQbKIi5GSFsbsZaat3PDv0Jyo1MZM4jnh
tDYODJ0TCpiZpqOwNF4XSDW88/kMdrDFYztS51yem1DowiklrSl+Gg7tGRAC/YaH44iULjjNcFf2
tS2QtJrGE81f7Wj6vdsuYRxzqurw6jL03tZgl1qXyRPp3XGnOPU2xhfdgmNetNsFuskVOcMfYzZp
hrws/xc8hCrqMdl4tBtVu7xFK3dczqGPwRetU7HHRAUT0DMdRayB7FyKbpknwFmve5AM7vXBhDuu
p7EpcLTYsjsif6pRTO4e61nOj3N2eGLoQGRsFzEARE4k9XBX/jd2NTCntSuLhqAGH88q5NTwPX5x
BhIeAyIxgkFTfXcaZVXFUjBhtjvmcjN3oqvwBaPFe6DvTq5F4t35mMlePLp0fuGrcpWnzBcsbI4Y
s4R2KRHj9HQ5koS+Xle1AY+KG1DMTkVKtGBSWbE5JM8aAcpCy9+PikLV6tm9JDqkBH8HviPAFUY+
qmy+aYEG7phnE0nKM2thNTbo9O0xoZUIVw6TUq1eJ5FLIEXnV4i7StMIa50Sojwr8H/PIPpWkBQp
rks+TWckB0zbgLNaPDS6cm2jNOxZlptR935eOvWMgpkQrPF5thomfTcgQt/enZ6MUsjZDbmTJaEL
AU1ohSuIjGhDkxmO5sKy5o6yPIsPaJUzYqF9AcJj9qufIduZpItYgP3NY+sCglmVv1c19w6IeamH
RkxiONWDklz2HibqU3PHgVnycKcRezI305QdJWkgioS4qI8jzpCmPiSji86ptiXrhYsLz7jBbnEH
R+XI1h/lIoj5DXjnl8jXDvXybtwKozCDdRVJlMYgo8FvQ+BpKRxHOy1snTuapqrDafZzoU1VPYS2
oFdTBcgBg8ba7QOvqnrTH/KwyilmJbGZlsfK1WE4JoaJWx+Gz8kHHWtO7OG08D6Jvcmr+mK9mvH3
tFJowwo3YUG6GuA4NiJGvviU9er9/mbM+rgPhMop5gea+gY6667niWmCZVaF3M+tvDmBC6Lkfi1B
JHdPr/s94NwvvHf10iXi58b3VsNQQ/reTa7/PNKpH3bVadRpPtZAgjECOucdzTTL3BmfOz9v4LsJ
BWojOFkWaIngIEsgZ2XGcr+mJNVHpfZiRkgm2n91m6nbmw6XsCOKUizvJboFUXrF61CIzK+pRr8W
WZbcwISMNRVsjxkTfxoiIU5lGFUq6Wlm+KyAAEnMyLyJqdAdRleqZR1m1tmdH8iF7pMJxzlFh4uk
BQnKgfXw7LkmF4CbafgrYq26h+VAZto6cpWQwRXnpnfaD4RAz3ULoWavsPq3NGJ7w27iDsHPzGl6
t/eFMyvBted5UUiRwZCz2O2Bw/ZaLu3kdiboG10kce+/ozcwnsMDxQSyCpbbvEfYmNaI61F1xeFs
WyUj7bOO0vDqwiP3Y+9g6bz+fGCBNoDQWEocTE15ExONcM9TvI692yr9EPk8nNDDLoe/5Mg//jEv
IeS4ycLw/bO39IQzqR3RwVaMo75cdIHpz4hPD6yIcW7f3S+DjvT6CnAqnu885CTsBR5PBdOAAX8d
icgAFoxqyjZvEAGs5UjkdvsiHVc77ZZNdhVxFe3Wkt6FU814
`protect end_protected
