`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
UOhJhdM5wnIGdwj7bnFQ6bY3hCpjv/Zk/+sH7+6R//zhAu53HCsQbHOZSrO3q/J2IoNWb9Ul/d+O
AibRJ/SU4ZXgCiCJE93TOttXsq+n9aYrZakViyfr2VCeYVI/HHoLQs/GAth+Ken7mNBcdCg1mYvo
7ZhP+8mQxNlA42ij8ngoYbo9+GuNAADSzPh7vScBi/iLPRnB6zlslSHaWgYO3TJtr77Y7YyP97bT
4QFNcteYFiUCIE5d8YRRDNm4cMekVBslwMtzYY5o+Ek11S8KFi74w23jF1+H9IxPqTEXOk7WrH7l
1wTFV/odi2TFpBEPGcTAb6IPis1foymexXNrfg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="ffIDfY78oWxrTLnh/vhAZvpX2letwY3zpT2+e2WgwOU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37488)
`protect data_block
J5cb//z7MjAhGXHMTPb9AaBQhtI0AjsWs+DjBgoxFuE5ZAiingUw1kPVVJXQMcNSCDxA+aSKO7MW
lCgFHVUMfIAP/bT8RU9HYgPfeWrt5GTEO03sUGlt0d4LGec3JVdlGwbBIccNaROnWmY1pSxdOwpL
CWVZrxOFDJY0mYzmzwf310lDNUGCpPgQMq+jZVkPI6Lywk38CR1qiie7bXBvoyJsIZEAkRjEKgaQ
uhfLtHj2DYsH7BMaVJWwhSxBFTo4dIBjpyA/uU2duEuhoDWQZaTdF66vtOHNdqvrI2wvpEiHKNLN
wINsCmMKzFxZt2AQUXhQTC6LLaB/DrZccqdNlfwFbN6N+k+EfEpRU/m8wPbVdPrN+WbqfQ/67g+T
EI+LGTUAlND6Ekbk1lpYBkKWHeLfrjhfCxZtb7nUiFBKlKFy7g6HeI+SgehtExp4pT0d8qP35iFd
SqHUoIyUYL2GvPZH3I6y7ZFE/eIJre3OTEMY8oF1l3KNd0p1si3H+h6vr70R0vnqmsmGYhH4XCKr
f7iwcjgUtEeHZIUQZRsK1NGVuJtKH8LOeXua7A2Xc9neqo0fkgNyyvQEzelDO4FQ+KL75Zb3N5EJ
tbObtNMPfkfUZzfXj7IigaBJoBHrRbEPlpcm8sgm0WERKNMQMv6pV35B8vxe3DZUKqBAbtXYPAiv
kpOk50RB+7hcFetkbJys1d1x4sj/M9xR0rvLa2dZDlG3cQRRJkz+3zXUFv02DZn/SZX2/oSHcgoF
cbMjdzOKFRIH73g0u5L36jntWeRKy4ILXti+CenxQGjsFRPH/Lrf2KNq3O77kb6x0ZMSsXrdX0t6
PMUSqzW9oD8aIfcCAMJnIC0gD+oGwjDWQi0TXJe09PvWg8RI/YDYVErDRYPbrZ5O5vB8+fKMkFSi
Z2IziIadpwSU1OGpjtPOQ2OwGYIzlcqtAHuQiOfNH7xqBBDnfP2USUDTNnQulyhxlurIvenOrY3v
M9zUC5FaBwwCrgKKZRczE8cV4HULX3iSUJTGAGE1uBg/WinUNRpPtUpjC1jgEAWHvMzxkWaR8xsH
Ku0v/6WSHKirhnNAHJtRgkthVK1TBZA1MvryepkeKCh70mx6sKYvnyZdkLHP2T0uJt6N3bu2Iqfv
XALQEVH8x1My5+eYlyzL2PJwJZQYrkOa2+9WyDup950bUe7c7aUGk/7Kt+D8LRPt7pBTlol979R2
nEboCx4vPKkoYcz3cLTynKupqV3MOR4vqnYqNrMlovhgTtII5SV8nhSUlTt6ogyx2jBdXCinQ3sq
WpkHI0NfbxSbT7GUFFNGaEX5cfwAfkxbZJI7rXD3hm2ZKQpngDuw0eMlVuXKFfKGbWJVNgEz/PmK
vNpXugPkT93BotV9uqq+rUaNy1A/Eer9fTOOv1JZtCFSPsF3LfHuawsDANLPSGV53WIiBBU9f6Nr
kus1Q5vfiqg/WvX3DXQosylbA6OanJpW6agiMjQ0yimqjwoR6hbGvhbRALtvR3uJKaoMJmnr2cdw
3xxoz0WCnhWbcBdELLulmoAyhQ8gVPADVi8MLvs9hfW4gr1oS6ayR0f8PNuowkHNiBU8iarp+w4J
y4V0zHDfChPjpp/QfxZP4W1NhMi5JYzR7tL11P9F2AS+mGtz8608C5Bt4m3Mf1uM65z2Hr6ftsS/
NbioOFxzwXBaVKZmLhIHO7ZMP03nWWXaxLqt6QmgMIOpkWbpgHCZOPrkiXdHmdYqM+K8RuYVOImR
OTXAMlalJj8TeITRQopPTVf1tqew7dZ/WUmiJkqnzSyJLLemEGYF/A0T4G8iW+/ZxxhK4BkkRVYz
6cOGDT5KjLp3DEp0YkV1Ieyh/gRHx0imXSZ4llJXaj8gs6UwumLXADwSSdl1EmOpHUDLi4zU5A8S
LnkIg5kC9G0cdMM61xASceBVovUNU8A2vBwsTc+N0g1XDbHZ1yywmSRh1vsANk1jfleXnnpdFJJu
djM1o5VRQ7C3V19/XvDjZzn+Zm+nG1fxe72whJHQJnCG/sdiWIcWM14YybJ+LMsIGTVP/u+BXjA3
oML2zclMJssRIJTlvt0EY8069vtQTqT14sp5QQf5b/px9RZ7zbjhk5g72VcN3axVPOh5s7OFLtfT
8UIMkkK+mA/sYr8byqPrDXfkhz5W8WORPXJAgrvlHNITA3xbMZ7bwCZL3DyjfjXUcqSCJHAk85kz
V6uvB2CYFhLBGD3MNPJzWIVUqaLHFUWMDfdjeA1tn/2EnhMzh+bDVLV9DxppcMwsCKaiXFHxvZDl
Qh4EAEcfM88Abvyp+6Tk0EGONUnDZlsMARZ8zPnqVjE36kV+S9hkxLdO3amThG9Y7FZVDwtVFsXN
CDtUrAIIkDv/2BWfd2ezBYkLQigDB9b27+W1UaygHnXWACi9ru+jR3gLGo17JXK6WBTdWR7NOFe7
51BykGlrapEigpwgKCP/Rc6MjhcNMf77SPVLZHbf6wR5ZOc8uGzt9WJSrONU8fUnbgLBgapJz7SR
q49SF50/1fGjNDVMgJQeVecnfHbIkDGvvX0eZAxLL+zAi/K9Y4hWm0OBTG6khISYzhUBjP/yl0hQ
Z/9X021CcSu2fIfGdB+WlxQdPjhj0y/rgsyZruIktMWugnZoPQAWWehbniZiGrdav2BA/0cvRfrR
wa0WP1kZbPQMxPM+nhmcZxv2Gs/Hqr/ugbmeZWTO3GGdXhLKk4S7m0I4YaVe+Bk5zPu+8Jb1HP9g
s115hKEuG6mykiCHZKouVqEzYMTSMDy8gElXrooLiAwjsy1EjI52q+A/oYEoyPTEuYwtfJ88NY55
I6gTth24PlU+giuzrG8AeV+Ys41jjZJ0Sefhvdipu2DsGKBCAMV14VH5sGzAdjVdOMkyObD6dsuY
40U7XeNtI4AslfcjO6XhGvRKNlgsMDeQn4/uiBmXoTmGmebRs3TJFZFMFbWk/+IpgpaB0ZdJj0Y2
iYLIfddRs5JnE6hwws0f1iKjrikur/XN3jVpNt2zQ2NsS1Pj+ZGhhmYi2Xg6wIrW5f/NoF0qZhmy
LqH7VhWtix1UUwX/BWYXyMCwKItrBs1vZ0hVcCTJOSR1AXPo6zVAxw9kBRnNYu6P1I8yTUQw5lGn
eogjFKw7Rn4YOK6xprtQqduR8VrEkG9WJHXqX/O9EHP2AAHympxefDDnI+zrxpKi4Lb3N7z6iC4I
+WPJ+K2QGVyIsbxoBYmFZPG3sKyhtuTLO+l0n70zqopsdqrEUbKzgStPOBf2VooHdh7iE6zAjlOo
+UJwLUKdYaOi+0/mpTzwRPFQVrCQOQKZFYQcZ2kle2y4+a9/AokB4dJwthBUHemVr71AceKztmTD
/nm/FXXmaoLENDgYH+qQtLoIeX6NhWJzkbHQxc3zsTZttZBoxaed7+6OF62wsIDri0XW6/GrtnUh
PCMDjFpjvs/cfvhX55Pg/pr3Io6CiMEN63vj8YgsBfm/YHXMP/xr+61R9nIRW7M+2hvaYdmfPZTP
2io2XdmRr/5z7N0stqJrEYvvNrheWKlVcPx3hz9voLQRm4diOXcE+v7jIHNzuNBUVXsfGZ7sWTlY
xxg7LRlOKyl3X4RZo4ueSJLgMk8SQfp1GPVojYUAGsswWOCAkHEuxiTcPp1hYG9kz+B8HhgwNsTg
DCI6vA8ojxYrkCV87unB3ytaHQOpIMUOUl+o8qi2qfXkDFl6r8pg5+RGvREsFU2xO+bUo3k5KGl4
JWhfif35HWM6npGdk1v6APgfW55Cmf4kY5WrJK7p+4ttu44+oq1jRNtRUYn7ThvtI4MwWT/2eF8p
GcFd0/8YpqsIy3zLkqpPxMzB1JxRQDwHnj8x2tvJa97nsIZKmn7ncEJ3fW7+9VhRegsDQyDKIF2l
C+FKB3x1ffcwEaHZMUTpTtNu/dioBp7q8EDeSFUA6BUwRYX8fyWW8VxHeSjAnfT97EWii4Iyl9Qo
PMogTH8WMcEpQ55rrTr3IQuZ0U1FDeC1AGPjiAH/DCYGLDrQ0//eoWfWYamC1JMfm6j/LhVFR+HZ
A9HS9gcMAV5VM5Rkpw4KIq/ADQM/CqBpy8VyrEQ07LJMDayoF6yclZigHdzCwRMzGArLMDMDwdBR
62orMHVAI7eDBwpbKE7t+FfqbIsJcoNUS6Zm4TPjRpbXUHcbaRSzXtjO8/Y4yJq2/Lprje2d1oxq
81yVSEKi34HiUhbmBs86dZbZQBSj6Of9WNCO5NQHOj5+Lo9hxYqqFKv2H29bdhdDwjFIWnxD2bvO
Kl4A++FKxPCc80WIC8GD2LmsWTRfoWPPV2GxYxo1lO1NFeZyskqifjPbePj2VcaE5FUUWHebrCTq
Zht7msakw918HitvX5uRsBzHPzdQ8cYfzpsY0cFhLH0sQmp3UHx8vnNY7f3sU7f9o6X50g9z20yq
edvx2tl9+tT0Xh+QaE4p/pR5z8Hknmyd5jwVblpk5Nlh7qHOMMWCeqjMrX9sk3DrBFFDUTk3qeUw
vYvmY5Rqxc8WkOmf+UxD4/BeeDlu8h6ps1sgCHZo5Fg77ynLwpBJaTxk0nx8e1nadkdK3tsqZa0m
ZrKzZ8jI9SUg7oNo+pZU/R3gI61QKHvwAwtUlNBEk36wG6ZiF2RjbCwwerY5lIDQCH+grkjwCZ4z
+XghAcAsL5450TGEhy3eMaAzoP/BENtrDuYdvaSKUNQ0G1pys9WJKiBXfsmUNwD2NRRbaTXmQI4y
RgrW9/whxH8dkv7p+Ns2k1QT4OiYtop7LFa+M53w5O0q6dUCAfX6V+kJCms3aC0h6hzzJ6VE+R9C
dgWKCZVIgqiqJNKPhd24mRbRxid4epruSDWPfAbnTYFk7QQvr69p4TnIn7YdR86zMcHslcrRlpyt
B9UakKCv4s48kuTzfweeNgXwHe/bW8x46nrPrxYP8r9melC+n1j2uDLkJ8wDO7xi0sfSZBiMDZTn
eRGfya0+B37Kqj9lcgXJaIkFJ4/zfVooBiksA0B75Tl2U3JQ4wuVCiTbNcD41ur/MoN3LDa9hns0
moQoW5WfdLJ8NXlU33Fw+QmilDGojaSUoE7culMkk4R/NDMoZ8gERe3Qyi2fuLJUsyn0vMQAnQsc
8VGelhrDrBnawAAF4bEHWU3cs79bPVJM9wZCzD+4h3tukRbBgI2p8PH49D7BCVh2hMZKq2TVdAAR
8A5goLyVt7/l1VdTO9zq7yQYIStLn1H8l4O9bGpkbhTk0A80S08Mgz/bhiagPv7VmfhCQZ6OA/RF
gHUa10eyvh7RhRKhb1nNACQFOoVK06XbfriJgziADpsONGXwDPBisaCMr8I+TQzk7VlGdMUYhabN
a1g374OctM2OcBclyGiZZVY7ZcWKr+AFuNs2R3lDTPkn+XrO8H9KsmhEi4rzajJpYaL+SeDrK9nr
32zQONtdvBzPsWggcBbpqE5IgZmB03I3+ZxaTpFy5EDVYuvUA4tGZaqU7k0u/8WyBRW/wSSL66vY
Z8ZStwOVTkUbW5n8+yHjwqe7Z3onltUumzgJTTVs+gPdT5cHD2aue1nKbIyan8VK12ABG9qjfF/W
eqdgXs6wjZ3az2jzfs04nih4SBSRI9N57y72iBwNMaTWddtrUCvVvFanpTDx7e/xZQFR0C9GFYIB
9kJr7mk8IfjnJuZYSEU7FZGbZ/O+pMxuCRfu9ec1BmM25RE3SXYnoyDdlsZ5rr6fwXbZIehOmimF
jHXioRNQlupuQOMK960jXkhw7dQ5Cu7cEA/JnhrXF5Voz2DgwbgrcHnPEFuMDs2gnOR/BIibMkZO
XqbAX6qPGSe1lLWIL+W2+2N9AAavNcaCu+ehimEuiMKAAaHjpqltzdmrlwpnV0hApAl2vJhslbGg
OyhzUxiE1MsHcoRWWss+BfWAfI/edwfOXFhZ2T5E/HXBGVoeow9n0JcAf8ks00btWVOCBYEEBywT
vYn7a/wJioff1ViU1btKmpiaqWgkbVp/P/9iGZYGKMdnZ3F2q4UNmWk5fJ14jpajBURagycrkjMJ
p4mIUjK5h5IRKnKJgGIgmW6h9gA7eCmVCTYCYBN9yum5rj/H2GuLFsDtZF83BTJmKRwjTuWG9yNw
Xrmz3U8b6n7b2OzbNdi4mm3/TRjc7kyqfMzog6A1EDtoPwjnMPdzGdm0WRtj3JtmG/aSEA0fzDtj
ZghFsTH6PJuY75YR4ia/K7hRrFZnEdymoxt1Qj/Fv5gdPT6txJdHcgYI7Z+fXgcEU5I63QoThBJk
kzbkgYnyiiJAusBA//Ry9GMDfl3oxbmrFrZsIyMcZLJ/RjUYQRXxJETBz2edX6UE7I09aUN7ynud
IIQoPPqdSrsAcSbT6WlJZbfX8L5AXWgjeAJo9neZZKZNQk+YDC3zX+YxHs4k61bXcTTgHgxwCkRD
eDtuWe0MJIZssf3g5Z7DXF16y26gZz0voXf7+EOXxXlJFvDSWDlgV+2kwQJVZivLjHZshS8VFNy7
qVbJLPvbpiO1Mw+1NnYvax7cA5LhXkSmTmP+P7rUuUK+r6aJIQ6nzWlxkrD0g7oLZrQulfG2iEo3
jZqx37VoXaiJ4K6gPYDmgWucwc7hLYjZdW7UuzS9ZZRrMgpB2U04aeIg3cJTljgFAo9PE+USais7
R3bS2fF+f55IacCNNgq+qIZcPKVjleqWzISAhWLQ2ABvW3Vyd0pvXOtqh3o9aoCR36bF6krWDi8a
aeuN3eD6nO882yQg2QUitmUxY6pDmYkbMVWidOTuaYHV7pXpv6qRgtTnKxa4+AtmYyS+s18kJPqx
c8WsudZhYBR0XMjbMpnYJ3bcJM6d3SoyxAWHN/9OW/LXmp2yXXlyWZ/QFljBPd6FmXxH2Qg6M7B1
KF+co6WxA2U1acV7bckQSRzOo4nBXdQS144S578WlBnNhbPrXPtKRFj/15D197SCmD/VJd0ab3xA
1NCAi/59xEoLX528eSnMjWPyYU82tTjUnUiKFILLpmpgDOs25puozQmb4AORPPfoNk+tzuP5MGxl
U/3tqwlW1tb6R8jjDlcpe9J5Ybs88kbh3U49IcjaZrU+FkxdUXZeX/diKFaHhtc8pWNJzt8QULi0
zz7W9Zh6bQ/0Q8HmHVPa4aZ2y4CkHFL1sa0aPfMw0rwndV7PMSun404uikzVW9VXEy0UQro5Ltjy
CTm2/HecWnarhG8m7wmnzkzpDiFTnbzu+KlLVZYkT7bNsr2g9UnI7tNiicE0Q+BIz07plQltysoK
psI9YsAlaeEHaSlN0nsUSRq5Y5ws8HActme1yftdNpFXM9wrNC6w1SG8aCjetGH31YkcCfQi1xOm
fubrRi5fHtgQastdumpTj6qOEf2Sw3ii1VGtC63wvikBgW54pt/6GvX4l16UWfjq2/3yFH6019hA
v8mYZqtOf9WMjg0tJsVjP5yZMX6V/duueIt1BigDhrIMyCkLbBmGJMR3Bb4Wqh4hN4nyqe8+d9iE
ZIXQ34fpBezPslp1ptzLAz0arvrIVvImYbxTMqH4ogz6dLpWEP2RIw1RuI57aQGPeDCV8msYrvoV
YBtULhM60dzCj8H7S5NPPvcwNMOPAXERyY2eb8tdiAYO9shf2wUvRa0aF91dGsyR6xcNPPbmgJb/
jxCE59WdFMGIhTjyf4+Pdpt8Nd/HkK8GYAmVEQhf6RDh6i4Iku9gMtrtYL2RR0EQMLls3uxev/h6
S+TGxiTaJyr68HiJN67DTXncgUxhX1bJHDFF5tTxKGyTpNjTSsriWix3qXlPybGnNAf+dyg9mKgL
CDg/a7MTF3QgRj2xsWP2P+XOOrrIWCw6jktQt18rtcNGvKRGp9680eUe4rXYdeOq242vSi7kg4eP
Vav17/kd9TSXojbjph/+FIVC7q8m4zxy02o8ddfxrHLZuI0CFSmr9y7Vvvyp4siGGldRS7ghH1XN
6zhuMYuTqHjp3p2/BnCsDeyG/JN/kYwLIMelXeBtxI/mwhirqTzyowbK5cRBk2XBg9HO/PQcMRRF
GW3yP4XsWTTeeXRBl8CdF3U1a17jBjHAdA65XaLdbaMf3uRSDv6a4abRMgiH6F4dlWDxpfj16MKA
CC9jTjn4qbEPzjp62Jg016vY8z3u4LIcFbvOIAk2DcVWQSbPobARoj790OuhCy8ZDZes/S736psH
WFXHgi8PjzMnC/p+YrqnvZAsb57BZ/G4zNHeOBHigjzYGGzBUb27FT57P7lBUctSiC8piHikCv3A
ORNw0g2re9B6TK3T7ak8zNMJ50NLl/anTzh58YaNpD2hz004Zmz0jNpPbOm1ybcjkFr92+xBudfD
CWBHoUsljS4UD2f1LlCNNh+BxkCxZUvfzuf5Yn8kaARsppTYWvtVjbI5lzceocuYqSs5e9S6bYlR
WpzBL+FD4OEO2HxiJKYJIOssRD/brXngpyUWo0Tg+XCIhcpSChg4eCkXf7MEMIeV9ALY6Bhj6H3l
dN3p8YYWhJRT/WrtJ4KaCWmJM0psryT8KLENATfNlxVO6OAbSCqF5AforEbevZTHdultOfmZVlRo
7QiE+CaWz7zzLqiTjFarx8wFBpRSGVT1M+mxWU5KYbZ2ihur+tTUBrEaNI+JiAVi/F/LSp6vN2Pa
hY6DImsmuZujkrl8EhiST6dd0iMpyN3SAx1kpmgB0boZdNgejnMvhKMerlPLzbNlelUC8aINOW6L
MZkJ38nzBBprUafCJ2XpIDrhsp55Fhh7bEtbg0sUuTDTGW6p1R/jQbPZ1TG7psZwyKITnJyN6dQU
RwcvGz1L5Qv0UC5ply8Y0KgdNLfdE36NIWKRfDCm/zAjj/nJEoOVcaQXLc8PHT9nSeKP4Sj46m/Y
S7KDJl01n48Liw2JJVXuu7affBK4PfJWtvKmgd92rjHJFHewy5HuSfCN52mXjDcbBIff33oXsgkP
CwX+fhIjiOzm5ZdCemyuALLP/cN4mbh3T8vkfy9FLsYeBVQd8ZuaJRS6Z5HBmhfWvQALfUfIBQle
MM+GVIQ9UY7sqAlVTDM22bTH8PwKe4FizVWpxvZwgT5UQr3/ir/CDJuCA4AJ1C+buVE0By8eWJta
pMK7+iq1HewnUiBoBZDXdf6EKh362PBBhtQL1g7xo2feHqoFhDrTkuanRcrgGoYrT7XcnM9ZIeS7
MHva6DmWlU8huyRv1CIE9pf/bpEfQDNNlyITafQodkrqCRfzRtXXoKLPQYIO+nyMj59Nwwwmi5M8
Tgd9CtG1Xmo0CGdyjmkkJP2h4wNa2zhOX2K7o5L37aBRkLvoa9jfz5whaNqYRMisK3rNueTxa/bo
tId7tLyy6NI/ANlNbK5ljFyR+mXiKvBp8bJUe8cXhnsfhpDzJ3748aqy8WOjypVy7gb4970pvM9I
BHGImHuSm1ajvTtpP0UpvXeyAE0Yu8uWSJifqbMyWKrBdWaq/4j9lrGM1AJ7HuCbkNN2x/7P/kNP
vIGISfbSUDVEemOtuRgoq072BpbLJ3KlfFT+bDrAxLe7i/X4V9qKW+NgxoxRKRqpg5SWmFCYGIyg
ZoLOHkNFv/tM0Vg0ZGnsbZyGzOI0ZtXzDlFP5MFTOCmOIaFjQJJi1EicwkSDjIxjneG8l0SRG2pC
k0JrODGKnSJdDNnQ9nk3P93fUkFJf8tpzh6dobjKxxDUFfzSYvcNHkAoZp6o0S5Wjk0Ik9yNSqXR
S0iY45THx0yBxcKn8PVJVbqN/GDl95tN5+zfdJZJ9mxxMqYjnv3r+Jw2Ope4GltN3sFNquD2Hiav
aCYKBa10+Ps5o0gxDwBBhy7Zoy1sJ0F5UOXaTg+eCjTKpH6ghFZQw2G1TIoO479LkvFjw+ZT2yf4
Rxo7dGktt5E/STQ+Svq6gZYkwIzf/UDr0l02SqiXoYuMwxg1J3jLE9elLbqCs8D6pbm0N8DJ5XzV
aXiVZy/Zg7gVUB+6EryvJA2DmHYp8CY0ix0d3lcPgEP6u5jhcYiUB1VJHkI+43DKwqP/jNCgfrBU
/L4Eej+7qItxq9ZHVfS/qvx6sMEOfQc3nPboE0xdde/Sg6cb/VhCAzAA+zvUTJNmjx3Wm12P/b84
zvC+Txstecytsy1NEVzmaIm9ROof6DGxchZnMfirTKdGPLrV9PB4DrH899SDBNXRPtLCNZ6duo7C
eXzS2qN+I5RPdW2tiTwdboDKnb77WeLtDTrcCQdWd4FazGFI/+4dg61St8fN2aj0hCn5Qk6xb2ki
jkzWJ5D/C+p+27jFDPf1Z89PwCabZSP5jLTZN3lEhuo5DQ9GmYbXDyL3IURiEkibTMjnHgswyASO
00CvxA6l11UvxSKYUb6XqL/tapknxNT1LQpuY/gVFKUqe4d9h6PPQG9KsZ8JVahe3eRoncWTPcnu
qaSn6go2ILaEiXn2GkSbM1idj4dpCU8g1awMj9Ken4E7EVp/6ZRR8sae+9mvT1ZYGcRalPM1eGYE
aEVgfU98P5MeZzdDa+8Br6Z+dy3yf30Q9PmV0UDO5Gjje8CZeG8NRq06e+XPuXyDJaP9nNYJz9eT
Z5L8Js7nzAuvq1qIP0m+vTbHV4xMRFryvv7zY1izAdfCszLlyEDFG0m6NTN2m0Tn8uSO3V8zb0Ns
HrZz+q6BljKq9nRJmDtnueiySiKXFrwXhByqkszvHJ9dhIBlQwNA3LfOuIufjPcYVoYM/cJmJ8x+
yl44yQDrbudmdNPWzMS5kW0GjRUKyCqZCObk0ZYeVWHVThdTLuH2ZVcykLEoqVD2xzSmn58soqa/
+DuEUpe1hwt6evdGf8BlpwSy/3Xo9tVmq/pqYTInKObjHeHKSqsU153c0zCV1bi1uXqn9TK1EKtD
FbbNPMvKr57+4WDpaxCnB/0AqwxK/oWuqUu5bXrZFLkNT1MKw1cjp7MalpvK+D4UeQMnv749iPGr
jTW5o14JhVjNCtN0zUrDZGkJXaEEg5/36mBNDNAQ3HIGUvXgxp44aJRKmhedWkS2KkPko+SQgDic
CX4i2VAnFqgPlCRrF5sMqavZfbqP82+9c06eVSE07eoEdwA/WSj3Zk1EiWMmIkDA+A8OrFAQNvgT
PeoLbwrRIdqqgOg1qML+mNAFuHNNoprERzYAEVZyPBv5wtxtu8h7LKVdA4TRSieRK0hkc/rKgvQY
bc1CgIGGuOYt6pTlF+uLTCS1DP3EYj8WioXi0NDhrtAO8ZW16tej+jITudvF5tE/ziarg+MrsUO1
AZ2kYIzK0OemUttgPPaaK0NCJE6YSfo92TqSzsNYwo2N4ImOOjLtJFeKQ48pq4uujbD7cWDKnQdm
l/ku21hYYUmCakSOceNoNQBLPip55nS9zsiVXtrCFlc1vPcIHRJkbUnJN4ddR1M3Efpj9BSSX4S/
zIXJhn2Hv0MoDWA4XvUkKtxRKoHdgsNm7ubiEejYO3twR5OhHvQGprLvhd3x7H4+Bh/+ynL1wC73
YNGXC+gLoAnp1yiRxSSvQRRfazsE8QgNJ/Tygy1gLuikdOJBVfDBSUZXTnuaO45AQeUstroOyaEb
gC1029E3y1jdn+Fji+yFCD0x8D4ih4/1D27D5yAtF0SQx1TTJBvl2ZHBBZ6fYWg7oz6AXDKSiMI4
U05POLcHsObkxDpQkPnrszIM5laHPEeBqa7/eVB+00FCeBfS3T530b7aYdROd4DJ4Rv+5Rq2X1dd
qQdgeI1cROCNK7EawZKL2iTD5TNN5JFCQVbQsWMhGxtyOlUwMuhSbhCRS6IBklBtdpZckdp9X2Kw
0+4dFip2GRw4WVUpd8WojK06hJ3CKtdOWEaTCBnKBb6YWxTsBErAcQARYFEX4CFiM2MDUnNxM0/e
5QO+pdAWtqqjC/JN3S+ziXgrDTaKiOGB6svoYS+bQ0CE2Ei1HHmRKRdg0th6BaVnmmur1c2qofLX
AKxj41e3KfNvu9oNFGhGiN2fLZpzoK0uAb8ZeMdJw1B/DFabqTNsxtUS7PuxqZr2AvMkoYy3QGY6
khulcq0dNoqmJGyByz6eSZsaeML423gD3wCd3TCiGsBdPGU4bhuN6AnFM3/Ua2OWCHgeNWjxnFMc
qmfxsS1amnhs2BeNK2o8pxLjyWpUMjYewPK5ztoA9CzQrorgzuqCMf2Yz/7J7iV8cxXrm67JPTLx
5V/jSpgEgMHfWZQLfHkgF+46ZP0xU2GRd1n+hy5l394qKuy54mkZIWhr8XZSgpppg6SSN/8OyU4G
/A4y4f++3/fPZIBe+EsNJK+rFolHx/Dvq841NIFI726Ec0yTbzSEQoDf57hh6TTA0rb6+k9161RI
6dN5B8wc1kFuYK5BFwriQNBsKB8iWmDi9ORBv9xNzHFi342oiIUURdpJClyahhKrdDSRmTfvX5wx
R5JWZWJK/t82ZteLOLItT5XjoN2+JVvNCv0vZVr5i4WfWcU7c0B0IWGkuK/a1LMYtTQsbyYF1zAn
7mtua0JoC3Ok96JPfigWPEo2ObqIki4CLO/FtFIAM8ihPdrZ75mCo/MlpVWdOdfH4vQ9GX2BQX2E
aKTcA0fW2SVJ8oc8PXq0RmfHW1FkxAG8jDOg06MBDC/ucf/hCsEd8yTtqbAwRzgpMeKFo/9FT1mL
fa3FUnKey+TO/yiwXGELmFDeNcKcUo+jJ2STHLnphru04x37LYsYyRfQgkOV0F/RN6aCHxm68RPD
yDBrCRC29hoAB+WNl12Jg83ymqxJxcfhDruCLWypda4dub1lPvRrnkQRrCl4Ob78wQHGW/vy4g9b
TJ0/TM6fVKjrZUszSYsQmT60eI/tzj4c1WTT2gnuqxJNkl/vXNlwmXP/i3zoNyIONsYNqs/CFf0k
gvDCWrmhC3dInVK16plrJLrdOefuPkueeKoePlE6whsMOwg9lAMJCeiv3gRTyf5bb5SI855uC4Js
q7ztWN4C85LR05UaCtBtCU84EQkpbz5nOs3veVuLpgB/0ynVooEdcH4MMvOtoE+3JAzO9L7zqcNu
dSbCfIX1dEPeqO1qqqr5fPomBQFUw9eY97PqAiefy6eoRjVFDWZ4bwQKRJapevem/pSCym3jOkmH
GJi8jeoqet6LuwOMo9P4DjKc0toziTGTbQQKWe7WxBXuhTgfSBejAEXogzcTdjGgsC29QuoQn1ui
chwF6LkaldFa6LWYFO9RZYZnolX0LrqAHvgte93vhq3zN/CMpqg9fRD9psjX0AfsSK3wW9svoAQY
6apdwgmxKynhWQpBD/TXUEps48wPibFQI9AAzULXPYASCrLu4Ax+TiPPT+sE4Nqtj8U3gIDdHWR3
kckcdXZyT97x+5LOvin+s1eRzNOWdCVMYYsEmE6VMgZX/O8CfC6Yob62gx388mofm39ggWS4y9Vf
9vHwx9x3ErUyjo9kn2qCQyS0zNP2CpteJiZiVmUmJSgf9JlkMZpiC/J05JrrZJDd8ps05xVYYCHf
xzNH7kqpRocJGWVle0t0qPagHQLlxXTbN1DyqS47afNxB3vXqROUhzpUq1oJb3rDerb30yRcLRAY
yZDvySK1yR/Dj1Q8GTdKuqVrIyxkpXtBaT8eT8sDgYM2snWVPiC4H8/q1KORAUHGE9egG6P9Adsm
ac4SIYnxmLeaaCoxcuKBzTttPaSRMr7k79fS6n2bRntBmgeXqpNunoUg2Mxj+OvmJgB8pOvSZSt6
aVNtBmxtO1l+WEQlf4iU6US5qOncnNS9963NZvUf202sI+dCZvro8xsnFeXmzHMvt1B8Q3fXnV3g
uApPcJl5IH37mAogxLIYZnh+nLUNvbtalFxoPtaObJJRiZ+QzLVV8IJSXxSaIJhJzWCyNnOFf0pl
YYnX0o2NqczHrUlTNmj1+dAuPh8y5fADi7GyKJo0+Y8XMVS3cSG4skL0YoyyXmMgtGZcX/7nXKpD
reppa46EesbfRvf+bpiAjQgLX6ZtGlBkZg/ZOL/ftMkp7m9eZO1FH9kpdmrkt3g0v1uV5nih5edy
qSXGdFj496PhsCZhcURIvkdgBPMjFDhQnT/z3kjMJ+YznQcKCZkLMloMNZ2jmE/jhSwvmF/gZBL+
Mwt4SDcLTXoCDZb+KOgpRTnkTUShzi3/QlA2BYhwOk7mCPo7DgkJB5sbCZYwLV36mlcaSSS1lZPp
O8PH6XqqQxSvtH6AShdgIeXzVfhci6IWZK0tYi/uiXNlRXX8Ouv747EEW08vgy+fHUC7sPUs+s/G
VC7zv4BR0oeot0h41WpRG1jVb5gL0y1+quIpm4Nd1hjAduVk9RPo9RHcng5cDeTbVi7dqwAfz+nu
XCXvoLXyzYmi1r9DkgD1AN4xuNfTLb4HshkrWYBdrRMbatVnL7eNJFd8SspwzkJzSoOst9kd/AOS
ZdpLVWcP+7ZjDXyqt2Ysvd9jWf3gh5zJl/KlmneIptPRDBRzlNU4TA0IWjFjAQY6DMn9q59S3alv
ACrRsLgLYspHhoMiGwGO9lgfUIkPfBB6dQziM+fy+yBw/uMI7AsEr987izUBHE5zBDcuIih4Z2Ej
irJGe0Zd5laNqlbhb4OWndHk+Run2KVQd48kblG5jJcdcwLF1hbSctCnfd22Qgsr+YNpDE62nkry
la83DLg054wiqbqOcQhhGMsej/tunH3+uVT8frIKufjSc3hscMHMyRT5ByOJ+M+3SciU1utL6tyJ
Mj0/QyiYguDsOuDqs9Y+6u8NoOJa8NkPSRSITlNGCh2zmQNPTC+ElZteVaQ2d/N3m65NVn41bvEv
ThuOEuG84g1KZH5p8w7ydTO3gd/vp7p8uhhZ6KgGUorQDvEGBpqI74VI+LYo7EnkUc+WZYsW4qm+
MDoee/WrC3A9+5tfDyupgqGANH22tKk5uoZjtANKbXnGbxPJqUF+3TvFtCMBsDWAm2VF+u4t1whX
l6U72F1p064XikfaKObsKjLJ41eoi8PM3VudSZbSKh/KoZ2BaXmmall2u45YRhewyME71Ahj8tDt
RPUfYJTZRSfohFoYxRzfhXmkmsHNcUrxG2fDq1Z6DeqkSu8Li9uhvqSzVXAK1/OXPYLRi40oDBpw
8f1Sqn3fnaQkR2xvy3ADoCusCOcaI9RnadiElWW6Z8/EJCbripaKTPYxVsby4spufqC62UuOF/dW
Op+fGOvnqQFZ9lk2tENsNxTyfsSA+7T6F5alFwt6W+39VhEh6Q3lYRLsDv3aZWMF6WDLkfyPq6yI
4PP6mFxoFDAvv9mhjiTrI8TyOEjKYgmm7/Rf4qnZlXhyeiebv6FSWBAo9KjW13Pcix8TqkbnRu1X
S1mXfQtIWac/MbsFUGoaM8AWjQd79YnbjuYFhqE6UTCDjA+3GaWomyI6kr4LRusWbLhaULZ1q18K
ujlQjpsmGbK4feeOEWopO4owbreOqcFBGgSxpWmAWWWQlrGpGvOjHI8ro7b9RicfHLAhHotMwwBt
UUfjJGaqOOdO32K1tO4V7Zh9akE26oKr/R0rrdCl53n8E22gBI+BY1oB0vlL875pSplStR+A08yP
GFHb01+OzxoFlm5Z4lAOfGLFPUV+exoC/aP6Ii4oZyP37/yCeoKdzJ1Dxt5GkqeY7HrsSMspVIre
9di/yLcRYqNYOLVNm1RrexHFdMdeOnxOhIpyyna3gnygBlObq61hvFFV7sAoDABAzqwINFwvvVnX
HaePnWxo1kbzVeodvjIDvI05uTmd7Psu6aFFOe0pCs4rus+9Ud8MJMHufzB8w9/iM861YToidHGe
/PaVJ9PpTaWEuen6VHBO6BaNT8BVFy6ZgyitXOsepWfO2f3vkcR7lDgkcapPde8pZNKCe5ptWu1Q
rSgjwDRpv+OCLRZ+MWPoMIIcFab6NdulOq0TkJ/1uUAShx+FHx4HLo7AxHf2g+ZuPUY8Apy2oqXy
GChjHQODbyoc7Q0HnF5fVr/a0edZOF09e9IIdhtK4pFJ09QCzQo60SjLvkvi0K8ScJjChkrudZh5
If08Z2SmmQsBTvjW8LdQp1nR0SFqOVlQ+R8222NzBNDlHpymh4wi8rfz9RC2eXY4jJRw91N2e60Y
jWwnPvFaiBlSfbkGEwYPhVCluihDFoExdJaPMSBG7xOKaZ61zQkp/tbXAZA+ffuCg5HpXsr03pbo
Ff3pN2NCt9TTykfdYcbCfMVWeYiTOfGv6iQSohDEw06rfd6VwjXaaCbgF6A7RoOVKhZpHjYFh3YF
Sp6wyMdmscaCGExuPJ9mL0K38fcYIMQ1qLlFuUnJQz/9Ig2xPxQgeexX36/SxjQU1hdfDTMFoEje
3dJ9XfY5jR8cm0tjbWTO69b5mBX7qpMWbj25pvDVKv3VR6XHw7HMZ9Byx8FRabjG95+aDZfuCJzF
gpHYNxk0J9ovnN380TWA8mrxNwjFWRxd2W84jzTlUpSITMuZmPtPvMkvcDWuFPtG7xAmtcBQf0XU
2u136/ZVKb2gsnOV3tfLiwfexgh5DHIGdvl4leySZX7YGvcvEB6yPXlGbYhrq/A2Mf8a/CDTuLSV
JzMUwSjbK8aPi9KeTgP1ny9DMK4INvitaOoW1aTQLA5WcIRe4LfkOkF5uAKUKGVgnevNCi0Kt0XS
ciEV8Sl6EJcoF1cX1LI5haZZpzasETyuAgOA1Q7aUE7c9U0sYIc9KLt3pEKr9sAfDmm2AlGhgaXt
Gt3V5n4DrFFCcaThmjXzcjXNUHL09YBMVrZNhROxLKkXXDBIGtAgE1ZE01WvNkYmexAmwl0zJnDz
E/PyE4ot+dul/MT+ZhoX3V4HRxra3WmUVtyHRu8ocGsOjjklFBvo6d3cdaeBuAlp47FUywNDTEEi
lvEN2q0jFoK1tcKD1K4BXLassuOPEP3SETKoFpSrOzdAOJNXnaHNgUUcRC3cYxy3S5OsZDvj8nKZ
2q/kKvKNyqtXGPqHiT9W2YO5xOA7zmxAIk1lt2J5652SZhd2ocwinuC6TVjpAjWUnctwUVlsVLbh
WIgEKgYE/mpoG0xlTVs+h33lVh5MdpLCSrmVxr0/6vbl0uHO9drkQfLmzfQIx0Ofr117Egu+qX6g
7EyKPYW5+Zq4LYe838KA5r75iUMvssWsLkDGpVdTN2DAZ5EnSuiHjgSy2f92oGFU3BkmZwM3us+0
THxTlXfYBn5F0Z9kuNm392I33TM6rnSXRrzyvZbckSD/S+IGzTfooXogKymlNYm/+yvtmPV5reZo
0hhdpesMc/OJqY9Vj5IOlBPi0Kan8RO6LpmAyUqPfMNaKXV6WmBvua3hFrOhbeMdtRscytQb4wER
tBSZuGDl8AFDL5sddQhsLKcfrqPr6Y4xkdOCVKJOPfNJE0ywWW5zr5SHxbWWV/D8s2ypXMtmT/qm
CaFNNck/MH9by4gax4ntQnj0CgAgUDk8+uf1hZyfc2VtpGAi0VLRG3Gu6Lwki1jN2ZzKDO/Dy5Bh
bkd9s7sSBxGu8FRs08PIW2lLs1wiPmnqe8QlWNFRXmOPpkLrbzUTg/Dah7vRlY56BHlk/zQ8HLfk
zR/5sEprLB7Twx0ByenxNPbh47Pjq2avx6TFD5HGJ8892mQRPEcSbCeds68ao/gHr+IKH1Gwil1B
P51qgiZIHS0Pe8yaFcuqYQojVEY6g9jMkyn8WZlxZO3uRXtSsENac4rqWZxnswksq47LZaNGaIUn
UsDdI2EKv4tbFg0a1tl5y+R+YGw/20xBkvLwbzk1bijKoDbe/3KcOZhYve2o3gXIv8tbNxn4Lpj4
3eNdxgkeqGf7NJMCwIxac/6zvbInPG9oaFoVzX97kCL0+i8yjkyboiAqP4mARBjx1fme5X9Ef+zU
0FytqEq5BIsStuj069kanWE16iG7bfDS7e3sXjk6OvaQF9rJ0OpHbk33ghMMsjRjFgVJoKGQsbqF
qFtN2f7IjCYYjC9xGUgykmrvcIkMkaPezLJWYSZCWYsj9eBohvq6R99V0EOctPUGKUJEOLLjqMhk
9rMZ/8RKRg+vk/mRpl3Z1mmaLJHK3YayNROic3KPrcOeuRlarwiGyxgje2WvKkR68Rvkt2kR9opl
YsXAdJVuclimAvurGM+zXQXNHUFfn0EyocvVAoBDq5dexPUFqq8RRUMHP/CJYJuUPHz3sMkHvWN6
2wxmyINs6TIvFvaEUTvPrMDLtiOb1l+gR5ODrFvfuk/np8FNCI0qyvAnwyukYWG8/pagmmb15H8N
RKfPsDt0apHEd43Hl5fR0D8d0Ws/joYSddbFCuHLJQnPz4OJzGszUtxPEQuYGAcK+hx3XMcgiHxM
T+HC10SQADKE22q8y+YdC/6t4W/oE1fFHKBb3S1Qz6t/rPKN4ZzB1jJCJr4dqkl9V74yMr1vW+YE
Ynp6NAwKX/Xk4hb7BHUvKT2yjEacqTZosDVVUuy3OQuKX/uFulsByuK+HJxPznpCkMcgPNZA3lrb
Ukyp/uN53teX1pQ+xb631Io4hbIqXO0VukDMbFE/ZO9u+qXznAS2GQdN77I5RojOIb14nKAzTKRH
HhNk1ZjzXkKF0QZHrjRyka4fY81VD9QHKPrSO6gOsA6HPUhwvVZyoQtRlES0xJkD3A0j+6FMVXAC
eTAIdvw6Bk4gIviCWnq3WRA1Gg7hLHMMWvx8EbbXvbNEBQU+G6q4WPK7y8vhFGUp65303Twu3nHs
MO+QATMhrm3UkbzUnd4JbykRKH1TC+099O2js01S/j6s/yA2mt7d1PDsVqaKL0JpznPYcxlveO3S
SZCHfe90zdH3XuEuuLyT6jeSFq6AAyk63aIsgGcRVI4UwRNQ/9OsVe6R+3HrxPjJQZXafUr7+YrV
24KeNPjoVq7tkj5ZL8hcJzmW+rCH9YvwtE8lkHqxjSQEoWmA+tL1lPMS8i13htb0IxVBdr+I5leC
9217Wcvz36pPD3dbNCFu24VAwvAs908qvP9Sj9wKtPttxZYNhYsvABbd2o3KHdkG73aPODojNoK6
aVf1Fiet1aI5G9NRYzTaGBVv8sRh7K6TXoqaLCiF5Xwsz19Z/fAOQ67I4k1l3Kaq5Sb0uNetWgyX
b7aQ+NnsjGfR2C3oTkFMD+YgA2Qfmoag7B7xm3aRaL65EvyAXkL7odDbm8OC5qh1biF2fYoZ82Jg
x+acobgSYVy7Otx2Np52SSVUPvO/eGYo7p1dZUYhQUXScgRPXdtfqpAjUczp2SyGCEPU7PVjM0ne
lLUTt4lnt8hJMMJRR4hOJr/C/shSEDeGShLuAAdhWhViKRveniR9gMagfsdA0waKJkxyyuSqQ03v
wBELKLgoB6edmc0Ftz+l7mDcm7HzIk422Y/CStzITvO5m2MhFOvsqFrCRhKwfQzz2WxCZDobpN//
CmyGMjE0/kF0OG6J38qoaXbZhxshJh1Z08L7FOrdaoBlPHY2iuWyYCBu8+qbTJI+wkJcU8sx+K/q
upzoAHJu57XaXdJrN2wGzFoqAsR0Wikag4t7nEQEu9lfr/IlWzloN288shjAUbn65UiXJ1w9WmpO
CexDRXUscC1KP/OPHDE3zCFHXD02V3eHoYG51qECWppT/zgMMHZjtdN3dZnp6k6tjs5vonHNjg3c
FTgAKWfBXsXSobgCMJvxlI/hlL1wRHoLr/ejUvfd3f8xRDlP6SQkPED8meSt2L8gseqijRZy2c/i
sjuE7QHJPOwZ0Hk/0EAv/y9Q/m3qs1rHgxY+a5ghePGYDy5owF8/vOSdA3Lrlus02JVd33ZNZzdc
KKG7bDtvul64xUfpr1hWM+WlwI7aOor7hiPpzkX9QYVpO3xkN2KbBNs6vaiBngzPsCPgX4szJHnb
bvDAIsryJFnESn203WO57fJBw5r1RYpuVdmce2lbjVwprdchgydVHbMJjTEN8meyJbKGcIC/MpCQ
mwmoEKeeS7da+5tuM2ILertdkcVG+B/8nxJc4YTTL/8sjhUDhVbYp40Dwh+C/jQMJs/GiT/1VHNA
hAptjp6TVUN83ZWXOuXxnFLZaqrt5s+AvKfOpAgTtTLnxe7h5ciIlijrymvKVixf4w5jaGGoMNXs
w0CxO4g9mij0TM1HFZxzO2+mtW056wi1sZ1t8pv3bY233ns3ayWj2NeBFeijsx/Z1oByDbfyRryX
DOtu8Q3EZhM7b1fpFu/pMMD4Y8T9M+FIpcpRCO/3Sz1wnsukRcMfk9ghD32e524h6VVTCxxnKBrr
rALO2s+FEyht2nVoLgabUPlwHiAIGjh+VgibxqNT8rw8oxGcstpoyi98qEyXljr3+lYOdhLQGfv0
P7od+z9Ho8JcDWq2qAhlLcQrLepc++YzatilzN6kv2L3wb05ozCKok1RsFZKG1GZ1dp4FChuNa8S
Lxf2F3/qxI+Q6ch/9CUoTv5EXAlgCqgxJbj4d7VgYehnnkxKwpsIEpdhqRp3PXOSBry7zTktCbsi
L0l3gYD2et/SKuasJuQq0ccXTGugT5c/lCFZejwgGdFJeE6mqvAjlyn3fMiMoLc2aXyfFWafb1Xm
Oi+fBAQpjdxxkhI6l7t+0vwm6upOmFf78cz/RY7cCIqdqqhTNYuFpnSmnb6w44A6FFRq5PQb1kk5
qenx5R8XyKzgKSuk4GKj6+fOCbJCEez8kuBAo5welBtRFDH8903wob7Qxc94rSI0zdoeJMX1m5eM
d631qqP8euEpAv2HPTLzgmE8wy/JZTJAas5JAigmHOtQsLPz7KfY5vYd6InxU73uF+dRFj5GTnYF
OWAHc6/r7yVbNstOQFHJO4WcK5JGny5/zbdryNMiNsuCLz6cuQiNar1uH5A4zQI1Cty/OtMn1K3k
Kk12ouMUDjdYz6vEM4xYcOx4bmt/Xa+vE2Psoc7KDHQeSW7n6Hc4NgJKSvzvdxYt7VgOwqh423gs
agh+JqdjRG5l/28i7u3cNCU5FYolKr9R69vZrl3QaAwK5qkHN9qKM8Tb7Mf5a4zHMRLyO9SzniKq
f7E9cid0W6/SUXKZGAsRZPxofVol75VA5zgBh6xJOJqGCK+Qn8DasgdBldp/OS1nrCiUOrh6b8GC
kjKjahRj6HB6VCdpjBnDg3lyZ//VxmfnvJF7KDrID8qdbeGWddaIzgcNUqf9ASaxbTpb+Z85q4Q4
Fi0/IPAwkAhX2uG4GgvcgYQqPnyVx9VBj6vA5Xi/OkTGinRXVaBQ2upbs4HHZlk+Tn9SuEreVgjG
m/NZMjuz+p8GTUXON7qYZS6iAeJOPPzWDxgGSalqS5QrrRJd9XMgfrnNoGBeOWRYPfG2XhGfYA5y
HFNt/rQAp/SKJmP9gYEXpVgU6x9QcmFUyuuqT1giDBk/IrDot8GE7ZBEy4k3dFgYnEDqU4qgWLep
XgVZdJHTYaCovNSlPhq6d3937MGf4uU9NCcUSl8gQjmyg3KyDKhKvvEWHmhfNUiTFevuwuGnHHr3
/wvmLeLFqd9cyTCPpZ0Gh6sslqHFs0Bc8MxozmZp1cW27ZIQDtCOtLMfwCakR96et7OkQbQ94TgA
YsMSTOA9FpSDgBJaamDuj4J3/7SWtAzlYAYdoKKgWh9/vM6k/UEwp+Rp4vRZOgS+xFFSV+fNrD3X
adx2W0SSsrt2CPdP6Ke40BKrt+NFC/PSlWsHYOYPCCjY05i7H5/FD5lBjFIu+ov/jHssoqEmmWnT
+U9vQHxmMnCHk47P8U5uQkahI4NEUcpO+OODmfHYYFEx64xgewZjEq34M3Ks0SrksIDaQCBcZPfP
+AdxAwYfTfDCkAnZWHNzf5bZRJqfS39kHT54W6YIeesMXjcvfVDa9YRLurLeA6+wZiBdBdObBPQE
ouSASnUL5b4y5Uf2xSC06wwE2S/6R6ETpFIRdAf+LKA64CuBb5esuM0CYW4nwjPkTH2neuwHpMBP
F2/f+IyJfkWKwGNbsXrPTb+xAcsZ22LRhllwXGpooyq9I49SGjrQeQa01XBQoY2Y4t8kV9x6spT8
Jnw9GcYYWDA+3yTv+X5+DwyFzQBEwSL+vOHx2HiV0HSrPgUtLUOjw3qWQ96PLHJk7lZv+Y0sCvq0
piB+dRmqT2+H9AxOmNGkXjTFGx3PMiiK+90/ZRHO2pEifa+nCq7va2d35/xompCwD230pjmCasHe
UZIm4k3czQW/cq2a+yhh56n9wJeCddXFM2DyRWT4dm5Kj/nR1YIamdsexHEhvqN18Js1R/O57M4V
CjxWt4mufMUnsMqVuBZ2QQBQ4seTkERqt7QRe9izqxrISUwmgwpCzk+OISrYSp3H+Ez4ScpgWhwh
Zb0FnGgdD+XH9p8OGMSM4aY5BeD4F7Dt39UGqMVJJ43jpV2SooedmeTkwHvEQKlWXz+QZZlPxAWq
kkl/T3utxyPBvRhPEil4wq/fwS7b0aDG2pg4v1JEJipkHRBLzwLLFStax7ZS68BRpnPbPi2kidQY
sgvX+Arhn6J8FqilZlPO/84bfaHybbhorKFFvBmSeRu2nHcJYamGceXJPvfuLVA0gmJ5UkX5W7pp
zUjArI8j8aNPSaicAVducHKiqmJSeFbDNDZp0ZL1kkPsnaTUq9OhIi7u0Gk3udklshYsl8epULvL
MBU75BXOtznu7yQ9/au1yPHWkuEcMjCUYxBIWUAtVL4R7psd5fkRVVaplXQ49OQ4cGST8JQGyPQA
j0zYxg4AQ+xXJfEQHZMlcDZmITYIFnIAzfp0UlpBEu+5EGPe7LA/qA+bFRWIT91Q/Odw7o0tYgYr
Us73ENXfIoR5dSXSB05AVe4sC7LYARywJA0QxxrV9mTfkwOsS4/8llt6+9ElayHodon8pcZ2BZ0p
owGbfHctppqUllh4Pgy1mzOmx5Jq1ylKIX+QTLUPrO3rjt7jYNrqxehwQ/nKr3VYSoorxjC7xPLR
t//LqzFRZO+iPqdRakmGx425xsrCw2j8zFiXFZZrSLpwm8QQUjeYlSMdXZWqILK/GJCjb11SxHry
PqVgjFXk6Q79JBvVUpLnnILqInTcJ6p46YnU9AHrsNoX42/3g5ROzkAWTRZOmFc6jlmgzjqs6bGy
8RbV+PSOOLvmv9fjQDY5T/h4y6ev67jf+gMeDLIbtqE4RRa6bY/XsLBKN6cKiU6iJRBNilG7Hnev
GkFICdjBFXEIHEe8WjHEAAufjwRRtrnxGPPmhu9sbh5DNqDIpsrfpHccrIzWlDvNevSzs8cjsRlG
ssU96rf9XrEAk1fCswtk7cH63aOjeYHxdSS36RoSEJTsWoecaQWPN8B8Hg0oPgZT6uruVcGZ6wiF
dFb4QyszHq64AT8scszsYPsP6OAPshRx2PEXYj461uvvGjOMWxwZMXy0b6kmtHo2ypC0dzw7lhrt
M2WS3sVz7jFWk3AUBCedewjCf+fFKEUE9P6paPLIoKDn+KU0AcRIXmZRxYt8fBcixejC1971ZqWU
RV06rDbMNFWalmULyVJyDs9bcL2EG062bYeCBOquSf293TSCprU0OP/m4Oj3KCzGOry8kfDb9DZA
g5CoCxnX0obLP5vhGbSgmWce5RMyxzfnbvxILg4PsTvWF5xy9npzqr/7LiE8yo1GOJY57BqEoFS1
eSiG2qgjeUUumF+pTZp0xTFGusL8bFWR5vnqHkDZUfBTK6d3k0T0MVwrIDQD1HKxMSzEqUaupCn4
sgjKQHHO5ZeEhUFsZtkQm41Zh8dqPjrEW+I+IkYjsswQ8XvckByEevOgV+E+qls33RrflWxEC60d
HcwYY2HHHmWockOUL+MHbcrg8nqWaUQIqdHen3s9tg3Q2A6BYehIZTXN132Ah44EhgOSh6D27txP
xWJHihRI8k9In9Q7rGiUDNa/4Acgfcn0NEEUxjbdB9Hi8mCHybcFi8TYys2DLd1/xXf7AsSQjJm/
w7Vn0BJYt5tDjBuaVYEd6rAuc8dhCPp6cux4SC/hPW5W5/GZlJShWECLIIjGRyqBicE/qYRTJxVi
ItpRZEpLS9dmM8jDUxvr5X92OL1uX4mQGXGC23kCtF2d9j0Xa/6UzzKqLIMEP81CetEQkNMM9zKb
JF/aZWgbeQMM34Y2dTqG51mZlTPwkscALeb5QNSFsNbLzh4WcBcVl8m/a8szin7QGWODTXfG9EDM
sq1XHr+32PW856xV/m2aQI6E8qoPPIFUQ/TVw1hKCBT0JN0uu7Lh4b7AQJT0t93qRny95rkwktaA
0xzr37xZ9Ag35oRq2GAXLYK3O0HQTS2AU7atyKRavdrD5MxCrcGIkSMwbfPS/5/EoGeKiDOrim0F
0WkrRjN2LoVlaQmQdBhSGbaEhIfi5I+qX9nC4QMeI6XU93QZcYN7RO8YPxzXK4IWsfyOAiviYcOR
bETjEOM9b4dYG25+8wfFXe49GlfX4sHMMnC3X9KH65abJFUrgcpszE59DlRZxgqppV+cu856UN8a
JRJiCbzJfZL8Nl+Z6f3xSOGvP6o9AeOM8XdSqs7IdFacfMaUCMxCew2H76tO0GRDpYiYM3+DwEB0
HyqM6KWJq7JF+UB5aa61ekNPZIzAc3RBzPnYSR0oWX8cuT0cDzzThE+fv5MRA8u1khLbAuDsKMli
N1+SblCyZ5uVfTj/pdMZnrB6TrFFQ7yBdSLa39tOLaNhOw+qmzq1/w3muZO2WCKCwUu2LrpjgBl9
ozjLhdNg7dqOl2gBgQTpIBp+epFvymGPx7jC10Br2yiHlVSJ7y2h5kcwfjraWviRWze1JZAr4DxI
xjt4BitekLiYPPqGtk27GiO3Nl3MLXsAcb2WBQIOdAXZQ4VdDlSlKADk6x+LUxO9TFxEcvAQnUcL
fzcsKS0bxdAT8GmZEerqSkewzTgrAYzkBfmNk4KdpKssv2SXnTr09ZHabIRULu3EGOQdB0JO7Tm2
ULbT3FcZxBoZYGUPf1dNtC+3DnrwglRVAdgrLf7aNlE57vzA0wjmmgUAFtzButhwSlnTqXjrzA+i
OeXVPaXbDrkZdIb/BUXNiWh8ykqGa5JokYKf/XX6cxWKZyo7R+gPXT5iSgDawBMDoiyTw6st8VCp
Hy4mAqbDFfraC8p95cGjeJ0Ek9WC7qBDqcXOLgTSnesjV/EbWRgtWDboibcLIYpZhiIZo4yIKdnE
Tx5ueK4/+3CdqeWHZcHrhe1S33sVgRIIj5xLrV8jDRmUG3ho42xJtXmx5OTEQHFIM0iz36RI8BJZ
9WJoX8QeT7L/8FCyVoo1zEKhaOKFcEIpdHN57Q1SDzdWx3UeF2HMRbhE2ygMNaeKbe0OmrNdXYgr
Rhm4XZqrCWpOH7BTMm1JsZ7C0Tpn3c5Y/RXe+zWZvHShlV4cGVkbznxfXNKwu2uoShGdS/8g63tE
SBJWVy3dP1hznoJGEIsy/aS2R1XfEnJ+4ZVxivlR8wEtA4SkEU5LqL/FLcOyRCcpT8nIOo+gIi/Y
PmsP2lZ+gzJql8UwBm9UbarS4HMopFacXaWS1VtKwoixb5dtQDdlYtCVbasx9yuAp5J8AQFKjeMw
jpCBDlK5Q7wcBfM+kWeZEekXYt33nBZKIEWkYUB1eR94GLfsKVDl7PnV6fKGzsqwhUKDz2pRJTEw
iPRVC2Ww5WLBRAxl/4e+2Bew1Fyg/gImn1XP20yckFs8HJrUnA6Mr2vKsOGSHuiZNyCAmI+VtQYp
o7pLTyopBRN2suUGkI56QifRVn1J5AbzySab3aA2wr5+XxTCvWpR255sObpwl0tfx5ELrfH2/N/u
lAojCVqDaVKKQ2/uz/uoyQdt3ZJJWMvgrpnUMav/IQVuO8iwdYTkdA0+jUxAek8yW1C79ZCSMr4u
19TJH9ZnJBBK1Dcx1NheRxC3Rfz9IPhnMOCaR/ATHyKTf7NCr1jUbRwG8iBAmfyyh8ZVmKqm30wo
jjpWUtrzh0rdXZoAwmnDDEk/shl2r3Ow7yqkUXj5xWStY3b0m+iY6o+nY0tvoiM11q6BjXFZXL/A
PBcNBEDe7IP5vaR+kM+gEzll7S2SuENQ1sqmGgQIHKamePPQNYHhAnGVhnMv+h2aAeu6pOTeUrJp
x3oDGXT1iJT5dQmeWql9SaZVAFqOGR1yi9Pe8ad3fTLWtC0iuS0deKinUgfL8NL7ZYExVTNOLLmB
nluSJEf8YpuJiAzgr007p+N6Q15r/MlfWN61vVHVkb/wxX3n5wrZRkWo9+/Q4ElBWC7QpWKl0suu
fjxcHYHr/DdqilnLkr7l8DBcLQSLE9pmP9n4lpvH148dnBvG6VWg7wGqyM3HIk301bJV65SJM338
SrVuNd77GCb0vrDoUCIIn0Xm/NwNkMWkXACdq0xyDzkEMK+g9ZvvLUgFdYv0/zkVbMM8bQjzIAVJ
Z4PIkRig96vlZQJgGwDuGGpB/Bwf2HWanp7xxL4cZjat5UlOkxfVdxUZv4oNv1yYtuwXwnwxC1+l
L2Ts5ywPxOIsV7uhIw9zXDNEoZ91ZSlqukUBe50sm07dCyXNxyzdUXMo1I8X32wgGaucX7lpKJkD
W+AIpPsCRf8/reMSHaDNz9J+nZ0tN/S8rdIykbMsGPnZurx5aiJIhjviUfts7vB7IB36Srq+XXv9
jilbW5PgfugmEbjj4bF308H2ks4wQXjaE0tjVud88R9k4SYaM+iaZMA/lSBJNfH47GipN9xpvCxx
+lVTd9VQhfUhhaEbjUt3Cb4Hy0ZONfbAw/SN1TnM876tR6t3HJD9ttS2dPwKHNLd+dJDyxh0bwc6
byNuJzUQxfBPeyixstSsmg7ibbgLP4b114AZOXOpOFoBWb0dmBe6/B4+S2BK8/ChJZezG8CjbjFD
QU9Q4kVj7a5NJ4eccL2Vm82Sx70QTSKDUD2N9OYCIfb5oZrXV7ktzOeTd9Pd1Z8jY5m+5mUZTqtT
BSWAiC+I9MXZGiUg2RLmtLT4y9bjl5ji46jMpeVCSaZx9umRKg22UbVOwNFF4ddpSGzC3cg7MAhJ
KOhCsb0JAzJuey0YlJi55B73EIiKouDYgIXUCTZ2Ui+2RlZH4PkDivD8khD/sTd8v5Djf0WO8Csc
l5NaPj5GqRtOt9taFmGP3Z/GmPobOEe4QTZTxQ/+fjdJk/31JQn9Gh8BQp44qcK4Ruvm0C9JBtyB
BklLbIIdizkFgHknyx097SSJviQarlYq5kSfOyADCx5rdI/5YYIoySn9/EngPA+BTOdfieQ9c1wF
ZC4UyiRFa3BX39QhorXsCdwHh84cTKSkpU/IPI/w3Rm/OHGE/7yY+wp6FNSZNB4BCqUyGsMGpBr0
hIG/wgAHP29FrzCphWCt1QOjiUV3b6XE5AlCV6E6eNX6NNscRhS6hv1vNWlVKZ7MKyMbz6mGgUZp
c9OYa9oHvz5xRXq+/iPnN0G+g9vtvbAMB+Z6FdLP8UR7mddxXqw7fYPHJT1WhOREw4tWmuVm51KY
dSt+20Dfuv+XJIXtO4N7xIliuCSYZ9CXMZdIIF17GAmxSDzWolEOLpM/nG7qXWbuIPwYFRX34Dg0
YMcHbsM9abJQHRqbEvxSTaUs1yht9HnBm2rFGbCmaDpodEMDs9+g6lKYeGxXe5DpDiSfQMPEp5OE
4jnwGUFuiaEg9LsbEKDtZiyU6wY/bwMZzTbqc0J9A87gjDKMbUq80sa/fJ/pil8T7AglDvw50D1Z
Zbu8EQHDxc6F2UgAN7czo0IRFmku9UAUp2FiuzlvkY07R4+dBU3aSryEOTgmYwgUDhyg9FoT56Dc
hvN2dq4zXGNkTcB56Pzh50zbIiewEIIE/wIukE5H7dgU2jVvcbxMHDD14gJzwlfRPh6Jp5G8m6U1
7xqFuvrqulODqsQDyArb4I632GcpzhO+riedeXrxJl++Pl16Z75r/P9MGY+c/QIISYhPdb40QAhP
2f2p9pchdmXaZnur5aqu8iA/UMYTuGgZfSDimD2o2XcmmPvKXLUOGMuR3x+/gOQN+sl9Emj1DEdh
p4Ds6zj6SyYfCfTmDWaU7suH9bHswv5JAxB5UWE3oI7yscNcBlirPZXa2h6V6csrb9h9GJL0veL0
SIlNcOhREcPmWds+CkL0TOkJcc/Iz1zNv+zkhzxBi/djKGQmFLH5iEgNd7rTZH+eKwFlohkSXzMG
wae839FsUm9V0BOZkvNQHVHDyT2xIbZQohJHhEysJNjQ3Ob4YMUF8kIFrZi4/iPAPJhjatVM7Wb6
6jYip0/767B8wnEVZLArKpp58feiR91dB/gGdSohbOxKtq7jieTNTkzAmt3U7Gj48WUfd5JWMT/S
OUtnNKCiFYYJ5J+FsW42SzLg+CLaDRRmSKg2JL8uS0JTBsMYdNbtMVA6HPy4oEAaF6fsJ/dJJL1X
RMazEH2VlcAVUzyHnTbv1sygMGGYqeU62UcsgKe+Uk63tq3gl+VCIeWr8xPSdPAayfvwITUEJp7r
hsb4Y96RSiyb9pBtWFQYWJv6RFPlQmGOG9WNrXZkVcXcuWxE9/JbSKxmm+b0B4NddgboWyhjof8S
bVq67Zd+US6ZVlf5iFpiNZ2S8f3gPQFulpHjxXqmsEixCvL9EFEDwa15ty/swy83wtlR6kRXKmwi
mXsO42RcaKBkA61N3i1En9O1flZjT4BHkYQZspgMbcILx0EzA5WSOgD0QPMz5avye9t2GAjGPqVU
ET57vPY+oC7/HkT0WIHHyN4npy//IjWTj/yUxRH6gOzVoUPoOdVX4XOUa80IikV5dSA+tg1Z3BJ6
3Q6mn0fzl3ilLvfABPgeGStA/OxON+s3Bq1xARPl6fQ218Ae6F1nZlKEfu8QYGC7CrNDqjOlqm0s
NVyj4+NA65UwYHEecsAKGdGXtS4anPIaSaHxcqrhhiY1DmGDfQwFOPqx3mjYZ1dNZcX1oLPXEVMD
4gneihGx0q3h6PtFfSmPbQ6ByhfqQIAG6pIbfvMmQowAWyXSwZzfNXndaN+DQrjt2kbXcalnNf13
wH2igDHNOXPinKBDHzDWsIo27l4hJToSIhK/3fNX16nnbzGUu8rxxYf7KuZRVtdHHlWW1AjRgxFC
UFr+TU9Qhl3+nBCo9HQKJVfQlaCTNUc2FDPSOr3LA5X+LFftDpJ1EGWo2zk1QJiKW2wzPOdX2Hhg
5dMvYt6fJ4yX0bLuFh/lctsFZ18JYvZXIDqXOqm/V7Z8KaB0ZVBrpIZe3dG75QI1+wuYKvAbv06V
GzBaMJzKzxSmIUovakzXU3SfcHxUo4v5o85faAN7k5m+XeQzcom/bCkk0MZPIJE9yObHi4Zt1LM7
r364biswrzwKrGneWokoPtFnOTdstp4+sfdeIRG8VtL6V9GAA++JdlfnpHRjh/tw6NZbrVlrc9j7
lv4aIvpVUiJK1C7x4muBz4cOwhm2jyfLnmH2pz8TNXw5EMtguDLWejlE9or5zVDvL6JzDuacvTgc
9vSkT4qj7BZr5yAz7f+axTEmknuQ7dCMMAVdeAaTREmoDph8xZPVokA7IX4xlt/F/WA88lJC6Vgr
QIDb4Pz4HIMD64aKpEQCoBy3pxjsaZ7UQ2swmDhPITpEfeoE4VaYFUUGEAqfeVF+4MmxEGrc+VJ5
klnWJW6TpUSJyYSDberrS0AwuQSkh1koanw1/5OB8ALt/lsFELPIYkIfDqRBRyX/N+0aXdvWOUM2
UHanDypjL4YKwYMoMYOuXOV77wrJ4RAvOV2kqMjfnA6Cij7DWhZeEH+KTYWtrf2f++EP+ukHucBe
PTtAzbts8e9jzuzsNuxBk/I7A/avRpK1MD+tW9fWHMvKgMiUJyMXV8L9ruzEayKaitHg2heBxq7n
A5kNHi8ZEgbpFpQfltSHAtvjAHNUpC9cWy1uE7/SR47rAmrw9Tz6ZXM3mo8vhWqDFCrNMriaOoNI
Rmd8A+1gMlcsNx25BCFf05UsRdQ10c0Z+D8cyYU1spR7dYTUNVTNI8GQuv8APvGX/Pajzrq50ozP
8DjmW8CKy++ytujHyiy54qaq8eDvAiPPTNLV8xfzpPf4vcqhgJ07kupre7gz71M/ix4OQqWekV0B
ywpDhri9FQjQ+MTkFf1do+BVhnqQyVzkbblhVN0i/yN4ofFdjgWjgLOAnQrAkNzn7Kg8qFcdROq5
ws+fs8ARozUUiGGwzwTF2oOo/o8zjYMpvWnNKsCKYhV1z7XxwBftvPST6AagW4wwmmp0KSb2deH9
YwpEj48OA/a39YUWIv+/kwkmi2AFkC0ueT1+9ICgPfp47p7xVtHxLT5EWwFBRGvXYTVmrUiCmuv0
d4HLyozg0N4CJXBOYYV9RYWmy3gVVL40ycOaNOokHLBnuymUxNH3+WHAo8s6veTQJaFcBEEYFWg3
YnC9EpjqQX5ozxCyDxLFydhb8mZj/3WwcvNZKt1Mvs4oc4kDNQazL/21VBce5aW0ZRtHju29jNkO
XwF3duwnBLS4lkAn6R8gzIPoQvxG8U9W574o4g75vOCzAEyij6Ll1RyQc6QvHDAS4bmP7sDTGj8v
Dkw/7J+c1jHrc6zBWwtUNH9ix8F2PRvfYfUNk21xmZ6aoYvozpgOJ6un1AK2UJso6wsWfAeqD47r
TJ3az9eYBk3oOapgkObRzzzHfXT5+XAwCFk/4VPLO9L33/WFyUSNMNEd/pRbrMTKlr/u89+dRMOs
XaCBC7TKg9hnxo0Dh96Rr9Wmlczd37cMThOo99jy/EHPas961Sh9Gkjeg0BfoZVyB6zYg6kMlNKF
FI+JavKH67zHpMI8zfoB8cPXpiqdH87Qq61+CWNvakLFuQcgUzu0OuckHCWnjhvBFWbauw+PpeCN
uaRRYyKKrppy1hbRZZv0f6j3leYRuMHEh2GFL0fmxIbGr5zKQtoBrN4Uv6ta5iPw1yiQrF0PRAOD
rPRp8Kdwi2xbZT4XZVV0Y7V3YdZ791shJhd6OtA2wfzw4zv3oX8wUiwn/U7Faasc9lI7MrQG+MEz
oVVUpyYtwu5DWKwg5RTbRpKuGmBSZsSzs93Kt6JV99Th3YaCsmp4qmfGka6i0avWto9Td44MqmcZ
nM8nD2TCnrnl1aTE6GK9mmmHg7Ua7e/T+TilT9vAgroKxDL1v/von50tzysRswzrV/l9HM4sysqE
EwsZ7QcwO8x5RBygObRd0cezgTz0X85YShX86nzfC2gFmYv37bfJrpLwCSfu4QNkQo+a1aN0/mAX
2obTRn2amK2ahaObWvgMzQ+yV7Mf3uYpVHyTqbBSEX3wh4T1eVbkSLcQYoZW0aOPATFLmQAtloI0
wtaivNf91KSX2rO4fjy4ypgWYZrmmsAJu/Q5ClQoSPuLhdZrAl9rX8LhoFQ14K9PkQDRbcJCcWt3
9zVXAmLAYREQYXwPWy9iMF4l0OvzJlw8a00KLZFe4JcGRFKA0k2tN6uh/duFvTDunLYgIg0B8bWn
0TWFXyMWwPNa48PK7a5NH/+Il2+TarRxpVFsK0KUuBIEhSkcnBntV0gmuqA3tCnMgzrbF1y8PFcw
evDllZ4ABNDqIso/aamo2ZLjHaeRwvgX9lIuucKhr9s2TeOKqxTNZnTMLAYrsvMRmg2jTmMOcfSM
XoM/eNBBV+/rG1CpWK/R6YwW5MsZxa8XoRt6XLQpPz5DdD1Pxy7ff/i1S8gF6F96uObuc3z4awr8
G8GMm2m0lXqsnvYdQcbyXHmdF8YE0e60Q19gkxW90icEMUtnGDK51/4qFJd9LkTz0iFkEKlaUSCv
v+kALN/ExIu4THd+73wvRh4isROARZ7Nv8vGX93eT9DMnLRs588RXi0TjUWuuVVWHAW2tIvR/YOg
6yXyeemlKa4NqEnijAAQnSKDVrsodjgh7AKfcvHfvc6MExebhoJYRwTP9nlDah5GvKUf28kc2nJ3
umAgerG/p7p5O0e9ODIXw6SJnDCrHB1007iyalqkcOI111DcT63O0SMgqTfnQpFP/GRwv4GrgmfS
tqGxwDHlNKsxf5QGkrzP84X+94ksQ/ijx5k2061Od4gPuGcIAii/V+3BVBJVkLkvhh/LO7MQbrUI
tE1ne9wJKQfRJJgeRYE4ooJpPaeziB+kla2VSfYxS9RzAX3EkP0z9UMvB/PoFrsDMLdVEV22tDxw
ewltX/O6Nfs6tgmdu5o3cmJeqdPrz77xVloODPLbibv5PkYCi69c+xyO/Uqs3N/Wigkjf0e4sDYo
f2OfLtaly4JVS/fHGZwKFNCbMSqC8SesD2e4tfWBtlsk+KsRGQinOMsQQB5GPb/Uvj+lAt/jsKPY
WX2WdEPC09R0awkviBfX6RdwANTBP9weHvV/qJxrrRQ+J9A8ED6wvprNPpbAm/gdk3L41THGoGBB
rvMzuL7rAFXUebrsCWMeRdmKxbTGblvOrI6LKf64iX7qFzQgDzXZLJzs3SQYaZtH518abLlSuB0E
Brt+pw7UqTzaZ1QXA7ylKlGq3Ja1Nkdc4+PPzJH4t/xc1IvbrgSipLQfoDg5V1pfyomSD+7OPcdo
/ex1KOAWky/QD0l2yV8kyE1Pd0g2DS7NMRx0D1co0Sle+uITP5VI9YTdOzLQBBdyjPBnQR7GVPkR
L2cqRQQ8mg8ocuLicEZoYyHTmFRWTmj0HzmDaN00DcFL42g2G8hwUGryxlEzO6zLyCh+kRnbilrg
PN4fTltzGqmONmXgTKRB9S8+eGtfMIJtFk/RKhF1Dx2gvTAZRC8VOIY9ASIo3ERdl0b2KPu5CNEP
yEoADdFha8aPPm9y4TaYxEH6Vo45U09w4ty0q24PjWLBsz8fzhR3eUm7IJ1C9xivIzC0h/uQ/jKQ
TnZV1lEaHAf6kBICb0rlL6pBgGxjuA+nULeuhc9nLaeY6hPoGVaspG3zziLHePGUKc/i4ToMYzz5
GMQ9IzF1mBAKKYldQVckMweHOI1jQnZBqlCRjdIuv7WU2YDJSQ9LoAha2DABSqVpOHR+10kOiEJO
UlI/bq76c01er7GgSwJrQcFHNFjXmQX38juhSzF4eG9jP/HF/VZeu8RwU7yYWc48NaGJZDtvLyA+
FJoC4tuKNQ9CfCaT/f4gi5VgI/wj840POj7VWlQGEchkAdQxX4XsnHgROqXR6Z65vvm2Exdepa9N
Hi0CLxJY0w+QL+2y/RHBxuYRtucW4uKsNbIl+TH7Di38EQ6UUMEGDDqrHHTQ65+lg/u27c2KSotR
Tt+3Ohvtdo8y3l/Li4OxF2L+qCDYMri+nWrIveeTPvHH2A7p5AVoY4Ohppy54sXaG+FwnwjWBNxK
6ExlNhyQXmtGuiBVjAil6bt/1aNdiglBdf3qKvi0zHBTLiQnMVima7d23skSvd8X2aolKlXdwyQ+
6vLDndWNmSNFQyK8lt96zTCoJoSHl5BRIG2jtCFRZDSrJyfAEa7SRMG9dM4RAoCZ95KOCYWgP+Tf
EER34bdvRmSDN/plOLxhRI6Hzxr9g+nTqoewhyjRe5muIJA7yrnk2nikiSHHkDDV57xkchHmsyrZ
fPXILwZUcyOzx9d2Bco0ffVmNnitaFtmedZrI3aIg4Df92czA5AkOrpoYPngLSC7iHG2bEtzMDy6
YJOjRDfxk0GkrPRmIsM5ZQWcwNPR2kiDyHNDIChV3Px1a4HMVH4KKA55eqWfqRbBbnIQGRTAZyzh
2/0o5nPh0thJ0J5tnH5jdmN1K6OTIRkzWtdgDTqCJthcygqUAcsBt9sB0tIW8FvC0Csv5FH5V7Wx
laWR2cdxkDX46rJLO2IsghoslbOKLVImlnGHm+Qay8ZXH7uHVQCQcXFRh7FWme1nJY3pjmHoBDPg
3m+1C95BUU1FzeuAWPQK1mYlc9r3Ow5Na5isRxX55Ikem4DZCApHcdeMeUBqzD5Fb2WgxThOMGYr
PtJ3tMkE69oAevNaWx00XRLIfl/Ad7jSgJKEfAGpZ2cLBO06MovOHxriwIGtweNk0DNL1Jg2Oan/
IkX+gpTA5svJ28NcqBbH3Pw/w+V3o9Kk6aphYRDFE67O80C4UcmKoNbQ7Kp9wi8xWqiTNMzQ6pfm
F5skUNMUZecgkv57K0E8Bghmf7aq8gXwXzEbVGFxxtt/91FZkef+PIdNAZbjgHn1oa1h3tKOx4nL
tO43BxlT9lRUKZUo/OwN/ERMvZcQTM1hxEe2P4dYwok3iEtYjps8wagEufZGPJyKB/ymUboD1SGR
/kixTsvDZonEeWmVNHEr9XTClpXBy1QrlkmYBfNu97Fxos+HT23Uf0VPyHPvy/5xm6+aH3/o7edJ
QudkQWibEYi7cHJt5faXrnKYC3b9ia2N/lpA8gyV6DF+zB8d5xQokRiHEYs3HGyaIgljuFhl6aNA
9QhH9A9M2ukRnzHBLS/hps6bOJJ6Lehxaw7jBkG9+abR1u+upjkhtb3xwF0TEeYeUArBZikH1rqg
AzSEGKvWh+M4/bXoPCDqnB6ln6fG52sIfNGgxut2A947ttP4QuU0I/2+Ic0lKSSgQMUyspH6FTHe
1Y3skikzdyPAtT57EDIqDI13MFEODgB9WBJyJOXd/8QrIpk3aRPjFLw5Tr0xWFn0QkegNiDOpn/o
lz+pb2v9Z4D1bqDM/znZ8XPIZfFYgNVaWQTHh3RDFOwf62G9L+T0kqCfZZjfg1vG+Kpjs5ZMGGU5
05heQPMVDP96HXPWK+9UhnTzz6PLDT9Gi/d8060UuTR1Vxj3EYCh/iZdJyyVnroNupxZx2w7u9IV
H1hgkEwXAIcgNlbSkfKci337821rpaU3c84v5GuFop/vN3+RkzioNFJ2eoEoXnAHok01pgnqBbtI
3dzBVNcr1evaUCewyL53b11xQ0yjgRUEMVR7RJlWQfH3pEPAY6WNLYdihTWPfaUWyO4Xw7o2H++l
zpBJXTUdje1pII3FxNTu2VDFEiW4jkBn30i/rXqZqPJkTeYZ97sOeBc8X63xMT+K9LXm93AnRDQy
bW4wMZQ/l22eKvrqz/vBMLb1BWpzD7V7iU++1rxDZQ8N3Ei4TlDoX98Wj+n2RwveZHjzunZfl4nu
tXlR4KN73GoaO6FmFM+vnms3f62vtzYbdwoMKoAP6BDk5H9ECL2OyO8uF4d1XbVy/QD1QhmmYilH
zzKWYaDAwZyadSK+tuq8xsr4EXRlpZNoRJlQwhmyUOkNQsqDYZj6R+moDJZsNhOEBIhgkWqfQkGP
V+ze0I36XuvXE2UoNVCiIlS9F92q9YZbSKe1RXMivz2Fgfa3oniFmYnv8Qb8KmlI2+ykvfSsy8W0
KTm+c0HbO4QmqnOlQfRGLb+A/u6gLbkQywA1mIi695mj86Z0LDXtIveGLXo8Hbh1eJnpaiqflVD5
ZSiKyqdvFDErRhVGS/43nAFYVBzlHbM38ZLCh1OGYPYARjQPGAnMI5OFU+ticxIlRx6U0GWGr9Hc
3kFr0dG4v7Xov30J8Z4l44W6ZKlHAUlW7Ky0NTKdumlwv8x90IyelpTwNBWwEaMtq1ax59kkdYpS
3aRJ24ohgN/Oc8xf8CW+OHqK3w7RHMATrPSXFtu4B4UOkbv6AXiYrBxUkWMBeBBQkjcftphhT9Qm
v1rWl9eMynAwc6SljqAb26cjWSPCAVD3aCoj8a+hZeXN/6cJox2qxd4Fo3vKuajrpJix47g2r8rd
hxAq/TFYL45nvfiystQnWLnqUZXD1kMA25eStAhRiaFvE5OOijxyWvsnuAWP0z2cVMkEGa5xUrM0
i6p+ACL2+FdfWWrjCY1TIl0F9CyLFRReZryz/qwxRKrxqns1aRKId/Xu/kbMxCN/2VyBrO1fZILq
Pc4zIQJIU6jQToYXMDOZ5zQ5BLtA4UnM1V4x2ijSzj5qqhY6qli9+H47eQ/rbZCVXpJkJGUZ4fcF
f0qfhka6Tiv6MrwvzowCfa1Gs7/9TYpyzcOjDoFaDfYNUBJHI4ynd5da6s8GJ/BeoPyH5sgbfsUT
eDYPmJIr76Aj4RxpquThO6vB4KDRHmVoCd42LOLwwfLbvOtJIhhWeLUzgfC/rcfsr0movRmxq+ZI
iwOOzuIKcFgqXHO+QMpYowRURXTYgSTLdOpR1Xklpq+Kvuqin/5s7HxrPjvIiUA+qhE7KcTEX9Uc
kmPB3/8dXgP5zBG8dyOiMxXOE5I+yJagOhtRwtE9EP/y+vYkUidC4RAs8GmzO4xQ6o4fbnmVu4+s
7FofyJ7vTxT0pXka1p0dORsM860PZpU/0aKVx0jAB/1fq8yZdOTe04b2Tot0FUuznsEWOgJleEyN
bbc+dcGRA0+4tNMyfAeeu1bxZMFRgi2Qt4FAOHHtm9oK2XEvoUngRF2OqYLfbZ+j6ff2D81T6VZi
bZeisr9x9g9zhGQx8DlvzNn7c7vtJnkMdl1xNR0XHpK+52h9u3iXFPwiLzPjDB9IJnmTJcxgjsJu
wwSpkOnkc3GDMLUDsxQ0gAuSq0JTUKl54kQpJqN0hMW46rcbPv/KZVTSOuhLAXZVN3SEWuInOisM
fjw9ORlgTeZ1YchTUt7bSnSadmJzLzsxjjlIV2/IEy5PmwRyWXJ1+7s+EGx+9wKm15aazd6tzm0h
YjkpmsV2GEH7r17gCafk/oF+QUjSgH76mgZlmsDpU/SBhAFd0jEoY0RrOXup7BgTZXfZeHmz0H/9
Td4rIwGHU2lt3RvO8IyAituVjpXtARtNBskdLnbzkzVA2KiRrJH0lpdoU8bvsEJ/QdQGOcTe6iSN
A0Zs7g7f5NCoOPWp6Fp+ncI18PZoL1DH93QqkFf1mYFALHJE1rko1kfmNKXOO8AXvSQiGOAqSxt8
zIJFU6BfUZyxOOX0/o98TRLS3dn3g9roQRFpM8Azpb6X1AV7VTJMdoZno3YjXLxwqYk4ULAVlXZh
fSXVUgYExgD2JqubfuaR8FSiYF+dVGry8wj54LpMobLcQz8EJ9FqkA6aAdpP4FQ2EuFMYAkEye0q
gkHjjoWvxuDLJFhTDtN2zwm+1SUnlM+/JMj2DRiqEeA6yTB9H8IsnTWdqOHtJPSvM91PV+l2absH
D38Q7nKV2bZMmben5Wqq+x+X7QrzriaLKag6+lnJ114SfqER0NpWMRWi2DkODxVCj2kV6RtWJuRz
9xrNoFqr2ZLrTXLXKYyjsWVk0Oco0tQcvy9fcMn5Xnzfftxo4aOYdey2hupakP5u+YZBRnT9f3IL
F9rfqXmP0/WDdFIdIFCeo+d7RW+QsRKsczEKglhUG3SAGfe6R/ibvxM2IQYUnq/3dNxI9KL/uZTG
Iv5bDWYnOJzXtKAuiKWI0U+yPq/ezSn67f2hTyOcUBJh5VvmQiwydWFUwsJ3HbccLVDyeXPmFSj/
r8WHyMlKLj0CKDVjNvKX/NhX9MN9jvruTtJwXkb5FTW2P9CG4X21RIJyVeBSd7A6z+TdCQz7y7iX
K+cvxDchzxJruU3GO8IW7YXPynVXxakv2NHCTNqR4PMA7psMeHCV6ndLnlOyyMFT9Nr54wGAAiYC
XkpcW+EIem53WBQYT8sXnPBShUOn39zT9DZZeTJMqUv+Fua3yqKqZHeUEnUubv5+50PcMMzaZ8FJ
Tngx4dGCBIyTNADZ5EHr6jExfE28Qe8EQzQLbAtlJ7kGA2UcOvCVSfK6y8Jap7WIKiRVSV6M4oNj
2bYNy+Nr4ka2CWcjEd5uL7DkWuRRWs6K+MmubS2WkS6Fy9OaIttcQQ2WoRO5V/2kgOjaHMS/iLCE
P2GQx6CZIDxk4ZGhmP9zWxcmEteWY3RGKxm5T6ZueiEwEcGOqP7XBbYnhdfusNhWwPX/9ohtTBhZ
D+KOilbeO6BLvKWrDrKJFKoYvILaXSN0G6cGul7kEKw8A+lWAKZXcunJzHT1HczJEc908bFR5x4u
j0KUwv9i1aUtclTzKKCP1bEursx7IVSOhkRFF1tmUVymMNWkS+RxhGcNIx9mc+CMnjlv0ioThnEE
pf1/qNq9HpF2uwK1W01YtSGbwFrfM3X/0iZA3M0T7t8aaCRuPG8ynkNDBKGloRjR+gRthVQh0AiP
1LjK7gPuMTV7UDS9ytF7SaY3I9eEX/PgfrI07lqB6OCLsVy1EA9bQCCtzeXEIUm1a52zOabN0uDl
7w8CZGWnZKZAO9/pSxIZFCOqQ4pwfxTbEw1gVeq5KtjnwDjBXvSd36FJvjGmqGc62dn/d1Bc8Sg6
fQd7uJY8i809SuGKQr8/WrhU6soPq4zUITJCmxsJogY/p2y5E+/oDJofZ5OOStczYgD3mq3ke3GM
BmbVK4gr6kFaOtq5PgcmxtPzv8jv4t6W9P67+Z2ZUj9rCXDB157rqKwR06va4mLOksL/vkphhiMA
E4ShJ48IDD2igupMYQNLD/XK8YCgyeuMlbEEHDiteCzSrFCrT25Njar5hYDVx7B9SyGIjUUBxf7T
guVDZufRtMNtf9Vij/DeT93KlDuuV9bg1DuIaf6gKKuHoR/63hP4/A9MX9M14P3nohi1bIoUoFRM
Kd2DzDydVfdxP1GFM6eTW1hNH6EYLR8nNKhaYhk5RokUjIE/puUhFLxsFDtSa+oTNOov8SRyqMKF
YpJqF57beZveuJG7/HK8G73AQO+0CZAOMQzRMSpjNvJNU5YTn2037rWBMUNIYDWdu0YmzBoHyl7T
IwEu5OwsEt7dfRvwnNJ7BZKMW0IrmculwiuR4jOR4m13dOhOmDxOZNhfLBQm+R55DzbSz9+TkvaY
hQb6cUVgLn26yJ8tZcENFkSTiL8dlqPaNc432eFU4dtItzZgwNJ1592+2TtXolKuwWCwRulYnFVs
7bsV7CW43ZIiC31vElMKilJYGuNTSbupGNQcT1uiq0yPQs5nmN31lpe/0MmiJJ+l/GfGFK48cfJL
Cr7XZRbzMnbmas2uEbxFHd4n799wJ5P0wg0SdQ/icQOKYTyF4VZZ08mVvHYZCwzftVRT3FM3ww6t
S1NS1AW9mo5Fgr0nb7UIq+zf7UxScCl7PLRkiJzoAMfQ5cvYQLaVn1c7nV8uFC1+wz0MnwlkRpwo
nw03oZvKGHGIknwDrmkgRztrZeJSRnFvSI+Jpl1UcETtz3wsMDHYGv3ryDvM7T949wNi+nVKA6nH
aOlSW0uEUrdH3poFZ3g9K6Ntx56AHebN/tfGxmR+Ir5OTYSAZTxXNUPhLXZq4HSUVqSY7lOMNKI7
1SUddfanCUc/h6jxCFZEtVoDEEZ/vd+wJYjtR0NgX4+0mXA23BYyYCyCauZr+DJPUOoO9uu6ohqe
gBPsFNuu+XAo2qqtPNkLxBaaVD5SVAM7Sk+QMwV3PLaN42Flu2irUYIlNfZL61OcvFdzJ+Kp6fA7
nxoQnFg5KDFrR92F+HvU2bEDuCQ+fICNpSYKXCBSn+xiJMXJ5pC23Dpaj4PgqFdNvSp8j30m4BML
Y8Z2qVd/bqeCpbO8jjd5Yr9fVpp/2AAOWvY1nmFoicVdxytTnb91Q3Oena19IV+lQiXtWsDebsvJ
aPiCjtHUjVTp62ng98LPoKk0nk2bnKF4DVfaigqXb3A3AS47S3I6zs8AnTc9zSZh0YdstZzdejT2
gd53YGlscFlEuoSVzy9OWO6wNHITov5xUvCMBT9DwXfxExVbcVwwNYWW+a6KeUI1BmqIkAEyU3iQ
lbBaDPx+CKY7EwYKG/6ls7AdtukpAjcBFqS0zkDyXZyCmoAX0gIbfg311IDQN6cYuXDr1p9KIb73
yCNX0sSTgPLccLt1oEGpc0F0WXBBAHMzrq/HcpUm8JyZVgd5TaiTLGRn2Td+pNAN8Xck0vECcgks
spD6kjfoYytSaanOLNwdyz94znFlWXKgn21qo2vUhQgeoi7pKuoZlBWKR4IpNrpPGs88JeUVjLWk
S+Lspq8vrVUN58IsjGmvC+pm2p9VqNLPwT1lR0ZkCOTJjsBNI6F9yxwq0SKBQUgo+YNuXgQBdy92
DCCwzD0r2zykRn6WjIT3jXPX2zEf5iL/jTbsz02N9Kk1cnwXnQXFWZ1PvlGQSxRspPS8Kand1q4q
JgkliGC+BRJGxfxPxH1DicOXZf2CCka79GO2RdZT25+MQfmMaMAWJ1V7oPJfCLQU1m5flzx4a+jq
iI0pK1yDRmiPd9F0hgqE/v5BwlxdAfluxA2V8DmKNJv71PsbBIkS6yXG00m+XQ2QWUOKblTGtdtj
BeV4xx0kYHJf9PqqFbQhiRgVVmpgfhOzUIa7wekdYcMSBnTbGBEVe/9Q0uymZ+MxMqvpOfi/HJXY
HZfTFN8M23O47gC0wll7BvPpSicBWAVxeCrMBFbQDl0tk/pwd7w7LoqiOw2BL2OPeEa2cQAjcbGz
JhqQBC78iCays4oyMju1jWRwXFMCKCGBRu84liB+WbgCZUQgnw/QtjzCC3F/NKF37eLH6Vmlwxux
tJzQltLXki+qdxWHXiqkWEr1HqfpicXn97vF99ZNcDToSkYb1D8hlU9g/FsounmjKc7bE+3ddywi
J6Lhr/Vw3BbYER2LnHHly5AX53niyN4z7ZJufetsvwBZ71et8mqIFd7tDzJvWDnfDu5UqoeQO+/a
04JLuIS+57IXn6UCpxZ8v5EJUI3RI9m73BvmrfSlfzog4RYYxLzXoVoVeJVTsr6ruzx64lvoVShw
P6bS0A7HUu39xx76zRXpt+dGzmYs0o2V7vVo9Kv9oLQ2vkncV8iIgPrYogSMvpZh2BZKI//QPpKJ
bPiIuAvOyLQY4r7kT8aTaDRptzoev9HAU3mC+OWloHTucRquqFzmHrIGoZITRXD4MXES2Ig7f3Mu
AgMqZkQEW9ptp1ntGT5wFCZWszkjwFBCmwsWVvxl/gKi9WDTqECFR0E4BwMmQ1qnzOTYR5mcn+Ax
PojORqpxfMXQzoHyTnO2xnLUc2MF+gNSe+fEYTDe7eNTmoftQKr2CzYLGzDJ9ociagaSLrtCJCVw
fA9FINDo8KwurNmSy+XkmXoGfkFAMkeKFOWBimTVQdZ4DchnmqEa7xD0DJlLXkG4///ExEx907j/
7vqevL4YtW46ytsjdxhl5aycY8TUPdWBl6WdxGnSUrPunxUpB/fE8HpxhTOIpBYh9rw3aFOfKTgv
8oInVfcFJpq9atlQO265iO+PaqefIFSkFkKY8IRk3Q80YV5wS2ell1+k7+laTdOaM/NFdYjJ1QE0
DSExxzYL3MlCJVSoTBuebSSxNLkFAdstaCdOXuz3TatCE+U6f7taEsdLw8HONYiiZkz60yB5NdA+
++eU69/faxYh0C3su/Ji/O7LNoF+b5/ADUpM35WWx+U0DTaVmKb7xlPrzVvW3F8b5CpE52ZUiPmB
xxR1nVW1PQU5xJL3GSVltV0cAFtYeXxw7FIxGMCz0K40bHOOxPQJCqdHummNJX1QZuKl/TiOjTZ3
p9TQ9A7lLF3EJnCJKLbLYBXRd4zA9t3DPan9d0KWoOJH9Vt7Am9nmHi2VXQqx01joWew8+Uz1yg/
MgZ18WfIutNy57CAl1PnZUEj5sJRDKJyXNU7BJc9q1UMReXEZ1qPCtYibCoQwdMG8a+lCVmGl/4p
v+aHbMWbGTcWPcWWaGcYqyX7wYY1IYYLFff1j8bHIkH3o5up5h7lSbhjC6xeMJet39sNSxOGh/7S
l4+qGLt4IE/iBIcE4+W+ipa6bDXzPwxUb2DQ1lNjjcskFEaocIuRIPiIE+7TVZuCCiYc6jvmyT5q
q7poCRi+lcfti+dmBQpWkStgUKWR1c8+RCoQPadLhiSD4fzVPhn2WYfOJ1SX4dXdPz3Is5tAdtIC
EVdUYto2I4EFTTZMUx3tmFEalllF5awpYZS+CYTqL07TSR+wvpVl6pyXFqONPNy1Wx7JpTMHyzGC
tSeDDvBufSXa34haPjPqvKQtK+JHqOvFku7BuIoG0lC8G5wXB7muoPYiLKRkkOCmqEH1omWyPo8X
fyAyWZr1FDL8OtMmj5vKvnSbtlvEnDQqBWwvC8sjmR22fxsN+ft5y8ju/t+UEj6R7N9kp1yPrB/d
5yRxim9yu8SuCKoN/eiL467i1nCZ5BHHYVbZv0PZYUEVBmf196nOZBmBSu35o0lz46QQ1856Z9cQ
0Fxzm9jSm4AJT6bH+zsFcbC4I5TCsV72D7/d/RyM7Nm/Gq9T/RzJUXYX8D8qrkIilZOSt8p571lo
hwSYh3nLLHkDMO6nMYk6Z4+tZinJ0hQbPEWYPDv5PC55UtVSIr9W/w2LjOq3XwUMdOQAqVa2wwXa
CoKZoeasNyYcY6b+zHfc9VezWjcXwAxpb4xzuLJuGdwoidAUyNii2KOJHOEbgdGlioYphe7vKBNY
2DK2BzA4QtPHjFR6VnD1Hp2diwOxu/4EXkiTute3MXK/oAz7ayCsZBRtUZAQOXZXtG1v51uG4+g3
tQ8R9WzxAR51CEK7dWl94avbUk6veSDswOCsYnJy6CIbtZRsyh0ir04YWWGTPHLi3oGSD8pD6NAz
4WnLBVh3z5NISMaTy3SGfG+1UzKH/+Aa4yh5IIYkP4AUCV6SiRusDHwDaxu5dmFfExWBeKS++ZPl
fBYA6+HiIA+vHByUFoBzx+bwlzDbPI0waxvphjB7PtyIE56OVjpre8n7SzAT7gsj5WZ+7mB7lDz5
ucSqeKCqsNVITJ8ADPTp+mE7W6NgN6ET6H8jjNWtBJoCHXYva1iAYDjExmgJq4YydmvOc2lNaP4b
HwgrYJuCfcSdSegdOBiIskw6FAuURMVtpcq7jJUy+2OMbej+xkrVoNqeI5mLF0exrXfcy+aW4DXP
oaZ0i6h6rdU0n40EH0JTKMFsiRLJtaDm6QcJhiRs4kYU2+UwyaScxvwsQ+Oxx5dfngbq1oe3f2ZM
mKTT+TXVROulogZXBxdEyfgIFoh/XcWEMVFG86T9dwRGZTamu4E5j7bRvjx+lt74v0z0MP+MmNFX
Eriaq54vk3j4N8fZnC7iss7WLEM68YYGoZlC+osFHEcwe8nGNl8BkPzqfakijcO4tJz7FWSrJTU/
w1HHyOYRXfxcisVsaHclOW9LCJuWApwkqv36IFiQrwzc5s79Ipc3rDvRBw2WKTjDUTHq4xUqXU2o
Hekt46M8gD6hV9Kwa+gNm3UTFETl7A8zmYM6iRIialqNpm9i9FBqsuPh9kOXBar3FXKc1VxwdrfE
axOYzpgiVQGo1UbBFfYjGnBY++AynYeEm24W4QgC+XftVtynTAJvpR4zkC8o6Md3Q5U5qU4QixUi
csrypN/GYysS9eWb3BO3rLPZcQZOUymJnJHVBXpvwTULJ5200Y/Wxn55Tt5vl4GfPzGAOGCzsDpI
E1iXRh7YeXZa7hDSFk35xByQy0oqXFajq8f7HCdOkQBHNCjGcuoNWkzQUEEJGKNSKjxyhc09Af5e
FP6L0xjr2ChXGHH4ii4hhXBLsYUDnajIV7FhwL4qeZxxZTUHnNf1ReNyRcSqjFH+2p/qRKMPEHvZ
i5llx5IkInAHzZFuw4PZPruQVV+E6JYqDm8sOhZG2jzCLGv+7YHAzITX4N5QrMvjHenziXIzMnhn
PhGfEAouzsJNShDE/DV3+X3v6kehrf2EcjPlqnr9AaFTHbK+FMoF4bAqsYKO8HSGfoaD0GHbZj2R
lFm/XfSMX8rjTIC0zkKJztQjaoHrMz0FKRWmTcoNfeWee5yvCTjr7rSoGkzZBZ3FdspNoY8mRiiP
GOLh/A1NHkE8zU3i0v5SONIeFlGYYoRG873vDSdYDJXrt7z4AeZKnkuZGWvwtke0BNAUdPRDEZNw
uqReKzm+yFOapUiONDojpSKxmrLmNSz1qcLtOwtYKd1hUea+wQi1UZ6AHa8mEFiG12gFRfm6nK3m
6fyKfUR2iem8GiAzfJE6WYHRcucIDYZfLm0EcFCLdoiix72vZBR0DIYc3dLAXx/+2HZnYnJJL8uD
ZOFv5M9axC49XVuE5WFNFEzGrRhRdBb5LWvFx3mYR/QiKFn1tpenwh4yMbq0U9BhdpFnvr3NILHC
1VAdctgTwSWCQaGJdu9gwtzCKcTYg240ZDTMR84G4dypjwnLo3cr+3KPU1V7pbvA0g7/nAJ/so64
OhfK3boYw7QoqPQ3kQse/1YE9QM9a9KfJslJFh/hYaHhY896BmoX2+buqL8GV0G8gd0t+20neLmu
dNBXCH6bq00CU+2rqcaUYgvVuxFmK6R6Zb7QeLyid+j2MGTl76jZ0XLviZ3Br6nyyarvf0MN5ULQ
YAOWR2EWva68v6RfthUDkG0KL9GCDdihWVoJbSIPaVktEKvVnYnQzsiBBJVpZuQi2lszkGox1rKd
5HQ5hQXO8++K/XRfc13U3rtvfgrhaIjRTk7vWWXvn4+4Rx2A3slu1BWnkV4EVbrEVmGQCPVMJsaI
O0mxDIAYZ6EMLG71bdBm8AohOxSSAx7CUMQOFT6DZD1lYrhXLnZ7JNpqNNgyZOS7NnQbqagpKwWW
L7IBHFZaESBCuzTg1mma0R7jcsuSFJEvra/gim7eRacBJbT2JibLb498qIfBCwnq24fcSIbPAbVZ
pzScLp/ksCYLeo9Cp8Fb1iztVrpv86hJtMci1f61QEjF5sdTMETJrZN7hizTn9EvVf2znOToZk3D
k27UywEh0+TwOHADCg7QtBlEd6n6AZx4LspyNvH/1onsbYqMXRB++udTh18o8+lWrEnnwKVHiZrk
JcsV0Wgidr1hdyoeW34cPg+Iis8p4a+vCtKMDgKXqJYl14bzuTbI3z19xLoKfydFT2l5QgNSoQz4
dh24AyFWp1XUiZh8ThzEk2Risx/kc5rNGF/74TsalZLupYVEZMM6yhXjUdTtMpzX8lCAAmLCiT5c
CEKKIJ/dOZ9Yq2xZ1okLFEgV6xHzwZgL7sQ8fhQNuX0CCOZ6E1NQDMVsoU0VnmTMd/HdZyNoQOnS
mNdA6MWFRlNWRdCtG4zC9ntTEkE4bXxSzzY9f8BoktkCtFms6P8kGcXCDAFBfCB87KjaO2bYudzI
ik4PE/O27sin18797OPa5GAhGmcz0aiTJzGDbZscho6Ypkk1ltCi4d6VSt3Tls5mTngUgBQ7EYIt
bFdF29MEmRnc7q3uMJxoDiWOMpgDLcDIIVkXzC97VybHUsNGu4rRbMZ1S30gzsAyJc5C5yoJadgU
gdI90YdC+bFQGSUpwtxNqAXgKdsFSBC9TN2Cd+bhZDGUgy1IDU69BGPfWi917MbXuTaHoTVzJ3PW
sni6hvDdjguRdhLcv/mD6GacZjtFT3XGPksPcIfZ+xbK1uEffEoAuiRSHBYps6yruHqIB1NEBmYW
AT7siPSwPRoIya+tp2bsU9rLI4Tbh1uLB1G5+/ipkiDeuRdYog4D3VV6rOV0a7NOYAo/ol037xxZ
CJs918f6DEPn7iX9Ef60da1Ehny0IJ4Q0s9hRrZybayVmtYohxljyCgfTl55P+QEuweIH5r/O3Dl
6r50xyoCokUPI2QOwJ5fuj1s+bvf3RO56pIB5aGoWtzNldRNYPnA0rjAoGbOSwLCpoQM3JYJUEOH
LfvgEf9yS6gXIcPvvkG/Rd6vdmKl6uWTiR3/zR1udMxNmFUenOBAf67iSyIQD9pL79iIaO94cJhE
8ik1lI7ZpodrmqHWJ4dOwbgQjv8JYn6wGsSbk/vBb2xqXE6BfO3lgeuX3V2i+ZJp5/y84K7xLoRr
IMRdfvqAVowwnTEYP1yVqQl8PYjM2vgVaHalk0fGM3cFZfmXT0a7ZSdPTEsdPRlaUY/FLGmZ/jek
plKCo02IohHLVVUosBp6IRvOfp3zQ8mbxBm7AJiE+YgxI8chqfw4TTcJkUNaFAXv2+VWkdXCpyOF
VMcRI2FCni8xB7HXf7z3PnJqoEqFOoIiIYTE0JX8HvvmZuTxg4RFI/UFcZ1EsUoZ6kBVNSwZJGe2
rmZWhQDwz+p8tMrHiS8z3MNAIIHfV3vQH7U4dyhIsbLbAmjMYZf5s4pPEZSWuy0Au9nipQmXDlXx
OmVvcZR23QZOc/MLw61BykQehiaPx+A57R2UA+9w9rylAZx6NWUboItxeD87xYzWdFQgAS1urIRR
EDeemq4B7QxZotFvA2D1KGLSXBgDXgnNSXL0DNPdgKYasNP0Pt01QePgZjRXksh06VjZzPm/g2fH
CKOszQ82zJ3JdW+4dcRvQ1ftXWGm3hhaLhRDjgi2qR38x1JgSNWBQrS7YvyI1Py9jl5aB4HJ5oW3
jgJItCdaLSzdN3wixQ4lP7TcGnJhkE15tpx5UwmFB12Xf5W5na2UtjsDHVPtT4F6oomq0/hrvk+x
HTOxuTE3xVlqoxBU1TcMZO6tfRDVDaxUbnstzKxJVGQIDwRePAGPlVwE2cLNZC6niTRzg7w4LSHk
QcHQep5klcru9mm+t1WDfogtHaVqMwxILYv0TLj+4CAWbhZvHCHFUqaX3naeZXCwES1Ajrt6vJbI
KC4cbxM6f55rK7w5aPYSlbPRCIO8RWapuJgqgU6v6OBGyWapi4IHkBUKe2FDl/sOUj2Vang8d6f4
AIDez3Ev3Jq5luXpouD+KnylCPK/ZN2Oj0TlQC4e63wdaf+XzqIP73OG/lmTDo+yqDbVTRp4La6j
2+tms7ce5rpJ9cnNOBCrzNH7QtdlMKJcav8ykMW7qhb0g2vKDchh0u7IIWsD2LGIq7QxBA1Djo0V
FOLrOW3Uxk/RIvIkQAgDO2/ihyjXR552xC1DVhvRGGVwkvo4lDILpJuPLAsR1ljQQZ/R0UStMIeo
85o3dl2pKgd4S2yt3D4Bvp0fk40RyFuFMNlKhER6Gh43GX5UxGIBlMRjzVyDoYHWwxAP63qlweXi
K1xdBDfNTwAi/LybEhfshRKwrLA2CX/Gje14Qc7CuORJYPj1h728oDnvZWCe/Sgd+eccW75Y5JK2
Q3QDZrG+lsQr6FlMHTpRpuv9gfbVQCxFtYB5iH7yDrmATr/w/GtjnyQMBXveXucEUajTibVp2SFr
VQAkCj6gLuho8aJJ6y8vkJPzbDSUxVJH5a6EbQW5bz7UwH3GL1R9NBoEQ0UJ8grK2JlilZJvQMu1
d6o0s5FWRWavYoeA29Mfu58Jls6JoZCItcwlD5IBd5c8LivjuQyXSCp/jobO8pYUuFSRm5SkYoZ/
HyMmO7CV4TCrq753zn+gYdMxvNAPbMqoG22tS5OnALJkg9giSsSiA4TAfj+RndE3ap6aurdVbWSx
SrHXzu+LXsXwjr3516zwfem8C255dpU9XKDjYsssDW4/skHfLNcZpAtDDAplL6qHPSvUPTM6Y3Vd
UfElkJorq5apr4CrVd8V6RIdajy7mrIUAPnnd8THOD5VdGqGvXC8DTO49VKqKrc7IJO/j5FvpQub
iyZZ5B9K7EUpxdixfG9bwNsULT+ELc3TduK9lhaBnoqTqgeDGSB7J4AKvpPAcjlUzMyUau9djUA2
O2g+Ai8S5IYfK1SeU5epWTIaceddHurcTRmj3Y31im2QQatElPGzkpCPUzRKmraMz2qGScAQ3zb/
H7GCZ2JsjJvnZypYJhnzjrkViPcMpreMv6egpoons6GxF+y0QxYfRGj9pvbY2lHME3uqCC3VRCZD
IOwGu0uJLmfuiTiSL2x8S3TfNHxuyev5Si21cVFnuzlrJSrE5yvUo6oIUtZ3E16KfS5h3EvEFz3x
x90UkoJx92bsqKF3FxWq0TPak+Z5cVMmGIwrZSAtkeVh4wyhXZOB8YVEBrSFEEkKe4EawNV98dQl
6nMfkXGndNblW7TzFqUrZLUoZCxdkJO/3mj8sER6iWXKn2bEiGTFbQlpn3RfbjGCM3ZiME0nmIEc
gkWN7u2tElHDLck3OF/YVFFkUDlmSQ3HaZP3jOHxDycseDc9SGrfmFFzGlPDW746GZf3a5LY29fx
6MgCvoVkCxPM8US8lm/phmmacnYxi4vzaDHlJXV6q9n4EPdheAp3/UI3P95QxfDxC4u919O0SrUv
wzSDms7pgAiIlFtZGLCT3dLgidMFTpm7dq0xTqNy/qMMW6Uz4xmlaBclSFVkoDAhUXGCQKiTocfH
CFRRj2kyg7pEP8qWEeEnQPzVdPqJM5u5ZF/eidjq/71qbrtB1Wqk1Yt01/rIOK8zqC2DDcVMTsws
+rgcVimZJ1Q+RxiSlida8yREcXl1Yz0pNuhD04ElmCPlZXg5UlnD35U1IRR30PpeYxECDQhtEDQ6
GKWSdAumITyWDCpkfVY4OEuOxwWjYg1q4Bt3dKJ0Vtl2kWZEfBota9/+/6qLzaIdoTqggyW513RS
6ThujSiGf9DAiA8StFPOFNWa0kviAJ1nXgY28yHTrcohj+D2wQP9xeNQG6BflfgHUSmMXVOpc5AH
WO2ELITxy8+ogfsW68auxxDphkiA8RI2uoDNruSzNn2Vw2UwFQeTs1TTPCqHshSCuc10gfY7cP3m
W9g/Kj7fsDYT9zRiLTNVrVX5emYcJJyNFswWWYWbhMz43ores0x2n+x2uWnIHSTKmaKHfmZP+BDy
sSF8CqaFlNkSCcQWC+spIW2xHaa2KgnEnxUAa832UIU++scMG/uekqdHc5reqxHqMpHMVsFA2Peg
wfopzsgitQm79FOtkomLvbZtCp+xTntM2VrlFA2KeTN0es4RjyGFYJRFa3U2KIdDkG8GffZqXfnJ
gijFRSim0AtVScNoo3onaELlSyZC4ITsvnbnNjizX0Hbwp9M3kP3ccblvMoz59p2vnkatCzthD1M
7c22HYH5cW5QXUE/5F/3FqM/GzakIfkh+GksMyxuc9mu2gAuiSHymeENgaBEQ2mRx0T2decr5xaZ
vGvHzMdVL0PvL2An/mK+RhpBk9pzzXksr1UTz+T3ccNkGtUlKgJtpdX5AVrto+icquBsi9zWOOyF
V2VHtLLjt/jE1IkZx2MhH0N9F+mKu1ySuXl3/GFcSCa/GQLV0Xmxxj5UmKzoY3b7PPoCgC95Hou1
PmJBRwUiQUZWpP8/pEK7Sn6G7aF1HjFhPkHPkR3iibAUZfLOiuoFTYz96siimcrQJ0CSC0Nrg3jR
KvWRI53Y8YPVJqLyaTXSfGczNYirualYFqE0oAkICDSUtTuqmXQ96Y37VVzPviqrRC7Otuon3T79
e6L9QzdwkXJValMLL7ZQOu6R+HnX/4BUn/uAzuqrCJjSFcB/HvjGDCQ1JtSXjvKyf1Vxb/3G70uB
I1+Wy4NnqssA9g1CE4FjCgthaZYxPZVHsFmXNF5X+bS0te0KUisfk0+/db2ZX7fEMCcwN2oNO8rt
x0PYgk6Xt7j5aVSgczo0AERW5M5X+RmB5onIytpcWvOb5iCJSmtBhKT8Lo4AbZi2mV+8Z24B1Ogv
djZN01ngYgQvCaxSDlg+vpXThQ5TIvVhOo2DM+Om1fZEQt9VmNnTLwh+2YJgSMqs43J2bJNZs0jz
5ovdrX/VABdZvYhlJ/JFY33WUEJ3mDVKRzWzNYosQcw993XJur3LWns/4yEQRVADzOIVFiBKgvsx
vMTMwqkfMXuievSV9W8suMfIxmT5xmNLHSC5mmVCkZPd5HKsc5ICuxmsTyPKTuML8kRLFulC281K
8X+tZEBG4wNjSyvPuy3w3gtSwrD+GxzDSY8dJk7U9F4Jdhig8YIYaedWX5KkVb3J5fKm/EMyFtX0
NwhPu6nqyeK0/c2Qu9FN/VeL9bVTJBDLv6a5o0npynx9wHf1ofb38dC2Wk3TtIGYeziAjdJeVeHp
GZNeA6XjKL8gDkQshWtl35QzoYXVSin0SQdeR/djqctKkqoEDIpybMMXxdHm8sMMPVFoM1CmkiGf
+MzrW4BK6LVsp7RNKY7iF6t8DW+VML3H3xrssqScNsdZYNNAVF03bIWRHLwpxQh/w26bE6mxdIan
GTGmd4djwBBcQyER4IziGwig1vk1gzwKVD2uRzXVR4/UoYYW5gtTxNiKW88z9Ly5JVUeH8l3nMom
WdKSFpK/hgZBgmIqsaN1bFsa+OJPO/uvTA15Rkvtt9Z32mrBJo7O8JMQZlFaT9Ez1gyoHRbzqv3g
XN7RuBZawZyvL1e7aDvNVXxmEWJwO9zMZe4Qk7r7m5T+RqryKNtkxNlvEifCDkgrtV4oD8xh0oMM
wcBhOJHt20kc8uH2svPyvuDUqau3OVl4NfB0IRlclhmTuJeQNBYq/8oLSTU/bKALmZ2u/d1vjLWD
k6e7RtRIx4bvgRMbePW/wxNH+Afd2ZzVgHnc4vnWByUVYplF2Oi67qlyWbmwec2ICyCp2hqvfUk4
7NyUMqEa5stud8EpyK4tTxuaMSZEevd9Zmvvpw2RIuKYEVKyju2x6vMDXD4CnTb3Ie7ymcABd3DU
wrTQIb2jTBD9F6rjwpxn0JmPXdtaibDprlZH2hIZgBKp4BfCSVSK
`protect end_protected
