`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
kesOF/CVNHwXzaV8IxH0xY+lJTfYlkoqKdnzLcdHZI9PwZkVdX6DU9rIj1nQPo6Z6FbwongTSHot
O0JhvQCulYv4PQWSTc3pptlAk/JY7Z6GifDOT48XNhyVXkVyAjTB/MhhddoJpMNHJDVJZaO3T7/B
KIcZNJTBQ2/3KLS4/d3Vn9T4jkhz55ibkU9wMBxdRchUEBLe/TKLPoQAazRZ6ajj3UlcEqdoPQzs
lR6uya/7XrY3Wk5xQEH8m6b6iWNMGR7O5c8ssdEV9TlF/b7LVctlnP8qPgI3A++qCnO3fG6XbvOR
GNl3u/59yIPY/+V+NECDSIuL9FN4oJx3Owbklg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="zGgYeTHCf3Gc+CvXnXUTF+rWv3PmKL1wPbsJqV5mtK0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54560)
`protect data_block
9sNfUXJFK+3d/SR+dxKwz31TxbJlK1I86NccXsNktOQrpqqvelRJ16KxXbu/mrgpx+bWnZOEHYr3
0sVNtIqQsLXfn31iwI2oqwGjG9Z9de3HwupJE23qJwinmoS2lETNigrDFH0lxf9QDhWM5+Lxl9ka
cssQ9ZXrBXvjS2n0827iNF6Arl1FcCgZqpMUe0wrHiHJy2z5NfRlUeXgHgem70/YfnKMy1O2b79Y
6smM99hLuEoa/PN4OZZcsAp2iv1782mGouRXheAn9xiCdmb+aK0obkjrqGkFzIjNQuIe5M46habk
j4gZyMIw3mUCxVOirsHnf9+Mo2zwRhsL/tSFUDeTIgXjCIdaW8D2vVDwIofrnos3J7m5wpPimHSw
C3S824Cu0OJwzY8olJbEHwao4htKVvpIMS70p/Ye6BNvX/RH9CVcJvl6RYJxQBsP4d8xqMH1+53Q
NOG9sA+GzwGs/RMFqpzIlfGZGpuxctNVgXBZ3bljTKXWXonActCWdt/LVQDZx/3/g/figCbWuW2W
rJq2fPuPOt7q3XvTFeBI35oqOAtSerHSOm1RKO8VVIFmLLQ90pD5OLXL0VGSrZN9n685jHTRn8cH
QgEyxYywFB1j3PMHsruXWUAVsUjrk78ttNb30z+oEKA1SYNSWHi5MBpgT8SHZvxvlLf6jb7NQQC7
FyvX3+nA0Nms0IaXSbdWif1ctzD2p1k4Tdw7MJe+A6hW1fRuYoDhnNuLzUsMSkujpIaWvIEZdkep
cvb+3wYR0z3amGcsmPGP4+SuUy6/a931hrASwece541lUFOWkn5EWlSq3uUKZM3dmE1csWBtAfPd
LHfiOghT7wh6zDWLXF/qNMdXcy20Vtz/UMlolAJmBFd87ucIQfmslHaKweV7YHxnahPI20/C0Vz8
ABDY62MlG0gRvBiWvOj+8Fk8EKURbMPW6nSkxKEC27qceai3hsVXWjdjAe1jOjAwzBXLk1WyF2yL
cuaiHzKxNsCOSNgwk3Dn89F5rNeTs5xoigWop3ITSDap78G3THfoCJ2qQUsAbFNXdaqyMy5sEmx7
Ha3mKUADOB4IUok8Sz1v0QpRnNf1AkkMgZci0eDN29iGTAM6+w0VplDN/L16i+fSwGc6osY7WuwW
LvxwGmFgrLVc0ldVAhStRl/Z1OutQMh3d1bnwfPZyfRGEPzvORubxIn9vXpdoE5bbggR7We6FIb9
2YGBr+0KkpGE/HQZNN9SPHNE/Okzy3zjMSuBWoowizQVg6aTKMwMBcHL+pHVez0NhX00ZW0GRS83
IPW3moOs4UWK03smNIdygKvm84Mw2y1jOgbfdz+FQ7A44QZJ6QbhZSBGmvyGISefIWt6mg9zeVA8
e+Uy6YjL9PQYR9lTb2TRJwuQ7ci8CoQjayjqcVeS9SRI2ACeDHxoP8jXYeOpzeZQSGoNFXhzxQTG
QidhrnUwe18BWHzrl0lJW5ienCBjXLeefEGTL54kXZCNsjLKUGDirPAGf4cJ9GvGebBuYycdFO16
tTzbLsBhKCSbbVsvi6zR6ZW4b8QOFasIGwKCAWe9VoeLsLDTAhMAofTE2Vvvn99IJPsQlQ026uqW
RsQslqEoyozmOT1n8vTi/QLe0q0zJzLhDJLg1wTHAGvJ5WZWcmsXCTHvSQsLii4g7GzKzadck641
ibezepamFUQqYa14e3gQuFe9zskwGXskGtp48ioHXWZ+loxOAbQigNYMsSxFmtTmK8ukcqsKRUuF
vxv9RFOCHfIzRDjarcS4PbSk0p8OKgPnGwUfd8Wv6QKMU+Uy8ogS2uYUnDizmU0WzRWM3OtZgprD
d8M3s6Nja6tYx8w1gO3NRwDTqsf3GmZttkhj4Rc9zc/l15HD6xTK8R9iIh4bjlNTBPy9lx06Kv2J
q40J//Cg9apf4N6UH/78BdEgEUvfWBQ/hXkUW7vklHO6kE5sIgxpxuz0d8k3fVAFP1WyZj379Rtx
1dWNNIgy0toeRTotDa6CrSume1Sjod5Uq3I2pQFl446tvLR8Cc9OblUPXJ7A75VTl85JUCvhwDNh
OHzkbGtSmpjlZilvRdUgFlG2Ws8NBQTlu2UITCcfboCVoNHEuyJMlAL86M/etzPkWInfA/8PKVVN
IGrzB/gX/wIkK0UxEdt2xqSrnKpqHHBmBijzAqQ5sXRLTH5d+VVzs4GNMa4UL27s+BlYYFOKg65H
J6dOjjlQ2slxjc3Ofvf21gUuyWHYKG2zBO0RitX3f+HPpl7AsPEYE44htuqqsnebH1+28qks3dFM
AsdbCuyyWWqHR1KApmqnbbDZnjaClY8O0yYHxV2anIzCD909QDsDErOFgqrXu3GZJOwQEh25Wh0+
8WoOC0yhR+nOnIagyWodUhKfTNYKrbrfrR5DbmUDTL8HrHS3ZESxyNsFqfkRwTsHJc18XbRoUHr+
jHeMg/XnFQyRvQZP/Fx7MfhgCWyU8eO4aHB6wPzFuE3p2vqotrjJDNJ4nfUCMeHuvrb+0hnro4Z0
xuSzSP0q5KCDyJ8yn+mNn4wlRMj9WbjVrO10UNMHGCMahwiGLIdXPZcoBklf5QbRRVQdyOO+ubY0
n4aeuIGcqP37lL6427pjMv4ztjQDU2ewWb8CkBWEGl9GGHpSZfHCd266HpxTPAjC0e6j8pmO0CyQ
zM8KuQXttCxy8pURP7AptaNqIL0Q1Jljo016aRw3e7UvXyWU/hkFbusLuGCigJOGsk1XkGJlCsSG
AWFN5LPTIlwXwLf1g1uLZW6+F/CtOs7CtjlWV4U4UOoe0uPoMKnDq4UZ+4NUaP9mXYF+aTACH77Q
QfB/fA2CbWKXniqos6ENionW1gmY2dW2HH5edq3KEr4VWR85rXj5SrhmYWsooZbO0wxq7ZhLkwgx
YZhc1xU28zr1OQ3SyLnqjD4CR1pgwR3O6Hqmac9tIyAjaAVFieNvDNhZixDl3ol1Rr1fDMTlqOPD
tr3KX6f3PMhsp5tWm9q5pKU9GGpzO25P6sRhhYKe827AGJF6SWqxVWspIz4X/LJOJ00DyRu/BJtQ
aYZG9vxsSeAdAFWiEO7gwzl3eDqA3IZv0ParJAQfnAmvbCqlZCr7tI7UNLw+KigR2HKEjCSe3iLC
AeE9mRljL1tNvJbN+xsWBA9FWS8nsTlI2o23agSp0WS8eob00q8fJhCNPoBEyoeFm+XZIyHHk18r
Rao0Ke0Qb/9e3iX8p/ZYq0L4fnwvRmRvEQZ0Mp4W8gKH5fiDxxmCy0+ubpRVyHV1HDSpogdLIpQr
heaq4g/8wz1/soAFUJMsv7JozZXCrFl/LGbJDUFUb8pi4JEpw2UyzYxJIT1p42slpdDHGKhgB1gv
aqmiNFmJpKhlK0ggucLkAZn3S3oTlB2jrtn+Yflhff6SoDZvU+aR0bp0kUqQn7vz+4ALPoxz9StJ
hJBXzbEuEQar/ss0WcfkSlf8mLLZQFmx4rvhPz5V08YO0d78U2hkeynsiLfHCsa4XcJHrDtZXnqy
Egz5pbzkG6xDN1iqciY0s1GXA374CilHuGlNDj8zATHlCcUJ8UcxlokKAwz++fZ4YhA+Ozw0z/Py
MHiUOI7eEaQuxbAFsNuu6n7sZqbGQ/rVrwtJEGZN06gff7iEMZYEyDPZA8fOTn+u4mRSvht+fF7o
sZ5Ns9zcJis6vsZgKy+mQyXERWHJES32vsRgvc2+SbSJOy5LWv2/wLpR0uVr5XoNFfLDjGwCgoiJ
wrLbHBP3/PVTYUcmZm3IVPfpt1bVLB30Rm3myWSf+xktv+Ra9WtNM0hXBjuPqrk4Q6gUEuKHWvfy
HZAa9ylUY6P2xzW4t8DiK4sZwRrHCmaKjaYefVNMagrWkGktwNj2sfoEnBZyFcgMXbh+ZwnNNEH7
E0La8CBuefpa6Ob7lCU2FT4E2DUjqB52etrRSpiHujdqmTboOF4qkyAwCPwJAxosUG3RqkYwxQZ8
GxMAjU8Km7Wj9TI2QRTBGAo3UEL2FwowBlnVjlYd+mCqRg5W5g7ut7NMguWuDU8ZE1Kp2oRarHqB
44GEfY3AOFwniXOd79O/29p5LewWB68Go9GN+L/tixJR0Ftx5OBokjsjygxoV1c0N0MYdXqX2bM3
lrrEMhksqcUiMuDPVR9qmvwfdUPr5nAxAPyzk2r0TfILFp9Ia1agid9wGtwOawFUHytqGAGuSIXe
higQTa3qGWeYKHcYPzHsxR5L45U6VCRf1Z/IDsN7tyPIoCFv05vqMFTZp68GPOJeuTiQNT59rFlZ
nouposUmJiNgaLTchnkeBTn+yzRSE3Yp/yD+9qGjyNnPnOdhJQ1jKCxpnK2XcTjuq9RQe3C61Wmz
XJVDwvTnT7YIR626PKFWGlrq7WI3JsyXcXivfiNYxfHPTT4xfMO4CoV/T6bE3QmV4ufyI6JY5gVe
iWErnvqbGJD5gWJ3OkNDmGZTD6NFAr3XwNcszdazq7vBiO70WVG1I6mqgPepFxkyIL4wgOs3DjUp
dzqRQhPlIgdn7QGh7pv8JaEdQ4GQCcAaRVz2NaeSAfupoxA8FyUF2UBwmFszTNmm8bFBQ+D6ZHQF
AAsh6h0BwVRl0mxVpi5iup/BWqkWwhxSv8R4QGmTe6gptpajKS2rLUCH7LpF5lOxa9S9BKVZtKEG
loya1yuL5Nk/ToeLcixioPGHJaeMQhTt+oTKzda5lhIEnmor0a3sl/TYMIltfvZ6BGujkvQMcFFK
T0wgCu1aZ+nle9I2cRK7VHKyEY9YopQx3DzVW2+GopaYIaEnGKWrNtrnHBMpNftzQxG2WDCn0LLf
N09jeojcqx6yZAdjM23Vx1nryLGl5iv0UiKkDXRSW22XkGfmAP8d1OXRBzzYnNkAJc89uzd7+crC
K7+0g3teNrTgeoizjeBzwsmqwvK5vJtkkB1esjhGW1B74zoKuG7IndVBfz2qZJ/gUaXnB88vCTwP
Au/K2TtJRPytsVFOS2z8KCVVKHwfNtcjGph0cYj/afp/3kPH8fN3MW5Xfb57Z0GioChb4L9IpvlG
xAGT/j32ecQ+6nPJ6cLbVUYEAAlIohUvrZXb7xEV/Z+AB9NyRFUdXR+ed4ZyWwMsBhZWmGlozHjc
jUZ1ih2ObyFxMZBdDiL+gsrEjwcfN0CBCv4xcDuh09mQOnsg3xTuVQE74q1apRo+2cyu3/OX/Xre
Qc/F/1zke5SWdC67hWKEWSuUML0Ws2wd5LUZR/2dFsltdrO/dOgfdoHSWx05UoCrhebCgx/DKL0j
Qp8sLUW5VIvZSr2KzCZYZ7gfQW57Z8lrm7ji7hpqVR7EzIGGXJXldPd71buzLm+giIRn9Yikx8KV
Ju5p5HJQN06NYRTxMOpxk2XlVt+aLOI7Y+pFv9CgDl1OFw9ndyoQ1H5O+EecG5OEC19xrqcUdguy
FHOsmN4AKa0717a/31TYHKbg51G442HBs8IpdKP3XTxdpDjF7YIO3B0OSbi5M1YS+9jUoLjuVDtc
276P8RblpbrqmC+vd4f/PRohw2waZuk4zUUWbSGwh33FzchW2qq7uyP0xYwgSkvcWkISs2YTBhyV
hhzMYq1nqsipqdwWaSgQ1pqgcNzpnRWvE2EPAhCp6LJ2lOpojR3C+CktvoQXhwTvw9f7WLyGZ6d5
0mWfJ6WYd1FgzdSLAI4uUXpPo2IalQHf5kTZrtSKZy03FO8zG3PYJ5UpZbz7X3+mHS3eqi4/TF9K
4j74YaIt8owB5fi3oE77yWSOjF6Ab36i8jN/vCaFvO0pYfgdtIE/gDgomrvNa/25F4yQSVCnY931
gkVjKcxciPt99lZ8M62KVsH01JLDufzOmjEDlxsuccwLyItpfkNsYGwQlNchWuHEtKl26JSwj51N
7U5yHC9rAHN4CLlrf1UuPQqoWIggI+Eyp0FFzsnmbWllxADw4lItGWCQJuMcwonYBB40PxAaOv0R
j2jKKGXAODRqAz6Yj04+7ogaQ6kIke8vu+CQzC+jO+4NJQ0oMBKCFyY+QxeL+HcDAcT36QdXeG2Q
lAmkWdbH/mawK2eJjsadqwBFvlp0Umd0hYjlCju8peUMnNJ/TY36+xqFERl/sjvqQCdMO2uItNx0
SMbjyE1maLBqG8AOGqvbgJLj9WDDIui/xce1GyPt5fBiGivIjiyuLaCK4eGFtTNIEKHaKjLCO6JY
1zhSU6FCj5rUT6Q+hKpOPLrFPiUglv/UKlmiu8CDXNMskJf3wUL3QEw8tn9dRJuO8pckUQ0mOHOz
C0XcKkFMD7P2V/mmGsrytUmdrO4epcXl851/CW74vEwLy2TRkMkqhD75kU4rC9yWCeliQbkjr+QP
XOko6nrDCv/EzuxsgwGN+7d3DKswK0wPVK+b0QNNXi252BKpdh0bKq0iD5pFll9kZbFCWrbj6h7h
KDx80aT294n3WuPaOsaXAXgeH3FUKBbcw2w7moqNU3rz8pWWlckknM0gN7wDmxOCl3pbgPnY1Fok
yRm/CNVDrDfedei8Emcfo3occu6GCn0piyqtT+Rixgg9fnQyoMWhL332cANZUWvGiyxTaMne0uBc
z+zc+MQSIGj6c9pV0GuOT2hQNf+dxeS5hIWCfxAbZ8WPE3ET0soOlre6mXSznU+XUUZi2zEAqGnA
XEjNVpmMu+gmbYx4Gdb73U6Kxb4aTu78ey4VSO1ni1N6VQDtE97M3lwyRVA3OLBaVuQBcdTqecTr
Cb97prvpmzH9XdaMAyIpPDJuKBo7n1sTMHm+05Q+3iU5iBX6NITvP9csJ2yTdqY3u2FMktzsF1N7
F/2FcyicPrrpLclLn3a+uuijEYHrutbBPbu4dP10UdjXhDi94eHgA7/a63Hq0fk1OklQB1n381s2
Mf73Yufy0XRU/hdKG1P8m1upIv+ZGKuSHtdOFcVcZuBIWASS/W5ofJIH2y/OrcA8aBBhK9dlENZA
PZzVjId1bMVfLh4S9bY4sul7ra88WE4w/vCRMO22q67p6ilCUhCYaGvun/D7pfYatkSw9RZqvpbK
cFNaq4yxO0794UgjuManzVwUNF6f4b/p48fU7hvxDKR0V14r0+lFDHDaOBOHocLOsnpjvw2WT1nK
gkDk8JN+gVPDH8VNHQgFw32FM2CVpaer6Y0t4k9zQdGx/XmCW38JQSSJraOjyl+mnHM3/7XSlmgx
3nZuSujqsH5ZApc8UXARtuaqh7dTcH6I0veB2PJIX8TLcc1rRMlpUghBp4vpwdtkX9WaLxKRg0pG
uElJ2IliLnqWHr7WsNy0XYkp7MW0ZjCjo6L5ESc0/3A9xjnitxZxtwouEhLVDo29IYay50mks5DM
G8n21Pv83ydOP5mvcVmsWEcmTxd7NakhtluK9AiWL0mwgJfHyYyJmcokLt7Vn6hPR5rPaHSNJA8X
aKU/gop149cMLzkAAjBZJUSM470RNYolT0j5I+KTtga5Jq9Qr5IpQNfv40yRk3yxdD0aurXOT55l
zRWAQcElLFJAAW60WKoAydbIeSo7RQfiNps8+RizZUsqn6hawJLueZhF2MVXWRy7MIL58t5Aymxh
Ct43XiexZDAKzOHB8AMLpOV1ZuD/adx3cQ0cTa+1HRSPpNEZrVs55hTxbyBiPhCMfUSK/eojsOor
I99N/Ppb/gq9EMLaSE5j3Sr9OKMF+2p52llHv5g/TkqXSuiDFK8COBC879GVhwST6OfxhJxzAoe6
FH/OUGrp5QC7kVUlcLfOTfEY24dVuC3TuJ1EcXSTEBVLkR18chUZiqwKZzYJjH48P34Q+CXwiyUp
1Y/hlcag4quaqNN8attHgQpPV8WD8PpBmHaZSWWSWIPoBt7P+Iyyr9q1cNs5Jq6gXvfBoTUlr8WS
fAAf2KfH7eRmBPMU6bwY9kQRl/Mq7WY0zEWsIZi4efu7BJeE45gOhvJP0WzvYNPKcQZ4XTDZqNmu
Sekk3daLWnxqbbZMv0IQLvAIiKp8NAznLAQcwklfzCO5kpC4ao7etm7koVqXtRosDgblsa5w5ZVJ
frzpEeX8y5vj4wReL6atPSkTOwnC29PHD6toajkpLPWYhkSLKLU/Wz6Zrvm7n8kCfp98EH7TI4EY
s4KCSwhrjuWtsxqHf+/ju9YOKzphMVA3BCD5fKBCW6eO0kz9ZNv+XLc7l6ti5slVcC2GDwN7qlpQ
bgnS1Rvub8XJcGxjdYSPc057KSBFuYGNHynv2tPlYKVTn8NWDQPePdsjE43S2RDnGZKyaEwXIbdl
YG74WUzbaIdolA9Hmz0oAX0Q6wRA83qLx362WOR2SIMyK17dpDrghaL24d+THfTBIFsMtVjSzf0Q
VUZZcg/oHVlLLdC2vIq6m/SsyRyABp1C6z+Z7B5gsrYZT+Ea5xDnw4hPqFN6GZDc78PUAEi7I2Hv
gARPoMfPub6zOifO8jGiV7ZVRNMfNwk6PTmajL+/gieKhUaGS5A2hWobabkcWX87wb6GLa7bBqFg
V4eKrlr9iAZKHCD4fiXuz98alB/tY6VmusOBr2U6cbvVyXUauA3OAs9NEOQWY+L+w5u1sNwcj0jN
q/ETSuyPLjKzAUYoTX9LHExPiKNJbDKHmFhNpzjhAdHubVkhW1qK5yoaG5/6/Rd8yPafpVdO0mq2
KvTOLxFjB0X3zdNxgfiTal9LkdfASzrnMAPr3Sk1/bh3TMeNSHUsK3FooeUX4gEbF1Gg0NM+P54R
aOGG69ayvPmArOBrSFPrEqO6XbPLpQMirfZgkyLyLKC+e8b/cso6eWoFF6hgf+WJkasspQ21Sry2
sMDQSRB7cd0HxUPljjVo1SlMcm3jrbteDjbRnsbq66me/W1/x+4KnevRLWmFrCBnhYY1NBDdNetD
1M2mYGDIVeTx9JFirnj1u5J8mKU0WZlAqTR4j5J50uqolbf4bIPhtZyR6kySeyFY3uWIoaD/3W7x
P/ZLL0LYNUMqEuqnp32s5w6ouuMraTWpEWBtZiuYy474pzFwgNTUOSnjSV4Fe769qX67MYa1WdoA
TZB5s8DjMb3HJ1Em7cI6Q0azRmwEyT5ydWLEaOYVAvavGzT+whF1/KKDQeVK4BT5ioyhbtJDdKdJ
yg7OvoTUcKqBrVm5sB/QOdvT/jReABqOk0My0BsbkbXRETbkPT2pMVAuYmdUlnxgXi0hY/FfkWqv
ItvtHR7sjZiOW+t/CuDKmGwl5DvsUDKbnccBDLZ5Ic2o7/E4IJJlacuiusg1RIlzE2VSytQkG41h
8gvDGDkIIkV79QqL4Y7khfez0YEfRhhmoFgW9NJYrQCl/fFbNpb/jJEDlH9AQfIbeYkncaElqx2K
9o0fR/Wzf8Ame2MNWlvinfU/h4zfNyLznstZYhce9J3dRM1Q2DP6ZBoYZpGGFlMZRKTYHl/RPmiM
1EtJH+rCipRWY6btog8vCcxCSEGOvFvZroBdLaRcT/5xvBXWBtKSdQxUtlEI6YRwZHyzp5bhyxZ0
0//rylBXfe12drbK0136UPjgp4iqtrpRUK8PWZ6l5fBhT1v8UxTyLlxf8zB2ZY6wX/fFm3cgCoN6
riguLMHkIa3sJUvqx0nI/OI0Ml2DIizNGPxEKYw+Gke7C64nyM0c9U77cngCGvRyrq4ebKdLgDoq
JTiLDpppOcT6ENHefW2Eht6UvbgsHlJFS+0WTsadj5MYcTVJzYHcHeo+NFSBOmdyLEHuwTTz19ks
bTRixmlA8xqadBU2rlPN3dr7BuR/AxLm3Rq9FZszHB80ANxJKNwVqcfBwPi5r1vXjlJTPCAbgPE9
R4dgRtificmuKmd0F+cdMRLg4ATqzMH764oQfnERQvwlAGcig/dVJ0QN2hEsrw8KjsJGFRqoFBsC
dB41HD+7nGWkYAQ+b1JH6fpj1mh2ZPVZHDRyzCtveBphZlVGlA48g1HUPW0Y/wDqmg73BlEFpnIN
A6qbjm7lG91INOhpgyKjLlDjKhYtyfOwWwYpCoTEjPfvb63zzsagc1m3uD4+RcEJ8dS6oLwwF7Id
K4mo53BwhEwivAGrvUZyQY1Gy+0VjsRd2k4vtmVgRm0dctt9u4H+Y8bBcFPRozoeDmYEKL0tPutC
1sCfOYhD2RAvjCHZlXV9x9H5edV0G3dI2g209hWu7ydEzIf+pT5ARWz6d9dtDuWtoSOPzBecY8T/
sVCEwY8EEPRP9v1NFVj6+xanEmYRKX1da8pAHYSYkFLRK60XpuT2s8aTiMgUpJNhRtPRUiBDr5N6
BqtF/k81gOWVty0THIhdgZN7ZMyHVbehy6iOLnI5RSFdyX4dau0uRRtHE2eBbdAWjuQmeoQQFqJn
mNr8fLjug7+CoDG1IRCB7duqSvj7gpUrs+J3bCpOe5ccp/Arto1eGODQHDdfq3xR/8UUfZaqWDJP
AKyn3qxNk3EKVwlN+FTvo81M0lLOEVVpMPZ1FE9JfJwHXLkbr8yiiFpuerMtJ/C9cJB9nq87JXjZ
hReeQ9c4TEc9wCkv/5wpnQryCUvckcWUD7WsMEu7OjMtprJ2KSZm6dfU/6SxasHdMOkao6t+CmM3
joW9pwVD9UEdW1v0sHCBMq51YPHPUS6zmmVqzftsp53bp5mNoBI5CmRt2Wt5rNLku7GFldJbVcWY
0xbVks2KESC3HIwYuesmYebATJ/1KtQYft/Z3TM2CwfPWHEaM2or9E0GOPWY4Q4Aq1wxFhwj9dtp
ApGS1nyCJftkmlNDlD2WJfU/d5px/1mJJtSBhT1rNLq3F5FBqByG6yXfduF8DEjGxulUoTBgqSPq
pDOCVmCG6SOQWVXwn9p8jk73iJ2K5Th4O5BdvL7szPSLgjGl4wanxoeGKvq8ZC36WWuZmeOU4a46
x+Pgs4VcsRmbcg2mQjx0rjR0eLhiMXoMGVAa+GX1ROhzoIPxk9sM0XQwvCw3yOxUUQQTOwHxD8Gv
Ji2d5XJ0+xhwJb65G1bArIRqrjVQSEljIoPlXNPH7ZCvNWzLporfl0pqnm8HLmkGFU6I9M5zBHK+
NGUpT6YQEJs9WmM5t1oUCbh+q14qPIVBZ8E2OjFM2qbzD31oj74wFTulTVg94d+W7f0F/U39NxnS
lFtunVDDLwvZRuxrlZ1k4OFuzTK9qkmE2WjhvkLz0oWn21KEfqaAEjbMEmQniYFhFpN7MDHqbEj3
J6/xFYbIj7wddrsYyIdBw9Y1ivQjTVAk7MylMoNQV5bedUVxeX6ruXL35Dnz9yrYxvqgr3J1yIzg
TDq2ZdOeIdapRom6EH8ptVme8jyBPQCdf+RnZSFaFOvjsNAiHM8n+U8WzpvAPaOTrM6V5ynd693K
g9AhgkBN/0drDSMHEo1Zf5SvQrbUsnvFpO6xwlEIQMN4Q/QfvbEWDvfEF6rvSd9BCZb3vJ2GDFL2
qLCzz7ty7+0BtNVzYIEmtiq/ogGe+IiFnLAkpoKtW+1FvIzn422aJCDV+Vrrgu0jyOTYo4+NU3zl
LvVyXEuKvuIkfovWIfSsQiaddYYx/z3KgXGd7P8nXp1IYhp4Q0qH9ybhHY3Lrz8CWFgDqXar2AYo
rKJBZUdM1OlLd4x09ClqcaaJ9tWsgXdh6Tvl3tJWNB89vNEZJO0kGI/c2XlXe+RsA58OlC1xu6eE
QAohqAcHoTBUfLb8jYPf0X5ti7IagfLK6vSX7B7IFJqqG8IXZvxApVgVyVgHd1a7A92xxjwijHUf
VM/Fia/cNDKZ/sAPp4PNYP3b8W/IDLV8cR6A/+qo1qtyQhh3QxS/m8oQE/OWDNWJjptkxwapypXE
p6HKK8cTvt4K5VPIS98NOgTQn7DCwpb2dSccxY1O1n1NG8dzPDiECO4pCZgeYw69y072hfFpACaY
4mgvQfHRUwBdg7cNMyFogLfK2uqaM4h9Lge632BzcK0fbMzLvoyvd2okMxbi9KSss+B1emnjWTr7
Wi0TQ7AXpUOjT5dN/FHrOkK7chawWGVxbaq+cud+CjjruyE2S5I+dKYfTPFTre12NB+kAZx1XJLS
0vZcsEiun+VnRZckjDepHPjvLmQKQW8Hcsg9+R63Ms9hHxFFo0kQDq60FJxdBLuDZkDf6eqJb6zy
Pqc85pqINym2bCYjETjjwpZ6IbWQNRWLYwQ3qoyJUi4lcq0UZO8Bnle5/tJuFUdklUbypWuQEN63
y2aTrsJa6UYRHj400eiUZ97KgFVL3vgmaryLTC0dWhYhddmFP3jNs+Qh/yCi2IXyILOH5pBoWoBr
c32OVf0gA78DPxxrlhvG3C5sfk9b3Ki0c3qKXiAalzzhmdZ0Ea6dEIlcFMibm8q5QPY/1wXL9i+g
ep2mK7r/PGZTWqVzbjx9D0NtntjlSCXMMcAAwNWK7V23C26/3Q2fUhB4QP6vFPnSEYphPNvVbCNl
BdjhWBxCOwgpWqGoghtrY97+wpOV3tMOg2yYOcwzHqYBERFd8DypzlETV+f+aY/TgFuvxJRGY1Mp
ebVCmNLCac4AbJbLl2Ufa8FfwSuzQ18zKxssgoTRtDE3f/NtvADMc9IXrsuOgEcbBLPeZqe3cUgY
9yGg6qqhtvUOnMMBNK3/Rjn4E9qXKffDejuTJ7FB8OUPC27ZIhxdYkG/xQOo6WHGDlZrRZETOQ1b
5yGJ5eXI3Hj0cwNwUyCd23k7wCMxtD1zaWHCIi1D0cb7MeTG/kiiGsMGkNFXsQHoxiWkpUH25mdK
G438PSmq9V71Pn2M15tAzAJQ1zbvDPmcS2iSb1dmjVzUawlZJRfze2Dkm7BN7CAC+jJkQO+bxIIb
4UR3mPtrqmVGEjhmSpMSh+r7y+Gc0uMN3NadSYBHhqfCmOHcO1uE3/iP3JIl+rRYMfoAize6lNQL
02hltxMmdzeta1d38nmCfFe7E6IofyMurQY7nuoWFmum0va1Pcc13/V80RBnvTkmlXi2MN3VNJ1X
4BXlKb7ggyUnIwjrLAzFCwk6hmqi2ZlVVIN9XR+C+mzQDrTMpC3go6pV5a47Vbu4GbVD6beNtJNn
lQUrCMhUUFNAQasSfJIUFoo5SV3KUrVoXVFo3U8gdzzuLpzkdaxoiWEF4V0h/EreGJWVciYFL4ub
HZLiVBTm2opzjOTs3bsMmmHwRcdiWLfBLtpD2zdztV5EXiqtAQIras6zJAv0X8YwN2RgtFOPKZAP
vayO01ehtGT84AehE2fwi2m0hoJpDAFAh65yXOb/8uSVA4g/Jnm6vkjzPRwZfGWe9Xam+vRKL2KD
18BqjXZUDqeBO7xNwHJPlIzbPT1c1SyZQA92ZOEveCvNArhio7CBJNR8mHK6SxGB3Lqf00TDjFU0
9RyVumJU5+XGU5wePiGZ2Yev8F0lq5WAyuDf+9Ar93UOHTW0UM2icy1VCh0lEzQJotNN3bCKsWGX
G3WRK6XVIyVnJ60Ne6Ln7049q1LLjF8D/6Bk0FEs9b6cqFfBr9AcRuv1nxtb0O2ZPTYk871wq6V/
mRqMfftakGYssXiRc+2U75Ffda2vtzDwQnj+mt6QTznuqcJ7c6tIEdZMxwIG12gZ69fH2KQz6nZE
1LOBbafsxA7ifvySQ6MEgOKIfTfBKkpDYGrgiNTurlTiZYIAszbUXc8uO3tPADkgvmCaTi59eqQO
UNRiNhaBTIDU+rYI2lDOoZdSsYU9aMOL2yT/UewbKfFGi+NGTqCyZxehDt8/osFvBWZMCBjNQA+f
rU6IPr4anl/kGbso0yFDq3GhXtyd41cWfFlsZtSe+jlV50AyWzBqWJLEYK/xM9rrMyVU3D9f4fiL
F6fNxRW6EDIBtOn8KdIMwAaTblLwcoh3uPvIJ24jOv/9guhjymPD3mx8W5sE6S5D/JlgTvodZqcC
4hR6i8CTSkS2BLRAC6aleL5AOTwoqGfgJjkeTenr8SvqRtVeebOTkay/exuH+v7LLWqtLPtG5aob
mAIYR1PjOy7a5Wv8ZSZoF+Lxejd47xfotKdh7S8tp91CRPFvzmvrClz3vsdDbF8ovwFfx/wRSI5d
uXGQYErUhK2WdX+iNYei3myfOb+Cvy+3VK9kcImkEJB+BKC731f+phMmKYfpwpuAHVcwJL4XqtQv
aHDyebO2fiPcj0qLALqho75T0xkpWhNM2cgKd1mWngSQz41jPERJQzsbrI4oFwrRSB3mTvNZuo1h
TzB967AMXSkfG3hUyMkmLIiIBn6i9KI8vStVi3YMIcxi9ZbIcQXGjPr/c47/ZLPzduMWMqz1VaeK
qUef4A8YQp5hbkYPVFcF4NGmNik2PhgM4zIzqabHNM6+mtViMV1gr1hY6RqeKBo3SVj/LnRhPvAg
ZCc7WbN9tq7ATbylpHO9NA6++FcUF9BZnneG/93ykwDL1tcH/b5dthR56o7vrej3zR2oSgnXtVF9
r0IrM3kaj2o9ny0N/oZKBKaENs0sWGccyP/tQRC7/7/OqV7Fx94kLGtvbfIuUhqacCf4a7ayLASc
aoB+eYHYbu7Hc3L5msDUzMWJCQtSvnxf7w/7lcYqM5r9zOyLzTTDlrAa+5RXkrVJ1rdnUCPLZq3y
iWiDAy7THvJOr0LNhXZMV2bVgNDS/or6XIwgzEvD37wk+Gq5SDG0pM+wqG/xXCkuHxJfjpDUAtOC
LvtrLqjzNqAq4XcY9lqp/m0xGnKbKuTFNJKPWNvmp/XuEIsQ4gWDE7LfHl0OxT6E5CuRMgtv9/OF
BUIdx1vweEb/0aRde79dZmXQu0CDnYVGEiH3eux1z+o7t6AyWeNmIPZAz4/PNJBXL7nbH5OH79iL
5pDjjxY1/1iOAbUSA2hOdon91iX9UDhqpBGpSdoZJZBqVa9LiVTux1i3fjF3to1sguBYXKK/xSeB
IhlvAhepWxFxNByxYTgWwMZ+RU5AChE3d2IQoz2tjlwJoixsnvrNsHp00G6cd8dVPkKGYATntEsG
gAnWNYy4o7PzJDrBYAEbyGImQArMfnx7V6otOPrSozq7xStP/03Ytxz0GUUjChfDPLq6IBUU7M3u
Fstd87BbIGDPFMsUiqkMipC4jS5U1Nn/g3y62gcXvTcavsbATUjE2n0XtENYZMjbjfGN9uCm/DSa
nG7Nbupxd+XajWTce7x6sHpXgIGKsGDSDp+eGHCzeOgAsIST+9wqSj1Szgtkkop0TYdO727zdzhI
+D+gWaDzCenJOV0M7EQIeciKeNO12RUEO7bAb3NDnJMI/LxbnL3fbQ+AdayIUcs+WyILWlo6XetK
ZUKbGuVu85UfnUc5C6+tmpncK4CzY0zApfGP6HfSLG5b4q1JBsKKKgv7oWDMUEcauQy8LfRlXMLF
zWh4muSrQB4uROyXg/1FcJyvCKL6sYfPwm5nESqndio8Y31sZkPqD4ubhteiBkuF5w9A/H4FrA6G
8OSInksYWkHZVUx6mIKEVxei5awspUYaR1+p4V7ecQHgToEW05yk5Ycv/yJzT2F/35SMWS5yTHf/
/FIBd1etVfwl6ha8sDmOKMp33gOzLiv1My8cgOV9CswcSY+RE0TAJvHVVtknWYe0QmLjlQzHGXWJ
G+030dzGLoCimOVFgEmReWu3o3hGKciCocXYEZdt89j4oTkSYqUs+/mmIgHJKw/hHIklkKP8FaLf
q2p2mIie0g5ysga44YExFsv6wgYEt6+yS89XYRslpityqB7HyUFTccsvEjMPQSxGB2WqStHuayKq
0EztsGDIZIVqExuY+EXdt+igTk11QmePDKexKNy16WXpIFxns5FLOt6UltIEbpsQ718vjYyq6I9+
muPsPPj31sqyWLYOMw0nRx8t8EwbYN7RSybQMkZpZtzKJ98e+goVD66nWYQE6oO4taJe0BAe09n5
w6C1s2Ny7RZ8KtCSS3hQVgsxIiZoX1OjYzbrwuvaKpYb85nr0B8+E9Z8Xbm4d/rTdNoevAlmbpji
lxCypIxPvpjYDElmO6fi+WV+37zH89t6YSAARvjwjazZB0wabDZnLRqd7NGzlw5o+tPQhmjoXX1e
G8BV2Pp6DCvm8Ift6cr4JP5i7egnaSJDxKHO9qaiixNImkJWQTSobPNPF1yg46SfbhR61OW6lVgC
kQicnaoKW9jhrdUDuGeEs5qwmPH41FP0sek8FUO/q8XM/P/7D+WoeYoYybt1M2jdCA8V6UIT3j53
H+N0HLWNOcN951yjDyDlDwFigesfLyoiVxyr5n7nKABfbzgrlL8WR6uNJRNU43CsRXBMqnt+xDeG
OkkAhMtJ+p2kIo69kWevVx56hgwi6/Q6HwxP9taI+TZUYVJVlPVVrHfMjNoU/bOHyvb07flFcN22
eJtgaL37ydJzGCBxG+P3F/YSp5YJobBwcaFYfkmJ2aIjE4M5dF7yZFqIqPQDE7Cc/5g2V5nN5ryN
W2Mn2CGJvJJra0aXhUj677xmmwLH1t2Y8z1kh9HKd6iI3LthYU6S/7sKUyCvbSnJXE3YJrAeX3OO
QxQIQDGYsntPrzUjDlt8iJorMkksLe4DqUNS4YLkihGiZHuyO2Cqq0GSkwLFvapUQSLXrRtOd7cN
ZcnmS0pazq+VsFftHsaxJRnMOaERwUhrysyLZlgjKft9jcwaiuF14Yvl76U+RbUXuQ7s4QsFFa+p
8MkE6W+KHh53EdWk3UFUyCy6Eo5/LHt19TA4x2oH8K7ksBelYQmSq4lNI1DQD5mMHbLyYdIRss5y
3qCoAjq4ONHBw1GXiy8HtG5lkpY4yuTTXifpeqnbtEgnh13sTSEAew6bfaJKKmWU+xZv3C0Ps1Hm
gebjc9owA2mH4jJEBUM4vmlKn8SRJdJGSiNSSiWNgdSz7vEhivZgtLX6Lo9793p8fW8s/ff6wSVF
h4F14xXWsdyNbjZ/3qw8ZlBk8sbXwy9U3GP3ok1vkdyR7yVHgIEkc6xjcwPri9qK/ZjeDUzMiEdh
DFBcPAiRy9I/G3ByS24X0uSiB7xX3jHLFzobOAkikD73NBhKI6NFovuPb06M0a2Z5Pb5+lIiEWvh
YZMm0aj9YDkq65buRwGu970z+hOdxGPxPnZ2cWL88FBImwbf/bS9E/HijAprvFeC3H5eifCuHH3C
YyN5EBHtoTi89PJJyLpASQZl9kXOtHIfz1rBc2M6Ea6cYqUMr7Z5qaprXrY+7vhRPNR7BLMFL31r
PkVF4tVzZdBXu4HFzCiNgtJrMXZPCmX2jGtYVBunks4L2815S7o1Js7K3gdCvgX6FfsivTlfCr3r
Lknf834y1hN8xUkGtxHGJjjYJkdSf0bGO3g/lyM0qNXus6c5h9LJKzQdXq77E7QnUejR7i1S0LQo
NSgWWuQAPahF8h4HTPhYcU4gtK6oyc3otpLdTabnOcW/sGqRQR+n4B5RyZ85NGTUbVSfUzdzRpND
1QGdcFMiJD3M8AXDGfSiQY477TMN+c0d77JPHlFEyXk3st13mQfas9gkONrQjvixN5ZKocKLDhxG
mqd/hC09K/7x2oi0qg7/WEoDbSdcojOe9JH8D+U5drpAIGfg2FmJLk/Yk/d7iYvDLmdzJIou6s1n
BB3pVAnTDmeXu2YpHwbTEkT7LloHm16i6x/DrX+SRdlyxU2ikCo3i0ypTULUy/9P7boJkutd9RG8
dlY4L2GjGB0CS79S2bFfVXLp06q4pnqtnTc4BeBxexWbfEExwUxLhR9MAK7tLhfE6JvG9NS+e/W1
f3QJACIEvEbMUReApB6bHvIhyrwCM6U7+3I0krMVh3g4jWE5yBvyHK7OYGGwvq7YuE6qomOga+g2
bi5gGW9hsQBfd4FW6w0R0ImKC3puxNraT6/VjDQtdSrFGYZuYwfixGPrSaoHa21Ssp7y0qPbzmIZ
7AJGiMe8WaVGNuX/aQIrGKAiJarEWUN50L39htaMXqjEdWTrS8+HAEg2nhwt3fCdMBbc3mYatac0
wVsVsM15N3Uq8i5vUToNtySHfImkxanw0u9d56gxKGkSIgTyVoH3S/6ZkSOzqXqPuZdgdaWKkpIB
TmEAjJKeO4BYZH37zYV11S5Z8aHxvJBHe4BbA3y6aPAQwf8CJPW4k9QsI5gulWYobWdjuW5ut9r9
8oci29No4AzWl+x3nFX6/beuMDDByI9peTchnkGlT5jfWG8wwXUGELsLq1d9iFzRExyYWiPX3L04
XQL5VLOPkfV4FaM+LNlEBTXtxAtGgLJDCZ1uKUpcaN06k9pU+bB4QNXqyLirPB85TRClJ+gpkWxz
TOZzjljU+RwgBhvk+Aofv2S3wXNEg7gDZl8+T3CZj08GvfNMKfukv0hdgv+ADRiCEU8SbgOYwrFC
yRHyLLe3vnsOeFAcAiJ5CYwwvWlY6NzWBpwpuIw3iYLr1GsqjFG2JJsvHHlZ1UhmfApeqatTk4FL
2bIet3PspsBhVyKDz71FPpbJqnVyfe/MOHzqRdqW3WB/YZ7CKKiQ24SnN/WWWravZVdVhBIBVCwb
ErSbDD7GStUiG+Gi1DgfEl7VtbdgvysI9zOsUJ3lwVcD2iDvn4vsiBikdo2YhXpqwNxDF1bHt7yK
MBHAjO/gWkzcTYD+FILCI5VSHX+2KcXTRYSctHCsCgigOz9tIfMJ5a6bx51+PQsbvrUWaUV3ZO8c
WxexPLcUewaHNpjybA4cfNXpF+GQGwCr1TSYoWUAH3dsrz+Ke0GaHc7R/4rkKRkomIATaN3pRlKX
C63Z48EHMLN6domIsaMlrTFb1FBpvpEOud2GqQ4G0netGBEA7uLHwIzqEC/SV1d4i3wCYkfVt+OV
O89cINxGhMLrXMmu4UutLscsfa7b0smKOIDDolTTYWOZTJDCCqbtaqgPBBAvAkLtwIN0wI/8xKx4
Bu8cCX3TMALVYNn05XaNyfUdMD6oJReV+CPNb8J/ppQYU286x3ttvpQN3lEU8bGlrcVP43XBnSiZ
Abim5rMEooJLx+RRyT2nScStd10u1Dfj6r2sgO6WTQh3Y7VZmK6jPQDaWE/S+M5D1yxRJrEY8MQu
+Nawqj/0JnpvUsiB1ngfG00ymITOr7O7qAdR+3kQrtdy5i/9aFAjHbaxRiJGJI/uEnKukGMktYSG
ZnaIrgGbV353o8yB3VjIE6Z5donXZ378wGK8+9EX/kGqtxO+Tga7BsSXkkTPYkO4C6POASUA16OW
DbjdyEOHwncwQDwvjiQ6ydVJEOOlQ9HI/DuT0D0JSJWvt2x9HmdDE7hZi9XDOZd2EkJSo55I5drL
Uli66TnvlGDKHwn2e9w5MYJNfBYDPru0giJdFU4rb2A+yNnqeK8jTMLMC1G7saFV6Vt6yWBR3SRS
a23GESYATucjFDpvlW3eATN0PE2ctEulZhBDo7Iav1De5KtXegxUSJyUQ69602qS6WdJPo/hu/+s
MrokMybjvoE07KttOjwXCN3IP6coMJFFjhlnz9P9DDSJFlsAyl4OrJxInBK+CcWpayVGCYVD4yOW
N/SZETi6rXoWNM7bIL76GC7jDJFuZMSKhaGA89QUXhMLzLWiWDbd7/yK42H2AcezJsTdrMN+HwXD
3wVKx2U5+K9IjYhRWYT0KwWIgvkh3xyUkj/VlrboTzkBLPnG3ePM2098iCFRnVqmgLqvsLB02NbW
7oZrSq4nWcR9+lkKXLmMuddPLRAFqv2Er/QtLC4dJzI7RSz7ishQUodrHsnCMVSwBiAdXxNYiayO
Z+YB+YLCRcZWgypWoZaWliDweDsloaiy+GINntE3uS5fig8uqFgiP/oiZpMJSqXfM8h68vxvCQbO
XpD1dm+bsordlBQ9emNT17IC4HXqSeTwJrcTaeBROCxGIazqnWnHzNcsg4Yj5KlnnmHqc6Il5ALU
W4a9DqDSRZeEQKNPS88R/6Sj0pLg7genbHyFZn7W8aY5CkVrxN2UOeL5FA2+47v1rsOkEsLHtdy7
CqRbY/CH6PMmEjUv8hMho8UQP+ReXOdHaMJNMTB2yNe7AQCxlreZur/rDAXnLTP5SraSCV7lyGIq
l0kI9SlxNLC5uroJMR/Lm9z+OkKA/+57DeAdoPcm5MTH47U9OlHKi23JD1hMCDAVVjfLhc4Rqj/k
1j74VsBg/diF7ExLWcWIFHpY99CyM7Brmndcn0CUVyTO2qx9ZpuVyqlYfWbGP861H2SvwFUfniZc
j6HVSyeWOPog+tTG/Ls6HsF3SqAbCguCcjnZTFXNUiVsi5yvjbaKGKXKTpQaudFzo/n2PTPPfKgy
e9oIHvTA+ziIjNP+FHDSkR4zecfVaV2zmWOQPXK7MO8v3GnrgqHT2DZNUGeciR/UOUryC1jwyd4p
3CTDQf60JBb2lWMwJuyABf6o+xtlt4D/kO2BdmBqM/ylGKs6ojUdl6t3cPg2M0xRD18hJ6nlGWTx
IT9/21qRn6dqhFK5FzHxCEK2rUS1QgOjnxs9aGkyCyh9seBhlWQ9L64jVN63JwwIRPFzMedymB+M
Ega9oGrAfvSu5wpSSetjKQW2HXbvsK7JUjyfx7FNy92NDPaGg+TuISv1904rb+8ez0RfsvxpWJqH
INio1z98SFYltqgjbCaQQzorClSYxnkQR+ALQFjnnjvzkCfIvFn6y50Bxk+dh5QAD8TWEBFv8zag
1+Q1YXcEtRzHy0B1qoHD+BysBWp+b/DfpjB+64fpJZYMcG0PWo5HREH844B16sSxA9eedWaKeJkP
nbfrLj2D7QHwP1DsClWG14xQQa7lvyUP+h+/GI0+gzQpeEuSIgx8VFCrg1euhWz/gPZRL2Prk/Rb
4Ru5jaSMDubEG2CMEg2y8umn1XFh6c2+JY3/jAJBnGHPJOohC9c6/Pmf1zG3OiN/C4/qF7IT6TvS
etylD9CNFH6Y9MFttrBxWE3UWOmIyDtEhGgQsQ6fwYzd9fnIcrk6ccw1hr/1rUx8wfDX+g0ipfbV
GGQepAHCmOXgrXhxxl4gbohWIdFrJVzvMnvALxvB1ScT1RWa4xrHYJ1jx/AbDM/kBZuSqnP3JrUA
wd7djufc2dZxRTCepIwvsz1pKOgrYPASoiRtYY5u5HetkfQs5qBxZgQCi8PMZGPKXXB9FooXNxfz
XEnoZe5EGNuVM5H35ofVwnRRGjociq8JEDWUEWn/XIvqorWBA0UqVwW9LUZwYVaU9VZPEfzKm0bE
309GG8emUj2gy/FYTpL6+qTB7IH6DeyI5x7TKyLjRMPDk9X27buY6QuS0zaHJsRr9T1vBAWn/JTE
emjPZTrEL7bl2c6AwfvJhJHQ1E8XHGRJZWWFv+9FRCEYpnrHIWtIFZqRntBBPGD9ga9FkGRn/pIk
DZh6bP+TiQAwM7ObPQJytIrKge2I3UPSLzRJrXOfJJfCoFDx/SqJmyjrisrV8nG6R4bbrQiD7rMN
XQ1vjpdmlN4dDTjpU7RID3eLg841phDAO0ekwmpwBr+88GmTBZIqM9AiDjrQVQEjedryqJuOD1Uf
vxVMybxP3weeA0Lj5TEhTNtqMCS2+ACuVafnsEBxBebdBF4i/bI21+gPM1EKA0NWgEHGHJJAkjxq
GCDOd8+zIRGOpjzcIYrn9PfQCQLa5JCaD+1CltOQmuEIgIq3q2vpmN5FGn+Y2O1futb0zcxWf6nh
ISONy1Sm32nem5WRUblAU5MS+4mWr9ROVRWF4SYI2N6KSlZESxjiDQ/qcO1YR2Tsq1ucmfTwdYDa
qQuPkVXSvk9c4bpMn1kaKVP0DH9qWuAmd4Mrs+6rRxzuKLnyA3zEOgUu5vlABLF71x22QsOXeOVp
U7mwFNg/Xya+fR9GH+7uBHs6D7ve/I8n0kskimzpRiQFdD0lXOvGA4ODcPXve6FiguvisQp7U3M+
ZfFp2RmrOEy/U/6dp0OOTYtW8qldb1+VBiU28/nf6yGn0e62KdyEhFqJDESqJ9t+Xq5ToCqD8wSS
fcN0Ugah3/Dq3UiMI6cwnZDEco32yCTJxFeEtUtqxvde4rMP9imjydkq8UBv69yUGXakgjgFqpXh
5a2BqB16UxGButzP5Geonq5xXrnuXVwR1qJ+Bc8/wUeVMoOfg1jxVdb1UBNMaz8q3dKjOZ+U7eDc
nwL+hxYOMbPAO4yxI41Ckm5677hGWBZd2+4vNY0sN/rBl9AkmvDW0SwNUARhKnWFUzl82eRTc2Pm
8ASXZwobwuWKmvIyXUEo/RfUrBW9RK0AthUFm1f+r/o/lN9j67IhRaguTpqfmQgWFhK8dQBVwtXA
F6vbTPltHX6omIHTcHgPMXU6SH8dRIhD3N63fCplgSMMofChQP0ixsLeLngs+ldDh4SsBoypXy+P
iP2WADOyVzwcAfdLVq0+/tOcxwOGGxq2Xu7PGIylJmjFVxa6zikgya7/7zZcmhF9B+0zJyABptuR
dBD4+3clZUGW7ai+KbSwsH4Od00x3UsKp/y9f/vRcQaRgzTtRNTDb70d5Wq0Vws4OaCnTzzawRZE
Qs1InWHNCJNfhNasYBbfXwuV8f3wPMCzLmknF7go4HtVy6DkqWyO9nxZFfBb537xt1rX42pZ5hg8
vsVQ+j774SVjz9ZDpIhtuXkPFqK9nmKctXqyjtzpIrC+gjLMgQgL6o+ZHHTKVvffZ3bk094pHcMO
WBhMGcJcTBWKM/Rn2UiJCJi/XoR5l9a0p0VCMCOMTVuK7gqha+jZYHTBzlKS3lgBmvob47gJ72L4
xEEerajFfcqCdpm97UFkrKZy9508WfwmEpC+la3pomiqOTYMUWGnQJW0XQkdbyLsQ0QypNIJTUyW
jHs+jiShStYo7ms4vJKGt4MPYHN/UkNCJsTahgVi5FtntVmHJ7U9z/6bGHnvlWMg7xjNDdziqoxg
pY4xX9ZXH7sUDMDUrOIzWIwdkSZGlVsRevT5Iw3lrhE6fQW4+Nfku8NN7KBdegSA0HLETNTOu8GM
pdt272PZBavRgXCAdIwA7j+Q6WP8JFVfo1EuoTlkTpUCL2cPhUYK09zW7sq6sMeRIKLf/oYfnspD
AybHTvzqfuVu0V52ClTHx6mRc1E8o5WDOEFdXa1jlh7IVBrTd4X5ymM2GdYLw27vxtKFpvj5MYfW
SREOagRlJ3XWl6xJDxLXLs6+Lf8y9OrzUjYxcjZL7PH2a/kJYfubNp4as+shYVH+EhlygZ5IVuHF
90v+yaeFMfuZTuJlzcYq7Wezlb33OdkE/gb78pAD/7by1lf3ylcS9F1XESE+u7rAYbddXgKanD0M
6GxOpsBRM/xBnV+tHCP/u17LTLaXgnugbGxHJiffkcrH5yO3NSL8bFk+GbkkANh3lBWOAwJh5/hC
YbHjCV0EDd7Cq7twk9Ez45bh8N8Y5V7X/us1o3xQ+Z3nrk83PwE4eb+XAr8fscgJuq9AzT+x+69r
7Fzsfa0YipFGkwV1HNoAskbccgevK5ftZCj5MgR7CdILR5H1VkYGUZ68dkEBQE8wfrUwz8Nw8Rce
LIYOZutIHDvxKfry1aQQ5MRzqWtgP+08oIVjsVfSxKBOcp/Skdh7CZhaPOY2QT3LPOnGAjQ5CkrL
t36zCntJk88h5AVXdCw7OTWu56VkoC6aZc60xw1o7Mu+UAt2canp5sdcAqHM5ymL+RXTxVsExZzU
cxMLorwqDC/CuwZNOoVFoaZ+XICegpW+TbRSnWxDl5VUCUgW5mi0vpnKtgASfRCMA2w65f0R6CKw
k0XfeCsCjNjnjhKLJEwGXid18EbpxN6h5mTP//1YXqSDjPBlyeNfL7RWk6p1XVY8WtbRvSfc7+G8
PpZ8urGLHj5z4HwLCzDtJ0RnZEFlqj6gWLWYou2BjOWLMDwH5n/VIu7sJKzEc8vvus10pqiP23vU
C9mAkv1hvxHOZe9VcjHF230Y7hkSN2nQicPfHA+8R1HNCMgv0xS7V1RcEjcIgA+JERbO6dlaYniS
KzDRc1Vk5WznJiRpV8o37fq4XP86Z/4Mhk/hWTgSA2mRjMmFAd84srzz2sXUAzeBNA5eyHQtG7Sy
e08DO5+amWWzRISdi5882cw6yqM2bpQr+rDKnauGUE4Wm/nSFIFytxcZSPOzU4ehioHf4Th3qzJb
2Ae7JvKVftRwCsDUKO9R+cCYLaFO3egRS1xtcn7sc8WbggI7Jbx+wmHC0GMWBneUgk+4VQ6jr5YN
ZHwaTYoOj9k/Szx9/nJ0qB5dRyCd+cKMx2LK40KPz847Qu/ev4HqTF26zbcJWeKcoGJgInsWL0LH
6Q3vtGYhwbdIzpGZqW32SrMwznvm4L7Wvkmapyht+jk1Q35GGT4wu5MpPj7ke+tCasb/35T6W5o6
nOK6tPA8v40wpcDoPCxpoZVPq4O2O0uPYTW1HOjPVGarUe404vxsgz3KOe7sm7+0PPeaPpHPDYrY
f/hUUKSnrk/o0t7C8Y5mL7iaq7HLcymXOwKHv4pYfSDQvJLTzL+DAAsJ2m08ZlIXIyRLvdZz8eEH
BFRBCCB+XQ5/wCIPWvnhTXT6wb2cSwgTUHu6zbrf5pNt4N37W/lIQi9ulqYd67WTxrIzDGvR+JSM
AHrmc6bi6DbmnIL+9ChsfC23Ri+eHD2CRU9CbALnfBuyFo0x5yAoF0VpKQ699TZIEbpIA+MJsyTG
DTNiC400j+g0GvCdbbugVbd/jXkoc/CIoTYLTxaewmv/dxRQgMcDOAVgnl1ti+iAPmtFYGw9a9Sf
2l0y6CbbWsBeFLN6OOH43kUE0rylSVy4cBM8jR1GnyFaznQX+uIUrDM01TtMQu5CDir3j4vHimAl
8tbjGOjWrP8Xd1/4/sb/RJ9Nv/Fa6rC+CTJS7Rx82ZzDigxB+xi4Km7hOyxJjO/V8pU/iaHFGL67
l58kz6EgqystdhIKWU6WSsNCs/6WSansw7wnU81MURr9v/ON17aQ3q5CNVVW9SDy3QmcSTWgYXQW
5DZjX9vLCZnBX5MXZ1aFUW/i9cYuhyDe2IawJulVpP+liK7RH5zJCQxjQmQ0RvI+7yAqoyZ2bFCY
HWd82A1+FZOOTEpIWf95leTH9kHr57x54gyp0glWH8yzKEEtW7a3Q41632fmWHKRPoqyZc+wiJZW
Y7aAbaeUyilgMPlr+NHurG/5x986je0PLUlNwY0iR98AF8uFfewb/0IBytF9l2tTJ+YOO6+CsWJd
BotRd9MbiNNa6pYNp4B8s4IEwo4Jye+IEasRYIgW71rVUQQlr6wIs5j0jePiTmQs6XIl024fpiCq
W7xhE2dp8JvQ++/1lNh+m3rwBQGcFRF2xe17j3K4Bu/O9eJF5ndmsTEitq0iT5RF8GzFOzCR8G3Z
/STPP+dOvs3sjN9NMpETyksietXw8UTMPLEBKK6Oc04f81h+YuP3UaM1isPRY6qHQJkingQF5eAN
ox8k68E+AXpofMrHyVKl7zWfXjdasWRqTcluCka/F3aZ4JbgkdrHZxFwwV7mReNLxri3L+LZ9Fyq
Y6vOtSufF/iFjFucIxzNsan/H4oDD+DPM8HPypDgCnOUMDYo/8njprnapq5VfEhyy/dOGDyJKXFB
5Pdsw09FXudBinzwTvpQawzT3suX/4Kq5gUygPApVLZgnQNJh2bHTSkT+PkbnQ/p+VgH1uItzBI2
dvE7BMm6s5pVZUg5R8yNQ9QSItL7Qgc9Ayk32mFap0nCBH/1gibnYx4YPmOSW4PvNbKY3iqZPWNe
6raI+O8yxJKLgC+oBkqu5uOoT2zFnYzV2DVuJ0nuvNwdLC6rlSpwZWMDT5yg98rTzA9MqOETjZ21
lATnD19cGniVTPoc2dnUE/+/0+jGF1UBYiiK/GAolomjMkEtn2TJjV0O1NfuexJKJ/HZB5GReAk7
BgSAOrg2y5pGzKmTkZoyfWY8n2I/vuvT1TrocEbmWKkERRm3zGwnqhUzt47BLZviRJUR9zP0oxZL
f7nw3v1gXHUjE5QNg8v9Iz9t3p36dmHxBxrX/sdcOGkFNz5PPou8E4IJHzbo0m2VcSORCaeWeX+o
Umc73v5/kc6Qfm3saZt4gtj+KPF81WSMdakr+fAw+MzUQcGHJpYEbUIYHfyI0eYJtfXCkxuMlh+K
H+jM2wClHHms5EF9fovRt07Jm+U8qgsEgiNFsQRiufTcTAfbvOXNxqiXWNz+wRuS6lciRO2YorsZ
zQzVj5v7j3fWI0EUB+Rp4Zkl6/9cjxK1daLGmwRn+QTzmzbyqdLGvAZA90Bu5VMMTo5QJLS5cEA3
3unt55UdUDaZoRU8c8u1md0LfYV1ZpdEHTTCXjnIRJaLvuu0DkyswaYc1FB89N3gnl74lCaJhgAR
XlEr3ehN91zzDiKA4RFhM4U7VXr8I9/YW4TZsiMN6I1zkhlH022f69z/nONjE2+r8PcpaO/CagoV
lveW83HRW4O2a3Mcsvr6//xpO4YuE22fkcDCONxlxLP+rCYAlUBLg5pL+2aOUN42bgB1C/SFuVCw
Uon/2GtaQE2PeFZ6SbgQ89OHBtSFs08k1Ah6zT8bcZqSe5DDsrs/4baJMjeZzlESCeOpLGQfNBTG
Nt1/liNASL4lMFw2914cy1sJ5jOMDS3pZvZcoIGk6poi87iB6sXX8AhrucO6MHKvZ+kXgMx0Khzu
6Lk/enr0a0N9Ar7Gaafrup4j9b9xH+KPqSbeUg8bTsNYK6z+Adx5ppBT4tG4j8rQYmDNNldAXRq0
l/7otUuwrK34bLRrubzQKWksNepBW4Y2AUsWbc1Y+QQiZXvaeTJi6OO9NZmzrmyFEZa3au7CzPUo
0uQenNbWL4dJeSGUzdaW2etx0Ipn0VriCal+BZIl1EcoWEIR74quBdji4RzMuKATqSJLsWAX1v1r
AFSDuqwcLZR9R8Z3iKLu5OeZvwWHxBtldU+1EQpV+aoqG8Tj1Co0G9m59M+ODA3oD1zxJU89wRlB
8T5ZhPgiSCjNdXdijeEw6Iq/ZP3Q3oUKWF2KhyUTFm4I0ZFjwXyOe9jXDjhjUemyGLFzHtf0D773
DRICVutY/jyJtYvXoUySs/HyoNULkShUgceSLPDkPPHxE9dLhPZBmVUbueELMeu/EQVTb6T1adqM
KLDQf/erWOPmmxt4z7upmjlBDJXZgQ5VzljF5mBveUwMTi/MtmvmbRN9OUE1+Ah0YpfrXBY4jtdP
kouVWaAhOAbS946Rt8G7xZGV1HcZ3MKRFJX/iu6YrnW69XZiDuI5L3zzEI3KcLDDHNJoesE84DhC
AI3CCFuxGb8Xknm4aAZ6Ah6i6ZdZDN+7XAfAwDE3IXMqtfn3ngBUCJMJp5nIJMpdTq8MtleFmcQo
0gsT2eVbZTUj5NE7qgp0hc+HT62FR98aTws1IAIRVMzKB9x0PZhzcH31zut7njw+OgK1Q8ZqookC
TFaTTMZf8fdUF/soel5hpv2GrCiEVvmQkmPGuKXzYLQZDkJSDTQ4JKHWJrqsm9v9aT0ErCB8YpHa
J+2X+H+JZIAzf7Dqt+XKAhYfvmPe+87fL3VfQg2rZQLFusIjKsTw20QsxeKiG4BkXpXZ+TJ+CKD+
sgXL1rZQ9qAoBUjHXWNNN3bnCWqtSTIk1SBjNW0e7wUDkX2tguxt+b6qDhvt2FucwwvyIh//1w97
bY0I1q2XDz4+DrVOBUDJdfy3XzirRN8ECtU9+IhrDJf+CoQ7vmcOIebnw6pd2UZqS9CRjfqtjqRA
Jgd7WH3hldDpG+txwWadZ9ea/Psax/g/+5w8/n6QyRTrdssrkg4Wdd6731I3yKjP2RxxYZeQHvqo
WOi0+RhE5Dzx6iPeG4BPT/cPFbeITvReKZy8lcME+HlLOJyvDKdRsH0k4P538xSoAgOkNVnvZyF9
Ej5Juf7shXPvkLn4BCoP/+Wl7ZHJU58JYUxVEonp184hKBak2k5iiENhRfS+2Fi1eZBRWW/o+Ik8
uDFZpdmRcGe26kK57cOowh2ET2N6XgXMy2rUK0y2fczZTpcdvNVEnav0YYEO2EOHUWff/hmyS0hD
mt1naB+lUhDXQa966QLl69GUvEFigkHsV9RcGQfUrAg0fBWfZjnP88eu9OyaW/0SkNgfamPY+qWC
wUDCegpvZWvstU/1kPF4pC7HJ+dM3nQqMURhQ/rgW5GMmxR91diG6KbPSOc1oXbyQ6YQHrKRjTrs
I1Mw772UGR2shki57ufEX6GEJXBgThiqtA/HrbC/oPqlWcz2i6lqMX0Cta4DrP4CsBZBiBgoi4J8
AxIPmHxLqDynYCZPJZnKj4Yp+9+zqebTrYWd75wRH7bgOwT+6LvfAuaA/2GwlChokJF6p7Oh5xBx
ayeDRXP8feN1rt6EmLLBuSB2vL1V3ix5oJZJ4oDQShx66XkV9HBaYW7lr/QklT59oUlaMrq3mhV3
iqUnXCCieeEBy29HAZkBZGvV4RIVWPNRDMYxbMNtGc8ByyBRMgMcxGQQcfzGnZkddkLeakyRiDLv
HqNGHGerIDLlM5d0Pi+CJP3nO9uz65+39G+Puk57n0M6pbO/v21UEh5jNOv76QhsLHOtje1XrAPf
NWJlXnxRMjZjFkvN5syD7ncTdYWnO+Juv6UxLZ3lwvD9HGtzESy2R0GqoDZqbvQFf7QLyuD3G48M
AJaTYoOr/1owlzsm5UdEhmBFn5EjEVP7c4j7/pPfLvDS58yZIugFF7eFFMaqs0mQcwAPsBUHWrsJ
lgLHGxk/MUWLq65xhMscD+WGvPKju4gQngtp04LixJQj6UsdfBFRElTNm47FtdjL0bK1Kyj1dh8D
fY5hVAywXctBh5n02ioJ1ofyg4RcakuKoTdCVqiObbRluk1rN/6SzPN5M76nf8KBYRTZK06YA8jX
OCuA9I6sw05WYyoWIWuTLnGG6vkltzzjCtVDXEZZD4R0xp3OesMkchyKLf152kd3R8t2QJtVv/Pm
qQDbIkU/PezWyLnp+dInpz6XBPfFTQbyAZvlAnxhIB/olP4qfhYqhy0as7Y+tO4oIY+0xa9qrPXR
53duLC4k7fODIYhLLl/+kFv7BZhon8OMCVpkYLP2fdrzdpjjY47mIaW1sgYqcv/lSst86jVbFPGu
Nt0u3j7tfHCjkSsqgEmE2YBplYYZbzM9ImT5zrTORbCpU4LD5C01guIJmejpat7h98XAQ228a3RY
pSr2lcjDwESD3POYw0ooCMXQLdUFHxrb59z6/NW163DPv4kuWjRXifu5K3+oeEGVjiOvG9O4d50k
78NWNvqoCvMnKJJcTvy4TUGD1AqSKnPOSKJu2WHSraN1cnzmhJfmFg5XM6Iz6kcLdidEUBmy9Q3e
FzCf/mz2WB+iIIZ2zYpl4o4IXCV4gLsBOlfj57EMojzJX+twvCBm6CZaYJMJudiACoVjbpPHwCqE
BQDk688WNZM9LDaqTkWgCk5XZ85S9IluMqkN8vylpj4lZEhQvVT1usAvlfb1uqX0nPeqRV7GOQAo
QQuTlwmUg0Rax5/jEjataBJh/CX3OTVk6PNQDpVVLrimURf72cOKLWrdFky3yv2NdTn7Lt4km/zu
WZGK1A/aIwLlpe3VY/WaHzIPGFPoY+KPge/5ytv/7SDW7KccY1oT40VWSw9VjR5D4QxKC9/RjbVB
gg5j+WnshI8RQ7H/XoWoS2Xsqy9vl2KrD3A7PMqwwYpPecYX8xMY/bql+LsEAWkJbBfBZ3t45UFo
t/p5XBJ0I/gM0VhIPjVfvzEVGyy+erLKJdVIef4YMl+edxeO3vKC9GrdC91hNhA/skJMWpU770SJ
bIvjPYuksZDlOUJLA0e9tyx+i+v3XH3q+k02Sdc2N/hp8oLItimjRR6nmPm9WfKMxponUF9w9juM
FY1mIlrGuptuePSLH1eGL9SglYCum2LBMgltq5Ew1dHDhEK1QIe9WuTr+d+orEIWKR3nPJ8Wy5In
Y0aKs08pT8B0xZR51q+VxwylGgI7gp2wksdWBfk7/pq/ujcZTv1p/Ct1HGWetbn77EX4ITUDwjSh
2kB9YYq8TJrSDTiqghOZzcduQZLig+ryubHJm5WZ6OEqLnReQhT2iUr1VS0pukTegrWIEXoBK1kN
d+jcGweSNMombU5HTV69wXV652gXhmU66yahN3PP+J8m/ffCQd0sywYYo4yg2DYEtgKi/B02fDH9
JQ2uTqCwzaNvXGJH4iOxBhGg+TevULzbON4BMu6mEoK0kpbVNzGp/oNlCg3Qiqdgsb6tybm7TJpO
5g87SiYULeMdjcstzRYpRqAYHMHGWKACdjQGeqZGhCcyGP6rxTo7P+PKalZacqRw6ymOUmGZiZ5b
0hw99Eu6Hiw8OgQLUVIzbVwZy7TVUtyve/LrpAOJkoV+xSiYgmlSEw/mW8n7dRb/ieT/pDVfyPXk
vJjzZpHgvYaqx/N9sCBa2UJPW7Pxpmrm4slr5k9WmrbTQM3kMHWjg07jLgMWEh74ot5SzLPR9vom
TzVLNnqfW7xy0C55DvupF9pLtOM5m3+BUBptxGpXBd7i82vZFdqtqrskUSR+b/yXu5OKhWymRAnq
98IaSoT9z630fuQWrwa7yO56e20Ut5VhguAogdJ12SJkovvrRuRqtfoTmDFIgkIKIB3tlSnvsGZc
yyJSlFsrJSkuZYyZWLvmVs2AZs7kO+rnr5qpSAuOXYAnqu3h827YnfVpjp0uj8HWV+/fg8rOKlJ9
PbVgsT3Mi0tdzGnXJnGPsXOMA+rrOvm1GZ0td7AxiIrb1zzjk6C6TvVQxTgSx77khbgWMsnRs3E5
2oZpW8m8Qmt+dvuS/I1MsG8xw1KIaTbvMqTidVOCi5wqTzHaPpCj3XfX1ngLR5dkmhCjr8A0kBiU
VnC0/ZX7tcJZXJpuB7j3RafydS3oCqR5VEz73Sc9Rtrlr+nPaJ884VLLojy/KbQN4lwtkl1yRwS8
vWIhGCCBG1b7BqXIn8+L8LC4g8Uo/w67WbdP5Sz0UZZgJTe5c1WJrJ6ZLR770SjoR+yPo806xOsQ
p7iN5dtfhOXEYJ6T7H/tUw3OqUSNfn+8UkYlu0hlkfL3D+ObNUWnuLDm7w4ZpCutE4O48PJYHnSo
C8XPnP2j1aG5C0jjd54wwfaI8o0Yfxnoxd+yoaWkyf8uxsc2bHWHgEfGjKLMaki/NTF32mkMV/aH
xvn3QZ/bCr+K9HGdvRxkCR0tnQcqsBx7l+07eMX7w7Q3AL5H7XTAgeKkflrsvMvdriPgUmDjv7fC
tvhqINHoM27VKlu/rbgqb3gnTK4IBoy59LZBpCzvhbL+a6Ibr2I7jhZFYsjwjK1sBQmhUkvul/2u
eDDbvArRu9CJUyAk3Zv1/8x7AywqBDve66GdWxbZQMpE/Ps3/ShY+yZqrW+rRmt1KUDs06kANttW
612SEFfbzVInZcyqXmYOGXwWm2fttBqQxdTGiIOJpMKNPn3SHyDCSyzrTMp08totwDJjIDWGeHw+
lQ9XrRwCDMJwzrexSiKizoZiycLTiYDkmZbubxd88YvlooyGcH1IqB8RwQbnnWbRu/frceJpM1Lt
ErxPoCjvz4xnaT0R9UeqPDHI1t2cwWjPDvJEkaELI4Cg8IxYOHZUKBg5VgHd2IVK6BoDhvZCKf8e
p7sgrVLzdSRfHR8klnA8bURxqjn6l2J9OPwz4xmMDEgc8OLmy52nnIfKj+BUUdGlZrD/sfOPb2gt
apahd0gPy+r3hwiD+YrJ7V1DURruMNRmBarEu1C2HQpNbbo67XMwapmMTUiGbuXS1oRusMLsQJSS
fSWq/87TbvRh/YQunYNkr9Vwo07U9arxBG37lheaFuqTjAoRx4E0X1RNe9JItaX0B2IL/EI+p5dL
x9q1ZDKnz2Pghfe32R62YexRFQ+z+wV3kAT+y0CMXv+FZ2Zwjql1pSnrw0VK3N+58fdkGUmK0EnH
9VEb6FSiRhw+CJyTuJNK7Z4Oikq3S5NyeKaiVsBWBrvLUAfFJ0zhQa8vzQ/9B0mbyJUcL/N4vlc2
YTDiLz1Ir0EMZx9ei63uilKwTIQXa5+f25QzXk4iHrEr9jYr4W8Bl/5PcPsgjW38EwAUWbHUxCxy
S2ZksGZXL3yYS53CLUU9i6OHnSm2nY8yfJt825e/08I/OvLpciL5SGU+PGcSOmgSdN5O1An/Qg3y
w6TJO7i7ng028VCNilUpvvHM8IPVKJMyLrIFmYG94QGBCqpFxe1LSXrNp7+Ijg+TZpNfqDamw244
8b02oaQ+o0Smp+kEEeaB8aISFSkBJMAoLMHgeREjtIptZY5kJKs1fVZ4qnJi+nAEKrVB7Gz3g8dB
mh7+f+6eMK5msPtH5tIQTkhChnIdM7e6Upjl0i3nMfQgzKas/QPFBm8WoE4+woPVaHOC7+vg3lgL
L+4yB0daAoyIesCGAZ3mSsMDZnAnbxcg0Llko+3EfiwN47OYJhqy+92Dh2L+qtaQHcSllvCXZGOz
/Lo0NI4GJXyd2hWLlMJuVL0gVS8MrOsRlAakpxBptiT7fDG5KuM3MwtpsMdCUwRc37xmLTIYDY0W
HH2Ore2ZRJZF9Q6/Glrq1VUGaPOPwO6thTJHdpaYOLgx0Umoj79ZMZsRGx6Ad2D72LYM5a/LG295
FniOA8g95wsOSjzHfKrl1j9EcyRMU/oG1ppkKZlAUo4aR2PmdXWbgdIh8HeVYvg77NN8l/Jw+Ms+
gF4uFvNqWoADa6RDQ/W0t8eO/1EyPzNigz9UhWWUT8HMR0Lh+FCQOzUmNb/KDrcBcqB3GkFsI4qH
Hzko1loYW44yBdRXK6Zs2E7Hnr7SI6b62HkKhecipSRM84qV6BWOUoEKIKfIa6AYWkEj+7399twZ
5BmzYEQQU7mlhtbW/hJiGIkdNF3XLW3hWgFYIHr7cHeHZl3lw0tVx4h2DDqYMC51GkS82yKSFxHt
k4K0BdFAEjZpBsELoXH4EzvZf7l4ckuCkE1VGZWvjzWhpb2pLY/2GZQ66+CpTP9YtT29FPMyVEvV
TZL5BBVyL8tLPKcfnhl6xOMmPonY5TVti9OyBjU43LpjJBG7S7DLU7fYOpDbX/yRU3IlJ3w6NXQP
QLxrDpSCCB59RqplDdOSdKvu0FQg9+ux9DkChYmRF2PeJwkpI4jnqAWMACvXdH0HucslToUrcMzo
YMc0UbLfCFvSJPq12S1AcCbP9g+n5cqlT33/WYkDk/h58QYy4vtLPXXjDfq5pItifieqgtP8SZh5
F9oXO10/bqnVpcu1cq5FnQ/DwiWyEH/EAHft/QTNIZRiuyHi/p3xz8uTFvnprvJqrToeA6iIm6o4
WaIaplufuLC7yhW9mVOdZ1nhJluFbQ2kOKhvyeHn3xQ2DzdoxSmkAvYTYA3FO3yKrQyPcS2qTOdr
lUcY2uTgPkk0QorXHA8jw1dQ4jN+0EjoatQH6SaLdFqGnTzKSx2lHkwZ+c2rAQ+guaAYAtaEQkkU
LWMn017Ojs8rbVZNMUTFH2T9xdKtvwWptO1Sq8kpcdNy8IvGCXUOIapm3nxSwF1YJQrtPJqo+m3Y
vQPv31kmrfJB+oELoQWRzBmLGXZbUKyJDe7vkBXGQgB2qwOf3YeK11/clrdiQiaMC6K3j8/0YoS4
RmoOhjfBj4bmVPBrjZXJaa8S5CBC1pH5WXVdiIe5uqAIj4dovsJZDI83StLWK+voZmNjFc9yL58J
fiMvGPzigi+GwaqTuYwboJTpnSb2+TUrPUqehjtKZM+GjHQaJqNNxvaTvB+4ZGsRw8na/eD7EzHk
okruxBNY1kxe9xpMpZAnzbYpYD+TU9isyUCadGc+YIVZJRhzrQRbvLi4nrGNKkq3ApsO7oKYs8Jl
pdUi4YiP00NMDwJrPBbqsGkaotwad6yJjMIRJUB2Q0kbdYw/27yU4K0RlTfvFVnvzTc/sF6tOdBZ
H6gyp7W8MpkkX+LPDEUKuR8TEP/xk7tzrGfvPvgXSaEhrVZsZQnDPDKe5TvTrhyPrJYaHRiBm5Zg
EpbH/rZdhgyPGtBrqWXPO43OyCI6WOqog2kIjX8ksI845YwR8QYWVHM6E2Ry8iNXkTw6onMOmrKg
+DDPupGj5ZCzJJbcYBryrEQWcJAjlWZg4MMYKTHoeAlMbps4xrExtCHkE+sQPsOrls2rgWX26mPw
b9lBJHf0/Fd1StjzqNhyswmamjKvfNKSga5NlMSYq0sRTLIb013E6ET9oagE4xxIxZn6HLvqjGU4
d6oubNhkgeWT8hATGd6OvKTsFjcylbAV7kPRjDzeftQI86YH9ApCK6PuE15ogaZo7aCzEkcUGJAi
ud1YPDF7DoRmS/zRwmY5l2CmWdirp5vxb48yNOBFUsjYU2VW3svJ6xUTulQJ1ZB+aogx7A196sGO
bIVKieImICBUrBSz3ZWvQjvei2KkB4Bh30f+Cj2d3mRSMODxnb0G39NgKO92ZlV+RH+UD1Zd5heX
huxWowIkXdU7WLd0yCLQuRTk2azSgVDtO4SXVQgBM2rP+KDZcD1Vrtv4n+dd3liyQeyXkT7Vv1eV
cq9DdkkmfamuRNJMY2bjxxhYteNDdZktAPdC+4ZiN4TiH2SxHGSC3fBfzBrcpmHTm/qqtM6GLB2y
oFXNIGYo8JKMx48a+PFdAzizHlFN/y/fi2feOKgTaakNNWuuNRa4FgbLA5Wf0mSKk3yLbd9guNmb
6GWdIe4ywQn+jsXBIpHg25L6mrHaDbVvq+0t6/TNmklCsft4HoDl4eOFquEEH7ky4eR/Y7vl84Ub
9IPmtXMCTzvQp7swHHQ9xEmySVnWq5hemix2ulilDULyWTgpG29s/UatLulfZIzpHkSWhIkRn3Cn
Xm6DpI4d1qBvNxGH4scnPLnqOhgiPVzhufc0knUyQs/O7Cs1B36f/dzdT8Op1pHI0a3FeFcjTO/p
LgU63LwMwBGy+q7zGnhwoqtvrkaAEe5rxG8gRAFr5nMpa14vSsJhymrRIb+7jr/0BFTjB9iw1oB+
5oidaX3XpKAfl+s4mUsR4LRBbpkI6GxflWy6rzX+dMoErZy+N1pUYXJgGKs9xiXoxL4g0H3PYiT6
UxgJ5sZ/LE0QbSfIFjmXCe5Y9BowZtLV+EwxumT3Sv9T7KQzxTD1j2xawTA/Ky5CREQGYm6j/XZ+
YlGL2y3S0nQRmOjJTLGoLc0iopEdZH2+GcGTQRipcL/oREkKhSMkQOuGRb+AjPJJgeRj9rnp0KhL
rdSJwl/a64CfOX3J/kDumvJRPJX2TroNOB7vtYKynlR267ZVgbwHTnUG9fNQBjPKz4bT7FKdUIaL
KA3SNdc90X1x7TMLqeDezEqSJuJYVKxOOFo5/UembwOlHMxwjuAs5vhW0gUC4/s3TGJU+/TBxpTo
b+FOyPVcMNOTDTwKg/HNeBgC12Hni6KNz809ap/A9kOuGU84YsG8tfUehKBeEeAu6DGHLGx+uF3m
dfuDI/xJz8dx/qaIt7gJ+2gwTX5qu2stHw98UVztTmHjxZGs1c3udiUS4iR+U8b8h848N5O28ga/
s1RUrExFejBSt1kXohyVzpbYBzlIjP5AxMm4DgqjDDce58rupWxs2xUMwvdNqFcV5EVC0PKOnVse
JOgjO01EKKvY3BbWBUoe4RAlJu3PNIw2RnEbvSmW861UJUpNktNL/pXleW+US6Q3wXEZazc9FeZp
Chogu/TU5fbaqbicL6M9a6bAzw/Wu63m073+CwfQ2JjQ3nPkMzeSADa2UqPTpbM0ChDlMpin3tzI
gvRyphwfZFWLJyUcX5IkJO1+Orn+JBXo8Aaf9KQezTMt0v/Eamh+amRcQvOKD3XYlsb8kFieJdbx
GyF7sipNzTjIX5UW/BmmpPm+q5SMWQRjj1k5cKGj7BplWdIfTmQ5gAF58X+Fv53f6LK4aYV22Kn2
QgxrzKaKgbREg5VYRQ1szKoPnTJedFo/iPA/slZFSO58IFSedu/9V3eZ0ITC9AqcBUd4wfzYsiqs
1sk8y0xyxDkZB8Xvhvx0WPNL71HDwAzRhbpOrQ/7WapoU8aWYzlz4s//JBZvSh0CxCtLnXi/NNHt
paQjejXRUNf4UOS/uR8ECCasIsmkfdJD+U4YTzqOnSBRLhKfY65+5CIegvauwDNmtZAH/O9BU2bs
zvnoFGl2FXyZNjfPTy/dIYEEv/Vnyla0M+FEji6Dez+ThqO18fZtaiJczQlbuU27gWeS6n42KCRa
ZBBCzgaWbI6JJzE/eTorhHraQszWeihp3BRhzPIgCNxJJ/IYZHWA0T+Ynwj6D2m2KsQoooxk/sSq
TsU1JPy5i8+hRclT+HL6Vj0eRbdZwruaEBdjr36Y/bFKreDpG/K/yFj+1nzgPnPrnTeVAAli7UKM
KNhQTtm1OI4n7CLPZmDMQugZTx1x2BCWc+pfXfpjoipGAcwnMDDhV/oY+ukf8eYCAks3n4V2Lzvz
S3ZWrVBhBOTniQpoyz8HGZuG8kIgA6UQPvvJgYaPwKpdL+GWKKlSPzL5lhNJzQ05MajL4oLTkt9Q
H2+CuQo1O77t7VrUix8Cee89GqockN2FUJMXs0rdyNX6cIEg0kqeSVIy/mSGxTgoMGUGdm+3XTpm
H/q4ftEXtijwEmBR8qL44u0BUzhfF31OhqMOhvwx8qGxfnN7znjy68Z+ySbF6omPO7qfrVqxdg55
HkUpzwvhpZra+BaBh81N3/RiEVhb9ZsHGrOYYYh/2WGHJOMvvA8lWqpGjNauV0HZGbWVqv4bgZIO
A/CbDxH6XumwryvY8s4U0vdfhfTPz3oUGijZ2YNSqlHi/Rx+FhwDPzn413J/86eXOHhwEf3gaCxH
VGaQP5ho2DjPRFNI5JXpSsXfWdW8Q01HWFoUspRplpQeDliLzbfjluJlpXcTQcGSNrQKMjL29JLj
oVpoWPXnH0PBGkwaEfPX02PqlrKhBne9fFTnbN/bD4HhA/9MFsNbh5KoLpZhv1r9D+ucXDEMoXt3
dBdY96s+S7gaSp+y/V0Kqg5FNvSQf3Ub2cMIy0KE0bzOUF4+Y7AAha00573pG0lGZG4XwdBU6f9/
0Qer+6tHEs5UuXQadsKDiqWtqQg2EMZQWZVVjr6OjAceHkv3vnYCJz+vI6R919cy7Idmfu3Mlmlk
+QzvRwdYvAoF9EoV44LjbWwKMalKfrgAGescirhpb2j6AleoSbkY35XgnXVo/cxA+IA5zMyVo4LH
14eqGjVEmmNE7DpSS0rlTZYuoADPsaosfm7Cu0f+b8FA9T1DjoaqJ41lPGGJOria/6Pt/1r6AR/E
TtCHMvJ/mhMawG2xH/5ERQ9mivjZMB+7xVmyA0oWwXnIIMhoq9eEwPH3VBvofigAQrzqI4DUsQtS
rV9LHJLcEbZC+QyL3b9ZmlIBDmeGhKe6c0OJ1w9UMGpcM10FrCvSq7HZ0oLhfd/CfoQ5pKjuoQJW
+agkwSVm98QJ488UpQxhirCOEp3i2IWuGF1YBXGNSnz8845a/EQoEx/QUlxauoX5G5ZFJBuTbgrW
T4n62XYTz/oS9Ui16x0gQLu5X+MHHh6N4V0V/djdQVk3OsVaV2TGHp/VmO2Op4pJaX9p73KbawZN
wIf8VxUg3tIMg++ROK8fWPjvcIvIs3WvgSBDvurbx21mcaitXdq4tuRP8B160tdIouAH7Cnnvpve
ouSeSpsbsMsyyBQa653jQgcRp3Dm5MXtJjkC2aHhuntnMKrb/GnDF4j8wFNIsIwC4mOu1xokjmiG
p3LR2dhkXCuJH/0ir9flVBw+QUSO4yerXcUltSMzR1jzonvtaCAXY1S1UMm0Rx/T8tZIUqrqWTjE
URmHI/hHrQzKjaLcJdKdcN+8RoDEiYzJbIu8Tbx8l/iWmSpi/SQMp7kujI8Rj33iYUlXlCMcnz1D
w5fviFabZzlU5gZ2ES9nHN4wP7xT3Ci/2FE0FXf0B9vcx0Ce2TyEtk/QBuPugfT/GhvzwrAWMch+
eI1Upr/3S7xU46Wskm5D8WKqSj0VNHZq7tbp02g7p/nMz1F5WZQQgODgC3g6oUrBgmoWKzD+8jSn
STSsKSPozhPsRLmg5NLdzw0wUQ3e9msFHdn+ZWcwJk2UjvsM/IodLM2X+Jlto4BpkhrAG3NMIxKx
NsLQEGEViLwgo4W5sQjXGgu6o4vjOJ7Ic5UiEa8hKcgM1Jdfjl2USlsJLnJFliXkOEqFKD5iCLzY
+VCWY8pvWmIVms8AkFaxjTXly07Wtsf8lKJVqzSXWbUKTflgxYheAEkfydBEhu4I5e0ZAf8xD/1W
EDHSJzPjixvLQViTV22pJLifwJpbTjtjArA32wuK4Jda9XqQ+sbv9nSpO1hQ9T5inQupO+ZxYSjS
Yrxw7UZn2ywrz4HfBHr6zN6LvZx0DE1GPz8wPWB40NmhVTF+QDXv8AzKt5WjKK7fZq1au3ybhXDE
B9ZNb+56XDH+FNSstq9+sHkrDY7Cn6uMruvnqhsYnlomfgfhBRWFFx1SX06OQRmvZN8F5mcqtKKM
3r/RYN4ruGpjtqcPShC2P2iXoEEE8wMdcqot+wZLVR88a/E+hJwrF/s9iN925j3FkKqrSIvnL0oD
uGO08JZlL7XUazDPL/bPzeV1EyQ/u3ezMZ3zlqRjQ9/zA/8URqYzlvZ42UAJ37QxjWcC4QcmQnjs
fmIvygytC+zPrDzdGAm+Mh36aOg+HxGrS9ICQmLpHhNku1Kh2FPl4D3GhgTlFmvJXQuFF0ohwXQh
267s6d4toxQ7xcB9ns8DWVFuBTETn4+TSWui4RGVJ85l4f5QBvIeQHxDAywW4s5kxICmtw3wBU2V
GnzP79qpqSe3TETm9McQ/4opUiAwtD7AN+jjGmgZqzPTXSP7QB91f11Q5CYnFvhdamOlnu2QsZ1C
HG1i+IuULwsds54rCFgQn5cM7NY2EkHSqidA6lH5OtxLBVf9nFRsAJt12iNO4hu+J2fVKOLC1SDf
C2uZfcT++zRaxJvhsSy2JvqhccwAj574wGdWy3Z0H152U/jEaAdccloqkOshnpBCDchM6DaHFNSx
eidt8MG+sDIzTx3qwEDD3cy9lafKoaHtyAnpUoJrpdXAI/Fn1fbfW2F859bVfVcb6/99zY7RDIvM
uSGV0bmP+gcFpEZ75k9+cWFDnpA4iMfK4V5b07YCW5y4J4hV9A9/Yna53IkYgW+LHIM3Sa0XZx5A
EwTjrFR1cayBRUcBw8BApZybSqRoKxQ2JuBWJ1imdvmAU38gGbil3sCGXUSYJ0wOqqndxgTLrXsM
59LWKFnCKc+SXnxiEQ/OtLIH64LTvr+TS1Ic3vb9pwW0pUMSy8zziqb0BDDZYFd6e9bnCV3nmD6r
oGy0UhJAxI2743/ddQ5hd9i7CKAEx9brQwVBTQNMUokZtGDS+RlBEOEF+ORMLcQb2doiJ7siJ62l
bvNm2hTTbnmTokcurXCZaRFQ0nQOTDKBj64dYmzBscpecdj9EefroeZOi+26adNxozXbB6+/Q5qm
BkkhgUdC4sXS6zdIL4TK9Bw+F+Okn+Q1qrhNaqGJ1JPkr09gJS/kUz8zu3nvi7JsYYdfby9ZxaOO
MrMhAUuoru2czaOtQDXJsHhiq53WzBj5hJwPoYMcilqR0yyx8c6zCk80zvhQL2eG5l1sq9VoZZEi
z3ZhQsG+6/RntmP2ArV0eEOR27aHu0U9bka7o8L9mqQZ/NV9r2VJK7s2k7ZJMpuvE02cl2c1qO+e
ctOggo0GFpeyHfCiTAXTQKxI+WSbxEZgSTZIjHet48YG42dEb+sBOcyVYTsuJUjPOdaHxVA3znxG
jDQiDrP8YXcxCxhhVrhLUtF2XBqx9vcAWICBBoVu2mQvtdGJH2SmlHXWyBaBa2ALqTwLo6yvCeKU
1e1J+k7NhbjWXcO/hWorKwsBcRGLCDR/99g13in6fE1pfEpQT52FdutcYAXfxc5YbDgYDNdLhptd
E+fcutScbVsWC/toU9snx8fmsRKqVX7ICooXQJgwEF9Y9gJbEt54CkaWiZmLCLDdVet8FdZr8ZcA
2D4RBFtjSHZ+ANm83zr3AMsjA5HdR1pRBCrgX97BJs8adSq1MDBBAj7J0YQG2kj+2KLMRhY11kmy
jgPIT3ie2/JFv5GdwgFK4XpgdjHxdVB8TgTqrToqokVu2VPpjBAxX/jReJKL3fGO6e16GQYoZ4sf
8ZcWrZzSWd9wXMMicVTCFyzsOiemk4z2wcMAE8ZCTTaUO1CVGeu4pW1/StsEC3HiHujhn9n5zccH
B+Jq0X+QhXS04vT4ZbvsHROUGEQL0bLScOCknVOYsnAqb0kC26PhLxH1ue1s5bWGb8+aXv8yZlkT
GKb8l4JnBYy5nKI9Yp8ujhor0LEKquLgR5sjB2n+Wvh/k7/oy7cvpU0+bwFZh9YTAX8d/0Mdro1B
t45OYfaPAIlwZAkmWTNN3NZm6Zt8e7MEe2PWX880pTEyT8Yva2x11D13zKpg/mQAdHlCOo4usjXQ
IyZ20DFu3CT7ygZvv59l3NKE3AERNpW0EwiM1VmaP2TrmfP1pvS1pHWKuvpyhlsk/+4+F++Z6RbN
5dEJSzQ3RxL3PTFMDvihxgRQWOA2oCnHVrB/XgSC7AA2n/pvw3+mD0omSZX91u+HLlL15fTL2Qq0
9JvL7IkL18U+BQQIjOrwf9Xn4THgxo/i4YtkhS5jSzquFqTi+jMSaTKjBEzjSlSf63KFvX0JtzDG
AVCoXdAh0cn9OCkSSbUvYh9EfAfW6aH1xGC9LI5e204yMIGvBg/l8cGX2UTw705A6XOpL0/46JPe
yyGSSqPIITXTRcBpTIOl4NjK6HdxlqdmzacZKd1oLA3RgicyhIHxHDGqVnIeFrc5YXkXDeL/odxz
YxB6/iA7AAmwYacmF0DEklPOEthacr9LbHZLnf9nZdN3U+WUEyC9zztskPZJoete/RUfvPR0+m6L
lG9U/9dpxknmEyNCWJTm5GR443MAZ1/fpDoQJPBleYzlTjJJqJr3+Cx/rv2DfzoMY0yutS3E2aoU
KOAy8LkQYV78Ue8UdIdmIxGzvxS4Tgo3U3k6WOO9ejoa1zvE0GeARP5vBPGAPQXdcEULwIKl3mXy
UpjVVZPbDhAWWsdbBFc2EvMhERAykov2i+lC0EjEJG6m6pGI2MsPEq6zalXOqX2qBL0fqQdL1gdT
z1LODbTrs52Zj1oEXzd+cQ9y2PhokuKBueTb4W2D1zmpCQ0UV8/CgVmA8ZL4U3CKwGvfEpSDr9cK
XvojvMSoxBBWWVDVKwzXrWrnYY6Dqy0SA3s+0XL7A2yGJDlFK9yARYB680LxOe9CJR2smYNZm4tX
5sbnkOvlix3m2JT8IrADOTRCK411I/thDA9oOpUi40kssY83mvuVf8vPoGKoaqXS7N84FOrY3x2y
Xv5OiVx2aTh0aouxlHnHHESFmQ4+uCqj5Sjhp1DoXCd7vG9q0rXbBHAFPu/qNEGtr0tiPX5/yNTZ
gaGlXGJ3L1xKNTQKhaKj5efcOpHWR2z1knZxHmFsTUQxl1tV/wbI+/91OQDGxdf9otjATbmcOpEj
W0K7VdaSLV8xRKOpUlUbvOo2NFprCbFMjmusQzBZl2vcBSm7Yx7fZ45fK7SAXusjXQdRgAMZqEXz
WZWp4iGC+8kDDwiTdfHqmqI2m3eYjV/EDLQrov0j4OjeelloGgmDbBKvxEi3KVBJnsSMuG7nsXLm
ML9kOEApVuv+n8jhKzer+SPgdHcegs8bDc/q060Do9KPXQjS8HOEWvRt0Q1urn5n2c6JdflyqrQG
LOBOtfRcRtcM9gY5n73LvD8ujbzIDybwEEAgJkUZA3k4xv6d0Rohcx+ZpBwmLRnzwm7B4S76lYgf
/wyPp1EtaQ87+RUEXXT8BKsHo3r/EeaYjYD7vANqkC97TBqhvFITrMhCCRb/0QO4MA+S2l9YRQo7
vvnCiZ8sXxGXHCbIh/sY+XxIGwpsFJKs4YGa0qfwzm9KbewcHkCFX/Xq0rL73tsvbDLWLiMRV3Po
ALNz4kq8ZdqJoOOcz0DKdn9gHeXA/Qw3aIJ1pN65qxKvz4v3rmK2TwVSehouvk0wv4x8/JIoMXO/
JWkmhjZt5yzKjRYNOnQljgC5OoHnn/9JC1kiOrSBabLg6RrkDq91N0qKfdtLNvec5lwscXLz2kRo
Yku3TSO2RepSiDHM8UgCFZkER0jGAqqTgDrktgbUBxl/j3zjy4KLDWngLXL3fPTBEAuLWgYS7NYE
N4PCbD6fiVtlBTfk/cM+FT65xPMnkGe5ZZlBwY7Xlzmnt+m/2mtB3WdCejePfTpz/kbXGVAb7/WG
SJNY7kOgPBx81TnhCPhWzksG07ThhDqLfhqJLe3gmijX7klwwhx9yd0ryEHKiWGG+U3tQm9zqrWa
gx9bzoInls1sMghiWCFlDQe+Maftu12l4cju5K/4a/Lhui8fjkqq1o7qZf9DKM67v/sXjwV7P0Ru
JlQD2VuS1PKde5nUuvpKT4f+czduxRBPNtcmeVAZALs4pj3I1eBsujkJBodOoaN/TEbTtAZiaEdF
hFz3LpKuq7PQd1Sx2gaCHxJrU/6vNtTCrGTChFlcSaV1Cofzf2sBoE6JGrlKMzAnAziFV7EIpGA7
6vEzTIwunKA0YqAuKNzsXK3DRP7/MzJWL5r+SyNx4GQXLkQcDa/7r9Iig877D6ATcj+yz1AaatYR
HcKRtuxCUpZ+uX3U10n/QQ7EV6f74QgK9Yay9WBs1bgFH0JkD2NJdOOO87VlqO76kEYskPWiQY2Z
TBdqwmoQ4OBaKEfn6EYZEmp7vHizu9kE+2+KOX4zZ1n+WSikiiPfoAIKRAPDGze66BSVQLM8/jGn
FwIkbUQF5FW2Uxqmy41YlOfJ1hBrPtrgn0pRF5dXd1vayr2fnA+yUmef0coKqtX+/i/w/K2dxUcA
88lERYm4Bs4P2qPQg8gjmwCyLzESpf0P/QjVEWqKsj5OsjL1t2J8cjF27PhfiejXC/MLHAMMeaBs
3yzB49dPm6OW7QcI3IMFf4TI8YaaT2Ikss7AfEZxOhHnETdKuMAUwFsh08PBk0m1/YTe/czwZp4O
AycTBN1KB9lWxMP+lj/WMm2Os5HLLfig9TgCYt9kk1Y7jQgwi8GrICGYSWuG9oNJPFnXUEkEQSH/
+y+NRS+0sjGL31X+5YgRnF0KdFFILJyPn15S0uPF3Tykqunf9IpKfLy5dLIge0rPIJMyoIfUf2jK
VAxotUS6MH7VAmhbEW+HsnJzzWhmsMz5gxa+XKt7xgYudDdytPjwah+QSVpgqNgpujvfRCGs9gy0
12WJrLfgILnpfIWC5J1EskW+KGKtYpY3WUEO3UPvfbwb3rwzdIWrz/kaCU+F8e8tRXEtRt17CYV5
c7Kc+TjkfoyzT5JKntU0T/kV5VlENznRkDqe6T2Kf0EGmT+ClqDNYfOVbX+cykbwXMBs399XD91p
5b2MsmkPY+rLFGXRCZBWlb+0LX3qZu8ThsKapWSDxeSUvyOxDmCuSEr5Hf7ZjNUP3eLvyDhRDzLw
LMdhYr7cSIVWuKu8l+YYVT0EBWmLka3A/jMkdQvYZ4KQiHVGSO+1nkYLVEr6gonku6ayPfAY14Dz
BHCOBCu1lih78f0IBFP2pQOlC0Dz3W0MNnjXEcUqvJ2b6DyD4NPH/oKfQVoNtIW7Zn3XkfS0xOv7
N7LW8rZHJbIyeyQU4Dsjic/9l9YY2oct2Z0FBi0++8M8Yn+nB2fFlPMTSKqYKsx6CvwsjLqn9Yab
s6cD75s6v/D+dFIEwxVLwXxnzcXKlwUVW6HMjxDLqZU/vn6hO/w3dFx16ld6Rvj/hhVeJOUU3uqf
34cOMm0nPkkOJW+oL116XVhMMggzHlXTc7WX3/eqjoENoGFP0pf0YecUIPywyq6FaJuSA2TXWNPT
GnplgvzuQYx5fnuyZuuZ1Q5Ct4BnCiyDHF+0DyO8Pm4nN71rc7szWBkq+TBe+sUqkY2VvB6j5wrH
astO5m1og50dJzG//3XPCDRmfAT7TBO2qlZu40KX7JHA5CTGSq6WEFj2ixgNYb6XQQ9W/PAkgK7x
yiSYVYGoDogGyX6akr5DYs3PcydalNHfhIwWACC/gZPb1S6dwqqnfZjqzERXh4UNOj3crgfln7Aj
9/5YgUCArSvWGNIy7BjalZZ2F2pYyB31GryFMU5OsNawjfQHpA8zZOti47jSYQgQwD3BGDFr60Ei
rae6u9mFktr7KDKK2O4A7yOj90pUjtWx6Sb7O5a6o2mvFTelt0wXaeq9GrpzuMTDt+U8h6wOjlAu
pZrGxDgGoq9HijwmRuXEbd3QJC28S6yFrjg9eBeYtz68qp2RlgbbJlcz4sQOmfZCaxIaS90rNrEk
jOx5SpSS1udFug0Tem1Wro8izI6u2ibP9SUk5NEHkdjrLolwm4O1xOz1CFnu005imTprnukASGNK
MRjKDX/U0Rg+6IgLkvz++GRmzD+aP+h/n6R1WVQ/CH0kiKPlp/GF7Fw9NsrNfkPqlq6kzQTfPCqj
EFLc6mPRVIE7xeiRfStsQyRsCHUHVjtaB1lge+hJGLVZgHCFm7248r4+gAVgf5rS8tMdIWZJnND8
DrTW2mV/+rX3SLH0D9c73ka44PdJQWw91zsrerjdNqqWd0slVxupJPQ3kWZHJI7lfL2EPQpo8GRJ
ufvZDh4bi1YpRt7d5QdITmB13VljaivqwUf61c8rTaQiebPHlnPmPhIWGMPx7yQ9nCrCcn+yhrXP
GBtwSXrQmQZj/xtYQxSf48cKePOZMnOxWMTOJKczDwCgWCrO+ZBLYN3FgRWfIAq0dXV3CvW/bOzj
duEtUO3FuaoJ+AcOn9SuoYeWs3ovE6kG1/X/NGF50Yeec1r5cL5T8GIvV/UkNPysPICIuuZw10wO
OdZcTPtjQIW/on1GMND0YPpLLrPnWOhsRbUG9ekDnqeNotLBGBte15DvMHqXk/2qR/zEZ2LMBazs
pPGfec/fedEqG7p58uVZ0seO4E0edvSsbEe5BK/ua9BTD/DVMS4pQlKik8e11d1QsV4rZATBC2Mo
mkIFxWMuYk/BidcyiorJG7aVubs/Fa6DmPxN+KZzT0Sr0iHqosmTc4l+EY/lg7lbXYcuBdvHxWkh
WZoaCKylry4SEvv6KBOBqg2egBMesFyEbanopwV9oZPyy/GpT7EbT4RBRICSdvucDZ2ZR1lWrI0N
I8mSzMHhCJU0/fzOS4E1QlRef4Nzvzyb625yUSzOh1Fdb/wAI81KcoZg6bdfqyk/L9Zrltna7P11
5rhk/9cjLV1R8im4khf3ggxU53cpGrc4qwi7g4eJlZWvPni+e2Ugsv3MZiYRPFm3oDhJnr3xlCnx
1a3VdV3MfCCXPYS72ls3t+Yv2WnGRn2TeVeMaW1vx/aSYYb1JPik3mdbxLf0ZKfuzz9cS72FwEc4
kndLtan+0+/4mAtkDs5dbxT0VGKR60fTS8JIXncPjjG1QqB2I4t6u6rOtpBUQvtmxl6lxFo0gaWs
qy8dz5OQ0FEDQr4rdgb4fN0S/rxe3tiKJNv30H3gGf6ef7WUZ0QlMyP0LkVZle8sN9qVG5sNbxuu
JguEhypp7deLy1cA4+y/XokjU6Bt2d1H6ULHCWIsHrNE2y3ygo6mrMdj30wbasax9Dl1Blepvr3s
JujkG+1frHJrVVwhSrW7ETk6wfey8h9t1sPABDflWifbj74MwZydOYIBtTxQFawMOmcdooq7R8ZQ
1teS2M7b0jcxnLS6x78N47Y7FrUtFrWRlnBuOpcK9hxyRkp7/jv0CEqOk/ctYOwB09nL2ZW5k29g
+7s+WxOVJ8iv85IO/XLf1QV5WgJ5rwGnTVqRCvtI/o0rk0jn3/csmeq+G3waNllUwaWgETN6T9PZ
j2SyRC5IF82ELd1ivWEG/452qWSyyfBQhzXjJUUAuiRReDHjxatjluxrJyBZj+FzfyJi9gu2NmQ0
oB9/SDwmw7oZQ0BLcmoVVKXLazg/Et/a9v7I6mepabVBqKDun2BZOKOamCUvcW0qM9tDnsRBFwLZ
hF9022y5s5PmLoD8K8ZkdX9aLSwS6vs9knPrjTIg9ddn3AI+O4eHKwbDcKDYBfHfUgdC4UR9Frh7
kXParbIJ4pG1tkmZr7nBo7CMYew5OFKmhc89eWD9H2WZjyUDzjB9ny1RZEU/MynRsh30KwKarlxl
qyWTcvOjBiLdsXo5hSlvhRxyTrtWgDp+oyd0Pu/D60vXCgZRiDt3B0Z5xE7fDWgdlMXPQ+IroHgn
RdsqOf1pnQiOzdBm36tYL7idS10/PvuqEHMA1YdtcwYCLi3Nom/0vR6ZOtrD33LZDEmu6iEI8KW1
xmZzPbERHv3TkOl2QSehTtBnsRh3uPHFBw6M36mDfRkd+qQ/pvLoAfvV6Zp+t0ClJ3Bejht8Vp+Q
Eq0bNKbV59IfKmZbmgzTAQweVQ177Vac7RPsOQ32a7qyJp/B8lMGT2gUWabh+Fmil1l2ontIXpBx
jiIwYEVLgcMIe1G/jnVTUUF1F+O4NHrm/WcBIklYYVXHFZSIv22PTu7v/8TqkvrXjrJ/qdGPMveT
x3GBoR8LS4CYOY581jpqK0m/lklskwVM94CbwzDxwXEPvzAh5vaG7ww2xWeZgfrAVzXLYabXoiif
tGEal1mUbBITR+Bs7+/hP+QaLjFN4j7yKx+PgI5oELJ311Gbg+iAbVlUBCFQbAnLnZWM1sH+8cxy
Bu6hNn9tONNorIVDwBciHpYlGzv3Gcujg+C3dO4N5UFcVKJQ2cT/ue4xncW4682eBiKm1KS+vpkR
jfif7v5CrpTHERRJiUQRRV1vqrLoGHCTPdCZXa15NVMEiXL8TuuFE6cNjjvHYJ4w1LNc7l8FYlTR
PTYMLVtnGrKhVMRtw66c0ZWXQiCmyPvLFbO+wQoudQs9Gq2hazaLCVLg+isWLOHLOXSj96H6m+LB
DJqfS4j9PtHCBMAXb6kSS03oOGwKrb1xAHQKY2s68eEVxFcBcIsV3G8+m2QbCiImd1HyFqpAgM25
HTm7xXksjard5W48ZDQpR4bQm7iP7NZWnUGyuThXnTtNmt4wA5iJo7nxLOVYfnpYQ3c68dpx/OZ6
MpXVDI3QoTqLtLT5gNpT7LNguAa30Kx7YONBxEeQ73FjTfb5tM+BKGQN9OrHnpnTejjQW4bNndge
GVJI9fWNLDaZCx+YA0cMEY649GIK5iynJtp5xNcYr7ublGeBJHUvEWFF/GSp92IVuulrR985OP6p
Cto6gMwc9TmV0yHuscMc1UJWfXTz/yBWbBc0ofq+xKr4SFMyz8aU/mF1jN/35ULlG55gua8+Lfqm
R2tssdHxsQw87TxyQcXdvqSDz8qFmVy3mj8+77d0qURJ7cjsoxbloLRKlhCFJIqHtyVdA0Rvf7L1
eHHGejUnuPIim7Xy0bo9eXPZPmgWrd3kN+k0B0qtZ6wZTP3r+uHlf6zIpvN9JQbxMDdUUeRCpdAt
mUlH7omy6P3JnNpZfBD1DummCHeWXoS4AKLXgdv0P9QQlnkNKE+tvyGp+gJXmDqfJJNv6g9SYFhl
Kbv79EYJKWiTLM2lomF78htjzw919zhHsfxAA2ayAPAP+61LC+vK3SVJD0vikz6tAugXTnN2ILhF
cVTPHzilKfHkPgd0TS1NVebYioSoqq6aAa5Xh0VKHUqdQj61Kphxmnr+Cztt4rjNNIGmbwh5IOt9
wb/wz4A6yvV1+9oReRBNyJX+cc/oT20Y67XUWHMEfmsE20OoI4dZXKIFzSn9PmgEG5/liaCBL6Pp
L56qhJMNkcOFVAt1lS28vobHsgthjU73rbP+yXAkXRJNso70CowOG+TfsvkZqWqyG8Buh8UCAYtR
+90yey9p+nsK4/FoAGwaZDbTqvbmtHQKPXEqQ3Zfxh3GvKE2zFqByzlBl01WEpBqDX60Uuq0elvc
xU+0WkluqlMxAurad7vkkunPIxm6KPBJnAhK1qSBERi35xPdoRAkghmYwynQsMjb/JKHfG7R4c6P
UhPSdx+qtrl1+a9OxUK2m+8EqXjl5x32TgN3CIYMwjnAONifR8qjIgsTAYw+3KD4ZVukGZ9jbrJT
kDAUO9UIekyCwCqOhaBU3nEvMOPfQbS8+YLhvKRWsOFBqq5LPdB4606pxT0RUV5HNPQIgF8U6rrQ
jP7in93BEK/bN2hTEvTft5oxjWzYewyJ2PYZ3Iy6vwexsOocVH3iEDLeigF2egGGPBHERq6t97CN
xbD7fnvp/ESymE3iSwdhifFD+gsBZhA5b08n+Ar0xIgiqyCLyrkukbfhli2p8ifpRg0mZtnxw341
0jeVgfzszN3vGYRczxNX1gcJ/ldH9ibmLUbDacnNDFwkCOhLkwi5zWn5kFXCghTl6BMQHfw8JobK
K4HvxinWLR4tRF3HAdJhnR1NSJfCu1LTDerM09WNpdAgcrb0hoLL4OuQwkA9vQhUWN48j/Jcq0OH
M9bVPns4LDXH9OHlOLHS+EhH2HnLXVIfvvSeBcASPJygoXDs10YvXcN/L9awVAdRUx/zd0eVb3DS
RAXt/nliut66Z2XWKClpwU3F73PIRW16+i0INjDMlWrOk8PoPLV0kE1U0JsiLNoZJ1IY1MTk5jyG
cPNbR/9g9PdOIzHjhJc6s8QvJOWS599Q2f+tuG1f8GnHeHlUHxb1IYq6llncCzBFILoS7yGi0il6
K2xMS8rA83FyLby8K+/oDYDPk0NWwP2O3p4PIOx+6xYPGRxYvjuv4aWekGzDnWvjPwtKbB9NXb1J
lOybmDWc9nhPFkHvZJ9h9u0jI6ISuZOhIiilUKi5s4JIXenA2yZFq0Qh76SS3M2C3BuUkmiWIa3q
TnLTOJFuMT6jBQhPeWkzyZ9TKbaBIwT+Gnvg/OmaD9Yxnf+bDnRpkd27f8RA+nM3s1mO8F1FkhKY
amT5+zc1Kqj7cytYPHM9xh/B/zzB/jlG3o0DqJf6TVZ+i0lmaDEqsE/HLhFcuasbFNWPX+Cb6cOH
IQFjmA4Hjt3lrq4nZrP/cOxh0270G21vxY0uJ20v2+mtQLi9OwLh6S/b6/oRthMFwTLFwPLfC4Gj
fexdW+Pc7hOWvXRfpJqbUhiKpxBiFPdIUA8kfIy9NW512bL76mBg8N6tFCU7FD94m3EGmmTjtxsf
LagyZ3FQAp9WG+y2c1WPUNOlM8lfsQRIrWgGtj2I6u4nQ7SZRD/ymKxbnR11Vr0l5D7qOf6rli//
eDbQLPxe6dXJu0eWdAMYDNMfeYr9U3h4G+/ur+RbdJfy9G2pQqyGGgqzF1YSR9SBg9IWbJwC1GQ9
tRY//tnP5peHQatL/HpnIGX191+YCHoud4YoqIunwXq7dMvFFEqfF7fpFe2SspMHoiq6wg4dmLdy
6Ey8f4QzSZrbWubtTRweo5hHhWIwv4dV31MTPypLUjRt41dxhAkS20wbPqQ2XmiHm7ITuPAyUvKQ
d6Rm24DOKhS5vy4SGKG/XK7CRaaDQzFbNXnpzYzTOjI3lgL/OVSRMoHNroa35BfSjFX3zmRtC/9C
LC17tJdWyPPSIWWcX00sw6GgIfeTH5qtSjdunCE91cyd6GzvFMsnSOj3113rJTxjy4iRnGz3XBL1
VMWOYqEI4NEGzR41RylNdmPXwhlCsaaVFbo2W6UKUACkhC8W4uYB+uRpvsDznxE6Ay8bMM5Nfztk
5CWcfSE8TkHgnJM8fbwpjIpvjWCJlVlgnGe42n8RaMC/ne7HysV5g3QA5LMvbFZwMF4Zw2ziA5T2
8l0tnzpixCIMQPzdD1B6Mn3L3oGZ8wif4BIwf+xlJsEHEz/1LkjB1S1PJXaOaw+FXD9jaEAKtCHA
Sx5FVrsBBSOrXt4pWK4WDOKRQVPGcRq7uDBqQAY0N2qsn9YT55RhfQmKqU2x3KVpjq9TBBLZmxKX
OoDXcQ7H7NiBaNrLBhGAEbZA4y1a1HTxJoU9FCMlGqQqf1EFFw+LZIEBbApTRWi22M3/PVxLWNiB
2HIW806koZj7pqDx+MJ9v0xZu1EqBVHS7TGgrFrkLSZplA5iRq1ZxUDRTWF6PjmxV4qbT/uuUTeF
IiRmvHa6b5ZpTGgdOJnmUr09S9pPR+tDJUm4mddVn2cdJuk4Y60mMIDcHSWD5QFjCk2jd7UlkRm7
hbJ5vkHxBxtbBCVhezPlDjYYhTNdeKh+5rF+mplppd5Wh4hyNnjL7FGly4ErcMp1q7Oyf0BctZCm
S1kcB/gcyxtIgNktAHJ84T3kKaZ97v5b9J6vTNn1OIlQlBpaBnCpltWGG3LmtZV5OHgNjQ8ch7k2
Vaq/8qK/DXSOZP12gdPV8lQMumbZqZaYg/2DoZ+rMF0nWC2ORVKO0wxbxY61cnxpRsAY6kZ6SMGT
wGRboRTuzJ9LRUIkVgMQyB9kgooIUqXAdYgGFh0KpsA3tkThW3mCQCKpYMk7BlIymP8ObgczDyZt
BqLytMjvfwSLLW741DU3t9Q8iTffsaPx+FwH4m9m/xdStfrA+/Z4EmwS3zOlqDkGb/njNC5iUssa
fa+iqRTGuLLRwwF/DD99lsycPOMKGZJRMqM5ozpaXBdFk767mtNTLKn5XjeqneOtlXBElg9FqwVT
3154UqoPKMdZphPxEkf5mdxWGEn45MZ2oxTyYj5ADGgcYqqqTR9CRi8gCExGpESEDXOnInAmnPN6
bJlJUnLcPTD7PuiW3OTiCCtE/wV7vWtd0qHj0VR756YZ7o/uRFHvA+fNXtEr0ihSVpv8ZTgspph+
G6x4EFmK/Tc7otMH+s5a+SM3EcaEilKsRCIeg19aOAD+k413oN9wTWvigLsjiFJoTkdnt9j0nUGs
zqruhGMWft/6Efj863mtCHFAvXZoTuYP81YrkG3aaeJh0ybyFq9+dZP6eo8rPllQIVKdClDJkfdz
+XfVbZ+HN7xL+/KQnHNBeewmxDsSrc+IhiBpJTPrmY/9K2Ph+C7ch7gXZrFEHNSLq0LufHbSUuBd
gIOaDzegynlYD5as0KXX5LNrnSsrBF83dwFxCB4z3GP6RZC3PXha5udCm1zyxLtr4LGTwSs91I10
vrXZQAIE0hBS2g5wC2IRYda6gmsDarolZFWDMWtB22tq6KanLdESOBWc4/YqQgIyq/It/0LFaEGi
ekApM52MAR1LQWsJQkynsu55UMH886+2cbYAYnYV+6t5YBEe75TtaOK55n/qa0AAAF2+epbHQpyd
WoYcORmaJ6kDQBO7S+/MW7tcRX0ALpYlgR/JTEiacEPh2CyV61tfmqg2flv2DgETb/V0A1ibFM7c
YZQwhRRabZxC8h/G4yrG+oSWnmcwAz3XMlHVXUkMhr/JAXSAxhZqs9VqE2iAhqhx7ZA5Ibe4iRvK
z4jgpqPisjlK54jt6UqE8fnwWpHsXK+LGqHLWwNfFDKeRHZ3vWGd1AXlx658NrycWR1OM8/6RLCK
lQQ8tvqlxKzfvk2BBd0oeqWbX5H4RmIaiH7mUD2qGWi7EilhsVuo/iWRQGD97sG3XqYmNvhCfKtG
kAJZ6lmduPUCbSNOJNDzeCoyoe53bVOv1/EU00jg8dMNKnNFroBfJWHrl/HAJyllcA15fgnpS9Vc
xecSK1mtKyz0crqDbTcKTtJ9+jx573Iip7Pn6hTglX/2GrUUpyIOj/sAemT3q+xktUxDaKFSy6Ex
ZzD8kB2xfP26+lxv35pJ217QPuJogLEjYuGFojD4CsybaZBBnLRTTBQtl8LJ2yzQZx/AwwTU2J29
UUPN9eLgRXWgFuI1OJ1Hp9k0PTaphpB+G10p90hq8i8QHkoDsNIUhW5PzqmN1Cc8OnnDMrBFYvuh
j60QGw+Mhax/UPp8lgMrTNVvUSPh6yly14Vx3G8MY51MFJ1RV3Dez4duZ8miMGDhQ11ExqEk6T7+
Nnc3WoBZIwm8RCWrTjRiG0+EexZlM/JlNbfS6sXQ3Runz8DuDFDmD82mRFMPGoOhiio1sREof0bs
1rK6cr1yRLMaG/Pbgd1FpjjkMXiWn3XIlUJbPDil7UvIlIaCMIja0vVurjYGmZ+xU0aPkWG1C5Pr
do1107mOXYn95G24GCJudxqOz+0+t4stVMWAouI2udsZDnoCkeuH0WcIs0KMjfvdl85hqmQFHziU
yOqly4N82JU6ZwDl0MrTlZN81inbiJPlTE7stCbcIEd7hRxMiLxXvedYusIzjB1YixqpSEEHKRFv
/uHnS5XLen4iCa1aDaJqZQ6vrf6EZgBIETyBcezHiP2eFW/Ml0rsAGlvEaSa/jtDOt5HNoRMLOX3
GUE00zv1c14vBLzj8jwzNs5WhMuANCHjzv15UllbsXUNBDvaZDp5ZNVxjL8OuSQguPZHTArtgh/9
OLXHDQ2CdqseaYxM8JZq8QoH5F2jqP7hvORGc4rnzkgSYJ1pqmR8NA7S5+LYJwaXyFl1TdIFPx/V
56ygBvTcM3h3TmSFmz0kN82gsx4ULKVj1HvFllc0WypZcErSBGKl3QlQv8Z41hcC+KtX2t1ihylk
2XWy/KXMKXznESOaMBAK5OS1WXQtiYE1RWXsF4Wc3ho6omPMyAelnuZFaASA1gIXMb/NlFQDHGj4
0ILoYbPDMiz66b+mCb/NhPeaLuMboP2cgGXcHnd5alCMg6ZO5sREQAn6w3cav8/Ledcvx30wCaAL
qJry0x8fNUnLqnB0Fp+wF9h28qzCMpsafd5cw6UQISUdQi8ZVK68V9Fs9P/Ta/7rer4gao342k2S
7KYnfCZXDtWVRll/JspeXLSRyQb2Gsb+ktYmAliJAd/q7ofKRzfiNloQJD6SbiM0j9SYkVMlTMEx
Xc1B/Dvl0QwcFf0rKHcpMssYoP2f0+bG5yCHG+9zs9fikGXXSTLUwHsNu6a0EaKhNKNVi2sgDzha
WlG5yGsWPTxbsmcaeyF2ixr+HK1ALNWZuL6c70//iNpcXpr5VBojdsqvaWy7O283tailSBDHncRz
Pm39BSY3gwmQIa3xVXRJC4DEkTCeGXHhnwF7DlXrBEyaCCFtT19/YV3dKCFyYuY0E13dhQp0t1p6
pKvhtAK0pNmxKTe0S5skNYSjT5no+yKBw8zjyF7rv64qhKltUEv3XsjVVcnUOZMfw4Kw58JgPakB
1ODFUf9sfTWBZFoJSm9wZZBXwhgWUhNlbyFancgr1WcjByq07m+VofCmBfLB1rIWlVvS/d9Z2bDK
QDo93gjkeZnp2DFUtmNy6f7EB+9/MWb6lwHHiogBcZfLkwICZGkaKNuHmSNweC3/CMQNjUAnMQms
WfvlCaujs8oPXzmfLVxuzjY0Cj98nqr5B52mW1MrMSpE6XELXojtxdmmNvT8awj7k1SGgVBzIdJh
CeQmZ8ZDCUwcGWEIJ/nWe8Qu2r6ZNppVGV7h2t9+OxmQvCg2jD/BpVwNsZ10CjIIkSF7dXzkMJSx
UBHOcdQXRoGL7+u1jiQwn5KPWk95NvX67b9M0xUVHtedtGUZV7h1oQEWIr5a3aS5tM1wxSEsh57f
oM5qFmr/nzhjrsv1JPNgWwamln59ac4NmqOh6derq8q9KwABt65fGdWGfZMP5p2g0vLGwMhZGs0e
CMuOCyodLEcrnYFfuFvny3xA0Ic0kw42x7YNQFq5nyKFq7u24dopIVj8xC4Vw/L1H3AOxOuP3KWC
3EcfnshlnC9yl1l6p77pDUtHJXi66XdXnJI2RZjayiK1zXcJNxArYz7eYh3zqqmCGrRmudup3aOX
TMBTHYaeTgqaG9TQTBvG5aXAIKGdhafyWwZDZXyY0425FiBAXmvOEwfkH7Sgfdro3bLxf5iN3zs+
sGhABq8Cnb5yirmM99rkilM4Lk+7r37sz5E4bDgHMhPJM8VpNX/sCZl9rqusWVJ2bdwC6l+89cjj
4wQkdyyAqWjDD2Bl7u+fZouDjQk78hpnVnNlUmWzx4S8i+q93UjhKPmTd7z+ssAMPUawLhVul0hf
f5d5y5Okq/TJ9ZODg1m91UKmmvdUYkV6eQ++uA7QIm93TwGMdcNNTk1gLhYbK5Z7cR+7Fshh0eRB
csAf8g16Xof+EEs/rNztFpxdiJW2p5gydnTHVyue4/By2788Mv9nv91ByV8WCSuynTnJkC7D//4Q
O4acClnycFoknJyCsdnkpMPnTYz55ythyZYB1MxAciHwP+3vooHI3Fsj4WWxma2s9nMVFyNM2jVw
me/R3jWAaTrLWeTiGN+oWglYB1pJhSXMay6+kyRXnFW3/wEykis3sK20P670AenEJAjr5vSDHnXD
sC1yOSijJwL4ki26aIRTFVhTFgEAQmDj8NOuy1wYfWaP5QDpwpcPwfsV6l6Dp1uR1BJ19rWdHJ3r
on5CpMpulUx2J6pQYOLRUoYEFLVhkj0QreYQITZebJRewLt/SvmAtJ7ApJpNmdcEULbuKZMxIpPV
y6tePKBvhbH7SshScOC3zrem9NMYX0WvXWB41oBmu69L5VYi9wcN0UhJpxllBKlzAxardCollul5
SzhmiEL3PI3SGboWH1v4T50mxGFj3oNBl7MhMDBtaoLxO0PC06K1I2my+AJJSRDW9r2WzQwvpAgX
e8cWmaBySoORJqdf0jKx1PA6CsWCphXxUMSCHz4L0pXMrC66TDUAobBJ3GYpVFnZqdNCR7kHYmL0
yhqKAGC+BgOF6sMdzYWJrBOfhlspmClwqMvnGwOzGOGxsSigV5wAlAalL8FrxxIDCiKDXrUaFUAy
RT+0fzbHiqWoFzwVsKBjy6HfvjPp0Dv9dheAT2tQc8esve16NzPXtpmyT2+Wk0+4yYmQGsf6gGsR
NAcl/Hj8jKpiZgh+Nkntil+NeumMHbb/CQJnodMNykqt+y3gWMrMi9g5ceD9YhxBpq24zxaDZiVy
pirlEiEu5Oh7xsHES9Ih4X7Zj1+3gn5T2wS7yCOzoHB3Fk1ohUL4eU/fkgaIwD+Ds27Nq6DYskQU
2+WkaRUrN0WuiAUNPFAD4ocIhSESFkAEkwjkVwUKWiTnY/ZhSjkdufWLvH+lwGS2SDn597S1GjO0
F7sSOTlMP/aA4Ij7U4vzVuiyvhtf+9HvtbogDejt9QpHI30SYXC/tJjUS3buBDcVlGPJ9XLW1ZDU
2wfskRWEKQQDeE/7cp2kdsi2h1OHDe01z9vNIDzBB07LtrEsYGh3g4WcVTyRERn/fkv8mTCAvB2I
HZjNettGtDAV0chgNQ9BT8lj22doBSfCaq2VRtbG3pjMMvM5WZr7TMPHmMaETywsaHbHLuzvOH+5
FjJXCkmMIlAXyU2IAz6wevSV8JRH+G3CiyWQz31hIIh3xwXmTxQHcBoSjT7AFPF6pcKanevsoJHC
WkEiJMKwZCHpzI/AWYin2umxnRTiS7tccpijoEOR44ztPS5KHdMXFoS2132Mb1Obj1BfUEodWizC
Q6U54eX16R6p5ZAP6HMCg7s7kLQPi80ZzzqMOHTHXL7aEyC4qS+JCP9yL9VrbkCAwD6Lc0TiSXPP
+QSzY57duvT7CJKWDRylCaRBA6+Y1yRZyKgl+5HSZ94mGRD6VDDFtP9jA7jtG66/94X9NMbYTCmS
DiN6mqimPBfcH4mM46CG26bYMZH2O9ccyXNkscgnVkuvgDOvMQbGn0q7QoNJXACXCNuS/zfEpdWQ
dsr4Ed6XZLLSYH9PBz94bD2SRL38wrqKOFaXECJzSs0l+KS0U5Vip/0MyEr1KJP/mXr6JjUncg9P
LUAzrZIimIvtymZ9ifAgUABQNVWCaa64D0BM3dnYlC8W3SyZu6R/OomsF2L40SFakb00Lh64h9XB
NX2IplHHNSSWbdz2Tb1HIiGR1yS8TqMdo2mdNUDVYaEtR9rXOugDe5+KiKXW1W3vndFWBUePCg5T
qhyvyq9pTfMoAIwSAIO7n6kEZ9G0YRuBILfwgdFsilm91N7avF657R/5u0c3xTHEPAWQ6yoZbHTe
nktMOCe2euowbB/wvaWjfiMxa5a1q0LPuHmN9/jH4TQhU/2zZ174XVojadS+OuwkZSFFKj6iz/Z8
Ffnj1IulO+clFfzn6+jrcp6yFHG6arnA39v/oSMY7WsXJkGf3BqLPvNDZFIeF+vnjbeUiH7jH4nd
MW70de2Fd0W0xImEc2ss+a6hPShu0CulbBo26n+pCQIR4dA8riJAoMZcAAuDuaBaSUdWlcPMr98h
E8w6kZ3pBiSPNcLY7M2uxuF7FedJlMp/bjc8q7DzueB1IVNCflabEfU2XdAG/owvhg6fShyXaD/a
ygczuwZHEZytckgTs0iQEo/cPAQM1dx1eTPjlCOOtjX9lty0hUT7NjvIziMeSQWepPu+dqjjxsEa
1WpTfmraTFTBtyisCk+C06bgZT59aClNthEUgpb+aKmoVFTdGtEoEUL86B2vUfWndi2w0EwXe5bC
zyMzRRk8+RrgqI/Ep1GUSez37mm0SE2WbY8UPs7DKQI5VhI4jZ/T1RnVDIYNF/6xrXmE3+DgtnmD
4hSB+ODMS5WnjKJp8oVORWwvBFgjV81gOgBHm5PV7DrHr8N0upG81G+SPI0xOdhexUoeyHyqXOER
kQ0ZWNvzqh4qBYwEn472ySi49G+w0Vf91gAKA1Fo4spo5DvFtY0ILaTOtIX/0yQNED8qfO/YDEUO
YVaSid5hsc8X+nJWdCCoZhbjPdbFQ7xs6VHRI1VjIUTTZ/wy6CKu/nBbuFhIVN4WrCcCBHvkY7uh
+mgGunpE9vPcxiJ5OKGQ5ueDixaSdyMSWK4AE8NlNMI69TXFEoYgEksv4rn7vNbTwSeoNQzk/8QZ
kORHFMPegbP33ufyAC8+JJSS0sZKPWkRfxE5Hx1dPQ5+crguYjbqnvz+zgr3pjLMQRUKqDjkWtb0
aLmCJaOf/7wxgu3Fyzddr8XF3Q4oi25gkev8JNR+NsJANLJv4D5ncwjA1lUDHjaw+HY/556c/PIs
0a6KNlDkjjh3YI9/zlcMpgXdoJJ/rQ79oaMh2wzF7pCwdUVSviTVdJOwCyuysd56Xg1IZuM5EJsY
0FGLgyxcUoVdrr73WfY/aAcYOaHcOWQYWZpi/oX7janqnoz7mn4/hDVjL/CM/xbsVrJdFZe2q5J/
z1JhF0ZfIPFhI5Jzu5Qq/8zXKl918dZNvl49joOk0kAorMUPOjUdLFa7Q48VYVWfjQNKn31mFmUI
F+btyBpFGlUehG9K5d/mdKXhyTOTrs5GWu/2ZFc6rb2ss4kOfjyIXve5fBZ4yLqMTv8pG1SAHhFY
F4vGfuW90eANxW/GfUKJjyESzWADszYr8L+9lfJWJhTKp5F90pQD76GQIyeNqJrzPGyOrhi3phZc
b3V52Zrzg3B41CFg6lu5IJ8RIoRl9T6ao+u+dBJyB9mCxobKvMup0Hqeas605xzEL7uxvEGBoL9v
kN7/m9Cx/7iO3pxn4IkEJV2uQ3glPVlBNZnRGNwtdBjL4aS0wRTTgpm9S5LrFVp7+ZkGaRWnk48C
S4Ds+GYKotbaxhP2eahfwRXjAoVjZqRo05Fzsk4hwp1xWaImZTTLgca9YvQoFgoa0lq6f8lUfQPE
Z8j/FOfjYQhLcR/dQu+m8dTf1ObkxqecPaWmSB+7M218C/b9CfYc5a5fQTCghrkNlWWKCq+Jzfyn
MOOp7tUMmWsGEs6iykv8dm2en6hfj5t9RvwsFouHOA71TwLisb6ow0DGAb7d0epM8zHalNve0RYU
GK70IT3PMThm5T594rcdNlhPd6p1N7CN+gyReQruSJB/2btHhom4OBvn1LW1Wn7ShMHF7PeV20v/
ksKHn6ZDJeot03xoHdI7jKOkV7pazk4yJlAr8XQuA+9XO7zaVArgresRLy/vgpAEN34Z6eZCpPAI
KwHSyUKDZAU67Mqs1c+W/qIeVCSX/+cWu8r0d2jS8vU606jcl6LVo7RkR4R7U1PNxENNVkiK3YLD
GEU3STsLj3L+zjdD57teAq4F1a4Y6k94yB1pVrM9hv/YgXtCpY//mBafg8euxmIXMDyLxJxNxRkL
hA2UhLwhawdmvEsydKxOwSWHBtPKDq+OzTfyPz62PyfrQjbSPHGooRKcn+7nxkm36/UpOFjIJUCx
hcrFXJyUM0ZzMhSUJMMsSYDXfzR+pTV1qnh0/MhHut/FtsLQIDYBQmGnuzwA9rHtT8+79EFDwzr/
WflVKVgZUUIZlZFvMPVTQU99xMW9AL9dLWcodxKdYvxXc/v2ye+ucfas5cWeuAojUGXFdwNp0RTx
rTJRZifFHmjAuX8T14wXDFDodUZAtzkrLGTofYxDqXC9ncq4lGWL4qYBfZeDfNU4v1k73//1ncKe
4gqly+c47hgTW4NisMlLaGZXtDwULNpZe1m6DzD7Fhum1Hv+4aOamPzLyTnjkRqkE9bjlznOPr/2
s2ZlrJAGhEcmga2j/bEgV8GMHISbnO1KQL9Te2HZ0iucrDne4uFy1PvLOftPccvABZWZWBFy3UXu
i9+BcA5R5sx2NCEYjfBTHcw/a5qgqSN/VMBTkUALaDpEK6+qwwja18dUP1NbDKQFO9RmGMWvs29N
lMN7ndBH6DJ/GGOR1JMBsbUiULOcIVdnEz38ygDJtChsuHLABMiivYLuTErvjtamCtlla3ojsoi7
K+Z9qlBN/WqFDjyX/1IntQ/yYz7nU5ogoMt+CbYLB4/OUKPzmP84GhXMwXqeTOIVfaHCNld/laEP
gxbhcUdWKU8TTGSYL1xXiuzCg2Xd4zIst1eRUwN5uxCiflvXlywZgtjXcqwyiGd+vPMYD8juamU9
7UVilHMnZGPgYGJmXXhremieRmHDnETKRgrIdI2TJQy5JLkV7Zv8OHaL0lqwc+RGR8SklIxLaH3y
gJs54bpUHT/V10PkjmIJyk8CUHqgF2j16Jg/8rWCcS21N9fa9FGS05mAP84sNJF4nARLeVqKkkYT
zlrgGykKw7w0Upf4S2B6o0WnKFOXulmCNEFmjiVg/jlAoohcDFXU7J5yYVHjg1064zc6vmsFfepm
Qg1bCD0FK0D7ZCygsKfdicR2VoM3nr8LpInJD6qnWwN7IwYQjkdfQAr05iD6EnzFvrO+wBW7eIFI
qpqLb25djpwV4/WmnP8uUYbsophIBw48QEgPi/GgnfAZoi8xmygXvyIaM+4O2N7YQTZgGZEX+Kqj
4/F9BXiaDCnOhpmTYp678c54WNQ31Rq/TzbWPvUp1C9bsWzKRZOebA0vRDUI6hupCSkJvqeHfOr8
RtB3i51KsrnRhbF2/GJaQcYGZNNDbdX474l0hkIVIFbu67XzZVzM2Sbg+6OV+6XeXwa1mW/RXvI+
F060Uh9d3q76gJ6dtr852pa4vHFF5J/N1W7mgpLbZw0M3CWwec1eV8AoUD/aGVQF6Mucil8H5VFj
bZyOCnkMlbOD0P5m9s9nXFNEsxzWeSho8UY9sn29T9WPiXJfU/6Fd23hvGznMDK2gsnQcgiFKhHW
j5OV4xf8+ambxIenY/DyQtfSndqq0hF3pecDi3x9CJpZl2szLdQs9H42Jf8veOCQyruFnVsgj7sy
gV8FX7AN5xQjlLCDitlOYLqF5mJnzaXfCoDZGNzLSW7l/Kh4akXmCOqY1y+8YmhSvCajHoiYRudt
pwM5+dPEbpWTtJmnEe9Imx9AsqxKfQEaVuGE5nSO0/2j6juDhtn152IkohWi22K+8z0WEiXO78M6
rUQymHrJSynMqnp1bfAXLW9jjpsZp/Djg/3GCXN1KsIU74jsQG8m49yCwyqCJ4cnRRK1qNlAEjK8
EOVRupEByU70Dpv3Q+KVUv42i/+d9PWhUld+kvQk7f1I1f4fcBL/SwiwQ99X4RDZNgk8NbkiVuch
Hygy7Dnj6gqEFVi6vugwscQYIig4x5Q7bsfox1ys7NzpGfE1XFyo0wxl/MVIz/GV28K0m5bosEjY
WL90SnTIvfXyjNsqTmJEcz4k1gGupWd4M4zT8pIEVTg6bnWKYiGC0C43rjShwqR/djeI69760yWQ
mMjvMiOt2oWKglHKv346p535iF7jPptqz2hIPg3VfF4dU9OCkwv6lyc9mEZJu5DjHRdvciK5FyTB
xeWIu/WpWkdlSOBDsg8tCc3/mMsD8McTUH3w3fpN+rfo0iJ0J1rn8u1EKW4kivAaRxBjAg+E8c+5
wjWL6oLER18lIalhXGaby7FJCv8AvQ6JQ16TZ+dMc4Pv9VBnoHnyaJKeM3B/JtApFVnZJ7cElaoX
ThNJ1XDSw+fjuazD35/vLZWDX8mp7wlFe0IbvXUos3dg4tw+Aah1+ZE0M+4LUyPmEx3hu4sZRsNd
H10Vv7v/hnG8Sr7h9+nH0pcGHr6b7YQL6PSeDd5r9DepxG2rBlEAi1kDqRIEZZoBYjuw7f+K3M91
Lqbr26rZvXIpXjJ7eAuq1s5Tf/CqTxmXjcVs0Coh7D3BrfGSf2IsdrATpe0FoJk2AbpKNkAf0dr+
U4fxx136NkVzZTCerh2WYMfnbflQ3PfLPBQpKSHod6newwsN9dkSc4nlaCJcBHgwPuNMn5ztQDK2
MsJfY/20ytB88WTSsjkNSrInICzgvVyPktYjtn56M7ujLPELIecuYHwVbwcwxR+HpjzhgzfIsric
MjEFxkvqvW4UyCNJXNcx465Eyj+eY4ZxIeOCrWiko5bWCz2KJRZfGR4eCWOLvDCXjC9929R03ppg
gT7XRu+X/7vL2F1JjagYAK3Ivy1wyFIHMMcjY8UuRPHI5swHD3rr0+rW6+D8R/8EF18yC9EjcBw/
V6hQkcrSvCpacNsFxyuRjfxe4nReS/zy118Bo2eL1vPLKDhBzTBNG4UId62oGXTQFQkVIP3ICcIw
BXsO2JXC3Fpryu4qc829AaDmoFtak/Mm9N+g+JNJYMEDFdGfMa5x2iz9g0nIIDrWsRF/PIOSK5z2
+//VJQYW2Ji2z3cXuhS6Po5L2gb25FDAnTvZCTrABtjKF/8QC+7Rw7IVAb6qh6GM9xpkVmmjX2EB
JZMEzSWfNs1/i1ZqXF3NldesR8KcIXjXVXz8C4QGMOB+fbnAapdrHIqrwu5pnPZx0Vmmc5LqeO8/
jDqLzvOm3W+9FGDtYBn5MN1ybMhVn5PI+scJ2Np33Gt73uG7CEtdmu/KQBWtXpaUDV0Ig1NiXkdZ
eEqzmYdnDrVFWvnwSt6z6vvyaE/jg+gXUO579Rh2nqNKtv2wvSHVlctZFaqZDx+JdKZ1Ha0EBdOA
sQzzzWLZbs//ZanZw5ScDxxe9k9Vw+xmhMs+ne+zA4vpKovcwT6VMQLAyLzXdLuz7pf5L4N9m5ZB
Ji661NKi2s3CUFUTVrEF8fFlpiVL9g7/Jv4d6cv3cy1HCyXUzCpHxd0JoNQ8EEXNMK1prrDtDPmP
y6Py+jbKr9+znm8Ma+bATf8AeYOyQ/bxU3RpcswpeHV64uXLlX3UJRc33YeDnG9cRpOMzlaKE3wU
Bgom51HEJrsqUanTj5lKxylRii6CT2ckuj4faybXzKFosOGm04I2GO+JKS3nt7QK+4VX4LJXhrGi
TG+35TZ0lKfOkmpxQPghqggt9shJDi7eh+VhBbZIXT+3GBTS9f/HXrf2chfyHL53hgtw/id9jCDb
Sehodj8QJxQORUFMm3FVxqmngSXawj5d/RkpNWU+2bF76rBb5AaWwk2pi/ucjVx/MJ1CrucCHAoh
HueXxKR9ax46wPaXECac8kKC0DxdXwbl1S+k+PgRTHGdkxab0KHgHpy5Jh3TD5OtLnk7QyN8L0iS
Vic8G4Ox8sOMbO4qDIlqCtoXLx/Z5MyTdT/CcylLFlI4D859nkDdLjYsT8PCEPyAJcRHPctjs/fz
9OtILMqVJFPmHDoJqCehwVKwdn224JAZJeD59OeHujSSrv8Ly9pwakUwkT85psJTyH/Z5W4q/HJO
m/5IFFI9ZZrt0BeOBAL44htOJriiALLQW8fYmNZIJ1AftKrKKCLr575Y9pRXlqfmpHJQHEBxAG56
RInp1obKlI+Z5m29J7MwRJs30xW1k4uZmi2Iu+PVc9o5DbCXbmAE8gVUbJflFmZGPdnLzsfFEEJG
gZrrWDEr/GlLvkzeSFmdvtrJSsiXV1U/tvV2CLnQCW5xADjf4BudYFydH23C8J/iff1Ix89Pp2AT
8clSoivxDtGqFeQlwvmw9c+F+FhG96iHceZJQBvic0Ctx7KtKw2hfo4d0qom6j0JtF3MMdNI+pEJ
dD/Nlt4X0ymf3ChvVhrj09ezi0ugjkOJ9eJ1tDgUUsmT486croiqnDgKIAIpCAkHQlQs0qZO2z2j
suokZf52OoQWYzaMfoz4GWZ3Tit7TtU+CSHHtWJeV22XSaHEZESSK860c7+VqJ6wOFd0Eoj4EcmD
QSKTSaB1faCJBJd8YzPtd8DL31Z2/0k8KSaNAnLaKbnVVpmtYzFh3iX1KKJTD0Ou4vzUlRkCXFCp
dRHmkcl5MtYxp/QWE5aK7fnpDRw71r0iLEC3UwnDwiqLldTRpSBleAn2be+FQjo7zSMTYDdQyJJs
uhZALh3C/u5vFt18X4wzxzCCCaBaNRdVNcShlIh9UPEnzoVD6IHU4uyp+jMZULsRc+E83QR5hOU5
Z4Xbx0714PsRVh5Ew1u27UvDdsa3z3H6W1rBV95ZDcp60bfPLmMHjW1aClZFi9wYQsf1OXUIXdxn
lXNcmKiYufTEZUpLxe5vTCdsLi3SUt+Bv72ND/e4uwawy52hHaEktIfXyZqrn0vIVaY8Cte5nxMI
hiwqhvgN7aKmfggM2uVxp5Zidhksx4XujJSPvmiqaSUy5EjKPQX9DZDHswUujHhI/+PWQ6YqNv3o
aEYtrgxl9aLpaiVdO/EpHW/QL4emvYjr64iX9IMKJCupRddIdQ8Py/XMuh12wg5Bt8eLuohJhPlp
ryjtHmCWO9DcmpLHY2JySQQV7ehBzBMfUB4slHTaSFQ29qfldkA8XJ4omLK0j+CismmjbjLV0Gb5
TBIkJu1caO/7zVfK9VkzJl4MD+igyO3zZsfFNyVyiLYwBQLISlzHvLT5e7sg41D0ny86d6RrN69U
B196FdSQH9zu4DGv287dAGkXetg79TSwnGQMNQU0bN0E9iNiPPIlsxj+S2DrjeJEITjptHSbIBOs
8ao17OWgRHevGpI5T1PVoJwFKJLj9OsZRvSMsl1dpvz3o4fp9cL8Rv3HSqcw4zY1oLfnLAaA+Ltx
UZLMfSb7+5wl+nnKEFZ9Ict+1Dm+BkWm0vJpvAGuXJfxAOFUt4HxJ7UCeTMGy2b5Zmo0wdGKQrAK
sgcOgsYwkrSjZY1U3ByrsfdjFG9cLIzw4rc7uPEAtbyIA40zoww8Q9/UEoAELOLvDp1xMb8u4yji
kAdXPkL5ss5xX9kup1ybw331gavZq/Yb9F9dWO/TqLomfYBk7bDJMEztRhzDXpcHwLmnLHdHIiaf
KXlu4AUv7EtR++wfTkhLo38vXZEtWSbiDjswRyURA7ZGe/6ia1zXMK04Iptn7lnro8/es8I1dFXo
xKMwuZm/T8Swb386xifNIQ6ExrQhB9y0FUI693vd0MvbvwXTlDDbWF+gt+OsU9bTzqE3SehHOkI7
nKHZID1Hzep+ocGZDFnNIO64HayK4M2lU+0JhNmY/yBzG75usjo6lpLUtBJRmn5j+hF9m8nR2LCW
TiNbO2bP3b9t+z2b4m7dOQjjleueZ0Qbrn0egcUTUSxUenQU7B6E0v6PuOorIKYSXOjOIUVEjg0d
hTUHeZ78h4zQaAo9P54jL2fXRL0iVqwmcfSACt0hIiL3NSIjaoz9wHnis6rqoYt6GXWCXoZBn+p8
0dxtEtAW3UrBgaECC1rg0egRNerecYpgdPx16+arzDg4pnEP084WUR2ZUVld4+bQtbudMCRo8y79
PNDZhcLjNQnAZV+Z+EJRqN8RIkJ/JdTZ7X+9t2O2v4Xyx1z+0lanAjBqLvmjTzHcs9tKf0WqbTbb
reTTS8UvrGgX+cqNkO+YAZKFE3ZmBfoZi6PDpMWjIy+YV6rUyi+iW79WymXhD+mSiqhMez32pFVe
u0SA9XHbddOa9mLNPCdbN7eq4Bawbj6e91zRcJn9pxjLnS2dLDYV244ybph57cTHfEbNNstfJ79g
NYL9+raap4GIypH65IJcg2cmwYBVEz5NPRSqXBQGrDHu6cqygGLX3L7YpWaBqoI7xMaKwISn9RyX
lFtjiJSznIRe9AYFNPvJGB3mqCHcaFTtkDFryOyIapOh8ZEveQociY2u5ALlidaQ8Ee/iRH/pmmN
wy5WIZsnaKrhbcxsUx0Ke4sFGZIQ1DGQ2Zt7xyPV3VENI+RpmBWC5VZGYm1L8VK/FpwH0YSsS4qA
V8yziYyFo3YbDeOmT6u2NtETf/x4mEYU2c0Rsp+kmQjJNkW5sFLQ+V3AOyEiZI0mRicOq7CrG1Zb
hFd1EVx6IZgpeJaHrEDCI/tR+wXl0QrcdNLryQ54HZyWH17nH7It+AQcCWbDXZttXJTFst13QTLT
RlF4sxSx+5fC09QhwLUqenmyViz3SW/uQUgluea+DcT2h/ASC6RoynjeXViBOyVfetVv21oVRSKS
ve252/OFirLx4jWEmDflRS4Nuz40pfKfu56xzHhxNPLXkQ7ufqc1KUWcmYYhypIwgBs33SMHOjaY
omvvHWoGCFMo7xntXcVYtB9x48VmPGB1FUMyec/ugH8euosBtU/xY+DwD2gwWrinRftNx75gLwVT
weFrBLBvUIar65G4i7y85rZ76tUi4z/TmHiciIoKy7ASlpSQz0KPvch3afKyKZ3eboxKfuOaQO3S
azuAYOCzCBNouemubQIgNVqLRdwiRST9PYtHwTkUbGtgNet3sRpmQj+5UweJMIRJvURvWoVvOAug
KVTetyYIcTnrEVrqKwTGiqGY/skIBMGCb241k8Opk43h63k+QMaOq6/H9v/aTcLCHywgtXEGdNL/
ugj/9NFlo7a1fzieD/Ny4GDjdih595BQNIMECkknAr+JtoSZ7uoL33TCXTUpX0yQjPzQxenp5FK9
GHH3WKFNiKZmEZObI0TaCzfZ13TUNAAhrJzjGbMoXnSRPM2tW21AWnbTCTdkHfSE4bN6bzDstdYP
UPMhlPday/IVS0nN4f37PIezMGkmBaEMzp/EBuTR4H7Jt/id2PoITr4qPndnHVlGsBizFNZ7EZd/
YY0yTVaMGh5VQrJXIppKVfn8dTlvHm2BvkMGPPOUUb4ot8gSZldcRKi09fHvtXWR0XGnWemKhOeY
bbedUuJh16yshy+X0++Z/QhnbomHF/dEbAtmqIVn7WG43nsGe0GNE0Ztm0MYUsRYDHjouqDoF6Ki
0SCcVOv8SkHO15XhHDGJZZUXt6zbmv83KZ8H1fucoQHSNvNmAW9GqX4WtiQvnwszA2uQQRpjvguf
G8HxlYSfEreqbXeI2IFhjJkyRsfAaET++fylYaBzyvQ3jcljg+9f42Z9oy08fAzsnjusmBV767Gd
+1FKzs9QRVucBvmeS1bbuZN15PK1S9wgMy5ab4qzsbNHNJZtU+s0jf1Rm0/bi1aWv1WLeGWp69++
bx2R/nc4a4Zd4fGO4lGI/Is0+y2NNeAjivo66Fesy1T5xSqRbPGBCBAurgcj599gUuYp14ClET/z
vC829evavz6lZ/IlfQdNZ2XY2u5onxtnRWEqnO3V+lox2L2uknrQcFCUJaiX4EAO5JG3w5pDRUxb
U9KGGf1tl3/Gm3HLHf8flx8fIB0/AyFuzMiCiOwBu3IE796QmuQn1BFceuAO33NDJnpx86zj5OEZ
O0VScudzHxLeesTby+y4PgHxIsaLlOe1nicZ99G0XNJiL8XtMpjK8fvZ+TYWOxm1FfZXZ/oCXrGo
eZ5hQ4cfKin/CFloYXdYGxixFkSqKgiVEoG8Q5SVsJeYKBLkc2uUZ1KI47s+QE+d8VIZKVtEAv1X
28Bw/6c3cAFXUKXRh6+r1AbBwQ19sxIsbPw3b53LReShI3kD4ZHpJPgvN2ZPjpbl03Y+UxP2QAd2
/UxFDX+agp5LPYzTWc4s7VxF4uKfMSSA03H5N0l/moIuyVLlarBsjrqL6mOTcXmKNKfaDuS5bPZ2
H1QCcLkv52W7eqa0MVBE95mRlKc1grjzz6G2OMfe+7WX7GjhOBj55Ua2Ct4LWTty+2JVR9pOvfhC
aTmvPl1jUlCDrXK/r/Hc0MoAVEqJvnT7LwrLl7gU3EG7QAY4cmVVoYV9Du+LKV56E+Q7NxjfbPNX
XrZFeg7VnNxV67S7PJvpTvF6FGOMDQcxnHb4v1+gdUTWCHr5E6SUZaru/P9RJizpZUkNgV6jp295
9NXMn86XZwpbz12+9mXs9P01i/yDIyozslsLVyAqbKtOTQCGdOymOa/79KC05qLqZGYYptt589J+
zyXB6PQHoAFqDFXAtMS6/NprQdSwv9mCl5vctDKtlYB0DG70U+9TPBqx7/CGKCJV8uMNvma5vh1N
MiYTgRLn42QFykJW2bZoxr8zrZ+1/fubPIQarQBx+LUtuQaAnNqpQyKpe0jDUbBskbeoswg1NFj2
cx9nPR71f1QGh7EQsttdRerEN7mtrKLpmUiREVsG5w7LcxLicvLH7cUJ0iPK4DC7PZuC142ScOJE
C2QNP4mRuIp1ytLDuNN2h6tA/f+X05sZlXMYVjmKczVS5JnaOLF1j677gMSoU+H4mVuY6r1r09oP
+wxyGWc6zffzUszLoHMX8PO+FNsf6Ahs/8y39xIImz5EH7hnGjB0TC223YMaKjTbwHBoAJzW0iuR
uvxXP1x9xhZpwEkWr4VRYAl1ZSoSC75lN7liGKUDOq1XZz2EjOPAhfXgdlKcaKwuJFgSPnupjgfq
Bi3t6HWGaVRGNESsspXcrYIYH/utDOrroQfdh6VzJePxmXaw824eQalZIyqqvVTWPvuduH3eRyWe
vGMEUvyzXwfHSwEUcU3bvqJVg2yqB2ItLzjtdSydRba3gV4so134jrHcLNpD8qgIq3UyDUMmLVt3
8WVH8pDOAowp52EdCxUYyrqo0Sii4st9RDQoezxpl/EwXE0m3ikOlY1zAuHnkuqeM5VPygVtV784
LmAhNi/zPFM9jkRyPMeT/bghB5C1I8LyXPQjAIL4UQeZ3C6XfPJ0CC4Jy+AzhNimToK3d8UVT3H+
rIuKyrE5G1P31wWBaRm7FzG+CAdsny7USAomqsdBBqnmhi32m0db7mJzLP1HQl362dH4UZY3wMcO
Gd7WKNgffXn61mH8M8fr3XavH9Al4El2GBnFlertbJMRAYDWeSS7yPt/Jm5WXhwz80EzyAuVxG+M
4YqBVXjIeZmTQHDsluy6FkxgzOMu86DQZ/M/hhMSEzKhg8JFWPDydwkXd76NZEJx3UvLi4X0DWLX
km0wdJxGJXoiWAht2FwP12yYiNgPs0EEfmt/Kz1IMnIDm8EoeI95X+1pN1pbYTy6YglpI7bcUMpU
rpqgk+BHbPuGEDQYuo0nTQu6CNoy9VyuoFbehe3LQ1GUbbSxXdQNQT3Uf/4ZuCvSBKO8BYNmEjnv
VzEcIsCuYkLxR08jv1KxifkttwDtIoXVEEW2yxdTK9UnBCN4esCsKHYzckUPfuOpjSRsNA8Nc2ce
G0Hz+0CF1gCxH8kQVqUhNZ5Q6B4m94F0tFP19Aa8cKSmfuDu7Pd+J6jznwuzlY7lvlva+0EKsv12
01EmZWB//vsjFAYFfeSPUwJKnAO7CBGLNAH6y3s8PBthiW6VGtTSr6MBUlTAULeB4Pk57CAxzd3n
LiGlIiaQon6gvTNjGyCtBkkw404FtZgpXAKSgV6Q+02pTYTFrn85JnOUycinq/KpKpe5e3qsV9Ra
gLFGUejp8pLWRhALvRqdTc/pQyVjFo03mZ0ZRJFYIb0Nf9cOkmueCAyz9eJjJgtC7Xiw6c3zs2Oa
VSxEz0CaRwDFxIB8SWwg+TnKr6ULbk7pi+ghP0W0WJ9oXk+wiZOEDQw422NptZSbI1WRbDstEjbF
LmSlY4X7V3Aax5z09s60a3fTxG2uqRHvpeGJhWcx9IFjz64tEXU2qFeyRyxbjEqAqLVMLJyQm04Z
AMxVgHHZFQNlg5hW5BwRtOX2LCDvCMshfjsH1MlsspC4jqtFq3o6sWlkuu5z4Dx7ffLPWfVmVf+G
skY64W+pxEmOvNWW83jU45/R0AKEzm6ifix7HN3WYEFXOQg6IIpfyVlnFigjRHpeVvGv7dERWajA
UgBcf9ZGQyyaGTPANLlJh9BUmxNIb+QPMfOPqU96lX9aunL8NA1GxfW1SWjG8tDhe+WahAaB/RuP
8AxQof6DHzL19ZKH/rUb0w8f8/x99NaskZSAEZ5qa3s3nQ5+yIQ/Qu1lFrZYOhP2ClDrzSguYYAu
qOqFBPp+Aeoc1Vn0Wa4THIhNrtmD2l9MEpuEax6nSnm6HCJtQ2t+mW1rNIULwo8anL0vPYDdK0aH
r1tjpFUrSrxQ08MrDBsBYRBeMetGYv+hEbjncenf1rv6ppKfN/q66JOKPvxHxyG2DCgZn/UMYRwJ
rYvqdDXeMHIUVqG2m71NTX9+GTWuM9IMTnRaJvgjSZPy6kaMiVqK8ujruYszui+wj21PRFgLRFfW
gCq2VHDJ10X2NUQJyOzavxwDbPaatFmimwNeYElD9rnzWBCNdg6u3n9vf4aSBYJRDrYDDM6V8fOQ
7ch7QMmbJQz2IUAqDlQTVKs/VNNxzQ5LAu15ErQeWTCh6m+QQgDFxoiF84alW7vtZOMA9qmSNL8l
jMsuWs4cD2/sfoqLsyJ1x7sA7eMqUHWzLWBnIav6yJ8rjkvOG/m+VVwtZb94hqO/8fLXrw4riX+m
Jcz83gEkE5Cz6LhDumqKOWuRsCY22ONxbIlZTCIalP2Tv2W2lrrzfAa+Y6KNYxcrdgajaaVvcbAa
N9tyRhsFC3Z85EHOvEZFSsvRGMXmCokzc4xX07gaXc7VLEN418eS9KULRX7OzGrQCZqq5TLSNVSL
ZZkki+nQ7/wgkQphvHz0gAUbxFU6/CCeTtPTCUwUH3dMwfRlN9696zm9Qcp1SbwGB5fjJj98oJ/Q
gF17BcPCE7cjKRtjErdi+hb1Fn+HwA+CwEBuJJbbSTJ9Ns1nKLNu6YHdSGpnpUn89VnBFP3vVWVi
dP4gJ5VApl3wk+5KUlwfIc1Wpkb8nksRZLzqoYesZn8jmLPzN7N/Pzp4w+Dmk7ACudsIwLkOO8ES
wOUt3RIFQID93fwLhebhtY7p2mjoqZYc9mpVp4uhZdUpvSsFBCZu6vVaJFzEwOQ9Aor2j2l3R+DN
icfNMGU+HgoZlzk1oLaM7p7UMT51nsZSnTql9uEeOqjIZqPz1+QUMYYC/6V+THSmuF3cClwlUb/p
0V0sOG74s2TDurQF2IgCjOxmw3SK1gedkN00441CYMhemtLctFCXiknclWQBmmBgYaSJblH02xLa
rzJgVxlRghnMVGwD43utNzHXp4Kuo/dI+Qwh9wXv02rnPuWJ2lBNwYpI9XKLwkDXnWMFFnUxj3ys
jtOBNHaVbAM9fvsmKldkPZdm2+cfrWg5u01+6erWsV7/h/fl3V3r4r9FaD6gssL66NHGGN0TXma5
pEJG/0T8sDP/1kUFzrWB1CBgg3ZEPKzTlk3PR7soAS/6fofRm58HCatrwCLZ9c6wOvHhdGB9gYLl
ZrCZdhNltk/CsU2NhL3OimIeTL3MZ767KEy+NKL5VyzzxOTg11uYXrnxMiKoRRyrnA2sXk1o97h1
t8XAyFicF6EaitxCy3e07vXfHHJLZ26iTyrhrVfg95LP0wfAzx4UHbSK/+HQr3aP5HOuZnU+5TBL
0o5ACy99GnnmfbMZvp00JN3v2x1AjgIYezQkb2PLSlm1JgiMoHaoEb1pj+kNszEQlCjIYMFqJ5yc
IhKqeOv0DVGyRbbv2BNgpMzxHQ1bHiDnZ5gAhPAIFZXuoOqUYO9k051d3XLJ8ox3/FC4dycsNahl
fTKEltsjo3JQUCvu23SitLbJbuDiiKUd5LGY8rNbMn5sMozJx6EvR/fD6mUG/RRG3xs+vttusEig
OZiWBi6k21gt5w3oXEqmI6xfdOMw6sYXnWaSmG+Gyu3WWZ8Y1BL8eF3+aGe9BI1T1SPzLjCpBHvB
BuTpWBnjXTvTEotIWi7oD1y3xCBQZ8jimNdSBQqDyq2XYu3oprrYN3yknNGuoQP7HCz5eX2koOvB
74dbUXtPJMc5IiR1olYHybxTtlB7d1AOyL9gl7BTWrqIZJZSTUUwSqP9NssfjKxo5JMkLGR+pbrO
2Sj+72sRdA5ZjoC4yFQTx9kWEeUj7mGJEY4uzpQ7rCg0U0Ypnc6i+yNUmyuvvEHR+JJXt1jqxYr7
EygGN2LgrrzrYWs0iFZlQRGy/fa1ExcTBJCNfqBNGnD5w6EOIdMFI9icZBKZBwzle6XX7nIu4AO5
KpPFE4WPnLQz6pba8aG65A14uDMVWbzOqExgEQtX4NiBC5tNdaFKRrDvp6pU2aMOm9MRUYBhXKC1
2q3GPBqNjudW/DecyHjYa/PIIaRgCwd6jbl075D7pzvtlzgraeMhh7vdBBvnjAPgPOqJ4p2iukSI
o6KOh/0S150XNLpu+7dtt7etLpkw6ipHTGOpziVy9j8HXSEQdEGaV3Hhar7w9JbcF0QHYrlAkT78
m5h3o7BREwCdk/jKGqV1hXuLTo6fkGpYEneCbsZGgYKOXlh7L1JG2n5ZoP+OlQ4yDO89e7tQqVmP
V2F6dgotHOZr4Q3aRz47IIh4Uu4pA0I9z5ZAX2kUWLnX9wJIzOGgHXZ6NkAi6vaLdZLQzT1GbgpH
HskcKvgDXeoyK5ksng/slCZ9UTfqsi1r97918f1V6M+g0ERwVyaHOviN6fQGp+UaI2rvBNQvY5jI
hJquZZWhkFhWvrxYSxykrjwK+cN8IDhfa/+N1zHLcoomV23X2OJKQcNt5/8mh4SfqEUgLYv5aQeG
LJKoFEaf51DtkU66C9nOVTyedGjFlyLtj3xR0Qpb/aOLjRWm7poSMDBy3nb0UHbKgj1eyPclIToU
pFnas5yxZqpHhZUKzF9k/Hj5fPbMhu/r2XxI31GUvMeTWxJJ6k8CtYEVm1/shzM5jVqSHddNlOQc
PdhhS0d/J33zNogkHqxhlwobbIBvN+CGe9Kks1gEYbRRuZ0N1PZ0uvB0ww5l2v+G92DmZFbH6kTp
pJkFZwlQwWD2Wm8HPf/5SmEQW8vQ5QQjmf54UWnCGfvle+ILn+VEDOhjxIQZIo7gw4hx55dH2C9e
BgZiPf8jaKefWsRsihbx4uZqpWDMiOSTetBWMhcEWs0y0rV6udoH+QmK7q5jSaBXpcjLGtoRJBL0
qyG9bHKT5wTqGcIp39VmadRxTOqWNrdE/lUFjQK2ifQqPKVwkAz5TwlcXn0v7OLlZtVhhRHT/YmO
LUJTfN5LiKvX1aMdJlvk8sZ8+1UYsHKwmBkfRhscpwveBQNTjsrlBQ2H5DNei/ufEaroJei9ODGm
QsiKOhDsFv3E3/eooqLDWYEzYiTYD5+qaDZzIH4pUZ/rbozItnnrBzi2rbdY6v3dhqKJSypXizaM
6NR9olsBu0g/ObYxWtqY2pDWVgjDNy2HZ6lpEpH8H1apUrYXLLadzrkPoRQguNYQn6rv7lFKThGh
cF3YhpBxxhRc1wCCXKVBOSoUvkaul1E54+fRifb2OAUqyHPQfmS4P81pOwgjqji2qSPmCEyVZPcS
oIJCgov7+Ar9QxQ6WuZnOI1BXb5Cj9xpPR02S4DM0onGXhdFGiK7f3znzs03Eqna2VW+sRJW20ON
p9xJSPt5T4W8q/BpRK++HPhQOKRB7xNGF9+Yyq+bSwxtu/qU1sIm7D7OqeMOl19QEp+DVhXjculZ
g/SyzqfJeYqVim97Wn/6E7SlPB7Yud3OTiEEr/lWfSzNbVO+Uc8zUdJA4k9AquSeZ/uASrIRsUJw
l4mXAQ7T3EOCsX49WknbGiy3XZyhuMlgK4RdvV/F8grCyS5zAw6ceVzcEfPORGBKtzYKKvBJYgwx
Ylgtel6Gy3ZjLr0hMP+x1k2jm4V2ejNuANpQdLtZs5HTml19f34v/XukHWpSSStl6KGGavomjLay
YJh+atehSUA9JMvC76BzfZ6GlJiXuaJkT+VSF3uK0fMq7Zniqujjll3UnMV496cPmNPBXkHX1hyv
xrVjqwL6hA5o4gKJTvNwCxgSXU2uoRh0PWNLfraLoWQvCQ04aRGDXNUTwtvn3c3xPXOJUTqmcEcX
eK9j68piFKTPaBjd2IVoQDFcKyaAnQaeEtFeoYn4KVbVmrvO6CS2aiQ8G+FHKtOLXW3mj86YYS5r
JLsNXYKr4IuzXECcK5VjT3DRbmqRlBs4jWTG0WOa4fJTveUm7DuTh9TIho3qmLyIW/gb0vsJE0Uz
WSJcSBIbsNgK+tEoHAr6PG2cm7pqNfUa/fRp5b4UgsbHcpmuTLMOHLTYoCQxL1eIq3KCmSEkaSoR
TBO5cnkOCSSgPxhDBbVNZRTbVzBLYSOvtvt9lIjy5kMTQsF2ZnzcnJhC71TAiTa4FZP7gQcYv7/X
kV4MMfQOjUONiFQmOaGxudiwQdEJYCU3/EGuEKJXYRtHJxgS3ghOffdxcdh6GVAKsR5WvFiSqRUi
R8IpYzmO+JvrpyVPHAiFNVfeXjGnzSy3wp003UxmO5+FTzMu27PZtPTKFIPX8rDRdZvTx9n/1ZrS
94PVN+ZXKOb1FnDBOw3nf5Atu3tN97FuqWqxItkgZXYwMxSFd8S5PQFuV0chKOOmHnqt19IYTDFr
1kJeEOxll7L6MVGsLTuCp0ubi3EHaOEv8Poet0O2XyK982jnkJRkYuUhBeHJTqUlpbAlfNrI9DFi
5npQqXK8rhfH+sKkEz8XQbuupSofjkmRUMHL84pbgk/DQ5bSaLSJgajX96pxwVRIE2xQB1CDJAp3
4CTK+a2uSZ72zj2Qu/MhTkGdfNDjBNDh/2jND1bC0qdeui0z+Cj5Kivwrc17+rilv4HFB7dPprZB
2sURGbHEjwVCCvqhivVSHM2SoYhgTI2i2YvpxSCSqsPUd2aRE82SXnjtiXxU+G/5UeMo+S0cEBER
5H1hXLMgGoGnYLVpL+qPAaN3xwsQgy9f3oI19MUNSSqns94y30+WBusGQauJzfh0MFEpdpenJyRR
sQTJg0RsQx57i9I=
`protect end_protected
