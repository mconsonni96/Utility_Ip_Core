`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
etZresF5hBSNznBZk9HMfuBmVQ9yKsi6DBgZJhdJduf0Oevo3yFTDixGAM1jW1H2MaMoFROMTB15
cizckj74Fs+OFsKBNM7+/0n4AHXUj6EuVb0JZIUFOoJEvPaZ2ULbu6AKMLM2Ekq9PJxwhwecpnfT
vBgOlkUdPgd7GxrbquXNr53/V8SbmVN3Be17gc+vYTUaq1902W7a3lBbmDXW4Y1fsVsiuI1siBh8
2PsHCmDk3Sxuxj5lOYTx9YbUt/zKl0sQ1I1bOAObMkE5tpErcceByapRJVFmp2LdGLrpO2fIKY+y
65J8LxSnYPmPKXMie8W5CliKNvq/nbg7OH1ZCQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="2RTF3c/BV+u5lTZnfr2fWu9ViX6nCx1tCkzvskiOztI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 139808)
`protect data_block
/i87smxY461DiFDtsOvqxT8UJxFe4n8BMlK41QsgdH2jRCWUr12AZ2gGNYY31uZ5f5d5bxNKLWfc
1MjIt7B4NmP+KOrUsiZ8fhDD+xAGcv6SqAlG74Rfh10PQc3UufuY3x7nLHdaC3boePkH8a/tcCTs
gOmy2WnXLcvm7iSA4QX2vQVynq6dlg1H2P2lHmZT7iA55yQIeQAje54MbFrbJmZAhVpsgU8UWDyA
q/p1STV2h6VDm27MdzSm13nB2jP9rV+NhcMm5CJ2y+V6Q5Z1f6LQfXIs4F6fnImfz+sJsPJk4VRX
yjDvbAOw7unabD6FoMA3T4nO3eLQF1WTLVvaakUXcNho5Yr2Z3ioCypYS+a8JqEj31C72xrf3SaY
xuat07iqrV+/gGpOEp1DIeEXbNl6FveG8nye1P2/Re0MR8d0K8x3b11gTM7+RU5wQhcm9uYk+ZCb
jg9dCteVPdXJYM9v80P/AG3h4HLveBvIZJNftgbq21FhB82R3rW0vU1/80x5LvfGL0RKYwKNIalr
jx/N1QfIMVpu87UZvvqyMgMgtPSnH/UHdw6nIpjBl1/95H27DvceMur4G9XHsRbuN3Gp6Bo7d9hL
pFnSF+wkb13+0OTLWWT+09kgQ/jMXwXzc/yn+SWYi4yaQb+bAFZrGmjuGs4iQanbBADIkSwi2QOM
pURXHumQZfhiQo2Oo//ZXSk5uHSyodTljqfExltZvjFoLqilK3NED4J2DSmDjSd4t2J/TVFR5CTC
IIKWRJ9jUDEjnaCVX6W5zB8dWCXT3ezCBAExh6691iVM9D4U6n/TN5g0oUBwp+wACd+ihmp0vbKW
ABdMlA9fhF0YK+mFFJDpg5JhuSntDRr0cCyF5ftpRvDrgdS4De95a8ImxjxlXFh89o90aWDD8vdp
32HFu/eOtBB1C3KP487XYjyM5m55jFeJImwZXdaZGZcwBl29j+tY9+czrk+ikU7uE3Pge0IwN10i
RSajqK+0nMULQQm9uE8MU3z/fUTuPmMM58XcGMG0Cl7W9bE4Fr/ojRj44as7+zPaHemh5GwBQ4Js
Kjyoc1AiKc0V8q78GeVMeCGKYYQUhr8YOOC96DrW0PJJOZoMhAMwnYj2y64L31Nths1EShmTSlsV
XyvzwVwgqXc9Z88k5jhsoqX+9BGt4B1yFJ22hDxxKI306T204EcJnwQLNWcYf3o8BlrkaW1lN2fa
ptz704ldY6nce6opuwJ/5RLuVb9RhTTF4ZilFcUd5Ghjl1G3rm7f5sWp8ls/OC0EMit9Mj+/2q6m
4wKKGZhC3eAQhZCoZijM3dTSWpw27Am5bDHKe2erXhvxYb47S3sNtHJIXxWW1VfLymh0sxYb6ez4
aQEuFx77r43csJfF7w8KkMfX4zsTb0Py0HdHAhzlk9iLOMFRyQLNdnw65DkGFLIIE5SIVoBWnulC
kDDdKg8xI9jSD60tFBcxk5z1pUDHbHZgXIqoeQAfvNlaeKkTPqb+7LcX0DC9BqciyE35z6XasWV6
F9M7V4JaRlYoNk5sKSdlfLwzhV4pp4wFZc2WcGzjv9MwSOtZg3wiKbgL12b6ekDX7br/shSn6h/p
7f8puVqrEmegHI9QbWmfVVxGJ8o98cIpI6hois9NOpePWlq8wIp8mzsnwVW8c6a5Xpy1gOpGOZXa
D0X3ETAp0atTEA4iQNHzesz8ihXrFO5BQY7HO7UjLUut5A0m0QxerWvNsreuKnD30b1IO2mRh8+t
z3xeY29h3e767fDLKa7ZOSKK2nyU7Y56G5Av8guMVqGTBCT+UK0FFqNYSysJ83IQNwJpFYNIuU8U
dup8Yxqi08r2/LcsnFY2yknoMgpdSGTdEZZIIFfjtDADFbGdGnAMWHnZOvCKXDZa+2NQL7Ud0Rtq
21yjjg/X3WbMRBuazr/WpnaANxAsbOXFBAhpNA7cHK7JLdVIJmqHVvvRKwQtRvxP031WMNhu88d+
CfIY3ibhFJEFyaXKjzbHTGLsL++fbPfSc7fy7pj4IjNNz7tIijwwtKAnjcsL8cwbSCtGHJiEM1xB
Pnh6BG+va0fpwLXMDWkhTsuYimQe1WDu+8iuj7vhLjbQu9I9wluoJ+vy4J8ZKJ2cvX39vqmeJpsk
wNea3KwT7s5CvYjkjK2v1xEc4+Zm/24/O91N3Dq1J6ueAsC5xgFb2FCJBwDLaiDEsQsTZq2sV9kg
onlmRFIIKUhsXS4eZjvRUWk1mIO2AkoVTJb/7RMlEgWEeMdTlF4Em1NKTlHvsh5bSsXajASo9wJE
/tLhk8L2rH6OLiuYlzR11FiLDytzj6GnM6uGg4swapEflQPyPsgn9E90XWw9o6m90f5Fd9Q8Te6J
Tlt2ErRwo+YgH8x3t7QlH7pQjCo4kIEoHtQq1Gz415ykzPc+Qlqsx21Wrqi/rmrbaGmXgMihbpP/
hPWM19NCi6HUj8gZprbSezgOldc4xBiIV22i8X0eBq+t+0RyjJDXicv5j2sxlPaHmYgLoub+wTLK
oxZWi2tJVnyJcAXnumZiu4UVWZmttG+fXLTBFf/ctg3DpNeX0EleIluDD8iduQpYNyWEB9PThFvX
Tb5r4ZGFUaARo1mfc4u656gL3GhZErXL4bRhM5/V/fo1Ol56j1uEZga75hzDSQ1/bNCVox1AdH8v
ShLPSzkNqwM3KShQ4xPtlRXNH2ctl15B7cTRPLTiLZyNB26qWMbGp0FkH+NgtTjPaIu8AYhOlzsX
g6FlidVm9mLiECiNpcn7C/ytwZuBCHQNr0fjyRGKS7u7wEZkPLQVwZ0swraNKJlCTpARp/R+E/4H
+BaAWUV3X0n/IVcYR26vLF6xdTBJjLxOYUNt7oTLzTpZiP3coqyjH18jhNwzRUYbF0I+oyLE5pZH
Wh95yfsUnCe2Dzvj87ytw8xePXpYL1hNMl//9bViilMSOkwI+Ui1VP1zDX/4XI8q0bqRzPp9wfCb
hjFoh8sI/Sj0vPwVnKl82hekzDuip0zobGvF/hmg+G14ry8zeNTXRFKiCiXMqOv9YgMnUkUCfjlS
adV/asKKbXRbcyV9X4z4YcWib2A9iWtRuSdZrX0doDZX5po1UwzUF275u7i/x9AfP2wjETujiMxd
MOq3CID+5URnDYO5mI5m0+X1FKrrXOefB/2n1xfOGpbKKHYUSkCTW37ZlRx2BgwzmZ5kdy6dG7rd
WtpeclhKpMJC1eDq2e9F60ADDV42O4FCfdUCP9UX1iqCyDwua2dK4oDiYJ2hGmn3RJYxpEOwLiAn
CtzJZdI9IEQCGd0hliZo+65BgblSMDwPmeDl7NvTx9B23OzT/j3MMJSd+tSdsfQLc64u4plRJWEE
bW/bxuJVY7y71dbW2LASkH6iMOr8nXmWmxVZikXc5GjTI5auycVl7ssCxRyak0/5x8oI09EBLeFX
Zae1m8WT9GCNoTXOXURWnsj1mPyP1r/EKhfTXDRWS9r+BZG4/SWf7zweymUPiT6DwyiPGWUDv75F
IVcYoGhfKC3VrHONvLVXedVCkP7soOKZnF6Pg7/vFiU/Yyn+H75oRt1sB2U3mLtHE2JUsD0kdqMY
Bu3u/9tYX9MNqHdqLX8QBf7hJCWi40bqesI6SgUgQt3Vn66974zPmOLoWMNh+Rqt4QpFBMxGIOOY
3DeE3d/tBo3iFf10cI2wQJQMayEXOA2C39/64rV746Sys3//w0IxI1BSwie+bX2Jxazrrtz2jCCW
Wlvm5KChSpShhZ4FOjKv0obn/0CSQzsRdyG/doKRBQgqmFMQ19H7ahL7dK/72nNwW0dyUUjC5+ZK
off9fEo+EeVgKvnczEwoQOANoZv+80ikb9WACc0t+iQ2yp7q78hpTROd250LJMuwTkiaROtSde0X
EmubmTw8M7l9dwEkyjnq/jmETUTyHc6KnagPBD9UKO07Lec5bFx3pKYwmS4UDKUpXBjQ6QEIv8gq
TU/ZzVniRyd+IaLPtJpAJCIEtkYIBkYAQawnxIzQPIv39+01EX68SRJvSxI3p/gIOsx//zzje6sq
Qoy7IqrJAtGxqGAfkvnv7817au1bSC03VoPPPO+8GHaoCgf9slPrMqohm2nW019tpzVGWarWHBg2
yrG7xNcovZyUdUNF+tL6XFrLNE8qzekGbFiTM4O4lD29tjP8ALA0WYeuQvtSrTszR8JJf1ov5NER
rojB6lUtcM5tapTBDXXYBBCQyL1Iy7xl73oQcZrbfJrYlu2qNS3j3IDqWlEBTId0P1APdLEJABdS
3T+6fu1sT8Y1vvb+0ukiuGOxRs8ZNYAMRGqkeLLw1S5BUMcXV0OYDXJbmjTma6zVqhi9i08qiFLx
kBnXDYqIncPoERMkjFD5qer9OBMceovFSLx89y0OZGM611vfYZ9vV2m0YKc1XCfVjHz+8q7gz+gI
B5plusYy0bDhP7vKJXAGGEtoUskls884jimpOFgM9FYZdX5FzR6oc+hxB6RDdpgvmAi3i0dyiCeP
NtA6VgfzvhXUG7FSfTVy0vlhYm5/mNSg+5pPlGsyaVI8+GTQzij+vnoKZJVKJy7UOHogsed241vz
ArO9vjATHQbevWUUp0Hmi8kNkE+OIKbR7OgkfB9zgzlfS3OvMBugU3kbcM3Dxu1AUxN64CkkN6tA
2qgqqLtxWcEfMSMQiLN559aB9OH32uBM1ujHulBXGOjmf09r4u3yMF5ffWMEq+HCrA7wFQsziZFi
Y4rljrEHIJ18gUv8lCQIMTB+KFoYL+4eW48hM/+y1QVRvKVoBCpDuGp6LTXVPAKFW5olgrylrRXF
byASGN7/o4P6WD654FmTWDgO9ibyLtPUeqRvmHK15zkKZq5bjAMcP89y63nqmumNGsHvLYIQvyol
WtB1WjNeYj5NouPTDZjc13bEiLVwiZAMWzjv859SSzXxZLP8pHG3NhJsjBQZ15M5mqOpix1KBd47
7sZAm3ZREqkEeGxecvft8BchEQagIKPdkXNu7tqh53+mnIlkxdSocPUEKrXNQNWq5lypUgn+xhyk
ImkWAXwjPTUOg0uggQRcVmJxFV+IsQZMdBORNMfcg830gAz2FrkTCCqQPNgL7+L3hTaP8YNQ0bvF
aJaIA+c43v9IIlcjJgSeIWkMYz2kmlM1BEsDFVRxLleYLmQd5TB0L91VZGlpT2mPrM5Jq43Bf+o/
3FUaojOwHYUk/55OFCAt2TX9+GAhgnoVLz4LgHep6Ubion0JhWPBTiUJwFq9J1F3msoWv2Ar9xma
L+coZAc40FnhR6wKHlgAHT4sxAJBZWtQXB2xwLW6v4yuEx5ghh7a11YnUUvKyFJuRk4EjgIfh+yF
q1bs8eOGhhAyqLd2lbRw0GLnd0jfeBDyCu/66jMlmQVMwr1+U1EYjMVERx/NQQIG6xMEu4nIxvSh
JhRaxWEMLeyRy2hpgGZG1LbWcOqRU/6K29T9E3Ncg56akzVgVSHx9WdE4Xq3+m1ovYi3OeAFOe3T
7jqvvqseh4XgYUyABxk2kHn7kAmuE9FFeX0vUHu3Y7TzXEY35AI2Ey+hcPAhAkbcbX87Y6LbzuGK
W9LfXVMRtZGzy5HcQkUJKwEKPqNqZcCYCqVL/wEG0gg1Z2pFLDpf5ocq5irbs8KBa40fDRVQo7j3
c4K1BywsEr6pK1En9STu+Hb2jl+Jq9+OzRqBnzfZoWOpJK0HxPx/gIEttoDwFZio/nqfYRwmGcId
A3dL2gRYnCjhYO7W7JPdiKzlVxunquGxT2hjYNWAT6rrindT+1H5wCdZ4LO6WuYEJzB1+CHoKour
FjNilcE4ITKi2U5D2mWLXi6T6GxxdX7Sqt1D0Ukt/4jcDIBjJU8W2agSSt9gwoqhvhYyGVMYHd7n
TTGamjSPPDbU9MHhRluguCa5WbxzB3jhYnb6JEeInDC8xIdFED9ZPKLfEklbzkPY8IZPlUQEc93/
IemKilxScUxHhrXCbjPaB7rWdGsrM6xFJOFKpMPX7J8SCb9COg7CgXxezpzrM0x1+kcKabWfmc19
iZ/m13h2SON1JZ9gCDMKYcVXegryVbnmMPAvQqi+f7FTDxjEmiuO4+3aDdsjCY9Q0zBBkGM7DVpc
RVYfQNHbR2lHt8VMIpOQcqNy7iqTV4gaJazNlmDebUAdvpz4/9LHUoEUs32+Tf6vw4PkycsqaO14
iqriWJawdQEVaoG0Oiaw6c1Fpt2U1uZk9zhNtJ1UqO7LOyiE44FqTIOWUhU+HnE0LjXvs0zowxFR
Ig3yA1nxQT5WbWWM8CssW7eUzkWP04gU7uEyxEQ8BzUAISc/n05dpSaWDHWXfHubdIhDtHIdNxuh
Yjj8P5/fcIkhDMngePYCA5WgucvhmMvro0i7/sFSWJXhCwNuDdRSwNycCtXy8fdkZuLbRJyBLIRD
jR3eSSIavbBO1WLW8IFPjIbyMrYQny4VVgPCoT4cekrRl/OFaDI+U7HqB3T9Ey2admVMi7/agSjN
lRrUY/OLFc+1VzpHNqsghU7a/wKV4DHn0Ueg9it+rmN5MHhGtetfei0zUaWzBYsNf2dFSIv6Bcig
z+x2VrW3cl7VZwhSaQctqo6u/sIayQ3k71rv+ZOq7r9JzZY7LecnkYQ2/go7DoV+1FjQBPNQ/ot/
f/gHlO4/2i4aat0P4Zv4RUpd5AZAqU/MucP3fbW3IOD4P7ImXsl1QliThUU0YMHvJkp2j1SXxiIZ
W45EvpMo+lY2mBVrStthg2AiaHjQvdTSdzAa4be5JezXPbZcA4VSkICXCpF809vSlP1uheXgzN2I
Bd8B4kFs4fWNFvtdmSboxYuwb0V6ZFYu2QqqlAntC61FeTa3YgAqTXdQzZMMt3dof2I0R1r0nPuG
6hujjFa19mqICHGL+ZWjEaHirEMwvopAGz/0YMbME76r0BBOzoKpXSyZtCMcKsmS2P3cj0fr+kc7
nt+6uT8YVKrByJDzFD3Z9fBJkGcO03XFXAO6G/hNQhjkwQE9/khNNkn3kAj5PgbozV7VjSct1oYC
ObXwWtRLWFGPOk4ri3O6b6AHiqNA+nJDZLVynf+whvofC46w162NfYxPJ399Jt/CrKHNF4LkK6pI
OIo8WR6aKW9DF16hC+OuPu++9wfw2J7V4l6j3vY3JVhemLzCTfWHUOKZugD7fGo2HCBU51/zh9Ps
04dGc9Hvi6gHEtK0tvRTb3d2bIBBQaQvE+VhoCxywCJzdos27r2u5VArpVXfd7YS2VZq0k7lFJ2Q
cE1KkdMKBl6NMZoerZrthcZ9aWzyLxuTOL+x8fclEyN8WEwVY62ywfyL9FjxbCJeIGPyamZIhaP/
KLUrqlZl6Eb221NiCUZ79cToDc6F489TA15vmbIR3T1pNoM2Roatm0IyI2SEZ6bxohsMWx9fSYs5
5ThGVZVXoxAEQ+0vXbJd+iEe5S7cCS0mIgE4jur0yXuWr+LHhT1htVo5cABcAYZLDvW7LXrR24JI
bDA7kq03Xc/ZCsLavvwsuxK4Fk9ZxtDa/VATr4KBenGmEqs5beHGVOTt6IxlI9P5JrLMPd1zBzaj
8Y/egD/d8ytsYLyVFMz5GH+o81NI/O3JLdMV/17CVmnbxgsYByuFWYaQfHPGCljE90VuJeRz2IOy
O3WSBBAtDpxA76JgGjZt71TSS/JsDOGZvzhK4R6ni8I7Na8CA8+uCP2BUDJmBK/BnaeG51VtHqr4
PBwABTsIFIJoaqOSId6mUewhCBcaHr1mnc+Tb8mEgFWXteOj7kIlA1sYExvltsMJ1j2VVdwAE5aG
iZVU0a4eCY+pNvJGNH2a4YKE8tw4LZYyz52MR5725gT7Mka8q6oxXMTIRP/J8TClvlif2GOf7oKY
Q0GTI+FZ97GbCHwJ9+aOMRMWkBvZZtOgLgjIBl6N+0k8c5nmAczAMaiI0vvj6NyD2sI4cj5vUIyD
zftEmVeIlTW33kVPVrr4v2FrTZhymqtfJGyFaduP0z7KP9Nbv/hnmhwqnhblmI4UakcZuKGFg/MV
qP93t9+Ld7QsR/7ZanrmEqDk+7tmhgH+HzcBXYBbb/BjLx23FP+8BCg0qcthnyDhIeYMGTYyADDP
YHN/+Td2ydb/kggJZiyEtHEiXwvujp7cm38b3FNIhb+hRMNv7FWTpemRBvd3OgtDz+N8tHruEzxr
mhKFPZPx1ExtIR2H9PqGMngJk0pu0OAba0zX5NxXWR82aafeMBltohgzWJyeupqhKEeI6PyTpKDx
ThxvMPnQsjt5q+Oc8ys4+zdWBjz9hVX6FcypQ2Zm22eZNRzfhcG6NVGAYPbo7TNLBdFk09xhdx+4
RM3gvppEwsN7j1puoW/vY02SzaKk+2e8NlC1DyG9NpKEuD9UmiYZz+9fjutAQrOjCbftKryiRs/6
CuTKq7h+dixMaG0vw6i125bkP/05ufGIxj97BKy1N7jqg1OQwamOZRdB5ZVRqGcgeBJM60beHZfG
6VdSFibkyx3sqkrpNMCZytBq59ty3mKb0ekkjvzW01Z/btPtX/2rqGzpFTXjUbDkfAzGTS8SbbTJ
GTDCXmbdfLSB0wcvzWWt6MCsQr65YTq5dPCDxV1FqvMNLgFD1lKjC9egs1rWXMTCTyhLcRu7eT1l
SdrHK9OXu/HAjE6GzjN5X+ZiqzrpuBWsFJKDcdjB4S1evSV5XHrA0yEVbDbETrj8t6Wt7mWL3CNa
e7HkyVIhkxn8OrKJ3ZghpqGqKRPqH8kjHZ7T5lWo2XycWTu0e+K1kcEHYJduuMDSVnJMmT+hVoX+
FE5dMLLIfwrkFhoto/RfROcn3WEkzP6d5Sy1fGVBi1v7GIj4EF8OeSbkYWziq++cB4FOL+FJ7FW2
8pZZ8m2EzAVGSC0FS/XH85+S4pyv94CvpN4l4JEQAAqcGzKiLUPug2kucI5H2spl8Yjo/aoO+LnR
pVomn0GWw49V6jwGXnCcpNOIMysUzB58RyBgDhzfqZFVUsniM/kJVg5XPu7jXJ5aseq400O1xlRW
9NdZjQcCX1SK+uxJZkKtwWN8u8Tn7SASfJfS51zOadeRxLyAe2kFOr0uiPdGh3Tby+7PvBAl5eqj
TZCT8+p90pm9pQgUBGMRGPJkxU0gHWOKRqpPcuEcqb5M7+W3ZIysYioyRKDEFzE4TBPfDyvcVL8s
Hc0tDJKoa7pR7JurqeF1m+ue2vhYW28bJLXG6FOKoyN8ecXzTU2YlI/93jvcPSkV8QjHiOgLTJDA
4eGBcNgwJMXBwae70g6+cAlPgwbPaB+/lipOBy4+zDpizf9pCkyFjiaw8XLNcPNo5NSah5apMf/q
DVN4mtsWjbYej7VcWYdTaRvrMhIVKvRRuXJqZ6RBP47v/0sIVBAZDZbebLNQ/BlArIOiJF6jJ+1N
VWxv2fRDlJPA2sm/B3YN87uue9AxBZE9XljGwXBR/ryMJAVm8BabWCCSJZR3eyvHQiNApvaLbew4
l0JTFR/ISF9CTu4rQiZefmVl3sOdFy8CzZGBTEwji7xMbgt0Fhfv5Zp+/llg5vCucgL+WNMraebQ
aLALnG4JCj/24XPtDM57DXeywyUyjdL95M6yjV732JMKXGVFZ9EbcWEjq9NpfpTCzUasACEohgXh
9iETp1fUzdqrLkl9f2t/oBLrZIyrQurLJ6EMtu9KG0itzbuCYb3vlMtDCq/vLuekJjq+GEoLCidn
Q+0IiPAipP6vqPuGkpPN+J/yAzuZHIzjt/bEa6qNyP9d8279DWB21e2umG2KJ35GzmTO/2l5u0UH
nhRHf+Igfzpz9hffarOqrO727ue1Vey5LFOWZKL1wCzeLXVDiA0Tl+JgRMGT61qRkXAvE/7AAhwc
prXnnomyXv8UGMn2logKCX5AiScwwQZaHhWHQTFpJA/0Mw8yRAItDtfuwUKUE7HsbyQXGQgCTHMf
irJ8cqjTqPcRc9NhPEpi7PU13yTIbZ8lR/mzigJ69JaDg4BOwxGmp3fPRjIbSqdqVheL277yHJRH
V5/RVmerF+nzWluMWpmU1DqzANcs9ZNONWwOUlcxRaVhlyk5VQXmLjzRWncUe/x4+uEUMtiRXNk2
k/1wA28OTHjC2Qz1W6wVKoFhQF7eqlCElSWVIR+uUtNHslaNA8i0dMdLizfv63GRX5KpjTN96IR1
BcC+SE5HNp+4Z7szR7cVSwmUTlQ8nHvyvOikF2HCKxbcFjo/2owbTVk66yIqz5An5HeIbF0/rFP3
mcJEn7nJ/8NkIJcDzp8QFTGY8tSBUor2SS4I+70wTJHm3HWWL9Wd8mELTU3n1or8vt3JgN5OSrId
rv9ErMVbib/UQiMHZsANBGQh+EFHccPN8vZo+hpW5xwYhB6JhCEbP1BOHYBo3/0QJD+kMcq3as0c
syFZ8ac885SIt79+SFC2hteOvkAWYC1xmNHLFC25fbS+Cdz2qGxKkzS3+kXx/xhwWFlru9pE2H1c
jZk2G+1qzZrFzsvqt34aGfNxRNyzJ9jVtcSaFhJpF94l2abIQzSS/Qu+fY/OGIKrFihz2hdozUax
K3asZDZtyvyswZiPvMNUEZBfgF9Zk7UIKGnUGwVo+TBN6kkZ6OXS3PVh9KiWHk8lzKtUmjwO9CRr
wLrgZawji6YJD6Oy04EAyTl7K0gmmpCIx0oHveGXimejirIDSWl2dJYy80H8INvk/Kz29xbx1GqX
1PWNOj3TPL565znfTBc1SiNpJzUUlGZiMDFUqyLalQmqQsWKtBrKn1cGH2BISxn3D2L1KgrjC9Cc
7sPcDMS5cepY7Hexk9zQmwWTNpIXdempFoLn3mT72CTRa5uVdEeruM5aTOo0HVZV0pRCEvV+4T3V
HhIHzVYA3mrZwh0qO521cg0VGYpPxv/Y3KuMTsRDk3Qw4CcKudehO1jrn6kmgFa6bANW8psXtURo
/5EqXBpjd+ndyjv30YxkQbnLC2CpcPRY243YK0xSnCJLQwHCSRNjZLyU67yPhFqFpxVCXJMPI+O2
k5S9eOOU0Fvwydv2DcZLpkTsh1h0xttu9Dbo3r0INYGFw31T/C3SsZNWj3t4NLHGDawC/83B/l1H
GncbLWRNNe1totI7xs/DP3C1TozbjbYIwbyduQ6YBf9ViGqC28MSZKNzz/oE28lEUt0zeiygN6js
TAlLQEeyCbVkeUVowJ31IK92J9gc4jCFuqnJkKRr6Gjl4gblMhsmqJl1TXpTP7RYnpFO2SRZhOmS
fes/oE7oz0Hx2qW9398HgaSRx/CugYW5RlgcHifp+Z0885eIa3hXyMYlANaX/spz54Zh1oqj0w50
PngiQz/iJ5mubBPbPBEYGma2oEYyvqZ8pW/wBxm4bkSrly+QuetQExmL7yzdoJ9QloYz2AtkunKf
4pLWvHf8wAGg/IrvJ9CoeXm46il91J3Ehrz4NaA0q+4zCTy3BTcwZ9pRpT1iTq9MyxR7oL2C8iC0
kykniwoVRUWqXPSghjFedZRuUKNeNo5Vq369GZWKsX1AbWRRSlRrbCZEm8pHhOysZSAMfg1q1wFH
4YIKM+JmTWEhJOHcRh0oNRqxGayIgRxhlHy4eAmsC7VndwKsQX2LJ3IJx7jnE7KhjtLM834PT3di
fQjLQoRPhC6zxUpJBe6/vNQZflw/302EPQ2cYq8rXxwG/HNayLsoD2QMVK0KEg6c320VFIEoBe4o
6dkSwB3hZkLJ7D2+/6kc0t6R7cBvAE1SDbXfLY/5ZgiO7RoQFVw0cml42c0cIbfodDONENyqRxGy
6wEUXS3i6wXvzkU1PIfogpo+Y0ZCLivva0Pq1ogK12QWJIs0782xKTdkZtRCGKhGHXz/dlkhlL0V
nBRkU5wMZTGQdMAvMiEn5dvH0S9xmPlwWJinCQfpV/Cp2lAPSQmjt0fNOIMZTW8dSRQzkADbFTZb
NuOeAWFtfUXpnidq7amJBXVNb5gVh8t/CqC8hOEw4Ybp9BlDggVdmdttx3gewNRlAT3WYigMISJ5
YEVoAi+N2Qize+wFEWYKKdJVOlZu46/Nr1xTL4yXDdczzsUJSYqA0GI3HyRKbynoHyR+spk6AVf4
ryyoGlAWjLFDaX13NpZ8SW3n5KwYBi5lv4siXevjvOdMaHLeRMNJ+gxpeawFBBOEQqyD/ihs6TBy
t8Bvt14eI57lEEGsq7CFk44L/FXHLBuh9gZ4Ma8Adc6PU9ZKwer1SKOmp4QpJB60S4f8r2ENyRW5
2cPagm/nRUZbMCx/66ZZj3p/o7G20zew9EOKXiZ4ejWCEgF9gwE8KJ7E3ScyO0iVYShwQ5uzgO1s
/gZF1I2d6YHaUaMmYstZ82OYI3b/c9adHgb0Wcj8O6QHKu1tuG5+nnHep00mTwlodh3GxZN/of5/
8hJ9+b8L1KIvnU+rjaFdWahmLydl03VpMy00vSGLzwLV7rIuf1qHUpbcnVfCqKYlqu79MWlsMl7B
6v/GXwPDiSJT2ZQHMzR/0SvjBB5WQ7XX3afNJYV0r+TmZBAa7IBhWptwccW2ifNgbXTizmvS8mS+
0yRAxXW1bsrimil6FzTSOZWevObToHAqsZjoAEBATmvz3Dnjvu5YOquQVe8WvVZaGL6h2XwoE2le
qxi1sz9BwCAJ+McAQXN/Ah9/iKzGmGN5U65e40qyLgzX3nsnlXgnOpYEQeq7Q94Ioq246Wtr6SLK
udaTClPQ7ZDrt5rEbcbgR6aDk4alYtM4ypR0bczKhdBamLAtKnieI6SdZDzh+vJKr9CpDAeKzeWO
4EnvL5TfQbQhRSAIvd34NP3USrSKuLNMK5DdzW/BlmrVwNFmYE+gg1zSTmBLWihQObgEf4RFJCHN
qFiTpbmLKyxbIUFeGq8mvQiNeWoQ9D5lRO4u21QRUvrwdY6D0K46EVz8McOZEBVGqir49+trMQb7
XA/46n5HB0TXGqHy9rw7a/M6Cn035a2uQojjua5Ltdm9Lx6WWCzfHRtEnNhx3CRYgWFlc5pWKVEF
H23N2+TtrRN5amgBwoC2gDBouCAc8NcCDNM618uJayXxaUjOkwIyzwDNC6WtZZNUnWtCfHH5VAgC
3i9tpeDOjtTGRWeNtQoQJ98YYThvEiQlVPJPeQNJSGAO+leKRMOAC6S6djyH8N4NkJCC/5r2IESq
3e8DsSp64oqf+uvIiHTcOOSCwR0AkUjBGtIq35p+tfj1gSmhfqZxqfyqHzp2UZRc6A/wHuv6okeH
4sESoUCYKzFjD5+O7JJsKlVP3ii5hMvZbyTj3b8tEkJ6ERoqCTtRQAmgbgMTrnZs3LVHjy+kIPwp
sNPPgC66Ulhk6EReyazbXuoBgufywHS/7MIflYCujdLExb5+VtdoEQo4j7VC6q2bq7+KnxARazfq
zzqzEbIKkNB7h1bX7yCfc/7QbrXV/dkkR1JK+3YY95qxEzMXHFBbavBqmwGd0ZTBitIb1Ek/o9VT
UmCI0NbXMVim1nJD/m/vcLk3aB0WaRul/OT6387xEVyvGMi61tEuauTd9GgeGwfZrig2b83f6ujb
8wcVUpw1MV9xlWubhglvez171+q3Iv1gJiMrjWZaiyjXD0DA9NgiQgrZEiGR3n9H3tH41Pzl9h+a
G1NdBEHcqVGCNlh8jkKjJzpNh8u784+d2tPgGSiKirQQ0eYBYGaR+9mD/MaeTjocLdtr92KHYz29
PgP3bffxWOWy4btEV5jT6EHA2TAqHSX2LiOaimCda7iFUGBXUiH0In/XWipvdZE5h2argRBOmXXg
Zypx3ehDH6FgY8WhIkTs11wmP2myVvVAwVdYqZty3jrw+H4ipvHnOsvzwnvf9lTuePhIhTDXKLpu
3QjKswtpQ0eVzMM1aO9Etd4K0GX0yDVD98kYLmf1/U4jn9VQFVQIGsvbHxmwf47tpinfNiYdkOsi
RhVM5N8CecegwW7HlrirfBkhI8I2vwu3ngjPj+ATcdX2HEGWYDf19lYGpeKumj1ZVTYyKclXw/pw
ok2jNluNqX0rtMxx+GcWRBRUC2KgZ0njDrgkGqXhTd8U0sKcaqyBfAMbZrCBna8smbaEdXe9N2Qp
ZIvPQ0DMUVxfcIDE+hKmIoim7skVCGjhYBG1oNnzP6XKQRLzJc/h5uZH6ltZOtMKdmewXB0zoLsq
isp+/MbjxaXb5nRTTT6xr/aXpZuXA0xKm/STLwXLub8iHlD+yuG1d/3LHejIPCePZcaYtH9e7V9e
xdwLeS1YazvPUetTv6CUDmHtoKxxiyJe8MoAzvN0pYmzdb4coaDSjXK+g0/GAA5pKJKyLe+AOQQt
YSIGkS7dNUiMXlDV0+PZ12k2a9ZyVXPyZeHpi62ymQ/QgY/1anad/IkH82Xb1yJMXrniWyZK+SiG
jfkL0uINFQsUx8I0A/XmBYSBtkXixohPhlw6epLzKkMkI3J4cpA4dZo6xOSyZf/rr5hIaTypUNyI
s1vaHFfjRQUGajME1RwllIF3TMafOS6N1J8P5e8F+CuGAh5EUplxAU1RWUF8TY1YT+qT7ZqhRGUm
g+ykkrMoO44OEHTWrZiq+1Jlrs3txgfFc2o7bcwAivy9TiX8EagBJwTL0GzfXAd7iwXWQ0qsz0sJ
NHQSOAyx8GNRkGqH2J2V3FEUNvUxBlLfplaCCYN+9cn6BWGapaItO9wBQUHwiSXXOyqJ/nyXcRA/
GxI7NiK6+EV35jiRp/xzbIR6lbIBSYMnyg/AwtxwcICDOuKRoAJw+dlnkaDOvwIeqmPGf7h1u5Z4
zuvDJA4+ch5O9npkYeyHnUo7pBo3Lx11c6/0ud7UQ0alVydraBE5dEX89ab9y7S40DhSHlJHegPf
ZcfI3fmt7ZYI1twyWjmvUFzhRmNT55FRt22VBuwzfWrcSpoYGVpTlK85saKT+7H4HixoOBrkiMw7
uVvblQJIlvWoFwuhid56WmVAlRoIh46Sg3ZULNBFp46H91gyBQxgfR/Z9fZiknGrBwbn67WE3WT7
CcvZoMqRPor1zza8jzs4q2Q4LdfuU8pqG40bbsuGF0brZOtoN/xr/JiAE0PzXFr+GXOJGv+nEVgC
2WjnMs1qKLLktysxO8vK23Gc0rZjSKg+SzGwr1Ab0Ez5YCHoFniTvCfBguCKUr49agMiPGTgWTBr
F2ImWNhluHO2sc+8x0Fgo+fj6CAD/wOQTKHh2FfCsgq8H0YTe9d1dqSZz7kZjhaLM7k6acehl6y0
nQfCoUZye6uS50kG2LLQbRH0IH90drvtk9kYbbXeVFLvAyidP4uEhp1PpMN7MF+1y+sKQffyvuea
dfyqwrfzR1GZzLiAv6PlpyS9kCdBOeAxoQGvP17FI00WIntVGwj88VPHCUm8PrXAnL7hyWZPt0Sq
7WV5x2taqVlqg/w/h11eXZoDxHupAZdTEyMXeSw4n8S34o+8hFynzGsyPHc0ngJ7jHWgb8B+AE/w
bQdF7+gatbwcy49fa7nldFMcsB489vtRNnnbmZBS9Pj4jYz7tcGbfy85amX3kNUd8L/GGEr0vqHQ
EaSOvUqHVijHoOY8oIt9CEY1W7avEytJ6KhdN+RHKWBDNxOpOBOF8pQ0xI+tpXM2VLL4H4zeKlEe
g5CAppfeCYy4xzoNN8dmtMXZBuzJX/+H+MvbeMyTWAeS3OZ/kV8jPpfKL8UKb7Vog6VSVl7IS1La
wfqbDl/7XUCxp55MemTUHeZCDAZN9P2vVcUi5eUs1EM2rGxDrLzRwLDSt3IpeMxFQ7Wto86CTP5c
GmtGmWckQ4JIX2qTULEFyEw6id9bgrZxF/dTh5AiTsDsM/JYEnF4I34iRAkFpKdQN8kVAVh42MuV
wbn5i5W7aD021hVdu4/zCWyUUWlM3eNzdrUp/xz4BQbH+YKxgB6AfZpDd/UNoiAw+W+srHeceTo8
NO1H46NuuznRldb1R+EShUalGwrS65i4O+yTA3jKm2Nb1RNvwGQRquuvQwoqeoeEIBagHmMWawkI
lsHRrX34L7bPzZ9Y9oJDS0MGp5r6xwnJ6ERzBxhzPzjLd1H5R9fu9mHw41Qdrp0dJfh6C3X7p1Le
KVlDo+UM4Reu3r/q4M3sTAac5UUvbO65d74eq0nqBArJvnTvxQCNdBL+tbrGVE127XOrBpjw3vXW
Zr/JjV5WfFWa/AdgV7hRo3Deyox4opp8v/BlDGDk4ZmyiaL2mguriKqUC4pqKoQLs6LgEXTI5K4+
7PAbiw8izMNL/8WVA4yL4Ob0wxCVW3m0XqGqvTkwFnMNdWayHjwf4U9eZZH5JdZPcDKsjZscjmHj
XsjyQXRjbxPGmCXFmHId/DTSmznI30kGy9QAULarVgNmcQ0nC56+GBanDw0pjSAc3VG/rNsJ+Uj5
JfnovvY/qygP07zSzF+KEfDg17b1Cboca9A0/wFuS9wI9+1XjhGAZTc+TMm8VxhaJ8kqpOEQnIfo
6FXaRPGcGtOZEUJh87LFeRpNfDN0y5lUQ3DD1zTNgGdyY/hhfr97kyM2O6yV+ibF554//sKpHGpT
TFC9eyby4/wYS+he5lZPCZ5ITmet2YL6QaikN4V69ZFFRgPeFfvg+bGIsEqUdebSTjHu/aL6d1Tj
FQ8/1gshliQTSid5aOY6Hqn7na/9ZRcNX1d2bS/j4ayOJ8I/o1RhAdmyUslqyP5e6+huYJPyrtWT
Hiudhwog8dmULInPM0FSV69R/Rnu1m+JVatGcX/7bfHwlHXuMDIou2dTEfhXaBx5oWju0Qadv9LO
bjqBbK40MdBMdRs2adniupJdqNcpJYTnpfl2hpMIUO1jZnPz4XOMx9ut3X1mlwDNrqhTrXvRrfOb
6Mdjzyqa7CZiOwZUzxF8ywuw8LkBm6lzYiSJid88a/27wwOlpQm5XEAltp570k/bXVntEexBa5Vm
JKHkpVKzatLMI9oHLmmxGh3QfUet08U7ktiuClSwhBiY30zZA98FRT5ysPyV8TTKaCGODkSMV3vi
VKTtU8lLsyh4Ui0M1W9UTeIgLlOvmfrYxzqkaEjdM+JL6aJX8r+/TjrSrvsRjtpMnqX48owMS1sx
Fhgkeyb2WFPd/pE2LH1s+8oQ6Mh4RY8umYCJM5M2tJPjNmRQHl7+cGw+5jEJpeF8Nn//OHFrG8hc
2LKCntc1NV1RUMKrFQGhVxUYCLVtPjsat+FMiEGljSO2kRPGFaQI2a5vg9sq+0RwUpZ+lsDrJ51C
jhchEnqRpy/HHz88a9hhr+ut9zv/lq6H97nZY3Mg9mKLUbXBZ24Akc8CXJwcrnXEbW55EufzAqNH
SF1+i1Yt1NQMPgi69d8u3lDZVcsKa2eQaGx68OZfKtRKS0lpSyNKpYrjSMF7kp1KydKSYph2GJ+e
r1iksoW85SX5kQPLoZe64DLPndypYrXgITMlsNNREDNWiY7Skl8rrA3d2fZwI9pf5nizwY3+/EYC
nf3Co9K2Cf9Yfwod+Zq8MOKUlvnMLLaAxc0yGFY/qzhIK9tck0UqJvNHrKsqgKFXhxqAeuRJFupA
tsP2wVe5dbCu7K0uQSpi9kCY6DffrwWSDHUozn23V466fytuDhvDQUPj9YKavdM6vA0D485SnA/n
kdwEsD5GDga08QSLz/dbQ5+cY9J/23PeZL/EX+zAB2HPOXCti4UQ2VCAHZ0+y8/7NWFw5K+FczTu
2CukoiCJ1WcBN7r7snvY1Z6CKCkow7PWH+BKhtS2a4k5Fj+OACAzQv9gv7Ta7IiZQNeY1yN2SNYr
5JUNO4PjCEXlLq2IjwubK7NDl5/3Z1MYPRpdgX2cNkhi3Do2uPoygZFlOQW35K4JanUzllXWOpbU
nOdNswtT6MiUC8tgu8eKK2wp0ccABzqLu/koJ/qRuy7ZElK0VUqwn5Ic/yu2s4SeGeWYEgxIVzho
4BuROxeANJ4sWWc80658VCniFraUsQGZmCPD6pagvOaP8hVPGDJ8WUXh5Kdin7Cq5ibpLMIwqogq
CiSJD5v9m1NjLOFbHjt4cvg6LXmRgZs0Nk5BKuHRMBxCQvL1bNuOPRYws5xZzaZc+WR0Gsefcqtq
eF9IVWB1MNHuvy7pTm7NONwRps1srvEqz9jSnsRbm7Gk0RTj/+8c+87y2TvF2F4SVl0sqdlyUJ6n
qfFLHJS4tnrUNeEfC0e1dAGHr+5ChY/EBV7EoA/1oOHFDmHYwUidY0KdPUZS+2meNIUypF4qNiB+
83AZJl+mu596IH8Z381btKnFooUWAPZMwYvMAkPUavCS1JDGr4F2DbfM9cej2A0L7et6WyejTEFd
/fpPbFt2Qhxpnp/3J9lpy+BTZjPVfo1VdUsSrKRnn5cK50nZoMGCazqTEkPmm42gJ/SyItkDO4EZ
55ulpDUqNf53676KEjrWCu3rtdGkFkv01fsYl0BB7OO4z+Yz4xvji7YkC8W6J9gwrpsQ8cjnBxot
YqA2AUd/PgQa5HDSvz5/nbfVXmMfdXRWZM/6+VqmZcA76J2/PSzlfZQUyvTz5LmeIKKw5DbY1+XJ
l2TaT7dsowEy3VqAgozNC5w1fm9nRW4XqjL0qh9KS61aXOsi0sabHMITJq3GUgps+wzgf7A/G4AD
gSR+UySdJaZ9RiW1vGvL+Ge6xbgH6rEyevDdY+Yj/qz9xN9q/z6MUymGOcnJ/Kk+mJz/YQrqcH+p
nnSgaKfUvlAUONwsPRqXHndYAUj4GnPPBQYJu1yCEBtCPYpBeYMfaxlq1sQFyZ9D24NAeYO6TW7U
3o+PzTScLD6Os4V4OfOjkXsVA5DAGy9MOFr7jhc2NOlIB26X/qy7pY1b1c5weqTgU0gDh4rMVFTS
MC0TH5na07rZHWJ+FC3lqxjqDHhxJPoe3jb1vEn8FNBiTY2VLgHiCw+IWLKpMIlR5v0qANk6nTfh
fhEP767JYt+86Xx7BeJq0lHzn1pijxmXFZGKs2vd7MLMPMCxlxsO4nBjslG1uFlahSynfRAh6axW
HjaBagPzyRV9hKKSZFCtTnEIcp4MU18QlZdqcbjNod+JnOK1xD5tIO23iW7AMPDlvrde2LoozaHm
MzJBzBaXDlOgy+SWLC7lNakAZHwpuGCD2aSRxWLiMdYef25aqfifSvQZjQsXfo8VLR3gKu8IP/ZT
I95uiaiSLkepyEDMYkyBJMYsBOZZdLokLRPZwgEZ2X5QsKc6+Img8t7LmWqbuVYk8op+K3pIa3ki
qs0ePQ8LXpKftrgYaPVcn1YJEGiixSmGPBMS9A/wsCfVUhh7pmTiHNpZxJxknxW0xQ9kVCXcOMz8
qo6tCcV+df869KAc2vZw5gOXxReHh7qkjbmYONd9HP+zpx4z7yMVpaiD+PucMRVlaNoAyHKdgavx
Q6EErGT6wycc2iFIE5UHYY60Dw3tbwXiyLN6Fq6ErCVCTlGrp8wPsBdFhZ4gWQUcTO5e7uFjwFL2
Qy2sLnqQFIoSEIYkWYezcEh4YmVghETVLeO5wxv18snFEL8zBhfmhHsePC8kZwMDQA1eJMgfHc8D
4FBPW3gCpXcw6QQIuRH3psw5YN2+y5eGo5sIe4UO4FpZsfdiG37dlUFiVE+Ju1dz4iThDsazYmoO
V5hyQFx0tCFarzo64d8kxlBy6ooO2+IKml+06rZNZ9BQHR8qrBM3AMrmjHpbmFzBE6EleKi8ET1G
eBASyq2OnMBR/iVc/K6Jp7+nVhpn5Zr6UBez80y5rFwOEM9epEww3vwTjWY94Ek5f+kIA4/aVyM5
To8GXY1zZGV7jZh3KadU8gvKBOwmJonV6f2EJyHHcnVPW0anlgLYAqdS+yu4ftOKuvrHYwHWx2iY
Zqag8iW01ng+WWXhcJw61yOdFVC6emzjOKg7jIG8wy5ueXpx/NZwKywVQIbRD3uyN2x5dKoOU3zC
Sao8W4WPXYhdiJZJRt/7ZRhnGSTuuBWKfiHMPOgeKNKCxa20hF0MzLvFpeAiARQfdnxg6kPkeUom
73SoVY5KWdcUCwRlYxGr4OFLtguO0/4drg2OPACj3rZwqZYTxSUUiDD7IeRkOdPH3VS0BPTAPLmU
X1wKngJLS4qJx1J/swcB1gZzVWres9SxIClzC7zMOgCOwpAXZLmotSCrrxBEzHQMQZ/iRoLfqg8z
na6NJ1x02xk9a8eiryDPVOOctkOmvW5ei7PxrBnJxKlPfGpqUx+wLLrgopQ9B62v+hfckr89ysQb
zLoL9pQAkI2opHd0/7cnGxet8WXG0hW3quAOJZECN8U3a35FGyWtEi8L0FwIMQpuJawDw6iygTHC
cgb1vBbZ+m8IXhNI4reEq1ygc3kDaXXCPcz7n2TxyBJ8wj/rkCjK7N3BySme4mBkxxtQrOxE5g9k
x/VlwxM2Y3kccV/M1D+JpSMuitw+EHT1agYI1HdkU9u0MIWoxaFSrjC9tdJ+rrHAzHbE9osv5YOV
3iuCydOu+Y0KZQWchw4OUV5ckiOMzWY4BEsr7CbVgXVW0zY45begE11kW+RQfoH1r4T6E5JDuHSw
T5iqhNM7IcAXAbysBnuk/MnVsfwVFKgcw0YClGQPUJxiTSnv3z3XHIJeZtfWVViJJTVzrkAlFj9w
UHIh7jgh1nhVWJ8THqwfChTF9ItXJ5/Xg17XYZ7NeEG+paIrlUHdq4EMaBioso5ToH4+p4FsIGsP
aCj5KIQm5us+7bs2WJfjkgwO1mBxYCMnQJzH7fcvH4NIcmG8JBy7Z5F0lPz/9D4bRHVjZ0pHaamE
2rGn0y3QX2l7WVjXbMdP+HmIoK4KV8J+5Zn2c7tmQ9QgZOSAtenC09iXl+shpV+t7nLYcqhMeY+F
lxuJdwfmIbM/f+gwrOzZfe9MHnPT+NhQOCxCB98Te0kNaq9n6YTPhyuPknncWrrwznp8CJUgNmZ2
LvFRnB/jtgUkIzRqCEa/VBZfDVsqIHxDx+vZyEGiw2JKtc8U55ol2WTALsakzm3N/gCyV6dyCNlo
C/3c0+eQzQzLSFnUkpn8sExX5mA2F2d3xXI0VoyAcQ7FqZHwpsvKcNQWS/fTcmAfyA8X6dXTafT/
hupBZnz/Id3An1BIk1XTqz7MUVDEDkaNN0dhn/txqMkGWQltpKQz3R5vMdWts1FTU+zwftfJnH/1
hozM8yeJ0y9hjKNyHQm5FN/JmMsDSU5pC3A/Js5I4laR+YdQV+jGVVdva/vhTT5M+8RA+zD3z0tR
9dkShNAruVF28KF5o447S79Ffc1btLzWdgylAfhB8pzDpIwuP/1YY9QjjLVudW1HaruIRuAi3MeW
liwrsJSIjk7VnOSDZjjTx9z6zJ4LSaO26HwagY+jNnYi3s4MRjjCf7RLDhWsRJPoiqnE/8ngvjWA
SMiQBwjkyQ2knxY52qJG26CG86Ql81tYOHZRCzSI+Z7L/CbuzCBlP10VQlmDHARhpG5ljxJ1My2C
aXjeOlw1tKmDJpu+QR0W4QrDesfQP1rwAiRttlSfYZQ2TbtkIsg3z11dpcg0o3LGP7G0aRvmiH+T
Q9BX17PgLZbMuPHSysKVAgfb43giKOFijyNPUuoS3YI2emleaHwjn45IFTN+1JojtXE+oHS/Jz6N
VLfr/kclDWD3en4V3amj3qQ1LAMjO4u13kWnmpLr747K+1MmLaZXNBZEpbnl35LdEhz6/ODHFKtL
wUcmvVZ0pTPDj/DdPIGlN4/SnPrbcPK1L9abT9/mmkJ54OQsIA3sKdefUP4qR5F1dBbOmX6RDwzE
0+YOfZ0451AqX59bHDXWEKVyENXgXxfmSnUaTY7X5LTVMual3k4xYcwzDW3a4dJTDwB5yKW3hJeE
Z29orcsZh+a0AHtPw8XcEAp0n5DWyaE2IhrsRT5A097Zsd/SOgNKQQTVfqMbAfjyw0CjMUEiC5aI
aAlPuET9if8MpnTjl/YpuTo7lTLr1GMyxtseW3UI2QEM4V8h3c2NEW8ebA4TjRqJkimYiGqcl+V1
nhwxprmP7/OAlQhUmAFHwUKlyKs/Dwa0dBLZwZVBtqAzf8Y8WIB9PPpuKU5RYEi80IGVbK3U2Zmt
81dLUTp4DDUu6mfAevTDGBqpnVxwTyZVhSzdAoZ5hKgXeLhhaZ89wRu6+nnunxj+wrB+fAdUJEZF
ozorx19x2FZH6WGjkfM6erxoh7EgN2hj2y49x+cTpUPhb4RmYiLFVuhTWeceqqdv+FcFUIcWRC2c
PPwfQxrr2qjJhij3ladA2wNzttoGqcd9NyN+WEI8v1+Vlm6gME7Q5MuGBlcUZ2MutVxyQpwblA0t
t6PjGOHLPyD0VE3q3sfSsvgKSNr7MdK110yOw0SYq41UNfkohiGDU5byhaoMKXogMF6EVVnPU55K
OLH7mvNTJ8dyZ2jPxoAPrYhaS3cI/PFYOClWgyfa9+J2ZyJctIx7I1YkisgUNIETg09Gpn636Gb/
npYXTAzCgRsD09uv3TkLhSDVyLQXBYOlVBoXgpmGrHuORjBeSTv73e8iu1IYWn+0L9BgarnscoWt
htEPzJzlu8aCKsdfQSw6hmZDEtYWI+G7zvFE5I6rI0PqoVPNa1jsAkP+J8rR55BxNtdgQpFys23w
gOI0N2Q8A3z9WLaGkuU2T1W2fU8Pwm2tEnWye4JhPDkD6YhVg76EZ7KgBsQooZtlAjXflAmn6Rd7
/zWzqhKt1m73KP7DhU/KfrtyxkfI99mzKF5gajZlydrzMtHytyRi5XzFrzxfVc+lbbmgkJfMPGG/
pgzR7bgf2+78kIVV8HDYT49y0/46ed+6/ezvlLWfDLc1KZ79W5pRkEYmW4flyjFdS5XiZtXiT9Fp
Burn20UI4rvkkPEpT4ncEg6dw8kx7X5uN0PbeFH67OjXZT0/WCHkCsocJPpdhhmOfZ4swInKQh+Q
HXdeTyoLowXdi6C2EDCAdqUAgTE92w9Wu4BWbOq0urXInpCUJWOjUC5r0CaREMO20iPTmEZPjluP
zxair+P8GD0t+DJt0ilD+8rP5ZA5jxrflZt2RRzO8OUe6g5YB4hHn+aJjLXMfmtxb++uG75rH4hb
kZppcZ6Eg3EznsPlTTooiwd7qexo6RK6nySj+YE8zPuVh2Jnvsi7yeZB3PQe00Icr9zgroXqG4hS
ogy6Cl2+Zj6FsC3+dSFkZJGGU3bH12CkE/MO/uV2GXU3yphp6oTm0rAn7CxA7Qd+ZUk+SSGw4n4j
nROGxCuveeRYBw1/oySS9Utp8up3FlclkUk2kW1sCEqA/jcggnwcnDzjghZu41zkaY/G7igXCJf3
E23jguYidD3LwrL6neEeLztJwKDaMgqbARWzuhZRMsqQ37wkzp0medkhdDa2B07hvgY3Pi/GOSYS
4QI59wYw148wRW10073EBgcFw4FZ+VHW7k7Qh6DAGAiJ76JHRp8C7Ds2oU8HI/x1BSHrkcybUlBY
xuXblwcmx3Vk2rLRv9S2wnvf1ZfiLiU+KiJSYC3uVEZI0L/c75uMHh/Qba1jPTyZ/UxQkLOvpo36
Rj/pS2GcOgqPeEKb4zWGwQXO8T/ixOgTxC3Rg/XO6fTOT3NxV38nqbgMIO08kqrVM1+jzDD6Vqyk
y2txbSV7a6itQNxA84eL3WUGhqdfa9W1Wsm3UslcqmLpiLdmqgZC7sV+xqUpoAp0UTDtM1yo5+Qf
7zeCUghe7wkcVtsEjSUUaMgswNo3iaDea0Ef9d8CKiD7o03mPtEOsLLlgPFX3NNUI6w4NChAJe4b
qQzCqJ365fb1nQX9tnz6iypHAYGmR0JpQH2ZuZ/scMiLXq/FNCMyVn8TeynO9GIbhphKmaM0uFNK
ppfA07PtZe5L3LSnJz3gcB7z35qiQE8toSRaS+ZQ4mOqA7Mdwxq4YIyBoCpajCSL8DR1mgp08FS8
c4PWbeTSXU/1NZGVcV7EKgcoU9ryVv0KyoVOtkq2cY2rSCkN2/yCoZ4kmrzvL3Oc2I086LowCUEW
cEZZGb23V6LNB2eQyhZz5kqLobdIvyziuiowf2YvR7xL3c6q1xxssDKnwRotfbnV1XwiMw8DHu6X
yr2AQPGBurwswo0ABStUQqUs2yzZB6v1tGIrkqGytCvHlmQ8P78IxbSStF8zFXjf4TL0ZDc1G7tV
Z3ZG6GTXnb1DmooyhxtkJ8+VTFz+uUMDg2NTpKs1WWhHunpeW7yuyEGG0xZ544QluXb2bZHOnmJE
fcGNgJ1xhJ+fyUcElRm2cTI6IaP6inrwck+mc/aGdwwA1Sg0/JG4bmY99CNAMP4xEiOQnB22IRrh
OZ3tLS7hxHMlsIXrxidICWsMgw13aXLMG0UaZqBq/x1F3av6Ta8N4eRnoS/+i0D+mrHNhcsLv9YO
Wir/hePS23jjgRRTvsuEkzVqEFxNUSdDf8YmN9jslvi4g74V5ooKs5j7E62ma1NV8LeE8vE4rbDN
CzhMWV0NC7SZSXLAAZFJtxJkZOcm8YdSHtdZNR1rzMc16F7Cts1Kdqs68CscO6UZ+LpJkQUxQlDh
AzQ1DRhxiqRA1l0LinUFKjftFCdPgAE5EpKLO33rghq8XdeHhW2vba28xlIwNopwAX8/59/IqkzK
pnQB7yfjuijboJ249Yjrgk7lJS4FfpNicoV5N+Moej2NnkS6RiDbhN4xMgk4kXKcbxlHMM9lGCVL
CuBYUusihXQAQqMpTT8+Ub+wpqzNNcf6Xc2pdj0RN5fKpg/1nGByxmHmWOP9rN/62vnGG/5l2Vb8
HHhEPspjyUsERWNHGNznCDkT2ZiWYSC2HZSRmni+oYxVhOW5MY7ru9jmwmMzI4U5RK5ib0yHggTc
dx7ENlPIXSOd47XrcURbPScegaDxO7LoLsnfptsNayG/LiezuV3sAFFsHnZUV9x9mRcXeuUBoIrg
6ksvdFJycAEZ1zq+IvpN9qCI6kdpbiuvv5Sk9KbdlGaurOt+XcNb0w+NWo98HJ60ygNsZ2eS5ZFX
ze7ZLjVTuXWfwIS3y0NyF7VdwctBZkelN9B6lZzkh+RIsM0mjA0/6qO/3uXmSNqQhMsQQV3tXONT
2CLrTwTFxd96PTsMxNjoYO0rAPdeichkcdWr+ZyNU9Rf1lLZTTbuWH5KKQv3Tpxmmyu5Gg9q1J/t
5x7/muyOQcHgtyoUpTEW1qEbIcuyDZm/5SX3g5e/ydGzb0vtuYVCmnfdxunZngTFbInwVsayLKB3
bzigh+DFz2Q2yN0wKfolEmyftkqlSl040bdFFh+1KmaILVrm+GmEy4i8sw0jBH57rsUz7pqE3yLk
Gkq90nPyLDEiIUGpdLtPmhU4kbFAUpAg8OQHhVpx9v2L9URwMePEAGIWuzgIx5x9V+jZ6qfTnygN
ji6NwwhGwZbWWofwYovUlqiMx6vVVVwICqDlszdAHr67ElxN4H8BbnYPgZvc4j+9W3lpYNgVcnxX
LwAYwAnx31OA6B1uO/hI8oiB8k7g3Jozs8IoFJaX3vm4BeLziFSvt+uYCUNgTLJidJG+PDGqZJpC
W/0dmihkCrJvv3VRgvw5losyHmAg+xP/CUJwP/eJQF72TKuONACPBNyRmltzzRHbK+4+k1JdO/Yg
2SZJMACYiZ3DpNWkoeuAM2w43AmU+kwSEBS12bJyC30ZcMZDZU7wtZnwgx6wcxuOavM0sXj8RG1b
+tfn3T8DLc2ifAbGls2/ml2ZFqDmIGSZrsXtxoswKE/H8JR2cR9k+1kPQ3ugOPXtQWiNXO3oCY/g
VKMW36YF1pN6yNW+LP8B+BVNMZQLnSeITDCIkVEs0dKfapQtNTfwOceIR9SZXAsRfKePHqyvsCBc
76LKRIjOQec4eiZCC+JTgl7hGqH5Gm1NKtbyIzC/q0z8UIEWzdU19s4kLEyrgOItIIqza7Jc6dOZ
Bm+F4zechKW6ewWpkN5JH4UL4TgHzoBo17kg5VNlPbzQwL7DUsoELUE/YED5nzQP67+HuKSlCYt0
GrPFIXuIcfXWGyKSs8CUpcplkpsG2ARfEZVYuHPVod/8aEu3pamDufEVmZL8Isl7LqpEznixBDnE
tL+hERqCJto6bZwzzbv69pIWNBdEmJzCpFZ2EL9KF+JropyP8AR+Bdhm9LAevVu/whCA7iYOzx0r
vk7Sjv+7iZrkhchhajWbCxqKEeHsxpANModu0JDjnzYXbMuX4W9dlR0UsgTNownZfQOS1IxZHMNe
biGHbwsLQaiDeSFtsYMFQHHmXOJhDLegntFQe1lkdzNjQVXTS/OCMCt8vbtGLPH7GjPWOF42f+Ic
cyhUdsDTvgaysmCdKoEOvErgOPwP+xeoBAXxnpkJWEESIAXacN6QF7U0Z9Ny5L2S8+Q00PBVkPRh
bMYG5vh6J0a/PYjkdvxs4lrLlzdXEfGbfICIfui6JnQ1ESww3vmTEGV1uOqnWB/ciB147T4AnB94
AXu2+zD+tz9WU8mziN+i2YZdILtjkN9KI8OiB07WcbmJhoovgoVwbUENOWvaX5yiYLQGhBZf0Fdz
q8iWhdOl+EcNeU4UZ03tNv79TLiMO+7whlHF5q2JqxaEKPwEyra6og3czcx/SrjyYoBR5/3/AQ32
BI+n7nuJ4ozozUMfyaOtFP/rBWigPgE95Z159Ucqdba8gyHfMjjRVXRQt4nfW5Zu00QWMvTJTghF
2KGzEMIUrjCod/lvrAojqhQR8vewRLSbgNeQAZApOjfb4trHkb+MwsfLgaMkYOeEfTcqwnf5lYp0
lvEzrmwsB4d7DOVGwrCsaqj03ClU90OT5TsuD/NBx+xQJ3ypt9LP/RoZfDlvTcBLDmNfutao3AEa
yngd8gC5w9lLH0QHZj2bLHaGHi//E7ZBa+OtdAQ4SRIO4oNz6uaeOW/kEL+Rh/qLly36TwLWzXeK
ElKX7mlaK2UKjl9omsDUKLVKe/h5LJ/+19CDfGXg3bq9KQKxv+THgPYGkBiMxS/CglgBXsTm4qSq
tF/EGF836W1f3nWTFVVn3WxwIrb1+tU9n5UFWEIGBn5GXVPmHYIOixnpLRPpgVnFd3GVExo/8Ao9
bRSoytyZVF5/+KUi8RpAZdn7yAyt6MLFie5lVIwzTgi2PyXKmEUyQhVmRNvkYDw+O17ZK4uontBi
S2cgHw7uxAajcYBX+155mru4/xpN2HrumNz1ewi3VothGlwTaJWEMBlWvONwbP9lqGrNJWyWW2VY
PdKqYocT7Xm6g8fUOFfXjTIlHuW0n7cDX9kfKgbOX4vTRREhJqJN87oLjDkomkh3qf6mVSLysjii
h+0XyVRwe2TKsKpq3ZTw5z9bRcTBwqmdqCDH08Tg2cgBlUi5Ui8KmwhKTZWDBYUY/hCy202gIvWu
4mzjGpo4vgV4H9IOAHlJb5G/WJSCdERrEAXVUfgpar6Ap8X4d6K3N+eDeto2LD4dTBCeqb/8Ghv5
fM/V1ExorTYwJ5jX3ik+kRwO4YP0wa15SSuuIdeR+ZRO36NQ1nkpDKvrJ1MrnfO14nF8XgfABEjc
8szDdbNMBRiwZ6GnbmTlQ2FbPjqSt/BLVsd7f3R2macfUC+jHdMc1iH4epfdyW2r+6zOWrpGMoP2
E8u7n5Y4ol4RmpJDEcxH1BcyPchbhwP3ZTIxF3k1oz+IBeM49fNJ+cTDdtdudPrXI1BNhdik38gt
eRbaZyAKSbwSXjFXAbA/cQm+/WrqbU/jjkdPhnt3f8XS4dl2ByxI8ytU3JBgeZHYsRlR3d/JMYg0
T+igOjrWhRJGBGShg+d4ooFuyBH63osxKr+KKQAgeoJEKFwfSc5CcIu00JQ8B2OzoFhIL9lTHRb+
1U7W1K510EnOCcn3Iv1SKBReTcNSkYH8L0Bb6zQXmBBcMNyKJAkHW5UTlRKe17feGNVrUASjxPOJ
93MjYYOCub0IGFyo/Psz2X+YRksomRd0ywbq+tVGBsEib6hsEYCfdnIbuKEaGKFA/ENFzXWuVLSK
/pxZ125T0/OqEmPeoXDHblAs95bb6nElDIx9lU3R09riGN26nq9kGMPGRDgySi97+uLE1cJuRLoU
KbfYWZkWEQM+qPC092NDMAeUc2x7v5Uq9Q59tmFk+FYWTCGSZodzEjcx4Dlz2w0UxM/0/ur4f0Ln
DapfwXGS+AmSTjgzLnxBoVrtnbIJvFPzXgckO18IiWDpq0UXDWL3e6uFgCRPxBmFWULsr8FjcqhP
6634ipel9Rtbh9Bhs5cX+uNaOKqRDtiWR9FRF4F3a9GOZpwvclsmXpbOw2OT5C80lfigDyiW1IHu
cpOKKqBAikLqUtBJBvJDOME4rdw/YiI1JXn6Kl0mZvUwfgvOOKwSZiSXYsRD9aQh9cDIa/6TA9fn
ai2ZUk0QVETVv7V+Gj7tjb55P4DLomkQp9jS88eBOh0KzdYT0AQc7aATXsxT4hG5YVkdayaA4uDc
8wxWlc1luqftWObSSNbdnkhEHQ8T/Mm4YaAENqZoBAtkoGXMSpACobsk2i0771+w6uqIkvdBUS8y
h00GnXuC5/nrEoB0GubsxhfnrWMXNcasm1ZbRtW6Xq08ZdF5DQkH6tre9EQzY8nlp3v744hNOrzY
P+1uD8h4V31f0jBma7wokx/LTROgTrp77FSnoOa0BE1DM/KjyiSNZSd7SALaxGpQRZGO4/eOANB+
RWc3fCPNHC0fnZo0djJO8QdHat/Eifk7upv8AYQXvaysA70WjCvaCAtdz7pQzf0MUhKz0BXVERUI
91GABZss6t5a6ahwmYtyELA6Iwr4KTP+5lxXuWwfewOzxkRY4PIXgGRC25XGh9EB7Q2JCgKeaYpU
S5vyai2m7nS6Vt8ZmyNU+HJeliH1EikTA/XYgg+CNGDAZ8Sh2yBWgXizY2m5eICsbY6G2R3ATRbR
qP85u+t51tnkX4k3OHYCx7uZSN2/gS7mFxrvC8ZjLIo37rU/xZR5YoqTylXTMoHrmbCYPUId0Wlg
nU8jWVpLJjtLZb3tpeCE+p/Ty22XliCBTlNqMhY/EJbaIpmihsUCLFMUwy6kzjuCb8cXF02bbaTi
alcPu9dkuKvqBniqabIyej/S0H1nCD3pavxuJOtpy2xtiQzq52iKzjFBcxf9jllAHQXH7gtnSE5l
rl7XiW929p697atl2nv/dA2UBN6m/ajSgxRbxzrws3zyVBgEoP3LV05czW8SLIV5D+fsOU41Cy3w
AVSyC53Q6EF+t7xcI5Ush0kwMWjjm56JPm/qSergIMwMmU19BS4GJy0u8K+ufDOD1lwRn/VlB334
vDlvfc9LOvGCaktL/e0eN9xZ3mHu8sx+i08gC2Acyc9bfLuL2fnK48fKy5NiDbiobq+3yGZKpEWc
WJyW/rYIXbDmKvSrzPM/6gercoh5qQt7YzftWiX4XXBcFQ8oOJ7DPY9/2xLfFXQSffY/NbU8aena
lM5EMVl0zHY0Ax6Hg9F/JEpBqNNm9COW4vNLboYmUI7cJgqdwMVrnG7OogUGu1x8rKRoek9dzRYN
dbQr+EVy4rN6GQ0VlJ5FX4MlWbeyHITTU+dnKDiN81RgRs5x3hRZJ0ySHVTRBqBWMEVzHiftd/8/
IYhUVZLlLhOunCE9Fl7weSK0wpPFqLy1HrqyH+TeQ1LJ290ePQ7cCZ+M6TYJliYTRJ2+LpDqhHVq
YSMqr5wE0aoU++wlH8gYXJP5W2eBgLcSwc4fiNv5NUQGy7bI4Yney98pgWQGZMSJTD0cvrHgEq1T
gvCEuFDdOrAOO+aYBOwGu+C7SfTm3XXFeYJjy4QPDPh7m/voFkfa1Q6Y55jhrZ8Xuyi64DlSErwx
YakFb4qSMfgqiH+/y+XIMVLTPrheHOA1ePtnrHG3UW6BW/CyLpuxx2QUPTr5NvXDeVK0D62bV26k
9RcMr70qBE2nDQRVw1Fcv9pWoGeKp9o2Eb6ea0y2HrBPFFFgbPLt2F3BCCeGB/UqPpMfN2pKMXQ1
POYrr/emcv7S6EVqgsYdDnjh7ikfNZiI5tzJgkIqbFa1v2r6rUi6s5gntiuh47rppSnHetnqSki2
d0naVeKsPlhacN34SfyxeDIj9VZFerjZdSvfJN8xo8JPDCfLbt85OVpHTiTh6inhkzsri42LTwd1
/t6XrhIrI9UtYi6tJhQ05A7SY2H+7v6GR5WlDpDePdq9nPxyG5rk8A6NrJwPtJ2G3MLRAe9fdqAr
JT0MCcUakRq9cv9lMzhK6E/bfjr4VKJXDs9tY0FMUbO75upzbMlZz4x0TDnKm5SKJ3+6hyx35YGI
8gdWfLV9eK5hHx/d8Riuymq302xF3nQyq7Q3OF4X4vXgdKlbXHbCaz4nxYlqdcFmK/IxkWce4mpU
6PAdUS5GHb613QTTxnFLcXjAibRNSMXOCt4LlpEs3pDmGISlds7VUwUOZ3wcRjL7Lsvo/lz9WmlG
HUq2Haabo70Y2BWO/mxw6aFUlcRmkeDmD0zOA02tP8OfbAbdL68KXmFboCZQNlEIGDueY27Jb9bD
vhjooaCkMLtnBYRvmmgBE/tJjH/ItqjufKJ9iytlGfhsXPiVlMf3u+alk84tpzw1H7zGpL+Iizdv
JpxH4CSAJ0nqap1/+QdGYo36rRxuuXGzBw+LTRavb9BWHvdh2rOZklqgSFxdWAFcwt+7II9N1nPE
eqV5NXNDHbxaiyxjmFlvyw/3sIRQiPWZaiLlzwaNSU1shEv+z5a26R67hT++b1tcZaZdxcCQNi97
7X/w5w9h3IaUZDZot85vGDV3T8fFFSQxz8drKDIxRsIaG60pnVffEY7JQEXw+HawTY9Q5ew/B9NP
ZmahHbINugTSo0bTZxlVqgsjg2XANW/7iPVRMPaHigjnb2F90MAEH294RJ2PGaMbSBG6mqK5Km+X
etxDrbIeWwd46RBP862nrrSlFdMw+muBbNRJOGqxFDMPLVWJD2+meXH+nt+l9udsCFWAVrUI20Ye
RizRtD9EE9Uv5TAYzHUrORw03IjcOFi0ZblkBGcykY8nJlE7gCCNmHKupumqCmOhFev1caEfXV5k
+S9ng742x5qbJGtXkvQAJ1qRrChGKTFzNNDSpamYpoZ1aWjY09krY5lwCflUp33EzFOyJXgtDh03
LIRpXbhoU8S8Pbc7DfT4/q2/BjD6b3XTMhLOpWiTgaVoEfqY4xKcuKu/bEkGAkNebXCddCc/PNlj
lVlxmmmeZ6DCR9X19rmhsCVm04+2lAowwzthEQIRFhTcuLBwH9h8NxM53aiVGyd3+AJPT2z6MchI
bak8Lksj/GkWTTlZP6ICiGNaub2NG2vyq36H+2xiUQ52jfQ76J0klP6s6+dvoZCHDBJ4FR7C6RRx
DYlOPETTnyQ+L725mLPWw4GInHYBec1Fc0QCXTF51sXdPkIN5dzzgbZiBenBSXc+/6zyvVwEFPzw
EGHofYfNGWJPwM2pdEoV0M1Ie+/K/EHxEV+QcP7gC+a3oMYCUsMLytmkrW9y3I29acoJzLkD8J9F
xIV+Uh2phssLRln2KHp9TSjTYne6JeqUzzTMYH5Ax08rTDkPPCEc+FhKFV+uG3IROT8CiNS15OhE
Cv5zaXrf0M5ErQGq0x2+Bek+SLcxZGNE/0HCIA9glffsW+Gbx0OdhIbEzXuGEGGrdKlbeoRRH12c
qFDLyu5EHXKPDwW+mAc2m8nVo6nbE/i7zoFHROgGeTxtVJLyvXgWdLSDkHFvH8LJZ72qv/K/Kf1m
BZIBC95IZhnTY6m05ZN5fhFbFJ/pud47bGsSzVK6he1pg6TOwnStU0ySUUYSkSCvzaz3yw1B7oqL
e1bxkXd4U9XQRvNSYaEXoN7nNct9Fm3/slhc0KMyIU7f7giSQsnxFCzSIrxOKCvSpDg0e4w7pEJK
9TE6T3qkfKtFhz+r/DoRhUQ4Z1/CffpS1ytV9ALWt6fl5t5pNmI16nKADMs55FIJ7KZlJ5hVqsfY
BAoeLp5AOj3Ty7+yFEYn2ruLa5G5IAUS6gs0Mrqb/B3mPZTs3yiWW5v09hKTzeviHE25x7uch50e
yn1oeBe0NgOGoRW5qGt6wjVfZ2nG7qPr6eCP/2z5nC43HPCLAvAW4d5uw78vwzptT+iLHwJi3NGb
p59CGHlYK35UfhhnvNTzfyWdvKI76dwnpSIf26qemUmkoUvbxOobfWuRWGZiLiIWa7taRSzVrbWJ
lzW071rKg61B2Q42J3yMbsTwhZkqww0MSIH+q/CwY5Yy5iNW3j8itN0YdHx0d0rg/8xxPx3YUEWU
+fFvaKSHIY0XMR5df0fVRVjXYhf8N4r6Vu5IqDuo3gtJ9Jp8dMuMmbvFaIATPORfP3GL+4pmvAgr
rn5FRFJeiQ7/D/ljUZ4/OtZZmDwNS1ScZYb6M6mRazFoxXkJtceLtmMg7loQIh/TnPBQ0W9DFz7z
qmuugOPauq218fp8Xh6jgmkVypHYkedVX5GtoloYeiFVnsl/YlPuHFOExM2uXSAt+t5mt0/VvfaN
awVXW+MQHLpGQ9825egbrqUM275STJiCapyU6fgY4cDh+VWfxzespV0j8PkWmQ1wbyOAhWjIOVK/
hMc1KWbUnD3W1w5AGEFR8G+flVRAR70WK9w0YRlXl64tfwj8s3i2nSTg1oKilpBtH916vpVSj9XI
Gv7RMLEr+QH5EUpHjgQ8ZkkoVt5HG6J6Pp2TGvHFadGem6j5kHuaPtYhMPHOp22vHNxz/A4a0PYn
2AH9XlWsKnvADa50G9suWkhnlx0ABVvinwJV0kt+FxjtCsPx24i4MJe+DdmvdLh7YyUQIbI6wuPP
kg+jLBZHa25aoH1BXEx1JPdR7aG7RNQCNa+fyvxvwPJ6pVxu8bjp2oZ1aBdkGWwoZ3B1wCRWll8/
iHwBjgY9LrcQx1LWtvMiZKSQkK6sZwbfujbrnixZyydyz0d+ISFxXAtuA8jtYdaxte1aoEDz7lw4
yejFYPARSeZL2+evbM6+rsRbiWahEiESkEERKqz3Iq9E9xhdswUCH6ia/f7FoUeCVobsJ/BbZuoa
FEpsgh0cB7vXJHNInjzjmhJbRrYvZuPENXodE77Oxx6eSyqvFWIedTEM/fFukGbNpbnf0ZnfXQyu
q2iJWdqOC+WNyMuvRMQl0sjy2MGCHr+X1bXNcsbOinO97rY09FIv4ejdlienUmh0fHw7+LWUopjC
LYN/kcr4Cdc/9wVuDtWfn09ENJW2t10RLyfmgwONqDUMZDQO+sg7XaRU+CCSab7ndXjvaoFHEaAT
8sPCNljVatxHXfSR8GSmulHxVAXk2yMdSAU77Lj6QUgF0D/U9Q/RUHVAFu4ng1YVOhexGxjE2qBq
6ye8eMo73eLSgKgM7rDiRBA9S9rasQJq2jVfWJyVEwotBsUohbvgLsIqBb81xkAk6DPMGUzSL71g
F1Br+1oXZMwuwjJKK2DRv12ygeysB+On3fdP9RBY/r6dyGK90vhW3z3CbPxFgSWwe7gpm+JRIE6M
n/MGVRedbzCS1R2ww2HB/bmYtGuKGzQSO0pm5X/mVQ0U1HsM0mMhRzJ6CazxHCqUG4Eu9Gb5xLgl
X4CbQ0n9hGiqAi0/sn8JRqG6xeP1xOIavaj7ofFESAW5gbk1v0O9KDfugT8TchxWnZTrQ3xmSYwN
7KHDqVgZYdL1jygNtPp8QOIEhyYVV4FGaYlW33fEhPxtutZuF+n9tTan8AwdAo1pjFzWjFLq/YvB
lXIf384q5bPIoUZWM8Ih1+wAVW2Gwp/vtu7YOkJbWmzh3TvOLXTM9QbTQSIPrTqVPgVCffY6gFqE
7nfkuc3qqnCQxYZP7eZHuajksFvzsO30XRNek8Ecq/6hXkeuPShLGOqD9TAPFNMSSfXvhesbdaOC
ATTeg8vuVDBQn8FXrK/39ZCyOyUqIaCblFw2R9XAGPeaXIHdI2iNLYzqCpsRAWr2t4KWXf2j6neg
ZQpWTmtFW7VuFSYGTivsB/l3nMEERDvQ8rn0YXHoteoiHBX2G1fnIVuzZJ5a3UGVzowbEyz1czfN
qo1P6C9PScekPe2l5ZAYd0Z152gu2P1EIg0rX1lOW7pjLqOYuJw0n7nx/yWkPmw06xrwb0mE2wJ/
X3BX3AsK6nHSInUlzF13wAAMs1ajjXKSYoxUf6Xk78rkZaAwM6ufXLnStORzXvsFzo14uT9FtqLk
Ahd84x++a5lc0d32vSvFwRQDLkkP7KV/jGIQc4EXzVYMkTVnCxHbCV07ejS1+9SISaR9GnEXMZqE
lyYBr3Ql9k7j29hbHns4tOJ22XhQWKf+PwRJXwwcYRbIIwr4oArTMky4LcGZOQ5bKHltTWpHwn3D
cwWwqN5acvoxVRSXW7fGix0vuvq8QcgEmxaMbLmLWoupGYNXpaGXdknK9ryJdAoZLlrETVstQI/H
zJQHOWesnFmZPT+WWjJcCveSfpENfciIAKHt9OHfIRWdF6znO0fLIJPsh3wc8W59j1j3ZDvtnrq3
ow+g14a2j3ng1ypXJ14Oqame3d0aUfObnK+UI5eAUw4eLdkHTmzHC3X4IAeoXwu+GTCugGqT9IYR
Xrj1dpPjP4KbNIEpViv9TD8+VOaaLZRB4SeUXeTLelhw72Ym2Wfk17BzXTt7XocCnQlJZMCKNkxO
oWXtgaQ/8RBJZitJlQTGRiFAgOx8dDYr5TxjqDeTDly4uIgwqTKibcPoCVsMpE00Nxi5mvDxQjfK
vcyiIpNdbAYJ6SVPsCDip7uRag9zxXTJrL949uDw9rhD0GJOJWnOQMtiocko2jiNUk+QiXvSIU01
u7PH2b5X5VL/LOhMJrE1Ym7yLZEyYHR0uG9ThhkY2i3t0UZ/dcIoBLeXnLPSG6n4726umrxsiraI
rSsbPe9DyPst/KNhKgvLw9QC/e+aQ4wsp28mbIQWSqZdv5d/cdYkqQxMiDF/knWWqDxzEKOqqzUV
JY3YJ0ybAg3shIYAC0TJDqHis5C3em6XCOnq2Jm/V1VRHTUdKvZBeJMP4hwlkhDIOddtjX7AYIr5
1uul+c+re3WQu0GxLt6bpdqiEJHIPT+8rOIKYhQIOt8M93jQfD/oFkwcYILLACc1tjPJw74gbiaW
mbT8d8Iui6s9PyeGFnuehOrotGJfvLl2lnT/2p72cV9SKc8LsPdAdrQW74Epuiafrw7vHVt6nz+H
W+TteI78mJxpYp05Sg/t04HDK7i7oRr3kDOoszXQiJsG02QchGiwFK99jCORFXbQn6y8oUSCV9yz
iYC0zHZzorLDHcW9JNwF/rxc286nmtJQtJxS0U1bvwNIyfS6eSi8F0jXxJ5s4nCk04PyHDc6Eja2
hIY90XGm/tdIGfren3BZqQY+NsDgOs+oNbWNqJEa6WnPhPcpsCtsgFxW4AJuoNpXw1S8MnKjdilh
eDsCZZh70c82mgG7OFREJMW0irssSeRAFJrqHW+JFFBfufGYxX6kWXrfeyMnYjvhyipy4P+799UH
fKfrXjhX2IdLLyl+uAms8jDRMJp0fNI/mkCOqFrXlJfC9V4gP4Z1aYGqz7Wk3Y72WAH0XgXjEe6Q
pcHkPeh8bkpL7Jnt1nbTvRZoTDEJgy/FpmCStKKEeAXI4jmCdz23sxe6B6oEWtDFVjKkJhXPq7NJ
pv9/T8UwralBwS65yDmi8xtjuifyNKNDjAfhDoozkpDcV0oau1czzWv/FtaVtKl/WIC9d+ElXJdQ
w60ogZksG/9GKRgdn2w7lSmJR0eQA1vgc54qD4XmysMqSuTySCLBAbMTupZbE3Hgfh9PtSZPE0Za
gvNpWderZ5JfuHP4Rx+i3iKYOdbzkdhoXgDc1qK9rHJhA/LI745YPb2C4ZnwfLesqOAOMMewx0wI
V2Fi8BWouuIFSYlW5mMQewg2UB31Q2lypgWLZboLVT9FglvepS3PgZkYjCM4Pkf07zqSZotO/Bhs
rRiTXQPSmEfTVGvD0tAegvFA/wNBtnfp8F/ocKlRlqgPZAzktDGXA8jTgnK9Z+WiRp37/8D86l08
O71oPZPnUBon8EsWYPYCuK9nYTAvSA00vIHUOGI3kPb8/pMTDrlRL5WVD9eBLv+VBt+CMRGDty/F
oFQoBa/LT9zFLX/6ZZ4RJDBIjaNj4/+btJXfiubLdnx2wCqX5Uv83bevWZanOmY6tUlqpT0imyse
NGfnAOieCQl7/mGMbZLCIJhUn8fERk/0KGGvUJPmJTUP7r1kfZmu+JORl/IPN8caPGIzTw8OkRGr
zRpyEq3Usgy1uTDKuBsN2NYDjUJyFq/0R58YGs13qnazqNCDODRAzKpyVbcf9sb+I9JJDDfffSYL
/SirEZ1+K2RSMLP7uKKhEVJEMNm0yxojmYQT+BVLrffkh/XoLtSrUX/W5A7tMlYRY38lpakR7fu1
6bEBKK6qJFMa4v9+FbcPtXLWZq0cWzrt/0+0bZdM+5opTgCo/A0fLm3cbhPimLCiCflUrADPPRVK
19QKChC+kyGTf6PU8O5MFjIsZXS8Bb1/FVDz9Wp0xC/U0zD0cPSe79VGdLInC6Ge0mvXWCrBxh+5
HWVDj9qGwnwFlSSGwnGy99+REFIGoVN5bLwrlDEL7XJQXyD/46w+kMcllAscukrEgRtLwSVG6w7C
mf46ObHxB1ZKggPD/xARXoTQthDNf7Xx2crNDjmVqaq9DT7rPxEk0FWHBc7Qon5SyqCkNUF2CxZ/
vGsEi9ITZPXs/CcZiblKiNy0qfE7RWorz/BMebfczXI0vsLArugp7S9IAlfn4gePdZJQmTomAmyp
cS8SAh/Yd7wrb0Qq/2ZctZ1DAd+l9sRQpv+kY7VpvmTjrkmPofrGeZ/oym7PTswgrlPZ2OqGNVnX
u0BqOlemTjdPhWJZskZjesWxdmjcLaKvsOFtIJi/kW4Mgvgle8n+ADPHs5SzHwtPG4VtwiTA9Bvj
TNySNUdX/JyJWfL8NemluwV68XniyNyKS0ds9/nGkZ9hrYHZ0JR0wEeEzu+g/rDEIRixSoItF0QL
cBsN6r1xBJHwXP/VC5eufwY0+OKApjV9k9nSOjC4tMPmyG5wslCM2XzfAaqWs3iOdyh7PCzdBuR+
TyxtvUjgLyBxNDguc43zuSexktbsr9OR1Bm83nU0bdXHLsMhlD79rfxc6IEBy8G3qtqSZA++RCyA
Iza2nS+btfb61oJr2ELroRZH9teM7Opo4zJ4C8NKCP6ERgxsqu1faqTYYi4shnG06+5Kaj6MQpWT
MvugNwdvY3tDq9UN4XJPKr0AgJ2zJdvaKi8+j49IPzSUX6XhVOlMYmX/9L1qP2BBH1hnP6/rsHF4
v9sgDQ0QUGg7eVqzGcdLk9IO/iQ7mt53wFMwy667MAB7duujsfSK2meJ3EyUIf4QWfKoIeedQPW9
s2tnHmuv4AJQheobfFxsI1MPNNr0iqbnJl+VrKqu8IJEES1NOH1Va9klc726XUce1NFs8AjvQ2WG
4EmfZ/fQ7ycW1Oazwuco2WjwieyY0ek09xPRjK2GfxoHVu9/KXcOj4nQ7ltHKrU0Frrsnc3ABo0K
8OM19Ku0UsNzGa037LYUBbQs/hdj5I4LVXKikwJkBfxYQ2MDWyaBqhcQtc4LOQo4MMhETC+K3prJ
ZfD+4BaEVAjszCkNqA/aHIIJurRX3eXzSnVMLLwVx4RdaMG8K+pHF+3yHHm9lRAIfGfCyfBtUnwo
/iyBpHgMn3dpWfTa5L+Qk5CSGQ4ht2GvPe4sPSz6hAREg3SYZD/odpyEnJ3epC6DzSM6BfVa9XOF
ucDaNOePdX7URtBEcF8F+6QqIKyaOnUcQae+zbOTx5R1wmAtprhoqnWS8zt0ZOZ+bqTFJIOEmpVa
yMex81i2znZbZcbCUJXIW7oZjHXpAC3fqTKTD7UbKJSSb+sMu/+TlR5LxKSXKBd71uRC1QMjnQ1o
cCZAgr11whpecL4br4mSFP5I5kjhtlTXjAXo9B21jVFNWLuFhYzn+ps8EUI5ypaEAcMxg98NC271
rNemqMwzhG8IJgVFNRVBHfgVAFjVv1NiCSKmJ12LfmOGMRcqbA+YM06oUJQTjvwugi/FGgndmMYK
8Q9y1d+P7Syx3K6q6dgXZMO0JPA2Pz2hj9sUbmVt1HF9lRqpMBRdiURqKXzhLyrIfTYbzQv0vpvy
UVRQmHuBiPBXaNBS+EwqT8wmGIomUaur17NtF+hAaRV8ZxZcr8PPLJNB2dxCjmm0AapPlkRq3sgO
Y9orlJrTpeb16U4CTsrSJ4mWfSYxO9ROX+mAxD4VhiaZI+pUBcK3eoDtBma75K+Z8MfOI9Cexp/D
I+xY8mHS94b68H2iTfeNXh7/lOUoAwfF+rRX4pGs8YnHhZTocTLgYKywRAB3jrf/IeAgiCGNzsTG
gtHfc9V694G8d0RudhjjpnnmV0PkmkHxMmArtMWaVPNtqVlRKTVHoMUH1m4c4uwfcD/xhUZMaILy
X8/B2m2nch1W1Lzb9z+HV/LUrnqFNJhuJyLCAt4IWWYFPSYcAfJa9025bw/sjeeIE6aLRblyDvSV
ASW86oKjLlZ1/gw/d5N58J7hHA8xBrf1YSBmB7bqRrMAi/FQK+KNouXwPf7OLWHWtCtUIJkAQAkE
oJZL2YSVQjEYLEveKbj45qbyUl0Ht2t/x9OlpZx4Uh43tLAZ3koLqvCwihfDSmbgZTnLfFQpPoe/
0eaySVlHzPRoiRk4Nvjp6pa4aWPt9Yp7NZ0Hya2sZunh1pRjUz2yvnElqxu3yuM9CsmLvUxwMifZ
tURqKYvd0/52gYwzlwNjjIEzVAIXzHRmMh6Lh4FmGhDwr5fVXBRkEc4PubWsQgyi4Ps85yJyb2VA
R6ubsLqrZjQFphAp99/mtrCsVu8ChkHO8E0VrOsKpB+GRmxFN1kQkklVYFIIkyNaSvCfiZhdrGnV
8UOvHCBiD+YrlbE1fOnLIdvf7a7sowjwCnD56dN71YiEU1/U1Zo1v/0pCRJy0l6kNaSUj8tH+U+8
tFbLt/FmAxObHk7V0Xl1+UQB9IRjN/n3HfAS1KWP9muQXMs+4RmXV6WSaKrDyaWod521yvdmHQhD
aV4wRBNDq5H2S4VtinviAiLMxlBq4IRCWR5vI99F2mMQCqcwnXmBAlDifhP0m3no47RG7gzoKlVJ
fSAW1SlsvcKUXCAAIM2rDkqRtt2cUf7vipdfBaYKJRivSEQx0w6ks8mRXJnJ8IDzACfIvCzQWluZ
XA5UlMwI0Hzlun5P3vWvE10P9f3o0VYNT77YErkmBKoqdBz6SyGItugWuBiKhP3Jgh5xUVZj333Z
w673kJ56rEzXLxjvVIx0PfXHcvaNoUlxP+lf+NxVyV+IA3H7fRd9wd1cpwWra4N2Uus1mZ46ikmT
jW5cFmDnat8PJGaHRpSGdeEXoao5EbgVlZl9KQTPYxXnrafpykKnO5z3CwhlWfdgnPUySeDlp0BU
bEG+BK+DovJen8+yXYztkPtS08nZBEZCFHFmB5KPu3gkvVFHpwBxPplJCKRLA+mKak8iwl3vSJci
SGzBqydApbNunHq/E1zPy0yy6ru056r57SiWVr3Np1YsGU9g21VN5q7+coZHi5ea2Y20APqIr6eU
iMpQuXSQ1PjQbYuUKQNTtoHdW+X1BS11lDKYHy0CsMi8AD9jf3VX3dvig90bB9HMiw1GNpeQwb5U
uW0v8wKL0rbLBCcDaMzJGp9I1pRUdwQhnR0rcdInVxyx6XluBZnFRNFw360BwFSgg//z3jeQmlBk
Ei4sFhUrpLXoF5XvswwLGpZW/KdrzYCF99x6dU536XMOiZp4BCXuipBcJpzfpsdizFkTryEZ1jjj
7W5pL0EYur8bmZtX+RHIWWHGBGQefTfB4OJyPbFMNFEbD54KCOe51j9nP4LDOwJFAncwDSMXrajW
Nz3GS2SZAzsuvRz4BgoOpTIRTfibLbdNQsR59Zb8tGVb15SPBAoTFxiKwTOHsSS6i8ilj7NtrGSp
0PjAmr2pQZYg9fgr4x5WAOQ919eXQZvmTAnSjQKpgo6xHMSRfc0faXcs0AT2aCQdpxMXpE9APosJ
19Du5KLmVqfVhY7inGQWidf9BflHIDlN9WJFFl5j64Vec8zs3AFqVVmDCSVatDikre7qOUNFQREW
Jtz1Y45k8PcBtbbYN6MfpC8bSgxVJLGxMKs/FTbwzJ6NZ+VKXyWzkGMQHt1MLcupffVQukommdoO
bC6lMJA5rScpFLk98d09GDzG9gd4KRab6f8vO5XRUfBmwNXdAt84cS0dv+lFLz3cwieWDiA4lCq6
G+jwzFHEPuxYMN9p5EVdE1PK4jnSGcDDQv63AQ5D5ybeKaKjqpW0+Xn/TF6CYBudf42C5yF2Q93M
V92J8q4oVWDFx2eTW9gOF0g/zWCQXaq/S8xq/ljN4nHYNsFFOTZu0tXR9r4gifd54xD3+DEzy8Q/
N+0Hkq4c6nbt9/6HEatam1sntirlz+jI2XrSTmYrX9D7iYXQo4NrFfMIUfN9OlmbTjWGpxps/abC
h0xh6tvTsKmYa60Q6+6VVhADPXB0MrKE60zJP3KKyBcSdWsAXcdDhtCFPuy9tF3vmZXnc9TEoRDe
/z+y7DygOzxW2mODUYLiYIeq+hCrwLBDvrY5r3Gtld0M38kDkJBd4yWiKHQuBnmAvpZdw6nFBexG
lQnwmJ9+SSC4OTeFfCoDdepYE1S2BRiyWIm8v939kjo1Wuw7VgnD1pC2NfiuggMplvZXQWVTHcMG
R6z8TPItP0xQXGZJYFbVrTQUM1MluZ933xxpamzui3GayOnVjnq6Xdjy41YZAgLWmGPM4lffbDNc
1Wu++1gLkcu3N9k7CLTlrR8Iox95k03rj4kpI5KZxKIUTuPYIvG/qqcP9+q/Tr4+FuyerHlyKh3i
W2R4h/7ZdUTq/C+HMt1CPLqkx8UJdKlCrjgt581Wo3wCybbOWKZbN9r+eB+iGvvYB3YN2eLi8ztw
tDKetDON6p1Jjh4UyO2AzNFILWS5Uhe6LTEelgyqUjU7hmxr/vbVTxsGs+JVeT6ZhgEfLZGfbQyI
FREpZk/vcoSdlbJJDr2KCHNReyKrC6w7h1mgCDmB7TggscDNQMeipMl8U0q/QalX0lguCcAbOuX2
3sm1Fbv4DF3UfqynaQqALL4Tq7J/ebwSnpZwRC3ylim/4HGMEZGqZzVmZlfUbcvgeKhNqvwt7ofH
dpw1F5XrHpizcVgVOYiTK+mNFCWk8vMmvGQ/X6tKhA/o4R+o8vtFCwr/3ZxPxWfMuxB96aUUTHpY
4RqLavOc8Xb62f5u6Q1T2Kh78oujTEKx0bVGkSa93T4j+L8QRAWNYPWBG6lxZQP1eB3HJM69PRfN
Kt3wQzAcXM29wWwoiXwvFO3EP+PZkDoMnPnaOuwaQU3bIji7OWudBosnAvNWlLMX3sV+Bv+JCyYN
Ui6jpY4YAZNgoMbF2qqxAiSUgbWf5eTiYRp6Pw7r0XL9V8b99cd9LIpbvRmX/yxVFi9/cLGZ2vyk
1xApSbmJKJRBJRsKWLSZKpNz8a8oWoYlQCP6SUD7kSqJDjCRk3PXeeiTYWEGhY+M/PgM7X9hHkv6
TH034mMzZyqrVdFcHr0fpgL3xA8fP+cJgLiu/xWRdDJlzkMKd0rZjxDWrl6GC8K4aK//krdPSLy6
AujwwxjUI+jlsuOEv1JfpmfR72RerytTimkxLs+pEB+FZoYeYgRN2tsnaruKA7ueIQ4YLTzb8awm
MPKmUFtIv2Lk9yw0+UKcqH+1evrTnBWAb5Mt1KqFirZdf2g6m7vJ81w5teN/dTzpZs7TnEO/qmw3
69BAs+0RNPOkmAyY/HnWa2ZdXRp+ltOfCFw4kN0oCzBd2EdHddRjHXWtsFmuYwD8SCa/dq8OoheP
Nm83GRsLF5Jz0GdzFdj/trtp3MF3TWRob6c/zOsyo+QRMwf+DxK2veLygE45lWIUq2FIX6g7ExLb
vBu3/G71nVB0CtnTX5IOHsOnhEf3KowrLWUi1yNoWbi/V5/CzfW6wgB8vGqj8jm+DLBP1Zp0LE79
MDGSWFrSksoEaWyWlFul7YFPcGydLdNsbIw9lnnIkBgz6JpZbRZuWWJ5rgYUgJa9j8O5pLov8/xE
1cuDiNF8Pn4xTIc4f0dUzLBtF5kS3uWgpqcAUWp/VWY+P4Gvfl98zd1FNj9+UrUweqAu40okBBMS
l5oQGoWmoD31S0RstBEaAIbLOq2eGPyevlI0oK7nPPzr8P8ShGaOtRdZ8gQEAk9LMkXbl34YA9vS
XWUP4Jw3CrIIClKfNdvWO2u5Ea6dtNtXDKnqCK7sS8WLhzLcpWSYu1qahVAg6g0wzXqY3uBotCVS
3Rmylp4usfu24GTg5AfOwrqU+v7EA//l8a5Noupa+N/hMUSX+nDgTXWQoh5bD0fWnvHGyI+Fszz6
LAuf8WpDLgAPaji7Xu6cFXEwFQ5lXFBC6ZEhTSELDBie5z8HdoNmECpeun0/5Z11YhWWT5X7z5hl
uS0TmaBMbpfs6fwv1jg+38z4z97mqeOd+23siwHMYGEFmpHHIOkpyBzdQKcHw8ygSVtT1c/2k9Vk
RHm+hsETZc1X3kg4VY3jK4NxRM1FC595pqBbVH40IUSD5zZ1FfVBusbbdu7j1z6PYboxoMyBICm6
/6Z6GTH3fqNmUHSxz2nhN5a4t+Bj1bI11km8kGXiTYHudKA+z8eyJuTwjPEH5V4DQKZfiZpZZXPc
/aOsz6CkSKjRURRbhyBej+32uxDK3cBlRznfaj8KI9pW4CDBixv4LRlrB+Mgot3f/2r9aGvEUP7z
1FbaufMAfMGNtuOFXfASFB7CvFTDCTzBOeSXdMpGjdVBu4S7Z29AL2jH/48MyF65VqHt1IMZxSbd
dpsVEoAHn+iK4/hIHWA8eqOTWZGAABsalzcgw+Q8962db1HSrvYqYGiSTzuIFSBpWneqjvGwg4iK
GHJIa8arf4UT+kqg2yeP6zqt32hyjzayBpMWAZRZYXp8GX/3838bTEeDtvEg9o0uWd7OD3EIBYDl
VA/DvILWmDK+M3lyTHhdB4u1IYErZ2YbmhE+73GBy54V7b5KYoOF+Ut8z0kHKUuE+xaUEzk/r2jd
bElRcLbg2ZSx0+xreQMgAKZ+6GKqs9xJMqj6Mb2z1jYd7B8QtcBjnCRYiBBncYtBvMmKfMNgA2R5
obCBnQMgQrNN02NglHx3wW9NDPm+jknFdAQTPAmnW1zX2WtN+inAmkDHT79XNaClBBTVbuqe2YDP
fbXhMyYyFeVW0lkhyNXlXAhpTGHHiKm4OEKxdDYZTTkaEiW9lbkIfWLdz12rIg0MFYDJXLXXC6D6
uOmHSkqMqBTemjiT/zbNnNnMDLA7MudLSvPtfMyCXhTMtmTwfWBAGufyeyBmLcdNNoxF1sKmJEBZ
YN3goC3NE+tFJwNk639dP/47k9EBf1r2K/gep6baxpJb/MS3sbR3EBVNCI/4/ZBwiztYu07t/tMm
jLZt6taHWbfhuXw6yCKk3h7nk9wCrhj/5oPl+OTpxacs4yufDNwaDl87Vcgm18heRsNwKLYbnTS/
cgG15XPocRC/trwDZ42aHYPbLT8YAd3X0+mjRLVvErGQrMT3pmAK0ottUWRSLNNR0djdhGUfVPs3
rws6gnMacJCNPITYveF+XTKYpah5Xj86FZQOy4bdvExBCN82fWbznwElFKxapsAg/D99lYQxa9Nb
J81Ko1CRE5oo8xIzCXIo+8X0RmS7YnXZkz68ygRTmOF0ptc6WuRLbI/TMPCnDaMUZLcpHrSW++AB
WMNcm1LIAV6MnhudEYp5qGn6mIgozuWVJg1ekk5sk+vdfIIa+BgWdkYb77ztUqwCyjCYaBPjG4sc
kv+2qA8rNpllOiqOSrGgAQKjd6Dg4bNdq3rZMjZKBpL9MkeyDXnaJWs9E/ArwKGu+d3JT3gp7NJ8
6knBS6fsKpC4tXDqpn49YwRvtiYqoQ9yskzmuC4b+OtdAjUNzeXoHeiAaAy6lReg0XWQScGDdbJu
uBawfhH3UDR7qPKmgJNnJINPT1L/YjdTLKalAZmaYnNKM5Aluj9hujOiLRLaCLtH1sgVi4QNJ+VD
QP2Gwr4glb6z5X//CnexCBOzo/bc/+JmqhLLY3Wgdj+XlocUgCeIod6lwat2Nmm66i2MIt83iyK3
5l2srHPF/Pe2V/L8oQO6Mo7ZeVLkM55028MnjySfikQgNldQg5zP9C/mT5vrj2AOmoCwY58C2Lnt
kKdTL3/mr7jipgEb0E8+N6Yo0rd30CjiagiMF4ZxvI9PisMq9L3217v1dVyFSikuL54HBFcjKOvj
Tpz5+mNLvBATEuvIq2MJr5QPYWpgLYiGZ7xk/cg8Dv1P0itieKs6wYqEP+q5c6zjLTag9KOIbZLw
x4GQrIlgmBM23lYOGTqAJYOEP85i2WctQ8fwGYLfjmGJEQ9QqVB+itjPdIslJiwtQ70a+QfG/yIw
hQBxivc+o7m6BOtUMOkF+tGpD3FqD/mk9IYFeojAsKYjmk87pwhrcGfl4TVG5rCBQJM9hCdqpoVW
DBJWyzTMGQ8PB2pwW6dWM5v//ZskcCRVK74cqM8vg8rXi1JKJRqWqXnPvftwyjRH/7cLlc0WE7m8
pxWla2J8JLH5Kcex+VS0pFGA82WtpysH3IGKx+Q0NHD0921VeZkJjjHYUbxNoat2ju5u86FPQQIE
8mWf0boPno24ju/HQildoq5Cgbstn4OvUH0hxWGbwodJPsVDJNk7i182wJIZSsIKf/jO+Stc4Vp4
QCY8vp2zHSflgI9XZqx88vFne1rp6I0RzMUHPaMiZIAsHdlGNlVHalykytlQmJw2kqWrGpMh38U+
VDnXrShNYovuU0oA1rvYhmhJok7A+JaHjGOrgWcs1MWATUjiO5vgbolntVxXJBoWJqW6G9rQIA+Z
SYGybdVSY0441HyYfoMN2iEk82tPraBCVitzPhkECOQKHgci1YW3g528aGnkP3h8WJNCfp7inI0B
TZBAL5ZvT0ruAGSAQVgtzXT80HFcwnR+RHmjvTD4RKsXXxU4Ji+MJBX/zKc5Id9p1938c0Q2eZcs
WtQxjmYy6uVwviNcKzKDnKlZ42Jod+bvjl+W1clw4ExqvJz3+WkWV0CJ7gyZFrO8npGvW4OTeWYK
5kxFf0QoI+VjU72BWT1hhPvtiMPjG5UxVUuJRAUyJ6qC1OFlhHg1N8GRSiHs5M9+HRR4Ka5cKqgM
Z/mDmmFr6jC/ULb0IZLFCn6Isk2J8erHGkx3aiS+iQH9ZcDRsMNqZzLlAUiHLgVSgv2TLMK6VIFX
UQB9K4QK7l23IzvmJ/yLuJFRPo/jG+wSFu92kXDCrEz3AQNG+JC/ZONn9c/A0oAIs20E+2W+tbAJ
C9hs25BcO8rw/GXiRcY+jKQjmU4JwoE4so+dm7rQie/8si+ALg+tgr0YPUowQXFMzny8d2KDbxQv
fLprocnwoXH38jo6UeKPWp7SefaW4SFzSdac7yyqlhhM+0JVzHyFBhiTR1plU32VDTj2oH9Dev4r
kgZPms9rZsCm2++OGqpNr3wQsfK451Uv3h2A99lUfZAd3RKEuRxAa9O6OK/hgMPQYkAPWvabbZoT
4JTdi2NReysPxSuEx5e0FpHuY/Qe6G5eLiS9oPC7h6XJCjJLSYfwQGItCYu51psKybyCulTG6z/w
/Ym22f68dDUvd1ORhRgCezrc3HnYZNc1GbtEh27QiEyD0R8nozAqCsZv/Xwoq56d+nxWVKSgwPUk
1X3GBMxjUdgzb9Kaogo2BovEdxaugsYH9wOGZVYgONfsDiNaq1jrI9ieAPL10Zi4HJXmKDmYYEsk
u2PHCeeZL9FATe6jLeSSpyldX7lKLe7EkLBj2cbheZ1I4BVB7QcWkjXg1m3rdjXpt5LktbGwpl6i
gyJEJbW35MIxJ76GtJaIq4HenzcAcA8JttOEMIGe8VWN61KOlBPExpFPg9O9steC2eLBE8mndHIX
xSUppD87i5V0RXl1yNRy18IeHs8eUL8pigsM7knK9FNi/oi02uZ5EPllbZSjW1Kjv2jCJ7THJ7ax
9JQoWhyJ5o7FnjI7h2NJnJP3316lPWjEYrWdBBrNqtiuSjIBy2KV0wmJ82s6sVe5EobH6FvbzgxM
AEwsJ4dFuYGE+G9qhVD3u77h7q2GtAv3EiheXSXZvMVWFafxfbssGTcYUJFPb8XjUqafqYeJ/EFI
KIgaUDoHivG1KXjxSUbCVpfXuJBceAen4Z9k0x+LM0qA2GZwNacd7sMdux0fbCe679j5HOb0dJZH
uTJqsT7RQckl6APK6F68DtJiMYvQqyh9mJHyzWDqwCZKEzUx+/lUvAINQ2IhW8HXDW7OFFwkm+zZ
cl2j2VQGbgCxsqutxB03e9FLhaBYHqCdFeVnw2b3lwNQtR4Jk2j5nt+qa4x0HZ0COzRa+0u8TmIy
lGzq6gvQqAUJk5PNMqLOiA1migs2EaE1fI6jCp9OiY3nuGOPEQuK2dhxEE1bw2XnL7Js//XLdjtg
kT6jzAbrIZvt4qVHspgo3ACnnvrrp1ubfqgCSUNPaYgUV0W3wsRBmBtBpNPvHRRWvbBMEOs6l6XI
IBbc6DP0AUpPRVtcapmIhtpieOwTDOsDaqQcbJ+ZF9aE8snpmxR3uB+AqNVBxB4S7ucTs1wV2LkW
ySrnkDv1rd8ho0j3UVTcDZi7A/qpdoN2lG/GYYj9rUS/oazFJRCj+eyIANY7G7m5B26oHzYczGNw
iwafhiRNmgqODetHE/DdrtZD1R4AYOAeEurVSir9HPLJrZsYmnTgoHnhKrGln/BWxlLPeh7vtF5r
7j+i/O1gMCmhS2Ip0cVZotSBIyHyZoHN8czsZ+lNn2L6vB9oo0dGqBsoc3dDrN2aoTzPlmjWAexw
EB5Uuw4NVuDdi/fLi7ZkU2HPRzd0bdtZYss859i2z07YFD7k6ohlFiLXws8bjIb3wvGuK355LIyY
yKobZxKlb2K6Hh+1zpMsuMoN8n0I5uxsvg0nDxhcJSTHHGaalhhhqVPFs8IYMM6eNW0JX/bI73us
q1Ifti92ltZKfhxgayco6jpKQ2M/ks/HnTL6XOC8KIBtZI8sTlTN+w/BpwLfn88GXtoneoBzdhoj
cK7yRM6IuGENs0QkQebdlCT/CF5Pb8F/OFFBXnr7DRh4+wC6Of7mN170h/ZyAsLwEL+XGjdBjJTz
qtZdOPztq6lJ1cmGxjglJ91uMVJDrd1mX2s2i29CAx33sUPdbWtaeuhJhXOG53MxPWymuJqw5BKv
mxQ6daNPZ7WCk33XDSGV/Kt8QKrbHLnYHmE0PSlgfAHyTtji4BfEcPQuI8JchUAQztc8fWSaWkjV
nX4Pw57QSvRZ02nTzF8ArNsAo7ERT+x/h1irZdYVkTDEFCoY5tFTCHzY5w0RDK2lnFX6lIiG890x
JMlQR9KR6f/iUeBddv4v0qGQtPof2dLMx0+Y05Uws20DFyQZWCf7qQKGvFR7Qb1mVfx5v+aAQXlw
SJCjeMonKBetQPgglrsueOZnTDx92c2p5UDO8lAF5Bb9ZhpvGvEUXKnDqWOOJjehzj9rI9REaY0l
O5ByGtuHsN9M5XFiogcrAx9pmEy4gkSgKlscZH4+cJooNTrrKIRLhCo0MgEZczUj8igYhcc/q7N6
b1N/OrgoZLssxyUdCaG9QpxpCKAMuF8ANPVfoR5UTvAR5Infhuutvpg9hFKxIM0g93eRjN8DAcTL
HG1L3ofoeLzGhcant/4jVJ/iOXkaU+hYeoWE50qjsnqcqKOYfxD/xytOboVBnjcincPjqn6AWJAt
UfNOqwBFtZsrKD+sVbOBVqcDq/w+zghVpxjKApWUYuGzz5J8DyRp38Fxa6ZoJ320YWh74jPcX87y
c44MfiiDdN6cniv3O6zw2WmNBePO0e0Wq2trHwcyBi5OTWVG1yHEOcpEFWOP+VsTTvGfTPwoeyk+
Nn+bxrfrY+Hl8IRF2jG33nqNCiB8HH4eUJOgCjs/YDCYt/dZh09ysOqz9znvCNPaVz1XukLDIm75
ufYSsMj5zoqPfhn/drtzAt6EmCMGFUrvt1qq2LTXeLmmcwWzOY/Ob5ClHBEQyJvwAowCYyA7Cahg
FGRGzEQ8n4WnKirGQh/XJaVa6oxeNhCX5hKU+sW1UbLQ0bEqRkk3SBbYKeSdtObD0fJLRDzv45Ea
VDTzrMnw7tI1UYIjAn/usS3IVjM5wOjmh2NQB4NQN6emmlmVVjJqN+rmD3GsTHaooR0a9uqE+w52
Dc3JFPxCHn5CtSzp/E73tDUO90sRIEtXi97iOJhCVCl/f7BAEN/OdRJuNtHOLXQpBZa/GmJ6hLwK
Efjuf1mdEECEKBVOjLZWWc9Sk2FD3rA1LEGmiWZ9flk+lABmq85ymdIBvn76lyCeWnNRHwhl/Jla
oaSYT8CPw4ASbA3kmEU7pxVbdA6HU2iURbVhzBUEoQ+aZwrbDkeo5fvMWZAGXBGk6Gm6eVXgj8Zq
VmsB+P3h408O/8joOrklEEx2DbaLpcDN7VUZ81W5YRWs4V/3HwNkQw8PGGpa93kNBaB6ZukLhEYQ
X9U848ldYJSnK7Hk4vhc84pMvaJWhieQ8E2t/N5U8buCLgCt1pIiY80+yRpeuYSbW7g6pxFbSdWk
TZwc5NRszIX0GMAJA09Ciima12Ys3qubaJSk+bR790Dutg0dC9uM9G6rFYu0Pue5xvojr3gGH/Vb
UJDCZsE1NYtApY43yEre1jLNPLaOHM2A0kjyCe5iQbVFpZWzXgXryS6TCdY609kbTcUg6V9oiZ5S
RKyZxThU6DmBrU8n2XB2LerQrZOBPAQPHrmxai+C9OOOe5YLZDjKQGLRE2GugrNdk/fFwTNN9bNL
SBEziDFl34eyXXwg/1gCaKIVwS/tIRZhUqxkQcir108G9EvfV9RIL427kCiPAwKFn5IDpJ6Ksr2G
WwhXNubXKodii2PSuY3IZj8KDZwj/3fG/VyR1xHzL6ycfs0RVXqahsA3h0diUaRJ7dFs59sfjEoM
y9PaKCY64Ta49C+ae6hbwSHGAuGSfh7fSpJPTzmOPhgiS4LH4Y8ibGLp5OKfqfPwKjn97zuWZ8MH
SCDHc0VuKd+OJCuKuMJUBkmBU/laFJRpLLlmUTSUjmcG7m7dSR2vPJ9JK5+1QI9mEe/N3XcQuUow
WdyLXnLATbDEDBRDHImU1w+gxCIgQoYCMDYi46KW6zJdCyZ3Zr4UrfrxJyXjTi0X+00i5GS/ZHbp
4jgyT+5sE7XLwYrUANpsw6rNult6SxzJ1fyqcAU9AMbnAFzdTDkv0EbjRldKyYjMDnZMwKuKV1H4
+FlQfLZ9G9Ug1O1h/Gl3tkUX2yWDfdR6AZ4O1hoHDRfq7HrChL1wOM3mkUwDxY5tvzdcnKnQyhyg
fC5KNhP89e6iIgLRIT+1zORcRcnRTbOIW5AObrzNrMdl9WopD4NmlwLD3GD9IV7JrHx6sRj0HB3J
5OdrC0Ucd0ihRikKfOrdvog8lwTekB3y77XbgEs5IhlGCU7ClgZW2lzo5tmpObbcIPT9qSgSBV+c
Mj3ESR/NSYhD5OcqjJwWReNsnFEPIHy6Wg3FZluC/YWsiOGfidoyh2GSBwsKtGyvrr7quIBw+gjS
RWNhuE1udhAUZY+3XC2pOSnmBZUJNUrXiZJt/D1ALf54iCcY9qCIU+SmdDMlwlVqu5TkhgIqoBEx
OorgWivLgwBGB67vwA1oLC5CfXgno8PcO0JtYkYCf1eIoPl844DLoo8p76P3SAwf56f2EkrmhraF
InutMT2j1CjXiGA8Y/4yBKzLlSZ72bf/Nn3b9s1JeVXNqFrzPAZBUr05TqPY8ltDDmb4pgKLf78Q
nn6dyz47GyZdMXTTqamXDmIm4xdCtSZp1Y2VWZUXuQT1OhL4SgqP9GcuSURaNnRcpdsxFtqaYrVu
cWwxnP3hodpWHgs3D1LT9CV5g/cztvbJ5VZ+G6PGXh1Js70hk7xNTTNnwiVN/WYNWNOUTID3sTfb
UUBKXLN7Vw2oPDRqJQ8qNxvSUiWbCLw7jidsZAkog4iLRDzC1OlvmZ46fv3W6qN0nH8PsYbQBzuh
NHuXrpt3xj6Ig+mkM093rkl7H3qzObEfvz9mG9K8qp5m/1kF5JSyueoIzXRbCU6SWdXres4pjcTN
XoncPKiHZT+QJsgzp6qQusbZKYdQD5jbSePjDpHlcHPS79OSx2a+1fQFMfxD29q8Emdhd4vbwmWu
JeLeVABeQ9AHUO+EQ/8+1OUHL/8KrHbHlOtW60iuPXlqC+mvuNdjsVg30QShBGMKnCxacT8XBgOi
uG9205i7wx4HwRRpfDIQq7zEkxbxqJ6ieRlqzkPkeINtR4urXqNrTHkhomOPBk9+ncWFe9J1EOxt
DLbwXbgNiEiWSv+HT+IEA/G/lIIOO0bH55O3kiKrzMYu4wtpJAmxdmUXfHolLVqphbRcoVakGMcI
KctzNfcrCdoo8cBJUJdJYh95wWy742QjZpiy9K6cCXXSoMb7OPtTXg0pP0igM6d+97UWCZvuJmdL
KGRwGsWcTU4xcfERiMZmg2YVbywLVR26hRxtrVJrabUeNG55Ljq6kSwwBml0qd//X+Fp9sUajcuz
UCFy+c89c6CgOrdbZpDTSh93Tg3iE3gvv3WLdJa6hx7cl8ez+BTvW2rvtGysMhVeZXfAHV+g2Nix
1/ljzE+m2PHEgYcv3FlliExRqLR5sLSuxCPCD7F+Zgj6FhCiTaSZdWG9SDESAM0Y7qesgZnHx6iL
jusNNrwEylumSCn1n3j2JxsTJ9qquAo1nIAo/tZ1Nm8vr4MxVP+6Wy3UYTk/Bl5oJURIZJbtAGe7
KfvptUe5L0ND0QhTPyTcB2QQT3GxPQ3w+Z/Q72KRKf0HmtTy38a6YoBDFa6dBsZ93r+A+pjRzLyZ
yDgE5Qkxg20aJtnfISJTszGxwyMqC4uvhym0+px+jOeLbXqlB/irONOyyulatcfm36LfGlISQVy3
eFxGH2F6+FTSgpHHT9mY9L7vS/GsaTtXgm68QrY2mhiThcn77lFAWYxIXiFD0ew5A+9WyBpLQeDe
ssgv2G/SI+zex14AkhOvieZQOlEspVKZU4S4WasRqJhv+l550x/E4FuQAVPJPcQXudyDrqYvEEjc
q9jMMwREBIOVwoR1E0ARAyD5ydUJmMn0A+tMWrtLkJ/2Dh/9xOIFkfiuodJZpH0kGkdox8zbW8iE
At36m4YJQXkhg3vxECACiPu/P62g6TMPZpqwTRmCWO5L4cecHWVzrKbMQ8HScpVre0svPlKukMMF
XPQ3cWQb7EsDO+4lyjb5CUygIj/GIYZYS+sluLgqu7qLMEFTu2k5kZIAz6lBnyvdaHicyYR827DB
KqEHTNRiJ9tJYotb767rTHRFOAUQwntJZ4xO/+luGKCN8SqocaBgORBoha18MRqkD4a5FuXOXmtc
UpBn13r3rFupyJyh3letPWlyP3HV3yrQ3jWki+ajh0sa3AJ4adRYsTP7b9a57BZX3bjSlR2Kaff7
BpFjX3wDespU2vTG7jr4KYO1X9Sg7MGLzaBRmihLtw9B1DM2TXO8PNF3ivkW3R4vZ9E6brLszSZe
5FMcHlD6HSTeIjKjlTZdmlbrSIAyGN19SAOXsC6CMWXBRCtH2Cx+qK1Ioe8b4eo36Ug12V1IV4il
DwIb5ztqmuED7kwjvCRLtkBaUJbtoans6kpG33wengXDXbTlyD4irJqoyWNWU8ZYlLj/4YAaU2t4
Zxfc5HDm7AVT/k3JIbD3FI/e3OeyHmjgUYGkA0j1/BzlTrgYbMtqwfPVn5ct6APIQFmmUHaJkbiF
kaYA6V8rJE0/wreFXtLvGEOfAKfoUFSSzbiic6WzrNXIHo0/nXlzRCcdspUK7kuBzU2OEa5hPveu
b7HPKss5GbQgZnF0CRj/K3I+H9EVnWaYbSaSsD9sTQUQ2wRriVx1ikKM0XXqgOthxycTusIrtn+k
NBuZcLkOVx4A8LASjY7ibVYzlARsOHVnf10Q5HjCGd2xdYqx2Uq7XB1m4zvZzvuE5j0+A2ryqwqJ
ZpDgiqTuIQg4vcAZdKsgDa3zhmEZSLripl5Oj8+4eh9EBuqd69vwoo3uXwgdo8FdU6g4PD8elhXD
WR1iJEnHpgqaP/hEcdAfy7hNpxKTIm61qb5xRIjEse2faoIqSXYW042CmsCE6uw85dqW8EmtyNWG
ws/g/yUPo1VfBrOWWhN9wI4l496RcLMEoiPObqRL60lnXCA2L6NqAnEpyHf2igDpY3K8bvm/Qe4i
ARuRCeJDErceo16rSAz6BW6cCCqbnrtU8Dj+c5nq8yyJo+1i6rK2iPkqNerAPxx6vpLhoVlGHph1
c3lwg3u9css3XnZSgB4XsNfICuzdSUfkqge/8KdHyT9R3kb952Hy9fCMBm7PG87msL7uytmHPHF0
T3wez86I411nOrF6p0K8Qx3RBgT748aQedNFVwpROCYuHxWsHAeYxgSKNAiN2wWqdgnahrhmqKbK
ozJA444C2HLd8FOYxB6dxwjoupyxmexN9/zNBHjYb64hULyZ3uEfBeSPaGufOjT77ktyoXmqSUqH
e1ya2IA8yt9GdnusUO0BR+SSeVFiY4c8J07H16tbb0q6eMfkEAxgJlU7Zee3gIv4pRSOwi7aRgVx
SHjXOsWQOK9dAyu+8OhXcga0zYMsMUZdhVaenrroeTYg8UtUg+ulML8kvO+PkMdenRszX6aKjr5/
VfMVoMFwSN4QQq3e3h5aOvl1mZvkLzKUSwsKgQesvDKahq61vMgV92YVQnoUYncKxQgcqg4Gk3/G
4zHqaxJOZUst9Rmt3NQYi4LbYo1lMB1EL8s7LuBaOSGopQSLqdKJl6A1BLcDTMoAOZ9UNeF22tqR
1S9HCCKwtyQZM8iBZxWpKP+yDh7+JS9ShWUD7hqHml4FoVUdBFOu6IvHgdDPitPN+ypib5jcXRxm
6mu8BWukgUObzDzcDBoBEcH7qtonHHz8c7XF+HXGb3keBsKzQSnxHtq8E1N5GdyPNZIZogy8wyaU
8z9hCgkVBIqRO8xsZO8IeFpXI2/e+YysC8TxMsBEvQXQFXSHcnYvF/ZHjlZLYadSPwGIm0u13kff
FYLgwJdm+ujdb/f9pJeV1WmBHxzAejbJ+wnI2OeiILpYcPi1OKUk5CHmTORqoXKl0IaM9D2xWdNn
k0DnwqExH7Yr8mHTQ9JRCtnMABsZwwTKpg6UPEf5fy9QIxKqCc8MoiucyyFUF2ZSKEH6n8vdO20W
pPvDGo90WNkCyDW1GDR7ThyxhAzeD7/PjP3dvDVO/XDl+iO4wylCedEqoszBvItVaPDYldT+Ih+6
0KXF13R1naesuKejLbl508igXmf3ZPRYhkBM3jlwOBp0NXWSDy0Ky9vBmBRLFddt+ndhqm22hEmg
rO4gAsh8yO2tRItLtmh/m9gZ18j3CuOjOjE2l5P7RZb+D2w8suMIj9imm+YoULUsAeyrMc6ZKICL
1nDu3UMEiFsxCd3I9gfmVOEJUW44iTq6ew9jg9JSw/DPywJNDJoudmkRS64XkLfDP31scX2Oopdu
cuGP20x/AaqXkzo1xJiTVzJXB7rjZH0lvMP59xPT51UmgADv9ncaALE/WBuNnvPlnSwagqXCY+ar
SA8O+W8XNudOFOj8CDK2JlfkWYVB6fxQHRoyS+L9yW+/6giYpIkpRBzFCHFvmha3llR55G3fGaPG
eJiZUIwRafnvoz/OSsXaGr+xa3wHYCE6qCC7dJxt/3E7Uqp8tX08BBeIYsFYqjQZ99WtbI5AOdHE
x1hC89M9goSFnN4r4yHjdM5aLlDLfCU1invG7ZQ2DZo3t7N6j9cbbeJPbu4nR/hDysUbJ5ttKZY2
liNPXDLUvTVzFpfuOASYf3WRGPdVEJkXB0LCdUADR+5DFi2qX0iHDTcHkcnn7il8fLzuSPTeOP+f
7gsKy4MRCepcHAUIdV42yyDLLaEfORD0xrhLq2LY9zuZzzK6nFVA/QY0IARSwFmvlmnqBDm02bvL
/cWEaum7NxbIzs7CPrmVJpTOJQfCRLFTniLxbEf0acVED6dHZzenhNL36cT1jGPf+9Soc2fkgfSX
z0u32SIOCDjJB8DCq1RpdYlWJZS03TrhcH0I5RX9hiRNsw09G3T1PmcSy1ubU8ojZ9SYYA/RiWWR
7C1HPDPwl5VrWE6dt/Ar1ipB+2viphrveNczPu6JewIBf3hDSofJq6OQ8/wzdIuq19FsUnqCIHRS
f58hsdAIePzZP1reine13NzA4lBD+ScZRMFHgol+nQsLn5j62Hu2SjTNrwZcJVUtDf02FYVrBeQQ
sogvjYMy0HHRDHYYEq/uRmGjnqtnVCSQ7RqMYJf3cClxtfpqtRKjKzVV2R6M14Sn7XbiXyCMpuzC
9y89NNztQ9OxS/RCZ22BVXqlj7/bRFkN2LAMsJZvdrwWZQ7QNQa9pwCG8SeIIhokcBqZJ2sFIO3Q
oPyEoPYIlZXHo/CpoNndR+rVhr4Jmg9zdyQx4Al2F3d7k3VAdKdRJU4roqD7VOb9ezCbnOocegQw
YoxdFOKXcqDgNegUCb2t2eksX0CCANkKKy3/wnR33s+dO/mKkIzddn+wKm0/sDKBtGR23xBtw16G
NAN/MWXLrExvTNeC23DhZ9dmnRe0oDGxZz5yb0CvpPbKNTK755hI61jaHdfhI1YD97Ai8qPg5K6w
ITGTCmw6CaYANerN2UO+m+PXXB7MeElR73RK2tuR3byKVCB4NQw7SEO/zi3ebLI8gdfkWcu1Bcq+
4R2vXYPU5iIKqO+poUVz9juQXTK2WR1Q4DJDoQlvrMuIu6O8fIRa35O9RRv5JKjcukO1U3dgr/LY
yQ9DHQWUFx4F9M40zZD9WMT7Y6MP666HfitfNcDLvGbeovdQ/Ho4Ii18IksEorgMQJW9XlTQhJw1
hnsfsUVio0+KYUEkUHk4msHaGQGxf2GCrKwfM0ORa7rn+s1EpTkznsWgO1NjXH0Pd0DTs55S9AI3
v7wLVKmJ1vJcsro+kEWlBDhunxQ73PjZzbez7iY8jd833NDH60niWdGOrfg+9x3IlOgx2RbacqGA
vMlxgGaHTqFSrDQJyPROy+BRZ97xW7UdkMnf9/Vsq4jzoQXnnIZfW9wCUsaJYUUPd4yyggDShpBw
7Z0hl65QMZ9wsTJOq7pjj2poRv242CE+guhk5qABjnacyDGO8f1c0apRlTbuUxV7XhG24wL4Aw/y
S5lx+41omGXDOkf8x+OZ58QyN1F6e1mmVhup5Zw73OfA2qLY3RyPLAbGl4qt6Bem7caXxjvqlnkY
kDG+OA0hkaWcXxNhbDa+SV6mGWJBihQKQi/gV66/wSYhUcCz9FOf57cP4Kyd0+8JroBchbZBvUVI
nBEPl/dom11lqXW6OeEvZTzJAQbKZ4HCqcoJ6uemM22AlVbQNwzuqL0YrW1os9QKgP/z5U90pXLm
R6IiOPbY6OKnwkpoteef0DjFaZu2NR12urWnnMhUb0FBcSIMwZB26yTc0O73V/RJ66+ySrgfVJjt
UF7UaW6qpeAP1hWEITdwFAtWxnTCAs3q2Lt1McjT9XybdBvW86WXhNp4G+uSAqghlxoDbk42PEQb
yk98HpnmrTBppdqbffFO9hImEtjW9yKIucBx2eINk2xSJeKiW/gPZGbH9U+1pd8YQUoe/nC7TVUu
2DBh6WJQtYoEw7KGkgNX51cBXUcTPixPrst+FiFB1NBiuOmmvx9FyeoE1QCIx3lMJNRl+OpgyIU9
vXwe/fSeMfRGAafH73wFIujkdJkek7eICu9PVpHO7aW5GdJqxBLB+zph3+qpBdgY6+04iJAHu3Lz
mjNYed5BUCPa6QZCI1HMoN2yea0Xq8LO5qlCPw0QP8sJbK+ToerhMh46c/w2pgPAoUiQDLFpoyF8
45VJYKjmg6o7K2AWR/qxWhr1GLem63yP2KuIMVnqQU3SxsTbeja8GzdDPGtgH5Y+Pmv7NWGYlqx4
awk2xTGfEX2PS89+esz1LP5bvQiPkMBBWSxVWq+dPkJzfkjlbJLPOf1S76HPJ1pGn1qISINE4q50
L+vGztDg2/DbtjdIPY187hiN9d6wBlhtj+yn3jP3NqBQtXIdMuP0pMqPLNGRZC8iWOOcn8HkB60l
7vgZLA2WG+YtH3GoqUN1fSUqCkjI8d7I9x9lUS0X+N2o6xCfEPAXncYPgvCno4G4Qa3fzxf2sPgz
d7XL4rfSprruP91OMVCvWxHQZFziLBIY6RzPBzEA5qtmqySbt74i0QmsTA2dyy/nZU+3dkXsiUye
TORY5oy6F2eS6ZkZNCYCgWxzcl63p0IsBA9rpj95Zuk+jiuVq/rliNbq7zExIwdSnVUmZ7nivn1b
jOpYi4yuKtD6ZVz7qJJOI7n7SKqhsuACrflxOo72j5qXVCItnv0/545CDXS1Yfu9o8/UPGvbwNwq
rVvV4565IOvJlEcp7AKJNSWtrj01CGhm+QPrsVX2AE+nX2QIPPGmhX5pCajh0587GRPAdEeovYtS
bMZYZlFmVNA++4jmJVP7wbFbW+fIQxVjVlLTycRnTfRlAwdS+G0kkxAt5JhA/83dHohjnzxoU7/p
eqVqGV/NojaDCq1XU4gulu9fVc2rnwHuZThHgLQYBGswYf4Gdy/+SqKENfyhnntzAOJcFniYj+hC
knTc2nflYq57FdTOEPlkxx94AUhR1zHPriZkGCxgTK/g2ijXkfnZQPibyT6IRpTb4nXWll/omcqP
JibOAutyv/yWQuzMOLjPegaqmDUqWN3CbxrZQNhlEdcVz1rnIj/hAPl/k1T6qYVOV1iJIFm4TMel
Z8WNYoySBDZO2cnP+1a8LpMwml4T4GaWR7B+t1fvf4usoxaAsDskJjHH83jZydGkAXiJjwwE2xo/
p+XuuyUhGY/VKeDul7nrreqkTY0VsdkYRmaaLn7ZvYwEKaAnOnjM2I8QCDEplSwS3Ildg0/VhU+h
qvjE+MRbqRMQ6USf8mkxw7I2ipw4i2sm4eapgxlC2pn7BiJ4tt06cwgkvXZVivyndGKADjfS+FQu
HGvSlVbaZbKF2pU7nGQN51T/BDIAnprmCXgPmDbx2TmNqgs4VStuwgOWyvNp4cHw59BupPXGaKqi
YN4o/K6aMQ1TO8Okv/8lXgx/Uuug8YDxVQC6rericQwWUVo/lXF1RME2LrjvD5eVWWnzh9he10m6
Z+bh4IMUZDYHgVPhgjM+Qw2zf9G0ROcDAXTQskRkrkSdBnkbRoVK1UELHuzr7BpQB+pu/kduQfIN
OSYobJaCOkkbVqE8i5L26sLiOZr3utAOFD9LUKoVxIY/3t8lEglyaAA+foNfsBHfYTaK6KZg7Rw6
Cv1OqT1ouuxwFp66WNh85/DDpkp5N/K46nkzGwjkzjQoU4sm1z9SKGhhsgbUIgEO/h0EMA5TntyG
+o+J9OiPODOScLNCvRM3toQpq/FaNXti/DN9Ou+FNuc6Zd2juXmIzQ5GroxQETsSz/4p7su3TRPV
mBFlLDXvc5dKWLbCjn8Ksz7qRnzluBmpD8xDaA96Oksre4FrFMT1cCd0mbmG/GsTjZKVJC7GugjK
PLTZtFHI3QIXf/2divPA3dpC31Oqs7Ki7DUAhXpnFnPvq+0W6vJkzaN+bRX9mh0bIqA+WxA0OsPS
5oGecBa1GX5oJlAf/tPgMkVg2kyP7Sz5SI+ayaI9MLTDqr0TUclXiQ9Zdk2H7BcAW65c777Uv8zV
1KDoTzPft591+PgRNXAzoeaim+jm6owXGAAP3hqj2Ji0MwaXYSKN86erVeWbyf8uNTIP9WKLnHIP
HBcEoYECn+p9elkDygVbFSzCUIn6VMJBldiDbM6Lj1TFa9kT2iQNFFLFfq6i7FQQrgfpMDsl8ksM
PVaHQyLynV1jbA/KO59lJpGFlGgKE1g3evkCpn3gJ7KuNUrBtIC5/RzFDkGaTlk0i5OTZipQKPdV
0PBPeJYR9tTHS0wzf/cPBPfuR554Qs5XdCJUYBPVhuxCSjiFvHnLnZldYTC2apZEvHWHOYM0qddv
IuTlADtQr3tk7Mr7o0Sslp3CSz2Ma0/Y3VD737o1NoRxodV5fffK0A8yltUtGtL8+zDrPmVcsaj1
liuAavrWqIesVg4VDp++l2se7bKHqkswtMzlqOoltjh3iI+labB081GJGv5ogJ47+xc6IlyraE8o
xZdK7u5QUd4RNkT6/oStw97N5yVtZT6Zc5F9lT/cb8A0FwGaDqnpLSPoOimEsGaJW46t07YvxBiP
O2B7qQ6TaIt7afYuggwtVr34x0QNMo+mpieTYi4qfIKSogteOV9chdhIwkt5gSPYAaOwtkPAf/nH
HSd7F7DibHcdEWJ4kYvzFztj2YeBqpg44b8kYsA+JhXli0Nq5axcWa88bwrPKBP7gjCuLQYORHgC
QbkWsTsq8WSvHZYwdNln7nXUiZel+y84AicepdNSUJXmkGh2fl0FOB1K/SnUkklOmMb3F8FjXB6R
A7qjgd9BmRQdJj/15JSP6qdRq/ZDCoj3GIic4ug0orte4MuE0vMWw+XjrWjpfVPE5rtpRAtWMHVg
tqQLYBj7aeCTOAwDIsedB+e8UY1Iu9E/r/3UuF12kzco/EAqBeW+8OYAtcdIyocZf2M5gywCabSp
ZvURIaNLf2bvvMeddwDnRXL8ixYi9vFfDLpyuherMvPQHW1CJ+VrSzni6oI9zo9cEyv5SLkvBjis
58/hpu8ZOTuxg6XHipgDbYInrWgNA/4AZvo4t11pmnfVOp99Fgjw5X3rS1ip+Dm+BaL794UxF5jm
yJn2Rpwd+2TeEGf9OMCrJ9pr59Le9fIRtHezqBLJxM5OR2ykl1a0MQUe7qFZqXSa8GjOILE57ncm
6WCcyCgITOrjiOrKaaNicEO/rXondOA7KMhv3xEWTlMWAWqP+COpuYJIiNgcFMoliZwEp60fL3Td
UO0H89cFhubCDMmAdJOm71zqq7Y/Z05W1yUz62lcIrMl8kM8Qw4iZYVaXjxIMkL8aDAwrurcyzKK
sY4HA0MKS59Gn2VpVHyGZ3teAEGuO0r+hq/ZGeHLEcl7k3bjRgP7+/p5goI+GMYnG24cmxZO/lQj
P3IQz3Mlr+euwGwN2AFnhOi2cBTSsd/9vShUzuyx+l7fa7LES7wpg3rFIQ01vBwha3qYCMUe/Ycb
Y9IWXPqYxX3EUtD5rWjkMvzy41mSAgsFjvXfR53H8mIPSvkgei0SSGTFU0w3a78YkpsQy5gpkkAP
IGna/mVIyZw1Ci2Zuc1+jZoqqyAkU9aofUjzHl67mZ0M6rkc9R/kkIVovm6HstG5QrjrxaH32Rku
sYfg9pHjwrjIuwHSvI24mEUvGaqTpNlBboV4RwsM6OKD2U/4kz01LzukyqzKNQJdVGt8GmvIuPGy
JffJ1iR3I3ex/UT10Bl5nlNCnOhWOhv6oJyrxs7r2fLBbiJXpFVIOdQwKfguGBQVvt09eEV2ywQp
aNDNeJfJkUga8yZdMzkjOLGNAY8ufRWvo5jq0oToqNg6xkb/eJneOWgsIYSFngKgmSS5JDaeJKPr
r8WS9dzY7Q8Xz0sebHzqIura0NPJlsBslNmUrEVVniwZmQ3phLs3E4/QOtBVy6jIs4XrFIgRruTA
75vul8lFQILc/tQqkr6fH/XXX30AYgN5Qr45VwS9THxx8zuImbgupqfQG1cT0Z478inASG/buitI
hzU+Zh2NcRgKfoCE2HWbNfDLVmN/nSviFE00STwVYJMjZA26NHD8t/O2QBWgSSNBNpkUCzZe8EzJ
9lJcG+xgEdOfCX+8u9J3buS1nGHcI0drOKmP5X9m+vZtuSctUZiJYN+oIfO+hONCPCF9M7ItePt6
1zJ5lDMT7J9S4lIQ/KyXNZcp9aEdFVFPMtr46I7hQ3UbZrpxcmU9jweGME1aGC0RcNd1iWps6ijp
XmEKefPQKPcQpAsmC1zG9ZFOWhCitoP+bulFDCFaFSe9iI7MvEHThKLf9Dk8jxJCz/8FG6CDNvsw
Dma5xjDRcagRhk94+/yWZQYmGZESh0KQLv7VP/yFqxNz1omtdnBp0deYgA1wmaPi27iaT+Rkcoin
lwvXQpTr3u8TOaRJT/ONJtS4ailbN0TCjfk9w550U/mGt/cbhPXD/YHcMFrdsefjqwAYUef/VnQA
CMPRqv9EE58/p4nbp6MkciNBKao4H+pcmG7oSVddaSyzGg9Qs650ZFFgYq5Lhx+56UtHBfhS4uTL
2h0d0mAq7x+sBfw14dyAnOvpJBfGI8OtdxXftah4TaOkUzeOkGtJJKwazCsdjHPsr+HQELJH1khE
LbcrxVBosQznvgtVaZGnuYN/89MaPMEiSx17zVIdZmyqljOMvRwergoBrd/K/f22R6n2/ooLub4P
3/ohvfhF1FnqgwIp/1NZIvfoib5fKYYF84O9UTCq/bfInW5eHCVt+gexAqe0+OjjlHTFKDE7OieN
IFzmwsvQmA63fAnOAkSKzb8HulmIuUziNWLuW+2T704FAb/jhKmqySyqpGgdogqu/D/X5cYhXpdY
68JhC/+mjgjavAwP9YkepNl5sHPvMxxpzKlzjpqWCqE8BrBD5k/ccOZrCIibaQ6qF/vBR/4HxqAu
looHZkHFOBliWRCYKyfGMgbLrAX916CWIyERQBkNJ/K+7J9ZBcAhjBHd+d6jlGNz0bldKUH2qPYI
+3yM1+z8Mv1NX1kzsfp05VEHSppCOp+wae+C1iELubz9MjFp+zXUY1y1T7uVF7c/BQ2lvrxFvvEk
AL7D/hAqAvzQI6wFkWe2Q4C0W1LMabBdcN3jVaSF5WLZTFEseb0dI9+A7VVUGssDW6UetrJ9dCiu
6Oa7LPN6f4fRFkJhTufuX85lUqMjSgbACKOvhfGeziY1/MnjWTKZ1EiuSYRA99VagyhYYBe32sHO
zbsd477ipI+X0dy9/mBvMQKFA+/hZvPD0b10p1PU/9z6RRIbo9DePlIRB0f/zPIcHU/3FskD7jbS
1yXtlgZ1mSXPqR/IQjN2JdxoE+8Q1x2CMo897FpQE6TKABFmt8wtFoNXDxNhpD3VQWElXnAQ4IsL
4b5x6gVoGdWhmFu6cx0G9D5egku4s2YD6tSlTNPNjiq69UBeWPSs3i5ZB0z6UEyT5ZFjXUX+SHpM
WepmxdEECvSf2uACK4I1eca3xtblN1XtuhriGRi4f987KJCnngI28b8TaE2G6teV/XHIUZ4+Bjly
q5WuAd14q79txrjbmqe/T39K7oBD6yCVJtj0I9CnYRP32f/MNchZ/QTftYrvFs6Bxqj9hGqeiabX
rzIpMrQQlU2N8+iN4YWc4edFRCGOI8Didge6HDz3ZcSB3zpx+6a3U5dGU+E7uPpmSKFuObaoAwkE
7nx3foKXII+jVa7/I3KcTOQFO6b3i9+EkqXZcKjqXWCMSyjJ5ZPZh8SRnZWbvAzWu8mCw6fBRVRn
Aalsrij8BJ7E9zA1MQb2UfuAqhgmiipIBTzB4BdawnJYZ7X/wqOtIEPDV9VMjGzIXNkgL/HvAd69
lq208Y2x7jfA6DSg/MTEAanWaLFs8sL4tkSsg3vDVCcYEPbrJ6EK8xz4N5VIs+wnGM+kviu+rzH6
/m67n2oGQ64H7ouLOfHU+sZVN499qj221GqWgR/0Lb3gKyZIGnbCHWiUeHhc58fyrROiGO5tx8rt
bHMYFIMoLNhuQohLOcd22AD+AlRCjcAg60IVwIJFfxlI3bsXsZ8yRVaNlXKJOfrXvvwD6RLtpLzE
D4XEJIn4IWdrNpQHF+nD7BzdcGqTM1y+XcSed1Ot2Y5pjBzkCGK/qmECmdmZVihnXhQJWtRpZdR6
OJ6836xEWPRWH22usL6Ie6k/0W0ZgQkwdZI0r9wni36GZWMcrTLZRpOrJ2nl8q4iM1IQCIxaSKq9
EIBhuLG7DwpNe7F4+bwIZzs3Q1NGFv9fzV2r/J85tU9kUP3BJTQZ6MGF3Wkd7SXCi1T0XkFCy/AG
H91GD98exTOMi97kgC0cUa8dfvDB181MfetrnaWimpfseXJ/TDtR6CCtVf9ZBXIL+7pyVl+UDkC8
gMo9abXBaGwzdio4Fyy7bVlxB7Jvlkuqdvl3IBGOSGMxSmThb5ESKAv8ryETedjIDebv8wB41DWZ
ziR8Pf91PgOAqbXspaRvLz4K6wSmy+1WOXe9MxRycn/edoYnS/zwX8hrlmja6B/qg/8Jj/HZY5AM
q0geqJxBDTbYTI3BbtZQXH5Blj2BB4nx2pfHhzk2nCuD/jH9Vq5ydKABF2soXDXM+D/LLEBdjlyR
C3PF0V4+7XcYQVuJ0muI4MM89i4ejeOHa+NxtjuZaxn5TzyyQkrzSmWS8csonsLMuVuCx0ywE/WQ
/A13jbwNToekQAlnOvYXQXU3jliUG4dY4/a23O6/4n2x7uu2BD719BTgenLV6l3ZqgOhQsC6vmbY
m6MPTq+JpLpfPbAVO3BGF3GzUWG2FWphIdhAijOe8LpZAhF9W8x1wfsJGITJ2EhMk6O1hp5Fm2D+
snrFt1SxUQchsoZD+ALdrBaj5NXv9pnQjkODKwRXGXZk4xgpzUE9QSQRbg4e6P7q6gbBJQLhNcy2
VlHuB5dxqHOCR0C+WnXTC4dQ8jdeemTbX4R7GznpP++Kzlr44kk36ll3gKK148fjsC6tdsajIIbk
9jp1x8TMfWOR+CKVV95fFH5cY8rBCJsEhif5WLcTiRE0AakMs4qfszcXImoHUPCuywGUpQrM+J1U
moh3HnbGtE4gSzGAr+ZrWky6BbP3rrQUpnncoHuV+WiLQi2BJzZOBHBm8Oh7nrCErNmK2inLkv5o
wjzPxFfdno5yTNVR7dHuStgr7D0kyIO48tDihfowLg28LfJ+K8Aw+TBOjbdecIhW3F9K64Df6bW0
8UgJI/e7qL0NYTjlIzkLkrh/94yqsLbJ9ink8ZzbbCUnnvXlR3WJcF2+utEGPHzAWg0I46eIycyt
MOE9Hu4iLc5ctV+TCDu8+M73FtVQnufKtvcz7oNvDKDKM+GMTS78qGDP7/sge7cdcYU0ZWABa2ar
EoaAsI6S3rFkNYKi79K24T6mB31jf500sxGomn+VGz8f8E9QROS+SwffnmGZPQrNogLUbPuCf8o0
ewjDW5E1ixbbw+iNYbEJc2JkQ22lsYbq5p5OWWVVciMeHPJHiO9Y9ZR2p0dw+G5nO7OseyFRUS1f
0M3WSrXunfzx/aBwrv5tjpFPIMpDlJdAAhwh75YCfcCBYSh4sCDeH5jJIksralXjLSjBUXY6muPT
PbhvegCe+/sVEBujucPCcwVcCJ1wva9HiC5YnrdXlyPpQRjCaNZAOgh+wL3ya48WDLCHWBzYWW2w
RITeSOYDiYOQ/Np9kC/daHZ2tjNXy7UkecP8wX2voa+M89XYc/D0/TFMXEa/9G21BHIE+w6CS7oB
pekEsZmi/G/0o/xQnzGUlCEjr/bDLqku2NUVLEhCRJcZfbIscpesTKMxfVM9XwuFcYb0ac6LSJxk
/0MKbBQNK2PBVE7nsZsmLyig9Uzqg++SuIbWRcX4GcjZWrvINxp20S2E8azPKjg98rjxI1Ln70uB
NseQwLVzDq2dtH4QSfpyAV/SaMBhECDaVhCptpp6P4FAcuC+srskzrugJUowDkFyV4M5smAN+FVo
lVeMDMvBo1LFr0gnXVU8ChEw9h/azrZT9mg30w6qr6EzvDh0etwRj93kD9S6jXqz1oPHap2rVD0y
TzreDBe0dzzrJIU29+11T0+7n1NrqtWAB84PIC5FFcKZTIkFagoRfLVKgquOHs+8Bbv6BrNu14K2
Key4IH650V4qoxQ+jBASJrMw/PPNu5bvwlOxYmgBJ5mBQfvHJ3L5o5WSwZ6CTxaVUz55GW3qVWtb
4zl4e8KZgaLGNNSm3jZMHxT3HDp9aFCydUPM8N8li/PXDYdBbEhk6oXYZ8iRC/4W/5vFzb0yidw+
RWPgQnj3vS4xJbh+iYy71berdMJUT0b/Fs5zgr7xH19eEqGztQyT6hBEM9vcWV8Sz42E3dzIHeZ4
ANPVST3vZLKzLgKUwQDfx1/6lZHsvEtsyQWIxuiWPRNtolpZBCzJT7uT6HK0L4jbx4+R/UYrrDPQ
k8eVc8qUS++hzrtH1qLorUcx4df0M5Oc22AScMSCVmxTvXYIUzlzdW8VZ2rcyotmy7JCDpe+dLYf
3Lwjh6hQ6Amz2aLTeSbjE1r6ymNoSXBlPPGIcqx+QLYX6RaAdcbRszt4F+VbbDSK5JiaPiI6X7ek
oAaBGXWNQeJJq/3eHmeayhpFLdD4+g2W/AP4XxqcClgGbtfkQOE9kU1oCW4qWI21+hkDmUDmC69K
uQkZN5xd856MaP5WgVAWbIjaXe0gOzLirxNHZtgqcRU4zDWAkX/uRn9UXap53Rn6oSwRhFcdG8zn
zF8QzDL8ZNGq95R76o81gzU+YVzfBdM/PTO9ugXj9ifIne8cqWJxjElilcalpbv+yWr/+f5qqDan
NC4GrOAa0Gk4W5j2WSdHB9zUrW18v1h0TTp4jUmkLBbsngqfz7uooa1BdKgt3+8/lN1bXtTMaLKV
NinaXB+6xfTZrp0KicjhdcAj5EuNvWZTwHWSYqA5xt8mBL/XJmp2ZcFPVnYVG/RHj3XJ+aaRqwUh
M2zFcGCqQ7kwbrMEGARuGLBBR9q9cWdSZf7UMi2fGpq36JEYUe8HKdPgwzfQJLFup5qa884mrmiI
HfnBVo6XlspnFEZe2HY8e70+3SqyMEL4ZddvH7E9qRjOzasjK1P4o3LEb8gYR81wzhvbqiFiSm/y
jgpmr3zHetSYMbaHvbemW0G4hATOpHilueZBN1kGa6805cb5XOfKDJ3Z98Vkx2rsJMF8djUR+gSF
Iai1ISWeEAWY/pQVMiOklZrZ/NoOXyEkykznz7qiSKzbFukaMFNgGc3sieFGKMH7gyHMz4Bb5AZL
WA5mLaelXNLVfo0VRwbgaV6IXsyO4+EIH9lbSFa8Xqn7oFABTRu9GuWma/0Hx73UlREqVgluALWI
+1VenqtxpNQ0XqOX1rK/clh87SNQ+TLUAD5A7LBeYQymflCFflHe//hi2xISN/b6BNXCrHaEUSrC
07kRVC8uB9hgVD3fKkSMRwVrOOKdNPCibFI90OyT9cGnD520Oa9miaqars2FgiAhsrEbKvCmoXda
7ojqB+FKvUwcIzu1EevtdG2DG4cXKTNxKI+YVV+WP57Gk6bfegRz2/638GOmuzyQ8GxtRrUy94NC
gAEiuF3rP1zhpJu1O/VmSLMKli+/dh7BzkMDdX6Dog33fU4PBQmgK04qQ+nbPgbzvgS7R7M11QRo
1dpgi1shSJyVnPzOkhV7IeXPfyFa17QRcBUKJMO0dz74zhIgHa2+KKTUWDVB3/4e/JPUb845cUvT
fikABsruKfJTVn2nI6Zi3egiVl8KJFmbUiIbuKE6kNIkMqzsf0xcGSrPtgPRSLwQhPkgTDG3mm4n
mKd6eFv57Ao0JSfxFMfgSe6lkRe0NkL8cPkzzuUJ34r84UFo6+Z8YUNlaxbNtCsac8oQGClVrj5F
IEsrrD81bQkfyUcFZWnKPTMKEWEca4mjaE8b9ZE4vVPHqWJVVnOVlpao+MoKNyN99WY7h+ZeRK/V
TzMsN2kenUEoCYT0VR/pOV862HDD/vWIijCOUHafGPlRfcpAKh4mP+xtqFtOCvPpRMiHeTfWhYkC
H9adwBDjnoEPP4moEIdIIVhGodAuurkkv7fPuDr4r1ISatMujFmy1BwwWT2cw5dmPsFj7buOfpXO
jV7jiU5oq9/VqbWvr1U74dNaTcAasnDNpK64Ow4ggG3613qlsuddzdZ2FHfZkOf46uj34uF8yE50
jDeFJLovxh86XADb43AVxiwnLnGQ9XqyG/TOnQzgCuMBLrlKlXv5D3ldlUuv/iZFi2Ksf/U4uRhP
XikdAMT/DysaHFM1mbN+tPWsgA/fGs6WRGwalrLzUNvlj6jYfNDDdlNv7G4yuJdvmsZ6qGaFcOO0
uHH5vgIkNRJ5C6XIF1vrdLK7bfzpny8l7nEQvRriSTPZY/NuX87kxYDLKMWoZAhM+gfmnszOSE4T
CzGbmEiApUrqGhKU36TLtp1Mf/fAexTIvb1DUI02EIhFJ+5ppkuY1cEUrPAlsU6H75cl0XXFuwKZ
koauFRHf1FrAvgzlX7KnM2KC/Bc+x8AuSFCgmLKLP1Mj8Ua6j+68ceAdob88DNs2kUsTdwjW34Ft
vYaXtQroICqbsA9aaKaTIB38MbN8xYVkCvAxoGIzoUrM4eJ2KYsYShI12BuFlCaguSi790+4KMMB
GB2PQY6meHv/3ChIGmTu+ed7T1qkKazONDpSWVf7IxJB9mJBcUxt9YnFesH9i5hFCujlotgmXDqu
9UsZdl6S0+tUoQ4+iPvuEGn8meXLckvtW3upylT+zmIyNJ2MnsFG4e+Jr7PhFy67Xwgrc8vjEA9f
1GgpHLG8T1WrfbajiDMBWckXDHR5zbB5o4pZVBvWTEXXP60M8N+X/9TfrjDtAPin3AsAIfB4+AkX
C78lWg3Heh0P1+rosIVcQpYDx24FQ23pleQDLe+Tw0HGPYq1WM/vs4p1imPHRA3+5kL1kHsNGfGf
2OHO6wHLpyit2hm471l+D7De3gQaRRylZtvqe74Fc3you3MEN182sf3MM6kB1upyXbgH6DnybhrV
sNLLvCk3Nwqba5XrjzfzdeQmTj1mG2a/UIJ9NRzkTYGiQ7RDgju8nHv81nLMZki8R7iG3yQx/NYq
EcGNILdeSIOrpKhBMcgkXwFIKF8gdJ6w31AlvEA0psinSkpW8vqr2a6DwRu8c16ueF5Njfwot399
YpsA1DRALySuQ4wGM1PV7rO2vLsXReX4RleDf0lzKaJkvX8wsJGQsGPbPzpTRFd3HpQ7cGGNhEXB
g/oiuQ9L7Racqq9CEqSmc272s+sONJzc/D8y/OuYXmj9RszpiLGSXau36+cx8g182Yn9GSE0ubqi
k2TG73WZkW8a2sMO3KkfQYLaeTeRYtxU4SEqIuXDrEcCpnnkHSHEWgKv88+oHvjD9gNDGEFb0mFf
LNeuUIWac+RUd6NE78Sf56mY65KVDwrWSf08k8AwC/+bYSwhe1ivDGbA39U+1N5NSp0LrhNGKnm5
y68RU9g8+20UH/GOL1qS1YVYYVgtffBlBkhcHIvfbMMZ3e68ATATMjhm9Xadydop4LyWCIUMYi17
dQluuf426Dho1HAXyCBB4fMwa0BR3Ugf+5kUzZS9G+NwJTTKD/tBTR5UFGrfTJSBK+/6PwSK4Kao
ZiHYBVg+59IOseCDZ8AL0CfTnbvI/guibG/QpIwUd6hBdu85ZyLkoomWbigFqeUrmORZ9rks3JHJ
5o0Ur7ZiRXplNpjDE7lH+zbdv61VgIfqCG7GAbPiQCjnHiRJ3HfO3A8bbz6P6AXgXWeHMCoovqfD
xtNumIgN160jbpVVR/6L6SvmOiud4JLvS6fuW8FV5jNcEPABl+UjcZiVz5nux0VF5d4QDRgqlanJ
RURVrRHt/ujwVKZ/VeJ8BwOCzH5ivXIaJy8x1vsS0PdPj6IATsUZASYcCmT7Sc+iymyJjnATz+hE
LMZUQg5ZXo+p915TqEWb/cjS4N4NPBM644ZmhjFDmpDFDGajaawVczWNur1halAMRzlZRRT8uZfR
o/oVX/Y4xT8j5pFjIOlWN3LB75vvvaVMsbx71ddhu3O2Jem+FioemyjcW+OnM9PX16Mekn9PGfgE
iZB75CPmwnweeTU+6aRW5LiqhXatQ//6Z9tweLCPl1GFGRMx6PLwy4A0+Gq9E1JF7eVIevijdHmZ
YAYYylBs5uYNCjC02v0D/ajFmOB3PXa+IaOPVvX35kXfIoq9MW0S4TiLCxqI5oK1AXJKUkzYxSms
ZPeBys7mpjHuseyVYtBI/fpPu5zCjMlMmxprx4eOvjSZKhLKGpBb0Z0hMoNp94pXHBSPxm1dNOSt
RmtZmaehGvRpQzXZTHMgiqqYmXA/m3dlr/OKz/XTWGVoo2MpMaxif/grFclFzMWjlO8tk73/21OV
tvNuD9lavL78eAVf3UIwUAy92WB9uJAlUg0MvdhpV0+ZLnNUWD0WsTxziZWKeFzLOeN6WJrv0N9/
Om+Mj0/WCcsyAtDwPh7QNEq3OqTb2YPYmRS2d8Ebc7Api0FFODTKUt7TJjFg+p6k7bfno98AD5cg
NHcbAFt4v5VqnxJvHGkMVG4Rd3cGHgHN5HKeFG0gVBFMBIucuuL13uBjDMcfB4rSg6VWvS+OsM+A
UCXqdn5bol64rMCSWm/I7Ie3I4zLBtkyF+rUleC+rSZdSuumglfkJmV/c1GVLMiUiIH2gwY12hIA
Qp2enrREdK+UvqHtddiUHxJa0qOxo/viodUfKOWNgyywRb42hQwuWpjz7e3rAoOOvKIBiQbPuFkm
jARqo/3heRyvVMaRoNsZN6gFywSphDJnNrF8LOP9nh/a8o0NWGv6QV8zWpVvsgspuVF8f9WqlsIi
Re4rTe3ho5FcMaba/Uy/DSasIb+DTZZHO4ve5+7fLP/e198yqiXEiKGJRGpE4pJZhIxUAL0Upb85
W5ptHIc+ptjobNvA1KzMuzNJ6Gx6uJaa2pbR9qwG8so8x0jNrvnn0i3ue9kC6xh1yVTS1lp99HhX
/RIse+Hwvh9rK+ywWKKSSmAgVYVG1uuq8AMfzBjftX7ZWVErq5+N7LEBzLMw8UR6qbhUR9MzjbZ+
gLC4rshtrfxKqzrDGgcVQ47hwwZoUaaaCab3NtBi83sPbGu6UkTb0kn7gRVvhzlf7u5RZf0/KG2F
QCwjhzsDdb9TwmIE5ptqBJGgQ67hlpKXoQOoywDffx1uMYgdmE4s5k8sZR0W5yugPAPeqTZRx54I
gIHmmam+gUb8k5ygtxg3vLYXvnnw7tnUjdmG9CCikVDRsXtQ9zZe4RhoO1eR+n9HvPtPEDIyzbAs
cB7RSr7fkR0rWumzdfUfePJBKUCBiZ/rb1CCxiq8veyeFrAytSmN45OGdb3SVpOxOemlbxxHsfEm
6jG5V+RAtv8TB8eYHssW/+tDxYmVIZZNd1hbvzrii5NKp8mD93D6jw4SQ/GRt56oKmab/t/FTtmN
xRcaxyaTAkdk1NVZTueflkHN3ujl2NVvErhUfpbw+uavowIl6kVs1sXIdfEgyjn7Eu0wrj66NLdw
UIiwW6HkaHvTPo4VN1rArmAPI9KOyATJ9QKR+bAg2Lq7rgnsRp1pMImxzjt+w1SXFnQQo06up4/B
R8Eg0yHFt9NR8p1pntlN7BTaDiLHEI8RFrrXJHV8KaSMkd+9o4N2BswTWO7Q4GUkdg7AQLcv2abE
s0iehfWeUnTIepab6a5ZdD87AU4V5mruTDE/IXBkk2Op6uXutTEBsztrIpB84Pn7xldL23vdkhcI
3U1MLZv9JnOFfIZqKizUjNPKHuRLcgLoC10puAzayL0hxxYlyXwHE4917KPQCwFJlimZGSNrwCKt
9ZG4Y1ambNpdPRb+34NTvE5H6ZKklzc41YdzZbuyxgi2ZKtZLB7k5l9BwX3OmI/GnNRdUvX3bSN+
FJ57WX92SwEc44TofnsUuzyy6NL23FFTpwwc9tYHXh5mXZsBa8WOYOGyCQ7qw9hMvgep3y6sTBzJ
RLUF+w4PgEFhRjq0b+ABH55vsyPELtcnW+i26Dorc9/x07ds/rXdi3SN0E4gm2G+KYIbxceRERf7
eCKHGSdEPTszQhNXEF6Ai0HSg4lhl2mq1kwydzW3f1YNOFu+F5kF4ZfjQ7HdKlHaujn55N1yoriA
ue0p0GGNoixlVrUAQth3eoe0dzny6crhvGFZ0lea/u37jd97xQBoXsjMRwqZIh8H2gB/GZYgSt0w
8ljh5p8eDghYqhvZK6MTelDtfsNa+CdaxIW+CVNGJVCWntaAK/T4VrcPdlhW8afo7TvLrpoS6Rpu
1jll8hq1wgorwbSFi3/VUk8CWmZCgoe1UZPnpnL7PYlaI2eHBAda+Q10uNbn7jb0ZpWpXXzmy0wv
9Myy3kOd2mtWVzNAhkYrSsjSnXHn6KWJiAwnd4BnwsbQw4+0bkUlmd1oflIDKn1qspAB70tDn7Xd
+HluT4Apl2vOTJDT8Mteb5EoTl4UPdYWwsTVSSpsW5Ade3b6kzj2n17eLwv8Ze10f5BDXAmGIri2
+VDTIyOEg+V9waKPFE4zVf36tDURgJ5b1B8gZl8H+AAZFPQ8EGMR2ZqEGmeqo9HpKWr5sE4jqLey
VeQt5evXPfBMAye+QRylHrhpULsePFLC1wqMwSXiuVPr6pCw6JMWbCU5NT2OLI2zN2PbU+Jb6yVP
C6ph2CeERcF2o8Np3fzSjwEpFACbyjzNaiRo4yudc1pJjYbh3vfNGW2BWVuOW5QX3T4AummSQekC
/3Xv6s/FHB7sTTE4886M/0XRHFeSTjMy8RUlkgvifw4yLQSBA0InBtun13jbpytfEhOwKxXxLuP7
2vVe2VZeDBKJFPMsbq9LqeBenZXYriQfg5rvsO8z0WqbfbRNqVeCY3XP73KlncXqN6X9ky7IpH6w
x62Md4ADS6CYv6o0Iz+c+6gXyUwTOlQ6gHdRszHafWx1cbJSiCohCT5kd2n3LfKufBZt9H9+bvwO
O3guI7n3X3hEUrQ1rOuUoQSDWgx1BEz1YWAhSBzjrm752QBWKiECRFlP6DaRl4WnCOnUbJ2HIw2q
+b3j5ziGv/AodpDhCuAwHVXOM5870gh9l4ZqIrmqj67O0b8Q0qJWQOulrp2qscWeK5rGHoz+4p4s
rDnAHC1qcdTLau9sVlNM+FuQduoFEAptuTzJbNgOYxJuNg0NalTDxhCixyOds6tsQGmiX1Pxe3rE
Bu17ZhrMOmAKjrS4KAny4AQNYqdxKXeQ8OzPDYU9cBWLzPlEKJfq8EFkfmzTTsGM4p3vJmC/F0/v
29V5I6I4XkHFvFlt6qHwKFrH+S9jrWJR2nRdenzCYNBQ7zCE7jgKTupAUH33+eTcSA41NxQtlPxZ
XkR+37OMWQ8X1sC53i6Vqd/Af5JGeZDexjtByyH0m1MHx1nW0zSCeTxCK28AdtF4/rB6ePwnyxn+
zhhRB7an6fg70zm2ZfIC81Zqq3Z/LLrhDIn9hnRuT3UgU1l6sg8+LCJ1mLdwdwTmH4wC8Ghi0p5O
5BNfwZ8g4bIht5pYrpazr3oqhxfo5oEDr3ljZFo0nmWo7a/0MZHOuZE3d+jF7tGeb7bC/dBS/S4v
Xa60+iu4SrLDWlCiGaf1u3BEvV4mjhBrsLseIXrE8Z8p83DX3zS0UMl6+phH0pXHel9GxpkMpyHZ
jdG8T3YSJtE/JxdS6NZ8BnmmdpJo0LXzks/pqgrtJXgPLHKnSsKBp4aJesHKSEESoQL0HV5GKuKw
7tXMEgqq2KCN73d/B/lRTLhseDWqXP7iSqYk4xoVa66hACwGAax8A06d0y501/6KLCjnjXMsB4lV
Ga4k8MREtQ2FysVsdiNestA11IIT77rAbQHGW4gqf2q4ecneLgOBjQ8tWf9ou/X2QJG3dvfNpp2C
pzvUKOpCnvt+/XJB8LhrF22K9KVIhLqRAqxXEKzIZSGcCANhrJ+3uIFwhHd5O9RgIOwjG52FWYwI
clGWzVUUYG3m1DXGBJEZFbMr7YhSpx9ctyFernlx4OX8TWQx5+botAMraGet2lf53ZVDNSN7CvNK
rOjaY9yfkilta5/u1are64YVSwRY8rJckOjgAlMvhUa7eDXTPHI77CM+IPaRbSwPZeynPs8JZuXw
HAA4lcbCWoHyKTNif0E/8iiSzuKiBY4bzuvU8uzlFmmaeLjH08Z5yZID2WoPfmQfYOmWnpGQG6Xr
y+OEQr4gkHDG+Th8Lt6/79oxWGVRUmQcY3VXAMpD04pMlzVFX3vTZkkLDXqdCZJldxdCW0GscJCe
dYk2PE2dp3zFTnQPLNgu+mTvwZVg33thfSIksN3RW/tymivs1YR+NUAwSSeCXCTIV0KGVG4shimT
uQrN5mWNpYZZFxs5JEd+i1Gh8tPy7Xmn25QeTbSbbDKdizAR19m/4q5H6owXwWSstn7EHnJp26ZI
C7G4p47k45ilecpH2jRG3wIhUdOsyMpiDIKdq8YC5/PNHPTH42cEyEj2SKNcat/GdETdgRw3Xs77
bn4Orvl26pLaa45mMVB0BDYMmEcdXUDdNswoyskUJ1nP8+SMoo3xmKn482t1D0PMwGjElRe0uSVf
dbkrQTjyqA4OjBTN8FZN7z+GTKejfY3OYT5jW3CNYNRwV10DP4qJWiJZ+tdknydQV8l9Uwa+H5j5
u07FWtUd3bWJNG9JAah2x9yaCc5qVtlkU2e22NGy60nS+Mw10Xy6EeC/2ULoQJmSUA1WouDXJOpJ
s8OZ+ZerCiwgf1ZALgsxhx5aw8dk+zO3axpSDc0Ji1DyjvIdBrcIO1ojbjIp+Em7emmZ0AwrnYZ1
LXfethOZ+zphKVt173tfJhawC9iKvtMSHQL1dHSE20q78V2vFlt7J9uM12p6UbHwYPUhG+k+rFqI
+iQDOOTA42I7wH9dh1D7rjyx2R5Xlkmuxis5jrvmiymW04+Hh1pr6dEEYPFez3QfTkimsWwdsfNT
zR/3dxveA89fXssKIN9ef9ER0Dqea+A9qoLaqihQ9Ln4s/i2gzMAtx1nSghW8KcPYCL8gPLMAZXi
E7Bw2Sluzs3yGKw7gIx1fMM9yPHGfBI3vAQXVDEhlt7Oaypl7OIVHl73ZRFXaYWecAYwB8B2JMYl
DyRIrWk5p//RNLxUVtx63n7wkZbs+uYdaVwpb6EaXrDIJ0cxpWEYcQGEo1cyX0pU+ErwwGCtpdVq
fRGLaU5p/oGd8QjGzH6VXbS/sSGgYkyigeu+ImducBrcoVvezCPq2pCvgtfqcoYalacr3rU0RZ8v
yXJiCUweOiPc92QIG704vr6nwRLFs+N4kfxgoF/HUydvSHqhA4pNi1Ud5GzKAUc/d2LwR7gUjkbF
lfYdPRdJH9V7HRPhWqB/n7lUuv4KZv+eOyU1RZVgLRuvKqWvDH4SUsVtFVCh3fN4T3vlssJCruSx
FUruy1N+Mc43SRtTGGlDO+XRGYrz0r7Lh4m0fkDJ91CN1gAwLJJiwml4KD106aXZKRlB7SG/2HFQ
aYXad2bT0Y84z5JmmscIjezA0Rx7ZxcBqcrW2ONK+CYQnvtJMXpoSnhFkzJeGVSejhJRxIs65bOL
5fp94OWuv6nfJoeesdYpZGepCO1uSvuMeKDiMPoTUGye2tCA7S97ypa7bmu+pY0b2oSzFbpoRUSe
+Wvt6Dso3WYe6iV24jQHPKxvz6AdoMeoh5r5L/bZ1g39MQShGcPZK8qTtHBLBpUQF7JIb8UtYWqF
fvdfWFHnUXc7k3hbkVL2/zeTH3xpbsHycXOPk3xgCQsSGMpmFaJ6Tkj27AXoLvEdmZPJAHAfY4WT
uBwQtXN8TyfpSJ7thAOPTCXHmrnrd7GbjLsTeG06rwJNvY493ma4eQt1fPllC832TwVE5oAN3U1K
1EpqSw539/rWuWBPn/82yZ1hkilVRF7IJibpacMVkmnxygDrZC3hnfD+FfdvrOK6YTSs3/r8RAKM
QfvmfRWYRtROj9zKgl2uoyDNzRIT6KAukkghUvScggB5vaTqKiy3JYbB0h4QogMMPk4j36BoTDhq
GsY3pkvAJEc4yHlD6nYcxGbQPesqqEhrmUk/ACyYhPem3AfOKdIrWsElaAqjjG0HIr6Sa2b+ILCX
/XsvD0kNGvm69hfIudaeuzPDyX4iToyC6tCQL5x0WoKE+AOUEUFt1dgixIU+wMdCrANj8eLdNGQy
QOUfzIrA4nXME4by7ZViS8uCRBp+N+M6fVDhcQa4SpQ9o+vo2vYQlWdWLuX3+G7WUr0dyA8Ncfdv
fnT4eaICraqRFbqHbOuAEUC6ChJz+RnOmQubsCXcRq+XOxRlJplxFsMgOzR1MEM7v3cRecKcvV3S
c793Z3ska8SLhu014MbZIbaNgefN4ijNYUCbGAUCsdH0wRB8iXzeP8Y1zk2eDZKdj5iCUcXyj0Ub
CN12OWvo3VU1lEdp8exIpOIzGq67O98w1YL/MBadvVji/fKLpz/hJO1Zxmua6dJa1ZIlrFsxqyfR
cxbenEgmpQ5RNP1RZrBu0kl4cRV3TvroGrqphk4QJG8yzV5KQ5DhG1nbXBX8HvUQ/SsdjrriwKYx
rYzwdV28x3J/9jqw2/UablUtryS3Di4u0qEJ/zQt8+Wuv43InSas5XXu58DOTLiRAJ684x7z1gg1
cunnP3OUylk76ewKzcWciGTnLuXC0hM6L8192WMQBEvc3bPrB8ttGIyMBvahhD46l+/JkzpLiMrF
QbiZGxZRFNV9ButBtkNqIcn3m3qXfIJL2G5mmJLLiVX/9WK28AYi0lSoKAaYyTDgdPQZaZQ7C9uq
rfPEhwBKoZv4RTOL3VdYIoUbU2xtvtU5ENh7HGWLm7ia6pdTwbDY+3ViaCvLoairzbW16NfABrgs
0V/QIESQNqr3KEUzhfrlE0cPpYX4QioBlVp8Dz2dsdtZtVvpGAQS/Ky/ssPFcF5T9DmlP64Epbsq
rfbC+7nhyIPoAeR2S/FB7kwtxC9bE0eJwx5VJ55YVaffV6GpPordi/vf8ixH++DVSgvME5hlx0j5
+Bs07xJ8leikFxZC0gr9M0g5/2unfz3xGyBmCATDItekiCDAjsalHLr+PUQX5MXGTdBCErKQS2M0
scOdf7tVnuvliMyQFxnLF6DBEpkxzMIkxeCy8qrtKpRZfHzmyx7B3gjErRny2XunSmiOSh3LKRzW
6iyiRbe3joxBierUCrToENfd6BrqHMxwnlL6SEtJ+5NwBn+1AnkZUkvhZNGnZfj2guhvKXuk/h9D
j8SaaKVS5RDkdtRQiVqrlgD+aIiLLfcUeDqWVCZVBJtYphRDjt1k8OhJpO822s/HikXDzG1JXGE8
Ml1ErircnZWQdC21HnX5bUZKg4ONwih2CYACCl+bixySt6IGGUyVoAljdm1gPsIjE+pruImKDKil
MlYFyhgbF2MC+xr3BIPvs+VrqSPhSdeWNt96SQtZPjR/DFWVpbS8ht+SMASyKyvYqydh+PWF5Sy/
60wgWL2LaGyjbYgumi3qRSVmR6GGP2xv37JfGO+bXZKRA4hLdX3M8acpzhyQtU7cvl+OCCn6RI84
7Vk5HyGNSBpDOGcT22M/RGju2ls2LeytMy1WvdeXXUvrLR3Vcwq0wR/TEUj5lhb5gY0mu/fPhgtJ
6N7wkI/DQVeERlJaa1HIgH4jTxWPODbrTpLgtUcVA4RoicqhAI6ejwtg+6r3eq6yBWrw9EQ7Wfwa
d1JlOcjcDYsJX256H+ujFgkxmT1H/zFC96mn+vRUNUsXLWnZiCek3FEjtKFRO0pfuDeK+l/S6G4Z
NGz1IMiqT6dATXjBxgZrDOMY0sAXiN29y+lmK+4PZhTH8KRXS1dtEXCL7EerSljLZaOf2KjLnJh3
Fm/Ek3yJNJ75+FGLEeRBsh4S4BGCmb123A+qgTL2ZoUwaJwL42KPLYNlUFtoRwjV6CTrM8uszmQ7
kPTZQ0Q6/HTgNl/ERdYIvpI/PzSfM+shj9yFhFqGGUmkZDzwWY0XMWIlnsdB/kM7rSfIUoSa+tmk
yUXPtjfwsLF0btfmUu0RzBRina6MUYlqtoQVRtcyTQaxmfMWlRbsGnBJPeK4IFYMk+5Yb7KerZ7v
T6hfxOjdESRR6TmWWrnJquTTrygGtjs1uYZVNuhhWaKyZTr/qU5uPGEwE78Vi0MFGmEev0oPXOYP
DMyxsiilXQLPW9ANoJbcgctWOLxSqYmhYMA7nDHamOCS1EMhGe3SGqQ8w2WCA0qvi7RnPceD5fKx
EFCfNrjI6s9KJ1eHEyiN5pdN/Jw2toURuc/liwTNzuy+qr9HU+Eh2SUI2p0hTSdG2mDlnE2SXkqK
v4ny+2jcSt95gmnTEfvG5/cGWxF80G3XuuD1G6VBiVwn3Iflqgl8yNrcKHcupAYtVXYCBkhxONNL
o22d6UsZLI048yoGG7VqnF0U1q/cYsveHNd6dOC754c00qMB67MgCbknUPrWp23aM3MWfZ4Z375M
Yg0F4GaP+dpDCRKucmuT4wMovCqx+ykxRqp13WH8h/lk6DzEpUpIiMWuTYptIfy6yo97AFB2kcGF
oCgRtgLXFEtU10rM62qBd7BiWCj+rqkssk/E6/IQyd2D8obDoWw5xTYwQreIUp2mdGQoYbh/KQ9T
Nyyb34p5VuyfjfOZMGGzdui7I4hbe+TB2LeozNo2zcG97i86NlU9p/4rEJ6uhvebquCOdt+s7Kaz
kG6Enn8H7tq2OFuIHy7HEvVvp06Do41zf1EWXHR06rLFTq69QGjWwPbuNsUsFRsl8qwC4X5y8Cs1
0GRCCKyBZTOLFH88z3r27a/QpW6ldbYMu1QMs4WxhBlPVDfOB5+mtoz3efgkk6IHwCWmt8ylHjvq
Bv0mPM+vPdOaaX3JPw6N220qeqY61lKNydrxM8XMpl/HSbtbTroLAEmPTiwEXWDSrDNDR7FZhRT+
aLPMz/bwNZ/6ry5UZMzC7qUv6cOguIan9q5BFaJJNFbfppVawvH+AEq3otdrqTZ4MaLE8Pyu7TBc
ZDlBzcbWZP3O05CXoV6SxdUlg8UChNXvDG1y1ZWIK9U3ei/YUZP0qXnfL3K2R8JmZz79mCwCXj8L
hp0B5d8muRrF1H7J8RFOuk4624j4PFWfTsHGnw9IWK7DNh2IGbY+zMbmaeuI7Zr+6eMlEBkfvPjj
N/379dnHr7aaeNCOPBH9+EU9PTv32hiCk96jAhKsQ4nXtJTwE5BRksuTyamrHE/1g5DVr+sbN0+h
XUMqqnHouyo5VShNwOocPP9nOqz5ki8MBjZNiJSbuGXdC2OR1+mt83/MIgrM78AR4MVpRYIVygaW
2O9eVW2tOIXDEjKU40Obi1j1wJ9gfXAaJ8GsTaEzLBMUmZhGQH30bv0YJPnPAKNAnnPb68z8wbyU
H6IzdSXcpL9X2NmCOQKVAWAVEnsnyqETgcXvgiX+tTZuHvKvpev3qaNcRayECryH2rWfZOi15xyD
Ss3VIACYJ1qa/uCGcCcoCHOVL/FLx7VnTdG/nydMJHUjLiradD+11mX/MwexBO88tZGEBvP1reFe
oAhrsk/UV+sOMuPqwAHOMSqQDfNqxH6DI1XJTXElw/iQ0l6iXgJqqqaIPvk1uhDAmDdGsnegxg25
2z51JfONS7zKVTJOwMNybIVV+R7DCLjSf+kp1XyLB8OZwltigYM7/tpEaWMDCLntFfE8BrRMXyHb
pArFkLUDFDYlaYx9czKn84vJ0/SUJENisq5v7pW2WwWRrEg3Qx80k9WEG6lgqbJL8q3Cxz73iWih
ofmrfSFXD1apNILocToPoloSis3kB0WH00ToBEShpTpxHVRWYaF4QmKocT1agqcxsUr1gffXf/6/
zwkB9lIX8eBhP6oAhYc5Qd6FqG50DEQhUH1yF4bLrYw08Uif5EuXPeKrWNLYVqk/VfyY3b5Tgj0s
6lB/Pgk2tYLn6DTwkij1IMMmvOEDLnyWiewtlZxP4kab3KyV3LatQLfDS4DY7YyArmp1ZKztjj9W
tdh0w4r+2MeH4qhUb5Cuwwi8r5WtKyC3laOOmS7XlibTGYcq7X7t0Ffd7uWYpGUvcu86jpT29/mI
e7d1K4JYbmSDp6I32MM7xgaZE/lodPttalhhLTVhIixT5e8BrBV8IxFVg4gh+PcGMfpwQcH4He+j
5tZv+CqZGA0UJPJk868q5iqWKYDeiEpFpCMFhCMmzY57g6EkZxgPCubhyX3U3bJfp53JZXkDgceU
zusjRB2J18isuZ/4tsQl3ZB9QjgwcB6dUFGxdFntQKBoAECRmrimPfsRj7/SmiekoJ8ddDepZByI
Tk4m1Nbx8lApnMqZ9CTJ8Ptz9Bh2wQFG1hZgHIo99G65A1O8P6gZwKUheHWjZ/BSvtLc7yul4gY3
drx0BPD+0uA5frFJht/KDE+j+2PY9FIMkXZLP126BzyBmhN3qvtwWkWWEOCL8yqknABHo8aKA98E
IXi3HBU0x+8bn8xYh8q/gIcukPsv1N6W+WqNTSVplfWQzQXeJhoVs3+S1bPET9+MATa28gDSC/yq
XdFFKVP8ris1x34n2Zz9efVMqg+KFjdRwIpwrvwqI8itdlJLN9lpODzvYcviUOH0gV33jJVMkDly
awh8W+qCGj28wJdraWKZY46tBnxcfES+RZTJtxlepodD2lsGyflyDwOPz4PS7aYym0J1Jv5zzkZq
xfYcM4XYn5va7D+Dt1QrTcOevVYX/3qRN2foyYCKLN6d6QxAASEttS3afC4w2glLqDHhvP4SYay/
yh9fqoHAiSUVje6SFFELboNgZSgVMbL4U5rEBmplfKU0bGSEMLDJtcUE/rAuAssSz0eLqLkX0cYo
/NIF3AREyQAf8GO6XfnZC0FmvR+RbkdLC+jFszF1N66Ai+2/xyknor0aP3Z2SOotuDzP1ID1DZrL
nmc2dc3zFI5snowWP06x45x2m4eKBGAJOKcBYG/ww5uG5/TkY6IQ24Z325Sh3aOwwEMNnT0spc8p
Dbf0bpP01MA+PC1kE5OtCBniWkzWEEix88idbaUETHnn3WM3i0283RU3j+y+fcjJ5inbbAUFX08U
dLJwUTVWLjdghnJKylIUQFXBWRDrgP37FY+eFf/pMtO7pKDe0GtvXqZCbHaAWj6AYI4I+fE6nsNd
vemHYtOl5iWvcR/YxD+MoLXcrUqZuAfJEAXS1j94S2nTUf1gFoBREG9ogtjsayK98gh2ecmDuBWN
XQawf7niVyj5Lux99eW6rJIwCQ2qZNazi9ZbJNUnvmfwmZtYAkjuTPRoQeKA/VcSRwhZu6T1TyEq
tH3xsSmLAiFK3hyTdwS+ImeVri2Z5iyT/ZT5zLPbuRgiVct8A6b4r+ha9R+aUnrG8t+k7Sc7askP
hjYujSY4Ht5v2Somqn69gi+pJAUbEM2SgPHs50+2zxmOR+sozca3W6uIwMPGePlGMoVz4hrT4wlW
jfvFafy6pTxiK0KzyXU2JzSrywrdJU3A3EJbN6z5MkyTErfk7ylYiBHkBLfm8gd0AJVldOZ58ETU
gT36YtonuRujulC57rvi8fB5IT4hGt9qmCmIrEqbRy5RW1UI0cbIUXS7TdFc6gciVdu4mjo26V3+
ykSauMFhA9oliRmSDYrxYf7NGUDNyZvNvPjnuNR7ZKDEcJh8qI381n9XPCp6B847GDggq0dnxIeX
I/X9ftnvMaYakhjj8OC2GrOW+aleibeSlCLgtpfrjC0aor2FKV0PKfq+JNnl9y7er8H3bmGxUixU
Fj2lFZEHqAigxpwcEDSboPT9EYi91Yew46HqK2N635Xk8dDHNjkxSFjXoQJm3V5iVjiW9dIwOozq
9a0eXuLIX1mzGmr9U72Su2Onk1qODSD6iCQ9ZyMOfcqxmpJqoj0wiXDb9BjtXJNwBb8zJd4LjehO
X2KxF9dRkNt2gG6ADxVnopEjtnkhG4/ZuqOJBcwTsDMOEaro7GnRwI2i69bpJqusIluWodrZtkH9
YK9OkgqqGIOlyYOvoNg8k2tfhjjgoUBL6PSkP9qVtAsMbaKNMeiofGUNTdR1wKwkgvl5iKv/C6fD
mwZCu9N86xtnigqLmdI9g1Wy0bq21BQXvdiJO+ibiA2ravnSX94K6NP1Itid58Pp0wgvfReBs17A
aiDvCOCiLtgme3uwg+Vo0cCXUmb+JR8q9XEAwFpnlPJxv9oaBEjMoRuiS6P7NqrXe1QVsqUTeFQw
GXLZfv0Lvrx8LFlEb6BpZxPhpicAhacoMEntE/S2yjBDzsQGA9ep6qvjCfUYN9Nc+qGs82ozw7in
kB9OrBdCRg0kEIZmlDj516RSgFJrRUj1u0CjX9dbGW1DMle3idXZcp9t167xrdNOkJI5yLMF+4QJ
JIeJHumJqtGfJXeSRr6J6K+2QT/Ab7412+3xTt0UOBpwrmTGjTxxrfK+qe5nfDlRZ3UWWgAy9vby
F9X6u+TxKz57H5j256ksMoWtDyxbFRp3fvg2On39mzNvRkGGQV3AmSZ3dUAfIQQDe5FVOtVzCjkP
uoZkY59M9FFL1WnC/3ZNHLqErqn82nbj9IdmDkGxiT65wpzrFy33WZrsJiKWCXGvIHOdrMGecVjF
3eNteTPaHuEOeTXRCbm8gxJzdJuFN1y9D1hfsuKOqb0ez2i7s6/aglBfdDiPTTCmQP2y0WaBQXCv
LDDq3KgT2p22+iBP850CjVhqmg9skgzCaYa+kOWe4ISZuAd5is9IX5+lipb84Et8WJXuOKS4OuzU
3yB7OatvEDyc/xOeND/z8h8rxPxqndLAl5dAZIu3SjtYXucXT/gqpA9dgd5dwWYSGIXop7Szuu/u
rO3KceAs1SRVOzGXKPAIh35vS6Ytik8vF94o+VAg785quZbkxZtedOB2WLchRAdFfXrVVYxnVuNM
EQf0OE3mJ4LVqEuVUwQwkw+R8pmiYn0nPnSi4XxlVq1UHiVBX+SImcCGfYslqH9WH4aQj15AvSxj
UL2Q4jWVfXMZplHjrqv/5R5m8Cctn8mn1GrrxK7Ryp6ConmuSdnXJiLHT229kSrf+C/rGnRXMU1y
bil7ldXsM0Ri8vFtrbq1PPlag8uFm4Sj94kqrh6e9dE+BzYvzSwoenVRBYOkK6UEvmx3bC2Hnrcy
/r0Sykm4ExvltPIvYl8cXFbTHD1sKcN7aN7vwQtIU6a2ZpawNCkMQdr8xG1hT5/6RNg0Fj4UbY5B
IoWxo8R5jLIUhLA9tvHPQGY7TtZtT6I5YyqT5FaSoKmXNZ0XTRb0ILL2V3dXlOKfLKNNxxYE/4rh
+q1jG+pKNjVAIUVSGcFBm2dsEbCcKcTq/hL58A0LoGgdeJxsHVI+YEG8PaCBPGPkW8hH7E+r40q5
qZUiukEgzNxQW0csxsQekjrhyfWW6IoH2uvOIut3iCXenoE/TSOXk3CcttmQs3iFFZs3XlHHXuCW
o0Ul0d4AYRzYSzsHmGyHQbRsqERUPuosEg4DXc6iyqrada1C+4d8VREIbP6YNHKGT5eMfThSoNAM
cM5yZv/Z69FBc+Y67z0j32vAbuxPsGXLJwav5KbUZJPoAC62W+GQLEEg4hDs6Vzja32cFJv4UNhZ
TMTBRwJOSAcCoFsRNte6fWf68tV2d8SslGuhhcawh3Yb6/FaFh9uAJXXMobt4zWB7Bz5ZCn9w0+r
ZDpy+rXoeXZR3ATWIT7pqtR08/vF4fOlpPR3L/zYmxwEOPmB/e+TP/V8yjMlebL0mZjR9AsKEZf5
mgdwfXlNFqFmZ5uUY+4e8gGqPIJhs6CtGVLWWbs5YKpV1tuHFaYwn8xP6YeaD+bzUl/U+U7XlZoP
+D30H2bmW07LX0hh6zVOh4KvKmCIRCFUVsUW5iXThDYpGAXf15jH3ClXSkWvSTdAiBpm57rkbrhh
rFdMOx36ZwpJwm20C8Lxe7Tc5SAigKqx2isLzezPBrFJWFU1OrXRhZv9RrUzAjSy/hwvfdAwaq5y
3VH0OyvKqkIoTS3nxVrkYS37LMPhB1UofbFrJOCi2GstWkXVodfCNnJFxniXHpKqe94o2zCzlxI5
fPyGVT4xXn4x3iTOokXaz7XtxACRbIU3BqGmdGqF6CExxXMpmJekSg5oCNcEHdazjmxJygoMJzlY
kSRbafRqqbIpiIZZlQ7ejcC6rxJXekepziwnatHJxW7tThjq0N0SIxkHrKQ5lSzwpQxCXRvUsjcT
eh6aXGdGp8TjImr/SkpJfYEiZazJbuYiFiTJ3LYg32RXPjCr0Dbz7BcG4EHFgj5g/pafyOp8DmKw
g+TtpoV2KZ5UmVuuzDXSkT5p1N8fXdvL5uEDy7pjjRQfAf036N0y4VF0e9Dm9ZDbB1KXdLf3lsz0
CQTWtKATqNN9xqgFJK73DA7ftpf2LPyptSdXQKThsOpmu8uL52JCPAVnfAMpxQD5S7ZdsQL3PGAo
K4L572Lcj29Y+npEORqYh677sHyslPGAy2fLLCiPydkmGwyLMLIswJF5cKBr+1MaEbzMB+5fX/aV
aHkPbYxQA+xre2dGCGVH++R8l9iDuMe+JXiilqHDnRrMk3DMTxisa+quoU1vyAkYA3iuTToC3Za4
PiGIGGnAI1We0SIQ34BoBDltC0YQuLGPBBPpktoZu0UbW3MiZMku5iaqqFIx5CeQNbfk547OfLYv
bS3+6CPXpo1hPxdJuzTqnJQdbx/xVjbgfnKSe/cZKhANcaFbFBDQxVByDzuw7GT0gVBR+NEueyUq
7X3V4zIeJPSLMEVUtcWKPjClcishL8RQ+6MkSLhYpT7TLK5Uw9UsZrwi6yNM7x7Ca4ZuPMOBdESx
J+S4vpjKvRW7o0zZyVIg6PBQUk8Zjddvfa3bsW71/XWFGQK7Lq+o6nLAOhNUr1J+jG8WSq0xZQUp
w4KFK65aDPabii0NEQdj3nZhKN8UD5DDijO2N7BOJMo1motdtdMPf4AqwgK/l4K3YWps0Gs6Ui21
Y5cizk+3kl5o9nZEYiPZBnkC8395I4yHUeIgc3AuB8lFVzIN4ELuA/Aa+00eihEUjR4foPCIE1HS
6hh/f7w2cvmaiwoB01LXkQ6lYTPz5CRECUl4ttQ+JtgbeXI0QrhNAeA55GeTAkcwpql9UFr05JYO
vlg7/f6UPOnbtJ1JGMLOb59lwnP5auZkg4aSXRPH6c7qTTZWA118rL+RMfZYVFqh3NIZYliLn9rZ
qlQdPOD0BuIrDjpBcZ2uqhnk26CXa9Q1j4XhHxAYRDKiRzIhKllZOPmgnn4IDy7fehiYptBBJCvi
acXbWXPKseh1iE64eND4net892HjcOuhJHGutFkN5k8QSWmCIqdE5GXhs+izKvFPR9Hnkznkw22W
Ecnx5SAxmDXXwlz9hu4+J469shdTALiwJAvNQhY9OF0zPH0hjQ0tczbUF/nhupuAMgTl2gkPPW9B
kNT79HCx18qKm/ZlCQEgEFueoOhz1q6DPJqBIujr/q0Vr0KdkBDOkFtDmQfpnjfV6OJObr85Dda/
Z+XEffAwPG3ZTc7jfiKUZWBXmeGGvXdswBhcOkeeb6OaxcgGYFE4+N+fxpkJU7iQZ9CxqMSLVFRj
Au7fGIm+X+6aJzQdWm+c+5BfRDm03ezhmx7nQTyihNGosgnkcw5qKJ083QucLdkJI0DrMgX3HIlr
SH05g2kbsmKtrddKFFmGZnWgdvkxikJBUoBKTacqors4xU0gqQ54PZyix/uVSNWFX5rKZBUvwpHF
dqS64qpjtnSJw4owmt6FIY5VBrQzKDuswcjPgOf+G9mi6oGxA3x7yId15pXjGeQ9SIjSVK4kwp2l
xuozJOUDbv3p3rwikWB91s/56Zle2ujpt8dgftyptxDdUBkpJLiMS+wfRbz1EYZzQA1xyiQGtQBN
a5l+rnd2nVGLYn6Ft7cj02SwQraT/z2vims8U8ruqEb3lKlvWGTOO7QliNUxnDsLMTcdbt6DHE75
Aw7Hd1mOstePXXxa4gXCjJ3A3nHOdD+XBkAQNmNNg0bvDTWfyeHj1ajpQUe6oz8tDgtsaZAP461T
DtIB1d5+Y1Fjy5LkgSe4TZgTK+JSTq6QmvyQaiyvhuIg66jFzLadotmd4Wa17GioqDPSXUJl99+B
iyvs4UaauOO+LAnGj3B6aeqOGDUJ01r5z/IC5+ZfNujx1VaWd9J6tgnruRZ57MuAAlCrzQhN3ibh
/my9dY2snwJs6mYwk+tfZl6Fge4SrC3Gyb+p655KPGZH2tZHe9wzM3a9kp5Wd3XF+zr79ZNgPSLZ
DdwfuvSpsN36MxL3Ro04pnH5ckZGCh4MphPCAZZRfSqr0uesl9Jf9Ax3geQzy86tfmyBydPkzv0G
mus9vkOgU3nMR2wzhoVCxs6zv5IuR9MOPmMXLnf623FFtCu1hNN76ALT1S8G7DJegvJYI+o7JiDQ
OB4UDK2PSSkr1HNvW+B2ZRgD3H7n8ukmg1i/QrXxePKMVlWuq6bnWxiV8wVXUuV9EK6DrWpvft6X
L8YrBt7YyAhOdm2C/zy0CSDH4tSKY7x9+GbA6Pl7pHql3U29ATa+3D5jNB42QC5sNxwNAXPTvN5y
xyzPU+XHqwvqGw4f4/QS6upuFXTnEIvT9S3n2+WK2DJdOmTm6lq/eRU+LQdRJu95XCsP8AvoLvwq
nynyHC6IU3VskOpsgrtWlVZJBCphJQ8oTsMY/HWS3DaQfwlTWDuJHCX9YJWo1CInvm+tisajeahv
aVExMtrPgnK150h3ZbPqUbHDXaoWe5tfF9xQp0HhDZhdRY1E4XaUNQ+UvrrSre/irP+6efbai7/F
+s1TcWq3NxfsvffETseXbTv8kBpqfwQaNiWPAtUbOGTQGZmIIcSHZVCq9Va3HXXQI7mA7lF96kbS
hUD7N1QKeNpOVi7v8txfVZnM1/esScETxtsjW3NwC79szF3g6+sdjIhJMMga7y/YvcjP10G4QenW
OIpsMHNMBI5xCPWB09nLIlpPuM5WMw8x+lXKo5hs0LHHB5d8KVcuPF4xB4TJ4vWCv2I068stw8OT
BsDc51Rwv7oODlCG/knitvE/lXePU0DUm6ntWgTqOTsBBZA6sl6GRgDUPatUjrSH4JJBYM+SxcMQ
nDdIqffaT4+/RFrVMHATgaHpWjwWouzZn3ZdkA0Mp1/wx3AmcgkMq6MI3PnS7sWzDhOpgqm78AwQ
i5xZYjnxNemiJQRPP5A6vpk71sXa13ifNiwVLxCtmjMOCxAjM2vuS7NtHOxViIUSWv3tR8BJadxe
RBSzuntRE3teQxGpoOotitGWJL2IGrRrU1dp2QKEOlRpfBGOGbQrmxDXfQP01cd1Jz0VzQmwqQep
ltrynx99IwqHLdY3FrlkiQWLuoCgCdqCXl6vZpRXpGCcTst1H59xHwh156A8YkMtak/8eCQynd/p
bC0bh8ob5UyPcez5RdU94L2AFy0Q4IzOvI857J7tRgNqiUqqRPbNoIljM4dqC4xTveeKPRDp0VeA
xKam1EOYrK7hxLYToMtU9a/qlAQ4j+YSvn5E30nWGNe11FvhtIo3f/L01qsRj7c5ggUkdUVkm6nB
xqhlma1MYXT531UUyFNRLmB/aJMlm+tWZizW+1p/MdXtbkP1Wf/gxlVMiqkiPPGsqTCDzH1ENrtQ
y0QB0513/CX7mojUP49YF0PlRUdr9nI3PkspBCgTfnWOGu4jOuY8ql1Ycw8dX5YlFiI3VnCZVCHl
SW5GCnYuoiBdlh+wyTJIjLYNBgxMxmYE8B5BFowNOQvBM+nncqS7F6nXNfWnF1VvUzK9NxOyIc7C
PcGGTmYDcxYGDvrAoRii+NreJ8tmJd00UusZKqyjSXXrJ+a/Z5l5ACi56jrU+9+7R3rSKyKJNJdZ
7gqLeBwZt+gCcyLuKhbgLIPlg39qvdAtpDTg9Ult89qI04lDvUKFHCVi2LZQdGGSjnImWukhNQEM
ZXceQE7Z+D7Si1ZM1PLBkWfDraNcQ/yzPWdL4bTFMykM6rf2MxRTIkCPhuDsGQBVdP86VcyTt8il
RYSo6rDzm6x8+eyFZ7owHFxL4ij+tF4w6lKtXOG8m+83LwX4eLvCETvW/hj/u/4ZGDGnZNUmZ+Il
CixuhZZfwqDRKChAPRD5Exi/YRQ3YGpnsOIE2UHf8YqIgy9arxmYlvMJ7gfBeUExSCbQujBQ/QFt
+jNK30bmKsiCHUCgPvkSD6nqf8yL/fn4cuA9TQUxHDq0mmYlFlGHI/Yowb1e5AIYLVaBVLJGh/fu
kb5WcIIGNd+OCrLVqlPfPagu/GaGE0lXLEr7n7PedXU7IxZBQCkX0Ok+JTkTmP9SvsyJS9UyxvCf
Lc/KMa39XMMszOwEEDHvcFvX87utT4ClhrRKiVSzQXr3NcAET+WHxTmitwROX9NzcLslIKgSPqn7
jDtJZ1/XjFIxlL/69mTXlggGy9HglpZC+1hZL3erYC3kS4NvbeUoI0mdWMl3w/avArR8TcWXoVSF
EL6LBgrAi8GTC3prQdwHroGxhpRJxiJJorzEsBPByMzq0mEoqgJVtS9feVgH/5CLrQx/dr/p0U01
YhEBe/KJAw3C6V8Uv8hi21vbn3MTPA2XtYKR9tyRLe01QR+YkXuM2pjKRFplIv6Kf58P/CE+eXg1
vL9CfYH7JaJCWukzrvHWxn2eEvo2bQe5FIDiFieMcLoRQqz51DFOV35rLlucCSbEWkaaORmicBbJ
FZG7tIiGjAm7Ptr3SPUTbVQEI7v0gOUHiJDgsEtSBpnqhv+gmCxgffQPASBftEDvk03htE0AzH+b
eDgH6co6rsO/Oasf0bX3FiqK75O/mtuWtKmjjeUe9lVXrQkaOo6W0tBJBaAXix7OY2MdzUFR6Zeo
t6+q7Vpk5sxk1caCe28kuCQSRLrjhg0bgrevTSWZWEjmgBYwjR/GljBYLbflcLNYQ/bp8vBBUL3P
2mPGDA5RJeAIiS4oCI4hDiPjXDjg2Apx4sWzjywRMCYaSoaa3vhjWKBxo6vSjoxu7J5cjG6i3xU/
yOp6QDSkoEc/XtqAUFhR3nvJEZlpgj0AXM0FbLzJbOyaLUq4HIuJjUqt/vRGXcY7pS/oifAFy7u/
j0zE6XNQ0bZwHY9UPWSdKuKlznCkwK0dCYNcsp6q+n2NWJz1J75cj7shQrj4SiAQsZylqHFQm5Rd
m1Amx3J+7CTBmO4XylYVJN9ajVdSEiSPOAnIX+fXMH+JqZ9cn2GLy+9ms3iz0b7Vo14QyscHuJpi
Yq0F5frse6EyZlvKx8Ij4MYFVyXRR6DQYhQVafWP0mZ4pTBGlVDaKdTUhVNOOPxbbUpj2vzJY1hQ
Tt2/kBirCbBPqr2XlY1nda/q9Bvwfk1gXFWte7Gt3UblUc2sA6wj+59IAPuKnJJZQwE0SiEE9Ge0
/+HC/JA5QBQZbhWtX1UKeovwSLUikXqhHNYDkNJ1EmPmXN0d5IfEuOakiGCzVgQBgnOo/8y2q/F8
xJwZ1Jum55DhMqYP2f70y3CEvbHLx8jADToKXshD+IeT1CPxD7zS5EwZhvx7qFs/+aOI9sAqdrKu
WI0J0qJDSDJT3mDmTEy652LtdNOqNF16c8FVqBmJnK+AxtlOUY+sGd08fr1OIo5UIezhJoWVBc9H
gIZWRTyeHVF4osufE3ZfdNIws+TUEXSowAO96VyBpZqLn2YODCbUQxedvN+30nJ6gshsX1Sfw2j2
OR+3FR0uc4PsK6/kMmv/BXXLJW877rDdOEu6O2H/IUe/xIGp3GGJYRWL5jEyQLfQITcZAcZXqZIS
/iG3QYHw4oDTEsiKc32IKAX251up3JnhZQGAXYNeB65Y7bc8IwWzYZTfaDL4t8YCci7xu4Lna39B
/MZtD73vHPlbSCYtfsliQgwCDLSAtzUEohQg2goomxPOkn2kr33WomvwcJTKPVEJJtMBIodzVjHB
9ShmBz9n3OtjeCzRqYiWW69FbrdcAtwW/TAbsquE4eF4dnhLT6jHsRzL5M6kNuPhjKuEjcD3uajM
Y0jsKG8bHABPcckVrM5zSc1kXREQak4X+gLHB5t5jVNA3WObe/aqv2zXlLaikrdwXBtyjJ8TZEW1
8gJ9LLP3V65iwfFafPgZ5oMYPM1IQ6YEF9Tq3p/yCWpdG/nqehpVtmdfQTvW41ZJHttHaHnjbfDh
YgCABgtnP+x4/XSJjWksHno9MCN01tPtOKJv0rs/ZLkNIWLZFCyMgoJcK+Fw1HELmgDkbgTnG0zP
HYKlSgHyOtMk36TaJnTldEWFV4QsSg8NVdUbvvC2UQjnI2ExB9IblryRLbK2EbRsGNxlrt2d0oCS
ip9VqQFxZGNvsIWqDbG18P9H2hWWrgdR84gTqkq/8Hm9Sd6UtJBL2WUqnQKVuwXJsWhzEA2qh1Vq
8PSh580h6U1Gc7ogvXUYSytjr9fqp6aOBJJxuCG7wl8/6nh8fLR7YqcBJZy4JbopunyuRlyuAtYL
yc4ZGP7XHdJQ4GBeugx4JQbCoPDGzaxvVhiSDroI5hYQnuXnuceqIEWpZvGINJfXK8Yn+9tPI7Kd
hFjTYHIJkm5SWm7R5EItWBaKndSDJa87/lXCJ1nzHteBwFDFJs+I0jVVQLklgszLhEMHGg4gklIh
Hs8SMan54Ro3GZYJbvMerhJkcaBiWxsCl03KMAGcLwhL07gFcMv0KDLxt89oKOdZDXFonc1T9wb+
V1e9/+FXianiIder1xwbz87F1Ujri782a7PYIO8m3eqlVIQdslRK+DXHCOtiS02MhoqyNgnxeXdO
8mbiSd1FVRmBhSSjzL2I3KXGO4QpI66zt5yR2y2lImu2yNnzOk4DZJG4qCVd9M9PTsCiiQ4feTR7
VeaVMpig6F3347d2JhxD7ElQyOl+mRivZAggZigCFDTl+G6WWYrJcIlknrKxPvB7KaL172TYgTBr
lpfvOgm7r5EK61MaayVX6M163tpQ0uetMcSH571frsYAmsmLIwMx8wMoIChhpM6A11VHizoNuhzM
ytmbqYN7N0P7eUmXGXB9MfVe9gSg8kqnkhsBjriOtQq3vljauEVuPpTEhnmLPMb1YoRqPYjfr3t/
9AFhMADkYzQuf1SlRArp97LZCawjQ1cc5Ix+PTUaO1HKNOi7cL+gq5ppMhWAAl3+qN9Jqlmq3YVN
Ut/S7lG7whC3d1S/a3dDoP2gBvRcSiygbqxDImttte7YRiRRv5fReEEwmNY4sPyjHDmcZgIYQGx/
/KOpSlnWuNjGAiPQKGUjzS7ml7TUd3M0GYuKRKJj0vDcE3u4bwl5sdPBa5d89eoQy+asuVB61/il
f8FVtbxQSc67YO7cUFmkNlTgIu6yGQx9PAbYhz359IRs01EEI/mcniXynWNxqyEh9KmXrlYH7VBD
KZ1v/DLiu7osV0+EqSvoVAtLAu4pcCPXz+qYJVyyf+z+dz/dh962Ipx8+G3ZJbpV480DwTxq/GED
f6mXk4aTwoF//vncicdz87H2DWOMOWcGCGRwA3gxossUmbJPeEcODiNh5Wo62QZpK1xF9n2z6+eh
WH1Q39S+KoDykbmnt2azD0NUNP99aH+0KbKuKuL3jY80viU9rAeW8c05Y6eZQ1Wua/LF9/AdbhuT
5I5ZlQiXa0EQjFQORXEdJUDEsSsfCbL/rfzyHUvN4Xk2Fpt0xOx67sa7R7JVQfpqIkRCYqcXrPCN
hpSoSKTCILar4WKzUNFJw0mlHL5SiXovc6emew3xby93R9vRh0m8/N6B6weWQtUJRSpimODGpvZR
y9YaNpSvQbMsRxCMFv4ERtO+/4vTkHkFbw7famUzgVOfC+KsqRB+Ppjp18mX5Cw91PxkbBHAk+cE
UuupIv04qPPLS6zYyjJyvbvd5ck/iMAoWqa63HslEKx3tsvAcIoZplk6ACP+AHGUOEiioIYBbmzg
ATD7rPd1Q9z3m5Gx6gO1m9mT1H9hiXfbDgCCK6DvTvZiQ7teAR8jwAThuAWf31b+BCGH4w7efqMu
79oZCX77GF36bP8oDAErZ7mFSAHjaAWwuD0RtHA8e+sa3pB6Uet7dNkCmuUMVlNGXfA5sPz0U34V
jOP8tP0kHNLlrf0hCqbYHKQdMjFYg6NDFsyTYQK8g6hlREEHVjM33AQODVXc5yBkeoOz2x3iHnwe
3WSQpAQIiqNVlt3ITjdwKNOJLXzP1GohlQ6Y7AQ+HklcXYCGzOurjM+sQLp+UtLitPSinf03wHrj
t8pSXwriqhVhuzoXlC4ZPLhAkGl6a82sEcmAQ/DqEvxeKpJMk6hacCYr627d/3I1yDRKx3FwbKlD
yjgv/Lz/FX5XO9Vs/1yXL16e/UIeb0EuXMIF5AIAuC0+tGhsXIQf3lpkz3H8Ynt4P2QBEIfFTQ6z
4TzXF0mtIIjBcBoeqTUyvvqiDE6bF6keYnbk1tH3XWIkZRfDWHaVsM0P5lA/xN2PUtriyMtCDEaO
WBiHHppzFqxY/QEMYC5i3YBXsNB5iZqZ8Eq+RfGLC0L76iADdEhSnUduHjIVzla2zEruxeEwP9Qd
T3HPPDzUiC94lm6zoc3ut2rYxPjfmRg50h86NqCYnXmuKHyRRHY2XfXEG1DGvOCyrJsJbaFvgzlU
y5v7iviAB+vZ7ABCiXFCP6aG+bq37O5uct4x7ed3J0CsqsqmOoW1tMGLnAgtd71N66IszH/6Tk2i
p9hPnCRbqpXhEFQT03PbJP50kBBorqbSERlgBqUGGAgS+go2rCI0KHgRWeiEqxH4+Oup9+JseWDK
JknSOQZwp4ulFvyybmh+4mW9PXpcLP0F5L8dcfoXpYoeITKdiJXIaiV2kQgnM8XdN0LHAkKI3dMt
SShAulyjHatVh09mqS/c2+M0MoJw/f3q+m9jwwZaQGHkF/U8zH0ihERcr8d/gs3tiVzGw9SYF2+P
4p42MVp/g+K9r5Kn3JbFtFMxJ4OMZZM/bWvPBMqTKGqdnN2p1zl2fz+mKeN5oW2OBwLZFjm66jda
mAP2J5XRUCGRU1SFH1AS1WgnIWMn7feOHns0LR8o83cIkO03o9FwkTTW4YcHbrpl7mQZ/DSCmSEM
GMnPxwOLyI4CGkxr8hpvLQqEtThIcGqQYYdR3pCIRPMUqbOz63Jrqw4uov0hTNuP1AUCzH0DEUj2
DZn9SrKSKQ6pdcIB2M/OWBk1qAKvTBMfog57wu3+nAVIjzF40wptDOzYRDuyeSNJ1aoMGO1FgENF
5PsWHpqEmVOTEhnotZGndctoM/1JjSlKtTnx6bApqijz8bvhJvpbBn1ov6df0F4JA3ScD4585Fry
cF5C2oLdWW0qRChtqIPkW6BuwpxXpnPcuupLYButUX2f+UH/fBVvb9TnBG+G13D8Zc1KADHno5ps
SSww9hWU+9MRlngCTNJW2CgAF2F1v7rWjI15gTOCEx4f/cm7T08Ao7XHGMEVGivoHJDLJXn+5tKP
JNtspDdvug0/uqIrtNLBEH50YtlA+Rz/WfUUbaw0fZ2zpWawjm+vKSPEqsrf4FiSb51AFNUxq67Q
cWhvBOee65Ck420cJuyim74dZF+39o+asKlBot5CQ4p5GYIXvkJGmHDvTY5EHNNPILhlUkbaQnaF
MpXNm1BjNcTwexKGgsWyPKJPHlp7RgRovpqBZTDmTXWN5ZKXaiEB1wztf9lYWd+S5v9EVrSf5f7/
IP9v3WGEKvak1yI0RBXE9hBUYt0XPVqclt9sCeFCVHSMvb7Ep7m/Y4Mjt6b+PB/l9kwXs9p1dx6z
Xebgy7COzAGeuqXGZ/ZSxt/ME62w5lXTtKZo8I/dAq4+cZtMaqMubsXKn5/J/2dCvhPJamXB7S09
cR8t+df7Ac10DWqJ8ZYi6Y+MmwKQGD24N6FFMiY4ciPD7g0jJZMX/N02vWtHEzm5YVKi2i0veOqs
1Ts2Gzm6iOamho/twbSYwzsJ+8b15YcVBw+GvAFilS1zwXFobs0r0wyVg/1RjshJ0pz+YzrmJdPx
4fnqABwJLYB8iZVzLHEeAB39T0R/72yY7KOwq58t+cRNYcQKPPwHEWHcXU5oY/8H63cvu120BNu+
y0NWDb0cv+ZaCqpUiyOmFEBZa9nQW+xwZ0ymF46W/quTKKcGY9OXlOVuCcW4TBSXb9hqEziBCp+c
HptWGTLxPZLDKOD+L8polW/j482Gp9t3pLgN39xIkP79PkLLs0hJR23xJj1x7HUNxemP2XGu6NWS
nyk8P2DsZOqK0TOqN5SN+JPyp7R28ngG271CCiEKRthKHwzeOYLPCSB0otfn5+Mv3Rl+5hPnBwnL
VCwaGraM3SnMcgPBt02v44iCZqm80zg/zdC0ZykOrlD3WPeDWVOiWik7AkVtO23Ry6IrZKisK0uI
DveiI31pcMMQNlMEsoZuODZazhsFF9SCWIo7U/D7rz5QeIboweexqBeybS6nIBCd6djzSn6mZ1JB
qN5RM+wtQG4WwgXHVqPpAqzpoC2w9/MCiEfvNSciQu3dsRs47ICT9WBc6oF9xrKguXA8wU39uogu
Hkh0jLsEQmyqx6zH5ONQLINL4zzRVdIdc5owDI08Ex9wlY83r80gxvdU7qZ1HDD2uPmNy4EZtUbb
ooiHn/Gya/ql27axN007ARcUlKzWWnan/h/Fkt29n/iGuCiUi8N8edyLu9gKi7PlKDch+U21xMPo
vxkCaEtuqVoR1HvSqvjdfd9cqcnTzbGvuCgZxDiMyKyUlaVGDFh1B+lwyQ3SlKV19wAStFbiaLZ1
NmbXTcqPAEkVbfdRB7RDlray0BgLnKEbaXPvJ97SyQTuu8x2g4/4ok8/KZLydA5PQXvYe2gvoAY8
k9i57/hetKnrc/4eFTcFsct8w1RoZeSAUgXKf3wdOl2kY0uv7safmSGszxaq0rZ1wDBris/WEgmX
yBASaDRn0jzIjssQB4lQ6h2+FwKTb4fpbxlWY4iY61oG8R0gOIm3fjfu0e0SWp+dxurdAzqxPLFk
vT1twxm+hVpvhBHxdlO97uI+evDRZ1IriCKUVj7ReRbOe1xc6uau1EbN2eJs+1jitOxW5k+tqumL
2hcEnMV8zLbgAIcxicCka5OcY1LTRO3Y4SonJbjJs2D24WdX9ZsKFb2c3ulR1wDOMFCJm7sj0zVy
+uvmIX9WptlXwBPbnEi1+NAAI9Q3tj9uQEdLAJVR3RJEUnaeHA1rcF1HWkq9DtTLl/dIhk/LP6WD
HtGW4iqipt/GSQ/F9kBz5byDE1y7zTPrvd9STpa8S5Mxb01UylQLhTqC38ndRUsJweCwE72ovTOP
ER/BKB4uz+FtRewbxzkeUmaTwJd7O/8GL4vyrbDAksxYhC/Mvrcin3aWqARc+qzDeKxMUvu49IGv
NtUZWN2W8I8/VyeaJWFmEq2ZPbRQyAHr/WyDVYfRgPHLKcZZRBmp1pdlcjNKyq1CgO1Imn4KyRR1
4AvqSSp2Wi+PiO+vTkvVtbgJKRtQXlNVuERuFM6t0Fw0AXC08q6o39Uq6wtJtyVv3vK2/8G08m2N
lcSWAQlWynXICnyeQCIee9BIuZW2TU9tCe/D8sFVTZqgZZghkPDOXn/f7/DOXIQlogVNGNmubnNa
YpPIhnZ7Z/zWYTg4GFAl5gCwm8sTHPjdLIAV/dsEWzK5V+H7aqHBZWl2nxtJ09DS0zWYVAfKCWEo
VMctbvkCDy31IMYnVl5V0TwAKWb3nkMK+yFEpwM4uOkMMCF/L+gP6XeLCW4vQOOkEV9dZp6eC9Sj
ezwpk5uv5ADvdpVMOjr7icE+hHdhIiX/IK/kruGhqMzO/TWezOmEDwRc9g88YlfR3M3wWI9pvtIm
0jnp+mX2gevUyeQOgFY+/QtRrDdg+G8qNqdncaQoSj1ARcTQOyPs+Y1gxJjpVsqt3A9Uj36SKuwY
Gbewotgp4q4EPDVOtPJGUg57RDrbAihGpK55dKwLz2rPVWf/UbFXlrCmE1WckLq5xv6cxWYvFOUs
3d2WH35DZIQ5wP4+u+EFy0FURP8xxFf7xnSEmNTqP5+BdryvHDtDYvmZkQBsvqusXkJsr58PRcs8
ilroCK0ZwMf3uIuR9TmMwcE9hVq5CnjOk4NwW5Sm576quFmN6RLo8AZsrLmTd1un5Pltpp1y2q61
lgtBMBRT+1UNJ0sgPllHfNoZLSZ/yWMDgminGMFD3eoI0BMdpddPvRmoB0WPMi69nsek27ArPs9h
7H3/O0j2YEgpQ35nZUm8EkVS6j0myhldkumpnD3SI79d+DZfAty/czgrhzSxVpy3/jw0fG9OFTVz
2OoPWXW5OeEKTEnRgYTIx065aeSYYZ6D2eAv+CUgI4WdwQ2ZRwmpSUlT6a4yJqG79YLRHlLw/7Pr
/lIP2QGw42DPvUQIs678TQH+6GW5lzj+LLbw0Qzthz8Hwl1ZdI/OcSAis8fnPVkn006vZ9OzGM8M
NCg3E0BZfuLBXDSl+oTQQaTPkRwmbsjXL0MA1Ht30y1CuCjc0sEF1iPD9pVXlYIiFAEasbPMJ0JW
hwDxPJ3g2cvIzmR8wMesNPrpth3B/HiirtYnt1lhjRB7Agl1hol1DoCIHvRdx4utpJS1kYlKg41n
vv9zIrcaDE4lj9EONCqrYySZyjxTSnyvgev/1h5TB8J746qRK+E7WUkMFd0LR4f3ylna4M7dl1UQ
PxlYP5+yqF6S8PrjEqCD/3AOJmNTsVbpEOG4yX4zPJ/zL4kJM3CcDgvK849l0rH0N43w9fikj0Gu
WGgXASadC9zfLIfR2ADQlZ6NTv7pQpGIJsNf0xO33efapvBJm+GLvfNIg0wDNnYUQ924AmfhL2yd
EQ7ut1FzX6dxfOd2fHpbYzY7mnK+7pv2ubvD10px1TPVPnN+lGXgxSyGsbF+wgMdWXC9VH0GLXVd
rQSWyybA/P9zORbvSE1gmvq1ah0AaIuWrcdOR6GU2tKpHyRgFAs+FaluPL2/Lup9sUnzmAf1yD4o
529zz/wbja9Jp9/HssSdCubEbUQ1U3kT2GisBTOrlWe69ERpAAU2/5wd97Bru3OhuJCT5+GjN/Yj
2EbGyu3UfDaPCVSEeqXtGT2RwOBGa0vpCzRtY+tjlpRkuYOnkb1GOtM5xd97kcB6yYjnVzH488AD
iXTPNcBi2x6xLlOY2juWa96YdDSO7if+PfVGHBytXWl5vLSyvJI7J97nfPLxqcLlyRQ7ekqF4y8v
3XU/FafOlqxIUrB1p2ottdK4RJTxHIY9c/RWYaowga3euh09Uj/FSsOqKbCTDupiMFksoBD6UkQJ
sFXN+UpNhUQ+6//Bs0KV4TY7CDMeHsdKOWYSKV0vid19CG3wep/8z3WpUepj9vozgA7TQ4Zt/dFt
9RoJPWut7EvYv8I8n2VtYJq7w45Vi9fMYklvndBPRWW52V1fPXv4XO43MpLJYqWHXlixphw/44Mv
SdRo4xpbuEQWR/qbtufInKTsrEkd3iHhGvwzH4gGVP1vEmlkRlNYULtWVYD2me4qQFpJfY5L5Alz
j6jRVzltLWmtCova+fxThHlpAL5X+jcrCrlcBFFEU1LIzeFvUjk5581hGjGeEJyAeREnOyTCbzAC
T7J2fydXJMA55XajwYPT77pInwYHSI6osacq7rgaq67qaakLxSuAGXkT3Zwr47b5QnV/n+fV6DUJ
4SwO/WY0GChJE0GfhaDH40SUG4EelWqlQjdzgcuKUty3wJphcuAx1O5psakjEKM4BA7pBhkYC0L1
PJ+h1v3RkHIkYQrzPRHv2Ssgc6Q4ieESxncfdmkeqyJuDRn5RWRvZIGZEuqwNS/lkZQ+o8bgbRjD
eTBeGV4Ju5HOCCwyyqWn+yWtCP6CrhvzTBwDc4xeuN89Yb3KHyeL2C6yFhVSrnMpN0PSuDQthRxK
g7Ew8ohtMaOi370gpdXX0X3lb4JhvUv54LQcxb1aQed+GzkEl0b0I6SqBhFCfZRwbWJNyLcbt48G
DpCrhHwSNaK55FPiHGDSIniWDCnonYMJGsj62g9BKc4mVbHtB017x+CjhtauoWFM01nV5JIm79O/
3MlPGf96SV5TqDv3ruwen11fhHeUL2ZoeDad7vAXy1dPYc9dr7JPMEJb1CWCX0W5ci8brOHYml6j
Vnuu9pW6quqpKHhmIWV24BwDwdhZF6WV1O/pJoZtMmXxp6M3gf4rWnVxopxXUFjCH4pkquU4t3gk
vtSEPizMbCvuL4lLluJcSya9eoLPydnu/OUAn9Fki0o9079WBryiNsh89WC0L3alTLQhfH4M4SGY
ypwQ5WOf+eOo1GsMjLI9evzR20NuMcSH+9onDLAbXDtUx3yKMklWHFKOrBjXkQ9xoXGbg4/KodBQ
0qSdDtC8kB9lfhQhhsSfWVUDCKqG/UMhAb1ltDmQKoLa7x/8dQCSRSrERXzTbDJSHvYdspLUVqgz
+GcSXpFruWtX0hFf1CZeMmy3H3C3QBHmDHqK4SAUzmddt6Cv2pnPYyIhBF0sUz7LsXjGUTolXcx9
NBo5GCePo1U1IRiiz2zssAAeWvyDoP3LYkY/jmVO73yb5jRJAGLfLRIk8WnmcYXicHqnbhNIub84
quNbYTw1hgSBPFXsscJeYfx1NX03DMn7fHaBHRNmDRsciDR1PqjhaGJlG65WpMu/zTj/ERFG/WSn
a4RYaHp1/jxZvHBZlmgCFuE/doDv4rusvUby4eBp24BjvoVAhmMKdIKpwesrYdZqulMsRPBTt9BC
BMo0AcY+dvGhBsLNi0z/AOsEdE85LTIm6ubqvcceyAln5QAhZSTqKveZXeoSRl8CVXgWLT2LFDtg
tjQEs3W0o0F8YqHR4Ph8IoBQ9UgziF3Vs9olfe20Dc//0djoPTke9ib324AAtPKmJZp2+2XQQtap
cyaa8StD987t6UVytBTxbIs/A/apfMBn7NDdhRC1qr/BA1mVACyEueckdw+ah6PUF2UohKn77ver
QlJ87VxH9YIjJ0xeHBx4BAOYuFsbs4yiwZWP7z6qJOWnJPQdIN18k0HgzuXJPeHX6yjtah3P2Z1B
BEEmHR73U2xweypEw3d+wZ16px6KKGF1p7BEdGpqyoRVK6lnBUo534ENySgsBMHR+Ya70z+ROJfb
wHeTckkH0gaLj91D64r3AaV8srgIq+Js+ipD5M157yyjvtLLbPBhs0z6Ah1DhvT8/s5TKWKWlcdj
q5Tg9QyymAJQt3aCYPYqx5JYzd6rYVVP9c2N4NTg4SyO3At+NI8ZOe12kcewr7ApTvGh4ySuwrLw
OjKKhL3BR0RCXa871yn4X9/i5Ab/JLSyF1XDszPmUlhjS5nx98yqYUDEbqDBY8S+ST4aBGvbSRBG
qWKatnIZgCwvk1NtJ6KFSFapfRKpcmW6M+QTwLc+nVzMCpMtWKAkMdAHM0BHrqHKe/7VUNgYa61j
n42LhSIUZVlh0zkUOUuvPJKFbWtSsOZdaG7ei0EgQ/nv5eFPB7RL2n1XJWDXy7iQSz6q5hF3Fh2T
oxNeY7amHkeGf1qWXFac8pRSH88HLodrQsvPyx2TludZ+hLmbrTzVphYU4jg6qUvDbY11ZXtlEbR
lC08ej8mJ9LRH8mGbJVcm0VDn6HvwvMRyOLFM0N5qiaZ+cMEgTveScwvBhRHvS+cPsCS9un3SUNc
cIFq7jwBUp82CcROVHAL+2PwKaVMrEtXcScWtfwRVqGCkHekP44Sb3JJgjlBnze6DkjR+Fve6ywA
OO7iy3Swr1h7GCAKnlFj7S77I1C+QPEzTSSYshjcgwUjmn/95dznLo1bY4J9u945N7kWk56Bf4sQ
irey2HF8azebDtOoyM1oitAGPRbKI90CjeDIqxbVTAAJ7ffSiZCm8+26LaOLiois3vOUnLWUK38Y
Ghss7POwKwkAL4lD+EhcgNQtcGRBuey9talV6c9oovaQKMXO0laRFFX+Z5HaymN0UiAuOjnCwOoT
pFRhk9dirya/hEUYUAknFtRnn9H7kg7jBZ4tszI5CNEQGZIPFzfHHw4gTjga9bjVURuf2XmmwNkH
0CB9ef8blIkNFAy2zZkuXhQOsIHR06Wf5N+wa7+zP3MpKP7C+3YlLD0rjVS14Unr+JOzofarq1Mi
mvH3mP23QONDVqgd1qlrRBw1k0E6X1V7JF0ek5wnFLK10sY98BWg2zWI2JAjqXI0bqIW/+vn0Jed
Mfa+ec5iVLSeDaYKxOBSakLh54J6dcYEPK8ak3Z55WRkQXVM2zIfe9P/k/4jZEXw/shO0xoVVu/M
3JAvkfAv7uK0ZpPMKgGf2MLHRL+TVsyQ8SfpjCB8S0gQ5bitPCdMhb4bvpVbfUqKCRN823aGffyD
oDHnyJqotWseUrcfWy8XDmDnV0+LdZ40DsdnG/Y5QpYmapWgTKXwsAFqpWh4FJYtK2EU4rabfFYR
Ncaa/DYfZD97/ObDZDrqKK6D5Y5e2rFb5u/lDnJUi1Xkzhk98FcdKycFRzgoY8hDkfB94EUd9URd
SqnJixhwMvjrMSEBjx/vatUcZrvs6Z90QiqgmvbnOGTHbl1jy8VmC65LdoeIZcP4LajmzKYvIwgB
2RPZ7TQ/3sEUhDgLuG5n9FbVSs20zZ7zLcrIZlxeIgd15nihXcDTJq1vXAHUrrGqDN6CLp4UI3yd
0hecDA8k7eW/fb/8CsPdOR3i2sFTm9R8NCqM3vG1wdAkQnYT7GCsjm8D/hMpCRnWpcoOJ/vTrCED
R9jkb/9iiRplMsUIvsxjTVvn55DpKQypyNjMLRqHBcR65X0UVtmeutOeKu+VumgwGSZSAq40+jXU
SAIS/HIyCO6QpEK61PXGBAsQsrlz5ON6XukyezZfSfqFWGmOKHTuSgw9bHPpkYQoY6P6XPd47/FE
PBWWSw+Wc6OPTDTLypPeOM1mnFPSMVamXlH3xuhzwJRzARmb4qPJwL+jCGwCGSDdOPG9Cv1PzS4J
/+jNgKoad0RWtvb612rNz+8e6pABZnKniIqEU4O3BTZS+e1YT5+oykus5rRm7fE7hE4eG6alLKsT
bQN+fVPu18X8+lMfZZQgHXiia8+4R6t+tzppW3xiXN1E2JILdyLJ4uvfAauKdIfz7EqBslB8OGzb
HnbOPjOBjpSSCfEVjWGib6EosDa4Jon/U0IcjtaXYlptlQJ1zLRjEyjXAlTjO1jx1Z6rEz/vXyI9
7DRBoHpPQzffj9jA9hjbwGjVmt8X9TPELLxXzOEjCutSg60uFNL2GOADgxOmjdjQqdeVu+rYkfzg
n7iDjQcQuQe/HImxkjaoIcHq5JTRFMucyQxvHATvu5VNY7ZuzfrW99mLp/6yNwXKJlmP5kIHT01L
dXyLxspcZKRd9J2iJGuwcIhgoFCxAkvR3dWPwzwiDG82TmvcKbWRWDMYAIJru3z8d0zZZEUPXS16
+J5mNaqy3HHZEAIG3gmD4eHmtVu95H0ty1TGyD1egZnYCtV4xmEsfpiqNJO6I4L8vVIAi/P7+i6H
+XvWr9UCR19UwAA2Qyx0HcUoonPGUDvd2gclZeOu4uCB/y6vdqO0TQMIYgU/7DqU9tYxHEbGv6de
+d3gbJXxuedE7qdKC/OXDs223jBMoaJ4wOPeEVzHU/QPNOX7sGx1PPHkq9nCUoIBhekxQrS8V9Iz
2G/dV5RDQLegqAluLtuuU0DDTEITjh9CaKDFEOw/DsOm3qyTq3Q78FcsHXp+AKxAZL4JQCG7FvSz
siS/UhdQrVdE05xgrXTjc+6LKkI3AK0y+/tQGFOUhj0FPmwQEQQ67cPqHb9hyIxjrXGfN0Rtms9+
Kw1n5BkuepT2WepH3HDBlGEdBDxuYhzfA4dbh5ijh+/nrQB403bi3XvfqWZ3UvZGttVlSk5/htwV
TqYjxjHNpIs2FYPajBZlrzDscmjnayxe3Jeg2NFV39HAla3z571eLQRI4dytdjcjnDNNyDeMgJ0L
xGBiTGjEvdeao7xt29ddn/Sgze6c7/F4L7Mrwprc+oh0GGPt92SVmIdzueg0cXpeLpvh/1F7KbfC
1Zya2ZKmx5d+6pdo1X4dPAhsHC40fRZHj/qwUjZByq7L0bC2XpHSwOeWPX6SNTPk0OtihKr/RX9i
HcgAgjzglc5JDga1pl23iS0nEBMrQkbGvqlaKckkpDQi6Q8GHhiOhLIImC4iK0BaMa63p8OFsUTB
DOc6t1OKtrEWitquPRtZWZ1ZT/CUtuy9U3/Q5sdFsWYd5rrvauzN/LSVUhsFP1z80ZP2l58DV1Nd
bN+dThwZWLllf4Gf+KfxV4gICTL9Ca28lLUpitF2Bw3GcRJGFAlYv6Zaq5E7daTcC9yMlJohhq6H
zJr7uun/ulhl8jlLO97tk4mV+zEWfkhvra7ATbvjUWabtpPUIl6iDB4MJ9n6RgaI9+fv8mqZjkiG
VyPu2Gik2/C8zzqE7axWxuKGtvRvXnV0ufVFtHED2r32otIqNGIKdNTbMVtlIQBb5yamB5TGYKt6
undN3GLDirR6Cl42Zp8+e5ar0ICt8wTd1M+En1jkHZIw15neo0xVMPMMMIPbw/Jbog0SbLfIDipj
/jJ9ZDWADZJSLTWQUPZynb7dwulm94y8hwJOfZFAQLlYyLnP7iIGaYcrvkmqsDyRn8DwbiPHwSBK
XZOnJIrsohPM2be4tm1KZPu+UUsJ3w0jBDZ+jrDvq4GFQvWi11QtEMt6OWofwwsBdRcjWXgloZgV
+pj8zaHDQESdqiDtxI46FGxRDehFJaa8laS0p8O+INk49m1+NMsg3e6PzSH9fs4tCtFCpsrZpRmG
1zgXyMyMVVBt6aa+iyb/+MNEWosvtCVcXC0zgqC80ycKJs5jgVFEUi4JKcL8URLmYlMRFq4aXHDg
l+dz3ML+8CBwZ8YifVl9nMo5QraTrly7e8Q/7tZhRUK7CTqkUrUsDMbA6SGlHxzm8VqrpXW0SJTn
nfBXukHa+6DKg7Id2UJrVs1trt3TxedvmajvenCry54s1UlokHLMZNwWeJBWDMDJN0HXHgq5KSQl
L1pemXKLj2pxyV6ikeezuRwAMEv3ZFPZjYTT9CKwTr/zLMe+QkynoLTQ1jUI8jQkq2EFfS0berp5
z/E3S4U9EpM+GexpfDzFFuNX/VPESSDI7bZgqQer5KwjrXk1N89U7CBqMNeeCUz9TN4rhsV6iR3Z
X5cfv25UW5gHkQsFnT792XfRu9rkRav/OurGomZtJxfKm+2XRiK+a6ObmIWWwV+wkNfmgUoCyx4H
GxB+B2F2iEi4CpEGpPJ3vEnEb7vPTDzKcXsYdPkcpNLCbJls7ajTh85v905WnicQAdW3v66I8cGW
2U4QGc2M/8trq6rW7b1PilJeK0hb417Efy9qkt9vaolRsFGB+i/gh+SwpAXOZYUKj/LElJ7COkw7
C9nam6Wd3nkCcGadZKw6Zrpr1Dv3AW35Xo5kZ0IDa77NSLyh7bHVNT7jCWkWsTfSbOBRyBzXIIBz
7Ntwqfw/TZ3ZHpeBuMR5Ws6h1D6Lm151cK8zmxyfpuyzdFzekCo/p1MV+sEMO8wdeUEV60Jvsjv1
EIeJLj51277NBxJxsvesb18x7QlmZns5zqLF0xUxj3HLRo8K/NLKBFmEQbNtwZyYemXGA4bzUlH/
Fy5efFkOiCOsPW2w6ThMA81f7l2hQq7DEajiLl+VWVDkbvC2TuY91+vREJnusvOQmDoLW3tES0JG
XQ+/jtKjEClOTZ4ErtibZmntNRrUDT9kZQ6dzZh+M+BGzEQoMs98OTgoKILmTTMyj1GTkGdj2QTg
xGwjiL88/Ho1i4V4QQ/oIfvB3GueZU8dQEtWdBm7kVOvc8DEwYDUXFIN9YQ5Ev0kpxG6aW/Z/Yu0
tMsI2ec29HpPD05rOqSYicENXX3a2uRfxcP3VHG7jRwWjAzarPS5ubC8OCEOI/kuPGVaFkoVNaL2
2Q2m5y3cGLt5iX2rVfAFMYRQCxKBRB9d7ECv6YlolQWgyPYrtK1UTLdkQYYk4EZWYzL9w4j+I2Ol
2W0FkyvDDya2J9hAVkuM6Dc1iueblZg7oTPGbPCP022ulzabmZNE/AAzY5S5VKvmdlQu7SIJdvGb
KZROj07WOGFBYlMK+nMe2nnPIdRNVSyrOrMQC7WbOnH8NZAO5mGJ23NODhzBdrkSmA0c3KGWDj+D
aWN6m+FCUuYoFHDx/0PAYZsdww7WKKK0AJa6B1GtjkOYfeX1JFd6ZUpN5SPLWxRxGVm0iEZ2KPsE
adaMfgkte6zwmo+lGGnNMtcmWNRMis9AnWYY1ds0GmdKC1q7RsUF3pGLWDSaYn10u84LzSlGbO4n
UzbHGoq4pyfDg0GhrTcuwNSeHP7orVr9I0Owlui87k+wjRmpiO4TmMKv59nDamO5PsC0LTCoWQF5
YH1Xjiub64xy6BJxZm3d7vlJti29D+jZkFu2jxfWqac+uDgu9eXD9N0K1Usy761ajjrdsCWZjNCO
iqHDTz1c6nARpFPxCpZQhZ2JyCozESy2ixvlVaf2eQwqAMvdsu8H9cTfGMNaqYia4q2dHEhFl9Ut
92+bxPmqR2YQXryPTZ5uEcmT6UC07eAJhrVLusion7ngF8SHvhIi/i4dySzA1UpU/83SYeTrOEdy
dJ4nu8jYMAxmcpJfNH4WspByO8EtKnnYErbEpJe8fud+pPAhx9VEpQPf5u+d3QPFvaeaMyTkIiD3
DUQLQHwLzFqVOjCQQNP/HWZKM66+aMfsPnVH1IMb4tXlfxGdhkGMqhenq1ba6rxumEntcVRPgxnb
ZBNQnp6JGcf9G+jcvu58UC+4DoaIWI9RoqXgCDWVlBpVbWYuc8+1GUJw4dNM44gxV6bUQWrytOX3
er2M1fxXVFjLv8VOLv9/tMT7VmUbl+kVmO5s6uQPqIM9ubWpMJzhSA5upQ2PNomH0u6Elizbhidu
BwHEfEfbLQwtCiBzWd7I0OdIrKe0w1GBxjvjh3850NOXg44JSY50QH7ZoAKK7BnJrn6vkWLq4GVY
AH/RnEen7Cn1Y2oABqQPa0aeKzmZVGgD/QEk+M4be4xhWVV1eBUeCauK1usm9mD/ZaKUDN3iwy8I
ldH/nhEyPc6Hzb5WuQbKQMnyYKf7tDEqu4SGx5g4hs5jYTIduECjcYYeVkqUAXZEhs25pDHLmYqQ
c4yG61dUQOIQBl2SK4KDZHYpBrZZaXtfbu2ROuIyf6SLFi+Ugwmw/7kjwGhCGMjuduYUhVKhDAwX
zUZdluRKlv8Eh3lYFcXfDHmT1llXJ+u+/XroaRMUgf8uYXc5bJ274/qnZj3wVKrVgrEGsSCi4ucy
fNF5N8A2W9Qp/ilq/RETmGjQ/6iBmQbDEUwc+4Fy6dMkJkUUpCrM4q6rTUuSKHFwZ7xp2n4tlSvf
3wQ6xL1UsNRbIGNbOeZv3Pa49pvsDZi2Ih4VJwGEYBeNtwVaYn8VodcT3rtPt2LZjRe6IJ+VaiJc
lt9WInaUKfcRu8932eUHsKqpIiBFYL8ItJGJzpPCE2M0oROJw9PzavfjuR4D81R26EkvVbYiqxv5
I7V2upbXsNsivhioiamZLDbKrNNa5HqFidxYEOjxVVKax7Ibqdoj5lZRXRyLiWw32SnswZEYb32j
GOBlP64Gbpujp/Iy5WlDTnDWQYa5IiJ36ESixwHYqEHVb98DuZJLiBeyTq1a9kity2gLJVTMJe/4
n2y4cPET/Y7+zpleuQA/N00bBW9uPvuOB3cxPeGiDOn8fHFtING1Tr6emPD44RMIbjvjBlMwrJqS
MKRCl/Ofl31ECkYwtvU+QrmHew76BzKZevysDvjpl7/qIAnbvP8kKmeBLVZPH9cC3Tl38d5l7/N+
mIyu56qvXX0PCFbWsw19llO7hpn0T43Cciu6JVBBryhI+3S5aFoCah6W9MtJgVW9GpQfFDGsZpEp
5xnSEjocorH4ojr777O1ULFhexMyN/OBIunn5vDFeAzMd6N449GnR4E4YplRC1YsOEwRqhZ6fAcy
KwlBBV2F8g9YDsXz1enhNy6uRLP5vTTc2xJq8xyX6/d5UvHkAXEnI2W7wVoS2vzZJ8pvpq8W00ag
PV5x7SrupChZd/TyyTKqMuxj2ZbAzTbaYnwWyodNla153xWvd5Unp/I9FoOKncvEJZshsIwRFGGQ
RdMG2STCAqkYj/jdU72ZBvTc4rI1kF5HVsO15RYkzpV/ws6tOMwA4uO2hcjw2gQ1iWvHerRdZLUR
t8JCxooOsf7y97SvWntloDBWbIlBHto1mwdOgppzUWqwqlDeBE2iKRL8I3EbI5JSORMMZ+cbtb2b
fN4+wUhPYzepDilW02i+jlROwyPfl2KTgxDALO/Il95gU6whJ88bgxHPGYBhYqfIshxSL80sfUSJ
12zcopiY7o91j5kKvOOU8O6ruFTIcbLQHEWXpd5SWpbXxmc5XoFzyVF0Xq4GPyXEO+tPxn1ZMBj6
j36kVmNYo/dVIv+6E/OP/Nx/Z5vRppRvZrFOA9fg8JB+BxABJVr8vOlYH9Np5u5i00DOWhxWfuPd
NuQGGaXaDCG4CoKCeGhLFqQJUR4Wk0aF0Gvf16psOMLmYPCJVR7SdUHYZptpquHCHfX8Py+g2Ygz
TaqdenJx/qyaI8IT3EAH7ZcXb+Gd+NGj5OtnuFWvllMbWdkeZbPMM7TM/3QD4JOG8s4oQfQrsBxr
B3mdqWSRN0kRsvwBFFg8V9RqlNPtyw2ExT1u0RAY6FBd8Ey4nLjyUIjHhBSxUKyDCPSAMG5wQ3B7
mowJ9LL/0HzCHkD0tpabFrbrE/P6J5Pyoq2jdALwAz3FDkMn/vkz15FGLGeoUl/trRS4PCIuGmal
otjBuW949/W6po73JIUCZvnk3KvnfJaCac3iYdpOjbCEP6iq0sikcBmdoO0I12pLd1qplHo6t3wt
jEjvRFoIhuLqyO2NqcvDj1FASM3251f86OLzoc2+zI2QHS9q63yclJvyon2DinlUWaYvJfBYQl60
IrP89y4v2sMtiSZIt73TRDVvQQD8CKHZb9NgW3YLk96YgMfWTqagAHP2UNv5KBVCiEFhtQdLl/sI
SWFGyrMum42sGpt6RIlij/4gBhJnX3VP0cOIwDIwfMiJWwToNlIsd1rnGzDaX82NPAAWPIb5jliU
jVVsmcmXjXTzHXO8QpR1ySgjC/TYtsqjzsw4yzeE3l5HwVINc3JygaZXXTL3fd2d2AJAuqhgbh+a
AxM0bAzQDGRV8Ebb7+/LXFlX7sb4sSexRZ0Uf80spzOa9NvSB+PUGh1ohqDep4xX8UFcp8GluZGN
+AfVCSx2OSTEQC+mFnejwHOnbTwDfsf/EqWEn7gRjN9uqAXxBuiYp3KFBGsbgx4n78e0WME1D3jV
Gj/RuM6L4mJjOpsVom1gi3gVjmWgfn6raYLvW/s/+c06WIUlfT+9jxOwwZ3+YA4iuM+EuZpNYh7x
LyBMrRaJ61sSTCRCM84HCrDtoFUAwl2PHN4q4Gmbc1pZAu0O7r1UBcLzdi0hZiz+mRvz307ErWI4
mzCqCA05bYiZdfO+wQp7mH4GuBaWoWknlFHjhYxhBe9R//qRwGx4JdOw0dIDB9opl5Jm5S55K6CT
XEIFlEmhkOh6CszgpH+E5BYHrc4/XgSYKUtutK3/u9BblA/INNP0yksF0OYXFgvqTmB+pG2opoJE
/NyqJRkicaUnwVz1D47FVYGFS+Z3foeOQVZBCEr2FWmOBqsX0MMpSmWSTdK1o62GalFihS+hba2t
YhjmJswuT5eReFAHVNOynQ6wsVCZtZb1Q9jGBCBLjlvW3dC1GG2LK3SXKJhOiPgthDyE169QDggs
l0XUTJnszqxqzfEm4jbUOXqRAOErQQ9Fm8m4P9ahwIPaFbYwBosToMWnw0+O+K6VpIymGAsl6oW7
3yu7u8aEQXx1KM1BDv+ApR59ch2LwRHjo2+V9VIIKYtO9hkdV2RthRxiSJ/bGACq2zU0beWYya8B
XH4aOuKp55lkas1pnxNbTNXoMMQJLIc8eaagXe/++fYoKt8RoUmLGx6ErsN/U+vUH6lpOMUwlOnV
pB8Ivevec9SMY6ao/BolT25T29og2IPMtI4Rrlq+6eHKFZrB8Ui6xIPqzOQwGPbx3beSghHqFZLb
kKOZzmy4tgN+1wSYOMSa9H1ugI4Th0sAUb9S2jkmb0N/Mt+nP9lJGT29YNXUnAzj9J5wPuuBw/nW
wysKl0seX6+D1IcdrAeh1MzHLwHsqHWxBpGYNN2obmB+WDotU3K944fp3UZMQ6gJmHvITJc19Ou3
S7+MQ5KYS2TrRDxkdz8JoqCAqfh8U9jD3c1DnmEimDqBMfpim35Ib7babNOQePEVlcuFO/xTQuvR
0I239RYm8uNu+rR2fFIH5DZVkwo+Zoi74H5lInH4nyILxf2hk+Ihca2xwEo4xjaYF1Wadh+YWsrA
qAXDPWtuL22z9DJXv0yHGb51cqDDyZpDZr7f/Em8puybuwkrKzCk7KokfolvubQUsEYvDtuKJsbN
YPUXFE+InO1NDDPJI+wfjfIK6uj2UcD9opZ+JtT9XzChInYUwfGNhv6Umt54xijZpjrmRJiUdDDY
Yih/RiWvxBNtf3afdXFHKg4Ezoq1ry1/48z/V/J/ah6Jey8x2W1Zz9mBkDIfDyeMwMj7+cvDjkJM
+4wliXpErgeEQPCyVkQH28o1YmAY0WPfgzFqUpTKQtlgN6rcNz+97V/GGCtfqd3+2jqd/3HXWqJU
Tgg2cu6QKJRtyiN1XDPhGkYbY7W7MPYkOypx8Qwp8dFC0fwxJ/YwBPMtGjYKIHsihn7l7RtM8XD3
ZujmcYre2fWmbJjkVdqtGOZ43nCiNLJ1lEtATN84RYlySrOdDNEE4n+N3fBM/y4DA4M/PFRF8F7C
pEEPJ7cdlHYsgQK4FhgcqWe7utRlnG3gH/YFWvKip/iqpj02Fiew1tKyOhV9+e+AtVFyz1EBdphc
CUN5SFqdwHNHG0zCXOJ8qaDGMR5BfBLc1INL28WQn4s9Aucuh1ZZS+WyZyQHd190zOaJIlE2XLbc
83IT/Zud4/s5/u/oleHroOPA2YhFwN+X4W0LGhFUNcKkvyN5smDW7sCdtmEQsSkRonom3lCGrRnY
fvPlBEAwh82ky28f1mC/PO4B4rQkbFYBbezbZwb8lqIUvIHYEris3nbCgF5WYuojyhE5VREFlse8
LiIe+VhfWoHUwnAQveObJ/QCbXsdACqTbIMr3Xq8bHxusAShSdeoQ3mueTWAn0KyEWy7Q7dU2u9G
o8r4g66BZaH2b+0hJ6j2+034raxwqnK7E2kuf/l3l4PlChu6Ni6qDfa6slf5idTkA8/pHuah3oyK
UkrPdwW871gDbXMWDn8sdAQ/h4zHortNL6p2RRAQTFMeeis+u+ay6BOEB8CAdvDIDYFLhQ9muY3j
BrtOXQeSsTn2swYebXNdc2ddCDvqY0w2VXtvulOrsvkG4LPMJKneQpO0XuJAzqftZgsQ2RaxhAup
bPDCvsG5LdA5Xga1ToW/gu0jHT6nRlpXs+sUzYgoLOyJ0+3LXnbKHwgpKwRvX3sbozu+anSxJkUC
Y1N9eLnv5q4xvQ5osPGdu37QFkzW4Ebs7icRBJ7gqeoutidP1shqzDji54PJCrm4eYc8pN2FvAlt
2AT0hWoY0dvGE99CWy/j9ijY6FYL330tlJ9boG5FG1Q8K0btFU8oIEbZbqhUN2uMQ7Q5lqMiqoic
O/uBSOwrQE8JCXOneTENMKM0v4ehDcytB/VZzPKMp0dNohuSJU6R0We6rynSLlI/0FThv4W1MucM
jxWsuh7NVCrEWBWFGUIlbUbqtwAyzZmvjrW/PZPEk0StITRledgA97Z/Tsxttm0W6YH2JajFwHbq
kpMjxiZYtG9HttMH9+bCYmxXUhAjbwfoo6vjkGbaftrtw/IrmI7ThYqXU4oUk6u5A6BEF+oK0CXs
wvUToljb8KdIkChdyRqRC6VQR6+ymmBzypNDk2UQl96R3Cy74d/7hueBLYApglnDT3ZDtIPKt/e5
etWW/a9AeNJq+IkW5PZBsmYP+kGFSd4XD57opOAhIfYhEgHRTUBedCzFH3049H4YVxXtEbdEqA4J
NmFCXZPrshU3X5w4mB7lDMaqTRdSP0k0YGX/ODpBTWkKzL6vuarJbAbYtSZYhDUqgH7NRd5YH6SF
le/371FBoD1PkHlvMF8VL7R/3geJNWrT0X+3j7WzV8bCTurcqgYlUk8jG/TQP0yiG8wI+wR1em9S
UX4GXcGvcQK0VGDjs5usDH43VnFr7QtgK+WvumwO0Ziz//D61nrYJW7LssdhJixSIswvNgd9ar4R
Gl9YmBXr6QjdUWFhBkazL/6yGDbwGdqkz0MZBTQgSItxYhPpu4/IjAvDVkxlVIbsYfJuS/aE6rwe
mbwK0Fj/GxVwAhw9MbKfNiOxQ3gmlcyXOBMpZoHURXrLbhyvgvoelCtwhUR9BUuQ2j9tKoW3O2UJ
+Dmsxb/0QYL95okZaVFzFYIu3ZqwLdDuP7eBcY7r5ohZrp80mgeOKn7pPgQFOSjo708EdzdgVS5I
9KET+nGF3febNYlEpG2PyLABbpx02gnubGlD+ELQzhrTW5Yu+J/rg0S2heoHf6ag4SY/4LhzRXiL
fUK6Myg/gqCKprdO47d8WbLCNOeJdMOTxviyVgJ7qttzAULv+ITVQxFvFLHnrCBKQXsxJjoQ/DOj
F0OUmo7SbVlqzP5Pzn9cDxN47L5y9rZqs9txFiApo2T9JmPgZFULRgHDK7IM/Q6NCKT2lMlxByuD
ru5TB4Z6WkWKDGKpRg8oyWE1jPQn9F5tL33szIOcG9MOx64Dxq28zXqJ+EKoPrEHzRQZ84+taM+G
fTDLJ9yjKJwf3CGFzYQsxV5jY2qm0H9dAAdq1T10qGN0gclPHlkeruK0bFO/iL8vV4Z6+q9aTrKG
q0tJdcWVyS1m3QRpDo7gdVufxJ2RNyKnA3KvneKxJI9Y1VEXybWOC6c+nnMmvoPnLzNRgKeziCDZ
IuUAp9DpHwPp4iU9NErFzBtyTnbIcqFuzm/g0yPYKyeBDpMC/TOyqIw04y3xiI1Ob5kaptDnBC6w
b0oQeGHayEmFeDIpxbwfb5I1qdBBDQCBPrWa7j1h1LJyeWNVWY9nIljd7Y0gO7ZsqamHdltnFUHG
TCHisZvAhQj2/UmA9fEFNA8UpgHyX0CarkYykkmkOdUq9zXxcS26hLykBJPzI2EH6GS2DNLrwK3v
llG2JSaFE8sWt2SYXrFojSOW2VKLsbwtYkO6v6REuKm9JKHXACNV1w7h/U1yqmR27A5zaRP/pr3d
rmXX8yOghhih+aVs7gHrYKeeiYQq11sQff1MyowFrZ8Xa5RnkBmoJP+2mlJMRaNSGphAekfM5C1X
abV4StZU3wiNgPGD19+V+q2wPfENiT/bTDdXJe0qpyPrYw8MYCStAErfZVhvcHmkBKt2dHwaXgqL
SeLrqQwvfcw1AvkhwYXDnSLEXr0keXy4ZYMJyhoIPt/b3pxqsS/OO6/NwJr2gKTHTDDQcl49RJY7
oQFsgEpHi1GhiY9YCN6by+yoAecz9GCpqtiIrOiU4paWFfa8rzYD+ckTWaW790h6Fldr7TbBaj25
QMidvFvu4bvsAcJ6XuuwiGedf+yhZ4ACc+LFwbHGW6TxpDuPBsZxWKQsvwlGDzZ6cCIvZIL4AAeH
a4wxugmcwFXdF4YpQ8X9gkQ0Vn5xMrT30u0Wf4/ySEdrsAwYSmTwVWYy/qXKNoP0l4b+ReQApLFh
Qzu25/S2LVWaCtLDADhm7+dShyg3dPK6SmF/TH2QhUQFbMmbupu/pqj/ClGudeGMcRvkCFe0y8+J
nx68tYFNIWzt4WsMNej0ToterOhUSDdU2wSGdxBqMVhTIsli9Lv44/MEYV+CdAbq9FngiXqe5XZl
QoTb/BwKpP2AK+bbnJx/i9kY/4MpvOwYUcaBT8Ya439es/UmcKZFo1KHcSTkvjJJzINTA851kl7C
07a5cJBRaO+XOuwQu6qNbmdxBdusLr6lHWwNi5+LopuHbQT9+B8oJxiFVvx5PZsz7KpODS/y/eFC
tKGRuQ2OLd9ltQGj9O/jIv1Xg1A6sgpl4AqgvW6qg8OLwvfqQ+BLH7/R7rDf0oqDsOug6thlf8fe
w6deKxlW1CFW0pYiqGhV3i6SCGSqdaD5eb9kNNUX9J08qyVBpMR49yIr0/BwVDF0X4vcTrlHeO4j
QwYq1X6X+y5JF2Z5ruSY8okHCKKckcQmWnFRF5g/KpTB9z/dxVbDDipEy0Qrst7JNOmDTtQRXxJE
eRKQuLG38fSqiEaJ56gI1AZ9QfaC4DDgG6hkjhHOCuuqtBFL20P1hg8s0Hozyj2ggCXZO1++90Eh
ckEPhWMkleqAHCcPM6JBWzy59mDJao6XS+xiJ7vu3tJuUDIptSDRbkca7nLif0jalFZZc9FuI5w5
cWPXlL7R/pHyajs3H5yvpY7gKC4jDx+dIQnFzMLA7vIdrr2QNElNdQqUQPru91jHngc3veA49RxB
2XYVpLlZMS75CJtVgB3nEVzPWuRPVpk8RmQS6U6tzBAhxDERCroPVMqPwd/aGcvLExwAK4h3WWes
iwGpZw6c12tj1Jwi3kQOLxezyYCE333ZJcXg/K8C7JladeXbRQXdoVRkBJLkj6yw1FhM+krkv7j4
Dr+Vd2gFfOc9GN1cgD31CitpVWZvyf8oRYlqWj9T8usrAtpEaf2sSZI6UZc6ZDi4LFlqPRQf2gx5
V+TNI9TKx5/p4KEOoLIac/9KYylukK8OV8eOMNb7O65ZUAjnYVsoU0AOyfb/zYzpJHbWLxSRT6ry
sgJ6sj2XsSyit1SJ5pZ+MIYYfvq6cQjS7wBR5USoQtyUQFiwFzGgcL/tch516yzsTMZDIZK39dZs
6+DFEv+8bpHWWQescN8xxAWMKnUY15/pQ0n8i/d1JhNlhPNH2dIH/8L7xhNHQVJDmJEk2++TPnRN
DmiRTbc15ClSwoI6EEfsrIMZ+31C2lXwKwV+sAvWLyUYUmzRWBt8LnWTI3u6ivcHIcrmsLu61czr
zwwX/htEH5t2SOXk4J7mwPhnYBLCk2FFJbzHOIRlbvr7fhKxdvww8RvSLXskAv9bSxlxeFw4QFpp
kcu6W2nGGY7xsaOrbCKXDyFD7bkbK7H36V/5IuCx8AunZC3aDKlWY20pMZh4n8F+CVadZMjjWbjx
dJR8XOOheyFzfaJr8iJKtxzD+hauVZVOMH1DBaNrPRvfzp/R4d6AxgSWVDPiIlcakC02Yb4hPJtO
nHU7L0ocNylbr5Oe2sE2WXdQtdFcG7brPbE3qB0nDsPGT06isB1z3c4F8WVtj89dm0/U4NuGqx6C
7UNZ8pF6nyQAXUBSIbPNalY5zyTpzB6IG3tkXS3OizVDYhfsdRpE43jsMTSt5IYfFkqVIQohOf/f
KlyXWRPO6S8D4VyniieZrD0J4sGcSwrrnqf6CPEe2M27nJh1jgUqXn0CtYYUaoR2QrW9d87JmxHy
Fg2kGuSVX4Apymjmz1HEI1dgi3pNj5MOPfkLWQ4QEhyLQHjaqb+HFn3U5ciSUsNBM7RKHvAxv/fL
iyKo/oEChdSjnpB02BxlPCppIeZHR99UJgI3icrQDp1yMNJjIIn15sMuxbAx5W83Fy9t/eld7gOR
q1euexx6LIVDJvZD2yHp/ZN1sXQCfsQZ0bgeTvtZefMxgw/xrboCDKfBvN2rVt9WIeifdAJu9A17
z57jJy8eO0D0Y6t+rQdpe7EXDeXr1f/yEk7IJ1Ehh45kDC/1CeGYWDavZpiye3pfiOHsQtR89G9/
VjfV2qunmf1iHfyPvGohkUbbl7NUzAyiYY6zZsytRRcOS0Is3Msi9AZvWB4E2zL4JEbgmFIYejJm
EB5e/9laioNVoPHw9cgBd8GDGarGJtQHHt2YnFRcoGOCGFdernfRWOl8aZ9CZFblC37pybzLgdHb
4Zo6jT56Utauy7um8l/tsr+0rdvOiSMPf1Rbtr1S1YY2fA+VZ4YkTo6Mjmw/GpEznYoNOWycYB3x
R8neb7k1lI3BMxwNrNJNMVYxoBngxr2Od5O+fxrisxH95OvKh8UXFWNlOdMp5pM7X4M/Jo6Jdoxx
wWFzjHQxOZ+at+AM5Zj1nY927zqRX2h9pKQyJzpLffEqcm9axwXzuLVKXMF9ts8xEzomq6yNmbjd
jOHj+d/WXC/m6Nt6oRfh8JLnZtiQaknFxR7qfgUhJ+MY3lBrFZrmKZhKnZ6RWe/JJEKBh1UgVAv7
UxBl5xQ+RGBzL4r8mPLZKLihd/rj91/QY7y42kgLxKA3nBeMdJRCyufMhSf/nxUWsgi0c4j5iGcU
1FqX56TRJ0ZDPUktJXQEj8LQhydPDnnhiIxbo2/80x8/WFFmsNEID269mHhoNiF+h032q5kMYVQ6
tNP/tW3fZjkASU+tJLk+A1NDh4LRfXwms+YiscTTKAitLh25nsPiYcaArY8BQd8BvE/DbpLhme9n
pgdlbAEw2ofX8dyOQGnyqfzhLzrAO+yyQJ80TYDtqLeGvkLX+GiJLxZkqauXqXF6QMZRLkH8oGG+
HY7KLv6WOHtZ2hmspj6m5hriJIEi93NMAjh4bT/Mvs6m5yNjZxLWY7ssFaTso8oLVGwy2X18skE3
uwgRx7GAVyWSUkXaHhH4AJI/w0+K5o5eEEByIyQLp/FsE0BT4nFZsrX/I3KFhF4vt+cNSFvwxzjP
lSiCZgO2br8cxi7Yip/G4UTEa1vM1/OHWbcc2g+ffeh6bxuUSn13DDoFyMgGBELdK04kcl5LKpt2
r35H707eUEB7NueCx1e0zRo09QqiALtl3g384z62SxbMvIUoCkfsp5+IyTQzaXo6R3AJ+NIY2EDY
WP/3Wlap+9VH16LbSMJ/0CpfiBTYKr/TnENJBs0ud1+EwU7ZMj3o1cxGqB067LiMm9qz4GR7rXF0
NA6eMlGT0bIgJuE27MRQkSX//9940dudOWmE6Q/p/pYqoRUAIgqbjJGi8EUmspzxhBqzrL44mgkL
I7y9w/6fUcjBfk7h6+kTVVj7wIgbn0OVGq+e5O5ie6lz3EDBdWpgGmNpOFhi0akqiTMJRtYwxmhn
qUVHWySmc1b7OYpvt3MI1RyCT+OcUuQ5uRES7xlt/Guxger6IJK5UlxXncyyVPqzwi60Ef8mSNsB
AULur82ra0ozaKHM8wznp7R9DlL5CEWlLMgYouVawBYII02pKZe/tyHyiLO5p+zIshIaL/wyF5rH
zb8+YQIQ7CFqjn83XAKBul6NhdJQmynpHbV+AANFjRSxdM8pwiNFyuKb5jZNNNIxmaBxbl7q2/cL
EiXJYT9/OcU8vDWtUvCsPEjHl4zGpSlQo8UCRDXVcsgRzZ1urtwDcJGI4/Qebg8vRqpIVUMFWiR2
IXDcUVgnXLjkGp48vJ5ERTx2RiYy5xCP+uY/rJPr9zltIPN/TWMOri45Vsq8luMyX4pweFoBlDIb
W+CJx8iSZacAL0mEWvPeDJZrKMb6Ko8DUdFnnDgj927KnqqAWLhUmuVPL2qfCqZoX9tvi3XW8lCE
vXEpHNrImileGjBCtJcFylLUBVlMlBKpuDhJkVzpA/F65EXFNdnHiVSvRen79ci97hb8pU9STbna
fGZ9QO1jsjLboFzhwQBMxWbh845J7vPUk/kgOoZEQ0hyH/7WDmPTM3YHlSr01ObdxJ/e0EAd0Gvl
gN+Og+nSOX8hI6ZeGBg4IenSgF8ycBCURv4QFdHKMokyTXsXa2wQYPgmysHxdCexv0ag5lcHapHs
ZwTWS2TyYeCq3e29gcA1P1Ks6au1xWdLUSNy1uIAVAyBEmdi8Slkai21UiDhoALlRH7lovDUoNI7
uZN3OCvWKWhUe3jZrmRakcLAek+MTmrlWcy3bYkXvUTh0m+5SJqTsyKYOca1jxuQSxylrSyjQg+S
JpDh0va/QeyTHugu//tA4YfbrmAC7qPpQzgXLgHvzOfuEUh8NbTgmxlsTdViC/KfSzAOhbNI3xgr
xOmKSctTFppMq6UrVHDVkIRmDeeMXe1/rZj75a/hrxsmJUSp2tq2Pxu5PhRr43KjbdgHa5pgEffY
4kZJVmJFoods+IGA1+0WPpYwaEmtSRbTbTn07thH9OPgQ0OIbIGcevUC0Mw74u8DRDtHakhJQ99I
uCKH4cGP3d1si/svEwZWKS334PJFSpUKBylEtlER4lOIVj+makBcZksyAHoF+Zct8uJqDMSaU3vU
6o7HysO24cdaFcuWGT6Dtkc577IkANGJVkIPVjyfl8NvyrLk/3276ndY42d6Noi7hgj6g9IBXXoz
8+nGXyMg3hf15XxzYVxImXn/znxGmPUkV6//6uFWXRVTqCLswcyfZbK6myYx6askq0HSuvqbSbYt
8tB9w0TI40/jNUQp0+ED4OvIpkP9MsT2M+uABhKo7msAjNH1DEY2Snx/3BGVtisPdsrZbblpz5Vd
+jCEQWWKmvxQmTzYDWtw4L5miBc7dOvE2VtymzxbIbvbU9Y9FGwfR2hcSbhJBRuW4tPLkck3yjtL
U8vwYvT5HnIs/TNVhGffj9cFbqkth97lpg6WNDSbqH4ySnYivhBe6ajCyHnspn0zE5N6au2GHg6P
jUPG1eYMhHbevbDoOrC55kh5tmFE3DOzH4QHza03LG8EVJuYXhiDlmkzzjFerh/xjkLAQbFpXrcZ
ejKjuzBj0IGN8xcuOL4xlTTa1LxGIqqcawvhEcsgM29maI5lyhlvEsi4VCp9aUADgMQJpeeqrTjv
lolFjq46UC6JRqZT7I5eARLtsQvRcG7PaV3tTfFsg2XQ19r4djy0ksBb9eKu25dmKfF49YqcX7rO
2Pa0D0ZMZIzEd29iJ8jyl0trEh0CBI5mXgm19ZHOGd1DqOVnTTAJLGPdGbXnw9AkuqP3aP+TEYJd
CTYZLkplNN+BkViSTJMc3UZxWf5XDaQkhuM9AP/0JVUaQgNme+luA/egJNm2vcO5fDUaISD4MS2r
21/mpR9CqSA7yI8F1LOTx1tByPgfBZhbulrahC05MgXLn97Uov7yQPCMSzfvrhQ/f4U4D0cZLCcs
270EcdLhzsGGlchF1QzPJu4S1JcNAdnMLUUYr+zMC6OXBXirWBXhvD7ZQT+2WlzfJyVTuiOpr3mz
7GTcRsV5P+TMxKAceLFONES8OvSXUsD2do+ks5ykV9lKxqdulwGr7k6KtcNO2UX94iEaEdOFcMVX
+sbff/lW6M1uOWR6WLjNavmSNgI5mW9W0ZKUyz4iaDxYzeiPCin3D/wsaUczicFe/yqSQSAo0YWv
dUYG+h6kuJp2hhEwuRemzlE4pGUKRY+b1OE9GY9/EegDvXtsZTAtkDFVbMIFK7+xzD2zyqH5zoqa
qQS9CNyG1aM5+dMC9N7KuQYWc4LlU+RC/yaqHipjgsQ6MgsUTX3/II9xw/AS6vT57RVmRqCZcQYq
5z+bntoGDD+eHWU08nOhUyM5O6zTaxB7pBxdBVKJqhj3/snICcb2GS4e4FZ8kYeDXTPu+cYPyTGi
yKOuANn1R6VmEoJIXZv7Ag++bCp8nYZ7enUGOyXknnsDBqc0X5dIp0VFeSmGjowMOa1Zz+zZ8gvo
h4MChLICweydvVmczXzmir/nwLNlW9HweTqhjkPTtVWgKcSXJcLmD6y3igCpFTbPg2fQlr7Q0ZS6
faJTZ4z1xgQJNgO/RkCxUzxkWIjYWqYAZY0VQq6TeTksbRjynyPuHMDlSWnwtMU24M+/RcOuLq1e
M1701IjGgFw0wCI1RrEMDzBd90hWOh/sW6RQBhgEUICMQsRVZy/bJYXEvptezaFAb1KPlc2oxs0Q
sBtuH2ZzmLp560gMgHRVv6tCQHtj50wP1riNMJbwbtHFH0vbpCl6cUDyF5gJh5C1IGNb1GakBTKc
DAkUQ9/5uzperVbwJ0X1IpFCOLFh/xKiwhb3lcEtWCF9PSQForzC8fhn7oqYCssgyu927fVOIESR
QbVUm0P2vofpVyuogBUhGQb5R4KVBsALpJB7ZXQ7vbSYcAHoyns3XALUbluqKwyuexpDxwifqLHQ
Z0wKEGA2qbeU0+0GysBlQneCLOm9ia9ZigXirnB4/YGrZceiw2BSSXbsb9mAPIO9ETKvm2s7niyE
UDiv9Y0XAX2PI8wguPajoN36k7ZKtv4ltpdA08Dp4jOIYFax4LC4NHGXg98ejFjUeZoryDrS0jRn
tMbZqeJghoyq2YQLpSA88+c3peHI56qKnm33TjCoduvcscQMS11QOWAWg9cJAQnBG5WKlYaJlcRC
JsbbK9KBOvOM2s7gNRuXkCdsZKAAOSowgOGpTg3R8UTOh8H4226lKLJTunv3MX80Z4ckA5kjtV6c
4SYfjBpwOyLLo5VYAvGxuXejBB2lG0vkHLqzLwGc4G7IXSjmVfvE5DNSyd9yoTh5izeU3ykVsoIu
NY4wYDgq+5D0bOD8aw3YVPdqmmNWqm4Z2ItwNuAfesSZBMpHeG6wvsV279soGU2oY4y3zKmsDnos
gAtq6MdrhMKWBSSwLSycE2FBKfMqFhF1lqRFq1v47nXEJqB17f1mKkhVyrwhPEM8bW1npo18GOAU
oT5QSSzHjl3DO81NhBvP1P1S0zfnCBbJd1mSmJDQ1kxpCP5wNj/S6h7vujD9vRXIvFiqwNwIiq7W
p/G1SSJC/OITFRUxRETZISpZHrYTRbw/LDdOZR8JcoEoEeL2z41YyOmLiPZwxsvt4Ugmt/f9cEZd
1JbWYX0k/0I+tyHvXtBqvWYq5XqTh1mKjXEaHqgmXRg0E7z2TsNXnoNH6VyWcPHV5+wH2xSq4Dkl
WTQrRJntdZp0cZQKlv2dQrwCqTdXOj/UiCV11gpDNKuiwUnkdftuo5snyEuFi5W0CnMQsAb9sqGi
cNPuZDbKfA6xfOoes3kgF3waAxj7CT1eaiF9WQuvXlBOEvUahOdPSIr5TiR05RixRMClVIMFgCmq
Gu8YFed18vgz4s1hSirXyoTtBb+t06cGsyFtm4uWeCCXYV0H9bJrhWZusw8gtU0TTB3+FcAWCJP+
i9k9Fey4SJfMPe1w097704Ha5sxDjItXMmFKFd+sHC1AsW+/tYSF/Pv3y43jeS0sBgD68+QxkOsR
f/6mXjRc0bUn9yBNfSccWvZpCMCLl1S+f8Xr2W+sA0E64h9LzlredxgOESBAbg8/HgQxFUlazxFZ
sB/CNEQAya8F+udXA1Oi87mWhKFf5YMmY2LE4HsQBwQxSBaGfomToKnblCYalCIcl5NzWVtk/DVe
yPKiTZClmXhhFKu2O8FdpcBDmHY3nAV5WNavnfGgOlGQMP7r7SJrFrxO50b3QdJGQMJinIGR5u5U
GTJicJDek7nfkmOaGs3lVCDsYex8EsXn0BrxlBMLGR8j2t3eXDBsEMnFJRwcL095dHa4V0U+ADFA
2CZ7J1Lbd9Dki9IYR3cGkK/QWmnoPc4JgsktGUZqL2Jpq4iAT7cf4aPYVKDnk4pt79fTajPP+yrr
ci/ixc4pOtFJXnnQH42FJm9XV2/4t1FPVsHYc2/qN3MSRsUt3lJVyMqL7mJGu0n06SitoCdDnDIp
GKamGyCLBNrxyVILsqNOKofqJv+f4WTSqiDdQ3ZJitDKsk0K3A6m3GJCek1ElEQllGOBfqUYCnHw
qfRZERW+3Jy0bfknR/7ZrHPy45cBWZgnIhI88BjfwJxoOZ8/UilQGsdv3JOVB3mQdp3R4v3ZfXWv
KixzwB6WENiUfVacqTqv20CjXUIB8khBKPSIiaVoncbJZVKKworZX5518TwH5Xe3Gz2lgYYYVXau
L8S2D1iQVLDpGfUiY+R+8L6aB9RrAoWEVsK1JW/IEB6uhexx4r2mOfJc35uRj7P1No7qMBsVvy8/
Zm/oXTaRNnWeETl1neSSZDGnKvOidfv+zz94YcdN8n93S7DcbMDRpaJQFszUlLdBTTvgo/U+Br5m
zRnx0jchKnM/0Ln8w57OqgVt9Jp3eCUqxsTwi8UEe5uTQjMJDHXXUz5I6XgvaT31+L5GOHJeGfiF
eHYCDF7By+3fenaanj0dRQpVt8j5TIkUkLobqLPDKJ1OJVPD2n8PIWaV0GkkjU1DAjUQULNoiRaY
UXsAR6BZS7qMEKZxLveQcYM4hrYM/V/RLoE1oznz+ydH3Oou4bkqOqvHJLnwn1wOJKbIwEg2d3Vt
uPp5cYVbQtiA/t4GsYhs1GHsYwEoGaT4x6wfBZO52kDJPr+I5/PL4xLx5BjA2X6zSTTMLSqMitfJ
CyEMAusLy+rn8u8C2uLAvux8IPDUzrhsESZwpdymc0mZc9PMAgb8vqiuiO8z/8iSNzLy8vkX9N7a
6Wf/fg5ZeAd18kY5+hX6375syMH6897EQquCBKEIoNqU4Enmq+glBX+YtO8X8/2xnaz36r+9bIaC
7cAbhV4CkxRGZ53vwdaJS2zOKNTUrlig8aQmewuBiHEPCVY8GiJ0brjaGXqHyjODnU9FjDOHOrvF
8oZFpsDBK8G7Ma0OluOxidtBXAQloyb8DbZNJRuvUGNAlyer5AUj0wYIo4SAMp3YGfSCbDwP0m1S
VrbzPau5q0ImWtAT8MFv37K5a9s2EsqgwYDSL66ltziZGrAluNxXiMSOjynGdCfsuGptAeM6blwE
5BKGuii53cBXsfJg0l8+BeWgSfZRzPg6pip+lXmALMsMlkopiE76tgIIL7s1pZFGeKZAL6QiYlIA
V5f9FMC0/8CKWtzBtgLBqgdmKghQ1Pm4hSuD2IMEtsV2ARNqR/Khdj+Sce9xNybf4StnxfhYwxR3
B9ZLWBENovjF608iJ7CdIcRrUHfHEiRPQqENNcik4f+KZNbfGlQ4SyZug5dxGjpamLGkthAGjP3S
KvYFh2T7WQt31LXX8TzgU5F/Qe7IoIxAK1VbOCq4TOwiFloup9gUhZlAupnZWVle9HvJ9zAU25zN
Qe+iFflV9zT9i0HAKG78lImfKx9L0i9s1u6iGIMEPRpjfTd1TIQl2sDunmbB57beO3oT07wl+Fvs
l+4R77tWbEiVSrORKpoJguMJ9s3aiitI4CQPjXy9zjOd7txb108cMqHaIUXYXM8zj5DeGxmu0MYF
EvVwvqF2bRPiLML4r1t+wmVvIOMeX8+nFqkI1EY/dOqUrbVKdp/jbhsUWzgpfhYkLJQVadN1O5/R
7EY5X1/7dNJJ88LNGYDFtk1RStmFwdICqR7p/YzEta2CCmYSFAMbY/Zm8zMWU7DdR0vHaszH86Ux
gM8VXsaKqpSl+VXTsnCiMvnof92uGEbuq782q+X7DHjSnMjOk12a/pO5RnewXgbD7QY1O4jiGWUR
tidZGCGjS1rLxzIjfQdu1wkoV5EezX7vTlFNQ3PYtb7ZEdEweymOK91K6+87XRLKjEPjFY5+C35o
xjaBWirnJxRPWFJRrfZiy8QdYD4aqdELYDBgv8pDDBhvSt4HyTI/mGk/E4DPMi56BBtNEIXFdGVk
44y8kyIoNRnMakkFiFnDX9h4/jTvJUdP9ORshG62ot6n90jWSA8A0Fb7oAOUCSfJxKSrd7p8MebP
+ks30VRS3zuBE4m4qAJASRtEs3aROIWlwNXYZufBTgzPbQIyX/Qvs8/UvgL4uCR6znBgpGFZmZL6
H6ewOYe/HRd+BGJpqYwkooX2dSrRJvXhhDZt35hLI4hpJCxdFS8i9G90JHY6r15bucJRphOoWvSK
/l9v+8xjN7admgnyBB7qEc3zfKtqN/ZU8s0vVbxJRpySXhcH4W0BDkE4+cemKHzqnmiIr0QqMMIb
FOkCooIe2Pj3UlH1ma8qKBdLbAP89oeyoJQ+fsEmYv1dCdAPt6sptAICeUBqs4iTSUVn8nkIWI0a
/MRDt38EedDCkk7U9Ztcu6sQt3euiypW18nanSd5fCxmGKod9WVbLpwEBOkzhFPoFuyes4bQ6DW8
SF56AiuZI5E7OCBochA+QPIT6e5i9cX5MZ+xfFeOwCf5B5pz09kWe56XUjdxiseKDNiZTN9xR88f
YhtognA8RvWcdUorutAF5Id4Ox4isd0cmZ1iw2nWh1NOoH56sEci1bMZoIF/zQE5z/bp4AZTcySi
R1kVLyrQ5vIi2CCdfrCbhQ3JHwNkz8KdB+OtE28RtZ222rY2eBb41qa3NaAw3hd8SU1fInSqEJUH
/+JCB+gn+dep4hLKE6VzdT6xRFsD5fO2rNED1zTimr0dfD7y7Il6zacyjrfzKS03DM7GC5Pponys
01DqIVvhehI8uYFyvw1DO1ANlz/NhV/bTPMO+gbDUcAs1u42NOw0vm9zT+NXS7/USDkMa5i3Dz5g
2MPfflm+AvvF+WgnptD440rD5M6NS5Wo0m5iL9wFwx/jps2JjAKPP+mFUeSsZq2nA1ow8QckVLLb
0FVAV51sC/F0pjO1Jy8vZxG62ZzWGwjS3m9i2w5BKs/tp/3tX+Fdcb96/DU8L21UHuu5x6DegYJa
b4NhGlhFuWJ/yi244HpN5kEzztkxz0qSaF1trMYxJ9S5pKvZmGAL/omFdrhhbUGj944vCKbH3HUq
oHGUqzgsAc4g3DOIGsQeLzyLHUd48643xRiG0NfeRLROwb9/zCDPJsu4btrSn2tWzAFb34T9skvC
cfZOGZRLQGYzbW74hCu/UJayQq+fm6x1aBYkWYCLb1PmBOCCNaZxz3a8XQzZkrZ6i7//sEQW+wkt
6sOlNBNr2D/vFb2X86OtqTWZoHEm96mc8V4JZmOXGoxcQPe+jEhLMCq2DSLO/Y2nnSyWjPXmLAnY
ubS6h/0fulqYpHNElGyt2LQB4EsUOsGiewaYzSsCLL3AZbDQ5K+eUxAvOY3BjT5Udy7/7daUNTBm
t+5jLFSKIR+Ar3bti886h/P/TbW1f72jiFKx3khZepBqSdhVFEkpr+z3WdWbs6NEU4T9snPxHMwG
E8qYzBUZsobx2AWkUcqCZzZ4wZrI0wMPo/D+dumTEH3TqgorUqRhI78ocUjSJuzU3FQY96f4npKT
C7+ypB61geUWM4k0UlRYkLeuGFuZ2C/wsm3+6pKZPCITIBQjvPj4kgeZlcsJuDBzfImrfEdlzs8y
tFLhq7CHw/hARlbPdT7E8JxSnMT9yn5AKLXHaWsKzhFWjP5H5vIB5HCORfqfBPwzTMHixvM9XUA3
N7k6X0rApgC+uXEri+Q2hy10rmAxSgpcSGTU+9M7fzKwvPfBsc3R9PtzSTQT21f1/HF0GgU7TUE8
m5kGYIN0o9cujv/4+7+8i3XJ9vgHG72jQURvcch7PAlSb7D1uGr6HekALTS8gPLEHLip34FK7TXd
c/pk/EXVJs7RpaNIzPkHpVUXNTVoruuY7aDCgqRsEoyoisKQjm0+mc8qpH/h3qOUPJCqoMUuZFc4
9Toozk2CwwDRJmOKc7BLVJo1Ia1ZCxLLIq1kYSjr++cRvyrqxSkU5W6p1IrMFVEVk/7eKGoS8MY/
9XT3esot73t5DzW8N6hcuM5LX4jmcQHH5W4e3eXUOEnSOBcim0AuqhnCxltKOoES6pUZg9kT2Pc1
L190AUwdCeTDknhzRMQkBUOV3iHqgnBpKRwxvRvreTigEnLXJd4aLw+TBgAfT4AIP59jvc1i8+s9
a2atvxmEOIL7dyQgKG+2szojo93VlKW1iShs9X/IHGMLoz6L0fV0/QivhHSJI5gceEV6gMHJaN0T
okuqlqJx9Kk7kpVJ/mCDByL/7jpaw+dF3DxtaSsjtNyeOtPEf1nZSeQA83Cq/HA/1VzSjBe4Pplk
dRaQzCbfUvXywrwv7cNI4qfW9zywPENByzv6cEskERWEG9nGyGPjzDr8SRxpvb4+SnwGeHRRGr/J
Zxj2Drh89Kl49HXhjDfWOTpbvzqr1KUlIDnuosy3ETS4gPi0jrhOZ5yWICO6EVrVRzl2kEfohDAQ
sS/H1KRzJvAr1L+2mOWUC5ga/cWqDzwWCFOBz+n/EexGUkbTPxq7EErQ1DID0uDftZ00Mz3fA9h6
cv33Zpa/eIy/ZdsqZOWKVIznV5uJHUnurP7nioI6nZsdmS+oE+h84+/v0sTTQEZXCOUqaD2gOX8l
sWDnfszwVgQtl6wL2PsOOZwYqGlMA0Q3Z2xQ5+CwtKxSnIVIW2SZEsSiob4cIyx+aslDsr8ePRqH
LQDSlrLcU54ms4VNgVovtCru4hkHM9+3sEplmczJ67uNAWHl9Dh/aVuCeC4QmJSQYAI+NpRc43wQ
rZlIPiripZfcL68JoSTiBeiY+UezGE1LZ3b4gUeuwrGm3HEQnxl4xE5ycFbF9cV/ESiIQt3gL3XO
L41cKqVIfKnusshuDyDUUI/lS8GaNLk8fz5ZmOXnZZuzyKJtCuCKoz7kegLz6ceYig0I0gksuEk0
gA1F2c1tELrkK1LMuE0nhV+AQ5yfG8py+TDzrUUgDKHYFRuqQBdcVW3beTd0YIgpJ8Ky9aJoHreU
iKm0K3/Gqrd5pv+2wXz7nLZG5UN33Al+tv1+nMTBjaVYXilu3JPxGqIbg4f5Y9898ErWui3gq3QW
0azggEee0qEDrgFPcf/rRJ8y4ZDip2Z3/qZ6r4Nt5QjR+6N4rBqlF9DHKC9fk9E1s04b+0tMFjUR
P/vl5RDKV1dxl99/7v+gR62v9VjKcztuApYUzpqhIzfy41IN8YqFP6Gs+XVq4T8XXlGgHZSMRJOC
lKV4wh5CETjZBIQWW9IHlw9I1x2k/iW9RhxMEqNPRyFkJAu7oo+9fGOCJosFwnD7gDbIvGl3ewtZ
J7h1S3XYOb5j9pqdqKxaKvoCUTaaNyjumMvpmU9XXVm7uqz3U7aja1N4/zp019v9UkhPYVcv/gN1
9mvpxFMAFx9GEjpEo6HSnHPZTA23UfXZpRxU2LF067IKoDN95kj9ZHwl3d3ivZ1rWxiFoJeZnDg9
x97eh2oZFQIwEfl7y0e6wIxfR4hXw653TULpCuVOLXSbvC3c7JEFqiiaxruTdeqr2CjXpuL29fd6
SdznWT1bB8+LG2ZG8v/otqrZgYYH3KWXQ9oCHmgpkK2uEWBlBZlqTk2nzA6StbZxr+W6x6j4aFTM
ZX0KOq7szXLmUmEX4EX9/jPITRj+dojBsWdyPINnIISrKPIqp6utGeZTNLQ2r/GkB908aioeV4kA
koSg3sIRqB/4+0KRrlrloIIavL7gfZrIHbFU0V1F5qF78S27uPpPlDWUoyiidWKo4PDZUv/eFbWr
XiThzwA4MLqJBZtPa5Pbyx/BlA9TOOPKM7yNWNmDrNmm42mq1vJCPaBYmh3kOv341UdkYwowSRFn
46lcAz8v/g682kwBqCUFfgef3CENXl5NgEmXXqz/4eQfLrODIHeTZtOel4TFer3UuNQJgU9yNFHO
/rSm0oEiYL4ZufpiCI1Js909KDg5cOdP0+yLkv2wrMjBlL1LaRNQrIGUVI4oano6eDL8AZZfaQoE
4UMK1rHTfypmk5jJ3NoLH7y5hPMgD1OyZ4RzWFlgdGby93H32ZuOvgFbiZ+ZqvcH1CAg5FLQ2iJB
TTa1lcejyJ0pHgTkwNkPKqI5VGguUYCy7VC1QrEVY6SKRv4n+lKrnlXcRgAu7jwGNpQeITBIMM4T
YGIYKN01Z+d9AefA0XabLXzTRka6B5+DlxCbsVGn8XYKDLL5xrhwughITUYeyfD3cI5HRVuQIamt
0clHjIBguEffDixMN2yksfUXbaSjxgq+waBkuNAMEv/T1aEdlcI749L7Wtd1Uqfc/73lGy5v6AOU
V1OhPxNu7vSA2+sObPdcvffc7FXo0z5x+7aj4+9mXnWEr07dGIw1h5DId5k9yNcB3EOMwbUZO3uW
D/ktGMeSeu5dws2tPVuGISym50MRA5XWYe6d3YlG/2JZ2AiuWuLxRgcSiWBFl5E+bC4dcpplNxKA
ETvDceghFlBTWWTIicypU0hePaVbtyQfL0FYGBNYGP+atihApmx75TiJzpDdypV/cgobWdVLajkB
W8CVstPnYxy8PyPdedVJjx67Z8zAlF5wzIkNAmulxt6aCrLdVWfLovZYq+cgCxtr36tKPnsGj705
+ExBWMKzdrZzpTVvS5DYWvbtxdiJO2M3+jt/CU5Mg4bKEAQpVvQqgNNNyApwbm1h9y3Tm5GQgx2u
qNLeyn2dUaTS3he5JZh7wFD6QAjtnSDl95ZIgccuIE//iROFvt1VbiyC6NnuHg+XUUJAQ/wqtdT/
zAPo+X0jhTx2BNxV70Jfhmbj144XlicRdX3EC0Le0Lh7/LO9YunUfWjPANy0FuOWRf7Q0vzSvvco
loDmf/3tclqNUwjXr+g422z8hoNXAf8khQzI7Rs2/CV0UghmFnhuS7cFkrIFkLUyTS8i+X7plH1q
Kg0i0gurxjKLTxHsnI6wiawlpak6e5SxjtaBzg5vDGAnUcsdVTXJqSQRWyKt2P4Wdaf+8nNtRLDF
iOKq2O/xxjP9VVhmz4x0Q+PMHIFG9v1Jw8P+elDsMsqONBJz5wLkOwLML2x5xMnvio6To0SGwMWu
+CsNAmW4caVvPIAlDrySRuf9uJ2NoA0LiibTicernlBZUVyEtDec0d7uUr1TQuopBhGu0mFUHFEZ
9nsdg7gU7jSnID4URDpE9BHFtDUK4KwqyXc/4YY0VXIQnE/uSPhr769fHjro+w8rWW86eI5vF7E4
J0p5HoGisQXDTrbq6b2eh46JxEit4avjzh5MGkq7qOTWFSKIJjDysgMPMyKakhCLAqJfVJNhqGo0
cmHg2kuHjsKH0Aa3TrENWoR7a+/1+EtccquVUtWFkucletHgBuJVGCEbRZW2VEbk6N4XJUuK6nfK
FJDmm5xSiTEAl92lzAu3cF/003lMMojET1ifPHgR+WGFN+ouh7+18UcJHDbN5zl1CEZynzO3kOYS
+WWqdXIUINdjdQTbtCuM1VET2oU3sYqj/sait9LA3ZIYPzX3BN2PSDMKWlwUkGD5TC2WNihDstih
BK2sNJf3axeEm6BcjsFXznE3LRTBKhq1hrAGJ4ewAoMc6DXg0qI31xPO+QMnkjidSjVouU8TEPp9
OoBg31hIWfJiIQGbfvJ4noDfD5QyrI7rlGm4mcFCYCbDdV4VSEbkg7oVS1Qkiacv3tcaiH3R1HcR
fnQU21Iz0L+IliDn5wZHSOMnLqyyfVPF05rSdByqFaZrrkCnLdHtiu0Ox4Nw1RiSqRk6/eR+Xy98
8ONsPlXDgixPngGXYjrYkoYtcrlIkplNQfMiIIliJCo3xsmJKJTvKyTnte5EznU9ZxXNACETmuio
6g/IrB/RMflYxWMxMCvCyLsoIu/1lMDdjNZJlLxfHHA+Vwz/OnqynJAXApmWkhjwqGqLDcLo4ZnP
D2dHTj+O1+QL91q0XmWwMiSjidaNzhqePsxXUp9EkdyjX2HkhvMeJ5BO9Vrq4mwYiaFDFsGV9mtU
+BXbD973S7PRiogOWSk/oR2zCou7VP2c/k4zXUJyhKDnIfCPx8l2GGrxRt0OSHHmrRksAbpaOBUJ
I0kBNOo3kHfQojw1cTDDIsup/XDxgC3DeGRSTdZMAm+DemNPQkFA5exVHLa0Hi9jpbqEnTqN+YbY
hn0XWCs79K5GsEOgwDa/ntI9YLduSyzGIYQDwdg9PVGVxQNgx+jJHG3jRU9bXuEE1vxR18VfOk1o
fdqgXHvKx6DF64fHp09+F6pCKYLKj09PY5yzsQyMMNlpYAUoAnml++qHVMc2zzZcIsyHv3cBiZNM
jAs0a1Izo4eW/sbfjQGa+gnowspu79IP6+pOjdHlzHHyDgNABgEtOjW9z1+3EJyRynAh1DlDlavl
NeOOwzQe1b1eydrx4qXfuUQSyUr0KpjK6lz5uXINQk0wkQEWH+8WPUhHSN7uRz00YBfNq0Ls3sp1
zTtr0EHlW/IKtauUHLsu+pmIfH/7wUaMTZPNT4mHey9ReTtyVyjPbZIHVfjoXmAL8CdX354IwvqV
Do+zfqeIEx3VnMz8kuMTE683zqREFwIDipZOHDoomefxgTJ9qL3rA9Sb6WwsEcIPz+hMYIvh1lzb
eBtBZSCA0kXgUwO3o0iDpUPFscec4IBaQK2Zhi5Q5/z1YTPDlE7uUOdwDE3p8lStoB4t/whING6F
x6aY5FxqJcXvXOk09A3VmkudWL+8+Eky5oU4PyZOt6WCRZEo8PkHCuSrUHKlm3FZsaeY4Up2A7bL
NnNxnKHrZWwhP7L1Y6FdTexWCpL3K9+enFDgdWLvefhzFsTe9nv/ZFkGdKQgK8EV85I2hCTIpTZn
sreZ6+r58V9tvQ2Z4PhUIv/4bqE9wLWREBN2Jlrt2+wMgopUNUSGbWKOsuGoc+ST1+9gealN5nec
kILsAYxWc9GsvhkUMb4YD8niXBcIpdgyXlZ89pJuOsjxciCd+mHsNmmGNkw1n8DoT5nQS/dHbr0w
zeqkHQfAQveXkuspoeBBq8KYSbcygnF9FuEeG1YNctu6jvNweNRj5zar6LnyF617xGGsVCAb5wUc
XkZWX1EKxISHcmRPbYdcb5fm21NroKfvmTDrp6+APN3ryKatM3tegM+eiA1FGlOASrUy7Pd89ZAj
T6WQDla5Rqaf6AWcGLlFzTVJxAEaFaURtTuUf5Ov9o4pS8ZKjjcBODP5hAQQN7A7C6FvfVMBjCh1
tda38UGBwykSTI4Ja25zIUpgc9IGldNe8nr6zvKFIw+Tw+TRTIDrLnJHMO3Q4teyVAbb+2UXKIur
0zuMyg5sW1an9MRE7Pr/bzG+yPd7kXmR9dui5n28v4N+JAjEZHvUriNhOGRbwym80v6XXb06f7R5
bpUTMaQRaknt0sdZPi4M1Xba6/jrCoras0Eiq7Eaxg2NzKDtKoISHEkbAu5PJb10qsViCg4j4gHv
al4xAh2N5Zw1jk5hLYT8HTctOrhTJqF6kF52rMGn9kWqPw1ElDDN2TOTTMNFz6Lpv+xTKriEritA
5giwVRg3QoQVM460RtAq/xJSAxRF0ehA6iO1IKnq/jruFwTuMoBsRQLnrr7qrfoPD7tzy0eyJi6z
NAx+4I80XzUyjpHi382199pS4drurTFwj0/6PRCiV+lQBLss1VEpZaNW3zCYrNS0zkIRPagzPLJx
qk1E/qNyPdz2qfoopY7hndwloYODoh4FoA9aNzaIrGo9bjICjrbodMuS6Avy/fuGUJ1TmHCzXIS5
CBaJY3QmrjJrBDSMbOXZ5GaVPJXKFvlRlLg/4glhh22JZKrt7QMkkIugHtCk/a5aI/OgZ0T4wcTh
s9EPnnCidKowlXEvw5RHqlZU9b50Effmucq/UavrikAAo9CxTWAOTrFXBHxU7h6EdCEpVoxA4kW4
ubU4irn16fjQQnw5kEAzBxOju1amD2rbXuLFJ+09XWbefdvBi+0fAblytdR3eu2tXaLYXMiasaw1
vP1mL6rsT3jEr4qDi+bIEJf0jJiujb1UVQMh3kQcuIwDK3n/DaWgyq0RijrMj2LeLfLbGe4xsNHZ
7/F4SJM3DRzYJVwbG0mjchrboMR5F/+z6JwEgWL3OMLgPowqzKVcV+tHOaHeqKGhB+08XiPeFkP5
eBKJcaZfCyPW0KcEVKKEMZn5c7vNKhQ59kzsU7qBfIxdqt0Axd/GtmuA+VDOniaTUoqW3rFw6nrR
KmRsNj5UBiRZyMNwj6PXN81LR/5ij3cE39YRAnglBo2sNz2Z40Ld11k1gxepak75AjHSwUKjW82c
8ftiGYIOJhSnUcIcnmCMy1u0blgPyRuf/1TbOMZmaoksYA3zZe4P0I8EbK4JJUxXt65pO7T+OizV
4cxE1q6hLYUtox0PNrYLyEwVAcGGGbsNdKQ+7kHxIE+Qlilq/AehoB0ZtBVXdFGsjSjkk9GfLpN0
OmtEB5phPE6np4L7IPJ+RKnaqbLSG4FM/XBXxD3QzwcqyaB2VO4y6JnTwfLGvfVGYph1F1U1FegL
2LHVIL34ilq4ltgwTyQOJn6feOndzc+9l7O+oslSTLxSp+abgITXtwTYCFRNKd7Qz80IoiNpq8pz
gmsugor4OI/Iw//rgYgOXMRmKxjzgpr3kzUUp23YAEZeCFxHa6OWQaaluBE5FDDeYve+xRId/xsC
ELmG6BmJgco8oNH4kuiCGoNDrahCVrHfEBQQ/1HIJ36JHDCuRU6SCxOTLJCkzrQqsYP+ldGl9Ong
N0iFibqh8bHXkiXAPNAGnDKW7MyjrpCRJSr6aQ+hzCVyEEugxEdbU75MiXXVLB1s/iLM1CXzMvRe
Ry9jxgr99xkpHPmNeIzTrLDDHIp3jGdKdO3jml3cG2vsmPHG5VHiYAsKXzZ7TUR+fmk214lPm+PS
jdwdNIB6TYFAe7Uml6ld1dBTDgx6vNHN+9RP7aq4UY3A65V8oMn/dRuvBKNh8lsMsU+h83ov6r4x
PZz5eCGL5rT/uH6MZMcc6mqKs4Uc/nvwA6lGPV4FkSNf+2XTSMr78DHSRXavr8Tq+Rc2+QflaiwZ
4uxLQ/Rr2s9Zglfhu0dHCa2Q3zcY+SjN2AkjpLO0ZE6nNpMVDvTbSeS4SI8qxMHy1adsOpgjpA1A
263bvHKU7bjliLlhoo9MWV82bsKjcwxUzGVh01yE7Lj1qKG/gsomHXO0+/8CIxyCMmlS3k9N+niR
082EPpf98drLCKyljJRbBgh9eEm19L+wGIo6S7Dfhbp17NsKB5c+lSCdZMIydlRYjD9j/2VgFlmS
vVXNpC7lO1EMfoFIS6z6GdiO7yiC4lfy0HYTDPkBPl9jnfcoKzzSjbt6jL8FtySZvuGCelJ+s2WT
LupBTJ4KTxkvqkpwWr5I5AhCWM+g6Iqr4ipYMAanpEIZRZwVvfpw41ZkZGjWYPpOJ2ix0jJFpWAV
+vPL0ej5EkYjS0vcb7eTIlfGkbpitYoJ/Z6/sY4IQapTtNgX/2kNmN7WKwc/tl3bPWAurcaVLbRA
+eFUlLXMVRHuoOZ3zGIIHIGNoW3I64+j6z579bkEyJwCr6n8ptuzaR7o4e2RaAqmHDzM/DyfzHn7
3vMdz49ABixuFrDn9Cf7+lar5sixP8AJbdTwqbLcbEZHKCoDHqC9ZqPhgooeFWs9BvLKWDadwLvr
0DIude4Yx9ZY78kBQk7BP2GRaocfxX5X5EdpXZEdf+BjXPa4BdHudhKssKoUqQWKuYKD234R3pIo
vbqivOoQoaiBySd3mjsNGpClvkubcA8x2x4Q75U9vZcgW3K+3T2+LqpiVjzyW6SShQ60UQqCNZex
SIiNtaCSmC8d3hf9LZsuIWWo/M3hFNYP1tZoNNw9O8OVum+tjBpHOxtrH/9TBGSvqXP3lRbFjVKZ
GL7SF0MRcktn12ZB51FJolBvmJtflSuXFtxuS/I1CTzRhVVRBN4EeuWbRj1Y+4pQC4Pba9ji51l6
3e9HQDp9p82bUOEGYORBvdlhn8O66WS5YS9x22ysjg8h5C46NjlpkdKp2zPbGezVPMY12YiiZFCx
A/vTpYBMNpeq+uLLQiW1KSQzdZuOq4FVMSsys3Nv2KScbhT3lQ7AC2dNAwJLpiD6yB3M97o7Uqn6
WAxsOmxgy5FdK+XWhXPG/TB47fftmN6GXSsn0PnWgDRkOrY0xTkqciwDXZRrxFw9uOk2A5ASzBOX
e74Ld7YxQEfOrSts/fRMwrBhgZ5bkCoJYluwDoK0L7PbWsd3HUFUfJe8frFn/0v8rDdRi9Znpwb+
b+j0Hfiln6qnB6EEhad80QF0OfZWJAtZ3CzJNS8fkmqmH4Z8yNF1I8w2jVIN33lcZuP1IxriMRqp
xdxp+x5AZ3souNvOlaXjgcXVWOBf7xhVz6HAfnfMOFSPDVc+txOl9vY0LLqGYjJBDRlajMaqUn9D
jNfCoVQx0EENoMbSAG2qeHmZ9AsgX59aIfcHleSzpFRlY639RPoLJu2Xae7ybywDIj6fAbcj+mMu
jSv6KZkk2VcL/h76uZzI0kh7D0+Q6u7gOMjfOYi6ucvtKH5dQPAt3cp3F7J8TSGrXIX+crp2hlE9
Y3uhcN1TRfV+6l70h5RC/xn0ueapbfKf+NxNPZviVkHgaoxFbwLLxncTbBBGD9qvFuUxuEYXJMgr
K6fIpLv0Jir2Yk6j/cv3yRl7H1iGGrrcYEC1I2onasgTdS9N5u7OygF7FOFS/K5+D8bzS7LaE35c
G/tFU0ONfkQqWUPGQasro7zR5dSdBuks8ol9v8t1DJXPDKNi3/hO9hz2aHCxMBs9cTfb7mRRFN6f
FD3JZfz8nuRv9TbgVrKGRjgtxLHfGdqE20cbL3HricI7+WKPGmBJD+cgEB9QojbO3loLTzDK0Ju9
5Z5ZdHcbilmuNHGLL7WwE0v8SAu92HxZn1D1gaeJpwxktpE8WUx5bSY0YRj6wWLHjJfWEXuqGo0Z
1ipF7dX6G+J7f1jqWRA9ugy1B2dIj+lRNDu8vbg3AG077pHciZ8TeyO49sjY7bJWmbgBVYTXRVx8
dWeLJogn3kYmrAd8LZvXEsEMWJw68jNOGEl3lsoTH9ceihdM52K63r2odZ7GCmo7W6gng7fCpv66
sIoOdtV2dryMH9f/K+NK4LNMWt1vkCD7Wa1FZULsTuTvG2mMUrIIHcvFrMdT3FkZ/qi9Y13F5wbO
ppPb3TGi59LznfeKlaXSHq1++z4z8HirHXYcdf0+Mbk0GmruJ9iEJrdIFG3p7DDnT4jn2pxjLd3U
/c/D/7wQuvjnfRVf2/RehXqldjguG/J6ACoU//HS9F0F4Fr8tWvjZyCl9x4v3mtJTu3agVXnIKXR
tcJIORzH9lBmkmi75yU923qdxIS14M4CKNletGHOtv/1GkcQAq78UiXMfN4uc8tCRgFdDshP7Qpd
Vu8FPJA+oCizWt+C7ZhOwAKktxyIUBexXG4NT8kf3QbDrTZpbPJ5ys/pNn9wx4/4gbTueNoWy9mW
wXdeNnkYyPpaXwmBvRfkLvbzU4PIm7K1v9ng+HKTcjs4/7GNilo/kQWtJiTfYrt7N6pibq+iexG2
QJupLfaVpsqDL5Ki6cIyI1AyImWjRu4/48voNlOoFOL72X/D2hDWSXBkjXTspVoBbXCJK5OU3AcB
dS2g2duoMWpP1BFGkI0US45D/ITao/h+D29whzXx2kyYYrc8aVCnli00cDN3foQnH/Y70ycF4FWD
OOJV5gi9N0jhvcx/AnurwaAE6c0Rh37PQtdg8uLJ/yZiOXp904fFvtfgXSO4meM0BmZpghiSRhwN
B9w9kxW48fKuQzgfn72CiyBWCHonKW+SmSpwtFuwdFAgUwvdDDrdBX+8r8xkWn106ouNykYU7Crw
p/LnWaLVN6GMQUyI9OCt6kmoN8on3oaq8GxRCcP4l6PdhJVn9tlSIMwX9W1f+9Zm4PiZ2pNs15Hz
pQrFMSycdUV+UaOd+j77F5i97WIB8eWdf67bFQtEDUT+hb3tMgH5T0uBkwNdAM93QHNXQb8nUtjk
1zbO87iYMaQYV2QhhboR5Nh6UrmhM0HeZJbxiKlge2Zb7CjpN7qKUmVRBkAU9om2i6V6B5PIO0dy
ukOsFU2y/Y/PO2pNVRC6UChBLHaTvxYZJWgG5Ks2IIp24gy5sv8pKp7Xjmy4BAKipBG+QaXlxgTn
hEmainoFTP9TM2LT+kLutWZ4uOamYeDyLHjZnL2OfTEuBDOi3S3X/u7AntUTXRRUCt96fbN+eE7m
rxPDQibpgkkd9PsdUWy5J3uX+U8AgRp9NGBO34dnZXC1WnzRwO61DJwSUjDX69pDWnp7yCMmNvZh
ln3LUni3MaxtEMeLWIaqUs/1yKdkryZ5WdJ7waxcX2s3fDIuHOjpiQdfboiZh3Ij5ygP0/PWqTbP
Lxb+xz8u2xMnlX2psPNK3aIqAxQQkEstkFWrA4ZabzgzwN6x0y3YUV1NGamumgNw7p3hYgiDkNGr
sn9c0mNJinzcAALUSlRNVlzVtfrBKYGgxd+PnKV/fQRmC4z7Aek8zBuShpiQfzZAZkZD/2yBP/7V
3IheGz6SOnJqSuDW5tM2jgmhPB8aTvcJYXWThju0A6qyKcn1QO+6teLWCroVO38MFryEDe4K77rL
4VNgJAb22oso9lYHNue3MBPmjfX4STV8a7LNnCVPTGDHjuVqFIu4KyNyoIxvLipvmXvWwQWQ5N7X
hI0h53AhKK51BcfYwqimM63cJPpzSqtvl5rBpfHPcG98pSxlr4zcIrQsFVAfYVXUpXmD3obzD3M4
Xt1BS6N2IYLS2u5cOS6bzXkVBMnEPTUjStoq3hpeLSdvFK+vbEwi2eG4+41M7HJ+Lw7qtklJ3kzd
IPppNzt0fXqbEcjTWvlv+3iLO8ksLytCqcScPTe0sRg+Nmj7GhwXJ1krj+jOMEjGhykugOKh5os0
iSOOSHy6HoZpx1dhmHtDlEM+XZDiHDPtj9QNFYazRNZsrxUUDKkf9gP3OVSOPtSOfnm16w1XYa0W
UTJMr5+bnugOsH6luv6kUN7svNW5EMS7Mpf22tkEoCZf3Uih4wznYPGOIfrDYlTYggC6X2KODw0l
VIr6K7pRKJouGtapet+iBMfxzRDS/2jvDE8AiDX1t/3Aw79qMeDW9+we+HMGvXEYWMrtW9xIDh9n
GJ7mrysyytxSVi97zKFN+cCPZNifSTmYIDdZoTx6YmG3IdX39ZpMgxHCsP73w6q2+tD7DNRXz5ZQ
lOBi9oXNwMnkDi7Wg+ZuUKkQaGyr5qlG0ZOszyVtn8OLb4wvqJM6klMbXM2nkTCWqW/aFKeKlSBz
NVXi9sy7HxGGARC8VpgHc8Rwas2ozccezcfhQld78gUkiScSeCjtQ/Eb9EBnBznZWtncbUOWlRWl
f6lSaQHZcEyOwSA02pCV2JU7o5kvy2igLNa4e68xKnJC/cAL8cCAFQErnHtphZQb4eQwJhK4TEO7
6elLBm5hVHN6+1S9nzLbItG8dcW50LZ9EsIFl+mjcAGaBDwXcpeiph/N6bFirBXYfPzPdDL3xfgs
9YFlKnkINQZPejfN9fK3dHzYhjKLrt9SkEhVrP4iS8kGlvlEx1e3XKPgSJN1l0HmhUwBU+EaeLjR
NgSmAOIQ6VCJ8hXvxNqe7fVefc5kndCqi60lGisKNjwiNMVkSuBKbHe8XzNO0YnIXHqL/q9kUfR3
XJkJsF+ozxHtOL+mf7Vis51ZXSDgqHmhWYoB9yQ4fnXTygeXtkgJtv+uNGVzYqeX/N2ezdmiTrhu
gEq5ckOaHME2Et4Lg3AqcKvVMkWFL2i2eatuEDiI5QYFNmbm4enFAnLMPkXjS4PLvhyQQdulUu6T
2Et6iC8tOPwCfH3/i4FD8j6nu3oK859RBQzPB/+gAGww5r4lecjm2+Iz2wwccFrjsx50lKkVVhZm
tMtXMeS1tlV2CttMK1oJ9WdrTBXlPyslhzL/dMWkwuxTMTnxvvZgF5OQ7+HI7KnzaWxwen9kJcy7
skXWaTD1+d+P/VhfVTkTnSPdp2IsFfgNEBdZjE1ILui13IyeWHj2CV7EHZEVObljmFDt8bQ2avyp
5J3uLra2jAgYoogL6GZef+XvNPIesbaSZpKOvPnMLXX3sb54+tJCBERUVLfR89IELnvyt8SwZPd/
qpP3JZ5cYXplrE0zYZMBbf/gJepuRedp8QoOwOmmf6G4bJ2nBAJg+gvCUEM2WaoRozwWXyHQ3LK/
xEIkDnL30PUSx0cqCBsXL7Vnaf0stI8bTdib4RuDixlx4GUk+C4hEf3wOd9Gwm0WhM4JNtEwLfUl
M3vBxtYL70E7L1BRJ0yr60IslMG77DJYiC4RAz8RYV/8iF+VQqvdymkF165btEzpIu2ESxlozW+W
8G5xkzvNT7QzOHAugZW2KvtUi+8m6M6Jts1NnQ2LEYzCh55CY91mXU5SyieKTs/UjYthj4WbqyFe
Q/p/nzKZqS4M1hklZpscceUpNm0nyi/lmYvSf4yJfiNILSrRLLlbU8gYZXi8+YfaUyL6rU30EZM6
psBaXfFuu+bCSc0LbsVr/UG+w5SzgicMApc8lDSabP1/nffffnKyUqpvrVeUEQ1olS7r0GCAUFqB
HBbbwVySvkpxl3C2oi2WFXzsCCE7LZvbpbB/BLh/8vxHLLGmfAUTD8yV4TcbzzZdTymw1ESY204I
LpNFgdWLqEVRgpcfJ9YMCErF3jA3V9701juvJcfF54pf1/sjenT+fKekSrrYHqZyg0zhRKqNN5kg
KyCBTyg3brE4vevm7KSPsEo6dI/+sA9esuQRNZ4YBxNgOz4eQK8D2vZ/w66miHjU/pIT9PKkDbTt
Wf9Z9/S+tajUEuj/KYnXHIOgTERy95uV+Zv+PKZf46igBlJV3LPgmJ70HqQBOQzaXRx8RIpJPgq1
lDTZAPxyvcRIgAlwC7RNf+F5Z3GBCJ35ghRR34rRLMOxfOJFQ53J2c/znCCtrqkaWBaOPo+tVfyG
xgzGKgSGj5KQefjqUHL9i20Ei9n5hjt8J4/JgfQQdqmV5qelxo3vt9/AdQNyuAaOUQm2ugI8QXZ6
DNXJSuwyX0LjczhD2oCnMwFVWJbOGkncGSCKksGGN5fW5uSeQVNWoID2cXdx0iyaqUN/ya/oDYyo
Yx2OmmMjHzy/aMd5+z6ib61XFk1Yz2u91XL0xKphADq4vXmzWVCDr463KsnVQpNGXkQ5xUv2p54z
JdOnVJbdw+yw+0IWeYzsqrH6Tl58h3ED3NMnqvgCZyk9WF7XT/Ou0qcdtGH/215MkUjeaK2PsjLZ
asTnE20ick6unCeZKkXYaD9UCjDCF4bqvD22szMGoY0ekiw9su8scJ2JEY4IlBCmyimnP4oHTbhI
VoWDOnyaICCdoiYpo4VM8u4HDGyWXhXm7FUpKnZhGom8xA5vYkBlMvF+k38a7M3UfdFaOHtoNhDZ
2daFsHgPvcO8QwS6u1bGnZ0JLtEe2C2GIr3SoyDv2KfCkFFM07KYZLNJ8/45QGE2rEA//QTfdusY
8dG8+3elGidkPZo1wGFrhqtto37FiGzjAiCS1cdk1O7n6M3RG6ujoXuoM4B6OYBxDledB2PlE0J1
SjwjsWskWLymownFu0PJ5a6osHXwbqdbHpGhZpbacrRmO4oNdbabbAdQg6s9izoDr1TA0QZYPHH5
YDnVy7++vYS3ByNl4Tsl07/I4omwKGtMVhOpTDJ+HtzTSisvL+GupGT6KZpjT/cYYW0iW+2nStmg
pAVuk2q7ZvpiwezMcUCCHAtwkqeZ/h5DI4KxvUIbbXuzAHiMBaEsm1iGOm2R42cSh3gy8Om/X1OQ
/F2x85vltgzMEZMpTA4nNVL4kpJTeWiDXwYQif8FrM8jVdI16HmX4qn7GOQn2mn2FPM1Rl6EWv3k
U3gjVCSZ4/JtQZ6s2uyQxcjJ5VqRCcmzyIaL8KtSbHNHmGrmH/QZl1+3pCLS66YOyqmm9qtxQ5oU
H567IuT7upNKvNKU3Eyvz756NY1N1yV5KdIIq279/VHQRk7mAJfgnidrJUML8Ypp7LYdjoBL1gu6
OAHfsY80Yfti6wm3RMLfBrc+Ss7jJuCF9L1kQw/An7thziEdiU/CX3Y2COqZR1eBifHZLzscHVMV
v7euXTOzTWmjyhaAEuzd+EZkshw4qcVh2itx8nP8V0hl/wU7+ZUn6Dw3DKwH5yI3Z9nJpzh2zPWd
Ol+AXa53Mwr2/V40msQz6a65NsxovPXuNkgURY8JeBPfxCp6bVXere8rP8SxjdoNbs9M+mKHktcx
FpKQXOu52d1LuNVBMbqjjdp8PacjO0SNiWDgmVBvpybhzY77H62NKhihXAU3WYnQ0HhymD/HNB4d
wRmDcsp9f+qCrn8qs8y1cJK0SoXWjRi5vbwhHVF/CtqQddt2SupPe/0D0LQtLy1/n1imYhCbZ+Yo
j2IpiTrvxkykGHripU5pvk0y6npOg6Z4eAJHOGJNJLfN9T9r9d/h7Goosmna4RLbiQTkWAaKHOlz
BRVZBvFGoqbbDietrjO7ygpzlsFKavGiKVqABXbKBVGlz/Qr1Qox5aUUfDkxnfkfS4VExyJCeAZw
Z/sAaQpKuAV1lCYHq1xD1A9pa3wEkCp+hbOJl8XvX4w7gyQQ8zTTmuZhjofKNgj7eJxZexJvnr5m
tHaY8fySKVC1AuY0thPNnj5bgpzsS+L6h8UWnMri/CG81j7xGBpn/YmQSum0w2Wc8gUNBZwq0SIg
fo5QvbAWWOh8AnVpChv4+ehsf6+fV+UgTMu71YLpIJA2UGcEvdYYoFfTpCM9K6ydMCwR+3LbWzT6
T92PMmJOrJZy0ZSiZA1oNd6dOzKMADNcKXDHlg/w3jdT6C56Vo4iMjXYSS0l1KS2go2uyNaoyKBn
nzhgXiK+rM5EXGlEKPDSD7YGhHo7cJxdHid+bNZSFBAxz0FTU3cAVP8GyCG0N6AOOI/nzhwywwsv
JB0jRsQ2LCkhXTzHhOs8AItygBRm7I/PwJXB4OFB/wK17ViTlyFdxS4Iz3K8pjHb+2jQHweeztsT
wxh97A1nzyL71d8C2qDMVQQrmLQXFHqQ4n1kJrzNui6O+4K6ySKscJbMFzYOpG8ntRvDl1BenKHU
ggScAGiHqyY40anWK4GuBmmhuftPbg7uG6Umu4PCh8F2q4EuCUXsvQoQC91cWUeoeHcjSesXX7rV
WqHO6iFs2PfhNVk2SdjKjNvqvkgc/7sZ1aI6yOuw1zdoQBDeyEPSRfiHP7T76Kp+1jSFfjLO4UQp
EWKT+X2K1QGSMTdreNRT/EAZ4/5WIbQgBASSc11CmbpE2QrB11oFEJbUW7WwAerxBlIQrP/9YO4O
JHKa1TDF21to8+UopZbabS19+IZaSC+k7ldaLOTr+uq4Piy+u+TtDEVTb6dKbx1aXxrW4jNdxGi7
LKuxQzIol49Z9BfEQULpt7QurfI9/aWQjJZE+vC+zEQI6k/BdE5zsCmzU0DqM23I36M1ixZIN7CL
DjSOmtMKmoOcY1xjXl/AC4CoZmO4SALO2/3vdmbrwOUUisOndA4QkEIffkLj72Osh0nxzVBwN4bl
f+03zv7ZnXCE2tDMWmDIxvi4E8E/R1Y0u3VrIWyQqXiaD+MSyvpd+M0HohMDDhAYLYbZlAAC3DIF
6W2JrGOIXNtQUvLqGbuuGhIjBNecI2CMsK7L26wry8oqo0A7MSueHXNebSHW9goG5X/DIamxS5Ze
LUnIXcqklGuIxLgipDTWi82+M9EzFGspCPyJ5ZF2RE8zwM6p795uQOZQOrjcOSjGewZGLAhaLVHc
tXojY9VblYpytUP+aUiAcjOqWmeHpOFDU3Wn0zxlfHreU2wGSw22a1/gma8j8dA/qHfTuBrKMThS
GsJpRJzx6KbMgAiV50FXVJ2nBGdj22J/HHRqkrGIzilDzWpD01Jt5k2kWCu7WENDt382U2PffNRH
npqGBUTMlNpd7EUVuOOq6PMrzVT3qSMHUAj8yfVq7fhCYEOyzNak0AThVe1lmZ9jTu6JUYvolHRB
cAFYly9VTxIumyVnVLBXJpAeeJZmMiZ4AdrhDm/5PPvrwUfPRBu1iiXUvjewn4At7f0GfLhag/vi
2oor5l3Lxu0TqRdc3wV2SkA+J+3uEyJCmncZAePNP7omKtxJDMuXsATZYN37pJjKt9ajlKRgw0hK
Sfgs7Y6FoTtd5nNu3FwerQnvjITl/O0oFiAiI4byxjE2PlPA/qc0WbMciryHya7rN04tMttLTBjg
jcor/pCnx5szPOtNrbDTSICJU+3nz7KDStDh9QZNu1VNNHotd96dS9CqdWXj8h2RwisoNODLV75M
rbbe3JImzOOlXCg5Dn8FE5l9Dce+cgZga8W6pejAOT4ctX9ieSn8KoNb7AZKcREkxLcEJWYZfAEs
jtksLvNyTofD0wLcBW1vbEAE9ip/c9LPR/kdmQ44LIB3KYeYN/t1tVZsNI/EjskJjTgrgyfk43HX
q1DFjHjE49OAlW9WFg8O5Ag+FuqCGwfdKWt2YjhtXZCOjvrKry0Q6KlYfVuw68M1pZPxBx4l2WLV
BtSqisfeEbw+NhbVTrdmOB/qiU3G/Dxv/jmzkcIkwCT64F3osjmoA8leyIH0OKZ7aP3H9Wcd0i96
v2ja84KP1fKS07Id3A38Jnt8hiHDtmWvkbC6UI8h1re1jvozOTi9K5Caqy569603aUYIRZVrY226
A3CMkhfuGgul2hDXbebVRYrrEEHlPwEQodNwq/d6MD4ClB8UBmKjvdx03beCjq+db1sXy554RBKJ
omlf2AApOE8ctCDhr75Ij80PeozY+sUMXDSKq125oGE/MlX96gp9AXJv5ev2gG9u9RsPX6CzHtbg
5EMnCCGFmBR6cbZ6PUm2tsdLWHXMe8gfydej1CLGxHramls/2w2/XsEdnd6hJBkdP7t8JBGFbj58
eyii08iLpHAA2Hhe/2SMfd2cQRJX6M5exYohFSSKb/c5Y5He20ngDhJaqN8dCa8xqGHWDp07ptYH
0tXpiWimLeERRx6SGH48Fozue8MnrSejZczNh5TUm0m9SqzBcFLZ1woMKXEDyqNZWlpURVdE8XYE
XTzfo470fs66SCLe/8W9pFav5ME41SHO+crrH0raWfYPm+GdhXC41hA6LzeW6QTWe57dvnM0o2fD
fhRkfK/yCRbIeDMpkm/eAScGBmqY3l6dxyW7Z/RQHXkmc9z1Vlc53OzZBElbODf+o8qvX2f0buTA
NMyJ4uwUy0/26sWlkyZL0trhVNFtitilgxfYoGaXNVyP/COFcF7pAb9xKmnGbqdKgZcUbxttqJUf
N2CmthAxgLSjN0pgsrOndraCQli2jelnHHhGH0dAVOfa6WPEOFMtbW7iwSG6Oyr4W4vwP6BRfPuH
T1SAGPqP6OGyKmtxogVSLPzXvHDJTNiMut/egkN5ZtUOkHW78JlwZjtV7xCns1Etk8NCPowt1QWn
FlwRNVDGOpTzREB8ys049BPdRB3AUbNCY7HIgk/uUn2Uh85xtKGErrMeOf7+CFC1JwgG+HrHPDJH
0oinD1sRiwn56QeDvzQCTkwGeDC6LbylusnEe+/Li2rFB7+yJf8LGZ9Hwe6dS6E6lE5vS1ZAKAQe
MNJ4Uzbai1Oc6Z2HmkuuSeAgsyiNGSHqMIS5N5pijuINRuz23I3Ot9U9oZJ5Mn0dW58/8oNJ664p
QJF26H/YvkUsIDQz5ldU7o/S2RG1r39HtqqJQDvR7B8gRCuqp6Xv8CTiodFr+SB7i94T0aZPrzsd
lBw44FhFIbw6t8Wci3SqV55gdlR+BYJPumohvfLnBW5Ohs3WiWqatD0UW5gS93ANH1OBmHHcaVwV
u1fIqsMJLodtlgXZdOYOvGaj8f7gVx05kQpiG0drKr+6QYJPl8L2xhDgqOgGYEtPOiOrz7fxxPkg
he3khAdRErzGRneDuL629NWXvHJZfsYleDaPr9h9aCSRyoi1+l9+w29mylWm/dzfMbmmglkGLlUS
1Z/YXdWmQoreiGxcnsLT3ozTtlA6BznlAelzf1IAfdPb82B8eNMnhbwS9Hkh8vbkUmLyq7r1LBes
8F2EVugFC4ZjK08LZLGFI0W4RXj9EE53zkKq8lHNA3vKhqrxQYF20semfWoC9LQHKLoiJwwSJ6VC
d/WHPyZ6DPygsUHupwJ5tO4oGQWWJYO7N1Wg8tcPwhJ2H6QB1+MR1ZtmwbkVIC2Vjap1P6QJ8/Dp
p4oMmDghNJoIy8YJN+5OBe5p0Nj5b9BV9xLbOjauW5DgZt9QkDnXFX56vPSYxzQo+6ytq9u8vS/J
H9u/DoxcqGkIdZMEww8TuZwpxynVUgoREXDcz2/TD+0t6zPluAMRVQypnDbeSxIdxdsVTMZYEj4n
q0JDV8o9qrEni0xEoqLtTYdk6yvAUw+kcQXnfowGJvAAA1Uqb+FVNAs+pyue02jPrBy3CzxctNov
6wXNw3GZglJa0ip0Fo+SwowX8AlORJZS/lhRFo3DITpnBQmHr+fwxYPlKS6Yn2rEkTY6w4bVgbbY
Ohj7043138S72IVq6jv2H/AIlNiz5rEh988N91bKyrInQmls4leAUCO6W13vO2NYMPziqmrZM7t1
zXh3ZhxpPW6Fgf99yAv6Qy/PtO1D5Tsy8Wx1DffWPvBy60mT3fnfAwfHKxDOsxY8ex5OTDEdnvWD
px+hmQqzWjuAFseVUSen5V1JR6Y7K2uNHqpMZUwm1yNaZIsncjbrsjYO9X186mD9is/Kh8ajt0ka
dFxqR56h4NlyIQ0fvvOhHNPYk2vlk3AP9U15GjWlBn4Es/EWVgy4CZBZKn+jEU9a/GECV79GNyob
VJpsqQt2Tw3OiddSRKADyZE28ofP9Mr0wOR7ydXUa8Vesh+pYUoytz4o0eG/RicNG64XCpMvIwgj
TyN7jqIckfswTxxMegsRcpe0SxDih0Gp/jUDzKJAQ3ehtfSdwjy0KYyWz/2OOOXV4IwULqS1k9/q
zjdMZKD+3Sn285nO6vDeO/6jmv+UMNArx3v36th+Iv60QhOcRDbXkcaMhx6IIEAdaYR2pFTKOXxw
nwNs7DruA6bR+a6GvIfEpTwsWTf5QZNX0ZwRPp1JIuH5H1frracUlcbI5N5SXE8QoevaOTe7QQKG
0mV8/Ut6Bxs0gIrhL6nA9DXSpJ971o5LiozmetWFZzF5A6Z+TS6Hi2SyeN32r2ev5L/HcLCbAums
Gqr7sR/nmBwZM4gkPN2d/M9SqbOr/fthgXS22DbLLXWWLcLF3Oj5r2FGK/FBShrHlzSx4RBpR+kJ
V/0EYHz3F//eYfwbS0TQLGew+CAAjF18a0puWZc1BGIOSudveZCZFaLP6vLgWhJ1eO1uxEF5g0RA
wctzfK/uPCJSKfO4tfdMQncY/qhhwqXuCNS+W30slwEu61mMv2RVFSkLL33Mk7bTrMmaWyid6OCd
Ul0b3aovTuE24dHFph5irg1wKrmvl8AoiVYQKWDn10owHibmifbU+7mqHTGVzoS1zsHDFup1+e7S
deA8huA4NyCEhWFHmkbuxaHdChG8RmgKG+uEcQcF+WrCsjW+KBB3htmtxCl6tviqtIkyUuLOxZwI
Yb3PzU5a3EE6v9HIl14xliD7xPBKhZ5vs2+x4uTBRmh61sDkRpF/6DBwp+rSz8XXZBwmw9omHXRe
1763LRmXIKsWy3aHxy39GvcqvuWWQ5YY/rK72NZ+sHbHJ0y9kvF9WSzThbr99310OhgY1WdBa9Nx
vFkQZpSSIHxK0+gp/tUgLCj5LElDxoKYWW5hoPmbb57l3SOoUT4UqjcwE1z7/4dPPeL9FeKdtwpl
a+7Xb8hdY2Rkrpg1qnWHHQ0K5r8QK46GUhph5+Z38znOI3Ti/YAkvin8HLQed3jpnam4Sh5K+atE
b++5dKi9qhUyyt2rU5793eJUqlfq2cjsHDlsPfpB/I66+nKXJJ5VgJLGUCpC7F6TlRhRsMIm5oui
r7jVa0On/GR8i+LCTPKNzIG4aJdk1uyM9iq2EpWYFn3stNxPWZ/vu7i4ZSShmm3bpRxIx77xwFvP
sfODPhrRv8BFKkrDY4bk2sn5dBDY1W3NndO5Pk6Q0sLHtnxoiwe7KsZfP7YI+7GmV48rPRKAp6cW
SZmP2b68kW+pfdhWDJhIWNOohBoqtwIr4hbGPlxBPnkCsWGoV+udCAYhQnDjLXMoCxlUrlf9osfx
33TjM8Ad9pCjiR/ePmMIQTb8NuwBOhs2kzMgEoOUnKybyUanj/P935dXWbl9SonoJOczlRXeg9PG
/hyKjBVPmvg18Ag+F0Aw6uabsaIg+9ANI5GCHgpsEEQzV7X28HyK9m3Gn9/OfsfhwZkliotPdAIr
KJ4aL/UCxD476reiHkjhYFdRtmfXuwFVZM4pdHQY9a9tf27RzlVXzjDhf58CeK8WZHMegmsRHRTb
OxH3ZCCc9KjxlQTyxnxl9pa2CGMQiahvyexM/rr8JuBXn0YSDNDW/7+uupte88mGYYowUBUcJGOC
NWLtvFcIA1HIinYVfgS4chhha9b+P6Lc+zBQ6qrKzb9Tn0hTu1ZhnFzTGKcwArlzAhkZP+Yke8v6
88NymUikrY4PTr0ZIUDonSegTV8oRwJLJZKvTDznVNGdy7EP2eBJ3fqwjaYRdpEe5vp4HToSSZF5
DUsLsmiVd3VNcXPBlxsQvwzRGRx3LydkTek9LxwtQivDoAmxu8rSHDdgiPQ4wzk6YKXaiHH/z6Ir
RWbnVbUSw1Ohqi6qVQIgt3CxQjQkEdXj2c0jlOb8g43SQ4nvRlU/mm3d18nT5CaM1f6NaW0/tFd4
+jqQrkiTagHgbVy5QyRH01Ag2OTHZHiYUiFdBOGLmm/pF+48qU6WqJfK1331IvCunidNookmsRoh
zBfgq71IJrTmiXttK3LV773NM9JmjQDrKdVAgXbRf45/QCkLXf44LsYlauuDXnh8iSXhcfrmcdLt
ZRHowjn0SoEktwgy0ga2fdm8c6AnekJJ64bcAlWnwAU4LBslaTX92WsA1hXFwfeY42NXBOg70gD7
+o41rVrrHaRrKcX12W1NRMUUdaPnnWFTnOSVy1lRZZ+RYQ82hwUkyCcXJ6KljxW+hJbNe31Famgc
JFFyQnAMDC4vXjGXlGxscLFauLYnaPUCRrvz093gegiaGUCc3fJ59qSevJPeTpvKt21ZoYN+fX5z
KYgpe7NwaP8ujLxfjjQ0V8W3DXDY9g8yk76ZoQ3RJ+QHVw5q0ByiIKgsJJ9ygtnFDbshn4bDxbc+
NnoUFPc1cPPy8liCAc3aaFc12WS7RI/yltES58GgD5e6x74Upy/23zQKGqxvVUi25UFcz/H4N3So
HW+9VPKEtjBWTjjw3hoXFI5oncUaTUTIWlchv1IductY2vXGpf+XqjNaIZWaqRDS8O/ReNJWUYhi
lYj8LfWol2P17A4ZensTjJe7kCZVig7qEh0dty9ZmMjcbDxw6cNlG+fX49W0CPKGdyP3DMdVB2j1
2FWFG9HQncJJEUkm2WE/8+DA3rIIg5C9gtKZ5t+Njn9baQWGjXiYb4GdidHuAuPi1H8FMjOMUQ79
JrHEaFhrxsa+rtjC11TBGj44A1O2S1xtccTPdselwVd8mGfF+oIXp3JfOZv880lFrWnEBlrAI9C/
AnV5kzdCKdDayng2JtE1OgR7Hvf+Wa/SnpF9sfD/Bic9Eo1s+E4sIIBZzyO/b0VgT6VOSm7TpGov
r0RuqG0pv3WvV2oSo3H59NX4BXWuC0DRd0dHXr9QWEGvJeRBWt+aFX1Cxc73LFkCdOoYiR0c0qjZ
/JIz6vuyAKjO5L+KKg6jQjYxf1EFZwSr9RYffDV2G3y8BcnNJOXD2t5NCBG0oqQ/1cXbSzoZ55KE
P2h2AirFt3KfavKKrK8MBZ5MI4gp74J9DduSyzHBIfhaTi5ycqJPgk7JFNLFlWvt+rSS5hbEnuzH
Oh22Bbk7mLv5lNd0JP6QZldc27hDSC+Wz7qeEnF6vHjdcK6oNFzBkK1ywuHeZLcnJfpKKSKib2qZ
SQtSp3SbXO4/Bv3cVXzpJ9ZAVrQOqbJMP7TdghGlW1CzfZa59Gg7S2nyRcAnqXc7t6RslKYUhWec
B1t7KbyywqnQU7CEOF9RKV6N4sZK6CTguX+Tw3IYD9nwJt92vuCztDBcg/46JA8io1pfNb/faSWc
4dD87C8enH58WqjlRkGA2QfxGNa6aVY5sABAwZb2/RvxaWaLZRWOADP7n2uiyC4FhSU+H3pv6j+8
Y/BwuPSGGEvwdoXnFomm9718YdIawBF9cw2lwc7FSs99VU1gORmiALwC8wTxXtN01EzjnO94vIwd
e0M61aMJqlxkFBOVTYC9U+b82YzOV1FEVDl4wRR/AWRN6mxLcemtqle7MR5s45Ul9G2LLDAJw9Ri
otFf/M581I3uz5vigP1xcfV3MJ4+dteFy5FL3KO6gF+YL7rFc9t7Gshv/TrwkaBDh0W5iTqn0zd0
OI/03IeXGVi+hXH75FT1w8XTLK7TsRWsYcfLQY36KyeGtJingzqBewus/w/hRan8UOoJBhC8X8dP
iPhvcHk9k5V+pX5aylzaAEHDVYMMY/e98H93TOpDPCXnPH3J1IQjQrV6ZdklmZr+s7OO2CPhFZwX
Rk1hKxgGvMYEdsUUwdp/fFkkDYX9GBRblbFkEdLLpIcMmOedgizl8tDORyWSGdfkjNqMi2Or6kIJ
wrSl408NmMHDtA2dZUhNcPbswDLZNqnM/7vhPiga2pYo3R2uiojgeFShBNqckQUFdIKqWtbx8Jcl
ZjoUwIz6/oTGNoq+ZuaCq2U+2T5bQ5zXVyGEvXKh7qLy95iPnoQLO/VgPK/pI1VstJJ7U71/2Two
5IAfXOuTsO9176jC6YujX2tbfcw/qS+cKKroayRSkIKFD7e0wHahbwXfEav/tZaXl4MDJrN3qYRG
u3IpiCNavXZDbkSXxYJuYzNtNZMY+gwa8pS7J3U+TkuvuI1ljnHrg/1TA4kP/3AvZxQqC/5NECEe
wRwDTBtSsvwexLU4sJJtcSQGDCdicy596/Znqay4wlqExIhT6ig45oLn4LJ/QdG2l21jiL3uUgsa
KWCKBOIPvkrd8dP5QFz+6eK6zpV8XQXfedAwWHzlpRNr3LAh4IWuhtZEo71LKCQ8cb+A3qtznqkm
lJ68xUqA0J12Aa3H1aQHcDP4Px54+aWp49yD1eh5dsB9tSdrjo2d9vYIbp9dyae5FAh9EIB5hkd9
vJE/uR5b08KwIo9z1vaIzhsHLAREsT5tOmPlm6+GxHh+RbLBpZZKVaBwZwrxpkwxSTogw5uPP23y
TnH+NCG+QeVtpoO+46ht9K6glMm0Nj//zgeInz4gTTmsz+A5ttNafBm4Fd2yxhGRwzthJdQod8Vj
LIZrZMITZqfD6KYEo0D4X8AF8pRzAbLDASvQ1I2GVcAM/Bq81ZyHn2QJPJoHwLaxoGuqwLd9xoGL
phmRJ1rCr9gXIFoixh6A2rn4TeZuOcMYvZa3yWnGFu2DcWdDckCiHW/khWWnq2C9cosz4Bx/xjjS
ACqm/n+ApRvZmB6Zqpb8GwFgdQyO1foSyHiMQ4smXLzY8OV+X+jB30sGbvObQ+J4X1bTGUlq+Fe+
ZxFGp3L0sJd43yfY6b0hWwysLtKtf4ZpW4NNcRhnRTsVWHxu+lnoeUaqBLDdSoWEzykCpqtsVo4v
hoXlDK5hJHddxCMPJA+/WracFRKv4uFo2nPE06DBdxjgZFOuE+CT2EVZpc/XcPplrGmSPPSdRof3
jg0WS4kGOuQcGPBxdu8Aikolwbg5x1cQu6OEkUg1OmZ9vT9XX0RV/ToBq3d38Td6WJmPvdWnctbG
AXc8+ULI2pZtT+FUwCdLo1ygJdC3R475qlQhlTAJdpcqERO3Z8aaOF2QlDZzPbbkvhdh+FsIIsPS
fFIlvSjpRioxwwz57NpSdO2QGqBFAGyAtZ8zgm/OOOpRTSXdflRykPUzD5b63rirnmTfMRtOebH+
mdX/bz+jyfKUYVIxRvyKnoXMsYhjMnN6X3paWYx4uskcD8w6IEb5wi434u0AWD1nKSoSfhZosPG3
LWwkyVV2mGZXwjXbVDaGcVZwikSPVOT16StyssultmNAycBG01tbgaZINj4uRWJBuYYkRNfZDLGg
1X7hd1p7FkpnDhSIj3RIM07qMPHpzgVXA6gB/CwhtXeX8cfDZUXMaIV5TElAgaPXe/BWufsySFDy
tw4DgOPOT23pyZxcVE/FC1oHuBBkNr90NsegqixbCxxkL+xVw6ZoXtmRiueARiygIolEF4zZouWZ
CBToHQ+Bv1BqF3M/timCeEiSdEPBl6lflsewEssj2f92fLa/jY8lvGDsM8Jb2DJpiTUQzQdWnMEm
UCKbeEtB8b3ez7+FxzFvMdF8sy8QeBdA72ZMnKc/iDBnqzA8SFc+IwsFbxqxsIhuTiWcAsJB2sa6
4/ix+XKpOfGAyYb+KFsMTqlBzFONf7e/oQKSEvWzfy9M4NxxIjrmWUSrM7/SthVC1Xt7TaVliSK6
ic/FJjzP9fSxQLy9mP56/2vuK4dt1Tkp7NarewD7aFX9RjajybQptAFXfs8X3G0yx3ZgC9cwB4/f
3DYmyOpBj5nsoev4qfPInCt66V12t1SSF967q7XS6/rh6LYB6X4FjA9r4Uc6fuM0rzUnoxYlePbC
qTZy0OfM1JLLbtxxEkYhYFWsxOeau6rugaW932eAFsLw+rKkOCGxd0eVCtBO/4rSzAEvrCLgWnQS
xA2K6ZFk0nTfNgmVsLNtj1jzFP0g+SPwA08wIDyQE0ifohagsfwPHkj580Lecw9dZTe2Rc90ixHJ
/00cq6b1mWulToZNnNqivtr5kGAUtzD6FLauT1I2Y2YH7lv+0wYZVBQ8U3WOxSmapvykf6O5eXXo
sHwWjvovzRhRH9B1CLQTY12dmilLMFyQZl+wyIqmeyIR+19khOISi8r4FM1N9JmZa2hRnfoYCFtF
94nIefoGERG93uRNkcP+oQJI2C+74jUZb6OAMIKklXcOpnaGl7u3bbeL+UiK/IEKdqk6MPOuEyVE
i9JJPSBzWlPYJolo+e6IxrXFxNBahJ+G3UG9ul/+hsr4N8ln9IgeNPKYkC2iuEUKrnRccWjIZ7zU
MMBrt81unWDNmXm6Z0qi/289gmUo2qzzWMaZDb5L69cuBDzeatKgbw4DEExQggK52LoMJ608h/+D
DPWF8j0wekh8EfTQIagPVXM/PyINBxwPYPpDfkid+ap1aQ1Wnhfoh9zALG90G4OV1Gtt15Ct4x8l
toCcNvws7TD/56mC0yLAtTuxUzG4TAITotE9usgqQKK5/CbQgkxnhOn5qZJUvtTEE2a8H0xrQvSt
JL9oKAPqgRWwuGAqYX/wKepRuaWhZXINBcLMeTn0yW2xM5tTfk9JE8MHGj4TkyVeVI6B9rXpJBw/
7FN4CBLk9QUtkPh/c0DIaGXFvVQq8qQBuGiopZ4Q0ZtGy0rLxxW72d2aEzKArAMZ6Ct1t/YtMoRp
9CpI/vfIYpaRrx7/OI5hbbBpgo3aDE6Ru1UqKgI6MKl1+w05ymue8VC5CGHNxhZa8mclnfO3Xu7+
daP+JLozRg2znNVK0uW1rf1ZiYsS6dCY3D2hkw4J9LNIlVtn5s1BceQmhKCShtHvouVeSeuO5aKY
xJ7PTZw0h1P7DC2MwTr+UN1dyNQkTDQisT9i3OFrV/Qj6PEu9mA6gOQ0nX86inyI9yS7uinD4klp
yJfknm7CHEjnmqjQzefo+GEJI8rzc9yclpUj2j+0BEPG5WhCzVI6v0ihLW7akRWrRb3PRHiVpjwd
g8kTx4jOaJocMS5A+ziGFreE7r+MZ1dqpTAeyzV+ITarPLw3p8mVxd5hYagkwH6LHlV7s3kYU03i
bjyX3x+nrE7lfSoUNETu64j9IfYIo04zykr6OnlwRiNzPT/FthCQ2KwtBmOGQCgaYk1ElritdbLU
3zmOfB5Dnr07tbNAiHqmV5M1YEJUtOtrXocIBwAiW6CEEJMcH2/gVL+kV58Ck3pcue7awHoI9y9b
HnzYofwcKB31D8EzYh9mec5NEyNJNkCvV8Mr/EXFEPvNElYj8umQdYwraCaBLzh7pMsJc2AP47z5
mAKoyfkWB2RudbU85cDwI/I8kPKdFiWe9ORGVOzubO7CLqG0pMpAdXbz7EIjzYOxJhieJA0FobRs
cDtN9W1xhe3EtRJCsoUP6x476F9eme73mRtiFOZhfE1l+hRVlL3aPagkpa/XTd6aFI1bZJmJyO1c
5zJDFjC12oH2qOLOfyWS3SU4HoUEVzqo0nI39iLKePtUrdsXEcJSUlqvotGFzsiUQrVxjUtIDG08
YNKoFLK9dwHwwseCigOLdm8Wy/FnUe903E8JRseguURBBOE7cA7fBDZAxuQZUcqyg7NYaoRWS7Ma
tCRH4mlbQ8CDGlT/pGR/zwM8KNxDp9EXd7VcQNsi77cW2zS+TPtbpsJyLfixTmkuB9AuTXQImDWd
g86WLWlPF/qx/YE18vDN7Z/tquWiCPJDobOfnzGZSPspKnEndbNSLO20q8URMucTK4oCCd0DCKJK
jsSV2hUTlGj1YMLWNrGIc+QElkuvLdSh13MaiRagolZ44HNFh+F8GWbxlXBm+de4bE5VhWBFeCTR
heH2hB65e79Q2G3cnkkDswrkHaKs0TLBgneMT/kg/8r025hzF3QPBgxG7GBx5Vy0ku8nIqDFf6Lx
wdj/Ms2SNb6y3h9UhLr98E862Ei9sYVm5pjxryqjXKYPw5Icx2OuU3HCo+B4tGYcAHTjad7Ax0gE
uY1HtzbyZf7CzqEElokMS5Gy0jkZ+y54ysWnvj9ULRhuLHuHGzaAApMAuKqMIN1r7snrcNIVbWNx
BWtvxedSUnfjAaKMZJxjUcdtdyB4SG2cpiUnPoDPP1ccMTL5KTfkhK1Z2ncbUAUMHwrMxCRcvm8r
Q839lDCXNJzrMbekHx+RazCooOf8U0KdHdqof+PKkbHpLGdJrR3mKFN/fary2yQZc7EJPtjhYq5i
y9MzYLbYwNIEbAzmhqoNNkBSqtIb1aNsBbbYCHpWlY83oRgkgCeanJaUpZkkOZ0YigESad5Re35p
uW1CUf6KSrF05g7bq7YvunQBXevVMEFg5uyLmd7w0CAMImPwE+Teg5fpChiJRenvOsvmB2oruScU
pheN6qe11BRJy4lBg0qq5PEs8PEMVked6X86uKDCd+Qi8JRavoVsNJuMQDvBtCBMJTlekoxCYceb
TmeJroWcFopWReonR7Oa9QXLwYarzYT5ZO2rUIeWo6Hp8S2F2TGgUMDiJUJ2e6zA9DMIZF8a0d3l
LWSBaIBuxegjq/B68sAYlkdLTQKXcyS7+vhTqvwpCagUOflyOZqnA+OloEbfnAWsZWC/4rQfuMO3
pNosfdt98VhTeiGw5dmSdgAnD5aKhk2MkhnWhulYrK7eilrDnTV8wuQ83PgkygJcyNlwM9m+WNdw
JdHvxOvIe1gEiq2Xu65iVp9sEuzwvqI1qyeLyxM4WBciXC+eZ07qnH9Z7lKoZEgjM6FzdmiJ7wwt
AG14+2Kjmt2947S4aGHPjieHgQCNXeNS/8fVMEtOTkswPTYwVQ2E6CZOhEm77SyyBHddSUw0iLYK
qr9+tVnTgqd/pYWvv7cEROPbu4hantmuI/y9zpsuYGxzGzFI5wLuu3deFJHHfssH0VAtI+hOWTQb
rvYpxkP3hfRxpBza8/2zU2XtrMQVTJgEsx6qn7B12I7aNVg5abe6R7HTZ7mZj5su7XRRgK4wxa8F
Xn9hT/QOT8SNF+Fryu+lpZOYpA8htJDXkZEk7uybx1Dlo8K/ClL+CjQ6MM8nPmpRVuJxyuIDO/e7
BUK/CkQoEYDUVJHKprRK28HmRaQGg3mPkvaPCdQmGkKSBCv5UmCDzq9M8WCyqlndHtlnHBfJEDdG
deNhdc8pTntpPuROGHcmbfBpnedc5+u4nfl6Ckiu61GNeIvzmiQ3eCLVYwPXGT5LrJ3OjtG0A5bt
NsULmYHtYtdfC+yxjC3ujMH5l8w3xVZfmgcC+krct1qj5AKvcy29k6ar0wSPeu8pr+CpGwVj0G9y
8DJu6uosi5OgyknEfMkxY+ue1fWfSH383BwSyJ+kxIF1I1B2FlZyRXJACL4A0RkTwnd1mXONALpK
mKFGY51s9nDQsk3WuowTmK4kdJnSe2IIEGEIDeSBCiDakL3BBnHb3hj2R4Pze2KXrCDbBb3++x9L
HmJehl54G/FBw2c6Tu079fc+HmMew2uh2rl2OdorhmnMQbvdOdwJBRJVwvfVBQpN0ZHotIhCFWeQ
4w0xmzieYl4CtmLSbiFmhYx7OOEGPLhmUctWibZ0ZDLnXrljyap8PLkE+ZpWlvGh03ZK9PtLzEJy
bG5AW8WIUhc2QSy1LZ3kgG6F1Yq3Y25vMjFCNY9lGILxCmEaw/FmW+J4+t1AtkX5u9TEgUFP4AJ5
LfF0WrlYfHWBUA8QB7rL0LWNmJgjsA7GAHt1RwE3kdPe3VuHeQ59BZ6IxH9TWBlMerMKJqueuwUy
C+xx5W1D+MVWpokJsc9dC/h/y8qJt1f5uOAR7HxmPc2sIwNFmZDATLyDyQmke+lVmwtbXGBmkCYr
WQqQiJ856UhX4Dt9bXm+nX8IQrzpznoIEMW8L6pwVdnMtPFxIsE1ivim4lY3qQpMxJLcVhTQbw7W
yNusrRvK/Y6djl/AxUBDZ4P59gp+vHXpIeX94O/KypEwKvYb2Bv7jyYyDRXYItuZUJsvfCZXgWwX
aQZxkFSNgbRgprOOtyfAUMPUwqH1voYwPQHdtbze1FMXIYZK6erQXrlinymHS/72i525/1EakziD
AAbD1N0uMOJ5thKihVdtiiEgGDSQgSHe/mmUYCoWfOkQ+PsiM/3EBaMuKvrheMrzKPaWskPZwtVh
Zlm0HQW3teE/m7HBLBlD5DtB3YpVYcGOZUVaEuSO9tg0tUo+EPJLT/d6exOjURKwvEzN2Lvh/qa3
E4rApaxE89R19DV+/HfU52IS3dbdTxCwJBHI01u2/qjh7T+AGd7XR4mXt0jbP1qNPlQdSyWx+k4b
q1cQjZAEMYgdQzm3sslxe/77kTyknpiEa9ZpTXONBUBj9wDuSlKK6J1Lu0Ew9aszmYDXgYZgQaUP
JzCl6GKWmoqK9Zw1ioGkD8TYgcM0UO9nQCBK1xn6jK7nKT2jFvCcy9OkfISCfHmtXzelC9cKLE1V
Mn767DKAwbiz3bV9xyQdmSqrGoTm42v2bYsIqMGfK13NfRVmB8eoWLMq0+w+s9AYwMCB/+3hVHoO
Q2biFQ6MX4MGkH85gpw6Y2EFj9PLxTPcaewiGmEY52u9seNYGiYj+jbeI6LULjc1gvvn69gmvvtC
odnlMEXp/w9WeiR90Uts5DPTblxoSQlcFa+dKGegT/o2LT3bDahkg/LQHSccnjBg7X8lD4R4uwsb
PZxKeevInLoHDgE2MO1T+CVNrcL0tpmGypJzS4xhXLGL1M1v90YnHyA2CX+vo8T7G0JmYL8vgqzv
YiHBQ3zylk4+ExZqem/WvCQNvDfwK1hvJSzYKK2fTNsfaeZBvo/VK2daIU92zIjeiLG7WT0mrkTS
fW44ExN9iYy3QXhpMJ39VCDaPaefttjgxx4J0DwysXxWmzyXiWVeprakA1QPfMeKBiimF5V85U5x
cms4OVPMjkkh8L3AiElmVoXBMR1Jx7EJcACAOlPEPplye29RFGgHXGLdeXp4JMX1k50tKviPl7UB
ZyDJSmW47CqDLG2TbZkxCPEc0AuRu6AN5vFK8nOjHfn5TRxjfbQAgE4UztdYEi0t09qY7IOnUlYh
rhfRaPdZ9lfZ4CADJGjT3XlzQnovho0AAWeYYixNftdU3ztiLjQKnvz1pRUQNPc321KC0z+k1y/N
WbIdHEkVYsVs3n4lkAf0jjVhMwd69pnUxwHYDoJ8IXrrlNX36k8WMjEaSguGtWbe76xy/I5uN1mL
kFQHecEP7Y0ETH5RJDgJD29fmsaI4WYI003tKqVCjgFVhBec077NLP5NZF3E7FXMtf9PcCtRyMZ4
zJ0OCFEfbOqDH25M8qOtGoiJiqjODZ7Gbv7222DaAc1Pmdiv/40jzhvCQm1PTvHzbUBIghrSxVb5
LtD1QVsnjpPO4t7B7Gt/7KmY8niNwe6Ew4kevc7WWCARStBbn9nVHge7im4Y9grUVOpqzq4kQNRU
k2agh09fWIkGUChLKTD84+tOVDp1kp2mzUJcnvyQdvoLTR2V0HABO9vIQF/gfuNXKvpiLstI0vtj
V/qK4ccbLo/wOOjSGPkFGWjUiDLjVIqMRzrO1nDeyzoOqOL7jvnnuWUK0Nz+8FjzO4TqKa6zjT27
/p9xqzXX6YnAsuulH/o5C0f3fWcDyK3zLWPSpu+RmLCEE7v2TTsWQkjed20v4nDDlogGs6ez/Bn4
zW3YOuNobrg1jJJBfqik7d9oaSOS4KgY8VwSaeikdgC2ZqRXrvrr2f0hR/secCpXnbnhBruo6oea
0sXEA6xI/SkZ+eEVAdnph/cJC5KOpQV22/2yHf5oyWXSi7NvAipBbE8nNqGW7ngjGl7dF1QSUeDP
bd+z+epoGeheFtks3kTuRNsLdp1OD7zTuGb5eJ4FjfhVhEkGhYmeKOXrJ6PXx6t768I3o/77I3oh
Aecl5X8gJkifi54hgYjImJRMdeUihA4eDMC89nP9VJQsE6DBg7DC6bOnY56r36+MAQcKbzC4LxM6
6wfEcef8kF+ZC7TdFwE0OO+EnK860j55vxl1Al9KPnOIjN6hLfZHH8KFJmLaYsMYHqdUWAHQN/Dh
nitVEqRK450AQvQHGzt/P/JDAorMNcLbM6NHEPnEXAlYsMnKE77bxSc8ZxguuhhXXak1p69BvT/j
+XbYdHbBCnWj/IT76+9sniORmxVHUUPO3PnrYs3pbqktkLbw0ON9VxwASp6qbCecnRycp5kPSd7i
rgYlTDIOk16Pd4cas75d+h0As8Qu7R5j1dRqcunlSYFzVnWEND5Dp9p1r70fi7Le58gf11jwnRKO
YNu/aiKZAfDaoOEadTrxxKtsj0+aA0JjWeO4gnHoGLMb4j092VdCuJIk3jhKo455vxQHnfFqY1AH
Domp3udA1RczGsX1+ORPF4Uw5ABcHkrrcSXDM0v+foLn9KTwpO6v9H3IJZynlmZzQgzuwhEye9py
JEgWogHZrHzPDC4p34PW2nODKbpe9yGtm4gWVO8IP1OEjDrswmj8hsc6du9XB3abbyEUkxlNjYnC
yxmWonB9+bP0uXuJe/0E07tVS25H0y+ThNrqe1mb8NCaB08AGew57afyQgsOo8r5wMb+x24hRqau
0XaJClGvIcdP+Ivi1ZBauKXsti/O33O3TlRsh9qyCPDmX592tnnmcbwLESvegxHIeyqQNM1A42A6
qjN98u0lGf8CSpd2ij73F/0VIdu2nomSuFQYdruGbUopAH6e+Uwl/Tp1eQncciFrLCVcR+NzXo0N
BV//oW73Z6laEJD2Lw4glCQ3i00bOqjdRYRt7A9nHZC/hqxUDx/0idgGtuzcjeU5Ulmdrf311gjl
VvFDVHPO+TpAEc94LvZrq1ArE5mLfT3C1U00uYPOIbxTmdeP97Qa+hrI85rOOLpjmkwh9KQJ+m/N
KklP6CI1I1usG2fWsGbTxqNJVfuBdJId1GypWPpATYmGqBx9Ui+GEABCSS5j2L3MA5VcwS5Wtnec
fxe+nStmPzBqBLlwxAJKE2IBxXnC3RShQz8lzMHnOItwykEb6dOVLGjAUdo37KQg29ARRuoKhrC7
vd5Dxk/jxvV+eD+tVy4GM3qe59hNm3QML3ANbCf0c8ldCSeqwiXBJq1QYcYyJy0az3GsBfRH6rND
Hto0JyXySzKtPL3GclbliP9+dv7pLnkpLfLnlgLHJIE6uU2JBHis1EfQOIGGdbTWjeDXd7oxIHsC
Wnuz/f7CoIN/YwsKGuNkpx5N+Ti7i8/aqdCTMkBisso43k9RCdJK5CkT9gUixw3azdaj0BEDO+MI
j/tmkQyl+nVgffxpfVlu3ZPfcpupKHgCiASl+JWWtVoW/BCjLRJVKhu5s3NmnYdldJNTYX5f4pCS
LCIa1SEI/cRt93ItLFRlcL2pLukoRBXht1oXEr+vGuHWJ61u+b5QisGtWAsZ4JWSPVE9PIjyqvNO
5q4cN0jedqpnJk1sImu/CyOwNQYGsb+ZH6oZMGBsIBD3oaMxPYwR/GmZt8NbM5D8TDWQkSrBV3Vc
KZJY/AVFGd0HRkHsahc0DIQfz6zBnYNsyySL4B6YFvhvfe6ZfC//ew24i8czPw35WhdAn9iG/sZ6
NFMe8eq02IHh/AOiZJt6XKJ9MlzBGx9ggeNIkACzR50AwqVikjDfPtCAdPaN+RjvDjF+JoRGNXVF
psYz/mcpE2szCmy8sCOGUdr+EX/RZ/MqK5pbbejv1vulh1glJ/Damuew74N5x5qiuMiwj6UG718L
e0DPGur6TIWQdpYRwk3RwfMYSGRRzMcmbXH6bQyt+zv3fM0F/4V6cB74Emc0xWMMIS0KhOMKnO/i
eyAkJM6/k/dAjj3BQBgFvcJTJaHM08y9Ec+fz/8mdr92H+Pj4PCqlLIvlikuQMsTJ0IyNAXBTpGa
l22lCyqkQBfQmv1L96UlLvCSBILiUewhqvLF2OmHe571I2hLnaaMMsXQcBvndc6spKswPxuxzQu2
R7ibpnpKQEPGam62bSXoPkO99FA5j7GEZr+FldRCh8Do6eQSLkZUO+/ZXUdCEX31SjN9xymocb7g
pYs9yFbHpfPec61iBI4wqzPHVj2i4O4pDruHdBlRSgmyUyvq8aousBOIfIQ3RsY6Gjub4EVxh432
x8knPJ+vGbdzdLOZckb/loFyE6ABnS5Cv1bi4Ti5avhdux0cfQ/IxNdlW10tiR0ptepCtfozjdHI
dUPGh+l+SYcmslAP12ToTGXTAb/5o0iG91TGxuuWoT9HFaRV/HvCUJrwCr0TE7c3NlpESRT07xB7
8TjofkCBWt1UQ/9XeWLMEV5MjcIpDqIaeCCcWlJsq6b4MOCahIAsiFOdLuQhgfDBBnvBiEQ5VuUC
y/hn8SQmWdYJ+nozj+gYTGGBoJsudr3iPsqtEkTBFRV6+qF3FpitERXo73oked6IEvJyqK52F51h
grl5iVd5leb0j1Q50iRUZp8rr9Jy/IdMxY4qiZ6RPEK1LolejeWXlCePppqAuiJ7qJF19VrY86aF
iK6P/5h6sy+0yl+Rbc2i3BCDt9VYd/G0p5RXoWsiwmDIGyFceA8GmKkkFs9J3IBgBeMIWN3IGVGP
qrNY2E2cpY8i0EgMxH99cKKCSZDd3f358OOe3uJFkxkjtDsAVA/oL4q7lBqZ7SGYJQgnxsq+qpZs
f6FGKgCr5qBsLd5Z2a3gf2If5KSgmHRAVsFI+RT8Ir3yl3SaRaEZLm/N3ZzdZZbodrwsugBACxTQ
M2VQHGH/fAU68rcml+r5B0+sDZHYOLZkyAcDgwmcqJxHgxV9qVRPvIIb/LKs59BHu31wID2V+F4u
j8zmtTjwLNAPsTgBRFQSOSXn5GTU3CYIuIjD2x3xZsWLM0TLntKFvptIMyFrp8UlK9lUPO6MzjCP
JLzyPaT1eRLOxTs2i/eB2TN+SsAHHvvuvL2tq/3NlkwkJpjNLiLH5IC6Fq7kj5AqkLVBS9OqV/T0
lcS4Xe4AHKA6f7/TATK9M4mkJrDLuxtuYD3fclMVOVK6c9XQAWrkzW/uEGoxUDpKyk0zriMD+5ky
cIrmptbOgX6Kh4MuWfZL7DXwiyV3x5Ul/kHZ7PY2IFXYkB5XfSuxYqPwQ6Lq6ku+VF1E/UZG4iss
TUmGq1J0Iw18m+PErLqsrb0hEM8/R6lQO4iIzTjzeWUadwlYcbGmgeIcx+f06OpA6T5BaSxtfsMH
1kheBny4wLYvDGRo/aStC6onLGzG/vQfbWDBLUEIERkoio3t4RjIVOWqfTx4yHzuHLSQu/sLR3fT
748BhESC9s9BBRYHf16OyLjI0ZxlofoAKX7jehsJ7Wx34ewnkNq2O39YJ15XNqfebWqkG8OBpx5+
Uo7I7ZFm5U9P/V+ZPvpftYvIDM4i1nrMpDuVvzGZIG6RDNg+hCLzbuyHvRYfX5FUu7T+Lm2vRbwI
nF9wL9JxvJ9vMb6n3enEhzdL/LiybPas1cUEX1JzH0cG39+Qa/JZ1A7tbTl9AaANqNwDikHFek6N
ujQ6QCXCMPDacUb+iK9jrwVuiVALPx21lj2XRiZ0Oy0a6yzqNeWZK1S1+3Xjl1XsXs/mR/meW2DX
CeL/KitgZhWw723/2EAeZLmJGSjDDyR2wZ9oscVIUwy9+p1HDCzNPYZDq09lqLc6eQ1JjHHrWFZA
rx5yjNPqN214dezMUKhQRUNhwVntbWGiq0oHHOGR4PrOGGqwZptvilt1WN4bFus1x7FUa4vPiBtG
qiWNGdI1DEp1a+cvYPCu6tNZZY3LBHDUnlIKyDNNmC6dxaR/2h31rZ4P2qpasWBikv7oE+VEnPe1
gihdDwaAeTVFvGSh88KTdqtUMqwHWSoPQOByw0NAKI8dA1IriPpludpwk68ziBU2fegb/cRYT/qa
q3Wn4nGh2v6EUhMuKTRki1Dg3GiVkZ1rOevcLA2gR5bZjvK6JH7hqDixXrVUJ5bwum7j/19cRmlL
WvX4G/LG39lymA4i7DIZulViwWb2EEGdbVJG/FjVzPpRq6f7lb5XLCFq9Tx+pslsrJD4DbF9yiaI
SK9xX85Xcm1BqqJGW7DtlPJ7cUiSR2afyDfPYkleb2CxmGDAVwHR6sMvJJDrr9PThUlyyrwUsGxU
AyeEFTu4zDRU/zoh95zryeYAWUqY6cHhCUYdLtTh42QKUbHIWkuqFRPpR9MTkNpiIWxUV8jJtnvc
F5ZkrZv3wpaC3ZQeMODGw+IMsoiopldgo3IvC6gwTRBtQffWDNrGIe1TLL7jQungVVlC5REvf1Fq
+0KHwRMdOZfEWUbT+Es+FhqZ929s3crkoO05j8ETXSTg2aIUjuU/xtrtS1eEzItZ2v6Ovn+fcTt2
TxTJDGvRTi9l4pU7W47IygTpNOLx7lTChN+wLA8OLrMeNXrX3EOU+3iLGKvF+SEkh/G1aiDb3CJp
7yp+q1EqqmPER/wkI698j3xVn8yy2Xd9wBXxqAyU3r10HF9B319Gwh0waP1gvcQirEmlt2NhK3G4
8hQpZ8XRmKZfpCsWklbPzn5tcAa0/gh1zAsiDO+5IRDd/haJB0sa/0hsm0HrCCQkzQPnb6B+8XbY
hdgNpgD2ZlZh87Dv3lOzmhK89mW/dSc6q5NGh/VvHq11ht374o2NiIP/C5PrkHCt4PqERagD+DoX
Xz2iqHm/BvvgMo+G082kgWyK4yRxNXf6XYEJlQUh/UqtWaW3BLJygdFLr44TIhddAlC0jOCq/XqZ
z3kVIv9dQWGRnWNaizhLMV74ImKq0gegoJ/05F7/b2XMAPteseYLzXRNAKuh59tz0lwV7s9H58RH
WxPbl7k8A8qynzwSZQh9Pnfwaw0eFzU9HezDsYSgf2BaQGkb+Khyc3DwPyPOEG/WP2l21NicbsF+
pDJyEfYPAQ8p0ZSlmPvJkqtVmbgXELZGS3cYsSJbhlXKiiG41phcM+yvraAjWB9LGVO5uszhPQWp
B+p9jNCwjskjwdD7USz1C7G1GfT8lB4tWcE2b1N1B7f2h3/BRA4adYXXpkG/s+UqrDk9XVciYqJu
6FEbWkPtcW1BZAbg1GKPEWOMy+8JxOMRxW3bEpNAFGmX1aLJE7EKma6Dn4yueUe83JRAfNuZcMBA
SxXwzsMnyMJVk4cZ0eTla6hdfmTQb3PcjZaceSCohRjn4zQrSsBvdLyKtVuDuqrGOtsgidMYWdF4
sSbuOb1ZjPG2yt/vM5qPDEzbLzzyOQ7095Hr9P6CHJ42DHLeOhWezB3dfbI2mfBTZmJCYhiBe3wN
Blmzp6xElW6fSyC3ca4Re+dOr6kJE8pfVP1n6MfcQbqRl9Dzxvbbi8qI/+58AIaSTAc1w9FxN+Bk
dcRB+hrtNlgAgmeObGxV0hiCSmoW6nM83iVzyQN0Tzr0Ruz+J1SdbqYLjBdIV3vCCrvikTmMWwwd
mCvWDwyq9SHqIID4F6CSsVEkGgDPQbD0dFGZN45exi950A3iUcznyLgsr0l8bGGcuG6FzIWtyJE4
wOc0J3lYEsK12uDBXb589xcB/9iqhapP5cOX/R8w6ogpI6tcd3QbSZQgvMWZ6h+jAZwPSOgPRKpC
ruKV5ZBSOPtOdVYqwwqusy3xjOE5AuHfUP6cNzAyNK/aWy0I9+tmFTfRU3fVIJ1QgcNNCOZSInnE
Lj6I4Vw5/VVFIW5wQffxLbTaHvLew+GegVwVLgkBfpkFHXTun5UqpCu/oJppNFESoYkx7PnPJWA2
/H2Yccq60b+WGRtajUKfHfj4W46+gcB3bWIY3KCyQwuB43/6rSVcJUlfkAHYEUyDy0ydxxF3Vzsu
T3ZHkxVa3PurWTanVO2TDyieunikhpEeGE2HFh5DPkRDFC9/49ntul5sP5ijkK1qyBz6+oWJA+hk
ZibJH0zUAiyk8mZorh01cgMflxyBaRmhy6z5oqOl1xohhtzYv3ssWAInr4BJ0W6AYd0ZciK+FJPa
IwY19SstALSuyqt3hTS2sKxy56RJLt82D/crZ1rziNOfEuDSqiqDwZl5Ry/RzxvLEPa1/Pb2G9dI
0ge3ErLJTeo4vMTV+c7ftddhaqe/C5206f/lAUnn5JAmL+RWNonZ0DrASuVXbCixX+V+e0l+S4rz
6AuepE3LLpAhFc64uOEiTo0PW+Oy3sMz46xUYCG6P+LmGA3MLFwLrseT5yU7rTSRhoKoAlW5VZ6J
u51UBoq6nByahjki1P8Xd3+eKCN+DZ1UmAEBJVx6qqZUqINMRyMqO+m7L8/L4oFNAtkGkyxMt5nW
BhDhhymtyTbL3Pg8QTKfThu+NXoofG81O/GLxZHOGgnihkqzaGhMpwOftqV1Q69K241ahAAaLQfm
xzNFn4LhpSP164u+TyWIi688XjaKxNkNlBkzaj85UHh9XYeBRkWy6sy6pmr/iX8Pe5I9+T1cbu4k
4RVo7t38ogtuG/GkvyueL3HUcOo95C4Vk5g8dziWBpGD2srSqTKC/0MwLnabHq2byBNmmZ1JdVs3
2kQ/JQKvHdAUV+w3J/0Ll4/enHjl7zwpa0lN39UpWoc3skq8hd1AxnEPwWXmZX9nLNCnKVF9jkv4
ZP45XIfTYOj4yHvOiFYQFHtLVfq8WJXQmoiZGJrJk5skmi5mrcWrUth8yH0xOtyuaLFNNn8BziXB
p9j9xF3ybwT0r4kbjHtBkOzpymrFDi1JHEqebPDkFMNq55TTUjXPzoJRvfZyWyETrywcubUWIoV/
O9RNIXthqq/IAe0mGpkD9VnxAx8ECujj5tinf14rtcE8InGLIfB9++p6CC/b29I4d1/h/XcXBg7Q
0jiXPXf/brE7IzqumJLldnGFUrHnJ+0OUyUbeGrlbHsx/v206Z9TcQjkisn1uqiq4f4fiu0fW70I
Nn6sXPa1zr/7a16vsLgFGV7900JGRNJSejwXxb4COBmT6VF8ddhAhc7t1Quc76M8l4CWZPgYlALq
95w8GZphuBSIQVps28JK9oFFbUDHPzE42Ou6Bmc2JvMAXaCEHe/G53SdF0gkJk5+CjjkrdtAW78c
sbZWuqitPZThBaxSZtc/EHNOrSgV/KEPuu91sgNNOmS0ui8H+uy7wK2DseRjHnvVBiiaZHFCzXwT
LyR/BSpE9vIsGuZ5qHZ2B2kl4chB4ante8ecfR/Ld3wbXqgg1hamIsqK2knbIu5PB+iKs4Z43UrM
yh4LHRBj7EkLyW03hAiYeEXgES60nCk60qtPCpBYrD89p/A1HdgA4STVAdxUkXz0GXzJ+MCEKSNz
qm8onrXfxH0yj+uxss4p7StvavEKThifHQpY1fgiYzZqfYlgzqo0kerDGhp9mPJXijyea6vnjNyd
aDkoiLJiVH4BigWLX5dt+zGPa1CUl1ir28hr6fslfzQn5y/TRwCf2bk+Ed3EoimH/giuXddeX5Od
JDP+VCJRZnV77R9TPqri15PBARMHCCTImNZSIuD21TO5eSQ3Mm4P38dzQyPbkZhzt1xsSY+4wnP1
UubjKHyNAB+rBo+PHP2gxZceVSM/fsZJktg1cLtaFjTKb/muuxgsEQkOxhVnm7c4eEbfqyw9rRg4
uWUhXToRN4E3UuEl5tMj5CftMnashJLLW9FeixmZKPOE2wqaAuEyeKw5ac0W2jkqoHsSGgi6bggn
21WGoYVpKlQlQmn9uS7nqJpA8HpTYfdLqVBYXd5PyJjDNcyxls9dEPIJUsUrVu8u1Tw94InArgjb
VV5ruMcvyWl63lSPJuqdpuHQ/CT10/aIeza0yRKLIr8TPCOm/m4fHGIfiGpH7zelKdlDqGzl6hwd
KFyON4b2D8NbU/L7IDPjpXVjeOlWeiZ5yt35g/4aSly6MHwpFNsF9Sivd32Y23Cstln18k1BdAWm
kxz0vwRqhcXf0m8A8l+cfjj2IdClvJk4Ue3dK41+sWJc4iV0OB2g1eaVKGKVwa56Uy/Z4spQYbsR
ZZDVIH0SP5eyaUcm8rJj4pboI0K6Jz0S6YdDiF6gma5z52JIVgsi4D36+O3y4i5e4jIcfhJVBYo5
a9M6xx3bVM9cb1CuwOUP6Kzg6+QxCYcmzaYpyq/YUcQvKj/DVjlHpQ9vJsxppDPkllXcGjQcSErF
amHci2Rf+EjmNuo8TjvBTqkEmyvbtWvQfFPNmYfMm6XIoWnSnLclByu3Z9AxLklzEQhrs1vcWq9r
B2AK3O/HAqAIL6awd0+kHzTr9HNRYq+sv2OvTHr7Zht6OMnOcuncTKKyUurre0bvr7jnhJgHU+5M
aqneOUrEBan29N3WuhCM2oegA/cdBsWxUTjIDaI65z50fE4SegnaSDc5G8EzgThD4F8i1aHd2mND
mXTs8q+CJxwSdc4ib9/AqjUFnxn1LNKSp1gTi9PqTlS0hg93WeZQ0m4gAGiDiF7P/TZucsWY3lxm
kS36cPohJTuoRFzNXqA1ZL876A8e6VfpXXfyVCMiNQlqRaE0li/OQZMGdDtnMlKAa/f9pihEcWut
yvKFhUcCq39f4s33yP2rLGFSzlCCnccwyRowKmgqrEu0pzf/ubMQj2Om0pbrXY+hWEX8n9zABIp9
7lWy9x9Wlssjag45BHUYb66q79fKHaYCtH2gO78gHCv7wbRLudoj8jxc4an2COsJOfl57zP7ClpA
NuYW+V2Z3/0LIfnhuFXOEYfYY8Qcda1Tj4wrhcRbmdHksmrhAv1zUjCycJ9y8f9qO66YUo7XfhPx
rBpXXAK2nGOCo62ELP+lah7ZV52vtERvLh09XHF8phlhxYeNYE+1pQ49t6F7nMldPQXEPFG/yQ8d
FZ+kTFU9egqABxB8ijjfnuKhuxcG4XdpcLZlUQiBjlZ1vs4yfsBzxGuXecbIxsvg8pLyj7egpsTu
z5+TeD6Xx0mp7o3C8wASaMGgGd7Sz/nYgWPLd5WoGbP7IAMGZoNYnR0hisgspLo9Q5Jt/EaA1DmF
enuX/+OFCvT+DlW4Xow+3meoSD+8Xeer3CFitlS24VsPpjP+PEZlkRW7hZtCZOc1LN5noDVzCRo5
vpbRJwkqZ9DmNjqHERKUBr+HiiJJ1T5pJo2Mkhupd9gJgn020LS0bivzOasDtzBu/qvqc5ztQU5x
VX+A+XIi3Pfs5MC1UU9N3xDvX+MrRZQY0b+sdzs0iLeQQHOFRb/KT5A8TZHchXdeoBfAOHRDs0V7
n2zjflwWDZmD10dEK9/QmiKvy96V8oNIZBdRMJJkWz9/lyJ05IToDHcXiKuX9fmWero2KV8G1rG7
4NG2CxviNzCfqqov1hKKqRXh/07wNZZ8em2ZKeIwIZHmXFRnkhubAa96Dl+4r3tvQOjCl6Nlq00a
uB6GUPPf9VstTTtB14DkZFpAwXtIAR9bpzNfa+ZUFfM6UVuifcD1Ra0mwwjNPhsxoEj56Pkyp+if
a7m44DTXIDq3C3txMHjTdByre9lJca6JKgLjKEmYC9B65g5RFFB25Zd3HhfhYQNmENnXggkW9Kgp
689/Ckfw9ioC7906pE2OMH767al3KSI0bOaWNDXH92F4BVfuROZvA2vCvYuAh+/rhmsFDu2H/Fy2
KN+6RCCLG2lDS29XgSBFGlxOm+HfdbaismBbUsUkPGBF5V1KvZmC/FBmKtUAoHsD2WXg/T86vUDW
01nGaRIWyXRBFZGrUUUYhgvaJTnoFbobmnugWvEABfQqd2MWL2QHsjnfqOvNHnn7r84BQ22lxhMe
4b2BUgKgYSuDjBoDcNqby3hnwJIW5mpegIzcqrLYC2DDD549geNE3Uwo0rcN4uncHiU37cPFSjqR
oCxLc/Wwkkb3oq+DiSftL4GgzusGs+UUX0sPT7fGnNvpI87I/8hUjG5/RfE/3rT4jnOKGI+nq8aE
T9YH2RuDl7blttqZpHQoMIVT4Qp+ZwcI57vJfmGBRhcB4imUWzYGLqz+rPOwm9mZM8P6vXvAb09Y
Gbn3wns/XtI+vfnn7IgTOVyO7+x08+BO/m/myO2vpe9A0ilInhgVRxBzzrIDC6GS9xI9uUm+ZBv9
9bhgUh0miRqSpFNz7M5YAqKhD04TkqrLcJCzzqieIFxa6ZCLq0GEl09NAmcVV2/g0pAmoCkYPAXy
gBdFAHW06gwYTMKi/CfH8tjJxMz6e4siFHj0OGKUXW1qEefadby6w+A0jVhdxSEYha23T0/Jr2al
qMM9iqAPLImVGJnS4znuodzBTpN9jJYeB16ip/386cJTrqz/6smcIvC9/jolrGn046XGEgC1Y3uu
YXKoUYOkM0ZVMoY5zB5MSt8Khd3+LDUCsEK8DzJr6sKASr41/sAtYuyGZhjMxQUPx/WIbwOGHjLa
613R50tyETYbDAycMlclnJ1U2f33PJL1RcZ/gZC2VLifdYte6FfXGZz6H6PMzceFuOLQKVC1YP/9
Kdnva0440teETqPDLGQi3uK7RDUHNJStlZu1NUVKWYpCGHUJtTUrl8GTbljswtxg5bKGFh13Y6l+
H045ZrMXVOsgqxOB9KHyh/3iQYBKi0+kADS2y8erTjJrPRTIAADfWGzhMFvZwLt7ynTXUbyPJHuR
6b8CsR8SES3CVf6LwuSRrW47Uzuf55B14jkb6iiC/4Y+1643aRWzRpPyt+mDILHOYkD4U9tkjdXh
eVZkES8Nha8G314cYYotIeTmYaUC7FL5YkE2YnG1a8BIDy0M8X7Ng29Fnj7lHQCUPoDLacs0HDmc
IoADkMYRdNVzh/PoXUhWP4JaW2g4L2f2vAKb0+1ZJCtCY4kmA6TnjIQQKYhufPfB37EQlj3GNZ36
EO4c2avciMGLsF42Aieh5SK/gFU5NFx5P5KvshgFVxMaVMXJCd9ZLDz0bDRRjrQjf2JOVSSj9C1q
qLhuqAOGsASYXrCKOgxPu6vd/YP7Vin07Ru2nGOpUYKWuh+COAVCQEEz8bkojaB+OUJyvaBz3F7m
7eOQz8XMDDhx1/VVj73DBEtw9aK9SfWm8X9CRC0jSc4+OiiNycg2xG0DTjsxVgPajhtMXlz123up
lo+WsWeUn/RjSQP31LVHDjAJ7O5hjA+Iz1Q85+KGv5tFuglCe8eJAVLAKwQIM3OXaZHFY8JA6+ia
oGWrJQAqQUvyskqKeyvQ1hRXwEiINwQY9w0GlHaWuXCegMEmkg6YBbCpCR+HX3ZfXIZsJK55DIGa
NR8qIP+l78sQjhKeOcu5dTWr6C7flotRSIhjcg3D9XPSbwvuXOYHe+kgv3VnIC2DR9sklWjiX6oz
4hfbKTZHmQItVkWqvW2vmHwMo9acTScyveiR77e00SUMIfMl9nn5pnAvYr/2O4HkAkMlmKk48kSA
xvbjzBGPk8U70Fh6elxxgDyDZLc8DyvjdHULVypoNeDCZnKV18eQdleA+qUSosXStZaC2sO1jzTo
pl3Ri1gzObI8XTGINA+nZRiRm+GCUXMhWFhHa6jsOECu51e5MpOWduNiCwiDjZkvPdZC7IpBvks+
6ha+n2tZSMFbhcFoAZz9loJvCeTWZ1k9dyRguAO3BYWrQKpPsPJlW+vKc4lV3T7l62YfR6bLcmRK
fq9Aaw3DVRGffKVOnJoEMrxMVNGuZerB2YX3JZX5g12AekO1PjNna3L2QBc6YkbwBL7FQ32SEN5S
Z+f4sVun/cHb4pFm2PPV2G0Bx4OuL/b7sNv71aY1AoSxJn5FSLDMrD0Ys+WFEFlNjBpF3vzUeYrs
fCGVkGByS3aMNS3u8Tvvd6hpmcSP9yqvsYvQ8Ylgy0C2ATDuIUrzeXh5FNj4qM/bZa8dn6KEM067
GJY+/8tG8OAWqToUxQffDH1riDvNd6mXxVEKc8OU6+/jvkL58dAyCzoojI9i8P5AH0kReGCb1O2H
JK2VtJFppNYGQb9oHVUX5WJZwn6frtg4keT49Jqwlucx9QQa2Uv1OFyFfDqEWvhBsdZ3Duv/0oeM
XkSfilBPrEk//deTBiXorbF/em9G9XC21ksLcZqY8zFX3Asm4Eun0IS3UfTZ81iMRLn7NpB029XS
JxPHBEjHsMRcnUHGfcXclD+07fqZDYA/gJEHALeSZUgWcWC8cnJC00M1op3PGvrOw3pQX8Wx55/l
SIJNJlldUGNNjFkkQqr5fRpJomVGd3azqeUFNvshEmlhF4pxLBBv3olnBM5/i7aqv76q9IfPTRP0
57vDPZCSslY0EwDvfLz4OP3JsKmIdl7+cTgigX3fJI9dU+tDvV4+/84XxcQ9FHolpAblCUwwvnvP
hu3C5zULJgh9sxaQEbeJz7mOT7WqhiUiB84FG5gsBqeWTGlRGnQ8QYum1DRwocWoQnMB97Qe2kKp
FRDw42u5wqxIS9OUpESli/5RZ7w2mFNRXOnO44gGafCy6RYXTGg34TTI4/CjGsBSYsIx2v/fsneG
TBz2ZZrV+z9twvDnXEC3V2uTUKLIb9UIAtVgDj6ReIIQPY+aRIu6OQPq8JjKQVIXsOwBdzcGAgBU
ubL8a+GTBWo6opwSANb8JLjdCoX3iNJbHxt+fVZYRfoM1mCaCnuHHg1WHaEUqly/DCtPyxWi2r0F
CWzozGvu/ZMVJwN9MXsnra16BFywORgqgEHnlTDehugyKyJEMH75/Y8LURv43JjyFJTP5chLPhJa
U39UzizKVD8dWhlMUr09c88yFMI6/+2C6lw2dCukzSy33wclMPlH9fKO+RnDhLjallChuMsFrK+l
xELIA2YIuQ8Zuccq7IuS4hyPwZ4ikVbW0cwRXi56DrXupUbSwk1zvU8vb8Zd4URZ8Np02ZOxuZGB
Pm695LP5riFZx2fVKHq4x0iOHg9WiOgQmqyUQ4NgGOKbKQcFizuxSEnwmOA7FEdgIsu+5pV2qJyD
LGKEsZvxJ3qfbFV7lH66ncWExJXYd4e5+Showj9pVaiIVy+EB7uHiXjdUzS3A7X+HVpc+ygrMzHC
ogY5ACMHzRy7364v2U2PBHncDPulnZuzTurJAyydeEwAeie5JTmDj4q0e7pgJINLjI1ZSJnXkn98
3bt0uqFFMnHP/FiCD4ZV0FbSc9Mlsn+rVgS92dBNYm7oZIp+R2O9zRoe1YL+rL2JaQxUWMVY14S/
06Xc7YBvgzAIu8oHV9Tvpwv58OQkZNSV4s27Bhtvy27hxt9vkLT4i7PzuBk7L6mutpHO2lQpd9lv
tkpqX5FHfqnugSA3pzPHATar8NMesLNTwI4HLSORDyabh8atWJWB+nmjT8sXAeWR5m+ax6OtvzHe
k6fPlApWJRM+EcZt+wZDaCCifMn+SVRcl05x9knifefXrST1P+EnJXs4MUfm5NYXhYHffk2cIRWV
wBH/+2uJiukZbQfiM/LagIL1dqpsAtwhDAxeBNjYcH6HcUoCARcEPLoauhzFVyda4H97B3ds5AhR
OpTk5lwuza7JxrqFyjOKueC4xA1WMUQimXoD8vFVa0dLKvVtMl4Zx1ilG2hYDedVJ1lbxwEsmqgC
Vqk00AHXG5mPgi7lBGU3BsODfjI7j8HErB1R6/GwwfUVcqCMm/JbAIOq2t21VbINSVCD9AbNzYqY
q4TW6bkY8Ev9iFXJ10gkMq6POVs/kzAuYjD8qKTskl++JkVaS/Ne1TZowcFVUGk3B36U9N19Y1k+
T8gw+jf8DrCOq7yGrwRxarHTEW3qSoU8176CILH9hS8IKlUxzys79IKsGzWYyGnbv6VsmvwctYZU
VsCijT5KMANv3wz+h6283tRKKcA3zo+2r292YiVULc4Q0Ladt6jkbMTnaL6Q0JFWgFFFj5Ou2VyM
YvElGlS9lUvAo48OcvXMnlK4PsMZ8WU/WWjjglx2fgIUzjYAyfKNKGxXdKzm+JelzGzYqd1sweCk
cqGnHW93lGJ01PmAo9ieICXqYCe55moiqBeVXxYY9szy/qAGvTVlUmYhys3CXlsSO6aJRkP2fChB
bgG7C/wlDhAhXmaqIu5cBSJ5XN95BjK0Q3HvyjJTOzpN9c5+mKDm2No9sd9dMhXt5oCs652hw0ud
N23rDV2X7sj137MKqfnWPB+Jn0vvI5g1uHu8JaZVOpGvJ0zhyjr26Crd5K3E4ogja9JJQWqFhIaE
ThGo/j8Yrb5PjCfC3Dh9FbRk5Tu/X03io89jaAjFP1TnSViN0AtWnKHh0U41W2yuFwkDHynreKoA
Bk8glhH+whaFD6zC2rsjEp6/nI84gl77nSqtVlGd4K84QjKRmTD++RutFuhDvMGXmBMaOpdN4qSZ
627mGfap1H58jMIautoIPViv/qWtim1iZ11VDh7xTcJeaa7etTyD8oWg6D9CBKo/YuC3s7VzHlmt
9REMKLrjJlsUfAOgmCswDJKmOrqP8bX/bAVekCmq2n4o2ykZ9UKZFzXd4mXAuaNRMVJNgJEyrLC3
1eif3Ljj3kg59Kvs918D2sWDA1FG17zMvkgIGc5cCwuBP9Q6bxKOnx0qsoGwUfA5SiFkI2Pmo+4a
ycMFlQX5f7RxhyaKr97UzJe7ofAdAs6EBoxkiuSuNGm9LyWnM9i9kARFm55GVHYj448Ogr5BEWL2
OjaUphWKcye/1JkY0u66+YhewbA0M9yR/NWWTdFRwAiyS/V7g+E+0WaFKkaU11N9jkrMYfN4VAUg
C0gDc1EJ49Wd3QkXP2Prac19WWbI4C/R62AwhK6MYd1RhyToq+itaftEeTCS162BcaFVgUmKeCTr
A1BAGg4ttZS3OxwwQ+096MRS+QfieaqE0tgACXmQiNl0RsQZ6t86IKL4QUIovEKueCj5B8Vw+i1R
PwWVm6JajG9q60jhJJoXnad9WJ8UoNoTcQyS/OuoQUmi7zmj2+YZ9LABeuA9OZipde58I6gM8tZW
Va/sUqPdElvpL0IWrMQ/P+fVJiBCfj6PnkgqK3e3UzUhD25ebXGRQoXVEwq3G9eAc8CScyALg9Ey
6r5LlbO3DfcLMAnkGLXN2XzbHO+5IZMhfFENf+Osbrb0s7ixGbsWeseOQ88hm7TpxpXXZPNGjCQW
s7HlfM30qb4z8oWWOgCv9qWBOsB9W8bzqnAkTPclm9nDhL8Sfsayno0V4yqR5+l/5UlnBgBByUf7
I032sZCRxe+/tzCPE7VLuXWvfgrslGqYWc5/pMV5FwH4Sj8IPC7QEK9kZrvtq3VmT0mE+Wc1Uz79
v+WpAbKghze6qI99LA69RHtqHq5O3Ze7zTH9APiOUZOnobYwOFUID3DDhbgFtPTlJCD2uqyb4ZLQ
BLY8v2bBDfTw3zcYClzs+4S/nXgTfE/EPGN9CDqin/h+ZtcNtj5esc8YqXrvmAYJAPWj8wZ1aFX2
ckmdO5kLZHtM4ENAXh08D5VRyMfUdPE5O1KsHHTWv1NqsSi5ptN6pg9TOQK3LqMpcHYFgN7Dzs2m
PdIp/1fJ5nShkcuUVa1QgGS5QcmtlkEPBD3OovSCNuu0hBCMYMCbu/9niL+n8Kn4e8JQ4ePxuS/W
3pzlvG8Xg2pH0S1nIZQ+6TrHQwx+0+A5CFWVVMN3bgWpzppDdFCwjF/TTqjWWDgvhuPgHcwnjczK
5z08+/uUY02LDRlJ6DsSPS2bPT0vMQHu9RiwChNdMxBc+/oleGkfF0SNUE5JyqWV/7QN3njWFQPZ
TDCubtGAwyUV7nt16yJnLZlfPQw50J2huBScPcC+aeVul1YfHbxHypdbqvdY7T12peh7l7LrUQVp
IG1Hiwt6zWs3GN5O51tX+VJlvxbXAGKicaeM566852CYj6z6w4GbEHjcSkntsdEX4V6KrjUXdgRz
/nvwPSbDRsFocPKgwEoedkaYGWdxO+3jkYhcap1fGwOY4e2j3nfmhg4wVPZqKCi+8zwq5KL4k7D4
2f9bxHss72fbUHRud43qwOnnpsOx6iefIoSk4Cblwa3YiBPOL7BxVEh/MCuqwpq2FkVIMESDXMOx
fP3qQZOqn4zUKq4bG8ak6BkgsnMrPj6uWhFxQ4DwEipM6leXU2XuQpU1neXgCfZMqfzXUJXOa+ai
iTmRY9PBlY4R4Da4OnKZLFciX0YKAaKtc9xk/PCMxPkBAFtW1QPeynpXiQMlch5zayM8OPttPLM3
/ZxGmMV+W9jJuolmFoOk72do7dZcmTNCeYHhScE+pILgwNihg4XiR9skk3hhmZtsiUutfBmOTUUm
sVvTdbzCvvJhbHyS2X45FZgUR+iBaBE/EGvzDj2M8fAgMR3f2L3LJHLDjm21/8Nnk+uuW2P8qOhl
gSuCVqjAVLwfYUPYiblezsInUPiafaCRv9JvubZHN6QnjN8QvHcoRAtxnvchAEleGRHQ0kgekg1y
4yOq4rn3O/cPsMJmCD3UJsClVVEJbpKKfvlSLEn5sCL1eJGOIa9xvaPpWzYHafmJPdBSjVJOc2tT
8qpSrdAwko3kFfR9U8jRmik1Jb8MH+9Semsan8s7Oii06QjoXqwYo/EOMPcp7veqy8adI2ddTIyX
mqqk0Hs0aAtZoFpwX5dz4N4CD+ZFBBnIUsWpSM2DOzsAiU+dE58ISzkSB6LbHuJKKFUM8uj7iOcU
nWPP08wuYCOtbngkQRby2x2YLljvI2dZ5c46uUAglv47kiCOIOGlw+NxUkkt8N+bIZ5bK1sxjQ7f
uRPddisNjUGHdAmEQNJ5eIvtobvk9E4MsWx8qr6cvL3SL0D+8y9gPqAHLyFx8hLf8AxedOLNtsY9
97wRlVgT7Qvrvj+MJvb79hule/AuVaVD8l+hs6Kf/MKih9oKcAgqqKvzLTcXbt+88hRHQUvT1ipa
shhbaRPOaIKq1d2iBV3ogyIZmOBBfop19Iuo4ungG1j9bj1G3lAHTZUqiRPzdbDhvr9CixHu3rmI
x/fg0IoGM7xTc61GkeQLkJIgitnt30r36L/vxNtISoxZDzHNFaeLtUz9jT5TruPBgZCWuqM8VnR8
marjscGUfwCTrUIA/7e9jKHGIpQiBy8lJkHsZavS8pzRnEUHTg4hG6mxSF6T6aoD9Vj6afmJMGoF
krFCBJQixLbIKU9djpuh/PCJNbfVbPNHhHWlQOxzlAPhMFIdffjFg+gBQbSCr08w6EP9OucZ40+J
S7ZcvR8oGpvISn2NB5rJj5YmwvUOyf+7QxY3kGPhxBeSsFrO1uExfSJkLvzYWV6194/2wWZZhED8
CDxusbWqYroQMWyoS8v7n0MskJFRy6xmt1k9h23yxL4wEOahch1LLfhNJoAZEmAlZH5hS7mUpi00
z7pB1CW0r9jZnJkelkcNu1sTEeeUWhI5d0/tDVLCokrghEWyzasibnha1/Q9qZwuav9yhBmsvVI8
xeqaVlsbmXbUtDxGsIeNYS3VrQ9lNy3XIqqx8Eh8oSbH5CQIMQKxj0n7LHYK9qoWehjPDClxxSkZ
aCfxn6nAoD1dDWyVs3J8f48trhJhA1uLtvd2nIUJal5K8vsaULJ+O7iiEMQ2Aydv6xUPrslrlybq
gnTx1Hf/7LJfssMD2wgK6inROxjSb6J39u24vrz/bllPrNR5S5K+yG1zxZ0lE7NCfOtdTikIMtrg
6bh/Ci6510sq/otpjL50kdnUpKkGN7mpWP3hUjMq1N/iSpvrN26OgBdEGqYgajR5UM2NEXVsNcE7
Uxx7M5V0fiHRzY0Gedfp9w9iZ70qjEQkTgrfFV3cJiuAEEKNml8ULmF07AxZdlJpRGI1ScKg4JT4
oPsW18tokt92JVpA9IBFYQLli6oqznW/6+L6MuLe2bSHN0DuJsP9uXlmMjC32HALjs0aFk7NYa6d
ygam4cyLQpH05ABI/iuyNMcZNkQzQaxcWOgaAFVMKQ4rTkfauYwa9cFex5a0+87jp061tGBxElV3
mJz7F2davySGWKh2cQLTX3OFCa3lgtIY2V3D8p8pg4Fr3zasngaw100u+2n3h1owBqcLGJnqBdJA
QAW75n2YfTGvlMKOV/9UC3ZR0i/BKRk5dUvkqb20NITp3qiejqGmrDMshQ25VXfwxEc0y42T6+TT
1VgCP0CQUAyVrAe+Ml73TwcxENahW4Z2ZnHi5FsbsE3MSuPE4XfnnvMmPPCWILwAg00SQIug4+DA
QlF4cvhMJ2NVFYkEMY5mER7MqXV7iUOV9JP7mMplx6O5MMYuThpjFyIoc2RqRz/oWqHvD3fPb2P9
kLjgANG97kXzpeK+YXSRHUHO3GAas1DyPRYDaFrlbA+qB9npTtS8lf3pJJTa9JEHhSHkKFRfARiQ
tbUQpLaItx7KM8paBVUKQaBtYqTMZcxWmIMfGMHHI3omzfuck8iSwJ9QVby5LrkXZTLtF1xeBTJM
eqhQ0xpqrV8xvhbKeTj9Fnu+gNqepjY1mj+wYgULq6tHB+zJU6BZqnyB5tZYEHqsSvXxeV85Q8kk
ISYGlLznddAi63aHnY57XPJ8/4gN8q0fgPs4pcd5fZbi06MHk0nWSSZkwbSNipevL51tilHOrBd1
ENwgq2cNy9hpuR+k/TOYITuxDqB+jFVsbuJ0BOx3H9lq1U8H8crDAUW/6QfUXOu9X1GDSmEDNwuJ
eVHdxzJ7X9Fb5qQOdwqNHJHkP/fjuUTwMvV50ip1EDgvrrkMFIYipCXR1KfkPWkIh/7W9MDwVQho
Dt4BcKcuY5jrBrEXQViYQQkvYtgx8Mhx8LPlFF1kjOZMs+8ZCF/8Vapk9aXlBkOsUuQ6c5Qh7PgR
zxtyw/G7i4nuCgqjYrQ+MpEE7Dc55odmn9vBrJ/GDWrqJtMCw/nPYhp9aHlt1RUe+34gVVlAxO+Z
e3oJY9mNprq56/dcxfiwZrlnLZi8F0Fvomu2WijrhgTs3q6FFFvZyGUyB446oagVF1mDJ5sIcIjm
icSR749yOrJDzJ3fMU7aUxANLe+hUJtK6h4HQVyxu7zF26DP1uC0wLQHwLfWvg16YA3V/qxDycTt
LuRkLg+Xcn5VqLi/XWPZcyYD/4WkVXr3aV+ANGWq+r8RSr6IaqqW1shMQDCZ+lKtbcN0gorRjAVF
oVjsCMwlOLFdyL/GEvCAFFWvtvND0d484lvAGIQ9VoRHqx6f+u4T2Mu7w4rfWpyaqUQ/6MMt20aZ
5ihaiWUtSKHYR0El/TOrOINIU/UiVsECr3mfGy28vXSfURqzAfPtQ8/cETNi58EBmU56ZG0R4LEI
A1R+WeFKV7/SLfjoVadTBrPtgFs6EWxVmr+Sf8yaKtljfmg9ADx4vRODq0rsnZ+3GjU8HCR6ME3o
9BAySUHiZmanMISN83rAtLioUmkabwpiCjoEhw41dVXdxPC9ss/+RBgziosFG6o1FZrWxiqPgdXC
MHW7beOTRLXAk9FlZOiJhTsyGCnEKKgVbHEUiyV8oggiXQ3H/qeo+eFFc+NCOZNrpRo3x29rM3vz
LTtOVrdIiF0igyGnxd+XYDnge7ZJVGNk80F/fJHXxGe6tO3Srw1P9ssp6FnXa3ff/6CiauFOn9MM
bCLKAYxxbWoNkrljiNCrLtWGR2ONk/urtw6CxmTXyDN2POwvrJATnRVXbL/yhXFs5r1VIORYJj41
MivACtItW1pmSrZq5ydXFQ+dJS8UAP5peJXV0IVLXUTLcU2JP5YJ2fq4oXh7AkE7y9u0dw81wWVQ
wJTcvMfL52th/ocAqyOO74JWNrr+DYYATZsbTnpKaI1BxDuIp+/Z1XS216Zr7fZMsHhNpuPziEOD
mfEjZRj7QDvfNYqaTMYyDN8x6zFFxkkMuvi44E0zkJLlJgpQkqsPcGasIh+a3UL8OVKGnXRUNBEa
wIH9vBNwz7vpVVEkt2iaHQaLIEhFaD0AwPPzjsPLHeh1G/O6PTVbMoB9ELIzBQKb1iM+8AnHsdqs
wuXlCfWwNwaTIngo9J2xbMPXKuevCcCOa3pokSzgYfHmtbcVrGJjgcuFjBuwjBTmhZEJm1yZxmV8
BYSl7OaXnnWgOTxzF3IyaNlDQGz6FFN1ymLSPIb1GpbE71sXCmTOEUKaYsmkm6LoTkizwmyrihXs
PtKkULXld4qDM62rutay1yB0V2EeNsRhCbr8r/KDZi1KqPj9KklVBo4eneOwvirE9FP5gSvmb0Tl
S6XVfmKMVcQNwFxkssw/3PgYVoSn7NgphYRSeM4LCk6WgN8nngwUcvZ1ObtW3BFBlBtVk/RlCzzr
K3+pNfj+/tAD3zXYu+6jJkZcy+gFylTdkbsnws+Vr5AriM7RHY6tH+t+ymj0/lke9s4AvdlZ053+
ozqxwYqHLbNERj3aWHWuxkiC339KVYS03uSspCagx1+lm4alVduRVQfWqv/8T0PAFVwOoXnhAH1a
ANNtwwBptLal7GsP6mxtBSSurJ/ug8Rm1lhP1wxEtHJ+GrkyHFjX50Rrqvvmm4N3KDsXdq6EaKlQ
XT+1+Hn4xZMOQDq6KLq0P/JcxaQl6H37YJJmK8XtkZBhVaItXycZJ9IvPfIVCaoYT+YIwS9UWPEj
RzM+oZoKPrlhkHppKZjlJmKYWHRHIE89+60uNgOBE1VROxTF2Joj+L4FY07zxwAzurbQb+BPxs82
RX8681JQrWfNVQ/FM+b6Yznas0ZTZMtoTbuzrdafe0+ws97oNubBqytEQEvmELe2zx6bfwpE3jx9
kpJ8GEzHn4+p+moEfscnxodG8D9iuCxykcpqE5d2CAEOjJw3iXBDH1rftg+JYMGXeFKVf1GL9/dz
8TMg1vn3lRvWf0HUeUUEXazId2AbMz2R9+j1969RzLr6LvnMLurZM/GGUNGh8H9Usjii1uBwdrq5
PQzi2ufyHANavHasZP2MQvktbE+d79+ndJYeLUd7MVc9QnSLbu1Zw94Gu3VFYp9thIuW2b2k8+Yd
8Ick9HOAJ21aKeYO8NH56h+Sm31WjbHdovP1It8j9LcM3MdPcdOJ0ktTx4rxMwBJvsoUcf2YslpW
h6dHuCkgyYC77TKvASy/nPRBG9uWBImyS4WsSKWy1ntVn5RkIOKgMBZ7JVT3tHr7AbDrW6tOzM8e
IfRC6q37XYOJFGCyXELHcyhXcwKY712bq+fY4nv5yZDLYrc7Jj0rDyB8XFA+nVNPpAAVc9NLtAQo
Zgr+99WV81pfZ3WhV0QDIrvh0fSA1AAsWLCUPK3x1zTwMpNsXTdTYgzOiiqoqAXmRXFZbc9EminO
SWfwfNhS8I0AeYD1spMiJZJnhwEPqHDfG9NL6KgrL8Wc3HObM0Tjje+zihZy6v3WZo53DZD96Tv7
ODzo2J7PWjfe+xk8NQX0AE4iPwX9xlaAw13Iwp7bhXJ7B/iHleP7BXKQCfVTp807ns/n2sB6lSlF
OdCEnt7yAXd7JR/XAmyQ1fDi67gYPtV5pagG9qzc1F/iDaMevbwOnKZDKD90mjBp/bbLLK5k0jUJ
v7CZeWlQk9EWMjhbFCt0v7i5KiGeAVAopjuaF/Fozj+yHg79AEa4u03a2MCcrFwCeqkOP1vccPLF
AHubT/7zZpSr0z04CAwVJMzAtosklc9UAqWpYhs2Tnv1FwOsCp4tmMuVoxFprvUvxJajZKm0IcJc
wrTtRFxNQ0Gv3DKFe5JkoOg46n/mm5j7kIFcvwY7w8lJOlRVHD6mW+idizLRSEr+JVtczdzixrO4
ai0t2Pqt6gELCsj6pRvG94tw4ZKlW8JRPiOI9EU3AqXs3mFvWkDrViXIsKZa17Yn0/pQ+18rjrB2
IcDM4lSES7ipQZIIxPq+Adfn05HmvEEUq9M/NDifVeuIlaoKvkQTog/u5yemwWpfbY5zArsbLKJm
Qr26tA4NRnV4VIz41jMz0WvvSokZ/AiY9BjkGj/UNdPjtwi9FWqLBl7y3m2ChW1xOtTL8T1zGGZC
5KHcoAieTJmDmtKhJw2LoYZfHyvsunYKucskF0zaFCQeE8mmE8Kb1PgWe30nYyKrk18jTZxgBh7Y
nnlWAwmxPFwQMOF+aJu4O26akiKb4lkpHvEG5WvuVs1MLa/d5gGqca5v9G2p5Ha/CeU/PCMvlHIr
GGNGq6uc+VWObX+0/GkKKrcWtGNLs1G3oM2qyYqWoMdhasC9lBTOmOMYoCTr98nD6t3RpYOhIkDB
FPDWzfxyk+jIAf2xS2CjVxj72Yjhs9PzKgIX+ZOOkaP0wOU8b84fTIKHcJiS0QZYdaBiOo7mNMGA
atiO0z8XAzQ66YcEtd6oYqgX4gBrXXExeifvjTodFxpidnnh6kCV3I+cylApOPSsQC3aUZ+ETftg
DFdMENH6Hh5zgo8QXjTeh0Wk4EHOQv4sW+txRRLoWRE4YnBZrDD346BzACx7IVt/Nv0mhwElg5FS
Zycc6boG/OVFx/t19hVypHK3qg1TBpCITiFsH0PBTEzacCGWJdDnVvE1OtUdyVoBSGGp76NGKOIS
5UBiGM94B2bNZzLGYDbu7Kcsqs5Tx65bmrSxS0JTC71crMZTW6HvkDMA8bdiOhXZ+9676CTxTaK8
4MLXrghKvkhoABj6kb88SAcajpRKG6cCAbOU/OuyzjsR7d7fLUqVZil2u38NOAlwvBS8I5IG2S/H
a4JhX0Mm60P9JYcF0pEIbFVuRQv5VaRh20v9Gd6AyAhhtorsLd560QUXmF+Mod6+RSKaZ7QZFScH
p3XmdiYWyU0dVGbDx3sJmZZoSVasE4sRo8nzKh83ob57cpCUROnmiu+XCSo1yV47taTNBiSBqYNz
JzcFXDUpHq5ESP4WMH+9egY9CXXgQmgFbAjBWKaIaQXW3tZxfpg+dp9Vzi+l+stnTg2nfKa56QlN
bIpQzrIklkvwXhxRlAHmXQnNgeQCRdptmu2npRBwyy/oQpqFUxgFAX1ndyax7QvT0kU+IanDnNP4
kvRXH6HLVyPRVxVfJah0dJrcVBqoqdX0IREIvFwlcWxpD8LXArzU/kYrsZhh/hanL0Ni8+MB3nH6
cHoblKv/uufeoxa45qZdYgFKEQB3rG21nslisMIVuI9toN43FLBmxa9mgCO8260XFLXiSNBP53U1
Njdfs+3ykZI3AytnPenPawfZrTXnYb5bVjpCltd8sWy4r/s7JeL2NRru0JOhhcUjD8aso8Y0MPCK
VT6IqWySTQMG6wn/7nmWNITHV8R9/4OV3sTpAiwMcKvxBe5EpYFwlwEreXGZtpaXJLhz16CI3Eev
pOwBQuO3kgySmcg4qnmah5VyDkH1f4c5qZcQPbTSVz7Ibu6x25WoyqG78AgDuHVyjnKd0PF8xd93
lWCkLn7inwCkR9tWOyZ+yLOZpsCUjxYIa9Xmr1a46lLz4VqoUOeJjQC+YEQDuZ8tSL7IsC8i1ZVg
NX5bo2HXz0IWJJx4jszVQJT6S0BwKQjzurokFCo/x0LShSIttU10nnyzo+P5N+yrqLg2wAHPQwfp
VaQiWNac1xSDZGI8Nt1HrlHKjya5Rm2Br6YMiaHYlRTjTbFyfMCSR/w9fXBcJl4oaA1YMuRaiLE/
Fn1ACYMHB5vDipYNozTV+R8Pmp7jzISiYHcTEI7MrW3+49PRnKrsB/ZbTX7Gz0sRSudzpvRAZWGH
KNc5ZA/N6gnx+VMYnYVAuUwKpTWXYBdXT8DUl0RIL6RGBbcwSW+6Cwk7didNct4Dj4+7fjlYFOgW
ch8FTDSp7fj1BQJgUSot+TeD4SLF99QqZUM8dZ0lWDFxKaZLXg4qBz52VKolI72tO3NZ5ueC09tC
PR9rRB6ysmRcOr9rBYdBKmSOIJmIzwHmJ+8cbapMcSjO2SP8ZtO+a+8DTdbGFa/F5viCBGUUOtmC
S/4bCxJJWuqizEGZKy0Sfz6TtQhnBNoXdK84/uTpSU5V5kk6PZ7EybOT4LlljLqqszM9nb4QwoMo
PeH1rG33pSQEvzq6IUG5/cwEMFYqWCZWZDMiAQdhrYCph+dWfijvi9Bwt0ufbMEs537Ik5IxOFZI
CnhEH+nG5e2aSRLEmJ4Q0el9P/mXKIvyDm7aNZyKYKg4lGmusWejjuQgqXOp9Zvrbd52ZOVA9s/8
G3hXn3K42JeXVwOKfttwhzCPZ1bGzVTHn26WoHVzPK4SfyePPOhDBxdnkUJvkin0CUnIUSwcrGIw
zuPXB70TNHlPhwm/4G5ikgFoRF+NQPsEKSp3/Oxy1j1MtWFxd/UW7SwhR/qK44pPAStRs6XDpQy3
sAC/3U3M6ZkvDYg9deAlkaBpEuwr2BgnVcrwPZlMdr4SkElWOWQCmSmhqul/+o24k1GU5hJE2pe+
PP4b9qEzf/BPLcEanyKXKcfMsXowxlgkkUssJqUZTBkNbqFS3AE5YPGaGAyTwdV9+gJiNvK3be3Z
MVgzc+r+a4lZI5bwFRh5n6b1qC1qDAQ4PtuWzoxhL8kvpZAfjyFOf0StFcMD5unzAiG5uP3oYCb/
doYx/sJIbWURLmQjpmbzlK1I/YRtr7ryfR/kA7SplWiebw281XLAk4GirNvWEGr085Nts6lGl6L1
1NUd22JZgvf98fGq+FbM0zh8mYyVwt5Wm6JeS45g9XTg3mYCOln8Rq6rmxk3ftfTx0/jh4biN9MF
gAs/7biIGmCHBzd8FqncwhAklr2pAbRd0pSekXb3XyHTqe6sDbOFPtqrf2Z9CmmECSomamf2p+H1
SVC2RyXmoDczqUi5IF79puFxrXyGDE2G7t7D/hMBpYj9qZJ+yoLSIbqJfcwuqOPiDnhLbiUFAw85
FggemPziInXwYCB7w4NaR4z0mUjiEXuAEVbJ+Reb5zNFBHUuqOvQbv9DBneAx2OcpxL3eSdKDRV2
k1yRMzxmeDbyOmRgOe/ddF1pknvFBqTh2y/2pABf7QDAb/DqLB1TRVWlhEnKvkl99ixX4nsMq/ie
z2aQKE0hQlBu8JQOYOhM+SEEngAwZ5rJCWMsCl2JCp+IdFOYZhLeBSaLgvWPevR3Tcig+JmjNQJd
/dRt4+Q1yoglSz69jLa+ouTPP4NY8cEuqxsw3+/T793edlffojDJO6rtNi7UxFMZEizv5NBrdClU
hXjO6pggrptcX115BYftvEa9bkqL5jOJPMuwUYzIaoy0mQyYkHmYrKtLfZ3XjqZNDg29rM5Ecre0
zK1U/buIoj9kZlYCfdPY0tbn2S5DYaHybgkYQDHrA9dP/EQ8GbeYrlkTD7+AhuLI8UfwukVbevrn
2vFkzOJ4JN3kO9fkiMwEgVkXo5uOZt+wTKg/fEO5pOLB6z49TGe3KjXC1f4Ji5KsXHw5Ofm7TRkp
TYUiBvMgqnu4//lROcgztFC9hZNv3tLZC6EE7JUj+oKscxFKHQ8XA6cQVqy8fFLO3W7xGJ+ZuxGQ
VLCC3pdfbo3pMPvN+INUVYgeQg8TAjw1Cb8MjxhNqIoE4Erwhxb5jPrMfR9uScuFZuIbejcdoh3h
qpu7vBOIM0dr0ks9QyT/Daw10vK0ZWIE5bhVd5X0D3uxkCAkmyfdQ4LV/+9mi68w7sdd2z6iqd3i
XcHOLB+CP3PQDk89ADw597Vr4XR5LLQDgrJ/pmWmG/nvp2dWF3uIEJ4lMWuRSNkw6GVDXF6mxDRM
E15civ9g5VRhk9GBuRv0YUi9Fh/Ygppfz8u4Oge03KSe7qy0uRORaXbxlrxOn0cS4F8kWb9z+qt5
0YbnggghGA+yGLBjBDOFYnTS+EpO4/8FW28F6DDBVYRAAqZkYjGO1ybDUS9zzsClfqnqDpFhp7WO
EqpOHXfRFm9+sfjLjK0QAx04F10APYr/KGi8eqTC3pmcGwD8Zj8DjNZa7EFagfx84hunIXYxWJEJ
qpHsQmoowNx8cjnO2m0O5C8sZ/5nvUw6pQxXlDIungKIcYTDRd1yL1bNXqZEutxbZd22LdtC0seM
6V4yFswWjV7WXYFyWoZ0SUfCOHsCxOLzpvQBpSOK0SRn+V+8L9wGFK+sFvSxk+IZf9Iprz4twiqv
7sasD+q3Q1r9eaffax01L7FS9IumrqjomWXKNyU2n1mMaEozlE4MBo6nsmBIeQ+y6BTpt8xgAZNw
J+AT9yRArQK0R80rL2YH+5v+9zW6tzEi6AmyqTK3g3idDwn+/SnG9sxmMKb8Sp6Wzpf/vZ/pYC1N
7gkVYWKuI78a0LxamaYZMCaJ+X+rPUvMcsTR5vO6xXoymOSnpRMjCJZiO5rg0OaaezkdJHUKZnzM
Q98fMG93I0FJgrhPS6J1VLCFL+tv5Vr8ENeNcQgHVAZtirRBGL/kvADWSyYCsWYraOFhNe9uU6HQ
pWuU0TLjUshFRnGgySsJ8+EHXvqOE+QLx4fg5uKXzCXxPv29w+oEkY6fVW30QVbGjVFpHivg1iCK
tYAy7mGemheBB8ioGwFVOx5N2LjJ1soju6TxNPlkP0F4OLqCrNwGA0qF/8hGZPCahNVRGt6i3PrF
xQNAbBdRCSIzhMWmt1R2ejiHKlGUHUk9gOpR1/Pib39tTSMGX0nA9zSJq2HLPa5Nv24PFfnF00vI
6ZtpFead6tbRk9lLSyD6djmy2UxeTNydixvOv1PQ2Do99O+5QCTPmN/UADS1MMoiVnL4EN5hvgxT
fV+32mRy2b8R+gu7Mv2OPqJmKhThKbkcF+njTk+1/sAuZgjSd6mdufAfSbd7EHBgoMsoW4hFUQ1E
V1Pb/iJYCGl7iPg1hit5meqv/7vbmslT3i+hiyAwsVMC0TBB8wMRn9hcv3sg6AG9DwelT23cr2ug
nSwfxqIez8GJhimgJq0iFO+Lk7xert2IVsbX8m0gw8Tdrj4MhUbQ1Kb3T/XJFLNduSV1EZ10JpqR
z3zk7CyneHm//Ri9lpmU7J7lFxuZnYb7pUYv5pwXIjRwrDnadNE0BWwhs9kkSA9jWC3QHrsY1FxE
5odA0wLn+MOqTemQEQQMbss9gCP/f4OznpiR8XXijJ0G47VhdwZyYfe7yiCwMU649JPh8MhjvL6a
yL5cIgR0Aayx0QimYg+okZd4oEoWWT0I7WhMKcJk2JgxxK/CYm0bZhr3DqMZkKyLyhS7gEwS7pbM
Li+of/ETBJ7X2fApQj7bXTXFwYeusXJN2PACIyxYb6nCL9vv4zzDTO3/N/tmXt9vKYxtU8FW+FiC
Zag1ZMlo2sgAcJST8Bo30r8nYlA3N0XFb1B4hTQ7OzGbZJ20YOZ8F6cnuf8o/CT9EqqedFninRog
LQrFYy50mXZRuHCU8iuOpyQMLF7kozBPpZYQLd4Udg6+6ERQ3VmXBylzygNx5FsYrpfzH7k8JZDq
r8xN0+EvXXD/Lk6S3x4/+OgvPLhIq7jBTUai/g9irvn905g21BQqho6xSUeCRf66utpxjb+BXDUL
+dJ1Wi/Q0gYpWbYW1qOudfCuupNW8g5eYRDMQs0ldN7HCzqHK/qYdaqChlPIS93IktknE9zXBm3y
JhXnM2fu6bhVSDHVxL5Bc4eykmJ0NbUmkGZDi8U4O3f8uvUJ/ND6DKBhWBWRIcqaOMhoIkFMDw60
K7YxooIeQf6aH4OiZf9SUD+XkuEv7mLfoQtbXIB5HqCyt8GSKTMw+muCOJ3rv4e5NCbBcv/yCC9K
pLuWhxEbNGAgPC0bnpo92GRtOIsXQ5TbHa1Q+MH7Y/cOVve0Yj1EhhdYApUI13qjM1epH++Xoypf
RMKuS6s6Zwj/BRrXwjCfOKkWYjf7U1/g9h4My4n3g8WmUX4drl1Ii0A6yofPw7GN/4Y+q4HLeNSW
z6ljr+SM23qkF1P3c/e5qEwDC6b1tvZDYcKJDQZYeZKiLJBgV3jOduNoMpdHTcKBXFRF4A6TIoXC
0WR6UxPtYO/+u2HzF4hkusTzziq/3eg5AZyRImGSYyWLfePOp2ax087Jl++skUeId0znaX0wtWTu
sKJgQSStBtGdb7cEdQ/zDB3MuSzvc2e3xDWK/VAJkSkq/6Qtm8z66fnhcyd1/+kRozuCo523plyt
DY49bIQcWwiEsNfc8/vFz6LVPyrROss3h6x/yvDl4ofFAq9Rlk5jNuawlRuhrPEeryA56GKgZkSk
MBhCsmrJ2IrRJLEpFFt28GzTMTb7m2QSojZJmS7XUUmge+/cIC45F7dxS6TGyFpjyYCS2KK/TUPv
gWpDVdfmN8b3dgBa3yjEeexZiYDYN+/oHagOO4zqc2lG/NFzBQFEydJqSM8cFAhcrn7EgEOekt8F
LzPSpdkTS59ZD7kffTMHUNExTxkfSjagDwnSNgeFhUgwyutXVZ6+25XGdZ86iVTc6SOBzvHB1DK/
3zd6OMZW1vqslXihkKuQdESaQ8U0zvPEgxPdEJ8jbDcnytFIsoNzTxYvihsKfU4rEULloyc9FSEd
NaVZbrsnlbS+PCs1JUF+AnCmC3QU0I+8GpPigdTMASjSsX6D5N/tjddzMRh6mWo4SHX+Ony5pXcs
63G/O+ClOjcQ6B3KtX9jjBD0fWvzGRVlIoza9UJQvT4BqNEPWo1AJ4zSIiFztjrZShiivoK3mQ3k
5b4BAmEv2oFvGNVJApgk10J9Jk8E/ZZGu/do3RmuUWoqtRziHPl2KXwVqZrp7ai4zOwJFMazMAWS
I3YdNEq9uGdDnfVxCQoyldhMNvKqwICY8jbkkQq9MmsNhVn/+zmJHxOBcztQPqFblzYtCnaYN+d+
2fuAULx7S9obUCIvSFVFF59nwQ/KXSKazZ7ichXz5yRstJCW6d2naJq6mkDHD9ly+dYLBa2xo0mZ
VXxAbzVzj0nYTnaCl3WFXx6DFxrwx3Bci2z9L/LsWmy/pHE2nMgnwz6QFMME+y23rkK0fnbpFvpk
YNaD/NEQg70FPpHrBMgnzYDgPi40P+p34+Ck8uND3Dlz66QrPaGLuiBMeZl9RZ2ZO/k7EWPaqb6T
h7qZHwUS9oluUYYbPYFq1dneK5c2TpiOyDIB/0adSlw0YU5+l47GsKZROaYcPXFD3svwakH1RGic
21MP/mXHuUU27WigRAPpowJFQZg8rmr5YT75mfw7gG54lgVO9uAvd2G2ewby7KjAABmKJGarQvk3
aoV4rcnJB3K+Gk6jAUhqdhnqNJDLFZFl0pNTcmT4EqFVS+xBB7WTt1gBgP4s4IMSrB/Vg+CAwPvQ
dvNHihgsE4zaQ22+TdkGoNWrJ0C90GAL59K0GnV+NpgxxdceSXHNVUM2Phl+RtRqbwlLnUlf8eGw
J+kNnCMSGR1BTyVoX8DYMTnBVrlOvZJzlCFwvzhqIY43v+08p/JlK3/QU+NkBtr94k6DKt0ewTSm
/l7L6Jty59RZVcRTEw5HpJXHKqES6BaazbNdgrC4hVM5IR52/6+yGzcunjDymFWTA/uVc8wJo6F6
9J1sKw+Tf2V88aTA4lG5ZBNQ4RIsXvsHl3i4hf8JILpi8aI4d8i+VSYdI3YSJtOXKM04oRkFIaAc
vDCpcsTFubTjfMBaMyvmJEk/dt0gt1aF7O1qr1muX7PO9lw7DxdRnkXUjWshuZBvTVOTkPc9sQF9
phJSY2pijxX0qP1uzSxzjvsprmpvUeo3PKPEr4PzhTWumggJR5Md57kR0dBruCZHF/oqzQk7EjNO
qdmlNUwvxAu+ZYe2OMDokq8bvRnTz6RqbQ/m3NqdV7q3V5tR/vhSaASPEs01NK3tN3OvzmfbkWIR
MmOEkUZUYW2/D+Ov5uxCVgXZN7TToX0k1h0wA93P82tdhgsEhUJOwIXX/X0qGg8fmbMkqyoYbPf9
SXQchP5B4Xhc/+TjmavYCVvCsM+quIPxfKr8FcikaVJXiiEJaWNRh46tpWlsK5PkhV4whNeOtyRw
DdTOrVqpbV54/Xjs/ADkeGi1RuBvJthxPKSR+JQraEwoen3FLpeOZOpHsohVBLcjdNSGtv189mDE
RAfrEEHiYMvkWgPkd/IM82Qk33PoIrgRbIjB3ePosIzsrXkJxHsOCrIm4PTPUHE2idO7HksowmOi
reXJaMcmh3Xca+HVW+BruXvZduWLaYeFzCJdsfG3xDArehqdlLdb5QsVod9t7+lg9RkzP2nGa/lD
UHnVe4NgEh3tMphk9rNJOWmV+sf5gFLEEPvmkZ9saJkBWy53odW2VKVS56kPiP+uAWj9VyYkeJEn
R4Dd38DNRB3LI8hqUVyWihgM5tNfNjlcFOFgfYYY5tQuqKEa87uCwC/i4XQRFZ4tUpenmFH/Sc8e
MtOZccb43quE2WZDw5n9Onc11J8vDH/jKwZfIuOx4oXF1rZjOnIX/gMpveOGPgJ4iT90Uj9gg2nU
timYvdqhIjl1iUQBVORgGeFGetI1TQJTu97QQyeYH4gxSc0x8TE4w5o0/fwfkFhEKIRNnR/lEg12
3XcBs1INNawlzqTmN/Q3SDDbZP7xHU2IuCwjPE3HaM9g7X3Pf5WvmLFqOJi2ZYot2SnV2x2V2M4U
pamPduGlp5ocQXXNjl30aI/zRWBpQeFLY+dnuo1uujo+yHh5jhoctqQcMN293ZpIt1lXQaX/PnYS
yfGDdFvB/yoEFSjdTzdDVHWjX4YrVtE9tx/HcvG8dn8ZCIRA8ZWK4XetPlO9KAvs2XWuTGzRzqDg
HhaHOPMI4zlUZtC84iF2mSE8t79ngNsSPt9YrRSE87VkZsXk8N1BjcSqWPPqKyRCHJEdTDgVfLkg
rVXHHS1M13y96jrwRQNkNjhHDOFmxQyk6CWvLZiowZ7I1x1Lln+L1/uJYTdJ/2UNkUXb1lIteVbi
qUlcJgBkrHOcqn3L20zCqhU7eGwAFIXtVUmk0xHZCis/oL4BvJccmH09zxckv6HklE4YN/sWHHtN
Z5CCnuaLA04k8Sg34XBZ2Gsrae3CmvTqzGVTnUCw6zKum1nammUYwZ4d3Z16OkpKf8OHr2pZsenW
tHKs1Qbv7o5SwCuJc46kU5KQCyz4O04ma3b/+f+/4JqLqwa2kpzCwO/lYnF3UO3YOyoE866DovV5
56/jp7wcc1dk96QLCOUAMD5bajHlS8E/blfYyJLHDah8j7rDJKfMKA4DB7yz3hvrxF69QEN0cfTG
iYndG1WePwCE24jUiZh9Y1SSAcfSETCvZPx2jIzH4IJEoVfYdAAcdsR+rEQlWqWaaGul6AI6WBwN
UbrN664xEgAKyKknqWWhYKxDTGRY6jfWkhHEDj9oEYp0T/Z2OIDpvoXCLuRjWL4sB9saIcUWuT1p
tJ3zfd2buakruTFy6gJN42XY2h9zmRAmD/9HrG212YpiEFOpHt2uZUCMWT2xx3rPdH5DeBsz509R
vlpJHmy0BfAQLjfsY6wj2fKqwO6yQKW7lSnrtJtLcBGk2N6+pgxz4WYwcerEPqk2gdRRHj56N9c3
xcHWiQJuEcPiDT1GB1xqYTuABQT19HGeGSHtgS1YnSWxqplQ9+VtcZMGk0ViWm+QFauX03bha1an
6BWAYMAjYIfo57S0xmcS1lhD0v3ckKIz2r7qzpwbYIuw7PERd3qU9UsJqPEp5/NyTMTrk2J6e0kd
MVh8COuGBbbFcxcBrJxxv4+8gh96K4J+PcXxM9DQy6M0EHo3IRAgpLxMK8/k7gC4ZScOVHN6KZ5i
RpHp6IfG0oGTbKJoqCGBaq1Nw2ADrwq2o9bmjqfKuk9aBa02csl+53QlowIOIWjnd5f4nxJPGxTs
V0DLCSQw5OgxAkWvo4ohJWLywWjxhjDzkQQEkIB85RyyJN3KS3uZc++tJ9cE4IaAR3fmsee90VO9
B79tOV4O7ZhgTUIlmZvAuA4DwzM2LEgOQWj6CPy00dk2Ba4JbHh3nX3Fbcd8AzyL5c1Pm3DDQBqX
bLctHgjVC9hcLPi7bKoO6FAWu2210JQChhHhOqHLAwjtL0LBKgi0uSQHlQ3HMKqBXH1CK4Oou8QF
htE349XfWSqGpMI5zCqkZzZKH3M3hVatprdSZJtyNL3yWCpehALfeyWFIsDorHpAFdRMJ0lA2CY2
95kNMWHh+vNPgagU1JPl0YtTHeUP/i/YK9VTnmhSFgDyzmGoOIDlu0n1wrinjUXkJ3HL5sNJq5S/
ct8sJ8DVJ8fu1Ut/YkuGtdYlOWeJ0O7ApqWWLEMDi4sGOax9DUDckEAVSA8TnRqoADnUCB1p0w6U
oBzjeiFGlTH7t/ShWr/CTrJsPlp/I1yR1MAIafPSQqwIz64BAE7QWceG1Sg+OYTBPPgb6S26U64I
zeYzZgND4zQJ0tU/+rnGP4wZh6RbRPdR7aURqovLrqQSLtl/67YUUBQFWC3ZKVF8Y7OySHyTrE/A
HD785nADcEj40Q7TXiq99JzqK+x0QnMcvLzn2Fw10WN5QTg81Kz7pSJCIA/u2dnVXfnOcT/rGSLm
t+quV44+qQvh+1rOjMOwcVOx2uCDtAqHL0LYLx1AoQYe+iKLOGYGnXiDLeFB66x5ySEiCqU8ngQy
eMTtP5OD9YvuFv+NI07qhxxyq/Wj60K3BZBE4LrcehQd/V83nYWtVNTxKlr3OYW8Q3zsAlWmGRyT
PxEfo2zRvspFpqPotmehVTbl5yjuRc6JXYGocmUSvMLgL3agMBTKUsxRNfmYK73uAj0PzhDwXD8T
3kdUXL1tVJ97Y6+ZN0JcuH9lBy+RZRLs7mXZ2P8ThPFfRgYC3A0/dpzasenDC4Wlu0DDVAIVtEfH
vNWLwK0XFz7zeKShrMARnrZetXlRzITtxuEsGYCYVZ/5QkG3znGAdpmqyPBevOBBucirtaR4CJYC
4Qgq5gnK9NFeEHeG2WwEFFd4+ZsP2mSCgXr+pRnrUZfStc7CGAI3U020fLF9Vau9pYCbjLr1UAKR
E4maKAf1PJRn2Ghs8D0kX0mktegbOrwAyDx6W0I9pkqoeHqFdFA52Eo4MJnEgiVNZK8iWTZfxB/H
XlTRzY2xRnJThHS1hE4YT5qjuxQHfxptWSxSQR4apuluaufRnzqg1nQtdMOtXWjJCuKw+rtMErzS
96Me03PuyXtIlQCwht2cRExj8qJ1sDSLRU9iF7jntGKREZ5w7kmg88Rr60Qr/SYww/nt+MKtZ4M9
NSn0M3Dsp8q1PIUVwDV14zc3D7q+sgqNBTFbQJjlNAfdDWdfhqKA/E74EcfjATsAkZ+REJZQa8qw
3a2ZO5CI6U2g0vxe0bdKBZTDcg5SWEMtjtFoQDQt471z4siAuo/MMbd/+0eQUuO0aNIJzfIpVDYD
8upNTv6A3SS+tSMsEotTG36dPdQ4kLdcN/CSDSByu15mcCVdJ7VXSfNKEiPhxRTVU6ZT1nf+lfxs
g2Q1WaQUoklkw4HpSJnmiPJ8LML0B0Y1rtwtuiRW/qYdy8E8trML6YfIAoMO4EuiVv+1ZkLcBDak
3RQ1dZgkPLziLGTtn2yF1LdXtg1UFgX6gp9isbD8tABhnJ5z5KzNTdKSZBy9+F89EmpBs7RMUsdT
h+BHLHCbQXxoDljQgqT7iWQE2yVgXVHlNO6+m63scOyQb3/D2/gLJ8gqtOYkGF9e1spSV9hYi63V
6Z7yO2alCuX2qokwZapDOuqEllFZ6edt2AAmao9lFLp9NM56mWAOpijJHPSLeQbYJQcOqrI9k/RS
lnmngbVq4g1c9lThrA2wu2qXk7tF1puYd6mFLhR+pEpJS0RX2jvyrudU/iGjHiwPoHH1zTStC6YJ
7ToFJsRWI03QtyINV/PRhpKlZyqXi/VEZ19f6o3bOae8xE6PSGBDE0pl5fR5APZW1veczgxPPdt6
xgiuZO1KqLyE5ZDYW15GEBNl454HjQTW2eAj8oZzdGyfKSWKHu1AKxpCm5nOJkSud7xiClY0kXRn
kP/qE2ob8aWzQIYTw0lgHbMf3bVweQ62O5od1lGy+HvKW7Bx4EAK62AouyMRtmiv+Lv0mAkjHlrM
zL/25CHBMNPGGQA0ubyMwJxN+7eH830KBytN4gnY2m5YmbXgdxAqA/5RxD38jteNYq5Fqzi0omqS
K3ztnMMkio8hmoTFVSIyf8XUCZrBVD9wxREwxlfLlh3uYpm5pKDe0oppAJ34x1IkP0vxCdYergqi
5TxkjnRl+jC7uxrKr1atcAhUAj89yv1za+oe0zM72+4K9oxqLZNmL6CYqKklIpa0wORrf3+0UW4b
tYOqk1LD/7V5yWwhxu0WepMob5D5uB35x6X17p/g8uA/hbL8fnl6clMVX1R+xuLuL0I6AzrVzAT7
AFoJm0DmARyCBGC/phvyVJjytR8hxEmhp7FowattCNi9Hc8c6DODYbmuRrZzmDTAXZFPC0Qddc/Y
I8D5Aa/hagk6iukJAw3RCFheGeYUUVWGHGl0nho7L3WwLiunvUXxl1jlO+mHGQ8D++hzM1nb0nKM
Mai3vh3th/eySOJyIVcnQLmHxgFq8+dLLeh605iyK0Z1mLO8jA45qyzT/3MPTEJMsovLh0cmzI+E
aIuhM9FEjQkJKiDQuGb0toSKA81OxbZHhR7i3E9nPaLroQj8xnncvbKq/6LXp8q7/sEu8Ugf+M6l
Rl/SaXfDO50QTL2g0AplMCulrgaL/2QRl0oIvVi/n/9XtxYV3MysoUetqV6oMDlpxtdj9hdKDhVO
p4M/RVG/kCTLieGpksjNp/ooQznuXBSMvmb2IwHrE3EMuF/x5EF5GdDy0I81kLgbUVlLdcVLrJR2
+Juvrvna45tMhsg+4jfl0hZXlzspEDeMe/1l/kuEBkDbR6JLK4NS2K6NLUfp97UnjMtLt0mDf3b2
rTNxzAaYs0o1PM1SkjTACpHUAkmbcZlyc5KAHryNiJevh1ccXxWmfA7kHXXBVT8hh3Kft0yLvLmt
2DJaDv1H8BlMMOllPZLfPEFtIpitWZuKIAcJVffMX0cHyMlNLI1hEna8JsMpCOOxnf1b4b5jHX6w
kgSvoQLq2rnbmuTC5Zw6DFyepa91VZ2Zi9V5i6UpzWXCcB68lrpAj+rO15VL2se9sKMmovBz8e6w
41df3d/KzolmWVhu9rcC6CLDIW9xwHgbJYgnS9DGQI4pFLVWBaQuCahNw2/3X7O7ym7ynGIn9jST
L5A4mYzb4NoQDdl/BkYMqLEtnBqCTuHcqiPbzB8Ii7I2rFGeBTKM8Bha/IJRCf1w7Yev2aNZ6wDC
KTRZvYle437lWIlB0P4scorZqh8khu+RmkpqPgO5dm97+PezGpdjw5AE7oE9ur3pkqkTQK0WpxHp
+cH5QWEiqRTTRWDGVG4QcKaqPzjOsNF4oEkQ/IxNTXePmqXAe72PjxKfuosfusCScAvTFdKhrKsN
22EQJJv+hEodLQDsJxd0y1i0GAjjDIG5zR3U8BGVXfq32WEnZ8l7mZPudf0Rw8/KLmhHdxcG5OBg
Pfw7PAuRNWAd1d5SZ2eaPo46F6sCEPpLwH1JB3nRPsPQyP19c+MW0C4jTN4=
`protect end_protected
