`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ZwRKrWU8XlvThQqU9nAmKQFh0CAC9c5aufWXAU+6SDddUAhVZlPUIkFas1ts016EelrbE26b1d9x
vwFbCW29LtudUsY9Mx/VakjjzkqZFVSzjJ8PAWPQJFrUyXrKUrqEv7cYGZb65SJOz2GF0tXFcfSt
YV5DLkJ8gOPMrk+n5Qdtm0czKYH/4+XsAt1tO2s7JfkB0xivV9COl+oAT3fEF+NBtXqrL6COWwyn
0mPndDf7kPQXoTSOYYqoUjeslbOuev1bRhGyCcMUhVfVgkujA0dS6/mRSZjtq4J31g9/GPd2NHgU
Ir/E8m+Na9/c9xz2+KaaeIJ+upOKzYMmZ2cwUw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="huodO/8HfstlrhQExrR8cpBPRuqqXi4HdSW5ukAarHk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14720)
`protect data_block
bPpwAgCOjgsXnQXQaqdv6eGhEuxwMMqpIq2YcKZVf8ZPVM8PF0JFfJxX4ZXv7Ce31OZsQjxkUlBl
N1dYumlQd5WOgnCo/ViZIwJSfw61DPZAkm+cy4G5S9IJQeGRj64djyoG1P0BqrD/nIfSYOc9vwaw
si3w3neC+etLARY9oeSiXFNjX7jFGQeZumA8c9Z5gD3H3z+2rVFX0Xidb5owMANLM/p31VzAN7Cm
Lz+rs91hZf3/RghnBVghjUEWwc5qsLEfpekIQZu2PfhcgLysxzMp8a3tkzGOlM37dThYi1wzN3vA
TUtiKTUoWk6WcvtQrKC1kh3uuPnBm5SuXMKCr86pQ5tmzi0fuleol/qBKNGBxdh4fW8HgWyXJceD
9ROexkfIjVchJoZA1u/vELFt7SinHFawVgeX4Voes62wrnQlM6yol8qhIjZsnSMxuPbZB/GkByFH
NkQeYDDePzFZf1OjcYWQdwSU/zhhHmIIvP4G78qU3tkS8aHw8JWoPsasbK+1o4WXd0w3y7DwBSoc
H9dGsivjpu9cth5NvGNBOYJm9doHLMw93hPLchEywxC1rlkzYGdEFAHumQFNSq4HZe1soDwKfatr
2UEcPQSQKBU1P16tA4BaKAuXljLGFp0kslM9dqx6TVTBn4oD+6kvqY+GhAcLHMTmNsR2YC4G7Kxx
g3RZ9cbkdBzI3WWEgR15PWSKieDs3v0nrHG/PQLbFFvP/rBxZH94uunZrMZSlDwnCJMKJ+ymx4TL
mBtDwIC/WSO49vArESkxtM+oVxCKBpLsHiPSo5ZjVrNoYoC7kBSIBdsGCZ231KkJaSRvzP81rvds
utfF4cobsWvlBQPfXXtuu+17nKgf3BIFxTNKCiDeBspmXR59InxuCGd0XfrSMY8KUiFkU0LUv/v9
sR6YYwPBWtK/jT32dV1Ylv7hX8ogVEUt/Kx6OHSbaxfAMSOB9tIXwljPfa6M9FzmN4/AiFAQx79D
BI0OPR12mzru65ENnhfHmX+GI+jMdzv3fUpMb3I5jVvflLJVSq85Eg/4x8qOq4xNoSVhPfpzqBMq
uN9fz/7zvIAM8ILFw/GbJ5rkFuuUBmFtI73x2TBrfRpwdj5+pJ8GHHuFMdRxOSi5PN+Yrmz/jkLp
jB7Paih126mAo23BF/SrsS3QaPuj/yoGwIrCJeEt7b+AFYIje5aio2uVUsUxWYBd1VrV4bEfgCFd
B/ZvRgcsMr/Wacw52R2BPnDUMr0kwNfs4z9XZCB6Gw/Z63yDyXMIEG6mnFuoQu9Ttaw/lguIx+sM
n4tYdzA0m+/0cem4mF0KbhfvLnTv87bYXgdgvwpUDdJnUQzRfrC3zYaQ95PdT27wXrnIxuRpKOW6
tOMeqg3PX/6bpdV+c1VcoCUmWo7x7HhZO3e6P4jO1vd8Peh4atNHGJ83Tt2AGjjpNtkclXMSm4Hj
SJRFcLX1k4qchHS/CWguUcEuF3/vvueqeXWdvDmlw4DGq9IGYBNNSio7IY15/h12ZTjgXUGkFM0j
PkNjRN7ESeEyreUfpaxku2GonFiUBNLev5KgEw1zEmKYnUSrnEwy+bg7BNDTj3O+ah8KjONtGSQr
Kt4IQYgxurjbdive2SE9Tq1jMThDYvr/SjNH8nXlgeGsck7TxlPedl2PAvQ6FxmLw/4pkQI1oSig
yU4X19GNvzB8ijfQlHI/11usL8QZE5OOndxLZLk3kRqzp4Z52qp2AqivUGn8pDASGkdgfYmaQhXf
+Ddb8grXC65iVhwVKMxyIZQafzZItJ5DiZVyJ6xAk0kuOQO4RPTOdzmYB6xDAnUQiHCHmGDtT/Eo
tgz7SfTHUj1X+XyBufGu5sjpLOY5PIuvO6XxsqA87cz53v9iyGUm06U4KlPYoRYNuxNDouv+pJDq
bIg87RMvXljSxQind+Ggl3CkY0pYILx/2oUlvPs1pOChocy+ggkJHWrtNaDTV8346mc6T/p4ZicE
geETkESUvWvbs21aKz539cbKuOqVmcxYKofer6he6nUR69rICFtjL4reKgdEeD28Gh7HN66UORHz
Z16KPQt4FRUuUVTpCaK4LJZtQh9kDwyA0G7TaItfJfZTw4wGb4KcdnZ6OSF6JYI9fk0x7PRMhtg2
rV68zYdYBrtYMXJDlHc8PmFPUjrJJRD/8ZrIVettSGK9KhanvXJbn74DB439mOA0cTx8Io+hb1ch
xIDm4/CQZn1jo4afiNcdVuJ7ekwM8838i8XTjdC9Rbqu5FILLmmV82uNiuJQuNMqz/TTjfs4w/xQ
STruEZHRhqppX90tr4EswhcnLwWtDyah+hHZRlKtOdLiTeU35hWjhyhD/eN2NHEU/yiMwbbZ10hw
pec3Njp4v71vQiaO9iXbA9JAc1zxD83CFxeND7FmVgiMqY+6ohKGojtirymRM7kwswNS3/PIEIHO
8ZmvSUzoEJ6nefWTIkdgc7M0mHCiAIBZNKXo7rshHkMXvf7GQcm59xnEuR5queCR22INHXU/wwnx
fMyCExldKTc4RAJ9ZYeNqj+s1YdH8ANni2toxbQHeBP0UgE28C/9YZt9dsT0Q1YlZPvzEvZjkvXv
XjG7/8iaBS2bia5wu/tG7CDu8IOB7SBesp4jZVdH8tw5lMhGRh3abvYLqZdN5ptIQ8cAYZ7ITwRS
m3rp0sknNT8YuIopUr2ZF8yHP9Z2P2CdYs0I8fe05IBy1IYCiSsXYuvzrtTd2U41lkJVUnnRUzFQ
OuSHDTbPkM5cfZ7WO0Er4B6Nr0jMnxzHk8zzelZwFKBsIp+NVnEvuN87Nr6OVW33vPXFMD6H7+PM
ROvUAjsfrUIuGZZCkQQVfWnZsggMuo7VfioI3jhxbkf4PVpdWqqGaJei1KCYnQJHdsxICLLjXFYo
xLpe5DlqQPKmRAxU+Hkawah7Srhxfv+FI380WHan/RJHKvmgiTGL4QC30rnGos8g2Ln7IMel1Krh
m1yRT1oMDdUBQ0vwLfr16VG1Sve7kEnSy0UQXWUimvHmA6H5FTLbT6KJ0xd2mUKBiyX1wZXZcj+U
l6IYP1E0UxkekSCeNCq2nloVGBKKQ5YJQFZi9ZS+ppnCVu8hrg47AD61BEC0PTO4Owi+DVyAm3E5
4FQB4ehDlgTu7d1veAEvzffJE1ctcY9p1rfqyiQJfVI156on5Zc7KGowrfUM1otRrHmVyea9RnAa
PVG+3t3Kb6wT2eor6Y7jxVVdWI+szdKzGHdNfs4olwpVSqx7o7lvkVgaSFpBDgXrphUqsCTQ2aDP
MNX5DQBFFNOw7hZE/xqVTwte1iMLmMGesf0zhSO34c/TboQhyHhG2dzD23F8asjx1HYtxMby1dlJ
0L4pYIJpqnQmsBkJPLR6pPeQJ0bQ//+PWwbGVs8P8BLQKG7m1z0ZIIoYi5ogT/1fZDLoxjF3hGqn
EnsjFqRsdtwX5f9Xfu1SMbKAzzdjWX6ofL0Vxbl2xHQvTLqiVzn0gd1+bd/LsjUMFFo9+t7tvhU1
oRtOISDW8KXN8Mx/2YxL+mne+2ukR6ZiXo+GgWhl0tCIuSZWEatdbK2ym0iu5h3M9L2wPS3+Wson
e9Mh4Sp1EeJERJHP5wNa6P+l9O+zn2ZiixcIvkpPendITxhYSo0lf/nLCZcLGGLLPXNbLB1GYSOn
Gq4EYSnEeVRp2OFqpCD2mmlvO/3pfBG4b9sj6xt/7gJvfHQnfHPIUfDGJHHKVM6mrbg1nFkVsnOg
4SlaReechg8bP0KDepH0o599Nau35mRgGS0DV4df8YBxZi+TC0w8kN1oIRY/uzLW4TO7NnSbX6Uc
u0HKy9Mie2D9ROmrMRiRQKGpM0B6rtIZQWnHLhVkYzjDpywIE1By3GtJ+Z2XDg+UGJYnJWfjPUrg
LwaAFhdW4Q5rpTNPc8i+k1jxQrX9p34ZFOTHGf1bd5F/nrQaCtrxvvmhqc2etoWId88gyAAeP5cK
b7YILEXQUrOaxYiQUKuSpLjNLHpClkEk7Xei7GFKUSQFU6WhnpsBYjmsRuZeIzyvDLoSL7pd1x/V
Cbcw4pRy1fh4qoMfLFr01dlgjpakIJE9hbFbiwNPtZcWgI0XlwfLY11dBduypwdxtcBMdlqZ/Twl
32+cLDNJl0eZxZLlbugLCmJKJ7ihiyl/q/Er9uJEAr/t0tdXcyMtOHeyhW8mAI3BgtELYthVJV5v
PbcWEJjA7LV66AcA2p3RQGRwf4/vYgzZ/vnK8/Hm1AxyeJ917SDMhEKAnT2/y300mcMygtp7Bxi3
wDQ7rTAfbFpMMQ6EzkjoyClLdD8y1poWGy4VgyT3q7LKNyw0/pvED7YgyxCNG7Fussc1kV3cGCcd
nJBU/Yd81+nXnKaZ9U0qc6gbT/CltNo015hyRAJOH92xYHwDB57ICy8hAelZMZnaphSE3wZsIO37
jOEF+Yrv28sRST7fR1004qxgxrQfyS7YtdMTWCYM2d2xskgW4T6eAzU8IC4uOff0Fvqw52VvrFu+
Mw7F0IYJdRQMg5hbwIR51aUoS/DgbbHULpDwHz1g6PSQqhImy0xqz3s4oWLXt6FmssDZvv61UEMx
O6Yq+1rSj/CBrPFvu6PEKD2O/eulWCZsRjIBrPoJ6Fxk2/b3vvLUdP1k0gT2NBiao89KpHQu2n3l
nceTvR89q7E1ldYh+0STqEtjlkIhvS/mQXrKOx9g3S8QXy/8ngUxyWMbR8BiiSzkm/9UTF9zxECC
W7gUNrDPDSu9a9ds/JEnT7n7D4IMGXlcHYsGkCNEMferzQImuUKUJB9tKUI19fX6IRR8wi1hWM0N
9QFXDOVkyYuHkk60U2gZR9vPI1YSZV9+qOEShewOVXEBhq9/JC/AMW9a0hj2RZvOeaAKcBs69wIu
hUaG2QOcz+jerv1EM2ji2s5nfuEzs2p27k7obZXPXgnMewQHuxQJueJVZ3tjADsf/lcgB52dQ5xW
XzEKZdPmqqqqvsKsD05EBPiFkK01u+cr36jEXAwRshkCYUJLtcWqTgIVONMVisnygBX0mB5XAUMA
Irm3IppdxSyO5V1J8ZUHFWyGZCJMknkeRJDNxaaFhTXDs+oLj6/aJx+oUBkIzP26lm2mlGA0KhoY
ZAWc+R9wMqu7lG+Y1IBWB9Apxt+yPwgmVdmGbI1+GykTMsFNljeyeLfrSjM92lQruesE79WTYHje
cVeObztn+KeTv3zL4C/E/qYDDG75tVNIEFhhML7cYqB3rxMzARi+wX+yYj0X+YW0f73kw6Ug4EJt
z6z5qFtoyrzppyxzG9syHadTP2y4QO9wdzNfYzmVA9JUbt6/sllJYpLTKvf8TWH+0O5YKLgdZDB/
rYubDUMwIbB5SmuNH6R910YM5+NfvEkybbSB9OMr2KJdBip+SQxcH5cBGpcBzNg7aS+f4e5QLjAg
8QAjNqAlKWBD0HTjEm1z6B1/qmTRaBQuFx9J7bNjp5tP477/OhB3F9DjGsPHezuFbAE96qOaHGYa
+8PcvWd2PDSYMniurBvd1vemvywCSKMMgZnhinVkEd5pG6rcS+h8Ixe8MOTrYozV54uNFIJcTpQu
0KJWLukHDEqUDTQAne/y2/+/RWOmoWB9ibAa/qi/1UVlYn2VZaW71xKo1wcRCb5ZMEt8kB7nbXVC
mbHsBTdYtOLOC4pOJtLpUjRMguQDHpPHuUVf38PiXLHcT/+VpLUCVpnHIjcgSeRw0E/s/nDEiLTf
TjC9Ixx+A9qUKUXVwcZtA7biRpPkrk55Y9HlLzZn5yk1hAcVVCepn5UdnQZnD4L5/ckAngz2fb0s
k1ONsTsuNliG7D8wIuoMKVhcoldf4xPsk3BxJZ34x1M5nBFKuwtUpYOAaSxptNBW5eZpaWhST5Qr
ZG7rv0by0SVSMKmqaX5cj/KjGtcajYpdRmQxQj+dFpshU/bjKeHOKOZiGEa/VOWvLXuD7UEn+Z0v
JPU7+VCh0X96gY/B3cihU5tJqaZr2tjGP6mvB7y9YbDDQqDYLgeF4DblPyasBsbqlDhIS4Qefrb7
W6NC7XYCcZBzGn14HSRJCEWODWEvk0Zg98IrRQSHo4CGWM6hdidUtS6tZwxTHHPF+ClNyxEg+Nww
LfomhrSGFxDzC9ywIAXpMIJB92P+fP3eSjTTgIdkOmEqOmFh3CyaF98WmbaPaHpHBIr1pZkt4F5W
BIp4uvz/SxAx1gYnDld2aOXJwOj+y9YfScvvy/EyzBR4rh05FBZbVH3rmTX6hLg5GwFTNsTPFMa5
0cmXBxTueZiOyn8vRTNLiXxALTdE18+6KpqRtnL0OXKt9G+ImhVUx31NUJlUCDANHBwm321rtMhJ
cG2uY68Q6TtpaKuI9N379AUFER6T6QTq2aMn/y8+7+3Wsbof3rVrEHPt9fa47jfcAoKOI6RWBLLY
fRAJBujOm6cHT4mAtjnY4Y03aiF9airT/pPZaHvfguvi52DG0B/aFax4hwK26w2yhoYFt/+nq0xr
g//4LayY9fr5RbcMOj/IQsYNTFCKLn3RKt6J8OYOITIKy0LLfA0kLssNTTpZxdQ4yhBjy60Q7xbH
xsAIj9XTOAoNDxykPYuuve1USwU/L5N9pw4MKnutxqnJ0tK6WPQqy9o6XZ4cOduECemLBSUFC5R1
nIizZrgHGuV4iOAL9JLyj6PEQZhYkp/KbKIbvcd8I+CdcnjyA4BE8rO6weDEyabqcXlb1hjfB/GR
xL83ja+CTvyOmrdEGAVvbI4uI4bCXutNqx9LquJoo2TYxjHL0kp4Fmk/z1cEb3WczbYTxB+k2EP9
gb4Xbpw5rs2D28walxCxK+udNxTRMekKkyhIUkQXiSVWvBrWWkjk/gHIx1yRMvEsF2m8v9dclPKK
O8ZPsW3bOKofo6MfkfY+v/nSfM8RbdDoufukcNXw5YHqlLhBi7Y1QWLcw4D2Sp3KkXSsx7VgjNbr
TM5W4mFcyWCgK78H2O6OQYfF2Bp0KS2KWDJ/Y5LM/1ishFFsznsEUmENHdOp5liKYFZbkbuBom3g
6WuFuhifir1g+GtI1u78jXXmVILYhEuZ1OLwKM3fodk7Cq5+ZxKx9AYKG5A1cFXDrHb26IvrI3kR
7a+GyrXCHizhDDzhId891IUDPtzMeAW41r+fXDx1AuxdVoREpaxwhzSPrz8no8SsOV0x8hAWjmds
CkiPQBVMkW0YlU/hos8VYsFHmAgz3pfuzax94qf1je9oaqGkDLTZu54JJ3lfEB6mJ/Qz5zx2x65z
OHYLYx4FPam816AL+JL6J9zSWa4X+JUQ7eFplOmgZvH2tLEAWgRm2tP0I9XlBEyDAi5PqpS0x5Qn
AWJg6CF/X02ss11BlvKuFKFMIlRbZcto52FH9tkC1Y+6ibEQuXG8mp9lz0HXj+GdYzNJRAmqZES5
rhdg0indSZRQFyh4oYEDqZC97HkkqFBUxKOT5nLeUWPC688zMr5AmQiL9WXZKBmzIGpylIRabZ9h
BMdeS1c8VPVvbzErnbsNbdKENOk7mvtBw0MfdcBCkjT8sFNi7A5uUPbiOACKsbS4/Tb6R2mxSuXP
iILJF9mOY8+LnZbcFC3bwl2/RBYK35/XFm47t1apz9xXQwzc4DYe8uzu8kqYRTCyKDEvZwh5gGUi
lcaYeS1EOvxVdaFnb5X1e0rPMkMdM2c373uI3M8GpIdNymxsBxBZJ4L66m89vyjdPX85ABAD1MZH
0KEbMYMBnh5DVOvwCJcJzGzFLEKrPT25kdjZK7I65iMn0KQbCFrQw7mF2X/D9YKnq/4VvRlGkuuu
rif0b8RCNYUBrbRoUJsweP/SFgd4TjP2Y1wsChFniBbfcrGky1YozNteg/sTOW5yxr6FxujbkcRZ
+yNbPGS+SfU0ttlpnCZBipqx8Z7PG02ghv4XY9IzWgIFh5Gag2vDHr/JHxrPbObXebsM15K+tjvt
Hq5+3ZtsuBEzBC3EdU/iU6bK9oHt8dE9oMzwv5T0g48BZEwEm0xWlSLnMeDM2LLjngslKieX1Zei
L6J9iUXOWxmQYNedXyPI16VJM4sFFIIQAhcbLiz7jFKNMZZvuSLHUCmIWm+CwDxTwGp1a5hTKf+F
Tgtnotturq2Bx+Cf8pA9aEX8V9VXt0IdB3suahUdM2d3+vRScPu65sKi1NIZHmm8DhqnoadCYAcM
aHoZxx4wGtJ9Aw7kwQ5eF+4RILdHzOxy7EzE6hGUZYhJF+Gz1J/GS8ienLQNVZUeIbqkJoWwW9z4
wpEH8SAhaWVo5sEUpUD6REWUL6xRiHlX/qeiFqshShYVX28+F2VGTceQfdEvba+Uqpy91FocrwVR
6hIkA4r+S6EyABNVmBmtnBoGKsdNc5dtLXq2KLNdZeZJ9I7Vjm8Ukelgd9Ed/gp143I3AVMOTyUh
/wO3HL0h0LrmNaVYqWOJVB2c8fpler1YTEjloT3B3WrfYjNbPak7THir2fKX2NfH07DQO/XEFOKz
kGfXldwkG76+oiVAXXZBjqDl5XJRS4Qq+CQFfXDXaBVVeo53v6WgUdvLIzMdmqFRpQW6HOF04Xax
0Ru5jye7UTNqCfseU1dghOZSeACmB/T62t1v703n6nq4Q7oq0fCGbdxDpd9gKRTBoeUB1vPcNUwj
Qj+H2E1SKLFORW8X1Y3vFhsgAtiWAsPig0P/Kp0VAVLX70UON8Hix7vuyVMdHkPbGhxWSkCQIv0o
kCMZSBLRVqO+HcDakt89e19GFOYy6vDpHOZB8ZtV6VPtLY1o2pbz8TBDOTsXyRmdRLYvuHcMpNlr
X/6K6cJTWMSqFvFDyZyz59j0ozlc9eTsV4nL47IoHZzbXQFN0gpYakkGns8ReRCCgYw/lYhFMqrE
Rk3ktTBqyMnkcUSUqhOUoNiMEpjR+LfQkN/jFayoaoDwODwAaXy0Hjk+Dt/qKrO8jy6QENagRaRT
MhGl0Zv99/rV9l38z6/lP1TjbBGJcPLXs5mlQ1GQjy5RNedZxiQB6Tp5sLRxUdId+ipRMuIPb5H8
ZhKTs0Yb5KxJHIiUl32O97lx0LSfSWoAnBqOTC35jwR6trC6kRoNfgHGZJ6ckhQrpFxqnrp0aCzl
S4QItb3aWKxZMYY1Z/PBDJgpp1Po4LNMUsIJckNupzNBoA0p+gXnh8bw3w06k+fJn5TWWIwzJ+OC
xPvI3TK3vG/Mpl9eMxWdQZuZXSnyqBzmOqcJLpMx12z7DeIs8N2Uqncl/n84Y0eB8k27LYWd4/aP
LGevKLwKHDiZ+hNbohSKq63nseHV5OX0NF2SCqG+2esdRnvmDQ9SIDfcgwXV3jNyn94y5d015gWn
yvj//TgETDzRJxcCsJUiR/1IM8uxkMk4IaoeJk4O0vl7QjWqYiOj0rGRZbRTL8VP8vIRblKTvRrM
cWRVieXQz46Q4d+QtOoS7YhcEvxCYsNKRvIQVk0mjmKYUoDvb7x86nqew7JeGLq9JTYjzuygXNsg
skQZNnrQKMsbI7D0cZ37E16uPgpsFmfqZskFgveIYFI/tLUSWXHD+pRqRY8FQb4rP3w0c9SHU5Fr
5zzYgqJz3b9N5fbFOwPAOXe65CzdnyM1yoHpeZ25v80k0YaUO0hKSPfqcSLLqgQ07UYRs6/jktub
dZhcknRnZNREtQgMq+grIQF3N4/+P4ZDkNsUgQNC194XaUdj51FA+5dByU+QJt+stgTs58LnKMEt
DQzfRCqSVTQIee1rRD0/eMPGDFC1Teqdf/Rgu+mVTaJLC/AyUBxycSIbqUWPqoD4VX2hvTrJB4na
YMv4Zv1fegJ8/X00yeAsY6+/vUbRASTx/RMcFxRhlZDxB3MqDH0i+MxECqYumthVVFFBCZPE3CTi
PD2Muuswp3eW6zXtT0LAMC9y/oqIxr2JENH0e2w5XjOHw7G+Fe0xekDVCqcBlxtNvFpEMlW/22zB
woQiz8JketRwDr3x6tR9Hfhkyy6/KsVxrowCwxWHf2a4e8op3c6hwMwHrxxeU2aouo+M+68WdH6K
wrDf69Aa7oMRw9ZEkz8EkNvCHKsk0PRhL+eTFQsv2RL5WlbZ0hTGTmZetXk5m19SblnBwLjWBESJ
vbCiCj8TlEsPitC/IplQv+D/FV+3BCls585rTEa/X20AqNhq4pUZGn6yfW+eNt3nQiJyrrcCdKcE
+djPUyqSv31jJBpZuLWYITaBAkz4D9iimN4uTN6m6klL/41L/crNR6af/p9pJWXPfDac+Wu6VWwJ
3yvAkV6TksRUAmJutP0XCLsvWfulq1fnlRgC6vmAI9hBMvjI+3IckSsx0zdunCU3udYYj3CyWunx
mHu/tRlwZzPaKhLXBNmccyuLriTR+ns+oPqcH/qeVSa/oTCuh+UKn9vczhjxJzkQkH7X918RBHWN
uiJ1y9RV3HHarkrJ+ijQUmrUNbPJHxqaPze58rh/TGGOYpG/N2hC4ki6VNABK532vPfzT3aYWtkz
uaWlCpU/9KlRp3lMbqm8mW1ndfU7i+h8vwlDqVSRVbmcYulFN9+CTvJhvII+esGpeLvJeHbLC4kb
XXf+WPlbqzgrOwC+poI/dnPn3Phqr5peVvtYo/j4JK8EeNRbGp7ocWTCaelpfPw7OLjXlgFEPmdu
QIWC6aVOk3ZDkF8lZVPNh3fmJjH9uTqfIhSHxu3VpJhWTufpgwcRKC83TIU1BwEffU2io8iqR0yh
zQl+DWxpmQX+tqSb5qct4MPFHBVKP2HnxvQNnK+Ej3wLywx1+SHw9vkKQLKOh7+AIAeL4IYa3UfS
fjEQHJaLg8EmExXOxbAe0jckY0ht+4kwa1ESyorlGx42vQaS6ipF+VPRIFIp6cO5P8woEFeBbG53
eDk3Il0efVrdYjml4DHCLI7F6Ka+F5giSjlxdNt4z5b7+XwuqvgvemyPePvPEvTtqCKnbH8qgAcm
pT/tvnPBG3N7undWKdfiBJ+KJ3qwb6XS/tb/HQ1r8O31wOWkZ7k0NrwRxrK71+2wSn9TOqfzsfgV
xWE30lYei+9mC69/+Ikfuw33XTns6fdu9RkcqQJg0CNtr1Vw7jJdfosM677Ewo9P+zHoPryCNero
jNx1ptI7tKx0mecMS8Kdoh0qVOg35KHizVmHhHehzNMWWHs+a7t/qx9zhbQsTVz1KRQopBjj2zTl
+EiBnKoyZekKIWjWIowC6T31qK5dHX6hKuuTnGHg47RZ1/dxylUUK44s/kGBF0XhSeSQUPim+aGc
LIMcUh+1M+owdOTn6CFh0HYaQTbFE/fEjvRENxY4ilmOPEpJFGWOgPlZeigdKRjV9VogWIVHVNvw
BYh1PVeQcZiyDLuvSv5T33SrzDVKGSPMackHEevcZ5aXy20X1cWJBiVFOKkqFUbznhGRD5Y2EdaA
cFS4eJiffT9EZWtxbjtCQlts52eU/dcPoFjgd3x13dtjRj/RcHu7JXbOTQIZG1BcSjdnNoOor7ES
GEstr2BzlMwOqeR59VbXUoCY5w5CTzy+OOUYAg9AX1EJmRTYRFkp9KFvR0M2x+yq6SzVQK2WlYes
0RwTN5AB77W0gsfbaiwpX1RPlqvdEyztYHu9rBGmduKabUQPWt51mR19i/V7EK5pKT2sDiLJSl1c
KNOydAyUPJeo/wBkkjqwTKK3w/EE/QsGk7RC7GQBsh5kCTarK7BI4J9i9Mdpj1OIj6oiOkrD0rfp
O9z7v8gYxj32oHwPq+S9tHJ4Kg+IKesOS0bg13C4TnBJm/zLRXj7DR4Ed1dG5yMqoEhHym92Lk2n
MV/4Ky1/GG9pHSsJNBpY4x0rTY8sxuq67Q1iHfzbwA4sK+z3TpDhm1lEfbvmAT0RZ/moHDAM5w/6
y24JrqWKvSNVeor1+kvnvCR+AIWFH/cJZBeuuznppHYfsNRYBbTagrsdPCmoAJ32nwBqLz8tj4Qt
v5lZPdzf5mzXk/tgYQMWP0vtDjS/g9Gj3VNB5hY81wVvFkE98Zz16z2kJxInex69m68eBTwIWqgo
exzUBmLgW5FwDULv+ao/J9g5Q+jtoYkFxSehCVyEJYqL3DMU8gphcIDXuTeF8Lqt52VG4K41jK/Z
+N/JkgUrjOyY5qd+dXTDFVNb1A5mORSRNg/IKVTi1ZR2hu6ARFDoHIu/paUvCY+AMCzzcqmkLr2c
oXidUie9G9MrqIgrSt966D5p7vKHyljkpf9UvwF4V13BqlwRWYXmgFXBhmdnXm457S7hAqgYI7yz
8K8Xywa8UUGWU1jTpbp+7d427Djon9WnhOUNkI1hjuag9xO5OSEx1CYbwMQbiBE8aOWKdxVYqsUA
GMGj7azvCu+Pkr1ZnweGTyuUnQv7WrpsvBYRq/gG82TxAad8ZIh63F313UZ2uW+vlDCWghXXHDxC
pNEUEgku0F8bJ08edp/X3YfOnSKnRmeCXTkjfjdwvdeS5+6M2r2tgte3GcPtsMZ/+HoY45FbA7JZ
sISzL6RPV827N8CQwCSdeZ+bmgiWIQnxUU+NzFkb/k6bKVgbWXJaRUPplbVmdF5S6E558AGMVQjr
tn0akRGclihvh4o3yoENw1DC884nfSYzRS5LFRKLkgitrhrMud9qrL89A+BRehdzNYBBN2WwKT/u
TbH0+hkZZz74TLWxTFpC+5bFFv5LAo3Pk1uy2csDv1TWO8uQ3K09ombUESW/aCrFUTjPDzo8X6OP
lAtm7WEmjpBzvkqPVQoJeRqz2uMHzdXNQuxZpCWRaSdZet66dfCVBUDgMocDBRcExrdO4qcxdJGQ
+YRVGoxmO7IMy1F/woc5aFWpppXm3LfExLGgrYuRJLGAM46d3xpmHA2mrR4T8mxRa5Q8Vp8cbI6o
sFZz7RBbj8NRGTxs80wY06Fbpvc80v34mrF1KZMEDA0bz3QNGC+/Ra5OrxSGmoCnynm4JoMuRhxA
mpAZGTCU1zY1fbhUJtIHt6w/WlZ5+Mm+gKIbEDSroDXejEZqMLSYZYCka806SLC67aC5j1mIjW/E
ETrv5WZ1h/c2XUDVAzyCcl3+LiGTNb2D7+O3rrPXSU9lGw51DDH+AOeaI9N82FPKUiyq8+SpVR87
vtR8+Nd0aJlesFHfuP7cyMyftXdj43wREcOIWfxZBs+a3WC1il6EQH5cHefC081wGQrtJ6oXZWTm
t6JEtpIm2DlJXztoJ+LzY/sRyH0UeMiZLcCIFiriWHKwV4v9efsYLGwhdES3J+eY8Exd8ttbXbk/
SNAzoAwPvwY+O5GtYs3FdM0aerRTajOxzN/cqu+NOSZtF8vx84eXhMklFzi8KlP6E71QQZIfJGxE
yrvskfU9gcXsNvK8giiiOLcWEoxIg/M7OE+NE9EMM3M4EV0ok1si6fcVrmGUBsqCaEuN2Pum5dtU
uGPucZrsZOgwO04r5oNGgUjrcTRBTCUgg8Eh1eSQI15NQnK3cP7gVtJsN2LDjkxT02ol8tZcR0nm
TZWUXAXPc1w8JpZ17qWALdz12GzunoD+XdJV9SsgH2ixUev2voVmGnEMBE6awVimS5/x3gJesJT7
w5KNxo629IHsXTEzTBidK+RWsbnVbaAa9DCLhjA2WtGKoLjA9LIGKLYnkIn4/IYlM0RxJDrVkzGi
2xLXpERR6+dG1EotLYvNCbQHqVXQhiRUPIsqKn74jrRK3JJkYi5NMyeopWn0f78XOvrTz2LBDZ5Z
CLs3qA7DbaUh7MclR82RCIOMElHsMyPa5T5KT7qr1ly/wTIEySdeGbLBu7qwBf8D2ihmguoFrNDc
uyALIv7EW6Q9HC73d7FK4Q6AEYquvopvQqD65h5BLy3NeIYVhXTuXPDeVeMBgM3e3FS/Ia6Lyo5h
ywKGKJLwSNk6n3KgTFipr2CmHs1RdQZc5iRrfQkTsQtjT/vwfcKkdAQBbHY0Kl5nZ1kmC6bino+H
87bMsvnDx9Gy9OwuZILEr1r7ggQheRVi5uRkNQ32gD8Xbh3WKTbBDq5oAFKrlk0/03KHDcCqAxo9
dlR8mA8BXNHpfHLxdasq3EnEX8hlSIvE9llDLFhga7rm4UXC41/o/W9if3mcUB1fFSoHT06k4B68
CzOYWmJBeBHpSxV5LGjHyNaW4C8XFsX6T8+EA0dBFFZkHIdEpdSiKBY0Tx4Ji5CP1IFXUntfef6Y
NXykKjvJM5byHgrkPZTpoxU/14KStEdPQf1h8xtBrU3PTgAEO6o6BuUsIeKeJQn81dZe29bpSC0z
+OIuMbqractlM7xkys6KP2jEEelROuX+pMQVrSo5kiS076sFYWp+/+IVV/xwB5Ey+wzxKaxKNYnp
vMDSaKj/1pvwaDSde9EYVsmdXCC8tTVIWE3cD50kkYyN+wD799gazMbjpvCItsV+rUXhJNJqKVl2
rVLRagJlt5WtoCbudnedP6wAxGL2xQUdf37RMuKptbxNaAYazw/h2mVtJP6QlDIli7yYiLvm19pq
5wZBhutCglZYbr6tdJIZUYT68Zn0dkZohoYiDn3QR6micJsXIyJSkUJqRGQbnxBi2iALyegwQRve
Ole81ZvNdnr9TfZ4hqoh6yQTzY2kr/zinz2avs7Mma/FNAzETBbqutbXzrRF6qMlQPvwu0DXA55n
CgepB9XiSfM/e8z2+KESV90DR6X8p6mINKOZvUfMuMlFqpXNUSEpEoFY6gA7LdYB1OzDluzZWNQT
F9PKZ6qyh9awCgwChBzOQ1jzHeNjRYUsg3n9kQ32KxNRCtNhGdI90EygvsiSOUZkkoJPKNbGrdnC
wqrVaPSCpQqqLr48EyFkyjB4Bna52VUrLooNVLOhDT2RP2Ep4AJhdtwUg38xCPl3NLWqBRfEt7m8
XpVkBof/zB/x6x+XdYjNsL9Ep4h/iZQgAXnoKL3lhYOI/i8AWw4Ap/L0eHviXdR3QTh+s40oXVNw
7gh9tSHgGv5aadJEqddvYcWWMGdnvlT3/t0vr8jCBLC8ML3SunGYeIXsrf0dMXUJCakA5kn70/0g
aXD28QHIp22kjw9MhrMSEk2q87SfNNmnS7NOp2862URwb0Yl3Xw8PUsNzO78qzo1oeP/4+Xnojnh
ragrJKtYdFl0sBSm1dH0QWviI01TKwEIj3/yYTBHYHSIK9iPh3e4aTRychrn1sC5ZR+nBxwvnXQP
R18yiTmKQxmnHujJoOdmXhLlEVUAXD5I7FVBKqB312P1fl7IuAg9xLl/fN2cy/aVNN2YRccQaDQo
eVXXmgS1abwsS0hUJDyfZFJTZ25C1zdR0hl1kjpBnOwk27eNW7t7jp/oZQMSCv1pVk79QXuEAKoa
QjanZygK965UJof0FZWfiRRhSWVZDaIDFAp7o6yuxfspxOx1z5LIvgprYHUYuujcPa+b9XEHtMAl
AdUHHc4n+JduoaxMAxlL8KCz9FaUAs/3bTG5fbzUs5Rt8hNGI6pOdew3HqZat/JuR4+4kP+XTkko
DDtAp3oOCY2NjS2EHJdZSjSRP3cv2uRZja6Lsnstj06XQ8PVF2TVPsPRZdXZE680mOkZWKbnEEVo
fSrX2vbcIcLfl0ViQ+/ZAlKUXgvl0OcQaVA8NCuDIY3u9TaOF0jr5JjSQobngjcyTPDqPfuKE0Z0
eg6U3ESujNqSVv3wpLfQz3RYWLe+gBD/S02mnLQ8m/rUwsRwmjVmmMdHAkYvX5K2JM/2ATAmzB9I
kA4T51GModGT1/ITXRFxkhHXWQkKd61X7ggHjVR92+2oiUle4dDqGOdEqBGdVwY5nIoquOt8L/zG
B7tH6TupzYTwDnvdWXPpU8yNvnt1HmroltDnq4GUr6D7j5Xo0sgGEew7f9fwflA8mQBP+stZDumc
iG829Q1PAiuYy2c6goeTvJpc0bUp433f3zeqTAAoSAoQ1k5CLr4QiYpuC8NM88O6fSTbBz/rVL7+
vPcmaHrhTRRfxTutF3vd4F+/RtDnxN+K5A0BKFwQ1j7Xe7rFRoJktMUvxxx86MfhwXHgVUH93PKb
1gm5+eMXWmPom4C/lK/mmMTQyMSTCO71JkThH2uCx022ZLLf3+k5ZVM87q1Q3BQz2trFSA0g1gjI
xIQkrf1tC8sHcHaMRlzKFbNKPEW6xvH3Za34daB0wW/6g00TQeBHFaJLwiMFYkqgHESRSBzt56Ng
FeHVO3ofZFH1By985+88hb3vZslpUzR4Q73yYUeM+m+49VPr3GQsKrTt6VfPk5NlejqQnboJS3ZG
Lo7RHpMYwa5pft1PIo1GOf0coZn1RjEYbepar7YDeqms4R4p+4Q3p4Xk/HRODepY0PjHvfNjV8xh
GlnqtiJljtFkAyxwUMOjoDLmis3qWKQhP+ZKQYkGov+iM69EmF8RpWmyCiAIbW5EL5D/jL/0QZWb
3tZvBxoN783tgOspabs6Jfz5Ol8m84auejgRBlob9kFh1NDGbT0F1l49AYJmk5IrVJIyoOiBc5yv
5HQDA40y7hb5qEwh7rJmQenv7U8KqNqRLER8GvF401Af8IpyZvkq5N8LMzLlJWAEb3ygw8N8hkq0
RWg76G+svuyvfDNIo2/7Q7EJpKRAwD4amDFSva9UEjCX2/1jvmzfHv2ni8Pj6NTG/ZfsPX7uNmoV
6w9FZ2cFkesd0bw3D8sdkXrp5TH5dyumMeJ8s8FBNDvNHGd03okIJY3hF2n61r0/PZ0A8bPqE0Nd
2zFvCeF+iy4+jyh5TCNxE5kHA1LzjZqgs58SD2JSZtKbtKulKybwlxZbHjtdLQAalHie9dbsh1Gc
KL7hzMHNMbvMMvDHUVoLrQIDjAC3sGDRTHWjJZsMenouxwEwUKnWxy3aCd7iok10O0Jrq4aPxsr8
KthiHGrDYJfRKMejjYfZ+YGQflVs8QkGS5QpnxB1ZTGyzgMOrTAtgwNLh84Fa1yml1cL5vL1Q2Jl
cgQu9gtTBJz9+D7zIv4hodMkM74xJ7gXtRf7SKc9oOXjoDqPkeW3ojM48PuplDHWEKHupgGakq/j
2KbQ3oeodjO59JO92XV1CR2n03QG2/T4uHmpeNDv7bLl8iXa5LaNqzCXMqhwvKHfanEuB/EPkRlI
BqHpQ4fRwDI2yhM4RUkgnE5XqS578mPtwzQv9U3XVq54kQ58rbxnEKc42ClV6vrhJZIAQxJi9lSu
1EcVvbzcWF4tMJvVgcC3XCCigXp1cRbGvl0pWNNJna+MEtdn4eyrTh265mxObWtiP5yvMmtNs0bl
wZIvq9IO0WENWLTfyZ2ZM8b2sMjbLz6bJOTggmb0zU6ZoFofWT6EZXEhxCKNUJDIpeWoOAi+f56z
+zs4C5HjL5jrgPcHUA0JH1JF6Bp3TDtaVMqQ0T4/Mvwq6BLU50IUzImByJZQtMG9IyO7ILx1aUV+
9IR8cduR01Pef91m1I1F6cKqieB9E4HTD78piZ8RyoWJlAhkbT1w4a4w4mSGGAM1hwYY5q786mUs
3xCEHI7BkgCEjutEbFR27zuVPPchm3VMdJTM5AKA59PNkHwOtty3jT1A92jdE2oCAz8YZ73jq90w
rpILigm38DLd/GmCb0gUX/AwJRFSUB81jtRThs8Dd/20nPI2sAFNPsvD1IzWX3yF3CdJIlgd6A4O
A+n76J6+aCDPZ35UK5r4nnhig/DZlwPpgCgzGGNNauVCOQWD7KCibubvzYI6NTBRPrSe0AY0Efp5
DiD43ncJ8TxJEILdxk2rBK3gI+vgA7fDa4Bo2wvDf1Z/u4jSKzDNX0Iw3pNDjPmZrBJ2Y+JUMS+k
cYZ+o9gsvqWOQJJLD1kQrLbOgurGaVsiXURKKxm5j4Ye182mSHHZWC/uUOEEOEzo2M4fGnZmFYyb
dqQdq09QQ0J1HY219LsWeg0Uy+HKwFmNPGl0lJFBDUHHSFey9U2yqLCmqY18ddGgM5U1AlhVp2n1
ga7yMi9FHKnlEMG5brajpMCp2w12yCCCFPYT3d//ClYuj2GTeleTuHclgI9LjMv5iLGSWbHwPHoN
fCEsPILK3N0LoRwWHHKTboqOvWf2zCkU4r6QFWAVQTupKnmBaZEEQ+B05Aas3GZNLyidYtbypu71
fsS1wSFIrHkUeFiHwjHsSUJJnFJj1w7DoM6CMSymNSeYAJbcYMIXah40S96UkrRqv8y+JQdAgR4F
c1F2lzXpk76xFR4cKhS/NioER/fi6KX4NqhSCYeufMteClxfAUZLMIyyOsvBM3dixvG6JsDYx9tv
+xQZ2wEQvrWWHyoHpF9qIHEKvSgAgi1zqvRfjXZz7+PTDKW5vFQTJ3Ym7KiIavNQv5II1AktG5j8
sGh0z3ii/axSMy3eaCXTLSvzpdhd54SIhFlrdFv92Vb54MB0GPJF8mJOnEouW3As74VkrCHIvf6A
zzt48r9fzOIR0yf8ISn5SuDgNWNDTdrsVbuzkHRG+waavnA+I5LGDAkTMlKkyByfyJz+jbYwWgbg
5MpRg47j+9sRn15bJewA9R0inAtzrBqBtRaXga0h5z11gc8P/3L6SAHCCse2Xliy/Vo/WknfMrGP
mZHre3n1PkdaAONbVR6DfZJLpnSUu3Ej7ywYm3y4XVxiTUxGSjNQZHM5uxJyrVpS1vSAuawbvlmx
F+YUbfLQad8crI1BCu2UiQyUuxF4s4D31DmEelQ39shkzzi+/6cA7ZYM3ZCM6W1VCH1xegMJXpRy
NQ5CZUG5Zjkc6QGByGOeELTZyKzayZ9oBMJcXpTZSDqiqjKvj1LCg160fAvNg/lEid5CTalYy84x
RqReSXSinLkOztlb0aL6ooLDoXbCnx8ysTUaUjawUMKfzWYpXDnbwjEJfvrxGIVvzKfGJTXORpma
iSYwNDtNbWesYJcBkG53yKRXxDskTmnquBAedgilVkerhXC7Acofm54pyzrOwHpI7JFgK6G9aVdL
9Ad2ME8jQqptctxuLHMTuVyD7JJ18IJ5hdQ/c8quSixQkLaa10Vw5Oxatfh5jKeErP2IHU29u29t
IRpb3nPMJ7QyUGlSgLq/eZTPG+5utDG2bjPFEbNlJEn9M0S6s9Gorf80Xool7Y+YuwDs9wD6VluB
k85LVbmpONA8+wLBINfGKCft82Le5f0cxDHBEBsoA0iR4L1vevCkG3c5Ajxs5cQZMh4pFfhe7K77
wxVUf1hHf+doMS3MQb/2NxYGguDYpGsV24uIjQQAn1QJ/La1mruLlfDcvKliHhf1ninSiAApCvHP
16K2HT64JXiKeqVrYopq8Vr2nnzUGYxW3O8E2PXI9oqwZs50xYmpssjVexy53HqmNjhq02xdWX1w
/U6yZsR0HYvUsuW+nuB8iqzgTu9G8PxiIcyb2m7SYzIoSsP00c8UNcad19x0cAzSRBuJ5feQ2FzI
8DrOrjRlYlpb7XHWqw7riRgO6SKbyFIaW+tF7QMhpIyjIU2vxjLjtmstNBPCuiPWdoeTeg5bFYdz
MS2+4U1lAyOUwFXrPgfvSxkyLDIYYpSBcSnqLMLZX3ksmIO6qePFapb318EbuKoQnSc7S+yp1pR7
e8f9DQLhFGjNW2+VPmDi+XTL2r51Zm2C63Jrv3Wy6EnV6wIbx8xBLTNZZ0NeNdfR6NI5YJ/MU16L
zfjqUUPcMs8ABE46dohU0hmUbtIxUhhCOYE/Gg11Wm3X8pWcCGiys2qZw0Zcqzs8gQppo0239t5r
QUG/OERg7X/eawhfTVQbiob0SgznorfJl5+vOBxokgzB1WWlFnglmAK4X8XGOKLQVXRgqvlPlbz0
TkzTd8iyWZLPMPeWOR4=
`protect end_protected
