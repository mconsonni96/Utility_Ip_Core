`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
FsZGBIErauGWxM5tEmy3hye6B/ks8NJ4MgfWpng2NTs89Ogqs7bT9eqTWtTIJcRjIFxBUA8TYVfe
+b/6d8Pru6M9pTc6LxV6QCvGot51h/TsJdVualiTx5qwC8mPLP+wznMOeCbkwRyCG1+srBijA6r8
AH6PXF8HzH0QMkXF3enzQly19VxAbkQkgo7J+U2rUlgfEXSZmhhGtT3ENK6PfUpGNYNH1JokO92A
Dgk5GDyD2IGp5GM8B5smqLqJkv6Rs7Wj0es9am2NYkyzSW32Gzx/IfqZnCTVL7+pNxAQOMvSkSvo
/GaaOpY+CHX3rKCxdSJ17t95LCyJ+CsQybF3TQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="XuL11lmrcbI5zPoR72dTm/3ELv3al3vovXjUEQ6drO0="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1696)
`protect data_block
rqgh400K6RiAqq36tPjsZ77reCg28nZxkbZJM3jR5zTDMinB0nI0AMzJZe6f2v8pcFis/O4REUmt
lOcwS4ynWvaH2kGDJD6hpu1e+dYPcCEDY4Q3VSj5eFki/UIAFLKHUktyFQkJx1xx3R8wgw9CP7jt
1B8A5AYiRdcLzXrpmQzQcKo3MZ8TaHZ6YYUbkUBbxgE6Cole/QNaalbk2uw2we8zPSzXylFZWl2U
JhOeYghXdFRodaeuJuCna2OcnEq1AEGDkuqr6rx47G+1uAPArcw1UE/7Q+iygUzrTbJYeHimfz/v
2rHxmOIAq+Ad29mJpTyz/PY3sMvxDwnqFFGsomJFAkjrOQTWgSvLLKrtGo+dYAE9vqqsEf2jaSC/
z+MY+tggQW0UX18QXiARSqGGW/++tnaiC0Xr6fL1VP11DLYAdeN+79CTCN1oE65xry34gcwZZbWh
fK7+xa95/dRi6dIrckqLz0OGUmQAtIC9j9sNZx6EWfagrLrNLkmVKVjhvMxXqZVNiRq5qEHIRiyy
B4OqNi3VNxq7SzEtz2awYD8HM7obbq3AOfX95MCkhfE1gMKWP9TwQzlCWveUQuKgRrNEcmDUiAeO
7P+UyHt1v4hkd6i+AwwpA7+utorBxgVbsQcVdz1pUYJ8b1n1lcciGQFKUJ6JFbchHsnEY2AuX/q0
uv7kVbb1TRL5p11w8+u4sj30lkQe3xdObrh0JmyvfSjvrXD+lbtSMU0cOXPkoQG4ctwTY0G01cpW
7zXzYGgJPG6kM4CBhWxdZbCR98jCHpJGQKQJkxkTDn8I7t74RVYesCb/3NyCW65RtVUlBHzuDTS2
JeIjcT2k4A18lhM0kWfVvApKcXTJTUn4fsuSYlqljT94P73HWzzZZ0VLqdqQshMQrcUTL6UE4U78
UChuct49Z67AXhwvhaAukqDEboojlaYGkpbOPmxPXt1x9YOs35aRZ7k16JCvatupJyeNj79lkT2G
7pBvbiBvr9ZrEm8BYiwqvKjIm+hkhcjddlk+X0S47E/zUNBXTEI/hYWloasVaFXzbqvpO1PHc2lG
OfXC4Mrzb6k6Uj1YuofSJE7u9CpXz1HHu/99vRIpz82fyjNhGOjqXlwvv1nf8mJhD+NGznq1MXsC
d3zwYipsvPuOqbGQyQw0bwWUk1xQUkXB5hRObsUk//15Z4nUZDAB+TVC+1ymu/evTovY210aS+ou
w9SUBa/Inod6iqv9OB1wWMbdDaAXw737/3JqzjHjaimonHU6BekT9+scVm8emw0av9ucpl0vRZs6
i/v0DNsLXXTD5YqO1cQi4i7RtPtP52IJJckiO5cBA0i/B0nDcFSm2DMQyLdQ5L3Fo2u1dxDuhGk3
/8Zh2I4MnuLKPAvDDdv0R9uTT8COOR/G7OpLpuNKuR+z5qHb0syJ3Y07AUgwsAQk/YQlev6sPinL
DekZP5VCfvYhQvajFb7UAD6chE+ELgyfmy46l/hSUUMxUwt9HO1VrhIp8bu8t2gcKovVGLxKvaZD
npv8jGH+Ax0OgpWO1E7Om1jgZv7w/pMLgbALLiHMgoizq+kzzxFWBBtkymDVhr8iX0CX/RAMzaA/
E7S0Dl8KpdMqgSMLHu++IYUBvUf4g/Nu/GOkgzaRzaADcnWWEPVuukbV0NBmSXLJfmT9+s/izC1a
y8ydaE3VMZDnOHjFizn868uLO+tU8o/lQ6PaigQKvUD5oMIjLV44r6eTyReKrKRn7wYIr6UMBFg2
qRZ5VcczSyyywsONUPrbYh5RNUgfIJ8mI5h7j8C0UU5/cs6aLtH4ie+uY4Ubbas9Yp8/pj3626Wm
FYP1Wv10J0M6uAzXKA6IKyKsKnr77f89ahcgca3Ns8WMxlyK6cgIsguPk/Hd/JSIhwD0MyQ+GPnz
HkJhjRw1jnJ43L/Xchj5z/bkvRKPxgipOKTlsW5Oq4AJiQVfEmVIYjmct9Qga1N9T7/AjbWm7pSc
Me4+Mzd6GI+g/QcBSFQvzAu8vEhb5eMHFMK484y1Uy4ukoBRSs50DidIC6XO8rMRkbONkk6t4TVE
UJ/zbDYyhk/r1tD6c6093Pys9l/JbGvY914A2fp4YJUXhPVRSqfc3IgcQDP9hXpI6W0jKR57YAgA
iNyY6k7Sxc7FNR8dIQuGUISXeu+c3pENtThPtLjh6n+7KeaPDsYTmJC7fg/qAT5yN+ht7YP7Pw+7
L0M0LIhQs+DxiV02Na8OaEiREWOQ4lJDYGgDukNn3sH90nBMMmrRgn9L6g==
`protect end_protected
