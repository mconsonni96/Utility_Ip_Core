`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
QeP19Qj+jmVNTKtlVRJXxN27tQV2afkNwtaI3xosQeL3VGYCGvjXjn+Yz/q6K5Dvwy8ZHd6JQ2y2
ji6YNcls5uTkcV5tkWoMo1uddYcoHCzkjRDDOHjY/L3tLsydscpYUaoKRQr+yrDrAo3f/PS+ZVhx
V4UXwaDZx4lLCqIR3FgTi9teSYIa1rgPJrWwpVTgrL3MY/Fl6gWt8vJ2dl9qgviaMXslXc+ms40a
DaJOI0F57UACzt2yeyC1MMBXyr8BkN3PizCdT417vAQS5Hk6rdM+eBf7NX/KjlId+JTm9+2SGILY
hf3EnZGOnVlJFFhYB/xn/r78ua85v/ZU3wgRWw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="KfpItwDYimKLCiXI1dkuhcXrRtLMVNNbnKfIzM31Sds="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10000)
`protect data_block
9SW9gEa1hcce4H3kc54zwh/KHWenUKFRFQeyLEYNXLBHZRsaIqORvPC24AzuT5OtHEaVXR1kHva8
hdXNtPTsEO9w8Owol8l5J59wlNVe+gbiGXx2R4rWG5e1zn96mETvze8goqT9nQFIYQtQIi+uRG9C
bl8IIfdHNbDpoD8JsKZI3jtHwMOBeFJmsz2r0uiLtLlFvgjMoM5vT4XGl+CNTBLcfqPAtmBkad2U
7NlSeBPi5CYcvK+HXcMclytiGeN8FO6AUg7xuPMQwveJEyO8TDjHILWxZBZfdTDKXdsBGRjlrMqf
wkJkw03pMM+jcDN+EIEI6BnemffOgW9vrZe6YR0w8932sB8jSH4h+Nb3TyJ3WB/Fjx775bnx0EcC
2fNzpqR0XXKZ38pmKcoEo2a7vuFuW8mSGOjPC8TN3GCJRezjFLVUaL6eZnPNYdP0R4cChTZ48WaS
TWEpV5/xGIPh7gJYAnv/uyvtUrUyYYby+dLqZUkJ9JqCRolTekTx59F3fsBXWUvpUzG6vWlYjqkO
aNurbc29AmOTkyu678r4qPwvXJIJSc1+p+ekCLy2HNgYUQ8oLwj8SyXJ5DNUGS1qfVDymF3B5EI5
XxWN35+NKrJ6j0eG6obOfSJz9eLlxMPm21C3DLqwCY3NbG37Cup9J4KtfWHiGwMgDPRsqJbXxRk1
rzXCg4OVhnUcD6nDfNkvFsrIIvcPkcLStI8efOKixg5rIDyAQnsphzVzPYG9MX3HCR8pAArgOMYp
ghlca/nCaEKCFKIWhN3/0hHJTrOwbFihXVXK85Ii3604X0k+l1Jgek4Mw2g6oibWVG5kH9ta3F28
R5p9VVSJS21eVjHpnbx13C4Irty0qcx0Ws/O653oXRTiqVUpri6+KXAVhFAmSvKMS3m/NNGXLwdN
Y86+JxHAobfoMmns57iJBx8Zsg7oYTakAfPZvvn2tp30nTX++2UaKa+TYHe5ADlTL/vZ7xUwnkXV
5zWiZkqEroJrvZ0gh8SyrfDEjzpRudjYqcOKwraLeipcRZ33Ojcm16K2b5VPor+Cr4TKX3ddcH41
FAsy191JsL95hBH7X3gi0QlTaMP49LsfvJqd7afwkTWapxq6uDq7OsWBfBK7TsyZr2hg3dcpJFZj
TQEgCL7jmqUTMxnEUqP+VgxnmdNXlCybjMt1I1SGn2t4xNUtjp3m3Kk2xdNg2zI/mzbOw/89npha
nXl1fsirCH6tZ2fyjCVigt0oBOL4Yzr3HjhtsxVrH+OQhi+btCZXgprbdIfeotpNEUaGsuyTcav4
Mlk6EK4V+Y3thmxBk248T3iNi49x3YXJCug/xoVGuXbF384FMdfQ0jWbbdOnCIOULh+k+nHJGCda
rKQrYbg4NeMnqbXYvC4LFDebafK9Tmm70rrqOjbyuaaExz5SamWTyMbSBWSnmqQ3GqjEww8VMVwv
SNnNmvFYbgXZMtPrYi0a+yohH3vWSvFyZ5DZZNSC0Iz7Faxs4v/tg91ZyFyW7fnE2QHsyiUBRo8w
EN6UyaiN+AIRZI+Xho5IChBsNnRsE64YTvCPTfGYadfkK139+K+t2bRfA94b9SRNcVEGv2AjVOTv
aG7pyNTVmElZd7i+Xm/NmRi1FTun/tcVDbNv4iMg7h/f51kr1uNUdVw+SPRapoe0tfmYfTtj/a0X
SEm+G6zn0MjXiRKdbqfeyx8OadohW7DsHM3r7NTcVkyCAk2rjYUtgNNl+3IxCCMgaMrvKRPuhctc
3SgLi3KfIqxidC3rlctwSyjY+49KVc7RLtQRUGZLe67GpiaYc1oClHYzV/dSQZxJS68F2L/woWdS
Q1z6bqJ85RHDRXtyQb+yew0MUmYRExRmEdv0vXoq3LamKV2jaTw8hV9NLkvXuER4GL/Ao4iTqPzj
D7s2n6W9JO/MiC1Q0pr2oarj+YWC/CQJuiTZvGbqKyTpNX4AQb9coecP+yJKJ4XTi+zHx0ScWzTR
SqQZQUd0JLEXCwzjWcpLZPZAYplgBd8Ier6lgEcwFdCfXW2aFyU0/7esNQfMfJy68x9wzdItN6cK
QYqhpGKCNWGAtzKWN4PnMk62TDle6OO7DuqHA8628GGTTw5pCuDi5wRBwjiw4DzoTVXhPl6y2NRb
yl0ngF/i4Zl1MpCbm2H8sDXs3inxJVTUpOvdfwcthU3xbfEqeCNHT5ship1kPWFl0IbH3psZfKvR
ZSXYK5SSJPjfCunhF4i10tLTBO++Vk41dfYXNpk8gApEXLtecnzdWfhuGt/5FF6/i1KVWxuE7efT
HGUwGAOGKTO5XQ6YvyBAZMXhqPRrMc+F9FRY54NpjQkXXapLEsNi8WfjpcLujWAdC1nQn/s14q0C
Sjm8MxC7E8iVTer1DZqVFBJM3YPGjGBGJMdmI7nB1YAqgL4eIwS2XjFg5mUld4+7hS6iycXv08tS
o65rVLCEX3BgKCKGRzy6gaX2o/13NFOxqgPyuATX/4snu9rN4a4TlNogJMlMu1HXMSvYIq+FMta4
dPiZmLoDTGUsDlqsfTrxY1FfXKm72WCwBPpZDs2X1X8sUutct0wJUu2WLWvRXkxA/BHEvZWqqSl7
h4wF8JR1lUgTYVrQqwt3U0jgEOSL5l5rirU+POv+L3lBDL6uw+3lxXXkOGbDS/pyLa48e7/nf8LV
Nqw57lZ1CDH1d7UwPx9qTV1QXti0f4N8N2xrc66naMaFhNYQY3q03rKTqIHp4SpzrMK0aC+rRZSR
Y8gD4eRYP785G9AhA2atMkYzYaNPCUzYEDH83cmUgwTNMPNBI+f5glM4b1q833q8Y4FhLVY7BTUk
gjJx/CHWd0WgTxp5Ior6a3ekpgmdAoHx0QRha8wtrR1i/09xejWAgYtegZ8PaGa6uTmKLM6niUuN
gwMWNRZ8yAlt0cipnnuVPf46LSm/dij76nfDLFJNzlT2ubEbAQdQEUwrVfQ4rk4Be7Z/fqSKAkt/
1frMgUSHxCLtuUV249ox9eqhtRYOO8OVrRT1fdx1wqDkuFEkfE9ahyiC7DluVvWydntJPehawsYH
qd3jKXyt3w6sP9x+YwDJ/LjZGW9wkDCRN3FGMG08uQ8MvN0H7WgHiOaB3Klhnx5dQy5LGVRxtMBC
OrD1L1VEMawYM3vca3wbfcSfTIIMIMGyyPtd0f0tABiUOkJkKFlg9lTZsjYzjxudXs/8pFe3SHEj
s+K9hqLsNek6YQlP5kfxPfvxgZfd81VqZ7xiPg8JxDkKc5J0DwHikWEaUnH3RmzMcQq9EpQYwLkz
B7yBUIhpIMXmuXIVnP2nNRXp6nF1gAFw9IhjlTuvl0TERGXq3uhMGmK/1VyDu61oJdRYeDzR5JoI
AynnP5iAap09wHkzxAYRWk+PkfyD4+4GgvF/GMWdGHzOizirYDsMY6JkuECwSZKnx3efDRlC2F3O
898L9PQmKcmq0K2PeS5geK7z9FC487CpHnaGw7j8o3w27lWlSjcNmBrnz3QJY0J1NBlmQTnts8Cj
m23CO+UMV3T0AmW7CNGvXxjgYftLu+nM6LekxKuIfO5KjJlN4CrkYyxtSCJZY5B1xY+tGcL73q+G
1zGyrdunbxB702FMxeuoWOCAtHDO1auqbf6xu1bzLOaI1NwJhPbwCmOa+n9nz3JUlKvETbwny/Wh
YmVIHNgjdA61ai0V3ojXZLZDH/87PqDPESLhNZFzygJM1s90Banca35aAGkVp3MmvPl0CaS9F6pI
dFXaWPQTCyL8eT76LgBYt37LhfSdKom5eD5lHutpgeShjj+SSB1l4Pdqie9ULT/y0Rk2MAahLQLQ
VLRQFgoO7+yXa3Sd7lC5a3FUrMRTj3VQlbwLFNPUuwrlD/S73FolMzVO8YWKolEpAlhuaaRrijW/
oMj6SfX4bSnPLYG24Cl3Acwe6OetpZ/qKzWTE+qGnDnBdh9XsWTPwhZNf/hdB0uSFMe/hMOZ1jAD
9yg+HfPUepeo06+Uy4CQwXcwjjpv+dcu6/rk/sLPrs+6BOwSbhoMy0W4AWBs8qs2FeWlNLT2YhUW
imQLzcXIz24YuZ3LngBhtMVvxkWjBP06aZtMdt+ljKF4XmNg0gxBCZDjAohHCsywqvuUa0Yl3USC
RfG6dXy7BSgXhrRLhTPgoJBsSOJwMH8nQh/pECwBDah//dewmiyZv6jrphvM6b59HhzB/KabZS/V
H9l6qUam7qKalyzYr4MnWc7hzIyhL6OJYA8bD1Qg9awnxgAAiZwtjgn84Clp8h7Qe3vjVYuAlwNu
4IH/uM4rzevAbDgikL942b65g7TBAOuJMOt5YeU7NwGsxvXsZHBfvHTNwp3va+M2VbnTcufpNpSw
cCi/GwVnipttxt+2ZAoWrOhfjWnUyIfejbFEi/IiVnJaVJ9DefzHUoFF1u1RO5vMjIMgEw1IzSLN
dySlcmswZIG/bQAP8cmRuUagzKl/RKZaG+cOdFJJ2YG5ja7yB6W90ME+1sQbpmsribRPSjkuzFLb
UOibffNTASl/IOyUEJmp/G+XiUyGd0yHaLr9YvG52g5qiXdimrfOqiVYijX2OAIAvsguB69g/5ji
OXqBGJjP+mNJn39InNlPCtAGeZ75NpZ2vyITuL2gv/H94erl/O8Rl4bNd8BUcZrPpVQjItUKQz9h
WLnTdBGJnL32UFpapgBM5gn8jJyPTeY+7UZlgT3TjjfE3xv8n5Hcjs1+hhYx6MrJ+ZIdutfVc6j6
WrJM7cO7SqXjxE4+1/tU8srlQehclSuFYEwOG3646pJOkPWXV0eFYTPNEkD8IqBRAsMJxvUIbTCW
NvG8XhYAc+HgCFnAQo8rNzPTtZi16k21jke2UUk2YzwngdCVztexNWCtovnjTTPirzS06Vrurrtu
5mKy9qGh0YKlgOfKWI8vFKNI2x9c9X9XEUmAnhXf5sSa+OWG+PYQmNbrQHJfzea2KgIg5fwKfAbA
YqvuYgaF5oO1sR/E4tXAT0+yTVhuHa4HSx5QewFbt7iSRugF4S6MB3fll2eG69x2/8HwoJDkxl67
SJ3XJcBK7M3nZXNxhGzJNT/Nrsx58BVH4ZiE1Iz15+Y/bML0DuU1EsaweRbli+gTyq25qkjMY9WV
9636BcJuLKq+hCupQnPEqaTBsHhl4PoEyS4csKY592hELrvS+GMvHGCCVdl7ZOMksX8+rxYIMRE2
9ERnRmxUqzXCQeS4x5Pdty0TDSg9k05zj0HDLk1cg+cIkirN/jcTEZl3msq9+CyFYHpuKVWQ3IJC
SAkkpA8EQ6QIzgS7tQw8AWEkhTIdFs4At2aLgtZl2Tf4fsB/sTjDO/H+2H0WWWyF6T/TSBOnZuxx
V9Uzpxrw1q1+y28HX8bMMmfB7mdmKNymchhRYnsNAhO1JmuyowEFwqhs1lUL6XdK0x72rUHf9kUf
dxlX1h89INnXLYTwogwRYMQpW87sNo5rBAOZCrqnPEgJS9PIP6q3G9jPlPH4DDC4K5GwwOOQK3ib
BR4SvG9m/DMAOTvKLsws+jLb8xWM0wv/pPb7w8xYuTVJP0cFnT0Hn38VSI6PR4pGpvbZ9yfxojId
9rFqkQOLRD3Vgk/pbdps6OC5TPPxNpvvTFoNIkgDF6PLHT8ptJydDfgVBGrdXSYg4727lgcPObTY
IsXfgcm7emJntIbGwcRRaZV4HD3EPJpDqisXc1pa+19zfpdgZ3U1XDrdIknz52ojTtaa+VTzfwaY
Of7eCrayHqZQmqjo1WGABys8ii3i1UrX1GZdRLmnS8n74+dtZXBUHvJhir2/qhNbrmgEC6ngKE5q
mk+0tLdrzJmlDoOo8LyPDndiCuLmvtyYdQ9LSMNvUSR4AZ9sKHmUyMVD9a+uwTo+VuDzCyhIRpUa
oPMOFgIWLTRKCld/ZN3IRcHzNZ0gS2vVGMR4Dj2fmBkj2/lLaetiNtKAnMlK13p9ZsHkeQ7BBg80
2UjFOQiu8qGCYp9LuuGBjkqT3/DMa/smb9sFw7rtHcUHxMj6qcCK3Xx3i//dieLQAXdN9AJ2QOeQ
6dyIUfW1spd/wf59LEoUOgajNnRIrbBOFNPsVdUHZRsGs0utTaRfZ3SREtDKjhcXAns3df2LbOX5
4LaMMzvw6ILRMa2xX5aA09X4rB75O5aBvNrwHLdAnSAWsL43ztbzrr9+rFbBExxwLbBLz2QWkRZ/
3pWkP8x5GGfqRJeHhKFHlasKNDt/sC5kctpE6odQyWCYoaZEvC0PpBEL6NP4yDh7eX3vPRFAze/m
ajYersEbkCGwZL3Iwh4sqwSDWki1Ct9gHVII4aZ8oMX1Hbk9+9BJLayi5vdsAjzLkyhAZAwKmoas
4kotUVgrYNouaGui0neERUnJOYVkRuBPC1o48/VwsPoprRxjRe75RthPP7DvavnfTkPK0ASCGB0v
ixYfhLKtCg+hh07Gx3waUZBHaJGFDlrEWgmS3C/cjH4csLD6l5NSZr/qSYkeDR/RcV8V6B0qyd7d
l0edR3toqjT7rGpa3K/XVGyaBK51Z303IArHXu58GKY30Xonx6mMSJSbNXRtkOt3YYBdrejaJ+8V
gF8mwo+jLZTt3BiLWMEkyqz/QyBXpMggUySFp14qFmL6Dx6At6FEnDZDbE6H7crahrtGreEPxUHc
3Ttv20eX4vs1OXjnPIUevPN83ymF0xphHOk4YD0dD3Ztd8rXptbUuLblPFyZ6M7Vd3r2JdZPJeVf
yD4byQb4P1dfioUpWxJLVd9ctnWO6C7rUuKS7nTmoETchflYCWTbCOqBxobGCGEsX5tE2rXWECug
HDhX8tBhNHUZLFEZZaYWPRyNR7BVWHOyaWeqML5scO8dQOpBY6CJzchLsDps9RVG3hdrae8AA7RP
BJvQ6fCGWYRM0r7u0MRVkNC6lBxARqM/n8xeOB4Y2I5dz4wP5cwL1gHM7LUIKbU7i/0bPMDw8TAW
GDz11tuF1KbLNLPwqXmpoe9pQP1PjNfSLKSiI9UC7KUpSI2Sy2YkKkFBROiXMTrlabfgCwAeYkBV
PCbPNHCCX1rNNlZXm6J5nDN+k8/EdVwpD1sGwtcKgxOnwkXLa6bdyxL5P2CXrSZaENw3KLVmeC5b
eyOeJfQ395WkDA6vKYnn6ecUe7hEnTZ36ygx4BfaRrHBNS+jDqf2MKFbtaIs0MfNZBJdzF8SEBrV
awW2VXFPQ2CatJUE50rZNBfOg0MTl6Bm8EbTtmbrMgDG3g5+j1rtP+ULN794gIY6OX31OZeg8/xL
fiu7RngWz8UaXpy6TzJBxXlo2NlX2BigvML1kqgAtwsux3dIQx596Fxa2fGOFhjrpryoIj30dBeS
c4qGIE5HrqYhXdybmKSHP8Ek1U5Qi4rin5/EVadxQuJyrgH8hnMUegyfE0JTm2ErscYBtoKi+mpH
nWBenYwSvNlhFfLL525BNvpHpCsenTPNI0zjjkSIrwpc44gT26qsDXluF43rs060lZ3CxnF1komH
Ua4JkvmeXk4qocPV9FLwFwlqmLbS5xW4K3aaZDLqVMdtuH6sZTVhoDfMKS+jtlzCp5lZW/qqvve+
nTEpmgS3xcxX7cpOxxwt2jbdOCjrEDVkTm2Fc/8D6giaJIDnQd1z+MS+GvR5ZNYo/J0WNpgTHmil
yOjff/OXTnX/SNeCRGg/QvN8fTVJnBWjjVeFBr4M0/iTFizrDCqziRn94F2IRkXpUL1M+UDtjFrQ
82k8jAZprfFeR9+22SzpRKWtSWju+M4RJehMd3GElFyw9bfPLqFvQXE7F013BgXL2MJ1i4PE7npA
k3UjnU3BNAdTyepytZE1qnPGp3Lmal5/mCf/xrLYPQ8YWDfb2sTHgNPNFynG3y44XJvl+E+7a/Q8
BKKTiOml3hyxwnmaqrb0tq7kM1MqOySlB4i+D94BEJ4cILwcaKPFkzun/ms6mC7Wt7GysMg/nnbF
A3I5MVvoQBro5GQFX+geBdTSbo/ms6vRIcp8gF372GeqRH7NowpTkEmkzRxvE1S4pdATTKUpOlPo
W77IjPYyTFvdlq6/n0oICbohEA5+CHuHB3Uc1lqJ7jGX5ghQUJrQliW/7Y4wbc7lhU13/CyEbCz4
8tafzeAlZTzdPVQOmWcMEx+9Jbe4ocniDKRxUF0QvrATqBbzsH7Me24bPAGP7+wdsc8b0OVFF28q
/q9nX5AL9XWPIrw5qJXsltsbvvbHp7h6lXJyS3tSbbomcdTh3AuS2yvwK+2OPEmC8tATDYtBEQrT
Bw/z9dtWjVuPjzEREwj0+Tj4XPfR3DT8Jbu8IjdinlbS02rh1/fAlDTlcku2bF/7D39EA3E2Nd15
fbGkkxRLMftajGy2ha8MS2eo2V7ye5aYHUiIDzz9gYLU6crIcBshig1GZQwLqLEaXmEtrvBXAs3L
LEKSymouiAgIWh9JbdO4xQGFUtz7SEK8BSVzrZjztg6R2HxdgZk+FdEBj53bfGpK5H/Thesd4QQ4
mHyfnqSqs/NhgLd8JIDnbk16PXE6XbGFRPSmkcUhFsIYzZdfYcn2W8WHEnhkqUnnZmBDcNZzJlLy
ybr9BwcsYcYeDwzKfP7W0cHbvdmmBiqcFXFl0yR1vxJ6jP/twz/PYQc8mpn4/UnXoDtY7yPavaxB
LemtV68kn2R9SAiDTp17i6S6MuSVk6g5xr6U9JpMu2gpQUFwZfBeEhO4M6M3TXHxvkX8SahLZLSB
CY5T8Z6+RUaHFSWPCqcxxArpj1fkS02vyL2yD5Nkj0HNLOB7RJBUSE4dVMUxsgZF1cNPBDE283mJ
8D68LFCyqJL7GHKQweN1RqB8LNujeMqS/CtTDuWr6gXbPeHRZUxqb5jn8mnHGRZbrxWI43A7eqYK
Q4gML5U0b/gqD8j5d6bAsA+HkgceuFyGGaqqJYNT0PNKvpl/RACekNIPGCzyrc+buG9m25nqLo5/
zLStG6Mrqh6sQ+BJCzVVEXOm/9xxolDAv3/EJNQT/vvRA517emRlocuA5mYKxcf6+q1606AKbLWy
47IkkAuXIqP+7sDGWcoE+Dz1vrKNeaWzlUZiYPk/ithRFg3sKwppXX7T7pOBU0wMWUMInhUO9ucu
E64as9IWl0eoYrj+dYQ7fnRKtaIHex8LWfrddDUX51qHMjTedDGaoFTaAx9qu0tMqjl5TsRVdtx6
nY8TtS/fFe2NGgwqHal43tTnNW8UuVs0usVlX4JCupE0xzju5w0O3iNHNNuYeQd1pk2zVgJ33Ggl
9HU/f8krxm4fme24UddSJ0AmKb26zj7KczdxsECKYPWKobg1IBisgSRrb4JZwEab97EK2yjU1u8D
Y6LFrBhV18pjGx5H235hXbOQ56Jt98USysposLFbbrTjrYpDElpudzYpZ8ng1zdXNGVv1o5qh1l5
7Pr8fqH6I/Tt9zyGtna5lVsrYztJrhgRGDEQ5A4Vhu0Uu8dx2sTlFodS2R2JUhkeHWUikpB0Ywve
jLA+F5bd6zCQYWHtSYKTl3zIcYWMTZz3xkPjv5nOavdhKHt7++tMlu+bNBLjQIFtHovW9KlLmv7V
QZHtjuI1Lnm2ljqeSd2tT6DkEu1C38U8fwK9e7aoIN4nwsXwO0NXSBSReJqvlCl5eJJDwsBjeA+c
pEXqAlCIgkg/iuvuUwMUHM3UKGEN9ZcDj/fkWHz6VmAwvgi54RYlmnuAGRqf6Z7HHSENRXdzbdhX
YGX2i+vnzwYcBzfG0PwLcBvEpCrwf7jPMA8OkMe2VCrKxRRr7xCYtG4MSSVU6dbAWcvBYPjJQ3Xl
gUzzVMgdU9oRcEUD25r4fraLpOUfFTws1LPuCcXx+BzguzApc1Z8bYTkOGL88ULLRBjrgIt3RKXs
FcVyfmz4K0wZ2NDdWq8AJKTl5zFFNW/dqYcb1DfckepXSHP8J5uly672fhZtzkCZ4qdWPawM674J
d8Kf65rlkMEJFqol9UZ5iTZZgMcDdiLE+1M+0123H627w+I6T/smOvUGnr/CSM/5ZeoYlvXEAzaC
43wKWNvm6U/7tuSDwDdp9OB9/TgmzibTEC+DFBFkwJhcFbwAaIJEAZyWFmK43RIUx1HRYmjXTxNO
AQPOXbuowNAsuDS768VvOZES5Z0SX85oQNJef5zG+19bG7xd79EO1i5rNcXGcM9oId/3eo1kvLG/
qYjh63oBvRJNeYA4DOb9lXa6BhjrhQN/hJJ5uVVOFiazn+bR0lvuKhrqFASlr/+oToD/nqC7MS3W
rv3V0qiWbD7SH+ZpogcoCzh79sloEjz7d5lROqH12JAbBhr9WFHntq6YRR11MplGLiDGZrh0nVyN
JT+kofk+1Dl/TQr4Nq0C+CDJ4NDLER81zV3np0L4GR9s8wKYXErdjRgN7C+4RRHFiqjVsR61e5Pc
Sax9mSsrWHTumM6CRIs8R+I0JSahkZmp7ruAJJWZD5TzMqY72xrypzsO/R1cJqMBygX8EpjU5Lz+
9ooWrTi5R19/H0i/32ISopGumQKOFvw0jEJJ+gVdyHUTvOkyivUqtiDYvUvnlOxMDMaDyDuxJczv
pwhN7FKaQ72408V9/CVbjpFF0V3halVb+tD8xdGFIdYMG91C0E4h9o0OnXhJX5ysDlr5XEA0DwFa
OD1tfUvxDa9fMMlUe4E73DYey/IgzNj6yy2A+bpaQXrlpW1FbDsA5G4jD6tHOMjv6hf9JBsXtQe0
tZatGMvJYNRuG8AMyUMWR1GNMXlDrT8vseShMrsr0KQcvhq+OMtc11QXBxFtceRFgc1uhBwJ8mk1
nVJPtSXu9RmTflX+kzN6k1ZomxG8I+J+ryFR7NUW/gu/Jgpp/3YJm3e1jz98dUOJYqio/yUL4+Ia
wgR/CMg7VKu/Bh/NZrcGxO71WeE35jEA7zP826URLtrOrtS7uT1f2AtGcAPR9brRpomSi9CbqwD6
qQksWkH3ziCpO7RebDnkY7Z46SRyuGdDm1f3g4/3TfqIgEAuah7XRMJ8ee2ZupS+apMFIk+dKnu5
Kkkyd+0YFxxobuHLEw/15rT4Mr3EBDB4xC3qXJcHST2SS7y83qn++fwBwOv4UUgduJVsF4pVSJ5B
mtD9pp45XPj+k/7QDUE3fit5O8EZPrxL7iLmjFmn7wRCX+ZzQpXqAxD7QyzV3qcKUn7Vcq8v5ukC
tJVbcoamlf0nI9kKVxszRUdyQ2B51EJM4t55IoJNl5LlUAplMoXN54XUc5IgbSasw4+H4x/E+1VR
uPjxxF+iTvxbdWXnQUU0av2A1seloUH3HPZRyupJwU1LItuhw2eMlIcFReb4+kmNMoh36e4NLjUE
4EUI9hWG0yO9g+ceHxhANQTqd+7OHVzdqXG+F4DY2JwT1rJj2Dk0LDb6Uc0cuBW82TTM60tSWfMK
mBXDriDPgcSe88Wc5/6Vr3WlWNOC6NMJo6B3cFcYqChViv1l/HDMmSJVqJhUMiICqJI7tgBJwKTv
LYyaGCLfZR9TQ3ZUFaG7A5DVeB/ju5/1WhNTUrZzrUsu3pQBRJpX6eKjtVqPbCebnh/JiN6Fc0CQ
th0jVPVW+Qbe8WjzxmzKsmrq0SakqjYCO6M5beUGi7kW0TNBq4PPk832VK1aQiVrgN5K2uC3XpAx
D+2Y/jlJVS1D1lDeWlA7woiLDpa+BEM9Ovv5SRh9LKn4DJTsOm8PG5wkkkyGGV7Vk/rJws7Mi/bv
QRpW2emN3Z+3BAq65Pk7iN+QfiZg3KH2r+99lUlbvMqfBMyxF28CaugoSRMbehE2fASq8kB0FonQ
d+lgU/PXqAYP5Ki4ALoAerkrQIR4JIioMb0CfX73CZ5t2eedZiUBist1CA0ATB97x1HBYDN3kX6v
CVk8CN8Af/Hxw0vq/klPJzL61WFcT536gk78T46yqoDtjEPgx+Ql7HgAwHDjwJcFUoFj1qBDHAGF
3ev0VW+wie4R1XawS3fD8Z+bR/+Bn0vBcxVgw1Kq9eqjtruxD4QxOWMlD3WYuIRhdL42CdD8u1Zb
qG/5Col2ETC8nnmcO+5t5JrfcoYORX1jAX27qyveo7nobHOdQk6C5718Z0fm3EQTh/nw7if8upWh
mq1Z9zWM65QCOAVgYGU21MQbM9uKlbWvSUcqS45jhAMvsjt6KfZejx5V4EwsQnqijoeYJexSDLhl
dwUSdb13pNdInJyDMkZkmQdGRaiAVINucT5xc08RveYlJ5EKkdiycfyEFRVdnP/A3JWOw4b+/tD5
ECodAzHOCFaxkPIBfj8dz3+B1FIhNAL5j7tG3bcM47n4lbGilEh1otbmcjJ4vKFtEJR9bIZ+9Fcy
5m9e960aRbnRG7bBnkdMXo4BHkooPpIonsNEoRTCloo7HisDyJ6FJYFfjz3V5piaEQVtB5QZnQRW
IhtGyNvNLbKR4LLFKmu6YIL1k6cVLUhUvGYksTpqMAv7rePLms6gD3GBm9gSfgKqPQH1eyIcxgnp
pUauk2X7jpMcLyrBRIq/7o5XHhTSDZFSJO3amn02BdCx3TJ5RKEYSsHQinF83p8bLDuotXG9qScb
9el5xf7Z7dEu/9VouliHKepibjInRFkYsTXThOYV1FT332Sv7lkrKNnAvS/udr76/Re16dgwv+N8
t8IquzpIIbPkBwqpYiCOhX4xSxA68LFjZttKa8hBnQs06ncHgttV2n04ckcUOlv566RIV4/GKBXH
d/CtcwWUus4yqJJf3VaRqWxaMmKhPoHAcRPvKq74XEoaQE+ZS5vOtU6BrR3ASkdjHpYOwrta0YrF
B9rE7vKqK2cHUqqDESic8flWgrrF68IXWZAYEh8FSZOJTILABqSuZCX1/KrK2PwhPy/DO0ud92ZU
U0NjdmEiHFCT69o7dD7Lggw9RoU56TAFYjS9AUud/CIuSgFw8qZN4y96WTYDq4fJ8pEAFO2XcxBG
dkB67IxJz6IEyXbQ+1Jb/tn2VbFL7cEm92/3+lC7ssme6CFMjiyAL+opE/hGfJyyxws8Q6GjYdnw
xbdEyTb7xeN1UMvaTl5ftFzEVtxGZhkoJGRUOBcm9kXva57WaT42ufyQtGKr9cqBucbZnp+acPEg
TsxLZ+uav1rsqJP3rNc7t4Isjh9UtJAe2sT34amrPllothzoP+BPk4OaV2oeUlQoCo5ocZNHTv5p
qcBirmFz8izsDKRpwx9Ir9fipZvVPn2lZvlwQUQynFLAknHc7Yc7/r/hlgw3u+0GoQRKHpycxATP
Kn9jf/y8KUdJ3wAB0L0PbSu+4C796WDZ9/I2zh4ETg8N4XpYuioi2lRooEF9iORqFuWXZy8ej5ib
82QM/xoOUEbqwtx5l8WHVn7XWejDGEAQFP+Tq5cBupYR8rjkU+Wzrm/fBF/mp9ZGDARwlHlghiNo
PQERAkfP/IRgh5w54JeKklDr19pYXU3/ag==
`protect end_protected
