`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
bkKDCdGzTWVi1ghehKQAa5goG73GCheoxx7hLf7Egu+EfAVEUigMhuC/lOZDTmWB/2UZ8mz0PmAR
vaGnAQwCOrHwo7Go4E5Mw7grUYt53O30to4ZI/FM5wy2Qq2KP4JFYIkDFBlLpI6coKxbM+LqV2d3
pGcXe0iJHRUqBD4qfr28Z0GztBrscr4GLs4G6HTJ3S5uO6to6abXrTYsaNrl0PWXRVD9lNtcxl3o
1sINBoeDiGA0gbbUB7XxkZ4QMHFugh3NFHce1UHmv7dGzlOgrTut9OvOkaYEhE142vVlKOz+ToZZ
zDfH/R8dNl98ti2h/u/gqMGp5nBV2t9hxr4wkw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="PPfQoYgw4PYNaCjZ4vZWJNa5nsG8IiWXaf0d80NBX3w="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 104496)
`protect data_block
hVpjpr/oCl8NFS0sR5X9A6J+vXE3XLBEV+aegSWbAAbqKu+Be4ugwR7Xzt+7M7zCa1OwG1DIAqEY
aerQjBbnScwsK/ywRf0FTVWjGQRG4Xxcif4dFoGAvu5Z03/02rfvUG10osw7GgUiK44KL2oGP7yt
lGX3IB0Gilzs7aOpzh15bKCCEB5x7KRPUi8WmXn1kHy2h+gdRMXmBHpj7QswVR15NkzoawpcVh/W
sr8k8lqr1tcAA3prrvr7YVU1JjwfsUXvnzqMGjtQmVrDeuQKjWIo1aFrNndoj4j22bNql9fh2ojD
/4NuXKbO3YdIeTwi5HjX+D7ThVW4Ajs9re0swln4Ddvl5WPNkaxAZ5BZe2Rx/5lk/Nn/WsOJF2CO
b0SsGq1sJYU7cFxDwMu4dxFs10DmMnjm2YCAr0qaWpPKRY/zQu+6cstqekDXJLVNKAlH0bKOHzfw
MrpdwA7Orjbb+hEQWC2B16ixVn+dkM8b+1/b2ayJcU544MkjLaRY3V12EwwVq3G1ZHOsBz9j162O
GrdQg/iIm8Omf7Bw62XVtEn7FZjxjqxdsj0RFRR/D/KWQAG8uGcqOcz3SDYFFXWu4a2nMx0T8GTY
BU/vUfn5/pENyoJOYry11fG/dmVbdi85hL2BasvofwvyTy69ADpvh4JrjPYhQ+wlZv4kRk9PMg8X
39rAV1PXoFLEFpPfKEqTeidXYEazklgTUtOi2QDqiR8abzWIAgEoaG5DSmuQGIIUhQDLeEN/8gHa
0JyWsxfGON5MJCL+aS6NFm5BkolBJeIJ0RLOTcMTT9APw6mTdfxVLnjVB4YgLdugFe9Z4rqim32M
OGBLg8dZbILqr3M1eK52EgISsyMir+y1d4AuG0SukdusfYA6+qzzZSw+Kka0iEiGhGd2BngpMhIa
dfJCqi6uSENoeLxKc/XCcZ/92l0zQgcA1qHpn5eDMPW4I+7SVX/zY/pSheBFISu6bHDi2Tmuhbj7
pLIpFNhA19YoK+fG0KXT4DetVu2eNx03ge5CanZ0A0LSoFJdk9ARTDNuwTvoNYC+xCwvOntGsm+r
k4/nQT8MNWnS2WY3K7IJH6HEaMf0Y398tpC2IRG2xoz+8dr7cz5vnim6xKpcXeNrcP2oPlxb1lvc
vWlkophOy+SBbbU1gdtztWchcVUaBtIeSGupEosHplLKRAD/CVRDjog9rkl6m/Y2Foiz/UHRQhVC
RFavlR+18N6lKwUbBiFvSCGyHcag8GCi4W/qO6pWc+lgvYPkpxeGQIkHMU6YnF0R3sVfFBz+nfzm
5lngAkLOxxcbksjGeMMH/u1OV8WG1odENb+onulIH5SErullednL2EKDrvtffygOH3BOWGr8cF0Q
Six5SSysfCtTiUX1TI3qTY1Cb9WJGKRYtKAqIw7UROF0HzDmkPUvFKUS2hd6vmwbUAw0SD8DYRno
hWU6I9Esw0KasOdX/43tCFMosVzYQPcsG+1T3xHq4dnoWita5RoPdP0M/NnEYW5u+Zgi9Mi1Kgjg
KfI1ovv2xX1cCcN6dMc5Y1J+BB9kgGziPAuC23Ldo9OKGT6347Khg8c22Qqownj8oeIHtr9Rbzm0
pO6x+//bEvSY6rZ5cZZ9RCtLP544XzWHkf2LI1GJKxP9RkfQLVWUq2nb3u0fZRE2R0LlAz5yLMSV
WjJl2H4hGN/bGx+Mrgh0K42ohEOYvQSwsirxirKHy/WBFCE0lRoo1hO5/Ckv4QqyxaX+G+PLoRc9
bMjC1MWsnZTopoax/soYo9GSGc+hZ7mLAzC+4U115gE9SxYkTnzlWaljq7ktk97AWxv3RJrADhWx
JAvhipS+FHaazQ6WMkxwkft54Y8TaWH6eweawIG54Zf4X4vF60ElDoI9ADxO4U3f3qcjNCEp9QHe
4DLFq6kk9+PluOImgHg+nGt9KWOaomTWMMqNqwxaByl0xQYDFCfO9p9ais3ToMWpnWIw812NwsIO
8+06leZSyr7nmm1nv4i06aLNVswR0+I3gLGhuFj6//y5xPVy9A7CW5Gvu9mhchUtfuzdfOUsK27E
WyKKck0dwliSEyZO3O/mpS19t+NaaWparqrBwM87EzSY0aWyzQT13vbwHNH3Hwqb/Pp53SD8Gn0h
O0rbwdI9o4837JPWaWjGxCvrK29fzdyVEqJWZvrs63NmKhoMcb8V8jaVmW7aKZMkh/M354ljI5bD
vyykZF2rPiuMzOdTIO9K4Zie5vOHAfNvoApZ91xRyAIk+jWzWRKsoH6Ig8Rjzbkb/zbrX16jP65A
8y0za5FfMptqcNA66YjoTcqT+qIIL+qx07aXCro9+CFpw+wuYSgw9EuwD8G/COEMf2K+HTQWbFmk
BaVMbA81yEbz0uzz2nU+JrIVWUn5XzxIbFC5HARr6mCMfikwo3IZvqG+mJyfRbQiq+/kjEZ/bEk5
JdkeQFb4L7aKwxJQgNhpanEQDspV9J9JJwD/ykPOEashbnh5ekBh4Dpzz403iGgI1iYtbu7TX2dR
H7qI4PxJky5tbBhrgKJwLAZuBOLiLupJgskQLDKwewwCmijtq31jYn/Ds39u1y/rRVuS5qPOWbMk
Zyl0O/VywI+8p14pIiz8rHf66kxLS2KtdT6V8m4r4hJ7NUsOO6jjxqZo/9P2S7XfaucL3APCVLcE
GBa3FHYhlUGbX9r/VNxmsr3qrGYso4HUAvQon7fpAe2bv4Ro3/yaGUdLJ+2TRpBLwQ9ZKpxoVjcp
z/0B6kxqT297mW73MQupq0DhSk+pM9znzHvt5LVLFh0nNCM608h7OEYBPXpIoxgm78lqLbQowC85
hzLfMzjioul7RY6v1AhBY7JGvQsEFRPuL5Tt5GUGnDPckKstK+jp3E9h5Sldt1G6UP1HsHeza1og
N/SA4jvFM42vbQvgy1VrV3GoXCGKJlvYSHA1EkljwM0VvBCjf2RNCz/a731qqM6QE+mqa4P3edcX
ivVBztye//lwmpjfMCc47mKvru0w1NlrBKA63rpsDDV5rhYXcX5/w+ZYhPFT9cCtP5pYH8AK9TyE
YiYHuv+g29SyRr0p3ZjECb2rl8Q905PX3wDlQbs2rKdqPlO0rmGaTBWGLxCRSfqvrkkXXO0cm+yn
hWzabz7q9PR3JRQK7+Lihq1yOAbnYaCVGclH8ucp5pvgAGo42ZR8F2Bu3NjFjA+K98VuUEQRllMP
8hxohxtttOQjmfXJgzVgHp9JvfcwRRMs6qKvaQpKzsGC/gzS3T87YC3pLd714znHy0pKe7P4iW0N
PViCzF77A/a+5KnLfblulBhPEvBnyhm00PzAtb4y3xmh/wcn2YZdwlAsvZobVgCAQpokfv49G7VZ
DBWBl65lelZ6KReAPkuITGzJFATnaGMWGyX410COqsEW1C3XAMlquGggC0Pl5FNFHe/LtGlHh+Pv
NPV50nzli2NwuWA4uitEs+MJWKV8xSLEGEEPLsE18SMHWIczCfZ8l94z8L1FLsKk2y4Avr1ADXCA
8R5wqgtFOEDPIyznuTJVNAz24e7bwSEimC1sAn+eVK0Xpe8BAYK9Kyc+P7BJ4M5Ish+N9GM1bw1y
72EXoKX2D80nOc7eAx09pUw/UC04Nh6KpMSpbEXhb3GqBO4enH7auvljFCOinsUTv2I6gFELHyZP
cEU6Jp1dhWLgB59Cg2ppwmCatVGVckTFtauuA85JD0zq5j990uAKUDCcDnTHbEEmF7dNMcaNqfxy
UAxq6svGLWaEL7Q8eAmNGAbq/FbolLAIQkzNG+vSYcdfWTFR+g9cBFeNR5jwpIU3XWCS/inEiKx/
mn4oG5jpcRNfPoMZ4/UbYntGIZAScFm0GTirbwBmIO+O8JqF2pobxZ2CV1oPpuILx5H4Mc6EjiaH
tu99un6gglrhWu4IUAGXp1qo3WkqQwyOS+2BoKaYz8OkrzhYPDTin3+r7YU0JmY+GOjeLftqCCTq
eue/KHlDh73WTXimuULGilCwJoCxMgoSWvmrqEAdRrqCNaYCFcfBUq5pzEnF1K9OBhAkE9bEoff1
VPCwB6DrA96HyWuCJmTHRifu8bRrvupUXyTtouhQy9/M/zr1BpYH4xVmSUw5W9Aa3TgheUffdsGN
YETwWAmDk0wk/ZR95PIG69MuHVoN5O1X4o3PlF+6E2uIAtCsMoaTPLYeO+2rTbehNuR7ty+KLpFL
zXZIh+noOKzDRn/i4os5kpsGYSkrRxksaGdsTSGY/D1vaq/eKLdsEgjODen9xdX0rdqYySEfdsm+
jF4Olx9/VO3oPAMVSKs9D55hdmoPxqRlA5SlA101PwPa2Hdj8heq9UNvGpRD/ukzJccNmLbBa72d
IYAQGQpSb/IAqcpJW3Wcr4Z5paupnyrtC7g152jjz8daQ9OrNqEwB+4426PZ/eUgRZVdb9KuNybQ
D4FdC0394k8XsK2+G/Gcua1e358xFnl4kXkxdvQ64XhPpJKSHCF020WS3VJQTTRXvD4bTQ3DOzAc
ueyNQLBTBXKjxEerB+m2HXlcUnjuzauFherFT5xINxBad0a2aMrEoA/7dOCFrtSZ5DHPugTveTMD
Hh2YG59bP+6Lj8oI/KtWhY18yqAjtLNd5rVNQ5+Yju83Y1+Dd42YOv5URbgZV036GVrA3M9wnDD6
FPNRuJwhCr5IP/0+5vjdaSwt82uHOdrSdGFKclLZ0kGhr+ecG3rVwJYHZV8ipdjLXZQ8HhWWiBi+
F/ovggkMvmHLb5pWObduehDbXH/yhRTGHf3YoEJHj07toouj0bWv3j+Xv2czjE5DYH8LXSQaoO+d
v+dacSCRpncebNtRn7FuPmSzxSLMmepbFYPK0JevrzlOhEDPbLllV2LYM3VafKzI/rNjwfbN+xmK
o9vIqIcdlPztsZKs5rPKy1vIGaytKAFaOOVB+EDYlMsWNqEro/GJLVakIK1lRaKypasCyPhNHQqU
fDCCCijgPqbnRg3zNpEhMt7H9fq4KHEIWin1k0G/CHCJC0WaTqbKe5Yu0HTdgPFcf6/txg32TITN
tk2yhE4I/Ao14JD6pZ9zZfpU4NRxpscVx0k+EEHpYyb8aaw6suC+1HCKrpKBeyH5ZJ3FE88GtYWB
6sf/AcP/rkGneckqw1NtAfBeeRUrcVX+0eZo1fztAjDLacxFr2EdMhcrbfrOuiCjTcWT9+np+do/
Ozq8C226G3YMj+Q+nyJFklpn/+VCZU3K8RaDFa6d1s/IqtCbKz5ao6tEEqiI1gvGhLlut6jwUMKl
DyiL+fedopp3kZfrF90U1GHq+E5y0GPNx9SQolwrqKt+wdsIppG1L1yoLfnucdrxAmbfbIaZoiyt
h2ttSnkgeTh4ZRmmQQpvNGu2f3JW0BeAOB5TMnHGwOnB+xoFODEoAdFu+T6Mw80ZnS42NoYigSC4
yfCu0fxBEUe8EhLtNtg8B7Otkpx95RCHepfG4jInkEDfbr8mamlF0ISJfKXXtfKPq9Zwt74T8ZAx
oAWNvWHS51tzjDpfAtTgD/JZQvI1vMAii0WHZWsYjM/18H/kVVvIY0+s9Mwby80b9klJolRY85kd
8rgG4IdJAqHVPIq+LOJmgO70seg7xdrJgT6eesGqZuSrawWlP2Nlg4Fn556QX49wma5NXGsIN+0k
1/AZyEyVSpw+hY+bmikqozNQWSI2wXQ7A80KVqF8CS44XDCwaS3TJ+SVkHyB3GQRnalCKPweuNvf
K7tLX6kIj9uVmlJq4OZegQGkWnuK8+LqBYNpAqhTNyLi4DqIjvx3ckcJJnezwvhvqnB4eagfjHJx
j0rxh8Qk7DU7/LxmcpUisPZBRDC9Bm8uBkT/fLV8tXZmOqkb5MgvrEZkFGqMFwRqK00Cjl3NA7IG
YEMvg/8M9TtNGLd9BM4OJFEpiYN/q3MJGXOD3hP4opBHODsNEwIgEJg4CChaII5Y7ZiztBOQTAyk
gPvN9Nwglno8hsiQdbAXAw0SwNV2gtyaNo8QlPaLXqo5DtUM0j7JVdYsRaVsHLW1WVBTgHODB+WF
AtJWicc2ceX5JGUN7P5tO18Km4ZY0/Bz9LaqsXFo3HxxQy8vWLZmTyhmcqkE+xOFGw57ZU0CXawJ
4GrvQ9ehR0ZJQMcRO8gePGgZ8YoAskgwvt/Ut59NpckSfGEQP6UajmiKIFxDkCOYO+y+4pn6D4/v
UVgrsw7d5qNwN/K7jn1IbTy3Hq0LgcIk77OYBMLtpagbcqhGC96Bl6cPcB5zeQYKOWwCSofz1hJj
/IXwZPKmaEjWgDp8Bq7cFuqFbr3FlbfCXRN8TbpngAoseQad79T7pZ29p5DVva1GZDssofSWopEu
itJp9HU4rCqMacNjPnQ/ZdmtC+TxiQKfh1B4fMoI3kcPWMkQI7cX2/SM0dKspBmDYRDA8xOuiDOf
fu4RVZliiLRjRHrs3qBm/xpAHresaYNEhCh/NustLpM48T6mwPTzeLYQqYNHpDVxyGQ2PMBAbrWx
Qrn/C+GY2TqV0gQ+pJjt29zwPz8ejckbYTp5KfbIrytGTDipYJdybUKvXG9u5gHAH3vcFuHo1dJ/
cmypZwUn2UAfW5M8G0Rms5/CRPc+u5Mfw7Xh1vTEooZj9xel4DKxh4LLAxOd7SuyMOSGMoRA4GgB
hVC/Gv+bpEzBFFIqwrIbCjZA4uT3RIpoerDQBeSuSZClYCpZRD/krLDH4rdL6Ua6t+gPJ9jUxIfD
sjzLdhxo+DPQfllXEP7Zi58tqz6bv5I/7K5n4cbMwpezdutpUWJaRO6BiAb0KeYOE+e2J6iYxtN2
hnz9YuprUmLRQB2dSZPOp5XN/Jn/IqP86q/hWMrUnKvlc4sp9zdFX1iD2Yp0+HFpqPdpwSTCahyP
GQhXtoQrcYTPA0RnWE9vsZzcF5iN+yCUrl9VOLpATc9e/TalZYeu5mthigudJeTPBmC/gNIiTu5o
OIu19xAbT20Q8qW+OvJvSKp9Z+eeSuQUWD0l6VubJ+aN7T4sVL8fW0G+0Fl7gj/f8AhovRZ6sFFu
0e/HhNQrCH4dDE8f4XKNR7hZRGpfebxjIHHSlZz2B8wilegi92in+lpHOfE3HQBCwEuomXC4t7Rj
+2zjQEmybzi3Ffx68a9uG4X+YxJLVTj5CpGQqQeX5oafqDEKvNphK1SIJiTBI09YuHgJphy+Tabp
jsUb0N3PvOuqetKIzL6sFm08vfo6btfW3slTjFq5FIt96Qcoikpc19TLok4CDNe9YIlle7s6QNqD
2uuxJvSLggSgC2vyeUGpykiMIAFJhGiNwYuOcz74EE9vHl24ocsx/xEnKV7klcQW1l51MSZYctnN
0XnJjcCfDaUVlAERTFzWk2Yiq8Ua81TjzUiPv7Ujx1c2oM6mIiqOysvb2nBjVpiCZcyHFHfrLuw0
50zfZZ6rx9FZ2/SNouytjOijcWWSxutvz7VqEuPsXIf1Wy5XICFsTFfhQtvQMNilvU6xTK/Ccoxe
heueQGGZJ4n7M75h/Wc3NRDkzuagzIhyHvgFruZY8NlJe2x7tnlfkv2BO/f5lWPNJqvCYf7uh26u
6gCzb6r1qOL0Yvy9EY6KRKSK/UfriVKSWZ8Rvs4HmkrpBpbmz1kWB4ngWK8I1BGGX6Zg4CSH48X6
uPaU83UiX0W5LY3Ka0hqGj30H2G24ZFZ35rXEPlnnKNuCjTYK7NyulSyCngVqNOZeFvzvAxnkyQh
Yc7J4erFMf+fH3JyxN/JNJsMAuHUh97PRpcHUJt2UdJPD9jy8XvdSBWywoIWRzH6atX+q7HlXfJB
NXDjnwC45EapQkZopqQqY8i84xEY8NuSNgoqcLW9x+z6kxlWpDCly3APDKDkf4rF0miNvFJGNTlG
lYusGXN2EHB7/BbzvoKLK/g1Pxz4X8lp7bEgLLTuuk0cyV6lot08EPW1Bz92MKuzUh5ai9sebcC8
Jyc2SVMjItCThAxttCQPa+cKDzLk+oEBtPt/Keu53OZFzap92tPxNOkeY6hdxT/LceQB526ob2Cn
oeSr+UCzjmnBxi2E/RJZ2M8sEKes9LOsCBKYs2R/qCKMX32QfV3tBxLP/hOFik5dM5IOtTYLInH4
XOPGYL4iS9dZAq0mcX76trbWp7eCpfp6pWEaIMTPzSFSbEBS7VBxacqgCWnLwnMhrKP4m2ilUg7A
H9+VZW4zZBnYFLiK09BLjBdz5RGJ+xktbE7xARn8paHVAzAq07CDqi4BA/+8ObKg6JdYW59khGmM
RyxNGFi776yAtUp0UoJCb1TD+6Bm4UkKAYN/WoO6WXt2Kbb5cGNTRTbGcYYtZh48CFNBD5zkORWy
u1OO/m0/Gy5AoJ+chf5dZHv9gdFCPUbOPLeArbuhwO3Zyl0fsyLa7C1WHiQDut2JHADrqqFzIhQ4
V9uq+lqFvl+kDvOCdEp5nmJTfCyHL5/Gy5AWG6i7mEawuD4mNfmsbC/jYIIpYMiSSXpKYEtOreJL
221ZNOh9g2PPgYNLO03b4y1Ugi+dLs8h7K90O4LyW52L2JKdLUN5uPkRTfqMjkq5Z29p8e32AmKq
81D9+04FiQaKrRzUGpCZ29sBH+WOI8V6lcYQBT7BJ6mms9ZRcIXo2tnt7UsBzNyJ7OObmjOMxeXa
Hjqh+m+xrojY6SItsChUSk5tTC6kN6HKSQR2MXuGjtpZWqT66CjXFtDd+65JlES+KwkSkMm6+IFE
O5ty29zao80+4kz+sl7Ju/GY2hlUwiRe/I1p9CtBgyKVqzQgPvpSYD9Da40UxmWdG9rHrOI2QNkC
ePNUIxPZaQs2KIRu95frvd5rnzZbOFFvWMDyiOFprKfiBPzqGDwSFcojNXLZgXV3cLxm4XOR3P8U
XbQQSG1/SMnAtX3dTVG5Ljp9QFhZSZocdvezTZt0R3b5+Tuykxgc3GVd+wjHnYifV+M5sjGWfdzR
/96mlhdrezScZOq993Yov/5O2gnS5My9Xb0W83tbUGI3x695O6nkdCaObi22CQ1QLwgNgnVnqkHJ
1wDDTlsCmV5lFzyJz9HTDLkxmDir+/TY8xLrNCwWJkhPsQeLhMYqZq+iElG4qm0TvlOlAm2atBtt
Ts7le2QjwPIyLaQ2mud5k3IvHhlp59aS2cam3s7K8mgM9/hp2id9fEarBak+rxB/P4NDksKVgr+b
G3hxcaqShDMmwrqQUL0JusUWBWxGS66/LxJ4BK6g+Qqdil0pcPVK+6Fur60rHsMYh8wXtBO6Zm28
lwlKwDkWRX8xDALVWxwjvxOrmRA7v7tfc0ChrteTezZ1aADVhhxEwTvBm5h8j53lNQyKLyYKouq1
I1waSc348l5qgdXCuW33O9BMFwrreS1VnhlA/v2fMNGk6OW7R8iPsD+OU5gG1b/rXslJUkYA5FIS
bNc+kcSX+mtOB0x/ps0KghlT96sRkBKwZmFMwUmNGcyw+kVhzP+wHIs/hllaBUtm3bS1YHt1IbrK
Sh+Pb5rzDYbNuo5UYctxXdRoHyhDcl1bqDcCm0v+zTAgpkgcoRQSS8zeSyHJ81bMGvtA9dXlzLzq
cR7P4x3qf7klvpDELBAPyMFr81mRVH9leMP5mhFB/ObSpEy7ZZjJpeyhQ5WBBMY1dlUnxDajgdj3
lMSyx1fDf43sxbjlbggdkjbJJ1iFluAcmYhshY3vRyU91mKNY8Tx2IhNTEvdT6ehkkJ8VOvxeiRh
EsFa9/10qmmDweN98qBFvulGSybBKYWgXBqCFPZYG/jDT/C1TKKQHk8E2ej7c1qj5zAz6QqjoPG4
kusde0huz/OVrc2XAq4Z0rTdwKQf53i7/VMfHY1W0ADpiNJWy1euTXGBsbsm0QOO/K14sL4KIfCe
RNmEr3rA13WudqUITVD8LJEAdeiN3rlFi5jOV+Mq5Vz/p++z6aw0upVEuyczd/ShITUeX4jDhMZD
DhvhtwHJDRbnVCQ5aYXsb6eKz16IQHFuSeG+HpmlJTpWztr3DzmIBNF2Vu8OOKjBEAjmOD9RzA7W
uMHDCmO3OBaUh3sgL71YEwoTwnNvOvRmTXj9Dv+gad5HOqYqhGBDS93yWNSGFy86/+aP881hDSS7
NgZB69mp6kPzrY4IS9lHeOZQB+Y0GXO2OpK96Px43SzH2sBrVGLkwIZPhAJx2xwCz5kgudcHpgSb
6dwOQSAbktyn/y8QOAlDUpI95FOR6LRM+aAuO01KeQ2qvwBamyecvOWUD9xQtBcEJSF5G00z1En2
ZsicE3QmzBU0xNAn6ffpZj9qeUBuhGbRafBiO11eSfmZccWFv9FleGbi2ixMxbizNJ/HW237UGG/
1OjeiZNNgMa6pbFDw+MQpwdRfSxpVqdQqIV7FDaInI+Wgb7COYrn5vIcnReCbD2VrepRniiuK3XY
hBlJTM6Up3lqmEU6vLUU0NfIVDcdULvi2kqWgKcjsMIVuH2Au9pqiicdrT3+edIT/qTHsNkCVvVX
SwR85zrs+pZ9IOk9bnrW1PwL/xxHULrkwZe3Pnq97KFeacoZ82dtw1EDDo38rJJg4Umh/20nkaRE
cL4BQmOBjWCX/tfMPAUlcfVvARSiCHd2lEok5WZo9ygZ3q9kfqnvIDQscIjpQQomubyGAscCFRnY
Ad3vdlBuXzfrQsSICS35Gyp7c6cmuFN+Fdxi9Q30OhQ3s8plX1hEVlCTshTnllmgv+bUD2CR9Ji8
SAP8MNZRrzO/Slcd4VFKD7YBPBBYIUJgn8vj/mJgJ6NohuSE6OVgxJGV3WQcghpriSKI6F8w9q7p
62ss9CK/RCU4qrBpxVNhnS7JmKpsT9rAicD/HLvCi2DX3tEV8mV+pd25i8UHinWwcI7/Q3KR9knj
b25yDMoXTyTMtoPlU2zzv1G5Pd9XSYV6+73p8ZCSgGci42toKc85oDBSPcnOlgbEFLlaSGpZSDoR
qNRuwByw/g4gb2uqzE5PimZ201m6oMVE5kkcz6d0JOLg1m8+hVDqzDFi2Z9pwuCJ2Rr9oFJUOu7M
LHp5iUngZjHGnWScMkKekNwqGV0zwMOnOZIFf/PkPpCntjmG8jxgktTkJ9KdhLwlPO3iKuwt4Fmb
0k1As+KChM86CNmSWUY0FCCprzI3gyai0pdVsuYvCiws99p0ZM3RSdpT0IVfs/zKvIFy1x9m2mCB
VHYcQOcMxgGfrJVfHdj0UlyubDMAPvXwwtpFtaso/f/L1C/Ej3xpQpFwwlTra1H6G+yBXB2tm7V7
APvOHubI5UWb7FcHyalLqFam9z6KDfsqoAuIPxcBYkF82elVyOogUKunPe5zDJ5jdSFgl4CrtYFh
pxvIe8gsKPegICOcB0ZgBvO5faHAQo0eAYjBu9t3sb3MZQoWrtBnuJdFSFD0z5q4kDPnmiMRihrb
n7+bZmlM+SLlTQ+DGcZZIZAMAdV1zdVtVrfbXZsUIM6mt0M1fGLmcAy9N5JaDMTZ0U69r7AuGu6x
lqa2xjcvoaVE8hA8XsAiEzETIR9R9Tp79AdFq6qFcTR2YCtHn1gYEojxvtX2uOR3Xv5jm2VXrykl
7XenMLsgbY5R+WCVPYtKZ8kmsQycb/m2mSB4xoG3ZF4BNHloXBflWImAcjyzabcLyP6KKv2uLIMw
v+Ghk5awAWpOfQPbdTysYRc6t8ogurQpkuaxnfQmQ1y678Jm0VcyjWR2AaT0ly4XLwVdMrj3ASVE
2ikdNrenP1nDECfr+zC1neoN8VNPMgJqHmtjFfMOeWHWkiIa3F9NijFyzBu4ZD7YOimAPwvd1zCf
Jhq8jBrSVZ/UD2gfBEaMQJjPo/IumYV67W59i3S6Ht0aTPQw4UBX+8ufPWkeI40cQDD3jMAUgia1
bJ2lhybuIDdfI0SAD3SAn/YCBFgOYdpYGDHRnLBg0IevLjcgPjuKQVRUpYwS6K9k5rFS1x4avB+C
cOFW9iCeD3Ay8w3kyCLntm0GZDBk7HeboBdNCLUeEFFOudFzdGNICHY8PyXF+kNyv2JFe/Ye3wFs
pdu4rlsBHGT+Y64otOf1+/29lIlNlD5dWYUnuaTQt5Orkoat6O6qdfPquvo669UZDAhF+n84dmzT
8VFPlZ0Y+vPPH9syPxKA4nmv5TNtTcynr20sRws9aniSShs/koL5b3raO+m8ShKN6NHSQhtaVLRT
Sb+UywLLbO07Pl0U7oGe7QR++btyLYVXsiGpGroODotGxRZdY4WUASwwf92rynheirQ1q6uld2iB
PbMz4r6gC1e517f/DErsXFWYuPPIoHyNIBS+C+Hk9SNP/If3k8FRJR7ztgovseht5erg8SjLnjXf
YklAKZ6FLLm97VhLb3y+ibpqohIajcYuU21vruM+GMuhz+BQTIPiDmtXJrd2k1sGKSm0FDPQjtbW
XZBv2TtG7cbIcF/YQI0R36qAZ/spRVgffIfCM0TTo8unv90qmZoB/E6bfaSkAp+qUv/NGH4JxYd4
/EZI2Rq+UsllIWlsJ45R4tA+q0l/gEjyL1Fve7AUTkyxbWyKUbzdjoF+6zKMsNgT3RQQ92G1+fk/
WGpQ4TJA7v/RXih3wtWqjdj9LDgywG7viFjrgdw4vp7Jlf6pmhQE0x+MhYxhzRMwS/pUkJCp4BET
DX10HpbJ2gHBd7O0mBDX7fmfVkwLdYFqWpzalxfwFDUjQA+/REvkxrEhHgrRmHPzvKf/X1/RqXhv
c+z5h2daDbwxl5+UL0Hq2hs2AZagxKvp+doeSSDYoXnPioeQkbeya6hb5M6qT5N52G5NrnWDby3Y
bTExGEZ4B+UEGZ2HxKWGCFReUoUaqmqeb2DvXgjoiK7J5GwP24H/2TGDV2lYcvhlCvxWAbJSeVqU
LK9Af5WpLd+iMIRQxIfkuDGgYWgUJjI1b3KIzmsOEBGhZUpv6vFSiFQcY+1ZJuI7/Px5ud+DBswH
m10qMrNnzMpEa1jnAGpvcoJF72QK+M41c0pLOo81jS20Po/bjGYso3O1SxEHBtDhG2aX6lDVCv+o
voDHQv0TH9ao3rYTJweEZqSap0F0tUeGSs6+E6x5ZqKnmFmfEtWwMSDXAT4c0RHHJg7ZMAtWRKEx
dVQYiNGSIW29UD+ta76icnKcXj8ai2WFmTbpgR/0okoVOe9ubWJ60tKh31+T/5BcccdQ8po2oVkE
uncJye/ClXFNxPSToPinsIjQEwIysfvXaCI3k9a4fud5+EcSmFLJ3Qmh7lnTevOS5JbZT16u5zEH
w9/9J/fjmvaYVawrG+kzCu7GBRsghVAWxIJic260htVEzJfzOVCr+1uMUDl2oOZRpLUlWrFrU5L5
dUlAXVFAq5BUZ381GHplowJrVJR11+Du0/avNjQiurqAln66KuEhH5MBJX8+mrIPQT++WgOc+7mA
MFrE+QVdvCbXTeVl740L4ezyAarQr4vaykzVXvz1gwhNPijHPvc461C6mzFjpudO/euQLYfhCXID
VHKIPRWn2ziPcJXKINOpZ8HIfEM5/QITvpZ60mA4IexlodsDrYFaadflDaDkUBxfMpFzw6nluuLj
twr7pRPB4VQsOLrJE7NX+w9hYQO2LjLoQz9mGjTKuMEDWlwGceH0WbaZmYMVK5CDyqBP7844IKUB
pPCYTBEdbUIkXukS6yf/H+IQ29V1JL3l8pEAtIBeMqXaAFpQYCnbbfhmRq0ef7ojs4kbWhX8/tLq
ZjnxD1rQruZYPRR+efI6XKBpaPE8+drKATRoMe9VNZsa85gvRbEvQNUwjxpu9rC1KyoUOIj5HCZu
7RqCnU9ByxDSpoe6LgFf4mLX5NTj9ZD6ZPYJLUF/EEeeBRemTBPlvbZ5Dy9JFjkKKnKB4BHaJCcp
mxI4l+2oF8DXb8YGkfHpOdE9tLb9YF8qfFCzYrdXw5WXI5DNwnKsS3n1334F4GDhK5SPiRS4BJ32
APtO6D2EjJ+5fVeyvKm1RpqivZeWFc5BnvR70mE3I74DvTDyQiBoOUAYOFC07/ledIFz90seM3XD
aWGV0J83S+47xVQUq3iWNzlDK93ylGBq0kYnjyxxgSUnv7wiGhVMOMz4DKzZBRyEoPz1lQqyFCtw
rfB7aXeqnZ3rRglByjFFz6xKCQlmvz09vrVlVOeYL8ehJglUP+9NyHMt65HQ8nqYFVFHxZVFn6/t
9EzoYAm1J46rR/60zYJVJb+cE9tkO9jiQMgfVTUIs23LrLHq2jm8O/1teghV/Vepdp+BzT1nfCoB
6Asgs2mnZujG+o/Ksg/dootcihx/LSg3nImEKsHfqTUKqGr2pIzpM6UdYW42OD+gnNU7+rbUmqLH
1YuQYY08rUFnGEoKWqMg30RzR0PxRhVo9iHEbCSnp+TdRP8g8V3qAYkSnaLcHou5oMi5hWbaIZdR
aa0qdjS6ZS2T5LlnfIZ5CYXTbt4r8eYZZKPEubioGQ1askoYktEO5ecrfBMLl7lAIlmkFDGN3hR7
nRPUxJCteBsXcpLOps9DcwcFfSMO1eCMqw0m39jzxjtc4F3MW8livpB1/awKEc//enkJH7JwEXen
OPdhNL2lQ14XWIKLt/ORQQJcMvjjRg+TiLRu8asAA7HtJ2JJv8WkALFaua2SEpMlcP0FYh8qthUn
JdmC5VtDOjelXmgXCnwcHokOo5q7ktbi4x2S4ywQox5nHi5ndz0ZWKqlttGEJlxORUDl8+g8GS1j
/4GrxZR/QxwQuEDYV3oTwNslT+21UUgGF31Nhm6Nkbo5xLZT/k0gVqStMNVHg3iKH3a7z5ccv5jt
65YMD2vDOLkZW2b/CDRsfiq9ZRm9BuNHyBWqOmJH03p02m3+gXL1IbgS9a1Vo7wSQPSOiP/PFTef
u1OkL43qAVRG1aqQXbJ7JTVfW2yRqPhhPQe7oeDOhTtoI8vNlk/xV0ZWziFqBdzpma1XfrquPM96
EOPSw5kwCTIi7OtsMTMVaw0WMN7knbBoC7w3SkWc5VlvejUkODG6sYuvME7tNHxASi/Z3v08qL7n
7IRTrM06ZaM/oAbE1ILXRi3Vr1UJq70kBVfSwKIgi15ALVZ7+r47b5+ZJyStYK+D3atONQwhKgfu
Ifc+Quadlg5Xt6MSA8Csw84+G4HIaodD9ZwKc11WJ9oQIG7GKy5V9z2zMNPg/phNiRHYG9eN8u/0
/BL0pLOTbtvtn75cUy+H3ilAI0QBIPFev7X70NlGa8zGQEbESmT2ATvbPJqTk1X35YEdY+0SJMyB
3pwjoHuHVtGv755LcvyhL2Nnxgqc7ltiBv7OrfjTWfbLv7xC7xcF1qwq/zJI1YecpWwsIfRegBwg
PKIgkf2W/Bz9x0jpEoFO+Lcnh3D62Pwt0+ieUfH+jzM10YVDHErPXUTmUCIkmsic0ckbcTMPjNV+
Fykl1j+WH2iND+hvOPnAaDdmNrayDQpv9OBWyA064Fz6PdFXvjG8aZFgwDKbDyuIBoHgjr28lk77
/HePdSbqSGkBr4ML8xwqAM7g6JvKqa+AqvhmYOlvOA5liSuJCsUOE5HqMMuDpq+mbWQvW+KtRDNP
CaRI6JBefUOZKRpSWr2euFC+lWo621luQ5A2NK0HSmE3PncXnJssfvJDpYeqZdowNr3lUSiEmlZJ
/UY732Nc5NwgzBS5KkCVLPEhA56EylsNgdm6k8HQM50AMT4dbblpphAXDEF5UFnyaRP8uM715FMf
wrFQ0pvjfHoknvrpfWBHatp9vW4+roeCF/ATx0gYt3iPhTnbe5wBuQtCn7L63IBqCLWEAn0y5tGZ
raczePZo5I6EzTzqiP9OMaIswT8h2gds59YQ/Yc6Vt6irRBC+m3h3HtikkFiCsN7fiUYw701hO6K
iP5E3nauRMaHGzHgiWf6lepkjhl9d98xXimMpHZZQs6aGMVmXC8vn4RVV5wNSulFwaikAJQOlCB9
wenOq7CmEycutN7L62kocODDYJ7vQ2AksQQ4v7aIaQp0Kl7d09ULkDLfgiIOnmVjPinIChENR+Iy
uEAfs8Sv7sUQlx9RKulVXMS9LgE6Ix/DSrtoVsBav6w3ctj6V0YikzePRkN2lVD5jjnsLClhU48T
In4MiUt/6cOFb4S2m2DFBUrroDlFUNRdkKLU/2QFinFQ3jxTu1mAsmoOi5c8px5irdOmyrlAGDXa
1o+vuuCkwDfvBqCPvj79KFRtG/QFQGSazklkPa1tyLBLK2GDcxUSNUDfnXSfASLWmjjgWlXRLmjs
O1p/DgjEnAR4CqzkyKhXyXAIagbV54ESFN+bR+o9dDJb6NrC8yJNxBvEaAkPqeiiydJgVGyRD7R+
Ot3WZ/1JjqrW2DbN6p2tC7uAA3TdCR/BCqxmh3AA1z8mwU4ZotZt0z0zezEGDsZpn/h+2L1J51Bh
LTBq0UVdZT6cimGc0Q3eXOiPNCH+2Oo+PTHOzjnIThmhgma6lBhRvazk/qYBZXjE8TmVRR+oIEnO
2b2equfrvHpaJV5x3S1b7wcy43g7U4ZuN710aMj3JM37G3SV5VoIQOH1nixVEqYQvVKv/SqKjkp4
TKu2daDJELrNHFLdokOTP6+hrW3K8rOmNWg7dylb3C+ao4RxQfLbTeqIzh3NzL+hTitai304C8Mb
xwICx7u3ukOw64p/fRyqjwTNkvY8vCbGcNtC4YDdOHpRz6UvBeUl7ClccooKo0609HB66kuFVs2l
CxMkBxYftb3Zn5Roqt1z6A/eduCv6u3rtIlTztAvwbj2sVAUpbvaWKgpuhcD7qSyucXzl6C+90bk
Bae3IZV+9cfoM3d+Le/Mfwe1bzrzKhe+2AYa6Zdqfbm7+wiWsjp2j7blIc9nUFblsGB96Cq7hIAV
WO7KfVBZjio6AcB5h3okbd918P2uWvsU4nAd27WrOEFyvK+S5lzSjjwTJ/lgXT1Kf0CFdj972go6
QCq1MK9UOBWpZwxKBQRIAfuE/O6StE8bd76h4PasDq/GSYkvsRhL49KGEJov2LTQ5QI7EmapzapJ
Zo1hBVSIg1zYaUgaisre2KMnWespKM9tWsO8arNM0QOWZieu6OeR8+H6xh2mW0DJWeBvYhXvy9KL
AHvtxcPgLYxIxddtbAvjKYbJR1pQ9CTuROXaflriG8uunXtrT1ux8j9VepAkD9aLvMnW1l1y4lyg
h8E2ecq+3q22+h5mjGnTgR5rOhAQejn28cdE84N+MnnVqywSFOXfNWYDV5JwtdIWU72BQJ9fE1w/
3JA5mH9iwFT/vozBH83ih/2B9BfqpqbXwyZXal8SzPmzVMT564yhaYWTTr63EOZvI5NZS+bIUSNX
obN270tdc1Ls95rUxBwi7pSeyFWkcsxhIfiJGpwBKw6IVyp2qT3kGV6IOBrqTmKbvTmPIm6im0TF
D2vKWOobkpQ9kLsK3jC5Vi4bM/L5bNSHkshyW8rkIuoBcY19Ie7mN9nqb9cn1ELrUFl0c1HO9hX5
aPqnJEv6Ec7BpT2kDdz5OJfPGEFDKPsyDY8fC2ojjCktQC5JzDeIlCb9LJ/mpBF+90U2sxfRqlmQ
SZ1FcqWwXNvFpwVbHCaf3Gpo+kxjm/sSl3cssqNscoI9LfsA22Mhyx4Y4SnRQh0gcvks77GKaPVX
nLV80sGJjGFo3jvWBU6FqeXPBODVESGGDCn+vHQH/K6xJN1ThifTYBjDjXOpn146kCnHCe+7eeab
JNNXbvRZUfiAAEn9QgA03eBzZadYoCbG6xgE9WEW5xzD5pEhrFJauSl+GjEhS4PIGH53Img41I/a
b35Jt0HeJRuulkIwbSPuRYFdr2iAMAvg4c+X4EtgIWT5TFgtqmS4zRrAB1x9lff5H6+QDjO70duk
6975B0naqh4EZjzsdTgnWGY9i7MnrMgQ3z2f2Ru+bT8/ZH4cnQ0tQnjnRJu3NGWXdKfIjjEuT3Ck
ZKzfU9h9OnxIXawS+h2pymfn9+tozQvBX0UK+UakBcPGXDlhFGvG8Ze8/Mv+U3E1ycWEiIiy+iyU
NvcbX/FkJzdnqS8MZmpr7aFLEqdNfJ01w/KDCipYnrav3leAVgf0r5rhPWyUEFFnsq5PugMi2txZ
T8PC9XtZee2wwpccleSkWSTFE7e0ohLNvZiVEKTLQDLvXMXjA9ykm5sPQWYx5W7tEwxPTfguJ9w+
mfL5SNEk3IsJNze6Dbzlx2XH8feNXP5MNc3f2hLFpc6EvccZEKMR88rhYgKcSNNhDUuDAckDjZbG
ar3UEhN84sxBBKWVAncKAq6AUVyeXp/QnjG3QrLRj4JzdpfnFwJl1cFTI1eHpvF/k7Cahdm0gmac
vtauZf6UoJ9owZGlY9Saly2pakf0t32oeV+HoeuY50l2uW5Xv4u329P9kyNLG2Sqpfj/fFCbSb5K
yKK4/cQ/seGsFHcQIMxScBt2JgD50I9ewXDs3hJcducTJzYpGcvRkC8J4Wnbsj+q/Cmt3kbWVRLD
Z/g3k7RqcHLna5cwnqYaEYw17rGcxMfgL/VnjT2l7BZeU3CXdECJrYy4u2ashfug7MhBYQT2cLg7
zlzDD0MoyqaJXMDB41auviEYiq/rHIt4pHMfE9FtcL9C3b6saQWRAoZnD6fBTs773USRb6KOqUFg
W+yWfMEL9zeKPdxquwrKIYJJFdKx+cnfI+At/tTdtmqI+WSqM1BKZAMVm3TcDZ1cy907LIkxy6P/
BQukYsVUfasTA/L5uOXYcCY+PtHW09pPUjACGddhMQFTS5kyxd7SmNroIDdL2o2Cu8s2pbc0gS6G
Zhp/4yB9VheX25oaftQw+ITjTqqxSXM3b4RSWi+RjRi1d7xv+oIfTjpJIgGMoiv1ypgyowQmR8Ac
Wldoyr2z4pS36fi4UuAcCA5UmW7Ngw2ANm2WTRHkfiQoCioFLQWciCMHad1v4FlbKBwU+8hGnqaU
PjiIeRoGJaP65h6jyS+Shg4ZphNlGtBGcKR9UVI2XlIUNMRa89Twvlpt9x6bIRzXfupJH5Qgp8VJ
4YPbs0MDewCHcUxSlJAWgekOJjphmxckfmg7i1YVt9OZBr/hByiTSMJmgkB5Na0Yl/IFEgNkqm7q
c2CcY/De3dwag19vNrQH6aCFGD4+HCqyNgMOliizcxLBgZ60x53wRIsP0g7e3pxayYrNiI+4WAzZ
T7WBwIHvkyUoHAbphQ8wNrneoOj6P68FEASSMeQPsgL4b3hMAl3JU3PzURdqOYpXP1UMd4B6CIcF
hfJ6EwJcWoZ4h4q+MeGfCQ1VUjK8DhPfq02fa+atM6i5bvpny7yhOD58ElP2yF9DBhFZDclBax3P
fC1Goo+HPihNj8yGQtHHreb6y83CDliJe32JSqnr0ceCNnMoqVuMgzi/v8ndObxqk4xzpUTpKep6
9pAwA8hJdrcdJbknL1eiG07h8KrJ9Q+5ngx9ni5TqAXEZocx5nkDXOfUHSfVch4hSIW8v68r6vOZ
lyiQ13RWzAMzD5/jPMZGVSZkTt/CvTzoK/saO2WFA31bchup418CoB+KjRfBjYG6Ahz7y9TkZnyu
t6vcu+9HGXkHC4aEXv1DiprxeC6AQAxa5itwbp3tlbB8EXk+5Gi1j19b2y9l+kSr61S9rSeROp8e
HVsOTo5qgAIHO63itU5pQjslz0hFyjD67IpgWcwkdiomTSBFAFgwExodDVXTRXlg+DhD8QkzTwO+
Yepq+iqcPkp3fi+ruzXRE5JA0tttN7WzL83TDmC53zmIO5qoH9V1gg6ikN/54qvAovCfHEFV56sm
fp6l/NWdXzKnk0A6/Mo0bchJq5Js3mmgXCT5N9sII6RIGYgXpiTJHZwuEoYQW/xJxqlo/EkRJHKp
2yPRRQN7A0Lx1SS354Ezm9HA0NpUm7bIhHrMN5czd/7/kQk9b0m5Clsj92fmMrPu/H6LwUj7bZsQ
QS39oBtoen6CIuYym/24g03oJ6LEeec9Ojfpc9LvzgEkorvcqPSl2wEodE47I3l6jL7xTe8rV15V
xNUdrWS8zvwzuWzHGkHdiF7+upuy1lz0DWtRf9Yj/1mmH3zecaKO+eR9AX6ljD1StNsXEmN1mzww
rpZm5zW74siVGv9HQQ4y9Ju73AImsepnFZHgA/Q3bzIaWAjNubMcV/qSTrlZKkgrXoH7EGjRuqAB
+OO9tVPsq4wkJuej54ZIs+AxJhwM4BVZEoOcv6DwEwDP5+yrUGheeQLDikMlvboW3z8AcIRiXp94
rFUgcm/8o7NioQW7P5C4O/KI8DjTPBPetSaji3fX4wJn9c+OOFzf0vIIpGV9ihGv9TQdAlRlPwvP
/BuLVVkNnlqqfKqoplHki+Yye9RaErbsD2hXS9wz/53XroGnwNMOgyKTQzf8rnUx33u4IB5qMiRt
YrdMDCKhs7G1+NoqLyy29UE98aqnxIT1HGpfG7oKO6YlzF0KKoaXKJ0hGhG/t1gTD5SGQ6K2gSLk
M235JasIhB7OqYif2X1XrQvf6Oie9NGslKoPaXPzw9Q9ySgk1hD493FnuvGkaMQXD/Dg3WnEnyyt
zeasQDkSy/2b5A9b1nDxs7eW/jnoSk3M7rOILDAQbqU6ki1uo8n3u/Pd5AAqqOPeRTmbm9gW5Sl9
OAspXQ7IftvkzfQ5FnAaaCwT22YliKLtTY+8GlpwtWUiCXOp+9AUyiTRuGTXCJUkzD0S8ykAAnYc
tn4qhKvtIHawh4nGAE2SAMOL5/HI2w+GoVi5VTbykZPo25x3YfZ8nfZHvObrwOQvvWuy4Ib+FzqO
bxH/IScTaSsewWUWvB8m5inAI9zWXFmA+7vXcWPiQyILhKGgTeFWDUey7qxdNmoj+WOeXferCw1w
jMLg7ClZBkA1Ial8gjzkr1CKztdDV1hIOwGi90NxZNZu1Y+mOt8MaL5Z41nOs0Z/ayrn2vD5Ipgk
Ohq+xjC9ARuC4hRWvIsZYPYsiHQ4WE891Ih6Mpi0Dcvkn2v2vp2IsyE4zFMcJ5wY53FiGYTRY+sA
mHHnRjOEVoMp+CrE2Elz7OzMCQXBhUrXB8URa+dcrbdpv/vBPz/NiQTNh9uapQc1irDa1CCExj8e
MhAomAbosWI4Qb4avAF2oig/LDBtphw3VqH4BQHY+wDIetwAy7z8fwo0jDNjtajqn5TSF83iLfav
fl6MInrZA6aoFz87qjfp4A537jwrIBVYtCoR1DHUXe5Wd53WzhW6PZcv6EmKV/sGHXKd6qSAYBO0
kg3doiDhNUyNYHzTWzQMj0VIiCgpnxXdK+qvdBcAs3ARAIdyc6er0zQ2VWPDvlWali+ZaPeC9Tiy
9reDeeKQIkyrdJQlGmhG3Z2/+iMnAI+A0MFQCHaWWdP6ATOc5FMmXItXzZx+WOCi6iZQsBUS9UYM
HUSBUVGBjB2rf4Fz6vZ7iRjt440Hrm4bu3XpPsbraT/pzY2BTxe0W+OEbsP47XyToxoHqRWZaht+
78qdI5I+i/SROrHeKS/5mi8yMkGcvM2X1VFug37oR4trcvI6i4Kx7Qz1rN6NeNAV/yOhEb9vMw5M
LWdcUs/zGXG+ihae6lCW9dXXCVbSAKrwfSBH2UbjJkcE+vm+6tyIMS+WisCtt7CQe086KSXP/6n7
Xt5Z0INgnHTVF8LZZ7FXbAnPopctI3P6WRef5q+92RO7mcdWIqnUxKdOaYxMYVOyL6U5ZIVEBOAU
PoZ3+OFJNgYmnAGTW6hDd/f8AQ5w5YuqXZOuvKhSlp2zc4x4SABYFwvp5T6Tt/z5gpk2iL9r/KTM
9DE5o9xcbMPUPKbPkVu5fZzTOHUHH9BYlmI+uzB/B+rPWuXfrXfN0MdoXhQ8HDTNF0iodL82UREp
EURhy226fR1jtJA0+Wf+iSNGHY8Q644je0v0qlL//gWZyEcm2FQNJRF9qWRdO9EdNz12PLk6xpEw
FtMAZAgpj5FlTZM0nFDq9Acr0h9IK757oKlgKArWOkFCdueJKu7F7RNNWP/qNIi/DAn6jRq7zK3E
SMHA8+t3L0MGZmK/49RBbgXDsS1gh92E00wH1qI7zmhosKy0WwA7xOvIDbtVFqvXMEoMVB0lvxOC
t3MflUaT2FSPcZuOwz1BRQhb+Iq5ZZ936TAqI8IFP/CDQtnmTFmmy+HwB32+gmEcZWZ2LPXvj/4k
BOrkMptR9Xz9mDa6qu9tABRPgsYrFweumnjmdXLYnVUWOggaUc9lPfGoVv8GmRX7Hmr5jtKGhuYb
ymfCL4Gnax8feSWlSJSq8m41f21h40oVjei4Ap2ClerBdwbNzl7G3Nu/HvFqZAIQ4KTx3TVxyQP2
XMwYR26UhXvqjTspP2TegslM9PEsbaP7o4FtVri7LvjfhfQejcg6n3YIwNlUf6jOkvj9A2DwkkdY
0HG1OmzOeUFQQBlabG4cHyyqobZvdvm8UsoZWselN3LBnICbzeuoDfrxBJTw90etvMsfp4UjdeJh
FP1owsk4hEecXDEYw5oNLHwKHPKH/Zsf9qX5tjJX/PglsQmLh9LO2Hxro1N+Knb0vW7DDSJGyI2p
/7XZJuj9lPh03RbYvVuOoCBLZv4K4lEgAQW89WbseZ5IoS4w2JKeEa1EvyUblAk2ca6vY+aXzR8D
izhsXe9JnWAy62SAuYXD3bceiX7tBnBEjBZB7y8IL6jOCTHayizbMvEQsRn72hefNNtL8iycNKKC
JAxvxw5Agem+N++gy58MaQxOpe+ToKC8Rat0uG9pihXujwxZj+XVHfiDEkKTPXQPMISnNX/EYFtr
6+hIj3d8vVh8mlrmgooymMtEeKqvpSMr12875eMi6fgHlKjZGjRmc8peczfIAx13hlNQ7SLxITet
tvrPpvs5FUpZELRoJD0nSN0km1qu0lgkYDoLyZ95IJzTEz5VZ1T74WHJSqDD+KOaDCp7ByWqxCGa
6VYZi2FmiuRgk2S3JTpX77zitplmkVhMUIZ/FAxMSnW4OCy4R2wS3LmSpUc4GsChgNeii3lVWw3S
IaKxmkiCqX2Kwc83RidH6ML9SvbcECnMfgFLlxFUhwJioYRxNFFd+dpDkLCuGeSefE1AtU74HFx6
tt8PzzTSTsjnUFOhnYUBVc5yFQvlajiQZ8NzgVbJRwovBY/R7Og8z1HOSSQIk1Wk2tI8h117qRhe
VMA0c1tPeIAT3JVUqrDUergljBR6isfRa8TUg2fIQJYlanbfH9jjgl3lct3fjgydU2rY7gWiZt5b
lE674aVgd5ftANEqR7OaDYF7fhLAAi3XR/eDu6DB/LJ1fWDfyRVJzTF3JhJPUVmttuuL6iLJ43VH
DjKg9iEJq2VvNLzBA9R1S+hTGoocpS9diArkrD+UHikGhK3JfJyM9etPT0dJnXSmIMJzcSc4Xos3
xmmkSQlxZZA/6zRYk9/W2c1Q09hbmFao8+K5VtRV5WxHnFdo7J0H+EHuRFvKnv1cYeR1RGN3JcHM
z4jtGXTbW4skwuyOfvUXUypJ2ask80etBQPspii+zXceCyFmGSffO3fgupo2ZX8au1bTfY+JJchl
+BXJOJ/VrllrYU/VWh0kjDCKb9syFPHClIyD9iraNSNnKrdM7jhlKz1aBoKZjbGBMs+ppLEb+q6J
erDYGUj0PcVwDac7S/hy9iCtV0faQynA24uoWnirusrmIo5OfKMnrE8npciHSIE5HkPnmfrVPDrL
IaggU42fNKj81ebrbrqJVy4F283fC33VD0MzQewcEPcFc9gQIZG+k67OdsqJLaT62j5zZAmt5bpQ
kn7zRbreQ0/uwcjtFR4arNBShwNgaANc6Djuoyw2zOaMwMo59ngKZy/KfGjIeWyiFkX+sMYFIi8h
NOJm+EzsqdjIb7heUmCHQqtaMAbl/kwo/WLpK0WEp1Ybht4IlqSUPsGKxjCUruWNNoGkFiJmVfvH
DwCKHaMbeCh4QjBwitBhrMVwq94OsIkoogAn2o719tezqKJ2fIAs8gBQ6t5VUkXPBiIyw0UQfY8W
5eaVLiYrWf6b7ozyDSDD2Mf7fsGEer1Tys8DEzdHw5NmdqMxo+vVsHTnm1lV17JGee+z39wuf415
Kjd7oR3wbDvkLlXt4Xts1BCCSHdFfbJKjDS1aYqtNhEainNMcTaQul1nhogNAlmtbphXJ6t9tUXZ
zAv/aNr5PVjUSgKxnaA37uYyyNGcFWXoKVTGpTNEA7DHoSU6Ab/zoQFk0QbXE5g5RrqnrPeRI6ya
TC4+0/qirf60IhVwF+CEjGw6M7lySAM46bL4HC0ef9Znnvj6FJyu3/DT+2Vtcdwk3xYhK/iWIpoG
Toay+zMro1uJ1vK2ruRnpvMunACUbzHBtSOMicwMToQPieKhdLOsex06BLx2nJS9huztp2JTCFk3
sw3FXKR3EDh8UWaxtl44yyeUaZo8oCY4OiTjQc2hivZaymWC0Os6tLi7UHq1IRqHnwkgSNGEWZxm
T0XdTBHp986fOJNBNBXpTehV+O1FXxWV6TH73xfpg/sSfXcu6hRaoWBsF3kd3ZWbE+jTSCn/iKu8
szol3s9qqvlavf07RURpVwE1kBPBmGHow64zp+beE2puaYsAamzmc2k6FAljowBr+B6r3fGr7cT+
184dZNSlDuphogombzBPJ2EnAb1LPJ2xh1hLFlHZ9A9HX6RUmMzy9OPpmWbG2TZigiM/gOgTwo3S
ZZv0pXOBuDWq4YdWqWgs1eDtPbuERXYqKysob3x2bYxAUVlHcDsWwadXfDwhLKpDlDtLyk72IHf8
JXfVe0L4924tz2qW5GeiciHR/IMzQIV+3UvNydhdPzK06RX/HK0tczD2jzhHkCqGfUTp/+SYP8ia
06GW/HJWi1VGhMX8rB+ZzQDf/saHCrvjv7pqaSgWev7OUZavw2iYl4jcRMIj2kce8nmrbH2v58q2
rsBi6hOybTNQh7kwNDGcpYaTurn+fTJy0+y+uu1J92o1GpFAVKhCBJMLvccGj5Ze4Hbq0T9umGQh
9zAOF/2DT0iAU34T7zL7KRcVcT9s8BA+A8mUWhq341SVcoy0kWBoBMXoxzujYkuVMzHOCMpejyfr
tMIaJQYTraBILoDkj6cdM6gqTqIqV68ub0xVBOpLYMqJunvILTs1Jx+VMylFUbnvTYHvBzyygl7/
ug8a+bcioljrSF8mXR8RxI2y4TOp/9cVacSldJmkLJ9eGy1/VuJ+a73ouKWhNfMPWNBriUGlcZb7
0k4OQMANOSUW00BYtHIKAJ4eQHTVWVHqXE3ibj3gxl8hIsrGqcekpKfYTvpxATE07ynrYfRLdgvs
oP1N/D1sbNP/xmPqPzH+UlLu0smAsGnFrRgyqsLp6AfndeX8CLaH5ggGkgpBv0iOsiDEjlAiNxI3
axbFN5RFthXdEGEN9ROqVfg06jMJEzyA8KLViRli+YNoKOFjmT2qrjVKDd3QGEpBoOs+zhI7qS6c
ZsHK7MhF1EpNhZMEtaok/shi5lfQ4kK0G9Ek1CqIQfMh1DykCcZedfLURPZxb92VTtmFEI5r/Fhv
qeM6RMP+qpF2F1Cz15qJRDAKKjw8e4Uyq5ZaSbZE/NQMg5WhvxWUGncipRQoUsUd0Yt+daZHKxbA
MxqOvaq/rsDV2q8XV+tEIxnBPrl9MxINZf8jnSRLzF15ztW1ZMqlqXZF/QxTm5SL/3oallC4199A
YD5DyIlVuFKX53tZ7/iJas3Mv658snU1+CoKwlGwoDe1eWOLs1ZNpSLmg5Nq42E5YzHialjU3Z7z
GBUvQxSpw7AmSI7fAvviIv3LCmt52TUJfjras0I6jikHF34E51r8z5fBvTXzHTjbJDDZqV0Ps8hI
fVcRWaKPxmXmduPqGReSRdEdX5FMvgcXYCJxYdy+mdzI72UPLNaCkjhXOv7lJRpOoRfVG5GRn4jC
k173V0Vi+syO1kAbFXI8+TpjTVhsfr+0lw2icEWmvtlfXl6pJR698bl7/w+tonSrmRFcJRd2i7S9
jFUlCQM5xk+cU94ZRdRxNRCiHjJEohBYKLIcqbMkR5UYDjFvSnYr2+jqEG8pLEJTy0iZkx42sNCL
4doBrNh/NzjCLEgozU4lVMWjLqJujktCDuCYRoGE4+Akc9AeAmPaefW9KV2YM7YbMbw6YdFgLCvx
QW5SOLRlsyOzDvFewcfLimmlCGQ/Qj6NBTP9i5A/qVxBfwUhuk0OVvxaKHWhVpZDzGxOL3xKQvQT
FYqi5h7lNJZcfujXEqx3w4WF8aJXx+XoIMSF2m5S8dOfzQXcNxfGGTlGrZ0nb3M3J4xt+8ttxlWC
whaLepjxcPVGixOyThGUjvPrH7qqoqmXrV1c37+sKf1TSxx2KzjLikKfBqAg19qQeqD6VdZAuiC8
lLIdi47aM7TGYGNY6nxKvvvry4dcFLX/KyWilOw3ozem5nIUIPmZtjwx3av6fBerlJVPL8g+CTYj
te4M/M1Z4jLHAoYsY8Q9o6RmBss6ythxDKcBgQv8YiKundsxG93dD7PR+w1+FK7IRsUjwDstMhSm
ElFwRalqXw2hXVg9E9F9CCdQgMtl61jOeKOPYYU9WIZ/0pHzYp4Qry07xPSR20cA5qRgX7T5xeZ9
6VivQRaS2T8X+putFfHKNeeSZ9IgyKG4hL+a0qj4sH3s5Zb/6/XOkdmFVjgCAMcy952NLHphWz52
dB6ovibo8uvv0xjMgv9dAkqfI2tsmjKZqXuFiHYjWOftLrQS3Fi17UAIN18OsqZP8Tpjiyw5ZoiY
dNl6oE5f6OYtKpTtBl/99Q7la2QOlHk/ZV4rV0TPQjmKtVtvo2uAsQIAFwIQZxlvX+9HRLQBrG3Z
Oby5QL15wlz+4yvnlyLgy+LBSZbmfYjLNAAY40TzoAMkC27FVgc6prC+e5FskK8p8oPK8KejIAsA
pWkQD7be5Rc4ip1QpeCaTK8LDQVh71r+CRYjAHNozN5BhU6Se2qYU/L8Z4c1RC6f5+E+j8rZmsRN
hN14IpvIcU8qfLksNX/cq2Nktw6UPOdXuRf9S8Yiq+PD9iI2aHP80OPYfWv0pW5umGJJuvRpLifI
8HRUyjW8eiUi0ouzF93K24pLU8raMlJJhyYcvcKPWDeLGMxo8XjQFZvsMJRwtL06TDI4q8+auJKK
qGKoJ9twiEtNpRyrjWRjrFg6Rd2eitTgOGLnXGvU90kMGCBD1PXPEnqD4vfGgkPi/dPIgomqgSLN
YhlsA54xY+B9lr3POv7uvyYn4dJ0QZPpGdBQ1JEh5IjCfK+qy4qMzCohQB9Kd0KoG1BvicaMleW5
K8fSfDvgG1umdHUEga+7qRlzStkXHZY/dswj0xo9Xmg0oTLP8J+VLvx3zD84m5FogTsc3DG3iIRU
uYmV9K4OHYGXz/JoN2Aa8JMioZYOQ2QP7OCv9Ir4AbfePYV73657O8UyyWaUAn+9TsHAkn8F05nn
UX36NMT0f6KeNirPaKXbJQLs0stnNNBWTSmDICsiVyYd3Sgxm8lXWDrLlCXIdW9EgRqOCk1lV92S
eMrFfjEUiEosiq3EQwG1U7aKV597+k5zDg0XkFGqCLUayk5sn5+FZl7YCsnxt3lnZxLDcaZHAbss
6mc2B426g1q/fl0eygC+xTKqiC1+HBSbcRPNRSZg47TLPabsiE0MeJ8H+6Njut+A8EDlw6wXDq0m
GqL5ifvGZ7Bc7hbOT2g6ECppSgsDOlt4CZoAbMWe7h+GoFlNm6FlX6LQVLQQ84sCBo1a+f5mj1zK
mkrmEwYHY+f7/1n7s/Q83YhXMuZ4MVKicSB0zsaY+Z2KefWdGyH2aYqWyny/PAGV28wZpT3FNbp1
HRtydr/3EdNaKB3Ram2Z6AO5xhH3sLchNO0i8ZsmPnJRyes03X3/cxZXMdTt2PJg4CefdNuCRl9U
uaf4CZIpRuL21yrua1RT7inl0+EMKhpr2WZxAUvxJbdqs1Ye7lW1YO0tT+fYlHZkZVCDTAtb0XXt
+pP6mZn5rBwlW4Lts8TyXAHRKOOmNvFd3cUwyqmD9qmTtuPcmXTFWQ9+lv92a5KzhJu2kYG285Cb
sReI2DUbxcKq1AWUGu9R5ACPZUergaF3+74LcxAyyvE8z9TECppNiIW5FIed14UmViNc1Z35m0/A
dpmVsOU0lU2xNrI3ME+xtefy8hoysAtRtsKRsU17QSrnpCG5z8axX1r3cy/GZOzAwWqWUuqUp5N/
2QxSc/VX3wM1Ygnnh/j8iU9KOhSbOAszen/a1wcSDXLFAnV91OUbB5sGC1M8qLmVsF5GePLgFPsw
LJPPnhLIxqUP5YJ3sPzXMC+DXmLA+7tQWxuRhfvPbbfsJbeDEPT6ytDcf8E2Eojajbz9tERuLl8M
wz+d6RX+rHi3XaquI1Sxkphs12wEmbGk7poramK5BPT+t1MBb5OSescnbRxqQayv/3/fGwY9rvjS
f7Q0APiu//OBq8CL//IUKt/YQvGzEjt5vo0fe5Qgd5nYaG+2e50BsaALmOeiTIB8ERobL6qmdRZd
ld/CXoP+rhYeS2qsXc1eQdYE5ihT0Irwp0pmLaaoavIRDyqTxYb4fMSC61C28taFLD92GOOP7EtT
1FYcw8vUGvyrCaz3hWXWEh7jfvi9cQ5e8VBZ3rntxHsbaeLfeRm30RPQnAanOrbKCan8nLvezifx
vkiLqpvfbHWAM29ysDxpoA/m9jAqS6xTItyYWmc2Khaevgacq+U5ci8AXVqIOQp4gGDl+8WT9Qao
742DM9pFLrknqHXplzBuaXZRoDbv+8cxN+ZqeVwwt0wdDNYm/eVkcfeD1vy1zeLnKvP5JsK/VBbu
f6xEvli6459yK8z5wLYykHSnTajrwfk8jAv1WN9DLziWWBPSgESC1V5Cl+ubNHf7cPXMkHf0DbjW
yrgWsbrUc1LVgYrNby9MAL2C/k79geOSc1EI3P6eyTwuYjf9l/fGLVpiz+MTK7lX+P5C4WbqSwQx
PNZMbCb3ZOqyMv8YbRENzLHojKv/cCs0h00CabdfkBh9I+bePlh7CqKt/EvTgc/ihLWjSeFRg07j
CWMWurLVpF5O2ZiA8e20ozX0uONZHNgpctEpmZjSxBBTeEMSi1r9hd1ZJs1FKk260JOqLPTWjMrK
06pCkG/Ww7UkZ1d2vk0+IZaM9hd7axRsdkmfPau4l96H8C4L8LtfH65wWB6JnZKoktFdxZANP8nJ
h8DklJnFaS5hn3i7LjP43AejfOqlAvQ4RHpx8FxcVcgPXS4VWnK9Sbf2TvvUact/KOIDWOvS9eS3
qAkS6neqbHdcIuPw1hvY5W7s1Ju3jDNYa7cPajrkTeTyN2+SewaPjSL7VEsAzlSV11dgEscGQB+7
nj92AuaHzmW5Gl2qsbQxnw2/gpLh1fSBoCs96Ov0HNKaq0PJmOrhp+3bMrPdG08WV7zLJs0me3HZ
+h4tEr9xi8z12Q9nXYj+KBfEgNzVAgPiNtXOLYLEp5ORbEGwJwgmbk3o5lef/qoCbM19iBGsoGce
hSoY95pWfU9buE69XM47ydbN+WS3EMJwESqq1kKjRWXzyJlnntZeCH6nP99geoBJ7Jolzb67ME+C
RmMnThCeUVAgfYJDUzKSn5cz6ngdcIE1b/7EF6yk6rrC0b65SWiT67gC6nPlk3ZWlNDcfPtOJKqN
/wjfhegbbiX89Vq8NUY35vu1otQZDzbCBPt91zvlTr52cA9QulMiXsDbVQY/qj0wsIRNbf7sDal/
UpNRgQ+v2GSYXAhCxX71DPY1DvX/I2wYVsqnAog8dg44k8gJ8K6gBSM/V7bSxWg9OJpWIvYND0aS
41eWEAM0yl8hhPkOhR5iYPG1rVQ+ABs0zGzAoizytzo2l+5tN1YLnKGh5LA2tHDb/RT9Nv7K5O8z
JMZhO3ngqlPL1YpjUySjh0pR2bmbdhkUjZyRzqiAknIG7NlxJziJ6xBABxCwMpaJ9aSSg2ePrZR9
+1e35vkV3VFknDK0Z1Zouj21Cqug0CGxiM1lb8kulquGj3lkHThjaOroPjSkctEh4sr1oq98/gH0
SJGJasAI/Zq7zX+GkWBG/vfEyiQNkAx02n8BkIU74T3MF/I5fvyN9m/QxD6nMY2PqVJsiO/LMKJQ
hlsAxsUk20VNuvcJrJjlDu3+ML5agMNKKW9r49ln9jmPcbDpY6glaeTxQ1H0jNcBZFr2YrVFMfmU
iPLL4hV7jsZlboWdCwaig+E40q5xSqy5R6fwrWhDdjR/QXWcMfjNErly00HDQqE7GKba630BCal/
QeJ2QPZ014nSz/uJno3zWaeX5woxaVTFT5za6C65qAkC+T78dr2yisD87vzgXB2vRVUdXGLKJuZG
kEnLBqX0mXJ+dcCV7O3CndCqr61H8ABBV9ml5gCpSajIBbyG5f0NMl2odFWWXK4B4tScXpVcWZBf
2925vSecmWs5a44Et9j8zt18uIVwhAsk8mOZdS+FOG39NrmtnDDgQ6yFzSTXbb3uz335Z8Y1cwwE
RRG6I1l5BEIvMF8cMtc+Oqj0gOcTpkRosviLUNp+W/1H6oNuS04NVJn5+6rSEUIR1s5Tr7fUdk5x
yW8ZElOutOFHER1vFcr9j7E4QIj9pgwNRqFYCLAAcXNsg+V1cPFqz7G78nT78Ml2iArCNVxruYPf
j1WV58AlmO7lS1eha+7XpWtJM4FrEjwOkvzPzPttOA4d+bv0ZBjpiup4FgWXIO2glZjbdfbCnaVz
vObR2VG3ajQLvJA6xEJo6DR2PeciOPs9mFdt316nZ8RSeLAJ0L41bmf8qmNifI4fiqf/NTwa7r+D
+rXy1f/E8BDmHpS3FaMYdQjtY0+z/ESyYlqkczRqmMNchgg3UZxyRG4O5usFDhAJ21PUcn2Mou5w
ZO2hJdrorzO1XtTnIYe0lAWDqn9kWd0L6Hkuq7cwSZ4Cbk0ar6gPhb0JyxCoONbQmklSnc7Ikz3I
5SMafhZU09ml69RLOAysrX2kFldRg6hRe1K4mAcwxUBmuukFEt5vqgz4Jz5veYBtUzgnMgTH5mOc
g7+EHGEF0hIi/Kir9A27KTMbjYKcBXuahdOYv+O4Qc7PSslbMg89WeUjozHkUoAxX+RWXp/z/SXP
MFemrxo4H8339JsxGZ+cWlYcGOPnXC9vupFZQ7QORGcvhy0Lse6tis/hGZWIZFYx+T+MYMgp/3Fz
v2Z1IeIIYuUT7se1ffwJcOryjmceaDtW97u3yHy5YWpP2xAqSLyxDbQdtQfq6rZHeCKKRA52nXVO
rgOFiLUFG2dN7/qOXgKi9P5w8t1GQ5ZIwKC1aB280NLRkwQxu49JRmYuu9TfB2Mz3IKC5xj5eRZF
EmlQ7+Dpb4BHMIFGNK7D5C2QjMw8n9Uq9zj/YdCfri7IRJRFs0dTGXYsAh4wxmnlfSDVaRvRUYDS
BeIMvnt7I4yVjvzantvhnFOeEyoELj7XsPiHogxN0Y295ALmdjaP0ixoLzsGkITtaPv+qsSUWzPh
H0rPm5GML/L2O2zgl3i67G/m5EQNBS3jxmRU+OU9zQzB89SB1pTYebxtG05ApHibGvTRBY6LgAHJ
sS+r/1dIc56P6dQTKi6NcTbCpuXzdZIVY5ecGFWcI54wt07vQRCJ8mGsQLvEwmsBAu8Syzlh1p+j
SQ7WKlTRqcOZJQgFSHblcVa2tgBMCBQpAFjIL0F2BEdv7uX+fl1U9/qPBaiQi7dwJxjSyA75cGL7
Z/dxf5qQtML+o5RTi28ibZkW4/W8qm8fCuJQi+Xy1lgZPz2zAR5hTkZb7ESLywMQHE9rbAvKy1ce
5f3YqSLButVwCmHk0F2R7bTohq7EcSxRWR1hmUnG4PcqVaTTB7F821KD4Lhc5mdgkErr0UM52RON
LVvdLiCHSDKA3tmpEnTw/YQe760PqSnYyLEa3AObq7HXf2XRiDfEE7gp1KXWbJgtrYC3C2I8obhL
llAiOqqL044NSTVw/VVcwBkFd3I+6s8eowxrESazwiKzBWFY2jOJGStZsoZxMYOqHcw1mC3tB9Bc
30WpCmRWV1cwiHN4hOf3i3xOiN//UuNvD+m3lnB1JPecf8SyF++rVNh2nUAAsmBkYz/7HDdLSV4p
4dtcpETQ1o0VKvFpmPjZK1p5d0bnr0P/+8sdWVrEtTK6H6EqWouHy9yH3g3cYto+ByA2MFI37Mq+
wcBwfeSHEr2r2FuvVO/io1ghp6siAWoceng5Tyqcb71UbVaQP2sFMZw8oJjMZGGbx906YNjY73Uy
NBdAirw5yXYRLNqzgV/acZtbuhs0SJ8tttwWLM8wfsTrdr/4qBWvn2O3swL50ZGY/AtoChvU4PmU
qunApfRt224EhtNH0yjgLWse7x92kaxf2h6kUbPreY905q9FHUofRq0pIE898V5zvww1nK+FQCuP
lZAEC/jYVW1PL4UaSR1RF7pxAaHdz6Mbjdq5mghOvaoIND5J1wR8VlgEiVqG53HTkNbvW/DJT1mL
SP4zvMsRX920oDwplnPbAe6ClvY5E15kutgAG0umVSwMRVWqVfMEvwswbpjDgA7I+uQ9mIrAgEBg
rw7aeF0rcS8ZyQm0PhPMFwxBIA66MD4MFDpr77iouw/X+r6fwVJqmzPBe6jHy5gW3N4ewTdofnUV
ysLPhoNyTapmtQMoBZ11fF4INfKfu98ZB82ica1HZA5sKlAjBD4pEjcfNsN0HfVfnI1bKbY26U5L
jUiAe/hA/rv/EFn2bf7ebi0NTcPTKrGiFPEXSGKmbmvxku3HOpzeeO+m3UASyL76JysT9tdYmMwD
vIhAhXr2Soa2wkFNYkTqnKiO8GDdohaLx/PWL9+JutlH0FtBfwEZRdhDULtwJ7dXw3k/nj2DkcoA
4llDmqq6/ncQBNkdbGAXqBmAuDLZ2V6BS88qT643P1dVzEtqx8yhG2teywKElZshLRPhnRfGOkH6
0auEowv/WXFVzgT2QSgkg0XMS4g9fir/pjdXryvKB7XbO4LaX8D/BImBMMsHmoF/Mpy/NbNOJb1X
oH7Q7XDAQ0FFfzBmj9Jryy12boPEpQe1J7AwIe1i1gximu+8RiDN+lC2VhBlQeoafUoBZmFPL6yW
eXp2+VTipdACJNwL38DJWme+HNciTn09wvw50wBYCXmS1742Hh5tbvgJadGJHTZhxfjD5ynmU8jQ
kzo2vEZRh/3n+Ie1P2YrHtIEQAeMKQVGGe3JiXZitszESsvcThI1+Epc2NZdrzZs/b8es0NK2wWS
SHnCYcgZaosiQj5W7xPbbbFD414k9+C5aHZK3PEVGVDaCfWJG3s/xZsyCStBSyNTB+7VllbK8gw8
a0SbAE60u5PNGWHBpI1s6FtDHAaPRQ80MxG91585kHfdNScrErObtjAbblIFZOFR5W18XaZi59IN
GgJB0k0mrFA9WqdYPAKg3G0Ukfzp5vRZudOtNUPAWfwMHnnkZ8RgEMErt/3cQBiUfOSPvoAiAYYR
+YND/KTGkg6ym9B0EhzG/mXNZFfXzZpRSBhyqxt8EArTq+FsMCpQXCosxGNKg35i1ARpraY6mZAb
9uFF13DbfCxxZHYbYBX2lt/UXuIlQUtvEu1xuSeqLgp9ExwuexEyylr/GuAtpFHrcx2gXIAAZMsZ
Jvewxd5FLxRy74hgkzpi0aP1qd/GUowpPgtnDpNTnpJd/MHJb7wIrdiNJ1MqygsSRMqvMIgduZ8p
P+e/wNYhrHSUgb5BF07u9+wOMLWZT+8pjDlxmLM1tMr+Sc8ZvjFuYrYBErLNwnOnEmwMo+faxhmf
aGYcup2Oqa8yKl1U/OVP6X+el5Bv/Ke6g7yR2OdUzBeqM8QxNWZLu3B23773WyGxicrBOjcH9lAS
W28zA8u2+T+FyhGVqVqDLkz2Euw+QEyzXKKn/TQtDVCrkXVr3DA1E0VIh0Okpn07uxQK12fcTnKd
FBD72RPCNdoL4xmsZE0fYqzA0HMSJXmN9IUKkVIjRJhGzUEx44oF9QZlkNj++X9O1bJwxNKR+imt
5ST+QqUjxN2aka8DqQVjkH6YmWwAv/i3jEcOYG4++PkzVY+wEyr15UsAlvPQsF/FJr2v+TuRFr8F
ZvKD2oeawkoKv7CLoAQPpxqw8nCvjbUJrOjD+iq0xDiGdqFth91bcX27pEIokDCPBjsoBegvxAtc
XsLeoS3oGCtAru2YxCn9ZUb/sBg0N7bmhJzvb5NQ1LrT5TfxCqGHARzLpYNYWD0F6MW0eF6kpixd
JBFIZDlq3xosRdRd5BVUBk1er5vqdFHUlYTCWnwo1vxNndbld6g8lTEGtxUbspBRqFJIq6Rifunr
z7n7Y7SkXoavaMkns18sVX6spfwRYy4pn/8n93KpFQQtgOSSB8e9lN1mQXbmSnX6UsK3tBxwOeWb
012/0SSkPvZ+rfdgeouJAavVuVIg1wDzMmZ1OpXqMUAYvN7VnaF+iLZ3QdB1dZ21yYWWqzkjH3ZH
y1Re324hQyDJTcEYsXAMK5GqIaI0aHuLSeX2tH/T6ovmgmrKxSZZLjSE7pfaZhH48VfmKJ4u+BIE
jRRcIp5MZQ7CyY0RkEtwVRzzA4h5TaTbKGtWdmJJaBaiDA2KbwoZVhyQX7nxX9XN5mulUrZ9599+
p4HSJIHE4u/vN3zVdRFFql52mEqVL3eJ6sQV0o1afkDbGANkDgiH4tHrWQpQeKhOZzAX2f9LDnrW
OwWASfLxA606p1BtyUIWGgUHd22ql153OxUU2IwNNn5r1cqOH2Gz6/6UPiDMj4+y5kTIwqRbQzZR
Ya4JF2vW//QtZS5Mfmb7I4ncahv0l/iQlAtnFkANeHvso6jG/q2sRcYzC/t1U1SdbRpjmR/zatdZ
E+wS4fYBt02xcAZM4IHpggX9MbThAflPlIQvHHGm6CvNCz6Flw6E7I/AVHj/J/vXjpkv3cU/dUIr
rZoZ3yHTHp5/hsMxfhKO8V9UA9SWKb1lQWzqI/9z5xPmc5doZz14OWZm0xq5WLcrCpfa3WDQ1RTT
QeHtEx8gjFHjVsPmVE97D4FUrZliMIYmXMhOknDc4nDaBw/WXT4lc4rumivqZin+XwvP6No2QLcT
QGWAifx6o6OUdC2/jcj0Xh8q5SyKidGBHY43IisPoxfxQuI3dxbFDXDEdDXZuwHqAuyuQgnuJBLY
OThl0sGixAWiKmFI7gy44V5aCbLMDddFRPcVRY/Nnto1kIPWeiKcNk37oULDjEXclH0G7MFyY+1X
iKAONfuLuY35ggFbU50u3QS6OK85W8r+Bu0hNqPtMuPWTJvOC44TY5uFLcRvW9QmiRI2hiVdyKoT
3/0MX4CQGp3WkTzjCm6wMpqgNsyKb6sX6dXwX0+RKSTLYm7CS71XqAKU2SkVkFM/T1JwhW90XsFb
P2P8XCjdZ++0szoSum6+fIlpVJzqGMNJlgt5N56+JR6TxHBscJ+dn5xJq0xDkPbd7W8jBi+y/4eM
5iRnMLnSu1dlQNbMzEAdWSj1GqKRJQL1HcEshOkmk8kLwLkQvJ4sTFAN0I/Rs1niZT9yRTJSxFET
maIPpsKKSHqbfRsKIjj5sqV6CkeiIJLfw45uQoKdxahQCNwMeOcmEUDbb7h+Jvv+a7Et8ADzobpH
GdJOEvmdouXyoyElHPVJYfCY/SzR5uy7BgietZTVGL3F2XlUID6CbPYaB0lt7l6zgMC/APLS2O+a
Xwp/MoqCbYvbgayr7trI+EgoC1kaEVxVDcRd6xEFGBvk1tSfd8WOl9+0ciLXdave7DX9+0urUGuZ
UlUVnEdAKxpKQ5LNErsrgfRwjhQ1ryN/A6l0lwlmzt6vzCnlWVdxkmGrV/GSFHdoIx2idkVPk4Ds
Ez8iCdI6bgTlRMw6e1hxjZNhGpnVKGMI5E3mBousEbeDbrJy7Fzfi4/deizX6jXtpuvZ0Bj69r/C
YIU4qke95TAuYcHIBPYrxIjVAnLH2GtvHMgtul8H7bJxuFMPQnHRDFB3S1zuWpf6ZQHXRQBGty4m
xxVE5bgb+RCa+zYiR2RdLnDmjzj97BxqOHD0ukPGqqmnGnMOJHiH6ke1N34KunyFrQlueQR827BM
gP57XGR0lfrs41JqPPxzRlepKCU15gvt9ig0hmgzcT8eTUgsXQuCCsTJ+yhDM02GWCIBZm9T/EPs
/t0oS6s3gQqOUigXur6MVIPRLMgSXuzH+0CWv/99qf4Fod0WbVRXSL931GnBa2mUiBDUqBSqFHcZ
sDT1weS0bd81SgC74uBqyYoKL6Q9lop3WsdyZLvqgPn/sWjFpRdrPLd0lhwCt8dHS8itgpmoverk
z8s81SHU0MVrujNCYlo59MuvQgYzwBrLaeFvKRDmBYWoUBhu5a8t6QW36Yzxa5DB7BfrurpydarO
HrU2eH3r1EspVZLn4L18bx2CNKt1PgBDIaXBaQdBdy/yeRiFnUJe7Rfs8571SkwdkQ8cA+J77ybU
ASKKsDQdZjr+Rn7SehCxMRkPUbqOJ4KcyaydH410NQHspS1K/1GmqH4ZzAwTc7ld+gQFDXoZwy7H
jIDYIZNC22GIClK9nlk52kYt4kYYZKwy70pWLIWgAIgSFWuT2v3HY/NLLkG5IKc/TOE3qjyqgcKk
nIrN4YPcxLvny8TxG2Z62RTO6C33U7vsMpmqqbsRWVoYWyKF78vS8HRJwgMSYwpw/iaZl1k4egZ4
zOhcY/ryIAMZ2/Ce+ZGu/9noP1SdHfPcfkJhECImfTNxf+fenLMu+BsVuXUWAfhU5xfeX8xP3Fa0
3TGsVWZ0Z3yHCxNtGw0vuNEqJa8PcJZ/mHbvBj1zypIVcKKwTJOFYP//PRwr1KfX9oqYzIM63ZIW
PK+vCeAmolifmUZDv0p96enFX5ElZnuUM+HfbYqvKQR+8dgMoK/oEWPD/I3mn5k7diKF3cHHvofH
EzuE57QlPief3JwxSQHGRAZeNDT7ht+ikxDj+Ea7M2Be7VYwx1TFgcHizbdXhqvkr96PDy/aqQPf
mrJl+c1PhuZa9haYtIhbKc25+kbAf0L19j/9paddg/gvKU+PgisyEFtIT9ehG7k3OtzvhDwX1ea4
ukTLJq1HZK/hfy7hy/PSweeBVBBTYtuEbf9ALIr3wArQd76KOrceLOEXN/AbASO87IXvFXsNRCCM
/XoY6GeO+76xVBlykRH1nt8eeaWE0t0JvVCG80UPqyHqD8lkBC/1E86wyWgk0zj6tBGYyaIBOVZr
iuwqHO62thCmzgtbcRnT+Wqv1SgXFtcy/BaNB7axuOntvj6a29Th4zBnA6XiFi5NnEAdhCG/MSi2
cTILCRPomGItU0aRbXeBdpoQ7ScG70fztF2UapdHMPbyLCuObPJQQUrv74+fXWBnHdt+9a5Ccp7M
POwse4ezsaBChetRqT7Om6BQZpbSI08ipX1fnt93s4fQXNC6lBHGv0O2o7fCZCVg2tviE8yEm+CS
RyHT+kA9Iy1VjMwmRCrUkGLeMlzCRA3azFjJxnxcTMBIAFKeLRpxFN9Gohi41MHzOSoBqKp8YrAb
tyN3bAlMjillvuCTzygAxskehQ/klqrt/427lCNjUywwQhNR9rdQtHdlZZ3mdvv2af+rvpeQpTg2
wcNL838Qw1TbWMSh90Rqeo8/9kONCTdSx/UGtJ+HNXu1qfvzdqAgVnb3NNK/91BGpMV6YO2MtOZC
WsI/TnTVDNyCMELORUfKoLLbMYMhYONJ/klKh/XO4TyvvfNawTdLbqeKzugA67J6J71W3qnyoVxU
JSM5NAj/RwWneO7669fxck2x3VhTnENR/JcFuyYV2gIW2tK5k7K4JCX+U6Os0jlboZbM11RWmmOq
DLWvPtaejessQBFw/YS0tIo3jQBH9pc/jdVQi4CUB6YufZav6rlC/aEKH+lut9nk7nR15zYyn8Jn
FZLCZ2QKWzocpXHWSezu3cLNPWesu3AwEQ2WWPwkV3TBZ+aK4i79a5sqMPAtw68DBVwNgSjGWmhD
2bWv3XcMLi3QnVx02/gflKHNHQBqhoBpJygIJ1G2GuuD3Jinigo55p6uzeowth8cX4HB1PGHe1fY
QRRIYupsavM6MZzKk/71Wt7wOYcwIPBOh7CCZUpNe5ijbaHPgWht1PsVdCD4bhdxZQvnNJ+9lczX
SNrQzI0zn1JKBJwaLkzUrvaP33p0/1w0OuenctM1qUqUFA8L014s+77YWAhQNJRNZQxtDBITHEK6
5eyw3Gr9IlCyhqQCWqTdq2gOCzUSPI4SlaH5cylY2SG4bq0G12X5W3+OKIiQMErsuj1k72sbHp8g
MY1luqn2RXyxUjZRuLSFX8bzAbtoDDcPEkMmHdeLTIRGlAQibawa2N1fot0G5165YLy7g2uJb9SI
huja5PifPUaHfEqx52cnmMQWudO6HFij9eL3478tkKnDrsu8ythF7d9F8TmFpISSujMr2HewyiDN
2yYjfm6F1aIfgna5oqw47up6+KrbeZqJ9TfaeaOK8iEb0JXZPskWZmn3TIR9r3JRA90U8/1rrvb+
ApVQK2cMJb00aarTVjfodIHT516jtoadwrZpXEQr2KLT5/FlClXpUkWYIS2UWeVzJvHRqmUlr8JM
JI5gaE1a1sZ7l37agWjVATbDqAPqyy4rWMt2bqy+s6ljKvwV9v38cs1fEVL5MKP8mMPr9I5fRNcI
UlybFr3nMmo9chS1GD67kmTKULucXl1iiyw2bgwCsGOWizcom7todVFetWD8tofBDXTksNXaAznA
NuxtRf+Q7OrQTYTFGvS921g9hhvV6uiJrNkpB9QkfIY7bxrKVvvaeBzYvcTtLgvh8uaCWQ3DJ0ZR
kUu9OI1kcHDyM4pAdoQM6u2nXRCEZJo9gSVW3pAD4VBnJ+WG51PiFAeVspqn4UUvMedQ+iVF11JY
oT4w+4lz58MKbGvjR+X9SJCTVJuoWYcwJV4QHYF53BbxXKAXzdbLti1tkZmpbTZrntXHe+hGmUb9
rdgnDn7DauTKUX+soLytf2bPARcCAV9jeZOuDZVC+hC5ASDzy23BssCizq8hayetp3KAp6aCbrym
isit0BlmF8bfzkiaRcPAdonT4YyuSeRY/DQ+Dy2tIga9zNaez1x/i4OwdmaEnErFvVy5Knn6Jvrz
DhTu6SQhM3xOCGYniXQuvLurzT1BmHq+roJHFWpW85DWwtOqcj/DTZAoR3B42TTMOdcCfydrvlcw
I/FbnM+D501yUJPeimfWa3dnkR/n+f6S1pmf7WgRuhRzBddQDtPu9cnb84GJ8VUB+3uF+q97qTpf
17FRY9K6kbyQAB02QjFpB85SAY7sxgXWwvQ21zawbl4IunyCOAoHgMXZ8Z2r347mL8/t79Ii2mwl
aIKfKThhH15ltLqAyqTzHSyXQc1zelBjn5xA2Kwmqf3YElzvoyftqbiCfQ/gQed886Dq+qReCFCR
ktRqLW+SIZtg3o5+NljYc1kELWQrgGjP6SAFbiqPYgp3BBUGb2/EOHbgYQfJARS2m3JfYP9+i1tO
JhZf+WX31P9H810v7cTof/9w5oCx77NWY3kAEOxAhYRQCiNnNN9Wfyo09ii3qatw+ZOA4zAgCC3n
xBcs1smWYImuoefaQLn2kCZzpl2HIH26QypQLA4Hxl4OKh+A7RWbq7inVTtaHAyhfHJR8fTpwZ2I
o0eCB2HhQxlc1/yhSjDTeTtDrAMw7B7Q9UxgwEqZYLAn7aKokAaaCpt49K1yFStk/9ZedXF6j7zF
LV3upvLrnAtSwrR8tM7tlCDouZV2zfS2blLz7qrgRergEnhAYZLDd8qGf5OvPEwbNk8JCwHaS9CO
9XJYDfAozW57Mu5stMqvleWhOtwZDVqYrov+R/7Z/hUACR7y6sx7uEgr18LL5e6Q05yc0bvM8z8U
OERdSHghF7+pm5lDEiokWs/S2fHp8Oxa5e/vOMbQoP8fgblXdmJZqqkelC4LzcNkUUFtrKWa2dQJ
9tr9bLwtAAyleGOTCs7UqVRPTd6E4EiHVovDjC2kXCjpoCCTwFDFt7gaD0HBIUOctInmO+OP4e1k
Yeq/VSMgIs2aK55IKYab2bLRR0uLlAvBY6Om3LjAEjvYiuJHIR7qbKJNybPLuwSaacZ3m+VgPxVZ
R5ZVCq5/GHOHPJbHo7LCtnrrKxSgsGWGADzcVNGYKAQANKLBeSnG+1hSntK3Eo7uzgRXC89PMFXt
2xhPYy4UMc1lTa4VXfkMdcGEK72vFbnIITzHEZXDyVcWDd89ovFS/2am71zi/aeHpfaxnm/ptTjH
HSghWxtMMxPmy+Y4EnM3i0JUaiX1/gvhcftP46cxRj3ZKa1Qw+4AF7cDyyc8Q9erqm8/r6D9XtKq
xUHtKRK05mtwUWQH3lsiibxe1Txxn3RZhb7+LRQel5GZH9uKrBEyWooyV/albuMs30DyY5w+oYNG
9TSaZb1TQbWAlkwOuohjp9ctw2cP+YLMVF1+EgSEiqY1rX1dJd9Gu7YadPZvxAsunN2nVeXJVj5k
dBv4qvliJ8BaoVg0ORvh2d7dtldr0VDRdqPD5Zc9QmWvmk8erMyB6FasBHOVLt7YU/1KGomiKfso
r4vyNYe9FcezZGFmx9MVIkLd4uJYVoF7pVXrGJYbL57mlwgEwOnvLIY6yjfxFaqnjju8ZCuRYIHS
0BM4gYDJNV5A45F7M45SBdBnw1naNN5DJhxZHlLKvjv1COnA+KwshDjWsNnWbtT5/N/5X6nvgwQ1
jIh90j9YjkcEjTk9MWr0wA1e1OPbPBPRaeE1u6R7hq9AJudvLRcr2CORoGQ8ZPlzcUau91pKXK6H
ZW4sqRKJcsHr6ynzZEuY80VTLU6FDdiropaMlrkTFHkRI2bpIfkbMkU5rLXUdnzyz8G/o9aXf5qO
l6a/MfVjzMCs5vMFNglxwyPpri/eW7Wp70HizIXxQelA92VFhzth7ME3HMM2zJ/tPYjzQYch69KU
K0ll8UN5mgjXaBzF/0oqzoh9wU/Ena2+/0evTf88WIj0BYctbax/LQw1JH6X0G3/TSorbXTwxXZ2
Gi782K2f2cWlCMeSGiQpCjm03WjvdHZHI0ygBB8KDzJW1jGulEsY9HK9LJiSkkFbpNPNRTqJRgdi
AIPSNk2O2u0pSIssILeWHt7y7RlXO8RPibIgHHr0AN8km0JMusZRzCF3A3YdqCdw3uykeOWzqgUX
dFfJ9xxyyAjT1DX73wqa1AFIl7mJwzEvqPWdpP5F1iu8MD8+9v3z2eFN9LY8wK1dYmReWaPQupT8
8znvZ/GshTJizpcRNQIdSWcd/PjjS6BvBRORt1p48d3V9njbZP24FHvYz2CGfTJ5v5/8R15sjICp
vfRK5Dt5LT5vhaNmOSfwc9bJurozwIc0U7D7LmLd8rO7HNPs1whgctApNV+akJZSXUzNyDSTGpXT
ZCoTn4HGFUN6lKuPopmJ3rjddwi12uF4Fj2Rsl0IPRmUl7A7+sW1PaCNr798FuYYIEiRZ+xfNEjo
TpkEYtAkPKDzJMZbAgeue1hVojUev+hCa1uXKb/3CMaiOYR5obvNAESyfnEKoMbbIaLy9gr6zUHJ
FjC/eC23ZcVzb0+1WaE0EklhWYgvZwkE5BLtmQk2DYBKiIcPhVuHTbqUTuB1nWE5mr7jylpCg+zJ
jQz9D4kvTE6WHkUZ55865bHLP5uaGO/X4OzDpwnUFAnkXpvYMgWJ3sRVHxFyKLLqeS0Q5dDFSZQ6
Gq5HuLRRm3c6mgWfFhspgKVdD98mnC82iQ5K2ZL5OBWkpHOSsWstRywO1Y4Pohyrd+eVRY7CYJZj
/afZls11jEw5QX0kfOBGdh6sQZGyY5/oSMI01evJkkQZZMfTB/82rdoGQFZwFGG1deoXR61Ov/iy
EXJjPLYMzdMnFyaICuhWelEmZeC6t+uebMM2TEkVCGPQeRLSUO9Ib2QWsHL+stTnSy1lU9/y6IQa
woOUSI3GSQi4DI6BUXK8V0peV6vJeBuDqfwzDzOWcPbOQLvYNid+4wxI1wi/Iwd+gGdZ+YTfxdfQ
vUmHEy4WWAfEhjrZ2XKr/z+Qotjr5y9SKx707WHVi0P9scKoRNkapI1XbBanYTfUgCVGzPI4c8h7
Au56jGBU+P0tA8l4g/bN4BZ/IvBsl+BoBXt2+5QMAXOhcXBxDV8sFj+Ng6Av4+Fy2GTcAH8eGBYo
HPwTbSBR15pIy1mz/cDW1JNoIp9BMdi18qTVQlAfaH1n8YzfStx6JpuESdi+4X02Ha1xzLdpYbF7
IPXR1snAettDxST85jC1FIIsg9Cw6MHROfk4NBI35E5FC0wCy0e6UTqEqUXMgYkegqjWaSOeZRFx
sm4dz8B9/95HTWRGQuk6dpg9cHWKdEYiFnQc+8BYdUECwIRvqat8VXSJA+ZwFuAidxg8NJQAwnf4
QFs4BK8OSpYYO3E8g7iAbSi89B4rpGAqFbKChSEXiw2RXq7iP43+sKb5jQ+dkW6GcpRXDJhEnUa3
BsoIRqxVAlxUru0PUOzN5w2voW99i44jQDwgctCkGsMoGSkhVCsJFFfW/lF8M/tIxAYIncYwdHbP
MLrSsb/w0KsMkgADrxsvsQLrZ3LihlYtQ0oY9HLdwgADQgZE9VRzDD5hUNipizHJqx3RDBE6mhr3
/9sQElCtBQ5PSrbWSV9h3A8jfdUUsHHBV41kxpv1q2XKSKsUoVEn36C8/S8yokTUjQ6mZkd/6sAx
UDWREAR668zCL2zKUp2PMSw8j3MXcUxVBtr1fhcPH3ZJ/5aqTBRpU6VVPSfnLbmE0jcDhy5cLtSC
/58ATbR/RX/LSp6aHgV07jYWfWI/mBI8vk+srVB0P4U4jwWIdLP9XqSRz3bMIaffgmnOf7qKoA7L
MG1FDHlCL+u8zsOK7/N4Ud9I8iEV7p1buRdulc1pimD9RKaVAYNc6O6NhbjOyfUJkiw1TFdiLibm
mTdg51aubNLP5y09R55KPOw+t8Eta94LT0SR8hcAWpacWm0lHkErindLOXGflHb9tETgw8EXvEoh
GZRMXP8AkEpkRFc7oOhg9o/pj/mfA2uZQ5SKHt2/mXr/Z+O4nzAK4gcIk8P4GLmjMb0AS+dlLLdj
uunkdvfVhhHV8ZGDXw/qVxhHfWDO7sSxZj4J3gse39koa4rXEBRO4MT1mPyuCPEvk7zIZwallGh9
2CbR8yhvtn7LDSV1GZLe6G0qtiAKIXACHr4HBDFzP+F3Cl7dyc+nm1k6KvOHYwtlNb5HLfRLVC9b
WnpvuC7EaSG5C+xwo/+fBYNvvkDmtDf06TkUXyq50SKtU08zNUeOvmY2tQuyO8bR1I77iWFkCb8Q
f8laAVP+T9wnt+vqaHIipTmiQBPU3dW1t/x9Mr3KyjYACV4AqHr79NoKhnHR47d3hzWGP0lc6t4A
CMcVDI/NUsqTqFd+92xsaPG8yQXByCFUBt8/0iWxydWUWW+tzVOUu9gLxFE4b/zq01PgyLDTjY7B
5YMMFUqLCc5dsCxbmEUvkHCS/ktNtvIJVxkkX+KBxkGnmseI4G5myBIkVxwOjTNBmrm73+0yacij
u9IpRD6dJi93kQVyRW0Y1hWMXrRN+mnls+SV7YMR5bRkEZ5SR3X0ec1nnNKAz051nVluntl+nodh
Hcxcs/7ueYr2zjuNsbjjQMG8HZMyx3lEQtZqdMdHMxTKgO1lNQNDVUOVu6OpZTf7mJqjWhaW4JnJ
9BL/vRixdsBIQlTQILUBdJ4A2CqLL+MJj7UeVRr9mL2JttYFBuiA7pPRw5axhZqOmJopvYct61pX
43puh6zray6S645o+dnxGQXyNjeO4/0vEAIbdjM/0uPOjaWdfzeRKhIhGZyZpGbEcCuX2y2GBROv
K+m7kDVnfB92djlYjdosI9VAziusRohsazB9KXroFYqkPfmiXPCEqc4UNwfqIv2gLKli9yLeIcD9
bofG8TFlb01OP8CnRE3RTywJai79rkLePCHvHzmRI1azAHRylRNw8687pgjjSP45QpI4aASj0bTv
sY30z2nl4s5QJSWDnyoB1bKE+d61k1XppJgA0qb/QGEZJxJUG14g5JkobpPKMjWEcT71hld3djl2
GjI4iPHXxUyN+VlWuSoknB6kXFHmgT2wT6Nk4GCN4BmMhfDM0qhcYW2mh0oJ95nGQwGNmsxRyJ92
+HJJ18awpJesoHIJ5mTMrO5D3WA4h1+P/Fl31tSRDcSguBT14FYrT7MGOmx5OnK6qBsdBME2jUe0
Do56tqEoeo2Vhc9zHvleffqpXmg56/i6oDX1WfnZz/3lbODNyao6ruC3OI+E44zuJkW0uGKtUnBV
Op5O/C+Xjq1zhrgWe1E4p46PCwKXBEpU0Z4OKeDL2iYvOrUUtqUk20EwMmBRgeCE+oSQtZYb+XbP
uek2PV/ouErXLFYmQ1CVdkws+79D84kNH9UduivuYbovp1uCY/YB64Gbx2rIM3u/JRIfM/GTvpWj
zBvP5KD+pn/0GCMjfCviSQPgZoIg/W101bulEGHnBy5X3xcmIa3U0EEWKlzFy4H4+xypBMmfIQss
18LooUA8y5Erq7wfKZ27Af2Mc08cEKIGYc+HoBKtPEz+5aanUr6cJmhjpg2XWkYheDCfO05YyCxc
JtykrXpFiFdBAafFL0AhA0hiGYVcESV+lTYG7McHw/IzQrFcRm03OWHeaHoLBtU4Uno/573csMkV
tUsdMjX9iqUlljiYAClYJsWkV9+Brg7lgG2iASwgCP2Zo7ZVHUu4arApnsKQHbi4r4Bmj26xkzzp
pnv4gmfE9j4BThKEnEoZ9refS1XC3hOxgryKpEJCWaHjxRNOO7eGeiTkufH3sKmPhWLjccEZ64DN
XWl2fvaaMktmfOGqj4vQpQ4U+vbelO1YkOr3KVR23J24xuQ/ueTqThFFI8EiFzYVZsWlWjI+QKfr
/011NbkdXZOd+jh775YcP4z9fw9OPzrgQRAKmylMeGASmtRP9LtH5jlIccLpaC7LFluizCMsXHnp
kJKVcNowG85RYeQzuvkHohGzV+ehA+S/IZ8hH1BA7kTFmU3tvjlu5WwRnKLZzcHw/pT7f875dL+o
NiOA5MhQwodIdMZ0HWfOu+TTZlFRmu+lhb7SFuu3K9NnG+Z6PSC/gzwQBjbawUuKdHLkpn3zBWrl
ua2W9DTsUvaHPYJDFEAm4QrRHYjnLCuXJG0tKr2Frl6HUVs0jeGgxuD4jtzPXz9YMNM0NZwkLw/S
LuVvpaUEuupfSK8mjfWehuj7A3VsvDCo0esZvZdT5BtAsHjpQDcfrptekZMFhk+HJAxEquU+Z4Eh
90pfO2M2XlwdHHm6uqcM34dimpdRV+Ocu+n1s/Z4vaT3SQobVqhRHVkiFcE+U0Sx72H+6llIGiYD
pbkx8NCTlimqcZP1S+mnr0p/sqSPPH2N7eWT5e54gHxOJ74Injvra4AvawTNwjvDsRhyQyy/7yfm
tbkLKiDAmeTSxQ6911xtwh2gcJZPPTvHSvo6iHg2f5y2ecCwWnIlmiTeBAOznFFIhR1vJicFh9Dg
9Q6zblI1GJLjsLFIK9To9Yw2o1FVzvBSGstTJ6q8YKvBBRnhpS7rifaVzakpdbdQCusnBVMN60Am
FYZlWD3YSnnu3VDT1XMij5wY4xGpOkWC8xBnqgWhud76JgiYqFTnf4QxXu6bhF1Czmu2wUFX03dA
rDL9/pBSLvQ5jhE7Fum5zqNwbtmxM7cVIwmYlleoIvGrV9qkSU+/Cw6c6BTtHRq02bKaI+BK6rpn
/+e/HXpQKOG42IDWM1UrKdk8DvRU/jIShYxHqcGAhKwNC05bI2fyp3bTWGDSA2Z876WjpFJa80T4
T80f8oMoYXMG+C6Cv7sh2VWpMTHENSG5O2rPmAK3hgW2xv6e9lOgFGJp1FurRbZn7VmoCz3JcwBY
evimhtrezirh/NwTE3hhnKTVO95iTyirhWTNnBMh0+hPSQTdaLSzJb2ySVqufp4Uffz7WD9n0O4/
piyWXE22d1QI+ksXV25rX3+SjUibd9rWp5L/IXBQ8t/AJ7z+/I8UMtMipjh2hpcCwfXzl+cAbqwQ
pNfnvvGtuuS7KQtsw/MZSSAOd3ByOcGg1gs703VuOEXwwTDgPcLTf1k0AVXl/Z9V6vKbvRKBHnMw
RAy0Yi9IBK40gbeP4Xdj2xTYK1IE/KG/0MYkg05CxPYMQgm0U93KPMb9mqHnnO2FDonsmL40JcwY
JqVrtZSDYpF1m0C+H7uFQ/0TyuNWubxuODFz/2cyT1/f0LsJswstZv8omuxRKlfPkVt3ysOXRdDm
ZDIuFSJJ0xTzNPA711FbbtTp1kCxVJzMTgIeRhIMCTbdK4ShliMjGp1aK8svLtgKaW6ud8ZFBP+f
R3Qy9JWl1qm799RZixxowDo6G4rr+1lTHHjyF2UzGwfqJJyhEPo0l4gztMjlEoafQG7ULxd5E1U2
WhxQVowfR3QIYnBeUJJ3L/uNYogLWz2XIN3gmXpTgbloviEcZ+v8yKTdDWE24MnfBvV4OcY71hGN
yMyrpY57gbijzz6//NgakoZsih+fSKIwaLMTkoVdZsAnVirCZUpxuwXZPr/rdlMZUf5dcNXIqaIu
9v5GkKqbKjrCq9BfYVzvSZ88ltwp1dOSkrCzr89OKNpM1sfnZljSY2QQAfYxQnR4l3crvNFDRgv+
SRTbs49SYlVvuVmxuAhHngJSxNF9b1wbCZ2LDVs9oxUJmPvbCxZ3VOHiTgj6Lh95WRMSI5QXzveG
a4p6EkK1Jz/VHE0tiSGEoaypSjioxofn5hw86iYZtNSkLvHavzItZbgfjmS+15aO0c0E83K2fBd3
XXCIufDPEcbebwcab9Lo9lHoWsT0nDf78417t5b7+S/IE4mQWR2u+XLYx/lJZshDiuUVBeRBrm4O
VIoVAXFbmQ8khlzvLnszWZMgPL6kqZk8CNm6bvlK1NpULGOgF5+pgvy0zZDLqAOjjrM9kWUoCYN8
xy1kUTOMYUI4AlHizAXsY3pVf1qUaxSbs2HBXLZ/6kX1uwQUrooQMQLOjlLRZ/+wbOuGn/mF7IeN
GhXSGoQMQGXQ7fILiPy2VptALALuoSe0lqAbnjACw+49wNvvnAQ8/2rSzqX2ETmq2AS60VaxWK28
aKH0T037TUfi8YukXjuQHfr5GYYmUvR0yarfVPMj7vg6gRbGPRO/aHM1b36cZvpqN1e8Rv3xNZO7
okDh/MzNcDuZ8qlDiL0eunRWgfPY1th1EbzgmShguiPSSaxjBOjIL6OlJ9QolOmAOWXB+Ju9nYXZ
/R6At3Cb4i9+53N5Uns8iaNjeToK4bXCE90LQF+JtDrMcbJaWyhjhgJdHz3LGGemyV6BKUcZ2C/g
w2UfsJ/wHsag4yKG2ZOnznLv1o2gBxUs8TpQBrmnU4FukARqCLCMU9gRAb+tLyZ7YBPc/U8HQAuW
idRfa6TjFk+SWbZY9t51EUxj6p0WSG3hJzLbbiIUoEs0SAKfe5rCvI8T+wGHKE6EF05Vham6kpXl
zfzYJq4L06iPfp0aAnAKzMyuR1Jc2YDkMYvtLUiKK5NZYzhz5j5d8WkWckHB9Vil5CNdGEfBvdSP
6uiXx/IVQEJ9z6pz+ruuTpd+CTRhW1WVrwvdcuAIGNVQ5E6Oi2yMY5x1Y6JRm0o0VRE44g32pEZB
VvZcTp2pQch9EZLG0Fhxai1b9uKisakOHPS34Si3BxvgxVkw1xddFdMOm3EMtF2ai6dWoehOGKfn
BwZK3etUHNrApUQN7AKjm/DRuPmZZP1iArYj1zOz3VdOtmVTKhr4zZfeHcb30oSEt/FGMNTjJ6kf
B1iCF2k8gYLcWv8/npL2UVfgVzJpHs3EsXDkt9rB96iOuqIeFQ2c0Ah6aa4FqEaMXY1T5soybltA
G+OH9G2nKUqWTNh2v1NgbF/6vQ8VNdDG1sZPRuT/Ivr3xIYCVrRb+XMKp9eMyEKn0aQ3WSWChnVp
RvAs2yOlNq8oW+jRz1O2a/SWPsLTRU6+EzHRiapfXkvPkV/8JN6KFTbSw/IVXj3chDgZsKuPlE6R
RgL85kdW8JHWozk8R1S16/17W7vTHJdVXUxphzsGgf5oECbiLs2Pu6SG0BPkXMUI/c3V8cTMBuve
BeQCBSn1tI9gL88E25Z/s0vHpTYu8h3PmoUQckJ1cn+7HuOk4sld6rYuUx85Nm6p6sniy9zQGHKP
Zb0gCtw5eg7LaKVDdHGM3eYIMgeP+0aTohlpqeoARL0Q2JJmbnnKXzaq8Sg5zFOakFIyr6CRcylA
uL1fVxI7m5Sjfkh9hwXxxzl/4k2xMg9+EwCAhFbHLEU1JTIJK1vljH1Y4Xknu/cz6pcwpfBVfz/v
RkV6nGHIjXH2mDcDTNzsfQIFnjUb4Wjf1Og+sTqTn9ytwtzvhPK4GH10haEw2ydAuarsgWd9st0/
DEeW8j73+KezXm7xcHYmPPEw3vuabFulXTF3oXm5D+jdxgXnmJziTDSWbUxWRgEvYGm+yr0BxH9X
hYxUEsHYuTSHBCiOba9P2DPrQRrKWLtixGmWrhEjQ6mxrNweTadPgyrBuifQzptVHytPP2+H+MwA
C0/I4nUPKCvGuxubozVuImtPN3tu2g4p5S7m8VetksYV/kzSb648AGf5wtfv4IDZYsjMyaJIhmy3
/HFaPD05sV8684pay1J6oMu5LusEBmX3pam6weux3Xcq4CycI/zV4A7F3LwkLz/PdNEwtHLrKLK4
zTOvdH33uPMcfezZ9eKfnuU3AVgOphBLY3xhrC/SXT72iMoizVnX7v7EYgZ2C69ZkzNY+wbX4EEn
GHktb6KAMWAmMw5w37r3MexO5Xi3SDGkYR2schIG0PZC/446OeshDcZBUc7/LH7Kv16TxdAVlTQ0
taHUUSE5waWTwxdIr5CXj5L7sWi1B2wTkxaMITV6+VXLldT7rNmHJC6B2S+Zov8Ov1ahKqSsEYSN
Y+3PPNm+58beIuGZUW71YzW1SlkRrQbtZuHevj8oezWjkw9ZqmphgpVJoPSZC2qXaiX5FbvALIX1
3ZkLDFyahcV9HTqtfu7AylPhKtR2oyszLyNyEyoLI7785sMiykYbH0AoZWjKzdrbMOXI3T/lghnJ
QGeHUe9YWvELbGy48PIuoI9Opfk75BkqhKOJfXmRQg4fKGZXW4MaT3ZXg/tvGQp7uFv9QN4QbiHY
QDAKBUZ+63UVIlZKkveyLPOBQvInOmW0MWHu/+40ZUt4wlOXm0pYLEr/KE29OICqpvWNcFl72H7n
+jXFrxFg8sV1mrqauSVgR4E+gaJlwiNvh9MyOqhuJ2KKpqV6MKMKIC3hd7Jd3MHxiOJvPb8Qsb3S
ti5Wh3lD1UdzE9uUaxujOOVkA0NMf3eQuWsLuJKi7vnEXRdF30PyiI/K4qBh9weMdGn+b9ZSec16
lbPudwJ5k/sNFhmXtIjOffmqAZcl/NHjrt5yoPzoTZBmjjCrlzzXK6TdKeDK1ee1oqC0Nna0JsD1
fqDHl4SM5BgfjJ0ZIYLj9w4ggGrmr2xoLlKWSt0WbpulAg/0sfvtJe7gKem5BFgMxbJehG56LFAa
L04EkutiUnNsjegyVe7QHLgLagmaQLC2za4kHqf9AI8/76Yu6Cog81oznneaN3lRP4BqZqv7SMRz
q6hI7mGX0w+58xwAplOzbd5BNK/fFjoQCY20Eun3kg0w7G6sFmTAasGB37mjPHrDVd/vpG7oB1Mm
tgrKtrG2BquDiW7RCa92tM0IoccWINwKD2YOF1cfPaYyXLk13HYw3MY+Y/jhpvZc13v0PPJgaYEo
X2Uqq70C6zmo0nerxCMo2yx/Cjt8t/tWlo5PN9euVvn7FcvnjQMbhA4G69gy8Jh5CVG1ccy2a+WO
qXRh6e9Ww3gc3p3iXI9sMMJFA+jaJJu1WsfOb+7jLp5dPZfta8vOwZVwPBi9yMqPQ9axbFQ1xSwM
7ejiC+OhZ3Ynw+7fIurNZyxcJj1Jq2Kld/0RT0jo/zaumG8AqEUDqoKbIjntUtkb9Ywy6C+5lKQ4
Pm9JL6fXZIyEZgOsfJmJoi1xWMTLQQ4/B775wWczWKySVlS+d1n2cn1w2ZLYksiEOXncgvfSspyY
m87F/hx4VbnqPhDeLg2OLifhoVUxzV1Watr7XL21nhBBJJND2rKxD6zhh8jW+0lNUVL6czhj27Wo
iP6Qg0HSaANeAFF4ZXeI1UYe0/1Ve9Dle1k5BVhqpK6kzfNI17WqmEID+O6MEA8u26ntJXc5dwDF
rtE073qhaHXn3ZSRZ2QAeX3a879HsadvgoIdA2UIB267KBKxrzjL3c09tTtJQJxJdWHUtGtAxkox
Vv+5Dvcrj5rRqB87WYBK0Iac4tje3U7D8VRLT2kfu+Jn5FToIp0eDE+7tGBmcZkJIgnnv3BQG52K
HiCOzIVEQoYXSd0/6wB8lWOLwnAbEOdMJEuuABh97PeRzdNWk74Ef6Rs2L6OC8GMWOabiU4wmX6V
EIuB4SvCqZkavPmbo6l5b/Yq0bHlB3tijLZhNWeihx6FoqPGJol3HsZVG/zcRulr9reA0vlS3r4n
/Op/6rZmH9DwAMZ3GSochzebC0yXmzLPUemOmgv7DJ1YuEfopu1fRPXjHNZPjjvt3hTXjmVH/BiH
WwhUJkorkkyKU6xnnZMJlqh6UJkmdK6cTNsRyIy6SIr7KPnGciiVBL82ML+nCUqGUGWpEdMjj24u
O24Q1EO4fwovWZWhLJWXHVZiuKKDgPRndzmV02j+IjBE3czmrCUjWIoL/NxeiMSwdNdwsQYx3VlU
XjpIcMh3njUqvL/KxbA0vTBJAN3fk2UBt4sp55aXd/f83NZGhT9a/mAPGcVAo1SRiQ0uRu1NZukn
oEmHAG3Isqhgoyek4bu8MGUyJSz/R5XI9f5cZpR6BHyMSr4sYVJolK5fxWg4GX+GQeT0LXXBRUJw
ZwQUSWKriyxccRkyyyjtPgNhG+6xoZVBNkuEBottNYKm7ak42Y8cwEs7yIeoZDst/gcecllf4H/b
DOdlO+Lcb7rsZQVtZvHqz2HK6oXpT4Qs42Z5C+BN61XH++nY6C6wYgVXGuGHtkXduYAEU48R8zdr
SJgv0ob7uRgMdLyUNlzPVHguMzPf34VSjX4BOZ+k4+QZ5caDgxziT8qrgvE529lDJMm8k7Pjei1c
xvkjTSYYl0Lj3vgH4agix/OPb5qe99O69Kuqy5dPsbXVURJ/ftrn3+DsDni8zN/grWziw0xg3uZl
4lqHTWL2UOe1Y4kAa5KQU4zoRJ9rGzfVEkpFLV8oknGnG7ou07PcdXHCsUvIDtcITpeOQOfEsNBG
Bb5cKfIi8SonJ2U9NLYUuPa0OAxQe1awJPq7LiTdr5fm0kVOHDzFVhrz6eL+NrX0k/FUwEZOI2e2
WP5lG6ygBy2Wmyz69Tam4XN9sgF5R7WsfvRIBkeLXjc9Q9Kl/LWna55ucabgItcDKf6m1L1q7L2m
/yOaZTwQQpQegDNNswvNR5AR9ZYIe1uDV8wQ5uqPn5NmKIPbSkzpyJWodXWz3YCOuPinj/ve3NS2
AWo3UKffY70ms4CsgSBqyx7Q6YlmGBKv1UmPZJWqs18QlNx6WvxcYWJ98HWEOIPKbmFhdLqgTVuB
plhKE2eWaiNF2/X0DLUt2MpHZzBf1VkD6yJVX8+E94GmDOfovjdEjJfxhwfTMhrJTGbsR1UbhsoE
VF2bpe6iVBLqHdUuq8QAy1IYqRbupv3cjV99TPi0MDmAP8cWzHhxBO3BE5ITENnNqgLEYrOMMByV
mFcE1B8tpJfvZWwNlJqr5pK+/scfD4xeQOf2zFtiQupLRETdIOYpbpRcRBAAMljqbWnZpg/WOPcz
M3nJUc4kJ3pRWjNDicr8ZDG3Sa0hBn/Fkh2RyP4SxzJ4waNwD+plPlRt59GxJRjmuIYZB6DlNRsh
HLExhdwgHOhxU7h60YC6Jc7hBvvZn5SSiZjSVKr1KvbqFnOs5HcAcYddRizhiNkn66qxTGNh7hOS
e9k2wXm/X8bK4NwiLHbsiQpyvbNaazI4+JUssL2T0hncRhBmRYYsn9lewNrEAOmlqhcn3393F3sM
rcsmKssYS5F/jmGe6iudz8g+ZtdJVzBiaOIXyJjeATQa0Bdt1lOIhseQWvQUEf4AVGmgyNt8P5aB
fQUz67eqDXsQZBhO5s9VjQ2YBD/2ZcCWfm04ZFJjoWdqxLCQ/NBs7vVgPuNcl3ZWdJtz3rqcJRD+
BV+Lp/1ExT0/wVQvJ7JDSw1XMqTsitOzCSKbNvittCCDwMqmdpH1gGHAvLEP1DdDeRFamUbW5uqa
xgFtSnmXoUB5N1zh3xnXAP4XhQJBYXUQaJ1B+O/nFZImB2M61xyOSdCUQSl9mBc9lCnFhXVzTmV+
Wx9zcl6amToCNPwaCaJcsoiQzMwmymqtByDiV+bggwwzs5tUPoY5PDyfA9PjrFFEWNx/RxpVrJhR
NGF34+nr0X31D5yn028rxAiuroJBf006XZNWpSalpbikCp8aMpUjEH3ufsly1oVpr8iR+z2H6RZT
TVf72QscJDHbQ1xTP05o6s42Buh4Rzi4QjlG4bfu/srVWFvX5D848noQPEUQhWASBXg5MlvD0UH7
OkjlyJZmJHN8fV3PPGzvmU2Vb5cwwdhs5pt/OSSurQuz0/48WbG+eJ9VuXG4rIMxcwQFiSvSb/Qf
GKIOBNMXPoZhSASMhyfIcHUJFzfwIMEc3c6CN2eP6fc1ihvAC85O4jpoOrQ3fw3QzloL6R/Ukgsy
a9os948Mk5OoqZfNFFxtlLSD6OkIGvvf4yokpgmFAdcLzHcsXqoZnPWeue1sTE+88qaQTekjN2uU
VOBUa3QcwDo9L9FeXomekLNHJYHqiTVdrYOch5IHzXAFmvnQOo70ZI7RR1E5r1FUXu0qybHbfAkd
JDwZfeENqxNkPWm4gyV/TKptcLU4B601hmwVlzlLEYl5yFmUKUa06OGiaGihSySe1bt+iQfXY6w+
TRYTLi6cuKDE9c5oVkM/9sT4FOLVEVsA+QY0CgXzDLSQ/6+hVHstZqfHZYDZOxwaNylCXkNFeNLe
CigJMU39KibjbdlJR2KuOZjeztt0HTsXqA4FB2ta1CtlYxJBI5XhCbH3JVRQlNGh4DMZGrcJ1wag
MtRQMkrK1WSF4aAT3tjqdttxe2ge19suc8dDG8/iSwRwtXGL4LCTuy+sXz7uUxksnBY1yXu3qPFP
yRi5Wm87i0H+1vm96mOLlSbK8EDfKzT0WxVyapVJhM00DlPGUM72l6MlyFdYUjzFpwEkBct4Og+O
nFeZf7c3zXvb0Z2WViXW/rXR/t1w5eldTbGfgCM0b6t0c+8TZZ9rFA60vJmiwS+mi+JCXnzyg1qn
i5lOFx5pY8UJdWdA1dUnz85FvA3Cwuh9l92okQq7xFIUhumgM0j9ETZ3Nz9J28WbSOHfmU9qShK5
qJdH8vugiUnGYfVsmW6Tsi/lEFgI/eTl88H3hTG+2sVaQrOzvGlZX88lENc8J38uQw4pVNxvNluW
y2hPI/diAYE0hpZyGXnZWOZmD/8mOE5pCuOuI/pD7G3fJfULI1+eCiqVJ8zD4/Lii3ygjz44frpO
tLm7leKRtzVeASWq43Ca/99F1hmbDdSkQ1PiTpaFwXWqQ7r2MmSn4a5U/opO7ANwOkrYW7zcDdQM
J1acidUEkpeUfMkHQBis70qHch/AbfIh/hQoqgy5MumzB1ZwaLdKpOLzf+mkedNUi3nEQMNKzGKw
nq5dkwXRz2j82CMRhvUL0uIuLsBl4TM7onGAapkvL08mhLRXpjlSBua2apYNUvGhIm5M7hDmjjIi
SETPobWikmGkP/BWOTY4c8oArZ1qm4dvSqHidKx9q6SthMhTUU8L+MIQPayZTq285DpaB39JEjlS
RjG8rfbwiNcDTbqPRm7fj9ger4hS0lqKsFMsLHrjVWpoAmkD7N3q+Jmm9e1VT+o7ai2ZTKJziAss
UpE9zf9TiSQ/X1P5MDRlBSDJ6+pNkGBIGVavtNL1rewgKKjNvVurkVWwptD9/SKjemCO0RqxclwW
P+2iylgn9+yVw+QdvHCuInMvKYt1x1BP6Jg1Zsp17XeEjaj1zaNPmh+BBf1it+8YyVJjDilBM5NT
2OhurhHa7kIg3bRmZguxXP20vimTs36Hq+LmXxxnhpA6Y+Vwm3KH4aOSb7frx/TwuatEXaxI8f1D
NcbVRyB78pJjxALcOPu9fLq8vuHKokS7QGSBIQKjLbeAl+AATeD6SxpCFWNZRO/Ru239OznJBVFB
TmCbT8H5M28K9mIkbixfyhSXWmcaVTno7BrRal0FrLX5ch0eCaDsn84ZWnN2KeF4OLqpeSwI0Hp7
gtx2imY8UNkG5TG9bIufzeStZfqGHOH7NWSFYQUNiVderiYwZ9r13sqpTaU8JIkJx1IvpvZmqRxn
VAtYG5kkQUFmAo5ppRd35HFcdN5SnWVPcFwfCMZcbrTPOhAph1nsnkgMtHOiURSQZhCQJp/HHYj+
6LlQWG39zxXJMDIwJ9fOqnGchU+LLcIU2tfQLW9MbOqLAH8F7Pycomj0E+guSR0XlNXT092FMj3j
8+C7VbovCgzrsNJUT3O+iXSsNN/AJQnzvsPYQr9Cz5yeU4n/nQPQrj0zmo2Yj/toX+hsBzkDoiFP
pCd7ZQu1d50b3n12zKPO8ZeAI/y1kCYYrCatsuSGfSPJI7hZB+VDn5iGKOPDhStQgvwBUHRuNTSJ
l6+TVAOG9qq85YWWiWxMazX0qDkko2gJuVl2cVX2FaQlmvUCAXWLbVjbqXDvV3x/flYPMb0Veq9o
euJ1nNP8/GrqTxmKf9NjKryVqNl5t5xrmc2WD4kBPh0X4A3mfgG7BYiE5VJrEzuPR8nrekwBZznZ
/TSi5hiybdWQMoxaseD33QhqTj2D06ewiJcAimykItVHchgTolFpTZgACTwTAvNebxbcV+mzhyqX
xmSnY2zgKOse1QBnYLEwVgHGwEmD8NOVVeRwoF9imeFbGkfns4n7n92iIPvikAqooYMzKt4uAHLl
Lg5TN13jUUwwEgJPry/B+kGaf1BeUqRM8jcpUJnCuI3mLDCwzhxy4KY9WLQEncpJtu/QvpmTV7h+
r1qJxrcttAPZeOU6fpWRD3ZTLmre9Lb8EkRk1kgIQH+HY6X+y1dWtVgV5w8rKv4BR2q6or2O4AGy
L3Zlu7QDkddI2ZKxkWcTyiw7LZ5aCF1QmHfMstSd8crQkUz0mpo5Do3qbWRdTZfU3Q4fs/0aKToF
TGW8zvI8x1LY5FVaT3Mlw+hPNmf93NfzDbJhOU/AeIJKclFI5p2OL4irc3fzgGxj+XY+Te5Dy9K8
HkcjJG2F8cEW4Y2FKuwZw6oLRDJuPPRhPKucmnvUQvtFRSElYV0qFXgQAd5VY5pVBbi/x4i/PXKr
VkgvTBqI8mG1sqOYiHuDm/knSc+qtooMBQA8kesnMBLpD82yyDd5rUwh9INOBOUfaEkTt6tdgK0D
59yrbPvE53a/CTfYkBCf/q/z09pECYlg4y3wM8F4LjAAuRFtUlOHrkmGg1fAA4HhTNw3k6wyxBpf
GgmK6ywztmt/bvWnNTB/LD3zlmBmo9Z8F6fDQICO0EiLF3WulbCLdZG8LPW5/TNLJmVXLHOcBmNb
Nn6Gx2/sh4IiaH7hYENwK0ZQZqhu7IYrI2+uPuLODFrgJFvgtVP0acc0rwxIM6Aolbe6wZ7DnTWm
f2dLDKH17yDjVYsujCbBR7g3EWyQ5bMp3Vnh4bmnkN1duPXy1Hn6IspbBHZ/bqJELtdlcCvV0qkB
XHyo7EzbhdctyuO6I/Q2l3+n5wI8WIHfptSPCoVAXAsSkNzu91GVXLctT6V0GExma8qxARnNye2Y
tH8bzS3ARdFwgdlmEMeIkzSyiRsPXs9qP72MxWjb2VZ+xX8hiHuiRkcPcEoKRdhyCucjLD5JzwXQ
K2azzky38kPmArvV50vqRARoC1HVGQRrsucinv9W374mBQ+OstzNEeVVkzWG610IPe9xBdFhpQlD
Ay/qNikWFiOhM8d8cDl97zHF3LlFzXIAmNmpN8hVok3aqh81U1qtWGjOzK39fXDPZVGsXJVaYpns
0F6RiEar9NnNRjDglB7sJAggp4q9Qj4ROZUedmRsgW6ZtToys1yNRo2Xa2mn2hOm9gkO+WwjBVSn
Yc8nW+WjmCfAm1m90trUjOdwDInJJm9PBGFGrvy1DaZ2QZjJad+/fXQqxQkXrFmcdYXbPYqPEZo8
pgotZ8F1LYJuL/ZG11Xsn+lJJw6YR5WXr3OyBosUN1Qe+BdJWYEP2w7UngpGrGqZqJrLa0cG38JV
kevfmgy/UazxUgG3u1r87+Z6VhqsAtMf+MJuM7jCt3X7le5lsf5L6MTIGirIbTxqnPcSVYQMDLdP
XtMR9EcHEOm9U97MsI5asnQ88ZnpfUQnhyzm1ORqeOwU9fgkxiJwF4obFX6D2F5Wtb9Y84y0QKCP
sp2ovQbdCXs4jFsXpZyoEw6u7S2Dvbug6cC/6zBrChmYsEl55oXtmbY9VPciYfvLTyx7Tfc6FKZ+
bvJls7FCYk752KDgDFYVJUSK+j/xw00doubWZ3bsYk4dmXr3ZeZqgGmeLq+sU9GpS1b7uAWo42gG
vMoxsHVOn2oH9eeYG+aEyK2XbtwrJosDZpL8jm+ih5q/iCWlW9tfxyhDBLMYr/6q4sG3uwsHLFIK
QQYK/C5M5xZwXdCxQbdPx5X6fex0nDbGh8EfkG+Gp+i0YJEvXZwB1CrUdDKc97g48iq2OZv3wlwl
x1ycXB08tkE9hVtST0qFkd/300QWrEcwCjHAcHkzvfGQbo8YZ43ozN9cJ4vbfC9fGDLZZkUw/efm
oXNp/niJ3T3eeXYSyKRFvrXGUbjFMS9uMXVlth5BfJI3o+40rwlJtj622kpQcsA37x/y3+brLoHi
6lwwFDJM9vOYBAPuHBMzlGMuihz1Qugwf2y0FUBXddkhaLzSuc4QME7sPFbBafgY343T8ujrapMC
pB91jq9X0/0v+dGLJKIHcYqLfEneWVdpSr0DBcZoXC8t0kq9qFdvN8GnHRbxdnwT9nXS/uENbUuP
6x4nKgWtMIGRTPcKq4/qdmICrb9z2NbuZcIh1AXjUT9R4zucI6vF0iw3OI/peIcsVrlZDqFfXxs0
bruo0geEq8b54soEGGPfvJqwk0T1hXjNFFOpda2rCLSfwfOHw2b7LZ3Mt2u0wEMKI395vJSE5ffT
l7k79+5ftc3FVRgCQpWY6a+bPvlQBrwQ8cvRxK6IMoBPZZ33hfbz4oUTmpQvTSCqKK+O9KArf5zl
MylKCHGDVU48ApCH1/wveS1ulhoYGubTXTA5IGR50+9+i9WyV0ue3FQ+0SMpGoGqZbMipMaHYJSK
YDJs17a1TLVyHx0FJpzRJi0ZiF8FZ0D8LTcGMo2rR48pEO9pK4rdJL7hW5poarxcHpzjd94NTkzm
PhWjCdOiD5sdTVTgNuhjyP6CjiEEJDsQ12mpQ1Ri3I0LS3qONGsB0TltjO+kwbSW62JqkupWVmXd
qdYGdjpTCVUkURtFwAzEOQX7+qrQtdTWUwzTBEnCG1+GZxKVSwa6K8H2ImK2hHSsNOHSe1lB72pa
jvaqdOc30i7iyyVrJa1yjcpbR3zOdCYKDNUDIIczp8GkUYAdY/eqtJQYo6DNlzQ252TGEsUnuc65
DJwWjkRef8tpSDBlj3VL2v/nHY/HVlEUtARyzyJSXmdqSamDD7Eg3qNLmLm43CYau2u+TOyoN89k
IfkT0Cw9IXAJErJe+hUHoq9YO5aWe6ph9tnYg8mIHn12S39jg5nFe9Tww/DDs44a+7FLUZ6Ku4bL
YWoKgteo1UXxJmbL/LwLN8S42Dg7QoeHV8eEmqZ5iICGiRGi/aF9F+VH5sVRZHKiNofCw+ON0ics
Hj5GaDO7nA1hm90IhE1U16rYU2ITKP9pL/4NcSHc7Rq9hzYd5c5meSNKZDovaVfasoHeMDec7JKk
wCRZG7Sv5czoO5YDDKADuq92JexMvgtMhvV27yi9/sNlADqH7oedKyT4cDycKSeaQ4RNcFFmCLcS
rm7c5SRqzFS0TfgVH1nO4agdMlrrCsSxDmXLaDxtMyJDoijxjcMyPBD+ApV+0cxo29fg5PjdLNQy
30207szBE32WeN6lHpFcn6AzU+cowTUlLM1q7whfB/ec/X4KSvSeWnCB6RcsPacryyZxKacY2vDI
8Nxw+MGrljAaDuX/8rRCTuTKRNWt0u/qUF5XTXH8zeovVbCYuF58lTLLPKnW9GcUqdMKflT/Kh2r
t6r3i4x4+BIrmUd0JCQbXqTDfO0ZUm0gZf2dmrysG3r/TnHIDZzyr+Yt6fU1ZfKMS0/xnoW30lxB
CgQUZGZjty5M8HcjUBwSCzSwg4e6q7vOPPS1edAcAt5UQbqefH7in8+KC/KNh6flEiRDBkHpNOEz
ST9N47bshyyjeAbYwuhhhl4BugbEHnimeL8PIDbcohB5HHujkfnOeluaGuEJ5q2+q1dC/+X/3LY9
MQyG1Pr7Na7IGyc6TI+oQ8r+bDoNgaEnKHVqYVfUsW+efR7tNzeTs55e3PN0l2OIg/ZbfnF4RXQj
jNEHmJOxXUrjOWIPXTlR0/vA9+LXBlF5qpxpLXxzrqby6/0/M+7AA956todJnvYQVDOEH0YYv9ZM
LbntV0RNj3TWROAo93vmAJGqci3eVYFhauKVz24/FhemL1qq5HciluxNA4/vHhqOqj5R+FfSmoG/
/lt61vfjcWvAGZ2XHGxCBQ/9riQLIfbK8kI4q2UKpSXO7lcQ+JjaFxLbGwj3XobRGX7UsZf0+yt6
WYNLeeWxSAcMHpzaODCp8pj8zhoh/CcfE4604GIyu/HtYkEqXu0/mfK4BsgxdgxWjcWkOgJIRZ4L
XElHV4vrQeEdSoSM74yKbp7BQFvJ2TYfEwvpEysDsNPC9dNWTkT9Xl+SOAGtgmL7DFUkitOCfEKH
VvbGpFAjcIMglnaFxDXYaNLEt7tvWh4EkVOI2iIGC1+T3UCvAr8F012aBLg+IfBxWOg0Sy7h0aYL
vC98xJtb4JtvPdgX8MUbEQGuSizeM4b0Q2SwufS+xjpUbeZpNuTk3FRTX9b70CU5u7XAytzsUaZq
mmW0ZfsY7uOk9luk1uPKpOr8jVT3UoZonaW8gr0i819CfzdfDmphtAvTl7a8B397HLeX30S+cml/
IM4MWUOugJYMxPyjuHAobTAR2j9WnJxJ2jgijm9ThXRQ3fVf9g34HYG3tSL2ZZP8GLKysPi+50aj
ewpY3x1oTSsV06YwCC5jTsaHxL8nvk1CMlGvWBjN/jOaIliXGRQ/ClhaIQIbbIbhLzrGZt7yGlqf
Fa2lQ1uy+sUdCpHDFCgYG+tnE1KLOvCqKF1PoyOetz5xYgAsGZLE48WpAqAus9Z4TWI2mSzaDmSK
/5HG2ck+RUJfdRt9+nomTdFfRRoOTMSZNzFh1GTQRoHBB0kv2tEUkmvjN2q6UeVkCwJGSDagVZl7
yB94nS1JR5Ft0JodIVucee4Cus/3ZjeQPufSaGvAZqccM4skhmQLPrY+QLpepV7yzXmDHh+YtgbT
fEMxUmXnw7123BUkcuF+JGcDKkSfcNwtm/tCCNALZa1hPUx574dsR4a4z/4f/lyrAdfGKOyWb7zJ
Wen8V8vxxuPa1E0CRUOncfizWnlVhfTumAvaTV7Ch5g+XIhvHQJVxCA0f7W8zEc96trn1odfh5he
ul+h7dw88m9HJ4dkiBHdUCwogmgegyJtKndi2Y315eOthXem9qhcfVz2PN6Ux1YA4RH/+IfKxvrO
yMAgdKjuxAdUfYUn6h3e1mx1uIw9KN7pUnDo89o/7dRW8UYS+q/js41E5n29qKtA4lnf4tD2Bjzx
p/nbOpzo5uVivtFgrv+OiIVv9tEYcjvMIx+SrpCkZ20bNRONwKlO7/JqaeVUx9XKvgIvw4sCj5ei
waG0P8b6nqau0Aua6UveRstigTu4C26e9Ajuij1S6KiFucN1p1Q4gtMHK0TK10bv2ZEd0GVVPk39
1ZDTVRsiL24C4PChuPI+NF9wIZSVhR4sBiF3Vv6/K+8L8o0NUTRyD9c9SzV52J+Sy1Jef2GQ4BDp
E2RgypcusqRRP4jHW0J7/sg1h+yDyZw3XbxN4/iVfGlCx3IBTBglaMjHi3VZgaQcGlc9kBeW5tCe
o6ZN0cyLVWzeIfQRJ+LoKK/kPr4wWkZKbeyrWVTV2uVc0jUFP03l1YA3biN6LDxcV0gM0kjOXQGX
9NoXKFh+Pazv5mjM8lJjPnFd8NzrLXZzEtq1533wlGcIpFgR0TWLdmj+zwGim+lTzzoSvIMwFD8h
EedKAjaA2qvEBz8SmB17crjmDWxshNu+WdQ1jRj5X3xDo3piWJqSz3RksSxvjAMB92VLPiUyHnsh
4iCeK9onww+jZ84wdQz/V3E1X5+1oucWCGzbqbc5SEKuR6bd8PG3EbPfExYPR+kED8AaFCK7Z07V
1gBqwVNOncvsQyXKHAv8HI1uzqSpWpyqy6EWb3ae0uimDXjzx9rdh/iuSQ0ibutjFR4mr4MbXqUP
/PYtyE1W7z6OFnS9cj602zCC+7kMeDZQdOTd8tufA6krkDfOQIjfUzVzYKOZk9/+l8SJCGe040xM
l03u8+u6a+dL5S4UTTu9cfsHnQDW43HViBeirXYcbDpi6usdt4S4gp3MqWaXsOj2eUs/L2bHOkbi
/u+Lk9JeFMhcpYd353UMNNrYeOAN2vPMFQfWARbTEgyVgckZfsCEbXxrG+uVkWYndcYmvvjdNqLQ
N0j9f4GGA9mdCulK3dwARMXxV3iWnN6FCoejBCnaY5bW8H4kbiO9umAJe7pzDi5H8VffWPJ38yo0
GDZt+o/u93EGC7sC59RsB2ilQEt9gWr+Sq2JRt1/noHkLXwFsCcSGz/Sd2VZvvX5Gie0N1fWW/MG
8lImFL0A5X1yzZ9ZdjZ44gLxq+l3GsAyjfvF2VNK3dalHSWAbAJouLBYujBZ7OLBFgqzqPF825vw
5y5GFwaIcMdsafXuqAtyoeHiqEe20Np1xykaB55I0MaZouQBm7zN2GIBhA7tP6tI79y221KTqhlX
wcHnNgBOd1lT3sLO2JV5v5GyWSUYRjSWqt4Pd7RNJ0t6G1+4ojR3PZSWjnMte0RjgiDcEugXMQ8Z
FdVS45VMtVflGd74wuvtKh/tLTIr1lxymSQf039bqq8USK0mTrgENjDangsAT1yRVInqOC+T3FIB
bwoUU/uLuPz2SwRnRvec4VBNM3kgx+Z692ME5Cx5EamgzNHDlhZRjiC61D9087LCjz6VS8UoL34I
/cmzHJ/izXywNvqHHCAgauLjnW5MU6QvXAHVi6FWQP1xUa8z4LXc+usx+YuyRSTA73bhJNW3k2Rj
mGvUYrenJA7R+51VvSJFK8L1Pqoq10vYe+yNyYNPBC5vbfjKA0O8ijiW02pZgq6DPXIPcI2qA6mF
OkJDgzG8c87+7siJ7Gu2MK0fq4UdRae5ZvlbT2b979NHsInep0IIPzHTxOTU4ZX74SEcrIRCtHbZ
478wyw9yn/ovOe74d23wAhfaSKr/PvZ/RRa9SwfIDPXnYpfJnZ4p73H/EeDB+TBs+97VqcUYSmNU
e5OQOifHJtuTZDS70CAymXe/XNEOp382gnzom93rt/8qgVJvvWWHlzABfoW//CssM0q94VOX+EhM
PjguzDPexlJOM35hrlAu81kyBq93/UQnlOxOxjc/5NTqRCRFl3XvWtJFVsK2eYIbbC+EO8uyniWK
J17ERrQvbOZChrk0cGcZTOstHb4oRBLlwBJacqjmUj3O68zn+VWAAclcH7sBQq+MyiL+i3ag6JyJ
hnPIWuh0LAK/H6vOrsazbvXJvF51OTQut9auzf2/2HGVFV7MRZrtACXHbEmsDCwHepNwg6Gyh06l
k3su4IZhf+eZUEXVlQS7yymyThZlmMj/CUxboJV7WHJHoHsbkfzrzprVAFXN3GIlE9zkrvVKMkYO
qhbz0FKB3J/ZTUEmFAUx6zRbh3SA0STQU19hjcAh/A2oyOIJGVaidsGZjDrsHDMub5+WVQH2gF95
cRx747bLhq2rNw/sTI13DoiQobVQygENsTb32xQZtjvDAC9qaBRGuhMJ8hLdl7YTXo5uE/G/Q4J5
PoP9BhUvke+Cvt2ubWyDLRF6+sejIJmXqPcGvFiA//8Vfld+JXitbsZpiJngCFLxkk2jI3qTSLn6
KtqdDzqfKLKaQcl6GA9l7S9nUIo1Gpu91t5IxhKuGkyEsSdM5f2QJt/UZf7dCOoay8B01ExcXBiO
rXr0GvwuM9NygvhRpgzpS4u3uMsHpHPWDoy6ojrDAyZkMm9meK/6EkRkOiPWwZQ6DT6VhScr2Oym
VTqQ/mG+A1O+0sJXVFxNLU184+PwE3NW9pEuMe2kYpHRAX7Rbq9T4x7hxhZ5Wx2OdBx1mFyh+pGj
B1UYqArpeg+COB26IH6+n54UldaaHrVi14XjtGgPSNLqUu0B9PyixTnbc6ZFMhW8r//KoOsFP4Mn
8lj3k4q1ybIYw/kMKEGAWHrbguckSJbBKxEM1riHIbUZGoitEqVe1XTpbBfN6USKMTOrIJm7ssZq
ShXQJsSLJGhg8zpjTM8haCtmziwfXb3vkj45Rpk+wLvvDks9B9M1F2fBGG8Pym0MRInHuddGJsxY
gRaBNhj5pMNCYS5d7YKMaxDlL3CKsrHREZC62mp6byUXwHR9SjofFk4Dub4IS3L9spXwueVU5JqD
mrusHpt3xTc4oO2EEG9V3+SVTI03Csqx4FYQ52WFVvym/1Z2YcWO0Dfa04efHNAYql5haJZ2nXh3
Qr6B3UGe86QiNHRJTIf9sWH8LYCuwPGvURbs5JAXlH3Ly2miVpiak05QmHsh8Agg+Za9YX/T1mBV
MZ4Pk5JHLeCVaQItET8rvy8ZpxQxGKj5R5PYDHPwnfnoF3B++CYNl8zFTx/jT6i8I3bA0NuHndEZ
hgDagyvpvpDVCxFwv9sVrJbTIsaN/mDHvv3+6usRsummSBcXuBp/dFgJa9yRxiGaeH1CrU+BsZ2U
J8Veq9xqXlAHY5wGu2oEUvnw+CoZor6xaidNa8mEP8bSHoDfojBb8fCnidl3bi+l0HVtx11FXSZe
4hl8MVBNx1c3DE9eb5D2tIlPrwtvsGbSc0ORBggCpd7vWRt0htuRbG2ek/ECjiibd+15KpM88d/e
wZlENn5lEUXEY6M9g8SJcvfsUA97F/GSpW8V3gf6pN+meB96emF5nw4EUgfn2jg67sGEHiRODVRI
UkuyXGfZBmkWuRs2549zCCKCH8S7puuujjnuVJvnUvPZKbj6LUqzzgdJN1z2En3q4uftt3m5plTs
ApIo4HXMSEv/B1NttRqa/qmQE0Gl3tle3lzCg1IbnXbIgcMWhDMzWsPXhHQvSyPzTslpezCC54VM
1zRtMZ4+2t4oN08JzdYgX0yrJ8mlRr4wB7gPzJPiV7I7G/s3oKYiFBJ2v7XWKKhk6aztdBvAD4lg
morqMW53dfmdrGnBEkC57pZafH5t03VXTxPqO1rHhCbGDh9bY7kiO7XklUBD/V8mBj/lMJV1b8rt
CS6r7+bs2tADjpw2jQ3O3Ec3JQGE5FbVlvEiwOdoA4g9KG8JJIE8tahK29HjJh7JWaDwiX8a8Zen
X+Ri3yuhwhuSz6Ed1XJpH3LJ4/37F15YxTau09MkcHXxq/AMqvnGldODotNGk89imhSVHKQmwnl5
2dYK6Q/UFFlAo8Jsy9mEKV7kV0OinA+pIl4TZChafoBKup9+g0WwmhS6/g/i71oYlsXgLGNt+C5y
fgtoKzq27ZvxwDH1QiJXlanTdQPdYQ/XzaNFnNdIjm56ixKtvgHuX9JQV+Zyy6Iyzj+uapg5uOUV
vGEICkjPFtlAsADJNl0EoQEyqKJc0rhTX9ioR0OiYpCbsPkjNprvOVIylxK+xM5XFEhHhJflHSkV
f0rA16Xwngm4d8vh5JcF4+/BYTFORFJQZWT5MX388SnlZEWMm7j432v6z81erJ+4ZvXMZnnBfdXt
E24H4kG66vJSNdVDs6g2ZCQ2Sbc6Vg94omlnNzcTmNGCZBjqNaM154NE9/1d5mYshTcDfPIGGqrf
+Xdf+zecTrn7TxJyr4LJPMfq03Nt++JQ9rQgHZZdfhx6CfDxMc3V8gVwUrgA6OQgsM4L35V7dEZZ
UYsVInv6aEBcr9k2kVNSRGa5+h3MkU0U7hzD/7Fz4ZIURiUkgKpeJNqERT/3YR/xjYdI5LiMqyjR
DDuTdp1QU9zZrpZZdDYTPtpFMkaTqHU3HnjbsiBhcC3zoEElEG7htyr4wjGsD16XJLWHIyEeRwFh
EBH+qh+5kCjtXt0GJDBlIzNw070TcMXAwdZ+lBhqimjHSEr+cYTaseYstXboTANm81ztViZ0d+8f
X5YhDekuna8834IsFrsBPfvK0peSk/aMF8rbIT4tIyjitN5lmB8gMx1qXF4T05xOooreqjavOvNV
Wea5wJdbDxIidOOAcPE0GQTqmgpR4pSGv6v97jtWAjfIl5SVaYV0ypTC2l/xDydkZrhf6tvkfapR
LRhoBTFKBySqJpJwgNmdzHT0pFEp6/1FTHThnlU1e1kI6MkpoCYdweNLWOybt3V2J1/GypRBy8+u
z4WkRmTP0R0dlgM28SBshXcy+P6Bo1R93FHoZaAxb+zWibyb6PH7KfV1DaVHRxvhTEyN1z0mw6wZ
fAAjmiXySaksIGQsroreCn/YiwWSr+YiGyKeKpMqRaaV04QdzJu7J6I+i/ZqDjIwxg4nmnBYB4bk
eBOhotukZuohNjeMTSETKG3m1es1j+iJG2OzLT5bCTPberNGhXJGSfMOSIV7zBwHIkbl3uNxJA6I
OVFhuIvwqGMHnXEMUKWXyRIgFzB7WMLAcPMs8iV8Jcdkc5MrnXH5bOmKYlQ02IZB6UB92dHtKzYa
30d3Wt7FzUTvmHQkyo+MLAO0xoO1a4/krcMPuGnb2h8LdpJDTtQDkNnmka1d6lMkrxsacozTEXyV
kLlFiwouMaJ/ZPLDQ2qJSOf7pxnp2qKnkOr7/yTOz4BPqirZratcWLG0cfyZTnTE4Usn3yL9sluR
kyupbdpziDZQyXpZ419uoAUkg+ZauaL/pvckUu9BRkR6e4sNxPmDMlr/Z1UtoTaVXC521aC+OqvR
Rh/wgwG+iLuaGU+OIiW6VxUZdjJMsla94sYzGqYxGOQnOv/AC1gp4J1kcoZbq6+4Q3hmykTXaoMW
WyOMqxi+OPTpt/BayRdvhAumQ8RJfiGN8phYQRdwZiCP4ihPD3C2dkbo/Re0wzfkonTYIB6HaKss
vCxmTaDN43ZiosyFlZ0Qn9JsUsbY7wXXqD9ULM1MbzBJAPbwQROq7bMpk2/sVbQr0r3ySUJow3Zx
xRUDkvP1fby361PEzfJtzK61rLI6g2LVKQkRxuBF0Sze5w7BcwdnWNp68g2Hj6AaRvn/2G1Lmoc+
mh6ycWUcPp4hyNU8hyvQosHOixUNgvNBMSKDSlM1pWK+EJ0ud3SiTCPIbnUsB4C5nUbVHwI/+1ke
iDDjiAwiOA/orI8zgm/DvCI47nRnRn0orY5zjeffmC1Bji1c3JW9tY7190u6zPLYWIdPGs5sXq56
ZFiWDzx3V3QyjTrE+5eIpTC2K2uWgBb/VEv0ksVwDAZBg7rawj7XNtwZjwiEvb6YV+lesev7Hfgp
3UFG8kS5OLKopNq4rMNO74bpT1TI4DpZLI8ec1I29ev9v9QEYUtQkIlu8OOv9+lxLq/0CUBy9LNr
j4JvcN1K68dAx4+svZ16sfJwn7Y07Z3oOSJQB8yYUSnJ0zsDaGH1L5yCQEYfVXH+p9uyvM/knbTJ
uZ4XE7ch9w+2zUNGPy24m++byI0Y2kznz1SFFJF48rEZ1q9eARynociSRh0AZ6aJBTwdJWjhqJDW
xo5t8qPH5hhuY7S6ayFc6q87nG5/xZTiFLHDZfbOpMPZb0xAyE/kVnQMnNXeTo2UiccQLx1lgyy8
8T9moUJ6XnBGUaLqCmakHhW/sz9AjQo4+cCmsKBtcmfICOLW6IiCxrfH74hZzA77tnP3PkOJcCu1
KbW38d31ZbNmPBEZ102aMrD14oBA2odTRf5+2TWKEEprHO58OmBa0cpFS8+C7pcKF219XU0biv6z
1rJxeLhjoRJYxrZnQRH0F0JG4XBFz/CjJxTTAUCSuWVwvR8f70mJgccYL7fi69pQ4qKnksM4170T
ogI5yvMbbY76KnUwxkaZXisvZN7QwXh9DY60/ZpoPwVb1wIFZ1qMQHjZOIg6WddJQaeEfVwOoWQl
u2z676W+CPcDteF/YsrfdT5vkN1IUAx6pjCFaWlZsMlKg9AqCDf571H1/GAWrf9WalKt2p5kf6KX
R4buA6OmIiZJj/Qlg8Q3lrImAyHr7ejMl3dZOZv1G9epHpwMlE5nErxcMkszNA21DTQMzqjDT7Ck
i7zREZ1MBMkCALLlUyw0L0A3cStd638jGnogz+oq/woy28a64G4o0sH+yNXO40LsfHovpi6lqzxG
X9ugoriYwOgeiRZ+Tnwn79TcKFIT3roIY4Ao2Yt5K74h8hjD5LaCEP7Oo3n+5M1JJHfWcTZlsET2
FrygdKKW+qqm93INNjbVn7V09Yb5erqMaK/P1qVOWf1c6UaiexTUe8KIQjwDa/aKz/7HJ1RaRXI5
Oj9DalJ9BAkIfMkQmn6HBypnbvMfOtnou5DlKdoNZTnBG8r6m5o/AIweKaErdou/QQgneg4LzSir
5aRespPn9xDRHL9Uc0xT+UEj0ZEdTtm74n9Q8je8z7//rMukEzIRjE0aEmocxB676CKDMh374sLa
vXCCS3kGJ4MzpUXt1fwMahm+2ghb+L5SJNHL0zYiaXnVlUWrfzq6Hvt159AbTAdwc143lpPD4TB2
PSPWa2wWwwcKh9rsU9RsiYwZ7nFU+uxoP2hgqYVN86egdQnUGAcjFUt+siLZmsMtGOgIID28qARV
TCK1hqKXpBTkIIRa5uvumI4PzqzEAQcE2Id7dF3oXf0hqR5U6gp/dEIqqZ8QggeWMEd/e0+AZmve
YGq8dfnwhEZ8xexKRJMVYT8XOvxx1F85zGBjo92zefER2tdfCZJvlLRlF9oh+EMBhtEASFugTeq7
sRxr6HK5dpbjC5CzyTeeXjftdYCufbQmKQX5zKmrpX7UaMssPlf2voygebOKE3uw/MMZe23iTvVK
75US5QJCebYqvEtn+JAmdhJEHSrCCnEVED/tzSuOwBtzP6L5AsU+7wQTdg5bshWecJVhW4HiGL4l
ttx6ZeJr7mE6SggkTpVaoyKA2BgzsQGYwxRclRxweBws7hlSxNi0ex3SsIlHdTBgSKt/01/hP+zw
Wg7ce4+oT66b/bLZMVM2LqqbiwLAm0Fl14DmZtYZ/YGjeQXZ28KILHTOv28kG7xyCMF5Um3ETOwe
ufWpXgkvOZ057Q/aIQme7d9HstsNVvx1ij/VIfStYNV+4wnAY2eTwKz0qx1sibeJCVVukF5xBdMc
8+XAtHO/SPA2FwVsSi9duJNF7bOwo4JHNS2XLzCsCmUcapaZ7RkN9CZideTHnkKeQy46DOhWwaM9
Wy3sBfF4k8oLxaIWVU3kyKoRlqGCSLvr5lNV8V4nAZruBtRMGuOb5OIB/248tfcA5FCNNkGAu8/s
qrH8p6jk5TkNeCBoGhH3T6EpoFIgOLti0KtYlPw7jPv9v/RqL2dzLEzVk+57k9+HugqbO2JTT4cM
rWGdwPQhR3Brv4hRCSSqH472aoGi/NCEqY0XovCa5pr0HC3CzKIlQy+M9MxDGIwYuSp0MJTMQHZN
6lbQXvzhsFz2eD7eeTZ4k8q5Gq1qTyt6N1W8XR6x5swWgBKZzsr82Z5xZFnnaRdA9x7edj0VYUYg
akHEaJgofyY7psVsG1j+rjmAmMmh/fwOyg2WRJznc+TWOZNJhHge5HMhdx0Lf9pxkft0yPfCLAul
CBaS/D+PN8low7aODaytj3ndS8hYmbfbmjc7SrIVXLLQcncc4u/lv4TjFSpEg2l/Fa8gT0z/Bh1G
0j4k7IojhGkGbJJJvWGlCVTZ50aW4Ahkq4bT4kA2j9UMkxXtnzb2PscdqabqVFjsu4AXsMRLSnUH
z42UuiRrjBSFlBRVCKjJomI4HRJ/RkvgIfSCqRGuX/t1RlPA2JpJRD4uR0M1HFGobCxmJ8CHnDvp
DA6+/LWroVbnFz158FRzqinGmgmJfp9ec7K9swanfc13Q2+aWFzWjD0UAuZXAlenju9dXk6T5C7A
OY3DESCA98ONpHhRSf9mHJ0r+Amrgg09wu/5LMC0ByTb6I9MFKDaEAyp3bWSl5XvkT5kWZdslyef
pfUdVvor09H6+bOl3HVTX5mEP5X+qWCihpMyxzEk1eClSPwji52OFzotfYKMPYXCmxte09dmvH1A
b9A6SBE0MCY6UlVqfU8oe//8SKA42cPE75iIUA1CHWTPBbYr5OfNnx3MOKWTwI0BeFHYNlH6DYVU
NwenWODumMHQlC3hcztjzekVmJbBVeqGzaFkTjDJtyYXC25YbteT1e+0kCMNikbQzMLNuLAVl2He
MvnajepMi0cu03lo6NdzhqFj95zlXsLt+wGk+YCUGcTa4i/GWgrTftIWloXH8lRo+A/5Mc2e3Vse
v4gswOOziTYs8yT4TKTaeYFWj5iR6ZEeUbHQ0aBXlP3n5tKga/Rny3ZEr91OxxNEjDAM+HUoFt2+
hOzKjAlcOqr1rwcNZhukK7QnTqoo8uPdizkUSmFEc8buBRl7/EEX7lTaAI5+CGj5TdfdGpzkaRxJ
B3RKNdr2BKiwoqKihgtbOxGNqSCtZsu61hwgWqCp/ap0nDLbxkHqqT55pYS1oBlmqdyBX5TBzKQV
e/v2vNOqkgtRKJ0pWHze/MHb+XTAnBCEH5dpGfoMC5y7mB8DPkN8BWAwmCKfOjswlLOIiFmfYZhu
MhQF7bTw+/WOstSDj1eKi+8KRWVifwSTFF8UqK6D4+nm+jB6PhynhgFrAOxbllwlz6aq1OUXzYi6
f9vKhuPA7ancpnPDCVKAOGnMbjmt1n6yrF8tZZ1+JVLgqFzYpw00KfWX1WhDyonTKRAD+BCGicxy
zSDFqdn543kFk7cvjaOAFApXxYh7bx8ErRoJyZGJ9BMYoWIp3airb9OA7E06bbbbniiViepwLbtI
08BavphboxfYYMvY2bsRfMaSRIP1gbSkMarssLphYRkqvIIzoKoQcyuLtJi8sBEfNhym9K9L/ppR
LkDanRZCpRdmra2Xg4KZfdPUowhDhBxZZ/0xpru8ICJFia2swAPBou3Oy6thWGh96OCt5WE6cb5P
MMsfBnD4fD6BXgZExTAeVUrktcHe5PyEcw6K4ZJYvk2sMtTA/AmBD+N9s54r5lGG4vUEk8XHqTXK
mfbkPd/TxDjWCz6iR2QiMi1WEumEXaQZ9Si02zLhc369eyGyCGX0CPgIifbquhWxXPhRR6ucW80R
vQPetRM4hAzEcGOBoXZPKI1csQUazpOj0VUfBxkWRdSh8Bka+eRL8YkcxZA5DyZau9IiM0G52Mv8
afOfu9TSKVc9/1F74z/bAmqGT2gy7/zj1r9++R0NsxwNxk57FhoxLFOItHmDxiMx0aafIVas7ZxV
ILxgF3m7uvuxlSBaDVEX77Zxz9FyS2nDYoMJ/WuRp3nVm2ipuvGy/gweZZxTwYCw6nAmHqKVJKY1
n+QDhEApYIey5ho3Ub1ftd6BIVMlmsNUGW7P/jcB+d45U6lb22eTf7qJnmGq0Kk9DT87DAWd5fe0
RUPlx+XFQpnGSRnkRlaZZA+k8m5pyxk2zqaCAM02IV9ssdsNtyFb2CjftpYW9FFo2Ub48jkvT/T9
gGz+VVEybciFNvmr71kNHSC0JZFZlmJ6uUgp44fKJ/RsqMpmIjVAU4an8HYHHskrtwFPpvwKjO/h
CViyDz17V+P0EKrbv658veImltsTB4aJUF5Epe9i+O2IQiJcd6npqjqh2eiQBi+YfmMHBGtzn0u2
MNN67Pkk1khKhikdGHz1EPXjopJBWrG9TKWhtBb03snVzjcKPeMcVG0vR7WoE5DY/SqF2eFgTkvz
yyUY48Ae+5I8m4t52+IYVruKuI2a3bCUW4dLYLJoGLL8+ZwP+dF3HHJ0ZbSwIXOrzjnziZkTYmTd
Qil2PYvaC7nhtb8HFz4v7hZnfwrSqQVlzUSxjjRDtdp1S+Q6THEzZptTZN6uqsrLyZKUi9idH8fo
PjoVSYtSkxFAtLS3IDhk6sJZ6DBKdDu4rtW7qu5JN5FIV18Eqv03qb3+nbOxt4Ae6sU+m6kRIvxJ
B8JO2OzEQxDrOSMKioUnDb7xrIjAPTF/UBs+lyiAjszs3fijeSa3T5jJuzuHDaOJlK3CPke8z0zP
tSQ+ZpFq0PtboyJ1YUfOu6P+fqwVXxHFJ9W+fGkDDY+mn401n+zWfzmN+MrdDIpD0ikR06u6nS80
hKnVMRxRE8C0+ODkjeFTzPtQrs5uu6RIS6VbUkqIfzJFg/8kBHsmnBfy5vZia3k6WjkksFB3+9sI
zAwuttY/3qFZ01QII91VaTvvk6KbfHP9Otp9nxuCmoQ1S/GGEgZSFeChH/fSuTfPZxJv6o1jy4xC
PRND/D2lqL8+WUTBLA+lDDTYAMCU/c/dd2MJ9SnVCGzpXs1f3B+J/KQ99joxopKwphIY/KV2FDCA
Ch8/dUgzcNuuzWnVhu5dyMSf5iuAdTvQiZJIq+cPPzZcspp/OBS5dTYS7vsM2iSXGzg7U1qCnhhz
UWEe9kuicOSjqHGVKV6ceGU1uM/i3XY0KxnTczdhsPR/V9NWnOVEhVbuWiROUiKOaG0b4PgHmlNh
9iLZngm5h417VRta/cpmjeWQvt5/zIJd3Y7f/wPllRXHA6fBhDEjdA3m0Lrmhzpoz9DQpIBs76Za
X+k+UtudMsKLcELnw2Trgd+E86dHW9AVtPcbJ26SuNcbG0/757LbA9JGaYaBYkS7zzRaGP3xQQ//
bR7b6im1kgt64JFfDhS+EsR50EgHvHizvPRPGD008ib3UVitlyGZyam2oRP1BQeO3Yw2KrM1flXd
eWzGiLMHBrzKd064tWkgVJCiQ+9NuoDS8LuEGk6N2BFP+T7BF/Bc9oLOroHk10PiOjg1w2H94roA
m1oJYHRvjyK8ES3KO7ylDJm5MHheqOr8v9rymI3zgz0OdpoWSSkgrQ3gs/NorY+V8Vitz57OCjUj
yRND2bKeF/skfsqR7uTzw4C231KsrPHCoEtHhCcv8C9fMQwbdy3IyFRknvkagsKknEvJ9a+vRZiR
q9cohVEffeHDK6kih2O4dJPyne1KZYtxjlqaTI5gbsj6HRvzDilBg6DlpGqXlhShK6InRJT2fSgD
FOqUl4D1F6QS0KzMOkwIyMd98UMpVNyVzynp5QAPsD1qiMR6C4ZZZhZHz+YndGVTUTR48TyFvEJa
/Rx+Z8np7tYV2jioJkL4IWvcnMXlXdV05VZNve8YPjsds3Uhzh0ThKTBZ2VDu32eLUhrs7lFgfJj
zFBBo/Gl32oPwHqvcMojAYmOvft/a+kNqRn4dnW012EO0ftRB58BkYlm+ZRk4X209PzPzKiDtJgB
6tOHyTcLWu4U0nXFuQtp9vzj2nkrVG+lmhGKJqVSdcmBbLMjvPmc+U3BsT45V9HYYkSAsO9AEiY0
yk1oh071iXgVb+kgwUInPRf5OSbptyxJ37F+S+Xidy7/xJzShuau9M2yZeMup4BMXLgjaz9K6aI0
9mYHj1CwqRzCXGjmc8B7jMH4HRSNZzFDTS5qH1AO+Ni2Vh1g8WFKJpIDRF4BqheNq5X7JddcmUZL
pZmJpXzCYJfrNQIuHHXLOMF+7Lzcq82kXf1twvj+ya6VBry+8YX3wA4tDye39E3t3usm834DCiiU
r5oeB4Lk3ctBvpCOtsfT/5Je7HeP6yTDrWUr0YKeRIEe34VUWs9a1jUIalzpn5Ft9l0TRXIw68f5
0wxOnLyI/i1QWahx13joG7DLDUdki9VSLRmC4XwO9vkEWPo0ME+HrXJlyyZxp4Mfr8X9/B75tOxy
4gRuRHHa8Zc6ijNcIe5QoI/JFEq2YsU949si0O0WN7vcyXbYujp4kzejLfh8gXiiWpkBoYYdNXdX
N51ReYNoJSL5aiRZnLcK+YOjhbP4b1N9aMNRfBrz1C9XF2LG5sUxyAz4XJ13v4l30KvNXfAjZ1gz
lij5RJ7DttEDcWK6xTbyXR0qxgmpSwyDO4yZtg/AwXdZteazI+cQXNEKwipKg1itPGT2Nbyku1fB
2IJqkymjccTQbEH7LnI2DQgKcE/gvTaykuvDNNIublV5eXRhXzhVhBMtdqn3qOjHTNKE883l8shm
y+oP6+3jUDCF8n2ZkvG7wMt5twOuPUB2G1vZDZnni40uYSKE4A5H2MOgGdA3JxVCr8Os0P31RLbd
lIc45Zs7aCnEnMhQsyGra9ByjwO1dz5efoeigpFAyJ474sBFPXSsX9hn85hxepSu6aOhULGCG4Ld
8CkzDAMZvLHEQWpQ3EDWd6aSFSjb9p+1XV0YUHVftYej1Gyhz1zrmEFcCgqeFWOFxaCTsnyNh+fP
b0L8fB4X+k87ltViX/f/JI5HZ3LQU79o99npN0wAw4QhmQmVaLInWYyuIpKg/2+wxqwLZrP1C0Mb
H9I9UlLni0F746KGCZvsot/2x9uQoYJKtRyxObK7RDEvThX7oOdcz3cYfg1bwQanjUhvBPl9oN3G
KHjCO+PJmqfYsmpWxB7wmzXK8TUwW9DdZ3RVpf8cS877Z45y56KaRLif/cg9SlNvr6oYvlaKzcwY
CCifunVSIIw39ubcSuVpDyj1iAD1vYAYM/E6rKJXRXf3SzleSSVEZwty4OcusSDM740K13ZpKOyR
RmGSW1yWAsWggyAw//9/bSJ87la+fdaqFjH0NDpH9CNInrqna1ugzQHt2O+/unU4+XazDOagJuvR
efTmXbHI/C+ERoCfhztohSz1K2hTQ/o2S+1QvuLYLxQJl+jTevi+T2UEnAtlIPLCKudSfVSlIirb
kk58W20A81NVXK26IMvzGI2hypzIbySoXFyF8kXeCAvfDWtoz7JjVaWC3CMXDra0iErmTmzAl7e5
QkVPX9PaXgEmzXcb49Sau3EmUE6jMGB2dqWg9Z4R5AyYxU4YmZajw1GIIun4D93EJ6wnMUyAdQyB
IlrKDL5ldabWlqDW5S/YaJqdwbtGgX48c5JfAg3BeL6x3/dFQ713nGEPAT6ty9co6qMOCVyTsnw0
RZlaB4g8vypIcsEncvdS9wgEftOxUf5Nsji+fultTCJNBZqL//dmbfqEdGfTAOZ1yEksaaQCnO+D
R9vxygzS1HdVcYc3UnqKatgoJWcqLGeDleZXo0bLtDJOvTv6dVKz8aeQL9JoYCzxlcuRHmWBp6HU
uAjQplnlzXF5sBcKlclzxu6gZShmUfolSDJdFJ9zq2N6yuD5vUHKR3vPnVED5wCcZG3XyWMA4MPH
LxR+cEbt7VwSmhUllGAxSnbuPfHluMvccIaWVDHUT3ZyScCQ+QmZxTZtPF+0nfc7w6X0z/zTIMPD
VhrdNoylAEoqHtkq0rKKZAZ8HytJMsAvgBIrFLHGp+GzcbVPeQBMqBdrlTUb49/O3YCdN1x4qCU4
Gh40lbW9ek0e04uB1jIgwHCrBFn/krsX6x79mrxS0gnRRBAX/tz9YSUooCQQNA3Y03mamrGendv8
A5NVztAK2YGV5kZhb+p21RONTbiDBDE1p5klkgbgY/RDH1yPFKrQIU9crjMMxZcvlcmAMyC0Lcli
+y47c9t008/0pIwDUXXLyd+/TXw9iHx4LyYkUk6IOxUnjD/GoVD4ubXwh17o1SxSdIRZW946gYqp
cyEQBzRiU2O3+4U7+YCEXKt0eVGF8q3ZW9sAb+qGLwpizguzU3z4iFXQ6gpgPx5kLYryUCN/9d/E
AgrCufFAolVnAUAqOERS2BTAYJi+g3GtFq2CXKGMwYGJaxmW0s44pzYu8Eff7DUE3Bnst5u+mxSP
435C7clO7sYwtA3hGxq+jufmg313Soj0m1TVIcBiIga/rZ/i3w6bw4KOjmd1zP8435UehnIPf+XK
Ob+Xc3GMc2U9OUX3o6OOH10f4kHXY69Jmok9MDmkhj67cFxNDkjuY9dHfc5ghodwtqDTKXKT7ni+
1zCOvNFeIjeDoOZg1KTBwfZ9587WB1L1yRtKQHRlP5nzLU9+rERJUzOn8YMEbQDBzpkctcCKEd4E
xhpFmmbfqukezeehlGjM4PEPWstxb9KFixbWGQbx5lU6KUPfonL3FTxVsQ0q8V6vRsQD9zaYlLyJ
aXpap0DLNSGW+IsjeRehb2XA3zRFQ5bUPKb/ywKi5VMhHXRej6Aem9OjrgQG41vlRY6pio2CZ2VX
qThsPJy/0CEwxdjn2qj9chnjIlq+QgYXLKLj5F5H8ic7a6hKfmt50Dss5xZjadE2SuUmD6jtzozN
2OS2TG5/gPsx5KWzdvVbAV/a/H+3ISr5JB/1mJKfYBmlV28Ka3ptl8HSw08HJ5byVw+i0/wZOeKD
mClRTWP/h6vE1YB9cShTq+MOa2AM1bNRSx08MmMyLynp4cB6Q91vZSxCRCGHop8faNaqUbZ3BDMg
vcRShgpmIZ0nSdRLMwA5gewTNERKZL2TMA7QPkyTTovGvjFf9aQSDMHxhjaPXMSxdk7w275+ZouL
c8jQB6x8WXZmsgEd49PY92qT6kHGcMUc2j928iSzWcB4aD2Tx2xICvebY3jXYt334ClsBXXgGhFr
mIMTn4X2w/tdNdqedDpg5HFjYo9jMFN7QPCox65PjsBDZNh2Up0enyBe1J2WWJLspGXHAgMDszmy
/Yx9XNjm2NQQB7qGW+aSvxG15xIw7UNTP0QbhCzNdUmbm+CzkMxHgybJHB5bySYiZvhfm9NTaHE4
OHPA+dh3PQyynIXEwEJTwIiAjienKOieeeUa9LvZRuFO7itZAYeNvSRmZcrrRIp3ZBz8bTb61KJB
iECmccjd2lwCbvesAl7liPLBC2r6eqqd4bOhD2ALXCyE6OuZQQ4pbeRI8CyP8CAz6wPtJ+A9MO0W
y8dq6gYUMLNkYxJ9xsnBr1HXrluQ3665rWOEXVc4lofA+yqnyuMICwWfYeFofC2ijA5Q1Otr63RD
lpsIDYidc4frVmnECAsW7Z8yhxNgk3fn6WNHkcAdcoMJh2FNf5Wqfb6ppJhCbH4PNLOQEW3G4lyA
IU0V7/H28jp+vsn4G55HL+SxQCKuhf2mwzL7wCvwgxek7Mv0a4+0MCgUJ1mSFWCxKPqpzfVw3cji
+hf1+1xTDZXKFAuy4QZSdDKwIhOw1A6dVgYZVkoT4bvOD927z+NPlEDaoxP3GVVVskNkSRaxpQV+
1VAXAI0ObYTUI/W31pLqnvjWbeAP9RjB7PwvwDR9GCiR1mjH3Ev+n9LGWCCn9gho3YdXMuYrQXvg
erZqxd5QArlwfd7Koll6XQ84gwLWUsksa1N40eBOufiE2Ts31aX0DfK453zautaPn61TRfrPjtyI
xarQFlulr82MnQWi9rcrk5qch6ZasIXes6ys8Uh5he6pglIHgczN37icN6XyGeSXYx4s9a5adteW
76f0akBn8UvTQjKjQqQgkJlHXiMIElSTgARVdvXbKWC8Fr7+uxif0apMgChABxroVCPw6uTACrJH
rhW5NYHQoXE0Pd7Dhl58uax3zqM5I8CYPguuEHJZV8t5fjuk62JVihl9gG3fwHPu3Hgcqd3+BtBL
Xp/vI97UJErpjrxl+tQsmtRq6otTwwlak6XIs2FLW6GihkBQbtISwDwAZ8cRQY80hZZ9+R0FRZBm
NDnz7r8kGbQVP7QvyWjZk+eGH3Hrmz7d2UXFPaFkRfHUlOkQ3S9N/fn3yf2N8CkScnzfYRscWLRN
0N3ZJBeP+wpeOrrPEGf/oAicf9Wq9ZjMhlahafM5vVP7TLIMdvmbNclgiFGzbEFDNiO2z9/qb4xY
mRLrn5IYFp84oIfdypzjhup/cFHKR0nhG8rP6iPG0ChaPu10Wg17KfiLoLECKeOAObWXlh5gSoNK
yJCamHYS/JN+EUWY0v/RNIAfQuSjfbknxP+YyXpl6ijT3LOnKFFtQ1zOdZk1KVk7ZKn/fkI1nQP8
ApFo7T7C7CCiseKqKJ103IMsFaeFa8/NVC6+b+8/ldmzFc11wf9HZ21b5AJn+8RiKn0ve4vWP8oM
fAnvvtlIKU6inqD0zgxYHygU2AV8a35rrGPoqvqJaxWVUt9zbrW4bbjp8t9IhuR1YwpbNRxsm55m
d+zG9jvKSLYK9yjVziweSvOmrmlLRme20jE0gOD44iIvQ2ut/t8FWm4LODaAaDeb0egUwDN/3CHh
1b7fu2bPNN6zdHtjQhmYK/kI2Blw0pMvKATVjIGKc5nft0PJQ++Y71ej74fgMn0r8CFq0kTYB4gZ
D+siWUMaWgKVcdaTmUTxd+ZLIJKGtmb4sRlg5z/8MdYMlC76+b67Yc+lCDskvJy8Z5Ru4141KT9v
MxahYd+PD3iwdDW7LgNB1kUmPyDOvD+n/RudFmpryFRDW109ku055ux7u8vHWZLjIodt5w3u0U2u
dRp9B2wMX74ePD3k498L6ahyAAY2t44xWFbQG50jBWE11PpHWH53i1+HlLGWWEbErx0xcJOFJT7F
VVGea9v2UwheMaZ5MGLPiqVSYTH9VdPuSugOm0iaFFmlBsuKKNTu1iVkwovehEjZBxS3pRfPoKxP
sOVU+bcA8qgisKW2v1OxGsBKQJ8Kymvyv0UWYZZ4fqfvzIZI31Rnbz+8abk7OIyCDc9le4pnASxP
0DmiF4I8q2Tu5AjDRwuDRoCmKtWdprl2zaQMTpfomsPRQL2G6VQJHbputIaDhhW+yHEHrnWO6zj5
XsVKCKF4xTx7RAR9HUylPGAoGjuIcSjofwHybmoBPNYxjwlqIrkzRyZV8hfto2kdo31G7gklJawl
Tnk4rTugUvhuYRPCumTH37pCLmDCaJxlOnEXwQKmJbJjuF51xGmnZfTyKOMHHGebp/qbH+me+WTM
MyjRDrM+8Ep0//nbnQ0u4hlOVNi/riSBwo3VA5E3YXjcl/tT6SBtyTSM9YzlFaIHM1zvsKrkQOQy
GEri6qSLgvYmMYZSXgswRgVaJ5uqNquOR4x8h91pfN1sMHcYEPQPXq9nFqWUgtEnxn3kZORUQVds
Grvtcn8ixQNwJBneq2ZepIfKfWY2ZAw7UtPLdLH8q5zvTfaQBFTNu6eAmkqY38gxYHyu8cSpGwOj
uydkUwBzo0njOrbkhvvAsJ7js7GTsVxNUT3TDXG5ElFBuFWxFImw2LTqfRVJ0a05pHL0ygFvAEJy
AHRctofFkUxcwBb/yHCw5g/bQBpp1935mLZfcbFmJf1I+4D7md58OHRcUc2rar16/tqwCFHjN5ww
Hem6CxRn4C8IuQztQblesUpRjM2QEtgKwtI0ZTyhCn1DYPUiKBFk0dcLJ7hXglwvVq/n+isJwl/w
rBURgm0s1zsEFAUpwrKzWP1UEpLCV7lnF7pRDyH5xk4sqG14G81Z2WatfNor0wCXQ+9PakgRzIb9
ZHkUVutTe90OzIyAW6njvz5fTn3+slqaRcNn4DWzbU/zItCEdqpZd1VKpWV4fdIqiSztby3u7JRV
Te17AiH5XcmiUZ5QZqfOxIgdzOwm8Xki1UrYwI/O7QSRCmTGLmsEtVhqeU3Jx+HXEWUTS6y32Ziw
AoB3xdgd5lP8UBAkrMn8S7qB80MJS+DlH/msyxRJVSJkRSpsTreB2qxsGygkZW9rc0lS1Rm4aE60
Y+sN3ERTRwpzMRHk8A/YAYQMKaljVq7qPNnusq08kUye8UVNZ2uPURn5pZoc8ub8f2BYdP6DaF0Z
XX2dOmesxgPG42AeKEzL4DtuYLwlQ/FgUsqPtN+3Ex8LTqbnpdoQFnU+wWik1pOtNsZ/4DEnYSJA
Wr7tJNESUDiZbfkgGmxbSr+PkakItKDoX+PLDnP0vPP3F8NUtD+V+pe9odanlJM7Gr5zue9K3md1
Ez//taChN3Jjv0lGAG/eSuDM28sESvtN9ncjQkTOvSl/FQ/4p0MWIIu//OeW3c9lgNS2EnuJzreg
eJcr1IKSwessEuk9WZm5iKcQgPQFXJutQkcMlulhpyBLb7O2X+lp/qEqnwTTR29cQFd7fv+ekzQ1
QpzVBgaBy4wa86csf0RaOr2SqsMEkKMVrIxGK4PIhJ7T7tK3680uHMGNaZOMGYF3/BcODcAZUZRo
gC6xuMNsVHkLz3hA+2cif9qsGAwSdETXfwZtRhwenKNGkWv2Um0iKJbMq9J7xHdpwWLeEvcvApHF
saF4ooJEzmO/dmzs/K6XK2tia/Ja+SoVExzPHCG9Myan1EDTu1T4wR1ppBut0LrMC3EWIW+fshdd
FzJRenL2/M+wvlS2LyoVgEw5AElm/Py4dctNDP2GZzLlVspSOv2lvuG1q2MLhEgJ5jQ4+4cBXr4a
bWSMdcE+dFcjuaRnJP/sFedr8Xdg5kqVl+QrW0JMSX7pVDcOIwA2lGmobTd8f4F4Mky+SGOVQjsI
YmH1iADegtzR3GDpP3Y9TGYiGkfBCds8i918kBUUog5XWqnpyfnpvU0qLU/oYsNocukI62Dl2uRU
9qtVQINri8aTZuRSJvGz+d5RU4FFEAAylTrr6XYKhdgf84xYWr4+nM/8aVJQZNQendTaHIUQN8D2
fjamGfR/vEzHBTZwTpVVNwZdoKNkJVA2xEKjsQCZbbmJF79wlUy4YwMCg3wD8NxnBtrM2sids9dY
Wdtbe+n9qdaxsO0YzYKEkRdyWIIr9omQykvj7e9B+/yiOdEv5zy2nY5WBnBlg24F2UV2pS0RFIVN
XrhBXEzKSDGuwM/yLXuXTbFjaEnRoMniq0Plfjssx6VIt64SgjjeWPuMLT1VeZoF1vcClIWtn3fI
vNo999y9XCfCIdAqaCF39KOWsDsRqCPzcFgoZi1TpgFbjfo6O6agTNbHBZTYdx5liDH5tZsGQs7w
RKAvQkM8alsBvzXPeJ4D5SNcYVTUPmpMicxqiljKWggCXAbIyx5NvL2C/jO9pOhkX6ZY34R3SiSM
w/L9L7upFjIDM5AKMlpKMyUD3lCWbEQDUD5J49pMEnH64I3+9LbUMTdtIyEjxYbnBSMIJ2qI2Vdy
wV9St1uc1eF2nptjJ1guatT4w7JGQVupyIs8JRMZ4tgLysx9r48PlGj3u5fizwHBVg6qCK0Y7W5n
FYb3SktOJyXfaTfkL+WllKS/rMGTPKQ14XqSDBSzfSr3qvRSnli0oOI+YU6YGiOBH1WvJezR81Sd
eOuh27XGSANSKqBM+nNNxn0sVIB2o1l0/9FL1Hvqj6yVv7fIkgmWv6gAU3S3x+ACFx1VD5+Y9qjy
a0vlMIKtuyFPYJDMcTK7DfEqd8ui+nJWTNzzTIpLdSgQkRqjojLGt2m15/kSI/mR5b6T4/sz8nZL
T7/xTfETMB+SPhZFjOdEDBpjsrqe+2tlfvJLozUtSwK9GzmaltnDwNzcUE9hifgxk1H83AR+g60m
33ZaJxosb2jms2ynJRJdV5f9/b2sUaqeYOjUueCBxZ0v1QtXe8pxio1rE73G9VAP7spAOoRA91kq
TbflSmaQuXlHP82NFTEPc7hNYdRzWaIX01tLhYTa/U2uCm4S2lhtLWT8YKMNMq5sPqjR6IfATvut
grOT2X8UfRQrJPOMxg6gsENX/xkNqukvQNB1JU0OIDtwPv6kc+nJoI2mcB92fjlTuVPXwSzK9eEz
i72OAe0x+Dy/PxLDpfnCJYMHwDzJegtypD495dng96LOJiO0Mnx9kgLY9o76WY6B969CIWw485JA
nwIjmF0nYdMJxIdW4Z5Vs9jLzTdYUUwZu172Amek11fXxdmQDb6mNZea86iKsON3YEruv1P1Vgj8
JPYSJ2JmYUvXkpJ/tbvquV6I/EJcLiOJI9PdvYBRq/eXrwjujS65cWUg7zMWi+qZXNFM7EfBjJBJ
9+K0S5mnQwdSUPU/Pg1smHrgM+nggpoUf2S5KSV+xhPyLTaxAfm4sknnls37pl7kw6iyGTRdvBTT
XMSzlktBkMfKghGXmuONd116SoINnMUYt/pWA0kWkq8t8VW2yazbI8SgaapT9avEUFmx3b7Vu046
I9AsDhHnCLiNN4NQ0tP4zzLyJJcP1wI3YipgFfSfN/fpwgaHm6TNBLjRCeFyBH4/02hkZ8MAfOp1
Cb3MI9/iHZ5+HdnFk40XHU8ARzcSpf5n7SgS5TA8o0DuJOuCEN0HDggHXyRV/ATVQPMMV1eKeXxR
GTW9Oxb9VFEacY7O5Bz7sYGPe/JB0O+lq17xD+dc+i5npfsRgV8q33+OjB9xqc/vslSTZRDPqQ9v
o6g5MMsvtE63hxbrPK1FG/u1WvtBuSDJA8cWxGFfrTO6IbLwo+hcG9gMwUDWfzmE9zyRVZi6Qutn
Zoyf7QamJf4QioiPhH60znpkpr2QuOkTTmoo1qa0YxBApQ5G3IwbKmAsxBKD8utk10maqw/KXOM5
1d98JKhUyIEoEYe93cLaLlkhvp9hqQpuwrBxHchykW+t1K20bR2/peO3BzLuNQmWa7xq0cuomgVB
p7XhQVoaGfq+bVvY3HFfHVsNy6bR1wfMYvpqvo2YzEe0djeo0CforQKhpVRHi4Q+bjxy7SNO+FNX
BfNu93AVh/3ryfYzqLbIkU/cfRcu7uajHEQZrrphcr8vV81ZBZEb/uyELDCsjO+2wKQPx83gOAFn
dC6Oww/q/vNlVOFLp8TUkQjrH4kxdJqeFyuf6MggublZ0SFShp7qI3VEcuVkikUnWts86ciFFUYq
8d3pSiBvFrRSGmB92bpXzrjay6J6bcvrHCp7BDymzmCkJfDsWSff4G1m6w/ceeBRgOVU6fkLvhPw
qqGm7o9Nv4cXVjPMawcDZJvU/oo5mIhSeOVWNQIFDTwk/W+LgP7aR83UkBPKrihqip19eAJlh4DI
Ug2EltqDOwfIimmqqh0h6ySkFDk8otHEX/Zs+TCHivHdUXQPdYlpL+3duPu/TSA4qVbq6wW+f7sJ
uypCZPUWxeqD95+EA0vuFQQgCw1hhQSJggWy2J7fCnI2UuJ75srGXVNVJCf7zSJNLC2epDPLndph
bicwzWiuhjntJSyECVESriV9LQaVwVBDS4yCGEMaX9blru59UKIypT4Tsfhl5LOdaldoZHZZ1Umh
IZcy0Vv0uXYFL6nkgwn0i1exQ8JiYAUN9phMOx8b5tY0K6NlSGP2Uv2m+p3c9A4wy3dt3TK+5iYQ
ZQ5DC8gX2KrJ+U3QQ23Qp1VYHb6vbLSTfoUrYXW+TKVNnKAdDWEzNfHBY/sBRpy+swJq2SzK5zXD
+paIc35LFnUBvKMu31ReLWvAs1bJ7ZjJlvfwtHvLpED6H9vK3AsMIsLlJITfzpBwKxSD6feaNNNw
FmWVqRamx3Q1ATu101MlaPDCN7+1NUtqh/zmDD4V3RxmuzwJfHx/2SjUb1gX0st0JzUjqxwO2Mfy
EcuEvhx8zXZiNBSBY0K4hT2SFvvJ5LYIvBcd6gH9akSCpIsNBeAZt+8uNZ/ffgCVdzuxmOHr8lmt
PzShJFCoRvhV3CNLTVeW53Q8DCH9eOCMUHGU3Zhv5XVLVRtrL0bCffQSYVmbVV0rRdynC9pG3lYh
RKSLoq9E/sYK4O9ApyTqbYBKTMjGvV77Y8uycM/U5UP1qK+bLJdBzIzIR1mnjcgBFWJCcFiLMa8P
2+PZdBnjiH8lZX+wezXSBjUpya7qwzc94ZucHPD3pua1M3tlN7JkV+7eNDCXuvtRRCGHab98VYqq
T4HR2YG3+jyIv5LNyPHKNG8LNWbcgsLDqBs8XrOWDpxLouNEYDfHrTHHL5HTT06fqcOYqc26yvsl
Ap5XVFd0zs7qo81fNAge7rYiGhUCQpS0VsjgMnkmWfFXssdCXmhV7G+M+b56H5vw17jweBsRfwyc
gWbwtI7SYERFULvvYiM5znuPe+iog9zwh6shJOLNC3Ln0DIk1ClbuZzHnRAIBU3ixJlyNsA6v0qc
g6w4zVn0g3j0yPZfz5v9M9f/89H2uTdFkQm2kinJyRY+q7KSICYHV3P6DS6xJLWaT3eU2g+A8dNE
gIcKTWy5qAwgV5KduD+l6IjiBdr5IARlSZK/BZhnPxr81EOY8N7+4W8jW2nHUaOsWex0SbOGwjk6
eYKBrPIaTO4JRNSqAYmpKyT+1oFPJLqjPMd1nX5uXazPVMLiJAvqjHKxfVS16DVRecaWmQ+iD+E3
oAxI/438hEGfDUXPQc0lp/lSdgbFIxkQAUAptAI0n33KZ8Hxu3wRA/ppPHlRd3k200AQ5BVY9syV
aH2gXw35EBkDqwXmLKXka7blPpFo4erMzhevmNc3CNKg+w68cH4gByXCvqy2TXdg1hXncGyHaHxa
q94kLKWFa5ei6XlEvSO50Qw/aX6zrHIs1NgL1CZWKnE75FqIlK2cb0zaSM29zZZH9LOAn0YpzJFz
tbXuZ1w81qFMFiwO5QMKQo8X5mMRjImg0jUx9l5n4Oc53q549Xp50e2ttAvuK5IV1iFuZ28fQJ30
PEdaXyNmYPneWnpuRFEzn0ybFIg8MbADwOZLLcHyPeumL0WbC42PS2ApS2+7oFwR4gz9kEgie5n9
m0jHIi7Eypk3xBoJE8Vqbd7Eo76Kti2+uT+t4qf+2T5rFmqOnGPGJj2hcf2txR9bL5q8VFYIergD
1kRqhY7tJ30vk/vYkza1qyZZnLuBffU4VmrZ29r7QwXbC6DMxajv7s+ROxnJrm8lStqTeNHTeI0r
N7mA/WwMRNJDERTUsL8kbTiDByy2Vu1H+Ef40q7xovbM9cgr2/HtnHEh9+CH3DSqp+fLz7rt0zAP
CifzwOj58G5ymZfeewgWPMzfuNsqAlPg/FqzPNGvcehNE84SvxQtM9HwB+LGOWXeaIPW7hX0oEm1
v5ieIxnKruFRHpfNg9He7iWqEQjt/MfzTc1ghoGluPeap9aq/FfuG/zRXmERRuIKkPfB32RaC+Vi
ViO4WtFS9vzcj8yocVx9vszp7myEHrsKedJ9u2+2Vg2twUX6Yh5yXVl0nWTu35/nGkiW/JbrDqp6
TaDpSB1qx211iDW124pjuNOoeaQy67+KP648cwYRePrZBYnpdot3lX3/n22TwVSROx33V5vB55JW
YS5urX5+JUBxOxuULsSFC99Bd+BNdeemzuxff8wt0rSqQxpmKxKXGd57ba7docqjixh4u/LukXc/
aTGIpmWqzpceq9iN8pbcu875ONwQ51Vi9t1BzYAgjwBh7rSj4SC8cX8OTwDB3OYMM1/3rDYgz29C
rDj++WhyjEETH92sHx4eEsgIeS0WVpcr/QHwYI22NclfPOG83lhoJW7Y+dwSf205Sqys5ePmnuHi
uT5lR2vqOqxIt5TxQLPkG+ykncwRBn8IHP/MbECvpKqSFOg7LK1Wg45bwSepHZaDZSvcM+QgPv8e
TTssXkCWeCSn4xnJ1tvRyWkOdqYvm9jHL3p7v2h+omnbBlZhXgENb3YAFzdoEShUVbj3uOdcskkd
q9L1H0lRLt8yUjGfF9vP1rhtUB0NQ6FEmEMlXpu33UxWty2/y0ZZ2PffCDnnMY4jCjJC0VJQ0Jyn
qME6YPlpm1mlZ8oxKNvdIAcCoJKdcbjPOtT/jsnxy2S8nmEAdeIX3rVjcd1cCGGSXZRvX/miGNRT
S8k+t3zAf+ZmAhHPMkIFLSUSs3/LYtYvxJI6RGZbLStKj88laADvydtWG0ufPY2dyYEU92aaXLgK
uyT6sqTKEukpH/ECD0b5KcQg6dFdxvHg+hRwA5h5hPN70BAW0q3CIka0TgsTjfODIu5honuzeQ4+
w246rtR5RTAlaPJe4KBqYSqNPkUSVa1GtQFOCgdsQJozzCDcMSMB2G2LIKICcVIwyqB1x0Fs9wkP
XfLa/L/38Dh5ehuabvGtUdvjqPDu4R7iigqrPVtrnNAdr1LIbiglTnWoUIjIV4dQo96Woh9aExVi
yRnFTMZ6CurMgNiWLI4OxphQbFKNM0yJ3fsq+sfjy8FgK5gV0hEhyuMUjovwTZXTCKZCHu8F8g9c
3Mxjg+2Lzg8z6/Ub9euJ8YiOSFi8uMrZdx8lCDRJpRz0P7pfP9werXL4YsyKMf95+IiTJHOVdiYL
pbW2TXJFyv+L/fBb9MJ8elEsDMmKhgDvuaBK+uxuGsPKxFV5NuudrOvH3qfJu6HIh1bFltY7OOsD
EHRA5+jKp5GJ6Tmi2LGtGRE6zJrv6VAvphiocNd4wh3Ph6y9utlKX0K8IQpuZfDV+iwKnOMvVSLd
c6hXPuBuZs3yfpgfBHszP7QmuS8h3hfbHxTZxS2+NNeOBam8VzjvYCfAbYKNaYcNb2qfbAwEe0RM
XmXUtIkURgla3jEpLE1fsNl+RQbJ3sJeAu1ARsPPR3fIhki6S4cLi3h/z60W4Bo1GDQLeRMnZtU9
hDJqJECdKuGVXG7VX5sdp5/gFp1BLff/y4J3Vbc28zj9/lrr2EqjQeTI6kUFQPerbdxr+1fxyll+
n79Q27sZnIVwiA8K+MksKZ8FnEzDyS7cs92tEMIUlLnRwE6vXPlc+scJSOS35cyrPntsMHEeiS9M
3HnTd972khh7AfjToHNCyKttSVKAUo8mYLJ3CTmtkEgamaMt+gF74GuKWhzSMh7h0WfA+MrQaKd6
V9v7zgLHJVLqPZgskbHQnh4YLsYxuCuQU+56Gwtatm+8d+QhvlWAPOK+hUPoxKY7qxaQZ417Gt76
Wr19fW0K3JPtvTfd5jVEv1RGjo+iyqmCgrjqeBuilil8c/cMhCWq+w59Fa6jV06zwNrqQ6AbMn7G
G4q/PiguvPcMxrlAhpT0M4vJJen3NTLXcheNTauan+dlFlpIuhD9T9Rnq4EfpfNpB0qELhuzSRUF
/FYH47x2YpN0PyOaiZvN80JG7zEevx12UYwvvS4M6C3f5iCBjh29ml4ZuuBnfmjlnx9d3Lw8/rsj
6h/aH8KD6QkOJOOfV4E25ecX3LKTeknMDaFl2mkV0sixtUQ6jkDQhBclByK5WGvOjkIrM0aSoDzx
c0vvfOuDN2njBJQyJOv2uVhgh2A2jSUEb/hdu4FZUNXpUt5A957s1HD200y0hbghkvw/xmL/qOSX
rBCSwrJb6ZHUnedBPl/6i8ZTETOfo+wG/T34JlrRK8cbwVItWEpcgKVldH6Lkb6HNvCEmnfUtOxq
bB6v4uFOWZ4llQutvqtonapLsS2FgZs4jDR2DhX8ZnbbM7rZtOOEHNIMef302LRGX4fcfZAdXx+a
utBLnpA9J6OLMVpowusmw3g9zxS3jpS3d396KYXgSnZGI9ctXtjS1AURTk0SRfY8JuqRO8LPm5eQ
/2CUnKmynzE6Y8dKzqr7+qCObREGNF3Hru4aqnvozh+bK49F1AD53np9cgGyNdfyrMBxO09EL43L
gPp2KaqChZn5xbchKxQ5bJEi6rzpQHPapzX7LxCR+Eji5hGc5TEVLKvy9hktD4MX6Tyknvz6cM+d
CongSxxSCeCpfPuLdOsH1ZXi1H7mjuc2d0s+jmXDj82QtikI7qWFEKWnWANcihrPFCiO2nBm2lww
xPhdf9hhmkxoRj3raBLY90NQlsDMx0an9Dg04F5P3VwjQsO80BQxRck0yZ8Vr5T3G7hgorEvjosY
cHNIPDqOMiaQqV0x+6s+UHDgm6MzAfw059JwY+nBM4cSv+aB9szQpAqJiMUPDDdXHuZ593AtJuD9
0vQXwnN2vIUh2Wxn+w2yiTfs6GwoSTmxWnZJlsriAA/QWQkkEagkZRZmeE9qKapkUAIYlOp5pgdy
to/MSkt3/VrvJaa4A7l2HEcW8jWgqKjoIPgJAelRHMsZbSpoddQoQiU1p4eMnorfeJ/vGWX+UCx+
3p4d3l1IHS4xfsEA2EzsON9VvzrlCdzMc9QBPBYw1jVPMK8WgOsRJzdaVcaG67zCs1/pz/FFy9q1
V+9CuYfHDNcGUfiL13R6GF7XepfQTooi8tHMR31egiz4wI2LFqfLuJSMq61UkGCkyfHp2aM5LtdA
T61JCaBvAihwL3qOD83ojrzkH8JiT68h7Qm+yxzp8th+wqFKVJncmIINNvKyE/FBOfuJTbX9ixJl
i/SMGgSnYUbqZjMfFIisqxfKFVoMGV9GzLYEbrRcJinztfYKuhswuywCpF7HqdSvR9WNP2IM0IyZ
JdwqoBsXQTzzRlmNGT3ERqbySiXmEprg5uNpXf2tvryFupowktArSG6xr6rNS+Oa5Zx8uLoYUeak
QJ8mF6OwaNLcXp0UJn1Lhe4am/lCGsybTGMjEdVr9+hu5gFdfuKlHxDJv8Sqm4Fh05OBKhXSQCP7
52uu+72qlukgJq2SCEMhaamuyriQA10qW92XFEJgHam7fb4Nh4ebO0dbeeEJUzPhYsHx/NSSvT9k
NcnG+DOwi2TnkKQHOQglzxdj6BucEDlNiB40a0de1UGcsQ/YBy5JZUOlzvlMddXLn8DGT1c5ycEe
XilJMJVudWahPvN/WvZRGi1u/h8etH3Bth9Dy/xCOtLcRfMzfuYfEnDxa7lPZ3VB0iI84WxNHHOU
Rl/ToCBL2p8FRdB/dngHuRGCcMiDA+LWD1IucW/HZBik7tQHyjkxkbjfcxJjdihx0AjZ0d9SCxym
iVNB7cgrPKET20KGDw2QItwbcWna4Hl2rQKm0LtHOf1hiQlJPeRuuOSsp96pkjNpRo0G2iZgu/KR
0uNNUVuP3NZOiAhxguDZ2lyuReYGQ0R5JzBrprLIAna3kuc3yeSh12ikiooMB4w7vJjBs7lkLYUw
aBWDh84ztB7XaSx8lzYNfoTMQJs3Y4gMwAElO+0yx+2OU8fC7YLZK+pjmJ6rgXuKXA+kwda2H8lc
cFMSfC18nUiEGYQHfeF7e8wklSSWNK1aveFfrXinEymPjJNpho2TqLHeuG+1L9hho7JDjGda4Dtv
6ZpIzqsQVNlUwfc1nupepHOcICtS/+hyuzQBjejrz1Jx8ofgYpaWbdjf7kYfh54CQXLOfDMKhrF2
mi1xtiG/XVFGP/iPGUszWoXqcrpP7m4dC8Z7ZdCNG7Z09b/Uucuo0kryP8H5Q/+VRlmITkCKrNBU
kM15Jg+CWzE9b/bvpIpzVxtr8EsSIq97WDKLJj8Uwf1/wl+Lr98se0zUucJonCptPYkYPswHXLM/
m679mjKE+4lWlhNy8qLMqutH/QoY2/7hNvUQyqSIXWWtegEbBVSmZ3sALwlMp/bC8EgaXvxp9VBG
2H+XAl5DxsquF4JzKvD0UT9hZO0zNeAX+dWlGAwfLwvrjIEv3Si2WcELbp28iflm84DDIjSm+mGa
Yp92+XE9YAAGTRJjKYirbwjJudGzpEe74qQyfMCs4oNG8u8P6UZy2DNi16hA2Wq/yIFGWxBFpEyZ
JOKXleNG2MpfS0GP+/6CeGvfLcoegWUMqSCRijVz30JoY56NPb/S5wRGMM57iCXyb6BHUX35ZUrX
QTj1cQuTF5tYBpv4nIvBffHDqMi7HZfX8T3iTLQvw+1jHKmoyxYCK9Oul+W+aQ4nOi8b1rvVBssQ
kmmsjGvPN2CI28PfXp2rN2EdNf+cSuIzwRmQExSUKcnjoOzImHN9i2d27oMLc7dcXKkFqka1uzTg
tF9Ue/5fz6nzyoRg4oYyK2YAV1NGq/4D6PMn5HkaIQTWEB11Tz2pRrYz39anGnLOPHTpk4WWaB+e
S7fbPR51MMhKLLpnEckuSLMjkRvHb8ESyK3ty109dDj3I6vcaSPLDqYbJAG3+ktm5ajzPtAjKHJs
irVAwetCsCNOuA5bQD9cmRlTeJNyAI9ORLcN5Mw7MW0p2ZFQwiT63W4MobYY1JdXWd+TSNK6Mjqe
KwyWer5jvspxgnL8iMBofg1Y9pV6g1g8Fj1i+COr4rk1az7KQzhj2wzHUW/I5YB5e88rMylpf8dp
Jk1bc1p/jxQgkoo1yqWgGk96Lk8WR/ME/drcrAFO14s7qvJ2jS25DL5dyHaBUa/mzPrxawzpWKQi
b0HKmO8EF5qFbNNh3yec9gcJ+s0jz55xs0TVHnL9Os+GIfqpxfzZGyQcXQVTRzIotqsrkQkD7428
5hrkNEvn919707TVxKGAXAlKPtPilDm4KZDBlm9bnNSDZT/hn8s/TYDcEFhPMv9PkGxlclDmSFzj
frIH5ivad5a1eybMJrYYZklV3kX1QrCIWZMkZL4Hg/EDXYlmly4oKKYfwMeq4GGrRDDkJU7nkotg
mJAD6UGfOJmF3Y8zGB9l9v+rolpu52mS51LhXyYY0GB1U+Nxi12iaWpQQXFRzW/qh/sMF4eNwPQm
pMj9JHCm1/Dwp9/qd2AxNxOc1aXKtAeRPsVNI+z6eqJ41b6d/C/gXRil3+JXI/Jrs5PKvZyNqVR2
ZIeriVHvMuDoNJ3FO/Wh/LAmtlLIMYaX5idFaJNNsEGjaYQPorAfHG9kPYfKZNcrIR1jI4Ea8G2l
ea6PMq2RzWFum3gZlnu5sOSwq6m/RFyDLr2BxsCHRkRxyh8FkirR66c11SSOAQwFaMYTrXwLSqz4
YTcEJhBCqE7ChFWtRW9OIJRYb8uktt0/ckh7x0OZE1QT7Dz1gNSIxcpj4Npksy+MffllQN3i+qSW
/BxcF6DDqBhAPOjoRyTG+yN880Y4xbR/gCp1Y4t+fJoWnf6r4sRn3jSrIXR0EUl2KihJsoPFabFo
sArGGUCX2BFYL/Kwv8mvTgQEkb0UkKtkk5hWEeNyd4IpftGb/qP+s9zvxGFQy3SysNDsUuVJz03m
x4HGLyiiJWztCtS5y5ii+m4BYEweZiSti5laDMMxGxad6B81JCSqayY4Hx1dEy2KOMYNEGCOIw69
5fecAYy6YUnr4/7wUXSfBycndfuZUc2u/sep+VQ6mCdUTAdJSfv8Zs6e1OJEkgaIkG+Vmg+7PeX+
iT9Q7P0wpymefCsrrjmXZli0TQNrKyXmlQQGmmZiWg+Pt+3oOGuSrbXkKkEFpYgPA5flZ2pKxyKF
lF07j46DlYJylvRica6Vl/tlDWxYwZcXgRfM5nZuSi7MUWd9ooxbYZPsizNdfunjly5H+44TqeGK
V+t1CnIE/kt+gjCwvJYo9MD5eUIrxjxs/S5CskXa+g4H4xUAUz+3jbqIQLVbN387WIkIn/0IQ9Co
efR3cCmjSTSZmqQ7DUcoWnPJBt7OJhGMbCSksbIs1/TXyKuh7EokycjvYTiLsLDZqTOsqgYjCGPS
zGVySBRWZETxhozEM69P65ltrSMlstFPnrq6WoF20jHok8CubY/E4MKhRLQXJT1twgucN/InsXeM
pXk2qG+u3ce6sjDmtnaDmpTGhRsNNkvyqIpSvx4gQFMJv6trXLKvN7hxFafL11fctJQZ0GCejfM3
SoUHygt2aquycj66kIXOboLoTQZrLv1zWaufpSSpO4FR7I1WFfls3NBI47uDwC2iQanPlPyUgCvj
x3VgNqCMtp6/qSX02AQOdlWux60Yd2c7+AQ4+ryE6pdKuOVTVqCwCjD4MYTs1lD4b9z9up2ERtKy
L5K1wIRnS0+5HgvzsVS1Bc14OqAhKBmRqB+W4/FLOYK5z0mrAMgize9aLerlKsaN4J0KcEEMdj1/
UNb0LLydu7Tzw/Iw6vWtQoJROWSKh33obKuYm7s+EEbslxVptau72QbZQz75nIzPqgRT5Daq+zzu
RXQupqHqOWE6wBlLLv4co2Wmn7dD7rKXNPVoKt9OjkOWq+pg0kbtF2AQnbY3TJ2tBdx3PeMvyh2E
juT4n6XHRu9888oIJVue8trQrAbe3KikttXopJ759jmuZCJ2a3fbj7zkvCkvk8TLiC62nZT+FZDr
ykdqudFq4qMYourrxn6M/Utko99EISQofPr24Lxp+pSMhUo+upeKlt76AlYBGm5RceEyn0NA0fMJ
YyWaDqJPUDgdraryJz7inmv61VEdjqrt1Q5bvZmja0MS0Fc8wc1lvLHGd5W9QkWzPCt+kjFomFgP
7EsENTWhVe28aUaxIjQxNGLOSy40MRzBVOIVEvSE0Knu9hN5tzz57ukinlw3G1FRmfrwnrzsB++Z
L7WWeZkpUCmiU2HHJiXtEMhUUmxqrp5gh/AarsTtWXiYZJBFQTlUBGPn5evejjfG6NLmaCtEANco
Cf9JZlcdlvZeULq7X0KDP8V8S+YCnmEEmcejrvNZry5TLunHuEJd+xq2yrfP0sxOhNCpd5Vn929q
O/RaQXV+1yVf8i1+zVGSQn0I1S3YcVQveAajNYDgyHim6lmcsAx6LGbgaCOIMNhs342MQyLk2tfC
TKmNc4rHyCFxqv7k6zrUt7GD6q62nVWjspfdahashNO4IPtfCM25HecusAuFbSrKmdm5IaIpeCk6
XrrwxORxi7utMLR3G7rhiB0BsZyecFuvKbbcdM04/ChzO4B4ozxyecf0xBWh8IC0AODnRn7qr58A
+7YmwkX+bB88UoAdpCkWsw9tbX8MJv2+kkafwhvvfGdlPavKW0fkk9/xteyaXbseZwfy/Je0fzYB
nOjnuPECFgXCOusbYNgNnWrkMjeDhoULQmLWBidRdYq2YpbRdr1ObXxtgwbhJcShoU0TzySw3xc+
3vLU1sm8yoDpnrOoG8TWafhKscrIK5TP+GECFdH/GU15i6Ob5t2kIEwe6HBjf0XMLTVxrJeoIft9
O2yJwXAaToKx0vP+B+yhyBwk65A54asV8rcEJzLeaByOV+z6y2POo7E4A+8bVFKuZvHymFec4s9b
i1ak7QxR4ym7SJ71AH9NWYLajd5V5/DKurGkfjudxOqRVItmK2pUakujzV1Xtbp6nZ4zTD4QE0Nx
fPwE6hCylaGnHLODsjINSQCLZdQzhu2gUZrlSocEZqeUQH6zGUt/HzS/xwi8e6FeLKj5lkc5LLQu
Kwo71PBIViINAzFEx6nq0hEaRf1sXxREDsbejl0F0181J1ImRHFJE0bm5viWVJEoBJ5L5dxCPrLc
D3269z8Fc9iMTaL4AcoQtPaQrBt0Xnmeln/3cWzFQFun3Est4gH4a0HjKgF76vYU/MTG46C4QMuE
HRBeAacVUXO5Y+shZC2K4cncYYrIbsC2KPC5UO1x0ujueeqgbLK89GNGk8esE9SwghdA0LgyW5Jx
s/qq4PKQxPfUl0BcUuJ65Qt69LW8HbmPFXo+KjOr6LRS4h9pU2k0UnSPssb+HOqZRMzJ1BbFJCIY
M8tWurHyMhV6XP83KWiUzLypWJLdN/SWv66HgLfm5Ue5kFxshn3bwobuT25/+Py6J2EZgV3SP6QO
E8Kp64pv7Ju48+IEuhrmXEZ9eTwwysBg6ynZ93wirwt87LckuXZXHSHBA8fVXz616CGh2pNZ3r1X
MdQT4H1VQ7P5vdS0UmhhnYCt9x3Y/gusKnG97scvkBhi5hHJQKwo2rCk7n8LRahexQc21IaIN/Gk
kTFMONL0ZlkSxU7dUBf3JHAzcio9s+LtGGliltV4VQcbiQm5/3PxBv9w+gzs1zd34kXABS9vPoLM
nYOYAKEetJ15MU4tA6RM8JXAAiNkbKuojEY6eeGuvrOdeKBcJjzbnoA0dEEmRRHcIA0PbzLZ3cBW
Y3iVLY58bTR/Dl524mKBf3gBfQfTP/MWT+eUWfqk7FHq+F91rAfLOIGFIEiKwWU2poCzQ20E48Uo
uPaPzyT5JlWtWC3utu+li1Zpjqy9/ujzHS/FOy+U9OCnbIZm06U91lpnkPvmvaKNLSxurP5T/hAN
Tg4NOsC+gOBLHjhxZr8SlTaKBOyfTe+nznl5/mr8tjki5y7keN4QjFI3SGpOV96klCc4tY+5nrHi
NihQhleDyx2u1kL6V6qxhmI10Z9x9/0ELl0Fh6yEUC4gXiVs6mQpW0Wkxbr0l4HjOTtV6gKHmx2H
n8srkXyzuJLSf/yjpY6C7b19zdSpmSRNzaiuoMwbEUlODV37M5x1Qdf58qdLcSIOoQ8WPqPJWp/T
3nJJwpHOQb+fsNF4KsEIi5Nwi2R91rk6OLyu/49hwXDxcpDu90Rduad1M8G6/YBd7PIZK2BaQExq
UfDK6eB3c+saF7ByKzOIo8NDbtGe/QKy/cvreoIaPNAHXUbQPbQHEmzm2hHL11Npx4UPxqwTGOJy
PCU/IywMJQje98D2OXtYIxzm0S1bkEvv+zX43fD6h2hEPSQh5eYpRLzVXsq/IQY4m7BYkeKU4qDU
ZrrJG+YYjoXqYJOb/nHhISeOsegB9ZzYhl9h8esKe9ICRKcSjMVW1jVJXfh2KtJO2IOBKSWle9xZ
M9H50chcWczxrpyUTadRsiOHp3nVdhlG4hGGdYkvg2mI+nTnCDaTkW9339hS6CmlDEeJSVunngrO
MLihZk66LDln3Qnq50c+ySQ7jc4tkGFG84ONgoxuwuyBnCfcaWSprZnWKRJ4tCi55rdCIIowM9j+
inqZTVOH4j5UH5yRxuZUm6hJOJ0hxJYmctIF+nudAO1K/wNUzM7+Zra/maCYxu1ANDTYbzbmlgbK
q4VIDhMPbNUNOPW4MCloxX6h3tqYd02CVSXpD/kr/5OKR6aAbUgAtfXgJtha1bkz1DPDE/KBF5Gu
Fh0PR2rEH1XVqCDMPwDr/VQURMqi+BFOZbit74/WFXaRNd7tE6V2hYSsw2UdBtvPUvpnsDwBRn4L
2A6/4p931He0r57O5g+Wa+8+g/izacyfMdSKnFlTVjdT6Gz9lfYs0j0hI1gyiR6JeuAnnORJk41g
gjH/zFC2c6J/Jy+Z8s3a+BkCpXvC4D1XMrLE9RLlcZUNTuSV/2Sr9G8wraxZtGTB/CuGcPaFIfRd
p9VfRpcbCiun8c6YEeovx9BWviio+LxaQd6iMeaEHsEGccH+9/sMW3AIxa1wl686kGxQ84Q10DHt
8k2TONqP2eVb5RNoVeuNNtqND4eVb2eEuW4mphi1+8FrdogF8pR1eCyV7d3dpCiiQ9w3trLtICGg
6b1i6gxldPE/Bdj4PBGo+s2mdNvcQ5LdpbTElX6fgSOMNlcIuHrA8/bSuVcxBwcE6jmFxUfs4ger
GufaEfIZBegLid/8nvfL3ytm8/W7kuXNLrXtpb4aWl4mwcw6vn2I++VZ0GGy6ijTLUGR+hfgl2QA
3WyHDTn37OtJaNgALx4imhZ/k6byHd/yPX+9Wo6bmVx7yWrN2Tj2yHa/55ZdFy1zL4VNV4bCGwFa
Hq4MTc85hyj8OO2PLB0VuiUgfJny/GuQz10OR9WI7YamVBK1o7dYIzg6VFg6z4Pvw3HXN2h+dHvQ
cGwKYNdjAjgYKP0L57/Kp9V19X9ngjBcTMAoK2A+qzvs9uGR3nZYei31biBuu4pZjLq6osXRWv8p
Kz03K3uOSy0E3Zs/7kV7OcPP3abXaSMwN8s7Rb2J/oKAwgNcmfYf1G4G1lF38RgA4kcKqHKsL2ih
I2/zwurdmdrUNTOq45VLBCDNZAT/u+u++99Y8LDeCxkalHDDfcSm7TZP5WD2uX9qnWjEWkr3OXWk
5S8dGBcNk1Fe+3LEBM9VDak8hpf4AX2jXKkiiWYBTGQvNRH/3qE2IKcAP9r1NSVbPN7bB67bLzu5
0PUQ/u8uItRuNwwy0ZVtJygSzNauBLVikfVxLOFShjIoQb+meCNKveI1+1qbA10f+ZUmUg8ttOk7
DkoaJog8FUK36ySheA1TFn4Jz/KMzE0z7rO1rszKQYlFN/8eJK6JL4FdNu22mt9mDY4+5QfCE4rv
cTNgFbb2B3QfYzajB8O7W5jqhsAZjtIOSaV9Udc0jdWudZxshzHStQx6l5NdHnqk7HhpLu7zXBZZ
/HaQ6gZJjbwsGKIpY8GcruL2SaG+NMGnE6ChSH83zpLJQpYopyQyR/MU3S7yD55vHAsnLZ6w72Pq
pdMfx/Dvr2BiENoz8qDh4/QUy+CrC5+n6msKlipYiPS5E717Bw/2/OH2RS39Tf9BGkFZgzk9XvNU
yQWjYZa7yVG+HSTJLFhZ/voNqd1qq+ICZERmOLex7HNGghLVsdr5BoDNvjOQPFPfk04SmorjvbOZ
rzIbejZpjQiM1naFfSqdkFEl9OWHyjUOpWfLndLYt93ZsTSShrzEawD5C3Oewq1go3ML21392HRj
Lmn2TfHrEyv0IBVOkSj4iYrT4IhF4v/uSdXnwSVWlHdfsIuJ6hnnCG9qvjEFr42I6GZkrPqnLJn/
3mWcE2TVivDZHFQKIqsp4Oim7JV+BGNXD6VpCfad/mTU4bUJdVZ0hN5mQdXBx6crbbtoRAjLKkp8
PrKfqeypSr0EpJG/2/zNcDVGQwtRcPJIOh7nlcfF3JE5iq3X7i3m0FSYmyf6iC9rFPBBspUvt/vV
MjyVvkc0KdU7Eps4rSvKDqjUHoDuW2ac+91zJxV9yaDkzZGm7xx8cKLJ5C4rCTw+B09h+JCMvwp4
rwd6jItkwG2NoxpHCB/XxxtIcqlOWoOxtAar6emUFcUGLa/4yh4szwR87t23TFbwkq4jeEnMyrYi
5zKmq3outAGimbKVkDC4zhX72DCILRyHbCHw3YOJfSt//uZyQmx760Qfh6eefEMkXA7SimMgJnU3
WgSG4OHTx6p8UfHuaq1Wzwomc4sAeTrIvtrjvqOI8GoYPsRmvPZAolGRM1ocmmcjyB5upVEfeR0T
piOxc1vVsVo9FuHyLBW9PZ3S1/sVxnyOLeYvTM7UuljPhgyGSdvpgc9ybZ4dzvSH1PPt1Q/Fr7yH
GJH94ui4tU9pEvicb1iMyvzTHX3JwQH6JgG8r9aV4LXJOz+7kpDo+j7eH+Uka4vc8wec3c5unMJT
A5oXq9NablhJ39Fo0tvxFeRtx/WwUUJnVefDdG5pDoyaCMnNG9Xdp0ruLqMwLVS8dUH0aGSJj9rW
+yQsA+QWBhHA5UqdopjBO6ANPe1tWC9arh1WVKcom8dHyP49BGcLvEuzN4uUlyh/MFLudcnFCZkB
Wy7/e9PESlGpbz0Q9P9AZXjF7o2/JGVi3Q8xYyChAXyl0vKPaPyvDjCLOdOSwJ+O6yGhLyEYTp5z
XBTYOy4Y3K8qEovxoumfQKz3Qi0mr9qX8Fa6j8Bx3/kvPXts7S5CMque47FGt/WB6/RECoeLSv7/
5M5T7hwCnJiuZ7qmIjtf75x98wmovAU4fVSOjTq5dhLx9u48oxBRLXZ1U/WfWIUiwjHA+FkHxefw
wKBAV/pSme03mtP4IiTuNpqCpHF4X7v6k5+nm+YgHb5EvMLY7OP3EhA2BACN94rh8ByNPVBtDH+X
zFkbkGRfS0S3nPQ4erjPPAJPs16jh+gVbfFVMCu07Fqs6qRu7qvVffzgXYLpCdkMtfYg8W1Z9rfa
bRwSfV7NdgTskxx3xt5BGyrzpZtyhNo6icKBDfWiCFctOa2YEiyn6TD7owyh2O4xmxhYm7/TjhTs
ROGuD++Fx6tfMIlquhYZAlDfe6BlAzwKXQ/hsxEivD/lDCjIxJ7QRtv8hwqNTDRTLWV8nsWvRKKr
7gJFecQr2o7MHU82RYuhbeGXKsBIPHZT9G/eFTiiNDCyCKyQfpnvbITswEn+/7mcpnDfL2UZ6TOw
Zu0JFEbaerAf9lkYkKichKPQ3RPctwtgZ3cNqlBzJCvUe5VUB0uH9W72bR7TWGXjJAa5Ys08WMAi
B9jpHLIYQih16Yh6O54BXkOnNzh6vN/Ey69FdN5RCixtAX/KOD2HngU/wUphuatk4Pp5klLU3mH1
VqYNzrynj4Vg212hQNLPfEvqKZZNNXA66VrB8NdbSCKn7JIBjA08ko6nXVxuOg83neSSZFVav7AT
8AawsqWLr6PlcYqaEVT+kdhP4N9dVGZ+hxF0pWpeCBPnqfMGtX+uTBqlvjtSslWaryqWa4O6yON1
vqn+etuPzXg4BGBIkYLoCcIQycAddN+8Z5AUCSzQjLtNAS2v/PEc1Y5X7gYqrHLL/ytYQYuaz5db
TfVhrRQ69nQlUeD5UqZQEtwnUL5eXyjVkqIckCkRIIdIgpv0ky+REoFaplGJHCN9ATNntyeXdaDz
bR46/ooKllmyRR/mST/lUj3IY44RK5XFqjQroaJ3Y8rzB2jOoAjmnoggrFfWYfmSh1qe/83gA9du
6G5yUdyz+c31EVw+kfq+TVgTcjunCxvfgdUbhAGMAgZw5FAh8VmSiUNBfrvd1qmSumsmG/n5C8iq
0SMmTPLj8Bj0WvnqylKuh36EMnWS2+jnQ3vAcL2XDAizaqLCvVjkeGNd+KLI2YrxWbXJabhWDIl6
uloeexi41qkJUNu3Z0RRp/1PPjkYQ7EVPV5+3mFUObauxi/fz0V5Hg+oKbfBfbNagGCCZ4jSKxXx
4ZSZ71ayVws1qLXko1hc/QaZqb5P0eLvDBE3Vgq3chZei4A6O8GAoPFH+sOWqjpQHdqrUdoRxzEV
wK6eA7waal/8js8nw6jcWOec/kKeWY1hSQgUFP0G56Rhs8L5yJ9G5CKq06dITMwK8+Z43d0DoyVr
MoF9tKpKzrn69UfVFbyYJxeI0J6WC+SftszQeCrYVUHvPe90x68rwrgJvfK3L2ihmmDzQ6yY/TvZ
2ohqOP0G1s2B0EMxmmf0QuqjY98XGyhechgnamETwkwY3PyhwV4iMSYPfaI6zHjyLWqjFdCAv4JC
0HW16n1nrOn9eOWNg9Td/De1OfmxJQzRnmn6XudZDdub66dVrINCw3ErFmQ5HlYm8z+7tWI/9wbq
ZgHQtq7tHbzaLODjm5TKY1GhWLNin4r6q4U7p3+cx5RFqTqldb4QhB6YnGDcMaZGuUd2DI8POEkL
JCwyRUgmpMZfQRquI1Qtj1w7Mz6FY4jgfb7pglbd8CEyR3wKtTUOXZhM5b9xjh94kksEPgq1Yt3s
10f381z1HtxnrA/ZF5WLPIrzTlh6DXysL3Rxv/kOYdPIXQbOMB4hdGMYANu08zhiE/PPVDLGBoH2
eXLx0NxNxQ23olVjtvlIQE/1frqIK9l0WOFWJt/s7VwoxBZQYdu7Ql7yiYE+XkfUPWTHaDnkgSIX
x/t9HWY2r5YvOOleZy/JAMcLAFOUKKeDCWlmemV6tPoYwUk3rizmph7wITPCyZQuIu6cL/gbCvX6
50JPYQ4gpTyOQMxYyTiVTSavg0S27aRW2i5mAuwnLFdbhmAprdB/jOe5XQuecONOUa+OZYlo7FYW
nBnYouLdfwB/VQjRdctwk8lfPYHSXxg/Hq2gjpS5jyoacBbZ/YL+cnpbzuWJi4focRM07dpx7tL8
ISlXqud33RGDR1TCyb2Kffe267ObH18FLNKszYpHDFt27ppS6roUryVZNmgN7z4Z0TOCased8RWB
om56FXWMRE+48dCftNOkLQkiSudgdi/uYaDYgVaHi4gSQ0a0OfRol0F7RSrvdwjK2RX8fWZEpWIf
Z7tLX5SwxrR59HvoeuL9U+dPvlJfI8ZuejibfSr5mfflGeGeqPGYc7JZtZhnuB3OjgUYNIPNns3M
tnK5IfWLOni2oP9UIbQlHaTygccgtwvpta1vT4ABIMmijLIM7g9wD5hW9r3iHPtmzBk4lGzcDbCW
zeRBwVKxXxSadfPSdmHXVGJJlD1aKS2THAaP7DKzriSn6dB2qAWqOX3SV1h13ndUyZUOXCAsbt5D
n7/x4CHaRh/kPpegdhs8IQusm+TgKR3ka0Uv5/pm54J0gLcMXk9Jqf5He75eV56elqhNwSqWeRd/
d9qvKJ57/n1IVj4V6K15r4oi6XKZ3k13TSiddVYPJTukKY5iYmLgkK80zdqq3NK/5VaKXFhhRRW4
Dleln67QMsH+IT+FFe2jiu6HjT7k5Z/DWP9/A1TqIyGZ0PjarWPP1zkzRjh+auufw7YQZ1GrYZMI
r0PBpvt4t4eKiJSnObqV6guqqP9d2e/FdbokviUKruZswmWLh0QG25o+PIOL0oJQD0+2x6ixgliI
EIV4COa/H5gJhU1KglPwVaxefLdcjWxuMJtyfWH2Pcqmd0xvH0IbdtsB7uj2nm+jW0FU2vLuitiN
YddbWEMjKKQqEAm2aPpwz3IfVAkUymVSpPZ9bA2xDLxJtOdoM7vtbuzVWsePGmNvA2oUNcNnjQHH
i9yzOfEDkdzM/S5EViwoJ8vgo8nZt87EUZLOoKQfOtq9gTwZ0H8FlfbRH3CxWyw2By3BmyyBCZfk
qGrVk1eE67Wo/IKxJ6pH7HCSwQeOzT5st+FKVYz6ktKCMC7iurHGPlT5a8QaWIY67AuotFykTiRQ
Ts5j7BZMWp12wKWTCDqueAuqtTMamsShhDho3hagx9zVEQ/SjVkvS5x9tP2AL5HyrJXGmzhnCg1n
N9x8LFNpdr4I3x4CaPXd5wiID2xWMzhITbtFyLcDaOiarLLtwKADre+x68h0uLYpEHvnRcN0F4a5
wssce55d2kKQBsUNsLR+41MuKnIDEuaI8w8XaJ6tKu6fzDtGagydifAfqM/zYAQRwjGTBl050Gi7
lJZTw2SMmxXcAnPBu65XZI2xZoAoo3rlHtwsD1W4cYAiJ63YXqBepNGM/azeOMJy4fq3IwZZok6D
q0nH7lHrp8Y3/t2dIqeHrPo7rhz6/4WIWkmHOVunVSQKaAsDIXK4bfm3mvxdjOn7KLBpk/ozTRVh
1BF3//ea9kYdUyc9QpVPPEnw96bNsyvzAPKsuP8qui8+VzWwNxFUsx6rLfics4VIe/Zjax6atDvC
jlzLy+USsoc1rwTQe4GoKI3hwKxYiXNIV5h1PjNbC9sqJZKlmtPAn+9NbgZsViRVm0ExsZX7hrNE
heC7+KKKoTBFzFrVqapegYlEEVpntyUb4FIhXrkPiRUaxp5Uk5SsJjJVRdgfchKqs6+eHlZ9CxnW
ej5L0MltNLaoHk8TZiEXSFOKM3ppQQVRq+Z5RUyeNPIyG5j+r/Z9esxeBJPvzVceXISAg/p4oI5q
N7nFoZL02aYdaSNoZdGf22nxx5Py3Cc4sq8DUG6mWrk/8PRnufPXFwEijPqBPQrfpIumuGT30jg9
qwv30cl82ACelhhCWMIsEVJ/XCQVBoNn0FuAtd47wXCI0lIwe0QwskUzNZm5Pvm5z2bHj8gHPdE4
wtdb1H6L7aK5oek5QziQgHryc4TUPRPIU5d9VOVVbWQcgtlu/dnrb5ZMv/5mfy5EP0OnSB9I5Q71
w3Rt12cZ20tRfIMdEArfHXyXPAw0q12MBDew9gasMstzDrIGQgVL/g+tKTqLJtLXGCsw7mEA78q6
5c64WLeIKxS5SiA4Td6ekm6yEUtr/gZfaTOF68Ln3MaRoDtMkDxBpD50XsTl/kk2rpswZRFODbe1
XmQ6BVUHRW/pAP21590G6v6kTUVo6g17fqxqUgTeZSHoeWfwBKd6+3CI1AosfurhKUfng/eQbLEg
yQbr8iOMOJOXqxhMlJBKhAQbcogTpMzDv3gOyuadA5o1hPimzE9dEdCyH4Li4LIuMg8iL1FjCorV
ykk3Mz7jyRh/x0ujiip70HoojdA4xJXSE/rgMWnmdSFltRh5EoDAqpRRW/MqIbS5jB8Rak/7LDg6
sBOioBxHwZnoBXmarThE6qOYX3qapd4Y2FsPPoZkyiozpSS0acjuyaObjbPT+Vnc6XWy5EvD/qUS
jJl1FcYocL1555hyoAqpe8Wcs8j5rQSXjIJJ9+9YdKfkv2fletgffY606J+SswunBDzoU8lyBhq+
QxOFbNSpfDBk3exmM5zwAsEH2H/XzQHf0fKI60TRDCSH3eIx22qzcjLXs7sRkD0oujM6J62JGI4a
Ygg4kqGKiIG5tKijlFYUwFVOfJZq92miqvmpG/OrpLtQ1QAcMh5FZ5uNnVODvYSKw959tjQmqSU2
usY+elFS1z9midweNHjRI4m7CAEhXNT8J79szSf5LIMoOwkkgaGwzxsnuFVqLHCz9/fTtbgUEW0f
L9TNtCEsp0wW15AF7WpjPMmVDtGolpQFdwjDtnj0F15nuK4/0ktjmZBaD1dwnF5nWtZNo0k29ZSl
MBO5ZbJnTFosXgqvMVzZAfad5V6L8t8ditsjHiVdTiLr/4u2k389h9SkuO4Nde55wGtDr4rCFpu3
j12RUs5T9HXw08wZyF/AhR8Yz/kiWVivkj4VIFqh33arOKunLoJiwesa5ihlpUo2jm9du9NQcy+O
Rvr/Qtq2n59JZlDmL7owGCkevoLmLcWDnhJZ1mwndVmCijM+MUZf2GW2PPfpfJtE09xR0L6RPl6I
FQFUfoBS7Vt+Vfy7k8kqeB7Aa8eDFN/srSF4metrP71bcfwgKCG8X4Hb5lCHkeabB4rv3gsfScM8
Kgv/zLvS5P5HulWaZkCsLSJhMliPrqW3o8f7SW7EM+LJk3T7f1v0PcGSfEbniYAGB8SMH6q0gCtB
xnYKCLNi2JczkpSDPM0dpuXK/yn2CcGVQJbRGj6KcZpVlOwSXcNVY0aGwAXvLxOozCpZc4V3mkpL
EmTXC/D+ERDKFx3HCbBh0Y7wILkRyXGd07BVEPaIMIOeVb2l4NAeESM6++6EbrSpV3S56yWu/vf9
hk+QvKRAcmq3RZwJII+a6zK1vSa0rv6b7JQjoyfRDlx997PWq5K7OpJJrvkGrqyfRebV6Rer64tt
WAv7sxRa4pK1Gvjy0nrWfLUjLQCL6C5vRY8BBvm1A8ua8TymPnyDVRzNYDoL+vy0Gnxpboc95rk7
J8sTincNHr1PSLSNj6r4NfGTsJXJg3IIaM8AuKQDAZgzALCpGJcgUHgxrz6M0nwrHAHwMMMVjFz7
r4QOpNuAvBH/nmsofszG0UoE6cMcs7w+IR6MVgF2VGrw2lwvrZCrahyZcTimptsN2l/l2k8woNdx
hmrGZPEbUo/+l8qdjMuePmzwNHre6Z8h00KDBisDCqfTLP6Vvgb7z+9mWT9bUUCx6BvTVmK8uhaX
6SWptBHFnjP5UIHcnsgug3/wMfpWRloUYLJANGRT1rbb9TS8zcvY2vLlzC2D5b95hk28AtR9iqEG
o1o3DSHjelZzWsaqLM+4+lukDV1LAyYc67zzPelPAyaddepPOBiniSlakIYpTwnSGg0Hm/7TEFSR
T8VPK1FlNODYb7HFWXQlSsaEsIRxUboumgkLD69EHS8sq/CgdnTcbH3muNuV+Hb41Hb2Y5K2vqvf
NT0FRjpeUPBh9EpQUtk70O7mWci15k9sg2MocRHPsYqkTZNn0TQnsVF3Nk7Z4Il3dtIMC7Z16cTb
S3qmt7eAKYEob5YjEBaOXG9ytqGeqtODas7/0G/OkAYeAT0FKLnPXDcCJ6i2bDgi/WvuEiGOox6+
x+z/Rt1KCIqymGkzHng+drd5dXWm7bTR+FIucEK3PnKt1WrjyFqK5UglBnG24WixIBRCgmKlthT+
rKzJObmDfmCAFkAW/7VFEsVqF+QTWigp/9rE/fhDfS+Fblv/j+XvlguDpfJqcD9U+XnC3cSY1SVH
GcpYO4Q3bvTiyHLjD3PFWP+vMFiDfUE/sL3BjyuR/uE8q0gE08+WuXLmJ3IW2o7vYbJOeBHEl/sP
n6AAK+bOqjHbXeCuBBIlT1CgiDODtZlYUppmMJ/z+DarSW+yXXAZKUoCvNaK2gu6eg+96/QeTj94
RbTokbH3Bb71erVONzsDQDTVTOoV7JmqI7ywXi3BOAxlvd/adz0DhicOeAA9bNV04ynylZ1WxGJQ
enDUcbkQzBQLxaUzq4+/rzPoDhUgz2HQBP2FQ0C5WwelZRu043tOHsw7wSeCXFTXlBKtpinfXVqf
0gXxqpZi5CtDqZV2pUBslvDLvN1UtSeF2acH63KrDfT3neHgfLOrO7YqjMX6spR/MlVx07Q+lIAI
UGMODQ48SpjndeQIke4CtdkBCHWmaNOWcwA356WfdDyRcBmynO69a7Zqq5iB5/7OhwIn1VvG59qM
gjgPBuf6cLVOOdAtI07sgHF1O/CflzmbnBAFuB1nraCzaSBktE6U8MLGwTmEchgiRscK3uAcFjGJ
Zn5Ex2l/+wx+1WzRAxz4SO3gbBadpEy5oDrDYB1xRUe+FJYucUUj5yVrwcII3CkNLshJRBtqj18u
u6TDBJQ7Ksaj6TDDKtjMGmiVk3iS4E5sniK2+463WMfptdByBOTQ25FIiWiiY79oXBOW2nPQ0ABG
H0c19CVPryUdsZh7I1FxjOLe0wI3oGcd6LH2Sfhygzv4ZyJ4ESX+eGP6Z6/VoFlb/ElP5LS6DTyx
YC5bR/Vje+E83PHWoPbzyJ0XrBtqrezRWmWqN3lTXwm/kZ+mOrlyWu2HryfE98vsmKGLWyYOzfJL
lxSLKI1IsVYHXo4bl+3vFsiuVJiNDpbe/9mVBMMC4BU2bIkKynoRJqCgd+Jl0odWb7GLVUS3/U9j
zjoyBYuJGlk3wHCpLefzr6jjTi0KFXu9nbjfAYj9IRxWpQ+F97J8dyAV4EpjAJ0yTU6g/+QvzRzI
pg+1FfpvJm3a3hoFJekl1Ssb9hb6Yz81iFcykRs1XdMJM1icbEXw6fDViA+ftMD6l4zgo5FsBait
5yOjFzn1DnMsqN29cBL1pQ+WH7v6TKPT59xYEGT7u8dnczJXF9xPrEh9qz5u3welshhtgEdEWyzd
3AEV38kig6St6tlwd6BAHLoGfGk86QTWOcOChCrhsB7Cvc41+xIXONqWQKBS0NmmLmkyr86q+oPB
8QnRkMAYjfCZ0RZGqfqVsfVPj9A4hZExk23BzIGPPFzlMAAmXN/Aa39yRc2O0EvvRpHqAz6kfhPF
KSAxzRhHjGr+Wj64S5OQlEH6VVLmnKC7cYnNqwS7G05xeW8bZkV17X5bMYKFsxlBfE2ftfRt46A2
5aSJZiSFZtAyyM0+0GCd1pKYeioT4UhsegBbmzmkL+LFGaLoWjbq6wPD7nyPi1AEAWZhfDWJbFN/
TYiuC83tSIoJRzqXVlm6aaT20d6viazSvBpeRD7DCzH7r05sbRUMlYKW85oHZ6aqI2+Fvgd0LOft
OovCpA31oIQ8iqW9Uyc9yZx+R+4NKiair9mrYfILWr3kB7BIQN5Y0jyQlXLgJvvlUkZtxz8t3Aca
vS7SSkgPb/gkasatMOHS4DxEnhiO8YtxG6+RCXHU16AiORkx1yGzIuojoArFB+G+s1g4zgZh1J6Z
ui4NLkJLgX2UZWBurr0RoywrRTMwQfPubKuPUcruLqTXaDn5OinTAHyWFUrAd9HOhztTJuyzHE0u
qmZoTYDCfFhUmYZzvp2R5xvru2LFh4aueTmUGEP04P2LQD4eI0IL2AxCoNIOCylNi7iUS2zEgCAi
9KUHvx0DcJn01soIWDSOhWsddSIcV7ZMpte+yIxMPX7fxhojBv4WWq627A+mVz5wmwogGNzKq2Kq
d0fH5vtjkshYF4Td1fgyDzNc/3uSQeICTUI7sauXwhmOKZgsH4S6+Tbmoax/4eSoeGbe6dKxntVI
AVlXIsYB/QLnH6ro8j8BqBL4XG33WM/Vro11ojo51zph0z0ADEVT4xs1GgJT7Vb0sQFCe3WBAX+I
UDVZFoyW5DUBRurJYnbnfNWy5TFpy8ZYMob7nANIlofxNXch590oZD0xSewDXwoLZwkE3TXKXjme
ITrOh+7RgNWz7rPlCiZwXxVp/QYO7+DQ4QFHVjm2eSEKRWN1lfjxCj0ULYw3vvymbsC41cLtx4+O
bcbePpU9rIDL4QOeUukwYXZSKmJO88mwbsts6gpzjWDk/MzZA5wfKkJJqkVkxx88CyVi32M0LGWK
9BtAHtZZQ4VwMoPIHfU2Rb6QPUdMFFrYSezIjBRHo6OMeg+uFISF2XztqJwThuvCR/JXieUM99KJ
7ykz1sKboX3LwueCmxlxa6vcx6Fh2/PaxiKwQjm0JeJsXYgqCTcdi0zOEHg8Nk1NwHgprtKNTt16
CNd5kyAcZONrIBwhyykbgu3adRP1W8Kvr+cH8xrekfFEIpdQxtChwio5Dl1HEYSnW2LWnIPaTkWY
dEobIwRkTJinyhuK6YNJiyWCoHXHWwcYK7sC01XGWfxTJ1CxpCTFYJtMz925dAC/sD/QI12pABtN
KTPlBo8NNb0aIuqZGp5piJ2Llt0E3uni2AfN4a/RncjkcDRoKbsL0W0nBrEZ8S/mjbl6vWuhwuO/
gC7IyQQMzjKH3nYfQxpfihK24J8h7JYJwCE/VLv+Ba3LdidMPIWyqbUwLmFqNfzZvuNqVWo2yaHW
lcHIDmsB6HactcDHbq+4LYD72hvdVVfQoQashgzviK76VLMPm51eOgD88XfwZVuGU0LBNtcnD11t
xJuLo3pyIal3QsykcLdiZ021pk7diO29yX+xcJ+d/Qb+w7PNezPGD7oXsEAouXssWC33O6rsv22n
hqIqXQN7QSN+TXYOBT+OQ89rZmu7BbtSJY19orxJdK9xxsTt+sdlN+enBrg5GCbC1/zbRyJv+7dP
TeB9mC8hcxb99jPvdH4HYkYLhPN/9so1YfDO1l2AQiiU5pVjpfdnKbta04KSl/k83M5Z9CEbYZ4S
D1JOU9uDRvjNay3pHLrQnoysxsfCqmbRa2GiSb8okHBMOdORIm2Upt/rF6Xg3UpFL/aUb5EQ5H4b
bS2boO7G2EQW78GxJL7SmtUdUEbZ9yqjnz1c6lEuillq8pyIkkIlKDi18qUZ2r1H2pZ9PXAP5gsq
RalG1S3xa0KLOwb9OYI6xFnD17IktdTaFmRECHkiO+TnaRcFBBA5udboKqs8ieRfgojHH7WorK8y
Dy8bY0wonxTY2G3bdn18eM3jTJj//AyYNo4MIT28lmPcH+Ma2B0PPHlu3WExMYKAf1MWOCveOVVh
GfjGH5X1OjwVAz75v53XXHNTKNosBc8o3xOdbsEBKw85NQQV3za+BIl2YEDUHLUZdMMINb/DIYu2
2a1/XGiAyK3F0Fxa8ujZK7k2cL68J34rmI7+L0YSQeThCco8IXcld9nuuxAZXet0NxW2EXjGSBOj
tFxyDCPDVZYQmMX/Qc5oUyJnvRbPTTMaLzJnXwuLvWVIIXKX5XTHEmRzY2YagKxRObOHiZhgh4NK
RAhWPOIVC4ABnO752VAZdjePzpj1XF+7pdzzvohZszZ6iWa/1ix4SlCr8vfhjPet0CZMnJugbs/2
WnD5nX1wkBtnWgf8SN7JHLbADAyCpisW38F3SbsuUnEZtfXS5V2C+YBMqXYLYGJwF+YO0TFR0vCm
SzRjRdZtabARECjI/qevczc4XyK7YFx+Ni6enhDU6RkfT1rO2vbTlpFjdaqoWfxmB45+tYV47YFs
m6I9ovy9C237GnoPFiE9KzwfOtlWvnC51ZKJG25n7jnAMoxpGOZR6S1oQ/+yoz8QDek/lTOgu/xC
F0EwZGQFNd3sbA1oMyEWq//7Yj5xpjSg6VFP4PBca1wCBGfFYWe9kPSa2gOr4Hzxos416ePtpD9z
iSErabBVkIi5If2+G+Ti64UEZc+x+fCu0BbkkoJB015BG4pCjxjoELKcKB+CATwPPSFmgSZBDVkC
Mc6YRYJJAdlOP2CaYLie4LQd/Fm5hVcQXFbffzPHKy0VdFqO+l+aECy5lNoD8b2HcoaAdo4Xs8FZ
vLftpce6eYqRqs8CS2gb8cblWGspavGf+TaAdJfhi/jM3D1T6BjE7GZYV4yfKcOE66toorQ5iksd
U9l7EEyrK0/7+JLYcvN4uwiTKh4XTVhCbj+IvJJnEdVuIeXmsd0x34ZsOfOPDS/4A7JZULfUsr08
Ra9NwY9//m8yH9vlwo8yBquA59yUJhx1ULjBVbooV/r3Ipf1DwTaBKEP0w1YoCbB1KPCO8UM66GA
2FSEc4/uXevcsZtvwvzAn1vItHaY20hf4U1FVrnk5tKL0Ihb1GT639KlhxI9Chl3iiKiWUyQo90x
hugiIuw8c9X0R4DwEX7RqjXk1KylKXxMm6N0t88501EB7tecOQT3gU+hAUPIZB4it5yU4Ne6LJX1
09qcD0MIrxa4/BkZ1qe8QrdZVv9niaJZz1Vp+5Z5nrS16FdSg8T1PIV3Aybk7OsqmXxIHV116wK5
GHaQ97oKUKXWj1M7jyXzIkzbHfbPyTuI7j+1lwRn7AoKwHuW6eU30dLKmzxJtq8AYLSCB06uDYfj
fDIg3j9bpSX3dLR7ZSPCrBlSps4iX+UQsh3vKcPfhWU9vtSgGpgmWxjp6MQlV571VENgpYPsr+ki
7U2aGs4si3xMXLT2+Y6JcfgeLOYrZu3wkJ9jW7WUymODvzqa2gh5L0y/TJJ0Uf0eS3hIStw0hPum
phkIK8WQt903GdQdd9xBscXpgcMBkRlMo9QJ5RecRSyycNoTIqbBPgc6U/GosgBY+ywFdn+GDaW/
l+3pfE0Rx334JFQ87HwiNJ/QBSlOqE8CAqsriJy7uOK5HXga1tFhP5c6zp7wYMDQ+SdCbMAkcSDo
w3dvBykdrxfmFHmgweib7IaWEU8FMo3MEs1Hoqa/nqqjym+tcdE/VZ3cZ+mcPPuVgaM3DMEN0hI4
5ET09CkzIhCrM4xJZmTdIY1ZmI2RNlBt8EcrQozE/lGEnnAKavb7cqNkSMF5Qplj+v4ZyO7Ng7LJ
2d5i+D1odVSjTTyN2b7JlnWPLmdKbvWdoA5+E7jS70U378CWigtb+GpkjeNcIMJFnVSOydc6EIlw
XP1pLBcvbE/yzNMYdNrTElf0/WRtUSYBQx/6Q3HtyCYWix4hG4oe+ZD5Zpx3XbsnEeIIIKB9J1tC
MDuyLUwFRPZYkWnN3Krqk+Ko/qPbXaQehxqI7uVh5lcn9V4hdBxq+zYpeTeleD+4G+Tv4mjkdG3M
JiRuu+SD69Ig1iSkQxKCOqOIYihtKMyPOixvTuF/iV22g5ge5yMkFB0fjPZBZ4bYZILgrm8nhv21
HyuQhqmydDjcQJqaqWtdFk8qrioejrHDO9920rES9EtATp/yHolQkoHpKGHcDYbYNSu5fCp6e4P3
+JLzZX+qXmPc9i9UI8dM+fBpBoppY2KBZuNW+6KmWpZoIe3YmOduHiS/RjVsIAtLp0CCf+Sbiuyk
sD5FJ6bojPe/6PfIxqzo2r5Tg7p5ki7M4Jo1VKGCSGG7tGdhuddXQNFst/NTpQqQ3zor/YLFNY4D
obsMo8p+9BEwwaauWifNuLn7bZXUbML57VgbmX6aZDVJcIPNiZvRVqRT1UB8NnM58bsjCM9Yi6tN
m8787HKjTMeU9E5A1jiLYdLs5dt1rfS7C8uUaE2IItGOHQQjO2CfTlSdCWn2pA+iVXGt3K+kuSR6
Lgho0CU1LhurYnZRBGr+X0zYArbwJ67SXnhlHJ2K20kZLj7WDF3z9zP7qwZhtq/BiFrXp39klQ5Z
eGwKysjxh2uwxMDojI2w3u5mjeb9iX1X0FQRxPp7FS/7J3CcJEp0/C9gqPzn90tFs5ONuJi7UeV9
FLCeascOZeAOHc5ZZMtAfo7pjzF7rZbdahRRqR208bcsHMomyIBSZXnkBmncxpWhGNy7uldZZ7Dt
dshaIlHuMgrY8X9vSRSOGh7rXWv9bBf8Ged/+l9eA2vL4WZhrWJdeBcm5oErMiWfrkFSUnLJhCzK
Yo7uOX0OjvNg1qYtbzrXFJJuzeYqy5oZSUqbc/hdmAae4GacczvxgxpkjzRst7ZMuXRfkphHjB/t
J5hGBhpQ0mfLkks8LwTRbAQtLbrG4TPthpygxTwmz0pS0lyzfnAR2XpZYkMdp9wpUXbsqnE/E23P
W9cqvUlRSL/+JxWWeCe2Hdi6hr/uOYpTkRDyS5tYlBZmxNERTE5WSDnQ0g7Kh2eF4VPgVYmOkBHG
M0g8fhCtJGD/e/6X4nPruMW9iv0jlWegcPyQwB7W8yTjLeqklMy8NkvRRXFSCmsyg7E7oCIcdKEk
L+wUj89wSzdBsTG6W115fLgwbbUGJ1hwRoxmXOaZ4KcS31uiG00CwnAzuZnjQRig7C/V70uuJyeh
e14YMSHrE9+VtONtXUcc+f8kFB6OqBksJGhwmaq0hJDK2V0I1vpGEZR+FiviJqiZbp/sOB8FsFId
yAJA9GZ+U2Ww5v/6Q/IvBUS5yEarPk0gacyvDUO64ujTa6XOhdNyKh30Z8RJAwxh76Xm+Tf73Ccy
2sr8qyB+SwnHryDE0niBQdb//KxGkD6MVO7wK5TFQWC6Q0iBwgOjvoIzAdFjnhoj+of50Jvgj83l
w11paPl100L9SjD5Nd2mG+1hr8rHi2wZNmhCRZ8JwPqwhYDJ2HKMU6U5eX9GfmS7yPvpMXl+n/VH
mR90HLIuAeQHl9ThMQbxkI/ZWhqtBH0A6HIDfQp7zIdxUCs7ThLVpPHIfgqgt6TSYtVMskLbFCkc
NumQcvlbhCoEf/1FTq0JHUFQfqQg41gdxyvOYDgGIyGV//2o0rIX4UWKAqYLw9ICeU/TFO12Eij1
RUHaSpBo+odShcF8A1oubE+h8B5Z5v9TlJzdVfUAVGTuKMo0NuaNFLPkmSRiNaUDmIZfaYdEC/rI
JQMKuUdx8se6VuemOp2l4hEp39j0WqiaF3tgk29DG4wdq3vAMTZAnI1sdulciLYflKAgEQpHEBKr
cv+Zih2uK8i0qJNQmTzZUgmcXbnn8HuJXNXWIDNfPL5JdpMzgU5ETFX0NQNK9yhLty6KMhJcZLBl
Di3gNNWLLRgOaQ3Zj2QWRv7MypDMnCzEhIKNLWH5EvrtiVKNwr5Xb1p2N4HUbAuJYQl7nMxYKsFZ
dzZod1leSItLJhfyC74LjYnRZIFyBeoPl08HgJo7JwliZYwv7EoZaCm+ibuIp7X93n0mkBDEw9ki
g63BQZofQTjCoDhREqpG2qBia0v0KdE1AY6kn8IqIro4daAw30wzCUvXmSblR8yiGlHyFidVNBK2
w/5EwdbQ75DCz0DHwyUj7YV+TlmimGsdEOhMc7P8NSQA+pLofhiRzzchfJt2eTChcc09Ef+XTj42
zXpG+cA7HawG8sFjoD/YvMwSWB4SjVnYbgBNNQBQfHyW2kgT/e0SZIBAhq8PzxVoeD6eQ/PXNUx0
axbFYB+tF85z8kqzg45P+xqMHFOYgfU0nL1RIDbKmkZFbjlteu7lqQDAwuNHi2q0Gbgrms1KskJJ
VhFaQ8dLxxrHWP/jb6RIAm0CfxRHBA7BUwwzxctq4UNuv83qACJJi4G9fZ858XQCWq29mUIuWO/U
h/cL2OwTeCy/iBRQyGCUC0pVKZjH7UpAJ8YjR5/dAl/aqFhLE/I4TJMC74suGRIZpcKSdM3HocJ7
fAcBIH8FI1TomCoGORzJ9K2w4KM+JfNet00OHKWXjZLIgX/smP69CZ3KWNP2vDHBo/hh91jHgwMZ
w5R4tQdFMUxBjjO5lX7goIEmbKgFN6WzHilvlvbNT7xwQMP+/nzO5MOa4SnbqkYdYpR+lOivlMj1
L0aKPaT94O6Xpsi3mk7mBOxGz70+iAlpRHVyQ09XtQkt7MtSaEbDEfjjTeYnIcRVWckZaDzLrZT/
fqoDchAotLdBoTqmUZCzqcdBsS7yE1fecqbYQ/LtBadfA9BlU1l3LMJFQbCO9j7Mq71AHNbgLXF4
aI3cvfQmwgH7dwdXC+Fcy09ObbwpVkY2DPFhslvxMFtPOVdu9wJOdoqFHMVzRiegqKzZzZT1rtiT
uLCP6lj4xRIaIRSzHv/xtJXr6ZBy52nBEA4W5CJEOgnMNC14P00fIJzdErsYJDUuH+ntq6oRdCC7
XBl0iyrp0OFnYVcMIKAhICtCJ1uQff7xhnqP0EcYwPkY0kCRxUSfu9+uYKDWiY8zIVp7qF+34ybq
dJ757eV4DQZbHzmMEpniDRNr6Bpf5oSbeN4Z/xJ81Or9eRuwkto5qwUw4rrwBYdwQVV66NBGLrzt
0TbH1gyBL77+RT87cTSFd5QrYqUzbW+sbwYywyg16sz1YI8p5b3o9Fa6UpNviY0WI5cpvMBsnnz3
ofqKgS7MiBOHxSwumNHiFx2LUCwJLjT27MVF9YuB9gIhS3/MPlN6FWbcSqKpSLkfspQwdUek9zzu
XHJfpYuODURkoZrSbzEZa4Da6bWQon2Kx/lg2t6YNlvom3J/eHBfkWIbS5nQZY8MKcJKdsLtKxb4
4jZ4Ly9wfjHwvjwVOyGguV/wba1Q6rqC3n/eLa3jlSZxCbAsqrSzZOK6x304zTx7jZp+Uqm17Wzb
GEobL+t9T1MEfJ+vPMhKR/T+QtMBtvK08bHVwLDuDkSeK8zLNfw9EHnHaFXyFN3f+puwmmkQ+yvw
12jbNFq2CDAYghAC6gMi1xbEFBnvQ6kBfPLTlGbxvydmlDH8CXMw/YuZEiVW8f3zR00twVkZx6SG
d9AXYi8TZlg3fVpdiNuojR424RDP0ei40XEP1dfJtTK+QIUE+zSCyLw/33UxdMT/d8cip5d7arJD
0LO2JLGejQ4jvfcLhPr1i2MBL1OiDq6BQLTr/ugpdzHwWbRrmVCb9KK+GexeTJhkGofIEk/A458m
0fLLhHk6HFUHbPURF+6y3Xaitw5N9jx2GQNpioetNv4HexzUWDrDlbJy/VIxOht0fgS7cSLcZ0TE
3S0VywQi8k+426VYh305Uneb2Bgy1PpCMtd/j5pNRIS0iMnqoqztpHsgnDLqP6pynwRYAGhp0BbO
6Oxmqo+u3rQ2ZL0Xm96NYwAZArPQJHyFJ+Z1HbKJC0pVykE74r20iLTpdMyIT4MipuJPTS2fHeWC
q4wMGOgKLRLuRKNlN+rtE9WNX+6AOym1Nvzp1qWEUzQwnuct0m/R6sb61NTVA7dVcF1opAftqrVL
eKKiRwUVg2qnZShoAYTvWinEOYFNLrSkVBk2QrxOCY5Byj9lmC+sTYpm8wjEArOnPvMNNmJsV7n9
FPKUsWUfqx5Se52wGHDmitP0qKMvIhILZzNu/ltWYjyTCJ/pGCv6iQmmQP5JVz/3fMAHihVL5U17
PMl996+jZKVT6fyLiAU5k2UQh4dNAoIHixE+wVByjIJM9Zn7Z1jx52HG10IpcDCsGyWOlJMfzRk3
B7DTDwL+ESQqrrcjig1bANq302pEpPKtSrd4nRbMEelCpv9ocdx/K7rVBYH4GzOTcUXMKlOF6mAt
gBUK1+6QUREyabBjwG5LMxEjQQxdRp7chNnrPQCDUOKZGAtDAuRBO3tAAUaFvYJ6b6HUFBwazQqB
UwuvFevKyYi/tqYJpcWvvbEI3uORVW5srC3TsaKlUQ02HYqS8FFhhW7C0nfzyc0ZY5Hh/nBu4eUQ
Rue7chwfZO26ooCR2fp72G4CNG5QUJxOHcjHPbboyYqNYAZzIwxY3wxhQD3uqIt164LHEZ6wuyHJ
8POfUTsbZ+tb/PGoyxgdq21kp8SsSIyta3lf2La1yEOkyfyzR2qZSBOt/Oc+obGihBUil70dj7Jw
Rl4pfSz1JM9FcltgJcJXHMq0lXAP1cx36Z6Zt0Wq8Xla2eAcggvoxfkX/e/Fw8WCqVH02br0T2T1
OkfepJzujj8r5QsmyciZvtm5gMCkxaQHgw5sBsoZUdpA4ivkMvYYvT7pZhUt9M6/LqGefb6FiJ3R
EeIj7FoNxmS6VobbbuWhZ1rg+t09w9qQRA1dJiNxy/F5pIkgZUj746AD63niE3i7IddmnLt2rOi2
SFDcQRj2GcVq+ILyvVX62sygkzvZl5lmsLoWhUNUhA3OJdbBZMielMpwUxrtREpmETOf6Fl6ssqI
J0rBu3nQVqPNhYLazcSkw9SanyKqWPCTz1f+w5/SC+m19hN2RJjiNtAJwNzza3N7b2nHOVifswKH
hqE4WT31cDVqlh6GL83A9f8sj1rZvU8bo9AO2uR/ZXqWcYMcftRC10wm0LUFEmr6uCia7l7VBLDn
XMoXHrZ7nhhzwVltvRHTfl1Eq0Zv8nPcxF+qnhLs/dDEPjHvrPth8UFKrHQ83NL8BQz+NeywInJO
VJKSJXj7ipO11tR5c3r0s5pEOc+PjYTlxKorFEq+eVqIOIrUg/veOQlkYyfo+cVJSCEAGwEfGQB7
KYcIKLo6WEEVlBPoigQTYdmKnMgkRUvZ1wSkcT1WTkIublYbH5eNVlS8JRRsiacCcp9C2YHsBpLM
rBz4pDMT6y6i4u62AE8fCQ1QYW3ECTtluLwhz9cbxcyA2FkkhXCVTCrGovZWRbytw5xmHW8K/YdQ
aaL662aWlO/DW8hOSlLpUiF6bo6ijqzaz4MowKx0jo6y63pYPqdUfr4U0XOl3nYb+FGnPZ8Sxibn
DZdvAmdhSt9CixQlZXsMOuEY/j1t/HHTT4fO3vtsIHGTmxegAJ1BO+CFZlIHcm1v2ofaZSN8d5zD
7raBuALGdIrGo4Aci4co8McvLA4bQwcPbMUWkYHgg+9kDEmKDSyxQgVuKjkyncMR6YA471LKrudw
s+cLmaYANrEQ/uNe4WBrpgzkzCdZzZ9ZV5SXS1x1UjdVpDfTTsjwijMpWpSAg3o4GjJu/wvoAd93
Pv1sOPl16i0BOGx6nXlmyLQto+2NiOdj+q+oszirHiJZEf5Ikv8GK9B5vEE+hRzU7Ae/Bn1dapnU
PTrnxqZrHZ1HSZrPo4mvallBaR7ccgemDr6MIgJRhiHRBu2NJ9xy2kOxBCntIhHw8cmmZ9fvqmKZ
5aPKt/+1DwjZxCRKkmrRaPYLeeek01Vg/N5T0sksDtPUPp1pZll+W5lFs7QpZuqeKc8iD6jFxtbz
1maoMGsAKgSkJgEQhyf3kbj4NOnILpriUj34dwK8jpfiOR4qdNgvYSc1OonIXu9GLaMIBO28GwJZ
vj9KxK0JA4O+pxELbsFfJQJKTun/uR94tGIfhFj2m5wzbW5GIbEZwsl5t5QWA0XxErrtebV9XWr3
JP8WxiO+uEyN1/St3bwzMRTb/kU1QPC1LZiXVqusUXmdqJMkSPIWz0FH4AvQADtUHy7cU0SfLyAr
vr2Ix9SahzuF3etkwqZQMviCtheHncrh8NHfFKsYzLA9xCt3sgNc0VChZlhXmwx9diYA0mGJk/Bm
/z6qOhCELEDMvcjeegTHxb2n8pVJBIuarPwbA0qEm9o4L0AE1R8RedrDuZBivr2II56qp+pOcY0v
Rdylt4fCu1+GqKLkhyDbE9jTaEZlG3CbO+fZfTYvsTUUnGZ/zg50biR0edL9K+qR/b0/fEQKtAPD
lmX1NAFfGLdwLD1FFR3fR+TVYomponnKsVUw1CwoXcqTmj2hoke4aV8H0pIyyhhOBCpSic0wEwnr
mXOu4v7t+c+90gUllv2b9nMWnl2U2msRkkNFnHkuW4kjl3L+XN7pXic0qNpsbSwLaT8z45mB2qKA
7V+mGh3l0oPCKqrK+12xF3ByTMQIt1bHO3UguF4lZXVsBv5MuwCGh6dA2j6WVoY98624sV2lDJHn
p8+P/Zu/FI7X9Gvm/3j/9R5NY6LCrcNR26Nm6VXcZuHLcZhdGkE6Hx6Sr9QvBhyQ4FwxiDH45qx2
yPGUDWDK4x0mNoG9hXIYXy2ipJAZ2Y7S//jcLb0Zi7skd11wUL3jPMyIYqmdbtE5lNsxnqN2FuVf
7wPibd9UwVxIYdTjTdbcEALz8Eo7DB4QvzlIk36lVJe8vE3lEgunCR7f4jtj2yhdPW4cyHXi3aS8
LJPokkEhOAKnqz1mgrgdLalXMmcfEPrqGetmlS9c6puulJRFpI90ztNvUJhvJfiZpOD6duGrqOMr
hhUKMmTZmbRH9OoxKfDInAxLi9swrjwZ2PSW0kvSHywO7nVoxeGxhZrF6bF01MZi9QgjTzcg1bX3
YK5iCoCAopGqL+cS880cAqRKlepPQdGfK8gXm2e7DrCld9gS8wd0ATOc5egdEwdel9cYwIwxDYe2
yJzdoSMrFB8tXBq7oBs9+KlazdYzxgA9HJubGHvqxYytMkhN7yrZZt3qWh67ydAN6DpaRLxk+L5i
M36UjCb6a2EdKozxxasGE4aHdupJU987DbuBCoDYPCIQafODpnRuY3g5YOFEq8fjSR5EzmP2grEu
iMlz7CQZSNIDu2kZRdWJvl1niasGQAEPx1Grxfn3xbdK6HmJqXMrf1xJY6wbV+oZi4gn2UNja2bI
syQJvkyVP1PCC92twQ0zslDWsHLMNWMbVJUvJ+nT7HAjlOg96znxq4xnbYRQ+MfGIqbQEy0jc8bN
sI9ZzwI71N+md0+IyEHWSlo8FDwa4W2UDg0eaxf9eSg6x/FBtYcp/5he6sly6EQ3Qk3NAmm0Sy3G
5PtYnOlF+GehhRGis1QqDw9ilMyS3Gpfo7wtu5CkNCGKZEP2mq+CQwSZsSlQlko//eT13HyQd+mB
/6u81bNJFVprbZlWNX1uSGb/JMb+epgIu1HB714QZfnd2US5bD9fv9TOZmcnFbFFeVzw9+D0IwZc
Frun5/Up8wD5xRpl5f0wZk2e7xfE5xOK8rGzo2DYFM8yoNYbiShRHyvh8J/R5s3TH8f74V/Net3F
KQrQ6O4mZEEax0pt7vJwMei/PZj0pvEaiZAkQ6CUrv0MGClni1Oy+PVtTvcPAaB6oZWQjg0eCckq
t1rc16z5cVvlkCjgquVTM74eSX54tvK7/ghlTHynCLqiXoetzmpGlKBkZMbE45t9Gs6STyCIQNaK
bRebdH9hZo7wLez8EtTQ2rW2A8uKnLaNX+HTBKad4PW5BaByMIrTx1VKDlt48hgjRsVzPoWzkQkq
hoCih3rrECzY21GbX66PllzxzBRIEmOCe01RBeui6y37PwiyeJIdppqdzTdw+lN9Z30y3hKQIu4A
QRohXt2tRJ7lotI64pomyGLwGomKp+pqgfRKmooCgo7qWuvvb62+o/4hqyJLyABIm3lOwyZxabNU
OHrP5uM2Wv6JEaUO6V8DMlinRhdYJKJY4ShgEZwlY3864KfZU+XS3FOPrW1yMnHfO0avmM2XW6em
YYOj3vs7mzkGPg0bI7X9iRDMJcZg+L/F5uvaGxxG0byHr0eUL7SvEujarQQceyPiQEpx4FyBPupd
lUMFY8aXWOqna4x6N7aq5cw88T+YjfhhlsRaTRUdQgax7DRfMtSGE3Bcs+QZ/XwPBiJovLfIevGa
wL4+2HkNhPPUhUJ+UBJScJm+d24Z+8Xk4PsDl3+3WBqp61qwkvxUni/F9a3NmsLO/uvQcZFuKYO4
DAzYIrVDZMDA6aq2lRj0Dpq8J7DjesXeMZiMh37zteq0GIUP0SGVjKVYkkuHnpvlILVSiG4aOp7K
4lF1Zc/eX9HJfz+106Is/R09l+SpKlXaavii9SW2XG3Nl3yrvxdeo6V/mdn2fe2DyfgDGUnGVAwf
6qDI5zNQxITOhwxBBPnYpyF7ph3wC9zeLLYWCOMhPaWS706TESwL/zX0q7URINbPd8I9tdTwUe4D
q4MMitIkvNDiW1tPg3W6hV3+WkEdjPr1Jj+vgLepEmgMKhfDeBtthvDOpYnXhxVdTNcTLrhYGWEp
3cLHwbUGTwO4lynv2fBtLTYcrxqaX/M0Z+8/wHLskyo2OOKYrVnztg9dQ2XmY6+FO34cMibmlZOX
9Q/sjMVEjbjVBq/2u+gZtXXsgHBpkr+w5UPMb2pxZnJmbDwoLBbNUQxc1rgW64KcKk6YurtuEDuX
wBkh79C+lGeKjhsi68j4fFYEhjj5XYkLJnN1YTvqaohI6PYgvmFf5csmTokzHCn41/t0WKBxOtCq
rN4vBODeoxqLTCZevTMXuaAqTdzt3utZfwT8KNFTL9T/kplq4U88r/9Y5s5mRPnx9aP08ul3rwd+
S748/uFgnP2hMOrt7FjLN9DeJ75T+dqlsZzwq5SN40dSp6zevkJWkmbf+XBUgO45mpoPQydGzNRY
L2Xfwz5ukoE5XSNQLXynZLz3E6i4hxpfY4fyusbocIIxh4nrS9DF8ggXnrJB3rCeKsgglWCu9kSp
GVmYQrkfcrJ4tu+n1gpwjG5E8pO1GFn1IiaRfhkCCZtK6+9SjMWjwcIDgkFD9UxX2P7XAZKkW5tJ
OrvTYjxYojf8aPG1nmb7mqe+KriASFJS1iMQRAhD3mX+Xs7FaJN38jH85vW61m3yIxBJc+KSJ/Wt
pWNfS0RND/40gkawD9oHFj6hx6Ugco+1CB+FYIqfGfeuu4purxGqlTrq4cKnuDEM+cQKPQ5HJK3W
PMDb7ifCeNOV7nLm9utBVFQ+s9nsAy+W6ZNpWV86kFztx0kIu2KjIJZ2LGq2UuPAyM04haFvhP9G
0gWpIsGOMjJMyOCXJPkR2m5wphLc7gW72rUBPnkWSaNZQOJI/vo01Ntc/On0vTY/yMp1Bwwf3XWv
IDkxxbrdB7yaI/jrGVE/kd4Mzm+MpIPVxL+lgx1df+Zy66Dnpynt9SBaVq4OvLaUg3hYD3wcbJ69
kH++bN0PwMvK1OHghTpfgkFyE3FFeoj+MDYX5IUBFH3jH84qk+Dm9aw6IXTlTEMYfvbstjVHuAg+
Cc8XqHfuGND12vD1jhvi0oljWekk8Oa2mWcjejov98jcs3DVslxcR3XEXqGEpEnsYuMBcWpjv7LM
cWnrlsWPa69W+tSsokzJ6v/hx/A44NXpaZoJF1XgJshiPNsxWBtwOPBwrz3WTlMqSIF3E9Xf9ptx
bSCYc4kvsVhByDpi1E443Ug/mcGeaoyRv+lg8lNf2eKbvcg3k8klP5ANsol75FAv2OtjqeWTQ8A+
Gb/0hrjKkPwcoMxjUPcUdkjn4swtP8+nOhtnsUa2ncJc9OX0lE8Mu6OH2AMs5z8CSnodT89bfMrP
0m++mC8BOOTXYHzcP8mIzFWZUt0Wxl/fC4Wk/EkCxx9JEjEQ67jE6Tle6svO8O6qQWkItOwmBXWq
2DhEo94+fxJlcrKsk6J4GQ/TyiJ/yrFoNh1Z6r2rTLlSt/SEuKf/ad4V7Z1sRACb/xKo4Q1yMtJr
aaLOqBbyuHCqlbCR1YvSBETFMmhTAiGQZbAuGdtjKGrSmSKhhvXnUZBpfEX/Er0eGDmuvK/ADPsE
6N71is5p+q97dFIbSyHHHrnhnjUmny68y00X01KLXhYES3v/wIW8OCMPFnFfnNzmKcltZVbQrRH4
oPHNlgcmq2B1xNM0v0BnE6k2HFQDn0JwroWIbCAweXEVIXKZJT/e1eSdWnAYC7C0DzHGoDqrEINE
gGFZUJC2KpzMNuB02f5453MzCgzNiERXtSsRljA8l4zpUTLa8WNX8mswjrk6ivqZlB9AXL9rcNNf
vHIe0FMc15cpP3xHOKjaDJag0Ix4TTVXrC2venRVb31/p74vOV9CQLy2cs6ge+JOc1KjfeKPjb6R
ozJj43ufiAqVOygkqL89Bfmk832NzIbmQfcZ5nK1B0k9yPIEgfgVN2apMQJ3ugwgfTEEXnVV7wyG
Pspl64JC4Uk3gJhdpceHfWtCALy77qCQVK6aG3/SJgt8cjs/5UmVN8YUyiiQNtvkKOxtZFRKE2hO
nbtI3gtZmF8xnEjGVe4Lt3Wu4j42DpKs0e05sq0FppMgyf5uw0sEyFDNz5qz6eJ2Qi4nkul/gBA3
VUKotFbeCZtQ5VlVH2otCDcxMy82jNVLYch024MEd11c2osmkyRUkGEYywaZVyb2yvk26P+vmX2z
F69taNxnTQm9MfRVmh/oIjs0rQFn4AlBMWVeBUFZhvMyvTimp6/RqZ9hXjDI/90Fzxgytck4cwKM
R39GsdkBXPvl4TQTX5R78zjn54TYwt4cIHXdo6TEeerCgbwSIGaH4HadxDW44yeAeNgMX/swHeEg
vkquGspxFCdOTDPX5EM9odZOQkpSmOiMxWPG5+mCnelqSOf5O3vIDUEwcVsTd6reX93+AaLvlCx3
IUMqfZdkakHprfG6+TbubBfns0ny8pSm7IZl30JO9Al3+5sYJNd+7m6pHISLBakdCoailQutgNLG
HijzkHm0ZlJoyeYGyM7XGMfXem0ig/wTIcyrt7NI6bcwn+JMtyo3tD+/LaTXjX+9jzB1KUq66fOw
toKhqQhAgmVTRDoLW/6CwMKwpLLe36PgP5+ZwUeH6OMvlVNywIY3XI/ambBmLESjrPQyTC9+A8XP
FLEYw14pD+Rtb2+shyT1cu5R2nN5N9+3mRxMizSz4pTrjIvRhB2QweGQXluvRlS/RYlJI1poaViA
0U2f3O8uWbvN4ldeGe/el0AzDnwzYtGevi5+2OHJVD/5UKmN9sM2vilsbadjG1zBPgUws88p6vgT
QrDb+E1QNYbKsJCaKVV1q3IOvpatG+GUrhcWtB+8lks5Gcb+KzxPhkoDqoQVRIZDQdl4DxDOGCef
1hp7RCcgWMOKupH5uPNEYan0Fr3g0T2HKV3sqO6fvwRcpYHiqSuCzXNRmikFdcHXNercmaFBroIJ
awdDIXV3uplMXQqQ9t3xb/XPxCZQlILozFHa8q70v3l4zZzf6UKukdPtqk9nDS7YvyQXo9cqv6Ee
hYZZdkykocms4Z4sAAIfgpoFsXgP2MBVzWn/B460igoZ4EZuqMYbYh52nO1TRCP59vwpSrGjLF9S
kFOXR3o8CXdvh5uMO0ccq/EFZvtUBo1Wsi8qKSpzxG88B16uq1k0I/jMK2Ri32skfRrxKkfVdNN2
XcGd+Qla0prV6LXodAzHly9Ot7wQKy8ucVbmPXvWhtozgV2Ww6sqCiS7qhCeBW5mIPCZtJcfZvTz
202MKDYzZx0wdBoFN9fb3FO3ORqnqr+DskupEYq3+nqTRG8ZatxwVbCP/TdK3fhGpHD1nwLG74NN
OiSOqQN70A38L0wyzSkh7Bf+FdQKPhDLRrL1BgTPSCE7k2Kzgi9XAtvNJ4mXKugf2ezuFshWIhQi
uRsk0qtt47hHpm5EdA8ZQ6qSxx5b95mbMyczAWUKuTxUMLhI920U8Cl8uoP1l77+DqyG3HJtVDMJ
bacpjh0R0o5ItF5SHRZZAr8Vqb8TrJ2Jm8csdb5zYBlfasVk+Or9qdWsxk6+rIdZ6hJuAfeiacyB
3sbow1nWUzLZthseMUd7L5QkZ4RahsIwZXQikgR79xqeQaQPjvo5SWDH6+jXtSk+uHD3QUZ7Rnks
nnHZ+Wpyn/f1Jt5tfIks44GNUWlyipoUCQt7iQ1G7EZQ1BD/iegMOyAnEf5likc1H8tS/86V3CVm
U8g8rQX3Of5seZx5sU+U+3EIWB3e4HmTThOfPWvtYMJP/kAeMLTVaP17DVMcqqFpUF1ejStvKk03
4N/ERfnZhCnUvFa2uJtH8Jo039kqxTCVInISbb+pPsykS9YZ0dTXPvaDDB79c5FomjdVHSufcL7L
CqoQvKkEDVTG4F4d7R4Y2bMuFC+xmQdbRQeHhXgxq3mh8cJ891qMifCz0/0Mt5c51kydD6V+WFca
JKHat25y2NCJW1rbq9z8Q0ZCtefrxc+1dx3f1/0jlm6OnKG9djNxBiO9ubjQcy8FTOnckEGHybwN
sxMkPL4j7uv+ZLlYvdq/GfrRjAwzCzwrCWTcZIMinL8DOiFrunoMAiYw/HD21x0X/jPs6zQHPwb0
MgFc87MAJGrtoyutm15ObBz9LKaz0D/1ZOMQyGVzchGmJl9BUR5QGY8r7TKZc8rGHgnToSWasZuH
Ya5hzQIuQAqvkq7g8EXcKnlKtpjOKoVSwR9g58cDygNYXrMhKEmIGythPASA0Mtg1jRScEc78PN+
oLwNqBfGj403lh2RgdBOkUZBs/vvD6OjmU209XH2epvOMqzDp2v/0H+vNUkl9hv6tAB6x0rubSjJ
DlC3NYHAZAOh9JQqBtteYygMuM4VtqWfZG9jWET6pnkWvfeZRe9DwWEkmA/a/UD5Z9mfI9uJnNdq
Vnv3Ni3sQT8mTme4WKMZ01d7fG6kyimW9CMT6HXTc7gt5DufpT7kvetvDfGZKSk3Ndqoq4ugzzcz
9wK1rXion6RREI3okMwd/jd+Jz9RSIEKf2Pki4pclew4WIPzIzT5VJ2UpuAMjlNVYsRhcPhl8YQu
/nrOF3qnFVovP0Ta2yY8oWJ3O0IQVI6/DraWoNCT1rYhXL3I/kS+TI6i2/Z8lxVLNoQnrS2S59Qf
vEcntq+ONB2y/E5H6pxZMkEFN9MJd7QKuEYyBFgMn7dhbildipmrdtQHMSGFB8AQKJdqIKNo53pk
ubzJvcAZ2Faw94ed945nI+iZ2Q7EuAv0RjMcafbSr590sGzUPOIqvT785H0UzUfxvaiU0gBL1wbx
QhbHFBB9sgM86EF5I3Ge9CrzmBJoKP/MKOqA4wbxncpTA7bXJSnU/XZoo1vdGxMEak7eSHvdB3Jr
fb8oyFPasp+V+hlKVO0N8usXI67cqGg236c9TsmpAyMUBREgHP6zk8P0KKfisUlDRcmr7U0/EpuM
vf/Wsb4LOmQvk+RriMvA5BD2PDl9IwZt/CC7zvR9ZSWtqR8XjolCAh56yCJATtL5ZbFrHp8DvY4u
aGmTV7Yr70QHuNth9hYJJ3SkiFcLzfqPCtxP2YgFIuoeXjmpnyreukmgLKJoSTpOswOO7JNyhrQv
HCGo4VzXV7cypr+QPlnpYQGNXQpsj5r0uzIhAMXJJ1EG9FDTJZRi2UaM6Lq6UHq7IF5VG5rkCZ5D
BbAE00vH52j4SlFCQnPUbtLtJTPQ6MxlXMJUDDQR44F5Mc88fkMpmiQPo93YJbiNXB5mjF2F4JAQ
JGBHayE4CSupCLdLy85mlWNMcsulKyTav3feUEV9qrKwK5phzbJPYx5+hQuy7ShzEcCISG89AW+f
uzl8ltvwXg8p91yVj93kEfGx1nxZMxx749uLARCiIJhUK+8dXBzTOkwgpJ4w3K2u2m7C+yGhHkou
5AAVoTwbdly/y2X8n+OhdiEBG4UrE3HQs0OEcBVohXsCQU/yUFNu8iMwcTdmWS8xWU7Q6aSBAzdu
lykz5/n5u2pLAaRcNiQRoACW0YC9lj1ooug9TRk1gVJG67jFY2HHrdbNe2PDO7yUI2cL3gqUIdUI
Oihvg9ZVkzJXVLTbZl9SKaos+/uSoOGY4bc6WRygJcsk4dud252gK/m1i4dn5LmyartGK6JmgWF1
DGA42u7QA9rbQNbnXnvHq9HK03dRFYXfGqSC5L0IcBL0kSZpbF58xd+vICUyx87oXIsyTOK95LnM
pVDaZ6Josj92VcuC45HHD43q9cnCR63IxaStDKENnniEYaOd3cSAYn2HAILYSGfwaDzJNOr8VKz7
o4r26G7WTBRXrqDKzy1ZfKUNyfhxGTo0qOTM66Rws8JWBEF3zItpeega/tqz0OqDcrtgwkKIZTve
yeRTt8UAf+woPpdVX4lhphjHJ9fsf18gkG0pTSZOb47rDtJ2Zi5IZzeKSS9vVjf0fQR55zmbzEOh
b9js+JM6+X0I7r0Kpg+v+i3l0+l3sLGses0n4hN1zydkq1324jAYehSXlCbaePHRI3iqsK1QIMSu
M9hTmxNYnHnEdMKRSdg9Rej1ZH2GlS0HwAvzCQqC3kg6dHr8+mOpvRoxM82+sICNeHBlv35sXxRd
Q+aiofv2xc49oYi9T+KUyMMUnmBwItrcqvw4tSaKs3bOlfRNQ9e5zzM45uTdgAVVGVyF3qcG/I0O
Bnphb2erv0R9oRc7NlgPiFwIzKE/z0LFhR+U9nOFu6mSEknsZv+e8oPqeMvGOmx7yPzCpHaJ851J
Cr0zFX0sK32NE+3Dwt10Z/24zV7vRPT15O2TT1LT3Prj/oEuX0adUITbMK7sLvawqiI3tWbl9gGY
qI/yo8Io8Tk2y6JGT8uCkC7qxFjzPgLGCnXecdRiMFdiZLOsut5z599AYJj+t9vM1mTNFCjzolAs
x8PZq2gw6dpqWdooSYEo/gWM3+v1pOOFlcRF4OUpsBt4IGzFF+JOTFmp8UG46W0myYKjjItRZyvd
Y5FjteP1ngoKEhaIQyeDfPoqyL5BI7tuUyCyifcAcGJOtpNdjn5PvFTwj38gwyr49KtmElrCTqsq
NmCTY+fGhK457WX/aXFQnAodeCUGMW0nJ3kuCwpj6SnQ74dg6ikwe7re4iudZwO319tzoXPLkIcQ
5NjKFtHRCugYwuVaRAUFqE1okL0CEzHpXXh/7ted2Nt5iWOEvdSr1502/c0KfEq50B7bN/bnpepf
l8f6L08gXqEPegfcyuw3qufrPyTHJ1L7EUF9CUF8GHCF9Y41K98dAa/a22JQVB1JWGycPujpIVEr
j8Bv1cIkBLbVZswViQN/SqohjkcYWwE2SUi3nohg4gDDVkPa8/e4VTMfF2kS6VFN0HVgMHwMPOw7
Q1sBfmFPZ17Vk0VlQ50P98RVcQGWn2MaNsQY2kB+b59MBHToXwWg7CQQWm+YWh1w/UYSN9QZH5EG
Gu7fHbIXue03ohtgPjC2jkxh491BfrJmREFjKBwl6LY8V7tCKnovou7Z+0DOfedFAWLbZjMFHLaJ
m+K2aKUMsvFWTh4Z/ARsfW7eFAuhjOq2p+xrIgjAXGM9MnLTSX3JQojClyQ/sl3b/ka2OklNs5mC
P6ieqTG1QDkfDlkjWAOyKljrE3V0SiBw0KbPH0abcrNFW5L3rwLGSyjMVMnSWOobi/QLveLEesI3
kbGCakqz2du6hT4W0ZqWQcWWZkKQS8bxReRaNMpppiwm83UEGxu+7L+hb9unnxsVLE+yOh/mqyS4
tsKkvt9Y6qp01zL3jiuQbvrehwmdg1rCyiU+KRRjBV++W+YeVcgsUKPeVDC8TEHitWC2eApF/soY
n9J9C3uG9Jo7yuKqVbLneCQPINyqTY6yNgKHDpTi6P4OItAK5iD7mTX3xrd+awdK/lm806yOxHu0
PKxQiC9k8kuH3oUK3ybowvHNsl0Lrn/GU9RoHgD945PGrMphLL8D7FEDBTUJeaOw4SN/99AGAWRY
jDIWhEHq3JdJ4tC8hjeiImlo6OyHmkI6EJV2w5AQm/VF4XfnqL89hndyR5Cl4570HYOen+mMlzqz
ZjOUz8J52nR558P8GH9dJhgSRca1AY5cDXCufW7r63kSR6sajtBSB4T57CudvU/qwDQrexc6IIBs
w7nV95ZDxHpZTvqyzK0jxG08V3y92+0exUsoyRhKrYFcMNvmL8qq14wcvEkzN0Jbnko2WIecH+j9
KgLWpcih7/hGcwGo0HlpGf+5Fbyhl8jeXbYFognTrvm0No6aoJ4juaER8fNQqpZr5heCZCwUif60
JN529nhM+CImg5g3W0sexspJ6OBWBd6VcggUUsS6w5jqCPlmQMV2ryivysTpRoFrR/40302rRMCG
UxXEFpZu7Pot+XDAnd0LKBJQRUfc8u8/LPb0Pvtt3GV97joVU41akY2igBicBPsnkMyOnS0kP0uV
dQ2TIpXZxh/zAAK9S+aApiIxywSZCMbbu6McneecvwIgvnxlYJZDyPngYXM+Dubhm4CEhAn+wyKD
PsdzC1rGGgiTWXUv8uvjy0MXOAYGaEUI9AYqs2hKszo5prd+IXgBqjajkOeMk4CwY+VMTtkrAArb
MxLV9pbZRz5FFN6w6eQJrXIpPyZEdUvG1TkE8DKswMewWXidRlvs50UTZQSAmnMftrDRxiHUGCmH
s7vQzHyhAo5l1aXF2s4RfdC56V4JKym4p0zDGUyYwH/YCpP/HOGbEjXMTIRjqY5p5v7LlfMTuBcQ
tfAadBVdma2NbSrYFhCz8zudUBcgT53H1DvZbE4Gxa9wud449dNDh5oM1pyOTujF1ggfoHMk82OO
+SwDhEdH4SAx0JG1aq8NjUlgESeAeu2K+HAJN9LWhFuwEEaAQyyEGMJXf3VwFzUeU3BCndNkZu/1
MgbHXkkk7ZrhzTBV4zZ2iyFWr1108aKWJ9HCFmtPGbPgDvf89AFh0V6J8lBxgQ4hiJMSU7GOPYSO
sy7B7Zwxv6S10qBuR/Onmod8hgSrA91HUgfKn0l6dONy75yViRw0zp7/zLFIoPF6PjWIr/6Z6ZJc
x3qWE2bblmsF3eHTq19nuSzFul5AzWN6chUnftELMNdH4mFi5qjxesTfV1WqzPEAzOhGpgvvSs+B
r7GXSzALkkRAfWE313wnSTRHIX9gAaTcJHh9x7VtRoLZ+0t1gvAJp2QOdaMg7yCYoASyAM3Z6Llo
iz5PQIRrkPPczDmUuXTSVJCXjBLhIGreNOboIPnk6VPnd31fPsE7d9QLpYsT83mA0cWJIFaVwGPQ
rkcosixUiJ2xnJ6CpR1cYkCm5DflgL/rE6dG5PCdTxN32o6LHotmAA/YPl1Qqb5vzk2cA4r2Z4KU
OZDVDO9IIYatQbIojbDTB9fZBUuIFVWQ5l2CHoFggLQiYIv3+v1XnhpEAexNjuPvYkT9TZEXJz1F
khVu1BB19oB0lkGuOpnU2k+wUlOuZ9Eo9KOEiJicyX91fIU8FOJwsT4vj2qq8UUeV66vKsMPHyGx
Z4QLPXtpcPEzBGhNY2I5W0vMsNsXIU3zrhGh7ryeOoRowBeC771YG6q8xD1YnjahXK+6IXGxEr82
3HadrTYv0eVOIo9W6fiS9EziPIzvHsoe1ohlGK7vKnXOitsqCHNs1atFRQ+y15MFuDXlBOSahuK7
tEH45n7iPY3wWOmp8sEPzKuEia+k4R2uisXxrpC0lKcCmu1TgqX6x7KmQI4cfO2zuhZTZIl+lfFK
JcyP529z4b8l7gctqUf8XLJra8Esr5c8p9xgTzYgQsdxVPeSRvsXNLHFNJCE4SgtQFumVIEnv+LV
lTUf6dqTkat4v83VcNt876kxybARryfxTeMaE20gkR/Ii1gN7I0OWGcEMnK2JOwBxgEFabFn8m3k
Wsv9gnLF3PCN4jCx8h3OjHjVR8f+x3Zh9yz7CMb6I3LlqNLHq0igvS0e+xx8aEKRbnVQmpPbZASB
z55Lol1GG0nM2J8ekzNGVrEcQRL2Ix1hle6TavrBp3MUSjqW4N/UDFYWbtCAbx8/LynwER6Sql4p
HNjuUvuom2vgKmG2CbQcCZFJTlcTSiecX0wq6vyjqdR8JGX/uShxjl2Qzz9cx4sz8nD0KrRfuCNS
YXPDbTBq2DPcMxb18fF/Tb3/9VoPdXi85NDe4nlz9E4AWM8hByEvxQti6CWA5j3fpBNhf0tXsJ8o
0xRXbrQ5RZHI9Ncma2Vz/G4FLErVhiK65MeWbQhwRN199bKdLFIvuo1jiXY9LaDiudlijUenwO0k
s57oFuxLv62u3w52AqwIYHFXpaeFpeKvSQJrsETTFPrXpf79SEEmVB3l5XXI2s2KLpT9MRoynyix
v8XE2fiy/H+sSsNhu3SH+zEzELenoQ4otNT1w5whm6TpzyIT355w3VLl6JDCqeTjr0LaSFB93VhF
XLx4fZ3VpQrnco2zqSsUBBud2wSzf5VTZUQqHEQjeHZpvdPBCl312kZN/tTWxEqZIY0NFAyTog9o
ctPStj/Bc0OFrAq3SVmMLOWQx9ovw2ih+fjpm1epmJNxYH1kx0mHHR474nLL/dKm6Asc30KvHOD4
Y21tlh43RtdBJNL+9VdC0+scS4pjbNPWN1DTyWoiN2FvNCq/MoQtGMTUqIPb33D4jYtmUsVV4fCP
xeBOVKvpfx5CMAqb1ALd3gndBoQ2kt7HP8EzdINvqrTZ3FL4JgQFod6cdoywD7vvVgJHQW+Et7aS
Vhh6BY45njeEv7my0k1IJ8GGl8s+frdaHykwhvghiFOX2fnfMSiGM1pGGeO/X9udegRj5ppwEdaF
a88RA5A2+rUZJGy90pB/k/fp1OfEtg3HpghQOrTNG+9H8YXjC0I37JtlVJbVLlXfSGqEakbFi2ql
eEsgC/F7JnYkVPhDu+ExveU55tmMxCnHGmNsdOkSNpa0A4aBOaQKfMeM453H4aDERbVvZ40mmIDs
8PDWS0fWdokrWHZRsjpy5DJOuXuq/WHfwQKAzfi2jghwwb78FudhkZv3Y0pxXPBVbHPH/qI45d+X
MHThvN/Tri19YGCUAH3qMD68wTY0y6Fyw/tMteMpPqESYgRPpCegDPhyHTNJquVY8wBlh35YoQ+M
Jkr4+qmIBlljGolkIG5LMjCIsJOjRVv6OkHA8rF+4NRfiqo/Rs9ko6xdXRlHGv4lYa+Pi3kQyTs+
yNX1Sqh0u0lFscKGwq3603+VCYS3+XSwhJlWGVEKGGtEbhuGktRgvL+FjOnbiZyt1ocQDikhsDJG
aMz+zKudFvJmTH1vOFNRy+ZtEPaDswYCZ7Zn5iVedNkyTcVl9Recxd8FAZmSI5J2J1UytXSvh8gZ
qAAG+rRep/YNtMcU10PbkFya3YGJAtzHD1ZXlofB0Bc9rq6ao/9A9LR6x0NjnAtMElFlGxo1j7AS
0SoigpLzMMxPgZD+R+i4698PSoYoEGYlNlzbriKr2PRYy120Ym6WWa34e8UKIlqee5C3bONOWqjX
Gf5isSCPcV0xPBR8vRWLNxehJj0q3KiK8v2NCtwvh9hwUqlkaztjPEAgE16QF+cQ5ux2JCmI3x8O
x7nukRy9XhnG1v1lCVZOqnqg6j7v1ksvj+EhgV/sVW7GLQY4V6fCkefgxC7Mvo07tP8ebPklfMUj
aySKpSCXbkWbWc3Dswbcsq9yATknDigXrO2iS7LDGVskYEGmBWYAW5Ez9/tllNMKvEsqg35GSPO8
r4fFqzD26e32OBo74GresRMeWpxscq37+wj3tOTZ/I32+0EAFJv6zwtiGWXF2wF8GfGqWcxBH09c
XF0VRQ/CwNNGUYA5ydr2prFQ1QqMA62AzWMX0nlcqzU70RFNhUhD4kbmoJnV+DnHEg0J935f1L0F
wZYCcaCWP14OdrSH+8ajLSZ3cno16l7egItnQgF31HnJHg6u6vQeia4tiGKa/uvTOtBTW5j2nAdN
rgSsBRdNUgQfGhrtFOzTVsA0IrWjG/Af0IhtrxTdBRxv9hoMfttCKnFWpv3o5kNSKuOvmYEN8drh
m+ooOhacB7DXSgINWxKJjVuko/2g3aUo1vEhFovpRQ/r2XVHiK0CelVnLdDyhfXiCUJ0QQbL2H3E
YQhnRPV+ni+LMD+hHC4mODwBW8GCXZ/zxSTkZKzUZWIsyLPcTZoPTTOr2qczNfIHiwrr88ytFx5W
uymEz4ZPgP/g5lV3RLZaZkT309EZpVUqPcjHneU1vnA4BVvHMOITyvH0XBLiVH7XHDOy5CiumsKF
g5+9J2E0d3a9SRBT9zKWRJjI9KbOuEN6lWTUPIGSXP8IfBRHHVC9Eeqh0RrdNuGHTOtEtufmZPMe
eDsr1cBn+/zzAK8XbPPMku7e7OoYKsfcvx7E6NBt2eFJPGjWAJjlkAgIKkxo0QidD3njvsnC7X2O
RkJtnPBuzkZsU5OM3ev1lHJ+gxSfBQWn/mwsXStihTCFBdPLeut9bT3gLFWwLpiFebiO7bbPShcb
qjpvTz3A8G+DHvRMRlGZnwVrev8GnTc9aWJ68ZqVvHW4G8VYLEb9wODenNmuF1JfKZT3nq4lJgWV
9YXv5E8F7yBCD92NpiiwmEb7pK6XSy33rQ1SOvK5naX0sf6MEssYv3BniTy6G3S0STcIJwG+x7lh
HrZNkULxJcddFtYGGbMYITBimKz+ZcdQHpc/uQlsfcQvwc44+t8itF8GDZo+dvIVsP2QpDrMlQuG
CTeTWpcOnmcQNCplzNI9UUui90w8g448vvjk4OmPFuaaxmXc6j+2j9GzmPAOLpROvpHG1m+/uxgz
T9nJ00CWEsCAo8a1WRFS0vTofrLAPRlWzolyfgEH1rzhJsgwnxdRPuh/sfn8HsSL9K/DoH4u9mim
bU2iKwXVMoDDTr4VP76nOeO9CvmFoIGdr/I5C2y+j2JKKSD0po0EKe1tGvnGwty3Z4B+lcyOWBIG
r9t7fIabpNlm2js+rvLMajo5qgY7cOAlFpqwcYNu8OagNNyxbJOABCXtlV6MFAlLzYCqTNRQIDLz
t0iYs8kETRdkWF/v6uwwCGk9zD2gp+PqAjJ/Hp5OZIBSUrHWYBUmydALyNo+XjbIZv7VLJhQnWAR
tDtMxW7jPpsOmHQ0txXOeGC+uDCLE/357t/osFZdXjYhJ8l+cc9K+kP2Hhj0OofRpgaE34hNNx06
ULeRfpJSNI2wmf5aPoojqsHWIhMgAA7j2oT33RW14y7pChbni3vmMw4XrNi2fL6rjoHTNsAybBk3
4MMKXUK+PbmsIm1SwVKSQS92FGDOUD+/54MjVKdFtQ08XbgZquyJFaXL7AIpkLBLm9M50ls3xzXL
gMfZcnou4xFyTz7YtK6JNGL+/ehLi5PdJjjTxDSzqQUV9gPw7bHkxtSrcAvCyFilEyr7nMEWnrQp
frnHTQCuVWS/7YzxfHDVc2zf5belMABylAlnJSnch5sNKXMxbXxKVog9YjI+oQ1OUd/EwbHqo27t
Ohm/8QXF6EjQ8w4nj+0fsk7lf8xNntKOXZ+83Xf33eu/fqaTYFtvzjI4bCG5JZ8IxiP3OOY04bnk
PsJNvXK9Kb5dYfJz1ngJ0nK8bOSOzL9nevsF0R2cQr0I58lbl2pjntHYnYrLQkqFlqnbpdJVSLI/
sTsMmPyjJ86kD8nEEZDoAlHOCRKmInoQj3BcaONMeixvqBpeIKtrzt6l3tvWVkz+7RXpSG6ZgYnV
LhpB2678g24aBeYVmXnk7wAtADO3yFzNlYva1a6Qz1750ZeNk88StYOhgmtcGI6IPbTC5Spw+ycU
LE+2zDuPSsIKo/NjG13QtyR+28GBZ6f4UmySNtnEJy/Ab8Bnj+42JR2pxUs/Rln4gl1WZx36GjGu
cQ5ImWgVviJkVm78BpnkbjeT3fU50ho9p8sgR3dEUzZOJ7uZq2BxV3elp7WJalSpnue54Loc/3f0
1cpgbYw+dYL3dUBDVh23C7u0knJs/rWNTGmJJQ1jpqO+3hRX0008Id05RVdlI8r+3Spf6FQLXKv3
0NOYeiYL3GNBE57zUBzvYiWGgeYcYoXXVK/tj7Z0Y/zwlE7XGUr4dLYKaU2k1trwf/3HawqgQNKO
lN5Snw1zVprHPwifYGxsy0jZT3DkLnL4PacwBc6HLK43D0fG1xoXGj4kLDDSxia69uxG7ixeZZEc
2Bg+esVOhAtBAaaBxiFKxnuDo8jfWCTnBoZkfEJt2n4hm585JAC44/acPt3GW6ZarYSroMsaa7Ty
IANc8YYdnbHnXVW5zX6cI03EOexynELRue0gqEfwtB32ZA3tEknw5TqyL8RGNBGpKxxeqOFgkQn2
dCiv3G6mpm/8Hf/VLf68E+z3nYlDbJOrgXxoAmYvZiYRgz5L8XRao7NlsDxHkHnw9kT93ZK40sQz
CFhXNI7GwGun81wXpA0k/1m5x6zpa2t2Pm6IesYovKtMQiawrfmgsxyH8AdR7heWsYHl4r7Xbx5h
vtYkiG8VVocfB35qtcwiRmpuhLpvruqyhn6BIlKlwaR2I9nNRufoNFCZ6iDOcqqxLD5vZkuhwZvh
UOAzSdubji0Szo+w5de3WYrmsijCafWHZvvzd4IZoA06WUf5rnnnQQX6fJKGxSkH5cQZhgsrtn7A
pGciHp+95aZG5xW9my9FCwUc1hNCFQKMtFVbsHFMvz1hEJwWOMK64lKItZ7f57BGL9OpTdW3auBA
esKTAlmswBFUkIUKGtMWPmC0TTtaw+bh3tO12XsjENVUn2p633Z114JYtjg2rHedKpP6nIsBPh9w
Tw3+L8SUJ88ka0a0Irc3DMN30ocZr1zWtN9FQBNiDLNZCAIGLG3KBNjaIj0dCGiC9vctbrPC8UOh
O49kZKWbvQCB7NT29ZpuY9ZgjFC6gBEfJN77sPOxButtVFiPopJcluDDGH9XbOXxGmOghr79mcF4
wBEglxkHbaTwpQOnIfL/Btt5EDcaN9Y22PlRHwnbSSnTxcdWfv9Xy87LK7cvq+DG8DhnV/cT/tCq
jTLyQenVxX165Y7K+SrdieCISjZNJ9aXtw4s4uQSL6G3ihqwvWWPSNCy2rBLzvQu7H9e8YKjhCST
Sj2PYPrgWxd13EOtp9Nyywtn+M6wNrjnweu7q9ozd75d2+pSAJSo4OUC5NHrSiuS2YfP8yZuW/WO
3g2upwhNgv4BbjvHHw2CyMzUSHL3n8Lfn8FnSffXPkUkAGxik8NHT4wewRiPLElRm4t469n7/CEf
+JO5+0aihKYXbI8IPjfCd1coCm0xAggCbZnLbYNntBGZrPcDiDNvxyMc9LThgmZLYfHfPbqQUSh/
YdXt6yZ29Xg5ammCH4sJRjMyiP98QnDHam4/WnK1MZjalnDfLKCVNFQWGS+NydWRQac3H3Mlz4/0
T9zMgjLOvPOTQ6gg6xuRRVHVmEPZDOhnpzihSjRlwc4tq3uydxgm3Tizy/xr7mvb1xkQlbqmLcm0
4qHvLEJ8rBvf8ScURuphgfdyiztnqeAPEOpdW4UbuAXIcNy7UrR2dmqln3bmTseIrrNF1vXJHwhJ
T6/k6qKLKlBcQYrE6WRBygQ6abdqc9Xo+EkAfXM8yg4fykt/Te2P8G9Tx5nQWFFSJXuB8lvcKJvo
ZhuuQvEevMkD3VKxC+SgqakuPsaKq5yABkt5NpU678A0onAm8zcErZdzhxbkf6tXHNOLLj8Dxl4p
ujeMEZ5W14VM83fIQciZKOCjOTTzOYCTvesHYFvXd8zyJmYELx4Qcm89YNgD1SYxLF2RdRcLZVpE
zC/WoE5V+KA1yCZpqHkq8kiD5noQ6wG2zf0HdIVqgioN/x7Gez3WPqhMlhJl/8977vKyRDMh6JSH
SP9C/z63MkO0Un+w304jNb47+9sR0FNOcUPRr3ibR7L7B7P+FDbmgtRBA0pARSUW3dxLC+tjb2l3
VVeMOdfPPARRuXLRvBGz1Iu5HcX49oSWWvL5il7wXpBJasM8Gg8oZVVh5qcnEtAMhuldAlvW8245
JxmnMoLjmvmTQ1GZTQ+H/1IVq/vuoqQaTqhgCwprC+djCEPraPaQybCv8KBDJ/pHxejNk1Q/zv3V
5P0ONdf5rOodJOkpo2zpg2/UrIV4NESdxK0KCUyh5FJEBI5LkUPcvjZJhvy3V+qEKXI1FddovKyl
asAJxodpMdKSpobDbTctWQj2Yy2UNYdByAeyEdHmBLG1KoCjviO62BZ/VL/gbitwx7VrvvMYNziT
ZDdA+Cxtz/tbRYub7SInZZUqyaWs4Bp8P9F/NmMBtpcFhjW8g5IExa1q/hQyIFwGibYm0L80ZovN
TqrwzWASD9ZOl6b80+oeR0nmKclly+6s+3TItGr2YFrlTkDAM090Fi9UFJyJ93Q/+4NKiUifOeVP
MfA+b3SWV2ynzqanZ59Sf0pBMZ+zpRvEvp4ym4FLE0wvKKDyQWArLdntU6hWyNN2DlcKUR3Hbzih
W/obr/inw+LuowrfstsjXPeAU0WPRpSaIou+N8LjhrQTeYd/y03wOdM1fj221k7nAPcNcmIxdA/e
efbTMvEeJFxAfMchzs3Qk/aJfgq9CKj51vmha+iteStG+6Mbz94OGWLwkteRJx9f728DEmtSjM3l
EyzLeLwYeA7MYNI4gHzRNRnpKGsoYvVI9Ql+AVQjiGUXv2xTJaqj2aJjenvn2FZNj88MpKjG8lOE
H3dBg/wua+lOgNHZFMEeCB2a+Nx7y2E8LkFLMlO9R5hBMJHpI5z7NW3QjO512ED4dQ7dJ1Eit7FX
q+PjmBwA0t0fu0SAxnQsOkZPh49lCdU1lduyHvt1wI9oOJ6rkdEKyJevjH0unG/DQtQmY+0GXWQI
hmuzTZ40BRzV0bGR5m4dXIzSYKp07n5RXeKnsRus4hHBfWEjAJAw6N/09XQExWeG5sEIyZQD4Naz
z3viiHHGLIClHyUacrB8EYUiLeEQ6MhW7Fkbyub5jZKqco19XRDf/ghdSSMaVmTsfUJb9ZOygUko
youYEQOzmdm9OgFkmgh7onRRIDsMOEnkvyv5ai+DWmxwGWgjklFnxkycTTWEk3rtTCvXZfeY56/6
eDwKjgf8fUx3gJdfV1LZ0kKEasULqY8RjYz4fmBqLM2YrqNmxwWblqRgOM/0Zfh263TT80B+/Exd
kc6VGKLqjzS6mZ0crgQZOH7zDD6eaHDZMlORWOQUprdh81zqAiaj5/xP4PfQ3404REY21nxn4vPk
N7dV4RV8T07VnFTR0JzR27XbVnns/TqrjOdDMcLS+QvJXXh62Ok171d28SYYKd08RrrfdF3qJUP8
8SAQEL+sstT1cDoATsx94CbbIGKeSg4qTPun0z6vjCoT7s7Bk9OmTyL8c1Tth/hz+xuPo4lwk6LL
IGuKcJ+SdnGCu0vpKLMdiUXaLJxzmF1GFa39gy0W1558iKk/6Q89LLNZWwofgDhw+SunUGPhWXCi
w0i4dGbsnocXUcYoDnBM/63DSCEm9bDDXe+IDxvoavSsau4/GCBlC5Z2hAPNLzDq8lZt1s+n2Gxp
w0syPt6XSg6kUwef5MkwsC7Go3ZHsCsDeLFAGSpfOyl7L2GaK5k8x0yvY9rOor/pvsLjt/iAToBf
Ee9pJcbXxC24nc0qAWt5h5naNf3uGUE+g+zv40kyvm27R2p4MCvH4+TJJqk/pUNCuG8VlGKDy1BV
kUiEeoCDnbCNUY8w1ov/9Z2iknQ46FdyPwxzth/bc0R3eGdKivlMl+VDtQ3h04p/au/N21VM7WHX
J+BiKY36SkPfGTTSY+Uy9EWegUaDpPN0HCk9IPd/QOY0ZRxEpLQMWF1vsDmJWOB1YvG/+tIXHYbF
V2fkKE5XOP1Qayo5viNYLBNDrqxq22fvzKgYYjp7LgaNI9swmJ9k8m90aYuQ51jyNjMSrFqESn12
qasMT1XyLiHUCgLtWP0i/5QAVNOu7Xyk4znxsS/uvJb7Ma7KR+xa2HlPIxXMSXJKGlk4yK3EExIn
lOLxCloXvUFp5casI9LnfgzMkP4NDNurK5i3WyFwwrKZYDRRqaA8tX4QaKLw6aV8ILIjlW6JQ+NP
yFdjQqKoLfmpSG4N+iG9zZaVlO/dcy+Pn09O4D+SoiOAFIWxS96kB1jgPxXPiF4zHxgJduZE0DFF
JJJ7zAtIm4kIHOYbAAO2FrkOpsjM0LzdRI2E3WSZFe1OGGIX5LhnyzQjLhIkQblQbx30qJZEMT8i
5ELIAIoirzR/guH2r9JgrC3JwJGQS7BXk/Ha89bpCMHc1xiDAxYXziPwLVM9lZnSxfLiu/J7VgQv
AOyAuzzr7FNj1t/TlYY58tYjRbV+YAQ+ghcLO1rmzmVIx+lPoMDKIRpTxCqJ7oaEYnpB+cbY5e39
iQWR70ChxU2V03Pe/b3mPl2WBY/kAPci0Q4CSbTMxpHJHH/PXNswM5kB0vIdt5vmE4E6kTL2mgIg
5UU/cvHbDRyf1Jnpre4b8dKntUDbTAQGeEQL+mu/6nZsyzXvgt3AzG9cRNhPZVbJjsiusPtRgCDV
53jJoB8iAQULvujXAx6g9pthOPkHdV41U8W9SM6XAb5JysakezYIPoxSv/uejVrrJLaN7MgT/ZTA
4rg71qFtXyZg5Ulm4T2+IhtbE5h0ACiNJ3PWDDpmA5JKUDrvtR+eRUgE4/2LG7kMhPMwVYTZ+uAd
hzWZbZb0T33EzM5tAo5MP8tV8FQabqC2nkNUkA19wKNyvil2RJm6tqffGl0oxKeIlv0mSnfl/kOw
7O8YLju2vCOCmqxe036ic2BGDxgU6EJ9YKn1aHPdpX+2297umT6w8J2/TPLA4CFHnsIDPSOMSphA
ninkF7nLZFQ/qDHNWl41FAHDQdELMJa8KkRR7qvju3bmwRAWPY3/mahX/w+RQNZW1WZB1CAMbohH
D5PNUBnoVniyOEOUIqA/JR7ElSR3GyEmZXmZauugzGhtDil8K2BD5VH1jFVb+Fkv0RDtlVvxZC8U
F+zsDNgQuxLYEdMTbVUmbbe6V+MnsieCUj4p2WSJ5nG/IvD1bKbCIML22FY25CfuJgXCbMx/z/v7
CRUzlazFmddMCIOtunefVDeTULx1EFNYbqBTgHm2bs9RUKNxLoAhb4NxB/e1UALtQ71jr57p2Va6
D7Ju1wO6XraiWlSJ912R+NuEP1wLDzadORzfFXtn23JWcPiGW/I9GothQhcnviPWKD9IV4rOqA2p
hlSr/wOVDvkyDjma/bGG7FVqiOs5zN14J04PSKXed7hj/KB9iuYIsBR09ATT7F15gVx4aQ/3l8MJ
RzojYjlkaFc4MdCE+znijbfAuCkEoyX0NBujwx8woWVYvW7Jv3eVkjvSnqagJXY2n9ybk2K2o1xM
59Zc6bnGkHM1yHbsfZC3FsaxU6hsL6YGYaGkgpaVvOTGjru/gbxKohDzytTojksB/PpgoMPpwF59
BxDLX71gsGr8QNYzrjLg6ovAmEy/KUbSQAI4Lig3+YEl2C4uPx7AyrFRuFuust+F4FfnCr+C+xBa
fHtEN3J8vj4YbsoGu/9E3Wjkd5X+IXW1NUB1+5RLlzwtWTj2ZWakb+az1GyOverkIyXz+2+RJuFH
25bOvxaV+RxwuBHLcDag4RLVlJh9f54+O3V80LZy0LdGdd7LRuWerbZye7QGAL3A+nrKW9ALBH+V
1XGo2l1agntt42FTDZ1SwFYBE6XY5X3m0YlgKDYiDhGwtdvmTTyNTppLQEQaM5ot2iANTOFZBO07
ifr837P6c3+fzRnhpKEH4DwK/1/Bs6ADt7nu43fmRfOw/pAFX+S6pTNyuvQ1fiBtBZ4YMK/z+2fI
DEOze0BIVAmwD0qb9wjh5vNvg922VYKsvbohAZntW/qUtiUbQeXLexpyj/b4/0ia5nyTxNoDpq/M
pi3cXZqrtsQ7c7W+CqWSPqUtIPCyc8c868gPjD3RygNCCMqOfumS2iiwMGKI/xYyzFfjzCfx4abL
JXAjbVM1qU1dMf9SNaOTa8Hj7ouZrq+iUy1LaIDU4OLUNfqdG/0SozlWwTMbGRnqHtdgp0b0L8T0
rGuxSAlvh4l3FhpmM/APN1M2/QcUijQauw3p+zJM6HLoe7B3iWLYdvLwFoTiPGRYP7V040Cq1t7/
oPE61j8F4o8JzcHyxIHxj8PyNTbhEAhdEupWQauszEZac5BDUTJlXu7IdcOOPCg+ar5U/NaZJDa0
JAlNHsl7OG1iRnw0cq9C9wXLWQ6JLzNLX/ar5KUv0/tCJYYXWZvD8k1KjekFG0XNzEliKHa0f2Is
3BuPI6tywB/80GbNw1Eu8RzmAUPsbNzh7oc2xgFfA8Wde+tGr11icqwqvbWdOCoqXotl4fumUSUS
PYXkULQx3S47rUaxRxrEBLJvcLGxwd188dA+kSviQVxRoMKbJdLrSSoX5wsZK37rtfqQZ1Ptr0R0
Z7fQ+Jlll/6p9zF089TADj2hB+bc6mkYqvHru9jQn6QwdANIkwO5Ool+KeGVpBOCJS382Up/YGQj
/UPC9ChB7ioioamDDUgO7x3A2QUbH+BJXNtgvtio3B+vfYyUmilSAEXPpnHvPAvBRFTNpUw8dbbC
/ZW3S+5PUziddy5gPj4IFs5Posp6KZKxh8nkpWJyW6+9xqJgMabVdn+CF4uIJod2HD2pobJwSSIV
fupwPljSp1G+XbB50g843DzeH0I7T7RZwkB1jHmwK+MDMTSl/xKL0xAFLmQQBkqwllSVHaH40phb
rHPjzXiJZEtluHDYPbfAkbd1Dbrx1AiveDexk23TOHRZCCxZmB1vi+FXvHgd+UYI7Xd26PzgGaSu
rFeXNNrhNFAom/45/cNHtAS6FnDp4mIw4JK5jXUaaCRKZTAi1MJpz/IKTZ0FywvTMP8XGXzQ/0vE
N9G2X0jluBq+chEwllRZXfS1i/a+7X9+13z+HZocAiboF3KXDpv7aC2AtZS/hOoik0aQ7tEs1p24
nFFHwe8i/S17p4ydxRjfQsIKaJvhD3XYIxNUDQKKJYoC7u2G+/ivzSCRh5+9pHyv1gfKJy3/bYLe
Vs0/4ijyoP0n7IGENT4JrWbTBDXXQtEFMV/Tf/T+ilcI4MsVAWwQhWh1A8DKHL9hsdJBfwvhQhQM
n7ncmtKZKuWQs7uiCfZbAen8MLXx3dl/rjJWm9jMVARd4/t3uqwjK3b/vq37oBT8fG31xKKcCssK
RWnNDa4Zz8Mus0UB+AmbYPVqYxrkJCZfCdEr81LQZryAeGRGEtiu0SDoryRiXz26tgAG3fxpNJ16
E1dwF5hh9DxE3QEs1R1VdgwKUb/kTDMVfeDYbB0BmzsITrS4OWH84uiFonnmcid5Aa1Vf+WCiuaY
3Ne3wJPg6O0oRqeg/LgBReJ5OHjebmBKIcrRykTqLNQ0MNQzCmOVBmCCZi491FuPnYTV8j6gFUeV
rGzaoVcwc2yrUlxNrKgcC+pXP775sPtxqeNqLn3nvDKPtXpoYPMpF73oU5YxzyGlDcqjrZyTvwAc
oqyu9vL/+E/+mTzkd6+NXXRstX6ewFiVEeVqxy95rg4cX8RIg+nnBuE6aT3O+9wXTy89GB0iAnLo
FxlTLdmF8k1zhewSa78+41wXAjtap3dqpyxSXs3cTffZJBWTnvpz8uIjBwfDzOZ8saHBvrKyY+HA
9O+S9CGLreG2d69G0Q91Lxae+Fa6l8UzndSu+JrVOmFNmP2X5MlxJGKi7Zdc92OIYIdH4/a0GjOE
5jgUWNwbEk7EiFpzjBMCaLiw9MzumSAxo75bNh7yaphC8+wGRqMxzD9viwRGZAiQnOTdYVLq040+
QOcwwayQSlpw0LhiumJfrALlh12CEBYer6WWsiu1tizmK7ALoiKgMiYBfGtx/etNJja0tVbifhBt
jF97sqZY8lnmYfLfGuX5DOJdTqij5nIHkDOIQl2SALHuwriIiKibXHsBcld7DL+VrBZ7eWuTmD2w
Ts4wXhJip00UIECr+jTJl3Y/3iQ9RJXLCy+RrKZqG/pWFqnOLnLHY++UD9wtd3mTTWs72XZS31oM
4PSS18n3JWcUW+C38ciw9VDHkwEM1jpx48ESylD3M2C3qrVOWWMLuw1L2TfNt9hbL4w8dELnEflH
O+B5SbKcv8vq5rRUiY2ywvu7fU+gnbNEEodYJ21mkojQVqJePPNde4NDNxTenG5GKCqzkvkc65Bm
LGo+2iAgs8A9/GqMzb9rIuNDFAFNjoJ2nQHphTjeQs0UIc3UvPFLWM3394jEy30YrDMmp7Gc8ovi
XnpmN5usBhWe0Uu8pQJp8D9gjSizr0uc4UKkGL9A5gVrejIpQLTUqjAR9dKNi4Ra3WDMwfDdclOu
muffJ6APt1n1YUMqsxFliM99cjPiY5hGMq97ZvwoEUKLG1w4C9nvP3bgKwMb0XNAA9ZWfYTIKsmv
+1HU3Nsj7HBm+JlyJcpnTSzeRVzPnW2uoguy+jeA5pOOUytHE2AXuWaier7XaJJZpXQJvEA6+4nA
Pi8Y/+gb1nmdsUYNqgZFlwh2eV7qkQsKz8w3KHcUVee3B34qvp+jehGAXYw8P92w75eDkC1PS3Wc
rm/0fZUVDiH+XNv4POBagqCoduoQx6yD1mB8d61xefRGz4QvXBTW/4LgtYQ7Q2DbbwmPkxlzFNqB
HJcSZAcO8nr4c8wSV4baHD0WVdehOAlStnyOWr0y1gzb4Q7+UDLD5v5UIpIp0sBJ9hhvZGzgR7sY
s41I9mDLY1g4jt8ztIR6aISrrHwMdUEYFW9ldyJSVho2rMpOYjcXiGlHFfVBDS0deehPEn5LDAgW
pRU+hF0tR8G6ViFj9mn5ZUwD4EXehym8DNuLc8CeGU8hBC3bY6UfN5MmHt54OJXlCk8ujGKpDEui
8Z3rWJLR79Q65VOxh8nat78uXdEZOkMYWPcQ3VgTlQunBZso1seyDi/4IkCkEmu5dq7ros+uJsB/
tdtnuosk31/v/AjmZFBRtyAqxLq+llCZ+SxhCsnRtVWmgbpqGiSQk+8ftDn/4leHEZmyo3aGd2ys
Tc2f0lDfxKfbjjXEO02dgpvbBYaOQm5DcNIwAaMDXQZzggY7Hb20a8SoReSzYdp3yn+9kjoAi+uv
IoMTYB9WnF5MaTSFyo1aETkCYitDGzc0AbXg05iMKBFqlDOoZbYKeDUCcNE3GJwv1YzqxYYmtXGA
3osut9eaYo4URLMIT3lzTnNKZQfTjeIP+xNPZOkTTlHZwNTRM9ZSrgNNCzA73lqQqiJuCHGG5iUg
NNykkFWw1ZYQFQxMWbI8qo8hF9xCUGqTEE0pNyG8/thVR7LIj69VnBn8h3SrHGFc9rU28c6tW4Hp
SH5rWUZg+hzKvGBtl2n8gFLXUqFQBlHXQ0s/lx82YipOZxJYUWgPedmgKQhkz01ib2322zbzdo9Z
EeCkYGyeJXO5AIWABzXP1ZNdLj/DXL2RUYfAgT4K1V8FNp/1JRokKhpMHvJvmxoLuacs9dtYKqB0
bfWq3cnL9yb7AB1NjuP7HYtp/WWqmqP/+X6FYH5Nhe1Eqk+hRHrOShvUs4X63hWtpq8OhJ3hLwxH
xVgRsJUdeKmB1V/KU96nGgB3RLUwDZPLZ7LqPWMtwq6XTT/O8VsrJwxWZ5yksBy1Kq2aYaCR4PKl
Hjv+0++LAgsvXdlpHbRKMODE6rGyZ9hzPwnoY7F5654tLgKeCZ7rfFDVUIdtX/c6WGxiuno5xcya
80a2tXrqv5VdSIBT1HucdxavdNxNjcI2ii03n9j2WPFrFz2o7qARlZ/b2dCTF5kc5WzpN2fMiozB
ZTpxph/9G1QF7hW47g7oHBfUYigT9jD72Zo//2f11eLTbtahMyvsHG37qD1osV2GD4dL+5KSDFvr
4dNbcNf6jL6KUhmL0I4BRVd0NZcEPSWbLyo4J3hNfcCXoEehwTRqoquUAkV1olvz8PGqiPpYwKNF
jOH0cI9LqR7E75LAEQEjpddn6mc9GKczWT8Ynk4LFuKopDM42OjCVSCBZU4jTZiKxJi1TFrdirzk
PQ5HIIj+jxqy1+s3c/YIJxkPmhnvIaWUSiPNHjaFGSsNn3Moy2M7qQv7ERkOCNEZTYJ80ghpyygG
Ub3US79e0B5nS/YrKo45OGV0D6LU7Z7XW1D7ohfFhxMqfZ6dtqh1e3p2FegjyEWP5fw4JFpKQOV1
5pEgHfL8v+EU+xmAA6wR7uNr3F8vJ/Z3A+Pw7gGM3lhUH2WbBUEEi70w3HMwRFXTJEPHkt0hjvE6
SSNZv36zjOqRvwzH1/YoD9dbM8hYccv/enwo5AQ14Eb0npb5PZ9/ZBqRz3v6uJvX8CLZzUTgE1Dk
of0F8wB2fqqYFpa8+j3bAVJSN/JE3AQ9dXM0ykR6P4TWijHavoX85COwrm2MdBJDujaS2Gjau9Kh
zr767eZYIA8uGAzba7x76t90xDoUIazG3Rk/0yi+SshnhkFP0A+koCkKeeVP8jafQdkI7qskbDEy
xPOS0xHlUbZrtwalXdH8Hvktl5xutjw9Ng+Kxvqb5bHqqZugeFQDTqIWBswk7Fm1g3hX5x3wlEmF
c28iOGHjDTG6gRp9XQiKueoHUNdRIMFG+03GwgJMtM+gwgNy9AuiwRNeXgmP24H5Uuo9GUhV7vjn
S7oM0Z7Ut4zqOps7kuZzwIp2iAf5UbCmqeZJDIa14we11WJ2JGAXNpDS9txwU05vscGTQb6rNVLB
DqsEj00u+Qw6oweSURcY3+vuM7XyMnazXLpqndsFcgGSeTpKLZ6G6eQhlHa0TxKjAQYALmP2o9QN
l9z9KRFzEwELm+xqhP+SGxjjF+UUVJfey2tSuCWr2gA9mzuuvk/wa38NYMmk9Q8ZF+uhUTBM6/ih
WX2Rnu4a3Wfu9z1aqjUo
`protect end_protected
