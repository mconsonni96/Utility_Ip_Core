`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
m5oq9Nxtopdx66GsZCbvV4JFco9KHkPcBtbUrZRnNakoP7vbsbT+EKhcdwxM5VaL9gG8EsWsTrtF
tNy/aeTA6mroyrZ6wLRrw2K9bLta88qZVjVcWY7JdA7ZFIZp+T0KJQV2ugAWr2/05nuO5n9oE7Ba
ea2lf6m34HnaVOztx9i/8o1e33bXFdgE5LEUmxnEvTNZe4/JFigRlkr5lbrTl9KGNLQ/aNulsps1
jvq80RcfG10Ic45EfkJxodPicuAZpKeu5GLbDr0c0ZBKxetKvs2tVk/0R36d/TmhtG2rwbacZMtn
c9Ky0VRpuWxGtjvJf38X9qugPYofMjUNVsljOw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="MBca5CU5mMy+6+50FmICimuLmbgF7pALxXV74ytYMww="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15888)
`protect data_block
GgIdXiOd5yvB09dWewOjDS91LPcc0rKyPY7/gmgw2djQjiKNmHkWsnVEb2CszqZvIEsw9/gt5BoD
+IvFOShxdUcmV5+lwZ/LyBMfc3HQvGJN6YyfaAB+dtypxiUMVHC/Ck9TvB2DvRPqc4Ee/gU0x/Cs
g6uKuxhZzHQKG1WyUPbaK8T0fgkRRndd7r3zt2NRoKA+FAhVG72rJ/KLcFsGdIxYcpeyeBhZzX+U
nN6l6i+zxYxyaXyS2hWxNzNHCP9kx6em663Z6SGWhUDFg7KJmmF65m7+AdPHZy+X7syG1QH9PsAY
buP78HPedGbhV5GAkOllbHaI4ydRTc/tKApvLOp3tsmFiU64Wi8Hm0PgYKofxUVUsQOn9IU2FjGg
8UoMSMNCx42CCqxzJVksBq/Tb6Wh+10nSL6SRuz8dHtNPlSQ7DIIRCW5ZWQ8OHaSWm04yi8FGnju
TX4njQUN9etk7tT3lU+VrG+B4wQEzKPkm5TBM7AkNipt/RMpBbsDoNJXjQomehiR+EGKEWELNu5q
ZSZ69ILJ27vGpbUWvMAlLy274pzVYuY/Agez0UfcAr4pKNAnhFjXw/Z3IujJbT600Cw0vIG9Bcn4
ahk8B5rCdeqjBaL+O2rSLuVv+EN/oVTglHV1dZP6bvH23R4AizX3fFzXXc9H7hbgPlccecp47RN7
sB7dJmTTIFXEZgVpR9eBgjcZF07+3u3Mu1PoUXUo7zA9GHfts1tfHvyJAZAnJOo3nPOdxP5L5su4
HI+umuARQvY0m9hOWFc/hUrrKPWU61aXt9u83/7zM0wT5Vo4fXYmp0q93YflYPzzYYVpV/Oew3jE
wMGct0IIBjXrMPTbTuOqvW22kND3ayrf4rIvTJ13FFvS6j7XqZbkeqXdFSb5HKZS8v85MwOWW/f0
iHgyTAoO5ZuIUend+RQIyYPiq/sBlgOIHqAcBKpphm17PJCB3dygdZViRgBxHR5AQ/zamx394Ogx
P/MmzOLqCyPHjfO8tdbeGGPSG4MT2DDz1QcEBM+GFxCcRhfO8T95I6tf6blF0MsnqnBN4vdCSQmc
5JkG0PQiuyVJJDWn9h2CF5gWbA7g02OjPhkcgdKs0snM/jsmNpvzH8yl0pxdUrJMu+NlmQyEPuFs
YnDZ30nqop+/rE88CUSeRuXAAVvOGZ1Dt1lZDKb2XlVGXAlj+7BUWmkqjaHOLJj+O++/bfUm9FC7
lUliitDBT17m10xuDNIrI7OyUvjOirPDPcWbZCa3zMWSP2Mmrvj+ifoQjioZpDrjbz0kP6MkxENK
CeIVzgIgKtLmqrYsbxYQX7G7Wl03f/CBTz/hAKMHUncMOm6vYZ8umfJ5O/WhYWjog6RzzPkfIlTC
gdXtDd4fu1G7HeJeg+0eu+nZw5G5kmOnCpCHsPzky75CXYwPkDzYXTeDAQot/9YAal1c+FjLEiWu
WNdxDNlii2I3ozYhOmE7Qw/bHXuza9iR5GRy/PdUpmHrqOBxKFxlfCFXLAucJv4rtWgH4z+5BZlG
Rcbkbqzvhu5zYQZZDjiatlEC82fIpWC1qzQ1LYWiySVCcWYZQdw8So8F1VOWtdttexEaCzd8omwq
I6sF6+qmp+qyV+lV0/EwvQ7beCRx7V5M214/EwiOzzziNxdvVHr1T/ivlDHVgRgOwaUqceab22L/
U1iU7u8vWCBgtCf4Ptm7hYGDWI16SRC0MmxdJmGlGpv1xJ6Wo/zqKSOnUOLgRfxoqj8PlApug5yL
dzJZekt6BR9Gfg2nLsg+GRmB0ZLVVTJC8SOzHhCQfB1HBBl1SGhN9eLgXc8P6UVcfqknJnVcm0pV
qceE/A/v8Le78eSp4GWS1urirjE1jAF7COJj06oODrlw3M8esoNVwVfhMG6zPamrBO8HSRja4zVQ
AxcOLWHvUaarS5HkBzudE/yvcZSuphN8ghHrFI0VobyFAYi7BluABLmZl7IhoAgcGNg2XTIDmEhk
fe7Lq2Po5LPOECufaykvEW5e9WFPJhzLmwqeXyCWTsk13WgFxckEgh1NO+jrAzGp75JPv97PPNHh
k5XMLaFCkOPeUMuuiuT7Tm/1ZsFoRajqJ3h50V3ZjPGw2p5GMw8NTkzZj1u14flTceuo/i6gc/NT
NzkVEGwUZ278f794dRVzr1fUsVyTOc6ShOV2bGoSCw+yUQnANRdh8TQq0RaF/Gsx5cmldGrtt3g1
hpkHOEbpqsvRNzSNkPo50kSfHMUzyiQ8uNLm5DvPHnoiFUMfHV0cGQPz2l2VDL6BXAq6arcDCbos
4WpBN5qBs+6qzR9VHPGJB2+v7VtS8llF0q/3+Bpav23hhziRUQlwUyLCDBc+2vW43wwtUqDi0lAD
iMssdRKBQCDLEEGWYD11G8jUqahXo6tdXwArbFHzjQUTHcWceAaaQZHVhruwvAzT2yEJ4VgbZf7J
UZZTwJEPRQefd4OR4LXnGsy6ON8LgH+allq6GXgcZDC3c053ZPLf3I8/m2T7/m2tQ76//VcZTW09
QoBoZLXnOEzAn6XS4jrWJ8kPcGTmu+5uS3F3Tw/Lul0Zq5s2TGGSSpr95AyGxN3nH/UzvCoCYckt
0VododbatIAOsoqXeyX25+WkALC3VdcHbjt/TTEsBlfG/FeKEEzJ499OEvRaEPGfmlK001aq5AKb
sk5u2eeJwlgpRJqVBeggT0faP8euEoB/j2NSsj0I4FF5vEWsMfieEJLCZLKVj686FVkc4pjSrD1B
VLkqwm76CsJj9HxBBLSZqXAEPgMYDBv5S8sUZ6mqa9ECHUjHQOecoHgOsvMGUjj3pcn3zYVKT2nQ
tJv8/5ri6LXTTNowiOuVrRX3sVcm79E3QiqU1ZhzyQACCkbA3RzVKW1kkJBKrPXkjdsuWceS1Z0y
mlVo2csV/sAj9NTEU8fa/otsHqfJuBGyn9jc3AjuNs6uc4I/J8UBg3dCOvNg3MmEqgyjMNOWjdY3
ooMh5azzxehEsstIJ5jf/DrtDKZn5CWdIEEat1HuPuuJCebYsDJbbeMycG1nO+WmRuQU8EAbmDlI
/tPc5PCmdG6Ywqf4+sMAT2CwembViWII3wRzY+YkmlQVn+tdVZZxWwnCs9ynLsotin4lWqnt+CdP
QDA0dNegl0/VOSCCzjZHSqZ2N8ZjIDgqSGrYapmdhXlqh2RIySKinP8pK4kkIQzXaglC8qkdKaEC
cSykEJJrdIYC4mQ51wC3gr3eRR6/Iz86tgcWmYaHUaLGG0CYZz+tq8MiIWfL9yzJzmR9MeDX8NXZ
PVV6oYAI9yLI/N0CGEGSArtw8tFNXRP2Gx+KME0gYuRfj7FWljoDO+rZ+Xkzma6xi+ZV8mXBiZZc
BJfViagM/OYIGtQCAHY9IIZFc9LmCLqEM1DEuBbrKFcnJsNgV99abTSFi9jZfrLIPyFzjGGtcEyF
F5nwUBB+GljH4fWZBptek7mM2mCi5sijl7N6fHWbZDZNzvb/O6qqvRMN6dLFpMzMxMyuCE9Nmt0J
yTvDXcA23ZoAH5zalUWET9vrGiCnsOG/hjmwF22Uo2Iu7CPa1vwzClPswmSnU+jKUwQQPZBho5Do
u1egngt+/5ivuahjGP3unSOmdOFAOHutiq8Kp7qv/DEqD18Esy6rjfSsgavVqQDrbf0Q6R9acFAK
HutIrKP0hWYd9t+HJnQOrMiMszi+xU77qVoy6qcOWtk+wjbM/dVoAPo50Y/hyrqj8hVtBPwlDVoH
wD9qfMGKHEl7rDsnBhDci3uFy7deE8sZfG6wLB6TaeM6CPNr38abRw5/m3swIkVCV44CHZJ8Pq3S
47lTgSJNhNWk4uFax+K/t5mfLrm7h+QTHkRhLY/UPrKlk4WedoMNTp/NpBbdOCjd+04wWz6Cjmte
hCWEa4gXlDCbrhCmLOINk2GE0aA/5h9+gsC68iYWaYHkumLzVKh0cGClDNmVNnQO2nlNrtKfE+M6
j6YGtBykrOfD7m9P4cXIr2tmvFtDeHquDFVq7O6q110fqGurUwO1d6SLL0YOCpaBthIoS/4l1mFL
DfY7wzDVIOYe2Zcp2AJMSw1DXC0lv3GLiZqC1pHzxj2w9w5Bwgu2oCp9ym1y6iKciMFVNMfbEJpr
Crrvl81fiw6BgS4sq5mBQcSUMR7roIUv3Xq6PC5UcBM8Lg04/UBKHUldwdoa4G9RhjbYHQk2VRuJ
i2tpFkkdKQY6TltQsDWQKYt2isbGDJJLRe8cEMOImkpljYNvtZGATdJ+O2F50kLX2o9kf6sfXZ1n
uqvPuSqa1WD5aVal/UkFOw+cgZlUba1H8MdWUZl9cHVOz74SMvdOx4gGXO7FnXRrnkftlN3Qo1d/
I6Gcl1em2h+6vepQx742KAWS2S3HE1hri4uIPBJrbL08iFsibbMaDym3IV7lnQRlHP31qciQL/Gg
NTPBSn1EpuhFRA4rKUU6P1f0rZ2quOb+GIDzcYAIA6wp48V87a5tixLKAwH/hLIzegGO+Mr8P8fa
Zc7NLZp9chISCntbHsVbOEiWVja4LpauDGeiaV8UmtuwQ39qSMA3Ug8hu2vshV7XJw12R9ZEFAzS
sdIrgesi7vEF2Ete81KZcbe1yDofSwDoyL3HsRbEu+UoUU7cOxiVTtRNY5y7/HyQjlmkgOMEyyWP
PisHBKnXWRCAaTpa6VndpZ8Nyu8ORuGI3/Dg7N88qaKyBBaoVRfq4imm0FV8hGeXR4rt0tcBV/IB
MGkVGkaOWKtR5ANxoOAPI9EOQAIjhWb5jRjeF69im8uz/BgMcVC4UmbxsC/EqVjKkvZwhYaVcTI4
Va7VpsZrRN3xR8ocx799CrwoVOHqTbpkPrp+AKV0MGCe+4vwvOC6dBZDK12ia3M1+bNtPzFeOvyy
Gs9dT2Sg3DnhFTBW6hVhW41r5yicVexQfE8U60Zsn30mpMrIV2tRTTHtG2eBfEzrwMaYGXEg/2aO
QlRtN6MDLwJssSNbRV1yntHNvFpJMX4Q/ythTWcj9MI3pZiV76Ys2cf5kvm7vQACdJMjSW2GDuoR
X2qDXMuFOJfPQLOwVoTsYLy3rzCAJImxeb+YHikAdvu6rh2FVS41sF/Vxz7V8E6dzhnSM1Vcmww5
3puIAOo4xccRrRtgEdRBHqSpyiyCW31OF8VdfXjuG8+vj6OXAAUbIEa8lDfyglL+NAO7OvfUNGLC
UN7jiOKtci3YORQ7/WJpu1PbtyyUwo3i9f3zdMTpDGnthRMuOBUIyLHjo322cieyDq2rCAgONQ4z
d0r9sIFh5PxvLfzH6OJHpSb4eCgHFJLyml9ZX6FQqvtz0o5Rw8bvNN7WgBH3k6JUzXYaiMO8WzvV
yEa/oBUTFNF0ue97nG1A5b3QwkfxIS4rvHwuDZ0u0ERn1kF847UD3RZ9bCF3bFyAmw1AVj4RElDT
rhuZNrhDa+dZf8NUvJwabJng9RgNVr6z0o+TyOzQPfimG0xsBBiXXxb8iboG+wUyQ2tVV2iWhaIQ
AymEssEF5BuGfxGXkGKxVc1AERGkBJJDo5ZJHloBNzvZxFRlvolXRBPbtwIB2XePdoBcJkc5TyPI
q0f5zWrrpIrz+jIIjXGK48A92+epTykhtjxJNROK+aGah5Tb9BlYsOeXW6oueuZYoQ8adJpK/94l
xHi6vFZfLk1DelaxGU3iljEsJjHvGs+jn3998K4ThRguKMJiS1MD1rBW+oGeEFDNVy4PIJHosuNY
l9SJ2HJMTdi87lLsAzkiKYMRn41Eztj8VwzpHM711/NKjNOUqRDxpHdI4rvQq34ZCnySsI1KOK7x
QKeTFyecZUz+liwVSC5X1jgy/LKhf/2jTNUetLwpbd9OA8nkq1eaAiCr5px71gDR1YZoR4N9cNhj
HrWlY6IDqacxGp3WDMRNAdxJcmixAArCuOwQMmFipbqeeTVireNTkoVeu9A5i+YrzZonq+ISx3OT
Ak8johb8m7eEV6QrxrvsNKapWGGrlgGbj4WypTGqR62IKc6BLNSIP4PGjzcK5I5VnHEJV6oGt2vE
wVrLhV2yEHJ7V/23w36j5AlwYFUFvyQRgc6aHxlnkjX1xHTorv28cDa8zUJlLcjyRIdfd9O97uoo
6XcUMb9MbIDPY/wj9iWFtuvE9ri8TU4jSicIny58MeTzkYSCWy6sweXDDezmKqMdRMDJHcNWSWUF
i4wZU3//3Zmb3gZ9GeYhVcGfsJkdZvhQYUHRP5bUJI129X9rQQclHylDDWeK2W01ib7kcZ6HO9Wl
S+DZ7kEOsBnyXQj65cQBk2o40+cE4cJGu3/qVsq+OllpGKiwMgcqboeA0G0KtOe5F3sbkxtkrDf/
td+fn3EorMRUGL6DWntAGWUsXgRaameUWlKMQCVZzTOllqtUU1YyALguoPbO6vHHwZSZGhZ/bQy/
GS73g/WpopyxNEFJ6IfFB+WhHVZmPVyvGh3YgjbH+qU7CQlnVbI8dOE5Cm1z0367jJ/BsnuZLcQo
7bANLX4lxBeIVcGmhYYCplt8AjxxGc7AwwKV93No5bdyNfNQ/9v9pDDF9vaT+zk4Qtb/6pmKcoKL
juEalz60Xezcgsx7J7AwXi+LQo6zt49YfQHzEi/1ge3jGz8H+8ED45R20GnCGsyVBXJWlD0wBwId
PpxcSZNKVSw7z0BSAgO1fa4wYPHz+QOZ5RzyHAG3HGBO0lh3ShoL2D8Hc9rDmjgr+s1bb93DH6sf
juG0v+09cnDxDeGwDELy3AhoPmJkr2vk8jOnicjKm/tG/f1BU3W2id4wWi9T4uZREGNbA7sOpfCA
m1F/s1pKqbG0NkNeHnBlIQk0GOI6Ke04KLxZWG3H2jxNm3hYbqQkj+MszCTNyjtx9GPFYwonVoD7
xtp08U3qY1Uxo+6naAXdSiC+sNX/X1mCoh9ZriYVTu0zULHNsngqPYDhAhJ2L6pS9fp7MdHrP3kA
VAjxPF/6TVhEirWKnEqv9bdI7siyPXvBwAFfcOKhZoiRaAe7s1fXMtPe4Vy+s/DhZTUZgtb3hbKT
YhJQ6c/YjQ+jQvsquZuTSvAltegaZDd2IEGizX899HcFUZzzWsjNe5Vr4VK+uuJrPzWYc1Rs1IUx
zKfnZSz2xV/pz583lZq4+QTVhtZszRXOziKXx5RrXGORwT1kJAzMZz9E9ayQkFr1Dw5GaP8jNDQK
Inpl+W2J7ikdyDeJzW6uFHmfijU5h29hD6IRraJMK02P9A0f81Azeo4YtU7fI3T0RJOr4disacqC
sW/QrSwCFXxzU7RG3pzf3RDjna2JnPUQwvBUqQpzEQbTridWSW9aYuxwqrVyGKYENXNEvJ8qQGK2
WPV1u10vr8yDXbBN+zvdjo+U0GLvDwEGB6g+EGZATe01r9wL9BIQ42XG5b4mfQ7wdP4i+Qk1u9g7
yl6p/a8ch5Qcx+Pq70spLDQaEEEDorXs0P3vdlKaglTJibYFWTR2nRv+HoGEmShqxIqgkqHUXFKd
Py/UyCxWerzGhmkKz7PToameI8ar6PxsMNNsRG/k87+IGJVPBdMVjP7oYvy6DoKPyFRfTjbf1InB
h35ZTaNWCi8bYHJ6E2UCLesJwYSkVUct6GxBxHCFAtC+S9Z7HZo6gOI04wITdCZHMYz2q5AY3lPK
UPafsWO06BSiqz0m60lQfOzeSvdIoVmNJXFcVwICUTf9SODqyg/79A7lUongHGRdHEgnp9VQ3Dou
iCtMRMHncd4aBemlGray2QRwUzLFDd8YL/xF6/Jze/dfjknnLM1D5XID4y9Y9tglrZDDav+4P54c
m/Jz4Goyk7Gg+ybFvd1+9F8twqewxwxa0JyRtNhVWzIiYbM4YMeT88imc5klgniPo2tNNb35mOtA
e8EEM7PHcdyTurHn3Oig43D34ZwKYOC76NqvT6AfbwqNCKaFnh4CzDeWOaB5n0+5/7S3XsTVBBvo
TQqt71lztr5zi3pmnt669zDZtDrwCblefqgrn+ogCbvi2C+/HsK7vUBjTpHR9KeTwo+m2z6gYUWa
SksI9NUZIyQu6t3fzNdiyLl9bktrYi+r1SzdsW1udKdqDWsnWSmnMFeFWs71JSi6h7FaNvZ8gLz4
MSkrFQSezNJ0J6VDtoYzLzEZnq2BncMov2SNPEzA+WTaUV4jHi1CKJVZ2YFmEi4QQfyZrOUuIIRk
cZw4/5Io0DzE0AsmOkSMTEJL/nEqTXfJMWe1bJVY136VFt+0GKbQJgftFvn1b0ete35fAFKjY6yx
jYfKhsBk6VxY7zOh/9t6x/ngybLyiohGUmmeM/EwKSm+nAGGPHB0qzddH1KRzYk2nwY3dMEC7u7w
SPzJObdnj323LgTPAmcv+yT0T1xzb7psGuXHhSnTiR7VyrzA1cDkoHwKosp0zcL4ViS+rt6pQFBN
Q5FSyOIKKTfhfaIaqzEr3znNA/wvvxhBNRPF7nrOeXKw5kOyCnzlkD6Bmw7zyTr0AMhfnaPIAYT4
Bzfdhh0ADcIIxXqJxsbtCvxVBr4fWdLzj9HQWfa2Egp36DL0hcJFiIYfiShk0T9VV3iMhTtIX+N8
QrANVU2FfOV4V/xevF6FIxWhLWO6G4kmx/l5k4dxufgcOjMhBrrCs2yYFttUDnmZx9iXyYlSB6+h
vRPL2HhgcX0Kui13nWKE1B7O748rO3SdsqRbeFcPRUIH8Hxz8KwI/zTnkbYtMi6A4oF8kIR9P7pi
q2kqz1dRx+M1pCCuonqizSmfp265MZtlI1puJgY6FgWoJ1gJUmMCYzsj6tOWGBKCuuYoGE0QYDij
MzjFk4D3RMsJnQc7Mz07QTD29cMr+HNOYtYVhR2v8UKurktdyVKKID2BWoaMGHa80n2JOX2copNv
WOjHroWW3l+6m1hSXbORgry2DmLF63oqbuAveb96IYeVeQsmCSI6blXexBQwj1BiBKZrIf4+XWMM
Wj85q2ne1XuK02BMTrQsLYp6gy78U9FwJdcSZ84lYXdZvwiZzcfnNUM82UPz4Bneg3ZEUDb8xXZ4
o+cD6Wfc1DpT90aYDMEaffkTMRVezV+U5zyFQNekhk7KwtXuKo9MN/401UObK/9kVFwfAVRzHnMp
/OGsPql1RnWhWRv76H6kmr1/LB9gwmoEuTAeM43hsTDKB3gcr3q3RufrOtfWF702zhLzFSfirqoZ
X8d3D/tfzg0BA3smQor1GB1wgSg1Bi7qzLPT5uIgRe97v9HcENNDreeyOK2xZOkpYoYsz4kC9omL
NArbb9h+w2oWzZHp4mgqejjdJ4qrAcHtDMq9ZFfue0t86M7ohcFVLFQBBRDr8qX/I2zA4rOeqow/
dtxq81EqEp70lTLaFTnwi//xwG9BArVJzr7Y72ODPON7TISjht9pNDkb4mfHdfSZ5wl3BVpDCEK3
pAzRAy18WAm8Q+LERMyjwl5Pooy3wGsfCcpHhM+zAs8D//jHM8brJvPSIQTcX7xqkwU4+aZe+V2b
ju/+VkuW9rT7a+f9mnq4ZpbQ0FY5wAtbbyfLaBpMk/RwEeKZfNbL7lyV4iRSDKxiefebvmNixILx
h2jkWmu1dRSLzjU2SSSJ9dgVhx4uHFJUItV07WomG8ZTDs3xbagrTAhRGb7r5oEcuRlfjjfDWfqP
wM8tbmMpzXeHLOQjey8mzfGvXjsyk9G99Yd7KPoM75P1PrKUF8A0lCgqdAcDFvnNUuX5mBBPsFWC
dxiNOo8U/KKc4HuAoRZdSRlz5i9wcoPAFG+sNogt1kF8hlp0TBjycWfY9MF8fz50d+27HMOed62H
u27Ai2KeLXgPKT29galw/DOzQgxv96Y0fHOIw9/z7EW5pPzfdVHcQ+NwOluA9UTDm1iCfkeHUUf7
oNmsobfLW24G2HCt4wWixTIDXv0XBgJfZGw47rqUzAA/MvqjhmfA/rsJivQMVHzthlPSuWfIE7tT
hgtSeXQMTBVycmNL5670SEk8eZV1My3zK1ohZvKFL4ubcCVyL4YERMjpsH2zLftay0OGZz4K99+0
LSpyrpqT9WJWHYMiE+zSWJw4nRXF8a0Bpdx0Apv4Ge5NvySN8CbpiQ7NyeOsouEH06n91DD3npJx
q87wl337rysye8h2ZArVF6E9vejilDfTsCyz/ca84VR9k2s2XqWWlD2pg8Kbt36+0jhJdLuUxfF+
xgeZ46oIiveZqJktJ/8IUwobDtG9/4nK8k6a6DYpIXh+hpAt5WN9cdBKFrdQLnkiOLUjJ7XqqIEd
Lrji7hBMxhCZiXEdUJiUY2Q0IWT5xB+HDH0N0UhzTPLB9yuRIK4/T/4by1ULR4YwkOZ401V6mrWP
xvZL/dGAHzvgi5fl/bG/qGWKh03jKbwjln01Ejs9JCgfx/hCFlXyIlkN0BP9Jj9LidCqmHRwlDob
rwTdBTK3OQWuKVD93eMAre8Jcimb4pqfpdBAQr0ceCk6xA4fBYvvo2cGQhXPQHYuma5cTiaXZxqw
5V5ZZkOOM4XpqIQ4yAJYvaTLxnXygw2H9Mye/aEjzPgwBI15hMSh/xEAbfOG+iOz2IbLyj4tu3ON
vKGAxFQcQlbFEhzUrr7bvKlQRqj0FfhD3cB0ee52FoeBpBnY+gcS75UtUT9+zlbONA8V89iqMM0/
JEJezAgj97jrRNVD7F8RQ7cPRManerLZZgtlHM4bGge6QBUyjLdRAY8nUhVhfL3f52MycV6wn9QX
q0x7cx0X8GijOnHGxF9W11kEZo3Q+uJO6PRTGGBUtPMLgyTRxdAF83aPNS0qooaMK/IrPfQZtLe6
6h3/FI5P15xtxB1Rq1844dR6tiWVgi4PPvMtI7/CLLJmE73bsyOWUOPWgzwzdp4H3A+bEvO+Vwj5
AlrjV+LA3yGM4Z8fRNMXTZQgPL+lUTJzycrCamjB4sO6eNZJFikRJ4RDjeFVMVCrbScK8/U7yG3p
6M+Ye8KpGVY6ualXRdokGipuHhE5/b/cOiK5oj80hfzNUHULwKyuU8YvGJa2qamNc3P3CNCN7Mv0
0nkqq/2ZfLW9LFI68cA1hQtnFv9mww3h/0WNViY6uXXyAEX+i5PE7NsB9uRPvUJLVHytYWU49Hfz
9mfXdBjTxH4FqOHfsIkAwoDof2MT8YGUjwqBcXSnrMVF9VJEXTTJ4v8lnk9DiK1yrgGZOBgW4wUR
ScH92K55yx3SwCD+qKkOdn5DtsiooNEUvOGz+e2QpXJvLig+Q9ejmao6AxBnBw9XItilRuVTkB/8
gd4p6xOTj3hTV8ViozxxIVguwt93+InkEhisQC72C29dNhyKH0KfracEN4iBg9jNUNt3ZcMTJ6Zo
MGFO50dBROfAAWtdm3LQt11gYwReGKqeRW/zu0wvPqdlw9bF7VAoXamvnfOYnA0XYYkiuuxluXdd
yWCdZ57AKUlL/uasrCjmPzXPPJh0FNX1llnF3/kRT4kEStxGhNaHwDfSu3iYXKN2tVS7qH633xLN
MMbwHdhgcEVV/YphFcc8ZELJIqHoSXDK/z95lX2AyzT2xIXqlgMitMgHbzYeGHAMppdjB/ts/lOW
LhsAlN59Z/ZXdZ0EqlTx3TK3SKmIDVtclz9cWca96ZA2mQh1LjLhoNpNYWJO+0UPXInwVjjWxSfe
GngXDD0djR7K7h8sW2q4+0h60WbrC/lkAGeimUuI/gPaYk8TlGSPnthJDIeNqQfE+4W6BRe5NtW7
yy9xXnQ7nPJa7FIoNn0FRoYWIeWtrxVsb+XmHWDcQx26bkgu66fsRc9C1qT8ox3o1jv0EmxCOXej
igz81Ubg6fH/AhoUe0yIAvxKCJEpPBV4XGNMZiAawf1nmIc6vuDo8iYrCqnq4TAQcIEGjEHNhQ3x
NiJlB9vv6aj4WTmXAWohR+CCs4+FAsuUg7iCCi6cPkl1PZRa9hxQZ4wNGW1L6idYPTVPkJe7octW
ELTYFYNy31vxjSKkuZ2n53ycpg/xAOLEZ3We/i/7z2cigNHQYpVv4Ue441cshKZ+ckKkTLHnLD9c
X2d2Al+zsPfNGvSm9svdWml4cqo8aYraPZctKHGQBjIjHg7UUfCffQeJtwsQQQdz+62seGhknv9H
ENdmjrGIrGGr07WN5qqCwwg07eFrndUwHOBfBlRqAaihJaahGct/hN+fYhzctz+CKQ6E7JEfn1Ic
dpuCNcgqqxVdNM6pDfI9jsjhnZ0cYnDUl+SPlhBokXKI3leb/WlNFWpoCrBsPAsQdI9/CzN3PupQ
xn/9d55VwUOHQtezsqk/3jJia/0X4KrDqtHFw4qQNsoUwU1cqUzhPSzc873XnoluvDnAoMrD7/TX
iKiOTWWfeYweqAh6f9kHJ8ox6Y+/N1ywDCvDvNnSM/j/wYS2818spoqu2alJw1P7c6HPTK8D2ynN
XRIKyh/NnJNqM1mnun6KlyFJ3mhv4eaF+H/vWB3SRyDCmfxCVCHvOoCSj4iz5j5hnChlfwPIAVGq
wFBmwkj/sbuG4W8czXRixzJMW9d9scNlUbxyVVInruXGNaJ2he6Llxv6IVowYnLJ83fGz/f11wzk
9vt93o0R7SAK9MxwFbZ65OHkVO/HYnKZK2k4HuAdM+OANGSyW/3tyhEA9YWIvLgu/USLQsrkf0y/
DSGWf5cH9rbk/YYFu3oyh8rsjFoNLpAPNavJDZArnH27Y170NfsNLyggul1lBhryVSjaY59B5At1
UgXkFSsQ6cANYWA5xRaD4DVmZYbIBqCCKw1Wv/e4f63MaX+STAC/I4Nys5C6RWzaMXu2Zp9CFZ9U
C9soZV9s+C8Gp5L55qGh5BkwCH4aQAW/cdWY2bX/AdFHTnm08ZBinHEy3E7bJauzuWniInv7YI6U
FrMNDjk5AioHMLQ0W1HhYyqKk1JuetKHhj7FYzttC2zf7YbBrgdDEhBJZ6/Xv99cV3pcGDAt9DfE
KCXfJGcETxAHI+VSNsJGydmcxqWk6dEwsDEZxpLhzdEiy6bMrwEL+19wnGrP/vvTnRoD/xITmk36
Y9YCt38ES1lx9sZZEAgYZQr6Rw9hFs6N4iT3mVwzYy9ZN+U6IR1SR6wRSs2mbEZldMF1HN4Lykss
A+PxNA9SEaN7NDW3Ish1hAuq2cz6hchNVU/eblT10Z1CXZHnnzWjCR0RiVe3nQ72qHicpLS31rtC
J7khzDz9GkT02ziDDgAah8wASjCav3HimvrbmIDuGKzvsQ6eE41p2IVDuXoADFU0WOqb0WuzHFVO
I63vJpW8OUObRg5j6jB3bgHNGnx2PvV/7R/o8yrPAhU2kGFeCsMTVxPAtlFJnSRx8/uuyW/2eipr
VO8XCs0crwlC7dZaK5he29BS6n7Bir5PIjjckD4ac/QtsBxyBFBgiKvEAF93uWemJuRel98MANN5
nJjcDUypZhoB9sLyKidgXSXm9EonhWEYGlJWguH3TVQV+K4PjrX9U1o5+k66TmFlAOesKms/qwP9
xaN3eNz23cSS36CkcxRMUJ3X2IZhVVSF9d1idnF8kXB6N0JxpmnyeqZhSmor5K7ZQ0L4KHOfG5gq
8QgOIoQ7XbNCnUPvDrDCZ5CPL/O2bNVNZ7Vn0UCVc3g5+W3O24Ms0Ba9800w4JTm+TX/PrYpkZun
pw0gEM2Pq7LzlczurI6swECKDBb/dmVdiRgjjz/au8eH2EBt+2HNPLmZF822+EVXvxYogMWxEMom
UbD5uP5untM5UFGKTLTNOu+yiR/VsKn/WjvDTqEO4RxPeXjdUowCAWUfC6CM1zgzVZHCebp4yRmW
K5B0xNlUPVt+TjAByGzHC+lQNSXCaJQGWnt+yYd9Hwh/7QTV5p6UhpOsa4GNBS4TTulUxgG388ZF
9ecrlhzz+VhHUXd18zvJ9m2uYQjlpOeW2lteZOWK8iSzIdyfhSf1ukmqLxPr40VSqUT+u34l9YEn
wVXCgPFN1mTOuiU49i2TpYsg/QWcnOFrj8/QbYWhKUQ9A+2GfTL5PKmjb+1zxbGkJAmvtKgfWU3w
MLOphcSbWHxPzxMo08JdFgzSYQYoKTlXgXalBPL/Nb/h0RDt/hTYuEXasaO7ezu0nL2ahboQ3Z3U
wBX8X8sQgzPEE1EiEBkRXZv9KmKmHsyrvfETVUQzCv3DyKD9R/C0S26TFPu6RPPlCmvIsZvteLED
aiSI8/mb7o8mvntRtWoB32WnQm7iax2N1CHPRhupF+0+vojqLg0XkwK83iObJ8KDVOxTA2t/Pvfs
ecDRFNA6sOYf+DG4ehPJm0F5mh3So8iZY5+I44SPJyKq2Q+C4BYyyraK0r4smQWmxYSMgWSV4wOP
Z7VGK+bakw79OzDcgQr2F4+H/6qKt/yU8E66k9bkVvBEUAp/5gs9u+ykS+TZmp7Ph8ng9OzqWDX4
UQwRrQdnHz9iFa1D5BUATd9XIbvdx4/V1aK2plMXcVMLYi2Z1gAY6nHzUwqWjvOqXTfpRNgE0qgB
nfOgD4UmBmI8zQbj1d5cRQVBTMyMfcFX+U7fnqIREREXkI4NeBh7EfDjEAXcmGvYXD7kSeSAYkGF
LNIrsK5hIQZl6MXGTSANdQm1PSYIleYJLc9jHF+Sc3xcxLXQa8nD9uwRE2nYFDDj7wJwhys2/0ZR
4MZX+N12BHbG8LROno45rtvNnjlK9mCxTg9EcwqNpktXMLjJSohfsY1sfGx2SsF4ywGLdzeLQrAi
nYHz+7CDfkZ7JDU9WkVYRKuPSgUSQeP0hE4Wjm529LMoJxrQGMSKUy9T7gY7fBtwhHUKH98LVycw
ZVf4ROitKcXcU6nv3zC0kQnams5PBTNWcpPJ4CVR51My0Q02z2h7TBU+47a0FIKrR1rzhwjm1hth
jjfScD2RPufd5sLQLZAOMY/XLBFDaTAv3J/Z920fzQbzm8VDRShsmEnParAaQF0yVC7Vaky9Qy7X
CdbfnxGhfbsIsxIaEQNJaxuTJ1DrZUIF8DZUHstIw/tLf4BdcIGE1LRZhearIFg42di8yDd+OL3H
L7vVIgAMeQB210dIl9JqO1/2/XYyPQ2s0PsaPbYkj+eTO/GLGJ4hVBeNTXzaFnXqzxBDL8la8s4q
jOMMup6c5ndPl02vMRqKTNHEpa7iaRfdIM31mKlIotcr4AzeHmUqd/1cqYDEdh3i/v3g0lQNTy6P
Xu9skPYlvBj2B/9pa0Enpwycu3aAxO8YRM1R+IksqaLwGwJGme200JvTR9quFraGhs9LyZ0uEv/i
QFEgBOc/LEnGaUSz95in/89MHK+PkXHFoknAa9C1OoVdshDfNaUy7qVCkZYZSElHAqWiArA3YX5B
JSABBH2A4o1txW6kwPpMafI7NZ9+2KtXRVUvkHtTQYmfSW8GajLi3iBn+8TQ3cms2DyJP/+LvMzS
HgKeZU8G1lFAHtIWUJsYBARNe70/ztQSmlS90/veN2YYzBY9ZlJX1+HYhI+8xbD3QjyZexCT3DMz
2D4N3GG7JlGFIz6pzaLnjSHvv+azRMHHRJzvaPzpIRplWB9ZyeK3kqsb2PlK67t9I81L2Z8CjQ7+
6mSQAaBBdh425xx6ke2YT3dYY3RKatd+dOxJ0DlJq0WRFF7qTwqaljVvskMz0TIa5nQzj9SCG281
HbP6fOhTd79kKBBQhpXEA2S2et3pIs5QaPdHaj5T+C9AHUEmKXqTfEIlv9SR0DA91arV0yHfdcXO
MGgtunlDst7tM+iWJQk2yTSsrt293TMoIy+QRhGKrCE4k5lD4VFZ5l4136kfklRodd5N25xj0slQ
bOwySThRiGSNBvN6erfUcxENwAbGgO086GvVVflGZ3SxbJC4ml9LZP+xQZ+qFvW/4MhaUf4VJzQ4
48GWrylW1lDwjxb0oQoo18m7xKeRtIcElkzZUyCkG+bY0My5UjxsVsMfRsg0MArel9mB7NKQbtMR
+Wux31TJjLpwerxBDBjf+AwSLomz2onO3VbKBN7dQ8w3i663vA3yNl+Q6cWQxwMCGBNKqIU8jjzw
gQcA2sZdmu59uFWmbKoGzM/IMaTwGZqFbgccoeU+ULK86FVrzyytDSGDBNFFvmo/w0FTa1Run7XO
Dl4YCeZzXwuLdccWSyD5one54dKe6RkyViY386hG66cTrVlHGzoG50rrDNOkxmjBDdn6tCnZEyZd
M0OSPMrnhyTss8AqMi8Lh47l7j2ekpP1EWX9uJOLgw1/mJhVWp/lD9S4wTXrMbahBrvp1FiseHvx
axhV0oGkDZ8FdrdsvdKLlIfN5tJPONGLSZl0/jDekzhhMZ9FqrCG5C2m5E8EuFKMFERRg7UXCdAE
2FOK7eZ1jROtEdcC0u+EKBxAPKeFKjc/l97izFKk5jfuFJ744viCpsydP0KnvryCuiCiUw1KMKS0
PVu1UMdRci63fK6zsmkd4xKHvYwzNTwzFhNsL2zuKSvYpt6siVBtpQEXeNyFk0/viOeKy3Qq4qwC
d9IFe8wwqlEFyDOtZR4j/he8t9AesMJiqbAQNn4cNIZ/Hpy/mbRSmlVE0blzjwviedGlGULhH6XB
5Dg1fb+rHnsjlW3mtt9gPGYV16jyLXODGCHYj6pqSB9V/hYvCbiGVHxkej5TspwbVxI7vmCnqSZD
NhOinC2Blj70sq3nB1ahQUw+djk37xfrCf7bUdHa3eQ7Z2Z6U3XnvVsVD9n0k94FEfg2IMhHwLvR
FT/j3GneUbE5pcpRccNKmdyDTup620vbeaYRh5nLgkMslhyOe+lrLLcCh+4EBz7Emonn8qYx9Y7V
w+oPp7Bg3gkiCyrvqog8OBSDgeqbGEAIcci8VKAz54dZkhiTeRZ70Wcn4BRhWvKsOyqZD9A3tlhi
y1apDT/Ukk7JmYMg67c+2slhJp9ap4psyDm0X+DzOZ0rwnlE5ZdwXIClFj4iKDwwA9rP+2QAxvXP
SHYh/giBc+hEf5A+S6jp38CVUpXoRtVQU90YCkhT50kjAPLguON2BfFjVY3nzbBdxJbBae0Xywu/
bsBnTCp8cRADZc5+VpJwH4tJORwHbJe077Dy1PaUWmp2WY3sL0yuUFNuCLux+GEUIjcrh8fFWg6H
a4O/qcvhnk0krrPN8EzNNPZFp4JdiYf+7hC/lX63JYBwqnFqVR4YsYnfXjNUgr/u5CdjR+RAEtkG
CO1J3EyEOQSiGpz2DpaMwa3ZVhNk52u8g3Mrwxw4gj+ANlst2oH29R5LPyNewcEO+15vGh264Wji
l5PkCYCu5mrnJ6tqdg2Xcy/HNZ+pSxJ/j2GzCtzg8SLtPKsRFOlbX858V+mUw2524nC9Uy0B1ISt
an+DcZP77sbficQOCQc4pefUhUHgnRUQQXJRKze+lCX39l1gHUKZ2fyUnLH71vo18aHIfqkQUmyJ
fnTKsNgfKeArknzKfyBFvZ8SsvfrFclFBgA7O3oYKWKt1gjFN0hPh+ZNPXC5cl72+o94W5I5Iksl
t7Ws23TuP3lfxmVIhNeeHcDPJBanPLHw5K8f6cDS5FiyymTC5sKbfCVlgaFWcHK5poYOBA/DJFjt
NIIdvD/lWLthSMDZ80NvDyo1pFRFl0bStNkOQRWNJFEjTnbb5y3KZhj6muqyRVwi62Wg9PFWFp2y
CQmpd4Fi3iPH5Z76CPvdFZcN9BdWzSoCXRQHE+HWm6nupfl1AtKU4k7BtAqCChq+DGQtD1IrR3Wb
0TMhkWLHMhiQ7dX0IVz2RMptaQ+Bb5uSQfnLHcRvmNtuRRe+1ryDLzOScO7ay+k4At/iUtO3ISeI
6RXLb/LR0JCU9wWuXgf1bLQDtkEF1fGwmm/jh+knPDcUvbG/A5pH4VrvvfUSO48UAZ+vBeDgi15S
/WLO6z591cyq2OxR1Jam1N4hQLDameU4l6aUT9khjlk5kzOgZ7aUiZAaQB+dcXf3DiLX8VLi8DDW
+YCb9uMkJIfqhLbTtkkfuCKsR+A4cDCMaMWNzWngWozZURYPEh2fZhaRN8wVnnGsvc3JM/dN7E2Q
XNVFZiaUzvga3IX77Ykk3R8WKawX7YvYJKXc6Q49dxZwDCAI9U+gHLaFlr75UHpWffXYh3i6SVR8
ghOjOiWT3dcB28vRRKTiGXd+LSdSPZyF8VgujFXgemR+hsgeVwQ+nNu34EnnQNRNRhgrAdesYURR
HehPsXNAZCySjzHK0D4si53q7QZN+6wF/u5n7p/9jkkwe/LXZu83/ThXDcd7cMnehI4OSNg9VWGK
56JRbeEblN9ai1J08ZXf8oL5bQud9mgn+vzZhit3B0ElUdQidOXXfSwCmNMi66P+IPnc/6ppLP7s
8gEi4d+Ku6MHDQNbLIDfngyfMGt3aSiujyC+Xp5ZjUim7Y9hetysC/jcZchabFOyyjQatdljb9GD
IiE3frBBlReeCZIQX0M9x4nJf8KiSpLsY94EIJI7BfdBkyZOe8vxKCwsYJOaif/K2u8RQ/WKFY4B
TqtKcVWfW0ifCrbcifWBCYQzXnOhLayVo2aTv6tMqa66KzIP+QqcSdKzieDSICrdtbYSegVnmLOv
d2dHZZHGs8iPvY3VmyM8wibJhUxMceLpI8ZllNBBytP5AgXgUe9KW5h1O4aLDAlPj8IspNdcXXEE
QwOcfvuL6pSFbZHcbLaV84RmFL8RvDr+NJ+Mxpunh+y87CSpgyAPTEgpzayeaL8DW2YVin1bhRAZ
Iy5uIe3apKs3oAnZbdOwSjr1pzwNAvTus4bsr/CRCSdyUak7ZktBlFpaag4nLM0aWj9QhAOJ5SRR
ztxob5ToXtj1Z+w2s31MdTiKDiitqbvFqjCU+AHU2Epm6SyCE0DSIDszQ4N/+CkddKLwgqLdb7MQ
XNwFS4yRLv0eqh2L5nqPd0GfeTazu5OeZPHmiZJ1A9lFL0t+mqf7aZG4t2iTKGRWYnLnTef4HqhZ
5HR864d1+D8w8HndnAoa/kKSr/FcgzUSuo7/zJatUESp8XZtzNA25Pa9csYarthZYckwVl3gSHtZ
iFEnyX+bjGnbYgkh6jVIf3Jb4NZrI3G95W6ezwT4hQqdDVacpUM6SV0pCjq4JZzEBy+/Lb7uyAUF
8bLsrGOgxBmmupaxtJR3ATpeS3IyFuqQAU1gzTNpdUuV+HR2VOP5qTr2jKbQb521zmDaIL0/oEFy
yObWvmFbC1O2lM5iUPCBPJkxMKNRlmkbYy7lvvrEG5vsu0yrm/1mWFbymCYy9Qj3sLHIOcwyc2LB
2uRvp2txj0OFLyii8ZTVKwI0MONe8+Hd1PjIqgS44SXZ+SDy2rO8r5T6YHcgvL//MHTaXs4bbw4C
YEv1d+rsz9tvyIvuN7Kjpuopa6oSyisLChpush6BOORhCgc25uCtCIb0zCrwxH6HB++e7ulQMPvF
0Oaty90f/jkma7GRnOigvNm9myeYKfhqonhmFr4/7rzECVqpaCJZczeXlHZRfuiX/5okhZYy8R9u
mM5WKyqzmoT2LmpU6INV4Sm1Q+eerV3CblPZvW0FTo31o2LyHjWM12V362NT9yBRX7/JhboalHSY
FFJKVEz/MD7AOWZy9EE2MGMmpjg3DVPN9Sli9OcOToZDmxQO8IXVBC+dMKIUcdufu6aW8rybm03u
4SFaNPbAQN09UppiBrRbxf90tk7UHIj9TAxwpnr4RukvtPZF6hhmE4KLkfn2HwfQ87vgXMa7chmW
FkjZG0pw2Tvfc76q8/gicrJt/DEWehhvnrFb6B+ZjIOaDo0XndadNP6hFNIt9OoojRHJswFkHSsu
2wJv+SAQl59f4SnhEvJZs331ngVkbJf9RanPZpmxMiRvAEtj4b6Wi0za7TlZaQfqQO52O+1DL4VM
IALPD6gn5/ASSq67pLXVlTasylxnU+yvA6KYOnG/OnZh6zU6934JfK2Gsh5jdfWj1YmJfwnkWfHr
kMZLOcRyhl3WgcObmar/Os3JEIaHg1xfdXFxMiEc0h87Xig7hV4aO2s206jiqeAsy6Jl3cwgzxhL
t/4GGB/ThBiw0b0M+IZXldtfVz4M8u1WFP1mMMaFF8pRlXe5FnlXmgGQ+HyQTPfbSSJjAZu6rXB/
LTDKsj5tO3J8nKVTDrbbscGMng00CyZyM3///OT/YOQTcKrN8yq6Ee8iGTXgcS1UyFXjTJo8juNR
Tnst9oh0t+kfrVDChWOFehulGBvt+yWRnIRXgxmlWuOYt2OOHuUkv4GZnUbTQB3x9KMgx+PjaaeR
1NND5Pc9ZoQUnlUhHz/F6wh4GyUqpclGtBDr3suEbuNP2bH0KT5TEuPLgDpU419ZYOGG2ngDyB/r
w/zu6jUP+qODbtS2XN1GXZHiXSW3997rFyfT19tRODIhP/8Bb8EgWqeScAFbCYnbxPEfR+mwQLug
ZCcbp8ut+ODmJN6N7VVCsv0yneavt9a7tvLEAXsX3GUsdskZWs0U/glJcVqck1sLMrLMe/uVSMo5
Cy2nskke2VS2D8hBLz/M6aHSu48DbWVNNA5y753DAdUsuFGRGHVRXmaBOPVOc52goQBEfAl/Numo
Uj02+p1OgeXgvLpNS5EbPdv0qxaUxx668PwzxzywODIr73ZFkTeUrLQoIlZ/zIsGXkYy0a/PszH2
Yu+8wZVrAXVIXXwKk5OOh/t82MvkOguR0fJttMRWsDKnv+0i+LUNMbZYDbpawOYIefBtrtZXKQ88
l3RJoBsqMzjNtuQRau+pqrSwthCF7MjOPnv94bfjT0AmEhRRb/dvjTxHfA7qmfrmlSTNmQHBbV8B
Hfi+tOExOBg5m479Zzlq/nElLl+g2Lcyi/+6T4aJuK5gP98uE12nHBRSPLBGZ+9T3sKlMoz0S5ed
U4uY7JfVN0GxZUSdWROIs5zuid9Xw9B3Xz68XIIZ6WYur98nC1bIsC5s/uqjudASyycpzQ5MCqFG
2gKT78RjP25eLnKPIEp4l2B61tTCPmU8UBc5vygAWjnnNXJYDJc5wWkAPvhZOPH6YTcBeb0gKHOX
UNPGKyEiYhXpeq0Z4T+fXJ8YKxYj9U8gDB8mQoDlBw5OyC5qIwi7OAmjLW/kq6R7IMZeoJSTSFtj
XGlGKqb0w2Y6oq61MGKOlyDB6q3gaMMz+CKRng+usMBJR0VosirilZmwRBFFLJw661k9LnqNHx3A
01/CTSYfdy8VsuzRmqDYZbmaBgusKD7N0rSA8P9AmKr+dcB/v1RTzavLMdY+25iHHy5S0I3pBsGt
3x23PaI4yC7ROrZXS3KR40wEO+bYx1auKn8szv0BxnyiD8febcM/bvpbQA/isELsxWMs48O2OPfL
aZbEeOGeM1B2IGrXRitQ7R3tGg2Bu88Gl6Emekmyt+Pg9Bsl0S1Ol/Ki
`protect end_protected
