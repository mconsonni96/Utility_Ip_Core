`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ExdmeSzx2yiXNTRx0iOb8x8g1iygngLerKelqS8d3BJooXT4V3zgid3d5Zj0PFORLIFpw7H9GnYH
HuxGAQ/K9ziZHHRe7fGbm6+FPxhhDEQi4RCb3IpgkID2OrD11XzIdMI2xnP/GCJAqBEeVCauL/yN
QRdGw78gO4WYM3ORyZGP2f0Mq8uvtZ/hf1JDZukWEOBRUH3mnUKpN+6FY4BdhtxPdig2e4OZBT3e
41snze0PAbDd5PfOMmz6QMySc02eSFtM++sWzuJDuAIOhb39BLPGTgy+2QhsVX+TfuYPyNvBOxWz
IgjtzxzXEWPqVv8LYPSse4GwxHyo/9Jf7y1Zfg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="oj/2n2Ow767vsfpLmMnoi1JxFdtv6XSocxNC83tvOUg="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12832)
`protect data_block
PZpx4F6kgLnC0w5cn2zEzNshRgV8wA8JM5rr8i7ETpeVgAG7jNkKpV4SkWcYAO43nCiASK7Wgdp7
VJG5D8uaywd1wUF8LMW07xIlW7VyWz8F2XemQQbQuuLpoqccN+gXy3QS8WBW285dkSGjyZxFFRCn
oPA+MRLpGVqoaUHgg7XsvwtnKBiGEUaE49kkTKEpI081oNmMdQ6CIDYDTXG90jlEom6mfNYdWtBU
kQuDZZ3fA2hv08kYB70LMggGd9SPzaqkm7i+je7N2Tb2npLwLt+rWTo28IRt0e7zx8At4rjy4Mq9
0b6EvsD8LWAZvaUEBJ4VtCZqmjfiFNO20XvrhrXMIVgkTWwqr+AQU89gKzPBAZl5Qak0owaU5wZN
Mkv46vBgUExZAcKr4cLU2aiOCAFd0Do3mFEl+V0HOGeRnft+x2hkiZWa5L/iambm0MHOhdNzTUP/
foGNmnCTUEr/EQKGWLVB1ngQJS8YrTSUCIOWRWTSRdD9aIpBbcD591lvng7BDMnnwnMl5M+VJC5f
vjR9DhjSRrVED+nhfwB6GlBcx47fhhDz8wjGjkRDhJngWemTSduMVHVPcFScW/gpqpAXUW97T7U+
9tN5y5nj9oQk9chH47x9fpRUAxMvBMkfu6jJ4x5pGn5yLUJor+AFbHV5ZPRo15MzYCNLpt4/ykMA
rJvaVWRV/jM4wUg/C9GWhrUapTYW6xnGcDeWeI5Y4FU7ZThxYNagWdktWSQKQ8vG1dtohW/HxOoJ
0E7OtR7DrDO7b/ZGb7yh/tLmEBo4qX1F359Hc99Fqf829LIRdTK0GPyHLKpYEr2ApU40bp6TjgYX
2RNx1CX60vpmkB1ziPa1KA/I1woaxQTjs9TSDs+9g6JUjiy4SyLqlBfjQVf4/Db88vJj/53SVuY2
1GXACaQ49XcYP61xXCzTbWRZUPoXVz2ChmEaleNR1lZOd0r7t/h5qP8UJjJIUIbs3LZ0dTWsJGam
OcRg1u46CXeV3ze0UDLUULbaeqAE8At7su95R0oWqoqU156YqB2E86I+mfCD+X3mtNAutDXe3SNV
Zg/6b8nRqolIsR2cCu8CE/6PuPo0wyNnDbRUYVKtKs5AP6r3AlU4xyPbCNLaFIq5SqfZNaGrUePU
fsJtZlGY2ANs/X0prpf951Zxc81JNWwkR9igBxVJgXLDdXKRfnzNRb8SpxgFRFiT3RVEIV5d0gbG
7ee2WqY2gB9jY5rHKyYhprtNbcEvxzsXasHgxFE80jfuSRe6tVVKyqoB6G7g6WbhA2zkIUTFrkXT
2pGBbjm9CgOU8M3DvOTVFsEw6tcM9MjtUKzhyqGXoHZjdnJQaagWODBjImfWLqoNKoODxxoMAwkQ
59Ewsk32ZhcPjyAf+/ZSKlF5Ldq+7ezJShWtBjsU/65DckdvLvUOQfcGc5tU1W1dIMVGGiKodLSX
+C2mRdiFLNZtgvk/Db4qssBHujp0oC4acTmu1ZzEzDNvn+TbKYiFxa+7J+B+BtSFE5+Jt8dagR2+
EKvoTtRkHTsKiRL8P6Xf4liyxO4O0CHvE4wXRLYRxs1ckw1d9aBBhoLHOMzXDSoCHEyEmteGDBL5
DbxognWbvWCw9rfu2bTlGQzYCSmJhyOPwnKMIIm2+qCkc/XkD/9OrNcISkLfuzMDVfVSsODngRXz
mLLbSSEMLrAZnGA5afzA0h7LiRLxOOzWPtSCHC8UrF5vAy+oTawjRzkeFg8XQqHBrydMh0u6FT+Q
ap66tnWQxrBOsmO38Z8PvChFNu9YZVM63oYzp3c4LPTxuKPX2mPsxtRJq8SsaTaH0rAXrVrJI4wL
mGh+g9wPKyrsLaMzMPW9DD5aUPxYtHZxZkwIgkSm7jU8stjM0macPDRc6JGrD54lO2FGCXnNqs3E
dM6w+ztowI2uFl2T8IYbh0cd5dG3md7Ak8Um3MSKD7mtDA2B60k8xzyQBE2m14Xda7aLSksCmTxH
SZw3NjMIcfthnxiwn89Cxs7UxcJdKE2pDen8ueIMMTlZyGgLolZbjvqh2mMPV9uyKGiZ+8FPaC/O
I+Vr+JmgSxlDtej/hCiHSd0to5/O9dq9H+0AzYo8gHf4QPGiKr0N2u7MnewMAxIcUZV+M4ih4Mkx
9gVoSSH5qbXsP1XoJp4g+VxGBOJ/YNdIqYXEoQx4mHV3vWgbsrMHhyRDff3/PgKzwa6/C7XtZjrh
ZhqxvdLJr9Toxi40QwFMRjHUWO/qYxe8ey3fceDNobOKRYWYuffVy82/LerZKhmrinlJIa1CY8/t
3AJsg0aSQLQx4QC5CyshekZlCoXy5n983DtEfIaN7GLKh+jQAQK9QNfRJhvjM022TEUz3bZF5Un0
zLLI+UC31u4lgmEfZOsfYIXR72shJircDg5fxK6nHX5OTA4TgfWOYogO+exRXzFJ2ZFXBIixiNqF
mwGfS3SiPRyiI3oZxc3+3aRsZyE6Mmaq7nGN0G9SiGGmtRNm3TI3sodD7K3SCP/JXgxvLdUV8R+C
BWkwX4UT93uXcQqCqQ5pQXz249THGd6s5oUhxx2GUF8GQIE0RwKNNKDmpcsyuKjcB32R+sGCb0hP
vH/hTesvZgHlaucu8S5B7UfM4uofD+4MKzlqCAyNLK2mAY7H60zLEzgsP89ppMYtCtpZT4iKFfMi
9gXZ4k/q1DNG+WEOOSuXgDE2meIAxEZ9PKYamz6ua48zkXlXv0R3LSBSbLPtHI6/zpLhX4R8rdik
9fLUUNtoObp2Mu3O83o2nPrtQhVKiJydEtEDP8uHJXYLv9JDkr8+3cQWvGUvkaHflyzO4Q5CPgPk
V5BuI6gptJs+RBB8Mbau8S5i6ejjoZeMk6nS12S8PJ4GC9CDUhqG5pQTPxGW/MrRMzNItxeHnHhf
fWXE4E6k15apoHjXBl/PCkYPinXzx8/uD81/FWqbIirzWBam/r5LCouKwAJVPRKDI68X0eLiyJKH
IFnPk6KGmb9EEc5quPiCeOxilbgugWLpYmiGBrIUi1fE6tKz+sq4Wf4AZaxD12vVEOLR60OHnGQv
NyDz7XcOyyf/Qs+3O1ogifPEvcsD63pWJxEIDfa1YIHVe65XW4mAnbe2WTsqGAVYko6dWQ9MUSwN
bFhirhzTjcuKlgZ0qUmQSk7uZyb6esiKLwKrVyknCjvT/Lt54LvsiQq8tEf/+Cu0kxKj3u4KbluN
8bpEWrfhvjpbQE+ygR+EzOGyMqc/0v1vTsw5TTMxrgEDpulZ7Kz17J7dYFUCMEPzLsJf/ijqZcg1
s7U4bpHtnf2IrvebdNQMPR+pgKfxHRwvC7QtPEpXf8umwNzafMkGBKGD/qdQrOvRBnbaOXsCDOXe
ke7Bwk+AGmrfYvEqLyoe1VAccECvieikuox8HzsEvkb7qG+CTBNsV+OG7w/LFldd0+IrB5f92n8W
86ej+gaRQDg5GqnN4GtG6V9L8Pn4YzfF/XAE/kkb5l2rY9dqmXNSEZYkIn5MdY7YMsRdTZGp3YAF
S/W9yejP6el/TBS0jhK0A/thmO7JMmHkessNSoT+05RtbhiVBWWcMBlt4GRJqUzst3ig/Ohl/ADe
edF1l/hzOwWs0TnRki9EJzSNt4ct7ypH+J8L4DgVhpyQ1ayDpvgTk/Xb1GA8hcrhl82WSi0yihUd
2TW/PVjmDpnor5iqxN5OdH9mQvAYd0ZgDW2kCX6p+ODQ5x16nZiUrlVBDTRfGSk07wem2Hoy0ntt
SOwfzaJo8JBOq2NDc4n2pFizOjvHvr41gROy8DAKx2P+5IImrxAp5KmK2IfE8118hC0tX4tHmLEj
hwxNVf1/1VUE78CdxWcGelLe6mKkmgXlKH/Of5rwgldPehGVWmbWXKSgU92bfc8xPul3xv1rAChk
YK+YKGhUZnqGUUv9KjgTGe4ZsxVLH5dsbz8xdFWlJ/zGNJh6wTvzoU7NdvuHe43H2IyurzANBcXd
f8IBLrSBqt2UPDrZ4FbMfjM7PT59GW5m1aYF3bAMeyLJqBUvHlg87Zz2y9paDG1QGY7LqrsXh6/Y
ZlGf8L4pU4awro4abGRZeGbpytDOV9exVKf/dyZWNeTauXg5x8jcNpktpybZBrWX2dobL5z8FtlJ
ZKlqKTQdPadm3U/LB45cos8ZDgdHnwvC9+AuhHZxEGnykY74gJSQyLqIMVgfPApZsvsdY3rjplza
PlxGtt2FVTs2bRRYTSzCg69NcGpAzw0MMyscszl6YtSOlu7U6VqX2gTDieHNb8p/0ypsfE3MCrUa
rDecTcGk6D3TEh3q8ToctKEwk4X/NsbH2s+aoOYe8BRWYsBUEZ39a1IdX5iEgUhd98fHP9dOs+md
9GdKI+1B087wQNB4PBezozkt7BTEkMAGHrcf+tS5+gEwnbI4V9sMz5XeQ/Yk6qmqiXmPzJFT/mwk
/ZIZkjsPinSJjLLEe4QAmDJ3BN3bRkor7giH9IeM68ww9RQwUpXFVaX0R4VN7tcryRaDPT+zXd6C
2xYY1cEeWnQT20ylwjLzKZxi6AnO8MwT27euULIB4V4RpGdG/q7g1Xr1+EPCtgTeRFd/ccOwAY7F
EepRcC4xHkWNxyW90IxB/7ineqktouHUO9IpJ0islgrJ2xqTIKUqGsqDHvorn/SDDsH9U229KpMb
mb14X0Id4fhV1PUuIM7WynqGjsAGlmPCy0oNuxrWKEC5X/0O+z/dERV348dtynkALTvM6jzTAB4+
62JfQJywCU8qa8XcRnGakJlcfwya4gJB6TSu9JBnt8FQ3xbQBLM6Wa4cztkJ++vvFysxauOhsCeL
vmMUmEKUcQPSIqhWIOvY4Ue6guV8N4CtWjDoYmuTqUzAYGj4QcvHh9j+9AM9UfbJXBYUYmwhbP7t
pJDK0/a3BEqNxvYAeJ0uYok+ISeyS1ZdHnkUe/06f9jsatGEDV4VYBY+8nHtKAcVRHKCYbVNeqfu
478lwm9WdXJgHMwOmUGybib/x+gDqXKsdVi3h7YNoTepNs6HTTrwDYPznU4QseXobIAjLRNBtzJg
JQl7xR4fkEgE0SY3xyK+DZ0ln3WKAAaLr60HFDUyqfx2MVSRTzsWt5+tz1k0sgg6d/TOlKS9xG2u
Q8c7mdXT02XrhtXAAoYppCogVnd6vwA2i9+RfCwa3xZ0rNodfX4zdwc20E4YxKO2trOx1v6ZFg+x
xINiRyVt/foWPOY+9rri0P9fxz7/U5ptB0XS4YPRKhO+gjWhOUkLy9vb3SVDIW96r20zwMOJeJxF
XLZNA/xzVrNsNZfpgUtFrPioYipIVkRPnU3nlC5dcSa8O1+nYp49TDZwl96wvtW36Tb+XUCywjH9
Zk6asVyOeWa0+4mh+rOmZVU+MrcekUjDq8AMAZhgQ3BnDUm7m6yHEYUoZ9P2RWUmx96JsWNPuai9
wDPqONfTo7KGwl6Ycak5OUS6mz5qSksxkHdo4rzVPABWe6b1fPhQf/Vp+aYROUxRF1ojIqPaN4c3
04q4rZNpqct4xsptX+Rp7TAwcEk/Q7eRw38A0DrwO9nJTZg7Whmowe/GXYgtN46RI+ALhG/zjGGY
PRYSugpyfRe6bTiVU8i+3aZo3RcnTkYAdVwJOrZJ10pd93Rt7vGfG5T1BjDoreQkzjkU5asj1tag
zF9qkkQ1k3KGRTShqjr9HUPUrxOMuSNHHK2Nb5saAVrFuFF3vs/uubq0rh0L5iWSdB3BZcs0AB9P
cqTtnPzopyI9RT8gGpT/hb/nACnYgTViSrDpTAKS09qdQ8ZdP3GDS3uXifrtkZKYx+exniRflYnm
6Rd7f0cR9Yl3uRGatQiC1HhStIYkXo9PMuPGjSHBnKS8JqAgKyj7jgvA48E30KRkco6UaJx8iP+o
02fBEN5k0QOyCdlpJrO8dGJrgsavliJWJ7/gFA1mrLJFjqonyBFqVJwjuijPSuM831TE0LiiAP5G
bAw2WCgm3oyfem4I+Lm30WwvYMk7mCZ2NN7485hA9lixu3RWIHZNX3h44kay4qioeMNngUoN5Dpj
zTer2U0lIz6R0emdxz77TOZwtBnxkKWsuJYju0BKy/gtBBaowOei4TImhhH88rGmJGgbwUkEo5Y9
IelEAy2l/j3eS5kwe42zU/C/d0OWtKv55RlV2/IsuZmB/qx8fE3NT7BvUSRCsMI5ACqYgjF4NFRe
YxEC1CmuPaHsT6XG58VmNKhWw9MQMPpUpW1WVypyHY9dBNNX4UpcbnHUzH5Yg1LOdc8geFnxTk5h
C9iqQc9HsWFnvKZ671HtqN3Bxk914GrxGN6Xbe+nOUNEbY25S0wwmKZXvvGEd+ca+ynRyoH8CPSd
mD+JWfInfwJnzMs1fQ9Ze5DqBypNSe+G6WFyYU7Qpc19hA5V1qwyyMdYPirZNJEDY8eD7Sl4jVkF
asav8lsRji5Qzk9797X+FU7Bg1RigY6qGSTTmHY9xP1p8oCAa3doy108qJNdE5pdOoFn/tZgiKdp
EdySNuM5osfAPtySFGSokkuJyBdDRlXwnWP73jDcmaaYlAQE4Gm7F8vQEG992Vf489+el3xAPcGW
zyreNSrir3Ni3bi/ml8Zt7HJxEOG++dakQSPV1Xf/UKrZvpoloQQzgCyaiJqmZ5/jPB6pc4EEeqD
3W+FaYmapMipPI6pU7Q+ybrM4ItAlWv2veezuMdVJadTy2mbAnjCkmaLB9rHoOgop8J2rAut2HbZ
5SV65st167Lxx275eUbPPooZ7rOXvm9fvCDylgzEpykkSGTDOX1MYSXllgs4/Ig4KZOPWmx5VlNm
yeVza9lK3i8la2d+8oOlUoRRPIM96DmwbyBg01F2ElBaP3oBirDi+4tSbuAyH2DCWDeIKrcKeH0a
h75X4blXu4X7Q/OtD4Ebo31ot0iOG454AEFdALmVoWHjM59R7dZEj1RW2GurZoXxaKFlokYpcvB9
a0GEpQstdj4URcvoZ8lHBLkCUZQIEatHDyrwYibA8bfdY70ap+CbDw3+i1Ed+KaGqE518JKzIawO
LcDa8NdlZ9PXK0MiEC/E0FIUzIrL2XNgqBcokYk2f7Iox61tSRDO8VleE5/rW1MaDoHbw3sDXyKb
DL0qPykTfzt6cGsT2aZk3jF9Ixcp0HWkYaq0ht/jBXmy7Er47HjM0mwkmjMIWeXggiKOnIac5R9r
wUaFVNT1SKTfUO3nH1UbneEjc7vUdvxip/yhUFpm2dtDrV9yOutShbmhrOC2M+FcQ8ouY6F2qcJw
4kkFfkPQFKYN0hEWQQB3FKUALXD4sp47r0tpOl1/OHvgmtRqrTqySpNmJeK12qN4VD545lLdZvWZ
J1GVsGaGuSfEjbRuCfQSZ0FINc7rRAblNM/YKZudB8JiNUh/TBz3qafo6jSYMRmaqaKUIxZ6NC7+
fbNvJSU6osAG88hYXfRtFGtLKQTyCcX9luuczPXauxWoPEQOsNQresgU0HxuUDzVpm8j9GoPzgqz
3QamrK0bR+uuvGPtulgrSd2ShSjbbJ+Lx1oCRCNVJSHlDVFwNBLoecBhyhto5ep5XkFiPKXWtqQb
c+C0LoKYM6wGYqVEmGNxc+N6PG9PEyOWQRJr9cQSBihiTONjKYWIY+x9CYzSkStkxoMKUV0DM8zK
BCfasmfOiSHxMFIx84PBPlPhQpOepL59IuD3vOpIUt+wx6lbx11HX3XYbE3g5/9RW6q3cG/H2kW1
b6QMvKzbdRrP2Jfae1qffSZ2lsX0z/UvxDDdmgECCpKB2hDKuXGa9QvC/v5X1M7SvZDe2wcRTepD
Truld3Aci7YJMZ7TNPbDh4tqO+iUvJwxyH6axeO1uqDUk3JIRDtHtDycVyRro9IszJk+2cQ15aVv
lWGao6owbXu1CFD22ijc7ODISNSJ5RZVfL/I5qMrVIxDQ1miJltHTUWeHN6ZhXFUWhTJFHtWnln4
FGoxVy1bqFq+nR6Fpg3LO3Yh+qrpObmDvzMFVRoTwzIeNQf7m8v492qiY7Qe6lKNLRTKzVBJ1F4N
J1xFR7izoaOkN2bx1s5XUws2aDpWLULIpk2+DKIDP7CFrk1MhuLD4pJPKpNa1jte/LuR492Vj9dV
/n2MVloQQ71Ruhi3+G/C9AppXrvJIKefG+ycjHOBwPsNKlMyVbLZ8CvXxBAhm9PG4lxLjCLdd6YS
MBKXGhkGPwampaTOebWPUIbG/ZfC5TQ9193uxpe2mwTcULYCOE4TtlFgxlWSYw7Dvp4WA1NolLTJ
y2f9uCGaP9prt93qQcTcxMtK2IYlb/spq2qP4F3q/6TYakeu5P87Uv0ahYgMvNvTrTxLLeevRYRX
BUFO+8RvqV3dFtSbuLP1HU6bVpxjOEhqaXXu+ZEPhVRULd67e+CbzvOf2uF/LCV4J6g2k3+qaka4
ZReNj65SwmPF5nLxcrDC36n/VjffISUsak0P/Gr0e+QtuwyM16THO5SN6f7oRPj6pnsDSk7R/sKH
1OO66g6eCGs0Sq4iS2GtArnnI3oaoDIOMoT7yzdQDmR+WTKRCjXWEmtt3jrcd4zyICFFEdgOUy6a
vBfKDn+hD76CJeOg44SJKPfc8Xw1w3wd8XOJshzX2QVp4um9u2XO0sr6iuR0ZZqM5HmOyZu8v42Y
DIwBYa94SEJ0jyiCCt9of6xD7rOUAtLmCIpmRQVLCbjK2cDvYdlG+RuCaxalwmSWbJDTEeKqgRAr
9tXaeMNJsnWJyG6tZFnaWgY7KRwYW+7BNSHXzwhk4Zva/BjnVDyhtGcT3DED0ygBTRDu0ZVhQTNX
KSgMwmhW9IQpDaLW3YV4ingzWrsYosSre5Dnsm01WX1wKwalCEFrMzhtkRUe1zxkehEUe1wA2oSW
liSIUr2ofledkOVFa0z5jp7WVjee4AxPcZS14bcd9uEQDyG8sJ2gyX9JtcJfetsIuLYu3OBvTZZb
A9vCyKKgoERcdKb30ZsqHpMn84Uwot+Z2RUz/Eegp3l86h5fwxxKMYjopsVVR93d2CxkOlyZ1qH+
Rtrko9hBzNfFjxkB3sBQ4MG1Le7PrVMdOmdcDZ7sgLKLbNwBbUMpLvPQXtKODx6t5C/8Uq1WenkI
+nKIl9+1xAnfQokvdKBFM+WuIohEgMjZrZnK60hA15ofvHhyGTyoFMD2I1KvhT8r0rLzz2vdUKUa
N70MjJ6QhVNjIHuh08++hZYDQR82kNcQgFt4NVIbvgd/3LNMcCaCmfsV0LeymB61cvS7iAeUdGTb
LED2JRL4hCBZywySIvcEUPPWfM7hc/efSz1VIN5w9yORCp0wpLPHI6KaY3oe0/6mFyh2iFAK+gtn
9wnF7DX3ztkP4ExPQmOGgjnEXGYDpn7GJ9r9SJjzAEWgz0MtOPbj7ccOEAbF9Mr+6mA8ufR8Idnq
7Bo9Gt01Pm6t30bTggOgjBgQXBV4ePGhDFnLoxTcRKMRwVNPjWlVECLxUC6MN3B7CdTRpp5awYRB
VNxTM0UWsTCWVV0Z21quh6nE5P8iq7mUCmc8d2bqk6Kslo0kwBkHYuBHEPPKlrO0fNezgH1VpuCW
24l6vsEeYviatAGz0zNIfw2R/PTdIfWwbLc8bizEGtcE/T0w3Vj6yNc0/rbYKkkYZ72SW6pgFVzU
efW/AjBJh7jSsqSKQvJsBIGMBS0nQIynW00UB1xboh35Pwqk0nsmZyhrhscQIQ8ZuZzLnSG8wotJ
WFySMPSmT7Clnw0gM/lkaGZeiO+gBcbAUk99/uJnG2j/GmGjbKgRksZkKBtMp2fO3yYBfJo6dskD
a4epja8NcYfqaz5ddXnd/Fp9nUoGT/0jWDe0SgQsghATgQIbRFHXMxFq/3rqKNPqU8ANf6kaXE32
PB9DSfqkZoiSa21IVdz//h1n55rhvw26VhhseZ/1AfNZ+BCjYCxu7lxQnGEhf0aEf2rgGsHRknd3
+gKIhjB5hADsZf/Uf5sIP9TFUm7+c4GCRchYYWSmpyjuAZYMYka9epYysTejvsK1J7YQPtLV92DR
m/1RBxDJHm3bvGaD3xAJzksr1vimp4ne+6OXdSezUpz5nPzUOcV9T77phrUKa5mlzDMptQuInwSr
O2Wi0TmkGPhb/VCzzt9mGTduYUOaQ1TrSCTc/8vAxCVfwsMaKLlZUeTau+GRD7DeviAeJGGrN1Gi
6/bIb/00gRGIPy9mkB3lfX+FCHLdoQs/AaFHQn0GJlvTYPHih8x4lZ3oGhc5ihYntEKg0E8Jajup
ch+uyfpvF3Nc/FjcimgiAVwNve34gwmT9O7ekyyRuzbs8IKVZRsXYejX2SfUjWtr7gaMSDkFQOEG
ZdaxigbFtGrC9+tfiSaU/cymKZK+wjCf2PFSIoLEQulU441q/TnrudwJGtf0uzFxt9wffB+rhP7i
Q4cOJyF4OqUsrLbr7MaJvW7khvh7GZ9yzSKEhkdDW2EQOrMfcW5T8REQTBciTdQWnU/pfrZxL+gd
mK1NkgNHgkhVKrgp29kGXjrprdTeRjkfvoWACyHcvPwQm8d7fGyUNE0clbw9xKx7vLyEHfgS02Ma
E5MhMakqErow7NvMgYBhweH5qCPzU939VGPtMqOAUWzjz6UHPgL6jPw+7dSiV/e/Wb76GNipiwUi
iThx2Gsyj5dpC0hWzvfgIIgwYuomu2oN0UpQFcvh/FxzDnDQDptq9sqdHw12vCZV3+hmUxayLljI
yWhReHsZ8A84PHnaNLudeZgW2b38rplI7KzBqQW8HmzS0E8Qm2unYloQBhueU2GCrLbI+Yihn+jZ
sqPKaq9FaDEhzom2pxU1DL+wRSmv7msE2aohyhneStHMtpSY5IPSzXeRlbrqOH9G7turHtht+gMR
zVmAT3pHN4GrqBP365Ihehpkm5C1Io/5q4F7d/kq4N8NYNwUjf4vowRzMTBGlhq5GipH8Jj5sAoi
eB22AOXtFFkW0fAOwPPfwW19T0jNfwN/hMBPcV0GH9jehYNTSy6c3EwKt4Pdw14/xf7JauNeej2M
jubMyn0NH7sWCuQ4MlwxIjWHkd2aIrWbJiQ8p3BtSHDjuujWZCp+o+v9GqBcrJJ9Z5G0WYYVmOvN
L996uYT7oaqUaUwOdGWYlLe/RZuR8ULp30c5gmQJ53+m+4ok4/jRjCaxAo5fBvPE56Dj5QSLEnu8
NAld1CM2axkz1KLCBvJL7pAB7l1Ka80VXJSs+NFvgIt78WasGWElMMyZw1BGafJyf1+5SHV8K69L
WB9ar8xSJKqFaGNb9koWlCXUWKhjqDqV+XhufqGwD1AAbweIdCyBFIhyWbF/+7xiWr51/hw/Hihk
30jkp3hTWDglZrOLDxRAc8WPg50RJu1l8+m+yT63Xx+2f6B/Gss54iZxHspW8HTWgLX4b6Qo8pFI
4qR5g7rZGpNjg9Jcx/o8BhX92On7WT4lg7Psf4da5m8s052ZvECrbcPxTg+GnjBTYOWpo15Xv+2w
l7AeITzGjoy1srMyTDIqahwSzPoVzpF3Z/BihhZ6i1ZETvg2TnKTEmVK14N2W90qyEChnsezBNp3
2Z3Etf5l16DuO76Qi9l1MhdTfFMMosHmfn/qrQD9DnltPsiz8ntr38rUIKWRDJs+rkeWLpl1C9m4
213PN2mzu15lGfqDgrWzO3qyGpDUa1k550Zf+r3qn9JSw81sN5m/yIELFNhinEDXg5NXQDg9sYLt
xAXK5ofAv7a9y4yDZdzSMXW3xohBkczUfVcxFTooX94lm9h9Dxv1LsrF8zbq7cDXgN9oMUanXspK
H6mz77b8btzzocdSGiHfEA9khZEmIgDGw4rt6XictGjXDJ9fRE+PU4fncuWrqaB78OupKPMIyGoN
VLc2UVvwBKXUFzTn0RbjRgwTCSJO6G5WEruGWf3LN2y15d3DyQnpPB0Wg1vUr9bgqSSfGiTzcAml
xDxNAlBi+GjTeUNd6RrN2Cpm98tg0LfE79HwyjbDBgdWUTkBlqsmxWPej4pcNdoZVF3msvs2I1+B
5CJ8Ppvytxr23KJJJOH0ByYDpo5tPelYe1fjs11pzVCLpf45iSgxDK/oTrWvLiGvOQ+p7QVmZByr
xhyVbbOzYGOw4i4lxxfr/f9uox2wHhEfnDvt+tYeVA3DGBD2a7XgEW7vdheu47/HgzC8v+jxwOyr
7F3mymekdO4hhp3qtjDY4nPpYSfqR8mRn9ut1XPZofqaB3S8g993Il7weNS29F1Immx48JgmvjQv
571I+5Vkm+XpbtgKupXa2kEGispichJmgM7RrmYXA+Pndr7Qh1tzxByfQAyHpt64z3ADS6twTzrk
IAg5uMes0yie684njYwZWbTuvC2fFVZBFdwhWpSRJnBj7rVfkrUPJYGQgI+/McXfxz3N5+T5PEdy
wONt6VVTiBOpUkhBHlXoYYauU4Lcz9MOLz2+e+NgjiTkJApmGKqiKO2wRNBvNCeoL+rn6QBtpMm9
CGjDahuk1XVw325CMvdWzn1oGwRh3CuIcmL5qf2br0ynIDruSikX0xPDChe6vpsIbG6Ry7+eaqNY
wrZ8MViYzglFb0KqWgH0AXEUYFi1SeUGW1rK0Mn9fyxeJeN3i0vDsvQ7Iy7+oPzlRbDUDg8Nzd0i
fMdu2dVabXYUDcbUwvUdABptagU1oiKfik2UVptpMw1QhP3lhFmGjZYmU0zectqfPROf/733dn8I
f3r0k2xfRIFUNP8FcZywQT6dV8a6q06BRqfhS7rswl7aLMLC/BaXNPUMr33Kmihb4X+Sxshnnu99
EBoMcuSWj0Tjdc+qCeTS91qxc887mDrKOufaAGKAsZeTfIl9L6iDwFJAdEI2q8yU6TUuDA97jXZg
VId3BYuqrAUiWpNYGiGyw22EnW63nphXbDN1nRzo1iAHRsWFZDYP3cN0iJOZG8XX0dp5YWLD5ZQp
tikeAjzqlAvIEW3Fh6lE6Skr0J4uTi7nJ7QwG/BRQ3PM6JSnvY29Fy+sYA3Ns+2CYXl0TkzsQYQg
kZqAZUOqnGlhSB6vkE0cZHBH7U3kVbBY/9pBlev3ZY8B3wIiByHRBLZCiIb3p1eHz5splg8BOyMq
wNgpIGn4IXv6LDjwXVBRbljDW0jAfNJNWxevD+BRge08Bt3mQPdz7EVnpksWEZm3KfeKWWsjO5zb
mi07jg/o3gP6I7FcaNB2+NvP67crVg+NTxVzdOnP6Fd6O2g9tHrQ8+M1Zwq1hAHiIyvDwUfQbIah
cvaS1De4tSxxbuiVX4g7Qx+mf7lFO8rNOK7kOetcGAXIwIuvfjjPoMrV2jqzU0cFT9P5K2gw2bW0
zz/Zt0NxEUyGjyMxjNNXY8qJaONwxJPHLrXiU3Ato0nN3iRUCzSYgLGdCpjsgDpnFOkfFGRBDEXN
STTg6uewj8l/7h+ba48RK4wmvg3eE5Rv8XgoZrJvjbHp9aOivvxBPtDdWWt2Io8lQAjXhmf+nghL
WHliKN650dkYSStDLLwqml8xg1+Ac5DPC9c3l1n2Py/qd6sY1PhYXme84TE4dEogvktjf2tGpOh+
Pw08RIklTTkIyIOBWHtpY6XfIjJqc9P91HUZ8EwNzry7N2cKY9DbKxUCJFDVE/3Gcbzqyxg37uG+
Fs80r5KsGpOUIxY0cOzKAOLdYL22AGRvtEYjXtg132oenEmS2y6qTDQwMxBGXlQZztUhBlcjN1Y8
GpTSgcWHDt3234/fcR/ZGEugh+YipSosuhGMVfuxi9xOhgPMhdA3jJKjFu7IC3Ezs/rNaPnkqLy3
AMP/XcngjPDh4zvBYPpRbQlVdQNaYx9lIOxn6QLy5yBMMgjqL398ZZuKcfTYcfQr97eet+hXY8zH
eThs9VN5gvEJuk6U3gBO6SX0GBQ6PAP7Oo68y8sD3i0j0+5+kWL70ABm19qDc/zCewBU6GpEWQ+o
HJZ8Hz3BZUgMjwkgx3OVYzp+WgTKI+mWEB2NTQ1hhqLNgwFduJ4oPW806arroNhNqOG4DsEoX+Dp
igLonyduLz2brSV6VyEaPnY85JLqlnKGSyU4gwnlrvuI3MflVuYHoIpI5Fo6FR0qUzB+kDqfZSKU
069kwIo45B1CfhopjZZN+ZxhHphcA7dhlOv2Kh4O39/frFAQPffZip35COR/iTdfNDBlpigWF5gV
Y0qyB5ezC+Aq8QX5s2FJjfHgSGwusDKo3AVWvGlAoOrrj6pvQ63h81gkfkmBgj3VgJCNjZtOdoI8
Iv+4lT1e5OOocFlcNnHIDGQnAeAFgzyhQceNsuf8fzXN6zzNq42sT1TBeqoApURpFWit0DCYFg86
RrnhXWXSQv3XUYS7EhJAXSm2A2RLbwEWl+JXqH7ghcUOwqoCD7xb91WlpGM2KMZP+8tobSDGLr0q
Edrm2IL443mwIn80jvYrPSun4Cx5OUfPi0lK1msNr5dwpy+B/IR29IrwiyLYtFVzpb95OIG/Qd+p
0UjPFuBS5wpEwKw13fFUDXLrxzucWX8kCEBxcsz+lYo0b9NqDSOtn2zSqD8dBPIb07ssLCykq+T7
sjjL+jnrosOLlLuXdCwGNYOP6qTv5OviPip7UQ8G8+erEaFyEKuEuUt1/PTi/Q1bmkNIq6rP3oKg
v53ZR8fJDKaidW1fPR0vB9NokIf2knRfL32nfu/HC3lZ9I4QkVaPqaTEwmd6kdpNaymS+bzXD/DM
v/GcbNgeOz9NGTjBAQtjM95FJJ2oFvR2BcJqiKNgkem3stijSdnbSLeYAdqaTHDRhkB4NEIPOSwG
QleyCxNAT1wHjYrjQK6GoFmlbf+cJgEbxU7Z6SihCaLhmdHbz/z5MDUpAwQ8hgiEv0CipRZPLJYg
vRKsKh/WmxPvP60yP6HTkLhMU0vI+z07U/rSBx4pM7fJVnDHEiYHP1COap3zElLdGwaN1G2kagI4
jS7dNEBBNM2IH4P6N1/E7clDA+rRT2mPX95isF2DFF1/wWHIFeHINxfA9yQ1yM770UcW6Dq67gZz
wSYpUUB6wvP0b2UCsoIfzledZHnyMChZ2R6gWpunn6KHmno+zgmvGC/UpY5aEtCDnUYFqqMF3pZE
3olFAdQw+UOsmOK0WcIrjmgCRvZAKiKEUvoQGGTqW2pce/ubx00mIbMLWGcUqb8CyDVsFa+GBF6i
/ehm91otZ4XB0DpbaNy+swnOVlueQXeECJdXmRSJReVFwUhMLDSxA3AJ8EkW+2gbrW/in/vWr5yP
QLJH/voz29ggfyjvH7h51oU8D7fazbfqnXrsTzWyFWpxCSEM7PulUWEQ4x+bW/LMskfcgSEpyrS4
Ug0MkLETXDtwgDWGJh3aN6rRKGoBilQdXpqq8pEou7jsp1otEcmXQDR7u6mYYXK1DfS0qJh7MGEV
j5GWcjq5jwfeAViq/K0ikxcKEmXLp1iqqG+88PHEJE0igui+QbDpHeOjHhn+XR4Z3dcrLuejxrhW
A6wCtuTXIOurxpCWr/u5ePg9jcPR/HON6wscu8ndi9cSn9Y6YMD9HcNth+b2qIuBPkG7V2saOH50
2CyG6Gi97lAxnZMEQHV612XrwEA2n5CUrXYpJR+stayel2+TgMuGcCCq0iCobXhN9aqThtY3UHXd
WODUMGWn5hb6uhcoXc2sue8G+vBGuQ6NBvdgHKMK5iSgVUo1lVukl1YMjN4SH2f6AJFJ99UpUJ0P
BtCJFXnS5UebTqEo5lj/igfc/wEZytPtkx9o4UyUAeolsHbGzQZeLJ83C0Aq7Ew4dgX4QWUH4wWp
FavePUy6uO1QYaEOOXV1JpJSbTb1Bq918wuLg750ug1Ipkcy+pwSyONtv/lI0SDiCUqmArJKx2U2
oSHst1z/M1HXiEZVY9ieUOYJTtEHKx3qeRQ1mEChiP5KUKpPNFfGh30Ai5vYwnDyXI7JPx0WfS/B
YhCLeznaHCe+LpqoPul2b1v9b58jG2IFy3ljVSbOOWGQXijCUWZzneYRvCRNG4k6OMgIBKsXyAI9
7jMUdH2uqGS1mzxpe3iUB8GyQeSqD+SiSNj+roC+9BAj1Et4Yj3qidB4k4c5cZ3a1GlwX0orYrXw
vn8XYq92Yf8V9xhLgzCWZQtBz3hZrd5J9k7IYPp/TAFlRU2gm5nptKgDi3u+VM69Cmk5ya9tQ7Ct
hCspRG5VnEiIb1ZcG8700jvhCqDl03KQbz33f1oX44IaVPasjqaMpNABLo26bTx3xukqj5ZH3hYd
LLLMbf+c6MKENImMNKN/EfjizhdKaJn0qZL2sdVSIvDf/szG8UsS54OvRhckZEgy813XgTzDBEse
cfY4wBIR4c6VLEuRl0IybjVqgmo08uIcNu4L3JrD3oWWZXhsCEY6PXabiA26+tsXnZGdja0m/64F
aShfTYVdBapSZzaZ66tl2Y0HAJ+IdC/Umh/xhYRRz14Ik1zVBoPOhaLPyZED8n1wwiDhmx0fYca5
TUCa9uWQt19XtLQ0p27mPsdiguxcw/HojtfJTO8FrhyzgyJmr0yTx9A8CJ8bt90yyIh0k2yLl+p2
tjCFB7UDhI2y3lq03wwqOI7nfpGsk5pkz6bflllOG8aSg6LYRBnpY+0yh8uW6krOW8rpjSKT98XE
2Zi1tZxUMPhG7s1hxPF9xp0013WoubOMwOGz5j9RXuqJCxZtkU+z/Zene4fCuhgk6Bsvc6Tio678
E7zavmzuSzAny9l6fDUcrGdAVDA+eH4J8YIwWS0JVvOB3L6X6tqM17/uN2umYHzRmz1fngFQX4jG
ibVjqIVvVMEy9lEgzsEfKMTPkv9w1+KRrqHRf1P3z49cfmD+I2vf2GsBAiOBmjimRkq6zvF8GbXj
yw4GfqQgyzHuxFAiOTzY0QJZnd98PX8jr+3+YCscMgHqyscBdoypGdhYy519ykJiH/m9qeNCNbCP
3QMWJADrKSW0facd0M9XvG9QoFPS37nYVWq0fRzuCcwecvpm2yZ+YO9jECqVC1kOhmoe72YNUNLz
uQ5ntBvmf690pkZtOzZXSPG4CkNPh8wCJvkdD9Io7ZvFIIGvSkgDkGkTuMPEKGZS+uKHT43jTfue
u2gsPG7zX+S/DJWGOnZdealsxaL8gVkUh2Yk+jlcm0BcGu+TbCYxPRWmEH61z986aieiq6K/2pmf
PVQ1+yPsSEoaeNNnLDQfXD/+hRjUVIdOCvq+zuyVMj7mH+BtjhAMNQ9FT6YUABqRpdn3Gog+RV2d
djZgE7f6Gg==
`protect end_protected
