`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Uo4XI7gfoX47J0/hroCNwXP9HZ8igMyR9xSuAtzSqgAzr1UPTbpRWGnsgC6HEjM48hN1tWyHDDUM
e4w2fpVbntmAUE+0l9eFJVhVjHm0yzsqv2Ugz/NG7YmgMVoSeQo8atdxsP4ZgYuRUt5xm90YJ/rp
2ahxK1xuyIyzJv/c1CnjERe4m9LQJQ4Mv62JJPnTyze8BHCapAUPJnx+UUoxlUqQIQS6S0aMABep
SwmV17sZMQYTVTfuSqthWN1KEt6Xr1PCrSi3LVEyvId2C21hmbX2tsdFMvToJpEeKnenwCSDJw9f
RNjshJBbhOV8PyZlDewp+2G5nFQ0R5yDLhROZQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="2bUKrXbKiU3qw6lveff9MyW5hL21sPk0nJxbhQw2RKk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8736)
`protect data_block
CkqvSng6rfCgzx3/kpkbxDtASLvmEM3BtCGejGJnAAjCz+0nqrTi2QbiFwdiA1tKqc2MbhfKey0M
9IDpmi+vqhL683U5nwkiIgszZnuaVwOOr2+kAHWJaFDmoQ1gfczZ35tPjfKFLQIc1fJY7dhKLH6w
dgoUQJ0B3M2RA9URK23hJfMTgUxIxg0XgQXsiGpEJNH0J33Nvf5wU+RSnxgPpaCsfJcQrE4NQ5SW
OI2vXMBpz3uW6IlrkzlrqOcNg2vekjm075l15eHxPAefO0UidyPIRgGbjzoqfuxc4v5r/bA4rbKm
vND/p47zbAB3GF0TeqoXFnT7+lzlGTYwLLWGvIoD/Vi2sBvAHBEGsMgHBZFonxyhBpt3lW+fSB5l
4EKSezTv+xsu6vFP5L+mzHACS7G4nJ8JNWHa1EH1r2+qQaAfPkKf6nEtX6fCqPVKr5oOEqNzGTKu
4F85uPDaO3n4hn3CS+o6k076h0rJCtTbUxPL3V6msPVPBkkYUM0RwurI81P6KpbrOhiKoO5H5jsg
IE5G0MUixFnGa17jIt9wfPmrMG1AAiLn1wn71E7EHhZlEBGhUH0IPykOh8yHF8nkrjtpf5YDTG2h
ubXWqZ2IlETJ4VvGOKRBq5HRYw8JiCFL8GFs/Qp/O3tN1PHGLoVYCBIUmEeeyyDBVMuZDNe93RxQ
qkuKuvooUfhpIqV1/SBaL6KQn88pxxVFzNZvmuwrQRo1zMzW7z464rjhfkhdWc7p+iJ/kl8mwwdt
/OetXp88wxfEzhDxFfJRtGCEUSAgXRKBwh9euazHyG97wna8aTjMk+8fxTOyyAlvAnFipIdOmNf0
vXlPFbnSiHSDPM7OZjgZb1orDVDpkkCXlfts8ds6A4ju6Qk4LRE0PvzWQRS6LznCHzhqMIGPxIPg
az/AknVpdVST4WqVPQp6YJDUL6ye4D1EWADB626pW6iB7F7wjJPy2IagLKVl7JfmS5W3g/lhLk88
rmvp+4Jl2IxLsJJXCyaeVD7rsKH5zs23wphfJlDh/VxnzZQYA9IWoIKV/mFVoMlE9X9mcuVJi53K
dFqseOZXDna/s7H/0KO225fz+MQWkfyqyhbkKHfEElMmNE020I+yN78dm/slpXoxwx3yO+w/WmFm
NWH3yZPYgIWUSnQovlvgBC5McpTd0Ri8f6X63aYzxjnKjL7/GKJ0v3y/JbS2BQcT0VPZ7h7DxIcd
68glIqspuDfg0GEAVv9DyHVdbIpTx0vXFhgHsSiC/CUX2n0By4wxIMpnWGXw+UyqkYYVF5YdInWX
J60DYpBuniJvMCBXYoRk/R3u/icCeKX9bJxISakppSQy4CYzlNtJ+iNWQcYo7uWvRWGWYcfspV3I
TOcuoU/UcuxuyFt5qhRWpIXP/4gC/0rSQ8U0nazEEIyBbJkKo4YMjsggmHHBGp8+vl5NT9wF+0qY
PlkLucV8jgknbm1IIujvQxjuLBZiueEwpkP4IrCw+AJhDNyudbMoDAvNZjfJn55bVbk7TvfjxCMb
4HaoNjCdTn0LzuztJZOkZRwr+4QdbdGUsSf+LqH0dOAcpaxF7mB2tYpESBtRLKt0Ae4YRPFFbFDe
fMqAZu3plMOYBLjc89RJxpdHsPmvEg8xtrHkSfa3Ckz4JdoqOBhoZAiZOcfLatszQwuFyVUADlRf
GfvR56MN929Bhl9yAT+/18GqWGXcx7KDGD5voc+58CAbNUKXOlJl0ewcUqtXCiAmvKSPwqKjNGuc
F2D4nRRkuBU8Ed94IkauPY9VdMJruREtjNUtpDbSTba+hoe1UCYvxZjxFAM4G3tZ8EvNPDpeYvbw
H1KLXmVGUmGvLqmSNQlQLxP2byGNdJ9QJHezbMmPglPyq3RxvCUSriJT5HVJFbR/rnC1Zbj8lfPz
G/KZtH23gE1o7HwIBJClEKSBaOgPeVXhEaqetbSPZKbP2vbS0G3b8zCsKxnfh/VL1zRaV9cSF6to
pVIpViqNKnkKcws6WcrpmSAR4WUHRXqxRj37y53wJwQctDqT2fgpLyrrNdUfGGzi2r0sVygoK7ZM
YhgiKzq+CtNUaXXw+CRBpKJp+t4Ppju7ayhnTWdm6pfKIrDSFdKH7l/++IkafzNTO/n+kyjhDiBh
TljkqBRNq6p4Ho/MFtkFrIrkBGYM6B8JAcqvKun8uDL3BBm0JXRnKIsYe+TZ1ywo4Hp4J3hbS0+0
NYiPSDylbRxgS9hvja+re2I5yM7LMloEiic5craO+4uquB44zIMvqap1Tyzws2uj2GukJ5yk+xQe
RmOt5NPEITBpyBgxUwHwgfPVLpQL9mNb39nitmmZZTD3fTw+Gei33XLRBHzbMbyFHkFtiK+/HOhU
NrfPa2ES3H6w1B2mkS2AGT8ezLMOj+Oyv6acAG0RFVV20bfqGRE8m902XsE4LtVSA/UND/d09RQA
vaQtJXJ/jpzXp+7W8/YIXnJrmHc51Tc2UVtdTCUrpi1KzPuLXgyGfgEYDHi0Gt1V/6nmy+tqp/Hx
mkaYXMPxiM5debVcuhG8L4HwcMABy4uP79htArHsJ5fbsoI8mJGbzSJT/hfxorUmIsnST6i6L2hw
a2GGAX0QKJH+MPrDo1Qcgs32sCqlIDEXqxfCxjTspe9/0EONWqyn7yecbUsM+FgmjHtgLWpwqnCB
RMP4g6HA3VkDiGNEIjXvS+mlVylShl/GNypo0OKct5xtSPjMJsJF/rOd7RXAlckPr7wlZPbt8i4b
tV36UlKqtE0ZQ2C2STbI5yX/CbNOj5A9DwQEhlD9g440vm/hn8zpfwl3L806pkIpvCX3mStK/EPn
V+pJOKoyxfe8yC6o54uAP0QIU8fX4YB78MA5T6TE6NObIuyOQ12MXsUPRE3DOIIPj4XQS89Inams
44noj4Nn+XcawXxab3jKF7Hia/c5+Rwe/r0phFplEQn6n2ZkHg4mFG7nHNFn/wcetFSifJdqnIZR
E25NZqId5+068+cUtcLgU+/WL+mmWxBpNrS3sRJDM3mfcBuO3gujLukETyp1ryA8vOUwdkGgQ8tl
p7IisEV+ulcAXogqhqUjRWavNgvLP3I3YnHUAGslOrCjHBEz3rdRGJQ2rgUuMNEJa+TbwN9VTWRz
OnR1d5QiUwIicQVHCji8kXRdviyLXMlFNNHedg8cUwFU9B53xu+CxnsHB2uF3JelmUbEeBwp9wRs
OPWLXI69BF0MSx7R6nsJlpIbVhUc/WCKlAaGL0jOqfZs9Gltz/B6k8tFSARbDdPCQMJ1LOJObt2b
WXGm3kxTpXMzZBLl2RkVSvCqQgA9zx2n4yz9ogXgLnVkI/oQdM8ctsJEDfVGi3iCGF0vK4f3RiI/
w82bROWjlYUfvzDg5C5v7q227H3FX+KtVzme0xCrtIrRP7Y+NyE7Z+p+Qf/fkqC55kk2SAmfdrl1
Vsfj3X2GsJEHkqtkCJ+ursy9rzu6uZenot9z+nYr0XwW7t5/pMcWdl8PkCW/rHVjYTL8ZwGqdxbw
G0DEDfnO8t9K3KrcBTmVmKLMD4jPuD9AkpVTTSgXY2iCVvqD2C2cCQvJIKRbtnJEQW63fylnLyyn
JVQcwXSyJy5KUkg4ldrYwf2iJ1LWuAxksRSjnDRUskbvwC1HmNlArN/iR/e37hT+al7nNF+pjiRd
AUM7MIfV9K0cBt5wNjFVExuU76lSTKla6caEoISF831TezRRI42ENsBtk+T0yotot+wef9osTP4n
MlNf85+rS/fITKa+K0HAsbfPYGRi3DxQLFTOnVcknSNZUfTSBhcbFuMxEFG2N/VsLU1As0/x3C3I
OEkIo8nEFU8zx+WvmrQX7Ox78yPJCYhZluDaploeZKRGN55GqlF0BKe2YaWn2IrEN4duY0jHE0Hb
uicBmzVGBsPEJ8qymH/Gsz8ciphPAedd+1enyDFVAzBxIHL1QtxEgEEScV7LJpisRRgsUMkq+NPk
O1S4gkU8hIE9cccbBn3V8xQ207hS6ML7mvA6VybTKGN1vbotOheh6/KzkbcJGT97kKsTg+XKhMKG
Yxe2YH1dAUF2ClZqm3zZxRBwdrH5LjkSuqbBklxwxuf1VcYiTjGI5CNbpW2VCxqPEFo+gq4zS0GU
U4tr9mqa+8hC8cbuw+x0D4FuiTvxSOuWmx1thA2gRVDTctff/xIUjXfaJNam6Ony+MVWvGqYv+3n
knfpJ0/0rS+yfEjhboEN1eIBcTviUQ3icsZvglkD3La9a6V6Tn1GDzPWvyqEarsYjkuGrPIHLgX7
F25yFfO0EWhxetqc0Odl3dyfVS7bF8HNEULtWK+rjHJK95x2hHDubkqJmSeqCLndgIfgm16Gqxqb
C684+hPRtrBSB1ebxQ3gul91VynKTKSDptiBhbAG5Uv4z+nhjusRJdOresHfG5g6XFhBFZ5ul5UC
0lXKKdXrCCG065flYfqrYCrS72cweSy8WBWF3TPdc8vv6nRjEfRKZSlmxtjHI/2yfn290sXXlK73
8sSV62hg4AsGEHDsw+6B1ZA6jaOKWonjYVtyoh5+HnbLB7neTACV+OZN5Yp/rW4ojQRFZE+BrqpJ
6nlQ1bnH9bYsxrz5gZKcg23tWyEnxncDKTcg+3t1/yKuYOMga+DkAsp6nMJ1ZBKJ3F/k1UWzKcLX
k53tenk2NoBVn/TKwJG9EcauOiT+6yQGeaG+wk58/YyNm5Xdjp1jSbF8zlZZ11Wg3Myr8l/JPpFo
B/eNO2YBy05yCiJAPYAitKm0Ns7l4rHLQBXxJWClkr9bfC40YYgxpxL7jfsZbksR69tl4+TB30mV
QxZYuL9ZfwtUwV8YI/RdQeySkDvoUJyGlNwV9C8FBxWLCOT25/AHu94iqyJjOIC1899c35IvjWcA
IVaBf5ZIfDZSjEtDSlhNsZApD6fGNybjcPxGyj1TU6jk+fFuYP8X097Sa9LTjweck736y/kbhDaW
zwjx+wSalsb8AmqNabTXyhmOFBRMPXM4i9QH21j7fESaA90c4s1AjO7NOPWIE25JNK0rj8H3shSx
5E7jYMg+ixYd/dq0RH6Bdpm/nBZae4edC62/HC4NPUVKMXFXwT5VyfiZlrEhbYeidNWM6WNBrQCd
5bVaEn0EEx3wyCQIL7EKjKCw/WlNo9z6ycVRKav/cJX+6Kquk68jSKtVsepS4kFxRn8uRDMCIa6a
wGTuMOVDT6hE2ixrbT18oZD0vVwVEj7wJ05+FF/LtBwupjkBuzoSOkFZEZJLYD5t0mHu/YB2tT5I
ULIXlaRTp96pbhPr2Q6zcfufdQ68zfxPgzfDpgI4ANCRznW+mwn7ACwE/wJNqNqV5yjVkbwbh0uJ
rIOIfKU/Hu8ZdMnQY4h+mnPxs1V5QAoM0VSo/K6nubLS1YZ68ZroCFc2BZL0rPf3co5IIk03J338
+Oy2w7bR0j72spSvx+sWTzq6x4gm1owxcYbfHsO5JU5dRW7h9w03iL076r6oEBk38yQ2HV6nq2fJ
EzO9LqcrJiEB2dV1YFM/uOVPfq8gRjxhq+WxTusNKFWsA8T/rc1Ob8PPTjbFGH9zlOXpIc4mlktM
UCMYJcOyMdFeJJq4B/adqwz9TZgMCHRdGBeMOjUpgf5etNvHtP9l9tgemN6PArBxRCD81hrf0FLf
w+LeR+uWlqCZd5bqoihPjf72CxQ/pB8jFT19u8hAlYOyjKcjdOVuP8Y+Wxj7Ce9ZuHRX78AXqtKv
dmp312qsytmruwUPyPMwPLYRGYsmy84A6PiI4RqWedr1y1fOmCPzA2bS2bToLPp+GhXM/vuTUSDH
lUBZqACK/s3cuCc75SZBjCE1qqN76Z+kFLy9aXnT5P+uu9WqN9AWWSFrmOz5SQxuw6D9OWgTB3sT
TpYDHm3PbHHGhlw+16RvsHn0yiijvGM7kdzsMNdJZu739y1gXwMZVbUj2VU/mgEQ4fWubOdsS+/U
IjMhMlv8lDwA5KCNxHB07RjD1YSkkxXQ+lF6ge5PSeIOyEXU7UWKzh0o041gumhIMuv3C6ZKlIb+
AsG5t6QqF9Pm2umcrlcCZOH7wdDx6r3TjQ9wmznWfDr9SqdsYYK6dvEnRuKUpcfGn1Os44TWob8E
lfIRK5qlPoZfczz78ilS1+8+V8ifvtZqf2pS4HnJeRsjTmq1UjV5WvJ31T/EHRKbjChM32MyiD+v
99HjRMrvYZvOaeNaJphF8Jz2Cox8j3aRJHFz8H2/qHnRbdCB4Mgptk6oKCcSR+A/Fv41vv5kmhNd
B5fGHRopbfAgjF1MZQO8RewbR/W0ZZCOfI5V8+m4Qh5ANI4qg8FolV+W5N1LCu44iew9y5IuWtId
/wwVUgVkiZa5a2lYj84CprmFngtJE8V7DyQpEGuKT3tC0GwNMwH9iao/YPy+GEMTKICcUH8QxFks
7utJ8iWHOQDL9oov9KTS+GFVh4SzFdWpr0/OIWERx0yGNzmVZsb0Dw49J6FRp2PH4BQKGPqe3LTE
tXdmGBbJ8Uz1/v1sVQijXUd8+9Viu450D8HN/+frd9rC6Wk0zToBzeQjOPCe8kUt+8E3+tEqMM5i
/vEUU968+QseMGDnTIobjdMf49dlJFPP7Adui4Q0iEk2WGYFSW/cSPbPL+yfb+PnRq8VV898wNfZ
kYnyLMMS4lWFze0xPzH1IegavqCy1lcTTE9AKzMur1DDPNk+9s+wAb9QIoLeCspupoqirHzcXD66
5HS56PzNc3eAnrp0/nZWEUDg5mLxq7nxlPwStwExyLANAR1xQ+LH8GP1y0g8HunmYx+w6+dmIuFf
9nklG4qjTM5jTQNf5lU7255uTKkPBWDqvoh4fSc5ta7DfSFgmVmXPjqqhVKE11AOJnFOo+FofiMM
Yk2lC0dbovJG+BGUpEHDDO83SIzRhavHAM5yhCJ2rfZqOJOmvnhH6Y3fMKZPAiRA+WJWuH0gL8Cl
CWrb+ZikcswxMNRYzst5mjnIkqJdaenhtux7n+gNe98h02YqSKNxfJmmP0WQ0RPDPaOheMlQCtDx
yTiDgNY2QQVS6oxlucJgcbaruUBEBJamzPfktuHkRIXvogi2Gmes/v3Xjienk0mQgsnsHaO31T0v
UzaU9ChASOX2EW/JJUkzID2rgoPz+5efPiA18Ae7slAGJZRhuaUJp68CIN3tMiz3+3j4BLxImSC/
vL5daUB9ZBPRNghLqYmn+77stimTTzt8cqHf4op6gatF7MMuejlzLlRGgkdzPkCfLtY+oKmFLD+G
p1GaTztAHHe24edGObHZMS4Juej6t7P1OXQG35RFw0UeH8yI0vpCb2WkqOvAG2R6thu3aIIYweEX
HtNS1cz6uPLnZI2cHmHmT5GXVzexTVF2UdrsdqHmpWbVJnwergAhlR1VCXJiIlKIhCm7CZmg/2HF
yMROmFqC8bFncBOLkijlwVITzL8wT0fBcmTOLHvfzv8kSXdQm9gDXxJ1QjdI5Fjgec0xdrX7vs7M
9A9ZZpZyOyNKdAmE7va1iqfo6RRA/2gHEnjhxSrfSB3u1MnxjUwBr8ZKyj/u53xcpZWWuLnlOSZ/
ICvlV7pHOcCWYEdTJ+pF+j2CuaOuRR5iGSDsKdt++rawyo21LnCbIIdMCYNSqbeFfPmoQeIX209H
gui2PHJJ3lcKZOUYL+YdDRGNlZMXsbCofb7lS96LTw+ApMusPZ99IyM/QfyNh8bDa9GWQLE6MtLA
6qQsuSpcu8IDc/A0E3CNpXes1jqzhaRCvRpb/bpx/Sin6WVUGMXY6TiWzhSiRCHX+u9iZr7IBcjl
yRL/zmKt2oz74PBfun++3HeWgjVeYFchxT5J5BW2ym8SFoHv9XoKMYn+WyLLpIeu2a0olc/6dOtb
0wXbr7uOOzM0jJJdfa4qQBNsSq90bRTJwe0FZ/+OVLartijQUmmKXZBSFWJPINV2VsAZV8yJr+Z0
sBx6AGcKVy+A7Odw26YA29Ed1tPEy6h2ipXV+V76XDe7J8NRNfbP7dyCMkLcc9O3q7dVOky+IY+2
dL6PQq6EkY36kc5MDEpd3+vBOa8TFlrQhmbJU8Sig72UL9qZmCVMCQ/YHCno6tl7tpyv5R4/dkp+
wnmUNcbLUWyOTm+SxEXXs+PuFw2aKOcdHHjIYlnygkdltisq6yDmZNu0JZkvfT7itRlR436lA9XL
7aZGr91LgRxt6atYLY8EnQ9xZdrgr6Pf6hdQynz8oX06dsKgEImjS/mWKZciZ6ZFPCN6pEZ3cpD3
PDqoGrNzwdb1PmZsjRy2dtku1EBhMjQUy4SqkOegNNir7Q/xZTV2BvCF/CyuW0J2Lx2h9T63LryH
1eZQawRgA0o6NnrFgxv5UDX1X+tuxJ6cU9VfDkf5wzyYHS6bBUxI8Jvf/0hvrZWWA33ROPogj9mc
og+Qz59DcdzQLMMlC5b3veIUIQbO0qY+kqcbtudIF0490/5hXuQKKGpIsFjUxFSVFSyASb+uDKHd
b2QKCw8b35IPt8ibFBVei10meIL7rPxVDR4Rzlv/1tLbrWOkE/7XiZCnsDa7JvWsygv4VX0ncy13
5qk1z+oPggc2fCm+iDMNQne2pk3oLHCLSHrWS7XCK9xM7Gfb04UOXNG7oyuobca+Y0fy7t5uRyS6
2aIZYwJthkRBHQug0Wfy02SWiGXalWzrMaW4m+UrGOCPtDntxXgKBBQ1ewaFS2xLKH70hufyOEg1
xH3lk+vNxZESY+CUTwAA8eGGdMYbkgSpOSs+gxOUJGXHd9I/2g6ZPBfOYdT66tw9/pJmJ1x0zzjB
I5ldWEj76oTc73y4CqHGnszk6uF+HE7fZsu/1r/gxjxh9pKtfmoG4Uvn2pNpFsWUl8JeCMTFBNsH
D3VnQWt4pI6yNOJiOmJfn1hVuUpxtcVXi82/rVer7BpsvKPRz4nCFzdyfuXNNYscz23OcWIIXFGM
m+Irk6LNOO5ykiUbRFLNreBaYd3WkPULjKuOF252b9h+IF0CFWbnvZEqtvn7qox+VwGTsLhBpf2O
pmKw9+vWb4hB1tH1OHtHZxbqzJcQwG6OJuuPpntAfny4FiaZj6CxT08Jw+2NAiqM1dv8OWZ9xrsW
V6BFehC4163iInOL5rlFs6z/nOIC1AMyg9xNg3qNUJR1+BXo3AaB5p8xDW9vHL4+wPu9miFLgn0u
T2vstR815k5VoS7Fy0MiKvo032ddK21QI8yjjkbYbEsdgYkwWmVD322hJZW4fW5vGzEn2smEXobw
aFbkGytwIRGXypCWvxY0P7FU7lceP1aGEhRdH2N9yiLJLVochdFPmvwR7zqHMmYjqc+h00OZkIvo
pznwX4nMQJeBCEyFtJivG3ft1+wJcgh/0xWfaDlnOEslXdJFCvAR4TtAWOmc2QTiiXGkiKQvSiyg
S8C09Ny9blv9n/jaHOf5sbbfKqjkrHd9vzzotNi7VPPHASYET77nttkwzLho4W5HG2ADgUHHnYwu
/Y9E5vEVcisdDlA7yCnRBdW8I971/8Y2/XpKj6Q46khS9mGcVe1rr98mcxKT5rUFnfjfWufkKpL7
QmlGWBZMliJdBXR7W4gXHTv0qK5qID7QYudpNbPHSM3R+CygpPD9pdwyaGD42fdxSr7TXyoNEVci
Tt1C4OycCtlIIn9Z4sg06GCgB8oNODXURoRMuWMqleCBqicMku6EecqnTBluwclAtxOITh8fLiA1
t5ESNLVoTtwGiJWDtTrwykXZpC6/3sVsNCB71Ah3D1Fp1vLZKkYzCgElaYI3RyFzaVkXrtyexdQq
pBfErxfyvZsXkPMuijxclfQx63Bxq4YtnNUbOnAEi8q71wz/4SBEHF5pAG0bdlEtIh4ErqZnDk/u
d8mH/k2qMXtN+hHTmxCdlRV1i8trTjy20Jwo5XmwOpT6RicpmiRY4KX4Xzf7HnBrnFu3ufwqOCvE
t4KWo3vZNtRN6g2M0UaGDciXAW5JuM3ZctryWTimAdgJZkV6PDumt4S2FFhdh1eCc//K6e8U5b42
pJLkiN3fCEfahnFqLLOhpTwSmWeltXfmc5ZDyNG/MVQJbJcCQDC98IwUMphriKaazqpYrrZvsSc8
0bdARpGxdMeHrS/P2k31zMqogFMwZS/24ZC41CvOrK+uqaO66NP0tnDj3tvyCqlXD2UoaZ8H9zLF
59JoDd9BiixDzYSTpaoGP1XUetSxFTGTVlIcvHMnxPqUk0+BV4JGVxFJMm8Q4CYiEaP1V4UmWp34
OtLoXmvBZITVCAdYjJx41Gp9PEVS4atM0oMRWLT0s/9E31S/+dJYRyrYuFp21h0sCBpjONr6pf7T
rkiKxMgdyCeOvf2CSNlV7xr/Kqqtg7U8by39Vw9KGV8NmMIaYujDmnxypxZe65YkUA/5eZeDp44+
9PAaUv8dUIncKL1mhS8KrBSi4uxq4HMomZ1Sxpe5GDdt5hoFT0oD5FKPUCdF1EBZoIA+PaX6faKc
fdD9wd3yat+Ep5brSO+/N9p3zZoEPXfJC4RBlb8ynsiF1A6aNdWbFylVSXdUKnYuxYs5PFPkfIcA
G7i3iopPJEk7BaENIhMQbo8GYQhAap0CQOaGq471I1PwvZPTAAJ3dDHAQ8BYA188PzxVKzr4dz0r
UrUWY5VRyk1Oml5HV7iPn38tE8I+yGXqTJ81rrN9+Td3PlBIDsni7LXdg16LcYTuBT7SCRu+J+tF
knjDRYY4LhWMHzSCmZNwRPQeigKB1n6wWO5M5sFE0KqvDXKCTQr8TxDNn9zVq50wiPdz1lBY8ntk
Ls3rHQB5/WpImvn9RSy2vqnUTC17oyWCeGXlKjh/aGWPGYZO6cbAO6nXuMbhI94GbKloKfVKI576
JF3L3k3HtJI4yyBfW5cOK7penDnYtKzvdeKfHaXLqDfmIwRIhp3MlcfpkkiCzkZSGjWVZrN7fG4P
kIFso2Dwq748fWxvOfolz456ITphp1IQscAPjEeCSOAjMLkdgVuiqXOClOoRHyKciUDOKIFWLWWD
7aass5zEwK2pEE2nVmgP+nd0Ur98G5OMAuSL5xjI56cOIBqalPkL/Ic3KzzBIJGxU9Pv8FpUAVXl
4tSE/vmwPzu+yH/Uh/45hx1tYySMCmVHdzPdWTrzOtegAi0gjay5vODp/WivgE5LBXFnBmSmhhn/
CYU1CoXw3yDzPlafb+mBW3w8oUE5P5pidVlFR/2zy2IcZQ4ieXUq7PGW3boyYaizTafDuAWMjw7g
WiFVCw/cD9eN7scYregKuubKnSVwUi7olFgAxrutyLqfJ5++CG/igCke7z3UgRIyig5s7FW36NqA
n560O+Y4iQVyuPriNo4hUKAA1UyPorRTBi9DlCGTCAPJhM9XtdrHPCWRPV1Eml1C6q0idaYxtlqc
w6OkFQN4VRrqWqQPAxJ3waS6IlwRQZt5WzCHF1+N7FZp1ofVHYllfXcZ59Db5Lc+pI+FqICZqRo3
bWpoHYl3VT/v+DxHBv2Vm+lzJL7jtNsXObUITA8ms1vcyidxb92xUODDc8ZRAmwT9KXH8AYb5OQ8
7T+/ZNgS32dq39jnqcn3YxH0hK5gccI/jUrxC6iRz4xNyGupxruTm1kHQC3GNv+XGeB8Bv3ud4t8
luYpptZUld2lfNZEzUyBGo188UqaSgI3A3vq/i0ztfz/2fd1g0x5U4RWeLq29vN7V8bLwVK0zGaE
A3rJFKCA+Gm6cLEO0NnY
`protect end_protected
