`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
S9v1AwiACeqQjEWmlz8uPEM1o4uf1RKV1xvw9NNo+TG5SczBxDct3GTuQ3XdsMejfNaVF1pY/Q41
SxOci3jbsQJhm5l8QkmHIH0RQUcOcNpmUwXuX0Lkcv4l+fcFUEgV/10Ib1+flVntcHz5piEF3AFm
X4woqntXwSlMEp6QF8Dr4ot83933gAQ3BHpvv7PTG16oY7VnvWAP6RvPmQ3HSdet/wleIlBPlfEe
NoQ0KAPAJa72Qruxg6Z9miwMrltSfVFDWj/xyxcjzG93Jz3RXjX+K6rC162u3tyPj9mG8gF8cwbB
ZgNbtgl0LlOox72Kh50JqzGxgUcoEAxQX67v2g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="lU+1T91ZwdhR+xHRFwfOCtaiNvVm3gH6lTe5EoiXXvI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17696)
`protect data_block
+nLsMtorisGLmQNGHdDbARstfXNhqe4hu5cGxl2khl/ovRolX2xC800db1mvJx6okIsgEQ7brRt1
3SgFskRnz4RhM5voBcSgJ75PHl8M4qIRluzm9VDrnoNz136fU9sIShuXKSDVb/iDsbg1+zFI42hc
83jl4/hi7AmNIfNnj1UgLzSRj7I76tp9yZs8zRTkyTtpP8b3sspi9RqDQQ0sYhv0KLqUeCv8GDa4
fMGte/zJMsXkDUJu0yvZtK/LltPU3nbubS7j+eNFZk+V7ARGgeF3i7yVvW8RYemg1UFN5AMX/q5L
/0YWlarwzwZ9E2GWjqgWoq++903nkU1UK5ADU86nyWbDrYB2EkY6VSBcId/GuCiVE1sEhY1cjmqU
hLuK98QfzMKiVpS20E4/RVm/25OsWVHfFZNml8PdEQj19luprQ22WxDSo0fKpJG/Qu+DdQHx2Kkr
BDRngk31StqKpwMC8PuUB4pMGgbU5nVsAKlxpivAP17zbbUij80KyNl49+Q9+kA8wrVpy6Wl81fD
JM5OBbhvRcfvXodZnlLH0wkOtZvIfAZwSOuHOqEX8fcre55QnLoO7Tbgh+AeOS2GHvFd4wuM3cnl
A+fjl9esCVE3qpiBMuwELFU1BOkLjxYWo7GOVgMhdv6M4XzKPnrap2ccq8Gcbz06rd1LmPC5mxdq
6BzLyj1th6eU2UdxlbnXFLqMCfMv2vqRToTzmKs1e6m5o4qvLUvq7d/WfSRHabbsleKqAxZbmJCN
f4qXF+A5axUFpuAyUf77uxWie1zKO0Fy2uLUmW3d7rufE4PJ0u2Md/7Fbhb/wRoS2ZmjIZGl77Mt
y4EnbUxn3CBpGNzVSlN3DAZ6L8Z2a8qOcRtckz+1QVtN+dX/b4gHlqOuyxVLzLIA6nefnePtbdxv
XY7/A3dy9eE164QUjmQZmrq6VTDFFPaMBELM7/M5UAkZgKfhHwRzlj34qKeDuBz2J5eJNIGSMcKE
L+h0RilgpYi0tyVAF3CjYoeuP07ss80cKcR+LZ5M/FGtG2ZDqMbhkY7p+Rnc1rWACqnd0i+nGomR
+ZQoDYyeaE6MM+/i0vzcUzkmy7zZWDUaZr87eGXmP9agb/aE1Wn/ZGBSQ8bfnOY81Twf1QiJ7/kU
GzSa+x0McG4G3yjaUOZFMXSQEbHWmAnbjtOhs/kkyku3QqC1E8Yvo9ocR0xd4MLe5+AmuUrhI7e2
yu/bITa/BkYXEnZsTjDj2T2obr7FztqYUW2s95lUqXk2svp5eKN7DZdwwj+OFNkryvc37Y43sOLR
lGBSW4g9e61dN3YMxK+FNtO85dlyXLa7nJ1SwTnlJSEoaD4AP8O6AeMjTfW8gjK5oM1BZvCWs9Qo
H7Y3gdHqD4JpaJdHFmahcVzA7kzJSxF1lp5E+Tcsh1xV54R6Tp42mR9sbEJIPGofsoNynp9gyG13
iETZ9aYE3IZR1N+029T0FUKkjal7BifF1mLLjlfJIH88pVeCjXren/Sl8N2pVgo6TK7VrnJyji/I
vIXncsR4GAS33YYJ8njBVc5f6Ff68xkueTnUBHp8R/YhwY0L/fQFgnPuzEzX4aIPfqZk4zWZBByD
fM1CH9ILuIIEd1dlQBc/YevfsKXXG4wL+YEZvg5RqtTStzZnsIdutc8igk0vbk3p2JmTJohOo2bp
cnxqpcxZgl6c6ot/G2q5NAhy7ZtVk9dOqUcRIlHZcwn1kILWD8amFTxISog8Bg9Czgb9p4H4a+ZY
hwCwecNrOjZU/c8nuGnmiZTD7PoP+mfyHqS/L4Yfr4AcMcWJrJ6MM1ZilO469L76NXcYzDD2T1MQ
LzF0QsHqtPkPV9x5k6VPaEqVjqNjdnPnUobOZfWEOvHSNtWt3xq7WojzZxPFqigGBBfrOLgqRmz5
jxhSkhT+GaMMROnCXrKh0Rc1jO4IFVqqh1FcYoaamlaXMEjlQb7Fc95+1eUBJ5FTeyWqiVi3SvPa
4GqQNj/UlHDtY9NiAYvS96KrLm0dhBVnoGfrCh11gWoRyr1oBEpJXfUXq/BgysZL4jZlb/tai99u
+tgjDgU/nJZwPcwUDvhkC5fc1Y9gD5gTlCfBid2CiEpiwpEMBuyUplS1pkAuf9FjiwA0sSclRI2J
LGhRrTZF2Nfc+DZnnG+8nPjnKaBe8Gi8jn80E8DPDs6jhIgD8wMoSWNljMP3P7SqaMt2PIXN384H
9X5NW+Bh6sU5bkiAPRbwxeUxrWJKKwiWBj3L/FJUs1Ja9P0XcCROmlNFcueRgokrhLqMiwTAQy4c
sBGuXdm9Fl+ZrH6usQsuIWCeGulhN5Yeyj1f9hn6EO0cvk7M+sqPgN8Tb0KzXbMt+yg8oGFGWB/4
cB3hGz0G5c0BizznL4Qb70OOv3vUgP/1MP3TPMba2JwyTUzRfeC7wt4ZLMv8w2Jy8xZ7+/RF5N0x
QaLpRpSchGdqQeNzae8VXgahS36wmVcb8GxYs28fhwzP9YhHdYbqWmT1uYJaTyOsFWV54YOEd7bN
3m24YPpSibsQ0o2uW9hs/eENPqbrEw7HFu/17ZI0TsL7nLyDdb0X8kp6dCxw8KuIS5oKPgCENr8z
Pxt8zMv3TffBokwqIvGF4Dx0gSuwijPGcWXPPw/MLwIS966ORRmAcPoevWZhO3bxjCVpHOD3SP2t
s5JNQjNKlD5vLZ3hSf2pEW/0MSadmlw8joY615y0b7e5x0LJ1r5mETqDGFp1GrMzNMyHaG+a17/Q
1Q3GCIYU8aObmCiTQ/tzfM6IvphLTQGimSGUA8A5d5ZHDp+ZCBIGglH06czFCbmSe0OWSGl/N6h6
+YoprFiAFHw8pHsoRwrk8AaWnAYSEFtRs0Z4Uii8QqJTuofPek6KvzdXmDUo6dsgwdsbTA89xEsF
jmfBa/x2KGXxBmAhSQT/J8xO0nRUEeyxx5lkRoGq46uJD5P8/miV1NZMv4nXosSEO5xYxbXq7m4e
NC4oRnLwBmlrXfxpyMP3meMKxWMJMOtN8nD4PSRC1J2+uL8FU0DHvHf8T2Vr149pC7WEyRsSGmJE
obDItGOAL5A0ViIhMr7TbP6JXqAC37ikdFghhLaq5Xkdz2zxcHVbUPKHb2iWbSbnILjXfNU/Cj6z
ZYH5LI62uvcqKb5VRJNYczJJ4y2i5ogsK+dvsR6NJxI5e7PKKfdf0YVgVoiLLRZEcfq6BoD9434r
EjERSRkqfz+6ub3vvFzt6VM7BrODX/o1RK3rL+hZHVqpOmQUzRhQNsQvcVdVg2VDVi1fWvbzocx3
IlKjH2sEhFQ4MevifLaywH+01TrX8aqjJcjqsWkfA73scjDcu9oLSy6L6JBDNTTeDHozkVX3XY1e
uw0zLFqG2Ur+unCye4VUosM/qe9nGHP+yqiDdOvoM9veNncgYEicIAhuJPHraeXbTHgaAZvdOBE4
zYkzCnpoD9R+Yyd4VSr7aBFIoggsP6HRSDJq8F0R5PGrjFtXtDymKESqDPCA/cqAg90GTiQuBxfU
ji8jlVyADwlfEDTtFceTicZIe+ajKCN2Yg2EEbx54LApua6GhVf6E+rNAtTlw++iLEdRF1S+khw4
Jdxb0OlhR8vMyiI9gDkmAogHYInkLGSmtG3fX31CYk0SXlx5ib0w+MM3837f9Dck+JC+kODrP1TK
5MhH2LDjKjaIx7Qcxt7eB3dEDZX3Lm1oeRGW07GO5+LdQHguuxGrmBDs7hryFekPp9Il0HANU3WM
i4KRqCaVLYU3sHEXYgn8G1ZZu9UFgO/mTEM57iKzErfRcUeInFONyaP1cE3c+EM8w7QYaD9A8aMo
gND9y4i2H1ttxX8m3VDil9jxXl3wkV+sYB2gj/OO81+jEBKSL6TNS/bq/icIoWslA1GsxRM1gCuE
epjOVZOp286kePu8x3kNHUUBNP37XHa6ywjDFO9LIcxMKWRqEgI6oy6inFYKKCLqZdpFhLya8maV
pvM6XFG7xrOAbV4j/kfcmxQm2nuVHrSRnCiD+/EJqG6JNDIgNbcU17ebQniyI/Y+IR20i8t2KleC
5fXfQBeCsi9dORIA5LitbQla91soB0H7zJkxWx1iTeiH0olFSM7kX4H9s51q6rQ2YjzYX5ixbuyp
wWYmdO/yWZL8HxjfgRp3uHz9RYjG+B19e0orYARRUkyzFEKOwsgBpICmC2GSDxa0S6TDcIOPinFn
D/Cx2/TrU4FbYP0YRPb1G7g/jX24GlJNZvY0RyOckmRQWE6wHvyE43QNQn5KB9/OHEQwBkVEt3wn
rnSsNl2J2xFreWIovQ5Ofwv+esCksfE1jC83NbLfINmFRnplXJjJbSmPArFW9MVk2eWa66Ha2hVA
Y47GB8OD08mTa7634W6g8b4scZmctiDrSzTGAuxsSrTQ7RqkByukDShk9dBqs4X9TRyXZ7tvgJzU
qgs3j661s7w8odM9/XUuKFkBrInOPkOnFM+8NTQn5galJpNF55PAs4E3bkt4ir11c4KDXuVFwmcm
3RTKa0vpXhzfV6MrNClj9fXUMoUMHa0Fb6lMGioBX+7qSw33XMME4+eXDw0TJRTdpKQWl+ZxJRWi
A32S+QNJ+W6/mbd+vyA9mly7Z+uSah6IxHJcK1DN9pvyXylm8V5gt3uK6qcOTVfUsFpuJFHBWUOz
HdMj/jaMKis5lAckZPVl6UeZ1zhxoP79rPW24IdPHqT1QG/SnTXRKssViwnJKsxWuGo3ieNeNkRh
dBFHYLaONhf3Pr80zES914WoAvWqxpvJpxYcCzd3JhiAgsDzyUSJweht9Nv99jYh4lTcYCrJmrBY
3oxMqHg1sppKOIbKvAelPjq2zQrWN3qRtjPLOHkWQXffgzeeVfSUWiRMw34Q8dZaxjTtpKQ8usAA
L8v1b9qe6IBU5NO3zcEmhsSk2tIB+IeA4/e5m52QaUr7FWogjMjQ2M3MdGHDv41fS0Kl2Q+wHaWW
wGX+qOnSvJgJpHc6FM7nH64Rz3BmgJWI9lgC4GCYF7oBhqQ+5xj1WC4NuSB4cQDJIsEyEVrNeyaj
gpUEQY9Ggof8PVKWMU1qekHiGat1B5CTjPTi2MfkF/ha0lYoOQXLPzPKH6b3hn9q39lgvRv+XqQH
GYahRN+0ceMlPQdRM2StEJbI4YyjLwqnGXmGBxDNQ1KlLgd7vG/Mx5c5O1RlqDKDQIWAJA6tNW3a
5Jil2eUbG1BlrsCGwWKn9KQw72Sbnxe1RS1pN9yAjMxxABgnhHG6AKiDRqJZxLfJxPwqPf+FSZxB
y6deomHrFO8zO0dgqn4dx21RUHJUa5/zlEFw9rlllSmZ8n8bNQkDP93w4IpgCJD3GqDhAYV+NgUw
SzS9DIPK6Pc7mk7wL3AWebkNgJDkhJFuYrt2DBLkvs7KOwKEvNGVaB2G3K5GKBvpprwvNOWQaW5J
MWxdMY8U8B7N0QA/FRqQDhtBCO/K9gfGR9kIc6mZ6KHYMBRPbRaZm7k9LgKOcMxtWKn5TN1M8DEw
DvX/mOAhycm5bDCCIWGaDqI7JH7yZZGUAEWIjPATCil6gJyq3wg3LofsmlxXs24SYQvUhYgDr/z3
p7GZoEra7UBrHsOjS0FkjH3eZzoaxX4Aa7PWiaAs213QpBDCapUkVv385geRTMMI/N4B52IH96Kl
N2pY4yFEiOIwaed4L21HPRHziekvmOxCJEXi9GmZrDSyBsRBNMZnJ1sb4ord4pEzjuaM3Y2gHhsA
ofrf1FQjH3h/XbEBOkL3tHgXpE/kvMy/NqBy+mnBylXXN+P2HwYddcH6gtULHgjswKOVczXKBRYB
QJFUm9eEy3JghUtKbNstcmrDNcjmcWytKRldHHI70jH8qUL+eTd9Tfk4WnFHL3fci3O3fjtLqQLy
ihUBi7MSparhfZRjjvRNm4lND88vCy0BuvEC0gRzoizoQRlEeSUx3jytPOU4sfuR48E62V3E4j0W
NkZEYnJzbhg8vaydpXzKiFNNLDXfWHH/skjeVJqYYyRJhZ3eU5/6oX0nhKdcr98zrUgaR86hrjIn
aWNwO4z1miM3enfAC+OoYyiiSRoQs5qby+X3PJATMg8a8vmjLkAwYUqVJapLgNMrFCzF3/Z9JwXf
vLyBRFje/HLMQkc8hW2jXrVyHdOs/7Cp7oKsQBNIxFk8lAOPkXMNQD/cBubrx84FFaU3fTVAq/lk
iSWqQp9zMJxUNFvT/wRW12OJPEzwQNgMtWHN6bYWcYAK5sIkFG1mpvj0wbILhIiD5HXpqn9W8z96
/fv2DKHPV6ofiTKI+fw8KLSM06JMYEVRBSO1eDOyxhKaahMEfh8bf++j0oPuWtz1XuhZqLV56e/d
awvPREN2/l+luwAUvOvAmInk11gXjwzLK+uamXDgdGQ68CHLWD7Ljbzgz/Igluimv4jlLyOMOKwJ
Cdn2blV0k+aH2ujGfIZPklmoZT6Y3pAc0gWDyxoQVvJ4u9jdDzO4YsQVFMaGShkLlUxNX3YpX6AJ
42buwM7BxVlldOi6MV9iDCkW98FzZSl2x5dW11WOetdweDE7wQp42fH8DtC4XZEFtk0OC7K+y8jG
w5J7UwURW3vLGpoi9Hr42F8L2WBf4kmP8WOypgADKDdzs8U8c1mN0/jrYmm4rALetfOU59SSVWOT
BzV016J+Qm9hstV1hNYfR1D69+BXa4ywNJXVGOyOWVIm46DRM5Iz8Z1FF0DEEvJbYwwKs9z1TfIC
vAtFmPcq79vto3ZO0QPYMvj4niqfDbGTlvN6i8feQ+sXakxUTpBl5py2pFgWdkaIYyUAkOuK9aAw
gWzSivBrjV8VVllPRuxgn+/HR7Jgaf9mXTsoIelQcQ4+n8c4w/2WsScYaDZmIO+Y1nUESPao5mmV
r6CcFzP+xRHrlhlJwvPldXFHeVNUxkuqC3BRjhV+jHCBtDOK3OekKihC2UJaRqFpUad3Qsg1+Bhf
RFnnjsErV03nr7Q42kOmuCtprG4Tik3ie3u2MxtHvnWqyCK+nimmFsngosz+FlnMBgbp/wefoGyx
kSuvaVqltr2IEydwBPyJdBHD4ve0VFVM+o5EsUzxRuyO0BIEiqBoH2/wnd8JIWZvf07BXVaDr5At
s4ZCcjijr/kbJOCl88ClhZ/Ua3D2ZW/fYe3YuSJGOWCOJkL0G73f79F5qdtcKRPwexLl8g5KgvSA
NIpPkxQGD0aDBY4qF54wKeYj28appIE4ll9ZMok74qj5degVLHSAEAtqB6lzYcIU2H6UuE1i3rAx
JI61G5FejkR6j4Lk9ONwlkJsNKALo6s1SePA03qaSAa2ZeU0oMFeaE0UPuY/nkaermaPOKQXUQgx
8bVaRZtN6k+oeaN0hqb/MLVUD6BFOIX0oNmxW5v1jCf5d2JhCopFXj/HN+q/Sjdonq5A1F+72l28
Ste6VmKgSR2wED7jh/p4icfrLaUpJC7hFcb9uRu/TMXUWn6MRa1BnitRvHKM+ZKo9xX9ErETaETy
1agZiRtWPmPHFEqOrnwguYOIW1wS8Rgt+u9+ykmjfZnB0HMUHX1/wiF8DkVyPhhk5pGQLBc7rkPK
oq6+I2Jkf+9cJO7GkRIVxYwCWNjSEzMcHK16hU+3o8Sy+L7ZvVecScSlbNysjRw9NSMfvtnO64uR
JfvF9AqG9ZOosuyaHLlFbMsRPBGxM+cCkqy/iJmA2LGjk2TLIij3k0OZ9l8aVxcR5tFQ1KETUIpN
2XI5rxHQFpuUQUxnAqmE25SXYqbb/+7VQVWhqXno5OgWleq480+BomEme2Qr8B8an41jKhUltXk2
v94zx6ubksdS2dPubRZlOjBgk+DnyBGgSbC3f7SpjoTBioE1zTaoRPOTF04msxgm8WwIdVR2YtMs
zYHcu0W0SD32t1ttOB+oeb5wlXz8d5+ckwf00QoNUe9PH1H5Deiit2UHi66ZXProLn2HDY5qoHzZ
mMvpM8ovWTN9WRK7TIgs67ZjjuXFmdJu0eWwyQ93G+quBxwyqZDdnsahj14Uov85FwLem3bklXqn
ZKi7kcUdqfEyYzVc9XVZenzzXPmtY+hMFNJNxFKZ2bFAF8uomSG82h4xWKhlCXnEjnQ+l3a7x0cK
4v1QHYC3XkYm6LaSBXANdVC5yokXOjWi4UkbmtmfGAMkfDC4eVsJ4lgor4JlOzZqtYn/mbJdO0Ha
aOt9HBZ2geBmKfzvbZ71ocyNFzt0PQ//CDEA9IuojdddxMq7hY3jF2DLFcRh8RusjP4JqoJ6qcP0
4HSO8MzR2bF891rHb1r2/ETXjf3AxDO1zlYSIh/42Y1ZfeU5V20/D+r9t2p8n9q6E7B8PmB3U0yZ
QuyEtvRkmTQl6tVTm8O5XhOcnEctZ4i7xVc4aftjoErp1dRaXPYcFXExFcYErpv08PCNlfTjyTo3
mnlTTJRbqJHHLMTEwhb18ZFGOrd3zc4XCcBrWxbwpdQPaK70pcakX5q/S9AEJAHpP9dKgUgJuqMv
Wj9TDhrGDyKAh56osn2X56t/mDkpzjfvmIesPgtCdoDr6Ty1Ts08R8q2JrIU2G6knxUStiqxmZ+m
UV05VDZ9u8oKC5xbMqJRUAUi5Bpk01ZYWXeGgPfEC9UmvVVWwt/IA07d1g5QBG8ptTCXWyhaBrpR
8rWo18l/QOkxJi49acANtlKgsWmo5PnbwL7UOHJKCcthu1eJNqPPK1f4NoElhWi8djwPGCw8bCUC
G5WNJvnUjnn8yXsI7Xh7ixTp2m36VNof2DiUKF88MQ9GEeAjVDthUndK86gqP+ThHmKIb67MBBf5
3fTZewDdAI/CFmYwqSQzzOU7geVfrN7mILsCtxwKzKO81wF4F2w+zibWFUP4oNexYYWhMOFr1br1
FxQ4vuCPX3Nybx+oYJZvOCee6+B3NpgEYAurShiCik6aqHrBz/4Ou0QG6mhbC2cUB6+QWmdv2sju
IqCm+c+OQo0gWN/3txxoeS7jQwCf9A9w9YRr2BOTyG9+eEE1cr9/DTiDCcjVrJJKmuZ52KbVmyg4
EsyGt8YiVNeuZDKzpis8PgdU+9AlW6wXJ6ITtQPqg8cgywJ6csDYvZkVfRUvDmWmYW6N6CorP3AM
rNFHXWqiSglEM3yGjab14mkUpaSn1lcA3MEi9GIl/sU/ObxalU77ZRCvTuWSE7DjtoFbLXsh22Zn
WHbZ84dnBZhcaddSvtN3hqcbDIf3WZHztSebUsQ3BSWM5+6nOreyYlBta24ANN1I8hTTooHm/now
dCuiMO7zUfZ9bXgkY0kQpyVqhbQz1UzV7/pu0MImd3B6zcDUbN5XocY2qj7syuNY5vlM9Q+c9JCz
ZPnhRZEBYrCXhN/8vtElEoNqgZ+1wsd1vpr/v2nhnPD4G8j6l2vI1K9vrUDEgVaBojqLaxxTyHzy
OFkVXDYNPJj4Trm9sf61MNF3MU007dJ91Nfm7ElFglhBswu8V1Lt65Kr/Fzkr54jCFShKD2NYL39
kXfUC1GL5I1RKDccB0DcEwMkHLde7zWWtE2iq7X9sDiOqJQJ1jCrySbq/2fNi6VcOOIUq7l1cK2l
+p42iBPo5L4dGFQNsrA2MiJ1BqKtXTmzylw+L69t+TymF0RUtQaGVnq0harjc2s02y5LjU/34hwe
iEp4Gek3tbPNo9CaS+McTqMFUxBzHNOQqvOmKzD7Na2CK+m10hCZ3wO1L787Nj6YROoK0BA/fKP2
gfvvGS4cwxa8tp5m3QBrfHIzukUUlHoD1+/K8rVrI5vtr71k5R881u3D0pOUVU+tOPzLkbInqHZU
dKSgoxgU0+W+DZ99+QTQGylnUKPZy6xtfPABVOt62UjlbClsaylDVAqN/uV1Lqy81jNbTFzylHV/
WafcD+KGJamecA5VE6fmCMBRH3+lxyHM7C4/O8vsRjmCOPog9NeCPQwnSObc/tRVpxl4B9N2Gife
9WBVA1xT7JWYPqUVcw3tq3HJl8dT1nKZrzFzvoDF0eUcbTwVprYDNJ+pKPpOpS/3/nm7F7iUnb4E
DPg2mQi0kkyVG98QgOuaVR4NC45oEeTam2vaBptAqHrTxvcY7c5Lo81ak6/D9+djhVy97iKHNSfE
ZUg5DOYFieCH0IeKlx8nvRK+BseEpZLA9MT8xp2FYGBSOVLC4Ux34Fs973OqFObaAhBB+zViEOBg
TC9dmQ/hCZk+xBejXJ4LQ6R7WwOxk69XIEQRsNozODl/5S5d/UZwiN0D0KEhp0TF8BXEJ81bqEFb
CmtOk6P3zCfTJPguy5hf9naw1deemveQb1tWDVn8plg/NeDUJbGjDWy3R/zS9Yi3o7JfE8Ohiy4i
wgROglM4Ben/GuuicnnzM21pC3jeG5jHdyUTRSzadz2u73nT530pkj/y58rMm5Uy8CrVuN3f8tTW
RjFiInew/xXmn9aBdu28Bsw95OD7VoGaU8dSWFvx5VaF1IGidJwo/IQo6Q8pWLN4NtHsdfAtFPZL
G2d+hRLuoBJmujwlN5VTRhjIpHJsQZ4qcNTaNnxHW0wqnBkc2k57R9pwK3YY0nH5yozroBH9wlT7
3WTcEyVFk1obPp2jPIZYu+3xMxetRoyjpNhzaYImrAVGguL7GQP6qXw7kB5u/tozaGpY0tuUeuxo
cJSQMcjEZtVPl71/Li1RqbuVS7hkrvcW+GTlzEQvMq+H9SmkGBOtT4hlmRUhkNQOQMTFklVJjg6S
47jvSnItxscxqxUPHTewqGEkxnMefA431wCE1ul5G/3nN1FJBmiSAVcpmkuRJyIZSvUdvpC/XLgt
wZ5Hz+o3huxkahANesriNocdhlCMlBJY332l9/CMJijIrrNBUjVzmOXxYu6Vg2jvrkQRnBV+hmmf
0QaTuhu+xbYm37TPJsdoeqmp9loIbJM6zfWbwcmpRHf0CJteSaSEjWG8WPTAeMx5g6JQ5cnG7dnE
9ntO6igMqLtar0kSOaqKM0fz1kwm7K/DAblPc2gmt60KPvhBomwS9jq9ApZqZoCNN71QdaMXDtpZ
mM0sH2C5pRKW58MnnEHZB0n3hUliW2YUAWpAtUAzmfMuS07R8BtR7KnBtPxtkkkdxDpIxXO5aEPZ
uzvkMPOFpDVgrvpDjL8j/1eIumANILPSXrcndKzGjGlKLMto0ZxKj/fBFBlER4vHlh1Wf4H79QhU
/Qu9npun0Ctw9SyxC5zyVmvDtNUckXzSpr+SMjyF5prYiOTsIUx6C74ECGLlhRneYyjS+GxejfX2
OeJyCPGlZCPgjTb9cCPcxeuJmQac1m9OTr+VILCXRgCt5Y7pk7qodZegVheGK4S4h6PGtOVRYoLZ
NYAqxtO71TC9BjC9yhURRoMMPk7nv75tKQ6i9vFVNLuPon1z/RD13h4T2OV1NkKp7kqyhBdwMhRh
uX/+1LHRbHtQTJcoFIdIUaYGvQ8tVIzqdW46GhRPfqKvNbzyTcyUOsbhKjkPYtBhpPzY9UAiEQPk
ASyuVdN7tCOeIp/s80IJuJyA2kR64EvRSG2E5ltYyaqrz0gOwfRRtJDKz1Oj0OQWKU1DRDiqR3kW
Ov3sxVj1qb8TVyPQ3JZ9Mjz+qkVRZhOKTaWqi710rVYhjXivGDs4KZYqXo+ZEd1q1MYATuHnx+3+
HQaFjVTC2n/tHdwL7LbsYjfz75h0xI6iXMbEyxQ0zmB8T25xyOW0EpY7bbBMfFeJIqCwpPrMnmMl
qSs4eF3Y3p+n5rvXB1Ik90IFwFlnLHafJyvWZNOgNNca4PWCqNmzi/ZfdEbNXlur3KTKmRLHW56+
KM9aFfTtmIcF0IK0svQ8yua+uaCwV9KqQuDqMUiDBfxAjoRTBLAYtQ+bpokaskS/A1OB4X6T1T6s
MWNX/HXIEAs1R8SVu+/JF5D9oJqINshSDcBOm2XDrIGW7SRvIQZRYCVUEx9Of4Zzf16RYvi9G+eh
mM7fYk2rg1va/LdsSTuRjd1C7kQggo0bndaPaeri+vLGxW10ZkKEbmqofpkAN3ocYHCxRtWJmjTN
uPXpj0lgcFLFWo0Lc68ztuYhtYdmgzGysabyTTt59qLruMcUqxgXpEZtz9Qcu36RZC3LEW5gIyeJ
NVrVVRV+g9SehgfobCIb0u/GxVS4tf5KGnKyn70rlNjzpGKEKLiOFuns/LnIr8lFDP+oMr7Ap7VN
Yl1l4qIuZ6bOFK4p0UqEmf0U8+5DFrR+YdfEraDVL6NrgxGjMHDSywupXN8jakZh1qeifY5oHPN4
YL0iYYi8NXwEaOQlrW2r3YZuOXPKgBC87MH30sLSgjrAnkqrfpcCqXfUsNJLrlRw3C7QaW8q6bxt
2aLEDRkGBwKfah/bxTYlnW6Kh4BcQdELqS0uqmNg+VO4/KInIfNt/ppaKeCT/2lV9eM/kROJIx15
5S08AZzu3pahSpyJ9HiOlKiVO4tcdugFPhWzY3XizwvyeZF+KivSUw+Eg2mtrnxykU9dMEnbFJ8T
08i7vODudkfTIVvmpoNKNNk1/wSu+WaEnLEkR2qC/CI+ORNjW0SdptFhu0CrR67IVPt0oFbz/8Q0
oWQdFrgLw4jlu6sk9G87x4K2udrqlgC6lA98GwexwKO9461cSpb8D6ifP+SOs8TI0FAx/GMMN8PX
AThLcaUDz0AuKfhwDg9pWxv9nlthqlNjzodxrkkINHcNqOV9TcPf1fpN3Gv8EBzdErqjX0FubV95
uidZaZWcm8FkBs3JeceMFSMJVM49UvGJ34jefw+9Zij6VPB5sHMcQBZ5L3xQQQO2aIJhDeeMBLJ+
50F5hV+gNWs1cFdzvVs60mxbP9NvFr5CSjlXx5MeHxtjsjXyQrGHGqhINzvk4U8oiNVHmbiOj+0p
/b6n3UCrZmKo7PcTDCQwXNs0f8nGudCvj+/y1s2jR3URLFYBzecQTMgno6fTxn94mpedPsUqg6+B
cpsgmHbdPPlwdLYhzVmEPMfYdgrcp/sdKXXkgVYcPrYSlLoocr7gvkdukLQTqpr3JyVt/S+D60HQ
An3vjxxI3j0poc506zdOascacNCF/lkq98JypYgdlMpI4GC8udeo8ZezHlzbHXX6ZSCP8V/ObLAp
CMm5NMJZJzvBzG/1wM+sbgTUeqWKfaXUyhgfEcMG5ZAsVDJrwbpmlmrKeHpz0C7WOfbLjKiV7cpw
5nOYwJ+aA5As4Z0yYhFmmaxh7SuIy7OmsShEjnM1WAhOd/xaYJH+pWTN2z6rPnaQZSZU4xViN6Lg
rV7ETzRQP4ReoIwPg2+IfgO0CW9goY1PhEhhbrQcMgICF80WTbSaEdmb+QwJlzTgYpoYsWDUfHkM
60EIP6GdexJP1Zvcqp2Sh1ZLweAr+bEqK5r6Ga3cWMXLrCJzjOPZZXHaR/fdoyt2Pj1p0+jTJ4IS
z+MIXkwgXlb5z0+XpvsH+pW+SUZn/5SAAZqhvs5Kh5r5YySGCuAFU3VbmVbsWVdisdhPZ46OmLsR
N2DbnyPfqjSFf+qAS1zv3YaCkJ3oLCYcDcHDoV3oOAqKdupIbw2ODbJDxIHG5OxcExqEzgjY1527
cY7uLJPQ18VH1u7RJBigeGwmvrcLiRfxoB8u2UjKsQNzXcqYZL/jfSIliQ8fZY6zlMN4MlSGJ0dM
xXqYpk1tsvB7ccV+jSaqO75vbYVqCDniNIAS5Zy6pDEQFcMk2e94qwpFzpWDc4hc3fbfOtnax/fO
+KM9uBPU7Xitc9J7ULI9xBCE8EPPSX6woupSI+0utFUiz0Mi5km5Wpz5ky7JqElaTqIlIlS9HjC8
bhuJ2NV+IugGDbN4wvGN29kGiEDvOp1wVGqwsgzbv7ZhyFq2uKtb54IkaY61d+OzYdeXBktpqsUA
0+REF8EAp6SdT8pfMxezomxUx3GNJPgAaxrJzOC1vun/WrwodwmyWWgHtc9Bl626CDobQT3+NVuI
YrgnLwbggEZJsHYQADiSwj0mZcDb6slGReLqcr35cSWL0hgl7ZU4+GY0rJs9n2HYTcTEKbBCNU3Y
1qF1Rn06UFjlMaTMIf+OAuf2vxNfy8BlkFCooZXADrj3fJ5jU+h2SHCH2Hk8eW7+dXuHA46dXulz
a8LIiegfB0nbL3V2lnxDAQlUzaovS4QFITv3tlAWjyBOQpfP0lSIv0B9xWBRuhNrJvFsAIY3KDyY
DD99YuhDKDqK0sAa/3kYCy5JhBGk3qnfgy9l0T4QI96fL9Dhfn67s6Xr11bCD35NKdBkmorg6h6+
YSd9WI9Tdwj59fHdSznDbDf/l0FWeDOqI3JAVAu9QiXazqi0rjktessm/lVuT2skyd184VhN0fFL
IeC9fw+v2gGtaGJH12Rf8md4h5Y6+sRwCX8ABxSli7oY6DTqYHzsAenoovTcM7PU0/aq26gKAYqu
06Mpfs1GTgFEuhf62dHJlZ445ZSZpgMU7dKwXbd0gZwc0ns8HXieS8JlgUyFH5laufHV5TNpojBD
JthlS3rIECyq+kIuHHv7N3OhC2yYKOhnLbQbSjGa29qfGFcq8s9K9GIt4cJi/3k1rACT8DrkRaaA
54JkZiXhDgwiwYyBIZWSMulG/1X98wye4eJJX57RuTaZDST9OL3TyDudVBR39rMk1fqTipyhd98B
M29jCAV4+zBqPSaW84wyGv0kKZLUGFx0v8QePLPDi/ftvmOQXOWI1MLftkz7qn7gua213qLuiHj7
qqbHW80MdpqpEFPgEkMQjXdvEpmzJH78gVMVKg0/Iug8Gt6XGv/d+WZnyZFXnYxOFDBIajDLW4eh
f02a6eXD/qRUHzMBcMwbQYXgallk0D62iS1PstAo6ML2NvScpP4eC6ttcl4Enr2WpSUfrW4hYMm3
yOKb0bSTew2OyZYhvvZdM8Gym1QCC9SoFvxoeH1RTvpCcr87tq73rL4ZXrhq7381HlHBCmvGla49
dPIoo7uoRsoCZU6MzcEf0Ku91eKddPq4jg6Hisk+0C9AHNbG7h94Cozx94kRR5OVIt54C8ksE1mK
U0b5tZft9yHzck6DDyH7xMkamV6/UUb2Cm76G6xK//oqi5eyBBB9Agd88lFIUqqWlqTGrOPfg5jT
feAsu2oWrNqqdTsLyJuqL28wGtjLbQTTZvvI67DPCKoQvk+Fjjd85PCmZKbn0JO9hdxTWoKx5TuZ
f2n372p0jPTJy9eqjo19kX3zjByv54Vivq7E3Pj3eItLn29WhlASLFUIaLewMOQTSFhcjrdUKjzW
l20wfUrNo7cAZhkMzuov8zHDy1MOsgzcymi1Qp+KSTX2AHNxr1e21bGXa8e/8X4VbSDNBe96uihc
xv9WXDoWlHDpkWbPOD4R6hjwuJhCBzwWlJA+HsTNz3/lqbv/6iOhLL9j4OA0t69cusWUyhX+4Yqz
yYJ+MrBO+SMQG3d3aFuwtV5T/RCefxjC4PJj9n+A4bDVYv63CGfBQQuvaiRpYHoqbIrQQWocZCUd
V6UbyC+COpR38j1hAxG3/J/yBRQ/Xgq/rrHVZGV92DDh/D9AR490I7g6eIvMIPBeoMQdtsVcn6V3
Y3G/N97aOuJBSuVp3iZGSQ3hMyRexZPCmVZVtZH9YlMu102NPATIJFto/GNx8f9Pi2RgvplFVZBC
EbIBiqHStMCtDjUe4gUzXOACZDfxpCDEwXll/a9gS4Qdcs2F92yFZBffMmWgaGGGlVjzg3Dra5R9
iy7/loe83j2J5qe7gWFpsWxfi72JWDFB66HPCSgeJHOHWwc8kQ6w8EYyu9MBMmDaGSk3M+dSOeZn
Injhl4as899m8hNItKvPhmKt7hjmpUdSkSKgJNHqXKDNtBJm1tll44WzHfjUeAnqwWc6NpMtrBXf
JpVkPlsSuyQlsnKYM00L0D8C5tHE2K4JPtmF9hsOHjbnHIRmnWNGbc7NOiIn1v7nUC/5F/NPn4rb
xPg3haonQ6WUT5AZypjkYzPS6qevHONDlFeE6Lepf4Pu8vLReod5c2ddUSo1rahVLCzWgOqyZ3uv
Y4fSHN+uQjzYawkMNfQ+vB300Vl9v7rLE2NQboet6WtjA0VD3Jf5CJvitZut4lh50d2Cm/HJAyes
OqimUB/XHbyDZirLvhCcaL1FcfwICyh+LGIrpQx/l2BwKhloYsui7E7ysQvPS97gpuR58CPwXufP
dBW8E+kYh/A2WvMCelrewCi7voHJKKqPBkE6uWYi9auAphmwpNC3QYJ2S4nHlGQRwGz6/mULCPd7
y2BfNBdc9XhVd6lP2h8oRJ4A6vfBlzfYEhcK1frJLxSAbVjDOKqeVZhQLZNwgDHyjpXEo3yc6uTw
N02xdkrUOXmo/SBgoJSk6On5dHdorROvg8Qq6q1hcjeCYz9+48og3IAzm1PKcH0e0MvxvhlvBdKk
Hnfr8CSvkjfwC54InWJTZDij2n7S+qxyVyAX6Fk9Sx9Ae/Mit3Wm/33uWvO1yadhiIcsjc3C91+6
5HIRVDyPZTFMrJcZTaDzdydr5M7q+bJCZfC/iniuhMzw+dro31/g/08LPAuiyR6TG1yrhdQx67Ix
N6W4lo1Yif3dBSXsLg1o3Fu8kZZcS4Y70OeuGG26QMhBlcH44BW5zHQHdwW2ErAxOlOGDuzxdWWb
g1fWgXDZ15cgs+YTyT8giTi003umj2z/jlppwW8FrzIzeYRPTekHJtYESV7d4qGTiagSlS1LL4BD
F4zp4xsT2YgSqJut1cqdaIKU8iNx8qh6u7eLTqpA2aN1j+2PUfS3vRRjJaf9aaJjl07dCj2Q8PjE
RB3o3Pr0BpQL6cdXHeJ0N0R7+9ZtYDSfuinQXjvccBMK8kQQuyjtYEUlrb5OlTOyDwYAevx7pJpx
DnFJjfNK/F5CxScQGq/2D33+FkL4zRmrYQCqa5hYOTB+fd7RQYhZhUGxltpTko8EOkt0N1Zg3kMn
4Kk8+ZSmFUEv7k5ZsF2WgmIVPjhpbYZD5LXdXdLdIdT0fsX+CGfPZIvDGGeqoNGHu6QNB2pfZQ0v
G22eL+47GPwOBeppwNWD7JH1fxZ/aKgwyqhH1MwS3IuRWDacFFNGZWS4AZI07MkMaUD8TUNpHYyH
SZZK4T7YI7fXpCiJ5zehtjjTB800LkGuYHKJjo1cF4txMjgZJjg/zAWgCb/yKBp2i6QE+tLUIQho
xNz7arEKS89tefxvmbUL08LvRbzORGCvaded/lvsfmZhBznVzLRY+saHjfDu8vifMko0delEGZ6J
PmCeRsvzjpeF3v+puDVyrETNIlv4wEH+RWMzlS0cSxRRyutQ1/FboeGYsfCo8oAjiXmKmCXAIbhm
WLMe24t4VbDANCoUUlnhzOvqWOoYWp56T31FMrgkB1ZUGyjOa+ec4ZOtIe3DeBlbq6NPvIRt3eme
veQfCibqR99x2sBtKJS4EgCcrzqQyHj8Pvdu0VaHE0N1rsEDndR0GXbKPUHCqkkNV9B1AbFyStSZ
zwZtAA0wibojNZM3id0q9OwxQk9dWEM+X95ciLn0Lt+PiKVchAUAkmIlGtU4rQnyQZIfh7BO0Hu2
NgMQR02g7BzuqPp1bFr0DxDWC1QAFNAF+ZsrnLZZTpOxegTXHwC3aLAVkV2wqLv6jx84bJF8c50i
fk6jqdKp23yYAk4Bwqc/5+7pK8tgUkHsePDti8s1PceKk4kts/Bpq1w4ERTuZyAE/yi/OI46sbyl
ye9vTcAITbDMVT9v5NF9M0NqMKYPzKcto7jWfIoCwaG/fYYCw8n4ItPuI3+fQYSU3j3XwGLColon
qPcc5A82vYWAixZ/kOg1sV604bmU/aR5Z+4eluDcbiaSdcMawp/nW5xTwynqFDl72Ja7LowHxveA
NhBRjytbucxLPL1zxKXYHf79vPEXGUl5H5xJpI4b7biy324PQn9fXWqNEwYBZLTMhQhEffpUytX/
VGP57+cxs/IBhWCZ7afkSdE4r30XBi2qEYFDiou7pHTKBFivi+kKS74ZZHr/rdWNPWY2h6TA22/v
KJNASOa9+YlOu08bm3GhiRP1RRIUKjx8bnfAXF/B8AfGE/i7lPp5C3SW+wiG/PnZd7HO0SmMZ5hU
FFanVqyRFpbETYvX9gwEPrX8pWmMaajaD7+3Wn4QI92fRfw97sX6In3IsatmuzsSv0M6+cpVuQT0
v8jHsB8KMhGXaUCndtwNPnZWt3tww98idvXQ3eeWp3uatud6h22dcdtZWZgFwqMOK7OTwmLe4aG7
8hjoXbHyUTeNKytiXUkIzWPbdLWnr/USvnTYrr1yzjgeArJJjzGDw3lYEi/aDMSCablmW4N8UNh/
9net8v7W8YnvOR+erijMeNSb4xdV9HyE/65E28IXGWWCo/Df6J2lmsu2gjD1xmS5uESxUGg1IUl+
jE1xWr5Kgx7zgjlVaCyx3VnJxzcURJ/ka4xU88Rpzfk4A+4qzLEOX6VoTutdmbr3Pddh6yR11lbm
n7V6ji6UbmUYWI2vujIxldwd9Fab3AgHk0t65HPE2/G2JBT0/g3Gy6TnqiymdLBP4nB0DlQC6XOv
f939l7erwZ7eJ+CnXk/MKR5bSbAElEGiM8IrP9ihJ/CH1P0HoRrsEDdX3j4nEvBBQKBhuUV6yjd0
czD0ROY24WkeVhVPyiFxXXESx6+aoLp1idN/+Y99K+o++9X6e4HeQ8bUKf/46hC2O8Row7llt6Qp
/LcJOn8vj0m9zN/Mgwlu5gPlyLGe1BtqlSgMzNKNqv8myR7mguAmyDyoQm5PWXJ7ML7ATY+2s7aq
7g0Mx18eaoGIdX8DwceaafHja/I87m0gB2EfvdHWDXnckP+PtXfClMmspwkjc6tmA9O9ExEKcs72
9bMeGxu4v35ujh7bRGIwylHUPWV0H5SdfEe5n419bmyg/bkwTmPvNKBxzeOEcK6AK60hj3oSA1ah
imPSEyDK/8LMbF/bhbRBE9WffwaAqdYR4iaNGLo4PS4cjt29y9ahR8ok1sh9GG+ocOE4GiBKjpk9
d3kNntS8pnRLCWd8qX6wcORKnfxYr80AQaTPA93TZa9rS4DV92262/2SldkvZG3BfNE50tNugR23
zZoyKoPvF0T3u58oysDIQDECQpXdFxKO2ow+KUYiaLpd1xvhMwoYdlRUU3mrcAVxNInnKnvupJNi
pNWStk/aKLhALWe4rBSLP0Il5p0e6FoVxqLuZRkPVzVk1r7+AKxSLMh9yMA4mO0cdZbPjiSqfIIf
IAtn95ZAmoO3K037Ox6s7bo0HWjVoM25j6LZ/7yNnpvVrcuTDazSTouFjpMsElJwSI/6MEhbVOP2
QwcnJXe0y5mFHymxpIMBj6K6zUS6yF+4IorFqexTPBKlKPYuXT64pIZKUwHOABQCSzjrbL1yYscW
m8Ge78yuf3TLXSTtNo4bZ87bjrY5bq9smhFjAlmP9rzY/32Q44MkH16tZpXqMlgf9aO7mKKpX6D5
9uzSYbAwzKyw8K54pR1/3ym66s2TcWKZlpEOEDLJV+rAHnjsWbbU2UKO6pVRzzf3ZYI3i4Fq1SCV
nPc1/Rs4Hf25+09FisvXvSt1r8P8OZNCGLOI0Cmp8PX8ADzlsHcg6Rj3Jy9t3n0Tscsx7UOJ89JH
KA+CCjAMGqnKqwuwdKhrwTUsYq88j9HuTiRfTAz+wCFFtaU6YVmMDh6Z42NJX6R5Kt2uFOEuTOtH
5yN9RV+d9AWZF8NBzFEVuP5kMyrA3bujC2XbuGoqJlDoJJ+zkf6UBMB8eWmN1jDb+a3js2rQ3ftU
bT75iyUTJuax9/FLAwqcrwkf3l5+ehM4VdVgoIM5kBmk+wCzQ6bBuLChMdIvvcTHfdvGTqV1yEEN
aud6Jnu47Og4q8c6fGehCptQwgB69geyL9XGWmT1rHRN9/Jurd4cjQi0kJCbhBkXCSnf4VhcoUA+
NeME0itsMyI6/O0MNITTR76/A0px6h/XM0DU4q92KTQmRe/DgSVyE5Dt9EXAWRxfL0PJFS0W3Z+R
mWD35M4E7wJfUKJeHoJCfzAiNt9opxTLjS+CVEoSu0D6v3c3AYJrmC6xCaQD+TxDYa7KRXnqy6td
FnjclVpvezXBz//VaCefvEMKZVzmPbu9fxgkUfkSYTYD3qDXrzc+ooobcKXBIgAI3sF3rh2JVizO
cQwLKURVNsGT+nrXOt4qMIVkrNItqdaCRyaF9hPi1XEO4zvdjpf8/3oM5P9ee/y5zBua2Tdd2o48
z/sMh2thW2NqNi6Tc5zR7YRtZVbKaMXe9P/FpJV6aJSOrClqklN0Ahmip2h9Uy8lHW8K7GZYLYi6
5oge2iGUi22AOfHtDnAVL7Iae9Kmty0fKthMOhvkoeHJJ1LiJnh1RXfOWDA/8GnMf3YakuDEmr89
4aL3ZrBq7na7VOnru97zNWjirpSzkVmFJtUrOxOTbaxvUze/O9hX60NemoMXM44FwOXZ0tYduckn
57MD49YFghNyeHUBxPgFGkH5LZ68e96TvUwGinxoML9CCeALGfYA1GHdH6VOmJL3qpt00axPKueW
Fhsy+5dL1PRVgv79kSMqEWejWy/erKyiEJ6CVhTkRBTkYCoGIrv3Zr6pAL79qbQ/aNRumY+fm4C1
jXjiwyZw9ZS/3EFNg6Czmm+ml4SeJx4nt/sRrruqLL2IBC2+z1X3QTnSvcV8CyD1Fbmrnag9xKnI
o6w4kLlLkMrN46Qo8o2xqqe604GdW9oBPoi2tI5i5ux6O3XFhUOao6wGsVv35AZg3c8hkTLeiJKp
0i4zvSW1kDXG9f532HxHc9wC1i9a3njjytrQNvU0nFjDTc0MFBSd/emPQbzLs/P3e5GmrBKSArVX
C8LjhFKbVbcGNb9t2deRsCckzwR0eD7mkXz/79r4MoxBDV/KKl2lwCaJYwD1cAbdM68A7QLnN7Ni
GEZxg5o7uefzc5FJbesnoDkeUxmoU2VF15r4sem78UE2+i5uVnj1yk1KRQqX+1BDkH6PM7iSzrAv
rHfuvhbpN7xaavuPnXbiqrCJklKurO4iXkvz5wZNNlBF1JfeEhLo68TKGWilHr8IkIznJN44EBRL
92R5xWoV4wf2A2JRqonHkXRrC167fLIrctdy5zH/1yE+yEATXg88WMrL9BvaPA36uW29g56PX5gX
y3Q6q9ihwY4HWzBFcyKTIfMOviSN50EOBd5zlbIq02wB9Tb7XH3r4SyyTu7o7EEhvEKLRiNDOZ1y
GmfgCAdRKpfs/HUkNZxdLzMiGPL9Zusal6z9BB1ksPP38iA96l87MWaeA4xtLdc1RSjzzVGV3AZm
zr4S/Oa/YIlGstUbHJ+H4wq8GQ1B0TR+iA58gXRodXd6br1StO+RKVv3ZWsvcQXvJz1hhpRmF1My
0OZ9hndyqTOexNwZa678bhVnP4mQIUeuiSGn5P36zxnj8LUrg/jMe4fm2zi+PzGT5l8CB85wySlz
RoHCRVbvpw4WQ6m2yVQXS2UueHrHoo0v62jzctGOl/LyUnyxpcReFkJ/1BsH0d+fF/iCmN7aOlps
WfV3dpY8kiJpJwb/QmH35b3kuG65tzQg6vSgjJCg/AJvLe7cyiIpPckG7UBBFuBwRe9MsiEMQPYB
kmPj4K1RcSucp85V75m8doZsyUGmyN7saaLyXBO0AVA1o7prqqdZ9QZMfe+c+ukMidRW1z68vlVI
qKCN06ShVIazttGgGJBCVYYtggsyTfXyC11LsQU8427TSc+Cl8hiHsphRMIYSzOalCUm74EjvzIR
YukwgPHLnXTYxjIcB7kjsgIeKH8Hx/u7Pc/z4XzX7M2hnMx1pyuaomW3DalYfStsTFhDPMP/Jz29
l+83wXKSC6KDoR1eSv2P+wKRCjMjwvsefcp1mIS9VDbJFzxBIjOKKcdtnkL/9uDcVAFvgTee89md
XCzZOjNMezMyxkH03v1RnYgaaglfQg2YGQ3w9+qjUanzakNutKjZWgu+oZf7/3kevnuCrWZHQJB1
Fa6LV+cdMDOnBapgwV9KIvNUOFFgPGK3kuD8dc+OSPUKAnBRHh24/UwSYAjpy64/E1hFpjGzC3CH
vggaodz/A9WLYZURqDLtVTRLkrw3/AYYyqVcZr7VCc8LxRhT3HlFL96K0uf61L/dnuSNA7LTlThi
sfCuI9/Z6+sQ0rnzxYy7Z6LIeWVOC/HsqwXRcywJ4kMQfEWKHrmP44MgKLDtgh/jgmtvP4yBlST0
kVSkrHxL/FBkJeY0QHRD0ZLcDJx9p09+V8K8iGFiStdy+YkutTeaEsatzcQpKMRqu30ETGmeOJKr
JSP/j9Kv9hnN+nUNrmiK2V1+gkWO9ElPjRjBAVlLGon+pxL4tSCPkc9v8gl1C4jrmmzTNOwcvtwN
KNe2KeEZCCftdi1AY/Lw2wZLRdhUZKUf2LmBwnFE0PwJGcazU6PfuZNMRSNAxoY0g+o+bHxyR9iT
W2j7A10BBxA8CBjFQhEngn0FisdVvm5GaOUG4nZpDGJ3Qu8Y5+P5IOOm0WyFvB5qbYsfJeVP2bKg
S95SVY+BMPfoBKzzOAi1TXrBwkI3gUgkEMGCTUm89AKcqK3Pr9xD5HropIMhDpli8KdciwNBslkL
kXh5B9y6QZwOr7r+22P+pp5cjnnTjdU2m8KqOrZ+XeZWd5P4tySA/V40selCEOoCb8WUU6PL2s6Q
xG/S+K14t4TlXFcJpn+/mxfeBop7X80Bs9tX1/DJwyWv3lqWIHVp4AobnblfTyXyCrVccPI0/i0y
3xAjclnrQlIIQOWQ5E6fdmD1GGgxNMtj/Ey2hD7/QANhiSBkX4FdC0eILlQFE/vEL6XpVPOI+5Q+
9dfzHbhPtiXIaV2ViijQ30ZSYVa0T4K4CM5u+v6AOGbvh3sSrNtKJaviu8noe/Frx/C1yHPTEYg4
S7fd4h2t/KxHthpkBBM5MTxcP1/uVnQkuiz4PhR/igio98Cxk0mi5wIsAureVLdWPm/cZtgcKRhR
R7X3+Hqu3eQyvEwcMUwlTLDqGPgjAa52URNlit+/KcCRTFtTzhSTDamQoBDmn2IB2anAm8lG00VR
+tPvEkXzCnmKH96oYk7x4BFmBiOyPGRnTk4xtItGXCQbJ0zTqPAT3QI1A4UFKqwrD/VnG7y5VrsQ
59wC82OdF1J+ZZseYmSdW00qGyuiMMQ3134Xe6ybeU7su5fUbo3DvVhbrnu3RY8OufMzwKhnN1sI
8JYTMN0ngxQibs+bjVJg8SZ79ZC/P6sVwrlD8biUbZwAbBSaG7Ojjdqedh40kUPO2i3i1i/EtuRQ
tQCCg975IbNd5BGtNY9n3iZWfQ9DfBqHVmru46qjjJ+EB+Gn+bfUDE1qhxETaodbFH8NOjXk4mOZ
hVERs+8lK7CVtqAcCOVedov/X3F08skUHIZvHT/wGqQsk78iLebbVjMzhHyxADdI56rpTcgF//s9
PT8J2gCp6eEYhCk+dehf3LnHbjU+z5P1x7y2f28sFGDpbwX24dNfKlK6Q1PHEXOQuu5WnZa1BPjj
9Wk02zLU5O23uoDmzmNYB87LZEqAzKFW28Cg+/1BbBGeb7KCYx1hnZhEz8jOh/HuSp8X20b1zk1Y
LD8RoA6efK/W/1LqlD0QqJc4DP8Gep2aUk18stska5q10btW75UWdYmjcyRTzcn+t9ubSbDa0v5l
4NZmyMumLbwfjJlN85SJW15AA0qkWFEib7n8lhUR2T4NC1x/EFnyRY/m3ZmhRleo33PMfz+ifFoJ
OnTGar/GsdpW66pPSAPZ0xNN8k17T0R356c=
`protect end_protected
