`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ROJdh4z4g7S2wCGsWNNLLZ/swF4jQV+MSi1Ipp78aZY557no/nhWLQdjyukwz7teqtZrJ6UU+L1m
uEOiYS7sl/WqLaiqPSn5Ntn+kA+HXarfQuLvb7vQRK88Rjf2e4APRKDkZiRurbugLyZ3MudvGApX
PWTJjXmiD1UpBd5mtLJz4BpUowQuJUvVw8jH3if/Y37cePZrxWoFy01ZkYMvqq1wBlcG05Ok9Z3d
MD2RHEhjosK7u9huj7AHBfEX6r+0x6YcNJzzysJ5j4pgN+2AQPZhl2x0xyg13rQs7EUZ4Af6gT5O
sxEHAlj0rI25McpXALi6LMQWsanTGLEbMRUQ4g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="XlIJ5H5N5J2b+D1VEN5fUqyYyUV+gfjMN0vaXG0IY/I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8752)
`protect data_block
N4GriWdC3GWZgJsctA5dvSYpqvJmot2Mv/G+dMpM8d9Df1Xj4qzWSIQjtWBAswn3ot4Q3zSlLoSC
dJ4T3zmxRiL21/jZS/LEYuAPjC7QF4cQFTxDi//nF+Ns6QI/v0qsrIPTqIS83qwgRmEMXIbtHLJo
0nuXmtFA518jC5fEWWj6QXTYBUTHABb98hMbnm8eKN+KOCQFT2wurHgHIXK/VaAEHcJ+2Xt1eQP6
u9/sEbwzzHWNu3E+EaydW6exdr4HsiZJYtUJXOz477aCPW1X6JhmnXWoqP7xSNIE3N2egE5kQJGc
jmd12BTJwaJ2mKfSRiI/JhVK8Jxp9H6RRAMqgyOEJt0NkgREpKx3zDHtNDQW5dOhONLFbCzh9Nb4
N5YHdXwqV2O73GxXqgdtdWzuBJ5XfGPBiCFFAatPyRsKf42a6AJle3lKmaW/DFG4A7p4MMpPNtQ4
t/BKqQNS/T9+IlCkB2xU5PWjh41pXEv9bvTaJ5Ix/r8uJ5M3V2FPjhYdYD1TJzLvHeFWgLjN3daz
9jv3aCCztWw+Rn1+JDRB8kNRG6hMcCI2tnR+mSXs5wcZ6vJ7LR91AIhmySAcuc8k7GFi99npUmNg
f42eCWMEK2w8m5aREkb8Vq2r5I0h6Q3njLwFxiCkGeoXEQwN+W+xkVvSI9VqK1A0NlHBLVw0Im+I
9BkD8EuUBSIEn70NPjRkDnNmxvjTPPFAUKE6SRUzxa+/7LBXfOY6vuQVQjVG0SsuOuXZMF2YKPQf
sAkHK+MLyt61KerfuLwKMSLN8spogXkaTdHV0cLVWSuDP9hai0ow02hkER4olRjyrRS31KeIaZB5
VBuhB/S8HSGWLF76+eUgEVHU0knbgjy4WFmfidAu/fviizigjwsat48b8gVDNSuTQMF5MSU0xd5w
BOgJnOiD+h0lqQCCXL2uSLrdCDG2zrkCrVeGbDfOQCaF/b1oNvy2j2TotHKRe/mCEv9GYqUZPydG
c5vzLkhH6B09vvEb4HZ/GLYT4klFxmty4MlemHUROiqKdwdYRHV0NLylLWibEsJJtXx81KR+chzG
O3ud+qO8+Me0/4ko51VJgDarLedqbJX5pGg5das6Gkv5BPfHFdv+nLoyBGMucb1IGN6H9CQUmmBk
PrL1unIVCwRuvN66NtHvQ0tGYEEKg+97q+6HyWX2a8Om4mgmj828IFsuKFuPUB4YHPSqh3Xg8W4s
KuG62PndhpSsIz2LoOpZ5TtIj73jBMo7E1lLIn50Q2NjlWy3YD+Xcwy9U1Mg5rswik7LOZzs3wRc
ofCDcS47j756TJMt9hBZv4K/TiiEpaRKkd3igaZydhf8QGXHSMKEHBVp072IruerZ/zBfWaaAoUD
nmlR/8wEzxI5Ze/HoaWhe2/GzfYp7SKqaXHDRzwt70A4R70KKY5qArmfQ+z4Kk9tQI816N1cChB0
69m/BjpRYjkaULa9G2WZKqSnF1FAgex9b6vpwZkjvO+cQlZjrGJCS85yDKY20nkBvwjgxW8zl/aS
5589lfqELiWhPZfoqPhM4bjkwERo1sC0tPQijrHkgWa9w4A+Mfpk5pIr2clxg3bdluNwWViHWL4W
JDHzu7uz72c5FXMAv5w48gNWa79dNTcPt1xnoZlp4Y/Gt9MxvBzEaz05EK3PkWpXE1QUB4th6kb2
SRAsrSNtZ0FvN2NOxI/rMMt7w6hYsRyMBJtbOFWgcGrqRNAteIR/yICSFUrEgdt3kTFAAB7/5QEx
F0mSb8lmYnsDtGKV25T2VLejLO5DTusrd657PfenEZVtTsEmezHjUuR4tFT0aCZoZ+difBtVbTS7
PJC28Kuvgu94sczBA95U+u+gLM3iU1DRR6UI9+zx/bmTOfT2zBLg9BMqo0YNVkc/dj674YAIHD+X
AMxDNAemOkWUxLmX3FptS36KMgtefDZESuJzt8ydOypK9SlhuCERjGU9XsToklCXoVmJNFnYxyL3
9+/7cZBb4sS48sDy2M8j4icHIG6mV5a2MK+tmkJ4hWxyecvDPmVxAHuGt0peTbzV3mG4xaKLixpP
Nel5dFgdH6mPciGRxVMxE+UbhWR8ZGahHVkHGSDQ0tBXVHz+0RYx5laf2a1Q2n23oJ7GahMimzEq
dMwAly/aLOeLz5ouLAL0Zdb/TyjYFzJbT1+uGbTNVOXWioCi6lXtNWKSTujTl4t468zNISyBH9P1
PPdoKBDwslAQw4ZDl1U/DA/ElAYyR1Jx0LKgW+W6F6dBzka9IHFUdtf3wVB/Fozi2GIw3vbf0HQi
oRtCyVAlL/iCSdVazyn5KpG6YwJ5AsXqSWm1RrKH4k6CRPdPuJ5dTO7IYvSrF49bHumtgbNMla4y
7ltwLO9OagpEn/ICbHaq+UPsMElgt9VfUsYNbc6FI+FBLHbcrWB8sq9QnuWPoC6yCtPVfhi1f3PL
Mn7rB5N9NiRy+gDbqAxWMfx7R3DZqo9B2OlzNN6gpNTxgOJB1KQFoP++rpVSPOrxO5RrTkm/2MdQ
e+e0KrFwgTBNTxvqC0jJ77Bk7aYt1+sD6NU71IzWn+1LNzN7u4vcQC2VpSm+795UwcfT57gFCFgu
9RTB8iy+P7qX9HegyxvA0NrhyvmWBaW3HiPO0rMBHuwDt5hKz/5cGMkk6rCsszOlwBoS2bqyiN4V
O0A+NJl91d+8oxBUY0iay0XR5pVmeGdqK7MxNtrRFRBZXxik4HdG34hxAyTjKIG7qHIWbSGhyUjS
A4vqCR6aI7GhkJk0bP4GCL1GqUeAgojxqaF+hU89Kr20H68zwT0VlJ1sDeQEm6A4iutqZnQr38v8
1kE4PP4/WSKF2JS6tKuzdEcA/tYZWC4lZR9nxXhr3/AFWiiuG3vad2NdxZXd/ok3s6tkwRCkIPc4
AQcwJ88ovpshwxDyQmlnPksd/4QcUl6rj4Pb1Y8rCNk2q57M8TzvO+oK83570Iem2B7KVRSqqCp8
gConkWvD6UP7RzmsEkNVyYxDwoq/ycRjKg08rUejDpUi3dEM6An9yuDSESCNgiIGRqwXjEvEsEMa
Y9Xb10lRvpeIDtJznRKhzNyQn9Y9r0DCGja0WOJFAFcjaqqpxiYFM7gmd5mQagIxrlEandVlylqk
dka+31PrRJvF+yf0+bHtMbxnG7GefhYCdL0+QFWusAK7UOl5adIKciSmmW2Dbh9fcQwMJNnqKTmg
DCmoAFZuufUNxrWpex3zJTf1o8DS+YPg8GUk28/Wc1mWzWDl29wNaOSWiDJi1l63mmbUZPFCS0tV
x/fkRNVRtSapnWbmHOq4Zz9k98lISErktfLisrOP1380V5Pfp0s5egmz16ZF3Irp/y/HFCDnTGGL
beZtrIm8p2kSV6jJo9ywe3BzWfoWEfLF7CGP1129xIWoTltGCynen07L2vfK/wp7/wnHWNJ5P20u
YKd0Pzj6KKmaFPMJb6gmiQ4P0UZXR0OL6lBYYsN+uNMS4vH2T3oZT8cFDXQv/3XATY/xiURH6PvW
yz8ed98GG7QDTwg/+/S5dLsj+fBHVIjfH83OPfPLSp4mn+uE44Ixpj02DgEUYIamHH1k/9bTJ7sn
EHeLfDrr9VW5fPXcT1yp9MmdpZw7Fd/nVZjAMLIQrXfzVfLEFYJCHepu/1mngM2aipFoPwLin5rY
UxoKM9x9/LH29O3H8ysJbrB5Kd/u2lpX2LghmOXu0YBdful853Lb/zFTjBbXKKtDjSoqfGbB9sIW
v1qMOPlPUHNp830T669jkPJD+thvjjuyfPPeznQsR1PcimJ7uoY34m7m05Jg/DdmIb0EJUqI+9UV
QSs717CKYX00nDJwZeBfOGk28Oe/o4sbqwRb5oahTM2hMo9Mm50Lk43QPWpuez8D54Dod0v8I3l+
6LEe7I2aVaw5CJ3SpLyncmCOcn/1JIlG641e5qKyEedLKtLpvmA1v2sSKpNa/S5VV8H6LUdsEan9
lUogdGBON8zK/a9T8hlsGmzIcfYMcFef7rJKxhgop6UUacrDUDSdoduLtyxMWuA5udZgQIAglMnf
cKdmOY2Ic9NqcaQLyG/Z9h1nkZ4aDgz7cIPLEL5JZw7/qntEdAfzLBzq7rib/GE4D7PgdO5glXKq
VbYlhGyd0uuTabHnYiSYNSTm9Ih0gF4+ZYWlTSCYbt4dt6tmkdQlxgGI1b3XC4NwzY2Vh4qVTiqS
13xRI8lWR2h+iOV4CdZG8Kh6pJ+XWqilRM1g5DD7L3sD5bSem/S01HW4snhUWB/Qawtj8q3oJrCW
vxcsr0abhN3T3rtixnDhknkjQrqNUmI75nAissnRuuJ3Entjy4ex35Bbt2UwS4hImOp+fu4U8Abt
ORYdFVvigcFrVZZMVg5f2JUp6gWQPic5k0pExiuuRug3QuAmDicbvmNwL//3Eo8///njEh2hCnck
OMN8GfUq6hrqig5F8r53Ah0iKyihx0NzlbMDOTWVftiHnPvhIg6ZamSzKNNhgHDYrWd58kTvNHfc
b3acuhhocZD6GvScV4qEGKGLte7JKTuMFuggFkLzjWn2KpATMAl/Fe4R+oNQGn13zEfBGAWvxg5Y
w9U7D9tjmB9ZXXLIVbuCb+g9s9byXbtcZHoEARPO8VMm0WZtbVVtb1FeSY5UeIKoDHwkHbW5W4rh
nTzaGxe7D5ku1XfTbLZF5mGkRmVDItkTapAPpt8LtMNE/e6xXPZQy65GceWOzl43tWrjmQwXGJMm
NwVaPsiXEH5xY/bGXzQKtUpP75gHkWfoGxM9IY3txc1sqajtEX74RZ++ThWu/BUQ803gutT1wbGA
omh/u7iE7XnxbdT4+iF93MPv15ZHbr9ejJi9Q3aGbDIDLyDG1KTIjDb4rvZ2pGsRsxkBf7e6FnQF
8cdhUn4WMbeXphv1PUV+u8SkpPmD7cwuymacjIxKB+XcAUyuqQLavb9NWTxuMNfxhl/90Re9dwRU
dn/262RHmELVO9JNSTrqBNlEFMYXBLe2NV+/CPEHUwnZgQxW/sWdApnrTOZb+X9S4QsLbls9uFPF
6sMLujZYc4jqWMlWcTzx9j6hDcr4Jb31csNQSqXp+gQ0H77iWc/IUddp2mxudvBkRdAC4FVjnmSw
AIt6N5RmGsOWTkKHGh2Fly5yvg8d1OhmCwoL64GHH3wolc3PWPYzGGma043VwOf+64VH+ssN+FcQ
WbquGQRBjf+Wb4C/Aa+50lG0lgV396Gs9LtMe4sRSxm9D7pttGccJ/z3iLHKH95W01jMt5zAcaKX
ICtE6d3GnH9SjvK89CNihve+4UK6E2ThSfR/3Y3jE0p4p1aqq46IZ1VOHXPeWKpSdsORQEe1GKbX
fD9MidtcwSqD4AqnQkhcGpLH8GlwCWDnFEGgdPQmGvgSP+YS7ovixrHaFG4Hu2kLQLZk9y0CaVAf
KRBoDVq1bcaCXAdD/QcLXJTTrzxWUDZ7fdG8NLSiepZpRPjgXy2zzD0P/LCc4YIWK7R7EwH7bpAY
gnk5+2GYN456qEsjYHW1ipGcZ4/7nv4qjdH8RyIYO0/tfeKGb+IdOHTUVDsk0Z0GOzCgD/MPyC5S
83baULPfyPYKDW3YSVwG8ui6lx3we5vZ5MuEOhG+0XiFrismy1f/Cmssyk+Pae2JmA+OIqfNP0Eg
TkvrHYggn1N3r8MqqsLo6UagQQbTRVRUqUj0Ojdt/Jy5aC0Jp4l/NIMkPJCGLDiV9PU/aMFLz5RF
IvJc6O7nxweEyPug3gqhdVL4VA86d+YuGSucPWsZ0bPZx8ewYJXsibljn9++nKpgQqF+J8JIo6fB
HqMSMCwPrCivaVgnB/M+rr0Bu4JJX2553Y8mXKWyNYgbU2MkS8bxiY9W9RWJAGjy2ZvPJTrBtT0M
bpNvix65aSyBtHTx2AqLD5yIfNR7aDnLNG+8qfbrUu3aMhtH7bOw2btRal2jCyo93oCONJlLk6Ud
O5bbeBJXoXHHiSpRcZiQF4xR7tNLy1tVCpxyxkoIbotzIpB7uMt5vr7GiXs8yfY4ssU8i+UosOsV
W6vXC/8z8FKi1TRTP1gtVRTnVL+m0++Q6s8nYPJMRr89eMwCtCXUfI9iHDNYM9LQhylgP4XNWltp
fd9Kz5DdlcrkrqaVW38OwOna0aXpPMo3Y4hsHTMQgNwuCGeYlKJIV8RS63bWPwt6oxdOmOtTNHhG
OxVxNIHK7mccXoRTN0pgqANX0MbBn5xphdrSNxuKGf7WRhhJtEwcw/SpNp7zAiPoFVQqqh0Pixe9
NA6cPDqGdqh5amimpdjN6fTgcT5qDZdeuwi3UrsuCRyule1HmEZK5QcdTxaMTY/sWlcnghJkJfKo
lKhh4ewG2xo4ZjV98vu1MUJcRIlTlR7EeIiAcQ3ODDEgkhpvdTMuAabBwzFOizN90mblTenqHTyU
2pM8/ZjjwxGnMlkB7gdxnzX1KJpDSVMmhEHazEFWMfgYgMIrW6z7L3NkWbn3x8j5/nhOZIJPj+gX
yJah76C1ecfCwuBIyekbTmGZ5l1iRJliOweRMmAixGJljQmTJ/DU+u1xXSwdg3W9uO19R3eUpaHp
lboFVX16Ey0CJrgEBYyBhVARaAXgRPzDqTj0TvMpcg8IIf5VNKcvF+VmEWVU4JTTwph3jTqv0Xyb
vWPr00pij6Xpg9WnltiyxkN3vZszKA5aEm/BLOozXIirKfqdn8ZYyG7LZpnExIyJN73s9RMnAd5f
UjSinIIAUwYiRrtPUbyvOn1vrz1AUCcjDrCQUgal8eAf9a2PLDNDeeOBvPiymusL2q7LtCUF/N5z
GhVKa9U7WzVNYyVTZydscDCLZldi5kbYj5OZYFHOwDifEsV4vp8ddDvE/Du/zMr2AF2X8wCUQfOp
thRzcN336BuqU/Egn9ZyI3mi3d1331Ty4792Bg1S5G4BQshcImxlM/JcMbY/7GIwGx+mX3thBJkD
P8T3FiSKEURcVbaam33VwHJHp3ReyTgNXktL1GhFJL1xuLCDzsRA/PuHG9dD+t3/QtSozHiMzWfu
9jiOd8VjZEgAYBrPJQDcPVsbcUMk+8TgpBgTLEqiJrO/6bBut4aTX+coxB2w+w9cglp38dmPm/60
nqsU0GRYvDmgqcF2M3hHUEgDs52Thj8tWJ7cR+Lu1qilLf6ZrFljVnzWdtGnjmLXp1z/4HR3mE9Y
v9tqRpEC3gIKxyJsXr7UxdQdrWwXKceKIs8/LDJJGS7ua28WgGyE1f/Mf5NhWVv9Zajx/o4Orsbm
f52kYB2SgGj07Z68lklObXTzKMRxbraTpX5Hz7BAMvx9iKlybpBF79sBmn2KlprPfMxb4AF/PJkI
aIRZ4GQP3js+ZKiLfWGMHnnmWmUWU4oK0hQDuy5ZHFNmW7fYVwP8VYk8Q47Efc+V7nSr1G3X1bHq
p1KyNv9wunf0kNzG7V6nIEBcjwg0iiX2pQMUyiKqGAe4+Z+h6f7lFdRTxVtojNr3t8sOO13a8VT3
g5vXQsvP9EHHnMscrPFva7RoGEDwBQAkufta0Kndr71BAr3ubnMDdmSRYcUa8doAnLIzh4G9WH4j
MJhuITkk2agoKmXeV69FxJbQhOJgFqkCV7xq/7VgITMKrk1UtaMhL1cCDepvMsMSMEt01mgl+q2U
QDiHhWI3dx3OVk0OWB0KHSrfNFC0sKDcVfyOw30SI9aSJCM6Dkjut7w2WG7Ba+XJmzC2Efw21/cL
qG4/kzWXsss3sQev9t12uQAYBJCWmLx8U7/nP5zGEdEtaSypNHpr1BfyrXg+Xg/vwn846kKPuAgf
OuutafcQpvSzCpsrQGsnwOtxlHU+h7rXxiBHLay8dc3fqIVfxrcXli4F2oGMgf6JCV/c6AD6qM3P
4p4WX4L9lwF7UL8MjjITOTsWqtXVoDHtbmkGAoHnevKdVcO/1JQym1ojrZQGsdO0nigHCGl13MG9
6TA2UbiH13Lgpnc/JW2iPTVOE2m0frQ/p66xi5LrjzVQ2zgS5CvuQRbFOG7GmNpXS5NuMgbUeZ4z
IiWKU7l5ASfG1+DznQ7dIwKPkROfK0k4Xiz7GLuaizq1we0barZUhuD9DAeakgBzAtSxZeowIRY9
5eUZfjbgWq86QEzcyckk3nc+fAMF9/QFd6ilYUo0dm6L3n133eZJhzRm6GMypz/Bhgvi0eGL7Mch
O1vCw5tUYrM4TbOpQ3aLacV//ctw1z/uZ6QVeZ0OIJNVvcKFf3tWPbPcZgfGZQa+u5ysdKLb2ll3
9LiT0nH0+/kID0Vg6DnCH77abJo9RGljsiBSyqkX8CsM35jAmaADBuPdBbNvTNmGMOkpQTCiu+MD
FUDjJxwH9Ud889cNnEb9nedGXowvfn7ZYpaappdyB65WoFe9TH8SsMmBG5hzEIHhr5ezgV0ss6OE
KJzfEOrKd/pqf7muHHETpoBQiKisUVaNqYmBAutmguztpRZFj6TnCRJhyGVn5RNhckIUze4+qVHe
isLmJCeW1leS6XvzwSsgjsRKIvOFoSAVmclLL5XBoa51+hd6G37F0OE4A6xtz4meEWURP2b6I8TL
sXoqiUp59dldBjgPCYzcsw0KyvlMTae30RC0ipU0j+UAzD6u5WVdR+nr5bsC5UmBVEzHOKLTPCZX
6zECBgbiRfvzOmprjLrvoXrSDyZFWCoUnJ4WQPsLkZuGTddn8SPu/Smv7/7xbtQbiBlyCWKKtcax
vgY5goVAi+tZdEbAfatd6NNZivZXpJd2XeSZiE3bDvFybqWk/TEQHhQ8hCiBCsOZ3R55MhdBcX6I
TQs2Gmp/bmrkwL4Z/2tGgdhGr5EPOiUUJUjuriijJDy83ZcFejsXgK1fmTuVzJYyr+DnQX86+EvI
ghfqVAWcFVZ8e/kfs5TksJUAziqbT92SNsxxkesX76vz64TM61rwxWMExRvzmot23jrlaVtD3U66
g+8k/oVTeGZQaXSymzlHAec0Gs7m9qswt/e7tENEkl+gx5hDCnGuWvTSZUc3BRRCfwWE0gTj+MhW
ZNLrmFym/v4HSjw8jM6/0UHxy7OBgf8rT9jULoTcNL05Mg1yilJtnaz6q4p0Rta8UpeaW+897DJt
5dUyStL7D3f7FGNF3QpUQFYHm6SeZP0CLzI7NqqpP2hZxaL1Wre6TdaSo8ZCkpgjR6zLeqWdODQA
/JyhqcXVCDD64VRka2HD1ogbFOdI3IwGgbQmovHz4E7eNgN/Zsoxv6jrVjLclXA6gl5NhTax1lvP
1+CL33UReWoNad6NE08bNRvrQzqOYdxRk0BDfZduEgOnOe7XU/7U1ALgddNcMRgTwIn4B97nN0h7
Or3tUuQZ6HO5/orfu+ET03cLqLp0gtuXFXPadSX/K5UZI8E/Icpc/F3NO2CRCRlpFiKY2CQrxmKx
V58zBYZC3isqwbZpa5uHQ/lmSMCxqCMSR7HIXYcCu6s+Hd9oLEfvEpxISQ/Rn0lavc5HsuvfwIep
8ueDUYiejn+5XoC9U7hsI1xUZkTL+CNIVQtYMFfAU8HoJ4M2pEEewHyo8Ir7Qio8DiPvAmvVl7BF
fACP5bI4opUQ+jmw6pJCwkEyYUe7RYBhh+41JKsn4zLPjSQY7TZNPk2gYzqzW4nzz883Uk43ExDs
JYVNU2d2PGyQXsL1DmsFQHK+a5/feaw2xLHm9X2LjcR17nRCnpxjYHwHdAD6GzgfxOqGRjuwkOjw
g1ClZFJGNGnWg2XfGZQKdB0FwHQr8XfnFHaXIyI+EhtnWXIqikQN/sJ3KElTXcGSI6FfXzrk6Y5F
RuCK9PklWczjYjEamo2H0heYoNq5E/6JHIYjSNxy2WGCXvZwOyuBkr6afGmbJxX0FKYVwG3uK3pD
YjscO/+xu7NWMF7AwOJONQa4NC0O1LA3axeorqQUPIMWMB/SACBn24E2oXYOAuf1kur/0czY5Tj9
lOIp7h2IPyItdVxGMZl2AwRcxZA15yRvZQ9A73AQw3GJR152aoRWSBRFlAYMeVm64x6nIqFxA3B9
w0C/ox8/3zdcKG/zAxCa/7MXaUdTBPtcirhFfNcWfD8ndi0vjKZa9m2/hrbxwpT0kVFHYExQD4p4
3yAMYy9/4KjwiP4tylgKJHvZTDtguSSR/g+KoyrVn6DFyPTxkqaoYV5yjZEzx3jd/kyrwGQbirsT
7ydxwU31lXVxNnDRivHkcTNFP6wzQt+M8ChjO/25Gd8Hnf5qzG82oNknk6OeagDk+Korp2XwicsF
VT3dRZqhbZyhq9UsOsGY52J8vY9ooGt3A4582XBq5RaNuTZSxqqyo5EuNE0jy5SYiJBw2YhTFxIA
clKYNKlLiYCVmQiLHrXmdCAaLUFrPdVhiDDJUkxnoZ1e8nZEcN5XRbscS9PzYaI9oRekByzcjH0s
/X/F6Iposg0ya0PkavpyPtfvbYno6EbYTFkJBiFBupREYhn203wtDN+RFzOOsaaY47Qf16OBthSp
e9ahIxsbblfu6S6uV2sTogD/CLjezLRZIgS8y/Lf1BjfBq0LsAh8tFM+F3PU9Gl/AXrd0TC9/+RC
VcsPfczB/mJ/gGZtLkCyhmNXn8i0jvMmT04LQ7SxPyNTrrdFCKzjLu5MlSNBIr2rU8HJsNYCOG8N
fjSHS+R3lUeoDWL8lUqOa/BJgRqnUPfynZpITuB3QpXyu4rI0SL3i6o28nJg1g2Z+0pWybuerUwc
VVsmWNO7NOz0uQ305A7cajrlnuRtdEegErEDqlOUg+ZD81satc6q3ZVKCHdC5B/VbBfmwIPvwChK
iVm9yLChkYl/8M1JZJ4t1nQF8Njf5WnqoOHXciNe4nW/XSL2HC5H9gSQS7hzq2JUFUdajv7DL45A
nEDa6d3Er7dc4YtT45VgF6x9XrC069HlS8y4JQI47vGVFr9IgINU1IzRWukr2DHSbTz5694povpr
1ZxtsGI0H70yrWjfQmxAxXLP9l0AxL57vsEMz9j4aHwvXICIhtx3HDLbBnuu+84DUZ4LMgQc9cde
RoGCGNtIVTBxaKvI2+pfXxKRLzf5RL/FBtMAEiYe300TCi3qh5zo7c/28MrwUO1jimkCKDxKuuHz
lev7a4vmTCtM3Sr899iWdtyhw3HKK7C7gIf+s64+5a8jGtjYIJLYBnK+kswndipWGFpKDH3BJJY/
gTx4ZSvucbeOaASuIdg86oALgXQzdvF8HJ4BxjDUM2HDPkW0+TPLEa4vOrXGxyxhM/lriZJBgwBR
iJ1NveRPwOSBQmJzr1Gs3K4wrHK/eScox/1McUqRa/6L3NzdSpaym04oIUX0kQJLl6F00iNZm61H
a5RTiGH2hpG4SVHj4t2XGEkFY8a9O3+C85r/23Om0jzm6fefyVEtbn8eFhaU//FtLNXMd+Lj1Q1w
SXBagFFfsyEOs//28fqBnwPCZMCoyhT79G/R3q6smkXcI5kNpHL/ecCuUc+8dMHzI8n46X407YnR
mHFtox+PpWcvv79jwHlTOERhCq8FbH4AX6zxCrrTgwWFjkp50xfSovVnvYklDxx/KoSlO56svBeK
h7h8p8tyXTxZamqlrbg4IvCQ39+JUkkBKXgSBt/LIvtiJVPRLQxk0ITIwmLtNDi/bQSNgWyF1eZv
GuSm2ePONF2Dytzs8HDcs2G+Kdw0V2PsYIIycKQKKdqGeYfID3VcKfU+DV46YoagWx7zStCLPkeY
/M8zYhJePksZOphv2GyPhW4zuRsTBjNfYEePyYiFKw==
`protect end_protected
