`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
UoTPQXuHoKEsfO+EqpCTw+/lSHISN8YTRluKlcoGuRJSMR3JvkpfZvb5HACvk+zj378eNmgfpl/T
mOT3pktjK8chkd/4/PWByj6WNARenJyiEFoxIMvT813jzBrsdwJXAXm2d2bmOcWuey2QkfZBMfvC
kfXtgzEHWuko08GtqffoHSwTlbQmHQNQBJrqots33uoFC0WtNTCO6yS1y/DayC+qUMK9g18upHLi
Yd+FdI+4wwdGNjzBRNLa9JEr4t9CmJqDgZBipjZzYlPXx4Wz5g6Vp2e4J92spm+pJQczXp+E7kF9
NsZxXeMQc+BifXxbyq096ytSTnYjG1WMVs1y7g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="EzGVEqBK1jBK0KhMTLLTVbgpP69wmUc+WRVwNomx07g="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 183456)
`protect data_block
CiS5BQ+C8ZJb5QVUaPB6gRkOdMHcmXrzMG5UNMjFgfZuWGFIotqJ5jUUF/DbvDJRl0NMA/VG/fLv
m7IqN32OaGNXr4wIq5dZy7mkV1fjj7RxEyFrCSrakF7WpYcAnV4jOa+2uUeaXu6ka+a/ksWR33a0
1PxE+q2/RI7wdBgora6FOwACts63WnPERCArHLyZHXFVIGgwk426yeGAmfKw3vYZtEowQTubSmt+
KkMjB+DK2Hfgp6XtAxvpkPaDEQEB4+5FQM+jVp06G0bzuaUQCwK3aryVThMi4DPVeap5KfKnjqK1
4YhOJtydXb9lSiosrWoMLYoavdK8qpWXbLK0Q0j8b2l2a2WyPw2T9/lshC50WPx4LzU50ARjq6qX
V9rrsNWvSBaq7DrcmhmqLbJnpvoACmxSU2acIj6UytUbf5tVDOAg8ny0R+qe/hGAcHPGpLLzjbSC
NWlQIA7dcvpFsZBDwWbHU+vDrWO527GBZ7Ax9IHH4rBs5fwjmGjj32G08ja2tAIB5BG1KhiywNjq
FVF2QbaSiVSFUjVW/aZafcvchu7+eRFu7+eRtJyut6AIn7aaj7tHercjRUW0vLv9sZVUxfxqE2N1
QP8ZUhp/Zu6u3/ANvViJ3hhapwRVqoIwnF7S8lksA9ZkLHBXsQM++vNPq6ccY4+8eEGAE3p7Dc1b
BE+kHeFlB/OKOjId00ekNq9S/yb331R5rfWB0nUE9rO7jcb4enSZ5Yxa2gOBehuoPO6jy0ugvTsV
d3ixyA+vDlCx79u10EF0+X2Bmc9/+mwEBkKjoONgz3M6UEwq5D3GRrrH7X4RpoKEmYqN1HqvNkGA
Z9EjnV8SU5NlUcNbeWxXiCAOwwDUcpkpRjEQLJkLpN+aMH80M1xgXdGer0L5H+B7C8SvjbVCyic0
M/JolyFjJD1AYGS0zaUUWMe9IKrCLbiM0mI+WXt6M1943zgTN7vH1l+WWy1faspzCF45fzo8wmD+
Rktf0XzdXamrohDLWlo4XVg3BtkJqFCZX4EgTBkVPle2JvP6u6/aTwX12UN4z3bvyqpwOuZ75qcW
Yhdj6umHKgT4XeJsxX8ZZ7+rdya+lYt1Sj3dsu+VN7MPHXVEs8xmkts6YPeCZ9uFDQtBwjyYRmjP
0Et6nJxxf90hRIZ3f52ptLbIthqVcPxUvVrlxd5QmCpEnmwyUG6sj0UWg1gJ10RddUzOUSOEQzXy
pmLdoz7Wk3RXzkJjQaYHgx0F3fbaMjy5Npf9trZaH8Uo49JvC9drSNsAXaJrBoHsvgD+SQhwbPhB
YmMIPvslgJ3YMRsRSvbUlqm+hdCtlrYqQdLj3CdzpfKbir83vZgrijHinwGm/C2l4y64N8vcpzAi
10gdd18xDS08n4ICf8DGlb3/Lvd0SSNXVHLWHENna5mj+YdkUrv7LoV7/Fpx4XzAg341qVnZdBxy
GxAk68B81a3L20Aosi1enyIUOsLLvBbtf/rw67WJ76MuPUTC48AecjrgJs9fcPIseo7F5XXN4NLH
/IP4vox81luCgneq0EInUSGxml1fRxtOOWpVF0vO+l5v8ui3S5fVB6cl+py99evDnoB8ytTbLxlH
anoIc5du6Y7K7g+odBj6vEVZBWW5QO2XCqKQV1skxiI8jpmz7v64k1IyNU/VN+zAhRtl1Wx/o33T
vsIq+IjpZIzl8xfVryHXfmTqIEbJR5LNwhkgR/KyMQMfwUhybQOOoCQPWBPfVIpZBNdNKAE3TILs
6PLfbH8HP3Q/lSv+Ow0eRhJDy4SGq5C1VYcD76BUuDGTEAT3qF6ZumLQQ4f4pXVbTs2wVR7MZQct
KVvtbD7NB48Id+w5VzbqWT7qdi0kA3NMsUAW+X1Rh4FCl08UWAW+SRycxc/QataF3R9Z40i4hm45
j4I9kysZh8A0McIss4Drq/MvaS9X1ak7bOZsMEvxoUz41c1cp18rFlpgSZIKz2MdQFIUqrg0Lefy
NcOXnRwdwQ4POZ+tRCvE63vRY7hiFZOBv7w3RBZAex5fVJ+rnROpPz46VWOLjtAPflkq4JDNm6v9
81YS2+BsCLbNV37a3ng1UBQyRwzu/5mKRRjW0lsUDBYVU0MA4iktaH26hgWKdtKi8ChmlKTWulvn
Fxi4LPUC9cwVPpIw+AcuobLkoEY2mt2N77BSpQMniR1QV/DCtnItL9Tc4PMwzDvZ4DIeyxES0z/u
Lg6HKwgaONBO3ZQWZYWmO+ENLmjtRf1nWcYcwwtRqZmlSyAanghNprekgoLKNoWk7R/uPpv0YDaa
PkUo/uOfrMNXWkH9xDQMIF/oMd1DkWveByiPyRCHwbaGV4aqj+RwjOZe4gMIydmz2JrHx8dsvPmk
69kwzYqXhTh4jWEfoynS2X3klf9vx1Eej8Ux0s31OfVZh8Q7why4xPlEPFW6G54KonF7ZOeHGqP0
+393eBn4kA+AUx8mvOS1xcHFFv9P93igYnhPeT8PEd+tvcERPHY/000M4lfYKA6d8eMXLmBtlTF/
qsmaB5NeNnFg9wpOK7h5wdsU9m8f2yR5OUN3UAbR7fNIxzrJ+6Vy+W6gmU/p9yDNP04RR69fEJ/b
F8tihUJg5sfbKz0DYKXJy8Rf8pSfVE2MocZwhxuUhpezFatJoDMeHi01yM1wQtUKekuNHnFXZo9I
23tPApuYfvepFLit7l7mf4t0lkg1sOBqfT3y/lp8/IXkjekE9OR2QI5/AJR5iIUa6RyvmWU4Gybc
x8Xn4kdcwDBkB7o7U2bkOGAQK8jmL/WqpFyaFtMchd9IQg3GIt8YLKav+SOtiD7tMptFB0l7vtQ1
PQsheJ4JedDgHnrNgv1c0i+VwJgVtJAEfIhjrw/UgJLUJZ1VzthiPZ6pF7J5XhVi7nFSMhIuPcCJ
WuVCtf5nFlmqLVuLeCmAlNDIQGk+YiZeEUL/RcV4AMf0ryMlEAVIvAjW1eMUbPJ0FOgtH9O67kZM
9q/k/GfQzKk3LTSYN3OIWlCtQFKFBKmfocOPRgrJEzkmLr3dZbw5S19GPO8zddiWeQcaL/ZNADl5
JDG2/9R1NmfAGx5tQZtJFQnhuTd0sTCP2AlsaahE/DbjmvwdIIKCuLXlY9ir26WRB0flo2VWgfDK
uXVDUdGDlPXtsDLUxKOiH2YbOsVd8G6ni9xF6CkODe6gDjheuv96XOLDRhblu2rc3SUVhfJcaGLT
ROUvVjxOKh3dSKkm3/h+Cxu6dn7h65M+diHYSdK0uuZVF12Xt9utyNjoOSpaUzor6z7nzPcty1Xq
mE3gEQKjAI7IfHJ8Tezwp681E78W56WP5FS/O0GqAa8iPdvQ13LrggyrWAGFe4nYBVvwzHrQtEPJ
QtPT/dRZd9EV4JCe7NvNc0Wmp0zZjKvC7GRpSnxe98rlNLQh49GpHxgDHeZLZ6gWVXc2/iXvyNm7
vsiu++NWmyrEN+IsD+KeU0Ust6pesNux9TBecZzN2rdXxtsYrsTnrw3vbp0nOelBg/MXqv7LzCDg
5jQWnesI/YJSxz6FeJnq3zVfyQB1YLqi/Bkxh5UvyjBZq2G4u1JrotGYr7JJ0dJBaVGm8JgkXx8g
YI3w5nPVJi5TPdSF5W0bKCK9+8nZ0Zos2fczl9PZsottA5uMwqA3rYeIqXTyjHw1kwxmnWw7vcEL
ObTnI+wGkDVQi86Kz2kjs6kVOZRjeb2gwy3n3HDQpktJsqG/7b+GZskNaeCclE83yt0VMisLIifl
QCmCytptFDandNnVoLzFmE1ku3VJx0PZwyMiHRitg1Oyp/ZeoMe889tuverRyI6oSvwA2xoO/4jJ
5LJE6DYCtL/HANc65JHB4EeBPkfZLYiUTi4ok1uAMUkxliIkGfISNrHO/pX+X8XxNYZQ/1VQ0Vjn
aT7S6D/IqCQSEf9HTNIIboytM5dBoqou9zDa2o5L45Z0AkK9g1OKlChNFHjMiKkVvoWXOknwb8W1
iXRQaG3myRYxp6SuUJH5Bqf9Zw2eGetu/qsbxkuGCNfZ+eUNBsSuLRDhPn6vNNol9dhEKHuEdDGy
LR2saFW8VzcQbElbqqwCeB2Z8mrnhiAgjawu8YM0aepVa/1/5IJJgcSZ1xhhpy5j1Fmxup5U/vj0
fSqja9a4GxIKm58TGcwZ5v+jxfsbsLDGjpzrnqIpEFzpZqdILxffRs39tSis2PSx+xq9DacERE2F
lkjATyolcoYDiF1LnVXplau6seRsogYjjVkSsEXMAGb5NiQ0lP1m+NY3D2CtOnIsJ5OBvuDEobDx
E5ubLuYlgCf7J74FGjR11bERjiofrLf3BY6dRFIQ2q+9QCU5npAjH44BAKkZyAqAFDQGG59YI9bg
91RuTvEr3CUB1363NVluwf4lI8MX+iLaYd0BvR34ck+S4M59lsjC6rwGax11zjlvHfd0FtQlntbt
Rl1qY78Fqygbxe3Cwjbwp2oJVgPlBxx9lcEdEU3dutIgVZUPryN+JsJPUMRrcp1BR3ZIhxxAS0wE
MBxV07ox38pbc4S4C9azG2b+JUY/GQQ6iVXR5J50OwhVM+DK/mirtBdWxkM7WTor8qE5dndH0sPb
1hbT8QsPsmfkulbGWTRwJBptD/8GGHNEUcxTkckStO3P+QBMTBSNVr0M3aaeUeCqKoVh0TEZ0YQj
bYWrG7tMesvIQnKKKbgpFNzefW+EaEnLbzv+pgFP7PwdL3Bwq031iLKje7h+4qQnviRizyb4YENt
5gjt1dDOI4Mml1iC39YrMW2qtF/EQqAYDNsYoFOrGZIq8mpZdiWSZygJuK1oaxNQDf/vPA4fUrFz
0xTOhdJx6kTpxxHYOc/4hrsX5pwvjh7DBUYb4l4N9mLnmtL92T6tXEIy8nlWxsWBylwqJtuIoWUH
MPx7PenHMWAp0l4zqA73tLsJUQ+bolMRIgdHF/u7smFkTeIpfmEm9yjH14OLm6ExkXQ4obycMBGE
OvAtz8vOajtg2RGoKi57piAvaayq12K3xLgc8qr0Yl2tHTtnjVcSAIcAlMK4VKLT2IK9T6iYrIME
P57u3EvPjbSpbdy2sQwZcHyKc1RRFturzv7cEw8IQuDuWhjpxk5Nmh3mJGrRsix7qwGNRsEmmkcj
w9+nablD7i/QCxnBwTt/MbFrZzFXlrC4c+oyknEK3NKOLivlCEebo8lapYJDdAirEvu7Ii8y9HXJ
CcZ+4tIs31eQprCyQs3JUhP9Ba5fZ8FpUshMHEbtLrDVwPD4sT75SV0CLz8EiqFZEbWKoNogQesT
rV13xW0i58sHS/7d16STGJb93rzFD91ASL17MQ7Mhpv/f6iBdFUFMrdLFzbgJ24XW9Ikq4CudtVF
EGIZcFrxPzumu+qAW2FQhJK628ieI4BVh4woj5x6Wn2BhyJL6AhC0Qhn6xXgWY1ZMVQex8Xa2/op
h/BC7ytNdeZhiBPjvpffwwcbab3ZTTACPLv1G4NotsEZMb60pKGXTMTNYONlyKC4fBrLOmgnqN8F
AI0MxrIlF1kpWUHm73zX1vWKMixzyRfUJWl05gTSnKEm87HA4J3d/1cfCtSLP2b7nLm+HASV+tQf
KRZzjETcjBmKyYgGKs5WUv485fYw/LaZqjHHQLAYxEWvw9p/BUGgar0Tkb81ugJy75LdUi6mFZ4W
Z+bnfLyk8VjBhRUgJaoOE5kS8axWBBjPOQZUz3dmtj8kUu/V6aiKGhMZARDD6FitIG8GuH1GIqMa
fJmahPz7UN7moJ5GJRtbpKApXyIR5sFmf6u5SFbnB2pyWfHQzu51uOapUVBZzErlmrCAa8WS8mqi
szqDorOHFS4xlp5C+K3UdcFMPWLCD1jOqgFmhUlMv/8FzNWdDuugGxOtQd3hypVb3RpKW4D2d/Ph
RF3+/5H4DnhowK7sVJntrYrHP6c99HiY4qufZkP8jV/AObo15e2A9iOFgKHoU5gEQQZbSm3CdK83
+SQHFyrt5vKERZKnu0vJGvQCKB9Q/11ZzGIljxHyNAzWVEjuPmya6SAGNw4cOC+IrcobY9Jx7Yga
a8LNVI+pITB5X5VhqMKBXCESxZQsLtXU2Oo43cf7HtWZhQ53kbTDNMvj+duZxtF5p4u1LRKnvWPV
neGX1g29lFarzcUXxfd+h3/9ZYbokDxbdE2b/NAh/3XE426fH7nEngxdGsYVR80g6RuBnDePw936
jzIXBrmzqbiGYeNB0AvMeGd2Zz7gX94cj5Wt4ggBjx30WYa21U7o2SsSYgLrOIDUoszWBYPStdvK
fyakkdZXXEjM+kCvyHpHLccQOnW96gJ2RvfVkleR0RwfHsqh36YGb1u1wMozI63JRmpltRo8zqEL
RRZrleph5O6+pkx8CxCH/XNnEfwvwJgR1DRiKxxBQ9+UH6cwXY56hFf+gGcEOEgsBucXTT023IaQ
HYL13Spas3OQG8ynfZj2EVxG3n4rP7/Cwa23rEXFQgyoW+PB/akSnQh4RafwH27kuIqR+xxjMZp8
nnicpR57x033RNiB4p2wwVXWQVw7IszeoN+f6zNV0FS2RUrlo3aHCKZFaKczzWdSQwoU1/YeU/wa
AZqEd5393XMVF2CuvEKLH8a8AB0hDxa3xoqUEFdUoPlLUebWIVV/4DsP5y4LRqGU7oc95ZW39dXO
qRHtX7OrulsthrUdZR9wLpxss7UMIOmUgjFaSyu5vSC2j2s5cUbCJxDPnVpwrlg2o3Gs33PdARUC
RKP0qshcTBmLB5J7SQl7/JYbkTfakmgDgJaP1jKvvm1ZLmU+bDKWd4SzBHAhc9aTp5vhldh0aH/1
bfpLX5udu3preB1YmdzC46pz5jyrW/6FcF5DOpCCF9jwYIp9LLmhRGyrLfSuWt/Imq0TOAX7r0fX
JjYTyFvcrgVowV9g4NFS8wGRD15Sp7uKGITHc8DUrBSKQdZK4tFnb5dBD05ic1NEpRZqMvqk94gi
yzGGrRa5hbRWuQNS+AB5CqmnmNBvQcesnKxneNCt+YiKz2vjGX4JPyTuEZ0Uo3j9/zsG9tluOcnF
efBYBV21pJuGeXZN6PVvZrm5GZ7565D6MopYU+s44adNeul+2wDfEpHMUQ4Fw1QOyUQ3MeluX1l5
Tc+ippHxsfPBQLJnb6O+aWA6I1AaOz5KWaHkLMdajDs08sztaWCMNYomaGTd/tGBP1cMn9Wsjy8P
BwSQhNccg2gQfst6AO4DmzchuqKvqS2b8qqDFiziaaBSy6wgJ/s3G48JZnCUDqt4K+qCYeXATmaT
Jd9q9QJWEtZJxK5hDvfk1MWPYVmps+86ynwlqG1ayoE9IAXzVD7A+qEsj39w0sHkJfUi9RGo44PB
6fpuiOyFgw1ohT0VvySfbSnM7dNDbeKC2uqS4HPAp1BUWFa1ccDCWz16+kenTUrAzSE6iwM6stMB
WsCNZIwSeq2FgszQpq3t2hesV4qD5jKkh8cAZDLOWc+tJ8ViB4yD7jNv1lloEWg9E7ulkZLGKLci
lTVYsvuI7FFCEsBbV+ygSgu1RWAzJxf2i/qT8NnQrc0g7uM+ZMxqQe7qWjJBTUh5n6863HYW9eIJ
HG/BMd+jke8m/rzGwUbXxQqn9Q9/eOH4HstdhWqWtXEZzVYjnqcU1Tv4VrJ6uU4y9DXfs7+vHcaN
yCrAKXme0ZvsxUIkChH/byUPYFYPjUJyo9vyFPdL/YYea0GY3pKLhT4ow+LAG1DfNPM3uI1/Ixx5
30Lf2s4RtgyWJ2TANHGdiT3MsuIbjrwMBrbl9Ng2u0uUUORSOrxEizTDlqqydgzKRhTBTYJDgftP
1axC/wrKqqi1AjET808yfIWK3LJiq0/9t9+JnKvvSrUpO+YSxRhdfrosKB9mG28KAb29adOQR570
gOP3hvP6CriCm8+vNFa08tZIbMwYLQTiv1pigMLlu6ef5LSv/cWsOLKSS32/20t+y0PDGCfezFHt
i7Drt9pYndyTt34Kg0gWVLHn+k212bZZ1sO4yeicfy626SyefPM8YpxX0P0NONOx7C9NiIgYUFrj
5Co6HBtR0c2+u8xEbQfFF2Te2lWh+zLUFhLswvzCh7NMMg4EkkVnmODhYqDYz1zcONndUlQPNmFE
EzxqCMx7AUxSD2e14B9c/40FmoRR49iu9dUF8m8obdxXe3rJEvGI23nOVef3FX0dcmuJtSsm3LR8
UHdp64FC7zDUKV+qnjKbeKMzqbHGR1U8sZemTI8vz6uGTMHJQ0rEIM0lRNppvG9r8URt+7/reJss
CB2tLMXcvADZSlKafF7gJYTyE5fq18Xxoxi5A0d5MMpjccisxu9EH93YixEu4ZxgEe+32IqAUI1N
rL46aHE6ZmshqI8wnpDKORu4bQ3EinOidk76y1gkjjo+CaEuSyWrxpxfaP8HZXgfzpTiXs2EciNf
43zlvc0Nw9UTMSFgLy5wOKCFSg280gu+oG3YQ2GdUkxFvnga/tJIztjM67rnA8lFz5zmBa8C1z4h
OsKOay12oqTOzNZdC5QheTss7d7bO3ybaPcuQfUBpOCWGn61UWziGhPHeaG7RSx0AngTKpWcgQgb
cUGuE1Q8Ohg0hBdORM2ETkIh/1yI6tI/eDYAkOLtmICyQR13CKtJuKqJsR4IzStF/rkqHG66d/WQ
ppBhbGPbeGvoLO5iPr3aOgkESJxxHJcqRFeYXZfONyNDRrs7M4KzXW8Zy10BvuGdH1foDpFXur3S
1qs0ZGdzt4HmxgSZCbTSTNDvF21EC9lrxhFwZRA+dluExV+cyUlpDyXS2heTsmjbA1s3WHpk1a6J
rQ194VDPrKUX791ORKAw5mbQvkSKH+LAwf7S4CZ/pMCUPAQUDIyA4McDZT5CAxI2CJLSepbNE2Nm
cIU8iJpvauj+5QSv5yvQXTZ9ZE6t7dFS8VAOz4PMQQuNgnC5mf+1ObGMDbwkOYpp42GuSiwdTTwX
cnqnPnvP7yxjniYwJyW937QUJUcPxKPhFKpKMM1kO/vKd/aGlKpLZwjIV2GLgDLWQa0MkPBEITfG
yf5k7UiC8cezvHA1UtPypmgrr2NZCeaxv3qtLU3vcEqvXCn29QrrM4QesN7SPm43seV/q3/JT+wB
ZZmQgjFnbHGWs7r6v9RhMaYDOIFUhKhhf+WLizvEvJDAqwqCO781BWkSexOZ0zrsRsSkb66S+FvG
xQM+Yx5FYAlm0MY0akw0Bios04Bd0vZ4YamAGjC7QHlFZV0/g0UcZYqgekWTHjzpXsY5qrccHp1E
1HILiykmTOC4rqJgPVIo37mC24QizQV9TuxMlfZ5eRk0jkpVYNf4aJ5fgTJKSyWYKo4C1GlJYC4D
zVRNoM+p7PSNPSOiYWF9qJedXDI8pHUXmgLhxj+Rewj6bi0o5s5A0r/wziydSUikWpaLC4huhMmP
dWVd+0QDP4CgbvMm7cWKdmXxKyU4xdDfZR1RiW9reXB4ximkfZ0OWvTJOLZfdWmdBP6DuljrAdo5
baWn99rfIDUCi9AZ6MgP3p8tyuGPsktOR7pfa3Czu1/1RpnL/2hQ7GQxK3Xq+bpiL2lA+XH/0LUV
aQKIBANMrYZ0MRXV11eKAFZDfr67R1CyHMOkoHwLsGCGMjmkKhzqejgi3DfPfmItrY3T3AzdxfvE
KVgHeAbXJtS9hk71stvzXl1BvPrHsnZsLOEPnq9W9ahd8iQP40P+/iPcCChiIUMfkEd3vxBB5D/D
EBD2X5uh1NbJKvys1IbhStGuGehYgLeTeFj1JhyG+Y9aPvPkrQLDSsD6oRfHrD5VmcuXAYBKqfJD
nLt3D2X+pf0POOpFT6pkwILcU1SyjPA8J9BJoiUIxsXjiD1JFvndMO8k/nCFHIsj4zfDKBZg24Rf
h55G9aw55wpriRusk6Ko706wfzmWfzyKh2iI7DVb8raQ5yGO5kaNu0ipbbZRn3VRivesn5xfg7XU
FBhIMIZyzWTodPFaF93KqieoBlZFEXcRlMuSNCTtk7DyjyucOGyEvYPxybZgRFuXxL9bYNy9W6hR
Ubg+At/c8iexQ1X1EFjKA5cMsb1GFhTH7pEhUJRiQcZyWa1tR3vLCiIXZ0whhAptM5dsvkp3+VJR
tFT7YP0QPaD18uyBDEdfFpIfnHnbWIEHSlLbXVKEuLGY8s65k1cYJxgapKckxwer5g5CPlusqYL4
NmxiZQp9219elGFzolaoadLN3LYPiNrbWJY8BzWNoEFSOimPclROYD0Qjh9n8tLACUJr+YGKd4xx
7hmhLCO3KsGdfEzKloIDaMJ9jjXCu2erqhHp5rPkDiO3BPdW2UWyBlV4uLayeASD/A56cXwZGTTX
qxiHir0vDqKyc/0+mHP92uZHbY7NkJfaIUZRvNzsFSANw1kPGyXB6IiNUMAbNzHW8aWiYdO+LdCL
B4XxMb98gHis5q2dUBBd7/WEsYc/ceYnNRAll1sGh9hkiZXf+hmbKYRSqOWc63kbJipF6725XtPz
c1WDg7J7FBobtWWG5By9ta77rcSJcWXPiBn5B7bS/6jZiCU/3b7nkwLOBq9y7uF7PA6JHDybMJ7X
phkkWAUq4zWPbJkQNp/5Dl7cnKiMXZLITHwITIH7lfSxLsoXMurHJ7YTZt2+zAk1jkyTa1GAzEO6
6Sg/vCurt2dJCuW+NC1h55iTVO3MUtKUlnCSq5/72ORUUJjkVBlOuly/yVGXgVEvGcGzfBfHzNzc
XfnxKPZXs6k1k9cCCyHMQMhqvW27L6YJodfhEp2rgkALtsabrzfl9OLhmLSYy7MijzbSYjgcpulG
yCpc/jBZf5nFVxUt52VM3CnzOLQ1p3y8zKLxfwn9YgCE7+tji1bmAbZlSpuIY2bJTKAjJ8k1CPBG
wI9K5M09BAddRABeQXl8junqQ09B/OX8mToGL5319qJV5tomHeG2q0z8AaEBegCG9zF+M9GP3E0X
ejiDWKZ6DttlyH/JnsAZjFIZ1VMCCw+6DBT6Xx9AK5JVv6dFG7O42w5uviBj87B5MmwQ9pZHh5JR
BN8WGex9tFcJU7f4XfvbVqHcsovLVoWbjvNH8KO0I7KWh5BgUaULTzD2uyBkd/2rgql1HIcMidUQ
laq6LlwIWwH7KYYEWFeG0wBmNlj+CeHAWjuv3UA7tiFDHRhSxD96X9C3btHTWNyOdxuuCn/EXPq3
+RLhUQ/AJDp2+CuFxM/79K+UCWLgE6rfvhYWLFU4ULopuUHj3dcnFsuxK3GKIQiAB7bU/v2j1Tq3
IQg+nivNkPt+vcLqQAF1h7aamYNUpVgV4U7zgWqorTXSjZKgkuZf8sXLGWB8sDwZX2MMX2ZuDttl
hyWPjinIxL/fsKgJOpKYWvoMBzvh5IcRzVwcgOxKsnKOhytD/jZxF/c3m0ajOD90EzTX+uLDHzJG
v5D61O0czwYYROK//o/biYnpd02Rdg+TSuuvfhsXaJgC4rO0x1VZilPt3m1P1lHoaQWKbzg8ff88
HUTl7rypXvuDwpcx9wLKArAiP+CHrZGNUV1Us7f45DK2M7ezGsjBDr6duWhDOuQS/K9EsPQCq3bu
CNHdsETLe6PAifMcsqN6u6kXJVv5PTcFSCAP8LsXHhTaXMBMgCbrf9ZR9UanccNXb1nWZWtbDg7B
3/HFXvge5vgpXBxOqIO+XvEUYEGUnJER1hvWi80NblUcjqWS7oxfDxdd0tUpM5YLjScWWLA3D3N9
l4ovtRqh0PnzV557F1cAO4mDVJXuwu0OAlXkSFnK6YhWj4ZBfrZwoiori7Z9W6sAUGl1G9o1kwdb
7h78YFWiCC0MuZN4uuv3rjM2b4E019ORqYYo8t9qu108ZzOLqf/dDzicm/aXQUWLdocEH2a7PSUP
cPFhQL8EGbRei7Ke153TPbgECjs3paEersyvzefBTl97u32pErwmf+W21FekCotoSWOdL3Dh9MEP
vsqCHszhY+3a3cN9MFMJq7ijFAwIpUN3lujXvAzzeASpz2mKauwSqmUWMUo69WtgygHJKd2S6I9Z
k7PrINmKeklz55nRRcO+o4zPb6gyeTWM/9hx9hosrio1N+t+tg2QMqgAgQr2pr+lU3kscj3x2KKB
+bIIWAcs/ZsFD1hCR+ouLcKzxQp+8wHBpWDkSClKhLNkiXfx55cjqDsTwgt7D7w85XMqKnMU8qDf
QjpWYYkrcbWqLz0ynae7TAg29o8r1howSm1t5MvBqdeBvq+XiCzLOkEGZdscyT1qSBnYWzIAnmun
vJePHkxVPzwi0i6h7RW9UIn0z2lp00JnGzAAz6fdS+T82pLL16vyx6OZ+72QViE2NpyQCOlUWsPt
+21vDDgEP9F18ndg0wjw4MUtXizK5fDMiBVxmIPf9+7/Yv4OVrgUZyevjaE+uCcHP6Y0huUgbh4L
jlBXQdi47nutJRfMcC+3vPziEWB/JkKkGprruaOzUh7IENkGLAp24oMQW4/jJKGy1Y2LPuQ/UVuq
euLz6aMAmOxt3RTiBY98x4QNaRMxtPXH2iHddEovAXJ3KsMlxspEdEx8KE1yC+nFmVJYG+Jgvgc+
bpeHBneFASeF9umv+WJ5cYpjI57zfwIe2DMaoVUgzqOS0Ii1fAy1fEGIg7SXCHzz067xAtwc5cju
Bz/R4ADc8Yr0tciEfuqapZ8zU2rhdpjZgM9jLML00r3XkK8jv8jkSnmyQYgZc+sigieLZvw4lv/D
Sj+AluxnyxBjV8Vu51F2AO/jzUa3sx2xIU96/8uJJsTfqTYN6/dDpPUXzwS2XvXwYsTL2cq/HfXe
DR8OTPYReagKQoLf84tZPdiom48iFctiWCDlhQUULj7h+Iy2IgkJjoHJRSYbmUw4RXCMbHqmsvc1
hWSchrHdpJqBz3mGNrL180qHxMK/26Ovgr8Lt+lgI8obOgGfviSYNKoHAPC4Ow0YifIrv1sD7zcA
CNJdkUGwh1bmcy4l+Z03jtthDxvXgG8cLZdGuSrxlJKsFSKmgBYHvEAmPwhZvlKRCiY0mTldBIoL
lbpHxSpb/kRSwik0PuxxFHrUGMptIHhU5o4mC5Fl+sQddK+gEzT4Gf2j3yQ7UUKRjl2XHCk5bThu
9O9NiYUEFJSBAnW+dddwhIu8CFYHvSXYxIFKAIqFuFXjkBG5ojsZIwfMxigbT2tezzcUysGsFaZK
IUz+pVjIFSl2xZBm0xAyM0F1y6YMdQTLduQ8EeXDzQ8JwI/nTL7s3Bri+87L743MoV+PHil1qeyc
ImWT5PRhN15sACidxXEH2/CP3wArQRxm+hqysH80rB2u3NjxrboSv84GVLOTswYplY/xCu0aA/tN
s+g2uy4PnvJMBAoM7UiLO3GRrYEBPG/Mgf8iC1W8ItHF3exjq+c0TArLkQpwAej6tu6a2qp2v4bt
49kBbxA5T0fB7qJiuGLXkQBDoPmcLJ+5xNiDV7NKovlL2YiiVmuDmajrYE6k1pKljxG51RUGpmNR
dkz/5LMTAENpxbjpTFtcL34T35BZ5KN+cYbd1xjd+KMtM6MskSPNS71gZ4XyiIFpNOdDhrApf0p4
h30w2oD5EWGDYzZnt2hwzy9aI9sboVeg208Tboa+OsenZAYCRZdUOU0GF8XRvmihQP8NkF6Iv/KS
dwm3Ticik65sBfblrhmzRquFvSwRfVYeB8JOvpFKCtAN0u0oqVf70QrUXqt7c3+1Iuwe//vOaDIS
Jome+YjLiJNgBL2reY0yob/K4AgWzQi+2mM1VlibIOj/shXpc84o0EYeM21s12Z/wKwgpPwHX5q7
owqvZ6bngfiuhKPpZ74iN0Ak7QildbR/rv16KhwdWd2tKCXZHKEFksjsUUXv3eZ7+uIlXS3kcOkV
vdGXbbSrn+j+1heNd6HCKckVN+ihoKtFFmQdSVRoorE5mpkGaqBvHlKS63DBV2O4gnPqBoSIJprw
KsWyGlc1oH8007tz6mH2FfZ9rxuGzG5WAG+QQ+Bhg4lJglLUGr6tanyaLXf/2VitFczibf5Ax3gV
jgnIFqoPPczj9jwlECdFomPzr2dbAGTvOq7TrHz5ZKvc7DM6PtlaEZUUOcY+QzJgk9nnGmx9Y5pR
trOSRXvx1fOG/odJCCSTEp3bl2hSWDMYK+Se7890SRz4qG7AaIEu1av0vEgjcZpXLFh88d5wszKa
MbtUT6VMOCGo1SSP3Flq2zZBrmap9AQlB1BU9E2IL6uJ/u64KfalPkQM6UnpGIKBJ8klJFxgwf+c
c6Iciti+RYAx6bkfuV0svE01ltofdjnizxpZlR3dYQpRnYEAmjrtOJH2O3/Bh/TRJhhp8ibEv8RI
3h5kAU0jPKxIwWeIVDzbmiw9X7cPWwyiujGseKTJlTXte9UTFgKBLpZtJZvMt2mnQxaXNp3p2sdb
ju4JrHwIcWSm4PK0soM/nZyM2fbwpyPCF0T+j0stVe2IygmZh+pIPej0a6ZExpNaPJ26em7H74ft
3DG1brtq4S0X0wOjEYCYY5U3keS05jukyUfsOckUPDTfCTVeiaDScGqlT03E7592QH/lKPND1Vx2
6FgG+LMLQx0j32PuRIdOXeMlVNTT7luVL7g7cuQlijacEntv7CMFeDp/2DLZmXacQLz04LiLjm/a
DlRxPENI+lKk/45CXlyaPFhZCSetp8lyoBReu8PdNgwdHUJFH3X3mvIN/Fe1Jo/k6jhTZ0FDytie
PqzASgy0Vu5uoeFXgT3O4+8fKDTUQ/KzlR7Iq65qfueSe3kQBVLSRiIhQwM2adB7Uhum8z4EH7Cz
leMxl6dvDv4tlm5LDUQGRVIsHzZXcXeW2Ftf69mRqrRMQ7EqBiIpuP7z7AxSD0sVNLAqT9xKh2BG
1esOA7q8TALqhdU8S5EJe5ewP1RW3Iv3gU+/B+33w2QWSPEFa+EwoBwrcLdkrVo2ogXPZjATAQRs
HTKQgKjITUEyYPh3JngYEhjpxc6NoVF54kR4IAkw8OyWkztAp80QDZJOJ6JVQYQrxpd9JNBfgsZF
rgYXiMilWX3kHUR/YHAFyCaIcOHlF8ZBUUmYzP7/u+3GzUb4cmXtYQYbmBBOS7fz2C9YuxuF0OI0
EBCQu6aCtPcmxJF1QYovwJtsFQ00IVBGpz14pT3SMo2UnNLYkZMSwEdnYLzlFqR/xLEZsdpXfjYC
0LLeNP+q/dOB8Sx9pYNflyo3TKDZrGpUf2+8fguVgjfvAvTIcRktImOxUL0IVH6PdCrL9pjVExla
/xmzGoKCeYEYf0ogwJyv9xzojNDQH2/5gDb62ka1MfB3Xr2vtJOlrt4KuGKD1VVA1CgDSNwoD+U5
kxebjNRyJgbkADWVorvzHaAIblJLhk75yBIRCILruRQKCInVArOitSAFI34BuOtwkjME+woTnMVc
HWLKHPNn0tv4BJ9e/HWMU433/RgWvu48J7AKT06VaUvui9UToqHSbTWlrKPp4+1pU4rNpKQ+0+/7
JfQr2IadrHvp/shckoITFpl3vjThzXfu7s279tzz9T+3rxe4hVZYg0yoUu5eGrD7Lui0iUW0lRFB
BWEQE7gUs7F34N472gVFqoctSSLyHpq7qDXjGsN/LHJZgwgaeRI6XMRtka/iDJux3saCeWVQQtm5
J5Qv6JZiVaVqjUBdMs/cq/5xSIvRyGhzVIcp9V5Eu4qioFe3msKzZE7jmcN45JuRx4vXPEVD2HN5
n28mBWvDk4OavRSquIJqNIF/F51WCVlsE438WtD9bXBpSuDjCnBPTgkJZIXIMjllXhnPqldyT7x7
oj9WsUDnvTnwq2esDKzBUBxhHjtUMX4+LSnvpL/ePrBiVan2jQ1xmLo3OxXKVDo0v91N71SsoHB9
C9ptLQVvlR6ToxgZu91Qu6bW5Nbmn7gxrYoP1keUVsDjxWlfTGO2pd+0irXbOjzDn3vg5BiGu+eI
vo2NahUmPqJm8580m8fWlGKPZAowQ2mV6dJHMBLo7c7HCSF1bY8zDq7LlKysictgDy0mFjV4MJl3
mm89/05Ln9Cdkb7cTmcubGbPSlDVf3M9IkcYQx0+AO6dp/EaqndavM5V5p+na5tDMCep22WbKTGY
6vMdCj5xVikfmV/TCSuSmzmewMO0jyRUe+/ny4zVSMmuRW1lJzPO6puRdq6525oT3/DLY1hzBiGW
mo3wZe+XIpefcBvDELF4a+dBCBnv/nHOpsSBRcJndvnMr7g7Udkg0xNUB+9tWnhNFpUZgoqHSumK
vLIc7TSqJs5lWGofeSNPJuGEXPXNmUbhYo+GLxLWFUTUkKVRYdUNhkpZpGaI/td8EHhzPalfaf3D
Tvajx3ksXG5nM5ss+Az/jzROq66H9JAlPpRkJddq9OHPVgtkd1v85KdnVKKc2YI7adwNzjjb/01b
KQve98b7ny2xJNXwMwfLirseiolDULfuJfhD4BC3DasWD5Whs2hQlap3zdYM6YapjLBVJKapT0/D
NqIstJDoI33N+kyE9drPrnaWBTYvs2LcOICzehCV1Gyb/baEFw5diSLEDPBOggYjjBtYy38fzT5j
78heTzsztbfiZJVChR1S52Qw0RpdpdWvYBlmJIzE1SjjXsw2X9zEEhkuK+FjeJwVlHH7d1LyzCpA
/QYTwOm/5rItzx8MXTgKJL9IKr1juwBvVcpQx3tgIHDAK4Hp/Fhp3IHCkAtTQk5TkFiDQxMwgno6
INObaqvnvUk/+b9PwVsZJzy9EzdfTtfznq3Fdiz0RI6885JUF0z/potMezAPTHnHeZH3vXPjoZmS
cG9kvW940O9nEdyKs+LhrruF+kmL/4pLgti7RV3vrY+uQQM4PjvXCg2KeBzonwHTlPnXREPFrZsi
2/XLk6TEjvuikgwh03GffqdXmBzaR3hTrovEAZbt+Iq5Wx30L9L5h+c04zsgZt/lRtMaIVlgN456
rT3D+PyWn5WoDfHZSedPoBZ3SXFVKtYdV52jdMnUK/+eJjktgcPpsL1Jro2qgJAneWrAgmoSEbtG
xAPCUsz1nb3RbgMxwa56NTJIwO5NN1kYNYGAEy7L3MxQmPoJVuTcV8wkv1bHB718GRSfEvt9Dub3
3tJASMc9N6bGS/DxAF97EZvo1/gk6djw2Vkh8UbU5tRY2Mp+csAi1VNBMUU545VYkN38NXAVgwYX
rrEHvo4W5Pfh7ARlb2WSeXiBf4QqwC0Fl6LWBJv7uyc9ZLCt6zDztxFFlUCaXrmeWUeRLzIsc5nF
kt1He8WrKjlAfGbRhDciAGD7cGiFVBjsjWGtk1qzZJ6FVictGi0gNwv3U1JbTITsEc4uMqbEWhjO
RVI4GHv/Nx7Hpj00tMHsvtHJvYu5cY1EkoZ8ESRvACbtCj47DcLx4NkMfTZJU/8pZYMprwL8PMGn
iCeenWeSVUJXXv9lAlwiViKq5LC8byOk1HgVyAmD9hK2dg8OwB1dbEAEno9ZTJhAlE/KpnW0kMba
PGPHsg4u66Qx4dAadBk0PjKVzxAhIAxUBYTC9FToVhFdfHbGGsJWS9S+OgYgctTOzjztViv3vsIb
HXuSQ8uxm8eBgdK6NbXn/9o3P+bKSCGvYNeZt8g3GnlLiLm4KQXDniAzgl3prUC35Z7eRvxFkHLx
96HqSUssi5BiC9yQRFKuxcBK18FQg8Xif+4meqFTADOmTW8CfFgUpWCLLoXKRqnMBuRDKZC8/9VO
88fM7uPn01vAbmd6Al+PwEoMfbrZV1ToK5bfT0EAqPseMfpaxFxjU13y32IAecgAiuOpBjXPBvTl
Uii3pb8HOP5eCDuDRY4GhjtIGAgIoQAAYon0d7qubQ82DaAOgIAncEvKfXurP21LFqN0gOQDCtB1
nS5eS4Zzf+HSTVxyfed0jIiA/0AGrns6tyU4YtdFkXru4mn/kbC6kINBnUOuKXFJFDFFqQZJe8Kw
43ow8dqkXasIuVYE+1MV7JHQE8zHe4S8T+4OBT4mYGHgJtUFXKc3FWLXXKXgk/UdveP5v8C9tlLm
lgrNjnUSKhocuFeqwSCodszLH1GIhAKYAQMTEkjJJLIt0D5etXC5TKcARlZFeUcaDRUxIznx5OcT
iGG8kkaQ9YG8MZgmzgI1wBLFmKt2KCmxW8B+puTj1y0rbSpUgOsuscilmo88kKu5YBsFyz05yaGY
AXpETx4YhHL6r0eScawA1HT7us1AOg4/jVw1tfRmv5kcc/ei4dUzgJRDVxv+1h3vybTDGKS6itw0
ni2NhftsnRAbxt2HM1EJic3g2SeaSv8Q8EXwhjiJdmz34BKpBkgv6tdRv87/9YupG92jlJUfhp/b
G7N2ZrPpL4xJ1B8sH8B5uIpo0dMPiG3cz45EvbZW9HiFJb9igO4+zrY4EmAqI++av8PXR0gxy0gW
VhWBeSEXNOFnyW0FfHu9ausHLIcuq1wAiydxnnkWl02wXSckesf2m2MpzWZBYfTOe1qISZoSd9PT
obhKUh+9PulSsOyiceozx2i9CxRw1Sn/SytX7m7DEw3lozoQ4gC6y7FCjyUBzar2KUyprMa7FhX+
Z0NBnzgRF2anGRsozZdf0Cu/vRogoxrGbSJ7fBHmBbYcsNLC86/LRaSHn5WVjcTJC+F31KAS5tAC
N4mu+up4f6f3vqjtrSp6TjA2dLRY0gbqhr6UBfUymeRtRi7vLxdN2BkCZ3H7C3A6ruN0Mr8QbRbR
0pDxsJ0XWXyH3DDkuYV9zgSY/5/AjW5TYa6WXNHazlTvfa8mFVHXZscJ2jfFWSMWAQsxhbWvrFPP
tMkwlyT6oblPcubpq7qUgeCn4ftkFbn9lDLxS+n6PvX5oYTxmmkkpNfAAQdePPVsBqFaZymdYU2R
Z/KVJ4wmn1f3QHgPkx+zQJCd3XsT8daBIHxgUufXr4+C0ajttRQOv5bYMbTSy/Qc2B6dUM3Omei6
Al3Va3uNddZ/7j9j8kUJX8SaBWG/qjK5/mh30unRk/9zN7oieCZhxxhsQNVqoIiveFOzX/MoNCKk
Q4pb4skWhb088FF7lMVF2ifCozxcxCBhAm54mQLNAiJxhiqef0oBx5vBZ/7BdyXczhZjuxKUKeht
vQxQfEpWNiLpZqeD/B2qZwi1WmKEVBip/jxLkEPX3GYw3BWBj4bCTLS8UvitWltUx6QujrpinT8U
4QHYzeXdEPr62y05jmhuIgn+LsSEFTwhlkY26atp39142P7uyD+8XZiS4nOmLNddmoEFZxzdRBEV
D2b9+HGxbw7VjNdvSuY2QyesO6jV0j15zhuyOGMkzEIzrLAgq2Vc3mSSp3evKJoCI1KQ+guY3sE8
NyAqXvUtntY2oSK5Ot1yQxqBO5B2qihPRf649EGIqxuvBAZy5obvxRwGmywnHftyoAdlcCkzNgSO
WWo0EGsCRAj+oP9rIg1pbiUFxsZOjN8SF8tSwFxaygT4QqwzbBY5F8ABjMqob1fWlb2Rw0gIYKQp
LcSvYNDJiiWN9zlTuTck8UcID/Terf0BNqzZefldgxB2pGwgUAaAAT5gTcZHlOJJGLOTQgEbmcb1
vldFn1ymt0bRt3NFCZiqKUKjxRBjtJ3zYok4gXU4m2BrBSh9pQp7B+5LGTIlOLdxoR7OtCbRoRuA
jh9FF0I/EaajU2CRC7UAUjbpBtkmYrsWNsIJ5caxxsyOz4kHzQrrPC6vtqLgMRIzthwgUK7DlYzV
2zaiZo58pKUS+QPJhYpEgP8eOYxhy8HkUco8RiCUMXpep0JiAQdIlOOXUGoHBnVtz9jacBJgxEsP
WBnX9qrB853rsk/8sVliQ5/nzXrNPn+Pxq0LbMuJI/aIih3vZd1E9RXN/uREk/x7SXIcbgBsvBOT
j+Edp6pS3DEehBM2Amn23RDom6DP/+xujUpD9Gq19watU7vS/fHSBNA1iVRn3G8Gx1xZGhAWKdGc
OyGTiiUniNK9v1xkLgCVM03LhUZSaNkNkn85/bShB/pB6qyCC180aHE726JpnzsZg10lePI/e90q
q6A+fQdW0ME8RB2aa5QFoqDUdB/A7s3k3j+iyjCXlq0mub3LJlhy0PsXxtWYA/5sJgqqFSMvZzc4
2/Zwdj4fLfV0jb/9laW/NzHtvSsudBzHsDbOO3Jkr3JkeVJ1VqZ5lbbVIsWEy3uNQOzCnw3J7f/R
RPaeXzi2YAsB59ItEGZ+WVViIhgHve7SA/ePx2hALn5ndPBER1y1ngMWOllbjeBfw3s0JW+XJvwK
V4AVbdKfiV12NMfewm2EBa3eqecKIDp/b0ydruDUBrA8Z0ShBt1Hhktt84NoLfREioinMrhnQYo7
ZEV5QgVqyN5RuxYeeyxY/mL0mrnonaCfia6EWYi2fV2XVNwrW9AYFHgd4sXMcFETJtnUUzf6Xy4n
sIBwR/5+lYf+mDamMS+pu9XsvRgNSnnG56LY8YBcwZYIsHLL607Lig7FejJw137cE6I0MaOneY6S
oafKxmwzES027o2Xrr7qJSp5fLDYQlxGZzBcEYD0bQmdeGSXMoigEUIRHnSazZtXUyojXrq9+4yg
H+lRq7lgNeI/1YrCK0z0bjFg60zmA9O9Z1U/cVr9xEjT2mQhjrvIBURS915utFivn7LWM6jVMO0S
RaSJLqrYd/yuP3LPQWh/HUoCpDhX2CL6o3lM0wHbbMfOawyMEtLukKWnMhcqT+pfE8YTdH11OHkr
F9HQgtP78G5hCRAJ/0H3OyQUcFE/3QiyLRYfQs/aQq/l9X8xjNvhGBhim/qMCnsz+Ck2OcJIV0HX
Zy/BPYiHxE/hfccksO6JokEICBzmqV3FSW+s6YbJfHr4/0FF8xNIBKNjyJGrmEvMakG1xLYV/tjC
bQNfw6R93Q8yNk2+PnJ49/AMpAQj8lNZl4+k77kmihv9QIlBkC1Mb+J5GeBeZVIrEx5RLLJE6HKz
snHUepxWTAfDN5MLb1a63NWYRGE8+HeBJKi6PC43r5NoHiDUFgu133qy0D85/0m6O7HkKznBjgbz
GRkri6nFcoWPZ/wgvwPZKznmylVTvOxWLL45QRYIptymaMBxZ6aU9mPbt58NDotaw2vaylyPjTix
LwF2PBVaMmLR+84S+Nxc5iRPZpyCC7ZnaL12t9o3ahN5UC0o5aQ6QqtArdR2LSdhrRsSHscEaJT/
yMTGlOmNWhYV7Qz8r0HjV7ytUI7dfzpJIj4cFn5K9HCEnx9eKQb7IlA2gix7iKJz+9HYKHpdwmNN
/xKRiseeBZpmQNr1HtmC6aqS8GQYdrvRZfROGMokQES9arknCi5m5Q0OHdN4yFq1qEcleV8Gs+Wt
L5d+srju5TRhssKzDZrSHF0o5aDR/IbuFZGbgJtK+jJO3Suh6jdkvfjCCBS0xnEdM6QJzHx3Ub6N
QfS2tUzbhIR7b/cOOM8aW8qWki5xunkOwqsLV1H/GDLTCtMTTNwTZlyKN2XadvT1oJUNu9ng02HQ
nXKBLHWY12WVdOOp3XVgHZ+RDcl5XrPfVBCVD+YiJRg7llU45cb6H8FmEFyQfq5HSVQ2GHYgG8mv
d9ElnIjgUDOjL4TX8KAlZo6pBhN6NUwgEfF/2MQmq6aIloNvoFemB/vTghY1n+s4N5PAiRGJ7scC
r6h9BPuw1QNBkY/APcVe+V7w6qCM7zKOXPMdqXfxN193+93dZMGXuIuOoPxekIKbl0kZXJOXFJsd
OyYnZL/T0UQbzt/2Jz1w9rnSePFKkBpC/Vjs5SNt2TJk0XtQaO8IEbUn5E3+Iptpd2wGJN72o1Et
g+ERMsKaxUUAjzsjNY3T0XbFblA4Dqhcgr33yF+GNVKdtjMA9Nl19MsdhusVSKWub67VCF7oGf8/
OdRA4qTFkzSYTrEFoHf2llO2yS6ptH/YwRz6FkijUibUKamUxgQRMKCcPSC7DugKj5yk7+H3OoP1
Tjbt5S9eOajKCBSEybXT8+mc705OBbvPUXo/8PxZO5kLT5uXGkHR612kjhdfy5EeAFrymq6/ISoQ
jfOsmsomIWVyU1KFv1cT6X429or3hrIRUmbIRRJYwMyJzq2WEjSgaJd5sUDLA4zt+H2ePmEpiXGu
zR5gA36hK9HOr9qhFUT6xmlRBks4uXD52yY9fxpv01+W8tK4I6NmU1B6dbEQ6QH5ts7648dmvkUe
/LEOMHT2G1rfUs+T2hNOcJP0EWpMaZOGmosatzhqUHl7Jk7uk0iOPVXqHCF2E3pk/dbV09GS1G2s
IUmvPNlLXoYW9Eaf1w+UGhW+4TKanYyw73/YG+a5HBP3ekYuO6Em5gddVHMtIrDr/tKj1rqgixES
nF5OoDoRzOo4ElDyJLgqOTet0zwNb63qyVq/tuUR1lOdJNX3JMLtb1N7Y0Mjb8+zjYTNsCRbVClw
FXwucDybdwj/EC5lnfB0swwHfpOTxw5/aTkUJde+YSpVuhY11VWi4y7FCfFX1CflHM57XfLq2Lrc
vnti08UnDck8WLNhi+vxcZ6Az/yeGt2tbaDE2DFRLOYuiIGRv+UblX1Svu6iXpN8W9eRu5m8zozj
uz+gy8vKsPB1KZrbDooCsul/96dt1+PjfCHPtt2gcTaXzigCZp0hRAff7vouRDlMi8Cv+EKnMrhE
W3vyADoNto31geEQqPJJP55TXZ++rVKnq6jzzjJUvAAtmtWrgnID8WAWXJXenT1MDNWtsTePMdPU
1LYlyJ53EUvh1v+5GQ9+eNL7p3luGLAMX1VSYvVZl3U0SLvoo4+jWcrYoF3QT9UwazE9OKfE2dd3
I5s7yQ+p4ng3CUPCm1kmTL9Dr1tPiw+B+JqNuw0HP39lH5A6HaLY2KEHfjBURrhOUnIHjcrL4A7f
6b1EtxP3WgWI99hbK5jZ+9WisjG04Q+d0KaCwAmSM+92fcfe7X8wA0huKVuAhZULI5gKcosNWelQ
M73IWN2hxgLVq/UayHsXqFdgoeIqO4Sf+oGIEdRUaixmEdJAyQRN5/wYVuNKn0NMOQXmRoiRTu8X
kaZSgOghzFdPPW+3Oqbqsj5cktVvjBoNDNixfOKw0+HO1g0bOhffTOFBDt7emQI+4uiV0RKt5Qjf
F/2CnhDmsWJOsKNG343YxARRot8HXBQNj+ScJzsxkooQBuz5fgPR7R2ybf6E9ibqCd2J5l24gDUt
mbIC2e5BxEgaG91CosYesuA/vGjvPPk0exYbDwgfwMucQxuClO6fABIaC3tnhXjF8wH5eoToWowk
t/jTicZtn4CsnNsra74KB6PdBIduICdSFk77Dz4lNnjZWmPRXDoR5hVDwcqjG1ZdPSS3Z1DZJQ6B
SsfxyeLlWewyIjDs4gCZ9T3wfiLqQdKnl8o8YHB+4l4u88WXjzL8fSESKa6xXOlDjawA+j8gIXwc
shCJzKnrdf/587Xl2dtmTQRslm92TFFywL/bvHMe/hLQBvwln0eHPAZC3GxEj41zeB3TZtFzxEFs
SD6R5ni4Av3qKT+VUK7McQ2FVng7HNRt2pnyOpjd+0gdywA9te42AR2JoOgCBYDobu9BQMc92rAQ
3JNC/EZYOQlqSYgHJrS3+XHyheE8XQE4TaXtUeyzIX4DGmaYBpDLlsovZRYFdhtFj/V4QFA1bjDQ
yKUpH51TqG3aVO9+BE9YyQ/7l5p2HZzfLayga8+yh9yLZUmjMUNNzrsnYngarHZ20r6bEObjmJ2J
2bSB+1ePgVniTF+m+AkuGaGvvMEnrFtBXgTkYuGDVFh+zMyL0Z8/js45xF+C8CBaKPQhdVUp+bhY
lp7v4tl3FzBi7RyxWQt1nEZ/sg3x33Z1VfL+UocgGmRGOic9GHC+N/rDo7ASJ451nuGcPt5tDG4l
7jNSqYQnLfVSB+KG4CpnNkbG6d5hyis6EKXMN0RjKAD4J4lf4+ZdnSavcq6uBWs8BJm2CN0Xtc6d
7VwkH/UpZT9kO2YGwz5vu13m097shGJuY6OhnNhH6SBnNl3j/lpmp095LdbJdm7aU0Pgr5UEZ64w
fD3JIhY0Dn8+qbaVD4BIIuCJfsaU49R2vAidXMokHJp3qNA+2i2zVTVs1zYwdC4GDZBcTSUJFuD7
IBAhqf4rRPR/fX3Qe8mM/Mru/s1Ri9nGGlYD04q3wOwn4Cf+uBbD+myvyXYVCBY+rDiPLA38ry5v
FNWiUqokFy4r+EM7qF8zqKejdGFrI5zxsyqXWJ/HnhtrkVynOREPY8JZGqhxHgxDM+qMV53Wyk/y
sI1tNAqVUbRvaqiH984fCZvLohpVtsALzHOO79g49yqq0x0PgJrsyagw2Mz5NHJqfeM056LYcjAV
HnlXYonE76y5JogGTw5ulL0MMn/+PJbCjzh0Sl06DQmR79xQIeu7lFu/2kDuaUFjAyVIpmMiwGk9
Jht6Nph+JtnTYTHFtD6RVnWUar8m5m0ST0PCA214BQmMVnaVTY35IXme3rfrnWaKdnyxzpbFt0eZ
0Qz85rOr6Lykvcb8EuIF3PX+/ZWHacbulAx/TGiAWT75TQONJefDv/eb0pHwLFGl2GtIE6ByfWXS
t34KPPCeWzjqK0ldycXuDdKIOtK/mEFXXNtgmp7VZtg1R7lR/sNHPjxNHuSxlK9jb19xWRbn86BH
BT17jydZAXOsSB7X2SjPaClJSLWwshxCd4GaCVIZucMa2549URCgo+nTQU/sd9AmjptPEDTSSXoB
yghVjHpHuJ6kMGwefu1CSzWqEOw+4CDOMq11PP6td5sAaYLRuEEDLMVhzBH2cAF0pgeJd2gIQNLI
IyhKMBaVWNCn5IwlIxmSGIt8fc9izkVRn9kjFLC9WpOg95vyRzSLTqSnBS/fXll7FfANxtC5DjPU
D3NwRuY3yNGXrhM9nuu7EBTRzT2akyhbLOpln8dSXp9qxys6E0ZZJgpwvbRHET7TtObxCFN6RvwU
O3WuzabB2KlEROYm9dtlS3/E483vYosCw4uNCOmtP3T4gT8FxZS4DFQtBjoXFMyJcGhjcbSfNQuL
yzs7P/1jT5q3+VqUMCmoTFImh+EfqDp8KT8bTLdv05n7yaiKjBbEejvyzsYBUPQ43dxWEjxOHBQQ
RZ4b7YS2NftLzRHXo4HMCCaklOskxuhvEL9DCIGM4pWdNbFDZ1mWXokgyoxi2fvI2e0Hz9UORtlp
MDF42R21z0mZ5kmRLvqG/nBWwILQhLG6LvWOHU3HdXC2lvgFVXPUTAWY2iMWKn4nS1jf+D5ggK2C
CYG5FlVEtY/o0FYl0CrwkCSCNIkf51rNosdLe6Y4K2QyfNMNZU49dDCAqtE0DvfpkTmT+dL8UjyE
fziY3+qpiZ4/JrqvRu52ijBGXqQXMrzFwQZZkS4s7dGk9vxpyTHs3kWQa929tnGqX52zgdOvMu0r
s3gi+vjIgUifn52duAsUMRfDwBlemO68gxMDunHW8FoCW3wcw9S5Id5um+zWh+AEV/YfRZhvmWmA
6DFdOf5PPkUkpe4vynpko5lVnuTo18EhbkPY3s7WQjXPscTnGmINxgczXOLEkYiaX+TqmEug57zm
U71IMigBe27WigY+TqLa30hFiBb/k59vR6PRPOD7l8alroGMXUg53cPf7lgdG/K5CkfyOxva3Udf
GrurER1cHOD+vcGMNN6EnkwN3uDWGB7PoSp8Wd0uToWpNBzrgQRFUv3WZ4AMtytE3X6b5SzLu9Kl
kV3Hs9qn6Sksj1SHypKNYFR4Vhqo7tKL/7W48vEH96uxFH99mveyHiIXz1YFkm6dBqtvwBCC63TN
FPyG6ZppiS7INuGolJQahuXi728TUGT2ysEK5rskYtOgOHqQaGb1KxmZ2ig1XD+xVRhVx8K7v9Hr
AyeZqINRE4IDyATxSECbQZ1oFhk4yEH7IgSU3hP54QRojpBJXOFdujevuKYEWS1O4ny0F/+rOBy4
dVBuJNS3396+EEdkHWJFzu6IIMQ3cEuRh8VnAXUlctd58EP1DNzM012BfT5rqgYkgdjFOc9EzToC
Mew556Jgn4ZLQY0fvqzTarqDVYGbA3/Wtn9x2b0e5t5uU5v3emo+Rwymwl5a8K0RFR93dYx6e3AD
1fkKgNsHT/pNOcKPUsC++wrmpKMYEGdf6lPXd89tAsvvbNb5PYNmg6wQMAOUDyOS7aRU5BVN0PiP
BPymi4x0iVk4mIRtvv8UNoqYbTyIPEIhc2c8oe+w2JETA0TQYaAjOtDeygCR9f7GGQaw/tUIGC6J
x02cev+HXtSp/Nbt0zSS/osWo/GIvaI3h/6P1/a2ZzjZ1bstP3jliNl7cS4/ziVSjYTiDkhGYLzk
2GYWE9BHfkWZcWV8AJqqt3o54RBWrch6rTWQduk3gsBhKhnhmV9hb3fr5bucsIDWuvNiNCF4d25f
SFPHAd+2K4QZi92dAeysV0UuJ9I7jnoDR1sKAZc9n4C5ZjIrB5kKXCc30wFNjhs5L6cgmsE3zWtB
bQ+cCwLqP7oPwlX3GPTbUww9BZpXq7aaWgSTQimcEYQI8B1yBlYAY4Rxz1y3r37U95h8JFthtv0w
eLdnLuvxILJr00vj7OFSo0JguwBcQhvtyr8mz5ymufZwTXKo24uwmpP3HJiwOaC3YJenH6Md6uUO
X/ca9nl9oE/XdNQPPKaF1cBd4so+Hnv8lyb78+1voKk8hInlmVeh1HuVxe/Z5nUUh1adiS7cSN9J
4VQSg74ikU3lH83Vhn0tBv0WyLfre5A920YgM1sDYHH7RQP0Uqqf6PSKfrRDvzDwhIu8LM3/WHIU
NqzpwzrczeZDsHWWhMWxxJKR13ND9qhPnXtfTYOv0xnSZX2cuPOYeAj/2D9sPkJQfwwO2JoP5T0B
oMittHPEixJqP0bQBYqkZCS1CuRYMazuUezVVqkjqgEGUXnEWSxjk/teqbcycJQK1bloi5qvrI2k
2od0xh/M+cLTAut8/0ojwoirFjInx4TtPojYwNxu6kgUDaYD33Q//xfk2Imooe5JKxmnxqxPP9Oq
KJoLveMJDr8yrzMaLDJFe/ozhIi8/3eAh7L4ZiJmKcDN8aFa3vY1PTxMRrF8P7l6zt7KBbYSMqk7
U81b3RuaFsPZIxdh8dSmJp4BGiruqAqwdA3OYE1XDrKXd2928cam9F7a5w2WUNjNWcJ0o1P45OCw
EPGtXaQVMrs0GmZ1gNEQ00d7vZKWoa0vijYaGt83DFSB6uDUmi8j1q+EXyPddkJDJq45aofAlnbt
c3umffuN3JO3zTPi/cNHszb7mC8gWijhxNTEp/MNwl27Nb/kXKrqjYzHoEpfRLVOdSW5yHMYItX8
Ok7yEx4hI5FuDdisKJpoPK5Igf3PFgjvYAXo6U+JyVm+2GzB4iNLO1++peGMo94jylT50vWSr0UC
KOtj50sNLDqYI91GXt3uSZo8LDDK8o788AE7R2GkY9L214bhokDDd8i963S9j9CX8TTFFRbKgLkn
QViJ4W84qRZRNeX6XSx8bckSEQDHgaaMfsLhcFtfjVSJRdO4LnqFStvGCMAhQW7eoK+mVXxMbmVY
tGkDD1qf2HHzbKPOMBHAC54IlEd2oVvaeDBuPI8ObL2UrhehsZZ0oosMBbPrdwDbFQiYt6r5kQ4d
JQi6sqD/Ra5AUH1ufipT2d3KWgmvQCw+RPsAakpnXng8wgCBTkD/d8QjMwOMN6L4dRkT24lJNBUF
1o9GlEnj9JW/QGjrmbIGpJPLuWT1pHMikLa/GbBMorlbaG2PbfihJfxsRp/ep8lEPR5RiM2A1MVT
BNXrRF6YLMEN2zv5vVWLnxPvFBzJS/P42ackX+kenBlT9vzs9qvkx5CZdAXhITYxsG4rdV2NvGK8
rTC2QTyO4WckUmWGD1fP+MKOYFQoBkyML2RixOTbaw2Mn26qr2c5sy5ny/pFsYUSJlUkyGIBLvRs
V2WZhGxWm8DKqV0i/HMCsFYhWBLa7HqPPA744PRiD/vL+gK1VqJf4ZFSQTNCOynDW+o3H29ABMRX
GX9v7gxqDH9+E3oAR2oxpNffmHjScR/Dy/HC4JskLrOfeLzg065mSTYIZPPeW1Es6kezvbtCM/Sv
AxGvf+gMpbj2stTkrZJmJMGxGbpQKEsLokuv/ejrOvQIJJNiWzwPLQnD8eMn0pP19xdNuLrKnuzn
JE9qNOQYTHqz9KdNbUv9xN/BfAYAcKS+ce0I+j9EiSX6Z62lmgxW8rH0KL9otyEXk0pZksSJFTJT
mpHv4vNkLLDlHsbpw2KtNCfLKlL+xy3lJfGUUPptwMemAupHP4qPfJDFq8ABspj0jsEIdQC0XLrf
IguJqxCxGsS7LsUEoBDxzKbvW96WwoJVQorkZT/RIq2CkJRRP97sRDKQm9sZ3EwhvCraGqBU1itg
kzWtaGUfwJqYcuCV/O+Ic7hM9lWmrKPy7FhUx320h4j9YlDU7itrpS3BOcXtRXhGcTaCmtjUJSp/
JBdhDgeRYIUHrTmCsm02ceWosjNODhJckww0bgoOzj8GK+oPtj0h0jbFZiHA481xE4kpMJoO2wvE
0fE7R7yaUHOZdy+E2YA7rFeYksfFXBSsCXNtiD/OXD/06/JK+3vD5Li25MfXKyMITXYNltoyukre
pTBwy1qdDLJUlFpMLxD/TGjQ3W/puWyZkcfP0CHfECIabB/O2w/6QSyIl88NcoqJciA70OUWkYqB
FKFsmyJ66XCVLOFbUnr1J95dtPxH9SoB7QmiY0XkyEfubiqNc1qJZQnNZ0DggfQ+yCozvfvrF8CJ
BKWe5xbp8bnqTZcNETnv8w4k6W2tIfaNmrMiMvu/9Tf/C/CBtelqOVr4bG/mS3Rd7G/QifQYaZkL
e5icZt7DY1ESTCHzWmDMyl5O3R7JzPvMZCBKc6aL6yR8euMk584rzE4eisjphSftJpAThka3JgdE
zIkG6OFrjKyX2hmn63Mu34ezuE37v+zn2KEq2Gb6q3grc5DJu6Dlmqr92tAqZY64FBZqVORA1JCd
c9ijFTGYa6ZJap9JpemlbLdCHDUT5EmpAfYnGsf0zSw47q2w8lXOpLUkvD7czZBjYblfAQ1iUwpU
fEupU2+jZdXykYFjWW1lOQjORmdVTUnu2tF8qq/tl78nIJnMJKuo9XvsjeXdEp8TAet7A4TqhPsw
SYKp1C5juzLwFrGw1Ui1DIAv29Vc4p5toEkb8eY7/M21LHFOzfz/54/hTTBNwWVOnpOk1h710x0J
Okd5uVupDarzHzatQkhOig2BoQs8h94If8XBAw50mBLoHOuFs4DIqxxZi0vF8WtOQxDqeK4kX1o4
LOoj5oCmxl76jfiH0VsF/KLGhGKZaBuZWT8f/DxE5St2NulHS5T/0Uk8Rcf6VS8WR/nJ80lTgLcF
jyDe9F8+6gD9ywMG5lniKXYJQQ4qScs+leZGyUQ02G3MF278D1cNEvgqGFpG6f1bpoWo0ZYsJn/r
7gARR+M1i69i+1JcWzyYOBe7lHLDWATYjt7c//BlEM1Cf5JglEjqeXGLc24CEu5tgtwtpeYRVDzv
hIC0rSUxi4JtAvhm5ND+Gms4pR4QPp85INefEGljWLra/W6ipUL5EgQXwTBvN0tgQtrqR7LOVIG0
rCHfBJcKXCuSvtbek6+pwfJkzv7X36locgRmTE9igIW9hdN+6mYW0e0EsU14VV5jTgh+o2Qn8B/Z
1o9s8g+YhqkA0b0B1YOVSjBFSIYidSy6KliFf8WJu2YiIi03ynTTJt6ahnYD+Bz6TR//+sSfPF0f
sn+fP71sPJ2Xf52L9mtvZNEW5oLYralWSZ6cpgiBE8j3ItiXU0Iha2JI7Q+dmpwOchTCrDZWoi4x
9tRjUVNaZzHoKGHmKlogH7Iq851Pph8sYpoRxKFh+t1h6SfROQ2naiP2nU1AyxBAlI4NSdmg3md1
OcDgwV6BKabPkRfdLGNkMQdHylQ2N1mIZBMCgrqrOrJJeCnAtyRXlzKfgidaP1C8J1jRON/2+xwo
pkGePSlWYbXXab8GX4v3FVFZTv6oUtizsilO0wzojcDgr26579sHdfJRL3qm4l/H932B/ep2xoXN
sG4HEepaW4V9Em4nFttwxaAp8bQ71IzG17XuaH30Up15lMQ2b1tIpTcvtpaNGKFSSBZfhwrNiYNr
Ozwwt6jbxfgCe0Huiuw99rV28hKOVEqf5eJIcbiliB3ywuiqYMlxwD1JFKHArON0cm+bzWOloEtd
G2rZiwml0z5eJSdR0bDuWhjG/pdRh1EnGiAbT0+Q4mx6XVKVHYQCH8GhsnTtmnrv+1Hlu6cxtcgp
dQRw1vpI7o/z5g7813c72ZjKkkQB51La9+qrbQMSInvsJb7jg88My91qAH4RpxiYZoK6gKDKXzsz
Ahx1Bnerf+4dxZQCsdUAb1py1ZNzM5xOhFMK+r8HkjNZlAzXonl8RSFWkTGO3pZ6PHgwVDBcShR5
kse+wdLDZP5oleXLkqqGdaARfe38552/lwP0bTsD0fByoffry6VcQQ45sbAvvhUupconnLF1we25
BvR4BZsGHSdoOnEx+uGz/cZ6Ja8RdkrzlwMU1LoY68zD05kHuar6o3/aJ5v2ZDkrejbxiMnWu7M0
1PaM7ZeKnjZ7j/ndaKNXx91vhc+Zb028py5r1qWpOI8bv9cmnXj+zObkYCxL2ruh11EkvfgF9OoW
vTAD/R6fj71Ybc4WIHAF7EwkrtjZRcdB3+nWzA1aiBATOEw9ljcS7lDV6dSq0bw4Khy8ZECeQwCy
9waC661md9BRWvJva9Lg4w9gTZ4F0BsFIEtUg922MjlsVCw3EZtuGb99HfSheL9nF8q1+7RodzkW
SMwRkhiN1XTN/4GttJ53STzgt7upd+28ZVRpDGkL2D+i4yEMbTrS0UV6UPMTl5mniWlj+yGfpXSo
Bk9WUj/PoWfTz5cM9Lwls1jjOjb69z4ic3wOFFVrDGIDJ5PVdU19icGZrd09QMWR83KTJ5Z4c6ZV
lopF5jd9GngRK2pXR8f1Z01TWma+/gPRLn5IAQ1SWoVeo8ehXu7AfL0DcervhYH2/U5EYGQFhx+X
Zj4/FpwoKhIKhVo0MLKaweVIgXCTaUhnleSaoLbOmaxQ5c+cdad2ZNA8M16CLriuDH00t47Ttk4T
MOUzsTjLqsQAlTpONOdqyuNj0kuzfG0HQd7FxvOxYoos6YOHChRjek64cvmKJ7R6iLp+evOlN90y
3sNXQLvW8cBYrbpKpXQDnE2UDbQboLTGLahHp1ZZtR7KLbKNEmFTOjuL8RAfxIEtHVmFp1l3DmmL
QuyZpMie97Gw7fM3bU88QeEeH2E16Hq/bEIhGB06iBh+ewEGP3Pn6TBMVaRkR5CSzs4h6Gg/oyPl
AsnOTz4HllEeBV8LDADn20bpgW3sW2KW5FVVdip0nr21JpiPkzApNPzzBaO8zHMe0Ei0i8PbM527
hF7rkE1AlnCdPSJu0WcilghZvBQJUVwzqubJvayH9Uy2U+uKR6HQvXFi4bS+XiAfhF0E6bZUPo7m
HFaPV3CrktNfqVGlquV3RP+7O6DYbnO0BTP6KCHhtpY6vLRYCJpIzdbevpJQGzKSYa+FS4NlSsLZ
CT7jeblpc3TlK/yl28RPbTUe97C6aihDxaJvrmFg1UezRbc6K7+cfqP7Ia3XkH7Obhh0YWMQLhM9
KQAA4oAsPd2Sdqs4K0ra1EHwLrP6a+e8EGpDvHALYMOT+YPact4bnN7vCNxqZUb6cWzqHERrbGwv
gnQrNXeDrDZCMBcyY9xIf+zQNaB3chvndizafe0nY0vxyWQUi0RWxoSZL2eal7Fo6OeEa6A9YKzo
k5VbTH6Fk/9KUo8m6l2t3oDWKIwtRDsOY8ZAU/yOoE+VFYKW5+koQ8bqKNJ3co5sQ5Ug+j+QsJqH
vKs8vMV29wHRstRml2V9SxlUf9/OCAm/YCMacI7TPaISh/Wc3AErQKQlUEhmNYcFgU/5bAFU+uzx
HpUqBjBnma6DFzre9uKaKMO8XZx0g0joOG0lAeS6q23WZIkuHRltfpkATrig+B2btche/mCZQ/k3
y/ugOQoCbeaQI0kVAPyhmc/jHd+KCak37i5le+v3as0QnPElF/8h5weVmhWT3sZcY24ZhXq1znjp
YxUIWYET4bx+A2QaVUPu68t/8RTcWEONx//zxkIIOH/AV9mAlSBvJdkOKE9urIQx8CuLhCPyIwl8
a1p5J9p4BsLpbQeCylhtEb0+BVAYhYqRpTWVYr0HjgZCYudU+y/hHF1RHq404y923R2otErkbAct
4YjdQ5SfXSHQgDMbHjMs43fhMtUTnGIM+PGvz5xB6jZ221RCYW+CgZRbMZ7Y0YKd3XlbSssbD5BX
Nwta2Cxq1xxjtrIvHywvMHl7Xd7+ClZ03TUtr4lP7uXrcWJ0PLMPs1kvmnLnxu8LnlZXQeclCXo+
h+Y8F4Gp4wGnJ5C/Qnvw5vn3TANYCz6ChN8Y9vKi6q2E5ChNMXbGupBdvFbN1SeomPg4YBtX6stE
c3kbaf94lbmVA7mFAxCCnxbSqBBCyWxDImUyb437j+KpYvwgTfNECbmyLVIJw1MuIrJBHCbpLbDF
Q3/g93NRji5PAjy10qssPzTL2TdE94zh+OkwA34m/6hQb8s3HMqFzK5dpGeVyqctMbyhZ/g9bYbp
6Fr7mdqYpBcf0tKzJzDT8gzIiL/ZU26hDgPcQRmtVPePoNltR+cKC1Bq9sp+KO6hfe7ZzZyWQL/6
HyTUfDvAqs/ljfLnO+GPtKxhsXvJsWSyiwQ1v0J6BVZEpdwLjqAmTL4sREgQkQBaCJ3GM4JYB8T8
v9UePj+qwFU+0HeN3GmgRzm3YfmMJy0hH2Sv1Ovka6baDD76td+tDzEZlU7iEZYY0pZ6NwJKOb4x
/PoYf7zTMVWv1GS1bV3/mZfW1pH5TqYt36bMdLrrUe1b+R6+GknVCZiPOd34gKoomCzpYqrmBEUH
fucdOZJCW4ft7eA1RrmxIOjdKXwWQhQ/PK72yr6nPxqcw82XXMWva+ljJtTkcsXgqhwY4M9OuoiL
pcRMt4fBoqlJKeL/zq/AorhlbLqmEveiADCYw58FDVdpBpmNW/9ASMsBhsX1a4sE4rT1+hb6UWTm
KsND+xpfI6R9h9mp9RNVGKQC+MuVHilm1eqyRjtskLG8n7Kmp7aVfdUrAAmHfHK4hr7qIoDnxg/H
uQcQj2OFDA0dKxiiG92VG6h9BbyPYda7VbUFpLR14WWn9wQr4ZJ3VFWHFXEO/tFDg7vQgMt9m+1R
1zRw5RheebpJSWd6z+vaIxgX4wK2aIqygh6qyDRXXPpaPfOK+KZfvsJWc+QG60xoi2qoIv2/cPAi
q3zQhtkA/K42dVlSXLo0VVLrZ7SBgaanfwvHx6fT0MYI+vyTHbJBfxV1Rf1plgP1WtpJ3sW26MmM
+0FalkOsbBTtZHMypbk2eUqTzfcZrvTNXn0WVC6x24xFp7WIgZ7d0poxPmwqn/NZgRx1rgOqT4fH
sERb2043H/fDQflazSZ6FxFIps4SCXhkM9RWgW2s0GJHzkbXaKZKVmsQlSdh9Pvu3QvXX+3NlSqc
B+MK1Fsyat+GjePsI5LfANQYo/QPO5YMxrkBXAcp88Ds07UIMLVoZfTAo+8/KLnq8SO98LUdClU+
c+TB8Gi19khwwZy4ZpE2JFIV2Bms8aTiIPCVtvwFDg1OIbU2+35nTaXNoYejdtD8iOaKlMmGcdcK
ea6fz7VRJXBa9OU+04UbnW3YjBxsp+6Vj2//LLEeiRGBxvBjHNkTSPxnY1dWDLaChFVgJK3ITm54
JbUFs7hYvMa6aoxBc5g1+0v5RQnLgq1C1hfvWFsavAfE3YNBjQqBdSXy/nQczatsC+P8bq7+pPmv
oHOFxnlY7DrKp98HFWhRoopQGcfTVM7k/DNWzlD/S79zxYqkAIj7owtK47ERjqvjaMdj7E4RjDs8
4bBdwy4ubAfdN71C4ajOVPkVImSXgtKIVaoDgiE9Y4nFXe01lx5rE3lyc8kHCXPFQ+eTHpkH9k7O
UZl1Dtp4Ub/zrr2BRoE1Xp3L+L1CYDvvWAmFhAkHbHhIbg8o1X4k58H5jY3Gnve7LLIr9kxCFjTd
jNwgDbqe9hFHpW/vxfrHop4F/2BAfKP6FLsyf6tp3YRrEuIPIXYqB8zGZuD/ygRXsxk+ODRe+Fj2
BLo/hSc9tURnPjeVSKbaWcUUbBVBEzjNAkWVPGZ/E6ubrCPUBiaG8Oqa7l1NO03A2S97DWdezRhT
kZjNcDTe3uOSbv4tx6z2UrR7UTqxcVdwjZxa8pXKNdMxF4gLZGp3adGIGue5+IjNDum8wBg/3dy/
dA+Y2PAhQHNQfq4ztzqixuivk3MTg7suthSXHkZqOVZea9/tS3xYFxurF2GT3Ira2cvu/i3MEWBL
9aQwP2TInI4CKntRkDIuKdWli6SQI6eqnOuKmIYqldidbgl+F7CNB3BQUEE7M3E1q62c9YGSunuP
Ri+NpmFQidJM1xvZgL8400U7vy10dL4UsFBjS0sF0y8gvZtx7a32UZJsKa88JOoxPZS2vHfXxp/i
yliUG9dfEBUNCLRvnGzGAufzK39cyz4JVkFh6vW1gvrcUk8YjmpG49R2EQohgkTzdb/F0sVmk1aW
vbYAOzZ64bqepz8byeJIx4d0f+v+xCSemlsH2ARxU++hI7/75ZKoODt3PxEHnVbHrxn2Y0uiefmC
NtZ8NCiz3Vn1G8vtkEeLvCcb0Y1/GoNSS74SQbcmpIyBSGlyDUKMckdGhEtlZI+D9s3z9Cd9nclG
jU27wA0EwGX1d42IT2CcrizWmuDFLIBOcqcVdeU9vPhX0o9hDvl9ymbCyvhqicnc+uQPPDdA8eaT
js6/IrO83/dY0a4vjDjW6A8AhQrMRZXhIIZKT9LlY5fdiQVIQCNCnUi1W4nVVlSezGuFa1HLJFcB
RBdKJqaIQxRBYrkIc/P6kPc5+tjb/ezXQxjyuy9l/hO+wIEwj6xmxwUAFRhOgRbYYpaf0pk9EonA
BFsRf8/WQHLESR2A7RBW6dx1v7Lj6N5UOln9iu+cPArjioGPs7FlVtq1hFQeeS3Uf1mlD6pNg+Qx
fnQDIj8yD3quKYtEXDEoRKkvAAMGGN/bYofjqwsCfpav5EqC5lmDijdjcyQmuLIRnT7hg1zZ5cnq
xjdFHPLxLS+A9AKW4HOOUP10qtzt+T9Cx41f3GYqesaOg3+3a6gWVGryQGrD8GCwKJhYQOcK29H9
ge9BMtJoV3AOUwpcFdGbGwtrrxS7T0O6s/0hmUD58PNHau1ifq2mxgyn5fbfaqfXfYpQw+MGjVR7
GIuO0xojVo0L8LEyE4U9VUI6lJxu9DJfUX6y65hLej5pos5CCJKwHPPhjqi3YuqjlIGXaiHI8Q7/
msCpzDkGxCk2R8LnWqeGDEmFPy3Lj/jw1XMq2yVAh8WZoJOJZbm+mBlQk7flpDMs4gJGSLetnecY
jXXm0iEs5u0U4PwmarKsVCPTYyJetb1/bD1aZ03td84cazPu0YFM3fenZK3XUh8IMALiUuEseJnM
UBAHdpIC/tPaFF7AZS460h5tQl49ybTxKInTL7BTK9WifqBE3PXIKHKaUaKU+/MGnmvD3pkXLJdK
2nLqoaWYd4EmKeJnRWMvC4TGoTfAHSeGL/yA2lDxI4pQWAthPil+GL8lStSzElF8aWcXOyQwuoxO
DyoRSfuK0z3ByXJsVcePPCiikIbZMecSVUTaWQ5+uX7NZg3VHgJuj2iDkeJcAmVbK2FDJuGHru6J
2pkVw6rPDT1deZVzxdNQxiarOPdnW1V2OMWGMO/ZeDlwkdOv0ENRFdCw4egM9swuvLGmwDU0YOHx
oBf1i465uXfDEpETdvjHOrKGdV3P802JrvSGjLAXiQO8R2xmFJToiZjSQiBc/cG1P59j3BhXY0f2
oHJWADt2kSEsUH4h55NdnOiMu94zM5xG9T5e2LVodsRV7Im9XvmqTUL2cbKFtvPnXQVZ2/ovGfuE
ahTlqdva5JSUgk+5e4VGsUoz3VqhIRsGlkGcN4UvxPruVzgjtCF0YpKFA3USBI9mv/wBdwVWp62d
iXUKtIPhnX8chuwWBMEJuZv4/cOMBGXKJiFUv6coVpmn8UK7oAmDZYOl412Iti9rdsd7XHfcKIvg
GFVg+mNCy99eHPkO8OTwY3r1/WvOBOhCHH+484B+9i4R227uFO4cei2jFNTfK6jBug45FaD8zaxx
zpg4Ho2nLDXzCGtx1KMOjak0wYi/DB2IL6v9yK80hSr6B/bAOwEZ+ogGKR6DLQHcTfXdnpyx6sOO
0Q1FkWoi9K+oAWQUL5xRvwOo9dGfTUotC5sV/g/FMzmIhbkyimhzlddIy0V7hZ5tbphnCal43yGL
KJrDDepf4qppV+fc9kxdTaYmrFVe3dnfENGvhlDnxjAOE2hxvzpdqRJrrtROK1dIBPRzzSGgLC3x
nB58AkaQSKwQdXlBgEWqBwLpqcrz6ZW5qYKjWk+OHl2tfO2edUofVIYg1PEbwatLfwHCV/XCpRZp
aVO/Tl3tEYa7Afi+GVxKIp2IB6q/h2sVxrdlBhaspJ3EEugU6hGpmvpKfIdp5FdxvOn7or64qHgg
RB3vd4KEMZPBz0nV0G3QeHEzNIj0RkKTWZW7pJfU3raFzpVPUz//uShyn1DDqlShVWuokL7DF++7
CFIYASLrQhfzn19WSUQzMt7Z5H9pxP5orR9lGh14SIUWJx7U7L2weDddc+Dn9+wJ7v+i2TVnJR6L
PpULuTWD0ucVCSYw0uAWnxHW6ia/+NMHAcvsRuQkfcR3/60hTT77/4Sap9jCHjCWj7lPMMt5NR3N
olGjLQKbATpjjYZtiLOwxyUu2lDN+8punxwv2FTVbKYYNFB6wwG1vhTeTCJ7zY99Tcc9mcwWPwK3
0QvAY9bdB+un2HZboEE2RbZWevUhwvz/IGj1E2bD72WmnxYOaW2QNQkiU4QkazWFs4HvbgHjMMvW
UdF8+MwQxJGPHEorS7wx8H68+f3Q+KtgJ+EmpF4EVK7KGpat5+5FjjnY0U99T+6Ba/G+Xu+oeBNo
Ns8x4rloccPECQTzTs4vSDLhXFjHfyYeMBzVg4g7PvYh1qgs2uVfFkWLL+zxFaIxvW+2V626pgVT
9jLR6A5JrXnjvvolNgnQ0Lsj9hqnID4lEZDG8cpoS82yccOcqez1qkIvWP3JA1qL2ThBGc/P0dst
6FmukCh41AWPDmrBjF/kdlxl6RIA7Gc/bPJvyXlWwIaa+Q3VDUwgcKbQizSO/sMJJ9+xaHVM77N3
6GWCKXlPruFxDX+n4BP9FLB5L7TC+co3woFn7wAOHOfW1fQmRRnvZyD7diJcHbnCZHqNmrTugoKL
4Mq3MD7bHLtQOgfBhkez96rhq5gYzOZNRY5/wK6eCwFRRhoSEpNO9unteI1hTBmT9mE8GfOdlyF9
lIjRdtuyYDpBNFkQ6vZ9cXbIzTQexV4wXdcl9bHhqPSl6s7Bho9X4EDE1QrceqT7i4J9U/VbZzqs
VDJzhziTCqFrVKIvm0Eg3XZt8tR8gs12U5wlXYzNzfxhzr8ds6heOCqi9mhebdEBZSUmQt+/lbLL
dfbSRFuq8IOy8c414cCVIyjsBxs5yl0BtxrQIXE8R9/My1v/GYDfpua3LW8TmAzBqp1fjw9RpQj8
lyDxFudMij3kPI4ix60mXv4x+DrNbs1TQTFRzqzeV5u30TAe7KzWn/Y2uLLo8O7axIllEisp7DlC
Ojlu8R1/01Vi16ZaF5qKjvZWuu4aiEaZFqrJFum5XtC0r/IIT/lA/xVnGY4rywbcvBsetBhxQcwa
wFTxdCW9HdokHPDtwHxabdz1qshC1HitzuskG8NqKeTGlEqAmFPldqnmOEDVXKwgV4LhExs9OxF3
ZoXs96YfC7jj3CjjlgS4NBtukyYOAYgAyDERMejW1oFM1QX6uuMAlchFoj/I7xofhXmfKr/Cyho3
oZgdRbn805uFu42kCkTJft2Z31GL13i7Y/UonY4zlACH3zCFXp0CdCWl10sXt4WOtZAye5R+CHfR
mkoeLyFpFK9jfLIMVM4TpOhUqSSiKqGlOeNXbWpZcs+sERoK9EbL7kfDrKZDPcMYBuKrHkUwBTGJ
HfpV3/1fEsmqeJySiZI/rMGongdFbKnnOa1HvbFPoyI9cQntTEnSFCOZp96smMcpyTNFYvR24kJa
ncLu2z8AOp10YqI2GJGUKm0ohh2T+2tRw8aUPvSefp0/4nb+I5IpGOqD87pNl0d5/EtAs1ZJRCze
aakMMfJov6Rl+nsgggVGJdVtNDMRCYo73PRyNCpbCKG7ia09uLKhSLjmD1/xiKrmfbVrFBnFITpZ
rFz27FXezTJgwVii+ucn7KLFsTNUYS9XdCVG/JnUk8iIKMW6o97j2s3p4wnLu4Llsf7pthAVT0gm
ZmEP/OovCEwLFCtZA3gzQz/38icNIVj3XH6gBaiJjeFz0qLa+/hncPqv96saPOdmluO+qGbCtled
rMys1sybaliaYtfNSzXKVPKy8CFWgZA65F6K70+Uze5Axs13wDOMX1C2gKjVSlT0RzGNsiF5CpYl
MMVKfQTbf27rxBOcffaBJ+v2ycx/6c8vg+2VwPmo6KtKdtjVyRT6/D+MKw0MCeW5zXvbEAfyhnYg
PmH1gz8VivnoT6Mdbh8zn+KD72FUVja8T/Em1VFt/77f5myJ/3yxaqUo7W6kucRcjsJoLae5Vp1a
M/IQTuQU05B7uuepn2ptECDPa9xlqU0pLIZnPTwmKqn5SIkCZciQKHO5/ct8WjLemgorVa7FxUfF
K9Td+VM+fpJVgZGJnEZNbN7pur3GUkwKdHaVqOodRJhOBb5wsmvhWH9zqFXc5GPm4dl3fkF4j4D9
oj8SWKyEIYjtUdh45mAZVF6/G887o/pemsP3WFQFNDESqjDoy0ghOYfnTMUizHXVxLnvw/TbDrDG
2Sh094epSkEdfQtZBa4dPM32GlnmfEt3MrM4md+2CNdhHcFxQ5S9eqHWJyBLIT35vBD3/5c4ccBq
iD9b1Q8Gj6jsmrlw0cwJ/BWd5DQtrRycrWSL57jAJaNNUmcDxTJ98zIor5rKTnf7eFgZl1gG7t3D
oph1IVh+CJt1p7cqnFIPF54IF1yr+Qh+Ku6d1swwpV1q1npDL+ToIploURxrnsnupqFBNXoz966k
R3BIcJ8vn5vTnoFx+KFHzWDQeJXMVZZu7oejCBRe9oej9uyR5PMikLdQxrEpGVYSdDGbsenhS6t9
3ySLO6Xfwc2/FVgQwJ2JWm9CUrg7HL8r0pJQknRMKQyDPxO+vAMxlI6nIvuApkfYgFhSRsOH0G+z
FtOLrV3pEN+u0HW8aA7fxdF+/O7Ann4IEFJBEyRCVERIFeP27lBN8UqZx54I6fvOXpy5S2DAOdsc
WleU+AWYWbb+jDK/1W1zQtUI9nNc7JrhgzPaIvVgYEH5aB+vZbwoUi/2qqaKNK1Fs7XF6e6UzACU
dkVA2PZ+I/ccBQZPru8cfET9wA44cMnvb8Ga+788J72iaD5NMJH+qc2ozEzG6wAdQivjj28LaX/V
NC3JCG9uvfHP3bB7yb7ilavi/QDT2zoBRioI97FI9WjhhV6WvGTH3+f6nPAT/AFRNqAneu89CxiD
kMe8wc+jRc4DYcWPN5zXc6seHl/0UDtuhBLOxG+dFlermlR2HHVCRCjCMhMnF6a7RSFdDfPTwwfG
WRFd932bjJPnompiRJJ6i87cj/1x1m+9TY8X0ehZS17gkmC5MmxtWUN+eh0/MthzjR4+hL5qmfXp
GvAO5w7ydgsNjJlHHymFl//Bb/V9ojDSUi5RUDvwWTjRqYhxxW5QX/AD54vls/DENZSun7XnlUPP
nkY8HP9c4B9q1jtOmbM3mG2KsYaXgyr5+2m0YsNUzXdsNk107NM279My0SyxXQr+ZQq44E1eTbGi
5vKnkiZtQD5s3zZ/MIkh2amsrKPG4bZF3H4N2sS2IcV+U3ZDypGT50jJP67021Prv9aZ874d+SRd
SNq9vCL1GKqSq1AVtU/JInUgZ+H0ako1CaFpmNmm2CS6lEcbRRE0NGjQxoO+Vu5GQOKhTbLBFXdP
MtRvILgV6WdCVqjZvyU1wycFlDtgpcqpl0H/I5VFc6lkhVAMKetnPADSLlb1pzUB2YIo/i/E+EK0
M8WCGY/+NoUC18JmfNqBy9tsCqXpHZC9aGmWURDSl1YDO9P8eLUWzqFIFlZOfV6ZYYW/VieifOgT
FqcDQqdaFRkrleLiB+fkypXgF6IHuBu5xwHynKmy8nKWMXLdTDqEq70cfZQdwfSJektQXVcXMq7r
xhOAnXPCHpC5nU/YfY1/mt//l0AVToX3Jj5rRRAWAIHLL1PmucevZJn2/RqxaFjKNT2NIPgzLtTA
DaPj83rAmzAWO0FqRBDmqjpnOd6rM0dJ39sIzLiuf00QsvW8D033y6n7vldKTL/dSQIi5jNoBVd3
9c8dGx07XMVdTO2Xbe+FBoZI1rzV8mloPv4yYH2Jm3UyA/vGfLelVleWF2n3XOsSjlC/+5lpiu/9
PAmRjI1nD7JK+ih54B4jaXMeAzTveUQ4Ionvl7Q/nQOoGrYE5vW+InF1Zlse88YaVqjlEGdKjRMJ
wwdAkbjuAgvlQeIIbWU8+SnmPAKVsx/Ix2dWvD77o1E8CVF0Yk+D0sNVzSzWtDLdveM7B3QqvYK2
rFuszPXlgM7TI8NGlsH6w/CUIyHebaN0XMIPKgvsThijagZKjdYNg/ziDA209pNIO+JOA0unirzO
1e2oVOzNTLv/Ycy+X7uDli6hWPFWaId6L06ccHIFWuoHEp4YQfm9mdiM0ZO4IoibYjziw4FMX4d3
Ywu1napo1w58jNhzNTBbLIN4S5Njw5/0pqSP59zEDnrctojeeBdrEe8z+z+gDqZClTREHCLYcTEP
JVhgUS2Ojx04C9ynQ1frhfdzqGWXlOVlvUDZxunpYrHkcl3xjrWDtX0Hf3ee+ofwUxemlalConqa
bd0WPEcvJjGlJKsxx6/7gwKPyZPsGIDJ5vS4owzpHfBtWRTNFlC0SbnQB6i5oiLUENKId6UeRBo1
dZnnjQZQBbcjj0apL4pupehCBG+r3b133ww/YBHG2V9QXAu5vXjHaoLy+h8i6xCyaf0Y+BiA2m5y
wdfUoPfFy0k1B8+8zO2t6D3ofnncb1G6wz060b7hrrTlrf9VBw0+affyu7wZInAnzWqA7rEpVJWP
rTjmf2wdzrUw7VW/wldqdygafx6puR9fBmZ5H/LSALVrg1nxqD0g3PVIK2Ly4vM3+VE158kAirza
zsvIk6ZqppujYhV7f5Ir7brOrv5Yy6tWZKB/uAlnS0EJm5A68cAvF/mtA11gg6QhnifPjHV8dOPT
iQi9+uQfhtocNimsdHRxCMhHFTak/mvMVkYjDysGquhO5K6aKNDI41T1/dRci4rJEMY6D4oH/+sD
3/fbnfvlUtCd8w0f40nhe5pnHfzcZp2jx3t1FvwdJVqpV5d6QioFkstuHw3YHFZ9sp+z/UfR0b+d
TpwClfd4UzFPwgHIAntLq5thgF8Xd59LaLH97MPjP8HQWWmm2FEF44DnzuaM2/kML0CE5oOPrVoI
yzzvF7D0H4E1TsWA4ImbnpTcxBUMq41n33e0+K7u/C+PCP4vGl0a3Ffc+uO3EPuPsfSQP3Tuzhy4
JMsPU968O0H+GA13vVhW6SVktJLZybhSFKXiUfuOUYPPFuTUz3ZN4mzzG9ysRRXNp3pQ+Aou89Dl
CthzLi+g3Xf1oU168HNl3ag91ZwBE3JDPcDHJ90f4/bkD9dxmFU1hI758wjQLBnAkZAGPd9NTmbS
0AIk0tAhRwTZ1rCf9NVcwr4Qs8dbE5s91BLhjdwCuj53synvG7Typ7g/0EAfV6WMIrgdr3gZBsvv
3RyYQiberjUamcqzI1L7cuaxEFcqI1+7EMM9ZAY1bXod0dENZKazZLirKioeHR60jO+XYdGtFWeC
y5o731KHYIUCQo9xQhQl+9OnuQ6nmVXZwDRbVv2cLPeqJATXF/9MSOib0QWkAtFFTzEiITB0iT1M
v3XM7PMbUsiQTyWz1r7m93oJJoWSPkCGX2WLqqmLXV4q7sHuOzgLYlMrbk+HMAHzq3uTxJxbmduE
zULim1TheQ94kDUfX4Ey6aMWWxzpIgsPiP/z+0tisz1BI9KShOXJ8QzW4+JYRsQFk1/+GZ4xwXRf
YHXo6xgewizNrbX80e6ey226IHiQYEXw7fyWZmJO/48eJV1b5s8Ot6PVXVt2D5pvyVxo4a3Hfuin
fS5A/XChM8gOcnAX9/DAyzjwIEbHzBN2/upcB9ra+VBjpHLZrXaw6qKiXf5ch0AG40NWkgJknASD
y8liJnnPQA8ZLpKr+B2lqvHmxYdRl+Ge1YHzMSzf4WW+NbJTibAGAGY4S8YPpyXWV2moUDFWiES3
pYWNNxMFqAUyqRNnSVUk0WhJfClx5z1hI1LBRAe4F+KHxOck/DFTEms4IPvyM6XWYz1OUBXQfI3+
1bR0kr5QStqWLEtnqYQRtxOya60Fg914kagc6WmJ3G6am4BgEVqutfqZ1StZjMXXxqN9ts27Vnkv
ovUnnqHPwLcfQaAllYCv+kQ1NoWXIZIv0kfMu0tMbeH5j5D7t7r/i93CTentIA+JftDOeOqtXEzv
Ip8zUykSMKFQNWfKKwgT0G3w4LqB200I/p8n4/YsdAvRNUV8NofZ+bymKY2/TST9QJrpUw1/BWD0
wQdGx2K3fITfE5qbnfGtL0h9pFHwljdVZjtQpUFV5IP/20a4YMXKplIMV4JIW4QQ00dUQ8D4Jq4u
wujTqt+IYeBDA7Sj6g9yvEtFPnrHW/L3JcWPWXzgxck27DPeIB1q6PONlD0hClDBYN23PrfXQyz7
g3EhDD4PG3Pfmkf6taMh9ojSLFNcArnVMK/rGa+EJL6b2uauXhHMlEwsWsIx2Q4ur3WoRW71/ydM
11raKyuSdUqGaVv7A1to4K7KQuwm8RoSLE0ASEVxZc2dDmpLnK7CT4vQ2vBPCC7Qu+J77J7tyMy+
349/we7vCZbMAWsNhVg+VDHoYNxnFhHxbq6dcDPD578y/v3l/FYO07ln4eN7P2P0Bx2Jn2/of0DO
EPFtE62+nxs6jQHyNkRGME2Qm1hw/5E4puhihG12ewG9GPPxh73rsDQj2v70UET6EH2QtQ+FpsoS
9WF6Wia0XTSMn2aqWnsYZYXX8vU/YFPmVrPgjKgnChldZVES+AOcaxvnkPf4E1OSlNO6eUCxDICe
K568Q/4gT0qV4yIesc2zLDRiTkwrRZfdCD8h4thpQAFKFE1mA7HpixoiGRZt/pChxMJE+h0NeWOc
QilHf5rr6al1TPGOlTjxPAjH2A8IxZlBoa6hhsEd+J9ocEYbmBOn+GgKh5VOqSkdF8tVlqTHIv2M
4Iezamzcm6TPBNJmB2OTEjk3nRzfTGHyWIMQLkAuEaIJvF9NI9Ygz0Zpra5VdRreuK9WYyHh1uga
WBto7CrXz+/pWMu0ayjf/VFwNWSEWBqBrve+Ah2sTh/r/MWRIolUgwa2KLEadpVJoEGA1a7aSUsN
oI4r85fs32rrkAuruSi7Qp1oyvKUQ6EPpYfVDPmY09NeDgGo9YnLI2LqwI5IlSPGiROBmYwa3mHI
E38yY8gTHmqoRp9cQ5MiM9+kLclxF/yl7iQUxJ4O6TgY7+Zi1utPC5Bo9mAjRc3ZdOb2hyo+3iRj
8NI7vjBK54sNMfY0PodPa3QWVXhC9jNXhhkJCaGmFJwUBp5jok/+VynQS9JIrWxV1ZCPx6rubyVB
p6T0t7ttb+r/XB/Ko8Fr14FQN7eKzpK69JUMRMXQtb3xbcgiaKtBPBckzwOAPVDO2/1dCYoC/wSz
7EOhKLmM8uuXALNJtgKR4/A3N64VNUbuFk9DNE8/fBuLLN5p8GVHJU3jvq24zRAlWol/wuoGUejt
ZR0FiCyvprbliKTw4V3A1y3REMYPx1Y6yV8KEy0cIMLQfAk73dsoOVIVCD/HyPhWw/wICM++KqO1
Ou0lV63OUk5BzKvZWSexgqI2DZn+xS1WRTK6+h4/6Im2BJYD5noOg5RAb5a/28x5mEtivNFKykh+
8c6wBDnfbSkCnf6s6zmKezz6vHnaMfJHwuT7oeYBLFmnhSQSDyCtfJ47JlmMXanKXLjJCibAAKLD
/HT85HvL7nr1qisYVgS7lKKuSdG+r9thHrvBbHcNNZuM1nexlC2n9C1A3QYlcExTV5FowVsfnydH
ZVhtO49vrJ+FZ57iYZ2fE9sOiYkBfzMl6rzUkr58GyihwMjBMnuGzrnQcka6ttDgxAcbt0DgGN64
z0lLMqS4T/da7v2NonyvqW9WpSFAmevDwtS3JHMXcyxZvp/kijjsN1ElK4WQsjm50rt0tPvJ0Q8Q
YoUAEFcRGVMFDGmaEaZDz16eXNmV6Gslxr+0btJQnnyVArfVdfEubB2fn02yCc9r3BRaZUroDIfU
KV7j0Q6JNibed+pJev4TfA/ey2HwgS77JaTzfOOyoBy3Ho57gjDC9qadcYSBc/1Rt+mssqntGTzz
ye23tlAJqUq502BDEfoz1mQT2H/g/7hBKh8uyTufp5s+Obo8LZbxY3vt2I4GPuMNlw41YARnuu4D
B1OUOrNsGk1+hMip48mRLitM2lzT4wFEIG6VQUoRrK0GSx4FSiv6IAO3eMJ6IUoAkPGpnHoagI9Y
OXN9ie8lrwkpyVCS30/5nFYi6GyZ6jxNmd9VU+otjz5D3gLk8tBS9e6AZYsgGqa8k8XEB62psxf1
Wj24xGQDpqQ+0KETlyYCSAkLBqOgKShACCkrV9UcmIiadPt9rSe4GiCFB1e1JvT451X1JtCUZS/E
T/Sw1Pd279iBD29zHqCKb9HZeKGeNshjz4p/ltPE88DkGfjY5zlc1Q5UtPxbgQnjTlexlZXAsYbj
c9qQpiVkQoKAeHj8+cmN0k4JAbmXcq3H5OFRGqztrOEX1mn9xRh8po5rWpXX+dxPp834+a9gvd+v
YDnAD5jWXyyxtjJ7nFdhly0gS6n4dm1OMX3Ep65x0oH8Ctopcf3yKzrW8tpsd6jPilZqOVRXlpF6
r1kQCfPHJUc4DbTf/9r2nvD1okKj4LWbeyqn1dfSF3P8JT8k68//eQOnTaLhVlm0uunBqqtuNnsb
032+9yzAtmyaeOlrbdB16wAr3w3NzbBnZik9zH5cAWwVwn3/2tYmoR0v49/gF3AqQI4KEMJ6kkfK
YRsimTvRLrdFEKGiMEsNj8OT0W+2l1NQKnhNW7nuHZh7bIlwjNEN07JQxuvU0pNtt0GKf3daEJ6x
1X4HBg3You0ELFykgJuwbwmOuQIawOQC7zpffbEll0nt/Z7cSYkMkCLiWm8QVulP5trbmbdxiV9s
SjHJdA02XuWeDu/QLxubCAZakg5E8kQjNycAjkhKa2H7t786I3ZcwxlaF7IvKTenw/7tHgwh0oOG
vlP5QFFogcnuymCGwvERpG62cXT+XIE6vdPhEluvD+XXndcbebLhU1kL+/GjUFGvxVlS2uXgUMF6
OQvEaE2CT28We27yVZxUuvBJHtzElamoNyQpwR3f6QC1oX517VaZSzkd3NirqNE7xs6ZtG/JfsgM
aCHbE3wL2VWo3Iyv2Z4WzxF1YOGt0N5RBT9BcBh0xuUVTT2gb5H/0PNtbfw3zwtvdueEiyDBy3od
tKNFvv+FVrWkHtJGy079ozVWE0uLRqFsuZj3waAnakuQuEINrnNFYDGgVeUg9Kh91+4o5Z/k9mxE
vJou8GV7KUlLKeyyea/7hBFm+JNDaHEOJxb9hcAespzsL654m5dRwF4fiVF41udn8n5nqM/892z+
UVmlPKFL6YnaMZ4Z2EN6JiBQ47kcDmz2xGfPYEx2zFhJgKRHpLrva8usGC/sq2ku9BcFNzG4D00g
uX/2MrS+UdTtQmKFB7LAXQDCru8KDIbxNZFUPJq0V3t1pO0MwbOke/1M95u2MAtq0SeT6xLDb+tP
9Hs3W8rl4hgXTLS4H5z55L/mMb2r/fyjrrKpC64G7o0yUvfMCBp7UnAWeYH9uChQOh/M4tF2c/DD
h3C+AbaY1nmDFyd2ngFfDDOrytsLzHKIJVNqMsy8BHYYV0O2oLeU0hE5+2lBjGjEEi+oIgxtXG9C
aw+L04IJc8CLzpYeHfSrCZuSwWHMKQzMt84eEnoc/v3nMhgkF6ZlOW/36JMFCbZqLHiF8rGtP4kG
7/J0ZoMC3CnCw1h7D2aZ9duxitd++YWAgOkwMeMKJYMsk/05AdMsKsTGjoCCpMK48HpcOmggXZhE
sHJcGOqs3VqQDb2WSiyQmI0yfR0PYdkzwRsxj+SbqaBb+z3Qnl7v+LZ0A8Nzo785xbBTi8KTFMLT
K+M3DI5+nsQZfRmT3ZNnCGtZWZ0ZPgtNMrs4a7X11vkxrFTOhm2LhxM1X41O2VYPS0RDvGnlGdvH
8ZB+lyYSLj+shmQHxS36o73CJC1qARB4BDQNcFBBOkfAO8rflnHxNQxuNq8QvpQMMC7cdgtRlBqn
cGYacL4MngEmMtXMLGj+Xwx7BWJo3NJzePTeD7ryW/PsO7w76EX5o9/2MSPgqZ1eFRlQD7qve/0D
jE0nUOvnwoVOvu2aT7LnwPTh5TgxsROhs8K9mTzTUDE9eUV2b2WWGVwQwHrOCDd1ZhBn6XshCzEz
q8wNjVgcmfbce87tcfrUWf5Ks9Qh49naQMlhk6NYQdEUBcHGqrO5DZwUGJFr0rEtN6NXaZDwISMe
eIEVeVETYlhEmXUZNS8cMUOW6Ev+PddiPQCt3TMD01OTHey6d9ZGkCN1Bh0e6uFeKORgsjqkh5yd
3SWMbUUb8/2C0HdwTITcPiIQNShVoNeD8oAVHiZ7vnp5idDGYAhjUfGlsuv++6UNe4StVXMlnK6G
DJO/qwj34dsPOuVScUh9rkTSsj9t/Hlog/ReAQPc4x9Mu6ZSg8yGRuQL7cApFSbt5lc9QfiIEi4S
ao64DUznfGD6SiAmW1weVtwOKakmx+v3Z1oWW/aGh6UHqop7QAzNEApF2naEpDOteBpDKlvNbr3Y
PgDLbD/JZ+wBF8B3i3E5VRTTof+ndxSnmwmwLcSDnX8eAeYqQR7t3v/ZzVP2XzIyaq/f9basOSoD
U5+960EihHpSJW7AaIiQnimu2UqCEdc2qfW9rpCYrVV7rGu9eDl94yOtjz4CGK4VyQHUB6rXJzH7
/EYBA0v0c6idw2O1J0EoKhoEFWKcQnEQxnwzqMa+ylz7Xs4tnIlAK4SJQ17b1T5WgdUW8ScQ//tb
Ttr8Rn0I2zrt7rVTr7szr1O5rwMui+SlhhA0V1Go5kWAah69OwnVYtfiB6ArFtDc0V0K8SOadeBb
4E40HZTi5EjJBnqGQ8C6rY7U16dj3e8ify/kwzB1q8QfCat7+kCtiG5ekeFFYZv1q8BOtnokga77
Oq/eJlgZvjHCCIlcM+fR5b+MmbvixSeRH6cK/OLFdVyCufYH89OT0GKMx501pgVfndtpLMu3gy2x
NAmCEz3iVvY/EZn2zLTbcymoLddWa8Q7a363erz4XRCfc1gXEEUUI12Z+ZcwuZHQz8nIC/Kb2Ddw
qNXkww1VyEFQ9zQhxpmctu8jnAbEOBIys5q6NV2JOgK+RRYLdoSyC2lqGy88fapU2gterh8c8VCv
TettZhwkkEBe1mBtKsk9399+nospmCA6qog1MJTisAqntD8nMo8kBytzbXED/GGWYD5T97AWgNBn
5K3MhDuBCpNDXWZleLPKOxwVsNtbh5zzujae4lC337dDUHs6/smwH5DSalRz66oIMq6dTdadIqeI
fbXR4uFeg9geWSa7J8DNwA7AyliJGybNQk49A69iR+cEw1WDJQGEkbBYVlhovJ//cozwBZkE4bVB
EshakQCEk46d7LrUxki5BRqBPAA/UF+0eA0uUWZPBaN4MNBWIJLKDSlwlZmi58nQ/XjP9+qSFhrl
LX+Oz1Ao1LgFkS3g+dSPEhF4rkpEnEpMRSr4rGu1//BxNppWbPw+PdFmBoiZKhldav3zUPbjR0Y3
4d/mNWz1XuoHmcG/sSljZsnTJ2/XXAj5w1KtUB52T+m+3QtQv/Jt6PrdOx8Qf5PZ22c3UKJhOH8C
IHF8mSXL/nXqITbGmhHUL1kutIfzMj3kUjdpmUtGZ1VDbeSwHlDYVxnpV5rUGksJWcP+hCp8zGcX
XrdTI2LmL3sFFbVrvyVkvOs77iX45YTtt1tHqfTyqNClwyaxpIL5HKG0rDmYlINpAZFsaQISDu93
1y9F+vVbBYW2MHzwIcR158oz9gadLP6Mxmro5/liHnZ/0Mj85EMPuzBOvf5/y7lHFDq4sBKoJiqy
2RVS/M/pFIDElHqaTiHbGmN6pm+qkeB44727MK2qPRYHTD0IXATDr24Tq9dy62FgbJHzNQcJjT3J
xAO0cNf878FrOzi1OqL2Y60aiAzAL3w3rXEroNDtKrKMz0XAPUG2xRgcKjbYKDw2BaXAh1kXGR/H
IYavNCPfUllOi7p+6ArXdFOhNOYne7CTfqOVuQFYCt2v8Msf+LU187yrMk54xm1K84lUO46/r0yt
U4zLwYBkqRW31HlnSQKlmiuaNLAfV9fVnU/41VFkfw+TFl1vEYpMglcnPvYqV/Hgm3O25CdJy7Le
7uh/mRAEEf8cOb0NX1VngHI4QTel27Q7+Tw1PhUcKttroNn/PcGU0Ns6uirxnvm59tVlYA7K5U1H
WS3FscLLC1RpfRmdj1K2OIHjVb9OG0Yq8v4/0Tcu/RnwbH0WsMroYmazpYXxO64qpMqOrYxCxz6P
O0IzTEBWlruBM+aeIraB9D4PW+vevd5mkYj1v5nVvu/cYHCcLv3Nbt9eUSnsjg/c7cWICepUOddN
kK4+un3xJI9u1h+xsJHE1x/aJunBkTqrvHAI0tQ5B8tO4OpAJ70dZf2ZF0SffkWvEWXwLlCSDGE0
bkUAYyLxmKcTysU9k79aBazIZcEByTItaTh+NsUMjc29pWp7/zFcl/8IZnumq1Q+dmQiZfMsfZH3
IgZs10UpDBTOmJczPhoj3NZhh1p+sbTq/PwZv8HejyYDdxbTiueO+NC70dYnFtw6ZRoOXHEuZm4d
sNS/gcnReE1yFqfIThIrSgNTV7jW1gIXKp1Gw+wkEx34S92mZKSuumykFM+kf6IsCxjjkTOgLTUG
GAnpVp8DxhqtYKryMyH84razVkcY9S/pvOPHdpHw4NpdJzWyKFdhftVAQYt4RBNxub84D1N03c3c
/iboCjjONWYDoQ82qxWdAMiDXeRJhDyJ8mM+QwUxMAwvmnxN40NP8v+gGvGWH8uk4ErXkAoecwKU
TtBFSkHg4m1aR3eiHNuBlw8DT1i4Gyb+4BNnsWFtLdixA6Bms0dk0ryvSlMX3pCcvKq1Kv5URPLz
hwtkGJ4hS7HuOR6uaSzMYUFpsta56ONRvqHdGgBzsRDA1unU/FbuUawvzo9d2wJsQ0eWsVYH+Wrm
C4VLvSCxsamaZmnWhPr58tzdE93v+wOp7hs2R2kzQcZqfy2bAZRjZ1ZV3hhVhWiC2B0yyfXQOR2H
B7r20dDLYyTfWrun2WPeGSfk+aLwZ2BRlD7Nk88ZGzHOUZaOkIZZcmqiaIL0HXjxtSBCF5M0PoZG
QY/ViqFS7+yE/+l8MQSA+wtxNg5XFFS/BnINxbIyijEQucgLhv4XJShOSdy+SPN6qUaZv2eoBuQl
UMzGDab+XO+gKYmouqGsmP5IDrEPXeLnxbuYBXx0TmPfJLXKDQ88c6D5BpE5TVJc6Gn7vMdM+j8s
gOr+NLL8/hlAQOKohlmIO94YaknHMuKpm61A74f/NeNpSK5goKbVEQhzVACpvM90Ocdk0pwl//2E
wJe035XhR2iPdjz4atsH/hrON2mOozqRALRXVCzo19+8nMGhCsLtQVLlORwljX5EPOob34rGqQFs
t078mch8rBlC1giEQy36wcAqN/EFFVxQXaauG6rH4AyhBhYF/2b2huOug7J13/aRCR6r5vuHXBfv
8adWhV0/WG4jBQrmCj78WLQQcBW7nJRhWcUlNsbpklFEc55gp+KtECOgrkHmg+pxPRdQyjeyKv2r
n6vHfzXjZ/uZ7RGORBP5vZyBXpeghCjlr1SP/3t1+hsUD96ctXpSwAced1Z1JEGO23WY00QkGZ/E
q2Mp3gZoMo3ug7jyGfghrvFmxSK2OPLR+NHfkoVHHPYCkhSn4W12I3lm5IFrBtrTgCHiKOmMVqFe
+NE8XXBRM4VZYpAVbdlpbEgqDZnj3jUMuCA4V+uzsCOM8db7HHulCZLcyUbt/+DmIB/TE9TJAl8Q
HuyFqJqeFxEBaFWD9DM/JCOtJOM2rJd20A8BfL9P4RGX9TRs9juXrry6UY81T6eCDrjXjRQLnLB+
UMzj3KySPHjV8NN8YMWoVZB9SiJetVeWrCQ84Ngy1OP5vM61bJNP22pWAaTA7LgSNTdJIOOEfRJ6
rMUP+W0gysrFmfsvXkrlxxiZhQ94to6P2NQyahzxHTCEjFnGMNUOTDH2RMRrOxElIcIaqIORVw4W
y3T7YOaD+op/fAXTFo52VIhG8dPvXU8GMN8tbG4e2UIdyuCc55UpXy/Mhz8MlreFmsgqhYwkJJnz
dlsAKRYFoBbBH2na1ysiuZeSoFpDvvdOhQSMQB7DPNXznDyyVnAXmHULsxGz9bSS8UGp46D5pC0w
a/ZBMrejYoZ03Tndw1kjhHeauoB9oXHLLD7f44B/TXQSRwgi2pISAHMDb7lNiXh/7jzSVpD4mfjM
6AnfWJjLhVmefI3tEZA0Ck/mlnmmTY7kAtQ1VUNZjdfYejbJ1gQBhuACvLY9wa6xKFiGdYiaTQ5W
j2+CSkhN1OgSxCbdhJUx+rHZh5O93fc0zB+mAifgzki465PNZ4u3Kt7ws1FjI7qSXym5w/MabVRH
8Y1LbmYQxMIedTOJw08cnJzlyfcAqCyt119XL4rHRQAf68FsYwR4vMRXCGe/E2FKajOinHna7tfR
j34+Dc36BxoE26RoIcEqPRfiBQ5fZJlHTzTh3ta4tjZt41GrkVbNeCLf9KZ1wwGPGhkEXrM64vaZ
AjxZaxALY1J6juAlkfadgq2jOhxI1dXHk1THfeQBM+Cm3CloXu3TSjfXtYBeaUFO8hzYGyQNAmMF
hKP06Bx2g643uZvoBhbU46X4WBbrSuAwww8oNT5FUylom8DqCfuJzq72faQ4VQcnn22LGvfWyuMK
TDDcubEBc/PLAHS5We2HLbAIFeCdajzkmfHO7qFHhNkNxBa2c73/uogh49uaTLkDXp4wntNiRlRW
zUJYxNJBGhr5QchvVm0/CpYwjuMhmYRpj4PJS+SCn0nLwjcB3adTDWdEUA9d/k7IEFg9FfeAWZqR
uaZgrrETA7mfjMve65avhoW6vZWJGKcUXSbJOzzO/S1Vhic5n0uvgFlthaT0ipBWMrdwxU/eo28a
+x/N+EM7ACPwgw+5R8geahQHLFHcJO7ZV6f0rm7lJ99V4MxUYeD7uolzJJ1+FmY2w8PqKnvXMsq9
YOnhD9274dR1ro4UGK9YBK37nLIoCtTn8JubmdPuXDZgoIg9z35/zkPwsnhFvASnsyY1XzTRilA0
rgbFkfy0x/qVnII+MEPMQgKUXIOmvGm4mS7r3sSeRv+Gx4jztM8CSKjOKVeZdFX4ZkNytFjql2cG
jXgkyZ/92u14MgsgnZyv15SsXN0VhTRsSAZigt2sVMWhvEQqjGwH/fJb29D3JBgdCLuc4XSecahT
82hsFtCKrOWCt5sNYvch8MUqyB5fhK6jSd2PfZ6cerskavZ8Ck2PgOcqDC0tftOIdCpRBh+YLBm5
ZsWD45P6x45ryu7ZhSEvLSs1YSm1gtmajNPKl39fNIwBmL3JW/mLImFFRHrYQpMnhltU7hRs+/Sc
vAcF/24j2IprzLYmKLrN7WdVFLmlu+J2uHpO8CKnUiF/PQ4i8qy1Ho9EOWY1K+LCfQ7RJ+q5vFBj
v0WbEnw6LamJkjhML3eia6NWkSbD/nLe2dgiy9fD7Iy5a4OMmZ+AEZ+/ZiIrJZkc+PaL2ABjgLH4
jWPJq4LPuuGDo9/0rBDP0v+vbH65E1+TgaB3dQOqZUDhhoVO3qU1fDbQhAMaPxlt8g2zdp/DGLVC
GQEaM5GrWxgALDOiVrm6UZXD7W8D+4zqgK4mZx62JkGbZNuHnWPPv4aZpwkCBMs9+poqGlHC3nEU
oNgpuo1TT2Ik1Llj+LlHmKn6jHsIQo83SsiQd1U9YJr0r942WzTLqRwFo3DNKcvpPJvFPtjwu8vZ
pi19Ni4Eykgnv37psyuWc5TCPsWVDkjygDgH+kO/mjHSb2HKEm3UyNMBOZqb9eCXAvCHVnleovDf
HPMMEv4CU2WyUFrtpx0XqIlDLQLWFHgUEbGtxfdsMMXhhhkMx/WyFgf9PU0tRf46OBPadCrJ+el5
eEFAvPQNGOau30JaLJfUGVK0ZsEoIOLOagLjr48Wvvjum516ZyEWf5FN1t75LYJUCd5tb7nE7cz0
ODCnZDq32dc+mH1cpU38wiLjG/DTg5mSp3GgVPk3ksS9G9OhOU8Kjgmo+otJgQuJUShHrQm7yjml
rpURi0gZIVCKVoWEPzfo5SUCDmKkxFTEMgX5xQdF3K//0P7U4u5Oss1L1imQbwnoVx3vBorHF6F/
UJT1E8eJA/B9Q+rKbBPtepbPPh0VgR5XndJCGvFxIGTG02JKRSUkOUo4GGVHGY8kCoqDePAmhoRb
6UOItSc0E18OMBAhFfm1frqGipAKaj1p6OALETay4VStiYFA9WgPsPK4xal3yut7JRauRnEw76et
6nZccgAIObEGT84vi6RNqPRvgqVN3mPBgPF39oUwFkA7IFu+xpRWgo/PPwW9dxexDmst33Dco2tT
y5T1HcY2GVR/OyYu5nWRn/j9uPUluIGi8+bNcNCsZJdIIiwLf+bhYaiTcWJ15txUsIMITjweIRWZ
7g0ul4h+vgmH/h801P4bcp3f9DlsGpJD5p3BNuxpZ6zWsTUuMgVAsAy0ZTTxENCuyYSxHeTiQIiy
rNSIPtNLdvlgsB78SEQWtSVHtZXUddbVbd+sdlBmhfElak4tkHn50kr2itvy9FA14D0TnT85Xxml
hNLAzedM+NB0AYHRg9ozTwX/QVXAqyrbuL7wLmKfok1PMHyXcib1JceO4pc5Xpcgu6d5JsGCz27l
fEQav8CKAu2z9OsKroYltfcPLMIUkc2QAB2FJgGR2OuCOleyRxfKDqeKEiIyYjti+Kj4VEReAEl6
DYgq6bpvkOWbsLbtx50b4PiBlKTiccyu0YvPMLLqUylPZf6nBrJXvLOo01z++A9UyOyM+3qOxfpT
7K+Eo4aMlwbnvbWfNC6ybzFGLiLfji1ZRwKvT7JKDnElqGpSJfyJJzX5Nz32T5msyEjPiiN/HnhM
8sfYt62FSocwtzpbPSiCzLLZvw8XO4mBZwqUFt3WYhxU3f5eh5BENb/9LltJb8Mdv6rfzk41rQyP
vMD0fs74mx1CURg2K8fsFDx01tVLBIrpflg/uRHxRyIvdUZfRJywBoQ7FNcoCRCb9aT4IJtPDE43
cBCCTowKX0LITeSF4SK8VLpSz9qDtVwtxl9y62rd2qcmqDEcMbUbDJL/6Q+rEgUeJgqoCxK1ajKq
QO8qFn/tAJ2GCLgECwzPIJGSeDddtTsmL/vyl55PbZ84DWbqnTptmeV2ZbiP7uaiwINGMOcvNb+j
3P6RWFmT2S+mOT8ETJvolSjUosjGxW2wxm+/H4qXirdPXVIy2OQ1tzHEUkTsgYMrqiXQoOrqEnDl
rj8wPHBLoxK4voBOAto28v1V/CPEcglsPyB6QYsY+LfE14lV5UHQRkwiCpiV/w8su4q1Mivo3DXf
+Lia05w4NDSZwXoDUZQCE5+qAbkqt+tESGXOs+Cs+wQ4BWNL191Ww904/ttkuo/tDCZprXXSEFoO
NnmlhqkVH1rQvP+t4xsut/XPHZs9QhRyhF2oPmSu7lt7LaZOr2j6FJtV0PLtXRbwoRvOedfjyO2y
oHAGcIvGmkMDKEDno2U7aWt7DsYHG49t/LuueMWuxndZ9fwjT7qhj7dGoq2eWP5yDMFTBb7SzFkK
PEAqCFmPexmTayRsrO3sKuoYc5c6UxNpTx8MIvRuN/NpLCOLa1uHzR+Lp96nWekSDAnVmkBzwRbz
3FD5BF6OOkGplECKceId1LA/2jJ+qtCXnh7X7PQC7HBN1i9AMgdmHXvhP3ZV3aChPinI/NgTKCe3
BSO/RAhawOfEif6WU4EBivDsIHIOFFIr+DePD0ohPc2Cf5+k18i/KXic0iY5VxAhNIwec9GVK1tG
03vEBwqO6HM1YuRVnAWMyq6S7rI+lOTBm1Vk0NQ3TaZ3lNLzJcLv761xXjvR5WVBYwClWjjNlhCL
B2STgANYefBFwGUBH4hE/P1hMzfU3TBagLDPQNxYxX6zW4PN41sHYgOIQfPTEsWSqzN17dxjpoEs
e0yU88ZAe0zDp5fx3odqsz7VX8GWM6Z6sONWAJR5XGUs3+6mfThv4ZG7Pi7QowP3++w+F/pY5KvX
4beq5GQLgSsYxqhiRjHTx5sdOyLj0RcN5YdEJdAgvVODnZFCZxMmmX4m4jhne5TV6bU8hg23atUo
ZpJZ6aOFXnr9Y03vEnSxh7BhDBk7OGQeswFEeCPfUpNsLW0rmNWArrEIXVEa+eGIJqhVu7Z0vfRi
wk8e7SgFjFWm+zXR8vniaqJxY+EXCcA+vwQa0mXcvM5XMIYT/12vN4XyawtFrDJK2vddnNU4MxyX
9kHuCU55bt5j4bOdPqJy7667seErERrMmkAFRXVYUue3WVpSMacZl3CaAt1vc+W2jRFGrmRcgVAP
n2sLqASeLIy3nTo2eySMMsui1f5Vgy7sOcuWRHoLJWfLx81tXx0Nmz+3rLLYsbiDVfISEQEjP8YU
JoDzLvo9TOyZxLdxpUbvgGGN+56ZmcMIjunaElLWKfEwPHqRKRYS/uIidyt8q4yGfyBc5fqNZLsH
vcGO5xUlzc6V5rqB/qd/1WcnLjZ23e2C3IqrG3D6IgWMio7xMXEahvj/bKDZLQu85D58Zx7ymS8D
2PDrhJJn2BalUCsDKzpVtF9iG7KRfCLsOV4XG0enR/y+Pp5qMUmbjjwWSLp73G2LgbQXB/uFRTcJ
F5jiPcZUdCHuZyhBFSaEbWKe1GD7ExQ+CM7fg9rK6me337BerngBJiDGHuw31Z5Rc5JrfDCoLv1/
66qkfJDvj73G+r1/bKu+aPuO7AENI6wbMz9hHitdUzGoRtB7T+jRaygpYCHTYdk7x1d/NPDi8rLO
lzWqwyqbP7rvwjeKr+0TEp1+p9TfsCsr1ZJuBKDzsKbtX/lRtHTpevzzAjavppLenISO5WIbWN7Y
9X+jMqyYJTke1FQvJO9o2VRJ6Rq5i7uu6KN8FxTdW5z8pchA1F4U9y1NxY7IGiTvlfGSU3tZ7et4
ovATJNky9fmp5Twv6A//S0cjfOuK4/K2mxZ/MLuP2Qb5PLy3IP+zDESUx8FTr6WiXmpeM/GivPAX
3dZ7XiongFMy5JM7uuFrx5JXJoWiq8ydZRlQ6i/deLN5pUsd37Cksk4EIe+Bu0M0Zk/P4FkY32yI
PwCPOp/99i9HikZgQhUmuRbQd4tUUNK7kt54QNQco0AJiXkckoWeh9l88x6uzooE4y7ty9qI7vpe
6Yd8ss8F23C0JrVELJfpji37Ajb5J8q+AH1daATrPrXqD6OXw+Ep8lMp/vA2AaJWaHaWablIxSR1
aUHPgI0EQiwkV19DBwkuxFn6l3siDg35UxOUT909lIAc3cjZJA7DuoYfUHUzCQKlF2We4iEDa3EY
XCRfeLZVlwOj5MwoLAeb7T6vXvirzeBRE1dEqdGpn2Esh9zKqGpTO2x1SnS9a54crCd4qjnCbHEu
TQA/Sq2OqIF+Kt67KxuITD7TjceILPWv7RSrvZTgrufGEmKiS5TZqLn8QjIFr8C0vppH3p1Wk8TJ
uPbNtsAiBFsnGP7WYoDScWJazGUESS/+SekV6pdwJwPeC0YUb+t2bPYCY4ZJfoDqIgYjRBxE4lhH
O0Ig5L0YZiMLZzB6bu4nZBPB+urD5cvjUeKWEHZf+H0pxsyVDv1/C2j8nQrtp3K6g9EaM422eJ3l
ga4K5n7S5H0E640b9md6xca6HteKPRVY+zef21aMT4iveBeXYiPHANv6xwPMHM4uLWX6Z8TBzqAl
sA+UmLFPSV+A2mGbKOPqxOsuQwNiKgGohizZP10WQwtW7niABGbpXNLNqR4r+J9R4UnHxjfkquPa
KrRBv+kseOuoTUIa2a6/ANpz3+Q4W3VxGBz+DgbuUu6n18jiME5CpErFN7X3gtlbaK5M9aP/2NGi
x70i/CI+KzGtIKicvKy2+yamQ8RXAtRMjxWXUG/m4i1TubE+14WAbqZnHA/1IwS8YVj0B0lt608H
cwwjNiIyFYMXLQrTrpFqwHc/pstl4zNjmEcfgDV0PSwXVfwHT+dvRTL7+J4/bKX1Mkyx7fJrXQo+
XQrguoa1qmDsPWzGPgYTDcIU3G0lQFmWz684B1J266XGnmFhWXam7vx3hv3aLZ/NQNrZo8Pch0ed
Aw+vE3fG+WM5trobCBunBLUlqWGQJaHX4Ev1NsDqa1G+Eey7E8gY3zVB6bJDEZ3wHqOR3mSc+Z+k
n7sUuPYddNHqGw108sohhBxyrvr0kCgockNqSCa6V2pSY8r2rBlYb7ckN1DG6SFRuX99GqnUWptr
cOEP3G+4d7jpA8pVmeyWkd5zExhwDK7xrpKcvflZsiJ7X2eyt+fpVTguJSu1/jn9HOMyFAP01qll
klYu1nVXxWm4j/nIa5ntKQo9Ufve0jA9CHfZC5B0QgRh6j9Cxfn4vzDhGFqXkg0zFnxQZP1HuoZq
JTzmdF2Z4lEkOuebH8Nt3q7jiS1WoSPq1M1DwpTNBLuZSkPBr5qyaUN2WINuXKyN0iQdDB/7jorW
lQPCVk25tzmwsTbjySB1SIWprl/b/a6UclgGNBvBjYCCcE8k6gA6cPGTh7RyWwK95eWjfV7CKnFW
M7g9Rru15XfWHotM/5D3OE4lVrVYi946FhI/DdFrcOs0DFLQgVM8Jp+4/r7PPeX+FhUUnmMhGnwo
aGdDF/7iVh2Xn4RXvdcnXWayGGH/pwh0GmvQsuTz87EFRbUA6IxKdcRobLU7pD8p8GorY6/bROlf
EH1Kt5HVSoDXr+JqT+bxiBxOvAEanoU2vy8GPHGpssFod7ETRCs6hdjvD5Zlh+6pm/yc1ptc25bT
aS8UvHZ+1/II3Gw1zlVDKs/Q28KEQ+RcElrhFDrt4GQDluIw+t5Bm9ce/Bn5MCfFftDJxoqItyoW
IjyHdNpkCGMCGPppXG2YUZ60wehbKVg5WE5DQp2EJ2DQUCN8uz4JWD5n+aOzhlcq0iKnvt7tFBiF
BLoA+3jd24nXUSuXEvQ5XSZo8MouEF95hkvcGQMBmz1JPoQpG+hequQxZMHixNh9oIsSgMhN7kKG
99/+RnbWZSztGXXia452JfApCRajSRfgTCchpqA/LUDexVncFW+J01SPkIL498KlJzVV5B/dYadH
ETF5EIzCMt+0VxoTDHHDjNVYXnv+zL/6P6iBrD5y+uzDFBi0l7sEwt6caqO+xtlY6WIe8qgR9ynF
V7mkeTtFeRC/AunsIJT+BZkhWGdg8kKIV20rMiQzNz+zw4DT3CjR4FV/MxAE+yhfsA2a9NOfuCRS
eY6tgRUiW1tKE4hPA18zbjbS1nufRD8O/4Vmo3CY0WOB4ebfCEOQX9T5k95p7aLiaje5h/4+MO1W
EPxmp2eVbgVwQQMIflZPmRC66Pk0YcPDSfQGYIntmmSb3/fNi33UctbUtQrvTD5TYpX1lpQ78THe
edda/Ffp7qibn3t0pD4uDtYfWKMAGeFuKyb+Z7+34Y62CLvKDCQPtu5+X3kd6mdkLj6L4bjYsXzy
dh2kUkKPRg597T9SKFSSkOULLCt3P2vFMMG++d80PgvwzlHmCHobZElJX+QiQowp7b4am3ATVL93
c4ND3kB0oMuhgLfS5XyljJi9SaHkFEwUVySG67VUgtYZInw9KydJYhXY/DFH6fU3hOr5qOISt+ub
iUQD4DrHNhsrBxKBGR8FuUsNRreE4avJ2FgiwrwDWawHJCRvSLwyRrufcn+IfStOV/QQpVOPamK3
iXBRCrPh4a39nNzNWO5SYOgeFvA4sQoCAQ7GtxW4ivLf3EsA24m9KgUNvylpgIXYzLCz3mw+D87h
U85NrLLTDKeyPGzmyn1M44OMbnOb6uvhe8CxVS9b+CfpSLbxDFv8Mxdbldllj/8g3pfFdMSEYZTM
GakTFfVy7u4xSXf6HUtD/wKHXEss9PwpCU0tpViRT1J0AN69dre73AErCyw8vaNxySD7jzKU4B0m
H9di6tiqfJqusU6aOXBjATsvpsp6opFZKMfXjF9cQYUQ6S/KPZ8BJgHvR4humkN4E7zEd/JzZsKN
yFLrLQupf4Vf6BGj8u6yBuJus6thU1ED+MO3k2BuuAgSipe64QPKH55NaHO5n3BS87oBaY6tLHP5
RRQWKkEONYcBNnDoWJnvQkXCqj2U6LmpM/lh298UryNQvjBykOl9WUX79aC017gnQGMIQXRYf8e+
F5IKQATqpDsNMVZ0Hm18QhojoIJPO7LagjkDDaek28IfVDKlIrHcM+Q6EblDNkm8wC+Sm7ycn19r
6ETNYEhMcdVpwKor+LB4Ba2AWmhLizlI9LLnizlnLdSEWUcuhUj+P/6VGcZtnxzf/hcVjuYdAGex
JxDOcgm2XmPYEK8J+pCRSJfvdk3NsqxFJQJhuTdwx3qes7cszCu/MhxEo7iI2r3d+qoUd3ZCCTeL
XsiJhPb80jVDhO6MzdoG7WIPFCSof00lDFi9FePawoCFdk1cx6chNDQXfiSwV+eWfby6CClfwWlW
lK/N3J+WVLO2jtd7g+RG/ppT3Cdxzs9pBslfDjO+Qvlwtv2RbdiHFxdOFoP7OctoiaE1tSJbaE11
M7Xb2hIkHOAMxZqsOnKJsGTrAIi3jlYz0+W3PGZJG3ehOGawfrQgsUScuq5DqiVBMdiqa+rPpvlW
+tjVXj8vwpOTseSv/Y0x7ueN2uUnowyytoaHQHKOFRmHObwntOXZjQA5IUjwDAYEPCDLAUW8Dm8W
tYUQR6usxEKsP7z48ZQ+1/516Zrp19pUiWPVqwxIhY7bNPBokxl8kAdRCYfUyRlgxaZ+eblNzZys
EQiUuUkqXpYV3fgHcDXmUTZNxtr8Za5ZPz8jhsrJxt0rBz2F5/RZswDZUUWCSyLKu7y89NDagw77
4h1x4aE3BNB4q38UJ6m89JtqrRcGGmpT6Le2n0Eo0+iMIzUEtiaq9nGkOIutjCzQOiSme2d9XgwI
UWt8SwREQUwoj8AJ240rivdI3bVHkMFBNmTuSuIMGVyjVuWfEPOxnEbwrObadJLsJEsEibYEo/EW
J6Z/Rjrs4wrlenCqNbN8vEeYtBlKye3GbH2C3T+/8N3iKgv+u5NKZu1kyTtGZB/Tp3u8ub6xezAf
mKvegTN1e/sVTmgdhy2YUzN+uniw+/SYIxsjkDvTxDTM1EgENitZm0Wxj51mg5ZrqBY+qS5QHE8u
aOcXMilz2OtL/zz12nkrC57YzszKcoTmd3z2zjp39DsSn2pZQ3LsY3LK8SEdAjqikb9JGvxDnjl6
h+O/FDPv9GHWZp32A9Md5pLqehFwv6k0Tbtx36rt+hr7r1UUM2gksF2RpAzPBehv9rnxAPAHO+Ux
Xgc9NykdK/dSmuNpS+bIs6RDFM492VeC+o14s0J3DX0UdwuxQUEB+Cr/qcOBJtYvhjPP97+xIUPi
IlpBjY/xtF48UmLR8YLqTh8Nz0vgUJVGCWOPjY4rbxw/mnkg/RTtpUg1P3u2YVDWAIxO9e2B1OFa
Q01quPgwrd8HNXes9QnEmcQWVZvIS7rXYd0UsBQ85Y/T5Uoa1wa8P1Z8jQIZX6y873YL2UIp5zYl
ltvsRVM6kiZd5Wildgc7S3Vfv9aPKtwIMpoGe/fJFMBbmEpQMR5Y6om4oaWMsvoyfkeoRFmQOv5e
5o72mqEpn5HW2aDhiuUrVBsu5SSxGWn6Ku5U3k03/PeeQAPrPIRPxTFvzW5sFM21kbQwOVfsgIZX
AW7XpuDkVMysgqjkf5MrANSlAzDzh/suSd+MrqP6ullUquagdkhFwRLbBthPCLFY0m3QOj1CzzlR
ggthbNJY8g4dSZdoO7vpEcqP3t/WGHFVKsdfylrjMZHSI1icIzxnkORNLTRwDUzO91lhRwPGh4IB
G6OVBIZUDdT/Xm6sm5rpA8chU760ZH6/ODl2pLLDohcE6oHc+RbfqBOpB3nPWdhJj3BoMoF+s2lx
T8gkQGEUbvd8fH6ZV2kPIAuDqLHzkhc/nmHA648Lxjv1xlzw3bO3yRhGWXsvwqMGCy/7miIRQGns
9YPZf/91GcLBnaEFLoR2Sxc3xqHfODoW7rQ00f2s3lM+dw7UeJ9cetKSecscvKyErYKGqZP9/Gpq
w0ZTr0XAi8SLUGOl9popi9byNZEbikJ1AcAJYZ4oXBNLd1ghV169YnZpez7MxV215+a+B05/61b3
OmnAx6H4cEjkR6ubVldutHGCDP9cDzqayRsSz+fND195nHA8O8mywVd3TreG15FELEIW5ey2/dvY
kTOV4cMBdL6yRO7dbxSYwNeY0ZJxjoHnygKMv9JWjIbvYcIPeZjo3Wknatq14BLY1f9mLY6qDS/A
IW6dj0CAi6vU4dH2zYUXvRBOA53SgFa2tLAIh1cbUUbhRFIwI4c9x+Djv7M4e7OE4kJ82RvrXUFZ
9D3WhOfSW7cjBQvRMiqUqLa6U0l8VTJvGt1O/kcUZXnrPPzPgNYaFNI5fjccLkNjXN7Cr6bg9MTj
9MfqtTG7zrGt7fSV8c2R/EkyT1nxJu0vaKm9RQQ/GMENP3t9iIurg5aUY/JBKaGU7ORAUQZZOipF
VZ1FqmR/JLqn897FEbXHOfp3qPW0S9vXKB+ffC7gPm2C8joP9rqUCQ0AoDy3fxK4T/Re0JiZdd9G
CXLEgr0NRR42UuH3j/G3PFCjTyv3l4DjEd7v+QOvC4s8tPU2QdjgRxKH+oiNBtb3UwBlA3kbY9uG
q1qXojox9z8p3iZ3WBF4GySd91w1xdDaBl6xYK1+ULEpgxWFZniDPaH8CZr0N/PINv6fvcmGjlzC
2nHbyquNWyNoV21JKD/dm2eJqsnhU/3v011K0kiAE3NZSKwahxymxLXJzZgyqOLFkEETTVtI1l9u
vA9SrIBqvCL8blj36w6jWyjQRWxJ0WCYAb/2f/5AneaTjox7POV0P2qTxECGOqfy5g8EZ6qt3jH0
BBnckxknGmgDj5oiMJZo1LbuQ3Zf0kh6E9QCd0hfdh1KWv8s3xROqrMsJQQJ4Ohv/d7wNid4uJ+g
em9ljgRCdKPEMdh/4dSi/TjU19nDaOUMFrN1TS7XYGjA0swWdawFQGKYyF3WIv7pzw0kgAKE9bfA
RJOoARg2AnpTH647FSKJdv8cOeQCbC3euWSYt4pZa9YFHdcj+HkY3DZKAVpiAijladUBC17E1BaQ
3cqw++/toFb8FPb3WJBB/EGd3eAWLnSIZQRJYh8wY/wKcg3AJAEtcfh3ZSNSEgZdMnK60RPkxa8T
ZhSTZLRK3nc4y7myTommVXAifmlTjS9GLu5ehmjvv1vQqvOqdx8cwlLGfHLyvq/aO7ihCUrHcYHa
5IXHZrsuYKcSrMzIt6OzoA9fWV23iIansihcw+03TQF+o4L1yz67ApN+30iIhOv9SjYEGB48qrcz
R65/hECtReN0y0nhxpeHZJkz3HrcAaymmBUZFWrjHOv2ms2d1GJae2WSBZ/xKepYJu0LgF32pMd/
NAPXJYSLjcRlOq1uL2saz/eEpQS3LGoplWub5nzINrbmdugVd5S2YIxvRxugPKQy3Jyf7My+gm0r
tJZOl0YaB11zVgnNcMEp9q+SB0gNEV6dsL/y0+tlC710N6OnBLP+8WcIJ5Kc64RqoUAxKyj8R5WQ
+QMDuL8hh+W7HLx/fGIoAjoep17Rqi0hquA7dB4Uf2RDm5SfRhxFTDUQGzQjXmJeOw6hdDkHjVDo
PBGYhtNg9Sw+U4Okd7q3KjFGoqfI9eaPpPcl2BAdOwYKSXPyjjr/ijmxagBeGVMBQEIYaGCwdQMK
qmcJnMa9wDPizfJVrFFO8RnafKTQFq9zD26fd0tlBKBaDiMgEKWWbwufOWt2kYOAjOwG/22NA3Jl
fVhHI9aAtNuy+0gCmFvEbjddXmM0soz+YE9UN2uyURzbkvYV0qt/CrJriWrKlDwejF+AjlTFJptQ
EGd5k0NTH5avWr+7zEKOoeBC8k0DFrcCVM8RCdmSjt0u+HCwtL4+0l2WeyGsCWbsxcQHL5ivCTTi
Pz3VeUSc4m3s6/rsCS6/58CDG20F6HpEJokJDrkudP3/Xu9h1+dr7P3uZU8M9KWxw2pcpywKMZJK
ljd4F5L+boLW4DRzrFVpDEBk/8EffxZeXFsVeTxldEMcGLU/BlAhpIG2kFx4t7uLEoEdhFB/tk3X
S2hFtllACzeyyc6T1RfDEkOj0RMmNbNj+LPU5zjSBJwHEec1A1YuXGzmiqEIXeHMTWgU+qb18V9H
0yPOb6yrZgiaf/90/ccHuPsLhkh8uns+ualNOq+5K3tM8pLJ8cmALaW+vBI/IDGKqU9cK0xfNzxZ
jIYP604HxWShrv69kL1PvpghbW2c2OvlnWPegfumijX665ve6g1iw8goXIWuzEAp8+Ker/ZRaOLn
ETUb1SnG0WoW1R0mDZQwl3nFqTzhyYEHQjdU2dJADWpA+g+5QyZWktRKkn1ZJ5HkiljOXMRkhno0
0qHgOyxeU6XeTY0jGwCobHWPUHUCwLcouB4zvyeRKtGqqOHHUe5ZqYOHQzRXotrxJrcUkHf1Qnxk
PTX6eGcZM9q5AnXT3Akmi58VMG1fAbGUZTVfYsz3t9WON6zso/g+VZx9spVLto1ytw2y3m7F57FQ
m4CHzGm+TD/Effas0uii32vCdL5k7e0IwAcfprIxMLfAICVCf27b7vT3oDcpOo6dWhCm08ydYI8f
V6V4UJ9pzmPLEpJKW1eGM8cFHwJ/LjpfxTagjfMSevTsBNzoR8dQaVcZNAs3JcanXPvCibztewGk
ldi7MA7pXjCayp/ax7V0SZth+zQLGs+rjkbVgKpfPyYArq2/A1hy9dn2Fv2uD3iNznH/5onFlmrk
nji1eFSAUfLZ49fvAeoPy8+eznffFNaAex9YXEOqvOB1yr45zeUibtieNKqiG4nJC5qL35RBQ5Ob
ia4+8WQPZullUd4j7qu4NZzqrIBDboDBlxYS4i1MNKlGb/aIG8bG+Ftz9VVBSgf1KwwxqAMwGByq
OBzAgygO6ceLFOWTmAKw5ag6h9Z8FmMrt7ftwmkA8h3SAM0SWjZXsDoQtAUnm46hJ8V/U9Wz8fo5
4iMeGMrFQ18QPz+BlI1t3E0gfxAEcgA3js+uqH04iG5szEPsleerCYic9i6TEn5kiSXGTRNHOAG6
0uIa+YI+CltB1vQuqbro7SQPRdtU0n1UDBbImBzjMduhlYVOS/Akh5t0wYfcVCVhseUG3QE0eI+6
Lu2VOc/IW5hD0y1LD+KYTX8UgkvYuDUHhW6rhO073f7Gd3Jg4iS3p7MskTvJHteg7aPWhZTmkfFS
b7/6o75AFfmFuHXZup2fUZhFqdXSanUCRWFkltx5+fjwNK8xTkaFQwrTWMSMNu2DS+ncFdbIm6Wo
IoeQ5/xEnlODbBBx73WkXduXaDjpskItShQWeJ/Vhe2BOnOkZ0TKNKXYnJcyLoztvdc5KJdvy1RY
OVhlLgaEH5GunB8QV1pNXSc9q+uw4Qab66nlEvR/64ZpN3jh2W1WLToTslz6u7Nr3Du7NG9IBryq
ugXn99WDuW+iJN4XG6LDJswkA+iUsAz0CCgbsmJMz72glk36t2XwVWneRYJOw9oF4J3U9Nyou7nU
av2BAss5e6hPZYEjFxfIGya9Yxj1oIruK0vmilpdo1J3wrZYKvHOwsklSS0iztMg5QV9wAseQinU
9tu1XCaMp6Nkvjq734524biw/5H1wsI8/0wyFjD7aU48u2UigVI6lG5Wt/JRk6ZWqwe2PdVW2GwD
730uTijJhiIRA0OD8/bNix3B4JYb+JyzU44ExgKJwc8O/zbq6PSZtQOTVcYp0Pu62ZYhTsW3pRQl
QxLmyJqsVErXnjE9kwBzep29OVzsPB1mEKMRbbO1UyGGRYr3kHJjs1WuhQjxPuAv2hCor3CUKvPK
hJB4fPwizMPCW1i+ixfcg5YzQIQaUS/wsEFIko9RHk0CwA0PYZZ+AfgKI/SFeE2cKUkiryEwAH0g
9AVr7zffM1M1jwrNg8XyrlRGJQ7dLn+9545HT63TBxTrCVwf7VA/QTeF6RpbDys15+a1mx7VsO4w
iE4sED2oc3fkaUdVdKD3Vzhy7v7stp9Nen92TC51PIP2+boJskRAgDsWCDAXp3fZsKYJR94mwvwa
1oxmPCunr1jQLSfg7uvPYa5Rn6DmvxD863rbBu00Zj4Z4my0ln07bulIVVGruGp/gO4IJ5qiE/IK
Pl6N4n/446ls9gOPN/RHj1C2BPQ9aqsOeBkq/E7XI1qhdaqvqYGXJ7F3yrjalm98d5k0Ny/I9bnG
WdQyfva8XXGmkxgC3sUv4/obHo4e5gStoixkSey08vbJwRer9Rgu9UlNlqqZApoWj6tk7NtMbnEQ
1C9903TWTKMQsp3NuWtkbmZ6JVb8DELznD4iZN2gZDgtYd1U8BEH5AAiG0nyPpoHVRl2Xrsk6Rsp
2s58oORRUGCplKK9HPjD9z23/38UlqqagWVH3HrPdTrF4UNO90T9C5BVXcLZjrmgW/PkWv9OTODA
siqpm8Sfq6N0RbjNyQi6SImgNmPKNW70d9HPE1w1heB9YwLTDWJQtPjBGk5GJbQlJB2FbuzaFW9E
8T1GbI63K8adDZna7yeuFEAM6cY2P7JDnTyR+JlgUNgZVBZRpG8K0ljUG366/5yJ6ZGSAB8i+0aK
7dL+62Rjailq/GOrvL1DRFWAJ8/ykEIGOpRRVjJkxZp0Wxd3SJOLjwiFBHMd5mR28GKVWyqH+XOZ
Tw0VT0yyh1Kx2IX5nadywP0NzwHjlNkVI7Q31aTwQgVXuQwYIB9cVlGyxXFtKNdHB+xsqqOlBVPF
5phpG0OCE+nHqaQIbrTIlNEov4OQdz8EubR0JpAMQJeYj4MeDwRdurzlcrrlGhXfzOYKY/ausd1l
4QAh27q04IeCknj/LAx3/QlWLawLIuJHhGil+VMA4QIejF3LZ9XnW+AbdCWpYjgWsSFg0sG3OJ/n
mwG4GKMDJkuVz05Zcc+QK5PomzjGk2d0b/4xveUp107Z+EUcJnzYECoRTh+XFPUcZptcY8EkqfFo
FKq/4Za0Z1VuJHXM3ovYCuqps4XWs5oeGq8Wz9lUHQw/vmPPYGVH+joNOlTgg02za2l7UHUta8nn
hR3cN1UbVNtMr07bJKp9k8j994wbzXUPfgCp8c6akdtLLKnKeDPvkpxIo00tp8Hurw5TxpfX0TZh
0fUJ1h2NDSwffk/AiwrztCiqY8g2uRjnzYaHfj8MIff1Sjx0zY7cvyNNpVKMnl+nZVQUGQTCtrhx
rBdGFjmlal0aw0ugn56u1gDA0T3HYX7GnU3eLQKtomRkTCUkXNDyTW/Sd2DZf4o7dWMZAJrFqZUc
ZO4n1Wn1cjJIVnkGWUQqwH7CI646p8HGpQGQpXRF15GL2iAwRcYQtW1s+M6kx24tlnVTZ+wHjyd9
hyaFaug6JLE5JMKhyIvDrl607Ym312MVH1OUVtu9Jgj7mGMYLwEYkk5v5yHIdp1ee1yvKHILWZU9
bvTKCmMU44aMOo9oLmec5AZSzhzxrfj7+17qda8AR/8tkGqZMcqnfrS6MJdrw2nLG+x5fqjTC19W
zoVCzs8VP59GXUdiaYO880oPE9h9JhGGZw0FZGOBURtzZE1lv7rWIod6On2GCPwepTAe59PkElQk
/BB1uGm1Ay+DixhVRmDTnQBExbJRmt//pz1XyikQxrWB+1ohMTkBKAmSmqXz3EwLYrgBfbSfQ4CU
kcgvXX7e+/fl5NrrCAK+YRvG2i+txrfBuTm4JgK1Fgoi4nU3qRTWEobjTTI2gjjrSYnnxfCSJRrr
Luv+hQCjYd3PP5N4cSoBoQUw3imPjw+J6Ag1L6MZ0SHUq8cljSHqVWXq9R3tYCu9polXFkLWh34h
VIDtIElceQymua0X26PJ2HK2dD+g/u6RRivcMgku929iOmq5RalN3epMqcPl8jwNEAlU6yirWfWB
hhw5Fzw3TerF7aQ0CjSHgJnytuSXuZuMBrrj22VhO/5ywMGEQ1KqN6j/Bm6livRXOAMjC2mW1YWb
4tWeOmV+EbV7vgl5w5uDtwZ3akL5aNj7LDnZgFrwNHSW4KxMbJYaYw4SRq+5gWqcIqSCAmHJtJNm
VJ9wemdrdwR2sRvnGbb6nVhSvLe0KY64ns4rVJM7CZ26F7PVyGrliaXjMxreexmFXGKS/OAT6t7s
r8bK49+wdnHRwptXxGeEobhHo2Q8HglPki6NQAkuNJ/pRcdLj7oxTEd3rh+rX/U+hDCeNYhfi1kr
1FWKI3gMBaCmHG8pbK/kMVCEN+J/S9FHC9vfGKR2BnAkvQqpBJn494Eeqi7n23lGNsUwFIwCB/B/
r2MVxRnVcojJeXOc0yoVSDXODrgd5b0SN0dLRjzojiZL6/8znm/jhabeG+NqsJOLR46M8RMA9+Rg
Qt5BrmV0M8D1rDYnhKPC0hBxb+Xys2ivGSYq4/YoViZZO5b4h2u1XFgJiYcJYh4Mp2q1QFmFFqQp
fl4bxpSy/XzjQv/OG54ok/moIHUehasqwrGsZpR1qhuExX9zP9XbTgVci//idV2yaQ8ZViT+F8nT
yZW/bCqTw8NIJPiA30o7qBn4RM/oCpmsbyBLIORCEseFb0U7YhV6+NKlYcv8L6ru4BF/mzakOPqg
SiAyQ4nZFO2RT0jqBp8Gmyes163QPQ0oTuqa8813rUh83ODTS8Dini01HpjmD8pKJJd+G2u4k4Dg
o42MRuYrMoFYFLb6MbH0h4l3IAIsN/jg+R604JthfM/NACs+2h01qyOeIozoqSB8M2bQH80xk1Gz
Yg8UAExsWVai8YuR4Fnkh6MI+Xzi9zdoSs9PWrcfYFw/YzqfG8Pwh2ujk93hHtJfMPTJiItyMtBx
3g1Vin2i/bsWvSppQrWvFE5FqoZEhH4vxoisaq18fYM/YYTl6xhFJOE6+BR1dfkD/u5+S25eT49n
sUS1HNwCUPDcVB9FAfyuuykjjZ6w7TSfUP31sMr5qaJH33ZTmijXTM9qco3YMywid7TfbSvEI4Q2
oFy1mWxbMCAjZB8rOpc7PU3KhxlBq4LQxnmFOqsA0CWJ9e62zhho7Bo2rlxa1+k6jzr9oIZf3CRC
sCLkM8GNyHtOrjuq2EISl796bb/jsdbJPXNWUVucbxeMb/Gk90l+GItsUf9kzVJNoYL87PH8K/gg
vvdZ/260lVNh3dHI2y9/clTRVgg4HQKm4HNr1oHmNDjX+mHk+LFt8Xg4/uDTmcE8HKSD2rH2vbT1
yOOR+LIWzqlKxPty9/95CKXNZQ5T15QLv+wkjqV/A8kBdjrGRKNo+I9jcUL+31b5lQMwuT/XsJ8M
Aq0EJrhl5ka2Q7BrhKcTxxMKlhOxDbL3GQY9TbVqT+z6o6zQaO3Zv0uUm3JiklHtwjcItbAH7JZU
B1MX3KiZYWLHPsrCzdwFWPT0hY6Jw3ETc1scoJjyUN9yF20jZXbBCMamNUZRY3rbQvwh8KuGIgQ2
CE01/XQX7d6xFrGEcM2pR1mqjayeTdPhZu/CnoTHQ5riJGo+q+ZUcuB4VRRXHjRJf11tK9VJLdkN
3B4eDwj8qlQGMoOdqhzC8ntEhRn1CW4AcaVv2rFr8YphIS1t6oqVmyBA/dy5k5ithvjk5rHHRD51
jkswSAYjRxfZy9aD0ZnH7J9Gz0DG1HAD1Ptwi/szPPuKoZJLuZXCOHKoaTd89aa9ApLtlbiIGGCA
qZSMLABYgqYte/AEQCDBUsiBT2jcktNi95M/9s4AL9WXjDOjTOhbj8S8t9fk9x8PkKOXBaDT9ZlV
bNxdXZ3VQh8lTmvdIeHa7UnuV6nzM6szEgSK5PG/1BFA/On0PZMTSBaY1xy4U1sRmqg8WZ6N7Mud
5AxFJHSIlCWKOlzchEJfxx17WRZl598+GFPqMmV7nJ9mmabM7t3JvFqRJGhdwxDsyzhdyDE+mi31
b7PCI/wirjrCWAyC6dXp5Gw5WgDRoLjUqH4Rc4GvvRWgmiTCjATpjg8E0Yu1uU3ucderaQ32GkMZ
oGKLdj6zfr020E4Cpgz5G1AOeKaWuTu1VCGPjkq7TH9DAlu+ZHOgJNOQ2GIBho3vlqxNuTTlbpj7
nHY+MeLUGI+jPd55LNO08DKQIIKm2oIAuJqb4wFGPHHLJ51QNXJs1B9ygPvGBy0qo3z34gmbdo2X
oQ7hhDActp48DMVZnjGnbPrzIYKRtOjboJqq+SVcllEyroBr0D34PVJCyEj6VletaNb21zCHe7/I
mLrUZTAepQn4TD72t6gwzkbfjkYyolzph7g0Agf4BiRmyy3VQPUiT3sHpX3ByUXG/wGufyvqRVi1
QAmsO7bRBDN4MQ046I2zhQLeqbSDhCnODRh1LXWr/YFeqYbqFzEgY3q6XRJkmZumpAIVS/m0n+Om
NKe9OvEzlxLkratzeYhmpCMqBTA/zsaDw0sg/ZA/tzccUMieAE9A7aXZiT2CKUlabBjd2N3qC0+T
ARdU0EddCizfXiMrv9I7hEcZ6RLa5iKw1qHsOrwzHbkhF96G+jcHJNqjUg/XbEigYxnFNbh+Fwzq
Wu/A2B3rmkMxBOwkpyg4e44lHQCT9812cQQo3udlJPrSn5yAgoJZakUDTkkCxG1MRHj5pZE1V1q5
K4sNwD+XbNbYMAV4qzj5gr5n5FwAXX3LPigSZ+bz+w9NsUHlxk0PSDC9o9fCS3oOQf2D03LTfrn6
eOOr7rkUpclrG/rxyB5j3LH5nhwluHfMyoYHn6aunv03HbRJ+s0hAzH0P+pMlkIj9KBUP0OnMwtf
9vNH63ZGEvr5hYSy/ImGpYFy+JAsc5w6bLjupbJ9HaGeWYw77EvzrEqoH7UJCEzDKYSVdokzFMGi
92uM4MJ6igtzXbUgtPZj5IvkpvER2tzlC9nBQMQHU2RFPkA0grr7upK/KbI50JZNmmU68yKaQTy3
WBCCV0hKGLk9FXpiYZH2JwNzCgsORe5slFDUde9kIWM84EHgj6f9laCFrA2hO8rIqvVm0aOoZc12
g/2y678gCP4ZUT4TGA0gQXuOWdIX4CD5eq9y/l2pUancHjTpm2SdAPaZt0u2WItli3ON94PmRR3H
c9KWuO4ByxUKibw8RgGCWf2ZAGI+ZbkKyBqo7tX+hCYKfl9zQSOMZhoTWywmrN7VgGLwUse+UjuR
IAsQjwPzKJJWpK9UDv66/Om46RJc4BtVzULyixi2WOZc5CpRQMj1am6WnUozmKIeTxIMH6j6kRaH
yVllxf8Yhahz5OyqXx18psZ4J9BnVFCjEdXRrCsEJrE72EIRTY5LIcxBC9KktK8Yyso9CnNd4nve
n6j5NGwl7OHhHpLeRaBlcEmeBBf6kcOSF55c6DcmaAYsP7197p9tD4IAlKypZfttCpCJuG24M/Ya
gEOFWx4ZxgWHhJ0UbouxE8v4v1MvBwoY/qikmMDEINHizXEtgzg8vXH7ekv14OILDOq6dqO3c38P
juGYYW8+thqqHOgru/4hzISNm6RvlgM8OSadDCCGIsAvw95mQGfTKh/Cu+iZI0LIR/+JyUvXfYYJ
ddal+E0gFXBrQRiI0+frh/p7tMXLMFbM4j5dO2UYN9rlafiANG/t+subZJTz1MQU2R3WPeoCdMmj
4UjbtEWnn09XZOj39kxiV170DaMNQn2I2m2G2G0F9cHL0Z7Q5b/kAKaLxQ4nnzY6opY2CRlJT0rR
RHBkLwXkjNSl/wfkGNuDuCtlcA1p3sqam3D29a/KDgqP91l2z5T72kWUvQ6+gOcygMGZpPSVGF0x
7SAKdhc5iyNO5lpKvy6koHpAKRUH7EZibt1jGc7u9A0Gu5f04+4HT+wJFsaasFpyr1iV/fKtNpGJ
409qVALO7tqdvjEwViZgyCg4nIwXRZnh9mZI6sdnZrR2p32Mwr5UMCqCSrrJRp7+bTQ3nSj8m2Xk
5aRBBhShuN5E0uOTJi0KOrMmPi7zNwD1NbS79Iy8L0OW8TnZmsnQrUyowZVv9B/c6HAc1i5PA/sS
yfepW9c/3WcXj+Fcfe9gBlPoCppMVcxb+1fde/jkXkmdHE/Rze5+yCWdR5+jhPwO/Tu/oQvko7zl
0tcZm5VU+FVzXyB9HxwKBKDA6P26B2W+oy8slMGuZRvS0oDUClZwE2FrgtXDOKqPnMGLoyzlpMD5
cqqKI06KlO+jYDeDBCK9yePlzszIyfRhnKbV52d6dwFLZ2LtS9ao7JopVB7zHX/GynnyYn26pIU7
JRr9R2mAQ1yI85z9hDVgVpKwuZAtrzyowOmsuu0GSL3u/yq+rmPqhaincsaHeHl8XAZn0fa1lVWP
ZpHXaUgpWR/hLkQ5UqOExCag+di6EeBg9yzRMvcbzWlZcWvAm/GSlMRksP+zahLHRNlA/FtQrs3E
48L4PgMEKaVFToJ0DhclEGpGgcUQmQq5ug+Db0v3Qhnc3cN/YJkRO8F0RegQJBTBfj/lfATXBbmi
t/o9SNrWzoUtR6BXKvTKmHjsCG+Lve7Jk/dyP5UgT/l3MyaBbQA0625ym3kip+xPTkLXbcX/t6Zy
1tii7He5kCaqCg1kiSNKwJF76EDu+7GjMCexKAA1Ygc/A+1ANUQDjQqIWKSNMVzjDKUPRMMdexqf
lNG9hriEOV9zkVhmMsfua0t7OOd44lU9JCLpe2EYP6kA4+3GpZ5LIWzdQSdi74Vu746GEORucI/j
mp4QvH7wBI77q8wz+KGmhjGeH2y3DZ1mcWu1uSAuR8Xgskc0S1XI2EBy7QCaupEZP6gyL0triy6e
p//n4E2eMbx1PdXSsL4YiGCLKLAxZlULvi2aeqGT++T3t3fOGs4ioiTDz7j47nVN6j+8iSueL0fY
9IGKS9Yinir9N5y77Ajx8njLbplAeRvgbsk1wJzqsM2CEhUYIhMe8rCoFyXnPopSpUcFDJwCAYzk
gXZP1FkNNWDftAeyBA31ubrcRDIbq8FgYp5cyykDQurk50sDg83pphvo/bWe24EazCAI/AHkLgF7
SvFPC1YhfS5vu3UgrPMy2p5o8R5LF5SHAloRFuKb02cPj49qSnZCNAqKRsXHvenHnBkR+LK6Ta5H
QewnzgbAEEvZaLqREtb57l0a8/yQHLe3yHPBDX59N0l0Xxw5wBNXNg0DwkQpoUm82FyAF89Bh8jT
dYkwsLK9m+NbMvAMUZ47eujE0EYP/w4mmgbTX+EXguIr8m1ODwrr2/G9Q5sP7RoK7OqxTZjcclAI
HSpHqF4B4iVEzVRNUDO8L4EvrRmsvMmZs0wNFU8yzun6mp5GObe4CIshCcbwZEsPngWnm+4rNcw2
UufUHgSkHEx2f6Qxqdsf0MISAtvF3CcZBJg5shG1zdwrLYz9s+pRQkUkX6NIsMVK3nDG8n325IxM
ZTSAR9b/kRsl1/5LgZDwZZlsVaqJAnzsN1rybrLyAoUomyjwG3la1CSRPhnPVL/TGdF94c2Rz5Y/
hX+YxnlMM8HbuH6clVGxrW4eFBrDOoi3oCXDDG8to2tXfKq9fz7e4A4Axa4O66zg1pxc/gh01CIb
kyInVV0PgzBsUDv3CZ55iqha7gSmBR0YoHyi5l8sU6/fM64osQ5DTzJurnkzjk9yNEWCvAvUuTN8
4oRdN2esxJ50dBkQU9Q1uqquuWV+nPTieD72l1UOh8IUgSfCy6Vd8N1RLOyWIue3JJZgm0Zpq579
6pw8Af5tQYst9KhQsApxLyxHuxvW0sRtv3EBlaHwU12glROXD5/PAF3RexHUH9aB8w4O03izw79H
8+ZriSQkfJsduJhfnKFIX4I91ncS1jtt8VNrcO2bsDvhsbdWnk+zZpHNksEJ5dlKmDBdNiq+TM/f
5zvxgk18lDiLtxM9PMRKOxMtBaVFX/0snOhPFBE/ERk8oUtV3um2Or1uCKpSARfQ81HlVeXdw6si
zLAt1d7X9sGhI/wdkHXlah/Wy15JeFzxrLgAkk7TJBBdp8Gps32SzwoFuz780V+G1YuDvUTropPt
Ne1PcIeMwd8qxgHbYmggUTq3KdhaH1pORds5ZFOcWjB2EBWo0KvoW9TDFZ787/mItAV/S4Mpi1VY
GaZ873F8WXRtVaBirEn5IYrIX2uhA0qbYDoOj37wbTm9zc+QYl6cnQT9lrW2UrNaPANsthZXJgoX
enR/WWWZrhET6VmXm/R2ggO6qBGv0yOOJS+0EYgAUwJpTsnYVaMerhEfy7mHFLUe4boWfSQgVHJV
20gus+GHIh/qUHMRO3oM5HztS8xRkW2oPiSxbf9VOpzpaDkhZj0w5oYSMQVNOlmxgGPQuxly+yx5
Qz0c4NQrr6P1Zh2UrjFohPiuGc55vJ+TDtJkPrXvKlVEKjx2hdtPsMnlvVygdsCvKpym7pwED1Ne
2OlJfIRLExUpgqpUVWXUiCM4ZXCQlnaGlkgtTdvxmXLHGfTFmeBxt5nnGN+Ayj6ony51BCJmTGWk
+fYBJqLIoFUk0jTJHxTYS6A+42NtulOgGthAXzJxtid4u3sDmMzEgOOUBe/U8PgRkkaFgfoESLLy
UHKmpMiDJJy7/J6KD6ZzSLIpSalxuvL/kRquJurC8/nqJKtP/aj2nEAw/voNDwDMdVGMmxZiW04b
zITcxMvnSWkDHEhFy+WJqFDFKPFQh8m0aNOPFvbmj/kybZrk4ukOTHYRoBMFUnVg2kHIXoKDnb9t
aOEUMZknXzRoeCxdXVvQm9MmlcZtFXnQD7cK00bOnooIzH4znhB55PAdF4wbs5MPXb1fL1EIRSG9
McM6674BYgKR42VSNVkenX2HfvsxnE4px/3d433QIe7Ft1P3Vjxhr4P10LNEI9VL4F9pQxNBGdqz
kvee5NainkYt1LoOlP9OKCSNvt395JrKfuDVWzBD08HdtJEPgsWq+vb3cFBjd/Fj/09zKifNXdKN
SXBhrWh+JRK67NXq+GCMZEdvyfT2AhJHP1tndS54vwu94h7Vs7zkrbcVLVIVSefj7LE9DODj80kV
eDPs+f/ThEhpGxJiEdtBd+f+3IaX1yUdi3gAhiWY20n9jgbCc3gYje8hlaqJzELSYj9RRpV/K6eQ
ufQIh7hPJLOZo7ni4hamJwLf4gUEAZMLzCABFWVsWjp/bc1JvsMhDHXX08mO2U+3NrwUmwpFetM0
t0y5Vi0+pk9mx7DhkZxg/NPivBkfFD+J/RNPz1skDpWk6CAB0qVLnT1ubb3EfQ9oRqHcaOFVCFQI
EFgiul65rdgBTl1Vqij0a1QCrQnqGZODVZFAWCal4TggVAzaI5Mp+9D8/WQ3VzFm/tytJxrm2yCh
pUHg0ENWp8ozHPTlF5N4LW1/XaubLiFjJBKwg8Hj8g0cStDQfOqZBjAzC9yeY/9hIGCHIwktzZDi
gNfJcdeyBL9xhI36CZ5QdrsI/qKYEsk0izIhPgzYnyAy8BRwAcvvM80JH8HgFug9iGaKPk9anILn
bZ/IJl1iLY2YmC7G7Zpyj5WiMrAN3tRXu8Z1JTVNBuPZoWCvuFvx7YV0O23FBpJjMKTJE9uPmNeM
LMYAltBuB7RmYEh1FoMfe3bv+/0SIGI1TNgDqeqIjXopUzCjq+gAJDH59zqv1icVNcPTzczXYdPQ
1UmJt+xMJCYAtR4WP3JN6se3KuPbDJmfxKtYH/fluG5yjwzjcdnLeE9KXCUHtjvR5JvK91eVbBt0
Ay6M58B+8kQX0E2pmDwXyVSrzijd+zUNn+14iDugfEHLKI1ckvLo60hQdkuVZ5j+X0ZyT6zOkixc
GDpF3y6udBYKSAC6TL+MDYv8JHuftQS+EBd7NUC4BSi7u+1jHXw5XgC9ysXGMAqbiYuS8z9fiVga
ioLhtXmZfDbyThx+NwqxPKhk1E6alq7gmEJ9TxWEBbW77y8gqDdUIDKF2bkhcplNKWOaWPQheXvB
2V/AOBZYw6trgRUuzyC/T4m70U7IIyfhMZ0NGoYk5EBO89XFE+LQG/eD493wi0fT2g0DNwQGI2OM
kSXqZNKOaqabPEoDZ+7N/rIZkSaQJ0hfOPcbmKO4DYzzfo3Nv+0sLA106QVvuoYGPoeWsZo5zWQO
KCLFuYWPRZxwOygFNL/Fuo9I+5siU11hvYh9u517R8anf8YyDvEqrWK3JCG/u6BlfuTNw5o05K/e
qOuIUKBMCEFgj1161GiSUEQGUeggjvDLubWyT22bOmqeMzCcWlbXPQjMig1LLO5okkT3b3/yjYvI
XaIF+AyN4r/2IaXsOiI92d6LpGMLM/LViA7xoqeDGmdwCymqlMppU3Fd2cU4ob+IYjguud66m5uF
SENtwH4nQKxrIhXPV8FhUowFCXt7taDKnfbYwgiuGTx32yCmLzrOzEUbTptQYSxnZ+Bcs7IWM14B
hIl8t3IcQp0OPh4NODWv458Flsgrmc6Vq1RyzBNJfu+III4bnlxZbr10bfaBax+FvfWAuFeaZdyY
RETFYPUWpDBawCdlspsX9UABE5urrSkLU903lHRkMszhwwiVBuSt2ApmKNAOpOXA0N+gHJdHM6Db
OGV+SRUIfEzgXRjcmKBpcZrEQHtnGKLyl1Ru3iNYOcRzTxLMJw/nAwwVkeATM0lCs9UMoXPkbwM5
wq5/g8MCfKTZOskorT8l/DI9ol/DsyDHaoVOi3Par3uuUnHEcfPePDI4IbCHjMkZRSzGlb8XKMjS
Bsb/ZJEgsyJ3+D/Vf/hYZizIbEXCZUXDpa4bBStPxSjIrUixq/dD3oO5gbZD0ZjcUhI9Y6lflWgP
3w++yMI8lcDJJwOOIAYnfILxqOhOIbqniLu1elvl2LGy8PlaqhpLiyY8M9L2bUsEbNWA7Or9XbKO
K9ZpEqB7O5OIkgTxx4pbvLP7fYb0fJeD/TdfWREpwzC2bCf0dvV3zz3JxrhnYetTN1CSgZo+CoH0
i7dBzS46lUXaDNvM/OEfdMdQH/gs0HdzL8j+tL/Fkc2tVqE2IC+LiBMNruu5o1rD8MKCCmEwX+Lv
yRWDDj9gI8wfB62X/1jCi8FBPIZ7/mAMQNM2SdgnF9T7MP7f4ok+nGRbHgHjMt/Mxjt+UUg3j8Kj
kePZ7L7sqi5PzX+vTrYZGHfu9201MBY8bcOBd5L6bXqdByVOqovrsQdD6InF3CmTzkpVFy5TMWtm
GdL09Gyj/sZC30mxRugpVQYFqjQnNVKHnMYmo0C+QtAqhS/rKxtJWXLI+BJndYagRFo0npnAmpYa
4f8f2LqWOUXGEhzce5kGiKmCokwZgGiQL9owZcGYps3Mce0gE1nW55Qes3CNzJwn7rbMoHfMKOGU
W3zYTfH5isKmDpxec7ys374AM+Xx4KIObUiowlI+jEoWRyGJgN3g2kUS8tHh5O6uvm+rDwFo9Sxa
5x2pxt9yTyRRHbqcyiTYls1BvsBvxflC7ZjRQtJYfXqXma76+Lgud/ZFWqDhvQfeDnqG2d9cGFeZ
ZFLyRdXs0wR2aOiihRmIGQwHeiVn65xeRCJ4E0ui9JnllezE0ABS53Sk4edLYE9FzvVJxEBZZIHU
yVMFVXickqLrQ6tW0JP8gUgQmqzXiYWna/f6dGfHY/nN5QzYY6uJIYY9sX7byGaRDD9msHZ9bv14
TRUtRGnwEtfH1xv7BFCL2/cHUYZi3Plhpo4iDuau0hw8asM2+pK7TKqh96FL+H+KbitK3PnpX8RI
OLgt3XNMUAMKHwiNVQKdo1rHblJ64ZLsNtnOd+grztxXmI2g8uvhI9seKmBKo5KrSWoA/raWX66c
cN9BHzDuPHmiWeeN09cHV5A/0JGDmG6SsasvUQqxFKswHEbMh+KSGS/FaivZJ6+XBt0dzARZIhBh
VJ/yWyZev82jYDVVF1j1BJmJ9yNUEXomO9EiFtYzlR36cl3VNedQYab6V9+jGKePcqdRBwTyseMj
dfty+lsbdVsHw5QKg8Msa/BAOc8CDcHg/MOQ2oWkBKaCSSjAHOYt4dsHQv0Hc2hb/1X/3rGxXwOL
b0B+JkOfsJZSCqVsKHSL9VYK9KTgYftkCgBrIHy/pqjz3rLXom2IY7R1e3fE/tEb6EEH5qsljbvg
P1lnVThlMRYnwV1AdDdpRkSRAe5LETX3hN5PBrF1JSQ1vFutnTtSOmRdNXlt4nJ1d1auwIPurvDk
JJsI2NSXNKaO8hxndrPAW+vdvRx+JPhpBM3sP0x+SiJ8Tt4I3NoWysKGAbeuqmsUSu5ctVTusgHJ
dLxmEg2OeE/JOjY/oJMKWUOWFvoWjzPq73sSeTGGnlae9cWmCOAmMHqDQtuS5v03oC+m5lsea6fn
yp72/4ukZWHUZBCs/Irl4ZPuE/jNWVegA2TiCosbUGFBZVdwdiO+JRZA8PXu4gb1sbpAE2ayE7ro
/YPxbqAXkSZO1C5t2V7/42t5vWNJ1ao/OdMX7J7gIZb8aYQhXaLTXYteqvPezaIpY62j+UbY/u/A
SijEf6koW0Iz5wPH4woJ7ootNX6a86n2ytFbt5kzIPmLaRxPkzJfH3CJYT27g4uyMyHUwGfe/H14
zoSeLHAWLIUdzaQse5ncaKu1kBEDZVr9ZE7895FhPG9klHGxAUU8lUjAkFXjtNMMe5BGXQ41gBUo
FT4DgoINFllzFp6Fd39HmMvzpOjZWqG7vPjtLVRjeAoUB7Bcli/0H0w/G927yXt1XDvN+gYN9Gmy
1OCXo8wlPRjx1DZvxbw60i5ibYDggj/CW0xXu8nVhoggjojhKKSSgbfcrMm5SPfGLJUsyMtb2iMe
gSGEk9gLiHz55udMrjErSRwemUE08gYRxb7yfQvHkEVF/KrerspEy1OGN5KciEEarxx3+QA4gz69
bYKfbGtVHRGx1ZoNh49ZYJrRuuEVxAXqDy3M66eNYY1mMECKHiE9ae2Jl9rtcPKfB/NSBtfj7SV0
b8QkuN72m6b8WEPVR2qu+/7K3L5dMEeS4JRAIzIOCx89Ii/zG/bpGM0N/9Diaib5iZdiGps0m69/
G0LXbjYhe7muzu/Zrcg3RZkyV7BJv/NU99BQM729Q2XFGdI8hNgSBExACI7O9x6DY4qWmstYdoEy
R4zfoeE2yPRDyFaIHCJXJW7xfUse154K6LIzfzwB8+LGx5/UfTyu5oDMZCoKTrR3UcggncKRHEDw
NgKkDW/Bc3eebwZPBPL1QhKtyq1Y7U52gTkBwyQAxPuZkSa3zRy+Vq4Hl4OZtNKVMOebylJG+qac
zxS/2Gwvrnzn3B7keP+mpzof+YoUH9UtD4oN7e1M4DaRDrgq8pX6UG9qXwng0dR6dbkqaYzkjK+M
r21fNAeo9DLPaweSLivmdTIzNbsuyVfRb/w3gt26W8X948ti0KUBwsC6kZQqUNM+OxwDAiWfFt8u
PIc8lc3NNhH2p9oIps7E5a3bHHK9uHJ/9jQn/Zmr+A/GX+hMinM/l+BXuJ9L2NlZQmcl2UNGzvzE
iFuyCrf8Az0uQYOrh9Bd8jm5G+P9ibqkw/xyaRnHOl9SC0QePJI+ZX+eVEaNVu/Di1IfxD9NiMIT
MoOQdEHrWsRmMzeAaIoOISfF6xK4+y1RcrfgDKD1CWtj72FHcXyhdAyrMYYPheXtMupyev3rPXZo
l/VWa0ZCY1YkqEKqVUxvpTWGNxx/2RJ8bPSYW0CRyZA38EaaFwqiAOq1iZOLYRDvUFcGS+BoGjcI
8ppQWPV2HGFkE/vEpbfqmsKZS8aS69ytuS8U652xkMje8YJ0XT91NOnFzC/s5ssg8X+zAoMhXWyt
NyI2u0NOh3poOmF4Pmm0E8UzIPVFrdU4iwwXUcW4B07vaMo8vEesyZCgYFlJwOr3/+MQFQAwX/37
G2xnbBR1JEtZxjvlAQVVhz6ESJLYUt0yX+QQtBxKFMf2G+lMu3LqRvIcpXVhkiuHRRVz+gf43uwS
uCOfopH79kwt8b7N/T5AbenCDR5A2z+LCj3skB8VR2icvcmd59ZU5JeL9RoGXVyg0ekxFOlcHoHK
+gvABwyvP25VCZD/ZKyRAJB5q8cKGS1o0AyZcMnnxm2d1eztBlh/XzZqHISxg75uKYHw2JmDE5sT
BDRk/94UoB4zEE3GH6oZryOEj7ygz3rJjAIRCXL19L5dSHPddo9ptAjKcc5rGhn//MFjSszRLgF8
yiOCeXIiqVYyOhHaf0Tk5nDHW3IlRNvyJKm/vb4bImNSI0/7FHx/g/LyA01HNWeMVy1I8bfLJ9EP
AKDOZEaMggjHpYgf+W6d4Sg2EOUx/wrMYO9gpGJl4wYGLlK3IgJeQYMEC1NBN9m9/6p+Q6v3KC4c
tmX8Kl6QM9WScDsKLJ4nsysNj5oGJvwzU6fPP6t3hm6YEXLVinhs6b0VnhwNJdYQOm0e87r8YzZj
n826RD10TwjHjs6psi9Wty32/AEwUGDQtkddAHKuPlEXVAnpXRoMeMKz95rWQmVAKbYjreuqTKbv
OJPKHI4OX3qNN/9eWjSC/DWrUi2JyXqtLjh4Lw5Z0eR7ej4TnplL1wbEmpZWv4pYIcdeJv2ckqOQ
NuVuRLfwY610OLBOrAjypiF2cdqxMW7Q+tHcuecA200x8b4IPC/ofFVbnpMDORZiTz4UbDKtE9CN
YzGBlLfSDHQl726rqvm2plLBKkHu0lqkj12NA91loUXaERMGecuotlohCJiJ1mZgwwFQxfmhk75D
mNKUiKGmNbMv4Et3p+Kzqet8wWKFumnsm/FsBAbsDsWPQKJDUO7NXqsQqjSpnB1vrQn7V1YUtFQW
OgH/GSxoS8hyHLFfPF134I8dzLzBIK+6JX1cBCjPmjc9/ZLfXf4sHCeM+nDwfYR1lFuLiFrXmbzt
GgqLotHtK4fhx5HgPRjtDEYH6Nk9l3OdieUU6wta57HBso/NsaZb7kh/NiJ/qRIn/Dp11cZQssF2
eT/A2ZjWC55M1QZhS/Fnf3HAsbrOPJCwKgjZRE0e3hyThcqD/Z13uM2O8BI7OBYKXLlsgiVXN8yg
pgw+z+0tWE031HyVkF5NI4Rh1kcVE4Uj4Se/SbpyKWuPwob4OFMNiBeYR0ihnjH1X5cFUjyJ742A
u3yZTQMNtP0BuHzp8d0bN2D+27px4cQhShgPALDFYM0QJb7vlXrRPzGe1M4gXq2Xw8Yc4xRF573t
V24VXonMopBDV4In9QAtJ9xdX9oaU6cuUJsE6bbz2f+aXb4eCCLe5Imx8TYUI0cl4cf39F18GE7d
/eopVNFjsgUFe0pFuN6uJZWSswclnAQCEzgMmo2fbZPpXpuEJsuEErC1fiLhmElLKUoHdnOIHj1A
Sy7v2yqMCxRHur90Y7DbmBeJQhSQIETVqdzht+KTouBvY2GSixtMaa0njjRyw1IvkjyH1phZixZe
wpcvN9BzxRyMmHhdiogI86PeVVNrZ45dsz2BesNjyZ/IbKW0swD77BVK2MYEL7jKzN6jch55fltu
+40e6N18kolc1LutjwQ0YYqkvDtVyO/KMbBMZngkNO/4LOVCeg9ngen5LLFPbdlgQze2mSgGQEjz
PvbEVMaPGY6+2Pvw/yT87OIqheafb5McyNK5Y2Iozuk7htO/3o144mgq1dOQEIlhbqt5F4nQO0j5
3OCX0+QAmtSyWMhc1N+uj3fl+YhOEWIFBtY32KDOEkvE/oLkW1tMAPimkRD1yIZXU1engn6dXiC5
a0o4V14uY6rIAz0yHh6Oul+z485sHY51/fWJIlT7m9uT0zl3RpUYoK7DPF8SrQl+9nWpPrJ90tfo
BmmksTAW9e5DqaJlqLhXESJDjtCocjTnuFNQCTxMZ/4ySydWSn9aaVwZ2D1rpPRS6i5oGbhdKV9w
ygOy6Wz3qPTxeIGawHg0oAdkaXcSn7rIDLtXteRf4noP2uI1YeoOPxcJPXHBXU6QYbPHRv8cWepN
dRjN9t9HkgM0SvAlok5HbPPJph3yKzwCUYNNf0G0ds3pIDPvqsamtkq8PYc57YyWcKHP73OX0SCO
QcfGCsCk0yU+Q8vaqOXeWMY9SNNgPbeslnRFGDe+azVeJbNqbbBSvyHbgXo6LJMbJxOwLcJatpER
AcsvLlx1Hv6C7puGiaiuUsi4xKqPqbyB5t2ZXOB10lG9Rut4mfm2YcSJRuzBJe+avQsSsqmdMw3b
d5qcyrs0gi+cW9eSySb8WS02g8RsShu0fpWaOqohJlrj/OizHRWns8MmmLQ8O4ZJRNi8WoRZJNvF
nT2TrUWDSLyIZ+KoGm8GDvASSK/qkTpow25vVYKmYpyy/BbR1tP+7RHCM9zFGKM4q2vMW0wtvdg9
lF9IwUAH90HVeuebsIZWI+dovoOTq0P6qF5hyBl5aYtWL/SvWtp4ObXSqS+drcLbk/vxb+bNuSot
A7Et7Z8ygd2CrAHPj4mLjl0UDbGkErI9xIrVbS4o0Tchlw1ePkCsI8biHjUlTZm/1RxCZpAxEEKY
e3Mf+1lQjSOUGC+GrdqAUN9emRXhj/8ue0AQpVHx+UvmwmjnDEKubG7id7M0tB2ymc4d+vP/qFF7
x6M+RPgZbqOWYK2Xf5BdL4kEUNK0AlD+xdr2HJSbYEAEW/scL9wUYSUcQ2tYg+XOSlv3m/HTEAiQ
kNOgohTvHXoeUFPUyXTJzG/jRCVfZq9rN4544bGlC2ls92DK2NrFSX7mbQNDWYdHmlT8elU0EUyX
nYsncrYycaI955o9OQZkAEdxDMhz0cQJVaNlcDwvXoQprWKbcJu+Dfc2W5MaHYixZNKYIUB73MEz
W4KKSefhlSxQLZQSKqBU8MGR/nLMhu8YS+B5YF4ovedlvMD2xdbJ5X9lFqO2E6PAf/1Dj3etA2RQ
gu8DPX2x/oI8a3UJ5LV332Eedv79mcGqxtrRMbaiPi/FNggkps7ivhNJS7UjXKN3MK+3mu0Z7ugR
+T/QFfQp3PFc6rdIU1UzOChbOKaZ75Vkemms+Rj/84Fj3oazrxSps4QCN5WgRC7EROxR2BRbQ/Xb
lRQepkS1LAYmMHurHeFixtGZqkGKT6f4/E2TO85mJFP+DFVr2X9ns02xjlgH/Ow4vfF98k2Fy9IZ
Jdh2HyUY61aD1y6fBoDTfheIdxVR5J1uF+VMLCXR9nwNIcnRgX24eMgZOHc5pv71PJ2c/R++pl2F
1SYpnOH0ntxFVrsMLVDHnNpImGnJBSdp6oqR5Eq5FCBA0AKnt5N+j6ZsrIAn3KOGfSTlN80czHpT
adevNPb7ScTDq/DhC4mz/WVM2GTGAOnU966/K2ibPFuEEZ6qZQ730c1/EmoE2y03nWn9XD2zSKdG
kX3H16QvgzatWre7Yfb4IyTSyHBmu/GFk11+/eQvsqc9Toiyc0ef4na1yVrLm2cvobRFyNXocsmQ
CKHqfcHfcsfhrnTFR0vNEXeuZ+cowkxFOJ+RYc8W/Gg1I62nCEjpO/GfmK6eJHWT/aUPpxfWEwPx
WOvxEVirCCen1hwVwbeBrNhj1RCZw6gMIfnwrLo6GrV+Yitcguy+fLPCiz6DbFfPDm43Rb2MGyI6
WKh0LmX5N+aah2r1pnwy/IZjtYWB3qmyaKvWwfQcSvNKgX0idUcl+E9uPELNUs56+xYhGNrD/Cn0
YtbM5RML314fSSHiMl//rvq3d0xra8ZRp1ibl3vfOPTNk++X4nhg5yoqRwFbPUJSWdRoUOEgTFXw
xkrWSRADVh98BsxX4HuH4eb0LLi/0N7F193QGxhGjoxSUegrwbv3dRE+ggwzJbRw02lut1JM+9lj
2ecKKFlqE8Dio5GHT7sZ6P/BdTboN7HqHU52mQnI6XAWklFxW5tS2hzVk+96YpHnr0Vam4QR4ABQ
sEtiy50+DuJ1Kb4RHt7IOr30m9Q3r69KeUJ8BuqX74KeWs32wCRRsPvAkxyie2IsuD0UIVas43Qc
DDnJiNGs778YP8qpp7OcyR19/UXb+se8jCYyLSvuHnqce0uSyDIc9R+Mrm1D1IlX0CFa00zuVj/q
K2IcCFARnPZTMuZGd6mLjdea5edzQmm2/m0rrzYJCg6Bhzzn3gkhPFHopHhDXoyM7ihdwGSEU7Ih
a5F47UXLJjoay8jMFL9lGlfNW2cxbWlbEgZQb7mrI/FzewHr/AGuCSQQo3qDo1IhVDX/LaUarUdc
00y4V7EDe6Gu99s+jy3YDK6wJ6aNlp2+/Ut+ZfEU6MBZxjdcohVkXFhVxiH+zkx+lPMpAshlc87Q
XJOPCRIiamRJbo9Or149EThShXBf0cJIGlo1SveiL0dPDd//O9K6FmoIvXSLPV5pW0D9qe9uWNhC
HXb4oFwDTnh0YDnp6Wsy1o+ZfzuMWWc9UecgZt/Wi/W+20Dzt7S5HhLmqbMxK02tpl0zOtVhLLDN
s1GK/JP6Zj0yYQgNjaSUYGkVCFbWPGpiYcs3D2UO2QbXrGXCqEZFe5oyCaSYFwhGP+E3q8OtYP2q
JFjgZBRYl1q6VHDAegxr0amsoMXWEs1mlgYk66VmJRivr1BZ1uTcVsbJ1DeShTaCSMs3K8yVWOze
A7pwCggcUAClZ7THNNniGbkxHsTAokd8nUCcn5K86bPmkHLfnWcr8Y+SVWQjMf0Q3WQYiDq7AmnZ
wH8rl3tjElojkk+pGdtMgFhyVv1E3Im4HqGcDhMe0mckuJZ456xJBUYzh3s5Yus0TYEOGZPqnnqY
idl570NClLvkfh6o9iz/yBcHetFz+Jdm6P6V8H4H5q3yeHr4d63k3sc7E9LN6KKDi6tgwhzvFTfw
bbyaKXnz52AR4oVRCmrv0GPpAj2JCvkXS/H1xpGoim5BfGdLD35zyAW97QCvWDfmUB43ZsZ4EAgv
vpYdUIxFkCqveXZ8ec/5560GefJv2lq+EtWP0m8QHzaN06YI4TFaha6yVgVQfrUiwllPSIr6vtDZ
YQzApq/cuKDlk6F8V/Z5Ctb8tp/+tUWskeA0RoyX5gTTVmEj3os8kakNCPfCePnD2tt9X6EXmGX/
/qRVBBoXqRICHxU2BzzvQB3r6/qegyTvxjQOWvyIHgICW1T3xrxoeqsilrQn6/3Jk9Y4V0e9YU7G
93jQX4i1V81gbZDRX4vrOecGv7U3Sh6QvKbPMWT51CDv/AsqPZQGgw9cwQiHx4dhgVCItofJ3WNJ
kffnCJV9Ys8eA479k9v02lDFeQ4wLWg4Yp70e0Xhy9clzCTHGBzQMVnwuPYfGpddj1GLk6YRSElh
0ClJlxrK3VjwX1FKcqtS/cWPQTglooHrbY9CIQXVa4n9A2ndnnfgF6Z+ZfR4UQTLYT5XcHNX1x4z
/cWRTaXmLlVXBrt78sHGMjdUORHJST0gTG7Zj0xe2KDRsZNG2XQH2oeF86OpiHTjdHOwvuRPtSpW
t+j3F125mlrq03pnIuT+Fpe8upBrOquTzBsjupQs7Lf8D8uQ9TDZWqP5tC7fsP5LXGO3QPtwmFtG
6D31yM2Ti3BUD2x/HoPJ0ACeUhlYT/Hlr4lZClNEoDOkfIZQvnc8ZhzPwUiedtQDIFmJ7IIxC3j3
gr6uwFoppQ9lFz3vMVbc1zO/s/Q6wvihQeW9NVm7mbcRjVJwPO1z6BT3tgA4VQlG3NXak9AiR7Qt
OUEmPwSMJTRqe27oha8/35bXA2o0Aq+jQTCNfTPFkcWTSg1IrVgsrStSyQjFh5A3IPMARVpgSGhl
FfmSxBfpGRZgjP4pxpH6jLEok1KKYPoWem1alpSoDoIwx7NFau/lzxy/P2kMl5wEpolAJsDSq1JP
7c9XumaBrfZjN5UwUxJl5gtEx0TAErh75Y0XkkX1YXMv+2nDM7Pak3rVGKyKkBeuLFxNjxgWbxqy
o6QIg7J3gsTgkWIQeA5CvKtTdFNzdih7eGy/pKKdW29cBb+pWGksf7hbIlfbL7Rku6v6I0upnDQp
0fUQY5DhdzkgoFBXjP2wLqz6ts7bY1P8HaVJ/xdHIZ84X2mur8RvRLigdgBIT9G0XC4yu8BPu6yF
qTBS4XGBTI8NP8W+dIrvseIh3gO/0Xi1tn+sqSEFNdHbWRntYdSiejMK7QhcYzpJ3MvPjHYZXy1C
fjgxOT2ZeL29xN9bB/5BD0tNVfNhx0fNYhbmC3lKgHpJRb83bYF5/HRIMnf3HvXGxk8mEtPrUdY+
y5bcOLlWrL0dvS3gu8OHDMP6YyJjp7q2D6ONvqam49yIrp83nuOveba8zV5Aal+aGEyuB3msETiG
e/MU/JkRpxDwjsv5DL1X4OnNHPrz9fRavTJg7UBuuWzRmDXwA+GtpFipFn3TH9mUCIeuEq81K1t4
vnHp+fhhlz8uWgWbSpc3LfvTF8e/q0GUDN0ZdngkdXERLIUq8DbGIqjJxaorG4xjZ7qlFXa2CTVv
P3lJT0NmN5U2Q0mS2ldzTkMgYYEFedFYVUrCsVagqoktRgoDSHcsur/Dk4nZw9HX5EDN9qVer/jJ
r5WCEUJBE3PUX6xKi+vOL2e1sQzA1/NzApMUR02C8psChSCbNBrUMLAUobPYYtlfqQTPYKxJKq94
U1QZBkc+TI5+Qd2U3m3tmy51kqaIfX+RJu+KnkGs2Qun4MVUZiugCFhfPrSS0aSqn0a/fCv00fmm
Jo4Hsc5QtlrdbPuqLCeOMc6J4H3TKZZDQCXHxZ2uMTpsFnIC2nv4i7ICl27Q2XhiMgL+DBoRz2ud
5sj/uGhQdtEX8sz0KXseChvi1L+w0Mw31VCqxiZwC9/og/jzHvwfqmOh5+HVbfqEtRFMZgLsxHk2
v8x3DSJs/AwP9Hjg3j9Aa7JFwDmv8F2KlkxJrabp46bXv6gDueibbZG4kPRimRWMEcTv7B3GL8TX
lu+XTfUdsyRqQFWQQtpl8WovLr0kxN21iUg9KtkNweVpf/sgD6cfMmyhXc29tD51K0ITYbtykxyB
zTIYsOmk3LAFIG8XtYM9shjoot8gkOt/KM+4kF8yt6XxunoYTP1eNEEeRIWdYv6Xu6vCyM6gK9Bd
EhHO9wo90j8DNzfUNJjuGXRqBeMgHOB8rW7Y0fV7pqb3wJ2TLhbSt6TVCgSkTj0JOrSWaBERT5QN
020nPnPHxKjncD71f/oZW3gGC+uxAPTeVb6jvb6KpXEAIaVFYUJ7JL79xlyhkYfI5vi8DpDA4f7h
CTXwVv4A/CB2QYEMEAzTPl7VfGkop6PS+PxXw0e58SKrBu2SZPBHBT4poxxyN5iYhBtz+IEmVSKB
e9sshwPIlLb3K+XS2GpkPnOyBLTavLSS22AVZ7gOAajO4FNs0GazCtjFLhul+2yiTyPbsGS35SrY
Vv5utB2nSBvsiSzkThiyOQmt9KAWqxBcVtiGC1htt3ZmVhYA0nIKwD2sxXLID7IsUk1ocUts7xiu
B/wt0nHCNLP7Q2DSwEE7OZp6OnIg625dMAptpwAkoqUaeVpCcyZtkr+5SMwbZKdGNudd7FSOwWXH
0DVNVuOIk8n0vJ9OboCDCzNB0ikyne60kHVT1rlSw67RlxvLyRUyYkN5S2G4LxpjgFePB6AZO4Bw
iZwBChqKaKkaOspJIMfrMAUtv1ij/KW375CzRRemS8eVTHQ20yL37g7ttEjDEPNeL24bSEQ/kYVI
oAZ6+zxxtm3n1CoUfy1na8ahlzrPAs7jJSwQIax6m/RsAoxn9e0ItvZXX1It16kGnKGycPNcc4mL
3ksncPnbbOA4xWViIcOT9xeLJ9K6UF6Vifm8K3ZcllYr5NOeYOba9Ox19zzddYnJFNnu7QcTrCJI
IT+U6EykRGEFbEJJFfjCSs63No8d2ET899y7PuxmTGZSMRQoV6keYHuM8GQZsEXc8C9gqVHDx3Q8
x8+S12oRr7Cxr5ySi+nFwgu+90CZ/vRz96JZiUNhdHPQMIh6Ualq+WLg809v1c5Voe+9KkgsOW1X
8mje7Dj1lqXdGYbSSasw4b1VYQs78Pc/Rg4XEkND5dvHaczu/uzDayowcb1B1TUW8E3bXFyXvCVI
OF/HqYjczAtSmq1aOesAX6EZsK+L+JsazSfx4MDCjExC2QjSatd8BSKGQgPyIVZ2N6LDvNJeiDA8
m5N3NGoMX2wA/hS+/3uAv+9UFuUAaHuSryL8KOeKRPUT8a/uWlJQMnAJa4m2gICko0OekvV6FGd4
vUxNlWdKBpMauIVete/MVSKGQXWg0oZ+kolifzR28grRKyzJsvxRKXdx4aFaPmUJjn9YJbsgtPvZ
6jxOZXvzOUeqP0DULXyiskfpueW9TW78kXhohtPay/rehppDII+1o2CbDOeK0QerDrCzaZ8nHf/e
sfSSf50DI4yaFd/fmcTQcuyGfbH3IAKTO/iC3MEWX7NZfY8bIUHZJ2VN6noGNO3DDK432n1X9ZEd
jus38yh5xZgvJy3u76X7KEYMmwx+qt4P17myNP3eDSB4SDY3Q7uj1SIaCKQ7n3AtlyYuvrrzZ7Xt
Ck2GwLMf6xpgQMf30eAUiAgylxvKagUAmCoRVMYTQ/Q5yla21wArfKzPlM7Qeowu9mYeCpiYd5VY
m0UkalhW3c9j9FbGatKdmsOugicV0uoLSByy58h85WehIc4HtB7xFOrqNx2PJrsqx3FpDlHN/weo
aoh24m4InGF/ijXeqhyWFwO9SUiyb4hGf3kCVEmcSFK+U1+ri69c1kOss//OKi/uPYGIlgkbRcFZ
d+nL9vW5UoLMiQaQtS4HL1Xa8vUDvuyNCv7QRyx3rgJch/L6BKTHanE+9zCTrer8O5qlXBHtXcj9
DOFRid/VH9vybjAQqO1/rWFtbJ+k3smitWjl9eLHdVn48RLCKb2C8kV8Nqe6vIL4u+oQHpVpRKq0
wfIQDPJ8ELrbVtZ/bd0EOMRl0aETjusG5lBAOLvkrPa/L0bB6OMqrKXMnVhJWDuHpVvwf/hM+n2I
ZI98mCYELWBI3uwEjMQs1MDcG7H1T2HVHikKUc8OAKeg5mwNH7YMiK5WxKE13Sv3dkppxtMtUuen
1/JghwppBlk+6oh9p+tdXCAIlzY6oCATQsVv7yLNGXDFhkMUQTAYKxyQIxQ/3+LcNCgm4Ed4ECRv
QPXxmrvYjrQClNYuqNIlIVZi7FNzdsSS1VdVUkahCgt9sY1HTCFcC3Fl3NHV6+0abK/qvNVQAjWl
9O38HET2uLF2Wb5m/dk1JRHbHBFEQIteu8XUDog+xhJewD7KUgSjW/iOCs86ci1nTbiiyVEe5VBU
bcVdSRzBWOG0pnNBfYmKoNtyMpvKKJCLqMY3X4Owh2dHtJ34zYSiRowxtNveAD5ZR9wSHpV8gTlO
ltmOERkZkARPacsFE3lCdh3kH3ACgxHsjt0t03aL/VAKmppEiGh+g5Fov+h++Ua3qkh5S+UReoNJ
xgffDVg5YVfn0HUJZFo2Nzf017ieX4OC1cTMdrlHbFMuDGbT1bivci2gkyfVBCOqibK8SWW8FNIQ
3zyEZpm+IHuOSXmtiSJBXKDtBYakMBD3d/J/tMNwiuGuEmbM7gKutljIoXvaaZAi3daIE67n/IrF
qgvuzmGYd0vScZm3qUkeu0+oGyW/kMyVmpA8gTBG+/itZKvhpyPsm5H9rgPFGWaE0HxQ9Tkfay42
k2Ap2GQXRRg7NL1bChHyRT4JktOk+P8eYyL+7G4QacaqkvpCBIbLeWM9YDV1VmO3BX10RLUh9B1+
S/t0wAvddDZWvdgCafJaVDoj01xaJ5ZhHvwt22XBgFF55ywIjP0pG0PvLHdhwEfPw/zJCfGr+l7m
TF5TquA80KnxW2+27phs2ptuQxuYY1rBiEX8b4z72o68FoqVoTBdKTPDYMpQsg/ERIi8D7964h+n
bwT6WmDhHParUYJ7XyDXYAueXq8gqTrD1smZAZLo6bbbhPsrqz2gtqA7am0l0G27PDoCichc2QqE
8K1ysxMn053DQBtmMf0qWSwDB9SNEW9l97uAdMpvym0noc2HF9A3/pYrItS/hcjcAIh4jT0yIglM
7U+HVo70zeicbJWwgk9EEDfD5ox4DsYZdjEm35rM4da6cID/UbWo6ZGomwcYwy0nNlBAke5RJoKP
esnZmM2L2E3c0Bx48UDdYYIvMtDtUQWWEeazqAr+5MlBWvGjtR7jA56vzAfoJ9Hx58Owl+IRNdnv
J8NxwkHlANwiKCWgS0DKLxC+0WjZPbyJoMwGOVCEb/uta6SjDkHSHsjygq8FNi1I0FkFSloIQrvr
GoG3o4S0bqBAGPOPsTN5xO0fWDREkhEna//oM5v+lvf/PDNaJxqykyX7NOZRr6LKVCrVuJ7TRw9h
BSzeGm2ahfmn/In7+olNLBsXA2jqH9SmDIJIRx1TK2x557ky7i2A2GLEatoxkFGeyHP33Z/PhZsF
QU/CvE3FDcWnRypOqoexuqH6Hqo5msHuXIRiyWEGN/vgNKGRclFcxvZmx6KMUiSnoLIQmG37FGG2
RYgIwLwGelozTf3GqgT3haV3v09+KY8OWabWdaG3TzQED/XFKi1PGTf/mVHLeZ6aJ3wACuKfTAs6
PHdJDDGiNmwHz+cgAi7yk+gL3SlF/P2uFqKTEPrUhk5vPhnFhfNFNed5u6ATrA5qOBtFt5Vo/an+
rIR/fqwlZ4oQoyBjKT6c+E5LFlyuyD7Qvz+f/+eQ+WErr5PG/l3gmZWFRs6hjqt7IhD45QlCWeZC
p4KdUpIcVJRFAdyvJntWJKtuO+/pWsCq6Sh1dCO045AV80GRTscChTOCYh2uUhzUj75jRZaSfj6C
wEH6oGcnRvI4fFNB9+2fjveHN2RM8AC7LGDoUGiGfW4/WwzCAl78FElb3TrJo8iWf5+G/4nnxF0+
SCg2Ho0SDop2orCu3UJlM8dFC+MuTTLJJBo6+AwhHRlmbFCBf15vj5ZQARlyeirYR+XEsBG8U6CS
T0NRdN8nHquzyRMjWdkndIbGrgNZnGx60PQwIx3lramsavWbJuz6bkIqgrSs+F4ESoho2X/rqQqS
ELJi6qcyfSmIBrIsznb6d9K4syq7o7ZmcgroqMWQaibixaCg2VNMutj5oWvQzpi1jvXhm0Oa4Zy+
7nRYDvkrBxlwwz1/a03afz1y7J29i96Xy2QbdvaaU/pMlf77yWmJu4TxRdUQc+OWkRybflCX2wDY
Mx/zrTBiyr5rwvsbn+7nI/FqrERWFNzWVikKQ0oT2LF17enkWv0EiYer8fWSNTLYXfWh+JCEYF+u
ks+IsZZPl2A90Tz8Qn5EHjlo4Ph+o0x2How9nuydnmEmbpH6vvexh9EeV1iZldThfHC49db3uJK5
xZiVaCCnEmP21k0/U8trzr2Uc8OcPplc7m30k//4bpGkTbMlPIn9e5oyNEsNDkfa7J6x0nga3aKy
UDI7lj/45xj+XrFFxsm9d4KxJvMS/gCwwF+1iqTYHvx7lPSNvyZTRGSiIJ5b0bppkxIkweD+k82/
j91vAgZR8ajyV5HD30FUUyUYoAt/iohkFiLT6jZW6c08PF4lsl0qzRRTXopJOxZKztOsD6aFazKl
cLssena35iqzypMdegzbBfymlE0wpDZpoyMYhU3Cmur65xrsrvboTOONGSh7Y175PdicXUwVnSLx
Uy2nOfZQQL3TNjmMx9wM+lNC2aZ4deB3B7uaKQ24fh9Hb4tWbVsfDhC44OVI3v39Hq9DkIfC13nw
5Pr1EA3NeqKFLPfGvhn59zftSbfBgKiVwYU+cMRjsJS06TXIenp7gXh5snKCEdpuckBaMKMVDbpW
+e2Jq5kx0t3HHghZ3a/0rBkvhgJ6uMj50oShs3u7Ga+k2bjbndFG6jZhOar0y3BLudl7KyDTNH4V
chihdY3nbHE5wfjgeH5qc8JQZNVhkQym5XMNb63ga17I5nuAP5UrXsrmjlJstwFhNlejccJS9QsA
y9d5sYpf7qK9qvihPtdTavBPLVBykkiC6EHFq9qebSdAHzpR7ZsmxjKPbxF7bUXiR0osbmOFnfrn
IEygrlS902B2BGw1a6ya+adc6x4Tub5fB9FNUCAfIyuRzKvB7U47JKiyQ/0sk5WcN+kLNGHAE19N
CMIti0uLNiT1x2cAELd3XPwWHAnRUO2QS76JvNh0W5RHYmeZoriiODnzTCVslAxzYozkbA0lFKPz
KYE1OISjaMDCJJBtl5ib/cWuEHaPGZRMTFo7YyHcTZi/xp1lZNNf1pYQRX8Mx5LVNCnFPamMJpn5
OgmEXJSXIo0ZCGIOwpy0MVxIs2vRR//t9ltqfqode+PzcZKGTutJ6aBJSFx8kMcqZUaZ9HluamFy
MPDJlx/NQUlQpdlDEy2BseaWDWgydJ7RzUteRBqbzw27NfTvBrnDaNm1NeTSjj0bkJ2gKq5BauA1
jkcz9I1Lm8xenY+w+bjkUpzdSghro87Ws69qvq9TAj21IqyDjKsN3aku8zdOnO4t0uzfIVmoxZGd
CfJ4I80XaGWZGoB1fZKlx+mouUqPtCUDV9atsWyLw2H/+pGYexwMTDhJd2UgNhxlbn/f1JygeOf7
LSmCJNHCaSrhPlb1fy0T6qJdtShmfgtFbp7oeAAc2mx02NMavrfIFzSUa531QM05oVt3/b69onDG
ODePzwyD/QqRkCO+gigObmEpHvuzx2HHURjb7w08x+LY5i0rfUa9sWrlcBz/1Zi7TDwU/adfm4m3
DNeZh9791wK29Ly52ntqeoXVgj4FTnU4IbuQdu+oPe9JOW2DW9PriKZDCVh2Bgw75DnGM318PE8P
knq7B/LvLhnHWQ5SGQF1RUzQDPk+h0geTDLuMpDdwpwKJFT9uyDv5ggamRGwOgVMuoxUfEqK6zJb
4PAVENAGLu+3PIh/mPAQ9HLGO9L3sTg90wLZ8LniT/NJQi3qjwkU3fEbIJajLsON3vB8SzW6uWwr
uWuvZCQQzS5r/+UNJFhCQaJRRbCvLcBQjEeE/nVpC1Fxu4McG+1UxvDaZD3sbteK5zs4fd+dDTdz
u8dZS9mMVo0tY3fZU88TRXdKxpO1+2HoJEoygbQrLFbRg0X7ZBO0/2kUsR0Puxa5mmmhehDxPPG9
D+bKs4mQ9ZoCKOszBDWi31KtT26vhTxhwQFgL4OCFrD9u1aFx2RaGqs83sFOlqV0HL2vanHejWHY
C/MHZbbsI/jIV82pHuJy5yH7D+5E/6EGdXfFZ0d927KQqMjeO+SQs1JG5CthAhU9ZCgAKp0jbBWs
MRFVTC7V5KDjY7HRQpKfZo75LTzIdcR/0IJKDJfOBntbQecVN2pd626fg2pwkP1JAIZWmoGA9lve
GJQbmPQ3e4ptTjy3DhstbFKQdaEjXbK8QWn+25utcen16URMii9P0VGL6wgfWfUHVtYxz+qTVeW6
2wIyYZ5IN937UB02KXA2gkYM7Fex4PDqOqKOv5NTWGEo78ZJsMvPL+1SnZ+MhPaa8dY2grJuaNhJ
aJ4Eeoi+BVEHmawCK3ja57/CYoUdpm7A7RvYevyIRalPILzibWU83e/9eIvKoi8JYmsbzWampWft
HE2BEPe18khM0TAHgtwRf4+lpaduI+TQpbcyC6BGXZykU3iZ/g+Hem2rD998vJv4KrFjg4OjCwYx
3XCKV5e4Uwluz1WqaDMoZKMJ/q0PCYUOrV29x8Qp8Q09OYNcRdDcxVmYA3VEEDZyG77Z4fIuOLzu
9Fe5w40uS7cxMzVGze1KtiYP6DJd4HMD2FzVKLuhsA9g9aTfyXvZy2ZZO8qdWD8C0ijlK6EJdAlJ
vNcdIyFpGSS6gap/1EKskW+OkU1McfZkLwyISQUJHTiV7B9gGr4TjHLZ1z+ZpVrCtHLhK4aHD7pm
DW2ZO0pdF0iJJD8FtV/5zVgM795b6+tMC34j6fZ1GZBUxfUVVLayZ5WHbng2l4uA+qWlxRv05aTn
ZfMVKRoZBzsmdShhAr/3IU+VY4JPbfXA6IF/uy2KmuNprzv9ulO9uo1jrs9K8bxTytAAk2xB9ymQ
nR253Mr4M2q7TcFN++SXtSvtoD0dPcaq5lOwKNme406Jq1t9GejmiF6Aj7085E6LCMCH0fYUItHF
u7R29bRT57GX237T1Rwli9D1USSGe1sbcxPDvAv0FQLh19e/S06+4Caj/GyAwpZjGHJK7dH4Oe13
0hVsJRZfsIWdE+AW4SSKReTxipnT0UOzMVxoEGhSy46ZtTwUcIb5Aca68NzhxNBiugv62VxFX5+n
0qcoFYK0/P4QGKRDMxqSzP6q857OX5hgMdCUMPgPdR0tmnm/n/6/HJ7c0ZTdN/tq4oyoTwMIgjPG
IsUBbno0LLIfCWOrACCl+SBBnp1o0Kg9t/lIQ4Ubp4xyLaTpladiQSNrZE500ABzucww6kMUluOw
+kmQHEX1GHFO9cVf3T5fFw3sUAOspGxbFJEqMnMZNknapqkrV5Gpd+DiRIcfMVStOsMXk2Mez8sZ
uAB9b/QQF0Mzlo9bgiYyuxaPfSQaXv0pCpoFHSzZJrs1zt42UvwE3G4nUoloBIHnAKzMmqWMQ86G
bph5vbMfieOwswEGC/RJERnOaxMFTfBP/K3pmjBPnvR/2PIOVJ8ceFOPqGjhtXaj4DDE+NhZwgZw
AoUOGmUNR2PIKhlo/buvyp+k7PstPZDwpbl/NIUf0bO2JML4pHT4PkGCQEZXfhb38qnx8OuGLy0q
0Qn6ofxrmgXHDh7Hayqfqn7D2CCAWMwCmeCzcTgJkjrqhlUlLBUu6x/PfJhYL+B36Dmqp1BHUrDW
w/ABixu6IA9BX9HGA38feNzMm5FV2Kp9MkBX2IUnvr7e8ZztSB8/UwVFq5+2B2pvbZ2crnGTj80s
fgJGJmLQba8QhxZCpYFjPlSSOLuLNYhZRXRdtKRB6VzRNY3nw3Js9OseeYhWYAc4T+PHWn34MYfc
ssuUvBoqxuSnYZ3cvIEzOP1KGtIbj+SWVHIzAVsJqE/EAmiyCE94+/aBzR2thD2YCfyA6gxcgyom
QD05nHrRJ5md+RqpI/4sKUuUiAo6gvwZGpI/JesOKLA+zBuJnfpq9/fBYXFpKcEpZgcG9nzhjSuV
CVXEKQtna5SiNdXOj7V0nMe0kTdzmulfks3mNjFgwK+kV/yhH8Sqj0vWfJ0EnxP73OEFBqZSUexS
iuZvGMIFnla9HYfOmkveZ9UG6Jc5/ILe+9s6mMJUxUUVIFoS7mm0JqdQNC33nYt1q2rjWhzAibqr
TzVuQq599/WLDt6okuazXV9fMIHRGOnORyMP7QOoMfdj6WD5Bb52I5ZdAU9/ieKqj3AP3rQeWPQH
njIZqEOGKe76WRRzdVUwfJM5Jr5x53XjLToJQahA5XpmauZD+5a+jHfOPLrvx2ZOci9NVjKH/6jU
V9Gfo6tRoqvLGmDeBn987ZMJ+TldsnNpg0q+yNRrjmCpeXCvNagLfaurmoazizTFQSFaS44/lLra
iyMEXJZeikH49Qs210MmG3eb14ruYJq2gZ/97gf99pnD1AIzm5BI7BD1GJBgn1ius1FFAfueqkcf
f9qayqTx6btF94KzvSglFKiuUnnv+vv5xJXae1atB7l3EfebD7KKnK15yWPkCe/Hbkf30/wjr/YR
sYB3O/7tQdYsWJ+kVguhmQVDzqJEHBVDB/rbgYpM+wRXGqfAinmb7lVcizA3lfeed+L/w7Z9c84X
bqVMAGodidphNCa6Bqnlqzxt6vMD5wDkVbKo6se2R4P99hy2iJcBAh2RJ1pL/u+Pj7ahGzZwhXqe
383Fya0rt98jbWoc9UhbNsvHGZVGIgHp6WOJQahN3Kh5uE53uNpLyLaaf3OMbZc1LnW4JeUfd471
SSskrcULZuQJYNACMKYJSX83d3YSWa2qd8yyg089b5rbt5zWyv6jknYLQ2mEFhv1pDutmy4R4N0r
IOoWxvTSyauu1F0qPzLOAutUEmUaVaQ/DllK4QpT0LXmai1A/ee5ZJCgSc0bA8p36n/nHeMIBrcb
mbs/iIAhjj9UhsOEErlITnYBnF4MVf5xuKq801C0K0nkUS/PMlqTOyHeDPWndQH6juVGXLsbCNgw
C+ASaUkBPO/kD4IpW2XsGdOUv4yE8lKbIgSSKwft3ZoK2zjVHVIi0GjWtLCnJnJuutmiUclX0PdC
fsWCI/d9/SJICfej4GgPo4HqGVXMaAtCOnKcocaDxSsH68nlZujM9cdSQbjWLew0rGPXSYwyVhBW
oBN+aCkVp7VoFKPDmyCqOFsEscr03uZwJCVMYK1QYSvmG07Qn6js5ffPcCUgnK8o7iM4JG99ykej
p/rJtGJN7gHSYYJRQf5CjohLacQoFH8r7BG9f1ju/swjmJIXlJbyOvqXVW29orIkY/pQymGazP6M
XWKJbzm722D+4r6Sx22U2zSqvdDBEEoOfbUxx56ee8NOygtWk07Ze4nyKOM4ti7F0j7r9UOWpRni
9lXqO2X0zD6ARBWlNU3noLCwTTPI/l2FdS0YCUryUcbevNr9jL5CvmExofouIMq63zkU/V/q6WoN
klILdBFMhuLQMjr7eUg86pRtzS/8m+09Ja1+IDROQN/UBisu5OKP5QOEbDY9aMkvSB6APxeatDAu
CQm0jYeBYfi8RV6vSkDArIgeUrYJpLcRmDSdcWiH+191EX8+udy9RXjheuExDukeXf5zXBf0CY0p
MD9fchZ7NM6/yNSH+wu3xLQpBYNX8hRi3ARKvNXBoHRHQrQavqrcxIR+VTsIYUaxkvNNn6hYKSvy
SqMk8p7+7PpRwLdnZAvaNqP6VcNAIhSgLyLbpyJqs2erohYeRmfWe+y8yaIXDzsE79MJo4MMaZJ7
9w+jJC+B0yj+SqybgjuOwsLxn42A3yqSnjXhzQM7hVDmVPdWRDYn0oBYqnEGWrx6DJgsVIq5GOjM
n4aTUeITYZ6GKqzWIbwm2xUiotzJ8pXYTDxq7PnqxlHRB2j742rqLmAyAQgJ57kNpYm5QLKaZ5Aj
U6/dbOFqqwHV9ujKzGjegmd6/ekaKLBf7CJFCnM3dQvsoON6zS5qu+wO8UNHdSzANUPc7gVR56XT
pPHKa1SCKxz2XhRdFfvDRzh7HIay31iwUErFoV91R4dXUwIihK9UQ/SGpGVyMZvBauVyq09c4lQY
9ztWdy5wU98+erLqBFTC5kM6hlSZniK2jTeEb1eNTxrkoUBevpmLnr92zxFlglSfSIWzUzInehT1
+JOqLwZU4Rez7yrdGcg8iBc7srYIlJZAYDZzWdtxQoUhUOsMVcdR1PngwCvEaxBJObDjlaBDyfml
qpS1uslqVRMCzWiLn5q3oSveTOOZzW0rt2tcJ5Pthk+vGCm+2JVXZ0Iaua2YOT3iBy0eKOa0gbz1
TCbo4bVPXMWHjmhc6G0U9aNZubWk2d71Luudu4LjmqvsboH7uH+Nxg1oliP4i9t7m52Z2mC8fPsr
hP6CjRzKif9nfrfIBVOtV8kwSEVknIkMduuUId6oLNW3UD45AOmMB180/rhmjP/UGPyyOJtBaopO
U5yCvPPC1McO7vq/AJlPXHHGeJTH2itCOCyFerYKZ6+bhNGy+Wqx1nrUUKUVE+bo47apz3PPJ9DC
g1tXuG8zWQX/pl4XatQi046floRA4jY742nHCZY6K82kXPdSmWyB3tTSeQzhRy9jjtOFTSduAuW4
JoGRFMYUX3hYP1VjAJs9DUTObYdo0I78h05pwrbYdU9dSvePfsPuhub1z0PEYVhIDHwcBO5ZmYeJ
Qhzkye7HKffkid/DvKUXg0prrq+H66V2KuNCvVYMMJ1ttK69a1xFdB5sTMzoiZslR5smkiuTGO6J
RS96CwDN733mlKOo9hHgfKzKpsVVUkDpfChzz4ZOOB4Yens9RsFCuFdUymlfofc28Tbu0e7bCQxb
6GrVsEtXU/p4O36x32u9vDnDtzUh0/L+ZExnP7Yh3EOmGFi6utPee+fSBQZuzC3rPSFLA7mSOeo+
j02PAw71g+fxnyEgnhP1c5eNIwNORAWDSN1CvUswUjC18ve41cycrL1dHIKC6G4ls+DRRvesqIb+
J/KjWM3h/pF+h1jSZqOYxM3tYFQo3VgfGFKTK2H1vdOIFB3PA9xiOQI7u1aTj7H7jwzAWcYcTSoS
aqVgGsgqj/JERmQM/7TyztNJcolFMlkcv9cs5OhIDJvs+N1CPNR4dMSFFBdSb5uN5TzIAhAdcMt4
LoG/uV7JsmiY10luDFhO+EIn7R92t8pVQgI+O4g3Zibv3XjsoNuLwDv7AvnoOyJv8i0PKFR4h/N+
a6jKOW5QDAb54xUZ44mKViYRZEsEv37URPzB+WvD1TrgzRaojcwxjgc4j8Y9JvFG+GIdhke0aEtC
J3RJT8im1cJrwBHoxyNZsYuRC8IHIxuQhon2H0lgrQ7yBcnhQbPcYM8afDOlW3V1RsoA+9bV4+ec
NEgvrZx284hvSzPMO5djuxVSYBArzDo0WmUFLXRTdfnZLWfDSVoTOdrS94XjQLbvgx5U4z8f1wSD
7ipRZIz3l3HkwWNAuVjZNUOw23mVr7ZZL3YGUyWsPYz00h6fI4yP094CrREZsmR6J/eB3ghMxnAg
9PFx6T+ugUmdKHyMghGCgLUGWOToiFDCPXRgM61bRdvMs3eKupFjdMouxBBDl3SUcePnL9r9X2+C
j4oU3f6K6jO+DfRywVg4hqoOH2fKd9w9Jwm94u4VPM+1M0hTbcJG1UREJ7OWMCDYCY0r5u7c5+V4
hDqDChUXg85bd77m04s09DxJsY55gfVz42Wj0SoBulEhjodGREde4NjysAzbQO1MJCzho1KaXeQS
DNsCmAOgmZEnlVvd1URIfPzxTwkWrVCtan82daDcFOC1Dz8th5F2i+yN+7C4scMItas0npWL8KSD
RdU9dg9qAKD7oEx7XlPLMQjIV1GubpJYRqPa3AvEsKdpP+rTer/ZgsBCfgo30PMlHTm28iUJUliS
WP219zeYK+V0ouu7R23z5OIo9rFAdTzEUJddbK8izvonE+xjQhC5trVh6gvH6Me1MCR8/bn8EC9M
TXKrmMZoW8uP3R3lwu5CDE7LjftT0juv2pyvnu5WkP8HvheJhrHEEyEa7GtLai1kcPDglEgPnC0P
jGvPqQv10mqTMgTtJUKP5/hBUIBWLR+7qwHlQavIZBc0dl8Xcmbe47Ig0+v7nuPXmKiQmkMXquTl
PZb9OmSfIaeu3XKuY01Hna4VXb1BCgRgPeIfOHzypw5R3Pcp3E1DwfNcGMAz2qrSD03yrDDFvpyT
iUA0r//XSil37liXAQ9CN/txst6km8b6tLZJwM6AVR8EjRc5RFhnP7hidyGd828OVP1blRcxevVs
rJ2hjTzKTk8MLcGYSAJmkcLyqsBBnYy4JZOOqq628I2CXr+mnKHmaHUtWze4QIQij7UW6u5hFDfz
yvkAQ8g0p/v2Kn/rPHL95eR7HgCke8SnrYaFkfBXAamWw2NsXjJCQ8Sq+1gVyX0Kdpn6/IIfzeVg
wy6ZZTrVdQKh7Dj5u4qqvaTo/KOqipGCaiArSJ0NNq/LxaWPvE6yoXJ9ZmrXZpWO58KAW2M6m4xm
mQQwxYldNE263r8zGXVGsdwVUz1rimNv8HWLK7Q1dKl7ooGyp+3HPmZgkJu+3dSJSTetl8R8J8gV
ElNpdDrm95sy2uoCW0sAhZOkieh+jsJL6Q+C/ao6ZA/lE6voL84IYrWDBDfaSgj6Ru5cMrSyMcUX
eaF1RTQQZmKjFJeuede+dfhco5iRIMxHwe1LBgf4c25hMIYBAwDnE8uY6mWCOpQvT+sepxAKwexI
TM0iCWJA+xNacmprq0qK7modHsVjc2SzZ6M9fBvkWmPDoM9Ft2gepB4HK8okfi7kQjC3kEdENaeB
wwRqpCe7/JA46v0v1KJMqWcJihVWTE85K1oVX9Nc/RYE3plXUp/5CZOyAzuoOYmv0F/6i2vuzCyg
2FN95NSuRRIuvcwKMHtyLDeykp6XJc5rjTNA8GH74nXeiofO3nIWUjnSOPDBbZmonQTuiNY1/8ka
peWKfr4alWbQTsyEzNWCUcqh2H4O54YIYSRozhsYRED2zg3sWCOR4nw9EKH6xzL7nxlQXTHCVMcS
sV8Mciydjw+Zsp0aGvXXiAeU8RndXvucxt23x/unpUWQVHWrUMz0MlGzh5ZsCmSDpo/tt2wPt0Kf
HguzJPJpvsOoUukuIsrTj8J8Yz8JytFD2Xhb9NXlwRPh01Wp4uIsjg+1XaOBRAbcFez5ioEI7+ap
xdBW68Nxo3s+uRNbFpJQBSw3OMaN5MM8b/UWU8/moHmwyw39yl+fz7/HSr4H9+YC3H7w/DVpvrqK
juAOsn9/pFpqYr6uMf1YBHU8jploFXXYnjx1BpkXpHNz8OR8GhIvu1648hWjYkCQpNj8oJ7C2e0i
VVBFkR78i1EdohiOlSYMENgPcfZOAhEYhlLQi1/wBkLk02YhAB7Mi8lDwSmbuJwluMNTNBdz8bYr
Ts77PxkpGxnYAU6bJcRxKpIX3bj7S3rmsQ/asDe39lhyzCPapWMFhgmwOFRWLc1d60q906suTzai
KpKysLlBagJy6N25rNnxXU662Kdhy84wEaJWmgOd4+rPfftMx/YZAy6DRvAl3aSEeRzg0qfCIhOc
87HMQMd2ZH6RxbOb684dmM743dWVgszVxUNKiCx+D5lO66o9vaT1SZ9g2fgOAhe1xgXdufIE7jLW
FyMArONDf6DkHlfy8yBSMg1iRPw6WMRNNXLs8TRbMUNc7Tyx8NliZ+7/1oRqqqbQKk4Q6v6BMQ35
T/mMON51/TyvTBV55SxixIG+vAMV2kEtS/ACNwTkRNp8/K1BdmUU4Y4+R7aWbWAa9xyAalPlCM56
vZ8XwzuCumI3r+UsqZ6o1kpqt1LOBHSj96q94HaK2nSY/RsqnfQOzzOrQzGiYeK8882fQo50Qvqw
cJM1uL2jvzO7TpKeFRdatxj+XPRIfrq5l9rBAdZZ62xJ11P22iknFGBQ4nS4xnEOg13yXoLEiEda
1/jYXfeomYPmwnzSkg9lZANjByJqnvZbbiVZstADueFPV2t0kT0rmnghwgvhUkz6Ni/dcYdFmdGE
yVEDaYH0kH0KnP8KaHI5ao7tuqqNK2zUQEFxOysFTBQr2qSWnb5xKzs9EWmUnLQtoAhUyhtyZX/X
LSVvATOire7I/UF4DVgIhlKdQPA+Vyll2OOFY2mKfiGCNTL0b1qfS3CDmxty9dacZhz9/jzA39HT
ccEXb/DLL8d9mLZqlRfyOnEHgD+PKCH+m7FzXMTRincPHM32JvFyKoer63IFTq5IWrSABai51JfC
XnCsNUHUlMXrr6Dt6iZiwcSdEOdm1HfSwMrCaxKBL4dTv9+iltlzqvMQfSyvNZpj9Qc7Y/9XaMPr
E18ueht0jy/KGViILl/TeUtEc4ov5ESWLzk5jwhaqmDGHo3G8qnUpZ6QPNlz09KXaS1APiRhXU60
UXSOQ4yGlUuJtHTWexEpUDeKzBsPbGeykQjsKlvOSY9JXZ4dWim/yFTw/IFZAOOWAYmg8xbS2mpr
UeMvzNFy8rRXl7qSdML9EigHDkvLMMwVxw7jDyhMqStcDbenwTld0Jigl4UZL4jcfKzj+ybZ++17
zHhPDYr7Ia8EX7xpwfaQQCp3wgq0pyCzD2NVKBgbWINYpirMbRRFNjgaJxyt8jCJLcF+TMADGfJe
w7dryNRlrkp9TuQgcnCOCwZWluvhBPtUnzUGEzWAWcNcWQUxUxGlqjH1C+kHI9Vj5JrcgSosPBeu
u4e/ep5WONiEzD4+n8zuf4UUTmyn5yUPD+qk5QXDx9eYcTaI1XbjpeFP2Ap9ijkvtQHb+poOWPbB
ABdmoU5TuquFyXFz39q/jhsUfFHPfjn0j9jaA+s0Qmmqzq7tV1g0i7oobAfvOuigUeSTmXaFT6TF
cefmlE6HIbxqPycSX/903MJQ0nK0bcNEkY4UGhV6o7dZC3LMz6cVM0q35uVkm5IiADYxN0P+W2ls
8mgbP4afERlOMSFZPFjtql3yPbdEcFPiIA6KHSShKf40Cd293Lhl0QnVciirXLA3KUdiXG8o0w0Z
G1IL/uHzKcJp1ugg/ecNCWeTdEGyb4QCKSAJ7x3nt2RYnGioSSh2UHycWdFL3AU0/MDJ1vkyvOxa
YuKD3lSjOfnv9Q9aEHgGRKofGkxEOVw/sYk8lSSU/hMP4HFQtfdNXGjo/eisVXmnDUny1sg04Yph
8HJqKTL68sQhSuPKNjNEXC7xjGPrWpHfSWEJvZyhHJyKG+LGHhrOR+KcjzKnfA9PiR+ZeHdH9haw
Nt5yu9C/s3+Eytd6THEWWfxm5y/fpN78/MuVVa39kzuAoRA3SflomWu9GUXp+Fmd3uIYjrt+Whkv
+0C/+fYN0inOUSPBQhmTNhmhQOJM38hfW5FGeq9LkKPwPMWrcE4HKTctKxB5HZFUuOLVA4OEZdwK
UVXRoFdseNOzUGKW7xUQp42zUcR+fFuu9jS8ReB45NSz4XhOcyEry7FiURK37N5q/Ucz9Bmr3x7c
t3ZYJiBPs8a93Y3vNB0c0v5HXsXjmpITqcY9+Hor0NAU4VDudoHlRuSalQyG0eaMOTGwi+ZT6v2o
DSr9gVsyIwIBR0FnctTcM25uklWQkHQqek7zKjRgKnCjot6ivOMuGOGvp7To+ERGKNkJ2zWPX3Gw
eXbmolG6QiLnfNS+djuUT9VXf2GHFlVbuvoIxck2C8ZBuX4ddh1ao007cm0EnftWvvTRnqUMFWqr
GWtQaDXo5S/m3sevVxIXszJ3LSyoYwzEQyF3x1AXLtCluifJbRBtK3kNKrH9c/ty64gteU9yGvRA
5Y/M8GyXjTNzMKY4/xJovL39ci5Bts3NtMwlWAh3F37GOiCSUPVM3yKRorRlzyGto+zjVVy+snjJ
tFl4zirUdydMUxuwHPuU3Q5S0AjhrlM3LSL2dpkHenEicXBB5bAHz/kgvDM1H5azPmpE/LP2GQw3
vA6q1xVnqwe2MZZuu84p4THLeRwO9T5JuaFLlAVwcSIaCJWB4vIoxovxLTBMv9Kjr784niHm0A2A
ir0pi/yu2R8t/mtM5BBjQgBPVmPtDc8MP3yiCpHuUACYZcdVtmxoBknve6ihabkmKUKqGh/XtPFv
bmiaPXip/KrpULyijhyshfqqYuZcWkq701CYAPGHCFnwOfqneyFeiS1hwjyfd7gHxRgcQeTrITwA
kiOuC9qbXgNWVfYCS6FPcTEIqRuLJEBcCSRlifwkXVhqP+tc+yCtG1A6766Z6B8lZeN+a6Om9ZkS
L8IFrm8HNvrv5dFgbxAG2POasO7kEz0EiuGTXFmjew6ZLC/zXmXA6vAcNdTtBOFSCthaWUWhxxgy
zcKmHgWHFGNU6APNZySiQmEQyxLQY+bzhVSVIIYPlBvhmWCT0JZ++KZ2MVgEmuId/Wzmt17GMvkV
1hvgkXiulrsiWhd+nBpTbsDGR+jxKMjXVRId3dk2GwTQCuzaxBySuEmWCrfGl7juAUgrFvVF3A9h
/5EQW/g4aFBGjnZtCcnfQ7Q+FrrjhSvG9wsES6t0Ha68lKQBR3Umghrb3Eyczj27fxC8Ugg95QfQ
xypjxDbi+c5rJKKYnUzo+4jlDmqJTR/18LzAVf6R+MKgKLkTET4RJfR5ACcLgZFaEUYALEMAaNBl
IJ7CFaHQ8R9SFfsQdzrGsT+MxWPjzJNBVGrNkJLPa7VAZ8dX4oXWrSyw+tWwgaZm4qQga/YyvEub
yFD4deQcb2sznstsmR2R7HIqX/6OFEpv/HEU108abDWa/BLxDd30opkPOhfdkR8FlznZ+XDCDoxW
0sWINwzM8Jl43/FS9RTmzGtoyCmM3A0IpFz+Ywod1EV2W2rq2HhOQJPVw5b+M7clEQlXcVA4K6FE
rNMt94cK7MNE76HRJ1MkmKfzf6hN3ciFQ2X/EDH8A3onFt2GD5Jr2lIbcaMbDu02oVjofp1t7NEd
b3XVTEdme3wZzEPxS5bMF8r7BLnyD6+aD77wbfaOVywmOm8vtjhg18Pc3/ehOH9IO7BicOcDhHPr
2eNf9Icbz2gWpSqNp9TQiZ0ci21K5s0Joi72/Tw9kio5fYirolBlZlNYWfb7cCo6xw8h7ZLg17LE
eukmevL3G/kJoYFQGAi6AwgtTMfoS2fb0hoiiz2AJlOuPvyhsOOIMn6Zrble9R+RPDvd834n0sC2
o5ozfAYTAKEx5wWV9lJz5uImDTLBdLKjqMXz0jA8uuJxDad9pwErPA1YHWQpRn4Tbv0kfB4wveLE
noMoDWIrkL8hhTVuaM2hKcJi7QkLNxRs0bnqljxRTzUQvErXcyZn94UL+P4K8XBpZZqAdKEnuSzw
HGX6/sjab/6dCvAPvIsqW1Hj0Jic/BGH+ntyt9U3Ch+Bv6MTd24DT5EL1QgTnxPG+3t2fisx7LKB
I8Lr5c6kMbHCGV3dHn6bjR5Z2mdNluEu9CQ57XxkCWRjSqkucj4pg9PIajkV7eem1JYHTJFJbXu3
xisIo4U8uBq1CBd/H8uU9u8hOyvRxvHmTWsN7SS+/5lQFLc+oPTtEn+ibpqooTAjRapD9t+OZMPA
raA3nXV67A9V+DsKWpcC/+rknBlNI8Z1sfIcDuy2Dmzv/lKU7RHW6nQj1xafSaPia8s9bkgbwKuC
qmMayidP4tGzuok0qfR4axf8egg0FEiBsrApKte2ip+6fkRqZ9aDA/hEzuKx4bBK2Yd9Ti642sW1
7hRl0uZLEwlpe0qJZch16NVUpXK7rb4x9LCOqrRGBv1Xjs0iHnCyFW5/YB/oFH0QmNEXHzIILuzF
Dxe72HRRExGKqqkHyHU2mEXw4zDhEWNBBmNd0trWMHOpgKMwN4CVAPYpFGfWJ4iln7MXmf7JEl+D
6mQtijiUBNUc4Bjj+MmKKKwZMIGW8LhWIjDiUTNDqOFNv0XyCsViZfYgkGvDLcpmALpBOuw0UFVV
WMz2aa6Cvde6/hrN0y8sYdbf0F+F1+FiUBdeVVAIpgcZThqQASGTVLyx8tyRNHYy4tvm0CF5oHpk
aUgRSq7RT3bhQDythfRBip8IkkTyQZF27mI1jxk0lCxOISz+bcB0OE29Ez8EyXm+AGoEt8Aip8qA
qHXkcRJB4ALLUYGEfswOxhXSk4Ycap9N6ZZM1AW9I09fADliyiFQchzyejJIjmCo/KU8yb3iBCSJ
CTEeiuqc2NxuoJZBA+YxHKXih+0KsKVGatOuMI+JcpNaP9D0w50EkMEV0eHV7bbYilxgxnQC8ZdB
k9pJMGEf8z/JXsBRx2Zt85YuDB0fd7FzdUKrXzRghQJiIST9ed5VQUehuxdWYZUfH6yo6KiM1J8I
hy8CQdP0L9F0g+Ak+Id6+2KFNykiuNK1h3ZA3Drmro7v1DkkoC9gKPgpCQfBa7xtYVgqL6aCZ6QH
tu7wVmg0Fnticdiu2zKPZu0ZvDQkBhR2qAuzDJxUa5ySe+OpWS2WvrME1OiG6tEfXwpd+Bmq5hOz
a8yYfXDl47De3TA2cKEwqOfMnpGCKDhhEKOf0h8bFn4JG2jpEXpPMlzvR5/nuwgC3J1t/Yinvn0f
8rO6wrIGyc4LAN68ujNuXUayYjqrxiHxIJHI4Pi+t64IKQcmlW0Y+twXjWSQVqieWxPLgY8yW7ZO
k/q+Fg+he/HR2rMggERsFftgSBpc7eOSDWCi7rjP91ZI3W7WNr3oxph6EFT7EcKoFnU/gNXFMmE9
LULCNywNpxOB87rO+GrSBVBkvJsuWM197srOD8fsEKPDh0PTo9Y6w9kUWae6MEVfYZT6KfQS5cnN
gyRxXBQ/6oPCBjzxRQQJOAL3y2rYwaReB7cLY5F1P5tYzd/PemWUMEjtb/kk3xRMojHWmCjanTVH
ManxmfDeMFr3XfwlGoqMwZ2w/vAC5H8dZsD0nsKNhVcjn0Bnv1l8RZ5/OkfTM5zkwzGcia0xLHJ+
tFnREUOE7FqIM7gfML3WuPsN9nhRCJaCSCHkSeDvoxyLWVQHaf6LzPCl7k2RWX5KxEMUHX6cnQ2A
KG4hmuLDFH2pjKgPw4fizISvhJEY4qqilyTW8QtgD4E1hZK3QzaRhfJ0R9kC7iqdSkShSuKXz644
Uxb7FE9vpqJissd45KqvxMDGx8A7vXsbvP4MjabD+TRNDEao44SZvjHPMSh1EGY7opg6LWzvHUyd
82MzQOaJ8bHVYO22NxZSbsRWLhyK6DBl8Y+qqw+kyQSmgbvEHngWMnWCnu+DY9HE0elGqm+qWUep
ICUDcZVocNMe2KA7yZRlbcDrXzkiJwhoSeB4aJmCeJwcJ9Ojjn9m8QYRz+lEv3WiOTP2yViJd17+
7EMu9BktEJvmvBNUDVrVoAGnbzmXWSAB8c03G+EgDVgktyMw2Lm762EQs5L87Ww2qre/ICBk8QVQ
8luWM6+xX5ZAVvfTE1jFCesaIGi2KsXzQlgqcgNNGGW7PLAcxRmhbVMYe/1EKg3cxK7fJny3bE2z
7BjL/+UUQEOUbNStlSJRE1QOUz5wcqIy+xOfC8GRL/ZsR8zNQDD8i+SHTwAxIWwvzVW8sTVaKQ6h
chgKOn9BHXX1g1G17qdblOSZX8r5C/eOuSGQdmTVUe8l9L5xTmJ/D8V9DoMZrN36NFsXYR7+OnvU
NhR7E4mnbbNjkO2BFMjuxdok3dW3hGQ9ekSkmylRq2YyD5Y17pD2NGTKkGi0CLaFAC1rY7KCqKv5
9oItCsTFmfbWelpDWczmx8/F5edM/GLbDhk+AXRU4iQ1vYQA2XSocxHorY//SClWPvKYkT7OPDwX
MLMQ+ksje5qPPLppwYMfbZcgT5buFMMCrsiYkmrn7nnNW8/z2HBA9YufFS4/mUrgq1jpUVx7n5qG
u6iMx9E+cumruZaP9eau15xzDjKFKewgifrYN6LdVUVE1+8YSA9slWE/ynoBU9JEdw9oYrfOBcZj
sdZSlD0MtnzIlEI2POvAvVai9fDlvyfz6EIBm2q/f2tg3GVRet39CITJj98izzLKt4nqPgo+6NRe
ZC6hi2LMJvj6Qk57AUvSa1AL4xSAN4o5nxiXbIM65hhIPGzFwrvjsgMP//ZbX0C4oFlNNpwo9hhJ
jD00e5e1ofcKl+y21teaBGhl+ajY5xGwG6KNDEgRbVaWX/+bCUiIY7ZeJ9xzsCpg9MaQRn/1x9nA
RnetU2JrImQo97G0uWzJzypGvIJtbDbNyokymMJ/vkFfNSujK8MfIhvoWRPoiVREvIPllkI4sWcj
qsAAWUpkFgal/Ys6823BadACSzHcRO0RJuqXO2IFAsAM29BYHleotTa/rUF9n8qLsfWhvxTb9yVa
r6RMx2MR73q5MX9+YnOxDp1nN0K0aQWs+xTwcNYmAZl+K643rbhuDwblRxcFbjlTvj1NkT7ct3qL
pvK2S9SPyC00lFYjK37MoUl7U6ekiAtTufKEvumdeXqJBeRsHHzgKKtt37JQlGiOLWlNxssPwbkv
RKDhEwyMTd/4Tjgyy0aPsUe0MC5XxmqftQjn7mEzU2Xy2JOtuPGt3/zJBUmE2cCayw39sF6fKuZi
LcX6CF/U7v9s8XtJWi6G0ElI5enn3I36cpExWNU+9pwW53j4zK+Ikh821SJI7WZtqR7R9YRaOdhl
yHvN9TnHy5KG74tv4L8CkefYC2gsBOtJdZ2VR/TrPnN/kK6ZDT/mp4zaT7keLbjvzqJ1XqEOTY7Y
VbJ/fTPJheqepJdmSI8iJgoBUuIowCa77Fugmn6PS6XsjrohYiCDNbjCXipR+BnTGnkw/vGhzd6h
xSv02H49sYHDQ5K03v5O3zbl9B18daSwcSLDd+svrxhHhjsa8fOWjVKnLDchciject8ck4T16OQ4
4pE8MPakc9x7+C55jNnummB6SUBE5iYC93C1G1CGR+jS/kjqTXb6iT4PE2xu6RRYHSyKEAQvplPj
gh00lT4yLC5j85Jsf9zIFVUc0PEGHJ6rQu4XflRewZpdyARJ6StsmmqM20143zTX3fUmz8ec8DrZ
Fw+WiPvNhMh9Pw//LjFUxzp48IzwyF0P1x7Dne8JpnCbqITaVHS1v+9qDNHqFVBqbyylozmyhTN0
tM3eZbHAMp6xAEnD4xl162R03DdeKOgRl9pCi/2iFO51Ipg/hFFfuVmDoTZAg4bwCqPKxjANvTRv
0XxzRNbqz4dqg3WHumbTAi1766IvVHWgo0TF9OpuR18zDi1IP5E91FdhRSK7NY4fSRFm9RaVUeCO
dmb5WiGiClo9SqMBHXnw11ytQI2p83fxHXh/j8Zv/6tGVPjOsNAla2133yes9gu4thCB+N0SsZLr
UUPBWaU+eLdge56MMtRHDhdFb9obJvCQZRBb0a70rDc9DVFHIfjxJd/4CZ6S9LZMWPKb5OU5mqfk
+vaV8BtZL4YBeVQwDvdOvKGnXMjV6iyrdnKWOK4wb8Dgrm/bIwV1/t0t4+mIBB+IUm+LjyASlHsL
9OyUelV7zw4PmDIfYeBL1FyASKm9oJ2BC5CwBTmkcMXW3xH4oXQ7QTMWK5KVG0VpjRjDldR/2VOh
TXCb/Ug9l6jhRC6+uStTwPihBIVi06cKkVUiUsdYDmFL44JtCY0qKF1uAAD53kwKxCuuiRa5ch5E
lL8zOIuaxupE3dOc2zKmlNzKDaXXnLohz6H/yZrCi0zSN5QoWoxawfYBIlY7e98aJE4pXDr0Z5LJ
XAUgLLG8e4af+Ch0wQ/bOVgh0/Zuux4WfbRkXb732xgUGoryy6loxx470Fu1wPD6obMJaxxRUlr7
rBmhbk0QUX6LeCf7K+o2fWv8GfKCkf4ce7P6gAczM48AjdHXa7cxrCjNaYzuMxy39ojOuB8fmW7F
w3FRyCwE1OzyxqM63k/YDwFUWKeySGXwmef9hCYk1qjI+SVMFKaa3fXB+yEKD+QtBoSqs5nRaePB
vCin31BVumyqfbq+fI48VY3KVnGhv9zK+RyrZ4LZvGiOCmWHc85OG/Ar+B9JmoEnWEvfGoSRgUjI
vE2A4WNjaPlJnlu8U/yIYz8bNg4ZLP1Djn8cvtB8ciSU0QPNG85tFvTq3N8TCg1TX/Vh7/omqbFQ
IDFxp5Wis+SBK1X5EvPOusCYSSLB8MWX7fvYpqA4Qwy9H5o8Ai2+Oc16yIeK2X9gJeDzBnQxGhGY
aWyLu1mDcVb14VTZn1jBRywBogVGkF2KZmEkTEvjlh6saRe3INjvfGNsoeWE+nt/Z/q9SJxMdESQ
wvQ0CKoYTYqFdklsc2pL+0V5GdO6M2y/RyIMBiiFMayJgwfhZdP4gxBnc00zITFedViAVxKEG72a
eKA5YusuC4luHLo3iNRCL/IpyP/ovJxt4ogml7smb/z82pXIFaeNPXO+h3kTgC93zGIU5HGyZKHf
oNh1cxtnZvsJDJKTu4OSh7vMoBv/8e5A/cW3M1ci+jebSBtK88BYfC2YvgK6XByZNqXx1sZrlhcP
b1gG9ybDnRPTpmQOJAMrCS8OFtecJ63xFAb1lrgy+iXYOI4DtZC4gpn4Ibkw5jnYZUZpLYqLIGRS
Ex33LesHVqvOq3/K0b8yqZgpNOm9xZKmo43QxqGrgXnz7yinWdrGVb9vDRwTXjZlSU8x1NtNQN78
OqfgcvieisVfnRHdKTt9lkb0VVlLjTmDssd/nFaBxmLXw+omTxSU+o4xFOf4+atOMkZtjM28o6Xy
RV+AjuObC4XfDXUOdNUMhRE+Pt7wZLGgpK0mewkFLGtl122fWOADYBs+Ke5FMmjh6BCLKl2dQAfW
Ux2AyvvNEbs3fMaDAQhhRVWbQg3HcCVOe9ZKOVfkLD3q7V0sFvWO1l17SE5RPBQYAfT8DsMBlUx/
Y2fT0/2uZcHWPlHYuvdOVFNtpbjLCV+nCEJrxdGS4qLOoO4qBwSYXEgJtlVs5sAzHB4R4T9GEpeL
hNms/+awHMxe1HwCXCDuXKkenyc7F0SxczP/yFSRrbMmOav/VCbNOHBwRwBWhegJdj3QGfyhCYc3
5L+2wP9uUnqYBgil8xfeLAEEMUs7XeXNhGeoNvtZ9IknqR+hL9Xt3p6/iG4KHjzBUsFavY6d098z
RAgrT2WKNEjWGvcVZbEZONaxCsP6E3JaIWPn6iQGKt9hcWrsFdq+9HVfyWxkxL47qe0yXN3ftvy/
2eFeX9r7j9b43i3/9OJ/hZJYPW/EZ1yteqcKAiXP0anqHDFJ7/m7ttrqgHI/sE3E6g+elQ5yB8e5
YrmEL26y3U9pU7loHAo64cNh3+AKIyPUXqcw96f70bzGPZuJF+FjK/K6rCnyVcUfaLDyqTiuajCF
tyoiplMiDuoJiuYTLXlLsY7OPNqM0I4+5x5As8L/PZG/Om816Cu3arQYLZSZCGYdmXDGTu15+ARJ
tvtr6ifioTsOYQpFSUUMzepcsWT0XPxPSzTsFERSyaf9t01xnoN5Sn0Ym3Fkbf47BSuIsgebFKbV
2QpXPnTlxI3tLY66Mmc9py0lTFc6VinrtVcT6QGUPsQZCMSk2U119VLEtu9924HkfSAg9RoEpPey
8gpoTwCOMF+pjPyNY3AXXjQQHIGcPuinYw6xVnZGuunkHNLA3n2tMOR6DYXeuuD6dHm3FGk1jWc7
1OEgQjJF/xU4JJMZGJZa5KYUsB9kmqNCW7jm9P1wkyXmO2rZiTlZE6jdLTMhPKjgx5ZxKkdS8Lsr
TMp6mT0C4HqXVl0cpHPr0p95fsqwh1z/AnBr8nSRyNm5XOEOntp44E3ScIHbXuvo2vLarNPQC2gP
h1WNwzsqNNuUPspjB0IUoaYLBjxXQUIbhIQ6ZTWb7sW4PbRkuVK0r913DYsfauOgDJjJ/O8rFo4c
qDmnf8LrtQRWicp7CoL6rgdesa8uFOnVKupSU8EVcw98sGwJ2MlXKBoNwRyfK+igdampvbwlPGsM
4hIyvQIpFHCoFf7ay2EaBIupjSB+0eufT4YCOcsZe4V7pUaXkG2Z4YC5PSXHRCnudJyHLQrt2kHk
Pu5mStPjr86aCSsTlWpXJgRv/7iyqwQMjjJO7sEox7OlbxhW/PQpvP0ifdNGVABFhYRQwcj1ow/m
zmtkPtUaC9nr0xMFhrn1lvWkSgfAeEwe4h3pZeBzqIbOXxOMeb60PrK73n8sjUiT5ecUaXc8XF5p
wNJlAJ8wxmTldtaoIR4eFHSjEWmlHkZDcgBQFmPf/D4J8oNB8gOggHpXbZ12AaODeIDvSeWx8d4E
r0JxPWOTBSj+vsbrVAsG9lKBd4CvNGWI3HBeTwMKUc9ReVLlLoYOEyV6uflS7HOYzcIR6EbPujmM
4MbOdupcASxna3IHHAIN+Fdb7HnWBBtNLS/+li777jXoaq+xXngMWicpHUt7GM5ydI+jGUs3PbWR
+dWZ90fGNMppF/uzmWnxGtUy6TSOKT2i2WL1vueF2PvBDwsDEbjjHF65usXC1Tkq0vcCMIXSGluP
SHauIIilImO9cpsLBc32mOd13PkEBZRG92cR0NysTmWifxOggxIlMBEdJtllGA4gLZn9aisE6fu5
Xk5jxYLU8+ID3DkfYSdqpg4c2TldHtEiLhs8laQR26IIE31GiYcaLzD/s/8eXnqvHS2XtZ73oIsi
D3IfEzgxcJAHfCpnnwrQboTAoTV3F6VUE03R+vHHC0NAoHlpoqMhoFSZu84C0RnuZDfdPy2An1PD
IjRZnV5AplJZ0OKVfp1Oi91yqHRA4+WuoHGDtnQi8lmZLW2h4IslVTdRGMQx/bp+t4Sippljc4lJ
nSclrg2aMXcvQ5v7hP8CdFEANQ5hUXr2HCFvdLwkPrd6O4VOdIrKUd8OQwuR14LOwd3Tnu7m1BtS
225JDyXUvuX9Z225vkPfdkascd+fBO71Hrq1xR1X4DTEbzWjZ5e21/nI2LbrN8QLXSQX3xPBF9TF
i9ScHs9JCtIbuW9GbCBn6nPiFb9tMhSwfWLeHtThrh/uvVzwQWTvBYzv7LvBPnkaH6JMVhcWdgyS
oFboKl2XOYtp6k8XBmHFcYQIwiq28S6zerQ4a3XThB6YRR7NUWZoAJ78aNYm/2q3dOPM0g/y9DQt
SSMNe4L0qncdoaPX3xSJQa/YY6FpdcqzUY6SvmmXFnc5+Dm62M7VCW1r/o69LMc7aJcNLuaotRb3
EwuOev6pSvuA8eNcNpJowwo6GJkeMX4jflmo2Y50Z3U4nQHtudZMc6HJuBKDH1oGcKIdU8wZFRxI
TmsV/85LF8a/mNFZEbzTmffJsN/GQIBvjmUkbX4LdUuK0NTbRDjx6zkiOmkSTvZSNhYxvNKqK9Y/
m7t9KUMp9UYIApQZtK1MenD/q6U54gKrkx4q/46ZONSQuE2VzYdEBxo611zGHPIZRWrABHmYqWgQ
4IACMs3wvFUI4PW9dZ9L26ueTUfUlWNjgVD8IaUM8SQE3DMUv6kMR78npmUGggVDPz6mtf4g1EB8
CV5HLem4ra/7idrfbDN0jxjP+5JeHgyRItm484xdLTu37LULrdGg6wvT16zZCpe8nAg67Yr+aBUy
1eFrUb8Y5JYJgJM9rXMTO8jYJfm0Mv+zD6G3lO5Ub1h8qGNffDCr1O4V9Gn6oNC2IyJ4K6dqWPMp
qe48GTKKTtxjJsbh+zGoqUF7xJTfCAorT/HR9Y/1g0aGDmUbpcGlD9Y448XUhaCKTe9NSKsyHhIX
YXYUuV1/GARhihalh4KZARR3UHktAw52VJiCUd31yWjjMKZSFbNLpisvsBx4/Drre40zinubnxio
Jc6Pc71PakrysYn3Rms8S9nillskZHidWYNmYqk4nFj/Dw1J9L3uGE9CB8fT//BUHLwp22ncthT3
XFlJc+SOLX1unzP+2J5AElcFrD0vqL6DzKjq+FNBOWEEvWtx6rdSCky7iQqYJbH+9psEiblNSple
AgfWmrVulhIfofhqCTSUXAeRvC4b4AAOpqPe3KuC4VsbNi4+zy6mNVGgnkcIDPE/I5X4ot/TAkiO
OWp1T8bluIvPlLcL5oy+JYcfm42RIFoVULxlh62N+2lf+akwrHXY1qJNcRX5XuuVoL6TmuyY2T3Q
Bi+p1KxgmfvGRpdaPCkcBXBqkIAZJovGckFaArJAJRkUzujY+7OqDg23ZvjofaAU/a7PUyb5QQ0x
BdFbxTiUqJsRTia51Xxteqn/6SgLF71bQy5FYF+GJpJJunWpGhWEYoTXnYXgqDAE2avRLwnYkyJ6
Zkf2FuOpKmqM3fv7TLt7gvly/0pewGXFfb0xzg2JAXfg1ItQa+qtBMJ8FYyHqntJnCU4CrLORQEn
+hAfckEvRt0Ey0m6fczXPiZ7KJLqxZeDdlqN+d7nkyJxgEFHluvkSkBdKVncAA3Q5X2pOgxeQsyG
rihAfkqe8QHz96F89IBPn9ZnWrTn3g5tx5dzHBEhL7vYwkupT3unQFbqqqL7QWbKIPoUk6sSwX+b
2mxIdjC5GMDLYABeAtda75Hf2sDbrT8PpJfX0mYFIpOilVWcgyhSpFjsEwq4p2AAn16hTkh44fqm
UDEFCGK5s2vma3OEwks+nO+0F4nanTKDhkgJ2wSW5MJZ2SO67tGlVlYWYMvAn3wy9CZv8Ju7xm3+
hmqO/tzbHJTRW20p1MrubMXSEN7m20O+cYCtL6XYgdLbX8AAUxx79dUX8OpTJQh+YLvM09bKmp+P
8byobv51pENoWrZcJ0xVnBT1AJet1ggjjWyomqJRWseqzGcQyEwLeJzgxbJspHVE0BRrV1pvl/40
cdebLduqn7Ws+boyhI8+hZP9Rt2DFKMgaLj2UcASzWRkCOvZDQMpO2BFobigy7ErTE7NM1t94t0j
hyeesL/k8O9wOiaNHmcrO3qEdsnYisq/Llxk0lqKt2+6YtZs5DwQNAMG6aN850efmaynBo121qTk
0fr1a3nJwxS1j84/3AtU5l6U+intgINDq5rvUG2gbNQG3s2JoKWQV6/4FejYh0JLjGJOC/envP44
6pZR0AoxWEJBg0PqfOpNugZQypol4/Wsloq0P2OxGIzA7Ui8idetrrNJ/qvhfZH5hxyTQFuFMA0Q
Mas5QgcyhT5B3GX9mNI4nFdVYTrNJ9VLLFpDk8rExr/r154ImYsTkR1yQUTUmiSsq9aGHp5ftSgj
xjEkilHpYw/1SoWzbHFl4PME/yuTgg998umq4Ljv/8CI8K7Cj8XH3jAy955Wm11P5CmQtjUPmH5b
VZUYGTYU1OZX3EBsufR5svVaeaI2IPsRZR0PsbV+DkSOTPgeZAi+kkyXTQitOwuClZakzhWHaoc0
fP29Q2c/nOtJ/DvVDr/6xfg8SqhWiJX3Gl4InE4n3ZnFGEPDj04qZkQefS/OmTyLmvIxSQgEI1q1
6BH7pMALWyEJ9SeIYyO4E1YdPb6s1/UQM+2HiTi6pkLzs5NPm/H1/MYWSM+wIR3Nn+dnDpHqZdxv
XST0Hu68kMyT4p3bQKtufndkWmpRqQI/flcbts3cCpFcbpRDGUyBzJyhXdrUf9AoBxCZaWU4/Hw3
Qq2aWqaSV23TA97MGqLRPFwl9tMslogC/LCpRcUuaFjoCjmKv0F/AlTZUphbMf+C3mvesKrC1VPh
O1UfS8cBZwVAD39unch/ec8TDOS6P+BWJ11iSqk99/QOg16+OOPvNo/kDSAbqzfkOwSCvg1NihjL
w/BorVQ8MHkeqXCS5DQYRsOADKYroQA880tPfkeMKaDwjeclpanmRj0U9Xkr32sKH736/r5rs3Qd
iTpKTHFXBw+Av/8mvqyZG8L722GeTjQPK8x3G+TMaAiS0pY3dLn/F+dIunUqfcHbLjHzhMIpjjOE
LQa+4uI9/tLvGh7tn8leVDkARSvE5NpUya5KwfcS20i8PBBQ/FG/WR01JGEm74E/Fr+NyuydY1E9
JyYLTKmwZyJWh47wrKiDeC4d7qfv7zoOTtsthjepxgP7gxLPhF14IOKyUUrqKubyAwr22+mCeeoo
qqIMV/74HewIAiG/gTwAwIbd3wilGSJnoeaaQr1h39Qub64bqZybT6BYPEVn41FseOsbZgQzwsLH
C7me2A3R/dxVoUcJLj/2J2llkw97ETOERtGnLuLgPfqJUufwCm+f2TiabIe9GksFhPjetHJ42yKH
oZkWwTy+VAjLj/e9JWdZA3Lk6xKHjSPeCIXn8D9vfzkN5rz/I8kUUMQnyCy/o6+uS5YZRgRy4W4C
KB5AFH1YbOpkj+/lrZ0HnXj9M2s9DCCIMm6c6EAZhZcspdJbIZsHyQYfu0lSNJ6FcwlthS70YFOB
ewLOdpZeC11+usgI8XLDdKT5zsWnlV7zKTusi4kcDevkarK0XX6M/ClFG6PYtdjLL8RZIbwrmRRi
lKiw1R3pOjgDcXT6FVpj0X0z5BHTYRNhLIgs59JIiAzE+tnTTTVcM3ltjfBMLdH6vKRtPCTrEyOg
GyIq/FfbfgC6Jo7YH7Yv4QVrIh9JGCp9+2wjBsEA8KfhgxxhksOFh6daOOQUXrlv7ufpff2oTfiQ
FnjQiJrk8rU8KnfBahKzPdrp4Wo1fntjQHdZyYkM8gnrYvDDU1oUtITFhufm6OdhsygFCyAf9S9u
UOvYTBbMtn3cglU0du0I4KTkOI/ZCzjpaOBb9SexgfyNDzA+6W2aWzH787HGG1KT3mXsynHc/3jP
e7FtQJhOkfxwiCBqxVSwwHFn99Jy3HxoYHXmGMUxvB/b8U3owA6iikif3LdwWOKEhDpMztev6ewf
GH+N37q28QsbDPXhV0Z2SxHUnGP6zWbFY3BsXB7Gi4RqNjBYcxSCXzoIdzWC/umtH3n1ebOT50zZ
Ze4o0jvJmiI7og4pHLq8IYBq/s7/9YF58fpnD/sLPXfPHVzo7V7l9WP0k24uDrAdpm0H7cL8++ok
yiLMb4u2zY1kj8510blKWumWKX/hrn9AJhhSq349MG1GH+9rWiGzzSiGpSjDPGbtlfmMbMMDw/A7
zHz/F0JJRc0lG1tslPeJf89MGnh9ue2FHEvTYCtg+yVnrmjxpiq34Zmjp0eeOxZ+DAC9XWVypmIN
qK2oa+iyzEVnvUi0xKe8Pfyki8mK0X8YccPzkTqZ45FOi9zCzfJ9NNSrD+ed48UmA1Iqia8JTkz+
4M2nQOePucOOaAUrkgoVzTEBeaDUij1aGa6DH6I2VvTugQodm8MiE5xwDOFWzPfthkBBk3N/xJly
BGqfPQsbF09ZWNKg9q7LrcCOVamwhubNkyOc600JR6iIjLPtrZbD5QdE1pwonfZ8nXZBC8rsIVFM
T6eLNuWISOFdZxKD8zmUcbrtPKdmhnx2M7xOUQ59QJO3tT0u8rrgouhQepfSjBLxkOreAfKud9Ud
1Rt1NmQhqZF3pV0hET6tOW4cXSg5RMFPuzfozQaNa+gICefd8WKrG/1wkIL5v0nyLW/EdgVpbeVt
1NMlKUSwGu9DV+5q4Ps+bVR6RWuZQBSdaMNEtNBpewunjbAURwmB3o3FkaQl7b4qVCrv9Sbo1i2u
lXIQLWTZatYGpZRI88yVLyb5oAyLYSVxECY05Hv2cTMeX7Mm8FQUDohLyO4czCtUw/p3OxSfX9y4
KG+TlBkYpSNFjGTHtD4b50ZCNQ8cHpW5Xh4Vq8YIOaBBqepwqdPTfsrnhifk19OqqxJOaDr59ToR
X55ejYohumcpeO5/TQZEGkmQ0EQdxPOAtnNAb4FWm9FGKPgeUYR9TlYsS3sAqSw9i4bsQxuVVzsC
BbUXJ8fZ+FjIEgV9Ds14XANepJ1jeTEZ/Rq9iLKC1UEb4/o0KzePzTYunwwfAiwPOi3SWGrwoErw
Ylm9alDMnEjANAlZtCC5eS8JtyUp0ENqXvIohveiY7Nx/tXcJaCK/BxCMfIuXSI76oV28mSTSx5g
BF7jolFChmTcXE+MRI1kFOWl315o1fSHxK+Li24ZYHD/D9NSJN9AoBWzPDNzavIbZYHpNjTi0reK
rqbNRYb9uHqn5KrMsXCtjIfGi8KfWGVi4AP5Ua2klprzf/76jyyb71QgddiUVEjAcTgOkXU2UFpZ
hoIdWv2c88I+J6SKuhPfPQUg4nN7K8pLMmPExcihA2bWpYL25waBGyQzPE8TPG+zPuC33lBn41DC
yhXXvJbcQefvNyXHKuvnCcXsX1zUm/ldvFxV3q2/1ZrVRaJ7L/ocCsOMBFvWTbaGVW8IMtdi6d2X
L3yBG+ZF+hlnpOhJUP95QBmxZN8p3Kruoh+nIa71jHfUj3I3NSc6vS9xqccRuSr9+LOxYrkx0Wi/
WOFaRp7ZmvTzCmKdu5oBHyX2UHrZpQNonQR47iMsCmeJujRpUFA/yMkM/Y/D7WY50wifoU8QTm3Y
lTJABhG1Hhc24bFonZjtlqN2Jj0q/MrKjd+NrDFeQXYDaYVhiX8DskIY5/odWgcPoVT7sENNizBA
s3wdvuNakyogcoDu9ZK6pTUdnwaaDMmWIhNE5yU3ecsCr6cx576C1/406Nqq9/h9YPvBdu5LqFAU
G670lCDtAFgcqJx4zSLARLgKZBf/GTtUuZHzaoyQHuvfuqY7oxkVa7SSIa9PdnFma20Sscg+SW0+
oF1U1zAk3cHJzKyjs7WoHDEMuRfbyQd66f1xyzvd8Dg3McJH5y5/l3MNMOUUGXMh/exUgTAW5Ld5
Uty+c6kSp1HhFl4Efi4QVechY+4E6UHLoj14i+YWJ9y5CqueLfrVhoS5ypCPQrXdqBMCZlf9H8C9
jn9Ns65dd//ANSauMXVNBkB5PTbYRW6QIbkhXk+5OG74HECMHol2Px8QPkhZqPQ0VAFoSN4Bi0x0
U1c5ajWruffdObllxGHUPe5Phs2v3AQzU1FcBcq782JhheJ9uGls2oIu+rmbRUF9jUZlFnVaJDCm
6id5XSM/xsnW5xDtsVKxwGH1a43gDefxTowyJ6gMFZyKyHt+Rk/ZmB/nG02dT8E1etE/mWG4br2i
BAnuNGp4NmIImLe4Q7QTHpABbe4XI0aTw1hxq4kfFQGcOAAO9eDNL4oN0rL+RL4ovhfBJb4QaLxD
CLgPa2UcOY/Er2rX/DV8FUpn5Piq4nEmM5RFVRIMqMRF4SWXbnspG5Wnqmm/SK1M7RoJeoMQ90Vu
uqHlqellG/lv5L5aKvENE14NfD3eHq6934VapT4nt8fTR5KTR3cthWUI4tGlV9oig2DG4XZkjYn+
h6J/eapV1WkwhgjdFpURd/LICY3HC1XT81zCzr8ZDyrznbCHLB6cb/A7PAiN1b5Mfk4sjb6xCe6K
PEriULayRo5wlHEZZEF3NMUFeA19NW9NTiys51cgEUHIc8CoTVE6SMyEoqwwCl352FzQVRORt5RY
JmDs9Po5Vt8teatlIRCEAKj8CiKi9bqvUhXjejockOMIOs/HwWiHrTVFBMVKlj+uFzLCyjfvgikY
/GnrPRmeZ/QxKlAJE9OC1agG4rLo+OqfkdxcVq/VNAUyIaNWRwI69YairXgHtkxo92vhhzPzydTM
xN3PkzGUXO5y6VSaMfrkE2abJO8D/KC3018qHinqtnDM+HgT+mtJb7NtQpdDlNVhkL6WorDtQaZV
Da4znb2fjFHp7El+UZayidDll3Nyx4G9eofPB1QNIaSKtRjemtyRLoc/b4XC+BcaumauhoEvJSgf
/G7IDAI2m6viyNT8glZ/Ws9MRdsk4RZniicDlmvAvBGKQ7Bu8faKU1l1M7686plzX1PGZWDGos1L
Ik+KOyA7aHtdO6/QQBAbiIR09zE7iW8KZ8TH/3uxJWRMpBifdp9fCkSaBjIDDNyuZd8+8QJtOKir
FafCkiQhYnXmyQa//BIs1Ez2kZW3HNMj8IEdqLdJlYwsHfGS+CbUzrJskvBrbID2K02nGvRdInmh
9Qtyye2sn2g/w/4V/Bk45UF4nYec/50pxGckItT2VvFzvJ8snkpmIABgFcmDKEmcCo/YheHnVO2w
hFYBuSDnheoRfPhRgvgmrH8ns7jPP11W1JG81iEhkeFcrPg+XZn/ZQj99Me8phoxs8Fp1w1W3WUP
/EhvFO55Nm8Hiuk0Uhha5LuF6Zc3M8WqNecgvUZ079CKdEv2ymbs3pvcJve9EaFliqkxRROyyvCP
hPWJgXZV6sgO4MKPegbUSiD9nX+5Ny0/M1mbpPsj+hzgYkffsYnGaUzywOX8+ef/SYuxfF0q1rRt
3V0AxObH3Lej0bsKmNWgjwx5XZxnzEVkRnJKzrPh9dgAFNKEYSh1UBch06ZvOdo9MsNOPSA1CeCe
RFPNFVMI4JauSqFHJ7/wFRLbsdmKpaWgTZv5IHFDhg9MHvgo4yvfPi4s2INEZv9NcXtfxchhd/3b
k4pzdhYLm0cNzrH25MlqE+UeEtQzD6LLpa/z50zIe6hiwB3rLFDfy4RSs+wBpJLw5DcDqGZ/VjsB
tDO4ZJcSh9j3qgHms1pox/9Bfi7OywJAhpHRKI+fKEH9JD6ZqD+p62A2c/ZxfAGOa11FrdEQ7REi
nQXzEF2A7noI6Vfc8XfwhSLFvfMK1pPmZM+VRIBYA3WVkKxLGylaFpSOTA0MD2C7ma4T3kq1QqH4
dS3xvMsyH07wB+FFJG26Oli0EiHalz0tO6sw4H1TNCG1o4OKWwk8KbLr/ddrwHUqXYmllb2vrJQQ
pa44TGo3kPtYYJvdwXFLX4FPxxxPcv16/6zRHVl1wYrSAle/B06e5F2upQeRT7xp+Z49L/UNGu9x
1NZ3OwIg3xm8QGIWfUh8Hw0sTG8BF3Nc7vkPSI9MBYka9MrJ0XVgrG35KYogoX0QDfoDCpRoEeoD
563XhxACIcVfY2poQPXxvYsk3ZL5uv50gQ/6p3VZ9oeynw4tMEwQ9wymNGUx5ZHrHlSP8Movnmsp
O1Db+V1+0hUxWct2FBtHdpmfgBEchkla5ifmIA+2CDfPEIqpGMpdN4kzzB+flbGiPW+NDee121OF
NRkpUyMb6ZUX8GJq1xD2HjTeZdgkD0WjCEjPLRBirWAKtBsfdFiLB79zzTI1CzIFKcd0p+ZdaDVM
hVWXddDTTQ0zfPAtP7MEYZWEC4dPlQhwgj2iJ1If/2TZ7E3WaK3Y8cV/O3yf3uMYsjSD9DXlh/vG
UmKAj+wWE8qCvtSoxW2LLiZngQYzBeYYXQ4L9pQKMZNu6EZzoHOCmDWr632/N2l9yjkfO90Ybzax
d2mksjdHfgFUQWOWFOb93pufcWwtfZZM9f3xRBLuOhLMu5aybY6pXjQK/xyBnQS2dsoAT7qYc8yF
5YGWf+M6pmkavPaNmxXaa7sPgxtB9PzmI+27Rp3Rkm4SzcuyYMzwc9YgECEeYrMOKJYKhIg/svW6
Fl6F3gUp1t9xKzFVQ0IH+5YunVmwqPjdq1zAsX6oZN/ogAUF8yg0a48uixgHM+Ehi7EQrqaE2PDC
LjGyTGuEjf93+jqFBt++iOzB7xAcWo14E5yY2v3NTt33U5T1MpdLbr9De4xieerkxSGcUXGgX+Tb
vQSy3A01ZuU5Zcb7UCW555UYFenxBRY0nTSidvuhaq+7qFBP65281wxVWXkrmWwy3v24IXQEIJEo
K/SoZeGY7tHMFeaWLej9Z1agFuf3D0mXDvw95V1e6rGz/ovIKnzf1N7UVLwX6WO0Fhab0Fermrva
pyBDXf+rH6XJlt/Ts0GjDB0fdJwhcl1VuXklPKeRCn5ynfgzUy6omEzp8faCCCNRn1BGPeUy+Ff3
nt/BoZP94XOK70p1EpTSyFpbSoXguNLIE5pEmPQfnm5INPFqWwvLf55pzM+Ko3tDYaf8KiZGalrh
OwGT6AEL/s/wj5J2PLrHAKsNzod1UZrdKz1TyBIbuJP3lwX0MOqdU98ZqHlqLIXLFBoU2vUX3N01
pzmoh9VMqSkoOPpgHCzKBf4g4bWDVlK6lC5m/Nh79DcDEFq2zTr68A5JZogPjvpWnvKizcpduPez
CmADr3uW2kRuBjTrCOt60ua1a3E5qco57aHeXCwIyxEDz/zRxfNRKfh0A8njOKLbR2f/bFX90v9j
60jSZusGSmqEkX1gNmobejG04Qhq7e3PwCl8lPs6Q1nx8yk655krqjqVpZK+NaCxbppKaTbhKOX2
1y6bdDtk6AUyv6POSaL+gmL/a8xiTRK1dcsQLWn0IsHMQIhQepJDIgghaHY2qn+HbfWeEidfpdtb
CZKN+PODFbNYnpY+reoGG029NmxwkIwVbI88KtQtyaoxxttDrvAoBwAMmKhTpyfWg78IhXcLwrXl
7IZrYQqczivbmOve41Kr0d/tpwu9E3lPidydqsmB6DDlzJb0Dldjl53mPHYClx0v4rlcjLLFpg0a
ZyH7mVi5KAI+aGStxR1lK+QnA8ZtSNEfR9ckn0LGyXYB6LePbeP3494EYpoSdy+5DCZ3nK+L3uhM
ucYIOf+I2HFtGnQJzbqcRtsE6BmkQw3TJqTVTdnQoTyuHM6mujaFqNjILKM0qXpe2pQI8Qr55e4k
0AqpEZGAGm1xeqZfAycRRy0O/orvqPWmT47x+9mVYQzEt4sWLg2U1an/b2uryCMr2UXZW2NpkHgn
O6VgaPV6KPHpzed1jJOmcpXdf8Vw09ZsNfO+c3WlX3dp01m4IGP3u9pCQCuHSeH1CGbx1bfr2Moy
9mMFIaDeF9/86soxfk3U5kc/QJd9GZ1U6vGtykDQaK4rfxTzvD2ULSES9UW0MHfIrzAnGsC/fROZ
GquQa1VpTbVZ+LLN7VDrJ3/om9Fp5kEECEdwOqXvYDSpEMkwHaFNsISd1A/NHG8zaKZN3dMAoTb/
LeFMcGl2Vh+Mi6hCHbSy2SHVWhhgsCfCDW5floCuy+KxWPMZZ2E5jwqqzrmu2P/jhx1xNiFe+nZs
W7Isq1xdhvavudM1H+J/0dYrBsc//7vvLrrF098VQj0HHv02I/mUVmGZTQeHKFV8W1MTrCMFxyo8
XEcU4ApPXm8IjzcQtldGidiYB8vjk186wTkB7o35nRGmYEsOXowSC6/NwYUZa3bENlNAag6Vt+ZJ
rixwILvw/DUXy5eBpiH70rlF8FciCAbin5bHBp2KfbkClgjO70KApHQIlv90mLsqvfhqPhS3hlZ4
7kyp8kwl7VryUPjiN4XjGxKhDUfuwZI4VZz9yh0FEhhHkZvvek62q4CTDfKxRUq9w1Rpd40mXiyi
3eM0wjghDnNZthsXMd+7sbkz4+peNbrvaPmIe7I+yaZ5BxF0eHKHTtrio5c68yxUEOBKmbB0zAIw
8XbF2tgn8VZNnOqDpzgGcJnMdSFHo1J3nWa6+3MZWKi3cb/usDjuNjcDO4LEYenl9VfYcbtVNFib
m2UlgXlAVvfhg6cJXIsuczMc0nsHxZiAwetyZolKktgxEpybaZ/dnNdxq47fk++tZSJ98TRUy7Z2
zL5VfALgxkPi5jqgvjngap1tBY1qerQjq0p589o3b2sspQMN5RGyf04y8rRCM44kALy1AI/AdBkM
l7ZXNz3CnwrRQVMdX9XnmP2ewxsVLkKPO+odFzGroxaBFVvCQHugOkksvIpwf2nKW3Lcm3lBPkaj
ccTjkfrn3c8bSn+MGpD8z8z/SBQGi4lLCxZtoYI/BMWnu46vwJetL3NUxGTKHhFxO3/k5ejgQVrw
62goGjIZxCWFmkAhPr+id5Qf86i1AasUgMfEQG5pfU2Xa+c9vQoPSeBNqTYLDElbMCx3DpQXweSF
edGELKPes16v7proS3g975utc1EeJ0UFx1a3aC/eyHd9PCxETcOeeQxW5wDfw31CZ6wUsG085tpc
D+OH5u7TAuuJq6NU4MD+wTCy8yIzMwTRjeVJhZxvO5rWAnmXXfYPZNeYZEaghe07l59yD7j4fc3i
mcSqpPoWXek8facx+8RuoR+IrzhN7sJOP/uIAXq9e4eLDwNnsr+BWRKAHEP+PGC4bfWQYV0wF6pm
KngUDlbRTjxnV8O5WOaurYEDKeWdEU4NmPcjrSexT7aehHOa3zv+nYbGsJu91FWdV+6igIZmXJog
X/eoEyDz3VrWGTIgZ5IjK8uJaa/5ohFWTdScMODM4iiu+LzGg+0+N69MSDHWRf5As0OVaOrirtoq
PW57hOWUdgD6vO+mSorIwrnJl/E6/1b2og0vKY5BZ4Z8KrLu4T9MWOxzPY3MrrhfbuLd0AP6GAnK
dhdPPVQRiYq9ZNWZxLtAju0HkJrJAGSs9JsyvmhQGO0C2L2lU+0oUJDqK+lEBcyl1XkpYjeTQ/2h
rtOvqtI8TTRs7Y6jnSBT9EfVBSD2NppLkFG6QPHjOBE4LkLra8KwIErEUTf1t0LUPg1u0eicuZry
fhXANxF0+0srJd6qiI+B03FMd5C323A/EWWHewuKzzXUTOCeYgLNZ1kZ/CPwtnOQpJfVxjlc92Hy
A8CeP8YyRJ3bjvzQGHS2iWBHG7by4c1rYzvG41Bp1bM/rYf3byiZjUskcV5RoT+Ql+sYN/SyGy57
/ZBm/CGb+V84Ew/ffPsZOuLpi//EtsYnJoOqLsVraVdDQKqRlhwBRyVjF0MJdGxkDxtHztvnYF3Q
tZdfwGA0spIuJ4iECOMwolmbR3KjCk7HfryQ1vHFs01IdCDYEyNO91zp0iyRnC9YeXvwVXKMvmsg
0/qYBjGm5B2RCDQUO6fRfHlgBUXSrvL50LYuAT45jvXeQ2+cHaa2uBHOBWixyiiRy5/RYhP2PXdI
VbFqFsPlnHwJVeOm62BCEDogJlIWBQF+wTRLI5U1Kb59D+ld87S8Sj8YlOPn5ks+LFjikwgyHxV7
j5Ht0MoAb5p6SEf007aTba4T82Sz1JU9AAD40rRX451NkNRR6Xe6qJmowuWDSlthB90qSYrONtsg
Jve9pgqxJguroYtnWvflr+KqEswJwA7HjfYlvKBAZrb4n0bCxpswF0VoL1tD4W2Od1xE6G+8zJdi
Kwjk5K5D15L0R/Fgnr0zqrx600X5XgmwXAEiEBvYB79qzMcbaM/8RJ1fkNJLGXrljBwjofKmjP5v
XjQhtQq5PTnkE1Ij2HfxCAT37cZRMX+qErrIdD2XaqrP69kP/C9ctnyLtHPfdR3u0GUHHzESCwOL
enq+HdMgVrBzj/gT70Cns7ANGMVKYF2pFzWFQ+B4lpJHVT86+o6RiDPdh2Di5zmxJ8bR1YodNyDo
NS7Z6rqSI9CAcy0zLkv90mCwmVn22qsBB5Lz4rRs+qEGQk/+QqxWMGBnLbW1A7I8uowEjCbAdPTH
wI/jaJs1u3r9ooN+J8rPtDXvvaE2acGVfhyGcFSCgszRynMfBknUU84NshaMQ8wyI50EceMujT30
Z5jVqk2tI9nBWSGt72zbAXcc1GCodw23MYv97Np1CFHQc8cH+TJt5HBJghsdayoG+VvDzqefcSZM
tXsKCdA4kpHLhlRWbni7IXb+1sTsXD4bMzsVesmfaKsQtB937Qihixz6KGyhUNyVeD49hVPewnSd
NtgGlvt3jEkkkfen/puOephpC39aPbAvOcy1Y/tArNmQEptVLUeLcMV82LSG/CwEPhsRypfeK0sA
XS9CoOe+6yzOZtcRByv9zBm5HBtDilHCwxyJZltBKQsTPcLNi4ttUpL6L4kiUGVeX24nJ3mP2jcW
D5UddoTzIRxPRBaga2Kt8omMJl8UbRG489Fb65pbgQ0V3HiKEDy9e+0lEZyOviOvQjOsdWiEngdI
rrIQVSr/4Qxqwna/G+VmSBthEPCAbjGiEZNJgR3XG4sO++co+zmGWogzk7/oVqPHEHhVasPzHAjO
70JqJGO6ZgyN2DyCkuvAYXRAquzZEFGSLOJF1oBeiPUlWKZkIyriyQpt13PnoZ8QBr6jtt9u7lHk
rzOXvVBmxfwCqXNa5h4Y4odT/WcfJnBmKOkaiKPlfWPiAeiiUkvjDJ5jV/jZTcEfhClyAZZ4msve
uMdvPMAbbqA/rg2ogsyoRbIwHmLMi+AFDTqEAOeJ6UDLCLI0idZG4HWkjH/Ds8btifNfqwNHcIUs
JmMll88z/4lf+r9JruBF0h553ShaCz3Z63a1YtflkpJa81U2WTh4MqGEZvkc3JWDTS9+Jl86OX3T
ziEa1L7pk6Zuj8KSWzVLCW3wWsexQx0h6k44XQiy3lr+EjxctSW36/jNE575ySJ7dwEzg63OzqdW
kdxN2X+t4mCglptf+cmOY1iuHE7XLCeINkoobTpSeKCzA5hIpkt/qK+yLQ7mFKdv40RhLrA8eUfs
jGAFcXmJoV3nJs+gPLTVMXzftcWFLoJMDthZk/GHVE6/UsIoUnrh0eKtXnYYTSbtGFRuRKTnUUiD
qvHZjLGLt+bnX2KDowWUovIq5+d9XFxdhVzZamdeEn6xuHStrCD/0DKe+HeHGVnB43uUsg5/JG58
RGQrb6CdvHawHOM7+VXhhgtdITfTQck3eLNGddNJwf5ydIuP6fzaztr8aUV2xoapz4tN7B9c5ezT
mZ1nIwOrhdFlwH3kQEoOnJLaJsRs3MXS8jGbQujkKwtIdxZAbk5s95pdPFepxLjfdEgyk9Tdy5cf
lni9KNpNTg19X5CHMbm4YVGt1deqnh0MmcewaZxvn0/HD9hDG6Wzvogy5/G2Oh7Ra2BqKbB+9qGP
zeUMhdL5kAeDzj+JxNA6EMmd5cqduXXT/gsuf9H7hiV4tnIbRf9oK6S4fRwRwcU+yqCbhBF2oHyb
A0TfMiuk80Xk+9KPjoiAAPPzWDiXyGXukcB5yCAL4Ucg8m4s1HUVXkHAE0G8ltrm71ZKlgOv6ONN
PEydForkiPKPYDhpQsLmSZQYRsvCl02gK1Zz8hJCHCG8G4LKhe+WbPAXXKuCSDceJJoG1Pwzqf+R
UGfAalJMaVSjFxXjQF6Sp8oHvW3GgkvKw2aszPQI7/H/qZbEOuB7BWnRdCyYjov/larbUei6psr+
3dJjuU+vCoMr7I2/c8hMXuQbW2vBh429dnZ0u8uHDx+7JE0D0o+Un89cmXF0UcS8q6AZmVThVHpW
MokXXWXdpo2wQz8bF6X4SS/i/kvO42wmgpu96j99Mjht3QjIc1y/aBjeTa6/5T1emeV0gewXbht6
oY3h18D30Pz1vX4bjbHb+h7k6+VCqNiIMJ6Yv/+cz6TpqhgB7iEaL3L6qMZetsmJAxaDCybVBILE
A4FCid7Scu9ImJDoyJh2YxBr7VzcU7IfPoY2PEVqmKPjNuGpitVFKee77y1twZW4atLAiKDfOHTg
Uax92++n75Y5SGz0r/WHlRsuhkJTboljQZ7Lc/1xlTSlWAzN66Lch7s1Lzua676ylr+OTYsdAImr
S3KHrvMGrkZALfx1j+Lodrtl2QCt13QJP097IpfwphfYSMW6R6kIGy6xIjIcp7g9K4/ZRji/8x9C
E1dxhCTPOHP015okrzzU+wcJXmjYczhT4rJLinr8rd/CF8Z48wusp7nM7iA0YH2PQU8PAdMElubi
2h3fzysfhMXNeXbdBZy6diYGhf8ukh7e+PmyjmEtS0Q8AOquoDJ9czO2ktwTbmWN7/ySTssfpTFU
b+i6xMfO5OF8Ce9r+ZTKCEdDpn3qaby6Vojai8abG9klkj/D52eVHF6dSicZ/NhCraizAJSW0h9V
6inL2Iy1sHAqC7Z7o+3CJgrRtgBeXEjFDZRdT3B9+DgO+UOsBVP7dt6Byp/5zkaTheLntWTFFz7e
87lg81qajFks0V1rLPUWGGwHGFdQOzpxfPXuBmNJkBhyhzdzLrNRPRf7sAAxZPJMsU/gqzdFNj7i
BHozgsWsitvStYIHXUvsFnh8erGZD1fnDI+LEF/xXtnmvnSw4E86tLWuv51MIaKPdngSGwx4COif
uhzMLBo8CnNgAX23nk8wrSzmACA9KcG52O0VYaeK+kc1c383R+CTuCKu/hXoRYIO7I3l7E1B8MD/
WYrmsGGAFMgM4jyFIPAElbq9YRli7mCXb5BJyOsSgXt/0PqIm5vc9ZF8Um53oo2qcSNU/5HlCJX+
JdzydOxBZQfTo08Yp434o/mx7oOWvXNSFfvgt+NXNqzl0cuHgFqgPYHTayBN/T9gGQ9ZdY2b9W+f
fqZ+t8HIRpJcanLWnV73T/LNfNeq1TgU3Q5klO9bcHjNn2yMycafNgMTcQFd4ZWPxyebNxthZowb
wXxIzCXQDcxGG/zQxuCrmFWiQkpKaFzIoIwgJKoQ/gXXLbamOAWMt/cpD5Pk0KNNAZLxp1NtUO/H
Fb7+X/GixoByboEUoDHfw8XqVK0iuSx6B8taLyNJensFJ9g/LWfMwGxifRk2PJpZFxDT2XVbqW3e
N3cFndpXmt9LEHLnZQjMArQiQ3q5n+YcEMyINQv1f+QnX99mOmMHS6nY6hNx8Qx5+GdoJhWnYRCC
LIIg6SrPHJh43ZQ0yYxDjNMlSX3Oddk8zHvOat1UkgDDUxB23T3UmVvb4p0/1dQotLgFYO6aY+Xq
EKZprnK6StBskS/3EwaPQoHXpdHBDQ8rBQexQvfosG9kSbZU6+tXejTLslsJJqVisp5x9BlpTSp2
GWEtUEj3MQXkAGM/zkRz/MVISyaEyVzCuG7KE0tl3V4uaMlD5sz1MXIYwwJE0J9J+Fcy43xc3AhX
rW+738hdgZ8AJ2ypwGfDlMPf84MzCRUB2vTRC0iqDOIMhOn5k1CHUwoh/VgRthYuyxM2PghwiiZc
FhVRxf6l2rPhHOV7vDgrTIIV2Z55mVHVC7yAeTuObRUc2gk3DUO5WMnbCZB9rmwYc+D6aqg38NJS
EGBsfn257t3NfF2k+g0XWSTwvl1p8TNV+/Trmuq0rID9J5dj4Recr4c5yfcw6iTU0RjC/8sNOoFc
Tw9wyHaGXHzpmIWENtNwUeKqWU7MpelB3I+Mo8z0yoQaGT2SZ/HuDZVLHNLzDI9LcxJ8WWiUNG1W
EWlMlbB/U1wGYgoH6IbMDx0ZrQG41n/JpQ6f1z+dpE2jl7dddsUinO6rQY4UJsaC4z+5y6Z4zmoR
4+YCqCBpRtxaSJwTDdE653qfXOPrxRAN0J6FBEh/9aC45VROEKVPCEBLIPAVIyNn0NWurombBiES
omvYPXGQ/oO/jwCpONWGSXmSuQHHwGPVBFZSNDb+sSQoK/q6C+NYmC/uLgF3zLs1XFmj+mV76LPN
j/rRGeobtEmG0Y5jPRQJEdutw0OuL0go3AAXkJ0MFqymgygFnsIsD6P2HZ+H7fQncXChYxOpqE5o
0q9kCANxb2gAoS/zUhnf802lZMw+7aG9+QMlpeXli7hrv8pXe7KskDghmS7jJIio0wS9FukzZYgk
ktYQZHPGvb22LzzW9/4JnF/OBLVsTrW2vHuidrwiEvgfH5wQkuBwTL9JdYrWKFAXfqFns5KKdsnw
E1cRxmPn7oBtM1hXKWa75swaenX1RbEHhNMvzW2KNheJOrBa1iGJ3Q8/rNAMEbV5cxxqQ9SVSnDo
1BqkBbPK+OAN29VU1EWfaB3YyFfIp4fDZknXu1c02mBSex3WF1tcncVk0328qgFvNqlzSwSR2dK1
7NCum3ee4vV9y2iD8BNQoA9HhOtpxdrVdCHLsy9t3NLWgPoHOYoegVIArc1eOIuglwbBC92rWncb
4n+3P/LLOmmS+fqMlUJwUDHbfOhM+YmRUb999xVUxSR72lrYTyOHeoDG6z5vEinE09H8d5bJPalX
UJ3//rUTxJMz2ari2zMrJu6zVsHVys44VRUiE1arUwTnohBee2pAzsrYjmEvDw36W/VbZ0L/qqvL
DWzpYUidYqgPduqTc40xQcHFe+RO+7v1nFytyZ4X2TFgvACNSTKlPkqER+h1XHoDsYSmv4TvuVlT
QVAsCpUG4ERSKyAgl4xLAReJEtRFNchBor7MACyslHQSj5/U9LGaHH9ZFsNoXm6U0oYVkWwx7F/w
F5ZCV3PbnssCe8opfP5U0OAoY4dAAcm/epzSh5N44OHiQ6c48LJuoUGuIZikurdi53cyXT0/5L+p
sTY89SO6qpJrwfv3XjOvjLaQk2w5pW2tIQjhufTWs7mxm57xVFhnMa7WUJpxiMhO9TylLYo0UVFU
Kg4mcVuVMKZSH9slCmWr0xV4dvTRzTM4QcHhczM0rpfPYicCr/OdOPrqv2sjlnQIHI3Dw2wR3gec
yFqy2mmW/6l1IbMa1FL4ECJGiM4mgrnK4WqmytRlQaW3vL3hIdGbKuA2xos0WbheI/nktuEZSVrf
+spHmW9i+hzrbwiK+h3gbgHcrHYIA1Eh8QxkFdRufLirMS82tCyCegLY5aW+/i0+w+e0Ifxvb+md
j2dsuSYf+BAsJF/uNb3KHKGNdLB8/CgZE7qj0DXVstejPKFgNqWherKAfltqEGQFn41EJisGU4Ks
UH0OO/YTxgT5LlYcaM0XzZ99J8ksrasP7/CzzQsEPJWiTXrYanG+Wm7Fi8qD1vTmnTkPvsnFq4zB
ZKCGgTasIJnpriXA5OZqhFpGC0z2MNC+qv7npGOHUJqi4ZFrM09xNg/pIdri1MrR70+NN6ufH7ad
uB059N1x3Qs1LCzhx56qQX35lSpTHhLRbAzpd32HvwByom9oET1iXK6dcGNlTJ273xdP4abyUhcG
8CAzjLuCB2O2XEokh5jbgMoPZrY1ZIObcl1WT89c2yfbjGnzYvkr7su70BQtJm0kCv8WRMYtT+3f
E6Y5St4i7j1vmDbongP+KS2W462fbvZ9W9skH4F8oS7w6EB+WXO0PtTjPaw0XZLeuIXHea6CMDNl
DhMUSEKGdyboddYSBSTV+ijuMgPgF3hPOgZJc04yWUrXL5ApbHy/VHkqSe8pRjw2lvlRc1iWWuGA
X2VIBgI4HjCOHVTHu8zTVVb5qdSjgsqSgx4htm3QlCtTvcVZCb93TwkoAQSLYsI6NufajlYgwn+j
/PvR4oC8dRLXgyCDkSkjnBP3kbbGkNumDLWzfokR3INi4wBsMkHr/oPU2AVPm8/HiKf7x//t4OG9
YANRDQpYaF1oGZ37dkWbQqElsHO0BK3vsNM4Mt3IC315EfpHgrFGMymyPSZ3e9mqhxnhSFEUW8eO
WSSuse1tuYfZdg2HZmBWPT4imdPY8y6iGwlIrMEuLIP+3Tt6CJ2P311p/wdNE/OnMOFHkzgLf0oD
mvoP1VdJRjxxoWUETY52yeo7YnoEZ7Kz6GS384W2R5GzyWkl4IWY1q6VU1AaXKMMTos68e0dm9mx
do5G8tiyPpnL/I2ohpsnQHrf3eYd4nWq99KOVJAP+xMyuWu+XXwDlxm/cA2ekEwZVPYbkCXOwopw
btkQw+Hr9ZvybGF/YOMpKL7QXGJXPMzLfPrHach8zXsz76EhkzHFdCJk+mcMrlRHBrg+HAZpbUHe
GtdnDnbsq/O09qvOUmXHLiRcCcG/F2y6q3lw9WcGC/nnvU9M294wCOpSuif5ertO9twG5DEEvWex
rTg3dA1kONr5EZ8p3fo7qecTmKdxMC/fcSXW8p/8okuEHjS/EVf0zve01vDh5fonH68Sl4Ehe/mj
NAf9p4So2rTxAFEZpR7DUhaxw+gWTeBAw/TWDSQIpyw5MFJJth97i6EgwnKSqZZi0gIfGnwxzz/W
QSOu0VxETD0p0RtZeJ2fH+eq8oc1Wuxn7Bsqfw+rqdQMINLljrp2JwP5wVPDDz3NVC8436xm5bJX
ueZ/RCEf6GTeI4mYHlHpJL87Xtf4YjneNKq2Yc/SsVLk2bMjZdl4Zwyo7bLQApkULvpBiIGRnL9R
i93+y0EpyGZLWibYXxzbv4bVW3oPg8824KtelfQyMIp6GwwIZoSo2ErqTU3yUAp1LoF6jziRK8w7
WlrNv/k4LKZKdrWdfpNMRXk9pzYKy/7AuKcnDkZvbejrKGcKd9L92zFpMhE/AOJTs2UU15Hz/FTB
xHK8aYhZ0sjgOOX0mx5WSMoNVr4S92Xpy7qmsJJucBqImLn6EUFYmW+AjAwug8+YNgXnR7bjmR87
agcYpIwufESzITZMGZOGoLiWeKO5uF7Ob8x2TIenmj/iXuDAENnH+Uv+Tt+Z77oT6PrRZD+HYrVp
GRWlLtBGypy27RkxZ92djC+2ldzDVEc3WtF2Jk5yF9J2jePALgIGK0Ra/lrk+2pQhAZ7sB5hWcDV
1YugOHki8m8zr+mKxYe0WtGRFvhvM1/FelL6t2fmMD3SW4T/8BvhVUDO9aGoGXxwW26gJFEzMCcb
+JhQqx1XcZxRQ0PluCTGgIkzeRPgfu9Nq62g7lIfDza0m7azbit7sQwT9xhAz11XNuANIqe8e6mJ
eZhRk8TzTnm3lLk9RMsRGyOE7TZ82BlquCKAK2ZWQFavNrhoLQIytPm9+Qb6gA5qDSf5QahcffoA
j0R9UYT1dVLRXKZ0AuFby2E0OPGQRhh9Q4aZ2zTb4XE03FtInjQ+pgrjCpB+HsE7Rq8vKXdmfsXI
8Bt9YrQxUmFejvFQW8l17CL8z220TaehOiWVcMxBK0WwsPzoN9NRYSaXq9wbf4KhM+LMs2jr/PoO
g2KmT+vVo/f7dj1M7MBm04S+5ePKB1FrN4vfhpGkJPVrDY8vWIeBfQBNCdTEVRvw1kl5yQw5FeOl
62aP7J26eoLWQQMvTvKdnSn6gok0s7j/b8P1M/+DpK5e/1vN+o7UiRTiUp1Vir2ZGQGqSaKWsiXt
e6Tb+4wCgDUiHV+FijQefjbd8cRH7e15S8sChSnYnRvIVyHq2wW+y1DUcjs0GM7QlRB6vjJg0l6Y
e7xi6tnSOSDKn93syQiGrynWzs6prg5mInAB2NyWjyO0a4K7abXMUxTi/nxrtEZKtccGpu7A2nbb
+2Q9klEtfc6rsjIMMszkLnjqTusDWm917U9byWVjNfyx4RXVmu9aZOvaQXE3jQFTNarMQFZWF3Pm
MAeAKM0HyN9YCe1eKHB3D7tEGUpN2gJcQKS2BByHA0+hCvuk5bwGM7uSMUdyh49+pzWH0EU3u1uo
1YLUuLm6s43zaziP4dTSJ7otwoH3TZ7uO3lecEkPxWFCZqBF4l43s2aqD1GgbPn7MvfPNJAwcfSK
t1IsijFMb5DTnq0ETcwVVeO/0l6O72wPx4PUEY5enxv138p4e1DCzTPjO7FDkBcTfKL3AxX+FUjj
C9sTKWLqcYY51toL3nqePzjrDnvWSQ8zgtkbLlVA4U+GNrw/jXzOzLKKzW5FFAZeoS3TrUWpMAfG
C0Ur3ZjwVIDfeD5PWlubOdQnibWb2Mwd3pd++wfXd7J+Wh8w3SjXLY9bZsuKoRxXu7/bLfP1XgIK
GmiZpMs8QLIgpe1CvDCOhaYgHMmKnlz51JUWn2+MS9BBjwnDN8wB2i5p8k61c89RGOkRJ6z+1TRX
a6zLt5PGPLn+eb15hZbkTDznovuKZhFnNmO/sh4kCLmEH19LaA1VECWsafyJnV2O+8e/ScQwLvIz
TU5rnGYLzyrINBx1mGld8p/u743I6z1xzqjZDm7+bXeXlgUpQycFaimphpr6E18IzIZ4vLI0Oeg4
9NTQK+QY2Oqv17t3BdNT1sfD38ajUOUwgByVNFAEnjpb84J84VanOUHwc8ilGmLDKO3owGo1P2++
Cm0zDvJWc46BdNivWaE+KCVGu4i9K6T21cs2mPjgDicB4kNdUjh0vmHTmLXO42GcZX+iLKQFIWTr
tPaY6ltrSue9NMK40Jg7xp8lnKfmBxaebWAFhQ5wKsKrOO+1BT0A8rJW1KvPkgG8kdosQAW5rscZ
T2nmjcGCGzYQ1zCpAGH5V5MtUq0HbT7o/lTWokkFqqigWir5t6BtCXb2x5kq8/kF2UzgGCn7+uvn
5i+Lgph+FrMd/cs/dB+WhJMJd5TT1Z+by1MnE028cLupbzkioT7+x2ZhqBlPgXrNPMpVbupLbXNr
wCrptwqtdqVr24iRtsJqZ9hnUF0DAxazABT1LBKcT/AD1yYb5QmDbxLCQe7tumIDqLge+fgimMiS
Rq5Oxuyyp5bgFeU33lWpmem91FdZtQY8B/xxjKUxacEyqBigum8EMOZOhTzGTC+QDa8DfAtN9fGz
5WZNhzKHpSzyLRTrg0CWnlo758GGfqBfB72jRwB/WXACKxhAZuWf6ncKgGxB7a7ilRYgRafnUpLd
9PTJ5hEDyqeVkFjtEGDvY7xAgTJYwTg2k0p+Dg7Ceim5BoKsGZxCii5z2zSDHbaHooAjTyCDbF72
NX17QZOtk2FqaCpSZSSaS24MlH+wn7EvRDYHdfbz+GBZjmnBqF3vuiMn+9suua/kQCLsd4+eE5kn
lbL0Jfrb4J3wiZCj+/RkgIMLuPJ6cYIEnddR7FDaQziyy1rQWhhHKLQKwciSyUARdWsiNTjdfnXf
HlW9o7bW6r8EwZorD5EYbiNDdmR6j1zz15FjujOYHHXNuGNkH5JHM5oZvFoHCtIDt4JBgE1G0AK/
05VysW7qx1bgp9CDAkQweXWW9zrFUgW+kD8vGfAbVW3IA9PEB95Q8O2R1CPSSRfPve4y+GET03+n
H/LUEy8VjfRmHf+rNdzIRZkOi2uDAHSJGLM7XBW6xXKpOvT3SFJGTw25ErLItqlKPDAe3ZfxGh4M
5JHYL83boDsFvR6l1mqkR/lchdoDivl/xykwn0/nUVqN1LN3aq4Cz8wQffNbqPCAnrXaLiPAit2M
oht5cTyNtjqiHqo9brRG20mpfKpuOL+dgUMBc3JO4V0o8s6zKDdF9dOCEFReV+sM8+/JBlcZFzaY
3kV5auOzpX3ck9iqpVosF1Tu8r2uC2vsCg2zJPU8Ogg1GAVMed3g3vyFiU0a2ZeObYlVbCfvb+A0
yqHhPlvC4CCV0GoRbRusmfEQJdxxjPK6vCyDisiA7c2wqK2pE1rxXZz+nuJfY8PWPjRJnWk2vtLN
m58STkQbJ+KclwkZmedhm+4WvJZjNxJKMM9eGlfCQhe7ZA0O3olkjsBcuhcYdCQIfa0nxH9iL1PO
l8/lw5uS0acrAt0/Tv6G+EnU386Fts8zILWjFSsZcGOUhXfTrlDve8E06C80SwYWF5T4DnNcrKFD
iyxBdxSHzO4bgvEqbMipawEI9MKdYoGgTpg7RPRjGHx+c7Ym/m6pkKvdvFT/hAftJQscMbBCdaRC
acLTERp0MxFWW4gTCwUE8kp2rneWhLmbcuJnT8wVJcVJPAztIxrv8go5bnzA1Z/dNOaM6X4r62e3
NFxnYQHPAlIu4WSKfPfly1J0ykNfBvfYIBrG87f0EMKU23wOkaUYvCDqDyykpQTBlwZrfSfjKJR6
rPaCTyvSsP1YwAd7aO+Ye2wGTvfup/zYejAXSZOjyAOVzsy04K71O7LW+ZrIMUbLS0V8gskFi9Av
VBf/LxfCuMiR5ngM9Xy2j6OgwsJKokBdzvWu1VAUYjC8xAZJJeVVhBUEWP4blhEUuH4FiJhFIixU
xvxmaGwSqqVYYeofD2gqPzf2mY8DUZGyiVK6kwmK4vv7LATCj0cDqGU7L6F0mp34ZSM67e5F7pka
Bvjz/3uMyTEbLn80iAKDSnO8gZgWCtpvOupknFX7zLUHuYCtop6u6LxX4+4jILYLoOsifuGKSemx
3UWyHkyD/7nH543V3/Dmc+JWMLHAs3QxA5/UVtFpSjI/clPMySJRGTFOn7OT6XWLCOAhX33h4IXd
jbSw2GHFO3ye68KChP2msqreRL0qehYwI9vhSnPzsUCkzSeksr6ct8fsr0BCFq4loeVTqXsEC8LT
9e6a3KwpYqwoAE1ja+LD/z5n0K3OyQ/38KS6f+ymLpTNj9rU0RdnI1tW9o746BHWBm9zogSXlgfQ
L+tckJQ4QbCDN1c4I4LnwQ+jMrOMazJB/fV9wMWiX4r5/LEwMkr8eDGuG0RBT/qKvAxSVkmHXCqF
yzDRjbd9oPa93j1Aa1TaFJ4F/lPlw34X/qGfgGrYi3A2nmYcxtd507sjKd+leaHCeExovyd+SX1I
jaQpzUO+I74+z4KB+iSy44jw4f/J/8roObRu4RDEvrvoc2bSzH8i2d+XwpD84dNlRIv1GlyzpAJR
YG8D6aSFBtnq5sptfWeHymroKwTHuhEuSwi7xw5JwllKmnFGIyGhdDxv1hcQtOPC/bwemI1m9If1
GSaQw5mn9sWsLayUvMsfhDqLRIncloHw2zBoEmQpkHL5jSfDRQJftfj9eFRRXZNfe9GY+VhStQFK
0gJWCM/2LgvlsXzg6vpAyHZsf/cC96yGSFyRGj1YaQ0UXbp+RgfLf+XTLEz6Jzz2jz2VaduNY+1c
Z7gNOkTXwW84ILFQMzD37h5m/qPBjuZKexMCgtVl2j177E4sYdPHK60+kSFdPkuM7apapp4NfUP9
C28r+z94od0jqYv/h3BP/SFdUmgd+kYIQlVY0i8UdG9LFGOb0Ucj7K0wTA7eah6FQIEh8mxr46zs
6NP9ns4CdZfB5LzL4SWcPPJswwzNjFldXBxrHut0czebBZBWRnE9yj8mMQWtIa3MqEstU8jtyMoq
l76dyfg2QBoijW4kLxd7BuJyWb9NoPJzFdivzSFOfjDm7lSAcIKvUPAGKYzVO/F6wOdkSQaBcLzD
/VrFX//u2pC8yw7jwjQ4CHXlyDsxyCyIvWSkmyhgLQS1oTj2QlEjmyjprprCHXnYMDxJgFn/dQb4
llMKq0FlekfQRaTp5eSxZu4pdriW550SJ4pwLkGH5fJb8LLfU9NTFGAlTiSFV2tVAAhwXq4IYo9d
Ou4iXZSsezkERe1AnbH+AEB/7tG9XjTZeyI+7s646TGbZccP8AzIv6wZXqZzYbPCZxIab4Jo75+t
4qMDX7VF41z4fU24QtzT6qun1KJl86bcAZtwWXYtQaJPU9GDAzZ/ZiOzhrilFPEh2SkMIUTLxIA5
Ck+lrDwiTs/OHxTa0tM1GJFOzulS9xyMuJvppwExQZjBUVsjvopUrxemka0/Cjq+tMBDwNfnB94+
UdkRp5qTO8BIpdyJx9woQ7WX3JVFfppsoeVv/subKO+tNO3qOUiCRpBH1qsBlrHWl2Q2Q3p9VvDC
up4VMp3Nv0WfrWwe+g4EJiUv/LjciRxB1GJAxtgHthaU/dDhzzuozBRAZPdc7De7oys5RJOGCZhB
xXuMAwtlStY27JT5xu/HUgvwemyoNGAehfSD9ZhOiyaiGKWdsDWdmHuK9IaUGkewRrplHZ9HflIk
4/STsp6XKeYLLZ4XgkAf8Qto5ndKwG0f5/e6QYi7Pk/rwZ/uijWwSBdl9Z7bWdpn7IIqIbiSLs2/
zOpeGeopEVchPuBrgr0GaCw52m986qq3F8G+YRCQU/GkDvlqTru2slMSRWx1OdCd/FoKWOpv8G+S
EKgStMw0V4NDEXC0N9XwDAFMBtPo4auAsVQhlIbhj6bbZ4eW/PekduV+og5xSHyUApl1xsZI9ccJ
BaBd5nb6rrr7z6URewQMQp5fGLpT3fMy65j5fSIejyZAOAzminpD5Dewd02BoD+U6oVhd+U53c7q
CvnQcCzW+oxdPYD+ARIXGZTF/vIhrLC+8Imbatb6+QOTXb5jGr2kcEIFXPphxeytqIXRytfdmrk+
nieknC5xhbgwOUJLqXF6iFTBFyllTK63GAAuVskLRydk/0S35usKIBLN+aEphcgeT/UtzybZR3cb
GHXchdMveHVbKmrIXP0gK+KL0az46rNMU2U4Li7Ksbb0FlOITCvHcke69Q3Iapd0yfs5Rp+xosjm
lhn8z53qIBuLvR9WT5PnmiuO8gZ2VpSztcYYkNoMnij6ATtTe8n2RdIlTpydZDPGM3mwTNsfErQI
ppAYM7+B1ie867jen8GQo5GQ/PCeK4tFOWsArLfkB9Ba1mShYu/jbmV3EsdJLEZX3Jtsl/XetSnw
zUbe83ZjoUqqlKvJUfiGqRPBPStK8S5kDpvCfma0iZ9EPXLu/GMDebjDMu3I6S5HTW5GG6r5L9Hh
kvQect+oXy6oq84QRnZh5aApMYCkSNSPglS0k8efFA57cPykLc0wxNHILfY/YL6szOjm0oDbkBKX
26IIQ1W4hjh3eHWR3IgVe1RnQY4MisPWlxSXTaFokZiNVgq2fPFOXaplszdsx99gbL1p+DJ3AyeK
YC8L9/DlWSXEbHZIxBI+GE0XCPKPukEwW/WTC3wG2qaTspDznfrtJ8SkJnJYvhQgTXn7bJd8QDA1
wuZdo6tL9Zu7Tg9jmpCoyp4qyN8ktswGoFhLV00ODvrDAGqWIdNWsXndkqlUTacocABHUtLnBV+M
ccApNLQWdA3bsiR2IGSt4aGgAmOepbe6vj60VH79oUbB/O/T9E7NjTwOWG7FDuSHajckIOA6LPv7
69D/hlkdMYjjYP4umBno3Kk5gQgSIgzwOc4x1ztsed7LFPq4ACpYtg+NavJGNHADbvR5LgilaOAB
X6C1d2IEOXAixX6Kle2k3xmkpODd6BBBbRgmzBHCEoLMbnYq1hcZZCyq/j17bYdrt6o5k6ceJ9w/
cJC0d2eeTiE83tWuv9f60+9eK4vikyakU5pU41UITSp/tVm9ifU4vQZEPqgPvslT9Lz0xZcDMKqV
CoCcAdgjAToWsyeKM7DMvzA9KtEHRHQXGGD25gkY/ffFfM592+GBEayFTNUSvuDklY/dKDawaRG9
ZndoCtAfefn9SD7yPIvFBKCD5J+EexVmlo2zMs/yECUikaZ5KySspPhm7XzVq7ns7+yrCH3aQsN7
1xo3RYccUClqQPPtTb/WpJMzl0xq6EzuGBgts3zD2Os6lY82P0wfp08MTcHqeM/+82GdGlIQr5vU
URC1iQtwfqTTUvczxq9bxF03zWiAeqf1jPz3fYoRyMNQExejwOcb/eG015xO3QcU6qtj5PitHKAG
6IgTHfbNEEAj0Rrzw2BnO3ubV1yd92ZSUS+eUdtSOWAr1hVczR30v4sg4h7M/qBUVEsYXCMcmY8D
xsx6UoL9eiX1f1RNy86JidU3Y82/ahfQyXw4pldi9gIZZAcw+ruwmFa9U0dBafi9jrbYejCcAjT8
xXpDJozSH7aTxbPq4419usyJ0lCCDVpj8soiCI2q2qy1ugK2ggIs4ehOn24E5+Nrehd62Fn1lqN2
/ByyQaluyQ03f15auZpfF3hP+DU2j6dpVKzfuHZfmtTDkxYMq8HgByMK4iGZkrJG7DXNciaCPFgd
K4qexNZI00fUBQD1Z7mx+ZBINOl5ZXHCEyTPt5acIel1jkwDHl1fhacXLVF/ct8LZXGXd+saSOwP
Im/KsUAG65d75I89uyTPp9I8LaMrCn6OMOlXxiKRpD0pO0x5dIZxD2UJZSXIwjLPi6amKVtA2qpk
bZnnhQwsjFEQLIWcyyaptoc4dz5nUczZNC6WQv2Do0nmDcpc9GQOjgE1pN8ohv13t9vcD1XGb+6p
codqH251vWyLR/j59TloCKNqCjPM7cnSFg1lM/mcKosHbTcVZ1AHg8itbkS41/hftM2E8yzb67lZ
SKb+fBEDcgd4mm01nx23AUDa1DcMBqOiQLO6kMYSDhb/D/LBRPklPqe4hoTqMrGZPkf6qjrJBdrg
+1+Yfj+A1rmBglsvbTqSsjyxs0u/hGz69Rd4Nm62kCBp0rxZ7pm3jHolZXn8iruQmUrzhslQjW5D
Jv+zZiAJYGLrqn48Ds4/j+irnOhoNP5sJjfwN515ACd6EoPeixeVfVomxL3BYo4Qvg/NPCy8teNy
GDNqtfIE6GZtjzBLz+nr8TghoC21gtgypcq5s1a/NpFG/VQLlsFmQgLGlvtZDfEfUahvDtdXcK1s
gQXBJbfXyLnfQGrJHd8O2RLSG99UJmwLO4V4wHFXMbPUEQ20P911nY5aw78nMI3i3tANxxlaZ5ba
62WuD4+/meWuZ5BKvKaqOnnopUQP0vyQ516PTssWHM/oTBgcW/l80cPXKCvz2pasmLA68WyxpBRl
ZpGIUcU6rOAlCs+EmFQSI8dk6MPGmi0akQjNx9vTHn2bY063UD2rJUu+i4Ss5Zj2QR/TzTS7zQv8
j081mtImXJykM9jDRUQ16ov2y0P0JM4Md5DSIi4fraCCTd74OiWFwip+oq1I2ZOO/AcwTJHQ7WQX
WFb55WdVsIDm4l+n9GBpQ6sfReNa+OlJ4FBvlpY2StNkbhndzxQTFInz+C26L6w0OUtPBwqQfd4m
I9WefOM7/3pwmyXMq5/aVEwPt6cOAk+4/aVB6DHB+MEJdS4B/TS/HJ7PibPEKavT6LYedeIqS+nU
J3XqjFb09K/RXHPKIntmRpG2w0GWpDPESVY2dXwOF92WBO7LNcL/W0B8ymIng09JFZx/WsEkEEef
GztMqISm43nMTolJ+Cvntl6d5qg2rtF1CJ87GdOSAwOHuUI1vYMLmgo/WvobV+eiDfDdQR2g1+qX
AmSM1mLgkgPyccMUOxA20Z3eFuVejVawIvT8F/YABnHjBW8NfLQv7Mie4AVBmiZ9mGcs10rANO1w
0VMG6chuhUrmXaHG0OARKQV1EkhiTN4NUHCXK9f/dqvhhsffg6FJTAanUjb+cQ+cTlwxR6EkCvip
33XDEcTMVLg27Ozbbdbjqncg4amaAf9kE6b5Jrac1kVm/SqKPLMw4jg61Txdta/wlMjBcv9m7uFN
eULmxNe60soUlROXOS9NTPxdRpyo2mly8JeA7jShR41ZM4JJCXrgjU79JYomHIVVOsZTzsyCGq9O
Pfw4UWTcuYTXIhJGozJAc9VN16GyEaBDxB1g/Qx5Cft6IeBbPGjmE3k4OGWEqu+/FJpTtiSGnRFo
nhAYu2of6iWLUhbGFb5e43zu5hYJ7KDOJfFHGI2kWdHfmGoA/xnNuk7/FJoVs0qzxcY1n6IRMWWy
99YB4HlnZH6UnmSjivIIeKLVnf292CkSkIaGi9ihzPf6phfOxY738yeYz/iwKwBdczLDpQNMMZ2O
LXauVimDiGl4PG68uJZe2jR7bNye+QrrtdkZ7Ups1P2VKnI3Lox4R5R0kg+PLj9JT0MldMLBOLN4
e1lL98rNXhLdeOkLSSYa+5j/H5tncJyp1TMphNpDCviKhY5oNnxFuzjZPzMAE2xqcyZ09G/1LT0f
TOSS6u77LzBYGoL2KN5Ul3Ieob9dxxwnu5opxfSlSvME0EimtYaLTbUIZR2F+9OAPa4YCXbxLN0Y
slCNuH2adAG2m6l32lysDOSYdcLd70sD9JG+NJ9pVtC8vBHhI8yoL8lXn3yyBZ6NT0E36XO/gPnl
gtq1LAz+gD8l5/agaredkJSl3q4r9EoS/k8J2vKZ8k3SdFp9JJRNo9BAyvzwxrZlJVT9ad2QhPwN
ENyO1t3Gd7cIBi3JeDvTPRgK+utU1TAPTDCr3gf8BhOEHrc00HF/b28mhmr+5D04aNUmbc+27di8
D3fuzJvnSNM7QThjOBD1mN0W61i+ztGl1+9y0T2K2x1hxKaIgl8UPcQ0OmR2oZv8zMtdivJZwtXZ
SNOiwQTYNBzSQblhex2hgGWvDDSdZ3Vx6TdaSkxZ14sziVnTcJGAXt8Gh2EQ5w5qNaU3fKkn/abK
bYzatM2kOAWhoTk6VGQFoEairTKPZgJrMiQHaZ6lduKT5B9VgtaS35Ijui+cAE4e6bfrM/Oe1eFD
QHZgnk5vCf4a5sdeSfbVpJg10PIS/LkXEQq9tV0351ueTMHLTbnAF5DlgVCs/Jgu1QthW6Wh19y7
MU8sQ9zdmdGqAXkNEqBckgNtmqjuawk2WyhkQG+WUx60cXMsb6aTsiKX03nf8dwfJrOIY4FdmqZn
T3WVuW+GVYE8WNEtJgYHEY2z5IAFN3/hr7cPvgbNqC80Vm0304AMDbaeowsy/qR8Hou0TCRAJQHd
jci5VZoHpVh2dV0c3yQrOdhnN9Nz7aqKZ4HNSzyoJ2xjIQH02jTSTm9lX3PCa0baNNmlAn1f89l/
IwfHhcIGwNrJsP6KEQm53+Hf9RmfQhPZqqtdWZCGFER00MaP9QcKTafLSli7QNqzQWa3lfjfHumE
ZecnSlXzjj/EXrQ7FuM9iejso8in6bp2yOX0JR0Bb5zREAhp4QYFO2/QBhhwoR4zTepRQYnJdnJ4
6CvJV//NmTwdmkqM4zn1HhNlo5IoVXssnIxRFFizQAD6YtSTqL4YUk89c8ISuFxxoGs5VJe7g481
YuZApUKOZyM7PJRt/HlfRa32j1zweMBaxKWWUf8/6pMU+Or+nRaHT1wmhpjZ2WtDAljwXwYJkvTo
SPKNwpImLyMe5DiD2hDQA8J0yybK6zH8GQCqKrX5wosxUcreoxAUS1yzPcSbfrOCudaQ29aOrv6A
AsvBnWPQ4lO8NwxNKl+x6N//9NgihXnWcuhgy6dDe7s3ZQYGNqaAf11MwPyqZSlBH5Yb7EWWua9n
JpNG8G/MicAmTRCbLSRAyXkCvHH0NVyrmKdfkO8XvEqAAWa12gpNTmM1005dQLK2vMjyPFK0mClu
3v8uKzYXGi8d9WrPVWDbPiSoilAMNoSJR9LaWQP46XgtzGb/JsNKLtYsGhWthOkpBbKUSSShX3eN
YouBY0mrq8iAv74IYhQBUKmtFU2LhuRoYcXUsaPMyVbOMkpag66qgkQvcefxO6WgNfRGqCukn1eP
oVCHt5Kfem+RqYOv/vPKUINFRFrSsywYIhREOQx6i98Tq3AFQuCx4wkxOgH8ypQw9RDGG8UuvNM+
Oxu/Ddw95ovLYo/6OVoFU786SGq1HSJZVaf6H1emZ/Kp8oyLyLWFATEKORrKoP6lgfn0jSPgs30+
+mx912a7EA91Ipoj/JllkMS0TXM2uU5swhyHJby+X8soDrVw+uyUTu/RSaMMHOOug++VbJk1mxOF
Q6caXK8kANUZuht13mn4H9/zFZqDr2thZKNLOc74Ms8nq/q1kaB6jIsPsw65ZoCFDd6BPzGxfPIy
p8/HY89db3RJZ95ox5GDzNIZUkAIX9/wOqekZkLoGCHmu8bgzNpC4i4HHYCgjLrtu3mufy7X7AYK
4XTQeWyMbKK6f7emFPEBkU+SttjVrqx/x02LDRmuXYlqvcMLYBkdbgaQCX7+NURFly4RjNqJ80ky
3f9Hf+/DH0DZVNizlU/Vt7xuBosq04Iifuwmcl9uI9R1uzpEE8XCrdlH/RfbQUrjT58Kcc0V0CH9
vU3i/558N6SY3wzNYDb6JXk0dB+TPUc5h+fExLcwVXCKUN6+MCl/HsrPo5oZmG6/4kSjztl+4axF
zP39FJ9sYjETZ+OS+tFNOGFhm3ZMCEA2CBy9BPd5ASvH5+u+/E25ToEJJUDEtYCgeiK4fBi2tLpS
qkAPCXsMbPYKYBJuVPvLFfBDFPPnEsrr/9rE4iuvnA3CRcLWWdWcDpAh0Rg7G8w5uisyKVjVGg+m
cej/LSjt3dEcJsnnK1EmHJ7/OxgJvzac17O73Rf78Zghd0lI+QIxldFGCqut2mAQxJpv5kVJ8NfV
6mvYm8e9t5PMRK+tMdabVsRP0P+vqIzrFK5WJimAhqALo9FLoXyowXX4gz2oAWa77IXVg3fuTWJ3
RfCbKUKvQGYutiFX0iqHNXbipLu7ghD9XxqX87KU0tdEjsX6/TIMieANKs+nvUvIZXrKgPYKD9Iu
MzcTWO6eazKeSWvyCofgRrEONiK25tvSj7rJRYoOvd1XikGfG515gAXyj9brrhQDvndjZrjAfXa4
DbSCgKEETaSUPnplR9a7jH7KTRHmsMwKCZbMfez1WFDLdLojtrr1rJxvtJXj0xJ4eNgUeZu+8igc
yB+Tp6t/vB1C+OGiLXbij9yfx+SxKzTfr7yGn4lF/VTptrzK1goLpQdvzvJ4oUqiisOyw/YYDhVx
Q4ZwJTwszMHnWV+8fToexcKtiowE7306iVTrCplyM4JH13DMrPxFh2Oorlh18vDu54ZOTvHLHght
X6CAm9cy0N9NI7M8ZVNU1kfxzuswBaCNDX8hX88iIpjK/4dyCOJAXVru3uVqtUr7LkitFitVCjIB
WAjhsBkuOK2EBKhPXsHmZIAc2tfIPAtkR1cSY3twQFPsHzSqaMJfUqmDMWGe25iSP0JDV9r6xAlQ
suS07em/5fUPGuikuZ7+q1pwRCUErKkulLYbGb9bFUSgk3UoZ8lLY/MQdNs+sJPufzAllRKfI7Hd
Qm6o9+Olun63J1E+G93t3f1TCZC9s0dmTuuE44KLAARjMImkABwhJpGfgyTfMcesGN6cFrRR9A29
BVGMnv+Ljes59fnTBbRYHEAD3AhDEs8OFjKyyv3NqDpcAW54/amhLjOSeXE6Xr/PAzb4vPCXDCme
zAcNw368+xzTojBlNh630q0+vY7UGuG+he9lTvkj7AQOI8zHFZDShqZJGRCCGw/MUPZaXriQvWXw
HRnZ61P82wfwS3lKJBWzbczIjBDmn94j7LoF5cU87fNOWjKvmgd60oikN4TNglIqL25g/iZ/wJdv
Mb3gRUtS87Hlk4l/DeIcW5ZEaG+Ihgv4OWgzDlmwhBEnLZSOa7iAk+baQ2ob03nr98u6MCjMUMLS
PALxfhfgzSJrlOJnZtBbJIqUnprJi9vXFAK3LqwOJKH8a2vo6iuzq/M4CsW7022Ee64aBkuVfc5v
oDBotUn4xJhQISX7HDlH0DTbESIdIRSQhHaVVTq9CqQ9PShR9j1AM2B6FOFZL1+9As3y0pxduOTO
xHa8iw8ew3kQF+XwJ+b3XZvqYc4muF5tK1/01sXSoEJHRsmsCYXMsIlBU4R22KW0g6un/2XedddG
TuMx8ostui+WTD7pzY0epViexCw8Y4xzWb8MpmdjCz+XIHx8yoO4QGEnIgKtXQfjOz/8s5a3tfSw
Wj2X2lxM01NmFA2mYHbiY8fRV0tdBEmc+l5OypVi/RadhlEhlWANzouT8hZD7phAZagxaNkiEY2m
YBRW2xw9HLSX9bMqeVVs/j+YiiAcvLYC0PTfWcH+WanUxY+P8vs1dEoQehYpvvVFEXoH5s7T/fzu
pV1AGVc1O8YAwYPrdNFr0L3ufROahB03jJM1ecktxXXJyYyd2CgLUrMpRmJ6mdTEzSef0M6Frno/
HvM8XPsPSNKvpTONO7qhoi1wgVfYIK6QGA5EfRvZ6m2kJSzc/VPb2t5ok4jR1OpiFuNOpk+hhEgm
XTRxIUC+ZI3/SO7RMhoScy0z9uCy2TZKs41eJ/63bOMlL5GSI22oNkM1xBg8d/lyNzngeg6tjBjf
WLSVe61r8EplVjhOu2IIO6zb3FEf44LN4r0AJj1/MAVn6OsaxOGtiEku2MIP/bTcz/MSomFsCSNA
qdRfmTT/9S68ZdCg1yCb/IJntiY6r3uW3FnSWL2UAz4jakEDZYyjnhPAA/BJEFZqRCo8pcaEjbxt
kEuXx4jqvb+pPUN8/kEcwixVcg3iJulTbJMap7u/3yqbga6EVrW6zzWYco8mCWyhW7z947BTPiNB
5flVNg5EyLvo4MsW/igTtnLTKUzPCoKlvCXaMRiqiMGmWaKzm0y6+WG+J1kA7uY12Q+fmkhLnL67
G6GTgdw7u/PFqeq3v2hg1k+3qk3LisoEfl4frq8cGjUvS1w3So7I+4FragOb5Z4SRYc7tklvONGd
TKPfnn+zl8WKIXl/lR9GmMvXGd5tm6vmMQyfUsOWwA/HKECHxHPB7c2P+aSnFeHS2LpB5Bz2HTS7
7SUo+288jFKzWpj7F5PXStfASYN28BCWGGfV1rqE/o8EXtZGkP5etIFXXbuKs9X8/rMk9tAgO3LD
CriUrYmyqmOECnqPZxVS9j2sE0bJ7jaDLiwRutzmpG7aBzgTC0N7+GQGK0ZPmt0YMnTnQpykOR/F
uFW1d8Fos8hP7A1XwNOHNVz84tpattsgTVZtEjzEgcfmH0aIss5XVoAWLnju+m5CzHn0trl19jEF
uu4UrIA0onSrQz3qK1sHFSWdTBood59J+UbWvaG1TE1r4p7bu/hoKHl2QiQ8wNFx1s6FnMbsXEiA
eBm3zMxLHgAPUSAfZOORkhV9sIn+Gx1h5y+yWhivSMDmZ95xYoRw7/J9xzzPXRdt64kqRFH3GE4u
rfxCfK0psrjjVyU0VHjv2S0sshCIUVNjiGJmM+yx6QrB0A1WhxIT0T1pQDS6njkCjAzjdrY3MSR7
mton6m2lqYjxeLTnhh4irEPLnVNidSTWcZ26q6r+PXb7NJVZukuTddXU33dP9GhEL6Cn0Jkoa3zG
tAIiE7VBZzJaY9nK6G7/U96QxPQFo+AvibE+5wjnKwb4IoDQ5sdr20CLr/4wdckjfHX/oCX1x4Cb
BT1cvYRl3qZs+KkoofHB5ZQt/tjiuQtK2WFUmUVvW+PzH1lmG6njTnpVvhrAzb5p+ElBxrla2tm5
2AgbCx7JD0F8pV7Bxs8bY4wryzB3Xy4dPQT7R8Sbpz1zLKw6J0c8A8bZh+6+B4lsTdYX2hmMhicd
TfRd/tHVyDTZemonrU+XGIbL9HQ01eNE0MWx1BV+rlvIz26Bl/ssYu2sNtmCrSCnqIw6V6T8hPdR
sANIZK1vDAgT9Ms67akT4Jy97dr4Ap+hkjjsjGDbYVnIAN1xTyEWfAfljdv5kXE1ctH4XZXvZxvU
62t5CIAzkzp24e4nOPlt/X4v0qr+Pz4MImuXTAm+fohlGBCJ9u/Y9o9Cf3P3rV6Gy5UK5D+fPG+Q
skdY3elgFV4yUPZUnMwFcBFj9Cf6v05lWzZ63y1M5n/3Z099YI7PaSbJCSBrajyL84rbBADtjkKr
UY8mx1QhzprRX/aOSDjM4Ha400RUNiNK7VGEtv8AwJeOWcOLIaJZvYZW7qOtvAV3Cl0W3E7/ha3Y
ffSgVMOH3jqLs5GbkO/5HC6+3Mm0O0KYSGI/HmnvpRkWcR3uvsmNFZLpCjO+zWXT5olrOaeiO5fP
qHKIFVUhsQ4r/RVbgo99Yv5A1Co2TD421waiL1bCp76DewM/4zol8cqd0EZ8BD2i4KgjwB4M2PgO
WfwkjgUce+DlJznvrTNhsK7JAIh7wJ47QLL5JED45IUjNLioNPtadxpMaG3DOQMACQmxF95xEqWf
2IKvxVJvMxoEVP+SFIbbd+RnR0T/AMu33VWwMJ412bVqZEzFb69kA6AcwUMhjl+7mh4ny1Ea3lyC
3sIjBydGmOKiE4cvzBJywLBDs7S4tJKvPAr82EMETU5R3JbTeZ2aemKl/KZ9XynEvXC70q0yUSZC
vdC0sddSTVNAkWzFBkYdD4cZnjkpSszA1pCVX6Q8pK8vmJcs/bpPcskrUfpGegI/MmEDCjx0gbE0
biQ4972ZZWn/XzK8npMbUyIkBSCPcn3Ld3up2JiFYQsBoHRmVfG1k4oszdTk3LbeWC8pL3lOVyxF
bDCCycqOZhljfbH2fFMyq/B8zkbdpiZdYKoihE23xZ1E0c6iUvd7jWSFgRId612bILlzCzVh/wOr
fygb/TnnYf02pjlE7A1FP14JRatmY8VBTwFx+OdZNBMj7z9p7iMBImx7bv5wKkeHqoO4qJknnIbe
NdwcnfxQBWWC6rjoip4BdAda5TyxKVS+5gRTw+cxD16oazBGoUCF/yux5vfQ056h2JkaVGYniph9
PmmRbkVZlaKQU3QP6BLGmYMcrmfd0WRxM58q2Q5CzCA2/yctjbfZLhlAg3LnaSayAobG7YwYSKpe
4qLmw8zL40+645jwh4Xj9W0tiw3fGLRx8HKrPhBTVQ/iYqdD3m95kPTnpkq+jNEbr1MONBE3Mxlh
7hbuYo8req2LnzKAWlmfyMqD1kws9dYmmFtK4kzCLB6Sq8z0KbfsH4WlZcTWzOsG2kt/YTFCKyVH
RlDq39myBiGrtBpUFPenA1fesll/8FjYeI7ds0kjxNWBU67h0dIUIB3/absn/KnkLx5Xauvr/0JA
xd87F214oaxvSwBp7xhyt6NOqxMOVAm+vEwXNZzcErLJr564cyjuoGAyMVFJ8z0bL8WvRQx9Hx5k
0CJ9QfRuKe9bt0uOXh/JYpoauhU7RlVZcoqlSCzWKITSrzYVEfrLhcVNNxQ9PXbdnlvVnD3+l07h
Gp81mMtap208p7Nzw+P2eXhKJkvkjiUoKB3yw/bqsRoYk2Dwh7rEYjxcOwRS+klHR5cOn+4HesJ2
pozqCPGrAbA87JTYx+is9bUbNOB6iSifU3vQZeDqEuZD7J0S2qGIctK+QAVsxMLpcdvYumkLdf6C
aslVY+bKnnMSb4nqgg6mZmV74TC9+Rt3yVE3t9vWbB89qdevNVfBSGUd+SQIHfRXh85dT0If8sS8
h95X4yO4OpbU1Ncc5dubQv4s5j0xLAAMR9H0aklsEH5LR+A8ugNM/TKth/MHWr4c3I7Hh8svFS8e
IACOyyPWYQ0hvdnPRs42/B5/6VQvKgdmLiNuKuQEglMOghmlzLZ8tL6Xdi080XKfFng9TXbMI0OL
r8Jf3g1oviQqyuvgslYb06dDRIzQjRN8JTrG6c3GvTu/WkHxgYgtAUBL46cZKLWEmkqvoEcvbcfC
6jyCSLYhszmyAiLehfRcXgNo1/NjGzLeJZIdy1AbHJ17EstazyvBqpl/tImjnogeUmI4wCZ3n5qt
HAlqBPAt74f1Rb5TgTgaq35bgVLVmSDg1zqSDpxvrg2GnEzicJtIsjR9bt1XGgG9Jy99eKII+Xcp
DFl0ewDcjrBKLeWlUlEY1ipP+0zPf5aH8f7ysrWiXuJt6Ei3mb3k4+Sxlo9KAI1Y+5NdZUT0LCSl
mNbRbGVv3cstDc2nFTAS54HBQga5+1eQaaQGJm+VjraqLC7dBt/E/7iG0ZehAKBvfyf4vWNgFU27
aihEP8XYg0pr6gMnZc9NwjM2o1i5ox9gz34Kox2aeV2xz28Nv77uZiKdcbLgHySlHSW2T11Ad8Jw
flmSxDzFW/kznm/N0mb7Bqm8t2dT2ekqz/2YsPNXJbdQMYXCDOfl9vdl4xOkxtawgcI4iE+W8rG7
KsS+YDdm+DTChcxxb0gS/HoVohj5b+eyoCRA8BpVmPTLtK/M9VtKrzELMQjxARsOnNZ7gdvVUYcJ
uSJqYgpuG4rd0lxH2zuoImHzsq0w7HTMT5v5bK6HNuO9P17Ju5lQRpJ6/JfIVkD+M2haR8B8nlai
8iznqgZvAHIQd1VdRIP2Ry2WmcAH2mX6IOg37qsl6+K96jcVxYIVo0yUbjBtt/1P3IfJHI3UXcod
35wYFIPe5OVTbXuydO41oJiDRHCA1I6PNwt1V1Xro0a/pvSG7ASiQBDr4b1r6qJyiwbmEX5gm0Tk
iOuuTsnASsSWWeQi6HD3knvl3a/ZDT3gKpTJ0j0HdMnqBZlrecyc4bZQL5tqyOS1wH55+PHeCcje
kH6XIYP66kJhWL/xtw+5vKxZbRqJJGUWBomog3LJERzGzP31xWnzVHg03BuAJrA/Kh95kL1hboWt
zKl49riUIUW5szYqbNIPqP6C6uomZIFIPaNeneBV+cPkiKEp6b2gBsPDvNMkl/bm4FrcOFnU5c7m
iwBLtoNV/QdxEsr8vb4HRM9bXRjgEmxeRCOK6Rap+Y+vf/hqWPth3rRYb37L7GvvEqLu1IFEIaH2
HJTUwimG/QUDELcMceeRZ2xCwKKmKAINsuhBYmCztqXXFqt4CmCXLiDht4GmsZnt3up9u3YYLLS9
AS+1sfJB/tdVpZBcVWod4G2fJcayJWIqHKWnyh5QWcvWXoVAAD4vth41ES3xnZ59LnwRW9ve+T6z
j6I4KheoXl8daqer/WakDBO1VtGY3B/ZBJXOrpyUKCv49AiZJ502tFIIpMz69Rpv2xDiMVx0EgX3
XK+Yq03JIdDNHd3fv4C1f0EzB5DvWPvwNy1J1lynl0P9sf4z8Y/BYRyCXCm8rD3GO7RgRUSHvKfz
Oa0ji2RLwykLg1CZfi2ELiOt/aHXiVLjXwIvOeBNQEZwM+hzeAKJpn8PGRX9AgDsp5rCbPUOkve+
3zcJIYOzcd6lceEruMsbtnv2A3CKfkFftOya/r9nKdZ2+ucr2OZ8u0mDgMZpF1MrrvSprY2WwRfK
W+RKhuz7euGLS+wkHqHGCc2Wnxm7IrePeArPfY0qk259MSZtTJ97ue/D+XpW2AwoGvDFFzi5ryEM
0TyHvFx1Y9xrzSfLNln6EqoNSnTJMFbBeG9ps7eZPDhUF0hAOGW7yUhGFU01nWEsBFazJFjhLERN
2xti1MR4/U0MxoFMfubpobXIpv0N7IEaWospafgnQUz8hpD3XfpSeuF9ZnS4zbQL4GAPm3vwBrIg
CRKXdsET7OUf29PzmxWbVxSgMxwPnRmKcWff0k4jOn+5439u2/n8WhJQu04ZXYmbuWbcMrep3L2l
CLmqG2dak6XhDYpiOzkezW0K8nDu66+/ndPsZuUBbEhlHWDl+PmydQPHUsMyDzuBE1Du30j+5cDt
ADQhuuCegYRILaQIXe4t3yMfn4Y5j4n160nZgciBKy6ABSpo3FWN618A6p60kG2hXeLqSv/zJLjJ
FpILKA36GfWl7d5mzN6HgrgUZOgWWEa9NbZ369ItCYOgE8Z0TPWv/FHkQMHjMVQf31gu+d2bLj0K
nL5lxI7tcjkdjiDOSAAWMid1nhrPsfa9wE9sH/dYYoYiiyOIxYjR6cmyAwDyDZ3Na/eD9mp/OTm0
5l8RyVN3zvhiAQCYlWYXxnCK3FljQjZRrr+qiFbJKjTR9XvOc2ihe18MxD43d3rJ2i/mXz3wFsNS
bByblbjObGyukiY5NwljruL4oRkYzquH294tS9lBfIwrS6O/LGQuyVx3kKoiXattKAFyG6wMez0s
W2L4Vf0kfQ5aOZ7WwaZsnfzrKlEWwPatufl56kWTVOg2gpq2D5Hg5jku+ifTEA7b5m9g8dxaL7na
TjeOzH5WzsWNfzEUqggfLYlSDInjtiiCO5ZLmpVXfdzgPVTpsuFe+5Koye0EZOZEWrK9WdkyQ68L
gOPj3JtWbRYZE4xzXGC5Z+lKzBDO/ZWCkFRXfdBurSZvo8NERW8trhO6D3iLJJ+c7DZWGZB/oFsL
3PjPPIL4gq5zZWGSWk5wR+Zjsl4WOWDu8uREOa9x5ophKRCH4zcXRihFPzhyOMOsuXrXHWiQdmZb
Er1XJVlkieIJ6xC2aFQ56b8k5Yjxxd7/EcSdBb6gvyNzp3cf/13i5GJFNnCftDox/spqyneCHAlM
5b546ylHYCGdcCIaeQMOlp74wW2FxnJwCSqaqWsZ9VwoDOxscvAoU+zP+gQreEP6MYn90+r4ytUk
dHsIbt/OLogJ8eSF/ABbb++X/UYwk4IJDNqwWubAbOXU0vOKWWrk6l5G9/pX/x7vsykAFOUEbULP
jZKrtm2zaGc0iCD0JLQC1OGl+TtkGn25SoJ9CKRe/Z/Z+7Jlxyea7lHXUqkwJynK8Uck8+cmT9a8
kNHppHDB0RqzvAEPZ9igXKdqTymD5wnF0/wLH5vRmIMgCEs7o15na1d7WfDgSgYrrRNRlte8lT3S
W62S1EuibrmpRbUTatklyMTkMH/I51yRe9ASzZOTsFyJjCWOxohIXLSzTQiQB7tCTpjays+N4gz6
+RTNA5ISrzXF7WEGsTHqdi22Nvz9bT4UHwPwWzoI7Nfb3jrCpt64eX0teMNueDLll9n9w0LX/IHT
kZvO68tXRlUpDv8s5NcQjWfPY9XBfIQzZ/KG8WH7+FYzW7Yi2KpdtQTQtvoZVYF92yjidM/yLru4
30VF04whPK7RzH+Ib8eJA2Xgs7iU/s34/u5/ciIgcR5KT4jrWwGRtsz1G4iFACqLXPzNAZuS1CqB
PpXPawXznWV/RzDlkKIwcO9D2sqb0vQz9OR/3HgponSBTugPL9U1i2qTtr2zHtCYBW0573PZVHY6
t4yxBllKpium4fw4t4o+asdbCWW1FczSILHcMQvmkZRjHGvRTlDYWCk0GuunoF04syUmdui21k9l
l30psUeXXAMVMsYzF67WIMy6MB4QHsthpzkgCuzKePtiFWPTKItxodGDx5MgXZHyGyoCqfOEEC4C
Xe1oF94F2TOarSYeCfzUQK/gtVw1oWqxAqXWMr/vVxTzqZj5LIlguPJd3edqCXTOKK3hZL3edPmg
T7tlVwThVWIKg9c/j9eUDJfY19tWvmetdCr5YcNCgu548mTNrhrVMMRgkqD17npd/tb90/7kYeR1
HjTbunDoytbcvwvg7n8hy3l91AgVfv3iBbl7MgBr6zmVdyvahsqcaoSK3O+p/2zm4+Oa/G+YMlYh
vMcQvP+ZfjcviFrZbZ36yU2KsBnw8fxFYOyjyum+R4SshNh/YEAw2SQ7S5oVX1P4Ez8NmlEVHnaw
TtRzT7TqAJUdJiPRrwupFe+I2G45cYlQlanODh8Zg4iS9EkH7h1WfzrEgnOuzybwJvVR5La3psw6
qBHAQuQkYlzig0jHT/jKRCtUM+xHYEbG4K1qEF7dH18XzJVx4T1B41gGqDT7sWIbDMwcmUAClUEx
D3EZ8ts6XN1mCqvGm2t5n+NL5+nKGAuloPMa/RsDvI79f/fwDw8k6CfN5JfMRQHz25oZ8YDM9KXr
ZefvhmK8ApOA4A16fta9j4mYAEYDaLArEx+5TJTOiwlqhtOQWFfZ6fszz3bhPrtltV1SwvgjPhJF
5BfApTzkI5hg52YpbHfUKNVaYaMIfOkBEEJd4npz0cFr4nVDK6BKYXEg8Rj2gL5OAlXetxr3dwVx
83dcoKsHACXu7qZk+tGnYtG/G/EFJWU+DozONNoInoTu+FSmUVQktUYwMWcvvQZaMcPPplNK9YQy
46SQLZJuXzWqxCrYVXeVk6uaQsvjVbnf2Gy81KTFP+BGIh+KsaYJ/yKI4n5Nd/4luv08D5kDkY1I
ij0h9bmC9aKOc55OBv3Ri18yF5SY4f3oyiMwfGL11/N5LOtcPEbslfFK4DUEHz1WOqbEd+ToY22q
PExf8vXqI9hP4+NRBSPX1MuiN7ADTwFEw/2PcdaHbaO9BkluAiQlHfhRExlV6ubuAPINUxxmbO1R
vLKvPH9CVgMvh5i/SGuZSBRfuS7ewoTM2Lj54mzwpS2azp4w5k6fK6LyFjoOMoU3ib18Z4RxYRLx
pmasGkgeB8bkat22gvw4+rsrUsy2zCICWhcjMILTnEDqCcM8ZxGpjsXY4Vz3+0cBGmcZLR+coube
Q2M5x9jl6Qzv5bTxtQkE8EjjGc0U0NWFHLuAKphnVlrnKM4cfcPcavAapKHR0KTBoY3lb/PKaFc9
doKRYUcrntENXeKDLEzgmPCxvRgM0B5p4cyydMV7vGh3qKsTG/G1L3Snv27mcLQvyltcTsHL9klz
9yZvOY2WbNFyPkUMTdnJ2lYpBiafLIyY1hX3qEfNnnhyPYgl1Vxlpt3uB2qKQ1SrjfQbIST/GZJZ
qtTx4uBW6do4DCxKP9NlK/cwKErn4ETkIJVY7PMBBnV12y4JpGI6ocy9T2NMSMuiMdnEA5RWV2ls
SDHrXnG0MFmrn607wfaiOro99UTL8CGh57scYHraJWy8Cu1oZpci5zAEBa7Ng5+z7f0ubOXmI5ZN
S8+81g+sjf+1qpObo3AZWriBCqGUXqk0urhNoiaYwEM8LExAS/C0oxbD9U0q4NXtr16bvPAIS6W5
W4KCIjH61TiySxP3FyWxtlRZv913EMgTXzfRRoeilye9V1zkSdh/qWKTeI+acJ8ZR/g3euHBw6Xr
d/A3Blwby2YfcznKHXzTvbyS9NTTzPy9J0vn8ml5wSj5pWs862CFbYRFaONDK7XYxXLavJC/t78V
1ze16OPmM+vk+849oHIXZguMKHtzlLx0UAA4A75VxS/73n7Y25O8WlI5cPIdiOQpElaLBGvay7w8
lDQaQtqoiG88bZwJp2y80RdPDUalJeJb7x6C/6Nzfz3DHqKTY0CE/+CMeqw+OA/o6LIZsVdILFNa
3o8XVg8U/ka59B9+qFl6URRJpIUwBxsR18DQMxD9RgGm1BhPBtGxDW/1+dFOTTNUwFm/GSGLDxFn
+tfbtajJ6z5KVhiUubrEA476ExNRMe5Z4zS6ORhCJsp3A40ij26fofPeJiM6ql679/K3mYTG5Nke
bFyZV1jFatQEqjKLEJIKuvdsdlaVk0tuQholXOmDg2MipK4hhngO7shE5J7vvnm0lD8TeXH07YU4
9u3F+KI+Cxvhd7Z5lDgjahJJqAjWw3zxyWqw7r3g4CEuXH7ba2lfFQr0DXLgMWcQxRtMelHzUcBB
BC1+GwI6xi+BxS5e6CHgIZyOHl+AEjHeBQg555NPbX/fogM9SScNWr52/RlobZ/HSPu1hyHntW4l
1KIcA6pv6dII9/DSTigyLwuW1Se6cZ/qS46nh6lPjmiVJ6085cC47K9nWboaz8z+2L7wvhllCWH5
Qq7hK+kxxlRjtUhr8sA8OHNENhrJuSLiPYcguQrzxyPVRwvEDD9IvBYh5aUzhhI1PMBxPK7CHgvw
RFwiWcSUQtEYraMVJqHYKbH/pLftKmOomWwSEvy0q4rUPC6Fwk3ihobAvHD7v4FY27m1Gh1okxGS
/TlR3ko5FiZEBQ6jTXvMbaQd/h/L/XxbceaDg+WodGrnTGIKFVh0PVw/QPa0Vklx5ECYrRm6Cx1o
ygTgVW7AyqLLdpNRAhRkKQXCHDetjQVhDdARzqswGfKoRqndN0OkBBqmlHRr+avZsorYcJRFcSNw
dwicmv+p7x1I7/CJIcb0CeD5UMoLpjl7Y0Xa88XTEBZKELv5KMJ2jt+uc4qNnP8Q0RlZnWmd13Du
iNk6gGKaxYb6zwQBqSqRP5+G6xyqDUg2Z3iqYB9sDssZDNgpQQlTqJGDykAc77A8vkRFZPf42WUY
RC3YUHLGuMWpGsbXU4Gal6buKARHKcJtGbM3/HQ21DerqTlRmqGvAY559CRSVAzmZlOjlVZr/cdI
ns0nzPGvXUG9b4RK2oHaFNF1n2ErKQhwJPzkZIeLTRtjo2nVlo88CCQCnHzk0AHYr/K5ByW2UNma
DvE5P6sYB+tV4cCw079PHRUAQVEv55FbjotMh8PL9ztPph+F/AnMt6Mh3NVwFN6WtkzjG8EY4Lmq
mjBbrFbxGpwphuht6BNtkaddTn4w1Qp2DbJ568IeOKv9vZeAQ7fWsZAJIVPPtmM+1ic3Pf0lcnhp
yatsGFVjGuLQ/PUOSqfsJ91Ef0ANa9BrTqK0Pf+ufTBjkc73fmPlOEgymI13X3v8ktVpMN/dl3qY
hcYhsKoatIapd/90srH7srurOS1lIRx2wGkbVF/2c+fGIwhwGUnD0LysfScf2UbKuMIMgX911pnA
zhkYrb2wsRWBTYSkJwXM228se4AmwyngSuR941ZoHRIuJvMPyL4XYTvqUIA/N5+C2cAIxXtEVdEa
91yokrGc+E0xLXsODoYTtokYCWzasuoNXX8npxSd4bKZur+AjHYAwDTYoqGEAah1cGRFtFnctMCU
Koq+rOKwhYyZiURGwe5gwqKCQJMU70TWMXqHOlesjojCDAEZ1ZMybxkY1gUB8NRs93BRSyvganwf
i80tzpQ9gnB33PnxISq1vM1TtKyyIcq2Cav+zFWDioE9VW8JO65AxG9dr6NVgrUtn3zuCvt/aMYS
EL25wYx2eIJX2aPLUOm6gtpOGSkHyi4Nv7vaz8jMK2UEQ0rNtXEW+giSnwwgZqofuKJQg6ZH5S7t
cMBCjNCtVk0rR4vg3slP1C66A+IidkAuSX66IykWrP0uv2sWbwgsO1lsnzjByd4JjgqcgqcIiysm
bxtR49V5r88zS7tBqMHqboJKGlGbk9Q+R3oFkHOipryKDGQDjBIc55LYTRYvrHXRkbBjtAIgKxBb
g7LNgpYT2+FZIyI8nadv+8xyKRv8gLs6hm1E71x82Q+anFxANqEfP/upx5m7d5Fzdv2Xli9kLsBC
Sv/SFnkUaGEyi8Zx/mHmR11AIfg2uT5P/r2JnnSIhyol97A9LIouAWdEUAdONvYOrX4npEw2PRe4
gWZtN514C9WNsVczsYpV5UkwCwxCuGUqNzVLw8m1vM7c9iN2pAUrgPmsjZgiYA14TtPWamCEbyny
cycC8gbqTwh8N+jo/zZoNdNLde/rwLVZDUqCt9YpH94aZVO3TCwcdCflL/uUcUkcSJ6hFIGfP/TE
5wX6t3o3jrIUtnl/kXbIk7rxuqiw7hxo00vYnGIMfE9z0p0u6SD/xtCe99IEQ/cggtO5jGFRXQEJ
1Hv524NXpNTYhWVyU1Lc4JEt/yIvb/v28CMdoxl50fnGhtKKlOkT15a68vzBi2pUu0TMH+/aY1UY
PcdmEec5cSwxom4Ij9Q7l3SOg+AaLdbV1VL8wowJWigANTHKV9vBIh2XWU9i08dLvK9bZghfr88S
vvTREquANyZRTFJk6h2cOgP0+7h4X0UDn3cudq41ngs46kvHtGGDxY3gWFdor6dh5Nw6TikGPn/B
k3gUbaD94cEDy73aOAYAFXm73IZC4ZIzkQPD1Qczhi+V3gi9UXevYI3FF4pxUNucn0v3cV126VQh
QBaoZeU0gAMPZCQ4QBgERkQ4r3neBb27CLOPtc+JX3Pm3vWDR5zMbVo8Vq03dGjKisOfRPoGGlDQ
fFXcqhvXdSVDync75DUjAVhApvO4Sc71Q1x4MrDE/nZII8ekY3U2sGmvzPUQKxknGQgl/pXiZax+
GoqvSSSWpxMwS+iJuGdhOJLwJoYS/ci2Msgk0zO0FRskuLt9d2PMNSGKR4DOgGPttIdlnhVmoJFJ
JWn5OARDY+LQtzYElKxfy7nbAbquNa/E/5Be3uH4r3w3rbirov7kycCn5dxguoVlL/kFJz2L9REh
2GwHTihT4V25yhAxMYww10oUhCzk4tajI2Jk4p2IrhyMOpZJxfSfO8ssx5sic55AHJUSLV3iUxoJ
lx4de8CMsp7AiUvYshxkFVDgzgTjZJLgRpTC+B2TU0qLjEzq1ecvKkScHjNUEL1vEbUEBLR+Ahrs
i+4FMRd2Uhn7n9CgoJIw1jTfctLreAcbLH2XtLw8zPisgqQS2iQ/kKLAhWAEJPfraCEnQ018zX8U
J3UJ8xszOXOGXZ6KQkNm7OI10+AfHJOOATkwyxEfPPrs2fba4iuozFb22I8RwxF6e/Pc+Aw+09Xd
X1PfryuFx1iYZek/FYeLKjfCuaanOoUfI3WgLEKXbYNVonZgEzBDtVhqyavcDiY5ovfb43otRWuK
O7jQgRhs1NIewdX1XT8wDTOmgquge36qFAU1hslBx0LAnLc25E9Z6D8Y/1C2hNL9WnofkhjoEoOx
EZKlvml/sZzKOyA8EkC5+DNg2sZVen7aP7z7ddhQRNHVwJ1+4Gp5n+hNTIJYuR5Fbm73jf3poGVu
L32NPCBtIaXI2oBVc3Ac1aDsK8+aJNhml/VmuynFaUTnPA+5WtfnlMO9J8cFZwB1ehU4fs/8m5vi
tk0Wq6L3roVzdAi1p+DXqPK0mA6PBTHsFjh4pObepAKIWB6idyCKN9uPXOHLznJ+//RqXYW2Ab8q
o23hfQKEyu6YXTrtytoUbllcUFrWWMsFKiQsXSOOQJ6k2SHcyCCl+S/XWyiaarcMNPR24gynj0a8
ga8zL1t/QqhC+uxXOcxhfIQL5BUhR2+dpL7XXRfXDmSvs5ZO1ADA7I2W9xPIODFco94NwI4YVmz8
IcEDOuz9+vmXtV8TSZB96W37dCL/BhTBCoxfIpQbj+aUQBs/bcEj6Iiqdwk6kcHyO6UC0YELMsJ7
molwIo+/C1/3EN7VU4sVERNhz9C2d5HU/G7t3nBtzeetyOLpWhJqRZmiP0lT5zN8NuA2jaIdtyeF
cRfMCRRKQeelBaJ8Z2yS1uXAgcc2RqvMd8NwV/lAdU3FAXDOE2NP9z97QyHgLhWdUEryNH/8ifa9
juxvIYNpVpvN+pf7lVXekFl3Ryr/gma4pFZFEuzxO5DV/utsuheUzaSFLj5TVaGq9XXtigfJtxkV
sYyIzyxmNgh9i1X0FoFkarwXogd0PlluFNMx+kycGJgbRJ10FpYM2bt0IvwaNeuAG7KF4ZTJNxV8
sD6KAQVcOZB2zDSCdYgE7rPq9zLKIHpmW+MC5gUjdvtR5cLaeV0nN0JMq3RiyJ0loqJV5w6DEke9
c2EEpSi30c/P8b4MDIytp5t8G5t32xZrmDbHSLwximdGXuqY0L9OhC3ZLypMqy5ChHIcMG0IEJoF
F7uFhDxhM9DMI9czoexRNmZLaFg+zllIxBL0wEtVCXYvxx9f7M0KZVHFrARWEntWgVv2ggTfPRKU
2M+CcovcpYiLYs6CIFusLJkgRbMQVcqn5wM6torlrs2OIwiEC9Cec/P+bhI3qOQjiPjUANq0MSAr
eGk3c7nHsdNH8HwJFW+aOWxKkZr+ftZGJs4jWnucdnJe3l7O11qpxwS8doQblDP1WBdOVydnotJ3
qeM3QFuvP+U5ui0lVD5ftGNbSDA6tXvtsMxFDvTVRTtazp+K4vSUBdVW2e7sh+vigDWuhigyXs+2
7dEajTpXkTrp3jzEX3b20nE7h6/QhvWX0HKXhEJCigK8meGP9HfdoMiuHl7y00BE6UXBu67unlID
DWqO+fgkZD1C5khx+9LzAxJssh3HVssZm+yqajAdglhb7Yf0z2uDXNB2FAPiBAa+8Ex1gg/JKQ4f
gwACtXCkc6TgFKbKIH5jdvLwaf6eyvIj2XTYr2/2ymDfOR6SmfsQGN2UAMHSmJWT5SwQr9KIUxud
6guvlL5v1J0X+yJvuYy9we75aAZNjgjWvV1B4usRoO/iKGdl/LMP4WM2gX2XfDQ0k9xTKht0Wf4D
o3Hc5764HQxXXU9JZ4dFetiSay58xruA+HnxtSW3xTHzs2Q1DKtWP1wqHmBxwZ4PCjgWBaDgWmyD
WLwGifZKGSz0YvmiVA5eAtiYOD9++IkCOEY48rGkhbsk3mD44inusv0YilIA4YvV0DFq4MBqNL15
0SezDPwF8DEf9HjcA1dVp4zvxcm6Znu+SF2/tyibwdqMBJCFH9+nSjrl1M1VV1x9Otdt/cnmppmB
CXmNMNQq7stjNf6pxn9cbKR0p69LYi9VBBtveTOVqppc0g3/CaUDYtJ/jeL539G83O9z0j5aY3X7
zmbW8vO7YJC62JtUCaq1i6nYN3hsvSepOUG80N5Q9xOK8Stmu6Nejy6aXfLmo4vDDeln3jyegZ2i
3tPZ+LF9awhQ4hHWH2gCy8zQ6ALdrnvkzCuYbFtYpRi2fp8tlR0xfyg8MAibzTBvkPIplhji8Nrs
pwdplm6wD9GRqUX0FZN8UvBrhTKReSGextQdEcwmfzMdGX6xh4RYxWKyY0veYSv+mzmG4B0Isz3Z
M40SgN21sSSxh0CdtXHllAVfzEPtdAXQON3cwRqEmKlVAICc9busZVCvtEeApTu9yDEF+aib5j8k
I0378Ob5rC6kflBmn/tZQGpGNubNB+bh9A+qbU5EZjK0CnA7Py/nMA6GyutOJeqDIaIbZ2Mn+S33
qY6C4PE3gcABqIsbOEs62oGtRkfCc6Orh0ZS092j3qPKaNjGdPc234Y5vWtOw1zXqBx3HBl52gZ0
uJSsMyuLpGKYxIIw/6ryCOB+MwcaAMwckKeikUCtgQN//G3lK610oWlwTEhfJNuXTQ6/8KsVgzr/
/9abCscAQzScye4U/jBw/BPXogdTjHdDxA5gZVDmHKBmGmya2UFffatx9riLsG4Of+nUwNyV+70Z
tp6ue3eGFxtPve/FH690liYot/WdBE2PrepWnwTXzVPAoDNRk8w+MK4xA6tPRUqJqXZs6n7McML0
xpP+vKb/kG7zi/B5BUcOt3aBMYky/8SJ1OEvLytMPnEz+iBVAPaFwW0ZG+KB36Ikl240wAiybnmJ
2eKrZBAzZwJlVonP0xtsj7dzOlclvfUO1DpD7NcDBAqVpq7suTyJ9QwtD2Hl5yrfumqbhDW+8YZb
s1FA0yHu3ie/QWg4RQlrU/tlcWr7TS+noNTbI+r0rnGpGA/Ey5VlgJ0x3LTZFkTX/2N48WJOgPRn
y6jSpWCDH5pRq/OegnaOXmxnCfnAVCytNukHOAJVq/9QKiom0vHQSw8ZonSlAuD23H/sJbtt5te5
aKAztiwkVMr94cHW/ovffVrly6NM4LVuD41s2VYpUo2mtvhfj3PmzY+eD4FhOJxDSR2b8qw4q30U
O8nTU+qCYRx4J+jnowhplmS9oIiR/K5La+bOchkgT0Gvm8fBnXZNc2m0Btt188dtcOJ83iVviLvn
UsbLk12ypE+/aMgPFt/d+l2SQW60PW9QBG5XSr6mVNgXpQqOBmy+Mh2StRbkYFBz0VcDRKYsZRVw
Glym84DgrQ5tlqS0ZeVHY+0TEFpM+rxeXR4JHD8I9dIp0BdmGc72G6YOSr7LJpT0onYtxatApc9I
XQKCuPNE4KVdIne+Ge/7OCmGY9P9583j8z/Oy5DaezeQ/hjabpThMGre7hDImieTPbKT511go83u
4XoF+zLJUSauFnB3qzZuq9q5pBMrlH5l7CJfSKawLRbmE4QUo4pcO+KKJPff2Xeu669zfcSDqTxe
Y2twaxHywkE/Cr9NivDnny89h8JpS9c9ArfskrZSUeHSAjHRSVVtut+MrCm4D9e95LZMAtlqfidL
3QG4ReQhKsMISzhvMr39X6DKydmuK6OPIOYjaWqL3mwxrVszlQ0mGc4r7m3hJSpvpTuTkO+gQ8gl
7yA57DSbjnG8qgW6RVqseqSv1fc9M5woBIEhtqX5WuVFRpaycIR/EQ1PFVrI5hatejAQhP3lP+AZ
GWfiNQkgSFz4MAz/Oz5quhROr7VEaEMb48nq2J9eCaORkEgjdx0tWOFiO4nu8Y4fFPj2y1uTHKuz
wmZ1cjEH1R6QPtwT8dlCbd73O2oyp5yzOHOXTq0l5SOsv21HzjeNxE/Q8mt0stxCqsZEM5i7kQSa
2MehVhlhgZH/gQiVGaMDiIGs5vleQ8AIx90mEEsG6EvDIE4XN3VZEMlMP6dkK+k+3Mfavs7PdncQ
iQBGZO8C1ECgfuQ3waE4zcqNNYxkCalvn5sz3d+6+bXS9j3AZKHKrNs8hpOsLTnAPcn4N6ItPJNh
vNjsZrSTHZBRWahzD1hWAlPVAmYpYd46kvOTs3PmCzlnABdcbGCYxXW4ItoizxrnWi/c1XLzq6KG
g6/Qf5kmNm4PU4ulay3kD/EpUlh9V5zlbT9jbHGetQXooUGNMZSb2U0od86e80Iqjt6bYiuKdu3e
PJuxzN0rjMP+kyW/UK91/1w85CoTn7GVC7Qx+EJFt5SCtN6gurAb/4JQa/7lb9LXtlcroK9Pp9fX
TtXlFWy/CeNOFUIEciox9QC7WDZ8niIDWkNhqt3E6tEJLSsAIEPt3fI6WQxfGxudYQ8WtoCuRKKY
Milu56nU3wZwExhBEbk1mf6gxZeIyhwPxfWT3Ad768YlH45/4PcLXaXDLF/ENYmrCTiLcf8lKnhx
kIp54RgXeeLCF7XWTeWBWjlPJ8Wb3XILl3JjYw4lJo2wQJnHHhH3scysgpDIEaTkAERU5Xnqv8y8
Wsjh6FZUjHhw3NPvrX9qujgy50kO78CCW1mNIBWF3sHarALjsrAQUG6y/O508RDKoCtDORGsVXYy
vmTi1DfoIogI+1Swu48+LF7Jq4e1Zi/w+rsT4rjGa8fVUsbKRGBOuRJS2bxn9YJnjO3wRXMSRxYi
lvxsUFefmjO4wGy0BsjZjdBDkZ0hfPw0D7HSqxOQaM/0MJfInBZoL3CqEx7NzQM3diJHaNdshesq
elzzpu0Tt89ifNowYDOJGrsM4rfioG4hqHdO21kNOvL09BF+R3kEhE3cvSpJGBwh+4e2LmYQC6Ep
pzwNNpn022lBT3bok8iGaJ7x17x/cHU39x6NVCWLef1pWgMPqTIjOX+gLKxEgwRlAqBdgvxuMV4N
5WGMEaiXf7DwYXseo37UfnD9uS0uMtroTtsKGhzH6wkfT83TpRof10UPlSD4icdd4BCexwA4bzcj
wgweXdxwSHAxwbWwXrsoB9yv514sAVOdYECuo8Zm0H3UbEVFZZHPGHatriwJqFlgAk11vAic1J/A
yHQUtyIEqYh5KixTKVPouIadnOIDP5B0ulDGU9v1xcq0qfQNC+2/HCk3LEZePnOKPpajzCP2aH5/
R+n4Nox80sGlsxb8BgkLyk0MRdj5wRYj9hCN17WXhX6YY37kc+xxDzv2g05LWC8KsULyTmjxgk90
bd36CU2WoaODotAxl2tthmxp/ZRH7LQoXLHa/llpk1E9OTCF4lC7kreRXToP8T3e4sP7YGr8Uc56
J35/auevn16Z/+qNh3Zl/1Gu78RNU15qZ76YAiT09bKxP7Oa8154dDKKi6Z7UO88MrcZytbsXmR3
kf3LwaNnPmsVNA/M/Ww7pPUCcnNjAJOQ4NhTjZy0SFsvzIwgT+t2ClUTH2yAlwLIJGKOkWZjiQM/
xowPog6GEWsOgEkgHn/qwN48wOUa+7SG9q49qOiEUAd5sEoo+1jc67SN1jlgx79l2V/y+O/+GgA7
pYNUhJuj0R4k4JwXYC+YQSII0GfwSIcfqSILFdsJPG6r4cijPzB0uO6gHM2+TevKAanVGlg4cXnw
H12PAxxp1kJPKyebw8daMUe7/i5JB5jC/vNj4Kew+swCbE9b8c7moJhywNqlzcoM8dmuTC7DWFvp
RsLunjQdmOZDJ2ByfRX4QGHSEk/S/GS5U0IV+uoulbxCBe4ewRFKYatUbV8BNbduATK+XiPsQzk1
9WYbh2gToA+8G1iIQ0MzdgvpzXyQbrzhIOjno3AbjgXSQ9uPHIMExatOwCejG4bG/OhPglDhgcaV
GxYMG81nzLQQNvkvOa2DcTlRu6JjAYPx4LRBQQKn4kyms9SackNV45JFESRBPlKDAnxWJesfHdnR
TCj0jQarfFcGDTCEU4Ujbzlpjjjx/lP4hFdia2HcSvo3KbivBtUi/6IjpwikdKE2Sx1DNxm3Abvp
bT5PY+wmH85AepBUVIt8D3COxg+80kB9T1fgg5wQV4j/J59ntziT+lVNs5gnsy6R+1jTTHiLas1M
dC18r1LWb0LPUlI00F05t1VYloTzWo1O1/ilFYBZI3RNMFizxhlTO2bcf7LKOnX9JVYOtTwX/ZaR
n3IvUjQUVrb9+aJD4WrBpDxp4IWevR5Au4ftfWjp+ETejhz4cxaaThX0mLAUTGPReNZJBLj9QKyJ
Io60sQ6E4ahnYhvr3yTwyhjKPDPBlDmsXbeNOpC+nJJgUeC09SfxDaX8t4iqIgSk8ve4HFO4YCzL
N+J+jWFDYSo8VZCxtqqP4RldJ+vasusiWt/xsK50wiFm9OjUU6uWlrOXJQXO4c/LoRsuKg/qB3Vp
ieFltb2ND00bX8UBQrV3xLqkccsT4/KmnqpgQKQe5hrQQrZr6D458QrE7gWF0Wyul+CxKF0+AfhT
XAoh9r0W9ECq9kdbg1Wo+tH7oRdsHVvDTPNnOXbrUDt8lRap99JRxqFfd0DMEisBYIzc/XvahjHR
ei8q3msIeHmII9CV5+qWRj2svUlP9MEK9z23kMmKLk1kDva0TlZ5x8MX9xQUhaXl1hCkuwAE2LyF
mlY/QuxYyjfw1ezVbVMa+5fHO7SCylEBC/TJdjZ3KIiVoX/d9MD1CHBV40jfXhPtMxAa1k1ugqSF
ciKSvT/NiC7YxOiNA7MnHW9vhhHuz7Ir1M/JusHzIotCGnR0uN4Y65WN/vnhokh6G1OdMmt3q7l4
zAXcOtIh5RQJtIhqig2AU1SEizcecvwNj/tdAsdsyUiGIEe1VQ6W/ysW4K7CpC4GMyI/MwkuK2AN
RmoCQnGSCcr8j+umY+cf1llv5NuhjK0U5Rtr0fZyXQAQG97nHqUZitkKJFHlj7wWX08WHV3yoJxx
MKQxDYgSXro/QFzVvmcWRHHU0YzhSEB4WptYE+DbAgpE3IMKzm/KMyxvxEVACczsm9V+q3PT8Vj/
WlDtxvYxVhqFBaKP0jiQ/kiXixuNTvV+Yjop/bVM5/9VIk2NLmQPTZFAoTuo1o5+yMsm7kDFIf/+
8id7G0cB+3dd9cx2OfeT5Wxir2SoMEJfXfC8vVuaQWrIwiYJ5ckk/SvtLgpwDP26xsqCW6d8PfgJ
1YjPqRTV+2BeEPVwW9TXL9o66X6SbFW9w+LUcDY6uLbb+hMBObAbSwaJRKkB5c6GPlVQXe1eCIy+
7D4KAIJO7KzrcKemAXAD1zDiuzlbRIelWKYWc2B3o/LAtHuFr8FPK7ebMz/Xw5xp/cM2KMIG6Izs
eftUT0vABRgMGampL0TSdS2Sak6dOznqXUMe0lNdvBuyHxYRh8JAUlcpSTM/qzH4JgRbsaGWhH+w
hcpfGhuPeGQ2bIbsnNJOy8CGpTZvK3RYgs3NdYYePYuGVc5SL0EdHAF/emVkgAiJO4wZkuVnT46b
8IvhhIyM43qBO3VZjTCvoBRBd9g5LboFt+qawHStvCnpkdNiADXbzofBKcoZ+wE5NNwOWwufFMLN
qf61pbGHmLTurCHpUZAupUOVD1GkYSgX7GIX5ROuISetK7iITb6XWXhpqVJOXEod8e8ln05onMCN
u+8xJ9WSOMUtLwlyxHA3XF2bxwONAEZkXO6ZehYanhrEGJD1vhccN7mRiHusixSauApmPc653e7p
zEIMtxZOYsr2WVHCr+tKBEhpK5+cqH+Gqge2ikr1vTBVNrWA6pChV1aCUGSyItYza9DTM9iw5GqM
o+pcZBg14FvI90i9/RQOqyNFFcrKjiWKNSsUF1dTzqPirU0UyVE1qo2voXImhhd1Rsu9XYRRsZfu
o3uNUAx+MErJF/N8IXlBnEEabreJUtmFbcdvxm5v2Rn0lKBNzJ+xqiDMLHYwCSvJtoCPwxjVT71d
MJ0wsC6HJke2VWkpyJkkjgbf0jDKr29+zIVHKfeYy55ayu8p7rlk/jup4OAA0nlzTLTv/2AInVNH
QQ0XCVXQcObLzS1bd8Pm1XMDcKqp0i9Zpxr/+mij+Z5ozJuYl1vjVu3BlaxgCLT6EPGX1/JgPXoQ
qQbCrur9TzhaH+5sIPrTfaybgaxFYRCDp71/CJWCcW1JkXEBjmgbtAsu81uLnZUMf5ffXVHI51/v
iCttOY/rCdQ2VGt1lr5rI0Xp9qb4XC0BCo8u4JdGdw/L4vSesu4uovu5SyDVm9nkTJhzgcaAb2cu
yKbO+13v+0415gSQ8QLy/xCyNQa1zk2MOcdiIT3CCACzjLK/3/w7Y6zGhJCfowhUY/TGRQqSmgu4
/FVhn6cNYeRM2842QY4DfJDd8OCfUKSSA+ySDgjNuBEmgWh6GfzPqZUqfZb/7gb9DIAwAchISpC/
cK8mnXIi4D7iFjdqHEss6J4Za6Hfw5p4+mjqS2iJ7yRvSC+YonfyPD/gEcRdeuy0ADTIo06wZxj3
KN70nK8Rw4M8mWupjtJh72UWzUvJcli+l+SGSSTgxAmwAtP8ZmcRgLpMhvo7GBMMLEC0tklmM5uH
ssUfq9XdotGikclI388O6C/oERw0CjrWXgC5K4fVYp+jCbJUedXaEYaVgBHRR35eS9OJw5NcjhzV
q5C/hjEheGPog7BThDIIFHjlmok1vttt2y/EQ+5qHVMD+M9st2u3fiT4IErX0YN3MmmK34f/CFmH
uqTrhfBSVai7ESD1PwfQeXPVENQCO/lCd61OBj2cPh9dcLj1kzXvheNhKzw7cqgsGS6F/NE155jv
x45kkVI7igyE9W6sfRVL+rt/Wqw4FoCSdReq2LieTmOqB6hNaOQZEEW+V9iBAe+hAwOX5STRKgVo
JkGG5wyXDffQusqICjNcts3RNsVtk5yg5rXIkdZKYVIh0qmRwCtjbZ8p3eAernf5soezHr6Wavnf
Ldm9FnsxCPzAJ79eHosNkoOnQmms96jbDlkQdCAJdk7kCJA6UpdSdnMr/bZ3AIxxex1d3Txt43yH
FawwS5+wHPEDwe2Fodv2X60XVeeA8kLKcwGW+2bHpF8+93PBfOUT7WYwl98+7oZRED4346VGL22B
Ggmqm2x3q11vJ7CLfFZf/Z+l/aRrWi8vl35/+pbhqhaNsKmAYHSMGLMCNQoFSsSlKQscYwSFIAcG
WDPXr1ohJOhQ7ZqLN3c81ktXv2DFTGgctvTu/oo3Tw5wfPs9qeWVdvvVtxyd88VhXT2wWZLRMBDU
eEkXG3EvJ1r9S1EXH+r91aeCL1rn8zVK2a7A+fGRRSCjY77jf9J+6Ch2znWLhFpKjF3ZLQnzzJKg
4nZNJbYaxzkev2oXhHkut+AV1O5kHHHYbHEFfgDaC6HSNImBYZCPkgjLL3PDxapqaqJoDZnujLOz
ZFq+d06RGvxY8NWOY3nYEzYrhWX1w9yWmpcuKDXSoikbkYv/vfv5nmx6HUdjVFpfiMwZS+etrlvB
sURrIvNanUqROjTWq2cUJpPduLrHPafHhdD8/jUr2E2bOm/0Xa2ApIL24smEbI9n74AnMWyeVJJe
jhHjVjCFnnxdNIj7En6eDprYhslEJxjh221/mbm6lEtVA8fKajtvWo0x309SqWVkbpmbw9Bi74YT
GsUylCwvzg+U99+M1kyfRCbV/nNRB/4ao0JI6fI7Nrq7YV726TrakbCzDaWjat+wbK02NuJ0t8Fo
E/Pgj9DsHSnmjGegrlMFjG+ennyCmaVOo+JSDAuAqZlnyPn1KG8OsVeJMrpJGeDnuE+F6JxXJnze
lv5bWXhpvDw0SudMsploSNKCPIQC1YyAHSrdzVljfWl/jFtW89ZRCHo365pV9L21fwKG1JPB0plO
hvwLIjyDuNvkST1ZNt9QqTaTdhriiPNNN6fnHP7ko811+UxsSjkpK+GaL9HURH/3MhAfvm5jadg4
tyosr2zvD9yEC882VN0lc81lY1g8MgVECz/96ktuxUbFToTYK6NOJw3cx8cm2EaVSBE3FI38dpMC
w1oU12/isKg5LeTYK9P0Noq2TdX6OcuKgSWhSxcJpJ3XUZSJnYXAkjHAo+lYdiLV4U6Pbwbmd54l
K7D/HNrYfPXWuPNlcb+ZzPq5VfD05STS9HXNaxcqOm+UX7oZefWbdcX5aaet+h3L8xn7/UNoOfYO
mJgJv/X3RoPKan3dTbrtGxTmOfLCT+ChXcfvJUDC/preqYn7WDaSCgWsmk9uTdNPbKTjT3h/5prH
LhBAYdgsAKe71hLkZcakTcLPFDPzrH0+fMHrs2jnAwwTIFsdf4zpGVfjEBMWQ1N/UAPd/WgBqabu
dcKzU3cJORIdAhtNWVetccXvKtQFDYIxzsFnl44JHuIa2iRMFY509npd11wB6hOlfOsA47aZ0zpy
wmZpRi2qeu6ZI4L4c1oPbtYy6NSotdPOoS88fkqN1Xzf3gbo1MGOclQ9X0RbTn6Fh/suh2UtmFOj
T0tVEjsn4aGwaEexNKR/H/z41lJjQzaCNeOjSVcGyo31pVV9Rpkh0fmKiNIvgbfh14ukUVDoHs7V
E+PSl1tAO8Db1sq8BgbaA7WNEZbt+EGtyzdqsJIulnuh3sVdDDA1428Y7auC+mHVHSUoeiPkX2QT
/eCEzcms76VJSGMUn+saHg9KaKMsLEFnwJCbKl7xIRIEH3Fg+DyjWt98OUurHiyLKJiBIvR+T3Xc
4izjEe3MhsJuDvN3cufSziUrUOg7U7ygD7l9p6ggHCUGGQaZiu6rJ/ouFfhZKd8pdwZOnB8Nl/mo
QijOABGh1rAAWuJIu7gHKOioYscaSMYrzbSPou0RDjfFpl4INCqDqym+hSkqnwaDNs5o/412Kkgh
KaP1Vg5/pFD6EY9b65b6IwVTztY1z+bzjdVI3+2uApHLfGhOkJ2c9OXbSaI/hx27e+mb7cR64i5Y
crHFMlmI6bh7yyKG0Jl7Qzp0si66+2OVSJpf+cy1mZykQkPbXpaFnp+Wrv9BGV6IKz4v/nAhqR27
5AE2qVY9Xfa8dGD4ntx3Z6O5rt0oZiVyF2FI+3B4qO8r6qJNS6IeJg/MbMfPQ51qLDevaeYtRkO8
M0EiPvwthkHC4fB8hsHJQSlq94MHwUtNyTmMgu/KDLlC+zU7GY67Q9G/CFRY/M6mI1RuUBilmV58
feOD6TiaUflEq5ctYutreggKa6OIyaRHZ6lgyrYbkirS/18c7hZFxxfW4v+kPAgTBz0jN/DJiAiS
+cjf3u9MB6D6ftFlBLZBIAx1nov3OpJqgvR+DnsgwWAKIRB1Y5JMDMD78DUH6vCQF0C1k4S6y/UP
2QnmdTOmgwXJysxcTpW4Id5UbEf++/v+v6eaVmOmhxQqby30Y8mM8j82pbo3u8MxkE2oCaD/RAZr
3ynOYugSTVKd3bufUOqs+//xBWj1oNrfF28TMD+oIx8wXh11ip0WyE0IK00DNzl18RIcbDOfm5Td
+sMq0jMU5WIdxiEj8/zCKmTg7KXSzHBzA/rBrFd3wW+7LOYq00np4mki3j7ywjIRXkzat054ra7c
4BoWzIezU8Poo8lDdDIG58S0WbGDwprmaTxCRMx8ZYVsrwjjUGPYah0kdOZNI7sUNspEQNPq3r89
rBk57vq8Z9SDHjLruvGb6f20oyLAFCaBraOQ9eZaYlTZdVOIlVSTB+J5/D7Z42rPoaxQXIBmLGu4
gn5voSOiq23JN2WOufJiz/EF4n5ZAk5SVO394ZuHqkc2bGcTU/M+x/jtvlTPT5KxT2ZNSjrEZ7Ef
yQMKrbb4Y/XF1wtX28FDd1NlnoIMIJBB7LAXm1dStkqjxrdGWOZpzj3N/dNzcbZTOjYupl6HCXBg
en7Hx0Zf05+xhOdemrBBWB0bRyyLsh55DruGw64wk3EEcG6r/wM1gwDTqP7D5VRQiXPUz7Tv9I7/
fJpuMCW56NsAMFCDGK4zcQreDtViVCmw12PqyFGOlRoDVKqNuJcasR9vPz2N0HpfBk8FhHoJRINc
8EEIsCHxEt+OKP1jkOHltP1plEG3ppwA7VzimohV08IajX2QttaDb2zSBr4nlT8H4NCqUCdtpL/Q
gtee/ZwkqisucYAHngvNCGJbgqwB2NK8o8DzoxTnTBypR0Vz4OUulV4PNShvA+Cqn+RlThxqIFvI
3htQD9LALeuZDDgT7ZkUKcl9CsQujfiCjN2EYNrCbZWv950L/qt50YN64XEkhu9rVyzRptLeRm1S
+WJh5eLLAYbAm4a0Vnr295o1rRvuF3Rkf8V8WAma1j9nEyJlupx7IotzKEbBM7uAqB1YvMKrL+2W
zQwv0ucDTBO6RYuVjRZklt8nRgxIzPRGdYFUCPp6hfgPgpS6QVkdyQY+zuILhz79toJ6hxjM4SdZ
G85kHdi0C7qQoKRIkdZ//Gliq7JgL+1FedjYRHy2acbVKX2WaAQq1OR2uHl66h3wmI1B9Jq6cbvO
vYzMpIZLzzSwhIyKy+Fhj6d6jzCavv+Pk2batWo93rwrKXERoLdZSFYV8yQ74NilRF51YDv2f58q
xjHU45lcdGJpRI7nWArPlG0l9ydLLAv2vP/aYh3fdcTkpVqqDMd39+qSdceghQ3Go5ndH1lFXKqZ
g1QwwFWUI1mvzK33MB91nT7wlvIE8Ka7y4fSzqCRcxa/cNY8U+s8UI/RNw1MYu3JxPG+vOOA6cNa
OPGbFQqOW2WuD5p4myEDZL0mg2UY6WkAbYJ4nLUov+hQSqPGKLj+ojKew/RUYitzPpzZw3Mf3ncm
7Bm4B2sgAvUoyvKMegtllP2FaT6LQEL4ETn2JjwX5mE2L89Dal1xo5dp7Pf+f6r23/RSXJmIp3DB
4oWA8g3rA/s+Fc3Q7f0Ww1kLIuZVG0H2bE0dmlXNLSWuMIhRe2gkBcEV5gTpLPTyXPyl32tTSdwZ
yVbUsVPVJekFv8N3EqPLgvaEQQpJBC8j+hXycI2c3Lm8jGkSMeR/C4kVI4HlGuFQQFwELXCVVrr2
xJAoF04KX9OhoJKuaYxnm6U5zpAnDaTKeuX1dqO2xKofp0gujweeLu/uL4QVfewxOEovNLxYHAvQ
Mt5s3SrI26oF/wPAEh/bIXfIM3d91QzWmyTFQGd49JTWGVKri7FY8hbxhJF45olD3xWPOs3enFDp
cWsT3LkIiTTj6IY5Pfn/9sYwLv+9EjNoZ6OOvV9iE6waUIdYhaErPVmSDvDGCZFyi6Kj5CGk6Siu
P91liiCSQYH7m4kPbjgPe3U/SMI9vQvoR1Yao0qyB5hq6hVGmFIi8WyUOS8CYC9VylG3KSv1+Lq8
z3x9KOhMOSzWjCUKBJqWcmwIRQZi+BY1SK1zwnQrmp6vFXegpWM43kXqoXCG0Gk/l6Wun/3k2G+T
fYleNW+PlDuT3v21AiwJOo2eX0/pWRY+LLjL32kjugENjTATvnkIVmKfSl/Pq90f2YMydFU4voKs
zy59LsUuVCexVuv2KAn9ue7+Hi5cRg90uc8cJ2GRpIspwHyb0g3X59DlKavXZjoZJFmqpwqTEmEV
gOv0nG6JcK8GAj0Aw8Z88uCIP+lIRXRwYo/CRvzCqguOfAROQuZLgb6GebKBOnmFr6HFTkI0H/TC
8Tq4J1hc1LLAVWzQt7VBHpHP9YobZgDV5PmClKPLfOAs7j+BkWG4f9c17SmNLPkuLritG6HyioFc
SGgEgbBDbOUrS+RN6naq6DUNfMDQ6RUb/R3LPleHrrr/1qT929Z7V7PMV4VPGBWwGnW/IxKGBzsO
lYP3A7O8ZwvOYVV4LgZY7EnK/KG7FJFJK7+Dgi8sHzlyyVuuP8vozbYunfKiL9c871SSadicULbV
ZvFFcJ2eR7H6VPKYbC/kDN4TVGMZ3jTgJVcfpvJpaZ40wy+u1hdCEvc6gNc9TNVWJYAQZ3L/WnaD
7C4FXUvm/sey7ASbWdNHSq5I1CftQ2U+7icEh3rUiMwIwbW0jtQumTnvdFHw6AAQZDofC06eTCc7
fRcGABPTU//uzkb0TxEVx1oJEwa/is779oVQ9zoiRLym629i746oM9NgA3yujzHhtooQypRSKMaS
5Yejav+SkLC1FiTo04V2czy09T0f2//1J6HYTVLprqlmevhaDmEyrPe8d6vdOwhJP0cKpPzBQTnv
KRhF7ep8PGjhMY/NweuHeQzGxjC1BC8CSsXea6Ekv+GAyDEMjQ3tpJO/jL6+ZLgrnHpy8y5y9Tq3
FKn8evy6m3oA0uw6AAGjHpf44XJWcvT0aja/+ecb9YCwknHiGWrp1Jd581tKqkj9GodWZt7e4qyM
NU7/oLAz6a85l2eI+GVlak8NbOCRroPGep6lZbomcavAPgdIAprVlOQ05Wn0fMdQYFizG4u/ag69
sHO2tye8rEQT9LxTla1ua5BCgPcdkltneZ7iYZZPw9ryfFjw1TJ0DishzPPG80cNX3XeKkhY9hJq
Mpq1OniYCwuRDmepCfdaeCnWxkZSJAUtA4oQ9kgMS19uR8SErmaZefWBemNremM2Ln0mgB3Y45yi
Qkdbu0Ln0gSxM7edGfhZUAvqIkLlVAjRNd6BK/jmuqSGRuentRIDm9IpCfa7iHuLcq4raeTvhfds
O5B5/LXoepFQvOsRp+kXentyLfUf12jpiXWu4kbWg0ig/FY7OtnNJwyvC2O9KOOZZvKpvildqTUn
hyooJoMyRKGvBdhosJfh5srZzOwoPkgvmf2JrypkBQiuum5avikDwCc3fy1o6LJsNlZc3pEi9qr6
MI//dgpsgvage+GoIeYH3OBn83cR8I2HI8uoa9d+Zns2JdIY3qVgtwJawOWjjcuT3xbuEDFUGVeG
9CFAEAPZ7117OUd7mHbFgCdQCj62H7DGSKcDFA5j6TrkoTUKuqAHiOeVKj8oHxfv3BPbkXxUurKR
6ZsuqBGqx4awcFXUlNSc/f5egYc7dOfYob7/NRh2ZhaG7Su1v/Be9XrFSg8OxD1KGViwZgvtPo+u
I47lUifgcDx2E5LYZSYeui/lwPfpZ582DScnKRtgkMMy9dQ2l50N2PyES/80P7o9/ZVSlUu+AQfl
wQ+euqa5t9JwekDWa5GdU8n75/x1+n5h1xv49DKSqYAkGRVPZX+S+pFx+9M5xDva7G1KhqCx02vg
BkabKj12l2tpQpe4tuS9LYCDFeQVdrJsC6j1HYEPvLAHOi9Kux8ent9rYEBDPg7eBMYTgevHVqkL
4dX/V5ejqumAZD4Jc7y+62+tQOMjHqOlTXXZwhtBfdCgiKRy95LGbJ9jf28klMVunb22sDf792hL
m/9mf0JKhKWaJMFZ3G+xV2BORmjGS3J9Ydu3BZN6RQmbr9ZSF7oDIFPO3ldqHpgk/hcwm3tct11Y
pFli/BRdZF4epHvTO39lMuAdOzC5ElfrHjCeymNIlei3f5oEBcPXQsJ1NUJ+/wARi1nFqCsr2Qfj
fvzuMz+rXc6D6VLsOCFqlRBbnTccnoGOOBgr2xOiQD7yAUAcmcxzeeZ+aJv4jLfvfL8WMMqOJvnk
U0CK/sMcyvZ2lqCm/aeQEafgEzJwOBJTZYqss1u4ZwW7h0Z7EWuzvY4/lkB316HICICXQgI3/wJD
TFe/MEH+iCT5v+iAXa4FWii3vvlvsCDVtqjum3XUomybB232xkdsyqh91efjsDOYfj7KJXt/9cSs
zFrKDNZJZOjGDJCZbQKicBnSWI7qW3ChC6DC2xeK3Y5209JszEV/lsk1B7stcsSd2zOu5CVL76Pl
VR847iatPW5AiXW9qfyWYUJ7uc7vNls877YzP32IpJnYTzz6HQ5+PLxCduSas51xSzMxt+D8J45T
dqpwGpUX8eP+w+PrT1OlJn/aliclhICqqtve1xBh3kmhOfmhz6blSP6UsGh6m2KLxoLERTIJ61EI
4RnLtRqGDa5zt/hCbxp8xKypzZtaCw4VKbUImW/QYolr4cUzUd8aE74VMobhe4iClTuKh0tq/fzT
YBF/7rBMA/JUF5Y1wSa70qm1PrNuuhKp0ixIfhqm9r8v19zo4Ado+4NqWdtHbQnCoCBvouZOojpm
VnvqXoRhMjUYlMs6q4+QogN0h3edZ7He5qHQK4d8HmLiTMiWdhCNTLcjkHGOvjg3Y+qUWYe32pTL
jguJfCNU1FYhyTsVu2n0GKiwq6gB+bsmZl+zyTFqTC7G0EpgtlAJGr6QzerIFyTTjy43cE5VPJJf
Rwr9h1ab+gyKqoDcUd4Ig2xyAHVsu0/yGaOwkGBLERm9kr9H3T69qLPXbMM4mx3+73QDFV8Of040
Y5AcIIsm88/cRyyyS3uXiLHJ3BQ5h7L+c3avor/0mvS6ExkIGR0fi901NerRR+rKcU0jqx83bdDI
ObDp6xrXExXCH2vCyIQUKW1ODIq5kvZAg8COAxwjW43dsi3su/ERPzIfEMh+C/an+s5DFMJyvfpx
CJDHn3u3Xvcq4bZhI5NPT/KuxOhXz1vmT7dxQa/xcX/QbPIT78DTSciikQ0D24+il9C0UW8NHYj0
C0QRIdpUu1z3/s+N2xJLR9pUNAdhp+K14Rmi7+cmEq3NVTELt4hIG4fjv1FLzHGH6mBRcF5U+KxI
xM1zvFW1RSnF0wb21GnO3Q9NVBoWAhivglnSmrdQvNrgct9fii9ZyCY1VjXwcjdT3nLfqTN1NaCZ
cAQ5kaGuD4MIbxQ2gB9scS4MBLbptjbzNKUhpNwgdQiTlPdazmNEKlScaIQ8ZkwKd0852GLCWoFJ
FNpT8PaXF++OZW9tZqvN1++71AF6G1gpZFMN3pP/hp264tA+kmthHnh0Is2ucJx0UCxhN+m+bFVb
3sgXJcyEV9NtGUErhV2MvlhdOQQCmruWM82xgKhlMDf1FunvJm8AU6PbzV6UBExk7Kypg3dRqB7W
kD8HZ2dox/r1TjTO+bZBWPxqnW+ZWSeagKQGEgE6c2fQtRAkHex6XAk6c00x5Oz1C7+92NczdkGL
RBjn8PgKzNvULQlrw4mwRnID2qs0B6JrtZBVkKYyuxH0LdFWZ/42Hm9MzbISQBntgZIX5N+oShE7
79QQDseEIJ4WTD8t59Dqac2ZMbOq+Lh7Qh5SpDp7DxJAjwVxySultOgoWIdD4FYC5PlPJjwV6pGN
4CxoPOYLp/ukPFHPBnd8MwXGp/wvAeM5UZi9bh83NATYU4FWVyuoVmYmmlu3ZavcIUe7oBXwa//o
Bg6q5R6GZwYmFK96hPQffgj0Vr1JLn498HuMsdH/G4T+ki4QATMj77+ezoY/58XKckbbw5mxG3O0
MUDoYqKeamJtTfcQUFvkgFELzaBOqjQjvQoz+SVyVIv1z0pHrbK8Q8j1aS4SqKQ8qOkIG4u0ujUa
2RzfUnnpIYacs8ZHDnYB0iN5AnY/p1VvtR4T1OOiAd2WuB8FT3f+kWzW0Ixgbd8OSg1cy6w7QrZH
UeXa0hDCDbxM0vmynS48EnjhFCSb0n+ciqYsAoYjLUjmp9JXPop7H1N+pcVAb8kw/IOZelMZBH72
XfCGt2mKhDEhFSG+u3Swq+AMngfLZ0o+h/uvVHmuxhnXAvk6d2O4MVVSQbD+oRfDPG9JyTgIvU3G
R4R5BjItDCFBem0s0dRh8JJ7EpeyC0lr0LwoxMWKUStqO/SL+WsH8QN60r8+G1KNlbNgqJP+sYzF
1RsKroJcba2q47AsFvV3lGm0SqyHUsyx+y5eMHe6+PO/m1R8cBwjNi5YW4daBhRO2W4Mj2McyTeu
Xq0BhjiovnP2HGABQ8/z4VLH+aLBA1tW25q844IxKHc2M+y2xoJCkQoDHrZ4OFLjQaVBURiq3rR7
mBMFA0vQy+H0JB/RFGWlv12qaYaqupYx/0K3xIzy0u0aIW21Ia0Gs8zHpLAfYD3OsdfhEbQtpamR
nQxElEPngnTW/MNwmqBXPKPysULPNmbEiblVLtLD+i4cme8XafVMTXV5UflAWsSha1ur+ujnTvzX
vqZWaI9gXwJZ0bg6h2Qe8++tpvFayUMXgNLfi8Qje9QuKgW0LSxeQzBfmqs12S+DttCTzgn30l7K
veb2b0atidJbDPw601jUG4vOKiCKLPlKiDlSZ3rmzpqfdV7kBGe3q8uImhQrr5iWEZeD6x/AhR4M
gzUU7NhQ1zx7xYXMPwWEez1b2/tI5ftU2Xq/OC9wClsCoNeqIwTJBznU0GfBr2pPlK7p+UUOtmfR
DDppX9QbdW1jvZ3tfglctQhOUt9nNFsOnLDvGImeRvoRuRRwiDpuKXKsKyOXx8hGoQmyxOLaYo0Y
yZ28xOGQv+GETxI3+MDjFNfuf+vH8stilxQUaB3JfPf/Fhwau5rAZKYUwE74OAmOWuKiODCFaJZ2
2xahNQVYqkFn3sk9nY/m2EJBOT+IvF7tVBEGItAGjfq5egOTmmH8t3t6+a/gjIxMTu/FnCRxmJ1i
ocfmW3i6AyWjvoUJZYWietL8+MonyU2pMLia82owVlKDZDR8zgrcnl6Uh0AVc2n5ozJCi+sKNIiv
FDbUUlAKyopAls0In+s59TVxRXHBfdlZDPsUSIwIGOroSzpUFYw2w/K6670co70DH0/0sjzWW2R+
eA9od+ZazI9jlFxkqYxjXWQJoieuUyRt9P2+O/SoKF4PAr0/v9VOqMh4V8kRtGZry4oHS+PqOpIZ
7BFRpKHTNIiw9Np0IbDMIf2oY/7vbl+81FErM/kMUjhKGsi7bJg03l6xeOgOpwrKMKIUwkL2mSWn
fA0jqmW/cQWJoO7RJBr3lOOKMTuZLQwT2rYOxclny1g/7EUYfcrAN8XBLyT7WBLF8x/I67QN1IBP
XF9GUK9HcB/ruovND524SqP1xHHKNRmLq0X+CClqVMXh6GrSpap4jl9Prz0OTETQNFt+ZHwrWXHi
XGl8BMbZagpMTOOhKCpbwK+76wvmtTGw7KCjz93nPkxncsA3DCjekRwgtv4WudcP/HqZyCa7cV58
MCpX440+x+83Qs98FOTTbfsVH4TVe4FULA+wOLn6BJwSqc00+AQh//WSqOKDZRFUM8cnJa8obi88
i+GCUa4Jl4sd2C4UarRZdOwYhYYXfyQ3Z/KllcTogH9hV34UCZbocFO3+OxUjfEQW1YD9s6JDrkk
sO5NCW8SRHTUif+rxace1GSAAfN8FwHzY5ExNV0GSMzQj6XAylUFI/4KfadIJnd6KyBy4GRG/rfj
B0u/7UTx9/sL2xXbzL3DAgQuzyp64uiImAJdsFjKxX2fkXNZdQMX2xmRQ0r5A08HXj4tC1564n79
KpK2zhRdvxj0X9urNY7V9QcHky3TKcu/wj0IUmt6l8OR95kprCFV63pNDFCg5hmaF2Q28G+rEn90
gOhyN+Lf4KEWu/ks/3sAHoHnVURCSuwVrsm/c8rTqnM85nF76Vurc1YfmcVHfOpBI7QFXTmANvx9
7eDvAOjksQNhY7WUFOBtZzyYULuuj3xQOv/bw3TqCqdVd79tp7rgA0b8lCktZ+OyLYmxF8rn0evA
c16lldb5TfQlmzx6wXt8mPo5VILOytCwdDUd3S3hrJ0l8e/gYSllCkmF+pY6EEU19D7M8oc9bBcE
tkEpxsl8GTgDOobPSprGD97uwx4hZHUMSsrko5yqyMAGd/lIL+4J8sanKmO7rJIGwWGIaNtnrXqY
f6Sx/9x7J4OcdTPpkyaHTSNM4jAjwISKAzHMjn+G6qsYDSvTWkONdc4Dwnb5y0yWpCAqPtPXrRPX
Q2E033ew1UnaSnozmjnNOeaHGwkv9oJ3f5njMe8UKRxFG4ghw7vKksZJNeYc3NLC85zI9Dxj5Bgw
V4uBdUcAdPB6XjsI3D6fqqZ5GJbrukkx/ocgm4QR9fXpjIDz4s+Ql2seQ/8f6zQsCt/C6P4lIt/I
rz9JMov/lRNeoWDjTcgBefMwTN6gJ2rbup7fiuvCHoccEYSM7Rm/oSECKEXDC/6O9qQD7HRmJR02
+W3HM/j8cTs/taQzNgt5hRM+Wgah7SZ5R6o2M/Ubw2yB6TBcejgvf6/vNtUui7pfyUuO1h0dGzI7
Y6kOc1izNzrnWlHhDNzu6AvZdSzUGsA0bLPpfXzAMVMNlmwsgyauTTPHcWHyXtUVWLAM0ERlCTex
K1vWyR8zBwlKf7zWQ2EhMI2YCQIvSUBrd2r+t2EjlLbKTqyXMCvn0zy6R/bwKMfojdlz/RjTDRKm
a27/Fu+k5K/pgZ5vVUvWISgNQkoCa4L4QrSbHXjnA/bxfhLa7ZR3d6UAd3nhFzBD/YsWtFX+pP8W
Le0e2XhZi0MFT0PlOHfGpGTgoFbeaFA3NCYI5jcQCgDjUqjk/8PPG0blNurMPtF94HZQCXxK5bx1
pMm3vNVC/2dORJs25N4ZZI4/NashRhYKL5E3zGFq35zf9RyIkn9IGSCHiSfJtL/zCB+AExg6EaMe
xvdI0Yne6R3qTAiPcCpLzB+uai1ZO6w2Vi05WRtoHG2j+nSceeqELFPqn/nA1poPNE4FSHidmlfA
0AjRGLsakPL2bHsZB3g98plEckYABVLkHDabyJCpiIqCYly7HQIxZeLv6wR39XxnXTluf1qx5AFq
wdUCWHWZA73ZVv37TbDW7sGX4IYkYjNrqUSt9N0EM3vhfDjpcn0+v776+vJGg5JgRpjNkNWZk2Ut
HgOa6f933kGqxLww8KYtn9FwZtXX37yW1y+u46FZFvRytLLaUSp6SZwMNDP6fTMZr+ZNAl3yL975
JElS/Wnoee+BUMv1bk8c3zP91NutOsTzOK0WjztIqE6vQyWskun6Ce3p+cQUx76zWseXoECVhlhc
OUeEleBAyOtzDwMqTLCvWa4mFknf+2NEeuiHGieT8Huur9rhSsIstQf+aP7mekiMQHEyQT7IlTo6
yd+i396bg4UHsCNzVd/kTa7q+3SmyCbsB4O8esog6rjCW8qLuLQ/0CRHEiDcn9wVGvPhMh5v7O9O
NsxDS9GoWHW98Ur4og9vHLUqXNciZYFbsQOQpAb08omqnEPKE/c3p/IlWmvNU7xOerY2OZFF7VaL
DHFmAqPtzjkkPYCOCmROgytZYwnm0hKb7b0/ExR35rl6Yl9fQAkFIzMtl4mMZvOhfd84zeaiB878
MRnJOuRwrIm9YtplNdwp+BHmyzjtcdSZiQzMqvvQYAdAMVmrYFfwS3HgCKih6biD/0Py84NIvcHp
zL+LKJ8ayUBBE+XqD5kFx29sSf5J1QEMX20BdDXXXI+zzXM2+mSj+umskQ92V+lXIJ6ZlENCirZT
WtOyr+SoAi0PZABp+99+uzwB+RHat6ei8Jdu8DGspZNiavyH/lNNesiUUnrEHzP74fOx+8qh+wk2
xK03Gg2RVK95s/oyRPs0tOi6jwIvQtoQCLB42fJfD7s7sIobEQ2/CRXYljtWg6K9r4BDVUlpYWn5
IBaU6T2jf1+CO3+jSZpaz+5OvaUD197duZS+SmV4txB/y/LNgDPeklzBV6k6LzmwvgHEHANSrLiu
ygG62LhCJjp16ucQGlKFpaK10qGjppCDs7v22y2EA/mxVEWWSISaqgKck8ZjM3qQ3kWxlmWBrpzp
gSiENwAkUUQP7djCb2DoFAkfzCHPI9qE88NoVg+8mu/g56PVqhKss8W4d7C8DU699N8J920A2SRO
TZL/EWwdjtwGrNAgb9MZ/MKNVpHmaDGvg22kCVcCUVs7gMuybvBzCu3BMIqSF8Eqc5vlntzcTBv8
bd7DUNiHiIgItqYAboBjeea5Ax425WirXFVXWRWscch47ZD4lm6JEEkhTI6f2jLGFhBEZEIM+R1v
D2Cp9aGLoZZ5N/sUzkOjrOgOpL3h4wDN/D2YbXGfbYe/uz5Y5lsBsMPJJPXjRyXUcHd9GLGF52DR
CBqPL7lrgw99a9Z9I+txbdt8Z94yGNEPIus7cL2FaTpUDibc3LIs7t6CDW7bwYDLjVSh6lLn5RnK
RRnKCMI1ha3FNep+yTWDK0A+ep3cMut9/DakWjLH2XbvnH7+lHB4xMmfV4oze/UCUtoK9kQcOZtN
fK+Zgm4qee1PvdVtm0os5GTmvtH9XR2sf15zvCarwmYGfDbV8CwgMbMSww/eTja2U5hzK/A5HfQ2
T3asI+amAfRlxQ3NOJ0KYvIdiJ//gl7EFz58ADZmGlq+eW9Gg9owTO4LkiYMvRL/1b9RuTWji2kE
c699iR0n4EOFXUbaRhPKyJRUfHoz+OCH7/L5sjwVSvRNvFAuby4yepoXWn/njcnKJxV4abQduNqD
fn5D3yXH4nUeFrDv8oXPx0j5ylVkqTuXk9ONuMCBhT5f1S6Ex5wF50Qiuec2z4fdgMclPrdgdw7E
IJLAyHTm/BKR/xTfC0bj7jGwlWwtve4kQ+c+hW+p1kSultfWfC0Mb66Ur9Wa9nAn0QSnbruEytej
SpEkwGWoqNhO9Z36jnijOyHIpSy9BL2/m73LSV1H2ZNTWJaj2VRKsph9tNWIbwFW+B80E9tR0DJQ
dscTnESmtsyaZmHRizKoC9WnPZfB8Gnm4Bk3rT4AflgFRxT96yrggQJ9q+LGRJ0at1KWsgq+gPhQ
be2NsNsVeuTWjGHlMqD7/J/ufMSCbh8AlE0FXT7Vfbr7f5Bn5uDXmGoAN264fgEloX3Ce7oRiGuY
oqY4XEJLpJfUNP9eRMfS0ULc7BWJW2PyUMM6dod3Fmzu7afheksYDJ1vcRi8OlgGFFsx7C5T4ja1
zVhdjsdpVwrrBE2m6+sFTIVsAkyhhOcppFvM+gFbum9EjBceAgUHd91VeQn9LFX9TR0j3XMluQPL
2WAZZLJm35vh4LMZMPXEUl2sjPWUBM55nM1v6Ga+Jht81y5TG+afPg6aC7d3BhxumrxFyDu0y2n1
mtf13iRA1ZUJL0M9uZaBdMJTx40OCGFD5uN74XqPJz1gfczjvJDqk1Upy//UUD5OdI6V+8bTaQgn
+e5LrLyiIPMcmcKG6ZDLnFZSVlhdGddnHYxEk4KyyPkypTidDBz9FvugqNUPcEWj7RZuq0YbjEK2
GrWInmVQGw9/2R0fS+YStOqML3KL6vRIpI5WqukeX7z46bW0LU6ac+eeiiGe5fXDmHt4PNrSvqPs
Q4w5ns8cIf88a4CyOumvH1UBWkoBBZlXSjiR4mF3RCILApb8wjQu0xST2/Ew5v1r01TMREMTPo2n
oV396gNzbs2q//Hg5uo3oTUr1Lp0YISevfulR4D4zCTWM7zSOjsRU6LU+97qsiLHiU8lADgY85M3
PRX5HF+vV5qbPeXTRDJ0r3D+Ybkzvz3Q5PFl+IJuMF8x/VBfApXPA0qUYJT269JG/jYv5zEGFlCL
SFZ+TP3OVAHiQezZSIcuAtS0CEIPIs7o6EEbCMvX3rwgnL/WzN/aWOW23YgTge3uXIwxa1bTYrBl
tXgHDkASwAHzXrCskkv2iOSjklqofHNEVcsHSRD2WF5K8YWurNB7Qvy7KBGPoR6kEnHtCNNj46Mz
Ba0EEzrx2qFU/5MfMhmtfWyRO/I81CNynNAAY7Uj176S0/+IVHGW3wv0rIX47z3KY9Ft88psARNt
Fl9tsKqma+tlz1ey4v1k7o5NVwakOVb/kFjtntoLXT3Su7aI+M2ouxPPGYWYwRR9O4hPx0Bv7sw7
6xOPQrNDaoxSin8w0dNHFB0Nj+AWQXOM6vd8kwfbmZfoV1yuhIfoD5yDZj/wywk0y80qjCoIIkTd
t6Pw/zcmz5hga4RD4iUNyeb6J+UbLNXFViqfCplrQW2pkdJo5eZTAOgot9Zk7mYJWU0F1/fGuwZ1
vLY5H8IxMBur4QyaL7277Vhuprvs97sbUIhDAFdWpp8hW20FFTY/iRYdlN+fB+ou4IG7Snuy9RWf
xAYetURGlzzlo1IVclWaxGtc2qo2MtofZFIudaAbypwXDcEbq3MNluSpsu1lwILxZY+gr8+0YqHf
mfKiFLn8D1GIWvvlYtG3dlOgp8tG70ARpRl5XMk9oJbQRJLwXuG06mPpUQhNMMQcfgUlDxSvzyL7
QK6YH7c+2SU41X6CDSRzGQRySWKnJWcZVeCeXpK19c1oLGbwIJId8FU5FFLHa1vOF6Pp8jqF92ju
8kK0OymnD97TieNohT5BWvw4JRQRopkRFdu+HSHyVZ/OjAbtMaULv4VR4H7KvfQoeC/LtNr2v9yv
E86XAmeFVjmemZ4dzjeLuxkAuY3Ky5002O5VsbBOHiAGN8k68iM+rCdzRDeXf+r3m1LVBBnrWZ4w
jsIs8PFsANLvyT1yltflfpgoBv+DsNjMwnAeJZfWcWcbxsbF/OvyUuPxBpcvgizo80n/XFoYP1FL
R2pAaFfLKcNiRH4j3FcHd1jQ/VBW7XuLZx9ZfHBEthYUp6J43Om/pY1KIRUrvypQzIaulj5B0tWi
qXZrrzOhu4Fns5LAMrWCM3e4zwvdtYxbWyJPllEUpLtQmvks345AUR5JzGruO8lga0HdeYmXUY35
KqwCR7lubX3fRjWhnZkYBDfaTzHWM/kWcJdVz4H96BqqOUIRqw75vAuqCN7VvnDYaEWI/Ho3GfkS
XEzcVl6wgzH/vs8TfkjqopdlNN/3A5Qa+oy/oayq0l0f7plLnmQdn9pWhHnso0mS6MiUZtnh4DA7
hdgq5BY+7ykJLEelhYhP3YOKS1Y2w8xc7S2Zl+Lx6+5AajmzAZdQzbQXg7YPEKkZSgDSp7x1waOB
bHwNdYkCAXIFc87h8sb9KUmg/EaDJywZJXbtS4TmoIWOMQF9RlLqLTp1vnG4C7HAUGyWwI0BVOTQ
lkr7QsE4wjQkChGTenEQSyF6E4IpGZzc1T7C3IhhudxNpVBc79EZyMLjFE0hC11ZtGTkzjni7q78
OUhkwhJB2tIBvvIUFbORhfmQhgmqiH/bXNoxEhmjMllkLJV81rBn4QxIlKHbUbdalfn7XwCYszqO
ip94QmILOSDaFUap4EK/UElhIR9FKdeNrODnRzo3ed4TJQxCZjzUD5kE1Nio4a6oiBssBcWK4qj7
aUC80kpjhcvzI+TZjbTjv+JIxaPCh0JnNmeRmElFK58wmJdQFuK9zoNFlywKeW1PXyRJyPa3w2wB
mdJi2/WddZ4H5/uLXNHQFbQY68er8DRp43C8mW1mSkF35HVE2uSEJ2S37Wdwls/OSUe9BzhFQbX+
1Kg0dZw/zD3WWp2a0/os2lZwkyA8/nvVtnvkOwzEAkj0PNStct8PwsH4Cay+fsIi2SBWjA7QJlqw
e5PgXPQplCjma8NnAZNetmZkMDtTTsQjKzdCrJwOZbDVjCV6A7HJ8i7x6FSXd8Oa3s2bNQjccKQn
mtaWn0477ncruS8ITRLtXpG/zyOEo7yRxFweYQZ9cYSEWzukAZLqpmPNNQ+IIHKGbsWoNHxKzT7z
paLRrVHoO/4BtzP0namQESg5Z9mSon9V+kbP+NBN94ijAaz/pxTatE0qJDST84rWlx1NIfwIbvOP
fuJf6vSGnBYpgnqvmUeJmMp1+A+BC9Ejb/Vc3KMWbNTgmvZZmWvbhzk3LYQpRdPfygh6WQxgRQXU
kCQqExzZAptMvISAlVa2vN9ATeIvdC/1fyYlwQt3WT5RGkmg7Z9sactS7pr+63/ACRNVnhGvplWV
obVMYaDsZlN800zSJgekCl5BIsj+UZuLq3sj81ml6bT/svDBwPVeXBpgRDKN9dRFDycvlctiMb2V
8Nsgf8SKnI3L8cyW73khXq4V6XC8V5iwtnjGP4b6X/gI5LJ7GKz59uY6LiH5InvYTvwpOxRhCA8O
Qu0QPQdW9ALWalazoNkK3Dm7kO9AOhGY0RzWAf50U7TeLiZBtFvMGysaIJtLKYLUP+6YfEAvcOH2
m99rDFQ/mkQ1AZUr3VMaXc8jBlInmCnaI2SFsS1SS0srY2oBrBjBrSheMTPngOQf3amzNsnY0zzh
zaZ73X44F9zXqKRRbRs+g93OCxCSJDGyqVlALH3cLhVqvupa5nBlS2pC9BOwDbaLQ63LYCFMCFfc
6JKR3mVPsJuJVfLbltWKsfKKuQY1V+yoDmHT+wuW7vbTfp7/Z6HimFqxTzWWWmJSuoGDPfNkLOqr
AkXHE/ed88ofI+KVq76YSELMhMBg2toUjvA452JVBktOTfrkNP1eXopLGtS/DEXU0ZOC0a3W8hkZ
EkuRShN4vvCn3uFeUfHJU7rhA5SZyzmRXqROanmabLLXDG7CJuXg9/SbL0m8SEFkfRJ68cex3him
i3yqmtcI2+0n10NAAYG4rvHXhLeV+h8hqMXv5WdeCu4qwAzinlgt2BkmSAfiFdRiVIL3jgPnNo5L
73bgjHbbeM1ibTyGPxfkf/TV4MJ37h2Taqb2ZWwhlMIHTLAZGefzg8LoFvSGGBFti6rSyb/Ey1lv
BduQG017OhARsPchJhjI782ILcW511JYfBy3PBMj4pTt5gAd6dXUQ+BV0qtSSuIgcn46qTcsCS/J
rwe7IHyvnArglYAMVAEBTNWoM5YkAgpiIdjjF0hwG2nK/yEyCT8OZ3vnAQZC19WoCmqudps/fver
T4CVNuvoMIZdwCPcsL7cy6c15DXAdgzB5dGCQdrEFCEXbArBlkyAHCE0CN58RsGffIqbaPyAqsyW
yskRH+8MpED+i/SGmkYAN2i22nQDAT2mvVMOIL2k6uexX0fySnP54DcQdEmPOAQJLBO+FqGQz+Ky
FUM3Oem6NPMMS0SFlvLZlxugzPmSpaVyI81IeexGNz9cdDOuk0eEWlgSui9ky7q4H0QiqFaMWX+Y
x6IyglplDQkQ7kkZ+bYnaQ+DApoiAVumcy7Bam6fCAIIS8prO3nlK3OahYEUDki3kc23ndtb7lx7
3PQ+mrgezenPud9uafIm0itBQo/c1vJfMct8iDa+9MaTq0KwY7SGJ0gUsYrLC5Auq1EoRVd23Gel
h+UFXlbRPs51uTYVDo9aBMr+o76bjugHOoQCIAoyz0+xJfSoA+Azfbi6LbGxWryJk0EgsTnNE5pY
gwUzvfrr60qJordKC0mkUFZ6kh/AZVnTjOK36CtI2XkNAAfwyU7duWAwzQpHv79K+qqwV+aeCKS+
fnhg91E/0FX8zlDoxHSgRlV2QYIE8MCyydL9Yb4savm/OvW+vsY/vhJDll0m8dFWkBgsV7bvmP0F
+CnzTAMGdat02MnlrDEKI/thl9sNEr6nGOY+T6x7wCdfLlXEabI1e9S1/BfK/JpdN6sdINoTVttO
ng7TY6bVNvq7fSHuxBSgUwSqoT/NVzmKDC9V3z1d4EGl5+qOEAg3sW68E0mH5wpUkhoHj4Cw2Rtx
KPPHaxzLbUfGrnFZZe06YP5SsegDu3jqYlCoSoz0tGC1Gkxuh77Iwlrgb+L9Np4pKNzQqx/oth2p
H1MOP8C/vLlGPnURzoj028UdTxwyv+ZkIL8uJNqrAi+1uIj1ezxdD+Y3mh5s4vOFzFkCJFQvFkj3
oAN8GiAeSGC/5JTdOK3GNDMz0bvlY0TttxF+GDA2w5HcgoSPsUehXIkuRaJqWbs8HWLDj9uwF7iv
znVpzsUW3jvTw1pBDwPsqtGFe5p2ZpswyLKoZs/ANeGnR8n/dKvaRw3y74Haob+WiemTNKKcTSUf
kWJBskfi92rfFrANcSNrUAz4tsC1XiOuC0+ofqgA98743QKOd/u1lK6KbuSwXwd9e6wZWSQ+YbAZ
RnJ6UFIgo/95Yj1Dvc7tZ61RMdSn7vmQhQfp8ESEN7YYg/7Cwpgz8BiXRldiKbnc5f9KLdu54cR8
wJRMj8CklP4IfuBsfdz79TLnYYSNH8OM76iAeGDSqCAgJIF6dojQ3dFlpmSUqg00qAuOPThXzb1K
uAeQ4fH5POd7ilZLj+kTicsskdX9MzcKIoRI9N6IBM2in+BoBcDbuN5pdEsB3b78Oz5KviRp3/8E
Kc1gcGiAkpqJufKxqNRtRuLDvjKlybhAQdJSWD0fXp6ey9HQ4gIskj31d9MQH84xZlu6ZUAcnkmd
iCE1HpkIQcF65NZeg3MTyloJpWZ1zufxeyZL68Ph+TVKApWWk2aD2Q+sWKXvuYPgMNNzaw3M/ajg
7uzYTgzkKxy73DaItJSQO2NVkEOjv5BW0ZtmaIh6e2R48Of6kZ8Avgm/ZpzIsNfR+MjcGRKdZlIl
+7jYnrqKD++epJBkr/9msm0bJXREQbGrgZpMV0KWrKGuBPWCPoSc5VEyAtszUoFbHlYAgM0kOD0o
npJvV3QPbqdWLg8CYSfPsozinn/Sl561vteY0qU+AA9XsJedGAamK8PHQua4oVvnV4nGMCU1Gzh1
tAC/YYt34vQyrzk4V7O2c2ttDkyz9ucUgUMGosl/rQQ77F0eU6ccz71r+FNKT/K80kOsOHb89q9s
zAS2tzP+KeKtH9bhb6nCWLBrf2yIvucTA+Bb55pdzYHOF7ZgjduLlWPMpV9ea0g1VP/0GPufdP60
7ZTgk39+WAA9ZLFPMknJ19A6oDys9ZamUqbcAgFwZKh2WkfvI6Z3Dqpp89sW9w8eV0yU3MH6Fdzx
qVgKhqo0fLPubFnFLEGEeKHoejzhb/eqt4A2bgvepp5+66hIXZA6ev6TMxXD70Sv4T3RmKB3zVMi
NyaJuV2x3mToRlxBE0GSq2N0jWgPGXkPPCQhDHz4yuHIjaGct7X3syHQMcPLV3LVHALJV/hXyQfH
tzzijBzrDeDRU80CowGRPpsHxOWFpLpd0CUU7LD1tw5WL00hL08Q6p3C9fxgUtr/D13LMTO2+pfe
Lo+Gk8azsqZpAGZkN0r9gnSE3Nbe7fNH670vl8hhCrsJpUjETjy6gHCXWEe9syo0QGXIsHTbs5w1
W7SNYmW0+M/+cpTIdgxSTSEBGgEJ6rd0OvpN6psAOrAxZZin9onWUvSyO8LKTcBzx8pnUnOQ+hUR
a9QiJQrITZFzkzJSF0CqmGysOVVXf6Pwe/+TttEC3pyqVXr7Gnu+w0wcV4a+oqKLFvAgf8uN0wGS
bdVq5hzoHJUO+TPApi6XdYI+NR1oDC1iD+X3rvKq3BeeybfoVv0b0dQfRxaQMZSL+gZls++48nX1
8yzpMEOzvpDdrxW5k93UoJRRkCZwOSy2F3q1Kk3Cdf8wmnLCtYMKf/iO3fE0eDUZlHtpiSVPn7sE
xe8RP7JQmRIbuuDbOYrPAq1nPb6W5WOY/v27DcRnzPDj84tSiRYNckD1cNrjGG/09BlS7ZcmpJvq
PsCqCuuv5IzzcMCZqVGMEJXy6Jjmkw/DnDYmGlm1Z+LXW0XgMdHVh3J+K0rZeKTsn3hF1nWBBoIS
BarY5wwPjJivqGG450NDAVwWlwAK/NcNpgELoRAMYjAk0LThMMm9ixF+/SF4S+wqYZ6WNaejw8Ak
cEfgFc+dnDKW+AWtckjqLp0wuHjxntGdGiOxWeHH/sRThL3i4a4WDH531BLZIIki5Ad2bee0Igoj
KhSog935UDtdXGRLQh13LPB2f1SIwiSdhDkP+0eEeEj588eJzxVp56yuCEHUi7fWp5mk8BgCKlmJ
KfQ3B2zrscj6h/E4WxCSwCnRs12uF1raWbrOjlPXgYi87jkBk+FYOU6XmL/pq8cJPHc4KPHTLVsn
gLpZGqUSeJupyKPEqh36repnTRkRFHaLl3ijvoXyARBcT4HrskmOYKWoT6gMZnxHyQbRNweYJWg2
plQuEo60lhsJ3XeNx1nwSzCNFaTiZ2+N4EPIEyekFmFOnuFNSWz9NM1mLkLetMlC9qANczim6+YC
ep63+jPewB1SkVkDMYwvocpjKf9zpmWhmLdFZ7939YqAT3vayeEdEufn59C0ljh4BR+hlrJDeiLw
/ZqNz023OLO5Wu/3vwNK2dGw7ldaWQuIv+HHEQgofRWxgq+8HT1jOyyqQ6touwe7Q2g01y7EO79h
F1XCkaF557mKv63EHtmwDJJzjAo7ImCIyPwRAZYAkum90AQuZ091+I82U/ZSeEeZAYVCzrTJE5qz
v4t39+855TQqgGT5kDgBSCGjQqdgkgBzdRIUmKoZ4iNst1910IeS7h/+FZpf6VWQZ5O5LMQtRZYP
qP7zonAxmOHRvZFLNcL5HCixVJBqWuJEI6StMSanIRJmoce3fOUV0lBLM4+DjYK+k5GkLmwGrH/W
Zgj20znjSyv+B2zhlPQKiHFJ8JtVxnRcrck3x5Auqjw9JLBRsXTvT682fFYcX+VhYT2HQVIbqwmC
30MvFX8QqJetMkcAyelDjAUVnyGXMCYmJrVfmbaPF2xtYws8LwmO0RvYIUTnl9aZkSZXNe032JGP
LeQ4/hkRIHjZLxPac/DWMqee5p18DSDU/cAjbfLO144YFA3OROrV7Ek0nfWPVe1FktJ/V5u1kn6Z
ylvtnOhL1oaL4U4K/sFWwOGkFBuq0mxuhtPrQsl3Iv75lkgZrgFhtS8+WQ52vVC4eaD0t/h0vt6+
PCw9HWxiMdpv2v4Gtg0tybVFsgYOwxXYnCCYXKdrVnVobsMunCf9jnTejZ1o6pe7MqOqSHeiLESb
W5fHBXESLahJYCKXBln/erR06vROSXZ6QnttqzXhklIugm+XvMo9q3gOrFpdKT5t/8rk2eE1Oz8n
GalDEKZkNVZoj9NNDuhWGeUdPgYleaawMSQKeFTy0uCZ3KUNTcekj16ewMJz49F42opghjwH6oJP
Xlgnm6WCVzOznEB1bjDkrl/E25LSJJUNwL6yvsPpXn/R+YzkD4/A0i0jLbwZRtAMhfm0hjyrrw7c
fV1itovlmmaa7mcKMUK7Vf8CJnqlXYB8d9YroSzmX/kxQc1aupRCnPmbYjHq0eCu9SQUzUX2wygB
XOs55Qg1mkDr8DO9mHVelyqRzG1cv6TgWmLfya4MUPoJT/qL+Upj2l5NhCUpIRWaW8eKepYuWvpz
rgK/FuLGaALDwh/laV/K0nLz6RjDvAaTtkvEeV3f80zCRhoNcEBtrIDUJntXw2nxDD2DNaVrs8Xm
9YsRG0nlK8g4YTlicVgAVmb8tNsQQiOF+vSc/YcCizZNCC38BDH4/s+5TWXSRo+95Qbus3nKXYJL
urQyXAF9racvFy2TqzmyJRKP1pOu1YDaCIMXpTtXrCRsoON6Dh6IKNrMphZwCbL6RZsZUycebNUG
oLRUeAsVHAjqftXzgMRjTtStOMIHdyBHvjub6CsLqYosFGWLiToVdEdqtmAB3O+thozB5B6t/jsi
YYutWEquEkrZsLbOs521Y2PlTBcUF/omMe/OJQlL+smJSZBo0vSbU1jLDk0iVb6yyE/vVfZlh5UR
Ow0pWcBNbMFtm8G4Rm9uxXWU/x6dQaCxSt8CPdx4HGhJ59OiTJ+xvNKLdmlB+e/2fe0qZvjVtkKS
iWvLVo6OnKb+H8+NVIRn4zjC2yasyzklZ3dwZ3+GwYVroWdrTaOK7ymatpXEGBEMjIL5Yu51MrIJ
6ypz2i9heQ1RFzqcpgL0fZn7B1cJmAlvzPdxseCw43qOEm+WY9k/NpdjgsWPzt5hQ6+pnbkZoaBC
6EfT1k1EyZ+sbexEpLXFf1AhUURjnR4byQtEKv9f+c4B+BvpdLdehVq2gncYjaqInr2mSVejpivS
3m/ceU9JLEhWw5HtKI1J8ZqkOeoy/SmR+CMot1i3uaz/1Pji0tFChb9K4qLLoK+cU8Cii9IUQ3r3
dSofDTkB7ayQi7jPD3bhhXJjij866Uhfd4sLQj3uoMuS5OEmXj85rJnh/HINVeEgNaypfHqTBja6
4VkaGXoPIIS2/MBoILpZPirzPGy0zYE58YIzqGP2jBKvSX0NQ04hJtjWMaZvyfHUKv15zz/3VoNC
225TD+fPcHlX3bba6V6xx+nbc9Za7mD4sz41fTYkdJb0puXayINA+ytys50Nbcf4cnxIf9b5kq0O
cPDtl8KnLif4hfNqlonF/CsKOxSJEuS7t6vuwAKWR5yxWK3IeV/QGgaiHNm3BWJEUkoyaEgiBvCG
iRYb8XLJots+YNrgWZbh6X88XWBmVVydztI9JSG4w5zLQ39fK5CayJW2Dt+hYVWPzFcnlWGroRsV
29DVEJHuQLQywM1dAgYt4QU2LYi0+kLXU14L5BpwADJ9722dW9mKz6fwHUn7yYNwwKrs2XxtXVPs
M9lApgbz9Bq4pxoEKAT8hl7FFHs/8bDWGZh6zGuOHES4ZoQgO+QdBmVokPZ8D8/HaH08gQ5qj1qY
PfMnqNnz1N5VqPj74THfS6p6OrYOMgrMkPecz/ERgyoYqUpCg+xKpKhvqw3G0q3l2+M4VZX0/Ro5
G4c++GdIo70hCoSPEmIVQejaTIQMI1jPapld+4f8UlIw0yWOhZT0woh9jl4tEDLaIOK16U86nG5I
TsAz4ffP9s5YOMCcwWDaCdHrQkwpdhKakMvnyhA9VFi+z2R7NBVQ7hsf9qBozsGYknzETDqIHISz
N3sZMgJIrR/02CJbM9210PiJNdHnYqvU02XQY/EXMtC3+/Or/xjQR9/h2UfQ++H5JwLIvwVu0zZz
JrkwwBDkMM5kMt6nr/ulJwPpa5AYPkgW+BQxQunHFy3qTUzYqS4GoTRQWLLRQ+o0xBop7Saxc4Ix
+oB87rjqZSyMA5eaoQXJkCSGzuAaAKN7iiXv77CbsvtXNcp2fBfxa4MpUX1BRApfVp44dEDS7wjN
XQi8zMJ/AzETgputhmSL72/Mz5Mo4gs5thNDcO+QkmCTPlEWBKjeItvnaAllm2nVh/jD7dEZWY+a
53Mr5sNbMJKVukMvcxgKZ8fgRfzb69xlVYtN8cT4qpUPkvSvhX0stew9IjgpPN0JWhxircxydvKF
BMhtuWPFbHiA70aq4rk112Q+vAI1jbvDKh0xIVFfCf1lbr3vFQ5o13pc4tf0iHjbmOM+PQNAoZ2M
BZfl4P5GLagsHb1x50FujQeYrcV0PnAItMhAKJdOVwZx1BzSVtN6jbEeEb1qvTq8X8U6ank9lAcG
VHcUZ7VKX98eHs7k9j7NNZJqTM+Q/sJkreagaXpukyhyDKLysedDSVvKvtJGOqYlZlwLiOGQcmx9
aNbY5BB2LN88eTnx7rbnTRZMNheNfxuj/9McUU+JrrFEDQmP1G3RQWJODPIAccu2XQgbneYWaGG7
SSrA/3SQ0QmSMIQeEVGKgGKXmCwGkTUsJsZa6dHjqZL/glEB8F2hbsQyYMuzH+2n5P+rxbXaWWdJ
sE5DAnhICyH7DL/63uyW6N+MZ/F53uU7HpPbObKNmGtgW7SAZnDHyga4BHI+ofBSPNw2ggq2Dv6s
BvrKW7p6cAFmzWyB+uD097yu5yrxyI+GlcHtHRMJuK6e4oep02RlCtMMHYJHscAfLz7Pahn8RZfq
yN6VpECoAuV/aScR/Ys5bCPXIRAW4i0YUucdNiSOhC5CmJjA4XxoE24sZlDdbLtjRlB2qFCJyfRs
AJ2Zwad9b5hh998SOw23c4oWmwZyHi8L/VWLKvw1oVrGE/57Zm/wpBfOZXC1ngpjUAzfyHa5BkM4
YsPQ+5iji6UFZEFBXcVL+vXcU/TOQCUY8/Ue6sQKJ/AaEQPnBklgjSzPhqKae9e31dwGcPeiFad6
WgM+H4yJblVHR4Pf9jscu9VmKZkau5SIxEa7a0Ola8jR6Z8z8yy/UvnCDhkcDv4UdyoQ/F9yQJX/
DOsH25Z9ScrS/wCfrSFvHA5QuK7f+w68ZgIR6FAnexMJ/3pyhDBWcjICasMScuBmh2/jEdYTf0Lv
+2myTHC17MStwIPB0JDltJWZUAOKi46WVwY6Wmn1T/V+BVV/3FibLPcexPF2wcpZP//YF6UMgVmL
8zYTsHuO7ccfvOScYrZJ17txL2l0jLnaa2Bj1VgnpDWT20i5KxzaUYuGFQU/F/Yxg65CVV1rXFqW
hp+Jq9ondxuEBMIl94biajH8IW56oD2GjASa45mr7ZCgWwRmKPXze2hetKU7hTzZUrxue15OpQnc
QcmZlyGsZMTsa5YUWU4sr0fFoZdyU6DS3XUwsNC8sqDqXxCxAguQS2abuW8hDxHigVWqw+ifC5N6
J8Wi65JMS42RKjQP+NfG3gCM2NS4KXtRh0bVeqdlL9qP4NTOU2tXnO0qn3dW5GI0tu7MGm0ufy6F
51tj8A0lxMduGVEJnxg0aviYOOYzxAz0XCykcIMYgAidaaDQuHkWGcXZt8SVIJtVhqa7TgH8Nv3G
X7nH5pmlzpQivMyCDS2f9LJasQxXm4xE7pvbFqgMVYY0ZK5qF6m7AhrAhgFK5h2Bng1hpMSI6zwF
ssrqmXdiV8S0Es8dnVwpeYCxHPRy6ek1n2QTMQTxNslcYcAM437CvdKerqViPb9fNKcVGrlPPBuS
idYiAaVC3Z6Rnohl99ZB3UayTwUK/8gUah7Yaqg0X6iwxGcUcEBE1Ig9Ys1mP9ocAcMRQcpH1ygP
2ZqDYpPAfE1N4j2OtdzDgLERShEqFv8e399XN2V1kw0LSr9soErSuUr+cvBcZN4GeLSmkWNsd+5s
A1WiIUu+zAozrmbHGGhK5P/51BU64nPlp4CZLeX9KQlwvTQqRliE1RhmU6kppSI/ePut7n2j5LtV
QFBfpCKuVqJg7wOcnT9vCxuQzZSgnNADdNNL8iElRn57Tg8EQc6/XBmusAS1wmltAdePEIbHmi4y
24SVY+QQLzc0Ia9PKBKZMlNaYfd6abVVBVvuUxHHX3qwdA2ctt3f6VpXFhq26Qo60XYEB3ib0SNg
zO0LVD+duvjyMUGsGt7QG/u14lEm6o8ejQjf5dolLqpyfm1MiEkVF9FhWsTP+8wJlNTdoGSEiVf9
WiG0pdYa6x1JoRoELQJOdJANB+6S9ZigGqZEYCr55R8JONPbsDljlwRe5bOLnoe2GP5rSu0q39KS
4Ff0WwaoVITomnQphGrecWr9jRcwV5J0G8Y0Mwrup4mi7t/Gl7OVPEZ8xCzOLZMUj3DhVVgi2AIk
q5JeucQSt8qRMQShzEVMMNuAGUytuS8zBhhmmzHxpmtjIxNlShhOAmifxT+7d9Qtnij+AZdCk5zP
t86h95/xOmdVFWPWyguKpO3ig52pKMhfUjD+K/9MMmXb6v+jFAZGg5IPMhacyGtFPuIQbYn8cdO+
l+N2+PC7NGDZWmF77D2wQ7ihu01AOIoAPuSLBs7J2qbfrMPRxf3j3afZsEHnBQ+fEtQ2LvhXXijX
qww3yjbRNJin1UXUknENFZwifyI9NCM0XzgnPU5OiipDDLXUJ1D/H39b+0haPdod/7gC7MMxn9s7
awkiGCaOC5q0sw5vZYCFrxNw1VKebXx9MTw0TJ7RATkrc/DgmUYSSI4Z77LrQPqfbPIt9aRSxSKW
blLmVYKwm5AJifi0t3cZrYvf152QqtJzFzABfMbDlozJgc5Xy7mUqZ/M/Zu7ogJnuILQUwCpz4+r
1nSj1HMskfqc8pu/Ajrvdvtf+3X7acJPXycp6VdR3lwpjTBsR/rJCbQjt913i0VivHVd5T6RSpa+
qtRltGt+A3cWoJXFGHele7hEfuo01RtwuqCMxNAYWeKrTF7zJ5Joh4cT/DzEVEO76w0IQD5Gz9rd
W4xsZLAc07tVE16eYp6k/Ts8JYEMXbx8wSUx4bJO3jmBJVCzTXtK6XS2vxx1zy/qpMpjVMr6iS16
X4M593Shjyv5tP1wJ8PTdvh8UO6n8ktpWEfxND10QWnW3oycInSGwfs8kjYFTxaIJZM4wRvvipOD
VT8FQym52OFjhc5SZ4C+v3GcuA57jIguMtPRY7hYMOAZuGVhoW0XPUGSpGbxwIMet62ad8d7gZih
Vj7ZKxISXKpaniU/EFgP94MHsa0fW9cWsiM1C3UPobqrAQ7nYj1OJkeh8L1v0jBbgZQhz4+QQcyh
6fXhmSsWpqP5g0fhPWsaWnKbgbDuuqWZ/fqB3XO9kyUyMEIvdV8AvUU/32q7ppUqsPMOAmmYB0Qn
bspBBsFuavNtAAh8nxrfTL43xv1DAt5Xishom6dt6PvEuacAqLs9af0J9bAQU3Keo+r+3DoL9Rnd
iNwHJ6I9mRu1qdyPHYjeqYYJf9ud7ODCB4AcxO1qgNZ5gIAdG2m9/tEFB4gXdBW7C1CRW7m59tu6
Og3UX6nUZfswni/oGRRjWgX4+H17F9+wh78Br590pfUNfSP3GWV2ekO6trl3ygCh4Lm6ArEPp9B4
whLY2najx6PUn3rmd9y2qyJhygyYN7FdGOvoslax6Tel834beewznmgI7M0OseU+D54q/1fipmA+
xM2XbtgnalFVTrVcBTVtYnv/61zdXoBBITtzuukCTEtJN1JHJRILfg9Oh0KkLjMMBOvv3eDWT6u9
V25wI+vj62I4fmntplc/jB4QMWmzkKouL0NzYfHC+i0humPTFnpzF34/9P91fbpiAs54o0f979ES
PPPzphOYNTicHLBMx1sXIH6JqYuvIkR24ZEzV1UU/2L46SfpVbMfIdou6pbtv8ky5KVzQmkvKg+h
xM2uoEyKwpQaL0C8oFffZiiq4HosjdqUzGtmJVyyT7nAQbfPsrTGTNPseMYEoxs2o148TN98ELue
rObKkrvhgGFfYWSBEIJ0WzBRaXgVklFcDV46rDKuiDalvHlv5grefVTI0eVUbikuIfbb8P918pnz
VOAMjINM0JWDS1r+ib0cgKwYNRX6LFdUGNZRXUtfhgX+YrzlNavZNT+PWYttgik/fWEKxs5A57TN
vrJIiYIz/8CD00uzM/Xi1e+oUKIk074rT2ZyPn6Q03SOrP17lUUy9DgSYZ4NQRETU/FgbzLFLtST
u6jY/jA1kCOabU9Am8Kpsts6DozgKMizUcYLcDh+ZjsnUcjvUBkruOflHAnjYlSMdVU1WD0n1JuS
FXwhrqGlYVYcyH334uYCIbj6SEkqY291HCOR+sGAb88lfSBqZBMTHLlj5+GWBpeZov5IkB75XhzO
3sPIa0Sv+a9Xrt2AYkmy4yalCpvS6FBbe2nAmdvol6eMvCP7nio8O/Y4JCDvBDag5s2USdTM33Df
k/6IlfZsVxOu+PgW3rkopWLD40WdYatoyC1ziLWN7Odq8q6VSs5x2LhdRkgBrGXOtC9eZKzsY/ka
GC+R/cYu85zHCxI9vy1MCQfxO3NU7uulTriHszorgCwexjlHqRcDf1p6p/jBO/FrcCUAaeiu4QVy
O7S/de7r6lMMekeBeSs5jNU8dkLaQQ6AL5NEVebdLY1d2MyfdV9T7p/J4F573BCkFmJO+fErOEb2
pbLLYtftHagTQ5nu47ZTYWyYyk1clhhDh6bDcLp7qCgZuoXkyZ4SXi/+FP4bJ9Dp/yMgTikhc3pg
0Wkpn5TLn1Y4jrcWj26qMyGA3Y2Lb6SbQPwfPxllOy1X0arHUMBBwYw0gDj8F3sC30bDQWU7zABR
WbfEuHZlF/p+mm2mvkqJRR00W2JfnwRAmst5Na4sJ4iPt8xW5Nloeox9mxmwNoSYQGPg7LPT5J9C
o9gX6lYXZzQjg0GORfo+tZgHrRtGt8U4McG10mueZR78PaW46Mh5CPllve1fNSQRXwexd+2nb+O+
9S3QkxtkNlTnbrRyFvjTy/C0XdzZ74Two1fuTSLKlNOgyEuSn7fT73ytRc1UD4++THalELAPXaSG
zyp4T6xjpEoxG8/KpuNzCoNJwNop/syEx4k1lgLRJtxK9jhE74LbUZXDa4SLHCE2qYtVIlrSOoJL
3ShUHba19aY4RrbL5umOF1l0AyvmBC0btTJ1ss0pGtb1Yg4laQLG1WuohJzK2CNQc798XKD9wnf4
R5AYixHRAb1+zKWZMWKV7flssWS/ySo5qydus/CmLW99GURmHh+xk/hqYmQlhOVMmz/MYEceUxqu
E6iOYSD8FMnexGIiXbcLdbuYQIKZYBDULKIBeWVXNSY0F/mkQoul6ABCL6xaxx4K6VlmaBnhHZP1
HXlCXb2wq3HOakDIoQ1Q3lOAR8uGDjKWTVVa9VmL4GSi2cpiveoqXrnsDtEiBtYaujPv4hfxyn5V
Ig4xkHEuutQW6JECU7soRvMLHwimeyjjAEhlPCtMTpzpEvGZIUK4EdtfP+FpQn6FlKZwJC82+T0P
cDB7ksDQ6CM+CUEXWbChisrD6nqXgP4/rc9MNpw0ded+gZ0ZMwJPAFqFzJqLN/4l4zc5eojg3e5q
6un46cCmmNTp2XKQATO4ZO1ZP3mcILHO80zKH23QlUPVQkMEsEpNHaaRirGHKi57Jyc2wRQ7usgk
xYvQBj/dZM6SGRG7fMC7FWEf0d2MUUYV3sgMhTEEcZs/BGMQPQVqFqTE2rRgGsqyy24kbmKh9xDO
iS2R/VLgpcmrXou3XEqNu7TDWTkblmswgOU19yKXZGqs/DdBCzQmaL2YS4yl/PLp4BFV/+70epVs
sz8DNQ757WJUapNaTp5nXpIlIBJhSBN6cUmO1DH7ewABkT215lo3ulRdUms582+b+J5Mow4kvU+U
ZlKHA8Us6QbNx6W1riolABMnLWfAfjLMPmy6csIwcBZ0VoDHyDV+VB3YNe26jxqvEKzO3QTr/IA7
gd2m91gGDL06S2wOwvF8XBb1sJVq/TaCun7ZvX+b4ki4uYToa75h01N/Be/yTW7K/b34Qe0yqYcm
IeJRQ6odtwu7tS6buivlkj4LdNNaDYPvJeu3z8QkPuLl6Jn8P8sEbjPIPtlev/gx9eih/OqhK5tx
tazLK0SG43UUHhw6po44BPoVqTxFbjhfBNkoh3DlyNf3ayrjyPwrpbwsbaWh/7SbXA5/Vjjv5fAL
sRIaH+SDmDMU3z7UrSlFwpe9uQavd/IM9qvwIGrtg9tmacmOnla8X311DU8u/TwqxwVjx4j74jV1
3k1gvWmy3VZ+p9cxGgKufFdK0rIyLQbFngELCkPVDsmf4aNbnYmTWI3E6y9jHVi+b1VADRcGVWYn
QJIZ5rxCDkrGLL3hDcf2L7BZRRCv0+zbFBUVLuLYgKaAjEs96Yxf1Cph8aQ0Lxifge4xIEEMgSIz
Ag4mC88ut9hf37rZ448IToJQU/w+Fnl2zmr1c7RDJ8pkDLgg1UruaY4fTNcA2YgurqKGB8/W5uFy
6KEOCvZLlmEfdzgt6NNSm5p64T+aJ55nGHhwbdhuhvFEdzd5H7Rlg73kt+wzt660mHVz4H2MtwDq
5vwNUOy5a1xASXSi0x0+TXIdY3YyJXW1vvRnbAZm/feDvhdvNs1mXoehxR3+Mrh+L+GV5kYeI+Wj
L5y/P8tMRCjbxgH0LWj1bPmFmr/kQLHAIfPDP1Bhs91SXuGIXkdQ7wMOuSBU8eTac9eCAxjPzuXc
29Z01Sg370nwNVPYqJsbKSxSIeuv/vwyjLYFtH2VfyXtyO0ljp5qJF3edcgtk8aVBIe/KUlpqWI4
dKo5kPI2WLKKmQ19xwAWNZcg/PQF34DLWVlp10kYX/rTmzkk7aLuZKRqLOSeq2Ga/dvpGdk1M4UW
mXipWH6bnVeTxglrMoSnZHF+GOjOjuPwFcmEeyNhRZt0SgJBnWlhaxLyfqV2B0zX7aSxU3JQL65z
nqPrnX2d4mQ3OpECNDKThguN6l0gbqDdOPAecA99t61klmIll7szeynABoNPf00hZtyW6bh2LWRf
4bHUadqBz/7MCSf2G2AYXEB6rsVQwKKOsmqZxXvOJNO84eaDYlhr1ws7e/h8Vpm04YYoUEuIZ7yW
VB5vaCEiuyN83HSmuGX7/RAhUQsTsJGVGt5OfIWfAs98BuINGwu0DsNB4aGV+Q8zPc1PppLpW9xC
8Pb/zjbc5egSCDomipwVXRodbWNx+csrXRGnQI48uRpvrKKaZUr9ASysBh8rJphN9z0tfDvNCPml
ehtoBQI+53iJYpyRGs85JhhHCJNroHaDHnSgUcSSszmWZW/b9nh48qD9vhk8JznEiWdlLDaIE05m
5HDrXsYhocqv0MGxI5+sKYmZUoexK+IdRNcwDf3vgXs9Dug8TfYG1OhOALM7N1wfjXConEB4gTeQ
cjLCp/M3ZhCIraYotC1LoXkR5m+RPilt/XeI7z5UaP1zt/ePzVAbenGC1Uk54paGhtdz6ftHnow0
aoX612DgOW6Nd7ntVJsItEAxpU8zekDTDKaNwAp7FQWczhEvmr6xssa7e4RgKeoaYJwYBVgmW0OG
gFlO4lGxzokF50z2BGGtWv1sZnx3YFN8nsADZJvbsHLlpdRf5NK7mTcXR76m0rfehMOxiEmwfvkr
wn24X8PgyeinKjB1BthCcEffyup+iXzZu9S3mGUMjmu/C9xZ9f9MaXqUYMjSk1vHMgVRSY6h6ZLN
9VD/71kRzwODkrVLUSLJVOM5P0qNIT4qJgBo0b4EJz9LhvgdgriwICaiivDo7F/GFPOokEryyo0d
qqwUigc24hIVZ2S96LXe0Ievov67WDI6JN1TNiUmkcxFwkHk1x0wZcJ6cRW0Dzb0kJiv6KopJcxe
yTZ+nLi1S1JBBCW8a5wGhEaba9bZYgHF5+GUHL2GuzHMLsbnnzqNfOG5u4cDhW9jqESHB5u6lxYE
wWdOa91mueThYQ2QgXmYDAXW76HKYCf1m0mVpfHEel5n/AU/G3q2nyUqZ2EHqLrmDdSiLmjqc7Da
wMsvb66FgHqIfqcfPILvfLSUzA9cpGygTOsUgMAS1MARsKE/4GzGpCCcafCW7tuw1CesfupJ4qws
fL0X4LsUNeAL3GHJap+AFULMaGsxmmdN1KEILcXb1ImgL7ifFNQcxG9wdRUIOgx67xX7hsPio+yJ
bnQrUAeoilONy0KlmhkzchhmpSqraVAfsLVb7K8izw1Vre+ZwdH1NpIqf6EL2zCahpGTUdPR5lYB
Co12UmBOExHMLoQ8GbkngEYVeX05wIxsbVkCL87nJKdO738H+CfJ9bPvyzL0yItVzm+jrokmPJn5
OLLKfZ5nP43/s7HfkAh9kv16MVyr+ca7syo3yjQmKVcy+0geWGwpNbPd9f6dzglqwMTXAXPbUgAy
Ew3T++ofrbRzC9yWUi3X6nam5rRVnempoF/LnWv9PBbig/7ZZs/WySDJsi0tHz64ORXDiXEuWZLP
NQVG2OEPn9aKrZ+qgvXrvY+s/4QlLsrMFqn3eqFOLLkZnD0DQAzcqCEEEIocGFfcMM0XwjiNipn/
tjTP2a6irYUap1i+V+XHsfPDtP3wyFC+MXW1idmvZ2mLMPySpzCLm+NIWx+ZHdki41uXiUBrHvwZ
iGcpVxOHSNHu5mKFO4gO7j66VB1EqMxV5SYv4IMIKNyLEyVudLLOI5qZtmnAlbGDO/uAfSHatsDk
ma7ptgaeFKKN1vnREd5nu+/v3d+Wi4QnNb2ImWb7pmqWGz1/U3IkXKLy+TI41sDVncwc65HeWOal
PJeeKXPz68nPGJgc/t7QYNuIDGQ6A/opECJlasZ/Q+/ZXHe1UDxCOmQFLLQZyYE5G+sYGNeSG5Fw
yEDbFmkPvE5GXsV9+bWvSLbPH+2Cw3hNIOCqJrId1jJc1CPg8r4pmIlDhFMhswQPNlvvLUcAvFwR
Nur6lUzMGxVEeeE2hsrTNNvywVy3DwwR/IoegHX+nZM+dkt821QIqdB96NO8Ux7ZhB+Z0yrWX5ek
2noqXsVX5gSeV+5FoGF7B7Ja7OncJLWbIooR3I00JCodeMgNhN+1ocdZ6Ky42qff3jHb5Y07vzfj
6iC1gK4FhiGMaX8RurkTnC7DYT5A/mN8/BqlX3unDi6w1n8AIwgozeYWK95oXSmH/Zx1FtADt/w2
ljAqn8+3lKAgUZqZgYswZNmICPNunWsAAoEE2qLh1U4WmrC8283aq5D+KLJw3eSBVOMF9WBGJe4c
giVM9EMSQa/txbuOp3cD01Ca/tHPnz2DGmDI1YChyj8hL02ED/G9uFckA0++e4Jlc/YLjSps75lS
2ZyT/atMI4RS43mD7DHM6/RW2iI7yrETVHj9Hdrgr6qSW4+/tLhIMP4qwPTBE5gJXWo7iUY/dhMa
ayQ05ihysuLTtbhHuh7Nfh+wVxv1ne80TK2uMhiOMAl/JdD55j0ao80lJyXFOfIm1KeHirYxr84Q
5oR9yucJNMhhC3Qa+2mD17ydmKSZVueqWqyuo6LvCGqyclM4PPN7QnL+ly7j0zQNApX45dwHUzFi
0SYNIMsx3oXM4SbEycAB0YitaGCWdWQ+uIfYq0rpbJ60ahHUBIOF73ofCuqTE+SMfrcCEUmO7rRD
wjgnFC9noVlsXh5VniR7WwDjew0A46F2y/0dRCPrAmQBT9Hb/v5mjXY+4UyjWEH+Zk1vmH5MAhwU
TX9g91jxDXYCBY8c+1kN5gusMQen+D0r7heNskcuAZaLTvTdoPD9BFeZqFtiXrvtvjHJChsnvW2w
c4s83Uou4IwXzTbLU/Yew+NEwAE2y+S6fA+3ZXPD+QceFTPRrjdlnF1tboa4pmID35Qtwhk0kTho
+vyb4BYQQ9ElCcmqCwEDVZNcsTr1VLDv8BE3i37pwpT/aaaPuh5bgCNRzhPNO6rGi+pU3lIzyroW
bCnja1oUkK9Ixy4dHfbvJxi0tU48egOR42fzspUHHRBcRMCIcQBmZaCpb7YpQrxUcC0D3AWQONX5
78nPPmRXZEF80lSYtR+WlUtUZSHy0So8aQ1LsCFD/3zPsRdRfkWYVVKT2kZ/fQ45EgP/nnRaGbwQ
TKJqrPVO6D5+EqPsry78Aj3A+/o83VLP9jY/z87/ScdVBxImGGXPx7GQO9XBib4awGQ80hPniylS
GvGQMdQa4X1tfjBYDWLHQSqb9oYtLSxfK+aii3oK/ObsnNk5GOT5LwhRNFSMaFtMOy/Wqr6md3CF
9Pol5ZuxWJ/k3XeEFslsL9xJnDraA888Es2ol3SvtHaakq9F6Mfqvp9ENo4hVaOSGTqEN0TEwBTA
mEWL/uJSEGZdKOMec9QS4ejyfKspdEd5koMF5BymlTjFyrKv6EQnywgjjqIfeOD/+KNj3Bi+t2GP
uiGVuCGGVGuef3ADAv8btjbzZg20ji3Idt4Ckj30ONcmNqFYsdQB6gAiYu5K3jYzkBYM8X/qEEaX
H1wQr0Rw9h0hjvM54nNruPNhgPeCkNjbh3WaHfehmQeJMPp1U5E2zgEgfmed+YZX7LU9V6TiVzgi
mh4IZkUV5qYRE1GIK8lsaXtbTKy9IybvVJGwToA/eeHTvrhrHUsgv7dsGKu7mlFpWDcYFKWpQ1tf
PXJ7e73JstwC7OgsqnKn0nQvs3VcgiRReQumIxrb8pEuaYnVIbLkDLLCpNHoXk16PSbRNr0qjOmI
7Pcic2GVW/nE6KAi4LogRN2w8pOay/UyCiKazmf3QwFW7oIB5nvUYFStbMNM4p53hqBYRcG/NtmY
zh0d5bWCgQN8904c2Wy0m9+tQqjBM6yQleTMe28aekuKilVBDXN9FHBDa0VIUv7mI8OHo1D+cv9P
nqag0LbBJrudDkIqVzLKBPWMlkDjxkPEHtnzd3uo0KzeHtnnlH4aGcEYYVBJ3WXlMwYExGovK1+4
s4ohadBgd78eZk7d15EnVJI9woMvJDuAXk7ooTpPE2oaG0peT3rt9U2CQmlItbYmdVkXXQzazPw5
83D+XQGCuAD/TA6O2bCJJdPoF4L+RPqqoYk+9vUWsfwevTIJXbw3VQFPgaqoIVQ0bm9K+rwcQNgM
Z/0aiF1cMCQC1k4K2/tZqS6ZmqWLdAXSxQfltpdaDrwf918vWFBjrQGxnxIptVGFLICTdP1KKMBw
Sa9XHbuKJJpEgyRp0ggu2OQnwnmk6g+bEy0I9iYm2JKX7cr0vPFzFIOQGZAw2m/WOK9zVRbAkqog
ev+3JawFZXgPvqDtW7WNJzxFK07IS6GBHTpUixLD3tUZyP0EM4lHqRTQO+cbjXW+NaJZgIcwUI0D
gJNN3zNFxXEJJ7NCsfR1SpeelU5GgpBiV1fgjRLDB9tuemeCq8GyGu99eldPCbv19B6rW8zTXPFH
Q7s3ocA2iW430R+st24WuO6LrEm+LEquXzanejvzpeM/uo4/8aAzvn9YZCnMb6OBY1zvCbD+gIXh
2ofIpuduTBoTNvWcWvTuW44K39A3mdhumRlMuKklczHVzh8A+ALFVIwBLvSZbcogLabZgWQmVTWL
Tc27m/Lo2ooz50R3EGbXF4AUkMcVPp+F8IGyygA53fQ97uSOebiPSklDqreBpO+zNy4wGsxBY/3S
/TSaIDoaOHSzsuPqyYTsU+rxt1eoZ0Q4+fyA1hZzUWrqeoD5FXEPzEtDt268flicUGZmd39ZQC8a
O02Mo3dgwHvRKqOfrBDMBatWSPRseOmn8s3gUfbIf2fgBwl5nhczsUxaWbJY+PL+2NtGKlJcrubb
jXt2q6KPHhkvTJbjwLay5OX+fHrUbxFggFqJiMkrPq/vjkMNOiNObcWPGeMwpX8VzhENXOWhc7V+
vCkwLX7J8D7LJ/usyhyLdylANvvLZHxOwGRww8MrUGkZ3aFZPsLmlpA/8VhidhS+U20bd2rFSpJl
MIQ3zAfKbE9W5AwiZ4GO5KC5jmXWM2jJTEpW4R/NfVkcTVnrAj68OT9qdH2zpLKj0X+gDm/rvzJZ
S+WnsfW5skA4WGG/aBYqIOTmeE+7uVx5QJT+MhEaI5etpmy7egupwhTtDg8HOPxQQv42WcVrWvvm
Ni8ShkzW5OIL1aXWE2SHtl645HpDX4ugV/qTOBecHCaJTvptRuPJHwm8YtdnsBfAaKIy9yycLurF
Bu9F+yoIBL+owMOj6NOZLcHZfyP6F+HG48juJqe94q2FWEJXSWH+MoiuY0wssJJ5MdmpsWSRaUnq
Xm/h8ui5ojUycyJYGMsFcZ5os5ztVbTH7Lo8jLPiYk0NW8X34aZa1yJJ/O3zVSbDYjEFAnNjiMLm
QY/8GDQ46qhyie4dVIJ46wRxRc9syMN9Tv+EM2noYrSe64xyoLJcC8kuxaF3MfppXAg9dRwBlcx6
qXKU9/gonEaa9ZCwqw8slPpzm3ZTi5AbpoBTl/l7Htrd3Jm/nfPU0BBZDyzzt191NzbMCSuUs3xJ
MD44I090+OjJVBmb2m0fWkCBo6M85pd79V3QWi31XnlzcoHJYsJQVIaz6fTGQ3rXa3DqEMVEGGcb
a/JqtOTtqHtEgATNCyMHgDA4xncajp6kKw2+XOIdNB/IIt/Ks3KPlDUba+SYdicOl9Fl8f79d/QJ
egx+w6kqZL6wSSvzGX1PPOCtUyJgxLf+LjvKDYOl4vOzqWBY7VyIze1jYhiu8IQwq4CxMW1DtUMt
XiC3Bsc2FEgZKmtjWUYL+I1NtLzBfHm2H+ybxRFj+omsJphOzClMBq6bPgP+7u7pswTrv7UZt0S4
j48icrkZXwq/FBsz2ISPMzaizv2IkgSGcCoOJ5cWTL7iyMB9OepJcj89qO6fSDFkOJ61WSjELIF8
J+AO9dF15U6sBa/33FbHImKP8cp/kXAgXpl37K8ZzFM+SbQSLGgc4QtEgy+N5r1gaQwiGjLIJAa8
4TonK1ko8xcEtxaLM7QLL2q8USP84h+fcsQrdnWU37r+b4R1V/2RWqDzhH4w1L6x0kDI8jZDRhKP
CEgRhWxN4n7ZPqKor0LyUQc4cckEAgJuJ76lChaNfkjI5cqSgfOoNrwehPKS5oY4eUzBI8jeDq7t
+KwAckhYHrOr4GCfFauQ7c0AjnyYROLAU9MUIFZHZGOzcBL5+UEAruzc9LRx6ea/PEcFs1a1T8Sk
gE9G8ttfG9vap975YvORIIXoppZOzi0fPZo3lQMimEO8ZgPZ9h+juDHqN6rUe7Fj0cmNBJ/3rgIa
XuqpQ/whJzhh0kXu0J4ycXSXnKdZZDX/bZxucVckth6cC7doDzWBP2RKhVh3ouRr64uV7GXj46fb
WAz7y2HR1V6Ffmd+HYLiaIw+Dtl0k8Z1BRKnJB2AFOLdhzAwDg+l0AS+QgM7z2NC3X+42Vdo8JPL
7m6e8p0KfzASUb7b86b8d5d4Cce3XAcKchjOfI8UJ7EFw1LpmH7UAz3c6vAnk7lin4DbY4IweRdy
uXZ+US7M3HQw04Ri5JX7GrswYduisTjD/x2ABTKrju3edyoAZjW7C4qMjDDbVGBGx90GMOMTGtwE
nxT30deWQ0hInJnxL2JWZLEPP/K70vwgjLDqAB58QLIt0MPAxJ6XW0E4yxaV+1QWuG9v1poEpakV
GOFPF4KqQqZSd9cK3OTX433hstW7s1lVzAAjoJ4j1TU0BCuAgQXEJrGpbvP11QyEfCzK4/ZIvPtf
J//jHawYF5bYLbHVj1TZzqtxBLbIJRtdPMUNvo+ci7Z51ekrrvvtsKUxqmYd3HGoswNW9NA0Mpzi
nKfTBvwEonSFr9OxrDdPNJQcZErXF+2Q1hOVDcwxC2QCLdADatrv35ceoQw6VjT/9pvykO4Varry
NYmwp2KLEpIMsmnU92zBwonGqTlS/L+JfV07JGOG45kPqTFXH8w4jnQCyz1C5Bugjk6yldFrzJ2J
l6TnfDcr0PKZXTBXdBzWqo6tz+v+fMIz5OXXYYFLCqAWECWAI8elNpstFQKVV6ZZ6V+8kVCrre0I
Y+HsA6fbLwRK2f8yAyAnoNkW3j6zRH4/vvw8eeliPKpqqe8dcZVJ1XCN6o+xeWE+tn/uc7ix4siE
gY52j0XL4XpmI0Yxn0Bsr4dT4BUjA7bB00zt950y/j7SmylfcG54s5lzumqgQZiGzAnbONGI2VDc
BQv8U+TMDZSrXThMoWYYBFOll2vt52K/6DoRTHQqKGlYcBhQhBc9Apggtc/6BL3X69VcbSB7EVfD
KTwe9f9A8VrxeCALWf7VcQoTNUiYPAMLp9j3PilGQE7fRUdtlTEsBSsGMHK4R3HIDisOvyAYE73T
FgCFvtjc8McCjIVo/DiC4E4C3YnQF8dyesJA35K5e87sKa+HXfYoqkeiLXtcxQvU9wmQ5nJgJLtz
dSG+6nPi9Pha6DXaRiC5aZ38bAUy/38aUy3v4+oBA7VA5eFuGeQSvlBvvuhnATGDrDnVZFCKcXFx
zoB8Yms594Ehdar3dCLcMwM5z3xNL0whX7j5FaRXRcOwjygGCroBcEu3+qONPdM08phtqVMKwsq9
xhoXIhRhR46u7jqHNPI+VdtRywG8lgtIk87UmA7ZtAK82L6lZAomGesasbK0CgC/A+5b4QKD7I1I
seqr0NI/kLkf/x1oL9CDlV3yYxqF3VEUI7dHiybO2askUQUXPjsXdHTEsiIJrhQNP4rPFPqEDrNI
7UshK3LobTf4ZH9MbotW5c6OBuWfJRpvLAssnYNlLGdGG79foahlvHOnyjvZCqPpGsgEMCu5zDnS
3bMPBLsBhBBYZe7VhXKA1PGxzxpCrqR74MQdTaTeUZLZUdAfBgmR768Q/GEzx3gzIvLVCplPwmHd
XtQL63w4MKqsx8VsNYrVLtaUJ2/7u9B0sUPamocC/+1YTfMGfU7g4MGV45JXnr4hMUqSwXmLfgY0
vtr7wsaVW7KQXanpAHPU9Vj9dJO1tvdfpItdR5o2pIhvuxOPSxoP+1zA68U8pDINAvVQbgbBbBlf
sBpwKrT546rz4f30r5r3n7qePfbF6LT83WOCtSIdmESyhQcBrSGYt85b2aRURJaF/1oH+GBnk5G4
OGCM2jEqFHJ7mA5QSICvSvh8ZxlpT1hTyUXLGhb5Rp91+RhyHPJmiGz09W5cTETVRZeanfFicJOd
MBGUgwy6Hn2hZclE7xgOgBSsZTMrN5KaOAhelYgcYs303L9+WL+ataWw1B3AzM6u1QYAcoJzyRMi
WDxOQEzau8gBV6aoPu/hL2RBl6nanQVMPNFik/SrITrY3YO/U2JDS0JrRosuIMoNVMCCr+FdiDsn
ZcwOT7y/QDd9WQxYvyO6Cg5rqLg1jZpAMUOwm6BOl6A3M/R6s0JMGsA/dScp6eH7bupCuB+l+Sxj
N3IHsrl1ssQbsade9OVKbnyaDRQilsDmZp1xoS69vGMrWIweJv3DEyhK9goKcOjIZlaHbyZGOaxR
gkSL/Tp0jeocpwz4whHZBvp7fbmo0fuHKcqrAW12eQPDe7KXN9+dJderzyFHTh9dvlzFKLR69181
W9y05GSAy5u/GnjaQ4LyZkTYgzSY/QB764s1uQkdZZfuXxOYDJoYGdNqdd2EVXylCtmqDE3ADffQ
yM6YHzwYS/QJkvnjmiEq5TgsLQy9J45rmpqV6gOwzeVlz0ssAp3FS6mlTyrocJFP66Hze3qMQ3s8
3gXv9IJZNrg7IMv3eCA/CKKKqpqtfksqTckNAGZ4TqxypfM2O5n36a1SHnUCkEb5teiKmBp7VxmR
V78Xpehhh3gEms1GoBwGYGmKvqHdfCTUrqy1JFx3O5xhFpkAHsBAkg/R5NuHdGbjW4yw398G4/DK
Wid5W/ejRs3ewBFzEmzYAJvaeipWocnFijQsCf4SgTaYGdC4nKWUXnxsICvZrBEut5rpoPuElS//
EhzucyqKTgBKnoyiwtFXJUECbsxTz9dHqvWW5sJfsSIXSH/ipGJ0/0AHeCsjn7CrdKFQ3NBPuvr+
9Oo7FUbSY7stt8anrVPySHFM0KIZH+A4fZGDGZvBsauRk74KcED/6KkJeuOPINCUUTR0YBuK/1p+
HgNZbNU8aGrMs8YzoPBH32DzL4lM/MR8LmOH+f6+l7yiulRaSEqzh7ZLYcwmLyXjFIH8VeaJbsnd
b23227iChv/ppoz8k5DABp9RTtfdE5ugy5BvsxpbOXyz8wdrNePw49i5IvKONoVo50WPrZiUYOE4
iz7eyhy5otALZZqD7PCRpzZtHi7IofV/41ehrJzuSOzg5sFHPDEWgcr6IwWtd/hUQcQtCnvm15/+
RIe6RuBzGTHtnzlaXOuOy9R6RYEea2WPHF69vnLTPyMNl/wKDGaNOXXLT9JSQb2Ic9v/Gx2/a/S0
ic/I4E1SNQ/LDWcEoE6kdYme7HEZSOYfWapmfYWfDBcNXhDVncxuRGaYcuYYhU8e9UOxYfabqIZL
qk/mCychEEExcWHnPeAnsmahYYqAYZ/jcZdeDzsWeS13odbZL+FuSHzTA069qBCLsiOiRcEmUV1V
im6hMVr5iMZezZajl/+Umd3GpejfxdxkdqYvkd96qn0FDdRrgldAEriOzcQ+aZ4/oulJig3soPVX
PrYgktJu8qj82GBDgY/9j8g8WMpAzt5rghTfJQTAN6QrG+uoi8tyUEeWwzKuC6n8fMX085ypqWJR
5VA3xiO2NFUE5e114XyBtSnbps3K7TRiqe3SBpAf/imkcWhEl4OQzCXxUiR/mc4iaxhPu6k5/Kw8
kKj93fiBjs4mT6l2CQywU8VoyG5X+aUC3g2Wd6SoRUAktlzsugnC5vPm8yzhUBc2Kp8sdsXOopwP
Gs7C+5m+YwiLmJIPLyJAfAC2mOaXzEs2d3L0NPLcT/YJ5ZDYCHZNiqLjjwo44XCFduAwyEbYz4wu
Z6ippOsCL1UScrQSojwJ1Q7IQUMskJrmpkqm91aLKb+nAi+Q4yJQQOZvmlVrO0frNwf8Zdcve4uX
X0GQhl9RS3ixMmcF8DF9HTeHW9uScXM3Th3xe5VqRviBSvgqiXbrtXlKPcuctUCOLVudbWnYgx7B
PJgGvqwqTjEXwrauX1QKtANAT8w5CtwK0xE47nun4eNl7pmB8C8iDXIZUgLNF9j0GazztGH9tcpu
ukUYPHDt3Mk0JzoLd4HZwQbvjiRMMp/xpmaRwQq+QLT+ixPiWIHbzRC86/zzlDQGl69w8ogIe5Mw
vwFQAet3sa+hpqf3dwV5Uw0alvcDgmIkJNapwWK9yKVn8pgEscJMCXHexerIY3+5uCqmbRcdKwTJ
lJyuZihccBehp0MKFfev7Q5YHw79H+FqyBhXQEbQ10WK3LOyI9rl7FwQ1ThniKczlZDJFQfIaCML
OQIchjYO4xO1KnC2ckDEXmwyeJ584CMUjliLKTxrsACTlEXtjuvwDrdbkYdp2Ghup+PBn/aqLQE2
sv5IvYTTUZp3FZS0SUiNezzEMtyibCbvLS9f2JLKRWobCc3ny2M8paUl2MI47CT34P/9yMe8upyN
ysnLVqPR0psPafrT3My5s1t9Awy4aVNmEJKTkY+bIWJzuf/Acjp+/UltDTNNo0D3iFk83otPeU7+
AMcCRL2DjMDJluD00CBfmPPB4+ypCXxBiZzDEQ+KkD2M7/phnPnBuQL6Hnb0usMU0Asyk+hZoE9V
6KBjFO3lnUDDiYV8F/FIpVl6nY1JyPpNhPdOEKFp40YjCVK9ZjxpvnFY44Fk+XIIovzCu8nayGFC
Vp79apObyATYWCe2B+UmvqbGsG79oNSUkv8xVpSZFuMk1505lew2caT3sLNiCXY9MUHROxif28Li
GmxNSrz/W4Yo66eaHn7J4W+XCnC0Kp/V40hrM4GP7VgMduZxR7Qsf02wKsZ+wMC5NB6VIde4tZW7
CW8MXm8OU+fWC3TDGzCtyUxlj3wpJA6qY4kcShpLSnu8FDRG3mmr89I17kIh5UvHY9/Vxx4Nk+0A
OQHPqNXhqOXrIsQShwBDuVa6CNfi2We3xiB0f1bHjU60l6q2ACndNbbe6QnsOrFPMC3Al38nF2Gq
4Ujx6uojwKv+jAPmckY8HQxr5l7WWtcuI/Dl7r58NWG3EIWRl9EERCdWpWkbt0xchg5usgqkFMhM
AlBpudbwaK42VcdIjg9Gh5d0trK9gMMcZpe5CLJxiz/lvgJf4AxDYvKtalGxhHTdE5jMCSExwLm0
uN4wAe5rUKlNE6BAb0KXckaCnx35qTjM0G1dM5L2RPMuMe1jQBKh+9x1gFH2MOLOzQA6V7TfPRKj
QtGM3mXi9ul7bZnzoM+Ifc0d2IHKJxsoOoY5ni0EeDP3WcCYnGHBQolM0mlFgKIkjhGcKob+au3M
rBprYUFoZ62G8pJ5kRJyBcWdB9SU4xFyBv1iZoExXmTMKkC8Saee43TMvfZTgvlvz9IDUoge72dK
5nqaxcfXJgp61WFkJceIF7fCr3o2yqvR41J2qHXLy/m+X1NYxAm5R7Y0gE5Dd7IbMsxJgMmDfYjZ
Z5fCWqtxzQPvCeBNNQT8mkIRxqKmNYjQpeMNFOgKcnE4OjEz7GNGEni3CBSVQOAc06tqVmMZ2bIp
6krrj3AEtx/7eNzWtJqHXqdIoLz0pzDttYCFS3uHFWRtoNmb5nFMwD1AH7jLUIQdoJOUhQ8CIDsL
ICLCSWGiWR3TY2/4DoaOWCi0t+U+FPEPrxA70qYaq6hWXAEfMsEOXpjhVaEX34zEcJswjJcpibH9
1dzt/4SIwBSC0uthQECx9Wq947mn0NdTJejnPfrMrccolFLq0iZhk7xIV8JBc79SBFisJuq7Bv2D
728wI0steGKSpD4W2lP0aUtSFhb0oJUYjYXgFUkOryZbFhqRLYGrKEMx7nay4qSnL7+SRmrOBvmg
np+Mk0+ZGQg0UpWCEMaJB4fXwZPdqPuGJapuL3C9SGw0qLM/v8of4Zm6rn9OKm1PPoSyjQkMn5vR
D9CfmFlS2ScMcQKcbsU/PZxwVR0nvkIvydMJUOFDq+pf9TKtPzIU43bn+Se3Ql+WJWPkjwcnxRZl
AFmU2QjnxDMqY7yecDWtj/FFNJN78gx14UozteV5n8fywOd3agag/QdrlwRGwjZAixPq37TV6g+l
cOFMTuHSxuzG0W4NcMk/6aoRLETWi6a2N2STs21meroomJcHVNBuaQhdP93r+c2giaytuE5fMNNj
Jn9wTMBoU6+F/auz4lQ+Vy9exqs/yaF7sxSxXgzGTR/2JjmRSoiOXUGPlWHEnem3otU+UfXhKBYB
xRH7x4v4q3FAL+eVzWKT7IxQLhW6xzj47ZXARZEntgk1tTgAdfnsF3IVWNbAQS531yD3qfviFHhy
P9OtDEVQ95W8Updd0W46aTSIzXs5La3ALcNrMXeDeucmDDlKERQQf/es7J73EoI9KOy7H9mlkDYB
mjXqo91Y4SCnxIbYUI7X7Ah2fXJZRZNq9E6LKbJb8qFQ0XtTjqbT3wZ3GXI7cyt+iY3iGBjBmtrv
0cPwzcjdYyxR507azNW2rroWVpVQ6KqTX4k4D9Hm11kS4IwjvmNpWxnGUiQrHXd6utubIQLuiHt0
evLpcvp7lnvEiTGAZELdnmf/uYWk3csuuXBXb/OviexVRdGW3c9pFXuDOMm7E4GZs6TaaRkNr7hY
dczvR6a6Bo3w1RXPRGrDDuMyXwzXGbi9c04ELGtWYtud/i+Kgh3qucE/xlhiFuBANZvgvUyc1FqI
X9HZwCyPVEvlhiWGO9Dua9UXEbcDLYTcSj9PCNOeLsADbZC67xFBPYrpftHVJSLWtvBbNySWwwMY
/IOBsH/CosHZdsIf/TDuPuuaWOObhXN5yfae8WDqidDl2DMfPBHVRQ6vgubwXk/H4EAhdL7SKNmK
+Vz7/7aj5bzqInGZxOFjQiDC0CHSr1r1+pRfNMwfz3qjsKijTS7lgDoO4gnHwctCQj9yzmd0uzz4
Vg4vEEWhZ/JS9p96bxfxFWAN1JKc+yOMaf8v+aPXsRrM/uO0qe0zhFFA56MG3SQs8CzeF4n25Z34
GpQ3G16BbYtirvfcy0Mqtye+dZZM3ISVoE1NRYryBDuiXdUKS1tohXUvenrifRABrDIQbnhkgS90
HU20HL/pglYHcVlB7JAqRT4sValbGXrEoZRrtiQbPd6JIMXa5MqBclgv9M4EHymXQZNZYuUzYnDF
LqqhDo4Jw08+vGw5HH2kQsWP4P1Z3IagLmaU3FtH3OMkkI18t/T5ZqjdZ2nylI+lRzs8XQICBwp5
X2t04vRO2wsErzzkKOrcflPUfUygaaDAI6GcUMWaD/ZVZ/79sVV2o+F19X8jmP3RHmHHrJgwCSly
6p27SkCTKdFDEpq5bZrDul8oVBei8zaFB003Ge4xbdNymhOxQLVyCJvDH26Hj94t9bjfP+lBtRi7
kK5aL8RLsv1rkeJ9cwg3qZ7VuDbcHUhBI4KohsOOcgMUEhkdpfV7bWE3jVnPdo4lGpJhoVht7FIT
muHVV5AdKRiPPF2US9u1O+xJ+KHoqaQoRunayHUFX9woWEzQ0rD9tnDF5zeT3xY36Vu6XSPBZ6ej
gc0hfiwi8W6MTAEnugZRPr2qUgDP406L3NHYMoiYoI5PaRmptjdA7pgPALWBIWHCiIubnhLFEJ2p
Rg40khQbZ6JPrSA37zauurH9o9ECDwvCoWcEUaVWbgJVQE4G7ojFLxwa8Z6HnPOujTPFIk98GvLa
FxSHNQOB0HHjlD9rLFqEwMeGu0nb0NNfTOSdwO2xCyMJVqojqFUYVouMMpnEOBaydcrmE1yIXIfg
ArUk1hqlSJsNFrBweiXkFElU09bSwShPsuDkKlfljhgvis6DL1TT2hQ0PEf/C3gZX20fg99m3MOV
jNBmZKbBwWJqJosarHMnQr0Mu/2sK9OEsnTL0ugrTaDrmG8L6cp3dec/uUSOCao2cdBI5h/30P38
/b3gXa/yplY45uOgraX/tQj+f1hgvga3ZMe5pP9VyGR7wUsU64spZbfPFcQqTaxNtAre5x9m9+WH
HsIn8ybviRKz+lR2l95v47xlEV4LdOK/3oaGU5zJ/lo9wgxUKmiKE8Xn7GYz9k+ms1IKsQ81tpy/
EWdmaFLG8IfMi4DVCAlwFXOl30DDGFPbcFkWD0ILW5U1b1xd3OIgIA+4bDYdbmeUdiE8TNK3EJqr
p2ULeIlBxVt/b0VIX9BKfYcHY55Lj4kr8F4jJMPxosOez0d/1dOrhuHLRRDCksXQ9C2yMhs9AG6c
iOZXyqEIGWgxUMIEBPrIwCONIn5BsKxFVGyk9PFpwEGdipo7IAzVDYchuZ38PY8njkdwLgXP+seN
f6VHfb+lD758k/+/iN/J6T0e/d6x9z07di6lkRYQsMrO6uEbn0emXl5q4N5bPYzn/OfouXBU6Sn2
IirVODxWh0cS9WLxzMb+DRyWzsEOEsEaZOR7rTQRNBcw5569CgO32tZ4By1S2zQqRqFARQUNQ/Hs
xG96QEgZBhb+QTmGp+g23k8ePpsBFTRkg9ln5wfuazqA5PX/+1BsXX3uLLpG1WhRKOX86plHIEWG
Mgz3sxaD+463Fs+iuxAetQiFvQTWVCwPlH0nvX3pn6GySyQOfDerNWljouZvouJnJXo4KNACndol
ZyASt9vMT/49girR89qQYqJs99v5BlD62KXElz1uhVJQ+qCTM++i8Uc02dhfkVm1I7GcxRVK2mX4
6pZqJF4zpqg7XKYEzM9CUx5JLy+dGOdX43kysyGyBp/Eb/nwK0J9jDkj2mvpY9yTLIEYDUKJcl4i
tBPG01XbRkTGgbLNtMIiTygSJCnfPa6/cFhS0G1Iui9DqYB2IVYi0/5rfrEnrBcwKOAeJ5/lRmh5
drj+gFw+CSxS0TRF5dj25ZtC3WLIU2lYO9LZ7QhL5yO96TaKUt2H3ga/c3TFKIabkB1cGYrLaNTL
ceZZU9Upsm7WACUkjNftQkAOjS4h9CKQfWuMSTxGdCG0RfauxQicAT2k/kPEDbn6NPnTtGqgTHox
12TrvGUjX/Y8EsqFH3omSskVp8sGVNtp9NLCpbQEtl2f96NtG7OSKC2uhSPptudo2/U4s+N0EdVx
S7wrWBbCJM4vPguEFtFCfqrDW/g0ogi5T/L7q/ULdrc1bN92+XInavXmhxY6Gn17t6WOLc/Ltk1m
S9glPQddOIuN7AZTNPJhXHzyFFGXTpB31sIxfAZEHSTTsLcQB3S2RKYK7w8fj3jfXWtafivSVjOG
4Ze0rl+2D+GIw4YzcmgUfuj9wjoRytD7Ebw6jdPajDUjcn6qGkbVXs3Zz9QyepNxreJmFb0l2Atu
HNvkBRE8eIxwBnhe7mB61dn+oBtI1AzoIl4E81TiFwVc5YoNGGCRvN38IHIQfB9O34b/JHD81si4
OyijQFFb3Esp62I6Uxp1XcaS9ervm+tyxFTEbiWzh8CE7ZF3qAZTDEVPGq5/Pldw6a1H9k4jzPGa
Y2t6Jxc0/dzfJWNUfOpPro+WtM0MjImE2iUWRLv0Ue3Put3ltA1SF8IO8gNJnxvVgFXGwiz6V9qn
uQpgF/+D9e83KX7vpN2byZsoRB8lMWrfTm7dcTsO+Nt2x9jwYCcc7Rxd1mfXEu7g+NAEBtbJgSJq
QUpvLHXO3aD6Lzd6Vr8AlS3OH7EWXyqBH1DD4IXVMzqua1hmoYREvgGiSSUcbdqrdmUCEb4q86sO
0wG4/ZcO5aJnwgPew2WUI4WeBrUSHkuq2TcYky4LivXIAqhtYVOvutSDezSXuoxDxzqmRLmBIFTh
ISFIvqzElZ6+jngknjlZns20uHAvIIoF4AzGdsFAkE7lKfR2MO3bv4mG4jVJSWyortYuGIZiede2
yNNptqv96Jm5wz0Xdfjeg2DOF6FEAwJa702C3l6TOSjAi5lvImEfhz3CW6C+WK1u3N58TnJQS36+
Hcv6Slpl9r2WplmF+Xcw0cYAferoDNe44RplpxfZe1Mzd8WEog9vCP0Ph1csI35Uzy1bsKi/+DQW
5XyBnOKjP3Tg1LxR3FCsnYrOFZ7gRuaJmdbKmN4heZg0zq017l+3Dv1qE8x6aUndD5QpuHrmYKWa
TzoEcmsbQI2Wfs8+IOqtE//KZHUBadcPWRR7KfCiZmn/V/SfHoDzI5RZ4j/XiQOqsSV/vlxkVqng
LLCQX2QSzllDCaXSagQk2jw9id8mcxO2bMagcQep9g06Bdfsb2GsDVP21MXc8EkZq40broK2TmKr
r+aDGYtCGFiEaL0w/mUhlbX+hMvtEyKPzW1Gztu+TBS/+18q8W83/e2EDLOy9TV5NXOU4oNPx+lq
5X001ldRGVt8FKD91k++ylbwtHjNWttQGOtoA8Iaa3iuSN1HF7gI7emYGB1lkWptdrjp80B8MNSZ
FKs2qrrCwIWXVwfr4NKH7GGn52FSRlkAUNAmAx/jp3SDGqIuW+Tkz1/aTlv4hWTUgPLqxTMzWMqU
bMNFSwzr6VflXYDpmj+IvCEqF9zJviRC+e6ZCyqc6qEcWbbq8QYjwtcIknLLY8cGZjKloU3tUiIz
BXmUWCuvRY2LgY6JqKtkIqEfPwxn88g3da5HblOyEZxkd1HpTKc3kVquBXnigfP101hguv2iQJ0U
D21496KFMt6yauH2Rh+X6M3KfqlPlOmuGs89cYPbHLMN+PuG9vHv4NlEA+FE1lnINl7m+ZX1wX1h
X1OJ0/COTLxB9cgYEgGkOhAdxp5WjN9CslkBZcO4WYt7WHlYP/hJ6RBDWEVlANZnfL1tr+34yAcZ
BNVHpLH9KEPGwQNoxgtkCqNLUMLYYPmQIBBCvMpAhNq0MtHZ9668ECl01zSnwN1uuH+OUUVdi3HF
rlAohWlPmChqiTmFbKo2uIIJJKjQPnSRI0laiUJ34x07P2DYM8Upz9seCIxZ1yEkxxf7sFoYjfX/
TJTVtPSANgzN2AZMgE0I5NakLGHnXk0oDtfgxKpHVyq2YrbL1vKwaBNXT5xJg9eo/TXHunPU61/O
Xfn13a38WeDZvf61yk2O6fFqMJ3X0MmxBXhqkBTkn98MV9amgKj5aDt4pCyi+xLrNvYdPwGD3KaY
2FvhHrJ32Ro4O0Dibptnfqz0J2XNwwmpu/duw4/G/JlxV8FwxkKYldDsAHwmhyxz8mBoe4fWSXIu
w2/DBz4jJPX7R4yTlWTeKRyG/nyBLG6d60Ew/fVGSqpIjQrCElHR5wa8/OmFItEoe1nzAYWf3L73
bf3tTvVKxHQ6xKi2inCszYZeZwPhmde5fXnpKMYtAhkowuQC+2GlOKnOSPqq4ADn/aFghcJDCF7O
VTROoR9/ImJv1nu0AhURidO4Z8vsrIRXqsH1kLbZb02YTg7uv2DOh0wTY51ZLkM5oahb+vrEUIsF
V8Cyr7C98cRJ/qWU5ec71h5ipL4vnRWfWpihGSnvQiOvcwvhvEHWmXJz/bi4ZfJrP1I2kH/Wt8/L
l25NEjOC+5CyrR5mKwxIX5ohlAqgdAj8zHgWFihJ7xQsaaXy1jARCNVvz8QK7s0McnyEirNuhAZ1
atrOCfaD+LQEPKSfw9gnC+p7aDU0BL4Sxu9t7tgLANFmjjf8DqLjvpC8JC/9YY7/EKnok74OLS8q
yji5sg2XaAC0/EsVYmduR76W1Gj2NprRdmIeWyAz/jOMfDHM9SsAe5MklbvsM3fG2dP1HrPjjI+r
7A3gQJgbTxkGApEp+/v0YvaGr2OOUgwui0zLMin73VePZj0yi7KxblnVJ7MtMivG3VL4OFIQ5JeP
JZlTylW0lLO2UmdcEc+sql9nNLmkgJXbUjuipegp/oj+3NoZC3dQVic59LH2M/+NZdeF+s1SgYPJ
gLArxIgWsjPNMgEMeW3Vn5kx5tEIS5WJEZm3r1I3eQTbCresZt9HyXckkM2/v/VaV/5Qsnpdb0d/
mzwhq9EjznZlP4KRzYBBuxG1ikdi2hltIndr4kvAZk4Yf5VDVWBbBrklRxH+IuGzlLW2DYNgTgKD
wPDACc17LLdsHNGWSmV0D7X9u83qLLzjLwF5MhI7mocmM+liRyZyibj90ssBWCBlOsju/UEqFQ0j
t5RMUeTqgIKohUvRAoswj0Q4C5oHNVjm1SPx/RR9Wgd4647IrKaeWSMEZErfyfpLTJmCEXLefwQl
3psAF1/NGwBtSS+myuX9OdawOeI5wMVw9kssrkIl7bvPyDEeI8l3EVXy5Lqaex+n+OjNR1h4xf32
vPnVWRHTTNjwyrVsbfd23iaAHdr1w3K4eFxQi67HlOGHZiMDyqLHAG0ysujD54gN1BpDvqxuhbRc
y2ojalgN7CjlJYvzl9BsVkdpAFYeCSI7N9Ap642uoe6FRmfTUKk8sIHKMiq4qMbph3EzjyZ5MAD3
tyLmxBAJMkxsHuekw9hNvBWz1vukHRHxx0SYhij3WcL7crUdn+YKGGLleSKH7V6n3T233wJNpL6x
bE4Sk5vOJ63fXijlHp8gttnDD9zxJjc70roBXG8dv3oO1yWpeaO9MwUS6KXGg96iYxxxlTs9aL1K
MuPnFmI7UK/8ZxA6uFGX+qD3wU8ou5Lz0PoU45rX5jfhY9hP1oR3oDAT4cO3QCffwxyxQUn+8j6V
DKZZQpOctm8FGd2gu15yqx+fvNB9FUSCv5N4zReksyLFhLPAjFyGCGkwC84fR6VUik6oRrEW5jDE
G0KEf2bSexKPEJWmgMHBXlLr/zSk9xtco1Hlg/gbw/skjXCuUZXukIMIa8OdfZOxe12ezbYyCoRC
2JpcFwlrgg0DaYLiGBwy0uPIei3ye+F3X5RUGoVYYaJIBLxZ08gpphP/C6mihEUBTU/6X/9aGnzN
dsyBDbsO6knFU+VWkbnKeMkMgWj24EQ0ZC8Cf3LeyPZxC9BXYnlKPO0Yq/EJeTSNddSu2Ob55hto
5zrdL4Rv2GV2+9tQPAHOpBbFi7k1d8cRhSCNCzb/ZS8VZwdR3D0hKtwwads9ZOsr4qj5XSDyah+o
/0shnz6m4jOgGoPBX9psPFu2wm5SipvWXJ+yVMwu4hLVzFCmez5Z1+9QA2spX3gmBPGqcN9nkpuQ
S3SJE6neojoyUMMtFNfjN9q1HXmTisWHkHWpCs4Ta+XgFiZsM585+hIc0sWOp13Y16yXNjGYmJtS
2wgJ9dHpmVGDLalh9UhBxBvCeTOgpZDlCCa6gQhH4hXEV38sYPgzcgBVlPQjVa7ozeJmmvgN3d4J
xBarEmAq8I36gD8jVs0cho7nDfC41Q5rbpbUIgFBUCE5Guyx8bJxxb28mDVq+GCJCXIZMWfOos6W
bZleuhba3Neoyyk+Gql2PqQur0mct2o/In7IpBRpzBEz+5qfDIoldyGNUMBP1rTOAsres+fVjEvj
DiOlTVCX52jOX9kXzuLArjAVYP8ND2Uh4OkWB6wngbWhtbAPiuT6biM/js34zDnicTOLpxqoYxv+
+KzB6aPJa4fXWG8W3a0QK9tE6IwnQtM9Jjj/1MusYSIBEdk22vMJo4/gXaLhdZpcpw1BoZ4fvIQg
VnHSSWhYhgK0qmfSc33WF2sG89mqHyfEiB1VIQS1FY7Z5KiJEnO/vZJ+jxZaC3QvEToGFvkERHuW
UJBRvDHPvPyHca/fmDDD9me/QgiJMMvtA2SD1Mx81SKnf57ZN1y6tjXw7Cxt5UAQIQmDuujsfTr8
ICcGVMTMHHravW8QCyPQ3Y1JvrHBRfQsYEOT874yAmSqctiRQa2skEFRalNKDEEwg7AWc9uSF25W
YDzd+/iUZbYVeKQF8DfET5QAWTQroziAyg9cgZOUFsTm9REYjjCWyYTk38alU1Y7yvRoAwBudC3p
gx0SyxZrlJoBTMTmAYUWCM9JB/YQzN+1h6eSZ3e3bnwQZ9lFeeWE8ziSJhYr05uj4JpBHrM7FIBa
Ek0aBsEqQM0FjgbG1Wl8MFISSMjPya9UrKalHWpHocUObQi11dMkqhBiDxNy85y8WOJlSEQw3qyV
maqknd2jYv6uixq3U82aCpIox6JSqj3W8aN1wDQblWLeYpt4kS1HEsp+f7c6VS34gHVepLe6pPzA
hVCteUE1NyNMZHRHPnojvqhX4pp9Hqix+UHXnzbaQxtG0vSPIuSqBxq6LCPFraqvrNQ8NEwsUXuB
+N/Azo1uhntnc0oZBz8ztG1Q7q26wfHpJ2E6MnyQnItVvJghSgAzNxlJ9EnmSMx75Rc+Pdkplr9q
Kayb0p/pc1RW3KMWxXkL6+7Ck0FZ2cuWnTcVl3z03G/Ue75Drx8hfiyXJltjY8mXbXNEekQViFUK
fAWGXurvvcsFhAH8eIVr6xxz19pDWEvdXl5fMfivTdRoqCH5j94XBqzDfyEF6xMca5yFXCL4LnzB
l3oRZqxtlReNgaJpE1QGUsUjcDyDsOtfKqqysSH2u4O0lw0XALs1WCT5cIlXmpMVGRZllpqQLirT
9wHu29ed82AEC+easWqPqn6Hvj5jbvBKOhETmA9Tb1bZyuF8UvBVmy0jSypnCqifkgy1QKhFIdTs
PmO2AxQr4Hw1JOYStr58UdEXdKuPMUkQPd9eCFI5bVVN66C4DXjPoKqCbeYDM60uvUZ3iUPZAr17
NEzyclluu8HB08TD9duQTV+EQ5NMI6jn9B6Yf+ITEfLNNuoj8FZeLH3TtDgskBgheLCzC6GAp5Qq
0rjeXqLUdal/HLGV+mdMMIobUCh37to3l1jjCFJd6dmGDSlvonhcymcJaFC9vY6nqR9zFKB/jbQy
e8UqZp5TXzK6j7DxQz9hnrZ0dXGqk32Zkn78WAdqonxtkD5U5wstIf3iA39qmiDD/i448uPh1H6F
7LSmB23iEn9AeOyXGOzWFoAMeWY1kkdR9B3r8+aIfp/y2cvKJNd+q0vtMmWuM6zEGFitOqmNkkSW
UeTa1Mnbb3L+ot9kPiLQC2M8f/0uPivhkHE7lvQddxpAwIx9VEDHy3iEXBQEsFNKLYoZqNhmcCdK
XxeSCOv+RDzS0pr/+E20o5DYaMe4yn6ROAvYukMKNs+qtWmzJm3/QEDW/Stu74dur+oXd/5MUxim
eNjcBvM1WSyujBJYUXmf7ik12KTcNIck0dKK+Xbi7YG1G/QmnttYvPGxfnCpnv0pjDLbn2DrCCUS
6gri05egvlBfy7+3ze7+cxPYn1REhQWR6z2X0x5skl4Guz//0Mly8SC6k7AJNLHdME3efTOMvvxs
CHDSOEL4kCnjwTg3tq9mEDVYYWbLCy7rF6+Eem74Pskv4bnCCCci0V5VJw7l5Xyq/oiimomNS94j
akzLPa+M9q+o0Pf/Ic8QHabvoobeJTNAXOMoji4UzqrW74rjHXITIJn1gTNN7X6Z/M1bqk7IpJtM
hyZllqgGnxtgKsGLK73SX4wLDf+FHg3Ou+EQbQJJFLRYbAlEIEUjesTIbfGvugN39gd79ztak/qj
uTH4wVZTRtwJ6f/olpUpklfP3H47yN0LYQaAKvUfmrxseDRq/89btJKY8K+gsn8PrqlKwmZkPfDd
cPv0sPYW84asj/PAoLsK70lAD/LXlqZwzrIH2NC1z5/z52v7zvwp8lgemELfXbVsnfCrO67B8oX+
K2odrnyyMFaPbPqhdSCc/fozS3PCYbkrIGWpTbaSjUl1vpmEs91H+jJkCEqycSHBb5O0nUUAVlhI
2Anpk+rTUXAnaTz0VDUYH0aueFeZVQ+RBmuBt6+T+fs8pXDdYGivj8AMF5rdHec9ZsIMig9oqQaq
OuzQb88z9JOheS6Q8yiQ/6n2+BtkhIk8yEmlDFXc52uUoGXCdgal+D0NnFrtzZ6RbPw4vbu8Dr3E
0Zhho5P9vqAhbjQ/OCozCOAYSr7CdoxP0ALJCe74fsX4rHYLmolENWyXRWTffSpA5nySNT8RbJc+
3XfnTHNEHudWmk5oEvSWbx8IbO2rj89Lwc9clevjfgi+yKotccp4Pl2r1nXuVqfJT0UADvk5z9g8
3fUF5VUaIukIL87gi8fFzJ8msnuCReTCM1i1XpdJrnozpifqMOWR21RDdHAk+KR/eWjFvebCMNzk
CZTek0e6+8DxiQ9+FQ9wRMP7hZ7i6qmVx4T++JzwdZLmRmwzQbzG/teIK3nzc4Rn4Lz87AFJ+geX
nK6YTlbN9HpUvaaemu4cn0oHMDFdug1Uo6/adPtDaKMKFzf4FxljNc/tzqMUFiH8uIqt476BlqzZ
Z7MxSAfmmpWO0oNmAE54gkmAwuL2J6yFnV9FGzYJ6uXjO4RLIBRooT/KyG9E8d/9vM3YA6RHehya
JjdGh/mQwWABOiN9fMVeQozPwDHd99+Wk4MTUMxxG+dp0TUJcpmId4cSPXjZoI6aIv0+/uoRjiVx
5neYKUtY+N4cNQG3UvEwMdN4Eqw8yT34IYdzEe5t+O0u9ma1bJMpnzJqGbnosBa7XFtKRDMJv3x1
qQX+/G3YklSWIkC6clVVFVkUyZH4rAhP4JZf6vkdKso7ho10wpg06fzYEpnzWMamLFd/hiClY838
IG8UfaKObCpahkH4bnw0UAwNd2WEfED43khIZ7faEufrTuJJ2hlB5DRyLODpPLyLuTHV2x6HELMp
McXI6TDLB2zeXeRB44H7srlDIj0i/yV5NOwGvjA6kqzdtdd0QL9cBsOMidnfCYXVoeF7HgwjxBdY
juRYW8eQZf41HhsLcSnV2iJGPE5j5WhHlKo3YvDATe02hzJMq7lvwShZc/tDD9MqXkElJMJm40ll
SEDoElYmsAKQJ4zukh6FFEpU1GxeIul/euLqmAeLhIStUymcGq/kXlbpgkT4JhhuV3erP9pKNT9x
qmoV7hhsWHK3PRspWzS5iYheZkZ3mcjjD6/Wj6b2cXdTTha1UtqbbfSZksCLgpoBFOdAExcgOCPI
UZmv22UDoDn7lk2j41oPREHEPkn665uYJo1IOlRwVvKksRUX44WYNfxItlu69z3lGFbXymI89QkY
BXAVehSU3abywq6ZeO0F3IntykbmMxu3Aqpi7KNz0ap6tILUKtXQ/EWbYON5prDPZfMzv2fC//Kc
4dg8P7NgPZ+DU8wevoPV2O7GQx1zwiK1V2uYYCEtaKQqe4JYzaagEWD2lb0YX0rjUPyEx7miP7NO
7JAIdgQaNY9TEFuOn/T1mIpepOYlgbNgHAicHtq/4xU/n8DKTTyoCTkaXlwGPdag8e49l46lzHGs
asXZdm77vFSLKot71qaqDV6BTyE2JKFDu03w4DXpneR8qRoYjT3mQJUb/tQdMdI8usHBzqU0W4XD
bzDIuK2cYcEnea4iPcsi/REJj+a8qzeRHTd0IakE7w2UuAvlYS27XB2qk86ddeC4pULhAoPX6D+i
tIT8ShXpcVmw8UDZxcl3zXym/Zdz0Ur6ge4uR0Kj3m5sZFbf38SHttbzvhiLzMl58jKKmmyPGQ8e
mtdgQ2NitXLzum2Zp6QUkYPvzvLQt7IsmdGm3m5OPB7chbSmX5trbN0rmdYTJslf9WgMNXIDSkKx
DM8uRLaqbFb5Y68DQ+jS7jm1Cej/+x0B+9QDWF4eM+OrD6FDB/cAhwsp9bSbNG9FVfuhCHb7q+dV
K1KmGedjkZa6a7v36r/mmTqvdCMxVwRdIQdd+h2mrUr94EYXt8PutiKK0azmuNeWEjY5gGyrnFlR
iqUBy4jLa5zQnPguRlxVJrx7ogzWRkMPvSwRuUwakokNFjG7/LIk8Thnez5GoxOEA4mJIXC+E2k7
noT71imL0fAxyvoqgZtEIiLHkjJAYPG76Jkgo0EgZvt3ku3i4YNBvUTbP3dTxJc7B6VDhhvUX499
+/ZAJY0VozXkKPKHSlEKepnS1YnyzGlBAysgCJNddppmfZRR4GL/kNYOftbWCy1ahus8hfEda+3E
igjJ+R9dgTOyWnu3x1lUUkvigDC/D2GqGNJRAZ1bTwrVZsHfB+BoAzINYhVKyNP9z1+ZgvZcBfny
klC6OPo54pXBsWsimnTpfHbIWGMoeUGtx9suwbu6DflKVWZb/++Kw8E17VBzo+5/vRPVkYRPbxE2
ss0TXNRCpVSXFYZDzcINF2u4yYHXHg4M5tVjOqjhFTelW0jOFwDR3GSwFlXdCKaWKjqZCkwN9lf4
JBaigoh3Zgfiaj3JiMuvF17KxK68v/TrJw1KbSLycIgiNypVywDdD3DqTQYkeH9gedc65dXUtzd0
oSV9ALi7VxkIohU4PiBHZI6IsDjDwTLLnJPLL7Xj7PELaAhB3xXfrWQy0R10ZRWxlfMZ/jgPuMEM
eh09eYevxlk19tcCiAhfKyKTpnUojwVt12jV0XDzGG3J9TFuPfX4X7TZx4+5aoGKZBaHy2fWP+vP
8bGGeFB1/R4Y/lW1htl5RYjnCMcTW69Gbky435Q022BJj4394xB61ZxsEJ7dY2g8t9gyLaJUg/n5
DIOelCisk8ELUs1AOzT0RiT/HqE9jw2k1vYqTQiFk23VvbH1DVjD+NpDqNJIQ1ASiKJ0PhfnjAUi
s6WnJwwWFpB+oYS+G+vsaM3QvWxEHO+r/caAyFh9AvHGuyuuKwX+KDe+aZCNPt4zVOnmJC5SpXDH
uOKB4VPhVphHEjKKJYJZBxqsUENMEkeJfI30lfDfDlhyhcaFmr8g+2aykAtVyQpswN4TB4kF645c
tux9KEsbCyXloXy/vjpinEQuWef1Bh2C7wT5TzyU8F+Eu6vdPGVdR7G9e2UvIdvqBuqEPuKYGuuW
xXYTzN3dXf0YrcvOV51wtGLsr3lHvARm0Ci8Azv9IiVUfYlWdqtnkCo6twqiRWyITRcY9MICUNI2
vYfH/yxyjaiPDhixZdsxg1wcHZwbyJHgOx4Xjd9HQHDaY8jGy0qAl3AO8inr2mnhYJC/dmw4Y09z
0AcOO69BxMNOX7SLtTsHLR6Fw1z8tgySFYdu6UYjU63Fb9eh740UPWi4Zw654K4LKp8yWgtZkcXP
4HiweKPApsc3dASg8fS4sIDTHGZyk+ov5oqMUHhO3yLseQLn+RzMU40++E6K+UyYPWlj5dlMO1PN
CVczdU5hTUiSb3CllM9lVroYSigpvm67qDwkgGcM+ZSq+Wgll47sdJEmE8UGyATZQVujTAF+5kYU
PzDx9kWdw3OA1E6ggNYtldWzU0fCtF4GxZbD5ErOEHUO8DPtmAZJbFC40B7SzBZYLWQ5B2jLYbtS
/u5WmeB4y8cOvzxHuYDEzPgUvyOQjOqbJTsqf3wKHPnNLLZUqu47guHAfNMyZEzJIucsmlwKQ8Yx
sL7A050jGSWp8EXtTPwaTmk6GAWfvSl3JRsGv0TQa4T1X/xDmWWgze3KHoJvPSGIr8QBbQVL37GE
xo907B3TwOrXoQibRK2ID6ij04j22AwkhKFuxs+x3PCOCt3Ec9KMoRX9Yf4fiHPieb7BZV27o+Hd
dlCWdqUkVKw7K11RB28eaMjGUhLIQgCU+cVWaHf6IMAFCsvUrHOpyJ2AyBwfsP+kBkD5+o5fhWM5
JsR+kI/pMei+4/2gRu/dml0ThFP8Tyvtx4R5YqhFVIkDFgctWDShSCecZJzLH/q8EHPHR6Piktpq
uBN1aDCQopUZtsQ9Ta/bowNfqpI37hjuhCC646v4EUWgqvAXkHh46+i8tINslGKZet3QHQ2enkLK
Jr5kLP1Uugitiw9USJEwVAVHY8RJUDFg3pTVITO4NgNfm+KThBmBFpkqTpzm8+l1mI62X3MNgptw
U21tjA/kOM3Qkcm12ShXOkZzA/7PBpquh6sLdL7N+Wvel7evcIn0aohWfaGQRuqNrV/xuhkRH46X
iYz6vkWZZlEs8Moetwj1vqkZ8jDpAcXCzrYIQsquKW3ZfuIacSSYbq8YX1v5Pq6I6H8GKdPb485C
PLiGPiDYyMVGWugmgXX6BLWYZViljzeRoPMqlV1F0rD0jAkxlf4vLfU0aaL/IZoItYu6G0Dqa7Ij
6uBMRlOR+QXai/7tjnI2EXstqbapFHmfdebb4Xe+urjptiBN4OZKlYG+TemMoLj1licHCR/onM7v
MXvBAUhb100q5OH4CHYyLlF0d9OSvGATt/YwBRESPCjUpGCJ8qK29ZSeJ3b6+P8si5D4n/qeX1No
UwD1Pk8XPrrE/eR7uOWbNGw5mllGRbVX0/nRovBb+D5E8iXbEInw2kVpcxvUXvIdg/iLYsdmNYTr
Vu04A5NBYNKaB0O6ZNRYrkeT/DRICXmFlsM5UIZDQEg05GtS2wga9sIa7zgcEb60oekfxwv1Q2JX
79fDxvbRK016yVXDZ2k0GmCxLLodcZoqIhH91W8TDEpxXoJLYUh3BgIR16T98J1yww7LSlzZmYsP
dbQS9EoQpC7AAHatQLQW8zQQyB6aFXLQKJfywMqd91e69u1FHflVccLoncyEGleVeW6Xatx+5BAT
k0hSGflPUQyg6ZdkOVCv4zDk9K3TKAXPpAXvTquU8+i9Fzkqtt7w5hMQd1M+XAf6zwV1ZsrETHmy
Kog16y+q5jRKbU8UZA8Z21AKOv83O6KIZxBYZioXZ/fB5hjINklCBU0lncDGvR9Y0B7LgCy/4ePZ
3U/muH46SeDYWtC+vvA2jaexrHZkaMB3OKCbBxbAhqcxLnAjJskTwlrNafpdHrr3ZLHbw8sMzIm9
Pc7dKkrcQJ8InZlWUBh2QS1lR84FSpcRTnUsXeGEuCdQQEtsh/fj/7kY0TWGIsaANdJ3QfckYTPB
DOrAtAuuFPeP7K3DNCgtrprZjgzLpTRWD8NX6z2ilZvpXkqlHqygKY+sTgzH1CvLSiPpiNM9BpfJ
vdJDoPUYj+LUtGQAqL/4BxWAf8ilGokJ1dKiBeOeG9eC1UaaRQvF/2sg/lEqETkh4WKxRq5+PtQr
vnIV+0cljP0UVY4KSfiSBlIhj5ZacD9twMmUf4zMDBjGNhdUJB8w5sBYNy2N4YPPVT57XdL9PT0H
OIjl2Y4WMa/VlOkAmwWi0o/dEXpQrl5QlzZKK9oyM75iPDurhiqugC/V94sU7B47D7WxdbbkRenQ
VHBmJvOtENXlIGcwcCubgsxBXkwRMq4xIO5wzNg5a2cRKttFNCO/eUsEw8esFzuDYCVyLSUeENed
uNyeaegkkYovJu0Da68BSOMTFEc1FF0vgZVo2bbnDQ0UnijPl/1vEWuYSv8k06OuSs1Tdi56m/Kw
HI0RT1uDlAHnv/1msnkISJV6qH1gTL3nMqolPf4Pm81CbNCU9syYYRWECYc+AV0RCnC0tP43NpWu
Ce5V4p2BjDlnEDgA+O0G2xG9dOvoes/S4giyBiGQ6MPjiT/elamc5rqDAU6OzdKtPaygh+cwdNGE
OBmEmrQIJ6qXvl/iQdJVX7gdM1a+Mr3rhlUrue6R2GHNAdgLTtwrmPpQC2nCoQ0ocNWh+/hecJHT
lntmxX+QEy4U+4IIu20KD3eYh1Z2tFBHOtd8lVxpsuvfUTz0SaOhqweUoYLLWQIRdp00AqK5seAC
WEhwTdAS81dyGzKl34Utyuk0iWIqe5x2MPrkdVdVKA7vfV1Eq8mGqpdp89NQVSv3nrUUtvoYUYFJ
qkfQz1ewzI5RCHxEqx6ddBn3DyztguMtwHw/xBkMOT38PwKM46josaVDQoREXNO4sg0gk1/WDYXP
vnq209OcKdJpD7sUaivGUloN4zKEJL+RE/TlcIQUvfx5mWdsXqshr2f6gErDdLZCokVjuthVixeP
9LhS5oIKbijhE6WLjs8ERoaWfW7qHpIzbY2J9N468032i/gQf6CR6CjIrTCwfxqptzKH4crrcWdO
3EzZEYL7Q3c0rORfIy/SJbLM3VArJLq6k1AUuKmHrdbrH0bw9GuMHHJNg7cV9quNG0QET7S8sl4r
LfWA2ughfsnw1VtnmL0ysoeb/D0KGKu5Ti4AxVMlFBSnAkfXpSwwrRTcZdqRCbz65c/YUvC9+3/N
O0qo2Hf6bZ6DY6J8/bMC5bAx5JqDUMpy8l0bJj2yNBd+83ACIxZgt6eAsub3XlHc+RaLJ33AE5mh
RWUa2QRa1FMAiCP2ccTXFjSLZiuNGb6qbgRm+ZUcaX4jO+5RiQGx2nBFKJsytBEUfAuYk1/oC6JO
jQG84XYKCaDzHKVXjUWXVda8EL8zba7gwWInH48WpFWClFdJZ8Fkk00HspFZcz9Qp1ItudB0rLYf
jJeTy7wlCH+5CtVSdFzQBxlonnpCq0ee8Gx9D/KugS8AL7bzpAqx5wulG8yt7pahpEn6HBSJ85nz
uMwfeOTfmlYmjctMyPeK+UgNJ8dvwJlOR8l8Se+deML0EC7ywr2oHGC7v4O8XQoVt7A8iHTr0DtZ
wf1zhnTj7GAJlOH3YiLGOGs+OWmiLx3qv5jENoXGLHRBRfJ08i8ncHavqD8lEKGoIsQSXqsFiIBo
Oct5AxYvj6KhjKm81ahsG+UjmYh1Fpxq9k5wat2j1Jjgilxv5+eR6ghX7hZmWk8XdV1qI/3TnAGJ
V19XucNHTdUcDaFg8XFGeWQsy/lFcjiqK8K0kdShwCOJHI/NP5QtVJsVg/sldK9BD7+2wUZGaWcX
hrAHxGFnaD9Bm9M6a1MKqpnZHonUT9A6lHtt0RXejF9hS13185yEE6OalWY5028kezmr4jGB8R9O
w/ESZfpnUfXhT+3VlzTF8+gRqMrWwN0sMtzzOwuuUhZybj4+8rWB7SkBiESQg1wqY9SQWnToDZUa
dz0IoeTEG4UX2+7uS5vh2je2qCJ2o4gY+Cp0CrL36RBLy9WzYW7qAcPGVPAbvr+Fqjma5onWaaAx
Wj+1K1r3WEIcBLLtNkY+VFnZWW6rzYqfLRm8E0a+1fL7WZ+8G7VJBq9tllyiXbJSys9wJZtRDSFx
H4ZNLp6loLLXneCkAWm6mbAB2wYvvvgOuotR97UfGoviBN4hiF9RQhmH+OprCKZly32pKZM/n3Ae
aIxdYVSD0jITplUADLG3dw3XvkfyQED+S+Xgw9RISarEFxmGEb/saXS+QHuU5G3dOAfZVZu2DdDS
osy6R4CwRgkjY7Odrhdg0h7kLfIr+704D7etgdBNWZ5Co3WRYr0JtTo/DtvNnZD5zJrLvctyW2/0
tXzNDdBQo5CUffwzv4Z2W0K2rGz13ljDYodeJOmLpiYrXNr9BCRE6TkhHcmdfKUwpHfbYdseK66R
EJlRLwjTjyP4MhV01EYCr2LpmvPbMOv4COjYKlnRrJA5GbHtVj9xNkAQL0lKtl1qrXxhfSGvmgR9
Uz5LC/CiRRkiwhMwi40/d0DkqvGHptZPb6V21Zvjki2OyPOAkyvD2H7U0NiSQOM+5/eDdHq8dlyW
mHvxYVkl9JuomICP0C/e513liuyFc1d9PqgBjVocrtMel1I/Vcyh1jZ7mF8gJiQ5yP3geRWRqrgi
M8F1onPLAjWORHOgecO2k+uoJl69dVyKCD4WssuqYobmvA4CaFOd/MvWUZsvn22PZ9WI4t4DVjNF
pis/wb/qsHny6JPGx6LoHq6AYaWQdB0Dv0GkudqOMMCrQ5UXaIAC3vDghnIkUoWbmelQoXNMAhTG
ck8cvxr24IqaPLDjCfDLYhWNuNg+mstXx3+EvG28QHvTnDefQhgpZQ+pzBwwqLvGSwuwxTTCIhpZ
1a++Nh4ncyjuCQi9MRVyR61xYCe2v0FCg2DR7KGGnn7mPVxrQT0rEEycSRjweEaKU7jKwkuB6KQ8
fX99GgVPTvVfvZFwhakZtpfuATKvlIuMi0aB1meOd6qfP/0AcF6URkM/nNw9P7nIPewuUVS7PxM7
woYs+GU5lGV4duXgLCr/FM6LY7Q9235AkC6Sxdhqg7RdYJ1u4LeSGNu19wLndZzkx8t2VndMbe4J
O7VbA+pFTlBtCKc4edXIJa+Bm1nA++KMOeUSNywpzRiJ5rXjuNhivNmUD6FX5oSGap6gHTL/SaYm
GJnELX1ZSPTMH3yfnEqEVx7xpEpG5261QyTBQxjvTiutGEPQOgfDIVkIqx7JIouLTQm5/xQio2e9
LYzKilgWsOsjaUkigSKSxHIAs6Jn/6CDaQW3qEtdVL+5Dfd/5TnHDjflaJtPZf/HYJzrqCg03XKe
du4gi/ZQH0rKwyshJ3wtTxJNkXNko4fRgbgpHyF+c+wny2L8kpIihRk7S1P3PmKtTJe63QRQ6oJu
ijpMuTM1o9+P5wuKrka35VOB1U8OnkcjfKIOO362GGL5cNppzssLZBxAXnoS4agVhhIwzxZuVRHh
CsChfjj186EO9qLsrXgNmDsg/tCPBp9L9qrZYZ3xNyzCPcJJqYZrZTpQYqjh5T63xIF/9EUvGqof
We7XTYHX/WDIkzdRsMmCX821hfL2/i1Mbf2yoBAvM8AxqH++mb4l53JE+XeKFVXVOs23knkRET3K
N+PtAh+qezzkM6IYK3kgLNVtdjTaze6hcf7FAO5TnR7KQphOogvKVDbaYW2ZecYXNKh3w4+TOw3g
okO2iAxDxmDnEVkPqgSlwnK39+Ne89CUxJ///yjPkdVtJIueu/Y2g30BLoVFW1fj0WUgmnUNOGLl
svbk7h3vassrZ3cQGj7su4dPisdy7MEi4zO++rs9cARLGLWo54J9IHaL5XpVTAcEw/MKBbUtjkoD
0pGMyoh6JKprEEpH5VK+qEG7PGYJg/pGV9n7cyS+Fd+3F/KyDBoODfgwz+8zWbRatr9BfUQX0W/E
q7TN/efcLg8ruI5AcTPZzhPYZFAzvTzgNJQmBgculz4HfcKXYRui/pW4ZEnnbiz2cbnMfNM4OUzA
7D+vnbGw3NkFRHRkcOPqH9kSdhyZqFi3PmKDuuLLIApIx303ylWRunGopXlDHsJHvdP9AsJfN9tI
lmU57mN7SfNCkepKwvasqGz6EN1wEELJvERcr0WosovWh3/O4oBdnhbw8Z8jH7Ko4NOdf/lOnlpM
0xPjzlWnpeuYnlYL9II8XAuykeg6HvelwzlxuO4wlx7ayQef92isl7DwNfq8Okbo1Xo6m5Sxtpkp
GUhstaD8SkoBrLw75CRxJwRDxGvGnn4Ad5iWazA5RGmb2zYYzS6vCw2icE3cl3MurwpqrtNoW5in
Qk7fHLPOewUp46p8oCocZYvU+YbwvI7+ZRg3zP/XoWosvsbs5UJPTSCae5IjNJUkvWcDq7Fb9akA
T+Ho0crG1go7zwTzP2/jsxL1Eu0+NRmpWh1DBPav1bn5SL4E+zQCKn05fFRln/n5S6XmQ3IlTQC9
CCcneYGYX5qv84cDMnt/6RRkvj3hzTX4goGXbjc0/dIYUreaaRKpdUZB39bg5hMvzfwiCRq1AsX+
NC1ZwJCDTRdK/bDmSg0VjN+D9kBxBhz4KyqEnQ+0qZmTRzv0r3gazAdmPWnIovHciH7ibgRxxWxF
/dNqtxzV/jSu6aT8XQk4nlL+9dDCueof/H1Q3qZy7Ntprt8p0cQuf6SsOYOKGrWhgRFiWka5RQAc
uG0vUtMsOVlhr2FrEbuEoojIcRlzVHWfgdUbfOnnwOpZVZ1SE6k29GZToR4cDbffp9AI4P/XvCYN
vAT/w/Bf+06Vy8XynwTLWb1rDYR+CKnStu/SgBmt9ckcRwkJEyv83jIsa/ye6h3DJxOsj6PRTCD8
l/8UPuMb09SDWI4cpt5yA/mig/900+neac8/YLI+cbZM1I71C+CF/kKU64HWr8Xgw0IVw4X8Ufja
RUwk+pizOm8nUELOscJ7L5vhrW1a1zzJOUPXpuC5Uiyta+W0ERUIfsv5CCu9zsnjO8I38jKy6ccD
E3G/lUeY/dk/BDhJF4lkuwYUyNAJ5wOQpcGkx1svfVKihzQkwk11k6HINlO5NcvolVJdWWVBTWG7
aRCB24mwrnRx4dQkYvHtcHm7+oI8Cr6btbpKsCyzJ17fKg6N2ByudwK1IJht/bq395fmuG626q8G
8wInC5sg51hiPTrMMWpKTJj1NuSPkndABrw6lMttsmG2k/1JOG7YGeLBBAuz3lcVgzETR/QT/MBB
To9S7sa4QacDKZF4iEmCcTXCjjZSu/2/422Qe0D4/e8BVmB1nCrnPElK3TLj5DsPddN6OU8fVBGH
n26E4IEvKvb3CDd9siHboNZPHbyJS729m3jsIUkya5njmG4hYTx2+2J3YDfBuhXAJ+OnEgVY69GZ
LT/jJlZG4PO5DN6k6WHZwHZtJml8YTRVbAwBGFQFK2WsfDcVBuIgYqUwVozItRHBNm1rHpGNJib+
7c5v4/f3uuzjgaKayrsyhwWOs4+cCpMwnhOuC/CJ0liF/m3hyXA29JULfcIueoJdOo7NK2wW2vUS
V8fXZ4DN4N/ZEelmTvNav3Itbo6Iq3nYfo8YlReeaX/ByRlf2zl0WypYNAygcRuHCc0fWYR9hR1k
K70BlzitrTFbSdYZLTwzmqXNYiCEQhkN4YgIPengY3WTP8akc4Ya3t8AY9EpJtHWvWafpVURId58
3RPKyddp4IUemwBSPWq6l6ww0oEk0oJnN1+VW28E5D3oCcrXOMXYd4qyOni68518wa/zpx0DD6B5
mG3WTpiB+pOSA8pCmTO6EAaXB7Zk1hix5yIOVtzjoFppIz/BheYhvpUKJi+AG2luBiImw9TKbLRO
wfPpvTUGpVmdDYc8kfjQTRQ96T43ua/wwugd4f1Ti+73yFy0snhzYdm6Xpw5tt6QDkqITb69o1zo
PmXcB+NIrp65I7PeNvYkYXKrGlR47sMcBzDqDx56zti+cWwReGY+wpdK7o6oz1TQPCiLlJeFjZac
K2urDCPMTBq38bQM5npn47GfFXCP2WZjxpUDPY3g2EDD9Q1UMVRhijJRHhEEZvByAEPsbe/iB+7F
sMY5eBvjNgEq6gwjsOtwJksHCjTNqbRfm/CaKoHPpUX1+dzpSiKW50L5xVicDEE7hz2pqaAzUk2c
tmxdJbQeLV1t4pUht4r4js/FblgcUvQFDrEA5sakZj9w/ftvD+M4G4v20ow9Uat7eArCbayQJGQJ
FUwdoSBJ8cc9POZOxT3FFW4tBzKthda3io5v8XBxqdUTJ812lLVbGJfh8/nulFH5h1lg35RBE4hc
wlL3KN4UDvLeruOUcTPXMgYBlfWSMngUJ9OGDOiGzfezz0QwTHPEjcgqzWQvCe/jzkhBAGPluFiI
BFfejHPZEVPNW0PV/Bwp9Vgl8AlFtEg/qVdtiD4Xm3r8215IRz6cRMjuMnSvcKRFkEL5weCehu6h
Jmd/2AgWxhqiJYPpEE81imQoYMaWw5SaQekiy2JrdClwGCuhq+2erX+g4vNifgoO33JVVWEKiki4
y89cqPlM4ExEzuuxIRa2LyCZdrR/ih8lm+MW9Vp7kO4gKBhsCNmKiqX9LIcnFHl/OSDnyHsLXsiU
kH4lPirJsldm24uWfovRHPv6ER48CzBZwcKY72nr6uHJUiMSsjzNRBFPmwblak5TUZ8/y6Sqpc4o
A+opKDqB1apQePbPT9nAdBlrb8NwpR69oUHMPn7ONUbAEhAcDoFy+FuOI8IeTcHxOHTdyUtv6s28
K5Ekm0e/pZuzZlK4CARbzFLry5Kaj6dEqSkLAF1X5W9k3pG+QP06D5ubPpVdtBU/Vrrsc23ZpEBj
KUdYbbeIQTrhvMdQui6e5KxbiYP4ebrC1zvRjw6sAuAXUdn9bMbpNV0OHmb1vyYUpjDtAius7bD+
z5RNEEfsVP3NGp93DzVmGxvxTlSXUwkR4cRdfyUgVP12W74k4C35844P7kR1nSWwsKB8mu2cIiph
qljdhmF7uagfX6UEFq5eOY6Xi2UcjjenP824Tfj4896AIpUu+HNfD9JnPsVep1Lg4XzBMQPUR4MQ
u+v+ufUY/ycGaYWgpY5PDRN3Ja6b/zWlHue8zOhmr+mPFuw0KsntK1V/vrY0XlHbJaXWnAaLhUfv
KtYBM6EzvzqeQKaWcL8Rn/cf2HSgNLGThvIIDGoj8Z4HdqdroGQQhZQ8TG18zw54EvUvyapawHEf
gR2FXIdWY1G0Q7hLVUFQ3K3J7Ai0OyO949jR9CcEoZ4mh2i2U1uoLTxH9sttQ6o5Mvth1YesxNnW
uxWSzN1G7Z8vL9sntuhILjWXvVF7PxE5i6e1iCljH3lywWryk7m/qIqHnH6ISfUoAxOQirlHLpM2
lqwO3008IW9sjW5r0HqmbvNC5TRUXv3wB4+qu0iBNbprEQjlz+I1z/mKYrzLpBEiYZRVanGyyGVi
Oq4PNUjVNvlEgqQaozTFYeJaxUYo1kezmeBSTB78OUyJ69nIHw+9ejZlIKAWSifPbgTjluRu8Qax
wmgQcIJmAZ3KAm4qkvRr6wLWUiaQ8UQLv/0uh5iGS0AWGNfoaU+iVW+pz4h2E39LX35sRISViFKx
0f3dA4ygiZpaFnQ8rNbKaG2ZHGuk6ID+2tqwAQuriiaYlgseNYhy0N9DPckh9L81V+z6CN1t0Z9w
Q2zrK2TBmYuwX7naVXXJULw+ZlS369h1bNUXnAKTgPUN1YHs4R9/1D51U2vylblGlegekt4dDn/L
kYEttAz1GvTPTYpyr+bI2MXYZXs77kQhcXPrrELk866tMuwK1gjrcy/0BpJ40LYC5vhOtBt/zDRQ
BUFOzC29qxgRqBYef+22qzRzajHM67BwzfTvFQMq7UAxWueHculTavFjN9zwB/ijcTjQN4+npkbA
fTPVY2eLDFyTPDvs5iFA8a3BtTRMgu7GuqnmTQQCkIgL936zmt76Vicx9AYrYeWCni+4YGRZeUPT
15FpJzvjhz+Yf1ciZizwcjJTmS21KqFE1ci17UYCCkpfxZrhcVw6zeDmNDSmNiKOyM6hj5S32CC5
h2CP8+W+ysEn8+lQTiOtjm1E07PxQM1xC8/U7raPhf2wOhhvNqj3ISYWSN5ehPp0+Tiw3VCWevEi
Gm7oeB5LGKJyVyy3ReH8eMBd45H+sgQHN2C+E/K7hbGWsc4R43M6aMlT3viYi3scdkxVQqfwO2rm
Qecj1XWTNysXL1VXKM8wDbSAYlXRGloVicwEz01LKPP/s3i8zd3u/vGCVZRqRuGOdO6dwu272Bqa
qtCIxPlFO++AMKdKq7tukjdRfo2aXsVjnhLxLElYVFEFC47A+0EvsyMk9XtMAvawwncaU7ce3Aii
T4KkwVQhjtUuKf6l3OM59zMB6/jVZktxm2MqtfXUWa7pg7X3cAsMqQRXf6lyUpMo2XiYnqNLdtpO
Hpsthv+r/c0Zcbb/TNyq0IFFSOjS4xmGLkrvD1szVmNmcIyA+9mBjDxELxdEt1lChEP2O0b0CZR0
BmkwMmG0qve/rwGWdCzBMVuQiZGXjGb3aX1J4ypbUSvBIcVwCbAFYVuhFTELJfagvoqPfoccDTCH
UB5tTqD2zQXHBoMy+B7ImI7GudoyBBcVwIRg7drIKmgCC+CvPt9Pii7OjxPTKt1axPtXCXpLvA6H
Cxawk2aYIeescPVgdx04wNIXum5NLlefsU9aHPIjKsWVpsQSEu28Uo7gArCu5jmmThmcUDTypaSx
UrUjTj5SWiQEcT1+WcIKISSb4y0pePhGobxLg8RuVWEptM/yewxZui2X2XffqsYzVUpG0if+ZpyX
AqaGJMwJbCquCrY4K959HdibjEIKS+v3Kz+yz1mPUaXcvtjQtoE3jb7Uks5XC+srZ2ZAMHUfq4IT
jzd7RLoSxBU7uFZzkJ45p5jsX4ZtfYTtgnuJcGblnjEFmMHi72lt+0QYfGgR/RLYa8Ev/S/sRR18
QphGk7QBnLHjt0y8OjHG5YQh7NqJ4y2LRhUZ6on60A+AY3s+5sx887wVzkU3Ku5ZD2EUyCvdynHb
o/YF1Bqz67IPKCiS2kT/YWv497wNDynz96OI7hknAMlOqsD3sVbrqOz3lNPCOR+hBp0D9u58wkz3
1Awo479Tr7K2uMu3W1lks3sctVzfzkuK0NfY8ORKQw40GHVPNlGyR/mQYQYhSwVQqAd2m3NP7igJ
3kDSR/LdEwjIAfinI0ZE3N/qibcJwq7FthJNzaRDAP6CIkJaIhZFTO6ru2IkoAfrU2e+Y7QhRiTv
9mRHCBbMzJGZMyZ+W/ICbL78Lss/wJu+ZM8gW4KOUUvyv08ssooU3d1t3VfcXbp4d9NZfT/xqlYG
qHGrC0IgiUuivO+Oskxro5fKUW6fBARzD55OvUbhQjoDh3faok0DIWqcWFWtbT+3gLXgCgf5lFQm
MAyQDlYpREdhamUqg02c9Vf02XZdg2wLZ1gB+iKZ42uTPVEZ9QZudzcFfrA+jg4Xt7G3D1BOVkTH
dE7W8uo20oYrE9Rv9bTPlMutOBfeCAVW60yPteS7bf+DmKF+o/DiNwzYzXcXUlkrdwnJzZ7+R42p
kDaZt9QuIkg4v4QX5eUJ0gYFt+SLz++ohuyaD/Bjq5QFafurZYPJVx08i8xcw5JsCHwzUt8f6viO
smFq+cwv//RPjWaKvJkKsaHEMz93N9VKhpVier3yW8D8Q5gWcr5Di7Sf8pGlup2NbxUtpo+fCySZ
/mKEoSMZYoa7Ckzj7opgyVqzX/mcbEPE7CmFsUzfhiBWLJ9fNoBahFBZnN5NnkFe34KX/B79ouD9
HXRIsUHW/XKmUt6obHpI6DZ01sgSrEAuIogTkM3t3vdPYVG7krv+UOwDyLulw7wqy0+DcMdwmRlB
NZSO2Pu4JYynHUQswFrGGwrkksRh1IOuuXo57vbXoj8JlIxjVtRcKYH1//kyfL1C1ZpyEtgIPzS9
xyNcxS1LNtgCLtqx/1lTDP+SNpE58Xxw8Db07rUEFiWR/o0HkumPtJzAEQfhLGy+DdIsUBB9Rlxp
Tcec0FZbcEEvNlADQvsgLK63I9IC08hT+dGJCkPm1Apr+oS6QgQl8aokvD7ptIIkS2k2NxwYtgze
BABBmhfp76zVKul9SxWpJZsIWbrhNMFNmCQ9TjXyf1iVUiJtEt+iSPMUQ3WYOYEvysHaH7kCZczc
82bWPCqUyZEEE04OUrEoWTcYJj5msVHt7YsJBpj3a48fdlPVRYVVscEA7okEoQKoMIfzkCYhmMLO
B2Zrqkr95sUY0ODiZCXuxOIvRIJuE8l9o1lfW/wweg67KbmrKUXlkA8d/05zcCe1jjkwUMhheFyC
3rURmIvzu+jzop5izbzKrMbHhyuY5FwqKabavBqVlYXd9JYoBZ8/RWHcfctg/Glx0EVLaojK7WeY
ngL079Qn12HQBMiaCrLgbi865hahi3cosrfBbbTG6DIyULnlM4jh/i8RlSLkfw93MkTVDx9hz5gy
vrXAbwXE1UNfqG5E6pctVYWBq9aCMvM/16ZmoAEGoNZxFGyf3ta65oH5+maL7o+h+HBQbR4z7V2K
+EaCxpsMPW4LaL4UDz3EvDa///pI8xh647jcDvsHXa/K/dyOMCjIrPl1cwfmBJHBXjjQWjlaYfrZ
DahvAtg8ECuEgM3afFYIfneFU8H8I9ynkEi+l8lTZXPIAtgFpOV/Gmd1oFtrhwxAtN70Cn4H4eBf
4I4nWXo2e2BplmBias6FQ8X462aikOwJZJ55KlC945tc6ltht/q51OwRJzbyOmQXjFEd3xhGQ2VH
s7phoF4prIVVa5ATa8J3Omw5myvfX8hRuXY6rYNkQjS5uH/aWGjX9qwjzZbObmrJdkjyk/OcvuuQ
UeewpdUGecbcfQU+L5541zh9lnIOmHdIsFqnZlWGQjnMZgxAlNJyRkatCbV8BHlqJEthiBObstvK
k82TDgR14SqLFqVvwiXXqqcT3LLeqnd2e9C3Y8+n53YW4118MOokupKDLKPLS3a52auiobQADOxI
26c1YOAocW7zFTkxEBmw/Qvn61yaQ11U0naU7rEekBPYan9ZBMs7DipGM3cDU0Fyy0XZoc4uPFU4
zxRvw41LHMR9oPpYhYy5NU9NcNFlVN+t6hellaAleU4davT+kFOYGDHmDc357BmeKY11Zt0k77zX
9i/33FZGoyQFmBknftiuquq4W5NNWL3CdDgqvbTXVsqcp0GQmQxmXgBiPoqvdYymb9+ce64H25bU
ji5/1nynmmLnru5g3a4FFFzeSZJn2roYqd/RLstY60EGVA+cBItJZjWDXXTnTMmBOdh1akNXaXke
rKJLbZ2z6Z6cmFZ4Rx827Q+jQMxGIKKAD/9eO10iWCIz/FfFj6oPvt99/IiGrP7HwcyUV26+WFiB
MTHn333h0YDiTjlqP7v8Ql15wfGAJXuIBT+n9YR4jIwPkcMiaHpCPgGq4wvxbIuJhsvFLSGCzVIf
8iHw6yEqAELGa07QnwUufeh6lfvopVHJ+Z6TBp2Jg6XU919UyorCshwSOOk6pBSmtdfZyA2IXrcb
J9lXyPG8rXSyvFjakt/gGUyRklx74FzlCvTHYs7hCgjSX41xgJQaA1LP763Ra3lFr0I63mc7WFEs
HT/Q6RKPCnR68BJa3NGxx+o93nLp3oLyDBYZd0TZeZiLg6plPMEo1YP9GgGS6ok20inzDwkkPK0S
s1aE0vPrPlckAryoY8Q/RbQ8ypAa2F1aw0QGVye6T8Cd7TupsYLO0eI/oIZdg7rI8HKuTMru04Ww
RzvFIQzfY7MpyIssm859vzA0C/R9T1kCpF9lCtaHmgIvAAlQZq1djRNFOyCHOn5TtTdzXb3jW/jj
yltNyNES9K/f8/AJgt+ZIpc/WWOwmXK+xd1h4lvvzBF1Ifsh6H8/ydHDQH9bSEf0Yijbydxf/Olv
Z1JMszQ6rQU9E4CwmBK4SboBD+mkp56tMoNDmwNNNC4mH5szg346Dw7+2xUBNipVk/FOqqNRrZTg
6hy/IiV8tqr8Fb2dUZol3+NVLtMjSkN5tjX/dqNlxz9LdSmSMae7QspuULSKZCZDjUr6WiIqAqYa
RgNGnphQVpilLG/kc9VryTMhUVIBrjLMM+2UiFpCyqHiR4R9m5TGg0pTNExHc/wTULPxKXSf3Sst
x8Z5OVDO5MiSO4Scbwh5U4VKk5R/BLjLilphA8YThqULwq8yRgWbKoIA8gSNxj07/14IjpBW9AaO
xcBc93RVxQ1Z2HAVY8rLamD191gFLLQX9MvIbs9hFPnvLqX+pJcG3od/0oONUvAJsZu12+pLgBIl
GeITxrZicVtLh8lfnvejoBQ+BaSyROKRl26AQ7yCNNel89iUsY2tqLX3ZRJxh8LUtoNkgh++BsyE
5IDqJ0Khpn71ZWLR3gnkDbU+aW3bb03HrID/hMyK8j9CTfKP95cdPfc5VSL9glN0fAvO6PI3ajyx
mVFebNhwocuozfZSqQYiDqHF2wF+WFwluGxXvZA9D+9fdjskpMc6nN7moMNF5QR4dgY3zs3KN9u5
vF93hTRh8osR0YVFgVmjeHzAAy8tmuBycl4xbouLckZwdMU3d7YUP7jplrPkfrDK4F0E0FQGaXVH
PCUrYKQzXSxm2o51Z69IW7IxA30a+cODT2FEuqpuaD3QeiB3RNqd4ReHza4hJODb6Rfzy/iR46iY
OF43qxRrp17n2o/xOXfu1pPuX9eZJTDjaYz3q0t5LIJAPQgnyi9HgqtYbf2Khcei5JTBnUfKNMWc
QXO6L01IYGZXq96KTwr08Mv2h6fcgCNG1bTzAScNm8/A9XHXP+JE/g1jt4lBTLgcaT0QWOeiSA14
ewcVnnDL1ooqWraLHkMgZsce6p2Gmthwqs8E1K31HhUYHhKp7oOo9yo2Y/wgt8D+j1DKa0PIfWDd
mlrMihCnz/B4sc0jzznvu8GRBsl5aA5jj/NQRzGNptalZD8YwLJ0V/XRaP8s/Oupsvs9D07KlQJm
eJhNr4Kl5hkPWSGJb5Z9/sY17n9pXWHvoirTV2/Q02dBIhTx63EFw2zj7mTh3/8BlY3LMPTvRwwf
z9NfdjrMYXdYTm7p0d+9++Vi5s+p2qTm13Q7t6Ah+R5mr5wnTi2v8DjdllvyCEJ3X5Q1gm3xDm87
TFU5SbMLfuo08y0CnKTF/HUPXRXLDqHIOGckyalvQzloiX7CWQn55zRSQzaeyNsKqtu7cheqGYTg
r682F2SLXYVRNm2c3rX61Q+e9U4+OIpxOEL5+4jbVHfUL/0ZgM6bGMdB8wf2hlhebDHhQxilLd1W
9zHKgIB20hBCVztw3detfiuC2nsoakmOzzyPUJ1AwF2sTb9EZRpK5KgFrrWOt2z5sB+VikgaNQae
XqHDf8c26QZIQgNAbG+bZI1qBMiAdAMhoIlfIEZu9rwNOn50CZld5X1DNkk3SLl8KuOaW4dyAJyU
w6dlsbMfF27voyJkUsftQnbr94e2USOZcVDwo82lYQ571Q8/DdY86qHuJVIESiWPdjkDjSF8CjMV
HD/13tKlZYJbVKSBxuGOe4r0MSDsxhDHstVtFf+UOJvtyDlC+QZesxMviqit2fX+dixog/gIR++D
L1BEOH/lKEARkQz7PLZUOkIjzeuWtjpde8kqaUH9XpulTJast19N5ZDYSKTmuGPD7yoOC7WzY80P
5OOUCM65OYgbs6+sByPH/huGWsa+Fb4s/RxFp/glTqR/I6fl5szqeb/rLH+ab5VXvqi7NIk4tQnN
6mXVNYQZU29RF3S5mW1/ejJWPaXqfhz7ofRA6QvsG2zQGHpeizCoqkX5o0SJjz76MQ84zOKYId4E
mjFcKL59gwHgPEp43PrKhOsgL46FxuScFoV2cObfx6ae2b5LbRi8Gd0RNQA/DVShYCNK0x7yLVAR
/uJ9QXag8u26qDwyvRbSZaTg0LGbdCRUD7pbTDviw/XxlvIo0UBFbNnBVyiKJfwBkKxBsegULXNd
Bf1+okvHwgEAU1XjbZV20Or2g0N40awW1L9o7Z3sgVimnf1oB3oZFZk7HzIRPPTf7Sssd0jBxApD
AK9XtCT7RpB4TaGZKBpOtyv/E/HuZdZpaHkGzU4Ld9TX8U+Bvsox0NqU0dQfDV/+oPDvguoYqOFX
E5JY6TN7mnGewVZiGozSPS3seGRuQ1Y+lUxJS7rBG56krJTfsdT199E5M64/ZUKTFIwRk+4xqBHx
CrkgfJBFN6e0/1LoRxwiMsvdCv/+KYFVlERKXWR9GY3oHzC3AB/79/G9Edec4zM3z45GNuVdHKUB
VjOlb0WWO0jC/se5KRj6Q83g+3QjyF7J1R60dTyLNfOWhzqhhB91bDTFQCfZk1q++Al9t5Pwwurf
6dIIHAMhdOR/Sh8u0VBxY5++fl4wPdkGMrfafSEVlRoMF6vs58chOPv/8DAQpzv2ccLTjZ5JbAhZ
HuHfFJbodSuz4rHWj/EM8JmTfl7MLBPhs06kocIRj0h/JQgdSH1PVIau3iNZQR/WydXUEzo/zmuP
Qg9p/EQKIC4jxRvU89rwJuWodXMRSnie/fHgOeN06haiSvTpWuBea7x5T5DSiRd3/DkAer+niLTs
5bdd7C5sd6xJHQhA3RZz0Ip48/oUCy2+VSkui2nRlsvEgFNJJf2G1LNk/KO5xDNliFH2Z6cBkhHC
jbHDnKBStRv6jcfEHNX0CoGwNxOE49w4H1SZnPmM5HKj0JHxqKs44FZCo1AiVU26tzogs+JjdFZl
V6+XR71Ei9ou/S5kJXcFJ6HxoOePFSJtIaJt7a1K+KwYz/6nm8BKVyIX4jzUKZcsWkSnZJUUSto+
pKgbUZtJg/z7a+1TO12QyMCdoqeBLvESYWhxxIilo87A/DCvMqUt1ObXWahhhTI+Rvo1ysO4rXS5
2JVaXAFy9rjXDwyzOt5pkRaoqDgsUfRHct9WTenHtcGdF/RVBEJ4ytqfo+SBsQkSCMLmUv3FO2Tw
XblgG+jV8rssSEdeeNuaqGkv59Lj3ckCj25qTbF33LBicIlnWbOoMwlvGIRnzpXuIaT42JhWkV4x
RGN+Bb1MOWwKe/6TwMnKAExB0Px6fxs7YtPcb0UxGkLbgwXmgmDPbq1TAb6bskCIpGZ8+dbhxBp3
iVBCtr27RzShaLvvJmq4hw0BixEqK8BWXQjD2m7rRZ8aJjwrwNljuxWeEvxC8zQqipxOC4RV1tAh
WVV+KBxRMa5005Pzl6G8xm4DMzmKiaG0/f7wvgXZVoXvzrlnBlXZxWZrDAgvndoJrOQGN41df+n+
FWDPHSb6dQEv9TelcLWCEOZClqRqurpvEr4V9RjDPAi9z5d2cP2c3T6O0CADq3RrFbCe1dXTICDA
Zq3eCmdqOwDVLs4uHGvJBAGHXipbM40eeeCo1nh/eTnTN8VrRHoOjFYN3ZkxugZF8R9IVJyH+PLu
7GwyNEDlluvm0ohhyGlsNw7YpCwJhuclkv19zJ371+PmlS3ChS9GlFUQ4mf5baNaSSeSNpfvXW+B
XkZDGymgVnci/Z2bJeoD29Yd7I3f/W9vrxYMsEEUCyltQ4I1mXzySUSTOWAqlNSD+1ZlerCkWfCd
dH2SqDHHQ/+qblvFoeX5jiNMANak5G9SVIVvwPcQ4q//kOR24C9DUojQkyQzCMmmyImCkSYZaObq
StyFXmPP9SZJi4ykX+Ky84KfYcrbtIKDeJKKgxTBnJTWeavv57owGLIaOgfNgTpVy1C4UOLg/JYi
JwXTPeJGU0HCK50AFE4e43cfkFZtZBV8226znxWw862LlC5NJFFG7VU+Ia0mxvilXyeSCnmGX9s5
BMJbHYjSeCo6UoSswUHX7rhmdbQathGZMX70LW9L1vmGuqdLDYdNG4hdUixmHNtclg3YTwmJD7NN
unVV4r9ArPehpcPUI0XuQJxOQVOOMVNDXoRx1dxGOKd3oeco0zTfrAuVIS6OnHW6QVeBgOaDcKUW
FoD67/wXLOyZPDB1uazaahF/+aldFb+nJ0mqhLU6eGsUJu9iumwI+qKOkOI5A6BCk2x28JqlnEbY
vyTqqX8/hlY3U6kZr+Dq4GT7IAblXb/d3OKGcXUuy6AXGJvFUdLWvsWeCJaQuo8ZT1hPXhFBmnzE
z9Ejt6gnW4OOPZatAkSvD9DnvsFIQG+j/SHPmjpP3kNjR0WNj3aiJaIc/rH08svl12ssWsvDHFan
OofcL3/S1cmujdWCWg6iN614rVSJbTJ3f6RQUwwzT6P2BLS8tT5gTfVXyXS/9oVffkAO382jOX2C
ujV5iEjzw6kRq23Of1Pq0e3/6oBco7Ji7doi/1dXR7A0Z4PYHS6bZUiy+SMUUyIdawzIcMFeF/xy
FCS7giOClASU9hmCUOsrqSEgWGxKq/FsdK7PaCI8A7pdIoYbU4UgE/t6VUtHxzctO9EP9apE4/If
/Z2NFsNUWX/YBFjWJ9YPue/tokVb6ViowtcUKoHV7RthBhPQCi64RIj+wXKxNEd2Un4/Vwy6roV2
g4+hNEbes0BSRQaGi/S90R8rl+/UBTt64HCkNo4zSP8bQtKmo6HvxZcAeEVotv30jmENcW/sg9z8
sC8wsJLiUWPf2drWLy+RRfwIp9qpt4R6XRvQr1T5D2YjQO9Ty48KfMm8YiKTkjK6QFM7WbZir733
sgyOD7nM4ERHeBQT0eUnQaWtTT6UVrWN8K91WR55gjJJx6J0PSBfSDjfCUIZuR2e0Pyu0s8gt6SG
X4RGGzCNWxtrOcPCFgWlyyRwZzszzpOiLV4kLw3rUNo5DKpIjEAhGWByCcHU1zCdMtlSTZQu6j+P
SYqtfOzMorHBa9Gc/lLg55j2QgXMVBEXq4enUcsnQfGRRBTFCwVTRqVUV19+gD104eRrXPyj2kaX
1CMqYI/7RbuhGuYpsOrvJUN6DFRZ8z9kdXO9uRL0lJYP3iBZi1rGiTR/jLQAvRM/aDWeg1/MpJob
+kuEWBZRx5WoQhvsQkKrCo2G6a9itfJA5PUy7c38CNsxH0wtpjOEtQhdApfMDyMkPEA+XbsUcjIe
SvmrztbZcl43b8arTN6ZundjkiUgXn6VQ7ahS583UmD/isx9NIYO4uSYfUD8CwU4TxEpdY9g+Otd
QQcqU624+2YAaPTp/OfnUyH12bgiuPGcig2vS+sHUeqHnQf1pyTkigpbWzJ2LX0vE0i7gP24DArf
o2BQPbvc0ZOw53TgjTzfROdYnTfBr6gpuAUHLib+SuTtofU76lH0WjyjC9nVIjnfA+O3YxZQ5RpA
I2rPXNIT0b1W758SdXK5M9RNFH7r7DoWsa0nY1o3ZXC8+NNEOaFLPBh6M0ierAVdBs1F8D4vk7QX
2UoZ3hU9NNiaZ5JpWT2hp8+MYzzyKfuC7iD2stoY81cnoccZ4Av/vOww12xqwobWQnDOlb+FQl41
I4vFnDb29X21RARFPtw1XTetglbe0MfnoyY18jz2dIkC7oU8OJeFpcsLTfh1NJG5V0JLNq2OVNZ9
FngfrRpKdTV/wqSI9OBbWE2B2HEj+vqxPS2I0KQ7ALqyiJJ/wLqUeQTR0ogQbnGkbMvBme0qGF24
DDZOBO99/Xy6yF0/wh+TtZq6b/VelZ0/Pu+0sM8W51bvdFAo3PlcKeSytgGWym1L90iu/3VsrTjT
Ft0M5qRuMw1JJD8czfRbv3zmDutrZCMKX7yhd1c/Of1TuajWo1fuBZwUU104jJWAH5KJB8wu/KWN
HqgSWDH7Fmq2UnO2GkIKc8gWROy3SE1R4Dh9jTQtwiUILZMyOvVLCy/t7rGjkQiaaaNykobFJorJ
8INQusI1etQyq7zMhHNcgZsGSkKWjvViHLaxO09JFXSscNMe7JetIvOb1oYcbzhqLslMykyZ4Jic
GL4gebeL39+y/e2OjEtArGBtj9199OEQ3PFIIV4TKhypjc/rZUyMjVElxOR4bWNOrjI2hneQUVuC
lQxRCyYZ9jj47M+6NxWF2kofGMnJ0DLBzSDk15jdquVpjrAyhsbU+5ZR8vZaBcdNJ4/hXXyaK77+
n8Wy3JR/pCF9/gnrV0TP9/QIlRFfRkVuwkLeQPtC4yMOVn52V2lBKc8Av8kjxDB+w8tLAeS5sKGD
DfE/nZQxco0MIEjugx1MAhGoDdqjL06++CV5u838JphEN5k2EC3pE3+XYGDaf3cVihWMHCDxmGZN
h1wi4EKp+0EMYwpmhD4mcgrGbDc2eZx5tQI6I+yr/cu9U0nRSeNmm8vkLYI/NRapMbJxf309ai3H
WkuVy21x/eMnt/I8zzELEl8wINEdksiBjor243arVtT1os5rwHVOIk6c/XRRhjeOL5rafulMZfiS
XRfbzYxveSQ10v4HErb4F74FkIuZrVc1xB+svvT72lKrSbf+MRwqXXf2+tazZX0iOt4Eu94zz0Bj
94IaBvSXBtTWlDChIabttz7fFkMO3JcY9Tk21T0TYmhi/PjYgupj/mtk9/Pii+HNBagPwdXlqCKh
xfBgRdrf0m17EWoQyL3lY/9NKiR5EevUz7LRogpwTPViIUV9ZlFWSG1Dy+qoEMozlr2pJusVU+P+
WYgvCs+azaggJ1A2WZ28xoqZipVNCoc2fzEbYD8377U9aZgmJHruW8PiliWIRLP/ygv9RV2OZXPg
yB9KxRrQZKspnJ2NwleUw2qlShZjlfkrTm70gPmN00a/JDL4/QBE02vpGdPwr/VOmNmr4WWMuEB8
E9VBR8amVzNGs+09H+jKf7CtOrlcnuTQseBh7MWKxE5ytlGocXurDMIOlUNSqQy2bhg9ht5XKCEL
I1IZ2KLLXO5QAaUOkBA+I+aCNlPpfrulRPJ+m7oropmHDWjUn6EgxXNBfpSBQUj5XovtfOKrUMo1
Q/8oMa2odlU2hwSPfPgRfevwY6xukiPgVkRitjp2W7w1l27WaT6rCrAogAzKK/643IsmIYzF4P2q
UI8MfBWTf9RAK83qcTPZlxHUaZY3e7YYE8nX+smWNE2dl2uObXYp0vybhAdvvZJvYlwSPNPuYmmh
/Cf4q8O3fqbibkamlSdm+Q7iLj+oaLAgDmfplrk6Vk/cpkL++B1BPbaFwwXh5KPE3ONsEhDMzOix
TYzEzOFGacJVY3OvSm0QK0KLxX37/EfoXIsVDj/FnClm7qgjHeTF6+JwcPWqtP87DRRGEyeQBdgd
jfdJDDyZhXLzmdePN9nHtq/x9BvB1PSNagrUFpi1VgU3JXgtJIW6I8cCEyAm/zHHSMsTqmID8Nnk
Y2DIGmCnoc8njLB3vz2DowP7vZ/WtWaXNYQtZ81Wp/ZCO5JrwFJy4/OvMVOy4llueEtAI/0dA845
p4o0sWbY0r6UxeT4n8TTu17uZq/t0nGl6Nh9wTVjM6FseUkRYm3fJf5FgakGTHkgOL0e8v48xE4I
+2FONHxlu1AQntluW82peI8O4FCjyPcvBbVqO596hJ9I8Vlly4a8++8OYg/ZBYSrXA2rcxeh92N6
fwtlmVSBfSO5T8C3K8Gz/wijoCBwWAUR0WyHEyrCMqsAYMV3X2ETRLW6ynEx+TB/tY2y7tQ5KuL4
0M8gHf3AOeyX8wfXdvLBxwPig7ejRUTvlB1tysaMGWW7A02DYMBg/izgL5ZwK+QU+Lu9Ixve9+VK
wiwAZ825uNZxIBIxG8hD3BzixbPbFxeQKtBXE17Oe3KQ0uvT4+bxcQuDOPJ0rCMs/NyYwqJ+SWwq
kemOENUFBXwGm40a5Xs5/8E3mNb5mkxQPmfa+0s+nBr2TGHXzq2REBg1jIQEofuozsvLgHiopnCC
p+ljihe5bGPSH5/qvYgqXj0NcDj0/2ub/Ef53jSXrg5ZW+TXnoiLe1Y4XgcbFUvb73nUS1fmbkig
m+Irz7XWHd9rMzGj52DFx5eeSpOWaw3+iiMbD5UITj/OFMpYHlEDVP5Ad5aWenwWpHLPqI9loz4E
TC93htWao0ZceAvqigb81Al7SPqbZH57uGE7iuu3YCUL+P3ofQ3VchuMbKYG9WbRz3iZWVtwaysw
fw00RTK55VLMjmArdavfDVIM0/DMkQsHfi6+r/ycYvV7mOfxoVoMLNSDpsBPcv10jJp39ni9Pd4X
bGpzM1DQSagnqTN0ZPDsq/vh9jbD3DbKcC4lvgHPqCzDbb2mEbhV3fHDXB49dhrssMymDGnkGP4x
73BqzhhuqB8yeHJaUJFisP/mZont5l/Obl5OdxLkK+cD1nUYYvZD8yvWuzFCF8XA+yWiAhqWu1fa
P7nUWhruggFQEyZ7qJdvWi7G7LATPj0aHn8UYhFCRNVzVKsLy12jJkkQwmjUug+7gOp8NHXrCqlC
Oo1MWNVVD4wdTHr8TAPISz9t9uh4FWx3e8unOZO/Ykgcyu87D45hx6A0iuMYNbV3y1x95wl9R5ix
rptP9Qr2kCmTLGEXFG/Mjadl2VuewedismAQSLyPNMWgf99P4+/dXVRvMn8K1/vL9HZyRI21lCng
4w3Yx6ypbbD49JI3ekJNu/6kztiwMCTh3OI5zxISRCokIezkWHr83US2SnBbcpMwuLscOgPWxIuk
1Kz/CE/8pLg0DPUaQEjrBL6fpfzI19Gea+yXq+P0RbWjb5OjCi95kZcfccerA3i9+p1HqH+XAL6N
I/Wu3lI7c6oAzuYgj7/jUpq9gu2zncvr0wxzJzjSA/pTZWorsmsOu7y8r8Ea1RtL24QzNyZTLuSz
toWNXIkJl+zkqnNHOS16kPmMtzECIgg0B+o9+/nSvVaZcz1h05/Qw6CYtvO5nEF/oUgK+2LZdyCu
D11wjtojspb/hULBFSyOQFn1teOuXO4O4f1SMYvMSe/vVHUNbNZqPWvjalPY7adNpjud2dd6Xgy3
B4Em+tjF3Yw09w/HaM6NpH52B/PpNUm7MwPc/biLC1o6yud9Fy3qBQFJZDiHPNmkddcniNF3SKvU
83vm20gTpib7YUV8o9Ya1yka5DKgQNrQLSarZUJCwO9WljR66hM1anna5zpxg0+NDCt/jweIJ1A+
UwV5GPTmGW3ovvphWOOXQ6upM/cv1MFjfdHoSw9PGUVBtZXZJpxdt+N4GmQVS312GMPMlYutr8Rk
O6tW3eLQyw/bX14+Ik+2ePr5XZ58ut8/abUZDH9z3QD4tl5UfG7Hx3lc9A4ewgPPFqTz7fyNp0bZ
Ev7OLMaDbRoqH1NmTm2I8DA6ZIoLQpLVoQxYE+gubBl1ygUmj42vx5KXHO0w+RxzjFVm+XSMQ6Eg
LeeW3F3AehtXkhVxQvuvIdsshfa+oeQv0TifyS6EvYvdwB32uyk0g8LyZbJUTtoKIYIvuIJg3jbT
rMlPeo2VkPM0lpO8VItVFYczwcWZMBIciMfvgSMGkMmYuMLZqqBFoGTyEcTC0hFjmheeg5k8QpK5
Rp+x0609cR9u6jM2b8ztuA/SV+rr5fHRZVscpbKq9hIIPJuwZBY8KtSP1dI3sEJBCmoKHK9jJDk0
ddiWt2rT5qfu3e9hoac9VWq0KGa/TacPxLRGX0NYmDdO7qKoovs2JuWT+meMTtVXt2lG12x+t0Sp
1pZuj29y/tEjwy+wFZkmaKT+Utx5NPcgeSwFvtDen7XsscsVUn0lif1W6ByKqxuCBLXh2H8qWSJQ
mSdmXa9vfWtFtjsyWYxHZ1nRlGF6Fz2PAyq6+YL8NvyDffu3zUVjA1j5VecE9m3ZKngzapsTSczr
fdkHpCRLRe9aone6/pKX3ayOxHwAI3qsy+yQwHxgfv4kDkDJGMmrmQXo4P+p7hJRxLhDTlQ4mAXt
Gld4CQ22VHWaX4IC02yDQx+93t6YwEKJ+Z0vBCiMU4bX1WZ+/TScdlb8M9j6F92GJQ6PfQDcns/+
aZk1qi1FWfj+AWOlfEYj75XlhEnrrjOA5cY6Lleghk+jikE8z7R1nezXUm/8Gj2QD5+ZbHFHh51M
OyA0Dm/i652jPGhVlGuXZGH78Sauxbm361hxRERUA4QQZGsTt//I1fX8RR8pHf7tskodfNHSxu9T
6woLHxCPnEdBd2e2FP/rG8zSZrm5sN6ZfOdyhD8akTCvBbXsZ5wws+KldnA9oK3RXw9mxNNhMD+y
+aVuxWzfrP9quqIHfFoGtFEwnA8+GBb0VibgZ6Kwlfj4MGs+Ojk9qgDGhKVfNFzLqhAkU/VcQFcA
EEmwytoDeXcpivw0DQAMJyyrHF4xKmjtA1Iz2E16Y6id5lqPTM/S2EVaxzrMmu3QNioqswqO8tMz
ODJyikk5YNR0E99z4gLWA4YhFudvAt0RJzNIUTMrhE9LXVNhg1jwZiWMGjPj4eco0CTuOzSm20rt
tWwbggH9g+RMTisDTHmURAbi4UYMdwKShQIe6cQBf2zWIWG2Ko6/T88slGyrxTi/hofSNQlNLL7L
yVrdFDGZyY7iNe4mPOLZQmLJmPXVRf2UeqNvpgOZzHIt0zf+x0KZKf+Srd3oYNvcBtER1I4wLOXe
IA1yBhEihFIZiyyRtiB6ZD8biMViTHRhj7afuW1fheOiXZWtxcCWNRQyJBfkd6sPSMI0590jCmV5
JQS3lkD7FPKJSJvq+RP4qtCPCypWOQZvvOxdeebbhYczma/3voFugCUKyVVxPUa+HCfTjpOTw0mV
VaXh9kgcHOzgomVCXlWT/vkMlYYuwpS/fRaODL5G3L1Ii4fPJOg2Ge/NEiLXWdXm9K0BN1dx7RGb
iLM3mZdpRD4SNzRvYqTnPzlKenboAqRxoeK9kM0T63acEYPjuSSzElElCI3jRHclbFexw3UJdD36
KRzZ8D5/Uw1rrBjhmkrB8tn0OA85kH5uJxM6ETP6ZCaITra4TtKWDRctdjrOzEFgO5B1cWBO+g3Q
b1as0CiVdyqFvCBrT7Guj/e7IYshFCEnzxeY0MZ+caO6RArCuTeb5VafEjZ4qE36DIFvE+xduZez
Y6sKrQEXaZNBFzIT8VxwtkYcvdO5p3eC+9hIBrruxp1Yv0UXcO4LpcuRhocV6P9cMwNi3krXEKOh
wqHmtdVMLP/9peuv3QmpX+/Le4m2OhxkadtkhmIbmTTI0TO9bgmfeWP/sZc2BAY5zgO9nZkC5bdI
kF2SX+KzZkvwe2u9Z84BvRb8ktpYTEuszhLfYp46mQUNmv1CXT1VHnUgTE+KL0cjwXHsYp8FH1sT
sghm9mb+nSzKu6A5/AgCfDhjINOoWyhvnvzY1/XmaLy23G+g4Rkx4gQNr8ZcwK8d5tofLOxoHJdh
zNAp5eysTNSb1Z/W+mJqEUgWWyWTRPq8kQBNF4qnMENbkcdtJHKqVIyj3fW0+qcXX8Eaoa8waE3j
41bhHWcD35oGmwDuicZRFXBi4cY9qekMBznvafwn4HAHo4x78V7utkFeHjktZbHJrw+VjP6ZL5K/
0VfjteF6wUFh4QCYzX+Bg3TkgrZUgLmp5a6urgbWhtXgwwZUOvxFF+S2TWY1YFuZjGibsTKlqaFx
2stn83z6NpSJfG2JLUCt2QCuuGMIxTRYfHOBLjBTrt+1NxBMnDqOpL5fdwPBpvRsp8FZE1DY/AqD
H3twfkWPck3Wup91sLiqRi2pxXM96EGaPSIORpqtTsIEeGbPYL8/PINv4lXF06Wam9CIkTzQUiko
5PW9SwZgWi0oJjqCNQXcTBKOU/9LzXloicrVQ22YIrZyIpJFPOaT6jqa+1kk4It5C45untGqoxao
KbEFynLpWwHDwhwlt6Wg64eYoPoNOMr0wJtQiZIGD+XCTk0MuODJGz5S0XJNBQsUH33JNjObE19n
Bv+4DCUcetf7t38F1g4YfCVux6AAawMqrkatDfjUJZJA1ldNdS4gfxYp9sCQF8AzAUmamohLEYkU
M5OwN5AfnYGgUIkETmugpMWVf3AczRTbBooeAmfUGGukjrDMHfJLvF3HOEBUCjcxKqPiwG+pFGcz
mRqOg2krfAHeQtCfieOYYNRtNn4tBkpS7r/anhI+x5RLEZY0Z6kEqLU7EPUgDFVdWC/BBIaYXyvE
vVe0Pa6YIW0tk/b8ev+MGhGO2oGjY0UkwPBBM1YC1HtGRS4SfFZBy+0HsoE99a+yo4hYPjswySav
XBBcu9G3i7+RlC38SRlGvJLrKlOCpSpO6nw4mcYxGNAx6pv26/APjktQ3p68rOQ5SJg5L4wLo9nf
csEixw6Hm0G9vLWcLlpZUE9C3qC8MTkabjTHd1HGhKIhB4tASUhAazkcAh7Wz1H4bl/uwcegk6ld
60DtAvsm5xsG/0f/p0FWQgk7Ful06l9LYcDuw3HwtB6cHc04Zl97a2xqFDzNr5HxpTKAZnyfRKkr
woz6ZKhZ2Z4w8OszvgsRIuxwVWuaROVmJP6LtQIf2bFws6urVWCkgJKIYezv2+ddbrcIfn8LZn0v
PwAm5/nBz0rWm6GRZORoJY0/dD23Fdr2FdDtRF2rcSwqixJANKaPZD12NoBVEMyXp8oKGPEXPRIa
K8TNFgLpPg4uKnsoJmdYSsufM8uuu9vx+e4gpYRK6gvQVMZ8PMuf9qsGdsjlsHsui/vGPfMT58Hv
u2TR+licCv8HCAE0lOeXP+qgaaMnG+VEQE8vaTOAqao5Tl3nbLF2irAUZ8Na4cTJlNRVBbDUiOXq
wGsRx9+24IY2WwI6s+IMqdMfxQaA+WYdHgzAYAVdvwHgdAu+KKZJEePg896fuZTpZcfyjhvQEau/
okQwkd6OEKS442OSeB8yaCc8hz+hE+8JBkmytXIRHN/cVzgedwO+shXTpxTW8Uvv1hu9vtZUG/hr
E+FQ824yqSOoZboXlyGqrNkUo1+23fLyODLDLOcX8LJUspJCLUUsmYE+goY17Llxyy/hTum/LGAA
Cfvzy6e3LPb2JmuTiFY490fECmNLziT6RwmkzdpxSOMNxPLVo2y6ZZ+N2Pi1muRMhKIlIseNAuNw
2GVjga6EQYjYTng2jo2XqXZm0UapMr3NwJg37CK48H6hSQMkYkZ3BPp/Z6Q2SNm6vRqBXj9XMKDD
E6yXsoBcu9bY0z4YMNV9TjtMpPNvoms2GOlZw971b3BvHclKg4r40cPbjcRybEQrX6CD+0nnuBqR
LrIdn4mAfB++wZ14WXbZDAz3NvzHYxh/3PWSnJBS9hF5iy5/kPBxnR+OTg4CAksanWqKrSmG/EPb
G13kDw1X619qO4i+zVdhWK1SMuL8ViLeXoOWlXca
`protect end_protected
