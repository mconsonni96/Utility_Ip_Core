`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
lj0wRIkCdYeYte2f7QabUuKxzJzQgWPBOu9oFwOWGQiNGeV03WjeyXjbcqFjv8Pa90v+vYETJ5as
pAok+6EYU0S1NA2V05+uLGv04y06UWyXck0BGwq4wTuXpDBwIwXoLbZ9vLbzlese80SWWKUif5gA
b3r0iKRIdp/yFKIpYfrD/NOuyFbN91aJnzwo8nWxITIrQwpjp1oz1ut1ZyLsmgy2qhGtjkTRZNI9
8idDO+6clyCN4pGC3Go8Jh9Mi/2LAQtR46m8bn6OyYnjkaa3Of0A6rGczlmsB/s+2dQhZu6qhsXc
KUVYWs64Yv8iZm02kOLWEljBzhlUfKUnPNSK0g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="voSqcP6qAajkbrnV6DrfrI/0nsAdQFk0UsmoX2NjW0A="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20656)
`protect data_block
j/V+61BFtFK+a+gvFft2eM1/aigDJ6iUg1AAKJQx148OZDOZYrgErvyZ6IRozj5fIF6ePNEFNJg0
L5R/H8gS+pVnUqcxLDqUkWOScgSe5hNaHksjWsJybSpOo+YZ5Jvi0+dOKyoo0YPdY6C28bq3huH9
TJknN6RPHoVQU9qG1CJpBvzfx5JdxvPWNW5G/n1X/Nnk3OjT0LGRUHqdtt14W+V9tWcfum4pJ6fr
YY1o4xZDD/vOmfcr8bO1SuGT+NHd6xxDLMta0ClU++hjJumeV6H8+VU9r+VdPnbOur9T2P01VViY
W1vQyqJUABW4/nEf1rbpXmQjP7zGBp/orDfC5zuBJiNrrm5wVHl5QTFo169uFek6oIiDOQi3/NYJ
tcbfC1noukevcR3d+p8L74DCgCIIS/rsDnJlXHr2p097MZ+ApWKItfg2ny7NSM7YcoWfXx4B2vo+
/LLBz1x9q/szBHlI2j0RNtUN/6TElAi/S1HYw5NUUK/09vbUo6ma4XQ9a9bMVhBJ5mQGEBRM2CDh
PHoRpA5MuALaYpLfbcVlFThY9GmSwvAULnz2SCSDtDTwV1w1DSxioPL2LQIIYEEm+LevYHNiN8Fe
FoMeEao7X7Z3pLut1Oht+/9JHz4Vt3cZsc2oY9Q6Lm8MoJY0Sc4/XuMJWX87BbEbH6zs/Ehr9QSI
oiFGJyVFuBH1UN8I9gPeZ9ca+ddWmB+eZ68JmV8e6PuBW2uMW8jBLL6wvVrc/d0i4XUdfJj8wm7v
+8Ydvmeb+t6lDDH9uT0+KYllwhbiD6cUFwLPaBrEbpdkVjO7GPSlHIfzAm3hU4NRja79YJ/WmSlw
mvubiXlrv6QVKKD8PqJhcPS9inZNcpnplDFsvERPOxNR5u9AnlGL7OLp6DcjfaXoVbJMsT2xB8i1
BCq30q2Em3HjYUveXVpg7Ed8EFvPqXADSjQYONrFhfihjaE+K8Rh0E2k24+6D5wj517hPus3Q94M
dWe9x5yZribGXC3VwEJZUYYDZ1TgKk8/58Aw8AwyiHHz7KbQQLcClHFb9MVfRjfp132xuyoi3AnL
n2XDnCv4kBgopfBYPSqQCYfAZM/2/7tnwCZMyW1Q+Pf8/379lJq8I2NZmDrBs1hykiJlT1ZwNMPc
zgyAF2zK/rmYAiDIrV9dhtGTiM+5CanA3eHBOA5O3mIxr9p5/1IWr5edBrG/H2mqqP13kqXqc0ve
F10q/thm8D1q8LElUsTIpOVIUFlBROyAo7ObFA1r5ndDgrGNLsoMIgsrrRfqrD/CRHls1Apg+nJl
xWojty1HpZ+gzMV6EmPSz5Vo9gM7sSUx2LIchpwuPoh+tnWjt+ihRZFNFthYflzQ7bhrzp3HQm1t
5M76pNFsUX4tNw6nyWFxY21emkiGHkXzrOtwa9u8myVOkkL645hV5n2BrP0yr6IMvQOw6MCiGDcU
BlKvILPHhHLb0skBum8eCFFDEvj+p6lZIp5oDFG+YRMlyE/jZ+EE2TpysvPC2/VqFP4yMpeMBenM
+tJY3JWt652/jNE9VqTMUhfzdaW8YnAJlA2IkQTT1PtG335dg051qHr5Xvc3G3PdCqzmRlKqFh/y
bJOXeX6BWh5g2n7mSeY1tGvY6ltBnNKYslMlC7Uh9eFFmPGSHhFV4LthBif1ZcvCqJxwaf+ZeTUG
YJ+qks60tA5YtMPHygwrqmKleq8yKIIZyKxFImJJXJAeehJdIDgiWTtMrme/wlS9dYPBaMj1b8mV
e0Ektri6WkbcME/v9TaFclhaHUWcE0KU9WdA3aMV0lT22/QNqg5ieLGEOmzo5kpNGjGCTyALDh0s
XexOsprYLBJ46nFy1o6YICBCYqsAy1lKdDRtiIIYzNsM2oYvwbBdBXziD7K3h8fb1zDiVWQwktzO
lYx2TfoPccxbhH98QWzH+QmFYbltcDCBRo6efhQoVm0hRoXySpgz+pgtulyhZL2+vsVGia9op68Q
ZL+hlh7qwBm7v2XPdptN/iWoYdo/ljjonSbHWDojxvCy9fWx7y/hjzsVgeHna5QkS2Iz+pCY6St3
kyD4euPbO1mbVaUX5zB/Rulk8Whz8zT36i68T7igE7BrqryLdymDd0aFI3jO+JZxq2jy3stPpYfZ
k3oBxI1bBwdQ37heb3aI9rHWcHpzPzHYrasuc1q+Zy+BG5XPvwu7K+JcwbWPwLPnpCuZSwZnCd4N
Mo0AmCcGpbL/dVJ7yTaiZkxw4bhfIRYSMh/9JqsrzywL3gQp88tQQDaUYr5VkGvHVfeRmQ5GJ3Zi
y+yff3SLn7EX/h8wWWis7b81oNStcmloziXMQp/MGggx7qX4YOdYyxA4pTGrpDY13NVyzSiTNOC+
FyDosBi5ftq6+qh0eMIoQgs5jmTkzYwZbk3LfqDUKj7G/P9CeMAeFzVPREnFJaLAzbTw7Psg7ggd
e/UoR46ZS2ha1aaCYDhVJj2sHoaZeeMDRpRPyAihCGeJ/MjHNPnoAJ9FmsKW4VE6YChLfYLMBs+Y
l6UqrvAphizNwpRyJi4v+cFQesIuvRYX/RnlW/Pg/oHbWgH6xn15TdjvE0YPuHeNk7CYhfXpp2P0
GUeJi+RBqwtrQw+MAZpBObSTIOeXL3gKB0n4uwaaDnWkRzL8sA7Yahpuba4FCvEUwcSLPdpEyIEa
lK1EFyZY3jlS4UXERFWhOsfGO6yG5mtw8WXFPofre0/TSjcGpCXhUJW4AW/ZJRZSA1o9/JpAnvgv
Dy2hB7JIxxFszlk3xLBzbF5QALRgNuyBoRkBHFHAomny2sU68JZONHks3E3SJ+sLQ0vkWN1Agy/f
JobyshruzDaaa9oiQxVZvGXt0v4Y6a/qeV3aaArNKA5kwpg95vyBeubH/kUyNH/eA59Qfmc/3v3l
DWA129ajOr/viipl1DeXuNMfLHpZx5Lbe79MURrC1NrekNyfgs5dsRUbpT1dd50KkCRX7rRxUlk6
RWTDqROuSHo2c0YGJcH+Cz86/+J+lvgDgoTUnWBAPveuG39b7Hz8xPDZkn3n8qpT6b7PJTOWPpPe
nf92fId72lECMGGvNStGLRQwRJW3EgQXzAWZYRmgf/0MNGtbt5ymCy7FWB398xRdv351IWcA2R0l
MJH02NPE2fBPpsNZn5ptMxFshS5+h7ePF91iYqAOmke9duor/H9YN5Vu50gsrxUSJzx+E9PUQbZh
ULIoBU9l+hc8LxxMAr43H2gSgsQUGZOzb92atjtfoH2e4iYyaQpMX8ZtjpO/o3wMluycxtzGEbpc
0GsEW9F+EkLAA6+XrTWjeMt0gXII6KteeiCbiLZhFNL/hJAyw3Z2qWtqUB+j0iEHiNMwDg/b1cJR
yzGL797PDfF6NFQhket+AFUl1+dIZY8p8r4QbifJ6qNWUPSRWKLk6P11G3AxQSbvMPwXczlfgIRQ
QavHShC4adbYVXkMLzQOq6ZIFG35ei6BJDGQ6f7iAxIEBIVzk7914toDfI80sIql8vAOmg9a+e7I
1T8Tmt1a9Qmsp3EjB8pUSDjyKwfnCKUTybvq40W2b8muTnK0Ypf+95N3m/DKnWiRe5x65Z8wtv3z
00cfGKAb4of4mnvL0eImq7H9k0A79VUMqC44RX4EWGLiGyoTc7hJg3AMazM8fj/rv8Sy2aAK00OK
wxU7OIygSxbX3ImD0Tr0i2PpxKA18zU6EEy74BY/KvX9FMJsGcXN27SnLXKp2cjiBkGqQRgDt2Fy
EUZF2MaSskLvWjDh9+F9BxVexg4uHYpB/o53hgFW4YXHLeIy+iBQ5eXAQ4zo7HPlkLY5MC4/R6sb
71A0nFpxEj8hFti/jiLu2nBwO3WofmUMKVoEGU9quTD/v0qhJeh8yiNnYNL8cAq1JGXRdjvcpXbx
tAnGYs5sOrimZHVBwg7cvyWKOFpCw8mckWW12lUvNOXltjq9g41uwEQ8s9S9HMTee503mQq0Sn5S
8YGx3aTpgR7lozCh+OaAZTT+VBGKLo3LP/gdVBZR/QqxgSSvJuK5IojyucG8176VE2CN6XRq/Vmb
bg5rmodP4lT36pW1hBxBSMLkOG4LZy0Fkr7g2ycr+n3rGgpYqUvhc4r9PdrHncKO50+MGKWz80H7
KPhHn0hrujb6Ir28oSGDMWS+JR9gGL8Pg4nTgTbgSM36FC0+ViMPhbi/gTIo56DUfY9hO/RdahZy
rNCqnKUtyf7N5PCPzWTyDsQRDKVPsY2mupw/aTXrjwfgiKLe/aNfZezOJfWwNtrnw+F2IdHp/kqh
+S1kM6aq0MuEwCmXuJX6yDXb3S82F/fVQpXfhezkV6guFSOxHsz9H3AwboYLQzPzXSKCiH3nfqq0
wL52VV+h8b86i9Sp61p4lRtEMqkKiWZEP0FJpI/M/wRtj+Oqtl9T4XnFwqxYEta0HzaSMJi2qaKq
VmjaC5RIdcFoe9Kba7OqEYYm6+jeSimJkUM86mIgApJFCmir0MakkVHACchDX2t2KeGuaMy8JqmZ
V1UGzKccHgFvrSPQ6UOPkMkE8gF5pYI7IGDuyHofL0PgSEzFrnqsNJa+oipljPirY9LRxFy/MxnJ
Lb2yb1Yg1DCaS5OcLPyuSbhc5GM8VxrpMnYn4GYlexLqcIyWxrAkTOIjHJU8DKafGlFSFbdZxsBt
OTagHO4GUfS+nsu98WFhGhcTLQYB8qBGrNCrZy3WK36GK93pjekWUF7SAxWohReww8RNYhatbYi7
J8tnxrsqCADlsx+Ox8cJK8yYUTUYllWkwIF8gr0yiwN3IvF8LxNgNB0AiGt1XyL+Rd0ZtE2xA0iw
AnV7WviV4oceBLhMS52lXEwXBfg9oYUTyZvnarCcnK3pKSqEKoA89Ab2lAiRA50GNXMmtfF7HZjJ
XnNJhpRHpQIX7W0YlFymolOWzvFdhtVGhgOQoSzMXXNnVofZ+u9bYcB/+F7Nw0L0H7HZIyNNLgoi
W1vM1oyc37UCHFaux2+m+AjKVdlpdUsnUOaxhZt16wIYrei49xCzUDl0lIT6R0jELajihgpZ9fNM
9ZUtaf4Sc3uT3gXSy6+pphTS4O6xkqz3qZjwWgYuH4KgUXJAtzAHlowLMjZuqNCAIeEMFM24GzWC
tEls6nKXUTL9xXhu1JTB08rHEHHVWJfQEun31sdx4KNFtd46QtMugPBSwE53UVwo755OAfoZtsAp
GlqiIZB1YjOAJZ+ZTp2p/CHf5DviuKV7a5jr8JTZtZ1ckiuHytuLpwNvoQRqWiPGRxUkQ7hdW2e1
Er0YoHN3qIJkMtAYoYroQg8XGH7NOSviZ2TLmF6Qdc8qhrrfI2Xthj8qm7cQ2OSR3UY97UldgNqx
FZNJAhe+PNWS1vVQEUEdv9R1tCh9iCGvZUXOfaQGahnDJae66KUBDgc2Lyq2NmC0kcgzCX0L9eFZ
B1PND7mL6FUvUBdtak8XqfSMsOQbZ/8FiCwNhanM6CCq8vL4V1C55/itukhbVKX3gb6VI0Sw37BX
/aSNkj6UH36CuAWMwF3BYhExUD1dHpCPNCnZJWVoTVLI9qo1RWvZNh+Voyv0/1vw3AYul/+lt+G2
fg69W2xaz3Omnm+Uj765nybwNxwJCT6shcaCMJKMBMKzG7bVspBQTSSBwluUz4EASUuSsg2ooMJt
m5AS797XDD52iA8QMoKj/1woPuGm6yQYJokIrw2SgqSJpI1M3uMbWzdkHzdv5fa3HnEvTcRkUyYD
UBPpQ73oaejXinFZTizj0tQ1uZLLKfDLkM5rDtln+y9ltSBM9ZIMV0BwTcRLA4V6RW9BWJUmUb5B
o0MAmGVyvQoIYNeb3LuOzYOzCHhgVi1LRPM5mXrQgbQnOMBnnmo3XknRqNZXqdXE28H6zcdyU4dJ
otRsJEyjvjRmHYua0PLq9njUtS9hUZilx9ODdZTe3pZ5LY1G2DbJCMu6OF3QC6ADi3Hp8ZLMKv3x
hvUyPyiFVjI0sk2goO8K9a2bDBnYngZvK+ud1oh3IX7DoDrZLQ2cf14iF6F0v3QFsEv26vFfau0E
FMVIhGIQnpcFGIDtk5bxAEjT/OOZ0eG7TWzrrlKacPT30THmQk8867AdTa/AziYMTmS8SLoxVt3v
7oU/v/fNt+d0J/X5DRppOh44ZoYGEp0dhaBTTRuojnNTFtgeF9BeQJqLPTwohMHk4lcD/D7g+wVh
SG9pdegRyEcOhc0WWDEbrpNcWTbjmaTomAK6Jz4KjI0ZMFwoji6z8C9q5qC/6600ZtkJw32/fdwW
gurje1Z5pEPWmkq3TO25arfsp+z7AJFbdEPClnoVFXwwtDbM+G5I+8HoJi/t2ZkbFCsjQ7BbJXS6
yoWUp1DbLx7XxZ9IPZy8+iHrUc6uveeHDcT/uwi8XplU3T/f6QYYUlsWynDaOC5Q1IT2wUz8RAD+
P9tJQMM004tVLh6nkffISRK6L/gOQC9F4+5ZGduLW042ZODEI9iJg23PmVo2OKbSCFryln9dzG8v
BtxiCs/kYI5ikzxHw/T9bOFTB/C8dSN19jVU48sv2HBtG3LsS6YVPk238zpBj+CkaTfhBiAzNL5A
3wq+KCPOgEH9C2K0mFLjRR6fp19/lKoIENZB+QhioyCf8mNfYUOrllMYWlfUMCXdUgzDhTeZUtSj
lj7vVlV7dFduBGsQ2tOmbnfDp7Fs8vSxW0NULopvSx5hwwyt6CJYGW2UDa4tgPcWrZuMytF1h8SU
0y0m/N2sDu+sPeWLDAz/TS1nvykW3gaMIgcKlwejmHW1WgyHAY+6Q+TmFjPdkBMlhrTfc2Cet3m7
0V19FyDzXYDD3vfhAlYPvLTDQa4OK6i96DyvgwFFneFcAm3EKs6f+evSaEvLpLyf89PgN/HVhHBE
ETcImJNM11V3LCdUaDH5SbN5BeaMMPyqoqCTxaMVd5Dh0mMWEZlJtsRDuFUjq4+0g11XpShA1qYZ
w5ute81+XjtLOWRqMj9Hsw+jO3mwQjaKfKTob5SiqswIBfi4QlKEmEyLl3iN5OY4u+F863snj1WH
LQaZoiUr+XahBp8D1qPsSjn7gaRfXSQl+/EPUB4uOStd6vDdTFO8UPonbMWx9QLQhOtqOhrPQh97
pFLjhiQBS4juTUEW72PVxY2DNkpDnnXXjruqAehqSll7JzETzmrJDUj0KsATOj9qX9UPKgKDq4rn
1vsn56uHxwLmnHo2dvL2WkpemIk52L3Vaq6QKDUG5IaIFwdHzDjBQx8u+ELx/Wxd9s1xAkfsdumt
nzqo/YK8zR+e6TlRypUXOyFyYk6gbUJPsSS2rjNh1BN+E5lQYuA/ADDDdEBxOlbGy8LpNM/UvWTU
aYJpzb3sWyrs1xzWXufK0p/vIq8OSt74ISYh/gwcwsVaHp2wnGLhaSB53TXkC6P/UTMFsRuDJv8S
qqsMC6Mo7cDdKw/N3fTe7EqmpXKl7Ft7Meq5dKDNhf97QpnguDCCfQrLy1oMxMQC94UFM21txZp5
76pi4kSxNz3FLNmB157yGzx7QQXbuIHaDUSbk1GyzobNKsIubmI8Tlwp3g6ARWACcYqr1xIxyDtp
29twzbUm7q0JI8GMTu1O9ICnWg6mXVCjFMwBoyGJr/rVMk+3rpM8eLLKRIAIhtdXjoChfGyJTEg6
UX4LSpPqKxu41zRzzQuLRKTqIm1QcZ0CS/rhlBccj5NhPsZdjAoV8LD8kXbDeLAxtwq7nLsiQi5T
tKQYiVKeLBp+0VhrmApIh63IPIMvsQ3agEDGBDa8u66N15YG40vxMk5IcPt1iJzcXKsns7Vu0CXx
g6Jx1k+OoFY+YLD2EJe4PieVSCgP7Qz4/DxWwE/0uo8l4iliQIxMHWCySAw+1qyTodoTU1DAqf8R
1D9X1UiXfJ5v2O63NCstMV64E7hLEX++PJumQWa1b1MKu29RoAsgGbHPQPm0J8hyJ6gHDyOMNuWV
+e2eq8OX+pM4nQt3C98/FuVlccbnjrgdWIuiYjQucxGHVViGAhwynOkxdmCcl0zuEgfKGZ/zeRKi
Td2PUHeErivdkNkF9V4TzarW7wA5rwBxNqwliEPp6bCQ9EUCwm1jX0H+OrddZLXEjqO9vV+bU0r9
nXKhYKI2NxORIyGBjg4fPVwjnnPskNhRmcUTbJfXSKqc9/Xdf0TE49t7D6z3YymqvfLmoVwuBwik
bDZa8ukZQ2y4s/ZmcivR//qlqKdtBm2985Pu9HGSZCjL9lvRF0X9X8o/RpMWWfik+Io2m3+0lV02
Zr9aRuGO+rDKd/vqkqFMdinrIBWFXstDSRBXKaFrwywqbh32DJcQjrF3RzTqvGLUMpIpktQj/5+G
UXRpcNlOxSzPag3FcZEXo/92l+NHlMEAmhFqGqSALaUrm3PSa/IEn28/X9E2Q7LyQQr/Ks61d5v1
CnWUXTU0iwvK7NtvrXJwOXEAWb8tfyauDqCR/J+KZgjRIA1Qn4YtLW8poN39ApRigaAy2rZzRJJY
Dyye8LcxKhwQa4InRjmAexUw51u14ABjoyxm4iDvKTJP2RQfSinbhbL0uQ/xdWxNJMiyNjYmxNLF
HZtnjBCschkR+kw/KrrM/WNHS8YyjPN28d4OEHQtVBdH6VisR3fB0Hj/ANGqhsmpmlU6qNF8TMp9
LeyqIkFo9qA2iigty4UL3GFjZ4o4JfRkBBwgR333gTod6GovOVdZC9R56B6g8WLls4uHoV5N/yEX
wDxYe9gTWwzkPqSNhr1N0wCXR9bo50HapNj/GbAbEtwOXujQDCfHvffLNVZxhYE1a5YgCG0rdQ19
VLrZTgsCRCcSLdJloOinE5e7bVHo+VvZSg1HuBpSSyyFUeI3/4VnwUEbdtHHnUH/9pJrTn/fdNvY
Dz66qKZMzwME6scxp7R3aMr13efobNTxzf9N6KO9IMw8gcdaJmDqB4prX5PmghDd+q2DSW6LT0TF
E1Ipdey5aLc8qi57u/hnxtT/xVHdaPmwyjJkWguYscJ/GiNTJZN+a7kfqCriZmWOcQ8EPQ/zFGIm
3seeXjh97JY3bpeGoZcTjBiMKMseZiQqrJmt+Mk2bfjoWvoXtL0lj81NrFH6Ltt/BUOBGGs5m/7z
Nc6cBGUxzrrMEwIYDZCRAgrBG49+mT770Gy6ONcfikhq7RA3vf/rO9y/4a6v38hlFOpQmagajgBI
UYPwBJB6g1fYzwlSGYtw2eVWqJMI5RKHeVUxYjro8uXQGXn8akfTVaU5HY0jEDTdZ8DfhGmfKp3G
WvzpGSNOi1uNsco0ErqaKFfHuWELJMuWiyOjDhq341sqo+jA6ENS6TbGrfePxrzAaB8FqpBRLmnx
+xGFg+FspL2+KbKr21rp4NCmeoJhhk9gg3Kjebl5AKjzRhXe1BwiSHRg9vwMO/JI7bN86FOuvQmn
hcwBO0+jWx8VyZQK7YZGGmSo6PhATwv95n3YK8zTut26nzPBB47owKTGmR6HF1ZEEphpbKO1N9wh
XVL2gtD0ePy1mNZDP/VXj3REuCwtQ1C/B9L8YTdxbi99HYm9oY0KokR5qnNmi42nerImfqKza6k6
QtswMikpgj0RX0gX1L/FRWT3bxYnL7w2MyXT3QCmXXliBdYThEhgGfIeAb8KcOwgKtmRpb7PiS2C
+dl9q4BcDHYOW1f+Jeq0SNK+J+Z6nh6JSe1lmPPRClOjdqU7ytn1Ij0drVfU7M5/TwuQymkkfn55
WoOr2I/hn0mM35XFKQ1chipCd6zZRyx6S7ILbxxFG0ECXfMBCBcnADxtDlRWqLwv0uuQDtp4d3cs
/GnDtFhlS2jxTkBTuhPQmzuXyb1Cz8ROojErk5vV6yUR9kejiKLZClOfArDjXStFqx2fHPlp645A
cKQ+PXGb2+81W+uYcgCTp3zFh3PxoWhL7cSk7G+3L5jG8fgrpezmIAcWZ97m92iwN+N/PjiHtOl5
QMRK+bFMeBBhwDug4I/eJ/zq/zzUXsNIBm2CfYL758JmL+AtlWZE3xuZt7EN9n52+pM9HEgOn1oj
yrn7pOUmjhOzGjvSQYFkaXdhtOhX0/gOkIDL4NGuIH44m2F0ej58iEIRugQzeJ9QF5KnJZ26EPIx
/yefxJSN2bYlSWviXSnnKp3Dj0v8PoKquiAwb5fyCcJNSyZgLI1H0WcD5ubQtETZzQqyiBBIxMZQ
AjR8CCpKp7gN5hxQLzPAnBKhIomyHt78jddlmFjMDr5bpLXL6U02uKkWo5u/KDueGqU5QEL70C7+
x1EYasCpQ73mX/sLRy8q093yZ53m1zvFBEoy3T1HxBFQdsLR0Appl/HUj5fF9A/ELc6yFs/HVvQ7
xnh1j4auUdS8l6AZ+7w5pB+EUxjfPLj+YO1X70gcJ/v2CuAg7Xz4/2SBsDhDXmZEHjXmWGtEflzM
SUDIlshUCNIWt/CF+D3JK06i3DP26zmovoFQJleMuL+JAiTpNVgjhN1jEI22hGJyWIb2Nq3CKA1u
HAnbbWbxX6/x8gh8e+qQLba2S5UogGOWQ2XVHeFHhK+Tb0/G5pc+5ridrVpSosZZpwld6iwSkgLB
ocH/brQ85SFsRq7BlPuXpxJMpe8S8yic2OoLbeFAU6FTcqUg0YzfIf3TerbvpIT+VuckZAqo85Vq
ZBwJYS2cClQOZwrA1V1vnNWUnWNcPQykQY990iiz5gxA36tx+/U6RQYcwACzU+inMmut9Dj16c44
zhH6qTAmo/ld1M/9TItkcrhT42Ls5AVF1uKgcQPga3xlJpAC/mfhkq2K3mQb6JGtsib6SkoTDluw
EqvW9ulIyIyHsrTAc6Q5YPThEB5ak+1+5Qa74LvTOJM0DtEyQeUTSNnMQkZAXwjdw6j/QwIg+G94
oA+6WVapo1wN5TyoGAC4couXidz9sEdiy1nABwtyzpRvvuNqR0+vL/yFHF9QMCvRwW2jotIwLgib
e96KBy9n+rqtr4cKnQA3fsk9UpRfJGd5WspjTVWZbRYANsQ/g6Jg9l/+Ir8ArE3CUGHCZ/yP+Uly
PSAAwucoLIWTmhh/DExLYlf3mIRhNWYcYURUKjQ/diiZUvde53hSGUYGLuZtgOV8cZbutAg+Sxt0
t/gZsid0HqmHSJX9MdLwAqVaLgQ6sDUmMH0uvEdtCsNzRLUgktQyzb9DuUUs7cEbyqKkfR2FWSYE
XRCA7yRbLjJcZu1szxOS33bvxwy7ncyzv6EcyaxEwdtwo/jQmK55LAv3VXur4v6/U/MVBJ9deBEy
6KeG2L/CVrWVBVAH1bm5rrN8ZitplPhTcq3YQbeEe1OCptxjSi1coA72iJdh5lVzOl8Ex+NDbqo5
dAiyYysnydZIMf7xjDllf5OtJA/kMsGzNFvAqnpB92lJuv6w+gWdoAax4ex4swbTraQyFC16w+ra
jTMO8EPjhqUxRUJRsv3Me7MmHvvNv2CmOlINBQo5aF1rBU2jA8J/ya+1Kc4XeAJ0fWZoo1+LI8vD
5QVmJFMMyUglUI9AH1OAOm0DqgObYZjCXVb/WeftvBB4jjNjoo90EJz4P7aVLT6awCPKu2OwHHCu
B409/5vx+mf55WUOYAEKyQhDicAyZ1aZ9Z7tVs8L4A8tC1ul2fwY7D9Zartc4Wg9G3/siAOOVdVT
Ufc/tLsxwfh0OZsZfS0TrAG3/mFZtr/UN5qddfaqGZHqCPhSSfafXrZgW8m0+tmnXakZwb9nHhnd
5uW+D1SUfUUlrv8wj58YDqdnRTEY28E2zNLKc2KmEm05OknK+O87ng5VerX6/RAlalzsYg+9Lffd
Q71sFOlHSbk438d243VAcnmoGVFAknfx6brPhIz9bWC+lqjZVhGoDybpbhcihQz0NUzPDveaNSFc
osgAAnmK8TDMEbts4MOMZvvVehWkCHhoxFCrk4K+o/1zY+tYZzQoBnndbSW0ih+7Tcz+JibLH757
V/WVhXEb2B2Qyaxav55yU3okKyZZuvqfT+Pny9AniVO71wrMSxCTHUa6jvyiQRpqeHA4BOMAQY6Y
L1inRbT9PRXwdl7w2xPDdEx2tXOvIrRl4D/kzX06tfpzsJcRvqTvudqKnOO11o/ukn1WNgNEWpHS
zUh3KhMfOC4122oVGk+e8ItCNaWs5mz1jwOUqRBGSQLj+PXsP2pEFbJXsuSf+3vltiRgCJOy1suC
CP6RTxGE4+3dXlrsMUSRCGobXKEE3FpGh77AqM0JQiz7IPTex5hx66RfebFfeUxU1K6vM30fPMc1
nPfFOOwnzb+F+2NeQiSQ9MI223kudPoRGIrPTY7DI6+UNlqNCXBXp+gLgaUHa/nRmRD0195iwYQx
wBXF6vKqRZK3NryrH5KTGqSHowsK4KTOx5jE1dkAqySPagfxxMZaSu2DFAPdaHJY4RMGgMr6XT88
usB1QSk7imVwhTUXpgmLkVcyYQkLESjNkdJ220Ji/mPpBxx6UQkZHH8GkojX19OIqsVFi3I49byk
L64WwjeM145xl94AANXhXbnK02zBQrEh5uDw1iSgb333Kc7LLggEiONeciwzWJb7++fzOHAuhPzH
RCS0BTMO1IJYAnBTqj0HAlOYY6X1+dyyB+r6+0QdbZuE2mTGJgowJ5PCKwIy6UuFjusmuLtuXtHB
ch1oT/4zagnIa/b44Ty48Sv7F8C1ntEV+5iHHRb46+qUkSCMUidSB+vUj00Rj2xzfBcvWw5sj/C+
AYV8IVRCcse7tauwS39XOrVAdqWai87msOGgLSjrn37q/D1HjPMZnSHXu/wr86fEYh5fT78fv/JG
FJQ6BzJsGM8vfbvv9sUrKp8i0DHZWYInatV2pNBViVM58ZH32rtgGp2RS04Wkb57HTx8bniY6DkN
M6ZCyZDP39F+4dUkRUVvBjMJI+ADWmWRWIobViIP+7wdkh54ul4QAZHPXmn0tWmKVRJ1RIoxjnsB
CBPOiwNnG4Ixno9nPZqRmEXOIr9Rz91LO/UDghEroOTZfPUN99fb6FaYjJjv9vG+jMnrtnM3ZOTz
uDV2Q2bNxc4p7buWa1wHM7j2nthzNX4aaaRbi9334WhQxeeiw6KmIZ8j2GdSWjknH5kdQa4qGZXJ
q1FEqZaJR3BUb67xiiMZpsTgMU0+zw3Heg7J2UVIPlVO+fUo5HvnBDUecV/rrY6yRpwxRDusaw+j
Pha6hw5RMZHOCdDpR4Ou7ZwDdvnF9rc3UMlo3xp23uEEWS6DRCRZqxd8nxz9mMpUfOolGYIpjrEj
kDVD2yMROPc2Zu1Q3A0lmdvYHFezCh5r3JUfTbQlVnavIqKhIiJKYq/hr7r8stPLtuD+1MVXixJb
L61NLQj1oPYfyRbxuR2isvtQKWwtI/ENM7e07PV3KLSqQ07hd7r2cEsAv4lGAmlo+B/hP8xAwpjH
c1A0whGxvTa5LaFHxmvJf589bxll8/eYicJPd/ovsJyremHiM7e6v0u5xXry9Tjj/U02U9vsFbWP
aLJTiSN/HalKuLiQmXwxNhOhDaZZ7lopfH+hkA8mUl0ajhk3cMuvca8xqKSocNM6KU2h/lWV0a5j
DMMoyIP0rCNKxRmZ9uA3Ns4XfPzas30CEwxxwnPWUsKgbFOU9MJGqtqpEGZuIOvgQfiCgg5RN+Xt
/6xyI11NdL1oITSPSyv8wnH/Rje6DhU05hpmUvjCc4guSsd5ZO8C3EW/3iXXM0ubvGouIL8E2sDd
zbSdvFIPFYI5BD1WyWCs6mYsLxUaY+PYygR870QfXsO95kT1cog9NvRKKbASyYnAvcsm3hMKo2A6
oY5mZsE5b0oHuvkFMXyH6GkDASlwgRwUhNksC+wUeApciLd0IB2FY3WHShy0BIKb4++ks0kwyVpG
0sOrBaD0l2jFa2fa6IbrMIDX+nhPm+a2qR5SFU0SNeXGv4VlMYhHnvfIxalthZqJdftw1YUfnq3P
XM9ZLVJd0Zw14mAZfHv/7VgDW+LikwFwl+pCau9FPnslh5/F5+Kfw4QzBbqUpgCHPAcnpDHxcNLt
4wjq1YZXG30RAlhhOmIF0opd+Y6osoi/2O6t85RuHE/UidSFBH4XfIIXQLu/ugatqkLhettpZLby
IYjkYCHMsaQT7XesFU3rNacHGim7tmGlChbELFmh+KyA13idNYFof5MLMenDeXBQCB3pZ0q8OJ+H
YOm03WBf2V2xH6xGVpCP45P86DrkiWesNkqb003t+dxutkPHUeOglZXl+JbIdLB/jkZxpb4nWk6T
OwA/xZo5dnZdTOQauxsnIRQpmvIg461pj4YIa1qHfHNv05yYjgX6Zlu5if07Y100VF0hRqUwpKED
13xq7NBe+8wMc+HGtGj4QGQ2wXYs0ORsU5dNohFh3RBpsVxnbS46tsjd8dFXcorjGj+2Xgah6hkM
LnLMKj1iHoMHrNEBpGW8kVhN0UqxlFpWcoIkH/WW+8erNn22/pRDDee1cNrk3veAtMMuBXfSYP0P
xl2Bix7QGKgm0BNB8Eb8bQY/qd+XL8iwswjyKNaZpEojzO7xhS85IQQ5Bykw2duG4OsWgsczc0Vh
YSHGEQ9ky6fYOXQcijaxJVnulcebYaA5Ozr+ZUDbIao96KnpgP1Z/nx1oVSFoRjE9UcJUJRW7yYh
bm1+mNMBXkmBb7gssBojWpotrm+yWdbFxpk7VtKAQ+I8Vary7HQwFf262rYtYIQQ2i5muTawL9+O
+pHLw7hX1sPN2LPP2ZR1rlJVqahvE1AaBh/Dk5BnXsp4yr31dvotaUIOTRgzf7Oy/TcD8GsySp42
+C2WBooLsSr6a3fzNAhBmSUWOYGv5YEne8ad4haNbEcu4n0UrCyvwqipq2M+DQ5oDtpZE0zTJEj6
c2r9DDKuLySaoz9vjyAO/j5Pfa26M7XJjzDdUhJdXMhkMW5H4IKfjgGmdIOCknHgK36RBUluFbuQ
ceOtTx4zhk1zD0CbYEY6m+cWmntcQ37Buj7EUfe4POYdqas4ukbMVaUT+HHvrB5FeqXNgWWPvsmQ
ZxpWr6hM4dSyJFUzacGVywT1j0VRwLex4jVpZN4UeZTwrMuh4KTCi0R+WUavanZVY3N7joxWYfpU
9+eOTmHtxe1AFQGlBUUqeFhxXG0yh1coIpvCaoQEv5dCkN0cCARiHKDelZLd1XoIuFgyTJp4PoB8
qcQ+jNJqWHEE193cQDnkk0MwFYmb0Cca3zYevKKUeKAFL4pJAg/OngbCMVmLFmpOJ7cLcJUqzASO
94H9GNJi/UeBzPuXJDypTF/ITCDKA8zC2FXG/M3UHI+8W48KY+bMuPCKw+69TgmDz9Ia9KU3dK1F
jTP0Ul4+GqZ4tWjx4ORKWojDd3rXByuXC5s+QJGYtBo8bp4hM4Rud6l9tChwT5OnIYE6YjgDRXTc
YS9dz8BrYRpnkZxPXGNuphkgZApLq5Ov6GY8MFkXlujrsbn0iwU6fI+SvvBTO6hi/2d0k1xfdmVr
38s0WZhnZLsyAGKZXDsUVG5CKaUVstNZe1VZvP2T0odfx+EHyT5FUd1cRuyLPEh4Q4i9IuNVkwOJ
jw8Sg0ZoiIGpceR48MLA4OZzvcYUUVZV7pfvF40xE0NY6gzs/668dsmmhQSL4a82Qw37ns9ZYrqS
fMaXO/mm2gFzng8/eJ9gd9bLiLvIlT2PxNZIOSOn8XEZsTdOZF6tjkr3kRrRbdZ69HucAoyrryZE
Qfzf6racHWOLC1ICm00DbRJGUti+hUCL9jHEvvR8NAObXf6ycVu5M++911hjJMAJAGEKx8HHf+QY
Gzpg744BN90phjmdG9bDsM236BfqB0k+PSbJHSdR0g5Mi2Vh7HlZoFYUVm2LmWrzQPqS5NK1XTWm
9lG247oYy2tS4U9HtHs0yqaJtfKenWtTRuF+lNxIXu6TnGj2NvvCQAyjCX3EAlVwqXFeSgCt8NiD
eqGiW+0ME7MfkUoYWRyLLrYuE/NulssAITB1CeGRC5FxVQ9sziWdN8dIcPqSLQot5HXYetUmUqU4
+m41mCFP0yQYZoFPWaN1lrRwjzWFlNbpaF8opy0q+N0I01XLd5HRzAMmramtbu3zPJkeA6kuXxKn
7KbCIIKLvq2/d/jJxTmLwh+aIKXsC9F2DNzqIR596zaz8BVdyV6Hosnw8BLX4+VOvfHSiB6grN5B
nrqO/OSTK2W+bNBjNVPAbSA9zU/wLHNC8mdPJdU4ej5E0ovlHeX3unC350FoAv2hNITzeOhAhMgm
ERXF3/HPrvL395loaU/g8zC0tzWm0Ictj/UuVwjdJ7OY6V8IJ/DfQWcQ0TWrbR7z6yZ411HVCLi1
sDOAcMht8Gpv88urSg6VoJ3Sl02X011b4BEafxQe/glHYjskbom2r+JNy9Kkv+e0dJBRpfyNIsqF
rRaEWAJG0r4+Dz3YFVE195/YWLvqHYsz9pb0J2rxlB3oOPPt/pI9YQbWfAsdVhq8OiPrjHMKzi+a
WgW1W4CXIk2OtWzCXcqlDotn7ab6ru1tuO3wdv9WnSDYdvN9QIF9RSBcWPyJR+0YZIlMgRMQxayp
QSFZ/hvIbBtITCiPo3KjsCWaW3h4Bq5OtmVXlHeib9lWn7Ksp5j2HxYdyvTsykjIa1NAB93lyI8p
5BtkpcCNBSgIDVcNVhwCCpz2aRjU4TRe7f05FZNMci4WfyH0y/pe4Q8qMEGR04gXnCfSlGz5x/Md
tF4h3d8bV1oyaUSnKW7Wv1oaJQrGoVwiRjezexNV+D0fjUFqJ/6iL/Ll9613P6WqhytfCWN/7YIK
dfgq5jzTKeHnKe8MQRjaz+tNCXDoSJu4YMo77uj3jCvh+H+rEVX+dsqFSY+wedfGsXft1nXYAPcl
0ldwLSUWVJ//TEUTG53sIcaNZofnOhudIULhHLAjdURlRcxJszIFEPAF6GmVonVEIx9T2ytlYlaX
r54RK5mEKVXWmk5wmPkIxcmc/ZHGNhyrlF8OcoH9KdCvsE/it6UGdAQ4bftQz9zTViOtGX4JdFXG
tMlrVEelBpyNEFDXjnztP2asmS+AS4JhEKPRN4SyFV0m5y9hIlJFawTo8UlL7zp3xEKURoynsPrf
t6t74CU4zntuuL3x75Zerg+j0A2awN+8c8z9MLl/8Dhh8lCSngSnWOgnNGl4KCqrxzzQpir5NOM1
UEnGSbBWjy7x7Cxn5JbFMldIEMdroRLseqooo9kIkNex2ZRKIVcY7RU86eNWehqzJKue8TBAQLbF
BDrJhMlxg9W9gE4j6pwW5IWDgIghc8JtLvBDTy2dZOQQ+wptDkiWmH22HJUDv6ogRlC7Y3YhtWst
hJN3L2jcAhA646dfO4j0fybjXMXQXVYur2Q/PlNTtBmBr/+O66VEnADBpvUSL8icoLYYVZb2gxM9
WJGRky0zPIaNHhxvupchmFhY2WCk5bSSvNipBhz0rVRVqhz84KYh2/9yNM+4uOMqrZPk7/esSEtJ
cMDf3O8CH9tDTdZRd39oU0tGHCHSmkWuxiRCs9RfozqNkv6coJ9GeIfUwF0seOZLnRBKClJ9XAZc
t8o/LRsSN8BaU+bXzFo2ysevln4GNEohiXVuS4WrTRnD6xVPAx/uhfq3k9l8qWugkjN5RaEn2Tqo
e7vt5rA7v+IPVdyxvSrIXZQ/1j1uQtNP5BrvzS66W0Z2ziASgl5uFIjN9AGfNn8UNtgs2Iud9+ZG
fdCORiU+m79W5NdDPyGRjYmx/jEHBIIIgq3Cf7ck68qrhyllNHLMbprKFEJkEYIV0y5os4YD70qR
qiPeLH2ErFgtxtwoqUQkJqpVi+oP+DPGr0yEIfs2/EBNm3cqbRJ7UeKPWQM4/ZF0H94O7FkoDvYO
8B0A2sHvZ4ZN5X85G++55tIFJu6SGkp4RYXo5qBtPVeBWUUzM9Va3Nraq9L9ZPcSZh0wkFhkSJhT
sZCC4VsuhtBnJb/phNtFGeu52bYPD1iSU+rWtdil5f2R3WnZ4qO9k4LZxsS6YMTR++fbwd5z1R/k
68EmWoQAXot9/kWVeyp0fX9JO0gzMmDb2VDUtP7oONVlhAMLVucR7JQO45x+Jx1SHfnSOjOvm+BI
vj+fU6nuYBqoXDIBTFWt6qcCs7LKjZMaNW7S9S74n9IfWy25q9e6PAkFE66Lxfe2RUUQiGcn15Mo
9h10S8leOwt6YB1n6lZip3IVek9zEvALRh2PY4cseroxxNMEueTRdRxaFYpg5q/bwzsIBcfMiEpT
i6j7HBFol7GkDevzU0P9+T8lIP/ihVjWW0h1n12ZDmycSdtevrjaGpVs6yOsZiH2tirbWS2hODnP
S/VJeQpMc4a8ZfFP4P2p2FH/+HY12fQ7Pe1lBAI0tOtG5a4/TzMGGRtujngjCVFR7pFDns7kAZfO
hGR+e66PIRifRuZqtCn3qWeBNOdIFaT26UGd6WU0sOSyN/3XaN7drWkm2BLTtZXSe8/3dcXUF9Ym
T0zEv+1c+h2tUi2XNXPjzPYtcuUY+bRj2BWodWyZxZFKdZ0mdpk+QQo1I2huzYt6Z6CuPI41Go58
hfwwcY6hl3rNNHVzdo+o6EBMZkG7Sf9ULugxNF/msCcIhn9ItToHqM906sZxrl/eT01ozF2N9USh
E69zMsCox6K50gUlKn04m4pGMunvs8I7Mic2Ur3vtUH1pWJWJ5/o/n3of9sxdRWJWp6ruJMtACIy
TcXjnR4OJK6CVqAfPRpPR43qciCoxDO93lhJQnUxO0036kKoWo0ueMI6aWfgCrrwjzjmHcZ6bqz6
SJO7qqQ+C1ZPvacGYEd8DUrtnqMYbp4idaSckXoSpuRlP0+UTQkuzx7KJ1F07y810AGJgjPs6riG
VI7L5CV2XgY+7V5EwZhp8tTTeCpAg1r9MOTdZIuLXDFoHOny4wKAltMGWkcP/iH5IjVoh30ftmBX
483SigJ+lmp2taCCXNzfAB/kTBWrJZ+04eWwgfij1937pAE9AA6Lq4A3KdR9pBf9eXyfG66nz7KM
Cabv4trIelgCjT+B2r4D8SFMfakfb2Z1YMFXCJ88+5oWWrEHb888BmL++8Pbbuv9anPSV9/SRTxP
2rdu6OIE9bOeZWqD7L7bRZPxzdmfeyhL5LyZ1zu9i2RiTomlyH+yvFiFVwWE8IGeXdX1mJka1I9h
w+TD0YSA9xwGJ0FyJ5ZZqAqmGm8zd52ILChhv+oHjHrp9R42t126sXupwpW3yWHwt58Me1juw2jq
JmL5aS6mCpncD8g6bQwQv2YO90vXImRvaBj+iAMpaDhHcmkkqcsxyaXKFOcCGbv3QDgdENdFRcl0
aySd4O8uR5DDe8yL7WlQt/F0drl1qtl08DoMcjfgom5cX2MesoIdKmUUVxAi0xpLz0zLiIr3otYM
svQq1HwIQp67ERN2ffKUwWvmxidbIqirQNr1th3P0SojNxfdSm8jaauu9RUDa2WN40lPm9/rVwCw
0LfluGAnDjGzB66vXfsHpN/bdL6xVM6e4gIDaPqdKn69q0YDkc+b8HNj7bVhTAyIJFp2z4KOtKTs
evOvts9+TFq5+RsIb4Mly6DtqRbIdO5zRlFSul/qJokFPyDe3vcAIYBsxdBT+1hiTuhR7siZwOVp
5ialAtiB4K9idbj8Rv/GspzFFO0fcv/mYAjnaHdF3O6QXPf8SS+HhVCDRscIHQfPlaM22IE8BdB9
QFdCUiQIuaUrY9tytQWhau7G2pCxUl8z2Tp8/tfemNuPNGfQd7R/GnoZyH61MFsqfxHu0C5vjigZ
eNEnC6KD+za8KNSnaI3BtXkMDR5CS+5L3BoWDeNcOikJ/JxxssECP6ho4PgVElmSGuPYMOiCjgX5
Qa2M7xut7xAz2LrZAKVDwmGSF6EenBmpBIQWNP1UcwpCAdnSvUqjkvpKQHIQYWHo0ezJz/Quwk2p
tqTWDDSnrYGLaNh6TkQxGhHD0eS0rPkCkbkuGZf2RwWHspfsBreUcLJQsSMLZUEwwYtIc40v9wbw
rKurxG9Gb7ZD9ROqCfgz8+eZGMeS9FaGh6jBMn4jTNzacyLvbZR/za6UGZJxine8rHvtHZqrRz/J
ooFx/zcmdCG1TESIXZQp7BhtA3MwKRr2lGIW0wtkRHrAPNcC+01kfp/kWJEL07BteOJ2oFt8qUV6
TYd5guJ4DW755BuxXiR8uLwokvLL69fSrAwNByMT6DI/aSS6XcUZHLV0PGi1aQHuq5rmngiVYiZe
8nnkOk3/mIyEvGnR3dxMuwK1FwPTDDt6recw7+ekhIXC0tfTzSDT5ZQLIHehLkjH/X1mdrUFvcvt
+G/ZEost7GXl8mcG23rQaAxJIsCaCtzobgdJtDQKGGdKm8bl+H4eT694c7rNKODqclGER4O35hTx
XhkYjpk25e9X8pMNJN5azT2O1KCHHxE2r0IyB8htMDaxUOVKhrqZnY19PDCxFvZJLR+QvSGuHzJa
SuOPs03Bxubak0gTqXraI92jFiFOTh0aB4Pv9S/e7Ble9bSh0oUDPyHYhydfnJwCGltq7XVzgOhl
9TpslnQAICpKTFfI1nODtlUJgECuurdgyLKMg8GKeWVc7DFKNXsbE/Q5af34SQIiMq9oQivQBF4l
PWkyTsgyrdX0Ixr6t8HAfcMNIukZ1OqpWCycFt66fHQt1mq+8aZEN5YbpPI0bgJIxPWt6z6LJell
kxB2WkEPojDaJrXeF4YOD5k2UpKk9pBM+HQqA7uIxxdj9HNeAtMEn/IiUs+Me/9t2cu8kDD3TIra
5fnN29nGDHXWFK2kWdYKLZDKGJeIzCacUkN2G9gylS57VCclZ9s8LsriOc91Xmxs9nointSFnbtO
SYwXSkcq2l8eq6/vPHp9z0zHPsgxFGKwm8DrwGtIgEsqnIjxselnef/8i61E0UPGuhE8z582nV6K
/7BqkC61i7WgZhL4c7shcISL1JH9fjpTb92EpWxVgwK6qcXHoxAJqYVLHAJvm3urwL/SHOzUN7sY
eFgKIi74Sfyqu0qsIuLFeJ2u1awFPvxaNfkhLuw5QPFVt0REL6kVbkGUXbnnLHAFj9HquI2zE0Ux
3juzfG4z6hOuuHxuN+dijV4HYJgaUg0n9JBUGQc0fqxFpr87tzvNDfvSub6MRflGrGghXPNwaUN5
81laJ4rvjbIWSElk2VEGh4v5Gq/up+ZIIfvYTkNYe70TVEf9nTLcPlYzyui0ou24AZHunjT83foi
Jlk6R8T7X1Z/BgFEaWvuu5vHN11gZXk8KqXLbh23MsVuxNVaBZktgNBRGn8SNCDE3q2kynyEhUxO
BtUYh1R5Gqi2jlLi5/27/Y5M6kHe4J8Xk3BkKdLmpOwr4kmtjyh/PEMmFRbdtdNAfMj1h6wy1DVk
gRabTFuMBc+K3LK4xKHylxsMlIMuOFmCWrGsi5p5cxJ3ykUexNS0LEJOuLhDMCIvRvAzMq+CvPdH
W0xpbN41HBwvMbjJ+sNaZ7CX9g4/6/F/NdjsjWD0Rn/hgJkeE1sF/kqOrZA2N1krOT9+G/MXPpbQ
vpiHQNS+LXGvaJtRqGvX65wg6kfcQyJ/J6eTeUBN/I7B7cLk/vKFY343vh2b//cR/yS9CltSaIsH
hM/fZMcgUQqnZrAuRHGxdwRCwXZfQjulebxEZY2p3UOyBjjpVbo7LAqE8SYnTHI/U83SHlL4fUmT
iFIF8squez6IO5/eDx3sXwTaBBZFFivt6jIs/XZDwE9Yb6/OJIpyirEjd1+kKFeQmJS/lS32j2e4
dCAjcIvH3SJrw8EpB+qX2SD81wVUUFFfKMpZTfVKUE7wD0DptLRGVEH43vF1ip2pTTdl1zt6yXB+
6GEEaSBMBJv1ISU90K29FWIXK1zMoqvQWLxYRNwZDT7XHniIirYvBu03/zJT18LYKbfvuZEzxMlm
toPiQ4r14/tj8BP0pNWFL5jMtNCXmKPySDfVuIgldgWfD+jLmPTP8KgRPheeiCqgJpjb/F3gdEDP
fCKuylSgi2jSKO1TIlKyOKIE+qjFcgo3qKcxksQJrLLnSNmY3BpyqbhkDGSpF18zK77uoDCexKXy
CccLLm+7OCBAiUifz9vWyghHYiiwCQwB4jvWVjTHni7Cs0wqAqTr6DEco7Jz5m2cjvfxB09LbtjO
Q55HyBWcFD+bXveGcXSzaUsKG+6O62vQRjtwHUvjLuypueDBOSTt0+mhLBWvfF4cx4dxiAcR0Ae5
IpFAvyZo1KVAByrJF+BDsZOHGqkAveoFCKwBNmqGZSoYxTRK2EbitCircwZFabPdSgzLZ3ktqmKJ
lMvKNfuhfmrBs14cvSkHbx8MaXMnDX3JLW+UtdfaoNsHETWbZgNax2k7gSvNQQx5geBSKJNTn9+F
TQRtLIa4LiM0guFClZDYwvB7d01bBWUc/wpC7aclz0T1OxuLHrI+5in80holeRJiYA3y+++oMeiK
AL4q6Ldz3bCXRjGy1CqJPR3ePnYQC5VPaRO+MPwepFRPxneAPEBp3kGVw0tmvzE5xL7C6C0sngjo
PwXrgJyU0N6JV96VmDaOWD1uMAK0MymJNkVSk+0dV2YXOiubgXO8/hnWBZTP/9qTp4eD/8ON31St
LWeTggFUMmWv5Dzq6YwX9DdTEFe5D9OWb6sOruq/fGDTwlAYZBHCW3rkACVAw4nTSQBU0podIZqx
Lqz4xrn3EicNTiwOW66yY5ajvz7pO9nqO2R0SWiMR+8kQ5Uq2QIRTNmm+4Af0zAWXRBuOt7Jc461
CB8gI/8eoG3uKQ59v7lKvy73o0xiqbzpzAcKQ83cuk2RxbOKoArsF74QSSNWYyjyWZ3TwHSMASm3
wvsDf3BoncZlOp8DZggul73CvUrQai2V567x0Z8jpRWuyT3htvpelnG/Y01EaWy8S4Ng3NwUYO6D
uTvPNTcYIeRPe7wKL82WWI+m+0KQZbmLxe4UQe/0dZRzU63NpQkRYw2OrmyAG7rkZCCx6LctWodN
JxxSf9WMeGmi9IGhc4Lv9Om7I66wsFeC9RXYbIstdNVyOawC6eiBABDeCR9iyjvm+Ahx9s6VCYLm
08HZ+sZwBEQE/IQ4+wG4ICv1ouUw5aoOdDnVJpoQCtub83vDvVTkJ+vlPRuLS4Qx6Ez62hOOJOZB
2wR7Tjn2X69TQ/4eeeyZaSoraGJocMF03RvsRN32D8746yaHYaTn221VR/ose4O2zFg/b3ptQ4/S
g2YGpqCgvNap8Z6WmMx5C8tG2pihY5XmNcHIkvyavuYHm+Jm70xYachycYSmhulbwvcAu79qEClQ
zXUN8hxr+YeuDH+KkRBJ/TS08GICYA1d4SQ/b7PUSq9Vpi4YrR0UjCojZpxgneBiluRR5XF3GbXq
gHhC6QSAhfn+RbjaQ09UUMCgnjBRdiOj0fs4okiwoR/MJOYDDXz1O9F56x2mQYdQPL1hExcT/+wS
ic0WAYM2NRkr4cOK9w+9mh+9Sr10/pscLSBEranhSaWvAHPnA22ba++9BOndjtPlYy6+65Hxi/PI
oQoXsu4wZkgBq1uV4rx1r/wqR5wHeas7r55eRrQdH3KveE0HX/q9TXUSX39qC24BN6ZrN8D1f0Ux
+41JtdA9Z1T5B3BnSALzAws9oNzODmoEhzhMLXcY07sToswCHFAJYPNNvNn4dTP1K5r6NRy0VQlV
JIXR9UbDBIK4rf7brPxdPusoMrYUGJL9BJQVMy3YrvNr+TpYAA13GA1JJp5TURqyFVfGcXM2KkUu
C0j8c/WRoiLdBUAAaL5J8hdiKWvh9ms+JG475mxDf/K53FYCxOet0qu8fIdlvTrOXTSesforqLKR
xb5RPjihtyqeWQOeqe+jvoHS7e/NY1Sy8xbNz+6/QumyfSptItHopTKYrFj4dsWV8sLJ0jCKaQOh
Q9tS0RpFYImkkKqPN/m5ZJM7FMyw2bf3JHtdU/9scDDAjROGGlOZ6zN5Uu+1wEAA8FQMCpw63pY9
r5dL2DnaWy3l+vdhUoJ9fgHZkoaZx4enYyFLI+pYrG8SzN4/PLVAAcRc4zZeIfOUbBCKkZcPqcpd
cCVojLNFWdiiD5DAteClrBZXlrIp0fNr2zQHPo32USQ7qv0qW3wPFKBY394gaEJH/neBpUjfubRh
w4tHStb7H3RhUY0YqZq2R8tpZFbLqGJPPZkZbjkybjNf8t0gHWtqz+u7DOmuwlcNC6syA5EBZ5AU
c4BCxag2Qs61Oy+RtTLxWe9AKiwhaMcJ6/b5yI1f+yvnEyvrdSPGTLwRanL8hUIpwwTzEVcwdDPB
kFxqUiCQuduvIxhQ48pQfAxBCO9hbahq/oMw1G7vw/+zK4acl3xh9je58Os9E/RwBNC8Ap8kew/T
mGs/DFxOTrX3afEXcz8dYcHg8vxcRf981ZzvUykOpMEs2+Qrd+/73NvR3J+QvT6724NIi+8UyclN
RJ+ysSN3O/c67IRSYiA4K8tS9z2QWyGEGTD4IK+2AW23H060hxFX837dBJdAYUDd9avXOI+dUM6Y
x2+X1lYbvHDdPLZOYDliaNkjKkpmWBdYWWMUKh7IZWpD6Mzbq4EUq2dOBHowHjlx+5B4TGV5Vuvn
ExBlP+pewp1POdbVJudBOgZdbOdgvbHCm+6sohMzHH68VMzUyKonxxJODHCGkMDbTiPkIAXSZZkM
mdDnX4PSl7GRycw3SeJpjHWVvNXVaRif3nIKeAqOUky4ZEINY1ASC1hKyhMfEtHGA15hV2qxLTcs
6gVQ5xcVi56v1TvXiY6b+/TsndiMJcUJL8eEQTxDxC4HGL9NuL5HVNb2YWkypRlBp+dh87SLBMvH
L9utXe+VMMKtw5Zp5hg8Ts5xfDotaPqQ9Em2cpaYaVC3CqXrJWHdf53k91YX+e0Pni7trid9ShGo
EFQpatJ3BOHtNBG05mOKlEm9ubEOI8yA6Pc8yhkTv6WU5C3n7kGrambAO/E/CBaq5zfVmwLzrvvG
c1shDj3uVwJLmXIW/lSEL08UjnR7PG1Y9bzY7aaX5Q1aoh++jPK9xI5gxSxFjjRcE6ZkrsqdaWi7
Denn+9Coh3vQx6PHnlHTgNrPT56PN+zJrrSmoaeaE/AjKlTwp8sVkngX4aZs3NE1kmLhVw33fTkZ
Z4ZZiwY92kT5LWM20QbKRLoLEGfvN2VKT4CrYwPnGdpVUPePAl9B+PtlzOc6GNIC0NJ+/65Bl0mp
8wCSrAqIZbjIk13ew8FRwHKwIGSg0yIsPnFYviohrhNww6UZBP6V0nM7sGA74R+t5OzS0FgS1XTt
vTy2T5Fb6vrMMXymB7BYeEbeOuwnh5OvQgL7TmMoN4ZqzvW6k/lSXqdaQO91iSjX48oMyfbfqDpv
tGCCWCI6SA+ewclhqfol1ADvXnyErEYWwYS+rQB+G6CuLrBdooaayU96jg3tD3jbkWeiQoWsxOey
vhIAmb1npRhxqN+JLSRR/blvqcSqvMOGqi5KkwgrhrMWMYaoG3ZsrGr2oEKzO23pHPdSWWuB3hSq
rKzTjzYJ9zoCZCjDyDzEgmtmbVvmOtyVXHOuKkaH8fBMbx9xpzrIXXdTsWBbdY2KMfaioBKl+pn0
loPj5CYeByn/4HflZwIMEZpK8iw9xM5FXhHluPXpEfrAIH7Uo6o3gKKLYn8kTBmLbiQUyyK9aqxR
n7cWhoc0QUEubeNF12jbUL1WAcs/3+y+HLf0o1iE/lOnYWrPv2rK69vobGbMf8ITVxl55WgYB48J
MRSJ09mKqUI5iOeDO1t9UhJB9Nxui5My3agLLq+15KCQIANVoZ+0OdVwmof6jt8SCvInkcCtOQX4
89FPGO33Etjz/D22MZ+pYg/Bo2Cgf2aFhWfchafMSpqme1okD8FLwHXLj9o8bATMhL5bzDrmq8g0
D1E2Zdz2D+jICz+nR2gd/cG5bE5jqdjW/1Y8bnFAezLUgVOa/lNkFwQj14hw1cHcycD7vKmwMSlU
Ut0wpPwV2uMRqG62OoPDHayy3fOaUtUVfpWSLt3llerofqRd/h2IYtVYmwIeY2U/xcZAtl1ifqrQ
I6jD3TBRBYKp+HF1Nm2FlkdjT89Kk5AXNeX9SiFANOURdySFruLowlCynjRtCzyMNbmMxS+Nck6t
BrEcvt0iioSTapnE+kW8bOBUcAPBpUIKn6XESZkqzGi/Khqu3TftcPvRxRp2Ko5f6gmWYaNW2ot5
O8tIAdj/SwglYw8f7vABKGvxCfxne3hRz8vu7s1siPJO5YDPXtbYrAA18SGFh5IkNGFegimxZ6+M
mcLATogQXvITSloh6GugGDGExOrlsadgJJwRjY1Idc+KfhBWjCCr9pdrcokpgiSY2pnxBuft1rH+
tBpD3O/7G/qUC6WhXDqSuP+M7VhAzs+A+BnhA6U1Tnf9i6udHUUh8rd9vjy0ZAELyUv7iUvQebtc
Fa1g9F1d8o3LiapZdv2BCqN4TBBk7zhSX3+TBwk24ZX0c1W4CfzxkTkokTwNdhdCP1+zJKdGaXaB
VVs6I8IR2wry7CaTBaMcdJu8zrL65xFB4cErihqVsYDN19xue2cvi140f8kLwUfIwfkBH6pG3Tu2
tQAebM5CcIMPyaXX7qK7B8RBYkzKP5dDgKrOMLGIHLdh4fuaofdG+9AJ+TRRMvahTh7MBOl2SQoc
G59SQquEnhtMIUaj0os7wucafuq0JVM4un2FU42jSNmXxgNlGlpJfd4Rsv47Gvimmvxy9Wyl1DzI
kve0WicedWAVArGt29Wg54MPswQR5uIXlLrDSRyAeGUopQEFeiLYou1Z+lacE861/zfD7MI2WxJu
diyqNz4EgNmNb/NoxVPIBf5HwShsrhoKRZ3BHK/C1gn4VK/Dm1/58jALn460vhY8B/e4qM12jwxc
s0lHpCCTkWaGwINb8T8nZbZTMfD1V3Q0d7hz8TMd860cXU8GCF7yIM0IEgS2kV2hAAH+TtmfpA5x
13oP8Sm/FdeL+/0jvqTlCaIEODG3++1w2IjbzhDhp1FCjePVpFUzL4Ei1fQslD33F7z7YMUD/xqW
nXlktLhN4Bic+bbvwbUzMaJb9Ukuob0V6MDARIdDuLSS9afpVtYkTngLr9TTLwBn5TVYZvTYjw8Z
5a9o8ubTPU9KJIQn/uycj3w66OHnXeZlUh1tnVmbjPWJs4+Nygoyan2cD7v+DxueCIo8pzutms38
a4s07C9noAk9AiivJl1WVcTb39w0ZXWZNROF+F1QcVWuThS3okgdKmY1fZjAy5XomNQ2XBoUen8B
fqOlCDyyVN8MDXvYUSyDYS2p80Fvn13xdf2xDsEbX6CwS/uHZO1dhknnKlB5U8+3+34LA9O71cyw
ayFXRizk+I+iXh5/5WXr924SrrJ4uH6Avjlc2tx9D6sVBjL9WaTJhOGlG6+NlHVn0g6JOo8IVzhd
i7Rc3UxTQaNnEdBNrfo8W0gu1D2y6oezLlgzo8lOMnVDCtMkO3fYqLuuKhUeskaeN0vGSo1/5zwl
fx87wyW33R/KXU1sa5NAAqrSdyPeKSCOuDpDmfVRiOT7mRY/uNyBZB7wt068kbtRfqA+1KVkfBSI
DpiBcWm1k/7JcMDUqVnjiiZAcLEkTuL4DOxGRHSjjz7rBfpzW1Ncv+oRBFj3xKRU7PcD/3GOaVln
dgFnIonuuwgaZ345BncMPXtqKdzsX/n8ZXTuRAdE1Vn6TDo7KBGhDNlqjzFw6QCcDWwVp+mdDmJ3
ZdKMYMXsPpuudx9rvRt7dGiFRq8j0Q==
`protect end_protected
