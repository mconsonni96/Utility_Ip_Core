`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
l6LC89LodMbN8GrVkHB0+2o+Lf4Dit1XpdSa95ooiEre/6W42/BIjtKsW4DHyGyckMZuUvRcnNv1
RLICvkVzhAwlIDMmjLG6DM3g1AOVEYte3Sd7r/+ohxA6Fogqetc9e55DUPNFJzoKJxHTk7/03KmX
12W1SGJiHxCdiBf8Ou8HMIaIg7n2/0KtuY9FLOS6q5/9CY0uydIbDV7pJiQcTSI30dE52rznR1/+
CsWrlGve+Fn3ME/9E6yRYvsvi/bLvmDEbxxOhJFJINr3b8/C9jAsBxMZgKfGNjAehoJimfvGRiOo
09R3DZ2qFkwjSggZQQOBZAh8x2XCPQ3kEBjAeg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="nT6Phv4mq8aFx/I7d6VyCpQSgyZtH592JDrTI7j5bKQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8592)
`protect data_block
JZdMUlnzyt+pKFKA8/Ov7rGHwMbPDozzdh7u0w6D5Hjg1rStByMrRsScWofb1ccvT+8S3SgmxhoG
3xTTPPdRouX39GHYp0zyFcBTzxApKTgpNnKhjCAUbEAHYwS8AAzyZl7FkEylU5BtAxr8PWvpqvX9
W8VH/ePwQ2zq6kcav6Y3xSUWTnWYd+fwjGqmlwPRWsxaO58Cw5LiLkLhNYIj70+g1BJ8Gpt5pdQc
W4qMfyVLD1FMovJ9NxmFVEMe9H4evDDRyJCZuZ4rbdUxJoKwRJN2EkoI9hUwIxdpC70sUQH9OdvD
PpBeSsqchgK4FG6RTUPc6+CgVUyZqC+sjwKuRxFLXt9TwPjGC3hRtdzoIdMpSvxFQvKvSUjS4WZr
h+kccY4sm//wouRtPzc5373lzzE8SSXlhSoyHPOXUUsF0ibSmq/1uYs3XVLsa0LEGXn47u4CZ74x
dUjD0vN363iqMPdCDaHGjdVTpobPLeS0sWsUTg/QEB3uRRWVcK3QeP701tTZNVdj++rmgQeE/Cqk
DPogrGgQ5KvUhmmA9v7qO7iPp6QLog7euVsbeE2tj4CB2Hx+Vk7Gfm3TrA00kYR1jAbNRkTxs0QX
T5A2cf0jYMNP7LotZvS+anSqAOm0T4KE7Tl9caeZXDtpIFXVdCO91kZgHyyFcjSU7RISkRPIupa6
g5Xs0RyT/dMfisjybBIVKsiic2ZAI8WmGqKI0HzN9QOH4/Lgo5+v7CKLdIK8nHm6/KVi1wx/RPfa
K/TFuayEZ4qpE/3pk54KlmpIg+/ngc9Bvre899Ubhmhnt42pHtylqC7DZfxtfBNE8MEb20SOgPcL
v+LCvBwlmDAuGomZBK9U0sY0FsPwRoQB3/qPpoh5HexsnUkprQlRRlqKZo9GjaMxq3Q0rjJ6BkaQ
F3huCd/UnKN2D36Dtwjgs/q8dxLLpoyPssC7zlK/H8pCBw7NRh6dn65ZhrNfEXDcWW5tnuEOyCH9
shn9iEKICzw88ML7PVk9905BHoSPfSrro2JmJJ0/Hbhnda9FcmYirpG3u1geAY48+id8ACLBN7PH
qBnARB4kWma4EXsAAvjE6L5IVeFwtvea6So9+lpuey4wFy1WfViO9mMcT0iqB8B7NCTQTgS/ZTUj
kgXMV4/6rnH4IryhuorxXexLD7EXYEz5OFJh6e7tadyzxnOvKv+WyCLeclOK151Z6E4FjqaBh1Ba
5N57pE445XT9nuVGWVFpN3ccdUT7UkXD+IjLhWBjubF9fZ8DJgyHj76fCgrVot1lNzmS6hM8p86U
uIF8bvZbGqpqqXLl6Llp/29nMq7Lt+X2Er32Jra7H66o0g2uLPT706KbRV8hRJkqYmqXNb6csEY7
kxVRBAGLPBinr6LHBbrjLXQ9t9CAQVIzNhLBhOttlOGF+49p2+tuebkLhHq/JFAtUG5eQx4B6S08
unnUixjjIOGzQTP2eMiWbaO3P/2WdGiPwSbI7gUTw2WRtMOjxDZs84/+QsLjJpK1verBbvbCoYRr
JnN8SKkyl/LzDbB895NMoJ9mNyUW1yBhSvwl4GEH1ZlSYe3vthdijMy0K+V8TwPVRUbjqoFDSZHL
YXAT6cFhlxephKbgKMlpzpwEeZAk9r1N0JMeNkNiyr54iwTC9g9G+xg2+WkMFfdUw9Ueo1Rd7Jz5
OjlYlCNSq6jLiu8nGQvr4DGj9VovhkF9bv/+VhHJ7UO9R7ldK471gxNfTSej2sQIhVIzULA+kVFq
TmUy566MOXC9xowiCB7Rhb6bZIG77hph1Oltbh3MUiutXE+ynGh0CTsLpYA5SeSwiF3DaLG7TnL+
Ejr1rwXfISWMbC1whO/dKcn7EMBC1AI3ZcdWkCTksz7C5GQTNUrn3u2EZgk7+ib79rrt3PnrARPQ
1uxx2WJLPC8nH7nlj/O6nXMDC+wgs2g1th00C24ijhKqM8+q0jDj0htAo21TDlOaWh1m83d1pWXP
2Z0o6z1qmiFp+E5Q9s6JuZ1i38DiT832syBjzmgqyUdyRteg2zOQMPQy2ipmoGIPalZKuYTaDHh2
+iWajs/nf6a8oYnK860gJcrmg9uOzfAuFK1MP6jZTWywOLlfUwiAMss0xIgqfAO+SBc4f27eDRKJ
baFomcVKEuwvJlzRReZUKfKewy7cxuX0GKLQcjr+OAx1pCByXlyqjktlIV0ACgdlIxgIRvbDCWzH
lsRiXs9+evkZUjEfz2swMDZIpP1gDEKn52r9hcAva8ndwz9DAxJ5yCGafKJeFzknZBTV/u3bPtWc
vssZ0nIHiZ8aKiZAXo3tgql8AvjoFZJXR5LucJtRQNqEYGP+EFJVFmcdK9++AfhRb58XyNU5tEt3
ujoXSHHVRj79/Sm2f62Gmw6hFKrBedSblu2o6+iBBlnM7DTlWI2WHMDz/jcsXgvi33Ke7sN4HkOk
BTk0cbopIvazORKkBF9Gb/AfzhCwKVgGmber+eAx3CYJeHzKemq04+0dSdhF5ySWMECE33M/72ET
ajACBXWuIXc0FeAw31g83oLdtfz2RABJaJwiQYkQt4yBMbPI3nHi58qt0T+Cxab0mcpGDrN6WfFg
gDzeINJssYS1LUdJvzAIbM8WdbTwx6Ll0w+tgNN67pv5Zu5VUrIncjb/D/3cGoUBLNaGCkrdA8XM
91VYLSzrga76yZqriQQwBt29OkSzpEL21B2hVpOE++oGaDH47bIJIxIVbDyw6FFDlwnT3uaOVcNp
dbK0yNL+X2NqLz6eDtbHo7/JjkRbg9R8tzR9xqGWmhpyH63Dva61WEAnANr6IZuSOgjUq8Ajvw9E
fQLf05wxO38uX7bqV+iOBiyNNk+lG0F1pvOYBlN4gDOW8jlo3WxIQiW7APnhF033qUj+5u3chL9b
hMPUGhCeHIBka3uqDAOQJVOp8L5L97OuV6sED0Rbe3VqFwVxsCKRsapHK18OyM3XVh2Kmo6lJOhn
YhV3alV6iL/Y9BuaFCqO9gr1X0L2x+Codg/s3KHjCpk/plobzNdMFteuEeoPHlnSbWxNS1NOHwDx
fRyZbGhTSCCpoeHyAC0wno7UvwaQJ7tR9iNV4L0t/R2ZpoLWCB4OjHZrL/KK5Xm7nzupoJlISnRD
QdrTDGeQGw4CvmD6VhFnsQoyAmgDR/hlTXvAlU49JIfAWeg4pyS8J6zhi6TAcAvKkBiZ2a+LtWbd
mWyF+9av9G4DI+7WHMglfYdkT5qaL6MwcFLJxCztfRR4PmR4ZEclbYKaR4PCmBFdWNuxlEXN/hK8
Jdb5p/MzehvJALi8I+FmSHr1uS2J8+H0RdipzHaT5fZ86MrAw2Of6Y89MTueO+YyMptO8Ufme+A3
w4VTQkXkXQBoL16SLggn8yZ9c8ssmUvDkjRslnyUjsE4JQBtUAms2ipARD9GKk6dl30ojpTU+gnd
lj1eqR177ubJlUPN0e06yL9vSBM0pVXVuTZEweOm5F+RqcApZ490MDxqOHqoyivS4Gn9R8vUvs/T
NIFndABWXPqeyyH23y0RC909Ieyri2zKFhZAzGXkazRZ/ZyXaktY94+HS9zYxCoenfgLdCoWtciD
b4ggWuJv1Pi5b6m8MewagL3Bfi/rox1G9LKG6xOR46hAYh8eR05OzPkepV28sLe7x4FEVwu/QHex
OVgWUUEzZt89AqpBMY5ygOl8Y8zJAmk/OBiMfl08DOMSQo7uq1LgO1/ZiD6ps2WsXwq+54P4EuIK
APt/YW/x179+7/Bvf7o4jUosqjEhp57jx7j0MmBt6BtlOfX4RfxPh+HTTluQiqb64VpCnHAgJgXK
qpF9uVe6MKsYJvK7+s3herOamk1I8NJjlp1NJi26a7XQy9Elk6NTjlCVAZSRv8RJZJ0E4EjGG/tG
M/0kBL1y5RijC3++FrucdnIWIliS559ILcPR54LDka0hTfv1ip/kBgjUMbGpr1NQXdKznhztUdcw
Ilu6SjftYlS/pAv58RUyvvMWCX1O7JMZS5fqygCp6SvSzgdua+lhsfcjpwYAySaGaXmIOVflkqa3
OMR82Os46dxzyI2bm65e0tNNZtNj4aSq1WDNpoM4bCfpttyWnLJWY5p22vwtEfJLAwmiWPuprdPN
mibfRrRkYCHa3HiyLCY3A9+B2wYGsNMp/gkrfmSWpZlsJ/q9ggW/pPcDk061v9ld2XnGPi12OXZp
uutIIzlcOwBB2mTP97XovmLHzM17vVULUvusgOfEATbV4zUM/cJ/N286E717Ec/QQX5l5EXVdEuU
DrlkCZPPLsUGoq9rRrpPxQezvkdQbaSaMMPebv9iRMjfbARoSGNwGPiMabCerTibf52JnmQDQgyk
EzJ6/w+Z41YzDhMWb9naU02xhur2elacS7nvTEzXknaHk23tWbUQWb+U0w52tJ2u/bl411cbGmjt
ojBX1RxKy/cG/U2ruGMpVxI+T6jC6XWXMz6Tb/VhWErNDD25K5amcbA0sbaplbLkpaWafjAGi0zr
pHbAKnEO+rlGBP3G57GYf4pHpMWVVZjnl6noX2VqBV6XoXF5ET47KREH0rAOfUM7URWjoMUMlgDG
nORX1kkIfrJ4ugdFO90IhgKD6+3EfW1hxWfczRsFtUkWtAabSX5vbRh/OwQ521oTLEhSzyzYmqXX
Gf0Qr9sGZfCYazv1RnsM/XU2xJDJ/SCO7CQ06dSAPRnqXRez0wZ4l3ULl4/HzAaiupMpzi6p1+u8
PS3shX9AoLkkek4UwY9+PYb4QpmIzRBDwdBmERHXxofJBaH5n8mVOajflOgbPzNwMKo/lIuXGXgI
Ce50+NDC9GBdv6LTsc394bxWWF4WrMhMj+ItPzuYa/prJ9jI/rSowNqKm8KxeLvnTVOfh+VRYRvq
Lw45RTadac2yQgcaeaaGVKv6uv6DAGFq2+XQbBzmKaLtug7H4/qPgQa/a2bq5B0v83zgFtoU6l55
6HtrBAokd2cVv2rMtRc2GCwTiq7KfNL+oLredojEomutV/AH5ok9Tly8Gxe1CnV4BegA6Ph0tI/2
MGn1p4v2zO71opIDZsl/ffoGoyx4lKzeImC1k95TfTvAfZyhTEBhjppSp5FPusfQbg+wK/bDoct7
zAf53L9myDRO0tQZPNvI7iWnPpCbhS8BRrbdZXTvIojx/9xElk4zyi7TWS0cnzCt0qf9Nz0tchfi
Rgs6jzhu2hU/1Od+8/8tYOeY/Li/ZmUg0LoLbXaUBnpkbuKzOTWWL9hMjVP7aoO7xPoEImA449Lq
AXxXaIoFpqXywKfgEwI3MwbvubllDrsjPq08tAVgVjxwoZIGlpKuamNbIegkJWdsAPH6S7D0j2Jv
kXaXzqwSNuA5kshH+duVzbAKUm0AnYwlXioWAq5g9CAs6L7TkY0ftMI6HCX8MbfM3Wqml2JZw8MQ
huubotm2OBQxQWPOFBM6UCmfwDtC2PdUr3oL10y71OqKHH+1MiNpPY0QPWH8q8FaNcTGVgphB5Us
mpOYM0kscsHma+lOv/H72Qj045gyh0R9Y7xK9W/nd5LTlAOei97Tl2IP9R5HMQyQNkjo7loI382O
Qn4NmsLAfRFpQQeGFNYkzLha+rjjuYwLZSVUF/tQP4XyXYVNXQz565DJauuInjK7h7RtiybKz5bJ
Li81nPAB1yXPQ+YyZRUPaykNICwbdcJ7I+Qk0nOxoHeAyyTqLW3l2o8IosK46OczQr516GzpuAx6
CSreO+rdYpCzDt5VKAlkzKemosvGPsowFu/qGCaUP3aelS4Kp7ABITtqdxmiToVmMFg0/XlkxK2k
T6PLvh8OBYuCI/XytrYIwyPLHggY1Vd3fITw5TGiyVQFRmdVw4H1eXaerbt/FgHTp6AvWKnAFy/M
WF+SanQJa9F/TLP3UnWA4a3/MKxxW4aCT89uEX0lWLcvNpGGY+CHd01u338/PFlnwzUzWxwx8t/m
bsslYoSEQI+zmi/Flp8BsWxxidFZoWwLMlvovrEsF6rIXrdbeYPmOgndtAChiWvxmq2scVCQUU/q
XvoTDBDudBrCGw6OaWdDgCWiQx8SgUY2vB+XLOMI8nnmsMRlmBM62yt6LeWwU+0spSXDK9tfWwJk
6CJzNn/kw9ZY2UtgCaqbuIe4ds1FK4yrsPzTSKBJ0bp5xjRUk6syjzZrFIrLyiNuo4/AHNURUoOR
SzmhLg3d7dd5AZlVvB8mgncIUtrhBWymKuOto+doQgt1e3wiW8wSpaVv+m+ZQpeM29ZMtvt3daOv
fZeibw3/cQu6VL1N2DuxuiFNcAa2rNZWGID7I+aTFiTGO+SmnS9ThnY2nq9nFwDGJ+KY0ADOIbVp
jAygJqr6Lz9B/8dObA75rLjp2+jkLfrp0JRWBmq/KnorALKVodPlXI0mQ39xDWc+A0C2SPLzXATk
eMalXWQ+HlNqN/u6pGblhU1G7aKJLVs5CgGx4x532HArgDOA6Rm3Wy0GL1F+9xsidBiHw/dPKKmn
sRTZvc2VWzUTtdSuwndrcyyTfqX2ovIvELiiBklO5NPQlVf+JiPain6zMJrRgN45ugRoS+0ndHiB
7rUi0MKG3UGBhnbqfk/oowc6YF+7YhQHpxh4lJ2W5vSEFHhVznZSQ5QTcXFgEzrZFaK8NtaX6NS+
sfiP86fI+gkTi4hd2J3x9wdp1/iGVIMHWt1uKxoioT5wMcBC5fy4/G4JUVLTalzygXcGJrFXtLI1
xshs2AjCbBWkjvknYkSyfOLAngimbqqhg66NsZNEBhunNti8yn3xjtp+aKbNRT5p5cl2344ysZnX
cZSqt0kOj8C06dVPELAq+FOucP5ZxlV1vrk/o/PMYtCq6Y0iTiVKitmxIJxd0ssyOBEbF/yqg7Ja
j/5JtLenqNh1FVc0osVDAaP1TN6cIpNFCal0pVE0zxj/kSO1wntFOpOTszPAVjnikbE28v4uLMf4
9SZNNoz8B89LJhhlN4ee+bBwT9tQH+WPugLttSQyQkC8SCX7QoPbMtQJiVbZ2Uz8HNKRPYasGybj
rDDcqNhvPNlNizWarDQaoFtD5VImFWAL5aDzTYuXylj8IGwpUrAjea4c1DeUVYWwCgB5P2BlWYMG
5eEpRgi4iddLRl8vqMjrefzMO5JLMH2j6wu3cOETlQGaxM47kTD548am69xJJ7lErWJ6skE6Ne8O
1y8lD802AVVuuRWjIvg7nDdTIykDWq0n3n0lCEaOiCfqedBXFQFpobWZgqawgyJ8r1z456YJ0GqQ
EgcFTO/PWSbsmBrNlRmLQ9fHiB3UVmCku4TkswgnaR81YpS8o4tT5jmERTwegSIyhNm+LX9hu3Hv
uC3OafH4B0lA60on7Y/e8wuQTkBCR7kjWBaTNnurjC3agB2hB3tBVkcCbdw9/4jJg6fFVPFwGZaA
yIMsTyeLzg+nJrzrQsr+k7EpHrfe0cjeZXPhqLabY/sK1KoARH6sXjD5XBmTxl5O9udpK9AYo0ON
1Z+JTyzKlm6NpIkR9THYN2pssiEXkT7ZeTugaaFCGer6zZPNjTksBTUnXbaMUMWlWVJ2epf+Nro8
Qni0R3vEzy+WTfDqHOA7GJfcjkh/BuMEChFHq2Uy57nr7kLfIJG5AOTmgw8C9Zwa1y/BIBC2F8T5
7i7WXlXSyxKwm68ZdTshQONrFLhxr06d6jis9t6UsDE1qMDWPGzqt0U6yT+t69JuJMLciOdejBQ8
bg3xPPN1T09QmrTiQXLmmbSTToOefdMBUXdbEVYRsOQc0XF4gIhrckhPhieW/mOxQ+ftcmiThhTV
5PIr2lqnReUHQcEM31AqGj91LiNENqLoxaWBSD/4wyyNiwEyfTa0fyU+q7uOCy6bJsMoJMdG9cl1
uY3KgddBvTlhH+OyB/cAnfxwqof1+8zvZyGqL48o8SenjsmZq/woNVX5EKlLIRRxuRsCOIavk6c7
zopyo26K7KIiacBkMFQDP+LHCt+VAt5JMWnlPMGBLbyY3ENY9MCVAR51IF2KDv9MXgi/5N9Eryb+
t2ZEOgsJLUlbAhm33c44hIOajavn3AZ0jSLwwYCISaTniEE/X+uynz+a2r3JPppw6FFKlS9f7o7L
eVhlk8oxVg2hiov5tf/Fa7HpcZkCxn0Tt0bUqpgxjISt6rx3Wpo9UQgB7cUT9Zz2UN/NoYeKGt+Y
8tXjnOih5ZtIy06pXQjn0ubhPCmhLnyUw4AiyW0FGUauN3n3mXGSn5WCXg7iepYYbx4197CRFnMg
lo18BrLT952OHo9OyXR64P/OCTV8D2Fg9TrMxPlcQ20Y3vbYityBQS1XhERrmqh/isqlP03XFU1P
Nftug33jAKr1JSTn9Oc4Pp7/HwTL6s8fQIBC4RirAv1uUnV5HwUi+RIHUJXiAgEupqfBXbhWSaGE
QFMYni27QEgWkb7KlKIC+3itM8v8FrpEAvy1zDTj3yWAMQWmkK+WzfBgKAqxXvVGLoH/kZVZ8+8B
ZaTK7JgeIcdE5f4fYqZYiL1pyjuEvmdcjStShXQD9GxXU+OG9QTXtPhHui85zDYZIaKWTuBGRFLu
MTnq1dAS4WfqIFLvjoGEGZO5HyZbGLBm1vFgpGHDSvSPukR8iNRuJHO7Fgr7oKuWQQI6uGaYApvA
SlrCT0ZxFe0At7VMCRfa/u0X4V6VoPSZHuic8GLGWO/ukoz54B9WbeKoejZcST04bCSP8ZMYNGA2
gtAFhJHw2N3/NndpZfvB12SW9e5JMuxxNhpSAJO5JJaH2W47ONJuPVD00LDqDgV/hp8Qri9zNv+P
9The3vGAWJvBP8BLY41EyHPjRmJ7p6KySqoSr+UGIHB5lvQsLQHqMfi5FG9CU3sf3yIvP+R0lG3X
ANQ74S/JDnYEkmk2CmL+Lzx4UonrhghcRFuiN++MdtNf/iRkAfe1qjgUfHf+2A9Z36o+3fo//AZa
xAI1FOHfgNFFWkygs8mWnCrvSOe8erh0RC8fpyIK2+H6doiPx8fApnS/9AOeEz/Qg1daxq1PIxah
ztMrn3Buu+XP3EHNblVluGH36HS6gC8IIR6BXdlu9+ig7Z1hYIwz/xH8ychFagV8GlOfOMAKty1z
59Fi3Uykz+ttSdR36B0zNhW9rfU2jBm6aoctSE4UVBpgFJ0I89R4jawq78v04VZdHu+gXfc+yt9b
3NWRWAfrK1EYVg+sI3Z5yIjmWE4+KK22hkkSCLVYQJi9gUOUq78K2h45fBEMHfh5a7L+QjwdHX1e
RoYfehfB8ZfxtSoKvEhD5f03yQYsw6nulKaN+csW1VI30tiP0GktBxJbUmQ48Zoa0BZlVjnMFVAg
uF+1CopgdvyHBUBgjuFeKyAFS5RQ9vOvz0VncmzjQJ/qYZ4ONjvbsa62VbKY9G0CQaRXs0OyafEE
3+Qu2SYz9xlG/V2NldrlB4ECZpELf93YNjlkQLyGdimQfopXsl74/1oHI31UY2bKdY5KemmLzKvf
eba/b7ZRGDyW1TziTtDzvfj7f1fw8dZFn6xpMSvxJke1nMtcku4TjYEoAdfIWnz1xqpuR87rDmnW
PjWuH0xdT8Aii+FzsJD3VXubBwBWEYFOPPJiHEK8LmceqA8pWaRzr1kFMFzTtXpj2e7C02bNMpAR
5tULnGKO+T9mGEoM+eHMm/aPwAjs2l6xWNaffF79yMjcE6ZMJXJush58cDU1QQEfj6gtFSAIGaFK
y0oDPzh8UfqxaCOJkThfN3hXl2EGD/oTOG9hw2iepYt4snaQfa9Tkz5zJ3JADy/d5KHeZOu+HD/B
rTKbGkZMsLdu1Gb1MPkwe5DWUMgoZAxj+YOMi8koWmcEPTEh8niihIpshNqqkz6eSx15g5izaGxz
heIz3S022naNOcJSVnfZbfkDZz6+SeGOJ9nE4EvRX/1w+AzB9oCRMeT8g9zaPYuLFpfGAuL4L5qh
iC544MsAghhjA8yZmrgVrJirCqGT/R5uLsuGUm2d4L3y19Dx+EPnppdG0gWQWaMeR48G6TZJRSPG
UWDKiwp+IE1DnTJQBf9XvdxzS3Ut6JsbH2wALpCk4DueEOCBZ9bXCdEM1F8U7N9rnA6WmngFhPUg
lE6n9ePNxv9ykG+NEASxkJQ+YFo42ReSdGjOPR3dq9aCWXUKG19kdjghrvGdS29hMIJIp0+l/9fj
b+va8znGY/JiNswTwlHjuP+ghjAYC56mGG06LAdS3lF/y8ulA+RNVvJ9D4ylbMQYJldsZ8snUUxr
mwaNYsnYpErLDOdKbcnuoxieSGFX+uXKlzFGi/ekvzlreXOz5PsK2o+C+xaUy62GVAXnUjI8ZLXF
Xt8a/oM5tHNYpQ5/r7bIuTEhxFSk9cGo5aqyBCS3kwhkkXHkhuRgGhhhO0wYQU7M2TNhsywaD3aH
qlIXhwu7TlEBBJB2zj36yxwVLW/38GedXqk0VB+x9+J0uSz3uBF4H6viSjexZ2GntslDquO8kA/Q
sAKY7gK9wnmxb9CjzqkZydT3QpdbDB3lt7Mh9/s0aUmQEBJpnYSfIdAI73NG4Ds7SQ6sYHaqZX+4
+vK2V2MisBWIZre74tfMP5zW8s6lNEKwLaD/0OyJctNL6W+zLkJjlf42ag/I/AQ1PRs9vZYnLH96
HhWXqCu6t0SuZ/atzirojAXp1wxnNDLhoTlrHcMtA3DYPLH+Dw9l6r8Scq3dvxo9wd3V1bFZnCHW
h4VJM8/YMQIKEfXDg37n/zNtCXKq6eUKvlgfCCpVdTiN3cOLBH/pTwJxz73cdtAqEqGH4Mkf4vYB
7dsieHdO/w/1ukoKJJtXuEnfIiOWs/jvqbTJrMIdIRJWr88+3g8SLTL7lyuPDfUVWh9b7r98rpNy
sqvfzjAMqQlCNCBvc8CkhnAnuxDtw6XfdnaciUdXNGKPTdBaGoGPmaqZcUvc0Ze8ZupBgmjOpqKt
wX7iF+2iUZEx/RbxueSlycxVCo2sTvrCIhX3LkN5fsXACVorhPZ0pcIE5ZaF9DukubVwW5ywnuD0
6ngK+ZdNBvuS9RRs3UKmXto1N4EmP6SSUJdEfon8yuNpzxK6YXvCgmttTkNp4WS4LLmsrjjEzH9u
Fb9HjWuVkHhxxoMZdRXvstHStwCIIk0WkeBFVjOOpDub0NCjf3AAv2pth28/xQgYOjRx51rctem2
KUBEyx7rTaJ6p3+h2LZNoy0XCCdYIdsQs5yUj88oeaF/QBnE+7dzs4RMMMCqZ2Rub8zLvJZFf+Jo
ngykxmyXHSuI/qsgaXplm1XRNHqIHdKzAHxOtTDP8EXYaabhTh0Osf7nht+RXsizFViBE9NDW4XO
2ECW4weDoXT9Ppfnh9/vZJAm9t0POWTH5/5DYH7tZuNOBqfsLmqFKPbO3R9wxqphzgke6S5tr9Id
agANtJmd35kU4BaBrJFykbJ2gnwbnEiijFBQVYd6zmApogjnZA2YPfZ8p3heWaScvhKW5a+8uR9M
Nk6hrdKqh6LK3y8zrbUNfJr2St9DVn7tjhnCNR/Sh8ZprCv1Xuw+t7Ey
`protect end_protected
