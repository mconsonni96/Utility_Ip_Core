`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
m70Kie5Jrmq4wqJYsgEO7mxsdkKilrPIXzQjHZOfNvoKrCzCLBMEAwICtA9BrP4dLwzxWX9azKgy
GbFprh5c5o3uBXnV1edtOzol2bW/dNMh0YpuTR1j2hFGf9yDEsBBKHKFNkqpd3b2T+QaqZvAJEY+
m1gdZEpXycuguX5GT2UCG+90vJUtm0yxC/Ah23WawjurWYorOtCvlVH0iJM+OtwoZIdbMUZaKCSo
wNIVlSY9LGxokDZ8F77pAL+0zLWBCD+XSiXCGaPyHs2mIdrt6ultXfwznyxt6kjiMemKynNR7cCg
74/nBeUvG708IWi49bV8kTaaYbGsdtz6+hCdhg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="bF9f4EAOAXSvlnt8dvPjrtDrAAFHoVBDK/UTHw5nJ+c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13312)
`protect data_block
7q77gXXvVoRPm+GUs5jOUIem+WjnkceT0F01PR5Nl0vb3xwVtGHWUyfQ/N9m0Y9W2sDFktKaG2ko
rdXTsbrhP9v5e1XwQECSVzmvNU1ONLYMx0WFCtSM8yD4I48WTRYen7WoyQGEb8ptkHmrZRvgv9NY
Ie6eeD6l19wIAzTx8m+EaToh6oAgrhiAZHedFgJmSjZiUy6ZYSaNMcCpXgJshPNAuy1KHrvpusnD
HGD4mLe53z4UDAD0LOyzMQ6uxtTxDKOcfOKWuEq/VluR3dQMjI2/Vc9J9c3d5O59waodjeW1kb1C
t5vwDEJX62FAdbTOU3KnnRiK+iGonxhwMzt/b6gqo26hMVlLs382uKhA0MNtotlLcGI8AtiV2y3B
d0tDwpHAjq5OTnBi00rB3OJ2NNP5K0zpA3OcSPQkcvtlgQyipUFXxw7VHvCXOT/QFG49V0Kpxz7c
hxQVaLUEEJ0Vyhq4t2efrlCs5l27RtGXkzMq6Acr6/jpJiLDe/+G2pTNxQoREiH/a8F4zFKZcKfd
zHdcC5lw7e3o8Cng+w53CdWZ7L59HkIKyyfOYtyHBcnSszbN/4+IZdoZ/EhVS+Ds6cX+BaKHbzQm
fG8dN3Ui3G3RVzyruYfw7FZEyDRsu8uz00zUPyh5W8+Rlis8cu7KAYVmeMYhLydI89smN+3bx/m4
non8CIx1QDe3oCrQH9cTqEOtikUd5Te/C5VMA00sAQJzn+vxvCLGRIlxRZnkRpyhAqp50pPPFl8x
4zxcTx9xjo1muTQp5XLlBRHO56j/k2/ywWsGWJqyyHmZZLpXSv288ay93HRzJS95VOGw9d0tile9
YYcywZLxSvn/fPiNeY4a7ZXsrJrYbHI/YdKIWbyBXmvUfcmLbMJq764qz5rE8outPFdFTyqL6sWp
Q9/48ALo3CFkOgf83VXXIdLFdDAI1lQYtiTP0y8LYqmFHu6rFlnMR+dvtiLVfPeyzjlj+nV98U0k
3cBrMdmySSiA9IHN6V07FqDpAldG69ESHUhP35FM71ySd+KJfk5rZn91C23SdWqso6TchbyTjfSR
uQO9WKi5p2C/EATqkdbpEOk7WFWT4AWVAg13VItBUjspctvCAer6lL1SGnrXz4eGWWTgeBUS0AR6
RqeB7AzVLeV82yOUsAwVgfPq5Gf8yED/IxnE9UQ0VfKUtD+9KBzkMaAaWiK4Np3PtX1VtMxHR+4x
jdQl8urgGf5EdVS5TVe2OCQJPXAxrHPZQh3SvLW2PrX5XJ3q/Ek6hWAi4ahogZU4uNqcZs/j9gxv
KOMrPeqJGojcOKBRg3OWMwH34NAj1pg6HhEqy8h+Z+1woiBl2WAx+BjTCe4ZDBFQqM1BLD/U5MoV
YlkeX8RJ0tXM9X2DMulS06UJ67Bvoun8wNr1vKKtLASkwBm0V5QH2OzK3PDl8dKLetuS7oGVOjw8
3D0ihbnCP2XeXC23n91gDlBkQMhoZHXzLiqnt0Y2hTiqcRQFRxLJHLwGNYKVrGu11nnDmvlSDgyk
OJ+FDRCwQfdIo8ip5dNMV8yjL5eTd0oY+X8lFbB0GMg3Q5JzWlm1qI8HBGhXbxhPeusGXEzkVKxo
HLBdStl7LQB2Dj5rs7Heb7UgtQMpnTtYysOb9fhE/Y6YG1tYnr8gSfEyFAuPlOnGCiQsFYGmCzr1
B1wxnFq9ugUPHds58jTS6/66TbsNlbA3kKFnZZ/CxzLAz9bbnRrRLTQRzyd7bC5CVADF5O/DVGgn
hDdeCjVDrKJs8xPndRquwRcqaEXIDiZv7QYXCdVKTkdq3XnPrEEFI3kAMRbSTo1FyRt7/dH6o3cV
CN4moqq7FncmHCVTzDn21pF/giM7txni6wM4nydkQGiDEbtv9QxEDt5hPnNG4YUuHLIzF2/DaCJv
52P6PgLyCtfue/gvOfY+LjEHSZzYxt1mF3v3qUs2MJKZTVRsmJQhQ0jrxGx99fNByoqE3sJ3qto1
z/jEahLMivHBixOVe1q8rdacsq9max031IIM76yuycPUBC3K4A7uPW5ZYSfHADAMPbym3xnKvT9x
JVPDBILHb0Xdh5belHZrLwVauq6i6r6e44aH9IIh0LxW6a73gqH7RAnUhMAdzgPv+SIzVsjG6EWo
ogbTrOQ0jMHrwDafz8HAFvNjFRl1aSMV8HJiVM5L5wODyI14dYDU8TLQGkf5yCxF+wv9OX5kqPD5
68P0dgDqttu/CzbyXb4w9+8AEi1uxVrvd2KROJrXCg9mr4c44xp8m+Zzaj95GxcKjorpcYSycMXo
Cwy0WTzI5FsseIfJHfz0x9icz7qbfwqcZllc88b66h2iiNjGJT/3mienb3r9IkFyibYojCanGETL
wijUUzPNqBxAuymarFAiiZUavg3Ltf968UHrOjaoqgDl4XDALCdYv+EP0NqqAoOCcgF+FOfVUAdH
BjtBP4yj5KiKPAQqeAAbpskQMtTQw9rZVRtQ7CLI7k7OqVd0kHb4037lanMWtXsByS+M/BpgLZOC
+/DBnmNynbacO2LZ73JYk71tsf1zbbx5f7gNUBIrYt9/A2Uz1DKlkYDt79LSNQpfyetSAb0UqeeO
bUguHnI3olFM5uisY2yruprFQzql3ols218N0+vKh/lzJlsjvJooAHvj9wPIpDZh453bWQI8FPH9
CD3S7WdGqret3uytdTJJP8QEYWo/C2+hVdmVR2BVjEA+7MkhWaf6xCIvhz2MEs3EMOF/fJ9ri/jh
xgV6TYbvprzmwyXQTiew+XFHn093PVlY4JvD1CTt0kUnaOMPc7tLf3EiYh2tDWOcYG5gRPH91as+
XyVvu0ma3yCXY10exOPjlf+b1xZ4Ws1C9g3n5z07w1D3EjUWuspDpdQnFigecNbFIF5ooNhei2pR
uVIZaxjeA1FHjGzcztcZT7ejai8hUJ0cSELd9t77hgfV+lBRzfSl3bTQlRV29msp+uQjiV5OzhUj
M/qDDO+MpLhNjWCBeU542oVfeFjp5sSeEebt+ZW1NaDCi8FurxozQWbgzbnIgrM7gX5WtxIga6Dv
cZHQ/h+zwFl0nF7dZ6+D0CawuEafG15etYwHCXpsp+y0kcmUpAsPUJZvrqL05RXuuSKVVbk8F5RH
649xYQQW3Dj5OII5xNmI18GRZ/mrkmHh1HtATHr5nZFvll981RF7kM+AIn9w+L+G0uDAKVM4h+0Q
0vu4fdGL9s7cxV/BsSI5lj78CXxccFrdr+zruDUh6XjBGEa0uM+HLvBlTlJQOJjrtL6s+fncQ57Y
wslt3DrPkhWHHi3uCkPi/cYDJP0yURgoSf+1wgka58R0hJ7VZ1oL2J1TffD11ttRPReJ3vzfHEtE
i72R/hVpJYQewZLo9SI8Ykl8wzTZ2mh7TKxzZiqO6kEDO6lAEJaH1GaKbhkm8ervLo6W9z6EZVUy
IsUra8IVNcKSkcl9yTTYmbGIvDH4+mHtlYd0C3j93ENG2O+CyUuIWv7Zy23uS12AmQAiWxMzBx36
zalfz99VXqod8LSDsMxZJsGZ+XUzfKgkp4ZWj7CcSTl7CQgmRJSuh3vdUDdQI8tFBEdjJPGQS0u+
W6h5u26C23WF2fppEYPkYdtOvPAHJL549/x2EzaT98gJa1zzRKW+Kea3HoEvqSzNMGfQY+0ceIAa
PTCFkAcGAftzyxhqF4FiUEvUBWqqLzoj7EyegJq6dlExQO3Tbxz5o5BNE8hu1JGDOXxhvnrhLMx2
h1LQHEBOpKH9t1QKA5kgoom088RzTcAFPjbcDOpaLSxfFroOUuKt54adMaAhE1cWIGH10PHb9J0T
daEJ/e9LN3BQ7BiOgpOmEe95q+jL3DoY67Yo3kaQ5bstfz8dLIjs7VS9NAIS0wlMVxfegvZyLAAI
E0Gh5FMpqQKxvhNPT83ih98TlORTRIhfkF+OhDovpLs3I0swyT1allwiW1rksRbHN4lqHa0xJTLo
5oQIcQ7Q1nVj//a3lTkegAKFree7CPY4/4bzMV6sc2TfuEC1oA0E5hn0/Q3+eqsodPUBydsQ2MCt
3TQ6E6yw70OKgMxWTIQnj8eiqL+rzkBzUY4KkK3Y+yI78oqT+dES1lCm/JFLhEPdYPCsMeeUgxpR
lH54FCFBfjqXoKGMql4VHMH4nXEdAFhe2Z/84MKqDlvWT7E9cCNm+Czvle8mdgqSCH29U4GPqSJD
PH1DTZboi3BE3DNTmzk42y6/W1OZKkjDZ/RKEOiaWZ8dsGQrSURp9Ljx06xWm24rMhy3a2rK5qd4
uGrkFUUXh+n3atbYqM0TOFimD8ZrCqmUaOaJPrfV4VJJmkdzVmrDkm27qvTBNsf4zhU9xaXP0X3N
xhIB4iwLYW5ymhPMGEqSpkAOXUI/6r/FCSZx4rlEYNfnElq7837d0nKJEwcjMu0keXhKik/3g2tp
Dbce17wQca3r0RE9qX2nhbntpBW1UHhPDWwvQmmtMD2m1BtecdW5dauN/a5qYcMQJ1RB4piovpOh
vvZj1wuSiv3mQst4en5HPPLCYehORbrkYfev2CGS/tFWfc9TExXQbKA4o8N2/wScS5Bq3jPPqGi8
s6Wyfj+rEkIkNt13ZmNAvZSsPFWHC3BJINVOuDdbCyzfLIBOhBGe4JZ/Dbmrqfa5Z7HtccMY9fGX
H0phQg0dHaJyzFA5QNcfrQkB1OqV0cFUKwGtsM+astTfL7oRtyckZcoHSmR9ezlbVhnpUOl+X5ja
azjE2bWtnxz7z4/fZ0u1Q3B0KlVJNKqmEccceUMVxfZnF9tKTCdvHVH1a/q7q5AEhVXgMBSNQJLi
LowH+PNuH9u6M8vE51LjG+362wh5kldf/zVgfkghbkKBC/2O3PYP2xSwJSGTeaX0OEQpU/wgzXUm
9UWVbfujnaeCK7BSlRhGxn6k5TPHy3OPSYi0bxlm/O4TZu2N66aPf74az9Rql1cLmzDp/PaFZqpL
xT3x8Yhy3U8Ol97wuvAnNR1jlSgR8VOWbTlaHIQGZEFHaQ/ke0SC0xmRjPT+868wZHR1dvxdb7zo
GJkl4QTkp1Mo6WSE7v5+pQWqjO8s12c5tqOeBtjZ7f1XvW57w8YapuoVNn9umodB7srkarStNnS6
PEzFFr0UuD4mq7jUQafpBNjDcJPsHPiibXiuZAddG1WWB/zfxIIi7bxe8hwmZ4Ohf4dCODX9IXEH
8dSWMa8EEaILS93v4A6fyOtsAyaUy2D/2Q6/dFa9arp1JPKsSuTgNruJBe8X+iGu1evA+7aUv4vS
9kKT+oXHIQA9QSEMV4BCv2tAYbPfHhhTowAjCnKUhVN6epjIe35IdVCpoPw+WvSIrIw0okLNuJDL
LNrLE0aFobyX3IA+pPmT5m34cI+vwEhBhNisHGXdxXgFo9+w9S9lzVeDmanF5OkBkbwjb1Y2Xx2i
E49O1hAde2ofPeD9W2OTTXw+lYx8vl4Sa4Z+w1UqYGZr5WVwdoUNxVZ55N/EaLRY9dAy2QHhKNeK
hP0KLlKEqhbZszM3maq3/QQdF3sK0tlCO/Jymh6gNP+Dal5K4DWu2GMVAZCjOgGyNhn1+9MM/8N7
urETZPjJmOomZ0nr+qsVZgpE3CiWF5aCwMnYq0xNDx6uayzMHXlR0Bgr17KjxQudjmoWRZhysO3u
HHHTTDx1HI9/KTp/Y/airXh5dHa1xF3XQraOrYkzpy07+xgLlmK8W4HKV/KhdSPaLJYlXHlFlMoK
m4+FmWPhf6eqT5BZBgUJfcCBW+Q6CyePH9QQBpWd1JVF6LoB9+f7CbGbJK5O0vt8Q30Ji2IlgxaD
baivDBRgy666/5+N0mIJ5Fmg9ylhQ/xnV7EtJ6hWjLIaV42ELl7OsKM729NuPAPrilyUHEQYNbL7
DSqae+XMItdcpExcrUxI6fuaIkQTbqBzhGRNI22MurA0/T071FbOOXvSIgiQD5sYhUe2+ItksPGj
bAVgtGj43nQkuhlAvBubFB8dGFYVR0FK0TqutZLaIzArLvCXj66G+pGU0BzWH0NSDbooz29RZbhh
Bnfu/Z9JUppb6it7MQMEG5a7Ws9/e3Z3Hqm3uyG326lzunnHTPcKVPHWXn74oHbWGEdbaAvxtH0/
OqGmsDxbBG5KWnqd697l/WBv+6g6LKbnOyLvEuCLPNB4ZAuNtvkEdycsTQhqpizrAjVVTFEAjJ5F
Cs62G8L5qYq1/N0xbrhXx4onXTKcV+3jZF63lGgjrwh5s+119kIE+T4aguRNqmCYLv3adswvJAWo
aHmnGApbowEoekyc+7wib7ny/Cbl5QKwXe9vesz/p15SgF6sJydlaXGXtMn53ctkaOnkv01rn6pm
jStYZny8sCEJwJJbQWVjgT5mSvTNxbSnxq/5F2jxj/oTbH0blzFKEhHnpj252EthSIQcL172osc6
xjgr1BvC1LaPjk4INgdQur1AqYXsL85JNtZDnP+TuGTGbaItzcNLjldwsDcVDBWWyBPb9DbNVXPQ
uDEScqEBud5nPsF7J4x47Ua7MbjS7gsFBZBTKAZxc7/p9qXT+fCdS6SOF46qUyOa8zIC0XwB2yh7
zd8d0XpoaxSYwWETT6gCSxQxbIsrN5pJpfAedj/bGaZIiJ4zJRwXrFdQVA/oeQ0tb8Ov7sePpibZ
Ys+PJl/G0VT/O1dS3CMWQQwo61FPTfNPzVBgmf52unaJ+/YIXCzqsydSJANQMDapeMUEjGTrl9nF
EDWhYnAWsDc2uCnK5lM4og58ssrkiQ/bJXzd/9Kmg1x+wcNZgVyHz+C2zoAu13D4Z3wx3ty9b9LJ
ncGoxkpC3MvPLhKoKKn+V+odpAqxBz6nRyHMllcXk9MdewZH6K9knK73O6vbHFNuORONwGkUdF9f
3hqY9WpN8QOkyTb6UDnM+rc2i3JEBbWa4I3ps4diuMTm/V8xp5lh5fkYZa6IBYQfOO1QPLLOnRSm
gmlbC2wRfftOR78pG/f/mqxL6oz4GrQKvnE8Scozcn1OGEzFLVQqIhSmmEvh81jr6JaO9GfOlAkB
bb5BXzXBJ00Sq7ngGJxuwjVu4mCLajuhEoZiWFzDFs6PznBtWnMfbYkw21g+UiE9KcMbZmwAvYsE
SMq0jdQbErmquacxDipbQ5QdAbAFOfl8YNXkhSdaqptYncEqRkfSuKIKr++e5FAv00htnBZipvq/
PYQNxU4EjM2pK9SFr+Tu7X0m/Mbs5Jc40oTKEiiq0P1rwgllh6mfBmaOv4a1eGJA1HKLUlW/HXeG
E/zLXQh1FDX/K4cbBlBmk7y/U4fkc2E7iP4uQCaLlyFzuj0jYRSKTNogAxsKkCOQOcZa3DNBOPZP
PuYzzUKGdNzsL5gJb+xbnOdh0LRubjymSwcPpRNsRIXex+9aosH3y1+HD6jaRiOfh9zhfiTK++iG
wsywhbIyK99jKIzBnR6M58FSy1aGZQqgIuoYBKr+hC54QIVBJSmdzPOcU0QOGN+oFItNsmaHh53B
Q78CJUO+e1QajX3+DK7rmo4Q/wxlV6YmwlqaScwxy9h01gIUmyb1/TKRcSyO/OrUW9I22mgogtpV
+KtICYlwm/fE9BRA9n5ZYSvW/dlZMpxlEny/NdMf2r45fdUICuf+ilHPDb0NMqp4mDTcEkcpdobw
u4/0g0SEHw1DTU7DI0JYNQdkBG2Y16X6IUGFndoFTVgBQ/JyW8WynJaxesmOElcXY0phqqpAXCbv
Uem5mfG+UlpVRNt/xotFZlDC77mgDlw8ge5d6ssxUucI4fqK0JO5JxwlEomwltRWk9JdMULAa1k/
ZS/uvM5cmBsFXPpMu2BXBkOkDokZnhEWzsJ+6Ak4bMp3+KgeTTG3Z4cbp/9cTb5Dhj7itXWLSolZ
mLBZjTv+SGsm8t2cr5iuK4EqewhfbGfXyjPJtnrKMCKUC3mIwXI9uVGzozzf2RG/aoRqkhx5oQrd
Ac0VIel8tWWYvU6gURKavTRHS1l7+zJ+m27FfqTNuPHyaDwR7VCMWDtYuj0q+uTqVNy9+xSKWHY9
2BURe1LmqPOmRitHMBTZIjaLwI9x/71ZwvE7RVR+S45xwkvZusZY0PylRlhudEbLl+UXo8CHk0NB
37KsD+lIhXmoKAS35kODm+uJFYQ2D/Ctm0wcrdqQWSp29NP/c2KIgbI0kRLzNzbMTuAxzgz6nAAD
2V7NjXyq5O9B+xZM1ih0T7aElERomaJrwqXJtTRVIOJY3/v29/BTXmwySGgD29bJjKCqgpOiFgMM
N2izj9LI7d7dZz4mjpMYEZyYNsW4wSt4xabB/d+CZ7osBDhhseqd+P5pxhtizJlfMCYbdgFPZMJ2
3RU53XTTbgIddK9PQlvIwVCMxXl6SXSlNIBJ2ro9Y7ArlSy0l1XvVx8fl6mNbJy8/0/2CmOUoGTW
4d2s0/yRuiAZl8bRtfUaDAP7AyGm3I+yLsklfv/QwGHZ2tq2JbZIPhBUt+/9v6VUBWJvhCypEflv
Nn1hbB0FWjXL3hxgH66vL/C4447v3hkKB/Uv3gr3Tfz5yDY3UTbHhEiRwoHz/hN6OCXxCjrXe8RY
aiYv6Ke7ldlXeV1rhMpW8I9sx2a7W0lo+bT/gpcxPYmc7bO6cYs8AP5X8QPcNk5YLMH70fHsjylX
YWp+l4q8k3d6qZotfkJPGnDINxAukezm4Ttwlzz+A0J3pEqvpz45BFITqSuvy01oFtVkO8U2jM4/
lAG/iO17OlrIjxceTVwo3s9SQdTxKHE80E9Io7JR3OvtQLphfMtNKjcfZtCm1+gpcE1RusQXAzy7
iG3fWZGU8J4SL2agE7i7i+cmOu5ud0FFdSYlRvgJvDOSNH524bJZgj9GxzkHrpFiwfXW3ephYfd8
MwYiwlFW+yopqE9XjDSAF5MZWqKzjXDEGGhCSjKWKmNQTtuPT2qcrsQ8ND/be2B1sWoR05air5XK
2g8kaHpruS2VjwyedQvFtd2zqBkjB4EbK1v1gU4B11xsFWqaYh4uAYXvHbYpOY7pvtIfNTPegY9a
ge19FkZKxJut0XTytq3In+N31JEXMYMvOHM9CerXb/ZxnOajslsDvBpwaTQ1qmY5bQNJ2Fciqz9B
x8Gj7K4sCS9soY8mYJPGfQmCbU8zzmHPbkB8LLfAM42o5H0chY39NEzNksEVKeEeZ8Fd12/5qW9g
w+nHrxoSXc6BYFaQwf2gUocTZVIlGriu2JWdQP6ed3mo1vTfdxFqWOvUalwWe3rH0RICftGs4yzV
F/DwPYgaLXc/X6GDPJ2fiZ2Eqd6ZUGkCExr17iWSfDjNAGnA4SWTUOgjJhpRKsT2xirE2K7ehU8u
SJa1cy1odcR2lCRPY8b+93SERX/QTEk8SNjA4YyMsa4BtPBHWqtZ3UeP2TSJsFOnRGOhkhKuFywq
PIaI0hIzwOZXTXdVBL7fh0Op9ONSZZgtJFw0tt+wMIsEHEenqnmGSWtYfmX8t0LLXoxMkn/nMJon
Tu7hjmd/iBiakRn4qCxmpM0fMPgw+A2HaeT0NNAuiwSw9xOetmi3He4sJA1yB1vqdowq9jDgkJaS
CdqBH6KjYhpeV9pHhMjKj/bYU2e7Mw0pTZIWcn0VApbzDR/PuSm0LZd4z+9OxCw6dgAO94fIjXNw
3FP7z+pBGYwOhkkXd9UVapaDGFm8x++gY+ddDhjEp+1Lz2yWxPoPc5E6mKINL9MLmpe5qJByWxnm
ypFl6hVa0iUlGNo5us6q7XJsyouaZQsAWrdztpY7mFnT5DKMwbozSNOgg+SwAzm1Q0VuRwI7jKJR
NVTlSto8AF9CxU0plI6gGIblfIHArceu3T2mpVvcPytDNw8a9q1Kt8lAqXTL4k1oaMloAsoe19jp
rqZqdeCQZA1OxfI2DQDNuUJVmgf4XLy+guaFhtXAx9nd+q//GCazO+ff8kVUbbVTvxePvMMsW9j9
OJ9MYnQxN6eHjBlDiyCDGSpQnn0u7OCbEuznEiVFSY2mpeVCHKw5tNnG4mrX8p+pblUbPf4eCG0T
ZLvWD2TB2Ko+Xd8WRnK7iUdyKyYJimfHnMD2bCpU5eQ3DoxWdnllD2vOVmWpGDZdAKp6+Ou8h2cX
5QnP032dObEcs5/LfqWVA6ccEQI6L7rZ2Iy29vnBHhJRsW2hqBVACEq29kRkJKI6ayIFGrxBxu30
RwoJrM3IL1QFIsqoP611qYxrwLOuNa6Exq+kX+BiQESTpF248gl4lt/nO0Nx0lkyh8F+pJqmkC+/
WUpsNDal7vhxhgbVkEfkzyIOm+yCvrRybZcEwgdrdB7ZifwPjJg1cWGNVXL8X2ZWhG9gSohNM6t2
iASpXxadKqpN/cTp+MjDOIqwXD60D0a+s2K5A3KHtNOnSuo5nKEK0GF4lXOA/nR5n8pwgV9trSTu
y2FAh28BaL3abIeqpB3SS5tPJUz1XhxEkW0Fn8768J9oL1BAJZQuKBEfXnoEoonh8FhCNfGd/x7V
goWIbh5cFLyTXpztVlT1bEU6sCUkWbi2RGhpldi8vpag6PdZjd8EkGlj/xmIKJJwgl7aPtRyskh+
xS1EXyr9x3S9/ydd7t9dUZLq4zLEcxRT20TV/tYUFiKWsh5DBnpsRC+Q3oQPF8JFZSMNGIQVD44z
R7vAhD2O42bl9mGfmOOw1GQ9RE95EoIygUwGsv8fMtjhhezaz6zMPj4xXrgh1eD9GAeweOWowukT
vGLvpsqWL1P/vK/vH5fNjAg5EttvXb2C3CoKu/w4Ww0+3MXszrLeyKjnmFDdxGaukBKj1HajvQwH
CNbFcPRphPvA6VIat689LUnFKnwstUSxS6QEttBor287rcYlOR4KXLm7kHqnOEcEgi9pdbqV+svh
coxG8uaUEID9fgWB0zwN1AnVfrm9iXPXffpuMg30TzBZfESZ32JLvwC5Yt33hyE/IQVCFttHLwUO
ti1DBTKVsVA6C+VL9IIVlmO3mdUsBXCHBeJ0SUnfUO5qlcQOrY+yIOdo01ryteTqABWgCDQEhxUH
6LEuY3K8kvCmnhD8d8Y1ilSIWnb5F6RYPHhJAoBYpqFNoFXxKrbEOGPXbbe5ZBjZ2giPqDmXM1DS
tUj7/11idxJyf0rgzR3j7GSy+slBYnlFgKvG8Yeb9tX7xvDBzXzCq3u2DKJDCvyS2KQpA+mr9RFe
BP0TxVhytDUVRKhp1PZiIu6Dt7wocUn0C+IGMI5FB6JvNF7R/Xqk2je+W6GrKfKhX/A+wKuFce+h
zk3ROLmKIe520EmpdLnHr1E65yf5FU6TTcTLPzKOMFOXsqVvnuPQDpoMMGsLmDHTkXb1qXwGfbY6
T8uqI0WuhQTv6EGt6JfHchIVkRCFVckmtF6HFx6rgjuDqG/sCx/vb6s9S1MaXGbjfpApJ77lcszC
zVag4XcBC7fDIzL+Yinj1XS4wlf54mvb9Qy7Z/vFGnavTzOcsP2I74n2+vZSjO6Hu8HMlT1RH1aU
ALePCPaofxwS4dwF+nStuQTS+KCU9bX/beKpnm8vw13NAJCPIWPJTUZPNdAGI6fMeeGqTWch45Ld
xQPT3+nHtRUNcgAzETkQ9OyI4bmBYBAVDzfvgBhCnDq1OmgiFHV24S8WOOtQ3AKkQDXpbwdi2ir/
Ek3/VlZlaEeNfF21WdA2JhY1AZbxn+1xPiFOL4iIbpOZwepTCXN9avO0pm8ZRCPan5sXgY07ArRQ
fZY6NMCWb0utB1O91hEn0aeRsOS0LP7qFc3wB3ieLUVViQhmjWhUyC8NrKm21N2wB4cQk49VVr4u
8F2go4T+eoU2d9j89iTLHmuq0GtIunKF9EP7vRIyKCA2Z0gdxtxiit3ayb7oLVcTNhF4PjTHNHWc
k2IGp6nEzISa3Z008yOobIdJ9yZidxfTF+2bPqkOP4FKfqpMOf64xmGOxWBdHQRlYqlj13AQqj3e
HlOh+QBBGYHNvJ3sGVMSTS361q/v4D1cMSD+T3dAu7oCZsradK0tHSOlWZ1l3885tqL3znp5O3lW
fhDRgXDdLdWxykqz7u9DP0GNfrzVjQtDZpg5uTRUQyE38vvafmcK3cM0d7hze0CIYT5D9sr/Edle
Bop8w7R/EJL+9jUhTE/Z7PinO1RfiI67HLM5hawDEO3+dbS+V6BfaYyuJhmrkxXVBWVokLpGxchN
oBpnao0axcRu+eoQzQEC/v8yz2UaeRuZq1XgUi9aND2Xd8neLyECMYPzJlwTIZcAbjnnJtg557tg
4Yw61RdUdRjy4uTzchsVzR+B3QwAyfQU2v5mHlnI2wSehYuqFoOaYOR0ah6eADuLM4tKmQarf4ub
OmZsSuc0sFYOklVNmHKC3Z5hWNbvo5axLNHoH+O544JPauRph73Lf8ErGqTcb0SXXhuL+WKkFYsx
CXYiCTgfTyUV+edYybU1jusEot3AFGRbkbIRxq+lkPeKXb9zMiL0Xuv3M+zUdZo7To4fAHRi25P2
6EiYMR3VxVwPpAZHC0fdjiT22uzGV1HcF1FUPyh3+Pa+CE2urCbLsR+Ox1ZBOQOiUIRB9vfRlwCr
wkCHc80UGUZ0F/Wq3d8/5wOelmmfg+QAnjS9wVqQwnGRCpoqMFht4VGPe96RQLhnRxWR/PR8BxGl
oLukItvVv7DF9tb3gYlhlTU+DdvMYZ3DYC+DMRvPMEx/HrIsHXQZwu1/YAfe9ShBt+noNlUbfTxF
BtFR/2gArX5UhpaEASKm39O+6C1J31auZKzEwoOOhK9Mm3QdEX6VhfOwh9ea6eNexPIQQib3WZU7
AjgTE4VnviWr37fPE9jtv2KgZWBaVoQiWTlOfDQlw2Ses755KwmuVrSfpm3CpR6AiLcrX3vmQOnv
8wWQXJzQhmYqVjgNpUe1Ur3y94KPifTMg7UXIXtKHqv8puok8JvwfpxM8bIpdHQ3Bak4GrOy6Xmy
1jqC+3j050fQWCGKKoHfhwUGdhgUTthLI9VsUy606YurMJ4h0TzRv4cJTqkxPfMdio5EfbSzzhIu
8csnnLRUDQ/DwtpSTtQgKSAQX30kbm6vmj2rq8RxROSeD8RAp8D7CWoJ6YSG927TttAUIpV4f5dz
kYNez960Xu3VD79sygdRvhXw18sYnwKlnoJAxTic5Ua9cATfoxpJESyJljSnTgQ18nDif7XXR73A
QlNTb8qdTrcDxvbsuOYpAcrnPuQGmIVE0qPLl3W4rIjCocyAJ4Iiq7jFVK1XFkZpK9/M8Er0BXXW
vJwZ9CJd/Z5syqAkzpDWex8AOhaXByaqgUDqqn4XhKo4mmtVrNVwfQlg6uUCcE0YnhWueWXV4BtN
5nWQLFncucPZLuQn8jSGo26GEwnGbusBbcQZkJguC5cfMM52zRow7vIhyEk1AySEnK96pBFbE+U5
43C7s0Sbe/LGUj3BqAEpjSQuquGZ4YCxhxxPBbLSuHh5rqrzriZBiblYt4q/+p4Zqj8NPLIOQz6Y
BA0u1+obZXIC4M1UbSBetNVGNJYx9lzGyI2e9EkNfRwX9re2z4cUzGUTxOydX77Gktj5VIhTeY8N
hBFk8Ncio5Jd/nwSnXwslrYkKC1ZEj2Yr9UMod1LXG50WZoM784kYNOu+T34XQnc3nZUduSpj1+U
OvnQMLOw0kD9YoB/1pqgEu5ZGMQO8VkPB0aI9CKl1fkK59+mgcMMAKlPCfptELlO7CEXH5WPw7U4
Haz1dK+M9nyhJRIiIKmsxOpmdNr9+3dLTnvNhQfiiO1WAdBy3auzIOtnuCR5g7BoAws+32FFrc1N
Feb2oteCRnwBjcsVjVMnutQD4H77c2no3f8lr4roT87tTWpOa0Io3tVNgLPpQtjVYp90LTd4FhgZ
1FBkMN189xIN2wSyYo3JHJWblwid9OGSNlZzE5+2nxkJMS5jYGDWOWXBk/ibyAbc7RYxpQnOou7q
eEPub9h73Vrri9vxOW6YWTK1Yds1v1gsux2+BiQhE/L2tfH9QOMjp5m/YNU05XaMlZvZAPNrBqQ0
L5tk2/i/8G6cUjci8qDd6lXt/SU8nxgKzc5s1Jk757u3gVuAQn/MoqcBVnf05DyW9ZZVvDRA7CPy
3KO3x0/z3J2t70CGQqw1uHBoacYL9cj+VNUpgPlquL3a441arLqItmVFArGgrbocsckeDXLKC+dy
P5AlHr3GMCur2OtPapf5W3cB9Ze6gMy1xvZKMOTyk2YDzKjW099vlLny1xSYK6VQUfYODrgl5jsu
vNLoAavYo2DqAq9neSZnN/3A/ZN2BVNyZIgcqFAQAuXQnhLN9fzXGSCuiXwpJABXyAVYsCobVrMM
DbT/k1GKe459ZBRVYl2izhq9/JZ1Z43Biuejh45pMt/2vKNL2Lpf9h2nD3lGbWuQtmxMGOYkMyZQ
JX+m9M5ZQ+eLCjtk8Hxg8UEXGytLXbm1avHdcfJE+UxvlKR40uof/BtPha/PdSyLRIl4bEN7EnUU
8UWmEwKmKafgDWzPG8oqTaVm6aENrxc4rDjfNaUA/oKT7tfksaUGAZU1bo5ZsGEIKW2MjfQXaqLJ
avdTnX3lKSWNJYdfYV+MlAx5ueHUg2kaP0yHeKG3PcbfwzfVLYP/18L8YmYmNxO4Jq4+0cJTuz4s
b0HvEkxdc4cwVsCsH+pcjOMpa1v4uDSTSJxKAZprt+Luc6lsvVse3Z0KOEZtdFGXdujANYawrUOn
gvwM7CNWAWW7NmAJPlD79kPdjqm8iUCIERYfcOS81Ti3dcGzDbdKjZ8lZFsDEtn1z3fl0b/WEWyl
S0tobx2++q2w1Pz252vuRXkaP+lB9bUrp9Q7Kndz+tOc6xswNG93jjemO0TJz4fu/7Ec+ht1zVUv
0as8QYD0bZP0qGX0UQtjSkG+YNUzV2GKpDJVETr8y/Koo/aIZiBCBxKdP9jvLA1uRdcQ6QUIQmhI
SiPOjVMcQZpAIKJTp/EYYmyZFXwsNh6TnV9YXSZ28kE6NXVIi7zOHXVcKuIsL3tV7/XPF1BFaAsf
2bcQ6Oyh4eklQNU+cI8pcj1Je0G9fqPBfto63nAVhvSVAivFjvSsvVjde9Fwlgruv4jZZhqgQrEg
1wGpTO5IwohYIdm3LyUimRE0Mg+9f3PBcAL0rOFrgopFhaoEXU7m58azZ/TmVEYzzr+bdzxB33db
XoaW649g/fcSwzSToHYuaoWFF15VjfTGs7A2tTxapQGCDDm2Z+h0N2siweMVskXXAKxVtH2Weqnl
UKRHFbVFz4eLww/dNlosOppSEkCMz7scgsO8cQzfRzVtMA9aRz9zAQs4Wb1wXu5o/JpPCBU5DZ+q
M1g0wMpd4L9ykM6nepP5t+7/HZ7ETwdpMl8J6Dx7qO58VEkoml4mxLhQMItnrrPn9/IiuHuTbcVb
q4kQDAfj3BVFxqcf7DTmriYJCK1UTRbY+FqDh6ZGtudiduzefF5MINzZ2Tc6DwQyXK69V/hSJx2+
jgPsRm8AIpInjEQ1UCJGvRTSWkySuc2z5YWOjTHJ3rRfYo9P7RlQMbldD3f+81owNsFcEYNf1QBp
U1FUvlxpQKp7CStsuwwVDOQocmTMxuVdMSPfAdz5xXg/Hs+OrEWS36TEXlQBKCZDvxP2sA+e65tu
3RkmhTFqRBuD7+l1/BKFRsA+HgpwvluCvk6UQTGD/zfOdd0mtd2opwWKdHeN/ti5XTv8MO7tG4WB
dq1aD6txiJGO3cgO1fbxCl5WZm6/M8tjDqdYkxUsCI7bC5i7vmqZoSVBddRxkdhzmfPpQ8PREgc0
vNhW8bJK6Yd1bwV3B5bAen69bKYPekm/F6ntwVqVpQU1fdnBlQcnvO4kkZ9YFpp56PcNqzxV7i/p
tfYyTMKB7TUvhyMsNSASym1cujtR5yoUxPyaCHupBwvOH2vA96i/21RZWZLryGkB3nQjvTKqERZq
ZAZAfKrTggok3/6s7o285QxmW0vFFCMYVMNP9tgPbNA/SJaHMm1mo1OujMidL5uu4L0AqGQ3iHNm
Yo+j+y9AhgX6zZYdlrFWkmMB0cAyFQe+AOagjo9lXEI1UNbYaTVJViT0wabICiCxX6SlRPfttGFK
vHAd8P92lZMNnKhqdlDhegxqnzCkU1CL/Jxya9Ec+hauKCGIAQqkGf/OazykWqbIgsld0QKba9w7
mCA/5Fm+bzY1mRnOLa5WETYmfGTJ5nVntbiPTFjKnBHH3VHcmHT9BDdA6+3WYpT6oSjeuCHxyNwY
BphQDEVUzkTk4DSpBuLAl/YIfee4F9UI1IEbg9H9jgfvVQvSgIpyv6bS+mDaGiJdpPU7YKqm8fnO
6xeAw2z28PBiM94lNdzxa+XAiHZrdm9oru+yOrrFTTQPDQHx4JUoPdIRO/B9dfQjEIORn01g7nND
vW7pkxuRWnZHO44DprM5EMgCnlhVEg1fld+q8WhRXFPit/uN4EQVMQDHrHtQqTNUUyph2S8lcM/m
6nM8XCjkB/slMJyY+eyibPWR8WDpdrD1ByF0NIu7WAuCLe+YdB1ObB2JiDlvzriTABe+6fo4Y2kx
EDEZfvkJKmqchL5w6hw6S2GakwXa8EPQ1iCsgS94xdIxruh3nMJdwSaY0kUT5oQ39AzE8cHGvmA9
q7jSASwyZJY66TvB/hIUjpZsvRKzfvYIyr7gQcg2PINEVDclU6WDOYua43NuzwNKnsjCkwQE61Uz
zf5kgdkuKGIXO0r28LGKrLE+EV5Ti/siNH0XpcYUWRRaYmNDvgDbDLxKUy4bRwRQpVAZBtYxg/kk
Em56eRoluX+aUNWdvJm4wVilwzHL1xCLJBAx8lf9rAZtkVz2XZwCKnf8ECUhNBxipz03/rg00PaF
3bT6RMfV4E3E5ZeTeK29o0/BmTU/GtXlx4EN3us7CLZtP1izh+AsiL/FE3/kQVMgWQutLAMem/62
3wcamQXcKZtKaPY/1Lq+fLpDswXGGfoQPcaq/CA+ehfUaF6JMPkPvdUtqDWjs6h432ICBx8iS3sj
w7BMuO1NUHMXFZfY48nQuAjjZqoQ/DNz0KiTMEsxpbbu6QMXwtQZC0fqaNdCXk18GIqiVaf3y8gE
BqKXUrzJf4BzKQdfbo+zWSfvY59MkOAIABK15iV4M+lt1mi5Vkp6QdmPQfff0HMUY56eOk61CY3J
YwzLGfgL0VG5Ij+MBlR8oWDeVo/+wiEKwq+SK9IhJjUFtzbLkjHqNHYhqVJw8VFbnIrLccjzywXs
72y731mERh0Vin/zYB1F1bsbE4Js9kAIawiDpTIDC0JYRdac+UmE6AexIVo1sxchVdYfZnL4N9oF
yEhZ7Y8QbbGoVF7lV9AIF1cNDyKfDUxO8kmU6djppB7CMgwFB/iQnZ9Bixlgsj6GtSnCjrmdXSEF
AHuUVE3qsVyaaf1oOJ2u2fRc1rhyBKqwaxOLeB6BBFM75Tg6j3+GTHr5hG2V8MnYvILuWSuWPHxB
ffU3gEv0y0GXUX/73rWt5ufj9LvJVBjsWb7ctRiUi8DC07q0wYI26i48oNnDfgHoZqfOJ6AlpGd6
PxrCz/0L4U0rVkjYsksBYvxc6wSogWl9okcNE+UkBWxGAWH67Cg+w9dZAAYpQ0lwrIC36K9UzVM1
+SrwDzLawmpKg45YcXZ7fWZs09LBAuoA6RJACpaDY5cI+wR+GhVY6LP3BD4AzLYUWTnw1UR8aUzp
e+lGdxu1ZpEqO59ocaOLDDyhqD/tEyDQoMMc5lCmiuTPqhSB4agW1RwhS5HiR56fYhOH9G23rhY8
8iBU6T6BBNxWYhLAgX3ra9JTanhrKOBhK+XQOVNpXTzcX+oIwpZ4Y62Xvu9gij/WblTLjyK11zIw
9HNob1G096pxTcFNp0ZJj874cYUngb/nSIx2R9U6fw==
`protect end_protected
