`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
a42/N3LwccVlBaY1sl5C1UM4cnOs/D/AtKC8siZUbHjoALUHbik/HZBxeZYLifXQlPTm0UTEEvXy
/sAcc+eCiUc6takELIHB04C192WOcZCJqQTZmjewlDGix1KvfqlTxSngYeyFe6UXw3zktR8JU2sh
IUNb5KgEAUqCIF4EBDxaGs85kvKSmV+HiYitAmLi9fpn39pbH1H9oOkr3Ld8PW3t7R2sr4oahNX4
z3nRZYuWgMzO/LNcBy8JzwOnBisG8TxnqYIxRuS9kOLWws57fMe66ZgoeKnrhzCacY6w62CaPhVW
iqXwiQNlwCS+fQ6mhsYyej95SHamSC07vpYQEg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="xvcIogMqQdi9NA8IDQILG2TVE1fP9bswsczBmYktvpk="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12832)
`protect data_block
QLksMOwlDUmYTlpFS+f06w9cLvrQIn0nCWXdWe3CnSbGkUZE2VOJ7a84sKp1ikz99o8Fcs1eEsde
WZ5TGiMV1m2KCEszhrRJdOZNKB2NHwuW/gzOd3Ansa3pp1y83lZrS5Vo+tSue07YciGYlpl1FMQj
2EAXOstGurLRuy+3dY+CMjhTgPs3WZx7/lYCrse74jVODz0slHxAy0xG499z9RCNJsnf2GqCwZgJ
QVd13xrV6laQoia2NkiEToW5Z97jmer2Up5y+3OSJ6/QNHyQd0u5s1VeTDXcyAqLM3i0RbzkBq1M
9e15lisHUtrfFzM8jCPniRQ8BR+FaIENVAMFIgQecWogKBH6FU0h0RYDp/nZp5Kmvp3V3e3IyYRV
ARy9nIb7K5Wgy11Q+BcB6a/AE03HtWtxDQD3FQ66zz93rVV5be1SbARXC3IfCvNvzOhO2oOhUJ3v
dsq47tzB4dzXdan/BPLISJKoqsW4IMDeO3X7RnRjiP5xZ+e4Mf5JstnZnuczOxVNHHnq21k72e1Z
L9ZssApjhQImvxROKgfjkK2PSTTFygkAzHjDmt4oHtLSYH/Vl9X5Y0A5ImC94gqI4KfUH3YlNQQA
xNtLvBlomjgm2TE8IYZoSsILG95nGHd3zXgxph1mGiSElZdVdEk+ZvKdZBY/V9tATCSnIYcanj4E
1zbPTVzwTLDLZC9lS38eToi2yZrtPawPQN7e4DsFAT+TXDmLYp+X1ufKP4uGEYf1h9QdGsLu8qFU
Zh4+T/KQaNs5H9pE/MK4uPCIlhw19WP+XSq/hrcnZRr4iTZKFLr/pMUGSEP4wTagnC8LxMTlqSGa
tMFtJ2LRcaQ0BkkZV/H4aY8hnnlI9QxUFf4Bv83b0p+o7EregdhpoOz/qrnBq9C0YQUgIPVA5RER
ILuk30dZmROe6ZmrPVI56m21YFffHlFKouqHc55/4+vxNaMm1luLEVsOBFPbD+PAseYiGDybhieR
GCp5x1b9kg3ccQs0mIf/6nM9YmLHgk4ZdREHqXDivcPk90UPg5r3XyuaRZswNVQZi9BUvPJ+H9b8
EXXO1GRAIF2m7N/Do9r09FW8z9/iSsre0NFWaMw6wNlaWq5nA6LU7+ejOhGX7ZBFG0eoA/OeQCDC
yvLzz2RWQ2z6USC+RQ2KgfxTNup9KmwjYDWi+Kg8pMuCX9DjIAOOLozvHYaD0Vf6Mgmx0PCytOwi
wgt2SoqN6rjkP+jwCIen/D7c2ZCc6L20tLt+1zebvmIVo1dNA34KtAIWthXUigB3B3XOVv3g4+ep
GksiIsQ6dL5V6wpVjEMie86Vx1sPyeFUGX5JnKuM6uWVYXgBdLSkSZ6BEINWSSV3JuKYw6bkeYC8
6wtmf1Ilitx/1e/ZrsXF0baGuWab2IWAYRdI8ELNjZwm/fbjB/yKKUWKJLCWo096U4+L2HUHTjPP
V0jUchkIYeV8hEclae9yTOO5LofS5iJhF/meSRpJIMBTOwHMcVJMPnS/rLk8m/haKpHSYEEsGMzy
35K8cJHR/4zbg4XYfYC0asXewU8czEQFlrnqQx0kdIB4s45CuBYcRx0IuQ3Ex24xL2x2cREqrQoc
lT9wYFg5HO580+7kWPuC20yJPGkj+52H9cSx/iUlazhkyzGGhr1v2yFkbLVz+Nf+naYn7e30kFUL
PBrggRMltscjBU/bVwiGzX4Mvnm8VGyZn2rK6LVNiei9xIssGGgQYeGEXGfTGMN6V305KOYsNXeN
8ivfydtfTUTPCnIepwXChqGDJyDGPALvzpblKiVrgkoXZ8bscWaF5tACIOrhwZbDUBkn4eFsGU0l
BrUhuoA4lGB8LLtIUjsHq5lGF+NHxwSZPAxBUL6z17Df5G2fRGmiXaP90YBfEZ05uL4Dm92E1net
54dulNleqLI8eI4PydNU44RN+nUS99lVbssjsqdQyfwednIzs36i466oMKkHVxvZiFH2W5WftKe6
NXBfbIW4ukY4v6X+brRrDjL5RM+gZLXtZZfx16RjZzn5HYdXmP8UZMTzDuTJ5+76+R8PpOvA4Guy
K3g0TN58kVb1Vgb/Lcd3Si9C6V8UsiwXy4zHzh9Kaz9aE1TY7FOPsnvZcwOJ6Vucr/PMDETEjLde
XVUl4PQ2gf4odfCXQ1toO1WZ8RZzDzyoNthsFjKmQS29PVSlbGlCltg6qIUzubqpFwcG72PsoYR5
eja9ALi4IjKhWEjK7QL7jZmMlzaYuucsvAwRQ+33WjJK+KJRpnizk06cE0LKldc+VMuso5jgiEvh
1ZGDbNdkBoAdzyw95sHfkOLGR3o7gZQgDfjX+6VetDteywpZiSaGKJgSxvNBMzpyPk1uxWxke8Sq
GHjtABl2B7/lCW3cEAxDiTf1oz3NHCL0sKy3tPSvSDW94nhFacZryRDO/HBzO7T5fOiLG34LBdAa
qBYpEyRiITLj4nlBkDyha3UUcQRD52eZxXqIOd0xz/QELPctGEqKejwNJyu+6+uNQjmB1wvTyGKA
UrFwLM05g8RCXMN4OM9ka0Vlt6+tjiioB70EeLHrc7yr3Qd9QCyydhnDQyoUxdS2cxfam4d6uv6E
7qlGupkY7/uapbzLfJqLk98S1mcRSXTKCIh5DMqfH9RpUBMCHAnUZcn6YoLvb4jR4IGogMXe4fpP
snYLJPUjOwe0PT+uOkJddGEdItx63wL7lEG043l0BrfPGkL+q3GQkQbAuRMLiyaeoFlYjtKLL+nE
VwMu7UCiViCDP6XUayzHzT0nnfunwxQ/7DXfXxOB64EV1WnO+YJGZ4+YIM8uF+8sjNDcaQjRORQP
hAt8hS2o+pAGJKo9VW1xB59CUrxLI58mjrdOP3ez7rwsQkQlTcT0KjsW4Vhoe37aFhRFSvspqOe5
P4bfgowUvP7ll6DeLaPS6FD+TxHRU5dVGlSI4YqjfpJ8JHEscXD3iYc6a5T6L7DydOoEKnR3h/9b
n49oMMDM8xmc8jd8dqz8RrtJqyFWkjfd7kNTx4+LMUYrrJkwLfbcUhExtBpKfejof4YueNqFCYay
KHlcTBBUgfYWf3q6tQptMc15JOnR9RtnsARg1U/w/GE/H7wWlF4r00/0fLWS0dGWT0kFj02cQFKo
TN19w4MgKouUTuWzcDcRS9pCBYngm/H+Xu5IdlENNGLrh+hjnOgMvymS97UJEiQWoPf9aZH5HzpJ
CiF/GyjLYK/Moc7+rjuIbgj49jsvtnyI327luKS5RUCeW5f22mNcJD0f8st37+mazptVhM6cGD6U
DWkVvKHObwjj03bFuITLWR6BpNLSfEKp+tQTLodOq0NdcKEhrjGEohdmwSraSGxi5RjdAxxCa2UJ
JaZQgr4JUwQJ2kefqtu3eCsg7pgZ8Wxplbm6cj8Kpibt5iC1lmfeLzmqdg9keW5y+1EGd6g65HWq
xYYs88d/N1zdLds+BRHLTueFQw+/LMTCG49mFJJvUIjsRhbwrjkUc7H7C+b5xOE8OrkHAZU7X4SQ
IHTIQY8BMwvilFVgyvzYFpUap3c9R4Yin9qpTkcGXM+fjCTx8yBxFy2GIZ2xza92IC15kVaHlasD
clK21SdpzJk9if3raxjlk+hk7SX5YtKSAxmwgZprEy8R0ek4XOVggLzO+THzL9PSuvcK0xeNnRxX
JerKBu888+iod9wa0Glx6tGhMOYJM/R5wvAkrxnRf+ymK9nlWl3WtRNGxN1BoCJsh9ZBos5RhO1r
C1+uA5MkWyg9Zf/TZ2KjzSQgI4Lg0nb6+tLVB1TSLGwLZftYJCosc97jgFMEPvvKwHnsOf0+UPbB
ESna71jojlIB6/z833VXcmusItYcDoxfj4RGlwWKFY9FbuZ68TkpPMlCmF9b165EXDMEpXi7kun0
HpC6p/wD1tX5DkeH9k/Xa+d3IhVYtg3fljes3OoHMlRNx5kDXTGRAIMVaHn9wFk8Q/d0mg6bD5rv
chmhv7dvLEn7TkRomb+Vxo18J6aDHqoAVdvV0HD+duRDA6A+mg1qu2GNrIuYWqz6QTm19KNz9wqP
qSB6gJAY30OofiOHEHfxL9fDF1RTf/FOOOFZ/EtPEzWYDOOJg4LK8Cd45U03olw8HFICuFrolEuW
TBGSuyso2H5wXEzVRVmTklRw/o0bZHD3TOzLbDDTYr5qDNRvD8Cjh2lDKnbaW02zuJy4AX+/y2gi
oDz2stFvnyz+vmjpBoNRBhMwqtXGSxa9Qbes7OFaMhiDn2XtrmMOm+IW4zQEKpE5bxIe8tVUNTnX
y3aM6TZ5LNY5WorWXNiRxhKxZOaR85t0SuVVX6x03c6qms/+IHEgfJ2klXbnTDsMCVD4k3fYRfZ2
8MusbameL+wJOm9MsVc8EEy9ui/x/fPYqCcjexnDOlWjg86paLn2YRgk1yCnsQJcGUUrRh38unIt
QS3s/B4q3jgfiVN/H0xe77rwFbsEhg/B9Q+X2rRHsuj5BC+AHWt+Ok+2XMEI/JjAH6q8RYMVute5
VYGOdZ/2C/BD0R3b/4jzdak7m223eXV88RiRM2q8S/yJOH6NER8B14o5jOyQGSgFCzO68MoH0Jw6
rBo1O6tqbFZpP1OV8E2r1PX0PDygJoQ2iHFZssZevRUAcEnAZBiRyex6yR2EfdJP1VDiq1yp4el0
LO4CuDmrsIF7LAb7M6Sd2uvwwwV1tMmRFrayzm98OhBDAqnfMlI9uU2YUzFMGEIqWzlfoS0rPI1G
lGh3GtiblMjlUfTQzETIjnDDrwjpaQ84sBVAfgoCQu3Dh8LoTo4t9ySqbZ6nw9oTeuf48w491j9U
gr8yz3fGQlBw4xG/pjdOuhF/6wTb/p6tLFNALOaWmYsz7TjDxd/E5+tx7c5KdbrRQbksApD3xuV3
6ionv9jFChxu/hWVG0NWdgqKuaj894JCNfiPLdOz1HlEqvjxrGKl1z7f22+qYEO/gafi2DH3YAUW
KusOFw37h1IuePC96lmOla33AFrAsw49YzYyM0qLAML1ZMnTtzd2Kcir0KcddFbodjcnqKPgm5pN
6jjNyAlQhCXFLuLZlwWc0KaQCn3fqkgQFJxAwO223ZMjfA9pCc6ElkMpMYCE9Vhy6xKZRs6bfo0i
oC7Mcrdck3ItDKkShCo6AuTBcmwrr7/wL8PCuCuOLaz+yVXxvPNuKBObYSnEugV28mYqbKyccC6Q
71NO/XX4N9AOd0T6wvDVPvBi13yftn1Jn+R5W/nDz5Kk5T4Imi1ZpvG/P5Q7o0xkD/cUhxpijkV0
MORheQa/wEtR8nfDjQ4TQMbGkCleHnsUYlBiG1Ksl3x3z05iKbzETTK6ciB7HxojdGuOB/1L1F0M
KwW/QfbeKrXzrSgyW+EQNVv/oJXWrVE2OOvGIK7uToE5uinWoTX6iiOAWX7yLogw2r62mIrDtjtw
c3cqX+1jJMWqjd93v9p1GDGuUbZZJfo0K9iQyCuXLRWuzD8Ee+zqPSFv2f4KDgR7asD571N/CYGi
/QlND1CBx0htSKladSqhp4kKmCcxKOlK+ymvlQNBDzcXxxPvT5isv8r0LuElGzsDrJaaz3xPFJad
r7GEKHjSIKuJnNlKokzpWsKtSSQcT2O2rFB3cMb30s8RTs73+apd7M6vPTNmSW2XYxyRoACDCoKF
78lbtiN3041sJ4yd9PdVGMaWtTwUAFUUCoBVJSsYl9ol3E03nVD1oXkpw2euB1I9Os1Z9tlTedvT
GYvOVUwrCwmkPnSEhC8uvmMjG5Fz0XAOQm1yQQRr5oPwgFbbGg0bD4n+JtmO6jso1okB2sK/7NS9
j7Bx/ZqEDHtflX9z4mmMna32AIPCX23zJUq3WKbX/LGeH5ZhC8fPnQbjWwLP2Co0vv1R0+g8yBXI
Ls0fyHVg19KG4G/YwybPPr9N004vOaaBhZ9WjcE8SXzl/wFW7lFKSRDybhtZQAntnpqo64gJZohq
KYbnerHh/ym4yykpz+DoWP6p4O1lRGfEanmgdFOsuczM9bNzC2FAlaw6vPnL+6CiTuYSIG4itMM0
+o/82Zt15wM9/4LhZm8i16LWfKQM2yCLFwEfhLuJqu2Z0o4Nhohvsofy93vxmI5qY6nspEfUBWKz
2qdfUeeFGLO88zxUZ89n/mG15cEBpwxR8RiwvAbf4KOtk+g/0zcECYvvjKw7la3uQ8hkBaOI8agf
DBKH8SChxb9gG1TMB4/0NjPTm8rK3Q3An6KRzJLB4MhkZazw5zT6yZYYcZ1wHUjljQRfLx2Kv0il
K9Mu6LLI5pWRNgKuN7hCSNwGNb5D9VtC6UAqD9+/wMyyEBXXleITQ6YGwVzWRxI51zuducVAONQB
ytUztAIDi21VTKSEsZH9+HTPhuHCVdj2bIv2+fL0dfUk7fyVaWCSMaElshwSzxN2m5cLennl/l/0
w1dcrLAEg2rwgCbRSWfQ7aW0J9wqttIemYNH6eY/X9QwJU2imZSh4+iqM+tilI69rtCOBGWQvXe4
vUhzhgnO39FMcF2Kluestb5c+7y/LnDaamGOgnqhB643DPPLGJP1krHbK0VAdzaq+7q6VZpzPC1W
fIinJXXcYqWC3BmtaAH95B8cP51ETgW/yui5hkpa7gI4rmkO4nJapisRJ39Ws8WUfrF7fiTqxRDB
GmteSZyfBfnCBF9JxYRyAMsx5UsSJORo2UmDLEr04wERv1GGL0GDGy/ml+hr4kJmmZRs440YBDED
L+pFdtmn9tGmCAPSnJ9Ald100r3/3cbjssMoXD3vj+UviKZbI+uk6ks2KTnOc3CoglRJQomRcd2c
3juNXkNhG8SEdOWfwE2qFj3QM/wOha8FXMsViS4utYj+eDVY3RbIq97ij3bEPZco2nHK3fLVSxhP
0BtRSLexFFuIVlSKn/LHDyHrAvxs8HwSBc3dUeDaRctzEJruYVRcrpxAUy+WJf38ZW0lEhO9Jl4b
Tzhj0dKuGTVAIFMMWHG8dPrSchWXF75IsgcS3vLXfsAHr7FmlxJJ2wMAtmKkDZsUIvVHmqFGx5XI
RnwdEvnplRorDPks5N9gf3Lk/mhQbZtfTnqGzEhp/Dv0Tf/Gffau/HTVD1ZY63GMSlNFd5WEPEC8
z65Ssymv4SxKynW81M0cbf6Ir86DFy/RC+NfXX7JvC7vg3S5o3CrsroQXVB0IKC50t6RzJKjmuDj
Tz8YRqRtECMxxp2sF6N0eNbd3wCDtvjetUQ83H2YeeX6XgM/VVSBfi75D+dA23Im2xxrNY9FD6SY
1zp1VKaidAG9b6SHW2SmL+xLK1stWZtLbshtTutQIPes6d0r3lILGXW0d3QAuxY1cq8/Qk2pUyBI
NpVTTfOTEYO6Z1oaqEv2F3qtmVs9HQoVD8w7+7T9+XqQK5hmHbeQ6pYgbQFWO3J5RoU5Jc/XnKIx
bNPu0YArWimki/ffAgLdGggj4mC1tibgk6Qm1kBsRBdO9gxN4L4HxDNFFtU9GuxdkM0CIqyrXJbw
Dyc+50xpo7+RKA9r42yrm/ZN5CDHU4BWR7BVTop+WbugO07INo0zWhCcaqfUZjFxykUjilvD7oKC
IPmQDA+q6dfqictsBd41oOWd0d32uM3Ij0qeRFJcROTTDpIhOGLP8paShZGmKo23OqrTx9urUzY7
M9yz9hmjj0gvLpDqhvAxl/MZb8mNsxQzwdz+ttqC6KnR6qS1ya/ShkZaQq5CY9R8lvkucO2Fhfln
IraW2k7q0H85qu5DG3jdlB91JGn1ZaUK2FI2D8qDY/u8c6cBY0pIoSKFWMNp/NtEuJ5gMC69Hcql
qN3nXaUm/9FxmbP3DfxfKeNodv2sC29On8La2k7PIPdYZldV8DyvcwVvWwfAFLtE64cLBgt3CqcW
+0Vtuzb4DQFhXEJWAVAag/npHNtRQOljvbP7FEBGArsiEGWgisfaNTMuGGd5utl4kys8Z6k9w0yk
B8iGUgTK0OP+lgehqZh1so8pUM3JqWZkz3+HIu1Ngc2PMoPEPNVvkoYt4/0+V33yD9PIX6QamW6L
at++ex17R5uYiYqhreQcG+cWswlfy7d1vn+GYqX/mzCvEcQgSMhIy97bSgwnzXiy9Bab0kTiKQxT
WPxBh8TSuggqI8BkFbu7xzi8AZFZp89JWXg0uYn1rpXvlvWu9BSlKHZsbU9wIrexClsSlM1wTNMe
0JsaaFjZF6DGeeaRKXLIm0KFkA/IC7F7E15llpBTOLFPUoFqFVKfVWaoS9TbdaJKVEGupGRxvqp/
GvH5cL7aPM5Tg3VIrG9fKBPAkPl3TQTNxXIfUwbVGpw3QdGUBZEc6Fucl199HtlV6jlM3+vySQR5
OHr81HhmnnPh+TnEPHq03A5YjMAPTzziTPqEQp3vqC6jPMOF+312fHHA1ccHj1LtUt7AzwopUAYQ
4pQoZiNBzP5WiZdnCdjiOtz2KrbdW5eZ8Bg9j+UE8JIUlGsv4RZ53FSvi20uA80dJ2WGf1rRffeY
1/NGmYU9jsgLP490Hg2NqGPXYbQ/bqRGbWmZj8cwjokaLMf3tzpx9ulVbxlYScY53kbHasYKb8Gv
OcJd/szTo2D7M4fbGJqrCyLZ4OXEsha/o4gJZqcachyvOX30druOWkXuKz0+m5ACx85ymfwo3dls
e7dMSdJ0XJkbtonKZLfCkw0TYjDlDuoAs67ZGi34PRh0aP27I4dLuBSXZ3/4SoVtKMTa9DQ9rmqs
ZOOhC3C2JHtNPC/yT5Q17tkSP2hjtJKhN7VZ18m278SNY10jQbnPTbzIxRApVCecsZtxjv6zMChi
AIf1da9/+0xU0MNldOuWGZGeiTPNrdmwveDlSjOQPJNayHqS78ijYK2L/dsSIjINXLCjr9OB37aG
VW+yi5znd2Tsq841/OnW3vzYUAFRD+itN6P4Tat0zpP4xLh1DEAOZ7eEcoseSVlrsVqksb9Z1DO3
op67/l/NP4XDyJFvtzOVUEWnc3M8XlcBetH4Iha8IJ4FgJHvf/vjDo0yQLZ31GbMlwBcje1pI5CS
j4E2jx8WQYYEDziVOljRGl9/ZfyZsyx5G5vjW6RuzqxLAcmp41QZBGgIuTWjMjWI1tDfcpFsY2/Y
7AKlE5+Dcbb6eHKe2e1rO0Zciiay6xbiZYHL4zR82ZRaPQYFMFpnnlxsbS+ZSk56HPB2tDg5eBpL
ElNvuj5vxHvoGjsDAL1VuLS31kvy8YGDfMEaSURd4715J+Y4LtrkIihF+I2TNcMkFAm10p/VtMWN
cV0w5suR434Dz/5pLpSJT04Yovq1FT8BFF6FnJrKbcFv0u2pO5l9IykoSmlKkyMKxOHJBHnhGW3t
ElpFJi7QgX46d9efPwikvq+J0RuKuA70qeAmjO8DDDe+YEWwcqM923sF0v/wdJeYBdEPkhyB9gQg
AtPAfeVo6xYC7H73iy9AhhF0bq9d4k1E8DzEgrZ/W29HQhW7rzvd0Mrv6gWPIisESpeEtWnWaQBg
wDX8LjfvzlhC1CyXrCccIspG0irsPPdW+HUh9/TXt9vWShG8+blVnA/OKbKosSBSHCHyovOKYMcR
Ayb32W1mOhzqoYYfQnuyb2SeHVyD+nB/jCcR+jpkbBjdwOgBLpikhqM/d1p91oJsNO3wolSL8XsB
X1W18H8mg//ljLAqEJevh7zoGpupDPhI3YP5/vdkoT/dsfGmi5Ywv6tncIgF2yxGZ1MHz6hc4zaU
vqTCXCdEYVdSDyBcWPbgf4UgMtzMGIAktCze9xNUxEzRfjiusNqJXH3cYxI4er4d86SRZtggoYUp
Ked7wQwHSHB8p75x5EHO1kcWbgHnvWTx6cB3hvgaUNvR0CActaSrDUZ35aV6bcVfsReGfDgMjXfc
Xuy8Y47hckiSSq5pmoW+gCN/pGO3vUtQqM7ORll7V8KyXq+Gl+PqqRJ9FesoCYsHW9/sOw6anyia
RX/r+Z5w7JjM5X1tPrG5lZK+er7cXx8M8INmnBO9h4lfTO3rfBgFDYW4y+YEaTHUQZScb2u2MA/5
faXkOjOI5RkTaUALvVXVdAzVtjsrHU3f5nWlNmS/6Y6PocqoSYJjaYRL5vzyG7eBfIzKK/uMwJ1y
J+ABRcgEsCAEJMj71ZCeLMq3Qq6Cc/Wk4MvOoj9UOfdMf20H/udSaj6VGjPCYcSBTggBk08ib/pM
WDKZQfAS0LHxhUFzU5xP/erjpyFPKcWjW8HRfcgwyHqMvbYLtNrBFPp5TZgo4dFGWLqQAdVpbaTI
SYMMCmqvv4SIE/A5mqL+CuC6FeKwZwyDBTcPA0gmBi7uiIn+DHLDTfaCV15/kd2Ww/1XGYKqUfH2
xRkmF9Ez05jl+Nd+zizsERwsWI16Sl8Q3d5gYc9BzzAIkH9CosmoLDxPWsIZhZ/v6p25+nvC4mOm
5SxInPtn4D9MOrBSdkxxoqHc53GeZw3GAVjad9ymP2Ukz5lqs3KISqiCKDxmnyjsOYcDIGLrbRSa
UZl3Rw0c4TrzIfX6mhxSqL2+6GKD6CoHgbaMpkfcEQu0ItU9S190x68RSnUm75Wfgzu54snZscJl
J2OQkHFizor6SqR99La4TY5RyZe9Cx8//td3T9bR4bm9TE8P6P/NrgiGW0Yw6CgqL1GP7XTCBJlk
W/sS7H+A+G6U9PfEZ/xRHQiDd4ekNCA/fKB+lGfwcrk/5tnxuMG0QWjDNDyV4BTCvAsy/8NGbdN/
+StPZ27+slCsbp2gSgx6uDNB079KzBJrOELynNq659vuwL3PTmL1uCsF3Pkj0qy6gjlYCs6I9wPW
Tyk1/LtQu1ELgCxJdbRqhCSEM8Y++Zf+RjhNzj5ksPXeXxwWcvPtCUthmoA8VCADMX1C5HraKK3G
gMzL+dtYki7oFHynMS5fbYYuFhFiJMojePfRafLzIS6guNLQYQnr3fqlOqF6Qujcrgx70gN/IU0y
8yNo0OMimfoLn4htkjhyft728q1Bi9ixZVcusqQ6UYIiZOWoAaAGPyAEZndKpkQORrQFNe/T1Ya0
WOWTu+Lx5P8dT1iOGQ2Mn8aFT2XVMB7z/2iikdXGRtZJfA9OiYeAkXYjeSOIsgrpP/n+l1FLlmMZ
XjSdeEAJpXF9oLWoVA8uPmEqKco3JZzKwq7lgoqxfqOL6CHiziLzMSBQAfnrwtsbcFXd91YEG3Oz
PghXX5ugaNAht+7G8WZL9J8d+G2KoiOwFL7R8Nyxv0LtTpCkQLIvo3rM+YBa0cdWcsxwo0zZaEYa
QYz1LGBIJV4lFEoYqxt6T+lpHzGDwuDiz67IC8Jxi88vxMXJumLL3YXpy1h426A1av4XlkBcCm/O
doh89Cc68c247mds17YVxBZHPN+E9DJkTI1FLufEN0B4ZUyPRT9yDbZZKawW0M/q7BtZB95hxaKA
jVOtKl5QTlhDvx9FVS/R8iw/M5JEmzT1oBllMpIxFww7RHo/iRnwhIw7wXpqXi5HoGC6Skdta7Jf
6550FWfRO3KIbZ3qcEE2RYoXl7kqZAnyhFpkI21iWokDwK8TsOG8bu9iL5y5YTViKMmlf4VtleRj
23K45NMAEhBbel9gZrwLnWG/zXb6fpgmp2qn21AuNkEKRAwb39XEeP58sux9s4foQfrH4X6iU5DF
30qIXtvUW/JfISMyGUdD86HyfJFZ/AlcAtt2pvd6NaJg7mZ5ymLiMkioh0s591CfJdUMERyJkAhx
iUWKpBVr28qi3w7ipgZcxMOxbiuK1z/3yq8zCDHWkF1FPJi59AeOb9g4BjP4+PBSYJu5nM4l1xUg
lc5tvgdtA+Q6ah9VaxxSgsrC7a9l3CXLrmSOSASAl8cKWXoZgxSxCxLhjKYY2CpNi/d6Po/xUgVF
NzLHtod2EDitUGI7mxvqxLDOulC1/S9Cyf/L/QUx1NW2USOltpTVtfNlTWJiTkGigJ9MfWAxrKMC
yhVu93fEvIGf8B+PTUcI1WOr3aIq1GF/qkV9tRuFvCX9kfgJxawPPu9RxK5/U0DYBlzhOF/rC5Gc
V7zIudJHcfXh+Sfb7TMfU8+ioda/qcsG/EII4+4jGA2NOB7+VFcRuNV8Ucyb1GXtCZp8s4WcHKd6
iQf+SxDb03RecCBTEjZb6/srtnW8GrQLMdEQldhtCxJT5iUu37fo/HNNnMImv3uwNc2nTq4BtnR6
ktGBa3wjahYlT2izwMRsKxFcxHZsrtj1fXKEj0cUt7KziS7qKJwjOV7whopclCusQwTfCL3a8mbA
w9ZokoYJa0l0yxM99pICDlqdHXORUPJOeMDshbTry9oIYb7lpJxcT0c70bceYaikiN4t3QBYcScK
aT3e5isChU65DvJF2GIfmMmScxP0OICWaEtjHM6gJAXoGZ1rNd2y9dMWioObYmKPOiRTz3+IZfTG
JV3GH7rSgh3TdEXz674nXL/UKMAWxXnqWSHjxP4aboXTGrSuAUsX9G8Di2lIu9Wf3aHklaP6R6JR
fvAQi1HNbE9etMTQw8cppFA8XGDV+Owx/gQNUKNSF9oQnVItLRF0lTsWTIABbYpTsRMvA7Q2+mpU
1pzyQHuq2is93dIxuGIMqpUh2Ejg92zGjvO2ggJ6RP9tb+lT2Jt8+b3BNM4/1AwQy+kvSovlbfMD
OXzGgBOzTDIsASuywU3g90vSQL3NlX30Kk4qkKMYhIRYuW1Pacc086pYK3agaqytU6fQUkdNvEPI
mb+FQ4a1N4qbb3xK9LfTB3/csxiQU6OuQ4CWmfc89C70pNoFCcFqRyqR3DDPSs9M5kKdC4CVrydk
eBlfIrHmlzdKmqpm+ZPMR+mCrWDFanG7f6WBfxVc1JOOMdq2XGkxYhWmiS4Y87habkfmpEpzNnMH
0chnKcfHDOEHtr8TeLY+/k9ZvOS0zYklbmm1d7XDwB+d0YzkziQwWj+83/2c754UI4fqVa3+NiDD
6e9QPE2RHCqAQF96BMzzmHnknm3rCbjU1L/ncz9flBtwytTBpea8xKYDK2DedFiYtPhLAo0pQZvc
dme2CtbFtbkIUO5vlii0toDfYW21ssV5T2EYWlWtO1mb18qxTe0Mgnz1GUHwgJs2Cu4BpCRnGIO+
S98G0aP6SZ/dpM5QBArq3SiEirFaQI78LSKzlP+6k+fQ+EFATowJcMkfvQuZwAUH0K3gQfn6dL6u
nigOdhkJnMzjrALYpHuJnHkP6bl38CpjmB85di2XNQhAd4hnJc8OV6YSdufDEofpiwEM7VLlyP3l
VJk8PUhIAbaWY6GD9pUdegGe/w9rTVglbe3QvJFtmAsFnKKduhydlm4wyFv63rMnE0Ug7x3jhjHj
4r251ylWJ2ZJZ/nld4TDhyW4OJdQmA/i6vh+gp9l+pFVFK3Fj2BnzBwZiu+659vzFb1s9gJqGGu3
QeYaZpEaoZx9pyGa2nrdhOj0gzO0jbGhGiROusck1pBQ8DyvZRAcZWbIi94OO/HYF2cN3Ya1RAuE
d0UglHWPj3P4OcWdifMWQtMLHaS8MqqZJnufMMChsv5RXFaOcsjjuxWIYyDnIjYyovo6GlF2ApiZ
NKE5d7RqkJXdQ2FR4RmijCFfOs1Eo01HZpqr7tpLvrQDzKUkhCZSEoE6CQ/mjs8B6q1FrZ7BJFQY
25SYEkJ7HkY4IrNqtDLWIgOHBzB1ifXAX38dYcuTRwrnUnD1H1YsZb7BOdXyR4rMOIiIJpRnN5ub
mcbdeu/XQU6qZewd8LxooJemwaiuqKfpvyQHQPsP07A1S/3FRLByciqbuWbhO0UdIUCSjijnrPhE
0hPUnMiA7UfFJXq0uX5rxlnPB57XuJCloN0bxg+PGTHzHUO3xxzQk+7sB/BSaWKpxLRG/GSy8FNJ
tbEoNR+L6l5mWlm6lfQdfbF/GNp1QpdBIiepI4uO/qdkZyDWIbC5Lam0RQStno6Nt4hgDpKG2vAT
ZEosBLf94k4VheTkpbBnYVxjo3fF1xtBQy5jWVixyhCGfXc62DRuiXpADp/Gc+16V9mo0ZoSgobC
kcwveRg2pfilpgFA4C02V9jWzMwITnbHdOmOnuySvT7YaJcvO2Tgp+IJRX9LKFc0ULYMrrBH5oZv
C60oG5A8D2GYKdkK48Yf8n36z2TAImvfcx4dWs+LDz8YZH0w7lQtnwyvNwreJ/zCF/qY3Dx6nV96
42ehR4iQT2q9tgbRVPpxUDF8s3S6zdIO+HiSoJXtueBOdc831x1rFU1ZV8nRQ0Clt9IdFqlH6G3j
B3pH8rbVwPwCqO2VN0WOVauXva0l2s7jc+byvnSWqWiASDceWypwEUC/2wkKLGVgN3ueeeHPuRyh
DWA5+epsOwKjsGS9V7X2JYLce6fOTFqPFUlCMKluE/YEXb8TZvWjrY44Y9XdA39VAVfSCVkLhnm8
eeDdGwfPcCtuuuPdmzOkwDbMNbnmupQsAuZzpJ2b+tMYIWJ127xcn8v+IFgPt0xVxEQD+okbiQDy
Iey7ponKZ9DWrThDeQ1M5xsOwXAoGiW0rAEy1O8TkaAjLF5/TrWmHfg2voetOoJZDtd8bcRHTJl8
nUyhyMVQI3oUTEEJC1WS6W68SumYMOUbA9hQl2a7+NMUFibpHubyYhcVvjdzso1sNUwLIXxdvJl8
YWM+D8myfwmIEU+kldoBuhcWV5yYheNbNgA+XUnkmcus+HKpCN2CT+R4MfoUSSQn4KMeimsxCIZp
aKXfpKzUexOQRmSWnJ9v0KkUY/sRd66OLvSj8aico2IoyLoXE41FU3TbYpalGTyY+NikJSDBCMdZ
TdW3I4vyMrdetJYocHMWGxT/XLYWZTDM+I9ixpwmeFaZL00RqC+88EOl3D5c/6xFIAQPOBal5ih9
cYevYpY6UTb6sFC64EtYwsSmlKTAsu+dYR/upzlxK22nJnnMwWoBySyZ7ELTixY+VI4HqXiNFbmm
nmacHxykxahPWPbY4pd4HRyRyyiSOvVKJlF97anUsfY/QdCsV2kPcbE3m93WqplWH3HotkgmEnQb
IBefm+RQ/ib6D/zOdVmTbE4FwDeIfXerYncRtZ3JFCV4vt0pcwoJ539ERtrXrxDk5whSLXrrkAxK
063HlG0+kz/sfsvjYVeLuVosICcjgsL2oUg8oXHN6/PhOVX90wPOWgC1kh+8NatxyHAKL5wSljaN
p5NwANGTEcORpN6+84CKMd3ZRqb+7fzX6h9O57jzumwSIBxQ/0EdAW9wUIKuAf3sJnwGQM2s498j
X7QPlDw8qgHwkcEMvkiwEX8H0bSJ5oY1vkZigU9m9SVVh4oLJQUeRUIpX5aQdUXhMnm7H0gRVPJe
uYgHRNmkMSN1Cf3zER9PiJLS3x8xJpA3CYlUfFx8JsKFlXCFBrwOrHfMJFANGad3nbaaVOsOd8yB
M40LRYH/nr0uFITUxFH2kzxb7xe5UQY0W5PGK2UKJ17wOwUheVZroNrvgr3eOoPrrH3K2vTBhXpi
dAaAAWamzSya9wVFWxzrNRgHF4uIexXVi7Uk5+ITbQ5P4oLUb20qzSAgkw0h4ZlQ7JNj8obXarG5
+CmThKBOApFqPEZWddnc29tBXsQGJ17pUbfOdnU30+Ut29dv+j9YBGwqHOtDsAI12PpnOkiyjCRn
qQyX7SVL/HWtlWjyLwuaoadAWYUkwFlsocBogQiYzF+NCsQWgDMKIkHeAn6UQo2Eea5N9ZZhlOQS
V1bcX9447y0Y6S/pZhbqiho78//H3Y0+lGHhtbDYxYFFh7hv19pRmsdJZcCpmFXOju04sT9IjOSg
J54yLh/5gLkHc/+yRPFxFEtvu+xrdh+29CnWO2pqeAjtPQ5+6ij1WnWPs0IWqsFjBnJynXEm6OL7
5shQzUnhIlUDcor0h5nRyBM/hx/wueCpRDP46EkzVkALAHDONZKXTdrii8iFpA49dbGYyh0CVt6J
aF20KS9H8SEM0+IeolimpXmz7S9bzv0Z28TWm2zyZqQMrqOLzG8gJ05dgNduNPL5BunYh2hjLxms
2dS3CimFXzntEo/Q3DQoBgFzTh7hhGrHUZxlwoPTj41pZDGEsITsREkvlnaszmDC49W6aaDZMb/H
r+UB1U1n8Dlfb9lrBq4oq6BD3P77eqPD4PdQ5saI0beEK/lHlrv7UqINnbZ0CFdPo+WYeo+tIjIs
mjPaIGFxK078N/RcC1abp6W1ITmxIO8k63xgZ+nsxTsAZs49RcauOYBC6gVYp5a2DTElmtyFEDaZ
6aDY4QF7N+5Es3xgX1i2wHSYinihIRto0Eepv/ng4Lg5J5aaHPlJGJD/aqFDJbU6j90INpxkixJZ
oRbbsYtsBUrqOeDhoULeAmlJivMc+ljkska31x/trOf37MV+UY2uzYygFD45gntrHfhhs3BZ2jJs
WUkHANecMxIxgFZ5yYNSl9tFoAGI3119txJ3I21nLIKO7VXmOgTs/22M/4eHEM/SD0WHqzXXyStQ
44sK9cKSzwZM3IoGtWf4XRQYrYcPydgfjBO7oumtxESrTpKrt9LVVXMi4KxL8/xs1oV8MNuXcjoJ
cuP2KsDQ9vQFJZ6hYPBE/OqKJcraxR4vyIkFDyNlZeBQZuxfpwr6q0mY8zZd5c5+36BW2rYnNaqS
yQnv+9+50Z8JdyyWFTMpMdmkrpuwmmeYgDxlDnUuex5QNaZKD7YZfIRA3EoiWQ2jUFdECxBlVURP
lwti938Yd1eVFR75wU0t4PvRB9bPtoag3rmbacUJuq+qc5ce2HK7BuuA+T3nMFQCopWaBG5MI0q3
ZYZVhsLQihalimlNBmUIm9UchVwAWBKtXDA1ZTTB8eapAdsFBdQMhLCiO9n9d+N6Bd/cZho3LvX5
SQ7jnE/McPSqr+zsjTgkr0Qqd1bd1YVUj30GPzeiDvjX1n5CwYMj5qGoko1zKpU4rmxIYkv8i9I6
HaEqcIAuMY8qc1NQxbv9ZttswmA+eMnjiy63q0BjYW7XDqd13Nl3qmmLW5vswx/suO2+QqY+nGiO
rg5iToTU5YiB3HY2YfJHSeXhdGq4do56eR2mS6/oAwtPjukRZYShM6NNQhk2YrwVwmj00+30eq23
cn06Ss9uW3iTK5HIIKMLmeulhSTumJEHcJZtiPOiFg7mm269Y+Np0XfbuOgYVEWwOhyc0/9nPac+
QBpUMAwxutClRvSR8eQtrJ8f933saF6FiunlYdyDE9xh3ScWuw67/lRPXUnLxCquGX4LhUf/ui0i
flu3JYZ+eQ==
`protect end_protected
