`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
BC3b5dqHyJFhVFDHEDECN9V/47l7itvil7Rji3bDgu3OWgAx0LSFIdxqwBO2fKY8Y3FtXhHrN1qa
oMQVGI92+draR4YvEWt+xzZMY7nupdkT+kGtaof4l8y8/3srJReOQthnB41ZjNpiWuaQCh9heIR7
OTgY/nL3bZfG4Y7IYqr6Siw8+eRZ4ahkcOZsPwo9bV0sKKgR9KUlSPA/3NoEFLF39alYAsFnh8pn
xRaseWhB3kYHzND95T4pZjI84b2TNwnAKmSADdZIbJTtT8J3NxTotseURexorhoh2vNRoONZjNZ2
DezG7jG2rHlmUqxAtlUaeJGw64Iln23gKn+vSA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="VwdPWHISkesAKbqZuUv/DQYMnVqXJ6H9YraGz0s8wyM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7904)
`protect data_block
kjG/fgNDkkBEYxhGSx+Yj/fP7MpWHlvSdA71LYgUG6M53g3rOOcW31UxPi2pSQeAzg972zfd9B+z
btCsK05N019ay/wWm0MmPw8O+OCQ+m3SZPpXXmi2J8UU1QX2jfekiC3v1z4cku4kQXgx3J0/YvpJ
JZsYfhWngub/6Xw5MlqL/2ro+7SQ9o5te3tvowE7oubFh+oA1bnuzOGmrgx0ita+9BzQf9Myw1IL
qgpMEK9mgb1PToGMywAdPI9oE1dMUYDXLB3jYp59wWX/gZuKF5OL5tzM67IBVDTB05Wy6p+m0BTb
3Av3NJXKlK3gQdepp4way5jDeAfZT/AhKQSfUOiZgtJlZrxXL0/kMKRkkRr6A7xNA02B0hMN9Nxp
DDc7ElXkSEeRrlgepdPvEEs5/pTUDeU7515VrYZyEqzAP6hC72EeUrIjTglU1/cUDLPtNRb7FqqV
HBFVtb5xouSJypIQJTR1Ah9A0U+121q1521oFD1pj3erbMxkTWwPt3jDrSFGS6wyICV7ol0mijrV
zrrfJ4oWUfhtvKoJCCI7ma6bGW65z+8bLko0Imf0MEqhEPtMtv9VKvQHfji82/ULEh6HKPGMj4qB
h2CZYSGPbD4cbbVyOF19K48PhkTQJDqXM28x5vvkoY/TP+pgF4mDDU6WpXVhx2hFrazMKgOhUoWa
FyC4h/7mU1YjhT/TLkUpuDakBBghppZyxHUsGilrDs6IyKIOx2Hnhpf5mAWb/CjGLVKrF3sHqWbf
z+e9fvfjghGfrBRj0Z+ERqNNYV7/+/Xx9uG4W18hu9NEK/CDIPP9sEEhD8UpSbWTj0wTGY17Bz1H
qVtGZ2ao1YtgpIm1KiUiZ+AuS5mIY78+uhNes071Tand5TADGF/GmfvNuhfkh3L6m3WwYadhfuSN
NmHTzUXGEhrP0v2xqkWA9dQW4ULMfu5+q9MD9jXMQeX8cWXg/D8XUl4WCUN+z8uk8s0a4IOXLh/w
yS3sukDj8jUNZd/tFDIiOjSX5V3helhH8yJGDuv/C+1mx7MYs7RruV0sMKbEAxI5KHwSz8sm2Oy2
KqN1nQ+IfzLmxcdfH3yTdUpnORLcnZepLn1m6+RAvLKkZooVtxr/NYHxqhGsY3vvq4FFUyiOZPfi
YJz39iRHFfMTaEF9rn5vWifoty8oz70J3yFxXKDE8mWwr80wFWrrwCb2dZuvdBPhoSmEixlIDyxC
/7O6V+sdlnWl85EKKp8095O+pyGeJtSNXk8ZOIw9apzOO1ch/oVTbb5mPsdpknVf7pFvAHeqjtRs
cwR5qJl6lDxp2HZVjkv2xLiSKLvSBURlSA8LmpgT78lCA+dxfubZzXig5XMuwmso240ZVk9YTKH+
ENeqZ3rf6vOrvbXQzVj74KELHt7H/0OY5VBOVx+rc+hdnwQ6VqOSZYG8oOpW0gfipnKw9FMTsa2Y
j1YtH1+gAHMjHl3YB5QwxmL1uzDD0JvObcVb/CXBKTW2uWg8Y9a2J3xF4Pm5b4B4gOb1raT1/d0E
xDDDetOf2wLbvvvkghS3Ofvm1nVDJDdsroz/1y6I9pN/EtMwmEvFuRoNta+l5S7jWk5NduY5jc+U
BjzbgS0Hj8amiKJM6C+JrOfaETuuGA0UFz8s2GyBCMzU7513mXi2881EAcO0zgb7YKwckfrbE0tY
bSuY6+liTW6MzPs7klD699RTflTUyC5mhzigRX3TdIZiaIU6Ho5D3aoPtCEHVEsb6VpcqqJ0lT1b
Q0Y6ijq5O9bcibRWzkhsmaXZRBfzgI/cnsXuaHZE6yfvjnGxHTdqoFBADYnCmivf4prnw9dtiZLP
dBsdwv89NBQ3pVuYGkmz2y11J7WSkl+bsr/2XJ9RiaGuHYyylpQo6UDkf/mOR0g/D7zpLCeOf0Z2
7mePt72rnZqYoKhhHeF1GwpROzMMGCdd+xsh3wFAjrWAgc7w/Ivpji2AE4o+bJKTGA1V9LPjui4k
rFLttuedwTj39MGWfRmojepBT/WlVP/LsniZ3j7w81sigPM5/VHrvJ7U6jwdzfurampYWF31thvv
TiqmRnjz73IPc9rLIeoD7SMa3h27AWjwPuxBrHVddAsbS/dYZC1lOt5ob5z0F3k3VRN4ICXitpfR
TY+2IZcLOGI0wcUie30qbGBre0yY4Q6MdQQ2eSyCkH7z5u5yZRnR4W140bMkJOuKRuBT1iiWLndm
p9Wqlx2biBZYYwX8C/4ilGcrrtNSS3XtnbfEw23MDWTRRm0JLMT5CXcehhmS3MCFOs1uEVGt9ryg
MzGD87HGfHMqXFFaSDEZ1CLUW+f0brDytXDOsIM3gYW1NwC3UaPtZ1MtCYRNoc35bQClqXuywWAC
hwCUjZVTNmBJxAUGkJ0TzDE3M9r/diZaaTTTxgDSRWJCfpOmUaJw49AVu8zGRC4ZBm2tLdms5Pr7
AB8wv/cXDrOEuWKbe9nXdEutRnNvuHR1EiUpjekeGyT1DXlswfc6X9F/+lEYjZShuzpbic05hX9q
c6Ehr4ADu10EJsvCBjUCQ5o74M8zm8bAggwYRgYiCqExVOASshBvBR4uKQMgDLQ+dWVSZmld39jU
bo8MvnhQlv/zRNgDi+dAh+GPKlwpABDxjgZQPnUFeb2twFRST4Iw645+VNGm9CWDlpfK/nEkudgF
zxCMbvuTi7oveV9hjLtjHpP1/KWBthis/P74wRCdqqj9tnZt8FGI4t4BoYwRMdafWmhT50ucI/Po
2CvjCxicbITUHA1O0LxzFMG12XmRBB4a+Ilg/tRuRShWRdUNxvBlu7wuEjVtkr0y3fiOzjK3e7Hz
uwjQ5q5gw34wT9JdqNHd/i7pIoG4o7f+BZUE+u77+lhA+uyW8QE5Jb7ll5mwKyeQt1IwbqkHmHoG
IzWNxbGksqobTcTAA16kxrdqWbZvPEdPVBC0YmTubQ4BM2riG2kdKlprrNuLdy/8E5SNFcaZNPpf
GSH6NC7QiR73eCQlQ0JxJP7cthQnBFB4OS3iArW6Dr/UY+a3lTkr4a7FnbiuDlViGFdn2Y6JlXdM
/A2grANS7u83ZGH+U7Tde/6eusJEf2mgBw9ShijucHLgEDTMXPrJ1hv03RyuYd5oAT/RbZzvYU5c
Z4s9JCUaIitt6TDkR3EpRXJGTw8REWhcnvKZ2Qh859zqN302//1xtaI+6ifMKCdaNnyuZWCHBG1c
VyUoBKu85KDvGMy+zlYMsgpSXruzcBTXysbfj298mmklgM+3ZvmyBG3jwF2pfN3d7DTjwcL3MeQh
QP/ijU6hDkgvmscjdzcX62RsG60CzkVj33UgzSo8ELnyJ5m/SQTUlS4J8FWb9lm6+phlNba64aHe
Va1MAxDbjvOLpzFvUwqCVnvPIrboI9ZnQdxrVG4pQ4sQWX5nutU37rUvOSY3jyQ+TWMOCkUNAXwS
FAjRIqG1q9z+U4mN6IP6dugpPOQrdlyjB1fl+4LPEwvKwWEo/wGus/Oa5lI5nMa3R0noodXEmJ0t
RzMBT8/KThKagfBOtuUDISXRrOhVPtS4G2k8/w7MBPe8iHCbAmwU0zX1vxUoxXmcbrVWdJscatln
qb6jWSocNmJivfng+F/K4iIroSSbv+UPPUVUnCr9pHXiPf6IX9YTeg9xlhsAde/eBkm1N8jv/BRC
0la6o3e0ouooYHD5mHUZ2bkoZ3o8Hno7VcjUScMKD1JFtViIjyxM7IB9IjOKtyPT6uU30aaNlh7d
3IhRmL6J87xNE9CKXFaXTyd0kuo1A2R00mRo+Ewmh/WIPUBP755noi0iOIhiOFCbhJb/OJuFWzCx
yGBQEQ396XufBwaRMsjyWkv4DC5WVhsF4ibHrJ5ZTIxmNi6wAPj1d18s7ukvc1VtDEZm7InZwKAP
PIvD7vU2G8XdQ3dbEYNvwln/PiYSrFJkpq1YtNxW1SwmxG3+IOmZRRDhdmtUH1mqQycOcflQOe/C
2ZVDEWkZIxZwudjI6a1epo6qrkX6Wxd9I6+whbaGl86GxYCEM7KnCDW1gmXzc1kyrX/TdZ9+bg6Y
W6ViZ17NViTxn5s/VNi80lsS3BhrP7EejxddHlToxO6lxMiyLhusDWB0Ud4r/FCQvqo2MyNimCLk
yHFC+++wfkqTllzLZyAyW1mdo6pu56bO1Sg6pHPEkRRO3KqDq1uCZw67a39mJUVC4sV0Pjrg6jZt
q56NxuNhXcUsM4ApUpQo9ipBMzj4gAT0FEqoclwJt1cqu/OyUkhHWvBmxSSt5xXysl94d5Nwp3XI
BIrgmsn1VZeYSismiQTO+bwrUdEqAVuK23HVguxu9YHvXsm+qCAShBdBNQfjkuIGtrHHYyW1lt3c
ZhnZn+eXGMfnFaqKcrDzm3eDbESguyewZ2z7tpd/ugxYZUVU1dyV0ax1zd7uV0iqxviWT3GfSbtu
VVSfQVMoUcWrd2ucIbSdJHqwTuulsxQNzX0tpXLZRSfE9dh40uUuPQ3ZZpi3iM5/vdpOdLLV+UTn
U42Hgo44zM9NhKKrr+Y/Pu8SpI56L7Wt4u1l7qUhjbhUO6o7UdR3enMLd5cb4517a9GIB+k1aMMY
KiorOsJBzuwy/we3wTRGLahlb4tU9xDXiNy5fsQ4Shs92mvbbE9ksEHh0LEWPignasWPxmhw0j/L
x6iAJNLl7kHpBYki/KYdlkbNjxy35N2pAheOKdcZq6VV8/2wX0Gb2EEM+EHTHIfj9NFRNw+/31Aw
PYRqTPcqlf8DgN8adQhJQCqYbxv9yn6LwFBczGKAXWYRx/UA0FuPMWvEJmDRYoZ0LS9haFTgvNPO
szEJLqVgxDRrkA7F9NaYHh6E1rNH5EKcCoYst+fB08KRhqpVS6z0FxhmvcpBtwWAKT95CZSQK+qL
1HH10PZMD2XYG0m2bD2fl+rsUIz4d3WS1E5xzCH1ejDpL1qtskT4V8mBfOmEQxbKerIEHOXWo7UN
E31RFyggC1ZCsQpMqPatBEMBsjjS2/uOq7bzLHk3hKn1EzE+ROi0bDaTMgmYnJ3Wdz6NfMlhQmtv
JQfrzEViHmec8RLY6J2knMxgxiHPDfhVBXc6l2XYUQzF3QFlabc5r/ALGtSUVOyOFFH3iMXU04Rj
TeVAWTQ8lkYVt52fB4F2xKNpbu0JjZ01LZtrOAW3ffGVjY5dVZb9MYULTf2h6txncucpoWtkLkvJ
0oNq8vvwiqPs5KVBOfiyA/zTYtaUcZmfAU72SDbGKbZiCgZsrAvzASMWQ2ksZpeZQRXoAlPgIoVo
FcFjHdh5bOuXeFv8Fi02ucOpgbvL1FzMEZ7HWTd4+X9Z/DECwe9kft2wI3BIuuwixUhtv2Nm8XMg
lH/5F1ZinejxIivlJexunvspxhLV3tG+fwzlKFB6tW/iZHyGBLWXcqFzqayl6/iOsaLU/+lCET7C
NtIGlt5tWDNr694p9IJZmV1OqkZ7CrR1Wqjseer+sdNxpiAacXbw3bnRt+zcG+AThirZlyeZyD/n
W/Vnf8we3lg827oIRA83o98lEmxAtZLeC3Hb2Y4A5Do+iTpVeHWWN0SWWJQM9ogLYzKjEfUn51/2
sFcLRdN/nptpW4vCuMob35C0W5B6nKFqQLA8TLaEV6lF8foClSwGFsNz/kz8x8GaT8MaHX8c7t3q
DU3KlyDuRfLhvUyDLFAYZ8COKa7Dhahuukow23U+gHRgVY9D2NCzp05QQo5Ftmq6fT+6GBijbi6Y
HCIyhDBhxZWfsDutitTtR9GRvuOJHPkFU91HIOl3wVUXJlWMeRtXgDhdQwKM138YrlWS3KON+2B0
MdBG8rLFzGWArusHKGPNpOXwWqCwELI8TDaNsGkK9/7EfkP3z8RRh+Loh04OpF5+8FX+LjdTkv0j
6tuF6Hg85HpS84ybb+y2h7DUF7QNCICWsTlJeLlX8IxGj8m7ZXxIb1yCALXCISiE3sABGOKBbWgA
Tl5SShYupK1ak/4JWbVTYPGGzjmID+Mtq/zYpgxctqjR8tr6JIGGYY9/SDJN/bQRHY0enTcV+2h7
yMD0Z3aM8K9qn4z7ee0N8iovwE/8vlxnnSIw1nIXw58HsuRx3ggWEjo392sfcPMNUU0Kjs58rkdh
dqysnnQN2Ai29pbdc/+y79u9+qIrkuh9anXiLgDSyD1F6U1kz5+6YEXsR6T6ztRWLeH/4MXb1+Hx
x0DaRNrT2Z9RjLi6NMN7E6rZNc0xDLJ7v/0pIrcdNSKJYxo4cR8MttENHWmc2d39EWBLAXhUhxsY
w1IlAhBUYrJXVrbRS86VmLE3tSHRlFjfK97IgnU6+LAGHcOmAquVgIWesjO9dtBJF+eynNGztWVA
h1uTzxU8JVZ8/UHg/Xi/mnR6u5uBYi/Q1FD7+SawDe1nWDZz2mAIBjVhOYYlOywKWW1yhjDfdme6
e2q8/npKRtUAPdNSJmcp0RLpsnmQnV/8oFhOSxks5udiA6quSWgjEHXvp7pL6Bl2rJvp6eEkXUuS
NVUkZUsmJ3WyPTi3GLPxYX/iDDEOQoTo/jTPUFzznolIgo7NH04Qfx7GvFp1wBQIYIIUaxJgwi27
V5Wtyvvvq+5Nc2rLKKUB8C/Q3VRv1yx3++r0f+HORYMtO7iMhsshXnGK3Ndq1gA3aYYyo91Q6P0m
roOXHz0ZhTfO/xQYj9vaidxmPvlDVxp61gcThdNysorjJMfifkVtPwgq4XO5ZnTaExShSpL4FgDg
tdrUbReX+QEJXOavLQrHkt1WRfcgzJFtqfUtH0Nh8T6fgHLVx/TafJ1Ole9lrpExr18oV46akeRu
TXU8QcscfbiSs2mKiRlbb0jF3LQHT6Ij4rz4xi+sxC6CE1I2HB4NHAmsgoPDPOM2wGedPLKHDUAL
2QMtij2jPqMtA5xTMfNJHUJN0Y+O7doCU7GLafdRjDChxqw0AHO7WC8HA/B6sP8nEqUi7CrrVm9H
FM+xRtq0IojvpW++mHVhMEAHCZ1IIfuIRpiLoLEueNLVEgyOvOpZ2PdsRknmg5iIQW81rPS66i3+
h5HcYJwqbOuLrDc6PSXEESc/6C+XyAj57BT8sqI1+cEPTeD8zRLT8f5YZ0z2FmUATfqnDJ4cx6jp
4cIps9srhvUWVSNbI4SWHiTb+1hkDfpB8Jdm9VSgmLlXJAwx+Dgh1Ra+0jWg+SSKFdvkhEsUZfwl
2ruxj9VjRsxVyXOX8uqYJCj11VWgKEfP+S8tY2LDlCVgKDhmm/LIui7dVHkyBb6/PWt209A81ksq
hPTh5zAYUpCp+FkAfZ0WeoHQemirPphEp351Pjios2UlwDAdJSqP1gd0uTKp3Vapjck7S1Kg4TSF
CAu2RAl7Y3l62Ue+swsGFihDtrHESt0ScK9+gSs/nm3PMqqxr8JUX+HlVVtrq7X+L8QLtwMotK+o
TWPeyzQBK1IIM0n3fzJkfrEcn3ZStnJljI5jhqZkFfcqYMCvl2GGTacGNDXbK0Wi+Xqy3Gyu8xUP
QmcQu3QgM4SOkzXeXtrQgujZjYE70TSp8fIZAZb17OAirs9iSIxzadzrKkUny+F5viVSkKMR7nvS
/wm4i+xPszn/uGBo8Z2WKhPnWeXJfDb2XWzTpmF5zKPIoKKeHK4etE8FCTa54El8LY+R5UlrP8Y4
FDuud9a3JCUowuuPT9HRYkX1pSfHzMuLkXhlZVOFbE4fywl7JpiMd2vVdsNE7vMSVgD225RIIiRz
absWPgXaJqowZnR+IprgZQgVHrFepY+41DpnhPoay01RFSOTY4Votx20KxAHfH1hCsAqdYu35FCN
l/zn8QBOP2RbROx3xQ78294v5nKLqm4jmtEyzOGuYthH49veZbhwKjzpf8Gim4qOgRsVmoHFU/kh
Wydk63emimXFz3Q3zrCVrUU2iz3jJ9MINQT6hDH4mKz7mOd+TPOKLaHGVbi9dbAURAKkTUBdILR1
4UkkDVFDi9Q8Xwghh/kYRm01hZyHS4nEB6bw/k3/eB7py2oBm+SaymT5K+HqOe9l5E47qLencj3z
pP8haoBTkAormWYM7of0cqHyo2y3LvaUWJyBtXpEHI6jk0XyblJQX6dSrFgiQQpGh90SeGrm2Xzx
eHrKJl9uHA73X/M7F7tYLr/AxrPqMasKGRqSCN1c/5XZy3xuvieXQc/+A4wAG0IqvyfQQFnKtgBc
dhH0Ba9RWpzKAch4JapLPeZDTigRPBeb51TJJdmZaFqlRn/qiIjbs/+GaGS0yt4wuI51A7/AbIRk
mNh/ZNLWduYf33/0AHKHl95+QfTGWQQ47fZZyS7CdExzU5z2H6km2lp0aKEQ0DwO0WRZOpq5asUu
W7nlSbLiKx+wh9uo3EzOdkd0TIKsIChZcuaouxuDpMrXYGsqSHU/P5TK/M+bpFAN49i0HOVCy10/
adr9LlOLU4R0qDCnuwpReJ7E77iaK7PRr/ddoBDYofvJ8SZJuqOyqfF4YT/HzSMQYExAzbRzL9R3
+pxwkP5hYQGB2eS7gRkRxpiFOREXUi+lOrPrClCoz3st6DIlzXWQlvRzDfaxJ2NYk6mxW30S6kZG
B/p7DXjdSQNf5O2DBNfci7PWXp4ZHCcZBrGAFzSK1l6UE6/qUFPupvvyP+2R26xuhEbvrZrUkWKE
pzoEnzjfeK7Y530PYYh3t2zUdxvE2We0vupy0WHWpu+y/DGWH7LzJAzH3/ers1YbrqpjFyWs4xNI
PIwLvOh7ab4fRhl3vY5SD1fyOYstNL/UFkJRYh8XovzcQYX+G9wjkJpnYh1o5m0hD+ogpUgWpUO2
v9Rai8cUSVfrwCrd6EDwr5jAX1LVXsoH9Z41udJm1qg3BYT5PvVidhllXiU+gWXAdrPnd7v880QK
BOwvVZvnnUpKwMlVvHdc8Gdin9AIlpwM3tAzVsdWS85M2xd7cRKh5INFvH78ibylsuDi7+nUdqkQ
eVIAzweQSYDDfOoAJ7WVJenIweUnjmsxpMJygwgDl3cqKJ3V/lxl64geN+J+0rImOcsxnn1xOzzT
iBSWhUYbotKmm//LblvOHmMZymleMu0xRI/xvqSVtVDyzfgQYn3k8DRKiE6JyBzW19q6MCgJ3RnG
KVSsj9jL0LHHlb86yQ1jJFXRMuHod2Ik+zgVO+S9yGez+UPolK8hzbDLH145Q/d2DP4fvp2HV499
7DEPxYQMu7ImCQberzb0DbV/qOaTyJqb2hAz+iJaJoOTVyonu8w4gf/yEMFg/CKixGy+EbU7m/pD
6zBjVfgp2NyVEkbeTKCOGjKk71AnRaQc8tgkjAPS0+LavxbW0/3EAqqSkIiv3ell3LvZK6b/gDNK
k1FwSm0kjeCiwgZcn6/mXXI32RcPkJmxybnr0wPlp96I7GLUZgfPgedYPkyflEDlfIDVZ/yPDBs1
TFBBUfA5ETABHwp47hgs1Gd9HhZjpzx3A+ISAfwfthG5H8l8wxm8kp1uj1ejKyDWwYY6qTuW79Qf
os0esrW4Ge+/WbIzzdy9szKmurHbm5vLYj0lCBIB+V1u+Xb3n9YeZa3C02OKVcdooD/dD0oIiKgx
k5+Mhecdbe/Tro5G8zW8GI4XgmctQHVYelyilgnC+aOpqx1dBvhG3sfQw69Rt5WDaUjikz8mmq1A
u/Ssc4ZNEIuasE5aVaj8k8/GNE3ATt0eJypI+FqvDmkw2aThWxlt7iJtdV2M/ZQLz2nnr4W97dSj
8JzbWLv2XapRw2m3BS1gy8TJDivq48vRoq/Pzf1HccUogJ342c5Sf2Od9hjj9yHhwk0MIXMWXeVe
1xqsHD/tudjkpyALGF+pHxKNZ7O/ks6YUNT+HqscRLdu6+ZPvmj6Wmnme8TVpQ+dFPYOWct5sd7H
TQu+GdJsJTOxpPEnGWDmI5R+QWIfwkttT/90XlXPSFRpU0Nytu+X8Ni8AgyKA63HDvHbECSI1Pht
aVJGQRfkOM5E0ISShQ+rTS/9dK5JE9Y0sTt4LkjpGWWfY4GS1+CPiu/xlJPNHn/zZL7qTjg/sn+/
jtYUBHyFAwW2JycAUM9jQaqtERuGzhpnySR2aRIvu07ToQxGea9v1+qS1iOXojYDk5gwpxp/x5rq
a1IQHEP30Vv4vzxV6zetu6UqdGRCqwfaQ4iUjxWRyXDnWYkxSc7P50Xi0evRQ0gaHT3I/LLH4W4v
/xAX6ocRufDrzFR3hjD1CMamKf88v5gDCtU00mhYc2Z/yYfhXu6OcmHLDH+e3ckx6humG9pqRK3Y
sexkF05pcrOUgKLA30+kn8qvkZQT4sIesLN8AW4Yu/XGgux7DmkxW8Zb/K6G6GrRr8b0Qdw51Xef
WvxTE1CaeHVIJcfcWk6nuxn6e70WrOSeDrRAHkqGBWaPCV4nRch9pD5FknmHv00dyMZ2zkiyM30V
De3ciF5zptSiOivsCIv1xa90Akd3cjZTXoElP3e65xvVYDzo9FwDiiI0qm5eqtHrURoqk/mveLiS
ZedIZMB0DNpRa0rUz7w1Qq+lb/TM3P/vw3VZYbW3NPGlRfKKQ9ED08r2mpbHIb2soMynoy+qUv/8
Rn7o6btjAEXRatIbSgR/1+/Zyx9e87dWk6htCb9cdFM8JhL7YbE=
`protect end_protected
