`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Kn3EADPKf/uMquAZFao743Wyu/Y8FF1BoP2ZVsKsniIjDzFKqObH8D3DnHiQdNbMgvqtHKlkk7MS
uv7HWWK/ojjXZ2AFnmv+svgZYgdx/txbzYe3WAgW2b1v89xIDeXMbwKs31z7gnl+pRTE2nzgXkW/
v+l6Q6B54r9Iic5+B+4y1QxOI33QEOj5isUhQqJ6jzj3CjGPJLY/vufcp0jN34xYLw0r31MG+l1u
Ok7/wI7Ayax87xxxjIqCClvpEpMh4A8KvQMXOZIlRuTf2rrdjmikx7brnakQu/C7JDXq6njU/Ojr
B5gyZiqI6kRFcxaW4ow24vq/6y/6ioIO9GcWRA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="zFlZa2TG1Ak95TfnxIv+OVTFB9E4np0aaJJ2XuBnaSs="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9328)
`protect data_block
5yo6E/qhSPlYww+tre+eAFsGgSuy/jZmxrhpoKVS/ZMC4dEVBgsoJ+bNXo40npDjZ1UtLluqs8RG
ad/FCvqFjzFg7TbI1GfXmdy5KDietFgGHFFwjOnr6w4KUy26EgYcCnUZtUp/1XW6ITPgjP6yl9Rw
UIvEwPj7pteSnfMkAOcdEmhHfiWciyon3spRCdod/kvrnn7lbF/UHuzllmAArVXzFmqD0DwXJE8x
NT9v7sqnuJnw9Il2C+FHC4OxIQEGyTQSi1rIFV1zQTnSZNtitVg9/LFPASCRVd6RFVkj2WBmlf4a
ih6f+nZF6k5oH4lEdmtonIoY31ETA2noPvI3m4Qxb5RxUTmrbjnC9WPl3/uxRtSjt5w0OtbrXe1H
/SHxbQLGXeoQ3KU2Ix/2O8TCTUt/EsJDVSEW1RM6U0WPsgA4wZ40nODOcm1nuxoAXztncW3Zqgr+
3ikAIw83cy/5Wemy4rNnqsbNTI1XHuKveL+vMPxTos+d++9Huvu+SSwUlme9tPC7SHcXPdTBnrTi
bO0pfgSRO4kcfsVW1qkq6WtvX8yFEQku6moewDzpmtZaim8lqmwQNys27qI8LtAtYqaA76Wt1r7X
Dwh2E2yty15qsrrpFNp6iky2bFptnd7+bZzGbrLePc+F9We1cbWFizeDNcZUUrh8xB4BM1YnMI37
EArCWYxpA20np0VZgkTXvCSxbcVMDjvj7UxNTJXarHgoJHfGLcGCc4+EaULBrAwc8uToWPLp8bL+
twNzAOSlLLEreFpgV7fjb2txkztm4taj4MT1ROM9P5z0RyIlh66xQFzSBc1AXDGaTKCQuRIxzaZI
j5ZZI01M36fBdlzo83FL0lgDp8To72je1Q+ZcYN1UhLTlI65/7Lr1NGfhvjsPxezGc+0VGrSYgzs
1mDOJM+T5pVKYHrjMGmuX7d0hN+NWhtdw8bbEdN81oG2Q7a478wLhcW4nE1EMJFvAY5luMDq+xdL
/Bojq/bjBv/GNnERhuoHpFgJPEt1x52klz3nQWRw9efyEVuwHI1CPsBByEFS8Avw9zT+qFs9x+en
/wgBgFvVhhYtyxlB/U3BAw4MwO/FKwhsxmJ28ZA1/cZMS61UbMbHo8hNASsVV3VqHiTFHMGpFizD
hFs2pz7xwh7WXyvBiTxU8WnMYviwB3Ei/WaHvf5wZvEgscPIBhO0H6ATDL0D9ntZSbQd6d/hYGEj
QxIRHGqpS5o1XyASeRJRXmo3FGlYTvs0HtULMldhB9rzEttwVocda84Mst71yWt5LF32x4ooZU01
QVoTS1L4HH7lCM/xeXp7PedIhbs0eVSM2HSC0Ldf3WdF8zrGy4O8hUpAeH4xPb/06R3hi537nBRM
EtDl9zaDtzEEiZNhQhI4wOTHNhVv9CyvHE+9iZ2E7xS5+sjpq5EijdyUH9foIVBgyr24WHjgqk0x
GJ7CQ67syBOFkkbBUR5VfmgXYzYWahaD/hjSssxIshDdINta1YNsf932Pp+v0I+cfSXJguVW4BdG
BQrep6RfAxcJ4c0OnReVQotqlLNCWQFOqO8wB8oHRGdhefsYgV6osXvu4YAJttwcA7ThqJdMOOGk
7RSpPI8eYkRjgQCVv7+RMguydkAMmRLb6h/AygS2DpyAdeVbQSHCSGoK5QvWewTandwu/H2uk8Qi
6GXe2lt4qj5C3zM5SoV4JC+UTnp5AQ7uVFSi0uv4zLHL7focmXlam0WEKZM6ZNwJag3BqgJF6Fps
G8ka++jEPlhsxrR+uLnOwJxkLe6GDr70ynQSM32D5QyAPg5s0dQCqs4lkJESpEoBixUlnCgckH8p
7Ha2ZkMlAujYrRBsTkp5AtApdhWtS8VaLZqqYmtK9IPBwwIj6w5XUCxnSyxFfDdRy1AOXU0cmhfD
VHHEIkXb0J+Xb1vhm3/46hnS/bEB048cf8lu2Ff+cUAj874Kx3L09H98WmGQR68IfKIHtyy6PItO
QAuQ9Vekkov7bzuIyiWWFWE2+Za00VCy7ppjoH4JiDVcHLiZMbKxffMekrcS3w6oWlG2SxVhb1US
97iUq001RnwUmg6dnahUvi4mtvaqj4bSCd8EbyTr/wtMGwDALHot3U38IEqEcmbTLUzhReUUFJag
iWrNdC0xiYIm7MKugYXwHV8YZQwKGwV/dIJmFnkf6OHPvtYN4wQZzBos38z2td8Nc43Z2mkIKQAC
kaCMHtVaXwMvaoFKOldig+q5J5cHF49QpTHhIamAMaTC9inrAKLDLYpcwQTzM4DoYIgPyf8LdVU1
GrmrNtEMDX9Tn5kIRR+4qXC4XjnfyACiWshcAvmeFHm1ylB+ZYJbQ0UyyxGbjU05yaXC5SH7JZSp
OApyFRsEt8LqJfG9YV6QkKcJhNe0d4crjFrv2gAj6Ut3Ts5PDxWGktI7ayLfw4B3dVeUfZOwCviL
JBksDSvZ5bFeC6vU6qHjsw7VddkRq+HxxN9VkC+W46/VfLK2GLmjjcGsyzzmtRLlwcsJSGJj7UwO
h0FVKSRrNQc5yY6oi02kvA/eME11GyiqpYBKuW31164o5D09/9SbtkDBJAvG31zAoMEoWuNs7gWH
SfIZlgwplrTBdJ66XsqQnZ/HuO5Clr3g7iZ8lRb7TM6wYrdrAsUI3LSqAkBophuuAxtmc7ElqoMV
oJLZbkFZXih59xdBeMojNgvUMHKa/fTXM1oK4Pc6aMJoqjgTbbGOWwtoYnfJRNo7lNk07ZOxYPD2
pcS1x9jDzC3N4U7c1H/GqLR/9dJFE50gtnViM7P/wfzlwWwmUgt6yjB4DsD08jeoGEHUw0uHinAt
r1rN/Em4GV6uTQm25RPMjVzquqc1KEuDQ5BFxGKxdzOWm9ilP8Gp5dnarm/s1TEgD4aCiZRR9D/Q
raqk9JlGKDu2v1+bAY4uQ/dpbwTBcWEE2n997hYdmru2sX31F8arghrq4MvV6XLcnLYqzX6OjQGr
A/T5UNui/ssOLQYIoUG/2fbH2/eKRXpbwcy0bNbqV/qKF8QlrojcEQx+x45X3K//ydQBpPiQJbaH
D7kEfSVY6PP1Txm8b+lKKhYPOASbRsKwfsTslZVJCQYnOLSeYypEgfnycRejJ5G5lzrxg8CBLXzN
7nWOAiDeQNlxS+jJ5IjfUHraS2zIZDgEclrFPNtlmPH9k6AAbfuh5NzSJT2lKpFRU0VBa5INyzIV
blQfs84sjsotnN8sYOei+BQ+bxJY9KPCI1eBg+FDwsYS0ga2xlNCe+/3jnJt+Pr/HhmJ/GwR4zsC
F7ybcHuymDDJ48U/JtuUxOuGDtbFROO9ljEC7j/lxod9ef98fBnEaB0JPbu0Egdxi+p3VdpCh1uz
ALBop7aNYtQ1hkoEg4E5VRsMPEZV9LBkTzczN9ntd2KH0wkuoh6xGjFOdqcWsWnNm4ESSWeQqP/m
pB4zjPmhikEejULRRJsZJCL2p/z8zo2u3M5p7GcZgeBXati4fq9N6xdlHXvo0wfD4fMvAJ568zWO
t4IGcPv+LXmq13xSpM8ZWnOgIBKTs2DnWS0yN14KfriO0ol4KP59cZ448Zm6Ce8/eFUAec1sb5Hq
ZUt0qQ4yRVyLRgQkviltTP1raEgefy2JQzDAvYoqsRNY3fATooJGSM5+Q3yZDl2SG6RrXOoslzJr
JuBz9FQsBlEOfOetzK0v7S3U9pRQmQhqCLgYRP3Gumz3PWyclAttXqsV0XZcaMWFLRnfm5dPqeO1
H3E5BxGHIe5whBPvueybbrcfs++ATqI9WAGGH6wt0owipbogzdwDl3YL1dNTWS0Uvg50F2ULMeLV
M9FUV+zctSqrd2k40vAstR1O1ccED9N71cjVMlSr69Owa6J1XwnJwNenPVfVdKJJ0wiNfXnxX0Hb
bQVXo3S2rgRC4A34diMMoEFnR9OXXkvZBSojzJWrcjycd2imk3ixtEeAuY/ehL/ljT6WNpoGQMuT
wJhPpV2UGJwR/rB3jjj53AemSrNYS3enYcLmNDw5huedpNY9XKz4CMcHozWYvuInNlmpsSUT3nff
kjQGWTKNKJSogUsj+ZXr+csx7hjlKCuqtp6yUSI0mOOaU7Zha/KioQdIrpF9WEp87mH6mp73oLOW
iSXGwxkmTdiJO458Sw7/XFKE5r1nJ14AOEfYr6J302c1aNvkD22iMcAMINGM5iOzEDpVocBWvPLo
q5iLnJ5dFdLP6w49O9hXDRazQqrsMoAYA9vUlBBLrF/uL1h6dafehL08Qk1FS6/vKIP8+6FyAoVx
p68ytAL8upNQKkwNsVKA7o6NP6eaCMD95IBUOWebOGCDLsyGNh1jvT5fvNSKImbRTh5pqcCAnVwI
oTIbXjKqi5rOp+9MgPbSt2J636NwOqN2kjzk2QJ4ksNk5T44HTkxZ0PzLewrb92v7L2Htlk2KO6j
PTDGxFqm5k6ddSWWvCOHTJtx5mit8i387vlTFGXLOjspJUfz/NqCxD/NvA9+N1s5inMgPPBOArWD
HjJG5lbQQwNhk7oRcu21iJS9ex7yvcsy6oRjEABrolxwSTsVaaTnnnZ0ikmypKSulB5526i5kyCo
sO4oK1+HFbxGdr4KQ925No9IveX6rz3VnZQMCvR7VDJiWaaTIJ1mFo0VjqboXwXZzdnqmaqdvRbM
iunTLuHwJusHtb4NTPf92GdBrJngIismjojQSBTfUD9xNinlBca9ZK8ffUl9VSWm/6B6mWObrR5U
FEC1GYn3ekiS/HUQBY+jzL9VFRXsRYe6Qp4vxWxtWlQY/20mBcn4IV5Qa4c5UslbjwVv7Hch+cvA
P2AsrWm+ajB47VhkSoMBR63dH9npY6uz2H429qIAytR2MGH4Rq8d6Oe8zQx32GsTWPPWl5gcWDWt
9hiDGUsBZlcH20o/aAKP8uD7J3/8NThir6bn39fmaH2BUL1qvmknjZQ1sbPm4gi9YAFkEmtjyegw
N8KYQKpJwBDvaU/cFWRMa8bUrB0LLUSTDlLH6ALgHdYZTVehV4Nff5QN5LvLxWJiheyob7+BDBN9
XKvTm+LvQhA609tJXuabpaEZ0cIsdTiC5qmRXc/rarkBIU2Xq9vtGV1LbJb3iz8Di6bBLe8Jm1Wi
OnWfNIALU1oFCw4Q985BESctU7vmREK7YBoxQQTeXNyQzTXMOxbHJJwsdt4gabAQyOAsYRksDDO0
l5eQkgJcIOSkz+0Ww+NCHyYeyeyqicWYIqFB520T2ASdE2pIKdWRAegrkMI6DrOqlp6g87fDPBPi
982ODtl7aY/NI7rBLSHbXr4j3KSDhtvKcF0siePUQGqxURfwmRb1s9IfbrWJqysbYWAZTXltpCX6
3ElZvsaS477w0Yewno6WjGyWQuZBEKuD//VKtjVJv5S8wB7o3nBFOx/QvtawOH7QYtoUkPMRKrEy
915ez4FY1013Ebg6g3DSdK2sucUTHZQwfKl3XP++/NyzUlrlKRutXJAGb4CHPE0/XfjYA74kIyDQ
JLdTk6nQ9G3o8rqWJdSciciWV2QD7nezqOfKKNB1RKA1C6cWSpkXUkVy6WhHXqcP0KxHkVpqH0DS
tWiykFy11di3uOC+pVop6UBQmQZRTSsQJq800q1JvKxIKAL0qDjThbq96IcPlIp1Z9OBmuPkh/Xz
XhxO74SprXy2TMrw/gWA/MMIG1S5EVZkDN8pkPrqCbzetYEoYPyKm2LCNqOZQnN0CQE03sXko42C
Cozaj8qyYvUJwq7gqpCgztwLm1Yx1KJ0mkk5/HVuKQ4fYUeyJWA9CZZHSEuUnMXegFJxtOtGRAVf
2R73IQC3WroDmIo9e6q/e1wVl3R1SRUg1XxHkfNKg3nG1zE2Qs38dEuu9Xt8lzClYZQ39JdX+8O8
0CjM7R149gp73p0p6yvwT5BRPNYy05tV66U7drnrAD7rK5xFPxKlUu62VxZdKPP33moxCCeG2X8K
6EdPsuXNzhKcVBRHMPn212QGSVNr/A4X919okt6/bNm0iDtMoYeVAXsIlKqkr2D9T1+RJlb+ABDp
//mOENDZfOnQGo7+a6mYOhdaCMCibCqlpWJXnYvDdtFYOKDikqs/HSDgg8HDKbwn2DEK4ZVPchC4
kvoXg+QkkyYVKhrt9TKbBV6zILCbojDORlSZ5oibU7Q26Pq+NHr0grMo/dYz53qX58sWEC5YxJ4y
vGitwph2S84EUtOigmSpm9auFJR/r1QRAbfHOrRFmfFDiQ1qhkNkqWbhlDWgi0S45Xg8dET7wxH2
md5Fs9bRm4jSaNpdTb5/7BAFcfjudvfa7UVQas6IFqco52+VVeqFRFkEWpuoCy1HYortuYOigA/d
STaCws1Y34dqAj9+Qo0g6wu/ftT0lqjhj8VspsRn8WXp32gmG7X9Fj2BbQwGD4rn/TFHWVMJ8ew/
r4qFi5p4e4NdODASdnJAp9zEzcI769NFh7BNcuagjgTfQxMwzfgRtbOgUtGZirGosVmwNsjvcJOx
WyQRKEpwPlnSq9bOntGw4e7MyQQ0RsnBbcbyXuzJOB8itZtYfjijOKier1zI4SLs5DcDimBxuNxY
2yBj7buGyVqbz7FLzgybinTJKbCwgaIF6xsls3BL0UIe0PFdolg1mSrIU3wctZ5011rOmn1Lv4gp
ziDONwEtNgY4gPG8XwmXKXmh09EWf9nsqaCK/71zt1+IMlAr4hQI7qUyeUpBn2EszGdj5jNNuu8w
znvC+LFBp20hTz5+gPJvTcGVXx+H94CQR5+xm3CsRJA2QrRCp8P7XIWzM/L52LXa0IZ6jVANMkwi
oMkY3Fw4h4GGiuMeX0BIuPdkJoKbAK0hscbmcAK+ISri0YXLTcYjEcSEK0FbKJ0RrSlRl6pjTsp1
HkamhWqI8IzBV19zDT6ehxNCsMDGpdfcr1gm7089NoZqV+qHoPcOegTRenxjsDLaA7NmaibA2TVP
pFSpEc1d0LdGKMcbwqxBF0DhHmBv7Nsmyc+uHxMDCWbEoVSM4WgRn8VJVgmxxTEKfnHpMS4bIjvS
N9Ddn9sG+Jm+tUxR58/3scjWOMEO0y9jkAMLHVXQdGZ+fR0722U8hSS2ECKt4tsKxh9kfc+cF3q5
IkFTb5TNMYG/3yGQg6i+znP6oDaSHcjcJ3t09XbE+Er7qo6IQQhSb88IyXIgD/ZgdcQMgpxCnZgj
JY7qQK0DRZ8AIBf963v5RVY1RH0b9M2kqfKFiiUq2B4AKclTIcTLht9eQrkhfOdlaJkLMP72LaKW
Uzt1gcq6WUNpIlgUkIl189aircYtJaLdRbxtZZKAVunh8rI0HrmS5fqRt9jFOoD+AfHXj0TLklCL
DJ9oyMn75BSIEe9BVYo1xcLXSuisBMaTKLS8xcHHAAFYHmYcWlswVHJGyN2oFfqJde8USTwG1573
8kO8mNehWNlxQjsIGZHG30teWMf0AIZQknFpwuv0KE/kf+P1Q5t8aopWLLZkRCd65FgluPrluba5
n5qOOigPmsPnVQCUrZJ0XQL/EGM7wnXHrpRebe2DZgf9aLqdctr9ahpkAcSJKUdkigukdeH3hH2y
vZ11DuCTQJ7xx0cW/uzJn9x+sxp4EiMv6IuhFH/+J3ksBNyJCMaEGbWEeEUC0p01x15E3Vpc4EEb
zWIjibzAif+IETFJ8KPgbNuJprw0+HPeqnnM75QTENIXEbie1y7ji/SJ7XyGzJMDpO3a4e8diFiw
ZC73GJ/XvhCSG5gaGJ6oliqvHjc9ZKO3c1dYXDA2uYjWtNKOpr8BM3YGhYOO+xxRaui4/XiXyphP
kr7K2BXUMAuusSi8zJq89BW8O/0sOtcVy0+8PkstRYFa2gp6kIK/8Wcyagb1X6BwNkqS1K2xSv/6
R17hQxdJ7kten/NgZRf77Y/DIuJ5/a4N5xoquTCld3f9n0zOFkSl7Eo+BE6uAiG9JRFc9yZWb9pC
4K3dpupQjPCVjjNBwvPh/h2UgWs4nuFruF5c3cE3bsHJ0ptElj4eAb4Yudij0bAC9mlCn3c9fLZz
cPHJBdDxcITp5+9Oug6BIV3VQoK1EMjWiSl0UlGilJPi7RiQcMdNGddroC/qhUSH9i5P9HRy1iOy
uaAw+t+UJcHjtad7Zt/IyfspK/XiiJp+3bTO43sLorejS89rfswkWnP63A3dao0mAmbZUlMxNhmd
Jjip5fYX1AvD3YI0hh7TUlf+pgK97Ol43C0AlbRdBgqgSnjrbK8PqQMbsIGgzWpw7UwjUoVPDB9W
hFx8ugFCo0JodBSQcwOqZEqbFDtQKUb482IueUbAfkUKeGMOK3l+TSyv+1YZE/NrVoedhg4cfy4p
J2D3kpAEqO2D3ck/MFY23COhDn9YLKXbAJK52xLkkSYyXxFISgXSCxF/Xu+CvT1Fc+Gm83b1oFmM
+gKYv3BEOXMxV/kXzicTjVAJ2J25/7/1Dfo7L2b8/VRfYHAxkEVKgbPMJrBWFBQLc0xZLAuPpzZM
kdzPEr6bfYzUE6IGYLYbCQoqe6UuE7xR/oU4jKqVve6Bfp1Jqjl3TVg8SZuCrausQh7Kch3SwkP7
5E2zpUm1JXPie5k0VRMOqlCvzOjJlc6xGzYUEAy0AadipHsQv0s/x4ZMTE4lX1dJH2J0AGv+5ja5
B2O/BHY7SzAed8BvDcDSA03Nx6HazVzQxJSnDnt8cbn7iiZCJRXkb4K1bOFo3P0YCAFLmb3qd9UG
/9cRHijOLR2YBlPw3jjdhtwWDeWGvrKmY0jH0a6ER+qMsOcB0aAlYo0Zw+TmjmPT27/ersaG+Cq8
FxSydCv0MyBY9LmXJv23uN5YKaqbAsj42MP4LbcIyNDAEvuuk4POPVeEP3zBBnn72Xa8fIsN/+Uk
9hdZ8PEk7Eie/uIPn6aWgVg4yOv+6NyyAPGyz6Pz7XTEz2bjTh+HpRXRSyzAUZdYNgGVxdJgbKtw
2aCAaGqHgHvYmi1IERPgjpA+p4dAmCGVcwXLCUy0763h+pBj3KlBjOMWpz6AOWhkq58QSSmDZg73
HE3zw42fD+7og69I7e26J9ylz9kwswouAzl2AfgnoJ408WrMjqUTEAMOYDxXTfLJKJlR8KW3HmC+
hIRwwIJirCgm+9Noh6P9/eo1sAOODDS5XP4Uadar8bRqUKQedPF3syie4FgEkCrY6NFaeOzH/6s1
jTWLGTVsT2i2udf6X4EFqc7Jex/fy5qzJqE2oZ+ynhWSK4WvtCNlPlRewdhsDSGUwhJqnqNe8ruw
tulr34dNO7tqMa4tjWDrcstA7SmZWxMgrlVIjW03CdxwFbeDHL3dBJNZl8nsQR/+zShNTEq5YM5R
szoxeY/JFIBl47M+65GfNRKFHvdkrAaVLsNPk1EH/lXONv8+8nbIThnYUOIhOdDXpKgzzDFjnKAT
nK+Mk8PttISy8LmJFj/X100PZjEGZcpggC2sXysDCF9Y66x0cW3g+AFiXPaWn33FJ+PPbex0uEx7
4W570jthyh6ckMH+sczgIxvA2peJOnV/dBKhCWZKKvoUgwVepH1LUV9bwwDW1r5FC7PvY7i2DtK8
fGWHIxBwKD8jvi1JyX3d2qyXfIunZnpef4YAZ4RqIfFWU+Iuln5v0U4A23Fs00BDiR4EfFGU0nul
zEX7cC/uqRAwpVGMXPdHB++2j/sTZgIOLo6ytq9BHUgrW1wvlesqTknfRs486YMATAc2fMeX3V8u
S87CA31ULAtPLTtzb4tV3CpNZsldxCZNB4x3L43sa7QBdWr9p+RcLhwwsjRqR5MYxZs51sQVmuwO
Aaz2BAauh8Uf2MD4CFSpgdmf+sijR2szTH7hMiwyQNSbygQEfCLq0rg36erOOX+3FW1fN30/cupt
VVeIngzeWgRSsgLLuiUubNq4oOCDwzuSeX9H//yVAgFrkEi36RchEgX3QOQKLhoWZRfSQkPF/qCk
e+jckli0JFYHMrDIwMIdJKZ0yfJ2kua+LQkFuPCgjxJJMWU+AuN6PwtOGvFgscbJ90qQAIFHs77F
nEVPM10U33Z9QcyXwEcX2LwrseXTcuH9I4hM9q2qWsqXW+oLu4Q5JeHe0ibIX8BMGQeVLZCbuiM2
sda8YskENTJgAgMHNyy1re43fJnAtwdPVfayFawNhVbdpkl7TAL9M4OUJ4F+AWUcJMFNXzH8LRu0
whR5P7aIxX3B7OTjFLeeVBMZvLK1RiAdOiUrv0MGgdcbUkiPT4RQLmMnVrPBXv9xBm702KKE2DCL
0uIGBVUNlCzem9AtV/nDeoCssCsXmhi/wE3aFn1DYRQrx9RToJUVK7TfFVElpdPfN+GmPzIZ5WwJ
wG0Xie+v6JALcoO23bmd9AfOAmr7BZOuXKbaME8lKsTvnHtfKmi7AEkoLaJQ0IRrj0AlaA+nCgkm
u/3PHQCXWURjmzA8OazOTpzaVREqIzrK+q3qBoeX8vToL9DongJTUS8wwgz90f7C7kyCRfhbeRrt
NtqyA1U8dATNe6lXne09N1iJfQi/0WtMVT68WdAym3r2J5E0VPSplFXpwKEkyI929eDuBwbxQ1ai
IbVfXRYQ7C24LcTX2wLXiDYhtcZPMlO+P9rFmnQe76Ar4tHLfTec9KuGwwm/6KyNoRniELD0lked
3VeCXW4/LFqjZcj3JdH91dxzSoJD6zCw2UKemR/EdDkc/TaaKVa2GdyhKS/V441mT6Er6kfNAEkS
S2gCXnyy4mwrZ+JOBilBQEvijAmX+7ZIYXctcmUbfVg8EFAtTWt8MtmdJVQe/l96f/AIQ1KT/+Ua
OMuxnydFigW3j8ojDCkH6bM1MuC+P87oK+oCKVaO2uSSNJ+dXmyJ2hoJKVkg+iq4F0wRn8nrSzRq
vd+L53KhGmYCypQbpoAuadpStFekWlv4fqHWH0nh7vqJwki1pxGHVUGtp02Z5+ctP+DcLYZLpoxi
WN05rAiqdxygteVouAx5v+xn2DwdyXKCg2W/WX9bjGll5ehBHU+NkYmd1ba1ewbwc56U4CM/tgqB
UsM7jV0Poqcq3NT/28hjN3bjfWJ/2AyugANxENiGwZGKShC3/PdDquPh9j5ksZjELmC+/xPcB402
2T7QLD2uPA+bm1og2aLFt6xrsA3m8YxS5ksfLnuegekcuigJWU2YyfxLflF8KqOaR5+/OUVua/Kb
OTeuW2+xzSegCjQ1+9/yIAx0g+wEWJW1qob67DIBfHV+/8dFfi9yaK9W/lC8Zsq+6APrWGcRO8es
ucXUi12N6NHhL7dShHVHc8Cg5EhDSi8y3E3YSN5w8L9sp+FaJyvbXC6ix2JENX2bvOc+TC0CcnAK
GiLwp/UtqQfqpJV0IlvDIHJJYn47I3n6+Z00Y9w5Ht76GH1/sz8y1QDxL1jqz3DU0AJjZu7wKzk6
pYWOmWsiqVJWAikH2Bn+QnNI43RlmQH1gAmbIB3AYI/9nQmXOneIEIZaAKh9PrErc2GjfpJwH5QF
2CrH7Ed9b749Nlnio/iAqBj2vcr8GbxwCfdi/yNV2tENpS8quNHkgY7Y9sK7PzRxloLZviXUM8fc
FABQLtBYLBI7JY481wGTFZAcWxVpgD8cSFLjoAC4w3rP6qtRDBWgpo5niZYT7ZP/zb7qTlOuVgnl
eyaTxJHyPM9kOHrcxcCe3/5NWiospoNF/TjavxICi5wDjchHeWlsWLwTsR3zOMivSC5gsoomrmJX
g0X54ZomS1TEH/NrIpJW56fg7shEJm9xqE8ILIDCAWXr3iPaUCFyJmogJHcZZI10cCDGmRRqTjSH
nI3NVzvd9522jvi/V2sOEab9D67qs8NVj4Qsv2ObVZ1anIXxUIu657jEIqel+OkjgDOnuWYcBjVa
mH+wDOLDXzFCL73zErnrg7QOAOqrQ41772BnMO3AKshO1uCpKro/QQr8e1ZMgKMqfatZAxAIEMrI
ugyzCUpqdtwEEKvspZTJqerQaPJQ2zug7HvtBJa6BX2dpjYQESzefXn8ARFufLjMf+KSIF1Sn/fP
yrIwqiToruapmcNhjnKe3S3iy6wbctdN6R+QYKCyhW8BIs5pAy2TASDDC+PwsXL3Fe31xdRnfW5V
17Qi/WezSbby5Hn1l5/NHU3kJIxRjQpxWKrSHseKfh4NDsP163PVrjrKq40BtoUDb9IBT5O8PuY9
YBz+njcqtqjtgt6VqX4W8bJ2W65Gx2zKIooEIVmAu4r+C7HANsqCajTd++p7kYtjtlnUb8Kbm59l
QADNfewbZL2BVHpnmQVRAIpbrGsqTO9mQUhpGuGzqUvY1LDNN+vxApHj+i6qOFfD7lhvBxZOKe/Q
Yl40T3d78ikey2h7qPUamhHXMMxtkS4N4Q5DqU/lp6pT8yg495JathDJua0i2lkZzBYaI5rdfylx
/7ERUkmnJlk7CWkAH3MDXNRu9goYOS7akw4uY+uG+24BF6GPRNCIqRRuxVC3/D3mvEEu9sSxianN
DVGmODbZx+uRYZQvu0lty3XS6KnIFU6wsx9NpeQQf0mtsm+SLQ==
`protect end_protected
