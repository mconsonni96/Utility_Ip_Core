`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
iei9cTKbCeyQfb5siJpxatpWsAwe+GGP6fhnatiO97rpJktwCgOwczOpPoFZme3dfmR7W3OH17/j
CA1hjAUysRADK/X4qJSww1Sngi/5DWtbVhU5giEYcKzYjkVQ9F0TgxEg1MP/ACrbKNicZwCqPW9u
FgMxaq4ayxSDZrgnAQc6SO1a35jatmynErvZLcxrtHRhzlN3nCK0ev6ZOVZDAMs9JGhrliDkehBW
lPriKUdxhVN4kIk+olfS9THxO8wW/iEwTksK9mJ/QnzhBrildoCV7kk2hF4sd/0jLqCFkwi8bpB4
Yh8e5z+n1Kgby6VN9aotpKic59jKdPYPjtfTZA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="8XcdugSfoZdsjlmaKYII5pOu1HoaDUwh89E42B4L50I="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 105712)
`protect data_block
VdvlsqkSM1RWDy/RJ8rdZh57fbFrBcXX/7xNNxqSK0oXEntW2uDH9TDq7ovjyB+kJnJBGb4OKjab
Q55zFKW3qX3ohPbswdE59kTBwZE1/duwi8Z8yjTkoP+qECwmWHklfwTpYnLTJgAbSYy4XAZ6cvL1
W6C8fm8v2bAcOXVhxk+DLH6LjsEzYq7Y0OKwoAtA70UCude/TDM4XFySJ7IFQJOaX6U5rh9Pxe96
Xx0UJBdHyxLAiWLyqJv6r0mhCKxff17eCD2HlsiUnl8XNV4J7Dz1OOYFNvDGvnybMsqImNkPYdLJ
b52YJIV5BbzUioMfZ7BFV/s4BruhRMPuRnqi8pXLLyMv4WymrEGD1E5xwCuLMCGCNg1jJRJVhuv9
A3stIYjspL+IQ7d9ec/7jNUD1zfkOCEa0bMVvocxHzYb5ngs975wV0KoUDicKnqht15Ef3SOG0lz
C0VvgncmgCZaYeVsvXyykFzWJNz4rbZqhnF9CUaH1upmS8MuAdNkSjkbpfSO17q6UcvUJNJXpN/g
XVRy+5UWB5dqXt2RhzAha2K8wlbkqSc7XVl0WO90uTDr7HnAw5gCKkp1bKkG6T1ds4D26OmuNjNw
CwcWJi5zqORQ5lXyjB8dCVzX8r61mrN9HoTIf+8eO4mpQvBB5UHVAzamW6SrzC7wzIIBCBEwa86C
exHmXldY/1Jna0MibDmREfb6/3dHR+qBIm+edODW+d2ycmUE0Gm/if4FI2E5KVCGfr5iWQ4QGPvW
nviC5DE5NvqrqDOHB5hsuKLjUw+DAxGXfraxMcLe2hsIE8Y4RlT+l64/vZVrsP7ujxMwhvw6lUCp
eUShIw1lf5Ta9x6+xohsJ6ftnxz/u0OKl/V0ugTMAMkyPtgLmBveDstRQ5h5iJbAQTT7bj+daBnq
1uFY2k9KI8B2xjQ+6ZbvkGcFzV3S8bjvL3yYiTyZIPCfD31IvTdeORxv+6jhST0iYB9JsrQ/7zae
4Id3dVXMFq3ySMl09NOnzyIKZsIk41LO0Kx/CjapFRCBIH0QWxRBHoptDj6g/sc/ZeJJyqAWEaNC
QCiFIbrSNohb7O28FcH/EHBBmkKkc/QgUR7i+fPhUMJahSu7owfHwby/U1TKL5eJ9qW7zdNiqKNj
KEd78eREVmjnMmwGOqdp5GdZ8qvNNyHt5/zcgNaovnSSvb0gjWNmZMNpz/mnpv2buWJhqzs0jGXt
viOqFt8YvmLcfWIBTg5Ix2JYQ6r+6yx+JSkpWq2WDxb/WU+UrgS0pBj6Nm/SzIncJzLvnstmlCZC
8xUrFRvV2/paNKS4t4BmWKcqgGoy+02/1Rem5qdQKizHuT0RdbH7ffUDeO/PU7YSh4YkFSGIF1K6
1wBfppwAlYS/CzZxqVuFYXi0tixydrDgQABCTnFdGl2Bua+HDonUX08UMOeLhxnyMx1WQ2AvumKr
+Z7G+WisVoGXIhgqYEmOQWef2X8KLBywEM0YXBPItczOhEwp2hd5m13dfkmmjX1UWJka/eo3p/bX
SMAvEO8kcwW30KRZGQ0DRPfRSwFxU2DqieHmGaqHlGLKFTX1dNZru3I4ZREcq7/+p7G7bRWOJnwH
nreV3Im2cnIWg6vYss0JIUFNpFmDq9eb/2ZyGH1vUirpY2B7mRy2T8mLRys4L9sWdXS020Un0ygK
GCc6ieJhVI7iSCAonErssFS3kcQ+Asy02RRXViUOsVOH9WQFKygwpnUbM/TalOYXIloBRIn0m7oj
vm/AhbBjAWwzvLrmViFKFwH2/UXNz50VQaGIC0KhSzljoDNCxzEq86T+CcGoRZOxTICgpvbvvEYd
G6JRukocZiCDwrfnnuLMNJRmH8BGPTtTfwUNBaNCLt7Bch2ehGkadJxJ0OQVKU8lkmFWff9OaoVK
SnTPs5nHG2KNe/HffadFoftaj1jjYx4PBrkDP/n0c6GYbNvWBkdw897y0KbLDJAYfeDog0T9lX1o
o/HB6C4pclf4ju0LKYGYhIEc4EotzGSfTtXMkKtZkxU4HcKbswUZvD6qBAto5ZQU+Ow/wLah95MK
Tvsvmapgek/b5tO+7tMsF2dYmS6v83X73gsFev8DBeERQ809NXQgvlbMvh8iV7Qitchq2aFBikH8
V9bX2aE8ivWTUAv6aO2tRh8dIAzljnN/XjGAw0SP7cuLT3tT0piZUnclNyseVWZdR8E5FGEDGJll
OWQzzf67p92KYbxm0qmOv+yd128/tnJmcUlsy5B0cmApTaS4Wd3TpGXVOE7Mf/4LmA88bJImBW06
XyhW0otGWFsFADNKpFLMXefgQy1Z3YRmrbVR+BlQjYl/3pIrbdpfzFyt3PSinrrjADepgDO+zk2k
qsD0fCQl9wvMJWpm/mUhZ4t32Xc0cobBVQYOCDeqaSxUMCK5rZ9p8w+bqEGblH8YxxND+4Mynlk7
VEXxxChznry7391e1PhR5ozf/l9oGusHoOKnXD30UCPwopkWG/x41zehsV/7hgUvV5wHCN5x7Y72
/u2xvaoOjxF274PDmD6Ou8/dpMSbKunmAzBwyPs2Pl3ltRjktwOzPX++y8K+c4ufkZAwqQr14vHE
E7DmJvmVurJHD9S+lzPwaMPQKd/65MEcYkKnmWl14V3FChZj5eXABh/j+ByYwCgcUniKsmLMF1pq
C3Q6vPrTq9HEYPDwBQRSNzWxvPH+T+En97/qIusamtbntv58/ZKbwwI8iWCVh7k7eW4sBQoLOg/E
YRI6OPPhZnt+BxiaDB51FxQL8AOT2zhP1Nd7WycGrjSn+QHTq3aye0dNJ6Xx50ybLT1WJoiPUIQh
jYkWqB7+05bpBssXxb6Z+hK499prxsiuAYIIEMvMAT2kr5sel4FdPW1TTlIQgKipU1L0QqTSOkU2
1oZhFv9tdP8xOR05L9GiQv47BpR93aLYIZ5OtAM1TU6hRnl9KV86wyQoOaDkv0td4zUcVtJA3u5e
W9Je4jGIXVygz+LkYhvuDWSPAc+t2W7AEjoMzUHSduuGaOM98SCsH2nRJgv3qlFHsrBuFG1xWYZ4
u3Bad4QkDGZvfeFTqJeppjiOcYD0zlkEBjjze+4R+5+BwiqBUmiTEOP8Lk5emSN2ZlZjG8kiehmN
Myo23E4F8276qEVq5rltAoDVt3my0PD16o+o5s+Gz0MgiMrlxLgYzeI0p4q6vOrc9cMnXnFxxrmz
+Dzqj1EwcmGBYQwMPcX8oY/oIBYQVxkORpFFQKJR7bcRKY8j18ERnZabZ8oJwlS5SWFGwrCE0lNV
5wIEyYGhWYnpRwXVZ2nmTmCUA0kvCEiFsBCfuILaGhMsA7lzyb+9hRYE9udJanHfmWaseI86mQZR
RNvo5OWcL+33H+Ipsh1T7aIsx1kN3irccFfTw9Dwg/wnnEA4KZ+WWbKJTaW0cTAC0s/blEtwveWG
k1Xl0Y/TPpZ2RYi3Cv6Pc9mrI619ySP/RJuNSFPP0vFxsAL3STwBoOSCt7I97opBeG2pgHYH0Yzj
lx2CKH8Wm3RAwwX5HVoSCA9sTq6pcC3hIGza0fOWIuY58326KGUsMoF6FB72WgBx8lhaz6AmCodh
BCvVF2UT8MW+FSyqO75f7tS+ajMuK+PydyvawqeQhpM/w0EnJrbs8Lu1f4Vr+9dcejKnZp5N/Ig6
eq5/q2YtPs1ZylIoB6hvfIFYyA86GIrdlbsqIlwu7gesQxDoz4YZpHcysaf+ALWuR0yERUWlTDH+
vRZLpq5GLwYLDwL6OO4a4Jov8eFFLSve54RBs529XMDV0s6WyOWcJCMo9p9gbpELo8wV/ZnpTrGe
uns8nVXw1Op4TwYfbQJ6Q328N0Obm1Wparu5WRPmwlim0aBUYUCgGl08ensDEBufB+SXe+IBHJFu
zz+vboI4VY8Z+POFTf+D7zsHpAiJ22Pr0GUDKekrhe4BXb31Yldgv8OsNdGnckTTUrvF0RY+Cxxa
qNdfPD8TIbjX1FHYhBSs2x7s2yOtcNsJ1AFnmEj9aiXAm0bPXXYgtI08xQ9PAHD6MVBJUBnViZoI
5BNG3FUDGkvh2q8rZrdxnc9nboA/aaabcZaWEXlhQQVWny63ZjW0t0/GUWY7BGvxnUC8C79/RGjn
NWjAHnbO6x5s4GXFv/J4sE0vi5t4BZ1IKVet8tsBxOGdV9et9eW1SrQP0gmMNQFCimtvNrAQdfDx
tOaLP1aq37RRacdO3Q1qcNiQ6y5HxPskrz0Ez0mySz80XGjF0//ZYQ4INGTHYKd4QP0R/+V3N6B6
+d6he9dfyxypGCQ9XRKaf1cp6oNM+Ds8CNtKXfbbYnRzPWWefUKJRp4md0kc7VyDRzgtjHpNXmCP
IhC60ZWoiER8N1S+24rILURCPHUJHy+zBHcgyTnb9jCP2xNLvSB58iqw7HfFBnRhxFatTK9UeivT
d5AP0OMpXwBkzU5GyA6zyzznHpPjpuK4kvUaO9nK8NVoIGdetl/5PKi63PaltBLFVjoj7GCTQE9Y
wdC6EuU70yzCuCf7W51EjLRnNM3zz/CtIw9S9GWZAvHNJMTR05R49CwSvVMBvtfiWdjqGkPWn/tm
DNSyWhTeoKwVZFJni8JLTK1tDuqNgNS3nKNELzJyRAnaHrh8lVHxBult+dOKpuR8SOn0k+vwJaZ+
+Zm7y9pnMJtv6jqv7vPqynEXWsD+jXb1IxVAd8jKVOYwM0PttCB73yzYwHgGU2/aZka5qkiJFjFZ
0yv0aLsS7wxh/UYVPtBsPUJZE0sjOuFnRR3gttFI4ABcDpmoMepAfvThNytGldwo01mkUv9mZNJ6
vfFkg7EKWXA5Vd9MoKpi8U3xE0cSjppfvNzHMcpQ/9g46yY8Ua4MxiyIDTFgOFuFHjMZsZjEBMua
88fogVarSyoy8BTNAE/mvQWHS25t0rmC452sQ7NUXbYVXlRRrCKOU1H+xSm8V3u4ht/1DZrVfDbh
UCQHAGXpdLJn1h8Rrztc8/P6GBkFSyBlkf7Y6oJAK4FUGcwNiJ+H3TGKVF3LoPoGSq2Wx0tFHCID
gPW3jib65q7v6QeaQSDLctPP8CIQK1cxEPFvFyPuUVLHOkqjrkXZ/N7RSLNVelEhzpPN9WQGoqx8
YYwiNPPvrh8a63Qu2D/WtPq+mpiNh/k1ELTgoSEira2Uk+IKqLdpSnzAInWPy2IIqi/dsKiAsWyZ
0AlpSF41U0EYIMdpWiOVpRUC6VaIr0tCsO6ubrvlZARzx1jX+XBg10jvt4xwO5K37nbwKrcKkHE2
mnC5Vwl+AUJSr8AgUp/48G32mkYPfzGCeXuh0H2qxMdMXtm9eyJayrkLn7yKbaipLt/JLDs1x+4h
6yOKwnXAL03kPT6HkrpNO5vIFGrPYUftQQ+9TOxm9nA18qkqEVkDGE3rxpu+EoKy9n+6qTUkqtqt
xdLDr0VZscR1RGhUNyu3NR/E1a9c1Nk3n22AOefd+Fpsz5MglwBO/YbrTp7mAKm6l+5bZl7ftHlw
08tCVuANWOhOstq5QlkEeY6yqteDGnpnXbUS+eieUSYpglGQSC1YDUkDArF/CDIihKgi3pa7AAK3
NQwe5tnAREGBaLWfghVWowecGMkGpA20hkLoHQONS2He01TWe9bMAgvlbfflfdQGnL7XopzuYuTG
pSmacLhKmyYEBE10bkJqddOt/dAJ5w86v3JJbK1vvjelgx0VFLunJuvLce+QY3Qxncb2H9wE4DfF
bcfs1zftqg8b+5JrUtnoX5byFpPo1w2uezipSl0VgfYFm6xI23ji8WmvpZfPTZpZiLJUZR1Vk3w2
RzGNxV0SSZwiv5y4QVBrhT1wQzaAmh3fOYRIaXPAZRdAk+0qR7cxcnPEiTEGoNF4oJ00J6KPDP0M
zj+Y8UrCjO18xRYV2s9y9l1XQR5en/h2op6+uScohxQwdiRXLGaj29rJtpqY3GURT4AZULNIOzRC
BB8FMIkuzCeIOmeuPV/XYm11CJntO9FeloJ32kbKUkoVnb+l4qAMls2LkHx0cIV/nZa8Ge3RSM8q
9AGtxq/3MgQydhMlx5+55UXR8z6Rf4iL7m+N/3doA1NKVkfwzmoaILIxTsLrWmXFzoo4EB1/faw2
UMqb6B5BXmIHbSSLZPejSeI+lgsCTNdGQEcMLQDx4/5Yrq94SSBg8aIxUxJv92xY954CcDJpXuRV
NZVM7c8/PgzrrUVz+0lVjNRQ4j7X+kIh1y2sgrFtV4XDzYXkRssK3asZCtqiNXsVTYtjHWI6nvbX
DRNQQrYies4AvInPToaImpgMMFeFwkaIc2IMGa6Na2GpRFJV/8wVTVA/SDRZHvuspUsJZ7y/9qb3
PiwkCcUGSDs23h1pGK8ywXIhrpuAURNcrwsos/JvLZvq+MypXjIevDy1+56A6SB7TzxTP1RcDAJE
9aJXXiSssWmrDOQ99M4TsgWqU8iBSs3r8usuzUievjUHXmdxxFfC12WYjH2LRZ8ijmzZjhwebBL6
n9luTxQMTn+ijZr/c7JkDJUHshO/TPbj6PPiWdomOdXz89gEevUA1aSHzWqGKNQc5KE7lZyOplUW
SafEwyEXkHli95xvKVE2k72xvThXP2qQaOtdkuBN1CCjpBaM+TSKW/imdw7WaDcs04amJZlGePOk
aS+wKS6pqCfwTbLLjM77Z4AiPSIKU0nkckIl4aly3ej0GbUtBjZxIafDePRlugsVUha1NpO+9Iwn
urJb4klKBtZLry1swVu4NKOfUwueH9tyFTlYlhJS4epIcYbZXvFV/olJk7BOlBihyFxa2P5sBxIB
qj+stPVxb8pqJU8fZ1FL6SWM45E5n+6sXrf7iCN1Xe5HXDvxRRUGjhRDOsvq3+2HlY6CAeuN0zrq
Yg/P+OZC44iv1Up7ImxnYXD2XdPVKEtLUXtUqoqrnQ4rIwUF75Tswl3i2T7xXqX4+frxJpAJFVYQ
MKhIkdDOWthUaEWasTd+9OyONnYHz9hKkEIxTqBjW6a6cCuthcCgUXzyYPJds2k5M5BMF24lGCyL
+NwNBh1FVKlOKb8sVDbF9g6A6yaOlm7zlyVGt9Knksejckb6ZiCLV/hLq27d3kFkoXFxNj3qktNo
KqdHLrJlQJ90iM5obr9UsSpGDvnBR+S+vEX6piukC+xZ20HQpHZCDgcYh7w+PJZqHUrZGAt/tQRx
UZiqdweCMTOiQHUuU1HokUGHstOhAWQ1ZWMN6nNRtR9QeQn8jhhg7kwmKYaYWCt0l60dELXsAsD/
xzdhnqMX3YsayGzuxV6K7MZPl2u+x6RWvcGiafCvigowKlE/b0IfiauWFwx+cWWISu1LrUhd4yZ0
3+CngoH+y1QQKTVHn1XBhPvFfJ4IXyorSNS6sZYYu0vHg4Mid8jpIXhrzz+c1sBE88xbGerNtSuT
ICd22+usfIhbkepV3bWsfMdhTSatKXh/9p6Z2SKaQNR5WCNDHc9+eP7XI/FTvNF4ocJ5SDbg9mI8
7s7bq3Zl7MbqP4NvX29UXOLkJCy+LXB1hNMPlqbmhHOi19QuSgSefVVvgUxpuiaVp+S6un7UWB8c
cutw2cAzk+UcYIVY9ufmdjsfu29+le7djHprToliKlyLbZys459XkDSfr18A5i0bW49kM7+Y7Fix
tDpR2I3+mj0a5N/foij8PYuF6a+f/2NJnjUZWkzH9YwitqqL/1uue+mo11J0Nt4ZaOTzRmCJfjed
xoepH8KJmdj7/wA2EOcCBf8hgwnOzIOLY7GzEeioL+cGo2Il94y7auppAKtGw5TlxHp/oABqXZDt
dqC+O0/AerVke2X4MkjAQT35fEbUEqR211aHpUhY+FIiTQOhO6HO3bVE/Wz4aVEU6n4PGF3/uPGr
UrAVSjI1zY9kB//smd0DbhL7BrFIxMU+qDacaLknpEhIoFRHtXiLrA8mDmjHglsUNcZzcUZGpnh6
q18e5HAJhGJhF2jwNdXSLLF/3NSpa/4k3Ir9XaEKNQQJmOljellQCLQ/sSCYJ3dlRfoDMu0dvr44
i+mV49Mvy4+ebOjVKfwU4pNcq2r6adcMmI3p1wVbIkGedCrGeerumLuNw4HpziI7me0VJexOy4qQ
HT3vrh6btIUECllf808qylo68XUlnE0QrbyJKe8lDMN1pJT0PY62CVaIiC0p+bDfTcmIJBWrWtw9
xK5S7+aoNmQoiDfUi6t1KFO5oJRHOsQdfIBeQzhH11fIxgT0D55d+CMq4j+zzLulG0D8IbgFqpYF
UMTHUVlhQxqiaESwUOtRSwtDn/qe9R4MXvd6FapSTEAw+O9bEDJYWN8j3Q85vPGaj6UINPkk6L9w
BtH322vs8J6Erx0CKZvRMul/XPhoylG4/EsfgmaU9swhIQD8RqJUVoQWvExahnumuWh3/oZbF5R+
+0rsVES6LUrYi86yKhpMTnyTFey7MX77I3JYljIo7AKOjR2V5EmUgAhiohcOTE09+3i+xu3//HyY
VpcPzHjPDY4KmmkNFHD8mK6TjCzs044N9VTBgUTdFf/YMTZR3bqMhhOh0RPzt9IcZ9R79zpf6LWb
CH47g9Txfsec5O2anTFuaOE5/GhRblJGcCOX51fD0y5IIihTGWRdySG4f8UhKi9Z9E8rhvqfhlEA
x98xIhONHgp5WURW78NtMPaLadCosLUXPz8WpgV57cKbnhe/EOaib3onkE9sgRrwQ11nJzbWBEhH
pXzHvzMXSdWPmKEmNRF/daxtlPYsYmoCnuKi9BuNgJ84xmEl+/pjfZ71Rz6LOAF44msS00WkD2tB
anHGPPUZ51g1U2eAweucqj2OXdGmEy8QzHK4zqEOlbKNQ9mAqLS40W6bDz5AomIox7z1c/XJLO2W
YPmzqYAFSmvNmNzkpN/aDkuy2NsbHTiAEE5HE8jAM/3ttPFnyheeWIaaOWBHkYIPEZ3bky1QcFWi
goZzgp3tozq3GZb7A7yyOhh5wuMd6JhQnwsp5EWZSHPMZUl0cFvVplkGGT+yiGtQSEtPcjgxjzjB
SE2sG0v9Mi0/oZMCUpo9bMALmb+a8mZFzZpCRqFbRIgYt+ORDjUyRjXOqcYeDAuInw+ix6ph7J1k
sifumBASgtZYsbvMpMjYYzcCv1owLDORf6o+Ofi/ZpQuwH8O0t4wAuNaGBJVzuyGHoDx+7xQQ819
lwMmiOnXBZNIcgZ+/zbHKiHVXxoFJRicmuPlEuTqchWSaKxpZHCan6Ku4XWkK7u7GqsDDE9C2T/z
3FWckFsR3PonqVoL+vVX2Mli23CWrSpWCjn/H4CKosYAAUMdpHfGFaRQ+lPpaejVxkHeK5gm84Sx
tyRmgShYhoT5hgpQC0mD0a8eQm8PMio+KemlH0uEi1g0TZH3TAfowwZJrYiZfrAZLD6LImjrnW8b
y/E/9drD9ZbIXifgiQ4Dhbzodnx7olAS3HS0MZ5cn1y5cabjHseQ4IZSNQGeWruZ3OEb5pVArtvX
FqpuRtz2Lp1DUenM2HFXioshi1hNBq2KDixppHnUite+rqWP1o1FiQgsa0KMH1vdN9lz70qE1+eM
ssOXt1CkhEgnqCgI9cHRlqzrIQ6hiHJ2gisyHHqm/JH3GODoSVdB8aJc99vKBUrQsEaURNeKvShc
2A0Z+5NEjTwdux20y5CEmjThKrJpNtuM7DheGSyNNSuMsGfW2LWsNqDBHurCOlDgFInF+cAfX+k5
GOnmDhZ9/+G+dhIDs24HK4oCtPmL3tz36MXb0fWKBtqD9BO473p3IvFnkRB6RBfCz0F8jBwr5ltk
vsWVgPgEbqLvAotLtoPgqk0yxW1excts3lQQ5/Nlm95Ve2cirzr2nGWGGd85zLLn6Hg5joTgcEe5
JHzyq+1lXzCJVdLnwWCsa4YQIdvAdsj+6UUTBHFnI9MXJHcP5NWcGCQP+bQy6at/cKoE6gbGxjWP
GgYBUg0S+F1fyHRr6wwFVIsU00WAdicMOhcQQDEfqNEearSGnWSFHQYSK9cJ4pCmmA9ov0FwWs8V
Ovpu2p3XoFKJhZXjmNKFGOsOqoWvOFL3U/GWg2eKDwu9WkgUqUG46sBohhVtbk42rGik5xYNduu9
IxgDRooPiOHHgmCuwORDVKV1v2svQRxtQ5QFvk8oWIimuaOQOkaWFXmrC87KVDwGdsXkXmDnbs/E
HUV1Xc0jbUjnUeJecxmveDSgGy8HiWKoLXsyMHMKqKqk8OfCxUZCDK+RzDPVuYPRJavZ4NrCmnLq
U1yKzMiTYhtTRhM8Y39hfaLF037uIhk+XrudVhOJHjwpC8Ymb66wuov02X6K7AoKY1Me/bzr727b
1nx1OhFYhcoY2c94eVnmeP2WXtEZND2WdFwRwRALiZCFy7MjsxHoYj9+dpOWLtSNJldETEUNCDxI
rwJ0QyrBzmvSfRbZvp3uQcT+/vk3sJ5c2BymvfD02rXNa+TdZSvSbavdgLECeMZPaPWfQ3vHtiLn
kfYc+FJJJ24kkLT1RGRAPtpLiM7JcJ/4Oc4xTy6QAYAWVVmRIu+3vxbZf020K+y+XWvCAjO2iHQH
y3eKbXd6X/hkpIy02/qfZwfMYOn6zZkWG7TcKbQdM+rSn5ZRknoMH3J7Xu3qB9Hi0vhJC7/BGoxF
GOCMphGqxNH3E3hy5cusKw2hZMN1pKfVbUBcY0DSPiOJxjyggN1yw2xpaHcLwbhHgrWxjN6RpXEW
6A1c1+ykHUNvIQFcZmQg2sFJjJV8dPMqqLaxZidYDTB/NFrUmaEgfbN+i7SBZI8vtTqVlnDxR/pK
mu5rTWFcJwbY8tJ6qqcZ3SnZ8j99Gz7QlpRr+Yw5CCEi53UmJQ2fEk6Y/3pi0DeRVBLUbT4zFh2k
Ip2auPSlVGYOymzdACRaTNclG3njlfgQss1fulB08YZx5iGAOYnGGxaaGuBxVMy0uOl3YzE0TAsD
ZWqZZ8FJCS/csyvI9V8G/xB1ibZvqoDtzUz9qIqg0Mr7/QHr1tEAbLA3XcLgw5LwMxMwypyjrU5V
+demO8yRaooxawkE/zwzOr0b5HM63m0Esg5P9glkFXJ1gUY1ZOWA3Orm3KH4aDghHdL/96hj0PWO
0TH0RHAIFcp7NwKzPKSTaAMIcIJgDuo3lyi6UY3Hg1V8gdQn6kYpMII6Gszx0P4UpDFoqCL49Z0m
lu/uySbctYOYy3Ajhgiw/gvfatMCChY8gD9Wf955DgbXXxfk3T0e2Xw4NzYZsR+kcnWT3afM9hKu
TCiVjPUMY9b9gHyk0gYTfS8orMU6R45zea+bqVnK1SD+LyoActbASThRFlNuCsdHS4pG6RYvC+Ex
Tlkiem/jTazxU6k3y7th4zaG7Ag6/Wx/SeXw63AkbJt6NSP4AMZyOkneuWphJYK1gkMjhXEFBFDd
anpAOLUHCpx4lMGaz+vJOHzw31p+UNleOyB83uWnIL61IDSw4F84+AaQ1oO/bIqHBz9Y6w5bs+Vo
nQAxnEGr/nhv8hmLUzpX3wKi0ho231BAo7hnXXfJ2qtXaRWjfbcgTIhwQQF5e4TZK36W0yMPQnak
ugiXwrtJbF6yNFBZcUQ8ztnvWlmxmg1BH51309NhD8Wa8I2P6sY8ErZZDSyfTP7sFrQRetwPb1Fb
cAHiQClYrW/LV9NRf3m0otofuZOYfdqZL8B8TGFnINpj9zLrZmFcP9wQJr2oTSQDSQbEuMpk+RQl
rFan7YUrGzaWw+DFQHOfeZUuqFNuV7OWmR7ELXop8oI45p8B0swP8Moml9WLd5ZyU1WrEW5QgOGI
XRElMBCKTc5AYRlucBEmv6jmbmmm4DQscd5wSui4jQeBQ1zcoJstFrFeR1jWNBm5j9xIjGP84swG
Swr/SnH1yRAlg5ibSEceeQh0a1vXzl7+nCncZ5KsBroL0W1y+yqVhTNTYQ4s8Py5Mb26uogTHQ9E
Eik/e+vKJU2WBc1wYjFIOazJoAxSWPddcZLP8WFE+Iv7NM42CLkU2dpVIQL1bwC/dl9BBQmIkZlQ
P0vT0IQm41SJHgW9W4MefwVDsp0RxpZ2Xs5I7gCYeL65pr+dv26QuiiO6nsLFMq29OgMnQyN7D8X
JGQUQwUwx8Fdw8Ez17iQMvyNYaiuJ9HvQzkQs5S9fdeUIH/JNHFZ4nHRVxkDxhXfI59Nt4aSoH1o
MTpHZeFAPKVuRk5qBruwygNp1gU8R1Wy60PL2zEQ4GDgKOm43AqEhUavaYmYiCh6oc+CjTu+MYqB
VFe9LJGtLy9a4enhrPOs7ZgSMjyjvFOQyhy9xg/l+egaQGd1hFyvbK9wPjJi9wNthPhdGuPKAY2W
uo6Ysawqn5Ozu2AGcXq5+gN8kCujpB5LNPz1B+OPrg6bdY4XM3MS4pIr8ag3YYIFRRY+BpjI5LBk
LgWvBJE08XIE/61PqFuFUfuSwjjy4Pk1xYn/LOnOTOuve1O2XZ0QGEwgEseX83tVjJr2xzckM3ib
3WROSeS1BEVLMvEwZncyIeZsPxnyyOY4tZL6HjNoCrmbaDs1bF51xudzwLtwCpbQK9Sygr1IEyrJ
b49xuXkTCxSSqbNYRt/BHHuRw8gVzftVL7XU5naEoOvWrd2w5CHMLHYy4qzwpmwziobjXaI4yTmJ
jK2EKxYTkdUj017mwmlhb4sMjmCgDAfExUgMfnySvAIWP+CSOWq4fQV7gGSZz7Bj44fj8+48FGsV
yhZzz/9R1X2FRhcD4omyCy2KOLY/yHAzM4BHFLZoge3REzCn12J0y7zP7uLNRN1wymGwb3+c8d13
pxEmGjfQs9brGu+K1FimKSp5qIh+AqkjmCVYeKbgRwXz2WfYfbUYr5XiHBPU/wYYIuSTXLkrKYA4
xKdx9xYxEmsOmAeL4kBLbErL602mnh6gBXMCmQNqxad8iZZA9fx2Plql0+NBQzf58l8al7UkGMUf
YmA5WmZCNHhgNc08h4MADa/JUu57jKJvUvPh/W625xV9ADAImR/XwTl2Yi4oZHYKmfpeS1aa0SnX
SOmRJ8NqIoIshjfVi0eiimTSPAArylkPj+RMgNOV4fl3OLOmfCEAtuOugsavzaRforazFGfUWCPq
PIJm6oFrJ8o8QWjl5e64ifigouMM/EW8yrWj9zSpT49mZ0kyTkOFjUuoqsXII7VpzGCai52o9Gdu
K8sC3poVBSxf9XPeYcx2Vemm5e14s2bONDqFYTshN2uZK7AY58wHd+AqRboRKU2amSKBSPWz+QiH
xFIa527AA1QtAakyL1AmQGe38emVba+aY2XWbIyKIS7emQhkZ5eVOuSVISwh4aZuVDECN0AqukhI
lsbi/aT/SPM+xfYNite3UJj5CHOz0xEHn4M1UvMK14HO+fol+0V2aZLADVFtQeWR39TUMLJYP5po
3AMl+apY+G28OwSLWBaG7xxejVjaSoEzkmqCfNJcFJxr86lYS1xbRpzNsZGGX4fHShc+cur4bIBr
eZI/FxQzLHpsqM5k7v7JOkhGNhez00ln/9L9rdw/c9YpnvpXkvyLz4nfvzqscmw5+uwWtV7xv0Ro
2FyQQdIMG2sL3dSgk8/qPJ3x9QRVtidvX4/LMXUr9bIg6fe3qQauHtAqqSfZ3OdCLnbxX/M/rh3e
c3XRq45O8530EHIVp1HVqq4ZtlLS5SafZinJVcA8wxt0hJANWRrf6GunibVNJKJTQM8AKIzoNrut
4Zl54CAF5U2hFuHsCy4zH5VELvJ1B0J9jpI4PL2If1O3LoAv9VFfj4q55RF/p8onvrzw83LzWLCB
O1ND+8/uoE819JpjlpJQWedzoPfVqiK+/1IFTNtrpq107bWsX8QnL5G9aj1zukEwlyVMQSTyHWMP
nXVaaBpgQJZTPczded7m+iechAMjiGFj6QaZ6hehwuZjqIPepnHufU3eQjWVa+Foa2rA7wR7M4et
saMbyS4moyxNM0QD/cOuZWr9hGL3n5EXZtJjIE5AZQGiJsavfiA6QV0gMIYAuBGHr5t9Y3JoKJjE
5eVai3+8eGSalbK7514x/nL1Is2OtWhu/cdbaPZ+0ErXxVFsuWBNlJeW0vreXEDd+bKDO7t+nC+f
YRMLIzofPWrCu03bwnD9oEmJdcvvWuAmuYrZQrWcb0zrCyXyFrtletFj2I6sBOj4+F61Y+c9utSi
wKNhmf3tx8zqP81Xh2tglT6V0zOCnJGQUt1RmGmB98DqqgLlbrxPl9t3iEO1xtsPFR54MEs1fE4f
eES2h82XcoemvqOsaWh+iruPRwPHG25ab1/FNF8xgi7lDhgqm6fOa68rIgjOQfeS3nZyCPdG9nPI
2mZF3n0OBQGibm3ZWwUaglwrzpkRENx99iChT9xmrOo93tRPV6ba/z/fyjwoiqPE6JIR/UejPRmG
wghp1K4nHmVQLzBMPCXhA6LIbqEru6QefLsNlXbfr7osKDFhvzGxHditsXRTAJFug6NMt/R8qvqK
UaxNUm2P3fHPNm2B/YX/aL6gD3r+usKtiwx8lamp0T0cGJxJ6YGz99Cuqy6UAJE9Sl9QJKeG1+VC
no734WDik973tFOQefU9nqpnF6qMKm5Pntij2Z6KvsGfu8ARQu7StKAxolfcinpVrBFztWVP1tq/
Cyu0SV054aXpEvtRTONJ2jXUqvv3SbJYqahdMivCKFmRHhtoXsNG8M1OrIfbSIKuK1WMX4UnL0Ba
BIligNxrudrGjIdkAwM3XqeKkJRJzyTbn5oqlXdM/ctQZt4vG8km/hSpEW8VJgDhSHjHH+MgTBaQ
swh6MtuXGM0+A9rdTzQgWbkWpqP1asHpb9sl1gfE2+5Y6Gro2VQd4YSrF5Yid71vrBIUYZIWfQLu
c3zkPw9pXDknC54/zs8c50EHRqfM1qBf9eB8BjTecbWku2DRnOvfrljvCLJj224rWRJlKEG8aXed
fcR1OCQF9BHGZP/IXMcFZDff28a+90IB3IqJyeViBfqGl0gTIA97yn6ItKD3ZYZqI6GmpCH+bFXr
bnrYunv5rm9VlsskLRb77eKL14qUlwiZGN5M5QCx7ndPqAEhwcNR3LAewAWyy65zd9WfVL0QdVRq
iJbWN1KK+DfexEvY9cJUTdz1f37qP2fTIb8a7GZiyTSMIztaCy4WsXD+xeViC/qOsVnzCwJ99rkF
cl3iTjWEtfmAqb59xeHI6zlt1+o5Yu64g/CZpFGbegjDEusAOXLb1ydylYm0VSIbheaKzSLZxvzY
XpyIQJvuKVGhXZ+9dc7jKqDMvIESjg0pHwVTkaKL+n+l39MLfA80vOhUVtSdzPMk/jLFRgtBnLeX
uqNbn2vCngmIfzBDhI9sDsj31TeR2W0kDEuwmzSB2OpKfU6n/BahcoUty6BMJxQtuxWN+jBhrn0+
k+zj/HUPK465JRAm007JM827JlxKF/vc/kqYoWx/6Rlkz70OcDz3FEySNo3PftyhDHDpZ0+CuBYU
JpWGtV2QiBxnQj7seVF11CwGyfGr3p9WJik0n7QFbWw4YKQN5EKnu7halNmaaX3ZWN/lPYrw+Pkq
UX/QP/SJWBDSjQsBuUVZ/x+8fz2henWkUE3vMKjsu8qIJfEhTSPciFW/JymemAxI8C07ZO3AkWZ+
N1xmS9zkpBhROUlF/kesD7dk0n7dfh+Hf0pLIgQyUztNt7vY5KOCn2+So2Yf9bhO/Q87lWnevUkt
RFRni7HwHoVulh//R1wh5eyHCkctsLqkuRBmL0o1NyHV+l6NnG+/DNHls3D07xfmSSBTj449R/ce
j3/7AkYHd8Q/rf2lYxsaDQNnDSK88Y2xsuOM4brCOe/bg144+oIgziUs0ayj4XTs/Uj5gaHr3X1O
Tr7pq9BMHwl0Mirg/p4Bbx//4Six7JlwpCfRdGQC51x0kb1Co/yLKO90wzZLh7ogk3FqxBXLnLMJ
5iwYZbmO+/d1Ou4VD8Whn3W4YC1knVznLsM2BETtNvS8yGtY0gYAI3N7QE/7pytsfRVQPYgPsJan
3wL22MF0sDuvfjfRlFoP0LaObEF1AI2G/1CsLicblFmJ8BY/n16kExzobs21xNu9fGYS230i+UzL
k5IRWcy2oFv7dgsqmfLdnlG7vaKJU6cWfXQ4kWhFcr1GHutM2iGoj/BrZkWf8xopMn0dINN+Q/iE
enmd6V1PYfu6rqIExbMpuU0q94TjlZHfoFk48wM4wmGKoXrDinlUmKpZQchcmQYxPq518lOSwM0a
7PwRRRQsXDT+zvRuFp3ab9nGltJLRPsmaBeQfpUDz1c9C+fG6v6tTYBYDZNbW1joKG+/brKO3AIr
C5lqTiSQdbSixviWi/UmGdfHBjml4ii6MvEvw/1LsvPAJ+RwbA3mNxaaknE9ToMp9NfceWjEUGlI
RaxJmUv8cv0C5v2IIP56xN6h6gePhrghpB6RstCDIHkMK2YyofFmb2/vlptWkkrRrWQduX6knfqN
oW4QJaN5+tTHLiSKXc9LrVSkWQzYBGEkJVAqR0T93PnZ70kdk048JdT4MnJJU3R+TTO08yND96H+
eDKsiqTiiHj2Tby01E3M08HL/UTWEeA8zxNGy6Yy8PmcGl/xF6KhlPEI4e24N0Q/7wOJIjLX7YxL
/Sq+bSRk7oPq1Q5ImF7ltrTnHv0uzwzNAt8fwYvPCbwe30Tku0n6XLWCQLUHuQn7Cz5nvH/q6W3e
sC4PWHI1ZllrjJgE+rMYPSptWU3j0Xs2y/qzksluea7Ly7UlMA7cQLzl1uLuZE6gm6kNRpPcHumL
mcVgVK7OEKYgRF3WdHnAxDd/6w+RTp7LysTOvHwlUG1zUHJmShOGaBdfJHhSKuIhBufcbc+Gem6+
q2+/39SM9HIv4B5F4KpFxU7EOcE6KgAYMpNH4XGWfsLo0N4Mf24090jdnhOORN90tKLjb7EIwOgd
oX7Imv3WleH8dyjRhJBrXTkMEMgRqwOBnRX6W6vGaVmagjJ0Z0Puik+9eNW7CGsgkZiJ5DA3e6EQ
2iPMMXZ94D3fkbExfKqXySvwYbDqyYB+tu4XRwrSkzfTUsYqT4ikyTV9RbaPYRrC9RqadPLGQY1X
mIBQdDxOlxMxnP/2h+15mEqmRr/B4vDWBdZ0eTnA/KD5l6gULPuSXPVoxQd0WptZHhDjjIOKwZK7
7ZhCT8Cg8jhcevLNJXQxrPB2wLzdqbOprRbItSy4xfcGNKiCLVqYfxjT5ntSpw4Opgx1YcZ926C1
nx+jHL69js9Kfz0L1eQTZo2Mp34bebyKYapBvuNkr4jV8I/xN7Rv8KkwCw5q6GW2QZcSRDxxUEn3
9bXas7sIFFZAFz9SXPH9E0K84VXTUVm5IOZMxr1Du4BArZHQaSsEXnPB5Bb/3ywPpy2lDXO2Ja5q
g/VwpRyNKA8pzkkaZRIUttjIlfooD0LpCi2ShmzIqfXGuQUwkSzPYp4ml9Z7aUis75EMqZWg1USf
IvDgDqGPUk+uKNNj1I3ri3TcwRNNzYkTiiqG6Lb/l7JhjmL1xcQ9BUVrgvwvNNQ0EKumSJuFeTjL
6EhXHnVg+2Yizip7lpYYuNgRemQ/R0FCy6eC/8RfXy7W4WWOWDhgJijB7o05NGnRJmiS6RQVOurD
seifzbYVmewiO4jSFeDhA7NpBvtZx5S6HIAA6nsxs0sY6k2iXFEYqXGINOQyLX5Q+xBpY1VuryTY
CMQcAgVNKfB9KyOyTtYp4tidS5Bo85gkSXDZ+Epz9r3oNlXn2Rwt7iOMDbHRwW1I891tTSelNC+R
5ADn7j23ETIgYkoNvXXKx77ZQKH5nfLHjYZTxFJxWONTZwCnDoRbX1Nqj92MC8iHcC93O5hCj6bT
OXrjpTYKdge0ImrgabcePTTLnRy/tgEX1CNsXmgJLu8FUQAXQJaoeAiZLNAjS6iIeFDCs/ssDUKy
zdZkWieIqLz70rPXDNW30or8wEKPlLk3JpDutPPaJnFgPIYhhHvyFHUrcVWqvqcsvRPdj8x4uX3t
9HZaBkpfoPxPHaQ+V09T2/8W9THkHcDb4Ae7x6Nf9Ur0Fkj90VgvKXyU1BOQ921tCIkPuW1ElyD3
8zqFNoWX3EETDkgdFanBA3JNWwQDr9IU8atzX3OLuP/ImzkpGF1V2BtMbYm839KGtfo5LrlZgIWh
jeTZyUqBSVB3sWHA9gM8VcyVpTeDj0ZoHd1dk3gtSsL2IKc3iuX3zM1IWtE5xutdOdipz7mqe1DJ
bAEjLDwAF9o4fGBZ5L/05TIMJuSKwCHkYnE6WcQwhBvCC7IRanLAkGmfXedgu76/hn/9T2nnCLkZ
Gi3ACDeIDKJwdzpDJFUYkiHVGlAD5pUAmh570EOudCk51mwfonVpgRmm95zZ55iUsrqsP02tr+/U
02Mu9D7Q/+RmxmSHelnmCer08M9n6qygmzsDTD+gJeCu7SVIKCnVP304qZvo4KKkqQrpB5STgYV9
ygM7WFD52FTJU6FuRw7JAj4l14Uv1sH+iEHx70g45LlnWk6itDNhcPofRp6n7eHI/TPNOyG+OijS
HrfpsTjaKmDFpcdbTXENG768ieiHeTOvAZtUvRMhav81hpDHXUI+oenIn6uk5mNHD+qn7zq8X7VM
Wp2cW0SErCn+0MaYffiIhU71zKs4NaeoF8NZWqGhF4O9mZut12k4hN+Uw2waBDioqisZl0ma4SBe
G658MdtDh1w6fSzKNtIT4QP8LGg66OVRv0uqZGTq9gzekIujmIO/9yciVbVTKRb3Hcbdsv4iQ43B
8bSDaw8D8pqDN9J/ZA0uTWhnkG1Q7KpjkbRXo3tieVUiGTtydULcZa9Sjf2XOLgUr82yijgwKLKp
I9U8yN/0ugB9Vj25R8hP8p+lZCoZP3HWQpimcKirSK4QKwT/lg9iRA2m8D4Zuwlr+s5Hndi4Z8lU
kSkCq49IXaZGPWt/yGw9IvJTBNelqcmjdrArCpBwPO6gfZ+sG/JGGx/7UDNJCMDvl4Y8vmQ0OzlH
um8ZmIS9xEZ0hoyNjFFti3PDDx5TQF6gsYHuxZALNyYgsl920Nzt/IVPav8qZRyWXri4H+9n2TsZ
w1SZ8qX45QYPN5juH9/bPRpEgnEdcVidaqIxOaxE+pnL+MUYdTDpAQ5UWqLo3ECUzOY/G+M2zfzt
0u5L1kCuE9BTVwctu631jf/WLeP/NFRKu9AxQheNWvM/WcLMKlTgxpLFf0Ox6Z1q/ePQ96OCVJa4
Y7twiwhowV/YbYXCFACOehFXZI8MG4fL1GCIWBbA6kQKviqpUzdxI9G2qKecSNrXZwA4QAYYLzp6
mr9cRrXYPypjbu3u3kydsixL+9S4IU0ni8ItfWE1lDEKJu7aXSCFj7nV/fc9PTzk3xaOGlKqTxpP
JqY6Wu1V+NmEHX9OqETTbZvBgivwjJEVGwdbQHTKWWeOkx305W9txozytn6xDC94i+C3VkDO9ld6
q31EFtyHV4VA9Yqry00OV4hQ8c5nZ5DzunbZcTYusJOUA5yS6/6xHkt0+zBB+PiOZ4f2x1aLZteb
k1TReC5S6jedLTdKwhKVsW9lTI41Ne8rBKs2WNkWHaJqMChaZyO9MkFwp9XlaH6yLIL1WRQ6Ikm8
yET6ef6ru61Vt5mBMVO2jpcp5cLYwEx3o+RuYyAvPvH6oSGYyPLcxeN3BmpTmzFgMoUsQmtrVRdw
48aNxQgIu13yuLkwfIM0fr1vBf83P4jmhMRkWWxXE8SY2PxbEtur7HTmL8Mni+TPNn5DuxGUK307
Q3IYRLZdfje4hGqBqMpvTKkDy91d99LgC8UNswWowGAwiq1xYgRRo5AdwLIZeC8HAY33Vtt4VMKs
LIWISeLSWS0Zv/ki0/q3/Lcv+zC2GuYrinCNKwxJ4VQ3Ack2kwRe2ZEJO7FlEBuMQqSYM9BtEsPr
StEDpkfLnf/RgthoRDpnAtFCCnOmKnO+5tY5hlovPn0SWo3KS83CL5jUX0abUx8C7hGpjSHOIWKt
vMhJQVHtF/flNDkCa9RUKflFFArPlE0JpMQXIZrWQeGYAW+vIRQ4qw/83Mj/bjJRkeSwmd8pl7gR
ikBJhgVofh9OdfSDLmvDoNcAsgcZU9NgEK1G+3F3VJmtlF9LXiMPEwwyuDvddgR64WMtjnsfBxth
gFF7RTOcrEFuakgBoX2zgmlG4de6lUNguNAWZ1bbDh/mmTVSoHKlFUeJHIs5f+AMhaGkKFiQP46C
o0QTy1Sqb6MQ7pZ+KCPF4XIJpKZrR2f9UFc+AD4XnYBoh9+6BlwGt1ZbZVBmfnGzfBjhB3bxksue
tj8DTiOfUymmtl/Ge8oOCZvifWZ976GYsyHkf5lUymE4cP+bV8q5ZVvdjjeu33QI7IyrAGWVn0PO
UnCeiHGxOnv0xCvqsLibG+WhYchk6lCRJhNRUkm+UImoYGbH3PjpWLdJinVwboD/jcJMj6HbiBPR
iOXt9ladnCHaLDyk/6hifRgzjNIdGWmJeTCKOVxZf1pBb4QdYxPCqs4pxSzX3iZL4rUku4id7rU2
8aMWZtZhJB74pLh1Thj1vaSKZIy8PxpNt7ocL/0zBwWsbl3u6Ubs18QDBNrAhUkktppwpgp9M0zj
NKxF3v/u7T6u9Orp4YwlQs5ge9ie3Nmp+LwO+LIWNPbN59oKwWt1FKJ98hb4B+zf684E+13bcvZO
Ydy2d+4ameFJKySxcqPtq0hz2/YoNpjSPLmraivWdM0J0jkKi4eLAbAds4NN10cHdi/CynbB+2Cr
OzAJG2Hdi4xa3zq0et2eDs71RztS6K351cUwhpHCUQuRTxAarXfxQpV7rIEQ9zgxBf7ZsEnrJJyB
bgtTiZ9hqe8T/dbQHO7Ff7ZmDxR6E7VoZvroayN7xdTELX/e7IMR/0YXlrU8JdqMcKnegBtWsO/V
dZpfzIe0YjN4Z2InPpebq5o4WC20tvpGjqMgG0uPkRqUKXROIE+iZy2f55cn9QdRLiXzC9R6qBdV
jJHPYWriUftE/58KlxSFzekqH+/ZJVwc50Gu1L1kLF4TSb3dyj04+fblAkMwpjSunUOm/dxEBBra
UtZIZapMrBmjyx4mix04QayY1viaxEGbY/tdtKnwjUkup1h7q3vvgAe2Tmk53u56rkyL5SwiwId1
tKdsSMXDYuPbeRvCrR1XPFUEVe38D5LdY+A0Oas2yI8mSs1csRK4nwhAybIwYFwCF1ApEVeUORjB
EOfBawSkKsHW5l2tYztY85sk/9DwxBLBOC5dtuXbDjGBeipiKRBncm5OGG/hXtCVw3wWLAwNfokz
AWpPRly6YTV7Jp7UhY+dY6hfyWyPz5PxDpYiAt+ijMmrqpIl+kLxGudKvqccK+5G2RsvlmK6BZO0
QbvVpnqpfP7OzjhuDlg3jLBQL53PiNBexkY7Yl3ROuJvMx0nEOX6qhjhP0j8qyGvRbVjcXtOhtOg
PJI0F0jIwcjN4Amj3QYz4LwOsucR24x6tkQ6iSBG4jKIVkiZi0WppGMthVrKufnNnhhW0IAWg0rZ
nnfILwWdk9btNRYIqdu/LAnhYvVYIKfMMP0GU9I5ls3T6YtXeEb3kyWDvfoCUKUTJLWKvERXdiUI
BxD47x4dY0I/1YkKfD/zGJlEnlcvxEQk1aGnv8uJMCvTIFl0wfrEiW5Rs6KVHnlspbWydinoCAhd
r0QMH3XlxrIpAr/RI+n27WfO9OlxRgcWJ8zwixrnQB8uuGbFUwe0WY8ZraNVu2OB3vlinJqW6PUj
RNeRzpLX+CYQY15AhEsI1dqqJbGcMeHZaUHmgaIVvqxXiiXJZpTlqiD/U0T26jDCWsA0MXQvdR5w
RJLloji30Ep2+TEvHrYkTiLBNb1NUmwwFUM5SBsNFuk2zjiFREmGrNumVE4spMwN25haGM7cil2a
X4SG2SgGfwck/4gMl2DWTzPF7nqQ9bfhAbaPmU6AIJn3Hi4K8t8ExIMLdXJzz+iaD1wHDIZo15gm
Mb6DPx5gvteaKA0hz14AvQ2jgf13igPjM091r8CwtL3XS39th8E1KUK4Ya7wGKf4cwKpZuDKXgw/
n9i3ha1ZaAuepgsK9ZYPn/CzeAY53Un8J1C6T/KbJP1UG97+WhDAG6lMFgzzy1KP/5wYra7Ex8Ho
K1rqLV+34TdP85whhK96NKQ3tRJQRKLDgi3t95kco1fax+Ussbsup7FhdAlC+J6Bqq7muAQM1akb
k+b7tgmrGDVczQDvw96Fa6S2+xxZ5OUaxtUbmBQW+SS5GpxN8YQpI4H0PWARPGZsR9EIirGQH2Bo
/y5g7mRXt6f2fgmP6MSuxlUKn68LqkkXOKI0l1YfUfYk4k43l8QgYtWkAeycLCSOgO7hgaXgGnck
sZfzZWSyTKx89knEZoaTjEHbhV+va1pwJYa+2UvdqI7pWFUEjjoNt/+ArMiqZ4zy9FmOzEBH0X5Y
UMm56J3AqevCvu/qlW4vSQTCn5f/ELOuIDAs+03l4WwvsSd7UZEIOxkGNL0ehFHQ4Ni9U2Qsuj0R
vEEOdxLV31oI2U6Ovm4q8RvBygrj7RwEgl/dLAoylAfSymv4sjh43mQ/3YAMGpk3jM4F6NUqmzhZ
FPZgUEr5sQbRngClPqizT96OkTo04FwOJzry1WGIFva/v8q3/tlG+9Dc7DiAQ1UFWr2fOhI8Vj1j
iAn7rTh/ROSXOU3OPyi0Dclv7BkTUcY8Ov6vNWHQ8VsAw5g9DHs7mONhJPkzO+tzW+zPW/SAi6lD
us9A9tmjdlFgR+AsQKx0eLTdP56ddglYUY0Vs5MSTixfmdsxdlnKmoXS3nQxW1AZqvEYRneIG0u+
osBc3lqf9JoZq+54FCfORFXLLz7O8ofe+b+cOwKGDCcnkyw1MArJLaJf0cFKvSOAkx5zeTuhVi5+
UhH+ezcRpsI/Ms+HJIg9dMCggJLeme2V05KsRKkBYQTQGb3AH6muMwwgxVP6yg5uBbMpqWT2tJT0
r+Mua32NPZj8lBOpEVPoTGJnSfe266pg0pHF5U5lNe9e/hhfaY0XE+8deF8nnWC0Z+1JIG+spLEz
aJKUj5KfMiG+POMDKwWgHMoBu0m4GDSCetjHJzE9dz5XX3auczELE+4smUo8Ld8I2DAKRLxdC6jG
ott/dBzhMEAZbnUifOCE6Me/RRdj9hg6hhNugD50AqdiiL7HVhE/4of5B013yEUZ6jbj22YtRo43
xOWRjr+VG2xcgWGLygrkI7QZkRBWH/VMVwnduS7qvipKUspu7Ks8FGuCNa36gPcyf4kWCD5FhN4Z
mGNYXmDo8AZpzk/yoFjz05kqUsRVGyVdZASkbt3FAwaXMFzvqXDrP0uQT1m38EuXfgw6s/Ab0txn
M/gVC0zBx7dcqyAT32yImJm3f6tLst4anFMsEfVn9kGLXm523r8T7MxbHxf6T73p+tERxqMQ+v6C
fYUD7qma1esoL9VFEKA73RLpIipmaeaQFYPv4GLHndpXvJ0q4w5ZWQAXyVuCAfomJXn0OsiCA9ex
XHOdLtqbJFnpOthZYReWi6VdskgbtSMk+uXjEXe9kdP7zyddrN9OZtPraYqgqUH5gYRKH5PzHU2F
tJshqYMBtFz0XjJJdandiZ3pLwcpkvxr8GiiI5xJIpnlyOHveH9vIrp2BAntvXXhWnDOiKSaMFvj
nPJe+mP0DkB1ljP0bH/X2DR+i1ex+mQSP9OfYp+qWQaRyFem5aCCGgeV0DJS4ySuuRiTkM9kdxhF
6j7NOix8H5bpAxxwrfmvCwTdhWK+2+X+6QlGnfHzPkESmje5ODngAwZvBA4RICS6qhgecnmQwEU3
OZfN0xXZWPOVCxjA0YDOI4YNj5xeZn//dyzta0elRd4vO+xPXJmE4dSHCdk0xgsBWInU0xZ/ZTAO
JKgUOEyY4A1NNO6PiX9QBfAmc2rYU6IVvBwBJ9o3f96NKzNPFlRcwGxRpGJu1xmUfxOSUnttZaQr
idl6WdOHyNUZ/p3mpLUfSVTD5oOoWPUjn/bkMXJeYIMcV6CsDgd8ZrDGhRtprfOdGegXDX9F+f1E
cRb/Y5W2WEh1/tvw2Gm9X35QMMCbMkV/ZkuANk4N1qzC8B0ME8OhPRQtXvG4L06gwVcovhuG+ZBU
7VtfBbHRDnf+fK3IVfIKKDr6fendXdblC1zey58X6JhY37sf8iSwTGJL/KEp7oQLve8kCAr8zafN
whOO5WXREgsikHpKOml3ENY/LDTVCbeHd1So6hEFMEzaWxwPQS003xMd4M51TjoTwjtmoDf8amBE
fcwvaeTvQ7gF5XZ7DTY3qgU/j2EdCsWQ9TMy9CS882/tbZz3fnLlKm/p7n1f6eNghkF0LREdURRw
IComw/v0JIG0Rg5fjUjQbiKNbgbzPEr/fL6zUq6+h/R22r+Rmyp78t2VFk5sSry7uwjOS8U1fvM/
NgmTU+lw/eCtvkZTHpCl3hJtvjAnARDp9H9HSw38u+6wdWK8H4EawzVPc1r8qqMUr8zTu7iVhzHl
vb018gyYZJuan6tkf3LCyw3myK/4BqPAa4t7hmlC/vT0WGDmZp97Y7AQbUhFAUc2JxToOfWbtGvf
oLAJtutYLe3AzpibGYxxQZerGHriTl+EQ9x2huZGXwor0dIuty2Ml5gjxrfPSJmnnq6l4YRiYUEM
b4bcSSKnlEqXbnTVSuB92ikYxeTeG4FSbuJCZQRxdcg02f4wXas63NYyXmNptiUyHCdgVHUGxZzF
jtlBM778zg6h5R1BJJOuRN+gTfGZKtp+VqM4053wspg6E0DvLiTuwmr2D6zvbvsaPxpujDf3wAMu
43+YsS8xbwVgjs8sYgvo/r7xukaqJ8E088OujCKB7XpUuLb9Q+TLmvvqHY1O2zuVxSUzVDDf4Gs3
ChJcsd9QauAtlz74H3G9yNxin/mDb3IykBuJTESuCGjoEuLdz929kEt5xlzrFNeW9/k0CJbpf65G
yWbxRdpRUq1BwSzGiQQnSUSGU1n8RGUjnWDtHMUWaz/60d3oP8g+c4hS1nm69q7bh5HQdvAMNN5E
GOVEECM5z0EXNjI5XsqyCbnKp/ifrmRArg/hoyLAO0+maPO+4NzZ+JLsIywYo/bsseNoYhuRaCbz
HbmsN21rLjy3FYyCw4jV+W+oRHh3oKWAFcuvy44gXumM1etCQhVRJYF4Lpu42ZWWXazDdc3XM3nW
dSYJd47JVYDWJ/ibZY8xEiHgy1Z+6Xq4x36Wrp3K/RkOuZKg4lapSo/mzTTBms+k3P7LIdXNASGp
CmPviF/RioTD0SUwKJzZkGsBE1vVw06KUtypVgpS+mUHxpHTx4BA3KYkv1S5f9RQJQ7jp7eB5l/W
Bw8vXdUNJoaIp5UE66LYx4AV5ixqmoqfr1ptKDm97vM3nlmynAk21TIFJwXKC85XxLqD7aQDpvQG
+mgdX0+vwRpf5Sbe87YNx7XU0IhVRdTFNzJKG4Mk2eRBI1rR+6yiT0vZblqPXsFY1Cih6Najc6I3
+suVaJoUi1p6m9R9WsL1Fsg432SRulKCOP8n9D3JRMJqytUwCJ1sYsWEbeAEUcga0wu0Ls0nL8TB
2JPYa0FSW4RrdQrMfD7RE8bOBz/PDY1Be/wjoUWNWoSC9JAYjG0Hdr6rwq6vdRYD83dct8sxjpiG
EgeorZ5Z/Q8BjA8npzcliQmVPhT7C8rV7jOwCVjkUaxOTge/XvAA2csd3dtMgCYQhNSSqqlKebNg
7R4XjXMjgjXx06VX1MUg3Y2EsK8ipQpV047OOiYz8aY05Q2HN6HUtjzJFwHv+GrFHjrZEgtr2Vi2
SoO+GPG8huqyT5YqHJOLIyMbh860jBejUMZnUn2imtGBFzVqd9bo+sCkl8omP3A8tdc3U0pTjppj
AVF0TF63fpi7zEZFHfHOve83wbOC72ELVbPBP1R7gsRzvaPRWgpTW+igzqTGDQj87izeggc9Snlj
5qpeiYuY9h+CD6+wOMeuM8Jujc4OXxPHRuwarpOCqJy+Gn77zue4jbxFLfMdpR5iVty9jNTCnZOt
dQha04x5LCJO0TqD6CJxzbqpqNWsQJw7NTiHkDYUIea3XQMvzM3mDQjUTrgXgjgF8m5G4RSkEcBD
j1jCROoHuVV2aKXqjrtxznNmr7rE4XQ2uVRMpo2Wtu/3dRUTwy6idMoOHkQA0wSEHjjt9hiQ96vU
TTly5nm4Pmza+rXRBtNEEIYEVEEwS7eNnAs0jtB9/CsltEzdZZNWzfm2vFgrJlnkj4zZuwPlQIYo
zeY4ihO32RndstenxDiq9Te8HZT7XHlj8k+7Li/B595OI607DsY5AF7OR+dl8PAusjMz40XzGzR1
j0094VedRNP5TJ1OnVAN0NMFniKLCA6Z+a77REuL3mfk3sgV+S47JcSVjFDIWK4YZ3Ziryvx1STF
9bZtGZxl69CWINX5v5eetrvUdXE5lYD0nQWmuqb5mS5mXYmh/ZTdKSCZJURg7KWIqENAXisOeYcW
e+wzhfUmgLZ4vT3rqf11eUeWXoCUxZu03JY45DAtMsBiRrhCMeLr9queRF0bJyKx9IxcRGecewLq
gAI8KnlKZR6GUxpkWC1OwlQVGi+tKyIhD7K5fGhBZPcrJgFNwIKAldagOH5Lt4SoMjHRAH0HULW8
WWj/2Jjw0DRq/t91sN4IJFpEEH+KFnkAsseJr9My9P3PbyPL45CoEl2j+RhKswMbipXro2WNvbft
CvWwLLvA7A+im2oGgAIHY1pzWU+5mlVfXfbn1N2GlDYAVhvuRJ/rOye07fj9vkNkmNtGAQavTUVZ
uXUzojkOjAQZiagzTJdrMyCz2O1cKheacGtLKZ/XHOaBfZmFGsOMlwUmo2VSGF9mJHOFfzBJwZOd
LW42HzVdbTgeHReeFu6o/M/XlqaSvDphb0kNApSAJlrbFbmvsFcujMXJ3/5HsYi/QtnHe9SRJ1xO
4D4ToB1EC6WJVVqtaYi/V+4nR3/gfpMQk/e2htpDxELXL+xqlZaxbcMSGtuAty8dr98p3Qp9Nz42
BIWtpwpLUO3TwFHlLTPlnb5hmbENOtk1T4v4etif5471NkCyGK8QshyTzEd3uszvDwddk7Qo0uh3
qx/GSNdk3D4hrf5TF8iDXikgtXCLZ7UlZKZEO2KJo+BFtwwo+x7N+Y+LkiqRogo5itt5InIuOoGU
y0w3QYbrZpCuFWzpV9ta/+dNjzlH5ibx5KMhbZnCbiOyP3UCC8QiRyg+f+y6Z99AEfUkhXClay96
4cM8PQ7H0I0HBd6Gges5/SizbFc6HTAfA5LidKhTyly56EKlweMHPMquwpRbU6o7pG9ep/0Hu7A1
h9OS9W2WntcAfjfUd/XjiAM/5pEvMDX0D7cjzBQ+GcXrgUPMmJrF8pl9s6E488suSSX9nF7kpZWQ
ByJy81Nd0fNia7yT+UI4UrLLUudkkCtN8muwlfqMjrZRhJCXSCz0fMSvarXAsr/i4vUZ8qRFGl0+
Xbt57p9JvxuyEWzS9hShD/aUKqitP4Iy9sKGr9mg0HB8WjFjlLbyJadhxGajUchWeYGxWSkv8aG1
i4f1cD1FQwVxqyw+PyEKiSz/lUMUzs2eApFvpgfbRQZmXhVGWJiqnX+bquUd8OSv1v5hW3RV47ei
MYwkUZAA8WvWoiMcaxbXOorsQPG2U2DS1rv4/S7hBxeM6OeOQTGuZSWcs/o8HLe4uvEHXlDFIOOU
nXOUQbmwgNhg68ezkngX+oFuDvsuwt2aAkKS+S9BAR1cWitCHbEnNWieVokU75kFefrR5LjBmyRF
zuAyekaqIMcruU5+ThvbMv/Z5B+X1lnefx5xFicE9/ANU7lr95abObq+aym/ZC1l5rC92PkrM7Q7
kI8EeH+ezs5wGHqhGA32VqkeU+v7lcdPW+DvTGQ9pW44SbeTV6ULYlqoRnGGYwEHxylFXCtVDx/5
AuKWSQvGhD0JGfZyBt3l4YFTb5zP2BYf3Gt0Wucd0GkOOc9U4qTvtVvkDkuTWqm8jszf2dWlT6ho
69zZwjpqw76Tv1o+Lx+lCS+ijuECWVaewWXEU5ovVFTmLkhnbsuCd9pncFMkmOoE8Iqh19FEn+Me
sFE5DWwcV9UNpP9d0/w89Lw1ePBEkA7fDXZR7E6xi8zvRB2wl1C+wj/sqeMqdQdPF2wjh3WVzErn
KDvn+9x+627x0kS6RUEVNKw3V0YiAqfgHaaplNPwxNBusgQ98qRoUBtZrcnRoLwWLVLNfkU/yzZE
nw30m8iZvJxsb56vqnQbrjAzPWBL1qdIwgda8mkSMlSQ567hYhGsOzeg+gtEPvanwgr103Gzzqij
eJ4UMgrwPM+tU+RcYbh/wolGQFMIHas5KWkW82E1TKtZkqQ6IXGRLM4j5HOWMimLgtVUGtUCfMg6
BPmXeFiqWISbSeEGq5GrdaUnZXZpNejSW8GqG2gTT/yxP3u29+i92PKV/HCMWAnhsO1MBPwEvMWz
ZCcl+EMjfzGXkESEfg2av+/2QIrub5hTByGaHUBs5PgrTA4v7EBXEo84oZD06g1tvWx2PmmKQNrW
yFBfQWN8bvzBU4x61BypjkhyRhxIj859wMaZbfRPcXiV7085amod1FZmoQGZZ6Z7QJ3GBKgo4tWD
fF97ZhQUG6VLq3U3GwqiGKMphoMPjgq2WlX+sI2GBJRcwAxe5ABYmRKLVTwY4tkCZXcFOEj/T39a
TWgTFxvt1wux5qOKRPccmekoz9BPM1SN9C0VE5P1R9jOZUr4r/UtWN+mQ4DzuMU3ybsgtQizw1mA
zaPRlNMapN8qH/1QdBzaXiLE7RJwcrsbUvfgBLOfy3SdriJtmv1q9bT0ZF94ZJZHJRZhr0mr+c0I
gVqNkUPIzicq2n/nLUD9SZpvju4v46n2y61dCJtVAhv3CS+HhwwitYdSQo1eFizF+kbOZ2Lkcx3D
Sfu9umHhQ2h6+Unp2+40l0Ci/rEwFaCQaHPLOvcd2rGlL7OT55EuhtuzvJum1qWSHZtSzBujyk99
vykGMTtiYquEIbwUoaNl6XtSvuy5M4JneZ08t0qk6hNI6geQ1ChvkZAW/ouyaIOd4EiqpJWFhma/
m4SUSWTP/vJM2+1in/VzwKH7NyDyiAB9nc+2qO1MQA18/951pCy/2KR40BW2WsZumGBh3GqrT/oc
Y2CeDpOufCQmu+VdLXKaSENRJNpNE9rJHK10nyue7+u3t9aA3+r6Heb28Xlq1a5LIexxk4BaKUC4
/QK8HKH5lTAD+vvYSdG4SkiTJq1D3I34kuWOcevFXh1k6zV/Xt/4clyehe7LzNW4NeCtlkDC8z9m
2murgHQjUAGrlC2O3fBmVfm3YYPSSaWViz8kCgExoV9oeLzzRL4FiN4o+PNDjYK8LTCie/BAMs7+
lqSYsbT2H5HmLTTyj21KP2qJMUbdTToBhny85IQrJ/2vn+YVBhNRo7NlVPImSgfWbU2mJUH65v8Q
PBlHG7QpNacJchGi6qN0drsXGDs6eqk7glhNwSjMw7zQI6+Y9sWieY7QOkSSttnHLA0QoZ8Z9PuJ
683ku5k9AKcKR78xibcy3c9Z2BvpudHI94l2vQGVtUg87dt6AohKYn6/UVGahlgb6PNYoYeX8mkg
gZ+USbzI6J40VKn7upvvz4hDdyKpI7MHgCmpXBzpA6KjHvAJy/xXAChnKf/sbHaUQwUea7nr5HOg
j4V2ts7chzUA2BYtYMfq+wLQCBc16XxgXhGMm/l4ZFkT1AFpduFevsmCYyOuy24+xqwyzgnJJ+20
bbaXuXLit8grmYzxA1BJcVVtJGWuJ5DWm4YsAAa4c0RCURes/4+z8KJOEBma/HveHylbT5LO/KYw
o66cDjBMVsfh12bAr7ipzVOzq81ZmeH4WsFk9T92NsIOD3qnFqvKnlfpePQeu2au1zN1oCUFVRqa
KRd8GB2zvSakGRg2z6W8Kx989vGkiK/Xgjk+DVEjUGjchCXzDqQWXUkVnLTRV1CEFEZa7AHSED1B
Y0YCPYAitOjFixsq/vBKOYMAKG+q6XwcnwF88hpZhzr8Sni5RRiVPc6r0UvCvZAZlsLhbNbXtSAw
0/eyMXc1CPuooQsL5Vmp3KhpYS0HCeebAIN6FWrdZZfCCqnj4246JwTWBFMepe1eEiNRCJ3DG5Xl
+l68PXIg13DuZgvWoaokGhJyrsrS4gz5lto0HxDAfMSLcQi1QGN1Sal3BIWz+y14zmWHp6gHlOB5
HvQBNCR2K5EGddGyyyLIaqiiXx+oH5k0Hr3Wpw4HgxdBYK/w80918u2/v2DCp1Lr1/BG4WkJOHZD
YrHpmrm5rhyuIrwufro0bb0otGCe3w5YomyjSxeQ1bymQnUH0qepeBYfX4SysQTjzC13opijGhIQ
i7bMFqS00GjzjTtiL7TxKCR12kWiAlfC97dx2DCdIShelG7afw0hyu1vPN64OAfW1C3gIqEMI2Ew
9UWjdAeXwgdLh4YtFgsvIX2i6KH7T+F9cy4Ua5IuqUZfO3o32ISbmMS3rNlaGnZla4eq7rBs82qn
1cta9M/7xKSejbEjyFEIgfNZlwwP06rCHloS6n62l7czBQE/ikkcL9cKoGMlsc9sFKeE9lro1p81
timRUau0DzZjooplvd2VQolFcqKUWGM0EPL1KAdvfEkVq0y7ppfYVSxUVeqDd2QTrZKXS6K0LhQP
4lTcuNpFKcmBHJ+ULneQ1oX83kEpuYR1vfnL1D4VRDpkU1UBGakE2ld5E3p7/kbFbGFbmf+GfuLv
ywVb3hTqk+t168imyV9vqD7MtMnsVEZwGSJu715zbDxegKEO96U9ygsANzn1YgAbb4/9J5MigG0b
2eZXwXWp+d1ZwjYX5Foc8t0D9opcMAa8AklkBSD+5uqkGnpIJrtFGEDiwBwD5VlSCfOKRvmK4z0Z
w36HiNDhhq6zvSnCH0lOzX1rd4DeEvvKaE6LsErSt0gM1ar0m06o+sryMiI4Oa+ghRSkXtY9t3Sa
NxanGGv+TwDJYhXWw1PK0u/o+CWKxcKPihnPEwg8TRUldVetkZm1Vsj59BHsHQdHhYtp7GBP8etc
HQBz7a3scxPFCkTcRU9wryn+kEPAFDhH4HKM0juA13GN4W7i/hmSm8iqi4tZ1x6TgjcRPLsN1p1B
pR7IxDmawjLd5acZW46nuke5ziYoScp5KUEKTqpqz5uh81Glw6WX2yOwhIWXtsDRLZhFNbGSRGjB
J1gTPSu/mflS0JZWTiJpUu5+3kbWySEmmwzBHakb1FrdqvYtjwnIuNZnYr6GMhJKgGYAWsobFTX/
v7I/dkEqGVP0vOQTVYCavaciqTaeiKpHJfS3yhq/iMJ0bJFWqSO6eH+NEsqFP0Nfz/6DA3VV6hMV
YTdaZpAJTMWC4yqQuoj2nw88qA301CKlCBrop7zYRChbOxSpPaJWUHldYpzH6l1GraJWzFYGoKx7
clwzXW/vSUUgc2KRCvXHOdSZzws3kQ1olZQDMtaVy3BJxYn7/Ah3k3FcFA7RdBYnAK2T0VITL0k3
NI2jjHAiWh4W92xptfQ9nFFqsiTWvqCVHLd+eGhB8plaKdUn2vvDS8HKdKqtsgUkwxd8zES82ecE
Yr6iqdSK72Ur19jGM1DaL4XpnLATiNA2fQeant8QdV7YtyO1gQstuC/FuGSpuHWvSw1WH8UctHT0
mY87ePW6ucnbMp6YjFi/0evDYMGjSWmvozHveXaqBpB8il5lUDoafDoiZshUIjAMxKVyPWWezEVo
DKthahkoQdLwYMb+4VUVgiQ09T1HTM7ggmCv6oZy4ZEkNdmzl3yE8+Oy7Ejvv+rODkza+Lgw6sjU
NsW4nTfxXuM4kzlS9gwEKF2YXH10HhT6QsLllJ0CkJnps2r7Wvx6NHWK1W1iQx1EPbNVsnNk2PyR
MEgFDs8BRLLnju1uPaC2PXK4zYys+eXbhr2NrbZpvIyoJRPr6x7nGeFuuOg7DBgFnWvEnKWEPqQg
UZlEVJjFbHRkpmVw1nOW5o0kgVVMUCelluwhgJWG3OFEIZ37qw1O8MQPLX/KZnM3KWOq03SC8AaL
SDGvhFozrrgnPa2Vx4mMoYJyfnxGvkMyzTTsC6WOmWb1i7FqjT6zCC2DHuU8r+wBIqbNHZAY40zw
HSdf8z0fHCb9KQBz/fGk+m6CBPRQ9OkZaASobYXz01dwiFGcpFLWMKWI7Yu7ruJHxn/Sg+w7kBEH
ku0AA2oKZFw4+7P95uhaRktw4WHXya64L9aWvc9ouZ50WUqCpzFQv2Gf3S1/RJZkfXd7ullX14aR
YVcvnU4Jg1T5ErMxHjah3Yb93IAPOxrLpVvyH6NurflNeborZrA5YQsVd6TYFk04zYCPcZwp26aR
PfVaSZBAUVpA1dTGwKVv/ZCaFaeA4gA6MHGMb+BL04QacAcX77z8ndWLkQcHp3dWXuMNrVAuApHr
xqbNMlQRtNWDGrIyD3X2H9VAci/0A3cZ7XfP5hvIENwb3uY43A986/MVDF/MVIekbl0ghhl0g9+J
eJzQCMeIe0rPuyaYyMxuuv3/Fw0r2Y/VSnmjukHo44hMIwNts+WQUua21N9kk3rl5T/h8ri34pj2
4RVyYIzO5fCeLUNU7vUpUAvp3BO0Seov3Yw9lxpdrop/Nh7Kgkv4a85DrIYJ0nVZxa7Z+aqADoNh
VeHPQubqr0RqgKTIyMlLbYlC9a94tDGUt+9HRc91Lz9PDV60iCWAD3rHoZNbAQyhcCQUSq3SzG+W
4kYx8nNXnoZaY0MHtulzvebJQ/TGziPcMbnYTBvkLPsA1JIso5R+t/gRXC9O5r4ZLZJQEMxLEEMb
D4Y+GZjFEzB3ZwvU4mIe8Nxb03vIHnEOp6gizWGInATrY5ZIf1Zr7Jw8odZvEAApJjYI0xVSdOV1
vT7h8GteE9Y/bSnVDvHoMdHWXDxb64xLSPltxe6KGXnh5VmDSC7lY5S91Rxgj3XwQkM+pOyY8Dpw
+vJLJw8Pdu64m5JfecuyNHoQTkOG15sstPCVPAC13l5dCfgOh83GHLjvy2Wqu3md9EwT2R4Fb1//
tN1zePR0GUmEs8xPJ6Psuk7MNBZdyFBFPGhFk5AxkgmvCd0NLlaZ1r2pOGNJOhhM+6gBwjB9jdfl
HBy1Do55xVYxFQCrh5R2XNBn4bJBhBnarJUC7hWbFOSRxy+QSWksMZFUAVjiExYCkqzI/02qKE07
Y+s+z4HkJAZbdmWCpk5zH4AF/WG34AF5ClQpQhUheGf4uxD/C4C2C7OgebxYBsAgEL2mdfuO299c
JTwPL6Z0d3cRqXqLkFUSt0+GQOI/z1e3Ps1zffPaeDOj9yBvumGesoCU7UHd5ygfJqrVac8Q+uiD
lqm8PyLcArzHmcCKcmXhWMd/Q7Q2AsmnU0DEiUyAm3jBLlP7+44W5sh1A0yEtTzoS74lDnvuCjpO
cFqLN88r+h7jSk24C3dM1cA+fe8Esx0rm+Giu2cfxmnVbWtaIx6kKwTgnpIQRDdL8CT8hmzgsYOn
uGq96nem2933hVxuOWPXiltqE72O6En/80mbXZyXoHydhUhZg/5WWTALkiqHOjI54FWDGQrVKyKL
BJkakXY7wY6sQ3VznODEif/GscB+jJPbfqI44Rgi/gV1MvbDi5yeVnf+kMTvT/7khKzoRZDjzoBN
0vLDM0XSh6jFXigVqmAdwKfrBA0T5NMVIFN28rNZ18np3xI7V+8pH/2E2EX6DI7c/W5pJwROJXwx
1jCn0TKJCl533gu2sGNWIdFugb/ptWHZvXfEb9T/ssqkBV18LnqY7r3lpLkKlpr/+cvwtSw0akPf
A5UXMhdjfBJd31yZH8F/PhdnwIy0YiqkPitM8lYkN8TTcxQhOh5R2CEye6+EKSKeKKU4iilHGlR4
VzbzTzS2D14Ci8obdIgGMn2G83oNobpTUyeDc1dipNwXFAOQ93HS63aavxI8C3X/WMhAtqbVLE6S
FHWR/keR9sFL9/2L3/NNnkMqVCYe7xRuPQbFOgwaroJo0sqkxb95OYaqetHLVWqj12cA9oYsKqQe
EZXBdSFNB0jpeK1rZpUoKDlDPuOtjtPnlSYrRDIA7m3I0/5YLfKJlo4WSPqAbd5AoOfhp03fx29S
/4WiIDklRd9rP6XK53BBqlBVMqk4+BJl2szWFI1uXx33e3iVseRX2F2HUSgBV4Yq12ojNZrB3vJo
OAnBXEIwjv5BWuriklQYEqC4QUmbT9ptu3aybNRugIyAMYJtQddheC962xQazFU9zQKZnSVn2VF2
/bJ/gbR/hKi0rlMLqa4egVf8GQp5jqhqKkOGvT6j42cJehbsdd9zmsQHGDED22AjTWX0NXP84Zo1
/B6pbsU2RPtBd6LjBwLU9fECTx2WiudOWUhXzGKlp31c5m8nYoVjh9BiN9S5LbqGCoJtaCLEIn81
D+uVKP3MHANIf5IMYTdDVS+dhf2vqlu+c8QH4w4SMUjwoy03wjHX8Gqj8wI52YC3xforNNMr0UgE
6ZeL3ChZS7bK8+qxCLi0lR0fAA+g7Bo8C4A/UzuyUswCuW/7w/sE+sRMQQEkJLRXOcPmfnOu+SC8
XJTXUhTYuJ7uzsFgRIeVWNGNMKxgs1vFOpQ9dGEMexEYC+Bvpma2ICQvPA1RjKRgLUKWFIgLk7XJ
t+ASKehruaLi72aDQHbUJIjqJJp055mxq5bLZjrvgCtsNI4RWXqHKJlD+duRuyPaXUk/bBDfQvOr
S2VbsvV+Wv7lopVvARCx+e1pgTbFQXQXlt7GqBadueDgUc+BBMWAYfHLFurJyD0rRRZ0rV9ECL8Y
DyNwHB69kQ60KxOndvjXCk+4uThFZ/ZHZKReRuwMM/rC4023kjspsti/FOxCZIEUuRVRZ+N1oyBW
r/LZz5QNCgj3qPl/G1d5HQXr74H/FQt5cPO66aijYAZrUEwj1JUo5EGtH8GvWrX3TQlgcSwY9zyY
IRjJAoBChvq9AFmFLzIYxclfJ/UHZNJ9RJfhTuPWeLDAakEh436eEp52+wpM57rqVunjh1WNCuv8
4lOLZjsopxsEwTqvTgKRDeV1AP+mJgZBrmqFHC5pj1Fb86gJFGHmd2LZLgLe19JECxWk5f7P6+Yh
ahzDnu4s76Xn1j5FVAd7j14QwdAeuDxyOFpQudtXKIbj8GLGsbjAxQVSSC0Y+kJmj2Tok62uRdfL
gU20gxFIhz86CQmTTtKnwVQp7pST6tVagHMSrwXvKcB5C6Q0aMuphGwsqtgnc5vRr+GmlyNVvwdM
gcxkmx/9sdZV10Q8EyJB57CIucgXWDo4WsGKrr82q/7jwdo19z+lyVwq9xmGwTsSI2Ej6az/V779
BxGka3CEGRsW/021NStbbBWCcu3UFv9uuSRgCDOd0PTGaujFo5IC1ZgK1Zlh5Dlzwaev7LmJTckG
JODHX6LdztOxmjDtiuwbmw9Lk+sMVgv0YMWA2ItnSv4lbE/kn+pFp/RimdHbHYh7fkCgE4yFS+ue
gLJtTH3ukQXOQmA3w2p8hYgEEVF04MRnrwSBg61Jb3liy0xZQ13eIGja8Q1cl2h/TRkzTnYnN52v
K7HrhibWeZcnaC2NUp1fCAG7xko5gwdir+TLMQznS9AccgV5UJmlxm+AFxsB0U2AnAaalDnCmXcF
c8U8p5MthtPsB8V94c+L3NO7i68Kr9MAF8Ek67ZQ3SB9K1WC6tRViEvO5p9tNTA0fd730escuPy8
+Vy6EG35/lXS91xpuS9YBAuzRoYfpGHJbrewr2bEmkOIXBcehKZN5c14POQKYRVTuzHLAyQIKn+n
29iRFXoZSqfo6jVCtyqOKzHSCLZ7u6zD4t7OBi65EtcVR9s432RYiAjuM4Ae9/OlGMaLHDgOxteq
1AqZeC4eraczQYyVXONB7fVjd3X2TG8+moaPoN1OKf3xgZWrdP8supgRbwPnQSMCrk2wSGqLsOsj
1kIdAPY0w2LDF8TBlDHV/4jcvLEOCG2mOQjWuQjkBQNC2czg5DKYoCTV0s06h6JoZsy9Kw/i/6oI
aGAU2RgO9ybkaNr3ZMO8k+oYThTuD1emv5CEOzmjUmw5HPY56bHtdfrIR1fPr/ecxwBF0RA2G09w
T1fZC25PyPzzUPAq3svYKZVwlLBi0eRSnYSIWlNoaaXn28wL3qLXByKsczNIf8dC+LoWNw9J9dmz
KPHoCtnMG2MtJDm+9hL1R8pOFMyg4S4cVmDqqxVfOrNYgzleZRM7qDaE14u6paMvrcX92GEwD88M
eYQBWCmY4J92skFB5ApFfp42s59PUKBz997uE6RNjtGiMe5Sy0gYf/juyyviuHLOGF8GTIgurvch
dQF5KwZh6x6jkB3mZXZdKZFJMUZEv1oZKQysoCLrkkU7fngWJ6sgqwLLR2M2q7WedSiFZIzabcs9
yTQHw2p/LNqtJxxn04nv3i/rTCNfkiiYFmvhyMJng2brYLBWxr5J/Xp1Au+J3+QbJc/hWDV7wbX1
JLL/8sKPXKGS3IHw9TKjc57ppfYSMRuZLeYF/DJl0VcNjXSxrNYjYIArb/rcW2ndtP3ZNcSl4uDu
GXlyUdDwzDh+C+X1xzwW0JZQwiSrjkZKgRMTHpdVHDtCTSolIb59Z3zYMLzdJ7olQZS91K1fO3QH
oEud+jcepqhsAI3ycuBpbrf/PZ1f1veKsEigC/agpCA6GDriAwHmUzvvYbxkQ7WK/FZ374/AkipE
qX+swp+QcvpsHfGEhvL32sJgn5Gk156U+HHBvATKC8L281/+7eXCPF6FuT265cKJqocQ/9rWTMa4
AlP4dWz4wBDULGlBaa2qI8gbBtK13RDIla4pFUZW3A0vC8QC4lQO8zUnISj5Qrtj7wd04axOLSyI
OL60Y1MIIUGw+mnK3CSMWI8VYcXHLWs1yXlAqmezxmlQOnMBihDGS39GZnS0BQklY2/QVe0MaQB9
l+JnDyQ6KAgX4g7c+eP5Z3THzxMMp37sYuThfClrHjGzfGvUuNPKRjRvosO0cBSV8CQPfeKC3dpk
o2fCQtvIqznymIDVUH83bcsdrfrPv6bZNHlhFcUMeNfP4yidK6yObgBXcrOYUylWvxhUhWiQ8afL
JIzSBED8Xlrc3rWdip5FK2NeQFYreMi2oYc+1ojrhOTIo6V9qa79DY9SobHz7llT0H71g6Ly2lA8
/CndetHehRLHzSwWSrteF60ZP2a2n7ChPXM62uCUgQW6UPdlUZIR1g6yPjzZzJwbTnwbHxBkKYaz
82X9rwJz4D/3WGJgZqZlyV5R1nLUizbkqB+cHz20cmzmDWe5KWnnwjhABbjSqW4RHrBfOgKqDADx
88igeiqhtyoz7epDAbDy+qTfTffnUXKtGvN5xtk2WcJdbR37IIeTvFB22Y3mZNEkJUAPMw7pohsq
RYa161y1Z3QMjQKwn7DgllQIDzmlvRwmBZHoV9UqqJdOivQTlJdZGqWIAxmTY6vX4Ewr3RUKbCd1
79QLepZgL1or0DD1fCRcTQU8Xu0Dkf0laNcLjvnvCpYnSEIITAQf+DJkBhcVEnEN0iIFjxzbQFWU
Yfm+L43OhzWVTAG87DcNYlTbboK3+ILlRX1iN+bNMLwNrDBwUSS2K+ajnr3XAe+tAJENgux2y/kc
GtNkcvS/0OuBDeJwOz7RNSFyr1DvdRvF3lVucJzVCA2BJ6BoIps2WKFxv85Ac1hymDdE1AGcGbBd
5fRvQcJD9yFiQQZJKInr7Q8EuXI6WuaMqtQ7sMRzHZbgTxy7/h2AfaxJOgVkQl1qwr2AZThEPItJ
pNf7/0HnfAzRuRvXeoALu/VA3/hz8mEfIgHvzdcbr0MPKK8sFpwe9shDdWI2xz3ibWFKOffbK+M/
k3PxIMt93FvtCluEupfvZ75neafAASrqzlV/oTLrX2Fx2ZT6g2fwFC1S8zjrSBR8Vu7vUPFEWPZA
9eyCUy0fp6TNM33GvO0KDxA4EvzgXhvfU7zA9OgXpBFKUDjBrn3mdBP/XFYjVb1HUspb4DRRjR4t
oe8+P70DjQpOgBJCffM3TWietDhiuGiGmhxbu2RXNEI2iHAj05WevYLdROWqSpj6Hkgw+OyQ2e0C
pp4xhvpg97eIbMzSRCeh3AMHdjliEFdYNMluPRHyv4NtYebup+GewB+gKNycNLH+CZhFdhTh097H
4iyjSbSVv24Zf3TYMICcE4U0x7x6AaH1N+aMmuH34V0VmqQIurc8ClSsTCSNz3A1x85z5SaV40K+
pyWfREzwZhBmNkuKeIilceJnQFkNDUKWzy60HEjynwHnpWUgJk/nAcktNFEpAYV/jVpggj9bQ+9S
CbqTc763vMs2h7CRXu3kcy959txS4yXi0BcbCuIlFrUGWnOVycunfmEUf8Py8atuyssTHjpSaHxu
nleyZYEwj19EZKMl7AOoI7j1hW1RC7GZ1bYNxe6auFEYtO5/8H6wkXarSxVFpzc2CPT+IkapBIkY
eR+E1ErM3yLECZwaCZU9ss2Rt+g00G/tIWBOyjI9yKqjNHAaDSkKEn8xTogA93z46/o5Z6co6d7L
lj/tUJoN2Xt9KyFGWDs2q2nb4njmkecJLfgIKtEybBRrSrD2wJEu4po7wqMfVvRvlab0ZObuw+zY
x6tD5f9OMOYhFp/PFc0/rHwybamMZCPc0eCTgFjjFVJwUCezsf9vH6wIfByD2LZmyT0N++dYPh97
xU17X3HVz0pNGZET4F/vK1BiQ4iGHk1MIn4QwO0TTp692UkR9Z0UwpgeXTYIaFVMylTFKEySCMFq
ZVDhmZDs6RLy7ehGLCfRfwqIVFDz8og0+3ihmsdTKESEkiZsqH9ODc6K2Ot1jT4DZRic0w5Qbx8p
KJDHo2CvWgLfTenm7Ue7HRUsojtLNPsqpRxjU9LJu8FEEcwDXtSKucnoG1dw7knmea6jbbRYsXrJ
ZoLh2YYr5dfp2n3tVOmNVkHLDuqi1K64EgDxBfMtVAK5jZ88A3aXmv7Wq5TnqCc4yprDbJBaiIXl
t7UookLTSpfksls5WYuZMwFnKyblCW023Qbu2iYpXhRIq3ONHcvc2TNYSeYgKQAxaZeM/tf5fBwU
0EU0US+sDARVJkZK7tGpc83nEyvzIesWm7i1qJ5snjuHswlcZ02IoFvcZ2D2laMLIE/Yd28ynvfA
Eh/+h2V5UE8NfmdxyKMPh7jutBQGFJB9a4Gx6dTsVyhi4S8qzA7rFO2m9uxAHnYW873u/ebZlTpa
105VZrfeRMCs4q5vtjbLQFUt9XojpmvYyFAhVwXLWAGCvrgcyBoP+AHE83JoD42Qn++SLH/k4Zwb
udASpuDo88fEh1PowOzDQQOWOx5x+y4d7qOBdUhkKos+PmewU4EqM1vxyi8cCWD1pjtAfe41qdZS
O4i+xBoRxy28VcwntQzv5snE/xQ/D3CWqutJFF0TgMBTQiEF7A8aA7eJPrydNIdLU0bUnCjc8KoJ
4twbCmVRNUNm2LKlsC4+IDAuFnnWq2UEnEL6JVI2EFKJIRy2GZpu1yhSrPMPHABUfgj5W4nnsafC
Ylj46+WUsK00fFKWxXYHM7OkGZjDgGhRV/GSdhrFhMEuoExi/Bwp8ieLN05jzLzVg3oN2xqvHJX/
4YVuKzM7dXKNqBtawqDANxOzYBqa4dkE/IAtwmRFC2+2A3gWRFjUhiJ5wbtjxFDJRaicJwI9Clai
GggiKq1mzjSZpknCN1Laf39SxpLuNCjzGztAksETzV0BSZfd/n9S7FiY3hDpChM9MZdwE81y+qVV
W6LwVADk6eOerHUj6IKzno5213tcebpkefqE228CE3YCwIYiVE18PmkafIMZQUS8M8tC+fFnoElS
IvkLfvqHVS+tBaPpcx1hhOBR4Mf7YNBpjzta06Q6XICzEjJluTZb0YeH352mFGfeJ61d/URsPpdl
vdG2gqen/z6CynhUXOm/yL7o5MvLdp8G47ZgQgRX0VScBg1uhoDaswQqJ8haDgeQ8NWY7088uDWC
QXNRmssBsKqYIA2eUIUKN8LZIkl9PweGmGi8RvvkExLnN0Zc5ZiRSb4QSzod4MWmKh0uEHYYnD0a
Con3zFjqjWY6A1nyiGYErfe571i3ElBdaV4pPz/UcKVPPz4Yd89z1zmDxnfSXmS6tjJ+ize5t0Eh
Wku+5z8gWtEihbnUXCz/Ixh1xD5/byKJR5Y9hSKVzaR4NGoO3geMvFNk/Nc8TFWyL9M7r5icBVL3
Z+0l9NqLCqjUIGN24Yb2g1IxWf1SWbTGvCsdhevtBF0uxqWaDBVZxKkDU9xQuENXp7AF0ItJDJwK
x4vFjj5J0weh5nxlSHFBf0K+G4gH6AcXv++eAYn8KwtfLSa8ouQi3eRJwQ9JnKM6wiQo+cWi+hM3
XSS8TN+QBvGVERy9unY9VOdCMcdMaiBlfhCl0pJBakwttzxqagIn7/CG46AqPh3PQuiBf1M7g3wS
z06OQOe4WuKPA87Oo/T1Nn3I+jb32tyNJpAxZujzl7PRC+S/KbWTxK5aeiAfpHFo4xHk77lyWxe7
OswxNPP3/SWS4qiOY+lzh7X4KtQT+ukMrfCXHVZ0N15RgcWCWtrQ0PJlZhqsEaEBBLAr4EJLlsD9
NItcV/Ml+A7H2Q8yzdjJhqlJfh+evowVAB/sq8/uz+wvz5b6g0FPtwbtCaVnppj7ljcvfQ4+bnus
Aay6dGyTfzfVsSejuPAL9ph9lZBgMt2Jm3/n3JWmw+YphcjmzrbIEXsnG+CsPR+VeuIsJIjw1uQ4
d8rxYf3WrJSoeEqd14XMq21Qp0n3EJISaI5omg20LX4fqWfdwAaQL75l2fFOE3v6tljuRD9x5Smr
eK1XZZLqAp58i+59R+qJfpuG/v3n9DsAtDtZFMC78C+vpYmYrUYDzDMVg5bJVs5T5U/wwduD/U3m
NjcDdpLQuskwpNgao8MdTpz6ActzUpvORyig3s8b2Obg8yBb3MVtB/rxi7rZk4qhWLwr/2tcOCzR
xE12dWWCbUqxZ4o8RvPmUai3aTW2mKW3a3iETRsFjg9bhZU4K8fcHOOppImZe7iMLFeKh8xH+Vmw
S/RkbTJl+Cj8dlM5nlMC/GoZ56IJasux4pPRORwxRZE1Nsk+RFhtK+HK/7X+q2WDv8ffccDvdDVI
9ow3V99axD7I1tvSHEUbcAP0s+SVv18xKYA+sGX8TOS0a8FCYTxyCAgM8XtQxDzlvHzPky9V5gnR
Qde0FmhFl72DLPY3+KRBMNU03XZgNL0k4LyCWtBqn0c6pwRsvIYwS0m1MH7Kf6QQVis+0Tr4vnpo
F12XzqgWes2kz0jAUw+oTu6Tdh9rz/9zsY5O+/24BlBzVvtFvB4OqO9rh5volmxtOvDEYgLx2Wvs
roM5fn450iupyzPHcWSiQFb0orvJ/4YC0dehHBRBZe3qxK+IU1lxIGVC5wdfCXFrFZlWAPaQMiNA
qTHCrwep4G7T0QIrOVvX8j0sBHOiGmarTui8w168b9VIF4/ldzDEwsx02+KjcK4HuLevZkNJ4gyW
j/gMtD4I2W8FS92Joi0IDs4Wtc0w2+ABesVBYLunvFY55MytQvpGx7OMnRkZkFxyxb812pODUM4l
gNpQYke+RIPETBo8zQTJaZPaHLZRf29GmKu4UJnNuv7L13XT3/S88j0djphUWxHLCDpRd0Yf+FD4
+ofCH/wKC35Yuqx90glrkKqfxgJF0Y+r6OAJDZ4jXCxReMbJoLhnzXChQMqcrrnFdObemTSCXTQh
nFOKslPG4k5qK7pTurRs0z49Z3HRvwc3cRzUwnO8SG/l6swAl6u84mOM1cuV4bUqNK90i3iMfUoN
w/YCwanNE8wZmiTBFdP9+kelE65LaLBPyePe4wWfOxa/EGeYqMTteppXVGdr037xZYwAUFPDog9Z
aZUpyL5sdOC6aMOs4UHq+fUis6WMo9E1j0sOGDsRqttgwn5IlwWQH96bxiEhT6STb8eEiuV+Ifuu
DtMgMpKiJrum9M6pE3EjpzgIWhyd+Dz9eFWMO/zG1nb64NXJ3I15+y5qZbeVbkWy82xuQSuCPBbR
CQc8PnPY/bcF3DyKrMhnvkZjhNrdTOJk6q4Ga3EL+kpKvUPfQ3zCPnftOISymty2fWXpfNE5LmS/
46ZJDy3RudlYkf2FEZdRFo+C9e9xIHBaZ0zzFtHXef3A+jzUMZ5lisuytlg9KGf9Mj2v0ZZUxAr/
1QJy69bFeB93WgoSLaDRep6MNFSIIBP9VBLiq3eVqo5tK1R4isZS+/d4NHhk/crXz3I692PFhybP
qri9QQ0q/gGBFyQs+a0kZamMytZWyUnytrW3RXP7+EGREHDtTBU6Jt5D9ms3bApcqE2TyzwS4fM6
CCZRxWUCAOzQF8v4QBwiNg+WakNcJdmC9jPHFsxbDFYFiR+zZ9OEQ4AS+KULZVkjXKqzdC/Cbmjk
YlmnTubVIXV045mah54zjH9sIjbb0zGE1Y3DLPOdYmfYRuyEPory87PghAy2pqWAiI7oZ+78XTBk
vd9rsOhTaTtB8U7ayTJL59z0Tp6TJm0aQf7dFvfPS0F0XHztlX3VOzp+j/J2VJnuFcRo6RRXRLQw
MQvE+Yne49X69JcZ19lydHu5yoif0au0/zCfUMV41esgsxasnRTbzXjJbjg5yBI4wdcMkQnS1J1j
X7lm4bsuPdINEZCyl0munnxYE7kxjxIL/sB5QBzjbECFG1BlszjKpIiAVTfDEekKSRp7379xS8Rb
oVF15a5ADI591cMv52IH0g7G2SdxC+zTkOVtFs7jzRbbdg8OFL8xet2wegMFR9GguHTyt+KRL1hI
GbUStgV9hfDcv9ZAiiqtJGeWswWF+BIPlCpL/LmmczHkNysev/mZ+OwvkUU1QwvMOzQbBwzoGish
+yOWd5U6nvGsMScitvFtgzcQmLe+uNyJb+zo6JT6Nf3DfEW95pv1gAGsjuregir2MxY/BAvVAoAI
Vl8vTgDsUN+jnSuhFN69YlOq/oVvL3YMucDYzGEUq+iff0pbe/8IrLXF/qB9cqSI0q8oOheXnc+Z
d27v6mziM98OOX/jEewu+U/t9foIXMvlsMCWR8zzGvTeAQ5SzvJTZ40ry67QF/lYdOiAKxxWICqJ
SsmFgtWLcuXTPnOzpegpvC5up1OuHHXSd1ImkxPLcBjJFFxlrYjECVtgtFylt3VFFaK+Ljh05v5+
avGh5RUOeJCKHjfTyYsPV6NkKWkPr67TfQjuY7TnZzrPLWNWt2fl3adI4EMZd4kWGai14lw4m4ol
Wggx1VTFJs3KXnOmz7EWifo5dTIrNgG4sBAgQc9W2++sxYESSZykShdkxW6KkI2X8ovbomaZcPsR
3ipMwSOEUZ0zlQUZohU+8uvy+rvzzAtZ55e6YXDqwmtx0qU/v2hP5yI9YBMd0/i1udL3O8khoFcJ
QrUE+0KaUrw/PkUcrn8MmsQDZPr2J+wIGy8UoghAjH0x1FyCrxnKFGi+Ga9NygzQbaCjfbki9lR9
jDP9GVxAfOCbnvRnqw7c3PpgjXse8hXi/ijRj9nVPTu7WfWHS5Zzbzlfu0gjtHj/1XFOmyBEQhe1
IJ0S9hLBSeRXybSoVuDZCxwZUFBZHR3V43zn3AHw/zfSjIDaxhA61qDiBTBHkXWwYM/Yp5rJ+ucq
i9OpyvgaKnpLA6N+raYXWpxe5VuEuIx8hp4QoKA2zrpXgG0dwl+NLxbBMH3fCopwICR+qRLVC4n6
5mH1S45ctn7xb2Nz5yLZlVElFadqpaveyMYgS9ed5A97GCjmtXXH9CL7P+Z2fy7CgyNWQ5bgNnWo
fpUxrzBitOTrEQVAduHL0QKGtxd5aNXaX+yMSx8ChliWSUZKGKMlsaGms5H+Z3Q1g20aupQOQOs8
/uFWIT0TzZ8SRugRvB8anyVqx6EDbA1Q8w71lX9NDhZgQnaA+krN5TbpHT+ivLoGP+2krZLCnpyC
Mt3r9vxzzACwzwoGg1/c3RMI4PnxIa9fsU8+4JDXdUB0e4Ta68u45XY4wfkKNbzVx9OizkQZPZii
UAGT6hGvy1psqbYIllvJ3St5vyrl4IH6EJyDaU9PlrCssM/w0TRxqyo03iiH5IqHIemv+UpACQpz
auPcoP0kGhPHzCTmUkTvev1WO1hhW0bMxVrdcAuByKzXLwqwP6Ofzbc4rfb9v7zB4BleLNl77Cuq
VNh3zLOOIpieQqw5pUxWnvzSNOMrVJgG740/3BR8OKVk7PwTjG/O2N2I8TrZcJlppAopwSLRThOe
zP0pwxUma9LvV1LDut2D49dk7tAC/5pPLy42Gd8LkWruV4p2VmhNnpgmsIAApn3bVZT8kYGgbUWg
ZO8+OqCXSgRKWlXPba0NwFtXIGS6WXZVfOjaBMxOpUpvs3jhb68na+jpPs0Oep0FykhCla0YgrsB
VU9A+TblPMqOPZ7q8MML2pXwNQKQp//ahk/U6BGp0Mw+fY/PSPU0hPCLSyav3NGdLueeC79bPHzF
tUAtGeVkKTMZiHS7OAc4x6v19dSQfZJn4FZJqz/TJExpRzgLSaMCrL7SygzMtGJK1gsJ/tNto5FT
3M3PfqwFNstCSM+4JoOWUUUoOaEWeim7VsgNngHnuMUiVWeSfG2/aAun+wXmOAhyPT/73AYXcKx1
bs4fHujczHRFHUkTsEF+nr2RUlsge+2p4BgZaXB3qOvbaD52HJ3XBn7EJOMT/CsUL+PiE5SIqxmH
sxhUG2CuXBrHD0XoIFz1MeqSZm/Dc1kKIjFI8WCk/7GFNeqfp1IQxvSWAs/gyClBdNj6D7uooWRF
APs6S1aHxWHFomZ9SkDF33dL7iXL2B7M4+ZM18uY7LVOTdDlN5GfU7QxMmYbFY/nJS3ohN6OXcoD
IHs8rjJ4w9GgskAisPyRPNTpdmhQiChen/8GFbihlvUMKmUotO3xw/ft5fpdXbCbjOb1L+qLGIOS
C/tKUz3VWCE2ypce7L0KEvJwCn+9kpE7etoj7P6n0yMp2lhiV266LOAp9bdVuIdoupTOXByG8oXw
oVBCi8aiVWWUc/+LE3Z+rCaLgmwIGZZrd5QyeqvB+xvdzocTd+R/iMLF1v0Sb/SsCrX1TgiMm0l2
NMBpoouXd1ltsDPjINbeUMDm7Adp6ie4p5APCVgQAbXR7NHa/qSEJ9vHKCgWkBc6lc47PNQ0RoTE
AC562uccQtKDoURUFRYTUIIZHj9pmR2Ybs5tdMFt4T+3HvwEu2mHdF7zdHCmFVs28Nu8vgzBE/OO
7JcoYlja8VbJ1jikqmgbMlqlxdQC/M+4nE01f5w1Pp0XYpV1wAdyD+ZRvQdjMyAJ038catYQ7VCi
yAx6wx8Rv8zHPiKCC4qcQi6CcoyV3aLOdtbRndfKA/yDYZ4bD+uwUVYmdBtbAP5W/hmRSIx5BEUD
rKq/b+tAsl0QqoJFgjsZAIx72Pe+POhJ43ceMOzSsHgq1+FgX8Q/JT7g+FYmIJqYcmBxdcqrMv3S
efav6yrA9oitmgltzb540Wf3G7gKQRLEuCNkolIlBLKtsGuP0JK8oop9sKH98x+rwEATcuG5b4ux
Fgc+zI+UvNNL89lhFSrHFgNWJJi85gVmljj/IlFVgVvoNdSbulq2Ie2akVHJHJOaMH+E6G9TnQGa
ikebiTOX+CAxzp5RnfC8dNpanhn/U8oqYpDRevjyjRPlbY3mfxEzy1FguX79eCnACrS/7eSmufMG
dXeNehMJuUBh/wIaD/bngg8tQEagTlYv1vklZ+VeMoGjLTViTurbeClS13h4Z/DZdt1gXfkbepDj
+GSKxrS+Ml99s9GcDtT1l/ipMrXxgl7NDTdtzzRL/scuivAZK5UZ982kY1okNYU3YYOzi4snp4m+
pxMZ2nba+zzHSebuEWR73OqlTecCVGCyDbc5xKqSW5txQiBfo3AHQWys51yD13MJSiGqDm4CnFBv
HTAuogad/jHpp9XBIH5rhSzr64+Ziyxw13n4rAv0wACusxudEGW/QAOtvGxVh/yu7OsnZnByO5Yz
HWqUXxaZFNpVGR8ICJ2LFzekamImXk5nRFuM3IDMnXSr8x+izzFJ56jkzl/KcckN7nWiGUpJ/N0Q
rcu2r+ynFaTaiQOm+HnRUVf0sOimvTo3KL007JCki4UeNd+guGmVuumEBE4mAPQ0KWWU5P/V3KDl
zurXatBeC04Fa9OJq+E983aSKoGar/pqpCxyUodRynrNZQwHke1KqB2PYs5wdVvbb42rd5OJqE9G
pY5zSFTsYxmW5FnGTGNqSfq9Qh5RpryHySYOnmJmzrG5gPZYQ4MmHDgG4oPTckToy6A05Mi1pTDD
ASo2Bk5wMKuKt+3LWwB0Ggxmq/CMp6qLCZA2MSHkQaj5lRMxgVcSn+8ezQr+/VCUObjTIp2zmxRy
lTLMppMzfn8iXqya4FlmLUteue1I2t7c9fu6PDGBBGYZjpbbZ7ZiVFHk0eLsd9JsE1WWjIgGnHsL
DK1OZXzJbDz9rBV/YbUpNEkhgEBghK0Td0NPKpwJNjho/vB7NbXNkgwg4o32xXxMEn3YFsG57aD8
wBqHANYpBWDPJcdEMqelQWcx36YNCy4uqOjODiqzc8/cuzRXTiCm2PrbKwfg05i0X7soISx2NL9J
ukLcdMpG4dKoPH+rxyUUonQPWemms0tj5LFamQE73IOLmbTka2jZUqFeHOGZjYOl3Ecx2LtkB4Fa
wknZjwnizz6abaarGdkJyw6L0EOxHoVCFfbLMwxTmBmGj4O0HGl666boFYF3AtK8pEX/nU1wKPVp
gssVYH4P7lPT+G9BB8QUwG4rtk2lbW9xEWGcLYHKghH9OEB+E6DgTSaHk3zxQr6jDaJXXHEIgxR6
T8xXxLSl6oP4GPusBQ4G7bM6HZlb5JC20grEcBQ2N1n8PSbUGit0zuzAD+O/mqtXuoQCgU83SWjK
9AynbMnLGbLHHsVjbUgPznTthcd7MK87RjMDqiBxoitOvBIYeDeKvIa4PDrP0bHPh9igJOGGEwiB
H2V//JvBkNKb6rzXJ1nFjGtYcwbLjGLDPh0Ai3syHj9ZkAK2AK53hETXdRi8b9YIOjBuss0nzgcy
ksoQFk7iyFPd5q8DkJJP9IEhsMkw+BD0eaYKyku1i2iyKcAcMZQ/Uoxx2LzYjfMaQPY4Mo0dUHnv
K9j29RJ4x4i90QyXp0azI7Gfw4XewS+nsej30bCv8U5pInYQK+ljPZahvxooBAUsieII1d1rFx89
6Ek7O+TdNmBL9LsAIg6SH/s+cj5w93Yfuy6Vi2i/RmD4OfBI+x7ZlS5CIloB6kcpqAJ8PXnXkgvr
s70gloznUzYp7Nor2lVgrlJSxK1XE1J2zVT35iyaIFEoKftSYzBF6EdYu111aLEVs68UMMXLSz+B
7MVso9AN6JZJfdQYOGQavXW/WEw8ri2+s5qsGsAzYqAv+N9TEN6uCqSwTG2OHXmHxF0Kgas/nV52
3inqHcf2jxapO0v58SFiaN/9IU04F9J+PRdl/NQATaiGRHo25aT6Nqyc9tqX0BHKWzEEzmXtZhIo
+wNGtuvAYa3CJVS7A0hJd1mxVu47PRxYMJ5SnRGhB+Tgq0DTWK20M0gzKUvk+L75dAuhtZqov0+a
IwxnW39MVAqb3MRFvMcZEcllJYRtekSkzJxqNlecOUALBzZFGk/NCV49+m3Ctl0wkc3S6uEknj49
6aBq29WmKFH6XAR2A+5rAWO/b5l8fKR4yGemdgTVyR8i/NW10PLgINGjUS+QHbwUOEFYYjwRtZ8/
mYa+OwbxnwpjIO4tIWMdY1SsGwDHpQho2sfeZ2X7WUhxlghSs1V2J2gwYY9byeTdUq4x5WHof4aq
HeDQ3mxlzX8gmdT42q9Z1X96sU3F48kn9ZUMmQ0JSyWAqCrkZpCFYjL1qIQkrcwev6OOfXIyFCNS
fV1TUlWP+AE4Dsl6T1ddd41qGsxFclmBXo5M+gP/4J4/DigGoOiS0HL0KwDpuBH5u2xAgLMM8v0N
xMKnv4TE0cZsBaUwz6E17S1X2DTBgV/k7e0sGPQ4zAtXXFu0fqX23mdW69JxQk6oyPog5sGzWO6Q
geRWTVFXrzk1WfrXYs2bjj96iteWFnVt/DPM9gXRKXW/4w2WK7ZshFo4PAP8MjIK4kt2lI56hAvv
854kODWH1BfwBNUDDZS2qU2WPr6HibF1v5VyU3degCzalHXxUB0qVquZFO2ehvEt6Kr8xuNkV4gL
1MJ+B3REmmqET2XCNoHAxVP9HAwol1U8jG+2ROlJtlih8pJqCtJSyxFXt2AJQrlwMZHEoBKqRAvx
551dvJPBYX8UifS6yis4gZGDyVBJ4aPaV2QCC4XwthPv3QkKbQruZM1iEJz3AXM/KjWAd6dJi7xO
iLxpUbDClKM3r3FNWJjrMdYr86r20Pr8s4tCoD5+qy3xZg/MvY83OoXcxuGn1vgM51/osMd93Gxf
Q+rJiOsPOwMB5tdf5PAJVW7ohcVPYZ4O8rV1Tph2VZ5D+ozsO7Gsvgmv/owf+f0QOLNMMQNXUV7s
vZcEFPmY6MzOPMHXE2x6S5D2ShxC7MqNWx2CDZBHpA+kFlQZkQnVsSsfPdzo4Qk8Ztl8XOtXUOYr
edrEeLOOa8F46nTDTRtbwwhodFSnRweIR1xDxpnicr+FuCr4yq5GUTWSAy+3GwiTo47b0/YiYVcB
+SxH7FlN6Qw5Qe4kaIG83/r77jFjs83j+z1Rz1DqvfCNfKVBaSJCYKI/TwjjH3zxEwONzxQIdFOI
6hK6/z2drb01Eu9kFspHLK7VmpPYx9lRy8gfDuT7eieYXgkLFbyOvaKiXwia8OwVKw8w+zx0qYju
JfknNtyXDNYIKbyrnC3ek6wAY5p9IPPr1StJh1SC6ad6QKkB97JHEAFDFvsNOlocn16nQcVxVU/j
tHk83JXWt2jxyAGX7zlqrNv+Zboqh7cuUS86uC8JKte+An4gp4EMsPtZqE4FIi8AuR5gwjcBPLqh
j5iUFzLcdf+JuiVsDnIsMMHaonnp77iSom51BDNyIG2tIte3wuTJEXfN5PP5NUpQpNLpZ7Q5+YpM
+O/0DViBsNobV7m+HxrPUj/JLXqdOuesa+9bdz1qHdG4KFsBrjGhsOlXs1LsJbtOonhTEMhP978Q
W4g6F3twprG/Zzs2IRtPU2GtkaYwxURKvjVW74UOZr4J06j738QsYqwf+1aiSalyAF4bXLYXr7an
xkU/UeIiSa+BFrd6h3cZwPoujSHPWRDze0pMwR1G5Rc1YW+ZdYwhi7D8fdVW7/Qd1Z6Tu7feyLUv
ndyaOCoJIj+cHVDY2eQxo78AL91i1uqzTNmgBDZPugI4Ku0dozr02LEre51Fw+/Y5txyQk664/Ml
JcXfWEooU/uBCrEMQNzAZigDJAY+iWC5i96VWk2KS/hCOfXPf9hrxDX10g0IAUSNckzy/dxPype+
IjPj0e7ke12eeIAUX+iGDdTLKV+FC5C3M+x7eKAGETmnU1hzf8Nui6nCKNlA/XoSOuTh3n4ez3Nq
rzDLUO2SEr0rd1revS9jmDDHkBU8+/G8l1rR/x9R0XpTM/N6JRfoEvaEFfaioqvuYHV+SG35V2Eo
0FOva6WYzaA5OPyijf31V3ZeBsXrOoSqstxPNbRnR2RiwTrcUjih//PLo66D9WwRrbvjCRikgVxM
iDFaHIWZBJYDp9bCfz5FzuvXo8CrxAteJKppaLyKmrKbfTVDmsyZ/RXqw/fN54/JIsp10jsTCA1y
cuQn3SpXygAwO6LVT84Z1sdiVA7d66HXGCEQ2LHI7Ycp2nPnXlyafMvzmoqwTvu3NRa4hlf4ma+x
uq1J8eguJQzgPtyspNQgoSgoUU7gJHrx21s7B4IdvrY/N27p3K7pZh9D0vkoQwmnc9NSkDqdaOg/
5OtPD6RHw9B9b5I2/mytkpHGLioGhTI7KgirUD8yb5+zcusteDshn2HVoyToJgj0UNtpMVJ8QWa4
zvit2Vt6bfh6T2CF2p9G9XfLSQUlgq46F+i0d5POFNA/GqkQQLD2cRbq5uYn7Gfnh2J4BNtz3C26
Kv9UPm0NwmSkSG8axG2VY0xcGeD8eI4SUYCvLhN4S9nNjUkfp6qHtohPqsG6s+JiPsT/1EATWV3y
vc3/ZDhSbJoBZpsagiRlf6UdMtDVBnGbmAzfyYBRT6/KMoQist4RDQMReHAMsKuFIx/m4HHzciKM
2PN1jwVLCs4R1OBR0bsgRwORxHg7rwfQcBhEQQv3uYWxLpqt4/g67KEPOiK6JMM5oMqu1Eh/LTPC
oQkKZVwRy6A8RP7zTaWuapmdBBZNFTEgy+q1eEABjdh15d0+XFuLY/1edcWO08NnvsQaxbuLZr8u
+uOYT3Z3CU9vSoPhWBUx1GLpsnw7Bh9w5vu+A1dGcbVDEowtWAoxjJHn9bWaPCcg058fZRwJAtpO
UWfCjwBYndY3LSE4cQ9pjWN78YkdAd7uMyAHvDFBcznGFRvym22Y+EJTNHIeeD2U8rvVyf058LgE
3u4Ho7xz7sX0cgDMyAF5yqiq2ilv8x5CGMlkLPZhgUstAMV1FUVIIjYsMOAw4xpsFGKTkJSGJbSo
wygW/cT1owHDI/xUQBnjW1wxh69UJT7E2gCPq5forwPqiFF3DZxv80j254DtICnNCLTgtjo5skAb
HMWpumsNvHEK+F1zBMf4LLgcbG788Pr2ai5qaovQkFFek3rbvrPoLQ0wWSapyRMfbOTL+Yli9xPo
WxtGaYVVrOQD6P3jMmld5xZKs0PkAQdWLqbIlF9SAHIH0NmOEBTL7kKbhhu7WZN6h7dEfKL92NeW
NPgRy2ITgDNzbzy3KqTwza4XBPkA8XCXPguXNe2KXM8wj5eXPhqZsFpmXQwKO5qeQ9yKvzf6icO1
jCcUY46ZvX4u+EEueoHOzszhJU4UlLYuMFnZZzJ6hmB/Z+3i7OXRTFun93HgEBSBEr1OkSwPJ38t
HmCJ3yNhj9eNNd0p+RvpqjZFnqhgRQR/G8Ds8Dv7ROfUCqn4Uy4ysGTjRNAzynwXrJ06iXXhVt8O
OPS1ttuAShsX7pKClEkoTMVzKz2fb4bEAhbyw/YktC9HTNvldjTy5NF4x9evw6/Ohhqa3VYTCCUI
4/+yJqfKcks0Hr4ZwWtXkD8zknPk6cj2PmfSip048kFE/Ab3XKOChd7rTqFRADC70m0BtH65tY3D
71hFIp7O1PP5L0qtpCKKfyf/VW70Gg3a1i4Phg/dPKLqIx9agogpFFvSZzBv+1euq+wuSZ9MCYAV
hRey2g4LWU12CiLrRNfZRwczuhq6S4ODm13MgRKmXldwby0Z1qvFkhbYbryvwaeu//jZiyTS4qWU
uAcN9wHbFRqjRqVZDnouusMui6DkQLWZpcMjmIXtuPemjYDJHAkmy7vcxpdwbEC0/4k2S04QhCGF
i1kjX4A0gG6WGFgyjwsKdTrilt8dsDkySJEw+/RDegtLP8RBm72W+DcsoqR9B3gfyVcbGsmmaKHf
RmNeH9XmIl7+gLGv2cGhfiZfCIvF61+AG1DnoMXw9B7OocMujVMdBTLVro1GTJiDtAVULttHSZa3
CHbR9oDCXf+BoQNeUx3tUUJ85Gsx0YKpbtpKhgVQdYKKCToO/Lex/OD9KfAHLD0cEy/c4n0OAeVj
3ad0Pyj28M0M55db+F8tsfhiCg/N3SIdIWki/8CfE+ILXjZKTDTaljYPzqIpMyOcxGMcgF8qFIZY
D/qy8tfjaqsfYZBBgr8pIh+xP/4TKCVkQ0UVj+vjQwIO+26G42cmbcsNOOtpkY6KXtclIsElmXrv
+eKkp53+kyH0M7Ja/1Q2bsqdu0eQlCfE6rX3bnCMNJAwvOlDLhiwcY19tlI69b3SW5C7PJmowaG/
kYOx+f9o/hsUehmh7N2ytM1PvlIJJ+pf4BD5fxpBJYdBUXgeUD9yeB9esr0xAetHck4BRe1G04wv
Wsb6yjkM1vpM4ZDlTkNwAfCgwawbvBO6MLwo1s1+l7tw28/W9Hlpnr5EPsRBg9C/2dfdTVY1t3v6
cJhJb+9I1bNvRt4mumiLOgOcUMTx7lP9NlihBDkTdE6sPxgVe9TZPVG5YZ08aKr1O1qhfayXfHtZ
LRHIwK6vvFE1qKVKJQrvP1HO0lMxgyuXDDvQmzOHCXrp5q3RUC4okrwfWl0/n9d96Eu5UXhXOkBZ
loaMc2Q6JhlmwEvPaRbRtYKMtkbGb3dzK42VIyzkcK5Vbz5JYT5A2P09a4mE91q04ECXcuIfENeQ
bDEnlihvvKtrMa4jUJ+yC/SqGNhcEfHZ6OnBVnSF47+KdEIW1nx09U08kSIVCNgt9ICvd/Qmubpz
Wsnbr53ntdtxYPDP+e7sR4zhxWThZ0ZY7QlefnJKB2ZKpiqfPP/kR9TC7ylvMh+GVwrNRcpRTEr3
3KgifNiuYyYsGuZGPQbHVFTmlUcW2ZV/Q+rcvJ38V3+/OQMx+BSAF5621FgwPQtHPy42jBF0/VWR
fpmHUfkmFK/UyNdlXESHGWhq7OoJtxyA32zEaOAw8Q7jBvOwkK7yUwf9mykbHvyv90AeRqabKKmu
iqU8ExH6U+ADcqFvdLuE6or1F1RMYoxAxDbS6BEf2OZXMOFRGAsB+VQrff7w4bg4v3VLIfByTFSl
8wf+AutrFuZnUXp/D+LoMbP3Z3VqZN/sROpEduLMK6XSGlX+Y/mdAjCK6BzmQwGncWodtIN8EOFt
Kyio29UniMJVfDZqs8O4uG6HOJ5+pOE1VAd7rGecnQ4hm0Pb1MzKcpkTmSmL+s6O44rccCRCFddk
aNbfum7smTCAZCPwv/9rUE2zvTDnTo5vRERZRNPGCwUyFLZXTVoBkoKk8u7MPowydXm5GFXIrTj8
hpSlcA4ssyYsoltDJrJFexXJu1+9rjrvTe1LeTBQcif1dFujT9p7KuE6kOHEzcF3WOATsydc1+rH
0ATmJY2g3qeWV+ZOKSJmH5phfK3OTa35Ou/nMqQbg4g/xQuXOPFVSytyXMayJja5SFkAaPvD84Yf
vRKTZKyIphBj8pJ0zqNDdBUAA1mx52LXShcrtxtiYTGUgpZPV8O4/2PwRm17xC59sn6kELMTH9fC
XM04NFWaWPUf0+vvREvQr+js40M71izkvd+jFTh6ZI7cOx2JkL31TM3oPayuzrkcgdId/kqhHNC6
Y0qSnZTtVo/H39m1PlOvxQx0KAcwOLmf5gWBiRVVuN2g2II71+cxBqM8T+DAIxwKv9Jqjqd9yUAS
/8khrliMRgI280/SH2yc2V92x8hXvQFxUS3eOUMhaE01XZUlcLxvXDuGQMrEPX+e9+sAV1mLHgeN
dUhWx8cwgzbGiDeWIAYsmvF5H4v3Pu2IVS5RWuVRBNQaINHVoo+Dgoj5AiGSMLFYUKkujm7eGQD0
7pfngy+3WKsNBSo5Cy5Ojzp/4+8bEeUvW+Unz9T9rtHYJkRFfNa8ygF8SP7dF4pnc+oqn8WIaAti
9lienOQ2KwY56iPpF2uoz6cGD4Y7qJiNcxVmiFQxOR/HlxcTzLQhQsJ06a0Y7NOh36jZAvm8HcQU
L41ooKFyyZ1A0+cIKSVdheIe6V/IuaWS4xg7GRf9SU19Av0yqT4rbNg78gJsQIa6tD9pCFh1IfcQ
omsn9ryiVyN0fMMX61m+Z63WCWvsBfp7T7rge39KjpT8oyxNVsjT0KfgGLQTqtl7jmKF9N0NMgaH
3G9OAMjuG2/YZJV+I5utdkgItG+vnYjnw5B8tsiVXOybG5itK86Gd2DjJww+RCp2XTzlkRY+Razu
6tVxtDRO0axv1/s2jsTDAU9mU19JKG4P2spMgz2kWn8cGgzQ/mr2ol7Jr60MFzLDsljXJ7bTdJv8
9pmqBYPGZ8BHSYs6M2niu/wSYjnlgKGEWyDlOCdzttUqFOAQJHJiKv6Dr9OTWhuEbBqkWjD7AYNm
+BMRx6t+ARooQxZnnRxCFSFSZRF3nvE6CRCz6jtzCoXpzjm2B8lj1exkqyK7D7KR7KF9ZyXEOUlO
Q/zF2kKFZeZGvERpHZZXSpyAMOXWpIDcdRyBwtQVvOvSJjUyRzv7tdt36FY1ZZehNeuIqmlb3N9x
dsSmumligL6lIamcnhLGX6xpOFoeCXlqqvoXmLAooyfwFPoF2ByZ5VobeYSPBf0ZWDMyzWE86FEV
PXCE4A+ewgF/tzYX6gKiPa99WhwB9vJ2WbRwrNCCtPhKbrtuRuCa1llt7+faTdKysdpC+P5PKwLM
GlzlWQkzzUOhZriouzlC80/y2u0G8uYtx9RDMr2Q+hJ7k8AUoD33xv8bpf7CuIMu8sZiF/cOsM2f
N98lRFUaXr6Wob53vZXL/zIwrl4DGs6qcKfHz5FAw6/aQyFvKcv3KFHGcEB8BqPfXrYGaty5So+Y
V2PY7zgtQ1J7ebDz6whcoC55JRmd539M5c98QQ3gf3vwT2+nlRY4mJnCzbqn81eaaJyxQVHbgc8N
SSZEDq9msC4RKhr47I+ATnxG4BnnYEW8Rja05F02XULgscoBOkdOnrG6vPBdlmBnX7NJZnU380ng
pWVRnteyWMVkgV5F3IzFketLrJTRDxUm7zw4tlY3OkXrRLmqK5Wg5LoMq9EeBSOdIUW7SPXKAOt7
pCxMrXsBROAkIqlb5XO01GPHxNfIt7BQ9beajQh8zPtsb+oE4NO2rg7Bl76755gvddaVqX6UwouX
Sq0VdOaMEjXzDFOnwzkcmEeewIf7GGY/mPi8MzBg4q0cCT8Pt/XvUfkERVFvT6wVEu/PoqhdbvdV
yNDrB0frLp9zeGFvXNqGwHmgdtJOf/DL06m+YPb0XP7B3RAnEkQbp5DIgDjo2B4lN49IprD7hs+V
RvpboNDAAS6yDwkg6qstZ6oW3uPY64NecSNeOAPw0wVoq3faxGzKv9Jets/4NDPu8M3KABBxly+I
Zeapg6RQiRNBdCwnSuQLctj65YLxjyUpI4H+pakVFbo/JiZkiUCTJvGvtXWglpm4xy55rubXLG3i
jEadnnCayGq6qX2Qpr22FzTf5ozDXQgyhlgypGvTL7nKZ4gzLX0txKCMaeVU6SHmUV6wXpNmyIxu
IxDGoWTWq1VL1cvvU9Ie08lPZOfjf1h9GwDnVpGVKgSJ3Ap1sSjbYsKiZdUbmcfPMlC7CmUccoC0
b4kyZ5zwZBUh9uRLqxjvOd7nUHrwMEq0MVxDJMnpZm0I0nMg4SPbpUFm0yDw5HViXdY0VFDcETA/
getb+2Gn8XUSPSWTl1vHi+HWDKun0crvMH62ZBx7Qp2vdlP+N3wgJEmOFwQbTj1T1VHOp7xkp5cj
GCJpZ5yuULcIK4mHNhj2nnOtvA4V31EDkpUn+KTToq87FVeEblFqvqDM3wonUI3pOTMJs1ZwgiYE
Tqkwxp3kUo4lzlJtFc8hcEDrLzC9jiKTdlqb1uuvzWUTn8Cb1F8wLfgAzVhq41ulznWPVeNY0MhQ
VdjWsSVMMfQ3ng7ZISJ5yYAehNvrG3LCBcdiOQVSKofEI6WJOVvNQ4WZ3mgvQwUyjAFpxoTiRLrS
GEFL+GTdK1NvrQpGkd5MBTUZpLAC/obsjVkJko3BQS225OeXztxyzrVY2zeSdbJxjwwOP4d6rY6v
DBD+3kQw1H7IuDrm4MraqVuL5HBcjGPwZgUo+MHTbAyDpUlarEuWJusP1WNdG9dO+neeAaIN2/9u
jzLkU7+Rk3JkuXAiZk1NvwqOyl6LUW4zi1yxDB0LrjXM0LNk/cWudBaDJJ9oLqbkJCWLLoUXU9lK
StJIJz3htJ6Up8s24NNg5q09RHPXYpEqBKZTRZNi3lrO6JX0i/DO7T2heXGDu9bFwLXk0oCK9+XE
sLbL00fqoipvczSvbjZ4aAJcM36mRj+abuOpQPMegjwoqGkymByh6kMXAaXQ4ZpAP1aTh1ETfXxH
axLNzkgsGD/219AIHEdiOVg4UxaNDGbl5WRhXpXabmvFLGn53SW2ZHK3E6us2JC3AzJCf4WxCWbn
X/4CXDPhYeVUjfu4SUibRd62FLGKRHq5XzmQ12l9+1DmaOMX9kcjpQ6dkIMBdKrI/S8ujuZ960do
E7AHXn/Da2TJV3Vw2WLUO5q7Nn0UoJjlkeIF6FTWKicCxFf7DoIWac4CKg1LYJDeDUw/F3/jjIiA
Vr9Ll3UD2F4tw4n3y/vxoOXX02OGpueMqQ9HviRd4F0AXzd+JQMlfAmd2egLN8mjX+UT2Tzd9z6W
o4RYzdPDX3fyN4tmwYN2KSrNUxJcWAd38xUsnqhkmOPeDzUvLQpfwtVmkv1yDEz77b7DtBPx5CXw
12UKrQW6qPnpemkzrhe8D8uuvtr/tjpot4G73Y28vtiGX4/XkQjAAVF92i37d3E2faVa3KuVZVgd
4bz6TE8CKnRDliXx6VEZ6xnBcPXhJ+UDw6GaCSy5foiWEsAhvsDDWpim7Vk0bZh6SRGXlpzfwYaH
nKsO2iUw8nMi7+m/Nn0yhG+rN40O6lhHF0kgNzPoT9pIT8lCXx0b6Rw39JlRurOupbNHDIbjdVPL
2nOMEW2QiHCNtqo8Wh7nnXfHWnjRWmXmYL+XMHD76gdySVhtMXpOwpATslFczTddl5JnhXDZmDKO
/290aQZQvhnOkUKGE/YDoAINeAM2NMILJYP1m9Wi4/0VtvtERBuMunenKX0wIBsTFN93yMacxvfC
uMxd8hrVwUSSeBnnkMj2PlZaKmQR5yJhgawHwVXcxwANlArZ4dszHy4G/WegPQ9rJNg32kIY4bS1
AVHD0f9ckXXOCsxjerEB6pLvTfddSK5XaHf7AlWLdodMJ02j1pXbSdxcO4S9hQoPREv5Hm1wgWXf
Z2QG9rAuzXjhNQWuomf8Pzau2GdFMoXIywR/vtS74BZcVNtDhLT0yAv4sjdtVFuwSxbIJo02gUO9
6PxwKh4b7KXrPMRLJSC3/w+DvIYh8aZzgaHenWiJXwa6pn64ZaeVHnYJ7dEqASJkor6NNWozF6JT
IWrbA+qp1SEpfGKkngo+uqE/9zdFBGA8dVDKJpC5ACniTXJW+oG+TIeGp71xPMnJfhCdIfIZZJIt
n2e1A0jeDKaP0ThaHtfAF5gamVhtmfubcd/7/d5CkHF1iV0BQdSjHRxlpTziQbcPT1pKnj20hWMg
DJoz4NNmLHucGpRrUsxOw/Ep/nhW74nq8I6jl5DcVnfT+FDxjt9Mc2AhiRh1DEBxqSzRYsvhpMtM
eE6fooMdmvXQjCuJ1E57K6PK8RMVLznO715xAItvF8ulbV1uQYrOkGpP7guJOC2UOqy2u0LWutgO
QOY+0yj37IHzWhHa//pttYOF5wmIVbLnpqKfjhP/yN2bBO0LdhADN9Lsa/1y/65ulYkRyYtI1djB
+0LV99eH3DPOgVKjMg9wMveT0hn/uNwr3TL6WXx0F9Fb6qGUw8F8fs7xae4AtgOeQqu7hKGeH/Iz
9x3ugPWewFVawm6SiBwuy3ReUWeCmAKEtPYPLuMtXtA/Mb9urDfa7n68Y4J5BqyFHsYWTPSGHC5v
lnwzXIvszn4Aohp7bCQL8GShEBCfPF7cQ9jlFEI30hYq2DVEd8GItU/KkyCeKOJgtubQ9jQ29b9U
rLqDnD1Kde1T4eWa6LnAy32XUfOJJ5p0mndxHhrOn7YeAzzbUW/B3jW9CnIjB/lU1swcp43y+m5q
ISqrUQEAT1ePv0NPJUg8W4R5WgV61XZGUqp67eJVJ67MB2+TN+mPNAdMi4LNIicRmqeHwbVCvTCw
D6NV8YAuQB7OCOVIB6S0o69+OybiK8dc3oPO5ETNSp6JRzdchznj0X4Yj7MrGLhNFdVrfD1V0Q0I
zya7qL/4p30HDAqS03OojWjPbdgPiK13CokINTpPtnmltwahWu16zYxv++mJi225/2Gm2wUPxH4J
+nb+XbTbnauk0ZI3ccPbJnQDlMlkICP38hrebUkpdoXJp5ahvq549oAuMQLQ0eODbEMsJGW8xz3L
QEvoiZQAKNcd+nzr0+XtphjZsFcolGDh1Zignp465V/HOir/pBonwblTmZk+hbCpbY5ZaWacVFgq
fo2A7f1lPjrugAY7GXJlg3xEhuIaUKyuZlpRhH9lBWeQwK9ZgYNAlZ1hYtkAj5wDzc4F37G5/s58
zW48iJ8fw8tx8RMdOT9VgM2Dgf3aEa7jM20EDFmA0C6l0p6FA3RH9f8HjSkQqZ6t6TpknQTuKMwU
JbVotuSCR6EbklDZsqfmgiG6wqLRgUDJmapG8hhzcSLZ+J/hBJbE4MzDc+1wv5ZlV691l2dY+Jki
gXAdYiFRXJFJMFWdpgYvvmMBWV96vj+td3X3LK3aQd6AYYnkxLrXovWvrvTQAGA7u6zsuOcH+kJ5
qXAmaUvlH2aVXugjHZS0AULsR3BOUfm006pW8fk2Fuhn+XQscQSr0sAXaMddW3rGAJXcm3TsVU8q
uhcdbqWA+desNBZZJm+/82jUALn1vhHmAEVuTOmRoIyStDIVO1oQEFzzM6TqNSh4TqsVRQsqNnM1
5yEGrRovpKOgD82dX/LIYY2HntECYIAkcGlizU71+kfzAWcdjW8w2fmDOVnfnLrGeA6Y/le26Jw4
/oMsKbm8cwkbaip+X47KuRwgFjP+Rdrzfnv7rA53Kv3gIpprQpIPJgCKoq2dIoAnx380WgpgI+Ra
vig/lrpnJDvuF+8iuErAQoB5u6Yuh+EmJXrjLrl1gq5JjmMSVtPY+a7MegZFQWrD3YiBRZlRHlj2
jdy092Qlg48faddU5tRzHShcL3qVH535dv8O/yXezWCvDV9ZeMf5dgmcwHrjjnlwRIeHBqinWYVX
B00DnwAlJ7DbFq/yvg2MP5TQRprldj//d4RcrKiXEh7dW1pwNWKB4EovEaU+5uFMiH9Gta3Lh27y
AYKW8B12zoS50ewjME+Flr0EdYhyXdykKxmNo+6vISNNwDKN7V6cJCDDP3Jo6UAC268IXwOsza9l
3d2oo83yYVk0n9wyvXiX+D/k7RjfDFfCf7xtXwjO8Zz9rembwiwvPMVzZhAKzVogQxrRrPetGoIv
ivqY6AVwn2CVzmKYVtfK8KnxdemakgeH4fYTXsmKpKtlo2TZOpByHJ48s3YZBxWrilV5mXFx9YHq
WLVxL88x3sF1Q590d3YIe7ZBVAOdTNsbe1yg4pM6Dpdly4uziDDyJs9MCqxeXHmp0QXaBTa5QRDh
FJhpBHZkDeshiD1xPQVp7x2LRvkDH8WfGaAyENQfYHc/Y88s0qBNYV8wYnXjeSfWIC7b/Y3R966R
9LXaAWnFjBTxoQTmyIst9UdSHttj3quRE2OnMurKnYiZSlOILXYFjWoMgtOqpyItDLvs+lB4kLWx
M/rtYXQXz3Da4QP3fnHA4kkYNxPcXVvCBgl8tOHoKJEEoRmMQVT7B2HSNj6Ys1MfU2pIcsC39P4k
Dyv3l87/4PmdLvUY8KJlinz41o9L3r1iPJkzaQZnQx0dMdQXmHv/vA5aPm1H316A3TwrEOpNb65j
xhdCExuxQU/OCEmGd90axnaxwwHavhCdCcuUyBHMBKnKpxKQx4xzrKpC6e40+1R6P6Nxr1j3gCsm
UaYR3SNulLgM/V1NtNxX/znqILGOiyFs/MkgDUzMMLuWfEtfXFA4Cc/1l7teYgjW7mnCe1c+pKuJ
jHn7/YjpFAX36eonoGl2npKnPF8gcG5d03ebbGw5LgXsdu+Cm3S3tdaxb2/oHZQC25/MG7aQW/gd
OBBs5kM/zkTFp6vK0nL1LYq3AYGgEA4PDVAwoOWIuh8VpigBWiK5bAImogspD2STzqaNiO1lbPZ4
DX589GzAEFzNaqSTCtm0SO/YzO9zKynyZ2LT/1bBC6l76Lj2YgeoRtwANUYafBSrTkOB+lqxx/O0
DgAjPsjpZ5fLRebzE1fwEfN1mnEGUEs+VGoYjVx0LeTjrd2ASk4Q6ssEyaKsGfBvuJ/hVpcmI6KP
p7rjfxIJzoPMZdAmC2kWdn9fTCJm65m/4+q95XUc9q5f1ptzIY4S2Zc+FPl4/xVzHZQtfPOG30NS
f8NrQ4on/mbEhmlih68b3AYtagdas6T3N/qhOtBiqKrO0kxCmD8Tvt/k7VHIRWMimzIHV/gyfqTW
c8Yrin8T1p0vFVTHwU0qiZn5erXFWbdSFWDnBvmnrcpeVWarSkWecWgZktAAjMMVXsT4y6pXovc5
jYI5ecctIdivgMIGpjtQVvI6Y8bNi8VeU8l9H3SfbCgdcNNxWUzfJ6szrVGf48V7Dqzx4ECR5wYq
NqaNZo4JbqOSH/TmB8tNRcikDDdea6hlsuVonyNpzn5DHdqgA8ZEVavUUcPZtwzSO6jfOPQe51nh
Th/kWSjOi9N7h3iY9MSj9sl3nnXV8lBDtGbzen4SUnqZunn9p1SvVcbj4m8+/ChylW5KcU8ZTPEQ
RiXTrrtNPZ5OwDXHfrrUzSswM/mJaP2MQZf8vL6XEqtxImb22067PVbgIE/lOVnKjN7Xt4omVZEy
41PVnMX5MNScMqvmZjY8Q0LvPoZ35zr9BUYyj0XIkCU911IonhGSc5x4EIF1kx40s6z8cIjBNQX3
xI9gZgOoGMAa7TKcQ5pklyv2oGY8Dx/hM04AeaNBdiCuElq9wANHyOD9JJMyfi1gsoCri2izUz4j
+rH5oK9uT1x9hHY7H8D0FeGwEnzfC4XiwG/vKb2s7kPXKIfSDT5FKMS2OWEVpMKdeLJU1bkgD4MW
2uXFyIyAKRXGVccJISHSh6VhQ+0xgFX/7Dnoz163mU0pYBw+bWKDA+vCov5+KrPM5LOrqkOLEYHr
tYs+dekVo4G4WaFJnB3B7vhrSjdCH8zUme+Rh+ZoAt2doMEfZxJF7t1GFwXa4mmUjgm0skanlKet
i4dtJK0j9qUQVX5ddjmqFyHuuewBBKifaWQr/EG+6b7KCrBvBqijtpw1mqDyHKc3V1uxufdULXwV
xmK3Nc8Ora81po1bwGgeXux1DZy4wtAdDW6vJOdefW2BNAmdcdToUjZB1dTkWlLtMiQFVUFWe8vC
NK+nPopRJnukblKoteLMN+vrTeF0vXbUd4+nuyO15r6Xxb4ewpyTEZ9lFNX7A9d6GvhbSlk6YrvM
1mmvvI4R2jbct34Y9dzScIPSfSXiny0B5Bs6SB8hPLVhLGZsZ+w3uUIfl/jqQaIpstwdOsgtOD57
v05qKEsNo+81kRiqQJju8snBm3KCs8vrb09zw++7OHR9hbidaVZ/ykZ+wSTl3/qhtQZB0AApz3JQ
vHs5eBqv+C6FaX1k6Xnfkwz/Fa2Dca+EBGKCKdsWN4FVDKLePTQq8A403Z8K7qsqPjWCbCtpTXOt
F4CzUjSAv+s/7qj6M4YcQw45lATW1yJprjWXipB+uHIZZd5OfSlGIahZ6z0bpnpzVTteagYiJQd9
Zs6cKZVQXdWntPnsgLJbRWCnUA/WnlZHu8XyjZChOC4m/fMuCP3Rt+pT8GTkTZ9qL4CYlhNl0+6E
ixsZ4q3VXi1+7LEX8D/OXUmv0bGCqKbQsOADCwIDtWNjz7TWoL+C7rQvzQA1Jucs5uhddZaBUUUL
4YONpVEpaUhqA2YhaUMFFov9/122E+EpmtfwlrJE2x+dDirCsXUUzyheAJGhQIK4QL8CX4qI3C7h
CAlUw3ftFhnVuUpC2fVSsWiQiPe0h0xRqEim+zbhpuxqOVx1C+WJ66/Jez8MyQCKtnYq7ltHDka8
KrbodTN+GG90RDoY5ZEYjGufgZYo3E8P6AzYu+f6sGYofmjs00MfS7/x7ikcO+JHkSm+Ph/GAW7d
fRtqwFkZ9WkMgzX8uIUjJvRRGCrU/VGbdDIf7xKRdiI+eGcurIiZrOpxAaHpajI9GeT7hXyBIXtt
qQIGFtW5O2n2lyFPaKihAsb0v7lkipn/NlVfPRvUQlXAGkp6CTgdqpS5JwflYVzSWXPHo37QmEhT
rTEW05IAzXfkHW6Ej9MS49xDtsqjnTZ9+Z/r07M/5P5V/+ddp/9++nCriALcrRfh1pguUp+nvctK
qEEaO5ZCYprRuV7Sh+DNjyW5sf412Ebn/1P72J2GgxWnJcT8a8ID5GyO2Qsb65JsgAD82bPIjNf+
jlFecT6PeCbqyOrWUBrMCjBsAtTU+GjCVKaw4I/quQgQsL/jPfKBzxfKlrkJ2fiUxmf9OnwHV8MO
YTEQb9hkhDJ7c4i2OpS+DeHEfhYr5fLMBJVooudKEfNPU75/nibXCi+bARBsm6mqL1n3BQoBfPA8
F34vcpgbIeqeU3ZFryc+Jfk5MCdPHyDlLXjPon+lXpOKYEU+8QCNIAkmbS5veyddgMRz7kaopvWv
4mcRXdT6G7uYq8zmLfFhmLmsMeq0M8trgm6Gw1yikEavawrskw55xtl4v4dQt1nSRbetMALPz2Ne
vf+5AOUz00rHFQqqc8TEGmqTdG1IDpSiaed9TdInngy0F3vo9RI8ff38wTiGM7Uly5LJp99eDBWq
ztEZIdlN6boatam0ksRQcCLiXrkbEQ3W4DOR440ebjDT+YZDAjdfXOlNxuO7ZEuhEUNr+tZbHYDZ
Undrz7+IZl9DZBPWQNeoTCcyKR3S4MslP3LgNv5RQ/abGOHSv5Tm0lXZu4zR0Z/lKAPvyxhnE/nF
SM1+4UJ6XB1D7j/QtWVEDDlyXT0cBYk7010WeVkr4jEd6fm84DIacH0i8tZ9onjiDsCL/o27WJnW
rvwDvFYlBbqaYF99FtCwUYawK9tbpTnlIOTPUBokhT+XxUyBGuN2hyr2IAf6XhfeQJb7iMMbliE8
Rb6rurpYUlliw+jfHLyTPmX/jHYaDbzjWP3WHzVjmqAA9cbbfjLgNFlQPP2L1jBFIdApJ2C8Mthl
GYMZqNtVwKGOIBOtgxTKCovVM31dOIhFw9sjT8HCozV5dI2Qi9y+thPK9rEy1rGcCWcc9zWUG1rf
JgJ0tJRfXwQE1B+1RcM+MEoCVhG+thirah9114jEn9try/e2u7ZftBnnetHicd0p/W6253DJmxRX
DzEzsINgtBGY0aVmn1dtx0mNpyMYLG98JetvM0L5MLGlhh0AMaz0stmIiFz+aO+n1k+x3XaXYCoD
HtuRUH1Pz6iGwiP6+byINErCaRrh0Bhj/ugt5A/bbmrS4QO1FILGhmgXLAUqso9Y5ZDjDVoGI9Cy
ty76pwqloaE8PitbREg9ZflfNfwDp66k2ORvmo3x1xA1zPBaL713mZi/p5Kf0zG8yxRIZOcpZcTn
fYAboFusl/yPDqVb39XL5rCvYUvWh3I1JRBNXTvSd8qKaxGxV3jwWTfngKqwvI4O6vdVxEUUzzcO
ZH1PMATnfx8upIhHZFBL0IlPKizPBsdm4UT+7ppwcFf+vRLGexRIOE8d4rEcOARRR1DqVRzfbzyZ
eTsH4fHNJ0ZGGk2+ql/VmNKe2z8ZS6XQGuDzkUUDBz04mhDfQbgvryJASc+hJXaywvU43f+BGFKG
qq+ZL8gSNN+SxACBzR5FkSMuL4OIyUACBJM3bo4yv44+B1tSe+nfcjbf4bHYGT8cO7mw5upECVnp
btgv/9JeJz+T91eT/x2z79827x7sV3cbI443n9C6kSds7tPXQjwt1RersqRGpm+PBQC1aN7lkvwj
m0uTHi87B/qMK7VKc+m84oM5ZhUMbZWPICwPQKLPCnvsys55KcO032J0Ls78JLQmaqki2nUm9g6R
xpO/hPfR80Q3A0mMM/sjIfCU+fA1jqTCUN5/wZgMIWdcnVCVk46qjsm25w4CVDx1Dmw8oNm2foBT
o4PkBYbDp1Lwyrh4g2Kd7E9+pabCgFrWg7oaxD6MxSoo//0tfD0DonHVa6S+fjOvCghobfLv2oIN
9J+x7I/YkQfamhAAbUNqkzfti9Dv7jRLgkWsMt7sUxg4zxwk4Eec4BicnFSDE5BVTYrZzRQR6/E2
NFl5R2RvUNiMAuttSWwX451wE1h6KUmlbW5seOvx5MMLiz1iAxCnIFX534yMpllWDUMFORlwEIJI
0x8UlH+6F1y/95AqG3fbVbw9CuPxV/3VVDsObqyog5yrIJhcqhcwViisr2W4hSrMW1dLbsXmV0PI
Bs+YbGoKkEyTsTad3QbUFtl4KCiFuWQRkB2iRp8oI+s+xfrjmFHYWFimtO2M+whefJkOQVIXuAUY
BvFyrfXowbvLt4fi1mQK14MoECq3JOO9ak7tYXkIAYPYR6Vi+MfUBceJr7twHfE1Zv33473UDDKE
4csfg4/JfD1rxF8ULvwvPoPxIPnf8T9ALFbU4Z2tXq/sD6Thr3BIVB+EsYrvTDOyXs2T+WZUEkAL
BLf7cwAskp+khHyEQqRVX/Il6R6J2Rd+UBbNQ1hQDrGEsfZIqFSGUlbRWkN6WG8kFpT572dAM4+R
1T9/1frVK8oJVRWpC3FxThE0zmsg7VRWTd94/3Cxdm91fi6F9reb5Itz/vjVDJICNwpVxk7b0Kjh
beWWyIyE5eAnjp76WNXC5ZpIQMr5PtCld9akxm9TGWUy1Ho1a00d09SeTbbdQZUs9VZFdCk/ELMx
4x+VwTzJmwrSjRe9565MyQ4vdShV0hvcesU6EJZCe7tDBPGHuiwWSlTxeaw4UFiNNEWWcDfttO0w
11bRy68vev4burbYXNviK7GRC4kAGf+EkcdEbb2GvHsBImvt+UyuBkTFuqso2HPCK08KHBp5t92A
gsN11fcJ/PXXMR9Go8ceM7skOIZvvQVYs6HYHgecJw2JLddRYOgRhC12ubOrKC/JCjMnEhdjC1jE
D08A+ORrWmUN2lWFf1IsuZC8fSnGRuI462HnjLjTFMobojCh7zPx7iTmLE3FHd4IsAkdRs+4ceu1
xISZ7juS5a5zbqTUaphk8CNJo6Lx1c/UDou7Jz565pd5FfYh6qb1LVYUYJQ6I7lxgHHEJ5P3hmNh
ts1pJsTI7NWyU4mjUpvBaa/2pIyRmK08OT8jlgMWDUjslFOs6pT0nkVwidJaCogL4wtfW8kKL+tt
/nouQFwqb+BKjBG9npKctL+8QYgoWsYMRAu7T7oBHE9Kon2Zk7SIN9ZIzkYNJW5gAVYS8CuhmXYG
2UjA4N8mgIk/VhVZwpfO/0nTYOFx1qHzcl+8nHYxZWad1amR0m2/dtF+PrHJ1POQGuR+EdmfsSl+
qsOadVjggUDqc/Sz0HHZd9QFQAQLjSr9EdxiYt4w2dv8LivFltBtJcqcnXjmsrw9VXvjTRzzFw0Z
V0f2EMO44yfxelpoQ6y2/hppOdyKCeHjOTaA4kx9ShhKw1GbUVlXyqFloSpjING/0e7j4Uxw7qew
WemYY4DVpK9sZqqTifwzNKpKZR6G85Z6poQqA7NhG64JDvggRepPnGAa+8I98bpIDTX2qyzTT5ZS
bDg+2xZq65vkK94S/xAG5YnNaIxMPYL3sBGehyVBxIbMufRvgNr93jAgkJKATKurId6qTO95bjB3
iRca3ebxfrV+StcoKXk6VsoTpZd4qyDymEWVIeX8lRBq80wmu7cILZOEarZ/xh2R/iK/A1zlSh+K
XCaGVeu4W13O7b1aeL8BbMz6qaitZONx3eEM3+vVIsBOVPH6LAC5briQeyFCZrg2tKv99uiODMw5
ozn4Ajk1AD9QL/jTMJs25q9PIQjC3+TgcGuGoJ2F9QP68Jv5AEth5s/oCpPkyTPhnTkTj3TPuUwd
GRPUx4ZUIJUPm9a++w0yAzV77nzrKFNC+7YMM3KFYD5EMeka0QtWX8uRVm51ztAxiq8C+bwKZLYO
LmMB7nfAeUb3rmpnX8tAqR0e/son8kyA/NlMkMGXW/kwJkSb388VWXYVh8v3UgsPG2NSaDoSCuSs
qrsgrtjPl/sqqj9bz7tAucNgXhHz+OIwQvHLMCZvzkOfgpnJX79DR6iFcVcFo7UBUjBc7ukLFZcN
KpalDF60+3mbboUjjUqO34bXEJv1rFxb1qqtGt9I9Il+itrZcDMpePMXAy5xbiQ48jUZjAp7uh2n
sjJ9yRs6Z/3Ry10jLJJV/EgOxJ5DS4mcr8I91/elQ3Rwmrj2GBhPu9IGIhzKH1GSlMl2gYVebYEF
WPVQeXAgJRTxI3z4GHUOjFX4Z3xGNZOso7fIR1LNBsupmWGXWHODE2LAWt63h4RdsPKPrw3cRlAk
76jmp0XvuvUyj9E8+NvTGMSoGvUsRG+hMTS1OwNsKVg808D7+MwYcy5bUCU+gViyYsXc+LkenWTR
ox8tvDH0J6V8D6J/hu2MJzRUlIPGoyLWFSSr0i3EoOliphvbOajas+6aOV4oJ3RePL5YONrd32d/
HzaOntMWQylLjXC9Yi2MejDoizdQ5q+XVtizoeWMCnFKgPVTX+Cbto8KTcRZTPHOUSj3M9KmPv9i
am4Lb+VYPhfpRnwohCTGZ0QTKZTnrvDBBBiHJgT5n46ilgP4HXZoiCfq8A6jMca7C8/aPMbhmCoo
rtpyX4GmXpOxCOD3j8kfJSJrjIvC0q8NrE6pzbBpFP4cI9DLE4axJZOBQVi/LwWaj7k+2Tnml+6/
mOte0e8GBncB/gujMp7q28yNwLrVr/hk/6YTRAwE2cEYPC/QM2l/NJzdbZ07+l8EMs3xOsjeR3kg
sYi0KTgXS/x4irASqlV9c0t23M9m6XzVbN3STVnYSV9Q7H8MnQTus0qFhXx7g57cHL5Z1YxpUhBs
aokh6Xkn45iRP5Jq2O0f+SfyFTgpGv3OjGGQJltr9PZ4AVj3cu8JMYe9ejeYZ4MhU0mQ+BjvCJRU
Hbghzvjwh85EcPEzp4sEEQURn1klNUdyrgAzgpETN3LttJ0Pit1UgNxYt9M+P8WgjU1TLJwfqW4l
YhGqHZLsE7gvI4dupdbV8xbB230/Iz+wjk4N7s/5ZNvkS+I930+NJ5LAzl3fh8IWb8k7DO4+x5GR
yn/9HOWsDmYhHVH4YqHDuO0dCseusfI1bpVaZx1wrkXcREI9V5RZZpVtq+UD/6RGQorxSZbQ3q/Q
iRr+lthtaQ5dsvUYJdPK3yS8AxVMwEpo/c0IjS4KavHvqG7tuH0W8d2+Dz2iRx61S2h/Lp1/Hdca
hvz0kemU4fAyEUEy4p9HPcMcoSukNfVTfZFiOsUDGOR67ZL/S3CogrJm31I+m9D6YcoTyKFRneTQ
r53Nei3pIEaNEemrtQxfR0qgK1AhunHZLs93ZEn7TcDukqmf8f1GuSeVyUmP4ydq573XlCLPenN1
HAqm7GkV7lm5G50npFtdtqWqBNh5iNVWniVG1TloFI4FYx0u83oks4J/yhQdO2wsh0wxOkNa0ITA
D7AChOxDelnJXvixk7uRWW9jzNnrIXpmpaPlbt5cosJcTxhpEBqts1EydhtuGN5i2nmB7NCYFLH7
PEKy5e9IPFXW/QFn+fyN2/P7rixeqAt+EtCXi0j10H90JW9xl6f6Hglx5NtIKNZdPjnf421tcLRc
cXdu+lu05rUWiGHLqkOaf7GRMf2mE/Xb4/in5C+YiAE9VyUYlz6TnFm24WjbILCnPdyRitBuZTJd
EghwOxS9/TkHtDCAi2AR1HMtdbM4tCyBQDwoTQECr+oYiUXm3ECRHWOWUxuabyxn4QJNHyh9s7LH
hQ2lKyQqq152UW7jRhrKAKj9/+e3Xhygdx/UKFaCCjrPoShxmU7rgkO7wntBfEhQoLUmxe90PM4u
boc3a3oLVXsRKBG8tZ1aDb0pWXqKDBK6jBqUQvwwqHseR9guK1HOS+SEyMhfoFEq7m/Kjrs2HNEr
y7TdYbPL2iTtzImNJY3yM/cdqyhVC3NCIKEpKkUjZS0ykJ5gCa6CAHTObAacEJ2PVHXBHh3Fn9OK
uPiLcwVjLUJC4s0BN5vfmjt/UisNViAyiDEjTk+ka2wyZyh7nB/cPCHGeLgaOBf+MGnXDADxpHrn
JZBh7Iq7jzdaYELaQc6jfh4vU2ZtLAv08uU5kEx1UIdkHIt/mTy0sxY+twxd6MGH4LCJk8HvRnSP
89H3kBP6w35BUfYR3fVkw894pPOgH2BHO8pPH519qAeJS02f4WAtKkZf0hB0ZFWZrIL6lQcWNXa4
rMIJIF7VIfzgQUsBrgRMSylWQtdAijtKexVqMTwhHx/rBNDtFa0BV79BAYvV3nDlXmrKV89iY86n
HN2jynxeuFJugXloIgujs63/IQyFYzDFDLbZdLhrQ7zANRi+lZXB/9dpmRJBwj1QaGxR1xi6LDvH
OTe2GIUUQJEA6j2CfswihRHW22r9eKJ6QtbyYTLe0dHMmrCoUQLn2Nn2DmfZPKojcH/RJSiMyNCx
2+Sy3MmeIHvSlfX4rBNfB2I6F6SbAnn0cAGkNlbRWJdlhDw4kl35JXr/wekGGPmQv8/6Ci8y+Y6v
OxRJxwhA7gLvPW/tdgfglGuUQZdB1alZCOXcPeEsiHOMOgIxJHXY2KrBFNTivuchM7h3UMKAJ1hv
584AQ1KbXpfvjD3LlcBDTSXZFX6EWhk3ii1J8zZXy8j0krNZ2vfx41Jo1JyywDfAYsgEpeOSxNiS
YX7QAnjdfXpnDj1n2APEsJpBvk6ADMkL5b4W6abl5wqC8mL7+Fws78h3LlJEo18Rb6dUuhuuI3r2
4zyagpu6y6EUG5WHBaDBNPbLBkk55a1EFaC61VANW1Jg9WJgBvc3egzmBVkvqTZC7Q1kXb0ufMhx
atR+QpumRhH4BRdsC9FXTNItvmiIIorvXMOJ7RxjyOyRnmgsb0Jx7IJ4YSWj/VbU2QhDTwiSCJor
6wJs3vrLAZTA7CF2z2H5nCWI4YUwwsLBZJuz1EQemH1+wT2vSjJrC0HMd0QQ5Oqib79tJKhsZ7UB
FkTcRTTeiTLXGNFdNmT1TUG2uTGvZUJiYaM5YgQqFqzPNLn3t9ESbDWCc48QVggNjNCHe/1AxJGJ
eDRSBkwbjaGKPUF6aoYkRxfF/j8Ls2tU8p1wa5GLxUIkgl0fWFFxFjCetgaiwOymJoj96gJaxjZ9
EssZgXM2VA6Z+ROMYq8b5ypKP3pHOsokq1cr5KORtvij1gtC/hkQr4ngNI6MXW9utA7xV+Hu4p8e
5LEs0peemyIpVNbb2R4JuN7//bJNuLgTyuOJou3bGl9yjbfCf37hlNESkrLyGK9zyLsB22pyakW1
2e29lxS4wCuh3rCTaNxmMwhxqZ7XCNb425TorNLqa7WLlq3Mi4wpLaM9HHADS9ewIsj55wpj4/Cm
y672XZ1kIq65YTipqJNTmW7FUC4kvUoO61tZvzRuiww44oxRb8Y1CJR6IPn4zGJJlJGQP0WRYEj9
u6HuaabKS04bf3ayjCYpPwpLASnxzVWPeZTp5J65IGReKkIMdy9zUupmpgCAQ/Hw0yMEM5/N9OZC
+Y7BAm5eFfzOq03DGgoQrVc/JUYwPntJbm0z9PkI/NWbY6q/UqS/TmIZPK3AIIWUNopWFnJv0fGN
1GCbBCZQraURlIgq6pEGSNGq3ZQgTa6aZdvebRcavr3OVi3jlu7zRXaeivvESWfvEfqSYuaxRnwS
X/lhXeJxq/alA+UxJLYHbG1oSMNVn8tkdTntEcAbFnzKJCU3MicHxtkTVMIud1awZRCbbnwQ2EgR
t18Dn5yyPhdyHbtlOphsjnaksUuMeMPKkmO3bz8N2HgxnuEtUrnMn2nFSlcmRypEM9sXNyZE3FPs
viYiYjtwH9sIyX92CcRt1BwdR9LgrhRdMp3DTLNO2Fh9XkzxD2JRsHekE3cQQDp3AH2AEieaZEBL
+mEf9TkV5kvIFfU7EtbdHXkIS0wJJxq9zXxiok08UQ/D6NEAhpUtfTjYs2pTPzWAvxaHPD0DXDS1
560oFmOVwQW02cJVMvIPi5rqZQJe2GbCZkUrOV7DdkbAZ5mXw3Iu3ug0XgWDi4T5BhLuJSBss77b
hG933gQhuV+H1V0SZmhLiPsLz2dgzMTaIUdyQ/Bj+Q8p9fV8SUfBBgBhbd8AlquTWaXkxCudc/V3
Zz/VXpYz49A1va7zhWlNzleYDry4np7vdFIgSjOtf0RyZIInqz7C45EpPSv7lSj3F4yJ2EykCFIh
daYiRmx+H/wE67dFqdzPc12OYiD4npesYYo6WFNtpYK08OwGFGHfCMm5+3k8w5RxkQOGu/1UOt0Z
sMkwkTOZ3qBxmn+pU35DfeeIXvZLYnwQsQ6HTAkV9gzVMgEhTYHwqzvXt322K2IDUFQdrtVtCIln
btgDSklMUIMaWecpTTImH3KdkfNrTZ14eQPxTeoO7dYt7TKZaljdxDryxN/EtCj1lwT1m6sMBXxK
UUB2yHoO/xfgaqEnGLH+v68LugMAHBbMb9B7ZqN8GNifBC8UWLDhFs7K3IJSkQDbfoq0NA/cA5H5
gao0EMeGbXPJ7k4sabQrCVuphazSfrVpJU/fn1g6PPTG3RGF8AZml11mAF8q8DAQid/hYEyY4vyG
8C4xF36xwK27gRQe2N2NDQpfzYFDsoeqSXc9X3tZTuVT7ZPm+3QIpaPi3mZQpGE4pjM9KQ8GVXs8
fQN+w9YaMaLOG+Tm5ckzXS8hr+Gz/IGQ8bp3IC7a789gIoBNB4qIYzuh4W3anHL2hebLa8dqacdU
q+urOK86st/9nb7Bl/Rtp+NAdt7J/V7MFEky5EFwsvB/DXTqWT9cy9e9aKFwRrx9QWBfxm23DGVb
bJT+CJ693hG7J1tOS3sUWb6axUfsZtQTIVOA82sZndGIfqVQyXY8M7ZirU1sRHAUcMhq08FqIvTO
tmSRuKcp68YfYj52SY2W2AUE1bienueuiftBuo+oRefXHh65iKxpWSW+09WQVeEX6/YgecDpM4T8
aAoQoWyge3GtNI/6e3XzvkOjThYUB3KPegqE5faxKF6AFX8PbWONBU8aujwKfYtkqN+QKk8KoS3W
7tO+3dJg+Kd0jb1ufCT7/DJHPN5LQcz1ZP+fEoueTCSn+0cRZiLqMzaSCmWPiGUFoZRyhdsCFHOe
L9582wcPI4jL1Xeymm+GIbTThoUUW24xWcPbgOnHlO6NnbPPOIIxt35tiX2ityvvg06ReN0XLvHf
85GFnzrslkAAsa5rtzrBcuOf+5EECIChDzyMuWZ1AuA3PXfOOY7GbJhiqqplTV/CcxBbBr+nQCbi
eY+TvO3sDemJibdDhDTXX6zzQh6Oxwpjjc8uljSCwJAQI3kDq1wqXzNUxHJYe6oRDx/BRI/JZbPd
4dAFCC+Ae5P1nujKBDZheEBq2tNTBtUsxEe2BIEALSwccHV9lKCKQcLrXwa1llcxgGtFj8ebVNax
CWWhO+liJykH0oYiBkF9NnRrmA5GJZcebPood7PA0tZO/wcYXHJTON14ivoentxKWpX20PlBAxkB
jTalqUbE2WGt45AowlovFp8v5UB9gG9/TLjteeLbGSqHxooELJC8wGxfDYcybEonYhGB/XUcNXHn
g+neofgml3PmWzZJxhNKTgdR+4cw6ka5cWNAu6r56mfe4Vb3fjvrFL/D0j8djYC9QMXPxtblXN9I
iwV3GTfMRJtvYDJoVu/iu6GJS6Ayv1IwbgxNQzLWjMwGuZbkV9XpE0gr7C2bY7IsZHCoux3wcTE6
6DuUWvfOEpttP18Hncic+oCwrNxBh1/uY1OwXZ6wWNNkU9QOWosnNS43RbOhviWXMuUM5s/JbeiU
IxBIUTEvSEwSFoQOTchbe20ymKJx9cZeB7PhBSdpeBZzdISSbFtXF/gHwqN0/3eesXoG981nd/sZ
NiG9bCChXfMmgC6XUDHNaxUR350Gs6w8T5mySU1Fpro5tYHqrelzDbPeaC1MDyMzcW5z61O6tEBI
qG/Rzh3q4qkfR+1LLYkyDXjvtPhBdmF9RDegDbpDQvAwV+T6ULwVXskSj+/+gPTkndaKHgMDPudX
wdahUbio1YWlzVZJeOuYQxImRymiz3u5C90TjODd+FqWXOuqH2kYd7A7Z9fTt1gv511259HLq4vY
bPLGdXGqnBvVbmrfWb6hVSMwzcK3afU/FaEbRq/dKImnTaG6tUNttsHchEX7/mOr57qygocEqwIe
lqCY67AUiIXQF1ba2sfd4BFrrxQtNGlmCpdu7wO9P/EbvHBjlKi+gGJZt4S/GPrsHkJ9iZ4ONmBm
Q0V+8zGhQwy0ylS+5DHQeETO13xi6uNqg+WS/z35HSu27OVTggOy26E18xaYXI/7AWZ1Aq0GBAF2
8N0M3bwCz0ysnq6FronT7O48n9vNppfmHykAzEkhRV4LCPqn+KdicEG6GZ/3humUWp5QxdBuKfxc
c6uUJr7H8xH3hPiCv24GuuEa5RtBNycHp3rVvhPb9rAk13tQWikgVaYAqHxq714TCEYI9cJTwkcA
naMTywhd83bSAqLo9JcrzNUiGUu+ezZlhUN/M1/0QjQhZTM8TCYZfdV5EjKHx6eTxLSN60uzvWDK
4kXAHpaH/DC3vkMR0ikJ8kjhLm02Of25H572pXQhjGCNPM9gDoTF5/yvUCTUzwClGTqLgwUyJ/O7
an/Lxt79hLp37MVbzn6IM6RSRERfDHPl/hHoCX22Y8U5Z1no82VXCQY/yCCG1t4hJIOnH7sUdliB
Scw78EN8vjXs00+wlVHpmS4s9jWoK8nsMtrKFcssSJ4fETxg/BxuLeQ5stuLDxMxbzZdN150hxZt
KZr9P8MUjM/YQKC9GbIofJp61P3zkxdD3J17Qd6sYXQXGMG6oYv1yCyhy9cbiUQMcSOfm1eBzgGQ
jFZ8rbUUv7jNH+1Ve/pe2zSLkanp57/Vpxran8w0B3PUmr77D/ejPFQ8o9KvKWNInI6uTfmG9w9Q
N6zYjK8+W18TvEKJTNozsja5/+EjhBUoNBVbtEJ8dlM1wyVt02Wt/4dOrUAJs5wimIZWlEf9gG5R
EUuhcw+g+Ps9R2LjSx6TYreNhhPc96MYhfmjhNM+j1rtZoRNOlEy0weCtbBv2XkCHKGRv5xUpuBH
Do22+A1mhDpD3SXx8VluYsDLRmnjWqVfovRPz8/gKVzafSMyykLQig3duW8stlK9gSJt53A1RM8v
wvcD5J4meNng7xft1dzSK7F++2DnyxlUNzzJQwQ1fYN1MZDXViMUa6ODYmgGGBiiAC+AgNmZO9wn
2ga3V1rSG4ADKoB1It1RetKSrQEIm9X6Rqw5w5oxZKmX2BGznmQ0qXZKVHyXlkOxZh3rsmBkDc6F
hH5AezYeAmhRBDWJHUmwMlO+nyr2LDdT7p3d5AlkwBWTpTfuCAqv2nRog0NRJ36Rg0eBH7VLdgpi
bLCVMudAvIoUEN/JpH/mkNEr3cHiixI3zxKh5FUE6RDU9FYDI7KJeqt6wSPFZF/Ci8SIjimjrV/Y
5eRITUsgJyH+HxpzjPOPJ9VaUERrHhssY7OeUsitKHwl6vxq1PJiB+0e2mNhtV4y7k2nRn4k014l
D97CC/muQdkpeLvLG1WNf8Yt8EmDuK1cOXvqsqtro75b7ZVEAMcY2GkPCBJzLI4P1jzWPpISBHVU
q0RBFudyld2SKKyBtJ66othGi6XI5nStMFegXsHFomTi0TbX1n3cPw4CZUF/FMFaA0h8g+ZftN++
ykLVu+lxQU1ndvlIXohMUjboeHXOR0E33s4KXMJwBr438BNSyfny93VL9Zmm1JwUI+qFv5oAt10O
cKcYPAwSBGl2/pYe3IKMj2nYbZBU2rdOem8JdEIv53KOGVHKaRpnJrCIE9wcvq24jkAUN/RNfqoC
6yGa6XdRmxr+sbNmzEzrH12FgsrLaD6E53nFw9Myp7mfN17bno6F8HmJ9TNCajp59mskiP00swGt
Vkz1zqx0giweL0papMEMhWlSZFQKvsxsyH5hYMgxGiw+Dx61ZdOlW685yUxNOJbGvHeOEdY4Y0t+
QTndJ3ms2RvGiIzF+Ze/b2pGrJiS7Yugm7QYLeNKPXa5tBO+c+8kSo9TsEOvZn+EqjKX/H4l3qxf
3Wq8hrz6IZJHk5M3JZenb648zutmwy7z6jt74LoWRlc7TVyK+UGNbq7F1DQqgU+h8dLE91Z5Osph
xlSM7xHpErMS1h+Jl+Q/Z27V8s5mytsdJ8dwDmv/xzNg5wq3O9k4p7VXxL0O/tfdF1JoW9eV6Hoq
qF36qGEwcJCS2bk34m/IX4hEXIzIXEyI0RQWz8w45hFj9gqP8eHSDLha366eQOwo9BiPxpqQMUYb
475SC+w051Ig0nsf0r2PsbTqsHfB57+jBSaiy/348tnf04bkc0wHHsBFq7v7CuKiukHp9TqWgdtM
xVezl8zgDO94PIQZ4KMI3ZVWuxhS13tfEXDykr1WwvwOGPUQiTKOx9j+pKPTU0mLaHIakB9Laq9c
Tpkkf+J3LFyTBFWbUFqKtMIY9eo2JXvzaAiOWmkZF3NaRHfHEQyiop/xTw4fwY2X4OHQPOzvIDci
LibOrGI1HdXIG3vx+FVpa0YxdD3ZNplH8WGVD5z5HLd0oyPL1uv6jgEB1eR+hU50fsU6RbB55q7a
wEmcVFEXpWOp5gnvMW9+aDnfbym7LWnXpM+ELxZ0G8H4nQr9shO+EzTJwGHn5bK51eSW9g8iCDiw
cFa2dOcoKEuKQL4X4PtR5bmeBJ1zbcwBADGd/GJARIiBfaUYmLfBw0WDj2trKuim8VDS8HxFepv/
3NEcfobstdDobblNDIG7mTCitCDylb5e6W8LljbqRc/4sDkJoyMWBHczhG8Jou4pERQ3tgOAoKpB
1m6ts99r3g0cXGiWKnzqvByhNNSTlxvw5fnTlXHaM5EA4CxS+68H+sbWSKbNcsBSAm6z+Z7FOm1U
Pz2FpCEJc20RNtj+YlVWc60LWwEVB8z7rt+4tAS4g+1/yHWTLj5AaRr8MA92xAX9xqZKzycuY4F9
ELHPR10YBYRE38L6Rrzu9R9wJ9tAnvjvxF0cd49fgKro3ewDSXk2oMKqAfIfSzE6kOSPXLvTZ994
Tsjwpb0WT4Kthvj3QjeQBT4aY4SHVCt7+1QVi/mxzkKG/Sqrbr6sbwfr1oivFFgCzVVJGcqbNvG+
XVbzD6koNYLsvGI4eTkS7l0uRh/8h7DXi8JeUFNKdxwRVNGksQl+iM9MouU8u1oI/hqPVHM5HeU0
mX7pQJup/TArESOmRubDNy+CTNtEyMc8YH5/YY55/MYL73PKV1T3waMdG+kn82CBvzOsgFbI1kQe
YaH4YE8FQ13YrG43mOqjXCWnwgtEOQq/4xiGgI2vz+dyUohZwM0x9kH3tMHtWxvP+jaY86cKB8+i
7Umw5mgxhN7QgA0xRx/pX/9wx0xVIApw54BN6Gx+kawHVvcfkpqh0jrnaOhqcmYXOen1RXW549gW
HPct0146F9bH05b99PBBYxY2BRaBvR9jxGwgqwq9hQyUy2R4sbSy2qiOZuwhsPFT8iiFTS+cgK3w
Vt6Vpdqa0T+xpM2qpG27Wjg1KHaxq2Jxt26MaN1PstgVWJgOPaurDJ6sJFI5ccP4sNCY6EMB7jhW
jVuC9pFQF6GFoO1DH+srqfzqZUxfovBgAx+DhSqjlC9qa2ZuBdXS1fctrvm/W9fq+doAoHBxheIX
SdcRr48m1K8l+g16h5Fu8kqc0WMbF3IaAGiGDr+dH3D959EwAv+RQrVnpu1BMtZTQqsJ1eBpJ5rP
YGJAldVed1HhpbtSzW0a20+bqQ5En5SVUNcHgonE1YCIx2YgjQxMvbe3/p0/Kc33tN0vz8f5HYYL
vbSbQSaqufFLj3KzqsaYiWMtsEUVASzt2hhPym2wGsR+5Eycm81WJe4LH0FwgIHb7mASz26mfrmj
33TQdlgv+0hSZ4siN7jxeGXn05cA5RVrnMpYUJd7y5herkoNbGu5utA/YO/FURzNyjAjjNtPA2qP
RAW2WstSXiMmZW/sc1cOOM9vCOMH/K/eL9JwZsvcaO/lRcOKtebr8UNmZ0BfP493WEgcjVuvgOUN
OSr/xZPi76MFBivm2C9/oH03hnkkKwJh71kyfabN4DH/THeqZxKyh04nCVmA2IORnW9sFpWD3Yq6
9Z+SYE5uQQdnqQlsfToFNvMqO+GycpX696eCEnJ0I8b29UvvV4SjmRiCYuwMtsH4UglbzdfkbMZb
CmxRyPYqd1W9GGSfEit+WAu3DuAfO6X3LfOjEx77odZOKAXlWHgUE1OD6I9Icikpw+u7JMk7yUfN
A2E3o7TWSpDfIinNnws2mjUzyYm3s9K5hVPBzgia1wYayBLdZgCw1c16I1i3MNbsmLh9gldy42td
jhMdNxPeWn2cniEVLbVPowJ3TAWXGn4VzYxV8UkIoQ0IhR6J5GCoYiktwdTScTbQfmGQGnPxcgcG
fiFgfVt7CgnnAPhm9AqtI1Mt7t/nJwL9jEWeZXPYMAsxboJxhKBUFLlIw5ujU3z9OltDbhaq4SYe
bNL77WoxwncHQi8pB86bYE9tIY7IPef3FIsv3sNrNE4OB9PoOk+frOuVk+W9m7A7kPdm5QBMFs+R
SErhjINstdiqQCjFcxSzumI2qaYo94/YB7hDBPnD+IdfkcJbJfmlpVJzrzxCPTLVew+dD1HpNnP9
x1p6yqdY4OXv65WIMGXFr5X8/UKedhQKALFWUh+qUSNKFSBR3iUNORzWFvcEw+qYfah795wmkBaG
LQczHumRxQvaFjwqpE+n6sx2fvEgODDSWZRZAFeLn9KpFqBu82L4Yceab99xZ1JSf501kgjEnZbA
Cq8xL39cufLmg9Bph1MNcDzbq1EF8JOn5ylHZIlVE85AOZadJy+piRX3LUBlnB8aBuH1hm8rZPtD
PjfjeAvnBYSQtJU9bVtZeEvoHUhoL1fYUioTx5P6i6dU3lkaKdfu+AyEhfawQloPZ0m9IWcc3l+o
c0MjvKfoCX/sNTLhgbUhZMWF1pICK1EXWHXv6cuPd2Y7ADk5V5BJIxnlCkLWLOkhXwMENpdoq8se
RIb9A6Dusr43PbcYgaad2B3ggV+sayYSCE6Z93w91NO2AGvLBa+62X1f6mQIDcSE+kxCPZ3GZGGq
TDV28NYnvLSep0kEXMaxzm3AhBWp+Ybs860c8pJNs9XoKzqPl5QQZ6vmcBjwkvqazmDs0McNo0TB
t4rD83fs6jvOO6CVs8pzgue9JDua3mPcwhKBsCaeIkbfEzabYRU6FurefywsVDillWcCfiFWnohS
Zp8jkzO/8TXADEZv5vlAQfUcZcq1108UsNmDBpqyTabdym/HXkn064YLJPBoB2LZNgu5KN3ND8j/
/MaLNI1qr+rJoPMs9IPKUGY14eG6hcH9rrd5r/dxbSk3U/d8+yD+Wx2tVY8tV61sMrbazHIco6Lx
Y057FsYMML4BCgsQ/j2D7l6KuJKfjUG1+I5TfAswO1FoyxYlp9NqLBJ6C5rBuzcfnKw9v8pnTGjh
HNzRqtAC1IyNyrGQUoL7nyK09WllQMukoiLlvKrXFs2aqfK9m+kXLTcYNkywkvf0lixy8lT8+2SN
bBvGYjqEIk+MRedPGg6UVyXT7Qhxu/f6/NZGKgQmqRnEVDMWpKOLU/LPQUs3PsxDBzwDAr0Craq4
KCwKssxfXXpaJN7Cu2ap6j4Bq9j/bWrWEU7pt2e3llk9HjQ7RmPXPyiCIOQaP9QhpbH3L3Pm3aKo
v0e3Wpe8QRJMrj9dnv15Q7m2tbELQ7cuEQPSQ/RJqu6oYfkF2p0fLCEhT9rCi64LGjY6I9O5mu8p
wrrNDNh5yNUFG10fIr2sl9wOR2+x7lycHEz7bY9VEZVPAks7eyYdzdYQHtQ+9OTEsxkMeVd2UTa/
WVSueogG1amFunSZVEMdzCZf8h/R4to06+KuTAswl5pepXhfLcc40IO3qIV2AaQ0rF/C8FHhYn75
vV8NIacFqotXzo9eUynQytP9CsIgcTDQRi6cHlO0Q6NwU7skXVR6VC8NDkwn8ce4bIyb+6SWRv8N
vpeoLW2xhsAqB2+faZPRIUyw0DN/PH5ZWiIYaA6GVrZsJhGmd+UqIkVdEgrrVrSAo025ha4f+bx+
apTjO1YIAv6hhMTtDXhmDKXJX399ZvcDnjozs8XtiwzEyFoPvzDB1zEiQPKrGKYxw62jesc+Fygo
lXbE50nevazMXWpEtcex+XnlcLEfQSXiKzc/ZjerNgqQY8g2r402VkOFLWgsENC8aXLkgOCCfC4L
NczfQfi+TIm0hD8VaOcdCv+P8KCLg0L8djRfmvdxx85zLiL7UXqCxFqMS1h34UW5t+YFyUpFTRbL
WAFBXRDLWifGejXOw5Xw5X8JgD6zKG+HUEnew4KID0mkSXdHK41/KELzyKqsrus53lQ+d60W+3pB
eWEjXFg4rfoU2K5r2L9GDgoMqEoB9OnCUj/IBVliQirXEX5c85Lb0xXnwpyDcFuqW3aw0MqBbZkW
rZ8QnAsDeqMqoRC76Bc6fj8iCKYaH/5yaG9m/W3LAfBpGhyKz8NWtOq6GwjS6xMsKgHIIKLjN3nw
WyoGEK5cBWASRzWIpXMKh/e0uc7v1wXF1P4EKyWDMtfKtVYTrLeubpxdODFKEWQgLksmIh957xSh
To8UFcO4UBe9mW5iLBbfzGrD9qadQZWY4yPP7z6KwX65m99kgRrLJcRTWdXFksvRLpyAWKiGN4xy
eRZq4R36Lh4MZg5ROtzfmwXiDpuJeIawPYsf5e01sdUR8vgG24eGrsOPymcJ98y9XZqXDq2sEyJ1
5ireTw1xtSdjUE9QXKFL6re7Qt21h/K3IJFIE5PxLeiM+K/KTqWA7PWEUz8F16jnfgEDpm0z5rE5
+3Q+XTg9LNfz3UkX1oMXlN0E2z6936WTp+w4st/j8FhnytvkF57VT1WHfSc4dDiooIDid2QKUwcD
ZCOO3Iu5dTUZrYcTCmxpgtLu9IUCdxGSZH2wQqj4FNFtQNEal2uLVAa2YlaFoStii7DksuSlJPcA
LW4oGp/rfmTqjAcEjUJJeY4me6VV0i6WWKrmu5roziXBLBZ24yRyxO4AotL4GKiEzIKMpQeBQvHq
DX0FxJ1BRLUB+wOfbrWRQ9RP9qWid1A1WtdCgJvU36pCK4JZsoNUYRy3MRieQYxjRBuroTzAOESQ
q4GWakJT4IT944XlINFYxnNk/etQKCdxcf3o6MxGdCH8lg3dcMvxoVNjwzsZ4ijdMYa8YVtgNfFv
UXrUkdmaXEL6BnFwd0aGm4be9cJ1sg+pJOJodCEnFkfXVbHY3tHA205dwPy1SD2tFB2IXgMeamDE
ArjhAhiAhmQ2p+H3GBJBlosoYRlNNidiY/N+ZEtdlo5HHBRK1ZulewygcPpHCJn3rOv0mcmWhNVL
o0FhRN6NBp5NQrzr78e5EetvOL5J0hxrslGpUmgnolHMZQC2Jl09MlLomemHDiOprzNKXwgStx2u
PX6P3dLkDfqkKcRwmQtVfKRfMC382ocA+uohXxJAT4R0Kc7VbKK+hkkpIVl1DQdQCAFGEm79Mh5Q
M96Nu8XwPmPAKkx+flKF1MQFGAkX+x4P1K9SMFvxDKRsSD169rO7qH5xnW9nu5U01AH9XaCP1KRW
lW0Ms1KzT1Xcv/EvcJBt+QlNncjbwrc7hgVh3kgjzvaa7JKzlWYSq6BtdR3+O9gGq89Ccr1sG2w4
Yr1HimJFPn5IqXDOZlm+QDcaeYEaG9z/S2gUHcYN2rkgNTdfFxID/WPws5ceDs5u40Y76pc9Cw+V
HOIN+iydKvlqjw6gESRPqknXkV9u9OWFidF8PVU+QGdJshsaKNid6pWrpCTWhMnyAe5HcxgLNJdl
XwNaUpIl+/BPfv8T559pMRk8k/JDMABB1+w5DJoUdHWiSzFWSC90VN7yRwpUqR5jLm+aQQ0PkPEb
2nd6m3XNSgVGkSgnSJ/W+nalQwCd0tTGjp2uWno7NnL0OYMd3eWL4AnGQ+J9i1avZLEOjGiFRkHZ
e+/4Yob8hw/4AgRGRv6hVSIEvUyoYI2dHqm1wtewSd1D+orkYvTAUsr/dE3eWVNWJP/Iw2eUxFlO
CW5wfDiCBpQ8+baU/kEj4PuNPXDCTMmcVqBlLNVEC6wZC6FSdqnr9UTayiqYS1qjVNy4TTf/plq5
nmYyiaR9FAf5KvYvJwowXy1j/dUBmwClbofPPe3EO/pTodM5F6EwAYPzPBHyLSXB6xO7nx58faKv
yIciMV73jU/12EiTTYTawyINLqv1rer0/Kz2ylCCzeIC/3oPvC2gkuFaEeIdK97rsop73eYs6Af1
eCXaDzrAS2R0GVFHd1+SSefVbLPSMkSmRzb2kGkj0R/6hzhPXdAwt/6nXlZnXJeosSASmEUS4NWq
fYLvAXfAmufoTWaYSba7KETFU35K8ZQ5BbsUJAnU/bNEBTPnbxtQIZDX1q/JaxEIeGjaHHZkMPKU
McS/n+5fxOAehMrVezcYRu35XUcJubwXpH+51v92QYque4KIpcRp8PgQpUo3kpJkUrWS3fX2F9Ho
+cjogX+kECipjsuXtIgEzDmcgsVUYWJ2DRoJWLIokkD/XgM/CsHYyr3cEmGLUhQs82rQ9464Sibd
PDmUnX7XtKMjHxeQ7nHOuOYgox0MstsC3chxZ4xnzb+qvwwShcbWau4tV1QW0noRcHtq7IpqsmrN
3ITNwSmiV2Z8qzv+i0AD5WyR2WJkAl9+OGs4VPWixvCUNsh/u404lmlFWhbQWzGz0eoGmSPuNWCo
Ul2PKOcRRVDbA/Nh6ExjfmQxNeJP4hj6bWkITEMgk4Zqvkes48JCYGDv/oAnmXyvz9dI4LZorhS1
cIxDHig896o2HLORBY4sGCiVWAowGdFPCoTws6AhWjtyPVYzI2aC/Q6XpZhQfIGpzBOaoOS0dOAE
LCWcqdZz563tTStP42fPetrkbay42xmzBSj4GfK/Y6uC7eGwjhqCisF7WNaYiaw6ROodgJn0+Noe
5EfjbSj+LODWwPwCw00J+ttt8U2q0bwGzT6gEGEovFbhy8R7oib7rvf83Eb1sGxPQvZde4sF2ltt
D7KV0sOM1CeUxrZE/B7CpCnxjriKnWKI+sH+w20REGtEkZkhwnUNHjGOElG4ITebb7HFPXlxXg3y
fj2Obprc+tniiyESEf3mYVJsOn9h1Y8riu7EubhGdGfh9jOcz5NhbHtjbu9pGlVQoxBPrvlf3nQz
WpPrZ6qwsQsfPwEVjOZwxRyvVSNv436I2KI9NM5vj7ChE5ShgSYD3Qc2d9D4KJVcXL3tLv1MkarQ
GR2Mp+mtMRmN0kIjQrC7VAQUx8KCxdymRAaHoCop/cTtGu85XOOPwriA083e92aUQjDquUhA7LiP
a+X7ogEeIqmiODCDqspiutT5AAZGIKx7nCyoH3mZ1ptizyf1Fh7KmDIvv+IyIg1PJgatamfqX4AD
PwhM8hYDv5LpC733d7G7cgvkaH3Z2TIKO7jSFQg9XBL5PW54t0Qwahb9qo2qfQPpjjNV45Et7k24
pOWNAIuaiAvtx+AlyJtCOuVLsk/ZZHuxzAu7uVoFcbyr+h3Co9MYTEAEBRB2zXxaewVQBNpm+Ean
8KTT39FPlp7Yo5ksLcoDGyUwxWq1KVoUeeSn5psF8HETWoEbeCLrPAVr62pgMrZYS/WXnqiXMhY9
zwmwNNfFcNjiJgU74UcwAJgtpmhtCTVbayvczLO8a7LVznwZzrkTslZsUUwyke753SIjlJ6gPF6I
OEJ0LHTyVStnsi5ZlTuSaHaxeLUtnvyYS+/2HWsjgjaUCRGPHKuVL+87SQHNrR+C54f2dQKOtPey
udLaypUo8fjF/Ia4ZttRMACCx+3uw4x++arXuyr71eMT5FtyxLOAxXXkITW16/pGz1fFj0gJhAzn
/sBkfWeEX8GnpgI1u5WgfyLKdcdEfSYmsB48rdkJW9BJYFhs0E0ViGl/yECTEVyvtSkqBMCn6PoD
kh3APjbnQ44Il7bekzM9hhkAWJElaVC43+iR583xVNrph2htqEx8L/jC7Fyyjmp3FSGKpUWtNDqz
SjLv9thF3UDntxj5dMkpkOkKuQ3suY0BgV8SU47BD+j+47tklcLy3JiD8DFL3LTL+3zeYUxIQ8t0
+J9tb/UbcaWfGYSxLmbM6nYO0PP0aPu2IdwPiXf6Hw3mREewKlrz0/YGBeG2OGXdgYdH/tb5RcVq
IkEVCmecjMy05ciaOXOpLIWta6EmOADISn3IOda2EJowP6vNzEpjWGj+8KP5YuIFIxkXJzWlaoCj
8QRa8nsRnkKwCL68ScsrHWUCgYSBwfylT0K5mwNiOL0RMs99wuIxB+3JHp5BymhP9cLNZv2LjP3/
BLY/gT2eqxvN2/ZYeM0zDNHtdfH0iXPjrOgdlg7aTeyub14zaQDvTFjBiMlGcAJttMnhfEUzdMvf
CArFHtkmPqo6qudVJnv09Py/yPBofXiuL/A0nyDItcUon5jN9yoOFTF85vD3RtO4WwPzfBm9di9q
RE5Ap+s2giPp0fQFccgC+1t0lJpyGle2w5N5y7EzNdUrsPMeVTAFzOIHugnVYCQXzK+6xbhqLQ9u
L+mvRS1gogxwkVqB8D+UohHtWbLWdy0641rdEQnQa47OhWNLc5PwrMX1jXEu8yj9PFQ/XlWXdIpt
xzrZ1ir2C3CRqVWW+4tHbzCk7vbGEXlnHMynhXbSXmpS5e63MRjlJ9+N2Bwyq0Ck6JMNpp4NwLjJ
P1oBNm3jFF9tY3utdqtV8uQsQnb/ymHTQ9e/okOSuwpSKraVbpapp/z/1sYDnNHbifmLebe+IutI
f5Km2133emrDcVHRRJX1IgKVwjU4DFIQTJzDt98Mzy8rfeFribAelJBwzDJ8ErwLbAjNAITLfyTm
kdCKSaL3UaWpRQCOdWjKHZ4j3ZjKtaiLGQx76pEol33xJqeF6HtswFLJGgDHc4TLBVv1ik/O5ltN
q7JSU7ZQkKKlIx31ENuEilCUEm9q2OG//zTpYFPjGdhjCHabRMpAwS5lIvupfhJib8b6NY0jY8q/
MOJ6XknsBdR14zqUs2EHTPqVhp0bv6Atz/Kw7fRV02q97/RaCxRb2w602qmTCUxXVny7OEM4/Sge
KIIAUokuM7iEJo4azC+sNaqMnzCwCcI148lYKYYqsFo5/QhLMANv0ASxysA72i2NyUKE2qo9P28v
rFqWeFHzUk3nifvLLi0zYDXpOMXkQPays72I9WFmu+u0SkHOpuDviYnFOUIIqffNeDSNsVVsXuCP
9GikwH2mhFYm9dEeWEh+q/8aQuPT1zx/VS0EZGP9RsGVhzg4yTYtgLky9xcqKK+YSlsxnkTHg7rk
MAw5X/SWfb74YmBNlifw+mHMwbV5K7znGuhIAbDJVb7JQoUQAFgMCXZdD+HmEpRMf1cop+mVmrjo
k39cbrl4h2njyjOI//k67EcyYCbgQPx894muXL3hCsYr1A/0q29zNq0HPyMiRtZJGDWA6lquCKUp
Ri/vMEvXXhBsVwy1SX6K+I5EKGOW9WIUBDU9GBFd13Yo/iutncYA3YSAGO7Z3bhkB3l3VdDcVZFT
3BhozroZl6G7WzOx88DdFZDcROdzgAN3kkqV4EJXh9b5t3BW5xUYssIcm7gKta2xHvbf9RFXs8rW
CGXKumgbeEyzoMZ7uqmoGHsb67WVEQbf4cYABqVf4LKpjRfkZMKITE0ocNLD4SS3aTcMPT13R+Ul
DYrG3obqfQMzo3W7mEoPqIn69++59ch1IL1vEu5IE2nGGsLy9Nh3NfLmmZhxwld3FIvlWtuHZb+o
UipMYG6RN+yoTEdtETgec9l4o2FPkng7ygMMeQkG8BMWl1mDzKCLgfTogolyACr4CZUiF+6KzSuw
lIJ/Qb19kvtlj/nOBM/lO8Abqm2NbgS2hK3dqgUTZaxyvfJNZur7CUf9r2r/BcoC+MogGjWEVclS
MHMvSI6ZDbX1RaXlrP4Om6uo0Tq9oTKirwSjhXCdj4hktHjN8MUrchFFMure/6MMF3QRaPS+IOPM
RoE8nrcdnn0klFxzRiIYvd5QdT2D1+Hr8OhDGjGD+8br15ycO6eUxJfiOAW33jM0QcyipaX3tEdO
utn3qwHD93xNjAqaK09cPL6lUqr/5E24GQdoApxGbLFqA9g1UtEeS+gqYPs6qqpgUgAQf+FvoTru
U1ojJyOke8/WoooMcYTqJlgxtq2rnG3e3+UvLPwdVojOPC/k3+EpV9mC3oD8tAyIrz8hmuCQNL95
uAtx9HuVcIFtFbCtNlAbAm8gaRqZnpJR0/chxuiX/0vF6RyJbByj0s1pT0MC3phn4fy9Zno//OYI
/JNJC3Av9hFafagtjRxCKSp2IB5KadLzQzIf6QYpsr2tsPEX1uyn2GQi3TAFYej4N3W7sjwzdFT0
aFtflW8FdS6LJ5CG7ohzBZAcFOWSEQa3lFrwZ/DW0Ssu0LLU9eV92lVA/ebsLuaKCf8KIFbm9e6l
XmNVnEhLs4foFazgnOqg2Y9Fx9k5PrH5X9kMKEwWOSVZ6r1FZ+7fbEhotlMa+SoOlriAW+J0iyst
sQR5ZpqzfyRUHm/UuPta0mlT8+HokrT9AyEuDPmPOL1yDYN75tngrihm3QU3HkcAvnaJKZYMIr/1
RzYHBR/2STXrIVATm0rNmJS05kxRncxoebOkpzYvcIWqJecoHknlucarmX1+CqFiO7Ooyx8izoqH
0LvVowcQcjHWcVs7ukmfE5YjB/V6k6vazuruA793cfTcZT+G7X5GzFYaBQrcbU3RYQwWxyPNk6U1
nNRZ0f1NFmoGd0Wus9LRAh1O2R359nn7zMYctS39/3bf1yv7gceIx3WzHRZXy+q7HqWT6gXIHzNo
EljGvlXO+UdldVEOr2bUe7IwNqbRyObL56bJF/AWPxdgoIvP7SZ/vTQEHDA8olxLlvy4XTOgUJqK
m1M1uvZc4d8R0ZLiT9/eN9M9VPn33POJ/T1DkiTC3O2Ufjpej+l9XMOgyXADMfJr3eXvbgd4xLwQ
tRjbxYOKdV3PZUZHm8q1eGgwAa+RI+RGt+BwrB5DPZAVeZmp8RXg3EBgd/CR3bgrP/ndj4H7MhnK
b6NPblESLeWet72fQja+DvrxeFJr/X6YUYagL3AJLPuMazlSN+CDaKny0ZyVJWNyj65xZzM2j1bt
KPX9/bNGqNSmFCxBzo22AFeixrhUJeDa96T/hLVA+gT6zsUJ1s/zHQ1QtHXLfIgH0XHdmlBDJm/w
1oGLRkEmV91+TplQvuJA0Xzu8R6+TrSv7jllTJAIfCUC/pJ1PlMe0ii7jbKgvYqeXSTJUgnftn0a
/vhz0XetDUtUagTGg0IEPBzrIpnNsCh8F16Reevg9XQMqim7v7Uz+8V7BU0EUwqTCBDWEZwdxDFX
0auZNA9wqfgjqTsTb4+FGvrw9P40M+OH8FhLJhQf5U+mLxt2Y3RMD3+pD31PVbgvtM8zbgZ2T7jW
iHDOOXiGsPLRCYad5bz3gL+2a8Xry8m8UOdpmefAKTmZcqCc151nOxXmlZHuX4dDSWetS+8XQgCV
MVOmbeuB0WqiiFG4jOEMBl4vRzYFX6VIbssI11xTO4xTt4dYuFW0d+wJtUAH9oUNUUWKOLpMzqRV
vhfM0emtuVL3IODzINq+it6zI5/gk9eUVhkXUNEBxR4DEBAjvCPB7wDRdE57BHFzTwErDRbf1QF1
Fc4ia9xKv3NnPeIYbMd2EO7LFdnAsMDlx9qLies/rzSqqy+mA28M4eJ5aFsXjtAMHZUQuuc6SCNa
991zqyduwhkvWlcXHcxxQbbwUA/vHDsQcKUmdlq68eQzqeuFRg/aqZVjg2IQE65xs+aA664GLiuk
ejYeNeFnm3zqQ/7wgjWpaqk3es6P8tI/tHiKAY03tq65seKIO7a0WjbSra8Y5427jVY+WgFY5xvc
znlB6F21PmjL5uhd2z9tDZMpXJ7SajtQigSwS8B/pyeqyCV/8kyB7MbKnaB2onnBKOwPGXMgZZv2
uzIomRiW6rNtgg9856srCo9eUBR7+tGWqfJ1jUIpVMWS7Ni6whRSJ9nMfktliOD3ln7e6j1M6xT3
wHRfJvNWM/dARg+KGvn8+kGOMOs1RvSFb+E6qqNAHmWNodoG0owG4G9XrTK11oIvlaHh3iuqfjyo
I98LoIZpAFIM1NfH7FdS0CWrxtlZAFirfliKOksfoCy/qX3mNF60ZlIbAKmN2KakGTeXVDnaTVDv
VH+N/NKcsLn0EOF/x87iXU58ix/kEd+HwbxmkDbh57puNljcN8PK1VPuxFiWFWSbK04LAcIHF5A4
NJ98lxsaouUIZsT5KruEIhBl7ISR2hmVPmacJgowaC6XVASRBe0pSHsl2Mu815pIaUotn9HelObC
dLad3YXfuMIsPoxa1Y1UYXACNxqAQ5Lc8TeMSaW92Xwo95MW3ON/hue4EqoJjaTWO0AKa3bOPdP+
2Z1IuhcH8cIg+FCXc1oYsyQyoN3eKeb348mkNztzv0aXtObPd1NpJAu17f7j+7WJC3AOrugyqSPc
NEGH//xyxw9JiGss1L+N6hwxp3Kj1pZt4WKO/e5A99srgV1GUDZir7z0VjwYiuvsg+rCU9+JK4zm
Rl52djM6OhEm3Pg1zlA9vCNObvE9UUnlhL5lmquX7hjyq3nlNyiv4HPXyNEsvzhh08uLmWwC8BZa
u2K+e2PkUdJdmvh1+CiHrjUDw+finw+/NPPCZQPUcVLjwKxL4/MYI2GADHU/qL3lc1IdRN2WkL/z
8uVDjaIkDWqp9i3S1NiJ9ArXEA0B5znkQii3ElnK3nXTWjQQ/zsBDVI9UCzzSNgFwCmbvPODwGPX
vQ1CMIwOWenke3EBvy3SzVj64CURxKMUKkpLgAKI1wPN2rEIo7+b51MOPHFTrDkLkeXHQsXZZItM
a+MLGJsAJs4hbiTRWdBIqM/WTZ3hH3p7DMW29ANXj1TRD7YcmMH/83/k07Iulg+2M2BTZQ/b+Mbm
phHD68K5YREfyKqxhLZZeSvOs3MiGxXkWZ2c306jmj1oKdkrREkO/N0+pUjLouyNFHwlgkiUzsuT
XWs3mOtswhXjz6lKIvTL3maq1pp68KGgnQaqCWtgik9CNOyqgka8FIvZ4gycLsbz8xYnjhlYRRFe
Cb0nqQ3SCHj/oD2DXwzMCudvDzYLkx6a4ziC2fnduK+GyzPXn817DAOryy0NU+Txbdgn9MzPbFWB
1zfrh8+JmwQ25ydN990stZyjobF3HRzCulcqAptbn+gjKApz129pcZShZPiwzkQaTbYIBuLWl6Dk
TrJsFunbLGChPhGTb3cb8Z0WIWWZq031w7arXpkq0iGbphVT+Uw0O5MjxgFqncTtIVVh2cP951ch
4Ia7q48BhD63tkfnk563MhN3ddn0+eonKU5Bi6KGPv8qePN+pyKfrubmdwPs0o+E3pb+lxoANkxL
V4epAnfv8Wq2+PonUCjulGOdR6n3H7+QgnzdzzrGtKE/WpvCCT7Qaqmmci+D9YxYQqxrC88CYUSg
KmcSFk0dTdlRiW0hDUUZItdIjsH5VrajHqjDx2bXhgf61650e91uSEtZQcteiL7Rpd5AB+ExyWZj
Vxw/FYkzIXepdeXNJN+W8LqTZVfRbU88UI7xD5jWhd+akzxv0Bj4XPKqUAZlJTt8UbfKjJt+xfhz
YJDhYq7zf0no+8LIqJ3nOj4DfBRZE213NSwYm/SR5s7JW7NkpG5Bcx841zeUKvKuq0VH9/8iWMXw
4DmaBB9uuo2Fla6jBRLQCr1oP8nuoTvqFmsB/aFS7oIBxOnkdHtGOJQImTw0qm0qR/xOxXhpwXo+
fmLbCbGCGrgr5p6FP/StbwNZP5TZDaRWxy1KYSXAunAxkua5RwPpKhtxZGh/9/mLA+RBOjgfMbrU
O8Ft3IjUSpU2AU/yFMB64rG1wv3juVaUER0Jftw+CTVNbHbxRcWf/tP7a0BZzMpu7vs91g6Ct2rN
J2FpM7PdKSDWDn4LyuGB2yDrlPDblwKjX1lJIf2cRgXsPV/xIFC9nTWjVPvusHeIyXrokNWbxVMl
jasSdyilLRBfxU7hX2u4Nml4sTmqoSMGD2Fb73xUYbPP3J/Eb0l78RfMHsT+rCc/g1geOb6jdKOi
PUYNqqlMLuIYe0QvcZPzuF1vDZiGJr2P8eleHB3HWGAtbJ9jZfnHUhi+mKeEbX0CYxWkApt1e2cn
krz25x6/9n98jsOIAcC0KQ8l9ZkneQ7LTZ6yO8eDqoxjY1HuyDAtoTxaFqcK/XXqS0FfpRQ+d8v9
MFrHziBqwBY16eH9c1Yt+gUUjE+BvHIpgZe9euTa7FVe0wthLSZiYI1UT7DxPqOdRX+hWn73FE+b
1YJZxP2FecF+V/Z8Bev80mfrwtR8jfbbPObJpjW6dE4WoV5oIq2LL1wq3YXdUe+tyC//Dkp/Wxln
OuCK3yZiZbccr6W1m9xYDy1y70EiAU+SKtPuyn/UcvyZJmI7E6uLn2VZETZmLtncjOXeVmqhVCtI
dwpnTP0Cy8kifcRXUggA9vyaMCBf2/iHxGJcSGTpKzK7j/roNIYgMebGOEopE0mrNYT8P191f74O
uh5wbW5w5lwOtmzuCMJpLpTaSHK4rhlzqvGA/fmWRcoVLeHa/sgjPYmFanibCPTcC7XO2SD0zY1I
gF1FHT7/Cj2S4rm6OAro/qUQ/bat9TFWIydrAQmp1Yc2wr0FSncdmOFJXhsgW7F83TPacbF8+30N
lRavb8L65F/A05ylOlZfZAb2E2WnB3AQmS/QmyuIO0A7PQGGT4CNVVocZd/rUYGj8pHK0smBKbAA
LSju8fZaVXhGykKACCtNFIWEOp5dCcv2G3CHAdHlP2vdJrfpuCtKHNg00BkE7+x1frNqacCYL4lE
+iFhcsmkkQOHTivQjaHKTbVM2FI6BVejlx4L2lbGFE3WvIGysm7vyhbXjJXEbJoeDJkpS6/SQQ1t
i073QQOADy7wt6QozfeWJXd6cyjvaxVPQbFifIeho65Kg9JSO5sj7zOsneATnj2cPqznfAOk+dQf
0yFWgyj/QkiHbjyHbUcoCIpLvAQTEGb9UJO1o058EaWPaPjAJiwk1wfn+xrjjXhvoyLCpW0OvKHR
z8JQxRh0Tmymuay0PVI6kC1S5LRFXkx22l+kmopJAc1jJcy7bUrh3scliwZqHIPsjbpBDFYsgbKz
1iaguRLmZ6+TsZq6MGy6a1k3KzRnQE6G+5riQiBw0i33cmpLInLw31lhSkbCDjT2hTA2ibXqWQFR
u0pPpPc5iffyipCnLppYU/NiADh988N4leM3RMErpfq3HIfyyaqN6M2BA+Ic0WICAEAZVuj/wqjv
mjXnDxh2d6V+KuZlWAhVCntncRvgywbCwDGy6byj92c6avMNrSpb2Y6Y7VGWRI2V1AEFrhYFvegN
6tK2z9YeqEDOJ1i+TOv/ku/uSHQRVMnqaNPnssACPTf/HntoSTQl2s6j/8uJAjdUF5ckWRE2v4xY
A28Kye9iPqdLDHdz+NaC82sFffFoJjPymByWFUs3MFStnwwbo91rdEdvVBK9BLA7f1+6BfewaZuR
KlC+JJjw7lZqDXEdkjKwKN5mS4yzh3o566cT1xZI2qBgrdWZ3/ZnhElZg8u/6173wDxIf8CxE/nB
v7xYgpDXXOkWrPaso4ko9mpj7at5tTSveWDs7XgR99YmeybzsK4/yRyZpo3BQxq7bdn1L4zuoZ9O
bbmAOSP1+XribR6Ruce6Hyy5E5z0Gq5UUJkCQ3hJoPNZ+pZC5r8qoU1dGoCULIp9PMfqAHKW+VvW
mIPsjtlbOYabOZVTocmljW/iKkAGFezXBL5v2WysEiOnTXQcSsWWxAxgCrqgo5B8gl8ZJAwSUILJ
adghdpXdte3sjeDIPrivzg4ch8/0PagvBBY9/lVWF4ESRnsun6WO/BGn1HEWHRzxUopfNSQmZPaY
yyJ4HtWafKFCiHsBT505xPG6kNv+kg9F+8XTEqxwT+v05AJTeRam0PIiBWN/pGmbRsv+mZAOcq9W
HL8/q6g9/IgoSC+oQJoTwUH7/rPtTnMYf+DvBS0Y/Wxn1Q0Hl4ungeaRBNDAdvbWDTWkSaxlXZqW
D5LzLdjmp/UzubttCXXnZDfUAKuuxmliP3sI93j9XC78EfNJEXuU1UfbkRLjwXWxHufGeGZ3k2hW
9DXwNi4IjifSn3/a7ea16ziGB1PcNVmAvNKfQUZT9/vBPdP8vPK4XA+BKiACzXbpR8g4hRUgFy6V
lNFa/HQA+V3Q1klYxNves1tyKeS7V0yq0P9Wzkrz4xQfFVUzw22bQpy1l2LTpGI3+6Ut2hwTyQdb
U2M/PRKVYRe68vUaDNJDeyRmSbBP99gkV45Bdmju1BYF5DK3cOvMQimOhbfVfeP0c7iIF4rDnkcC
L5VzTdeXcw9FvQIamsZpJsDNlxGgQysbaatePBa1cZOwG5ivgQddZqQXSuQf5H+F2tu7P5wql0hC
0R0lqY1f/Ivc2tiPNbFB3prblA1A1yT9DTX9RSXappnYkW4yTUaakanPHINgHmGBsO4WhP0lDlPf
eAKCkUqkBEpClacDhqk6AsBJQWy8+mltjWVnRMAuLC1rmsk9SYxrAGw6d6f8Z8Sk9ahmrI2gp/Mk
zgUvTTv+KNoggMoxsuH9Fs7rY/CALzG+woehwQAjwakvI3epe22MStykQWJZZlhe5WoMsaaAv35Y
LljZK33sBYfRsugCOkGs1eUGkKiVzvxGQ6Oo7gDHKqkRogqa82g3+R5d1yRN3HQRq/HnyeprAZGR
TdrQSzpdVZtzTLLWkNvKiWcWc5KJTkAJpUflpeHWbKgVihElBkcFSx4DuaDJgXzN+U55OunReKMi
5x8fCVHgMhrOBrVXPnVaPiTyC5K65S/tR8xsjnfytKHmMvUybu3y90ZM3dLKUzuiQuqBYf9ES+NU
m0xglqQ7zRy2hVgs0I/FVNAagiCO8EE0Rpyp1LSNtfsTVQW6x+uy4pzYaeY/IE3mQMPpjh56DwHQ
DzrVtCw3J0JVNXHEx74ZkL7qkBvBHQ+tlDY/Tyg88LhpU744LQL84uta8LfdACEOkZmNp0TUjTa3
n4FbfeS9ATNqQNLiwjmFho6fVuqWFztIV8ayU5q5h6CTaZGhxhhn7vaNMietOi408TUC2AcjPlGI
CqXMkGPXThKj1bvG95ItRlBZl+3BWt5rGU+XZx67U7T2NzPeJkqEY0K/OTNqc1SEGFQw1UU6mb9t
f1ar3FRbagLXhUB2bnoZyLDF+YZjKfFmvJuQ3kdBYXUyVGe3h7o5+PpO7p0nfRuH9AoG1kYYUpo7
5VGOrxht99lVk8SbDlcBjwnfaIbZHVWstMfWqVo2+buCcrjMFy3XBc9f2TZS6wSreAr8zzQDgxHu
wvfQlv9iDvIFu822C5GtxKOo3Jcx7cyZeoJgsQaxoq2jgd493C6maS7o+4+qdjkbeyEyKvhgJDlt
AtmYcAYMoqcRN/2emLlrGHigK4TtzwSJlqhLZ8YJJ5VxjY4FtZzAfuq58IvKaf9Ncl2ohZkJRh52
ld2x8ikTepaONO6PQzB5KPfFInjO/AI9TKbEuKp08g2mcSZtsRFijlMgKc0KYoYrrHOtgJ4GZP7q
W5Fi3KARC97CB25ArZB2yUet5phigO6PHx+ZVqzN0CNRHcjSf6XJQsf9GZtBt9Gz1RrL/U2eQXmG
kFuBRNixBRc7+cKZPqz9vq7c2bLHFjluElujZmZ4eeViG3SMYCsKAWwifl1wd2rd3BxFs/Tzjp/Q
BhCupVDHKy3Kf8gE4myknqYkqKePqPJF/wcS5X1a4oGhn/bpvFBXhJ/bwUM6kIbPhypEq1WAhJMx
ohHIKiIHB0PEq9ECVucPM8sQkK0N3NJga3+hTE1TYg7jsKm4oNTKJ8wsN46NsGfGDZFqmXD7Clqz
RF2d+rkuqlo0P4sPfU0Z3kRTOc7pJC49ndPScwqCpOHx4KEMig/ynqeMWomDGJRgZRrymDsn+PFu
/7JgTeYhWBYS7H+z9nmQ6ey+NU7OEbMV0QEanKh0fIhnNS4h17VKR7pm6J/OqH/oq29kfn39FJI0
YANXzABl2JIDN/iQ5pkNuu9dQaq3HLu1t1ZE49gEivBQL+/EFoJA5cBxKFkrBZOQNjq6TmA1ku9u
wgMjrQ/YBfJCRWzTVfaj6jWKuTEYMvmkdT2aB8QrI0lVdk4oPJ0iW8RfTeorAS8rnFTtxfs+SaI1
1MLGNvuG84MsPXVZ+blqEv4F7W5QOIsdQHFy2FT24Z7nVeY6Qm6poM43al5vttVHI0yFdfBg7wIA
JjMl8b1gRFB75dxPYZIKibDeQtsPeb7r4mT3iKUJnDnNNyLqgRkmgvna2haJ6MUzfoQQ2LkVXX/F
ZnwM5IBQch7jkR97QSOROoi4MRBiSqM6TSSnO3ZIcD6ZDBcpGvvAk9bgWlHuoxOWdnHqbbmzt23z
3tjGdbqEgFgfAjHmv/9RTWg6GOoJISTWt4gKiaHMqp5Q/S3Z8NS3qHzx6PeyqMpYyGa2MBjrp5tR
ppbxeY43mfobBad90Gy3Bpx5jgbWtBrKvjdeAuUWE9ANL945f1stZf+PIWaHmMAtnbTdipUAOx4k
Bu2krUP6SScwgUayOJS95FNr0HLLMk8sKo5Iis0guk3sA9shnCTQBuvVWKJGqBRkgeXWPai+/zbT
8ugNLBSkYnxSQoLKMi+mQekLF4MrfunP362iEzzV+G1W4ohYJrFtPhZMXsF71kUoODpVypRyJrZW
Uedx+IcBiSJx8KrPxISBNmGJfsq0ru6XypfRdUErjpY5GMiBQBWjexTTtFjurWNkTK+IPKyrT+WL
SCmvVq1W5A37CQVNcjp58U+AECSDnFuMDgAdApQmbvCjeRUwc1GjXdjtQO99p93v/zOBcsBLhexA
MMEjUURlTKsYRARBXQ/usAjEXKjzK5NIt4Qbj6AmyL1jES9yC+Y5/eltomSW/DVRWBvKPDx/3yNn
H9TlvdLYjo6PJD/rPHtanztpg2936DNwry1TfvzZU57+w6YXauNQE06dSVYCKUZSlmuIqxzdx5U1
s1BSHVYimWfX9HKJKZL5QfaXy6d8+sMO4M/9x1ogx+1n2fqoINykc3PoPCbKvqVeGCCCjfZO1f1q
NG9kubvh83tVyRc2xPLwpJsZe9wJA0qCa3STdhVazvpXHBeThn9vDgq+YRTG2bzY+Olb6n7BSKZw
loZ5weBqVG1pPPbIlOvoNXi6l+nqjQCX9XjH8FgHZrAwsABMM1FSSF7GTr2D+s86Le190ss8uG0G
Fv74qAyOPrgDHogTwAbyLyen2ZiUWQpXzBw5qyP3+WbuKMgbYjAHFb7T3bEhjbhgthDS83bY9Cqx
OQwHxz2r4BzkBZ1GIGLP+6nWe9JCbSBYz3p0ASXAN10b+AH9dyMiUF3tnwiqOrVVIFS9XO643hPL
y89fIhMDcGChmTDQx5hCQEoomVptlVXJR96O8chVTUmGbl6ZGp7zfE4Bl1FoCchbZbjpsRwrw4nC
Jf9poLNKylrcaIq658nONJnqQwiz6cTuE7+k7jPrG/XnlDCRdhmxSKXtv0ZYbTkqkXS35EZXmR8e
CSCxNRSHgku89Fb5rd9w5GEgCnavA7vq5vdOS2FoQFoeCxEA9aARF2dERvyjY0wclkw0jiQVOWsf
ce5r99jk6f5ErmCo62vfTv1iyycByTNhxCQnj4l1oIHbUBTJFv7JGy1kCYdfKT7tQM07dbfOK1+h
C1s8+nZGcSnF9n6RfBUrPIi2xrSpnt8v/H9jnHL6r53VfVTacQg+cdEcwUfgUuKBm5l/HPXe4qdK
TiOrSQ9QmDBnjO1DLdfYaiYehvwofmN7b1Ycfb8d6utnemfAFzVq8s469WTzQzdHpGoB12dEH4VX
zlZwFHzX+FTTOwLD0NUBsyom6NmvzktRoKrs+7gPAIggLlmmyPg1hSp0yw8ITaTch5X4Dr5BTvZu
GwHJxN+SMhpYq9VGJDKCnvzqo22nXGRU94U5/pT7anUGNZnMPg2G5z2s95nQqmMz7Fpvs3BdVpRq
xMwHlOrxaN7V7hpxlMpPfjhB67KjW/6u1dT+xctbHyPTvVz+ymHpNRg35/lKmpuGV3NxoM0fy/Vr
1NRrSba2EfKNnZJAAAAgrgp0tEkiAENcqng74shaYu+4di659hlYpFH/YG1do5O3U53NJD5w6GDk
SRrF4kGL/T/sCLp/72RldjBkAIUbnOIg6UnZDgYvNO0ADa15C6xtIU7bRPWrETqdsOEJsCyWSxqU
YQPAGvXTOicUpxeQkjVz7LVqjh+XKHU1PopyCfUqdhL6gkB3+r5AsQFn0g2RjFn5SspbvpNlDd9e
U2A1Qe9bC4nOL0tvRjsfh/MX4bzqZWDl6OpWB7NhQ+xc3h6zpdVtxiYC4wfIofY2Jp9SA6uWycMw
83qoX7Dt3crwP4UymNwXp5rLOAuLFGrrBSH640m/iM6T2VWr639Go8xvVIK/mfOJuH+6idez8a67
OpMMtlZbfO/MkTjxw89WAJju5LO8A6bofL8zpjMBTdyrHVB3MYpvaLXAvtrzRVXg4NrUjzkFriJ0
YDkt3hb4HrlWq34PomlcAoCvv5Ow0U94RXhTJLKQrF0P6L12bKJgvUmd2j0xwibvU76+YqarTx82
No6eqdOeSUYj7SKwoYFuUNB3nWuKdl//jeAu0yHGtdVtuK9JB9a4kyeDaFdHfzPOKS90yf0QCqTV
rspgukl+eWBuM+nOQUt9/2x52udD7M0Uj7Wz+T32vLnj7WuxZ9tIft71pOqRWGzlmWT1U9GnTeMY
NA5tPFa288USQzH0M1ZWsQ6kJwef/1cyCJaJWwWfav1P9LnbCPOKy0dcZ3Dzd++iVvNNpsQtJNkR
LazRbSMNLNJX1I8g1wNy/6GSpltuMAdOlgRhGJO06/JPURMy+j07djMSg/RDE8RThVj+i4H5bTZQ
B/7lbqwrDC8JNnm4xi1jlyNQ2JKnibS6gY9xXGyvKxjVNVudV/rgEk2ehEZgR3EVbJDsa2RsYgZL
VKcW5ttX+IEl5oeM7kHWs1sXVWTujoxARI27g9V/P50N2tiHokbQpfYmTC7PAIrsDvy6HLO4wxLm
a7zFH+HGFgC/+d1OgzEZuR6GY/+y0OWLdPDTFI8qs0eMUz7+/aGatDhsHNR1nTCs4QJUsnQVuvjV
isTWqM5paGTUvyxmMveRmcZibgAlg17lWVsIjZ8gRccxfRBY5hxk9CjRTFgHsdRnqxJ61lm2SrFN
hJfjYIT4AW6f/wmYGDqh1Mw2nHNkDDD/jfNdL8f/YWtil0bwjJ/Ed5RN0id3jIAM4a+VjA6/YADH
BA7qcsLNlV0wsd28CjDDLcurQtIVb+S+wabaGMNNuLwyXhOkcXppNErVwTNWibPpq0R3NT8Kevau
4l4wRi/v059E6O5+qznEeU/N/CT+4gggFIAlXIYbXqO9Htr2Q41XCASXEKGNoUyEmDz/wH7YHTMP
G7g4YVhzXBC/tLNX7T56C7njh2WBOKVJBhcCIexiqLCH71gqCJ+utW0sj1UMfrIiqmL2Ru5lajao
Td8Uz2ipu6lFP87BH/gKYrHyBmgP8U3r+wTxz3fHlqi9iYl9yTp2aCZNHOqmNxPpxNWenooM+8tM
Tps/2F25HYfBIujmDRWeHjeDn7weYfpjpFRAMHJMR3XDrLzZuTnGpMCjhYyqVjhYITLAKyM0myeL
ZtVbS4E5ke90xhQo/dwWTnFSQHABGXyCzN2qyB1GCSDF7ZpHG47VHvdiIHINRzqdwhKR7rilkJfR
BD8Sq73y/gIH56qLYsaq/jc2f+CGy+oiVpeAS8CZiLOBnZByF4E5NnpQTZSIULiVpFRrLI4nNCvS
18IXZRHPgX6YFQ9gps5qOTWZFqdBXzmTtNJy18vpmHsF2luixvgtUXNNGRDXdvIkZcUz5kqBk/mw
jausEO5NQsOdiXM//rz/HgtHQ2HtAXTeqa0Qno5zAwwuWXg7YZsSiTiE7tjWaVOFp13XDdOj1Alo
JHYgL2OqbsU0S4aUgD3RQkgz040gKCsVdGZ9qDzsZuACCvXjWSR/CdRinqv0WyBJ+Zpq1S2XiRbR
joR0703v6QWix/+m9ZL0sUo6KTVcVAOk6+xQ6bn+YP/UY4kJvb4QjuejPWGeQCNgtddZaOqt5LMX
WuLjO8X4PhFOZ4X08Ra8eL8kKld3utCU9UA9HM6kL83w71p35Thiax+tt2Fg0bM+yrUmbjDJ7up8
UUCGll6zlVrcnS8igcntp407ac468MXt70SIdUfcw09HZZfLtr0sBp5kkUudCCxKVgSHO/U/C+qM
0hS948vDySZTECOUtyz3ZbMWzhylvzZiHZgl1e1qZe5JuxyD4IX6ylq2Vv75ym88lSQiE4MbwtKN
5egwNiXQyJ5jOkJsFpajSGczTQkwdx/XlJ3zWDlTrtexdDnxDLTGasyd++l289p8u5d4PPWo57LU
rp00mxpUxaCcWppn0P7C6khqaO1kV7jN66ljben7hANvvyiMNmh7Bly7rojlTYMrN/L4NiZZVCHy
DvU/uL7uKnVDS0nCEmN2uqH1rqUNHRDaeTWvlFkzb98AbwBIzqx7uApqwzeXID1xUDf8pxpHdqiC
HNDdPaKil3vJRt9khlLXPBB6rV3rHzx5fYZWNFn16qRz3FZEyPi+JdgvZTcQS10qdPkaL8MI3yJr
YPFkUy5BireLaGPVUMiT24d2BFOQGDomkwaovNvbXb2X3AptEwXjxtnGdKPJgqsOKg1gtyIB7SOg
ajQcC8v0PVTbfY1u+g2GTJ+XicCMle4Li07FUKks9AK7CDlyRgNNAuBi5j80lYzutVzMzwlRWd5K
KTKKvY2v4PLDgTHp+P81cvfrdDjcu3gKhBvHWYc6CtHcgtwR2M/PWJvbTUA32RfN1Btwe6tQVnt5
P4RFYB+c6tUKF4GICzWTSu4xYXGMw0+Z9Tc5vVhkJibCvjUHDo4s4Qn21R1QrTkyIIQAyrV7Z55R
y9BaJMqNatNULko7jsaj/MN1ecRszsXxZpewhr2B9lEUFqqWleAfZSuzUqa8K/o5wCfMCebRZ3gI
ACtz8pX7Gi9q3JhpKmbJdAW+oHaQxwDaL4stDCOnLa8b2oQaeBnB1ZEFDeVw++EuvwTRuwU9glCI
Y8wevhqrnEuwOxsYc/8MobxVZmHhWAFBboXt4eB5ohnyNUCmRAU3g7e/DyIxnmiDYF96BkowitT/
1GG31c5zXLGlT0803mVITKD4AQysMKZniMBr9hTYXebyS1DnMzsX/bg+L/TYI87IfgHsxXR96SWT
/SowMYdiIdUvqxCyDsvQmz2UzNIOdfdR2sIsCNNM7n5efCKhOk0qU8CXApAGStsxBKdVxx0apaDA
SzVb55o48ssF/iM/Kk553AZXHgjWhfR7hnUJB8uCtv6+K70//ztiZQf8ncZCpfzQwPbIddotykAa
XSOyUYcsGMKlhW3RghioYFnQN9Y8ABlqI3dZ8YunKN5A+cqhpWTMjUBd4LruTvL4DpCkF9p94J3G
tZdR5w8inKXrGJUutrO7fdxmejbBhoIpLHEExtA1yY4jrr5NKdia4utCwCOU+d65bEUbePWvYAZ/
mmqBZOvsM8vop/4SfeATSg5q1GC8C3mo7r0Am2DGps1f19rG+7YLNqictXkpCHsISSGaxjicJJ3E
FHQnAYzgcaeep5NMPzSBeMqO0gUxMNPBryn2acwrX57mncr4mLyh/WDn/bxmL8y/NBSyASbI+KMh
4H2Yp1A5bFWSkb+aDvjDsE5vmOc36vC0Hk4grXqrVUeV6Zkq74GaaQe85U9k13MooIxAPqtbshc/
z+fL1BYObj3Sd7mpOWLRu6bWEUQGHkzv/WWtOKMoppDH7b58V/WTeZpYMa7NWr6Ck1Uwep2cFxHt
o470GE4WBU/1JaqHWxaI4CZGPFvgWF+nFFjp61VIwpFx1n7hiRuarm43aXA656HFpAqBnmHKJ8+Z
GyTV1Aq1GqAbmV1Cpa1sB+xJlxp5pPZlFnZob2R4jYie6i3vTTz4x/Io+oVOvHqa8FFvtPB5EXAr
jeGNbbYTJkA+/hFuqs8IH4gxphMcx8TQty32jWOnjUnlKfShSGTLsqlzDGDfFPXizNIbmUa2aqRP
r7/oZZsrh7zum05leIQRJOoIEA4NXnW/OwqxG7HV3SHYiRhj584w3dE5U2MZdklDbeGtV4XWIWBA
AnfjcmJG1MASqx0gWC3tpzAfxps2WeAgVZ1WcfziWC4RpBBxqhFjQKPaPuVc4ODunmLNsr0/+g1C
SFMfc67m/n1bap/YIKte1YWL7qT2HMc8Px4bvHmfBbbawP7q4XjHwRlCdeSLM0mipk+GZIgzaZFu
a83tl1W6jO0TLOfBY/BFG2u5fnd6ltVLrvC1O6x0dUICPq5yAtR87pDeGPcvJ0/ObGF0jaLfuWOO
1pxB0PUTr/smWj3lgK78DMI/ejnkpuCb/g/SJyPvkNnTSlzQeYeRxTE/kihp4pGg32XPP1Ax/3iv
6CaznslGQ46FAXPbGDHP9oqu3fBjRDLxkR6dFRaGMsinlkNe2XX9KMRYmKd7NEVoaQnAGZvE6CQR
ApdnCwrdkI+E/epe+mhSZR3/H5CNgCKGc6NqmkRzBHCw2VGYBmDJKk4v89o2grMpB8HaZfZ9u3xb
BjTkWSBS5nE/rJ0Df3NagbTEmC0gkA3Lt9FOFRgbsRcMIfbSoqRYaV4YrqxbDnI4X6Y04mdg37fx
uF8GTAocH4WU0pjuCMHrVR938a9YAXgU1GRLMHzuaidUSc7TNWltqEmLf63CQJcQjWj5v5PEFheN
PnJeDaUsnbXfoKkxFmNgBtY3JDd1yCXfr8V/2Tx7+xnIgCrSQ1uyODo6/dQJjwtriyRKRBFel8Pa
ndN3qfbvFNBB5vTCsuwo1oa4aBzhN+A7GbcQemZ6wjuHf33BlG75pwYaK28akQHazRCsRYkMq0YW
VEZFlc4LBQatKZk6x6b3Kvam+NOCw/zz/QB7Ri3i9P2E7g2O1XU2HkwP74RYdQenjqJ6jrC6j2wl
WoydOKZqoOCHp9zzhZEl2OT38N2+CwPvsmYajbIGUAsKpMmk6nGpZirUa6COXguBR008c45p3k4q
Nk60rJIErhS/aWBAKv4kr7orha1HsUI3+5cB6NZI8tmj25eYRG8urdtJUhhvAO6ugJB4rGnscC+u
bOKi7LEj9RhB6VH222/Xocks5yGkaUE9Oa1tKc+Q9sIE0mOx/hL9eS/w9ReYxUSbC1n3VNW26BKl
6jTYkyuO3FjOUvfL/P4YvK0YsbIy57xEYJ8y1kvPt49RtoFrNkf8GpjjBepyZjLPcNkX6EK/2HA3
xwdnVkUZO0HbYrfHxFlXqsrnWYLwxsz/QVeB39AkRwfDk0EanEpsemhlOVoQBxxhWJWZusT/EsKO
hBulXggSzER27iLly0+rElcJeGuifCro8Voi/bY15Yy6P5M7Y23Xc9vop9H5Qh5P/WqesYKccTln
V2bttx27/ZGYjsmkNiwwAIjDpZDYJQKm9cO+T8b/G1GPKGK22cVe2ok7be5gDwkkHIbLHYm9kp9O
rnVEigHu8sULbUidUke0s5Lk/dmsWJ/DLSXSwoQooVek5tiXpZ46Jx1NXYtUVWVAZOvOlarZ6gi7
pvHsFli05QhSI4sgDRcHN83sF4jhDWuEJvo7Ue4lXGFpqdZmoSeGvqGVeEXOVddZkqnoRvrTOa8o
n2/e7Ey8GogoalikdEeiEqNTt2fAkjvjB7ikKoQoP0LeJEIH7RKiFD51kSYY1gZrBbLlTC9RHNh0
F3YBD4lOXEAg147PrYoL6GWYvvzWpRm69REwSBCJL3E7peaX2ynKQZLBmIFMTva/WrR7chwt1iFz
abqr6zov3iXGZ4V/d56Z/9f/LKRS87XJTvZyZz8Ho2iQbQoHbO4fVRpr/rItM4C6+GNbBXb9ZdvF
FqAAGqiPqFf9n4S7mgWu4Q48JMxpg58+GH3F1TytoMbDaLiUntt9DJzncgn3pZyYn4ygjj/cu3SH
udMa/QI2nwNChhoC9noAOD9KYceCJstAE/NlpGKmY+FDPQXVdRwEx66AJXztb/vuhvnayLZC52+4
yJAq/F56tDK2r6oAmUhjCBPJJk63r6Rsf0qE/fz7tRf3DHrLN8zI8lrLQxZhUNIvX1GxGfg4h46S
sVMnIxt+1VseApU8BTpoop2iB4OCnBY10zyggyvpfYfYiWVKUasRgcP4aBNpCMj8uR0rMfvJ+K2W
55BVqtLLjWx7FaAqhFB9enkNwW0/2cOySzlJV+EWDndHpP/g38CMsOCyWn8ZrXzAiCyt5wiR/wIY
Fngx2dddLtjxtgDhc5YoW53e8WqnPyIngKbpf4NdVF5/kapATs8HIDB/XYQP0k3Djqa6NKy1b62M
RuYZanYIiGsUeSs9ow18lI52gohsvD07MNVsjK2QBKhsJ2W7bQOQMoBgsgPcINWdnuqSZabvqf2o
oL6xaDqKaGIUUGJiSB0mcAYRvCCVPzgNIfUp7b9Ds2gBBkJQyGkmE81izXla+PWmDLRxMHcPrsKK
8C7zBAVBKhpgaPnpffj0sFYjEWeKQI5IlaRRAuqsNh1tlfcXp1q27lKwZSbnj1zPOu7nXVniuLdF
4hNbJHZBylxSwJN+D7HLLx/cecPzTexJIt7Li5XeJxtW2kTFDLGADT5gwCFUXv2/x8MuNVOZgP5x
/htgL9WfaZJuHIxW8bwJ59E0epTzYa/vbfGgEfW5UP7elz6mnAS7ElU8hUiMzKhyxTKE/wr1DP4w
2dXRz/CdmG3N1sy2I4YF7xe+DLFjsCNKNAup9OJJvyMdpEy/jI5tfOL0uCATEicd/Qx1aJtkeawC
RjgJT9MKk52JUV9/y7AXTjM31tRauRum1XHd3aw0AsRjv6Ti/YyIzg5CA72SxJOfANvJ11Diks7J
D3rWkoVm/OKIKEGmIVGc8l022kX1lXJ3dVCop43MHZnuxMDaaVUB9qgopUiZAbceFX7Cr4m97B3N
OveJriuM93u5/L2VGmOFCua42QHMRY19ZC2wvLwp1IEEEiOyyyWFKuT0Azr7W3s/wldsOcD44YaF
g7AZ3r1jQZyCpnJg/pJa4zFPQ2kOyTjwQEqmEdSJ/mzJBd9062hYk4NmmkIcEK2MUb9/Jsq06j3x
nD5tT3TN5avnTfyF676VQGkVYi/7noF/i1ThR+5GdzYEdA8yVY1d8AFOitVZrDNJ/OHE2AJqJns7
rUWLusJQdUCX2G2IaBv33kN68+/DNGy+1q8SFUQ/yGIvK4tMJPUr/ytY+d+6PKxjC2WckfdZdYFn
vnXY97R2Kb1xTmDZHoqr3EL2PmdJ1ZVAZvV7OwCLhPzx/8rjKQmwD67uaQ3x3O3l7Ts3ZoJN+uXV
AoXNpUg9YBCzTeJsU7JV7xym1vYbSD1PqhEJecXJTwn/5/TTVfRJ1bPlhjvXVA5Ov/eVHuUtWTUO
uSFo5IV5FlHvC9Remf/gC2UWV+r9T4VvfT0GHUtrsYsAY1TFAd4lUPnMTf2EghhoWMT/eiH18/cU
KSZzjpVP3DCSpXCPW9198eqSUDD2c52FZto69VgSRczqUNWd5DS2LgTLqQOu6kQGMeK0eG5l7wwr
3PGvkIHTsw9puuICZ9C9Ms8U7yiQutsd6cmdqh1uPmuycqiYjGCyGq0x/rXyTJPSL3pdFZNZd3Iw
v4UiehINXphtT3VZ8bDQqtNZwo1Xm9RdCUC4h7UyDAYSZlrIW9nA7BEPtSkGzlL85wRogfX3qEaj
hboGiwKgn3bodTyboVBm38bn4TnVTOGTkLCt9Gvr1wHKteur3l34ZDmEf3fRUqN61MnChphFVp4q
uUOzn1UswS59pxpcbiE7cl23yWQCNrugfwOgj/hq7H77AFlr2+MKq4TvFP2RS0/dkzuRIOiom0De
1Tu/E685BWM475wx3dBJ/ri1m2S/YbsvHdhAX4WF5MxNr8qh89tSm+Nc7o9u8tpG202NXW9IePvX
xdBZRi1rP6bvFyZUJv1Znp1HIhNYf559wbU6JyK4TPQ/YVdF7sI6y2mN1lVpadebZGyDbdkF/Fmu
Ofu5yl3HkKMG6u5L1xB4n96F+Loo2PrOdCIqFlEA0+9SAkQ6kZ0xoAOXHmI4kFdhmxs9gAw0rtZT
jMG3ttzF9hyQgMWHpkHRcqs3uAcMtFaLfqm+ve/L+lCyil0JmODY2Q4IW3YarM5q1BaJ1aB4kbC9
A6ci5pyW+205XuVuUiqjRBTslSDbw4/YbBpIgGBRICBRzzJeo15vFsqBuw60Jyql4RftUfTD5Hoi
UNAQJZnB7MD6PikRlV3Dq7i9oD7XXIdzxmdfYkemiWS/Azh01Aq9dfAa/xijBTSnHIXYt5SRbMqh
Xcv98xlpcY+GVEBVDrC/G864o9O8nNHhD5y8MQzV/Fd7lwAZBAXW1KLsWjy/VML30tSaObMn39jw
q0/SL2ape2Vf3lqdX3DhXbGO68XDAZ3Zb+gTkJf9f+9FF0cEG+bNbeSGThQ9gU90UiS25abi/m4i
oQVtGm7JUnV+vCdwpf2FHXlPaGiqKkTDgzguOcrDkfz6uNMEmFp1lW45Zxc21BuO/uBw8+KUYiQh
7wEg+y5YGHeYJhTtyAyLS4Mq3ECNGuA6MK56UbhoZXVnGRr3PawYL5E9HAt9TtWcAP9VUvKK/pAz
pgc8QCGNLW6COgxlPb9nSRKGKDE5gfk3fhy8B24kvwcACgJaUr4/D7LP8cvXlkeVlUdYn2aB/k/j
IDLz/x47nHLAJndDrKjpfeIUU1dhIOTTUffo0hrpPbMKjXa+fY2ETGol/jN1LkMAf71jQDH4QWv1
5pLPwu2syZolPtJcwcsEWWsNqk1vWzJwuezDeVjzfupXyoA6NdzdEXsYberrn3TSXWuYn2CO6OJG
Srg8t5rtnveLxoyFXzB3OQ39oBeoc3qQM63O/eJO9IID07yy+IImHvA7IIQbQCoPHylC6QB+2OWO
i/uU+lRNfX9wCVLpVy9w3tCCRc3e/qmF5e1SzFnI2GErhKvnHedvOlM1DSrP6FmaTK/zo8dxwfvi
TuHvH3Erf1BUaDbu031VhMkInpUTTrXaIZ1kLP+uIJ27reNsdEEZ2OrpuPd+pymVpOZOnhvcq5C3
yVTUttng7odWbgWTsDv/7zTWxXnK0UtkRa3oCqSFhwcp0YwZoQ1vxzEchdvF7XQxAE7sH1QuObUB
r2yJkTW3JLDLgzsbWtF5QgHV/CJiWKM00zpMoQIvjM+YMVDTL50VMR03IwC+yenBGY8xw3d01d6R
8jKQBpX5tl+8W3PPEw3pc3lrB1Uld+9Js6dm/577c5UXGEGoAyxwNIekG0nzOaGUwUEU+l9ZrtlP
CA2+hUlFSuscFasaYfbMdlmPiSjG7MqQ1iBB5ijLgfEjcMCb9xZAgZgAEQUq6MAEJWt1pzFpZaKM
u76yL+c0YKZEHDLxAqVnpt7/kl+NBi+O0HStqw0QpfYgHhKJb9htvNDAO+lgYJjx0aaUCutbBV1Q
XWS/iJjzzW2qqOygbuQAzV4X/J7LeDd5Eolvl+PCCDpw4pcjXAhdYcLgnhY7MIEpStp0ZqgokpbM
DHBeX/Mdxe10oAYHD6OrbFKa9gHJoqrcu7QzQZBRRxYKxd4mJHGAg6roHvqtZZPUjQ+YdyoOtQB6
nZ2RMxm2fcTNaHGhbDTVp6QqMOosC+xR2YsImwfqF5rXjVQnWL71fYk1iuGhEtccnuY1KDjH8UQb
sDd6Ymf4KQ8jx8LPs99B+QtnY3Zr4lXSUxyI0tqufStYx/sO3AT6XfefrjmRA4wy9HLqsJfAcyXV
7faJp8CpqIWu23mnmEttiJBkBw5TY/KZQHfzotTmmZ7UHbI7RPtzOR9xYS756HXcPujpgF6P5mn5
nl+s7tCwLM43lA3z+lpcVJ5gG77I+xfJlKRS52WW4gnFQcoDf12GvWqaUnDmbA3rMhaL8mA5UhXF
mSIithTvLDrVUbuNHlM9xtHWfOGRWe+ZQ3C1OohbQ6gw8Oqt6fEtXoRRpktcKGiQ+UakfxzDKULv
IPlCkxD1Co+i8lTPRWudXS0eauG7l98lDUwo/lxDcwoIkD0gZVD1IZWlUUrbFvQlW1JO0Le3hDC3
emPfyJhhYQDNpYnXI279GgCB1ZHjhATkhBSWa1kLbzZtyb8l+uEZD6m2yF5hZckNrL+pTMtC3T1i
wYWBc+VeDy2/Lw6QXMewSdatMnC7tA6SrvQfGHXFfJGNEJCm+qf5nNyhdNqYrFNJXXumqW0YIqn0
GgJSY2uh1xOwb59DB/hQB8R94rLXbj632GoII4yKNP88Ptu+R4oPcgypOPZ1/QOJ+8F1gnrqvIGV
6iR1I5Z3PRuOO+UP+oSfG6PLOdGE6NVfbhLdOHtGIM52LCPd1RxpKUEzAS2bV4wlvYsUsGrHE8Y6
ONUTMSwjF2/o3ANxiorqUoI9Su4bn2dGR0WDRanUzbBbVcWsY1jF9qCnkEj0qA5dtgka6cGSee6+
e5KDYpW/48unW7Tie8q/pZHstb+rT9kfYJrA8fTtsivgq0owzn0MxdA5uWKjUteau2O3ys4uekYO
UUENIoYXvK8W8imLD7k+ON7UV0VNUMKTpGwYoSMbjwVYdAHzJmF7k343iVpmYHvuJP9mVF/mmzQV
lKQ/o2ueCEVzUOwSSl19dRuQYg6X80Ihs3ZbIJf1xEvoeKRnPCzGL4Hxl5mVgeKcanj9Ym0T6ldR
99SJYjwJOT9+bwpjdqY1QvOhHNd9l2iVbdL3wEXR9ixCVBJVe9DSYz8PES8tTx6WzYHIPktecxtE
rQjA+N4BwiS2eVhKhr/rYWKrySojr+Tgp85ZznMUH4cJ3PbSoIm8aZfpIQtKDyRnlRh7wnEnLvsQ
fvKaRXH38m+gfYxmFAZVbbkX6MtmobcoQbgp994IRWgfIBEOrfcj+8KteIUjGUShgDWiy5zmhnDN
XZQDCJ1p+mhKaWw2alZNiv3BmhRi5vcvq4r7Set9rXTsDo0k2FZudNe8L5UN4Q3m4mAJWqVSC2zH
NWgYagvtrz1G1ZWf4FuSzEOJ+kCUr5r0nQ3wA6ywTqERUBeJ58/Xc9xX+tfpPLwlQOmYNdVaAluI
Do4wzp64XwHwfKzcTXqXFWdFLwgNBlbyqVtdI/VQy95m/TgdYDzeZ7dLrHBqK7F+7t+LqYaGsa9b
Jlqb7+FlBwHc6mODea8eu6rDorjEitjWsv5mZ9+MqsbUoNamRSgbDM4mnN0QnkodhhMiF9vUUm2Z
xeEOCrFt9Y+kCKufK9xzPEoaK72brJ81f/JSo8xLPsViASEDM14yBVVdrJU+pGeKG0C5SMzYnt/G
oqXc0w9lGFLkP79BAjEH/415WggkYFll8o3z1EcAIMbkfIv3zSqqdnJXS9m47ptTbMpqJYH/4wv/
UX9pVIf8k2ovfJuaBqwyT14/es4hkI0lMeStFSAyF4cmcCzsy3/SnacSFN2KVQX5DhiLrz4vD4X8
mokV5C5CXS3kBlsNKGHfRzbJQuvmwsLQzhc7CSlaHiAXPPu4K7ISy6X5vxPPljdy/2TfXnV+pWIR
805jn/9bbByB+9INISW/xAi+/0LAt6dSg25hZy1HBnAap0gjozKy0c/IQPQ9EI7tmjet98r+UeHP
I1CoHsRtjiQkrCEFi3qPSWAyZZmqa3dYlXRC3cDZQRYma1JedakI9z/Bl5A6t0yb0j5tOeXQL0xE
LL8CY4s5K9sakyyiI327WdV0H3ZoLqcuhvL+ndN7Xir2vkyEvNMSoiMU6oz8yGSnboHITQ1yimTC
CtXyo1aFHlAkuOGYXYEY/hNabkv+K3PkSzxbFg932IThs6Kmgi7byb+UCU/ato27jJQaf2vXTlUT
ZgMt+DJhJ2nbgsDbpRKa9qU0Kr2Dn/xKsPf58pp7Gu2maP/wAGwn1NzEqs74R4x0nEsgVAV69iP0
EMc+uiBUcDgFkbUFhLve+oL4szWktGAPYZpoCzNJzZH92/tZcVTeCA89DqLaE4KgV35v0cfpeGBy
EG14FwB4rxccwe4NmdT8gTZwYBNvI6qT+cDfgJB9no/LyLzaXMRNXt7VxUcOtPbdwEsE5LxVUv9W
R5LW8XtvwV+yk6WG6f+TNkLRF2VMyF7aYm7qjfzXhHp6GRGVSzKF1Awx4GeF2B8cXzrJFSTNhxFU
x7kz759Y2HPnhuXfa/WHXIZUFbI4CqIDkdq4BoGIrkDjkTBug87j/JVDN36tQ1cbqWdE4xFmT3n1
clmYYtY36B9Wz40L+52Eq6XNpXW7BPmuI5lzD0t+lbFgMIiNk2zt3P6MweS3B2JbQG/KhyAp50go
B2y7mV/1XNxBr40rdGqbre511Rw6TcAZTMrdu8CZbVUxOvpz7+ZusT/eur2EhbeZgnsXC9YcdRg8
pgfFKbLmRmu7c6HNGiMnkpZyuVgAC8+WSPuYq37g/WsWcZewwGsMItaYx7siuyzfuwXk8ZL391qo
qCZlP4I0esIn7RCJZj/TxCmRt4us6QsndlduOQ3vFAs7uVm+2BPjGVBdWcMbeifhUtjQdkY9x2vX
ZzkBjLw0ZG0jiIbnRTxSQxnh4094K5cj9wTPOj5sAtEtMCQ/jwQ2y8Pldwfg/g8NvuQapgzd7LVh
F09q8bZk2KsQkjjmHzr3TSgib6db/ncMq+xKZZE85BLVb0fFIbWEdWXi3GWjIHbSCX+z4aE8wksh
iXrGxil8aluRbnA48TvKhtUn7EhJXnbJrjiod1A1mBoYfT/iX7qTaXOHaxnu3Ye98SfVbYTTE9uv
unXBpyZMPdFbhmq6Pl0+9RbdSa8VY4M9uAa3cA+q+ltx4GL8GN8iE5RU/cyMuyj46kbe31zSNG1V
Gw4Ulf1lPy+KcY2Fu9PNUsqFrUGSxsKj4Ug5qPB1pLmhNsUNZf14P+lI1UMc1YvoyBJcHxoV6AiD
tMjNLubim5NrCSyUi6Gy1xFK3XQ7M0PiYiNEH+B2BJpXZOsqgwd7LnlLwNjEQkKaancEP5rlKmQ7
2EEIKzSMr6sOTh1YlWZ0MpZqZNCiU6wMWpPxBFtIIE7cJ2o9bdZgFHzWyQAWvpKcPnzm2kD2hxbM
qEYNFppdZHwdlIkeBrVZ1ZRE2//9+tcmUSY5KrQXvv6oefsUpYYV0mZLyhHxIaF80izxg6pE3/OX
/Dn+In27nkE5yYywkhUQX0jHcnwOZvyeKnOir8Jhx0Hgr2kLcS/fT/2MD/cg63HVIjSuqVdHQ55u
RQw5PeNnQVbe+9jG892nhZR6UOygCMgJ7A94W57qI3F0a2RNnLL4Pe6RXVx5b+mkl//7wBYyPXlD
l0W5Lcn4vGn5bICfb7CNejQ62L+7EEtl0TgeGGn/kgzwyCsl+UknMdoY9QOQe/+EPfJmC7udFwV8
7ZMS1+kcI2T081K0IsetsCRtBDNfbFJBobyF/zBrX/XnrS2ycYZh0iLQGPO5j3/Mofrhnk7TkpUk
tf3imd7h00SLLCshPyKf6SRdk8vTOBjbsK/NOOr4VPczXJRw/iFCN5e3gxiaZflOeh3iDR+RMD3B
mYHkixZAzasNVeWlSBwQ2CfRkdKVsD94keyKzTCQ+pKMGzqFQXO5RiVHn9ajmSCS0KNHFLoEackw
gpqAo5ozhQ3NZI9CpcT5hMFi0v8g7fQUZ86XnJ8b/zHRMYoK5z2ahwBxLb1Zkn2BEAjjf0i7ROcy
x8vHnnSx76M+2dredkwRCPs6Nlu83hZod1FT2Umdcd8jYC4l3oK6bizhYfwwOVgKOsuhL9tNYxVr
cI3EIVIVw0jjxinBOlUaHO/0p72g8zi+yOg7uodR6QxG328S+j74n7/JGHkg8EMZ8uLoEAy8dak5
hwgY9cDphxKjLOSFAzagggDEWr0r+WYp9DdSa52/LU9vBjG85Umi+VTLp1MpmeeiptvXleCBnjSv
re2ouMZ1rlhumbJf/nYYC8+kfXvLCTn3pHkKqqATdS3xh/gNkI7IbVYI69VqkdJcS1cqpNV2MYJY
2h1bjBcPsXbWA7MBzHoMh0H2We0+RI3Z7+QB86YiXnWzvmx3KjtejkGQU3ojpI4XZQxmp+caipoM
aW/L5yp1sTBy+aHXxpGFX+NaFEx6b3yuwJ/T2suNc5IdZG2CC5ngO4h1+017jXD6ReUC2Sll7TmD
5iUQzgzR5TrBP01IM0voz5N4VRvkXWkS+16r/dQu67jcL2qDpuAenvFT5GuN+1VGzrmPXmBCOgMa
aeAx2rrMfvfF4XfIak2C9/opPW1FgV5rGf9/jaNij+Obu4MzpIvbI99quxkFrogRGSgSJh09u9Nt
B+L/SRAGI3e00b38vJIoHtTRU8RA31GZbaGxDXFrvZDYs3LwYtYy9+r0PGRfws6O8uoT8WOFBN9e
e3ebIYsy6+UJVyAFZR3rsV38GI3t+e8o62mfNha2cy1irOs5NbPx92FRJplRnrT7Z8NOI7UC6sCL
D0mvtECmSEINsyuNFNnPha8hc1qL6uclEjqKiuKcICN8DcokJaHjVT3/COgFly0gYehFfE49lXjl
UDvbCK8ZfT9/QH07Enti0LkLuddSkcVdfxzAWpO4Eatpc4e8s5bxFadconzfzH5zk/UWMW0dBdlM
m5DN4F+AhOd5FSbdgcwC7lDa8OiHH5uc3r/1ZhJeTYMesxbSNzQkGWm1mhK6Nn9B0T0SHkhmtlL6
+h4aGpI6WRMkGozs2zWa+XlBc4hF1ky9TJ43y34PJFmfOHsgTg6b63llBs/F1qtcHu8Djusu2HkL
IC9i9WzqvYZN9vLpS93syDblf4iPqY0zk0dES1Vwzn0POAAHkS9d/RMCbfsXD1+1IkiiNRlKklK3
EPp4mgynJQ4+vNvNANkK9AExsZeFoK1rhJv12eVDGFYJsqng34NAdrc3VTCBTSKWhmPGRaH1tQVp
fbGUJG3biPQ+ngQarYPTCdzlNY1bEjcr8PBkAzPprSB7Nxbl8VZzKmA03UYSyrji5dThqz5bXCto
s4LbaS5fj6b1Crr8igfrBo52OC6Brrjpopn/X/puiplYf1pGEaTbl0esLrBJX72HRe01lkHbvrgE
B1854+hpvRmYqBuU3L9AJanvWo4sdaiMm/pIVe50v8UJdOU7x9+f2JvuHokMY4BeIop6RFKMvFQt
QJpJRVNwEGnXaheLaL1hZDgXNmZudkQkTdUDf25tTgScQU/ukt06v9hUJ5cNBlQ72R4m067nz1SY
iYAL6Prb8C6EtvdSp+RbAjma/qPYSG6rX/qaJoBm4VVfaGwSqpM8D1yjeCM1jzMF/po0u5/E8OSF
MacLsUJr56XZlrsWJe1t7o6gWf2MlZSGeZXjsAWrvOA1l2g60w3SqqOnp1weoFvj72vADtOVpzzQ
y0q89DxUcthHX4rZsM0trVEa+9xCsfc2QwT2U+7UQTCUy0ZPrLyCIoGXBCbEbhyqJJhv+5N0/zoe
aVd9ShOUfKZc85auc6vLxGxMvOJgMvdHq4NJV+HKcXP1v7PbA+S/+Zk9SyXnPuTeW+zLe+cDILrI
De4U2wPa2tiE/8LFg7550692Ox2BjsCY2lAcfdYAkF7zJz8uL7VdhqO7SyYjntDeRya9P9ImOtmL
tEEjrH1S/QpJcZ9VUA7XmFpZ5gTlxFpN1qm2L5lGYHuxL3oXCi7GYYCqMV+9tRT75DjEbo2ZBpuB
J8tN6Lk5ZQRB/Cvqi5cpq5fkxibhq6UzpZJqphTtx+K7IH7Z5tPzsoeaxKQnIR3GAEAj+o7Brh3f
Uukhbjg66COfpCDQNB6Qx4lqEXzTPqAh08KoH9F+/AV65Evko2ps/E3qExSrZGnKqDJ1NK6+Si+f
m2TQ9dwGWvlGDCMuH1tH2kKlbKz9S/W3oYwzGKe8Un1UbMJiRahlbcgnu6aD7sZ8hf28PH888/vw
89hDTgOZUVNsuvfX5zSrFBV3pnDfo4oQaYF7VUKU1LuykDl2GowJbGCj/w8RzWP5nko4YFzH9tYA
9tHbNiZDzD26MUa6NDHj1ER4PRaE9fLpwGWFxv0SznR8ZtiRLuKaOg0+/oSVRLMW6rTFNpFZSMsz
3g3tvbWq6OgB+XvIB3Cc9fEHK1NvjqZzVWVYsaOAeIcoolOL+wU4EXaGxr4Us3msA7Ztp0Onm+B6
JOuF/UKUODfkBDOJSmf5+TD6fIMoDSVQa2pUfRehjb0sTpwNuvpbqw0WqXH4w9ePzdAONDcVmmo0
QLXjjvk3gBZxIoqYV+jmlDxGpBE/DsqEQzHJFrrLudQ/TOZ8PIiPZM+xMck9vEoLN2D0C6zinZCv
tyroDcIg05kZp+8dJ/lAvbDUa/dzbLkuh/DTV20KBwpSBAfA4fwLAoL0O3jCWTPvwJnugqWfv3mK
vcEoJOgGs+jenEBGsVBOGV295UcWatm9Ac2+aqHDXxmVsNsF2RkEkpPgTde+ZkpvLq02gjvh2I3i
rNUpAMuNhY0MJJgIBBjntkr/0kN7VnCmyN90IGPWD3sE7FtVIkmrxEQeeObcJviDgvZiYgdl8bUy
X5dA3D+yuNpuHvQfRjSJ5NiWY09bnDgroPLmoxWRNjeCelkgwsraab2MyeFlbRSuGpQdROvrAIu/
NXs2/EPHEi2Rc4HLMI3zsNVYeVf3yrmRbUfaU85xm9U7pGooPHj1sg1d1hoThgUxf619urtxetCo
ziDRAqv/owEZiLS2Et3PgeuOtwz26Hotn9JiLsBj28UQhf970VnxDE+FWGcg1EACG3TvStpW7Dmz
q0EeDWVD4LpTF8vaEISMTTYjVtCnYuc5Ijl6gNGYkvUksQhLiCnjbnHP99k413C7+aW6XCoxTm61
24TZp0EBpgmM/U5Xk7n4jHf5Jja3+6RjoPHTYdcoGHwQPKVGUHgH7N/aVlws4+U4S8k8ymKbYnK0
2wnx1v+6OeEDTLfNDRsSzmDKROwPfCPrRcUeubdABObm7xxNfcmBzy5f7fp9BPPgj+lrN535U0/f
bQitXUDytZWibUcF3u43gnn6rRuyXcP5ZyfHO7SYx67YobhtZ6TgWp9okWDlz4Q0VfTyX/gnPmvd
KbG3r+mtEQSgKHsqet8ZlbenBTH07AcMzWSEU9D3fHbuOn48ZE3sFOIyJssXMjtlSHOoupuzT5WL
daDeVyP6h7UKMKPDJlVaEa+BhKFCd2ff1OJuTRI1WmaHFZ3+H9JuPPM+dev7EC4jL4VAqMduk7i+
r0T/rNB1Ugg8UkhcE75WZdMM0UOhrxqW6/ioV+mVKyDVr+N0xldx+IwQF7ZNzw/HJzQVkzW8jp+N
ZZGImFeyxKyTX0a5y3DUeeErALhRXhcP4WArRxdGixVCsx9ZW0Pa6hmoUXDTPwILP9LcS2/1MAkN
91rjD7C3ihOFq1cQ5yuTO42LRZ9U1z85Q/A4GYjmiRpEBna7HcLXkke0W33MZXYJYgpDXpqSr8zZ
e9c56RNBTmyN1EFEa5qALQw0Y1ryzj4L85eNvNyd3eqOkC7J71DfntbEdADaVnOz+AjOhwQwWOqs
S/3NfGZt851FsltmIzS9WJyT29PQYi/I5606gXR3bSxa7gLRyRob9O60POag83B8VpdMiIWp1QRl
xhMKnZNsVmCWY1G68Z0NKR0fLLE2UbrMbbQzv09xtPDlFZDPr9HKj6g9apRAllHMpnGnACQMTwBD
tmNk2HQ3pX+FoQkXTfbUsdvhYuH73NcRfCvDDYqpU/6GUiAbK2ytSkiS2venyLM7Ud30yZHOd1qB
sIwPz+BYaUbUqO2c13j8THckjEm9TsjZbH85MGyiMM5ExIyIthsTI3KnHNv/Tyy3ISyoe5n4UV4k
OTpGZsYCKyl8y7P5IH7mgJnPY5kxkSD5VzVPqFX2p4uJtcrkwk2YtgEjD59Fr8jCc4zgQglBqedj
TlOZ523qpNxbOdjtK30JbMrP+FK0OKthMd6VgIzk5bubNm9A1x7jvsq8EPNBouk65xS4wrpnWj3o
UmVkcu8StVFSu828WxIhS4sKNtd/Ywoe9SSN4V4FY3qA4BUfjWKsOmI3mLUiFI20FpKGe6ldznf/
H+g8vb/S2Wksl7BvkbR/yYSVDJCvXaqaXsa5me85xvlNmq13S3x7WhxGg2fPJWVo2gkEsgI/2e1Q
3CAD8PWCox3TMfXBRskOxcobqzUQhWmr6fyvh3r/D1CLvrhn4PrniYhRvtj7M4ta6UUjz4yTCWdE
wVsHsy9wtY24s2Dw9F7wCIaV7RPCmhRs9PRskwKdLVnDeUpMB8vdHHrka9cW/Zko3hX7LWJNLcsv
UaxILmXUSyrt+h4fEZFIUCbNo9TQ5xdm7sRKOy4n80xLIEvYQlzwUTkQ/MC9HXDOCjkR8Xkmr8nN
0ir9cePhzp0AlDdTny7OfFkXdcwgLPxLDJosbBw4YxGrrs4WKMydyVFgN5ZSd54cLOMAMVl2Shya
7GzEHJWCgUVwz5O7txNvOUFGCzOAf3o1sMcOM+m5fSw8nnBKh+kU3H9I8BuVYviFezTGWFXo4/6F
7w5qc9jyG5XjNktf7Z36sGGHRg25p2lzznkjztQzjhSzBDg8ItchWE7XYrByEugCRzPj+bih2ucM
wjQ+gObvPA8RjcVN7us1ys5PFiUxfMiyYpdM4C/iGK9GZFfN8XvZs9ZssCSgvLf6aJrmaq2QvqQr
Wow+wrUsT1yFctOPr3hdZuEkC27EdQCdjvZ4QmI0NB3FfvAEYxDBasq58J78K8DQ4nLljfb5C2+N
wLLAArRUDj9R/OvBp7UmuuoclCZq6TWhaCOuwlR1JxnGDRMRl7o3ZWvGhAk19/P4GTlND15pZFQm
MqVgCSZzTDZpAI6+/FZcNjMww0JEFmGiWtB5vFT9ohwV5JaWO92wgB7P5P0MCNtrGJUrl6PCYrAT
F5wbojN6OAXs2DBhL77LT0jtMhxlCTrhiEcUDsBGHHMWUU9tgmzWWN77g1vgHEU0FuU3ZfvXQkMV
6XzMeYzq/d8LJGK9xmMVfpY/HF/ZjC8IunAxas/OB1UNjoLCbwTSknTNphkjyeBVfPZrX89svnmx
IyVWrsDYTkd3Xx5Vjh6S9Sg5mIdOtI63yrvU5JuV7j8gdC9Uwlkb0YJ6979P8dG8pGXikMn3kACl
A+jB/OY8r/ed3zwRtBPFPD0HfH6+gpMfWwIDSviucUFthqe+6a8Qts9o5Ka7wEeB4AWLr/qRY2s7
Uc2AYvqjCl+ErdG4psDwe3goAeYxwCBY4F8iyaQy6q0y2t/bmjvG/TLGfGGI7vkEBO8VWB2iernK
4x3BWK4eBEgOs50wi2RmCgfU6pVmWcH7hKuUN8BPa8yuV0pTyLffUv97ulPUm4fvuHzxMp6P7Hiz
NbVSbqMcz3WCLD3/nG4AhXdHZV40/+MJ3TiBpXTCxMDBD/o1LSmQ6kdT+17lmbNE4GhYnSyMyd5p
z7RtEeJwSw2xusoF8/UsMOHvv7vkwpENByPG2P0zrpXM6owr6GlY116DDVSyg+u6O8/bjQDlJFMq
B0i5/n02FOgIdyc/aRz4XrOZyd6vRqalpy5fbNlZ6QmKZNWREv16+M5cM7N1nqVLKel7kuhPdhqP
dgo55NGxB+kGq5U1NZwOwzQNP8/nctxNr9J5czkdjB3woSNpdA1kjXk8KPnQ1zEK+oqnJRGGlDzq
MpvWAoeWr0CvWpO5EsVC3IstiS6US/G1pdC7OpeLVfYgWGVzSINZ+r6HVtMIsDgkzcyppn9jhqf1
PDgOKYHQggD9k83+M0mctdrfYy95EO3Qq2uGXQEvd6NyMD0hl/LG2lRcdmTzcoCdcWPSqWqxqS0w
NQ6UwCENEWB8ySK/v+VduzOa1+SeO7VEUZN1cgyBqeV3ePlr17eHlZarXkxLCftEaTH7Po4cWLLH
WwIu7znYL0WHR4RbbtEUax5L1HdVjQ9JP+PVLtqsw1l08ez6C3HjoEhZI8RFcFZk9xkh2m1A+xgu
wNo4IHqAn/JooD2ODqXwdoPvMqrn3cLlyXGrPbDVRgnacgWh0TN+9May7Yx0N19Lfgm72qR18oIi
04jXaUDf9PdvULW9dYGVoUMQKVjku3kUzW+8waA6geNT4Zp0vCpTD3lp6hxhAE9/pXpizraXi/D+
Lu8bsfNwKKgiu2Akux3ljXRVuyvlIhTQNUgDTZ7Gm1eYZf65Nlcnh4rKhNfnziVHiHv0PIEg6I9O
TQwHa2a215Xp3eS9Q1iFDLpUK7grihrjAet9wPdO5DSoerUX2K1CtQJuY/lNm1U+ns0vIi4DbNCf
xIl4Y1fZWMycp7dP+L7s+01Cw3tYg30jS66a6mWivc0Y9e1sUIGV9QWdhnkIsakyv744AF6bKbLn
Ayi5bFlr0M+PJEfJaOOsnnuIUsd2SimCnklf5eADxJzJ8KosrIj/Os3A2RViU7hVfbanANse/Kao
ALDo03vG8vdh7gh9TgqpX9q8w16cFiRGh/Dc7smK3UboCh9f53aXgHl7zomt2/FAsbkJ7tnBNZh7
p9thVfBnsEODqCFOP9zD/LBLwVdRf65v5MwMc4r/4XRAOmqNDDI69yKZwmKls4mHiqueqi2vnEoL
tsxdoL8pMqUCOWqjyQ/rlVCXGrSajsQc+Ir4BvB3zyiwXPLImSCLQk6AWzlzspd8HqVy17U6LpQI
XfrzVUUAiXe/iOp5UXU6q7nCAcStaoF9RUzU5D7dLtc4ei/ITJxrhDKFqPkmAwcvB/LoSGqN0Awh
W0M3fH4uqn2/UTIJyT14Z70k8YzUQvWr3a+exFVVlq2Bj4lHGixrH5edYjXbkhUZkwJ8pRLYHFLR
/E5inCToqUvI+B/qz+DqtNxBYN7CW9Vythf44H0AXyGhZ++czCywqr1UfcJNQB/4Z25VhH6MFkjA
iZphLHtVcd2zGt7a2jbLzg3IaOkiRolhURIUru6veStADg+f0bzdXiptdVcxx+5RN4RJrJ9ra8Az
5len+ETvevBJwkETCcIKkJ3KKwc8q/h2keBzb3SKX7/lRwDdreB/K9XHNaLW/4lS3UM4RHhn1TlM
IB5dDVft1p4Z6k9VLveDn1QxY7BhrKEsiVQssyQ2OZyBiQeRRoFtSl8svmT7yErpVMWHhZDinUio
W5QyhcboNxbMt6oKfYRQfYzcZYMBxtLlMnV1+O9h588768YXYLF32UuUvUBcD69cFO/YwUtCepCf
ueZqicA29WlWzBljdo/yPt1ed08UBpaZskwdkNkG7VvXrLXuVZCLPiC0UbxdrgQvdP4Ulkgbux5U
wC9ro93saSQlm72Go8LSZ33UYDiMzkYYl3aGYldsSPoMH5alcUVcuvN/H1MQdzHzeMTB9Rmh+R4a
30CZYP9YUqmKokFUbevsGjMt/LHin5Drv8bgVXBbslBaHkwU3hHHAEnHN1OrmOy+/7EejSQMOpix
mpw7X6kuAM7ETjfOj8OxnRZJfnrxR4NpxAouxPHJ1yCiuT1V8umNSrNSv91d/8dwGz7/IltF4dsO
fhXYCi8RgclQ5R+ouUx8DVnSDUzXi4+UW/L0hB/FHjO+5w/TlbWdXWF8bLLYmNslXF6oBa30cZNL
nwrMjlCpCL74qHj9iiJHU1MpCvtFEE+adX68fLRTy0LJ0YWI0/v1Vl8lbopfKA+PnixKdou/ZT5y
Qdmxt8DBH8JeBJV2ixQZEcWZmvI/ivxmzcj85mxIId2afNz5PVhT7mQ794X3nrF+XTUoUGT2qgwU
gbb1oKxJIavDe30XxoJZtGJEJ85thWpTeSFxWtOHBtVIFRLUsl+uXXpHv2zRB5xatFmODbxAZJqO
cWOXZmVLG4iIKId+gswK2DCvIFbrHlS7o0UJcFO54IvJ2W8BFFE+jfSfV5oETvJz+4PyAeEh3Fw+
1J3LU+oN+JtHGA0JaXe1uZUML8qjAvysmDe6H0YDgjCLjmpYAeMNwP9sCxy6iJvK6ikaLzD9YpiM
V/Dfv+/fopMvUgOrvxaXQm+OSVng/2dTQVLHqIEmpqc9YbWiuHXbRiEptZQGXLe7t89dwH8I7syz
UIlnfvAKEIrge7LMJ8lQ6t8Vr3yGn72a98vQc4EaXIYzM/exwOy3KixrsxdJ1+tRSRpQ/VdTp89Q
lxwKTNiB+uY+fuD10h7hFLqost3NkFmOtS2xtDcZAc30bfTunsZvUlgBoKlylMtOFR+qJpOzCdL6
iZ69Z6jbcGUwMvJ9lVpJ6RFDtla2s+sdyiXpENE4VaCqtypXsiL6I6KM1WiT7zdjQlqWJtFKEjOn
efF8z2MG3bmpZ8+XHXmhR8sjnBlrxVJc2y9dsL4BUhMp36f4BkpyhhhbZWhwNHJiwxrQ4bTqK7GU
GHLBb5yuWDTGCR71wVE+O1Sg2wP+6yrclbjpTN0tE/UVWyfNGGUoaxJBjCapcu7YlTIupyHoKvb0
U935Cb9tHvCEv0fgW/mPuUKvOUAqyHDXNVwLdTQsbH0unIBqne6elx5npbfJruwGG5NljDhG8IIw
lUOxcH0XTMQ5s35Cc3tOVxFScPGhGnqLNVJbKjH26zzbrzdkn159af6zGjB9lvY1rW2yqfPBqnEm
N2OoaYc+HSGWGXajRNwUzbpqRDqJZCaICJQFibwWmx6PrK1/459KnKDJqgSFO3qjy6FMhk73pM4l
oDw+cPkW9FjRzJ8GMW0JgVzK1dZG8qnDPUXAgsOC0p6qrHpGphvDet4OWPK4jayztgHcQl6NdWw/
mU4r2QOPrn1fYFDx8uv1RIgwOzpSPMic0VJSmU63YO67YID1L2ptgtjwcENgm1fuxdABSznyfzVf
iBR4bVTaqX2tydM3v3NIVrGMi4/yYHbChKVfLg0H5pufFh6TAGMzoUdvvIUG/7WS7GBAvs4FUF0T
XXSN6JZU8IWJ1oo0mCQ4SpbtTELbn2JDQLdw8Wj0XbvOLPPvNvxjzP7wOKk1P4VuhgcKUWd5R3QW
jJhD1gYBo65Fml3+MwwZl/RaFQprbdr0sx2GMOUZp4Fm1ClGLuMAICgZdf33TE5aZImv36Zixok9
I7n9CPTnQunZ+wronc0XDNIEi6S+Qy7U0sAYxpdJhgGjVBDFjiQIIzAEajWZC7N/SXUeNrU1WswY
NcYH1U12oaRDlwWSB0a9B4OTC5/LrEiFYe/DyxmIIbvJej15sYNiYcr22TUfOE2jGQ+naxX/iooO
xY0JCqih7chE7heKcrwxEb64TPak7atd3wa3VTWZgy3nYkPvZytbR3tpuNwzpKTYi3l2l9sFPXnE
mtgXjFjFg21IdSZNDW+5ZKAfUIM9rLUajanTzOf4ApFvkjr+swGSVFmSAnIa9NVb2+amRTPGAk1f
yrzFmRA0UAIfSSnCqTw8pXCfpogOc0j83ygf7G7VEya5U8hcAgEsQzOIBiJ94gk17thicodwv5/N
pwqCY4Qw8k3jNwnMRVd/XNAsK9bmb5LjW7vqmCrMshPmuLARJJrKFGWxBSckfWW0pvSG73SOq/2w
XXboR5Q8iQjTgDwMc3DocL2YXs5oh27d7u+Y91KOQ2jXeFNV0+rB0bhl63E6FdtWBGnoAR7zAAew
U3tRadxmnGFpjez+t3E6GacdeceB75YkqWEeT5YTcl6AYFjbwOQRI+UkhxZOaHx1IWmY3baBzwPZ
YrQf1b0E0xRDQnS7oW7EGZ42XW1jy4EBTcxZdEnMSLk+T+0z4T4C0ESdzvtGMTtO6BaUmI4SqPyk
jSmc6h4vxbzwJGJY3btuekTko8iysU67SgSucCOQ/2JeuJjCJcaq2L3T4WwMxYi3FMj3ezlnh82C
GovOcnoXTfHcNwkFK6XkLI/eognKdvdOZsgX4F1mSxynX7IYQgD8t1k8U4CrNtgACPargHuR/7yI
/6h5hIbxQOWgN5tcgwIKSsHwwLUjhwrtgJO5m9R35I1rmUg2CBRyPsSK6xqzn82LvORSLDzaT/H1
Ray8hEJSemu9E5KJSQNM7HS1txssNQc+dTlsj++Yx8quysS4PdN5xf8bRcgat7kg1KmXVL+hkvc+
fhTwQF+D1bWavWBQraEmrn8yxbc5B7eXr25bK1h6ST5wJPgLiG++u7xOuUrJ3sHfrFAKz4uGMreP
d0v+lwzNpSOuqxYbfweNP10CblLBnlaAJXe7G1dGvTRF0E+RFN8qGoGqhDDULgBj1x+er1MUPtz3
5xNe2e7MXsq/vmA9GPrY9bK2R1e2i5oaRjMR0vvytrFbmF/M399tWLb8ZtQc1GtsNbGxGtkeD8kF
fq/ObJxo/39xBGRqQxpj9ksExG1DCtopZOVKX4IBW7+O/U9uQ4s/vrIfJIH/Uv9ZCrVjRIScfJaK
oBoKns7Ene+TFrmvY/RQK+IlMaPo6uVcwYtZj2VqXepb8WGdJ1mRE8wljbQPMSYUWgO63ao6B17D
dzUHIcB8jZ03L7in4E+FnT56dW/bIx6hSf8xdMtc6ePjGvNmCws4KJaiyeydHDfcgzgXvp6shKNm
WaBjqnfTPlcM5Gz6FBHw98rbuE8pBiN4WVQJkqk7ww7Ea0OF42BUGSStb++trBMznUmFzVhEHuXp
HS1vmgb0wluKfx2XDRZxgQj3O6158L6yKnyAZLR+uybOxbCzLuxcOdVFaJaMWlra7fJGYN1XrBq2
WIztduJGg6FLq0HK5HaLZAgaxVbAAaiwmYvd+2yBZV05ie8JwWLt6PUoIs1BjLY41nhXnlAjdJR+
ptolRI9EMs84h3XUtgjwG5mTycfUWy/RVxIQ2y5P0repaYxch0IlFL/SK/UaleEJd0GWMFtp7je+
5jGT1o9WdlxYDV96w3H5B+HflB0h+fzWSuxC/FRDmu063IUkFca/1TdhQKk/8mRCHw0b5rNDhZ3x
N81jAuU6zrwGzBYfa0G7Srf99lOyEwlF5JxDuTaYe8EUOlrmxrMyizlvqW2ya2RDPx3w5pgKOS4Y
0bvIxg6PvwgOlS7BOd9752XVocZMS7wNVt3eJXv/5N8WbXfHXS03Ml2lY2JjMf/9aUbXKG2lsAh7
OXcOmxPobfbqKHNIjRFO+o/PIU/aK4L2p8+aBEJL4mmRt3EdlYZ0Sv7wRPMLVbxqsQiOKbeXff5i
ITlfDvfLMK+gWFeRTkcK0ea9sMJwBwrhjaG4JeCDvdZtk43ezfeP9mWppPopLxBr09MppfhwsSth
TE55POdFepipwVzV5jiJ0ARS4I2uu9lNdcJz1oTDvwLJikOhPbDLmP0jEhHuBjlY2rQrrB9L8CRe
p/GhqbyPzt4YfeVmNv2q3kJ5HedFhOI6be80fRKYc8JOnYmagNTTFtILM+fLWa0AZMeffFapoEGE
iK0Hb6vMozFWxBJ0vYchPouXnkdtUZoheKUqONq2oNE0ckKJhMTQVjWviFbro/vDdEdCJk+8GgeG
awJ7+FDxTJ3fkyDOL2sN0ro96j9Hom0SG+R7V0XhReb5KMqXLc2JTtgZvJdZNyiIRLU0chvDMi2A
HDJ79ce/zEIgOmJrzs4FWSuwPYpvGD3hTGnm1TTXErj3fIv83SjtE36WGH67z5rDuf4Bv25HYx/V
PMxqK8U7VlzdGi2fIVY7v9b81fn2XvlgwK3dklRpZp4r4GAiQ8DbbJAUNFyc9pMVkDN5WukrmBxE
xXJSy+N2mOug9pjZJwxM9G2oeuAFFK3IvSNrIChKTq6AQFJi362AIgxBbHNlIuecLcX/rCL1oQ7C
0cIORfY+jPfFxYMyaOPJrF7w2wo8NxRTWwdLkdd4uUQn743VXrTSGZtOUSnwuabV/8cOAfG7esVw
fGbYLpJfxDBFQpNaYfzv1yKtBV6JbRTXJl8jY4/YkTWYevkJ/EAc7ARC6TXcJUi2TYyC043Z1bvR
qAr+W/zV5AJdCOydqHHIOTezrM7y3/BcxsqRudV3/HXPMEhaqwbTQamO6y4YlJPBImTiIt6f0efK
Z1ybtR4JSjOIWwYXzEWCj5AbY5i+Rb0hwEkIZOa80qgVQ06nPZvjkXdEkP77vT++zqblQOnjVoa6
AUN/xYoTiqolL6pcc2cSp0O6fUh673ki5Tb+6AUbJR1BNZjAwNkstqrmBpKQuEiBNikvlCfoJJMr
1NTMsCtWhBvyqgMJ0KKuu8OaxfK2jgKXmoZ0dBSLw6BVLkbKDF1a8VV5JNUpab+ws+09FQQVePb9
dvGYTATN3EkUUG9MJ66s3u5zXVF82xySzDO/oJbiiQn/2i2OsaYxmk63h6G0r72vCNaj72E0aIQ5
qt2zlNqggsLYB03zBRl1PxC1UZy7a1hW0jXdg/TtXkEqwzqP1DuVhSaOlKwF03hapuCZXXHsqvzV
CGPAcT3IWMf03ghYBVyhNYTX4UVbkblQsSL5KA432xsktAdG0mM3wrjX4YOFCv+vACzh3kO+8QjN
ZampS03k8fB10AaM2nGLeTUV+SOSSncLVSP2ViQkcQyuyaQsSZ4w7LchxUMd25uPdmYW8yz0A37T
OAajvnEbM+AlyKSz2oMqWbEu5sTSdcxR5UTN6fqcbIko2JHeGRHDXqu2swL1Q/+jtRWEJmqcxP4Y
0XMFZRQzd8Dm5CjmlUyyikxBAFiS1DLAv9E2IDSpVvONDRWICX5xWutoKVl7J3Ck6B8NQ4JCOdSn
viCtPmjd3jFGWN/50YmKUgBnPuS8xERHK/VqUTfF/PeaRTGkdsXwa46/BsC2PRoafv5mhaJaAFF7
lks+USmlQh1mElGWSAFpvATxgAjk08kB6LWuHE3AEBcCahBZV0earaO5g4c/V3KbjgqHRsjtFkyj
rURRrJMxhg39NaYaf+2APq55irQ5TY8oNgI1dGWhZ5qMs1ocnB3GYQgZxYhaQc593Z9jf5iQZWym
tKalIDgU3+8YZme7IdiSvEl1x5sthKGKfDl4046C8uvSppM3J7O0L6hJ6MSbxdYbb65RT0vecy2j
qZ6uDTUGFqhgMx2kvbAL4G9nFkRL5ykziwujvQxCsfEpuQ63m2BSDunoiJZp24MPtNJ4daQJ/yEk
K/1m+1XaCBvW0/AboCHyuZGahuSIKPcwalTv7San6f7kx8RhvE7cEyNbvBD1kLlTzhlCRWCyswiG
NKZdAeBn7i4aIR8A5us+Mgyk8OibWCWPKQxuEq48zbWe3z7RsBGqF9WriJK3PXh79ZXHuzdbXoFx
wWhJlnAmo4Scun9BkgC9jaDMnrHemVUibOt9itERKpnLEkUd2Gl6wHF7m5IMPAnSeMoGHbDbiLiS
C40UwIs33mnZdEiUc4A18d1NZO6r+XQUn7DasomTBN7Uj+7KVMO9knzVVOXuWkv5efqIrYhkrQMj
GYkz5JvaryIRXD1CjHM/+M/pf8eAf7iLUz0zeUUxb+oUoYWSiDoe7tWVMH3tao+bTntDgd5MWvH2
sdtl5Gi3mru4eYCn69BGH6u/7PaEKRXQ6P55LXJRO6z6a1BXkW204qV/q/3KA1IdsmMywPHg0dD5
1M/H4DeL8731hIyXLEPw/ujO25mr3I5LGwwFH/2+F2AqnKxH3UiFhLjjHzECs+63hzJhq1gmty5A
ITOKW6JNp5fz6CTd8iiGUdZPa9sXvLWH24h/P6WkgGDCqcehJhMiKuSdT2Izgn5naaz81lIKU4n8
Pdu0bqeJJZQObAlkkZMyBeu808tJD4mCKPX4sSDz2MVa4G+zPHTIwa3yI6PzlBVfMKgfYtqDzUzF
RSGassZuSVXr0SCRytYMQukqnTJtIkgwBBrNB11TWfkn94yyPsn7+OviebT1TnCt6hW09dNH9vxY
OfHKTabtotxu8+xolwmaAt4KNhQscRzIO1lhUs0YTumw02SqQ0HS66ZfBx8DCcwCozUhzmordVvZ
Xl+pbpVwNoEI06sMJp1WlHkxNFWyIa1874ciAwkq8kZHcoWWbiLJDWm8kLcoQns0kVRVVS8jw9bL
IAr7K4DPQx66yANkahCGeV7WpmYS75nwAB3IW3mMI2TRVBBVOZhwmUvDxevDRR1uUx9HLyp7PApT
7JOPGEX6cRjigUQKIN315iYCo6SGloK6VqLHfKX7TTwtd6mw2i4eRO1aqUcMiWA0f+2jSM8T3zvf
7MTuuPzsh3NvUd2n+EC/Y7nlMx35UrVdBOEXwdJC+Ol7l3Ih+0rvB+Zd0dPb6qj8Og1QyDpzKjPw
f1Wlsm1iY7Xxn0QFcb2rZw0dtohCnyDB6mcWNpZ3bG29F8jIfaayxtO6A5cDSZrrDvYVU4BgpeJr
Y9BXtETN5EH7oIh2LHLRyq1RmuULXVfEgG5lc+8264BGBDHzfFeF6vYRJv2UJBi64YUAcGebWbfb
IVQmgbTpnNktSOSzGdELqaBoLtrQ01gH6OSPkFQ4WnD+czPVss6xIdmYDBGwDdkCMLwskY4pDwvN
m42lLQjUUirlcR3XJQqBJjneNK7qVnT5u9lUY3dEKZvttmntgvfktvlCb5qD1uUck9Zmf67didDz
RzEhA2NSJH0TEqqghhVFpOPrMBW9d1evajC/CL1BeNXviWP7zOYohic8vChA+X0D0HgbxnHJ9m1c
BIUXaYCZe8aVgNH07aBXaDI7NtD6DwUN4KCG2Ej7Qs8mT817ph0+28wepIgo4EZ8KmbWzwigfWHj
UvjNgvOcdIbqrzY4Ri9d13dNvZxbsv2N7a5Y2utMHdSb+JpIM1ubkGjPvCKc+Op8ciYaVD4LdaHV
qrNaPDKO20LTssB3ffodOfYaCr73T01HcNWo8tzluvSctNR9XzgbAcr76OQ3AfaiI4MkHU65kfn1
BmRJ70QdGECv/x4/VUy/Hq7l3S2UjbinY9PTpnzDyDewumDe5zBAJxCBbEjjozMlJwT7rD63HmZp
1C6KsQ5PBYMudP7e9DdBL6/HLPBX/xyUCMPSFibcdFmY6GKNuK0t8Ejwq1toMpVLuMcC+xCGh6Rk
zwRhMvYR3EDoAVlaX7WAkZKD0BSyF3p5TjYDKdiFylVfEv2/wyaIlQFKCGanuL3U23UvZknzzkxz
NRBjemoJ1PEY8tfM4jRFY2heO/RlusCiAQEgXIMrtyRO1t47Db+pknJIMI/uIulRADHWHiL8T/ng
xDQ5sT6FoDoBy6eDUGgxBSzeX10e7AjoEJXRVViQvMobtwMCLKra1dH7GGmfdzSTNImCkzJhV8wG
jJFUTCMsj/qTWQ7QUYVSxVxqJsIby/ZY3cwqafIA/8MDEXJz8JNhj/ssPk7wibg5aeYbkkgTW/Zq
lW/jCCBZgr7d3O7aInVRWhGlDjVgXry+W5qsoNJyIQ8KdYapjUfLl0va10/DWjYTTUT8rXlX2dqU
w1tI9aYCTrvaQi/Q/VcQBb1Ag4yIXE8X3M54oYTfbJB7afV6ynob1AMciJp9yacHzeH1FyMOogCh
3jAFxjHdGoW+1gllWNMjewGWhA+6p5BQEARnmkXUHu1YlKM1zExTvoYfnN0P8RMv3y5/ZQrMQ0zI
1IRG6AMxmt6mZZPJj4a7EOmvQBChHoLiWlFDbK5tvHKd6m3+HCOU3nGSmCSznHqcjiQIlS4bbf9A
ieThqvfAK2jiASxQ1jZJ+ZQX81hIIGQu3RG2Gm8lcjOZETfb0M9jsWE3eb7zyQgxCieUbjqN3nY7
NyPRlAC4clzJ4I09B9sH9NlvlmHLwS0tnAHCk0g9VqFlD81xKTM0aNu5Usu046A34+1pFCazyHxu
rSA5NC+Xi/v46sDFIY6+d6sWrWEiyky1qDqcT3WKIIv3rG5wX2plRqNnXbj3VYI+1WoBkLhaOw6m
2c8cX1paTxV5yuBmHnAxPbawSuzAZR83MtyB9TM8p1WG0jY63gng/gwKNtoL6hgb0bzUEBrK8v+y
LHjl4iBoWz5LBijdbKG+dGn1+HfZ5ZfcyrHAhcgJHb+oRc3eFfwp7JYSHaFjIhG35GQbur//4/zd
nwEABvRFuW47c6j8aWmXF0YdUFelKtpDR6gsm1KifUDeSlRPLConFIVxS6vvfXTABkBKvbBny9Ai
WSDudjWxMEkT4HrAJL700h1ssZyNwfn2etWNTzV0FAidLhIVBBofJlSaRHAIs2tWgxN4PRx8KOI0
MtK8ZkWTPU1iXVrn/lXAGfszqOYktDmaHvQT8p7WgF2gUmEQ5GGk4/I1B6AWYXpSkEvkb8uR8kIV
IGdcpPRgfRmOoHkzuksj/KegBEUA0Vh5lcKZ93dkLao2nOFVbkSUg+yT+ZcTIsNLjAihIWvajSCB
izUBg6RMwnh0LQckyZZPMm8EH37/jtQB2OPe7J17m6Nn5Aq3cL2m1+QNOwVCHSBqtPwXE2rJZ+U2
ACLjmaZEVAUPBnW8uu6A8fkn8jr0luWvMzQvsQCGWY3h4L3lIuLheWjBJW2XH+EGYJcVK0pUaXmq
/QJKoIcQ8a4BbbEabcz94oyEmGAnC/ZA5FqM81FGmhUmBSlwJso7xrRxPVz5JuTZKgn1ktkwSOrg
asyEeUuoYWNk5Ld0C+BnR/10LKux476S+ojupvUAo+D/c/Ee9Obx2Px2a8f749Tb+uT8uYnOR0S9
h3lyCJ4IbcRsoNZfevsH1da1x6NgfjhmRMKsTnh7720bv+T6qkCWD58PpWw7crDDUkkghkXQWDfJ
kjnRKgyc5MNepyeew8MNt0eHVHDTCGx7sstG8mi9QH3CF24Y+HyS3n4nFRB1kOZ619lt8BKjbcpk
jFFU+fp3KADQx+F3FLsANi7eK/pQOaF5QTHFPgVirFnsi/Ea/bqA9UENlqawnewVFCW/+nps31zU
MrrUv6NDvT+SoRow0uNhx8Q0pZAEeCNJAa8pOS849TLRVkyhMYBmGe7YDD04LpjC+oNU1rHlHGx2
b/iyJyHBkEMExB8/RV11dWcpSX5Yo+t8ESh0QNsEIq6CmXus/V+MNknsTQ5kTbOZPoqyrkk7Q4K/
v6EObDHFMkkZf9S77PGwQm2rWEbLcTqZn3oKlzfgT7AuJgxDTGlL+97hun4qkC5AZMDw4aXzf8iQ
61DYmwOYngu9eekafm+fWbJq0xObkYOhsnxKT8T7zETv57cCMF6eXmNsHLT+yhUu8auS/nBrcaBk
Ekg18cTUsN7TKmmIhbnCvMXXXS/szscUk3WD3p0/x4hAc4ouc4GDI03iPzutXsmdsCItHyeZBP8r
dtSbnLhBVQ26mhNOOEa1sOu1KeaWgrgVsOKni6+yLj/O6RyoLMZU1G3c8Od03e+I+K/7XeC8grH6
DHGLLwtFnZvS82dV4R3nnlvzQsYsWntfLTRVnViriUr2vl1I2Iy5l58OZ9RqzOCIBTXjRlZO6xEi
x565Dz0aLMGBpq/HciIIfxKzfBn2MBzN6tj9IZQkYZrZgooLyTVYF48sK/XmkzqkifcvbvkJtDgx
+/dp5Jk5K/S9v70mxJfpiqkxlBv3rxeS8SDi231pw1r+S72bUoxXIQc4CkotiQIUXItojY0aq5wW
tfjGX0i1kN4WWayCjb1lYX2BYmXQNRwDy4lU13bnoskKdwRfMoBYGKST4IygWBytde8XF6AEuR0X
iv4dO2mCwDU45ERCx4KBWHV4+bJPr/v3EWG+cpVPNE+5mAXXr38xrQcYsg+GpuBy2hLMhp6F8iac
5dXsqwpf87KkxTT58JrN4SCugYwiYx6odp7cohFAMtxd0NlWKbz/jkxMBGkeUrJMAAkJ6z64vc8s
lfKVGo8l1pCZLh5+2VwQTltp/kVMGuyYrQvCCistoW8SDUnpikkjWsaLBffobQgck53ytSex4YLe
1bMoim30lrPnECs1pLOwNzbZ0DS2vaEcBeRWutIBXxW/UEaj58eI1dB5+ryYQcVwUWek2vKMTGn3
vgiBj8VHwAIDcagKMuWUyx6zLad6GXUn3WGBjwSUP677JdkX0ndRxra4r436moz8q2KhK/mU9Cjf
4ir3+Qurrfd5c5L/97AZF/AiV4PHMsgahJBmUMm/Rcq9IskCyAC/ExonXS6Umj8s5g2+q7NPxP/B
PMvPF0+hC58lhGI4rjbjxWqA0m9IYu/wXK58rGZ2k5Oag9g58XjXCzoeZqSEFgrga6FwCa9j/210
lfvXeomlTsEutTTMl3vyyi3AaAbWnrq90JXOv2xj1yYmNprz1570RIj0z5WYBPealIjH3NR5CPVQ
V0rGz7WML74x0nmKnFI1hFJMnWpb1I3TLxOOEr00KYEH9L7neY+pOvP8xS9A/EFC7C1/SakD/LzS
sI/IKI7dECPLxOUcDTF4HEVT012qfcDuwwzGhbH4G0PiaYyLK2MNDcHRvpk3I3cPiLwffDsMFL47
7FKZMgZ3jXxOxNZDWQzoE7B+MbA8B2/xP3UzSRBETdVmJJP8h0H0jkbYiAGRcB8VGMoPhAaaxq8y
7VNTAinW4eqk0347+G+V+PPpdvFfFE9MsBV6sU1I7dazGD5x0dnyUq14KBB6qVZfa1dvzgx8Jyg/
vHUDCsM4qX7V/YB3OuO/CIUsvxGXJK5DrgNTTu1uIIgABnO3F2VSHb5MbIFtxCROINhFItPCc1Fk
b4D93hh9Fuewap6+q6OH1Q0ULAuuZnLHyiwyBxcdKy1TE7MAmiqPJgAmEYfwDnFDx9QyFiQq+FUt
qkRw/AlKkiUYnTxHUZqy42pMLq26grLL4NwpRLW7MSzylo82tkeW1F39YRjNusjLHMHhy7vLHBM4
z5roDLWBnSzPZ06J0q7F9XRe9kToCrS9zZJzUjTtb55noGFQZeBC57EuOp+DEVgFkOyUHsMtkSvC
hRf1Mf9TWx/7GaljdbxOGKUmSytvBEq+ikrnQV9cIY9fnkYczYEYUvwjwt0qifw3jHQfvUlv46tl
p2cIHTxLv216dFRAI09bXsBStaKVZXqQnkkER+BQuNAU2jr//A4HEripZXN1HlNMhYEVLM81d2rN
LIUiVEs1DNU22nCBsXu+pD35nxUXePYVeo2kZ3Iaf+iqnG8040fWnn8Ix2mImJiDsmWQFrzz0kEE
XJQ+cQdIAnj/ddBG7YKuN+UmC1Zz7Rhq4QzKtqmIz/82KCr8Yd+0hUTmw5us4CAY3zVRF9xMHyDw
eKJpHGWfdecvNm7iL7xnAuFr3Cy1ie45kWgn8fGf0XL8VSK37MsMWTUyydSlvxVDcvVGjGulRjGb
dCW6a5VReCEpICWfS5nF3taUS3EXGwUkL2ReLZJ6TKxblUmgEypqdNNSWXvF3meaF5U2rLZ3b24f
2exnbV+QAe3ALYocDqQw6WeGd6RDLZlY8fkVsOefyf/99DNePoAV5xSZO4tubsBBcdPcsrUozGyA
P1YyK2MsMyIsjio8qjN6QoTKCSjtWOy1FJKjzz/RxoJ71BYXdQiFROV3+gVs47ZrJgtL/IoUhA5S
p++m5x/j80uBt3+MEWbG0K3k+D3xCwLOx4YgUO5OhsOXQZrrbB94bTcMGgP96jqjXt2Sj7YkdgSZ
JifLZ8w15rvSKLlPU71WABzFjMNKeb6tB1lDpgsoNNqHleUHJgzQvbOaRLFrDY+lL/5uDB4n79Ge
+fKbJk1H8PU4YKRvCm9Hm1otWtyXr4rWZhwV0dxrA0PoTUUehdcgweOzbYAwwpAW2dTf8NddJwp6
9YzkF9yTfPmwUnrUcomhcircn3/j+zDcVXa/Mn0wV8335eD/8e65Fy99EYsDqQsfQRzb8tLmN/e1
gdBtWjqShQkgNcQV7r5FinxubbZ0RAkj12/KxJ3Vg9DsJ15LeaOukTcCxuHq/P5xtv7CyuCFsFpC
B+6Bt+RkzyWP6w0QU+eCV5H8hJCpuI5ITIQo0IOGKpxi20uPBQoLkl0zylUIbv5N9N+WM7Ntnonp
2coFbiSaiYN7VfzObCotN9oKD0s5IbJZ/WtqvJhionUsrDHoKBz+nOSBipJet9X7Y4gY4Ckohy0Y
b1iQ8w31/onw0WeH5fJSSYFJONnQ5TN0Vzu3Qk2OL1tVMJlTaHNhNzzujvXpG+wYGrQMxKmn2VUF
Ll9sI3tlHABtXru/0SdokKkdoBJ6DJmBCbZQmhvNVC/shxM5SvqXeEcvST5A0nVxAOD8nRPaSxQm
XfuaJcTekLf5zIG0UnQWjcFpxAzszBBzuCIVMe3Ycrk2SIHDrw9PpoWyNyQ/bzk4pC4yVhCi5uIL
VufgbzrRARV591RzJqNE/mo8pkuWQEWhsD1cK72lUNpBgC2yljNXAFuH4dDOfGcX1ApgvdKYIbNK
sa6I5k+1NXiCedFyhZPQnDoKe9DsIh1gmT6FXYVWBthci6Zmf0cLTwntldQjgILC2ThchVWTQ0pw
hCEmNpbFBYRSn+1/+OQiOJ/CDruGyeMBggg50xYfc65lhmDVOGtsTmRR3lfHBlCV2/jq/z/KSOhU
4bU6hrHUX7NdoNWC483/mkS36mq8vZnAPQDjL+N/fpCSNTR8ewafg+3zMMzpdmbt372VNcvwXO9C
LhjpV5JBzySwk6xxsrW/pR56ItEJgtm7J44hsxHX/FFZsnNLs4Q2+P8HlrPKSvO3UiWT79u/KTpY
H6bJq9TvN/cblBFGGecBEz9VfHe+3Zov6n+fm3F0bLhfGfm9wjE50wlHGpHGu+ZOHy39oH6gBrMl
V16hac+qY+zawGqKfH4cbFckQgyl0QHzV0Tbf5npo/k3MjZnFPOQwFovJNaxMtoq0fy/50B/B/rL
6iBowFQlsE+evF9YUpYkpVfsEviwARcPyjDP1cgujtwvnHaZxbaGXeF0I1yEgoOw1vOZvX3HM62b
w/eaEzhQcOPvGHbal32z81/s30z89MFMEgop7COEFOMrmSSauA6NgjMxGge5UJ9VdsjIkKGo2XXM
qGSVeNB60WLD+faINPA1zjUL84gWyOlHEbKluVd8eYKWhJBSM0nJ37k++Z9tT1bzTxNkH26bLwqB
6bcnb2EFet9fsQcMrBgyvq7QvOTmVxwStfoYLa0Y2A/tme66eqzkZ72r32ANo6mlzddGj7YJgFXb
Nt/ONEwpDnV5W4WKhnRsClvQP2Ez7GW2B7g49EOkQfcT0EfIlT1iHwmtcOr4+4F7JEHPloezwb5X
2J1C3a5jkEujMQe5NjnYRzMS1I3jM7Bo8SIrDwBea7tzENWwFp4FiuUwJlplIBVffUNf7cPb0q/f
7fxRNdly0LPBMQyGsepQCjBA5zLlK2vPdZMrgCXQ/aOfS2WQc2caSEAmH84KZSsgI89k/wWTLPLR
2u60bgwuQO/RweDqfH9rEfEEEXDXfd4dVm0hlbNUAXk28VGp14oaW00Hu04MVfBMLD36m0j38yPV
+RN1ApgCDVLC3tGBYFmlEtf8BFCar7j7fBMlcJQ4FQLBJLIbcT622p8UJVD9SzCoscJNruRIhHtY
a/H79hphaGQMHd2iSdWldvPptN4WnAoS5KtPmvGtkI+DT+e5tIB6/S0yWVKEDCdu4cfVBxmKe1j0
lBiMT0eId+u3qb86mPbquW/d7Nwc/HyRsIFWRjS2/honNyS80+rM0zelSRVovhRcDY2mnJSlYwCa
2lo59zcl893rVj/bzEl+CcOQ04YZ6Akz+z++RuMrkKdRtvLMposx11p8OPjS+YRqYlXHzgrw/ZRC
Snrh0ryskXrt6hn7I9jhihZzlh0wBI3xMw4a/ni8S9bGQaAF14MQx77iC/cDI+S0ElpUfAnduGLv
O1gkid+k3EzButXnG6L5z7yizRVdNUl5M6pWDrptkIrSgwTUo+MPheKTz4aR+Y6akxU1png6e1Tk
do+jvvYbSis2PvWrRW+lBL1IYrT0RqtnMzw3b1oQmSeL+AKjFu3TZe4ig7d5toP66JxzurjFwVny
squPuUPQhbkXqQ+xNV1J4X8C+HdJXKexn2p4nHtJHUHN1ZoBRcEJsZifSdOhJQ7pGQ1eks1ALb5l
dUBB07ojkDv57/3+kefSqIFUZYZbT1Dukq9VNnsaRcq1oDKqKYc02/X5o6XxJnk9UPP+yLQxU2Kt
DJjsfPQugaZRCUUVNSpBDd8I8ODPVC7QGvsob5Jsff82FcNiuhFMIaT88P2J0kUb1Z3SB88HDfF+
BonrMarqVldZPKIp5xLHl8nAADJLjn7fVmPZtk5etu4WOz5aNuF5TC3bShovYexF++UYVmaPMNNQ
jfBvFRoSZjtYKPdDzKDyCgQ1L9hccL7qT5ZVLP/PE9LnUsNHZX4x6fdpYmxmXpdmCQFpK8aMQvRI
OwZHElzDbGFB6r7/43AkoZTb+v3L19f5Q+keA/RU0IgDZ/qmdovkaoG7pef6oHWFAiKCwQ64sNcM
LP3XS3i9jMwWiMPJirDA+SbSi908YaXuVP2V0mjN1SyVz+WMMGVzqJcb3V38YhVx8WqFneNK4D7P
01Q0KOqOvBcHNQiaShtRu97JwcaBYqtwNZugHqVCMxrIYziIzi3TwLRdzTmBq0hpx2f2rfi9gQoC
SzhFqYgoSXzXLCG2WcpWGeaCELfzoeyPzeoLdUt4QesI+/85jRbPygI6qKcHRlYRueds6iGU+ixa
FEV6sWsAqcCaTN2AB/TFKDN21dQdn1lWayDeEEZupBJ8ohmmzprjjnPkKfioFlGdc5A2oijgIJGb
t/sFgR5SS2kIc1Fw3xUvPsZKJmTZzYeiXp/BRKuKVcXKlzbSPbGPcZF8/1D7fN/QqfswuvfPoez0
ekDiBBSxAcx+ltvuizN9pPldZaI2ttswnLMfE7uPFJi3D4FJ2ihnTOsGKo+qDY02EM82h64gte9B
IRjrnTE8bSeRGa/nEd1WYR4JEpwzf79LWNOs0FlsUY94sgJ2Yl44OHBsCqgVnGmGl7qJPddBs1pq
ju3CIV8F7QOVvqSSEL1b7JSnAlU2kiQFgarq6IMiHojjk0avrlVJDL5EHS1LA+B2IiR728DM3rmA
VH92MxT0N0MxRFA9RvOhksO5JwkQ3hLtoU1dqeYYcsfeJEzhYXGaY64FMMtxSYqhqRpyQPQ5HCQh
+jpQpyCBi2Nk/8n6eIs5yGCJ1AtZg62WE2bcQmnXaI9wFa2saJvFlYdwbluJC7yFwoTPp7pdw7W3
jYfDv3IGm51EO4mIReUfa0MMBEboXnutUiErFtrvXV1j/KDmUqLOEC4+xdXG9mV4ko2Ty8kGVVtN
DrHwOJLIPATKpGPGU00hFAJSvvaYI+pz1CgWq4gLG6Fk9vOj7jias1PpEiy68+t268TjwH+CzTKV
kk3uoFq75VtHNiV/1VfROaNq7iDFM4Zcu2QLcRAFHbs1CabIo1F+SMfVhtLVafVJ1w05ujDQJteZ
Ih9I2W5q+SYK+UFcYhV0ILygGwMEqUfzs/Dtr7VRNqB4PvPBQ3R41TU7te65gQwa51vkkTS2PyDt
OAY4PqUU7MMRrSOAswqB0HYLIzHNAp1xxocE4G915aqp7oBbo/3/18byxEnRGtO0NFWnGlJ89R++
0Eub9LmHueXPTfkAAVgwCB/f7+t0V4wLRaaGKJogsD8m3JVFQX6S46KDf93u9XvK3f2eca7jdze6
97KBGZCWgI6kOVJpDUjc6qMbviLw29S4w4Q1lVbytEPSspwD+8QdzshzrdeEo2k210isC0m0Acla
eWpewbeCBfnJzmKP1yckV6u3O4HGHTUQ/h5HjngJjnqm2GpCPuqltLmm4RFKVe5kkAJUVokAx3Kf
MXtvtAle+/wkpbO5tDIZsFXp8hm1shxHSjedyJTtt1FycGowcKAve25LPFNMqAWHW5ecjuafVN4R
onNXXzUSphecDH6kWTRdJJewsbKLAG4u7u793Cc6l/xC4LXgqdZbYn2u0dGBR9sOmtDpM24090BQ
TkQPPLu9Nw+MBmIgtsUmKB49Mj1ZvEC4Zc45fMGaL2wu5nOiH8RZ5hRBpEzg27saZDxFln4cMCaK
fXsfGEW/HqU1yQhxrlb7jHsmCHyG4WQPGT+LmYa5ol4WA1eW6E+iOVownhXQGxTPNps5+NBMORVX
sUoA6I0fVFG0238YmvZswrh85px7Z+V/F/wj1n9W8w7sjaO/LV0mKZ8eMCKs3z70FekbCdPh4XJ0
h7t2gnwu9AVOIBzc616WdhVpg9ZKJqamf2ddraqImbEG6LRlnAZkhjJ0/C9LE38VwKmIw1fogLeO
C7J/fMG/YQTg2Jvvgms08qZV1H6Awf6jQ6xbmCQUtEw6T8be2T8GBztKYDevDzKionqaolFRmWMg
9bjRAfU6PloLXa4eYpO5nQKnzuL0JYZ323cigh9lPvuf6braXJ671xx+XyJ5Q46r3pHN0A1BGTxm
PHUVUaQ8NrG1/bluNM86T3/U0VwZ55hS276yFgdmKMIa7IHsxqKDZqndIPj+nM7xw9g3H8nB3kh/
dG8Zq6ZNaEPsCfHLFHcjO5MTYeJOzu0kkjfKJzTzQMAl6kCNFHXNFtRBfKb9WVj/gF5UTwEq65w1
jnUofxnH547CO7JfoZY633dZif87cRYQGBOc6zNiJEyGjz52pnsNUqcHFPnpFqXwVSjGCvHwHYWd
9+PeukgUPPL79jKkuOWdoVeOvtVCEJ+uwkeY9/MPSSKdzPQfg5BQ1Rs6ApcveoGwE/m6lZ1LtbtM
IfyqIZji0yvvdlfOFcmzNfN0KAndkG1M1uZY8wTbhJuww5L5CSINmuFeD7DMw2r38q3iCgy9Nado
XEBlACERB8Ytnp0WKXI1l2+G5z91BHF8CPyZqKzmm79JC0roIfEb+R0bTrgvEA+mUtXyWhRwV7Kg
+XbiPtbSVdjRMwukQ8SHb2P2QUMUfiptTU3UoNSXxPFEq4IAtmT8M4nTu7t/6kqpBUavxdyTKOUV
CW3fImqTqLNx1FA8PXFIBMGne2Z4qcuPOnwDg5YiIBeSHJH4OoMGQE58Iz5+1iXgqiV9Fu9+n6X8
BUfVZcEp2RkrTUwrZaHXhi7M8N15GE1Lcso5E5o6UfXH3lunf0xPvDnmBi2kAKhAo/eQrGLt1xB6
+Oz+XXv6sQy/+dOKSXlnRRyT9mxx+U9H37pIRPAhD3Pk6p9pbCvX/+2WQ9BjqkrIz+Rcc++bYddJ
oF0L4jrL0dQoOQA4nq/wIuWJVgSvhkGW6i4iABawLC8gFUqxo+DYtmZhTbk10OeZWWm/28EBX6SK
qRNxwJnwzwl4mKR/4LVxYru8xvDplz4UPx2BELS0I3bK8Yefh4/8RipGRueQnO88M7glfmJddajP
0oP6QipWTr3EK5+wP5ADS8HW89ZYFTrBH+w8J6e2DcaD91rkKr86Fw5QHtfDARrN7coxBWDiMxMi
1civ0rlwf2XeWeUeok9J3V8RzXYZL9YRITYHNf33aYXjfWzDCnwMMw1UWtE5aZHm3k3c1Ux9ajev
nTqcCa3pDmYArh2Dkl1PkMz/WJocS6U+LP3JlO25h+6nWl4ndsRu52tA3YolTzOQKpbBa28UMQTj
DUSKioBFdZYidIvvFm0UDFBd2gCFekcAGyDARUI87B1ZHgyQ4KERhHbowaeyF7tPgtGszGQ5jzE1
U76AkVPwY7RJOXglqm9ufACxdf9UxCiNqubu6HC6iG2lOadYsFFpllFA783CehmsLUbUKL4XP5bm
nGObohIa98iPAaoVlhWMEEbm/Klugtww1fPzXqrFLwCLaWqvRgOleSWOv6fC+Rk5hTOy7W8SvyCu
T0k0Z71qdhXptT5v2ImLvtsN3JY4FU4q1gUHkcJE9SHAocf81Q312fTzG1gP69Ia8W87ddo3hWqx
uUVS9Qe26DkixSQDoSVK7fCXjaep7WcobY2meQcw6JZtgydplwDPJBoNYnuNvLYLILl9R63Ob12A
UrHz/7L3CeykwEW9o4PMxAj0MP9v6gL0rnBhd0ha6GpwoDQSPOJWaVGsalBKFic3+R3lXjpxMqEj
+y6G1/fKkO6uWdt1rwvxXqr+gLRS/5Yf3eXwprxAuJlSC2MZLzj1wQtP5b1EjOvPLQlSjToBgegW
DYlD/cN/BMvsYjUW59tU11uHyr6ElaY0m1SSgb2jV7HGlCoybGS6K61HEvzRcEZu2VZ4z6Yuep4Z
q2FPaygSzCyUlVcRlSsRST/ScR+CP8D+o8g05bNt6921ADR4Xab6aRTw0hmD2LNw0P3ZvztcOp0B
JlbElSfS7TtVcRzsjbxAKuBY4aMdzPdeVceCgowAu1MoBKqUwaad+5puji47B38pwnLzA7vopjX9
VtgQr95WE3Ij2Bh6ykIAjrXBDWxaS3RJsFS3lQZaeMQrIjHQ/KML2zSCLvEEZ0v/bdSkH4NYFEgH
8YhKgS5UowhdkKKPW7JSfal4KX7x1UQLPCy7AZLejXA9l7MRg5GzZaUmw9kU/yBJQB9HDbMxo8nS
KXRMG8TZTg2ijaXBL5e7rbeFentIJafuljaFH9aJcwF7lKllPiT5I+EiwskJYMJ9NgjuWkpa/sYg
AUZFgd+NahKKOEorsmKklmBhOmvWtcYz6gQD/EpUI2I506fSqEQo99O8ZmLxcJhESIQ3KknLs40l
Mcy60ImdiFUazitVp7wOb80PgxRdjvKeDpDkyf5gtdFBN6t9MwuStBDZwr/TWCSdqn44ko8TbDNB
62hgc9H4erXzbSuNMAK2LnnpNUwkQzHZQv5aU707MU+CvoBUZZ8Uj+OPehQod6YUpJS2if2GndQQ
2b6Aa8Kts5Q+4TPTlPT2ghME40ZQ4i+NCnBUIiT2to/T2R26lk91YaMCgn8EFCOM7DgT+o1a6rFg
2y16bBYSuJxSmP6uopIjVfa0PvHm20OJqwLsdW6SkhY66Vm4FOy2NITIuR6SocHKBMl/eQH5HL60
uJhGp5fX6+LZqNrFij4LqPFUDoWuLy8wpAvxeMs0nPmIjSPebaketM+YYeXjPi3ywCSy+WB2Dnxl
5XDxQFgy0h12vN2CP+IjKeN69eP4jIBJnu8RHjsfXWS58C2/tS/c7tpqysNR8UO2a5TrxkLgXXC7
qMIPFhXBKhv199wm0b7S0LwQ2fQ1g7Hq+A2IB5bMIag2nkHT1VPa0+PT520ehblBSHmtY9IwocqT
qEJtFzGZOkvwktLgD2NvNuSHPUSLUDdoeFFtq+lvyTQwMHxhgD8pOURlde80Ln6Y8xEvQOJULXfK
LOOd9BaNwCkdvuJmRhnofbnWCsOWbixOgewqGvzpqaVipl2trW14txsvm8zSelN7nwhHVpdA1AJc
INWPty4z7/Urgzo3Lj82sMeYheKyRmHya2msVCRE2pG62Jct2x1eSPjjId6R2ZftFSvMG4B4eGiS
mgtDNogZbmlX6KlTNCgCpZWP2DyfiHsresr5LSapG/0k501Nd5T5MUdzoSnBU459s4c/ZKzrOIiB
fI59H4x8h+dkgLocVjFpu6uU1p6MrA/Jx8DHCPR1sqrH2QgkWSu+t6okM8fHRcFrSSieP+KPsqhu
tbWt7oMEuq1GbCALm5Q/3R2mTRFlpt/f6UPTznqJ7hzOpAq3PaK0Mz3uJO8YKR9oRVcXesr8knHb
4oZSCoA4aOMx+CaalVsh+dkra4xPW58J1Qw+0G9eYQDg63+0LbSUsF+Eo7Y0UjKOzD/5NVh+RrtI
rQJb1ou6dvMZsKhQyAapJxhX8OzUJV4+dXL55fe9SRGuVNzNYuWZvgYUepVDrl+jk6h0IemQMP8T
ud88FraypUnSD+ApdCuBALG964esFewTVvjli0gbHl+iev/WUIHBviduZ42OCbjWW+ZsQOpjeKFx
HSd6Q20Fl9YtF+qzizPOFYh2CbhTHmWUYoWNj2+pdBvVtw05LWTppum6vbaZ/wjtycrdlcCkICM0
hWa6zQgD39itoMCA6jk3rqPtN4yWL2VPPT7Cru76SkQPWtwGufNYVOpQVfkNow+Ki024Wf0a6joV
bKNOjm8pxzZ1460h6w/ewyvsQKzG821Zz0yCFzunIIszbBv+BJLZ1/tFnDu+juNWxqY5h2YJ38Tx
BOaNkSnSVOODYySPXRNxxLAZ7SU/5WVJbBW3rC9s7nMbLzw/VRTOYFUVS+C4hN2sxiTIMdrTQ+OH
+n4Wzs5V1boPQjc4GOJsKWp4SlK4VpEC+k+hbGA6WhFcKvwrccW9wHQ767yePaZ3OvHMFQwie1q9
qtqdohmoHfvdM+vXpe6ZjIXgr/rDOiY702aRIKl5MbM5Df7t2JY3VW29zuBLYFtDju0lyZn2vXqM
tzREvX/3Gcgkzqytue7nPvcxgHXmWcVvXNQIMC7KqWCj2GIea/s9GWY+2wqYUf7m41ZtjimfI20g
Oq7hVu+Ib2UNgXRXvkMU3fUzgRWBfdIjraL+BHMmGD9G0aifPUTOvgLUPRzEOk1wEBGIvKbecAFw
6qYn/89rZefEeOM29YXWIh9kn4tBRhedIkPqtdffJHtrpN59ofg9KSIQPJ4pDX/WN/TU1w9k8nYl
6F3u0G7mcuksyPUutEQ58Zs+QWiOG6GUK770Dab7LMDFBmd4ZmePjQ7A3cAdFwW+fKxuPn4agqNM
OH7Wlh2qmIcQAmGEJ9iWW6fmLBACFqa5QRK8sYDpxIrfN9zEtym1EdRHT9PZkzdz7AK9LXZmqirL
xeqRZL143nPnjs4nWUHlKj3RRd5bPug3ujzQLzJWaIBiYYoct7sMN+yY+/kWiW9HK1pFKpVcbMAT
iCJDQoIGOdlVxqqrV6MAplAp+Q8BfSIX1INeEfEWbiTRxPFQiL+MWqd/lcSpFEeG5NsXPLmleCLS
XTYnOG1QIoA3vUz+wwVJUbnWhl5Wh93mP+jcisBctW2rL2ANuZhCLGmQH4NpzxbqcmB8gTbdTNR7
DwX2QB0dKWrsNi2Qx6+J10bp5/JBqOAeWAMxCoMNkF1+QDGV5OdWcONxLKw3u4J7mCvM7cpkIuls
LFez82tcD7o63hiDY5rhEga3IITLqoN7YJC8sPXvhbWgsORDm47Ehrp5gxkVg2KQAU6h9PG2cZAS
y3jDxRapasBswInnDzYsHcWk4z4rqEngKN0sXIa4KSn96JnLcwMcGDqyg3Lc9vDnpw5fnV5kLJXP
GHf4biLGE8y1NNPDMlNSWXljjs72ulIFu/byhFXvrFd603NSEA0ccgidXduDhUwER4oImknozZ00
FTY33ILcF0bvibMr41/H//nMFyXAAEjpCVNa47Xvvz7+KBSAXtMi6Pp6yK4YQz5yAr6HLJWVVr17
cEzBzCKkzkT8MO+VTkVyJ7i7p+g849MT1rSuMywv1o/+QbT4Co2LQqoZVVBTNKxMpKienkEe5J29
pq9CnGM2o/ujgFKJ/U5XCGE48QIoDrHZhHYOKQZC+km+73VkRW4gLEtlURGKua/2TsAi4yHzsrVE
krN6+dz5MXL2H0ZTcBLxyetLVHXjauIcbeBgjLW6Uwddj9F9V3RuAFNj2oQRtRcbI1ipDrZqM8oB
Vd0swLAXFV9j4hyVscndBmN5jnnYGWObeHZnFGYCPRci9kylnAFgsqNLZTsb2/wrLuZrDNKR8/LF
GNJFK67dB8nvAkwwCC9BWFfB49keAF2MfEDYZQsOnR4YUkgN72TGarhs64eTFNrhbJJ6ZHP+Cs1t
fI8ekkJMYkHmhg2eJzh54n+rwVio6Fjr8vNu8JzjbTf6WjPznoilEof0+5IsVZDKsBTa/58D2SAY
Et14E2eB0RD+NQsZlF+UQxJdXbVJscDc8xLeS51IspexnfJKol67OfqwYSI8wWAjCrpUKRv+k3T2
mrJnoFwXANN4aL3PH4Wme5AtzH1Jyqx1I3Ss4iTE3jH7sDUmXq/WtOkoXlXtn7Ejb/OE9UucXhy5
R+FWIN3MCevcZ62CYOxPYmNPHId6A+VDil5V/X+i/kYuRMiMM7IF3AgfIqG+AT15gJpIKeO4BNli
axEe//xEI3BDIormA7R902DysobAnsghzNJ8bXktPyXCxiWtStgOlxHzLkqGzAxIbbvfS5pUGfx0
HjpuZTBfAYXzX11KKaF3s+LibRVoPGm1EgfjK6nMBgFZcDsYcNf8/VxDLR2ZasuZxMj0HJLXMPs7
PdPGpNkUc+a/PIuNlDlHY1NTFrPXRIHxwqI0Lx93ew87LXxbqS+gSP9zA7M3PokI0anWlJllUOza
Emk61+++f6qO1NJ1HDFFPdgnI4vBiBbPGIsJ5MKh/f3I8Q7jr+D4HwfBgo64NCdRPA2GPxZ391mA
748Sakm7PHRZvV9B7jUXlrhQtX5IgojmuOAAQX+oIX7r6+T+0FyOOKsot8KW3hJUdb1TmLLMip3k
wu9DuNOVi1MJ34qHI/SJxwvAkQQfhczxNl0aJl7k2iZsOXwRy4ZYQVSvDkLA//8ZsS1vMBh7EDsN
x3bb0R4lUrkSja/49crXYqCuaVUYqvC/ctG8METVr84HBmzMSHskp4pw+OQPUGR0ZABARQjjKRDW
ylyRb+JycnToUHVOXXxpUSPtow+00MkEtPVuAYIt2uXbQavkqas35wu7EDy92146X2MRF7IOATGe
vOl+eaNP5LGZZcLtgNXcK/v2+KotVQU37d45eyju8E/VbHKvlDb0WWfut7NdbIM/u/NnKbPNGKfQ
6eidRv6yZfDafOOdffNBYG29bgyzSMeJtuG0gl8//zj4lMhxkFXrSetIJ20defy8gpLU+08ZfSr2
Ips6DWNH/J72F6ChkF+YsLtWBbxEqS/nBiq00DYAFZ/ttc3HG+b4+aii5eGpMJttuXA/P93d/kHs
asUI9FlSWEc8kWZLEqsQnwwBJCQw3/Bx47oBIAN1lPEZMH0hLXG2l7+wgcMc7qgqE5cl5s4w9Rk4
IJFk+P3jUKBRTpw3aFANi6of8pqpO915anLM/N6K4CSGsyOJtXAgIltPwNd0k8Nu050OXNFuDekA
RlJHOuJ2Ou8PZ0fss+Rt/LPRktQ+cOu2/7z2GCpB2hwYAXIWLu8io9QJVUoACQUxEMH4SeNRr9WH
W0jF+fIkUx0jCPlXYESGWC3BXrxQP3KzKU9J5oOzBhkpm4Pyc47DuLcHuoYNJChxGh4nOeFmn57N
jk8qYtNDVtQiMbUEy0W8wDnbFHd1/RRJg94m7fJlLvLygbnK0XstrUeE5toPfdtdnFU6xwG+/mKl
mn+8Zb93xNJ0fda75TobLSQGmJqtVj0aBTVKspVvvW/WVqDCDk7uLeSuQGahtxPJ51aG1NlcSefW
Wm9G1IytEwEQhSY6Nz+PM7FlhXrS8ms1mHXbcukGDCwfBX4asRklDp28M3qNPzE/BDt/S5wxifbb
ki+VmyGiX5lY0WPqbqph+TjEBKEZUQtIz8AbTyGRKqRUKocOVU70gW2wBvXHd3fh4njtmm0E4iy7
/IGne0zn6YhRjVpKBer7DyuyA7JEu5vjbIxL3ZS5CJeiEuc7lsRLDwVAB7bng2e1RwN1ZJx6TfWr
LJKhImkZE6w4xtRpEOEMvHJiKtl3d+k8SGr46e4VviRYy7B9WkOuU7jiM4Cbwzj4cIkO5DSjpl3b
nbWHSkBCHwrIfRUUxwYpoHOo8tLWsBsOiaNb38Ql3Cg1wcu0AxVhBv6zoVlUOZfKAm3JSD07P9GD
pZsXrNwuvhWcMATKXYjJgz/Te3weqxyxjTT2kj15HqaxB5dsTPB4ofJSXxY2iFLStsHMBAfITUJb
8kcgvsEM/FdvI/AuQIHSm2TUPGFHnw4BmntJqQE5rFKQRsxijyVusf38jOps5VsLDgEb+aqJErG3
QuMAFiL8Eb2iwtcActd6vYCuxQrvbH1sBxUOkNYCIk4Q/VQd4ucq5w7QLyLsIt4adZC7UkoweDdH
nBMyat382gpgxwqPrgNPy+BqtFvcrwLIUbvrJQGCjp+Pu0TIK9kt0ufcTo7N7Pih9s4FkTOla5Q/
kCeZJwie6m0jQq5CGD7kVW5cJH+Ltc6u345KuKj3gE35TEtRUHuv4Fqsn7ntxU0LalcSDMlATXPk
BiSCKwPhLgEUxNEJvtnD3FV/1EuxjvacdYsNjRu7DX8cwVaHaq2NuzSC1/QWI4eU0EkpB7J6MOkk
6f28l6VW5AYd4VVnxrvJFUshVo8k4YXRqO7EdWALxRO8rAEd9FkbeCAi2eAply9qkkoalY+G9Kv7
3TCM5gvL+xsYOSyr6oR3KwJnfETbVPguPSopH5OdCWhB+GCXW5qenaIu1DAkY/bafLKRjqdG9Pka
X6w2inSbUTyPgT1+KCx6Twnp38vLY3kujQxn5ytmLKcn6qyZYDXaPNHLlqLxOdcIFLJF/dsuq4ZT
/zSG6h3zTT+F2FWKrz59Qt4O86gBrt8PM8jEDcjvIjN2uJurpViy/E75LH1VGwD0JywZ89AzwIis
DMLtJLkHaM/uIQPsQTRQMQu79qunyNPB1TVH1+91L2VXbBStrHkNDYqCNH4RCy168MIt1n4fqz7u
B5ytsNycWkFakN8pKZme+1FDoOwKmMkknAKkP2qLhT1yLnynxBIURKST6tgbZ5ae/yHqsuegYR++
/tW9qMadOAtFdXEEIFE1m3U6eC9YHVpwYvrQPHKv4Ys/o46LhgWt+ZWK4vLIrtsKOpaXgUhGvFwQ
hYVyy3jdIKVu7QtClL8sSgvrwyEjib8VnxKCsdvav9y715GTfHDZDmRtr71SVm0EQ29zlbUtF0Y2
GVPwjBOTRan42vJhScisOUFw82okNehrKlBawk6MY9ucW3n4ExIgPMgCEt9pAepIinj8VPUESgQa
nQ3SnE4UgdV7xoVz1nVBl5SqSuD9xaBnVn5to2pW+AgDFHSXVHZFbjwy0ApIIE3MW3/ja6gqAl6X
6mmI+B2+SUHTptnGSscmbA2MvetLy/CeOj+zzixjwyonqEU7dB9CP49WHKjAWyxJBmeyS/5tER98
gweoHHA563beTfaiAbUYgweHjYKkCltI9EbRpSalsogfeKkDOQtTcPe48ldQwWbHDn19qBtwBRAe
3IeeI5y6VR0fxC/wht8Q73e4ER/DKSp5AX19xqMr2vt8gGpsaR0loL7+UyQgkoeJdeIbFJZnZPPU
7DbwSJ8JcFf22XUGuvfbNDGx0PeoEdDV+w4G3q5etEGj+mmzAOrUH/1XbZ5eyy8wPIlyljtNkTBf
lt3GijXRfJUHGPfao8aBI0voAmsfwwtF3npGUnUofNr1yxn6CKIre5S9jXqTQ6oH0hNOGEx+VH8R
xYpxqUmWCrLMyU+xC01ZR9WsskX+V0d/ktBl3yFHJp62+Ga9pZYSWDNbXzZTegonE2O7Cqs/OLY+
zuaMuPWPgl1Cb2N62tSM+sR0+DSCGN4lB6uxtAVPIuVrNuP23jZRsECaLrcHOB0D6IuUR8n7jlIM
vM9Ez2fGG/M2p73kIWShJCLjTuqTv5lBnHIJk0Klp5vq7kAnxWxm3paTfvrR4nE1PSyf21XaFP+B
kUo0bHjnxtPDT8qPr0C5PPuMvy4nMSOO50u6RdjdyiMnla87d23/FuFgyf/1ThTQqA0z/zxTxWFB
KNeP6wlV9mfIST1p+pqqbnQI1SoCFo9bNG5FJQHbN11aeLs/CGvzfZHA8OMgzwb2OKLoDvyiTsNJ
YE2nHaDutJci6eNYUZX1vzLznD7iWF9fqHNCYHhi5GmUSKEfC2SdKh76aAP0kH/YOzcBPbNQxQJd
lqbbxnyRc1Hq52wMt8l1f8J2psToQsOVp+hZRnHK4P+llA==
`protect end_protected
