`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
PdDUJE3SVsklNnDBzX8gn2evUOzyfnvGs/jt/psKtDYet70e0lJUhAOuAxevuHm1FVSynSHuXk1u
oDloSqhY+AhvKG4wg5eMzfbehpggQVX5EnPm2u1Z3Eg4kaGpWb9fpL8Emx8mKq16vEWts7ciNRu5
feIAE630DaMo/d0sczipAatW3BMoBTTSkwSiSzz9q2X1G4TQevqYORf4sEKkShe5HQvajEFQTp0R
q1ZeLDZNyNl3NCRXbBwYGQvW89BJ8+SXtBo8jqo1YyABW/L4fDKvFK0hnLSBmb6iP1nW8KOMTuhS
gWjNlsLXcAAqsh3tMSMp/3+hHmsYruYCfMbmvQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="EDmeAmesH9PZ4msFHblUaWmtuCnQSIo/XHHwQpYUeZI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11056)
`protect data_block
3dAHeKHRV9/7zazofUcgcE6LJS0Lfos0GEx2tq4mNrG18mZMw/PpbKye0Sb+4CsgCdNFtxS/7ctA
HXq7T63MGutt7qzJsdfWAshDKYuxojM3GJ7UXt8T/6VcbzRJTerPK3V8anSKwxRJ6Lw/yAJhWChB
otoDUxK0ppCaDep6myi92+YdVgvdrM5L3zX4wcjKEe2r+cUOpAlPi+kClTyF7exl6/L5P4Rg4dw/
4vnoApSo7JSL+Nz+XlYNqNyNMcHjivWnu6RPZLasDbY7vLh/FVuZSr3QFJJVoZHs7j8+7urCCR20
eDIWiBR/KSpexE2+Z8q0qzlWkGPw8cb20oiHwncCPB83t+qSafoAGCfMuTCAfIv17ifGw8Ocz7fg
MjvkaKtZIPTAMUqeMeyTZuQihobbUdKhM+GxNzAN66YrdeIm8pNt5HxLh4on0BzaNKtpo5/wasL/
eSrdGTiVjuZvQp+VGUwkMDPc7CZ3hLOQZL72wVYm2lm6qPob25G85jPV0ila9YxRh77EVl8M6NAG
GqLKizoQE1VhZEKI5g5LTtIbxrJCb8h9AyZS/YPOSWf3C9hhPOxrfMehcYW9g7TJkuM+SfMZbT1G
hl7KQyKs8/MgoIZrSxaYYPkkKRDqDe0V78hcJMo1dh4eVKz5sdcQ6xe/sIwrATVzCe7UVZ+Z8qku
l1mgBfyMS4fTM+F9Pz2pI9Obm9D95GgExznddgRb43oUtu2nN3czmQeOi+KotIFnOjmNLdhklK3+
QkcB0p6ldWsX8xYkgU6WHa2OBJ4PvgdnOFsh6F0BvDTvM+HprwZVw7Qx5VbkgjRl5EXAXjqcQWyB
jgDSNTbujz3FSkRyIa9YRvdB4EGh2eEX8MHer1MLlVmTpAcurlOvMQrboeQUhpT6dGSNcg8n0T/q
0vG+L7Q4xU6YNhVjr+nAx2pKg/DJnYvmC9hvCVpPMmbvnTHbrezNGe7qeYAzIH5C5UUX05wLLo1j
XMhNepDJeT7kC6zumwjDR5vOzlX3vPn/5Frr1NMcxXvVkrVLViAdB5loOZ1BLMsCQ6sIPXEtk4K2
Rwcrb3NGC8acve050DG431/FoIUgNLV0KGlyZyjNvNJ/o2zAHXoYRBAXF+VT7fj8wn84q+8tEKJB
XjnqewQFrS5Of8pB10I+NMCj5TNHkqprTZhAwUTQfXdnnrTIMOP1WTRwhmwNSBYmPMgw5Wio3kif
oAmx9xh2xC3TbEy5gdiNeJFXvwJOjqEzhcG8Yc/3pPQsecYNnBOUGR4G7y/vgGFp3vZRp9+VPDQI
afIfUmEQBU+Z9/uIqqOpRJkuIMKY9Cc9F96Q+Sq0Gat4SwNzn5T3fDAI6j5PEkLNYHxSxtEMXMiD
aUq8U5CrkxV3DEnlEeg/jXlsJMfFntbpk7vI2i1ZbSdwfEqkkuXRpRtryxPISNzdNbIfnNmH5a85
VIlAY1e/NBQY+kBOsHZNh9MCuXFFCi98Fg3ig5icwtBjieKRLlHsffinuc0mqYcrUqPm7STGZQbD
yqhh3Cwdnw1lB4q0Mfh4s4j2vYdMt7kMdcVpideSJtR8J2ae+qYgAK4Dv70vMAyU8IeL4PRipPT4
H2aVftychoFIRv1anwb0RGfpOWX7HT1fNKkQSPqoZEPMMIab4mZxdHvAGetV0vMZp04h81n8Tyys
Oq3YhBv7oREdFspi/G9UWZm8xJ/4JgkonKNfSQsJzD0Mspgsl7b/cu4buKAp/JjO4eKuLTOE8cWq
aWSfoBcnLaEugibAGHMOqPyghai6ye9Z57844wGYBoSaJ+sfTd8PXJW0JgaUzsBPWXv6io0xr0J8
l1+7ggaq+X+Rkz0YGfushuM4stsGf+0EnfneX5Q+fWDR9GEhqmK/j7LzCoiZxxqMbB/eeo1UdJfn
2PHmhHVfT0xIdNigNFha0/szlRxud6YjIZp+Zf+agu12gabjc9O5UTOXSD86mjOPgE6sqfAaW41e
/ab76NfnDEo2o0aXYFJQdu3yFEGXdFvQBqQRB2vWs5WL+R+EgsvW7Gd2y9Q4MYyWGmZIjBqpky0h
4tlkUU684vQgLWtPYpCzm3jg1o6DtquNGtdVnpcFUgiKVOTLP8slkyDcA39EDeredG1Hf5LvKLjI
PCHPwDmwwoZLx5q68gO/0umk4mwpFD0NsZTI2lRrcS1Ayt0RyRXT7Tr1n0KKXr63jW2IoJqT0KhE
Vkvvm+GHS+FR5YpSXjOrLzJuthJJE7Ok7PjQiKh2ETsBm1vMsqub3iHRUNueDe5gUbz0wbCQ5MRz
jTuweIihVL0K8V2axAFX1GLrdK5LMNLe5VvceZbxzmsBlEi26fqpxZOKa3MNKwEjA5KQmztu3hdK
8DReGuQL59amZEysz5xxzlZkDVMbzm5qcA1LQAN4452MHZwa4X2lA2q5WDbCHDVlrmtkwojS+wpz
7WfUuzbOoA9IerB/afbUhr8UquUBI+XKmh2k1TpxP6+QQ9E94E53MkFy/7Tm6QEKKI58pjsAozVx
p6SrLtTBeQRDobV7LMGJ+zzCkk2ove8tagpVAPmhtF9hnseecYQZjm+6VL361R4CkRt/gpKgHMNJ
Bfkyl8Z1LFm3h2U4txjI5WEK1ypsG9vzaDSiQmYyVRpwt/n6NuHYdnkpXOAJ6hwz40w5htxAwurq
W0XduaU5fLXpeVYxEVGfCCzK+c1i11hUU/eeNCZYAUy+PtC2gdZ8aVn7HRE2nPkic7yfdP2Ddtxe
qQaZwsvkfRTgyjHdyxUxkt713FYn//XecFeTZOzFDtG5TgoLdZA/zmhMgmmxqSu/CQetPfaMHt+p
cMjWCWpIPdqAX/x5SbZeH4YWp1uWjvUIDGGPZol65TAFMbtXY5dRl/QLavqsQ2KWERnKemsFvmDh
SBd+MspttaJ69qLCeNHuROVAn2U4oDH8iKItQgUytszUhWN3jDIZF2CfbWx5RDf78EESVsdZWzG4
A+Jjpv7ge08WZFSIKp4i0Kg64ja19ubf+v2qGjSfEPMXN0mO6ll5+r3zFSndspOXwMIG3urjmZTs
xEAtRP5Oa8AOO2gpsutVhWaIE9dBWpl2iLusRzToN5jKbpz7/2Fyes2+lzeVaobho+ev+hspiHCz
om+/yax9qVUmERZibRgw+FRSNQj36PG5VObea/8nnZIKbt6h7k6EsVx6Qplo7RoDXCzHMrROytCX
xn+aP9F1fNtIkSYdlHkEm3X5LdKXvGXbFRyCHx8LplBCPPerf45jG8PvHWx2rOCe3zyUJPSxHBu+
LehJSxeAKmwGanS0DmBntb47owxg5Be8wvI6Prf2m0hT4D8pqGtvVxDPrtYu80hKzMze0BJkeqZv
A6o1hzn3PLYK9kGb+4nExpqt3l/aXiBEAi23X8AxgxYQXICzu2bAJOpr96SPzY1L6a1xpyzP7sa1
U5qoqAuNg/qmPEKm3WtFY3rEWbiQ5EPRl8No7coQLZJq1bcL1zW9YLnJhvZ1X2Rjw5V6e/4uxLEG
EI5NRHR+3Rt9Siv11jR34FaKAKbflYRz4H+8VdaQwEyw7mZSY4WYrj8+UUAn0TliyGx2mKY/Z7Xq
nWPARWGgBbmD76iP3zWnfTxsqc4Pr4vUdHg/KqD7FMeKdISveGgd/GohtxhXyznDXf3Pk66nC/ku
akdyF4Zro8bakf2QnLMrRqnYPHWlkfMhffrNap+OiXdaliB6nSxBz3HWV6pF4wBH+L0cA+rcuSPH
WnanpecRLnUtWyHdsOqNCml6sCj9k94kqMIlc1RD1yB+6TBvlvr27SZAmk8z1uLINnSgjrtqc9Yx
X2DgxnU9j2Ix4LNBxPuYoeqQyGA2XrKtkwS/cXR/SuGbYzrzae+BRuCzFn4QPIAeyq+yQMGPucdt
58E2gOP4nAX73rfttUddG1T/Lee4xKQGiitNhnFjkoNOLG0V+nuBLwKk1mSbMvn91823rR0fK1wm
8FTRblo4FllUvaEFWe5+ZAfZp4gHDAgs0jbrF7GE0AAsRdZOn71t+a23T16nzQGacAT8W0Six2pF
5TWHlVR4sdcdBsrV8hWKnRtwkBrkptw+aipZAD1PM9u2XydYANrHeSE5pe39HQR6Br+lsEW00gpE
a1+NmdU3KHK/TILyTRV7vp0kB/50wpzrN1oRlfz6lO3n7/UHcBk+wR6LR3up6EXMr9PV3/VT1KsN
/u0Am5aP08dbDE4CCDN8SP4UpPY6/BmVALDkTZLBJuMg5AnuDv5WX1FI8FjRHZvqV3D/Eomz6jYx
1YZVtOtmNb7tPFIvfTpI8bAMyRTN+2SpYT0bsiWL7esAGUX0oSMriKPf3oNIjb2LmIepJVty2u+A
kxVUnCuPVPx2JqYUqseuEVUWyrwuRwftkY89jHPWNkzq8sOp2k892Q6cY8Kzn9x1yOfKcyB6hXwX
3cUcYxotSibu+CQEoUrxSEWz3bGZEmpa/EKgLo++8GJHkfefeHSES5o5IgWihzBrS0rI8+HXQXTX
1odJDD6rd6LHDSmmRsy/wkmqdIBEmxDKeDV5NuRjqIWrW5EGif7HkCi3bzcxeVdTWREHYu2cAwHl
k58Ru32KwpI6W8kiHejn5NQINSAnWQl0Ane6ifVcsLmSZCK0p7FjzkBLUsMox8wA2re0r8omf+gU
saYpOXF0HJJzHJtleGwReuyDK8Vv+FYOzVPhuLEbuSGro/ZeBQl0MeyKTfTQVlRpuCYxlDY8OrS4
Q33H3gIxPBZqTKJA5HRhamEfbN5Mm4qjZQEnjkGzV2Q+EEaGe1z+r0BFIU+2PsoNM7j0ylMPKg2t
e5kkXOQaVnrSThkt6ZqBsjIRxFH2iSY4sjYLNxze1FVsL0Et7VElMHgc08v5yT33/XaORsmmnQ/8
dceBYB07MSejAXA1sj9X2Y17xYdLFlMzTFx4HIKV4AaLSj3TvKwrbPFj8qmmgfvZ1E9127fUVGYF
A2Vxo/b4tqrDFL5VZctOHAi2B2F4rgYtkkgDKlfuOgnMLEP++sisI/JLUIMsv6V1297K9t263zQ3
fZA2DutRiyWtIetilGY4pPSHy589N2BwQz+y6fREqs2ZYsWM+KvzqG8Aw1HPdi7KBn0mm6QO4Qyl
l0tXCq8ThvufyDcGSRtihAwTrvp0rbBix3aYC0WxCLvvlCCbpJ9Ow573s5iEPXikCC+URwtnuIYs
iazcoDt/YjUWuYmjV1HNaJXNi1NGHgHRUaScDU3B2PTCDSTTGl1iGsFyx5KCnD/LxCuljVRH0/mm
Pp08d5/Cq4/YQOKns2+XjlMEC485KjarpyMmwWBP/VGj6nhYGBu5NoJT59PqwldVlf9YHh3BfvCj
CMRI8gzPLlkOiC7/YjdExbfpDn+X7wHYkG+ZL0hphla9cYYYfCr53UJxbdY/EdrKfmxxUrvXEXpU
PkNu1jOrE+YUInvzR3YOu+6G+RnJBqYhSQWc1TRHFoDDU+yLLWxX3qJih86+1cJ3En4sLydhOxWM
mi/a19blBO3qmgopof2wQ53P11C748L8DWgmPzp62uC6s6kLLA0D8Obn3EZZUUfFPLuPkWlIGN4d
qbQmD7MmnshECgSVOiNpTEK805/0E39dZZ0sRsPdtUaZt0fvI4wt5m/owA77egEJru64U2WbPlOk
0nUIesxudiJAM/Ibb/SPxQA1mKVXZ3cJxf/ooNQR3HbfbwF/9H7hLT1fSTRlN72H80NTgrrPqE+m
aBEraKtBuXd6loHnoZk0yHD60Pgk7H9OOvHGRF8oRB+OEo2eR4dfoFetiuFPdFBKRCL3KwaNsMO2
BiKRxMVUqQbXJ8ji/FYQvVllBWj7/TalD5kY5WtiarZqq/3Vm8rc/+KKOfghMivpfw25Q+6R06WE
MLa4bI2c7lM122NNYBRHmxlk7CEfPm2Z/gqR8ixn7EhqqMIe7SGIc7XoakvTgR4XgWzvY8TuiHHs
p0l2AJgse7Ur5mjjoUBo0Pi9dCYXty9iDQGEtMpJRS+rqHpSD7nSJp59AY4wfH6Y6IEpEzjATu6E
Rt480fKJJjEvtPdG272fgxoZn730ZF0P1XfMwXiCAi+PYY5h3mb0MlyayEeqtTj/WT22+ZFURaFT
nkB7sjoiuZ7sxwGtdzIFqLOT1/6OF4EWchs7iWhJ+CYCLVwmH/oK8Rkz7Z7xaBQS+vSo2yeyB04N
I2zwauffZR0wu/Q0nnw5paasmdv/jV4ccAKEPq/ff0y7AamPH0gPJLrroUIlEna2DF05reK46L7g
wCJgyqRQg/dBGGYYiZCYX+++a3Q7KgylCZiXGXtWE2KyQBlPYwzjLsUiHM4dXy5mQA6ufDL2rbnx
K20OZVGOmwyV6qwgFcm0dc2n8odhkmfs3cBHJUJgSNleuNlqxjOSGf0v2/j9DrZSt9RlgLSgu7NF
JYZSut56IC8hqe+ocH00/v8qE/SGmNpYyaZWc66fBboc4chYvM6oBUuT8+jd2MVP4JGnvgC3HQhh
8X8M9HinG5sVrk9xii0KCzWPkuLQnFUlqrkxPRRdBrKHK4QhMUriFy+2QSYvJYPGiRJ8hfrb7C1z
scU+vNe5a6GDWNHHFLchqRqxSmBfFIgf+1X1ATKs00zY3+GjqUDDPuUd0QMD9TLb7JLHgvdFHB95
OYzJfrNCb/hkc0+0asWd2s+7BjEQ4IqlOU5KWVUW0gpn22kH+8Xdmbsm3ex8GHsjDhvHGtl5tBiQ
PrwEi7BpnbxCSBvgvuZSgVj9EtBJdxV9Hh5fbI1bU5LdplGy4+VCswew5UcAMD1SWPzVgpKQQ5AK
ps2f66nusKaGlz6mPZucJSA3Vl/k8UuuNArVhv2M20+NM1+O9nc1jKGVMkVam8vuCPi1oy6DumM/
MsJU3FQjEtsD2NFO4/k5Q+P0NRFV6kF2hgiCGFD6U2wSqduuS8LJHtAhsqiITmeDdTXwgGScvKEH
36I793CBR+FpdfrkuBHkoyg5KMhaYRVgnkPSok8Q3ClerpgdWj1PPPgLbGUsNQBuXObaG2lfPnp7
UgemmThpzmGH0chV3c40Lm0+o+PYLKu54l/DltawQpesFy8WEHY2pRX7T8hi6vKrA1E/rRYPOnkv
SBlG8p3wL7EMKqa+PDWFKNePxSOwV+kKEeAPToC/Qq5qJ6LtE2oLcSOuIw1pmzonwcvSHMgj8D9T
JiJ19+NCFMUk6f5rNAtXITtG+wcz0LLy4prvN15M0BHNOuAjhCZiLV6OZ4pG1yBcbcWJ6op86Miw
4Ie8mTVgFQCOEoeeAg6TwkgdWNeVqaL0VrVdlGU1E7wKZRRoDxe2jhYuxROtbPW5Q5nC5Mb482hD
zX1DO6o6WGvN1BZnLxP3fiejFQodxrWXK7VGtdLQPtyIzsGj85YnCupi9ssic6WQUa42XvSJJV7r
OiAGQ8+povrYSsokUuhnZ9ISzrLVJl7BEOxiyNNYqOH4rDJ6Cf2rrReyUl+VCGmHzy08WCOQGaMt
yUIKFhV7M6VumlNktPixbq+mWLOTset981+fzfTLmTkHlMGUyUHn1OvM6Egcvkk3Lnb3ziLATDXc
b6SI0qf9Br50pUJuMy/B7uAtIEBsKJDrNIivxfDWTgnXXDnkleDSuqwg7LBpGVAOiiXO8eKwafZ7
5VEC0NLwF9bARTBwSui7CN3j/SnXjGBe8uxMffjXVTjzekUTBdTnq43YMeKlj4plCwsSaNdc4nNK
uvgmCJoDM28R5DEXu2KlrrFXZv9n9TExiBQ0gVpRThVo1LHRjI/dP4xnyfZESTFOUltvswXsYR8G
ugL8uqVwoY38pdr8kLuFygplw26eZPf43Y6iS0CO2vP26BreZKuUYidVhROi7WH/M3t98Rku6A+t
PAsiRyM1QWWvyl5qq0xzpOlokLSNcTONOw2b7hAuM76k4l7gvFJ42+ALLj0uutYEf4NrKUpEttu4
Ekgr8Dspb2ZjE62rsV8luipj4qdv6nmWvPPuGhQmbYQIQkOAu9PMbvsSde2DlTk5/u2Sn1LsAXf3
vUatUjr1Gz3br9mb7FMqtASZNMGAjkbg3BTdu36Ay0h5QTz7mDeCjyVQrCMZ1IUQBEI0SNJN+Q4G
hO78FVRgxe3ZuUNJma/7odcHSvuNDhpGRmjiIfwT/bv2COps7sra1x19jwSJPaHEezU/9isZ3EJM
oxbUuX6HF8CH4HsJ4P86OV3vovmXuBRu0vZJTCtYpGUCtVwyseSAqRQ/Ds8GgdVbq96Ki6pjMvnA
nDRs6LmGsaDdG4z8e7Jbkp1LZMJpWITRm2jM/FTHIvvQI6EC6FeDEYceb9AxMtrYAD0Urzbysqsz
H1kI2O/5GgcEBaVtejTnyhXAi/NMAWsXz68sage9f1WyVr/Osh9dlTLFSQwzc+RsxWVraBAz4X1q
iyIQ0KueZVU1GKrUqPQ3Qmy8ngB/B6zFLYO3YPLiVmv5v4fIgyLu60o+E7AtDQgdPfNveotM6rc3
srU+Uk3gPwt+1kbQkrkFDB11p1buY7SCnG4/W2Z/tBC3gPFexGycge1loZWgwtnTSt2Ik5aaArFL
Kqj/xevpitjf+Mk9jW+4zrUxpmgv3aVopo+illlKGUxPhmjUzmZF83KpYf4AmTdAOWuwYS8RFlmu
lCCUJiB5vWgkztYCLo/EcH+jBVnXpc2BQnLrTJAtfGtdXhLY43E/Qd6cuFskW3OO3aPfGfZ9mZia
FnPpkgKKLZCraoADMnzVLvUCul6U8UTcuLXJw+rmdzMMU8qN3KdLpQUnL+m4zMESTDQqS5ycp8uA
7zjuZq5NKHrrh5qfstB9cX1l4otSQFB7nl5pVXlOguZFSnPdJgCv/nONiwipIkO7BY1C+LWISTbs
wC7ccrAVq0eDIY6TvomUqTicYAWufcMy/LlsNwb8nGsZeaEe34BakY2t4aDrdyh9XX+WZyPvFqEC
2foXUHEDiqS4eTs8/DjLw1++aeU7L7DWCo1dLI1NyEBByzLTCddPM5c4ubCjl7kjEEX9yzjx6AV+
6y59+3k2OQabldJuUDK/TT0fOX43KnzMYeozuO5rNV7oSGHiWIF8d66BImbXVDG4fER4u+YdFE+v
FYI4On76Lykp9IEqxi1z/XllepUH9jr78So9Fufh+Zgr9IfpltlBfLAdEqyXdgM19H2qstKccdEJ
tEpG3pUGhN4QG+GEWd7cMd1Fsuc7vZ3FsF6rYhWAPxhGzxarFVIkSpmSyzVzdAy2EaMp2ODN/m6D
caq7fZ2znEtd9jdVc4tOV0qhGbGU2+B2Y8KCwBxjdEUt0NjHAB6QHE0WUvJxP6yRewoOW23KOtvA
3c2eKdNHl1BSDaeEhh5WmzqHEfnrDPR0W7MhJz8Vp0X3rhvRPo4oQD6TjJ8E9oEagvf2VxUs70Wc
57Z+lXWD47vnLhKoDph/rmWJ3GhuRKSUUYZdq3wrp3rDy7cIIt8mdcHvW8maKG1RacLEkSyB2jQC
OZKyapETrKjLHwm31cyScpQr7Mvd8rcaWLq0cfgmUE4IWjaecWwXELAaTf0VzXJJb4gyhX21Z0Pk
ouE90M5cbwAmuWMs94CpY3mgRq3+m+SL8K4LxJxXno3AUTxlVGzCe/dw2vzqHbgIDyfn3GGmjhIs
N5hR4l9PtVmTzjx4cs1vUpu8pl+CPmNA+XOGdhDSR8HezJLRxykbELP3W4Lz0meyZdiocAK/biGl
/p9ySOasgG5r/2ogvYXqiMZhHqxvoLQY6kdC/EpItlBaSWOAYz8V5I/huXJ9J2Dv7YMLHOHs8TzD
OcQMX1bjvsLcWC6ySgYgM1LvwS7+fQLy3HEAotD87GcLkG/FnfG9nU2jd1bX8OA7n0uG0nKp/lqE
r4DHBqpRRwvmBaGwycYITt/l30iefeMr3JsBH5oFIjVK43Py4Fw5G0ao70XVwAIjoTXHY6+RILG0
ubbtW1RBrazkMKzeGS57vaHEEagw1crqEGWM3oSFui+EJNPTmC9iE4d59i+c9jx1PJL992seHxee
i3AEcxHMHTZ9DY4JlAlRMDwjpxN296KokGY9uggLSlo1znljx+xTB/lOwxqkq23eama5lLuiYLAh
9t+XZmNg0cMzIdvfaBH6hIsmlVXWtkK8MUQov/bJMjuzI8T917GpBbq3q7muwqscDM2CJe1KEK0L
p9VeoHR4LdURABM4LYrWW1wBXosvKdj6B5QrQWEdT5E9rDLDna059YsuBH/fUFusA3hS43hm8ojG
ZmCIQLz5q+VC1Fcqx1blQz6/IQ2OD4MyDXzDd/vq9OfYVrixGqUWnS2TDxNNzHA8yFRupriCm8ii
m8LtYX81OHVfC9WyXnYFkjqK8IDUYdNvEiD+czXMwxlQV2Q8OB9Vng/n4o8fIdjrTiNYlPpQiMqI
ppYNQwK7lRCj5ibnxo+LXL04c2GjmGIgNrShHZbqqPGGBZqFgtk9s7yJfW8dnrvm7jAZ4J/4leA3
XgJmhoWKtj2gPquveOPOJBZePzE55AQzaf1tYu3eo6UpVhSs8paLIG7+tyCOuO0pB6N8RF2w0Y46
/DdjIYa5DVqBY5p2Ljtem/GOsSFJdjXA+iMjiU+nGrLyJ8tXCHAWjyB31ICRazwUjQaZty8xODZx
Bii3JzYlV4sxBAHgW5oiSQlbBXvLJzGKOe9CsB1Ipxubjk48+MdLeOIIDP1HdjlUc10jTEXttGBz
2SQuZyK/8PjKyCHCuGoNpeJtEhsWTWrnhCfdRzEO5f+JPKXYPwT/TSHBqyJBrmYsfugUA4WFwvjG
HmJyN/aB2fygvTpUpJYTvV2Xe9cayVzwc7D2VaHFkPjQduMSfOLG85nbo1CYuWDG1GKuyU4QcuVJ
/PhuXcBdTPL/Q0u4kME5W93QniEg6mTfz5sEQRRmRTwvDlbzYbXSQ0U/RfFftpUKgvQG7rnyrxgF
GyQjV5XBQv2d/t3v73aTqPDzCY+MngF1elwjJV8GWrDtj8jr07aL2as1OgNLkrba1O0WmEzW9l/T
MOUcp2qJO+8d/wr8oMp/mTm38dOt5OYmlYYpB1sBoHtH6SxuSCJqWCM0h1fh5LDnHBIARqKr0wZ+
aZbov6AuNssd0aHkH+0f82XrDxH0IveNI/ltvNYVDRS7knq9/Nf29V8ZusPsoxRL165dqpA7SuAv
+nV05a/HM9G2Hfk1T2szMOiCxVpI5OQlc8g82X44M9RiCKef6xewccuLdrIgPIQmS94B8eqpMGX1
6aeJqaj57uK448V9qQIhKGrg76iXNgb9O6Ta9anh/WkYaXH0EMyvaxJoIwTLfkZQ8OgHBqHugjxG
xsABH88QdgLeY9I4yjwxB6Cx9MYi01DAv6IYkeqqQzQb5Lxy5sIK9vjpDbFBbmXXdTzgm2+Oppoa
B8W5DVwQG9p4OLUEHOAsxBFLYMFcl5OVYuN53zGNjHmP2qUoh72aRg/nGvRGQs0QL7XGMAoX6hca
xmSxh2P8FDir9EHpXO05cGz9ZaRGq+bVenx8WrVoFfq1o7Nm3L40l3HmBpIof6oZpGIZA3Ig7o5G
gNB+0KD3dhqTrEIBBUjZ0osC5Sp0PVfalwIBegXUcSP3quHKvf7EaqW2VAb3nVBuifsnDIv6x3lI
AWZRmv7X0tzLwV4+XWDKjI1FCFMzcX7UETkb5pMzVChUzSQdgIVmK8sqUJZtuLw62TsNtBXelIA0
E7NF61W90TNLXqy3eeMBESgDyN1WyEI0zHIc2ivDd4CvQRKMAc+W+vLVtMZvFRyVhHiaXaU1pZRV
wjykv2VP8EA4HBmK/3mRAUClBAo3cEm4x4w6iZjYRi0xWnryjmT1xwS+GRQFMuGaqT7g+doEISqv
1RdW67kjl8EZ1a+VQdcqup0t/+f5keiaqxtOAeLP54HYNjHNqIJeE1/EeoYFCMfb6EQmvavRygms
2vSypTxgHLJAApsiUzn8FSkYPEBUFQFKs1Ec0B5JovQsjsn/h5/n7VvlKqeHavdBI7MyrghCZ+hi
f1+wN1bANmw9f04asUDDiEWuPjBEXPnZ5nF+fBqxlNgaYwRBvgzWdISZ4x4tyjtYKtVP2dOR3AXg
gn4vJPelpWxpPOitxTBlc8befuMiCwPTvk8eZPbxH8ucqXBpPJLrTTVhVe5u9dgszGQXIgRCpGFM
Pg6jteI3HREFS4C4L5w2osKuHlX1el/QaVEAYEUmtRheN8Soqkk87vtbiJta3SBnGXNLyzd80m7L
8O67lB6nzJ/DUGzP65ST/P9H88WUzaxXaLpkcq9iasIWXSdVBAgVn1PK9xaJHMz2G9dZiuTHLUgR
/awFzXKGs62DFmiUid/JPMCnxGxLk9ednmGKCotj0jnAMqai0PqluwmlQSqALjg47UB92V+r+Rjy
knadRuTQAup1fkW2yUF7xSUnlrg6EAM889nqpVj/ZzmgphHxYKm+75EdSqgYeRW3QQWKpj2QmmMp
IrprtaSRAy9EMcyeWzt1VpCqC4YYNthVQHA1BM52la0UETIY0MrQNd4hRNencjPEbtC5EAIBUIBb
3YbB0bTqgcrUnZLblJ4xi7pesWhM2B6DAguRgQo/z3mPoqnJ6dXVE3dyWgNGhnzCTHEItgK37Pm8
hQ1ravP892j8vezCFXMee7hPgVdQzS7SymjgeIGyxbpVPuIaX9l+QwKHaA6GNrhZg94UXBraqjOb
01O56JHZ1JyFklBxZbQZAH3e60piBF9iecLunZD29zfNmVctWvBT65OS3Va+Nbg1UPO5nL8aoFIN
og38d/O9DGEm05H/Dv2AuOX8n/8sYF0vuJmmIqdXi6lPLJ6GYpSpHgZrywH5CB8YHaJDmEOy+A5G
rbpIBOMCN7ZPT5cmTiewttor7So5aXsqqYO0h/Cl71iYSVvCyNdA1dICy/XjM+lMYk/TOZCzL8GT
T3KDgE1s9Y8vxfhSIXn9/i+4hJM1WftyKE0rxWYEPka433Udt2p4v/O2DZO9+9Q0SGjGdf5ycl5b
orKvccv7reHhQybHkx6W9PVSgT7pQgclACD3jod5krG+ynQ6KEWuVZnD0KPw4Sqz4eyYKU2V00b5
EyA/IsVZsA+bkyl5RltVh09Kle/ZgYcXXaESDFUZYsUwNv6aL/JtcbMofFoAytQS03TVxaXXYazR
XQ+Ui42A7icTwOdrxZlTni0orEn+NmOCqN0Ue0IjQdWVNFAhH1Ovq4jCfgUYGeaVx7l8UE5Jw1mz
n0rXL1fTKRfNu+3qIEdYS3dP6eiHVPDLf9TBypHy+uNf0S46aDyMXvhK+yGytB5G0Iiz198k3+2f
X3yhcImX83N3NpYY4eaiek7M/i8nyNhClN9jiy7RoKu8Z2krmbdYDK+WfkvmBtV7BPYycZ8tfGkE
YhmN7KViey3WgCLJ70uDWVXZzdeZhMqnX2aJ3A7BRDO2W+apv1+bwA//tXM4XmCIyQ8IZPJMXhw0
X3crN5zxuq32sJ5yd9Lc6x6SzUURCXl9P0cVSZn13v4nshWKTV1etgJpnUs4BSegv4JCRQN+D5nb
CqM6/qVLaVOu+CbhzmCrUhtRZZDsAjHthrTdLYq5uAwuJckZBdCXwcxe4oJnTi+HkTLfRnlf4CU3
HsAVnYz5SpBseEKsIYM3KxYBWg89Vvw6w7zSoXtBRHjRa8pg4QVSjQCbEvNkOJgnzfM/CvJ/AlHP
cgRk8pjAMf3QNJ8+FatqdojLJHSgdoRnUOFjRqX5IyG+H/3pfvk1kHK7eQZZJCOqxGRtPHCLdDq4
v8a+KrhDp+iG7zeQZ1fT+QtdZuYawGxZChtBgSlgDEizdRc6UxjYRJGLe3LpQYJnJxr9M+d3bRtW
oM5CNNlIkqcTMYRKco6MA5a9q7G2cnomUiHEqEpPKp6n5hjZqAYzoIF60K2JmFi1b+NpJqrr52gQ
/QYzTIrunrUa1M9eTLfAQbVPZYhBbZQVmxDVzqoVQ9uuBVH4FspIRjmtfq64xHULBSYC8mh7ctex
jnS+GiDExK1EFc+ryyXvPKp+w1rLWXGDTt+GrhP2eDYui83usrzn3yPe+BKxmXFWIKtjAIPSuQWd
ofpPI9LOTwlsnyH+hiVV7WoxmHTeajbd8SDd84bPZK0Fg8UU4bBfWZe5zwHW/yy8E3Mj6cfpaV3e
vf3mhc0X9EWe5RPthAI0HhX/fqzOEJ4QwvpuEtmFndUHfz3Kq5yRih6d5dYcBphSLGR46WYXjkol
ALwAFwVVe6wVXmr1KMec+CEQoY1wXhsut36fw8a5uEp+X7ngM7TCTAm+yoH++Rl6agq5dDOD5lHI
B9WN20kxN1eavDuH8AS4cR6gC2UtIiOHlMHNFevBkN8siJCoOhbAydTIWdxqF4pNduTmS4JOOqQ+
WRFof/ak2pr4zpfBY22IZL5OMChyX0Ugs08MUW+ljYzCJpz0gK1CYaLWXbBn0bp250LiRGFm/k1t
OtpLaR8eImeBI9Tv7shqbGEZIPND8GBdNb7u3Ct9cGflebif0+8nPalyaKHE1zh6Hsmy0R7SBiRn
L0bqm+KuKI7czb3ief1fqmbXmkJ1sHECHyZCb+gqjIZ9Gk/7ZKm+hRFVgpQ2h7/FsVfjSg/ykfn0
gd4kOLbZZqYROYcwGcWRJxFYD1V8q3uYGMtNEun2TYnSSOxDv8+eAXOoquY0lCoSvkXtrTC3hpjl
7bYj8rTTx2CkZFWNdSA9ih9A0497QMs9TnHZrNDLEbtcUlW4vOyhSnlU3ECChS9lxTqf3wJCvVUX
nz0v3P5QVUJ7W2XmxVrDP7emyOOOewu3kIJiD4WgNqVzyalZcQhhYY33vKCqpwHJfdhOE/bsQA==
`protect end_protected
