`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
i8F1Y14h+7yA38j/KyOBjnqQUofey5uqa1GW/qkWtWPNz9+/3cY6zsfqyTHRbwXPM2wNlBtvoC1w
JeewMGVvPQIbGBGapne42lfGiy9P+GT7pYbJtIEyjgdedjKL+pM2+QhG27QYAGV3GVvVZk1zoQlP
FgrHuEUPeOAbBQUJTqNR+PU3r3eVi6yBXFRjqyhKHic5Cp1LY4XtXvZ3V/gKFcrSSIvr/YgxWfJY
aNqcZcLUQ1RuxUqSZ+AI28F5+XauzsjmPc5QXamSXSiB6HHcCFfXl9ck891rwgsKXuNFQ91Nb2Aa
ak48gJCmspzvcE/1NmDSSjtMOyWyR7Q9ELKV9w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="D+D7Z5/a+rGTIszPBnDmJPg8S8UTmjY/DcdrDfJY4PU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37200)
`protect data_block
UTUocy14tfS6taL5yFK8bfPkq62F+XvBazSCQWSQEgt0tuyanMq3DaqWOLJX69e+RtrQ6mFYjKUb
BpwnNFxGltFuM3UmEa6GdkIDE3t7rlnZAgnsIZGAegpP1ZQTPKrYVt13ccHWm5zCQERby/8UC+/b
gkE7T7fYyfq//UlVds7X+AhXl+8ywHjjy1O/DzLQVVz0qyrkudDvf8H10hleC0dZGO5T5vkmqwG6
B2zRCtyIjalmQxIef8aXlu9TOay7i2cZgzZmOOygIu1jRngg0aTs2HsbHYbk4iEboq1SJ0G7gHBJ
ijFedznP9LXXVuL0WhFVB6nhR29WHRatB7IoG+bq+r7dlNpIJGQU/lVyHJEb/Z0dozm+x91o71RH
ll3SAuaMEe6E+WMid0TQogu4Up6lXBA6+d99CnwsY9DX2C6xHyTwiqlDev4X/1Gk1wqprDjlboCg
6BbWLHUUI8cQwCvQlsqpPmQP/QGUUgX7V565ijfzky2FHeTtbM7queliZtxtqDU30lAsqcC6uM2S
NmYm6spFceAZgdItt20DjaEFm8MA3SIVL2paAtsy9yfm/SgIhg47UrN9EBrcMsVIlm5msyaxhYUT
NGfPQaAoipocSVLzgwBuKwGK7BAMWKVHyLinURRIEPEpsNcHRXuYAJi0yOdQcagKyLgGGwjOg1Aw
wQ93L0nBR6Eo7sYzRRXMjPqnY9LT7esw2axWMpiJteJty/2fCAM+asmC2aHc03nEgTkOEgGmXEke
cut4huSHXw0nMoxnyjyeBcVDU7V7uarZOhsOxUxxYDmDwn+KueMKR6thGoFlkbtZKp04fRE+sjys
lpCaaiBCNTk5YoFomdwHi0UucGsRCgMa6nalcUJcoE+NUd8mE/Bg3eJvRZKmxWiK+rchub4w0dH5
6aQfXxGfrH8QEsU49BZcaFV8KxPEee2wXTSseYpHiu98QV32xzL+BMSG5ZvxFYwMPY2X+TiEXssK
aPNENoreiSw+1HNL/aB87BFoAxNU2aCAgTK0ecgs4n+jR7+RKwDKzB/h4198BilX/erwKKUJEF9T
aXwhWtj4ivt7Bax/UvNSHXB7AxLedVSN1w5kxQMj+tNpo/osveQEHZV278Q0abvnxQXYzBusHT1r
3/6pqaktTrdXVX2MexBiNeRFAjSrK+Qiht7brfKGto/hV2TiSxJICD35mXHvv6UvbEDGNf+GkrZc
9dVM3xJhPSLaqjyirH1MejnrzfYzJZbN9xsRflFvDgMe7BoollLS3PHLx+5Ue1GNj8VSws2ttfOa
W6adGmq7LCJDrLVHV1w4X6l7VzCdSAWJUDfmFaEoslD/ngeMrgtG4L2B7klda1QmYuYn+2jn2o+T
IYk681FwJwHnoqLiL+wHNVBaubSxNpRlN/5XN69lADvv4kCWzUt7Lh7xBNV1tv5iMYKj7MWkZyYO
dpq/zPh4XHfnwYvyps3EsU/o6fsZiQa++w+28Nalti37j4ML8rKKlHMMoC5Fklz86Jr3j0j9PePp
JSsMiF84h3lwprMAwPn8neKvNBbJ8wSh1h9HOs2Sml8j3XJb5tsjFhDqcMWTg7jnC8hDsBxv+zaJ
IcSOjSLeBprcgKKJpiAMv6j6eMgwv5lhG+N7AY4p1/JU9LwTx/kJzTXlV2q8LJm24h/fEVpN7LlN
RnzC/ic6CduF2hBnfXmhPiWgFIT2G4fNI8Htw58G4FaBAgQjm4+bqdrHiBIaG9B4mPD2sHsJeR9N
y96qRnjDqnZZ1x1qbWWNJJI+3Tz1R296Qa/us4ecJnstYFsB6XLKZvBETaOcqMXxBQFUGJ5cpe91
7Ff0YN2M5qaK68XCN5mr0L9aD1jCbb0NrP9Apso0qgQOh85FWpZ/aGmIpbg0EI9H5DAwwW5tpKCh
4abK+lLN1wPOIVTzj/qTZodexSapHdVLyOpEdN5MFigjBdRezmZg68R7hCgeCJWM8oMk2hLwzos9
FVFy4XsBJbX2GjhLQyiKsz0zZVn0rTwzmxNed4kVlxYxilqr8yzs0brKyipRwkPr77n+QH2eug0I
OGxMLcQzHMD26WLy4SFDL+9omWYYzJo7KYx5b55lA/zeRAjt3pChdECjU/fNWQbWsqq1RMA/ADTz
evj4MyfGDi9pB4ixs5VSGhHSnZXCCZyP2WVTfmHcHcWum6bnZawEPBCb+lHGJeXMi2AT72B3UcvS
V7XzG3tt/au3Z93O6sbA3tGBwVgxNerWrjhihy0sfWT243u7crv4ERgTNTLgqh+tqIz8LgzOp1nU
DC6+bu931Q+0hr4W3ExjcG/ymbJ0+OycKZMPnhSB7R+0sthVAeLgtfzMw6d3zggkot2ln3llPAlZ
5iBWdzqwMAJ/iCoVa8I4SihPqA7J5x8Xi9FBBaUJddjek6aIfcXyPSMOI8YXG5GUbvgeOpQ4kf1m
QFmUXiTWpiFF7BsPQWz36tvG4YvhsJRf+dTdLnNcgRdKEjqyFsWQSgcraDYpY/Al012KJlc4xHPY
deN1UnH9GCyuJ2jtFRErIpruPLkoallryC5OQNFVI2rxD98zL+/RwzrCzc1stRX9DUteek8a23F3
xfvANl/ucoPvTDdfsyBHs+Y6FPMk3z1m0k4p7io8TdjaGHl8Fdx6mlJR+7kUqItApdC457RFloZt
uuagtHvhysOntxkD+2+dnXBMnz0my9+c1cIuc0MWVcTpinkp2pSQouKIKpQH8DghJmvy3Xh02YYu
iBIoH0nzL9PVcYRngzC4nlR1ejToUZWuigY5/IqGP29/KI7NCcHItQbs612V8c9F4CGNBSZTPdmB
6l2N+Pi0XJ3kKN6BCqgv3d/SestBYX5IXDUBVkPZmqUk7vRYjNneJ+T4t0yzlfnSG2azIvN6NntI
o3FfAV4oxqu0hq3mY4eQJK7pNyv0xc5g0N+zSjS64IY1fmxEME1oPN9skK3rraae3Sr9LNlBlCSE
lIL8aTC8qi/eDwzIfmBROuHid967kOxvO+erUUwKGtk+0qj2dXawQaeImqxDxzrmdYyngy22JxqJ
f9RGYGJBLkDC59r3ZuDMLiJMGx3drdDz7gbeyjm9AYm3IxKf/Dv2EJ4fJZtsXowo4009K1QQUhNg
DQVXxlMja9DtCArYrK+b/pESlAQjTgQpIb9qD+fVWmXZnaKsjDIBb1SkVJPATc2HDB3qpxsZKlad
QzT+/YJrdzWVQuQlj6MKkK0d8jBqfBr3aYVvwxCiyohsV8sJ30Ky7U0EmbEybwdKWSkCA6lLVAso
JE3dOL3+mL5gXvciFM8MX0ZgKJ8y4fN/Qtfb4QkRWdmwSQf9H3wsr4+VRDrGCdoROGFC0MgXxfqu
ykQ73KxNG6du2uy+yD4p+a3JEsdI7roc8x3IyjLuEiOOpWkTP74nzBI3EurT48V7oQ5ddT01yfK5
PwW3OGwavLLaejddB2Ko8hOpPkAweOhr27qaCzqJWyL3BsAtVB4Qkbciv0s15vfyL16QS6pW3iSz
HQnHz44zGdnJGerootGs3zxNkb+VOTMPqlzqRYOW8ET/D2lia8Qmn8fyXnmYB3fTl34MQa+8k2vd
C8gejfQ0TgKrpaiQ+wLU+cyaTEr87ltCuXULKF6L8enCuPSOHrMXr7yevOtr4VvCn4X+3e7m1CXp
F2hJwdm7skTs5g6PCQDxDJOqhmHXe1dRoRgdTlsUCdpwVg+K1J/Ey3LaUEbtkpBMmBEnSzJMtotf
IX74ToMLQ4w6JVWgNv9HZkv6l678daoTER3r3cSKPKM8P8vNRXVMBSAU+0v+IIU1d92muVCB+ZJt
UzghHxQc0+XVmK4lVJslHGOQYUD5Hs6ZGQFwwjelW3bws83d9e5uXIAGx4KGChBrkAI1YQv7ODHD
w12r0uDyjSyJyO3DpRr4gtBab+Un4FzLYENF2fYPwtVCj3NXIxmsfnLslGw6n6KPqWk0yaIpSk9w
HTorQ11aqsnYJHfmpnlCN1T7M7LbOkOVFWdOfHkB7M2wTRuBdqeIxFmjCZRWA0uuVFawbkegXEo4
yeLoCRMJtEDWRGWoTtSxE7XMl7mD1tECR922LGuOci/4PYhoooYAFI/cC5zwJt/E1Cimij5nGgq+
O+w5jwE7OtI9xnht0hnSV7UVypRvtZIoC5/2rb9NeQRkam9Ipkuet5q+EqNLyflq5aOrr7uESDCz
LGDxMoub8vd9/M6HnpZlPWRl8f0Cv+qYVlSuprgv0/cOwt7g1sFEhqLgJ4X1I+vtstKsqBZkr7R8
BVzSr7mgpUhIFM9LE6WonJcjC+SGRgGvFy8vEa1ebE0XJ0+UKfApe83GuXkk9HyTIucbnWCTjgaz
MCLRtYMu8n2w/81dZc09QPZqSBRWRNROu8TqbfR4FAj22sMZ/DwUidA3Nrvs595HfmeJODr9tjVD
7fcN0Low0EWoK0FkZPJSfRLhOByjSnXKmIk+k31M0LhUcCCJho94sCkzrK+MvconeGnpvjoQZp8v
PQI0SSzh4UrwzFX1CnkBeBAz8Jv24YdYzJCsI6S3bEn4IqN9Zpo1+ZA7eaNu0mFnd0ytjcNdyMnL
tVg28/P8GMaTdadNHwAEs7+fvq/d/B0yRHTjWUpuwLvcfDnISAn371r6mHJXEWqmjmpDPRoYrEgc
YGo25pQtGMhCfIqvcs9mm/FxBAd7XzFaxgX6kWF+XEts5vbDe2zsvhTv1DmdiHUbwN6goi28mV9P
aYOqK7XcLlb9yEEQItq4AUpKn+6bahz/MiOUCgW95hqrsGYfb+khGkatMOf22SmLbugdtSqEJxO1
MawRZzudIsmEvB8hYAtSEfo9xA189krhg+BfGM1XBNTwbLfyak5xZafn0KNoiTGy5Gs1KIbvVEHx
zI2z4yZ+X6SBYQ1fG27QD6IhhDIaQ71144wYFz1A+vehFEOhjBfnsYf4T9pyHgHbxrpwrfdK2l1M
Wy3MG5ue0zRssKL3QQI+UwHKBXLpbkwAJtKtmet4FAYNKG0bVLhRxf0yswR2zIeGeM6HPlGF26cJ
FX8bA3aYPFMtakHVyvJL0yF9rdSdNOcHg2pXtkb7Df9hjNPNyuGyB3m3TbiqId2My8HjurN9Gsiz
jMyJJYwRt1tz+atF5mRLyQt1labDbVhuBpAdhrDRjlWHzgwm8i9N3xA+bmnRzo13OaWNe4QLhctR
90TiWKHeuCXgxiuswDnubuut1bSZqj/KhYECOSmov7jzgR++Prbib4CCs1s+tyDqFU72wj4pTBcj
GYc2bFuS+oYew98RMWYRVkcvf3zY29XN3vA0dW90more4m9wK4F4rlkjVP/yZ19UJvO3iyBqADS6
QbaNNLRRbYYUp+hwFk6cTc/f5EY5bQlwMjD1bawTOExrZyyjwLKfhqmR7cRjbOwlcv8I3tqR6hD7
epqWpyxw7v9L0K0kuCVJ+B230UUWfWrvDvUI8VU3EqsXHRMf5p5eR4MFCYdw1nguTFxYfH5THnEm
xp93Tl4egRvg5UcSrABxALHBbuC6bQfAN57cllamRnL8moEjsYIwBxD9Oh5EqMbdpcIJ8TS30py6
5AK/JsDAMoG+lwpTGyfdxrBlH8LjzqHPSZLXmXxw0K1nSDyI5M5L/CXd9eJdA8ZDvZOFZ9D++ojZ
089bJ1cou2qyT8d4ikO9/qPbOYQvLyGbW7GoWSEY36kRAJGpYw2abxBT5MNaW91uPn/YF7nq/snx
tNx4Ojz1yTTmFViRyNLWTMilN7QVktHB+86wl4RQfiTn6LkXy7gJpoMeijHGiY3b2uLOzJ4x0sK3
/C1wXeIvcDeW5vmv8bAZ4QVKrx9KB60yw5I6JdkjSdxXgNKrVBewSWbdCs96ywz5nenvkBkH9tE5
nwk+0Ab9WiRH7Ky+1N+8uMDmeXGFATCzadv3NilqNhI8P0jckj3b4XM5vh9+nIsA42KNctIzQkJy
Lk0QJJ9G7VECJ89YeTWQhdTPob4D7/91hCY8abIxvCSJT0WbOOT5eTQeoGH8eyQKxf9ztg+Xit69
t3Ffuaj0Q3TL5gJI5fGrK84K69nZZLWwtnHidUbKGMFD/NeEXkjLk/tDldgAaHcGBdP5negwIRni
JrIXT/UHpzTXnLEfmgvaJXf8JGUGBcU3wnPcRFrKxqL2UpV53VU6LNRuqkmhmYqse4hUm4PufET1
ZanTld21JHGNESizl0FynicRUE/MYMmDssQttOLOHhmqMlkVdAnNHiWl2YYhqkBYeqfg78KffpPS
0/mwORkTiPzyzJMYJzUS81guQRKiqkdGWxfYBF0ubH/ouEACPE9EVeI4cHOqGtPNv9aFY3Sx8mLf
g3moGDfKPSm4ge9NEgZ72O4F9vtUnBjQbhKI/rI9pe78JDL7m6XhTkpD3rolhPbxlZcCjBpBiE74
8R/ZpViCUv5GEJgrEnHlQtfNe84n/0+eoc+f94J18Fu2cq5n59xCBNZZy6Qqb2wuJzKXwB5MeQk6
ggEjMraBKWIFxMp3x/A60ZHgbEmNbQwb0uzyLNHyDUV9j4MTlJX7LaJoZGQzE+QFv5WX1W+Fv+Dm
TGJGRvaXr744fMcLBNuj83F0SvATYbHcwiiU7VmjkLzXF4ScsVbFyjyQy6pLG+bs52FUxsbDERpA
DncXQkfbWhxumo+Vl0rbBbYAn5Y1BSlkPFj8Q/66TEQRdKlv2PnVo+dOur7tI2dEL8hvx0FP1Pdm
DjFZjYTIQplvrvjbINdwQNPha99n2CN17UoW0d9S9/meB/nGBvakzQch4ajYyDr0YkLaAF1HLtNP
sCxEFLs830Xq2T4/iYgTD4i5Zc4eQ9Z51FwMLlr8R6XTM/PTxh5+Py9QoCJs9Kq9B9PQ/i/rpMgb
ED8gOnJPTzTI6JW/BSfdkFWhFfx4iiMoNCtfx3QZYWUvn00lt7+rRNZKyZ+tZ5UHk8Q4s33wRRSV
g+hswf/wr303SEO+BM3RXE0eiqY9/w7Kk7x2V5lG/qTD19GjnHWSXOVp+y7Q38N9b+Gqbetj0HxY
ItNF+Csbt9AilIkrfsvp4hM2ABdbLPykqwn3ai7VUdRUKPpUyKPg2PBOMJCXQdjRo0kDTwx8iTWl
C/t3bLOxatCG998iZixCMCvHtVrkBmCUro1OOIn8rFg11XY/nlkMb9ZEg4hi6Migyd5Euv8iPmTC
3UIoIHMUiu7Ty5xaRJ5B/v6ttPFW7rn/euEXurjAfJ5c4yXPEGYGo79mEFqh5xN1+y4nzUhsJH/o
3/YSH4omKHNd4cfoJYu9ULnvS5e8LlsIIwHpFkZk9UWNN+VEPiL9p3MJkoJson+CyAee3qtCpXQN
YiObZ7qLUtpd+52/RVMy0I2y3z/hFPfyHc5VHnCDjXv/MsDA5eHT3gOFCp3s3uJ4ymmdmyU4JUY4
xLMU++UAp+Acmx8rPEi9qdlA65OVL9iiLKt6Hze/umVXjm9y1bl93ukLqkprSqA2dkw+aLqyUIgG
VvLaHcnj/HojULAhZJ9sXXzVKncFjvdfKWIgdncOtJnikp/oLLbbV3Keo+GVGgKlIYEdWLL6plwA
yMZyjAPNqc+Xbm0igr1R565u9lH0e0EP1teac2ACmHzvXfAw3Hw3A+Zuxz3Y74yXvMYz0EjKI2wA
PFfSZYzN4g3fDcU0yR49iTu8JV2PuGMtnUIVpdGl4FawZviVDKL/4O+k7g0n9GdRbFxmvd95c44Y
SzLooJsmWV090Ui4Wu8ZCUIkK/ByaMjTyselTgEkJ3NTSBa+4KRS+4m20oxWNnYEISS2ZEPF8ktY
wRTLMGZnmIbxsKZGGNliwpBa5Zxr6z0xZPm1ycBrn63KcHgN/br9Ly3LkewyxyLaX2Wwy+NyS6fd
1orTy0hqBovuyRCzQFkxIrkOzYGvB6KRphq/JNQMOxocGf7QJJddscuOXPIfgrYQib5AxgeZYIA3
vBXmSpBlW9lQEy/lm3C+g5Mj8J2l+oyHtUFnJQ2NWYRo+h4V8iiD61KRfbmsRSrth7g6jbfdvhEx
grQKVK8RJKm1oMDzTlToR6InRp1LfzHfOTamX0G38dvxlOe/C5qAeO/kD5laqvS0zq+pRdWrTH0E
LbiKPSuTdGY5KKi2I0zYh5UGOj+CNkHXIFI7zuIGF65BrQsJ+yfpWvPX0gcfdej7cYFwt1TREa8/
ThpWsQqEMMlxD1MQU62RPKrywoMbUQpRQzp0yNMo1eC7rq6AWZKSbz7P16sxJW7QqU4N0dxa6pKJ
OZtQrc98vseIC2LPiewrARWdaRAyL9kX+ilZ7mj0Ewr2Ya4RPwCgZcRYNcvc0INI7XLLgQq920vr
o32xwlgtjezRA86R4RMVoysGF+lV5OTrx5AfZ2WU/zLuqIZa1d/heA2nUQzcZmLJoA4pO2RjFSjQ
PFzk8LvhJkUFAnktk6fBgjndkyvDu9/U974A5gRF9t60yHDSYdwidgHpZ8kwePpOnPHe9DyxDvhN
IB8JxyIPgQpS86du+YzsO1JfMgXKssTPYPA1LLy5q7+yRQ9aNk2jr71qnaMmbFULevS230mY7iTy
+aLvCpgG/kZ+KQPtIzYXH+mg/HEZYL52UpBK/kor4OLjuWWTZ8DzhW9UvxaqoGBMDin0dZu+lfk9
+P40jNzY+0aaRoq5hjLnVKU7GSbbYgGEUWSfBbaz3uzvcvwhUKI+vOUsTKOiQwcqpcmLsXVFyG3d
luWuRtCuzc9907K5e+3bhsfGKGFzJuqt1kamVwWLMEl69FZL9Ly5x6rCqCAIpK7N2VJ7bXbs3Ps2
NJWhl83FcXaClqr7pB6wldQRRktUujlcKjm54EkRhsjG4qBX/Q8EzKH3jQFGDfO9LfWz2Fr6tHUW
ifysFNMF4Csl3Llo6tgjofYWG8h41FvkJpEgJg8AfnbrXjKG16m1Eevq07XXV/XSmll7yIQw7sjE
KUNkqrl5nu6T4OfWUHr4JhJ6ZFaC74VA3o9xwcKG+Uzqdbdcjwh5ac+T5eSyTe88huS7N2hNpwHa
h7rc/XMAb15ENCQ5f7hJ4rhJc9MrP0ffCWnMzSyYFXSg3pHF9jwEFtlB6TJCrV/CrG/GHh0J71cM
l6f2hzGBT7fE+GHUDOQ75eTAEWozfNN/qWChj7Pg+fioAvohEF39o/ptppfpHK5zTj32fhO1ZxLH
q190EIGwN/VdiqW0j3crO9kSC6Yq/HBrkylm09BWqqPKeJCNeHVraa5RzZ3H7U/lzwwRqBExxOdQ
H8qX+Q3estflth7v5eBUjr0a9Nny/WFVVD2Xh1jmsTXEY3zXe5dGW7ewQmzA+7c6QLNOv5P0qBE1
quM5Icxw5DAr8Nc8Gpqt8G/oMOoue1lFqW/5mUWxSmWSrarxWc+Ze9lS5tJlDcf3DnAXhzEOogw4
zgpqWn4f7ky2IeHV8VSpeHHnDcRkdgLC2czzEKQCWYXNTVtwY+65dkHpDz4naodcZ9OSqOIq57AG
ng/H5dTJ4ZBxGQl8CdhteYW1yesUkaGJ9Lxl8wgI7bc7PDyusxgy45iJ1HOYfAMdJ/V+XR4CN0dg
AzBMv39tar3Ol9hWDX2zeyurTg1wShl6A6KyeXNp8UUxER5Fquydj4Rzu/Q5zBgIPdv2P9nN5rlj
6lXC+6ISXyyECauRWhKFugsdK5VdrSP37WoIzuDaxdpsI6jBq41TGR+k44tVpJitZsT8kI1YTb94
U3JC5Tswa3ES2VEDDiGejmhbxcK37HdpGAPiTh5YcpMbnoFBIzwwrYE8QuINZ7YjG/QkiiUJwXjJ
1+hLECMF9g1i/I7md8hSUhg6uWAD0fdvSmzDMYvY3scipoU+rD68wB1mEihyDV4GHKp85XeOrSzJ
748LWFYioF+zaCccct/h5i2pY9HyeppvTtVO5tVm6ZDGXIIvQp4QeJrcQPFPSkVpvfTwWiSIXfwb
seEVl10+0p/0KX8V55sT2HjhvJS3RX9Oex0Sr2Lpxf93sLFxTAQqhOxEvkbudepwvhar34b0jiJ5
M/B39OERi+Xu8PXQojEyGTl1nyX+J7Vy0My63j2d7Ww1P98YLj3/4KxQsduAexB0ovDzRwpG4Zwa
6E0Yu6Y3odfNIsP58PX9YR3vTsDdqvkSmbbSML5PfCAKxil2JS6Oj43v22TAvqhn+rJB1ev61YtB
JDfItaaOA2SSHXrVlz2Htt+PP9pLZizxqQtdmef4PT11SpigSZfbZa1uHx2n3iMtYnCNUvaee8aV
GVJAtmVE/Wk5uQ1QbI2J1D3sv+RrrLb8deJtTjr7p9iqnF8bbwa+7nHKy+AmQG1GKVnLK/ewIttC
nTHXGa2y99lsRB+PxCPudFJERHmZXTve8U1L3vxYbEnUMUmTriUanPfmZySbG1sxexC/76+JO6EZ
4BvyQmjdN+0pHw4MhIoDZmXv5utl3+ET0LAjqfoqXYEZPry0ISPzCnzXO+hjkyVSoANVhv7GBjpm
ijDjv9srDZqQiN03XKk/uwVjsNplHHJtSvCpETi9P/Qt05WQr3WyIFYlHQkM7a+IpQOjBi9HFZ6K
zw3D5//7p4YAGixW2mDAh2HzP02RhnvIfIDoim4UsQL4yC7jYBrdjg3BmTAlIUEApSqUw9+g4F6n
a7wlGhxJseN0UWsG5pGfDPFDsOtVQRFBTdku0+BmxvLY8KKNv6PWvsfi5gL8OsnVyA4X4xekRAmr
mNt4V6ttwhlHhYY1Tx1VosZGqEjxwBSH9dlMZRe9zAxuBgyipudYYs+FvvTZPhr+w7yKeE+zLv1k
H3gzAkcmUbdaoTeqXsGD3GOhkQn/n2bLpbyvIl9z3Ww+iZmJ+/rd2iuN8Ljvx958KQxdut5exoPj
9FsUUyXK6qaHU6vTmrC38qSU+G8V/ZVUNBhgOvi4pKs9ZHAs1u2txTfC/ycEhBkrj2cBiRmdb89W
VGZHgBIWGdh8itazX9VSt0W/CEjbLCTg05N9vqyoCkAPwQFNjTKQT+DZbbuaSzgazufVoNB6beEE
QG4GrAmX6Ro+lvXpuiGVSt+7Fz8sTuY8FArqc31nyy88JyCdVsJKlgUY3rT5P5v0fQTky1rYKbZ+
l5M6IFsKGDpyDQngPWdKwlOldZasb1SbRQGPVERmv0kfY+G0FbgfQk5CB+QQ43alrTnpFXRHg7jz
86BxzrX0ilyrbQZHp7VVtENQNskvU9VjLHi37N34UV2UhDkLCNuDi2lTGcqKyet/BkKd1VESrT0Y
xJiWf9FbhwlLMbyyjmE9zSsKXY70qT+LHBcs7UihloIjcX042wircue7h9W4rNHfY6dcYvRG9nQI
DitHNUJAZ1VFbIcDLAO3clsaOZitfgH5t/7M+wHJ7MRBH4dRAbtCPsYRjj06jV7e4XXjkx+lJfuH
1ON4ZEWqf5wXhmEkUC1BgFY6wXqbEKIgyZhTbz90dRZRsByeWqq6EIvd8fvkKLB4hsjdMPm6bqvG
p9mHxYBu4xhEuJeTestR7YCvFzhH+8cQhaGXsjy1a8zql8iMGccMbVSbk5mvh6l2aQE1J9kwqTxd
NakOXyFMyxxhF9C7pDiT52IksN3y5J9vx5TL0np5eq8NZzygssIWZQLQdZsEjZYBpLEebBnsv8bk
TJDdxsXbdcYsTypqIJczqWDiws5Z08GauzWcCdcuhaNRG9MM4eD2hKsqYC982BXRmTngSFB6Cs1g
mGPIu87yVs6vEmjKxO6hnY8t9coRT5Ed4HJve/D1m1RzOmN2Wb1rue6IZ2uC5EL3JeGda5O4eLkK
Pg6v+OgFvj834Nzd1mGz0s73xK+ufYthyScMNRQFW1uMz6unQSrffbVJSJL1LTJYUcxU9HI9k3xt
n3BI4d4DQj5OmXkHcqaGyX4E/LDZ7mce9TFJatVflW7Wz58mfCCTBrxi5RV6sw6djnoauwHe+tGD
m6kkwuhSqyYvr32NqOHJnjIRds3hbTfDXsYMKTzU8lYnCxD5HiJ6Ei0SKAsFDuGHJ1LczK+npSuy
U9cg+tvjssM3x0Jq3fJ7iH91zFp6FR02zTrYxmCkbHcqE3zIvGBrLc84mW4tCWe1Y1E978ztyaUb
f8olNpVElHj3sQe25gwHrOARnii6gL/c/pvbqhgMne9jmZS5mOhE8gzs3vAc88Nzb74NMzdnmAv5
KSNG59JtpUiUm7pPqvmdXOp5ASDI37dsdrRdEoiFNLPfSVuGRHKMjmL+pPjicSSfqPVedJ3Mju0J
LPggqMQaJEK6uzKsdVdcxfyD3fayIVYAvLtIwFnYrD04mwjQ7/fsVUgzF7daPeyFC6hXy4yhWxsE
XgCA/73kahdzAmGJWIiO3eRpUCHiMrpUVxEqn/tqceQSKL0tJi83ugCbex+AHdVfek9zeBeW64OV
qJy0ZL7cw3/Fhazj1SYKk8BTOE2INMuvcIrmNpVhGY/Bs3afWIyV0QuYlLKVwnH7VyXwSzud2TMV
Ffjov7V2tZyjXksfKNpbcY7UkZZ20RYeftV493Nf8okdqpp4yGXC8zLj3K7d1ccILsBMkr5zLX8k
//kp+9CR1KwwWdOFAFW58aL3lSqdNDAO5Srjci3dnwQcySo7hOLgwGddPnXmk7nx/r2BcMaTcUzF
gh5tninTp0++9MLmBu29KbSirJ7HRnP0YieEO5zffCKaHRRuaabaLNlghMwgLJUq9jmM4pJQPFIr
QldUrUDP4VpGWDYGaOYCS4ntQbbmVQfyp87CpOCW6w+hly+wk/+dZPccAiKbs8xnNeSbwa7MLpvH
CddmX6sRmYLkp8ObhKQNmjfLQ+1Dk+jVnQkfg14C3nCnjhQ8UL/nLovEi6NqG0RhlHVC5u+seEE9
lNwQHsY/fRcy05XxAORVecwYRmDZ0T1CdIl+5WaZ7ekEZ/r13kIpRkJ9taxQIVd9Ct4gItdz9xof
Sh3EbQUJ/ETPVZn9xkjbR3wrJhm7pq4xA8CMoONSRPYjnVFO0z1Ce2fqYT7lXFjpr1mRx4SXEK8x
tVEvo6M3T3g2kSFzg2+TLOtbolNot8jTaMP7ZyUqA4/Y1/rO3wCwJj9oY2cI9H+Rv41zPzE+OMLG
k4FiOb3+VCCwE5zcCo5ELgpOTFTsDxTXCSr1qAIBwzppGwTTlwLR6gARZN3M/3wFRywViYtxtEOt
lHFO/gDua/txUtX53yWxFA6hvBW770ZDxo0Po9RHBWVmu6ZNXZS8JBo4wTKSdYQUGrmH/14f4oaF
1VPh2A7feAzTaiYUD31Q1+TxawZvhi+Aw+wGtwQ9qg+Xi15fXA9zNrMZgcW9DVmdS5HcUD5UfUUI
QK+Q2EpthNdUnjOL6w+VkV0GhJHtjj00BIW9wCaYJFRwNGzAa0QrqUhmXc14tJdkM6QTxQjiKJ1y
gVl2Tniya1Ypd77gspdEQ9SkssWa2M4KMGVDHYXANTfkqKk3bkRtL0UiDrqIhRrC7J5irDN2sp6+
VNUxwgqqsoocSDGklG3RDDNSbGSOvolyb75003hp8zC+UsoP6MhzA3iJ8H0IV+JZpeaR77S1cGQX
9KRa2dnDtJg7FlOnDqhitel9ca9Tr9GwpJYjkz1IZSIU1xHSwqsD+I/NnIlXhpQhVztscObHy3/V
zImWoWXdabL7d89hRQzzVG90go1zRa+ofzO2aLCKlPQX1xaXlpQBgW3QohXp65xcYIQ/UKlic3qf
I7wAWhoyntsDt3RRAFOCJ9COdYxpezjBM039PErv/P22sGMbrdKrXtjPG9VRTu/wVYu25shJR7lP
HtKP3XfJiJKqCWgoRJ1NEQC+8x31ABVcW18XyBdbEWas+S5oRZVKkUXP/lJx10fJ3Ql/loeixyIP
/e6k06qlwPNM7pVlOGQu6T1/q20Gix2aTXnVMbj6l+Sp2rcopbTHjL5r4JGQCaKWkQSB4d2oaWFl
GP9BKxyPrG8q77VPkk9Fzo85Rv8CdAD4XtdHhp8ABbUARI5itg1UuB2FWw+OZm6vpGYyMnSRqQf0
Kpeq+xIyTrj7jGC083XWpft2G2BaNhCGE5cevfkPKiCKSLw7qo4cFBQX/TAr+DqR+vwoRVoP9Lsq
vGb9K+EVEqr4dCX9J5g+Tvs0KGazdLE0kNm28WzSVoprF4Bfk5RoCyjmA4YlKP8W0Mqmcb4m0N5Y
SqZupYyT4L4+9rmVopGS66QpawBDkCqw9IHV76jqV2SsF/oHKQYDgkqaNlAJE+M/vVX9S2jVKB4Q
mCcxQqpiOjwdUkzw1kW0IHleKhyqS4Ts2ouSyIBlsTLJM8+bcuW0JdWyB00zJMbO+4E6VDv5EfAJ
4Jc0ybseJ3uqzR+d292G6NlBmG0/mzg5Mvk451liOl7kZUEDBirp4gzki9Q0j0anNbS927Ry7yfE
2SZqb3mX9E2BvWsIIDFCATMm975LWKJja25K5lcrbQoDzm5/EUdCsrYNNnNtthziKLyPHurd7K62
qGMA7zNNWWi2N3JUl22W/pPVdPzAsXtUmqoPkV4bIL32wkyKXI9SoOQoDWP8/9cPECMIXsE5YUV4
RxBsKJNozxW3Z/CudaogRaQCP5kHytKfzO2JPSab41+P4zoYaL4q8+S5BWaEnKCo9DGhRHs0lgPt
trToTKOreSuRIK25XeLk2c4gngDwUdeq8P1kSzyl6d84CwqJVTQ+waU748VIdvH+/mUm5JIaSPXy
xuUcXy9VJa8F2bCub54NRvlvZ3OXpPgpzbmTCpEKWxx57j/UIUWzMlKqcLdCKKm8Ea6HJ+KyOeCF
tDOzrU5flR2IxN6xxb2p81n1uRr1mn2zyuti6YbNqChTGzdzlIBHBaqdu0oiXq8hZEDOuDQIPBcM
M8SCaolNherQzUbAVDmiWqFAbuaTYnD2TJ6mIvoDs5YVc2BbnaPWEMyjpBm643+KndqtmNxMeUpx
fb6BZ1LfvWDAxK9t943NA1/Lq8fUptKMvy816Ekp4OakYzVhSjF/yRwywbfBYfMjGViYAl65bxwh
sc4YbzlQxlKCgHQj/tbvLsKGFdp6D6um8PopM/B6y7DEp5qWJH7QL0YqmmCsS3C890KJ9m0IJ2Kf
r0Bz7LBEt80qoGuzCDmb6q4QVTvg0i0icV7whEP+bVZ/tjDoR9C37ouB5RFqi3OicYfB2PLxO/gR
7Mw7Y3+Yhxht3GEgD3dq8dxkiBLjFC0Zwb2TFJSQQcohfkhB4qvUZsUv+/Iq7FpXc4xoowOdvXg0
DWhehudl+A1AfO3QlxXezHYsOtaRdtovfEduoPMgmL1G8f1ljvwWJRxxipA1li0CcxBPQRvrK9Fj
JJtEX6pCIVoTMcEGQ6irJ0eFDL5FwhloIInk8ysXJyAUN34AibFSOvmBIX5NGv+xS8h1m87O8B+1
sJbeiYXj2UUO6C0at+1kboIX10wYA/IXT9JmaV4Jv+NeFe3itEawAsZ9WwjbsuRgU7p1JqTzj31C
sjSE2S4YJ2MkJ2d8Hbywmvs3TMgDLXgLaNfdkzinwbnXOpY9IX0zrWFjHIsRmXDX8DXjO7x+PvxO
XUj7+qUlaJR42Tzzco0KYKWlRYua68JCWx0dPdCjxAGmUYmhyeGOkR7Xposfcoi2B21yIeRdejGd
b1tuleG/+7vhuc/3ptGVFjVnnVf461JSHQ/7kbsTa2FgXyCJjr4ouxupb0LtDYj0h89/UdaHZI0v
CALdozpEpo2eoeJ8FKSkb1KloKYFf1h3+U5CJtEdKpQiAARE4JVnp+ZwkK18wa6Y9I5EanTOWo3Q
ljdR7XxhxcbRgatAY8KhJYE+8wgQLKRjc5eb5rRd0MN0plZg/e9ioCyfV2gwMypoNXAoJcORAnKa
PwyW5+u/hYdDd1u5AYU94vNFAcREONrr2R8zYCeDWFhuVuLM/fMN8+PlDUNBij8Ei84VtCHyHqME
5ET6wIu8Glyo5IJ7v5CXyDcuVxpbF5AvtbSuGDPmFfCEQcazXPego9P/SWBKtcHiaDCs+5Fyv+nV
rSgTbiHV3BnnecavubyNgiBV62lnDRkOFMM/7bD2rLiNi6FS4zv8jGjzyyepjFFcsMZYthokJ/qV
MdDASTcplpiL3eXgPX2tP4VdEc4y11oas2zk+twkP6RcOLwjoy2UmwGI3w6vPMQvzOhOL0p0R5ra
cSbnJ+IE/id4NDndkYGAJaMGCqfOcx3RR+h1jjQJMg/R8VTE9RdevA4jS8UhIO5FiRb/lFXaIR6Y
a5VzRwg1orGk5f/N35yOIiiSuKZIgtEPfkxJ4gcUk8GEBweT3iXoCKCM/x6bu2BE4tse5ndaw+E8
MzQJ7cZ6lNReEw914xhr7mnAkKq7lcmVBMaEQEf6Y5IZjg+MgStT0ftyLrTE+dL2pKBrqfQLfAzq
w1XinpNzmqT/VCuKkPkqMUqaWeKhgbUiPxqXElHIkdPGkiTWD5xwnm7BbtMAKr9FBM6M94poEeBc
bRfiH/kswTOlkEpK8ZJNGpCEfsjZCc4Dem5puQtG9RNS1gmFwE8NdBle198vXoLw+oG48FQMMUbU
SbMC0EHXZQSNKzWzUZcp3uEVPbPuZfDpXQmhkidPyWV6yVvEORThF0jdWI4nPQU8X8XbBHkTZQXC
Ss+UBZvaviSlMAFzCMjm6nIn1yqrvGTMAPYl0sB3ZRBWFTYSdaRTB+6bFCLnCNAbHU88C5eXJKCz
vEfwxKz0WmuE6pD1kwMIBItDXeSPXY3vGc+ZVHo+ka0YjeyIT6oXNS9l/wXUQt5CHFJ6qfnuXJCt
ebHzqs0maA6MP5aVwxsBJ7pEBiGTsjuEGZqIxaNdK8SpFAadMLAQo/trminiGe1gyeLYJrOPmewT
GvLWjzPcd1A6cXcXTtFP2d9q+Khm1jQb+JdifbSXVeXkBxNsdbKQyI5WX13smPKeanlYMANnM6Bn
87urQwEmCKlM0FI1zgVzr2OxF+k134XyUez5I4WJNE3Bx7+WFbsZ8u4bmuwt6mksSDcmCXG9KH+K
PNYPf4fx/wLlP6WnsqHe67U/5/aQM0kn/xr02MSJ9VVX6rdfqqICgLNhOOOUVCn9V0SsflVoIMNp
/uqU/Q+p9dLO/jib/+areWsoAdBhK+sfRDlWMfFi3+I+G1S6a4MFbh/RxKQS6t0APXsaLiwnfryR
mgdUIYcrZc1mdkrIRwmHqW58ZAZKbl8sY2Pl6wWlXQ3a5NvFVvnZ0xdK7XZ0GIsQMwlt4TSxTfbg
eP96xxMqm1Y+or2zeGC62UsRyl8iMekkJmuIpZKtJXsnxovWD9oE7SxcV5PvsLOydM72FxDkvezo
iqBXVI6iNe+MCeh7eiNDqO4P9ZqFxcfd9vP5jrCxHX/Hn/2ygNTGCrG8wq8PA3H+vwNXOW4Is/Jf
EpBV8qf2BPH8JT4XxVWsBMcDzGbtTjeHMuydBS+c9tO4qmKkbx8O04Bgz0uo/XLJTJA5B4NTXuEm
PN3Ewvyqt3ZGi1KIqHegMNumoaYsrSeloWe6+nqMJ7kogP3EVBzgnr6AhktRPtmvhBQje1QQOWRz
ID+kfeVeI7WAOsas+pLNNg/KsRIf/KaeuCa14hWBQ6PYBK7L/3BpDIQJGe6bGqv4V3rtpJ6DXTFI
VNh8gymGtVFGFSj3jJXe3jS621Pgcx+kaTXf2BFJoOOKFIgn4ar3TeTaK5pK90r+1qVWgHFupVOk
lP+hfv/mjJIuSyu4BbbXRrA39qnLY3VW+Us1WV/diBicZrDe7bF3TymGtFcOHi34naJXMPFFwrQQ
AFOeQ2JCBDEreB7VKoiNLpuwimJRf47TXZ6w2kMYwEcCAHhB2i+Q8Z6svmvYZVgRB0tiR21g+MvT
Rl8N/uLyEZ3QbSaTHFrdYi30vu6zea2U6ubq6TsDn8xqVO4XzfZimIbyHUcGBMNaUrhxyE3nPAug
W/SqHIAzwT2nmPs6vx3lpXdyd18MpQSGBnBMCEdkaZfJvcKBKrV4PGXthTQncoSiqiu0yRIt2CCM
3v1YjfToUvUpOmwIJLxEr/WBcLz/JCoiCMskVsct47y5EWmn1LLFWzKC83ctSNh1Eqzw9bLEu9R6
qdX73FYZx1h8juXUTYlRyoD/1isWfvd0UqkDCmQV4zBRkHUwU2DXdfuBsNY7q4ZadX49EvN6YLx/
OKk85NxPoJa8lgTcSSe97rL02JuQvYOhY9Iwu+w6eIZ4axFIHXjqEuHyXvokpjHBbeqJ9rE4sods
DtqTkycclC7CQNuGbiaI3msFLq2XkrS2ykbVH+pC8OGdW5Gvs+WhI3jc9me7VUcbtOowODgwFGLw
dicTcSsE5nTlTLUUiYDzWVdQzbpztZhKlLav0ql0P1h2Bc/xY5uu2uvh//z2mpu6nPDClCSMLb22
s4depWV2X2GMg4xUzlTNTxhrMNtjXQmfrMNWBjTEe7aSjQ/iauzcZYWIWbgrf4hwu270o5IAQ0rK
u4nwpEGx6gFDf8M0f0GK++dIY0qLzvkkIhouhO9xyrauLAwnjyG7us19KEzS348SF89aod6rI8lU
+HNyTcygCbyGuo+hfEtT5bEgsttIUZNdiI7tXuBuNEgRUDuQYQcp6h3otz+UXql5v1JpY8uohFRw
UO3l5kPIkV2apTiCOaQPz6G7grfGcuAS9MTjKg0oVKc3QDaN63tRfFIY6Mv9gHE4j5aw8PKhZ2LH
xrrtbykpXouN/OhfkTDAjgB0Ql9iE0UuPVFrPjqR9wuF3Oo2pG2XG1f1I/luhByJF4t3nRp2f9W9
kbIoovxKXXeltNXx9E6FFzkFqXAEmhNgzEdPHnDg/TPy1zHGug60hBw2L56Lvqx0ycybvW/5bP2S
DYa2Qd1PrFYscJSMKk2bnoGjnu1apd1C6vzGN+KTAmZHyqOlOyulvHLHjSbEbhz1QT08g+O9ntiN
xGJBBskOeIvkCy3IzSGWMlKpO6Ur49mp/NSx65+B6TwO9uLtq6he+Wd/Xwpz3VrWv3i1ICr9zldZ
kpLTVW1rSt/tYSuYGoMQCTugksZfbXkyvJotyCAYC5dx5TPHHI3r5l0fopfDWA42zVVwPBuLz8Gv
AhEx4t4ln3cCdwQnZedxn0S+LzgCCLMke1NTDEsYOTEFQFxvD8sWPoPi6Bjrer1XfLCAryS6+dPc
oLBw9wqJYmKuwYGePkX7QyMDF0RoTHgh/xlNgSQrucwBum0jam7cnOaFt5iobnRwCmrMEbWF8x4k
oF+JIB/MczgkezFWrEf4YKbnfIp16S7obPrWB+CWF11HEjQEc6PJMIyE2JNp2pJIQj7WargY/0SZ
j6r4efWGO6stXSTqXsNSRcW+vNWiR9FcF1dzijE3H0lc3A2mVGlV/mQ9/rlZR9gmcqjMUhrhkpTp
CKXV4dKq6TcNysppeP83MSiPfEu59rmMZlp5ESdlKMLvd4uLv5zz9jRzZjtLBRL0EtqBCNUnZGd4
2DiQPcX2YMYLOJeWVBd6t5Pd532ztObyS+6HN5STUeEps7FDaVkng1yo/1pfN271OFVKiourqffR
i8qjMEjx63h6VMO1lWciXWiDiRMc2I0wfYFuTqSCOKS0pT9G/79ThC9V3N4i2EH1M6w34kruiM3Y
XzDiRomdFRkZmfgYIb5J6a+Vg79BsmPuAupkK0svorm4ygSubfUgegr/qTuHzlPOokbuBnY3Kbp+
cuspB+426LW720up7YoJe+5U0dbW14RS2JcyyIxrJ/n9ETo3FrEUN823vHzWJ7DRwsV3mN8cDTyo
Dv7TNzRm8h4c7OXyE7v8ATcUKjyrbY/d6ga9tvx2NTWlIbi0ANAKvbVRAe0hM9U1kVzyazvSYILt
Q/Nj7LsxxDlflqF8xuElwK/6JVMRDHptbURIHbQGRhXZH5vEbSUfzbwd8kOyup85AUfpc+ecNjr7
Cx4M6PBe+VpTnnsZLqavmQ2xgwZbM5pnygXK14OZP7buwsEFaiNK+dYemyQiEn1MtK0AeQCcloai
N0tlPYinkW6U3urfzfJ+2DwEVRpW5mS5WFozBnHkYSelUDuFQc+21twHo8zaYs+tjLW8BLDsWbM2
/AKjODgDLDquYVbbo3F6Vlhb0tV4vk9fgt85B38geTnA9zOAghkypLiCLNuvPBUG/zKQZBpTu/Bn
hU8bxr0aDOHMF3454TJ6HA9GvSGNOSINyPoCU2D38/pQiqLTFYC6Y3bljN6dtKWPlC1FRbPs8lf+
q1/r4gMWAfoRDFh61jJ1GbYDmRQTk6wPUY8asxTs1ASVhvv78MweQvUaBZyFhN09bTCQsg/H8J8C
x8KhqUm9W6R/Jia0UcqAXGvXIVZI3hfgqhOLyaq1+qWsXudurtapAk9JMVA0j4SxiZegrfy91M9w
HHz+3D1RmdqV0r04LQif56U6N6pzaKwfrjXlCNKnHoMn0R71TUpNI/Btr5IVqJPuIdFE+oROynAh
2WZbKOwBg5jQBPgLQn/85Bgs85RMozSd7EuM7DtC6GJhIZ3p7s54L7SatuQ9bvUDQBFaYcIvJ84k
r4JwoDe/jLyP4MG7WDaPuaq2BuVvxnIhhVoaEu1WWT04Kqq7dWL5+vl2aJrQ59X8wYsypggT7UUT
UhQwU7s79W+ynSqM3lOMRM1TX/UTItfhj+ZLrlXIy8QIUOFDcdZ4rCtHBy7zhFXr0YYmXysgW3wm
Q0G6b7aXcSdJ0aoC0OAdFLtVG7yTk7LyXnAf/65Q3W9X2yaoPpOIvTtoc0gCeOTUGZn75RMNbJ6l
zG3bZUGWG/rJRUaKdxQqPBzUcuU5/dMRnlid3QxaX3PKbS2O9c4OOL23hf6c0VRtsZ1AycAXl4YQ
NxXuyHRQzgONMqU0Eg0YDvpV4m4+rX3CTxBmfUpT4zvpgOc+iFETNacUA5kMvObiyxdVO2/xeWdO
p0b46vDwm2L9oRh2gOzM1hrq6F1C3rxYwfRDvCIjic326V6kuq/imnW5nJJTKf/vA1o7ck2J2kSk
Gejz/2N8mQS5CGqfP/wTUOSBaLaUpKgjLGmpi1Cx1peCe+0IVEDK2rhVdIQdB4CNov8I+S0bDn4J
4KzAJJU+WJeSrrcUY5bGtQ8ICUmbVEH++Opw/V1Vn/JkclypPHEr0UPbQ8cKMxBhC49Gm0X/23a0
oRSvg7SA+DTdKKYIft+PG9xVSbShyuwDrUpShPXV97VAQqqNx3nA0C86t3hHs4XaMtNfxagO/AqR
ExH0HDfqzPUMf02PS0Mglg4joLN5NNut7O+bCBgdmbqZrsk1IvPzxvXDr/6cF9oZXO1rEW4Tgc7I
rkwhxjcMT/rZvc6HCvdGdkoamzYXR/na7TrxEAzfvSEvQwYLaDHVw/HpVrZ1svjakt8AhrkAaYNZ
KM7Iar0vo9/Qd9lIw7PJmybeJXdO+XD3s51/ctHcBalrrnxrQ1RB/3vEnA6nkWYBvg6SFG1yy8vH
p3mDQQCxr64UwZPfaoQxHD5e7eGTwHu7ddYczzYo3uZyI/fj0G83ZvMGHVtYAH0fRnsafvUe9wGX
GdOOaa831vG2VOVoVAckutYRxNDrVay2y06q2zkRe2fbNV+He8wSHBOViNMGJ1ME+V2ZS4j9wlNi
/staSNg7hRCe7Y2GeDTWdS+srvBLbsQahfwABl/g4VKSnkEG1+I49k3YwSR497nkvT4KScwQTVfo
+e0okFdjO6Wc2tFFaEi3aPnG3rfmAIEFf12pw+oVHrPb0BsL0R5i725FXFDLiambBL7L01Fe8xaN
/zWgLi75RfhbS118gsP4sq1x/+NHhYhGs53BBLLFE9KyWt4gCUHDCKptrQYFF7r3SeRqqJSqj5lp
Rbd2NduBAxoGP20oaNCAruUkp/Ul/U/9FBvBkQGE/vvNZdLrteyEqwa5g5cJyZVOBvP4xX6UAuSP
ZVJ+0exzanybnkDRt841qyRKVcUdoVOMgmkBkSQg+Rt5AgpVv1/4BLBKhlD9cMkepukNqRpys3CY
sSpzDHIhZg1mZHMdCAGNfzXTWJqqhZ6Hw52VTxmkfuyQUzPiaUti8RZNUhWKN2KV6BQnr7cWhwmK
CORPWHCIPwCW0L4AmegNrD3xDh2omyj49rPHOT04FXa+aKeDLmiZVfcP13MAI511/WnlZbY5MpEY
jtua0zHqU/Rj1GGtnN8u5visg3/dY4oJyAezyjwVcpGFt/h6EE5rQBPsGsoVsKaIwgpq6sDoGFUh
ktyBxtGRjJmIEgZTaauZTwoEAfyWu0IzPFkqpt07MnJByXR4EVtFcaC0bSTWkEbZb03AA7IMaSxA
D9Ep+QlXKyyEprpwggtq0Ji6iuhZWIJHCmhcwU0dHWAsmvbVCxPeNPlGjUelJZEI9OlFfLuznLW4
TXp0zN/PjbvDGPnvaAwlHB4MbO4ECriOnLhM81wgRlKpk2+8dnMvC3If78XhFtNVAp93GZfNcaT5
2HBXSz57DobQurkAXaLgscCoQOhRx3J/+iKBMs2np8lxu99gNIQfSRn7Cf6jbMAK0oEMmQzh6uxQ
GNnXzwvMshh0UVVyuNJODoZ3lc/BJ/kOswgg7NnVCySrQmfAik4gJWqqN7khAhxf4r3focMQP3K/
epNy4EDkGYaqOv6cFAFucIWpe0pRbSNgvRwDGN3AVM4Qggbvu/zhS6tqvsvxKEzkGfPK9jhrK43z
Y3ralxBRNJ5bt3dPNW/dkAgTlTVsKtc6h135dCt9QtGZ27V8iQOc2deNv5GwyAWwVyM3WGAEZckn
b6oDrorTsNoP+lZooKFeZoBzwpcsLmmT2lQuK5QhWdq5X0meT1gSTtvo1VOsIlVDtmhPEjhEULMC
I8Tw+qdSySLX4sY7zZ8xXqg1oydzvz0iVOqnPmnYIqmIXxIjdA+NxaYv7ocaD9QVRABiWu1cTQJe
cS3NlDoJZ7oWy7YwPjl/MKlrQbpFg26s/zMbRajd8cQhwMIayGmOOxPJb/bL2+kKUBrtB401XMxG
l9K8Y3IT2mJn04XEL54eZk7rvNJP3krs8p7B76gPfQXlFNZTwDgXeFXFmFnDq8Eml2fJ+d3ielRJ
jyK3Mch3rGwFSx+mRE73YulowmUmVnHXY3fqkJo+Y883xoOpXT7CjNy6mo7AVp+cd4z7+u6GIrda
QTkvCe19622q+2bnYgqdnmbJMAPZYHCcGqaBMy1VQAlUXO1mnst0mLDTd6AfHU65sT7xBqTdpI9F
Cf601S+ZkQYwFrDMFLMDryRG8Etm0dyqflhBNl/L+xV39D5yX4CTLjH8oGEunqVyXXYS4gDowedA
bwAJV1g048a17bbc3eYEwxlH+R1ocreR5G7eFsUtRSmOaAnTO5kVDjpfKe/Cy0RTgwZIfWJDUnr8
cwQLsO4i34OBCil0ZFITORpM1OxtINC+jOzh8O9z3v8ibtonR5v2Re3PL+QKsNrUv0t5hfwiGGih
4MLnM6fX7Lq04zm6rXC+H8i3KI/sOEl1Fj83Tn75DwmlWtbZiGSNEc0PlxZa/ymlXpG+g4L0fJbH
egZfWPlW525MBKdVxGvPqEkI3IB882siw5AkWSHVeLB5t1Q6NcD1n9/hv0EeFDyccQjIyXPLpIex
hy3P2fjWxMPxoIOu2UpAnFuX1It2QHRCxxMbRBwaky2NvaPEf4DPkROJBYvGrg+Q4sx8NzwRl+ay
+R/CkmmNH39WXcZFouvAd8m8Y2mdStbcB8nGZ4Oz/w/pO7yxJdESqC0aougGlMdel6D58Wme5V8X
Qt66yJejL5Wien2YJwDdYAMhgOssVAg/hSdyBqVI4zK3BGf0Ntm+Hcx5WPQHhfe2Nh0MIJCdfQtY
9zP3HiDEDr77qShby7VdMBwfm+Vs1EGfr9ZnFG60JK28HiNJ3YwaYmiLN7bG23GUQcGYneLeGjYL
LTBimlyxXRikCcbJmSAvOEv027mDm69+6Fln2DUj2ucrJc6kjFOkqI3qdK2gQF6DXh207ENycDuu
RD15oa5TIV7Dg0cveL6P1YFmTmHvfPW3qBXyRn1WKaXwxaVpxAlUQWtI0y0bdSxz2mcOi2SeTGox
idA2rr5qA2rSECcfu1O/gyYNGP2jB2BUzzwUJDS8euK5WVRbK1LSoUDUgLqLFVUQbpFdA1S5B8QJ
5guV72dVnqg15esZCxTdfEhBbzEf8bma05bfEYLytihYJ5Vng/OaV6Lhdxw2ZwPo+W8/Zc938ALP
xneS2bnw849WMUMsKI+wbtNhcG4BFns6I3KS7HsuVuh3xMXrmWb1K62uAylmTTHjGHCkbz8wTAKC
g7WQf0BxWM1bcjIIc0vQ+Uoo6wOaetiKgMuiJkeTon9tjCXChBXGwsJVc2IqdcnL6Y3K6+RPSHS8
/QFoH25ylVUJ7I9wJ1SQIv/4BugvAYjg1zHQOOhZVKBHDx9aj/HgOtlvTDsaZFx2dzh3GyuRWjEf
U6febuavYzCrF9HE3eO7vUZ6Eu0PXJQ1cz5iYkzSQMXQxO6XnIh9IVcfwRPcj3CAVXI7h0qemUOe
sI0nKMeABsZxTTVcHxJaXxVJbturDCEO0o/ZP62WcR/N4moH45nSv568KXMfgLhB26GKbzyOc1Np
WZWXD4sxfwVooBVgyGdA3RUU2qGw6udsFkvsbtN3D7I4gcQ3rP8kUiPRJOfQHEMmjg6JmI4s+atC
rHM63d5C6lO/iqj5VG5q/YLEXej3vgu9F+FnrdbYUStTe3V25P7qQzyq9rGV/7fIEdmwwNAdqmF9
oovdo+vy8UXmxmFLVTZa0VyS5thR2tJ/1wV3NxWbYMiqGzyIg54YZT8y3AzYMz9Io//akjWKLHLg
dPRFxEjGSMZCslgjOaQqyKDyjuDpyTAbdWoDMHUqvj0WbyJZoWsGcfeseKxQ1oKLXf6lTDDQSbZP
20KGYonjWsSDBF63kFOVJdOlYiceayggEyWf9lhQv/nPFyR1GtC3ko+L8iaIqt0O4kQjKkyUldWI
y9/UhejUV22rWDZY2uN2a9ojalwDFuBK/ok3P3uoj3F8T26wcqDRS9Ge3JeVPk5l1ItODCzfLYx4
pBe2dYwYtz6HEVs3dbrTZpIIC8NLO1Z6j/haPMOQ9/rIC0/I+D2fY5+4dIRfr/q9aiZQEeAr/FwP
1eRLpqM6zcYlgXq00RNHwxBz98rEh8222Jx0B9G1Srq2giMuwrQkLqibIZk5N+Hf53L5m5TWml8/
fTOD2FA6UyW2U4M/9RJj4ycCcZyiMc596mg5Q9/G6TvioNdjREXALyWYZvobMO41XlFwhbFvbd2E
konanzrU3FYNAy/sLL49BK1uPtcxlufEmaP/0Bpi5TBco6o03Wul+v8Dn1BB3dEd0p7/KFRHSZ8G
t0HCGeeOiB7nB4bf0g3yKzB6CvQmWRIyMv8X5YAmZN2rWmz1SrYLlwD2FqLQrVE5F+qOlIDv31sA
iNLm2hmvhq9nH3Esz8W/5WTfOG8QQ9i3MIMryRQLQ9Ypc/jxpNTeP6fPVypYIXE63Du/e4KdtOhL
by8UOPWQV5Nx4S/su4vZtnpt8Ga5tr/V3pXwkWpZP9gW1RuExBQNFFjMXZLqJ/hUpG9Ls9sfxQIh
f4xAnliuyr9U26PVDj75yrcrFr+Wn0ycmF0JAczDD4RwB8XMZOX3KLqiHtHpJPIMWQUxSzACFO6l
ITWVOz1myVS+Fa+NVGV7tM7haoyeuOkjaDEb1CKTPDfgisWVVf2THlstuEXwTsmJ17Qv76LieqyZ
aedh8RsfPoKioGuCYP1YQQZlu/7wa51HPtIwwTBxCsnFjjmMenq1N6K/DiNUNgmLu41UUWwnj9xn
UNCVOEeV3z5O9dMGcnxs1KK31RGnI96Q3geYhD/zDkvV/LWF3/c8Lxv0lobKHMxm3A70JPgDKAti
apvYBYLmB+TkLq4mEqVD8IvKK1bYYuGkS9M2C4f338Uwfo+hRkBJgyeRBU/0ISvdjlnihL8UBrh6
jsDvhZkEIh8DT3nbEt9GClsAqsfrf7sk9hQaophi+NucHz4lr0bK3698TbeYqVoSVDrx+tVnFBWW
x6FU8Ez4FuVYWdI6wH1SAU2ANxb2lJbJ7uhMyaFtxXX+cE/2zyKSCg1XowqFdpQ06gwC/5nHuTXc
CmLwgAZWJogPLBDNZ1xi9EJJT85JgHI1mreyurxhxOhR6H1MtBOBXq9T78hc70BwVRPXedGxTqMW
uzbbQZQQCMMpSQ7Cb4saLG58qfTWElQMlt+qacb5sQo8LLeecXRFJ+U6RGZkdJlW8Y25CTA4Y2MU
inzG+Kou9DzlKxi07rzCxyb/yjlHggy0SRO/dIwYfG72YLz/Znje6Y++33g3NVt+afTtPS0lsYXp
eqiCXnEfFynqahSo/9MlDjvbGWeZqAY7ULmclkVWPtR6c/rOYT9aorq5g00R/J+rdcvEqtWuBl6F
10nYhtLdc1CpZgPdYSu4Pn98VgmZYSPovuiSBquiMPnX9HfOezo8QocZgkJWEm0tZG9yuYFDHdWz
uMu4H1Ovj3meLpW9HJYMTrm5BS18UHYV2yAkw2VCRHs7XcpvTvu7M0IPr6PD1QdRfN/WgF6xdqJ4
FS+QM0SoloEJRrhYHp0ezZ7ZR40xIKewYyfq4aofgfmKCmvF0LhDVDLlMwUECxHxRaK1WvX18UmN
EhE/eL0wKKWlXgQPOGVpzNSqPZ7R8WgdNI9Py0/ZE+n9tZi3bHuJWmGZ7xd5QcvOs88bu09LYheH
5LWoiGkfKtFBBgMwc/u3B2ms23COUNFc7RlrcG7gZFENmT1y6Wux5xwYngbtcrWhcQDNPmaXzMs4
zWIbaD/06hLP+RWEM92Ywpz08XrRuJv7u34hcFLS8qZfBO2Jshu8KPuBesVPiccEwvUJP45yxMxn
j9kCkdaVsm/7Tf4EP3f6iDXRvkdAF+fPHsNQAfPookmMw9gH4Y8jx7v/p+EPmXMRyqe7+W7bQ+Jy
cJXbvhdhMHsVl0bbGpDm0BZR3TJINEb94ETBJ7GMHSogxol7Ho88Em4rH5D89P2cdB651p3HCiSQ
aByS13Ci0hiiaKGIdIiQxWPX14cXp/9Keu4pNWiBY9ezUtYYy7iSmyJntHsZzAocoJQ1eReQcgM2
q1tqEznu5LJaLogM8WV5eHnQyd0khFaENmb0wC1ZkxcM8nJzwUhXpWUhI1CebZKe/K7WKVSzabDj
dRgiU7r+Bl+BFMZHCtBsT/dxN47+4wn5WCSuACr4nac59xkXQWcWFIOTEWk98/WiAwM8+QYOcNhe
jGEslxRF53gucAapauTLYSUWdlXc1AILgyPs+gqSipOCX4dBNUzYxIlR8lrevrw+xWacL51QuZUo
1ZKEscxB50K58iJLsfrk5oEUhFoRzIJV8t93I7XG70/nOBHZFEXscdOS/mb0sMI00I+exXTKV5Mm
cqKfklBcd2ci6KfFnsY88rPT7P53wBnOrCLaXglq0nGryva2B0XuO1xypxkAW21raZ6KA2+SflwA
xZ8Y3rgSx1gvumdMcgrBrPtpMkOE/c0iG4W9IcVe8pCA2ea8+ghSzKXC/WRd2Kft+WQU0dTRN8kz
K82kz8Al2QhUsBXtwrk2q7jtMLFmq4EzWqENIYkFfDZeopgqpSk+Joq2EcSugrE52BGD5m0tY9TH
/zfEL02l2PFIvj8l8FAvBzETZ48Wty6waorCPCTGELXYmLTaLss7lTNd/OK5jeszshZ3zn1DyB4L
CwYuMb5m7Mk24s9E8BXeZBhZBS4nMhKvMBm2CYRVJ4e8ROIpjhaZciAepDaalbLnoOgId8N/q6Mp
nCTNAa6aLSYS3gqcG7eFtndQx7bVWsvG6bkG51cfWZ7LFLCHvt8fP50Kiwa5xfRZ1TaG10jvehPi
tV+mQ9qUHiQpBwc7rtPfJIDTb97whe32jCnY3YcRpVsKsdAUE2KbjKPo2Rw6WRYF15lGYFLtMWxt
f3ypOkZjOV19/pCt2zoP67Qo0ZBFRHAhe0tD1M+3a2gU8PRtI9d05OLyJKKyVP52sqMWVJYr0nrp
IhgukiHRVLuWUpKTepjY4dQL6yEP+iLl2dgS/UsVlBOaGRTyJEGnugSv+tTwFUFMpmLo74/Kw9eV
w1KAquEY7NzFq6U03PYfF4D1nfoZUMwbZx+BRj78zvGYbh8Py7VX/ACSdgyfLIxJc+9KJ5aKa0Mv
JqP+QharyHMa16bbmlkkz870uCgD0gDncM/aJk62NQE//1+Kq0zOFOzvtBkz2eLwug5AV4r+IcCN
EtKcavrGIWcAN9sbFxZknof785+iGYpZUAv/PHv1AV6Q0ZHtK0vl8YdxY/XFXABajQoEd44v98Qs
Gk2B/OVVO48tmCIxiotnnRcbdriAcDLn7FQKfZMUB5ctwgYtgYDqnQMTLtIpF5HJN0spEonLLG3e
5oahIT28yk+n/rKePXLz+dLNhjIYIVCCcGxd+WEndeQ171Iy1wnNbm5FW1CB/gL8JOZ7gfgWHuZd
TnH+m/eRUmWoQl3Xx0LwLePl1PPTpVhVnTsi9vOMqVUmliZP3n+eyGuUGeiapPi+oBsqwA08IUvL
xVVUPwY/XPDtQ4hvYWIT4AZaEcn8b7Wv4gLhI3DH2MHY8aa9KAAq0y5BR0vReiTVXAo38LDHiWJr
KteFx+fHMwi+RjUmlSqfPqkiTlTq8rKirZpe7pWa6Ad6Vn+89cdRCutA+UpCqQbzG1bXw8udpYDU
X+q+svuPMLp8orGS3uuYEkvHyytgD2Ib199hhg5LxVhSsd5mjURmmJIqrzomhZB+czC+JtxM/E5b
X3KmLmQN3v7sEMPEBJP3/GHvqm1yBAZarAqKQ4OJPrzOpigxx2GSH7aQZipHEfDmy/oAEEO9BDGU
Z4Olpqa/pR4x7yrsciKpXrSrOjb9l5VpR0vm4i4rlYo8FCN49a4sio1oXFDkcdceADEfp3V7k15o
oBnvaqkgGFzWS1W/zAH0OgV9BemL01Z+oa57TILLx2udQO1tZqjnPK9iqbmrICCeL2f3b67E9fsL
8B8AtNL+naIQ3/PtdnirQyRRzhSgDVCHCKJMiB6Hsa3FTTzosG3RroGZMPkaIHSQqhKkBOwOUT/k
LAMeLvDoh7SN9MmqyTlSDvzIMzkcgH6iQhUZGkLp4j3dTVMskX2b4B2vUxfx9B98FDkIphZcdxKR
LUeNvD1hRY24iuC1gxl+LqeS0bjP/uSyxm34sIzZb13ZXWXIOv1/2SxZ70ODAbWX78Xrh0vkYQld
7DqqdS+bFAACZVdOf+6Ya2gaw1cf856DhpC8ZZ9AAToQ39a1klYI4mfhSWUY1L1TQZg67xH5P1G3
GS9o5ISPTzHmKbnNwADlIv5+uyzUS3LluM4zwMSPp7VuNRHNdGB+k9XzvrRG5dGKcV6Xyp3PrRPX
Hn3tIvvWEEDH/XXwZ3AWqjpMsRBiOvuHHaWUm37VoacBUCQ1d1VOVXnYIgZ0PCowwDkQNPHA1+AQ
QV5er4/Dpb9bUWfesGNASvAPqSYsWwndJK2H1Mp9OJGI5lXMlnuNn0eoIgr2Z4CJhhNQ0bJuRI9i
K9pgWWhyfC0vregOQibb7MA/WGNdp0XRC7VmOu2w7SqSwQRMwf3nCxVZPPrbEZbGB3l+OHVOp8JP
IMCktxlrQs1GRD7TsZGow+XKHGwlRW/H6YXOx5HrOqwVwdqxlPlSt9xpthlknxykHEuKLWZrLIcI
UJ6ERFyzhQbb1VFWmxIuRzCbmti4cQ1VJioyFsmnUdSHZJ3GmOmvnaDKg+kgivOxMRp+8SF7Fo6t
GKcw7Kxx6YBCyy1b0QpZn1g2kUuSU4PX2GEzCTn3w02CpfYW93FbiJnDMuc13CQ526h9sFZqF8NW
9x0sJixRSfgiYEKxSs0HwQRziyMTNRkNZZA+3FoO/PjLzhKigkRExV8BG/M8Gj6B6pIlLdUUGDw7
cftEqCAQYqXeJoKMMFA0Xx/13nmbUNtfLKMsZabswlwZ75ypp3aktjo/9KEqc85cpQ1Njq5no2TT
FYQ7hkn36+3ypBRslV41U93w/7gcZWQzEt//oREfFnMmnzW3vW+eo2UPIejqONDRcwKi227K+0fE
iwUdTyLFp3APmMgSV8EYGuWlUY7iRLmvFBNXg83lk3E28ttpHdFQcUOiDQvbIBGNPWNi+PUwWWG9
cMEaoL255KmUTkFKF6t8fXGZl3L50GGDctl4gqjsvTtgQb358DIeYekvtYreOOoA6D9A3hHTI2b7
bS7nhCs48SszSDtXiHQDFv0pMob55Y6L+GQsNiMa/v6ObBYZaw3izKf4nI3JvDN2rXFvYBIK8M0c
+fIWD4ffVmGdw5YYNHFpShOXlYVY02rzuOCaGlKd/KntF8mm3C6cfhx+DDtApdlxCZEwOl1nUlZN
cBEoHDzr+f1lIZ7HAh7x8T/z7sSWjkeW4H+s1cuRXg5BQ9AXwYmlS0AdhCCsB9AkSOTrI+EqVxCI
kOrh5LhUCzS20ZCiVybR57W5FJLqxsgvLc5Vpwr8asEM6dkGSt/asXBwU4qVKSWZoPrVALfyJt1/
s9D/NrHbUDHAxVreH8EtWedf5gUziqH8opqtBzKQZKOrXZDN9wDF41gQ+yr7xVrbHkzzR5u2UORu
JopzVWoB5AAXi5YTPCokHMbvdtoW5Ic7uEbAWGs3OYf+zaaiaBkk5G2loGPdWln5iwNX8+v5+V6k
A+O/4iZqlmGRNlRIFxO86UjaPd1s3epLO0HF2L9ymIhr6BEFAnGSn+5xmeDlxaICPTUyW7Svt2UN
fjI3PVItV/xFst4regH7ta/SO0xPDBd9x9Exwj+bzi1N/j+hK9xmem6he3jquujpvkusNLIZxpcF
yyIEsRuvH5LNIOveDqhoE6llwuTG2L2XssInxIZS/wlDYKp80D2OXWtBVvyJJILfkstNcy7wcWAY
e5uVX8JJCXsaTr07EcYaFV76GE98dgCTmc9xEjnTJ0Cff1IdPmKF4qmCMdd/1WXQ6NIqYVvjQhtp
Yp6/u39wKabVMpreMy8bDRpULNJtzuAv/I8CtrFygutQhjh/azXiUZOt7i9UIw+XljPUUTglOU4U
6f33oTwo6eAmZkt+7qXI/uVd10p2YhvVZMmm0rdc2kcY0AM28Jbkk15X5y0IGOvLQ4UZ5CcHp6X5
yvYcY7TwfDz8/ZvqwJ3KumGcC75IJWnKqJt40u3rbKZmD5vHdnvKd7G1gJFtkVEAtDRAAP3UsUYX
QxsOYSZGl8sij9ChJhfW537SlKANbhFvdk1R1D0mmw09oVooofSI4NkIIqSQBwCs3spRom9eVkgc
Q2g/+O7Wsf6oOjoWDerm6f5JjW1QS13YL3iyLFSrMSTHNk1IjcB6TI6Dd9FPFmiVqvaZrAp9oWZh
8zJuFvgnykwA8y+U91IVgx+uS7cHJz/8FX45yFp/5ehD7O11/lKpS1gVKU2P0TpKrT0CZNRe/BdV
KcUufN537SFtXBsw2FtNP6PIIcKthRISnEVUreXmyuVnD8XWqAI5ysei9lYOLLP3rPV9OiMKOyoP
5WBXgMh5zDSIV0LjIpBeFacJFavjoZNPXgUEPuZvU7MRYp2NdJ6jhA4DEyLL4xkS3I+GzShdWpW4
P/hBZlX4hmcQTJAVX4SxQYoyBN5531CMnswVsLizwDUZ7fjm3zDh8YWC7juDshSogs5B3We3/Xcx
FBx3RZ2jOXc5z4C8vntcy7fheFyVnLCfDn24nXDET68ej7mXjDXB5r4W2FSqQ4rwRy73/6bvAobT
lccQps8pq3Oeg5IKtSzakeIYgVA12G0zAl68qijzBYBwVokIdVI6FKOCcYduKJ2Ss7wHY1MsvSwM
SlUAPc7mgkyeUr+mhBrMKx8pyaJu+o059RotXVFPJnmy4L974dB0IqDzU5XjMnEd1mCcVeCA+7ik
REqVJeMeAasvQJV7F7owyS7kZkMs1WgzpYm5/ms1eyHNiSl1I1WMvVoEYxymYSlXMyBDULpLFwM1
WwfvuolNHefrXqIlf99sJ4JkQaff4wqW6aQSwbVbtUYDkimepTUATC03RniFXnDmw6EJXvzKn6Jz
wGcrRmzvzElkjsm/T/LPfhLt7uEccFt3Lu7I2AnonibQpun0GNlk7w5SQ/db8IvRaOPnEHByVBze
B6+6tKqvvtG5FonQyXzSlrZGIEZeXp9sy9vTLNwh7uNl4CncsXsMPZ0aSpR4xkViDWw3wW/WYJun
+wUjK43+JdJa0gb+ymxr4ncE+VK89U+hIEBe8L3NqgBP6eMb+Giwoi7n1XHh7cflJbhHmZmKD6Jw
QtuRvuS/n4tPvB384tAW329PGxp1pVTC/6Hm+yqagWRxWZ9RyQ3n+gA0AQN6F7L8T8HgLNvQwBZx
ultnTya3a6dGi61zJo7fmijmVl1GsG/V4YVeTQL/QxU9KB1UV1BgrhC75P+JLAhWUyAdcEppr+So
7Fqozbv7kbJC5RgOk7XG9HZ2HJ6uDbI0cJ2C+8W/GlBtcW5wpaEvKjcw71fp2SvCqtZyd02RACtP
JbHoPMRXPtxGbuzX1VwkSqGM+ueul3wNAfdnlclSqy35obrWzp8sKY800s+VkvtoqH/99ctjgHcR
vk254arojTA+P9e3RmwXpMKF347096AhRFqyq9YIp47PbzWFU9yiq4bhVkjhgl5cX7Xd2+1uioXv
f0Oalf+JOwC2JTsw2UXM6lcqHy9u84TIin+q0GcbgK+1HCAM7snBqK360Lyzvar8H/o5/td5JZw5
Jf6aXqHDhQaVvIiyGSUJYpWs/bhNSEDgzH+Mdk0y1HbW3L6O9cGBXAlKlMPQXyNYku65zveCOysT
TVaICUbmbobkbpELY0oeTe4cft5Xvyt1K98sqWbpnQTxoZOwrx+4Tj9q2RO2HC9mR1tkSGWgoFYP
cWye0BU1gGEKsJYwM2NmzqvC+XMG4bzWYauLhZQ6SSVJuz61EdNpJILhCYdF+c2GMwfMVeGZuY6x
sAmbdhacmS/oDZDmKY5JKN57lTRJrJWWokqiClRSuJ0a1PFKuIdk0kfsXgHi7EM3ACtDZaxjDP0l
rGSlYiLnNTo8SUantu7ON1TvD9zBjJP9khqTFDsWMHR8jXPDawO8AffoctyBt4za6a5SUH0O+7AO
GbnIy221uq6IkqJQG1ooNf7NuWux/EZSacSJrV4vxpH1IBpnSfCeWovJNFzCqKM3LFu+98EWKdbw
huarfpKCisGWvzTmW6MgngBgWgX+Zqeyebkkggt6Xwis/lC9qxJfuQowzXCN7yXhlm9X195y1B+S
rF2mb16dcWXSSpf6ymkE8/b695ADhrFOMlFhfzggVyUaFfqc6X0pjXRVJ+h/dDTrX6Sc5dsYP6+w
BOkNcgRf+l38q27W+ZpG7sTSLruL3OLZzUQwJH2CjybhKV5CpDx1iP3Rc9vgD9Jd92fAZQLpWYE4
AbQIST0fBH41paEeDfCSO0OKIO3uuPY5M7tcOv7LEDkJ/54YMzphVCq6/fRknruWPpQnKJW8NagN
fZAUBL2PVjePK3wQGvvSzWiYfotoY96gUxNySWsqIJi/ADmBbMFSNtTn/Fmg0PIO1srATlNQz1aJ
ujTeCcVP5LapFT8neDwEK+pliiYqc3xm9MYfiKIZLHJLX3cmBUlTLnrAojI7eCpcHXA3csI9IlrY
MwAbQb3DOkLiPcu9IyLJU2ll3DBizJJgoO8Vleg2fp/SR0AD8K/g9hIq8zGzEpJ8CvouSKxkU+w+
deHsISmojpYMKGNRvfMZKQ8UmdL/B5H7HJ0NH73E/r3RG+RWFAUCQ+4k5i1qYUSLgoqAq3OIb90H
YNg9AJcusvrXBChuGQ1R5ToW2WUO9QqK7nfe3OzJBU8cX6fSfrWBXdGr1zU9EXaHdwR0y90pJ2fZ
22OoZjDTZ5gwbruMasbgWDs45s/ZJQg0WXIuIqEE1o181hb8JPVTiCLLaHwBsSHE3phzEuqFGfNA
7bDxGcYmC1zU/ouy6PzYI909OLoBIJ63TF4u74p9ze3VP2qd2So7ztVizPrYVyHadl6tN42Su7NH
mKkhjyG7KVGuZudNDsUVZz3s0SeK1ewKzjJxoyjIariNcjbxwtr7PUn2y+7T0QkwhGJtPjoErNOX
HfiO/W15Os0NxyOwlkH8+ImVWkQNFNazMyVdDb/OTUQFw0NE2qBVWXDoRkQhPz5zjWn0E5EHO1Sw
OmSl64OKVXwuCQjEwV84EMA7ZgoeNfILKS0K5okpxHkbsNmeco+arBaGmCFn0qgrNvD+qtUI3Rnv
Kon9CBhJ0Yvrq6JWMPbLiP/jNHPfIf1GYyM16aQ2GYd6BCsTbU/VuZDWdVxf00Cq8kBiMPU6B0jJ
MUJsaBv4gX3xexvMV1maQdMI5S3IWl6VtqFIeCUEau+GIDQbRXXJHB9aF6AhQdHDNNMex8qWCgV4
LMNSKvASadw7IJOb7Q4H/ltDtxp7rJrwO856pLW5ZEMTMcXVpVRaxXU1eRAYzJAPcFTgtiEy3UQT
bIfND72mskWWhnzMs3kx3D8ZTl0+fnJJpn2cb3uHefT/VDyf8CHPVfsJwhPsb7C6YJldzau9H0yC
LK1nT7+hBhqsZC8OjKUJHri88KvKKheVY6/08JuND46eL2TdakJ3foS3+lrUzi3HDP7RVxiTl5c3
jeRYpkdVCtDzBjjXVmU07wahiFti8lEjLOyTTGkJ1J4+OtMHmo3wW6EeQ6iw+WobaApFu/8+h7AK
BmICtMWgTDPignreo5ivtQd8QZQdiKiARcNn/Vnr6eGil5sC/Mh+UwQA8TYkFMOfOlczwydTcvyG
5UTgaa2oxgwgsAbDrzXPvDWX3/RPZ1LD/1wmFBtx9XY0I5RJHWYEllNG2zu8Xqsotzq1GsXWUVky
Ug2A9+vu32CaOJNV6fOoorVMVkXCjBEedivaBHQpesK28b6wWH0FI95igXuF+vbARIw2zTZ99OwR
dKNQdvv1jT9PKw+u/xK5835Tn/05m3lB6Ww4pnTDExhLxNLhm5zo1yDHk3YTmrRXYq/Xr9LaeA5E
jBguqhwsTDoapxKTafCT3kP/UNfds4QxBttI8GhOLfm5Vno/Vm9qSEZ5olAt1fyJt98MuJVa6acl
a53+DEC5b1I2BvAGxW4EOGbBYaivtFe26euyBx7itLJjJ59nY2FYZpP2ci0dnSCa2vuOanTDoW8q
Sf86u1WgPWqhI/OU2Xk2TCQivYhC3lnpPv3eiqfnjVaob1iFV9uvSyw+z2+oaVzZpb8FnuUuwjSj
uU8661OMiaDUhX5gzY9HyBzxrbn2A0Wu6St2U//YVT/5nB9al7ZK5YzJZOzLugAulktE3Y0+q+vC
8SeSEpH7e/sdABAmOSr7C1Dx+bf5AYIqAZVE4gvQ6BmMJfhbni/u7z57msgZFXJM5MjCwV1cE9Qz
ZAFZ5/FN/73XWPStOthujdpNgfdhpRLCjB/OR5zP4g8frvo2jqh5OcUUHF9zQFYkZaX59L7H43e6
HjJe0tXWDH3VuJsfSmBK3gLaBaaafGr7YdTCoab0TElE6/gPkFuEtUQEFJ/xoQnvdmJCq/RwmKi8
FDe5+UWsL8yIEX9GThb55deojtx+K0VJeWu7e3vCpuEu1YpjKiU4P+fckPVaByO7L+xUc3McExmm
gSDGprRKOyNtnN4D0UIz1cQeHAj8Gyit3FOtVOanp4LcnmNgO2QNCqr1j1b3TC6Aslsc0qa0UYZ5
ClNVb5YVBkcpUlLkhyUWmZqstgfkTsfKGw/SM22Dkma8NYrsUGv8ec4oC2jK6GkzrfFEkeL4vVzG
UEfU39hZF0EAgrteubZzEQ4rayarZ+cfsinOeRyzxodx6CBoLpoE46C5prGSArJWkawEUXbXbpPa
xie7yPyrCUYcAoIXlY4wHemUsuDUiEeD6/ucURqnkfhi/VMppNixj7HldyvS/0fv9P8xSM/fJvd/
lrvz1tKokAaQDtZqjjGBpXx6MTJ4Virb4Xz/AULwR6avSvkvPsknsNbX6hm8qI9rRX1/pulY3QNH
g3cL5b9lffvns/PktP/uqziANTzMu6vjL9SPiu0K3xXEGNK0xxY9All6oby39Pn2fN+d1LXMCHmY
t7X8eN9hclDBb8V0fl29BUsnHjUJcFLnZgb1FPTOGp9VebU+rvctOJNKopiJg1GVVM4urm7kaBS9
GEMS5XmfPGinzoe7xoCljPTl5sDS6UykIG+XKMFwbz8fRmHWPfBbGOXjXsyo/CTb/b1VZvIsmeCg
o/hsPELwiyzzkv5B2lsLNXfQgflACZ6gJ+bGzFtC3lSurMQbkNLlB8ZSxih4VQ+037nktAJPckFc
CkhfgDBxvTu+7nZWuCsfsFABo0aBdstoIbUB4nZbKzmtvYBXqGb1ajIk9dG8qAOGwTF7jxmclxqh
Ml2ZR/70a0KJd4BCIECFrih3wXEUc9/1Fh6n/MnYD4pjT6LWTd1DNeqYvGyKdzqWqG80uX2RsmAa
VzxeKKH0ya+n50OcvVJ551pcxBKZNVx1XKYl0H6Z6wQOyC1CVmA1vvQ+9T1ObQbFfgtFE0kKSxew
x7yeQ2P2wnQp3aiX3FYIBF6RSRu/LmYPFGdlCaKPz22R2tch2rVf63p9Mgea0A0xVhM2fc5HPAEP
nymDaDSN20JK84S2MHeA1nWdvjWi8F0CJ2cZeuANTflFWMZdZej2JpqR0AqnomiTL31Q110gKQdf
1/ok8E95YY9idAObNwcwgY9DjnPZiRzx5+AJgarZt5UHg/SAf72xxSA1AtkU+2LXhqQAIvG4E4JB
Hb5N+Aiaj81p9I4A3gg/YLNh+9ByV0KYonCnduQGR5NP0XyPCe1Fqp71OBV8hOnZtEabz/IhNum6
Md1ctzZj5icND2aRbhmWruwMSw4Eb6iebxX6lHclbCyMdwrRtSe3bxU3cb5A3+I0TaZRY2RnP97v
C3jOE/1RxF8zoGLIYvYHjyaNs1NkD769yR7odVRNWh/OsbXYjsUE1RHTU76rBlGc2bzEAnH7bTXX
c/YbKFb949ZHy2WsS78POfW6dm0ghqbbzwAUIuRhREJJaEDxG5oetGTWaTafhx4RzC3wVgm4J0Iz
jijntwUPQT8SYkZ2xPD7iPXOgY2ePFGbHy2h3xPGqj3GQaFOpRF7JeYX6+JVtW2OUjFsa0xsd8WL
DokudsIDD+3q5BHpKzJPUj8KJVl2trUH4wAARu5oBBIGS4HtQNqOSNbEB4d4j/2kyvoskaG1GuOK
x37worH2RA0evXwOPE4P0J0ACOthhEM5FZhjrwaupp1yucw6QLgRDyzitbSDnojIzJHHG/n0QVJs
qSlT3TjMbcrmxb5Q9c8Wpkhp2kF7K/DYg+eaEBAetUTMGXC+Q8xPUXu/9vlgygkK/Wnle0mWgFlG
rtmi7KKiOADfjxHlNQnzNLWfO+0yrfIFOhuR02xQwNstk2Zn+iOutPoBx6wLZ/AnP8fq/5HgMo0U
6mpfRGKo9F6azz95R9nrvBigMC3GcZm/VIP2b0wubQh4mZs3sCnGrNaW0hUttRq+Wq23KQeO6Pnw
jbx5RriouilM023n8rvmTHxjz3A2CazY7Ood8KmrK/tullYyYNBYXpWX6M9kmp8e8VgvkYq7U0wg
7KkPgAkBFS3So2YqVjYN4GYUqnMqcDfZ4xmfa2YTkiSJxQ3+y5Ny1tpeyST/LlgVBP8HvWgL/rF2
BA+WqVtEC4FdGtBeShHgvQHQyPYGYuNOmVG53pDNnIIzmhgqMj0I76jWXFZmlQ+jAcaK/g4IZ4aa
6BrW7iKtCIU0c1HH+l+OrYJntKBxu3A3TIKV/D1ubx1yHwP7lsG0z+LedNkmqrYMRP5mTdj/fkes
Nq4hqq71HnQrOU2cfFmhDQE+phBa2jBoo5xluaoGAT8F2dpC4mlXjAF8kb2GDnXfGHtgrK5x5VIW
lDKvtif8mOPZ7OYWTp1MoD9/AB9edGWtlBcmgHrkspy3dsTZIjgEJxvjkyyyP5QOkNG+U6iO4EeD
7QXEOnswYo0g9wgFaLgY/tcb/1kZ/PIigMJRiEdK/Tj0ZdB+LZugvU/yXyVbnn6WO/r/twO6eGo5
6VjNkK5G5+wXs9nRZP0tvgbvUQWfHOIMc9FQUdaZbiPmAQ8KY/qVhPcfxgmyQHkU71bH7Z2o3ju6
SUU+MyLWUNEwSoHKLMdEAppS5sfHze3AVyQMSo3Pn0UAtfFAP3m6W9ltksgOTWO+MvJugFid2jkW
JE7I2AjvfHmDQLXWnDSh+xOUxSuYALPfJgsr/u0nLXmeL2DU8krYG7K7G+BF6QfPAjlQrrVvyNWy
h9z/bl8cV3GfQRrxkCCuwg8HEuTQypBn6zQrFkeAtdG2s8Vr8+2RmHKAAI/mSV4f3LZ7pEFA91kK
iqOf4My8aplcmk0Jk+PLi4gvLaANkYNyw1XmDQSOwV7uNAdruuzYKvXE8PRjRhqguhBb82Jpmp1O
TfAqO7AnpmyOQMBS6I4I/TfFg+AiAaLEf5Brgysk+Ko2c4Z/Nm7FpQ2GsWHiCt7pPzjx4NVyJwN0
KA81eR0hLo+fzvajIGEPxgzBiK1irLozHxPjaUHPuUvFN7ZBa8raGus14Sm2ZS/oc3qGBKsGTB5s
4/W5m3e12Rjsff1Iejm8BtGt0BA4SaIVrlk+F8z+hYh5qglB0OITbXDwsDPgn1xlorWDU4+ycE1A
xCzxv56V9fcbI6TokjD2nUpGWqRU6bKaPiZuaMRgL59ezhV+T1qpeXWsbf3xNJDd2QJJvyr//BsM
oXex4686CYSQ0QjL1cx47FTnf2MwU+f7oxBKThJ3h0kL6b8uGNbLcDgiYyOKE+x1EJAYIHwjDN3r
3Vabj1jF1FCCo8bYAY/QE2tnt9wcGsaDzVaW9khSeQi3Y6SC+XFqlNdgGjxe90y1evtiPMTyiYFC
O+74+7US/ua0D3mX8T0XEZyUIGRNZsX4x9yhkH6sXM87VNAZ5sLHqmiudPjFW5vyN5f3/ZpCA8ss
gsPdzBW32axur4+ELLD+DIIog3iPJ5p7s/Qj979PjWlHWzCHR6gVDPGqUqVs5fPz8HYcGKXcBEXI
vhY+x02zj8EZEUOo4SDFkEMTUpw5bA90fEWGb/imN0u8SATk1s5dlstyoB867JMNDediTeiy7TbZ
R9rtQa7j0VrYmP457ehUeoEoJ3dmDHVAhzuzD9pDRRuKlDlXW4E4qn47SaoftxNG5G6qp0JziL+l
RFvdDZmYhKVRsaR2o+JxH55073aN6sH7rVa/GkbeOYsKrBsJfa8RU7o3s1Dk+8OchIRLDG4qe/ok
YFdGotF+vlhDhzJwrkUhj5XKSfe9fnHl0ACO1TobQo3sIQkFsBNjZXpl783at6z4227rHZ8W9QKu
28hrUx5RnKsyAsj+Hd/4Hxr6xy1U8rqyWk5vdXZ9WhDX9iWJ6CCdyZLIo904IGi+3+WN0rfcuAJC
aJ2w0Ptp92Rn2Azq2xkjYzdL1LFSfWtgJ4EkRHqtZa7YkGJBiJPhzBlYfPmxkzCKDy0VYq2GE7FD
6nFdFK745XlQmMAdEp1vaVoAnZAUkupdnQI9OnUqKH3mdE0qKiQ63Xki1XL8/SAzl1xhN/iI1DrD
FPPFYX4LzvEPvWc3ZN+bdcGVohTWXbVGLxZuAzK0kWJWqoPQjY8n+PxMIIii18w8mgsv6Ho656G8
iOcnMBoLtchulnp+CABEvsjJljVqHBL0fYgVTI4MrjIAHycccuE5ZH/Ud+/wQ7NfmVxboz0Yobi3
KQSi6HAFqC4/uJY2uwhbsFTrcJy4SUnia+082RI2AzbWpljqLC+JlhA+f5YLxU6n5J8YKGpv0gdJ
AUaij1QVZHY3Y4XhaFeMe6lqtX1ATm/WP8ejAVsPH08tqF+Arj/+iZzzIJfH6UBN/JrzbsVahXY5
CcjzIRADuoy8NPoXcZAoGyUtU9AM0Hi+wvtTvew/bQa3NzROZamma2oiTGAFdP5+2snvgAP2JIeK
mE5QsGtpjy1qyQwfX4XjsE11zgZ61qH3ctAySg1GAQcWJf/rKkr2z4vvSaDVGNetTx0aTo+16zt7
3wc3hVv2yclDI7u9B7J3OqWcSg4lhZkVqwkqoDU87LyPyDEY4F7rRTiawKtbNE9lIyn3OEnkMXwB
MFupfyuux3qUOdXrQZyKOxdkobPsEB+D9S4Z44Xfm9eNnIUDzYseIiaNQeXyI8EeXSDo11x5zJR1
Ggtbsb9P3ZSgmGRE9zkJmAzELHs0jtzgVuY1rr4Icoz35BHYVR0tFEb5re/h+papLduHGw11ndHE
9wRAwWxi4+TlVNgTh3uFuO0ppYZWBrc9qVTp9ZegdNwbX7g7tieYNh7fbOM/8uNF1gsWk2lXWim8
0ig+FvvgMa+v39PtjrTZInK4BuPVWc3tCtFd3nLSkQZr18y2QnFabVr1wsZkyNStnz2DXiFMplzc
yb0SIawxep6BJN9Lo2i83WdtMIWkA9h4Mo93MpkD5BRQ4AfMm/HM+TD1e5WSv2P5G7LSyN5e/LRh
JjrWbCHgu/lr5vfUnkgOwlHThK7JqBt3LCMRnW8FI8Sa97ichzhi2ZV18wbmgyHFMB+Zzqa9xlft
1HcNMcCyMy3WSa8FoYCt4ofGwYHNvoL9YcbtLwaddp8PbWu9WyVCzB/5Bu/1ntFJ/uxUyErj5Tty
9+xWl6pefOOodJ5dgDcRBG0TngksTwShthtb0RM2uAqdwZ+EFRsmXFOpDkiNVRkUfpFYgWirZcv3
AaplTsbJ9/9yCL726XN00+zPoOTOUNHeOll3SII/uhjpYoZFT57eyYmOfnyBjQ0s/Fr4RWVelS2t
edwFtnSOfdmbofYtAHBm7yg9PxSyIeLoWAB7mBA4ENs61ySCNa8cNZHPlfkQBXp0p95FABnDw4jo
nLPxeOWqRJWAybJK2blEVM2WOYM5dDLi6671pzchbq+l4agU9+PlXbrhRGhFDVkyH1jet0uFsltK
XnKalEKuoGjIK6iZnjwmSfP5MKau/JM0isvTRMnO5umFF+NNc0Rrn+o7QgjAtJT02vq1Lh57xOM+
tI+5FL/8eOX5WjFAv1VuYXlXBbPvtoK9teivnb8WfJZEkYBL4WQ+f23CZHGHm+9RppL5sCvvP5us
LXL7bsnM9BBCjR8f8Mx/N3s2gOtRikeYO3MAS3F3fMMdG/iSZpI8hvqz+v44/hvLcGXO1b4MgmEi
CzShqXufHzQGjdstJkTIxtbFJJnFP8l3KjT2l8nFsFCKQEzF1LVWHcxvR9ZHQKzMyqy+/SXtoo/X
gd5isdYQSCT4cIv0/xyhiyjVxW+RtCF1UGGTg6o9Tm46mTFgxesj3E6W0Y00W9th08KbhlW8jHOB
B7ltC5l4iT0wLwklOjhvt3iX/7H+1UbUajCV/ZzlgHLw0VKeFVnmgDq5NmbIHhg2BbF1JDaKLQFX
cDkNg3QUT+W7HobjQepe9kQcB06mfGMsE735R9bmtAmqkEfBeJXkCFi5KbS9li9dZPyiWpud6JnK
3FsCxgYWsPxXoi7VQDR+4C14ve7cyZEGVnQVnFgbXLt4Dyl/i8RhUFrIp0OKOn4YGzctgY5R7Oaq
WJOChzLxXzflV2kSGZQZVOwgXUECLELX67hklK2TiOANcwPaNLFqkcGXQqeJwu07U5IBX0GAdcOA
om3NyRv51AXm9FSDw2ZY8fs72OkYX+EZebj5LIUc7pEsS4vnNUkXRnGhg+J7FCUbyDEEDson4UAf
Bh6aSpOYoEhBp3l4oon3hnhAKFLqigeTmCsiVgMgHVLRC5isZRKDcMp2q+pq6wDONwI6t4LIYFZZ
X0ynFnKvR885zMOiebfsUNywRiy70m5ooDhj4m3fWF11xviBDKfyKeGH2OThfYEykL5cjzS2U9Cy
ljHaulSPSuNU+mLRePBf/nF2qcUCNIJIqINIHauY3T7WxgHh0mtxoBkg0px6kwKK14j7BAzV6OLz
n31g8ZY+DJ8I++0aWPIwOH+vATJ9BdkZ6NUlUXwkIRB+Rq2kUh4z0gaNJVSsAwTFjaSIbkLZVvra
8yhVxtmh4DqUKBDPl7IKL524xF5m1aiUOpUosA0xuROCAA2j/JIltHPmDVI5Z6UQdUfeUUUjtLEZ
+LX8LRGA8EoJkUATHFAaN59kxwV5HpLhwtkHjDGP32/hiO9PLuVj2PLZl4/lMQl+Pt5YOzk87tPL
jl3Fm4Tj6maZvsZHSxkH636z1iMUA3T+kCruAKogQAwuDV8Z0s5aEFsjmocd3UnJhj5BqsU9QsG6
6/YCUQerzyRipn/1arZHceKmDWXEA/C9bF2gJqNx+pW8B3w48FGOXjgJTa82EbtgQUz6fbuRda1z
vfQ+JMKKDrpLbZm0C0FM2t2y20eZByoCNMM36zY0PeWzTDuf2nU0nLXjuUMi2sPlTQgTHGBbYtlR
7E6BtGEoCeGaeU+kuoQ2iIZcmhx77otggpfZg5SdFj7cPjQevFbUX7TS1dqawN4KYWxXFBCZrSoc
sCRxHwXMvQ93x3ReMMhlNHyTUoKkGz/0YQz+iDDg7gkxjZiF4pcvPT2Wq40XfZ/HIikFbtpeC3E7
BctwpFK3OwyXK4QZM0EA4AU/8RAhBLnr5tp99JDxLylGbCXsRXxHZKnl9aVNVT7nHdoJ6T+4S9oh
NRhrj03hIUVQpgrtJSe6SsXxBA9cM5ZXVHk7Nom8cDJ7AbV5RGNrvF0/thr4Q8ax23otK7dwrIws
v9vzotZZiIUU2CjUdpp//EXXBrCjeTDdxhHzmrAg4jx5HjaSXeqXtq+wIymOX7QO4Wmkc57u825W
6MMP68rjuUWyPwqGKMIFfuPZrdlHAAGfkhOLXQ+LZlbNEZZS8oA33rZLb4h90qAkY3ZUKF8SjpyO
YBuaR9Wgv1r4QKmw3l14+pyddpD7fD6J/V4ALcbo8sjiDOCLI6qwQnZIgkZLqitakK+pUB2LRgJD
Bu0Ertzk0NwuRhRAi3U42YLU3Ta7/0OHTJ4JoivCcKJPZ2RXOxIDpAxsMSKeCfSGFEatai5OTQ0U
9gxWlMB9DvU7DLgNosxE85IY+bSuOmFIuYpJU27nh8ROmsqx8BEbFk2LtWPTVnOlPekl/s5JHtP7
zZiYwgLTyUl0ZBM6tWwK41SCgt7RAHM9CFxSa4NzxJQ/N2HVBIXF+qEPZNC4dKNBPjIrN2EAX+2w
OmHgW6Q6rYmB6NUqn2yzjkYMzg4flZj+hLxFqEDitUieM81SL3JhkU3Iu8zWHbCeupeXKupymUDi
UId60+anLcl+17G6D4DgXvxP4oEbngRZQmvYGzLN0+ONSZ+4KiFiQZklEnF+Sk7XMc2fYB9MUTAZ
5UioGa7GpBGaT8X4rHmz+gt0jlL9fetN8b249RJRRwz7bIlmyjZggI0+bduxR7VPIvDL/0eVUoeX
OCPLDN+kr7njquJ+r/u2s1XrOTWqJ8euL0YMHkw1X/T7d4G0iV8xei1IYawxKXdRmoKUFUy7LEsB
WzCG7BGlpI/YcxSNqCNBdbVFiZhloslPNkdERKhsL1pAy2SQ/xqQVHG9Io1CsXcexEp9ocY5h6EK
3p6Vb3YDRb5FDg4mv82oS7tY0YpRYadT2/s/IXOq4vyADI5dvwtvvw2dJBLq9bx4NuiJzfri58l9
wKe3I1RRqhfQOwP9ouD7p3ZA97PU9Xdr3gg30SRSliOtFa8N56xvTn/yUxp2v23+MWgp+E+f1BrP
nlHFoQM2FjzIfpB3lwRk9+ZMOysF0hIjijOtXZzTqcT3IFj+axCSDlJIr8/uzBhwlXeGpSwYBZtm
n+zpP8ij5acrlficrbePkcGqBwpBsuh4/G/1YqVDw+KqBd2N+D3AalU/DBuAzYDB2WJYpAKk90vD
g8FSDKSOtNywOoTl8q+RXJCHbviH3AoA0GGqdlvg05d87msLTER6T4taXue/khriiyxpwA3i8gNC
3ZkyTZRGa8PvmfRbo0IP3RcAb5oVgrM6W/l2n79uvi8KZBM8qRRSaBGQxs7AaHN//xLjao79kTMa
A3U09fHYXGlc5NNy4Yp4pbSrKcNoS3P57nGUDjAVI+Jym3PwWLOv2B1N221DMybwvPIlnuouweCb
H6aElg4c8ErtShUc0ZBzFzSkgaStcS4YORFnSfb5ehwlrMbji2HbwLVC15kbtmf6MMnrnIyoCB5o
emq/yoxu2H6YN7TJVzYf2jnH+y2PfAY+04eWds7jzzav4yvHPDo4Pj+JmB+hcPNRgYo+WqiroUNb
SlYEkObP+lRFoAlAoRpSun8cUyFaF5nU+t2HFlwFiYgUgyMvrqNYi3zTih6oJ7nKxZZnbWFAgZ/3
ghKahbgY6+nCc7Xfh8IqrwEvwWrZbT/f8tdaTzwztBerVdCPE+asFevBSqcq2RiqvTWSNBIbiUAK
UOvgtBItIUJ1nTzdlow9yGmJ0K16jT4Uuw8Fry3gC5JD6GUelA29ZfTim+QLUbFFSv/qGmW4XCt0
w4JzeF4vm6zo5kYd1WI5QX1KOGDXjMbbX2roOCkKuG7aC+oZXg69OnInNdNPnHlOKFLU7Zl1dkXv
5Hx4Lnp8FCrHX/x2ROK2vHsER+DoIpdOdJo+BHvgEjTiKP+sHIbsLF2LVHQ4z+5aL1ReeMwP2WEe
asiOtCpywxTViszIyaWxb3Rh4uBSIKLMo8dtGmpx9ANTlikrMfgAxNvlgBV1dNJqbwqsM+DDukGQ
654p8wjfUR9/yKEFMmznaZWFuzsglVZV1BT4x8FG40Z9vbBvPHmNlcnQxCuyILG40obd9I/67SpF
b9ETqBAL/uTCGzF+BTzcVmolxhlcjfMn5JvszkByG3I/zjNtF3cuREHtpWFTcuLR7MIioiHHYc7a
6dZR0369PaFAQQCp68Iq/VdCBEeSmSNefPV/h//miH9kVtUSZ820AgSlxE9tL/Nsg8zQUh+dXfmT
lONzWkxr4qsYshCpqG5UpzSxxoIM3i1pKRaYinmM6yyo4wXZw9zMYD/25uCA9hPB1+nP3uPPc8cu
phGj/7OmJZhbNKSmTy+xi2yQJ5Eck6O4YHgYoBv16dazUd984P2aa5kBZqKPW+g4CwWbg9NhqA1t
2oQ9ZXpUqzwY2K/EviI2jZ9TBf55AllKK1yYgWnCgf52P7jwhzQuLbpaoRiGkUsuUIfHvcIT1p8s
oVrhVPMMngl9dA6BKQAgWCS5R2WN+W/OUhO6agtXZITW63fUXd3A7unLfuW7sxA0LpzVwwQ70QN7
2tzqYkL62+/zLtHfRJyueZEBn9ilQgi31pNUkrUfJaWeLQiPoA98ECbbYnK63qUzIvwlzEeyb7+5
qY41W0UedalkJJYssagaVg3BM72utS1vWuDWcQ94zB+focL5U74fadHk1dsYdBpqKbPvWzVAZA62
WUZpqG6BXCBKxwWmYFKk6r/WREgotoNJgWMFng2YyzlBOlunYJc/E757xEKKUvfvlOMZhLbxhJlR
+x1liSCk2+JjoVSvz1etp4m8YV54ui5qyvl/UXcl81o9/9D21BqMB4lL4HkUiFv+66P4x3Rh+Ms2
ZzI9UYkjeRxRmq3q6oEVgmMRliF5mWNufSfw+7lMtHc8gMLnfVh9Zy/Mbq1HmTy9DZoQqUXUZVBt
z8hdYv6nXE1bIzonZeKJkfLE7nU1oLgt2jZF89HH/91F6PBvfT/AyE6u/zqbrpzSUieU/1RGvP6t
72xETnm6jUn+EWRNl1JpuIAMVDSoyoRKlVYCgT/CezW+bFrCqvih12pEPd99WV8cVUGNyUF4Noqj
UcdH7uCEoxMcxQG1oDFy8f2mcWdMHf0WeIkRFGj9DxoPU+YX8eLoz5Rbb9q+ZPGNVc57OH8CMdGz
YtrIihXYMqwVFxjMFRWd7kXe7REZGKQpUP34KVgwq5Q0lfio23UoxZlpndwa+Ss4cJ3UaQRNgY2R
LHtpv2Pgc2YGysKi+xZv0JRzlmX6tUnNAH5Uvw5XARMY4cXAUSNt/5joRIApIHwjPJ8TWsSL1V2Y
oOrV9DY1L7iSsecvl7Rg37kFGNixBwAFVO40DgC81JC87ZUDd3pQOueCw0uTRO1DLeh/8Y+JJHZR
JFfA7qq8nP9Yaq1S3CWve65zkFcP7go7Yp8vrilfLymgo/rWcPPBkHBN5FSRlKsKKhKnXuGK4Ef3
oXO+vE/SAElRjAbNV7i7224X5chyLcO5w/i44c8ZNBveb5sL08jEPKXEwAKHz/+htPngvQoeHzWs
vCmmrsonCWlFOXBLu7zFme973yXMg9OHiQ+eheWcHevrG4aT+LZl7hY2fAmc9lOAkM/GwU2OB7RW
51zm1Oy0eIhR9qb63Dk4WmFu/m1/NmNOwuUpImsIPsrMHKqeoR7j8DVfzsCRVCR3IGqQIUhbzbNY
RpepVNLRE3ugRl9+OUFtwsRgC28H5GDDmC5NEYNk9bObsMWjbY8hZDQWcmXkRK3lwilYD3sw8Ak8
m6+fxNq7pou/DnBPc17F9CHZoLQagZYdDAunHk3y28P6kVqHH1ESyB+KEObvcHsRtSlr9KycVoJn
DkGBFsLrmiLOPpKT3//T6cwE8Nu2APBDcaFkiSRrUOeAeGxiJuiDmk0Jsa4GV8tD8Bms0goMtEd6
Xi25bdLHD9pWgGGFwIgbzdp5qFVOosqi0C5dz4A+/F1oBMSMalYBo8e7vT5hkRNCM7WBAvEzzPBn
0xSnFV4Bw22FtpJuTsMtdQj/WfKYbifjJQ5Z83vXwCC/5B6Q/57jaaAewksoxtR9CMVHXaZFSMXD
AtLU8WnOLxeFELkAl2LupLO3s34o+BZiWdyOG5Du6mcnmEFcttvzJ2hBDR2rb8YIpToNfMQzxn+C
YIX2I6FCCE1mFuUfFROcgWdD5G5Flv0l4AvjW4wUXJUdQtaQVMv7C0tmWdQUXE1Y0umTG3NlPkdl
QK9hsMXLfgJRrCI8KzMNFSb9ky0zqF22rw1agZnLKyB1VeNzMDUpGiS8NOO49Gw1Y4vsccWrbNKx
a5OuNnWVpmGN/ltfTeajP1Uyc+b/jlvB2XAKJRReynhvmTO/AktI7WL3Y4Pwe4++tkc+lBm+B+ST
Nb2OdKSiAEtueZqqcD5VQrGOTsvhJdiOez3MPjTBVRT96jueZtQWIGX/LNyYvfLvRFnE4756N1/m
9/SQRS8e8eKENGRtijbW85qxVHH0tE6NXJrJZP1dFuDGFyDQjmc8482m+zegeGoKTACJEDz8CeHJ
BPoFpbJLt4gnPLV9juJkCySzroljnMrk+pbl2R5UV50myOT6QhJTKNjyK2CpIV+Ki/i4gZoLYTCB
NNHrFv5laEQ/vxrkhE7pwvUwCDL9VSsNtDIA8h9RWnt7OD2roXYLuabnwmIFdXL8TrQS/nQME3Qp
sayBV3ob8m0qyHqC+EH/tae/ygTpvPdw62U1QfsyT6lcxs/sxWfKV8pkLTJkaS8X85tYUFUlmhCi
Vu8VzJcXx9ZiPXjEORke5AybjY61icF+xWjQPtdoDLpao6MKqpULZ481QVx6UGBdY0JvwSwsJomr
6+g7xG9eWpnWvWVkuhLEUGBycP66/V3NYvX8SBN5wo54JPsdsOFxuy/zPRej8fg9+7Iqgham4Vvy
UatzJkcD+VJIpyizBckJbmXvXEOmGD9lDrFVK0VO+aQ71Keqf1lt5HcC+AdkiLJ2ngk26t04MI3c
OF1zMMvbJZoGXKi3Qb/8biDKaIltFplUHP5fHGhQAgWVsqkOvTHoKIJ0myUPVIOUxLXUDUlz99dU
bw5ZribV/+MAObbY13WOioyKg7V0BItPwQFnejpx0lHxhj74u7Bzsi1R12Nur0CAbeqkaI6m+WfT
paHvcja0WEXN1cJ4cHBTcdSHAEdg7HP1vqyybj4AGWEC+N8ZX2xu/nxx5fiimxhXj0ZS3HDBASOb
37tC28rKEem0/7VzlXMAinTPWtmxkCls2A87SSkpVUSaW+tCKvIZEOZHagmaI8M7e75yo+b9dciq
MMZw4swF8lv2Vrl+HM1UlwZd5GUjFfc2bni4evdNZ3EmH6KoeIY0Z/TmIvu3i+1CPpVeMXuc/T5v
4ei3isNpgi+aSEq840NnjXg0DpHY7kgkQoSg9Bgqd/wfhFa6NOT8r0Q5xsW5VjhOWcxmXqCh9+nV
ZJVJQEH/F+LnPWrw4jdQR1hvLPkAWRzcgZ3+Xac7CTFUQzw4Y73SWD+YnhBqXxQAyfTEF1+S6Lsl
2n/V+GNgK9mVjdtufxYjqoWzjJubUij9CKmFWJNIE7UIyJUOAhNZCy6DemY3RKiGX6Wyk9BsiViD
bgRrilNgkrkR/ZT8XV3l7e9FpjEQQQY+HmMXAKZuRRl7qWJOufwRSHsYEWv2jfAbpL9O6UZDoSg6
fQ0RoKuxQmCeG+Y2NSNaHiSsDclXtErgRYGWQoiFBS60VZrUl4/jMlegz80VmKEXgu8EItlz05eP
sQ62L+6m1ZZ5vuDlOkmOQKFFZ6UEg5Kb+ap3R03n0aXMp//asDINRBlwx+PCsSIwIdV6vqgyBwkJ
itS69ijciIHvxX0QN3fx6KGkeuocB31v1Qa/zUYfsFWmB7p7d6pPfRdZOWWtuwVRnijGKuzADNE9
5ifvablP9UKI83lz8s+OgD1TxeVBjgGbTwQQa1YpFPndtfmnD2iNFaMJd6O3SnjEYSotCgLtc/sY
yS+dxfn3LCC9xlpCL2OSWUChpHk4EaI7giA4YlxlZ5ZXOnz5y9CsLkeOxs15kxJJxslzterI60W2
bh5s8RZdtmvLorh1ZEwBiTQFrQcEQxmPJF4n8puKJNVjkdLqLSSkoJwIt/hQ8xK25kA96K3U2BPX
VrNLXbFfWZYVGsJozkWqSQVM4ER/m+CFg+WZVBQmOctP5jj4N8iYgwJ2RbsiXkat7mRec5d4k5rR
FFoYK7ylG0d62iKkRZxT5+ytCrrijhRyqK/vUzctcmssTNr+904kgjLbH8Uo0BC0+Z79cZ+Hb+D5
EaxLK6dBHCjvLcWe5tSqNbIyBxv1zsIC+Decft2rWE9JGq++ZLm+8TsYo/NaD8c2w4JTh8lLrkk+
/yNdv2KaDESkvAgL6L0DYOLn7wuVf6JdNCIpufa2dExWRlMOH7BRRAqtNG+d4mMO7tHPJwEnOFE7
7OgqVM3pxGeCz5cQtCHTZP3j4A8OpEdhp0KjcjciaTKku9p0KSCv3aRctmHcQQOPLSIvBWZlqPJX
jHU0B+Gh06usNGH//K0iwDz3ptEnUs9je4GKdfx31yW+OamE0zxWkxre4+/wMv4pZpx8Xj23p+TI
c7GYeZBy2LpjXYOGwuI3JoRB+KmUqBl3kNi6eEpF8tkEWcVb3AeUSSpgfQMmof4Lhe03WpB/Qtoc
UnWH08hGqBSnHZ9t1Hnyw+MWCmCYzQczpg9fibvQGjH+wHNEAuQfkT45w+Ow6YrHbRHzVHYdLdRY
Om8K7JJrdIx1/jycj8Sy0t9GduF5r6lDccJ7G8+Bw50AT/MChH9Eyp8GCc/osPZXnpZO2EwgScJn
QH/ZdwVhkHzwbElgAl7WLswEUG2IyFA542swaLUVUTqRBYsNw/uWicFCuUHlM4A1vL4X7eUS5hul
tc5sn73Jzpr21j9JiPa0XX9TBnY/3vYB8g3CMbLgClHrySXl+f75PSPdIAa8iq0VJlO+JqmYjxUI
YBT4u2vvY/rRLSZbcJPcy9+oR34K44NQE6OWIebSy6ooz2v39Ab1mtDPwJUnnGTT09LnL1xZqYgx
LKAL03Uuq9/tQEtasdPiCjtYfxO90e+ehSSjeuDoCv6BxMKf7YXAWf1JiHUCzs+sF5tqN7YPtALD
gaEXFijN7C90TLeCx9c8GDoR4ApJvcePmr52GWQ1W2sJQ5HQ
`protect end_protected
