`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
HAglb8QgA5iOr9EGEC38cL4Z9Z6XmzyEvvvLGA+92G0X0yZzkb9U+emlCuQgL+dJk18kqR+gJ4NG
G1mDJnC8pEkn5BYHbOpn8wHxafwEjMLIt0TYLSkW4SPTpc4t7+JwoYM2kpD809V4kW1Lgh5uBz4A
fMZZELT+rBJXD0SKbSa0rXTQooSOrTTP2gTNIdVJYH/m3ZeAfdAXxxwlfFtLkGN0i+TnaOynvOmG
7Ezb6av80yoIglSyxJcuKV38loMcfUR1z72Gpn/iTHCDsaOEWFxwNAl5XJYRtqKT+dXGzd/kPcJm
+PHuG2GgUVvRPL29mZ79UP+NZ+xewd4Ruv+l5Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Bxton2JOetUlLWDy4TROeBRRAnOzCcdQkeTAdYnh+iM="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13312)
`protect data_block
/z+1ufpYZTIMVjbPf2k/bIIio5Gr1cR1dBQ1C3LENOqiUr+B09M64MDZngFIES0iCC+3UQcw1/Ut
7XoD+XTemwZSmw/Awj+O+yPAiI0sdEDjtXeHTwCl9+BQtx9ywP0DzFYKy0Bke8A0ulOpPM20dkD0
3dMLfeH4BaUYxcKnZY6CiCWo/5KIUBFzhWEBoT/ESC8iXpLGJPhHo6GRnO0RJJ+5XJzQhg6dx/KW
3ypdJWo69j/bu0uPXCJOQRB/ACCmmXOsShIYbH6r/MeOR0Lzp0uuJ8gXMYcVDXerZjMGN41dm+w/
OdId8KkPPcETSrRHrkoRms2dCwHQBpWyz3KLBrkAAVVVnrExemwrIYP8v/bZqLt90EcctHIoLWhN
7klGJggmU5JIEWit3o7VePJB5bFN9mT/IojudjDIUeqULbRQpWESJBjdm+htQqlxTVdbpT/BPjmy
AtHSEQ/f2AtggMen/Kwa2hPjCugle5dMbOChGY1DwRb59peVF7O9bfm8uGJQgvNmrLz8xePDudrN
jeqN+OGXI4r+N7ZHH6MqNLLEFwiOaSsfFdQIPtQjdlHBSy3F8Ez/V9+mXJ/0jVEiwifvBxJrN9OT
r6ZZQoW+O48knHQWi9oItoykj9Yw5KLkDo+KaCe+qvevERhqsDSqbZza5ty+Qh8LRqwGxgxlASGW
zDwlewcsRlhosJ9AC/4XLCoshOgXf+kvXzSguDSoFLR+d24fqqSgS7mJSLBDVgF4L/B2DVvI102e
W9AiCV9KqANvzCoG1AVXzyoueAGqBfMyKJZizMMyFcow3ZVCnC9CHdUug9tdkO7XH87dqIgaSAi2
bL1Nj/PWpLUSLGnxPtaNaAbVoeLV/+ZdaIijba6O7JSgS5Yi0RpVN+4fRarqiB4fmV8dKh41p51T
XTQiIUxbz2BMUnYxSDmPnRG0I3rdvYD/ep87PCiJ7DFv/E90nWo/00vKRNTnXa2AloPy8TlN65iP
m6zTvA86RK/TDojjO3L9QQ39BRQCQC9ndxdp4gygOkQRUVDEFwZQUMSaOrFTkZ0rmXeu9Zuq2abv
iRNzbc8iTYTCB9GCGv9kntQGUrmjYm6BqxD5QY5cuVK2XK66GWzoMS9oaqbpOWY5XtFkO76YWFnl
CqhGjFD97Zy1d2yBUmF2SfiMFcjhEZphEX6rVpzjNSl7FjYiiaKBEoWj/cNLPR5m3lISdltPJkIl
CCUce1RT96ZV35c5c2D9SkMz8ul+QwN8eh2mvKZuY36Jvw4/UVXFndK/m6nMTq/2quSJNC7NGWkt
J92yBkZykIlMcZfHazBEBAdCnjHsOJYS91Rfm1CxyR+FYYZQ7O4r/9rVOyr63ebwDC6UeVn//nH9
iSCT6+i7i6nuiNFkHLHDu457ajXQYF86dCKznfKOLM3sj7tGCjm5cao5gfRzpGGaDGRDKFEAaIDP
FRbxUzuK3lyv7KWGvMetL5ZhOzcMUDW/1NQrkJk3m25lXZmPs3Qa7lXj/0XcyInI25As1cSt7syE
7mtHBzNStpE/Vf7q8aHktHill3P2eiktQhz/sG2F516d+xMzC5tsJ2WNdklQEGTKvjrFZUWUKkUm
VX55p5fOBV3CojwABKb3PrgMlANDu67DmNRIGxsQYDb4PRJpqfQaClpcYZvIEeS61P5rC89tp2ci
a606ybAfkWqqtFfN7EUFvJyFNvAJhloupAghFZOPh7bV0JyH9DAb1vzBpTaoSAzjtAxEcAVUwNch
VjFzEQDj1SAKPGLpXh1TSrnsQC1xS8bpvnubi8atu08xFABVqJHsisOyrZT/PySSBsn5W+N+PIeX
ycJyk9AG5ds6bwHy6St+OoQiM/Sx3QucOtAPabI5nlKWqcVcP6rvPhkGWF69y3CspXJ366kIOZ3/
62RC9zskLBHULH7uvlMV5OndITcA36ARb4XaniboWmNDuPmIuPjGLuWAvBvMzfKrJJO26/KLEzHo
cGawB14QWuxiU8D4aqFXHl88QYYZI0Yrutr9T34c3KioTNjHaClCUSxhuJ7/61MIApeyrnDXkrPW
fbFepZCvNwWrM6CJOGX9TkoF0qAYVL/E9YtwGqtyAgE72HiWRKwwpakfUW0YQEcDNfsigcWq+jnI
d8qWhek8EPkAdElcspDp0qwjd6/k7oE5uZqK44dqV3GTEi2HoxkCkZ14zaWfZWrDryVrPO2rJE/A
3yiMECDT1tPdKbsVZlWf2FZ000QsUZUSVXvene1J1lrh5hF/bHHvHTYj844XaarYFHy4MZN2gvGN
7rmppWjsxAebWIxc2M6pSR+fSBFy+Bwv94ETmsFH2/6jscrFul3s0LqF14hggEM2Z6SDCC5iMJri
sEZFMq+kegiVSEKl9KwEgB2ZA82E/7Uie8czTqvHMULdqKXcqB320RcLtMNEXqaz7oST/OYQZ/mR
bCe9f19bP1VIA+h1yj2zQ1Fn6FfTOwLmpa/oyER5ikC8CCqzbgFwOocxX6iPqVVZgNy38ALjXXfw
VweMaSnLaQp2Qzx1IxvcdE2ViES18cOXX/3WlF9LSvvRNTdiyaTCES3w5Rt5r7Oj0S//3Qnor0Ol
fxryMPnD+Ev/Ihd4pvr5OEJNgnXHz43GRHOV43O7/NMu/iU0hAW5zY0BEOAI23ys5pfIgUB/hxa+
2SBcYp8P7ugRgXdP0nrnWkpaAn/2stdPAn4YLH0Kq+C1wAzQVI5/dTV2rQDkwPFnkZoyGsueGnbG
WipmMJjgi29LWZH+NgZx+lKoePmBz68LptQ7uruqLTFs+irJuBIAWIUUTQ0pFgh53Oh0tu3mQwSa
9+qqOfUwKChRTp6hVL9cBB+dcREEhwtD2s14hjwq8hG51dB85Bves1zyyYE//G08QnyydpBv1gGM
5aVQIJi0XTOtEYasRqAkwRGcPIJOJFqD2N8kVRm7I0hCf5FNZYCyGBrQvWtao2bexuJ+BJBDiwHU
BmivjmUDOD4tswgpi5471RpnnuCimPSxUPmqswZxg5iPLsCOMVnQijZYlzy5XeZj4AQDFsjbyLMr
mXHYrNtKr8gxC5XesTYcXB2Y5Kcg0+CNHFJjgb/Owt0x47B5r3Xi5SrvH3tR6nxBixCBIilCdZ84
Bj/qKkD6VkSZQ4OdxwKmmMy5r9gGxWjmRKoPtigZfBXIWlexM84QAEY7k0GjcAEjpUALibUxJTl6
08TjFdztB4EsNe1s7NyRh5/7Iu0gNKgXl9Ppxvv85Eli1NN5H/VqLjD8kDGrVC4rTfW/8dj1tEzV
RmahRsMhsQGQcOApeu7zMm/+fZRqk4ApszHROV8W0g6hCrI/NloBv+xmIeDCoJJRUsZfue7RlG5+
+DBYoi1JjWFkk+SrfPXZgQ4Mwj9+bFWqGjHlvGf9GDQbNLkiGion0tvRtoQuQwf1GKjDER5BUy7k
J79Uc9TkEg4BK45PtqLybE7CJ97/u2poGst5HkCtkLL0DqMr35toCGLdZMFf7yyOQNeWmqekYS5u
5QWB8ffa80P76e1NED/gEGs9JpqhA3UPLjyiFtNEbZHcJwlsV2FObzF2adpBBujEqqn+c44+9utb
GMi2i4i7z4uqDQOvx0DPnmudMsaYAY4znNOSZ0G9MHGYoMkSGK3Tgdl+H53kS4Q+56gT8754uAMz
yPhu7sXNAOC+ujhUxenrp+huOWdKvhXJxj/o7o267+CKiYWYITzonNfcNfZEqeOOyt8z+uMwEWDP
lqOc5QlZ0DZCQZUf9ZNnHjOOGqcx66btkPC3Qdz83pGoZRwT3niv2oXJi0mS731R7WLJSYfkaX4m
fZLrRbvPLGRuYjGwWfrOQ8Fj2Vy0m58sb0uGx7gEwuWaz7+nTjamdZeJ0hDFULuz7VYyy7XumxWC
AvUEd5RTYhKq7BmcE1To/5HxrmuuIEorjRMDsmTLPkVuUyuGjC9upG3u9pFGX3LszIb2k7iut+qT
r1jpj68ROoRWV/SbNBv0BPHKr/LWeO+ulLZO1n1lpkdgJIx92UgycvIVBkWcGzEpwkzkYrgc9d+P
c4MSC1KsMFUUVLEz8h1LWPmSh7x22G7JhbT+i/gUnAqbUBh/4WXL6MQXDxbDZDaDgledqyBvSKsU
xiJ72VBSn/6crDq+Rzh9F8DWmNb5HzP949h+fGlfBq4n5ZvAzhHMifrq+z4GkioDi6gl3tKG3zs9
HBrHVchFWcAeh03/+3HIJD7d3+sMSDJKxhytEt+r/i/Rxc+TDsZG/hZsvtHlcWMgHajNvz9IP3zu
UFiB5Nf1Vs8n7BPNPtuGyhuV1cBe74iS2b7zPVBsZ0sqtcKJh89XZbez4qXdRibK00r6yIotFlrk
sq9OgILHLI3GzT2TPXEGjnL1jp1FWjBPOjvUyGDqJWECZ0DdnzUIg5yiGhSGBxAPJ6TVhAiWN1Tn
ppF30K/NGsRUkBvwvEGsZyJaFBAZ1D4eowceoVMCtjetRLhJX8b7I10G2yR1/AD8N8M+h96XOuBh
W7tUIC0gI22h7eLTiziIFEy/6Ew1aRIZdlkzqHTH1GfehXn06DOT8KdOOhxO7pwybYGmaC1QWq8o
3QXVM9bnw5zPTHV3L2934c8IHLSnCdY0fe05VG6w5F621/YRrLv7GDkPMBJbQbsyisFm4/7aW6wa
UUfVlsifgcaKuY8KZb1euUQHvqizScwrT5mVCztmxuIwekcOny1XFAcqzvRVHsK37ZXZzwYMyCuT
jTkBthphkIOPTMBiTaSluEjmLWJqCa04+8I6EvZNKgv670arTi6l6mX7AfI1pXXQG4hTyOdFKQH2
5C2LuWY8TbTd+23CdiX7Nwu1onAEpbNYNIpNauzsK0gH9VBbolOi/nv2fNPjVyChCPsF26FsnWTh
71X0mcFRLkPQV17t9CgvrmjshnhYX0HJaFUDfGi6j2ENW4dLdR99q6l9+Y5ke7VwWId4sud53E8/
B9EbiPjBHpcaLzxfglsbz/OYwsuMErOAXs49UmOsFtmwtuUtYtaWDj1+UJpTQsujPK+PDGjnVOeV
hnz5OoOkN6GduoZ3zrXfUadTqNRaZO1bh5XnhUaOQ8qoxbfPVuldAPtZ2D02eIgquLdRMk2Dc9Ka
8vBVcHC2dmI9RPLXRh+3qUx35IzmA8/Gd3i5uUzt5PoUp4d/W7D68B5mmkX6x7gBSQkSI84L/Vnh
QDxPgRFE1gJvb5lW/AetRhii4Gc8NLerQkG70hr/V77+3TSyLy9yHsQJS94wrR4ga0o6H0zisXwI
YEW0u4RBxudXaTQL4L/9FURy5uW8Rai4zNoxueW7RKnOABOjB8gAhNqqJwimmILNxhbhnj3hhi2W
4EiWkv1HHzaNa2NljNd3yZulDkAqY5F7uYSKXz3TLeFBot8DtWwyuzCkkrI+RDfUJtXmqtpM9T/P
hqJTgMSL2EWyH+60ZO+3bVKPbsG9/2XYkYGahvbaNk897oSc855OkJc77ikeOkNJcgXDrpfs3DBb
NxUp/hF0UbHWFp040VB/+I42dJto8c1c2jLuNXMlawXgX5N4sO4wCno/i5LhhuT5GLNFtS0UlFRj
Hpip//Gj0ey6eSID6BTUNtT6WVXmihijY3pDJwpGGufPM/uwjeYHgfrRY+B7vIBajIMgslnurxB6
7BRSPPoC1rYV2bre1B4HMYvpo9zRSo0Wx42II2ohjC6O4cP+qBkjYKBUXqeo7i2vRyKFdeacIHoL
VwrMEccdaf71OYSTwtbBnY2J6VhEk8je2TNJfUv0obttluT9lzVqZ+f4WlmBr9E7hVR4SVDJE684
HbsYKtpZP9k1k0a8JdAoZhNxrO8Vxu3TwMkbj7Lh0wZpLgFjkYLVtrk8TqFdsPjo+atRp/R7hbOk
iv8b1H/JTC01EjmF6np1qZSNRDbtQ1qFrOyKcIzo6MCW8Rvv+xq2dGLzLNZp/M2ZzNbHfndemmr9
TBx+0hlCruynehsDlcFj0voCOVc9fPli99dYCEJz+QTArDkrprL1BcPPVreNZofBguTxvB2lcymb
NYDMnTpQNKH8CGpNFhj4T6ijHHkdng63iMtI6bupl3HgDSfVDFlH8Pnm4FEtVmgvozhOCOzN4Bke
sRU9pPyflJItMcK2iG/jM2lxDc2Nw//1GZrGduc/UkjeY4ZRIZ4Vsm5KDhjtFeBa64bFTGm5STEG
JLIQVKpp1Cqn4THXNQHfp7a3SI2N2NThGw6XsdxhjWz2vVdqz8Y+T0TBFQqGdMGbvUzJiuVP9WGl
ZlCgQAA7/SJhO/nGjdqqW5XXL54bFz2a9znykbI/N+6/cp50MDsDftbMI5dS6y7Q/bIE4iCvKvtX
gMEJt8N0zqVpZvVjEi6Np+tJqIoK0lAxr6mee3rrEuLBBQQT4MNZ6QlBq8D2jxeShEZC0rqxUJh2
eJdUpI49zGoxeCDROMMx67b+7+s7Kj6m3cQQtRLF2Z/t+TqBEH92x6GPF61cVzUGS+FqNkjpUqZL
8+KzygZUnigN4MBymjnmApL6E4hEtIcymOTKkfaIYW3kcRV2ZLEn4euAUxaNLSPWxTjg2Zckgfk4
zfg4qCiG4ZepLllbHiKoVb3VQgu5QIxkBKLSMwtHYBhseBaEVwKCN0FrBvqxDRish+3YOhKcL3yC
9G9SK5X2vYVh6BUluJdHg4+ezhzzNSWL151qfqZY44V+37nm9sFjl9MYBA4maeqegCEpY0z2U0hf
fuMSdQjk3BU6aoKdNHXBCZxP+27vYAuZvbNamCHLzE8tZDYOv4c0A1RKX3NEuWL4pu0clyqrKNc1
iz2Gt3Ko5IGQ264wQuMToBQITNkBXzu+0TLRBkkv9ZQYkemOIJFdSNwUkBHaEPDByXwE+3u6+qWN
fKCGPK/I8RrxajztNQpQdowgbZOwWhvoxt15C7bw3E1ZaFD2f40LFn7fsVgIeM2+Ymk+xpUbmDRY
pW0PPtZx8xnWPz+qSB4SdSMTywUl4EUakokiyIpbLGwxdG+7Wkcd8dT0Z7SiALF920QfcigEPDI2
B2MDcpkft6kG/R68G9mJ+B2mIo1uRhNcUzv/MVWgmFv6qaRovpQp0F5uL1byHja1jgv3WrBDQn37
E/wmkJci5fDo5naI8icN7/5fCO+9FUU6IJ8iKnf/YxcawowLBRz+LOhqRnS90t6XfsYUXsdbbyGP
qHrwplNnqQyfRcO054LrycSqtSr7iVxB2q6yECU+T8fxy/S4H+W3HdqMDU21kuz2lEXHP8lu1N/9
VJaVer+zCannaOvvUpAA11CEKImsnwXIsDjYF0lAFJOhq0U5reoV0PYBSUTTxT+WuMBhdOx5oIGI
/Ha9LwP73xUfsv7pI3e+Kw19BjXdxU/qmxJJbZCC1WCu+zi+6IU5RkDdq94Zr6tjULap4M9ZFH1U
A7kVX39E6ShSScGOPrcCT0MEACBgdglGB4dPCQ9vrQUFu7k5Wi0TrJLSug+ZvMtHrZXHtf8p7ZA3
SucSC7KAGwDA2bRFzGKK+hJ7Tb2WFIQmGW3eK3fMiIOf23LhqWW4yUOSm12k4lhd1LAbofSEjyVM
onpwpsadUd6CXHpk2XSrbIxpdytHuy1L3X7VkVqpgi47I4nPnnyumv8C6WKAvX9YmCp5PxUlTzvG
BSbBn/qT/mnVAF47bE3csa07OpwVzcKUhw62+Kf+QEnZoYA0SeIZZ7FZcq4gaxc3aLksYMMI2CvF
GOvu3/ZUWLIbmaLWH1idr++sH06LR2qj6dCt5SxdiBCJhkinyvxSRvmPvKCr2xxCIhEgOAn/n7DW
d2PpalKfqEmV4tC44D4OpzhiLXTxDCu8H4D35+vxFGTov/QeD7I1YyxXde2o+P+8ir3HKUoc1J6b
Ioael4tApHOOkvyaaLRBbpHczcmcG7H5+jssyXSx/0sZwKBDW1WbKVliqaSXO7YEy44Z+uhBFIjC
1wVc1t51FF/4fT+EDfRyt135pl81xiMZ+e1vKDKGgfx23QndXA6VwawjXt/BWQHre+MWo98FFFLd
yXUhuQYTI8hzwg/vOiR9cxavlip5XJZjNMsSPoAxQhF8+NEW6OHO36sbrZg1EAQqaNZ3H4jy8l25
E/ZcWHfA2PhBA2+CwKg2lbcC7GYKUEG+/+Gq/cKwsUphhpZOZ0kOBCyZyc1bewR2ZcBJRcQbedwr
BNqocxnY+5G0GYrFI2RUw4n98sqWRnLpcD023lIznPd0FwGMc+/WPqqI5Pdewj7BywIceecnwOPJ
cKBGR2Uc88C5wU9uXwVNSDXL8Dk+FAs+4Ap5Ec6xvs7b9UZLYgk3niRXJSEraHK1U9beBqqqpuuC
BIHeRSAjp7NUtuufMk+BwFg+P5Tuq337EaEhimY64qD6g8oMfMbGi0RJu/L+pmf8ntVILvRG729W
DUPE/83V9yRUQ4kSRdKbKgzaDzkbmlOj6vE7RjFPZlLgwykVdB5UMmDqN1tAvscNHh4V2GQ7K75v
V+OobkEAW1Aa1iFi4LJRBUzGVncIo8hdDGx5yXiekPMVhQRNBflsXYoiT4iAp26AeTM9x0lulqqv
qFfxy63/sZSLvIRkuXQUQEfrWRlIagWq/FJV42HXaa/we3DPlCLz6+9M05L/oJ5UJdC7FCWlxxyN
38Z5SS6wk/+9ea5M9LYshrkvyDYxCYZWiog9M1SVF8L1tVh9lV8ksF4K/3xRfzYoIKJJfrRwr3u+
m11hmW9V2dAtjwphZzqEWGIPFVntGMSeKqLJMnWwIkmUdANVO8xkVyJtHhO4PoAgD6O3E0EzMS5f
Y0V9M7inpEu47Rp/Rbvk3cvspBqlqFL5eg4KeME64lub+D9kE7DBfA5iQwFKA4mMgk9LPAo+DWF/
6/JfO1Po7YiDbAhrtQHpSGtjg0ZsJBjOPt0NI9qa/eq51V16x5rP4YMIyVrotKYATyOK7ahvDpo0
BKwmdEpBfWTE4jCPKIFPPdV8QOLwP9j8JQaNIUJFC83EFVnL/FgUjXG0j9JM9GDF1F61cIgJl3wf
nO9c9w7f0ry9s73AgEY3HOaMO4QuT16RnoPJ7i00OKUdETxa3yccHZKF6qgSUxob8GJKgEPa+2Dq
GAfKL1jwp8y2zVTrZ0dFM3tzgxRDI3OKohfFppn+a35mAM5JXWJEcbV8spHAOyaaBbdOIq7XR/zI
nmbMh8gLJBQGtITm/Qyq8ImL7SBk6lDyJ//MSF4TWkoBMRdXgHEuSDNy3Fdnv4E6BQbjKHedRI6t
5+60T9jgJiSAB7ruquyJiyv1Xh6aE7if1vZXd4Kc0D4Iixd5iDKuGk5YYatO9d8EJZCO26a0Z0Vk
o4XWNVHpF1tCwWpnU84lzRH1rrquMLnwQBCc13j0rgEb8IMvKhqquiLki30rOy5sp6IUVxPGxl1/
Z+e9XX21dtX1lZf1dm5f3v7nYKvlQmppt8hrZQsfNGaj8A0UKq6xYMWSjYFAHihEwWG/VMKqZvB9
111HyZOk5ShvaCRoSThQJct4S7au0hwztneV/IWymiETVvYEOVVWlAZpV0+otlyW8mLr1SpZ55Ke
83u3O+FppgtK7ldrz3GSrkN6/oCAqVePS/asb4+FZA5PoKWEJ56UuKd1IyxPnUd0ll2WFW0qxx8W
zFX1Q8ORdIELON7LBfbzNtlo+T2L8se//o5kr8KXH3AxiRd4LQ1TaL+ukYVU6lua+yegrG9CLyXk
LeZGTeEsKLJ3TXw6MJU8hMsbipyIuTW7duLGCbFimgXI3TekPMVQqzkbAbC68OXPYm5aue5WP3cC
OUVjdiN+6UfNxwp+H56Jaw4gZl0a+Bs4WQJKklzAF5SX+IMvlbLzFeSOGzUajHFnIKWXVsBIHci0
ZNQhiaRvDXfaJU8N1dxRJ7MOvMfyhcodFgk0g4drIT/oTNAW9j9Irsvnz7QEOgyAeZdcV+cLVqEI
3DT5RcMMZN5R0I8nW/pnd7/lmzZC+o/kpzPeada9BrMeavF6nCWiz6rS9sSX3xCuG5n8bmVIEuLb
KWIsdzCX7tVOdD87Ij/DNxbiXVjoeoHjMLgD3m/EziBHmeo1Llck0GvNjfsnijWPoCkuyzYM1VWr
C4NmgMK9Df0i1mpZVKbbAEoGNAYsOTZdZeYq+x5UK9kgFm0QewkGsFl9N+p0s/uX762zZvLffXro
hBRjGHC0XvPFydETFU9SKQAxCJkRUgBGzGdJEwQl0Z3b+ICcWBeLowvH5l6BZjlpIfJu23iVk7Wn
KDFyGFrYkMrjVUyBVnuP8RnyfTnO56vmbLTzAsvzF7WGnCgPkJLSBkFbNXM4XTnagqIC5+7wjb9P
RVs3c09UcpuJ1DVl4XVpfIo64T77uoJu99NB1IZvgVqFWwEz7rYBoZSg7D6Bs196ZIqGzOfilsmR
a7EAo2qwL3DFc+CFpg6Fw2nSjQB0VV71WMqjVuPZ99fFmv1/Ko4OFGzDzg49K7ehPIRNg2piA95T
lKezK0KL3JzZhTvciIoaRmtnP3oVpb8HHNNaLMTuTfKvnSkRr3FBBY99c6nnMJu5AhU4vRACy6yV
oEwPgw2lg2xvqeQBNTx56NXwG9nyTiCDPB6wYFjDxmJBCk8yafs3q2R36PaaMUjIoDjvJ2skucQK
LhW15g1OGyo+tMmNGfmPPIkszpvw+w3PBrATLQlF280rxJHhWvR09n6l80qdZeyhR+0zZc2quEnO
+r0sekapOpB6KhP+KfDtXC+4E43FUHzGUSdD5M+xgNpO0PQibf5DvBeReA0cxrQW3teM8bXpONM6
wiO75KUqnTHZTdPsOUPuVoW68fiGn2hcWffdWmuJghaL0dSuBTlrj09escXgVo/b/xJCiotnqcf7
UhPw4mYcvZyB/8eqiOkZjf1jdD9CdnQEuaMNHL6/aJAGcJZbwvjzQDaRTzBIcj4bcYiLejIB4Plc
Z7XsiPiWA4XELJPrZjQrltjD3d1DkvA4GLkmzXAs7MiAk7OafK8gTjMX4M0m5sQrIulI5P2kvyVm
Iu92X1t6ST61ANLsJT4Zw46kj0pcJZIY4Hj+KVFShE0bkuNRHdSSZnZsDCNjJQcAmZSshFAxMZsQ
62rfYBX2WEWcRTgqkjhFDSsH2WHPajgdHvcqCYAfQhpkyBeHFsQQC6X7yEfhQd59SQYVnbKQV/6L
3+Wx9TDYHTp+vU01WJkMeh4aI7gXVozM9HLDEKqaxTaKEGsp+ExdjCCQaFjDLT+F8sIyluV9nWB/
DPsylp35G1dI+HCzd9d5vpzjd7WvyetDVe+B6yDcTFjjA8cVBJWW4hHYW5Qi8HPJrDEKLpjtebJY
0uMbQ1i8Wvd8luGsFTZ56FK/QtWQ17kxX0iGKc0zWKf+3Syb3QMKdOF8zSKcCfS4v4XKViDGiowG
K3iNlcVOpsYvEYqVHXzHr4bwYe5jAPfQGqOwkQ1nC3kgdjS8pRiQSzHaC1VYN509h53uTcpy2dUN
4fHlqg8H2qStlrRyKsPjmDL/YbSTFXteKNTci4jaMjoyImg7/YctIKMr3cej8HLLZtyo2V/UgS5u
JHsxw2XT7RSbxgHyJQzEHMA3Fk5DYtws5+/EvubC+ugm0iLJ4Cq/A4L0+U/UfvCKtXFf5XW5cWFw
YCpiNED2RJRY1nXwv7s8R3DyE4rSHpnTkMg4xq3lt4KSA5CyWae9ZCD3AZPK9tEmPzc1jENqg7uL
YrIZZDsfdslWGNcP5NMgkXG+gQLhtHvxbRLlvTwjKgC84kPInAVsns/URuBlkIaXa4YsJBhrpHnn
rcdIk9vzu9ILCEZNhyaWOIizG+u3oJZiSG6/10SVvmO2n0s1rfOKU8OHoY9VGuOWjbs3bzhyMUZS
1bvg1UN7bCTMRaZ99S9MD5nxudnS8bn96I1V2+zglaDITmJ3Y1hN+yXdY/map68FmDuimivt9k8K
+JAe0nq34V6MORqLFSvYkLfW4NBzUBmIOZ1i0T7o+varUiOvJShIlABcZdv+J35cm2rLWt0An3z4
CvISGl7BtJV4IBNFXimoLSJkDeucRCbgbaiBeV5glW0Bpj5Ipq+youPLg8AUDUUm9BsYh1kGeH6C
I/vpDXgpd6BFw/YD1gmFYZOT/pIgFxFIWLcUcUYTsIbMLhvJmRTrK8IrqsVFSyLdXhy/hkXAk7cI
aZO1561YVt6amx4Yt8E3iVCK/oMdjqO/EuHuci4i4JJMmZg7xP8h4wZ6kqG7cdBoxjc4YblVQ1/e
JjZJxKnKmsWp2O8UbuibTr3l9vP0PCq4nql4Ok4dfwMFmY1PDswkfpJHAKRD+gQlwf6Ap3pDvi4D
1+L37qwK7ZAEyfhumJ6PpKfjhe3ksDBRAREqjW+PfFPjjgKw1jz8UN6x70wDZrN+hzTFMV3JjIgi
4YMO1MvukUuvvFEtog/K5R3dLmvXe9qOLEEfpw1dbjR6gljw38CRG7k/QIShn+HpL9+tV0HXSxEl
P2iTN6NykhbWAJ8mvuMetKTwXAle4XlmNxEplzW9wT+q4JOFwtTXXFbjSjZUy1cInTAkw4AP90gq
CPo9UEUJJJrF6lnvF5EDpEp1I7/P2b0OAyAePzxcgzxRWo/efaIdn4eUUL3nGEahRqoxRBZQjCR1
t/AlFEz98EosDJaV9I+rt12XSKevNfOkCCtalWiBDwc80cpOlrY75Rt1JYLboQJecACbQb3GfKPV
/YIMZXyOTygRcIpvR5uhOxjy6VRWAXkRarrgvgfiwJxz7rnGsUgD6qsZx5xQsEHhnNunY1cATLFw
i/KHTYJ/V4sdwPMCl4xC4uU5XMrSSw81ekc2yWgMS2OsQnseWslnpax4kh5HUQzODymv5rVpm1TL
cA94kQOHLAo419Mq02wx1pX/TihpJ9Jy3e+uYfGhN3eRzQP8hNGiOCPObbVTh2LBGtErDVv/kbBI
bDs67ROkexzfBDVPec7QybWOgB0MA28ZRfUnmCBXnwhIsMIV1QcIL/DxZ40Ut5bcs4+H1IA0bfF9
IXq3Aa2q5duBfURXE/lNDmfiHFnA0Tk/SAK24ArnfX0H1JFSluYvGPNbybXM2YvOFLdn6oMlAKQf
+TXayTrlXZKk1WUZKjNJsSo88SjTe1I2Y22f7FzRlGu/lDcgyKduNcx3ac7PgyfWrxio8piFF52I
K9k6wEqO7pCyni3ttxZkNVzyI8q3ZEsYGhQGCwUcu2rbwVZMRJXXyEVQ9n2/Zi7UcLUO+doHTZAL
B/Z0z3hehIKM0kwEEn/Jx9BrWVdkiMAkIbL67ikdvUfrRk3/NpNq5W7Yhp5fxp6Hh+p+Jo90XxVx
il7/Oys2ALYoxlLvP20KtjkTFJL03o3bEZz9tYcRSReukMqxJmuoFCSF+a1Pc/6tMI1uqH85XmRA
eFPaCZVSbBwPH9g+gLdlq12CMUk9CE+NDyhB5kvxaWiYYVf4Bgy1R7YCA3tiuk2AvgsA9Ou9aD/Q
ams80w6tnGGD9yzLygyXySNSz+C4UqFqUl6hgGB8pznG2+6lu5uELuDbL/Zlm4S2mJU1fWYfNgKy
mqwzSqT7h7Rb4qocpZzLSk8A3w+zs5U6Q5i+nuWT0Joc+2AXE9LNn99F9brljd+qdDtqyeYLjmrr
bH5lGbb5vaGBQbsfGJXrBx7kZKBX+SnIqccqKTC5NnBuUCV2KEPeR8Qa5xV6tZK5/XXQsTvXwJ29
0kquHxrJ7jkS9hMHO/dPFXa1v/iiCGEapyl93/jouxncf715/10jdiT6iXbEf7H42NSrQXjNf66L
cYMxvCp8ULFoTBc5SatmQLVXJxpTpnBWdv8LbP5DmaH5DUFkkFE1LTXCT1dzFcmZuofUXk6gG4U/
i1RPDmx55PQ3OVj/08kHBHiG1Zi8E8QvBmUvMNHKQv7VQJQW3n87C4Wn1mT7ZE6dXAxvSgIt6o1+
8pKxYLoU6xoFUj8GlmDsI1eLeIJQnAQQAaUNoSGVkYI2aGJDva5B4r5bAfPPO3kqzXHH2wMHfw2X
mGB45UCO/zaFBYtHjv1w9q4isN8zaHrqMCw88hokyyNj5gmRoN2jEg0VeyW/J4qDwQIYTOwtvidd
zg6IefvZMZFwfzdw/sWmUl314Ofy57pDN7RS4SEnO/zCLw4/xrnWOghd2W7tC9II5f/HGb9+ineC
DCRRXkJujcdunyMdmaGvrgvsNIEIU3ZmHEoWbHl4+kBs4iIEzEFyTF/RawnC+2a0o31VF4bSbm0B
e1Iad2Amg7ClrrfBH8b2HkwGbD6yEfVOqETQMfIfteESYzGcudnypo64mhTqBP19oT/Mq+DF586r
kFQVUKXrgDGGKXaixgMHQ+ebdfmTF9u+GcsHsVj/uSH3Qr6NxjYGx5LbCyQ0bbBVEXFm/ab5uS30
FhpToLY58PL6JJ6K7ZqupDRcihxuD1GMEgE+vxKqDjem15kdLWufUI2TTXtvhBZatmZ2vqAX1eOh
FRu7VFWl1WPrXe4w3asg4i9aacdIAFElOoro1snKy0NsgM/6r3JhQP2XUqoOjU5vhtqDgev7LSYi
ZcRoa5JbBS1wIqE3+XVpiE9jwtqzM9y0EsxR38bl8jAc3VkMIPKm35FBZnnkPoRqyQs0B6ta9zYT
3I2r/JVp+UVLdevE8JQELpCqSzkT5jQLK418WTLeOtufYXE0+aF5uSK4refHlHu5JUeu8ka6SqIo
fMbtoDnz+PtaYkV8yCR8z6PbR4WFGX1TZAU50POTQF4FNnDygU+ZMAJ5YsGL88+D12OHpxgnjgmH
ybQB0BUJhoJEdDe5o1JYc948fKE6gqSrd13SQdEbj6cJo5cjiFBJY3AjvhLposjES6dVs4Mwx/RK
IL5HyS1xqL5MdgR42IvTN/TfPuQdNXvHKjnNBXe3D9ds6Mj3alTj4Xv5DxgplE204/DiYRpu5rKv
qsoNNtS/LTrwLL1SdkfwHPnulfd/tZBvC1AHCyUteNXEy1lIRbnS82C1lH93ascQ+vm4fu9Vm3z9
CDeJkfYulicwDV2lLGPXg+zuQQv65q4cec7j3W/InWsWfp4IQWNB5zIOUTfpz7UcuRuYg0eOzZ+f
zo8bBqlAwd11kZtKzVSMIpSXuxnZsobAWUtglcOBSuiq8XG5R+wnwttJdoZqEE4eWurDc39UHtMj
MpAOifWqO+1b32fxiCaI00A1N424suXWCJzwKnAanW98AEX70II6qKhTX48lw/UZTyW0y09Uz+zE
+W8nC0+UqTRKp941GEZ3xc3Ok7HVZA37LFLC40oQJRlD4LUrQyN8KzlfxVcrvtU7+Sj+ikVy9r7d
6SlD2C+V5oSsC6Y9v6HfzLLwOwtULZ2w5QWuZU+Wt7ApVkgaSITjt0pyduJaq5iC9PPNYDF2HtQC
bjiwuoRJM/sZi89DpX1zATIF70OWrrSu4f6R2l0izz6h48DPIq7hGCta0NJNT5P85UjaD/a1Rqbi
9k7PgBrowpL+PzGSbFgxo/tdfD7YM7nRowOhvnQNrjvZGgTLqTsp5J6oKNh1eejjQBG2ws99yvJi
kh0y2SC6AUnJ1hyf4E+VqkwZ6SI+WXSMlZgXLi80svkrCZBI/mWSRt3gvBjFDEslEZVU33lrUKNr
t4GgIUQuSdmGC9z6LxHBkBR80/2i3uX7QOh6ebk5QOQpq1hvPh4CpY79lItFbXwRj491c6+89TNa
4Ou83TBb2qn2bTQLHs/L7RsXxWJzVICG1clxhz59vQCp4flCwTjYbqLqovIlGpBln+p9BGeO9e6c
WHQo0UKvm4A8VJ0k8SCCr3p+wYcj+LQiSUD2T/zDP83jl9acVTNvSHSHW+EmeYTJXbrROqymZSgx
jXn9tT7KGNVCG7SWOnwkIymtTqw+GnI8Jb84nR5up0DDDNYST1TairQmmHHUEa3kn6JoCBzs5wdj
lcxHGFMA3H2LuA7oHmbV9meHEC6seE07WPi6EgmVGf/d1xmyFt+42/Ib+4QYVGI2s8+UKAZxI4gC
a6uQK/ALZ9OAXIbPixfKhBvtE6MVnXL6lVly2dvJCC7S+OyPiY9uLzTiougz2omWMH5Q26IDf/Dn
txplxdOcI4+MGWgl4qSdfSFA8cNSUEuL4AetdhP6Wk6m+armglMWOK6M6fdg11b0rcZlJNEgjyVQ
TvcRwsW5KRUkZx36UcilhZ0/c2dtGxm+uKhtPYQoa6FVrx2HvSTeNMgwtDhcPxQjewju8VBb3HTN
h9RC9/+fV4oBG9YyYRimPzt5nFX1PMWNYIr4rY2W4qmhuyLcBu7dO7hPiI2QUWXwHVu6B3UEnKjF
qWkyPRbqt86uND7Va4K8U4uXlm1E7doTqo9FKG1HHgROrIYa0gxqJdd9snQkWSsqqqqcudLbo5f5
9CyjruLbiNHyTNv06AlgXc33tBk/Og971Jfne1vD4nHJMD27drcjh1D8gchvPi7yIYYOencwFUbz
vrfcRU8wnkXVzD+sXiGYuKBOGRCIosJbg4NJVVtV8488C4AOKlUsX5ZbYzT/Qswodi9KqfoKT7mB
J96yU1q5mWuhNP2XqaFFDBAJCmgElvg15Wbc+a2vY0fsanDALPe5xVR/6aXmcOfYhDyGhTWCeisl
cmpC1VbuZaHyohlj5y2OU54IFY5vxA8a20AEgkoQVy4wZKBBIlk0RrqXS94NYu4eeBMG/Tf79oVs
a/GidvTD9vRuLI0DWrI02QGE9oVEI2dKQuKy8L/p6bi5U8Ejzhl+1Wz1tEa4gv1tPxyyDXEqHQu2
HI1o3gcZfyaTiFq2QAm2oREFrcjZuOqianVT/G1C+Zm+4Ew8fc7VJClaY8+nKZPbERDV+TC6YhaX
3uELfBJAQmdJq+6uBXoN1BnaQdDmoewURWN1C/ItM9AU2iBEC9vyDljUcvFWm8oXt0HbphezWxgI
LF/HBIc5Crf++yHDNty48dxREPRzgnKryXQP5CN1wnriogKe3fhlDqFmxZiJjgfFSkDVytON2lHl
uZaZQg7GqKoMqS/EuvgvHCLuJiGvMFQSfYiqXe5iDkxGBLjT5P6vFxNYM2XiHphf4cKvSkf9j0v+
nwvsE0H8j9L5t+w1HbDMdV8jQwKzExyBsqzSpdLD7M9FmCbbXTl8hG6NECjS/9It5Fxnsscu9yly
allwFntK2raAgr/kd3Z7GCASz3N4D/OJC0BDBmQ+F+6s+nAtFJm8BZ/M8HrU3CCT4fOPRk5lYDmk
6uURxmeRGDZqA7hYEcg5BPWW8SpGxRpOAjB0X9HnFwj813tofffyUXs13HoxYyA4H/qdfYTaDg5p
0skq7cqLTAdTpNqMrjzC9m3mNF5y+O1B9pnojeB+29hucXDWm8HYJcvpd39G+1XOeJisz6qU2wYD
C0Mz/421tAMbxRxMOyIkF2sIeLAv2y/LnMSJjSP5bc04owZ7mLeVOOuord3MlVX/3RZSqrw5y7x0
sBG4CPQ0IfGK7yNvAEqbBghtbazltGBJTjNXRLJtO0veM7Ig2X8XioEnlPVZaksNdWjkVO+4wzbZ
lfO9BkU4kZtBOcgGsJQzej/kNTKCkB5GzNO3vvysa0dEx9Ug5a9pM+jriXKoKtXcPu51YkYBq4/T
0F7+b4qa8Rs+reVLERjc/D7oB9koDufAJSfRy96Eb9Dw4JuPuN/ghpvYGqXyoCczuWXfSyzDdCZs
lYJKYIfIt/WrsRG5DavwsjWtGVuOcf+pmr922Lr/d76BYUlsXFHYPescnpehM1tz/maTlfQB7h0U
r5YSqqKYPQyKRO/7UaU/knhZGLbdR2YD4lfby1aAzvfDsqu798SXvHM/TMV0cIyJnS/mm2FYkyPg
zJQWgdCbZEXRbTY8GoVsQkOI56V6YVnXWPXROzcgsA==
`protect end_protected
