`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
QjuPviAoFHXDFbhvRZw09ygZS9PizPJ/QnECJr3AP5NohQwamjheZGGA/K+DZhdzWFfLkljegrcr
iYStK7ewm4qbHFdeMiE0YqzbtARje5AJnAOvEK6NyNedXVq3OXcUNjVS2tsEajn/+Y902PJZCTEM
rBXawJdYI5QcWg7fq5BIo1jmXywyAP7XxAtdpBlcR6fNZH1YqnjFOZo0dwv+A9mwFxtODmC0AoZT
3mm3QkKujH8O9HHkT435HV2SIwKGCaNBJ/57pLInukqHvxb93g1PqNqitqyXyD5fuLGNzRUVxJdu
Bqr/+r2y+YGZJrJXbhpoFzyAGfb2/kJQH/CpEA==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="dLofVtki7KqE+4AmF0RT3i1iLQskXcDc4jupUSxFkSE="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11968)
`protect data_block
qw6tET1kF3sD/w96T5Nkx11aZVgGOvF9bjJ7iDT6Q5ty2wNZMfH4BYcDBvdtz6xTenJN074O9qLZ
cSQeSRzcSY4f08JCeC6YSZ5tQ5mrZGh1lZdPFkAqlL2BuvvIGhPweSMO04/VLiehNRpLtdbZADaS
PsoVLCGAx3fgmGGVxC56iiDNtmZu3jyn5WJZLaAdSi/afPRExraclQPIfe4/b8EeyQU9g5U6BvHa
zq4JwRJx9T6tqlnttdrlivZ21HkuF8QqJmAaA4sq0IQJnCiBPfHS0iorNrZmfYRjwa6PG7yUgOpQ
XM6cjQcCTp+S4PBBwN+LzvgG8cTWxb51o5xg5f2redI/M+JxNRqLv+xLgpAlPltOhQ39Gg4awtSk
M352NFOOqXYjeDOPLJJf/H5X4tXECvbYQSL/EXui5dJXgQMK17HeM4HUdeiM7syVVYfkOAAdklA1
H4EJA3D97vwAJOZ8rWallsqPBBuJHEVTyGxzVfIhHlcKe38l86tUHOCbn/YDcei24021zOckzvr5
IBIFuksFJ3ZPnm25NuJhg+DOrCsFgJ1Wd/ki2EG/L3dp1D9TrfhRYYAp58OkcRF07Pg1TFJAO6sf
LRBmvybHqobPZgEJNIWzb64UTqmncfsD1KCwkud6X59TGcaEJJB9U9bSOqhDi2GUY0MiQHyFut+e
T8FXqoxoDbm91FJvuqSP5YOkiGoGCWSYohq3gQx00ibh8oLKNtHaC+whhMxsqE9IVpsv4vn2agjh
NCchKQfy5zCzjYUxT3H9zSrdE2Xft3/DcVFKp2evCo6aL8CyNsre+srgwmxILgB4AqSgDwpSR+CO
NRW+QIKVDKZoqLuq50AA0JcNA7Q4MMJGDdRoNalBy8/07Qrb98/1JTDu6Lb4WAlFr8umQKoadOBE
WPte7lVBdUJnOZUQq+QCbs18e75JERBsi1FFRFB+rjMMNtnpYZN13hu2xj4rtr31/mFA2M6ss8R5
up6X+bnowejCnHmgC5NRdBC/Khv4k77Vi5TUEjB1xvN6EIIOyXsewbLt5P4RpOs2EwV3zES+KoiT
5mW0QV3sTLnKcz9PEqlJai/n3TupOLFhUPWTg73UFBaK6yQYiZywkTQRqQB2E8oNfLcJo5JISVKG
PAY2aMRZotkcULv9mB0+4ZnU+SdiN5BqQfxK4b92ACHzgVwkdVt3/JdC8tVI+py3ds5QuD2mnbmf
x1WOccJDRaVjf+hf26FIXBZf+oQrIew3QAclnkRjiOZRX7OQ2MB6gz7skYiD0DCgj4f0u1eHrcBd
TmC+mJ/YUNLHizHK1GN4r1jnjhnq++szRJcyIV2bXuCaVlE3+F0+vxew+pvlL/ZrGgRv2Bq/EXcQ
5CnBf25GWQ6aOhtxbgz4UJ0baOEbIpbPRig7LVhDIePOt1FIr9zfeYzOrt+nZigI0KVcFnRkncR2
RqY1gsxp4/YK/nVizNPuxpchhtb5hZrSb5vpApeBO9GN3IQbE0rCBOq9Cbkz2Gb3fr9BLTfenk4f
46vzEh3cOCeHmqKMGEQTe6c+YBusUnTXrAQhVJzaqsFOXzep5yMtVU7oW+G6lSDeXi6HUv7QjnoU
XZcF8EeasF2G5xEUrc7JJbvXhEo0XDT/xj6joxYsKD8KO4cRgkjIofhhgpw3F+c9p8KjsgtRZxij
SwnRpJia+IBYjL12wLWKv5X1BaM6kuMrPiGm2rolyXkNqmBfucbLzrRyqs05RbtGMs69mJ4Lzdjc
bfYQ7KZCx37UeA3Qw6jAoedbQH61g/g8uiY7CuPv1o8msES0LvuEk8gghhlvQa8ZVOyJl73c/iN9
Wp/TLIPyrnodWUe3+OciU0kLo3Ak6m+4+kOLED2tWdxiXY9OBZVGb1FKgV0afWaFKtyNSNK/akgm
wThTevsr/lF/viCpBA29ExTwQfVyg0HHFYCkCIIzHgpMB0oMON34KVeJOdKPeBW7DdWv0ROOD0Qp
iPT4w8AMjAzOikD2jSSXmca4FSTcS/RfUsnCWVKoHk9yeomeqK8XtRDyk3y2NKMIuduQTtYvIyTK
b2v0NkQBrOUiZlNiBlqbOjDeAhME5Fil0kY3AzkqOwzCxJgfnimgXUfGhStir6Dojs86f2buBN8V
Bi9KGiblCNhHM9KFRaBlZ86fpGJ35hlx816qjtI7Vn6lPUqJbjjJPmwtCWdIf3/V08jLEH4mTl71
AAYK6I9KUIR65Ie0l/HspXRR60vS34c9r92GxCciDUJLBUR29Fr697jtmNo6Ap+JNPhhkB7wR4Rd
Z4WOD/PWmJxJ0zeM3VqxV4BAUZHcNFFsoVJ9znmPjIgfgIGEc9g6gVX5rVHBT78AppZgzQwaLfxD
xGReXhjBhOdbMjvSz5Q2A5mFZpHHWdQ+TYFUeOHm921vGQbSE1Xv5WpktEdVCTaaZZLvGuaXd47o
tlSuNPLT1JgA6T7+qBjzg/jmkmKAMed+3ZwncR2m897Oe6jAKYCY7dDyNCzLmeczSL5+vM4BiMTc
/lr3mIL3a3sId/pTH1cUIfY2fNoveDZ/NE2+cLphN5RGTzdxDLs26y5Xj5seoYhq8aOjkzZ0dNBa
5eV74pK16H56KQOdFaMe8HX/zMsjVD3qoq6JVS9ZqQdD3mnxKX/pymrju0SeaZx1/dgmE2oF0sXr
atpwTnmVIyJhoT9NJUbpaLCZ0bbJK4QT6X7EG5eO1QyF4QuxBWPaJ8r/2sgdzQQdDXrNYwNBMtBI
8xEq1vJ5WoDeqMKdFfey+waoVyFu1YVx2woivJd2tJRIgJZu62AtQYTQkvaz86OTj6Z9pOUXunOK
pRX1SC9W/4xRxuzjYIovRDqbBcGJoJuKKiOXi2QxXEPgzTMhy4BI+HHWTPX7qM87cmqxaI00V0mB
GlvAyH2UWUxJdp7EmfY7dHonC0ifPqqPIE0OZd6Zw2aVqef57Qc+iedK1o/yHWFy0YgLeryr0bXa
hTjDcV7eOA1IGY1gC/hai+FoS3jHvVJ433DqJqNSZcMRVviJQPsNPQ7aM7cHZV4csGKCkG8x7VFX
YhVukB/bPzfFHPjCUMNnAspXbM2cJlUVerfN2ZbKcWTJZC2U5GjFV0FgvuC/xUITus0adACHpuLS
hAonsIzrd9Uw/sRfcBjvU4qWRerWYZfwZ8aY2DrFwfy5hJrArejSQjNPDss+KZ7t916/HHRxuQJu
59geGM9qrtDXIir0gNeYZ1SRDut+OGckt8FxzSDtNKm13lX4vwgoFEcVG+KuAOfRdIkgTPHiMN4F
Hd0rGciSRR9VFnxLL6BzLag4BuWFnY7T+7QN+vbmbewgylgy3CIAimQLUGiMzQyv5WdWvNxGTMZf
5wplARYeUCjPc9O5wvCvkX80FDJcNcS3Mqde6ZvysrgfDGc2a8QFYZAF17SwRLMiUeZGMhEU/Rzi
ftx8zsjDgdrPzVEEsE8ggmilz/h/0PbF2mpSyEw7H+Cn1ckaYY3Yt5mVfGn0A5pwCMd/XO/e5T1m
IWHKfgrWPvJN9Ymt2f/Y/fP21W++9rBJA7bnBSEf6t6YZ+DQm+I3wsRY/EgtStB8fdaJ7mFhMPoo
9HV1FyP++p3dCkqrR1YJ9jaI8C5Wv64EsNs+LaEx+EZq3IAByrUptTT3mYtS0tNfv6sgOfggQeKG
YqlyULu7MVmqjUeFAuGpwYUVyJOS3Hg6gT7TO0Cgseok2xyY1SdzDqsqXmFwppBZSSMqx0RKMI1l
zNsAcHMyfyzFlk+RYScBni8VBn5dnDia0nYIikxBkZh5uPoYlu4ZQey0KjG/we/qkiQuMKxumTvy
KlDUwXxCGV1BtmNy4xYunVclXvl/PhEKn7t+NY2jTt9pH87Cn4iqwHYdqXIjXRGgz6xQ4s3Twnpp
yUh3nuApDqtr3YaHPtkhXJTlqwvQqEAr2geFCBZOJAaC0P5QjNO7U9NjCvanZGJuASQGnxQbXI1M
K9YqAJFGCg5JC+JMyVCEfEO1kbuSDfixJS/kojHedN5GdRmv96SjBNHEfdi0kxuzNHiKCRvx3WnM
YD8elgYi2QkEWST+gj2nmIFdQF7R0Gfyw4CMQsxwZcrsC6XO5cWB6xRzxumSowh344tRBuZH3HJt
m4x7kBrQ8zwGgzjDvdQtXRhGiUuxiU5i+41U6e1aiH0/uyqDHtZMcnewn0ZFaIaJcqgZZ4XO9tpy
j930S7lO8zDG93YfHqcep9mqh17R/4gdY/usZetosFU3rpDGFuB7DFv3aKvFFtM2vJaUJjndZigr
hMoyTFTF66nj1vYfltcafYb4r76FQnksRIAy9bnqUdQUxzbhGAO5xNq+K2cbFy6JOby1oGdCBm4/
vQQVkyR9aGN9uPzsKnpiEQz8SKrbyHk2II2Yl1IUg/Hu2nDJ4w8I5GREL58mWK4S0fjC3hXh+bb+
H/2yHtiLBugKpzeHA8Hzjm7LU8e4XodydMLk0VV+TWBvWrq6m02UkLK9HXHfRZDkWiS00fMo+JFF
4ix10yr2DbMg3FiKELapU3cjIqTYPjLnHrDyq/uGLxdPZCFwC7HxlEVGQ8jx/OrAxG52oqiftl+l
vXg6Ka1yPMTBAenpdnZ+gBQB1FKdufGoEhPUgwz3asVHnWj4lBcBgNlpvt0QkvtTOAGxNBIUo5T3
Hn4Rp6LjjFxTGGqOiRepHQk1r0eWZd0NAcZ8zZigpZGVzxZAZHe3PxaSot4zAUkj3jAobmpDWJgX
kMAOecxrpoe6wkcBoj75JD2o0tUR8ppxTJ4v+LHmmg+k+S1KJndmYTltIDJqTiIlFb0CPNN4Erov
Vxqv5PVQTvED9DYu+P0wXZM02W4TL211eGHU88b5Z53+vsCEMZV1l1rTibOY85Y5qHwsajrccx38
maXSJvxtLL5aCMp7LBxEO7Pvii87d6RQ+RNWtN7ktvkJfX2M4Hkr3BV7jda5m6ldInNpYcRrdKQO
Tkz1NKEljLWuPZjJvfUQOVf9mwqfqEXvdlnDTHLHl/B89xPWnN+CSl/XFEOGfjbSuZEqGxf9mr7Z
SM3n0cKVQD1OGsuSSaePsdIEQh+w3XOvbMZEXpDaDL5aaJliAHDrdox9AiGyOqy0PGqmIkRYPZpW
+Tl4KX7pR5qm8vwVFEnVYmq6kqlktuNTd9dadpuX+I4WZ+qinp5b0favo/K8Yrb9Q4ataE3Zk7yv
lEqt8J+z0N0qy4YXGH9uJVCL3V9aiP8oDRbsAqsp6y5id8tiy8fgUrlCcdV4oEfwfwdD2BOFDsj7
sTTEWpHWzjGEudCPgzH1u+KJGQ4tYBzz7VaPBgu2tt5UUtM2Vkt4H5nEdca+occ7p+mDfpcZomKD
zoQml5OY+JwwLP9uvl0r5/ViBKggxlpp3Qh9yh3l8E6zS5xImuUBqD7pkmPsYAfXo3C3Q2R7pQsX
17v5yvlyTlNpj9/BGmleHH6drLutNdx/64hfFulfqBxsrJ+suk7iS2hTFLEd3Rz031MpQB9JhEQM
Vc0VuS6oDnMRzxTLrhbf1JPwn8/IhZUu3CJBfkkX1ZRKcXOa8NwZye+fDDuc8JcNGwOC9yPZoNuy
WsQd/Ge9lDjIPXSvvwuYzRDs9gZweOrXbfnGBi2s9Ed50NIoN1VYlVNAMKlSVgbwZSqeCNh3NPwN
f+Q32GKj3qs1nIvqKuvJINtPRj8DnYgA4othMefX6O2Wt12fJ1lW9Ul3Ub+lClUc0v8wxH83fJpy
m/M5FIuYAV/cnlP1N87IYygBP4o2lIuX8mX+i72JSobHLrtuGeledHLemhtwaCUGwCTg7FvQzgkE
gtsyM090QK9fMRbSMV1Sfye3z9VpHm/ft2UUKNGfw5cHUFNks0mE7HEGkgN6HGjtpB84pfj9cPOH
VS4NMZ9N3TK1eGaUkBuPrWM1TZEURHtqYA707XtQc7lmXvTXz6aWJf8lWgwH/BgBrSrMRPR+QQjf
0T7DoprWr056oHUGUWfDz6u48rJtzP0O0swGK8gmYB5LvhaU3wc+F+r6k2NUPM+kJFYULBN7gHs6
wnhyvMkLwml3796iuurdOb49qZiN0LEfUu6AMiZQBTDHBL6VmeRsvY5jYqOXCODr59bDd2Tg4Gnq
KIxwd0EEoEo1sDbHkHtQUSlhK4SusTLBxztN+/26VhvteTiHiEGEt3jzbj55QNs0umFme05tcLqc
cFF97gSk5TJ6shGbETGCe7PPSR0hxVZbB/rPqPHYuR/QaHOoU58MGD5fekXS+9M/5cXrlir89qTN
cpd12pHsyeaiECaXjnOmOVgSHaimPJCevqOJW4PRZ4nCENMxp4uxUdXLX44gGgNUrsz9l4bw+eez
yHStGqlI2+qQF4ldZcNE/PVrFWiw8en7luDLl3XoKU1qeUb75tjkL81SaCN8mje8uyRMe9FYfge6
16W6D7qPTuKyNhHbP7Yee2v++1YL505tq0yB5WEWxk2zW9DqdR5pGS+68ssiOxX3bmAiIDrP4mu5
rlWJIR6eJ3vc2tXurt2Va2I3SC/YEVoEP8WTzv2IdZmh3pmzkNMUEC16mw15a9ZND2MUwVuaY1a9
GvLCh0JM/+QVfT3wHWFqHaUaMnNPDctiTnURWiPn74zSpF/CmIyI8cNiAe5eBP/ZuP4EUqly9TEL
k4EMZKOXTI2/YsyH3qRrsEc5AFeI9XPg0KUW99gyg6S4rUihSKSXALDscWfyYqQ5IZL8SBwd+gZe
hRIMW8mY8TeiXUbKyoCx1Q4t3uxtGLiZxKGfRssUtnDq7P6XNTmHD//Cex9KLWymLDb9khrSo8jK
WepFcfceT9UFW1yzU+lFfu1QG7qFj8G833XlR1vRRZ5iHOXNxvCqBLsVFoxpccERl9Av/VOzTujo
z1A2tEQjd/1JEB0MHgECxCwK2AUTzvWmiHflN7PoQdsQLEijWSis8yd8XxAGrGEbJpW0AyYzH5gL
5QmGpKPmkulIPnG03sNv+Nrylk7bT7tn6fSwp9x0mCqjmU1Np4P6SXyove/Wj5CurxaasqqpoKvY
UW9rFNUukGJKL0F0t0xd8BkkTOrrLJkAkBrWk/ULN1m4mBJZXiSBnz8aZj+gomCqpXVjRjEgc3mr
iqgjq/K1lPq+48N72VX5ZxGPGIg+eTHyFEHMU6Ag5hsv1kCFNMkNcjYvGY5f7vx6fcYBh2szYkBn
XIcKGKnyC3tanjLrrr7CtGN1V/qog0IxrbWqqhf2rNNv9TsoHdYrVp09pLlCrwVLlzh0Wy6DJZqq
peZapwKvUkg4zwM62nsGFAQjzUePiUx+V8nv1dVaCM6NV9ervWNrK1u9V8EWkB+9+WkuNwbsd59M
IxvzIpHJZpNxY3mOWZjhNivkhweR86KtfbRS7JhwrjuCMINdw8UfQS6GU40IGuI6Fz+PyWSI1sr+
nDVTLrbdbNY6VFVJziI2O+Cv0nrAjJG0B4qqLjhn5ZR9IJO56TP1xJmMwJgvjjFyt8jkzhLtjcJ6
5vusSH3wgSbW3v0cq+CEQhCS6aFLRqQ+hhsUY1rNF1ztRqc1bmstzHN58PKZPKD+pTEK5tpP3amu
kwwvNT34tGtGWKN9uduWoMpVZ5409LCapQ8BEutjUcTiheq3hGhS/cO+QSDUdYf47KTWj5gqLlhk
ya0dBrdTx9OnFkJtSkVXUkxpFLn9gbLnx1xIgYl36iv3Bk9q9o01+4FuUcWlEa54U0OxI/sEu6p+
GR+B35wHv6c2lqTd5clw2VO/SXPf8p9ny6cvIE9yvzNh3SrZ50i2sVFolm8TyQb5702VKJRmEBuw
Oy7i+FoHNNBJppeVMgz47F4v3GFeWqLCowVJStZdnYpoVg2a0se+SxP8rsbIiDp8jTgbPYFiwNvr
BSMOu1+uExzMezQFUsghDCrx/G14KVOd7lbLUPki64p3RhC1flzWjwxqrmEGcy7tubTgGtkK7Vhw
02hCHeQt7m+Hco5vZTIOIJXQIi7HlRC15PlKnnmnZUaI9HC3Ij102bbBTYRNlA1Gkmpkk184VgD4
E68oUcfXqTjkcGU+0m42EAztw5KPBAjVYtGG7mlDTkF0N5D8p+KFkwiOUb4AadrJ3TYKF1jx1488
TucYc77G72t7YnPSjM03dfXRcjrji5WHuOhqIM9BULNFDzNu3rMH4Sazq7aW9jf+VuFu9olx0zbC
x1BX/guTA5UhJioYYUrp8M4hhj0psvnLsldRiDIy3tFirxceuupwMuL70BM1OU/tet4uCd/kwj6c
l5ZnDAgXQRX6jNe8lKkxwZL1lnI0DNZaJ3ZC6vz5xVVfUI2RALuJCrpX+2oFqOov0AX7Se/jfBVG
pt/Se3KysxXneuo/WzbEGRybf12A1e/uf1Km79CikUnLyoVWkH/CAW3XtY0fS1ccrKkI30dAmuwG
w0Up1Vc+NVK3q5pDbSaMQAoul5j02oO98HvZ4ZmIqAskrqAICWNDVwVX4IxG2kD/I3fXeh315oEX
qhU1AZpYqQwBkQsBEdYz/3xphL0SDYi1/mQABtDrSL+L2er3MgYj5U23+boeNRPnSqP9RAQBSaYR
4Zn24DCZwVsbNFo00dZQK5gZ2Xnz6YiBHNnA6QhBcaFYHmxfT8EKe4rkadlJdzUBhUWEYIpAIjyc
em+8eBr5dKptH2Se75zVzUNu4FvLV72rcyVwB9LNsBSAc2qoqnwjYThdVI2f8lat3eHKIDjcjSXf
ssnarcxW6+Zv+HGexdw9QmScp/xJBg4k6P12ZSoJemhjqxdar9piTQr6VSst6MQfIMOkYbIMQNcI
vPX/q8FtEke9girGcvi6yQywVESUw8Qe0Zw41zj0rSfS10k6AgcxiVEvWTTYl67zcv5meekCHtKm
oMnca4uoP+7B/tQljggO4/jP0Cs+H6byjDvIGMdEuRG+WIh5+HB3aYStymbWb07aqulhwQWjMxu4
cMJEM6hTG/xnakyN7GYuphFqcytJZMfwbnkArs7Ca4MxWrJkw72Nak7bIl+qiqlA3fQ7fffEJCp5
oS9qa/gRTHNtuZLDhQtLiG24hSQwMYadvW51eOkC8ksrJf3S3btH1lZM59wt+xv9lkKeEJ8SIwAt
epnG/cd2GJOQCkQx54Ky6JLnJoqGfk6i+wQo3mQTQjxldFENYpvJyVpqYYtDtXIG4+4e24D7or40
xhRYe403TP/b/oLMS17b8B/UBMSg5hwcQwCyaRChDEWOaNMwWe2NJT/nnMPAW05thmaVrVz3gtcL
RaWaTbyBZVV0HPJBrvTm6qNoVas4Fqzb6g7A3znDX/ROQUoTUF5K+2jmCQW2EQidwbRBZ3HNejYb
EK/f5TCW2pcW13enkiC8l92wIg1O+32v8QL3beteuHIy2UttYgBHhSxK1TLTlDJ3ENgbn5wmnXlJ
f5IhDUfaZXxrNvmFsbTQ3ZlWZNR6kcA76VjVViSMGveLqzP/OVl8Ok12izt2i/0jGyb5ksimm7W/
GaA2pHYnzzMIA471GdVi61pu1RIFf2tTAjJM28Bpvu8lTaHgUmLXnCS224dNlW0cOPTHXqOSY1Mh
3/MvNGY+Pa5TJ+r9jfUu5N4Ix6aSXYf1KTmq4N9Etl+l82fmOSJysiBcU9oWGmRl9JjkddL/UB/A
Z6/tOQaAsREN5oZQVavui9ssPyEQFEwyM+oB4AUXad4kYd4jZ8KycMoj2haUxCJM4BJVyAq7aUpr
tv0kdlNJDjuzVnfkTHNZrKszMMFZqKzXqT2GPZx8IJRXKEYb5IKZrTIQNAv9FpAs4Cu3RgFV01Ll
cVeqx7tFbb5v69DB5pDE2ni+nYAfAaB6KhUvU93hnGbfz/Ahqy5LzgWVGmMzHGM9jftfd2jHksZ7
Vg3tLTb/MuVBp+Bo5yDPNbZL/VFHs/6iVYs1tqrnf1YmoaudwG/UmQMtcMY8oXVl292sYCb0iIod
XGu/w+gCgmqyGbNyoy2z0PkfzvxyHlEdGFX2aeHdOm/GEXtn4p/HgqjbtKUXPzYLANN8HmWqcCzK
tgOoBL/ZcvWuuYx8IChz02mb4eEBdoN/C2qFvMpic1vUsAfltwpf2cw5o2zp1d4ik1/jcgi1y4Lg
7oOJSOCoQ96ox4dBx7X8YiB9uroEWTBu/H5VgW6RCOhTmftBtaLO4GNyJs85y9q0Dk0LrC+MTyvo
pfCMjV7pNDpa/s/n+eHjDPa0NNU74haRF0/XPwpvKoTFBsmI1R7PHaF7xj51D0whXY/hZSP96F3T
DiiYy/VzukgZNaRUbUtGrhH+o0k+vyGL3V5VKOtSy8JphfqM/UvaqZIB+1T00lRBA5PGshvjTmPm
9z/7gjN9S0jq8p72iR6csa3gLe0D3tVMYksj2mt3cZOGK0nfQv9kRFmWsPjyYLrSTdWZITgcYXzE
c/ECxhtoW8hxs7iak08aNu4e5MFE9B7nXBHtKnDMgKVKwgisYr/O/g9tTXdsFMEB3v/cS0Tdk4sB
xUV5lRIvxm5wgaAngM+UzOKhUl90j+vqeW/SiWnlvImQSq1GyIgPY859WOMsRExeX1pA9v1ZQtbP
hhpJo19ksrbIvnBcMVV+NWyqD4vhNU1V5w7CqkYKunjryuvxLWXfNJhxXX0tEkPT7P8GxRl5SS7W
li+11XytTm1qISUiQvB5Rudbfs0tMmCj2vZsevBQtPYqsGxhvSQWpvXRxmKY8pCSXBQ8gCJv1jCq
NNTNJdIUnUOqdFQBmTnfBArkP7PRo8UkCQjxdDMBXpeE9hvGC6OAezRbyAPZWlJbkfcdSxAFf5K3
H7b663/syno3qe/89kYTFNJ3nU+Da4sVHFD4XawdjKaxK+kufpY9BcYn+g4kTHppyNvZRjDxT4VY
aR8Zdb8MpOA8HWgx268PifY88OV6NSEmNxJu0ArNhYNrB0B4TvBM/YUyDvOCe3jiIRECeCRaNrWH
QbUeksxG5KVpRrO+rWmVreUoco0fbOhV5i40ZkgqlaZe9smG85CDk1iIxBYu9//dznWuPABT601v
i1uAgsk+EH+TfL65ILsa24Sjsu6DMTpLWBhkc09FXkTByKgujkp6jOcUGgpW2+qb5N13nY4fCYp4
5tI3pAwmWnmRoNKE19XHsGgFWdi6dLvF/3ay2ZJFWTUY0WVRUTnFujCmauf+l/WJr7a6BGC3fzwb
EtS4dulI2bio8q7iQOD+7zuUjbiHzHDxOioosqgmWB/fm4WPKB053zULWogdNzLUpDkRPCdpcH7E
wNC7TKNQOhv0XAugNx/VqKaJgqh/aahcGnVikdC8b+FmTXXTzgFDHhbL0VfrDDHT6ifVBug/CnWu
4EjHDwvp4EklPm7k9vk94UiAC0+Is3HhX8dQb6nSzhIZNLXeuB1PJeYPY2U0Hppi2WOubmmCY5wJ
jkRC9R2yzaTDKSrtIQoKVPCQ93fkJFgCfdrSDv+29O1EPPKj1D4M6bhmDLz4uWY/IXgfHPKvRxc7
chlhAWyFSA+PY3s5jGMGgQOddMr2QQ83OpMAtDm/jEU9CE1kSGpmlCpQZTodbsF3pecFopnvmLRj
NUAj3ua/Bzn9o3y8bYoc5vBc8BKStlY9IQrvHd5F4TYWaUn91CzU3B1/6l94x7QmrDBh1fjUsCko
Ul6od3L/hRl+DruWT0MmrHRME8faJL4aeIr24kIaUfpi1qNcn86XaTX6q2UqOKaH6Y0EG77xN2o+
QKtOVKJY/Br65Cqwk/YFpIvX3rmq+eL6Z8SfAZ1MDhmIsaI4tiZHIO6mnvAJsn5bZ92Sj1bsGkiX
rI0OfMQkRZffxg/1zchGNAqs9jvkHSLUUZkbEXN4hTVc71fXxePIKWr+KTE27gOofJwAJWaxLxhl
c1ZaKq22WX37IXBeRHsEYoOS5f4tsjszbifqAgBjswwmrix2BevyZAk8XW2rv+ngZSR9Ys1mDZE5
q5Lcu5X+J37dF+KSQJiRpr15eKq4UJyBA6lAvo6IKwBCzwsLk5o9K9VVlb9dr4BvuVli7A2OcaWy
kZoeUY/H811eIy7W69KdqjXk19fFvbn04LRdJNClo++3Hs7R0Fhi4/EZxrydRpB5s/6X4uyMJ7cA
ukdrGQ2HF+BkM66CSkrkWsUzc6uDTKZqb3TlKVVYberbR2qh3O1Zwrmm+8NYW6xPnyF7D29yJyQM
JodjZkPY0GznHe54+5Lfqcr/UE4GdERx7hNgVTOUAQfWb/qnd/eUEUpkszOh8u5o5W6M6lUqKOAH
9Lwwa/h92Sp+yfyaWJ4V167qiH9tVgZfmXUoAWvbiW62JzVQKsFhGKrPbxX/N1M531q1qoUSjFtH
/KMPjHd4vhtA3UW2vHWNk3avlL1oLzhXTwABppXWLQryfjBiIbqMynAJrGtofXSmmRepPH6fMg99
aVTRS3+KLnBSTbd0FB5qq19iW8LYtUJri8r2Kjka2eUI1174c+Lo+61mewCDh6A++01/mLiqDL/c
AZaHqn1K16V14pemD6VCUK0niDdo1iizWTEGEri/vchumuTHMktqwSEDrkXCLuWgfkZZ+UZEORS0
MIctNQY7HdYCOppSWDBAJ31MiuNFFGtqDT4EHvBI2PNfFvivB7iV+I5FgIokEZLpn1QtFQRHfgut
CLJHVHzMNtdvBhboHP0kBmbuZbIzWlmP8V02UOhY3wPYXZqPEFB5l1Q1BGZ3SdiCoSq1R0YAHm4R
HEAMrj1c/1hpPQjMHTmc/jepbZzLiswKx4Ppw/2PVryLw8sVj41Kj3vZ91KVfeFPpP/nQh9yOrlS
fOZuZ6BMYoanqqLFZwfhCbU3bg7ucchsONG6Bj/mHZiQ0qRStOZrf+PEu2oxtlvk4ZuBIQuMaK6C
WkOO60ZWvlkYdrtZxQWnBfpkdBn4KV+2KDgouOU12HV5xDLBDDLwZpiV7cVRVVHfGGX8vGBTMZBM
ycgI9Cxc5S8XpJS3gGxn8hEM16A6wQ2PR+wfqXrbHad82oQeTWbNcjIl1PwLcbrA9zAmwecJ6LKb
RgvkiRE25G0TgRaK9EDFMQpSotF4faQFXxOxCo2bj3ZiwZUETa1i64ldNC4uLHfCMB52Pt1YffYI
cP65OotVx7dOIystHAebdsFXuC0uyQMAJPZtfo0wJFtJzR3fjlEjLhVsmjHdHR188ue3Eoy2zeYP
2ud9tbhbxapH8qcOOEMFY9y1bzi32iJr9AU6m6qAvA6z3sTc7PEgH2qqrArFNWw2ZAFSF89Oavzp
wm2XIrYW3OL9JxpF3tNuQqbrfDLILtEAU71lUQKc7ZzirRLReJ2LUapl2wOwGrcwX+tmkkYASi/t
ZSooQmPvVu3q6gZBWN5RHQ6BYKD7I8e51r85et+ADCJdl/nGvCV/VUfaLC74Yb8mUBkzTt4oezEt
3/hb7qWN6T/quKQ1goC0yv+QcwTGIFgyHaxzBCa3D0Ad3Pv1Jz6Jj/9U4jLRTXsmEgZD6ePgUW/7
FlgL1cGolKF8XomL63B9FMecr3uqtIhu/7YCXOjlPp+cPKVHdGFW3xz2jG/gSnsvNWi3dfu4Y4zO
HDD8qq6cw1AjtRncv6TvmuMtV5mDWIF56NHfVCKqEHfUup96jJ394T5hmlsOpACzaVV4lAFB1v35
u663qvoxfbwDZZNUmB30wlkuD0/2A7aG0eUBM0r8wdUu92ei2x5hs79do1yVkMy8EtwmUBxDnqd6
J4fjvGz0MHk+omW9gjhFKoEmzf+fMMa+O4SDpHuq4MQS/0WdrEJwLyHIRxy23AXOL19tIJkOyy+3
cA6UK3QrKQ7h5lYqTx3DMv2mDpp2u9luJDBwoWb58EFJW5OTDVhgvHPa9W12o/yxi85/F3Q3Kesr
LeMSllVQxwFqkxuyyjz+JGhSwmwH1oM8ZqD19bAPIVKsuWx9iym/UkaptkJcbZz6y7r6mNk+Ja/z
ggc/COvh8gZS8Z+Ln2/S2kjAHr/oq5GvsO6C0kCU5ryMPMVTZmGE+vT2JbTyjEnGbEgVfFhFxE+7
NYQzs9YOejlMqg4Zyh4apsD2xijdBx6AR7M7hccGwpp0bGaGWDmjl60TAMJRJGras8yyQzVQNkYQ
ptBa9pElBCIDJ6Vo45CtgDyTtKG8n6lfaWhBtWCX6RoxmLzskyvrabM5vLCuqOGMtEq6Nta1n1f/
jiqijXZ+T4K+wq7iXSQ69/yhsZYlvmVfFXwh9sv6gmwUXgBniqBJkPtE9nkL1L/4exdKYYywJRmo
j/Wf9PCUGhAshkPNhqRvahhLpSlc+H0mqoc+sBBBuBW+OofxbkS7/uhpI8U34rBSXx0D0j5Ngf4i
H+5ZeYaKB5RdrnI11MO3euYNPIhn5B3p2ihd70lHZVsehvCQU4l+7CAWLlRiSrxnNF1AqqdqKKZ+
DMi0mcFfGX4L0PhhJ/NZYTsugdAkqG9HgFwHJnmNMLNijQhjReHFFrOnXTchGRknCd5r0Nk6eVqV
PA96EHwxH1FZ+eBYOKEVUo+ULs/d6Q0bk+V7+Z2u9ycefuy4qfpW3UrTXV/RfqVyO77bj5tDN6Vp
hh3v3I9oYSjh2FlUs2b6fLgrIHj2fp2NAvjsM1A7LOoLXdhA8/8KzMnjk9ZgbngDn9VoKma9ahIP
mNE5bmi4mSe2KBUx5e91x/uGcYBrYcIxksZOIl9SN07ga1k0JU7GFAnhxxSwuhK5kpxN0zFwJE92
lNBle7TIazKdn8fMjIyYkZkfN3ay4M6s+Lbtg00mwvG9/QAR2XtuLFVRYK080C0P7VRZWzqFvZKo
XURLYpt9u8qaFYNJ7sOcxTzLPDW6RA66u2wDsBtQxsR0tlJfuluM7GsUqdb1mHpeTdPZdl/peZnv
fyun3Zel0KU/Czd5liFTZlC7cUGPdpAofyh1UHQw4ldmk6kT4QWwRQUjxLR/TeIo0EJk323GMWCA
4R7jVP5Sya4+Y0zPZK3tT90QTaMAxI07IZvxL605mfThJtilwrSenSLB4EQYYGWCELdceELP+BGx
NkQIMC2fEf2GzPCgAMT0fVRH73pwbyKZTcFM6YrXHlxNRZWXJzuTy+H+YTPtM885NJu8UiANq2X9
TaLv40jDyjS3A8iKHCQRsBdlVWHcI6WR6ll9sWH9a1HywnllUeDhIn1gTiVflE5LlIB4ZgK9XcAZ
qPvbIoWp1cDbQ6lk7RMEtljkQBETfB8o2QfdaTM0lvlTMIjAnQQVVfXBMa3orBlPtF5rgSVvm+19
jP1EBNtURtf040L754lVK69+VYMZb0+jOPQKas41Cv7lDT3ddNz/f/oOb1yYw1rYoW3kMcegoysE
xRQ0aYDio/3E1rScgIKdqCz117Ev84wm2tnMDzW1PFPTfdafYG+NFYgrEpCcrEGBekCUsH08hsmF
Yq4/VrSZALlF82Oq/QKJEpokkskrn8x9eM/4ntx2L1i7WjsaEfbyW9zhLc/62E65wKnIJBtnUsRX
JRibcEmbGY9Z59avaiVx5hmGJ0Oo9Sjdp69YcJVCxJ9cn6ds3XHwy4Sm4G1nT43mW3ndTt5VWbJG
Tx27SwKNaZcsT14Urz+OM/a0GkJozHmOQ2cLhmFZcXQ9zYzE/UJeMQvpn84EQ/WyD7BcTp1Wekz2
k4usg6LHAAZ9KGE72BstXKDGzgXQDfxVvRlMOoRRa7roM4h5Rr5GqbKpzJyUUCnlAoOCSp2c9ijV
NLtCXogpRhlSAOkLoLqi0GBqS1OVZeDeKD7Wk6lugJNx64n7eA96bwwOmNQDEjHp5sAKk/yPYMDC
8X2TURWLFYZdctuZepOvv3LaNxcVKSvfJMLbg7rNN06mTAliuepuEbkrniyBbkAKlYdX+JOLVdWe
7KZg12b/nPA0Qkrus3vV9hYX3Ml8lrH0nVL1NhT68UF7hDYq5PRxFW61jo9NjRysfOC5P/TYPyoD
IOfHGjJD8EOi0BQ9K3Dfm039oTMTk5NcoqGzyqFJkdilDs2/vl5SL/o/cC6Lw+bUcEyw0v9QrdNp
DmFoauzlP/aisTSdUuOx5tLTHYYBuTJw64cb490CsZW+4F1R5JwIqccVqRel17kcqfl77CSptA==
`protect end_protected
