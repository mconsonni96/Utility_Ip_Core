`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
QASMEgZPoFgeh0GYz6O4a9m2i/FOuk1bf3Gg5N3BmLNaJXWNn8kq52c8th62Oz6G293icHaO10UC
V0xIKwjWNVUaxu6G+YcV6fu+OVvlvTWG1902WNyLg543RtK2uhXn8SJnf0IW8E9nE2Jt4Sr8X2z9
36EHbhy/9QGSI3PslnArv6X8OwTql4jtYs2N6r1cqBYESfRD24BRdO8oLAMazSQYGHgWHxR30+GO
1cBi9DTR5B9k0u0D/QygxAhAyr9Bi/qlwnmCP0w21i1iM9wCre3u9UiwikNBTCh36/ujAqwXZLP8
ufxdHoO7T5MplI+MUkyUfNJpoUITXqdEMSs6zw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="+8Ros6SZIIf5y0vPppOik5t75/tSeqZOIqP6wIhF0fU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20656)
`protect data_block
Vlp3YHawScSm+ve7zjuP03sDVCjjvJvGQmdYZJgMAQlTbZZRp2ZRz535PEM94wpqzyNowxv2MmIl
NVg2sLawyVtgVlT3n4rjwB+bHBsX9SCH9oPPyLPvow78P1FGNXvNFoh57e6qgHOanOyRh9dMbmbD
M78j8EQtoOiL8a6Wpmh87EmAf6lP6cE7iSpP4zS9a9qiVpM0nzITtWh2bqjbT2vEWHMUx/IB+aBr
7EC6JlbxsI5e9j6O8hC4+AziD3/Ps9q/iflHueD7nfX5tLQXqlq9HMZHDQN+x4tJoFEGzNHJv13D
pPiitaYTnRWZ5NVhbYBLOmRUY6ZLR+ugqHfNfkzUF4SgeQxl3rEjKzdZXpqYVUNTCUxVT2YT11MC
Nv6hvlE/RHcOZ9lVT6Xp0D8sxrOvGuBJMiaw9FeWhGak+KMQzZpicfjHilm55s3flkrW21LLc0tQ
GXl0Z9VYRkrqEjZCTWXFcR3Pv/5rQ+r4n9LhuIPNIEQQh6Y59egskQvPWbmKAevSDmiwXtvaxHXP
rYNhmbwKpYmROc5hs9wD61FahlSrbbDZt+g/UoVX4gpMWrmKXneQkwmRY+7WObW4nsP7LwFGYL53
c2IX0OC093kM6CFbYxyH+ZEdl2qKUhc+27igO6zjPWkQitglhCQnhrYdKw+Q/aJHoRRtSamUSutC
q5ddVerYDAuXKB1QQdJUvAc4+vH7HCLAazfU6vLdX/fJ5eMJGMDACeZdXnY5MG1hr0KoOQOvWjjB
rCORloUUF02SxTIy2evE+IB7FgOVEwiRE2XNYPgrGQvg4MF+uFyKpSFmBJk/6V3vQ89hcJ63PC22
pAWEZYAYooJRPtOE73vM09g3N8YQ/cLqEsvsWGtafbNEFDZ5qvSiPDHRyxA7dRyxZLt9ekixqpdS
RShDyjiblr8xi378jACgzLLIG4QdEAdZ7aU3p9KdKPyiZFVop6Nnfb2T+AZL5wyZ9R7bxPdEBxTQ
gOFyjDUiMcwgBoqAZW9zSt1BUAU8HVwLQKg5w+M7HhwikzX3z9J7tHilebNUcuXzQ0p5opkYvU10
FxFiRVg3wMmlxcebpifPNHyzBFP2PdIGVVE4wpHc07vLRhqPUdnHLhRy428k321IhcgFprcAXJz8
+ZRdlT3pIdjOSgJhuUSiFtoQ3/fKkk8eNabrd+ByCW8hd6Z/PD2lnBLvjyUmopSOK1fINO7nHUhd
Plhq+XrX43md+4eUuF1XUk9k9cq/cAoI4VjXHfW66Pn0QcxdirneMiKgaiptsen8NsOhKbZa/3yt
WfBcDKhR+PCpPK2fzta0GUM/NQTvBibW/Jq20yJoYzUO1Q1EoENd8j/n24Rp7hk+k9Ef8boG+lNU
lkdiW4dAYQIq075ZvlHJBwH09rFOiV4wjD2yzAwBaYmfVlG67YV22Imaa2mlJnP46kkrI2Uv9WNX
/++R2COP1pqXOWFYg8uuonn0+eCwxT+4e7pQ6891WxDLo22729b43Y9YRvbwi2H9OEDEHFhWsudR
yKkIvFal0lfMOkFP3drKyF47p0NSRpOtwfmKSH/quTZssUWUlAYsvnB4OJ9L8GubGh3Iu95SkWLt
+y4KviqLwVzeB4pOx+IUZz4F/Iew5KgHd9vmjfBsvGculVXHYAVZEJuzzpBM/utvZnsHiVUAQecw
pOzXkQ7bRd7ujRtPMoyV7WhMlCzkZtN6ClJR/7CsdT5HyGNc3U+9sEKg/0krmvEd9ZexgYLue4Xz
Hs7QVAhdxOn55pfCznji8jQ2sG1XPskIsIErNt+Dxm0a025G/PuUqZM44vus049dKRmiTuut95Ry
8YXgt7wgTegqvg55pQdTcUiM+hk187czdPwpGl4tigvUSd2kEUTIASZQ2UIMd5kau1DA3vL3BA6K
Ytsa7YjfaIu2cFWZe7Vv71KzPw/79P5SdDz4E8+OZZTxkg70xtSI8oee57LCJDE/4dpbGh8V7gxk
3W1W4aZh+7guy75TeDk66ZsxldoAFjGhXndxJH2UPnGpnSa8+Xk9pCQxiM8j/tR375Ng/xnnsj+f
fJHE8/zheZYfrO29HmhzlB7kiyT9lbbVk9ZMLyixGE6PdOR7mldkrEc3qlgrXb7CqZ5B30dx0Ma6
VT11VfzlifrK5Wfeqq/+Wmfqk9bzIRAFhZkugoktWfL2TIu7iPMlX2N6SMoC2t2PBGGlm4TpJGod
BOzKrWw/7xl7naKNQqPQ970atVeT61FHKQNwI09INXQondaf4OZqtXjjVbtFuyEEyWGjgGSFyVPZ
ErmpftMSo2ESx0bhqbRcCsYX7haWpnzz6C6i+Z4QZWQTgWHb6+hyNnSNZvVEJ8oOHjaQgKpebTVR
XdpSr/agiZIAfyKLBxqy/Gcgs/qr8DMFZkxNkcGRWQUd1flatCRnQWVp1+E4XNmjN50SZhR1xYtP
rwkwC3/OmtCkFUcLC3QSwmmA9jrOdFVGreRO1zz7VekyouCq0XVjbKjBppVQ+7RWTrHhpJfrmLGU
UvZ2Gn1FXK6132WI3YJw27ESDDDHjdvNn8BnlwWdeaiNoE84Wv3qrO5kOjRG1vvA16LvxodVy4pb
gACWztSdNPIdhiijiUtpLJTZJzLUieq4ALw8STBWvzSSkjWt+HB7EeMUncQZvRBouXxFvSn2eIde
/Imux7z4yWNBkSOjdD6PcYzrBi+oUKYLDaUICJI0ecDVCNGivQPy4Sx0q3XvaZ15F6YC1x1ZwsC4
lXI3cHcnt87acob+Qk24Fo3CI6ICu6TL67HNqw7MXbBXEBWPgJDpUvYY5MIo1eg1xAnoo8eLOf5Q
2moj7Cxt6wnHgYK0DwA/6CA5YciekR8VQAKVuVv1uZcoxykG+QthnPNThOtQpvijqQP1nAxsJw24
IOs5FGZID4O2MJt+l+nxxIwweVj/kpVmEWm0hjdaLJPdj9NeVIypBwKe6nYGi8pjtEkDpFODLbAP
d95h7cpgbRtGPlMMaAzwk6yyXSHORcRmiIf3NKcNTjnG93M56czfbzhOa9lWMk827J5LaeDH5bEU
HhPb1c6/5n2gdpEee2CUI4hx+PWTk5PNT4N9STk3RYa8H2mtrwC6DjiJexg/9C+B5ANsrQ8xwyu3
+j2n+EKKRJTq10ImiHkbuwM8ELvWd4uEWwgIiKiZI74dsuFNixLgJto65Dcg5GSVnG+jLQp9QAUp
LThJ0JUiySk8VEsAwAcM/QcVFEHBnUf3QME6Q0Ch+v0ARDhe4bUlXbBG0/gTLLRl94Qhp3WOrPmK
AfVfIJhxSKracQromBmCpbbmvV0+4x6BvSms+WCWU7G/uS+ZMroisXoSUYrdizG4ubks4ZibgyM2
elGuSVjdMBGblKiGUUP5wgs0tZK1nXw6bceA6P96bdGgUDEiAy6bnwWNTi8q2ykvS8hF9ugPjcps
r73hsyYe6+CbU7A9qhIUSl3VfF+ef6oaep2GwEt9hkItIbaRI5+MYzPAsAbuLZSo9ZGUHtyp2yLg
zBPSizVw51JgUvsYA6x8AVjzOjAjuA+MhkQ84V94fXR++cWEyn5yGvj1RDiPMytvGJxVJYO5/G7c
lNTVZP9TTTpflpHclu48piZOE6vU+iy9DbOtInmc2moeq7KtT9SbaPrNWxpeRfIqWf95263kGsjw
I0xn82rufM8b22WoHKi4vrT8ScUixq6YxVVhYFHK0HgDtD2TSKTwYVvXdPbwXnzPEC3j6X5wbxLx
4yoJsdQXFTADpYG9ojoy/GNq1icryj1tUhw4qbvARgxCQFRbe2t+N9Zb1LJ0GusZbi7YDRv6N8Zt
AgtCHrN0HZN11ERpXVRz0M74trqZwbwF2EcVLJ4pMkaZfYZ1QXMzeSc51+A4jDvFkT9/s0BL87Vc
EdhZzMdZNirxKs6GoJeRnEaWvc2GsAJmdwefXwtv/7SRGEkJ8xDZTWppZX8hWI+r1LsbqjPqeqsq
vFinZnF0kgauWl08SDGt1aePTQezuBx1eQDwYui+rnqj25Je04yrMCw1bVvL3ARpGem2eKBtfZCJ
Oo7w8AuuIbmWVj39HieiHZII+JNVCk2ynPQWgzChGxDiPMKn5lnHSFtNnR+NIt8Io+NU7qBTYgKq
0ttivszIGJ8rRSDXz9U2GeEpzltTpTYijzYNQjP4ZKHVQS3EVmY9U2ORrLEN4wTfwidIpIv55bNf
U92zIEgmTJkbpOZzvL+44fX0fablwnfeVMTsovWp0woYK8JE0E9b8/gHYptBk++JZ3Q2E8cxW/v6
d2Or2dCjWb8f1QBrrApaGe+CJMsT1Ic854/5yGgZoeyixIh0mpfJ9oJLprayZ69cP+Oebbt8ZANw
XK/Nl8ffSRo9TzQ0uiU38FRV441j0JCIdkV6UdC0zsDNo7ZHdeieuG5JadmJa6/2ZuhYzuFV149m
isOBVMratGBBOfSnbw5GTWNYlM4ynr384kJfOe8B7iZdnRtiwYAwHoOlY3UcW9vFtVJ+NWtfoLvE
2PhgI4a7Eopfxu98bPIQDvnlkV8Mu0QQBddm5TRTzbbKJbRr+53jHsNHWH0mIAWV1StTUAeryh2k
s0j4A2dvzzYdD/q1LmbasssUc/WvAfNuBMvbZxGhsyf1y+HVuB8hYe94L8JiYPLh1idcZLw9xs72
DNSA5zXvK7U2w2oD3tJWS6pXF62crZLwUBHFomimelphaaW9A/y2L/2r32VL7RwCowjppVbZrmbi
Mn/WFxeVNkr4COmMSWKhsByI/n9AsdHwV3qLNcugyiJH9q0v9ruU4h3xkkxZMTOxE7Au2ZdJiezK
HzOmIMoxoVwqqqFQIKKx8V4BIlEBlGU96NynKSSm7kW2CwhH+ObfKJX2fUAJM+/Su5nC5LSUt+Ts
2PW/27/JkpVP3IdKNOBrIdXuw5XSGnXfvSa5PkQzq4qfu2DPedjLTIfquTyx87l6ZUChIMv90UJq
63ciA4gpRt1pdJO0FRCpYAN1WwYt6P2bSSxCi4HyCdZsn4G8xN624cR2DyytJzNLZWFbgB++p6rl
EefnYFW5i6A3eQF9dG8Qffye4EhtFuXAuCJ9/nkS5r4HOFYXxOmgaDlrRAIR28MWAKPxVhZqXCV8
+hbyDlJ6+51/jmWf/TyursLt9H6eA4PXuqhnfOG9nM7l3Thj/SjYizxHbt7/kqOrYuQHj4Jz+NDj
YXz0m4Tu7lqBYXV+ungyn47xOoDdMZcx4ZbKr31xpHNKuB/uER6Ul/hvKAIHUa9mQaMXDrv6GusD
mMS+d+8LuGmBFYi9IMbDzJ/8hqyr9WIhBvKimc+3VM3RY+yS5IfkS31mA+AV8Y3R4WnHbjHVVxJ4
ZJlunQjULpfs/XXHJHAdTNADk+gLfTAXlsb9f9X9bK9N9oemOdQVw7+RM5XPgXxU2ANDFp9JeOYx
zBUgS7z6qkchbwCc9jQN2GwEoseTTbKoXgbVPN6BVRDErWE+W5Kui8+Ofm0It4f71YvBd6ZI9V1H
zNOEddYgvXspYTBhqMGejZGwivt6x8GF3l5np8IK5rhlam8MnrZaXcpg+6N8kL9o7Iz9Az+Fi8cf
nDMBguGA6cTi2ej7NlnnPWqoFUFLHWxXbFDWnt+VtckzTcmZS0FnB304ZHfStpu47xmYS6CqpJMf
oVG6wkje+bYLfUMZOf5S4bcnjfUzVH2s69rM0kPEdTFO3vlRPHxf8iuALN14VC+4aA4AEppDQi8J
eKclUQrLsgnyZzGNEoCSBtqwmybi5duuvivZ4x4J6zkkVWdGTMrauggboT/YeRgqjgjDOtK5ljDh
eRABn1KEVJ9F1TxE50HvXQ+phad6kQD3iZd8W69DLnKIdcZbESGAl/lzqWGhPopvmCCVtj6fp66H
kB6Pi7gQtE/kkFoaFgMSYBMsOkDLCELHO9e0dmtn/NbB8CAEvEJiFASKjjC9VfY2TLIigh8sIixu
iGhAU8coJvrzfhPebcTTVvvmawVAnj4fHvA0NUWqaxzAG+BuqVHy1MIZVGlrHd/AvdhvbpKOcPJe
+WcPmEom66mXOQKufNZVU+D3kv5VPAOmR/MoL+yO8lvL4dnSt2eMPzWpuhMtUW9SddXXcUFuzPaD
JSsBdcP7HHw4xqiHfaTChSPgQOBA/VcBosG1X+eIJG/jfIuu0/SnwRaAEeBhYuE5UcmDY2i3xHxk
haBQE1xSd2lWN4tfGBIiRIWJaJZU1OmN9Bd+khZxTnALE+T/2iC8k2ebzMaAf+Jj0+AgZju7/awk
EWWoVo2vewhhTw0l8EVL6syfOmKT9ABfFouZou4Zq5P6wotlVST3P5oRNH6A9iB4DRhF5mjDzDcz
n50MSwRVumO12R7h9dpLYEuVqPItdnbc8Ht4K87Uj657V6PzaFFtuivHKXgZBltmzRn93mgMWNKY
8F1CXetOmMnMB/gTYZJ99lq4AJJ2R4C4yg736N7R/c9QzZpEkkwbrHIccfJfYL/kBog74se0Tq4N
vbDioXr+38ddxoganD54aBGxfNlFAiFVQ1HaFrG+ATEehScUKfT/6hVM32jQdV0Kv0pz07hfcned
0FQRc7zs6+66K4cFu0eUWp8+jHwPg85csbPD2m/IUlN/AD/I/wP/iEJgooom0lu5vBcFKaDYeKlE
6JBbvSPb5vCrpBi/7EwVzIebWp/vmz49TpmoVyL/IhsiHSKcEx1pqHP29aTb0w0bKCYQiQmEVTw6
T1IYcGeN41Trd4CG7VHqlIIvS98naR7SzE4J4jLyxhARwYnPRILb8vztZPs/98oLLd/jHd6sfRuB
/lObjr3mSzpirC9lw8zaIFkzmdWsygvPufBqaykJANFZtbTVmA2DWwj10A51aEgzznubsUhih1Lf
Ne43AgF4wQ9VwnWDhgVg8QPkINMydv5DpgHAaAR1tp9f//KZi6xTiY5x3Brool3ZWnkJgTGODwdj
atecakXy0+fA/6ijKNbGfZTeE0xrIWGvv4qDfFL+aoxBgxBimI4kV3SE3UAmpwZPrwlEVksY/dG2
0ky67KKtZ7IU/IE5Zl8eyNPAAP1MzF4ASqVuLU2jtte0T1JnzHVm+6pYceyCcT5/tsbDb3o4Iafk
TTROfpjvagrbz8kLFh7vlY1atUR9yPgkwD8yXy1Sqhr6z875z8YZpfL/SI74Abj+GqjvoqNx73VW
w2b6jLZ+XPrfPnS77sPOIY+5m66XBBhRNYZWRLpwfLeQxUxg/eYKEHimo/0u2nodY8f8tDVa0v8g
vIAIAvxP67zzrJkSjgfnRCIoQnGdf44cAzQpu0sd+A1b17B4mWWWGLk/gj9j3GYcbe6W9uSeRml7
sHAJfWMEqpRLcvns2HP65568u/qt2BOgwf5FiURm0j/sHTHa8aE5M1d9yFcEZcJ9C1hQlH2ZySGA
OxjF/O9yZ4A/ir9wod3u6WvewcHmAQkNDDHy8lghzfcgA7ZQ0re3jeWLiPSNaxetD7cMh/vm8Zxv
y8BtLXU+1jIND/f+Y99dDjTbtvgAkOF4ib17kdrS/zx4QNVczgf/HtXyk4Kk2ZiAo09wvWvy3TyO
SYpSGqxd0SFi/wR2a8ZyMUWTwFbKHNbq2TYEEiEfNFaFNnd40UBjp8UK0vCJ7uHKZ+3/6zEgcZ24
erbfMm12EuAmjmx4LzPr5A1IYd7MaQfjNZoapPxPrAdb2aPiWCoWvEwe1figp28gUrf4cC8Gxax5
CWjK/YTDIWTZBGHUut0/f23w548DZqEsYxRSG7JW4agfAiYXj4f6z5Qb1QajxWh9LILe0761UK53
pq44ZQyfylXRU8VjgFTk3s9cLuhEj5KR+of+XTgn+KJzwJxuFJJwTLkI2dpGooSSJwv9UfG0rEbt
HQHNuAagMdBWz8UOuODE1Rn8xzRXn1cQyVTXqTwmk/9/O46wr8IE6MG+roDfz62bodiIjyuJ4rhb
bsX/WiIF1uhUgE24ZVW8dIyjOeGyrIeS2Zod3wJJ//6IPzo1WHK2M6vtHezlAQ+KPQ+aiut+h0x1
v2+pw19EmKlkzZKZvlJsGfe92gpToMN2hxmQrT474S+akb3DX6x1XcTXR9nvM/v0NbaCUCCUKZ+F
tzDY4YnYiWy1N39bFB1MjBNsV+YJAlT4GQh+gRYfD8iWu7wfKq2xX+7KoTTEVW28kbdymO6+tUBS
QiyxzwyU7CKHFub+7CFlY4xVxMxJ1vk4Z0/H0p7pRPQNDObbGFEDMKccs7/dGYfwyzT+lxFChmnP
eJ+HzoQSDKkiEPQ2kVmhI5FE/zUPLefv7mYP/q7ttCFBN9jO+DzxcbNKGODIoHmLb8AjtVS62v1a
0xx0ncqnla6LBjyh351xY3IYl4Uuf93HodFrrtPkPWy5lDlPKTJq88LRDUKwgyFBL8pV5Vy6h5ke
0wxyMOsbV7f0rT0SwXMWeCmj45BeEN5by7/HAaemFoNxv/Kkx+g+sZVdRSGISxsaIIahixZCxsbG
MNUbXbPuxJXeINwrU/adnb91kB65JLuZ7TrlRuLnvPOK3sdS0H+f4gCReGCCH9VwxGM4JuZH37xK
DsUhuCFR5+nlR9U7ScBsaeGTE05EVSTIcFA9nkuyiChaXlSuLHkCdKaIkWwvx3kpTaUAKSzxCkh9
cVHbroEaDYfqd8UWiznWZWYe+++iwZ4C623T0N7FmJyBOMTl7NuhW+cD5vhHsniWRl8/5ap2id2B
h9ew1RChN+ZfvELRWJyvx11A+X/EP2uL0hEXEexjtVVmoHCAosQzOSmgIjIavnUSrLLvFlZVyuib
d0xxeS5coOfhZKy4D2THfMYocWegPO9DpVgSQSlLlxrlQBer5c1wCvY3c3q9dBCF9LIm5iAYAkCO
7NAwavvTjNu8BT1LhzC1eS99V1yKjQW1039qgTIE1HsDmsf12OyjZRM3goPEDrBvYTt2sYk1892X
WBa0Pv4IrBABlYqy7rCgxiV4aNNYx9AgsQ8+ndekxtvFDdh+n+udnpPvTZcxhfrWhZYhtqsQpRdz
9hO/7Dg+WLTr6tPvlxtyuBUMMsLyCSCVBNYp5Tpf1M2mJUEPJtgR39y46q+cE6SSm6irXVJPZzuF
d5auE8QYrCmqpHZzlKUwDLNNNJ2yJvSBQDYjMAJkCjVQGKvMdmlv2Hg6Y+kAWiYX1gRTIBG01mdr
AH3CteRWYi8biRUtfZ74vhYcyBz1NG9XZ1fSY7uEB+mohOUTJg+gNBNMxfvdDgYPMLyV228a5+7Q
YI3mV+rpNqums02jAl9l168vcRL4nKFmF32LFajczMOj6RxHVvY+1PqIvdmO43it6NmByKUKqodT
n+bznsiEMFw8CpQkIhMWf2U/rEBGyM6Xxuh92A2DdLSaNINXf/XTWWxApZLzjp2eEuXU3tpzYwnB
+BmbCx9VNW693rMz1O+gac7DFNIQLTxQGVfaxDgcjD17dILUx1wTojDLzGsvQRAXhL+g7zXDsKTd
OCmRoznbhenw8XNnp9WpzufGHd7zuj8U9G/CWbCVjHraqgdl4g4BHhMfl+GMvJfiaUd9OsPOYIO1
9ZXIEUrQcGBEoQylbsgbr3l/zbAGrwIxui4+6gvufhA5FvmH16PpKBSbRlC5+IHQBWSwbIvYV4tx
0BGp1R+P1gISaN0zDV8I5I95DkhhhVumqaruwqyEkgpZ3/q/GvQoJ8Vto2OaBEDAkn8mek9vw1/W
wACh9wOsCpiZbknp5lF+g3X915fRimK3JZs7y9MaCPi9Kyymb9bErJpX5jqFdr68GsP2Jb72RjwA
WdveGbCT3/J5G4k+PEi99oO6HNPzjBq0h7fBJuPLrIbZ4TKLmgUGHg8fDaYv206N5p+hF+Qq1N8H
DNMhw0WNFI3m6NSEwVjMIy/61/DWVR0HZuLbh6auPyu+8r9yszXrWtfyB3aMhdrsYMU+jId6S4em
uk3kL7VOybPb7pWvuFoWKmBzt9PtN4wO6C6j+rD2n3lSvhYbtHVffY1sa1K9XHQFDbT+IetEwqsG
Sk2hXmOSDTknYpHQgZ2B2JBYsMBKfCpcUOafbffaBzMZwccpYzq/dXfRWljM9zDfGpO2CzcUJh7h
lYfUsNJb4W7njI705maoOUrUKID9U3BIjz2d04OtXehAULyh8iRRqw2cSifBtZO8SosI0w914Mqb
DsVtDFhLkZycTfZv4QUHN5KmWGl64fSr8Zagx+vcUTBIZT76cWISGzmuTBWbr5FnHkU7w+M1+kub
SRza85GOUNCD/5gwsU43nGjSoWUXkpxYvwz2cf5b7uepWawRtLwK2rjMSR2jYXSH2fQMqAmWdIrA
ewcbM7Cznfx9FFqoqBTXLmmoPxojque2NmixOJoA48V2TAy6kxe6/NPXwUmqbNlff7FI03FmzCZH
SkOh8oU+PZr7Sr1k3jryAicm+7WXWyUQlWJpK2w0QpewnjqFjvauH+nRFHjdJYrV42ASS8EikT3j
4dVZsbM75+uCtfHf6Lp91PvhXoyYGuaNGHwySyBDBfU/V8t++V3wmpX29u9MwpfLa6KBXykIAA5c
04sjU/JqdkYz1kulTnrUspCiDlNJy7X2qKqIWFKJQoQtiR8a51vYeemUU7nHdo1buroHC3Wk2fBt
ccKmThsLGgiDZa7jIGOCJ/+m0LJbxO9Hg209nJlMAX1/qu3OAvrSJayQWT8crKCwPitSjnCGhXhe
7jzRyOvjdYWrubh850T7LaSZilPBNyokH06d/APFh/K1nAmgtq3cbfOZcVv/BoT14MqpmzwsZYFK
rltM5zbnyLoB0WCpa1HLFv2W4QpAoZcdglg4OtdeVJTiPRIaTIJXo3i3zRAG1WWAsujh3fSsac5O
rLJ+EwfTYY+t+XMq/iNDVzu3PeCm2qnINRE394jB152s+sY3UBCpk7mDGPxDEosy2QkKLqHqVJUg
jZ89QhYsmPMOC++nASfXCGFAab5p+GLj4l0794SJbGRYM/UQo3Rj8HmDsq0P3Xv1Iw1Xu8DvUJWs
PlajKWQKw8PUVx6ASxUg5PL43N6us5CtgZYoFVSVX48/wyEVgl7TItTMR8RB4oiExYKKhqKP+LhG
Hp8VqvajEmIbS9n/ci72Mmw+3X/dAhqa+q11Rqremvdif2cCnk39nJNMnhOsqwZQTbg8gsI5iJAC
CLWw+aNNFZwcTfEELB9yczSHzgQvXY7AxLXZUqVGMGch/f3NcFwMrdYRVSws2lIO8P4pT08LhyYQ
sHVkTYWEVuQGEa9PAa49yeJKt/rKB3DFUo35+7meMmCbz8DJNfJePLbK+6RciAlqxKLfKIktWakg
4lF+N9Jd1lCHenM6r8CacRZrDJthPfkuoNRp9Jr4hhcye/UjtB45VYLi/F2ZL17dVKsAUzXcrlhB
OQdK3PyCb0F2s+uCAwUI7fRAiZM6GUQTNHH1zmfkkdnnKprWYJXy32sCZosJRyf8JFXTyLjIKjlL
Qr5/EXAgVmAM4HPPDW+liGu2TxyPIvQV+cQj/8W0X762rLMsFZUd0ltXajXT71ZREOwEkvCtdPr6
lST9sBBCGXAOkx0xyh5mGXAyqSiJyrS/ZwfXRmvNZFj4nQhaz5DwdFmkIzKWgxXKde38f6WckXry
ZxVaGxgWnPhQwWFhqGA9kPe91Sfs/+Cfqh+FEFFgJd3J3aE/RJNRyWPPSJQZEdCLuosCXfJn0dHO
Ykb1YLFyK/8HlppcaL8MiZ+Mog4VcFXgCBoUjx3t1oNqMG39tQRZrS81fVwYXOHmML0eNFSyRwU9
Quyjm9i3/b/Ev7GcmmIcF7i7RnBpFtwVxgth2TUzylvNJn4J+0Hp4xbZztBelUo1XRSrczBCSszX
NqMYCiWo24hLpcM1rcfUzFy2KiaNrqWONXnvARLK0WXsaP71Kb85UmLkBfvnDfHOq9kp+ARDgNZo
rMtWlMzZkoTiEcR9zHeQWrj3mZh1JBllsExQYTqW0hm1Qh5FHpkD8ccfc32zABNDK82L9tJooPjb
MYr4YJnLvJxRKBnk3T3UQpN1Tu3UqLvxoMKvnVRAzZUK/Ngsar15Sahbus549LWHxhYckxRBQox9
UneSgn12oixEL4zhl1xOwI4Wd9RFZhblpCrmx5p5X30wwxX0kUTM3BNvUCTMVfxwTBdgRgPXtBru
GLH0rvYAF8tYIgtZU3tgM3WEeF7fVm9ph2Q9PDa/yUD+jNxYMkg4Sr3GMf3kTqRR4SGj52xcCA1w
wEK7Yc4n/Jse7/oWiexf/T0EKoxkMPpgpP2Zkl21cap86l3U3R/6at2s4qQmVk1m8KfTe6ffRVLx
QAGvSBTvYez3rfjE7JxEUMwZIjGAum2NBdwJrVjK/Hb2knWMEgoyISPTho2vM7LciOfXblUhQRqF
rVUNXKZxeBIl7r+c7Kett/mV5ABITWA2XjtypK2cyyoD6ETJ3h5h9wMJGxXXO+be1JSnzldqo9mH
e4x7MGHDndhlQ9G0gboPu8blO19DhIulUtnHh5RgFp9F8j0i1WvCTChnjJjgvXJwfGX8aVgSWedD
9evHS8pGC5yD4pnhHKw61IonVpN12ig/SQalFEb4WDQCBu1WpGOeSStNeeWH0sRjT/sbt2JkvnNE
CWllyEkEn3LGdtNRfNIs5CO+cQWytYVCzyTLhxAPa01axgYeEr+Apq+wBCNhcVwOPE9/k0/KBv2q
aqGUXlgF8z8KZLPKQ0YQt1d/Q2Xp7J/Xp4ByMD3yq8EUlblJWh6APZZeTn4Sdq1P5QfGcKjbmT1i
TecNeP0oQcxflol7tR8t9Xw4xRoj2cGq0jWN+h6vvro5HlNm5nF7GSYzUd7b9h3QTdus4aCuAadI
5vo2mT0rA2YnUgA0nRLM4SYUniua1nGGjntnN4Q5oNejyw/3eNfriT9zAssq3ZpjPxhRk8GFuylp
Fq03VQJfCXiLMNXypzH8h7elwD78uQau7zYVRJYnjJ7vUQP01Hxq3FvAkxVC67VljsLq3Sw9nVHt
HxHXZYq7FiBZXH9dMeDvvkoJDaxcNwHap1L5irOHXb1Ib7KEQwTYRdqeh0f+HDYE8rMxYyogpZI2
dh12JG8a2yB4KV0IciGfmK5hQbXbtkVwrTiKwI1vVk3vR1Ek299LsvVnczhrAyqBSIJcYVRIdzPQ
b7kOzTCEn/IkXtOgAxfDwMTNt07U2NUGPK3YxVrp9J1XCzj3zqShDu7bhsVourpFSpcuvNTOsO7H
h5v6j1mJOjcv4IrAHZQNLznhLY053kw1ez2v6TKvFLfkRXlC5ONSze760dnApumObP3tW9j1avu8
s2zCVpuM8szdLWIva7l4C4dtM/uXNKja9vqUX0ZSipzLp3cNhGU71p2KlNqxckS617lOix69u8IC
8CWIMsuBtMW6N/Y6klkcGVOc3NFp2aArBr4arhfJlwIsFL8s9LWwQ1GbLdEI0O76K7DrVgZMUzhN
C175GsTEo//JidN5vBn0oP+qxAZC4RK5vx6qv+0aevAQOrEwYvBKUBNOp8w34k1XKLf5jz0QvIal
KFq/131y2ByPlfZH2wNlfT5bef7gmyQVUVcDjH9SQWFsko0vDwxi4XlLMYevjktpCJo9mwwKaiNk
bYzif9JQP98td5BIY+JZFhHPCU30LB5BnaI9u4sfEVgH364REfi27pHoDBqUbNVaUMtnSo+gdQr1
zytHzgscfQJIgqUzbHqmnSmN9ocWi96qzrXA8Btrkx+GEPZ9uvqQ/nSZbq1fGyCXs4j+a+a2d1yW
cDId8nFFGSBp6yM8sayDV+Oyl+E2KVc7+VqwljIv+3WUvQJdMKpVO22BV3MdPQyEthj3hxH77Ibv
w8MkIUgwtVfSnM2mu8nXocw4t8KLgD5D7vVnTvaXqS5GsDsSanv+F5K5hfr5FK4cf32d22gz1NBG
2eD66i6I2Jz9VFU9yMEIy7yhxlNeCkYL/nLGuutAr/tDEuxrjOWYQABN6eCd0yYnofszaL/8fgKc
J2SlyMgaq0Zz0LwI74JQYmY835O2SjvBUgrRiI9TcnAt+sglLC2cNs6af2GEqjfKvriKLwXFcW7b
U8ceYRXwCn6yz1w5LcQtmSYigH9znCUTzwnMKESBdKL9YtJaPFXICKRgPr8iCDv6TZX/fpE+3JXa
fnyN/dcG37dp6c0i1RCP6a6kabtVgGxAsAqrDGjMoZ+CjbnJpo3x6kmP1Dd54T7lTRq80FJGrUnz
b/4oYHINg866A9xTIsglk92d2zC6WX9UzUZDcUzL50fpAqaVe+7FCx7uSTPpKIR+J5A4oYfLLJ0s
haIEdbfNe+1meVQdMxq1/th0PK8i09R1RrRrqCqArr8zsBHF1M/jcAstAF8d7SwcuyhwOwkl7XbQ
17rbnkQLHsxNcAPleVdaCkCbwjymhhR0ORQCOpdVW61UsRUzvhQ3q3mpl5UzUqcSCJ9w9RxV7ov4
zp2SsAk7fGhfYnM8xTtXJgxvsmFgJgqYHrN9AdH9aT47RvYf7183+rM5/HbPR+gauw+WYTDLT1Bu
0BpM3RWfG41yaYhpi4EaiANwFvrOee3GUMR4TWvhxfucWI5GNsNI91OR3a+tRYBM2QEl4XKIO/Lo
dfILQQB742zTvaTvV/nMYuUmjrdnc7wfc3SMRQ6hf1A7BuLS+650MAE/recDdBtOzGYnAXKsvfRV
hWMWHif2+tJ9hoMdpMJds36F9noIGAanljjvhuP0VXadrkgcqqu4Equn3lnotWTYWL1ThvNla3v3
D2zPXLwvMSRzdQZqHt+kKIcwEFzWktp0KDNm9r8j2S4PWxOdWdlGJfVhGKQiC5oBkzzZOvh0N7hC
EPHaBXSenDKPYHCTMv/YhkR6dFmpxSUP0/sdpRjJ90PzVSC8CuvigSibf6sJLAE6VskuzMjBOEpH
xSYUfEWWtS3JHmOkwCQKqk6hup0aRxFIhLxwDNASbiHTdHoigK+BEThLrlc1IvLvPlWwjjxIZYfZ
Q7FL0Hoq9/EMXuKZyYkqciK7ksWvvTUb5awD33GD9PDteg3W3j4d0Y9zgR4n6s3b3osKyY7PQS4O
BF4xf+Y5ktDksuu9PbbA4ffgPqqRu26XZYPqlXgNy2Y+77hOC7oNRnN1UKGtnJpGr9j9eUmFBw1T
QobMw6awlB+P/SQiYnGt0QgSMSBs9v4fGBu6sGXki0GIUCmIRkqpOcRJvNoalB7SSpGmL3AF6iOM
Ab3vf4+pbzjgvimHP5ySyOOt0BkgfzP64vCNYVCFmFYNiTdL6d7FmoBx+z6jIPjQr5IpKtxK4+hO
GZiv9vO7+pncLf2zdPcSXPjBLtP/pkWIUvPGp/RVkqvCVzxGgVEgoYAVhwhVmIXF/s/ilsYYOK0l
6kV0jZwWSKNA23odMdVKbR7KRU2GCj3SiS0890p1u0GxLK2nXgK1EAlE0VFwZ45TeE/6p4M2s3Tu
s+DiNJ6A+R2AULy97i9n/sSvg/W0tfOEnZn4s+YtEn9R2uJUUzGdTubmb+DAb4HqNegjE1nxErLr
eVEmmKY2CLC0b/BUmMtDaCX/kECPQu8LMmP8xzhUFET6M+SXgVQzUkFcKm8uXEAC9ql1aDp0zIir
CViajrqGib4UYyl4rbrvEXfzN/o6ivEPc9bimvHHRec5gk6R/Ks5V6kF8aZPNa6hzVOVhbIIivRd
HeyT3SPxVVzmM9e2XMNTaqQAhcKu26H4pOJHQm/hYX+rpGMgEftu0LeRDpAv60liIjjjEm1L6Dx9
9rulIu3hgyjYnTbsqz+CZKMeoZoxyvx6mwAjh0WJvro9FfyGZuq5ru0ewTFlqQp4tRnaCnzFX0ox
5HQV95pK9rPY9MpGY/EW7B3OcQ5SSk55aq0NdZ9rbxNZ6MYdy7jd0bdSf77aDN/UOsvvA7rdU1Rw
WIpeJYsvxfTmMJtWzeDeZWU+SmjsZu7RUppZq8vX/anOAThJjTEHMcRresHSS1dJhSVyDh9Xxctr
0eSzXoEI3ThZqI2KB+Gm4GoIW7+vWNM68trUdKsA9FjXXjZVnlzLnGQDLquuZ8FI4/dk/cRsW0e5
rFJf/OSXzBBsqtIWyItnVaCijKztaYp9AoitehlXzt5px7Nukk4dEwd6WmOgHHFwLBrZWZIiDfJK
xTHJzZ+jzMDhUNM2b1B9gC4sg4f7iPp8910/2HekwsDP0nIiACTa4EK2yNu9f0gkXaxqTNorbAii
6IObz2FdNlGouegLPfXsc014YTPVIXNwmFgC9P3mkSxoXdal97x6zfOHLi2VLpSnWibqCa/o9f6h
mwkWg/s/6oLIiS2DGfy71TQNsrRcZ4A6QxUCUfNVxpNK5pP9MNjg+hAjWzOjpbWz9O3sQLrv1zJY
hpB66v1TcEuLMAF8Si4ESU8pb/AfmyV+VlOGDhzKrY8vZPDu0vIkS2tjLzQhWIGBOhHATH5zjZt9
cHTfIE76iQpceys01pbHqEphg0iZJP3YRE4t9zuUIaD32ZBZoGkaPBqMRMK4e8pO1GnEJWsCGgTg
Ka9XckM2FrjInDtvlLgak/9ZL4V95ZAnwTZ/jrq99Yj8E1yoaGQJUxoZBUW17N8GyjH2TBPkv1da
hbadvdW1dMND8Wsv2CEZfPrmC/ScR5JTPPZUOQMkhB71+ng1jzS657KDMoedhw4ISJjCnZhDnu1n
OOhmuf4PY/br0QAXTHX6GGaPXmm5ofWbzhTgbrz+avvdzCAjH8+0QHQSj4sAs+e35gg2cVCUw5BK
bobFENydX1d8ykuyL7/okyemAp8CeiDx60coymdGGu98fc0hLI4x3IrncL7PadmgXRrUVuESqbsY
aLNV1fm+JQ9vWZHLi0qwwBAfWyBPLR/XCQm0cYLtFZO/VLY+4/Q6IqaXIny/tw36rx7/Xtda16rF
WqppRPjBdXBRWymMG4axtYQd8ZNbJK2e3MBf9F+xqueILuj4m2vAxcwLaS+XGtapVYFEY34ZGFaX
Ko4ZvBUkjvX1LF5qGLE+FNYt2h2oLVFU9eTfuUJqbV5SeU7ZXYRQaeyh5YUgd6rwNGP2WJ9TntrO
4wlv4jwE5QQQRabXdkPHGISzQxcfEkFfdgnVDGK4h89Cnyu5hRxwWIrdr/GYsEF95qRCtJk6Ey6q
Du1zsqJyalv1Ep5rLkNkh6jvOZfxRv2xtqN+5k5qTBHDh3BjROfImAJzCZm+MAkN00I11fhzOg6r
973styXKZ/4PJ8TAes9SOExvPn5j0uMsWCxCNUaLFF9HrpN7UsdxGG3uoBYJnCA0Rn5ML3rMQ9Jl
4i7OFbJ2A0eXK8uGQm1ewh0b/NagVQk+mAWIgRQpu0dF1Fmx6pFjVuPQxh8O5MLG8lUfiCIv8p8p
raC3m34DKuLys/mm3+VgbTYM+6NptfgkQNjHmCUnM/DdLGhWGFOEX5uz8PFhVZXOj6EupASkE6kP
Qd6HFZa8akux1yZzYJYsaDPIQIiJkjLA6aw1UPEniUWYqDQyUgBdAv+tFPyc2uu9k4qoCn2dUi/u
WjzN+6ES4RIm/0WhcpaMV8k+KVsiofnI3JKnlm4M2Bvm3OUHqwHsWcWily3+3qJj8ZYYKIhffpXG
cpnVUAs2Z6CMaXuaPFDVqO810yRSpERUxiVwGhtCZhktjHTBWMIMOhdumeim9WETrdkq3gpxO4cC
NWzWawNziWjGteU4MF8/5ZLmP1iRD0LalT1lUAxWhXjPfxTGUXeKH2fAmt9ZaPC7NobdXTAe79a3
wXmAWRqCZBEwU1JEO5wmhFgmK+UtaSB3Zvsfz+QZKPfbIUFao0Ch1xDI/7kzk7tlqYEizIzSX29l
ExV586WPJdsrt8skVbw5zDG0bqAsDD3Ua7SSi5U6bZqi7SxAUkB1J9hyqBfBsyPpxbwI/VLmpwgW
7IeGDofj3z+Zd+62Ls7wHasUl6WsfPQxGeHat68ZICgEnDTp1tKM94xHUcQvp2iKR0+yoG9D/003
xQsv3E+vjt0ph3cB4ISSRFO7iCaRJqqeU0kGRzaVDdQ5vccSaoQfj+C46DRNdw7DvPAFinZMu9en
o82flQSBnNgpPLtFG4EayiqGF4XPFP1fTsQNLGWyLwb/CwSSsPDv6GsDObmTsx1C4ItrBzhdWDXU
SJMeIuh326Tm/O2ISFJpIoAmBkl1OdyqJEdvOtZlqSo5mqQHduBFXuWO5SPLYXtw9CHJs9k1wtKn
aJtNMssDnHIYT+WxMhhKj2cCEbHmkYWZ+QZSMnSHSickTdeQs3K/zT/eOLjprtSvCTt6tFy/yLpY
fERjEgnRd8/32ZqArg/RHvr5ufeJyx8p4mVeII21q9p5a4pLrjbVQarP/cIYbbxvR1PPSazoSf1A
XVCEDiBe2S/3m2EM1jxtuj/fZuQqDGp/NpMajGcNWEqNpQ+lEWuH66Lq9t9mqUiB1AQM8TQa9YMF
Htmuv4X6zYXm02tv7cK+Ywud4SVbdbwRMgCZwGZQJxY50xIPe6U0W5mNxfaomSVxYXq/SQyau1D6
ldJ0QU1/KdCbL83852L/DMk+G+gPra044vi6+gM/Ixm39iolnsm8ME75D2qz2/UZt3racGyocgVs
I1vSZ8B65BYVkaD9/WYErjkLCMwRyb0GwdXgFDlW7gwNHevFlKi865zUDUfJxv2JxU9+freYyrss
MVUGoE/3haOHq2iuAp9WLJyL+DQhaegcUcGsCk3N4/02HxisiersXzhVw2tRrD7ah54yLPLZgD2W
twou8cFb0IryEUqOOcBvwYIkDdhy6enoI3JaxECoOHo2Bpgi+Vk45ZHqb4m3gNoI2ZmIknRZdpS2
c7pIR9vsUz8cZJPuEDGnAr/YcIYJkBXobq+panUl5jDq1uPS9XK1zDmP5XEE4a2ElPOULqq4LDS+
zcVM+/droR0nPDT4HhPuwTsnY7/ftcokvnM0ABQ1VtS1/e66r7foriar2FxeDdE7+t5sBwhF3I0+
RdNqlBMQ7ewFDCm23gnGmXJY3KzAxZ5IOf3is/L/zCKnivatTSANDU3zoWdYLIQHbCFjI86Q2Hbl
/vo/gvXKt/HzHiMxKG8tLKWesTBVn0OQESCHCjuq8P0wtFoFqJBT/P1E1LXOm0o+Rqdg/IhDpgxs
NcR3DWqB7UpZlHGGA+M8RaGjGPZBoV3/es0tEesDmhev22QAPwynZhPdrtcPpy1OnpJXJsPupytV
oZoWt8Dm2jnDFQKtYDbOyBcMhwrN6CeDTcuqNKj8FOtPZ7KQ8OCyl8N5aW74MjZEgvrbDoMVX5oC
SPklz3fYyEfBA7+BvqBmkOlsf4kkPc/JSdKS6pn54LNCfA+xHe+hhfbCgixoJnWbihO9ilVHL1G0
38JKqiTZnukAlW7N9j1aXAkY1ZyCmkx/3jzJd4yceAtvpB7GOQk/t691xt6l9QGDYVfGMonnbhBl
ef4+FLCt1qw5BXWrWEKgK8JMKtek2ThKx3I+Z8TEQNzELZAxydlwUihQ4xuZpWdBTh7YKdUQ59qX
x0DFueMRddj1jflqCYOhyjGjvcw0p9klaXf3gOnTLDptyutbVCceDy5ZW0Zrmqgnbf4y7ywpuglV
6MxqTIaK9OUWMh8oaoShQ173CKqfSnlsqMi13gCZgcUpW/m5Ci+m0fuJC4+zwBU4wrm5oXx6Y+ii
P5xjnmEO8TeFPz0j/nnC9FjjbSb3aEJBB8Fkq41sv1bM9nwjPno62UcHp8Ux65kYSewJvozvqO6q
e1eflRu6DXbKhOsOMagkjELYoU4BwzF8OhFIEjutWD9BtmtjrVX1jhcxTg6UkY0/64e23iXd/af9
Ghb15jGENppSyV0rYaC/hyRSksyjvoReDc0f2MZQrQtRx73gQDUAOCu19ryjQ3jkuOiUleQF2/QD
KARqc8OOuQhN0O5p3vVmv+UryOmAEXdGP280rwLiLxCZLvQ7WXYHuaTu1dp+ZdrwCmaexC8BtxCD
LvkROmFLJTKqknkUdTBWHDPiVALkcLBiwQKx0ez6uOwo2wxEJJdazolfnRQ5rNg1HYE5xrkp3PvH
0zDqH3QJyJqk1zX27i1xWEwZIC/n5JN/l16zwf139tNzLRn3TpsCYrn3/zhhHY3BN62el+XbdtVB
nuTk6qn31vUVIQhoALVzhIJO42Ydvn8vZWJDMNwrAy+3ZaIBI04CL8u9q1vklqYR8d00YGgWLqSI
Uu95lV2zqRTwlLSBtdjzekinHGHXIkJTS6OymjHgj/RTPKj7cnmfi6D0uviyMdwBNLzApheKM4NY
1tZmTYaIwD0JKPfRZ1zli2zKtWLghZneZcqJ8TvMpBrQVH0rxQLRjqwyqvk5+A0VB0PRVVkqGysB
OMzHe3lvEWaoNvK1TE35rhVuQOjAg7IaViHN+L4L8imnci31jIiVCDRZFOZyYGbegF9WT1a8F5ci
jX7/t1zEhx/Gmow/ecnAKDnJqtzFzn7NUtvFYxX+9BKf0y7+cA3ydXCV1ZejeCUj4K9Cjs1YJTM9
MlXCA/JQgRU5SX2Hi+R44F2oeSGLJTOmHdXbvxQeWZYX/smUohlWktu6vONar4vNrQJhL4AF01hg
twQiJ37w+rTAhc+Sbe+YHCEswHMBtQbxOJr17vBnQr/kXp74o4vzhHP8pVymjgkVyQeQMFrmaSQr
PzxcIrnlF1NeCeb0H4EaJGNhNhzRtlCKHpO+0M2t6tBRQpVwU+H69QNlysKPn4aQRAhjb24yhW03
yhFC1QSCQmon2z0chaszvNeVKBmGZedAtMQXqyMjw2nRSNbC5/LX43JyvhhL96m7tIhWNbqXmXBX
yiArPt72hEpNCixVxPkaJKJgGPz8097y9cUhS+pcPYvy5b1OGbYFnjAcqqsI7A0mhILLclZ4CM1Q
uSltq/hJvisDuHziJFekjzSB+O0hgP2oQrr6YOavuisn67KcSFc9PEybkPrfq+6NwPS3G0T7H3q2
tv8EWbj0hy8r0y4gHMr2lgOx4JsC7WUpb+3Q6AnGmVlP7F7sooGwiFYId2vNSOLJSm2wxXrH2Vx2
QIc1kXXKkNfviX/HKJ5RpyoAZcL/xQJOCf9oQQ0a4uXDe7mnxv+uh6szLjiIrHppabL9K05YwD8L
HP+ddMP/mCA8ESPf5pJRkk5sqNh23Gaz1zcILK7HNykrfnDQI19maZeKMECIMDxUT9Bfe68woh+k
gWHMTM3YqhaBWfhmjPxVy1DNTbgpxZoMFjxK4ph48nhdyZ96W5aP3pC5OE70EXr/EPq7rBwt4u90
l+lxNylTt8PxuJigdf7Q1UVSN7jJa7tapZgGDKZm2p1pWk2O9zXAmurWGqzjDQQDF+wRUL4nCep5
i1qZGNWMud8IOGK5SOkRXlNY9vQrmVigW48GvYWQyu5j/lkXcVikfGltoxWPbbG09uK4z8j4D9Xx
CimjMVvy2EyqpUlZsFGmGIucqCnyI0dkxlWPFfPzGFROw6xm+UsxKeqtuk0D1DFxwKXR/6qg7JWj
vNnAwWWyFwBEy8GMKM0WfVRabcoIyImiH/sasHIW+glZQ3yf0Bru26FQrgiU6aLZ6rkaozBTldrd
Df2HEurEaFQJ77NtfSWnunc/AFmIuX2OeukOSbMfgNyGQVyOfyLn/toGqdKZCQ/sQIkLTFs6WhPf
A12m7qmlQ0AFaXvgp49lRjJRBQhrTOxj9Le6AbVcTjjEVTRQjqqMeGjEg7NCB5ktI6WgFTwlPLeA
Czw+CMmwceJwo4i4QnBv0e5xyoJwfG8hO1Vm2nAkiyEKVK1KDGPNxLI+nn0Mb6wscs/ZzM3E+yM0
z0WSF1zbrhUBhqqyw1X+ykhB3UZsYI7WkaoC77Q2Bjlxeu0yJSAEFL4dz3W/RhvXetohNmb5Lm+b
DMBVZS3rET61v4/6tbNGIpshjYGGNMcNS8CHdwJvctt7xNPM/A+gJ2OWzcM+8HuLb5wMPsuilS+i
jWtMO9UkGb+gttt0EnQ4HVBqYAK4IH/KxZVfogVHgmLgzWm2/5Lx9EjWrYrgV3eYov6c/kqIkvR5
fBvy8dQvt7hfXsF9WExJG1HGZ6YCoCQ2876Xi+emXYckt78a/K5czg07iBdlp0xTubAnnEafIg8o
vFIXLTse/lHcJEvbcC03mIbGfcsb7cR2TFtkBQYK5e6kjcxXyQT+JGWfVasRGPH14BKVoIt+VxcQ
ZUVjrbxP1QaOidoG5JkoJ1FsukkQky6bEBN52BQ0y+Jp49s/XpuWY1wcVkdm3WFuqEEJw1UeAB7A
k8S4m6M/+zw6EVwTpaJYylAUg8WxL06/qHTewInlcEbKBkjPgPm2mYC5SoqWwdcFfx53z690Mn4C
qP/FkPk7zBqAVt0Vw9c2VNBkHRWpdaFBTA/+Wy0RywKyBN/Ns9f29urq5MWvjoIWEr+Tvv21FHmW
nCjCPUVQGzxzyQU2dahjHfUssnG1/O3/50megm8I1ocnSZ2y3mhSYwYFx5Ldg+ZLW+0IR5aLwWFJ
+aZdCdYfydJLKTOhEhL7CtTavOwrRJZmDLkqGSoz0b1/Pz2fCI1YRbEg9tS8Z8rMkQzmjL1wcyV7
ovrqCF+psNGBhfq8zGBgp7uRzZfgo2xg4icaxcsTGGgHbxftOvgTWcuF39rAB/poptqLkOwWwxDL
OpPSJJOIgSQ9R/V3Uv8HhU+rBKPC4Qek5NbvkSN+uyEs/NpLABxVUCKkvax0hUa401YDlPTK6Pqb
JynxlXwFz5FA1b8eHsYQeCRtOLwkmH74zShaKTJvFfq7IvgWshjMCnNEVPxOezqw2/RKVCi90cYe
VwsyQLm1rGa7Z28SZeXpURQqDZ3WBs9yp9ncNzwQ6JBnSBLR0Z+tUIK85Ze+KWccqQSC/UtVimZQ
PdAoJDte+DelbiEOPa731oPGB7sZ9RH4X3Q1pcyc7XxRMCkLQ64Mb43U4AjhvPb0IzddHgoEDP/K
OIZI4vr37MO7uIpNDImKRHUqRMZFUPgJn8LMRVPOD6/vRGOx/ddqeno5zAJJIFVi6V2JZOsnCxcX
eXknx4Zwty4BbcqhrlZo4xxTDIeXlPzXBmo80wgLcfC0xAn2A+KcpHmfJSL/ApeoZxCP9WrwZEBG
lhaYtZmYzsA8SKqK+cS5QZoT/QgBM8+Mjedv40kof2ghHBPP+s/ueWJBWIz02G3zAS6n3aDLkCV9
mY/NOo/jVHg2Xr9qucWu7uqb2AdwPWuKLyAYtYqITYqnXYuqWSR++mtda3gN4V6JBvtW65uLyyW3
JZCS7CL2Jx1nQoRPZ7RtMbmAE1QMEulru8MB5Ag4n32KWq2bkl+4xyymk5VlbhXRuEBUx6a9+pJZ
xCs9lG2P1rNVXxA30ZJsAfQkRSRyZna720k+IG0oDxxfnQiehrag1T2wP0+j+4VyhnnnbWkAPu0E
soVjJubAeeusUTqfIaoXZXoUYsHOSb4uBelUWsEqgtvPwDkLa90qmI6A+rKs5ZKTNuLWR0FTZEMn
fcP94fZrpViaXjtCfcNITNAr7ZaqUWgHoWN4BnPmvnwCkyT89AwiqbXhsLVhBKATPYk8qDMRDLW+
nxKllbT3hVh1sILedEyn3+y6bql4wiai1TZW9IgddtXIhP3XhBaoxK+PQhLGS95gc50RZjpgIGi1
P/8PmM2rKWggJ2BZSarsVvWpHeIAdlv6wGX6OpsLFOVSOfiqJpYmxZZJ98W7XXmiA0udaLvI3qUB
Jafk4BdQpTrEmaHhZjX7i6FNjX9jxQbFH8ObSRfDc90FojF2Q7GVS8qxChFfvXCZWcDtK4ERU5XB
92wP5ZTIJJVG3izOR8DlFYe5G6BoaT6B9PWAEBFCC0VZDAgNW3RfGw2i4EN+s/sr0E5ADL/Vo1G4
M6wypR/XkL0WIwUPImGCUUbdG9xn74iR8Bfc+vNl5gokiyCB1WRn23fTunL0iTxTcbd7WM+Q8eAy
wHTPP+7vXi6STP3wi7/iMIlnZJCHY21mg1FTsXSdaw6uDdaHZ32SY5IxnEed1nr/7OOj4U/FNm7H
uXdUppu5TlLSCb6cvH/kdc7D/mqu7FQ1G1GaagKIExgjoq+Jn//1P2yZujeh+6emAa3Wqnj26lU5
JP9/Ao9T3jNQQ7WIY5ciaPo2RBDAXLIbIxHEYYeHOOFV/8e34gavEGrQtAO3xmiom9OjY1/65x/H
fWDPhmjGhoRj6ttXirl4fSProm/wn0ca2uF5aLMqLMMqGb1uOjRIwLtVGzpq90pc3LdSrGU5xVcZ
BX6pGgIkbmWCTNcE0lp4hIL6uVxtNwbCw1sIL4XY5iA9iqAzpXkmM1XYmWlzTcAEt/7cUv7h0932
YaGSojL9n+z7XSrBhbYJexmQ4P/ULEjEIWn6zabLwpTV0OGcc2Efju5bcamA6IpzgFhupbqCFdCS
hG86ME7lZPjXoMH7zJrf+oLA41vY7xBZFaGi7Urh74YJ7SD3Hq7q3gV2rYpTF/Akq5X1uKhfoeBZ
jb90aWP+earWlIsINtksBHGeJsCQOIf5NGHjyN0VsTv3N9RitAuKEqcEgcBahOnp8sNSrCIPRPQE
YmcaQiaj3h2nKGg31NXiDz1sIkD+8jrU2d2QN1z2Z4kIviGjIhYBnqnwyciLZP5OVmRbZLWiFoML
OI7bqC3JXCNeAcl0O+b+NmvWoh31jwf6YIXqp6LVyj/ikEdBuKtQGQwe9AJWqx02CGaaxLlww6MN
Tk+qsKhRth1Eu0+sprS5kWfgQ6EiDaPdLH7R+Lubj3vCiSFV+hHMXCyMH5XGah9DgeA0mKoSFB4x
J+bg0muAcQLEUm2iJb1aBgH2Zqpyompm3WiMHdqLOGYJt7GoTbz95X14+GgG3fhtRHuKteOM1Qbr
Ht/UVlEwn1K9qeP8/ByniFyRP15zLF0t+AsfMI23BSUiuyUv2tQd1wuec8JJp8vMhqfihzGqEJcz
GVSji02PoON2bZAOHrQwRwjK0nFYRb3CLEzOnO3PJVqmQP4L2zM0I5mv5QVwtquiQa5EFKbp5yJu
A/XjndzFbUhGAUKLbs5/8DYefqqdtypIanNoiCVhL32UsF0iYPr/BrvF2FpKekQK4aOs7wWmDlnW
mIJ1WYBM5rkYEo7Mr4iimE4x+/10CNf9JOPIqNpYxYxDEWRjjU5sNeRkm+H9qanrKIO6LWt2GMtE
txmM49wtIX5Y4M52epoG32byFJwHHq10GYDj7vTpXaFN508YWZ1gEheev+BTay1KvuF50C7maqXC
kO82oi13TvS2Txpa7rjWkCX85asspH3DaLWoHceoJkvNnOcaTC27bXhHtyulRbscWjn9GWNedS+5
1+b2B+CTDC+VA/capTRr9OgzhC6csRh9VRyBAzHSJEjKBkGvdOdmvXc9QG8s7kYGucZoqC7d6SRw
BtMKG0FGhulGbk0/raZ1+PIA738z3dUFsPw3ZUKSS57z3LAxiYAQK93mvuNEtD2/GSaiHgSUvInO
8YaD4ITm6yZa5zk9KLpwIBZBQluCclOzMVUfz6sIM0HjJDYFX3V5FJbwJumuV+tc0kRAVwVertBs
ELt6BL1tDVbNGqVZ9WVwLYV4SvT6WpoFyHB1kkeAiFrfWGQG+Gd2akc8QEd5JspXNVvUDUuA5/Nf
4UO5sbU/4lOx6POhoB9hNJIu5OWZIpye+DqttK9s7PK4lkZULWY+zisPkPmpsEWyWT1FyM3fnF3A
/TD9M8sdQFQvk3Nr4m+jTXybVYQzDCyOHGoE/vYtB7gsH7vbHEKQpTiIprj/JwrCANUM+hnfNe0F
q2yR9f9D+wBOyWotD9hTL44X9NgppzbIoYl09fqF4CCEQYVPDU3Ul4PL/cC+qwTgDOGSwk1GknC7
PRiDXM4ZFWYvP99q+56CwFKsvMMaApAqOpL0ZYd9nP8GjnvGkw0QWA+l4+foaLGLkExTDJNfXzUy
kdVLM+0iahIxjaWwnCyhQommC1+7W9DNl0k+EneCf5HZ3Dj+UsMrSMEMunzLcbrEfGzHd6olBzVn
qI5CLFUA5MdJWb0plymJ586lZo8A5q4X5coBuEzPBwGCl8IXcVyuY5BkCi7Ur3BmPZ4jFmO8qG+k
KxUkZ3e3essWKLevLn/ByUBs3McEjnqlI+juiIvdVJ4ejy//CMc5UC8tDL4fsuC9W5ve+t3MY1UM
uo1vNzVK06LzH2axucsbQhhuwRDj4ZXJKXO7lKY+oCWZdlBmyi7WrJo2FwvfF0vOO3MHcJjKEkSR
TBP1sutxGvVPh0P3d1diooIr526iOH06o6t5Ip6GWTkHr+KiTUtmYMNWBs/PmdQul3pDGNAPfCNy
Jhe+4sQdDE5Gl2EqUG9PK5Z3IuYJSp+EZ4t5eOZYUL140Kgbjj31Dj04PNE4AhUcuwBqXKUBRr6h
UegI1L08g/3gH5141eRvs6Vvu/pi+x0cM3gV1W8oHApmgWYpJNv6WyfjVoBeoVqA9zrH8ow89N1V
JCrRCf9Mm4oq/R2JBfRGkTTZo4w4z4Yt8xJgUxiP4ZpfoEPnhLrkHx0A22ApXeXN7cHPW0uDj3T7
BMuQ8q1g2Ewbk6ICdkhWKEAU5ivh+ZiruDOeiFfyBfrzldbHcI7yInt/30yQRhbx5uTKc62F5iaq
fhwkRskDpGSFIjngSXCZju+tdkcY3zXjMW9vObSVqo4/3mdTISR2U0zQBJ85+Y4+X+hPhK76TAIe
sovz9p1isDEo5zgWHBCvSYDNWZZ1KLJI/ep5mQMVooV0U81dkLgj8YEbrhv99PaKCKJrRtWBWg92
va2ZHjETHxuzYPelabeK3T5tLUyPFlNRNWL8htAtMAK5HzpkaExcjqk3WqkoHPXAknZSUXx8mFC9
wATpjDXm2cN899onPTd2A7U3vAfO0e0hPitlzVaHx1+pir5A4Q3MlpvGhNBQVmmzanpLbQXJKBVw
h2igjjhD/DAHkcrhnIM4LhRw01HCBojulJtti1xJoQSwfoxbOC1Q/q7T2k4eawpeNxPn/mmlyHmr
y2BuR2H0NFxgVdRB3mDzvco7bDGLQ41f/8R2y7Av85DEV6osVEwbeaRiOlLWAb4wdEbLtkR0Dl0T
9qQtG7uGPZmy/gphiEs64GtMuZIx61RUTObKGa/pWt/vtNEASs9OSLJ1/15O9kW6Wl3oREwNKlhi
9nzLHbOOSivEf022zO2sU7VPg7LC4AESGeG+sYRVXHxaorjiSFPtsFHgYgTBbZvyMhdorYVa1PIB
y+rTFaUqCKgtvp8axzEuqJZ0gOnNJCp2VFcVd0hZttm8UrV1zS0bI7yyIIhHcM8/rfP1S9+dvFNE
/aDf6OoIWH3UuVlDHNLQuw2Rog3Bqq+1lNsXZmwfZfxo0mKSi76JzmjiO/2bqarLYgiOj1zww3m3
+nx3AIXzGIkCMRi5zhDcwy+sLROwIZ7f+VSa9zfoo7+P93NKT+VTK+BFYCcS+QJbikWS6NI66u55
SiDnsujiuh12HR9xxVn8OKeTmDytARvWxcVg3hy3SRifYcCPpGas8ux/Fav1oiZDFsb2Kpoa5GoD
aAI54BjotseS8hJ5Pslln/SiwYop/B6YOmCkQcSv/rQ8VNNrd06pkLs+98wDtGpUwiR9WrNdRSmm
bn2KV1RJNlG8/Q+zOapTliHCkv7goRkzi9X45Fsm64YJvPrfgBTm5QPluklGqKb3ZfvdvLL3vShF
1zSHmJMD67Glm/r4cnXVkqijkApP+Q==
`protect end_protected
