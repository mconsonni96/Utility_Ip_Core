`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
L5aH1sX9ufIzVNUNNTcMaVhDGOg1MDvBhGuGLWqhCLD8UyMi9zDIDZF1znWmDKYwtqggXofBHtRc
mDtJfkXboNVL7ME6R4zw+WDYrN4IZmk/70ouTOLHj4nrohe02xkfOS3rsgUPdGgDlgQpvxVKtUV5
YO1+TO9Yvnl6IaBuO5TY6obhq72CGq7pXBkFIj3+XItnD9I7xKhz7rA3kudJ5WIhP6mxq7INGhMJ
+z9DMnA3M5rimc1ss0Ukfk6yCsn8RQrZCN2xEydjB1+1ExbHCPY7ZfpvBMBKtSx/FzjBbi9hRSzE
LKsMWr8mqsqtT/u2yHGLyEZgDRKGYI+Gg+9yTQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="P/uD2qGaKHGxbtZXcL3xR24F0LDkRJDGX55ZTqXvRpo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8752)
`protect data_block
1x7wTU2ghrFQs8QOkLoWrOcPtP+Vssmw/bloCUrRcgO/J69/8dhDLn3U67piDxrouHwFL9PkdGe0
yTIdd6riEv2g3ylUZqAVm3hR0ixOtqL4YPSGAwMCddFr+8ldBMY2SAnPKUi7yR/P098qMO1kDZ1Z
lnU+8BGAyCpXR0FPorGtC5VxuEQNvNLIB40iPtF6qg4RFQMGXwv9v6nwzCJgo3sBeSZ8dLEiLsGn
r9NCHakKNwZbH2ifS6/iD3haNDBLBKYjSN41jLjb4spqC6Axe52paoda+0hJiZOSLOpJXWAgtFvb
7dawBJ+o5Uwmd+KwkPo6slBhAABTLCjLaIabWxq+8M32rGWTUZB9dq4Pu3Z1IrH1l9tVjmYkFryp
G9mvpK1sEnISccW863eujF5xpIXrZ+mDksP0FKB8QYHAGMhnNgLTyg8VqMdjUlGauB8QJjJRWzd0
yI+RjM4R1aIXkLkjpOEDIhbEx7WnZreB8ZXgrBAQXXbHBlMdpBKZvUjfaotv8nxO66t8EzlAIgqb
mO/5nPj27nOz5oRqemgfJLKWYv9BTSUG7VXQALmVavgTT9wDw1ZYfrlyyxD5y7EkW+bV6PJXRPrX
eozijTk4oXOVkx1dEHQ0+jstPLRjEwb6iglbCpO4LG6JERfapbkfC0+/gEIumfvztb2lZ2Ns8C4D
BpA2jk7CL/9KrFnRL4ddO0tshaSJ0wyyovKPorEuTmN5D9ijgBUMuFIgDhS9SHoE8YMmfqF/tfsV
fIQjeTBHzMijS3B4ocOMtp7S25oJnkhzq+gr7e1qgNXUKMBUJdd67Wq64oAalEw0m+1g7HgU/Rhs
BUAqSplbIHEuaZMges3m8PLY7mMGX1DSTBo3jZ4MAat3rdNvAu2JzuEL3i8t4bbiiYaSKu7knyDk
FMb/EwsepK/XSJIMs1zcSdIYAWzG2STCT4prXS7NncufOYDyT4gLBG6ask+CJv62RUorygm/XdMQ
pXycLko0t60en5pn5nEGC0QjmBh3usaBFibuSLQyxvHQkl/4I6PhiWGk2o8Pk3sBXlJENdf4ZOpT
vnS9o2cZHTUNrXWrVvtsPpwd4WpOtpJXTcgeWbz2NIAcB5bIurhc3Vg6j2q2HKgf/xxnYwr/STFA
e8GxnVjFP+xQOQyuJfNElLwbYmU2XWTAJaliyA4EaO83hOcZhH0EVhxUHTlJkflksuymZDiO2hD3
nhy8/YTGbFIZXvL6hNlv5dAqfTTlD31X4fqlUw+1rcNUBaB02+GMZdylHqDr1vUPaGYR8z3a7Yrj
orYBcZeUAzC/XKFPyXjFA7AmjdM/Nikf5MR5IYP3rXcVu3wTSc1vwei8f59wKTHVlFkcDcl3frno
Lj+Kd2ex8kt8s+29dwyRF4fQQsHx64XU9kHIZPxUL0cQDg0n2HW8/tkzz8A+Q73E6qkfBF2WUA6+
CoFK+xEx0mRY4YuhFsYQRJuiLjRJIPlkzR7We4Sml7M4NSsj4ctg3ae90LJFGdw9jEHqSWaWSNv4
S4zOQRrNNE+mRlROvbvy87n/iS7L/pQVetBkjmJj77lRgM6J7LAqB88CzIwyfpdLFjmQTQljX+VT
EYjHg7pCI+5CN2HTjR8UMzKPgbn1LDcwdKI+WwJKslHvBqUgvfJI+k670rBp63wN0yf8QRx766Ne
UtDVHV61LdErB7J8IXNzzg1Fgi9pQU6+/Nb1vyUlNAl6e7THUMRObDrmf6QTLtSZwi74TQLbIDN4
Ah0AulVfH0a4943yj+YuWFOjXSjBI8tsslElCDPT6LmjjI2GBUmRlysmim8Mho/YtJtyzsS53dtM
QgYyFnzdX7fLL8ma20Mw93f0xReOPKThQjHTEIs95KNh3jSSbMkuvp3dXq15qfR+VZm9RfDe73ab
5EiGN3jmv6GdyIL/xfup4U08sMmudicGw02L3iYOvr9n7fwLWScJVTQqgbdMvenod0I7F8CW+/sz
jPvCa8ktSxV48E9/tywX5Qem2muXtRhxxJK05ryEYZRN1SMfNwOfbS9PdRXKhqnBjy/BLshdRIV1
ShK5SZ4DKWEYGE1/0trdAwLcNo6Zlk+pwa0HbAU0OExiew/Fh6cDlrOMYYTJpTXEUupnpMWRukwP
Yh1sC50xf7Nk7RtswBt16E9BsSDrwpa9MRaLHaG2q2MPXhemcy0HZiLsAmLjayIdu6cxUEjafYs0
s1e5kKsYT1/Qu+7Lxd65j9yoE8JES7ZAEMD4ho901sgVqcoXXckSgmh+nls5w0HLR0t6wP3qAInE
LY8C/qbtKBobWKOYaKunqueCizJQbzLxZgZZdOeHzTFsN2fmmGbDnOWwot6VMz5Wdae4LGeeBm1t
SfAVjUamBR5nzBAPF5mXJxp4o8VSTRrORJ/7lSUJTB+Q4OxgUuUmR57C7l0bkRYtbzOqIxF/6xmC
W892k8M6zV1Y4cd/UCNXZs43crTBT2M4YpdPQ0uSdjORhu2enJX3mWs9dC+X4tSREqIrmFG0udfx
V7nTV969PM2wQgUvqq97BsQHa+dbBPOIrn+Ez/cr0UCSyoL9WpEiDpWQ470gI+344mvsAMLroary
a91Jf8FooirDLpyMb6zttXyRUr+58LdWV/gr5qiGol1WlnfiRIBH/OtvkvNklzB6wZum1yqCE8CM
H/1kShSgjhrUhsGSMMXyFAhHaum6jRXyJb3hh9NIEH7BHaAKWs0NINz1lNymNLH3NtzLrD+V/OHf
gybH0xzq+nQShF9PWAaVAamJ76H2v1LbeU5SzNfcg5Xc/tbUWmpkxD2ZswVWLkN66A+5u6v9VBH+
8yPaJFYsNvpzDw5lNjxqrzjxhiynzJKQJ23zzbZCSU8ayqKOdisM2qVFgFamixJXzqzBKM15OfPP
4TNQfrq+uYtBsqIKn4+7lGXocsHeRjgynbSpjz588acwGQsHl9FjdtjbGF9iOZOKN2+pWL41spnv
8YGNzqhbhHn0bKw8luTs4zjNYqVQw6qFFj40gXGJdc2aJeWQ/L4blwVxO/SaZfdIcs6erOSn0Xsk
W3I3mTWZ/9mfjAI7+nDSjS+fnRP+sE0KhHeJxIOP620iduNXAhnf6MOI31uCqWnfQYk/co6+7bhL
D6LS4gutBZeDv8P1CiTNBjTnMYV852oILh7An8VVUktNI7IArofaJlvyxZODmQxthQeBsOoOOgKA
F8z6krGihpdJ65dboWmYbSn3KVyxeX/mW8YTpU7nzx1amjFPhDe8iIUXgCwa6jz3c5NpZIQyS8Wf
KOJfDFPx2+vvNqR/e1pm15X6z2UP9VUYojj2nIrmIrsJ6B7XshE2gsIZ7+OJ2VGxdeQjcwc/dd4W
KhNgMwWhB2uGfyNRpIcp77lyD6FB7O6FCbAbKaB0s0G/M+uIA2GW2i+zqhtMFiLpIPjLosGW5DAU
7ZzEXzTs20F43LV+NJH3qNC6ArgkSJtdYFj2dEm5T7K5rukoQG5+R+EJmYyYzrjVpvtVFAf5jQ6F
gFvhvhHe/OLfyiEfS1hZE5nzRdlvVVeBZNEHEdnlhUwMTdM3vatEgRYKlgU2GbJ2pl7rqGHfRc71
SybuQ+b8NBCoAo7DMoh/u7oRrFkwf1iHycm5Pbt4BEEFz8kkuXLp7qxMhH55lLFPz6FW8uI606yB
wKyy0Se4XD6B3YuIx3Kw2d+ydYGBrhQxMXx0p0HJV07sPk56s2e/eJT+kop6UefXv6Z6rRAQKQBQ
V9JwvmUhxLrR1XfYe6QOjytftGzZi46N4W8yAQA1OY003MC4VGr+I/es2/gNipX9XdjT4tvuDs0h
pZWXBPaqhcuZby+IqAz6Iyfi0p35hBXwcd/yLWRxVsWIHzclcfgkhQgLMc5hgwgQr4EIreymleQB
onfGxoVFD0TA47BotYPquPN5EPBMPcPMw9lzaX9KrdyY8SEbrp4brPibZW+0k+yFQVut/TfzKrMZ
miWoD/WoOjdLHDCvXHjG71ZJJTDr1/tvXZ7gkiHFXx3odIlOj/OKSLPH0I4YpVoO86Bq1tlM/VIG
Jt9wQD1JGJYiCd/sFIK7uZ15Jd8mUnqMefamrB6JwIxu9zG8M3PUWQBSA8oB9QwrxG/5QqNP0Ggo
wYO7qu3JGyqlJ/NQfTBluI6H1PipzSr5fvmlkUwtAIyAyBekSeQ5843rxvwxnnjbQEVsgQungKn2
tqZ1e7+ejVsYF4dihezRSFrq8gBy/wTqon5WtR0ADGmZ7yePazpIeB5uaFH14Ir+NGZGjUzEbaTl
BwmwYJlaUWKD6Sn3uXKx6JVZdgPMxSYKAML/Itw1q9h6ImEbJVjeI8kFPnhHNUhPoVyc1IC8BaFi
9bY5OUabERtUaSk+DQ9ycG78/HWR2h/ZWJHizeOVOMaRNkFgjX1O+41P4zyMevLA6KU3/gUQ/G6d
5x0m/hoiP2+0JgdZYXZ2a0jKOfjHTIV3gyRs5MOgqxwA7MRbywxir4JOYK+9ompaZpHfuKfPTJOy
VIJGDkojp6rG/uOhunr4kg8m0gvzvF3ieV6RX/V9MSFdQ6KwSmuMhrS3XzpZ7Gc3RpDfEnY1+BVX
kGgoWxNPwnbWLnAzfZdogDb/zkiiaqUqGIv7UpmDxv9LmvQAmWo+wBz9iHgAylLYqQtvKMmaMj4E
zBoILXe1GHcs7MCVfMW3fQ+sKKfEpHhB0hScUBrqxeXWxlAHahgpfQx8Wn6J9OVPFx4zMpVJU4NZ
u7U2vBzSBgNJ4cafT3xV6d2KmbuWByybqukvbq3A5qlmW0zL0Q5/tGHCiR0N7klX7IbxWtbWjLx6
JnJf9C2ZDMDCOFAE9lDYmG0g+gr2Rkl41Q1mk1iR1Rh7z19N43PfSzIthaqG+47sO5UUCwXVUpUI
EwKMwDqjZb6XVEZCDMP16bLtwVOGdWJDG/jm/BcNBX8N0HItLsw5vXS1COo4nxKNha+IbsmnaVRP
royDm+1RzvbR7c4Q1c5++PrqC5vS+Z0L3Y+5tjfcLWL69NAcmDNBxa71sptXQoRgByiamf9qIUJ3
/bYOSLUhUHvx48wp922fBR7BWr9i0hUV09fyR0m5e5LMlhfGpHU2JXIeGm86DCK+C1SqgsqFwxdu
cblJuzXKxp4hQTZflpmzGDHT7LVDSBD4QXQpQPzJvoq0S0JiwIDbN613YR3neU0FEw+KUXrc2zs1
nc0tzBPmma3kae78W61N1CzUtZjO4XF4epkwlR4v/u/oEJcWhBqtJ3Nv2hz+tMDOJjIcP20Ern5s
u6B/R1Stx32CWwqB5vMfXm7pX/3iqKAtU6hWhggqa+/Xi2L25FJC1kwS9nFN0xWXjmPhrijVkrsu
nq8KSSoC2ATSyFgko1ucp60+ChcNUALM+r96lOLpXsNUCRDLn0zu/V7eK+dlcwtio8JGHHEhMycs
L9dA+kAKOMjnVhb+7pgmOtwgXIRnOjreS7gQKJ2qzYaHPWyePx6f2KTwMWI8CFeVodmYXYPFsgz4
GbX6zVSYfaWX0XIH0B/kjnLM0mtZskPfxU2mFRkKGKN3mdBepHYMjuloBGJMLqJKrOniVGBzG2om
/foyJNgiY8+D6/6RySwz1qfQSxg8bCf5OedWG+NN7eCpJsN7OgZ3c7l4j2a8F9w0s0WVkGkJzEh1
uRzOZnFtUHnCIRzdpUgVE+wOsNYN89AasbEF6u15fI+tHgxJaXrV9gW+FG1aVJTbgtoZa7vTNvAj
QVeDA1M8LMD8DeKmmOANNOSJlT8IVYVDU/pDhR4hS8wxzl4HNy/efF1rSYWXxD4eZcCb6QYVXIOd
zkjtzHA3iTlCivxsBRz77NnlSOBA72vPbPxVSxMF0L5OFj8x6Kfjsgn4GkNHJg0/X7zPf/O7LXeF
gALJbZsJSKAMwCHCTjhOA2SJGTLBDkbrLABeE7bZSJvmRJkDlwcJANodOp23AU7DH7I0d2+4s/IO
+62JaAY/SUWYT3lr6kbYqefcWBeNDvA1pe/ekabaKwPB6Y8O9q2jJBF6LQtGv/gnTeG/8u6YxW4Y
kIsRPAKHi412M0khSW/S7m/j/pIo0O6H2Jqsy/1PM08WMCVecpYmk1q0FzYex4lz7qdrxTPRBJbS
gL42ql6yu2MAesio25xobohWHYvRoegsXWR3ipVJBwmoEvXSt9Zk1dnJvfP3CnUqvvzLlEZufTEh
i6G64mycqhYuPAmAwtSrB/SKHnTV9ocwYCPsNlxTlQL9+Vw4w26qTHsdjkW+uPk+wVkzOw4Sd9Fu
5fjy7SWRdKl08vGXLivecu6jiEp1mgNZ0OTZYnAfKgHwKjtX2ySRWzpavtWyhIWhOGRbRlpefJ5/
XCWo47YAs+unB2LmRHERXof+8PDMOsIXLV3KTMGrcWdFi4TmdmIERxuDyqKydSMvdrzKWLMSRkUZ
iWBJSl9SSo7Q7rAuHdz3jBzxQqTm+SBn+XFh4m0C99d9FPaJPy9+p4VsXwgvxbfsdGKmFrT657p3
TMkYjx8TtPXFef7ql0kzD8qg9O/3N50VamWnMCpEhvSZQgNEBnycFZ3H0MChBH+Ox8S+mT28Rydd
wGWcKixH98Ng3g5oPRdqU2oGqWmEaZY5MPOFAklcia0NBowAjko5+3Yl2t/8WLphYd8fOdyNrkMM
GnnC2h0DuH5xUTG1IVTy8eHd9FzbvgSHNh/kOiwd5CC+rlmoJA+STfeLVYSAdbLyMQMTZ27oziGK
DTWr98reWohpDOyfc0qXQ2Vt4kXAzFivYaEHFUio8Xn6sPWAF6kSc/14poEjeMBYFgokQfZIaSEe
5a+XeyXVpc+FjVs5oyVXPvCBNAED8xlhpgOOL3U0pv7tg5LWTHWH3V9D/CyOe4SQljUUd4EIxFOq
qKxumksaI//odO/2Q9UtPMtc0jQWUT1XvBSkVHQn6V2aTyrNRc3n4UJ90i/AaJxlpikKTDBv5zUS
Os+K7+R1LyggHDmhKUGKgTLQj9eQrHRf36rmiVow9k00qWGQhhc7SE6TTZKzWu/QPF3p5lYaML/1
PVgegJm6eXssGaJQXUiQJhHzq1n2DK0WueuqXOXMR6rOBYteHQ0vfuqL3R1NSCiyV3r93fpteWk4
72zxCCQm51V8Mtmz357Ra7RPX6kTGhyJ2ZiiR2kKTtXkgJLBkU9znH6+yfjTolo/nX9bKIa5LOFw
IJjHMgkRlj7xGp0lRJKnwbNCty9dcGq/2hWRwgDxJd5GLExQ/0ZHda2GiUkMi+gRqguYitE4Tn3T
6dh7ESC7CzpjokLrpo26+Yyy6B96m2/XDAcJEUNCf/YA8kUJAP+ThPd2M64HI9wndvgFLtLpx2km
vxWnsWOk4dAq+u8q0OtKFR9i4P6zcHwOG4qcXZ3Wwc9odEKgcttGewgiDKKE/rJAjdtcKvGZecSj
3Bm6of0IAd8GtZ03fFlb6Lxo1Ve0k/hEGIpkIoyHzYMz6wNPBG/z+NhuIjBqnNZrOwJGFwMIgHQF
GcUvRw7UnFkM3DMoHZgMyGDZCYuXH3tWWCfF3q3uwgitFLRScFQgPrMT0wR1HXvxJR9Hb0eUh67n
JhsfO0U1ZEqxFJ/Ub/oXEbe6qqI4qeO9XdrK7H3BtyDfvhppnnfbiC3i7+8QqedSNFUaemq2lc1r
Z1pSXDFDllwCDSlGuWcOGr3FR/vRJAOMGSy46qe67cvAJ97BytGQVdg7xODLvMiczzH52xCbNWav
IPTA8qphlLmHCgnqWU3xYk+V3tXpPzoUUOEip6gbgLHYZVZAgJ157AdHwDDLo75cdFfAW3cBa8rs
yOuje3DAm2Xz/v33WgmIQnOqurnRPHoxDtBh4QjgBlSpsHLt05ARO1zhJLm9udMEzFo+gtCHtcld
nPDNPGKtgfq8wIcuBF50srKjO0l2dugZsL/QYqsbiDDDnn3CCdLS+zWDcpvoQlxhdifAWibsZAE8
iq8ZdhgLzr70vIbx/8vNZFVRQoRlZ2jPs4tMOsmm8ZsP27+KfEJRXNrffHLFScdZZNbTJ4/Th1A6
4TeEgcmSAkqc021uI/kFaRH6jKfFYUjhXzl8AIXeBvFJDpzXymUI4ymEUvaBIL/I6pwwoZo14ocK
omoDOdvpXltQOmrb7WbhmxmtP2bG/aPIyy/ODScu/AExEEfY4qXPuzCSni3XK0jlDR/FHc+OG/AF
ICgoB9ElzvXBzpLPCYUNQgYUYduVQGGbn0m/rdA7WAIcX87MHReTVX5wdo9Nztxk+t/U0uoZ3j64
PzTewJNkhY1ylZ+Qa67diFBboMYolktTLe667wvpRQtnfxyBGeVqTdNWTXM/EsF/b9KBShBEcsOx
goHRGg4P6HDE3Lllzqm1NNzFiyq1+DyjlKj3TDc+GpqVfQxxDhoWCiPuyqq0CbiT7othQLhiqTVI
6A/WkywnCRl/kPl55JlT7E6x2iw9EAI2HKPoL6kPY3qWhuRECa5CTryIEJz+DNV24j2S0x77WMzT
/LubGUJJFhoIr6O+zexREy+gzbHpBbHtwF9KXqBZGdczHEIz2kH5lIoRUeXJ3ReWBzZa93d8svug
iS8XXGGUsGnlncXDS/qb1YDkz+JMZX+P5VgVo32CIV0wR8/6Bi+PbANyA+WptRnM/TEzRkRPtOGx
FJnMmKpUbixvkbTUHzzNdVijHU7Cn8N+T7K+3XyCRmZnM0BSnOcXjhGy/L44YIHk1yKAsDPlHODZ
mMQ8FGDkDB4FGAFq2FBx1N4/bKY/O71dZKrtuHr6g+faJV1DFSYYXH5UdHvukvYYtbczII9YpCoQ
sm2ViUTCYA9rSMVl0cZCsGWw+Z2KATUPqBnthEcpLCrR7zrK/gqm/mwiAA+WLqT9+s7825S3cmMS
oRI0DlnxmlFlPdME1ZjDVwE++wXAYgs02zTFTeAZojm32OBPXgsG3w3lsu6IzjpKK1PPYMyPPylA
mmZtH7DCPK46km1PQR9XEfNAZ/UDH5+qtmzd5tB62QIexr8Kgk/gKR7prNrNDAtnmYMSEx7XoRRl
4RL5lrR2B6LJj2Dqno20ZEoc+YVi9bU7AZXgBOoGmQ54xSoMz6dEeG5H+PK5GOWFOP0spwsgSPVv
uMaNDtWZvPVq0MJRdUgLVEeA1sOGQ5MH8Ime//2FmxKzUEFVEHJlCZ7kfwMUXgRbZ6LY+mK6LnoV
QnagXV75n61FMGf4zmsP8Mcp/cCOitLTrrDdX44tbMNftCISAMd/S+wBS9RPJHc191fEHVuG24K6
1SW2YfYrH17B/d3UkdODZzgMWtmidDUWPgoUuEmIs5/Io4ufyvtqN6kpg4JAOKsildzULnW7qWxG
qi+ZrXMKTOtrE0AM+vKBwRskGqsdnfRMbNnSEZAdMg2Q/m8/nmtRNNuawfwH9QzNUbFsGBcEvGZ6
FGYosws8Di9ukR0cWvrYXC5299rEoZqFpsxfXt5+ntdvNdZ4hJKTEkdlKNopXAWypvjGGQBTTXC7
4BGfolwZHTiOdXlt/Y0C60eNDo0OyEEgIjlf4G0czRrWgRfIEQ+VkQvxN4TnYxh0g83ePNePdFH9
keTk00+RB4OCsbyt4V1OlcNdNTEuuxFFInZ7L7XrK/OY2mOij3PAIlhDMjTukB4xyv9QDZFhSWBH
dPu4wJhXEBnZX6L/DqSDyIDXjj4PXvaK0N/WRJxoHdYXwi3J8ZdWGqd0tUNly+6U5zudObUQETkp
2mmQ++ONkA+CdgoxhHN/aYnvO2WhJRzbKqquxQBu0V0NA0mtwrXBD7D0BjK3G9UG9dwEW4qcCKp/
/bWxsLcl9Wzv58mJP+Y8vwiYzJQvGi13K8e/fheO4Ygu/Bo2jSSdWR0YyvGToghc49MKqcoQkY7c
qxVIULTtOO3Ixc/U9yYEFEQ6/4qcX1bo1Vhl6pXaH9RxQEKbozGOyFBaUiGNUEey/7Gq1KMy6C/o
hFTHl1yZ+elg9/WAo0SCVZBAuYV03b8MNa3vqZoYsl5MNcyljKQTyrL7xu+1XZQ8izMn6z5USrHp
dv48favbtrY1AWnrSr+4rgUwjPcC6ldNrF5m0cYzsO/OMReSSlQI+7fhloJTWVbehDgGLKztIoJC
31ZMm8nZAG613NdR8FIRIq7cty1eoBv3w/2eWE8oLvMvvlRQG9PaI+pUKjag7n/o+CZ/AgwnHEYP
0b4cQFHBbWGuyb+9oxr8Dd1/w3AR1LOh+4IjqXd+u+TccHmRVm/02eHn1KiBHlxFYTOPR2UbpUAu
6kkCV0Eoed+AwRAxGpkA4nAvEthv5B5jNoF/VvkOdEQGkOvxcliiXoQDsU7tSc0/djUIYsFS5pdN
En07F4tbV+KppMwkNjlMSV88vLf6eC49fz0Zq7dL6zRBSrNAecQ0vVjY8B5zEvT+1smseHqL5Eu2
S0LPMc/nCOftl6hsMjJa8Lgtf749rrzNBzqscIcvB4zCN9lqJmJcN28mfTUEAzj4Itpue3w1UvXD
C7pSXx9VQkqaw+1nXuA+YUdRMgGydDZUmcSBNdmtOax0wXPgp2aNSp875AcqvYYUUfKulX0p5fZp
N0mVo6cTgo+pFkjmGmtX3z4jktsGaoTxrT2S0uvd4pR8/JPOa4Mt9qeppmMOyNUQ8bJMwuaEk7wi
LxSfezGdbVU6fMi3RSPTsEueZqI6vTMr5U+kOt/ghpmx0scka+qQCtVcwHPoFEPBDPyG0N+NbiQC
cHol4paCn4oKOtehjXKV6NgdCncnEEdLt6+IRldtnM9sC88MAZ4hufudcrq6LjBTx/5dyEHlu5jV
pIH6ir7P6ego4GX4LcpoQmjnAseSuhD0x3KuBKSRYfaPSTeVFQsgAk55Abg/W5zT6NHr7hH0Dzgi
WP1/pqxDK2T6rPST3Rkb+MJSBkBdzwkvQtp/DeWbcK0+s9izpFTPbR+NipseXGP207rx/rRZxZRd
cFqG8AxGbYajLMt09pKbzQzEO02U1RJabu0X0Jc1r+RafbeP4KGKg4Ma1k7P/K8QAoQCGfZo7/xP
tmlNljtYOkLefsPPdrCvva1aUl5CeJgbUEoeIOkExlmKRQA/E66L/BbIplc2/PgjwjKAVKcBUrYm
EuTkN+oOHGll5qUgK57P2yG51OtdOhhUtm6nFvUrN/nKeOEt4S2ch0XPVQCEHsCN9dIR/y/ljp+U
wwBU/BVIyittUshpo3QHsK5VU13nSnMVbJhO7Y6XJxALy8n5Elib1ncMSJFhb2tkp+/DgT44BV/k
2kKQbR2FcCWCvnSRhFGLSE7oXH2iF/o5jlfb/8Ue5NGv70OjiER+EKHmH7CaIrcGFb+TAM9fSLIy
q/qv/aJjPcCSo9oXyD3SzYXXoc5f5GOpxgPiY4Poig+ZjzBPxUa1mn+iHgU/JukCdTIvmI+6EDPN
hPWL4Ev6CzaOoGgV//meRX2lsMeEH6Y4m96syEG411rdI/k6NoKdqPrdZCeXmM72TrLNlhg+x1f1
rkWEXs1KTyLESxWRS9N+TxbzeHusCmGLHhAE2MjiCg4lh6Dl0PMd7aGAQioq4qcRyaJRpL6lhrPr
qwwWKXAmCK+w75kH+rn7J+4q55WKnSDGilw4uWYO8iBDj80WnuXnr5WZSgzmS1POlDVFIkJDR4Y8
fr+CHTh0oSATkcvvo3pAfmaawZ3ptR+LQ+sN7NWiHf8volSmy3kx5k+dkODMYAnHHrE09wL5pDho
9VUUX97lEKsl8Huu562TgwewKRiHATR/ArER9I83ng==
`protect end_protected
