`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
dDfFWED029WdtWwoRwQ6TauyaFaSQWE7Mt/lIFbwzX/lRxdX1a/9knOlJ+AMbJo6v9crzaqyOG85
f5Ru4x6WvCvJPCj3ejUoloNaJUgjvHr1pTeLBDwfRa8qDsRwcHGebEQ0jruXd6x+HZKEYBbZp3C9
QTa1mSfl4sXHN/31ADddnS3tb0gd7qM7Np2Ou5FdCm0V8bewdOy/vouVCWSm4BtFGemViy4xFl7J
IGmiwvj40QOopBCQ01gPDaL5be/S/RwTsswqSpjbTSlzLg+e7qw2lcKjXtBaPAH88NZMWG4UQP4J
BkkKjMRCuCO9S/0P9qSfMQF9mTRb1e3gIYO++w==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="Yis9II28X9AnMHGHycjLH+BYv5FHV40nkBQlrPiXC48="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 104496)
`protect data_block
S8XhrHdSSzlpL1YZJu/xul8Om+JmMJBIw8l7J6x1b74MLF+501nNeHzQbj5trDZWk+PTgbPy9NdX
G415tQl3P1EYdjmQofsyshaRQcbnxWygk/NAzPjB3mRBbs9eMog9Q0RaRqyQ7s1aFGdBvVMqPXzi
ZPEuaH/iAYyGlcD2fN4YzU6NbEFDJhIZwNDHaxAHqH2kMrbLB+4oa6xiNTcEQyILqFClnF7DFDYg
9SN+3gdzOTDyubLPPP1H5cMJRb0nTzuuPT8m1i4BvTHtikQ2PkEgx2e5sJKF1NlCzhRTb7LfBhdg
ORlAbBewpb5SJincYlVYzvly8P0g3ICbBvV+da8vmKF3YSSeIV6l+b8bwwpYDBOAA6mdDtpigOiN
xs9+CJ8VbUCKCSmBmukiGb0eLNQ33kZCA5n/XPS+Cc4p7lVKz6UTfr5OuoomAV44gSPrwuxorxQQ
eif80OaGz1FISzcbfmptRUuFX9mjczY37nTYPMDSCSCpKvLqTQEjQRR2nQKXM3ssGdfGSaM/R7De
Ma87XR2wtwMaBOcBKeOioTdBLQPgxfTJxTOMav3o8WOS2HCJtmTmrwYcyxOWwR/d69v4yde2SlOg
7MEMsyuBxlC/L4uMY3G54w+iEsEXvEiXubSkfGUkT3Dtez08YI+BBJ47g0RXOiewzyNvoS/qwlmv
v+YLKFCausnNT9Gr7Kqs+U+yQvcCqp+ciNs7y9hbHXgKiGB4MtMFuzcs23kTGkEeCphmEI2BIRkb
L0jy86fmCVN2Dh8CjocDG+4FO32M5Z7cB7e6Dmka8w7XUl99dKyMY7nRfxdJKr9j0gblxcxfVdBG
htXgXCOUyv0IsJryj98Y5l54RNpoBe04/w1Oio2G/LIrJljrn+6HmkljNDPk+50bSx7nRJ9u12qs
Z4bfQ0zGnQSe+oyzKLrmnZFjHXfhcrliNZiASUnMO/IIFFlY2ykd6GW3Pjkwe14w/J/v6xhx9+kU
5mLleUH2SzfwYmzmMExPVqArG0axbJyGxugAsccBNGkaSbKZ9gZKDWsEAWtuKXQUK9ohwViNNmpK
ABCDsxkEp0MksoXaxlHY41V04E5FIrspMi+tcnVnzxE5o41MW1ijdau389dDVzweZD09QzMnTFgO
PEzbGu+A64qJNOCDzDzK6YkmvKcEvl7OmY6HeUndkJkxwNO/i5KR9h8qe6SoRFK+OtlWKDf/zsZU
+8ccNmW1EC4p7rmS9VsPRZXL8WV4LE3oflc+TFZ6K/C3II3T/GAoWO8K8TSCAWn6Dro5qQLPsGca
wq/1jxL8Vm+95oDmaTrccot3r/AiCt6Sk035r7gjdM7QF1U1ZJz4sTsWl561RHdOcReBSu+xejnL
K4Ry9a5LLfUEG5o1aXQxHxdmFZpTE0dCs+GLfV5qIl8HXdSP2yTnhdWgJeJQ33X6d71d+oGyJOch
Pa/CtxeTMrQAHjHcscar7wyitw3nVDYMDAJ+swu3Lv6UXRKb+Ye/JLwpAI0oploxj1iOeioNy6/a
ZgNVskUY2h7egxPl8k+cPlJgeJ1JdyZMIFhWAxjhKS7Thbi76tQRpjLmtJmb/J3JdbJImxWBhAvq
5nvyDsIGOvw1LjTuzejuS7KodUN5gbDoMFdIS7dka9fQXZGcJgcqrcfD1gTx7KgMxNMgTeE8H3Tm
LkUNNGJ2114GrjcgR+XJ5YjPPtLVqBbpRBtLCvpRl3QaaH9HnGCVP7Mnftl+S4E7GjYYpqBwLwue
/imVNlI/PfogqsQ4ip/vHRksAWHh5cDEZBltVQ0Urb6Xf52wMgELnHaYesGHpEMSR4XDJlo3GZ1G
t6hffBiv/3X1KzQllU1NSTnEBP9FrYl2QnLyXT4QcZx/nxSDGIf37R2IV4r24NfT6nV0WmCpBcDS
fJwrX3gpVofSwOJIFUTSvRrbvMjFVheaTw0BTJL6yOzlt3qDuOlc4wE8T3azkN6KMA2KT/vg0ueW
l/s4Adl9BsnQhfcW7JfEW+/CVsIO8LrPodlJFPOUT9StF1Ao8IUPN73Z9kMdXyOcnQAlOQqwZvXk
j+p3jTMUJIjAASPCdliV0oG1oMdthU1fz4QGS67SONWRZAnC3KN5lgRVzHwYyPFppm1R2lOTkOFF
O0W5tFiqJtZBpWgGI5wOyskl4BDjJND6exDX1Z5hdnrnKoqeauNsIa6zYJWqnVKrpgzqzVgAhOvn
3vMkApXgDCr9xqvD9YqOSfNKnaUNM9PU1KLO00umY8XbHEzYkQPPZSRT5wSOAkSdvgIyKQKBpUEF
Sl0Sh/AlVu35ShR5k+pwaU4dgfEOev8NFLkZ4gjpcAC306b3l0nwtqvleEVQucRXP53ZOVggcVsp
2zsuiRUmAuP5q1jlySZCF8T+fuVZsPKW0antTLn6bC74ht2WdaziqcMbyeLV4rJThWfsZ/kdfRxe
mcNiG9aObfs3i1PLDcEFiaPRsaHEDI40n48PAeevQQUoAB8OYNEe6MYHZJwwB2L7QqJwgoCPd5+0
lqXzP1y4AIdg5GfyqajNHLZN3qB0tGz2h02ySAU8veThJL/9IoZoIH2moQZm2Qo5AwM6ANQEpRhg
oNppKPfiSJmPt/o3Qn8mCL6h86/SMbkpeoxnmVaE9nRaG2KdnDOMrAfMrOlfgwmAZctPvOszbTK0
duf1NDgdYdSyHVF3+ohpx/pV+2qi71p9FIc4V2fj1fL1EbhZx89JUbEynV9+FIJOMmGyROhIOVPN
aVxQwq41N9U5NHkf0s9/xtJxUe24kDz4jUz5jgzkLEljdn7HAhVwAf7TGp63Qxk2rIgezVFQqyVa
8vUY5qh5/MpJSto+hWRTQOAk2AKycYxveEr+3g8ZMYDZqcbpCaLyUmjRcHgaIVQifel7EejS6l64
iLYLlQqjG+BnwVwuRzi+64+ysZ8+4sOthcbjJ8inyVHr4Q5OIySSdL+SsOEKbvIpnEJ1FScdtjYq
xQ7sv3fE1mZlitQlGtH2lep9l51eyPBo7tifDKLlPSNORgU9ceG5tg6Xsn/dc3fkvug6Dy/8rEBJ
400BbFNL3a9LPpynjp9ggeGighNHDgmF+35OSv8KfEPRdxiplVA935taNdhoFw5VA5dnr5udA59n
+jmMEHAfSYjrE1VJDL0Vp65T3mXk88SCqoi/uPH5VyQw4+MTdI1ToX1B6EPqnfFNqmI4UAi9x7/k
clhJzIyTrlSbd2L0jyumekQWqL6u92UWfd/xDUm1SAN2cpbvs73YO+h5kc5C1S7lfYIOQK1amymt
m0Zuq6cc8ZQL0Cze+352lHEouBMY9H2+cGaOIzbpXvljp7zmFDVMlOi/ovxWUX6+J6ShDUPUhl6H
9Wx/T7rbjDrOXtnNTam8EtOG1Nl/SpvvbamS3Lu7IgxAhyfE0Sc7uNKrTO6SggCIzKJ85B0qBN8i
gQMN0CgZP52upDGMxa9VIdhxif889+pCEngTcVU0PN40R7rRxQTTIGea4uoVld0b7+SG12NV36Pf
bObjkuTCbTZ+4xT5xj+K8JVON5xXjNdnVZilVNifeFGkDMszHm4GCRZj1bvw1U6la1rEIZg+X1Qg
DfJrXcUC2GSzODdSBlKxPn648bPT/Hbsk3JW/ga+hKrGWIRRuDn4xI7YUkhUm1YfKpY8+qUEcsJP
gSRRcguCA0X9G5U20Qs0Xe40UmGNDQo5bs1J+8S6KW/vS8ja1A8Cmc/E27OKKIlOQya05c8Jqn58
XunUQkJD/EuccBAXSQFx5xbRMm6ossq0XZiM96qwKJgdRd/9ub3u019mlwacHtEP6ukxfWpNkMpf
3I28VCqZLDJovNQytvhetvgptYzJXAqsfNSbFX2a6YeFQtesCC6BainY4KCIuCmmT6kvrelhsO6a
Bm62rhu+6cFDxMQBMVjqgg7dBuRN52qV3JMJnPxlKQnlp8XvxcZGG7wOyB+weIYpJOxkmp6OINZZ
FlU2mI0I8oHtJQrXFotolxcfh2GfjirpXObKX5PpD04/N2M4FA9Tyq9iYXkI2Rf7wUpFRJd1P0ys
sk3Hers21j9CQe1l7vYxGqfw6dmoi3Isg8LFb4Nt3ANcQUmqIcxiLrZhQ07F1nBDqrtXCB/3Sz8o
A7Q7QqrJnSn7Ey2dvs7wwtEKO0tguLMp7/r6QPMbJpf5vJdjqdn+NXDyponMpLEL6itvfK7j5967
zv1DmNHwaF4yZc0TgGOP1yxEq07QWDOZZgiFGtMyTHGeUP696pG1oFb15M8DVpzJiRxuZI9xxiSJ
zka3Atne7QQDAKIh47NvLlVcFX3jXD9UWjjuERPWeDPSR1cAv0p0owro+0VwwJxMJ6ZVbs9pNlUC
Eagvao7j2HhFQGK+F4ZJ7Qb8QyovkIL9qq8fs21q08k3P4mJJipbSoHJnekzXUCbM8IaX4s7mAno
7ae3ec1BzMQ5B/CQ+rMUVvC20OAL8GlfHEOX4EdE9nLLrmdYIZnfVT0RBV5+36ighGYsx44J4OkB
L3rM8OArbCGBqXOCjoGQpfw/eF4hLTkLHvojYx3uwDwkMjlxcif8zs/VEjJks44KLVKP85n2n+CG
svLx9m8PTQylA8bPFJQIdsBQFNRt4aMC6T3fqeOPyEoHUGtteVateqH1CmKACiMkkaMVIYII9iar
crIrwq0Zt1Ru+Nx1ZTg7WsMMHZIZ8GYxn8YNwXgqKM59CFl4inp5rJAiYLdM0sv0ytHjQRpNfO2F
gTPT6irulLYScNCBbV3FnhJhua0SyiV6dUZoU6cXMadaIKI6guCkKCJMAtMGIxcoNR3Yq66kpEUD
e1C3RSKO8lt+3WBPS4qzNYLShxyxEXbd6WN6lCHRlCWTC1pkghn3PGGxFjgBtdu800WpWeYEnssT
cGiLeySL3zbil3uOkyKWUOAY+pX6p1v4OjJ92/CDx93ttn/LRCkM+sGMzRjxq64fXqYOUTLyHLQQ
uFnrTcMn0SdPfRogXwDmP6BTlkvYkm3Uf1ziTG4/hnrB8abOoQQ8p+zNvROkNosK/u/RZakPVvJU
UYwcT3Trk/pMsfFgS6WN/6eeYi3TXNWGlEU5iiiL1HSCQTtVsX+JZshr+rzD+z9gnwqx0FUWkfBp
NAKEvP09RaDzwyhFYryd88PUtgWpiKL8WJY6IdquWK9aBLOiXz7IdJ4pHP1RHtfq+8TmgpK/cHhx
T8Ckw6RCjjBFAhQseYUJbnRdbIFrjPIQwvNeHLoxW/1OgwG85bTwohTS9jbPMHg7Cd5C8pL9p6up
d9T4Q+/Sco8iKWRrEvwQb5FfmbeHa+06+quT5avLR5vJfhDXdPn1xIe05FLCtgDuXR2+F8iUooRQ
f4bbsIr9AlMcuZzgiRWXUl2hZ52ONsQPy9g1FtOZXAbCIr9zbUAnSVSqfekCDig5PEwTgP/IlQAl
qmmGEdk9OtPPMiAGZdmbI5jqSaphQD/pHX825MXV3QA6a8qAslyh9WNx158R0AWW21zBcP0nskws
KZ9fBx/00enLVTW1drYeNTvhFhcVfjFHcZtAmJ7jCMPsy5Y3LiIUEsMfFzDVQX1Rllt8Wlr4lH57
3S5o/6eCo5nMIjQxE1uwzzshqkYtYLFKccSdVBWYT7w7fNYe9QC0h5Y+Ov2JDniXFWJyKQndhb3b
lIbGsmjeoKGIBL7bolIITeZlFWjpHuUWBKkWOup7oIEzHoS3wJe9tVP1imoCRTPr/52JCPwzRw84
6HAtIKJxz8TJvVL9+BXDI5LCIM5hWpzk6MM62M4xMoxaRE598OXUeTtaULb8w4dYY+DpiyY5nKj4
DCXxzWnK7k0IAKE4MaGtp2YWvfYYJtoCTkeUFuerKBAc5oDjheupLTMKRNJ9dUHB1Pnv+VW5cXUH
MpsZ1sagJSk/HOsQ5vdbh8vOkUCB7tyc0RMZNZIAoSf/BlwlBUri55asagrfooLiQkKrYFGNjnjm
sLMSIpL2GjQp0EvepDoxI2yQeLWe9+HKb4lzhq/QJY4yEjN7flekMt/Nbryr1L3sh1D/qCwXBooq
+kaA6t6tXa6gCkgC8kn6y5kncMNmYbEq6BBWFvcXtRBTOdoXIqGCNkYYUj/c+R3on9PZftCJGmtq
vG+CbnMpThZfwuwj9dDEkmu73KoUxXWdoL6a5BxT9nyMjAt02ox0UUsMK2DVBwKHzJSlgq4ACVys
qHczyq4xHbQaowzA5fArZOTQca8O4kcrv4fboL9ElQjbek7t7SHzprYvPMH18sFlEB28U9L7Ku4T
hoiH6olmnw7d1xfgsuOWZiZuyIC4FNZT/k1KNgGhE7icnJjCB7mu7enDg7Gaz9BZK4XgAME1WVov
vMrHzNpRf9udmG9oykf9VUp5jAqPwTp5g8N7i9CiNanYsG2cABDHymKzovQe6xOEQCvvtkhiEjUH
oYQUA7IFPOIz3WC+Eql1IGrUvSMp6qP7/dG4Rm4EWbskW/uzZlYsh4/cNe8n27EGTfdWVrKD8LJw
gcehKP+FbXTuyRHFqp/pO0N3fLsFbH8/AZK4RF1B71nWNl2P/enBDvOyP7vwVJwJyRo3i5jliIoc
Z0yBA0qODp1iwSiP3gOFsoXykoAGXqEcmhFUIGY5TuvIY+FyfIIA7nJizX9jSbVsfZBIanQLO5lK
H0Upv1isBBIeIJohVXeoK1B/OcIBIf8ku9ct6E0ZB5/1TJADroZeHA4q74U6WmgKsVPFNO4LwppR
f2q8JhG+CEGTLViA5yrXtuAxXfg8T6681bMB2byPGSOWtt2GQPnABcrhrG0D3won286mAnUoCuU/
j9v/j25tQSdFozH5c+s7g4VtjYhSJizTQpi5V0G1KGZeFWZ/u628JUXR+xElIT43zOWaBSp6iASl
ZmKfPfy5Ecm4oedRv8mQYSZVtRU5SBOZsKdl/HvkVwlh3oBdiW7+dGdzugPfia+PIUh+iZZfmZ26
y+Gv6kq0mlIlmU7IpaXdW34hHN44Zlxc2YB2Ym1AUEz1o9O7YoTP3Ey3ysx4LsLXV2dsatmqy5do
AH0Mv3Xi3H0zyFLqyDNoSCuv12AMuMzU6/6CcUIQ5ot22rKmlZJtgy+AuWQKKB/BcaUsjC8ZkEwB
cE+IgSlJRjPRIj4v/rq1GsbjszMIJ47Zz0GNtkCCbx+UMDZxS43JTQ/RChBEExE78Z2l6kkau2mL
piDY8xYNWX3C+zAipi4muM5U2usFjlj4Rh0QOieqT5Yy0wW+txp54cc86dH6MmbS1UjiDr0p5e8i
0WagAb8DVoJIcdCJfr39DvL+r+3dZJOCWwfAOSCUrP28EcXTkgXWW+bhLB9h7/uSJiNPg38E4I9S
5CyXDhK3zHWpJBwvMo/xvle5us7OYsShEIWjtE7UoBPO0rbAv49Z43M88KISBAE4nt289C4PtEWP
qNzOwqKx14qKEADq6A8PQcwKzrkMWkXAd8t61tue9CAUhl1+rfA2SqSKjxfd33IU6PmXylAXTIoc
suEmZNybbvftJ/gD5MYWshu0WxA5SWZmmuNq/kyrs7mEWYGzBqyKq5+sA+DXFmxR5Wl/bdsfnD7z
MkmXyw4A9f9ObUW13mrteiwus/w6vo4K14giBnZZXGNsUVDBmsyORa/QIJ9p3iS3cqqdaMa3CKl7
vNqVZxDrh/DM3VJKbFRwhI8pkwrDdDeUEDGJUdCQBaOuEV0nZbRfNbtLuZuhFnPmr6m4/8BX830R
jT8RwOyTtxoOVWy4/itapI1QhKshLEqWeLNa7BZ/kjh9NtMBSEsB0uwbuAKvXI2uX97hG8FrZdEY
Fgc6RmpZEJLBrrd8YDWgSIoOc5ubhaPaZd798NY2CUndCbDQIdMlEATnGTJH6OLlmlUNT29uLgyx
heQtD+F+hkjZTlTAeHa3d3TuR8+UoVVHfS0XBiuJd2RettyNZHDZELjh4ICSFJq9oXOjUpyIzT4t
+pbvstnM2xH1kWWajm2FWKYYcy46FogwFRVIklaeTSv4lyaInf7yBoeHWq95D2MlUeK+7q1pX05p
Hu+jSToCAZutdEa8AoNTbbO5SM8IflzPDne7d/a7rAzvzEQgwdfB7Q31zgxiOgI0hsNAxh50xzlo
M632g5NEIztA4gD6uK8lMdOr0Mnik1tfyQIdoTM2YSJb9sH5IRvdTibzPra6qaLEmOxF/fEzZZML
SuR7bOZ2OXB6OTlOqs3WPHlHbpSlUvmsOKwZIsqmAGhQ328FA6Ml7XArOnlSyl6gkK42Ty7wGJkr
e47owT7grAYRsG8sSurlJT4L9LhAlkdGF0euLwhoiwlHey0pvBLPdKC68QHdAKWrpQRIHYGqK+SW
eKkxfTd5hiAgv0ZxYEOKAmxnJESP8ZgS3T10vsC7CMewIuvrJqKzB/WhyRACJRayOF7sg+i0+zMP
iTtD2GM65s/wzSQlztLYyQvqdzYzsK95wsoiEiFhvl09jK4ShAVZuheHR8a5EM0GzJxbwdTDbAFL
ymThhlEro5TsoCZEC/7xMiSCpxfgVOBIrZbniKS38Db0IIc409pjwBtc/adw94hIrjP4Jb/sMs1f
EHRIJ0o1QChriMQLdyo8klhOah66o7dOrLaxCuu+6Anut1d3UtBTr88v6hz1DX1MiMMOKZztK7qU
eZZ9Gy9e8c/3ulZ9ctImZYLdp6tz9uTFEB8nVNNLsmuNKi4r7qCWp9WiweylGnhIMNJ0FMOgdWTp
h6YkN04DqWbOOvb8SqYwaj2+GcofY3636Oza41YPzdAcDdXA+ZkZM3gk9QGsWRxaKTfEgnUFCtVK
Kw6m7ns5dW8QJFpJALxoGjJIPPEsMQxTIKURO6uvdewwVQrWGOoLj+lpaybdD32/t68K0HhOZVNC
28LJN5P945nmjeud8spxnImccOoVaAp5NmplrbduhSl5VqlrsyfoQfKMgts1pVdeAN3IjpBUPMN+
zw+cRkGhuwZ8hQI0fTvb7qVQ7b8g8CrcmpGAijvHiC+ZhqtY83xiWUIb+b1ca4XA1SU1zM6dArrr
teQ/A6qmj3ii3+vSxCTB8/BcGQGglgooOUVVgieaPye3vCvFx6NXFDC524e0xi6HW075riCUpDav
szsq7WZIQfZmaPv6VClLTg6KBOzDzFc855T81q9nQ8YkaL+OIAhU1EABVpnugs8oPMo8UuEKuWVy
/VD/ugjA9FQk+ItZvBGyxnAKTSK4edDu38Dx3TDL5h8xcvmnhqCPs12TCpww0B28vmgpFbOa3l1l
2tPMiWjpxeu8IXXSQYF8FQj+b+BXEu7OaOCZRIZmxhhQLD5q8Z6xMIZZ847Eg+041zgSm/LjJZLi
Yfa+G/3nmcTmeDm3s/yiEADwG7M1rZOSOc9tU3ckEjKVi8jY71gMzGkDCFRPjeQQq+fQ94Zz83M/
D1ujGlMn0TA6xbKAFs0MLQ7sv2sHGuGBJ9BNFNmJbop2K9Efu8qotI6O1/2q5DxjBhRQ+ZRghVFx
xLBriOFJtEVwrRzFiaOI15Xmv7Ji3wBLIWQhaE1FpqVO7MikY80s/GFAAQikWBsKm2A7O028lVCZ
RBKIZmBk76VIOWjuuyrSlzNJbaLzOSGgafTyBsCCiXN5pK2nrNe1CVK+MdKB5LJM2QoI9p/ZTHUA
5JMQN7rUyLwiZdax3Kkb9h3R7WhN6MypAxRu6jT6yQtsPm8OyR9DzOVOW86bVNN5VC44i0Ea/uCi
cvWBGr0I07n9+pTjjSuJCN4r20c4XqCdnU9J7TH9ebJzvm81HRD7KjHCZH82lpFwDHGOSYDb2Ykp
ZYbl7f9XIZwSLmprMhHrului7USaaCWrhE2XGhtTWVSgbOkjhsEYzP7jNSFoXERMXxl+deg4a61F
BeIw35eE5QDqYFHL5s8nYDODtxiPqGSgMpwI/HWIs2oaY9ztecm8ynyDkoV3TIqzym8fqufMd7ly
/QwAySfcNqLc68NBOAhiJMWFY365uRriDcN5ZfkrJiDBCfBWUs9kESAg9B7An+Dbzr5mHNKmyxur
Yj328u3fk8upab9xKY2e14mg6vW7Ge5fJ2xAdoyawIgnsOJ27+5JWDcuAeuYhCTIAT9W6R4LlZUh
qf98FTAtnMwo58Wr1NzjJsTkARhao2ugx67LGiiXQosWtJNX8+xaGYSgODoCFPwnewGSAwBckHss
0SB4izIM2E0bMv7Yp+w9peY4wVIbXJgYSZ2Ir6p7yvI3ksK52GMriiTKx/9SqeIAuoAfAfkxrn58
0zAeqK2I9Kz0nmCPcSIqdeINz9w+D/wZBycHq7nuoXiTjnq2q3CR2mppNlyg1VDgqmN8rU8rlzr2
W+bu7baRsVhG7jOhkHakX/K9xcY02y3fNI+U8WzmNCLjSttKSLCKqQ6SIOEgttEF1vK2wpQ0tdfL
ybgIO2SV+wyweG+KRBLI6sF/maJxSphVp1S16K2vrUnbMLwHA/2VlUw6QgCuSfwxS6XeFkRQrTnt
ktmGb26QUj24AXu8E1bpyy15RHrtyiwSLfabM8ds/SxS2yGnFDuHrDyv0N3tYoQ1pcBLjiOGY0M4
cyuEqFl+d7DVRoCfzwypnaMYV1Bt44inFCXfyhBjhNHG7LOlgZnt4yY93a6Xu2D8s1keLFS/sdJn
V3EPTRRTywfvmPc0Ob78Dh7M8XxanWCT5XHXYWLySy+pCNp+B4kWn/vrzXOkSOqlVKPxv2dEBsIY
DpS4XgIdYzg0H5cpLQuLZ7mRjGw3ED9WxxWR52uxYIomESal9/Bs4Dkcr2dI/DG50NJOqE3KGK5t
NVW3xFCUks5gdAesGgCqfsX4pFYqOEQVbX9OQnicaXPWO8bJYXje2hWL1jiyg4FHnd0F9pYr8DSX
CXZ66++7JA77mqbglZZHD+J6IfBrVqzOgIUmpZiYs3UesrV4dy+Ew2ORF+YAfGqYCfgKViMRqMhb
2JMwzME1RW6HntZSPDN7OzTiHUVvVtc1t/UJHJ5V2tCAbQRAQkdDrLdU6t5aOyDFqaVNKZGOyErN
Ac5m11eXVRg+/YAk2KZ4R42Nd5aLfsBnl85xv5KEhvrfcNcDeM4E2oPZpdvAnvZeBC7J/EPUwSbV
RfoPKw2Ma72dAymNoDNcl2TiTOptOrF1c+PW3OtkdmSRCDHluf7TunKtCNovPdint8MiV8grUYGl
QHnDH7utT8TmUOidl19CQBVq1bJsMjQbg4gYfHg3HVuQ2yKCOJJ3DxtC4DSIejgg6we8uEddVwlO
CFw2quRbYze/1/TcG49dRw+ogKL5blITK6XwTpgku+dQnvCbt9yvLAVe6S9W4cfWzoum/cA3Odde
UTXFkl2OpYiYN5tE0jLFh2IBUmjDFrIeBg2Atnd+i3D+6I+D9ZIMX4qfXzY3KAwy/V1FFlIk8pJI
RuUn5OqIesVf3qUnbf1ExK5ojm7cw087OHc21AzQf4PRabhCpzGDdjQNppHo+7JzDTwK75VAvzc6
GrivpB6AWFXmG9XW0PiHBWMsDNiGDBRko0LrIwSUQN4/QB8ZXE+uaEk1SewMCoxQzyQLDASwaVI/
Gnso7hj8EKIZm7sZZDuCD6PqM/d3KgTVzX3yUc5IvQS6830VTma3oIjdLczGdFOyhHFbbWfbUntm
TKgq1WCxnXJtsALaXB3elyxTawhfTvaY4Hg0aEv7AL0ccSiMJS1hY9iYMJwzj+MO6F0CSt0V7W7/
UuRicL74Q/OGjpTk5XJS2jCMnb8gt7rCFeFlDQittKvlxAUlfI1xz0x1QaEYIRGHqb633ut9VDT4
BbRtJ4VPk/zTF+PEaW+i0NdKXSEerGNqjod72QYv/xhH3d6Rs1a1y/fqlRlSj/bHud+KBIegvSgi
sL5BQt4dw4Zrl2YMTL88Ml2s1tHiKhQ6C5ZlyZr08LdnYn3uyNafxTTeEE8ldGgm92rVHJKtOBDV
Xcun+F6pCYZvP3WYgyT4J9cbwCiBydbwLfYKY095TTYDQn0hTFw8dyDAoeOUXBBiajBdbvUzx5t/
pAvgTVArU3djg1618NlyzWCenMwvJ/iA5woJhlLVFz8JIGfii9ZK1F/ZZWh052R4PM+LnWMj45es
Pn2M8PYPs7JboZn2gj6C1eVSlzZljTZv58OL6Ckh+rzNMiqs2xA338l+8Me8BmqocQNW4nPGf6TV
jnp+QKuJeL9mwADnnIZX1vHubqIDHsSfcl7c6VhfqLuDCehOkuLn+km5smJV2MvW6c2HQ+efRj0Q
p05hoQBUY4ajrLFCf/Rk3BVSkn9rN3BP6gdap+J1BxJxfZpfaA5bUSRCnifLHFRWSw0oHHKrinOY
rBBNkeg7ZFnU6pjeXLMYwjKirt1DKlFgnI8+4HqyZv73LvfIeD3agv3K3kcn8dEa/ETgKfwCU6Nt
wdBiUHixexd9OdQhbAJcFu0wbihuWL0stjSotiGO19VhubVbwXQ0AhCdJGVXD6wwZiXv4GGGomDR
+M6KrslBVQTfyhiZp+/TmadMkP2SDe+P8BhNbogPUV597QeXJmA8ouxOro8FnWaSHO3Pfiu5OtiX
5/tV992tB4bzKk7Fbt6kV8cKqLhRMYMacnZacEnDxJ6VzNft62DASnnv74ps8mGPzf+JGdz7hlox
1qmtSZLc/IoUhp7PAjtwTUU8ixLlDZm2VpD6Mke0Nka/15W8x7G/WPoz0N6fcGth6jkObwI0ceEm
MERMi3YwSCroPRLrPYmiSFLbVE6p6u3f32FLA38jx9wBV+pEbLW/zDqCwlodPO3RIaQj5yzTlx8H
Hy8ODZdgKlU6pc4LUZ/6MCpfiyudZKZxn1/Dl30UrygRB2P2xilSxCT5nl/E4U/wJzF7Y6mEH0ZY
LyynS3WlSRlSpazAnzKWYnGcnbAbeiwbxSdx81Brpbr5ASnddVF8rVYoneVv60Jopt8AF6nD1643
2f5Tr0VHO83ZPlHD8r85vIgxjOy9G1vCNFjMqg6/5C2OxXXZ77Xvf+cpYTe01qgmD59vq4E9VAEA
KAytp4bXQDzl8+junG+/Qy8vL7hS8z+N20wFGlLzX4kO5TEyhOgT8jU9hTvxlZVnIhiOFE23aU5c
fI7iwvUZPbEEgXIMYWAC8r7q7mJCCJSlv0LltaodKgMaQhX1ioLdGx5asm9ICI9Zn+sQhM07i2H8
5iR7LbeX5zEOPPQ5cwH0sJ0h+hBHrm3lwa7KQczWU/ilzsZcNKYuODksKdx6ZrTWJY1HCKzg2r5s
53Fj4g1hDHyfn/6YSTBEmTMQ/WwQJkQFi/JS0c0iXm7YyVs+GFOBPi7dBiemP6XL5D9RMgvnTTYo
53vEsmM4docasdPF6KH0LdEs38MiYMAzhjZA6y4ukgZxClntsI1jbcIefUxWBtXVBN4iWYptEy6M
hRdflyABJGcFAPbqOVJ8Il5eH6NvIoP6sLXgGa/x2EkAxdydgr6EubsZGbPx0CCsZB7uHbObU9Ve
iN2L2VDtPWj15Cj4nut0z8DSqK0pe/Vu3kVV7C0KLAeyYEyGMSSCckf/gxpr0qJgV9bPGTs4+//p
9X/ledf47nN2PYyriRo6JnhoOWyS1QUd9/KwTZPwF/H4QGOLSwxsbLWTvJy6OoJW1cavfAWnt7Jp
o5tJqoHPeRM3mY098oW85jQIQf3a0pphGIjiy4mbon89qMNYHW0iDsFT5zgjhtiaeXXg3j6bB5eo
0GwEXICmcb6r3LLHWAiplSvCXi8vV9D872YzHqtDBmL6F43n2zQyDaBHM1sXLTkblzdEpwyMSKDq
Y+mSlGRErxI67psdXVuWoOGnyQayoJSPC5lI/u43b7XEjbQzv0DisAL/ZfsJyTHHFgq/+05qdY+0
ulHnyKs9bWQc7x21OorWJGX+27Ku/NO+oJKWRHuNiZ4lXcTzt1M395imsYa3TmTTjIuxs25odSCk
GbC7bmcUrrAOhVG2EoAt+o/3ny4FIoBbwO6UsJJxvy0DRvh2q1zwT56OiG6fOCW86sZphCaChX7l
L+XUE87YP3TdeI2CC3FZNzEF2sc533Tqhl+kcPfJx65UDQ1qzSqhAZXGb5yXzeg0ol7GXUH8Hgxi
4ArQOh3HU8S3Ouc9qdqrJoffEveLj44e/VmZ0Rz6a3HDVfGzzo/sMPU/55LBnjPzS+W/vtkf0gQY
qTCYgnelSjKeONxS3uoYE99R6otAmpHi0PLNGQDc+jJtO6qwqabMjEa3DyoTxvMPhgsV1jN+7LK6
t6NHbTCZpeL10rnis6SUgevAJH6RJU9ZBvtldzYE4LjH7stYrh1LrPLtjoW+A5Vm7f5Qa9bEjn70
JxQHl659DgWrXCCAesIPNyt38THhoO4suEGEBZSb//HoOLHf85kFDqZJ5xDlksoo7WSD1RDPFKU/
tZ9IyD2YaCaK6fMUNpnLFAff1oukLS881JbIYr5FJxEfEWDQ5sEOofEwGSe13zVMy1tLKjki9jRv
XBiJTa8RUhmDTrmCCRCj84s0TaL94+d2YzYOrURXWmAUoOqzJmohDyr6kvf6c7XYp3WcPH9rx+ms
3iZL7vJu32e4KqQVM9eZaOcBBTaYJ0DzjHN3TGAMwmzG4FOUcjqHFcJQtrexQxNpAiECLqcxf0wM
TxlHpsMh6hmxyGs5hJfdoJnhaYC3qzhuuwUt4X/ZucHfeH7nDlUdCeT9d+pkl/I+zOLAjDFWglnF
QimkTwiOo+kDL9kYnGnlSVOBgRies8Hnjgp7hrFR/Vcwq3nJ//5//h7ZUotZ8bPdVa/5I7wFjt+x
A0oZR0ogXoDFuI1AFw//4MUHsjNsSZtoa4/Chbi5bTTG1+pZaqw4OZwtDq894Fqg2vnLBXfbgMQk
7w3V8jirWtu7+J8c2lMQZ6eTVAd1L85r0faf17QhptjSVQNkXTY5sOp2y/fJVB7aaNgq6M5VtGQ4
xbVwfHrDa+Plnb6/a6cIoT0cIwOE1LSBC8sxQ9+c+T2SCG7pk6xUCm9QDkER5Z3uOKgog78/heJc
hORx4FnKI89VneS3vLMt1Z0xummpo7b7gc9HJdWZjySxeyNcmr3D9DcqqufJ8yW31Flr2/nPQVo9
8wFQ5ttTB27uTNac7W+vY7RAR/ov4d/lSzWtkvTVxHMy6spXnPjxgLx/wjdk1nRIU7gErhtR4g+J
wz5tIln6RHgEnH2uZs0SqcjyKR+pjN6hUim5o/1NImyVW3BDngToPyC8jkqyW07pXTN2k5npiEC+
bRMYAgTYtQ8PRDdOIAgc0Xc3yd67TBTCWy1xJZJuINRqZFMlz8vcvSsgLXGUMnr21t7jczqPHcRe
ofeICtl6JZ0uCG4fLDDUOK9AvK2Yso1/hcnNdTbSzdh8epQFaDj8rNuQMvRt7g+7vBeKxVBHdk5N
1R9bf+8BLGMVbqQv8DNdTsQLiNLhByFPwDgAMxO/v2TGJdSOt5NVc6rDVXqvt1Zdr9OjhNf+T5GR
T3jQILF5EpGlMiaXbHE4B2e7lHTkFlMywmveQ73A71hdpjVlH0Bl4ZpzibAoG6zMW31SJOMJV00S
3imcQchDDpUMk5k+40EOLOJrnu9BnLJzDjAvy9+saEReRyE8Rg5oqbq97yccuRjatdGNXqXh7YoH
BROaZRYldic8w2hFjXyxpBug72232pltCkLG7VwSJIdVHIq51mm1XYeEsAdGZBi2FESCGFMqd1DA
HFi5b9rbculTfMIhFAXgd2M4Girg48jh2PAtX5SZtUzRAhtau5VRYI+vYtHOt6qWIc7m3JpIuzin
4fk+7NwyX5TTEoWPHdZQIEBMpvodNmqvqlyZd4R3d9WSvF49NHcMAUFhZbqzq57mO5riOo0ycdSM
aI5xNfrwQEeqvsKg5J+ffphrwo34/bghN7o7UMdK8VoSREf6ijEw/N7GTCG0pjP474Kdat7YpsBf
xGtiyQb8nf5moN2yXTgbxXtCf7+Kg8XXRhApwsTYPAkGgqNpYK65hYFQnIW+RboK+7r5vQyI5SAx
c5Mn3GC1oGmhiMdSuAF/gBcpEAAyzVzfsZkD8SP1a9VTJEEt2ZLl8ZuqVCZ7xMwefrj0GBPCuxQR
fi3blghIsMVVkF9t5iJ/s1mCfiUdpjtOuc1f2Ii5PymvnMzyCbZtlBOZgobS8ysy05lC4mC8p3/I
tSq05PwT4PG92pWAg+4CgwIvZBAu3M2FbjsAWzi4UFVyOx9bi4HdYFXHoGsDI7ULntjF9osyCFQV
MFHX7NOCbOrItOwDdlSB7xFzEEJGiW2oTYapoIJ/p6YrFHQra5x0s8DrVRoMftJnmIvqjlFL5+oI
jEvaj0AhI4LP88xkTjOMSGYtU17Oe/xpcoTop2bk3BYcqZsDaj2OYuO6dZUA0C413hswRzARDpd5
bGTBH0PR5Xtk/DJIH7IghAG38qdSqgNEG9d5Vx3T+Omq7chxNoIhAPx1ycY5uJtBpGNL7Ze4vEFg
okOi/XSi1zolbEjGgMWGs4+h/l8dc2OCIyy7bpVL4x7El4sF5vWfliD781mZ8qp6jZ/SyerrMmZn
c0jOcdgXeIXrF+aGuuP9f3Fymx6vpLCd8USW2xHr6uJAri7KqgigyjPK8qLSfkz72oOc9HZ09/0Q
Q+b+5ieZZdUEvfGs/90SvRnepqhNoJVjbxplJ5DO3mJmYvlMkE5gboDhu+z5pYO6g71P5pBDrNVs
LqDRr+zTLef6BkfO9QzyaOYXTyU//7hpwfR8sro8wk7a7belMHH1z7RNpML0TuOggnnXCb8jLBGO
DiCwq/KqdnZptv5kdH2prdLSjwoa5B3XL4G2Tc6SCoxYVt3EVob/RyM3UVIAPCm3unuP0i4ZKs3l
8n4lQ+VV8COBgiu14oM8aqJ9bH9aTsdhAKahV+A8oeUdz5ltiJes4uUOkpELOYR8qNe9Emw9mRGV
lNKd+CBGp861eX+wTmQBi8M68cqOIb0rhZUfMdGLM89UXNCJ+yAqPj9x5q57wA0iPscdiNIfufuU
ZhTv3iXZ9+iqfhroBsqK0YzasA+f7GDrgK62pA10JiK2GqA2q6vDgbyxdJZZTdQNXvE5D6Yl99kp
/l1kyFNx19OsDhfkVVSxIbeZIpNcKqb66OIsdl4HfNsy05a4GaxfHfZE1Im2lK8/LLJneAYgZ/bx
NfwBmc5seM8YOSpeV2j5X29+Ghj8Xa5MUYj/NgEC23mzaUt78itiCNCeuAw3FyYsoGUFlMulcZz4
ql4lGCiZT+xiJFN+rlKhSyWijGapgILSPM+IXy7kiRGQyoFD4ZuoNge5/1MWSXiAB7+yqP6mCq+3
GT+AR8UQOLR7itZnp+Jv00X2LuLbNO8IfFS8i7uYFy9pdGJHUu1rccnmkqZO+UVzsqcx7q91QtF2
LCDJJOXk3jOUHasAT19AvofyknNJu46aBOIedPWki7tXdU6/9ud40o2Xkld0lspu5a4MKAt55guy
wUuv04UoCbpyzCxoriWYax8q61tQIFUsR3EwCkTVqrMq2nHPOeR8L6r1wbz0ywvOnFRQwCUdXNJL
7cuTqtUP5WZSwUIHjbbj73NF9GNGbFIogH3IXA4AqU/ZMqIS0nJEwpIUZSRSeRHCnlXX4fDDQAav
TY5ipOf0Ra8hpoutwFYEvSf1nYbM2kjHvlpqcsq1myjBaSDIYsBl3I3SNbBgyliD5hdab20fHsRj
pnUx/xkoHMLLhy2luEDHTGVNWFCZ8BUmEC4K3k8Jyhx2oh6THQswsCdBg8TEs2rPV88kxWY6Oeza
gRmNU9fl4aAZrsjnJpbW+DC8G7tx/Pv9Ars0+XAY/u68B935NngHumbPzM48RT4gDW+AGOQTvBoa
QEqBR5n3KXwqJVM5q/9s6Txy7+OzRNeXS/FEECzT/w8/8Qezbm2uNnN+IBUvaP+kHz8s9Q8gIpg6
aEPFhXkU7zWFMC1SYVeu8NNeUL7nvIDbqDvV7cYNAy8KwWi4D5EQn0ojtB+F8F5bVUvETdtYS+rS
cVlt2H0X4IR1M2LtqmWkbLASI664a8nf5QjeSM877TsbQsGKsw0D6X9j1kOlOqr9SPhheaROHxRM
M0J98FCyH/61AjPIRN5ame2weFIu9GMtAfDUFiw01Wo6sW+3CNGfWDXFxIPIFOnur3jte8CZw3RN
nFk9p64IDCE/SASG6Ouv+0xBYISbi11+fuGwoHtIFyirJcz8Ulr7e9LMqJUZv+EPOWoL1JzW3dIb
S/C4L/kixL4aSkfwR+5OzO1prYlXovr78VqJUl2hBxdIjqfCVSb2sEIv++6bt0aGVKImrSyBILH1
7+wEwneBsprs0aVwEvb5beyH/jlJP5nuWbDBz8Oc8v5Jqf4D6H1hDfsijHKnfIIU/Pib6QOX1XLL
ZzJzx6ItrU14801NcZJwOReiblSN3qS+HfndV8GTP2C/u9ypcdZh/Sp8NNXO22FPZnlVP/LfPScP
Bq3iKjP8Tabf7HJcvhlOPo3geA/nRwKuJush+/UZgYgzCySCZlOTKu1rPg19Ol6BzKuAHwAqS80V
vKjouSvogLbpAPB8FCZneKnnqQpANrxcjN5kuluXhMeVkHlcDYt4f5meed3YkAYjEqmBuVJnNvVz
tDcJwc1v31XhrPp2w5/qlyhtps2VqKrwVB04GuHtDIS0C/K5ANXvBLeUHqEyt2k7qW9hA/mk0WoR
XcxI0/aPaJX11KsgsheaGX2LKmAFj7q4eV0rnmKLDYEhog+eiuJxzzKpEIDOt8VeSJs0WHqOMvvn
7urxkZaLIE62bK/r7Mi6pH0ZMcu/td5ITfvcuYvSIsNry2+c42c5TEbelTopSiaaep1MhVY8q6Yz
xuFoum1F+sWY92JhlhvrWpjnWLF/Np5FwVBHFgpqLf4WpFyfUOteAyEPJ0vjWDOtFZawdvm0sHMC
zlvfubrRdDp2vjhYwSeKhDOCwmZgjarluHytfaaS/EKtrE1bM0WbQBBDgwLNgg7SnQH6BMp+NO+Z
kN0vS5EV2f6EVjhJINhGeiZOchTXVZ1ZWmKiQ3lBDgLYl5i9Dg13JnwymnYabU+vZVzP/kNZNRQN
b9MyToUCanjQtnnihOMcVqXaGfA+dk4Zv2twGFa64l129uT8oc3vaeXCtpEGC+Nk/TjYhK4MaZZ6
UahgTZIG+R/Kgmne3ZpMsqApbb3YutHBbI384vNnDS5kXdsD5ftmJAlB4q60FUnw3M84wmHyLFbm
3Lo6Gwx5pqR3rr2z9/vJubTUUMs64NX8Mk7Ac87aOeuGoLLWrp2azKBaOWS7+imyF0HV8e4++Ji0
QUIcdReKzX8qHrDLmThWvGttnZFQLscGHQmlRnMr8moWAXiZBaJ/3qHx4Dm5kxco8PwzDkWJXYJH
GhPXtI+Lff8TyatWgsFmhsvZtgbeuWlKY48IYUHZTpoieWrsC2+4j3RSbfxQJyks/0KCSuZ9zN7v
FiJPquZNPihTPc8niVPrD79XKtXA/aqu+brPZquEcs6x3EbMuS8MgaJZU4t/N/DlJm56Idb9ci2F
wwrDc/SI+LI5qVv7l3DMYT2yLyieANBdJh3nrJR9fAuyBkY2/QVo1qlkQc1JF7kt/BBi34DQUGd/
ti/uFw/BXpibMVtAKCWvqArec2bVBNfNPnfvkHxwYvNZFdewOj9dfAkx5AdYh7qa5PjSJ/oTu16J
xI6dzLIm6uUKUhsGYR374JtVJBQ9jejj2WrU4IjSCPqxnsfg7B6Z5e82v388PhoRNA1xjCxy14oV
p+2rccYErFgY4bD0Y54h2YZ4SVeyJrQimN9rxxDX5n9YNGTVjTa8qHKgQiU8f4/j8bHtDag1ur73
l0jiv6ftd2XjdS4356CucDzMDLTuAvAAZPFFAJiYuFNp14hZBEepiPXsFMd9h6HXqTZOSPJpeus/
cBXSXWO1ofK7M0YljsB5KkMCmobyieX86Vxw51cjeh/zZjKvmT2zpY9KKFfQ96h1KGoe1Kksa6+w
9mWCAoALWrUssM+HTZFClUV8t6KGUBVZa9Y68cuygUQn755bFCunMI8FIX/qrPh+scJ5HDLlg3LK
dFYJAVWNfoO69bDVPRCGJtDyua3Wb9hmgU+759Z6MfnVqDFK+VEI3LReqVIiw7y66s2E2Qfb2fDH
r7RiC06PlWoQSXtwos0hU5aMjyMDqeWNNgPEqb20iJxnNMcfTa7tYMClIQFXC4ihU0MJMrDQ8xwK
GGP2CjWq+YqYoapBwC37N8T5cVL4GC4zVcxzhw6gDO7s4HnuJeHDaCFh9+vTkpbMUhnTRR3yoypj
hT+gPXYGiNSodukAefEPEBzPkbQ7veMHyiGzuKTc8LInnCZsyhUJ6RyIxn+CgJCTdT+2dhesFdz0
LjAqsGvq/UXfG1vkQatgIH1w4qNrbpwEBSR6q/FBbs141KnvWfXAHyQSLgVT9rTddDd4tQnCg5DE
f6snWoPMV4Pbq1d8Hs4dUlUMD5afMEQPowCaYEzlfY/hHbEXpp223gbNVq2IosnI3PZNTwDWuja8
nC6Xl4+Z+b9WjCEWX9TvV0IlSKI2wK5JAZRL8rnV/0pZQwuk7U7OZ0rVGeKo0W2/IazLMNvXmvXj
/Tr4zmghSBY4xa353VWEhA0CCahmnh647kY46JJrx5K+F63Zn/Li1Ldd28z72B4kMkVKZfO6EczD
jUXR7om+2UVkIIKiw6GzZY1gV27BtkAxaX9zGKJddxOeOkWxZuyfYrbro9k9gRU3VTulTjbmkitE
YnY96BQop2Kt78RjX5muSDSzeP/StOXNjxbkA6PaqUaVerVu7KuHCRBXplDkH5DmANk/MXlrFvmU
gRmmTS27epXZMD3TNj1TAh7YacTIJBM8kaLe4ZDlsgZ12z/gJr+7OiYlBdAaofB++ME12BoN73ZH
9NbcKKKjCIlwPayxWDeT2uaY07N2mFzDCyvF31rhOVxUw1rBes3bAYcq7ezjo+c+KsFrQmUD1LGj
gyMwBXodkhw0bEsCy+Q2xq9n1vzuKheYqP2+fiDhVh6SFjhoAt0BAlFFC07g8OvgHBu6YNE5+s3X
e55/wDZ5OFyboa3/hDkanhxHfNsoVZqWwAqdoeQZiMFwbRQtgpDgy2KLYS3tCEAXBz5Q7l+S6icC
tUxUAbcOAiIg/ySpa+OxWS9Uy29LBOwZEWRfzKmf2nDpGJalW1rRhwE/aWJfngofJa26e6+QCccZ
5BElWWIKG9vnml+aJNfGWPNnzXWb8GMEi7WhlbZPPyeU3rCTlft+FQdCP9wJRPY7D5qW0t42OqIW
6kWD2vQyLcLw74P4Wx3tz0BjTT8vnb5q43bqgjJz4VttHRGTWVA9OCPMcFm+xuGi/euAgPsICsv+
YaI1Q4ricVcpjocETBYuOz/gpTV2PkNQ497JVI8asWA9VBWDF49OQh3FuQRJAN3N41a8tO0emAUK
jWjiInHOfKr6kvzKBtsoMO6siqzMP7HKly26iaeYVxO4k7lrEp57ex/4kQjoqr0OTRpqpsEeXXs3
AT+wvYlHazli6dbEjSPCp001Tn4rtHDm0w7iBySGx5IKhGgQ+PhLoKuvu9/NzMwEYiqgUbboF44V
arJIrH6kxcmjIowGvXFDwKSsEhB2V+J9l/OUxfVjnSwoKNBn0GBhnIb8oNRhw/9ixCS7pZmBHTiN
Abt/WwQD5JMFsw4pZkrrNfTL0rFI4JNwL0yhcOiqFg86URXv+ONbSswpz52sef2atuOAs+qlnT/g
n6xazdVWPpgScl2G/hPP8PKVUHoXEBu/pbiuOoFdQSr2U4COr9hAn9AhsSMhRAPQ0efVCXc3ptUH
7cG8jV+2m9/7CmO8lQXRPJSRn13MXE60Hb7RAbei2YLAMdafLcny38bKqiWDif/49WRX3mFPlrEi
677gNT4oYxuH5mJa8heUximUZewK9I0pNbh/IM7UBgFdjHSeR2xCjdye36kjQtetoXWa/jZNGMkq
bA+7Wg4bzUQ99pYWA9LC+RxYrhXd9V9arQa+DegWHQZTklx6LkpYTzZwHtdIdt8tzxpQ/jq21txl
CcC6hMxII/YxreszxU2urRvYDRYaPJZvF2fI8ECA+zXTV++yvg919KgntiznlPyK50Qb066ODqV4
nkbKhhgijNH0RyIzTnQyoYpRS9i7CxM2F3aER81zPPYAlvT1iaeYaOQkK+hKpO9PfcZsGNUyvlXG
9TUrn39pt+IvT4IvE/ZuNfMaeiYmbCmeZx7/kyXVI/rteZs2qNdTmdUSiWnqavFlq1a7lNWYNwUU
XXPU1ldei3nyQ73EMH13XBLzhhhHNmM1QjzJOYicbzvmSavbFWRsowW1uy0CckSUSh4h8DVDF2LQ
TdYo4iCFbu+rciftyc26yD+C0bGPvKXTxvNQuyzUEi+TRE4SDz/XrQuL0o/sqc6Lpr9hRFfXbVqv
LQ+qw4VsT9ACAUOv9WZq7aOI9hkhjo/ZqpaDrAyGNQ0HbAYOo9dqI3axalUuIZIdQB3d1wBsws7r
9/vOfd7pKuuc3iUvTmfnbpinbBBRumZV04d7uMpNBocxxOr/Wg0cV8hbC/f+aRIg6Dv/F5sBAjX6
WYe1/UL51KA3ay1t7f/NkqEDWh6sQGm0Fg/rqYPnABrcSYeA9iDvDkZdEDUBDn5Jsg+y00uSmbQy
uVJj0He8yFC95eEGBIvE9LVbBK+m2cucY5JrrKORPf7xrvDumlhx9dXaiYEpDEAmXTXZuuPlfAse
DoXJlt8M610ALo37PpEHMLz6j4OindNn7Ge6vmvywvBmEQ33wfKe/V6pcpX9vbodxztxxwI7USNz
zSkNvG7qu9YqVp2ost5tGo9gOldq5lMc6ja1ppnQsBDl7YSvfKmaVzice5Piy0M6xjdxqHyE1kde
LVUTuy9iJ//0Q0JTy8OY+4hp+0L9Ii+1K/Xng7RgVPQWj8fvwyGmHWCeDlFpJWIhgydgwVwaO+HL
Av7nH1+ltANzbZ1ikgeLNLMgORcIzxjvT0ToehO3UDGDpKNNGNek7qP+tohDfUW5nB4Uk5XFXPz5
aCUZZ3fHFX+0DECupDoYr1taHRgUK5Jm88bIN1U7nkwHuX40QxKSq92xgg2ZIpuTOZGcrIcwaXRo
w3diKzzppXcL/jRnVbwyivPVU4RzuW+nPNRHjHxcRHmbMFZU2A27YSfhw00i6/wpO4+4OqlNjYUo
7zaZTDbvRjOWwRGpu7RtGr8AeNQs/0DGf9DD40OVDoIp9pWa6Qj0ZUqNTC5zOxXryMVIrIKMTNuI
IyyeSrBD3Kj0j3rmi/OWzaIWJ4CxMtgfZxIrRbh42LWZ1bSJadolMX9ZtJWdyxez19VECsu4GFqa
LJ55kJ2mVba1D/KtkELeU6Fhb21hQ2GcQCdMd1LM+bnRnK6j0QdmoRLa/Tp+8qRZApCW8cwIx0R7
QrrBIt0tNVD4a943as/RT6oXPnQOGFs2NjhAdIXW/tqAQNb8Sv9smzlDNAlGMBMvrGc7L1FayWV4
tG6fviyts8jLJHOe6qRXTEXMcE00/AhfBCZL4FjhJwRIHiyjuHUHFvGtS8vfBZMzqGa2uWl55j8Z
GSaktQAID5aYGRBykL6+14okUYEfQDzPrul4Qnr5tLLMjGGSR2I76mZOY1Mzauws/uIJKj/acYn+
ZG2qiFf+ggFBXRuOQzb2spfnCVVnE3bLgkTTN/TUpArX7Al7lH9oMDZxb8BYy0wxIDFB60Cze5X0
kaWWcMTb+JzZckcUS/Hg8uS6xXKUv9paHXPeZgVJx/5CJ9A8ghEoWk/rtF7euyx18d0mUl1DGW27
NYZEDdl6AZnUtV7fRR0W3qQumQxqY/MJQnunBiZCnZp3LiouW6eae9SGh1UTcBzLmvv+kBzXeqZa
Dz7LtMhqq0c128bPsPgjuntA92k8GvoArl4ThPSADRdRCssKXUfeX/WT0K22Fgjjuxgtd5DY1wN8
k4SWFDXQ2f/2upWlEtWEWWPWBnC/eVnqFyR099/iEjICfhU98Lu1a9DaAasFVcZz9zcwzekfYhlU
IvDE2uHtHgi34U2iknADjt0ClH6cVn9DTxRmRY6XVBsibkWPs8zTNC8JlFUB/ohQPxoqJ54oFeVg
tFNf1nJBA+uQ6n0wQTYbTbd3gGZWAv791ZenK1CP37PpquV/xls2gaCVQIP3/a+TMMdZZS8K8IZF
R6MnxorrAI+ouM8Luqr0DMWHezV+ZvaAq6e9f/DweSlV1gJ+TPILqitkQXeYb3tcXqlc5T7DoSMN
ikGcV1lWh+WpzUHAFtXhG0/9lLAX+ejwih161dH2eCM7JS1rRDLnpJEmkioErXBFCPzf+b+etD9F
3+Uu5rcNeMvc+xUpVlqlFPSVBuPn7dxYBdzaMsokuuNrgFoA91+LHSTNXdFHMzPf8jPlpNbBgdXg
dSR9kuukJW6AEXL4GY6f6oqh8kqMUbZVsrUFgVNqUp0Y4aFtCrUa5HBDbqX5/fPLy1LZT33CNP6B
xrqwHlZXmYwMmGj0jtcpKsbbk0IA3RyNkxI7dDPf54QwTU5p7KPDj0DtgT3FAiTLVL1LldTb5sgM
N9Qx7jyf8G3LvVX7AnSNTZVJ+qBtrnUXJxY/Nzl8Wo8tH79NInmvftEmD8y/5KJ7MA4Zj0DuSAoK
/ajbJVHa7iff38eoE9lNG/jyG/REmpIAJgqvfIPZBobU8hVIWiWgynz7bgO8LSbn4QoT9kKQ3Hhq
IsuZCywdOdqNoZiFYYEWLCMPCWM79m6saStHlBumY8O0ZCb6u43yWsdFAdx/LRznNVqqWjdeEn4N
R5yoO/yv9bol3tbjq3uKbteY/r4N8WyxJa2VCoqym2WEFSrj9L84R6NMjhS9X36SEWhfvESJlU4d
0nU/77cgQAeo6NND2M+enLFr2bj2ULBn/ks0URSK41cn+JR0xzxjz6iC8Qn74R2Ou02VlXqv4IhD
27Y6z9pgob4DPIJfdjUdJK8y9iJ/Y9jconm/dzpPVgduebyPupMjBZk5cKN0ckbOLL/db+RFDBjb
35pzbjB5YdMF7rZPcBIeSiIunYy4wiFp4QyvzOlm8aSuhLVQ5hsSLDsVcGPK85tBGnP9IuvI75oh
9QQwXuPJysXqnmVeh82zHR6t8/VyxSQwiqzlHshbjPr5Hi1DBJdg+qGMCC2OMGZIaszH5TXtlUXO
LRCMfpxra1e8twpG7auJ4L0DSJINqX/P+g3CBcaUH0Qe9XNIfaXjD+Ao8+cGDpglVi72FGOCCDM9
k0UAMSAH6kqbrsR5ecsdVbtDQrDRc/Vq/d9IXaxS8Q6r13zdGm0jnVm5mEMu/f1uT6ZI/N2xhEI6
riPI4F4b03pbIxEqCMdRdDXTo346cgL9FUNkj3gI448hAwGeF1Glh4MGzZdsp0VnpqaF2wNy7MeI
y0xAc47+y0VIAVPfg1XjJxc0clAIPpgYo25FDbfPxJSG2HH+4+Ag5+7jifnulXRPxCrenLEyt9vB
MnVOvju5NGXRe2ssXjXjk20g61ZPXxvSQMFPfjCbOrLfO/YlfBv0/Oo/u4hfEU8Y9wUmZVY6SgIm
q59y6w/5QrgdU2AgcxX4XVCY8yJ6hfg3UDN2Hml0UP/dfrQ2l8YBgCGc7PS7G5zKv+ijxjJEe71C
ErqwbXOXhHxczP6sp/TvIm5TC5V6b6vy/bY/uI4s5tccvd7ThTeYEEhpIzcDBm10WmgvOrFEi8kT
q5uuW3GclgKg82hs459a+XLNaROykEeqe5BC0NFSE4wqjVRr/fb4Z56eTNrdemwnWOdzQKAPnG+l
v8LcKRR+kA/zc3eTmwdjX0XSAzbTwr36bP0RIVetsV7Qxxw+dbtAe4JdaBw08oyZLAQuZneTX32V
bzGtc35/w7+3JRz8z8ktNxcQ28dBy2OsSu0lwkeO4nt/tvtHZOKmEyIX4BcmmNdKazr//bE+kWyl
VWi7kOxrrwV9vHMTvQVbETT16Ju+gK2u7Bb/ZggC2Sbh4Bf7b8OPRDutr9RYqaNp4WRtG+havjvv
idicIo+auguHnazlkbyXx+2e+oXi7q6d5kPuVe4A9Rhz0lOp2COqnIrz47yOBMUNr7+wtcV41rje
vOBEV6OmKA/ugLdVXb/pCvsQe3pDIvGjaQmengCO10F0rxPBDgI7ubYBVsoGFrnlbW7y0o5OoZJx
UpDWiXbv9WK7LJfcuMNOONlzi/DIxa8K+2SK+xKF2pRpZrRxqMx2JrJazChtS426eDNvbIaSeJ0Z
XpzIZi5s9+YKxXkQTdc64VSEz8AxLLdeufKLWKZ8FoqeKMkauHuA0/QeQC2vZ8H8+uVbyMQH8VCx
TtUKMTBytzS9YLQoZKZ1YdmJQyt8X+BRIjn3i8h1KfdXcxz/yJl0U4pM4XQ9w+lp2CQ59HqcV5c/
HT0u8IL3OQW/4ItD9XtOjHR4xSVzmNFBRO2AHrrz/DZd+Vo/NaFgbEDewBtY0Unn7ydTmEMyO600
9YjIfNMLm8AQrw7/iexZBsSpYT12a7eczSXi/a/4+hBna9xRIJwiZ61xKgPB7gOZ1oLugI4WmYBr
ksvFRgIa92moX4qTtMyKHE/FOpj7P7SLy5DH5k/7jNs6pwBV0xmaXB1C+gyANawrHHTH+rsNCqJZ
VpdL5A2C8mafVRDxALqJ/DaGC1ZxnYLm2dmvu8gm8iHcEIQzKF4lDnMZuA1O30Kt+oTFS/7f0YGc
AHlNaFy6XnUg60pxUz2dnG9Kt1Ohj4DP43noF9qHlTNhB7byHsDYj7vGOoMwI7oa38lQw6aTDITQ
5v4sCiJypWClktW6vMs/H4jViB6jxfI6E13Fwhkl7V6E0lO8AJlhZGbn/m06NoCTYDbVVECyEAq9
YtKdncKxMt2z98xMT2I5Zh7sTr65f2kP7Zt1v7I7wp+bQiq9LQ/PgJBa3McY14ij3qKFF+szJEX5
DJiHzE1Hl8oJL+hvUUKPXVpJtJKYDi9PJRvqusjuemr/F1d1dGsIvrIzWeyAh+oNNodAIn2jCteb
kymFhZndgsUszZtPu+CbJKACA6NK7m0/1JoiG36J3nOw8BSThG70n5QzWCDFNVbd50qORD+dWu1A
dGBYaUdxCXROajUeBHk3UuWYxAyd2Aa20Q4ZNPIjv7g41SGa21fsB3ji6M1CXL8YuSy2fjcSquOo
stGqMEqwEkFSe0Fha+dNDMsC3c/9tKwTFa7AxeqYdgM9/IUnuYaMzr/bvnbOBUpfP1gxtI6Zy4Pz
MmX9nKS3ORmHQPgn9QccgDpr8KVe0MkPvySLtNVKhvHkNCTUXz96jwI4yCejsTm9FbWJoRoVOB2H
hWQhdCRRbPNQsdieX6zYa4mE4EgvO9WxlyXH8w7r7SpSpSD74EcNJU5T6ItmPtumvy4h/shDjdL6
ScsKbDRoylZvBMZNaK1w5kZ/cFdt9C0o1aXBXT/4n3F/eaQEnzMV1yONZin6Gj7huk+gkxC9s6KT
j39v7N4Krjhl74uXrIchJdyizbPcqDftjWDav8IZLVw0M0A6F7WHUPar8FeFKsx89Kqg/8NEVJNQ
dZJ0O6CZ8CATHiV5jrVdQ95dsmRggrv9eDQQmSEyXQRPH1QAvlB4zvYWlTtQGMyCySeUbflJiOZ4
zr0TuGqQgca4TOLOnwU4wDxllLv6qASaoC4q/zW1izecz6gYpPmM7P2wFBTMM1y6Qm7eceMtQsta
he2M6MUIJLMGmnuN2OsW0BHSd9q4vNIDcXqwCf0y+Td1KXGZH56ZPhUYxBZj2a1E+NvoglXv7Pa2
qtbKqEIqIKFkouQYPo4Sc1+9o10jGI3ZWkmNmLRGOMvxxrfteiz9mbA/CjkKcdyx5lzti/TWXD9N
wewwLyEL5xrwaZOOtPGSHssMm/CUzrZ7wYYoDbQsBvfdqj8sU31iyqXQ+msqI8sQ8BzJ7V4GVr7r
q8DFa9aU4wSc70exMggvixKzu80EtXIi562xBVrFXxzfGQhfTxB+exaKW6r1Upae47lQ5bS51wIy
LapbH5zLeTuZRwg9pcdZfGgEuhDvAdPT2ol2kkseHShd8u2zlCZdQajIsk/GfxuwYqvbtvSPBaZa
HyQuWZXyFViQNGqSUlb8SciUY2I09yH4WN0I5L1e5XEKQFKd7hUMWxOffzQD9DKa0pm88qRt5stW
cN/r2CS9/9je+XHLLOdmdgjZvXXJZFxUuYLxk/6kU3VRdn6iBwr5gaSkFWaDtLf+by7o9SrN835F
fGqQNdfIabrf+hf9G/n+p1gJBmzVnKydzHBGvxvghbUCjquqmfPn6af44wuh8JWtXtS5Z4XtulaU
Xfr6YAhUcuI4T1j8rfO5CB3uU3tj7YBVAr/RCKQvhd2nse0JfTad/8EiGpyCAeiofkfm2dPendNi
HsrvEQfP9gaemQ8obC3WFoWYDL0whNY3j1SNQdUwZB7+Sa0ZNiAlmgd1ZSQrRgGykSSK6lAAcWoM
27pLG3vITo6zG/02CNpwPlFHBxpJuRKMQonHi0gAwMX63rk0Uc9/bHmkmJgJdUJ2LSlQvUzkAsC9
zfCkeEu4GwrI+wyI3EiIJ3YD5szqoPfR5dyWJO4QF3MplAn9itz5Mj6TauI1vIL9Mjf54axvl2u0
m5iq3+F8N3zWn/K4lBY4B4p/21+9K63Q50Hg6t/h2Wjcmj7lx1sGYSrlr1Kh99TJQHyEEAkpiyWu
hndqSscKI/jGrF1dphsnpnThboCHHo8DTffjWfWRqRJcS5+KeYxrBdndxCAdDjBgxjgYNCnMkg4w
6oqXCX245nH7dmtTt7ZLhQYFaUmwWS6J3fRVp90e5E+19jFAoJqcLVNOWO9XVjVx57oaptjOnBHY
jefcBbKcam1KbuWUhx9RPnk3a168wMmVwjxLBBcHDmV8LUu5TkZFrfFzB5I7M0GJIX0fUr486kkb
hiRv29bJRfbcLiCa53Bz360u6s2kpwyU5fBAEs6WI0CGX2RDoGVXZwYQKb7GBSj857FkMJuRWo9G
X9aL+IBR93fVBxkKsgIab0Y/uFnX78BdC+Fp0qqBb7UUXAa8CoQJf4S8JhDf1HEjryyaJ5UQLoSm
d4Mwcn74JVHvAj62c6w4pHQhxYZMSyVfsBL7o+8qEWzbasHSorLT9fYa3tDg5tYhjz49WwHrC5ph
2HmZh7QZfV5DHzsJ1WcsVi6oI7oCEJAtW1gPNAoiQ2zNWBjBAIr8lHD6vDOkIAN6kycVh0yDV8tf
Uox6UUkRLUm9nTGkWpTBl97o6iDAF/jh6Qy6wF7h14ulUST4iG7SYatSrDFichd4O1bKQM3Vu88o
9Qv42wG8CkJx/5zppNT0gWKpEaz90YiZ/dRZjlaO0GV3eFFLzOuPwh9BpbYNMZCltgOS5uJuZkyz
5iV3Hq/I7kB8ndU8tu4VWp168GSCHpUGiYqBx4RV4qHBGevn8jtA4TXB8ChaML/vEYFwyUU/BjDS
lNe7DrCWAHdTm+LlEd+tnE0VGsBzMdmHHoUIdIwtEwhj2/vlFfXjr0EiMDRxx9vhfPRrvkHFwPwG
r3zzae1Xh9oYU9lgzpWNNYnYqxG5cUzobjJMA/Nz5+5s9Z2haZE9YtxIT39/ge5024iN+0o38SXT
/Ey+gojzb+w22FUwlvPAdn7nl4eXbt3eKBLIpwoJG9XhfV8FeoLyUAr4upJNxVPnNuIstJImIETT
xhf0Zh0yYCsjjLmtDYovv6rg6tLiQ7z/OZ/rV6ZJv1X0XUqmRShdJBwifXse19Tzl8WYtVBC1tF0
3RUystS/uUej1ueBY+Geaio+PefursZ2r2zTNfT6X7S7+EIyLerxAV9lMLLJeyu+lVxQV9s4mSm6
RTtFf9kmWc8o3FBqvSVZeqbMMR7K4HXmLOevl4iQgnfBzRosprpXD7P2YHWWlH9weeoHWupshTFz
QAhTVOGwhHJr5Yd3ld8YF4P4KwwuZQOuWc74rX8Wm8rgO8Wyi5I3Z/BG0ehsriGMRMHHmKAXOtjw
iNOJyxNUf94tWTTv+NOSs6SpNVbq1nZZzZ+veHuT0Pz3jAPGRN+h9EWhCeuq2hg/0r7cskeul0Hn
N0CVViIxUH68tYjehNgZ26bl8rn6AsupCCaIdkYYgTaPMQ+v+oIohxzG1MwZcVfsGzcS2YiDBVpB
u95ThqvOde4K563AaFHjevjEV3tvfsWLxfZFdkoINJuhDMlCBV53ECMkBfig9i3aBsO5tHkBrU3g
7MPR6di3/fXEGobBHJTnKKxrnU89B6WTuOP5NtAsti9TktG63xOLl/qZDvbkv/GQz7kMKuR8z5rd
8IsCrLIqWmgAnkWCRdzuK/VSevCr9L9/WURK+v2Qmp0xrvcCQUk28L/7uSa0LbP0pXr9eD9CMcdv
e51L6xdYmGlSi62ftnduahNz3mq9dz2fN0iuJuko7A1stx97U9D9qIHiORY2K7idOme5+UudM6Q0
FD8ny0lsKlw0b6uNL2Hoh3ZIUx6EC5TC6+DTAktE6P9e1YBbUqs7WHHlZtxjOvctfkxROvlrR2s2
3NAhvytxANk9nISKPLEXIL2wsnKMexrSRGENDkIkEdwPQOW4D3iM6eXnKKNfklNzNsyTviknVL99
LyNJ+7o5tWa++yboH+X3mLeYfG1/kyeBLzVpqD5m+Af56IVS81vA52PyFTNAnkWN3ZO9YvHbxy2O
0axH2BxU4xZMv0zp4/Kv8I6TgLHU9U7jtEUe5G0nCO5rlluByEXY+bdxXy61hkq/US6+q9bVz4wq
SF03x5yOH5BS8+861bt0FBMXgumzB5s1Uf1HWoqzCZ04Lsd8AZGWzgG/1b6NE6AIV5EJ75+WaHOW
BS7wP2h21UH7O0wTj1y2amhaaDR6VkFARWKOqw6cC+FUdUyfKIw2v1fndUHKwAIZgE2hRq0yFi7f
8Eu882JW8K+b7cERvrkGB9haoFHXLH1T4QuJ3E38aL2ztZuyShDs/fSzTe73qpChrCdG2vju+ag5
5ou9H9S2cb89mAv+tDh1f67nmvR2E0VRvDF8HaiFOnghl0aS4bY/giMwIgm/jwpHZhtWOw7gXbQF
7aPxxIfhtBXsMO+fdEc4aOQ3vXSQSksTRcoUI/jQNzJTUpaEBDyutXmQvF7Ruv3mqOlCC97VLZvL
uP0GG4fLD3IQfS2DAAfEp53pIj1lLd9oDUSQ5bB6/9kpDb4tF3ojz+uLuKwnyi0wOTsdxsQO6zAa
CM0ieQ29Mn35pq1hWpKf+7J08k2yNcvlVAMt1Agmrrtu5KK4jqfhOa501Gx9s9RctaJsbihwaY2q
tLZC+ykdP4Oxkz/LPXh/bCbuPXRST17AUIdPbWOoLBKVnWlMRFDTT40G07nQAuaMQyqOuiEybXRN
WYMQ6FRr95cpDNqxv6q1tg1hSx7swmHp3/R8YZDodoAopFGX4ODrVKqgg687bb/3MxZ5CGON66oG
7D+OziWFnHPebG0Rl6M0jFMx88eSw+LpA8RFnwBrSx3cUtbEjer8M3UNvXA6TWYYBaoUHCjCBp6X
tLJjaUDFzycK9Ny+K/N6ewFsMYD0Y8xSWLtgUD7zHfIiKBbrW3hlHtMLjUuc74En0H5mem7HgT3+
MQ9LR554lKz/x/KSoKnJ0VqMDlfC19CnqryJ8DbCKZbmWFy8cKAsmEtAfXAW6BiBhw2NMvm9wsqg
Jsk42mhY2FTEPghK8tbljqmrqsZzb4yozPqYRpHVIbWMPTa0sf7r8NMwEJVopzeQBPfnzhwwru+5
7AIrVGFDvN2nScjUlF+IQDn+La1YyFjzkjoi6YEbySTgsqoS7XQnXTgM3E3snOr/CXQkz52FHGBc
NcPyCfBPlWNEZ8rCjw4YCMxKsefnmtmnRHSq2XFkuZ1Rj/wuoGLi+EFl2KdkZbeqLKw0JrKT3bQp
HviDEmwYqAlmMeJwxCOygBJIttpzbTHAx8K2qSnhz78meFfv5KgCPc8QxtZtU09wthynkWLoYDbH
7WZiRZfqsRsgGTEpbs4n1EY0p7cr81GRN3FbaTeWpyNJMiDVteFVfDmtaLPTahhDYVDL7enPyJUU
N08ANVcGEcfaa+YHE/QvnCTXkeWRNq57QcIMzLPwqClg2pK3eJgxMMKQawg1G5b6c9xwoFSgPt5D
yTosT/2i1yATCjduSMoURLwEr26Vp0E4G7hCmFHdryeMxLJr1RxELcOKRAAU3ePOBX/JK2KOFDdQ
DreuG5xXkjqkfusWY/XFDdOZi7zm5e/JIYlO/2J+8th1LrYDilEV37x8p+ZXCJtAj4neZFclSLRu
7Sznx77syzfoGPbQzyn5qYOuqRVgwDSexTrxTbafxmwlfWn9eGo75ur0l3MQe8gLpY1F6VE1uWx8
tfHWy8ruZDPpDgBNKDPdt8J1Tn4s5IyW8PUhlmVtE7KRXxb7dZajPrpMoFs2WtO/hHCTWWWsSYa4
Yqp2/csqnPDrssz/lEGAncHITaTxc12K+tx/dnH+IJZsOfNh/xmiYJcciryrhNPPcMDWjs9U2KWS
eBRRFkSNFss4t5V2tDA51t2l+6d7GHCYjA0g+8qharOefohFFNxN4SNVrU+a/xOx34cQkdqGJFLl
nd3fiW/F/U2FwAlVA/eAxPZJMnBMvKCirHwtu+Vac1zSPEiM1cIY+zXAQJ9IlXnryOK3j5cjQbDA
uRZ63eYNJV/hiSPGDSfnmjeVXvgzpAorc8HULOJ9z0P7gE5m5Ptiz3lcdCyn9QXYskEolWYc+7Lb
C+IhxMcEtbY15CjveE9KY05Owci7VcXBjxeWvl0Z+bhF7fBE/tyN6MEifFFOFIqItBMhE+TPLTah
3enqbgHh1Q3ehmT7mENzqhykAIjGelqHnLv18PZdr4Uum2smO8xxeiOhhX3D6YHkJ5dxSt8Alrdn
Y5g6ee6vi7JJpT4r1SaOLhSSYeDTwZwnueJHazjpwTEMZ4oLzAz8BwN41Yyjt379VguhDDT5JHY8
UYQ5ruhLcfxkjJ7t3Qq3dCxoq+KqPxR24+Vb4skWG1WJhX7SW354fyXpzJxDLgZ7OEvInUDY0ea8
lj3OfJLNSM+Dh8oNmY1ulWqoag5Xx2myBYMDqbfnIUmB6yzNUSCMqEdiTo3qxXbCQB9M1M5Az2zE
N39P7Ww2Chtm2MnTiDZfbRDD9gL5SZYdPA83hzmo4I/asoFCMKnrLleazUN+ByEUltSg5KjGxD9d
NY0EwbjUVe3aiWF/lzIqtM7gI4z9gaAOplPJnxbF3Yxzh4h1daAD+3y6wMaDFS+FK04m4zTv/nJw
90nCCNY3JNncCDUZDYKz9UQKaavjOjwv6zfEdYyrzcowLf9CNJ04eiB0z7wZy3WgLlM3D0ANAlPc
aCTg6oqlxzCCaLjxNEzQqlzOeg/L70vNmTtEOM7Zy9lbuUV/6QwwbN2FJYG5OZtoTnvNgHzR3Hxy
2Og6gTnPqfcPrErKXb4Grij7XoMHNszY5ZKK/I1qCbViFCit4wXLtSLm/1Ulh2ddImUKRolyJGZJ
tESglJLMmQYSa9sen+9zflIUxRBYN3gTvv5KFJpKmGWGkC7k1TcQMvtUri0daMK3gggBovg2IRjK
daGwLAPL5lTg/KQ49yzzJHTGb437ErQR8FsdL82bHubA4N7UIQFPHYrGwGvVqTTnNai9BHybq4J2
j0OPZp3g3OCfGeTlljIQXc69Sjaw7nHKEOKcXwPeG1HedsRFhe/xAjlWRxSbTb6/ZGX4/j5jevyq
mIFik190sBjoWq4BG52Lby0RslTYg/F7BvMrMYZ/RaTJgK8wAs7DxgaHJth+y4KkoZ3ktZDn/ssy
ITCxijZqfAgfXKoAa8DRUetBrIaj6NHTnPN3eUMTh1V3N/U9hhx4yqmaABJLSeksYcQ4h9zLq9SN
0AMvu0ACQBnmRbgmWtr/OXJHTIrcCT+gansOZK56SDZJ/ro+ABTbDrMgnCMfJ4m8oK97/iXJbJXR
SDidnN2N7dpGOeaXLosBpN0A12t9kdvtm1EgbuicvFi//1Ma7PjWh72xPb8RtB/WK3F77EmiUv6G
gpZgVKP0p0TJRj4k/9zcRRLu+EA4xqkwNP/U3w809J9c19gU/0ddv6zzw3VCcqHBrNd3CFixjmDV
0dZtYpZ2W/DPNQxr6I86NaclJhER6mUPj7rKFqZXY5rA4ehfeYVlh+KWCn3ttTHNI2RZQZ6vxpwJ
so9Z6E7ATIYoziSvxrITJkAXKBmVQNrmYiijZsJYLMRH454IZqI971YXJh+q1CanWWH1CsfMSpVa
WShCGcMALBGKrZKAPtw4LYKMGRjny9Z//P5SLDLZ5zoR8uo9ReDw+kcaxd4b3UI7npE+h0GF68nS
XDY2T09gCtPzvHvjnHlRNn7TTCJNMMmLU/nmdekZjE+eIcY1oN6xbRZJ2ygDw5o6ll1FTzsmYR6S
1jCcS4MpN8X1ORbVsem8t8rVdQfvhdnGjzv0XtwcxAyfuFK9fBYRVJvHf+geMuAVxwFZifHWCBYE
Wtoie7ntg/3xgozO0Hdi2hFOyBELDqovf6bNbPCEk4YW9Z/GI6FFhIcZkAH29BnuUg4+qrHSxA8o
nL02TJaMkH5RdQ0V3rnd2kfvqE7b3SXrl5X3pWN6/1wp+SzxyYgi2DzQrEBPiYiep2dhqjzX5xjl
CKfSs0MlfapIb9TDcehGakZeHJ1m0TsdH7lvGu1FdZ5mac6M2QWCjGwn7ep99B4m/BxwA3N1RowD
trFwIVwhp6Cr60PkrexZel42QmENNXSlpWFXfbrqJxZzEARAkVLTkFf9ysDwMKJAKucx0jgrKeFt
/sgnwC/GALjv2IAVh33wfrWR9msA0ON0utjM+nEeRD2kWX4devPhY7gVXf3F7ZlMI8B3wPEpqMj6
CZVJdaq70OuiWUq38l4qxgnbNU8SHz0dkJru5l7D6kD2Kq684qOAHPp2kDxaTOuuZR9a++rfH3fF
hGaPsbfnK1Ggt3zADAMfyVN9xTrUqCXJRece8xdmNMXsKK0TjLruKdxumSFKrJb2bgkvdYjz9+rj
NxmzLQiMSa9Mz2ZGCkDigKj2n1lbENN7x4Gb/h1m4PnvKzPcoVJZBVz/gaCt1fl56wqNTUGpzme5
Ef39fypC8HUKpeW7kcJzqJY1pLedgCSH0IWyOaSuFqbU/6REwCC6qyGsLVhZ7mkYuiz1+d3MzEEh
Hflbc56g3bwBvLwJdk/fjVnslyE6PgQxA/TYY6b2VP13TkI0mOUXS9LQwx/yW7i9AryyGPE1yBFV
dXmXz45TiBN2i2waU85aDMkDefNJaP5hoCqNLOaKEcfDVh6IXgT911Z0rV62lMqcLywWI2lfQB9n
sIY0lQtFmuigsIwvrSi8dPacpf+YUbN2Byf+tGQDT5LC7+7CHQwA5BKXXICCCnoWAUal2PX3sTap
oc6vf0iBjiIrTq+uhUyBucSx7ItK8ePA2sW18TF5q+n204FHNVjVpMpfrtQxoi2rxGmZLHfwbZ0X
YHOzatjXNLX4EhuT1GJ+8x8NVZcopztUNHOMQHEEkPlE4HBtI5I8hrrHKArF4uXontAmTeOLAUDg
8aaDiR68K5kGaH1LhdIY4STivWTV0a88Q6MX3bbwGgLjvmb59JcP76GGclxh2nkBj789qzxw33tK
ty3Xo/7CNhP56zntKs95M8wB0+JCEAhmeU03UYiqYBJHhbpIC/JrirFEHMDjxu9y3id4p9EYG+j6
NUx2NdLgG8YLsDfNpUV3USLyZa4McY24d8VnI04gr3jdnamvpKmaCp1/LJUZzqPUH4cHOz450vpZ
jIb02PtjRUTo7TBRl0Vk9HNTOxiQd9n6ysp46L/NkNFhOL94jgfD2Zs6hd7raTq58X4/FUgGKf7Y
YB7s5KtudhuuIJjpXmdhDcFX0zKEo2vdIHl9ht/lcPV+8MAd8XPKO4ndQpqEc1h70/6zjsIBaBR+
qTh8pqsvc4snjilImMxww6EcRLMy+CKKXEMtlHx5mv5k7fmSvwOn6G5IyiDJ0GESQSIe0N268eah
5+5+QX4FwOxXaomwvHKsMAfT6HvBj+mmNaWtnjjBj2Vc0ZDgDFyme+N1fA6I6ZusvFXNjzN3Ob6z
MyKaYnlrp+GEVPHuByGgPEZ9ci83szpPtX2n5ciHPsIdWqM8/wNW6/xzFKXz3io53n/iFI6UF3/K
RSJZVOmqre4vmKK/89GXLn9gVRKL/SUp2wvFyu67Cd/TfO4Mhc8W7KP9PX77eMXS50K/V14+NkfN
ifjIAf7vBehwvPygf1qlqZAjMwlwud2Jjsevw3EleLOLc/FSIvvE4UGXeGEh0eDEutWtET9tuEfz
wo6olyPng8yed3F06u36EOnjYo2IX4QlMIHeWv9+WJet9i5ny9/5iRjfsjJmLdwE4k5rM4ZoG8cQ
m5zjvEKLhiFOY+P32gGZzncJfZbItnc8xYgA9lU/PpQkw9ox9h4ai//OaG0tXhxmMcLS6l+3FNX3
Jv8vPgGEXT5zTlPpSfSriNzVXDI8x26IWCs3mAV3V3UclVgSMB2PLiXxMQ7dshLWZsgcKsRGjY1y
rRTBMgRuhuJskM2Ux2SZ4ym5oGtvfDnxjbilwAOQZET92pv0RRjRa1uawUpm+5TKXonYipcjzt+N
Vr+q+dA7XAnRU5PzThps5XcbLlT2GPCpOXAJEvAbJETPvgt7/dTjRCxKrT2vcoz4/TlSO1jSPPEj
cZKKVTAslWZskawccNMJ6dkuwi/+ynbBNhb2JH6Eap/zo61KWY9+kV/I1xHFRBbMu3gTj6eE9BZR
n9/TN3HA5fDHUWsaQuIQrOmh7R1P3xW9EPL+glqlrVWIH+GgvFky8SmzrpWF24kaqRyHRt50X5UU
EWg8UyrAjcn+9FNy/dDLG4obETSP7hi2XGY8M/xr64R/K0g2v/ngkImMTKI4G28lbPMrlaj0Euiy
sEuVfwwBaddHSD88F7/qAjgrDMN6IC2uu5vweBEYku4usGKcrO3+cq0q/DlbTl+RZ5FaUpI7O2gw
+XGdOUmKuM1Y6cSxnA7c9C4Mu78WQS5Tk3HfnGnjETMJONOvcIdCyqUFUnfqgRdAjpDlRcLTTn3x
Smgn4XCYoX57j6fbBc57OU52LFUH+nvzQKeycB6UbQibU5KaWvydg9gYZo1ansblztHKv2PEgWVi
eXvHsA6Is7TW2gEyiWMt+Y/9sGdFM412zda6wHYa/RrtyoZUsox/Jj9f6SpcX11eCj99HN8xB0vS
ln2A9VGs64YNYw6SI/GK7sXk0cpIu1hDla7vHFwaYUDDm5FsJ4lbh4Oa7uhOHf6EWqoB91GZ35EP
hzJI/bQyhqgG0x08jiOvzDmj0PnD337Dbvd7dxg7se1EGHTjSiwEW731KlNvI6HRI2bl09IeZkyN
QABdAFG/iHjRHmugi6D1BYJW6Tqz33aQSz2vA74R20LRKvngmH4Q1adE+9Ug6bAsoy0/1hJj9rpK
+AkNKNggBkq71wjD816c3G2cbOtGAVp2pDN9thPH3ttG4pr6HzubuZSg9NjQzESNtYg8Sh0o4+bJ
kfdfzednCY10jc6tFEA1Z7QckOeS3nqKaSXD3Han7IJr8TS12NLDAvQBQB+fklXyJM2F8y5iAIF7
c6Vh4pnlvJEz8av+lPHUsVf+2b8nnPpj1SZdZBbQnIfuB60Jq+Vqg5NppV+fkNfz127895JZ45+p
eWCW92nYU2Wsl8XUtIIrNcSExk5uiaWCW2c5cIfT21YE6FhpTVqB43VMuVJXcqwJE/2YuD2RueB1
B/nvNhTWEyW+Hnkh+nEdXY60YaJTEWvwJQ8NIM9PLmFbHXjzPgQBpRBRNlGDUyDDfq0fUvVWSsjr
g+aZ9et7pZBFz0w62cqqwft+H/CIXtwZ1es1te9WRH5Ai2r7XC9KRXPPFRqLeM7/Pdf763d6BJgb
IlBGAfyzyVjiSwy1W7IDvlf61qXaiZt51C7L8wwfKyiACqAQZ/7v5E+EhbXbKxkoRX8gn3Q0+PUw
y+NEnus78xuAvO+iJV/C0GSZwHlMAKmVyYPHQmeUxhS94gpsejBbU6FpQV2if4e9ZUncysBBx65o
adQHpFQFYpTqxI9x9AuGF8/tw/ckmiGaBItuFBDCKN2H6fD4iHcjtiCh3KW/BnurRsx0Ykt3zgwm
tEu6Ujo6v2pgVNMDk6QAROuTjqKEv55l+MnLVhUShP0ZMLLBJo3jDTnC4zFpzic90xkgltswyRBJ
oU1uVK7iAQ+sTNbm2hGav3vSzQR9WnOFX+sV46v30EtpuamS3KmgtmX7o1AL/iYHoH9JIxZlJrPg
4wT3Snivdvi+BzHUN6ianAH7jyTQmigdHIUgASCpNZqiHSLC3ZeeBVKHm37NkMsp44i1Y1ICidj6
Gwc0J4k+iVyH5QQwKtauzbVc3bKOrkUzWaz+7rPW0R1EkCdqDhoXys5ibop58Kz58L7AymLOC/vO
6o9lN23tDkg3SJDEeg6Lb9bqJ78MiT0Fo8SvkJ9qvsqEmusRHn+uQl2YbRUrdG03Rmboy1J6/6oe
/M/4dGy5NE+43Fnnt6pgjomoezRWqFkRXX4sowJq6rCF6U0ANaPb4zbO+XV3UsQeR7rTD3vXO1YS
BPlYwZgxQDZ+p/pKIWE/DyswTCsAIndvnWvbqbTtiAfZP3jQFXfJJXlph8OQ9O4P8IThYX9i3d+z
n22YP2Oc35s2kHImp6JcHMihBk2rJnsiduNaNavXkMLGjDs3btziiujDNqVi9qg6hBL3N0807X8K
V8zfcyqBC73a4aWGfmU/oFn45sZfBw8q7syOuR2DJhVvomxQ+crSMRxfJAJvWTvxTJAO1P7GJe9l
og0+Gy98NAE+c5ExO8MRPcYwDpFwSlHx1abUvQdFT1gnJa2Cs4qiQY3FQyB83WacNhys2kYzwISz
vdAF2Bab6VInrRrbkyQg/5Q+bveNB3ANWZR9wppsmpg2dA6vztIEg0CR2b7qlkA3afsVjVgyPpWF
7YYz+7jD8iJCWJYAUdjlKOzNOQa8WIDF9pT9FeHzJqZWnBu0VSAxyHBufj0HGfdz+8UcmduRwoFB
o5JvjSDfDVfNRk3hwIM3niRVKrcfo/lO3wvf4iEbQGGZRutFkijunlx+uuc3nZG/EWB4JkW/UFHs
oUhNBRMYDd9+yq24gQHxmnuZlaci6jGRUtAaO9OLfaT6eU2g/SNNnC5QBDe5LChUZDP2ph8xcC2a
dVaq0UPsW80Cm0Nao/oWbVymiCuFTkYpRcQMKkQIK+wNsmivPNvANqzMSUEofvP78/V9llSc190j
+nScS412N/eM/4D02Rg26a9Kw9h1c+F4qMQrVkd26NyXQt/2tGTyL0LQ3p3PguMvOJjpTzPFegL0
XVINfLUYaHixbl7f2JvKlnoAUtp2ntje1snCtmrp1rgYNRiNZpocLb3s5xhwT0D92rgBGLfR3Vhk
s1hbzBndOmjVGUrtuBXdD5IPCgkDRjoJTFTvtlpvThd9P7riH1DX1Mhu+B97UhHOLOocv3m9GtYI
k0kvhznqbmf9nUkTQE61A5sxXn6aoLCTzKjEr30gcvWOw5rKDqS6GQfuUqA79xOGqOe1qXWkKvu4
VpfroWWDA3qO7uRqIntucwR4xzFr9Y3FfletSQdnOY+Dy2rlbjM1Xyy1tly+jDkMAaE2nZfQZDCo
2xyvnBPYrBzFKoq2aHurJmikGUvnsw3wY4Se8Dxu90ZJa6xlHS4rE5vxlo8NUi2C906sDA1Kj+Dv
PoqCP8C4NQ0eZf6TnyYh1PMRXNTkZ/AFI/a3RMggWwrTQrjcf8LnnQRHeyYD/EdcDbmNwrNFFl37
yTrWLCMvtK1XH/v6Zsc6/aYz27gvb1q862lgY9ADq5TghSQHsb4j9xDDzSmBc5TFXrTC8XKKhCmu
Xf+Zo96W35tTHx5d5Uoo+f7moXryOz6RJ4sHJAqiY/yH7YII1PfTnaQCzjJ+n6dBSCCtzT9uwsAQ
ps2nYnfIr+G4eDf/VddgNcRnZDGGAGqeFEl8SYZtLV4pmbOm9D4We+rZowNy9gYfH1HOCIYF4pzF
MhuKKj7EzUbl8Rbj1mvlBMT+Yjdj7W3PkHgAmRbve29+wVKPsehXN5TRQxUIreRxz1bZjvtEfeYt
t5zXd+bKhV/Ze9UVPzDJ2b5yJHhNT5y7ReA6w7NA2uurPuAH5mOIbKgpwowcg8T/FkSTEVGuJJa4
+fABCTGtHs3gjK0SRAyMEGsg/BwdPiRQ9EwDKqapTt075ExqDY7BTU96TmrNbnMOWRfBsTS+do9G
9YXnEVqmId7ozCv6pA6L6COzI50HZsWKzsOrtsD2f4KAGCcQpJXbYa+/V79Ms1OX1EQ7B8IChbuW
WmdI1nUS4n77DABiE91cu7zoZdQ5BudwqJ+4jL/z6ny5bbLiYpB+Fq/u4RTXsCZmSeaSLNr28dUR
r99eYTWqB8JdKLuboVApAalCEebNYxxwPBZv9R4xFKv/pkp8GxINRS+4cgANNfGUhCv1dGx/9uv3
oKJu+KHXLAMbnCTZiYLG0+nGdmGaT8E3F/th4k5X3HsDVjdIjdqIy48UduZwKasaIEBvgOWGAtO8
hCyZ0r/rT/RlggjY7iIASw64UwTe0zhbhDNQEKsf/UFLxaeBkPPIwGfRQpTAwJ4j+ByV0mCVWDBF
vxAtCtD+DITY5U5mXeiBW/MOcrh+HAVl4sbVdKmMP7ZRAHC3w4WrdBA1xq3LPn0XpWIOLFfC1wZT
k0BtJehTdwL47HmtZ1+/UcT9KALMBHlbTBvBDYaS85WmSGf/VZYqoCPA22uUMbpmDMUdh5swja8H
xpLU/on7j6YAD60bmqW3heVh21yCqRJYdsyzioMID5XrUBNbYCy8MvNeyUX80nBlneAQzMS34b2q
jrXJHNrlO5j+G5AabpnSxc2JmIiG+gcgztNauh6AUr7OERBhV2RU+0fdZKe9faiNz02+A+ltIMIi
+7aOPiyhwp59T37kUmAHyeIfutlLHY1T/Mgs1LCjeeY3OnCZSGn4Fg1ArQNLasF9fNjrXQWg+J7L
bU8c5AresZjP1nJxywnpP10b2wNXoN916B1PoM65XwW+jSuEf9Fhhp5imxKzNy9fqXvXd2YZ0uFk
T4D67Ld1buVNfnCFE/FXcgOi2uob4go5klb3J8N5u2jmaMu/osENawmlDSqsbvzURxDDA8QegQmZ
+TXfPVMdRj2N3lmBJmaJY3w5yaTeyu2YrxWYG03xoGbtL+SKcRcXOzJf9wHXcXXaQSh9qOO9ReqQ
+uG42qKcyxTZvG+q7bBzCmht2YW4gDsLaGpEcK7e0LUS9FlxXGbvoNl3tl8uPWrMX3M7n/aE6B7E
JT+EWx6BJNDjyaZB5rOxw1i9pBWEsJ9ywKfc4MOi2JBn1t4qRtzyL3ijLqbMTwK43lN1Ok9HZvtV
EzxQaoB4MsVna1bb7Ccb8s57BPhmnT4kqUebW7OhCrm+6MdD58yM/YOj+DGeVRUSnyrW7MKifup8
mKDFCyiKFB7v+eSwKDaOzeSGTk04ybjvBaVdEg4Oa5vgT1NXP8+8xR43Bc9Pt0+nlTMLJPlRfknz
qcmpptDOoKPSOWhgmkG9L/omUjz+oWYHx18P2XCy0l4DrivxlcWQ5+otbXKG4Nrh9tdZh/XM0Tf2
k2OQCJRSPXXwv/dLC+q+e3gki2aWzt6OAxyPK4KG3JpaN7fXlLzWNX6cT48myVRC4QlusXgzXceZ
XfGraxjJuqdGLD2pAgxYW13eulkZCNAu001MYUZcSkoRB/rhUiTiC38YD0wtVAfYf6SpUBISobwO
RKlXZNWwR4ZMx8IfBL3hvTUYBnl5qMLrCqUxWeBr7YdHw8yPPAXXdx2g2VqtOB5p0EYOJoitxVAz
dnQkf4lFd6A2LXh1DgVMRVHLCi7GDKvy7Yf3hWOe5HzbyqgcY0F2OkETRJLh54RH9xEyUzYw7boo
oUtXrhyJn43O0k2l2v5EY4IQ6h2Q7Lclbro6UGswS0+R3CEMLGoF7et4Kw6O/jlI2cjo/UFSQlKK
8QiLjVMT+CaaDset6zi54VqOKDjY6HXHRMFAqvqSJ6bs3yG6IaRR9Q61D8Smm1DxXllykBzRv1Ag
JeoJXPI1PzitY5DPrNT8hCjt1jr/HKsFMTuV6tRJx7La2RtrWP2GssVlLphKfdihul1xGiv99eDI
GDZZ6OQhQTxVT1iUJlYh3+zgXK1S9TO+cqqAy1L+tg57Bh7bmVh7WNJUeONvUW0rywTP8T/SIJmu
5J7uRm2XSy7wRsR4joA7adnw7t9yum5NGcKYcZZwggXZ8NNJqIv4RXQgBDRoaFsjSL3jM4mlyqRz
1yIcnn2nlJc0i8DNjTWpOcRGQ8Wy2jvgYQVtHfebDz0i1E88XvqO/26PttbVphAf2+gegyHcHvRv
ZwPKtrKeGcuVDnMt6LkW1GmR52u75VbJaHeC687WVAIw6Z7hum4mIEqkilI0nuDT12MPd3UGtfxY
+XhCv62iz8OIow7khqGIXbU5+XWgznbd3ldJ+G4BKvIoAZvzhHyfjcczIbT4t/ArimnN4zk4rw41
2NtU1kkq5T9W9orgVu7QMBkUl6m5xDCFUwoXKjFe96IHCMowAgOJgprFMPlqRp3//B4x2RDBX50r
j5COMfjYLCcA+bDluuvLyaryQFCd6PLScrMq9l7cD7FkVJokZ1/qUmuvy9DdEYZdwbuq+n3kjjpd
A1OipVc9crFCqOyg8pUCHyk5j2nhDb+YvhHM2X1m9vIdB+nN1m/mC+xruJh2re5gAOw1FA/1C5nl
wVB+h1MVZOAGID86Hd5m15JWkVYI/YLOYR5dghHCdj83gPoDy2Abc/8LmsWEs31dOI3XxssWIWaH
oPJB4EU5F1qMwwPIHGJy//Pv/pmM69oF9fBjJxgAGUF0o06ghYQ+vGUHsymM2PAoIfA5iEf4iuXM
NUc+MXKztTrXM3dMJZ+LBWuRDkSH3ibbU9ocriti76+x5cBlv7gIXAHbvWtxd8QheFRsQO/NKVbx
s8GnXa4zN9ChR/0CejqjA3lwdVr3bsMXP5HJBwQETSbF8hsmCiF7PPcGyYlw+HuDCyfUYV8m5bHJ
Kd0gFkpe6o83y5saITSpO6gpFvadvUlBolk6Y6rToX9r7H3x6qWeiWy0vQ/8f9khW2i6MCukWSj+
LK3A4Q/1uzFQJFnxdcIYn+FWCGhFmX4iVtIp6NuSUegYOE0fh+5+Hm1FuKCaVr/bP6rX8QgdDCcT
r7uc6f5wDhbVJuOooeFo13jhfJMwFb3pY0vkAn9ObktmCOfpKZJC3pVwoizvuPQEGvErQ1uM7gzC
h5tfXZlA0qgsqAkFiiiXWVB49eSaXLo0WAEqC4F4uznO3mXf1rsEbhsLco9gPvaJW5REYrQ0OGhd
eZr0Vfwek4dJa4eHDWxrw6Pw67mmKzfXq/1UTdZKt3M3e4rVeB8qTTgkcl3Drq0azlbvISnpIJbZ
sygvQK+upZ9t4a4DURy8HgSAmSrDNDC7Wy2uP2oEAt9e1ZqKuiROBJig8HUrQ7DEyR16L0S1Pnhk
ze9NgxrbjFXRfGMJL9238M1J3DfyeciujcwXIyAd2V8sTeEIiGz/awEKVFmJy9Yw2R6ptjwNyD38
iAU7JVbjsE7LKllvUDz6TPBoeFKfuBd7PIKMVi3tRF57JmVYOHW/KfN+BpV430/jE2hM+GHNpirL
aRMMy/qXUSHDXXgq0OprCb0ty5DW7zQToQaRxwM2fjj/H8PoJwclEqadG1zvNUi0rHsl82yKKDr8
wcrMFSxEiy+cO2GvI5kBC9k9axfg9wrr14CoPT+87BlyYEbuaJQmn5vTiGmz/5CPoGMIlCCLeFn8
lqkGtN6I0YlG3GWfYfowE+LD8gq/1gxnSqRuzZpp02y07WLkbOZjWM4DndZTJDyk67V3OYaKZyvT
1XwQ59fcYx1bBKjrY/x5u8834JS97LB9WI9+SbSLf3yLVV0/XXCWSGXqI8JfZOzmU4gvQEaBxdby
zXcJW07stb1Jehhd3kMF35uDrlm61tn12fxrLN89QsHhSjM3jl1KRXOunCyN6MdkDQc1ZbYz/3/E
TPWZrXeegxZJxVS3Pawd8QfwP4gILlplGBFmPQcxbSgoJ3YHUvnGV6RbjY/7DvKcxDR+SSdwaZbI
xEOLS9BjQrKpJ6NJgTLXWLGiq3OoVYrXsTLls9n1RiAUssIu6G/UDZZRc900u/2HM2IA9NfPZTFi
l6m1a/BnEVedStSP5SjsxGS4lEWxVdyH67Qu6wbt2/qeW+HqgFKaiRBYrBX8gluzxELqoeD1VQvF
vPUUlr1Fsk6SjnclbaVdpprue785FzaaAh0FVnpYceaog46FR9GQrquCcUtRraFNHXc1YAN3aQQY
9hZ+3yzjW5iHIt/VP0Tdz9OvAJYu4FMOZFy3t/TcR+LnPcfnjnkPxUJrmPIvQz1RxSWZquBeNvIV
FaZW0vVR+mp8EH7NfcBTkeDfr3t9xEsxK7Yvy+vm2fnrgSZxRZmqj6c1eQXLBtS8wYDJ2TJJGHIz
EvJFNCQy7yxOhsdvVnxk+G3TSUoLzHAUXA2Heiesgr4EYsfrfzAh1VpqJuqfyyznKy2WJlwdGYX6
IGt5TNHq7MUWtFAvDTvSQc8AXaqxEW2BcZI5wPwxn5PVoPb+Ke6V+QMrrC9NTJpq6N7W9XU+0Yf8
277uN45SNv10BLSlXWJvWgdKltya0QV0HFOKaWwBtC5mJa996r8ZZo78ZBPIE1jmSA/MwII9MBVK
HyDHFA8m29IwWp9UAE8rsWFQfGabrBI7fJ/UA8Jq6tUO4K+CZmghdFzRTi5V5ElquuPZ3y/NP9SX
YCD/n5nsO3hmSkmHhRA5pfmEtUzCAe8vRtejIQriZtL7jKjrtzIHmxMAJ9NuNnq2EjNtYtizEqoa
0LBRJqGMv6AInBjV9MID3bOHh6jAJbLn9Cr4fLWskbnf4Tlv1rJFrmuZu7csEvyxaxA/Yr73Nlgd
yDTlvqI/Jc0gv6nxgctOH1I9LsDeKP9kLW30/fLbP4Ik8olk4dl0uluYRI/3f5xM96j1aen3mxne
6oBI48tlheA2WlTHHb0h/+HYiUwxee4dHM96TFMdtTb/9koZaNaoWJC/0VrA/P5mUb1EBTqvaSxj
qxCSmykYhwcKrPhNitLPujdg5zUYuMoRdQ+mLLSoFMOpPvYTW4ORzemYd9VrpiZru1/NxcRUIlvO
7qBjWvozpdzckw75Xz6wJivd5FhHp89pa/AqVjSxgKc+OTFnIYm6f/i1w8BbAXCTn8sR6ipYUTfm
j+jHVP2D4cQrTS6c3B71adnws47T7xHPfAY7Iv745Mo5uXXwrRxLylVI7VOWaenw0yJ/6/F+lHY3
RN47WSSYLPIoDier0bPHTyPtifYY+umXBmp8RKz4HqK4E2u9CfnoiviecmXsE1pObXxUKvN6rjCv
+4inQ35efILuACKmD9vo/ZTHXQAjkXJxoV7s2tvF3gqc4Ps7W7PkR8zVa3Fly1B005Ahq0EK/vjz
pI+4/NXhHB8G/lGlayse9aZMe4GxR19UYRIi7eD/DoEl6M1IaLRF8HWL3US8IX29DKddlu64NZEV
lBq0SXN/9LAW31axF5CxA9DzQGIDpQ2gMvRZxCPZ7LGOwULyBFrXvisHuwQ8Ufq9T1rD9RUpvQAQ
5s0jF5KI/4kZN5TJmEJos95FKSEl4tO40Enupnwt6yWNTjzrm3/nZc2csMW96NJJron+W3cpn6Yc
2ksO4PaJUUgQIKMCuaThNfeBW3SbLPq6m4SwBbPQW7UZI4/0vc1MfCov7XrqeAgy51fXzKssH8kZ
vwJPk8uhGwq56/E/BIDQajMljevXpsjJvpJwgv9TtaLWlWw1PJpoqp3D2R3pmrPMz81rCQVQLO3r
E5+/+BGtEGhGPEu7DnP7JFVbQKX11JrEPvy/iYDjw/xbMo95A3MAJdIYgGGBlZJ5YWPwCfd83FuJ
VivNTfs4HGeesWJGnDyVTNWJBhixu2MZB7DPYHUbacCmuQceDqVub8uyQ2t+ODR96nwWsMICkn3m
PGapzu9zjmo+OSqso7+w/Ph2tR9lsZHpbRgr/yBo7b7E9VNIiU6pgMUFtXQcMRXEt10AeOD/5cBI
A5c7C3co3YGcwz7FKjSm4JPwDzDur33fQZ27/ARoKXzfX6BgSHXY3uiuhgqLp6QYBxU1YQjZ7CeN
lAvjtNmlDDcYNQpIulbem3bcJ6FB3ehpozt/HKysifcOUtckL+33gTez3zB9xXV/ip9ThMjKKoLA
yYve71gJOQaXN7z4MfUAUuPrmVySGWyeNNPSQPOHgh+/rF9HXKOPx+fzep0ODGXQX+ePdyxzJWu3
VrlaOvC3fIfoJFJ9xnIft+ziL0puga3vu65wM9+enOA4wN+7MoUkvF7ZbCVWS9Iq7J8SB0wcrxCi
xCtuDhr6stqZTAGGvbA3UzFcy22KEU+N/hS6AkRLzcsOqdyBo2TsKWp2kcC2v1WJOO304k/m+Faj
Wz8jGCrhoSEWsRWKmwaVsbHQmy+T2itqdPmKMp7lUSL8A53vNMQTPB7Ghjsfjn4VeVvHVaZu2oih
GFnr/5thaUvoHbTvgqYDRnizPQU8F7X4M4Eea/kIExoKlORpnJeSvD5e6IqOTZjR9BanjjScxQCm
dWXBxui3PTzv+Bo7xoYkvMGEGiPPTo9XhWUSSafjlcNbpnxkwg0Qbp7XChAuiUtzWXYVkvCcN5oW
I9KtbfQ8o83XzFK1DqGkYK2DZGhB+U7AdqlnMrry4k8MX6ZOxNq77bkunq9ONtHnjPdOb4h3P51j
TyjTrYz33qKoGmx4g/uvCUK575iNX65UhZEItsqHh5DZppcNIRtyu4cwImN5ytEGQ0aknWzfg+Iv
h6YxKAT0LUDaIWCk/P9niOsBhwW4aeqJvIOVv58n0tT5sO2L9O7qhFZgD04izlL6WP7A5AxOaX6N
9Bhyt68oy2w2f8qCAA/zz2ZjLup8TIHKzdDMu9/rVtvWLFruoncrs7NTkELQvOnZNw55wx8ThS0n
AEqf7o6Bvr4C9B6LRJt4l51RZKPtOirKXRylTe2WefxI8dDRJyvlrLrWvV9gzD8v5U5esTfdLGL8
LQdO8VN6wBjd78TvJTwpXRMOTRXmjUcO5mSpyby6uGUmo2C/sVGUxLjmbDG5LaHea1nvegtydtQc
HfvOoSTAZGRiHg7b2f8sBRL9M+AqZcwQAtzUSQktUDOGis+aFeRMeUK3SAOg5hqvqzDom2ooRZIp
+1hL+SSxBEiSi7AOPLBIZR8YjCAmSBMnMG9M7+ZL8MDGlATKFEpYxK+RWfR60kZKKo1yHbrkncYX
rOuAMte5zNNukJk5my+lrjLZB+Qo2YsC35IZ81RU9Yrp1f6JlU4tTBGyFcWJisgvMHJkehw+lE4f
6n+ABd00YGK1r9ofaQNGRpdpsceYyzhWM3Y9DOR0PRJ3ZopKd/V7EknVUbhP4Bolt8/yac5surpZ
LvrIjvYWipJtG6a6G016aZZnpyJoJjBlGPWRFn1HnOLLIWz1aWTvI856peCfJw8RvUDkAiH/Z2V5
IReLMTHW48sRYWMItk0HZ4jK0R0WCEceXU/Ik59cWcdT7vkUc0dNRQoAq+3uUE5/EYwN8TYztYow
Te0NHL9DPHK3BvLzxUWeGbPxtHOdytMJ9+NxEDqCjlf3KKV7M5bsdlYkq5Yj1b0r2S+QNtDCRBMx
9J+b8zpkrII0xw8/mP+yiS7Wu7yhdrq90C93MR+u+serv+gXl6hMDSSJT91bAoWPmh5XT9xE6XuB
WuujsTO/XVq+O/Wb3rtW408qhbcwroGGv5G7f53752dmTogUV6IVBWjXABdqSMrMJ8W2TMMWFvoe
yDx4GR9WN433b1BZn78labss+MFPa9os1NsFsTWLejrOOMrrKHX0ux6bKcbQnQCFuP6turttKbPM
9audR33xq1Bm12bFVFoXvFkPvnW8j8YWre0v2ZN1PwJmoSCrxGZkaHgR281ynCirfmjvd6d9O6eK
o3Bpo+zVQ5EANEH2zb9R29ZlPMVg7BiIaGClNAXUHE06QVtAgi84ICxCZ9ulrSsFp28ISkd3sp3v
XwPJ41CLdpxlmO0s42LQc5FoUV/ORZDYXkIXra9kRZ6agZ+kpBo+Kw+AGO8C6e13NoogWcdkwf+b
U8MDaPQ19sLAfNZcWeMB7+sWgC/mnq/pWq6tEM6SvOV1k5hEXk4x5g9aGg+wbvmHjh8OxrIgdmnK
U7w8F+w3OGjejiW1k/2JPSc8DvJs2j3qbP9QA/h1biN1beLefl1RivrVObCOUzFGznd4fUDJIMu0
zfopnkfPQcyQyGDG1U6pGsdo6Nyu7D6IfBxxhHkqKrJkje6F9AqW6JLNQ9EUHb16j0sGsqJ3Vw5p
3TwtkcJBdS+FFTq4vWBk1vHAYxMsupIjO/K+TpemzA3waJZDXVb4jMef572MCoFV3DFX/6n4cA+l
fGxvFp9IAhmXvK8Y6jVuJCRFBKdlSPPYSK0GuaUGMoRLUH/5EFMB3fneO9GBfzIsiP0ixdUtstYj
k7PEwfvPXmqqXLyZ6r+q/GQnwz79E0x5huNloPDTDCAU6wy6ai2AZtHLql35pxXx7T+wGyF4H48l
vDK9LLXgdzaYanVi/m1qowK8ZZHiA+ZsBbLvvRtNZYCJ5HRKxVXDAZmzN6B1cpk0JB30vtqRHXyA
YQ8+6ssMUIUOY19sTQY42Vh7UD+yPGJHS/TSMQp45zy3R6BOVCnoETcYpHTL2olrGMCed7xa6OCO
O/SbPMq3DyaQRwKh1u5OqIo22814ShbIHesd98psF0jFeEWJOuUCxlMsk6pUFoLC6ApG4/bDxZUi
QKhTGTigbjVyo4WlzhUoSnQ1Gjn1jmw39HoC4rt03LCLK1qhKBXk2pIlKuJKC7JC78JJumHm4tG4
SB0Az2T1WKEK9ksy8BRwgkNYIJmSjs5UhN30B0B/w3Y3+99zK+srk+P11lRrsh4mIIDMIYZfzTX3
73IANVI8eHZbbMFxdynthmA6fjTB5Pr8TQpV8fCO7DiYuqMciywC6Yk2XRvRmYyl3PS4IEFd+jBb
Z4vg6WVUHbiLKUbzJAPsDTSz6IC2Ak8BlS3cMNOmW+k1GHaKVzakQb2ovWbOUN6p1FpnS7zfJvgW
9gxgHNiN+EgDmzaZLhpaSb8EalFkaeykzZXA5VQAkuymWz/owy/r78WSeNtQCvHiGqvcMdWucRPE
oIuVujRSakM9Sr0bF6PY19jkYyQhVmaxieGYyICJJcYC0ZcqyO7HPpim73aN6B3AzlkqDHfXAZQg
enMwDNftYS20fg73JAF29XiWi7FEqVH+1UGqPr+/pmHBzuWswYqTlKpjN/GbBOGRpoKajJUmuisA
mCx9SjQOmIROPbvs8QHWWDxGyatqPSGviEt/Z3VGFh3Dea3ZyHlM1z6Lyt0HIeUQtPzlDn9/exhK
SRPoJRoTCeNNZwxn+DkS1Y3t2DkJ6mXjV6e5H+2Dsyn7df9WJet4AsOkaFaDiK9Q7Ah2d4ZJ6Gjd
66ytaUNKYrjdwM01WCY1sYb8dKejU+OgF7d0HWyf9m5fZH3kkUc9/orn3hJWUhh73Y1m1Sd6Ecm8
CtXEx4clqBjyP7ZaXkWpILjl8nItmI5j8dqwqIhf1Zm22sYE7ve/Rqt4EdkbzjpXA11EOGEcMAk2
wg0JPElW5Is70GE3uDr3ez6lRx+N5KW4ZFfVX2AQ6b1OZ1dafmIRdbwODp4bIbP/Y++ZcyrjyA+u
vOslbPYdym4wn0Su4t4nqkDRDtvY0R5Bx9rz/FYP45XLt5/P1LPVIL+vyNPuXu+X5t8LpKUEs1HH
gXyzi6jDv2zSckB4TzSyHmdYAzicDWkVPFI9Ah8HKKEyIQDO0itma2kNkRGTicop9vaZpM9bFlyv
KWRHsR4rVFMTGazGLjOIcrd7uQsUKhuuFDKNpErCTc0PabFM5JvM15GaUBUjeL2SG9s3GN1s9JRX
4Kf81fcY7szlDHbFHf2Rlj3sqdwknvTHW2rO2pTHDYAyQJcPW+jgB2YTvmN7V6HC+cc98628T8s6
Nt9v8p6Hswis4Hkv5MPxflZFBy44Q4tUC8IT+WQLNK7KjY1mgBmy/J8SRfFPNPQUVgMqIXb7p4Pk
fmBPtuLiw6o5n9gY10QD6P4A/69EySCR3rmWdD3i5yVXR/lzW3y/PhvbL7V4ucyCxQRBVfnnMiF0
raPndqZ8l7OQlW80A+MS3088yAjifg6Y2uVRIik3nJ9ap1wObH2tympeohE6M/tgszxDyD0D9Cyh
l9oJfhwAVZNd3FCtBvpnYe1t2jPUfvQTal34tQXz/Vkt7CkvGLgMka3+cx1bBobF/GohyCX+QcMo
6YJtTnjP6FRA+atk5hlqoW7xHqkNnVGKWuzGl71zMnp0B7wUqZHd9cabn000jmp4D7zQpO7cvryf
HSjAM0OSWRA5RPsSiX8l8pP5AEkHblcMXSH2NEijvJMzDw5CYB/TZ1FmFgvK81weEdk/zH6wYUqp
86308u8PTcxwreF8q+VOXgmsuYM6l7Psm9nZHhmIAOMLs8MKG0CFf930yiNWf88Hr5Ttv27+LDfI
HNxI3R4MeLOefeJC/xATqJP8KwXz1qzmahgx27ffLlOPr/X1ryu1WQEWjKlGcnbE2Lp7p2tk/rDj
tTw7RR7HLN5uzhO9A98jpPN9oXUBu94Ec5M28A0l/MKLUvMZyALDCU5IPoul3NP2sbFglQ8W/Tir
QEE0q08tT6k+HpYwg6DL7lBfkIHtEm6yr2VWX1IlFDRb3SpBwFp7EXmgXj+yRo/Cii5OFabs6Rlp
g8JGl5Gvuz1goPHXEh4qgGZMwT4gldF3GI0qxMH0vIlFQY7vBakvdUoZsGwdecoBWvCLUexS6Q7y
novkUp0LKYRDQpyrbW2Wg85Ht3GLBbddUxbQD5O7SCxOFx7PK9ap3RWoRVNUZmfxPFVg8OyTaxJv
nuEtwTLxUeb1xTToGAzz/r6t2yf/OMlENmO41/IdAkB+HYgFthYRUUAjxxqBs3JvwJcD5ffwvQ+m
t7iocVq/RCLIfI3g3R+Id1N6nD/bqnLeqhkeaxtwBeg0B6C+SPcwlHdy/jwjEOWZGv8talKcbnLj
EKbRhOGZQKxq+6CC6isKyh37UI2yME5LQFWcFRqgR0E/5su+VOmMEOkr6HAFlVjTbFL7O/o9f2Je
Hi8+GZc/C0UUliq14UeZsv4tuQUu2lrgxxhw4hSLpWMLmtv64ShYMjEcB6Br4EDzLt+YYzwWrsz/
nIs998t/s1Wiyowj9/0suWWirwgnDMAUbpW0IFRXo++U57pyF5n2f/IYNmCv9Jypp5i6foLuAubl
wfs2SU7jJs+QsXGxleWIAhg0tv2v3nRuz2LTxpfQXAudl5UjGRSIBMEjeQRCCtHZUqU5ArqW/LWx
hfcscOMnwi8s6DXSGQl7F26mxVCgBq8omGl+k34lG4ANXhCTjveOiqxws1NyAGDyLc33Mh2ViuO0
5VndqhXPZpF8rN7mX+hOXx0dY9ii6MQIlbNrkfgihiHFF9U/q+ci7YX+nO63GGKE7FGLTxL5n8zb
gD6pNfLejSxIt6qRkJhRA8p73mugUiBWhnNEKtGqnqW9LskJC2ItMBSWWh0z+0AqwTPAFAU0U4fR
5AmEqqTaRxJFQIrRVZiShjEVHezshPZeuXPQGsvEG2rORaVg7XtQlTnVtQxnd1KZkWj7KAR8An/p
jkDzUz+kZFOO9e8QPw3vq93rSHNu+0pyBEv9I34zt2TgHWXcY+rbDwPG89SjpoSQhh56Z7MjY3o0
rmV4/kHuRqKELxppkaS20oiPZk+ZWWgeCW2whiNzBOqhHmsFCY1YktTjRQk3ICJ/KSTPH3sWgzK4
QKq9AAnc2K/DyegRlb5dEGdPP+8uZGZXG2CrBsK8Mrow1u2kKm+KMFewJRUcR6GpPeO8oPOZdOo/
gUewTGyzCwlPgDwcKrj9zj5eI3Twva2CioHPI5v6ef7RKP4Y1n5gXfrWYj1EmIPWSovVLrfWGbpk
0NR+h6lsL8ChW3MQziDWxk/8dIbqtpYzxYE668Xn/v7K/MGMKf3b2kJFVITvbp+54zZME/y8su53
IZrFSC4PWP6RZOi9shzI4weXeT4BHKpEsXilKKzY5lQPE3riWgrNd41CQ+RRV8xfbnt6zh1AdBct
q6XefKN29ldVPU6/KPL14VX6ZTsxJjK68nXOWcrKbZt0GIORaNCbZy6Rl2z63Nc50CovAJAwoOOT
fPlaomBLCD68Q+jywSw/xfSYNN+1RiTaJ0YvCkm6y3+YkEO+WX+8ZHCPyIEZuAxuD2881twuiJ9w
TP9ZGbob/aYV/MyMOtfMc0KzQvdedaVBcTFVlYJvhbywRPVhHURkERaJ3oGLufylKqGTm14YHnZ1
pepGNEWZuUbyxhHW5ydgnS4kVwoWCzkQJvq3GQKD735kSD0TufbFUENapa9EbRYHVJIm2EQgCheS
jx/s2gyTAXr1UyoF/fMEG2E/Gb+aKoYh98nLS6Qj0wYIT3ikl8kUaCRT7hlDxrIIKIcHC01lxFwB
or6xXdNP4YfCIbJLATQfYxPWfa5BnVsjULGjQ6/oJLV6D+9dY79sQ9lOwKKIoIIo3Yz5je52qiH4
O5Lf4FmhJUFbsMXpHb6oAs6qWlNMv7Tn9xzsD3D8e5zK7G0wdKx6Tn8vXxn96v+ijxch7MipkYOC
wp8caMEv1C2CCM+SYH94ShVi1UPlTS3eL3aid/i8toC379Clx2vaeWb898GfkGK9pSruC09igRgR
Mrybo964Uxhtjv/QPOaj35+NRPAfB7oM0RF+uFrdTOGsPpAWDbTJNjm/+U8pHiB0g5qkZI+RdDFr
28HaVMVOPddzb1V7CcILJpRPsh/rs20gipBSY/RS2mBvCkrgOwmMVuawOX9fzMtn/W5lmtRcRTf0
rfW3xl8GsVbTRsQxj5J5j1bn5EklUiNCxxgaUIfZsHnvU8cIo6gyKHqu0D6pjR73ZWZfhQ3SDbrL
dqWG3rhcQMHIClOcKSCHgN1dsPA28e+kplEF9cKRMiZ17HjT4zUC6kAAbDTwR1hcMYpvbbsbpT//
uRJSVlOendIzzMW77bdpGyOMNHPHrQzhK9K4oFy6oIJD2Sily7k1dOQ5lfB9KR6qb+fEhH9bTDm9
hMR1w80d3/kg0XvuPoWognUyZLLMdZYG1sQmZS1MduO0xOJnlc3QnMoMWTRBkBix8E0nxmrE9cfo
Gg8/JKDhV0mD94caGhoGSuo/7sIzllp8/+aAoDrFsyEOzjzD8YxRe7oFqNhwFhvXUxyz1/B/q45k
11JYTb3m44bDzYUYd9keBXL2UpICNlkGXDBa3aSYDMK3qDNSaYc7LmOV4mPlJxKp7yhn22oBoglf
5iBk6p0mhCYOAiLZPqtv8muTCkf3Orkt+sxVZprX1nfdRhEdNp7hJIKkNyg5EXXGXev8kSSMp69A
9UcU1zkmbeQGJpA68aiN/3jK/l0pFvf0jg9/HNxSx/sVm3QUh5ngtMuyH9Z4alhS8No6/E7BsZh4
ctreV5YxxraLhNa2rw7gAT1LiJd0ip8HBwIzOrV2TZcOADlTSnuNaWM/FAFBxGDzNRP9qJ0jxi7C
BzoA+gy4WYdgbtRICGK1bEf9t3z69M6DKb1fqvncTGPo6DRjkuO8ZM2/mX9QdCi+JUGUB10HG+uu
mOUhaZjjyoy7D/l16nqAfiwbQR4ponMkJh8nfsiw6D5hN/up4e4EXyUqoELn+Yl1qJP2WFz3KX+R
vXaBCDHzu96KZQlwEW3Ky/vbgz+M+zhTMRuNIwbu8x+NL1FvcjDPBtuLZ6UMD1QqKlTowq6/EeUg
up13HOfW+bLgcdbZ8VmamSbm47VL19oU4V1wFvJFKUM8ZghlXzy0AaeYBp9R17iY2kw5mGmts2xZ
WxHkhlVEqzhK2ziJz6XAJwBwiCaYm9aLOAxeDh74JsYzRPtD39bjaUzTVqqvQpfaTsN/lNlcq/+H
Epp09nK41KlGAchCwrUDe5+bKoOG4hdbIz3K7lLF8sMzTL/4UAAIJ53TZsd4BDVrAPen3Nbp2zZD
8VE+oOpNln8KBdTNkOXVqSHFnOvkeoq24ggJ35DzuesUC++1gWArSf6jD51b4ZsAdV9IV6hgigSa
oWTTm9K7fA1FqO50jDn5EWaUR0IJYK+DTWBRKmIUJ9YylUCHuLBNPR1DyupEiSomDIK6qdPQuXNY
IYEVE/cCLFA009WFxMkn7Cvswm9RP49Y7xZcKgbaJuzjx2KE97Gm8VXJtKEKz0ZElB7IgaCUU6m/
xdV1knezKzN7483/RCYEGTtQsTeeSO/xg09RFTQ+CJ7zl2gx9LOO/MYqjHh4epjEd3qzuUcKBPon
IaecpmTUq/ZuOjiDzG6EGTs7skMM4/aNHNLruW2Lbwj+buD6kjJxYSSz8UGkzl/5JdcE3of65Km5
fBSVIFRGncWFBFVKJhbrufZISe0Uv9ApFq27gkuzZXE4ZHmshhpoehPKBmFyAdvHhIk/4WOd35Tx
cfrat8XCMRb7c+42eVeZMAhSZuwdzIFidXr07+rHCw0OlWnToYVlFnYzac1XsFZi+jepBVRWTut6
6EGCUZufdUs6wuFpr0HqHq1GXq7C1uRkmG6N5e4Vf00z8WSfZZzIfBmVU9KIpGo0QVp14kQNGj6h
WrR4UbVXc6zINEkIx9j0UgqZOjsxtRgk0fje5bFe7snsIzZnBpIq4G2LhPLK7att9z59dMUCyTay
yFb9iR5MGX5+U1iV+Ry/jRTBH4koiWLBtlOSIS/v7mEDexX8SBk+ha64CxTlbFgckb0jJlP3/Kqz
DF5P+j1j94PvRdPpBbSiKrsg+NnYoPglq4iAkOgL9pgttN5O982HZdp2csfajp1lOY8uEsIdgGM+
7tL3RdYj1fBr4iKEDXdsT0S4RWcmItplIUgtfDX6iZTJ0nUS/7RLRZ/zSlDN5pyVvx3dGOC46cbM
zmdKW07VXPQ+y572oG8QVFbeGh76NdG2fCHG/2Qhs52voPq+8Jag5Ja2xyrBXXIhT1vwBJaWEXob
6wcXUcgWBjZqs2T6z6T2FIAQoX3RJwh+omuoYf8R6sQGndxby3zAc0ahu50fCmfZ7gZGZTXQ0VUC
S37CrXyNLSrhTfBvayudjUaQzCNYfscUvYia+qVlmuxwh99TaKuScQNtb6sObwxCaMF3YbtVkLe0
JTbq8/kPXUx/A2KMleZrn4D4RScpANgbM1hA2aiXNnBJQ6S5I2k99PE6cGRt8RutknkfWeMY/pmv
AUlExfdOwLR2z9CRT6bgYk/NDbNZroOiHypDW4GemupxRfpIrkn1z8DxO92qdOJwRWm+dbBloecP
WGHfxgOb+jtxeZpmqFl/K4JVBmSm0HldQ8kZq7ogqwfrfQGX9qaSfm3Tg6pnc04KV9xKZVC9TLnk
EDgzQbR/cKmiLd4uOPFWL2FgZ0zyAvcKl55EczwNSa++rmrgCLe8W8creqi+wYtWYyI5VjJBzWi9
rRBAQCX47u0lCM872hjiNT6dgbRsB0LMxlKFXb5sMXu5UyooiCqz19BF4Xn1SkxpJg+vQZsO8a3j
QTmy6zsPdkB0zUzACGK8SwxtEx8HzA6KXW9LWTuYUdxlNhtQL6rb+FSzyjBNtJwVzGFdRhZktDSp
h9TywyWlouPvn1LO9Frgl5VfdOccoxWjE0YDMegh0of+zo8MvXpBm2iT2NypPnoFJcDiLMF1x1zq
p6g99snWq/3FKvZhlbqd4ebK/HPVOp1gI+B9c76alP0q+mxlbYQbDc8ZUhraStbFIuLIgQnHnyD7
YXk1ZQQDrkwr0m7KsrxqmOLKy6boOOZK10wigJb8F9p4+TvZzUk7k+3xJmwh1fdeb7+QFIZ1nPLx
2vFaXvg+cqdBRwYU0boPYNe1LfU2Pe87N1a363wLgb3fSeUKOViQpb9hd2ft1LWrnEkyRtF7xqUC
DKOnIVHwmcfaYbDPdkvXELrQ7Fcg1W+mQpMxnZPulYEn9kH0VgiRfeYjMeuJQEm/CyxBSVOYf7qD
SRp3uqhnwQY+y8FjaxMXmOUdgMk4kiPsrRDvgtjAlutFedGug++5TWq5QEnFt/NIlKGzn2M+T2fp
2Gtn0YHRESlGKDVts54fsRUM1EQYippkzxjjudYj0AkDHYhN4egfG9Cid8SY1Tp4HehZIw6IyivR
khC/JW78+52eJfB1v1RxWQ6k5OKmmExGcoRIe5qlUFo8jeMM/uigyOkwflYOoNTI/5fbhU4s5I9b
NayguH5RTCJ7se9RRWkoYT2CJwgaQqa+qkqWMM5ah/0hr5EYl/r75bibqcwYR4w+ifp0oQlxEHtI
hAwbYdvq9RcEFJqjWuwr8VFbccBudcFzlLW5WS3LkW5V9aAZO59iBYf7ZaI2v9AeMXkt0SNHuEua
hdmpLAF7pB6rFOTDhinQQTpC/PyTEyYW1GP0GXxa73kgovl9/a8GG4v76NO5cIGPmD6rkJedIKRR
dsTCSbZd6/+1S5T9knKKGXanAWlcPAjSFPB+OpMxZ2r2EyUmR/KY9QSOuoOIPe6TASf72godNAWH
ysbrzYeiA7BqNuvesYcpphcr3IfT9+tO2TnRpwSuerRo1zE6jpqKJzPKZp7RFHilmImvRFV4Lyvq
m5dWDEiXVrWeR+UjZzMrCZPJRtsOYU11VsUksXU6ib4Ic9uPf9GwxySC8MZwv0+3AfquhMqxfd6A
IpOpNP4SoUZ7EhH9S2DtQwQDhIinp9fhw/Hwhi10Ybyj68ZncRjVEaxFWTXGlnJNx6/L6et1lOWv
gOLOeiMjNKk97EDpHZ0qrIarDJp1aZPsPRzpoVLSwjaIVZjw08n33albOVwo4vFryDQesEEp8i7O
jIvpIa2Vn5CB1mMpiF7B2ss/YkhCu3RDNEUP6El9LEvHOVEihQq7R8dOXw//BNeZd8x3wOWfAedS
e6tCUeF3xR5TCyOAB9jFxVp8u+xM8CxxvG1seTP5gnXND3Pe+vHfNf2eAYL1Ngg8L6gmPRBAA9eI
HKHOkwCjNORub/Tfkh+FLvZbckozXmEsr36cU+0CQqRM1QZ6vvUR6uoHeWx2o2sFG77Ks05/u+Wq
3FzEMH9CKRk34x87i8hZffnLAOLnN9yXGVUxIv9Vxqb0UTczTfK+JX+ijPerfJCm5EQAjzERFTfH
KP5wrB4JgVnt9Ex/2j8qVlOxmohDzZ4MFX3cr1dbQkHeFjd3y2XoSUWaByHg3wiCtJODmt0AXK0z
IfvgO7BwGayNm6RI10a2Xe93dgTJ+TwzbQEYYe6Umgqwam6kNu/bhAK7AYwMarpV+DMjDqLwimR6
gui9bOFQJ9rjN/8ZE4i2avUlk3fngwF9xA8LPczTjM2jk9eCN6wAzsHiJcwqLIWK6FPRpXhRG3GI
NHrc/QfhJ6fl752ywq8wd0aDzUNm7Rh/BMqLtqo+bLOGn5OJ6sv8a5Pi99mOlyuLAed16FS51i4d
7g5nthp/appVB0fIiqHm3s1pyl9vHZbWBoA3njXt8LYRZ1y2X060SHXYD+QSip6RlLGG8sJNYb3s
Cc2RLMp3GfdX0VuPQTvBbENmT6b0UMjW17mEagK5fX3gc8Nv5fnBmcL5Qv8jStYygxuawFFVHEmv
DBFt3QmhSH+/LkP9pWbxXVUGpC4Om3ScaFa9W4tgUIqXDpz2ivXfVyT9ml8D5OWzJ5linN2vDwOl
fnrUNIzFiYqQQv9nRahnvOQ7PuDkGz3uiUFFL8eZMG+wViwmDfHhRBUXnqcf0tZ59vr0LStqov+4
8Fd/xRwn781N9rHYCBlKZPJNrPF75XBV+hz1rTJDEfTM8AY8+sSRvkGJUP3bUQerHVaSnxzhd67J
WL2xv/aVWf2nY+f9tOISU1p4R81Ba7OFzLuufjmE1PKgc4Iw/ExJRbTWx/sHtQ4jwlVvApY68xyS
gGBzt6QnACZEhWJUpqApK9FwiiKrLVp5S8G6U6nHHBU9vnqFq5fxlpnPf0RlLk3IltoTGEh55k2z
LT8J4zMKpBbNa1PkiDp+YMH2Z1HyU1TUO4UTFb0aEC91hutlCFp/OPTAnYcrymMDBrfIu56C8Ehy
dLaXZYVgNtF/AWu1KpanK7+KMP+tseRyFenj40ihzpkeRT+alMKC23Saof2xwDm3bKlTLYw4fWa4
6BHy5He1UplL6+pOdxGDvsdxGT4iAss+DMC8PkkWW+hlqd1AoWSrFI9jYs9oF06+iBSDTLhasWoS
IuObxHBltU1JmfDKtt7XtM6geKUrUg72dgo9KySubdpJsbluiSr4sElCHjrY/+Am5GDxJd8GFYBD
/T2QWGDvbKzA+ya+yTWpZ+ldcEWIuoBF49/akgVvJ3xiVAWDt0MY1i4MBsJ1759MLU1KChFkxuMW
ILGuhiFP8yIDoP5GTPsl7ud87FclhRm7y/d7ZZJF0ZBi7AZUqOdcpW7GNMfkGkCTAPb6Y+7u5Lyn
88rZRHBtGQf5TTwU3v897JAEIhyDNREzNTQe7sUESneSQ/lvPKEG/Bi7RzlbfD3E5Nvm0QNmpzxT
TlygyGmZWmssetwIYLoRktanO5OfausT99XOCPF6fn5P1UShaoQYAHDoGDnlo9TlAaDXQF5U9dCp
5i/C+5NxG9B0ZyIKaZ+cU1gtLqubKHzad1URtjZSQGGJJ74Jd7uJbq3KxHO2jhDYALuuqV/w0T/Z
WLKUCI7AfcgmSp0hYv85gLe6O5o9oZ/J8sjOxjdM4xwkiPS57UjizMlijDqUzubdtOr0dbGd8uUl
70v34c7vtWckCZrOmjNhnhl9OPCfLQZH2kXf5XPaTbKP0ppON53CHZeLujMsRdqCdJ6cUfBCd3sW
4tgnKphDAsRFiZm0QwckmtM16s3we+ICz+bM8QyvOc98D5IITyC9Zh/mtupNfGtI594oBbfiGc87
wLf+NcqyYJxNaipaVb6ryU/I4W8o87H1GNTylDFRi0oBBi3Jz+4pC8Ijd07Kom+wrmS/hy8d7aOS
jZ4bb+li2XEqyT0QjIyftLrUxIuRZ62U3xazXzQOPyRfZsMyUG8ah2bW+uXBlGS1ajAnQeO0iD2S
JNHM3QRiUyTWnsGOF1ZnEsPIGUhHN+Fi6NL6+rrXmB+yp4hABLQ+fUJVCfCljhuk0IA79El/m7bg
A6h6ZSvZRNj0oWIJZFDOZLwLivwwWMWB9H5pweg5+h/UUIPimrzzrCGKOCQqfRHKAYFZoFF0jmXH
+X5edvrIgjGbPIV0Z+R4t6HoDdP53btERj2AWvsmxIEmYI/mlivq4VpfsU6yqFP6vylsUiSADRWF
nYsNQjNZnsnNeh/qDVK33HV7OBDG1XLXEwrJn0vi2iC44mxhF4ULeN9kIrimoF8qD5iFhHCtTVbM
AbJDlVlZyM7rTlnh9d3Zxd/Xzg43tMHoTLdCqFEIMlgB7p33NY2J8ZfojdvXaqN4Zf9z80p4owUi
wvRUlDrb9lboA0KU8tccbszcWTpENrvnKkZjP0AwDsb3QK2uCs6WtJZM6xm0YQsnameGe3Ke27vt
u0UP4XoniYqLHPFhKUkwQ2Zqjkv++62yJcFg6Uwwph2mK3dZ5ErvKuDxnpZiNaJsJfk6kwYdq/DN
xqo0EPEIsjgI3WMRYQU8nM9/IBvVlyuJSZ1W1tCg9xe6joVaMBAO855+sWCOFjFUtWUMahFFR1g+
PCfsdEpk4zBjFAhhzhGPWNGv4NZE/rEy8C3h2a+7//hWKFpVNKaM6sTKC86CBMdnmrR0NBKJ6l8+
VuciOgS1v9BOAFyg6YP8WbvSdE+dYJS7YPw9t0AIP+/7JN0ZFygfzzlXaokiJGG/uWp7NEVmizcX
Oo/HL6ycubYxUotxoAeJ3/ULVyOgoWB0xJ2067OsULd5l8ny2dMUaBrUkWCzdl+eMjYVflxLh6hw
UW83uJFMLpiIpQr74k9BW/2VF18wozF6nq4XKUYQ7dhuI9WN25Hd54YMGmlznCjDXBecEw/zsoLU
VjGPiVFO28AkgZgwWOHUqnTXFTb8oEaMIMCjenygjaBVpvMdrKr/sN8zKvM+fcHGdAcoCLXGJXFp
DETxtTtw7B2vS9Yitkbp1+8S/y97Glu3ocCO/Cg/kATsywBlg0kMCW5mFXR0iDfbOEQqJoyZMJYC
hiwZR1fDh/AGcFCcu3y4ModH6VsclmtSb3Y1maYau+SYSEkkPBjFprkDau3G+kWE/UoALk9T/0cu
XCZ4TRjTKOIrRcyDTk6u+PCNUGtJfRQLRXSkLw6IFnfhyaMEIqcEadFoI2YeSPpTsINtezenq2n2
BZCkUDMx4G2IhSF7lqeztzy+lNOBxpz4vNOLlijCJ1B2OnHMwGL3I2vWAQO5f9q/PT7TL59idwYL
O/0wngfTeQZ+TokMpevc/sw/DtFmcmofXN5xqGTDt1DYACS8L08uo0/idl+D5fEO5gK3+c3xcltC
jRjdSadetDEQMBfEn6Bjdcvh1H4bARL7IipY2nDy9yaDnrbFGRihG6pRGiW7oUP8HNcigddgRn6j
cgdzLAdGESL+VRs6HYJlxjvkqV/J4hdxWloAIyIkUcQXo8vquH9PwHiQisawjqcoRlWIf+4g5qDq
KQQzTkDdHkbLTfHjlr5RGDidQGgtwp4tQV/ELNecskkkvmf43fGxPuZVPWV0c7E6DHqDRijAs0xW
5e2d2WDMj0GmJnanzkzytvPWEqalsb+svBQjMbfRl2V4ljp/T2xCMcLPD0AGjjzg7M7x5bUpneo4
dJ1N259rQQiY1EKTHFKNqeMaZQSRJNR5+IVxmKdLQmoSYQr8BqsoPAtZs00OW5hDUldomttTZ9T4
nHcH6APSB9MgwCS/gG8o25uzbgm3rZUV9dZ0szfwYniSsuUHHXyCP0bymsYR+tLDDHp9eiCuUDqM
z0J0x0UmEEokSraPvJik5qxn574wKlVQ55fRbNazcdNZrW/Pyy040u9GQC8NsBGBxVBQPbyB0VN7
GxlEcmaQbQouYYLdH/Zs6j4JI16tME6U68vW89wOS21SVCi0A1cESAZnitIyOhI18D3CTp7+fH4E
koFZRDToI/MXdIAdUMZ/Relh5Ey7HZ/maZX6B9eL8NIzaoyXyeNj7oyOH+sCLnR80rOtuC3i4o3v
8JNExm1QOVJ6zLb4mbudrio0X+LPlDmW0n8/RbOznVtgRmC53teHT9ss95WHvCr529zTZinXKi3X
Io2tWbb1vJ2emW1CUx5KdQX+L3DoUOfYFeGHZLHSVafQUccd36DfizFrwaCObsgwF1X6yRYF6l2X
mSzAeOgc9rYVeXxo/VQA6JNwR+LKPA9fE391W870RujFnSkCzyaMUkOJA/Xdw16M/qlAdMDx1lY6
o9kEcTXZy5rY/8BesQDYs46oUhvTbfiBJm0gZT1oNrlqLIm5uvMLh5vxBiMMfM+RKEywnhBJue5R
0q9ITwBJrzQa2leXbETrnppOicKD4wUFMlLQRnawp4WCjfGWDcEni9OeLDFVyKr9T+W3XRch9glG
DbeNoDNreKgEGjQpxA/DF19FYrkiVJb1LikwtiFVvt8T9kn0ppz/bsECKzKNv9ZUUOtLfwpAmOQE
tNRJhAhC9mZet+UDcFr5EGNOSjK1koWuxac3utykhI7fi8f7v0dbpLDql4nui2ysuzzmU/FIADDy
ZzMP8GzXtz3w9hTEQGV3tuzJUoAXCMiYnlbroT+0eeODwGe8cXHU2VSeyKH+nX20dM5kTQfaYcUW
YeKuyGffxcJdck38PMrQ/vX6mNzama2OzCwxtpdzhiANKiSxz2uZAyy61Jh+v7OemHbO/fUempiP
tjmSw98JGGaQlyKTYY339JszoXMdC8V/I0p+buOXxC591KkfCjMH9HhxpAc5QHTY27/AEFZ6yotS
BeM/acRpx2HMSyLyXl6gJ4P0I1WUs0T+q8A13S5cR7MlwYAf0j2qGtH3FHlcfz/j48WOSbNiyje1
qJ7jM4eH6LoPbp6WB346/4L/FWScKOMU667WAkP5/DSlYoy0iXYRxOkDE3EQUubVPV2q/j4e5IiB
QY6oSAvBpOdBZK98LtqPelCWff1paGu5xnn2GXm/6LrGs0EdayHhymwwREEM+SOnkc5knBxux0H3
7SwBzDlIG3b1HwppC/kS5f7o3O/Ydjl7R3PPKrhUD9VB/ddCg8PAzSUvaN4A2wUSCRMw/Fb3yI4t
sjIF7sjwtXS34OxIKRVLBCoBsalUY/Gm0Cj7t6QOiqw0pXFsddICVkpvA/8r+2yPMJ/9rQoKWEKi
3XDhzrZOPbj6eLnWzFwnF2fzzNtHcBYRM9s4Wk0kecaPOgor71GTIBof+lSbssn0Ji1lfBKl3rYE
LB/gZKTvoZmehPMilEVr3uUlHboC+s3pG/R7FQ53lHgpR3RyxBySuwVmnu2f5hRlSmQMnzuBznfG
kp1ItkLGwrOQhbT2kxfD2TMjJy5fEM2222a0fmXJtyB/g9Q2bc7dADV9CHC/C8hVLAOSfZkze+o0
4wxCFf9K2q6N590jgf2W2TQAiUoc/Z44fSfi1CrjWwMoer6D0fxrapfOyDDoJ7nTRxgWoN2VZLat
GmoAoE92w6xhgJF/CB07HVxyUcjWtU1lRvjtK+aR1m341jUSyml9m49fh7eFVU+vvXPjpNLhO1jK
GXExKwIClM6rjmP6vfFJzRSBBWSUTV4Bgd7fa4nUnQDlamPGLU+CCyLs/4Fx0i0IUo8a+UPmpTSu
q24/O53OuNcSPKSgrO5KCgRo/GlAbvxydjXjxUIqc60J6S/a3LpKdUCtYKBKN8aR339iRDNdxeZ8
1aYKo+LnMZ7Pwh1OS1K9nGeZLMVUHcy/YVk7D++GdXJ+WV6Vr8x0QeL5urRSNxn4TwIOdMna1yVq
NqBQbxqQDQ+Ggb7+wLTuhi6OcIoA5dwPyFNydz5fVm1C4W22K1uBBeEpkVNUB5TKJqepEbDRI31c
U+S/LEXQjpCfvzDhFInzmts52quuJkFRctYjQPfKBPM10+N1C+KfIqcxhKNTlP17NXKRrl1nPrWg
8UXKoUhklPKmFxV/OIyCB/cRdR2+C0Sds3l09chAOiOsV/ZQpgRd4toCu8q9oHRs1uQcX0V3eMCO
gg+PmReOQFx44Z/QCQZfYb2sZsyJ0nLZTk9bFI7OdYUlIPtnrYSsAKsWrKSd7RVzky01FOnIlvVF
l7r3EQuaMveVOyhDh2eOY4G89tjM3F0jFHsHjIyplk//Pd/0HUNfh7yb2Rh7fI+UD21gaHMV2eMN
XmhY8oLgdRBs5xUIE8mjXVEnCOly2IX8r/KsjlRi3sTAiR0pWpdQ21LBe+wIW1yFcyQR+yJ6Di+o
ZLKLVZAcoPEZ4nDutqR/RR88eRtBGSpI70tv5MWaDYntXK7U2X+6j9DqVnCQEbXNwFohMMHQ1ZXr
i3LwjGjpWfv3xBqZtwUJlwxRCQXXIvBv7uEa4m2Sk44l4KfB/TKPxbI8pohV2Uc5S2oHrRsCapZO
26oGUhKeSfl/n1O/pu3jmZUmetKa67ebs4KVSjS/G0IZ0KPJF2z5IWNKQGPO812/PRyBn44yYV0T
wQ1ZlYpwxdC5Z6+tbD/cV0tTTu6ICu2wB3xJ5lKuwj50FJLJf0oqwfsksf25vtLBNve+w4twb9wK
At6Iaj1HGWRV1O+i6TKCR7V5xdaGQP+07NJjMh+mVQewzThnVhkWjVov7kNzInGqFiEhxdXY0NsX
DCbDcDBrQ8pDGS4VlDkX7E7jCHmPj+4K4CfUbOs12teR2A8x5ccnUuZH9VAZ/FtVxtsCMDo5i+8s
Y5ifDwT8fP7OfHQ625Nuczajpoe+1VXTMAV++iaYz0a2+wlyFhBzWAvp4FKhz6xolaH2zK90ItJx
tJKErtuWD2YMCg6AWSKwWNNyC5VvqAdI9Gq6AdkEkFfbGh8UYbMjvSICTt5IrUCBDVOrHLD7fB7Y
9J4j8CTWj02tNEaXLBYv7XVTY3I8mQZVYVk1Ih5p1fgj+CNqzzor613i4kNfO7nZPx6KCPpoIPNT
qm0j295aJWYv3sR+1nYZ8aXYGx9fmFr8PWnvo1PWbeWyky0royR78Z0Me8Wk3RlB2qQEKix8pT3y
v+q3ElbEwdPzlwJVoauVeUzPMHulx3um8XrBIPM90quxdhHrZhLBeYsZFCk9rR/SWbFQIj63KPxX
jvWN0++AN47t7I9Xo9JJYranyCnPar+4SxhpBv562LLQHbrojSL6sNKoO9oaBeOL8UYNX3Q0wESU
k3mEbcGDFzAap0u+HZ4KzAo7yIGrxuzJ+Rm9CBkCsQb48L7x5Y6KCqTFId6ib5Hx6eWKbcqiHIbd
CV22bYuWN5yMT1wg6VwFuqqYIdlk2uFmGKdWJF3nxbvIi6RuWCZbfVc8heczkNUsnmOxPd+t39Pd
eiEmlLvDaGo726cn+MTy7WaIK0eUxnjZOR5feZVZuB8kWhrHyRnCSqWXAI9CW5vYy72M/tY62zJM
QodlxzUJn8dRifBRLtvPPH3cwhIdGCoNwb68D5XJ0/WPTFhqTTGa7peHTJi3cCwIviVaMN5hXDF0
SGmyBuSomwv4Rv0NoyzJ2CahmHtHXXPo2ykMSltLsVaeWlEWyxjDv6k+Y6UsCpHbz+zJ7FmShjHC
gnF6QTRt8o81CPbdJNrgUrX6Pyfffs1Nj12U3ym15EMosv6MuaUguzu673m1/Tki+xwwLuEnbj8N
fI+oY9+8S0ctjUTbZz9qPxDtLcxpVNB3oIeqiunBVQYm5zrvWaU+BPlS32fDEoeH4bL3QxQT7cE5
+zL3HEQyga5ZyhU7132rhcRY2Sty8nV2UJxVZuzj+w9ZOgnhecwSOlJJeXD3Vixzzxi0MghCTeC3
NsvOjpEl11a1Ni0A+6exwcalTwf/vqlBIuL/h/+uitwoYifZ3cWv5PgbcTddFh0Vqx04k6wmuR5m
t5iEOgp5FjHu28hoDyJFrcNA1fLL2N4X/kkuuwfRo8jKYE+aD2b/gDOdhdzb7EMCNtVu9Nilnm5o
3OohEWAXfG+HPKY6zNRd9qbjX4Pgl9mCy7GLY610gjdX1IihkCXb5SzqpYHiPmmX91vqDkmHsvcn
+NQdJ9MtTzQFTr/jIq9o4QU1y479xvzlbHIhMxO2dCK4yyHoYA9CrgFnB4jhR0195HkSGM3+8uwh
L3Y72M41FrWaoNzDS1ONmM5m6OJhWysxp1BdsycGr1NEaPBjYjsHNgPf6P94jGInRgdoLES4XfJK
QWjNIhGJNEOUjOgkidJRyc8NMA7HkXxNs1SgPv4PpSvyGrjS121VOgTZ5OoPkTzK3wjlzTIaz4/o
0Qz2r/PvvSNshzg3N6aB1a4DJolcg7wmFmWxGMQBjibEyp5ZXeaXatjEOn95v9WhD/jFnS+s97iv
D3ITfOw5AwOGzfqNoTIpYe1I3ATwfEez7/qGcD+pHx7eGU017+eBRQZRcaliicOomofiy10D/sSp
NazMkSy8eXZaD8KtZYTR2G1ir/2Ry4jQ23oycPRtIRM5+6s2j6nnzvjC3DjaA/SdibJyWvSE3q4K
2A9x8T5t1ruX/oEjp1Qv5uEBvmJvCEpafaPydOgZzpX8QaIxoco6SsY5rIXKd92+HHe++klR5H1y
xKbaf0KcRfOviQY98/Hq2IjqpZBKFX5YvBqMGLZAz0RqwLophPfTU+oTG/lmSzpimxhZPi8wUzXh
wNqPvBKa6KHN73lHpnFANrs6jhXMSTQ0UFO2i1PFpAcROom+1gohj23xHJlfAQ5uoWeUftPQIAzz
IDcCNOXa/iYssr5kH33WdcReivLzirzCusbkdgNJaEnYUFQB3VBE3f2HbFDlmyiho+vLt7UatIWV
/ZLohIKLLXlDBsSEAEoOCVuZM0v00KutptrnLKowQJ9Hr3oF94AyW4v5nrtnM4Okac7ZZ4jp4ZF9
9dYUdHL+TI4mw4Avbl/fopmw4MIkiHsEk0li3vrIDVT4uCTZrwlG408e0rEC05xfSrRS6tB+NLf3
58eqn++gL2TV0x780h0LMjNYdLgcpjaAwfsoiqiVmQp8xmKHnef9d7KrdgkkRs9pCQuUFxV12Zfd
Lm/kqhi9MQNybweXYAZfbBKPTQsnX785sjHwSl1DW0aFdNmw/GQFUPDVP6rpuslyr4nzGp+FGG3w
dHZF7NRxF+EqUVyd3aI0euxdbiGVONkxLqBo9rEdkC7SlxhT02dCkYlDE1bp+J7Y1BczTSkVoYIv
4vfzBZwopvxGNv869vLQ9s044xEPNZmKBGKXje/Yf1RrVRLtMWVpDIBmJvL0P0KYuFun/BzVhIyj
dgAXik61SvPT8IuKhvdjyFbQdTPl9x3Vg7byCA4BeQTGo9VLJ9oCH7eGy174tWziweQ1qiYo/wPy
hL4aaa/aevYKhjSL3Q3MAH4JhM5luZOrgu7mkQx/czYpomtc4eL+Huck58szYs4rD70ZAFIPg09S
GGlNiXzx6l4JOhzHe5YZh/+ATeX1m1BjI9r/L7F60/gKnLz8h82ePWOy0baauvrr3oeSk1Mwwd4x
2Pm1FWAfVlpuU2ZQpPnvxGlRkdT4GxLFw7kDo9+IzUWVRlArnDPeS83hn8HFvtUNfIc6foG17xbK
Tgq8ftbYHTaNdfBRJ09Vc8rnEEbzguc+ml2s7MwCRmgC6XtOUKEhUzYkJn76T311AiR26pvhcFXa
tnkpVaaU958bkeCdzv8/1gG3l2uNZI/ihsmYdNTVbjltdKC2i/NpJYoQe81Ly8t8oX0Z9YzekVmY
uIlxhLJr/ghLi9n2ZnYZPGzel6qvYo1gUdGxVA6twA4+Umc69eFaopqFnCGyaaNabnI9tS3v/QzT
UlZakN+1rWCCp6wnyt/CSc7vkb3C4BnlneS2wqolB38I4bv+zrOEK1CcuurXXrKuIfJ68j2qh2Ag
vYXmZ5auf2FPgwlmQFi6qzGjHgMk4iE26Fctcxk4dWxNDxY6fIG/cQvaZPehGMH4/SMPGQlg3NLw
3MGpKpRlHpBsVLKtDhQ5Y1k4fiSlSf5Sx0DsDrKSCyxN0LKUj2C5s+JEGK8et5o7JD1OYeuurk6n
AXV/pMUss7dHAYHgWt6n+FMtzy30GF8H/sUP3vRVhBeVJw+S9/s48EegPQc78WNESdH6acRdcCft
tzfKrUCCG3ho6rNoBHmm7W/V+flXzUNPIIC6d2sMwiulMeSlRMRdK128Z2m+Cdmfu9SiWZMdwaKJ
hiLuIgyfLFiYFBHJLYrgp2QMwa3X6zfqDzqJ6Fc9xQwX3erRZHxZTFGQnA5yrggM6IjEcGeagtjn
R2pIAobEJobeAmPIdAEqF4YkcVwD+O/wvm9JXA7N0Bwp3cz0vLaO76cR98yFHlHNaU8K4r3GrL2w
xBJ83VCEMslW5hsnnU1bwHYrAzxRdnJWfU3WnqhqiQCZKYVvn+OrVh0MJmIuK81noewc/hQr+NwN
hjL9Z5Q1Tx9zlC98ONjL8JKZkKq5sQg3Y+WUF7Tux6D9U9anDbPtRRbjcI2eZmfyuK7vIO7ZEMeZ
lPBu+lgnuy2V3KVQtJTlmvgLBIA2n0BDPYPeds04bvxdDsVnhVi0coYXiQvJLfBD+od343JNMx7c
n5KrTVPTjWOKyMkeNNUr0OeJ98EAop0I3QMeP2Bw7//gKaTClfDp2se9WubPk7r9SbKMXfiy2HZy
dJVaSeLE8fjtvMO9asO40ki8MXNuq9AmfeJK+hVGZkWq6uSgBRntlLrMgYJNQhMxdbJ/gCzVRgvS
88oAjsb4W4CVLsWerffZVn6LaYRz7ap9NRkiEGAkTMhgK+v89yBxvel5iWF3mQyzN2ZLU7SEa2kw
r+kmOcMmT+j1jDn9WAyE+M473QQXMd0IFT8P6Kwm1UFJWnPoyVJ9FC4/EkNbCN7OY2IeEETAi3Al
8+rbZt8ZMrIk5zDnat+edyEwWRbsis9lSAMBttiKtwSJ5Rq8u3BIWUclv6+fc+POAewT67Yp4/a0
Z22d8l9QWayZhakjlw0VBGHynp8sgvhu2fkL31Ye76LOmjybiZL6BSf1456jG+THR8xiiFihTw1o
aj/fAFctlDpsKr0xiCeB5m3oHtqBofbes+ip2vLjqE9WgyKnOEekOl9Db/9q22mLG5xJ1iOIf+6O
MRi1wJ4eKf6c8tn/c/Au1ipiczumj3Cbp8dFTRYkdRmdxzwlhNS7vGCm1U6UZU9pzD2udCBAnEqW
FIFwwgph+gsMXnbjUYWepY/q/0df1A8ZPKOPQiGoC+QxAKOGjyGOBrZNAsdXVt4npFNPfRaAVQ2n
3zhkMGVsM0xJG7/lpotQNONt72SsvLMXFrkTLsNucpf3A1j3RFb5cbVdgFC9ylNdOOe1iTa1EERE
A2OBsK5T5ewZG0FFZLziSjooGjiG73uYEVRkxUAi+MTUnWtVR9pV2arMepLV8aB+Yb5JvcZNwsTs
dq0wmCGD5JxpiZ2XA16IKQAeaCEnxdPUf+/zYZGXmYiSPUsZ5klARkE8/bYoUiWeRYecpFDljpap
ueYlu97nY4TrpvV5P454rx9wjRrMt85Z4lhW5L3oNK9nGfX7q+vONXSbxaHPqjK5QjWqVPHMHqnP
Ig2ElPHBMbvFg8C53h2LxqxDQXqgMliRNCElQMok6OmAhXnCfSGPJKMVKhiDePnS/hTbnwaZUTja
dOsCZNe+FAqItF2FMZ0x8LPb398PU7cYlW6qSvQMdyvGpfqaBya5o+k1Nkxm0LqqUNjaip7xh94S
xlLbV6HeYD9HIAloksEGOk+y0ua2fXsuUn1cWpoIBq93Vxh1tzJnMb5NUbzLKIIrZM9wArF108U5
qx1tMvLypLi2LCADOUgiIiGTLeRK//RgLcQacdruLA7OENbCF/j8OgWSHUabP9q7F/WYl1d9/h5K
s1fuulZ5959Rb2fUwRY22pbyyemvS3cX0DTxYgxlfBIYConDb4aMaHu4HpwrA81bWRYb6ruDjnEx
JudbYGcKEk7kPTlZXDMfDVxS9mzD7WKjiiF6icK6LjL2hKV8Yu+CHdWHQJtQbBXTGrX8fmmDi1uB
5tOIdBhuFDKkR3RO+PwVLoByjANdMlvfU4ggNmciLcGV62l/PrTSDwPSZeKEs4nBK0CYI9l7al1h
VqE3KDGdOdB1RkGDcd2TgOzDt9HKG6cUUiy5Beaouh4sXuNnVE2iFjv9g4ZjNMyJaZYGSCCsqxtv
EuO8iEWlnS+Xpl3UtSnfTRJcddVQ2D6aKPwC+9Dguy1fdEBM8231LCKF4WdSOomWsdfnIPM8C4py
8v/qL4ZPay/bNR5IP4UO73FRZh+WrPJi8kRC/Fss4Ws4ns9pTve4Djt3l/8QC6IouXa6pbsbw+0o
Ba5IxOlU7MKTByNhLhqf7jyqt1eLa9LhxqinQyv807oun/OWS4YcctSN7wawaMKLiRxHkB4saESz
luDk+8ybRmI6cq0YSphtiqwEoZ1IE8zCbNfcn03++ZFwRLLZGLppBo0apa9UVMXHFPkajGWKhqcx
xHghTvk3ka5AnM6oOowyyd6+zf9YDz0yu3XDLd+exByeR+wi6UqZ02188bI6OHCw32jpi9odW4WF
uAu8xVIhq98ZK8ypzzQz6QTox80ECGd1iaUXnhodiCcGkcxNlSG29vWFJ2cnyKZILwaEEECKI6nS
Rl8PEqXHhxTYVXFu5gGA4SwFmcF4Edk50OwSTQMS1ColkX/s/bk3oICjvKv4UTI5Ku8GG8Ek92IE
tqJIenhLgBsATAfE1KAhKmSSAcemSjutvtUPY+EIK9zMwKO5VAeBaZbIHFyHy5xyqeDSNUFvVzuS
zl71RH/2e01F2o0PfYTh+RWkfpmvkb3hjwktzzfJeoivccYkOY4uPYLDFQHdGsQ7SnDI1QNXBJQk
fU4RP5MXD0CBRe30dl1gbCDHtdwpyBMdjlS4maQpe4IFZNae8PobaKChV3POp5eEpTAAazgGt9Sp
y2jiPrSJCLvXYV5D+wIM+iLctsbIYNSFXc0oW6Ed//pD+dCH8CIW73xsw1uItwZD4g/mSFrLEMVw
TgrWAZD5FzY+Y7cM+vPEU/bTNTrsaMEO0k5NAVKISr0ALzznq2lVkInou2ktgyGjF53Q3TAAY/Go
TRNFHDOdS0oHEPAsRbcEaUG6KkEFVtg6fx70EFVKrhrZfpVXwh0+P1cbNfgt1Apsgu1pjyTVLxxl
imd236+uRxx8hVu3IQWzXaYEksSXfmWYq7M6haBu86aaXGXR2og7FPgaqFqSXW6j7arUv5ktGc4v
pb/GZZHMMKr9/iL3wuyby+hzjuqUui3/pvooYh7A5wNL/Pef+6LRHM5zs8cC+CYjeviEzZSS0bLY
fhAfJ/SVtUE1c5R9Z6104ofhFyXCSevVh2HVmOa6O/FKNLiB/hUNDh/Qqn5OEJ1OEFftkOQhb6Uf
ycosGGNk7X2LQy7ptL9pdX8Id/QtIfgIt09WuZn0pyPL2o1AdxjoL2J4hun9kAOiegsuVONY5GcQ
u1ADAzXxKvozc7uJk6QVKv9NAw2ozcZc7jQbaewGot/b3SuxmbK/23anjseoMWKKzw4SRjOYC0g7
adT6MpLsFeUG2CWy6z9p3XkVGW8Tg+W0LGBRPpYBMQUWOW65QSznTqTHHv+6DCMrs3nmiQVCEIlH
/Saval3DOBN3Ge074l+BVqAG1VV+OzYnK4D003ZBkdpfoSQhw3r06r60Npv+7tlVe0DTDMlfZ6Ol
CkDhR4V1riBQNKJEXnlFrZ0LKvxzCjZU3sdZySRyEutqGOqHqqkOL/kwhOc4OABG/u0Vs8ukvId9
Cn40EzklgMmRadqTr6x8nTjHBZ9P93SiA51bmOZrKNNfRUMaYDGq4Z+SLo2UillIcpyKmNX7inEC
zSoEVFDzz990gyzPdtRHH8GFXQHpRGo9PSS68GMcKmi0X/SrzJK4IYubdlW0ujg8zV2uu6XtTgDL
J7/dAzLbJoDzFpcx6r/hXWDsROlZY6PzVNc5pHUiZotTd4Yu1GsJIyiO7b3va0HQqnQ/PABdUFgs
K2p+lUj4EpSFklegu5ZkQV17mfZfPnWypQ6WsM8JuoipztzXMWecWAd2DslNU9uz5gxV/GXGEGUu
wTf6HYpUHUV79Y9LSDQ7z7CiBWAYcwnQRD4jHRh9zSxuW8/SZSXFfudcIa5yGoKVO5gwnfkcbLFe
A/gJAhNbL5yLi+DbIpTyKq2fJlb/odYr29THh2ybUKypB130LQYrYVv/Wvl+IqMNKsDR+fHVvZUt
JDFsvOv5ju0WCj5+SkJHly0GJ/wvQ8c9lovLvwjlNqqB/YGH4LUnTRUSAaYOkrDyMXO2J9bYuqKY
0VuxXk9xo2HZZJlfiHzAP3tVfSY4OUiq6+2S+u4Zs7eW4ioUFZ5yidfY77MHKDnHfharqrYB0HCX
7YKBKxxMk8NM4vQwN9JG/o2ER6DzHsy9RUq2b4hqUMatH914AqJtjM1QYC1M8qhXpDhxL8sR2L1m
Cny8tv/ry5of5gwtEiq6/eYgFH6ZGcw4QXHh0gfuWRkuYyrxjdveO6Jalh99qoOcHmfnBXmqnOHm
NuO2FfojCUr6jJhVyN9nVc8xXPQGgcDaYKxHTFD7L+4B88MUSWpfw6dUTdQrZqD2r0Ei+mIMkyAJ
yx9/YpaW8bSxI3ytPF/ba6BvRSidAohtHIYmDpiMWGXkbURTriVXI0H4+T1Jv54Uvnd2qbqZ7JX6
pwNk9zQAXHRkD/Y+1SbzXU9mzdTLXHoCxj99GTY9agKEdnqEqNX1GCbThgsjMZzSLcmCzECbyJpO
gN2J1EJnt2UOSVt9Xj4rgYvnom9YnGPhSVF+/Tk/ddqbDt0k6AyGKso/We3U1HN9j3/a13P/wOg5
0PSLFY2E883XvEwtNMBga6wylRBk42X4DEgPKO12x5RmuI2RfLWjeKsyJYWFq+uuIYQ92WqgGzQn
kQ2a4yPV2rh9o34DnnHTeUs45DGwWsHwFSOCEoJwVDPkHZnrVraCqDDYvdsQ9qy2bOTFJSlEqIoR
0N9bi6ogJ//4ExtcxKmZOMw/OSg6jTKZiJi4P+eX6CmSZ7YsdAIiIijg+cmrK8Q++7IkoENcz/1G
JG63Pt1CMgH9PLCRoXU+UBmH0Z1i7ySDWAiZwsNuFA/B967NGKe29oIOt6ZGvQT/Jo0T5aHWTRN9
oFqAWeGwEkwFi8+c+wa57K9/Zy7Dfn0nstlxJVAXm6rr6/i0PMg59i5bZx6jRQMwIGmZBd+1KccD
K9sMbCtTP2SAc0tO4/d8ped9xMk6GQR4Aq4PwiuBoeMnqkgl8LKNKBBNLQcKs/6Zy0ZjOqBnxy5F
p6SRcQIXbafkwHJCLFOJJDz/YNfDOEo3PS7mPTciXt+TUOUxVDsVXqtC8l8sl9j6ftdjIdPlC1tt
3CO2qOqn2Vebmf0HKwex34dUX7DUab3oZT+TjEn6+h/Y+ULl8qFF5I2GCGMkTpunET6PivhLxLLP
x0y+dgrao8Yn0JrROFrj0YcvXhV6n3CnCPGRn7rmTlYeW6k78HvZR0CRDlb/i7oHXWvCLvIRTD6k
C78gKHhYqpUUU56CiDUsGbj4xIthadWwZ6t3z/UlhoiUAWNRxiyowAItm89KTgVoCA9SthLOa+IP
UBWMqJQx0SckcaoknCWOd8AowPN0BDHxFV1pMCHptO4lEawj+kNgfRKl3XDBj9ldiY9+VeNcx3CV
8VL6wRSlAkrbzq512lqOmg6Mb0tghtK8JnpUuiT/zvoK2yKgBFAMx+gDqDlV0zIuylvcc1k9j7pY
CjtSY6WiIGixwCn2jG+u76/W51n44x74aqaD51ncRVFLyf3sYwx9oO0SPN+ij+G+Rem1aTn0RL/w
Fsq1mrUn+08AEcRlm6uPWjPTWEcxJ/DJUN2N7QxfX8MA6kKbaIUKVGIBCeWw0rxHuSbuz1pJFTAS
jIvXT910Ey9SKKWm5vqVcfWlsUC/qqeyhXj9bcVQH3oEZnb7Q4Pd+KOnVVDMTXNsmBRhQOGHFWlm
upsl2DBnlN+IHa+yaVub6vbO//E+IbIhDwjiBYD7YcRxdffYFcOHo2QhU4HO/6oTpi64oOZHfpcW
+BXUyap9Tcqt5g50kEGTl3DWO9lLxkw6Qbf/kPPK4sw9iZJh7kPF71fxrT7sNzuUTleqCAfohjin
TovFXgnqLPhM228aaRd8McKazBNHUNhnpaf2Htjao8NLARclPe0D/rWZW+UyF6XsYVUmnhTHfx9W
Rbk/DNkRw40IqAZprZ12i/nxo8sJzvE/gvUCRRXNuybZKiTr3t3iVtwaSBg/0eYUqMZRvHEguqee
zeImBdrOpvzh8FC5syBzTpA2xsOr2EbukAkrImhxgy9cdr69oTfPWijMojjcxg1x/sX6Ku0xClX9
OyMZnQ+WtL3A1xwyYp+HxupgHl85/Zb7kg90dFuxzFQTf7QIIqo7SMKKsRSqOWUNnngyl6nZAlZm
tq0+1q3dCsI0bThRQbeygCP6ttr58dPsqML1XNxlvZ8BSMQp7IceYUygA54EBT7vTXgUqASB4fUk
Av3LXF4giVSvYVdcraJXbGS4ItBP1N4039H1/uZ786VOzvQcjdS7VQisDVAElQkvIYgCYSNW0qQ0
6AjqtRq2Oy7YrwyEKj7Bb5vwD7qV2EsUYGS5QWBYwA7MD9e6rfpcm0nkP66yAE99tfCr37Okxpj8
UQssxrfrAO+OlKC2b2lNJxPVb25W2ouCA24N+7ZdxN38xEA9IFL+OXEVMIJd3XN51Vl203xDycnJ
bXmvhRnkL2MM/1YQAajqUEkZ/W/fM8KUViUZkMHPS7NjODnGa02JtXAIWT5PcBr3RtmxlplCFd6d
4ExVSQmHfIkE53PgDFxcvjYSfTpH1S+M4m9muFMJsUfgWXmBYsn1E5Av9fYTjo62Tia8XJZcYGt5
9cIsSZ//9AjRMJQLKHLp7xHdrwDRKoHL6BAkCHg78YAAOQWZtwCf5qTj6d0iznrvav0GEMTnSRvr
FqZDWZOD8oSLe3LpvxlXhAduC5ya/Xq2ZiuxxtvW33ZIRBa+ZzuuBZcYS1mkCBxq1a/6jV51+a8D
wTswFmtxNy4s6ofwmk987HSTkO8f43hSLPvTG/Ifr0Plc4YTWqbxyWAvIG4m94JzwrD3tBDDVx2m
6xzpjph6/j158HnyvZ5RJI9N/waRbkQEUmmqcVFY2oLE52/EclK34q0zZX32PB7zcDsNt1XRu8Xr
1QEBbc67nW4flCNsSae5qJdZNpaqiYcb+SrgdQ0m9i6TBs8o6ZlKqMkH4NTJWfMcplUFa6ZlFJPB
j9kRrmEMMKE4MfvQMsB2jvu0ZIgO7l1Zm8soheb0r4dnmcaruf6BKq0/taPbYDkBt3gwmv6uVG/e
JT7qXh8B4yZXRYjjZqWiMyKewpavYFQaiCMjGstC/kRcpgBV7L8q/FJCSnfSlb1/K89Ad6GBxo2t
wXyPfiRRHD5/PntoS2jVxtRYyHxAGmIWo5WeQmnMEWJumC1hoddc+HGHxWLmv5ZWO7HxND99somr
p7mi0gueDbbr3jnBRlFRJZX4o7G8njKI+oIVFLoJ5ZYZZVSRR6Ga0uA2TNttBTfxuHSDsJh0CmFk
IcnXAyoP9QZH/WEam4G84w3Xl+D3jdYqeWPSFaekCvA8WCyTWQxBqMlMFJWnsLJvnc0bx753XAlP
LaBXV7y0qSLB4T03pTLmPlkaJf9q414RyZbS4L+6Gu4/L7CE7p5Nuhz/ydY2ghfHvSZcnI0mjf3e
fcz64wi4h7sK4l2F8h6oiAznHRmR5Y+xu5XnCeChk2EoHHLF+1tcArujqRx5Snu+3ngnnl4tZ5v+
o3WOeTlX27ruNuty5fNft7EiHUteuRtoJqpWqbeAXYmcWZXGvd/8+sdMJTX/ldAz9hCt8tBuOWaf
W/ReKiX7M8PsUvZvS2CzIcVdJylSgUXAEOMbIr7+syTrbR7bmnyV+QRXr9pBEzDRTEYVwMoDePzI
69Bm4RhkDa8F8iqRmOml6JDWU6Gl8HxhyrdoBddBF/SrHQJkcn4K5T91zCS+2btfjXzSNImBW7j6
ZNHnuaPySCT20FNRPMrJEj304OT/vQoirKt2B+Y03NzZIMt4oQp9yNZTTtpl/B0H01+YTQpmBmw/
z4WKK0LHF62/nQfKanp0nVwjy5DwGFdz8nsqpapmn3tz+dzYktQUhIIVzr9pX44tQp8XKo4X7Mh0
tVJ58GhsEqexINqXbCdoJDCAod6Nf8abDxvfNg9jUtRecLHnSberOMlVFuG13chUEnovoncmUTn8
v7lAaG+OoLerMlPVjc7OWdaI7KD7N7+Pk5yWfwZvSvqn1MYgX4/6RuwH2ypgaRuZzvqQYyxi3702
UkDvccQxMh7L8WSnqV+eKjvullj25tPY3UpP0uEMeZDndD1Dz76x2WxYY9FBfDPrWCnUgdajUoXc
tVdahVFeEMuTNIus6FYAdaXR/njIotvDGqNoeNKLKirwnEyDPg3+SzQctvX/HCDt0uCzNu9PHbMn
TccR+xWpqtQ61VKGzA5waWLlsxxsoTKaEW4WWFfGKqKBrnhlx+p4t6DdNHSMLI5H0+kWOKB/Uarb
o3YyqhykujZMr2WRiSJ9DU+sK+1NgECu7Ewx1oeZ+4xAq3/nfwBc1ft8OejTrsxk0N3ehosNNRid
RPY6asZnwiOK5vZ3tKOmbWcS0svjAmZzVk9zrkJg4YKx84PqpyXRopCnB+WGj1L9jcPsVb+HBR8/
ShL0oq35tOiv1NiIClMH+CcaKRuaGide3YIUJeaG7e4Jz4XsuiIES7Kh+7n2zXsD6rkOxde7JUYE
u51Q6S4ydvJjDsjduPnZKzsbBXTPw7pSkf23cPTS8uBG+TA45E3SlePucMuKypQPi9ILJvFp6T+p
3aCmBJ4JoePMensxN/gda/Vp+FfnNUvyYoeYWDqMU5dtd32r/FbxmlK2TDfMgLvuPIh9SoieYTyF
Y9euCYVxQdb45QpVYVbaBOoHOZxLWB1XpSEVBrM0PAYwWZlswuoDsY51JI8VN7wbBqo3bCK0qJ13
5JQX/hfhddA3buYbAtJ2nUFsR+96ngMKBRxSA6N0I2YpWBPLYfT6uPcmctLIey1X3YR/ByZtV05a
gkFE3XlWSZbSFCfMFLyw+/l3R5Q8HNPphgx3DlJvKSHQ4sgimy22zJ6h8G37fTLEVyGKYTgYKC7d
04f0hEg0W8e+J2mqMTe56qCIyWSmzALNlw/xhKXY+SWEZZKU+vmkBkdfgs5P7jKXEdtgMM48RQu4
mSEuKV2drPUhlnZGtAT29q2ReVn4ngGQIkvzCQQQoZrjIJ5rDhfTpVn8nTUjDWukBwzQ6g9IcLgj
SwhDEK8VTihj2AuHdjJutD/qG0NSXULOKye25VhjB83yg7CuNsZNLndsSzDUFRpJ+Lii6bdVbH+P
KgnsQ0psV2fCyXGxTe6zFjS0NasuuUoF3gsT0XbYGSYUAR/G2jaPL1UfPwm5S4/pByxd4iJ1LIkQ
oOy9NnfwDCkuzVLYPin25fzkL+5ngy1eRZYRvIJEws2HRsVsjiwL3hiszpXsnNg4cARCX4uc5Z4B
/GPGGaw/bpSUQK9UUycgZJDDl4rkWYZVCYyu2QGfyDO9o4Nz+aZlrb3KUY5BxbeJws77uvLuxmsE
/FQTHg9DuBbVJ9kbY76BkMoukzMlf1hk895Y2vlAFrLiiOt7D+qm/Xd1XfOF4xkzAciwgnXebRxN
8cldcvhZ4mn8mnE9mQLXSlR8wuaW+3M5Dfq8mO+3TfSgTQRuytoE9QcSJWEvoBuQjk2cffB6apo3
z6gGVcqCBmwMCdzInG/HZZAx5QVPzYyLTXhxxRhobmDcPXpJs5zg/AD1KFvsAfZvPWPsm4zpP0HA
NwBUEnmzmk1ZPhBDuVbtpwRNKCzL9T2Lz/acti6uzHvb9qANIBrdClMs/BD1tQV25ZvYrQyiOIHF
Xl0DKmv64H4/OKV+dntRoCFZKLBhtA/HWJnfhE18VDN8Fog6eG6Lr/0zeM+n7VAdmYDc0xEGVs2T
cwm360P9s6sQ4tmG3x6uHMnI3CiZc5AHsjla3ZSCALn0QRZvWTSJM9z62Ll2xvq0JlmWX9/24Qi6
AfGKnjUxZqWQmIEZAWN7WEs3Nh9cEK/IGlw1CKH8qt3Ae1dh448LF+Qid6UwZT7VbZA2+AtWy02q
oOnyBlgMoTjZ/73E0M8Uoz6ifSpO5nFpa/ObEmb8cUfKQSWfR/Ju6t0mbJsl4Tq1SvEZVdc/uxjo
tdvtvx8S6gSTUn/WyLfQpN0OwTkNW01ITE5ORIm4lf0abvj3GQklQvTU6QOHzjfHsOcSSMpjviOT
oHN0uyQA4ZUVBtl37TexkRh2zOEolW1QxH7upBBHoLTSyExT1m1iuUrlpI2XeeqZPDZDLgvgiCi4
OJB47w4MgsUSmZ1fMEj4G0BbPp1cJeHarfIw2vKtw4/lGYAE8RSmKVqgmJE0LT1MkOya8A6qnLJv
PX2hGS47uPp9cRHESHhjOlf+RDC6Thu6qztmPOOlsOgWw43EnwCBOotCOXcSuWNJgY1v8nf01IDb
ALfsP3gc++i2wA/FanKvuBwNKjUK/8+3fbOI24cmo/hyPzxXt8wgqOISV/7JHeO28dEaPDTbhYS3
xojIyb3XdhSG7B2tEdnMK7oW4MfN8rYqAAPjh5/MhR+skQEAJdG7rMKSVatHCRnbapV4EL6cFIoL
JVkdAAKQ+/weOi0ym0g7KZUumXssagSNcMB/cE32G5hO+n/RwT4VegN3w0+h38JrqnRtT2+r+9Yl
RJkypYr4TKfXMQSRL5E1av2ij6UOncSUNhl2bb2V5WDFilPlDpkna4iVPTMdx/XRuF85QMrZru64
NqMAA7sLGkuZeMRlZKj1LEm/gVEdzeGLwdggz5EX7uDCZo6/LLTDMQykLrsMjMDhQOXA3RZiXQqk
3Fibp1YZfFyL7P8ofvS/XRb89T0RIT0FyXxpxohK6VXIbD+HeDOS7WiXqV/t5uKbla7gWIb534q9
Zrffa7rEPxWf6rRXiKgUZpfo9HvRsGUFJkyAH7CFUtlEwKa8NsP27K9Ocy8VgWQJHFnNvGO40diI
0WKuQ5P3ge6Iu8+nQfr3uh3eVCeGbBnEOG8B4q/zkIx47OMTv9yedqie48jICgYbVc81KB0TmOmb
TCvGRauHXzJIKaoQO3ufkGNmg5w9bl8A6hPwu/YbJRN3zWhHS6xIkXw68HK+U5pUchDw62njXLll
Yr32Y0sOYbteAODdX5kDePIdNkfwYmaD3j5iib7nNM4Ik+8/1VkvaeEa6SQ4Z1yUvzllfED5Z0Dj
X0rRAUZG4ZPgCVFoYEHQGX8e82xItzEjJ5jvRthF/kOIYSkEIuOzM86Be/dhBalLMToUw+6ipEAm
tDO6MZT6g3G0MvcGZNaQiNZ6J15MhsELUKwMlvVxp6VUPlfywaJZT4VPa25dAu4FDPGjN6l+/DB/
Vfrpv1wDVReraHf+14Ucu91meW898ac83D9DPA4myAsr7f+3gldLuND7Iskyfo0DpIhPQI0gg1hW
c6fBX8vQjItvnvrz1jpIi1QykIFDbqrJ7Gd61xiDgBlS9Umb+xWK8UlRHkgqmEoReRbCNwArN6uv
mMJr4+PBXybnugO5NXCgBMHB4iZl5f0DNCgLZ5/P01gupsm/2AKJ1ZBiSJeaU3Gh7XLKofCcSmUI
SztwLvcgYbRBRzmVW1eKhPmcSfXaTFf3YVafHqOgbMtcbQWLNWhhM06/PW+T6yuBGrA5rdJDfwmX
OairxnCOs1aCBqCrLw0qm0a+q8ZC4ysGCxWXjyz4S/7/F+2Bh1M/gN8mtA1KVte0/eR7as9jHKsH
svZ/XQKW1E84w37j73SDdIjv1yQbupxTrurjyPeo7xxbr3VZu8s8mb7dgm3nzaaJRzpQrnR8w+ZE
eCzNPXv35XhtWWKHMIufvuu0QU5igF2nstplorXVw55cjz3937qgGqP5F6T5dZg5Izdk7X712BYE
vqgXeqHUeSKSSJmEr0gPmq9taRmb0oIDZp01e/PVbVh9mEhjhmQYK0R/1ZkVwQ+HHYNOxfk3DC7S
euQ3VnbiaXkM9l6Lvg8boyMoFCiU4vW4k0S2zKkDICuHBVsMrULJhBfB4S7yoR8nPhs6TcjPOTnM
DK1q2mXU9UM53OAEVwOXQdjMPHaVXhnm0vw61O2G8Ms+L12Q483Fn0j/zQlpBl85yssuhRXwfXFW
HEjjmr2t8yZwmwQKIYwwm7T0NCZ53z+86aVijXbwKHBQtnMlBSXHu8R6fAkWlsXFJQYtDvluKXBq
uvKlZ2TEJxb/7VOGWcc3j2mlsFaPGXL4+XIlpLfETRW1048AhtHQdEbQxt7bWxbwllVoTWOxV5CR
BBRQKWft114BL3s2adlHnsIyT4NmNuVRnpjEo2RsSLtOEPG6SDONjLvKLhCEMUlT3B80FfLJ/EC3
nNJ+pxyfa/O4McDZO9UHz60hWrRTAG2hkw37PXSkKxaJ9IVdN3XS82Dk6ale/XjX0abBqJ2HbAQv
WWIdCvjZaqx8UEuNxAdGHSxjZNUoe7ahzVVEZSNjhjW9jG5BggMuz48ProeChmULqcBX2Q8jcYsY
DYm9H+7Cbp9bcM3NquBQBzZVraLk+nloZ4rTeNT8TRbH74zLh2VlkIGJrnd+VnUHmfNfAKblVpvL
o7adzyan6rx1oFLq98r92wkoOwjft20dale4wCALQ2d7pwAgoKlClcReOG7ip0t14qk84O41STyY
aqNWd5kDGVwoE9LVCQOym3Ky4pySrlZXZ7QNsK0D2xvkifm7OQMNSncsrSPB9n24g/LVmXtz7527
Um8QP9vcz5F/94dvXxkW97i6H/Hg3xxOaGY2EfdmGp0R7B/qB8TjaHWqzi1SdxBe8q8Vpc813M66
rEuSAmBLFKWPHJ+9DR0o6dDTljn10BJj1i5jPxoTjMuGfj91t/dcya5BOWu0xzXxwPKgAdm0Sj+O
plp5+7hT7pkxnTZjQP6YIu/C72wCxnxpVTG7DtPX9u7DfnzaNODAxMzs2FXSSKVnDB3fHjqTsp1H
1WizKZgl50abDAOwd6KivWWXXJlV4CougvTk+6OFDj5Ch8OzJHAAIxpe4FxdawTbo+ixKjBHibiQ
/1TqLBNmfVI6MtNyoqSxBy5dVzGNP8y51mCG5upxgthRJQzSFpcc5od+1lhwQhjX9f72Dpu557qF
WhrtsWgI0u4lq+Fm2Hr1ycgaABOHPvqwb1/lWGDCfKbWozqlgFZBbN5GbAGnF4goAFUMZPIunVuf
NBegEGVqH/OT7W0DwIlDSS/n4PiyEgfyb+1fKOBtxO+856eRR2XrEe86otIXIKiF5Dr8kfy5f7OJ
6xBPublJhM4Y/2gHsUuuBPD/xyCBL5UfXOE7WaDSo1BeoBk4Q8Eyt2FFC2LkByFkVm8rdvoU3ElB
Qck2s918almWWciRPR/C5YvaNi3n3O2Y0i9X15LDOG2gM881F63BjvYjupnAsRwDPk94npZHsGJB
FEnHfLFzCOviooVC0J7Yz1q+YadmqZJp6RtELDhmYXuCR6Fp+GbwlEDWlvUesQL3nEhTb64FtCHA
cKDTCeiChVzgwe5L+ZbjKFrg53oEZQu5P/46GxNm7JGQDDhj0ZP35tBiQj79qd7rEFFK6RW3NuJ3
mENCuX0MaddJHzS0TMLtg7mXdpjKmqiDnjscPptzbVFbS3i02ARj/cge65i9OBxMKGq/h+R8yjXm
EI1oyo4YqbpBvbuNeE/vIYL72W8AbMls5rFI7lvZ2BpqfDPQ1e2dgPjoz7Uj2SEFEcWh/k2MqrSf
AzKb6KjuDLyv+z6wx1i858LwFVg+F4iWoJ8mq0m0JpyRvuzMoRnEqPJlgnBkOkLfT7p2rNVwETW7
bbsLXDs3R1UPBrU1adjrpFKL8A2r2scR6qq6EOrjSCOrhPLIa6znWdRg1KwrQnBLp1hzeJshGi7l
cjYRAQJSta/cQumfdhDjnBqr6LTvH3Gb4DQ2V9ccq0UwpyJbwbakbxBoYbNPqwjCd1gVXXd0PT9N
ZDpUUCh+Yl0IixReY9rWsV+cFhNWs+UuOGvubk/yMkT99jJWfRI+K/TY2QkZMvnsVi2c4F3lHDQ6
VpvkIFTsGYQza3zs+/5mW1r8y6ebLzQuyc4Q+jPQ+vF1KNBlxCykwsdPXKe7KMtabF5XR3iHchuC
kDWOJhnNYN8TPx5TMSDq27ilonpqe9AlmmZBrkXeLuuz37EezVikLK33KKMSIKJvoCPekiPf8pn6
UDhZJJSwq2AHXWJ+TnpFyBEArp3sXEzoxGHtaGbXTiJ+A5qyFJbPpFfn4zNWF0kqdDmkiZY0TGKL
An9YSnOKooNSQPyY4MWT3g3VMUwnQCmHlUYdUULQlPDoopTTyhHrrb48Q5pFOrI+1MEBdcszjG5E
j/drERjUQkXTpMSKNpb6i55/DFa59k4hbpOlMJ5I54y4JSX1EkWj4XYORQJkW08L9FjdPQ0fK2ww
O3Dk9PF6wIXwaNMPimycdBCyiMFiAREy358f4Q95vm9fR9bRh9qakk+nTdekYQ80MZ/Xr7hTU5Sk
iucx+WVi4Jro3GLu9iE/1QbajbleoRJRAfaX29ceZiD8DW+EGuvtkM4ahhu1NjY1k2JUdMzegMg6
3t6kJVnmY5oUVFr48TbPhoXUotr1ncRJZ7lixopF0LWefYcWPHB/kUBpDCk9nMlCBhSsMPaO2gCA
mZsII4Snnq3S7wCatP7r8i69Xw/eMn3GUQim2ZCxOFBNAGNVKl/SQT4OfL/+GI1WTaseq7Y0K0Dd
E2XBrgJrDPxGsLzFmovsLuXY51zWmUJFDL5u+Wfb3htfAFlJbqIIxmak3yfYj0GW3AKDurUYrIA5
oY943KfPWDO7KA2tA1T/dd8gWpXNGuuujC+ncrqLWiu7dA6owFfvS6RsKXtW1wjNYnjnyAzPYwc6
XEGnA6BrPvWxlgySBPd+85lh9mqvGUY9sN5QIMfpZg8mhkoelZ4QxrBYkz+bjv8hRA9moFQ2KTpb
bzs3D7HQP6m6a92G8xS09ML7XB2Xw9w+JefaA18pRcWF80cvhcEQvSTPlD3+Dv/kvIkXVJk0we6X
HALbJ2r1hD7GRG+yv6b9Og4I5MJGgY8MeQ1uAAi8P9AeZMM5JVzXJPI7EZiySiYSJdMPphDXzhDI
j2rdOnidtCVLhKiNP3I1mti7M1cGoAQD4fEXCh9t8/cZq8qoy7or9Cg73cbMno4cqC06LfbT57zF
mzCZHEp+RsaH/p5NGwBEjxV08se5oMw9JV2J1gP7ktMqSd7JyiqZfeipL94Lx0dLt8HxZtWaIDUj
efc+Ib2VVe6zihm7kmtDsqXRN9mJ9dMd6+vYqYc+G/jSTxjV6zr7HUWJail3c5mxkEUh9VyqjIeR
8j4rwvyyLmvfSC7IsWUS4rQCWvUtpI8cvfbjDs365tzC537GmZ8WYmzVhvCbWHe8LJRL5McNYnZu
+Uokn2MbAxiiAsQgEpZEQFSeMdI/UdPrSQ/BjLicgIrW054MhxBNNS+RK/fl+KcBd9XUi4vnaLLl
yNNClb/gcQ+2Vnurx2YvbITwTl7N5B/hmcnkxQQ9wD4ESzqLpRl+Ucc0YdU11WZF6PTDlS2aysWt
F9g4pJg/+vBY2MiHHDNMlWzE+Rn6Xmkoze5AiTUQ8yei2kwh1eRBwE1Ox50VZEwbxJhQF24Krlaf
uxauK31AmZoO7KSTfP1+y7GHgSBAd3YNVTD4gJcO5rrMA4zIuyR1mDFnGkldtvD++3hKkEM8WKxY
OAanRexe5hhDMlEfI3VZclGyOqfh5jXsKuxQrzoRBwm2CvkdSoI/1O/H2PlHtZQvkwA1E+wMC7uo
3CqgQq3aYDoyBHaGKigH8DGZbG86Wf7+HyYqDU5XKTKs6WCs61Lq1Iujvrs0Fvia4OveDdk4KA0R
9P9FtjUpK+X4qcBoZAt2oQLe3qYmSD69DvgfWEoTfMEtHUZcLFdApmek4jzXOxtEAG/ajzoYNnVp
VY6Rbvat3JJRi5HGtNiFSIsnugnF9B2INQN9H/EDnH4WMhiIT4P1OIauW5GGV64AEXqEeAnDR/t6
CTrqT14g4velGVhfOzgTCNcCd1GGmC2zaCCHomLvAaZcrG1zyMX1jVfrry00GbduFjkndIwUFrIR
/zeiHGMRdbcK7U3ws7R0c/EatUQLbJNNGAiHkDcGJC3YRNB/G35AlxcCCp4ZRU+0AZbAI3eKZ9kY
Z7OGa+8PwXRXjSrEmlAsB3mdQfeY24w1YJDxc/yMErwOSEZDMKVWWwPakHXmHoZR5XprOk5nZNql
kuMrl4AtjT292eD9E8czEbzxZ+4sXmSnfBd6uNLK7Ukn2WyXrPXkM9oF2P6Yxgy5UZJzKdxJzqpx
1RwPsNct7qRFGbRM45rk0eWKSN4BiY6AAh9b/6sFtn5CmCFLeGP1nF8zy22nSG/u3bFEmol3dezG
GVFPKjkmVNRiYQRT/7V/WOpPGOA8PgJfILhjIzeQM+jpMu+cmPhi96yTdCkiEgKGkaM3Jtme9ccf
wqBsbrmg7zPZQT6Lnb/pFfBOBRHAv242yjdKX/qdyKiE3vXv5e5hQE0EvbNRhq5nQzN697ISxY3L
rva+PtskLp6kSgOLcrV65xRRcW1mcYIek4N6iDcdcEKOYjBxjesdtz5nhih/FnxKyClDMUUZgvHO
Q8zs8bzudfCAazzMankppxzK90V/E+zGpCse/HmUk0ZNZGnnaJIv3xxV8Ym3oF+yXUEQS0ufcYkq
ooswadaanalAvOP4+ichK69YtHGMHXLwjVGILS+gS9r1RwWjTg8GzLAzdU5jEnnwveipoWAYJtAK
x5vte+IHATaEK8BJ885cvgpU550ZdNLKqEl+eRxpSuTXvHFQ/FowM16aX2If1SFamHD2LHXGnmRM
dFXp3MlYd5Kn+UKZkUNQsFMD2G2HgHgm9mkcFsoZJrfUgF8rdXQxlYabnRr89IVrd6tC7mQ7HBAo
HWDR7YAalGLrM2hqp1p/DbxNTL6uzkWXNLHD9eYb58bhOwWEJB2DD/iHfuVSGM3aGm9Q7YEueSrv
sUmTC1exa8nWZVuw+U+e8quKP9YuKqQuBiDMnkSfoP3AUg48YUoRUSuLhhnxap3j+T9g5AQGQ60t
kIQQB7weBpJ/4rYb3oA+mFCuRN2C0LXUIcMLDc8PYN8e94Yiq7y9RVrr6mmXrsv1+q5dqScJWAbs
PVvMrWlO9npSdhWpOkGY2axDVpgwATAu9oiRKW4Ay/LN3R8MT3mfnpKztEp5evNrM3hRgTkhyGCS
YjST57m3iMv41K5QQGL8IYyOZ3SYBHA3AAK/UaAJCjRpz6hrFHfo5RoXMs0Ylj15SinlDMvyVbHa
xjY3aQUp8ZuEBu2o5falRsI9j8D1w4lV8+ULNDD8tkmXaemsEWA3xmdUyi0chYrLOKe02ElGR9eZ
VqNa3MEohjAWBiZ5/u1KM+PTbFoIsBPNrovDaykDmJLaCcMnFZmCJoCiVlS8wSUZMJIkHEoR0grp
4AuxOV3vUUmN54u2IqBx0IMX8kVxXYyp7GBc/4fLURd4JU/A/+9C78PYxP6WRVR/4ASca3c2Jpjb
GD2Uo58CdItnvm+VsuP7BMM6pkfa880537dGEdYnch1EAp8Mh7/k9qJZafMOgzJsKbWCQsxs8rbd
kKFa9yx94w9KmO4GFk8FcsNSdRIWJMpfOlksGQ+5Pam3McmgpUwn32YJoCiyrxZxZy5xUzTrUDny
2J3Clz8hdemOlrLu3YRV9Tx53vOK2T9xLyUhWqPQ5ipRzI+xyIr3n1yrz/1EFVpK5sd2yHTRAZ0h
NkHvmeZzdGwGqaS+V9yTKRtJ8b4bcHlD6LigHTqV+bJhKWQbSW6W0DSYo+AcL0Vtjkq3U1ar6Gjw
m+yh/ti8gMMDrl0hCfZI8x82hPT6NqGhXs5mK/qPNs0szA2zuUua1OEMWwRcOoIvDoOSTv8F/UWM
8qlEPWFgqWaiMz3rwi3mMU3U+2igqsqhxh1xfGxj2bW4E9Nav4q/7AO7RuLPCcjYeWF8Wu6gmoZB
50L6G2sBWtp44rDURiqk6ZdEGmIoIwUYDXZrfoTgaHyOPOlHgvlb6aCZeuVUsA0+jf0+5tHsDQM7
rT8r9VGUk2l+oWoqBRoc3L98xIdoGZ+ipXj1N8hJrGz8fVl7TG9UNRLcWZyeCC2xi+ccXpkKwfHQ
ACH6qv0dYdxRwdEb5eRWpdzMAPNUQbIpx0aFtZFxPC0QR/2jC5YQmQcPxZ5T0D0DyibpL5SUgyjz
isazxh/j6VNPwD2YifuIxRy9Nag/TzSBIthGiPFLrdD61HtW8D7XtokpYkP3xHbPWOJMohm8ZfUi
uXi644Y4YhCgdDz5Z67/xY8EB+dWvM8VW1l7xK8io992MefZTscp8QA64kGMcrHg4RpEiAinauVW
ols058bRymSmZFx2ayv9qU6+z8GBUhaPXVtCI6t9JwxbGniBTFp9nxVjnvLH53tIbDTbB6OzI2Nb
2ClJpDuWLJN1OlcJ4T0qjAH8Esa85spFD09Qf4LuC9KA52tV9b63pIL4BFBPfzDNXFwXLL39NdG6
Tm8/WwczksVps3NOaTESkwL+0Fk+HJNY8HwFjlCDEHcxM9ABnP3yZvLFxeGziuhw0Bh6QYd8SrJQ
N1tEPWEiSv4KNFfc1B4MO87leFGL6NnKPilwTqZjXUMbQV0Hw+5CAU5LRujvVnF0pzJw8Fx4b9GF
l7kI7v0n3SSTCN06shcS5e5z6nHJTuRjJBtwYPJ/dCKSTrX3L8YKqtj7sBblpXd5v5vNkpUes/Wr
A/G4NvbtSjxzXxTWD8/o3k313sFTsrj3nKRxvKUAPIe6ay6XTHGM8fpvfkPnQ9U8D/ybxBlEeou4
AqgHDt/Ui5Aa/YB0BZWvWxuCB6twreI/8AHYQwzYsimSgYEGZdBQfy7/AWgDEI2/DmGWNcrBlQZQ
BbB9cJGb03Hcxmml1xAAeUTMX3gg/+tbIxDludxdJdKgR7MFwpnwJO2bSZQGbE44uoyAZb3D+9HD
o3LgK4iGgkjcfoUkry4s3unNkc8snb9RL4WhVjvQtW/q1VLFOb2O9YdNK2TXQpBTyPixaGSpxKB9
Y9ouWrRLW4qRxrQWwWSfEvWVF2lCG3QM5u226pcr49urwWH/ktbNhcd8+2F346JoqJ8htt4TFtVC
D6Pdmnxoxij2QX54WONNAtwqLPUmofJ0ALcJp7MBhanoIMsag8VcLTr1+55vv/ARQLKAkge7WRul
18/RoJYBrKyhTJE494N4jOk7EEEf12YDkkGENEoVMmwXOfYohMTBHz86yQteIH3FSFaWGzJcESYh
qmdHlaj+OBay3IFGXf7h1+UuL1LfuW2B+I6mLYi7gdamJF++mZOCwVQeLc8BXT1YTo8E+NvOpFkr
opmpNrUbt1E6bD+EUqaekoITw3FAKJ5RB9NBNt/+4uDi5Fmu7aKSEtjgp19lWly2h/X/Yrs8ODJa
34zujiCMthAx0u2A4AWXBulPZhCS/3F+XWh8AQppHge51RoeFQanxL3KWPAKH8BKQXdvI2zJ/Gzx
aWe6IVpOIp9P1saShpi9LqyaQy+CrWHVOtkO16nNNSkFVdP+xpZGnvyPJ44felrTGIEaNAEi0Gbm
vVNhouaz8hnHU36M3prcbkT9dCXkBjqRIlVe64zkBVupP5j36lsIoM/EqSML++QLETlvs9gaPYGx
5i5KO7HnEHP9oHeXYV0P7cPnTNiXC2GUlI7bnBf3FNjstPfWmVptCClDFQh69C/GJqfcUw0j3KyW
LeRKqqtaYbYXo0NmQBd2PxhZAoI+Ea0eVXbW1Y5ieo/wR7E2I7GZ76sK3SZHC5A+71xAwnAhCc1p
SRw2QENtUi9+MIv/vZRadjmlf/TtebSTbgN/K4BFi8Kp+MxrPLZQbjFn6xwkmoECvLuZZmSPEjdp
ff4kI3txdn8bOY6XzKA4fhl7lYDDVi6pZlgM+qV6bvJGmsiqUNZt6oWDL6r/yJ5IxoXArY2w5LMf
CPzFkUMSJ6d+UoysOzDnBGpz269Tcn+gb2BaLh4gwGhUqUyKsiCri3SrRu/P9xISomStBlLvRLd3
iAosb9C7YNP5taiPVJTO3PiWIgy7p5u0Ak1vo3TzsyaasP2ldOAolDRiF6o9r+f6OHsXQN4XuEgf
wuhe18Fh6sHS+7wZyT/ucF8lbDV0LBFbiQ7D/JXIyGx4p6PxayGkz7zMx5WriwmiqSdDrbbTQmTX
MzbcOsauY787Wuu03JL64AGA7tm0sN00g3dEPAGhGq8CtOi76AQ6N7Ln/VQzU5zQU9GCdrJSUOGz
9FbJaFg3o4RwJc486LD27DmJSchdLaLOLURWJSDbijQMTQL4fEdR3bChmki+z+lHXBSF/bXOeymZ
LV+O4aNyIToxZ9BN6y42ipmHQ7nGkAr8G1NEYzitthWWa/o4gc1TJXNyDLn1mTkcS4Xdv/xUsCmg
6AkliCXRGCNbsbV4eFY0efgTRGZs+nhpjjtibiDVd3BzjYxkrylMkoCTjJOjJEeQ0ASFvGGCdhcz
4dPQ3apiR0Zjc8TRmx4qUAeO7m83wOiWZdR4sSeJILJkgxnzveQgWFDBH7ibokBWl0TFkMUNrHpo
eZTKlZaIl9yT8uS02nNvFvKwW0HqLQIQuZd4vtjEK63mALso6kgXdZjyPK9cyNEbTyCTMssv9fca
h2RMgGl3ERkE4xNFkgvMvCyr7zn5NIVlYRieW1BR8uATRqig1mVmgfbd71l1808HbnFwAUgoK1Ns
8e3JMQtL0FFnRxeP+UJyDJ/IyOB5GVk4XKtaca9LEDH8EfsUux6+a4m4IRZltx/8vcxgO1/zQbg1
xVvcXiXvtxpfh3hYBwaIlRhqpUbrcf19Fmyuvh2xhsx5eNDSWhXFflebyLsNgwTtzgno7ObL/2Yt
ga01n62oFmlsKTZahgpyzLd7rMfiDV4nfEqPtKT4Le8OYDv8UgzWbsgFWvDGQ7bE1Hxox/Z+FSxk
43HJLDihlkwYUEJhnm1pQbkHUn/rOhQUU+KD1sP/v7CTTuonxuhfR/Rebac5+QsQStGs9wUSh6JP
5N8zS/VfDAQkBSBQoUIkpN/qndYlXFmSEGmnpxwq7lAM+Nt8mRRueLi1fApfF3A+lCwTlojUr4Kv
9H1b1Ig793GTgLG4JKhCZ4oKM2v8jKUQl749P+ukvRH90mJ7wRCaAm98pHzqXxnWv0AmhdE5AUVx
IMo12KCG3fIqbwqDu8GMn/sASy1gJ+YOhsthCVhCt5xsrjd9eX0KMhzrP3c+WMyoX0cW/IZyMDHW
e1j5NVfddnOPuzp5BOoedsmdm7d9gIqT0w6rAXpM8XnsdRfj+9YyAm3vL2MyXL4MC6BJORAnTB0S
NLQjnBThe+WIDctf/cLrKctqvdXyb4qvH4jezMtd3sNU0271K4A17pMdmYRfg+G1vZLd696ECGSI
v1beu2akG6PYl8a1NP6mf5th/sdPvYAP3dHrv00+1qN3s/S3E9d/OAbcbsIhqznNdauDdSYWKEAz
tAh9cMYQha8B3qsnVwxP4pKvCkhxKaidLS6QlY1I3vACN6mWBA8HHnGjnzG7FPciJEWHR56w6UGK
tUzktPY77SaP8iFfDusOt8m/4gS3arf4ApGLeLmYnZ8s4HUHngF1LKR3WfmnO8q+4NWs+n3ri/wk
w6vGq8WZT8icb97wsuk2nNkdEduVKOcEh9BwrtXFe1cMFIA9tSba7FjkvQkIWulIQZGocTchbGHy
kntTwFVdfDxOtzYaOwju7U7p0zvBZXVSvS/u3poprk8q1Ax55r4vnu1hpbSaseaGT3r+ESxsrVCX
uYQ3oDk1i6uGGXPEBOw5GEcN0+cOdQXGDj75iH3ntM9nS3s+8ppNdww+/+fRX2k3JQg725WrDPdf
1TTtU3zO3952Np3O4smlaoFUPgELXof6ffsG/CPSqpVQTtEaPKfJ+i3urZy/obBX0l+W9pWr/0QP
DUmOOZja9Du9BHaa+8Bl/6tuoVua8xnQxQRYwY2Rm37yNcV2luTRmry1aT23BpbNvRz6byQEUKUc
00VXd9Jw2mKQp2WbFdlPLesCYjPffwsCaODbw6Wd8xc4s5NLJH38hQF3QUqD7mhoB3Ji/45/Az4q
lul24Ya3CS0fuklm+PP/z6lklor/EHG/KT9rpWyzwHXbDbuDaNSJxHXLeQogA/DOCbs9j6N0PbbK
i/wYPlP29Fr7kiZ/iCC0Z5cIvY6RXtuwOqj3DA7lSM+SUBUeSNmKkssLPh6u0Oj6uVbsk2+ZBDMq
dNN5CekWm2dDCXZmeo/FBB4k5dNx64MeRO/XnLcIX2XidX6cUID6PBkasSM/8fmCXvwZQK1oS7I7
J6MlE7jbacqmPkxU83rqclE0Z5FLWxQn0HSjem9f+BB+Gkv8utZXI+JqjEdmSVK9xet2iZA+COEJ
uUp3l4xtGt8v4DziLCNDKq/v/+1art56umP+LQL/F+ek2gojJlPYmivGONASplGwhu7ipkxLO6tF
kCqxhD2xYOnfeHsgMHQau9LQhzwahEddqn5mGWTm+pye163lCJw1SJGGH7JEANAgkQUKnBODuXCt
GFBkQ5jwaTCL7EQ24O5NEpz5wXWWtFU4HG+FE6pXfZi72gmuweQq+NPqumVLpBvmUFYdBpuUQ54x
482F15RmTGMGI47QZ/da3XZu24V8XV5AvIz7pGRiTZMUe1fipA/p5VpHUbDMvMkxWCJfe1n066Zv
LWefjdwZG79tnfQGaTABq8WHreOZzpt2xyV1x0hhgRSfGsiW5FLZVnwkeKMHIskzoU/oUghHfwPy
3hmAF69rkWZSrn9Qj/zHUFlMOS90sWJvVvTesAlM/c4gwoihpLn1YdQpeMjViBK8xlRDa8smti61
xPr4xSy+3GCRS+YwXWJ5K91H/29qDesbxg+WDvTj8TMUkny3OTR+pypY+AfWJ/2twEaJTI7U4s+z
Oq9NdyZKOt62cfN0ysq6VtPxrF9AEtVtaiOxxRrSteAOKBISJHE6pgFfpbV9a6WqzFEXeTKngJMd
ghFRGori2crsdhQjaKUQSDMNZbDp9myAU/pRK1EPsH3F8U8vCsS8Bil04GBXq7KlnP29HwhHBpEx
DhRtht8ctRVKnbvYN8lIiiBXIEL9ylJ3kTFBZQvuyDbKA7RdKQuiQlR+ElJSe4TDW7M9js1EOAZy
7sX+VMOJRHn6X65lOZXAyaWemUhxzxdPH4VDKT/QLlOj4hLh20HRRkOO+xIkFU/DrM+LQQcIGMhv
RRtCxzAeqQDpBfMv/KRx0V6cJd841lRBDyMdaZ5GShKvbG5bkQzSNh53Uiq2yYYTScP1h+ROpMjk
olMOlzRHmm0zSHVqzjIojUy2/q3DMV3TvhZUGc1hI1ZvQgKUD28vfNeA0ThjlR/TQqxS/WAHl9HN
VGP1T7sfpU6N6xHxPAd1aN4zEwdtn/8W/tFTVvCDso9PDLMMCIsPDGR8e3lVY3Qs6e/jJSuzbXBq
YOMM/6H5iZinba3I/yXIZEb4OreXV5D7rxP3QYJuT2BFaXg8QqocMCUFj4ierS+S29C77oYn6ixR
GefyYDDjN7neYWHK+RAY+yVW6pOo1NhhXai2v5ot/txiKKSbYIhkSMHgFjZLLgyLTMmjcVM504EC
eYPr4lUvzEtWMGqVYImP61C867YknD9L2GU94Xsy+i7fU+zGuDhpgkX9t2I7IuXWQvkUgQ5+k7y7
es+aFO3fW63ti4iyA67p9UnfftDW7dvlIx5yyWWS3VAkdqkmINY7i+mh0s5adnOkBdX1NWWhGQHW
wZRqT5+Rqtg151OXnSKKEbyHc8jg8gC1JaWTm/7osp69aGh/27EJU8yd78860QKkVis6emPytZzm
USDh154AE9Se3lrQYbcsuGDY1SfB0+FPUuzuAaW45DcbQoQcXz4QHDz2XM0VnP4fuImbnS1iW4iY
vPJz4aJ0I+NyyGbJQ+XUgkEW2KRoNgieRNPhUeGHrKDBwVGGaZ/juU4yOATyfq1kaWNqU1dZR5fs
P9C5tHvVXACeQfyRBrgAxVqleA4KuONvK++8k0KRAUom2MHP6UZF435HxvYv4uXIb4zHoROE/f5E
SRDVzhu5e5OjNeG29ZPnugQW8hFg3NrSi2NE1KvKaTIwn98S78hWJbrxgcYj+HvbRhmrvFh8sEk5
l+toETnKJclPgYViIVGCsZoHW6amlnc5MVkxjJdLF1eZpGsopkle0TMAC/Udlasne2ioH7+iW36B
S2cKTyAvkUYAhZD3Ec5f1cpGLZFeSl31OTDbhN3S66ppMYpzM5r11pmZn1OR7a9eyETgzKXP96Yj
x+3W+3b9QrPk9OClBOsCMPcpKlGJ98hhFKwOZub6cpnF4R1aGw4fyMd2G6blHRTdV/e0Occ86L/O
dU0DcD/ZAhjQhazuRop2R8YeDnlRnpxgG0izAHXCAZjKEsvDSzNhPrnR9DAmJ4VDCMMG70GUcpxh
Smb/F4PRfTZ50+kWvkCB4Sc6FE11tlf4Xqnype3FjH+GJjX4hWJsguo343y5iyJQxPUsxOQrIdmH
L+P0DZEiDWRPRrlpYrsJKp4xL9JpvZhRhkRs2PP7oBcZV95i4R26/7cY0/9V7pGHyOs3quWouXYo
9+y7DgxXlqHGLDDK3zCT7SOMGfePIKVIqJwamOUCQaIG+PFYdeEsNE5a20Lfj7zfCro8coVaABKQ
2g1GJs1VhelhVMOOADZ28KrsfTajhJJ/WBvAtxl8Eyaul6TzECXT1Q/tj74OdlJkeM2MeqmRrhxV
WC2kO+YCtXAVOBFZMArMJ+EGxIsTBk8qNQT5y05flqgZdv20hpGTu/621thpKJofbQ3+7HY0FFY5
4evfwAzIzzSlHirdjvE+fIyZzBJ2ouvNoeguCI++u0xd8OjPG2lai3ozQTC2/Urt/+3jy9wFiSUa
uaAUqdy06YQQwj0UHI5KOip62KwlXwu1N+hIdGrk/A83TQSxA3D1RKwrLWPbCkaOmBB7wtABLqur
ylUbO5C4a18g8dkq2W3ylFm9q0CtJebvKrveZu3hFWbKUgJPP5++pt2AUu6X2j2nRQND3kxITdN0
upinTSkJOfYPNMLjS1qDe68e2CQFx3MndQb005IqbEcemtr40uqwY1Z+FqY4g8Jm9ArT61zoo9rV
lEWK2pN1ISZL+lW00EBDoOshAfDOErqJtL8p+2MwFaW4fbDZ6Zv0e2GOij6jYlEuaELEnGmwuxRr
56/Vkz78Yq2hQkFr5cjY8IusggIq9fzkkmUGsBiHOONBvVMklREww5DYAhsbqiG7IrgDF/CdouBJ
hQsJklZf9dj+n5Qb0Hi5zy1PsGYI1++TKEFwxWdJyQ4aAaUgwWx57bX0Vvizoh6YlnlvlIM6zvrz
2rCmTR7wQM4FKep+satJnGsck7uQYOAazkiGHNQwL1CLEe1aqKSE3vU38MxtU2y4+MzOLW9j/TZB
Tpz2suWgPTqXv3jzWLb4VafxATHX5O/al0emTSxaUQS75X2ej64y13IQc7fyzqVc+qYj1qTWytJt
FRFpZmdVPDPUDYUFf0LxfHJAZ9eVcexSxSOjEtw99nmnHxK+zT+03J2Xvl1M4PD54El17skqUdIX
W+8bthUEhlSjNYIbBiEPo/c3P/h3bJakX9F+fPEt54N01OYPS12Pl3unEVAcRzeMDdSEbAdnzLq5
cQvqGvXHE/hHmGLZ9q1mfho1leNSBw3RgH3Z2Ujmr7vPu6uXy3hwir4p0lxVBH+/P+rxKkxTYKUY
Ooy/c70gDG3FEsTFO6Kr+GJsQ6ONyW+IGQuOHi9uLGSATjuIw/KbMeI6i4RQorBRbGA92SRGHbqI
S/x8jRmt15OZeNZ2Sq3rd/mQP48feZtCKZjeQYPSgVoQo4WgDxU3QHsnf7MUT9kpYzHLjNHeKq1t
rQLbuAul0Ysj+iTfeTW1pr6Kkq5hrLxBEJ6KCtscD/+vAL1EhL7j1UUj/JPVRu9/kujtIxAFeu3n
as/D9/Z77ql9/Loogo3+tPb6RD0tAri1BeM2gfWMmubNCBflHwzEu96HS/O4+D71oDOrrFCjKM4B
VPMLYQUB6IVYZlJ04h89DiNG0HgmBqNqHoYiHlUdRvfgPK2VlqabW2aUv3EoMjtw5Xc8rpYxTaZQ
Yz3msV9hDey9WFUUuJNnvaYI6GrWouMRmx/WOqfW0samC8F6b7lAxZAtdbvyqrE79ajit8lVhV6d
Uof1YVj65XQ/MFhLaa80J7vs1pWX75W3b4DJk07U8pa5U+36UyON4PDinQ8/7l9rCD3eWtRxB2dN
FNqj1DoSM4NQRE6/DrnjEMsaMZp1qnjOCTUi0y3wRoHq42tswN9XABeHrDYe5PmIgR4TJcQnOPQZ
cfhsjvsiiH9V/4kCL2lF2jAw5hjOQZl/eUj7mKZzeYUKDAiIz4ADtK0DHfXOOmrK9aqU6jrK5vPM
2N6KIkxMpWVfS7Z3SkNsfNMfh2ums5tUL5Dy7uBvhK5N/IM6Tt05ywpxe8ocWN0OixKQVVy2qS4w
y5cV1RaUh4h3BMhqD3g6v9Jii2/M1p6kd4jMIGgcALjr/ZTTKzbHhFn4dv0AlaqOcFyZFM8UPPc1
ssJQWq0FiFmbQjA5bheexQLdXHSHn0ZmYGSJiCFvlaNOdCUrbpng0uIUUY+FSzAAR9I1qmuxoOzy
DoBKBYJQRCckUq2DrCbZ7OyHNdWqtDpRmxBJn/a0kIHW5Q5Z6wvFEGt4q8J5zkKRCVzPkywh/dWe
j8B1siw7+GD5qjun5nYK57Ss2XVxtPmLxe0w6HylcduLcKT9ii0BEI+pT18JTarzPK//x2Xzp99c
ZDq2lKGTzHr26fsPcxBYLTarzpaGs0iiN7HiOrfkgZAjA3q0CXtmbmEVDhbuz3Rwr+MklMn0B/nk
jQCtli9C32S1slDB33cbQ/W8DV791YPinGVsTpFX6c+R+qkm4QfA5ThPDOtRwokOYUwd5TiHl0Yy
idPwxFAEPgrE2jPc0HkFYExSt0T0J52+ICt2+znEY5Q8d2GA/o6N4FLDMLZylpc9DOyLDyMXZoA8
yhL6OEiUNSL+008vjrHEtX5Il38Zn/T1kbyPH+Bv1oMChvejzQn/6sKf+yzoEb9aVEsy0IOpM/OY
YSZYgFtCjSHad32j1H9LKSzeljPiQralBa+0gx0QefhsRWc7A08Z46mhmvi2Z27dp20iu5erT2Ya
qTpBPkWwZjs/1TN52aeIdWWWuhqkcFjNsLMIFbooNwYh2NGCU681BWrGAm/KHh01uaCBk0Hwiu/X
lPlx/ZBrk77NwugEnTbuwtDKmcWcJpe8M/d9PQOY3JwV4G8zd3P0jfKSUUGJZU1SAWY+uzUG2F8A
shXHbjE/dESfV5pho8+7WOm/f1S434SdvVY62SDIQVVRrgrmp6/LAo1GBFV9FmSEKWfhDDNhoOIV
DDoicJ3XmZn4+YSs6vPo/rlm4fy4602clSLrNSo6dNsLrGNNaEj4vIrCMVeK+B4+WSWo1FOe14CZ
+w+QSnviJtzuyHh9lZ3zzrUVT5oq12vQPQDy0Br9lxNcfUqGSx285pxgtk5DfLGGdy7vAMdHYIlp
iN9Io8MlTgqidSm8C+6ZEeOoAB2dRBP6vyOBGNl15jzFFujziP945P+BQuFN3hJL1lU9YIkWWPVA
/GnGb7RzMg3WDqGveQ2lecDJEspx2Wkz4v2DWUZTvqQ5NBm38lkRfqqLEnrGEjP7b1EcFcrJLBMr
qm3y/xWls/scCzT2iW31mwq5bKD4hFj0OO155VTYeeeiThw/2jeb9CF0uSeHmY9Uzvgo9a45cQ+W
YloX+4CfyL3fXxI5Kmv7NSqpsuXGDf2MdvDsxGSvTrJQ2PEzvAsQEcccQyqQc+QKoPH/sX8LqqEM
7rBj3D2CZOi+NWrU8pjcDEriXegPjkvaDIo0USUsfu9TjsUfEXlxh8zaT3R2g0qvTnARw6jT84UJ
+DWMTCM03gYeLGWsusEfC4K5247Ng/+STt7OWsY5h9eiUi6v7P0fV6p8Itieni05+BixUqP1qg3P
WkhFPAyRqfGJ2xYVqkt0BybPUJTBwXjMcX+aAWCpejZqp9iIqwExC3VTSCz3Spw5bFvYYvu3jWqO
bibdSBGHhQs5Zx2+sCVTviRXtz1GhAq/P/NIk+fa/rc5EI4F2pSn9sqWBoknXXX4rC5l1CAWahK0
yH0hsUaXbIUrPkMVfqu3YAzrxORFse0Q/wH2q1phi7NGKpN2oYNZa0l9BCIpG5ANcJyPhV8MiHAx
P68Z/PvftSq961gfTcfBaAo8bgb3s7No7zbwxN2TAStpr5AynYmE0MgttQu0r0B2Tw8GPY12Cl/+
qyhb+CNRa8AU9I3Ebqqzz/duMAhbLDw63/cGAnE+SV39fQ3kTTI7V8l4s8xZ5IfeEK20KF+z69s2
0vY5TFCjljArXPLx5cII795h55l33ywU5jRNBFT7gyfJx9UxfA+sp1FkKXlUGFwf3pYiW2C5ecaq
chzY+fc1dLwRB8L7hV6b/DP9o8zxx8Zy+mztlE8AHPAup5wTanQXof+s3wbBS+Z5OFVWkA6I67Mj
sOWC870hLfos2Sa3AzS35iAW4CIlOwo0j25CqiT/tAa52tkdhAUc1daAWkW4CCCihV5zFteXtgAT
JEOC17NYPV3kdDnWkY/MSKizToZf6U4I4uuhrix687m2u89nXiuGf5t7w7A3ZyacHO/z8CUoFXGm
JSEH6KnyXjNhRdyT/yvslkRPXPL6iD5oudWG5l1PT/nPHp1xgQ69ZQHjypopUXXm5RHHyDctLvBH
X6zdJYsqX0a4ELEvitQjAR/t0aHyNzbLcfsoHRngJTtD7PB5aG8oSFZ1Dtuk5Q06BkhBDwn9UWgq
XjBw6Ydn+GXgV+hR1/1j2L311r3pRKCzIPpukr6EUR/frHmYNRX+yqK2URi198P33VIMEjYNYt4u
WLFmVvw/ijoi/k/sOXigkz35NAwNwWqhCoOXaZaCElIMRj+Zo9PiWV2LxMc7an8l7VE9GNqkQYE8
c2STaJe8tq+eh+5gFFECG5F2MAx1JsucQtfFQV1D+YGjIZtIQst25wAdVYZbM0se08+Lew3FhW5s
WP0j9DKAs+yR4ChFM1Rv2ZVYNeDCTzR/NbngL9QRKrV8zptXCo78CsJMaCxF3zEPp+exTu5HA6tg
+ngDgsYeVOsVdhWlvqb4jKIVgt/JYyA84jbP8bYT2fhHbsQKF1jZii9JmTVJ7N/byb9WidRT76ef
RR0yIXSA5yp5j5WBK6RtAAfG/vSpQtWWWYb8PFZdWuay9vEgK9f6pzeBc/vxMrA8VcWjQKLSeu46
NgjqXz1ZLdl0anACDjEMDfgaOmX6w1o4cFaVAMVzZMPca1omkhEq/YHC3snL40i0DwUD0lkA7x5T
jQFechSdaDI7EBDFRRpGxb+PU50MVDX5ybcs9CHeP0SukAh/IciskWm3Fj3u+GEp/ylwgpHcbNA/
qEntHce5GtTilcq4p3E/h2OqOsJGPMCU/V96hSvg+bQFv2C1D4whIfwrzE7bjw5NJt3DsqthuPiT
jFnSaOeo6DANXoIDJvHrrDFNChI3jyWU4VbhFGl3OK9BtT8MSbNarzZMPKKHaFHBIJ21MvwU7e7Z
3VdOcAaugmVO2MDCmqCjToCPQ0nvUHXO113DQpIfuWm0De8vBz9JA9L5+LzQrPJyw7JzZBY0b2hU
eI/6gscTZYnNxxcpgReDW7St5aoBkHzgeoZ6TkyL6JIiLG4JP5Yv4CDM28krtCkNuRj2ngR/xchJ
4R5x5s+/gua+KBVghxMz42dKULDR0qZ/zPcfq0tXRFW/sWcEO9/hpw5V2B1NJESpaza7VDYKTki+
3xL5znt8qWyzFt5bNkkDRTGFpJyR/nnkRxx5ACbojYGqi3dBkJ6ADFDGYKfpg1thQM6e4SJB8Nvm
GSlDBRAxmSA4o7gMF3psD4QgIPeJHKi5NEZIvHcymferBjms7EkTocXcSOoNTfNzR41U2F/70wrP
75CBKhziHum3jq154W0S2F99TdeIS9qYM0oC9CtQ/+dzHLKnhbqrpXZ7f+jRWMhfr9I4p5ej3Z5S
s7hezA30X9v3JS115BF2SE0CRN0Zo6Jzmk9+xmLw+bnxmq0IFnVor7nqXZ6ztp6XkqpWfmoCuUV0
WIgWaWpiO4iqF+SlRa/0UnCYO8pzXgfmean4DxRE5TCMg0BThyVTh0ea9hCQfaq3YPk4+cvaxsJq
5DG/yQ5GZMETl8XXvvbYYq5hCjK8pBlhHYdSzSPho9wYnzapFtzWSIkd9K37lLM2ghgmO45KEnNm
/moOD1wB6AYdSiMjlZk27nRiiBTQ74gznYESoU+KYcQAgu47qWprmiY6SyJVVMNw2vUlUNRgthRN
yBvD6uDVCT1hIUyD0a7eDBm8vRsuyrfSyvI/eop++TELDTrnA4kV4R9kSXOkv+DqPvrhH9fM3yX4
30VnD5GnNX/mJWV8g6AF7fweiAz0dBGUUg1Osl0HvDx0pWVjWToBXyB2ns/3iTMyaGL5+J+ufsZF
YoGMa7i8eoeKenVB0QwFDbddp8utKzI34eimS0BoRTzk6uzvFYXMRLRYjTgP2GdULBIWRX5amcOc
jSfHv9EvY+WbIUUfOPfkAPGmSUJV+uL3F2oCZkg5fuuZ8eXi28dZBGoyOOarKCMM4h/EsINai3dU
EjNvZ41z4pIufL74ak1TbIj5SH1l25I4y2WWSIuIgmhnoBjuFB4MMk6oqkFcA2lPn7F8x+KtLfxt
y8EHebCgYlwa/lpI7KpgvyOFRhieLfG8LBUG6ITXCCH/29ygKeuSzmff0KrDu3iCtMuw9ai4tUw7
jjtW23Hvx2J9L9ak/NEoxS/Eq5KrJBpZ8wU9hszqzYOlhddokZcIgIGDH/4dfU+Qlek9tmlSG11j
duCC25479lxRi4LoOK8W1xo0xk06p+4MFCfTbEn/sQTDG365/yiuNYjA1TXLSuJMh2XYl2XR4hL4
dEP5A0LXLFPg2bkKUJcaihIU3cHC/q4Pg0ZRnVSdjcvlYQdXXzyHZUF5oKJ+Rq/4AYtl0dKTxh6d
K6y2/9ebWHhkN569fAdhZD3wZSkf7KAQhNsUPt762IsLoK1ypTVK7zGvh3pjmVoCrMFw81fY+rhg
NabShNMdUspShpfV12Y0fGKomYdYiyGyjdQqkYDdajG7BQ5BTixQZtqOt0VIyht+fCEEh63Z2ZEX
IfWAcqcqAzqf59ZvTIhTPzzg3PLreqjZVkAP3QW48AJUjfucZA2VA2nHrowAmGVW8P3caZkJmjun
5DTJX2nRalciW0ZZJ1k1BVt0Pog8FMX5mxHuEkV4Q6ANQGOz1wK7xb93ZIrLxooX26ZRnQnYCZ2Y
orizqouO4f2Ka2g8/12mZFya4Lzk63CpxzlZ6yJobfnC6dTq1UdHoBpsmGY4/QgS4KhSdR1dkguO
CK7UqlT4nQaAQNy3drqgEntUtKCQwtxpb44mxZuhqnkQFtQvYica5av0ZLp/4LhjpvCeEO76y9P/
BifOBYbheOrUOLq8kl6xBvzcOBc2klGQY+CDLDgmelBu5Cr9aYvNBRUnqV3fYQdvSfKa9MrKZa+B
bIN43f+pkTz3FskcFAR4nUn68K0wevViaN6wGA9uolguiI+lWNeI/G1tqZ0fpe7jcFangFNTb1Yl
9kCjmIVgsx9QM+PB2IPb4Pmbq69CPam+UQe1t5Yb+dAPpP8jyDkElLeOKtiVRI7k4IetFWwqFf5H
z2H/BecPVApaJ9WbqBVd9Og7MMQ+hHs0D5sS6Dm89dkqsvDy7rztYAoJM//ceDyk5ehH5ZulCIeP
XpNzAlq83o4tvGqO56Z2DLemzlXXFMJZ/SilOZlDMyiPp10rSvsDjqUweyR4o0ZRuFTofLF0AIdF
uE7ODn3LLPUx07Mc+OYn/+6q5MkHjuLf0FoXjvrnBoZFr3gl5R4u8gH5YzeYXvU0zamkvlP2VXWD
5TahAYUkog/DMWT0Ows+kcBYlM56r4ST6dtBPN8alVjmDWaJ8DUpP5anRwNa8sJsz6AdwndDzmQi
Hjm8oxQYS216j3yUVmTKb2eMESxzHP/vU7Ldo8SArimbzPLZqBXvrZtlxK9m3KhCymsKfjRIJMjR
I2HyAbmieqqVZ/410ihMmhEw7uzCThYF4HddEMzRFCrREMg9ioWCiuZVR4xLNF0gQl8c8TEGF2MX
apaWDBcqt+dfk8yhv4f2mj62mvgrhPh7sT7UXeAZYI1W11pPmC9ZIPxPrHqMBIvhnokHqaC3Cjgu
hLGjnYaAONZ10TWEncmdI+jB2TRnYbzDHQTEKpQxhlkZWm5oMlBH241fcfQraLOPEhHGF2/LOgd/
r0BWV43rifdnK35AjewhecjCTOboEwL9C8N7auxvdSk4JwJSjYV7UqHZY1g5zmdKiVNKWb+Vl+x6
nWqRhKPDyihJ8SHakGVryXWQKiJolnoqj1SH6BDcYhzk2joxLWOsiMQhvXkzJk6Y7Ei5VoYPcA8K
zFdQHzEmbMMapzpnt1RVsr3BfrjEKMrSH5nbCtRQUzZexfSqP6KLbrB1VYmu/eQw0GiYQKFNBxTV
4/AEP8FzVfkVTbPfFFwLVJq3XWEw4GC1bMBfJVoRl+qh1mK5+kl5304OFacJiJn4J56y4cO9rSm6
nRt/Q/rOLy0rIN6xqjGq+ovJrqcdWtS9vBmZ29tYJPJp/FTJ2KqJYN96n7JvSpMe7N1qEIGxK9g0
MNl/HsenSZK6MW6RqnMVrGryk0o3BdbNG2y7wJ8EwjVxmaGBF5NOUeNi9HO4vqzSJQgVuf6dsS5k
uhu+PebP+cD5b23N2/6AUEtVTpnJ5eaiZfBJjA+injCgfSlOM/qVZ4GluU7tJop7AAaHPeKXozFe
EX/YULLgh7si4ziryiEcPNgSjyMIWB3Jd7wgMojunvk0VsVMwdE5tygdZ/rzba7b6cdzXgKYWe00
QLbP4aaxrGNXx5jLWQnQXi0vQ/y9bfvqlhO0YyqxzaV16USeR3ADxqu5cusC37hrD3fAZXST7Lkb
uy1K6XI1rC1lbkYACWANqkavXxBkJTFxUpG0vDJVMz7wOBFwFYYL8hBOhkYM/f5nQwCJ8ZMKRni8
9d/e1E4izojab20GK+DUrH03P5Gp91HVcdEKGtU9OMopk51dd1Nn8SoFwwnfB1isXZMEB0fpdzcn
CFkx0Fkb0/PDHG/DUnWBWw8TkEcRs9bBzjhEL6D0Yy2OveAMfciV2aEa6NsnGVeNE4e23ekwM09U
cNv6sxucmgzLr00mQ3kJnZiSa0LMXp/Aq0lKSwYXh8MoEXB2llB2kMiijOc48AhEcSzQrKMpW2aE
wJF5LXj/xWcgSgi8DapzZVABAEZSh5Q7rS9AzboyQkipjW5J121nof/z6FTH+KHFM2tshuncXAnw
XkOxw9u4owu3KZKhzFRaQE3dDlTUIyFeHcmpTbf7GBen1GyYxgKaGY9YabTLN2G3scDF25he7Brc
MnrkV0s1e/F962iD3J4M8fXxiNedUjwv7tPLxhkS6PD1ePoKJLde/x0+z5Ql8/EYkvps6A8F9a0e
hcVlQW8jSBXAuadwhAOsbH8i7skPHoDYfrYQMaNZzfubQqrurlLCIpn56DPKTc31KU0x2gXqUDGq
6b7BYNuPw5LwlBr/XlVV1m94RqYG5tYV7ShmUcq3SDhQIbIPezUMJb1BAzIr+fUlDBFFMmcvNJ5z
FWylm26/SkqCawu+txgbmLcbDb0stLnVUmdbrGhox20QhTtPvhLwScGMxRAQCh06CiG+LsL3m7Ne
UMAF7p5v4XRpxvs46rxtSBJoDeHmEecJViQr8y+rSI1acaY5d9QVHGhUm1zy9hKFpGvFZay+bAQV
zGtlTjAB2fBYYAQdobrBd2h34Nv5KB0lU23jFoNZbF/ZUWdNejsG2j9omVaetZqEr1TZRzdtSGSA
yvjRQU3zESzMdfWm/c0hVhKfg1SOvZsl7m+0r9CynwqoONoR+wstllw/UcgNNKEYiSRKhdzolWzh
ByuuJqtEbC3G27npgr00nz/oS026wi6Ctazefd3fKEwcdKbn1bERcX1QmfAgOeg+Afuy2Tk0sO61
45rj7169V0XQM+XXO8ckPQ5MaI1d39Eij4agGRAXRpFS8nUgcbK7Xm7ufMfSaxu+NeCcokbn1uZZ
9PjbZsI6Ij+9lL4i5oH2itxYLqOKUWxWxXNlvUzk16uAD+chlttSZhcY6nW0IgD25aiLXP3nhe3T
HDbuoKOVtkTe5erlNLIKgNBZUw+MIjXa1A1cQbfW6BPBsDkvRuZG28eD5xxpdqHgnWZ0HNSlsRiK
K4yy8286Kd40TxPfIuMNtuxTrgqwBwCOu4NThJeoNl/nz3/9e8UXvK82Y6kN0BxI1KFESnT+3yT9
dQgj6QoWOuv1aUzzuDpMBzuQIyiyoY5sQxJdofHkAEUTIsZ/re2jmULSkKU/6W3QFW1s6XqjCexs
H9TdJvOE8KZfySIoKth650a+WcIcBnvTmqhhfUxFETqc9CaYzPMoiX6XES6a8AycL9mGoVNUSwPD
AIqC3Y53QAwKy76XMWoRjtc+OPHikBkyJ8JknoR+6nuBKs0QX2JFbbmNtwv93qqEU33HH1zrPcDl
VCNyRwWqaCQE1mbUqzqy/58QSIAoA5OsXVPsMXlLSSbkgKssqLoJxUJp6/8O+Ocrq8S/fQEe6NdG
FGn9coRirak7J/eLw5sF7ItuB8PDGD5Dag903ogXYFpAc/zhSCBiq1rqVev9Crr0xyTe8pCTfc53
Dx1XOo3YQk5oZGyiHGlx2yLzpNizDMZw5yJywyGHnPAxtt4j7KDsX1h2zcLPPnan7tvqK/CfyuCG
ujdXuHbXqv8EGlbG/q8HnYdsmazo4Y76+PnuCiZ9tpoFzxmThHlvaLFL2RKHLWGROkQ+RW4ivFsb
9Jd8xKjv29gL1pyzdBFlCMJgQ8VVbNDDZeDxQJtsYmCiktZ7vHdRV9XxZYWfdKk/15NjU4rwzyYT
DVAt5kU0FHlcydgo3FBMCqnGZRniuRG8X26fs1yIHfSOaAmPO2SZG+D6mzr13uMfvw2YFd+v8iJH
ZoUuDQnoA5ms06a/T6rU9L3uNoB8nH5fR/6n1oib1qPwAIpNAKIM9FrYC7170ki4+cp73fDxqUIj
9u8lOQUTt5SrbSYuAp4cuomSd6UORlZDffuBucNsH3azTJgQRHNCaWIxFXOFXpkzBi3VWCofp8Bj
5Df7JseS5Sgnrb5YNkwcurw3yeGxXoJGv71nyhuWAp8dF5t9CrDe3obHzSCdHUeuTH7yNLb0sqFA
KhswsxMTeSLwH+0Ke4GNOrVprALa3iiT8hcH/NYOeAeu7lUh4QZOWYmNgVwgXI+DedOBUuP1MmYI
5uyzvbJKsAjcor8TVArChEIPojbGlxyaykKmCJoC0C9zU0x7vEnAYsM/xx+z5KcC3m0bbhBB5u96
fDunzB3BU7Fkuo4FTcAbGGVLYQUDtJzuQ/R6I3g3h1ERq4pc+ZdvGnW1UAT1w4qmKDXHookC5DIG
6F8YhZVAMmBSoZtyfnJyDucnN5w4x3mBvQBTzaur5SfG/G5uPBP4pklLGFQwXGspm+EmUfEK3l9q
wZ79WWZo8QHwy2hQZYfhf7++BwbYMIjeKZTvIGVWeA8lnuHzhlRDYUvWwIsga0Ugr+3gQQ8/67ri
6JZB2C/+lo1blEGy0fbdKbMnh1rUQ+pb6nG9g5tfZbY8MJdoy++yyaX8ZfC8ZwtVGLBExlEZz7wT
DTg85oBGTl8nZ54AGKyQzSQg5x5oKIpfqN7RjgNBDDVunJNL0nhk6Xr75PKyyvyBpg46r6zRWaEE
tUoiE9kqq8dotmoHPHZeiPKVAEmBir4lM2pZ4VZKCTGtlvQ6Cdb09m6ml7pDU/6pLZ24GKHAkhkO
dj3r/7tmeFqx7+Btnr+3TnKG4ZciQV3i8Ibqg7xCBdz6gVU9sFXiwcHKww+hfFwhh1iq1dqYp1Yq
ubElSIf01RUHuLhzK1FL1LNSphXqg1RBbu74B8vIdudsP3g7UdTxRcSgJzerOPS/3Fq/qqZ47Tke
e3RXVt0h+AmalOmztb+3OVY5XvYIN8Dz3Ga11ERjztVxOEWsPipfigFp4di4oWSmpTKo6EC95xcs
R40DVImYz0d9ZfSyLiVTQf8fP4dKzEXsQCuPlcV+cQyNYrgWFbiUb5G7whffTvZJoslitL7V0xrW
M01hAHM2XhN4OH8URDk9QsQmqUBYljUtSFAmLL0Xsnu24pIaaAM6Esq/uvpjdveeJ09n4PzXS9iZ
vDnB0jSyBH4GqVxMcWcXzZ//ejSU+ngedS2E3VxNQsp2t57LqPO3nPbBz0i2MVFB9lsWbG7+SbCE
WmRHS7Ot97iIO7uNdG+RXHC3G1aDvV+oDtTI0DWhTu7LGW1CyigZi6xpWmymfiziHnfaIgxRS750
hCg5TPKcS7/Rsfigp1N86a7mdcFohqOIy99hCFgnJ2Y2qycX4I+Xo02/Ip1ePjiJl/6Uzl+IY/Xa
YV98+0JRNqQbJ82Eeta3tQXA2WmOLezPw+2k/B1bqrY93L2t0u4mcvAe4WMUnmCnVygRaF32ak6q
LqRDxLd6GMA/I8BHBpIQ3jF62sSLMlGVr+AvWMz0B4oU5PhW7Hjh4WArgSYApNl+URaeXaZ8x/Cm
kkXrfimmjTU5d3sOYES7n0kzb4U781xjpru3EtlhgsiXTh352AvAq+vA1D8xTtx1Wi1UIoto8+c4
YKr0DjlH+CNZ07sOomGYPBRKAbAt98tXAu7vPklfJacv9CCNtllam1r4vTcEHgAbPzKsbLQFV+U9
YMaAFJJQRwVqRd/8vWZ6PtVOCew9Ii1cW9l6p8sxJdlm25c+yBfku4ihqMney6dfXNlyxLbFBkMM
WksEMPqDBBr614AW2NibK2edd4VjB8brzzStb9RyFBrnqyGp7qhNcTGb4TAyW6yNjGNw5KTJr58q
26ciOFDXFBMnfTI3iStUQk4uV1rxT4Z+3bqe62p4m9YoX5kcl+Iyl0wzU8FhIX8Rciz0l8WwKmTe
deITUDl0Gq5PnQiwMH5UiJ0kJKLkh2tpScohwxBQEiCv1nd1QauKvwiJfeeF8vgTrzqyeYdGU9YD
Z9Qx8U6fw6oiskxMw2Wv50GzgJwWvRlrdjEKQCGNdYBd/xmQTFLZPQXaT+ON4L1DazRdRqt9yl7t
deLI7naFnFyYFPfYvAS8hEo2DCrDE442TeOh9+VhKSzkm1JIQFax0/8QIuVqRDgHCVk4aEMsmSEn
vCVCi9MlD6wzW/uqB5DcZnvr3I0eTgfO8V+k/S00kCZr1PnADbPWFdwKzvtGA5eQWKdRsg+3nHKg
pB3h22hmlMHvcxc20HK/yNRmTy40sPWvdGhew/XGAihBMScWmdmPtax0xOepNiTtzBfyCAWCfcK7
iNoetD1OAkfi/+9L6wcSMYH+ouU6KeP9cwmV60WDOmF32Pf+SCDrlvGXGrMsWWmVSoRG5P1MjkQ+
qsfDPg5QdHswBrPUJBN0atYj0HKzf//vgRt9OErWPLP7t4Qeuq0HrmHt+H5X3YVfmwP7JMfhj0vE
QiaeovtLnDNRxvXgiE0cnmeK9LXOkk0+VejQqeB8798iXOEJvLlmzc3GmlzStJ6wR8ldKi/QJSGO
N2JIxr7MO0wOZx6F+rE3L30q7rWdKPvJTHQse68u4irgQd8EzPhbvZRNnK5F9u51v8tIuxiqQlld
VV11AfbzJhSLCZrThNBe2hHL7QMBlkS/t0SH3Up42TCku7Bpn2c5SxOucdTTh1nnkU7CvjoMYuFM
e2p0Ncrn7YYrgUxT326tCYihOIeVs4oODfb3pDtRnu8rdakiefkMTXSfkwVDatz1YcPYp7YmGy66
UYFRi3rUWgFIoa+tf0IwQXWpSF2vKYnVygF0Jq1/0CL8+9Gy2zmJaYKFl7GLj6ZR5PLzpKVh3wyJ
8xIJP7Aqj6kOQLWSBHFkS1uAplw2I3GJ62T7ilxqMI4dqgruVOBp0mjGaj+iyXMTAt0w5fj/Q+Hf
Zzp5xETSJ2/nO+X7hy2hNFUA0YsZJd8lwgYJKfx9BL4HXFjzHEa2mYLP6d1/dCKuQhoqZGx/PIup
kOYUfFEAYqgGU9ymyM0lWgAs3/571Y3R9BbeYYoVmi6l+qRxxLmcnktBboEC1qyKs+gcDQqing29
sfRdDMJ6joKEz34JFzHw6ePIWZp7K7Rzh2afjVRITBU4BPbYCb+AUx3FhrSXw13RV+03jdm8widI
ia5Gw/e1VVLMTwGGYMPFOYbj4+Q8EDYBT1LHZIZIi+9yZiEeBPnQsrz2+Zaq8GGCQD4uBApt/fTH
XwEpRiFaN7j2ACPWiCBR0wuStKmmmxhUOnfeH0oWynsa6ruwb0enmXU6eydONNzJ0nbtn5bLn7w0
VC4N9FzP1rLDTHz2gR+24LQTPHFkRD6sl9LIHHGXarv2WCU5Cz71bJs4a9ej+GsHjxMI/Wp71onE
U1IOAtACwfnnaCdmHAlCPFbEPPoic7t1lbiJif6J6Cy1Fstd9V18ImFP1SyHo2wSJObAx7yoqprG
QB+jIzsPyA69lvcLU61JWZt29RG6TRK6Y6kw0FcxxBVZuGK6aTrX45NtkR2oyXMVm8ECri8G2cd/
eRikSC0Gqe/XbUraRTACtSqL2TWFRUhT7WPsxdQ+Tm5xEbrQ/fpdjNx4RZA+SOSBZGiBHrFN47aG
u2ES2E4g1ld7/RaVKhXh+Rxt+gQlJoChQnHEVDIriKoklZMARpPvTP734dU06gsxeRHntCAEmoFB
1maOmuU8uyBBVjGxp27ffjoV1Jitn/Gm/vfbVyd/mlwSPZxFC5gTnOsuhYW15CwkNb1G9UBTiwxE
zG0ab8tMu1EF5S8nLHfwiMUvLXqmfkTEJwU7RSSOPqCW0ygX2Kwph43kKncLiByin5fIJVr1q6TU
MFsmQUpr4PWvNUkdywfUgFfGkcH+jj2Cthg2dkGffRtVM6BvdihtHT+JLwn8Nr6xZ3/mccyNJYsw
6EmUpy9Kuf38JGQZFvcz9ecIKo8e0biBfI/r7xaNkWIO3rm6wAS3o0YGim2BDW5oqtumJIFgCs7s
EaB4DNKmrv8ZZ9EsT5VIiTu4qMU2HaEu/we1xLqD2Tk4HKcDl1bZBx+PoxX5vKCoRhJI+pFWNXz4
heGPcultvAvQMEa2yqbqi4JF7oehYlWbDvCS/HNYcnmr/3ZOyFeb6dC5J2TB3ITcG2okHD8VWAVI
se/OKpeCCEkbafS6KYdpo1RiPn2KEz6zl61NGR4AcaJFp0S3S1flpLgq7dMhrAxQf/liabEfAsll
wFLaufIlUxHoLf0CJ0vnLjT/5eXjw69szY67lvWGhbsNNfG44ltLdxVSFnBxcyYWPo2WV6Ggczfj
zj3WSUKrqCJ8IQ/kbvxiZ2UoXd5rZkWV9ZCjsBsciYew72xpV4YA2292+2NpWFTZv1fJF4wStEMb
9exuENIX443Z4OvTbpyee7OcnYXbwi9YM7wir/PAQLfh48rSRBssUE0dW80C2s328OEn8F5BI44D
hL36VxIAkXRCLkMJAQiOOo1/DMRvUQmVC4F6oEXEh541bn31LnC3cUoCafDWcBFz6PhrICywE8i8
SR2eUojZUV2UjeoAISODHBYwcoYCknJFUl2lNfOObe+3qhXLxD7hxRq0+AMcRzNxlWSn83ZbKvQU
auiMQHgnxwn/Q1kcPq0wi4b/cbw5/5eQzRzR9CzF+vnqEpte0Df8xRHLJKEk/7lkkdenhnpQi7Lk
XDDkzdvTtGk+ZjseROiTKzVvlbtlBrzSy2S8hegSF5sG1khB4sPIkJA0QhuCEovGw0HZ/Xw/0w4T
qIdbrhvu80cf+uhvektXAcp21b32YaPhtk6yBk/2f1dFFPv6ocpdkgFJn941V2bnqxdyc2IO8fF6
TQ/7Y/NOXHXeSwrc0Yew2ckKATPivTUfn+rVZ1jQUKnVrZlviJ0Nl+HkewTdYaMWDa9dDIIEhS+S
sGPUGAt+4xnNoXOxwcRXeRNN+tPCxZ/C8dO0zqR/2h7SGIBOcXSAWe3WI7G3yaB12aS2YUVgucr3
/CYYGyy/xqtQkYHsklfF5xwAk/nHScciFH0EJzT+c+I7TMYWu7r52JKC3aX6kU1nTFD2xrVHWgWj
jmr+bOiB6TPedADsihAs6a3UbxhIktmvMYRUOI0Qh0cnZo8KQxp2DwdEUKVicwjPc/spVodDKyfX
+Sz9byDl0o9rWKszRkMMaOEJoHyCVjBQtxPlZ6M85ItjICFGziLjnUxhJhrQv7NJ+cQgF4QhXDO4
ngC10AO8ihnMg2F3sL7T3C5/ZP8K2rQU1XAYYSdHM4bpb1MOqGfaMnQ2XXwjDNqYjIPACpCEBYWi
T/jQ03lR4rn5CUTOgraJrTmvWT/cGUeyfti03CaGwmvALw3tTIvxqa8UcG+DutBc5i+5lBLDn/FY
V/w6GA6szHrJJBShk8ltIl0c7vyLs/W0kBZojjDNsA00MoiIZh7EtMrdfSEMpRWsAO/H94OrlaLI
kMRmWKR2p54qDs+6GrH9ks81Hle+YioIChzoXesMNnboLPxp+tnyqBNCnw/nsHddXxXh+YftU/mq
ov9TnQ/5iW35JRQed8gWLmNQJGKl7ywEq5imopDgsQR2RELbUrIBWVNAXEei+DV3YxuUQXKJPXVj
U8ZBsGZmFs1jr5aDXMRO0t2l/VkVyExdWu+xDjkAWBr3sBMMhc+SL3M+595Q6Ey2YzNKAxtwDcYd
ffQ7XUSQ7LdXqMRclo1dshI5Jno/6oFrq40oRar9mTNzniFXjV48aOqX1zRp0ZHF4SZ0P9/fgvUp
f6DgwVzOeD+W16E/IfMNTbCMbmUaZnsm+NeiZOT1wPuOttKQuY/a6csc0MWPNRRDhNIl5AQ0xY+J
WKrPL0rVeWLRFE3ep21r56KqbkZ2IYGfYzClaFkAoQUp+zV5tOQhUSe8pNrDysfFFhAFo/aEVjFs
2eulIsK7c9b4m4z26cHkMg464oNUjbesjXzC+ww+S8sohhRTIMY3Xc4qvRxxgpyweeiEZTUZmGJj
7E1QqM41XnLMbwd4mSCWq1SmIwBu6mFcYOjQUhE/5kMTG+jBdoh41YY4p9yOudDEnGd52OfYZtiR
1On9lQLbENB3TZ3XdREyyn2WxJvTsglFOkWZ/WE7rvYtkmYUsI+w6ZC34N3kdCWtBRMat85Un16U
Se+RNBo+CQdKj8DoJyJRIDfkBM325H63S4nHUtgEUCnsXxDKEZuc54GjvC126ILZEv6ErUnmsw+y
nc/2+2LiZh9SjknlfE7PmcDSLnWKBsIIchbRGuDCRaQUOB+3O9ggxjZt6C7/mWKIqg4MKMD5lxne
9qjXyS7/W1q/mT+xxiPva5pu7o3DIfuZo7O6+QjX8GPFQPq5OSnsv7F2RQhFOCUo3BEyJblRGCYY
4+pMJGw4JAjUs0g9hA64GnCZgFrhUk7lEOkOFuncHNzNFD1KpV1DD5YaSm3MBIn3GjG6gYFpXJEe
hzYepvYMVPZ0qcNAGPzAh1v6vUNC8uU/R+ubD0DNz3t6dgAI/fiIEhX0o/SgnQ7A0QDwf2spAeje
gj6My+jmg7uqoIlluX7OKqX7REvvzoMd+bb+KJ+SkGcqokhyBAb2XeTmZmanrTRP8C10AvDA7RFY
O9NNuPXHOp+t37cwbGf5Alq0L0AEozF1gNlkfBPfKuo9FQ9duDzVrJvmgkzcBk9dKoVfydyuNed/
KBhYKnFoS5JtsaxC2Mp1hfm5oc0+PhZzS8R8EX4zDfRyo1kRQFIVetLU002UiBSIaOpqZtW9ySQR
gonPTm2LdQFO/2Q2j3IKebhck96L1wAxaSDmBlst4h63ZHtt39EXy830oqdKWYf2vUlLr/5I7Ag9
We0D5SeNC3Yb/Tvq1uq1DV6iFDNLVBJJVCO8zUT3fuDXX/hh7aGwjbHeOaQrb5TB7ZwVRScy595w
wLhHArfFtYogf//TvFf4mDR6oDWCpKU+UFvK5oI/a+mK9Pc/RD2LcD544xvMN1014JTr1EHFgC4L
Idzyr+cqbQwWAlf++w9By8Meqp8TdAyw+fj1/pgj5Xq3rXB1oBkS4fAnNxpoYzobAj/qWfMKJIn9
aROJ20Qxj90FT/BIjWXyGu95jG8u2XbF+eyqLlCNSSAHsvG72Dt9O/9fqhfiC+kjfIHK8MGQcT/A
4/9xMk92/1q4HfSZl7u393Paw+ZPK4TmTaiXJhEmiObWfN4/52T4dQQ3auNnfESGRGDXE3/qu/KF
EcGu7xqAWRQh+LYRZYn8d73bgfZAlfvQyNy5XCgrfUnRVo4ifvh3UZJnK1up6MocCWo0nAzhCUxc
nY0yOTQ5gCJ1iToF5WDVcmeksXpMiHg8mzWeif8HbK+OnpHG+DZEojh+k2WvBRaZVMNv5uLmYPQj
ulqW8gyD48i5J77zDSj8g//M+ODLApiS3yM9OKWN1rTK18R7TvdWR1diMNcoXDU8qZpv7+9Li/Jl
dXlUI76DrjDAJb+aNruN53/hMoZ4tPlzlQ4CVzOVgaVtEwrC7AtEpka4awGmDEER7G/y6CDpm08d
CflRX5atQoxeGN3TAcVlwvjFkOopjpG2MWjztfN7P6TWdScVGmhtqxuNkMvRqtSRTGN0yut0R1ZL
TwqoaVJ+EeUlkdAImExr4GlmU2MElmbCAV5iVOgxC7v7ezgNuKulXdY6LVkujleH/iRfQmfHYvCj
0tUM6c6qmzBITn/HGpXVV4kAAbcrXZJjd56ode/SaJwnObZ451ClUfmOOtErCjRlM9DTyXmGDH4C
aVcc2bLlgHGhxsGA1+mO89rycx3SWhHj6vg83P/42aSD5hBIwewGmisXShM9EIuEAZIrjuXePxdm
Vu2Io5djv9lvORdCvl1Ww8dZ89wrMJt5weOgvN9ePQJ7X/+aq2rjaAzVP9MIjnVCaOrbKb65ucSB
UyvZJhfr8mif73JiM8TzZBX0sBztz/dU764aie2PIg1wvHnFvDx65rLC38TZH6LQ+kvcsXpfFDdZ
OnRH08n/OQola2Iw3FYxW1a4dXkETB0ZXMgO0gvaB+uebcTj2cxAaV66+CHXcF2v+qqeFEV7u4eh
a0G27fzMBSKrhyhj51KNh4xY8bdd5eJSzg8G51pWGr2lbtzy3G3YqyQeaxvUkiZTf+AIsk6k0XzW
HeSPeGoAU484ggZrXoiAIRWouwvxLVyK39tn5gHjfdx4JXyRWqATqvYvLNORmWPkzJMGIS0t4wCa
ZIWv6qSNMRh4wxqfggoSl7JTOzQGSlC2Ev/Ipmm3+VjYNJAKKeP8lvr99ZBu62jI+kYIqxDaNM1d
pinLsC1cZGFGLQ3ZsFxrMu7zADHZ3AXmYDioH34OsCOOmRsM3s7yos+QS1QvC4qi41SZ8e/WPCwC
XN1ihy2TFBVMW5e3OYBvIAiMDWx9Sok6F3y+mg80G50F1gO572Cd49sFmlpJ4m17YGDzDRfBhu/d
hrxiyLT6k6pon7d157dP4V9/0axufQzm+m4dGJdc2XgSBSYhtVLyp3QV/8C3AwKpnAFkUHg8wmR3
DlosvqzxDajNUfJWd+1SjX5HnGC3ouucV+ls18U8ZFAb8gk5NUm92S9+A5hG3Cpzg5zHkGijnI1p
kdQwUR6sEJjFC/Ap7eg7NoRhaMK4VG9k0LbcH9UuvqEQT4cDeqobA31+fP9GjJjvzyCAgoErdnMT
xo5PuEN74DxQ/2KkT6OzUm1hWBFVjY3hckEVmXHgXAjDVbbh1LpGAZsrvcdpDkkKIlwZLf2Mlc7m
SXqckh1NJhW7htzuyR+bjHD3pKjgtcmwv18XkSLb/CQRMZ92qelPsTX4zHTJkg2O3mbhMHvQTyHG
Mbx73umWQnzLNgqDzS0SoOuTfnZSxbszyfqH0BFwmaNzOI4Ruc258ewILmwf3gqKxiXAdEr8eq4d
mZd7+R/+jqBpXU+/p05k6lKJsQOblRsJay9ehSxPRrw8Mm9olQIcTVq9qYSEv1oGv2aGgwvio/jH
MaHhbI61y1NJADZB7HgIMZdU/3/FkjEJaBvc3Gg1Gb6ADpMh0P+Y7yyc9ebYSDuLO+9bqLoPUtuw
Yt9heyVLk++JwCvHCk1LAyv49GlAwY1HAlZIrNmjnoRLDxFZ0ITL0iAbc2tgdbNStCIqM3PY8ko7
GReKWBPE/tk2X/88S+mF2XxZKElnwK7/TNkbv9kYuCNDoGypUO2rSDZLAk9b3Fq0AKYpb7KWWiFW
MmnuGvKomIjMybApGKxtZlqMMik7CcLBcjPUeZ05dFJ1r9x8X1rNGVwmekEvSqw9vaHjRiTs05Q3
3UM6NHLZxxnPZSMVNliNiHf3ZZRbWHwQckX+REZzfAMC7Q+Wd6LkSDiYS7ZfhPBS+g6z4Jg55ARj
0YrgUL623D7A85etgmX+BaMzOuLGqaeI1oEJyOTzImt+Od/qHYTdeVo0z4o4huMRpERmXGWENqZ5
mIAQ7Oxlx4qQZy95E4qBQfVtbX7Opg2Fmb0fTbQD3vQQThKbvPNt42TEi0V3PbllP58ftnwkv4VJ
4AB85NrTubj4YdpaCtqxgoXKM1b0YzJqIQ/eLKzbRC6bZCeIUnPKqFe8Jbp9RblR8sUpy0kig+Ay
m4CGtD+kPUEtEmQw//Mma6zya9dunAH2kMYcHvKMZ/ZbUSMbuq2kUh+kWeM0n8xat+z54E0pq1lb
RHK82wPYLxvcwjOsi03b9Os8aJfcLjXCljbNnDIIGGAcPO/nrxWRYMFvOGeNRFhPPEfEXkeum26o
xoLfHUyOq5BLA1yJBjHWaDeoQ7ZrNjIATjChkEEog2fHPWQQ+x6wH8pDcBpPs3Q9LLnfQhOLv0RJ
cvAoRRiu50E546lJeYPier59nle3OuJnwS3zSarSudjJ69I0K2oVRKOnnaBcgV+g+LD/4uO+7Gi7
pN3ewjl5E403vYZzOgeDJTOOvD5B7NXzmoX2wd4rFj2/3enyW1nNjm5/+HpZr6EVz1xx0TizR/Lu
ubtT0MvB3uHlNm7KmyrBaNHwJmp16d2HxggYNsBwiTfuaBtdQZQ0nNCInlpzPguLYo+/9Q5qKyJf
mfx6Z1kWWUsUsMHFDkhta6exY51FiH1ptBw8yucx2lyB/7mukZz1p0k/x1RBaMOSAC94kWA5VWsU
wFPj7Zgo72msUvZg9eOCKy6RIt3BVZZqoT4I5pfYuvLFDxSy/onBbIzu4LSPejEcjrxMUrN48Dbx
ffbFhBPnvlVPPCBo0AKB5ulhrs0olccSoPDe6pZdXeC7W0E3E+8x1WHMmY5/zGnHQvmDW8ZGq1fb
UOxEXXq0YXXTNwHqo0FfQbgKOhBaSzDuJakE1eCQcTlD0/E3f4KHrUHoA2AbizYrwprgmSDbCL9P
1rAMGY+x9tod8baUOb3gI/Mrd2On8q3b681foThHt7KH3UHFry/O3uocf06XkzR7gtQoVgu45e4S
kbZl3QnTVimdift1/5Nk85JbmqK0wr1RFRjytWVL34Xwvm67mek6s+lniQs5xr1MRD+VcrBtInhg
QhdlWwY8FCRUv2F7mj6WU1BW4ABuef0OJtnp8Ope7WVGlj99Etxpp97hxQ3BcopFDl7NCs5JlobN
OV/E/PRWc+ZdEak3sDyLKvZWCeN37gK5pbzpB+UHahxORfhf1kvdRbCV/f5z9k5wyO6htdB5I4Rh
yyUSPhzAho/OImvbqi9gnLdJZZ5zoWYgRJuZj7AzTAOeswMbjSEyHi1TGZ8xRUIg0JoNHGI2JHvK
d4MVLRigICl0fmFCJpBtNXDGxOiX1u4gECmf6jk420J7NmGbYrR9tj654CeMpRFCMNStg/C2et4r
eUrntYr8P+/634wSyr3Awp3Bi690AetcQhCzRf3cEhaOseUUUwcQb1WTyBA+0SraEXEYGkHqa5Ed
MVvP1sAy8ZwR4iQmec79ahAnwgWwcIDWvbybqvtGZdpkZTgpghNNYD8cVWNDUrAyFoizCYki98F8
fGlp5oDYn3IBt23XWrL5oy6PnmIxglGFs2k/JCkXObwGAl1n2+GbqyJGZf2vTa5016UhciNQsVhX
98cM4WCsua/67OzKSfcx30OTJQmBIhcSg8RwL1CxRFlP1DJTuLWe5uHbmfCdf+imhF12NAYebFfi
D0LI6njo2yHyyly8slTR+XXwC3CArRwvl0S7h2oR45F98xr5qyLQwxYJ7O48H9ALN6dsWZ2QcoAO
BsgH6nD+tojaOMl4r0eTvtRIEhiRLek3RFwardLoTAbmKS/jGX3U5gLHmriWIKZxbalm9GSmYhOw
IIUiEtmYeYePp4LvYvV010gp409L4IFRFbfTZ9BAFM4BQ9Gt37LN13RQBCg5aC9HjS+LlO/rgsG5
BURcmsshjwCYBeJ16mCsFfphzY0ScbU9d8zJ9bk5ukUBwNjRu960oymggKUjariSwMnnAQRpoTi9
hIRL0PmVNatNUGnQQx1yRj8E6fEXuwRTsiBMNnLnEAY1mRGg5J5Rnr3iPg94WRnR7zjOGiSX/HnE
xnLZ3sAs/5QctvLtnKFHOX4qSPNxzNbF2X5gBUTSP0hYoSEoKJypNH9NLBCGQfkV6eji6SAEH+zu
cgbfZplRpTKJi4ZDDKIXbWcH4lgU6IV8+bwa+5uf9w7eCmWh33Lxj9zXLtwQW+cScQH50W/qhUpx
SSzDN0Ys3Xf6NPj5CntkmruX9Oiegx2Gw8aERFRRTbESpidDOHEPJB4PJjuMCbIrAGFQZWdhrpaL
4CG20AR4YIaFV1ZmOECOCA4BWH7+s6TvXUfcVz+3sk/PO+dAnXegarmAIeKrbG6DSPxFhwOBFwfU
j1Wz9ibB85oTUPY8CHMiujFJHfQzf8EdR2P5646vHplAkHOZCmByhoQYR5f59x/LgyCOotsKhSmr
8omiw8k6uJ+8u/ZdQzfjvaKKdoE+mM1CJr6saY/kdb5Z8rVE4YWZwkfaKriWUEuoW/0KcVZDl8o1
3teq8k9G8liGWTNyj7H1Tvo2z6kDTPrTjihWRi8dkTbicJ+V4V9IuoNzNxLEnRI3nDZFJTv3yLpT
h00SZ3VZP0FAwAyoQ48bPWXLWnqI1y2UIVGG3rvaMtYv04/xZ+Z2cioGlQ4B1JeV3IGM5oZlS2G+
RsgDdNPsVKkIPydebRXd3R3bx0cjGMIJxNIou/SPU/RgZ4cx5rNm/64dhE3Vf/HRz3JzL5gHAUt6
ML1Q0CxPP1JtRxusXY8n1uFsvOm3Wiw3HuPY5E0XxTWvwNh6viEBf4No+GezEdq0KIOWC6NCfds0
DS65soyUsxtiOImLPNGAO15x0VGNC1ezixoA2i2JtoHrKszluYXMzDSv4gz4HyEEhuXvqag7Kb+T
VJJgq1GQGD9SWeNNKVC9GitGMqoSwCOEwsm7TcUS3pYF7D+KFLHQZcIru9TwIwm8qFV5GqNTorzo
dScHMpSwwTPZSpeSNuokfSE7W11iN3gxFzX6hu8wBQDu5IdDZJ+GDl8zCFKgn0Tcsm1gLwZG1WL/
q+uJy3pu0+PlarB30Sf0VNU/jtPP2mGMWyS2gsFsUWTjHEFBM3Nskp4rtV1LQEz5NsDS4HTO6s9V
W6U4sS+8TNxGzCtkxmPN4cVgWocdmUxO8+rsakAvOaFHM1OBPbZk+bC9oiM9oQVS8oAmNuF2RW3c
T+XB3wh6ySlHpWCHR1Q9jGp3WG/um1zh4Dbbto7ezkOPW9wlTQgbsUb3Bo18OO68KXe8uvGQiFGG
mKKW/4jZLbFunuNcZLvQh3JYri+0woOybpkk1GWGb9ZmkSEJO3s9CbnNDGUnC2kH3XJZuSr28fSD
y5kLz2KLTvRKmqvH3cpZ6JEHXcM7UTcXF9dSFRUCk/tNAVd4x6ZC3nexiP2c+XKtIKAbRsol/RET
fUDir9+vSVFKBTikYmW7X1+QBhRMmpEvvPlncfbt4EkmTldSLckSx6NbPsT8rrMk8M2ooS0Ci9Z6
0iwihARIk4voACkqRZFbhB92xlj8l3NElg4nX5b68C5dtNJEQPszzmMrJLpFCq3/j5+SRR+yxgaO
/HHSC78I3AI3JIL/xz6phzCdLjsIY4jfsIvW4OvuYsjRMzcWJWiZiyVG4Wdi5owF3CiWNpuaE/Tu
88fk5KtnIExVGLckVQ+0U6LxZmeQTO9+Wi5qOm1hCaxUAQuzJLiAV5DDRml7XdTcqDuJqUSTlEUv
gnV6fkgdMrxkcofMmpKvl2QRWW57UETitbELE6f7LoKTEhjN3khx7ado1qXCM9tCZpPmb88R6Lln
m8IvVf/p4fEG5M51WOfGwZU30ziDA0mKXa/yqj7L4fOA/X/14Hspyl+Qv1rpbw/bh5f5qO1iOgbm
RdsTur5evtPlmLpBazvTuWUy7EQ6CUDXB5QJeY+mc/QfuPr45RBDPcZbHvkwTmgXO6EmnxrrHNJ5
iEFSrAT28NNX2CcqKwKaVDjY3gVmJjAbRDyRAEClN8Sw6a00rj1GLJjsPCa3dhqqDnkJ7Lh6uBuA
h6j2m5D31L7bT3kPNqTT8/QyDMcGch0eldyU2XWDy+MnNt+tZZVf4k1mjPaHAIrw4ByRYc6Y8Z5P
NzetYCyJWtoON7VprYdiDaGPCGvGsIcGJhJ4uaLeEGfqfe2nEPXEYheMrGbq1qOirsoHcU663U9B
MY1Nl9ZhBKTOgLmMB3D+LERG2aY0dBLzVnnO7zyCY3rp4m1qxmOBuDTDCa0qlW76s51Q1PnF6UsE
oQPzhug9uMiTwu7kQFHx5B/zRiwyuAWGgXzz162QZxwoYSeJuAcKWpuYYRNez0frFlGjbdjOdGg+
L27a8kIJI5ojx5UbWUCZUQLvUleZ9iBBNwCEBlip35ZjMfspjp1KtgXn0f1aSSXUea4wTP0qY1+T
FO09hVT1aaI8R9y8NSjHIP2pQc8bPZRV59hTRbDiRskSZ7JSgvKUBdrRjSvCqqjyEouM6xXQDdK9
wUWf33+tDvCFY0bis4JOTrrq7bJBEo+HY30jb+k5i6fXEjwYZOFrVt/8yHJI3i3Hzjm1/nBt3Rbh
K7t4PZFuRi+5wp5WgaJegnYMu0vARZgK0wVqcJT0TSCqFywvR4Pawtf8bW40OYl4JGufYIlY5vPJ
I+Q79E3i1kiyM4LMlJNReIP6Q0b4E3ZusAydh4SQ/jx6YevqsZ5C+u2XlkY51nEZwYLK5s0FhX60
2YGLHHcfUxsRDpVCisizUxxzax5jQkTKuHbCK7cryzmiCgzSaVx4jsAdIaP5mNV9yzswBZc8HTwq
PMtF/By7rLJcN5A2yG/gKr0Dg35GJUh/Oc784MjcZT1zR5EBtK1bIflp/cSdmezRHIrbkSf8pPVc
Ot9zwFexH3SWszPmRPrxi6aaZ2W6Y0D4iKs8kMz/ShYXGzpwTJmU/e26o2+yHW18iDeBGSJ6xmLS
z3UVdFy/frc9KOn67zqTynP5jScNrzFyxdwZYrI/sEyRTTizbhCTWcNkSAh0m6bOzNQ6eRvg88rB
WRKkVsZQsJOWCXiDA1GDY7wATRyeEafkwXxEBmVEBCNJ8nyPtglJABW84qKLKQr82k5U7WkNMO9i
UokV0omnbt1ROwiZ8HC9myCv61XVZuWrjtALICJJSXemd6IWzWuZ/D04BdiiUxBKrozPdSkPrDfj
VcPQkHpyefLo30Q7P9nSN5s0R407My9x4Okpqg2xWX0cQ1KZhe7KFdE5Yl/5GC7eMLFRcHGxkQ9H
kNYC5qcLUVoiwVKdnhbGC9mobVWrbm+xDWR343ga+bdpQJpm3H348J92JS+l56yK4l4PJSBGktRq
iqQISFu7bSZc37KPF/Le+ED4elN+CPZxSgsrttck9s5ZT2sjJ+VK2D9gkT/Q134Z8CZ9ahHkE/12
EqT8liBvNAWKNo6vtLjlodgAKrT7LTd7X3Q7VSzF6LaE3yRN/MPY/XYrAYkOlsOKr7WtM+3bfUuH
pbJVU53sECT+xS8bsa/nC76zUbLDiR2LQiQ1fj79HYNXvF/owYVJGG+J/d1FCtXS6YHqacJRfGtF
uvvtLFNzGUJNFnWFMclYkl0fuUBHPTTeQGiimKmlXIb6kXjrlyMmoag86mfsnkvTmoWqRBNhPsOV
rgNDUBUzu9X1HFTBknxLs6EOgN45U+4w9koYWuUcGeq88a43V76gPU3Yf4uTKnXib8aY+K23GABR
qSyRFPGO4cGkJ/AVPVS8CBQycn8HSxgbPCHZ2XqTlm8ta6iHL2XYdQZAoqRmdl8NT0WUThbmCniM
XfI2LazYGeDM54/Kzp/sWbVWkb52DOblvfRlanVnBY6qkhQwDUO2qHQvotw0sAZ9dXEPQ5ciX/ph
nUcxVhKf9dtX9jwUt6JuXCyqubXD2rkUR4SnEuHnVBEzXDu29q/UhXQpCcABAuNzoywodEwPuFrf
lN9fvOF/2q299IJu/6A1qH+Rwg4FqhUN06nuzr8nKa3fauqyHiLa/6Bye+8vaGFDtuEKwjN7Kw+6
NM7T7VhBpFGyLAQDDx1/dpL5J9QrcrNHueD74/WQ4f1eudSIVEDRrS/1I2ef8Nyjt/WE24Cmj5yd
wDdqAQwae7bJh4hgwtGRXufZ95D61b67xiV67XOWi1CnaYGk4hzPsCxygU+KwzfGKcSz/fdNZ9wH
pG37O0GVZmho0GcNpdPijEuCf8Q9Bna1w0f/26oPo4lG3wTPyY8TWnVWq2XQIsyPsNVtSP7QwMTo
cr/U8b9uiJj5zI9Fg79nItHKOb1Tug8I6HwJYfVaO8JrLBn0H2onSQOjBC2AlwAqepLgWqU2Kz9r
61sO0JoCYmTz/E4S3oPGqV12z7Ddp6b0tEoUxHoLyf5m0Y24YaNrH9jEG/P5cSK89B/1ZjQA3J4h
IW3Wg0o0e163F30FP+jpMdVRaOaYqMJnvBagmFPTwj1lve5wsQUqEFRJcvou4lR6vzx96fQ+syT+
zQh+lEBGl8yb/VaOgrMFRvFfK2ycLuy+g9rW/H1f/GqtU2xRF9e7nN9LwbF3djWXj5m0aRiIi2FV
OlgrIDy92DRiS68lhw4mxj5oeqn4tqEmYcKAyb+f1oh38chUx1JuR9kZq5/zYR5iQRk0eXlLZwKn
V6A6PGK4Vj/6dTJdvdVzXXA7M9SJZ/G/ESyUSsxLYsSUNiIOPAQO/zj0BBqBTCnmb3a0obdys8V1
sIqt26sRIROPMp4paxEdZSE/eij5tDLWTvy0vxrVEvil0+pgXQ2k2He8y1kDd+WtYEWnhXanOBv0
iTit6m3y96Q1y4pEpXyWq2I30VFm+qsUmn84GNu5r5DD83xfOATsv0L9n6h95pICo2mNaq9oW1b+
twY+dDVp3c9ElI/cO3zKWR3gSGTUeDE3R1EvgfFhoDaU3YZsQoOeA2al0X0iw3w60uyxPHpPtQ8U
nnH7a5FW02hFUJEKDLz6h8O6/J3+thj1msNc3rWJWfIuHdQ0QroghlmNJJikiaIMy2rTMu//N+JJ
UizTFivlFaY7HlpNreT7hcPw5ueJW1Das3uyFfCf3TCwOikZFPjfNQK3VnWCUX/xgth4W/2jogGH
DL+cdCxaYZuBladPkQnRog79IYtIBpsDAkddOyweBLFOT/wRdm6VaoamKz+AsL9X9dtIITt2PGPP
kWOj4Z1Jq5GqIRnqVXtS4UmF0l8kmwHza35/lW5olLVWlyl05Ixjea073kjVIrIThvNxSi6a9ZzY
qzG2bm35dYW5UPb+Gk9YPu07Ag/3LUys4s//nmdigNZpnIzN3yMLvRNpX//BHqLyKIBn9nkfqe37
rdsBls4YEtmKUKFZJWHuF0cWrihqEXkneAK21MgDzD/Oq7+9M+mOsownlFybfF91c5it+lTPeYkm
ROvIrcHjpASJ1WV+KgTKK3bpehZKBlhbG7pCLcNbO01LU7yEHWrA2ULVfpYlgSpkr0H7UFJI518/
3bTmAN95/fUCEoKWI7JnSosX6GrAlKkm65fiSrP4uo7LLH6QFnUk1OHDIMaLaVpr+pkkFLlFS5iE
15nvC5ogETnCoGUGNAj/ho38XfgK1mvK8W2df/15mfu8eAMlGH5ltbvoesbFI3nJ2R7H6wQr1IHx
NqgzZiSyB++gsYrky7Ar85f846L2c4AHggmjvMz/3sJVU/ei2MkX4yHKLlN00ZHiJsi1t55STlaH
oIm/F4q5rYo5/QZn9TaIkmjqYk4mih/nvrYcuLela88fKXLONMUb/UFMOqRznt+78dhhUmCUy+nn
zf5qw+Xej+9OEi/lrcsI0syf9i4WA3/2Zk9qe+s6er6Ecrgd4tIg8ctStQ44bO7qUIrSJJwR303C
xxzVkjLh4ByCdwJoWZiXBxx3a5WgfHbuBR8Egn9bd9GHtygi+kBaT7m+bo4lX07k0maI77damLgt
QqScQfIYZB5RhsMBk6yg1cqGNUpqCvKVOs9vpj2OQb13njDBD1uSD4VA7deinLFoxbTfehLk60B6
Fk3eZJcjuaHP40wMu9K5yjO2yRtFF3bvQFRqc6dIyJh/PG7cJvOGDo6zj6tRKIFhPzKec2JCFOie
ciLh6X39KeJe6CcBZQqhY09HWjZR6gEbDzgPOBVxhKsoYwUx3QZIumzBgQ0EZa5LS8VWazcqpOsw
gqKfIJpUmrBu8OrTB6XAtsNmVwFR0dAlQahAYXPv0Sm/zdUIz9hmgiFMVJETLekDsIM4sRJHSgzA
PDU202dLsK4XxmHtYDeVYLI4k+iNVKyCEVJk1/OZQpudStAIKSeA1VCd/7lugOWrexP1hhXvqEEf
Ve1LYF8kdfMjviXCis1N0ai2PeKagfcdqa4FO+HsIVZj+HzjRELQonQOzlV/vWpaehJtwkjnnyKY
zY7gvun2uPvi6vTO2kfYWem5XIprr3CH+eosSrjIO5WOROeNxR+oR4+aiub4uxiAgEdEb5Ydop1x
NOZ0zM3PwOe+4rvU1VLYRw5hWk2+OpiZDu2NnoRdAHz9Z8RjotWOg7lTzRVbiOkZ9fL/n0EVD1b7
y9Jduh8oObSI6gTVLSylDAStd3wW4mk2XSmMKrbzsBYSotTrgsEiYQbRPHt8nz9n7+Q9KQSFkIv6
KZViV4tXAjtC4q5l4VdPJogNI5FshuzmkqaaFZEumydeiuW900/hJVsif495s5T9pLJLx7mKKrR5
JY/H30iaX80P2lC2sA/sdvdyBCMmbRlUiL3J3Bz6CCrrtxqDq6XXNJccaIMRTP/rGOWC3JbGzSqY
mShueMN2RIgt+/ps9F13D8S3krclfH+oTwFW+D6w2cmYxq0GjtbXPFk891jh2T9uj0nUv6nRvXvy
rJDS+/rAMUuCFyOWvg47on6wbyhA9/zhtDMMGNGZE+QgRNR2w48qZY1XoSorrzlWusIFgEApn4YL
yogJkmjQTLUQIZTCHvBvV89dtxGcLSlQ9Z/usDZCHu4BmNg2XOk2vanKXHs1kOhuVXGMa0uUYkk8
eUqJ1I6JMJWcvolQbrBDTNC+awygU6beyhDVIUR/Bafk+vdHXu+c6NbUvGyrSdBVmWpPF7bkX0dJ
8XYSV7oAgsIEjhum/QqVGU4a1NI0iRUDjZ50LffKJBeaFBwtN1lSDeAoc1xvHXlUYQnOptGLmfqe
niStvVrynaSeyprpe7biTSZr0JNP6lRuiO0hyrxaEn5R+mphngIgByIiDR++AChyprleGkpO2YQ8
7l7XA+wJ4uS59qUDW7vFPOUTIvYy26SxG89cI8LNc8gzec6r50nPhoT4rwpxTTpPWeNUNGZG7CPM
kZEJz4K1sC5byNP+9Pl2PSJOQsjBmUuNljIZDnSkkQr535a6HFXjuluYB2nQvbUK3XvF3fuC3Hp+
ah2bS/nfSkt4wmm0KPc+ox5VcXbjLL3tL75SOn5fR+J93odmsM3DDYR6UmusGZcOuWPTztlr8Lle
2j7cBqthvZ0Yrmf4m+NevHHCb5IC1LyEFajf7ODBcbs2O5YQdZax8xiIt8oUYfZaE4dgYSUunm56
MD70RncNGqLX6aPPArmfBRmHBJ42AKsjrvwjrCkUqhkkMdf68N1NfLt9bfd2YVRMCLclYT4NB4kd
Y/T6n+Ff9pA4pSfXyjud1c0gYOODmtLVhrLcXomk5LCAAq2tQ48ZcykUznwgfeVywMt8SlIrkpVt
NQFFr715L0RwBIgdPcY+O7a9mLZmUXhiKE7XVqjdSK2noMWhcLmd6Z87kBoNKkQJXttMbf1XNKzl
FkBfTeBTrpu0ncVZyPCcm7ORHKQ/9O/mp0X1A86LVEBWtgnyt8wEnAOyMndHxIDDR/2UlKA/RJ3Y
sVvvb1Svm+ZnP7iUwHD2OKoclYj3NFuHklUCfeprQdkwlKyLsK4XJnb5jn1IPwvhLQKIutKMQM6G
sm6tGpHe7pqrR2viSyTi0Uilegbl+5XLgvp58arLiAIaJHp0epUFCg+p0CrL5ZpIfosYwKDyeXch
lHrIVHIiYc7bjS662D5+mkuhZQHWJzdK1tf7wPs6cg050KgwN/F8JWQC4foX4tc1OjP4Rn1ig3lV
YmKmkty9j75FSkEzHevKvoF4tvClRztl40y2VRzO3zvvSZpTAOQmxj04ZaQ4yVmVqQvv7ozp5/oQ
vyUzCsyocSkmqJ+jj9557wpcUP4789ywRV7EhphjWaDX/DwzjLjUhT1wP7PpxtCaOB9vT6DUtuTF
1hI4IsWFLQb+TZF0mj0+W+LrwskW8xNbvrr+VyFPOsLwRIeXqjH87+d3U/yWrMYdP2mdOW7YaYmx
rtmBIU4jedLSV4RmER5V4A7nW1dK6uapgdXNi0Pklo0jI1llXgLX/1Axai67NpYn9Y1OfD342AnH
KgByhAyPrsiJdq5a3oAgYdfF/mtt8RYW+bxrrT6A96lfboJ2j8vD+7Lr8updJrYzkdWAg4DdsQjk
hzb+ECA7wpGVKflJWQ8IVIlDoGsD5rAqNH8ZYRIZ+ok4dzz2LBP/2XdwIahZV8aAdkBdQdn8OwXo
ujEsrf/hqpHZOwzxdMUe9dJOYSkGiU+cglFadlEbtNS9rmiscaijtPC2PHtUBm/2BZcpNOLISQkU
qS8m0KELab3lXGZroUx1itO1MEpENBVsCcFkg7BOuNk3du95IiPco8/4kRQ2BsnY77esRLras47e
3a01m5+yEPSZzV1YIKiDPKJvlV66ouxPpWtu7PcJrBwK2yZVuKxWJSskiwHkQIqeuZ51oX8IUX/u
s9x1bbyPmmBFyXT4eviKcLbZZandCl0V0vOqOhtstTagLDn6CXBA6rEysy8kC/HuRl3A5t4IbE2K
ndY99tmtJoXv1M+xo431b+soDbyB6143wSseooof6499sDtsCgVtBC9RpPhXeQuFhha+ykiMllqo
tnHVALzt+CZPa2cwtNU/tTg1UWLRKk5FiI7NeUbcP4zM4JYx509UGVa7AiQKqJeNCMr60SwDIJ6K
4IwSNJZQDU9JrDSuiZ3BwEDMaPfyErCq1qsavTYnrhk4lY71V09SASUrM29F6xIXasYCDQSpPJty
74v1B68ay//jOvecejI4fopOXyu+jvWZNlkPfXCBljjVn/E2mX2XzGrObx1BmNNrt7Reyhh27AGt
AeJ2dCmzjYd+DiIMg0GtCVhUt+qtiXu55mTQBGn/vQ2lX134rkWxZHNveu65GqlpWVELaMNZpFt+
RQl4cxmW2ZhgSriwjN4rnhWxyDDXpDRa2XcyrNEQaRxp8xGqftrG36pkeQ0ixalSabhy/+IceDaN
2mWvJsn2Tx58NuaVuH3Nnsez5UOmyMsjExUJlo3hPIrlc6Vd+H9J9zsEinoxNr17R9LrnFw9UYRB
ZbkI3rNpRoVsGYCDce8KDm5AQBKvjW1cfgypwGm22wWuCXVnzNQsIksqg7F9JrfZdaBvHPVjnp33
8Dys5ifKt/Ynsahy2O26NJduxM+uVqskLdfityzlDcXetEeWXmYPGeYL53keo7lMD1F/I0W97QR8
9lAPEA1yYZ2X+w+Y0uYuyE/QrXhR3FAOMGx7FKIKReWf9/eU/rJb5+/DCzqeBC4SY3JfOSc11IJ4
YkIV7DQXf3xnepYNZYYCMcnyqclubnYRi1VZc7E4Ve9Tbd5C4TD7NoJTdpNhkphA5JhNNBYFyYsy
TTH5pja57y7hKS8Z+4QWZEwyPlM8/yb6zl+nB7e5lqwOUSgbkh051QvoYd+0/cgka3u9O1izGWRk
J3RJ8jSJncjse6z3WvDcn9l4gfBNc0fqMoVC3jTpO85ml29whplsbIRUIFS541SdFYJChzuSB7VT
h7jrA8bGlofupZUtXp99ICeiIDspoTsEoWaIFJ7Q++ZRY+h6dHkPPYVmaQB5eQZFwBPi9tWElSPh
KPSAOCv10GKSvfiyZPkLn29OEXbfLPSDxh3MXuONCAAZc8PaVWC74U7IzP57ITKdAlOxcUNX+Rl4
EvN5yvyhis7Hzut72NAbo0DQygM+dldzwktrU8uKKr8LzD5aOq9ry379AbBXYSvd3k6CJw3zfp+k
NDQfdvC7cwyJHp3vHKu2cMymVgBBZi9/Ee1Gb4gO16cxX8uEyJIFHL4/jEiWbBjrApFV48Y88JPX
Rw1gnkcf9R5a+wp2qc4Vq1f5XCMJUIaS72lj0MeesleZIzzqGvaGrpiNYKiZIs+RWPZA3+VR3Els
88KPfDdoe68kyC796ACnaJfgm86h/wLEr1fsiCX9C1LnTAwheX7A/goXt3StB8udwmBFjUfRGtIs
rxbqarKhcvT7L2xbyLoiYEgAv3P+GH4sKKA7XAyBdeLoeI38TSRZ2cVqeqv/C04IQdJDFTbMY7/V
jUAskisd8UsM+B1adAYYoInlYpLtp1erUzSt5YHRvZelL6CzLExl7URcHAe/v1XIYNvIsrz6KsCK
piY8suNKR0zsitInMvz+zWkyhIynvMiGSHfDHF96gA8nFBD1Hn1Qel4VqgML+CE6NuyLWjdJ+9Ji
WGDXQpzfGHPUjIbdJ8l6UeaZBadzFlafoNlTwsULIv1Qh3L9wNmXAYL/peVFg4rnoF3+9V0dTVj7
wYKVxQzZ13vJQkg6gm3/Djte3MDZQFlqCHKv8X+Yuu3yqxdWyG1sD2P98RSlL4LfxlQvLjLrQzrJ
y1XSJvLhmi1PFrGHZjtrEzBR9G7i2hT2UxTPMu9F/T4GREVKgBjsw8HKnzh76M0AeMDd2ksicRt0
zPPBQjMG3+tLm5g++iRz3tdL/TAwWu6SYo2VyOeGvoUR4wijX8ry9FSmTrAAAVZJlmeCoHM/LKrr
ebzgTQydpG489KQmxMEXRff4ZFfbjCPso9PhrTqE5v61ZbaO0eT1EsYrC/YO+zmjGJF0pfewmpCd
zPoptVPjNfPwABVVLrOFurkHv7/6pu6QbNDDIMOxIWJItNAFkIlanw8JTYxOggHJWioqHQTcfVcF
/2D1/drJc/N/VLCsrrV1LODbb6IqJyTfDsfNvypf2PJXmP3UP/4qTsHBkQIug11RnjaTb/MUjXeP
bjzvjrF3xO6NQbOq3yZdhi+5VyQsjm9dc8EL0FU+jBqWL9S5/kPZJo1hEcKdWWWpy/pgI8VJiNXd
iy2jn42VkRKGVF/xbuHx6MkDIDVI0Yop0rA4RNIWZc5e9oalqcQ/XJCZGUWZmbDzjLx7RLBn7DTX
TNfDZz5QTHrspc3egm54F0uvAc7S14QkLr7Tku6G4WwvbiRqaFGjzYRyLCr5MGfM4mNuBXfll+jo
4ZaXnPsGtuvW6wYmF2WYH1JskgsbGzVdBs2vbOhCjGiECB2C6APvnSTx2PPS2PZQuj9VHheYfmvQ
CqHNi4CNDkIzczjTMrm3+2KKAeymHbb3tbwmKkaFFtKNaFNza29Lkh456m0IsIpLvu54brAiljWI
S6YqS7ZR8krC5vvcU196m7Nl5JZVbjDdUt5P4QHddgGhtbHT+VDtfTDOiZf680HaVJfnmbAByK4r
q8ms6XKEFDApsATLtxSfNSRoKfBo6wj0mqWdIYC1AgA6fYE0xRX4c/5b1ROeBfbyaJNBIiOAZPFB
rvo0r/BG7zi6JXyc5HmcLTvhHE0CZygJJNPt1lUzRD+PTQYkM7yIT7ku3zjlRWOETj9oYFlCX0iD
jnwqcDqqeyth0wtkVYAAAd62WMWvYrEgViXEwDlV759RNroMWPK9xcLWaqKP22cAURMmuzfEhWDJ
sAU5EsPmQbSbJZREcD/VBPt6DN7Q+nXljq3+9uG8Kt6NAGM+8BRXQISgI0y7Vt9iOGW9Z3JbYCbr
mT2M9udNoXCbo81IszNMquTfk3+hFCc4t226MoAk0pFj8ikHkRoHumhu/UQmg3PZPyMD84fKZ2XL
eN6FrKzMNxoFtVsMkZlhe5mXYstLoqN015M7RFsdKyTskuzQt2NplfTOrmZJs0FRZ6OSPp7QolGe
uyVh2FEh+3+H4J4L8tFAZToCdB5TLG0bB6q/KmeA/P2+tQhk3nGJwuh43iIjj9YWGDjRRvj7F083
izUSbz8HShe3+/HwjaydyRMw0VY/SWPb8zEM8by5zUQSMtTN+yjTY7wz409Ewx7MqklAAqcvrVJO
7AKytyyPwITlbqza9RsOmNG4yVK2SxG2n0aFdvbqZDfPHUY1AI82fvxYc80iV8kX9FVLA4LLxd/g
CIIBYwi01bwEULQlbJ0FjR7R+f+W1xFjji/BBxyXh3yK+ud7o/lKNTufMnedwF51+slMeUcJdQbr
w5w6/z/lHlUMVbj+doJlV20iTgG6ctkR71MUPeJVtA/IzGaOBPvZeOYgP1IJl03Pa8gNnXNF2U8e
M1kX/CVADvziDz0gSqH2UavL0mAsh+i69KXp2miggiw8/RAB70iXCQTspkwFciE9amqQvXVP6cB/
UBJZo7WtM3/fWDTieLLDq0/UZhpxnTTb6Tav4bqkqBav6hoLYHhqvWZ0Kg57JvqZdcceRn/AEsE+
Pg+Mstnqwmo4L0ISX+gxHVbQQXpfufMDa3xPZZsraKtxncfqiRUlvMqgO9e2kWCRR7X12e19pcK/
cJhyhqKe7ZusiAjK031Cq+HF1eQPzpXiVjcuGT62d4+yeh72YnrTcwRAwKHESi7N8ZJpk6zFA/nb
2NLpVXRbLKLOMZw0EIhVsll6Kw956OpMTTwxjHNG1Y0//Ycso7TL5oeySo30HuxO+0LUEvWD+Xu/
9lXFmKLgxNqOjmSBNI7J0XFEyX/hOXRl1sn50vRSRcQNMMkfMNcV5c6h/FcnIHQG0KWnuIymSVp9
9MRmr6EtqM4N0gFWL/1Dz2neRuvoS+vPIHsXXxaaqXlM99WbNNxsdOaXpct6dgUq2xx85ddj+NMq
5t1wfeR2W12VoGXX3R067PrGIAeb2p/R7WQPvbsYby9MN8Z/QysqmVeVBpzF6PCAbCvjslWid+LE
YmRIdgqEfTjrfXJt1voMa7ajNO4+bF4gOU1NoyGwX4pYiMsP53ivUs509TK8DbUuCpnweY4Adspn
mZrBk1lCOlgZoQ1ZP1syXyZLd7U6YNHXRhFE8s2Rm4VMioOOK65tksKJaab628Y1nf3hpXcx9/So
Kw7/alk6VvuDYPzK/6sCexM+IapRfU7g8JbOGxOCdjUgJuKMLvpgRlP9Iop7+clACxMTNQVhgUyF
2ndF9c055DeLqzDv0wr80EaAI5SmO+odAszXCFFQsBfy71i7EGmH2doQH4YpzAwqWHxQwnMbo7KQ
R9S/nmb7dGpzgbiTMeIWQHs+mzMpF7fheZ4Yr8chRTKMdMU4eF+OMUAOJfmR0x6b5AskP7vofjBY
0SsshKZVGAffSeXqZnu5CI7fb+ddaaxMx1BDZKVy4HMWqvw9QzuolCfgbdWYeEzuVQ94/pjZvIJ2
CuZNG3Psx4cKAqgBtWQpeaMrqor31tmvsEoGldoABw/Ao22/Q2Zh7qwH90NpSKAxEc+LBr9wteAp
Dvi9gNlKjtNbQ2V5/Il0Yn1ydOx3DKV5I20kSazEBNCvndaQXspyVP1rgD+30lX45/xFFqD0cunz
8/24g4OnWHRKtE6DErABj9FBhlr3aJY23uz9AyLTgIPU25U7Y3RSADmjsZqUgF68cZwVtzJhkqO6
1IrQfDfdZzgk0CZVEvdO5TKrqjyRtHkG0d38+OA+HD/v/3riss3262+jTBuqbKLjwfTh6RUKH6hB
zQFnGl9g3d/K8fdlGWgIFQ60jSV+v6gMcyQdEMFIFFuMsh9dcCi1KXzFbQWiRyNlQjmzaqo9aefc
YR4VobKagwHFj4ekjbo7gy4GvIIHz3yJsD+oH2mbpGoag0l5evGzxDCf7PxQhkwn2VHvuoOo/vw2
UMjBKEghN9/TnU+Wt8JrD2mqYhY531OYLWvVyixJ4OfNvnvJZYO6ckV4av1PUouDXJ+jNxwfoToN
vp1cgPOZiXMyxq7Cq6BxmwcsBHClptb0NfyBc1cXwFYH3W+dGlt5puuGxWFlWFbqB8Mk+nEotvbh
+GAsOWnGEBBX2gdvHGHbnnzywjl7pixOvVMPTvb+XY3r1u1ZIWizhxbE8cphzIuS/n4baKBpbkHL
csqMmBSQpLoHAPbUYpW4UVWElGwVkjb1oCRC1xRUjtsvCzBnH/CJij/58fnM3qA1fsQkcW0YDNwN
8dseG0Y7TTo2PzFx44V7UpLd50JAkpkLSk4UyVrM9apzy0ppIJ0QuT2bNuQ7+4ABq6iF8Ge0vlHF
VzFrokV0qJIKrZCDCbDJGuPvA4eY8iswBMD/0p+H3PsDGuJbDHViIiXu/Pd+bHgCTBkPNa8OAaiC
rpEbPANmRTeC2zKG5BxSu9SME4UcUg02S9k7205hHJrLGyL3/drByn4c9wcpcWHpez37zU3JSxuu
kp6H3dVD/yJoxfOmPIlHPqho4WNLV88GwsvRatCNHuPlR4L5SYpbPEO+yWYp6NWk+ELNqQRJza41
/pU7MIa9bwo1obllE0mdnX9vxUatOzEDYDkCDkzQB8vaznt0TWLhE25SWxrALCbGO83bxqlrxAy6
q+S/Muk3XDeh/31Otfc99bAT5XTTuYzqyFiPkGDwTAB2pnyKxSrN4Gj5taK/KGxnNOPpPRmOVK8r
JAAG4Ya64KrlP100HeOvjMhsi8XixsVrRFQZ7hsm1jKTfoQz94cRorm6exsZZ4StKZgUIrv4tMGg
rds8SSZuGluspXBk9rHx4Brn02w+XH14kX2kk0BT9957MDS4F0YqbYmEatMC/3HsdOif7oETCLwy
MmGoQJAK8APXrjlaKbyHjQm343xjNMJoXFRVz7yE/l8FlJBK1ZYCA7uWZY0iiqZ/3sc9rLE9N2Re
RzSviWmMA7xi9vFktCM+LLW9EDWiPcTE3RFV+KkkTZXA5yAd2vakpTr31GSAn+4U7uTC6Htxnood
5RP1hiIHkK5IuY2JraoJVggeZVju4Zg5SwlN8f5Aq5wvoDOxgkVpQ2O1T4EvvP72Nvj1iqKq9uEp
xjnukXU10yxdafwe56qsfJ8VhHmm1DWNrbgGh4VAWXX7fp1TcY9iNiHaEkiW7LANXU0Lr41R4CBj
T7Xi5mEZyjHlR1u7wjLKTnv0e1OOEh5CJTPGd8Xt4REc91FJQIlpPS/UkbpeE7uNF/IUn38oENlX
7HckK5nj1wwFg35lOCflnq4wbITX2dQTeWhsEdXxK5Z5Xdny318PlswHzu9iczp5WLSXn6t42efX
2O8Kon1rd+fvqfDv8XaFZ71XMDA9RstUmIYt5nmVML5lQ7bslFfoWxtNhiLdJWxJlkoPp8BFuipz
iR7Fq4G9cTGZi0nyoMda4FNjM9Vn7SwuEO4rzI5f6PNHS7Srgl9n/t3sy9CiQVcuGlis/2V2DHqh
4vLe1dd5Rym638VO5nKYdc+dSScHnENzlf2cKxTMYH33bBnkV+6SIIBraHGeojhp8IklzjdkhEMH
VINZd8u5nk6FyiPQQielGdmqAMCIlB7ZJ+mLnTPX6ESt3Dx2Wy/fPtZ/AgsoPv7KHQTf45kNbRpR
SF3b0i5XsiiFz8so4pigTmGTEhZmsvvg66uCbkL8k/BsZxC+9jWf2HuX/eItfAffzbMuSja6uDtk
6d9DI5jp560KtKle32oo/EOtxz/S8XVOdij2njyKZMiYhVXAIYfYX2g5bVj8KpmPFo4aCAKrhCbZ
c0JDwZ9xF2pbr7oMet56fnRYpbPYHJ3RjC2e9m3ZpepVnQpKsOpI3plWXjmN0YYBiPN9bv7As7Wq
wBl9egb22OQEhxFEMDbMXlmSZMS0Ry4AfSXX39fjx93KHjmiRjGFX0l+1HcQ4RerK2yBUR0v/DFi
AfdY+rudhYcymXJPFma+v+7uLoU3t6q8BqntihyOs+tAzUNvjvNf0Uro3VaZ5y4im/KszKvtWWja
YMpVCGYNKmlaYIoqoCa120g/0NX55BOolzf4Zs0+/r7p01I7qL+9/Xt/jgcK8vEISkFEkGbXokcO
AKRZPzhUDGufuh8e7aUKZiRCcyHayk7y8/lSTad0AwIpcMzwFPeKXnxTXTtMBbGa43/l2QWWof3V
Cr8/1VBAHRCwc+VviHYzgWVeEVgIOERKZH9XYy07RaiFCb4+5JshGOyV7x/2jH/XslMxNBzsc5GY
fOM3KUd5Ma4qG2rrpDcQ01tRgms25gSoHmdHP6R0dLFeBgvbHEIHzhsg0Ow/p6UpFPqIcox8s5Nf
MskIsWdc5JqLvM7X8XiaD4CY0+lJCTFM/D3urRbgwjKtjr+4G5hJygzgB2fG1rNGj6gxfx9Noy1a
i07AWjFvJW0shfmIb5W9MBiSM+d8Th6H4G0CQAalx+qyUJC99pYFeUdG7EfR/fUMqUGqwJslfwUT
vicJzd/MdiRGzQvTID4ZAZb+Br0IzaL+4fv43ErfPPTn9cLNjLWvQjOxQU6XilYuNBSsSJyi2fAk
TkntNO+mTqKaW+GYZVOYlrC4u7FFMKCHS6lU4FPne62u09WSaqlqjDOgXyCTgAolDo4t5wYwHrtV
kfy4fH3+9a+WJl73BdS8cDylstQMax9TQE4dIPi1D0w4sxxtl7STNpiN5fJzPkmAGaUR64NPOBnm
eqVpbNbEu1NkARJtV7g4G+UcVJf9HfnCcimRkqGHsJHeTIATCXMyMk+zfkgh1xdU76tOhXA20Nrb
eCv4jZB6a6M6APEw5lMTGT6Ft/Rdz58DpCrWxHlyrTElPJDuQ32i6eAfuFXfqfteVqFHVwNlH09p
HS/SdGN6fFnniw9Kb/xT8r2YCuOvSLgdxK2qENlMXvlY3N/c42DiHgCEtymesrsJm465n45YTftb
H6/7I/omPdatW3f8pQirSNgaRMrdYWCk8JxmPFRoM7sdc2f96Lj0uatMXZKQQfqiudxEkM6TPWzO
wrEKtKkD4Z7vb2BZTgoX3xIZEFM5sa/Q46bCxb2WnL5fm/Xgjrw98Dtb1VFsUtDmvd+e9H3CGa21
HBcdTixvTQd7R6rMbAJBgOmsiSyHpf9z8MnAYwTPEHFKJ2M6quTy8ys8aZXz62WBKV9PhONFk0HH
ShEytp3QaJNS9d7rdgZU4/XTX+pcKJdh2jD7x98Yjbet0W/8LSgwppSroEN7FTjtQ4VU0g+MgXHF
nyb2SWqqD8P4TAJD4ldjwrDu7q8JWMw99cWvb9bbLrww/srDhM0Cz8a6sadDL3Uv99oFls6Yy57k
vAGXf/MAph1lvGuPoeTHW+AF2YmTz6566PJq9AYv7eo3l/gdXyKJ3A51yvao9YVzHPCfQFtsJLwV
8SMZAqUY5NQUf6NsgCqJaqp/AAw8m48REj00mTp5IbtO0yUdx47tnEVjf4v6fr3qR0khSAa019Q4
ti7Rv7WYJ7Ty6BHhDtNIE00TyeUmFaHUM1IzJgdgvDDdoMRLXol1AWXnAe3EYjcrraSA/h+cbGT6
/JnM+7G6SmdKnwKVmNdQ2ehUjZK764PgIkfmkpXpdgciEXxtGGHNuiq8gGZASsfvl7iNvotdHF/Q
mk+GlWHCnXvO8SxEfO3nIN24Hd/TTvlgiDavbJW+EJoGcHFEEeGbnOHyjZI4Ko8IGbSUHAIdqWZH
Q4dkoyPJTaRQdkLWf3SclxVH89MdZWoqqHbRCkOFHHEMzHyRNpWA0WSsEG55cNsvsYTuTM44GL7c
j4k6ob0+Mxq43fqwTel5Zv/LmSoHElsgaW6wWwNMVbTMKnIswHh8B+KDtZoY6T65pFWOcb8X1oer
1PSX9FD7QjvOnzmo54qQROAINk+lNT7NUN7vATRy7FGk4p48ecIohf5xYxTY4fYn/X/1QOGsLpXv
PQSlbURKSIo49Sv3zV5m8tjzddZKPzQhkOjn0dfzfha3lsH62HWRAIj2SHzQ5r5y/pSm9Ey/jTrN
oYfbvuGywCCJMPZmpDlyM1sF1QYON8MVOE9GMjUjVqoylBxcNAn7lq+3UilTghfs2ZG23gXgruir
Q8S5Ym2VH8XFPRR+OYCYmVIpy/PKPcMPLx675gwYVleIS4+13lD4viCbA8wiSuXFX8eOv5BI7BOo
7GwxXNcArOtZ944HNbnDO5uJPoY3TfH1avWJ0YUvOJekarnMN+p4ysdUxdhsl7WAIPq+34SuZmdv
BFA+6tAFpkhbvgiFzlooTfEwzMyv2KPCcwew8bDxQSsYF7mA2To5r3xi4et9VnwCTf6J4h+dZ+w7
FdunLTV8WcHwWW4JPu9aWCYfmJbrG1Pv3HMR+exxZG/hUSrY9+VJDleNBo0WtTxHfAJ1e31vw4xE
93SFpifZqzGlPWBJXdAwpxYPRsyy07juh4Jqxuvw5/lFezRVZHT1rOTQigGxXg3IxItzDHbPlqhg
/iGVzWVzbaOySmcS+mTQkQp3NQVd8etFKV0rAq/GXQPVNC+BmKNnHdbHA35Zh/7RjBVZwrooFlCn
KWJ0a0eU724DN9xpvPRjd2DgNvVwlyoqIcFJaFvdjwXWIn36Ba401EfrIu/KMb1uZzbGl2Vq/AK5
Rd8Cv7r135QWWzy/NrTdb2S9ut9w/9jRK5IpmJ8X8t0A2NFTvfyCYk2h0Dnr8/9d7oboxg0ml2+D
dXLLBb8VqdkKKpfL33GVTqxFUd68JnFuTlhqww7MPBic5ECkXZjP9RhFvCRqNbSQIsHULFyvfbUJ
tqdokk4IYvraxbIdsQJ9PlgvSL58wiad3zfkrhobF/rPE8pBFct2iT5fcNoFkEo16xm7kC61sjCh
C6JnP1VqgpY/++3LON54erKawokvGsqy1IVTNqujLwsm97Vle6Cwg8BkllgT5+GKX0Ynqsscn0Qf
uQkJ3i6aXZ+fLTPIvq9sT5isyMRwEIunYXnt7FWewVEBMV2l4N7MyA9lkfRkRiXC7udcqAll/a3l
irJQMCSdbqNW1wLuAl1/eFRpOjfD2QCeVjXcQVYLI59NSIX2IS5jsCnKOiKKQfS8CD3A5NwUHtvh
2hWkCTlQDdYl/HbjI+VXH/vmJ9fPREdmSPDdBgLsTYH4U0/I1SFS6aqI6hiZ8FERVNmypMsUvkZD
OPvUhrnkyMHAQZsfwTcdUctQox0a455ltOWzqd6oJxqEgtWPToHj79GggHiyc/atgvzsyvYamJDA
dZ/+aHSfbcNx6xJln835W3qQl8vH1sL0TvguYKvyeVm0TrVgHFEps9FzyCvJlKU8OTBaC03HYruW
QOT6AHn+9Jj8aY7NhQEuzl+1puW5qbGjQ3Ybv5NEVCTtYmemuqJ/3zE2Drfrf3pXTrylKTz1LUyx
uIV/FSvk04wJFhTaNh4UBjvba9ZTAzeAibp5osGNl/yyFRAMmBVnO5B73KdlPpEUyd2hcDBqzwij
1JUfj9um+hYCRRIPuqcGObFn3MVvipr+vwSj4iOUn7VjbRUOqDFlIDMWXbTvg+LIu39uyxxepSKw
V2835z0/bTv1bbxdBrZ2r/+p2zf2FIvsius8q5GSGBCDnBpy+0d6sVErtnyiWY28nD1YyjV8GBlq
x+U0xRpnpiq04VqTQRdDLwcloDV9D7/2PVTfPM3rZWVZY9gJlhfqTTacDn21zWCAp5RUrOZqfFWN
YRkk27JRYoWtRMYKRfjR7b6Fhk8xeRnMtEqRsXBU4ZCpWJBrJ8TqF8FZul9U4/7umzt5i7yEf/Kr
bzf9IowfsMSYtlaxkyBW+V/9sZkRDMvRuSlx2sLFHLDhkKsUV6ofaimEpXGLHwA5AeAXciYAEthM
RDgV34L4byly6QnZY34dk7xjd382K79aPrgv0TEQza7nKkR6cZLsWYBXFV3rXVkEZiJJfXPwe9d9
wuehgMJGJ85UKPBTS0VhIvu5pnIk48xVwwEJCkpMISnf6kgY1hlkWC4qXZl5M8B7/4AFrrNGjGPt
g8JzcMWextP9Lctn+5zcAHmvLe+/c/jpyee7xUetOh3AZ17MFGxb5/VzQBjN9Q6AlqWQutsBbG55
MDBtSo+6O3Xve4PasEE8lqzxoRwqNYG13VE3mpjklnl8DtKWTq5jgnowgtmT7OctXMB902rYfh9O
E46zuXdOw8hOAZ4QHx1a/jatiUO406O1zUeDQuVR3QzKoPheiU6Sratv/oplp8L6o9Ih9XGC8uLd
mksbg9HEStaAXzyvQkg9JEIPxEiQ9kD3drL1hfEyMNjead8kE0qcToE6s4qyXhL/H7kP2kATD1rJ
rJrNTkXpeptFi5p8rQ/3P+fLacpJ9tO69v8MvQV0ugW45QQ9GbFxMXzpgK0qjCyNGu0zpyIdAlY8
XqvBNr3n9dG1zChVs+Q5dvtwHyRaephefE/RTEm3fJK52wDwizluvvmPKeQjqxnk21AMB2Me17F/
uW/NNBr1IMCPPMsEw/o2WhHkth0nRZIhRkC1knRtqLAg7vbGiXa/2oK52G3xIj0B3nyVlywtmePX
hxZod3BDkNnwaGrwZZnVPDrPLySr107La4LcI/vveKfZ7Fo+QevsqsZMAneu3OW1PH54+9xHIMBg
mkp3yjkEYfhT9X3VzwRtAWIFYjhWpCRQeLoa7nqjo8tnur9m8Kl2/ZFPkR5A4quLjsNQ4jxMQuay
TUOdq4Zp5TFAs2PWVcQU3Z2hxUh03jQ15xWFw1iVAe/QXY7DbNklEWW/U9+6cADxr0XeEITZgxbi
7Ah/MQdhdnUxoOA7XNKoOnp2EDgU7dC3TltFqc57i0BinoTxvTNpsCqPV/Jt5tP6mmWSs6cpPo4O
bJgu5OTQXfeJ80xbsPj1jfPv3FikyPEGS8dIvo99wgBdiCQ4rmi3MWgHdQWfIr2Zu6a37dlrXHKT
tnhE62XZFe4XcCrVC0Un0u1eqGOCKwngkliPwK8nvfWw0ouy8Ws+zgoX07OomHb127HRUG4msUdE
jbcjF3IUk8nry0GRpF//BLAOteSPy7ehAenpy1Rfyyb9kPzdFjYYeMgD1itBHkpzB2a1cZUgDjWt
A38rX+CqOufhPoatrTrtIcQY/5Z86SqRmejbk2m9yXemCGgLCPVgJ3klvHhC9U2H6tqdXex1+gnU
7015XeQWeO5Q2bgzL6a8OQy06mbBaw2r15MFrtSGehnT4Hb0XMTmsDgMSd6lPIpJb989ciZFVZFf
tVswfmB5WWiR3/pKbPjlT9lYeoayK0rL3cKmvlQ6mOMUJTzA1sV3mRqjrLpDZrpZPdw9ORqmLXZe
Vd97K5vNtHT7raUBPvQtcDeaIldGMr/sQyhm9zx4h2aUDHOecG+GA1OvSVZjgF+YvMiV4FhZ3mRz
UaQ1UaDH4WCyn3QdQNKfi6hC8OJSqwGMmpnnSwzJgqdwfd8AjR9uIhPEkpYOBEA9a2ORyErUX40I
DuHb2qGC4BfHgf9K+SschoL5cIZPPn+A0VPR3fyVS5V4KmoBP3OvDh54Rn59S8hJh+vdbEimjVVm
3rpIxu8OyKve3qnR3xAio6tbUm3HN1PAk6+KYW8ocm9QqFnOklsUlHF6aHB2M/DE3DjpBsi8nenl
AFesIxz4h0mw6rjlocZuraDYv6SpoVEEahW72RFU5sAvhOYqUGAXfgxewe+XOAjoAfvvEYBosjva
5bJ19VxeOEVW69BgkKQpdihaxj92vrX5OUkcMiq3sGd6fWDsSO8X5RSXYLkmKEUPQ1ZljpJ44bmG
8L5Dm31weADWLUonncWfPOHMX1/SA2EcmWj6BhiWN/COanvqPUOy9BljswX6QclZOgyvT9e1ftlb
XbTW9jGcLJBbfWOqdhipxC8y2jwkMDSBiOluto4gY1Ij+92dI/EB7oMK7d1GzgTD6QCsxpvrh1AE
MBirVmGbSZzuSMXHCw8MNmTQSr5yVQCWE8JpNyO/vRfy6Op/Hp/g6tmCHH+nJL/iGDkFXcJWtlFl
lmmMjOR6JWUsqcFrGYj7pfQupARB1G5CXP2zQvC9X5ifiT4ABxBYkEXRhUzhRBMCgklNxeyXxbDy
7l626Ap+R5E+zkLgOEoTVr31xIuC7pGIaVuYW25vZV99FFo85Xw5B4kc6sWOb+iAFhXUg+f2XQi4
wPpha8TasLYdDR1mUs1iMizyqSOLN9XLT4KklmKL2Rg2PVHnkxATLjUK94t+FkFO/zTN/NqCEwf7
0uVCJZKx3C6OxFUUNTqNY+NPzCviOhflaEYiZcJr429XS+XyeD8AphiOzcJL1QK510mEJBvFz2nC
AgeWJRymQat9dwxHKjDrNa7PsbdHWAU7ejPn8BZNE71H3TGJIY7OobkhfmyoAKtAwwQ7vtzB1H9F
O2oOVw4WcZmJV9UqVXIitGSBtIIXKZfhtt3wog/osYDFwLf7PJ25H9y4oBSGbPZHEVqhLCS9VOyZ
12BmIC1JzmSNFwdr/LA3e14u5CSxvbK+wwAs8u++Zlo/RRg5LnqTL19YwSr39T0i0+0A5pbWza5T
HWd7gl9CfhkAhGeFnyG+wy3cVQ10Ytcp43kplSwwnWhYQ/7wRgFz5CPo/WYq/tkZrQjs159ZTDTe
2X+iseGLFuUuPMgddJz7abAl5IuA0UbpR5DXUAtZOD6/l68xNK1j6gYY2+1dJQPoYSUnAaxOCogU
rdwIE9525ousCzmenDvO0eFOvq7v9NMzRHdmqgB2OWsVloqn6CyjwuDIqYiOWuOcNxApxIstqCVD
uEMGGwGXM6rKDaxI2fwhqf0YWhCsBdasoHgQ8toGM8xnjFOpsa+h45QteCL0/v9JgXl+GuqvDcuG
Iw8w+GO0b1jZJMw2Zx4W9IIMyi0O7gyFFfsz66+JbmJc756SbOFirCojJTI52Bvm2B2lPTFOMJU8
ZltxcchtGM1e2NywEQyiMRqbR7rDPKRs4rYdzRHQfMqa5oIXT3hFsHEv5qaZop8Xs0KJN9r3x09t
a6iZJxXk0jS1ZuTNVJMiGIPhTGe7RHkTkGw4g7+cLVgaBNHQkXc2U4iDaDhQDHBqR+3VPoz96iWo
zC+3qJgQypmosITmwHg6GYZlepTlJnn+1XPmWOdJOCTmpc6Mlg2H/YMXgS5xPSDmzgBwONRMMfvV
GXf3ASlRk9BQqYgefJlrs/G8CrEoLKLVHXkQ7ZpChTKg5Xej7G1hQ7rWQ2x81pKs9QycWCn1SE9M
kudEKhi+RiCGUWdJVp+R+WVbJV0qROKGGh2NV6HBdV5AbMf0MROvc26Xf69q6ru2BJwQp19TQONe
UeTlMprE2isLen8Utmx8CxWr54fQHMmiqbiI6A7liKLvQ3YQE8siUsrfblC0i3QKaFsGcaX3VsrN
iJ4JBgtIMoBxiBNykvChPrIed4xmhjjSEF1e1Pnf1zNd3LDSPbAZHu/EuRmlH7Q+2RrfF294epLK
S7oMowyfc+JA5sxKw/7OVkdf0BD+F5+Noca1vV0zXQ/T+X2zloGI0OIYpmES0EqtRi9ug8kpYlqo
iWF1/X772lc+193iAD/v+lMfRN4r60nThJJDaxmJKwbDyOYBrNcwahkWmuih7GwzYV7rZ0F7D+mV
yGVt2VfVsIDwtlVjHCCdz//Nfx+7agoYpVbZ/jQrdpsBRlbfNCz23gxcCHcY9LEc3ASMOGYApGAd
Xo6pKi5JqKc25IrqvImA8y+Ri87FlGeFRd2+mxFvrTP3+RTMTf0A7v1588K1nAV7lohQ4r5P/xFI
uslGUlnXWYnvWQg/0RP52VPwChfnt5Ih2R5/gxmmSZNUBoOGE+2BIr8vblilKBAqmD+UBwa2i1B5
WX33sytAOTIeQTEdf4SjrgrsesiSZ7+yQ46ADXCD1QxDPDzA22AUa48gwiCRM/he5ayUClPJjHTO
uluA+DCSzKSxxuvhA8m8DEedAaIxef6f5slaJp/LkgLKg1zXhEnjSyO3mI0Jfj675P/BwMEeJa4F
z9YkYS1RP6m119+FsSRE06iDAtTFXCz/Clmub2o/9mZo3q5SzO/6asOwgT+sJQawgRDNmdspOS+Z
XxFwlxEHmJxPQe0G+9i9RuAxCcuS6t/+w+hmiKM2feKII75hoLJXjC/jvdj4pi/t9FBS4/6owkcB
9v1Na67hvNfuQti4Aue/eHEd7LmuUfVg3ACvRxAkKTHlF4Fn5MJ8vnr7sQ773IFxZ4XUI7DNn2PK
ruq3tGQJueeHUo9nYz+BeaqAiaLhxEbaVxPu2/egC/S2KloLmklRdtt3z2D6c0Qi1ozwecvG8oAM
0x7jrmarpwEb2pU5iFgxSnsGUwEinODql/4Tnd7u/zc8o/wX/lHXVqb4gbc2UMy4WE1+Tif66TWL
zr/MLtSlGXlDJDBjeQ4N18YCkMesDaf3dl/knerfBgGLRPTxW/olid56Wnu443Pjq7+VkW1NoBWB
bdio5VnWJMIhmZmu+NFg6GXGDokFZvuW2bnIViW1tLtjmsyzzw0E1IIDwYdQzHrnENpt90JjQfqD
vhxUvhG+TCglPaoSivBGvX4H5KmDRA19+yydPbcID9ZMDCch/fp2IeHUx+wEI7Smeu2D7i2Fu2d1
BDqxs86HIklV9HXnM3ZJy/6YAek3zQ+0VCo3X2JvdRk7zEOepwwRLPJG33brrJVH0eUp2CV9dRc2
8WLMYdo0LLEntHd2cXCncX6/2/FBOqIwTA4ihluqFv6jnnSVbgeRbUhErNnafBZPg1UlWDjmZjVm
aYT6866ib7locHHivEMJyQhbF2ZdhpFDJeX4Kfil+8TFP4PMv3x/YzfucXIzDkcHNSJT6vFvynSb
L8L69SRBmxW16sYQjVZa6GXryGrs15+2jP63fehiWXtQpuGbPP15hLy28qODI6fcsI5dwnsVI4q9
y2ylSu/Hg2LE6+xtKtcrIloiBUaw+eodSM6JfDgi4rSJddDZHbjPhKkqiTD1A3kcZuFvp52zap8r
1WoBflDSA+NN6PbjXXkb49Q4j8a9X605JE55iA7+tPuZIY0aZIXWI+zqPNlINelXiTk5aolnh0Zt
iwbcRkwrH8H/zI66X0axgLA3Wdg15pb7WUhyoPkO4pd7gEWcA0qqCdIp9Y84qdDw4w42WTuxTo/P
WhUj9KywagjkNkvRBuvxlsV3Ncg7qBvXjXsTmXp0WRH11w8S9/SPJDTXi2iof17FHRx23kCON9an
290KxTzCYxYcCLWZ6GSL09Kgnb7OxNhKiAq+E3y/0f8F54MBfvXWBbCFcIdin4krQRIkLc5YYsJ5
P4nIOKo8OZvt61fcRvPMmKwg24Zz3EVsXI4E5hZLzUMAW1EBs5xD31hQ57BqK/eqmE2S8ir2stMj
GrMSyg8K/MhCnEi7H3PI6TW44rajLwHgwp82f2HZaj4cTcQS74arOk9vTc/F452/tvFFqczXnh9K
ddLRlQZ8XIImCs2IWSb9KCP/wBJY/fdGKRHfJ2Gnt8yVhHytIbsXEVOBh8u04juHKQCyoFDJSyC+
XOdDAkheIlkPIu8S1/yWj6sEkPwR1RCDRRCM4ckaY+uVTw07XjqcblOOn/BcsTvvbzPphk0fE2Mi
4/6nty4geMsbTKwhH3kPM6aTb8QxCz1ootOfOwWJF1BqaXuO1MYseOPZTnvqKYjMApAHL2UPmvSV
EO33q3dRFkqgSWpQ7rNpGEdPMTYOsCnYuWioJs3eWLrpxkI+e+Q26/1FougK4Iv3SYj/mGDO0UDS
OL/zhjOar9ar9QEaMRoAaKvw/YqYj8fMH/I2bPIRHEpB/Y9LSbJhD/kbaUdsUOnl8IiKYEBMjSkT
cP3l25tF6rgFxvp8czUUyxyVwUVeEl6jp/8lkzhzjvldRYMLEz9RKJEHGCLqWLqOuL0JaY4wW4kZ
FDzSqVCZIR4ufuQF7VAdBWG3Pb0EURpb1i5YjucappJYW4TD7zRaOWthWIWJdwz/5Zxv4U1Dimxt
KJb8B6EJSwrTzR0maJHYb8ds0gs9MDs/MAT+/5iuC1zJ+s+QrshaPj4H+2Fb2hcszLqoai7e5Nhq
cyDhTKAzQjEWSkdaJvjUnG4U63MTUYBs1OVw61Eu8GmSH138IdS8t7Ndr9+gADbd6eatwPe9EbrY
KbQXJ2f8eGTUVun+oam8
`protect end_protected
