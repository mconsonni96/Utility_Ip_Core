`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
MF5ioD4c8VgB+qQWL7qjTZQbJhO0KPd8nuNsg88zyuoMWReK+xlVv0ZIIyB6nthC/1Vz1ObArP8C
+ByCBPER5rG0VnQG15B+e3LhDrYih2gNEiUBAaorUXah1m0cHFdKYQ/SJ5TwTfbtrFBrrvANFJnj
CxepyKWZwtYCN1IUGdW7+ClqaxV9INOHuNscdoJuEnF/0Tc79iqZEenlt+8or3VCat/2rO4jJkR6
+epBx2xFhrB9a14dhaKTqxcnCt6czmlPoIFQQFKnJYQBy5DSMJWPyd8PYjDVxwt8Fq63Keqo21qv
6iJ+LRewaKMWAk6RXOguAQs+Fwjg3/Wb0PTAsQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="RsdXqm0LBwpicoiYG5MVftf/kauqZ3T1y3+uj7pt4v4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8592)
`protect data_block
+yhROyVMdDwrS6w86o/HD63SncoG81EqryIj1iXufO6gzm//kmr/7FV5ZQXMY6CoNtprU3aIXKpt
pAaVxan03IDxLaCbIXv58PPzbyT8BGmWcARDaMb4asRbOeforXW+9X1euisM8IwH7qvX+JtzIvyB
3sYrpQ4ATVU5IniYU+aD4hzxzmUT6F/aCrsfN/DrcSaa2Qa4mh7BuncE5tIOB29yuatjAPFAbFQr
RlQsfako4slDHDrBZLfPC0Y697oxZxaZ+/yaNcq/81seg/jc1uDypTiRBAcescO+DO1gsfFjHphA
C88lTspKKB/qmVPf5SynOJngUIV9mGDEvYhAovADeU9xvhGdEzbQdceRj08VzBsjVYt0GFoonoPB
eKKnSZYxf/ekxdLgPIdEe+NlOL9UAQT29xmoo9xbtw5xQBA0xvsc+XfZKGO/4xEs3rigopaqqJV/
ybbGAQww5yPIAUeZzYyLd8YncLsG0r0RBMwhfgFlgLBFuh6wTkg6aQ6J5ImecXSxiBmtpoJ14d43
PjZbC6nzutIV717yhbzPlRSM6qSkrylGHEy0svmaOERmDm90IviYWTFbgnTt01Wfd3VO3RR6vmMs
N1Oa3x83qmOxxTKnjzqhB719I0TSu4sEfTYsDpjdCE+mCPai+VQ0BFUYdhsJQ6BAcs4gNOwn6U/3
xL7ue3MhujCMab4uNMsRuboSw4kVtZV1TfDphy7qxgEnLkLQKg4Uz3n3qqe+ROPZdYKgCKoGBq9q
7dpPDfBndbBZe4wiEIo7oZQEim+QFozyxEbJFFNCf/U4x1VNmCV4OpStrp32tlXjJbVsV4hamSe+
pfu4sFgysFrM2JRCF/u6Pq/4/tjE1OYH5qs7vbcmIFbilGgWVb2wNhNZjtoNegJ1rrLvs4u8PN6M
v4ixEMhIBtb/Gs0oVRx9/qa4Zt5Y5DDnkGo+QFcdZyO/WS+hv5wq5KRIOGvYiJinNACFru68kYVW
OhXpCMCp2LvAvaMLcj1ByQeXKEWrScRrYu2kIknr6By8xm7dafRxydeBURyGo0vqOkFWKVrmDrKj
gCKtlztRHNez5XBIyKaBUhMX6FJYq8nPWdk2OvXwJ8GGECjlEU1FiXGeq2sZRyWc1njWWsd+Clje
iuOx56AB49GsARpN/5kDduWGtAgM32UHPnzP9RKXfx2meVi816BhnkqFsry0IDmhCJ3MC+702lhH
crXTVsm+kJQ4A98j/HGCOrO/ZIUVB+V+5wyUlNBL70qOFNf3fH2Byz2QGmrVJAPi9lUlTjcfoIv2
z11XB9112OadVQWgg6kiv8+n/K4tSWNgI+9jf6nf2Gh140jP3T1rRie1hiFXrVFrVQGFs50HZz8Q
J9rArId71t+KsgS7lHpUdvDYSVh2RO14CIBDd+QRhY8VwN8gHpJB9AEsMaH5mP8NOmSDNV9qBBAB
sGzYEvoHduw2SkiD2Bhdp/bBismQ85+ByqWaXYiC/Y5AhhYl+o856ccQBtiaFmcfGXyg/fL4GPyO
BFhIWCjGep2R3gtdJHEbKySgEf6mAJwFuqbzBQJ3xGzOganjxklTerov6KDnWEOsropx/GeZykhc
BjrmrEjLkfj7RAcrVHMCFRKXsKmrntVd/ORS0+hYl0H2RTGeGKFqh5NGJvHBmPF8hllyDsR7v8fL
PqOp9VoN/CX5XBb1qZ9yqQjUOH63RGP6goIJAKUfSsSWlh+zgbXTur7pMsqNOTzChRJ5EG1esa4W
4u4jzV/XHpXEVjk774kVrINQsQTfLtbastJ+5dT8256+OlkTMHAVPjB7uSStM34mEsiedL67G5nW
t8r3TngrFMzT5KvNHz+e6LKevgEOioYEYxDRQ99CnsWd1efRVN7XUUXXpwoOCHQ+YosZDAieOLv+
CmOFW0w1WiMGBIxCakG7DC/hIe3TC55SfoJgzRRiljIGEOKxwWKRA1cXmNq7ltw3DIeDWPjRq6vF
saE07YaPKKFI4PuTk78msGDyY38XuVVFOAw2P8rl5trmjRbW6ooRgDpvYNMcdrKcsVtZA7oOKo4J
WBSkYLddlk4WmZir4mV/rZNCPLznki4U7pUfxN2Lmy1FwerZoUsFbrg4PsNP5BccWHB5Q4+Kc7Xh
HtrZEdkc57myleC73EsWlNoLduPxdU9aYAoEOtXMVxe9BEeuqMdIYDj05vQEE+dHM/obmCZBKu2o
jO6LcG5crOIWLrpw5u08rC2AGGTzahAaRWVAkaVcp7PXTFwUAQGe7Hr+Qu1Z3V2K7TZ9DIuwY4Zi
II47VhTVq27W/c8Spvh7jzNdXFctSp1zuXkMLbbDev3iF+rB6/++vROGBc+IjsE5wvREABemR6TA
X9NpYoqt5tUvNDg8amwWXZzHKXbgKd5dMVn9kv4keam0W+gr0On2ojlc1Qck2hypu1kpXq9qq9t9
sK3BrvxeRva4Bd/31vuVtpLUxbDK1ThC2vfBdeP2gycPDl5Vz8JY7qwUeL4SbFKAH3L4Rshxerxe
3jLaCRtpqa5zPDjw2pDSx8YNXLiP+I+/jPetyY8LfGTjYMC/dse1WKtNPM8Ts6ZUsHmp5BZb/vkr
e4r1wThbJ52uXhuvsocO9w2pOtJGC/9k3wyuCwXj5fDX7amVosGiy98WsG1/pZLvjrACerR73kGY
N6bUGzmQ11Ayv11rUoUbbYqv/rbcp5FYGJhpFzScAT4cAQu7r88jxwY0NwXBVai4CNPTWB1b+osE
mnmGZU6Bi9IjgsSu4Pz2ox2KHOP5Yvn64FWMCifHL5Gv9TTgVNEDmNoc2ULc+EYiBa7yzzyL5U2I
15HO951+uXaouh1zWi/ZOnbl+z3l3e9MDG1esADNhFNkrY2rMBwaNGStzUcQkYyNlDJt8MBb5CJA
tW50DQbLCDzUwLa1nohAyaoRG1h7YXttNApoipZmIw0CIJ5jPtlTXnLoAEsCa1xGXzYzqIVi2vyg
SX7p0XF8pfpqhGDlrdtgwLmHgfgab0IRz4Q+ksHSwm3UXi7+HPN6T6PXcrMVSELpv5i+nSMF9kRE
bnTeJHtuYHb2mf0TGCLgYj8d0VLDRMwwiy6KsXD6d6nnpAQiXRmF7eEI/vmkzlH3YGcOpJ4l1Msr
S24Zkqn5fGiel04xKWged7EKfy4JvRnkbauEkPUs5yT2Gi38R8nWIDM1iUHQLX9nTwl5Utn1I4tc
kf3pKZWcbYzLCmtfocCySuHrrgG9KalA+ERGNEfxevVhhPruS+S0sifJf0cMHgEP2BieY26a7XLD
sbX0qPjzjp4Gus1a0sE2I6TLNeLTWk2Kf2St9V0qt1u7ejADGBq31FlK98LbzaQL6x9C4JMATfOT
MGNRM+8pz9ITU2g2pD+EArGpxRA3lc1PpU4S2lEKn5+7JoPQbqINmDzcLkjq0pADyioZ0up5rRs/
phVCb8a9Q1UL/jCmUcDng1Uhb6mirP5edJN58K4ngFIjenJykCS3k5Gx075IoHIvyvuwteWBtQ/L
W9Sq03uclhNn7h7kE1ppKTG13z7IP9BKxdtuEknk5+OTS1O5gmeNRVQc07deKm3zhV0drOkl2M1R
86cQJzjQxotLVyU9uQhXCEuFA3A0v827ktz70Bqtwk2gC32jvuKm6KjYXpgZDw/+RT+eUgfdjzHG
CnM7epVdDaci8WIjUHU8Qi/Sld2Wdq0JPAwDySgQQ0cMo2e5yUvl+r5y31xI5usa2TQHdz4vo8Ua
FM+6iL5PaGXH/cIPSXgeHVworKAxAmqLHD7ZvSJ9otkoxEjRbcoRNusowGq1ZpLGYX8BsXYlo/OT
TF38bgBvbN4N8lICDuEv8tI0adSM0jbQH562WnosDxd9uAHlvo/8htnw1rHnrpP/r1oWp7NCChr5
MJMODrszXsV91zJS4IDnegHcVQCGWDXwnECOWL61nORhlAHnbn8vBsmvjaQSoLXistYO1xudZKGK
HIU+9X3agBTsSR2DQvaHIwo1ukhenLGP9rLa1tjM3t/pfGMj70tGwD0xMCCnEHmOHTTIE6k46fcY
OMHvVw1hMD6eOij/hzOUSUzR/4ZwlAUpUqw2GVRfIQydjTwDBhSJgjvu8uLDwQTkqdXVmYwkOxPA
3eu1qKcT8XcKa8ZJQEvk3tldTqKe/djkrk3tour9agnsvPBiQxyZhqJ7e12BR7/xIp5/rJlOZwft
aiXp0a1v3m5Ff9RwchbrO5hiUNMHdy9bZYQZnk3NpnXiBaYP/Bx+XYhjNbDNqW+ZeMWy6KJUDqG3
8jXIsvQBYAPmfZIEsAIQVu+HrCz51jPJg12awJL/EejJmWQ2n7hq/MfmBeyjU5ejNM9hqgiduDwo
XfBoL2VABIEPvjZeeiIjl+JMeLWG5p7m96cSK2Jec+YGaqJBdxWYkY8Ur/xdFAeyQAFyHdz9o06e
RO/EhnsbbfONol4Qwkw/H0/Jb/jvc/iyXMqnLwlfy0IhsbcmEANypaDmwhLCklFIfD+RA+B3UQ8N
om70m653v0FqhmMCBXaf243d69oZuQvjTXKAaGICILwM0Jcer3nCan8TEbUWTaNerR85ZFGHFT9x
dG88C0vwOP5i4Yhl5vn8DgsHc7+IWuzn5a2T0gJ26NpJO9pU6JpLre+YtRDWXIrwWmsHUe/qBBXI
0WumcepSckkPjAfEVVylpWYKuOX1XQMhZvFEkcS3yNdPyEtnwtg0iF4PsZgX056st4ITeVmf2PvF
M8wJHaN0Wgi0iQ3DOVmZGRZ0RhqnVj2PrnI1XpIgRS5flh27wkQi/+mRCPp0xzWWQdBRpsqBbIjE
63v0ZPat4iY57URMJFO2ZWU9beDjRtHbAjen140osj6HqYBRvxsd0K+Bti0q4n75RVGq5BgEM2Ra
jU9lNJvOE/O9KDIhGKkdoXsG/OefSWakU6XNMoIE3yfUpTskxkRTg/ov/dKKXB4RR4LLBHIW9wQD
a9JGlakJ/Vf0VgeTjYGslzMVJjFYi5TTLMXnwH3uL8yfUulZQ6NF2R/GPEeG3CsA/Ths4PFcC58y
x1O6SQE072N5gt/zFyjl+Dp8SD9NMqAVIUnru4SIsMpcUv2ZKWBBcH2HSBzrXbkWFbjYUqQm+HgN
QwHpK6GUQRyRNYaZdpDgj2obPuDiJaw92ncKL8zABD6JUrzZu/A75VmpJKRFkLO10ECnOUkiareF
1y73WihjhxPoYfb91HYyCnVV2MV4zePhwdrSKyQrVd90kcfLaBY9TNUUlvA8VrKoycx7t5NMfZlU
0pGVczDzBJbPZTe9hklOJNpv0hqFpNAuillJTTGHccsyN6Hek/CTZhNT/BGzSdHfEgTco78sm52Z
7zWrMJnyMQNeSjYhjEEVzqQ43nc0ZV0tMWFrqxi/YUpsznl8fyStAYrT4m5bK9Bhk3IJKTsPZR+g
0UW4+3kt630MLlbV5LgjXjB5mu7/k6Z3G4QJgJozXG7215xziwI8qRFnffOi+M/hSr0p4nNDNwNe
DP/DD6NHWtuwaViZyUYyUV31kgv7amWyzpWMkfjfi01jixTQKGdlzhPG0bUDeSFcSpR9qskLkQ9Y
uIz+SGQ1/IV5P3xJaGntmE4TRdoxd29Ja73Q3TPW86CAdLaHErrxH35HBMAkt+cbDSfq95vFih5d
LuH6YRiubMf1WnodrWNhpL8K/rr1jy/303Ou8cc/YAfj/VyF21+Zp6pYqrLfTiRIhYuGqZ9UMiVz
7v2I5ZZDNNPdRJDTsB/0+RK2LsDO/+isHmJcBT9gPxSWmFN0MTnozg6Ay9dgsOIg1hG0DFZ8nP9j
oLQpWK9vVkZty02GPqZ3pJBNhX/9A2szBlFflPn/4h+OVzyre8DGNK5OEX0yTz+rXmYHFl+GhvMb
b3nRXGK2zRwQa1eEo0T1jsFwK2GMg/WjYaLVi0Ynfl2E52FrZw1JCHYIllla5XGc9w3vnj9bN1e3
6KGMifcEqz/w0nlspN0sAKc5pZma25N0mpA64TlF1ZOpB1oP67o0eErd2uRrVGYLuXMzZ0dlKkbU
O3d1ogoLGpBTzY6SyGasezSPu+NCDieENsNLBP+vY0GcOxKc3YvrVh3Alp12mOpZFh55epG/c+5L
4C9wDlgoOnNthDTRKwjocLoOTo1E0FAONlq/LVDJPtF0ZDVi7FTbEj2J4XvDylAzoH+UNNv1iO7C
OLzDIz5id7kCC4YYkZHL/m0D7a9WwKQir8qCr/E/eOaTASN7VQcfIrmli/45cMLQxQH2n5i9GgRX
5ijEYiZTs4LVzqROc40EifNRWj4191abjbRN0AOwD2rAiSlmix1xqhfZDetKD+2f36ZPXwXCv9v5
S8Wm6Z+8Wp0C25tZ2B+4J4YMd+YVvVida/fFYySEk+C199yGn9xGgkjWb8yOlorwNUleuNH8svNg
yBA/+RTuWkeqhlujDNZyDOEK9NVZkmytv+8nEWtZtikRrqYSKqlPwpEMbCOU1jGMjRAjbm6coIAD
WjHnU4v8uoRs66IzRJPOwTeR8LeiSujWCwzm8VJuyYU9pb947sIlQ0feOU6ydn9M0P37uyb/nVF/
qg0UBK9/SaELE8JXIDTILmN7juJYJLJr9/h0zUOEHLb6dmFuT1iIKZ+qYIgL/PUZUCqsEqcw4YY/
mgDWu8i417cI/am3SXDsNBd68z/8hgvQGnLjsKO5zlYiGfiMgtedPfI8dpRAfH4A91M4LZ329Sqn
rc/LoGdA+mP+Oi9NnPqp9TxWhcv5HAycHH15q9dERwHiS/rCi/WHJTcBiuZaCZxMeYENCRGivGkC
qEKyrS51gPJVybaMdxdDkE2HAlE203B/PV2jDKoN2jpBuHr33ixh1AFPyX4aSi2E4WNjM+gun5XV
CDD9REJl+efFKTlL/Wg+Pb0xl5my9LM6S6Cto+9XfzqETxZumA6hs2mqSufmnPJH1Bwxg6hqRQho
kMA+4A6i11HhUGFcVkMjvPId9jm/e6jLWjtv7Dx4FKxMkuqc3ppUHXHSPDT9WNFBO1HCgg0yxoCE
vR2edA+K+Ampx5WyLTGJkNuWhLV+GKo1cBXiPeasB2Zif0Nc417hN+J25sEHhpsivHgoit+pN8Rh
zDAseB6LZ/nTpvrT7wkjsyz2x3Kh5pO73sgodfFvXoT3YJQTSN0XSzEeqowyDkPCHdiKpNf7Fpev
+sxnCBaDtu2VXB4WlzMfUMi746b1a3QxgLAQk1Dr44b23jyRhXXQQ6xs18N00E9HQtVyz32N9mSu
NxCP4V4IINuw5m+7uClh8WWc64/4L5EfDCQlB2jIeLrBYJRmgf1/DNhAFm/hvVSPT8eAnVk+gQf+
TNFj588HV1whoa6f20mhjucK7UZXn5a1vDq4uKGgu7ILiIb1hHCbL5+82QAIKhQAJ0Onu/AIYRIk
vjxf2ogtmZrmKTcQudXLU/P9h10rJuQr42958pA+QI27M6MwqUZJ1R52dgwDzqzUunl9teocosWA
g421RBrND+2ixTSk/wJfSXa+f47jFIOsWfk0J+KQbbrtXjWluuAyIf9al/piS1R52BnXpveRZTii
K2i88q9YSNqEU7GZbEsPj85di4/T3Vyeh1k+65cd0VB+ZHtbmNZruzloCBeo+Cw/yc+6r5Zh8y6I
ELer+enR/rKRzyZ7xB0+6xhOVWWVy75c2NnERCaWcF5ZZuy+k8Q6P8qRQhEmZRVCzUZzNv6Tri1J
EEEuZPsZn5F0OP0YrRXdhOfIB1SNmYB7H4Fze/M5Mw+OShSqBlIM+VPAuQofbdmhdnGiQnZlJrBp
EgXyyLEn+fnVO0JPKDFRoW+tMU75TJlcyxLf2z8x0peB9RRPQYVNypBQoqVZ2OevuUmKEGodbnRu
nS9p4P8KgDRvn3WnJBZhP4u58evsY6r2oIrbYtmJY/wJlmQsdTZAe5Xp8bL11WLbOaYmODdEacAD
MLmfce0fO5gc+goofGv7TCsDqSHy2R66NaPjUsk8Fy6MCMGbLdUwd2NztaooBL2IUBju9njRQdRx
1Lw7R0+IEs1JdVercdFeWkzicMom4kf3RYmgxaQ+WJSxyz369tFYLaosz6o5xo1e+bClntTFCHgs
fr3WPS1zFNX2xhXhxEQZOCHCevvtn7PjK1HK42daow3fWZxYyn4SVIiFtHt3cUiTKF/Ohhhok6pP
ELbuHbE1yaiREeGBDK9qWOAg92dWnOSjJeNsIcjo1EPS88X15kK3XKcKtS4Ph6ZlzhRPn3QrV1Dt
12RKuYhfGR2gTgdXNCbIsKupKgw4PHmss8U8ldr1axMuQfNd/qeXOxqmxxbwoqlJ6i/vdDm9/DMU
aLR0SwxPfbpEBPKnnzHa4x3Sj/T4cm7/yM8+l3FDJ/QrgLk/N9F+wGOkw1fsXhnyMHWdnpLM59A5
MhH+C+HHepj/ngTcZqT0D7AC5SRLARHSBLqYXJuH2LDs52KhkGauNDD0PR2dmqpiiRMj7sN3wyeV
d3Y4THeqHwoOGrL5Oik0ax8z64/RyZ94BvGJMDRNHMk89sPMFg5LRGTwTTTXrgRWhegeYsXIYmo5
o1aosYSs4rjG9QrvJ6X8ZjVlWLdtt5QNzNHewE0qMYttj8FDXQrtfnt2z2xXdt88KV6pXnzlIzhN
A7xX4mrNFuZqifoHabD/VEJ1DC7AGgoNeZf2udiyNXwBzBQdLqtn18yqAaqSvJmr2xhTS+kR3Sen
6EV8HTCi2wAxzOIjd6j48Zk9JTkjlS/ClrEyAXoLQQCNZVW61fUcjd0NRdyZX03JYACq/StF+Ko1
HfX6jd626vGQKc0hIh4A1CgumesZrxUBoy3WS0NA+b7kG3cCkUobINrELQj0TGf67E8LXCFeJZUm
i1e0ybCLBfIc6NJL005dqfIq2eXrR7ooXD27gNlr3ky6KzIn8tedZMGv95nes/3FdzwJGvX8Kc65
fG2aJ8PUVXC8TfA5P1VkO5TM/KJHFEv96OPRbdDINqkVDnGOVJEVDA9Xh+uj8Chk909ojndLqofn
Zm9+m7cXjJtZNdpdyIKoWGvvykOXvSU8MVKOwcx1mwnowSOURe/4zHJgd1bHXL2D4UbZBOyCLWsZ
InIpixAp4+AasuxEBJqZrm6TblIyqPbnZDhxCrnjjbgJfyzSCyCcR3keQi00DjaqHNWgaYCV9FY3
kpUrzTo16tPS2amkoBqVTlB/BMM/fZrT/mbArJQ19e1/WVpKgv0LSadqWPpOswjj82aNRXjf6AvV
FSM4A5J8wabwBhjzPbIBNyydCK+pWZGH9yaCJt1rXbps1iLHmelSIGCIULHGrTaUUNyHtAZMPdHB
23cK2cmV9b5JlUpqOfvvyVN60tJaZtZdLKPvILhCqxyeChXEor63ckScKLOecxb0OAg391IaYm39
M56/D0dEMdJQWEcOQXBVwgIQLVpCkDINw7N3n/hGxsjDEP0ewTrojLCdKv+IO+rjehESMESHwqDz
5B7YofmSHBYui85QmdkQcFjuqN3f7HHYozTHgY5JlCuzeSTWrtVechEtCSvI/cC97G03ptl2x+gT
Tk44GToqPcj7uOSeCocP1q798Pb8smeJEUkz7aTcXK+1mkhiEGHvv1ws+2Ps9WdOV1WKaAnRuoWb
AFeuybUw1RRBKbVywVHsfXqXDHNbZ32MPj1de+4ADM9+c3B/sBhoZPw5idHxDkVC41p6iqmHoSzv
MEfFpM+iOdRfCUwpRjGqNkJntAIEhcCAGhbEpqLp26Ozx7bSP49k98PSoeIHsUQcSzjcscAOAf67
KbYlkNpyPTqejZNjFIfPJcDPnjnaQ4FgRdcX+fS2M0aq5yrzx1NFeZUp8D4lApdXj7ngVwuj3gLd
NCMmQbbJ4Fbr2utdanLh1Nn6RDutg9tLKvu3lJ2sMQATuJw0AEVpUOgSX1D5wBNXgzrdBUd/4s4e
V9kLMFfD7Jil/u0COlmnnTGsxEaZAPv2LtHQizdgaiXm2yQFXYNabTuwk0tBAuVoyh/XZXfkbhOP
MmgKUa2EFX0yiG5oxBUva5/t2Ef+EcLBgTJmMaPU8pAG4gzNlVVq2n0BLrYB2t9ZCzBZtn3/sOmY
69QVL21Bgdk+wVBdC86m0JczdfPmTapuSR1tefh28tpH0GAX6RfWWXzf1qLC2eZuGg2XXaDpwduF
mPq6hTzmLkA/wJNNg0RWjX81qEolWNa4Nis0yEdJKH2iV9rpY70ZFuuabQYrJifFycXun83JIGPS
C1L+Oh3hZuzrzQMRGz7rfLW8LgPfFqbyUTnIPvF9NSOOQLkHppE3ANfezXTWbkVGTS47w1TfTb8K
zD5yhmB1qa0SRNvpuv2ImchZUNvSpViq0uTbHm4DkbUNFbH6zTMTxHB03RjivaWNmIMTIHMDjBQy
OjBgMfsDOpNMU7DzlMHXnY1tmktrVIzcmtT72hmTr/BamsU0V3zRX2w+OAn2GBxyXKRUvFOfPYuQ
rlQO9P3dmUgX3IQua0XehBgNuVd2wDKd4jMmlCQLmY8mM4qPoGa332j7ubl1zP8YEb20ccA+6Zvv
MQIwRBykwSBOYquA1p5JqlkBh0ujcxWF1jieITIi9wcfOwYHbUAAgr02qBUsXVlocJKH5Dn+4VSr
O262igJLpIg5jG2PNPnM5yV+4zDoPYcfFq5R6HgHw7sYghA1j4ssyXAFAPgXYXdfDKhX1Ky7biAR
/fggDb4mOmwPYdSG3YV/amjU/e5nwTkbqFLvF15j5qPID9KJtges7P73DwYRoZQafeE9UVdUWdRF
+AALX5pXaqpxtOkoiGXkbZTYYQNB7awE4GMK0MtQi1Deg7EckZbPP70czgjOcd8VYcvY+p1M7e/X
JUefTYRDi8Ti9DFAu04J81QoFyoGrhQi5YZuBQpm7THze2/gXwMdxNgu3iqxqAWMR+Pftzqu+7V/
cptv2K/nBz2Dqp7dpP8EwTw5E6cFJmyS3JH9L5pMVR3M92JmkhF1Tb5GRM4oAjeXvbzuINLOEhi5
jU+wA+kargsxW3zoEyQe+OIevJmYLe8bVl3HUa3tb+rtvH1fVyok5pkbDvMrECSipD4A/wIArsqi
n0/BTsU8Z11JXzD/ozhTJ64wQuqjG+KbFZ8Z4ynKZjvooH/WQ+U4ZFw9EbpYwjWpx1vgr9c1u135
G/tdT+1ZEZFotKsYvBHO6pMO69BY4gSMdSq7ZcSobyPnk1a6GoLK0pN3i247w5pbdMZdmOt1RRVh
wzNwufFGdNjrVehEg18roQRHRdWW00bPz/zkNiuj2xqKpzBlWYSevIeyOlFkeo3IPVYOKTGs6cNg
9qMqVGubIUFuEe14yHCeVwM6JtdoEKcVsfd1hVzkZviDpzV3MDie76wnsv8SH3pNxHn87uljjsPC
CkUjgSrleBwKMeQjBHnLdl0pf7ZWhHM/Qi3vq7KB7Jr2StFjaCy+7tQ017KHqRgfM0O1jVxE1c9C
pIZl0EwG8OYokwDDt6sTekCvQFpMw1LB4PHdEmoYiMQayIUcB8eQ0sy6
`protect end_protected
