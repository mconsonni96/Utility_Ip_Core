`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
e5/jbZjDQmt97CrsRtm/wqSS4kO3decaPgWrKyOsLCzhbobp6JyMUCocLAtGn0Jkz10FqgUWqJIj
+YhYA0A87eV6nmKnjvfjB4GPkbnzRysbDBDnm4Vc5k1NTuDrgYh4sSeFH51ihyXsG4gbTK1L4Skv
lUmcMs+zB85HpWEUDcgeiBgDEjgapNZReMCBeNBGD8Z0jpEC/P1GtOJUJdagrl4FaUf78tZpJ4HT
Jlom2pCYnpLh8asYjw6UL2zBmlDHf7W5/qRnggKOBFLRjav5JlsN5Gf5reLuCK3ZIPTClcN1HDon
tVU8ZDwac+ZagijR8saygG7oMFExh2ZKbChbWg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="l3kZiJZZ5b/RBFSIY4fpMb6Sosl8h8inChZyfSbCbOo="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33552)
`protect data_block
WG6ZfX6/ukTaI0y64nykpJjuOMk+p9uoCuxC/pLdNprJH/+9Z8NUTz9G6ffF8JChADaIxHm8UD8u
MowXGKANdHM/F2ioAzczs5cdNwVzxe2j3ky+YoFNM1I/6NSaqF9vE1nOU7bSMXaI8NYAuqhM6zBl
GYz9FdGZ6tHQk2yGnH0VchUw8/6m/6b3yV9pdpTmNUbEae7KpeurA96jJWedD5Rd+f9U5eO0RAXV
pIrr95+7lfD327ZG7fvDEE3529erBzjQ5HIRH0nQVsVSYgKnTf9KDXDeJuD9d42LvPgWJ/WbhVeR
cq2u4bqjKpoytgagkE6nPVMiE5oP4fG1sohKip/a87FVjUJVwulQLg85dLL1QOY7HNN6y9h6sury
kgZHhpHYiVSgDTs3D8WLFip6MGA8hWXtOssz8E6Gyvmm5+Qux4bbto3PLPtQrUw6NGtGKjf51F+x
uGw5RDhhn0DfEostS7UHsgFPXrNHNu946QQoNuT03mxvt59JZQd23zyr0ezuukKwUNeueXtsRW3p
v6iLHgHbu9miI9BJ8uUfjAdyK6O24wSEyH99TeOar7m9vwh2Bp1tGo0DvCkrgN/JRuhvqdTJ4Cgm
X4QPaD9Yi/BITsiiolYbDFCUa+I2ewsYbrV7xK2WrDDCcjJU4gPp4SZtxgfKwDIzia07okwdn1CH
H0ufZvIcA6djhL59WWtmM/0zS78xo2koL6ViYLu7TinOzBFRLfycUudQ5kBjULOOhTgHPbuXVKnL
MTFJvJ3bEwGumpZi8SB7W+d8UoieWQYXc9ymFZzoI1WGJrfFoQ0bAIcajm6fDoNBjby8Ap9ju6ze
VhZB/abAiiKHPVABY9J/tQmrOJRJGktxfQZfa9VNrueZ+KXQZhMH2JPKkzHwafs1LNLIQV3sLfpT
CfVmI/IZYsFrK90DsJXD5Vrfla8ldEMslGomqC/X2DdcYJtG5/U1agBEV1404R8EJK+jfcvuqqAf
8axwpn2jaCHrZJeXPOwcYvQiGneTcfnEcKHvmp3zIgCxKeWDGmyKE8AdGKkeglGCScUHDE5aii/z
8orGSHGAmlf3mmFkJeqcJivGaIu7RBWsy4EywwThbycbE9OON5NhA6Ir8dFSTCwWJVD/I4RLazqB
JiGuLWdzfy6m1o3DwHErBmboZ88i25WxRG0+/KP+PPKie3sCAdq2CH5z9PLefStI1By7MKbAaxhh
Nn/0Eqy3ZVYHQNN6LtYomjFqscfnkK9cNuPwFbfgxrWjKcVeEqIiVUflx6rvS8Eeiy7Muc42+gS1
ii0UioQhkajToA+9YECUsKJLj23lLUXp/awOjrPl04pXeguk6ByBCZ6NLeZ62VvWfb9xZgA32tfE
Cla7dxvnNOhcUJ/VJMNjwJ70rQumR52WYs76ILh5V3587NQa0C/9n4dqw0E5RJNT58YQCEgOTLnL
f46pP+MUjUhODqsSqGVt2wxxnVlHCwhtX/b+k/3HE+mWaBFRfQmXD9j7F1zwFq4R2YHjQk+YDR2b
qJCXENEMW+KbNSXL0h/psze1xXsftJJEKTwd3j+f11garcQo/IUU5NNhizJm3wKF47I/xu70l4eI
U8mQXzos24RVl2Luf4k73Fuhqlr3c9ua3CsjiZwYkSGhVo56/eQ8o+u7w7OGaWyisNEwa5t0jwv1
VM/klhrR4DnIjW5JdxeJf9b30a5qz1wYLYIve+/RXyop+U3wC+lCtzc8uzQ5vHPEGUNZ50qAqKZi
ERm2W1U0Qiu36HFeyMmO2bI5DelGx6jMQ8k+QbxQyemBqSm8Imm3zkAqga6zyXgSB6jVYcPr67W7
dYk0FqfmAvxqFAk1h8DUGXPu60Td7QRY95r0mdjOv1xDRC0vDrEn25rRNRAm97a7hmyzqxlS1mXY
Qx/Db3wNsrEXHt/RR3ApvhGIOhsSylhNs9YpRd14D2Ms6VGBt732jE0u7SVNLkFvrKtK4V/d61uF
6ArrXbYHTOELwmCu1IgYqAjxtQsDMnuZUyMI9/a2EprTtG6OdtRbGcQkHkW0AsflLYESooF2lIEm
q/mx427jd0+YuVz3JzZMGV6FWyc7YPcDsKSYU1ws098MqGJgTgv2sztBH8TkrqH+csvtnULo5R1H
EskOBCjL2/USJGmtiiq4VwRWOlQvp3T2X58UoEnoYx+bjE5IfxlEDikt7F8DXH0kwLV5jcKlth+y
/YHVitTeDkugKiAX4jtYex30KSXjQxz6tt5uaL5NMdQBO9f69y5lb3nXXhkb2NXjxpc7zBwaaHIh
7rp94jnkkLqxmXF+f//zlM7sVD2fSR5ORAD1lh7idgBk8N4Hr61qu5DSYWK7OqCbqwLuj3bG56+M
ziRdv0TaxYwddqWdhoBrNV/+xsVw3WfsGPZEk3vcQRzhL/XOPcB9cs9ZNbheMy+YRsq0pi2ArF98
JHW2fsZqmloZ+rmhFIkp9imZMYNZZbh7/GRjHTwQb+Tt9UV/BIy36tOI77tIZCsWcXnhQGqzOaqR
g4cUJq+R2Abf4AhG1uC1nb4e4jpos4Zt2XNtrqB9lk0y5sdB9nwxUuyeM7QPiiw7MLY38kcX1Nwu
Hr0edeCscNr9HFC1IK3LLj/BPr8LH3TM4RrPstjzsBxnVzibiMzQt891i8rdIjB/9aMBBIHNYu9P
9sFOX0NbIssOPpsZwkiy4mPhAPd8CPEyWyIjefqM5W3vPKqOQP+MbcATMDWQ4zTpFdmj6/UgG4k3
vOW+N2vZ2dKA5LWo+FR+x7yLnnfvfU35wHlq/8Uk3NzxaqDOu/3wNyMU/3F0ktGhi3MU/qXSqw2G
eSyEiRpIm1W9dw0Ol6pApplSwZjokpu+4FCJwyleP8gsM/LytkmgMRl+aaqXUS3Bmxd9z5APUazX
ogLVumHBLn2Wc7u6i0vEUcbrzWm4uS8Z1Td+WaxT9WmXz5iHtT+OjLEfgCRFUVWjIwoNl6nwWULT
egQVzWr49f95EjaqYu4u8unWzvLjlEIiMQx9dJjfhFBKfLZzN299MucaFGZX9QoUjzE+7J4Dpt5+
XGJMApRHHnorzpPzcWltu8jpOoBkz+6BI9hMI/rIkdXF2vsFwZ8aVhn5kOsXnDTcDXAPn0KHioft
WrgAKaudAm+D/TtnFqyQhC959tb2sxVTdcbbyrZ+SaElRXOBrrKL6uVJEPm4R6jBhDZgojJ8o3Vw
dD3RCSyyE6mrVoCDrNjRDgPDALgcWWfKQxDkerbXnyTsEZFQ1fcw59g1P0BAus9wAHEB0Aps/oQ9
tsL3OMot7Jh9MC+EqSIaCMoa+iazlnHH1etNiohqXHuqFYvJEWdE2yAPUkaKAITbczwAxTa+TlW9
SDoPIPkOIymETvae7tLEm4hJNyixuvTRI9bkaTLV1j4n9LL2wDHfqCvIjIYW7LsmOUgjuQziHBlp
RJsNvRGjArVLJ77TTgLvHP+fX+q4hnDCJRq3+4RLdgd4GPjE69KsZ1SquO4HPa5Cg2bhOaxcQ04R
0ORzeJO5v7EaVLMwf3NM1j/N8DS9dTja/3tYvXQ7wlmJ8lSvOEFx5WVg3bxTpU+SeQ8NJLvnuTRW
pdkKgp4isYRD++zDnvKSnrzrszbBxKBleYZqHhSpoaYmyK0JfMEwZdQPo21g5w9aP7iy3UmVd41J
3plkiy3iLypPX+bUEIMV4uJzckkpvgX8fxZc7GhwL3acpIZN8ZROoTPiQRdihwSdrj26WpUrm23H
pO3w17zea1VGYezrzUK72XPvaahnaCNMRrhwTNaE+TINmKUxMlXJCFBtxGqtGKVzjLB2sHJzqgMH
z2HwvlrYc+Rv8YMVXk6gMjZnFi7ovOTuEgiVTzYfdX7FGcTg02VMLR3pHabBDaXm82c2+zEtGBfN
9F3tDQoMZXhmgSEhP1KUeUTcU+l4YMt1P7CiDHvoXVekjiASxHZT6e/MZLpwyg2GMYx/1/WSl3Pe
lhzaXJXX0q5dG2ORLFSDIobWdiLA366p90XuPjcKAs4I6HgJx5i8QtIH/q8djjfm+iDlqE5evXKu
97i3yFPAPuys4CP3u583ET7vjrKw828+VoE89QjMcSpG2sbCWg0wzr8I5I6w3vGW9wk/62cORe0N
xVIhxaaa/1j1C+EWAet15pdbcah+UCpeXk6tm8pNdtghQv8zkwFU9f4ERPP3PEUXhgNlIMQ/8EKB
Gmks0rYpEBl9rmrdBa59zBZopSrcZTNsIC/b+vw0QsAosD71o1CpxnHEjnglKDxCzUqKsbZtz3cB
s/KfLRRAU88V/hmnsYeispeClThbciQWce/K+PPG7sN2G+WKdD3NdN+2wxNSeCBDn6aNMXBhpD2k
SnJnt+Ff7OMS9orS2mTUIW8hOXu8q9u2HGn9+kQxSIhw7GbxGRxZC+B+mIuB+Kzh7CCgZKRtMrDA
/dxoudo43v+OeTKraxz8Ev8t7E1Ybs6JtVyKMh4Ios6SMvscLBJtvBsFKIRv1KN8Gzn9Be06+7dD
Kg8s99W690OAUW6jmVaQgmglErtdX8SA/F+RP+t/+mY8+htgV1p9gyhF+r1TfAyC/q8wRtY/odm8
Ldw8vQ84VqgJbCBsFMxY4pjeQDa+hBd5n0eRKQTtrzhJyuwEJwmqZY8p3Rw+Tne9dis3oj+48S+1
8+yKmJmPBTQYHv1aFYtI+mx/aqUGZPkYo28Pox+atMN8NSj15rVSxbNFjpxx89OgNA6WH/XfMqO3
FPX3Ay6WdbGy2ZgKyWmGZOvZsO930qKOJzVTmLB68smzdq7vimv+Hfhg4FuK6CYT0vTXsoNJRUN3
Xe3J31VgYSlnBAGCbYM2XZVKVqsCXhQIRcMvL9laIW2aq4Wwnw1xEa67f2Eubw/6W7wqfru/aKtG
ZQoxk+vvVWmIzzfBaX86NxcUBKiSB7R8+gT+HLgWqLi6hOcGaGg6FseLikD+V9D43NkWqAahxkjl
5hLAG09Mgd0xzbHiy+RtSifgH+NrxOpX1MKLVsadph/MP0WljDjO3xgJcq98AH7kghR10J1LtcAY
VvXwj8ds/HY+DKu1TUJcpZzMFgieroXF+C+0jw8as1CYVdWi0bJNBhSEH6zZFVVPGHWxpTuTj1rJ
itddMbM+Ato+kd1fArWK4NoE4uXjkUVM1ASGQJthPdsZ5ZqhT6ebb1+STaee08gInigsjhNZ71Q1
xeA3Oq3IjUOfrCUTWokCnGn0sQULSoEpmvIF1s3iuiGpoV18Dghi5p3lminX9ViZZW7+6fm+cVZC
SDv8W8LQq439YuTGgNex/pKeWynBOE0Ksn4kOsQSV3JC2FxhwUVzjtM4xATyJnIRRiFg/R5wSgT5
8vew7jFqlYZpjr/lZmvknKMoQzD4efRcprecOXHXpXDSr73xaj89Gth1curwlotPeTm2DZU9PbaT
LaDH9dt5dYb4rse6JifF4FtbD+hkwyqPuFGFYD5BGpLspTNRDVPxQCEXGY/LKouKge2BLCp8sVeF
H6+LUaIm+zbgq4AT+rUxyLpPBFf31DA50lshf5VvIDVahol6P1R5B1iz7FM4JjaEvvZoFMsLAC/j
+Wg9N88KTBYy7I/chgSUZj3GIMI8vgzIvwgb75/8L3xRsX3MO6jO0kUKmGEjJ4AY123T/9WqXQ7A
nknugqxeVgHuWBsDBTshZUdAl7yPXLlCzvL/8+dlN8LVNh0Tm/uBsPyu+l60uA+qfxsbiDWHKG/A
Yhu+i4gnkLF2A7RrGiQg/ymmaYCOe1XBS2VKeQIOUls4m+e+7cHQyDOacqJzjsv5nIiS6kTprIgB
ww8u/NM/Jxs90cLFUUmfwX7lhZrv0+bTXd+6L3G57lSasE9bbmYuMSeLWXOSTSMtsHb9ph9eFJn0
fXrTN7Z50ku23pOWwrWZ/dHCGyg6CTJEe/pXTxhn5GC5czxUQSKbYfE5PoyQ7HfAHgWh8np1BPoO
Sm2ZBE/KW0Iw/jdSODs4ZKgYHw5tkPmY3kwMVUhLt9/wCIrrJSAdkeN4grDsQ12cCDaYKobiamjL
ndV/nkhBwkwoct7nPYJ/VJPhGpBGnjKA9DhRuRXLufTvSrLon45VUENKThJGY/TVh7WorsRxgsYC
iHJNb7jQZvK5kWNknGpYJ/YAxglSQ+vet/HHf4pnxXQLvi3mFyrJO0zH1iv/3jfFDaaaKkUTFeRX
a001zAs/M3pTIQZPFlARkyElFXoB6AkK2vcGqLBAVvxLlvqnv4tkrRha/Z//ngLI+8o/abIUk5a1
SIcPv5mIICc3sNUr1X/qlaNbMI5GhKOi4Xfo5ZNzGeXAviqG34M+HR7SDcuK4esAE6N+SOY0frHf
EgQ/m09z7rREnzlTjSaBSe2O6crlbRFDn9xCca6EoL1K3DxEVxeQfoFMb1dJkCB9VBsQN1PPtx30
c0CZO7aRnRkIpnIR/1wYJgv4scXKv/QQDE2Bd3sW+9Z2GzIsWgSE/U6/VXm96B540mhmnR6KrOl7
ZZNRGbA8VfZ9amB5lWN9YIhzhKGgkAbtf1jLGjfe26+/Dc2pkPFFCUs+CrGupBXDmddayzOhCiby
o0ACr0y6U7Q/HARQLAxxyWcwzRjHxcUwVPhlohKNj8L6X5C8thtISinzBypj4pJ37IBReA5kzEqH
7E9RsfEnnBqqknLP2y2c6Sb3FAHyf3ENexPMjNpBXkT0SYxYNS4m4H8pBRlPScb6ByfzHhO37Bg0
JAmY1LkfUDm82nEtFizOZQ8okddGb4Qvk4L04Hh+fjNem4PJtwQvhwHyk1OpYPZa/SrhbRza9DgN
sF9L6/qBkACubUs07uUvDnsBvFDC/4C7Wgb0yrHWDm6Q7MaxXPEVc8XwfQpyEyNLneHTqR/hmrOg
V86RcYVXVUqz2Hf+0zoedmZGVtJO88pSc8Jl0UueXCB1kEfFaFhO6dGegTYAvAJni1Ud1JuNQHS/
t8H7ZhPXSY6Wi2wG7G9qJZbsVXA89tnTlInjxfxlRUChP8nRFCfBOTCHKPuDCVvsMxTE/hx1Fb0Z
0DlUAU/0xaxvz6Bu8bymDJeuoGyecDPYiqYqy2/CF55DJFv899e0tR6BnMcm/xxOzOonSFL1QvAi
V9lskCJq6JqJvIZN6DJsEQInOCT2eWwjfwY23ojwm42Eg0h5RCrCNBQpJphvR6z2P1TVC8h3inuF
y8FxrbV2hRntSBxnPdLHzkonI7E50xHtMOqk28Ck3Mv+SbAL/SmoRmaJvbZ8bey/RUYCHqGQT14l
NeQTr/g8b+Tk0WUPiEMTWSezqUfB+CNYwmtNpTiFFFM6bJx5wvCpXJxXWFlJxEfpaRjHdzjhgRV3
UhNdxS9ZWw9GXpa5aBgxqTbK9xGczsQQNhl0lgAFcKq/e9XlAaAG9Pw2NIzUAunw6s+U3vK9ixge
75iGD6JaaaQHADSlHFLUBH0qNq2t4WPjgLJPT0hBBpNrnk7IDprcK/EKKvK1LmbVUNkC1ut3HuEd
3Wobr1nkUwC3qmsUq213gtFXOLVV2DwfcbnrMEEzLut0O+uJ8bVXih+FNewN3KrR9GCHYufDTlnP
ehr8jnAXINtAtY2k08dZXWAoyQW58dXfFUZcG9lHf3AL6hd/yO+5I8EbBa1BNzd3Tf6XR7MhTWMe
gvkUjWRIQ06T6AjdrXdrzlIO0yTAjIA2I4mvlzrvY4wfSepPCvp4T2vPVhTW2rJYi/3Cz93O90Lz
s2V5oy7qMbnvG5zCoWHVI/M7XO9eTjtZE7TwZz2lN3j6D28P2jNQ4GJpPSRoYmx88S4H8JqKH1Ts
One3qCDFhr/5ngZ8nyuRc6zqCpQR/rIxMHuYelZmt1J3AZoAdFM9CrCDqvyiu7mejj7EwRpkqawg
oCeROP9FgoAcFGQzZIKAds1K29buBU3ARQDBL+KWeauoukgl4KVCy9KBZ/ZzrWTTd6AnCD0IDjEM
QjgXefj6n4vn9gE9+YR6RHaiXPYamQ1HlGK9JqtcpNfxL2DzlzLuyT7Nf24SfHOs1t2aqzWARg6t
n0bmAF8aj7LiSmL5QtArVt2TZkz4J5DoTdCSlDlJBJQbFPL3VHSwgsX3pgzpY4nhrhbKdKFxgZH2
N0T0EJAymdWFlGrnYoMGVw5DpACiBaU/+riUSLJB7lmLZNuunq5LiTVgPxZIu2g5tJd+1ybYy0AX
JZDiGM2tpxLg/efDJ1Ie0JWsrc5thkdvXYlnwHpErY85WVw80yh6kptQ5L2eqSUo6INPzehCrFMj
qVi5uTgrKDWjSGYvDEJzSoaOeWR0Vnh86mmZdaRwoyjmx3/xPMqiRtMmNDy6PiGYFpJa7hh501ig
/t2SCWflT1/eHh+xTQhZkoGYW6q4Akn2AzuOSdqFs46ABz0nEG+HN+I0eRWhni4DppVjp4LSW84w
cZio8kW5flYWFeTez8b5JxHNFhSTiNPt/LwhuDuR42tm1kiXUgx29xCnR/syGI0f0TqJIhRoH04u
uoPoAUNG0KHLZp+sOCDues/zcfs+mf/zvg6dK0AbrsSTX4kI9WR+Q1/Sd9gLHl6yY3NORm4I2HVL
wM97Ihqz9ZgC/VMiQO8+5aRcE7qom/rKbQmI4zIkdRxlb8Gyy/0/p4Veth5UnzHVQxFmf7DCqtuS
Cg1ZUE8pepS+AmlS4b2rkFNrCVquvLxNU9Z8DgPVfnMX8/Re6NkmfDVWcsHXrA7EAy9j5GM5xxrR
Jpxb/1PUlOgWEQ3aCe+bWM/SHkfv7DXtk4HZt7E9qOfk5h3a9QeeYn/s8oX5Cfmn3pviJ5ThXPPG
kF4R6xWshQv4iF9XpuBnhuU1Eb/eYwFFn8mbA6OiIhFj22qkpzyRDJFDayiW6Y+YHesI//RlEZDw
zbFhAv8gb3XqcPSwW/3+yPpOyAjy77AusquTwkVPoXorhUiZWdB5279y7j+GEDAAwj1R84NSkLA2
YExBnFNvD8kx2bP/jvNVV/aWdz4BCOwTQnL6xfy0PN4NkRTzevi6MlX47cJUJbQFf9GfDcO1c+FT
4FY+DB+dzifm+6RnyIrApoG/kUirHPt7J+YwU4NHnwPtqdoFQiPQISWAxE/zgmy6r04G7GWLIxDN
qjk6qp7VMUR/Gik/nzIC3FVDuDLIRnESt0sDGbKKx10+pgbpGkppbQpUECGFA0IpyoJAAzXd/vnX
sqkDG5ZRhXQDHIzL8bhPAWMD7ocllTMui1uq1h5daQlUC4tvsLZr32nShf9I+JcpZhaeLzUa92d4
iZ4YcmmfgYpEnTegE/jd1f7yKZE4lG+4uzdS6pQScIHul6aJs5JOB1XnFVU6HCFH3mF2aZTMaIcP
It62HOn+Hf66FP0NO8xiQwwcYJvJGk0ChX9/00TI6lwGzTKbyyze8Q2WfLXzTz77kVXFOlwK/eSr
tDNlWtlPAPeiBT07LOZIdpm6zMTFflG/jGTClkXI7C0E+4HeNckeHLc7ebQNUJUlAzu61BzTt+/l
zt8iiQB06H+K5jS2B4Tfw19cPVjrXu52XwBZCuul1mYNLtV5scC5vK557mUlGNZ9qYH4389P3qZh
4qjWAahWD7kGxTJDpLGN8GU5Zg6dzuSL/g5v5Qnj/NZZhNoumUAOa3Asld7wzO2tv7UJPdT9ZrHS
RcG7suCag3kivJygWuxSUHLN9wgxMjV56r9h+SetE8h9Yu7Z9N1nClrFTExAL1hAPkwjXSHvTMhm
HPN4EEh7F2Qy55ciEXV8IZLjsdmbItjxBauNU0/JQdSJieFAWWF8N0Bdia7QkGclcgwLzt0kR+dm
lFPmLEANUT7JaK3ZK3kw8my4RdEP0BApXDy3mp0s3IfjYxJWjuRQjmvqj45W3P3ii3B5wHHBPr+p
Ywyg64V5s45V8Oii7B5CskIPeR+Yn82NuVGRib3ix77w/X15r3bXg5zbULzgL+Y0os7z8bKo308+
mK0f/ckiDgbpGl302ujYn2uqJOm7bYsQt1/AXNroPrLpsxgbrmeLNdQHU+d55etiMh0tJVryf1wt
/kCkf/UbU86wbzak2Em50mk9z4an4nzKdba2wy64z+l5bCBKXmslaUgp6324vJ3uZYWtSwwHMI96
uBPZjF5OPGCVmpv99R1mglke++9uZL4zCg24EgOV0sn6j8gY1Yv8LGEIFzXA5jiLUo0IHYAB1YLG
xp8hRyWuvlhFmvuvtdN4IsxbU7xJK74Do1IEJDqgCbc0XHpoPifyFq8faD025ChCr3CByqYIAyfc
FZ38Xx74C04I9Jj3EkNX1lXwoI1huO7AKsdtE7SAkaiSU2uLu/DqY9TGl2Pk/v87AclmndOIa6mN
HOXWqoDFTf7R6mCWFPahQWr+7Uaz6PvmM6nazmsY7RNk+gdUlfjbg+x/NlMJso4NOlQwb+uOSg8w
/Ms5iqzRD9AeJLMzbWc4CrgJBa68JUaUyfvmUjCaJdjG/QCZge8C3eYVMymqHjHqRgyNp5JqN5gu
7C9rj0ASHPoiG6TmnZasYXIPbHkqfgioOMTOHKsnSGkhhp6qfrey9Fh4JLV/J2XYaxuLPi/vlvRa
J2W2GWNfQC2JNLlR1QXguoLPEDo8X3A7YBf54Yqy9KC1Mk1903/8zINDTJ3krCGFKubPXhC3UMFQ
1G++2kI8G96z5bOWMJT42GpOMIIZCaMRA+HphELKpLNt1UC2qS3WOofIKruI4zPdJErwf5WZn/4b
FpyncRGGiM976u/GqxjwLnXeFzQPHOXo6mneC4iFPJ0Z1iXp3ZUHq4XSSgbov28CqaRcKeZcRyJA
Ab6k0wEsVnliju4I3IN1RyaZqkAkzkHWb6dRQs3DrWK/qLVx6e8Y1JLtp9OJZiIRM/ROaZSDu0Jx
yIxNJTa6baLHeqD7zxpx18qivg3nVb1lSxe8CzrMmV+tEsAk5SoCo7+HiicXdeu+h9Epj88ZNFl6
2LSYqRKmH/r1SXxzIqyGydPx6gsIkkZkxgWfwboq4JMUZHhnDwgyNOQrhCu2iHES3Qj23LkhPCMi
cJdyfBsc2AqaxiQxAKMGW/b4FeLWeLRChewB7gEBbqW7/qEetuwZ9QvhtkMLXfqRy4hwrR2+6Ui6
s9C4OY1HjS5TIucJT8jr9wPxFY5gPTzc7nIbcvyb0lGJ5Q9EnZ9tD4SozQXozkNdazrKlrPeDUlh
FfuToXS1n97XBbheoInfV1EtphfXIb6ajAHMQX3Mj7JfwgZSs2pUmCMEKX9UK65iOPQtKfvdu7/S
ndVb++Il1kaK9PCv2DouhGqHAvwnw2+G4yi8VVJPgzwXerDShFl1aismQfWrrt6mGYFhaHo0YuIo
bOYcuY4T8GPVb+bfuRYmYzLDAoCjJfu5BB1voJdNOw2hwZ6LQ8VTISZReNHbe2R64BDhInK34wDa
XnW3O6aSUATHA1EOoea3NaCw5jJT9RKghXpj3se8AACFK33DRDEPmyW8nK1BeKTRylblwRrACmV2
Y6o1L26DUgnVChG5QgE6EdI6J1uW3jWqSJhR29VwhTOoW+Jl7Y15PdJw4OO+nxOVINBEgOtrk0wH
+5WZVTnuXfgS+LvySwsbjmrot0q+ul2qvaokcdnSSNTzqogAG7UCCkTKXk1uT4osl46/rJaMNeU4
hmIOqnfb2JF7ZnoMM0i2xaKJ1Ffwhr6TYVgCHvWmPpOO6KI32/3uHyggx/nFSze7dw4Mr1D5SGep
Nzy1dSTVQ2IhI2LJ1L7GGgdP1KOTUxievnqBbVG6+8UiCwr/VxJzBNw0iAHHDFlY3/JXRNYNKKsz
QfqsTnhtEs9aEF1sVlA1msPZ420ahnVQ0Xd5CKPXChKLKVoGtFyhk/lcUtG/DEYzACHSV+F3FsKa
B4m7/TxWZPgzAGtfJfzlE8K1XfLUigofsaSqFXBr5EVkR9OHXdO5kaVF9TBM0jsRSEJPuSjyk49D
kfs02lUNVld7BhXa95Y9Sk5oSaLtOxZXzvKylhpDYhUxmUki+r6YjJzzH8IgikLfxRmwkwxI0R6p
Yas+HMjjQ3y6IUAswwbOXbX2QU57zATPQwGJ9SXxZwq6WH6bF3QSEaDh+mmBn6Ct0wmQuZebGalP
5XfneBllvgyUYlP5VxhkSBXjf8NZiRisaZ1ElcBWxtCEydQIAV1+xaJhi+Up3+0dKxk6ujX7XY5l
meddTxNrbtqoV2vv1l0P/iJV+xEkaNI99WTCxfKRPH0zr8C8+0garr41wqrta1Q+nWLbOB8IVrNt
Ak810bFe3RaS0N66GTERg8f0ZFwmIad/AbiZDwTTk8VQqYRGhwDRYcOkQL2+iyWiu6poAXJj8fPk
ne2pbSij0hVZ2Z++dSRSZTh5eYXyCBKgK1kgt2xGoNLwVHsAaaTHBNLXfXK7O81YumGkHCkBJowY
zpnglVUQrj5BW77nkRveOKDKJK0x78hnXaverttwCVO7TwS4sDlxfWOBdKICKHlJQXIf88S4NM+I
ZhdR0Qva8hXJYTFj+J8JRysPp5Ly9HlLGBDQ4VM1Q02tkYjFXPivs2aCm9EhxZsHvdbvPOw+pC06
K6DkZxOIxlgeLh9d0WxPG1py5xWi5GgLkGP9L4p5HmXmFDzqhNbuKuZAxMdWKImzGtOLdONabk/F
Z/Le0A7JgXVhwV+Pg81fDMGBxaXLbrviWVmCjLvKm9d6CnCAMK68BCw7OtMDMed8wBcBrAkLT+Bd
nJk4q4lGuMchXLCbTDBPngLAJkwKK491vBnz3duSZu6m292j44yky0qPHcxTsRox0Q/1FPwiO7Mf
fqIXjKP6sATPDtFbh9dkfz9zURikqtKvnHjzswwyisU0H1+kcrxX+FD412RkmCZFu2oj/RFVS0GI
zvvH1i+vUnxiYTZ5vR7N8oX0VIjCalvTsyxIFKD5HTl9u+KItLcbDRXVFYXo4WhZYxUSNAMGMRxO
v3mNql0qB7u16G+ZKG9kEnjFX3wlMHVWnvCFxJoTY9YdUHJA/5XEY6WtvN0oQCJ6vlgakwhPRMAx
rckKGciuXuZES40XjShVYctEYvyiW0RG8BIFEtMvIHI7OCsbjFzE3Ij7v5Z7kJERYdt00gcaEipX
cxqQUgrkRuRti8RFovwkV2G2o8beAOiZDOVgfj3c7r5wcBlANlFgpCPTZqcdWTGZGzQgc6Hlmx1V
/F7rJ13ZScIbnWAFvucGe0ChUQtEBW3Uxb6I0+LpYbh2fuSnyMNsmCfCMh0o6AB8W50okj2esRAC
2OmOEMciMP4AH7r/JCVmaVzNhhwG9QlgchBj6PhfKMr+IetA65+RZwYtgVbT4+LXaqZq+cHC4RZa
OlXNWf6o/wVEo3gOzo/QOlCIGCFjB23UJ1p6KF48qXdPTgNKXpd/auTpZaQZ63CNv+wqL/EW6b+X
L8e6VKSbxK8L7Tlozx8N3EQkXKhsyT3vcqY/+TlRQ/1xJnfjk57mYFiAOaYE73pd8UBY/wjH3Zaq
NdwJ8ZN6uRi3gLeuZ7ZIVBATSKsVPA6PmmvTtKfPR6KBURD6GZUa7oQyZv6x5QGiswaDEo9h5AUs
eJgJzICVjm4k1oNlHL7Bm+d9RCTxuV2vN+/tk4mYxPqjHVE6iSu1h2TBpdwb28QNZa2g1cTQ/hrl
/I5ueZkeVpxb9j1wpGPcJTdv6huOiXQcJAIxo4fEvN/7U3+zms1pOL32bobV0h8WJkZyxKSoNIhr
qmtJ9cjTn75s9dFX3agLPPu0LhtncDTCR6zbXWVvpSJQGWFcmoaqs/FPb8wpH997B7jcux3b+6KA
wts+2Aahk/uh+URtVHnY637+yzvWrIe/sfeQi6K6rVfSfeO3c0NhrpyEjV+M5oJykUii3+pjgbNn
f6WofRl1YWQ0KGUVIX/j+1XnnpmvRpAl5LlqcKOPOSNZw0jRp9Wz5hH0LRZ2Tc5+2zFPYRSwjgit
3JOfze24k6eheaB0U7OXcdcHQcsgFcldZB9ufoJhUjm5D1YHUV8TzuVBZGjJr2NwMhTcuA4M7+k0
v8M/l3V40gQHreJip2zE/crZKii8pGQZFZ9KLJA3DeWJh/5yrA8qQYGdiTgvConRfJmyq3FiMCK3
Um/FV2AWs03GzNA23fokg4RKbkV3ALk239NjDnoFVR5PnJSlYfAVe93UiLkQjCdYB8utpwsRuUhe
ORcMIYa4x/kl0TETzyXt6aNAo0AaeTqCQa4t0SyCk/cSbEnZnzNGJQHkPapybbdwEoHCf3khKdxU
Ff/qCNFiapuOCuGPWDuAi0Nz6F6UeAx/C5SIKokgmLn+OY5LYybAVPgKb/p10/UiQJZ1QDPqreVj
2pzLvVmdRvrc6UdnQOUC/WJHGu7BuNTK7rzvHu+hmEGRTkzBdN+q4ZjRX8LT+VSS6GJ9wuPdJuQO
JgJnqkJbenChr+dyjiU2ldY8Ww73fuBd+E/9tnOtjt/3n1SpnhnIcCbVUjM8XZxw8sjhuqEDHqvc
dEH3w19BgWKjSqJwZPTFuTDQKt4Th4Z0OJ4OwVfnSJcdkXmoeiNdwqQnRpESsKvkWJM2enGbm95r
Xakk/btjgEfS61UhqH7lW0cm0RO+8G0driEEUY7LJHGArPC9Bk8eHBiz4r/p0G6ZF9VgqTu0WRru
cVwn3ImgsJnphZg7XQKsR9+Jzql5XYUBVj0RbLz5tDa1XqwxcMPcBXVCZ9sMmlQ1UpAxFTcY6+mc
BHiYQ0P9MERo82usz+8ik5SuDsqDvAbiq6fxQFz6Hfhrzk0GLw7W7NZFBuz4p+BSX9rObnvGy8Sx
OUtM7ZxX8lLNGqmo2jrAuAPpAXb8Jfib2LQJuxt0kjgnL1V4rle/uF7lqz0fbPW25FNt+pUTlbvA
BvEU3atKlEiqPH1ZgNaBCN/V3vd7AOB+ImGUm2KiqRYgd5NyoHbgLflzz5kskMlFrcDd5YmBxeyb
VgkMnpCgouq6Wo+pek9gr7nq1M0qz8Mpl0037kLxFKBMgfjK2NxcFbQBS2/gLgLc292XkT3L/wy2
81j1Of6A75q5PPtkuKvfbNUnlpUAdKB3egP9pPOprAVry8kgsNkux+K/VKbDh1Tf3XOMt8obg2sH
3m+cM5ZEm9LDlv60mOFjJ4jUoNC2OCCywabqr97BLRiGm4dEF8+UProkR+Yf/ersqv+ugxrBmiSr
GzmMecinEAimCLnuOhoj+fMi/CObHIcsiMDOtY2eKTG6d27q77uLiueTT8vpGbRo1VogWMVugbm2
XBdjYU8UtS1r31D0G1URuqJk6Lmo9t9PhsaHfiBedAT1cv0Pw3wsK9OCOZReff2QRaQDVbAuym5o
iW2Qn0WxF4q7rRcNUw2bw++Pc8XcxcYs/EQSKdGxZfGHQc8G/vj3VA0iCHoIGQGFjcfN5wZQl8MD
c3yny1Euk6UBauaaNbobAIK1GCKT+R3bE5A+alqPVeaUSxhZJHjZJNdI5snVTSV3P/i+6xCVMQO7
SEzCZHACbOUbBdr3afaV/bxvPnxVvXV80vYJMVbF3fpO+L8SEeZ3v028+4BraaKxQHfYoTPaKxh9
n8vaVxbvwOMQqfsUr/mqHH2a1P+eFFmbTIhk8nRa2gFpU4UwHvE8kP7tjhEkG0XLOKgKdTEPpWrA
M5UX7pT+D8NbMijhf15dquC7cLq04iLapbT5Q+qeykHkTXbDqzlwnAPWdWRqIbONvUxTb7eNzi2f
7O4uNcMKYkSSfh62CkIbcdYZ41+6g2gv2dZZwmM120Yj+orFONbY0AWkRNzMWBdmlPA8JtHDSmp5
NAZitqowWsvt6IrxMl4s+AfV9qzzQFAWwUBI6McEhj+5T4Cxp4DEaDX5h4rpGP/tUx6hab2TMc/G
Su4jsRbAnpa2eqaiznDXIVAbAJp0GaVeSydwORN4ZlJE1naCCrnwhKAivQHfVtWn6/Xo5keB4j2n
HAjTU38ZTxP6WItOTKzF9farFgGyXUbA0qUUoBaZkb5HqbUD99y7G9YVxRQyHYITLyhL6ZAnN7K1
SxuGzNk41CDoj4ArzFbNbem0ZPRl9b+CqUgAbQ4++xu3KmpcJjOTUpIxhocuF1qzsNEkW4GruvS+
bvLOdsPejz2aQyvhwMryJDjWquG/537w7XXDdkhB9zmVwqp2aYsjEO5v3PnmUZsudHf2cZI29Ttp
TWv622m10jNQmjIR31CGJFRizz75TvdiJ6bwC3/I0jm/J0icvE2IatG3BrP7Ti8QCcKVEOyMC3Ar
OOKp4ghgxZfPNVSa4Xbt5aJ1I5M1OtAqOob64nQmvptddoW5fytCLjDkBahikIQx1ykIrr/ArE49
IG2VEjCU8AIZaxc3QzFqPTr8HVwblztqz5k33n+TRYUB3d3b29r9Y/y9xT7BhszEXLB/7SXly4tQ
5m2bGdZ6Yjzb1YkatEJPFLADo2qIoxJ1IEzIP5+bNNy4vwcpsFIL+a+GbsHdKNCrGOFCqu8yBbif
rpoD7EYEuw3OQb2auoT/naN+gVgnfSJ5MN8YQPz5UQ8Pw3f8137t6r5BdU41O0EkHneMoEX6Dlld
j+dw8md5CEHUgtIUrYp5+q1dh4GT2HTI47hPre0XY6/Z2iuaOYvaJMHzvXD5q1XBB5PcErU7k3CI
MzOhN1CXE2nkxW1gVrbYUEaOtuQtxbnNOaEwZn5SBnK1lCXklU+tFl9qmislJRDc7eKmvtgczv7r
DDVVPSUFGqhV2X/toVNoJLFNQZNcGzguDKXoUUhGJdRDDqVXwSKBQ/HkdNSrllgv9Yj5tPVYZRQW
6BOSUmTVx+ge+Zi9P/s5kG45uDue8jQSk0s/m0zwQIGnS7dfJX1lYIF5aMcG4Bt0nqV+T2CpV2O3
9MGDJIl3gswVgjDqEZtkWc6JZty3TtKNznXCRdWUo3DVIG/UDmnN51vIn7LoLmNh5sLwELGGMSL6
gmHVhwPho36MGSJ40sbnDHM1/PKnrvcXRgu4WJw4bWp4B2FUvDygQE+WJoTxDO5SFqPXr531zQsp
uCtC8S5na+aF+145hcQBgTHqDR4nq2en/sSov6OBmDrIpnmeXfd/XgMBfRzn2ucBXfSuUMY5kUv4
ck6+vzFm6VZ6pNUPUhDtTYN2uAXt0NAt2CEybC+I8qRf9GQifojLcizgNonx4aSemJtNntJf1ufg
1CKY3qt1o0itf3XkONCIpEcRtY9BoJcCSNy/43RLz0MXX7rfCI6kPd608d+319XKVNNJ9o7nDbwP
g8B3bsQqK+LzdsGSqBUJNQRfKtQisOjx1a0BZTOrrOBEu6VSCtH41CA5VofrVxIThW+1bHLyHrdO
fm0AkHEYUb94vpLjHCUdUKEmq1cOX4a+PYreOBJ7LRzxAGhEcRQ6QHFAFuKpd+U9g2xjhSjk0VyG
MAurp08pgPoKf4F0Yja9mmHPzkPPLpRgKWIGFzM/BqzYMjMiTmsCaCjXlrNIjjk41KQCGJ/NCG/O
1QJWA4007S+t2i1SanG+Bqg+B91nSm2b9k+NpRv617sEecKdoUiXiInpI0AJxWi8h7RGY5AH+yMg
Z/RzUdJWWN0x9EF5y+kGs3vFVVAxHfO+Elwmlz5uSPJOGe2VRq43fhtk+NFan/6myVhjM/IHUU/F
jgMUVhp3CMZmy/074C3rSzoZ3p3lUAO680AXNFwQVljEJVF5qNJgacmUi0pv3mUVS2c5z965+SK5
5flPmL+7jAKZC0nYlI8YWz/dI5dKhBPs8lSsZgPOrn2dkCMftEtWV0sAyNR54i0Qd8AV+6Ic21BC
JLqLYZRM2hd64FJw04FCb0uds5NCyFiexnvP5QiFhDDYpZuyEL8h2R4b3ng+S5SfcOKo8Odc9Rmy
GqAbPOw1x0p4vyKENhFTy8niy43qqjtyaM00O7l7K1/6gTSU+yYSx7FHYH7gF0KvWPUViW79xos5
1qSf4A4/dF73twMkkyaj20CFzWoHWBgJQasSeQ8wuEufpALCxQgOC+MACqOUm7XrJVKmeHsf8hK6
hN0pFTPPe5zpRPuRmvc+BpTVob57PGa08Eh4qaKKbkHur+LCTUapQUmzU/ZlPiOtXZhFcgDDUPT6
5kN3kzv5kIwJUlrrMaN3UONfnzZzXyNwTCDJ8MONAaWNgMQ0eaKb+e6gEGCZd/zlk3tJyLVqJL5+
GUAMzNHPpX2QESnzgi2GfO1E09JoiDKtiPMMmaGFpjCJQGhbIoulhrI7E0v4AlueVUulhKd3VIsu
3SevZMhEruXk1j5YABsDM/c7lTrIRNYnpqzIpTP1gy0AOR4Dd0bZ5zadjvDC9FM+Hn1H5NhuvTxm
UKCJX12gJyXb1V6ibmMcTOM+AKRdie1kuCZ5Ih4EDGIDlpY+0rsnCmU1oL5C6M/mSdOXIRv7Iuh0
HQRbhZCxtGzbrWl1MQwg7kZnhVgS+T5DBSYwa19TnQCFrAqY7Z2O3CA/0efrvkS4+btMXCdpQLLJ
hjXqsSuChUg1PA8PhxHN+s8L1TbOhrhhZgLPhEcxrW72jf/e0EmE1yokzDkuJPCH8VyzYyh+1SUZ
8TivjL6sOaXIYbiaV4uVfPITUVKgq1Jm5me7bncvQSSQtP44yZsLjmJlXRYC704u3dEsquNZzxWN
gJLPigsqaRv0rTiJ7pRZUxdRYh/qAgmE1M9K3FKmu+X5V8FnnWsiVgvQF4c7e7oShZdjRsbB5i3x
AIa7IcaK+6HQ3ZUYs2gO5ycdX7Kt1vT6W+vZp6g/P0NTSw+4aUOMoRgK0vgGGwoLtH7NYpf33Sjr
AF32YlX8OuvNAJj0sQeVDAURl+nilm8RCGHLsCk3YixfvP00DqL/V9Dl2XmFu8+vmOPEj/o+BWCF
ZHqyGzQ17oVw/SQtZ4vnQ4RM7isGFn+w/LnCCczr1ogM7Y+Fa1gAcDkNvPXzA5QvFq9jR7KXlZxH
KUFPbzSbv01+u+IOJxTskhZnKOmblPhO0FeXCqFvty5JsrQ5ShLfoDzwRwLQw+lTUkkXxM0TPoa9
ohaTNcVqVVaLeZtdkZGEapr19v4PbYVpH8Tzin28yDtV+i3ADFMPo2iC7cwbnO6bYWasrRPH9qhp
0T5cDvAxZXZyJysn4OH8CawNVvQoy9ZjC9gILiHv7PdMxfRuqWjgriDX5rNrZgyea0R9iKCPl3oE
afXVTr8uRU0JfQFE7Qjc+W/2EQR9VS2cs6HkafF7yd0ELG1adTo4l+QWFrbyvGalshOrFz7ISOBk
q14x6JHh5CXwukbOqdUjsiS5v1CGx83ADb6RCTv++AAWQbpgp440wTvmBzAag+NGZRYwImLZJA1r
u87oMeRkInftqN5dhEnC9yCLGk978EJTcigIShOxX2ST2CD+DLnN8T9H/38EWKahT6yZICYPnYVf
Y4+i2ILsVUcvKcWb8H9nGeLAc7XdBMxDQXZA6PEoy+kVgSOP8mbAjeU3a6JXBHpI34b+ALN5HAIp
O855Zj8jcBJ4VdmrfwsiztrIc3W2f8mDKHER9JlTzxzVisPPgpl/qaAm0PpBS+GSNB9aTDCAWaYu
VBTEmFl1D8TB5I1d93GFlrl1r99BULRrnjE9cZt1rshEnptNBxaDwxs+kjdvpzPJE6w2soHhsp9p
lC6p4VpFWKUgNFhdOsBwpCEeso16uvsJNvRD4s1b7AjF0de2B9FYn1QwypXiMjN/EovQH2YJP9UL
Esn7PrsSIcFjUdGohWJ10XmIACX7B/sxALhwqBK9YYTNMHQBCCXZMtPef1exBvh/FAPQHZYzuZHu
OywU5JCtP4yqshHD8ujfafRgWXZCxDNCczCoCAQGFruVo4mByJB3nulLQDMWU7VmSq34Jq80UbxS
tJeq5SAr06p3ff+RWu49wqrnDUpp8xNizcqNWqAHLL7b6aITreASfe3WsHbOR77yJjEvFkzhdJiJ
/Co3LjF6UhsdPowBo9fXiy/BAWA6ex/+Be3R94raRpHMYtpi2pfGGEEz7jJrvndkkTq3uD8UditC
+EsZcqr3hWNqgaNthAIfwBkRMNTG5jdVVxraPphm1aoqeECuH0oHwC8nIVDlAjOvN/0WxEAumi0d
jVFEFFbDZXzKUnsbw70gdwEoRzLjYRxBUFroE2excDupy1ujAh1I7mjjrD+Az4tqEJ7gbeW+Ru6H
X9K0xHTgbuyAwlV3kWSKoMdf0/+5vv+dUGpfjYVvhIdOM4uy+RAa4OXK3T/IHMgvKzawZ4Ol0rzD
isKBM6lNZbBLUGQYqEC5KosR7zoaVinN4FqFTWa7cFezisiYxMDErNPQT6hq8Xm/T2p/2ySqCwP/
MaNStvdvQgbwXLYCiBYsA6xP0S7aI057O9O9lkPuBUblbQ7xHhHqlq6T4dpSIdIuB6ykpAm8y6uT
wrliyN1MMVH0QwGd5CbCQRWSV9Lunds9nyepqJhPB7oSyW8SqqwQ0Dx79HKXREZZsrK4k5PGnnnG
As4L8dE27Gx3mLhNwskgPlXjwNV/xIGQd7Pt9YhfHvaKOAC1H3wY3XD0MH0j3GQpKDiB51gm43Gn
a3JUtBTun31rjfN830Cy/0nPr4O+mA/oB4RcNZogRd6DTnv5oR/HFAa8wgr+8YC7CIrFg9iKRGl9
vT5LTTNa/fRXreVUPKh0dX9S6ZBD/5KsIsPDvusr4Hq4TAc/brgLotRWN01BE9LgfVYA3cO95k8G
onxLLi1eBea04zEDSnvUaZEHilfRSgaaTLX2ceslAGFoufrREmThpJgZudv4ggN8niAllDBc6pve
WvZr09Bm33LI7SFGMacS8EFtm8BlZjMUKXqFeQL+Ry0ma4GxRgksGTAHPv0Iahmf5tA5owNr68nj
3Smo080oAWyps7cJuAvZYn4bojnST5Q+Yd5kZtNZaDE/jWodU6Wlym/75Yy+1fgDkk+nU0ixdba1
eO4A723mjqpgyxcxVN+DY01nplN/wiogkfqZN/rcD7Ku8HI8fA9Dj8JpYXr4EuVql77YU5MRuPTv
p+8p/Hd2bkGa7s3MfoY9SqyjW8OwJSL+KQdzNx3dIKAfGBlPzLBDGS0IvzDilmIXjGm+TWsFIUgh
F/vRQ3NDNqvFWHEgPGluR22ic+1mn9j5K2R9TV8QfHXNkQACZNptfzsr37MbD2/nlv6k2jOwQoIz
9ip8zB7KYUa9rkPlH4akkYsPbGOXEM4SseNZ/7SkSEycXkrsscRQXpJCKbq4deMQT0rBUU75OKCS
Riq/E9QxyyjTMjBOpP1JdlpQT6jqYNJ0A4rcNoSMiilSKYvVlmUQun2bUurdRD7z1ZBP/RLXASEb
r2jXFUOcOirl6FQZDbCfNCN2HN+ydSO/+uHrS5A4V+yw5tZUK0Ui5jcuY/jmyCmlB30GPxNqCoL/
1cmWI+OOy1uY7Kp4cj0KwuEVEwnuARkIC03Ui1RRRyhzbu8OCx5niTTauGuUtAN9b57quB2neSbH
PlC/0VXKpLEtu3c35OyJBSIfrQzsQXX+txWf23uda6Ms91O6ZVzb0yVPtnzyY8wKvbbNPbNWs8CO
iHgPdqcBJs18q/Ua5D5TjVkgBOFqQs4OBhUJU4MJvvazw6s220tt2da/j9VA8hIJR/h0NEiM357i
/gRkyykVbbCyPj99rbJpam2mpMWsQEkRFQjXmoxOfI2xsA81wGfMqCOzuThX1q78ShiEs7Z8ct5d
8HyZQfYlikmWUtHABapyyN3bCeKW5iDBIp4wo+Q2gjciuRqFZB1T8GOtPPAvnFAdZ2J2dPXarOsk
wrAaPRSiGqL+1RtFmQZW2jmPBofwH/sI8OHrQ2jz+tJJLx/RUVKmykqHO9MwCCRYiT6XhjE3EI9t
ld2G9WesvzuQk7JcsMywWOeJE/6bxGoJzZoX7oA5M+8ipewXBOSAxtJw8wsQNXjPKV8gppSbvgrC
JyTZOj87vizzmMY8KZTJMlhxWrAAAVEY5UCnSP3cPmG1hK+94wTo14pzjreGl3gLus7bl4SpgLRo
vLYqVBhJoAIFNw/Cu51/hfYpkCYfizvOA4yYbjcCyr11VEpg+2ZrZchgbbImSRT0rRrE7vIPkvpP
nFkD0iiCYhu3ZCbTnXK8ZZuWbbYbEe/UAYtxX41Zi/X8FZkYGWaO8QbdmyEL5BANO72gP1UU/TQM
rL1x/92OtvcefAu+FNWftPySx0fsFqwIGSmcZiriBYBPggbEbHbe7xt1D2fDFgkNq3bXZCTvEndT
dcj7NIM6n+zA3I8aytmZsDd/4yziLhbJZS/jq1YpZ5VS+tWzL3AdUETLithONAoX5aspE+gQFH6c
7bG+aqhBgdJkFVpy5N9QZpS3/cJwyh0PASa5X/9rDCpBQJ6kGAMe3H786BO9QMyMPy8LDUuqp5Kc
RPQnp0Tj532zYOUqbEjQjpxmuk/d/K4I/KsM9mmfTd5HPKplfQxSEOuDpLiotQx5uMKhYmOH7g0Y
zBhTLbFi71swPahDmskYVHWBVFNoBzt9JoMxyP3MgwieD6Ozvmd2cR0vfIRjIXlTVDxFyMtvTQiS
69KEDymyQClpaj0dvWsKtNEMhouMyDpGuAZCmDIe3wAsARAT9T7pNo4N9HJ1VDYGeBliaauddiP3
Tq5LxmlpEKB/Fg928kjeeNPMgHw0our+Sgbd+MY0jnNd2M0+oSblbXN6j0NKWOXEvD5N/PcYPBQ6
kGbLMdCsOSdbXGCAbd3otqWYowfIwjNwPzPBFaz0NId0W/D28JWNmJE1+Hbsqb/QRDJgIoCDw7AT
pp/+7puGrOD2xbiCh/sgtqp5bT+QYqn6BZejpqIt3WfSKVyGQ/RZOuiD/wBn/291+I/9kYFEzvv6
Qy7l9ptyb5G3H9R+YcjHsuf2+9uMbcKANWCg19qt+6FnRQj92cP0Hn20jVpzaTMlauyQF0upr76J
RgDGHOaeSMKwA3xYW1cOrqMrrPDsGM2OwRPqg0hduBsgpnrZGSkYQ4FErbxBafuWeAlKVHLx/cxS
5gI7y2HrK3xtaKLdeWOcEJypxdwtwGdQbPOl2rZOtN5QPAz4+nFtv379OllVVr6Qox3i1/q8fUuK
gJcGwEHU7dWZjY1ZMJccz3GBH6hmY9mccSrsso68PAIC8TFvKID68IHKzxrgqlBIrr3zM6p8pmon
4ybij+k13Cl1XPIZja+7wmOuXkpu465sq0gseMNNLRHo+XbItRZ0rrY+ICtEGDHioIo3J6IBpbNq
M0CKy/biCFT30ODi34aOHh1bGJ+A63dfu1p/3HkJ3eJ53+ganSsYa3Ashjtwe2b3jhaAUx7tBFY7
f1plXBr3ftG2JDHmAHX1gzHFvrRhY3JFNHwRaCd2ItwwvgTN+RzXmGT9karrnpUJB7sFXaByFona
hPfGcqkozgE2XutXZv3xOX/87qovR2a+5kui30eU9zUS8X/sQAylbFFMLblXQdP5g4V/JJLkN4Hi
i3/Zkats4EcXgrtZo/cImGrm+uQKGCKN9PSCZYdhmjbK1ttyhEY1NeS0+2K2kRbnVzzMdoAk/vZR
WHeUVM/KBCsbFBCkyjoULi7m2oK+WwJ8PXKbInx5BYYPDI3jwGmoLKc8xpfMFhhon/oSsTiYldbX
VW+9e0JJlelB8cdtrXn8detLiVlcgHuHJuDpC8GfpRyIYUtmzh9KLNOcMp7WI/C4E7LozFPepGxM
xmGy3NLncmqyVxZHu7GkkLifQILgQV3x0CqvTNbcrn74hSDNhH7uU2TNRChxpPzvteinlXcM7IH/
regzGLZxgrbLwxG1QhMNfZhnuyudrrO53orRXyFEKxZGFX6tDFZec0vP/PzRFQ6UeXKVJyXIHeBQ
LUbPCMcMvi68imEsWONYHVJJxxMZvF+50BMz11KZYAEfIXvNGJi2GuOpp4Ixblc/prAV1zBHDbeD
B+eGKxYsH3mRyEPJKpXwVbPueZate1/OKuZAw4fwyEoXQWHSYzOmlJcLeljyQW6BHWSB6p6lkO9d
bUFc+4bfF1AyulstQBwE7G7kXDM8GY2CBIMg4cwar7N3xQc1vIxXqk+iQNsq7zViwKBcTS97LnEM
3WcEGATAv4fItwyd/+1Bg9n2Gjkex+Gm1GELl5+PcaBrMVGu6RNJSIRFQlzYloPALrZfsn20vOIx
yfCsSANixgv8sAZPPGgFrSik9p3RYrYjmpHqwc3+39VNeKxAH381lOJliAO0mezdaQiSDlfwyj/g
VyGraz00jC7yPmAdDJCj+CtIfv2DRwyxpo5gx02SWW9eewaJ3reX6/A5J44RUWIob16xWjFRAe87
X7YixKujTW7u6CNH6h2Rhy2ZS2l/gRvowCqsXqIsZk5RTzuOwAVaV1aqxPGAt5NIj8a51mtj2GqM
yK7DyNVef7ckGWeMLsR2QgLmJ+6z9P4dPSSw3qG4kAD706iU0YCw8UIggxEeTG5uqL99dtfS2kM4
sXVUlV/In0fYHGheDCqdRZC7JOPa15/VfMe7yogY+CHTEymMFeIr9vfR6FGxlbQfZR+urQERdgXH
tPIynJdCnj1ryV6UZkbbaXssRS/81+ufLG+jhwgz6aOi1s0OVfLPqMBe2ef6Grv0AP7353VaW4xz
vq87b8RC1mDeJ4YDv1QSOWqGSOxc4LHBxKMQ2f5hwPKKsoMrnLirUSZJd2eJnN5OAtSDqobl5WPv
+eyEZGGItqfXYgtUwPXRJr2ttQoPZ1xPl+0pWd99w/7f9+yz+CU04TW0GkplcmIxqHZD4ES2Gjoq
fOZ79PZl6ZUZ5GpbXrn0HYY2Ug2m1bGel83wcoMeeVn0puyXYbm6698Tq4ocrkPVCopr+lPkcHO/
6/NizL43h/hVO0br3FXygJyNFGbaoIax4MhdRpJ5foa1O89rWPbftpzR+FnXzCtPwvoUchUblUUu
LohRYUzu3VPyqJIT3t+VnSSu/QVwtz1fY9QG+3/TbMmMXNDcOQg9vdgaGFBt6jW1pApD+cJ1dX5M
+lRH72A4fSHK5uXnS3TN3tLWpG8vjKcEoN5qS6NHkNyPEjZ+Jzcy6CEIZ3Mcbl4tD24K8uzmmoF4
EVBqbFfUWgzTSeJ6zXtFL1J/0iaTGnV3dEGfAaDMbyQt54aGkEzMCB0xJiAtEx4SCx8sRiOxTTsy
1LCbi5kaSa6ZXof3AI2TOr4uHBfbXFL1sYTsZgsCETsAVmJBwaFlLHfEaUb1aLiPn1RWnhk0qdCz
0sRslh20O+zK0l8AuAiyt9l/Gk8szDuLOKwmyCCLyQumNhDyvQzGUuAeciZaYypIee9BkU/mIVoH
zYvKfwj7Saz8sSFaeUuEzCN0XKZ3hS4/RAghqD67EZ5uGyEJwu5VmcSmParOePhDDSxhbrgDEK+V
QsVqMoJealfbV7JNBKmiu4ZOiShRgU4K7BWjmS6GZv6McSuDI3pHuFir4L6AldR6Gfh+VIkjjdyG
KsWyIESX7pbagWEyKFJOZGsLbIz2GDWN2jYVEUrs9sYv+gfbFUXBg1gknXbUCoq1SggmmvzY1boY
cr8lEhlOKFODiKYyNuqeqQrkKwHCzF63qf/voW0iAdsDuXc2hhcXNlwq8cIARlIpMlpEMyqJl9Ms
mdT0AyFZ29eZa5uTLWk0dwbi0O2EP8LTw5aXqBRyp+DZd60BB2uQM0rmYDJYs6Wzg+soIpVBg7LO
LurgILtN6wAR9Py24R3E81bHFP8P+/2aAIa8GnBX5ssoPK1qmfts0UBnhqg7r+7vNE5JOkdRLIMJ
bkcxOnkT8BOyurXvaGVF2rML1bobzNs0ek9n7jBLH8uenowLzEF8D68mvb8SNhPP7yoiFgP0KZXw
zmCJlAmkaJt/EvUocOlOrc/QVsrMPrlM7rHhjuNzLU09GeRCAzdk9LFGN2cn2QTzURjdbWafVNXn
MiniN+UlIVPnp1zIws2lK/88+aT5T582aQlc2KeCiTis9bcTsFcAZ44GFdxK1fmksUmWjTeVJTxT
aHWMUN0/8PKE8l/RAksxPRZL7exmsoIH+bLpRmKY+8t0agfxEpd0m3sQZjXf+zbYb0bLKN7yX7QZ
vnY3c+KD4zrQrYyCCG7+KcNsGNYn+q9XCxzcHqEuKjXO6/DZQI9Ppj/RzgBQE7s8kokaLF1uc8un
/o6UZDM7GWQ2IAaXrP6+rFGh8HLrKkLh/Iy3YJcKKxcRsAn1r9jttKyvPXw9+els2mtKXLDbCrU9
KNac1QRx0c4SEZlT+nFc1gbEk+ydZvSkWng3kUDsRZh3jeBozfpdjQKwV5OosZNbWSixo5DhmDKj
WGokPg45s2Juv4b7ke3V+PW2lB1TaS/1qhy9aCSSi3XqhvZfHyfB2yJFw23rJbq6KYuO9kNbn+mp
zKGRyY8fMABOyk+dY5dKze94emHHB6z7T9bH318UqtcIlLccCOhDf9UhTaQ3vc0Ctda2VK2eTXtK
RjJbpbPwJiomxmBD47fkmy9rFPYWL7JO8HCm9XYw4Pd6N55I58/ZvfJyBB1Dc6WSnIEQQpbwHphu
turkdnex+kYDCFDONCfabrPJu6+sYIvuWAi3PUkDDwWkmx7mv9VIEwWTpoGWetojbK5c/9C8Ji4G
KgZIGQcRNqZCrzXE+1gLY9qbdVPjrcvIBArAI7WwK170FST6jH2Bg16UMWrTb9RbXVGojllJ7uwD
UYNtodaRC/Apjdn3gEJ69XWJ6teL2T5xS/lT5kJcFHJ0xiQ4loiKfD0i7+tXluRdAP23J8If+CQk
c5QS2gdL9+DoijA9EGCWin0TmI/vGV7Mma8m9zaUAgAva00tajSRDzeSimxqcIi3Z5pyR97lsUTX
zJM6Xo8vLuMwKQ4N+VD4Sf0rSK6BjY5MeThQc61oJ1AsiQF4fMZukXOaIMwimmHF8VxV+bQDSDm9
SA0Kff0TGsHNHD7KvLzYwnmSRM3ztDQzr08+5+zPdhhh9rxVmYdf7CV3vjKa4QHQR+9rVmy+IL5L
JoNU5z9PYaEo22z82oT2m4ZfVYZ4JSGL9dEjeH+uWnA/g1/qs8rgv57AV0hgD14mNbss7OL9BS+q
EHZwzJ3NGXjFsfGKUdQGPps2Dax85kS54DIus9D7T6LBnCwWVV6d2J/sceyZxB3t47im3/XHzve8
mkjijLlzXaPKifuPIPLn/7VieuSyfOR5HEVg628BQyndKIVY6M1cwV3n5copSqYjOnIoNfwGW+oM
tF8213dqWlg5LJsusJOFfXunA6Y5S73AC2UYyhhI0idwjHu+xBULTJzSPiQvm3h52UnJ1eKPtoHC
vDbDF4XNsrqjX2QVmwpVUbCrCEEcJOqBQ5B4c5byovN+D4frHY2KApVday4Fe7F+pr7vgCe//9sO
WWlk+loQpkBw+dGna2HUhUN53OCwvVknJMUfpadUtzjxZcQjP9hg6qlzAbKbpXRvEQyCgSbGrFGX
iqNSzbnb2W17XtDT0yWF2VWztqplzxd1ZupYjMhSA2PWt+RJwRhEvx6zGBwzBZX8z1aoAkb8aP/w
CyHSXZ3aVahe7B6dmHhcrRDG4Mb++yu3THRcBYpak28R3yOL9kUlk5fcEelJSLmHqIVsQ3VZGxCT
MFpi/1DcIJ4BDNP/VbehYO9kTGU4wLhGmJmorjLdeszqaQY4o71CQfAT+FLylLLaSk36xl1glZGG
tRd43z46oudjz2HOFOdcFvtngSfFMiclYlMiKfZPaj5qJnWZ342qDs/+XHmuFIAXVXs2LUQdrrQi
rLh0D6RYvBSmEyPmRpHRWTG1cKTUgo3hkji5Jq2OlJvwGzUEpRd0m9zLKDWlV6iJw5S047l3foks
R+9Co0oo7T9hI5T+lcokIOeXRIKCb6MeGUcVyT2zTPrYxsI0LF7gZshQuuxhQsuB/5CZhhaNMcQn
JWsvBeVoAXPpE8b4CQ37trXksqLfDDopSkVf/bfFVOtUt38SkozF18nUHBSlwUCICN6jOrX9ZAkW
i3YdC5zIa7/E8aC2SrY1I44fudZPQk7XoC05IX1wgbyJ1ue3lERCdKZ36GesDhIgXMroCu6S3f9i
SK+2pO/CZzgduGBHpIXn1xuVr6d4jqA4S+EwT2ncMJBo9altHPSwboSdX0MaFCZjxlEsulqLxpAv
Z407eCBAg3kOLCrSCEnXp3CSSUJs6xJff/lGmDG8AwHW7XLYPaeiN9fqVVdXXLq6dEX3dpQKlsvq
fHQ++2Bz09sLWKcAtn6bOsdZgSaAjHpfC3I3Ow3nJ6QUc/yeXTpRg68Guu8yHw7lsriI/SMMubjk
42lTDJzzzwBJL+r+tUYJn5bDfDS1d/PFNI85X02ovTmYAOyAmqPHbcCBjFF/SVgIyfMat4Po0T0w
TZU3TEGzHvTW5NNKmkXAZUEQkrx+wqlcftAJIb9A3UQGJUlCe4IIKe3ovctw7R4zK3z2gSrxZhve
HKyX9TvkOXiUTiHs6NEdiLqZXz8Dg0DoltkDy77S6KrAsyleeI+JgoAJoqlZ/M4fdUwdhAnR4vSz
mzs2N06tFz3Y0sO0TN44swD3SN5gNEje5hXsUAUINV5uyEXj24WZ2Yy/B2wlGyFWQwatzW6e+wUT
r0ACqos2Qc9tPCA5ffGZ7Wv5HdPNJNWYzKMKm6ty9Ra9gzjpICulY12JKT+kKRM7J7ZZQy0zt1tS
cYT8/Dl+dgHGx5V4mGI0kViVoKquIRIMVgC0/8cEDO3pvKu5ti/u9lefhb3f14W8ga22mDowDxwD
9SpZzRdTACsEP7cmmPPRdCzO6EeMbHZOxdO0nbkV9kQdihPTenS9AKlvo3NBgW7AK5Us9LPXQsnJ
wnYXs1FubEHyqHRH0ZGVCXQDw6wk6nhGJLwO5obZ44yMqMbK3i3VxBSld/Pb57QCrCGBfVrn7xD+
HaX/x2Dz97O4sECWVIMVpenlpqFQlXCj6vw3o0JWSNae4GZQo3Hoa/Czx4QChZ2tEIFoJHo8Aqce
Cu01nUlSdp7BTe0ur7dBZxwmiRfjPwcoDQ/GK7iHRilB0DLtQcXRhe+uBSjrOdHXK6aHMfJ9ABAb
x9lMvZwwCR7ZLZBVgVHJ83oonjaibOU7DErhY7XFa3e6m96pxC8vUb+ODgdsrLA9Liscza9CQqw9
KlHXcJWzam8iHzpT2OH42wlTZmCniEbiAiUzKliJKtdpdKmKHXIFHgKFxRp3aGk9H465Iu2QzYMd
AUS504vy7Vl8C7GgTyXocS+Zn3ktTVg8JfQuyqug7dHWA9VknlPpy2NaiZEwNcNllS5v4FxghAK6
jrGHfXXBUQhrh2qa4vXxWtTA6R17numayIHfGFaL50TM0uuGkg3itrIiqNwqFguPzrwlYpHSJm3c
1NdSHrrzcyQsoCQffKfsJH2ZjGCmHpZVHpge9QJK5Vnp6n5e6Ui3s1YjQanM/Q9n8RT86V6Vk7o9
tH4bpUHER/Uv8ShISpLdRtrFh8QUYpVn1rpsqUuVSgrj9nrUXhOMlIi7oFQDHdfr/M8OBsNIXQ3m
pFZrccc/Hhgzwk1JACPPgrh9s0nxpkQcH48PFiU3QuDuc3APv7zS44Rnj3DoTXGukGNZqYQikQwK
4ntTP26oUXytkCkz7KgcCqUhrnDjGiWMXsQ6/LWfB30/vrfblqPvxPwBpGD9srFSf7ZiP8a/FPpx
2thCEVxhk5ijnSO9fs3B8el9n644sx0cqeLemD56fekkFJDW84flOCAzNmKi07NZca1r99UVhUCg
vWn/BwjfbuJIQDzJZpmnEAZsByXB3Dsyi+w1pCK59GSmiuwSwDPBL2B39OajrGZjibKXRCnYPYO1
yTE5uUVGocT9bkED9L2HuegU3FcUlIG8hIu4CZwhVoRl8nh7aUJoeyRKcJZjHTVZawXGy2mB4CM+
qKLMNpWke2zBqDgfYFadwQP7fcw7uKRsbMP3OSdgc/kJpzLl/EWE98QUb9sKH5h6U8xei+6qXoX6
F1YRELAsK/CwLOs1wo/2ft4PXJ8PTjdmYrDhZ5qa1NlYFmQSBlHHl/lcfn/dQFZXBx+N5TbkcrLF
yMH4nQW7Oeqk7IEmoDPxn/K2EvHzhiiN+wIPUvarJYAUJ856I/YdCNlhb7bF3TLC2N/ksDmPJuRQ
jOcfDBLjmVQ2V1ketCSo100FrUmS4U97I3d9EIGFXVSm7XjBYGlNhZOK1Hv/IS0eWxdOPKbwvFCH
SkVvd+dBnPX4yuwEgIHKV23I/zXT4G3LvTOEZdERL3HiSgu2GBAZgt0Qzcmln9ghetbrzXAQFX9I
LT8frNqUpI9eVqLFGWw91uGtrkWQnNiwQuaQu66aQJT9BFdvq/qAAiNaP+2TpI1tT8m4FIFpSaHY
cxbFpFRkEMDomdWHN2N0+B7xoQ7VEYXxohvdJ3fTClFUJqJq9/RDSp1GRDLIPMD1pysl8oLYbPCX
pLy+F6cMwtr2KLjikRmxqwMmDaxUmhvKfwUrcEtZlFFGGIdPNFN+d6VOi8X+gqjuzRHgYQyU1v7F
0waDVWBv1s+QFID7k/DMfsXRkbHYjuis3mwnPqpCdRlCrYNd4Wp7XVP5IH+rFKNp7SNLGmhexdvY
VcGGc/ICgpZ6FH4CKXXYe6R0r2GpW9KadmPUplgnxH92ljbMX57iaSp6GfJxjZ5wNiycr5yWUes+
HVaPf8AwfDvHj1IRvzReoNzvWOfh4k3+sP6KLchQy524q45h4ZIL8aG3gEbKaGEt6Rjg87LEQrQ9
KQa1jDdycmDi+YV4Vb4+yrXX5Rib0Vx4MjAcLJoD5R1QdRkKa9T5q0Ymv3lBYXq/uk4QaB0U+je5
L5VeezWVIRL5Ob6g7OduMCObNXewWqD6fOkiSp3gZ/lzVZY4ustkC7uywqxC4s2b843VIVXTZBqL
1fAMPAJSCOwUg8OmjC1ErlOfs/0xbwVEjih6rE+L7KXQOsnWa6TAXgLE38IUGLXd5WlpXD7MfalN
OQ/tqrDbCQKIMCFtpGOm855jaN3czTXZkkz9C0DbnzZiLZgcnnP7Y0AZF7odGITa/TrCB4cg8slJ
TqbpkhoINHD8B9e5K6aLjVgXAux7ZygkFoYzD+i1gxUXGE3OONfdjrDjUMTkJ+O4Meop9F9Z1t0A
nQ/jbxcywguvj6Ko7zKDCYkUMYbLvy0Oum27L5ANt1U+KPs2HeMhgmIqL2vtjq+fXOjS5GCFwrNX
ocSZUEOuXlhXX7A7Wpvqutlw9gbGsyPQTYW5NbJa+57AVrUJJn0vJVgxGGsLwLnfWyahzDkxIRC4
Ay/H2TWPOL/vASEsLYEySZBj9JJmowVTkUQKU2xR4quAeH2QyDjeovkYTYi1UP50k8T86CLJ6HdL
fdcloDSWbsw5VngxgHKUzeL7zyzeuHfHC8IFyIBdMRcsWcyZdHiqhx3/pBkJjU20DAEkukII+QVa
pvQvLWQ2hEHSEa8dc29ULj24zoMVSo0FlO60YRZvUrpVKZhur6L25fCJKSX++xaftyV9g2Aj/9wi
aQBip/H0fQ/SL8xAb7Doyp0DMBbFR5t4tpUgXl6v8/k3HiHO2ZRy7ai945nqOKWZmHPNPazVXF9b
MYkNsmdlOMH4b2cCsM44eepdn3T/qMx/HbaURNYkSMOFJ2Tcyo1EBbOhmghS2hFMHX4bfMO82sUf
hw618POH0cu6aoisr/xzAOcDzZnuHh1g2I9mLpO6++tESAYTzS1d6avxQepz/IRH/AnDx9iISWS2
Q0NxiOG4dCEWsRkjy90/cAHOBZIghTAuk6wq1PMDWguuLa5O6ngqEmapvA/+qrAsTQ+SDxd15hxs
rjcN4xjOA7X6NRZGd59ABmcCw5M5vUE7I9zv4ZRZLyqIvY8a+4UIq0jvwaSucGnGAsGmwikO8FEU
GmBzt8zCm7MdlNDZxMvLmlxy/yqLbkugkamg3UmK9YwFC7DWYBLGHWx36JqJ0V2/dSBx9JqiVWV2
k/wAqKZA3t/zG3x6XTgLEV6187jkEReMMCCcrUQcqlbZu5pDgMwv5pz3mzMTNcW+ePkpEuuUj+Nc
FJ5lG4/1y7xr5ySn9dkcW5kzgy2977TIiykLoelgXLL97vHxBKbiqgAgHup9q5pwSA7pgGz8v+IN
0MVN1wKFl/yre152NN65pfagB6NfYOlK8Damo/1/XMfJwdYkPWy33qHDYyHe2ANJPcEGOilEUxw8
YxmX4uosPPm7+lcEFmFLsp7B5Gx4LNHKcoRnjHAuKdZCuhJ92i3xeayeOKwN1oELgryZ9B404Ja2
tswtaej1gdc6xDXEQm6S06QyzLmPbU6KOX4zHNxo0thn38VAe2+nt6yG4d0ctNM9qEg5jgq5n0ZV
2dbh2QhzWNRhjqZjy/mEUz8Ik9sJSRgAtbtGvVtqCSvGT0d0HChbg0/BJY0e94hkN0k1z+uwsICS
O6ITQvXN9wfkP2h5GfVAYjTH24LHnIFVsUNHSZkp6bgc9SAcVDpamC7Y3HDYTjVBCo761s53MsP2
0iLOLlcidM6B7OkC9TZC6EN1yvXWIbHQ5Q3xowtlfmwEFE1OBWPXlfXdA6PVAOgZ/X4swWa5tDjN
Ysa3JbSXXfo+rf8hQZCNfP4/uv5DnvJX/p0X39vdAkb6JTGQA4E8efVpdAAGYsbJ94L3ANynONt4
tNrPcSIHWZuV1RZPUTeQjN/I5seZ5JI7vUpFLRpxL6yAEfqMbisjql0Pt1F1rGCPmrzoWYIwlJSS
sh2hrLa1mSPlMzINVINRXNdwD5CtA0uTXUnzji12gm9iG9xaBeWBWzJQyXgs2ffxCv/vsM3ukUrq
BWQyXMj27EMApNecs3OvW6XBhQI/8sCXVgaEHrv9TE4yMTbsx5ssHPeIm9JOWlltytqZVGY/U99U
UoF7K8/tqT74EajUK85XmRcM9VOp4YP0Gj3lxu+uMh2Zs9zEfgMd5g1bQ8Qe1pq7S+92dkCldYOT
2EMRfn3jA20xZiIOZb1DU2TY3Wym8ECJ3Pun/7sS81RYbU61vWwinUDmg2eRIvcOwQim/ol23aRT
MuxP2mp4+A+MGqgIGFTXoYejsr/RsScxavFqL+RbwqCqN3CQ85P2EqdkUIIxu0By1WBsn3leOJhx
Eet1A7gjULqg44O/1SOc2yzqXYrdThIuKyY9XwJNqIVSxNkaaynanGruS++qLYXe2gjhgFQTp5rT
TX26wn7j2KYdQs01rIhW+oWPYPybvwgDdOn0hd29pPcNTQ7ncMnQiBk6eKZoUhWdnkijp96sB2Ch
Mzh4HPF+z5y6khhv6HGhh/nfww+vEv0kczEdcFfFSZ5tT95h1/AvLFKV+uHqZW1SserMQpof4pfa
k0sFpAr/LwyqtsPnOFGuFzVOw0P3mbSVSZRokIidfM6V4cuTbgXkKYe8BnlCu0472hFtC4wgKqa8
4jiJpAZDcT9haDGSBvv0Zhrgz4vXfXqYlO7bCwD3OL/Xe5bNCI/UC9cOp8NEYlX0kBM9aigPxgcP
B0Upy+MLpQGMd/hJZzwJJzieBzJ/6kJnAtm4h9DfIokhi9Ug97/kfz9A1lWtX8r6s3jzoJgSXdQv
WZoaHao6iQnUYTdjdm/81c9EVUtRJOhLz5X25SCWfo2B9hzPq8MQxzbhwfOhV+6ybz7kjEo6dHd8
62kEJMCu7w/0OuP8oaF5bcklbnBykfVUu645WzpsWE7aRtCRyNShaynUf6li9Rz8aNacItsvtEsV
8nmkPVPL98nuE3QGGZFkz4AmOCcVHrff/zjFAk+rEo2NQggeq/zZXiDlcuZMvQB2/rhJPfTimcU+
4yo2KC4ybHPraxYV3BtSHuUQWaD6QQaKbljN6vnwar0zwGc6JTzJeYZTQxNF1g0QUMukq0KDbZkE
cKhJ2uJH9HkQu1M5/gbdEOMHIAyuYzzMS9JGtGZ2JiIAOdpFOBKQr1QhyO1okCyVnPzKvs5IqyGe
hXAH2a3fj7LWAjVREl8r8J8gN0ufPfnzK5HsJlSo3nTBz44XYSwDqGY++URVcWBAxn3jqxaNy9EN
ZItjNyxbaYA+R4Tw3JkAeBfwL4d8yILS3HDk2HMescFAmltfxYLOuRcOgfUH/DPCtAQnFFlcXZrJ
TKP0tFYxEPilcpHvBlQX0qlXg/xG/pgAaKoh+wxRbXbJavGGj0d/sjmCmhZDr21bRG10ThDib9Zi
LRgQm+AJDfdAHBjgI751h2JLrBebg/qWGdQna36fUtCufJAVM3Qzlsr2Camk8jv3lmI4b174HNW3
H24ttXvziimjxc1spYe+lc2Ol5Ly30Bvz1ub//o7zyPU1qtUt3ehlmFNzNQ4uFVYvacdJynL/NMi
WmaBlm58pC7NNpPf+udV+Ny8QMWDfFx0HV3mhOuSFad0Gww9EKyCoGss+UJT0pjgPRP9s5PWB/Yz
VQbxOLj07AWUeorjfX1NRY4mYtKFMKx93vTeFSpEMn+GnM19zEkxMtp1b6hMjZp/v3G+2FfXbA2b
aT9neJ1Ak3ZDjXij6RGXuJKoE4Va2H+trsGeAqk6HgbEVygWzPCl7B87VE5StCFbjnsCxngBbZzB
EwzJWdk1BRyfmBrjWlr2CAtdRq1nc5bnqq5DuB1+RxU/3S/8V8kXLCTSpdoDJ6KLMkarAFLRpg7q
iJh7KnTie/TKv+rJieKG5HvwnFyBFg9He7yDV1mvvwOFw9fs73htp/fE8R4aWQ5yCveoiqZZQHog
+wf2DPHMtRTnUCU+0j2faw0ZjFeFg+aTT8skZWdr+QpPrDRa1FxznwwvkVlykQoqcFZ6/gn+uRu0
Qtzam6MxDho3Niqud6Ay5/yu2PO8BcsP3y3JR6ahol9wyl+AvFwhFmFXRRMGuFxG+GOj29kuOcgK
1qXumZIF3u+i86DbsGxMgTCadayNTwMXjm7N/GBR9QVn3DdC5qeyKuPWtHUvPyk0gf2HWda2bzSu
YFnoE0qieQ6X/qAHlehurnKmlmklHE5Dbqhg0ZbRHXiDTMp3fu2qrOGIXnBL/Iy4HG7jx+wdQ0+9
DbeXb/evu6R5VAXVhRVSB9n8fnjQU1I9/xqKtMFmZxbdROiubzIpzyr1DRGiS8LK3ACyhr5mYG0w
/QWEtjIASwbZIztXJMrx4YXkQrE5iv8ALPtp7uAzMwL1bV2zNg8y4P7CUCJ3XewFizVN3XelzpFZ
6wHW7tO4IDkSkBsUkvAIuJOiBcHO+/onImzIVzG/Iif0zYcTy1xvA95LQBu02ECp89bWqKuWK8Ah
efA+VyAEVyl4TXOH1kXOu1Mdl4rv08klz2V1AigLsWyx+O7fFgESuyxfcuWGH2wm7b+vSeq2tYO/
EoYyuGwTUUNOBm4zNo9Wdh0LSwwJsn14N3SsObppXgUtkojDASOI3gQGL8+lVlUusONRpIP+gDZL
f25PRXeKkzky2ZajU5KD0HKz0hsLfGuRGpP2dAfRX7tJyeSE29jqW0sCLt38JOHYFNhT79jFFPDz
PtjL7FK3L/CMpHNb2yxVkk5yDrtxOBAACgQzAAv/cGM91egXFUUomb7DPD15PjakduOel/c4O7dy
xpL5TyX1zWp0xPze0Xddq0O2R7WwWvbXxY3ksDeqYI74T/8Xkdt8JY5dNP0ajPA9TIDZDWFAiCb0
RFp4NAAuOm3ESppzsEAkhEqWe+CT4G4ZyOV/+CiMVQpj4P8n96IKx9svDxIg/u7zxpOl8VL82QYv
fbKq2dl18FXZTlytGn5wwzWyJVi1X7KPlIlvvhQ07+m41p6+Bp5RSp79svYuFngFGlXgrwNEAT1E
AOgCjwE7NPhmdve/p2KP5IpQy/iAvUSpxh6u67povBTo8xDCpwlGNHMP8kqmfHk+jmUKm2rH744N
DLi9QNQkoZMmNFCaIOTOpsfkJNNFEvHgo3/he2tJXNC8TjejWiYouZkF2/CH7bYJfm2N0hbbVMDw
lY/NT50tMzZP3zT6kjA2yxMSapoiZdScX36kaJOLc/Cm1dTWRDHutTaVHQMUlzHCqnyzoIoeZm2M
cIyYqywOmNUptn0CTNiQpHDaOZRTjorx71zAENbP3CE4fc1PmtmDoWE5VKPYSDkRK0N7/Ckn36Y2
8yIruMw2JXtmTgVo/y3bjsBifo2f5Li4mKvIypfI62Yiz4XuaKaGNSw8KQs/a/f9iCKGRYui7WEl
hgtiXruQcNiArgNW7bWoOojILi3wsTXk3hoRJogBdPEIxWJO8IWWx4HmiTdkPHB/qefArAqIbdX7
VJAL2LG2vYDTlPrtvtGYOqBSwrmNqWevKZzPa7TO2qGyk5fvAHw9IJU9nxW6pd36HgILvdxaSvVo
n70ocHEu5M1+SzLAV32CS231DDWIejXdrnlaTTmCGGQOTdpsmSBW6CMBrWcG5Um+Ieka6KX2A6bz
2RzGaVHL32LF8Bvy1fPiGUTduR3Jbw8h7GK49QYGMZD8rSp1ZIWDBoyI/rDDEpYP3X8YbcyR4D64
aSgDphCpWpg55tS3B9poWpNxxMhejdwMk0dJEVkhaSOhPXuBwnmED4YsvPbtYU9gldx+nZ6bYtnE
3jiEuIHdrHYMd8x0vfGd6ZesDzP0V9UQrVmiZgUTptDBgUXN37LlIj+CGoldG+XiixscmW1PYQem
3RlPm0v5dNP2+wHlkTmMbNRDSz0CNIy7de8zvYqw+rthcPF5POp+1QodZNX04YJwjCnMomSkIDHJ
8xBIdHCuOLlOHZrD5VfVOHAwFdgEOKYfJiFvoBJ/67YRO+VXMHLvz0UYAL6FzmAON3X/mj3mvbaQ
U4+duaBH277V6m1y5CO71p6E+PiBCE2QIcqWiCPcpn5VFifdzWkq6uLONNEtSoiUZ5dFVoZ1PjkU
P1gG04MCxh2vBUxsOcwk4NJ/IZMssR9JfrzP0vNdXjfr7l16IWZVWI9eZf8dRDpCHdpSznpqsFRI
7tYGyzyZoFZ984W/q1VnijVo5A1da/Wcj8m3MGlAty7Zvri4aCwa1vvtYr1qYaJQyW62rAmlFZhf
qmORnI0QdtTPw9ZoiY01MzWg6YKC9odbs7BPdhrHu5Vi1JRDmvjE9d/F+2oGX4hLe+e6Cb73EHut
5LkAr2otxPO0eo6UkvPVcQE+FqUFcktZ/kmD+EZ7y9ZOxOr5Fl/HQFi6EwaSxph4dhoeJghc6R87
IU/CRTkc50JkB2ADfyiWk8SQJMpc/6lpz7Gl6ybx4WfgMHSXMf+xXzTT4RpKGwhHMrf+v/cRoAH2
K5IO0jEBzP2nZmEVZE6gej/8HdSQsFSkfEa0GyTcVu3+z/Rnwu/cxFIwXuGUDfFC3iE4A3jRQHZK
Ex0eHae0WYX9s2BP1Zry8ErebEraGKu/tUHiy3AGEu07eagR2jAflvRFeqHOq6giEcpt61v29yDE
v+7TdTY4AXun8BhUf4f4kvSkcteoNHI4rOlFh5Lm5kwLgUb4bgpe9XpJwlXvQC7fnbIpKalepi8N
zKjJK2dtQbRVGZOOMZKKO7LWD8kFQgngJ/SGokibLcJGE/Kzjd5F8kty5zRBFI+ZAujeZXN5UYRM
ZS3K3go13VqwkK8lQGd+4LLGi2t/9HSxZOO6sg58LuKpEaq1nU7+2Wac00yrfpCVQv5yfZTM1pSl
KWe0OOEuIZpDaQ22go0Fip2dy8Ky5/cHlDDp4nTszc+Nbh6VJqsdvwP7iLKfDnTXJMnOLAPuAgyv
SQuhFraqbJb9iD4DTvZUt5qyahR9nLNLo0Urupg1tFTVzCpOuA+FR9jBkNCdtHB4sc9TfQaalOx6
AH0A1XGhpcpSxtqCJOiofYB16Juo3jzwnDJRwxxcBCrbVGkUerlboIbwMdPJ7oKMyJw0IrPYoJbs
pfsj4frctdjxLXmYsC+uCSLxSPKme4hsAN4XujDY8dZQZgMQmGT/+bEr8iolhaRdTIQmgOpCpn+M
3UPK09SW9GfNlUqF2FQyByWnVaA3OiMt34+pp1QV4ByTBayH9TobHu9EbBNyb5nnmbzAe12afHGE
6HOYlOGRKOLwaW1c6v352vZ0jy90OsJSjl6nVfCJ6IH6X269vxDVuBoVGxqGOUpcyGbuz1tUIqIF
OZqk72S9gH2myDG+iBNg7G7ZrkRqKhIsuvPbvmbxp0UAcchA1YvhCTPMNGU6WEk+iPLOaDiqHkQU
z+XfjaJFpDcKKcJWMtFyvAeIPahgitiL+hwDfZfhYVPeULGDQND622DrgdTycDqiPTlHY3F1XQSk
ho5ZCEdeGFDDNDjXSW6u9wB94l91+jtUHiOf9nYz7vMgVOeAmv+/ecHVxF8NCVwwFjYhyx2ljhjI
TCARxq+kfASSFSWbbXwApA0CYrS7xWzt+HgqmGcOxV++0LXRH6aLonkVdnTpUTcG4sJZehQ3et3e
dRn4tg06yHzridzBn1kJMuOMtlhvlgEBEMl3smfYSOzRTK19Coe3QLQt5VM1C0zqirYqyLsABJ2h
mi+a3hmHpRpHVjjVjy8hiBmqJALfbB2TwS/h5kg33y4DlS8q7aQZN49S/bN/GI/MrQl8554Q+HYM
u5N0xQGHJiV4mQCWoBl3QHF5h8laSt/GN1kAla2t6tzk3PZSD0BfSY0gAw5zn6t7g6lCHWVX/eMT
j7hUSF3s/qO76quoXdbsIQwkorw6TehUKPFlUSzSgGgSP/Ln7jTc4qtSLL2Raki8xmlkvURFzzOW
5akxR8/hXwkRyh6/bc8f0Lqze/2hCxo7AFX9XLjkc9IBR92M38aavrYv3id68B/L6y59M78oXSN4
WEgEnIPQDwfhGLJ9JZ4zZIyz987jhBRxOGKZLatWrCK/JPY7fFarB8MuqyrYsLsMB17S0fM5cBHs
ljRAWS7jTTlmG5VasWcJHZYN28ctg0VOtWBZBm0E77CVKqblHXvRFPICbXHPibtGiOJRbObTZUXf
MCkQr5CF/TiqcU+fKVxLw4QK4JsiD4gvy/1HUNvaQRKGYo5PW4uZxR25+ESMcOypWzbHb/iNv155
VfpuTdTw2pzlB6dzLLKdjMTkLE70VnISkjUHZjrYHgkG8602EoHuIFObOc6M8bCLFWSgzsdt8FDc
Hn7N4cItp/rOO9vgbnRB4UPAwUza0hHhSLY/gmTtCJZITdBJDj74zzfntM7e0GdnqMu2Quc8ytvq
XJq1WYcFu+ayuEKjRvnPZFJdjxek2HcZ3yUubkafJvER+fi0DqAwDgp0punroVKdlSp3tli1FyMK
IoL2jdcSfLtb/Qr5Z5+j0917svKD+8Q6dbiRQfRCmZnISAeAOUG/OqFQopdiMVmhFtZp8Rql5xew
xzlJVOTF5FxAxAee4wlC6QZ4DGP+OyNwB9ONWviDJJ2dTSb8Tw1psBdFEcHK+LSHOovhO5VjLPrB
QWkDs7uuc0DK0gzeiiMPpNICSnC0g+Oq4wbdoFvgo868AMZPO6eMx9VjzMa60DchclrP0tkIou/J
9iq5alvYzNvfSn1LC4IbC5f18tStBVPdJyucFPesx4sg6xSsD3UdTL/FKG4U5304imocHoVbLnAU
/Bg/T5wTyIdNijlhEqq5rCqYu1bN5VhSjQVwgsuCxCgGinTT/UiNY1xVMaYOUIxlwMwFeMmM+Lii
jpkEGuiT7op1zPPVeUb7WAs+m0WANWEctjxTzkAWM1qzOhXXpbUtkDl/B6Ms7TlwmvL244YgSLhW
jT+PDh0yakXSiifvDQrs8l1JSz35m79G35Uv2aqonThj5dXzfaZsBhha8Z+myixgmMgwyVhx62sq
OcBY8YoRevqP2MszGuQPzGD7lFzl3dcQoLsUv7xave0X1aKimM69csZL9HU4/XOs7bE4GiDmLBvT
VEnAP0EicKaoRdm6wUXG3gHlxmjwJK+TvzWRt3xf+1kFyYRR5vOSqMVrJlTy7rIzL3STLjDBZOi+
d8QfZNVwEwW3KbaIeqxvGsAYOrkhJHCbPAtAbzi+pZXXr/UikeRBuIztRlkwIYGpRPsBADC6sHRy
fgJuo0p+3VOeZR5uRZBK7tCA3rY291rzgp3dma5RxMGwp8FtOzZJh4T4//CD4riYQS6AolzRDNT5
k/nOqkSd1v74SFc8oclT58CdhKmSQ6l4/wT2EGISXbWrNH66OzhfkKgvudkDRppPILfwgZb87XgY
yKcEke0K+gw68mi6835ZF2S2RF/B1wRHIhA4Ick3Mp28pG8TSAqLfh91irY8tjC9YAC34nZBclzD
aKdFDJaVk2Y2qd6DYrbhTc4Q6nyIlUh6+bLmfhMpQM0z+Z4iNnkJiBGGsz0UJySqPxRz+9I/Hnju
WHJdtmfMlBiE9uevZLLaSpOMthcqJB8sI1T9mLzRBu2nPlihlZ+HFXVlhqHA7W180IFTwcSZFR/D
G8YXuKL1RAw+L1RXb3uBtnyMukSi5Ok/PdXg3EFHQyUOs9VRF/rjWxAjgAJESS7FT/j/c9SGBkxq
kavGa9Y+bfi/pW2nxyNkoEO+tM1JNaqq1Bsf0QjMS1b35IQt+Su8dw6IcTPMHpo98fyrYV+TXmgE
B/lp8BD2bxCXq22wNUePlFVLhPSeSMshFFZglSgtEAW2RnC9u9Jcf6ZaOb3elD5xyR1PcR+jlerl
zizd/uteoeAaI4qhs6svKs6NyidICzULkpAebaZv/X/fOFMg2ax9V16ovMRNQBKzIU1TP6U8JLeq
dVczM+bw/mS5ruDXffz0G3icq5K4RJHf4tax9OPTt1WZSI3WHSZL0t3i7QPWeKydQ3X2aS0fX+0O
kDC0vNPIgiWOyoN1zgg32nXdb5K6d95pyCscGfu6Nc2SeTAi8/5fguJiHbf0SWxXVhiDZdEwiHQx
56isjmnuVMK67+VsSpck3lep3vzyA0fdqwsV+za5YsUJ6sWSr285FW7OHLUrEuwmt6MkL0xy8wAF
/ZFTjEl+bX9TLywpQed3Z5vGbpU2sXxO88zLaO9Dyem+yTcdkpQvJeqkSJ6nLJ0iVsIT9tqcXLHg
4DxQyfIIUNAkLpMVaM1LDqKixEB0LIOZKqPbhKD+Pg+AkeBogXFS3pDIYl++GE5OsnZOzwtToKCa
5gwQxcU+1JCEeyUjjTZiUWFDo/XOgAxD/+kP906sdbJg8G95Qu1P0vqaCfnxcF9Nr+yCC9142y9Z
vO7mgL0wG6HZBOdofX4+m+VGNB/gQBH5BUUt+ENOVwWJFvRr4ITzz+uvgMzrqeX3yAx5DOfV/j98
lHAWabxP/TmUBjdEgUidEtifiqo7cD0lYfIZybS31nT6qBif6e0uV26eskup+U2W7oN1tUbBwdEe
r18ASETiUM5s8fYrTDWJpFi6hM+B7XnrNuajJvdAIctHcWmclvtJJi2yOeXQg330A3vz6fr605DZ
SP6JJg5k5f8Licauc95U+NZ71dchyy/LgKkz7GU65Id1cdychX8ht+3a7iJMpcHN3HLNLtQ9NAHA
C3sl56X7ioo0QWQINCmx8vzGaYGP8FX9dYiUS6iwMUOvDzrXEFfCETwgau/X+KWqB6vhncFgEXiC
jtjlAH4Lx/yVu5WtKqFw7Fm7uuG3PfsZOdmmAJxX7sw6W46ltGw1EGNtwzXCklHuBs0Vh3+FV4QE
gFuKtgqhtKwDZJTQqvNRJxRHkoJNAYXrfgBElWQT+u3I9ZwJqrWJ+2eB66R0S3rhJuWsckF+xhpr
cU16lqkGr+ntnQl5FFNReSK6MK8EERvtzvVmbCp2nFML6DfpWbi2AJXz8U+q376G5cSmNnNV4KuY
/tF9rtz5pwlSV0eU6Nzx/5TCczLiOuqV4XuQuIhPfyr4PeYUKzy3iorepMgab9YvTdov5MxEorVV
p/86eqzZdcvBY73zqbNSZDoWv/cRLby2pi1IgAsPCzPWy4Egv08fMG7758TEqXfwcyIP4iUM+u8R
W5DPRpNwitx4jkf//iuP525fKBTUmZd5VG1jAz+kcEMa/j2BazdwnsUWrBNOq9fUYMaU0FsYj595
S8H92rVmSvfPNkk81PHZn49zuKk4MOz2r7MjMdW9EcWMu4VPBayptQNfsqwQgPySSURVq4nRZtN/
ll533YduX23kiigPGSjcCmo4m7uUTKbjHFqiGANiSC1M7Hunl4rv5/tTfUqye49g7Z8+306ehzu2
MSgmojGzhLID9rIvcGEreizb9BAYFV+Wnhji3O9Z7M9wUj3d1a8WC3lkEhO0Seh/Wvrk9a1KITmz
kXUZ1mbqE0gPIpkBZLkeu/ceR72PE4HzGOCARLVpvDzlhRAEg66IV534OJyvjJceQ/Jx1zl34KI/
5zXDOiTn7UTVSyodAOBaiA+Kkfs3U/V+PdveGBEweDYtoyV9Ah/021RiKZlmSyFIO8U/ry0lIZnE
1grZQ4vCd7tE17Y7FaAos0RKEGrVOrvC8okFN6UKQJkvYyVTJ7CtBjgVc+EErKjUHW5RAzf8QdNo
iEV9qz3eCxHHsBxNxUtX/W9XI680HCo4bQz+R+QWIUpxi1PklrcITVcHtpQoZKOrlqUWch35HWIQ
cyJk6+X96Ro6PSjJzWE+8PR1VFJiLDUYu2VqmpHguT/R7wtUg+4tdB/OrITPRvdpk054H6kKDyeL
GrLNTD1rDNHoqk+Oval3OCvrdjsa+Hqj+L8zUhTz9jR9s0g38k6CFUp/H3tvTA+UQH80sWc48GMo
CfXYxqcoaZlpUyYokEOX/ZzOp1nQfHP1XmdQ/ztFfsId947cEWHSur/wD7i2FASTIzQBlmsp2i7J
Tgh9UxWQFw8hpmkRC75waRdIrKZB65liSZScewgi4b1F4YaUqc2qW9wVTt0FXnD4r/DK9FKtea32
1CAKrpg/B1ZrlGVwpHrEAqoImFwG7k2fIAHeFx7TTz6rRXiReCz6PibYk5zCZBlsH+2mFKDH06hT
v2mNGaq6i90UUf9gBYVpSK9bLyflxuJV+IUrhGeadiwfNKnLWtxuVKCBr7C37pabilkYGzczpV1Z
gvsBT7HoleT8IC3fhwo2MvYkJX1DovHRExhHolBDBA7YLrU1By9KJtkvvIM1fx2OrhspEnwm89DI
uIQghSC7rPPEFHN/a9qVJp79Lspz9aGptz1kGSK9oMCG3LHRTTNK2h+uzmuJPQvdEQ29g0U6BFjG
yxBggJgoqt6ZwMay3PCfNCJfizUaeLdebybx43iYK9QZxNY/sbE80dvtrcGFc/HUs0d4nyRW8of5
6dtKKfNWMihaEoCYPffB4GdoSxvSUF3HHEUokWhGkwMDQw1mJQaPWWLpIU3W083nFuyGYza9dKUl
I2pMahNfOebdpCEhCnbSBrfOtyrey2uomATK/Rt3iA5ozGZcFh0my3RlboMqHW9pIAKVK8g91m69
F/fnRXQVWAG9umLwckT3/iOoP3dofSn37DtWFrpYny1jyc73lmMHspjT5t9bO6OabV5XmHce5FSR
ot0JjTSnsWWrSLuLlgiF/TS5Ft2BtZp1BuWFunVhaceQQ05H7awudehHwJZF2Fzm64G2Q6oQj2c9
eKzGOO8vdGacLiv6zEvLcM9IpK2P6Mf37fFQbr6Wg/GsR86x31AszfIANLQWUqbogphg9vhmuqc9
RHsBExHlFV72ePQwoR+hg/hODAO7GWMNGuUNnlftIPVTb2uBkH/gIoeJ1nSkpYLE3mqgKNKSl7yD
t2S3Rxh1kpxJSpWb5QRgoNEsTRaZr8JEYBT8YlCmX8QwwmRlDhjWZNZGFqV1fMJDWl7wodwx+zsV
zigCuImdbJQw95svS+rPEpbnEgW0UiWPPIWh9GVCFcoCDP6X/SprE8ERD5N53LAd3FfO1UM7lWlu
ZaEdA1KqTTdM3iAjP+zxgqSR5I+gIR/Gd7hJrtOzjn0rnQlyAGD8nn6St0+wBlGK7Tc61Ec4Hr5y
lWiah+aNAtSLlatvJUGtSuoQGlUdlKBzTenGL9V4X9TvQOsSrF9zpApYhJlyYAsJ1SyXsTC2rQhB
nFa09m3NP9eX7bMxCDSikLMNkOTtObNq4mDlF4seoAJ/7nmkw/y9IOcZTDg2MKwDZyr6EVW4yYuZ
MPevmZ6ONOIr3DcnfsGfktlf9e2qP44ytKUGI3nVNMQD12i/wGo8KwDtdQ2LWp8AAN1meqaH34sw
3RW4xsWiyo8AMcJQgXsBC3Mpp6lGHd+AGaEnZVNP+wo2Fx96KhHp6ZvODOlFaz2m++02LTUHzK38
eUo8IalBVNQvW/GoYgmlgDnSDT8796yfv/C1wBSeOttkx/yKl3+bn0rYA37jDS5nydiw1jWlzndC
qJj4/pAqotoEzdZzQrChQbdesWLe2c1S4Uw5AbouytF8TqkJeRhhtuQnOE41TVaBtwD3+N2Tvzmk
jzduT/WYNXqyPFGhvNtP2vUAJtlpiSHannRY7ZohOS/jwJNF+8mXc4SFkjxVpymnVIW6cvQtakfu
84dRmNrm2L8W7UtL2Rf9f0PL+TtmyTg3eHiakXhsfT3E7rIc2Ruwe66K45ni57vsS/PxPzViJ0Mk
spiJ/5C0OfyZTf+tUj7YqAfqQQgjZJpr1YN2u61+aJXwLEuBvmeHDDHBqKkNVAU1w31/yEIic9zB
pEM1OmjrD9zVP0zkMUbr6IDctCVzZikGFlyqjOwXyID/hfW9rtF4zzbevVeBrp44qceXvf7Rct3V
z6yUeqN5f62+Bs/LFhwoE2gdG+Wnv2ZcUheOXwpQNKkwH8c0m1z6D70It9KUhcvjjAhalBKPr+DS
4f37LRYzYfZBPUr4TcvKNYOYTLNM26CPj+dg50AU0Du/Ki+7p0/zi2kMxhp0mC9GjNMdZdBdx4A7
3Ld0pf7qg3/KNSSadfRCfkAg19eqSOn/HSxg43qr0RJVDNQoYm6wEjJjooSuCpcPMS/eeHZyx/wl
jGuJMgAxLUWog80Kn7FiQSQvqlAuS4hBF/lI5NqHi+XJlYZoFSuVYcg8qigooyuX4R5LYvwbsJXB
vPN1/vnhDnLNQ2BtU9omUWomZFl7ynbIixgfXhZ7OY13ykv//ReQTGVK0Wp7t99ly/hR9RNqQp+E
7GOYBGMgIv/zof6huQowqzUzOgDZTXFqRp8IzeH+IKNtICZm
`protect end_protected
