`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
SXgP07X0rvniKcSpFpCBqxVFZI/wJ0LAQzu8a8iVHZ/WzjhXG3zRKGoShC+EvSeLoQOA4r0KT6OK
tRKhk9iaAUf38K9Z1Cco35KSxYcAZ7Xaq+vB5rVDCvgnDGqM+TtW81V+Ta7JYLVygMmtvIxFSulY
fvF7C0nRQ4It2dKijGNaztLXsxpDFa2VEIYW+Y4+swyUngz/IebGwwvqZafYNLnatSl8JGJxlXoB
m/REY+ewnVbqF9DzlyS1j6LDJBDrOEfgF3mAShJpVIt4jIrE0AV7dzNF0YW6vsmBQGxvDZ9uUFvY
8LNSxmdkPUzkuAUpPnjEFc0R9yrAuKpRIH5phQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="tg9EKhiVh+k6KcOVwrkJybobr6qH9ACed2IulwtQcbc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7568)
`protect data_block
RO/1PuAAsDhLdXaaMFhvd7sTvsgJoRVAYNmPBs/beDoIH5HcWnAghOU5Us9gaAm2fw9Af/lNQXhq
I5sWvEK66Eh1uI/JNj7MIhbYelFH2eQF1yLdXnY5SBMuN8R6zPsU9xKLquuaIpHYsrab65HKPEgV
6WL7woqcXOqlxAO/fuKcF0PrOcR1UNNH5h0A1aOORmqkBOIePnkdcS5blTp/YdxmvJ88pz83YRW5
wKqGG+gXVeDPKsHxbe9TlAa31zGUZrMYmRA1clwIdBmokMafCAonLbLehDsZj5SN4xRkwrjsrjLf
JCgNgIF2tYwnpiLOme+tDe7dJp9arxl7DAMmSJTtt/CzxMsfPeglZu96R1Tsvz5nAIgM0vQ87htc
qLza+N1RDwrEHYAipC5ODRbPBEEWRx5UbXZnbAmGe7vWNM9PTq2jjqX32ElIvdi9fDXGPFhhaO9b
ytwSCe1T4p+RhWzQcziPHeVD8Fuu7zzxymDfMil2PXgg0vzkRewTZGqshGokPKxrf8YG+XKtXVmm
eG0BSxJJ7acaGTZeI7Ii3sO99x9JOuOISYY1Dkc1dtQjS+I+yMM0saL6swFNGdIf4DKffiyAGOiN
KqhHmiIseUyg9lNaKpIValZDe/lfNAaQIY9rd3X0mcO0Ch2VRTHql4wbLc+58EEQrfrnXO77HwZy
YHFaNhTMEEFJZ//D8dDmguoINEIZaI/mklRgf+CWs9EdlC2PmlNnVQgDyH/+pUQKIzLuKwdeoqcC
AZsSSMO+2MN+fno2pwmIbg32HiA8jLLI59UKiefhN9ugG8bihoOJ25sRsGsYfMZgLIWBL0qUycXd
Va4/OFuvJFK/3fNLbOkk+TorLvS1X+pTFYUurjsgcjH+6gLS6TAOzGNCQTw48+gqqoHsqaXjBaEt
p61iDFWoyEH4Iu10TZKmrErZFz5cwJi+zx/RTPBg986uDQo7SCgCF8GSZg2N2uOtWhXMtJfzOJLW
ISWKBhTm8hF2XLRMhpDVqFeeC8YI1gT98eXS35ZwsRCM5pbKRq4hZeBVOoljizI6zrhiRNORjpXj
4D9Mz/NX5Qq7egpEfgO2cFlfEU94bAs2Dep9ln5LHGulAONeuqKGugARMjrN27H+xWJ2VURzjp9L
U+pyMgWtomKUyfAUWOfnij+pqPt8/HquwFs3d1E3q/pzyXbdt1gD8I6BiWwjEp5a/Z3V1RkGbWzP
B7+PV/zCKZ9BnraLsCfbssjx0GPvIvA+I7UC1a5vZwj+P0WHmC97tXuipWN7xb+h7wyqcT5poEpX
CNprrzFHzY13AMl+j1Mz7H1sT1ed3UW8urqtl0fwNdkaDHYLdnwPqDf6ll/4i2KgVmVIJvaESwhF
OV5/wY7MF5xVaJ6+8pSssQjlJT6h4n6A8XQSa7Yyru3PX+3VA+9ESlwU26zrOTfCBAFYx8v/vp2T
AP1cp+jPSDO4lwaTJ+qkn1T468XlFQBlZ2uR6HiSDhpIeaM6mNcvBv2jWaFwtLhsfcPWkb8UmITF
S09kX15wUb284Zg3euEENwr/1TXrMvp7JN8No+yaY1A5+bnO93R/Kd33JpuZrx7V1SUC4xpo8Hs3
C7wmrbKcdcnuRLwPj8jyDFKksxpHj43BxjJxs1ExFW8ubsRuHPeyDyJ2oVJRW3YnpJucKlMD10E9
zuV0t8sgiMWPLlhf7BiWf1ZM9VBhbX+umLHgolgXoPcKRFW6oW/T1dYrjUoHUF36qzAnX/tc9kB/
Ov6ePvi32uhFz45xcBjLsypukOskaO704BKQRpaB7DFymJFdxSfsyXwAzFi74U88w1d6hhtLIim/
zEBL8PKz4hFX/uQW4TYOlw7VWGXaH8a52xxHu2Wr5dmz0r373R+BN5SK2AdQnKCg36gtA066kyjs
540ZPOe7w/B7353ClaiupP7J6BkE3+K0LZJtV66aWM5F8xrrThSKTkX6hZgMIz1I43LrieDjX8/y
IVE2s/hidgL3X6zCzhi2KGp7f/O6FVrol4JGwkNbf+/pBQkr7ii39bkWPhAj0YZjfitIepuySZEK
kLbKVb3Phi5j0ZZfVLOe4A5NUs4FxQsuEzVqkdjAtqTggbs09HgMMtQISYyKfsqTOWCQxHfhOxZt
lvghhgMFxd+RAOL4kWpEqD20usu+4FF8wkWoCgcqMBbt8V9rVsbvJULZzTAHafBpyNkj2gHdN2hK
/xVaN1N2V2HMkaca5oM1Mf6gyeOno5KaQjnQ0vlnQASofD9MoWjqB5ZvyCgTXl2FS4hSK61G8p+m
aVwfmaOsUa2p19qMDPQgCFWKwzjH4VDuE8pZlx8Nn0s+qCQjB+0hoC8qdogfCv6T1wlIgpTtmj0I
LqYo+8Zsd5kQQefJ9uWjl1YKXDsu6NE17bH5JFSpPYpBq8G7wlGSqsALCL8TwDBNLGzV0PyDsHME
jjB2fNpCU6M7byxjBWM4v75G382diXynLbkYL5WuumsODiQ9/m0lRl8sw5PoYO3bWgG3YQ7NDmy3
QURp+n658DRQ6r1KhfxssdEBCA8eR9yI54g68aPGcJo8e3hN7TKZmGQPYnFzjVS8dM6XmI7t0Y7M
43kdMNKt3W9+p0topKKGVkaQCnaa7bTVHHu2jN3tGGG6BeFAbXil55cKrlVHVKISD2Mvob/ytsw1
2KSWZFBCSmj87ugkgsB5LuOamAB+BGy5dbKE2isNys2qj8lVUHPCaAZeSxvZJ2X8pbUIw7WDyjfo
GYSzQISqu/7mBGMSUE18AOa/xDA0yrZIWoHIiKM3RRdjSPKy3mglMq3QDekpMNv305AOdKo1ncsC
4uLCE/Uq3LTtbzZY/hhFVkRnTkdtR6jlMN+tjZ2lPBtkJPQdI0F+wqiVTsCSsMjkeTu/zAM+1bgH
QG43Y/0p60lP+OWXFQwaGePT5dOtUdi09OfLfueOVaCLYrq7P5sMBjr7AHqa/bg4OnQfSDQPrEwO
2lqHNvixZvC0LVUU9G/hMZ9FDkzF1U5G81mf2/UsSmMZxPlkR7riCCUgTfNWI8y3XY0eNuQB5Fpq
ZMq+Mrk4MflDHg4fMhmOTZ6w44nKN9SEvy2+dZoiO6QXYkQSBkkr9//5jz06mb7tebi2GMVyFk7s
CqimPxmxwHE3WSh9bwjjCG49TxrIPzAe70CMuP8CLx7xv1AcwoU8ovS29P+9Na3AdNRpkm4Sl3YI
nuM8dHN/sBd+sN/RML9CMiLlmgITbtNCESLRw1wG4MbbVA+nhYF8IgFC0Y2oONnbVKB+L4cSaBWn
aTEkyAU7w7hZfVoDWjvkoMEaKh18cUb8fJBHbgI20e4g2AsGKtbQDXFbi7QiIYCabstRcysUpuWZ
KHZBPcEEqigJrzlg+ZKfzaHivI7OG5+J7KTHT9xURfMyUk2X75xMhCDxjdhJjA1sIr04koSe+j26
gI8gL5ZQVG+LcjC56rUIF1EeLIRVP0Q8qttj6IxG+NOh6QCQ1A5YsIyPq/H87rszfEavA7l784Y0
n+bTMwiH/YObvxEAprmQZy9NjnNaT7fwKnwExjdRjs43x3CNJdaSFFk9RSJ/afwH+9l85a2/6jV9
S/zl9wdkgcujStlLbko1FIQIeJ4vnCXJqVxLherYLUY60xux8gptmhUNx79JU1y5wbX241u/AXF8
2hHOKYa0LppBagHx12RsRvsb4iFSBC9F9WWNP6f2yj2fjVXU3XGNtbyswcB4zpRZ3O/n//S0InC0
blHZoaMeCAUnEvBOczdARG1WeiX5k+AMifcVZVAH41TG+yH00nlhU+I6t781G53S/317ra45BgPi
9Kc0u/KWAgSaUh+6zwGn9ZPN2IZpSOBqAVBgYsKWUsUcckCatDUEzbC2VHDN0ag+XHpx2TKnLHDs
B0r4pEweYv2i+qn5CKhkKLnIQXvNFkM6w0b3W7YaHPx5ozHikJfObBCM03yOwb55aIxfg/xkWKop
SAmyfa+Gs3o1YkHBxFHefe91uxLnF8Y/eAxDgLtfxn1Aap1DKbQFhrmlQjb7iL1K1+pbu9dl03Yo
Rx/u2GfvPQgkjgo5Dkw9BGkhrMBOgoBS5Oqk94UCatI5qEpsMT2FlrhQSW1e/2GM7s2P2X0dVmQP
cqYAtFCD6Bc9hCr06paBfQ4XfUBeUVseHE826PSKD3sj7jedE87P/K+ZL3fiIMME9sitq2BwDI2N
/AczmWKy5q4s40dqHqU6wTdn7crWypODkOb/rMTInF1uU5Z9qeC9z4PH6RKAZQ31EPdF6ocp7fjF
2PewsSL8wpluVYlG7Dog6TzzgSqE7pr0+j/QPAC4TISknoHDaRXJSB7GDEq4lJJPZoEgfU1ouQgd
4UFa4f2fDjsB+nslLFwJ5EYdDCoJ/yZ3mFnZgJlGfZJ9HAYPd4ADlrHxsNxv9DYmjcA6JUgZqoBh
BpndoqqGOvYB/dXHlaUCDxZpCjC3wlOJ3NAaDn5Yk5DBL/9Jxg3CXNT9DAmJBhgvqn4G3rrQvmiU
IEzoYm/eKchTzf6ShklCPSQBWahIQZhAJu5DdAKfa3zbNLRZEJoMy6rYtxstr6OXeL8glyNzOqvT
GcDAbaleewsvCQpIun7y4ze1xDkjwEOdaBudcA0N2UnPsQpYW/FfUB4RdRSoeenyG/fgLnE0kd3l
D8rSV37yHATKvLxUnxPVk64FjJOZBj/911feRr9kE77rYgsZdbMOLNyfnmIox/5UkKv5ogo8FQqW
yPuzMNlhsP+yV4NwZeIGUj7y7Nu8LoasvaDQcN1GfSNfaPYYe/PbON+K5ZJpFqT0bbzOYmRzLl7q
vx9Hum7E6+DstWk9FVWGfhOpjK4/DVaQDekZr6+ZCyUewExauyD45eLIun35v5T0rXhvbcxcP1Wi
cCieCmVyDs7dCXTbYP1XiaqRJwBBM44gCRWbMayPSfvS+oXjf7Sc9chSFBpQugkuaXbcGMiz/NvF
uSlkGqfn2rDSECx3IWa9QY3AsSYQCNMzuwbfTdsvNg2uWdLQTiVBDcHuI1me/Kc1noyBHpxwHor/
QaCTiLdMPAXJ8/mEf8PbzrABMcNkt5LEgST0ohfGr7dP7dELpc0EnvuNcQ51WOxycqNMPp9N3t5P
RobIJdcp2OK24OkdY4/s9tlCIw2FONG17zsTgVdfLf7MKet0JxtNSCfS4Gob2tt3tgzM4Tu/j5sP
qiUPNu+/jUgygPpQel4OYQywT4zV5hPELS5YEQl+cnscslG3sU6w4W/XD72Gohyz9LWhgBQVkZ1P
frjDeXx4wfvGC+YSSOxYys3qLuhOpXgs2uzpnFF+t1uBfAv0pp/Iq8Zz4EmWHP14pPRxKLTWzUoQ
adzvgwVBFPYyc90J75uIJ4eQk78PtytuRLxWwT0eQ+tdahxeThSosh+zwxrSQbVFp55mkm4ACIxI
O5K0EmxAei7m7n+Vc3u31+/YxCaxsSBXgN+cHBmWKxLorPNCDUvrvzSCC+ZI65I2HKNCJbatBlqP
HVqwzJOaUqy4Ws1tRbF0Okj6ddt/PdqgdWaM5wkobIpXqv3YtD63EIE7w5xcmvo76REa/yT6JHkl
eB1Nwo7BEjwI2i1atXszQvM782+wHPELHWvOXBzVlK4qpWAF5nF3hi2lX2a1aHjDZ7hZFrnBTbdz
wyupZST2P0OGCRfu8df3Iwqe+houQi6rByLM3SLZaO5NN1d8p0Jy0dA2qn1Mo8+S+GW/zS+8390o
+0F4OGcg28FkvscQUueX1/xke50X4OKn31YQZQvh58wbrhDhY+ubufARWDnYFeGFrqB8WKNks4k2
aJiyYIiJz/lz9n/91FGo04QnsUw0HNTQufzOd24KXgSk44khonrhzY2s51SHu7WINOjMj3dziyc/
8LEUPLFoXY8ecdtr5anB6Yd2yJq0mH4Yj8dmMbaTGfP42KU9vm2FVBb8e9khZy96N9ObJ0Y24oYS
ME/BAdpnoX9rEEAshrj8J2/sxnGVfft9GjV2FFKiOHwDeBX7SIIUUqctSkMu/u2cCIPrm8IdS/Pl
ChzoTgOyASwfW+6OKXzsFTPkx08YnR7yUOld+3UjSJIl4RhUkaMdKLyTuO+AH0bi/cnEaHccfu2v
UH3a8+p5sl27THbLdWm2/7iqdxAfnaQgk5Bsqk6GZFrEQipxJ2fMIYl4hDX6hgDY8sXO0py/mEBW
jGBxkNfQfMtN+UvRjWnRji9tcyStjHpLXKovvKqPDYaGpc0CxNHPfXJk8vVZsPiO3iaGz1nJtqaD
7PahUs2SftU8DtxlCV1zXsb8c2U1cbC8dtCXWRXhhEVJ8DsU0Yk6rtZsXsm0tG7eexasNNk3SBFN
hFm0ZwVIY/l2w0aeacqVaDkQ/SbTtvYJKGpXlUoltKphRPOd7Z7szv3uU95B3MfVAZn2wG0UGPFm
kdYKXFuThC/OeseddI6I74LUnTrBvlFuJ41amRktXksuGfF/g+ZpdV6bk38xWQSpxn3zevN3QCMa
XhSjUaUnk5qTwYoEO4SryC1jl7wCX8iAoG4ipV+7xD7vytOGc/AdOZGuJjqVWKhKoscD1yj22GBb
ubkYyOi4Wpo5k21Yn16KXxhG2Uh3AdCA1p7O5v0QKtGdbITtrCPRvri/zvmlNSeca09sc6cPhi1j
7QxW8hGbooK2GUuAViQHG7wSmh3C8mrDTUDHZkRVmI5F/Dmeg8jevBf+GbwyyqUBPCJaKIFu4mZy
12Rp+CYRCs0bXdH8CVhopjqXDBkbSp+B+7FnriGru3/ZMxNdChvW82OA20tnw3dNZ/iuOptoxVg/
y2zMyvZzxlAFz/N0+yag6DU2hOzxrXSx4FXEgfIT73cMdIby2dm555FHy6vJV3dDEB93U1GGro7S
VOEmbM3XynEC1Y2+uXQ+asJhQlQoWGS3HoZ/pol6NXYaTjyHWSNS4o1zaLAPaUSzLmbqCDv46LRk
BuWnyUM4yloQoAjvPvz6VthTuit+4nn8GkO+KIbh9cWg+6JknFH93vQ0Axr9C+oHdI0wHzOTflF6
JWHUIiNg6CZhgPOL1HOhIFDPJS9xQ/w7YyggXwU/d01r6SAZfGhUa1vrYUwTuQGyHDPyFAQVRs9U
H2xeBp7jD+ONTMH8542Shyspg7VU15ANM9OS3J1wdHwkM8vIlTIgFKJLXUW9r6ySLEfdKd/It+ex
sQy9avwo20QkJZO4mo2tlbxgnO1jq38LPRGOHez15LyrbKyMqs3+srf7Skv9obWt5w9zqCwy6aLg
34D5TVZDkj9jrhRIGfW5RCPxGgdl97dbqtRwHy5CcH5ZWeyWJL+b+Owg2zNHC8WJVpG6tAYeQW33
4ILquAQopgO5f90/ExX8G1bKnfGBAXWZZgX1bASgXRJzYCYJK9g9hDDCv8TdBr8i3vOzAyaRE+B9
nmKqho35fkaRVpeHgu/OaAuQ3i1HFwinwccS3f2YyB9MTt1hER+PY1LFqbbP/eXonjzK7Vq3Sz7V
ANKsbjL6INnZE5sIEt451F8rK+G+fkyHq7zCzLU0a5C9ZfgaiEWmJekfbKhc0T+Lv23FDFnWg2IV
FNconkTbIkLXkTD9sy7gCKbhYKQT5ut6CczbH9hUpuKIq+Bc6y/v/37TKof7sqEnxUMynCgRDNAD
h0YmM1ALHhMjSCaptc8IDUA5fyePSjFAyRogxg7BHDagulQPTWsDiW1Z1VneGtnHKFvolwh8xblb
HBl0pnm0eEpLmuYrc+JMAzv46bSfMOc7NO5usH7idZdTg4K4avRWuyIc0zDcVKhAVCulM8nJpRZK
3CS9je6V9XdTS1cBASz3kkXqLYabYTS1tXTyI+CKCQDLW18AMoM6slIM0BWp/KA/FDdE0deYqrqD
YXpPm7OfKpWp8lOEJJ33ruW2gRqKLYUeBEP+A9oXbA6mPh9TyXrDT2NNOSpjBV2qhM6DTpE/2LXY
Fm80L7XO/Bs/X6Gq1bJboRxfD8DpJXLgHq6+JlqvwK8XUT91RAw3pQQsuZ1Ph5Khrjw4Y1etZmGE
oWhxqFqPHHUaSghDSP/v2Hs+lgQPnh9EVXmsRyHdwlbXhT1JmpFVvkCRTGo5UBdZRO9HA6uQhRJV
PSlDAK6PWPlRCUe6rQP5DLsDzPJHhGHL+U22VCER0e/syTPGrUrXpWNM7jbG7vB1lkX7QJ9Av4ba
YL93uU0EHqSyMoGA3d282ezfrlrNz9SvdazJosksrwwVk59ZVC2cw/EZkO6jBVoFf0b5uHHhP531
c+GnLd+GeUi3+2TilEsdNqojH2Ra4aSPWmJxPNClurJ8hmzxBt/zPUqiLsIlu0E/seGE8AuhosIF
JcOBsM7iOn6WrZ+AJEkzst+JoKcugdXjMw80o0wZZWqdPEk8bBoMpYMTaIbCWgFZy77BtMmWAn3b
dk1UG+QjjWT8NFg/PYs6TYs6NQaID1lQrSA1nJoAvfj+YeD0ARw9KUK7d8kZFCNwPm8ZLvWFHnMk
5dE/2pLgZsJ/S5vGOCpI0Ub1G85BCv0dnOl61qh3YlnNgP/P2nWBj+AE5FvlRoRSuDFFTRlYQTtG
pk47Js4SDaC7IIqSJdkrB5XmuN+gzgGYjcH6KzOqFQEp3FToQT9IHn6zh16PwZsA5jyIARB72ISC
ot8IwSlSZBnlowAjZKepdrH5WhSlAH+DxZpfSW/XTlwp7+1H0GOakMNhFiX0OZNq7KmTSlE2qx7T
e7/+Fum3G+I8vveVsr18eFCtysdNvv/WkKw5a/DeNxNrx5B1U527htZwICEQjQz9hB4rDhhGROkV
om38inn0S8R0VHAd/Wv0Cw2fUO2hCpBZAw1lTVfnQEB4tuYLeXlYPGLkpaIFCyhYq0oEF7uup/Bk
P08rw57rutwEfYyVbYY0XfMtyM3EcEEVjTg+cei00vUJFKqzcFIkQOHEQ/PtZpb7BOm88oHDUzdQ
znfGG5MxYRBJIwS2qqa0sKOGA8r9kXpv1qQwAeGCwBlCob9zLLga6dFKqWVqn5JWXbnibWyUOsTw
P7q/XYeNLc5LFh5bDUzpthpQ7jGfErh51NkydVyiE6bbNVoBiLl/Ru37W3BT/0w3a80tHG8rxCDs
JOWtkk094KveJjL6FecwNUWrBwdqhyvbElj3x4N0q4LxgjqbMV7W/mLaWKtclBoU20iDi0xwV6+X
CC2+EFPeG0ntC9I7RnCx+4yuCck0ZbMs3gkSSMZLUGnD8NpVzhdPo/j9viGdq2v6wdqeoh77GWFr
WeDEd6UdAdAH8UWfznKlDKjGnYPrVQx02LIJdQueUA2girbkSk9PGs4QGBqTDsu9f62iR3htYC/b
s0Bk+8lHo07vUKzlcteFj286xpfqmX+xuOqi1bU0SfosHWZiv/IczOtyX9hVn0cULIBcrNxyFA7i
v6QrU4e3muDw20pbUqdzE6GVFNL080A3BIO6eS/Px1dqp/78kv6ntMRVlUtuOLgxPDEOvpZ83S0F
Rs0pF0qO5OfZ630JaekJLRKmmrOjkQ3oJ/y0KEUBdpEIAfLnEWbB77TnacQhINPNxCbHF9wwvuBF
aFr/8eui+OP1rtztOJKIs2CIjdtxl1eq4/lzIZqV9a8UEHQVIrtWSBgHV1yMhB56R1VRJNRU/z76
UGwYvuEV6gzyWoll9t9Td1c4oy755WGQjvO7cjI+3Dvo8nykNd8+9kEQP71Wl7ZH+8RaB2K6khzx
ddzyFTNgscGoK49r1huwHxWakTIwMDx6ybMrnkmlAvMtZRoDd3zlXTTuGdF9tDPxS3iDH5oXIDYy
HCvCNzHC7qViVpBp5tlYFEoJxpE/VBgy35/YtLfVyTUDSMHfrXhmwis0Ec/sk/dbCNcEAsBrGMXQ
fDa9t02HzLrf7GFB1fSkib5Qjtik2oohqJ4l0jmN0KmkV13+0ohDr9aamLWImMiY+vGRJDZFbWXV
Lo0MfK3p7dfJOTUODJ3jjikZK0EMb1mV7W911bBYbWelBUQBmmpApKw44yFrjfaA6jldEZYpn7Gp
CDTbWhFaGsiknHs7m1FE6BgWlV23H6caGyKr2CjvSfEOJ1dFmJNlBECWldfYpbBB44Eooo7o64pD
UGzVU6I1aDytRnHxEl/mSqG6/fEGMTG87RZ2xP8OGd5G+SkUqPLIv/TW5y8=
`protect end_protected
