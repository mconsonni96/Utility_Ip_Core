`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
F9dQCBxRQWuDAkeI9mYrpbHBWCAjr9UEeaNz6mxuo6Z61mExXhu77u13mF2k/+OTLPDmMMqQzdpt
N/Gyd25ND4VPFOJHL7aKnVzZXusQBkV7HG0dgep0b9DampX46rtuksWd6RSNw5d62drVdRlGlJC2
CYHVeK601XyxCoDr4FJ8j4fhBtv5JRNMNHAOIHTQX0W7bN2EoqNRLvPByd8Wfvg8o2f2mYdg6yil
J1VHzwxRLyP2HEJcjJSzExMihsns4trZvIPUE8RGL8IOOKyg7J56hErbKx1J2e0onKoNpXikyyTz
XcvZyJb9Yzb+yK4Ag20zcppAXdSemFXEMCu31Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="RbAUxQ8+MFXxZbiMeJW247cBBGfoY2je2tYp6J2m38c="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19408)
`protect data_block
FraeFpCC+NduYIUXk1WpHNeelXWNgRfVUOryMPqudQgJG76Htuup38eV8kRqjKXkmc9kyXK86eOU
cUW78g1155AuqjIB6Ycbcf3m2S7UeTrSGWi7VTMEOpl6qMaMxQw7WMPy5oiZLu43MVnX1rvFCgmn
nG9QVx+nzx587wSDse29M31PH8diVLfJc+KUTQNXGm+ajxL5xR076v+Q5O3zoN8guOGqQ30BzHYv
aqundOiFIZwxr/G/V+C9CpePwlD5t4H4nnWn3qMtGNKTL3d1KMvsJq4i++tEl3Wb93cHAL0/twbQ
O/lOicoWUPvpDxDupuoN1SXy6Hz/ShQnyE6jj8plgCvlhN4XmI9i7cNibZAbCqkLtebyjluFvJgX
YwDxkNJiXKkB2QerOqYjiSOotNztzkkYPnU+vL/KtKqLmb5KWAysnc5ZgxLZWRcol6RHoq15vF3I
3FUc7kxiApI7OwFufbOroPM/69KutReH/55gv/owxNPlNa7c3ENY3pM3sFqZdPDq5BMxBLd4+QLl
HQMJRAsX2oIOU1s9NNuVCwJb1f1UNsQO2BFxJvQlB+nnZEeEQIspme7fKUR6Z06TCfiikALH/hmM
jOePxfzpwLEWfq8+0XwjRM8rlMTP+GgetqWmo51WT9qOy+JgCVo773SObpEjgwzGtIHlwyri0MzA
KzL5SJGrZcFD6054AmGDiLGuhg5aHTJeMa63ooFtTAt3ZiBsaxA8yZaKv+WhXX3MnxbL7pxFkLCY
Svn3KBOgtYvhgJqPpdn1iElb+dWBVBKQheWbTJ8QmkhvaJ6M56NSXFOwYVKNBl3pSbFGOxyiLuS3
4Al7Bp5v69CCZ/q8weDZDslpA4r1IRvMa4ri21HWVgb9BevnJ/1CLufURnL9lmdtrAZwxxxMfKIr
9rZp6R86ACIjRyskuAOp9R1Yyw8fa6dXCGv6f4sTHzpyhqJvVAzwbdp/MXU2Y6ygGe9a+shUc+5U
Fr6jl9V55jvClCq70xopzetqOVgcV+lCiJkVKOCXFVtK5kNIStNW2XFDaVfcoZT0Nyc4qg0zhsIX
jgld3c0J+t3X6C1z8ZDCnbanYtezFhxuyYn4QpchDZNEBQKYU9ouHntM5uHVGpZXCnJx9POzl7Yb
/XgtESlPeKsvLyO1ebLge4gcCXVxRsz0kOHfxmK7/D554CP/QVy9yCrSXN2XpZfFiVteuQGYbml9
gsIAeftkOp+Iyv3G1RZeEXtu3hbLEGgo0Pd2dsyyq+UO38P/GQ+aLoHWTX1iog9jCtiA4lSD8i/Q
+e2w+eptKcYqDpeHn2w5fZDABXvVH0S7d6di/LXDD7gadHe202GSuMIK5cyyVxperTHZK38yEPKJ
Fda5oTMtjc4yjYydf9ZOustuLlVc+VKyTEuWqQIXYLy/Cs5tIrpkkpX1CMA5wZNn4eqzVBBN01UQ
Ck85em/h+dJed4uH8+UsoDLtREGIddGO6OWrFJoeN6+eqjFSsKVwhUMLkV9K3qpBU2DGY9S6vkdk
fRrbvG02HhmXJ183cy2RvjgF4luxRhcvi3+et75xHRPKtbC/hijsOZ6KNHwNrs/U+jgqmObFzGK4
hHEZ+bGYvQepRn1+Cz8fUGk97576QSGbnybKF61JmTIdsGtRQgTWfOXDejkn8G6pLQ+v45urcDdZ
fdNPMIhmS9CHjCJqLbWKkbSb6mKaWu2sq/SYiGNIQuY8VpskWnnMBNdiTydjMSk7KjBepBZ2uyLc
xuWdZF3VP+Oo68tgFiDb96B+P1gr29IYlZRE4raxFquZmwNKtc8RawbOdGth2tp0wWgZdr/Bq0jl
4tBWo+9clGp2Afw/FwM8bP6AeETtLj11BsxO70eJEymTxw20+N8o3q6LA4ZOcrxs0k6PBYo+qWE4
5Wg9c4Tuosj+/M1W3XoE0M9VejUZ0upp2hOFZEKs3SDplpe/YRBVr1ZPEd/n5JNCjJ7RuQTj1xk9
gJB1TGI+eJfYzNSrAMVsi1b81tzC6Q54kMpqtfjqEjK/kqGJdGZxUMjvtisM9pK8qrBk4V/4p3So
R7UkSCt842HHWMgTjoJiHbRPOTr+qEOUpd3gOL9ukgPqUoW+C4NsveBMhvnY8XKH9aMt1vLYue3x
bXWKYd9EFfhUDboI79SvghROeNpiiX2bjJfHYySJ5Rf9bYklOv+hd+j7nqMfqX/V/0coxLDjAnZP
6WFkPgbQNNFaGwLrI5ZIzewQvS43Zf/Df/dbXUtqXk7dgOoaRvECeCvwpmk6zjE3YKaY41WKiTZG
fIKVvTKoHhEznPX1KmEndM5DKfsBuIYBF+LmLQ6DQA2x054M0Wn5tuJJAhYxpV6DOoPH+anSAy2B
m43jB9ff/rvP1OBxUD5c2nqWFtes06bNleu2waWlr6fPUpJHpLlMesBH7hV4Y8ErpzPkr2PCMaF3
okzYb90nE0JAIi3qwvu5s9h02Ve7cXD0M1qE80qEOCSthZ98UzkoldgExi1gqBnitfIjzmeq1X1L
gpv0gISzgEA/AgiMWt63eEXHejoOWE4bP2sbBhQWEp8/nH4diQoIR3+xyNOqIh7ipW9kYBJxKRvA
j2zWdhxfpp85N1tZ7ZyHCrkTGrOm/dzkD3HI1djhSi8P+V6kSPSq9YhDjfuXAB5NQVdeqUuQQzGv
SQfHNzDETzze3IOuAW0Ibn/PKiyhM64D83sxvi7n4dGLQ+aeF70UADZ7DQwtFqQgIKaIU85noynS
uaw5iT5eewXkjTI+KPZFWlbr+4gbnfnAJr08VcJC94ROTvsULYR0xBplDRfFaNlyn1y4kFkw60Tb
z6v+ApfMmdYt++ORhyyyiQMEtOaKeqcMd5dhO7xZP9aF1GjFMWqESdi2hAhBV9Gw6L32fAdGVW0F
Wuu2egCADzDjNKwVoYrBjdD4xQ7lTJDefaBr3h+NyhhgOXb/Sk0zlpmFOdLohJiAR1eGJOd2Kb8P
hWI42PPRFajvKrJsf8I6DQnt/zO69tG4AjJS6/zHRwyDrXhs874ShHaA7PU2/YBQUQ3T5+0JAQPS
RiLXnNKj0bk0JxhSEpFZryos1aZOjk6mrT/0UsK+UiRxf+gLWYU7OJU5PBwf3MUc3V3xSeFHx9Jk
CZ3ZD7nzG6xn+ICvZ3iQJROU3fwnvT5Xk1KY+9fjy1XeWPDvBdRq0mN1XYQIuU/jGpWUfCatYWyL
thIhAn0E6fE5cQ9LR8PHxm7slrljetrRh8/DhcSncFuXraHkwKYi5+rrxza9QyXU/6xGE8/RT6AN
y/5ph1IDHUy5J+CnhvqB7HFVF+jAojYLAl4nHyTW+TcEwqLEg63QOBHy0S1jZQBSlqmaUiIm8/CD
JdP0PKE8t7slAg5ODv1ddGJP+73UMlyJ0NoCrW5CH+AKjyFRpFIzSzTOWX0ktDZQ3jGUnPv8KZiD
lzwvZ3zQrsAGiydUL2P56Z+0Cs4hdY9C2dT783iy5Kn6ACA92zdl6Z1Itkqdfo4t/w+AJqm1hdtC
m9K3dHiaotEg765Hk8lrkWH/+oyVT4JEFzpgqe7JCuz+g9AyAgyzf9btCzwAQovHm1wo/3HOO7j4
zTt8f67PHDUb+a38fni/NX53bG9Ob72wZI7V5c0AmdIkwkbTKEfKupBYAiqcFDRP23rLHCDyKEqh
Qvguw3xuByzP9nCyx3bsQqvc+Dtxz+n4ITkICc++FLbf0zbK8RcuxcHdzD6UHtGxhHFGZSg50yEg
eiAZGHtuGbyFNmZdHFlAhDtwOoAETvp9GEvWdiCJh0ixuU+H9e0K/xt0VGAF/4b/HyofIp8o9Run
om+NUAg5G1Z/05e9Rl132U6LCTKXw9vhjFv6Ft6kNKhiL8US6FJVQDXc4Dz/lfMLcfp1nGmrDJ2u
24bndFpO2+2CC2eWEgk+4sNi8dDx2ynFxb3o3Luk9QF9b4d/+uQUrLizGJQ+Dp496oMaDb+vBbx5
9SRyiOGJkDQs0BmEh1NSHcnBgJ+dqNMtggmdQI7NsRKYHW5GwHTwTaFK64g6OST+VnHLXqdlSlT5
+9jMgzsVGIQCDPgfL3pIZO/KNouB4fdQVs/IJzzGnm5gi0O5n0UGoFumGbD6eUAEwcCzWEe4+zLV
8B2mApPQpSXcYZjK3F0+br8MDXTl5Nbn6CX0FEnc4tOlA8DQAFQWzHPLHj56DlRipwg0qBntKQrJ
P8DYDbIjWDkqJtxOMWTCilwg6sbIMGwRokOpoha8y2wegTshTNP7BpBFkkgkIPPH2tbepR7ODrfc
ZVLDkCPC5Y3NyItCfDyCwMSmTVDm9d6hcxrmT26Oj6ZFfBO+OcG1p9ZRYn9DeXXDoYYXv97mDZNJ
cn05Vbe6i+X5MunGq/dv9+259nqz2NCFtFkNog3nYZzevfx4f9V5cFSODaYSaCZCZqPZre0ssyfC
cIb1D9Vy2U3RrooQBNmPSTcO/SWsJAA6zxq1wwjOTsfbLCD1swd9qYvJAu8ES/OR2n3megW+1krc
OHdiDFCDrbulMAGR/bkrKvaPKVJZdvi3NBneDGaF7Y/rVCZbZ5xy/0sYCIACGFmh0Indlio1wpD8
zvRJH6szmZCPRVZkh2qu6NEVzj1eWe2rjMQYPFuNe7leNjmc8uzujTd7ZGYeWhkSaOuSMlkv+rJb
ZYBArlKnXEey/DTHICF2S3en+Fza1xfnNMBmyOD7onkKGBj+sXQne2bJcCOZIQEKqqc35mTqaA/X
fJdO40mKWwQF8U+GLKa1R5sEDEXhntsqc7/VUTcq9G1zsGgFonwBA6NluXVvyptdI1nxIddt/ylf
HQLEDu+6QJiER02mOeHnRkdsj/Gb5rBTaWPtR3FM29FWl/jAB1lahc5/cZxqho4+mFnOy+lpcIMu
FXU9IiT5pp2RIQu9NKYXXUtB46IikRtl6YQwlFvXLSun/v+khoYGhn7R4jbNhb2Rl9sJiz7HzWhz
HKBoP6vof0/XOk8NRrYGCxION3iwDIhoJklGOKe2VY/Q/9GpZo5kTSYKoScW5xp1Vt/R2KreUdfN
rpQ6xHHodt/u2LvlQeNZsNcquRVNqzGBckDDt93sZ3YOjtl/GfiVBqYMafWFTaQJjzAE+a5CNUy8
1WMfcQipUdg/y5R3k9Bbh38g3StV14nHHSs70BVGU2GqtYr4n8Z59xsKu5tL/rIA7RtbC/Mcqx79
HFWREN/OyKsXrMpAlmYTR2UB7BJYkkkEoOFYGpRzb9wb0MkF7QHitNj2VMm3hdZ8isM/Ba+YpqdF
TdXzqgDBGsLueAu0Uy47IiD+7Gt3kTiaXxPUGTFF/+RVLD1QI4vBBjJSwAmZwPr2X1kJzZZtsR/9
7BreCTRAey6h+oajqI+shpmroJnEH/isa+ORp61jWYoYK8UQIQkaL9dwSKpgHBxL7Sz4HaF0im3w
tbbOGKom60tRcOylyeKgjAigzkQcx8COQ8pV1zmrw7lsH/H0n9CGbpKIjQ6E2gbvyrjwdgsw3Asy
AI5sjIaILei/1zEVW+5F2JumhrLkVWQ6bWQOlmgJuh8u7kFstqaAmW0zUWirpqp2oe5mOjYuzxmS
bgs0Xh9fa5NlAts86MZW9wG0CGCWWb47Xc48MzijXfFMEY23i30WU6Br/QbyKT3qzihm4dhH13o+
Dbf1NuIyBq0PEa7A+tOKZCNlWDAIbES3KWvp3fqg3HcgKB6HJfTh3qT61Pa/IU6OBRSGK7tOc6Yt
NODxqg2qs1Rq+gQeRUvCqh3/9Hg9vqwyNk7Xidz5DiLvWSN6OcNDZqw2Ccd28aDwHJXHCq0nzVnq
fJwYswjacm1xADYtDS+K09hW9Ah/o1Qcr5swKrjaFWVO5KEQGua6NobLSDJcgnK65slgcyyaVbum
sEx0iFFxv8uvqqWmyYTP30yeq4JQjmurLPKwMpmGD5Fgquw3XEpfQ9PzzpIPuas5SDKmyNBV6X1u
K+QZw4y5R/W9r6onH2HDhKrhpp8+bpJ7xQt+qcqMiGwAZpS0fVzvyTii3t2prpHMLukECDeulDWX
ZiuaB1QD480gezfixpLqLRcxvFeGOG/gZ14y9YAEnVc8/XTVOxZvhU4CDIVdEg2WWYnzDbnt6PRZ
pmykMcY5bowUsWSF+gxiatPcrZpC55NXOZQoKUJnsXgfuqEeTbLqb02AHvO70G+JEL5bhDBeOHXa
RRRViT5ZXFExQIMqmR5IqERe8ALtCGgi5Y58qMFzAD2A7EEEGoytgLge84DxXeFyw096ycck75b8
/jDO0VqOAN0SBWqGEFClE0g6Wr1FdLzDgB3if0gCuW4/BuXuEwbGM1M8u17zNO+AgC+c2Kv+XFsd
RyqmSL9wj2MQRWDWhp7BwphycSTHp6uZtxDancklvWUaizDOLmmM46I2FMx8JbfSTh4Qvm4gKb5D
oWQ5Twf6Mk2NFE4SurdidwZKz6IxJNmq00m7Kbyh8nfSrYDGsnftCv3yKoHuhouQ7Fz/a56fPbAx
HJFSwVOGvIKXdWbNae7YJPGmtON6cXqSSY2EIO/haB3vlzpBDkOPPu6kjYR9NBioJVrbklrOMySQ
A7HTcvU7BqRVE/YByw1LDxrapnQnU9sRBJz3v9PE5RnPPo3D+zCyn+ul0PSH4AvkcORdqnk75/TY
fNDARyxrR/zH7qKqWQ1/9waR6fn0pzuwLtE1Z38Z17KzbZeODfI30KParkce8QrClIn25QiCJxaE
7YeRVf32L+TYfIxvQ7T2Lf7POCTHn1rIjip12Q2i4BVSywnVdSOOaDJyfBp3JP5JnUFc8+wQWFkj
y73iO9LbUW09Yt+Zx6VUiemEMwH2Z1sOh6uYF+kXa02ZAe90fbejIO62cGma5u/QborTVzK6s3YB
ox3Fg3eGPhcFxfnSAaurD5491s9apgnq2e55dK3vjd5PKg2h5cLz5WrlQZ14iSGDVQCFC2YRuySp
cpLt/xsKzg7tHMlTNVIlejOFstjJBZYVjO7qP05eBdEAnEP6/4rwb43vshvar5W1pO7B5cWegoqk
dPGIlgXeqa4+SRi81YKkBQ66FJtuS/8TqSKHqrzoPe/qNkp70e+gg6qoRwT2BF/TRquuJaz7aKZz
xfIg7oSJnHqWk2P1m1GDRvzXG+Q2uCM9o/IhghlCDBDZtKZajHKqpobPohfBK6P8LIeVVBE4j8A0
zdc9If7Ig4gsuSl5IeH0pTeexVbN4nrRTFPdg9wPP/mqfGBOaEPcESR3d58vaYslpnrd0H5ywyVl
OKWiPnPml49jVeD/fykSqQO+pFyu7TN7/tdefylypwreaVfmesrY5AU3d5hn2HQ/ksgVb6JFNTO8
tbZqD1Y8fT8S3r+E3Qz9usGCd4UM72rJnUm4AVJ1kLW7lwXiqgD/8BxzO1ay1Ow5ptKPVeekX4sm
/I3yd5STbQgxQLBuBe6cW2cdn52W1QJjjF5ujyUSexq0bntQBWsExGT1Y+4uwUTpHWA0T02SwFqE
9VTb40XkGGm1JV+2tgEranBMtr91U3FsX82iDXZ2YPpuDjkZ9q0aCeem3DmKzZLot2KpxYZkAlah
O+9euTdCAnaNlGAyyZWE0FJys/qgmO3jv3WnygXSTw0sz2Idc0y+xGE3f/f7BRkU087k4PblEPnk
Lsc/ajT3d+S76OW9Fy6sCXf06FziNS21+BC1mDJMX1ZK6Trb1sTjFsQsGfMzddmY/bfBhDSc3S4k
wgJmuMgyaDnIDTuVzyfThToRsr34zGzOqQw4As7G7mug7inuWhh2zlKl7DiBbV8jEba7RiWLqDfp
jxd/GVaE+c7D1v3TlEiv51s2YxG1/Ny+Nard46RORSLYNr/o4x4RoRDQ1x5dswVl2TWlFIr1yQ+u
Q2uH+e3KLK1RUdnuaSyf9dB9OZuWRGLCEwGcj+5lZ80MXwrVkuOIrO4OjNypmddFYw8DWYwu1RRO
MGi44OXfpKNPG1GTOHokr8DW3VAH7M4udyCy6nbWCkuEXL+9WkcN2JV8zcsgy57yziTjKqCCQl3w
TNfsW+G/VEMGs0CsgZMSX5IbmS3Mecfg+e87VpreZbleZHYbRmQ98ri93QiSs4czDn4uhhHX8y+0
LWPGp/jdsmoCJ0DVDGUJCyBE5ddfOW9sHa88ePm2CBh9bYePxBxbMcC3Sf7dAp/rGAhcJm3Si5jc
lmJCTLGsUebkTEaGgX3B6Yiu68IT7ex4yIHx3RTZ5VY60yuFCZFrdOwXScUI1Kl18WXisPFE0RVS
+9RgjpHEtprAIu4zwNo2lTJckxkKQB/+LGFhl1rvJBjQoiOBUuNpGmCm8ZGCNMS7b60GcTJHaIEq
D51swa9lFUuMKZpBzoqMoi/sLBtgL7eGdbGbDgA/7V9k37LITWTw5UTB/3CeV3l7mqh633T7BaBQ
2hIW7w7nYMw/8jsDfzsDOzb2xdRtkh487wdmBNBfQyeT1WNLgVcR7vTntI2kVOH9h5N0ePqnmANM
Fk/LkJ/QUq0Nbw/HDpIfvKgLO6wfbnfwlFbN0qNALtVxbD1M/Druzg1XmCSnX7CAE4uxSzlsCQLp
y02nSuVZLO8aX8FpjsHTX/W7SciKe0giHDCiAreUdBC0HtnWr2KyzJI5zrcWGu097Ac2Ejl2TTuD
cfs/gPLKV7yj4HiWAs4Oe1Uk8EeRlGfsVE3MKNPcqkqZpNp0//oJF+HO2luwwHXicSWktLJJvOrX
u19iHg49Hk74pcTPu7a5vwswlBwRwAvBO7Xxj27kGDo85NZ9GJmkGCkphMHGBBmE4hpPIhZa13DQ
8j/dWEU7puQCkG4cwqmiBHbrwneJTmzNeX6hlHN46HNK3RXaXU9pwHCloUMXnGau8C4IqsPJ9J9B
YTiG/mZGmM5f0Ommo6YyTwFSatSbP6i8d1dQES9YZsFzqE8KHCI75VZjFxn9M2NK6dXJFm1FqUAE
tCgJta5Ej1LC84WcuLXgPSNuKrLz+7+9ml9uoAx8emRE77fSw5UFKy8zef2fQ+0LrqYAmrVBS3LJ
VZuHULtI2k0BKXXiYK4lbshKd04PMMZnT5GylMPuKRIaGSzSBO3DtWWIgg41B95ylfjwdH4jsUyj
pS9CYwdSiun5J7ltuG/PRH03d2u/5hTpHgQxCTs2AIRfcl3Zde/ZBJZlsVBUVJaG0jP7Hp8A+zDl
t3D/9BLEsum9NBnPGhmqME/R5oLejNBlvToT+C+3gZaq2FOFanalpomXHbK72H6chqlCgJTDLLIt
ZJcxMl0qQIJmpODgqzI17uCrH/d/E8a3XMjxXLAyZMUdS1tLkJDS/cHqQo1RkZ0bsrZ7roGuNyWC
18hTnOhc+8Lpa96eCXK6UU/XegI+1WwhMjpplraOuRYXjK7vfN4NkiS8y2tbGEEZW8eNpNZjFx39
0e2N2ldIi2EgIDljbBcBWdw36bf4av303EAemzlvirB55bSli+9XqnwepHC7dNz6KhBNU+d45DT5
0syyqFgVcZWzC0fcYEjYTGbLk1PD7HE4ik/Ff1QUfioGdQfs6MykLo0YqboQm/ArRFO883EqrH4w
FET79RplbcRNU2uzPlguX3/WeTl/S7BGqLWKzPf2Uep5i7biW9dcWxj0yvcsR/0mZSwyiGWKPpCA
zWowUUXaAQ8MzNVt52yFrDs5PowSP1+iuQ4wYQThxaeKf7+I6yF9CZOLYR81T+miZb/ipkPZCvhG
+rh+b9ddm0LnaIXL21MC5m0fVPrDakPkVfDyiqFTrAY6lhoaCMzRv9vEUHr/ivMZulQY+NbeqTJQ
qnYUB8ycT4iFSpiR1OiFjkhyJ6cI3Y75VweHJnqwmJp/zZjH42Eh1snZcLDBP/4m+gt816uDRRTq
9OMfd1Zs5vdPUYd6+NK8GlTsq8pO9RYC32qmx0j5lBZMI1swzxfkvPILyaAXCznhiy9knCSxWYnl
oq0RfuFTWHV4hIC4mO/JfczjxllY75SkwBPUcBh9NzcgVxAp09aQrs6BrAxTaSjOpxt5Q7px/9oJ
voeIkDagVKus52FQvKqrog4z7ElHnzgXwPewju95Hva7GQwCUC03ATwsYUZY20L27we0qC5f6MsI
tk85D2Io3tkGHP+qXJI1IQR/PXegFf9C7/5tWAD07VVcd8D/bogTDutZWIc8yNel9RZiNBphdmwz
OcS/s/HjdaFSqu+Pj51EK4o4hb8ql8FbH5rbOoz4iWbJrSW03rV+2IoJQNz+c8vBXdCQcXhJpMsH
i+MVFwd1GY1NEq/o1j96n5vok/stXjwWMf2+GQHS+vlTviKT8X0SZeSJIxAbWeEYD8Z8f7jK2lQI
2r7wjYe/qlqCAcGeCQAW5Q94dcV0nquHcWJmHjRl7Wc82MSkNUlQKBbEKwD7gk1zc7rclx3fUsJH
rkyisuKLzhQYTg6YueImEcCVhZu452Fitx0C/w/uEcMGM7VkYrXuPalsDoXPnE/FcMP71mN0h4oz
/t0k6SU9oMj76Nmjs/6UIKb0pOWEGdbnw3x1GvFdfDTmSDUDJNuZi1+r82ie8ObyzzDTtdOf7CN7
b8UAnd18wgzhlda/cpTTyd2VU104Aa7Xs8lsuIvPkILuPRgJlA4wKY114f0tkMpw/RIEvK9c60Dk
Ws86xu26HyoY/DGm/4c/NIrcpEL1H89hR/KuKz4nx3qaZkua99uMEBvXrRBOv3Bx7XZZSZ/jL/7b
l5KIN8pSTZ14y2pUel99Nk9rrP5GSDiCFbZguY8YYNjnHAYeGQ/7dl4svMoQXclpBNYA1DBP54Br
DiR+v9jKcmFcDFpQ+v5g8Bx09tpJuUaK2E5djAy2skqmj25+AMGiXTIQzMP9qYFBeCL3XFZeljO6
TtCbmJ+QsMhNzTn8vhLWnX1CmR7stPnymAj0toPdiN4hoOXAuQsv1F1F2rf0N2BNyU9xQuL30Xrz
Ni8IgQ+4NyHu8l6W61zrkGGr0TG7jtCeQPya2V5fYEE7vF/RDmDY9/T7ECqYio/9payyTbuR+LiR
bdilv9TK6xEFPxkxNki8oa95B9hz0yfNxOUbNJUyXMItF3PvAeTDGEJChotv5H1/zZ7XyDfsYHiC
imIpiPLa71LJbFtKCU2g+zj27O76UW8VQJC/Yxj2WGM6ebVL6StWMOIs70+UJKuaIVx8k4yU8yrt
pnxNR7HDqzjeD+GfYrh2wAqp0qSh7UrEe7qYCfj0k+14DNrBxyQeRy2Ogcwox6d/g8lDAbWt0dVw
MFANyYmvzaTxNW2/xDQuzhuHLFO9Ebm8PsFLQbYWGWeeX1VUQVknamXzkDKxFtPmYUrZ2tZDmB0g
KX8Guv+JCrVfS3e521651tzXa57VK0iM6dqN22u7auPD5WWkPRYdbK6gUq8scGHI0vqHQofCaUZk
RXNdFwlvOX829dJsB0979/qotOgF+hOizIn/wE3jBDMm3QW9e/92Ly2em33gz0IdouKfn8a6Rd84
s/ShFTUixV1gw88h0Ys09p6tKDH7FPGnPI2BWDaeYRB3nO8/AoyEZXVW/9wAUtY9Zmy8St9TpIWj
b9lTGJG6LtL7XFUbQjdGRvpber/aEeEh7gsTruRDldgbbAhHw9K1FQyMHqT5Pzc+tSrhzM0KnVHw
NidAXrLW5C/Vsnqk/KJlu3fUr5HhmGugiPZ0tPc7tiL2gZyXPbluG3cs3KKbVyQPoK8VkJyMNgMb
+mEtZ3PrR336BSXDsysRS1DRGwLQj9k1M/GhUH/UlyK9MUO3/idHgzg/5vhGs5oPIcXhpRgRK7ZZ
EMM8afcck7E/MkrzxFb+zuEJdi6gnFZxN2nWF8yl9rUuSInK2515jj1vByb6VsNeF0j/DoUMeFFX
XqNWEy4uFNmbSvFmDfK7CPP4TfHZaQJ/pgmuKJJy/0fKzf9sxhMjCPg+K+ivvSQa/v7iarYtw6R0
lA6QHs2NNR2pNk0aquFjzJoVHS1jcwlYpznHwf3NkYp2BN4HxwSajnL0nld54aZEjB8w3qq959B/
9RnUKzS3bzK8Now8LVXca2MFdgsbmUjC/i4EmQlrDLsQSsF7w5qvw5WoYTkj1xerUE6w2qkg8NJd
UWU/jSPxX89uF+l4P6hVcgRuGNSIse/aEuNfsnBs7yVNBgN8EjwUHsJXdUlllAc+JcfnXZFQj+4n
W1Q37J1qmmP+apXoeAqY2Jfyex9NJVLKZPrlUDPgHr3OdmU47uiBsHW15M4M7yJ3gNDog82d+/0/
jZ9Ew7//WzTqRSPpurm+BBBfCuYuhEBsq+sns9mArO+su1q6D+Zd4tWT07sJXWSq1La1MiCX7A0Q
g+eQrsd4+58jJ8Bzsc+12u5/+W36jU3+KrLmgEKpvtRMYlcqRNzAw7gRfGCUdL5iPZWCe8L6GMEo
k0ZznSM6zHAC0KVltE3cWSGGa2XtrXDvPKETXsrFmK9pc8wwRK1uywYD/CXOnEg7bbhC0UN115B2
paf8qti0UmEXLY8f3CoIq1+tPBs/wghIzyKHdzo6gm9kQ7P9oDw1GdvAlUKMqzjBQ6rJzPrKaepP
99OyHGvBw0yj+Zzlu/Pn37RvC7vYJQnhiDlycjPrR5L+VH4ZhRqXx35nKg6+mRz161JqE6erFyGA
qJBnUWzVF2168iirfHPfvLNWBya5Wt/L9p/TVwHR6i+BVhp3W7k0RkvFcD55FzprnoMZ7tydDs3B
dgKRyHXho/ZDI+Qod6odkU9MF2sUnLo9akBcUPV5x683VroGgciCnX399EPyjzkYuvTf8zOmK6E8
TFSl6kgbeLuyX3o004jfwBeznyO6eK1DAFCZ/HeS5p86xrEcwbOAhSonEjcTnw6YHW4WWnRcelQP
tywF8fy/ABKbQu8GM1Pq5MmRdRgfulraKF3AyOtmSgonM4bYsRLvqHLHnyKY7lb0GG1J6XYgV+tc
K+DifAInXpu4s3rtPVYyFfKxY9sHT7n6MAxT8tIW6KrTUoBsGTJ+A7GLyyrK+Omg2R0JOXlkpokB
5E/MrZdCdFN84JpngMoXFOSKRIG0mvER3LyWjPFT1sMFsXJUJFY4AlsVzr4wigvdQn3oHa8vxe25
D37fCDLclLF0pfUX7a9m7n8beFh188QEy3EyTs8lz+hbTMyfOB1N7XsN4M8JAsO8P8oYuAQyCeoU
t+sLZPTCqvtqWpwnwMS6edwz1u4SR/8M8NXWaTCkmEijFQelRPOimOfdVTxayh7lWcLqLCkrOg8q
t0NbdUqHwatq7tprQDbvNtJeS0z6fYcBbOT+DJQjoNKSazd+TtWwbkTCEUBMGuf1x7asvT5JuvVc
bqW7yLrw5BUeKjg/BWl2u0gLxaiPAuOlE4cugC8tZMQdN9C1eXJasNSzS76yKbOO2VA/1ye4zLU3
oRkDRU2g81t7GuE3kSFB9n2D0LcH/hPLjgl3F/RVSzrWIZrZ6B2uIkfk0Ot+KuPdbwFULH6+uzx9
aCxkvlUs15DYGL8HKWREBrBhoVALT04fvsp5pXj4TyLL4kq7vQJvW4reVk0ZzVQwNpgbtm99w/uA
nnslxfl3UAgIzlI6EiJUIOLkALfjFIrnkRHPfJ2YvWpbwOPkgHgSo4weNpHF808vPsqBkuhYhU+/
R++ecdiIoSAWt1K68dfp/1AJ7WPlLF7eXBTkRZQ+OibC9eVQHCH2GrPwr41H+SPvFdokhWAXaTNm
1K2/83tRnmRM/s9tz1jWL/9KP1lZhURk0dmWACebaaoEwlfvGHrUuXDIoSyAmxUUol782kFyeUiA
mk1LIOayvweYGwTCoZm7Tho5m7TTKZI5f77pAEkDxUX8ttMh1NxBE9MSlYrsqdn6hmuoyHPkuQQx
0WNDReNFUavGTUjUp+lntllsBcjlVNJo/5mBfSZs833bcTmio5ISw3tK5IKBlT/p+ze8AV8PJoPo
VbcMRb6haC5kOHKZXOHl5lJtjy2gM9qFCqgRZZH9e36rJbIly053R5tZt74gvilKl/zRKVoahh5P
GtG2b5qOivblPfm5qroElhkRhlj3oMOHJLiv+vVNfq+NJjXIMSUu67vpkKAgh2gG6xpbxs66wECk
aabv5Piv8dL/BoVdainqHNHKq6aLY+ULWWk1EW1Iv79h5YCErYl6g4Rv+QuHEvsibfqreDk9C2Oz
CQeIPrsMP/xkNi7gCTS5yf3IX+WJpmAr2pMnMIEeOQ1AXbjiasq3J8+WHnFO9tJiB5RV5zfJ7b3G
3s9VBEoVn27mXhWOnC1WbMF7qYK5SHAfxLhKT6VfD1PccAQKRdZkc5waDWGpcb4BFWBDgjKa/3uE
wFMax8sFfugK1U0FAzuChOLWrXyC2UeoQhUwXaI/swfj1/rHNX18idKfCk4nG1iSf5lafuAP3KoK
KILwRSb4d57IcO+ICh4W2pfDAnL5qHDOpC4ZQsvhG2+AhbThBL8Bbu8u5itJpG+EayiKNWdmlCnT
xRriXh5vPQDoFMJ+5Ck6mGzowaRpiL9nVzfLkGWna/e7XBCwsgQ5joL16OqtA+0BuL2YxqkDyuzp
48H0u0wPcSdWcgWZ/Y31QAW6waBKTW8qzl2i9EhrsBozvaBC5GLDAhJfnYun0ijJ1gt/iQD/nFms
9u8PbHJOYjt37CW+zokK6Nt/MXGMfFsI4IVqpBcswS2C4VejxTMZUC61oC3MK0cdwqLgUOUkFQe1
dr76Pl4hwvXUpf3p6qoOxxWqi0w5tHHoMUbhRNUwFNNuJw1l0P5RFhu743G3Klmc0yGh6t0Jir/Y
XQlZmsNrle1fg2oeSnhYYJmjZtRqAW+vqxVmMBo/IxzC1cW8YjmPBepzeawVfCLC+EBf1X+h4YT4
/8HYnLbM7ohl8riymrlpafhATELmONMo4MTSBSzMDO1RkLlsLz9CC+hBpCX2l4Aseac0mX9iV7Wh
e01H1Rp1R2IXObwJXCbv+heEw6HuhQSifbnouN3knFjLv2OgtZ/8amdN9WHtMpI/+8J729y9hjyG
HdYwW27JJMamKG4Od8bR3e6cDONTpUcH+zTzNaDDInQkRItRsNfCN0FLuvsCAT1wov7v1/cZMmNc
fSMS9SBpRPGfWM/G8vQ4VjyUe4bOkrvJqfKmKyIZONyt/KCEfSOio+sBWZXjaqqZtIZLivJK4YNK
XR8oXkiU1+WnSe4jDzLep+28qfmm6Dt/7cZmYTg4N2znWdCqyoCmjHMBOlu5NcjvHiAfSRGKN38v
9T6IoHb0lR/TbrJ7a4nFY2Hlb0H6FFqTzKLtZtJdRMhKACDMRweGng9zoQouMFRkd0c2kexwpbzu
d1ZQJAgBS8Sb3FHnnEFfRxkwBtrxc2t8v231uCEWvlO8AuhUmwe70NEw4ybISLIoyPdZzuVaDXny
lvofBOM9vPAh3CMW5+EBMfKSHFm1IejmfPM0RSNYj9wOYOL3JM/i1oyoiFuOLT5Oo9fGhzdopVxa
wjCEH/LBbHp4bjrWMy5XpDsvE5AMt+h10RBYZVUypMEHI/Yotzn2ol0he80d10zF9hZVn1ncDQRc
fjiyQt/y6P8UgGcSlBB+p6I6BG08rrcwpWSVf2I3POSb021/IIYq9kAOvG0Fy7Uye7G89+u3M0oQ
v6Jaxy3q+fqq4IITmIpPPDemELaJLvGAD1x70rrOcN//rlgjULS6cLfhcVxGfJGo6PYFuby+QDos
wvWMViRdwvSjFZ544C0/n+3/HwB5ttQSKjpfyzyqqHQmtHr1OOBSqw0DbVnQHtWXxUFio5u0ZTsf
2K8URPZUpFHVzFpVpW8O6YRy+G97MPsp5VnweozTCNxKW/PaLoLnvl5aeJyaKX04DZ7SkGG/kglS
4Y3PV4126Xev7af7p+sYCKdvO2SdX5x7vV91uEngRcpzOVUQs4mdVUNqGS2jTIBgnBlsYIYfQ74p
zPTHjGEBX/DrdRRdF3tgJoG4hZ6y0NPQFfmDGmyrm0cdbfFxa5Fqr9ZIctLE1F8uH6wMQCX3ixSa
+/PQfHRQIVEYjGEpt/RqHBAq4TISdOZKWI5HZyOv8dPZsnHVB5BG+w2UM61KP5VLj7ZN2xoehph4
vxm6U0FQ/t/6w282ypwwbV3OuaRszaP7aXDt1+WQ0dGPM0RkTNRIIDaM5gpM3aNP4DW+dDV9YLa7
syPN0IkQiyI8fVxMTdTvrmWSQagBauT9UriHZ3/rkjPup6UgIiZFXEfe8fobJAU2VGJG7AIDWb4L
gRofrvNhejxlReIM/SARokdJg5+GJ+cNpzScrmLM32kdlbCUQkFKpcnJAP01EwCa3QrXcKgviZmb
DR0pJlmW4vpdUCGFT7VNHNpvMc4jaeLNw2lgrbDJokEaBzdNCW/tL5xSypfsvgVFfNYZLWCMlIOs
LFgmKRUIFjKj5Ia0frShuiakGb6D1zLpcYGa9xcu2Lutm9lOfn/9zb2eqndplWayVHjB/AzkqB36
Y+y/zkA1A8gDUb4RrxhHozI+NWCiJtZ2coO0qJobBzTnJiXthHCfTPSOGz++wJFqjsFdY1xTDqVS
HU+DB/DzPk7pK6gqd9r9I44qNDW4+lzIWCgNmXN7KyOEItXDtiQZFfWdcYeQ+E4nPbDFcleBNfvy
ymOe/GfuFVVOralwo12llX1vV0luw4bIVLtuPCqrLKiTT58k1Qcc/1tLmfi4LzU5ueJNAscNz6kl
BQ3RIi54aqRwjNBV8VEtOuov/P48Ot4sQ2M+5wwjki8v2exfeDa8dR00lt7VtljiGAm2wpmPW+3t
bW7/eIZV72MUtFFXVUvRcYbdtZSlw0TeOd2PfjOP+g394DBjK9WsSO6ha2algJ2ehexMUFYs6Po9
XUlx2AU5hxo91eLFWpK9joWi9YgTSwWKNzbbUOIiTpYO2Nb08SY/TpJjSCg8Rwd9pT8n3hHYwZq4
0mVQQWvxURsBxPu20NRlxwuWBmJf8MyMRzpSaFLEWTzArREImSrE7102m8iLKvtWBbzvzOM68Gct
8w0G9z306dPC8BVfsX8UaoQrh6Xph7DOOHEmEgiHbRmSftJgn47kK+Plr7aFrB3lbfTAtx7dhwph
7Ok5wSm266Vco9SmdPIxYHPB7AiC1Zw/T2jzmkBb+PySXbFzSzoSkYsg9bwAT9hEcY2q1/vwymip
KnvQNcSDWfCIbj6GPDCCQ1PhSk5Ao9blD4DGYIE9nf7MywTsDM3Wb4BzAIYvm+CPk7aacSnKigYo
24KmsfAkwGXsuC2xBL/xzAaghzO6RyonHlTipBvTQgJWpNknZuzL1cf7h729pO+y0n/wrbkKf1gQ
2gRkgGWqhkcHhQPo/A4Uw3iyJosMLW79r/tpXrk7J8Z24hjDvSveKvHGJER5ZfxgXe4zSbC4YF6B
fPctqlN0BHF7U6SYPqO3aPPLKoKPixpxLmGXrT7GZM6lk2+rg2RQQMmcx7Nrz+pmV2q13Dj3Y3sK
F3QdKjWZhxSlPyYaluKs19BhLPyOXYze33HEGOr8mAv/bSI9DaSopcMTv99g/Q3UUwXcQ42hOTKd
WNVKMd5ZS4b7oEtq0dohHnhWwaiRml9xDqE+TJNY0gezg+vvB8Lh0OOL/ufDaxUFs8dViQPCtSa8
4YgdRQM2yUQt9Jp/GhqVcAqjYqaliedYYg9Vb04JIoKN2FDtnzq1R9wVBuSXGA1LUbl5BnmA1b1z
Hr9LL4SC0e0s6dZ3pT+dDaknShr2toFjTEOAhb1n+c8Db0vnnm7fQt4ilelVpJ1JfSr/ppIaiAKf
eHyC1zw8kNWV5fwoHIXy27BmT/+uvIYSaiKtLSbWIpkOcw4nDEFJDw73oKuwDATvjONTjr4JvDCm
OWDpf7MHJs9oP5t6MR5LSFGxc212OYRnqimRFuhxmi2caEhMcXKEsyxj4KIr7cQbmIE7EUQkLTZN
fnIHltin8AD+Gp/EvO6fnRKH60Ydd91byEBrq1/c0t6/o69EC3xVTToj5BHMCqEO85tpMkKFimI7
sImts5V9De1z2VvB81n7O8nDpM4nkhU9710eTlb6npcs8F5uBVJoMQwnSxwFeN5jIMjn9tyDRgel
Y5RJct2NuMFAWEP2G/cClr/1/6oWhfVywO303w+lLh02UnWdrEl0ayNhEYXARkOHeEy68s62YvGE
u9sWDSin40GCCCtagVjF3h4HLLZ6HE9DW2t9J0YJanVBLMf9kw98c1nP3NRiPdwXpIAgD8nNWzqr
2H7eAUKmuFB/Kr7nBlxNwrd+na8jQjnE1k6ajq2cSGqhJ1cmsUgoEMdXhfE/cdcbAOyJZqIYOtHm
AJMlA46WmYT9aEGQZQPU/pld+vldGP1GuoJZeFjXL4807OPto9TIC7aNQStHA4Ilr2JudNGuxCeB
YHh8YbD5rBVdMlVXSXLpMd8BmUuLTZGXn4JB3giHBsJmEzczGosMFUgzM1PeE0dNoQTahsAyBG9n
tSKfnj8fBUG+yiENW3HqCfcEuxrZadbGQV2brdiM6WT1fnLtg9+qDU0a5GDuw8gyATfsi09Wugk2
JFIaao5nfTN8p7WEk/qRZgmJz2IajSHHsy5VfGCiK1TzUXq2zAN3UgT4VXoK7GCd/Xvxqp3uJcwI
ABfx4PmW6tYjL6KSzB/IeQNL8rqEQGeEssssUdspBjK3xpnI55qs8P+G7/I3OUwAVpnxX9xgQsiG
TqBQ2PDGvgm9rP3giMbMMPSPiCKVaxbMaYtCjJCnvgtlBLmENv+E/dpMaJDHDRJTuDauuQkg2Ske
1eOhaZJpc5xs6b3NKaFi/v0mDLBorhSpT/SUQUFM0kZauMmw4LHOIH076Q9pb7hUn8oFWQYejefS
ePbjDx/vg7MHsxU3TTpAXyjiKrbrvkd95+fFZ30tx2VwlpoF8Y9Lbjgf79IGwFvj5fE8TFlvZzOc
9Tl5geat9GJ1SuThbjF3fxREc3jYL2jxHiCm2+GvpNo125tRE1rderOnxBaYkVzmqTyOIPdYEPI+
vU2DDXHy+rfdANbWgp3r8s01xpd8Wt2CO+KQFJqGZXEjgl0uZBbYOnjCqGmK8SpCpA0ryg714kIH
bbfT2/K5e7/+EkbIF1ByIRcVI5NvrWmfqO4htArSJ2R0IYASd/h4gsfVeTH//4HWeAjV/1iXXdnS
fMNcNsiFg6Q1PTklIyyQghfUPg6ryCLxZPLdK/xzBOUTzG+oEeHxW+0zyNe6UuCR0NFCU5yxwkIa
Kg2DAEx9wVoGYFucCrynQEnMT1gwSc5MnXVpnB/MssBxAbd0tMZL+YypOIhLOdWqSXWqkRxJWwlI
ZJyQ8FBaozPmTpnX96pd17mYJe7b3IWIDWRyRmNyxQh2wSSTgHDD+kbFxHwpx98Q93acf/37tlXM
7y8VcZ6sqMPFpiZVTOHTkynru2unhnDyyzrFx4eaQ3Ck9ibiZbwNadW8hw1corxu8LRbR5iMpuyn
kLWKNqc3ZOUBqnQCF08Tn1kL6DEjCIetfJank6bIHJWHXkCfoEgJGeDyS8eoNRfGbmbniS/AidnO
M2h62/ib4lYNXs0gcJVK44BZr9FO8Ab4GD8puY6Ck6AXiIAGaAnB1GXa7BGp15B868F2BfUf3Yfq
dQj6z5SVymSgL8A5hf72+NoLkdwDUzFulb4DDw7RYGcXwOk8P/8rgNvU1Gm2KsQJJN3IdBNNODLC
P4Vqiu8bQaWLI5n9+vr/yYE8Vh3Qn2Qe+r5rbjc+qZGIBLymCPLpUeqLvPcSm5Zje+AHWbsX6Tz4
rpodJHhTKy9vEQz4+Lg7XZrW7JmVSAa+JeHv6+spKBl4ugN9NKtnuEO7VOmreQx1G0eZ51vRsbrR
ji5HwOrUeNze+iz/4MhdsRRYrIkHZGKx3IodF+/8nfkTGJgC9n+lDBByJQawz3+stt+rh9lDKWBb
1q/cj5ikkZzuJOK4H3yE85Ha+lI4IwZXvltONzCoS+Hn8PtQbSKItCd6sPksUY+ZgcJlYckPlAlk
QDMy/bKronJ8jp6xfR9+AQOGt9sYHCtP1Tp/XTc1wFC+OgAXQ1ITyW55ZAiZ23uAMLCNGg0MCqhD
+T23HygTRqCP1/e1oMbjMbux06D7tGc+hYQYYG2W9Gc3lMg1B2SMY5d3PMBSRXb17EQ3uZ1mJOZW
8L/unNV015hK4oYtlxUN/34RtneZaPbhlZMY5ZNc72zKmeqUbXGtBSFyRczuF3sIo0K7gRb0GoQc
TQjqOTWpcXD44h39GBtuW7xWv0th0hd4m4WldNhMwxO8Wav2Azu0E46h+2tiJlz2KjklzX0PUUFZ
U8V89oU/QiA10OmRMJXdQtaGL+dw2bUhpc0xsiCZPKWk7GFix0pxzpTCJQ2F27QOl8/txY7tddrq
QAWjn5JtAU7ZcwZn6SCssunY3Ve9q3MxGdkqkkq1LYKm5yZ2FssWNYet/R2ZWKi8TtNQngUzebkD
4UgF8DA1qgQFRcK6w8zkwDOYROtnQb88R1FLXQ85p0wxlIXXviw/xdB0ZgIRo/ShNskFRE/LyOnf
JGDcsM7TNRJk1RRNFGJqxGu5ueF/6eDZJZxyXeFwGZTw2jjN15j28KRbNeVlw4jnvXNTV0b8KO5w
yJ7gVn4g16LV9Icumwr5nvR/LdkfKdx4pLnwjY2XzYzoKCifSBjeYSEVYujzizfgGV1GV9CoFyQf
Xslqgdf1rgHhefD5ZjPYvFI5DEMJuaeY7vTO2BmwXeN+M399TjZxxSEPRV+KEjfP2O8ZJEp239sS
cdr6x9WnESkkBS89x1mLZZurbzw4GuX+CHUtolyXfR0ZDDYhK+cRPG/7FxeY6tOQoZUt9nCoVj/f
CZmS1Oc39Kz5P3zj/iToLNn1XLI0OzFExAZ2ZpmVthzBa2G+9q0/wHeHE8xhwFhMiXu+Ii9erXrW
qLgd0wmHvyXfGRS7kyVY8pDJHjghQxmiRM4xB6tpTZMWapvp01qqpZlaJ9GjY790DTfyEfUe7YW/
SZA9ECHCC8eN+D3s768B1TGuRyOel1l+FQkeio0E41STzgPTyOwPqJ/3qEDu97ay01zvRrCIqu2E
eJ5m6WXxgObV8Vcc3k5hQO4Mpy7NP48bl5GnIpXYQjRd406zTdKqhkqBaqn2G5qXuZOhtaf+XKW8
/rHoSIJl+X40pbIl0rxF4gDDgnPv5HqHAD+oYAFF/sU4ybSgYCBGqXHscCjQW6VqF3+2t0qV5KA4
Rc2wb0ATWLW75/qlAG/ernO1Vk8V7Ri5kt1BZLu2JOmFedNCBnCGrR8jkJImmoyYoJODn/kpeGfW
4N8bKLu55fTmcYfFPfBNRRaGpbyG3f+FlhqEIK60EoOqZ/XxA6trAmRj6blmdVvK3J8veGwkbkOa
SYXt6N0Ltn2oYT+nUc3v2Q8GIVJViYHvQtdMRmqgjvjPJ91TovErmzENh4EtTErBs1x5Motv2LlA
F5tL6zyNsc5aeoyApKHXgvwK5U5lO19t8nfogGvOGe03mRT971gbtXk/aDLHi72bPnWnzu6klt66
ILCprjy/agOnq1kBA1zUB26pfF4IwJBjkN17CXYNSChRmyfQeMw150tXooZ2spUGgzjVN7koLG+u
7/IIwVe/pbZcTWy/vuNzUS0cVdrD0DkOVrlOz2M7CM2qnN2AEt44BjwSE7H07MEvT6Yf1n3BasXJ
vqwntdrSVf+7cxM7xa5Gm+7J+8dmXxqmeZKmmlujoCimWv2tK3k/Duc0IFZ4zU33EEtE1IA/Unhr
xMohRYENAUloDyAJNpKw5zNLieSX/itSyyRZTnEAEMsDd/kDrApauwDDRoxoDDuwlMCyGvNREj5U
67yQ8IHlm76DlQ0OIYMVhR3H2ZGAOdVAax8C0kzkCDa1RQmrYfzO3Dy+ySbgL441WDdZwdn+X21E
AqJtUNUZI/l5amr9/p7eHYVuytlljQVkCWfTS+QMoTm0TyfrsuRpZB0Dn262++8H1pJSznXHWS/z
zPZzs7O0MQKPZfTSi5LI72NNcWctBS935ak20RrVEWZAsQftBTadV0pjcievMk0RkKc3JFkDHzpH
3k3d9i8flyiRLZ8ry7MGn+19mP6KUB2squ8jfrug51/lj3L4v4ZlM3ekEsYzyPzMXguD6N16t/Oq
4FbmkK0tSkv+pOSHxd3D6p8XhEY+TaCkfa0aIPbmV0yExUqBUnpLxqYuoTPZU/a+lUcRjMtruuD+
uR6j0J8Hkv1QodJvwxzcWqjVkD0AiLADc/crNz8jXs6qD7pPCtgJGohBKoMyahBLURuTzioG+UYq
PrQYwThZtssYwmz6qSo9KnGRwQxExH7v1XdsX6EKyNUwSGDfL4uhLg6dONAYFwO2+AztymOpEeO7
gJSaeIesdbFC/6m+aHmNz2G5v+RRwKK9MF1gwq03g5qlpCTJsYqpadZQQkR9N3QsVBHB7eDsiHNH
Jq02NrkLGt53jMSUeCYIDnJV8X0+dPv8B8Kvq0d7n6Fye71Hi7aERs0yRbie/8KaKCxivWeKRKb8
ahxkQNXgI3u41ivcnrALHNyGTTo8kDAfclFNSRnuxQzodHyhtHw47m+GkksBgjkXzBHCkE2EB8RH
G1VxZvy+MhG/oWjU1L1rMmjTpU8iK4KXq2zc1QcyFLhitwNYPRPvNsoYoxFxwfnnX/CAUY9ycY2v
IaixPBzFHnZApTy0AEZ5Ky6IcPaVWn7OL6UDrZAYcrjIRdvGrp1EU7trLX/tNOvIYbTDI3FrY0vR
SJcIpgRDSuByzLgH/HG1L1KXgJ6dFgm96G2Wl6C47+XwyUhK2o5h/BKiFm4UsqQAWiKrtVeJTmWO
s52Hplq5wfMwZXvUMHTceWxEv3LjtvGyWPGzznWm+0uaXrvMfpjB9vF2aoDmKEczbcfQusefdrXL
LatdN/adr4poZMSxaM+3ihOuqA07UZDuaIjQlom+FFKCsnebLDO9maBrSPyG4fh/KSOHJ/3X8qof
KSmuHjLohuiebX+SsJnqcBky2N3bOszpZYDBBI9AGR76Amcm9uH28FjnIL1/f8qml0R75UfrV/1z
A+aCErlzQNcSTIfDluVSG03vd/jpQBvvqh4ErNMYzg1Nh7UoiI8UVW4rNCCx2Jl+M9X6YKJ8fnSp
Z3xMp945aKoJFxe4w+oSU5nU+lcS1ks76X09JElLsGXXtKMKrXqhuuC73i1doV/UEsyWdh/me7Qf
GYudKr/IUb2qqJQv/pNe/6r4Mn4YAm+6pvqwm1O0dqjaaSB6yWrxoqUXh77SxB4F2LpPuU3gMgPi
jPnq/YOGXVLxxnqLFUJuiu5Jx1zzIeSny9smsxuOFcLghjVRTJLWZMV6OEfzhHgcRTRWDBpZPBbi
iD7FBOQdfXee80CzzqEPZpVEOLlOsZxLT3ALF8xZ7JJrRKeH23F7VrHuLn6aMxl0pmpuLM979PWd
+QSNazizBLJhy6n/0SqEZVk254hQ7kVSqWMfRJf3GG1DFGz04DCIZTd7Y+jZQpCs5QlL3qpfAR0H
PH+VgbbSZidwvJZA9ThlUnTq2i4/4FomBsbN4UhA66xK3dPUce99q7iKggLRnx2IGtj9bPg7xR52
djbbdAP+GmtxuZTUkX3R00MGrOdRDLGZV9qHL8NlUswJ7sqYUwLXgEUPxJmmKXsLp4nYMT5BqmOE
tMBOYbKhEisg4rWUA1GMOqR15FUkumaGHcrhciS4mzn7BmKa3ONI89sd2bvApuLg/HKI26J48aO8
HIKSinbxFCpx72y6/nMU+vpHxuTuJSDypEv81NQs0tJQpGX8JZRDEAntBViZ9/u4zoOjA1M++G2K
QsJKcwfbYZWlEi6QNNskDtR2Y5CRdLf11Lh8UZqQn5vgxCZS7yzMzXhWawaBov9MV87RuCh3qdOr
XVe8bi8dUIAaAXnYdxgX4YMjCvVZ8Zn7KiVSSWVnYcOiYSPS6Gwr/n+NvhOyFqYcArFpA+0driU7
1gtDod8EW8VzLvswtpfC5Qt3FfaLXwubBljgvz5ilRgOxlTZbVltvdfqiQ5JAZOWPZWBrDR1E9Du
xv3LRpXcRuAWKGUlVlwEowqGP3pwegjAWjVSU+oX/QMJOyzXQlNDZz3/Qa+sg1xC41sODhEBLp5F
d8aqEG2u1nyKroEdmufVlSND/3cWyALImB0PXhWqqcR5oFNn6n/xZBU511a4fFU38L77mUVI9HF6
I9vyvp6VQbjhWDQeIDpVWbJMGYuvKI30iKgsqUaShfi/KVUKMUGXaPUSDg0qvqRn4cC33EnP0PpC
YzbwYVvZIYwlHlLJ0bJg8wHUMq17exT4/8Lczy7bYSzMHyGLCS2rH3tFB6K/c0ZqWghgcv6OXh7x
kiL70Ox5zTyK3FU5Mszr8CQIctyZLFiLPjQs5IqPq1/YwjJDrIfW6fFhgn2zoc/2RNjyVqqmfGtR
SJ+VUnXDRsgmdt8GUdroQWRvjYEdq+FrC7bEHZyizYhwHa9vOyROJkhpycDEzWoHBru8MWUtm/Rb
jKWN302QKRK2II+llYDPPp79j+WLajlaQqebsS9B9L/W18IipRIPpN1pwPvKf4AwO5cOD6mHvrir
6xzwOMkKewQ+HAR5LYZL25VgM5svYTZs6xIaYBZYd5HzfZZxDgv8AnGYF1wvSP4p+EhT2HwgFKim
C+IcjJhdoBQG7HyO81ijokl6X6rhs4oZS6a6v8wi7gxHj7IRD1V9hltZ70JDobKMYIh4acXmBXpZ
dQ9gzNvFX7Jk9TIvtFrQdTZ8Qqn3qalLIRIbuVAHwNCwMpc7iCgN2x0dAN38ZxidZpbJZ2+KG213
9LR3H3+pVJy9AA6yGuYfptaIkdMMEfnTW8pGqkxTKJHWJSWA7G/mGSTzQtHClHmJGgKZ10JC4Yc5
f0UVFFJwI9lE55uxd3oziEGj3KoD6kCH0TWAw88rLX/if46vaVATh6yclwgsJELuCtjDjdrxLNTb
/E9BwmR933xVlIz2mY8SY/rhhkNFsm3VOtXzcpHyCRf9DK7reYuxp1MwVoT1++pyuKnoVLoF4bu0
gcGLIDHpK1BHNrm3MdlF9KITEi/zrfPqrw2HZJYSZSzEllD401SsrJPwKAkpvEpoMzR3juJ2HwIx
ky9H4phejCnyzxaVZ1tjAuaYMkd8UOioD0W1onRxPNjo/MOt8g03SXMah11DPa1Ha6t4Dyn8IPFZ
h4xecwBf+B7x9auUmLZ+rL/0pQk2/7mokuhn5ucn1u9mzmxLd687dw/NCFgyInoSsWKH8m+GEJJt
1pIkeuKVkeE5FqwJ4s5U84nQ9/d9+56RPEiQ0Xs+T8LsLkqHn0fmQnM3A8Kf+6sDA7kvtYolUW+0
I/wiD3mbQTlHS5GX2881TuqBY24Y9mZ84BHt0EK/W7zkVbJn8iX8OeSk9BUzhxQBcmCPOatCrNrQ
/n/UdJROp3L9pfPnGieqEiHNhpHgkb3GzsqVwxX8ULrzA8zIOSoP0pC1wnd3QvU+thdDctijgPdS
8wBQCVjSfiOeTnKVCPsacmYmIYulGPbNTGQGeQF1lB7oWO5+b/3p1Qr9sUCGjSTpUEEMM6lxkoyG
05YCmyKLmTp96d3GkB3mfbyhN/jVeGX8nFUhZ2TxFJgSZvqxcKIxXx9TFmAduh7u3hqmL60cYqDW
DtwEJ1LS0roGCYRiqadU9jzmy4bddAAMLlVXcnQsB/zHOxZA+bxeb4tpJAH51jgsl0oPb9yeE+04
ZoDYWIcYR9zzmjGJkOd8/JHS1qXy47fqDCqktnQM5yG9HyGR6jdhJLN9exBRStpucVTKmRoPou3h
OXlsOcI9yxEe8UzJTflYRikox4WN4adVUWJqCgk1V1i3059rcAC2GL/mk6VVs1buEj1ZgalU+wCh
yUh1eLltbpqxEPdgmzxKzDd5PMjdxCK+iThjNpxp0U0T+VY57s2Qa+gkTQM9qCJoc3IyymueomwZ
rSksT5+MVDxSCGLs5fO+58xJqgsYt+5p7uBTzcjhXZUNUND7IlT27OgVZjSWuPfOmNetVL+9zb5r
yx1aBRG41TiYUPCn8KMqo5O65OT0ZZrIK63y5w==
`protect end_protected
