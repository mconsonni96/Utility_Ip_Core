`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
EWeJmelyuG1/1Iy+gGu5K/G7FvRo5ohgxGHE/g/UwqZ8WEHhKZmWCTpgprmkHjDGWGn+9VFs1JbV
Wqt3MQgCz4DHvLsGXaQbskj4sxeXu5BkY4cJm30B2uiNVB0k1VgJj7BWlqOqXkSIIx2OCBJ4VZbK
eSBSsDwnvpZAmrq/3o+f7I/b8v11ToE2ySo74Wuq9CtMBioEWX0rbV0LyD53sdpPb6RPXRU/ZkPi
3/hVKW2UtUy86kPKzTyGcro9pHL6Zu3ollJ9Ab/oZCBrx+cEXHmudHw3Uzzj5+VpGTDqRMN+0/uk
Xj5UoubF/YMZlMKp6zGXtaNb98ieB5FNDg8sLw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="vSaIA7Km2vIEmzsXg6aTmyLQY0YDNzhwczyam1D7FOU="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37216)
`protect data_block
Cdyl7TETJSEEfBN9YvfywET9OXPvz9SISK013A0ycfwhGcCcnuZi38K3KZbsANYg3+HCNJuXfAsf
PiKMdutwQwiFSvm6vRcI5SgSH/9YXmZn/A6c+/sn0b9sX9etLE5m3FG5/UD083EkatGrYuGDtW8E
d1h8apCvThfTlqjsA/gVMMZFRia/N5QUvuidDAn8FzMjioheZ3jbKuzwwJNnUTC9YGWLrmqlc321
0MWIDel3qzcZMQwM7vDRnBgAbpRVcHmI+C85x9sb2V0Fk9EsoFwfM+tIZ4EIhXs8LKjXeRWBzJYv
FPwV7fNM0qRNkWmvLfMJ6uaxcYqcleSd0y9TOwi/qt28xVP2yn/Ef750PX69W1OfJll5wjVIpc4R
Ud1F+1nJcONHH2bqir5NK1P1bSkr31cvQ0PMLPHWrG+MdDmKZxRxPcUSD4aKTjUN0XELQt0HS1N+
wG6Z7a6N4uvWdO9AAmutfzeV7bPzuJj5sDQwQSfJ2hviXqRKPpUnr9KdKLM/GSjXFBo4xYJfrb/r
EPEuslAgia9qKR++8q3WsIImL7sD0vzXx7GaxaKIlZamd+GP2AYC5CqgcaSNW3EAwb9obX3D+y7d
thaa8nLx27NojznNridLKDu5G/ZCWlg1FC9elUmoeKHrNxcYXagKrbQu07CgF4s7UK665IYgcqP/
YUrPPwONUsfvNAQNWZmDcVYw9er/Z7uTxuzHBNrjliPUZCvj38IBoU8nbB/64owfVanut2fezwM5
jCNGqF4aSOOjOxTMAM5qcsZeFBgBV/L8wr0foPuKfWxhqCiizq9XNhMwksF/eZ9X98wgqOaIRVf1
Db2M0OSHpSwNcOKXfCHoFkSoHvu1Uy3kSa9a6SFdbshnuOnZhDh4UVtbUpqkGLtWwE4fz58aAYI4
TgaY3qwEy3FvsaG5Q83UU/v5Zsx5mlb/x4MWFi5eS+Z/DwtRrZEOdPh0sAAE+8WmjSYqv6bK7XmB
1VFw5zDnwKQ3+Po7mwkVHO9Z/MO5rK6ooh/Dxi23zjS++Jtc4TjOJmECvYKFiCHnMmrCnrl8Nxqz
Au+9RNG71R1hAzlfr3GGASlyJdJcawsb4eXwMgoZKSOKPhfhJ92uFfxWZJLhBx4USejhLmEZwaa5
t+2JwNgvQFDuWr3w8CzzmQvhpSFOqo2NhLL4cJ8wIlEY/rxigTb8Zf58VDEKlWZ4INsYdgpQZS/N
Qow5gTRfbpbBER91moYlQ0FeFkPHs+JXKLZGN2F1LieIVXJv9WZjaClJDo+I6ndeS0g2dFety35i
TWvHUUEv4If+GZMbnG/otyRlzZNaugJG9bwYiXwFQh0/qAbdfVE07ZRKF7Lxsoxl379qu8K3Dz0X
Tq7k8C4fyXxMGJ60WebH1P1cwA2BcQZBufOQD1oSLWIAwafOkT8Kilxjb+hGKd43Wl8Ogk0Jk456
fBnjabdicfrq/ruN4Br87PjLH1q/0YyvsT+W1LJmd7xjUxpFIFGo0I1yqDT2SoSgent7xmSUQAKQ
KUowg1n4kRwA+esLnYo3qxFYAF8i6nxt4egIJAMRtmGfdom3tqO1166ysrSHt8Um2VS/O10ZD5vR
0/liWtE/iL+1vcEUuevA3ATc4a8QANGAR+dwlBDyHkMbBVTYgaXdTrfjdUdus/HBhZuOWXuB3vIj
2xCWjsloIHjV/zOVh40XnrPFye4TfR3ZC1o05GJhnqjAaVef3u9VK9TnsmPasZZHTtFA2BZTTgxZ
39bT143tIuKkTVNWjfnMim+gwUF1HXB1lG5pmlm5FDn0cx+GgGgTFZZ3KTJa88BCZvHGYj558zI1
F8wCOG1U+/1bKgsctyEhYzmBUyJMU9oeVTrOA27+pB2uGocpCQNBCzNIGw3nNODKR6zp2vKmFe3w
t/RycQhZqfr84PAXXnBQXs7Bpg1Do9vzCPjdqZsRSrJp9bhkVtU+mTfdDrXvY8Yxl5+hgNPxRX9+
TwBhiBQwNbAe+QrxstIwWntJ5HrHnswuDxcqei3Q17kKr4VOWSxKKeF7n1ZFn6LFr8NKmSD3nUZt
rZpytCEupgAl0wUZ8i0hfOucGpnoKek2wB5HBuvORZvfdq6KC5gkwu8rr+5Xilc/TAkuE7cPpaAh
OWOzw9oS3rDsFL6DpMQhe0bx9OD4EqvpezmEU3NiQNNgd5qeb6+lhZbgxNHYEgxlK+EkECp3q1f7
mIiwyIPe5dJcZV9bIJZLCWpRe1OnjMtu4jooYg8tK34XzNHUej+iWzcCW/VyZu0PNfygU8WJ97B3
+THfM9wQ7ynfA19Sfu+fgqDhr+cDvl5sSNsarXJhtpQXdVCtDEoWOxMX4K+x/+s2fu/rWFwdNXsS
rOn97bKMYNjOWVsfpdNgd/byqawgsh8XM59eYzRsp/S4pQ8UNfyX4xh1kuhsqGNS/wBsDJ4CLUiR
erok8bJxPbIL40V1HZx7CW6ZlR3GKWcGUFULzY/IS5zudSEIQSmMAYxI8rZOMdHLh88jw17arLfz
CgMbypdLMB1IO7shcfYp8AhxXYTgg9Xfq9d1bqnFmp/76RuLCGR1aNg8LIlPrTXbwTRWT0l3w1F/
kLwhLVt9IdCDA7FJap5JPQb6LBi5qRhd6mebmsyHlkIkcYAbvrdRwh/7ZtfRW3BfR5+90aX4UBHE
ks8nJXjkFCMIIPUsWSAn21TDUuSS26zVHmADuOaRmQfyV2lQcY5Ael6LgyvHWqw4+e297tv9kzBz
nVeQp8zJJ/mMazjyeFej9BknH0WsciCCZ2I5yBX8pwYj8/z6P6Z05UdVcq2B+Y/nWCSz6sC0Mi6V
FQYpsmvN0p/BZcN1Nze6bysv8TicPMz9DVNUPJGcd+5X8mGBsl1/iwxlSBwsisYd1VdJx/9kJ2nA
8xpH+vVBlZ5ntnmeCuIfCvnH26bhNp7st4IkgcNt1so086CFKSwABqazhA7aBCskiW/fAYCK42GJ
cEWlCYClxsSLlpMcEu7YE6cuUXFOgpFWExM9UlBGcgcfR4Xir4ZtPXINpl3k4v16GmDezDkzcmPY
XzqKlZhX9KhqE0sc0S+rOuX2tvkXGfnI2ZAIpBS4FBPhN68QPGyVzd1q3zdnVzdEWsgSXNPD4mPs
RsLqCFr9GrVdpZWtOHMZ+CNWrvla/4qVMRzaaHLpeqHYVdh/7wVgKL66241v7+cWvIe/sE07Az3h
bQ8xp+Os3rk4dvgblsi1a5Gwv95N+3idDoaPVOBpDD45+k+Vus7sSbAwMgvaJO2luewYLjZdtA6I
PtAtVRZt+oXpNldaiLVLTsOZGVV/sE4y78WnBx9OSq15NL5QaI10GP+fdQdVmnG2psInIOzCbcRg
I/U7ZnOtf9SoXmeVqTFTPtZWmylgHRhZ5vGZC5OGXgVrvZ/PQSWBMqtMulHzwUhOEK6Mr9nInZCJ
7jo70OTutpGp9m9k3Yk4LGLJ7mqOjtfjFg9O362epJU1V9Df+6+Q1Q5zsAvfBVTIDcEeVNBIrX+F
QUdzjLouMQmqijA/UaoCCzO2dNtMtGMJ2TkTmALYHPvd5QLL50S4kiAx03ATAKzM2Ru0TzDhqPo6
e2CStX+SUBm12F7D+9ZOROskSfRboQSEF2pCJyGNabIMfa6BhpwHlYYyCmWA99XQv3MIjJuSU1Y1
m9Vl5Z5sIYEF9HJMb47jQNwi5SeypZw329KDQx6bBb6h2Mn7Q0lX6IikiLnw7WNnHMjvg+XDI3Om
O2wmqcCz4tadnaC8pgeTTEXxvrt2tp6YE4+tAjhZh0x7eLB1KGTjJFditEwd/MW+WmjjI2VCdyxF
ca9MVj54AToZHfnyFTzhDMJFy01H5Ql4AC3utp26BSnoK5CrUop4v9QMIK4VMzFQNvgA8P/V4LuK
CS1D0Z3o5gA3NBQ6CXq9KX29etsHLarXvQXEnttJbyssigsILI8jNxSJMhuYqsrAVFMsV24RfzMF
NF+3Gz/he2FnZLLo0ANeO67ms/OBqJm3R/zkZwcaR2RQ1Y2Wc9VP7PR0uVhlfo1ZsLdu+hzCgmQR
kE9H3Cvc/ZV9OVWgRwc4gxxOhOfYRV6fxiZw+gtqN+3RCTAW3/9dYdnAm6YNrcw82ggDdTwNbrKK
IwnuSKa9+WN3YFFDFzWNRQ2lZCHvomQ5Z4xZBdBdFIOkInb5nqD7ey8Ip1X/gWx242Z6YqrR9gtG
3/Uc9mEUtygeSFqOVhaM266DBpaKN0aJpacY/e0wXemLsrZOSKZeAa/Ea5GbZzK8y0Bl/N9wDiiq
tZBKMyJrxyTEkCXJl7OUGDPVQKq5rDGVkmZ9wKtmwARUPJQnlR6ryHN/Ld5rQOZmXSUoN0/NHxxh
KdkFnvXa7fqDxsdOHUNxXFXmbM7mSEsWCAaOObAq18BnlOTikQ9mggqgoADXjFbVxrryR/lbQSx3
Wben/5dp7UcHlm6kZumk4+15HCxXEPzD2tdWJOAh1MkJPRdB8+HO/G+LcqO0yZRvuJ88wHusLck1
c0xg+FTV6uaiEA97YaqVkJ+eLxHXanW3EGJh5a1zCDBZDVRbtEj5MuyYVU/0lp6WwlvpzHxRMCak
BLX0kPww2SLRaaz96rO+BT4DYEiA/OPHTkDZ7xT+hTTkMN5GqSBSgPcMaYJs9qPmMssTgwqKxfT4
wmga7QbOETs/JQCrSN3C/On0NBN/t4/ms5ryt18ch4TJnd0MLny28g2QNYzHa/hNaALEqw+9CmJY
q/s/wFvAYq0AI3ogsVNvJbiX8mkcTsPuANNx41u7MsJKwSHs8bmnPR/9++VtFt9KiNc14WqkZ/tQ
s6/3NkaQ8DaWTcc385O+iUH8VvIB20FKU01QNpLsTeA90N2r6xTmfyHYwpf9hE5R0gvdPeUDBqFi
GTrea8fwJPwdSJvyQUk9qMV3aSZWeMHiZsNGD9+UQUDr49YpgtQhdEY+ElhXNHi9mpf/6HgyTX5E
wYqOtYC65yo3bEZd31wEekFxLy59TCdhMQEwvN0dbp3bucXi7kQ2JR2g+WzpbB3tmFMiUxdAZLRG
lb95nCecda29z2utEcAKut6Z2YSuPCQqquFlj0XgX72RXrXUKSjqNXmhET+pyc7jdcfG1cpC+91f
2V7Mihl22bI44gkmJPrrajAtjQtQznDQ+DB8AArv5Del6oDgcfv6i3k1cIEYs4jVqhwcnKCP//ue
OWLrZbwG8FjfXm5e/BDerPw9Wu5uGe2/F55f0EjhUTqkvngkrUSVRvR139g24NiQ7TcmD9SenBVW
91IFacDtdD91m+Y0J8VN+yRJZyYCQuXNC+vbR0YnwbIrwhlucwESu47pRwSIaVLvJ1pqJ2hQAiG3
Qu6RRctx+XkmffNEgny982XRoiCd7CCqX1gvxkAS/SoZkzEX/r1DqB8IzUkoc0BP41HHKbxbOpZ1
gjrGF+NjDJlZezvnwrR65Rq1VKgoQ1D4pt+B0jbMfcRSCb2pFJSHsp5rJ9pgzHG8wG9FIgGgI/JC
jY2ViysSeUAp5eUG2Ss9yUC/ViZfhuSGLUAjVYrx7Dw3TvC7xfxFsPNip/dn5jd9O/aQa8qdNFt6
sfX5cRO8DjTuNpo7aIP8PvSm/Zsepfha2UvFDQPagAuRzn8CCgs4Z8hXbOsTCtgafeJJ9wZikqq/
p2GirNOvx2AUT8EXoiZ4hUfFbE3HeCEsbRrQ7ievBT10IcGAM5QD2E6yjUlQETaPW8edLW9KXRyB
As1tADxzcKOcyCYCbK0Q/gfqkM25th/vnHAM7idjPzNPivukM8dfUC71oBwNDsSUJetngqRQMY2e
VwG4yz8SzOJ5rsmQyQ2Vomh/naFbN+p5wlFe5MWy1ikLIgOvv7qEAKu6Akd1wMOG3dXnERj/0m/x
PzOtSSo0oq1RZai/gOZI3pnPZvaw5sb9c7aqSZK+0EEBfK3+C6iJUFCjYsRrAEd7U6sVgiwsi7Gj
S5RTVP8hw1VQuK1scCilenRR0DU/+UNeRLYk0jpBun3a5SEiDBvGLnH7DMRINwpFWw2iUpY+DvYe
mwnpcIM4DuyFXHBU0SdjWHO5Tr9sBVDZ3DNcOW3gXP8T2W4YIe2jL8oBIjr4wnvopyvYPGwdL9+w
r19XqmopGil8bFL+za/jjifLk7IjBCn2z7rFjFblPUNA281IMAIQKSJC2kITK7dwkuihoOHFxeL4
YK1xBgK9ewm9oRkAc65s8dOHr6hsQXY9Jif3nyjDJLgblx+XWS6xtt5sFMFJtgPk/qO4HbuU0nWt
yB8FgpE1mNAQHBxCxGT4cE3XeKm9vAf4ZQbeH+VPcnymRe1+dtS+HGxnGkFJSC8YO3lLDpmNNiZ6
IRFROEgLWIJ81G8F9QYWH5K48/uznvn36029w2aiQv32LDbBiFLizbGQTv9uFn9eO9X61pIVLQRm
RgZQuU0RdyZ2ujp7IDgdrorufBBIiBURU/3yX7L29fYCvQulRt0oo0OruiSem4dGcTmZsQ4fN+/i
dxFRxMMBjRtujEwhs2LhAVc5qYAu1AYIJBYk1fymTDlxKwAhtUym8KoEFcr5Dx/aW4mSyWkNqoYG
ZRAMO4kEF3jt5U815YCqhMHYkYZJOas7Y3RbHdp7J4ShOztiOJSTdDYMYAS363HvcbI0lDkW6oFH
qcxiF+WXdKTY0Qa7Vj40QL6K+KeO8PIwGPvFiJQj9YwziQH51ZKSDuW7TIEUu0jSweas/euu6/Ln
tA+dgBsZs0G/nTm/V+XMH7slrhAM5Sasah7R5f3IWCUwTnUsGICluV55TDnc5wjl2IHNznHM8ssu
U7bGI4xAF1kAXYwI0003SZxycsxW0tXkMeT+8S9FJHc9ONpO0kOTcK3bm3ylJpxFnKNdWJN8KvN2
qz0ZD9D7Ze4QPDdcSvaWP0Xbw1UzzbL1q9fv/S4sPohywbwWGu82cDAs6HzWVARJmZdE8efioFFJ
PQg1BPc+Z4DzwUirnqeEbRPNTEo8+9pknbgq8njH2eng3uPKAtSZeZ6br/TCIjAvAez4LHKcXk7/
+CmmD38Ace4z1w8ryLfeR2/9dj6/DWi0eXbpbAWKyRM00+Z5cWvgwEaIM47abDatluW8DC577+Rg
uhEY0H2MDkgpnedr3K5eLRIoMTZ5pXDeQQaU9rceV2iihd8/022xrR61EWpfSJZ+UDJ4EiO0OIGd
38IetG4I9TkghoWC673BwRHYmf+1M9kqqnTE/TLIHy1h0zfRPL19rGMFdWSuO0f+odvZZ5M9qy6S
Mvl9mVhxh7IbyStPC+BuRkVUKS4j+KYW50ZNf5QvML2kUGELKa02S4ZHAdS9C2rSbk6W/57Zodj4
w77KlJtBPwBhfq4B/uanz23LKxdcXiOHYZbKpLq2SzINJdO3oSpdoEc10agz2WRc53PTcw/0pbbK
nPnBHh9MgNKlMNp29DQxfpwmmKorU6Wa7OXSnl+RiE7rPTAWTvr+LOya/TFYgrZFIffKkgwY8sRP
9OVLtCQUobHJ3esmYPAbRhwkgt5UuCFUYxh42QudK7loH6dxHfen31wBg/HP70vca297l182XXoi
Bu8T+mPjJj22zgo5YvFZyc0SCYbeeEoH73+C9R4nMpRmWKqJescO3LzH5ucRXIaT7mYlLTMij6Lp
iYw+0Hmwhy0qf6p/301EjAGokLe6oCGzKkHzORoiNCdG4yRIteEcqVWAQtcc8XrLx7JiCFFNbH5j
+KbnMr/M+TOjpSLE5oeuRwztoYIACif40V7vlrE+2mJw8WRzRI/IGeXZ9s7C06doi9kneR2fyfpy
bSNg2AooP5oAFSrvDdMh+eIVNqYmGUY9n514lhcAfee/e+VI2BFXGKmXtZEEMdcLh37dzeR/jy3t
zc5KrAkGrYiYcom8dntEIrde3VSP4hyj98bSfb8S7jaSfgqF6F0gRbowAaOJmwBo+/t6G4ycgfEz
7UD4vAazxUB1V7jGQfinBitdhLJ9ZuvsYoaFOA27auNDI73vT1nZqk6If1WVx/jNA/RiRwm6qFaV
ygQvBscXSFm/NrWFwjyeGaCWY8PfkwjfS7or71bhfdRD2HLwKUJB5saLt2Cb03DscJvBvoG7zJLy
vtFv62XDPVrOL6j7wTFre+fIIquQdDhl/ni7qVs/kPp263jcRAtLIG2VeLLUwWyG6osuQSIkuvUK
PWkySuNWK4AQsKESXTHBwFop7dmHJDVPYqmiuEtGEU6RiU585K0LJOXyC3e8ZIB5Pe0uATBjePsg
6Yt/XSGzRVuRNxdyqxB/mV66BxGVodFnowa/rgAly6JGlqeW779636sNNZxJ4COnpuAreOL9dumj
65W8nkUB4G/gkoh6PnnAXC7J6eIfX7CKldGmb4sQeyGPfeD4OGA8CNWoELDsrik0KPrNM8CduvBs
J0oGCbrWI8aZ68/gByYZcwCBmoi2uh3mTjzMXE4rQQj64MQYKY8/qR4l8wSPvrZKcJkej6VJ3hlc
RbcgZccfU2Qv2vf9ErFTF8T7ddf6oc25v9fs3UWa5iA5OW2vrz1kcwUxXsTSL/GOEZvzZV0jtK3v
8PldmznNee6Jxfe2siSRE3aKWbe4JbwGFDMbMqJKHppaZNuIT4W/SjHTQSCnjI8XwPfeHkuO9w4n
CipyglZL3mJ/2Ygj6XqZT+B1tVItMfqffJyDEVHd1QR/HmZnsGFED60xPaVC3eN44LvWIHjRkx3y
QwNXiO5porFgG1kLcpCeX/gwaLz1ej4qUX4GhXZF31E0ApCQtnNKMlaybkEi0g1GWMTmY82U6ffe
ANuNTA8cmA6skmLsW+hqg7xzT1u7BkeRcmodldmAPhVVL1PC1BEfGBBUJ5yxMSU/8cOi7P2YpxZt
6WkhkrtQxFSqYmGHmviRyadku9G5gYsRCL7uK2/5qmoOoEghp3O2dLoDZqJVy1uVoM2gj2aG6s4b
fRgctuXHwKfm+R9QM6naenVYB2AzjYw5LUkqoEbRgvG6iWeG2ezuzZWRX8VhkwrXDi5O0VZ80W+5
QRh/5chqKHcjYOPSpP/fjWbLB8uhoMpgI2F1xJiXJp8yiMm/ig/8nXQuHE36ohdXbHy8UV0P5i29
kEuZ/uapIhwPm6IkmuWqvnLeqdUjyY0fJlCIvz+8aoEw4FMIQouI0O+uhKe7/InlOoPjallz84ML
4E586tBd3FtbilRs18ETHoRGF/d+vaMtn9luK3vARA4Zt8rkdC0vsW+agQUQ/oKP2FWrozeXhquO
XQlNn/hSoGtzjr4oK0bkf8t5P7aIQMAMQcrg/ri3uprmqmCIgr1L118lwPcqQ+o1hrLZOWq0cMRO
mlrXGLgOeCyaitHXzjGP0u2vFmdQ3wPEal2sV5sFtxrD3eY3+fTUnmbg84XeH2h49aCdZL4Swl6u
yWftl3VQU1PvAZOkk88e7ltrFleWW7VGAJmEawbww6HT7xSKIe6HuWjtGAJgqmyg2OIlofUhB3Dn
7ey5KsN/xib7M2v2xYHX8elDCaY0RINQmpcEeSeBBk/mInpah6F07a7lTYoEmZnhrN0XUW9oUhEw
SjvpAOAgams3FPL7HagMLw1WrsbREEJc8J2kXd1y/DZZXj9jqHk4MS9AVWgZTPrHkY6R7GlgsCRX
t8uSyE1n5/qqK2dHv8CGPSd1trPSGB58Bw+KZWACQFLPBD3skt7U6GB+D+dW+B9MN20hy3Ym6kXd
RLpFD1IcSm9QOY/FeIdwxoJf6a7M2SGSLRF91OCD8ho62Jp0G+eTPXMwwYWr71WwV4BSnfNNvf8E
lWo6CJTLbuSszUh1yifGRVgqZT52QDOFLCmwl9jhABPxgJQ2OpAqcgPpBFskeXI7dFxjgMgPB8YF
cCXSOgpLIqdJcYGaRX3A/i55sdvVNlwR8ta/qRrK099xO/CRD0wrAPZT6yatTpGpf7Ke5UNE+REy
wmPvSpPVsA1C3XF7n1sB+05ZcQRHDIk1lw9Sf2f9pCxxeiY7zMuhrFU2xki9rdntxryQgoeiYiV/
8JRIL5odHBMkmKv1boJLcLkYCG0Qjl7i9x7ON08YqnjmqGrTM/S8IHI/N6VVZF+zcXFZvSUwBSkr
+WVHiEgpWyW2tuQgvjIAEZTYlW4514d/fx1yhAl/BFZJqYAJ3PYN59u/WrMsnVBC4gZFNXkGw7nI
b/fFbXiGyJcWXPHdjEAPs7KdM/9bRBfc2ZyTsggZeS3WqSbWRz/VbCekB55DvnP9u/TtnCJ7osWS
ZuGKxo7WDKy49lWIsorMboxxKxAo/bWaa0+xSTnDbHfifbPxkPftMmAQ93wy41xjrVn+BvXXVp7V
xbJaxSe8WWgJ+EWruBoEjLH46PoCsZJcOHua5BHhFcne41z9xwVCKcM3fpcDVknLFRDRZaQ2YcfF
piaJSUXKGbwz/Trsre3TxUEffGQd1UJnhxIL7wzCPJNVSYhsts3aarRzN49af+qjHU/IPsGQSsJh
y/KXm3/Or6ZRlWplwgRh1RFmTm+1FhB6vTgnUem1750TOYMtckkfZVHj57IlRTHu5YRzFh8QJTjZ
cnZr34j9UcwzkinadLNPRRCt8ifoiTDdTAjZ3XvMiwHXJYUW7bl0hN+EmuYUzsEPBoRJjj+HBd1z
KJ5EGPeSovwuBAOeuCWloueUVf2P/LmdrhYYWWfzpOI7neRG4lbuSc8AaNoTrE9QvIEhHKeKEueR
d7trb1bOzQ3agcBwce+RIzRjw/Bi1ugUJIbOTQQq6iBlxuaZVZpgSCh6NLhKFTf0MMtwlVnJ0Q6M
9/NN3fbOUReIUUVHGcmllTJZcrv3G9VGHa8QYNh4Vy3v2n63RWUwOcxSfKgWf2iZ4m49XY87fufQ
xaIRiFqFrsuDx3hPE4YlxKk6sk8jQXVXMtH7AsIf0Yg+zoQVUFCIbbsH0qv5CMZBLeNXUXD8j6+l
axD0ib4laeo/+eRCfUimtIUrqu9KjpYJuML1ZS/XFstuPlnCFls/qx6UCi+ppjFSMF5kol9fIDnQ
B595YA/+ynJJN/RuQYURm4j1wBITwfrA/1sGCHlCHXcOPZKrfhxArsKmKLHWhKPcCjTCDK0Ym70y
QcMOLI5RTBRKV01thzMfJHXkHyeP4vlxORm8Xmv6qfk2OgB6LafVkThSe2h5WHMG7bDvkofvZZdn
/+v2p8TVT+BZ5fr4hMZIDHotdGO9nbdAR+mA3XsNLr3b4Q2e1GtJPMh5PLyKO9cS2bB4i1zA4Awn
BNlF3zeyVcXABStdeZDEy/us4M+cu4blxO9KVSM2qEOtb7OanGZ8+7WwKvSSDneHDsV0UzL1YuXp
QmBqy4OdZ2M1W1EFCKH4ODDVMwtg0IR3+uNxeVoW8nP8PEiH2sAGqxnTdwpLHuFsil988REMScmS
JTtfOqi2XiVpo6HPMVaIKKHow4qW3DtAQsY9QBSWuj3Crcr+rGsXC1S8EVSy9Ih7wSoj4s4thZm2
/xApvrJfay4IV4/WyCUcCyb/cRS93wrLbkOGGM3onFTbRKXmvQvuTkFSN8EmaJe0N7r1zFrypmcN
ZBcyOB0dBgJjs3EMCrFaj/IklvNFmLWjh2ZpGqz3sQO2tl1O+oBp2zxqLNED3z3byMaUF9oxWAc0
fz69ddCspt7q3GI6nG9El4cbUDdKdgOElj/8C0lK/RsFqh7RKvoAASbphta877fGtEkeVQIYpBA/
0zxgzFRs3fqPC2T2V2WgP9J7dQZ3fGYIu5RDiBXfNHWSyrcQvNNkx1ZfZG45YG7/tuwgNe/Ex5aD
DXusgK90ZgRIHNpP3CUOAsD3k2KczaRA8cgH2Wi7DyuOj1ZxPHhdTZQtp8H/qdYBAIwExnyNfFGX
46UYUjy1q1jfgbbRBF1YmEew2wAnvVNCORHSV1OHS56UvZ8V/zh8Mylw21J42Aou97xmdOE4w59O
XD5EcK6klbBXU8z3VPD7FN5AiIXKQ/+C5adPGl3zpqnvyxms91PfOKL/Y4ESKBqCmqgQYJgTGhpg
07avov6nn7zFTwzPlZWG+EStmbX5XQBMfKEfMmHX7rTb5YjpMj7+en79W9/ePkGdCFngFyAKj9xX
dxVQC5mcVCbYJvJq3AGbYZmIyhlmjl3AvHYL8EgenVicuGEAbIseoCr3yFyRQD8oYpbh3QuI8DA4
EUFf4k2IQbrYWu5B+1wiVRn/P4bcB5AaEUnAt3Ie0ik2WMV9PQ4k8DLk9lGfYm2fJqCp32cLJ7fo
+ZZHt9uhx0J+Na5kQMYm/HNNtUQTxq1Rx7ZR7PB6phRm81A1rm0jvaquxEPCHSxMxouzyWCz4LZ6
EVQrYMGA35cTSM4uVeCjQ+Alfuy4S+g5Ullu58sPGPhoDV7SucypZTd8aFCn71FMTBrBiK0sAg7+
JExalZZrUsEE4yRbNWnWuciTjR+2RVVVchfVRiR45R1slE53J+V+eGbToijAxB3Pq+8XDf+cmc5L
Xnz1YTH8bSYTuBu1rPMy9c3ZEfix6JX3CR0PBdwhGxY4xM/7Di2PYdssMbCrrnPJTS+bFH0a7GyG
xugGYMCCSh9Ou0TFjNPKsYi3iOONZTEUoJbikj2VPtLcjooOojXdvPsEUKKDV1cLl5Fkl/18GWbU
fgfyawaNAHfDnYmily0ixLZlTuuAWBvcapEFEWi0Be0FHKSD7fbcnRTybzaLA6gtFyfA3g/TRkVY
EhtmRZj+ITSzYZDabJa43vcJaa0Y106MYPnX6Sa5oPctxIyXeFEtkaxiwMPbsa9QYKjdQYPYPTCy
cg2KlK8Fs0RHpq1OYcrVXTdxYxmDXUiboJtxZkyEHRo3yI3JbgxCXdaaaEefuqkENfaVbGiwfbn7
XN/GfAF1dfzmKVsYXpvJLMev/Z2Cs60mzIWICxH9akt8sH8BQ1QlMU2XUpeLSuPM6a7BPx2iJ8Z3
TAoqVbuzECOF9UowZ4ZiGH+gyz5VKed/yX/uOJ16ypXZ1Sx1UvNWj7FQ8xnkaBNNED0j6W14dgEj
saej4tzC8y6GGSpJW7NpnTLDFMloqAh4xoL2P0hl+FyYOHBhA37sjnlB7AgfHAZGfMszyoCuR5vr
975Dg+eunmLf0R4NoZpoBQUK/KFvVhKkQRqhNdhBE2NEkRdsQ36LEQOW2N5pLE1I6rLYXBY11xyV
PsdWVtfz8H7LRvZgq1M4WnjLbFKQKNX3Si9+Ng1ECwdpOa7j7wFEGIZz41QiPRMxBYoPYcHMDblM
5KWXhnx7ijpeHKR/Np6yh109aNq0zte9ixIFg/2oIDMgLfbC7G0Q8Xxf406o1TEAOhzXQTdHPGeC
rA50YY0hoVl5qlTIUGxk31wp/V6s574K9mNxbHhVO5pZlUlNKnz3wFhxF4WqCxtwPYuZqhapc1ST
BQhg2a9+AICgKXJKZofKTHDK9NieSUmoErFhfFYqsXyWld28FNSlJSyEawptaZS1ye2l9PUtgN39
iQ9EdP4GujHLaH08Ly3J4vyAw8MSmM0oyo6EYDbn+yH7EcFHMQJbAFjti3uEmflWvSQSmxVSybgl
wUiSr6BlTcCLvufWsYi/6TDYKnpbElqW8NUbXe4ZrGgS6KCQkbU0RT+BJhmJhIR2pdrMsQV8mST+
iE1z3Ac68XtkXyjLK/8vLk3KrqN3j6zLWl/BpZxaphMcoWPHzCia2i4wOej68UEi1KGlIvo9WGXA
gCxnQh5Ow5/UoOQfE0XOYyRenuKbOecfTwbN8pqj4uoR4yJQgBjUalC6sWrpC6jzQ3DnJVdV8bN7
NBCzVupu+I3dEpOogs/f615ob3yCTJXRssHfX1UC17yheumSx/4OODytNR1oHdpvtT3NfMU6Zqhe
db2pW5sT4vbp3EdFhzg5WPx/4i+uPytLKFOwqKuG+WmXjl2L+/yu2or8sfAHtt5onmzJZO6bnBJW
1h7GmyWVL9me+coLOTyUyPEeZHMP/tXxjWrjt83+8EEKqZtJpHU+7Qu7qbXprBgZiPyd6Xy2G3Di
8seuH6Eal5MvTE+1EXO6FrDNgOeEbiu653uluGz2MgUudhGaMJ1HfKUnraOszVkX946RWN6mxpFT
wHpZ543Dlcp6DoJ54yBn4AMTC/VpCU8wrBN8naZF00Y2FGL76CveqIy3NhDbG2v5ixSfPkT5aP+1
5Kv+GQyxa+34rwp4FYun0m+a1YMKMRFNl5PoKYOpLlA02KGzR5NJJCOIQqVQaeuVhtroGKPjZo+B
Wh+h8DczCHh+NVd243QWIvSdXIH/Up79nI0HJy5gd/gahkZt0aRyUs8hnNIAE7g+pKsZ88Ighoey
kMQu8/PsSbTyZiY5UIohxXsVEMpsUbfjMI7bwTdN4wTRh/GprmJ/dDfeEsUYVSmKeV2MTHEKUaPY
hISRHBV5JI6Bn4CHgFzqWy006aXAQ7IRAoBnnAPCqPGhorsp7GnN3FPmKSmibWa3uPGxNKgk0T7h
U1lN4TN5mDOLFrBRrlf1ZSoyvbfAe8mrOplB6OcYajtR4nPsWvVN3BXBTXeo4PvLuLFgaZwHWv2K
KvW+sOxspcYMkboIZC4G2fvrhdhtEW1RbMp1H40E9biWrqgYI95WwcgrUxYldRJa2HDZu0005ta0
opCPGRb1QsygJSGO1X8c1ot3I2yCPLq7I6ldcwc0iTkXB+xq9cF8GpDLT9Q07QROf4oAZwo3A/Lx
Jei5MBPewVPEoY579vHIaVR3In2xrUA1HhNBxvz46YgulvjGKXKg2w5x6vIbI+0Cho86a7D+6OHB
6CFZ50lOo4txVXj2Wno10QEcF3/FfBFM/h17VtMq7eHYc60rAjmBch7M4TLX/ZO/GCiB+mPCjzdP
o9okLjuwXxPWTN5XYSBWNYeKjDWlj09RzHrjjY3SnaKc4XKoYJtnj9cu0rj1NoB/VFrkWg2FvxQ0
5+DZQPzkubSHS+/f2Ma4RTSTMAiv27B2dKRxvHk8VwA5KhRdEmPf8R4UJRWIVQBZOjoAhfgAO3uc
wo0FSl8vD3FUSLa3A0LAF7D0gMCX+z1p15dq40laP84xOys3MkuQYUjaN//BNAwDcponHaviI02d
I+PCa0bgA6nHgBkzg6K+gnvmraVM1sJqX9Rq/Rab/Wyobk7kqFLlWupm24Wcwux8Ad3+/vwRclB2
KnIszIRrZFz5ZzhmqoIrZUVvtrf2cc9I+F3TVLjzQbckBaZfrq82HEGaaiwVIvR0943De2V0zQD9
2X7rv1sLWg/U9Crnf10EfnGJEXhmi1PVydu9elL1n7P3W9Bez1iOVUgruGIhnbpqrktiaaTU74LF
kXOS6tjkjwWT4VnAeX71DM2uQdqcP9mEV0fV8Jk/3Gop4NfXbxzZZrFHlfz+mvArATJibw+NFShv
OcW8ntghWb7ZXDwU6a7sNxyo0CxiC1XZIxYuZQnyq3Md7G3FWtPhHwMuH411UmGUIGtFNIoMuNLt
gRzw3uGxSLrCBpDTJvuqdErFkoHvyrY2sYpG5UzvFlPj/KsgxeTWxOl8T67z5ZYOVxJ6xa0cImqm
1g4pDA2bB0qzJa1X8qvRGA1RfUzUEwhRgo3b0M1HQq39XRFlL4s4iTj3P5SIfBsZby+EgkEMkbIt
q+gmEaQbVLH4N5/XLLW3DDSnK8VufclTWwt5RTbe+SSsoxee4H+WOox/jQP44JNC+Hd8DzbAoJGh
pSrP4Ub7dn2/Zzn/R45p21vrS6i3gH0oq7788mtiXgViWLzxK8Z5hJAz5PGFirz1vQTHMMxKp9Df
oDx48Lo1lGGD240QxTdxRRz9utFG2okFV9c7fedPKibYby9Pwt18dTk1JhmIRP79Un3tEFIA5Dzq
7FrxGYx2UFT014fSFI6kcSRmE9mn/uRF9mOZd4zLkrDvRmoo1q8ESBQ38PyZR8qRcfJ9+iTEQK/8
rqHZX51K40Aas0eSgkEJ64k5XcJf9OrUcmIx5qyrA60g90zKNPllPUcK1KX20c8YO4A7pxZH1aHA
9bJ+WVxk/FA2rlo3vYW8pklpqEI3a2UwndLmFvaCMHCuuVAHyai/FxtQSvU9thXJyLMWYWHtE/Rs
D1ZEAV2pD0qoAdsb4uHpT9b6QJxrIxVhhytagHeV/NXyxJ8B+/0xQlW4Ao/ErmYrI85/SUQz+/qZ
2K/TaMxdrqf94rXGbSSu3XbwM4+VmVgC4l1Y7yiGHdjfUMqQPlcPfDstXd/hjAbOBVxZkW/XYP3o
2ogRo4vn6Q2kSq3RHYKNPacjOqQ+arUTKeKMOSlSlvkX16FQxsKBw/lVv3HUouxWAUm01kqI247Z
mip1L/FHJfLVi4Rtx92lZg3Uk4HL/tLN3A6Ak7OtyIBjnRr0fDdEj0ECFWo/uR+ixWbxeOJ65s4g
W3Eyil6LP5avTH6H5cbMU5dmzN01Hys16KqukWbLavDP751T3lGgof8ifiIYumnmSyj3AhWwLkh4
IrdD6KBodOXMclwdQOeQB4hQFzgQciNXSbkPXKsLPJqG4IKtJpPoOwpKCJEY4Gw15fzIB34+mbAR
b3Lbqg65NZmwW43PHQhuvSR4sdoje9I15CD9ubAfp6VKdf4xPmJg4+x6Ng0Xl6GBXDlP68TmcpMX
KnUDC5iRxC/bH12ARidAE5DfkNI/GP3VsnWkgBqLs7isLrqF74dKiSrM7yf/Nafc5wEujdITIfzz
8FOt3F7+jSAzPlHmWuj5cKLN4iq8FAyZAgrsod1fif5rNxzxNAHR21ydywRoZ/sRUtAn0YZC6jcc
WRpfD9eDhGyUsKUvzEoDBcQPRm5/y/f8PAMX0tE7/pZIFFChH0aRoKnSfQrt0qGRPbY/zlnhPdRO
csMn/WQ+01SjXK/4S/H5YiWItdRuv1sIYh9LOJm9v+yRgeP7gWSjoauHsHX3hLfZHbqzMkn65+k8
DPJbCp50NEBM1Qi1lYn71cSkNriCMhgOQcoe4AszjyG5fFRNrDpK5GqcnGuGmDEcr1dQB7HNj5pc
TBu37vBAYFXGiHt8jHV7Ivnj5Mld1txh7y2w0KU78NUgk8ksmLW/k/nCSeX/eTOSAjlxnzi53Ln8
5iz+/43cZQ+39nEYLZQlC2YiqE21PSfGujpN2SnAlfYz+y5E/Vv4lsBCB6a01JpYNmgvazu2Sb4f
8j/UPnd1A6cEsB7hcC+l8zVoKOZd4MAHVjqMyjnmSbWKpopk9rdXaEONFeaySwDfh5xE0GrFKsEe
iH8cdCqW3C8VvTqdQVRfgw4lPMpH/Z+mCJjALxm8l3QyygQ3wUA2jXqAoRFIlf2nEEU0oaTYpi4G
fBF2e/F1mLRkGiOdwNy6CamqjVVFQ6v4tWCOM0NqZCQRacHPBSIZfDkz/O8JCyLjgnzEhNEM+ous
dGUjy1+CxcV/rIv1XUkNWj6/yiuDF7eimzfPk20TXb0NP1l10+HuUC3ZI/ezszy368vBdb30+PFR
QTcMEYUvekL5Fftp7mEVwTd9tpTr1zU7PSPn/kZoCFsO2Bsh0zBNVziBFiEGlzYSt5REGGM+KdWM
yGqb2Dm6+D+j9NDMlLIPVqZ1NXTa3xkRUK7QlYdacvF0deB4YMWueM+9ix4TsOgj+WFROelNfHx4
ZtTQhIzzJWaKgUA0OId4Kp6AjcPEq6dgSWlLerIlzN3YuoyWNumqxmN3l2es4eY/09lZTQ3DkxcK
SP4fMXu+vEau71lvc6lpWx9kmxQKq5EswpjkQS2htGz2x6znFUnLUUXMzoaInNxgdCfhX+MP6QF/
VK23IfBoxhDSDsWds8wuj83qic9dgRQhJLq1ZPhHZtI5w/H/z+p2SXJS4DbTgAq3HS5PKBvIsdzL
gJHv+BHLLC5DRCz9Bp5zF+nDJbpmkEk8q29uaaG2EW7D22MhY/XN2GI3fNUtACJTVxOE/w1Gcg+/
qSIj5f+GSFVbdpcq6QF36re1uPRv3nt8bZQoLr6kRb0krF20Ym9ezpdVgO5h90aEBNcLfQcN4M6r
+8Z3+06vGE8gqAyUw1TPBF2npp2PiZelsPC3KQB0l9VgL4HCGvS8zxiG9BxBQC5HVX8xBxX6IIlB
0i3lhWKqbXG4X9GuQvNH+Ho3CwkImZ3zPIzBOAMjKk3kcw53/9/rcpispvTo11Ur3+SBO5i/L/i9
N39AZ9y5EQgMGsuE1dliIVepW6bijdgg8E9IT1pPU9+P7Xl7lBi76XsnI+9J+LJIbfy7lr7UNAZZ
M0dOinzOYIq59zZzdHoUGiJCCGrCUWSdzRPA4CKORw8Ov6DTAo84ashVlbJjsnYie6U1Jpha/YI2
jE2FaPJVgVO+o3R5DRhEYZwTqS0ZIoLwIKQjE92e7dKx3bD/fX6o5n1IH65e1MENAxJdrZ8gh8R4
JxDH508w1uN++pdf8I9W1fTGbO2Vto3Dw3Skq60avIEADeERDM3UTNurPaeXn0ZB/2qhb+Agh9Sp
rVaOvP6l/MJT2P4ljUVbgbBMJNpLSoZq59eb+UmNLKzD2eXcn1fr6tZPjdB5WxPcaZ2Dtj5qD57O
sAxCL8qDavj6X8x+aTveLeJm970RUoLtumPzXcpcY6wkn7car9ARKDhCXH1fpWFoNS6BbAbHcKAy
yuKrE6AX4D3gR0sxkoTh/aFNjspFrCnqLt8JHnB+Aru3kIqVlEHahJ3TBm+FBI5XicBSBaMQkUae
PJuRUJSgFrnn4YIZ2SdrIIt7UvWF1k8XXzbObiUOq5IHj6fZ37ErHwdPEgTmR3BuCdRJHa1/AHeF
FmjnHyQG4imZeuVTwLufQyC/+TXyj+oF9OXjgcENl85ADYrYmecvdShOA97seR4iwFt1EZ5t/euJ
j72Ou3Sg9CF89Eke0wMkPYHrTiSUHBubeiNvB/8bZr9brf8X4YUBI7c76PJT5gFecUbZcBch/pbs
zCB8YlbUEdkj/IqLpckolIlIDH7iQvgX053USlBCr/8uxv5KSBm7Q7K77lLtcnU/YKb0nKhxclOP
dLwF2SxK4WQjv4CCMjfy2wC16MF208dXVktPuav2+3xnvsDVhz9e6HvA79xC0lQ9CJsl/OYtd/2O
o1o5Zfe1oBgknYacf9Uv0/+M0OwFoIb4WrgxEG520R0Q1mZ2AN5j6rPTeCI6i9tq/Vur90PkYxOm
srkN+nSjf0RHwOHoe5hIeXTfYRE96TuA7IdD9StaBi2Qw9vlbO+aB7z+/iomgUVyEnTQEpIsYAPr
Z+HSGZwP6AwE/F9YAE3YWutWsVenyvFQzpVfs7OG/4cj0rZzpBNw5hVgTqK/nI8bYU5VCJSUc4rc
zpbxrjzaetvP/dkimosfUKxnpGkZLvD9e3Dv9LzkJp45N4yEXeVDwHcOkIaWdgQfm1ATIGZQ63Wv
EY3/TWAoHhlzLTguiFKtikMHOosuF/X1MYKrnu62eEUvlAovaEuP06Sm2s41VjOl4b6JiuLwUUcb
7EduNbVJer0qY4Fac8VpqrAaslvYVHlw7esOvgBoBhdCo/rsdwipxoTVZ48r4IY1O/FrR9zPsbvh
xdDEkR2jG1ikMOdRN9RQpzq1TkpWCxU1zkhhSRmfDdoLHVTgMS7VwSfGTCtwwrNXl7Wa8RK4UqVC
NvElw06zdhKoSP87URjGCd2Xp6MdxidzlFwQnyLGwTwwfe5cS4IHVGLFKRLeLlN4oOJQ4vFjBgCS
g5RzMC35kXftYIm9BCYkhQuAaFGQpl1x79t98L7/+WsAIlZOBxMGqf6iL9zxIxylkwydZrJG+H2O
/1dvNPSneXDsfgR9sVUYYzxTxvjtoMTnUtZkgG7UloOGmyYKnu1RCcV5BGMgKP/9X7IPDSHZMxX8
193xbJRhWx+NzXUgVW8+tV0GswXsVUSvLiVHZ41Jesr3gJXfbcuX9NF7rEmJK/XYib+kIQjrwqnd
0aZsdEHHOMY2Q03xwU4hcgVt88SyCY6A//I/iDKgbhDL/zgrOy2yk/4ao5lTadjY2LVA8yb2GDhB
WPkXKoLEk4F5NDz9BiMr8aJLVvGEUpVA/K7WqwR4irnaM1F6fB1kBuRKXi6bP+OJjLZnjL7gWGyQ
ASyZ5K4VrLUeXM5A8GzBsnyo/d3HE3e0WRDg6wZUzRoTNRuyIdgFMKXiKmZv7WKEq8AfbcJ7rJeH
6MJDgh0ofAXg60owi94cAm9Wd4Xh7jj19kwXJLX06/6nXvn0P/uR/Sba9u1PApAIg7GaagKGbuZe
MD8x0gKHagXcVZ3hwEE/V/Q3AAMMVwZMsttaQGO/l8mgS5/T4IYbdB2tVDn1uJADc9Xf+pKQXcGE
NuzW20FL/R3mk61OmT8WFlhlaVVMyoIBfY+NfTUC6a1YohMRhc1fthLWz44e7XKMmnTsP4HNeG2e
362pUOdr4FxkomuvMal0lf4cNinxkZ5OfSyweo35lZd5bQySXcBA6NcxqAOEfR4xWti+4YZNPBUw
UdTOLql1GbmXC9769EY3svfEiNqawNbiKx2jtOA4DhEq3LqwiOP9e2jJvMEW1ipCQJ22a/UjIYH/
2gvt0XsXKEW+PyviSgtF097EidhCXhYg8vsRzshLr5fy+nocFZ69Xk5Y54peeNQCQ1+VM64BVhPJ
VLi6JS+3joD9kiln/PR26yvAuMNj7JERT0u0HkHgrfXrTt89ioyVHWQ6VGqjNcG3TvGEFFPX7es0
2X7NZ5vTWVt5lmABM5ppwSI5NFIgLN+aEwSgQ1zlvzCCnDGb6UI0j4Hc8avkO0revrrY5Ygc2BzU
yl1jLH7MGdrKyKgvlfi0EvEcZIg3K/JEGcgs0MO5rXkC9xD3OlNwPsExrPlPUvLFXgDR+yu2m24b
pX5bVftMZ1A4TY9ksthpsVJJus+0KgeCo2MfwUjH/hha7XGzhHncVYgblIDHHsbpvzVtv9JxsqUO
0YJoWEJpziJsUXr0P8fhWKWJTps8+o0paa/yglACwJCGDG+0WHyXdePBReT+NgJSI1DkxJ/z7yfH
NwUC+nfoI5wHxgsyZ+aWENfRNBMuP0/WOhsWpAdEenzEmP8lOXdlx04VSV2fHG3iMkZPegwB1YBJ
pUW+X6evKZKfGp7y11w0yPjEtcVULZkYJVT6DCiHsPPoO834eb1NAfpQOoRh0FsCgHZHxf4mXQK4
m4LSm7NaMtaQnkJDnMGTMr6QeBe/yXoxol0YaTX+TvlUNo8Q69he6VzvkjsH3eE5HpDcdZEcj9G7
Xox/tMzYFpeSAUr1oUxfWi+uRnB5NS6iGlV1gopXpQ2d4OVG9bWYwJwqEj7cOQs/GxyPiiZxgBR6
a2IkUyqAOWpVYMsNMohiMjKt3FkhWl58kG3ZKzorj71BFz4q/fa50oG7YNBjNUG1+LQwEY40Dh5z
CeX7cwrJ42we8e3wOOG1Z1rJG5W+fZkI74ZJChvR2pxELil2v5oVu+1wwz3+HZlD1mjAYgSMCy01
BY8T/uqfBCUh41gWzdivsWwFe8gQ2INNZ+4lTLJXdvn3I4itOAjqIH9nGkAk9yXYyEY+qsNPQxQj
C+RMZkr26ebQ4/5yqsMGiQseSkQb7rFlhqi0ODVIu9AQvFz+JwvqYQdi0/5QKMlFyl/nFbrqZwGg
zQF9WtVdIB6Y/rBQxxMuGWX/eXlYBKMgBPbViY4TQcGC1npDJ49BBvJHZnHYrEPQgNtlV9OJR+bf
i4MUG+EcCH+/Orl2r9zOkLHOEKk/544jlr/AcJSSzqU3tP9ZCDK8q0MzrUvm2nlcYghHyw+lIi3Y
1Rdt64IvUPG5WlXS2yOauknqCrMygty3Q4cOv9+W6q24tLqCWVAXhUvI5pruqNxRQTuowF3gMVoK
wHFG8LNhR5R/hfc3BOIeOshGbGCoUuj931Tk12nTATopg9UOX/WjUBNm3LcL8iWJEpEpyDyvWFnK
RCj+ed4D8mWrZqR/yM+2VwmJeeJYV0O2puCerLPOAZI/+k5JTAVQnq/7r1Yr/aFiR/4rWqgp5OmN
iVPaxcSEGHujJUnxqtdhxTWQWwxDkzaIcQT+nOT7HaKQesWPP3DXIVksVjsqnLSWkrGQh9d+F+Cf
feHERjl7DYDv3pf0V+2d04Feb8MQ5YqFLV053ZnKOPCIOstl8BCL3WBpqvyfI17SitwA5i10r5+y
dbQu3NuQCBv+IjNLX6tF5VkYBQ1MPbGMIOwtJUXC2dlG1ssWT88rIHI1QjEthtp7au/ENry2ifR7
PKvUPYO0aalp8S6rZDRpzOA+q5m2bxMe9Zij3Kv5bLVoZpTV0gzLqHf7TwlnBVBFPHJYZqwcXhSm
lvswdexzsf3c1fzMwOV0trbA7um+HpcXeD6BrLZ9N9PJ/B6z/QQpEWQXZgCXdJimClcmIgXIncSF
olAy0YB09oGytd55EQa/hOMJ+sUcUvmcRjaOgfbCj6/7rGKGYnrCYg60ikfrVgeiCbtWKarW4uKS
Qw7SUuBXBQs8cyGXuU7Y8r+YuQrC5ncZ6g3olRi/VDGODRueBQ0FSK+PKbPfqBpUr3bGVQYkfQIw
xJ4xwNE//u2JBNUD8/pIq3Ohg3KSloHQjjXHmBdsMHFyfbmlHq8o6JsOX6VFWnN9AOLoukFAD8KC
lhXNkqv+PjFxEUOOWUHbML0O7bmvfHGbQo45ikPCs05doUKcyA8EwklOB7UE6BgPwydhBmkLLidK
c5bnNrexnDoFkgfA5hvgImMxd1bx1zmsbt/Q/s1uG6D089exHInsbLLsKM6q6OU3cVIZcbaD6/I6
lGBLktF4FEkucsEBhhD8zQ/dHylCt13tFPDnddV1JFN266odrtpT9DJPQ0bI1aFyLYlhTFVBHSt0
3GJDZixxahLiLYUZwuCcnFqA6D8rBVbXjfDf3awVjtA/CVj2QOFmxsrB8J30RFfthon+uUn6WBeI
rRLXMOdR5Cr0U2skNaWg1PR+0OntQOOhiePvUq8X3TlW3vKDSKU9VYl06+9xu7mMDwdJR++0DsBd
R8IDls7hZARQJVokvbMOZGHUXm9RCuqENQC0AhHvlIWK0FQljvO94yNYGcn8ERw0wn5NqFZg/VRn
9aI9xucm/omkGfX66Y3XdEimaDug4GbSECPhqv0R7i7DWW1grj4E5VSzmNIIweolFxJn2BCAfO2Y
szfeNq4LgVjAogVwfh2kTzxroU8Rq27z9jcysMAEHzfNoUE3uKebGoT5I4Q0F2UnI5gGBQUongeH
fNssb9CwHw32hk/FZgjEd2ZmtKGRRhLRvYa2Ldwk1iQdCNbBgicRXRD/joA6TX61sJW6kA3gbsBz
BmFP1/fsB3KlkdSVP7JoHDzJIXm1P5rQQch47FrtldI28gXneY/e2IrhqbREo/grcjZnmcD2fand
plKQH1+oEErxOS7PiPjl1W+zXH6oN5nQ7MrjfwUlY4zzKndBVWw+wJ1Z7xpU76PWzLV8aukkzGxr
jiR4QCUQLgSGLuUVMYrz8wWVtq01u05V5uKFqt9JzYeRsCa42itQKkCGYkDNfM5VUUMKnx524jbu
Yjq0ae5Mu2vLPZp7/TjC+ox15llbnFoa1INsd6b1TCQ94RyvyxM5isv4EKAOs3tXCxnuWCbQkELY
us8VnC/R0+5gcy80L2jt7N8WqHkJzfEJ3J/xopFpciH0ZiBQiz5kTD3rq22C7TRisdAkjE1+ZvCB
sA46569oodmhqVbK9RxtmmZAphFiQcDm0vjgNaKun2PIHJiksbmTIuVIdjRa20l5PsGFDVV5Ydv3
Mik/FLLVYhteI2PZ1wjKEcLAwuIUAWIlGh7+dbZh0y2H3MiyQQMQ9cXrgJyRlwMYDMIq6ktX+o97
SEXN3omjm875Gyi3DlsgRWsR2IQx2d5w6Bof+6eTIC8xW+LgCsGmJ8OzDjeIFZkLrFYFq9nWVy2x
TedDQDwuw2ilLNns8Ntn8GXuVGpKukQYdFzShwx6Xs7PtnZRrx7XB4FuMo9kN8yI1+fpqaLUkyYG
Ken4DrJfzP5amNkTWODIKxnihdijkctSntbF9tA4V73Uqce2i59QaoJcQMsd6bbxdH/oSx65Cexo
15Phi8T842tuccjFNtQPP1l75ZBBJ23rnU8joswMwyPwmzu9z0444jFoBOERxUlLq0WtGUuajJJ3
+cw6BTrx1FO1NxPD/+qZxz7CUXwiGvHwcQf2XTzBrw0skeChqK+rk4Z9aw1BoxYtwXG8YbRRW1Bh
K1iSAfH/Jw++EW2aZULlVeFutn6slOXwQ6gvpsKv/adlJkmLOTFfTnPPt8AgosBvg3y3XPVA8i0i
Z/mWX61dcrilWYXopeYE8zjpJekqVsjryx4sRTCbSiPYd+9V18kcuzDC9GwPk5+idUABVeZ2kZYN
pg9Ji032ChzLZJ6Bz1TTqz8MfePuQHCd9I/8jWVHLFAiYiK+Ho9RMymY4lxKkh5Nh+vEv9jH8mKD
ZyZ2SVeWHNDqy0cWabuVF/munOp6+wm8hWmZR+flhP/XO7ESC2sBcTLW7g8Uo9GYJpR4eLnZPIJA
r2aDoCTP9QD8vOr467IU1/l2gDRgtrnIyaxcN04eZD5zuPdrjucHCaaSQqhZ7eohwqfVIiB2VBY8
mYPKxBhiCIxEQ3gw/GfhhNTvfcy6wcJyHcuSLm0lWji8wmp3ip6PqRT5EAexAWskkRhkxEeYdbsU
j3bPe6BsP1msBeF0qIc1Ct3ATNKxLqkC9OU+5GI/TUmy6XaIeYN7qateH9SR9WSfp8dxu4M9cwuA
UJSsp78knidnjAVOCDw3XFS5OkKDJBZf76CAoDBKkSRQ5ww8CJv6LAAxNFfVvQSrx6XbdDMcI1rL
4lyqk7fGrj3Dbti5ez1ph6VpcgGt64D5m6Ejrukibp1OQYJ920s+WYCgyUwe8fY0WjoN7gSzmgwP
wH84XUrA456dQKqSJbSZ3qhTtS9CMj6HhKgNmqvpSuJtNZTugS4Z0wULg6w4WpPMa9PLuJgPvcUy
T40Vm7c0827f+UhozcS5DYWhgJLEjL+76ZnBpNJCqSvojiWJJUadsKQK60KbbSwtUtCOIczmRw+X
hhGZxI8WWETIKMuL05ptyNBSuqKWZFxBYqVZEJXR6t5NqXl7XqKYcWrpQKVJAdiHbh25Kgkgi3Fd
iYob/3Unk3a3EwCUiEqtchPOh82EE/KXk4FxO3RiOzmlZ2VUGxkbfMtvo6zTEWVHXv782RP3Xtm7
d/sgVkCjmh3JqWI5xh4NqPgVUW5NVKCUX1C0zKuPSFSw2Vwy9IakusjIeWLNBUPVlH2u1McTsetN
YX6cFmd7NkOn4gRmMkxyi/wBkfLefSO2ysCK3aYo7kkFbWNl58YYHSTfa/DGOOTHS2EdU3sV5cJa
tUO1zurmmyk6BJNkmRq75aMJ390KreEpC/MmryX7PPjiI1GRMlmNm4Yg8DOIl0o2zLQdiUOuxnYe
mczIgDpg+fjE1PaCq4oaao0076DXl5Pf1qXDtb42AP7u3DkVfBp2Q0jP00UIGRfarVzM+P2r5EJ9
gBQENmd5Hxug0vKbRobN64FJOZ/i+AyKRzG24l0dcb80QZ4f4c24CnjGm7CcNyeLXeKHGq1fKlW/
Q9jOSeKHcx5vbxeTlvferwzxcNAQxd4by+8YBGAj3/4vkjq1FJIJy+B7yH6Pd02alDHQ3/G96EMF
XSQedNwWM1XFi9HP1wmVUtMvYcK8V/ysSY3SiofdIoS3Fk3738v2jnNoUTH24NIGxkHQ8Al47Ghg
0CHJws59RdYf5E66Aoh2eoPlOKQI1y8ibgvr7qbrrKvv9GnlGACXNJ1hBiDh+GW+rsjKu7VJCqEu
9ZP+0hhiUPcFFAQFGuscQ/qcE4xrO43HfwNGvcG4pReJid1wc695Zttj+E6/SpjE71FEZbwoUhr2
aIjleAk1MJBUWSmZKLc25mJ03Ihz4dBxLROANbghd+IWZ87l3GqjQ9kX8n/8JlHwg44DaaUHqu/i
KUfSPS4z9dbnuJ3VLqXzPwKmCdl7KG2mC3pPonoGkeH351Wtboi31SocZlrg1zHKBUHGznHLw0G8
XW0gbfMrqpXMPoK0A5jzR2E9ndNtXm7vpp8vLuWBOBPxqimpfgbJEuHURJsY3Hd+tXA5eel9VdAh
5p9HBQ0fSSSYHmKFdGdDNBtggg7Rx/cEJpLgUc1O2zH+4elPTH1eFE400sNw4XFZwxXV+oM2DdG7
9VLxaAcMLjRnEdtYMa4n9E48RTTsFAERmkQUVil4IagVSfaB/OdKb0se8wbuW3iNW+nzQcYmamtH
Xuhc++q0XSqtnFZemeF6XN7FFQeoj2aZGkLsbfOfLQHII1xCTzgGVXTcO6lh/uhXMkBXLtBULWN6
dB5NRyXUpmyNuCl0Pjbw2fIU1/fNx4EB2OcTFABeyDCNwdo30/Pp2Ef8PwUbjKI2XVRhpEm2ILT9
/kko2CTZNStpuiNJTu8LEDS7teO16z69UQQe8HlSXiLhnKLfAfhQZ9o1IczFxvcdziseDtZiTXGM
/rshnyaYghrZ6CKHyxp77XIvQacgXXx6kXgGH3PkHLvHmr+4T6/Fdb1MM/6zF05sL1fgyTtbHgyr
WgrgU3SRW6WnIL4fBUr7C1CaMHZux56p7xYMSuLSvX2oI0SaqQFbC6YIcGewnXbbDgvUfsgErpcO
wdvVhN5YHu2Y67G3MJ8KLSeXk5I9Ouqvr0j9p+YEdJBBAQfV/WLlc8l/qcxnTTk0aFGlcQ9ZVDDQ
9PLkDbO6GcXMZyb6Ck+FKhEvAfqiCu0CCrCtapHtKNwrzENEOYys4Y3s9ytWEbYDvKloizCYtF+d
rTWoD1EBwBRHSAvSTLC/W897ocJkZmfGZSwwGUW9HJ3VKQCc76gnALlPyaiSdq8MwOjcg7GBbfei
4oUWkdxdgdkQaFvtLFNe5oOXU5D63S3w7IUUmcRArLI68lZgzLuJnucK1I+ulJ2kmLdioH+UneOb
ghyc51nkCQv+6gKgYcWDa7JBN1Vg0c1SQSxEjzLXiNOpIYZL2I7Uz/y3iTpe1VMa0pDYAfc0NDNK
QKNbQ2Yl5kAn6n2tZgxoeuENx5wfDEXYz/wf555Z9yVCJ9L/Rofb3rYQ+sK3bW+atxyFiXaHZgrv
AxzGOZ5tE624A16a2b40hnWHm3TxbUlhdkqUpM5Jm4ImubSaKt46ISA21EQRWWtG8UCQOM9dJFyP
/WHAU8TCjSLYuPIY225UlsoI8ml+1+85jKTbuC7TpEklcOo5rEMNqxO8AqcSVskWvm+MRvrzy3Od
xXgeYuX+YkaSkFzRfDew8liMhXn4t9Sg8tFJPKjMSmanQp4pddL8JUPaMdcxX65O3JuSpwx8hc7N
Py65GL9yGAE3OKasfcv/Scv1O0FcsyE8lKaXO9uVCkvLg+95N2vhf2VG2hXF2Mq4hyYgsYS5CqyC
Qv3m33HjzdVYC1Uj4GW9prOdKVZfvAHURcWvJXwbb59Uq+qhidPtv1jU5B71JMlflI14njIH4Ekz
X8Ge5Q7UXc+wEMpCgs5AxXsJYYYExV/PAjb02da5MDXmdvHlVluLbTf/YV5ZTsIxgffOQL89j7Jr
+Yw2AsJZfO4xq/Cl3NaS/yhmFVXfMk1Sf9i3oIs679bxvNF9E+4iO3MGDC/6ytSySRb6DHvyPEP4
d0iyCZ8UYB6bb8NnsCo5SV4IHUtwypQEyHojpy97bRv7ZUvv+TuaJkdtFntdDv6YD7eKzQRyRhPr
UzMBbJkIR2chylsVuPlLgstxa51Hh8aQkZPpAjPEV5jryQm2dm5R7CwaDdReRuxDey4pNdzPE4yD
4V6MMZ14WAlcxR6kOoFTTeqEObNy+D+rnVbZRpnf9l+zs4/FCxX1U2OJGkOGrhN5QSdrf9YeMHBe
61NGu/acL3WbypQ12GwxngnndYuEmDDUfVAEWCjo1NTqvVbpHekfEeV7wZ3jD9EAmAZQvXwclx7Z
zKw8eAYFlE2+OKAh8syj0tCLKBLn+49BH7w8f01XYNQeCH+Ton12JyzCw+jvuxHfsuRl2AiMszhu
FBVL9fR4PR6JaFNaYqjwlRwIZvJj0uLqnBfe85kc9R+SrCJ2CNP64nTiRBWq7Y1tmDE9kPIpQX1f
3kiA9NRSg89I1E1VQoaMD6Gx7i/OFfEqW1HvrG3v6JTfEWVrsOitcCgwsKSHS3qZEgG9+FbQ9+ZI
fP+Qz1Eo2xnu+RBYpGfeGsqyjd4MG5rzBSqEeiOFdDbprkK6Dv53GZj1hrRXjRZrExLogpDGWu6y
zVZFk5qiEM85YiTfj/7+oGJzr4gX7vKvOZQ8MqufxP8deLfI8qHXhaLBPjOoEl2PkQlTfP9VbmPY
NuWzISA1NvlzPQF+0K6QjeI4kCGlh6bItn/Y7x6HKHw2LzGEZ80IKjwFanBy7AtZ9qr6e7XiwX9f
omvwKAHgaaxHVDOUr2obZsprzj1/qTkHBIe33fuCOeTdM08vEu77nwZcYj8coV+sAB9VrrLU+4rt
9QU9aNFZ6w6sq92i9PIQa2Rd2rJpe55BoPS/+jYRLNA2NIShtdfabcO4lL42ncCOlDXi+IColwyo
nC9coO8G+8s+D66mRWi3wWT/LcFDQGHPF278eiYDTB71Pa6FZy2l2DrFqKl4yB908c5oClwQvxdi
PO4RNYCI0unOV3wf24WyEE70/WtWd02ce6+1X3UEDKQ7d+TLJKr/5VgT0O9wLfVzaNLECP/QTHdP
+dcmhZApF30gm1FYNmVz553+THOOD2cnWJPRGpn3BHH203mXmZPMb8k0wejDKrfB6KfD7M5YJqgv
LcGaveMh7NxyHNZGip4M92P+JpIH3bQSf1aqcsnUcTiJ372GMDLuQbFJRkkIfsccH5dn8x0njR4j
+L6+wo9UlrTCyadEwUhCNeLvlnk0a4Rh5IJ/O24nBPnhMj77fySKi12tJa+/fcrRZsaUPxq2jID0
ds+nPhltUv/RMG7yPDdpyetfT1r66WLAAlyUUfX/yyLVXA/ECzI6O6i6QHsMcXgwFZENWN5Nd9DR
lwIUu976tIEKWJyTzXMpwOffHe3c6B7dfjfCtcOBAsT2Sk0sPO9RaSBtX5OTnoNzlYEEo+ae5a5n
WxM/iMy87JpE1WdOWtoTtanvcKBJN4tfnghKqml61kcy/aidPVJXOY8vY6e5fuoyJrtlEWF2S8ti
i9B+vOKgm/y5UmqsM0IBjxKpVg8YJF8Wkgqz+3GtflkmnC1shEjNgNPGwCCioAhEnamxP90+BQMe
n4xG42N37Av2eZfKxpwc90KXKPFBiUNl6bqW4pZ1INYNtpYRWd+0/m1fnqhFYFbnjA9CxqG1VDrv
1R2r0V1L/BQwkDW2uHL4EPG1rM57LKyU5tpaLKjVB/DBIDm1blX6umNYfs8qb8eaZCIlkBV1GrkX
BeSg5HMR8HQo+5pPkAcFQ243QxcOjWfDxfJ3FupPIB0R1yMaD9tqtzsij3LFfxl8TPsC10cuzye7
Y9sSrNXa5qZ9xTERhmZDmAsdRgMpFQowmDsAvjnmhOC4QOG5AKRztzt0fV2q4RdJYK2lybG7l3yw
yrgJDCKLMYAyKx04y2quzpKiDxfiJDKNa6RgLZvP+doqyVM3Dt+YdnXsS4L8yJ4YOcyqQYwd9Rvh
O+XCB5lU4j/Mc5QaenyAAs6E1wUAQdsda5ZD6B9vOUjIJhWwCiV6n2QBelzHCkuUWnGGwZnVTCbG
vIKcqjmI8YLjaroxG3JBlUPtA2+8Ate8UFM/6GuDEZAQ9AGsDWrTpc/xRKI+4x7opsEI+0kVnirP
bDKvBHZ9CZ5vmB7RkAofcYoPDTn/ZH8+TIv82Mx3y18gaYIWWYdHmHS9GDzhfu4ChOI7QgGjZDjk
BNubz/9Eue4AAjs7HnEkkplWClKKgQxuD2chWCRrSf/BKumCm5hbul/ZiKzH6I/HHEmz8iWbfUc0
+8mg/FlxpeWaBn3khr9zy24BhVuznZAtLZ8FwxedFBlDLPq2/Ld2HiPwLAKqb4lowuBtyNMxztwf
jAl7AYFKguwmtsFXYHGJimQYe3HQawLkvqLOPoHekRjHmShxLpS7MmV+OT8zZkFEiOGby0EEaik4
edyKCuToZjfB5CzO0N2k8tT01lvI8KwccK9NFVHARomB4pticZcvGmxPciIAz6KTLvPIruRw+m9p
Iy8+qyCQ/6swJx16SLZ1YqG43VvSVWHgab05BZcXKj5ltXhsRM0LzihH7CqgzED46qZCzaEoLFnp
+jeNbLvnjxsZV53uY8cygMCeoUIRPvar5lsviAYB1B6aGBYcaIaN6rPQhMJOuNFRW54Phldr9k7s
hpJmK+plRAripBK+9u/PWs8V+mTG6VdnkQJ0W5URmAuOt+2g6Y4Qs3+aEkkE4wzeaOZ2t8mpkOjL
tz+jbSkEO913otVjeTjjvaUJ4NJdxTFq8JvrEa5OC5FhQopI4TO7sNf2e6f0jE8Qon/ssjs8jp/i
eTJtONorYegTteiJSqqMvWDJdobHLbDuJCHVk+C/dGIvE5kpbDlNEcUYst4USSpZC3eYm/36Y8SB
DzAP7Tb4lJpHBymbevfh8IjRh4Ac2O3kXjEGrwh7cjJvyhwv6f+w42Cv5FGv9qt4pcrh995qfLOF
mRPBx6DPBZvODZDXMs/SLZ60SP3WLy6jnuwhzo7L3yMPeIuJ7byuOezdY7oIDduvSlr0ZJCQ30Ei
qzdCSg4MtkMENbiJAZmvCLF1PdG5Pu/rc39szOtxUf64TFDD8VfPVylIosmylBFW9fvV8JZy2KTG
xewVRn58+msMd8e8HVHTtjXuugDyz/kp0vEuA5u5QEFUwkMc1HFHzwE1F+9kLjoL+cngPInfs4/r
n4VfNMtl5tw9fNxxu0fSKbA5cVgmvCbexCqHn54cGs6MkL/vARJl0d6zXttlLgipZRXZvn+430BP
JZrn64MYhcIvtZ049tP32IgUxSO8ZpfQ8lhnys3AjL6W53zp2TpIPIp9uR9Sl4lAgS41KljwgCuD
Ow/Yrtr/bnjdYtV+ZGoNf67+lsp4geEY1Rv7hQxr/Devi1EoPF4JvHJvStID5SX/ms3djYvxP3jY
aYIrJ/ExkjS3mT7et4Z3yv5jEU8I9oG31geobIHBwvXdrehAwrYloxduekCOe3ZkickEW2kRFQFI
p9vxf0fosHjeSbEk1tLiy5WnmZIPywEk70QK/vvR2S6umI7WM10QM2RwIx8lq6JxDnXYjQRU84bP
GSQw4CbyHhGE5w3SWBZCnMdpgTccy+Dv3DeXzHU3DSdbAW58Rv4T4PVNNR0Q9Pzl/0FQC4ifG1gr
zC1hqonaQYGMbvumDGXazFVCavvmJ6W4eDwfs5tOt/2mz+Pp71HoTFTCEj1C9Lc+eUFuSvez0Glc
eTAAROokZT/6sr5q7f6FyKQEjXkzqcCFdzs+wbgqyqDwIOPuQf9lOO5ygu14zBLG252rGcnpMEUy
gy+s/fDnikxytuHIvWkZ8Lq1EllzxCmB6T8U36uWim2GA+++dB9jIsTvcyEPM4nGh62cu2zj11eS
GKHPzR9C3JnYEU3dfctoNFdAOUNfeVesuc0naqtJxg+3mIqX9W9uaDaL2pSocZG+7PQKqXW6jfv9
XVTZAh9dU+veHwaKaqIhXgg2dLp9kXLPrc3Fpb7UDPoj6ySB6HgG0uPVXeZD97Xc3S0/iaD0T4w6
ueWycy84nCQqPelgvxQxCGsOORpKlh0Cmn3JTTGTqNKEFRtRLr062bWt1rU63mDQj66X/fsXjvXu
wmxr/zABLeZMAzE/rSY/G6uoJwRJ+1G2ymtVgieLvdUmvpEtzCLbMzPKsMiRkE798k3uDUj1h09h
ifhRWLWMyCG36Jhh/0kpz1XnBXNH5T+VPW6zKQeR3BLqf+2WLD+FAAPHwM7Yud+ymG6L8BugkWCa
N4yM7i4ie81suMl9Q6WQq3fDkZcevnqrav02GnqM1trcIwrsVkDe/xrSCqPyDKjfbPK7J1Zje63N
bfnYsqsT1BFZ4IdBsDLpd9UKgnOfzf3rwuL42zc2f3Ri0ZRU0eQJF+/CTDN7n1xtRlRYXB/8WpnO
V0QrGyFpeA1D+1Gx0uMEbpvMAnSSH6z3z9PNuW+gjWYjuPVc3gJdgk8UzkReI6MbPADMeJgGHIT7
e+USp7vYcofIygyQP9bkaFMnWdsddpJZYoK4C2tLJb7eb6uJsjgipQYGdMOywaTj4a8aoDYdVnVY
p6wxpcMHKPlKuiTadh/iq0kbMp+rarEjdPrJ3Ld9n2b1TYh4jOPmn0ETwAtE9WNR7iownxHpiqGO
HNc5H5RtAlsuKfhw0Av0zpt9BQHI+Q/0ernL4whYatRUj1QLvDavM94QDCaA0YR7VoaUfj0T+EE+
Bvf5eYNp7fwd2hQ8f/o8/COaVb9FJqPAbJSfqrBgRRsJqoEabSUwtayzRuhhQkDwmSVO0yqZHxBi
R/QUh2xSmAVAT7CIF1IazXy2Nxkdx6kFTpF7dxFgpVMaaSAgJ2lPeqV9jPYVjQUHbqVSr0njhGoD
NwOfZI9OcxVVYhrMT8s120jLaqhwyhV4WX1UbXwKq0E+jqCBDdq7m5nSV3vZyDeTmc0EVFBauWlz
zz9NuO8zPGUQizmcOo6G4vOL1h4be5ZLVn6F5TOJHMxEv1szGhdrkaxA3Px/DkHszrf8YNugL5AO
w99EeibrzP8v1bF+FFrTZwOY4vrdIV6mzI2VQ1eWzUma7HiYqIYGahfI9z0J/vZYk5oQcXp7rfnX
kSAteR1Ut+2lZJBtOuIoM7v4aGMvopSxc5WodjMfn9vKSzXyptwyEfc2o2qD8/XolXKpQzMAz6wz
QKmGhJXGW5u+ToxbCTFS5xk/qw9ySX3R24IY3d3HEDeoQfyKEvtLaYamP0vym6gl6fYt8DD/jecG
s3VfTBmVc6xeApLYkUdID055yLISOs5wH8OkDXaLpbozJiC0pwzA5mBoo3PKHHCqYEGTo52fzU2G
wp+4cBwhYFtIciXAAVf/eYDioCURTb9JaW3AEX8mFI4DP7bxRexeOuH7b1h/V4VOfD8CJ/hH/BsH
j63cBI5UmhN2M6KbxfljtIfvaUVHBEA+Y4jRka9uGTPLo54AWcIcfws41Hq8mUlTz+T20V/hZfUx
syt9wxLJZNox6g4zEzsLPG6ZWJSmWlxBM8Fp+HVOHqnUzpuZaOha71FGuJOKG400Po2bBP6WqvPS
ZJitxQ4zDgvBiem8/I4oc+y9s6boe4Xn6I5RfDwGg+hU6rqqWYQr4DVBXk27XNuaKuzcbqMTPGpi
ihztVaEKIOTs/21VW3MklfJPMenWdCc/zX3AI/h6nHt7lV9MnPi8j6btOevT7CX9NDg4C5J6FJHG
CkZV69Vw4IiKPh+YbWbTddIe7nuX9mFKt+ax4l9u1LnIfHVuTzmbLlgQmYVTqws6QhAHr6BEyApA
ZgdFeRVmaQJI4xuCjvA0xzbdd30W5Nfn/6VNls7aCbwJ9voMx3rvqEvWcqJhjd5ofALIuuvyYYQS
uLm/kb3hRt/XhgGjMf3xwuICaKzUbWh2rs1SanT9wpum/TVFkD4iRotlW35V49nJ4aFHWivBEtqf
Y8luP/9kCXVu7C1+oWwM0pP9X/k5aa5Y2D/YLK+K/K9wy3ekn5L9WiQy2k3Wo27BLuckLEW02qWL
Qx/Y8Wj/nJ9CjIwnexkmWLHQajD+55IOD9bFFQ1VTmgHWyrDwkZ9GAb0Hy0R0mZJg1hvuGWh8dqy
3ScFpXwLdo8WCzwnPCng/+0BQbcKHo911cuw1b9TMrz1AIYtRzpNj6XSqTvthFkGfDYBinaS4u+p
hqLWEpx1ERn3Uitr/Q7KHld3uKPBI/+Xsidey1taUcTFuBj6QyR4GF8aegTnCwBk2mmEov+Sc1yv
lOINPDpqVuimcyg2v2bDw0v8eokpeP/Z/X2kOoJGZZT3pYnGOVQIBcNGPjM/O0z0630IB2EWaMs1
o9emmTD8CIeRV5dAStG8jjBFhONc4LpqP8Xof2pX6M5e1eTgllFDrI9oeC/Roc6sTrT0Ep/EIG1i
87PFez6u1EvHssZUkLPNz5IPpj+0RwPGLMYudHVEMZywBEFrakAZbBIkLwsJ9X0VndcbGo/q0fi+
WId98Bw5i6yCcNVLk9qyddPUerPTA3No/rf/vtEfPtUI1r1wY4g0D3d/bJij24gmnEeMl0b56fHl
aOhfr3UHZbA9gzGNKAR+ogn54ExMDPjY+a/6XxIXkENULNac9JfW4Hw/9jUH0i7W0HaN98LIfZKs
ip3ZW6Ujv1N04FOSlM+jtVCnEm4qekXF3XZKD2PDyB/VDxK8dSTSSlmsYUTnHlRNwp0UcRlWRLmg
/6d1Dfkmipr9BLK2S2IkTNxlRHxjqF8qGTIxQRNnQbZ6+LkGy4pAcA3TceijvB5TXx+25oPxzpVe
NmYznH561aDmEyTB/625O6CqYFTKE2MtzsAZNlKLtUexE+S3fFYiLj2rVyA4WR7fBli47SRLccvM
rH4XH1xdPDELX8WA5iDu5oJaqE42blm4O8l62T4lWgvYM2x/1KynwVv0XD3ptKbCsH7IabS3rro0
fWkG8YcVbHREnJLjgynnxVOFtddj7eckYo7V8nYIOYlpqC0TL6/ntSfp4hPZHeInjMsBneqdzYRP
+J48wHAUBnPIfEDAzExJLqw+pBo606cEa3NKmCYC5G9BQN6FCkdaGDdJsim89rga3a/lAIRe47++
VEBxPCP6fquxysxz4Zzt26I0Wdf5TwqrBqwVxlEsl7bbqWtFZCos1xkulB4o+4TA0obxpWp7cWfs
fFgWpkBFPJlSdPvOCDNIwYU/S0waeeVxOgEBIoPpCkmKt8we+XAUaahjLFa/w1ZZh0xZI3e4zlnf
2fIXLSe8saw1oCTs1fDiui6ZKQHkcYNhmVyS81KY/uKVCu01LRepnAGDqRarX97OMwN/t3jHNHro
tEmiqkj5Jehv7fXGGAp+QvYimuZOsHIVI8sdck+NQL/zuhCq4CfFqsRsdK+hfR/URxZzhON95Aca
f3a+DJU7nj1JlIytJjZLo/DWNLiqHuvQ0fStLxea0YXz+1ddKe3VRckXoB4KzucuDLXIqKWhqema
f/mw32vGzcsoE8GPv4Si2V92i+hm62/wCXYo3bhsOQuFDSo9p8+2hkdMI3PeH5N4vZqQsAHYXa5o
RETn00dSi1k3L4qcEAd5mkrze2+tOa2YtGcjRXlFYuWTDgm2AuvK78d+jGE95sh3scKo23bMnJFj
xOhw4oEd1taQOxpH8xaunnbetlIkdSBAGYcF9XvGtU377JwrQR31I7njmp815515mT5Tmq92aKpC
5p3onkPdwvh5/AKug1rDEMVd/0SkYjOB3bZGvp4OEU3xaIrEDfEcWeHTEDEOuR1bZuG943l7K5Xj
DD9mIqODzmuvCxsTpRuCsfeSilzj4dXrq76WYzTepPGHGLqaDl1Fq7XDtgs+ftaH0VMI83xuI5LY
unqVJY/LT/cWyNf4XUKGkLgQs++nmh3eE1XG4+jOLrGhjzjiJtdUHdAXd8MgTtNqW4voKKdNpZL0
18uNJX1G13BPhIBnsW/47OCRdJR/fjCdYS0uG1h5V2OlpMPa+oT9u/MHdr+f1pHbaS9/sLVnORJw
3HSQtre1lMuJu6pgj5LWgAz6TpT+TBXOLUU9ATd9KuPZki98LWuT4NDfz4gBuwP9w9AMVs3sqeRy
x3WnGI80C75cnYr1rIQL5r4ZCqEZKU7IkTxugPkkdIV2xqA3Bie9AZlxHJaFkjI5wNiNUxckQHnA
8WV4oC+bMK8vIL9jqJjEXPAnntNNGeMznArsiZ5s89jsQDV12Xjqpt7b6s1pRblhhBrl0gTNxslp
MnrrfV5QwJeCO/nhUgvzkTJ6FYv1t2VlAthUWqvgOWNByVkJ5t4mSuIrw2nrMQLyhBHQksvKzyfU
86l6ObAzuRq2vLi8NRmvK4ckMeuUMOiQYAPMj192Haxu6v1Mn5i92k57O/Tb4CpiETwNvOYGAPkR
E8tKSZr65U6oT7k+xeaKOaUGEFi481p7ZNoKmwfs5JOLBBn30kiwET4KY3dlTiXPEF0l2PsSsfLb
HhKzOAIJ3N4kH4e9poeEvAvyahtQl15j0/zNUYuZigE4btQfGYxzuakjxgsM+sZblV97xyjqdVRP
Rq57p3mKnKvy15RLTXrNCc3yE5sETH8OTRVru7d5PHxHHnhR0oK4QShEZF9t+Dxe1ZWDRoWGNzRq
pX8ChuZ4RwbQ/OC9GXAx2qPqyHQ+Pz3grA9BhigwqxRChVJ85gDANGSOednm/2guBTXb2kJdlqBm
yDkfSWR/Wti8lHTj1c7kQBrmMT29V8vaMtoJiwv+qXyvNCDqwXP8OhYzyVMuHKiR61DaIVG3a3/8
ZKLaaZGqKTdfZ9BuxuZB+hKK08weJsGE4LiQsOcKllXggqdFBjjZRej9FtnwlkdTjtI8Wq0EBxdl
FK+kGA7zmILH3ULJgNcGt/S+/qyKmwZxg1o4G9O8J3aP9sLSgRSAtjoWdsFmx2cEv602tLqySXSz
Fwmxa8aSKkf9mEGNuDIe4Gwb+s4ogWd3i+mEeagznX1wJUq+XcZzsMDct5R7dTkoz8z8dwbZe/x0
xRswjoDJGHtAy+99uI9d/Mh6YMmLwg378lCi6UI8HsJWjkk8P5O+h3mq4bJG5VogqQXOqaMco/SL
SDybQlmFQlLGEAwc+baYxF49ehWtT2y06td3xx6wrSJ53KbyvuP3iVVMGK4zVaHLTTUyZuF2QSx0
RwYtKY9zx/yTh0vLAWP/I81QxSQnZtKHTwonFnvPWJr5f45kOy7g2CF6hveaFz48RDfvTdyEWww3
DOe9MVcy7L4NEj5lldh3qtHQIw+psiYZUk+fUowz7RQLj/0vx49J5xivVa6upl05SwvIF/FdRe3f
fiUVsYz64gDI5aNzyOaln6tMmSe/vCfF/1INhOKmGJnQ+SpkaM4AUlj0l9UlqzVxB63/AYCVeH17
x0tOKQkYWmgpqqUQTedgvuBUslZBB+ybMI7v9R6ZjIiurnyxQu8tTyTImru3QFGMwaSKB7c5WxTN
sXhGmbGT6IT0ZNhcVqsNvOASEPQ6HOleTQvWOwy2kdU9WSbKNgm9UJv1mr7stzQ8tnYGGAE8puY/
fApPnGilW+Bb4YAOs4bs4eZGAJAQ2ko6YTTF5eEXD0VF0ZwZC28fQQ1pVpfJknCyLluKEHj6jga7
PufX7ihdugqKsbcYCID7eN626mBuccIuGJxZsf73qbNXpxppY2GzaAULTm638oSieVuCDYB2Qcol
67TcY+4+pU89TFbVXDB2QGCyrcoU1QeGm2+jx1EMfN/9FXt/YQHuzHuFDMy6rtNY9k26K6Ehscbr
5mWDRJ6JnQr+OV6/5hAzyopeMraxvK5ejufTyrgslUyjkt2mtJpZGHQdlR2gs8KRhd47WlL6gff8
sG/ydoFyy8pXEfrZv0Gf1Gq0LZUYqyh3FslAXoBQyXSGut0VlIpt/hgbV5s0BBwyKW/QpvJR275U
mzpBxR7NqIor7M582vL6JXEPbfhrryJitXAmg8T/KuRTYkf5lpo5LkzUxKBMJgTGaPeU3IfNnev5
bgZzVIlWEVJUHeNFeiCt0mKrfpCEEXQmf/9qer8m5wQBSBIy2UZX+aB8TFT044gmhC+1i6KYZKG2
7v2visVSXy3biNV6Sw0xt2NL8V++8jeb4957Lxk2wby0agNxkwlwno3eMfCCjC/pN4C0XPtwFBeE
XDhsPZ2UfP0aR+u9x97f6Zx+culqRMSTkL1E47T1vXccx4FBh1vQvTYvufU8brmcNo3syeKGTyDm
lUW530fpBzWE82OtiUphWVo6KfOUFXhNWGsJp0j4djBtujf272YZGxIHia+EKdyh4sZQ0vT2Y3Jk
EjwjVFWOIdYiSYL36r6Bnau2HIJ1OZ6AK4FK0XB3tf1LYIet8HG6ZgPZgSjH9Av6ZJiMik7Pe/j5
4DWTvdwoQEmKW8VnM8PXnJwPhS0qfKzme/FBk21HLoI1lYQ2qusuYxbkplUZhSd77f3X/wfsbtr+
xqqXk27tpG1ilezV2QGz4BoT7+89yAvQalRy3sGZxjCeoG78Yr3Zh9NaqLM4IehskdeY97JaleRO
xBraW26vluuAl8OIvq4gjeGWrtkcb6SqlPch8PMPmIj+//AjELzAcrLXUoqXHNsYtIgFDu0k6564
AI4iA6lJv8I4RMiymSpA6xIXDxC9h7Zb8CIpRsAuF+6xWS4RnN4QDuuhwYe2eQMQWrO+YMQx7uKv
/4bjHeTuTuEjw+WlVTsQm2BTVxmEDmcFFTKMMhPgvL3svinrd5EcoWJJ5ekSBKeFVG1+sIZAjjsf
oav6VR7qCzrQGVcrV5+9PxA4eokwXOevQJeEGYATvz2IBEIEkkzgXBnoz/PAANtWUDZ/Tf3qZ8oc
T6ykZGW7IoFa/oaFE+9yQJBti/okv75yYYrSM6iJt9Hixbswv1UqjQi1IWwE0XgqxyAKAofxr50C
to5yncyLUcP6NGv+DkAaGmZ3vk/SpttvnM/3PmHafp/rXEWuJUksXfnvRe13lD1HQYDUFYsi1iNN
MZbjVX1k5hJy/rsB+V9EHXCJD3MkF91WXsFNk15ilpd3tLFAsJDNNwzgdIe0xUJ8hF8f0INHBGW+
7kNccA4WPhH0rgdDwOvYae71tYk3gAEVxrIYKajY568Zgw8nJwkHhCjN9LMvk+K+Y6Sk4znUFF8J
h0JCScNsPUFAbxRXZuGkQqM4M6hy0IvTFvQzTozIrzGQRzBef8GP0hA4ojVhQb8mzC+x+y4dlGKI
ysywYQhhXHdQxc6oU3ISsA3LWgyFnsVnqUHyNnHlcWNmiT4LQh189XY0hVDhVXxmwKPDvmpNaBd7
imEWhP4Pw/VvYQdlzvEB+kg+pQKHP2j/VTC3oQtxIYGnKu26sgedWX/LpvNc1WO4bJp+HLSoOKxq
EFHmrQ8HILpxWuJeY3O4/KY8NYyhd+8fxuB0j1TxlcmQRypeLxHtJQH7BpBZ4Gg+PMOGVBNtgLPd
dK26dG10E+b2jrjGK6QbUOdO95EGO+gZkARIGiLmkwdW/57UY6JGWgvNtTPWbcEh9cUVhhXV+P3L
GsGsWrLT5kYNS906zgc/uE+bIUDqbewKrr+adNAUpeYn1dHENk7FAfl7EtHW6/WTl8k+NTnHmgy7
RkSoI3Yfhpilm0bdIsW0VwjqOBEMIscra0A2teNXS9SkhMsiEOIF/ULgJlC7KZ6vHPnp3YhqAndr
AGyTh4duhT2UlTZc3pBOwEUuaB1wdml/53Qix03YknC4KSzFY/t6TrN1MENvidueUWPLY4sjnFOe
/f23rfzxU+GBDzQiG3xUOV12S4VdxGiSMSn7Ul8bvGEEgNGh6cjSZOgztfQYsMvlgkAWDbYK39dH
SsgHnbIy1MWgG0JJWeWopgAw09Q/6l+LLEQaDvYiZkyuJ3TWwc9XJTvBeZw6IGbhFXSFdVfj5FZx
nFYfi2TNg17xovVo7HbWVxPR9CpROd2rxZ0jj+f8ByNKO6Z3XI6rtggiRxUihKah1l5dsbiAl+LX
QYE3P7JkK3OL3Tv40j4Tyj+5j2AlksN86siR2i1UjywElMJ0Xny+qkKvlfkikfsSJczjXcC/fKxg
9PY4cnYvWnOoFCsGUJHDKkJlLqd1uoZAtLgy5jhLhJaqPiixv3hruA61+dB9bGZ7vOafYI0VeiMh
znO4dpTsy1vNqHvedt469O0nEcU1AO/3Q/S6KvGPSv5CALsQ8cqthOsopXnX63aXlc6ytBfrZLIs
e65kLES3rRD4CN4y69XrV84bK0YVWzuh6JkYzg14BIO+gTKqQKyCBJVf2qcc9pgpx8XQ+txMSXPv
GWadT2DKvkWIUqwYS25ngmTsZJTNe4ZRQ9e5iCflOejL/532lan8dqHEGW54tulIIzxrPZgqLVHK
F9r4Yw2/a6vq5hUwf+QvBjgRavrpYHO/uirGayE4muYBh/Czg/CsYVuBlyir5TSIizUw8Ji+pzZk
f58oRQOTEsBO/nc6Bp5CipxYBL9Gvn64r3bbSS6VUjPrcatRRto5roZ14mGokYQUb47fvGj5aduE
QpnUp2bOiCv9h4Sp3ThRdrakc0gajYdaHVQtLpf242XeSpc4tnNIWz0eGT47518hEHsdwAyh2fg2
0C592oAhfWKvMkzlQ1naKfM5pC+t9PgoW9QUbqJTRDEp0c5u3AC9M2TfDRSSnObZKkclmVQt4Reb
2sML/aw8L5mPMyYUpU4VlZ2GvR80iNYCTTTcokY+jQFRW4s11pAnrBldN6BjGVM+V652qOpP3VGY
lEHaOpEtJok6s899gxL8jiOJl+ijaUBcRTiGluln6KzT6THrwV3WrAgh3bO9SNp4bO+Qd7TD4KVm
C1kxhJyxsyg5atOU4mmyeOzdKOtwVG2r5diUYj7jYOS6ZwWrTT8OqCjCJFRBKNzw2WZTPem3T0cp
1pXdtDK3efSzwx9w+5Q0U4Ltmq6l5J+OfboWaWCExWoRbulJvuy5bLP02IZzEWFdoztXnl2sXGl1
xo03faFVQmnOyH9hqDm9SlIxoQCtZ52/NfyS7MmLBV7vXI2OJtmM3UvoTzmTxYoenc2r+N8atQQg
GOQwz29Me9IJYJeMWNFiK/rph/lE36G+WF9xMpZyJlIOwGvmRmC7qUXN/Z1cTJPA2VNDmKxDlXXF
3c3QURgXfjuW2hUKWng5kOHszvX5GzyKmvRhD3MwQfvnr5Hfz50TaYDM3mH836PVaoDNDDoJFbnC
FvOXkKr3iZj/7jYfPseBUoHPSDcN0pd+qk74GcHZQtxYhf97qMUfG49gzuIUIMN4YPvwmcSQDXqo
CxUG84k1PPMlqEiWP/tYP+wMY/LdLaCGeuiWPbvu83BKp92o2ddg/5xQuM6gbd0L8lAPsfL18fmp
6se8wuIa/qGHfKkbP8PhpynAYOrJsqhf7Z5h08TYqg+IXdcRdiY7A4A6JXpyDY6jWYJjCkXiCazI
irKhdYaXW9XgZglDAFcJMf0aTXeFlUw+Rekhpoc/PnSrEs6rQwR+NWu4iPODQJSTnxNaAW2Q1vTY
8U0+fHVxlmVxUYT5IZP2BepLFXIHt+UmF4VNjVjnWj2Uv332EKV6UtoNEIbANc+sTMoIuwIr8Evp
iMjrHNCwrWlzpEm/Fkn9rGGuljtjlj06Uh9uyhavdLrXG3g4cwLqMHh/hEj/2oEvNK/x3okH4MBi
PWs4x0j7ioee0hXzadx45f5ik/1WF+6iwBQIGldo742i/ucNhih+LRjDQ643UkLBh6ZvEbKDn5Sm
xyOtHsQ7h2bJhVCcU+UvMAVbRc40VQHFtuXd4ibRcI9ozDvrTfoJe+gdkTGUoQTaiMqr/Gt0pnFn
o9o26CEHTHxfHZlejPaKJjNax3zfnloN9v3fFIXr6YLsXlexBc9/lADXS5ESRfnv2wgPKNAjs+yT
cIhoxvZ/pHZOORmGarw/FMXO/PMdpxLzxt0ScZ8wlv6iKbl90SndoEWvcOGwY+BZB/DyosYFeD2v
HEmxAec3MmvKvotdbvjJSDGzSzIGNYixbWnx8TB92gSm8khdOr7wq0Qn9tuzYRgwtgwRRkSigJqE
j0mY/gsKmy2anSFvV1CpS3qykIXmCtzeGRgUS0MWR9G3ARB23Pjksjsa8oEAe07sGz1PlML8GV7V
q3Z6exlc7erBlaY7bkhWAl7wNIJoO2s1/4G0c+9dP8UmdPwD3KX9BikvJTbwEj7dZdw/E/wLLRxR
2R6OcrxUQtoAo3LZfuhfX1lfBfWwEJ/x2x+Z3kBjgMOY6z2ZmL+FZscCaQ8GL+ejexcLDLWOgKWA
UIHhX91gU8blXJIQkjH3/e3FDQdemm/pB/Y3gdabLyDpDS3fbT9o8S8GXcmBAgDURa+OafnRodta
PniSPuqkAJFvLpIaVIhNsQTjU/iendOSUIRmb248bvhg/ZbTHWZi7a+1s+/SD5A8wjDK+kMpQo+5
9gMV+yhavH1qR1C8CGXgixbvAAPHgu3GFZKyPQwpbGQh49ABFOTafe/7Wwc9R/tYJmD5gRSzx2AN
8S0EN+jvIHiP300VLqm+kn55rP8V54YgDCoMssCqzyQoHWYffymGDdvvN77g8AP0+Dltv1P3H4HA
/lMPmeJOJf7n6v5NLRidvEyCXFbMaYvMjFun7GAYitV/rldO58/uXlkATuvg/K5WMpYN2vVsrjij
QqNUnw58lnebEf2ETzZlrzOuR/s8H9S4RvjBvcixdNzHTCefkP3u/SRG0+ffKik+Zv2iHNCBYjGg
2IZKXWNBUD6ILP2sKy4fJbZ8Yr66Z/ao9mUvqYgNsbGThbkCw59GZ6ZtPZWRRzFt5LNcPIXRszFM
fjhMcXj9FPbM0iE9kFvLKHoGfHbM5YRaCGyq6xaba5578E7IhxC2SoE0y76ast+QXnv0zSfCMqLl
x5/EMbzqC89jDVs/ZHIgz3FiXYBpCui+zT/V+aYy3s1f7yoNF4LAse/uMy599klDyP70HwMngm8R
R6TNeTBF3ZTkWfVR1oC9rNkzhbhk59jChnq+v5P4tPvv3IKnsAJPGlpsK37Xtc9PshQBlJt6EKQz
AWQqokRixbezK9ZJj2c9IC67fbeIGDrvzvZcNGLDYKn7TcQJnVUXOeJOgl9zvcbPD7kLLC3wAmPb
kGJaPsRR3z2HLd3SIXL4tPnbOjhGRD2G2Ohx9QFSqY97K6W0iyc8IIxisHEO3u6LyoENPUI/Qe2J
3hqMhDULjDIm9VG186YEWAmvVT8hAWQD+KDUdnKADGB+nYoilyNg3wVLocPL2IBODP7jFg5diIPk
NliQmv6mxxRwQOAyULqjFAOzVUb0S6wF9fugwPHAiRRq0lyf1NPISFXDqFTiv4NbbkNIFXBRrmPD
2hv1/xmbgTfe/cRI0eaFKzG4no8eWKmQZeO9NE4Kh2qUvObYzih6YDogOItiJ5jPNtFJzHaTj5TU
XKTHxsvTeu+nBjsdZZOKaC9+0v+vFbQB0GHEdMkJ1sHrFQVfqvCHIUSStNqOFIp/GAdFfq2H1eEB
90vw03sJTCbzv/JxL/kjWEwq93gr1+3SI44doN/I8YzolfWrFVGCLzBxUFi1IgM7KlMR1qJbz6l8
W96Gq4chenLLosieN8M8Zp/LFMqIH4xhswki3B7vgNMENSUsc0DuVxg4eqyAZfr77EZpp9t8U/4M
wupOCbOGtX1Tk2iuY9M9pKvRXo3lEpGr/WOjVcscBMdqL8B7NbVC0sZ6wwhDaKSPuuLr7MMf/29I
1fJeYORoyLwmzh71Yf8iJgwqk/+nfawpPKF/NqjUFJrrwCb15Y7eZoBWKscZv8EUhkzPArYzKGId
KA0Tgx/dFEJvbx1i4bXQvLKuR3zGMGV4NhRjWzbarrd48C2uQgFxElgLMHPb7jmXK/uXX7b5PSa3
78XTnODbNftqGWlcvpeb27Sw/dsKI2c3s6eAUYvLSoJgMl+LMxTU79qhqP5bWvRmE1cG3Rbu1aob
pdqX83SM/4lB834KvWo1uB+CJunOyER+fptcfRROsOQmzjqxoLVG8AFBdClE3FjBKRKI0FKZThs1
HTlisaDcfxbjmqLeEQi8k3vddSCHUYtKl9CC9aEMy0eke2+mfeyqefVQ1pboOqwzCIFaouNTQ9i0
1kU4inQqWm73zsnqIEIpfrsc9kgvzHCSBKmVRLhozy69hDFDlkLwsydxxH4aat7V5NjdM8QSVD9y
C6xCE0fjjZ8j1Z5mqKdxdBbIVILJQuX7uTxO/m9YktI2Yncanedixvt4aF8kCXhZbAOE9zezMpE5
tdJcNBXqOSYsJnqDxbOsEUdPX22wShxkQWmUlfYUMgtSUHRYhtdJ/5QGU0fDWZugX1Xfd8Uwd+Vu
19to/bxOK1wz/sFZnqe+e2NluHVtCzXzDjrmnqxEmNAMbPi3Ez3IKV1TfRLSRupnuKgz4ZZty03L
3MgDF5YXT6ywkIsQDN3n0Gbdwfcxu512S4KUMrxeIR2YwZw1HGdgeCsXfHH/H+IodsQwjSzgQmjY
NbROY+qf3F1ffjg20QwX+nLWExcTO0mWVejqslL9wneTJEnfCWnZODF8sfOAe2lEVT5jBUQ2FqR0
kiGgjxDtxRwVnEQYWUNwjd/YaewPIdkvHaf7EfQDfoXWhmF5Z5ql3stAl+OQFm/np5k2vLd82sm7
+ByG24sd+TIbBpp02HaSnWX0cv31Ynz91FsPk7bFTyvgdp1DUpPomGL4HL39tZB3LrwTKvWJEei1
hl4YOS4w3QcyhfuNYG6zh99qUeR1Qmiu6ih/iRj8b2qUMP5da6o/GaVibti5yMHOS5gRWriCNdKl
qTlNPD7ktGGMM5gaU9wXmPmj++8Eb0Ir4raiIWPqWIL8Q3UGEZKarSUUEYbaIch8M8TloBh9CKA6
BvfG8WtEPTD+LBw/Ww4lnt4mgN+BEUt7u7zij7a3fA9UHJKr4H3uvrzujs19WBVo3HcarRbDDdzt
qcV5Fb+9+KhQaWfvLJZR/9YpcWUVX3Mo62VNXfdqrxc4jYAJRPhHrjKJbu7IXvuDZnRzuUVtihi+
4k/B73bcBZ3cu59DFPEISFPXGqF2V6aQ4gnAWCGbv7VGz6tMqhMVvCj9f5HCpC0jMF/UzZChXZDq
zcbh+4ywwlvm4TTMFLKZMgFwbeHa5XkvteHQDTGotQG76kwDovicLP11AF2M0zkc11OSVrxmq3B5
7KflFMtzS2L4ECc+jbb92s54UHM6Q57Q4pENiPQCnRW/eqdEeEqNUyd5n6j0PQbHB5ApvKrQtGmY
+e6V9lLpgdV+YP7HtfSgSff5EYg2UVs1s41Kc5xSO4ze+2swuy9qgrTEY6es+m7RVUQRc+nX+E3t
QilS5oIKWHIG6kNRvKRwvrOptu3IdzD9rJpdi83h9KKQlLgkRFBddOiSaWH97Td3ycwWjb5ALo3X
AZsRrv8kx9x6TpS3olO7yMFkgJZtqWjeicRXMH76OfJm+ZUycOJ3AnV18jfhFfXFG+ZxJ3R8iBvr
mgstUFQmEPjibMVHq9+cGosUXIbGwIuk1mRuHdJ8KJtZSn4eRWNE88uF2qlxSVNehuhH5tUFp0SR
NcH2X77iwzhe2GCRwhF67FzXsC71PGnnWz35ORRlCXy9+1mC3PATDNhxURFTxhZIy05vtpe31gzv
L+ITiAYApTLm4qUswn6sE7uqt0tlVVuy0RvmzuIUvs5FwlDWPydzREJYkH+zcJnHCD15LLfUeIoP
/zfp9d5jdywRarVL9RDJAAUaMoLIFUhO2x1CEZp3P0desqsakoqYnzODjZvjibr225oC1cFUPO9Y
MA686U2cDMSgAHQkwI2GBG2T/MSXkApYyUiQr9iYGjXm7E2oSTQ+i2P2w7XozMDPHvvtlCMQsqSg
3sG8YLmdDkpOa9JEBAgufV3G3jZdF0Z1V0vl48CqbMN7i2RI413JNQ7jnLgMKf+h1v1scj33ahuC
IOC8Gk8Ww7+KqO6mlQmz6uCaoWqNflA8D4q7aGRct7IxJ2toyx8o66vL+pvDxLwYtflZGGIkZjK8
sjvLMT2zFFyQQ1ja99/JphvQI07gnu3ZR92iTYngbX2Fns6VlO9I027zvYjYGeIjOCM16+IOjKYF
q+OPwTixv/LG9ZVCyS2EOOVrvOiEezpmOrRv+6pmvG3bWmVxGpNjB4MYfNZm1RUxkN8h6iNPyXYB
R02t7I/tOwWFGM7e6m+NW4DtaRLsmF9K+8F44XPY6XuXsG/O/jca66jyLJoYg8m38Yy66UrYvQIK
spAyr4LT6F7Pp6RcmiX4tRJmgQKm1MOpq8W6TTMBLiTYHVrg1h89NJ5ueiUMUNJaMqmyblvDKXx1
CdIS1lCkE4ooV6PGMJ7/6BIcrmgw8njyiMsnPD2Z3Pr+ykdNEyX0SjdLdUmRrUcDb/PNhJyxi9i5
POb7L3utFWMzCZRLa0MiJmFo9tzTf7r4sme/g1xsMSQv3hPlRtoIxUHF0sLs8ZAn8rMq8ZaF5xar
W2RauMRVBtr5J4n/UBDkVWazhyg4Z/f9LXKvgS/A+cLi6QW0SUBIp7fa8dHvTQI1OB4H+tDUSYBW
nIC6bmz1ExGO1a27+CVClpHRCN70hESG+sA7ILuBw0bCEEgBYtmVLp8j+sy+nSEPGvCTY71qlLAI
QVjaEJsw6PJruyml4lUAB9MdsNjcN6EAwWK55GjKJb3oWtzzE3NRnafjkzrJFhETRYkAPrWSNAXN
9YO8+lHTbxEx/+JMPK0Mh4rl53mESFp8yTsgamc67PQa+pUOT4l/yXyyKlqoV7WdVclsSmSLHmFV
6ywyTl6m5lEXnia6XCQbdrY8d7xTFof3LZt5+yVF3hcjbiuD9fCK+10AerMxi15LeqUMspj5T5J7
YlVKUdhJprxN4RkS7j62+jJkW1SzkjTPR6EMY/Y5sRD6QhPheM9WdeN6SW36WN6DO20djhHmLHnk
eNLwhyS4Sdqo3Qigar0nBOuK7pCLQSmVd+6PJ3cRzHd09GtbeQ6hSqvumSjp8Ixewp5yWMHHO5ZX
VZ1zBqa/tfGWEsqb0mAeX6uByltXXfTB9+aalhOZ0YNIfrA12jthutxICYLs13CsM2l3YxAvW6eF
WwRqU1gKCrNqzDsNRejHeCkNW//hpJh44uyMYezgoyo9y6umeZmNs5wbSM60oIy4Gc5KZT9QeFUr
OugxzpLRS2kBKS19OOKFps8FL81dYUiMCeK1jXvpsEql0kNqNc+24oOkT29/iHGlQDw+03raSHbl
fQtlJ7w8fajUVG1ZTAvGA6l99dyoPX168/EoJu/YAwDwOxHl6ucR5sZof15FA7edvl0OgnGiInCf
Oo5UI5m17b1KTU64Ey7JTEi6KTOLxKcz7YaZKLMFm4Fs3pCxnsVAK/nd+kpD9Ej0gVrnfVXzV9be
D4PXtf0y/MPYtunLN8AmWcLdBzzY7FiMZBi1GUoUqnY+QnQQmzhFPG+U07qtZ8lZ0CTrOJmw3uaH
pbJj0eJOkh6gQwwIyVfoGUBw6lt1jQBwJNnzvzJ9iFPgrwkNKxHKQjBRtjVUQCRKQDjh1xxlwqD8
cQ3U7ErEAGEcNI0gKVizjnVEaUgeo8sQqclnU6p5rzII8k8SM7Xm+627/hMrJGNNawgd9koD8OOJ
12mm6NKn9jRXGvpqG4Sb8hK/sbUTJuWGVUPnuImfXaJXSXgo+uM5knLADp0lmEy3pt8hP5I6geQe
Q7UAhHL1XG7P6KsdINvnIQ4KoU6RW3CG0dD4anvi0KB/rIap90X6R1NhTXofdT+QXKs6dp1Gx6ir
2Z4quTER9f9/a+MmUgYAtdn44sSIb+8pCLj60jsLtA72VTABDTJB3+y5jTMUPxvrb8kqrRDcWlQB
E5O59O3GKbMgQj7bMLe/Chc+Q4ezPwv9zyy6v946wJQRGwGoeBL4uGgwjPkcxuxzhhUbp9AKilgc
iwB15AI5Ye3S/nIj0573OQj25YS7Tq8GSwEeu33rfk2wg9nAnovP709Fxz93bXV4DgRQdF0+S/FP
RKI+qhQCFsDWS44zb9iPoXBGkLuy2qQ2v7I5j75oVefPwvii0rEAUK3JJNr5XBLmE5u4Ikimm6z4
ok6c2ZX3V3oanR1SXuAqhrEjN5oMuB3sigYIG8hrqtmp0NLVb/LzCjplpb6qXApoDAeCS1bfWQZK
bN72GzGxXCjcReVNIxh4DXwZ7q179fLHym+JeEehmBQatGYfSYyRDE1R05B3leGVQ+iqMA30yY/D
Dojyalk5ZK3/NstiL6/zDqvrmxZjhQS9ooXmjRPI1pSM953zOZD/6S+v/uW64rvc6gTMTFvJx5D/
lBkpd0TZ8T4JyaZcrNTHv7CsLJ2dsG5kMUj4cQTB9vdhgdFH9dHuq9VP8iatjuUjWBtMzPyno0PG
fOk3tssC1VtWLjDRlFt4HCYVYGL9bLn2wo12wRqnak4B3UFOY5jNkX2VHUCcmuNLAu/H1qR77Tvj
yfprmzC5oOFL65qG30QY12eWflwfd6U0CqPhqrLDUMjX0UeV1BTrjX8tp5ydDd2MdmMIbLdEg1BY
tDYWFq2AyTZmI6yIYEiibmORjkrgwEJ7c0GvZ8P8vgN5LqFIAv5YTeSVIgDJhzdHFLmtr9t8qAi6
Rpvmr24h0/3dl0vwzh4BLbv13hKuy9DbhfUveA97QM3j6PYSdKihxPqvJRmETiPuvbqsiG+wgtIA
GiGHeNwu/kCw0l0PBrR35Rukr0q7TcEXTxC5HOt50WY/n2pSYILDLAaX+V/ZpBC5HSV2D48qTgFw
1L6f06vIYNXgeD15ZSxwGrERjlIELvIBk5X93Xf7SoddjGVxYGX40AD7vak00CSuCuBFdgYT6mOa
Kl3dsiatQeISYqzvh1PPsFJLa6SUScJdO2JT0UvmeMe9BDI9fhh8yRHHf6plu8CUMwx7upkcXi0A
dG2YkyZGTHr+4zezUashj42nDhi2qx3zWAK+ZgEW6i2X7dxUVUKlbayCSoVWK7u8vCTB/dj5gG/v
P5qxdswjxQHNwJG2wl5HSTzYEVdgTjNcJX6YwyAhhjVcXlxNoBTYC/nJAlokFaSCdfFkhKnCNrPQ
DrHFjYoT6WFsCXX6ubWQP90QRSoI0Cf5eCjEJDugWOZCz68IUCehDtitgGxuVPwybcOJPXlrbs2a
bes1rj7Eon88zXd9IPMXUxC/hJP/MGxElTAXuLQXge8Rgd6rv+GMGZk7QnKN5ywyRi/ypMn/zR76
hzIM/xkfCGgF0FFmZOtH/JDdYR3FCvmGeiLAS2VAZi1WrPwTsedcKGthlqgibF1BnboNZRV7t5Bu
6ThOcTrHjQd/qpgQ8FeyR1CjO8ZUBnmeaK9Cs88CuqkDW45uNBWKUg6G0AdcFL2IM2hLbo5zb/lW
/WkcazKVZ7X6n4Dq9CsGWNRmDkLN5KsFCnZoy4Vj2dstr43nok4KrXqjj49OJKP1PxSrLWUlHbC8
o/tanLyz58n8uO5KAomaL/SlbW34LhQCbLbEOg3xYXOGYX+OK/VyJUty+Fdqh5t9En+bWrRGnTQh
CXKssXdn7JKKabeWN/uBMlb26manifYcZ/T390XCAHBw9aZ02FvNP1UUa7fAKdeeQZhsXTcIcODC
qeZiFjtuCQ3WYnXDNg1n50gEmEh3jFOk0ihdQhk3GrLIrRzjSP/zVU3URI3DPsJ7KyIq63N6nv0R
dcUrRpJW+fVNK4GUuJgPj1qGq6uwNp568bh37K/T6Dv9Zme2saEx4VIeaH+duHZm6/dR4qPU2PbU
BQVTTH28bQpgaoaKZ5MwSxsvCaU/QL0VrMAzhPdU6Nx0hzRY62sWZalpObNBrfmTenUGEnsUUe7V
gwHbS0tLu7fU7fQnAk7e8Tdk06ZiPYTdzKJdXTsiSN0UsFhWsa5PSHFlaVW3mDyvvA/ZXO+UOhZS
d9+fewtYx+Yrnr5xM86ddWtB7VyjTadBce6ldQnvoBcf6O5e3w+I/XxDBN+ZoeT8QFxif8OXGULc
6E8fKz2Aeqslr2BjeROI7tBicI0HVRdofjLdY0l7myzTOJRMyFJFpQk4+ATnZR+ZP4ZF0pAjX3Kz
Oh5fyRtibivSlhlXBJki+Zu73URCix/rwUPjsJy6al6H0jGY42w6ZVZNj41F0cHQISXW+O/zSnoj
hhOgxKeul7EPYTFQ4yMcs9v3vaQIRHzizMzQgXf/fDWLS7rUIy+ivoKM31OEkiRmBrQOKfkHsMZz
yJJYoTGQiQWQ9UPKXTOABNfD3XZUe5nKxwTG4ghCWwh4JcwGz8W3VueIVa0/3KKlxOsOFQ==
`protect end_protected
