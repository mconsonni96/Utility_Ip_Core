`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
teW/h6zSV5cVjVnHIxs3ukkLrniDjzyBwJt+/aMmQhl09OahHB3yK1E8ninOdR6N8Wm/100azzGq
0bBw/AV7u7QZIp60h/cgtbULqDCUYGsqqBoSQNBdPpQFaC1hpTQ92ANlJB5PCVwcQtBpNi5VJZt3
Gvy1xdfPtmTOnZaNBIEXbOV4mWBRfivVAi8cxE8CQeD2/EBCzZgy2YuE5/bvGiYTku8ikq2YOT76
J1//3bQgMmVJYhA9IaMiNjttmCfLYZtNg0Va46ugC18QTHs5QPl4Gqz4i86lUY0HuWsmt8wDxv58
4h2xLfaZ1WAagqoytQuL1S3GyMox1Ut8ugcV/g==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="rfKUR+IC67YSl8ry4XuukHYaBNkGgAK+mkNNvr50etc="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25088)
`protect data_block
rP62sQWR9HmTraETAUv9xZhNE2a9GdqzhbAKedqjaY0qZPdyr2mPXQsnmHJhZK9qkWhYp0RbcsyF
wdCArtzO8xzv6XlqcGCUc4znWLrsH/WEb/hp37zrJz7AZ88DNyxf7voxBMfYHVLeqW9/7mJHdsbI
Sft1d5GnRjus0Av06yuVtSoFFgW5tQjjb0K8S0ncepUiKI7Ask70J0BOax1fsK2ONpQHHYrcdeTD
u1S+eApNugJeYd3JkVpC11MJu3I/x2Obrp2q5h9hFz6iy1mG/wiY4FVX5Tz2w5oOwPrd1vO/XcSR
TPvGuv7afc/RchQIS9vmk754wdFhyDuWvjzZ/dORhkrdBfS06ilbZNuPYfa7w3OniNRuISidkXn5
/dQagyGC+r1qHbomLzk1AhhdQBFh0SpNFV45l4jXVYGly6rLoCy38UkyYMtW4pbtIhGZRGt6Dqfi
WdHw62vzJR1CFIZ5BhNTZFx0j/fGhkCxf/fvo+4QNx0djc2tH7hFEV0rZRvqTT6uEI0B0nyCTbIh
zOUNr1JS+cr2k6sTq91x1DzCi6fhTv4WXFlrpjpDxKZjRXDMkf3vs/+7OBATkejcAKsnk+fdejAQ
Pd7+/ZBl3J0Mjd+3WU+ItEXrpyepvnZUZZNCqHUOtwLri9nA//5lWPDEONBHyHFHmR1mevW2h99H
GF0tYn2TF8/qOFIVm6DbE25zyddyckmW8Xs9z+5SBAjroBLa0SFv3zxhSVQyJxdyCXNJmaTb80pj
CxH/5Vn0j72hjO5AF4s8lOVrp3xoOBAw4czBe9RyBTv3Y5pWgNkqGL5NLvK4b5jsw3AEwbBzakyB
soDMTwF6lxJ0CdEqytO7yZO1CWCBOfsTqO7WvEq5xvpkTDs2ujz4psZ0SlSQLNoWL0P9htgy6uQB
89Byr5lI/8JoqoBP/lZ998WbEqU4IAiCovKyBxuT7oL8nMB/Vgurd8hX0KIEW96sOLHqDBtanM4T
60ayCD+ZXqW0jXsDlRLETwd1qeG4IbVSCav9fgcpud/LV09rCSoqHSl4IoAqQd/g0UQzIlMY+4qT
MJfYyFvlk/X0nWVsZLsNaXsIGIEgzkc7UQ1/8x8tQXXSqg9B5X8hRXWGqpuK8xvBg0SU0ZdvO88u
lD3DucCmhgsp9upSvH3ecY2dAS9xuz1YOG+xS4oLAGZ4DyywtC8/mGGyKUmugWIQnsO46OpMLcbO
IeMUC1myUD4UrbWIZsWV9lG3rGOENVKASBRyPI/myGr7SNSwdeDw2hLCX5y1jswWuYt11bl1ylIn
xxnJ2GPWtM8+YYFRcdKH9B6xJ5K2D7ny3y9YpDzMC9xT7q2a9h2/cUQdD+UENUmMi8D4yxlwMwrO
M8AbdR2qieqsDQcsXl8H3+xb+rSWP0WC88aCmzjoRO3krcI1EOKJTBV1nJd9sP2x6g+qhPMG3OsY
q2zGFBcAO/7XhBPdbKOVlryytEJ0kBA6Kxj7N09IC6U8WWNcCCZ8GQNI7S92CCth16Ta0m7rda1I
timy3RT9KqxB9Wcpkk3gJWEC21DlV2kSLi0e9oZaDR/C5S8BYJ3muDxJvFu/ZTKMCUj9gvwH+mCz
zm8t7jxjOiSobuXv+LEEVfh564IZ+IgjPckd3OPX+2Kts6+cW8CO9DOdS0GswcM9mpDaKZ3JGfQ4
epPgzJEkDeXZZ5NfCbyGQ6l3AgtZuOT4cRJZF+MZzm/+Szfo48oCW8tFuwpHIqyNOD9K1gPMS4cx
/o9BKWhsaPrMqVRk+PFO369yRZ9Ss0QvPP+Bbgc7aMbnE+7vXzDsJWNazRHaIA+sr/FqysqQXvDL
tesoLg8kJ8+LydzY2LFd/2ic74dEbV6uZYMbfEc9nF6aqXebXaZdBmiUSugY6HH6joHpvI72Rx7D
AcBDZ631ET0MFMLCMn4RlVTX+P/T7KNmkeVEqhKmk/Qi8/HxPb5HSAhMehrxqv3oI71uhX3DugZk
8E7IqMcVNjWIitCch7tLizOTtOQY3krMPLYNxyjK0s5U5Ddwz3+vG/01n0qFrrCsC7A3HLFJw6Mw
1DoS/R0YCTKxr90JR9Wtzasnsvll9+Jky1kCuKzwAMgv9S/I43nstdcFtLz74hy6gwGiYdzorLMg
pF2FzEoeDSTTEI+ALYshz3xuApjrmof9GcCb2yxyJQLWSptuwr9ubgiz1X3WcCRlWPYQXKar2s+l
ciayU17F5DF5+EfkhnRRX1MYKlbWXdMH5c2DSg9bYIkuFqprp6qIrp9GJal4PasKm0m2bDdqY1BD
FMy7qXyVDSVJdUNR30FSi7sO63ElOY01/fMIVCxVq9kC01gCkxUTCAvZyhaZ5u3lOf91OUDJXY0A
teFhlmK2pgkCOr8RfAdCtBJMaR9OOupQ1dZO8tRNnrCQHzki/5YGg2pKvqJtGMuXX3pjF7i5ogRE
jpjxIxHain5eJ4oDKyun3cJZmsRGXvSCLFfK2zwZqGwpgUdsrTQ0uM6nQJSqUXFcgb/G3I+rRIrf
jTpaUQbxJ3ehJvQhwlv1J9EUGNPEb6WgVZstR5H/aCphxjyvvHgvsRRjxCH+nercuyJg3NT7EtXo
pe71W/3f9o2Qg6Cu/E09T1OjIb5kLOxOKlSy/I4q5mQa/aYYkzre13KN8smNxr530cj7WBFtmCUz
Oa7oczpZNIyP5J78DZHHJjI1K2L+KmBExtDtiJpidG1JLQaTQyM12K65seyoO4FMC3nC8gUoN9qI
X3MjiII4+URZtFUefrZQ5gP/gSZmzMVzfsYt7nbDZa6CEhP4bRfXp1Yp6zHZW3U/hixeHgB4NF1j
uFmGl6yMnB0zldC/047ih3XHHJTZ0FSLrcmfh2KzW/ezMDu64x2Y8LgP93QbShac5Rs+CC/u8jb/
03aYFO8s2LNaFFiYOoIPqBiOtzA6m/pgFwzFqtaY6tJ9LFVfdO12xmJ4y6+DvGCAfy++gmKhQkgb
rCJZ+hZPuT3snMmcQGz43Csy96VRIZxep9182oXhegGO6cmMVdr2EcFPfRa5Qj6V1oKAcvJyIsx1
O1KuVoalXkyddo1AESMyBYcJO5dQTDAjwC6OiHCVAVwdAb0Wz+B2NHB+cpJalKBH/qoX1YLNRetZ
Qv6B62yNKHDLrUNPbVKIs2XT50SYy+2Hf//HgHSsWd8t6DgNLC5ujQuaMF8nfzvJem5Wu59Gm5N3
I7ZdkgJ00KZ7PhVRozBy2/Ilffb9joSF0sWXAn64NhCgD7LwZ07ATNUxuaVf4aQ+LJVOBSfH3Ti4
bn7c60plg8sRAbVvcMaWWJQd1tSoFMgEj4gGExQW2WOZQuAxpykt0A05NgwIzgfBbbNltMzgsW2S
1PYR+yEAjmAeTMyq86V9rwl+YTHnTmwMhMzan1QppBQRjvV42ZSPFN/6zdtmyg5fju8iB6Gsh/hz
I1iHATY7+KmCIurf2o/8SCa6EXUw0E4qindWj4YW8Vh2h+s/Q+Q0qWf4Q/YJRqvQZBCyTbVRfrLr
dxBwEfGV44IIC/pO7gYO0sK/vsslk6ppxOsTCAWj1H9b2LAVHxVPFmKwCAH6vIedGe7SU4QCPZMH
rSB7JzrPGqgPJKGTn5JFXaBMVo6O8neOBXVv8ZJ8GjBN/JMAvPL9EJattw55jPaGtL8aTqNWZR8v
d5oCMnPEAuELhDD/vLBMhP3xKvG21+6KmT1EZTg+NFWUpmCXH7OBjDBtaiV8Zi2INWBaDE2wkOxS
RrAfT2uAxS2kxEjJ8ZQHW0sAZxlztGIQDdqNhDmhZD4rUH4b10SM6T+Ownxsza5BhhbQBTeSABHu
Pb024qezNlG8UogtWjXDL3EE6yWu89LaJlSbH12Ndyz06xlMvpYJucAFLo/oYlQ3DI1B5iAabyy8
8vsScttS8ENinyTTulDCqCzW8ZQ0nPJJmFeEyQ8rhlTuNapLFYiOdsQq8zk3pI/RFwSEnovtA7dD
RjPhEaZEgtQBnR5XSGUZolMZZw/I/SwM2iPUFDuozMXubedJ7LwrrteoKNKihvcbp6pOxPctcCq6
jdVU84b8I5EdLC7xMEtkfGvVlC9wkh0P26fWmymprMoIFih+xwoTuFDxo2WLCcSZNR14LQhWoaKL
A+0T+bN7C3TErfYVuHvNdgEhkmvoRDVala49jaAiRlLX/rL0AfbXg3Op6dcIl8DZCaudEBUqiOpF
Kucm57viwNpFUsVIc8LEX64Wxko3UVrUsGswWrWWUQrr881G7QwAgB/qqj1zulP+8Jbg8ACffRuz
Q9dfL/gve7Vk3MYk5wmejuWJ3hvKfZfP3PkAvOGeycqCNIvlPZWzlQa2y9SKLsp+EhdjB1yMSF8Z
Wuxt5BjMojm3pCsv2RHC28YZRrmBDuRXNB1KWTuAb+DF6sgAJ+ekAVf6f/M5Y/oUCnxJxgklFtX9
EPBiZDz6vljue7KyW6aCaqcZRAMGGye1U3TCXUyflE9x2cXzLtbICYzbh6ynLrB2clhFDa+liYo/
ti1t3wdumJq1ZLvq8LSl/QqQYgFiyO1EI3e0tZsdyu/MpaXe5KTLtexk5aKQG3O6ibipR31rUgh3
cm2/1rpuGhPjxn+WzGFH+nEc3BgFlnzueHBkm3nbWsHwuoCrrmfYt8NDZ15HBpVYeQnYQBS4ozhV
hggqZj/Jxmx5R21rlLxumIGYo8mIYwWkfh4AHtxM+ijSMSrTD8YbhzZAEXorEuUjQagBmZrQnZV0
fFT+3bq+nree7OVj+dPdZSm553PN3Sb5140aKkAh2gDAY4SzFtozhkvX145VnFtNPCmDvVWs0vK8
CmaJHA5WdopSPEcnv4zWnWtmhgISYzF2JqwAoaxyOLS7f+qJkF/cdbx9/E7sn+i8MNoem9s0/apQ
LKObiU8h1tMyV9vEMeDv5XxPelJB9wFGrLPLJqIN++TBbNc8b1u3GdqIAAo9Jw2GUMsky2i7SfXx
3Bo7FKYMm2ssuM4rlTfEZ/3GEjoGiQMXluffpRTLpmaBCPV24yBTx+PdrJ5PNyqfQnS6Id+nxYjV
t3UqL465J5Ow9OTrPWAfnrgZwC/ZkG1xpiIe29Vh6PaMSFH85cTBhjH1Wvhtr0fo3DvBTqZGRNMl
1eeLSc+9jbhv0+SAJ89esueEUcGJ2vcxHHmO3GYoYcvUc1odEgkVXkc4apwsFOBpOI03E9T+3/9f
pXBM6pPXE32eHtsyE4iDMSz0HnwAhnv1YVdnzBqoHrhsicigyDvaA/0FXc5E77GX0s3GDpkgcjWC
x39PKMKKaEs5jXkugQvJWxWXXysRZAhUUC4PLGqZAIEVl0UoiQ8HuX2djzhN3ht1YNF/9vC3plla
8K7KN1DOszgxP0HjrhuXg+6op0qqt1RZPUWoRLDm4G6WJ7un4FY+dkyVifwRQwkYCbENIy3o4Eck
OaZSEnMTdzsWQAJ3FoofMynqh94IfxlWVGWyOgghwotKtH2wNfgK4jEuVqHeoGewnC+peaUwtsSZ
r+3zUab+kPhggWA6UtLqqUVfP0eSoFdvoNJ0SflpVGNQZjyCNiG/4VaLircfsrCLKdRYSQlK+XCx
zXPHoVS5UNgMV6qlZr2YEy05HL311BHfDIqvf0Gaw15OcaMPEJr6TMlYgkPID/oSSFsCl0hN6zr9
KO6N8bBUKgYa/SRAkX2tWEQczHnVRAExBsllry5Zx1jAGbJ1et+BgcRUy+yWoO2dv4V9YpMyPiX9
0Ez1WvhkStqutVPF3ZwJEFx6zuGscswEaTHXXLoFL1lvv9S1LABQrahaCOlnM7eqCEkkV66MqChy
3tBmVWNfzs6RkMR3h/QZ44U1bbrPSyD9txNbS5LhjYMV1czneYo9FSxE1cvzGzTJfiNAjBIXU9Dc
079ILAduxSRntxiKzR3qTCUDFB3lKR0WCG0+2gq0jh4IGHFRH4gKQmu61tMVd0JzXkUxwli8Fd6H
mAVdGvRmRB8VUV2LBstYwxoPNquFIhTc24QLqNecjkmwnjTtfNAa89mZdMZB1UwbxyiTe2pyLHzc
tj9cMgr/o2Kq2+sYe3i58hkiLd6rluGY7pc3Xzb/o/CpoDT9LpPgFuEjVkNhOrogAyIgUu8YnKOC
CSdTA89ZA+2j5A9IbYqfNciX0izWI/ORTzD0TWvCPN5mdhSTk7NnzAvVn+OIADMFFTNOX2lHUxBk
wdL9c+bCAY9HWaNL9g95OOE8u3EcBzAJniCqIM/yzK+yOdHlZIPFj2odcGCD/BA82C2Sl4bDlXqD
QWr3japP82qKy3cv4rSmFyapawbfHpKhSk0h1Y5CtCA73WUF0pAiIyhlH0QCOxxluAFIcWmhLf2/
vwoi+vKe53rGpbr5woXuGGEcxHK6bNinl3iKxN/5rnCpDLZoBE19MImS4b/4FBKACThFNGiVcjYt
wroRhRz5V7Cq5DPJUsTu+xk0WsiZpIcr8yHrStlAI830ooBQNmrpMDV4HBAzg33pFriefz/GA7/4
hi+qG/f6/77Yx+Jc9UFBCa/RKLcPEiEKpgxgS4GidTJ2JH5PbOyafNRIEdJgVgLVRWn5Q4e71A7f
KhTBVZ8wWoXPQzZ5w2mEXcJjOc/b7bK+qrEWUhQCQ5uXHaOMHFf5Gj46WecCIbiolZL6qkQsT+wD
xilzijJr3HSp84j59U9qUdmrFXVrMDENn3JrCGEtEB1suLrh2+gXLdyhko8dnM6jwrLESfjElr7u
PPqeJ9pD7H95tFjSlJZv8rjZFR5zalUMZfpsDDcITp54Mm5gApAOfRt0+pHSdx2fS/9hpCtJJ/vs
kv57W7hBWOKXuulBWwo+IDxRPZoRBaQOhshi3PKuTexmQryjq206ZJN3zyY9frnUI5RYHKixI6Dv
obu4oV8BzczlZDxYl5UWeBXXkbQd2Uih2ZrlJ0t8pNY8DZG6zlsrhsUsyZPj8fB3bvrQpBPhEpPw
CSWA7mg23jqxQvyHpGiciCfwD/MTlvMeIK1SiXMZ0ok836TXXFS8ohQn0X6UWmDVQMVeQLx66Iqy
byGpyMHxYmkoFVVanEcw8P7rWi7o6X2KkLYA0Qi/gOeHFBiXgOONfWwj4oulyJb8Falm0WNXzZLv
/Y/wFIGC2r3GBH4mgvOx3bb+8xLkOmp3dHiGHQUg0rhBpvuXVNWbXe7qHRTy+ofKW+yk7aZEHDlc
DbxcoOq0d+wpJCKayRIFDWHed+epAriTQmBMJNNC2yMEw8qEz/1R9O/JVmT/rvITHk4jMouYhTkM
tQ/quMAN16l62gql3I1zCTSXixcFxP4Ux83Ri5cTADM1hTsmTTEL/lCiVvDvkS2kCHUq4eV4fxwJ
l8TcAkdchjbmXGQsTDWrZWpJRqEzYYsE8VY4CXa8ObBHUCDBJQrHRMYQEVCqFXsTfSJHZJOLlGuv
yhDRIIYbCmbRwsJVVKTf14maCrxtuiKlDTarp2VMDEOUKGN5LeznQ36YqioEoGMeqbMkyazT/CjM
EZ8miGZp9//BIuZnsiyIXq/0d11zW752eYnODEBtJ4NafexybdOAQhOmQf3DpAHqqEtBekl3w5If
d6jy1NodyiaVYFY009O2qHgOyQMV0t983ktj0DOcbexWwl+QijrRU0RicDPA8kD6v35aWkmiFGMf
NcSCZOQf166dQgmXUDKaCRwvyiNRKunN8kQHkYIFyBYCLbz1/v5q2KDsVSlg2EvSFkQ6v2GWlki5
ITCb6U402GnBPD/uWopPgLWeQfSkDXQZUWlw+rOKFWTYKiFQs+YBrWwHhDnxj+LHXhlu8yRHrrZg
DSsvqxBdN8lZEZzDK5DdSGXh/Xmezseu+QexaaLisgR6XQ2WIs+nzAPdsoIWLAZVoIRq6IQxz/CM
zhVZOxUzcWeW0Vb3sB74mZ3hCMGMGSmZFbrinL9MbYElCdwzqvJdgtLVekICvtDOUNGH2xbb1aEP
F6CCW26zV0pAxGfyM48m6tbFYnbdXJoLSRCZm7iYuhrZPBXc25SjORzeRn5S7SKKwvZ2K2Ys9BvY
WwR8rirf2rY3m6j88Lod8q4FsSFRDABESrw6ktIbG4EnaXQt47ZLBXDbrrpsH8sNzNBExuqehAvN
SgAb7rO8DOvB9VZEoUiYu8/CVFK9ypdvWCOid7yRBEx2oJ87gbEaFQvGOWq3pHsDOal1YAMRDrEy
kVeECfUuvIWavMPiZjoXajtedXLoq5pheZMZV8azrAsJBj8rAMIGVOkvsEqQWz3BrEKU8o5peNuv
cmD3pu2f29l1P4H3uNLBINQjHvq+FI0YTZSFQaqUmHAoSDu6jCiqdO3fB2JBC0++2V2T1fOcmp+j
TYXMCkQG0jxuk0ESFgeYNKLR7YFsUoA3BZt3WVBW2FH5GGA0l4E3omfUIyXH8XsVHjHZGurt3yoI
Xl/EFXfC6ygBbowniYnyX4QPG43rgMbz8IYDqG06aPfCyAb8GqkgQ6p17b8MRsSIVpDFjuE+SgcX
pHu6DdoAjHDd0kf1iYP8uQy1jwwb4vYsRIYz6zVEFRczrIwauxeHQyEv54aY0yj2YxM9kIkupwCh
j+inmwg0YGIf8ffIeM1uc/6bdyfGPX53KmnjFOu8/7qxkxzqiNRP708rLEcBj/0/WGnkYeFiXVIA
NNja8he7uRpucKFfPHJT0h7IKAfDRdN8fa/7jzjtgJ1k4TjoMo/y8Wz1mq3X8jx5xVGkdG9kY0O7
hLRolNcOMhVwNFf3yfB+KNL/b9S4R2D9zBYQYslHKIHDYGfK79AY7WbO791mvmFd0t9CSbhlxKfL
IBSPqIcshrhc+LgvhNK7SJRF1yoMM1ea3RDp6CpEF4i0OTwW4ZwEVhFKZFxMgUqlwQmy19rXIg9B
WglCbgN9XyzfGKDtSkM/OHrU+vEtd0xZ3ZKFvm/Qiv2TQcFssSpFPhAZpptNAN8wgF5fD6Ju66v3
rPraBm/zvR+9SWdLt27V5qWyszI36eoEabE6o3lv9VeoANgkLbx/IJ9VNTVjl+L9PPbsOo9hpQy0
qI2wFyJmyBVb8la3vg/83vX2eFVi+lqZWMxgZOOVNw/jsMe9WBqX3C0cZ1LZqxug2zsbnlpfRdsw
BRxEyG5EMvc5GBqWLYJCOI6uNZJgZG4JSqnVmkL9el3DB7lmDPxkTUzQsY8Bxqdl0rrKp4lsLuux
67JjKtOI/vToL0E/FJoM7q1U9uBT+QqvQxYJOfT9Yz4+X3s12rLNAuQ09pRhT0nRJJVf15dM9yrY
Uffc09IA61QsrO8h8WfktDtyu4EJ8Kik8gSsDwJUuIu7tiYsaZlp1cNTbsyqal447kDr4UAuQHDe
ITXxAZpz9u/yYQWeRnTBZ4Z6MtsHi8z5uuBXYsvyCJIua9x63HbElhntkilsTNeeJ92MxLTYGCTy
KHWJnphX5LGohQ8qW4nC7qbcjEEEBR0yyDfbXIAyf4o1rSHymfVOfJJCDC9gsMGsMPr/+ydFp4FF
iu9Bon8/hmmf+G1YRSQ6k1A58G0OCu5Jvwv5X8RbUXdZ1kADB/pSxnrj9mL8L9vRYqt1V8tzPcpz
lOzRbuidOA8gipivhJ28RfePL9g25hkBUzeFJFv1P0/3lAjnMwTYEvK/02GqdSUaScQmd2wpc28t
ANak0Aiau4fKqnwj6DOgTRjGM/4IPdwdBADT7H6oO8oDurxil5cDcuyukvDv4cBxArNyWj2kAr6b
CxAIK8iNpiaCwhVF3VcBLLImy8ncRf0df1Pdae+KP4gfMFyS65rL0T0cWyjuFtl8z1uKMoQODC+/
iUHmeoca6Z3mQjxBsxVTms+zerA7LnVqw2VlXr1XjM5D3TtlR/tuizIL/UVN2UusWUDil1x0sAuz
dCA78T3UvJmu+LFfwPa56is28SroW6bHVyY+8/ayIqUJMoCgZm99CqqpldfYje2N/CeiZhol1jm7
2w7c4jphO3saOvFv5a4G359JKxH2GACSqGL1tcBJvU7mE+siDMEmU4hxNsHfmPCrT99VUsA8CCht
YLP2yGiWUlRbgijk/OnfZ6weyeW3Iyedgv5x37nWrN9z129pzD11C9Q7fLSLiaq5QUMiqXGmSz8f
Zg2yoNBGNsH2yftxAIeCH9IZTiUetv9k1jpZT8/I0rLETCMhopURKoHQW0M7wZ7AdB9ANsVUjYYz
64TbQccQH11mQOJPpoMbVxkRtuBsvLYXX0epBRttCDvAE9Ynq8vACtZTgDtCmunZDYFmfNKwnEuM
7w1OwvSGTdTd2cPlF7Dc/faT+jT9pQbLPAZ6H/I69lZUsB2Kea8lGg80fmkwFN0ngTlMITOtWczJ
jF9jjn8CaaKxTt6Y4ErF0QMokk9S+ySy5RObGrs2bH421Nen1sviSRHheTrcPCxD4yQy8pgiGqIG
TAJYR+gkZKPAyAQbT3+jfEXIGOxyAHfe/nGn5+iBZs5gpv1uU75vjF5SxLLRoBKK500eVWEUxhXW
/qqhoKg/rd6w+r5tWzO99KBete5VwY4ZjNVDY3lCukmBhjbdkzMrdbn+LTQfjgFGkkldyUhAu8v4
oADNUmxmNEBqn2ASbpuxnYPNX119S6g4BWImYA6x8+vNXt8cu7MZhbXA5yZ+ZMXD+ztBBF9n21cZ
O7w9gTjdNDt6arGUJpOL86W87PdCf74Xr6RPvHB9PbQPEaDne+/TpMWOU6MKSlxkIwAZwYd5Q4S1
s08I1cHhM6KnqCxKmOLZ6HIh+/K1fEmyQGqTDTJ/1mXXUbQ8alm9TA/tuXJ/DqLTo+dOaDiJz81N
pw8tMXGNncR3Wsb516+ztoRm6MFPuxfCNfr7ducbbEu+pwqai2xZl8YODhqwRN998L++sprJRjrm
JfURU1RVrCJ6oLIYWohPKkue5K3YMGV7E6RLdBeFIPPo0vvieD8X3QOMK5d6i6C3DghjBUhnaDtZ
IfvpFURhziS/c2Lm+DUjhkKz3/1C3JynLdunluF+zSGWieLUukJJ8qmEwPJL6XZqWWEuBXJjvFg2
zVH4hcr1jVSw6KOED53ZPw+SXV3C4zRViFlwc2MpeautXBA5c0gdkdPPh+HaWw0mbzDLZ0p7Of0g
A0JU0QE0chC7jBHTWyXOfunw/UNRwoR5TKdwDNyGXJVAI1iVV03HuKNmaI43iUkQ/N9VFgJrWKtL
PGQvqJV3ug0v208qFM6AS0T/teWtVvIBK2KOjZWXHMK6tmNNoOa9zb1uMKwtdarYxXBIBl8gogeQ
stLpGyxA4GlgLYkb7+MyYAFIaOCTA51UJdYwJEfEp+KDf4hCZDZHzFp6zV1qSTQXUZtLoKVnQCnE
QKyN2CYtx/OQjO12n0Dd28e5CnSu587Hfr8PZQiDaQbpXXHyqs1HUlLbs50SbCAqYt1db8oKbGlp
l3bXPsaC68nALmKxaOHCcBPgR6NDqjHCAvNYYX//qf+ntjsX90o6Fph8W3uhNWIQWlZoSoJrXgPm
EpsNGRnxj93x4qWI0v5zjNq40y0LnV7rAxkaclINiPf0jFhT5skmgacyFEaUJRN+4SuZOaR8dZac
kBqrSKsOxE46YczXOuTCF2wujGkrhGvfmTpBq3YaC/frNrta5S6YMradWtrwy2G2cN7qMi2ZMWEN
dDpZ9zzIKzP2+xIzqHWlnY07b/SW/07fKEzkMy/7w60oefrPoaCaocoafp7mbeZ6GeI7O0Uspb3X
jS/p2jKRE1IxU/nlP80iEXwThWoo6e/WbMmKV510iH3nuTJ9RR+lrwZkCuRqwvqhwPBoF4w8KnOE
Q+aLQfWNE8tdDjuKJWfJ7loPKPx1+yzJmaXhMuChlykRC/+0ffgScCQeTlKUzmsj1OBiKw2ghFwX
1vbO89G20qsaL72uBi+SYCAxt9+UZYumZKXJp2Q4w60/r9JtPAKDWl0DMeIC/mXc08R3KjAkXgqO
rDRo3oNykMdmsWIEN21L33hIQXeaR9iYnhRSvGM1h6HXQfIuqG/im/xTblKUGhdFaABxe/quB/fv
9raSpSf7bB774Cw2FNIIJIApGlu6MrvhCfSfyyHkL7uBTY+a4KuwxD+Lzs66OMb6tXBTpURL/xuj
kQl6MNBoe2lYlLDMuGLB9Tfksu3NlzT9tv/f/VwyvnwOzsDDzpavZokzq0bnJE/3P+POMHQ2Xabn
bIvHCCGSKnOlm+dTU2uWRHKzMqWoB22hybBz6AN2zKXQ46t2nNecjpKAe4dub93y7jIRdELpNK4M
3yw5H52wRjoA3FdYqgSHHaH4/us+78+rhUMLT2kOQbkLtykgokosaL19cOh3eWUora3oETPfdxmx
K1LuzuxCE746C1J99RYj/g39FX4pnX8G/5zITyjvjfs5ikPTEGpa3SfWLcRFSvz7jmuotoMFfN7w
DfuvFG5K5EsSZB+OPDpekpH8UmMVyCeJaeydTw20XDBBNzxaAW2Ao/+NR4orGCzvWHCTgCGh7Fbl
/wzsDPJy5r5eOcb2GLIAtgd7CsMZSRj51s5nwxeQTeqEroTFn6wSwx+aPkNfND4tj0bzg4meWX43
lDjpSuMdD5+cGDJDcl/oYtxxVfFqLpz/ARlUimuGg1nDRyTBIDWE0IzyLf9clMe96Kvs5NWcD3+A
NJ+LE3ZM6+6x8aDlU06NtaXbmsC1vY0pFuhGnXyW9raw23sWQZUTAbF02z6iW2A3+hvzCJvnxPAF
9IYUYfIDa3ZUUZmKiW+hkrwGV6eS0NvpsKoNKswI44DKD3ikYnlToXfqdPpcaayKg6zSuZDnKTUP
5fR4EpO9oYLe2oG/N7Frssxg0N5yi56WYaWN+Js1tVsJUfqNgGvhleKgxQmQXBDn156RaP71Hcxd
eUEXftC0jShmrdjyqbYIw8n0N7IDUt36rMN78smMuvBJK5uBU1ogdijV/2qN1pcIUdVmQRlkAqCs
+JUVzwoJ574mmBWKVuT0zCuGcIzFzQ7cYCUF9vYkQuhu7KrwACR4Krwepy0pSDoyR/A71MXl89Zy
SATX1RO/KCsaPe5LDrudz6wVZ6NOhR6Z3+Ug1IZwwn2W0hqvKGwuhe2agXV8rWvfjIQWaS5CSdX/
e6eDTAlYiJiJ7sflELmAgbKVxQkyfKdx3wxGeuraZnTPZdW29v5qap8oFiE/Ba1gj3O6seUkqIBo
AOHJzsjXYCvUCYyvuWH67DTGH4ap6BIWv+jgGDHUv2FKTOUIj6hfC5vPUrmc5efm6i82jBY2hW7X
aZscOd/GX9tAnce0iZJ4K5NS1FDqjQ52qtcLXPxJ29H3JYe6Btq0upZKiqj3GQB0Oy9TEj6Cnu2e
lsUZkBExkKLu1kqJo0aEtZQEzQ873lL9mquYvfTxKC952s6xP1voZj7es8MfzH4KOeIIX9LU45pC
dc/OJVYT00oNuk6CCwjZHyhugYVB79jrhKI1aPGbQxxC0/EnFpReQ6HvZcJz9Up1lh8VFJcqaY65
ro2fpMGVN6MfJfioJkXdLApxOyzUm2g5M2l6N1V7GBYFhQW6KDnxC84YPan1+v9k87HbRoC6iTW6
FOVU0iFridpPCAK4QuuV5xpG3GYlKbLmYx6Wm00XCKYIXT1LIGw9lnhJvE5ZqaCyxWYQDlA4YL+v
/LTaNPkethfZedN5SadDFFjNrJoKstsR5tMaPBqMjnMyL+s1UHZMkzO4kr74LHo8O/1p8jQStjGf
lRMONwK2kKIwMxa1k9ZXqPPi/uhgAt6+I15lCjHFy/TniRx8aSHEuKDoYEvqvmjTQ7eolpkQ8aFI
MRfBkx8a2Qm5aLtCtAKhnf28qGOWTzc6eKADPZmGTQX6nUwLehpX+5OCYXVELUG9OuGbjKllj5f+
8Tr4+soF/FG3lpMTv1HlpKCl775KQcDxtqwkH4RELtNqE7a5msIaoFE5IVSWqonwhYDWIC9h5krH
PlDUI8RXsVPcvarPno4rjd2JTIT2zxKn5KNBFTLuogNivNIOLRoLZMwPOqB4xlFgxX4eeHrSzLUH
t2RLPLVRKZQN/UV7s0jEAx9836HuF/kui5aRweXubhTeYoBDOkA+vOyDEdTZIHqKMTce8Lx6VPiA
N4CdixZ2bpPFB3XsvfuFvr+Jw9BgfbM4E0ml02uF2N8ZZVIaNEivasaeJcSsI8eTxn+V/NG9KVhz
VlpUUR5WjRb3YsPrsE0KodJPugOJ4cvZtWtOHExhpRkzGt0zAS0qaFcPrC+wJ/0vo+DizG+n67qi
fWXPn57SBlv+g2gMVWJ1x9qMbUh52L8E/dfHOTQgL1qR0IRisjmZ/shbttgzp+h7qkJ5q9o5L83U
HWFjolUoJSZLqXeioqRIbQSSGaWnJxRxQURpawrhT5mvt5WQRYT6EkGq7wbUYDx4mVgqVTUv5UgR
bdqShsYtYXFEaPrEcppakBJW9j13UdiVsyDHey89bOFtD+4luPoDiozYE41fINbT1L4k0mI7iDBS
22Gmsz9XzKEp80nygnZeUmgoZ0kB8D+2vvBiKW1YiI1BTLkMzfAdlZXgDJONWIZbMOz8/7IBaDta
nBZeqcs97IEJfVpUkgnLNtHZbAd/uKODxLJJamA9vP0bMV2/GPjBddygkcC7CpDbJgJAVoAfP206
lLAtdj1hR+98jrinev5cdJO6a9YhuyBW5UjifN/HUv7aq87k/lHfOLbJP6MWY++/YOosEilbvwCv
wVT5CIeOYHckWejjnv8a6IbGNhRplG5wHh1erwbAGv0iLdBA8yw9KtW34lidWHAYq82v9rzVSvAx
BxXEmGlMdMPh/BVJPHPfoDy7b3SZ41hHY7ntat6Tql2IIR635WbxYoeaRT3yKFTyG1Wn4SsFjGiK
OvYbkHPOCiiyX7VdFztmHX9HIxIdDoGufLhzJcw2nmVRkXxR6zunVXi7UCAuFRjnit+29BsPxCxM
BZoDcwfQhu8p96RKagyQmvru37nhEqj87tmibz3YnZbmGkrkflWoYjob9aPW/zBqSdET+KbMcv7W
IogQl3kPGf0vTsqiLBEBDcklHFhIzczQexFlZeB9o26cvQTGXNTi4tj3VpaFG2U03QMxlS5nKZUQ
DY8g0H3ibkCatPWbN2Hkfprhhkm88Z1BLuI33cvJ3C2/4ZWIV4es/trrLNR2uVRrEBPv9xIcA7LB
FeuZSsYAAZ6GqRQigrlYQsfgChZKaNpJ2SI8gXbkJ4uv6ciZIoNDP7fmdNqk19hfjpO1eiBhMGzf
b2f2+VYgkCGbJgG1cx1KZRJ3ul/8JxDhS5odLrxRdoBJjFGC+eyKBzRelam1NT+EArzgYT9qmOxK
jK+UKTBBoTpllkqeEhZELd1dBOg8q8zIxhHFeAUWBO1GwlZwdwH4s+EOnGHoGDV/ijgz97FPmBrd
/V/4blVIlxNPOfR4NfY1Bk+S6WlOyN0+2snyTqHlrhYbQsuKq2fL0Iq2OsAJemh71xYYjp4+FIXt
CPNQeeaRd8dZPeg7SXze0v/iOw9/WwHBeCO26kL3nQ4GcjOmeLsMlOWEqQkPSia6CkRsRWyzUiWV
0ah1sLxfRb/ERN5MSlyF0HeDuIyySBbk4wVXjIx8Sg7Zgin504NhWnmmZqZQzfrII0sriR21twSR
xjKrv5o46zZ7YuwMOAZj5+ijFGBWujm4P+hVWi2dWmcXRRQbMeO2dR2bBQpJdXC6UaYxYa0N+eL+
hChF6cSkH8MeCbwmktfbLIzRaqjMnFx4nMdHdunN+5dZFO/gLVmZUfu5W7ZUj51PpNWtbYHMkrQK
Sla3UOR0LozR7uJrOUI5FHBeLD38Oaodar9NrLizfKGUu9FLvWBNCRFb/WYKEhe+v0juEqeyUfzF
alYWL74zFK54uAbXx7Z+lTDKPVUupXHCUcJX3varlkoMr/rqsyIFI+fBD/T3yaKDUWbexq83oPDg
U/QwY7ZtGqJr0chzEKvXmRjWmBDqSkBk8d/nAcC0QLpcq9AJL5QycJwq5BrfWtDhQ984QjjTEFKU
Isc5/lJG3wRgCvnAMwTl+lSBg2WFIJeMH7PjnYWwVT2Ea2vae2cd0ea2R6qAEWavdqfmiOwnxLDd
jo+dfPr/vmLR43MlI6Yzljz6mOPdqcmRJ34oqcieGjr6qumT17QdQzj4dAtrj33Ei+0wFoEtrPXv
vAezzgUph8UT60HXJjWl5r67p7dKMGdsdekLp0POJIpLfPopc4ywIl3yTauQXl7SEeM5AmvZsIXi
bHdGzPriszujPnWhB4ORkDXBGIZ4gYLx6Uf/jAJ/XnQHNTSc/u0DOht7nuoGuPDSgj/KfM//mp7w
dNyVrQVeuKUR1s1cBlWfsSaMmsx7i7TT6hyM+9UsGCWJwwyCmKiV8HU6wN964BJISZ8b/xjJhbUs
Re7ZIzqzcCa3NjtQwv5IOtbJJmEF6ScE2zMlBrncOeVWr8W1NxeK8xrx1YJaTUZZF9YbSNHRoa+c
fyr03TRyn9mLqAiPKcrPI7B++XVweiwSBKRAlE37PNc7L4RKWQWgs/0VPGrbkuuc078V/C9Op/id
jPX1gRr+yTSa1uy/pzGUsGaLZELaxBsEGNfSdZ3w8rDLNnHDpqxKbcyQC1iVb+xLC1cj+puS4nkf
dFmpoA86/hUsYn5dTyCTZed6XFLngPHNlrQTX3rr/+ovRfVeC4ZsATHebP7c8wdHquWdj+11OmAx
A0ZUMrtg1POKc7OIgaXx9rvUkHbw1+NHFNJKPhOFw2BT5x+zNwpEg8NFzxeHyx6XPPQ2019bc9EY
9w0e6VcVdsq77m8qMELDIsRjNt+0xeuOLP8W8zm0GbLvWls6/ek92/CwGdEh0cNsEDwpyr2MqmmM
ZsxjXkbHOTOofsfF5JK0IyxHqmej9SxyMSy/Tw+MP4BNG5SiPzuy73sJw/6ild6t311ZZ/OJ2VCn
b3+6+FBlOWtdu2lhELFYT/Uq8VWTUfOEYWsNNA5bmctKfTn64HAB2izndygxW9LE7NiL7mO/xLHr
gUicf1t+BjbFZyWC9xfvKCHaqxtD3d09wwitygTXsASlPO5+eW9d6+cGLOuhtm4FXmtafaCN+9LJ
5Q1Dw54kasYXnOIZawLmudebZVlKj9K0EWyCp4yQg9n9a+Motvq/RD/PPJ/hJf/HtH6jOR4wnAwU
nCA//ejqmB31N26kJ3RZN3gMpGJgYknCLxYI8bHKQi4QHTPMEmW2DMizX2Q3N2h759VPJeS2ZPNJ
6CLr6syYw9GcrgZnZhq4ROAeBmQRSvLDraWrCAeeuTbBRLDLJ/aB0T0OyWikRDAE23glwMy/Zl7T
tzyPxx3UL1xRS7PlvmghJV7cC49R0Ce83s1yPjFvJ4H14ZONvqaIX1CaL27WjZId76ngDlYXeLsg
SHrugtknAdkKSXLhV2NcqlUSrTqIZuW6DLk4ET/NoszYP39Dxiw2+bTECRTnVz6RAZ3kHAg7WWnn
wCL7JqvKEQvWuPQJlv1W4+EXLSFE0i/yGDC0hLJpHBdlW3fU9kcGo5vXkJeButVqz3VWl/1FA+LN
47l35f65js+RANrwGa/gysPhUqu9LlMFwZ/PlhLjbqLGh0m6wZekfMSk58HtaQvXEAApqqEkmTWf
0UWSwY6iTYPmOI5YegBRob/jtwNVfLzFlYjSsAPOBKTZz+dz0iakY/AKTiD2+W1XjkFpWuX/bjsl
FVurRR56HcCgudqF/ULfRhW6gn5ZwP3PGM9Vx2yqAoxYvjHKy4k5TdwJU0PafLgo7KrNBf0OqrYo
wVrgxs8SN0L9CMvp11yiMWjsdSY7tX8u+ZGcjGFQ14JIU8YGaSRVLtvKfifJ3IfdXMxzzhU2v7hZ
ezF5ASRugazufwmEE0UOIjBzqY27RnQReQAPgZWRdlkG4DgJlYXPOFrLD+AUxfhvNf3B+Vpke04B
je+oR4A/YGJJRTjswAQ1YQo9WHWA3r4RFk1hwKNZW617bA7DcU0WaTrOZpB97SW2Ae/RlFiExOS3
8ei3kl7BH1ZmlpWizqPUDMVHp9XG9ptVNIVczoLhjKDrHAlLRcqMdwgrnz//Qg6Yib32TW22r3sL
ipsi79RLVnNLzhliwE/vQQEEqdDTapBmUc/SIFNKxY0q8HFvNeFkQD1efv2uVd9LZkUTuyTCA3Im
uhZs6ceJ+q9ZWl1h0h0CmXLSCyWNIWUiC54TrPLLcxwnP2dOTCgF6XbzXVdLBnPgziTUlHXBCKAO
RSYBgb7Rr4bH9LaDWSmNWmXJr3cyebclJcaGe8j/BeWJoKI/2U0IZ33d9VdDDkctWgEDjaJBp1a2
n4HDhdnuJhKZUdnFbNimvM+hEgMQigpP7uXQ/OFUBlbzrkjxCQCgheszby4pxazMHbk4L9zd8Xxj
ChiifavQvYi4+Sfr4yl+geQ33d4Wo9cxPmNCL5I2IZEF4+V4AVWI3B4CjjyydiknveuEzS+vctZm
An2ofdYagNcVA8uDvmpJtpH8zMMztXXF2TGLPfAKFmC4b/kTAs88+wJxRNY6LIrYoavhzQnV8n5c
xNHWzvznF2sXDAd3+AAhXd27JtMeWu37/V432BK1TXkz5i+mMF4J+ecNQTcqPAI/c+HbZMRpUw8/
/zj2cjcLhYzf0kfcienzspVCDs5Y5R5GO9HQF2mCM/Es0uC63E9DebDEgrOq0mrGlIm5BM8B0Ulp
f/ppM/AIYU43nJpkl3JUdCdRZNu8NdQ7Msc7A3nekUAsqggg4Cku07Ymg2qfrM8sxZQWoT/3WED0
I8F3dq7kPiZpe1Vd5CuB3CflSqEphkvk5v3mCvooUG9Gs73iqgicXNku9p+IZ/7lQN/JRUdq1C14
p/KqiGqe0pfgzjLI6EuMTLMC09rvKgrAeuPRemPnq2ea3DBLAZ2TxVKAbSjuG1V2DbIQ3W7TGi5e
9Ahf7Da6ihGIepOr4PhBH4dgmrNc8oYOzLehwFAGH4cVVbAPUV5G4WcFZFFD5w4whHxAcx88rSdX
L8/AxviaiHGKk2ujNHei4RMaPFuGeE4VDpWItunAKuhTlyB2Vfxzevrd3+ZmT+mRea9TZw9ZQMFE
XHPdpeJ3VfIrTXjciuFEeMj7SMH3fZIg2pI9KHnLL7iBAG74zy3xBx/2QOBTP/uN7M65VVTQMhKZ
HypCSq41HdkmDuNkKf4uBhW8sc3EAjEbkcNaE63TZRvQaMxw3yJIZzHxOgfcWA3PzKOx5+zpMDqW
XiDOEnbLe0FK44EbaFqFsDkCsl30Fjp3JYqCVU/KZKno3JjcqgfMqrRLUl9mGLYRYoRAvoRQm2d2
IX0Hm9NIPRnVkvE6PbEeE+LjmeeemhgCs9LdU7ib7hqPQXUo4vrp+c5orpSHv3Oy1ADFd9wypV8G
yDF9soCg/kptgtNVokTQEUsRiuM4hL5c4KDfG22Nvt/qtfstVKNh1g7Lj6KAnAV9Uf+A2EuGWcct
lstMPDFD7XqX7BpKp0MYeA7dH5qeoJfffXNtdEqAP815nKPS4HI5EGlUe7RF5I2zQsK3t5wps09j
k4JkVsINmFa2ba3MvLzk97Jj5wTz2+5btsXcXSI94Ibp6zjSJ0hsNWeuNOrOhpNmN9d53kx8pcYe
rzN6d79hzTRuV6u/UO6NaMX0pI7kuKdVtIqG3LBipqwtSW/fZobYp6lKXBkyPy557LfmDHMSabgW
e2VIgRotmBY01fEhzSqKAkZRBnn78krxHwXitBSaQKAPW+BhrAxEZ8WeTMjqTCO4NkhN/6k2ghyv
Vpo9NNJWwNLzseJO6Viasw97nGmpWeNp1/4K/4f1sgFxs90rM+urOENEE6yI8OzYIXoNLXoW2rqe
7A108kVlQLErhmLlqcLDSjEYDLPfKV08Uq3Gh/NLK9tdiycVRA1ucOyJLM1deUecbQZP4l9KhdvK
//epR9tAOW9YA6gTkSpNMtTGJS8EgjUj6AFSA+ht9X0O/NNy6WVVu+J1Ktyrm+T8TmOXnYWCdFOz
O0FcFuQnLacvKLsx076IT0qcDj4juGreU2SNFA//xRzVjb8aPUU3Wzqe25cdbuTsDHjRF60UfYIz
T7QZpebsxuIYDENsrlKcZ5VNIP38e6Y+f78gwF6hRtEahk+PC3ELpPayMvP3zKgo7ZFip5E3tiLt
daDRhjMQWYlfKOGDW3jvEGZAsD9P+K7TeqwjJw5JBJgpDEvl2OvXuCBiTcr9z5kSGNDyrDWyd9ah
AvSEpoM8/gs+LtjnvsIF6J2yEAnZ/9wyADGbyAQRvw5Zom8pgRlsjCut2HwRgCR13kFaABXAx7v4
zAE4v1HDwJKYdaPXDnme6mXeU3GerdcwAGwCu5cudbs9idiEAcLplfapKkRDmVBrngGTN/4prc9W
z1QWTDyiHVRk1O93WhZCbnmAT7I+JA3s5gwsxqF/CEjpVT/OzAAXBZTT54bGjyKIczfbI3Km7q9q
gsekOasgb6iTb1zWSYkEwNQ4/vvw5H0jdd/NlwSF/eNkoC7dk4QDe/dVV5zAkiuH9Obe0Pk3vQ8G
+73ZrMBSkw6LQ44Vph+2+DYuXo3wwUM52kE/+ccWajbynPpucsAgTzcJcQYZykX5RGRiR7/XNerT
PGzL9JgSNNUkIzOds9Pws/8/x3DV+l9BbyuPNqWluJAsAhRGU32M+WyyP7EYiJUOJCggoAyzv+sc
mzuZJ1vqkmWO1hasOCel07NL/JfxXwhNrT+c3p6+P7cHyr1A5ksuZvJplHiD+sfCCIk9Ov3nSaze
r7RPNr/ZNXD3ZNytR2RJqTFZR2xKi8lxcgWjHRaOUSaaQj5YORzLCYTaTZYFHqrEAu8Umo/yesuq
rkwDzxkRRObXCEuNlBubhaxUSXlkeoQ0t5r7g4M48KYa8m6VUiqhdJ0naqTu92JRNk4nAeWNuMov
OwrGcefDGzhPfYlrkoZP1vaFDU5SnmaTuC5gKRuo8BtH8hRGY3hKRowiNCXHWsgPmQZ2YvRpB36v
uGyqQ0/eKjApsJ+GWXNToJTGe9/0JAp1Lg6t2U3wx8xx72Nf9ScAyjKgQEwiB4oTd3cbMMq5bNA4
AF4e/+y5CVIDobikOMXnLBTeEz+SGwJ2egbG1pNUMyjXLl3SLwDpZs99RgV0RoHJCbjDwDXA6TbM
WH73zo3X1+XVodTtQDRx0Gw28tBHGviHt7scLEBt+ymfKDFgoUXmsV6RDYz1y+UDIWZDJVNoCpv4
/ESc83KzMUhxE8bW+Lqoxsz/flBfxpsKvJZghDErLNJbiIApXAjsLQRIGykftKSd/hBPHLv/a7Bb
+5aphSgv3aIfEGyyonpybzW0jkesKoqU5JIW3wKSRdEKkOLjSor5jOLtvwUN2RCPJbGZoeuhwVXH
TPxFJXayPiZigYY+8t1iOAD0dx5RgKWXZ5ZXw09mLwGIhI9qVaNoN3c8EqYAq/PW+og0fuVL1+Ms
t0f4k2rB+eU255sDUXkxmzCgLf3nQsyPKi5ZlTjTM+6W6UUX9pMfnUMhaHoQdInOREr63tboVLpI
s6mvu2zMrc1q4ClEPNeA/nAxSHNBDK9vq4VgheNZABOVW3qDEL16I3y/VIJFGFUBSMTsL4hWuEJY
AyKo9HPJPE/JPQpkQV/Ss+Q3ELzalAeEEKEoGKBDMv2OaqEz8FsIdxiK0G93BMtYgtD2o+940Vp0
soLuqSEwwFz4CuO2KD8/zqMhnPJZ56mPHbvmyC3yJE6RA9bbT6NsgIwkuegn7lx5rriqyVNqxCbM
u1gJ9TE/6Gn6xqMxIYoijsH4eBXZNEQQDGRWCXMTpl8gKCnsyZler+ZKnm0PFe0TqSZg+brSnII2
QK2EIqitiEaUXuNEfmDFRN+I2wW03qg6TaTn6Rqk5wz1t40tACBZtOy8xFRr+4rgkeVOb7ytZT1z
eRCh6rxxRN4JIF5gcGNaUmpmj8TtkvZFaeiYo2BqAnufCpK4TWe1GPxaC+e11lyet5q8XAVut+zk
Np4k7z0ufgXSoTqbB7GpjjbeL+Tk29UxmxGqH5asddKRvCNgI4Y4gfiZICohz1SeRoNb6BRx9y+x
umEu4gEV1fwiRHLWhr6D8+6zPqwGDB3QtHgxTu/K2oHjvdxG5RkzxMwK7YNLV17UyiHSElBq0YEB
Ijbzi5b2HDMN2tXwmMqH+zpkjQslkViBEXAhlffPoiWG1xae6m33CtnbuAFJUS2McLbKCGFw4V5w
93QZLNvF1Wg6WZ5btopxC/ETmpWlX8sFgZyNRag+FIxidmKoV0O7CbEEF/S/AiyH3yAjYSwqrPS1
f7a5LYilOXbc3x3nS+6oh+lhygj9JWFEiZPAvW1J6Ec4GeoXtgQ1n6GyjlMEBp15OAmaPJ73VoWv
9TCQqem7VBBPuJRqyMbrbQ2u9cATHA12jKGnon/Ni29oNzYSeyaHo8kI8djoyYA3A64HNNeiqIiY
GGYUgxd+635S7OHVTrusAza+uUQiy3p/+IkuyznTO4I5E+D6JBJMdgFm9RxkezUJBWYscKAAZf95
SNTTFmG7B1S0089YwEjjdqeCAUNRVEX6lHsIIwr4OprlLeBa+HtNz/5DuHiy7icCEciZU3oLHfaM
/0DTFHiilgBCnBlRKDEp6B8QyZEem/oQiTIuiMfW8yRzbhAyqP9LoQrOy4SS5Nu+MLsxUnulJFBd
r1Yni8/8qDaOSICYrF3ZRryI2lOXs5cOp52FGm1GT0OCKiho/xFHt+tSmSlB/qRGV15WSrWh+qZm
UsMjyNKE2TLJULZ3U6VHIc+e0iDitkd8q4CNOyRH06DZETEFuJnS8QJHvQSmK09scs3xE4j72MQa
lc+Ht73PoZ7VrBvZE0Wph/ivxAX8bSIui9hgb2k24jpIQozl16wN3Tg6FUveHuXIYPiVn+nD/Zjw
itNu3X1rdo3QbiUCzULGbIFXETTTp5IzmHQiZGezQSIFEAds/ACsCvmc/aTa3R2HQ/tE/d6WvYyl
YBgqvfKJr9HIobSoo94n0lJmpeQxkpmqavBy/kAvYU56FYfYq1S+iLbar9izQlEEMHN76UK5nv1i
I7uHkqKkQerbYKmBuABkn5q10o1IQHcKhjR2up/FrZb7RdvRq8lGVspyXSrwSixI0/rOpi1V2k6K
YS3VMYQa2HE2n4bkkVcxSZV3NowS218NpYN352B1AdfeAb0YuvpNz1DgA3u3HoX6Se0uekz0SAft
c577bGuHPjhrpzMLpchXLIAZENxJv9q7U/AXHL+nQeOPzPw3XKAYUmBdcaN12VnbDF6NJQawoHCk
WvcQHBNCYp45SUZ5UdzpHYdIh2iZv4Fig9HqawlV1ajJPQ6bs6hE6BzIwTwxs4QknX3uSegQ8nTn
7xWz5q5s9MATFfOAKBLnZ6wSb2IYcXh7T+i/ar4FhyG2ejbyXatDY67NupGe115a/c1fUNOMJ9o3
DIwKsFv0IG9Xpa+72L7Hgzh3W3Kbgv7lOVNQ+bjzsTb2u2zRn7c8rllXYSlhv3qJgH8BagMk4K/Q
46YWjVXt3P6XRhgq4+AC2jmP71jA0Ss1Aqu9pnn0UDp10CCSK+hVBvpjogOxd1LdXFpmtqoHvjXB
cV6yEzAwRH2urkeYbJjfexyATG0Ve5b2R9GOVJjz5QRt283y2zaqLjUY4JbJmYfxv+/QX3uofwfN
VZ/BJQ/HfrYxD69JLR/D9O4ApSJaNDypirfNFQyFtBrmq+TeRU3EeMvzmjqXsamHyP1BFtZEXqXt
21WGip65ceLB0O/Tr9wFQp1WyhVLB5j+7PaWBpNfueoaJ8VUYgRZDO8kAxoiqKHPRxN1Q3l8xJq+
6d1rLmOwvYhEu/G/GTX8Ukr9YZiKek/ZoTdG/+lNz8RPu3dPh+DfS6pj/mLlLE/MY7XfMyD15nC1
ZSvqm6iu40JUPY4cSp44G1ThPIIZuhh7vbJJGGKRFVFWNKOedjBRAejVxzvzujRdcUqmfN0Nh8EW
9v7tYmMDts7Gl3aOhwGkeOQizcla429Q37mUa3DZlwQzbR7/uzKJt9yhDc5UpCIHrBEemlqrLKqn
OIvZ7+WtDIALiRqbbfFe4uPfRDYDIvEVute65GM8avUpAurLxgWVrw5W9sZPqKNQR+Ax1cAwqLOU
tjAGc23LFfl3H71vw/hXjw6/c/Dz/MPQmZDglM42bDe0gsO3sTG4HyZTT+3e629eJoNec19DHENM
hE0bKWbXzm1bJ+L7jKI9aC6AQrTtV5pLfDYrst1i7p6bqhSFBbw52ChYiPdEwZWs/oEW2czax7wZ
YaG47yUKycZJfcElpV+hNocTHzX9fvRFx9Jcv9SGx3g+fayA2alM7cme11Sj+KGMnVOblujukdpG
5KbdhhMHwdQsoXFuCZtryA/bEcLtL9FuZGEyUezVCqDQab+vzxdPnyKRjcNvNVDUx0F3SXkboa9o
NLG+xqTo3WFqjoFs+ymVRS7/i3fvI9ZNlVeKU8bnP5hoZpMnm201m/srZykLNrdNhDCr+ZhOz/x6
eTkf3h9CzVux6xr/Qhw/fQyKezrmMnVgz9b8IzLM0v2ow9nNr6nd9kpkiN7CvFg8P5xsgWwc0K0F
QsHbuYvc/Wq2dIuocXYMnbxHLlFOeE77EP6w5uwEm135sOdGz40ZROQWbn1f8l8wa2lJcOVhMirF
dVxzvfKkd87C+yubyYgbAcQ/UrKSYnZKP0FEzJxnnCqnKG0hElynDnUc1u9IuLR/szexXwpR2be/
oupl6vvu85dPli1v8To/BFjcsOiYXEE13lBqyASyHNE+XDGN2ajmcP9MNANHE61eU07ZsCStxkD0
vgPl/DHdyyPKDWKBzjQUSNgx/OgUancEOWKAoCIkGVDuafyWydlCA9H/6BJEEsjEFyrk7Avd4swo
6NooRuOZMSyPHkIFAIutdh8ohf7qySnNusv9u9+8hWxAy7EAu4yQKa2qR2C4edM2L/CxbG6EQH60
bPs/YERYpwHAINj8RhdL0TfGk3skfVh9bFfBUV/Y+O1zHIFsfTRiIjoLcDh5mp3CyxKCM/sdFJcL
0DHzO9YpfUOiIoND6+2B2MPi1PJFUS7U4nkP+bJk9AEjMrCm6uWZKLelp8wPKHTGohFsUyGMROH8
+5chMCDwTosUIMKa2MjHdYhzNPGZtKbo8MJ8+s1oriRVZRk8lnitdiNT8FZ4EO5tzzEiPW/Co4As
xm0zS52FdcOk3ZOsKQ64haQ6nlEeX7PDG3l3BJy+PupSXhkgtFUM7TYzu6gDCubV/KcJFN8K1RTg
qvrQ/b1lkQFqYU7Um1lYI3uqjZMR88cDRxfyOf9rYsaBxU/VxsROEeV+dZqEPckhHz8WwsDiDwRB
ja2Wcw8py7Ka9Olzah+qmY2AsxRbwzY9q2CmRpnNbIZStCnkpRJQ8EpX7dmnatpkleW7oKaSVPNH
o1mLylJzwRbub/QsGsg8q/wGchT5gCj/Uf0u+Ews9SnTBXQPcl9if5qcXkEF4E9WRcczBF82dCt0
fSrHpA0c2Ms64uAEnMDzlwRLwhcqeE7C+9fBNuG/Lxh8OLz7GRwoXEBjjMlfGpR975O69KWY/TFP
YZt2i8DKYenbvz6zthkwI/d4XnptkwytTgLhWJZB98CJUhAm99W/7tmDBnzG9tT2rEfnTNmIWTiM
uxR+nPwusPSZee/WwLKOTK4+UQ/Ffwb56XbiapTquk3pom4eT8Yjkug48JANErw363m0LWrziD6D
JxB/RDYfx9cQ4tiVSEAuwLHyHSWjVUirXXRYuqUyHAeKMb13rUSpuY/kyht5O4wXPGsmqOVqOJ1M
wKn+0tr6DotNH1skfDwpqJ1PtWOKnFvK5LpEAanEWWEX3KUtHIPeu4fop6C/vaPcPCANc9eJ5LCa
CabUtNUotn+NkhB6lx1+y2jqron3UhVWw4P7XOBUzvSW5tN+Teg5RPY5KAsAZfbAjnkhWf/Zv9EW
DKu716BSUgLBKgg/yWipit/Z+DA60MaGvhLBqSsYEw1dtHxeB3B5sKNj0t/EN3JoU67CVzbp6fgj
cFlgJFqKWPCqeRnCz1nBXpr0GHOxfJWZjcM/BBJnPDg7PXaXhOwf8FgMtk89ByQrhP9N+mxxL5/C
bmiSIFA/n/kZy1sKa6boj3K4ReFOzvEt7RKsR3zx6gvs7aDf1L6PERAJy39Z/l8BP6gPKgS5tdHz
cUHgcQ/ckeY/CE1+e36IdkqPdG+rv2m9EeThJAAOo4zumytqpAFZzM3IZXtN+kkQU28PrHpfXLjK
dJWcvcTHi9VgFM2ked8PLFxxnRbjnH0hnGUdJ/6Vb3IZmnnnzHUHqdCQV2jJXt/0g3kbvEsjTGP5
kMOFyt5fDR4aA3iA10dfhGfrXz5t3bdr9chZ4NcmkxumR/mZNr7Z9DMXzpRKCE7qA/Ld4F7KIWLP
h2qMow49DcSgFB5AUm8sJvRD5CFMw9HdSiKo/kLSiMVznMWVXFvr3j2ExbuZqra2gi1s6JKcu42G
43Ds9onrMVF53cnlPU7XIm3JUKvmhLFlJxqzQIgSQE157qDVI3uUiLFUrgjEhoW+5XtuGvBpewZH
LJExSDCgpkGpJUKryIsYdpKCiJvRpu9EngKkFhEAQV4uPyMrejdrvJLUnH4zdoy/K5DbXlaSOg9w
5u7WvGHx4Ke/VrgQFVqkUfJfcSE41zdL1Boc2raQkdVYGGkE54TDIsBVgDNL8o4WVSHcO/LNVquE
t5lE3KMH8mzkRgy7jcEzTU/SyvIjXz0kmNve4e+o6Mq/loUfTY3fXGsJsSOMFMNAFiuwIyeYKszH
TATRErpHGlW/48MnWu+zGHArP5FufiY9f6NeJiS2FeqV/XGFNkfmOELaOMC4fsFFjZGm+FmwF3WH
63POQQkc0enV0Wkh6orqvYGgs5aJEkM7ARYdyDqwboU0oJ4KIS5yjJtv8odFvAVHFSJLFC6Cp8Bj
4vCNCBF/7e+YeUIJUPZg4xgYX6yYEulNc8r74K13cvifbE7vDzeyB1vF/ZT8EQE/6bR/Tg5VconQ
jYej8O/8MWMY0QMc+EoCB99xfR9TpPxxpn2Vpx8xE24mL1Xbv2Jt2O5doLFBthEVirhI/+Xl/6wt
QNFT3DLhD7efqbEDH7eRucaVGtAHQKVGgyoDFPkqhdpDS328pMFe9wmJIc0kUvAKQ9AfJ90IyrRX
3GFRtcAOkRTVFBoCb8g79zJopiKZqwPZ4PxQG1G28Fb7sGnWow2IiKQhOJa13ZwUJjCFd5hkcyCK
Y0WUfeu547A/FLpzWTTfNO1XP+qYborRoG6a5ljh214vFcdx8ikdC7e8CIdvm4wU8NHChc/etXJK
rEcpOz0Km232tDlW09+O+RVCIos/jsJ3+i4LT7LEka46UJH4hx1g5ZXFkawelEKZUTLM3OcWgqpC
i2K+csuqctrKzmspZZ+h8d8/2XCCHRT0Iu4LWszEoJyxsrSJd6FkAeVlRDq0PURiBorHdqB9ABmM
06NvW1amz82sPaSNBE3fL3ezPFe8tpfym4TyeNkoazu4qWgVXOqgGvSBrVSaXeWvbUi1piZ5ypZe
WjGJeq4wQVcVhGdABqzVxMQ0VEOCgiNnXnBjC5Oa5KwSPql0niY1LRqXxS5+s7TI4A3pwKXYPdb3
nAgndZhjYGG9CqgIsbmtT+tD17fwoZ/m3xYJ+g1RyYEit0m3o9XgJtp3rH3l/KY9Sl2e7lG9lxMd
sUBfVt8lgGZWExO/ozjgcLJwYtjfvfmfYMA0GeAkv7BTVX7NWz0vWFHHiiEu3CFxprQuRZdZhrDq
7G5hoe1qJeROUPm7pxCbIZNwaqq0kP+NUJf59npsJaG8hRLeLxIxdSjePeDyCFjMwz1ad6PGI9lE
S5tBLH+R17NS2ltLyTW3pfYV2hahxt+ioK5AbgUf8CQmFPCibPaqSDbh7XeR6jv/e+kXNchbeSU2
iolC1o0mgaTuO8r8AE0VHDA3GIGqO4zXAkx/AropdgjLQO+8V2i6yOpNleHhPHyq4q4IyeYyK1yt
Pwosib7eqnhDzpib71sBTw6J3EeXkc7r6kEpI0pvSos7vnBusxKXysbKfdBWqRfAVzojNA8kJe72
WON46ndIbfHYP+WuZT7EseEb+Iuxd7puMpQCr3MCU8QsF5Xnx1jkVEdxv5r/i+2w0+KwFP/vPB/P
lxB6YHOUb22yGHtkV5brL3AO4Hg+s9aSdbELjb8gSk52BS2r4HgrzgM4YpUGJAJYwxafpuCUG0LT
toaqj8sl4OoLTr/AuSdzk+v9aGWfk2CrvJPnmZlHkahgJIXmyX4+dfA0ggE8P8mH9XuCDX587jSK
cWDQcB+HwTGlFlt1RncZ3FaBMVIkp1DXpyyaoc/18wqp33pwCaV4RsR9ZsISzeiIGjM6uV2ZpAK5
SeDcMuUpt/HXM8KIaSl09da6VxWZZ+YJwP9DZv6M32+ow7btq8qrbj/a2XMFJSFJ0aFZ1qJAtTAj
lflAmtpBi3wknDJZhe2WbXNtkwDdnrvfGQ/XDPPX3Sm4iqdz9050KFENrZ1J7Gif8a8+DIIAbnHf
K8+QibsQ9SONfuYH0st08kbxtcmw4fL7GLdVU8VPEKGBHGiNgwYL0RHY/VkDItnG+VqeyRr3C9dI
eDnVL9qQDeD3VRuFe8mzrzt/lXTmrVy0/FF9t5apguntURKsM1+nu8MASWaRB9/RRIqpwUnsqliG
FOWLomBWzmsqJzAdgM4g5a2aHDIbzuw73AwQIbqcayxZPrP/CcT0nnxmCaUCFtJD8N102xH0SOpt
48nx7p6SUgM9BudrCTeZ7O2N/w58xNZt5ATbqZR7mdxLz0LGtE2M2mE4GZ0JOtXfC5m4fsPRDlcv
Df3TlSS8n35DgtcUOp1+ukw/4OLhvFovbrWJTIC3XDFLQxm3U5jSC1/SFEmd2l8Epcm2DDy8j6Td
1LUzZkUdtGThDHd5L15uX4mio8Bj106YKmn/bL5tTPfwkz1wD6dYJLmV8g3eSzg002jIrWrKvtKS
sTYqpwltrfn48i1ZwuY/OlThUZtod0uxyFIf+Lt4+iMZ4rniAgc1Omziyd3+ubs+wDKd9DvB5gBv
qsB+f2sBKWlXq1uhObsb8H7aD3m3VZmcTVlJXtSUB/nFxmR2RSpTRYbgmlYOwGp8AcOvEYsf1IEB
jqSojB3hb7spJpeaRa1hPRRCYBe24S/uTn1AhMBKVQT8joUdqCfpar8AKCfXoGEeek6KYO1NA9vV
7n7L/clgABcOogRU4PYMfcZ2McCqw9S8XVugRq58cz2eigdDUYGEGyeTzvhNgka4s1m48nqLpB7t
wGElGxPY96FZvw3cIQnZedImCLjs5ltdXMGyZbjLJH/Yq2GR1/MBYttpP4A1rRfB569vVDrpTHJ0
ttT/4P1kKdFK0p7X7gpjnMLr732XNhiZ761RB5Ym2JpLE6YMPyoS1uGYQoFr7Geb5lS015KvPmoG
c/Y6ba35XljJH+XYZckZYHlj1FEfivSOuZ+HlXGCn/SD6QIGD/Fi/eLK5YUVAAH4iZqfVRg6Oy/M
FDLzuuMT97HVku0PKjwKMkTNuXdiMRMMHu7QJbx5aN3StbK1fs+Lrx//OZHpAChMf1BaSHQQ+3u/
gr9kn2cKFOsXsKsSgtm1YDncpLQ7jy0rMnpNExuBrQjy59g9amJ90CCY1vywqYUw3xBXfpvCuSC3
mC+Gv8h+/U4OxnVZhVwEIGzF9eY5UPMoEnSnKi3Bum6MB8jUgN/f41k8RpN3Q9T64u1Z+OsTchX8
d6jCwRK8fiGRkMpCfSiNQHJQo3jxapaGM/k2iVEFTQo/NNpjmosc/eZTXl4eyhrMTQMAw1hEZ1dS
6BVDM8YbK5LveUIg+91muPI8rZUDfrc73KQuIgiT9nVVnJ2U6XXnx9IDeWsO7jYz8lNmMl/tTTzn
f3ErjA8aJyG9YPr3dXGSPvS6IeqrkN3mAod29k8VFtL4JJNyqqkUo1iaI6LMWVjh5F++ZeB38lRv
VDowz7CQmqWQOcAafB2aLq+fQiQTDNkkZkrK8S3QLmDhVJyMnuwgXWf4uLS95Yb2kQ3WlNnlPGt0
6FHxAMAGWCG5TibnYFefw4/T+3AAcMuAa/1x3yl1ToSytSXIR+D59neiQaUqQskf1QHUpttyS8LX
6ztQkBLWcHqp9MimK4lON2AriO2zUhWlnCOjVHND7TKc1AUYYouSOyT4cObuOYYgvJhIlx/ziUaN
VSzrGxYoWYy8/CdgpavUuCn5t8tXbjanG56HPIr+w5P0NLesrV/pxSykhwoa0VIN2oRcD6TFGV5O
Pmh/ncis5sCS+v0Ldbi6fTYbqEyoHtQs3U93+HxTLHsmLoyF6fTsN+xT+HSpPKZ3E5N/xWcINjVh
pB+ViODrEZW0NYJbNZa8EANAWoxFtW/DdQU61Oul2UcaxCFIjjm2zybDLQdbPKGxdyjJng1+NRNa
HUzwS1x5pVEmQqZ0wzQXtouDotllnMTJP2SN0JNBP/F6beApur/XUazu/FIMb+sDKdo1pMFKAT1z
73xc47wUEMuDF0GXLuOBfsQcsBZrgMqaqglOROxlrtZLZaFNe2Rx+TZlPOSVSGQF3wyec6Q20MGF
ByC3p8lS/Su5R6mEBUS8jE/fjFxshF8IyovGbRtU0NpO5xxglgQQiEQvSgT2F9vsGXeCWvU2EBLX
Uh22S0uqC5rxlTNPix6Ucmysz5VUKbb0N2T2jTH5I9flzMHs1H0PTMC5A7ZFLpoXi2DEkmeM4yb5
hsq9gtIOkUlNJE6cwVykd/tQ4MzuqtBVWTG24E0PEW27BlaB4ZNh8D8tj511fZmIpmMCpMtlyS4B
D1dE2KNfMDSWi+wbWcd1PnLQ8WMpNQG1VNS4ihqwH23mSq5DPgJEDSqeJH6z6eHpEiGdHwLe7Cu8
Ffql4U1rBiX5inE0p1EofAz7TzomSUDP+af3EpyBkEFyoNjOVrpNc6OuxXwvg11zS632fVRw/cpu
jCMdFszUCko7VD4VoP8Lw2QpaMygBniXBVmdrS6TqBcJmKMEy3HEFcC8sYBybUiGiPkGGxNeyBK4
wONpoUz00eM84fOLs/rndN2KDfjA6htn8CuxjSRMborb+KqxuFKhc+F1Waix/OAyDroJvBofDlKr
Klc4/YlmyD23dX/K4uPhzlnbui+qG5fiDVkfPAkRhfnGap5J1XJJ7pUVr9DwyIru8QKIB94aShdT
cbdPUAzh3qHL7VdkSpkHCMggjMduAbwTNiJFshrQpoHgdYraHP/YNv58n5Mi0hOvPTvhNoRc3vRx
llcy1GBYzfKB5WrW2xFWoAomDS7cWTMrMVkUDtZqEWKgXwACjPj3BY+evwiSZuMnZJGWQM9j+DTF
KD9o4oWvFLHBoIynfLZyrtR3tO4QkobnLW2qkhmHDGH/uCKXYZ/G+AapP65mSKIJ27JnnlKiW9nO
7T8NHZUhyr52rsYUYp2e0P9tfbB5hK36a+VtmnWll/3D1+a07W9va6kYXyNWV/PU7qN0lUy02oRt
P82oB4g7YyH94wUShXGunjLNa7EsBtzKBJNT4COrlX0WO9tdpBLp8yLA9SSMjpuUin5oxXgNMwnu
uFo0e/hTQMFlz/aheUKXshXVwXTmZP6hDaG65SGirwX1y9+saRowrGzX3Gulvd4oUIG1ywNFObcK
AhaAJwwDUaumXlEKHIaUZUBTaW7SyYVy7/hkMwtCi5sT6AlhjG/RlgibO25zNX1F9OskSiTEw4zA
Szre244z62RFZ2jXHvtrLzoLjm89uQ7pFgtH+RGJsMcgki5PjDTGUdi0OdL+uOWA6R0PI0v+CTIz
++BzySQoWXrW9IqLdarN8jVxSKaN6mojUmA5M7kuUO70fOGq/WLU9d4AuQR9PvOnRbpzxEgXCko5
bS7fl+WWvpA/Mi6vUJ3VPvb5osE+9FVdrA1nKLF6WQiCmxLaOZlewiUaIKrlhKTMiYw9UMRrC2ZB
TRH4CNjyKrfg23FBp7z5FP231DvUTDJ78DU6kNYeeZDuzGx+HKBw9uH2TKdfjapFcEFtVT7HfmDu
IGjqgiE9c6y50Sk44yp9VKHHFSaWcHnXJJVKnqV961ktTHdtMeo7p3M9KSHBApUXvW0UUx1w2HPk
UuWymkCHWCMjRNV0s1YoazcVtXAXbYVqGwOU2OG8Kgg12++KH8kqbeuc485zM4Ig2tsKFWJR6Mlq
WAt2EKFlh9yMAAcmK8HkRDGuFJPkNawgmvJuRH1THfceecjImhjwhC17kCLNcbHzxiMi4TjYbnQT
kWSgoply8aIvFpLLYcrujBGESWRUyzSjDbiYUo8o32GZ2S+BpXBgSqElBFYfgAnIZfd4qXm0oXsm
u8MPphY/H3DHb6NQxbAl07FW5ejQ/s9KLyODD3RQBejsaekiYnnEebf8uUvpQHgCAlzjdnXgPPEi
L+aCzybKAcW2y0DTr41m17MoXuSa6gPnOlCyFAzFKcRgAvlCpDyuJksAlcj2Du87PZ4sAZbDi1xt
DR2wFE5VoPFxjIiZHsyq5ehrYAGQay5lSoM+gcmSML/jmVn+fmxgDy02NvhLboP2D0Q7qYKW7UTU
v1brQ5zYaTfh+sTWkPVyExsdOC3BxU8HCZLtcs2r9N1oGFCyp4TWrLyzIt6jA4lXIbItrZN6c5xl
Ude+oZGAg/Q5LwgZPl+w1miCXv/3sV4fYsRj7XBv+NT1y6TAHaAKGbWF397jMNo2gRVckgf1/X+M
4hFmmviYOhKM/NQM3tZfUWUrBE2SGnlB9DmQt+C27QRYUm18F/7pLWCT1geH/9HzV0j4PBoT2I9r
dXpwIZjul8ahgk12EA0WcgDj48uZRdofeSK4/cXOxE/4HbB3oSOomLhZeR73wmtj0j6FBJstRsQh
fg2hOHCUP6DYCkHrYjeT2IFggf++6N4+YOP35oKgr7jU9wu0/TQo1OtWNPLYfbD5LgVGKCIH6LE8
78UmiJmC046iyC85TauemIqaa+6zuwpyRSuFe6ptMQMNSKdQSpneqYZEfII58pMXGvzQ22nBl7mG
d9M0UBqRuE/uPmZUrB9ZFLDVJjVQjjLhzNujzskYjf+S54BT9uGoFjWltgUqRCQ6Q+Z4Z8Zc3U+w
iYLUBPq1HPmG4t52DiakD4knza0bOyHInGE1DweUGjTq96Dbq4wP+n2f/4TIBbHWkAlmg0YBwkec
0Y1jEOy7lNjEXUoYYQ9hKbo3fjnbxbzKI3b6oHZWZV4fa9LFanJFmzCOxKNcO0Go2vXL9kj04Yxp
BBxFWWen6K9HuO66dkoK0V59zbH5wTMyJxv2daaO4l64DlCxA0l26547GrQQ7jDpQ4NSSCj4uNgR
NcofXDfmUGqCFhGjm9Pvz5FMZKoRtSUyNPPtM/1YMj1odWR3BXFzx+HSImeFBEfQxehpUVP6HWWo
fOF5XzYrAv79OFj/+NbNQSxNju2Lgv/bIuZmN3Kp26g8L+IQcxaKwCXGVoC6Qp4TpSPRzCOkZmlq
RP7ROlTTwKIXj6TBCUb0O0YxOE1ToEXWhW22HhzfbLW7t3wObiPMqWjGANhocbyiSG2mMCe93JKh
JvMmz4TH0aQw8X/t0ke6cVisyP+rCs/swfdGUT/fuEwBLHymVMLeqbTZwy8zgZU+4pQ5C7co5Bpd
24PDfkEgO3c=
`protect end_protected
