`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
XOJbTFlBd/zdwNVcgqjZw6nV5PKHcoWknN+9sfgZQmhXNjyTkS3ZXXDXPp9szlicn7NcUIHqLDoL
hA2mqyvVGjH6HDDToIf75jp8eF3qY21Bw7mHpb63Li95bKWCctNtE3MQCjrq5oLgc5MmhMZG5LqA
yPRoElponubjrwZdpvjbbeKwPo8CfAHP108rjIV12NZmealOMfaFQ0CvtMijvhWEm1VaPHI1UAQK
EMUYCMQJn2BTZorPTf/5IOCwZFDOW2x5b78hteO/gF524BXsmbLC4JvsxPj2LJgqXQ1mPRtDgyik
b1k/6ObpnFVQHF2niXbGutJriTrYiDWS+P+/pg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="zvwpz0ZwbFyIJb4mwAB5Lup0DU0q26HymJr1rC3CW+4="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 205840)
`protect data_block
0rt82XrbusFyZuf/T6ZOkU0MHS2iALjGKLoLSZMHzQB6ub3Vwiz+5pAS6J62j05JHFVoLdgatPTK
E1nRpBxLqkyYLug29B6HYEcKib4oLjLT/rHjXXTBDNZbmNcla80h2fV8SzM58+PjTuLynscmBkA2
rk1VPEF+6rSIcvBp0NHhI/MHM1AvRUivHvehp6V0vd1j932j+GaJPAdl1i7f+HvbPz+3pLe6aiE7
wba2jFq0nL99Whjm5IVGzhvOA8U5Qb8n+LFVjFxeQlmR/HhmvcNoioCmmeIaVvbyTE1PJ/bVzUjx
GCTfx40320ZHgyorHnpqdqFD0qre1hm3HCBoRip/ibxdWn8vj2xKilFVNSj4oc68bMC52g+6SPTa
1xZ0s3kcVIBuUr+669dyKpvDX9mh+bRCv9vwLzW/djkO9uZv98ZDhgZKIAkRlXZ3Q89hi8CljYR8
k6xBrbW1EXoizUS1MQQd21/WnV3D3GJWHAAzbdt0/LtiLEcIGzOSDj4SwTVNg/GwCeTALUz7noOZ
/qtMJgSBJl3Tdlv2tWVTBN3dq60N9uyRLXHxCvfXxitE/o/qd2iE6ADFqufE+8Zu1AI3pBrGFpVO
ZAWJXzC07pgP50lrCE0z9Gl/ppmrwcyHWnoGxWIr5zg3uQ312raZOHg7EOYO6Pu/vm9mMKf0ZNhX
lHOenLIuyIswg37+Ry8Nm1Ej98BH4+14vq2Gyr9DYQTFtxFjnUKN/gfeimXTCl0jR0JX/Zpp6uZt
tlGi11A+aRP++ni73AeqpD3WStDTKLOYtnjG4QXrYvvEhw5BeUiOHxNKhcE2+kJPB83MWmrRBK7c
QAsTq59bnV1M75B0a1vsNzSG+tnilMG/QqOna/FWZyT+/77pY3LLBc0xlejetWn/woqrULsNnexC
el7oJHKBPaSSnrE6UDoKjVjyK1xd2ylw4QPeHWSMTlTnXw/0ohnkLCqI9+RbwbGzpeFsTtjPxvpf
uQGxPV7+vXwns6KRZTOHgSh+Jk+NRPGtyfq/6qupmKqp3i+nBSKYTxAm0tihhJnVYXR0T2WvxSK+
cI06QpPRxLkJjk6nhggFF1qj+lNnlP2QnW7bGFodRyMydHCRE95i/f6BoTu71vg+kz1X1ct6GGi2
CKf8c1yOKyN3v2gz3BHhYxo/gzNejMtJEbjXAFlf4Fl/gJEpLzcxL7n4jCFtcoY0NTN072iMD61G
oUzztVDBQoCoArRDAEciQSmlfKCb3g74DqYfQ99tSnTwVW/iImm9HDd8VV2KW8Z411DTfKUTduW0
8ws7s9Dt1/yWX6ILz9GS5zZx2Kp73z4JY+jSLmhKgd7ThgdiQqpU2qjaazC6DWTh5Az02H/ajlhz
SVjYpfx400bbAZkmZ569/Vd0jmLS0pEeuoUCtlX/5VwzgAudqnNrXtvTH6agu4EjxzFammn4AV6C
Y5FxUhncLHoVomhCRplOYqhi12YtS4Aljk0CBrWpv+uEBwkGu+IvoJdUgks1ADHxvLox9s5lrCWs
kHYEGWv9bSVREgfl+QoyhG4QQrvnMaJsj1W12O+Fmn3rUM5+5HDgvN5Uzr6yZvBhAZOtF/kOageN
v6Dj2yT6LZCZXVzPGxBbwhOa9gXfbMZMFo20Akg6lLxyF0AR0QyrmXsq3GzkNVStFu8VaZgghuXq
gBSJBUVhGCO8/x2ddaQQh+M6tjVv0zIChWtmH0GOBzJGMt2OZBfh/YcumGY6ge47jqYxjj3iUxf4
bY+6DviZ756xP4d4Fmywn3UF1PBeNbEpKyQJVpTMasyck58qpk1h/RXqIiAAm+ZwCHHtxngLq1kT
M2oeghm8qxbK63pTIRY/mcNkY776taczLDuEcilpyeZgDrBpzBnW7MivVP1Q3Hn6H0FO8zrwMdaR
M+NZSfeYIgN9Ur2GK9V9LenjmzTq0ujhhnZwPXqTKAOtMHleQaqy6jhIHpgClDxiKuOVq4NZp/HG
vv6gRqD3TO0jRVx+WAXPl+IwxhZN8waw4ouQlX7R5xFXOTafOZ3TYG/rDicbm+uKuWCfHiAsR8ui
mmA31R7L2QUVegwbX3p+W8nGltL6WBuThwXXwxGo1f2GPGKxF76DrR8cDfnr9lQJxFccbJ8FAZnB
tNMFIuI8muIEhweIUD0spI84zMs2/rPkYdbDRYFY5KtV+bkKXhA3u9MXR9Z7FdPkY6ailqTx5zdF
Zy6Yr4YQFlJbPP+meMYqiYAqVre99xv6sJwTc2pMAJBRvIhWltqh2AKkxhlL8NhFxYk59k5ByIKh
GMqI1U4puPn26pkY9TZlMva6E7i2BaYNEA/I8u+POz6tmofRH7FkJWZQbebHcau/pv2kFt/n5y+x
ctfqZ4zdA9kMznUHjvI/h8Xb/GwRc++P/1wmojNb/RrI8U2wbasIghSMibPa+WvCuQPezkey+A1/
41FNsSbeKI4rCHj2opDSs4EGnTABcf1+z53dzc3axANzL+bdjlIyfQRQi8BsFLY5/cq0W0uUdqGi
+Fsz8NjTFdMrn/9ggk5qMmxqORokhdnbMu3TeOgrZVgfOhMJtMtb76W+IEpZ7BmIaAVC6ZYDRxLv
yfWUVJY07R7FKhf1KLsyIq4uS1guinBHzP57crcbtUKpUITMEbUiYLc3yQgrehojhpZ4vwQDtRRk
l0CMOHxgWHE/+zF4Pp5mPyZeiy5IvMN1GpVyF++5podyVeYjHn3EjXgvIIHAax2xEaw7GLp/dVdb
MFfEVqdUlkGjvS7776odZVBXR9TdW4X+vT9GB20UjKeBxS6cpSvEuhsddK5e90OUXmWJuTJcLDey
jo1vz/cp0SSgABD7/typL9Peiw0EJ/MO5UuaxYJ4u2Bhhd3gDOyuAsdJYGY539yexYttCWcrPP6E
NybbKiOEyu+I149OfkVETrm3FALAzl5ayAJ9lvY1gex7E5ePrXlWWrkZxpYEpq5ygMaBVAaXmmf4
XiLnqzgNWBpRu0G60rlruhbqKh6LG66pViKpp1sgLa3JpnGTzNXEjQplkPPNJPAnSBpgU70vOg14
w8NfaXq6TjhYxL0FuJC8jtUoaeFf1tQHPz2wtJ1JbesilwJEmE7X28TTsLgLFJjkuJz9cmS/6dmt
YIWOiuEssugzbzDj6wSIOMIVXkt8WA+YfHR6VUFu8564UGvq9zJW1vM661+U2rmQq5JVcH8OU0oI
tJG6ogZ9tj+KlYY5vK9Au6S+downp3eG0UKu9J5OZ4NJdkLvSaCokCcGAE3OuUswfVPOcsP5Td4t
2pRWmlB5uiEza/yV/OTIR1Ky0MMM/A+QCXvhyQt33x7P+jnlj/BTQ+cY1UaT3V91t02VpFy/09hY
thBpK4e+MI7Tj3N2Pq12kPHwishg6rtTTWFu8Fy4sXI7D3kpJCAP+wu1mGogMqAir9dFPlxDSbDI
yfKDY4tSHu8MzqEsBfWp3IzPMm0+9pRCtQg87dNT9Q4Uq05FL82OiDcTL9r0FLNNsSEk1fj78dKA
B2B7hG3fk0Qfvvmx6kiOHZrot4ziuwnaiJBmEZPcGdi1D7MNKWFS4+ED1HCngeFjgwmUvfjH4XVy
5niAQzJCpE1Lrle7SK5ylwt0og5pxPep3psR2gWCmaG0qOW+WjMxU27ZIOQd9+WpdRG5C99DPW0q
C09Bu+UwEqiOkQryH+1wdsNV9eWxl7SShNHpU7nkuJtsNEQi6gucBY2wjmc0OJNoqBlHFBnEMWdu
aCzxNLtvureGyn6pLoafHt0iM9YO9aBfSlZJHjoutXAI5TQR9fodsxHaucqfWLkiqX5ORo4UDc8K
tBO5xoGUeW5+d9V5sAu6fAGHjPsr+IECHT8IB93eKAh4kUfdukknaIkru5HF3x4MMCtD/q8zkMue
ihb1oH9EZly60K62e6Dvx42Zz7kol6VfOXEcAOaMQ3rIiFQMdO/MMiEMHAeqC9OTY3I8fTJ0NR8U
kTvx3vDm/VW9qd5XHErNvk/RAOi57VILqWAspvmyjbs7OBqH0DKPNqYruBlQRAl+xKZ3DRWGaN+v
tAZ++LH8/RMBGkGIJOP7rGBQkq4BVHgn7jeyuZ55eIOIplWMzAKyW/PlFzpd8z8KU6UYlZuKJhc3
1EqeAymqzVj+9qgI2ucsX0KlK87JewRCAjZ0SQdCBs2BQ0lsoc3SiTszVXKNvIydyxxpltB80zm1
7JoojOy2h4HHdwsJgGZaa1IyxArPiM7aj1jNg/SrHDsOPrq5VFaNzXhJ/oJT6sBaBS74khXeCXoN
e/FOCo+5XybzbYeKo+Wv0uqV/krOwfnViwrfV1Era68NecQqDG10nwGyYOxD5tZJv3+DRJXnj7u7
KsgtfGlMMr3OOZX44uBrqnyXSQdkEsn4HxSLhCF4Q+B2CewtFgNGOWT/D2dNaohPvXEQOz403fxR
P4qbARADGXq6mhYkZAi4PKi+Zt5BqEazrwDSL9AvFTb6Stl+SmU+sD6U2Lrda39wLsg1dmfH/Deq
USKNpgrheA6JKJ8M39umUuvJMTzp0/Pm+xLoxb0BHjGJMwm1HaGk67rSyJ+O22HRgeW3CTToxN4u
93iMIGn/U2FzoPiCaYm5wfDzRXTk4b/fLnbDV6kRvagV+ec0rTLzyS8TYqXtI5Wvy1OmhtkW8SHF
1Teyl+YYade2vuR5sZz/z3i18e8ZfyPYocF3K/CfazuunSCi5/JUYImZDawRBYnkaX/BgxHzWhI/
fA6XKF6FbScrXEsVqdvIzzg8Eof3kdXBU5bu7RKzEVmjHGnFxFBYMHJ+6+O3o/QT9LTy+z6Z1obs
tgPu0PIql6E2duqlwfBkByGAgvb6DRLpaQO0Xi/sbMVGy6KHdN2N9KgZilIXwlYMc+PoyffTlVdK
neEPF8QewGYRHgsDky/Qe9bv8k7WzCrEPDgMK8BSeM+5ALG+LPrUq9wjTHS5YQvJqnUvJ6Rfpze0
cmypCPv8Qysyxan6Iqd32hsLlzc+HHwosbKcvVrYhDgbV2i+wz7biSEMAhL8rMk1q/CM8a43fa2P
VnuBJlyXBJSbaUhFqaZJgPGrf4UXDaoH3jtzpqxq+5KaCroD4ciR0q6bwsxv/AFZlQF050OgtmxZ
WamcdUu/LpP+XioJ2BeVYi/eXpOMyqqfKv7GY+OE6+QARkYrzRrXB5mhuh/Fxpw287Afzvj02JwN
wpVgx6+7qbHpqdmDfcAaI/g+zqJ+EXnHiizRfN65v5eECK+gBwcIzIxov4IprABhvAuZpJZnn7Tp
Eu+p9AYaDwTZnlyL7SajtUBWtmsHanOVNjFEHCk/WgeKPThsv1Z9MtJOH1Zz/29aoQpU8LP2hmFV
8vGRJcRKRPuPDycK2y4C1CVaHuU9u9+Fr/IsqGpU0Jfi07HQn8PwcZjV/Om7MwRKARl+UijMi2hg
nOcek90pEAJYvS9PRFMV/Q69xrFxSO82QA0MkGQ42SCyx28oxSkOEFWhN+q8y/eutkaZ3szppJz3
u8SDpbZhNMC6V407Xp65I29w5r+AkpArKBVd0NMS7lJiXkZ86k1yhvoaeReum4bQNKZN39gtT6Fs
B+arpD0+MRsztUgF/P0XLV1DkAJYTQKcZBfYtRwljLMwFKeWVOwaTIe9EtsRDT5kCGb9QJKfkUpF
c7oOctA09z63TTsOjXEkurv/AnXeAwQ+U4SD2ZkJwxBKzgnESI0N4pkPqIPmoyGB3TqpkmK6t2iR
2gS5YxcbuEFN19di4Sqe1uYeNmzTbO9vxE5oXgLXt2V6qAsB+4RAKkztZosobikkLkxYXsCUV9PY
eA/f/6YvRwZ2iKwBFikCuduaAF54a3x2aoCmUUFmKQSl3J1K73BEQLQCo7TSmP1nI4u1Qi0CaeGJ
z7kDGwWnCy568XrEo7IezONBpwbPE084yUNxt8n4t97VkIoqF1TdRy1R2WpWrrXx6Yea9m+9xscT
wd9Gw1FunwlUX/ltRA5nxKF2voRecUljm2RoMeccIhcOffoSCoTcFr2pfVCEQDp5QhRBeClBHZV5
EneNtnbwAT7a7nr5R6i0NQlVqwA/RpPElj1jHb9UaSOvT7VaR5/dhVIY9SFByYhV6WIpRPhoUvao
jO4MwJrthQ09aSPlOSiHm6Wj99VXEtrekyVVFRWEpmVODFnWcy+e9BjpFyRZSiRHzIedUIlIkq+K
NjA7HT4rCdVxixcqWavfiROfIgtcMHqCBtR91a7QgqHByUBmXW+FPKWUfEDSDoTnn67l1IAnTUaB
s+NxgDR7lY4qR8WWVFM2qKmF7p0mcG5r+YFRvX6SKAA+P6TTHUV2+9FFJf16ZC9V9iXFw/y6+XK7
guAwd+h1ZjX1tD2QQlAyOFzgZGeI36ZXcacSS4nydh3Ol8CYhrh41xgVz/m1x1gFsod4U12XY4rk
WyxYtDywhPT7hOthPTKty1pO6VN6p2aW4P8yPMt50igVEol9RvMH8crcnX8v/x+STt5vJKmQZPum
6zfObcbrPqO2rbY/ZnP6ihkyWcDLQMX3Hq+uWnJ6Mcj9mFzTcZmZ+d6CehRSNvEABFHqst3uHamg
Epra1ThVld/Ypigj+1qAg3pqE6NFsWlGMdH7suvgezmU7iTZBi+u2ICro22NU1I3Effw0Z/FzbHX
zf9TMa0X39huABIqhUM9L7VBNstFeOidAoGqpovNZNCXZ7GYtf3KhetYYIGEyruf3yoRsfcf9b8K
XaLtUb9mfAjQBQPweaYQ60oB6bkOWKT/aUjIvbbE4cR8P6DZhl8VvqiwfUmXDJN4/2Q8q011tkqw
c3yWNWarp26YbcYV+j12PJqmQuwkWdlmins5te7cDm3pYbgedUB/W7QT36ccEr1ENFTP3oKGHg++
KvATACPuc5b9lAbEzjjj7JdVc4mtiFsgSYkfI5lmccSELtv3P9Q8qwumcLo0ZPbDiRwktAyCsPWS
/tou9GKXfRltlvnNi4nDF0/ogPkDGRU6qCosGGFLeMFDe3YOQT4kowyPZK8nnNpVkpuM6JMVq/lH
S33k/p5NxWFPLHz27BfjRzHyXhhw/g6AidIYVxSPvC/+jPqXW0OAXySOYzB5fqBl8ZgGGxCunn5r
jg4uG2Xm2rcufbf1A7tD1uNepbo0/eVlU1ZQ3DrEhJHZfX52sh5lEvWrw405VJjh1byjjmX1k1KN
vlhoREPvkV2F599R32S2bWJ9TVLu1F8mKOkPSD4DDp/AYVG9oW3bp9aaMtUhhBIrgIjwl9GSQ70B
DBUt6gcywxqmLrt/PVQEClIeXyn6LeBUvSSV7418mb5veIXEjjE9Vmt0oR7A6D+dr2U3y4oyWt40
1k2WlaCXCLFxGuITC/65LUli9GekC1UTEwvHj2JT17efLK8NH54HCVSkUiLYwfPXZKx4cycTFUqP
/gvI6qbO/1lmSRL/9iD6InA1NK0QDB+Lf9ZbSRnOES7jsvsdVLtGZ58nDQ0EnFCmh0cXH2jYvpzY
sOY2QRWcFQzTvf/rjUtVO7uukZOF/P6txOZtNmnkbgPHpEU3uuOMMkKW6+xXxnYKpoI+YNvCIgYi
44ir7qNa9m6d4qQZ824KPYpCKrdL7z7U5e0EEAAPV8x0DyCV/WURtLcv5ezBG5DNqm8cmekLHHDj
vmEiw4emP9IQRGig6SInKoYKsvxneIeIA/YSAkBR3lvvweQAvVkma0U2RZWl7LiVvxcYGvxPu9Z6
DcRPVJjvWy4R6hQ2TTbXRgczq2HViy2H/nUc6KZ1Fxh61z75VplSQGWcSuNM5WNcgUKd8wXgmCBz
VWioz0jWKX/IVjfoXpnZ9ibL4Y647Irr5M2UTShof//P21hdotCMdZPwQWL3GevGTJMVJqX8XerG
ZnJtKFCShISMdYwwbS5CCr+yWAhD6OyM28zejXeNtZE/UqLSUO340RtAKZFrjBlqY67VfjXsB2Qp
QWY2oeSPS7xcecjS9YQtxEv7pSE5zOxN+PFN/A/Os6hqk6+puEPjxHi4kiwMyYRDhQoDT2PIZhpZ
GYRmpVmiyNSRO4hKHv7QlHonRo/TOaVINhMZMYHAhNe0uuw59BVK/E8BV1/r67AxkAq9R3ygvwiV
jVyRFuj9Kd4F8JJ4A8AVlgE+ftt2XNCn11M1bi919aZhZYHkPhd8UpCq1XZq9y6yElRbG6syMkCI
bkXft5ebKMWjsI4QP0zFKjCh73cdrMRIWn1po3u1SlijDM0nAGH/kI8z5B64ZywOwkzeuYHQS0By
j4/pzovanePcUWbO7lSRYXAGfKYzfE+QZjI6KLIYxZM4pXxY7Wkm6buL+grepl0zkeFmm0bHT8rg
2egabjC8DxUWqi/QkH8aZzVm7qLw/7n2NEU200pGIK7Epgf4H1DRUcukxLTAsZ5WbuxDM6sVeic2
Oag73/VrIWwcfrTcT9T+cl9Sa+6ztg1H+cPlUi52qDFT1YsEbT2VEEVMoAWiwTHqbNzaEronMQjM
PLYHBl4rkNQZ0tLvS4NydXT/MxCB0jezqSiGfnijWxPa6cxi/YWJCmW4oNZbG5Rs0D3Wc9hUi6VG
RKcleU/QCTZvdQ64iusbs7zXbHEu0/g+E88fyhjrr2OlrahB65dcD87F6ybovvJysyrD40mVuDRY
AyFjuJpHZMAhsaODWMtY7g+Pd/d0yAOBQjllYJE/89mkQO+aHhYYJDBTSwTCO2R5cQNBRPv9xx7i
LuiT4KrEUhKl/EZZ0rGFfJl5JW7blE3xZxtaP8GfBX3EikGtynB1At2x5UUenABW3WK+hIqhrUKx
3dgE88jAvPi3aHsWQM9UI9z0gUDrTuU8pCD2y8kqdOwRSyDFd4/8Wa86kR4w7vuuPFlL2ZoEROGM
Ph7h1uIOwk4rduOQ+LTdxKMVaaj/tTD25Olk1TO5sQpbnZKtVEmkWv4ApItGV1HwNkM/W9f87WDh
lZiw6wK7nuEQKn5hE0cIddyqWt/Gua5vmxvaMm6wiJCK2TLQefzYfD8zw6BPnlKdTD4mnzw9exA7
hMsYDM5G+Y6gdLTYWb5WX7RQpyPZM9AEbGHBHXhjFyMKecx5bah0VWNz3Q8q8mkC4RVYmY9lnXwZ
4EnePJT8P010fCF7dCc6tx7jRosUxhEZaDRqLqyZDftlHWRTI/35dTIRfiP0E63HCm4LOsyYLf/o
Ro2eixqZkbEai6LIocdWLnO8N8f6vMl5IcOSife42pUdow9UvIwFKJ50uAmweC34SW3dYMrco61B
uNesGfoOAgpPc7MzaiuiGhqLmGDyI1GEF8LICZtz3uSqOQPPCgawfzAgnSnLPluPQLKdeu46sLJS
byfYS0Z2GzFA65CrgTdU1Ba91e7KY6y6X8uwQ+rxCoZDgQ9J9JB8OtbnJT46qEXGWcDDFcp8p8Et
xY7cOJrguWCYjn9RccnP/WEsqUMfXAVps6HAkY5zv+nxlhP7VUt+Qu83r+3D396hSkti9ZcezrL0
GScw1STSExCFqBjGc10Nk1Tx/ZjMgAtvW9MIi5DqvMyHNGgPLMKsYerDBgJfpld7llfBiacYLji2
SiBbRLA9TnSiNcFlRQoz6lLX3aZ6DXi5XBdj+0fmWvBVRpJEknYXyEegvTiDSomU8pR9wpWP0UNl
3NDtiPt6JImtP3kXTHniZSNJ0IwHnhKEnSUFAmO+hgFkc0Cg1+IoXLndUib2vBvyEClCDIaxZ4uv
Rkfg/tlas9Xbp5bN9R7+RlkgWm38XD99PcVpTWh427DsprdU8H+2zXNKuNWlGJaNqrwwlqMdDn+l
WksodiXPMXhGbUS6Yymorp8nlPq/uDSj0VAhp4WphYayXyGo9cvk4/dg8rV/vXG/KxTxJt3otGC1
UQFAMLXw0X0w2a8lQES5ZPJeoePnLePkUq7zwPbWQ9DGBvoVSJXzssaIsUHilhLAPzhqmsBLksQJ
ntmDg7qyxc4jJcAhS7uPjTKMDeMpcAskuNF9DlYfFQ+uU+J5HtypkneApwYxaz+eHCWvTGft3dDM
ZZwSX00em39Q3yq8AmnymnfWQ8DLmTlOrKUaVk9AX3AvwW7nDNAlJyK71egRzbw2Q+3uMbryyM1s
uFQ0jgR/aJIz65MhUxbf4BMZAuM6Jy7YF86g8RQE+K2IGunpoU3Sha+QARm+dHFkjRa1mcbBvHMS
80T3eHSsqLj9Ba9Fv6Zb7AJKJsH6/gl44Pm85NU4rxEtJbNBEL2Zs+ugdDWIgwh1VBz4aU2ui1ZH
Q0/ASV9m1zzt9/G1spKtiBp1nTBfbfx01qINhhTjBZH29X6PuEfGK7DNEFf/QBREbuFVGDNGaz+L
t33xAKJ04wNtPAZbSq/o4pFEbiqhC0uY/vg6BRGfEW8QSLLc/ickJWAcMOHIgp4bpCAtc5XxAk1G
Ohbdx6uXePFWXqacJwsd+0FScOTp9iY40F+uDBpqgDqcMP6N7O/jfKFIQcKHCgdAsedjCxIYejtt
2BkML+7qnI4dnNq0Bojr/ZH5UH7p3aSH4xIjMvvixsgHbGNxbDDtQQF/huWmALuesQ6M3+APKhle
uWIALLeHjRYHOULsoTOyy7ZGuM81gbhpYGGV+zvxYjMZPs9kGQo9Z+vGKJecPgdC3uWuBMIkQBM2
UnOEKHDhhbdcVFCSzuYO7Oe63CCNQDIsNPTimyp8NuQCnl9w84ga+yGttwRhlPUVa2tKfysBJxAp
Xyc8o7eWIpbQy21JtItv8og+8QBh0GQ6KchhHxy9GduwEM7YLjLa5JbdmngVhJHiyo4hbM2nYKXk
X4oOsaGa70wgg/vPCf8gJUaxi5z34wGzhyn2l9qPtPW3zJ6ky+AzXKkjr5MGqx+9iZyGeVdWFmx3
lEZ9jQTO+An2enuJ8zVPR5glkHA+TjId8Lro546HXTKLbJgxMHj6SUXSA+Kv+Wihd3C1JQXgdBsl
SIQhYpzp+9EboXxOrIGHwwofmXGOvwLqqOao3HU3xCsJg6citm2iuQ5l2K25up0iasZd3yKFsL6I
Ma0MG+CII1jv5omzWnJlaDlmmeMGOT9zkX3GqE3onhiqQrvY/H48593WXkbiIqGNZK5g4b6/RxNH
SILIgInpx4tWjV6qezhU1ykJt9lLpRorrFQv++8vku5KEYZQqc2afPQRRvR5HKQRvmU9zDdEuXCf
TFVRes6M0QXrS/X1oNAf2JRqGAZycmjb1npu9zLreMtSx+Suc/ABjjqYKcxtmQG1FKcwoaBA6d3d
zIUJOenfHP+XPK4jP4twpy94CcwI5P0C3NAccJNq0SvFxL3nx7i8sID5MXQzwA7wWqbnab/XXaGu
XOGxfAErcytB+DwKyc+dnPGbc/SgsWGOX/uSA4JTw/+d6Js5HNjg6l/sPFGNAxlTayu81wx4nFP5
0X6CXIjtffW/ztWu+DWVHFBrh2E4hNqDqAn2bL3OqfMw+YacUIaHfz0eqJtre03RJP3RCtuRxzhT
tvg71cUTjxhrrj3z7JSEcscF7hBBkTB8nxFEJ0M3tCvebJHxZhVoUzbzgFntrWcSQMlHryCftv4V
yp0LmFdSQbD7/O6FSCNCMQpWZjrPgYT+lcoM8ENWEngZno51j0C5vVXKj82GDCTenMS1Y+1KG+t2
3bOZfio2kstHbjWy7FNoUhmXt5D61vNiW9m1eaVQFaHUsb/bTWA1T/6BciTNj7Q4jg+AMMl2GogM
fAN5qXxY+/a6+KKuTXnDKikbN75LHIO0PQFWQCkYMtdXE08SM973bsC2kXVwDiTgdE7TukqBfNt1
+jRvRyWPg+k4MElUFbiWJzXYHbaZA8KqRLDZOksIT32qMn+jbTDKKDOe649v8Z3rzcRsEAqSEscY
JhmmGI+MFiBKZ+fsvROuHCc15Poxg6A3K/fmVfhJ+uywhGk9VSGb1kJKjYxh4Sr5j2n90FwJzDRC
AECAUqxkzoj6/6G3IJUseT21whd9jszpl6uBqLFNMgO+Ne4Rk4yEHWlq1nI3jujBu10XIVJalFbq
Wk+cKsqG9VloR6J6ezocxWgJbrH+R9erBFMzbbz6xfDqDTGz3KBuTC9k0XCF2PjGgPhbDYrA46mQ
jnCUBxklycwk0oB82zUBA8FSTwdV6XOCnbiENtIiNUuYcRm4EX2puXHlQsDirAnePqPMDv3qzoDw
Ijzc0VLVAvOoGjv7rawe6atMM57s/IOVlb4dJkFPh1XbNiBTeJUYXqEsdMHLLsSpIfOtoh02mxz3
E05V5h/jSxW06335YpqpmJWw/+DE49CYnouPD0SvSr9TiSzg5Yo0G8oAz9Tk8OyWMlrV8uuKUC/c
hgo/Ui/l5GZOmvNoL46My5cylWj2KKLdPz5YxFxXzCcy3hxXeIuXbebbXaPojJj5op1JtIncU0Q4
zb1K0a2XOnwD3GcbR2wKPNjTQXBXPz/Ou2er9ys9/s3+Ccen5o3BhP5Ujcqno90pI2ZcxWPUmIy9
zKbjGp9d/yNPczgeZAHNfaGy/UCis4SmUR+sOw1NwmLndWH4RROwL8wuNX3C9ZFZp9cOPTDmQQOe
hp6ZIgfVmU2k3sz0dEGcSdykhDBE6jqQCr4JgdSWmZAGrpFzMY/pV+43U23THsGcnEMpRQACjJ33
ix+OitmezYB1XId8x896Vzz1esYcm3+f3bGdmtV6K14TVtt3gX61YIKawaenKNGTZ4F/1AUZxAwe
2xvi080Uf4FG6ONFKubjBEaKVp65RmejuiqcOAfasmHRtjXuhOxoRjItoUDXV8jpYX/O2wIEr9de
/e+HUNsL2mb37Nn951LSEWwuWDBcf2XuF6oO2BLqfNQHaCH/iqkbzhuac9oNOnvbCcT+rg8gavYd
xaDefCI0rfmwzLRhxDvR+BfRqUUE+VpPbaF1KAuC0eYJL4dX8uABmzqSwk/dtohaCmlvSAHMyVuX
Q8xKLJFO9kybx7spoSLbubuCTu/DVBJ49PAM4SYsS9xz9RsHSWaITufIeOYZ4mc9/I+x2P9ZtfIJ
C32tPNnhsg/XXwKNLnaeGxCqUinqv2+AYeznygC7uvm5AWlwT/mEC+UOvmxKujlnhl4jD//lIZCL
ckneZRABoKwduy36I4b4Xrg8rRO4aqXnOVjTYvT158gV3HXQJtd8Hq/hKe9Y/NA5IHWW/JUVvz2L
P65fQp6NS/8/ss2IYz4ku1QV9s6CogiKuhJJJc/r46WGAoZkqw9h8YgCZMdNAZMAAzOi3Ziv4IXV
qRSgsYZuhxj8N+bUe1L6AwtZiVqEVURKMM3DBNdkYX1jEKjvv023cKhNSWn+QL/ShCVOsvvH8bT/
o1/KhRGbEGrLoMONtnbsV/YWthMTMHEPwoFjcrTWBBsrG2E/zEo2h8En+iX8qc8y7e+f3q+Xa0ZH
2Oa2l2031Qben+h3WpV6X25jwiSqzSawrorysc6CBWRBjscBTAnz2AkTLo8x0i91BoTqRger8KFJ
UWhthvXVsxzyFdqHv7thTS+i/NvGF2hStIWC8ky0VSJbGxfqER6ijyNsGav+slZ8mBpSosHTHfpX
qcd8eNJFHOQY799aVF9T9Y5u02145DS861dAinN2osAT2cAQXCbmd3IBxInyHtO388z2XO+Qog4w
clq/bC547LJ+qV13w9HBNErnMgmZq86vfUivmmIWgg7PuszW2WOYGRumAIBPblWtBIerI/XHxi9u
spl5H7L6bCbf+920Q0HUgg8Nh9xbDJRHkoK6dRuC/bc7jNremX7XEid4PLc9MUhij0gbMwm4rfKT
nWmUSNZ50o/Tc+jvOdKkrgouFjckXIVxIxJniQTSz8UJDNDuBl/3iC9zqhM8KKrHV99NsnUq8heV
VX1CTq7PpO15b+i+pWjUmp9zkVfKPTFavXpsG9T0/Z/MdmBOcl9egNSYTRsHibd33ap5feHyllov
rsiGsJFpxKInbP42FV6pLnaO0irXh26ud+0BQnhZAPRB3nTZLd6Oe/Rt2beVsd2dF93lewtjMPy3
CRqqHXEsLx9E2OaY49eIQeUjW9rwSfqfasSp3N+eRytJyeNLqBcF5IZn7dfgNztwkF9JmzV5S9RD
CVxOniqCRS+n+Dfne6pfCKv50d9m3R8dksXZ5PqrqqDxhcdwh4U9fz/ZXB+d5ou2cObODKN5I0RR
sULA71x1TQjH/H2lHOXAX/7j+Q9wZnv7GmFs0KccMMiYBlvgXybiY1usrGQIt0WwuJ9/qMiqh8Nk
V/pZa9xhay48/4cFX2jYWEMoBosSpKSYYRrRpwkOrtmerGnCWLmuWKWslZ7FE4g9o3lVBmTY9fxi
d942XgE8SSm2z4oe7xGikiyj8tyzluJNAeoN4uGp+5TZrjaqfJGev3WalD6+asNdoxXS3zwkQla2
5QPr7kU72Agxv4Hl39HXiKQKqO9RjaCvPFhknNwVRki9N1g7cD5L9uZDlhtQv0F3tG/+QX2pS28j
KH11mUMdxhcAjHyOL5ZdMOIkTocBAlj4LY79jRlL9YREUClYnh9OhLsgIkzFVfodFRnnkZh9jPnR
74EmQONIW0FxuZ2PrpJC2vHQa5jguTvhV/BqFyjr64l8EozoxF0+YaUsXOoFpg3tLBloAGRiJ3fO
Ro3SSesGa3bksr67jFmSUXNAd18mupMb+iCC3aNrTNfimdROB8goszz17Axl9e1SsuLlCHxux1cd
hjqAsBTha+IwgtwE86/qsbWH9p7zCSGCjZgn8QpVZ0nFF+JxR3QUg8gnEKNktqFkfe0LdnvxtIbm
9asiHmSQwZ50lILFu0VIY5eSewNTKDfpPgpTpO9gVIDDRxWB7aFAPJFeD7zpUZFREGT5ZIdq3O1x
MgQYrEY9LV26J5KNoXZXAI7ZX7szDdR52O0MtwhLKYYYB6s93mqEASy/d3Q7T6BVMX1FQsRvKMlf
xW3PJpbyz5nx5ZlAoO7W42Oq+5wrjb7vM52KgDjrLeNHKxPejQLOe0dQ1hD3Cu+JsjCxNontwm5s
nWBAcpXqog9cHUW/7QqIC7A34WJzq4RqHl/UJEafcJqZ/nVBGaDHgDtmPbmL7DG7l2lC6SSDRByC
pi0XsjpEXlHlL9OCM5ZM7cD7xjztnlK69aR5wzGTUI73u2VJmn6bEsxuVgoXqlYO/BqoVDq6wv+y
nk1Uw24XMTDqbKcip1jBgH4Svjx9rZV5AOCf3UZEbyofeoVZTdl5eDqDHiOEeG70+zjGDINwxikg
mMpXSH6Qo/7i2WeFRWb2y0XK9zBOpGpuCvurpbzWyq+jV74d8rG82DONw3Xb7ueZXwP44wYumLjx
QaJgVZ8vZBwVYPwNzDGuStGaDbvlHglQ6DcRorR3zkaCvo1ptR5fwF/h42X7yXdiMTjO+Ujr9zZG
lSllnHyb1MNUKTS9fIV6mQ6t0Qnt0qdV9EZoSMAQHwydAFWBmB94NoIX/vwGvBq23qGCq3S5+P/l
sSqhzDNYAzP9HK9n5c8AbnrtxQTr2IvxVLRMVQSKsttoQRMH6oZwcOqqeR/JVH8ayxBokESF2eNM
KxEHWOrZzZ4yQdBr2vgxn3N1ld84jSI1zoUfCeOiotdSE6FYqVqaKJdfoqAwjjJxWu6FPm7HMVQX
wBGh4fo3HoStbcH1SevWHozYMGxqkJich9REufZ6NmKfkDhhj5fUaCCdS2fB/mDSd1IRWC+HOTJW
UhpQ9OERsKlRi6BWI5iOUl0PMihlbg9PG2vYTshfQCnu3pA7Zneeaab1EARcFxu6OcIySaQq6DrR
IX9J2Nv6ifj6ZT49s4XK7uVcSuiyvHHenmJLvzWeutFlXdkFeLW8AQldSsKNB+NX4Arx6vJ+7INM
rQ4SxbmmkOzBL9y7YjkRmhwIQNOvyKSg3EUp1kHEvz2WuVKDBo6aFGybHtX6Ef+i5xZjtmuk4UrU
gvUXKR8mBo0fOYM2o+Jyec+c5cN2owALPLOe+SIp6kXGSnorrv4l66jVsnNPM9Z6ROfgSPabwfNq
y7OtNXz17sxHJvHw7uo/yjTvxJ41JpAsdJSEdZSgL0YdmsJkgeQKdEXFHrtMXNNBJ3KKaRwS+Lht
iTXB4f9PbTvDlGsc1bjeOIoRDz+i9Q5S7xOCVyc1WuCmDc8HFqTed3es/8m5pxC4ttBlN6cQM2Nq
SLg4C/+vE7xlbu273o06mqEEw+8nOYnTogHad3FvHzqLmsn4gA4UsPzY+laRYtA9adt5DNE40ebw
xlcCogsaweyl5ZYcFMbyw+u026yrS0Xm53mSjwoo2GtA9nmZE4sMqvvjb3e5BqfEl8BO9oUVNlzJ
RZaj5tlW/uLdu2Cywvk17HtkVYHPRpZqI26M6Ilti8WGX3UplGt3DdYU7jRcsoaczBrKea0o9tyL
qR9OkVvOSWR4mqvTtGWvnE6CtoN/gVI5Xkxvz9JW6HBhqrrWcHLOVIXAEN7g6LxD/4juV3WM1HO+
4zaUv1b3PMCeEbCIftKkBjYran8DfTB28wWrwvE8X+7IwEcFIXQr1ErOglgCFpgdGiAel0TZxDdK
hM/OTp2QUQHuL44mS6JE+SQPD5aNznyOtOOBnujyET9XZOwxrYwFLVd+CoGWjCQWaMWVcDiM7zmw
n+CH6Zju0TRrUwnVfW2Zxx4Az0Usxdo07EqADBIW0gEv07GnDs9g/F9hvfJutPPx5XGIqc6znSm+
Zd+Owxh7i1t+QZWm+U1g0dNq0KjeMQ34K/D5toHvW7Ya2VdbL4C0GGScptfaJFhXCn5BwrV2pQTg
Ixq84LaAk85+65c4tPMdaGrFiNVrsBSIAkUjJ62Nf0TBOwtDf946nHRvtIsMLKb1EtC5dnNdfwju
RXySdC6WdzJWSFjWwe8T7dud/zzeKREWPQDpSCouXsdiKdzkbDZnsOUEhsplJj8OZkOfRrFMhkne
SaLQ42vMqdd0n6RMUZ1l+H7+BB0u/sI/XHitm6rtxX6VVheW8dcgKbJVGrIGOgxvzOnC2sC1fpf8
lueUp8EM7p9vAfEiojId6VsZeUF171/lLr6L6v0uHl9ieI/eHeUI469pogHrZ7lt6DALUuLNw24Y
Rx2PDubZ9+UcjMDTNVrJrYxDEEAUD0Bunpfg1+8gV/gNNVtRALPxLwvTxjddofX55+WnxG6WqQ8r
Jq9sxhAxzkPM/kUbPu/S6w0B871Gh/wE9g3i0xh6amt+KkIL5GL02UBgSTEsFglg3/6GmDYCP56R
/HzX1AsWKAfxd+OmMSgqXuO4HpJi64WAxN6C3h+cvMT0GoB/QrRC2n7ES8Jss0aflKS0Nhr2hsWf
WjLsDgYmA/OeBdFAi1lgfRhwWS7e1pR1eapxq/YegM6hZnQBb89Y5YKjIiEeaGS0JemoMRO12NoI
lccWPS/QQBvXOLVJKxOgUbq7ku0gLNnJaXwDmw+AuT6+rWo8t70SvrNlDD/mh4KBzxXK/saJEK/3
k6djZ1Iiq0f5SDaPuz0LPpMii8cigDjuW7inSTMuipzHet9FKEHEZhzsTCrj6IxJlewmAmKbx1Rf
e1pA/6qjX4aY89yo//1hUlVG6GpgN5RBEVCRaYeNIevWAAi8tyHFubSW1piAXwRO/eD+pBGy1jtT
hjlzCf7GkY2dxtXYqg8jFF2bL9t7Q1vIeexwq/UtaqsoezhoHiMARZDO1FvQhI7ccqc6/5A13xvm
Yjl6EJyW1aJ65lgm7SRxZAEKY6zl7BB8v/427U5dAhcvFB4acYy8npfB+jeQ0duCypZQU2WpjgBX
NuF+cDdYP5n+CxtYJEiFd/Oc4E2owDv5rqaCvf9MQp4/1ZxMeErJj1pMeh/NMEiOm31tGLu8acrC
5RcvN6TfZ85hHB56/oi9CWsQynegDXX34594t3tnWDAzrePudR1SeILk3RkOFztgkW/Azd4wjykJ
OCH1JDdqviA9FuMmqLyhqGLw7Gs1f5bR/PLlBEp4YnmK4DQn2v7OfXBtZvMA9kcHEZRn0H6ZfuUi
58cCwdYoe+YhbgONFtWV/ToKklC+/wKh6iOXglNRFUHINfhYQcLi9t/xd9cJpc252+Suuxtq3WIb
taprhH65kDPnmCfW9pzpUEaDt+9gDoqCC9a+QjKp90bK7hIxLlD0EyrXWLdzc6GJ6+hLK3oNoqAD
f2RDxfUkWFqgpeWJeKH9gqufAgXSsaP22Iu4ZmClLqjzDAX1PXtPhRpJU0GiU/276pIGeZjhgSdV
wRVgYDrXu4BwQ67rA5YamNC5eiYS9UmKY1Qa8pq4HcwOxf1Hp8HuPrrDr4u0Lc1jniFZExAWYHxD
gPOOY877XOg75Jvr89MGggpGATq5cknd4TrIy+63uBjXxLDp//PTsVq7SMwhsSTk9WFg7+9T1Q90
cZ5gktkk+QxDtCSO4ypxyKPMy5x+VcHbHkqtVmpodEoZPxq0Yx/SGnLyjq1ZA5xPcLLYBnkmYJ9d
6wKHfCoFqFnQ+DB8PJvzdgI5qNv95MYeyUHx5I+kPoAZ4vCkPWDOvlRpIq1jMBRMVr010k/2fo9Z
+8vd9hJct1eZImRmbliOv7a7xKyKVBC1uvb4ReeYtjnqt6Nocgk6HM0zj5qdjDp3WBAPPH1ETExH
IBOhj9RelvOZC/G50ie65TOLEWp1/K6bKSOkyAXgiccFG2/3y2PaWc9p0FXRLne2LWe58pUjLKlX
2dROi3Jygyu5Ok+JfzZImFSSM9ZydGkFCFrmGAnw+bCR17Z2gbUWlB42chuEuj2t3rTiUhsRuGUs
E1gp2xWcrB/v+KIQU7EqvnX0ZSbddE8tJBUdx/+/kD6k7vjfxuUtJ9ng9kjdWjm2679L5hOvlli2
bOOYjH6/N360eOQ0TvOHA9bfeChSFKmc+Y+b+4SURMp2l+Wh7XDxKLsF8P0KVvROw6T/+/pS2FuR
5/zA6FqHqtzaSYHUPnjOaIKv1TRESrbXZhUJtbIR2PPUSAHn2ZxKCjD3imTtJRIseYWVzJIFZJmr
gQgNdgJq+PgjNwTU03R89DFidEOXTKBheikT6pV8ub/m8XziWJhPy8xEMUhN1+oTmVXFMp/NX14U
PlcXb48wgBOsE8a1fvUGwu/Ym6VgnpH9bDFyhFjau9tXkeAkWiU0ZHnUtPTIYMWlx6fFApAYWAT5
dO3uTH7Oiz6KdVPcE9/iiJkUDOYKD3/O59hC6unW/YhPnV38OZdW4X35+AyMUNYtR4O5ah/ZwgNY
XPSDIxXu5Mu+35lg6DEAzDJsrK4Lf8xeINR9w6MErUKCJ1/S1Y6m/rZu75YgMfeC/Z77JPZJZLBF
CGFHGn6IOivo8gwG+bjQfYhiMG4dW6QjYsn5N5u1oDWr2FggL9jX+0aBt0uMBN6c7v5/yoDuc5QB
1kabUEHvMuyFZFWHsaJeosdzGlQe+TCR7eKJqlEBFr5Kbv+8MGHAJTW1ICStXHobzUq+hPbvNqbJ
g6KbfychYc/iKoLUfoNwfvm+a85l8dsmrTtWFol3x3FuDCiaAI0jGehsk5MQSK0xbK6/IWonmdHf
brcSMVdFQN4k0OiGpvoFqDmnh2nbXG/gxhv01qFA3xuo1tAszMEJtXjZG6ukuSJhyNi3qbejL20l
bMu2LzPasGQd4b7VnM1AiYwDoK9HkhlTRirGvTIdvZXX5GLcLsDuOKE1OLfKxeic00MpJHeuiIHi
T4RsTeWwcyR7WEOZEgj6Zdxne2x+W3/CcnZ+Ph3+RJU3gbBfLVw4s8j7baq8Q5MOvxeSOWpbw61T
cNgZjm2q+EEIe2ey3MDD2d7HUZLqCMLty7w8isR5mpBN/w5cGLWPOhU11L5bWP3W0gVxdwe1fGmy
1NVnHEwaxHkZ9Vste5fOjoITNIbgXzL6mX6ZcuIjxmzVNAU+qIYVpWBx1zw0wY6Ol0pXOmEXvEQ5
29u9ftxWmfnWO6iqaZuWS4lXhSlNzmAjr/n9UF/vM0jG+gbMo7onP93Dvkb1+CZXRWf65Nw5x3Sm
v6PZEixn0nMMk4xC2xxnQbEFxMsOUPSdw7TpKFPWTfsocqQ83m0m5gRY4pIphVkoij1kqWOz8w4L
JfpAc7xNwtvmtlA0ual6V/DvZVQBM8KP1XGrMPGu1p/sm9VV2v13YLl9JtyjwoFMACpLpyw2e0OR
+sbhWOV2sca1aVAcXPrToxnLsPqYpHjARh6yJRaByHu1OI/MBtmuyoabUbxfyBolLwaa7YmMTbmq
ZVnz9tiCS1g7PffkbMUAq2g/MEqEDw/DstNlB7CqoZqGstEwKLQbbdkkvdl/TW9mUUTwrKQfGr35
h9Al0YpCKTc0PRWVIoeRWhp1FVrbz7WOMDmSIYsZQWIy5PtMSq3UAk/oEsmrKXuYSOF3NN57Y5Gn
l8GAeo/nG98sNaTXqCtZJf3fYSXoKGbP89XkxNuoBBIZQMMwpfqQBZGW9tmxBeccCnOrpOuCkiaV
qITtOTsLjMF0JPSnK6xzWAwfUJ8oneagNxWVGVx4Vq6Dhu+3kBTJOp3JYE0aRwn0PJzKH8q9TdVQ
pr4HQM8kiMr4NHW3ygRw6WySk+pOcPgTBAXKkNd/W7IaenrK1uTLDiRhzwe2iQPUT/PSKFmxiNQ8
3M7kabPpJFfM0UVfsw53s/hVewgbYlZ6BKGkIZqwrCMuMJoFuz9gY4jxU4EIRgRUnCyoytVtfi+K
uWrpMEBZ75hXlceQIN/CQKNwvrXzWlj4FfDJX5k4pa8Oz0OW9rNuuQpV1JR5RXcrsffJyz6/rU71
Nvuui0grzWJy+BLsLnEVkFLw0TDjw6oTEpqof9J94nhe5rQ46MRdZTJ+aV7qZPwGTx1C/06iBMP0
D3tQKGJqfU72ZQKP1oK56quTu58a/uFVa2ziNwK4V0YldQ65EF5GgdmMtqB8fmv7WAAt9KuVHO9f
1+w+4WRTPNZ+RQhYctC4IbjFrik0qnssG/Kp7s/kt5mVcqc8t0ue+ey1249jp+M5rTtHu/luJ22M
7fWwa9ZVrm2wS+NC6DnkNlj5fbPwEaoX6EkU7ltE+IZb8rf9IGQmJj9aGj1tyexhdUPAQBLTlT+B
xQ6Ew2+ubQNKWkQsskz7BYaDj6XRkWItDA+BKhY/513g2axjGbPN2J1JA391PqAKoFr1c2EI2Ejh
n89C02Vwhz3rsnbIeyUOfKcA2XFDYiT/lYxnozz+EubLCbWVYIiAXmw/BfNc5TNmEtVzDoIWVsfN
NZwLeLyXTrjDW9lgrGHWEk2l9/3TBSC1LGm4W/X8emI4FjyZ+fDtJqgFHd+UouNlJ1NF4MMGtlOM
jilrp9HHxrBoh/giNgIblI0u0rf61IN4fsmLrKeaZ0h8LZdAuY9tYD5E5urm84nyDXSBDJkFq2OK
AvOHx8egiqmuawUhPj5ArLc3H8X4wSgMPwr9aENarurIhCkGDE9xgZeeKhzr7Q6z8ZjWQPPVezNX
E5NOZdpIfU//CPoXyeCYYRFeY9o0V3uL9n7UKd59j8NZGQKOgknr80ch9jz3+62nWFXf7xTRSCbp
Q+YBetmEg+yDp82w00EITusi/1s6Swc4RkvB79gjmrkkC/doWmWI0XlpomYuIDm1vQFNJy1XVuvI
zUUbfe0CFVg4AWHY6txB6kTlhJwrc9SAE5MFDpHaUWnhMpAw15g68hYpBEhy1iUg2l38G1M18erW
ZjST6fZpzcrWZj4H10IJuzsGoMyRmB/ju+08LOUxd9UnYplftU0Zy+0FgPsWv9BZUUWSvzHuPnpp
nbWhR2fOmjEPDZLuuI3lgNMRhnTl8TpdcwbxCeowC0fp53c1vgv9kMBmj3cscIF3RMQRCELRlpXA
SMqV/+rVggkekGWMZOYMM5mcvklIhADr8RMh+uK4EPQh8ggqr8eY25z8Z8l1pmwJlCaJ2P9aSV4N
Lr9kgqfY5c0QI3ndDHNP0ANg3nkK6PixvIovaTa7a6DNa+wgGykUJGOwGUXf+HPvAFbQxvWLY9kk
YESco2+R0AS+lg+ant7soUwItAlB5MKU7e/oYC1Ni3EAcK5u1tF7lN9YuzV7D3PcDkYuuSt0eLXn
nNWIo6yIRY7npP5EtRb6ygxJu2Q2RcupsdUJFPKdiMX52CtHaZmacPzWYoxMgdA1DOVDOun94Gcb
PUV9aPPtV48plRYiRJ6sFPUEY5kJ+DocsrjDAhwCENNHEhdGAkAueULfY13EwO8YX6mMCJuvAzzD
RB7ZlNb0Py16iRIiN4r3tnPUrT6hy6kN6a8vFrfOFkoZ6tYjxcO6/9+utv9v98QWBy13/y1uoV99
RDXybGwWvQ27s80PCmUpSOz9V0ZwuJ1NJihAxhLPDR/FEPJ1b4ki5hL5bfPCAGi6OTNwrjp8luKL
Koa0JSZOZube1z41AEHMzQR+ExDfRkFFa+SYGwPplQD5UNfDGVjba36G9nEgr934/gPrStCq4Oxz
/XLYlXwEP21Fsun82h9AjrGEruisJYAhVM3md/mOr0tvP5Dwzzbv0uwoUAG9lqLhu0wgNGGAgI3I
yIZK5HxkdU4ek2T0MTXQn46gC0qAdWWhR+WL0CGn5+c4yUV59UoU4z9fDMyhyT09lfTH+pB9hqJQ
tzjoqqT5YOCoqE4Li/X4tLSIvPnDtXLWuzHhJtw+8gVONNOYxTXF5Tr642Gu1yLzYSEl8/qT0OZh
zpxEnkcY3F0/KFUXs7XejE7pKd+ZJ8o3VUqyzoToPMBVPiNdeGTfBlUVBn7u/8BPFYKaWox+sebR
d603uZbohmYy3iPvGVEhNa1+BXYJMqpXZJfcIX3AA9nTycAaH74CVou6qY6IwRhWZ8/uUuqN8i4m
6xiI9Uink5vLuHIBP1QFvWFddBanbsEVUmD6bTUtDAx84iK+IbpJG++njZJ5DLGO5g5fMNXqk4C4
rKW1D+PzGk47wMuHJoBF1giiRTsVdN0l3gnCwsUmy31FLSrkQfVGD9Om69U0zo4uG3hOaH9PwCwF
Wj25Kdl892vbIk/sm8lEGA85dnXxRhnYBP/be1motJXpsR1/6hxuF/kxAauIbrCneZ/t0+oLk+AV
DwZDKdPd32uQD1wmyEgtAuBCD5pgidM5QIDDpCAaS+qk5HmuAGhP7+WrWs3KErJobrH7N/nAvxzh
J0dumNyBgPJhh+EXTTLGfFBA0Dga5iiBz0RP7Oz5Ht2EDiUJ9OKtOQDNaGwtQ3bQGwIjIy3cTjhz
dl8P7755JqwgSxLDjdERRPTFEceO+gq1MQ39qTgTzAM/odvYPp/vyziR/TuqEZVA3P7rh7P1PKEW
CROLsBWzHtsZ6QrINvi3KMAVr45i8ysT2up6WglCK0ME+qggVfMjXihh4/2KXGkRriY0xnXuSfYu
TfzTXCZ696bMQdK+DS2PqVUjmITzK2aU4Lnmec11Pk+BgK25dm1a3038wC3eaoKGB1owQFbrFjie
z+9IoNPQAEFAqomTaA98ZMsQnYLPPBS6X9B6XuBkeSGqF2G9PxJQ1/A4pSLDPzCinikfxedoZcuC
bX3gCd7j88fiQYeMf5IztlodRUSSLAIJy8ZGyOZ9VgsjtR67GpyF+qqJpUQvo9FY3l1dEgiq6YZ4
ZHBw6wUzrWKNu0W6Q3b1xwOL15dY4gpDt7nX9fFgjOUlqaXeqQQPEbR1AGyEM/70mqjh0WP7DDmb
mWASLwlby9fXB76yBJHZmSQTRvhlK9Objw/ROIgHbguyLbURszZ6ezYqKhkcEat9NaBFxsa7l4M6
ZBrcYOHrvlhD1e8twTS3YJdHa6aVHU/Zv19PwcrLwMK9vBda+pCSjYSkBr0hyJqZZFD2bthfYpxR
Y0IkkWh/EOYFrBpuocWwSnqfA4/YLGZBVU3q4ekLhMpD1/CjSjVSVvRHqesQPOjA4Hc0sGdwFvnr
BwfuK1nYMn/Hy8uw5qGXAahefjIBuAf1h7+VpN/jjeQI57X7WnQ0m4cRDq6o3npMo5VTMoVxuh1H
Hw9XT5AV3x5s/Gay0sj52Ti7mESQ9uyectyWgbzQjyXDEePfev4lxz3QN2vTGPjqjCPBYbfQuhn/
Rr9I4cp7rzHVfmE/4U0cRwZvL5PjsXIuIaAi8GwqTHkdaEQKrBsXXFVm8zb8Z/jG3pYuO2TPNTXp
G704yF2L6eki/BbrD/gid5hc3v8+8/ewLw7Fj2k7DuSC4RxfRBcotxywU8tZDa7/WJvUX0Q0s715
C7cYfSjF1LWh2yiD3eCKIybAFk6ieUSti5b7HiV+T1NQPup3EcdnDHzHikQmC0pETogkdOm3mkOh
By5q01rXtGe1P33xHuAC8N8gDbQHAXDzyN1XP11rH1ljyxMEuRBMgYzS0vDU1Qns8HT6f93YZqU/
EwmVBGO+Lri0jPWRb+YUovJqifHhWLamvCRUVpqfj6xsblkjXmdX4LXkEj3phVmCerqHYl+Q+X7V
mtMqV1R+i2gfPaLhJlopBrlJZ42FAKFlRPZrdYsdcGgNm1GYfpC/h3tcR9A6IHtBQwdh4QFTbXsm
ccK4BiTA0hato83BGDnP6GRq6OBAU5KH1zpoMLO/h+/9+7WuZiCOWXqfLMHKSfm1q5k1KN9dGFKY
DRhEL64u/ML0dewj1ueyOtxcbx7lZ7TQJqizXMOQoqD/57HtxnCdevSP9A4mXKbPf/fVjoXUT6Vx
tesWnWJdJn5zjZi1tyEHHR9UTFCmod9tSXCHm8NRb0gaM1h14Th+B9tQ3+oGXQytsI0kI9FI//VN
qu+ZCrr+cvfYpSty7W18S252dv1ltXp0tlH6zHesSEi/MvZmB9psds6tQLLs3yCNB61kIFeRQ9sk
o3K90m5Wjea8mfdzPrLM5FAN5rlmxQyvcM+KD8t0op9nhKLZtq07q5W9EVb5GW2gUsD8xvD0THgl
wUFDO0Kiq0R+re/0yXLVJDdcojteWx9tMF824qf7rszXNqjQvv39n40z9jiti4ors4xbKzJv9T8O
/ihS6wak+cdL1AtickhWrDUqtd0GXULJXzkrmhlgH6xNZFkOySjMztWt4rH32XUnQ+Q2aZVaQGI0
YnqU9ytAlt+t90XLfhnWdfGke+JBZHLiabj2eTOAu/pLsUmUGRe5+OBA12xtZ9wC+bwsFoc98scD
AyAt8G0iB3nRQlVWOim//OtfX/wYpKKV23dKpaL0mTM+z47BZh+/DanjQHLZE6x8YG5l7g8Is+ZQ
JK029LtcO7r7nsMW279N1XTUIf4POk1kbdMFF4vK8WZf9m7PcYABAMcnDxHawZwTxyKGHukNJ8XB
Qh/UGM6jKgTY+OKAhUwqOD6LqypQOXqFHbctjGNMyrMwySvOwSVHbghALJjChVcJU2vj6UDmPhKh
CMHyeaLBDtB15Ypf1CehH58nbm4KtOyK5SOft48gzg6R5PsMz1zrq55d+wIneXKa9XnyvCXuuU+G
GuBivYR5MHVyIp/y6uI+6hNpFE9V8qYlAR3gzQQOJhN8wh2RjmJAzLxsfqyavIUXAhAxL7U6Vv3q
YwTmYUCizwZBH/zmeMCFlug6BkSIOsemL1RPM0M74ASEB0vqxOKCGcsR6rcjTnldusSPZuUaXGL7
3iEcurpZDlkfx5yruBohiZ1vEiVtMtCWfLm6x/WcjyaoOIlP2Ry5izfns1JUx6pkhYvWvLFcWDEh
78CXHcwNcfw0AhglFedu+Rq5LAhLwo1Sy9qhVd8CDx2VXus0IK03rLWKTgTX6F81GK5w5rpin+dg
9EKIQ1ba7uezmaX+3oyLrgmtGTfhxKEwkU8LYWtodm+YydcU/j4skYRHU41yf6s17poIVpdDtK1Q
eAfw3WW74Z2PghU+iPKrZpw2C3YREwJTX0Fwzp8nbXAipH47YIapTlMKVSA5pwang7FZkkzRu0kI
3YDAPWJ8txXmoMtCnsfnUdSHYE9VgtrXK1mGTdJvIdFQeXNKOai1Qy6WDLT0hv0bqaHFkl3LA4hs
NA599e0Y/yT9Eyy1KAYPzWALd6Uv1IIVVw3FYZJ+t/QxxxPovC0tQ0V1jhek4Dy+tjbDyQGqEnyT
08Ybaple/m+aUMI0KZ0jGIPJ+0FGeUoghqp9BDpeJ++8NYEe7Uc8Judrhon58QXfzzMMf/xTsPme
8rRl4iWjRHL98omkmpXeURMYQ3MYCFXhvUvXCbclgQrGX+yPTS0pYIuR22U3ygra8ruqooR2oPae
VV61zbgX9TigEhfKLeRSGo6m4/VhCbx5a88d4XutiSC/2aTo5HRQxJKxAH5N5/4+/lYBeq1TayUJ
sOZ2/vNBHAdR+BBVeyLU1+NrXqojpSmpD7ViU8EdcincU+4hR4nb6Z6fOSPfAh6+qTeAFbRJvjXC
JIFCYXJWG6eDY1OZk8fFZ94jC87y3SHca2WrcPWE32wNZnpeAttp+8tZlk3hng3vGsj/PwQgE2CT
93H+ju8RqZxefYjI6GKosvLzu9eBIhn4CQNFmygdLrtitegPZ6gVmrLtFqc7ZR7nIFfzZB12Ex7p
B5rCSttSTHlYMOsywWAsD2AybqhsJ29mg4tcDzYXLpFoyIJYeUT1NWpxlaA3HJNq9g0ICrKywa3K
W47FKkA1qAeSNMz0fV6lkJFXarK/xGknbx0DzrK0VWCrx4lLEqGawRs8nhCJuqFoW415TAqeytIe
QJ4bcBhqpY7wa3Dng8ujQuYXcOI6YQF+mexuLniZwlyghK3CCT0W0Su1LlCX3dqYH3e+C8jo0GAm
3k8YfNBt60w0DHBYGsB1tjVfFpi5L/Sccbn3MlZwfPnrrBx2hPp+0X481Mh+vBjlGUYYJJX5eT1u
poxVj/ZSgZboGC0bEpWNA3DrTtZAqLKWkNLzLlmon6Mn7TKTtIKgv6/c1u/Ld6yEc2T3UELpMojv
Sgcc1XrsKXgeCWBSV/aKsuxL4FjIj7x73830SVuGfGOJBpxTLshX7OxQA8sa4yFIYnAKulJQMFWs
uIcaaCg1rpUUpUUqzYrcW+ip1h3AtkP9w31opiYD+CEOEGvD9KM+2qJVhRuyjZ3dz7fkOoAN15Ok
Oku8H9edWG4ozM6EjVUPIaoX1uy62jnNTc3/iBytim9wf3eq+aBqc5fpS5i7Cz/zql7/C9H0X4lF
+mynRdSq0AOlHiSwKvmwoAOIBQCFSvE5EQTki4j612XeOoD3JdjrsG3OJzjbFfuet3fQlshQNPB3
QbMJNwIQ0s+3sGKVL1ol1Ytl1FYEe13RbyVu8ZGdwFHF3ot7a3RGWQDT2svU2YFA32XgEVzP0BfI
kmwKU0riYqkXDOB25T/FFaJS3Yl22TuyF+uyZshGegxwQycUGQOqWrfr76w0BP994iLWcnU9572y
YXrIrZxPGCzC9du/8JbTGTBXdMUoDrM3kG7jJPuVdfdZ7poiSAboVsNXA1mrOMTFZX3pJpDV7qAm
A+xfaShp0IkIm1Y0hi7mygR1+dUEAtqyB5ze8nmTiqud1OtWMRZ+XaqLKZCmy1vc7cQ+hLuLd2Xb
GnNtYcv+W2jv+fzhv+a5QDVkVFQH6t0X2yt6k+R67Y2pIE0FcGKO8yM2Zs8w7xwXRoNqER6qmQ6F
Ww2mWre0xxdnciXJzRq0Xml8BmnGXnjsf/wSkm51sgMwV00M/BeUx+o5dHNACQGZC9sNtNEv02or
Ark449+LzHsj/nEyPl9CtynmLr27O214oCpMM2nU170F4QqhqXacx1nrOqqkIdvMDI120bT7C1WR
lJ+IDiRuJeftv19JZUxlmEP5SSEwB3T+vlKkGSvhDLw21U2HIIvh8NcYmZarCQy9QV5NhwtLpOCt
ikUJ0dDICR7dKHBnAD050YaLVo7ZC3HSuw5OblBSyx9EjPycp+7pJCGNTcmgpJwCcSpJkgY9bND9
q1vgV0G5hdf/cpSdxl4dW3mq6jciYJodyLxTDgz2kJA4eRJ3b6BdGfyK+16f4TEZPTvDti9IJ4x5
67oBFi98OjHnVWQdJihNvs2h5GvQxEmO5mfrFiB0S3JHe1rPugJXLxIwbtHaYs0QOYg/QkPRCNv6
Fac7otUG5rFz6aJ7wMmNJLxR+09p5XY0+2jOw+DuMGBfvK1ni0mztYJT6U9s5UGTPZMt/zqeoaDq
yIiCAZTHKtq/Wh3pADC7wis53OlU1BuyUBT8HoeilNKZb/WLTUqoMRNMZCORlGR790bFcc7F6KSW
g/2MbWgtZ8JuXy4DCV73HcyuKc1mmtmjFdk4WdZSSvLKrgO8lgEC8W1OD2GiIbuqNob9qHxGUtQN
Q7yC7ZHyfnBk5OMLGG2or08/6YHJkPy446vzkxN/iSNh4hKNn71ZTLmdZpAdxOL6+kpPowc7dtvL
xZR+Ss2cO28CkSxBMe86cSHpGF8FaFVmiKLiolfEYYhCFY2HZPPQDslETf/O0s1r/QFAfdsqdQM9
/U3jy5ePl3DFvx7NGlaDKtGWsKC7bNz1XtMcVl1/qhkUWk/x2EziNXglt6UG2o8ZFBUswxID+R55
KnnSWzZEPHw/40FR4XYBKVJOH7b6tEwBMUuy91igMua10heH5BQ/CcQnbvz4q+MgdXTKDnEsgg9i
XtfBllNKlwCYZ9p564ggoDtkWwf6Vq4HjgF83a/FyaJgkUJEA1HFTVdSFTIRj1PdtbFspNKrhq5u
rWvElvlNHBw18gCDCDZm1pNsiI+VA6kfsdc1UnpNU93CZ9MuT9rudi44UGLlK3YUunCWkgxXBAyA
llInbscBs7LPBzf8cmMLwrIJC9FsHGiqE6oGghA/0Xzd5xnRU6HA6W7I4i3W0I1PqCXLqCtaR6Ie
bgqwnACoBt3qXr6f9cU/3XqT9OvgRMlftgvMAFP/f6qDw1ykRqleYadHDPGl6gILSqFD+418bjhJ
ZgBdJsyoHFHlHztLks5WOWDUP8VuMCtAaX1VVzMYaymOdtlDYW0sqYuYDSgvfkVuEgIfTnGbGHKj
PSi5F3pnLNXVTNrnBmuhIqcoGPXDlJy1x1IGVhborqN7ahrqiKtlIpVgvzjawy7esm++fbIQdYkC
zgSLq+9ZWPy/Mp2Z6qfLn8p6T6hk1dqQRWQ7ksGhz9wzMwObx+OTAr8Wv77vLduo6LFnJzwO5ZXs
/r7yvIh0sxdnMoG/pyBsjJ0vv7k4BicnzJNZIy59PUIONJS6eSFaG2RH81vfbjQxsnDqpaQrYbsC
1M1fEETtHzPjq9vbb7XKzjm9UeaD1BHbe3eNZX2w9NBD6qAaSFdkpi6p/M1oR46SKnvvXL3qC5cx
ATIFBrJak4Pzy4kWcl81JgLj7bFYk2yPhLoA1rZtOIbwY+zmxMZ7XS+IpA7YUlRyedyjydQQiAwO
XE0FVlgYixqsUWhZL4KQLsL+K+kQ4R6UUAeI70xtNmwVS0hFO9KoXrqJOxST4YrOxyZjBQ/eBpRJ
QDRyrXFJO3ng0xk+XfLjt7iQiSpGmVG8VfQa/KK8yzNL+5DyXdDPdRYMYeMh0sFWSOrlU2ILyR8T
QrH8rKqsb+fPBvtnPi90chKAR0VgWFeVj+q7xOAJVxzKwrzHKV0ib8QdmkoPGBOsZaefw5CIaRGN
oniSZSh+PXGpGymTHimbsHFVn2rOEsT4v8zPoDaUfNHKqOR3wR5sL4yHY9UdFNM9WErCjc+g+0h5
E5l59NuzNnBvc4agYHP3eB22kLfxNwEFpLYrS9N0PMdVYy/UdcgnlcJrcDtSSdFZBjEaV1MPw9eF
6bluNz7XhxHU0f9u/vuUqfMGLYOtBR75OT2IO4FnnciGMbDN2x0gYU8lnlBp9pfbz8memFSCgrl1
NzzM8/frQlEuls94Uv/cUw4rIWZSTj37Je/RQv2/2AD6TxyGjKY4dXMhYof16WJDnSxkuY94io6M
W6NAuDn9Vdr7S/bc0sV2PL+XMKzCicAs4Damni+lqWABEswkU7F861rgRVQXfZVsdv1ARi8FDWNc
0eHQ+QiFPaZCNW8gkavB1h/75tcETl0LE/3TyMVpNdM0J7YukTE2LkIt/Nze3bvUUANZ2AWQU3bY
PxPY2v+K7DRlJxmV1j4f0tZkBtGLQpgWX/2OUEjIY/sBe2Q5mEv7Ha7+WWTmY5h2Huc0V0bSCbwh
eXjq/VAsRrKI8ZO9hk4v4vA7kTYSKaWPm/HZvw2slIHNC3QNGAE5d7OqGBqs0nXynyrU4h7sSu72
GUyNAQByKLD2zjcMAu6xI5wghH5Op7IgP8rWKnWxWiASspZMOJYX+v1oy2bGtWP+exvisBBIYsux
L2kTgqsMnjAKcZRr/RWuzzF9ys3uNpTWChXbLenB/9jbqbBltQVfN07v21SZQ8ia07ZS85wgTKx2
aowEaEcQc1l4QzNtW/njNOf2XuDqBS/DQpXdeKxOMpoWxBz2fVntrEeF2Vopv+ChSHpazdVZx9hf
yLXk2F+pAq2cEKSg+ZF9FC3+rewAAUmLkSpiQ1E8wgkeCinezbcS31rJ5He6lXzQDp6nzV5fEd41
xgINMXoMqqyPUUDXYv0nydnyz/Ltl2HR6ZYyPVjAwC/1EC+cA0LJujs13G4vpYxGMcs9BsG0a3uL
uz97AdS2d2s/eXtWW/t96eVLDI60B5HtbtbZFWnRU42IEYcIlN9wQGkeAwKvZ46h2gi70dFhhul9
Wm60rB7QjmZcrSvEE2joy8gjzcpqHMkoroAgqn235IHoL+Mmyradxis/0hgtR315Y6p9tMYIRL4/
74aB3jiz9zl7TioHgs9kcZp2ZjddyXa0Nkbnwlu6II+2YT6/LP8EwdMTjEUQkm/h+NHhxwqKBZkH
kYY1ifTKZf4A2yXiwReKbzXjZcg6bceGr2JCRywv+oOxAlb1x/KYkRdOm9zz9HDOPNwQQnhSD81b
wu1iLnwLUg7lfldME06DLgWfpztEv7uHri00Zrwrnw5r+itxGslGG3bo73ZT0wmA4aEYyQ5K7lTg
YUkUtX1zD1Hk94Q62roErjLLa4Nnsq+g8s7RZJKZtkFQQ/TclbtZB4n38++FVAy3qLRQTC13q66e
D4Ci6cR0tVRur8wBFGo7tqQhtAhCzzRh7jhbzDaU24Qy2mBGXSk6FVcqYktZSLJHbTjXODYMzQB6
6SoS/n3pZ8fAgcQiJVaAkr8E9qC9TEV6Wwdl8fFKcdwB+XZYkL8IVg52DJu0aWXJ3L1+ptNlKZtW
ESfJiPC5g9z/7h3JVDyBIiJAiVQcyYoAREP/9/RIUt4YqSBx+proZc01Q5IaoFAafgMRV/Csdd1p
AmdUc6Z0AN0/ylAjbzA4zdr2L4e5ajb1NOTTpaVk9xA3Fx6AJR4lwfCR7ueuMg67aKMtziF2j5oY
3gjBpYS2CiWAEaGmDLCZwI2gb3wUgXmtpvV5r4/ZaIq7ma8GWv7bXPEwat9lyLnIc6vKcDjqWz4R
2mTfgiGZv5NEtj62ks76q0BbC7UBHrdEbkx9tDzYu4yPj25Hr3LUfE1Iu/WK04rt7kUQ587B5EEk
mDssWkULyOS3AmLbfqelWCCRK20IvN8NjstOuXsk+roKtua7dVLONSrRglt8pZBxYsousBUesRA7
PQdEiLGFdtF9reiBB0H9ESOVOiCCxqSFzkIz77uRzsjvylDMlp9OR8ZC8Xcw93G+f/qqgIWR8Row
L3HFgQUphxhrIIxGvDHE3PWM4rvnLd4gC3p5dc+u+OYtQAQ5/S/0KgmNplP/AhDaMreOddwgZ3O+
5dKbRowB9E459nOO0M0lQ6oIukb4QYRyruNmCGwz/iyHZW84s3tdVFr369O6X2dkcsOiSIhBCWUy
jBrrIMZi/uE/YSPzmN1QZlMaNh0QC4zmjcxnitCdHrxlGIHdyJ4kG3YeV+N6wARXnbXZOvBi8WdL
IgJCOnliwogM542i1ETIVZrAJzrBegQvIi/5eB5ekFkQC/tkzQVbBEuQHkEi11RBp0KPw9uVCQVq
rllOZ9TKWTQUY9ODCTpLWfWKxqEEKCRG3uLz0gCAkyeSQyYgtSFbiM7tkM/yhX253eQpARGZmx+O
MsnmB17ZSH1yaYmmkl2NoagHUjbc5TvD5MXLNiPLKUKsIROGQA5M31t37Ez0LyfzBfFEgtwxmDCk
WeqEQx00xgSy9UfW1pg/u/6NRmTog0ufy2R7YznUDXnzXAMWPGAI5c0dTBGX+9ByJU0pujviPu6t
+UilRHpqalk69zUZ77CIiEdt/Kts9au7Ie2UdouCTei+1uxO5KrRnzoZMG3NWKDiu1/bBe5h98mA
MqwfXXrYoBfA5U76jPibizwScuh18ZybGWzZRSsV9Kns0w9a3LLVoPaLSyEJakbgNRm9Vb9ISwJu
KIX9TeFjw8To1yPs4PSneNdphpl6xcdggbhxkhK85bKs0BFrSiMfZ+NuW4NGOc/A4NYOQZqSa7P8
UZEjsCFv8NA2uB1V5LTrnOD2DlgoGp6RFJS2JhKV8SoerPcpJXAxZciG49EW6twZB2aavamzQUOw
3EBMPCvRzq8woWNiY1EyQd1vTHspLQPrXZNLbFhG1nMMhpmQYDNw558YgOrq0APobTAGJMYBfUew
5ruXM4YT2I+9t2eTMFE/gaeBBJHhuq2OOUxLsgoW4lwJSTmSQlk3XyIWv25xmIhay+i5h57A7dgM
03le+LJp9gSY949To8Mp4DdzQNfHPOjU1qtks3CQfKZlc6jG+Y6L4uTeWvTAQsFt0AOnK7Es9lyC
Pk1hhyljps9tNncs3FRio74jxCQ+nkDNpox5tNGWnf8g7egwhuQOaZQ/cbY3Vo+B7zX68td+nhqd
ZWDlHLNvfr9fx9en2KuoiE/DX6bCjJPYQ8fvb9+MsoKG4MH+lcB7hTzC6vfLGGPL0oqKR/cAXQM7
QPwSHsOU0gi00DB+CjEFsN3tKYwgu0aaTIl0niUPo6A4zexm+6Hj5dVSMiUYwZj76stccb4YCm40
1qe3AEZR1ichRbHwGs/q+isOqO+QTYAgPazOYWm/wX3mnvabvcDp2b/jKHwFOndN21y7B8QcIvat
ysJSfdlEzPxXd8MP/QbZv6hFJNfWY8v7ZY+W0ipFuJqyPtDyGmXQVCaOZ+ZPHwFhACwZHSXJP4hu
+o8fQSKhGOZ8xrVEiIlrgyotGL+Pfqt2C0c34DWyiV0vqCzfXLQOhM7zibB8ulp4oqQCqAK9PydE
loPZWfay80ahkG1aPNDzGQ+pZJT24S4v8Ezpb5vQy/yl8bXfYCKwkSLbGFuMRZaIUR4F4pBuzsr5
kjjPxRe+IHd2L3vGfpfwy3YcCOeGsU/Mc0gI84RjwQnj90CiPmbwAS4iVxkgry6INMyc0fI/GEb6
zDVlorZoE/24nLt9haXD0Ue7Cj/0W3Qg2w5/7U5vHAQwHchxDmq0lLYOqplwEah8LkflNwD5cVFI
2uBohEOVc6snzfboLGXbeyEvVvwHb8lL8Un6kdN5jhwoEWefELxBFbdHCcwQop+i1vxQrws1hMtd
iN43xx6mc3W16FlwV47vLYDLeEhEMSeul7xcjr3Eg49FYZDAbIyW6POkEdIofG+3En4HoZvCcFSV
WQtsHQ4ZqeTQAWxRyps7iTBqHQBqOTBMwj23/i99PTbk37DsXHiFow63q/5qZO4UFWUna53JgMnH
e5sdIWgA/Cf4S4Atzc9a97aguHfTcZPESiSgEIbErnAVcDnMvi4/3Y+iDXSj5zLsOPZR9RORbjm9
71qWsR91U6N5tEoXiMeSyw8JocHpZadqA4WgpR6sW1cD+8VyXZwmfgqByY2Ej+8Y6d/DEPvlLdrW
KN8uA4ErK9h+aZmjEkVJiuHbmZMINFwVBhEcVjLw39fb2vm8qzXCcOXIjX3YkIMsVjLr3IlWGPaH
VF+YFiYya/GjIuzNbr6If82QLEgY/98GlrFXZ3QncFDrFOzer32l3aYzqzYUa2iyq2J4m2QBmr/s
nA0CWaQCuq4UkEnChxv7chSN1HaBrxsjDdqVXQcb0qqLugK/0mFFgi2ptzBg0bta9NQqcYplwjvJ
TxIB1SZMgLHhnD73lN5HA2vuHVmPgQugG+wRq2iDujg16uxY6jVUrzjuHtoLQGT9bttcLFt/e03I
XY4JkosH3CowybzHGKp5hwbyqFILl4erScHuOuAqbR0+TTBzMwThKt+kJjqxAwHRWK9APOTSntkm
N2pwebkFBX5BlXD3dbKaoxua61tMDyccXdZeRwC9FeVBWTw+LR5ksI0gvXp61UWUbYNkRlKhsoV0
Mh86BCyC6WwHqFRoYpE7U0rpvLXpg0Bjn9tAQheP3+wSTiRyyyNYACeSY01tSDNuwnzJlH7da9Vp
bxfbTak50UjwLt7Cm0dG8AmPKWhTN45g9n7iu796rURCkLzPSo5vXokoQEBbA2j3BieLLOQi+rig
Yt4gy1hsnIJxf4ZYA8uv+ldVMlYWUi/M2W0197ysSBOWqVpQfK756WqlNYDJ5hSAvpdtg4WFSnZR
L7i1RY3NMCe3OTguST52dlnMqTj01TKz2OeepTvL0oqCJJgbFlPXril5QjzU1aCOz/A56QWP3CYO
f859BW/xuS2LDg3I5XqwofxNHYXTR8mYPBQfNhm/mrfhVhCKCfzPgdXsf8i+JwivXx4UWtXJARVP
Vy8paBa/yoDSgxzEMztethxfkJd5ZjUCvSFHt5qUK/J1YVxM86x4gI7JbBJe9ycrMQC3P08qFQSr
cWhT9XpCGFMcwlfkmM3y3ZhWtZHkyT0VvMX6kp9OWuCdzUaDO14yVI/+0l8O/4kz/tRieX8rtyzs
2QAcxe+wemcQmVQq1uYHEZG8eWrlharpCEMahhCNgTU5P4X6GSgY0N6K/uB01TEGeCdmFnAJu5O+
WQlPdun/PdxO4omlOY8Gmd3UxkAWu4ajzEdW06Im8/zmAdm4Mx8hrEluZoobb8YDFdZJ8aBqv80+
dWl5Tde9seszFvwuJu3ivpC14wX3SGSu85SPnP7RcgJlmyKxDmD9GSQ60+rv6wasRodR9+cz25pG
s0xswRMY7jP1SWkrJXkVWr7mLUlrcX9ipiIHga65m/GUzvIJfYwStPCKddLQFWcDH26Siu0vlhyX
n5wPIBTqoKe/uSDTxNSMXYVxcMV7PiOWCDuUN51eRv8fSy1286xoBtqpH4cOswM+ugagNhiUWN9H
2Hv5woAPyXwAjx1/JyDQ7dfwNo/sNPu1xnvD3mqIfvATjIzVS1HfIBlXaGX68oI6a0eGqRaDCLl8
Igm6wt87gbbhALiUB3nXHl1YrKVn1icAZke1CO4dH/9DyB+njBZna+T18TMyTr8FUWjWK7dcmLpM
cVPa7iErMfqGXWJo3CaA5dbjLI865rbKzk0IB7S9pC1cgGbN2ROP41KAW+mPumsiVl14ShGTNGdL
dZoAFCp7vRcaHzYkgtQab84yP62T4tVoPM1bu+83s8Jv110ItIJyTydfdafU5ViBCZcS0sbNIol2
qM7uN9ceXqPMkJDrfO7jjCc1Gn5A+Itx6GgmCLv3imVEBBMbS2wTssG7xhRwWkgwWKhfZRrHyX7U
GgH0Uxsvr2adAF7JCLLMEElM2bXgyAKgXa0ozob8WRbn9EKPJ05zL3/JP81Zvk4NTUVuNfF9uDt5
YY+/lrNTc+yrm8fYRwXdMM86HdRCr5aT/KCuzlu+t1/dzwElNwsk/U1EManq+0bxRhnN8mCSR1j2
r+QZ9MXPCBHooyEgLYVDtE2CC8fTlv6UqWXNBvRXJWAGYbQjMXrMeySYiy5us1c7RvVqOxrHe+OP
7kc97uDjiteLT5wX/ykK3BFqhx+F0ATu7XKzjR8o8wN1zMM8FXTE8tJuHNGlz2qUGJcHv8VsK5tx
fe17VwZr2S/xtA/BWn0GSEj9qMMVQktGBcrRAODbwRJNAYCBgDe/KO0oYQYJiVReZJKBccuQAFGo
kKHfmSgVoIxJeVIR3CJFuJwDq+GO/s62ekVnKlrgCE9FczcqF1lvfDodTy8/hBh07MgujiwCoTWU
6b3CRD/AQlgiLtCcx+vRPBjHKwWyF1X43sJIjDwQpl42qK/UIWFUd/SDLTnzRh7dCRWqYxOc1kR5
BwlT/Cx3A3z3/5YQbV4fxkoAi7JHChX9X9kafb1VqIJOwZBI1tq4hHXuu1R88TfD5iCc8IK1K9Db
wokpqDfwEYKMuDIzXPORpXSiRUTCekyPeNz6caw3R6R5KOGqEAvFNNvppbjW7Jems0gKXgD6rFrE
vIDbmyPUSSbL1HFwr0o7hgKE9TD2mS15iqiMPBAKqcoEx8T1YlryDr3rJEyaTzPC6ZEa2g7dVHe6
ez2eELMMnxc3RzWTm1Jpza3HP2vdcFARTnIgJGwMHsAbIOBNJVOPE/7uYWZ+Gi9xv+mwN2oCi+R4
xwoyNG/Aqs/b3saqks5Vb9zKYxQk0lWxIWOrKIvOBoudNb375EwSQmmsvxjbM0hiHE6dXg6BWvj1
pl4txZFqZLQG+vmzbyo+9IcDtAePrZ30Wg/MDwTNkkSxvm+IZPWMBj8jFf79MAVp8iHc4nJEJnrL
NumGaR+enx1uWU3asC1Hds6htlcLi6OJFNAgYe6aJedyBxlDZuiCUqUCAyKy/BUpb9Z9D5t4X40D
k8yKPWBFTk4uo9NH5UBw5f2sQDROxqTon4hzzh+vYJPZD8g1KRZyp9+DYjqknZcnGumrLUi9/35d
NmnKh7KECw/vT/kkdWOJ1C/IRdfi4D7rRDegaGyaNzNArPePr6SLmIK0ruRl8tlUlYF8j2E0LkIV
0UsXUSN2MTQxUSkHaLSxLSz+wbrTAXBnaR7vGBfxAaBVPym3+bR+5Pe5k4vwDmsiCcwCw7fKTLxF
+zjrojQfu9iXCZb7Joj3P19+eBm9J7ufOruWx3lqPGPzBZ4i4jaQ2uuEXw0M86RuTMT9hVm9hm9u
Ae3iv4cCJ1izPwxxHV7NwwAy9PT2wh2V4y0JA3xTEZ/1nuedPJ3py/drU+ATc+6v8/TQmY4egJRd
x5CFK6cG4neC4izEWKuU2AN1LnpTjLIr9PMh/5DcWeOb3386oHujGVeF+lOsKEWc6mBXoL2frTCE
O6kdNPSXTrl+gjXBF5grFljAUoxE2+5B8pYBcbDMj3DxtT4dpjIT6DDCICtAW0ukir0Oqu/vDKfp
5F/RZkWJsZCJVVzL/ka+AsDNIEsllW79XP1OC+d/CswGm/iAAI7IU4J70nujYxb0BVIVJd59aE21
hpEjpk8ZEmRX1t0c+UwxqBabJJzSO7xxz95vuYehd6ibi7WeqiaiNRhpPDArw+n6bT2L9ohxAsCV
Q+dTA9QR0Rnuc4XnfvjUUGka15QKRyjcvhLU7EKk7KCUVeQ9tF8e87gne1M2Np1WAiutxaJE+j1i
tWCHmapOPSxIrJECBCJ39PITMsUT/zpn5xnBQ8MK+8sTYCLMff/VeAHsumai14WKnMABYa+rBBRU
OEllVDzLaI573hYpcwheEdvn3aSERbD0dLcqXo98qf7ENY7KtUbOXUtgMWuN2LAxBglv43U1fv4+
ew2EjmnV+QiVFlWEHaJwqWFc9kMK3JdOPMTZ72hcmrc0p2yHuqvaCJwjgDqbVyVfGpU5P/nWS4Rw
5bXfSmyhm/kd77cSxyl2hTNZnjPmIFneJVkxPKCS/mQwH0x82N01H276jU43VYjtQF9JgYrfuFsZ
fyYTvSXfsIxYs+vTgYeD/K9SxEVyQr9018H6IeCqOBL4o906DfHU1nUTZm9zHx/hAAx36Z82O5RA
eTKQ+JabTy870s7fTjim2hO6CYcwhhxAbYvw3OHNGVLAnNXt31XCOhrzwbCqlUYBIAktuEqamjgM
EqAKqA/VhJBOxaK/jrpHObHE9BmDiCTvtd9Jfb9vVwhMIBvqSKMUinlYCxl+k5G9fTeEJtH7DKYF
VWNGeIwqdAURrD259FYG8dpH1uOB6Rk1n2SH4oqjt6TyrDnFd16sFQlmr0JNdFaz33Hv9CPWFpXw
VWrz8fUt2V6FRvE5BK2ARI2x1QDfuzb0+/UXqh4a24QkNMxGrxNis5XIF+t1c1VK1OklD5RFOV8H
HVvulGbfUEWHHgAuDVzri6jSjq1QIlAHjQV0s0NXsLUfl998o88BIxQjr7GMJtmT8MncFJktHtgg
VDUnZ0titvh5ns9h73CkW69STaJp7xNyDQKyJo2/PTPt6ZM8EzduWlyENhZYDt7EL/RYiIRntAGS
afYk8tK3wddhGm2oeflL2Is7dXCF6UuY+rHDmUxCivcxUSK48YNeKinZG0IaeVm/+MFDWAnyNPES
QagnI8B5ffO7ye/gxqHmRnDVTDNNF+Z0UqA5VxUcOzRBgsbGlwTUExT3B/LV/6z2BybN0rsE4IYM
gf1sSMtU2EJFNDJzOS25EeXplRGHUPCv8QrCTqgbjMH0MTo8Wi83/vs6rJkAXCZY3Opce0DhyFYM
ADFbE/rXefXqceCA41oUN3qA7aXcoi5hwTaf8HrKU4TgEKtXo4BLa55b2FobkOZYeX6hVTfWy7SI
LxHML7JsWmTW4+VY8eJBnylpCc0qC9D9BFXPTBSqXG1c6TqJ6PfA16Rmrmif8tThCV5BH0WUT6NA
oExxQs0KJvuq0orZ2bWIOlu4yEMBGmXTwGxRf0LYEbJoRrV1OpNEx7pknMIXyGj/8vNdulN18/JZ
2lsL8lXhoAlVFloMEdrYz51zW2DEsw1UXbyHf4NzLkIy+K7TcvpMvuVfJtDxId6Bho7NO7E7e1wo
wuBVPiVYxTqI8rtMEeaFr5Tu+MChRQSmwhp6tzdoOgArmz4qVV45w2M0wVQoW90su9UidKkt48zH
FEzEBCY6yu2NBLIg5iAfKfBC5gimprgX6o7rTfX258/P5d6XhXz9QN2+l+dLyw6StTxmr08MwPMK
RbcjvjWgQt2TcnNni/AvypPN70OifAAhMNEEyXJBz/gc50499+y47Vt9A5SSom7+MG7OIAK3W43Q
GRlqRiitP6Al6EfSAXOQEm7CCp++lLx8OWIIlKHbYHU42v880KfbwjpGa6UhMgmH6wPYz4jOEFaQ
eC8/78F+WJp2T06QSV00BzMKopKaIchoa/yAqkLIL/ieO3ZhkVi+Nn22/ZIqPgYOhg3stPF98d5m
dspXNoDObykrjYD6UbwGwpS18xKfjcm1YFTg/R9jIDOVN7/R02thSRipVnuxo1UOuUrdrCSouyyv
jDmYlOOLuQnjGBUKQCuqL4pEe0zNYXGGeyv+J0fLkxqHuiZ+WaFLpMbQg3cH/bVScgEceP4MsOC2
iuC1dnAp7/4i6aiJ7RhVLyRsGjwf9JggwcasZ78L7jugjD8SaGciHR+yivBRLZ/dcPfY2Il/zRrl
ePkVRr033Utdo2HR0rzIJZ1tPDpNeYma3vOBTIOiSMNAlu9f9OoYI2bK0rn9EAMAE55k48/DXOji
nKWx+JnpVyS2kmq5BUPNziOHeCNrBaCZQwycKKvXdQCSBylWfru5U9/wGTDXTSdbfKUywAJKFEnH
PXO5jDaL95Y/2Pxls9i4RKo4WWhA1DEWb9bv5Kt6f4VSPpgHrtzQNTMyvu4SIEy46ZhL/OTwuxgu
nn4pbt+4v7WItANwzQd0QYRHy96Dyux8soruDEnqTXzFt87r2XLAi63M+X1npnIUkt/Ws0T4M1os
qX/bY5S6QuTsF/Fe5rMPvo4R3LkH4GvUwJHoK7+STPqVuE4T8z8orrSdvCPULH+HkgoHCoaOWInS
pgO4ZCk4COFkVHZh2So0G/d/XVVi5ygKAnFwmmnUMc2adt8RNi+9A9Svz+NGt/uE+XHX71PH0WG2
gMlxQpCtxYWigsMbGSrhcNCnAF2iSJop7KlmVWmCDh6LbEB6KdhObavbryXjWWOBZ9p+fUf5tHfE
QM3az7QmJXWkBSHLjtHk0E0LZeoRe1Wm6Et12+THKqyi647ICRY+k115On3qGQSzmWhQzA8Odj5M
N9LcXzvlGW3HF86wGkBd4E3hnQS2gznEYv89MTheJNFztTPS+InxW+DyRpYtyz2sce0/MHD5IV1+
F/nsP0NdF6D6M1gvUKxm4TD5vmxGRIalccM9bSt2VISHfDMxwqlP0hwtHQoO0y275YNH3KDxi7aC
57X98BoGw6TYrHWkstKllCwp+g2R/Jh54vjxENcfH6YV+jqxI4LgIZ/hzoosCRc7SF2iLIRAb0fo
HYLWMsnQ5QTr4El52Wz06TiMK93H30ezt1dRSfm4tCx1RURQDDUuj60+GGMswuuSJL6rgvVv3HM1
ocYX6A/5+bUDxxoHjZpyVhjn8hnKlpGm7d2iaMd+s89GfjpMOE7HRa8Apy7F3mrJ7x7gUdQa8Rmj
R3f1kH4Vkhhqn6pKfHlWAXTx2ZE3F5SO37UeLWgFj+Gup3RlumNh+dhvTrkfSbfyoF+fzEpm5N2y
YZHOBfb+2qWoXEqlpIiZbxYevQGpKEU1JK9fyT6rDQ4kpAL36rfKteiPGhRZ8jTJY7XWmhVNlQ+s
PCvjiqgSAaIAvzcaWAKi691h4kxh0tZE8yLYcp2rrxfYihqm85r/udWS24LdzsY2r3UspBJ0hIy/
AToPQ6tcylSbfDYGOQyg85mtHAomIMT49f+DuERcDJeX0jB++/oBUyV90OGmGcfNpbItiwj/paWE
mDnK876JOcOmhkm/E+O/o5+Nu/BF0E1pfa2eyhNoDg3XquGqVlSOfyaojDspUee+8ir853os/09C
O7dAdqGyedK5IzuDKYmynAXuXJLIhjbpevhob34aEPV/jrbzHJP6ppYDN2wmqjThFZgmFZ1g+Bt6
prbYSdnoBjk4DW0kSRALMn4ny89zbYnrn5xJPGLduWVeCg0EcOILu29p1myij2WPv4XEE0480PmV
W1mTHcNn1mjBLns0bMbYPUAOBHOnoGbgjrQTuWXbgH0LvbQbW7XhPi46LwEt+Snt/0cSbT3vs+Oh
czBs5UOgas91BiyXDtOZ+oDhv96QNDCUYVnKQvV+NGxqc84Vkz7bbse6Ea5ICdWN1angPojt0uXJ
rFk/2gHmTav81IHz4TzIRvrW1grmIPqPAsnHyKtc4Zrc+OGvOAYpJoGhgqaax0rsHNAv+SP6ENJu
QOG0yfKxlVpPmB9Cgv7E9k8hu/nOxxxxLRqPUsf55mDQR7GfJHWcx2N4VIYSEEYiBkT3knp03dIm
SszMtydsPbM5Jp6jjY6ksUeYMCNmR3uS2kbq0CWFxjAs8K/VY4uXfsXmzZmtjefDI1i7TQFouSLw
n2YiQRbdGywPEbiGaesZ1buNVN8ElWVwGPVRPNRaBYU+yU3WMYMFgrCGFJlHlSztZ/b3PgXbDAmo
KbQRFoNZAmTsV9H9T9hw4IHMR91gdSj1wWW1EIVnfX24TPBAbhWXGTuiHH3gyLnbLpqkTjnJHVEU
Dg++TAfek+XXiU8ZUakfExntdhm5KED3ILFlrtaryCWP9mQEnOAxCXuc0ddSr0VCPAPLE9rbSFOm
GQBm9SF61tvTBZftU+9zF3hECU/2C+HKsO0TU47j0/x4urLZpFEOtYp8pacl+GjOuTKe6ZXh57tE
DMaR99x1MyohG+hoXTa6M4r+W8g7vJwIgWGGH/x7PPadVOSBaAXSrWS9rTZqyVG6vqWJ4PnCV/st
gkr8Ziey4U3KdEQXkRRL3tdRQ3WxfH0uIjkjNeSyvWc3wwSNvpA9YhMcBdBVWFpJLGgS1aQh8fST
rZiDYqr0ShCyhE+n9TxIDGGWJY+/rYzIPS1+19BQQFp1JYL05WECFhf06L2MJG65hvTnEHLaq1UE
4DyhCW6YLxbN+bshxVeLYWoRzBBDSmZd22ZqC4v3DIUjPBzgSSbwwytAkohR24RTnCwFw9g3Ljce
dFVHCWS5W52Pb2k62QG1IXESaWiTFK2B1d9KN4YV4OEXz1SvnWvf2CUj8MRyrlIYBgX5VDGe9xfN
wQdpjrXgqSAEvXtgv3zsNO+K1mF5BBGhyxaVBvO9BCo5D6jtC31IrgPpoQ1HHQUnBqnI4V1ke36/
eBdj23+m+MGaLoRel08gAc7UqhjaRQcpbQ1Y8S1P7gRXizywvO6qYAuMrMVaBgTkpxxPIsIOdJxg
bqml73yPK351qoZO5ZE96LGBh/ZNXwBu3AWKDKatE6eoa4sIMbxaX4VbvUP6eU/D8N8nu8aVIUll
qFgrI8OUbmZ73ZKYk0kGwFJ2m6UFBtnNyR/O/rpr7QEdqoyBwly111WJPqo8EgXHsItUXP8UVnL9
GFmzGv7K5U7xn/kKLMvtx4sgcwMvNTQYjBTnhxX0N+Y+GZR1c+pK3jfN7NmgPx43ufO8Eg7zTETX
wtR5S5CYS3OmuCKScnvuD0R20mDzvm9FonE8My4C4viLsGWNlCQZj352yt8sgMaIH2sPe/g+uBx6
FMSWBsyur/HNXH4FlKKYksVRUjbrrvEuiV0MMDzBzOA8vSNWSSdNNqB6AMYRUPTQDrEpLd7RTDJe
KEj7oxtUT1zUv/rj6NebFzLAFZ1Dki3R3FCApuzWvUJNOyKThIjVqKzeDfPa2Nj3jXrHzObVaxjg
JzkSRAvFrjXYUwbd5j9nCIthL0qB3EuttAI/POLnb4YXxsbXk3PPLH4r2e369mHgzsAgD4z6UyTx
55J4iFnGEpildXKwll4H2OjWjPL93DrnC+rrOwJw149FK5YhjXW+KEHtTLCXmdNu8g1vftS3e63n
Fmucr1WN6dGF/zqcrBeEAW8wEgIRX/0eBu2b2qcFEVfF1yhqcqfZXv38+11GWm5V0ORJzCo+esis
7H7kRfGCf0IsqRm5SfbDsj5CIyWIewstXtuoeDWiLWUugFuamFqTI9y02GJTG5Vw4r9UmSEnh0k3
pHKHz7obMpOugwObnRp0I1qNC6W2SaHGs3WQSdwjFRb+lCOYv9AFDDtpWbSYJ7RB/4CX91Zbvq2D
Y8zSnVYgQJFUYpO88DK7FKP8orrHe4ki3ERC03/t5xgpCSpRPg+NHM68XnkqF1oODJsQfMK5rif/
/vHK39KwWbgxJyR0ulgw6oG9tphaVgZYWLL3SsNSuJvlJWHbzdZxwNoPvr/mrloTZHFR3YteenD4
n0rDoO4mHeDvr9muD/Pw9F7Ox4XIftWZdPaBJdtKWoZtn0GF1ftB0RqSr4dVhVFogWwYIN8to1Mp
Nos9jdJDOAu5X/QJJIRtxS9OgqQAoW8bMS5HEXmB+l2tH7/xl5iDZsb/jQ2R9frTLcvW1wljayML
2XqGyDp6vHhyRT6pnYRnhqKCNQIjDRN0CZA+D3ku08JGPsdHIhqiwL1AxBCwygk4+8zvag5t7LHB
R3aeecOggpFNrouAtK61kYU37SBuw54J/J1l53N2zuDApt8IY9MctYLzuMVeaTpVgnfUNc1gWgA3
40+/3BuTGbAYaLkcKRXad3vMD7S99XqT/q9MkVfUHT3sKb30pgtKAFFxdrgKxpNaA/bkEZApo5w9
skzy6SNzibOXcjuJlRr4MPxxCBZmzwXy3/qZW9a6sJx4OAVCb8RIojlo8B38njxDjqADEqsxVfIE
e318MACdgmcuPcUGEsWZOqY+GlXyiOaLxrBtG2+dd2oJZnRAUlvYlBAg2l6AZKbYS0z086gGMnb+
NobGvujgUsUeSkrXG/pVpyb73j9Dy5WqY2YH43BeKFISZjOKJgYoJZnddmXWN3w0Le6TJQ8bed1M
SR4gCvJMSG8QhTeSWYT0vq/IEprAufid9ha3FTR4HXvezWFcgmB5e8uoqKG52D4r7Z/U/tyDFiuU
9LHUzzZUTGrK+B9rO1oRrons9dQps2NU2i4MCm7GE7blwpRO1nzkmgEcy+EYLru1AwTa/2YuX0uw
hHGsZOcaxOEPba4Rw+fdlWxGTIJMlFXHaJBnmel+6H4/68GmbJOTo3a5b7VLW2g8QzwKYKlW/qIX
vlCl6X8Le6ngOpFxC+r/OiTc1/WAtAqD2ni5MDh/JQ0WDtNlqRG/SbXBFwa4jtZki26EPNLSxQr6
wNk0TLplD5q0W/FznXF9U+i4FVmlqEhPmMmPOuw33IRLfVJ6pKisStCgtZpM8CrZs75oDHvSQRWK
raOFDFthekuIydVr2IeVOP2d9OFXgNIHOvm4LzuM4YV6PVaR46stHtveZxoriJ2h/lv3ivVIBSGs
9dMCFHI9G28PCMKMyJ+jBIznu0okvhap6BORFcl39loGrw8TYGk0xUyumU0OUedzg/S7G2/1I93s
d4bYEeEtqmf8eznCKEXOUgAnj45qphgnzTPTsQ2scqZjoYs/6TH5och2HKIhr8jb4mdsVKO/VC9V
vY1IQzBrR237ib7A0wqCGqSqOiw5dAhlbz8coZPR3T3kd13CByp/mVCI4U/FKxYgPZkOcqOoTldP
/V/TfXNTOkEAnKm1lFKW04m+LlNE7K6FenNWHkQTEGvdeLFFIKTlYCu9iXjB5G571TJJT6nz1UG0
BFv/CBXA83dN+bXrcmAV3+Xm+0yGPeYq4JqbVBhpiX3ohBiXdHsJPx9FPHxKWLixIMxODtyApYuo
aT3YFQT/NVg9uI6XjRw6Tg5yS1gHqjf14UmN+BU/bV7F7QHGXT1k2E07NWfDyT4yB6CgRNsNqwbV
ld2hJhT/W/JHgFXdHndHYRDK3TVAMx9tPeV9IuVSDvyC0rBRdHNFTHmi/1JqkI8zxsJy2Ih0ysmW
Gt7I7bltj9UQNSKDTntCfQG4batva9cqWTASpU2jvyxK1RCKUK2y+vIi1bb5TfqQgRsbdAxGyYCK
Vqle5RLKjZLovjJu80ks0S6sWkHnpfS9/nI8iFSpoOBp4JUb1n1V/E1sEKuixui6U99S6fgGawHD
M9FfjSKMyEYf7U9oixuFEeL8VYNzpANn/DDnlwoZL9RYGCI0oj81o69CRKgJu0gRpGE9H0L52orW
BdTXCYYuDs1fMW5NGjkSJUZmtCOJjgDEytjGpaV+Pz5SKn0Fqfldb3JSO1OvBWKsVxbanLRWWdxa
miIpMyBpZljEub4hwEY5Lz17mW726BGKG1mvU7DbgdrS3DcyA67yb03eDZHlsmzUyJeellEfrOe5
sElTbnvO6HgWibueFGh++i6DmTc8r9Y0Oblb+yQnOw8RPOMrSjWBk39oKbRqh4U8dIrS9vH/uBdO
vsMIrqsjF9ZLMDOPwDfodjLOzF1II1w27vhlNCY7pTOuthbvdZ0F0I05y0GZ0Bga1vvIQL890DrD
+atFT9Yai11Wyd9GU90L5aw+4odSY1lGdEjua1jIxPdXEA5Hvktr6fgCSt1wAE60LYNIk+vFmi+C
jVj9wg44q2QbcT9TnqEJt+DIOs9b0MDa3E6pDrVHifSiG+O7AO2ODeE+VlMDpy9Cq5Zw8RpZ3bnD
BCILprNZfg0/JCaVr3YIndp7g88j0jzmcukfuCTFBlD0/PLjU45wX6JVyDKEryX1LFHWftkmSCRA
PPRmkvu9dHbJ319Oz7iorpdYUOxR4oEHh/qhGSPXk2cOkIeTjtUFGAY6cFlCTHB+y1jOCDdYNIqR
fvS9VbNCUXbnsa2Cl8WAMjBcBUl3/drxkk7nGVxz5wNXSCgpiUfeYAR7d5MQx0P8rB0ABrvIEFVk
C6Km8OpowFVY8n4wQ9Ab3OFCSPgNPTkgRD2Ff1fGJcEOmC6Eqg9TYY+agq4e64P6haairzA1Dl5/
IMeHjH9KnVHKioET9yCSlKCkif8i7uYzyYFeBOxv7X9LmSxouGCruCU3UrNbE9vmn853KfggbUPG
OQrVLV59wnZBXWwuaBZdlwtT36k9sECAJcZdo52HddWY6ej5CKu1ZEYuEnOrFfXBXF5JtsOMdF0y
V0c+diLHyqKDmZ8CX9KfT7hndvYiL7sLuY2jh2Ntz3Vw9Af9PpvNXitchID33MOdxzhjXNh24lne
U4VPHSm34FhnGXAwNY7Fg4M5LFDwxI6ZvqeO0F3mXwf4fO34j+LHZeB+WkqRTH84XpZAcoWsE87l
ZKvytsjiW6noBxRiHQoaTSMwTpV2mF3JlfHSU/8D49K0rIbxfpIE4DoslqiuWcmhvCXCCmNGRB/g
C2HG43QI3xQLZZUm4Lm29dN8RkF8zst+9eKpyxSk4g/GGWHyuyZCVPjhcvmOov+d8GKAjXpjgM1H
ZBc9h2a8vAYHaluZiy2lCHujujy022o1KwYqE5yxH3vok+gddk1duNgBAqFOeru7g1Z90vVhHSph
qyV0MJbDtO7IzidlPpvUNNoK1icRwbmKBrk8LngiGtLCw/krvM7F7DXN9nrLShmjy+Re3XUmczZI
xquFjAOr5M8YnuwV/PdMz5ec7aUT8l/jpc2/ghWYf2P5Sf9zGgNk4e6PzERXaldXgPb8W6UB9U9w
MQUNupLFOO2vEd1jegIDYYPV+X7KJWnE8slLH3No6eh6qqqpjFMgkvfv15hYBFLujvikrXTKqE+V
/r2FW+1f9d5noNgzh/EE29IaVJsno34MAjCeqG6cWyc0J13ygovzNeNBkJl4qJBpBIzgX1nogMlA
v4rv5pg25Y2h0o1oEJq3HWgBhecVMSK0hM9MzN5gCDElz/5jKKcOtXjHgKZZQnD6VUe5Nt9zZAuX
ZukRkj31yAcppHbwMT0L48CCuOYnfF3GA4e///ifJ9vT4Q/d+E8rd+s1k8zChN6V4Y6q8BcJMOdm
6RTrys1y4kCBaL+AgLLiMWH3DezP7D4aCsfUq3u5XPrzejnNynk8CyJ9+yZvF7YyVep6iyN/GbZV
y2/KZxa0QCHc8gd/Df0t5KrWeh2xEz9xks5E+jqK/httXiCzIl4zD2KLub/mUpwfEzNsea6OwDdK
zR5ENBD9M5s2pUG1CVuixK9iYYdv2OvL4b1Oh2yqUpmdHMj4D2cSg9g65ZRyeOE6FC+UoOUxhXcb
/Dph3q1kuGRL0mWT069tgzd3Ru/LCbX5YYXvVOhJGW/9/OVKlQgWEkqRwo+AO38VjAJpdW0Vohd/
gUJoE3O0Hl9rbwXRWES+ArGKZ/faeY5Nv7+DIKUeXe7F5uv8zOOdHDPSuzgcep/YPjvR5q1uAlPo
1620upuQZ7IPT/RQr1q64M6oqbi1FcNINUXlv/VH/2Pk+T7K8RIb7QlqRzhNnTLXh+jdyV0CJN+9
C0phX7Uf0bUvPeBS22XUEetlgBwm1bmtt3CYE7Ylcs5NhkPoA/Ccd3qm7B2y3x5O9Ve+6UAdwER+
CrH8TKxQZ04mOzBG7BTMyMZJxomjmQlvHIQdPJOC82lh+4JrkHVgP8H23AAMhRzJpjyTydMKl3l5
ZL8CiXgTkB4oNnuhASOwdUWMafhdB5BBKIujRd9+Sd9H/ietLU6xQUcSfME5t9dz0Lp+cY1pUJIQ
LyTt1m3WTpChsHpLCKHrVOXVK8qR00JKUMrw5PkK71nxysIYht8sn1BHB3dImYOYbX7J57BbVJ4Q
265TuR7g7xssTUbLrcLg1Hv1YqazQopKK5O/SoWyE5a4QUAS2HsbSQAjjl7dCxBw5fBFtv6NcWwi
1m9cN0sKAHzLFdzy4AeR0IGkNnWeFbRxPVSRQJNRVZNB2JZxcNeLZhLK1vjAcMEH+5/Yscalxo17
WfTWbONjl+hn/4g+cCiyydf0iHEJOcXRoPrcUCVUJz1G70Xc2PUwc9AKRHzGdVd4m8+dmMAwbl7S
kI19MeveyxS+of6EHwrKo084cA42ramEteZ3KSQZKr2tTBdh1iKxrGxB5QRtMaGoo+hD0j2cIR0Q
i4/E9zlMPkGOumDjQn/VdAOUpkMMd2XoNWv278PYWbLvpxma7mNuL3SUM/z6wcy9Wj5ACAQ8VgFP
aHwWbYU23b8UjbFPbK+GuCXIxpsRDxgwSK3z3fPXNYWQVX11s9hAJ0fS10N4x+3LHw61T+RXCGd/
amGdVCZ25rnTgLuqtXESVk2Ss8FoTZdJ2XPmOpvSSdd+0MeE7667tb0aPXx/kXQqA+bV2m7QtGMg
YT1BPEGXsm1pY8TtgZl/UWl5kLkS2v5CR9weHfMYBUWY99QPgAweOgYZ2uCyvkMAJq24TFy6HDhZ
FbeGUPV7i33Swvz3n1lRFgrXEw6bF+TPdXOZGZNIfyRoAHFTcmFtWsaZG/9EXhc5veaW3lXRx+5W
+dJbK8qxkLiuIMReTcwk5LpJ6ck2lqnsJYmJX77wCY13rLh9LyD4S/MrauCwuC02I5Kq9EhupgKd
H1IkGbUBs2YuojCb19O23HxzeQVfmXDO55j8KbwYriZ+4MRZEUhNbNmIgcuDhnZFs5juSmX4cJZs
Mn/Due2SliWNuzrAlTefw+mgLJjjVykHgIS7e7aNQwa60vWShwwCjy4mKrkiAuXHVP2nUNIbWV4B
1T40RSNdkykWymViX46bbvGML5hL8IXVkZuozr8hEsne5qGW7687prpncQHNRP01uQdwobTiIDxf
5MUZsfU4JC7gMST5EJ3xro3JrGVTKZhnouxPMb1/ugBZy4zCDUAjbMAQwoTN2hJfpxoXcc++3iU0
WI424ih2LPN1qca3XXwrxhWu5BiYf/4mkLrkg13vegErOEiJ3mEzjcjXlWa1ZyCdkABvHqL2HZlB
xWAHXT4X6QpoXgta9l432R+BxgeqY9arEdVjZmasKwqQ6/h0we7sY5Ju9BllYNS7GmpxSo61lfXk
I+8Kjab2shqBP51M53K83G1kHwLPTZUnaOrhqf9WEiGur5HZermt0tL93XPf8MeQscDzkfMgssXB
Yo9TbaBNCZt2ihl88lmfrF5XVGfKqu9RCjRZ3wvT4/fV3bavaYEUV6AmBhHE19CHFCUQQ84CGuhl
l5Nx4uPw3O/eOVhvoAc8zZNe0YCP+tMx8brs8gsENeVRbHDVr2oz///N3dfEZOqXkGrC/lTLqOF0
8W4Wn5nJPzlYyqWE8lx1cCuq8dZWHYn/NEWt+ahsivoe9V+KAT3e4vcm1KmMOP5d6fJpQJbaAkdb
6Ib0bsCmqzRCJa/WQ+9+lDS9JtyO2OW/vivuNDhSbaBPVpdLLdG/eEOQCOr8Slc/7K+hcFvWoGUO
JFilqdvnUJNpHuVfcKNQU5LhAcRnYRuWHwM9PbT6SGuPG5YQzrEc54tagBkP0Z6gTduw7c/2ajIZ
joIaQ0vPtInfOVIgQxhVqx9PZFByOiNiVpm2irA5AHJzwqIFdq9/ui14/PdxYCmrioCEa1YeRaGi
k7dsU6nhlyUwnc0tItYRGbshxfsH88TjaghM3cX7eMfFky2b68I8uT0HZZIy63xIqi999treDxp+
rhGXswJt9NgcfJvT/I3MC2bWzM2D9amO+2Ypxt+17yybsA7idrGdI3wzuXAGJB2Qr3aEE87UowLz
88jCuvxjmxZ6mGA24ZgMyfaZqtpyJTWUKCyacyl/BnZDaEFO94j8DmdbZIjHHzRBdJXnTlqYYf+g
nEpsPWWm1K3AVwBd3h7AlwAdME+PR52b2YJ+o5Fs5M7vrA8y2C6cC8V5raPKvhiHYLcbzzTYl1GV
euKwKLZJ8MquuwQLMZqm3h/GeEC1dupfTa8SibuznYIkBV4+J4PTnrXl60/djCKCsyxiS1+fj+zC
3fOc6CREBuEqq2AGff8cLlbMTYSGfExaIgr0ZsKyRct+QjSM7s5oHOXo88E7SLTsgdtyE6cPwKRY
ij1ZTZ8HE7Eh8F2F9wyag9HdncsdViMB1EBUZI7D5UWQ3420Z/sRJ9HHCkJ+z4XMI7VZxTh/exKK
R23qHl/kCryYhXU6AjjyqRC6MowGRyR7bM2OGVfkuAr2pXOhrOYeVDhJnI7yACh8pSDGwBxqp+6g
cFKPxz6ZSg/8udB9pOgTush1FHoN7zpPgAQSgecbf5Krpn9oWqQSal591BMahkEXQ/QlwZRfy7jI
7muypj8IgSVNtdE4dKdfKoZGXBZek4NzqnkXp6aqckePT+9XvW/sm4d2hcSB0nH7XLmIyJQpG0x6
DSB8Irp6M3C5XJ8hLxX6XNtuD4ACBi4dJT973VwI5QUvFqF1jViat0PJhvn6rPH8JxBnEcJtm1Qm
Xc2sZGW65IkRM3TkRPoQq1EsIpOJgb7+axd1ZlDboMq2/1Fzr9LQzbCIzar0Ed6hwWCQFPvgbyW7
3vHkEYY2UOY1x3BHB7daqZWEOWeTTh+2zaCCbtQyCBlEB5EMLzqB9SY5vguasyUQjzE6NnI/4+rf
o/4DIgQ2hiDu2yvW8r6cLOJka2qfjEVbuM/WdWlFIsGt1IddYttv0Nl2OpIM9NlWutGYVLKgZ6pR
YJ7tunmiJrchWK9ltL6hwL+/Q+SeE01wYff198KceOkTKYgmh7kuEJeVmaIfvXhBlPViauzOpofK
nvxlCjv3dhR75IXGn85lfXIjxR4LgH4fdKxvGC51U8jwSgNX39KnZCHKl/jaqLWL8e7D63UaXURA
KgAIbd1VvYLhWvwgPbpbWv6FEyNwXKi6UIyeI5j1LcxOZm6hyLgai8ZNgqLB+r/sA36QBbHOUH2D
VVqr3Uc8b2pQwMRwZWfXld1QC5/P1nxFaPeAElUj5e2HKw8wNhyFSGB1YyP1uRFMPpMuKU6tGhsu
MoPoyKlMxESJJDvmk3J0wfVmJUqg48s+ZP4nsBtm8D114zBzwAZMHF/NtIgCtvK72VNR5Nbs1JDP
NnqlM9hT1Ca9vYeePfNEHhPtM/KVF1ijFXjTMf7VJIRcrBXukidswcgdo3eJJ3+br4Vv4f/oZfls
J2yere+D19p7+aXbM8VGx9mkyZbdyjsrGPnddqe8jh4oFo9UJo3s2jM27yV3pNqY+mPiom9TEAzo
PkI5Qx1ZJCJthXvUSiTG/8ieHhgY2dI6/Vv4ZIqVDqz1q7NqrpeImg8eYfdos2Mr/pQNXDQ+f/uU
LRLAzIUQkki/vY3GHVYZ8xP8xOzijRhU7lowk7vGMPLdLR8t0NxiSe1xGsOfD2ok1+n5MjRNSVuM
Wj2c+0Xnc8ASPNtwtUrqUYSY9UlYzH7YFRz8EIuiLMzuSNhVbWGt68c1+9MFgqBUNajv2/jfAABL
hFB/nl68F1tkEAur930Fds9wLSxP8/tZ0Qhf8LRusaBJtzbhIPxct3c2Fnd/5w25hxT8JvPLt4z8
vTsuPHoPEgCoYQEoE0chmuj+eKYerVjdVJPnM71EmrLB8brKDHYsKe2grm0GwXIeqsXA/QzYHCEA
vhPfADuF9WNu08uaZU01MYM04SJZvUUAAUbhiIS8jxUIdItFebvB1b1KoxQrTCPNGEbZ+Qz/l3t6
qpHv/yZ0kF1U1nsUP2JaR5QYNIfky9ry3Xy62chxOxNyOYQviWIV7efIaV/5IWZ0Vq/wP0KfOnVf
NUjS/lGnogz51QchhFlARdkdlnxmDJVc+rkAbMy/FdnLMHK8AnLN5CCD/2Tsjxa4MLSMfC7hBLnp
HNdEck3Bo2k76sr98OaiE3wpO5rMSl8ml/SE94YPHtAlVNXZyyUK06e1Mx1FK4eYTn7qp4osKRJ8
eFZmt9hzj0cghbZQxGA+gcuP/moDoGRbPQ/Zfxrc+v0jepl+inZFne/gJx3ep6Oi5MCSEqx7uk5i
ACa4OmEbENOXwKnV4SdimUA/kbOr4yOfGLxN6Ou1kNUOMXzgbbks1DdBKDrw6t0YJE9toZ3oG6if
LGmANxadpGsSz1b4oAzmb90/XMijj6/TUfZ0+lQEwmkhHnVF+p76SiurFrXjwoxuC1dLGIilvHBh
E4LtwE2YGNJ2Rk9qLR45kb4PJeqvxtwGK+KMuOe0PpwXaRfPnzioUOGBKWKj0NCWdol3WpqdlQc0
O9m71zkBbuxyegKSpsfQdTiQpBeCX+kFEChihevvD0rOPkMFnh6fvur7bflTsry8nQIBJOyG5JIv
aEtumWgZIrW2mLr2ZTXiPHdP8+r8HhedLqT5T93tstgueZP0lhLoUIkKrU0tci0hXrZU1MLugqgp
PDHnjs30q1v1IUdGZ1Vp9bRwd3ax4bF9ftZNM1ec66nIlfiYGonoxI6Sg0uQvPeCbYg4odKyGvWZ
j6uiWfLOvHCNMR6UVqx8g+B77BFUTYPGPpG4KDquDHeYrvWA/nZsDG4NQUuq3ufYBXv66TPNv3du
xduDUl1eK0zs2uSErzWU4EwI6SsnbTwFqxMBD1sNmu9+PUNWu+8V6wnXpU6CAEZ1Av0xfsf8jZpj
6MGaHiYr6gcMlkezgMVd8o3JqTQ4esbObVWyd8t8bNrSgQNczYYFamjDBGtIAsW8jCNh3YcvF5A7
B5lWWc+snmgTXUdF1RimWkdE/JuE3NOoY1MAmhyQiM0bZ0GS0Uy49mFyNPN7kcjfAvdOMBghXLU4
9lGkeNxIk8gGEndVdHy+eLSLicJSZnhw/VnDed4euv4UxZZ0AaKfp8/gkhHY92c2xQ8T5koZkUbp
R0+2CwovKydbMlMgH0PyQX+qYc9heSZKyL7VZdVm8/a4IIjWuwTT14Tz9fUwO/mC5ujyEJXPyi+c
e9Hq5IgisxURs1/q7Zwf4y0UGQp5NfaZPKuzlM81If5qu+y+hAYJY2FJvwWqKOEaF8VU7aTqUM54
Y72e1t9/D0/JUveCyZGAvpdXDbJIpndofxeCFTBbfu9q7XVkq+UHL/DMq1VxZe/vWhZMlKTseHH2
o0zhfrjUfZ/i8zHcaQlchi7wWlffBRJiU3nwvdsuVDFFKdRBRAncIicWRRNsbA+4f7wfflqUmpMm
6LaWzJeupX8y2QWhTIthy5XOlmFRU+LZucNw13pFaQrw5g7ZMgwSkOCV/TPBx2BTFZXImY9JV7N+
8oi0qpJFxz3lIIK9jh3y3af17DVI7KUN6pHKvt+Dwfh5YtGLhWRgt85jGax4H/nLVTc/dnjDkGLU
/bJPKVryLYxzjw41OEcpl/bHszVZtg7Y+XoCwRTq2u/kjj40JBSIQbuQ9s+Nffj6HbNjCAawOg3F
ODnBDPqsjX3bOwO/TC56L8bz2xtCOr4J5zlbSriItCrBHOQ2XgceI9gltM4cas0/7025iPyemTTX
lcZlPM3zXZOJ87al9qAaBxMpFYpqlri7uP0Y9vb4NtkBPws6vvh2n71nqHvTm2OKQhX6wK7gw+QF
jay1XDXXakN+ElfvGWva+YfPNNPCoZUx+YJaHV+qT2snvaQdpZfnpL2gAAEZ73y+sT2eemmHhnHn
BB38SCOL0FytEruoZpNBcU/iBkHP/JS5tUaQc0210EeHDiOEqp9rQZmx51dgBeSAE7sulzuwP3k+
nDT92ixJMM8wj/RVGVcCTSVSM4ZifT7KtJGkuw8zZCaEubrxGe+9kt+i0LV4FLOOGpr9BMcydb3w
mhnXT2BCRhYE6DvTzrxhwKRv+ORrpcjvOxT1rkq+dBY0tjL+VaBGR7Fa2pxvBsO/ypIn1zVZOsyK
Zb+Mkt5oOHFN+rN2k54c7ntRszytY0pEZ66uNkiOLp3p7v/809q+jvatvvQYa/fxRXt/lJVQvSi0
kNcG9jTPhMWaUETdu1nVb9Zfa+SGLg6StyL6hqRX1Lesg/ezEJzr4o+sh1KFBBU0Ci5dm0+1UiL2
rMgMNa/1GCu0+mWlh9bbPDGmGvO1IhxlCAlW3r4l8ZiabwAxoyEioa53CWXlgmwmKddBcW0niEqB
67ka/PpYLmSj7Quh+T/xRSd3b2YT4P+O12ANoa9YEKI9CBQn6xV61bhnpuQffmB4RKHzp+nZx9WZ
S7EzIda8Y8dV3Zg1Ul5+gJiHWKBya7LZlIU/l7e8qfrI+fpyulUcblvj9Sj8BavjG/fQZ05eHBIU
cB7sN5pj8JDy1UjSQqa7JBRodTrlihCam9tlEGRolyTsllDZzAk4lUHLxSLDww8IVwPSwQTqZKLI
aO8FlLA6tFDMYgFNcrBT3gLcfDy3vgt8Qxid0URNdSy3EGs7ac4tC2C2XfUvtLHhVemCbW5DFfjC
lPYkLfaAaOm1wgpFDKEiZOWw//BKpdRc1sHrjYrvfh8Wb0KHuPTLKcHWyN061lC8uFx/g5B5HQvK
DVK8PXDduN3AjXzwbhG0lCqs5gYwPsD66KVya+e5q315+s/mwNa692B31U/egoqqLy2Ctnb2oLn7
5M6zVfOxl1UT1YOpOqm84Rl9cqNQLPcsTPbKpxoexVuYspX60unUADpqap8FXslUzxSJDbjKWn9o
LKbs9QrpjQVGnrHgkS/iEzQ+ZinJcecKxfbALpmyBtB5piNKjt8QSIbfMFnggr6K51C9+GSlqoY0
YVDRYesdxugZWATRm37M6JI/UpuSPmxOP+AP08T1QRvn9pxWM8a+0eK1AroV0qGNB2khlMiJom2B
Io/TRQW5Z/pQ2Yv8beHlPXUxTIXl0H96rG6oDk+IYSalc9tM3VCqDjYzWNdaPg9pbli7NzepL43C
Ghapb8bsh6XQm2khh1fqTqAb0oFUlBSTxDgF/ntwzqHnslgnhMVDZwis/27xM9yqe45FgsUE44pT
rs+4KssH7cxZxVjnrhBixFdplNmuZ5vQVrSVSOB2ZooJjVzGWet2KRuxwHSlYDH8H1C0fkmd4s5t
lEiR56SbN5XmTAXQrhhul6ewTp8Y91ascZKVG5/Rs7JLeaRcSpkZpSeEDlK4QX1E2/ltvTlvPs7B
VMugyMkPKZJiGIbWK5Z5G+qOkT7audH2n5NM6Ga7gHnRf9+iRdMfJazJsVmt3Rw+OP4kJtwDMpFN
HgCLLnxRXjnqa0d34kEYM8GS8r7f2jr42/nYZKFIPJ/Yocf+2+FHEYM+p4efELJM5+SKajGrMt9s
Ol5KyCHTob7/hwWSHuM0p2fC1/M/Wt4v1e4gv09hWMQTJGAvvT903tyxpLJwJBIvHbjuDvUWpvay
2vZKwgZFW6e+aoFTXd3hevpycEkMizuXqkQ6XqD/mm2afkpLOtDefcUoOgLXxs95eXbJsYNIMwWe
kxRWOH/UaalLuRBtnm4kL96pohwtyn4YlN7fPQOLNzckSv0NPOocJvdhFIPhQ3NVIeKhd6qjApw6
UnSV4WkkaoJ0/b0WJKQ52zLBiPreV8ZOHJXt5fn6RCml0wFtYXB4nY2MZjUAP29BVsPIWJBGgBHf
zeW84QpFixLpvPg+JMWg07FePyTkLr8UZocDLOautcMiCyQK+O3ZlF+teUWnZUl/l22tiC8GSXzv
AiaYjRO3RZvYrjDb+tjWAgoPkrbBtEzkhPyIgRbGICHzUSMx2mitR4FTFRhiIqB26KvLSUGAt3Ih
nJwl1H9Fu/8wr9VE/neiEAxKuGSoaUyj5bguTHi7kA6or+crzvEfzqmfEZrtkPvqsifT2WqtyJmu
9noD9NCRn/b0g3B7iTn2YCDaP7RXI8gcFyQ1bgGhSed0plf81M5LyZiKD4R5sur5OdQffYcKVrCN
5XewSU4Be1N6ABkw6akqEWHHzPUq4zPMKQTCqtqztackEfXvVDQDJrNA1WfRJwuAYprntOy7PCzP
HGuTVOQD9ZTl+QBoN9uKyWFpIVNfok/7ht3omhViC08uDODF/k6/+bSgsCPLGhGrdqvwYHq3+8wQ
i0n/meIgZNGo13mV943R5MyjxmyKe1cPjfXuzKNmGRtGQ0agFaWpEaepGbedNgkC48ZgFTTPvmQp
5MQWmrTaUjgV7OFIqs8//uSd4w1FuPQRk5yNZIQihJXqfZbfspXldKNByXUWYzGVeWtsVsG88kG7
yC6xHUo0igP9Pf+SQq0uv9dHErNBD2tIX0/YYHpn/LBv612iKnOPYGFnk9P/zxUhHMzWbh8Rse5w
TaAsmp6fXVnM0jg+gmDH3pxD2dVwVS2WZwxH8nUbLTBLPgRHeMy6ZKRGHM/hAD9pPYGCCUOq9JT3
aRPsnwkIi6Ck4ZhlhR1LgtsKEef4gtxYvI0FJQxchNConcBrZ2xKTllZEbmJyZ/II/GzomQ/vX3B
fQqMFHYgv8n93o4HE1GmDL8Hyy3rLAGgnjkS71rFIo8N4LYZn2H+l38ZjhsHvQfdYeNUDmA6Ysmu
qpBgDuZTWazBxVoMTW20hMMz7AFrtl8cRAx/Q3eW+dLDCRgql71KlgXCrQ6OE46h0no/czDuKBTd
GuCQnufXi0SijoO0pG+/oPmlLaDX1MI9ch+1/alic3XRZi5JOTOPRbq3+zF4yH5GHUG1VpSnxsjX
FRuKRshrwcYExF7VO/k8KkME7MovsdNiw9X5BRbCTMo62u8ndkte5iEvWUhYf0lMdeTPe6dFCy0J
xXHEDBDo4iaPCA76h92ICRhKym4V9kjzKHBt070dOaN8I1ssEG/8So862NxsndlC+ThbVQbbTFQO
tEcqrAh9uLzE72oN9o+tEj8ULJ9EYoNnGntWKaPVTvBFEN53a4qJFe7WTnsltRDguxui6YtSb4f+
OwkKGaBNfWZQLBnGW6AzvOr+yBD/ok5P7XqDPg4tZ5X0zsPVreOAaVAevRAMZVFC+Bz7FMyhuHGj
pW7Qk7mMMfHXiF4wbeDccf4IMystX28p4+AXNAbXP4Mp1WJ9iC9o40gavYrH9okSv43MxHzZQ5hc
IwOq7bMr9SDuaG1Efa3l8wSxAS0roGV5Jd9DZW/+nTJSn4GtDEtTJFhJD+HQtA+Jhz02lvheUwI7
85Nt2A61+KBUl4WSvAGRfjwzhL2qLKXZ0UGJWqG4Gu23OsrslZYo9KU5HnlQvkEhvd8C9Loj7+hM
KwWLT3/1akRSudRGT1KubVMkvDyEGIPBMFTBIztC5hPv3vhofjRkD01oozaqJ0zIMjFvnla98kYG
hxVfzTul2Sw/mO54a6XQUwHtSFi1GHV5iMt8PCo7ppVRo6Fcz531TQNj4NeaI5ssJzc+CNkk9TiM
1EXfS3/0i4t9S76nviqCH9Nl+7z3Qt7d9x1ZicOZMkR1CY/TU9HmN8dlEhYSSOulWqR/7hBRd7c3
4zYc+MGUdhMiaxvR1x5JXvbyZZCtLoAcvaC5mDysExb6DjGESTR62n+gy7vSvjbBFD5nMOt4GNBA
8LlLlBI9XcfeiaFoJeqk2+5Xv/bJFCySucACsQ/1RLARfcyRhZT3OaxtouNv0NpBtytJ1v0elJ+6
A7KvLDIvRtfdQlEW4tBN3QWLnl4Ymhiz2eISh6/4EftMDVLGeSQKW44LgoD9sdDZN1kfw3yySYDx
tZTr1+Pe3gNdCfoNERvR2/S3c1MNQA6KBX7pA6D9jty//sYG/pbX1JpeDEwwRTGeEiV7BudW/Spn
8ZKYKCTJqxHrHaj+CXHINDegvFK4WNYI2ZmezXMh2zzMvQDmZpc62IcoEjDPuNmhXlrIfYJ+RZuC
TFKV/gUgmnVFlUC8jdOF+kclfZ+7jx+Hi+V7OIkzCC1UbqpBeCfwqr6xzXNOnBtvk+qlvD+5dnOm
kahUx5HwLVDsg4fqEuKT/AxcVipH2LLA9ZTaEAJ2HxroArpmpW1QYH2ZlI1llDFfmLLkjc08LVD9
XhIYjb7UjafexHVptNb2R2+quzEaC15zjYLKZgFM2wsdu41zN/rw75EiOlU3qR+0EwNd7xiGZZ8p
SAEx3hNDkC+iDvL9WHIMxTda85DTl01z2s2rq081Yj2cpPr07USjhzc9Pzm2vxljcJPdUT4X+qJU
39DvH8SdD7okx/K0PPNeJZZSv0XgWGr9qN+/nJ0ew7GjR/qqKTonhlFA5mxGsFrOtj5d6RMwqk6l
tJXU2HDeILyuocKk07uUvfG4hkBmcsgaGwqMckXEBVBQ9c1uPrQxIBFJVNDeqXOv/G1ZhAHN+625
QxYRRPg9dhSvX7oqsHbUR9AczlhbJKhVpj6JFpGqUi+xE8r6ywkyyEr//ig8kDfCTL0E9Us9n2sE
BRAtcVkqZ3bro8ENlH/mP8VMBRELDdHENNk+pAUIOFzxKIZmxbVJSNTtl1lFwvg6xvWQF87sgfcD
Z/1b70tsMKw3Gd+2yGLgjCbYeWGNYwnPEdLjGY8xouWFXu7wXOL5TTlWnZZCUK7Xx81EjuIDSAMf
1NUrrjSJEHmkPVkmYAsJIU0VgihrY+24u/KtpcT2K+ARN7UkB2aFnUUC7rBio2kUz5PFtaKW3C7T
CS0lzbDzwCE3pbWMr6dwezJhHvljt7a/vB312mwGfFuQI0pDb0RQhD2g2Af6PBeCzi1L+z3Oosr+
S6elxTpRxsCACWXREaZp7numjsVOkKXpNhAQnd5kmvnM2Dz1Zp+xMvAwYpSCFgjtapW/zlzcQkcd
m/lJPWwhiyqU4/8MZRqmND59dgAKIAGbv/I1qM8ZmcF9rEr7XBCrJsB4s9RKu6DahxQrp5uy3Zi4
HbVbUR7bFJyTwJFB9nm2UHmyyIKu/W9sCs03FpyX0WKytPtCBP5vJlczEwTDInYE2qqZzKem3i9J
xWkR6Batdqc+0FPXRwMAvVzTFXfXze1Yi+VCLa7hmyUSosZxe/WQMJbx3w5KekdL8XkVtVo/bgNJ
G/EdtxNLC6mkgMIi79FvHOwIABq6Yg2KKCbbC2FJYHTlX/ylacniEXlsnQvcu8XDvc5+WY/gKmgV
io5HSd/SEp15i83UBby8DrlZ45QDmkoI2ipOnhUVEQ4LXnecPJALM41bBgiUU/eVoOwAtXYQjMvj
lzJXTt+TSDvYlQipE0xq8GjSNpiElazgIcmVv0INQtCtnPXBTbkZZF2QyabvFn29MA93pQbXsyF2
CDSxNPtozEJLHd8twb89C7U8nijxbYFmP37p083QvFOgHASY/tmW8t1KmeGDvjxJYIlv8TMCK3zY
rkrhHhf3nkQ1O5vAUN+sGZqWQo3M37QuzAb/fsXaQCehJG62DmpXZFkPV+SkBNAaui+M/N0g0qmB
auMrvHfh/9CM7bd/a2lKex2K+TVmUcElGlp8ppsrDO4GmQsrDRt4ZmnNx+AsrdbzBNtXelcLx0Hq
koFxA7WHcmenAOqzkHLm36gLlUMfRsjijaQk4ukX579DxfvDZ03ecWkJ7HdnVfaZ8svjN+0Z48+4
aAEGc+bMihA3ZxX5Lj4rCGzSMRVw7eDdWkRrIveL7R1QP6ZfROgzhvt79QGX2jpHAu8rg9k4AS8d
lv4I8Vu676NnqDNnDVfIxOAjHj/aEBcIMIJyau9Pk7ipD5q5Ldy0yvEBm3xvmfSfTkMYcyb/i4kt
brMHZSoRFFrLRmuWhP+WheMcBVYQ2dumDyRF/Tc0I2RVG0qKE6921fi4Wi6i6e1Gian0UWB3Lyk8
pGU8OB/iPz19qLMuZggBFD7UKLtwS8x3N/ci5lI2IhhmaSKW4CEbvgPhdzU8O2TjSt05xJn1qw46
VXU/bDSs1AWYy/wWU+h+lsJ59BRP952+2yb1KinfCNEpLexDaJLR9nBsS51biabVflezHFjynQOn
DCPkljel1C5KA8vYtMHYPhG3XKcVj3juNpaSWB94gXwslKX8yDgGXQOEJydYa52iMM3+3oairacC
50AXnOo6tpi/yBr8vl1Gy13o2webcuvuVmmmHXm8KLaFR5qpCah+SvgLtPBLmZZR4Nz8uK/rGx0e
whTiYJiw718mpa/HEdxA66A9QMR6MVm9ldQYxOfOuZAj6JuGWchFg23ioCZVRuQc24hhXtmloLpu
nD5dtv5ys2xXVwWg/EBOq/ZjFBHv0VBb+b/SatIN/0bJQf1cPEH8mwaXcPTxhrBMSLpYAnPabV3Q
+3Lrnx2VKB8Rnf47hRO5uD6LJjQNriaVA868mIiNaN9C7zMpHX73JSGM6AXuzVrdbN6vroRFWnY/
b8Ne76FTjgrTLNAIFpxdfUsh5N2/h6IcmEN/3mN6t/9ELOpIkJ5p5Pu3ss46dkFq1dH/mhFD5K9s
Ocq1IhKjELLeeSGaaKHnU+zsRf2PmjDNc6wr+cwucTsmd7mrGOrl7z2KzNwA5WCCuuW9vvlcXq6N
kPsBDm5KzL0Cddmze23XFhTX/PoYJfCrfy+OiWn29P6wBHM0fgfDMoieocuOVZ8pYkzmSdvpnbBB
kMRRlrNifI2fh2qkjqtcM9RC/KcTxZ8QKJKmMGgTtZkmYcw2789gkdCRArJz8PHeSDwWIYg1g0m8
PO3bZ8YfmJ1xOElBLUVQjErJ8X3Kn82GiBD+zLkxVptjJlHTnTLqqcGykyRkj/12z1BRVZn89tJ3
MTYhkIO8LQ7MNKv41E/JlI3p8OCHGOSq0CyrJA+K3FeyQt9MBrMoSYDQkHC37TJzh1YZyWQd41HF
wSFwnuxspPgRPDymQOcwCa1ItDqeNPOyFA9UO+3caUVAsKDB1gYBIteRe6lPdM4pgIFT5dgTKyLR
/97M+05eqQVeHrKudgZku3sF2CbEtLm8JBxh73LggobrEGootVGZStdWmrxuUjO5o1gMGf9Y6WXS
SYQCfybL2EOaoPw0UP6vB1hPIRC6XhXhfTrAKwPG6hPU9rdeFaIdlxO95dto9KLNewhzs23wANPr
+PcKK94b/NJP241nt1EwBVJt3GNnuZKLc+W9KPC1SLIH3ubNHKGv3NikD5GtCrt6lfGeNrNgpACY
C7nZd2UBxRDBfZNN6F0lmFGs39Src9lAtwxUm5Rhl1a0ahsgjyHLPhrKeXQikZ0CWOhH9qS30VKa
Wv2xJ5TtsEMWcs2aUSBt/AxBeYeL62ZX7o1Ioy3s/22qgB1Jcgqc+9yFCNKum8zOQwoe1ShbH+k+
AN0K329EG8YEkayKAMPioh1L15gLDn9hnzmScRpcKdo1ArKFmevKe3mYqNF+ltoSV6ADnO0VFAKq
vS8lwy8TEtjrd07LmuDJgFNOutE+7oV25hwX0pN/t0OLPAHfdN/DPD5qqBaf/V4DCH+EKV9tryUC
i7Xda+pgX0LG2WnZIM3v34beI2aLY+z45lj0hmKjd6a6qG1reZPs38BmyjQA1JA5ldBWMdq1w55H
3Smgx+EiyjuPPBWSx9bl/hYFU5QP6v7/bp52FfBP0vCsuwiZaTJiq/Ud+Zc0nKxYusNk36jsiHc3
zOUqCbinXSvBjCf+7esbre7iIMrFF8o40Lh9KyeeHqkS6ZxWN/R5AIANXvxELEVTgv+06Y7f22v6
jWrq1zAv5M7Vgznf7frQ7IdS5ejDsa2eGY9M3iiJwcTtGigk/cN3yY7RLtW2CMTmMdyrrLKjJu26
9L0XwsUe6J9Uu+U6NLfyMye+s2/B/hzQxi7IMglsXzQ4uGlq+muChyZQkMst9onXmlh0j6cDy9Bn
cgVPS584aGFJIS7G8XHv1XnJkRBFvCp2PmO84Qqc4BPFHpLJREvp25lktx6WPd9MNXESPoGKbE99
lshKrX/E+7QIzJ+qrxDxcMgx542W5vgiH/XBC/tWtYm4ZlAvyA/f4IXOAItALndU1GlfK19my9rA
sk1HtcbX/1gLiQ2lltKOsfr0dpt2MKHXdH+S3fsI4v7KfrjI3pFaq9v3x2boj2+M0BkKA2VforTf
98tTkHe2u6s7Ja9QiG1wRPSu1MApeSQoWmogeiVp/Hun4dC6LsAnHzSxmYcfPy+2CkIBwtyl1c7g
ooWHvDlYV8PwRjioOpvWEig+SHteGZxhHhTzUEvQMNyOLAaceGRjZ/K9EoDhRKKj0nkJtrNJTtMu
hQtDwhhVRJALQC6gnFujWDvAG8sY2acMqXVRnmh8LHI0BfgLooyXub+5Pil7dJ1G71xFcuagkx1u
KdDY9xPcFN7psXLhq21Upd7sKDVjDq2zi7p+bg1BeivQIqzCUYoYR43dMWgIQQlS+f2wBn3N649M
DSX4tl1DqUL/eddbhekDt/FuvmH9ZpPjPUhHzdQJrSJjOFAlkqsknfPx4V5aMxA58M5JNQNvol1n
d6KhPgsK9GTZoYyRmfo5GUH1B0vTD9dop05GIvdJoBeN2blb2pOx4OCtkTu112FmqxqIPartWurK
Qje94pqEz3PQZWu8sFqwKU9QoMob4fvNdvFYg7cv5mk43Klzwmsun9TXv7vaDyDHd/9Qsh5MGsR5
iLDT9Kb2oXMP7TvKsJzntZOO+2FJyxMubNiqL3JkTvK8kjOLnBdvdDxTbVRBEni80pVln12bx30E
s6+Lsm3mPMKY59Y0uMs27ype5CGugpr4Rs4yPyXcSLy6zBNCbvCaC2XC4JnCzawgE57Xom6H/APn
loSSkyCcjs8bu7b5BH+rbugIePn/mfmhtiWQns4s16P4kHo6ud+GDAg3BIWAMG3I0PVJxbuZJ/7b
AI6KlpIWbnJAkDrfp4Z7IcxTD9jtfY0U5K9Q8uJPolmXpT1chlOsdIZiPgB5klnwnigA0d8qjxVJ
J6ypOsADU7pRL/sOgIMA97FrxyWlja8TiXkhzK8mn6hQoDXwGj2eX2Oqzc67aUhwJypZfg4uBTLV
crrjBjNWj46a55mXKd9+zXyJohjJt5YHPCE7zXFAcgJZUggbyGiWGAd2qZ0B4me3WnUlK79pr2Sy
A/FPLxDWbW5/9Wd4UfxiSFRoaANeS3aMVlyKJrV0as2rDcNh0QSYR9R2SZYe9DhzBwgX8wC0wSBZ
BeNVdv8bhsgu8ZbvDFe50bTeSijqqOB57e59SBjsHjf7Q+PzgaMghuA+mnofvVK20OIiAqAA6iUD
KOny992Ccgyn9sTQ63n0sDQL4SFjcfxc132UZZg5DFSA65bloDmYrf1yTsEPGMA6seHxHrNY+gse
GSjjTFRsVt4D0CQAJ1KL3PWM8Cw0qn0YV0SKEfB15A6ulNpt50UhuXT5/A8EiCsgcJC5dPlHO+x6
7xI8zenOjtgK8+6e/rseQLje7RprbzNQeuyCUuAAe421T639UDG/QIA2zyCi9TyEXYh1weg+I2d4
+Yry0UC7BOa1PD2BlJszp9hrzbI0fIIufkM5cmpYM/eNJLFr4YxVWBGJF9JYOJUDLYO2uvMDgvf0
K4Fk6hDIsdS9v8kpcqQPm98j50LOZLG/Kv63Chy3JrXt3JXA5hwkLgoIPO0eCwNxCiMGCNEkM2Wb
prliyUADhCM97k5QeB9zrMlTG7hOsxbNDu2iUVpxyC0VWE9c/EkC277aXJtuBqa6edKjjiU6CGTi
WxE/q0eEngd6kp2VlZaER7NPWz+NBEsOken7ReVDSFvuwFVxZwPA52/XPbBf1n1Si3E7NFDMgmmG
158gIo1PgTU5CPcGJ4GaUss6Qw2HkyDRohTrTtP82y2ZJMdKnbkcuMBbItZAG1aBQvp/KHgue20o
vs4svwhm+tzOQKuXzEHU5Aqr3RmCWwZ55DJqnO9/WxNGQrwqzw6LSAi/uhJOT7yGIL4wDdoKaL9g
hax7L5o19ulVrF+bBdmxZDVdWO4HIGEU8VsFwyzvVuLnqTWX8aqAoMVIhxIAOIVeXDZDGwwsWsdm
JylLXSBZxhRkpwlSJdoulwADyF9qVHCXRRkNtC1TgOxrAzlnG2vCs5nDCvlM6uBUYFBTBjWPJ2z4
ptMmRn15feXgd7S+79qYk9JH4hifqbexSVH2aWD8kRNj7NTY7MrCyy6upPBHGtwUmsU+0S+ZtziJ
ZNRBuNNFLO1yD92sqj8SLbTuJB04D04gsBmjwdzYI8MizYIj0+03LWNH5eT0J+swfxMd+QFSxEba
RyNQ2JIswNXMPu3QSpQU/cSP1c3mxcK7yhVcjP2FRl3YAu3yMfbPWz+mFv+QPHXRYI7YMO8qsT/i
nHg/R0bmr8ODoFFTrU1eJM4+AmD5c4z/oZbi4DKMyp4pZ7M0CtuyneJkKqVNnEtkhHP+vnu1TPL0
h3M4kWd+3uMZPQJSAhkWZ2UGkbQmPbyWsvFXpeyD6C2cEc8zo5iI10mZq5LPWETD4kOTcyrDAeC2
jlRjfwjQga5xprIZbL9xyDOQskksSc4rnlso1mzBBGvC0o4ozCXvZQanmUUq4g7bQuZJFuYsyCC6
rXyqqfzeZVseG8s8s9HqXWd9qSTOib9hEnIN9J11it+/H/8s6zREA2Cg+EsWYJk9HTd7smdbuFX0
U97tuaOiRq6tVt4MTAGuWOK1vlVdeWwhBYa/AAsmCu52aZcWSEe68JmTOdhxLCW/R1+ccVFBQqal
o3pS0gS8417kE/jnzrlQ4N/m4dkSVGny3OP2eemacIw+KymvOey3yzOElVBj7RiGtT/XqMHfLbRt
plttiSEs53PgaVn04R+L/fqYdwqkZD8TJdHRX7Dyt9a39btNfTrQfNRkPoY9IIbYtXChV9ONftvh
oXoN7SwwnKbeB2+RD91CFGd0X02Rs3XIR7OD0aEhihlIKRSwdT6WG6mAUSZsOFyN7847yW38FmaP
E0ONVvQvJXCMOwG9X+NdP3jFsn0GPX7D6GdxOxyVmJ9RHA/lTJ+SV1GqnGDXMVCWaTFqhjJ4LPoU
nPhYocdBzEk19uo/piOItHl7avBOliTlCyVwZJoM1lD8Fyl+EI8SrVHVe7Ov4ZgmC2HLMKrf0fFk
twj8IAbudHOjpW4Y1N1o1qJVxpFly7lry0lnWCWJH8U2XNikvVbOnEQHZ1mlHWPztHSgcEo7EwHB
3T/ekXwjcmGlO2V+I9eL7cheyWBcN/JE/pFov1AhI+SFkm64/yhdkchwL1EPW/zkHbYg/mcDXdf0
zptVPawtHaHZFiORhp4Wl1t7sf9l5MbLpXYep7Wla3UAvmxSY0+CnuBNxaQpWrbnQEOLHY3aVImM
x2OVTNpM4+hYE7FcAOaEehl9UzmkfXbnMreMdPHQtdTWTjpP1kKE4oPOiDFvGub0ojXz0375DwH2
1w5Ze6D+wyK8aVwnRvHWIxrEwQHI9ppKrqox8PsH1hw3qrDBAfNW88//z1y2/WFDznoy2LEQYIsi
Jm2Mj6trMfWFw/8CSd8xCo+eS7I9K5spbEBLasUZcf9Cy6P8xLdHTBUfrlXn9dfFNaENFYWbhftH
XAO1gTPx/BOd264c2ZpM6leKhBKqGB5zEVp3j4Nz9nRFcH2Ow8cwg0SlG/Pjgq5ORfJujoqz46fF
o0fr8fwxJSkmJCF9dCmMid3KlXS/5+rQsSjGCxLaZynWjiQgM5mGDlpUj7F0SjJDznpXIzW2N5Td
gE3WILRRXcOkGL+QNm5k1CxPRTocscQLim3A7ep/UieVPcwAKfZdlI/DuksNXjIG38S4dlJZ8iWD
IoSvjPz6/X5GoBfRKzfQCH8lI6uBiWxtS7yE2ezOWK4//voAl6vgeAfMHPEWVpXmOuCZ2nPZqV/G
EkqlKuNyNGOYf/dpz9HxtEVqiYImz6cJ/QKFWuu57h1facvClbz73NBfkR2vnu/A/+9dqA4Yz4YC
ehy4Rwp+irRPq1tFwsLEIDcmb9G3Pdr/XqthP33SurJlTvUGayK6HLlzgXr6IWX8PwcK7yPeQPV8
L+YTx1snEpdxKG6WSRTqYNZOMfsC2JkOcmx7ntmEI02QUIpbdDUiDTpMVLZP+BHfkw0lDgh40l9O
ZOqljYQqJVKkmfWGrdWytmf+02aI1X6mP9gim/3aGZqQKTTJHSInmlcl3Q9SX2epp5Wb6yvmjjGH
iy89Tu9FkFrJcaJg0XeGi233aHDdvt3UkFtmZ5uoUPXZylLUgAibfiP9RCt7ewnxrwvr9q1cJ9lt
QqHfdRbdEkgwItu5POxuPjOaPlBeEMP/nFHk2OgAZgNYzLeSU2RjLApiqUIgZC8bSfsIUZKWNp7f
lWskEmptZgIorRZrZBQ32TPLwndiSkx2PGYHRdwGvNqdREe44Wf4v6M8/+s2rz6ApiXK5VBxx+XF
GnBD7cEKkKfFhpgyY4dXj86psJAhh2FG+mUG2YNvadhEcbrxQMlWCjLqlO/ZHPi+oX0nXJF9bSLE
JvqJ4Z+8Rw7VR8xX3k83jNxc7aWQujw0L076YspCwoAfZGMFW9doB64hp1EkJmA5kiiu5NoSNQ3y
L6kZMJ3A14dy6Hvr6YmdR+vsei5Y8YHO9K0T0rteas/bGIjl4/dP8D1Jjm6DZF48iVEly4KYzyTq
CL49uNAfODQLprC5d/jOH+JNrOlsvNAUN73cVbk3019E4HJumvaICgSWqDC/3G2hw/TBbgYTAasi
by25QaxgMC/9vYJaTJOwKNuqstYTLJhQg5j0KJGdW8ni1MV7er6EhhY2o0MyMWv1e/DvSsR4qip8
TT/2EfbQw5w7IbrpAgLcGgOCO0B5yjY3Y19eE8iddJDcQ8NO8+vdRZaTIXaeOa7ZrLFPM+d5SLBA
zz6kvduZXDaYBs58Bo9SQmEJ4go4zKADPiF+fqP6YERR/6/2sHlTwCjNG/RlZZFfE7gZEHKgOuS2
d26cCHud8DrtpFqXBDsjKXouHDj8rxBsFcfh44c7qCRx1Jnrf4d4If5ydttnxiWee1KraD5YsxSZ
h2yr5IJ2I0fbeKPpOM+Qq32sWm1/35Yw7ezilimRfOFqehCJdUDjCPLzdNpLs9CgdVYStnWa51SL
ueA6HY7jKh/yB9M6nsmhRNCaZVwco4vkLgWrvM0F1GwwtPnuJSj2oVfnWounNd1LauDl4KXtHTwX
da42oczbIPsT2LisIX78A+9kmxpJ/MNDlZwJI627GX+BIE/wLnCYVNMJOdFY5G+75wYz3fjOhgb5
l5EEvLIf8SI7/WDiH5zm0ToHCnKJcv3RtcjPfijn+cBIvNqffY6c8ZWrmaA2wQsRPhwDTjvC7Rj7
PGer4R3l6Cq1d8roj96bp4cqfCSQDaGmixkE4wY+WLcDi7O8AbMEWcnFrZeWgkfl8RivG3zC8Ook
pDPGlrLfe1LI8mWsL6TT6scIYk/naH6wyC6qDSzQV1wwNgAS6TXJhI5tUvUjgRTWw8FKJ3o/s4ZM
7aDXuklT0G5Fb4F+V+9fdZDZB0UN/mRv3V+GMKVoLhyCCybhhCTsqJ6jd1XeeLy+nI9raOOohQuU
22+4L1n6zywyrv6mh0hxPU/eDcn/PUe1BBi+Vashx8Upe+zQDXPQF0vAPPcPLKnVEn47mKILqilo
YIHen/j2jsmFoDvzQEwkfvmqrIX+gUWvGPPSn4l9LZkNhOEP7m/zh8DEXKcPhYoLzaFl8uV0uY7I
vONaPLSszEOQGtklznImzcnrROnFZE92GwDDsOskySEefEFR5O3vtdWGxm7o6Wfe454N7dV79DHz
GshVnycNpOpkZjK8D9JEqU3B9quJhgPbqLZVuHxx8LoK/nf5Zsja+05FjYesu5obhfsRmGgA7z9R
msdsL005DVyXpkqoj+TurgvAcWwCMMG9xs8FhxPV3E57Z+3Ci4wB1xaofjq0KeTkNhsMIh7Cyh+F
Es+lra6DkA6OCG82WAG063brU5b8P9KQRqHdiPWMcc3iWpWd6UKuFTWXoKjk62+nxVlo5zv0e9RP
sYt2ur1L8IuEv7EPA0yHz7pDSyn/6QSclz9JtsGWC5AP0tsth5+wPZE3mfZu0x4uKhPyQ62Dg2DY
ug0cldhnFpLpQb764EUDZn5s69urTdbnPX3+H/PF9etc7Gag8E+DYgGTWKMXM1gwncezYZcpG8I2
fctRPu09jE+bC340vgupl7doeO0pyH60NJR/icFKnn1Tk3x2TKNxvaRBAUtmVF+ESfseqO+yVTYQ
jFR0pjUW0QUBz3qVbpcv0L/xLT5YQxN1DPIqpZNI1bXjhqaK++UwL325QAG7mtfOVvT55HvKjLJk
4EhzQhIMtCIT4wDUzYRCFTbrB4BLh0IrM08lta1320YhhTZMEoJuU2co/oCSq47jcUu4dAJ5VxyD
PWNamOkheoedbnB86r/A1x6eeeZ2eaavDe+FjcAgY2+RStIU5Su9yobMK4BH6Xm8u9NvFQYP1eYx
Vm9lyxWo/2W7hm/0DsIwd+ZstlclJd/H0plPbtZixT4viJNkRDqktpsMmvs7coN7rMww//sw7waV
vzV5OOs0qrX8q6U10ee/amRylIRA3tvtcEZnhOrQyoievzaEweUFk4w5HexZ2mft6eqgrkuYd9re
8jfOAL+oIh8qjTEUI1v8gy36PmUw6801M1yyrMI0CwFSLJkXRAgjRne9744Wo5lVS7HDb2Ls6E0u
9CMRcydBRUvbNNTBKWqlBP0zJTB1wRI4XKD6q9+1yWVErNTaHh0E/EXo75JzO7SrarOmoZY+zCiB
IFoJt50gD8fOupNwGU3vxFpT3qQ5gCf3VzvymRX20QZhVutDM1daJirqZNf/XsjyiLfnoR68hSjv
u4RtmNknCRHJkR6t7d5NssqoxLfxEkw8YjZ3zCZHUCwLaYOyXdA3oPh5kIo5YLNH12bK2KeFgrXh
aqwSAPDlt8f5x5YR++TUJYocnWu2J08yhNSub7JK8JZM4DSTmVHDGUkk0cSzPBJUdBcMmG7mKZ9F
Te7/O9yOrfhl5C5uW1TdhH93+ZrkpnblGvavlYujj+xX/L0MFvjBEUhMT0Pl0Q01XXVF812vcwOF
6uijSa7C48qvmt2qulPo0xjsXAXug9WxSTVIELJdpZ2SZ5dHX02HnycIKKEf1Mc/gu3/BhjubZeV
qmp+RnChIlrInMDvLq3NjHQjVaZlAxEOz0i3fKzkYH3xCOkJtZMhixcQmEg+IpU8Hsl3I/DkU8kH
dY1BzKItZMS4JvNq3i6AkdFukNEAyerh5/JU8zRPrSn5UUvjV+ophLkudLH4ikBbp4JubXKHOh9f
iqHCO88a4Z50hKHfi63p/+XTgOqJW8epVXEtYCP9wFnzKxhAJG8Q3fBJHnQ4lAlwnJGHlyjBszao
1Vqe4zumkorzY7JEo1a0ZIR09GayBmpdWfik489We/fjMHx0GAxgiQ4dw92p4Uo46sg7wbCFpV3s
OrsgdirNHeo4gEATG02Uf0EZ5jF5v+Nqd0mO89cmkgj7C8OdlY5X/LsJy72vLah80m7mMp1XYRtZ
3TJCsoP8E80aB8HB4pyjLA1EcehRnHOkbsh7tzEorbUY0PMYDw8kKpSzD/ei7+0oxhCv4CF6yLzW
CcipFMYs53aRcFLdMDm/UniNbtLVOck3noi6hG4plVxZqyJlbpRr6EwSajQfOEj/Ue0sAIIlQXa7
UUsM89T+MLwSZvB/tCtcJSQXFNSmFo9fyTqKhK8ldr0QdYZS1LZ0Gd2Jf390xsFiPJ6cXrW6XkzE
RKadLo1ZKC1eIGhmwg1Lo+DP4b2WYRPyGaprkoGWgOnaK+usY7sNJXdomU1aPBnvpShSWEyefmU9
KkjcL2YEwo6kzz1XtxTkeb93UvNFkxQr3nmKVwt2zxB7HwDrnmpn/B4vHKbSBQU3Y9W4E1IHA4tv
EtMTj/6QktQHqepzi7PvvoazhoiYVzU9MW8prJRZjKwzWowt07IFio5ehiblt+e2j+4986VAKLDh
34i0aUnmIQreU3QaUdjysUdXgt0U6t1Ip2nMV08xaMomhTOh0oH9TJL5Y/S7aswMp2cdgroHHEiZ
xnc6yygz28F0bdYl70c8JJMckA+Z6Rx9iBBfLcdUq7ja1ghpcLCmKSgO3G8Stew0Fp114YdbsYT1
c2i90qjy9xChjFwTDXEWNASFk7xS9oJMD8XcQ6IQa0YsAjD1c6V1s0Az988OOBRml+BiK8OZ8LQp
sjq4qbcSV+++X0+qrhF6LywdP5U9BUrIFVAwuewY5f7m0ITXoU1LfO9H4JEh3NVubNXrWQvY+QYC
zEoPRSQ8DvXD3IGBM5eOQEWLBPxNABv8zxlxiIg9/e8+s6Ur2yhG2Nr6vpl/wozvqyTWfe3/I4iX
LUe8HGKc5+UQyoGRRc1WC7m7aP8Bl9D1CWWY/Ubh2wm7ovVn94zOgpQxqRPppZ6LmFYpLlTUmaBG
GiAl/s7LiH4WVSEWPb7SsJVaOCNmBBGdS8Q4riFXenhnpZK8CjsO7npM+2s1/x0HkUA7arMDXAZV
9gpVL6nNw8mDcl+gCwsfCkkL2PDoNMvBNsTFfZyv4zq9obt8ZGD7/hzsrbapodn2c0nTg6ckv85q
prR9CSjB67+/MHgrjZJ1op20feFI48RrIOKqo55cqnZ+Yn3eTrZozLlYpVEVZAeSh9+GWnBiB/4j
VJpGHNDIobY2RGZxC4yoiIBN0MVJ+SdgQaN9nDUMKgp/KexEY6J9gRXtyHPraSWgEOeOg2u0Z81W
fpBeeES1K9ssRS1BRsBcjnTrg874VgqO5KUIK55DkTIgdotU3QP6w/nT/ikfXUNwAgTq/+oei6l/
t7L02r3Te2kISHP8x8nkVcNzwvtFZX3bFFW7mrephK0FO6tXS+jnz23wMeisuBw0uKjkTxo5Ihvo
G787WPwzRLnv7v4eZYF0iW7uAU6TuRtyIv4Ea7NKsPtKkuO9MxJh6KCh83cfet2y3Ep2OLnrY+fT
lLtXbHrLiLjPDr+ZZNFe+yOM9/sQldODIsfjsO7awaie6cl2sPfM4yMYwd3XdAsw2Gx+742JggR6
oz9I9qkHeHJrSARbjGB3devPvh9deA+POfNGfI2MlV/YB8xcmuGiL8RXrbrU683O90D1whHetiVT
rkpCMNTP3ygIXXWlp1fcUFNtYlSsWGMtemSiFJYCkMB5MEWhKIX0lQH/k85DDTZd+Mb+jlOQpXZy
hvfz7u86gqIpHoirWZOOsXPvXWv82xn2sqxIpQQkI+cE7i3/nuNcIDprSRQyqLUXbxAAI9UCBEFQ
qZ0GnIpMWg3aMKNCwpTlfZvkK8dDLZ/vmKkJpx3Xsa5MryCkuF3T5TmFrc/5ZUgaUBbfGnr59Sv1
ZUuW1bDN3Dt/SI73tr8sCyS4l6Ab6N+rbwfVFgB8Rk68aLPE05NfplvLmzfgItF5f1fmhAmTVghJ
uxzolEMcw34J9j7HPIlXeWnnlpEgimwfZopw1wnDqpYtMhMbXOcD5TZE8TBLkVcbU+gOMXP2nAuv
2L9MMM+QyJpc4NhExiQCU0+aVylHMeqW+KNn8nRB6mJPEEMnM78rAOQb8zmf+hccmr/zAYczQAqa
D+CAbHduKTy7hqDLGq5UZl6NWefZGX/mpvnKO/AkZPaVMXcopsj0N9g22KAf/DL7Bcv86OWeQ4s1
7aV1AJXZCnTI/UFLACXz5Omb1yum1FG3qvXz4YVV1+btvsaDyCO1JtnfxZerlTd1ExKN4Z86Iyfx
clKSmuBfqDjHj70YmTQ1TRceJ2YYSL8yd3qsrQ+vvEiryk38rbNV/Eud7//7E0cp8LvuuTEJBEJ5
Ra/BgoDq7rZyz5kecI3o4RYA8ymHpVBqc/4jYIopr4C8Rzlasl0jQKdnQKh9rgQmPjer9OpWvT6S
h0WYJgrPVhKPXi3RDwM9VvK3/qRXH0TqtmPGCxJDBkZAEX+zAz/diBSapt3yKC2k+ZxTxUvujogX
9pQ+IAwOIq/zhbmYoyyEghECFS+XCk1/5MRzAU9zdnzA0KMf3JYIfxdKdPnMqiFeHFSC2u4CP+Aa
kxNGf+dpdEXFL9i4CtALQMqb1DLPaqTW+AWfnv3azyCnXv5MlqLCBeuR2Xw0pNXmy1/XOYE0HbIf
BvagkFo0/24mIYbEswO7eIFo8tiE1Wmazs6CwJIXCvek19PKvbi4TO+ewe/BztVMpkShSGh4X7tT
pf/0Za/4GH+LagDpA+pnzDgYtJYelSRhYnKCF3b+hCs+RnXX2AJgGJ/sIWZGNgzjz2SwxTN/CObA
H0dTFsI3hGyK3lFz7RVk+a8IkyPhJt+8siBzQYF0qIU9BnbU3732bXyWM4cJuBiSkNW/5fDEZLOk
Vn14RYyviAUNQKx1ITelrc0d8y8rATWfP08KYpu+cNca5iAVtg4yn01OlFhQa7qdn8USbtirWp9i
H59SMfYjE+aNC41B6HtHZxffMqLk3HgAGLfBmKBgoE9myIbS5ZaRQmUUQgl4njfJDdJmHTIr3oCr
WMxI8wVLg/LqP5WdKFJF3MgIMQbdp+A88XDAgNKQlWTLYPTu6pB3C1MV4i+GLSsInPjcG+ImN4Hr
uFIaO4JCASCbdsUZp9NUAJb9rSOZv/BIzPddgnB73kxkxT0I4Vqfh0X2ZvL//DpbxmHhx9KBdikG
lE2fdVvFGHP5B7q7KGmnkZuBkNURBXSBUsnmiiNQqjPWX1Wdy3V+EBNVWJaRi9ahatzGbzGhKelL
myMxPnk1mqweA9AiY6JNLPuYtaYiBJHW7JvG8W0tQkHnA0PvmPy06ZsAks6cRIY2hsNkxa5ufoYV
skgsQKRqfcR85kgxW7cuXFRE4ulgcaLHluGI61P8B9Q6RhkknSgfRWaOCTY8eLmTWwE6ULeADp5v
SnC1w7Siv3FGAU0V0KpUUiRQGWiF7PB0z0rOnY084yrfOyZDbpwORfXLdyi6pMRvmpLEdvnxZtd1
BErGf4iM4GxL8NASTZnPmVSsAolsprreM7HmRNjQ1dIJaR221iFI2lqbkdHUB5dip684Hoxeefbu
SaQQFuMVi9wXhlJEnOQqy7BeVRHPDS1XPMZsxBTRzfwp0qYbYqjaDgw2Jx07OR4ME0ySR/jRy5j2
iQ+cpxip5rClg66mXOTFa44N9KhaUkadM/SgSO9zUjKrDEl5S74o/MAZuOG2GkOk6coTi4neAzXx
ymmoDQ4nwvdVaxUXUmgpezPVsoVF7nWbnZ7jMmcSStm2tUQf5tU7ZfdNv/JUTZTEeSKkWorfIVXu
LqCBCj7VzwRx2QmHzlVK2LkSCacYrFr1l88Lkyc9v2M0i7npZ/Qlg3qq5s463Bwa8th99bu6jjd2
4PisyIyR6AS7ikVLP/96K9R5lH8cvyZc8WTrdmQUPAwyhLQmitj5lin6JHaKk0xk8bC8FZAKO2Mg
emHIVNW5/2nJogU3fAfwSmgO9IrPCpSEkC/yzr2fIGaknjs2wIw0JQkYMFZQgckuerBXIghxqahm
hn8Yl5vypsyn7hoCEdwTCv+UUdVXuc8dAK50nzyJGBF+Slv8NvgLUjqFPs843uo2LrM9CbQFAk0+
RISdrzADasihKp+3csgAxchHmvENVnFNPmLv7FI2lSebEVwg6NFIIPjVIkJUVYZesrH6dp/k559g
VmsR3H03I7OOpNldJXrPmUsjlw+XNU0z5INuijIQJ9mSj/3ThqO7dMNxqcBSxiMzc9gvta7P3sZo
evqIUxZKKYK+hRoUIgsE8thZZicoQr+VCQt0nqloT6qPESjS8gQYoRNBLq8hOvVDUnDMYPE7XiLl
dcAmke5fnreRW2w4nf6Od1ZwI2TZLzJtpnXUfz1BNweeYhq/mVdRj4Eo8lQ3l8XyS4gGcMm93+Uk
eoxHZ8lvHxwftqcLGzyH6Vn+Ga5bnrld/5p21s3majPheouI1IU7wllsxbrVywOWyGwT33yDbJxZ
E+PeIAAIiEnLPVvSihR5UiaQAU3nvuP4EsqT0fq2DqaIGh4IO6oprin+NeRHbJZTrDoTnwfHRgaJ
zzX8ufi+p61pLV1FBOemtZAJelWh6AhYaLDtyVEMg4GbL8ojNOtyGtKvBiKZZWGmrqbnO/RsUV8U
sShfyqy1IOvSiC7WMF9wGdPtKVkVA/2FRzu0QnWA9VD+nQyuJsU8NqYkBCI+H0Mb4omXw/Got1uK
1Wri0AH8fu4fy/vDCvmmdPAxEUz2Sr2GGkZsBZeZAHa7j2rxU1KmNRF/1NYK+nksZldLWkaDccPN
IjpZeYVh8tJ1XbuLUWmCz4ruRsDbYbotmqtJHyR8mHRQKdk0l3IF7E9ADNESLl5/6DYCs3OgN/ap
INJEeBAZQPrNbO2go1HGaSsT/H6BI6I2P3NvG4NNahyRFfotgwR1MAJq1H0py6hydENxnl/5Jjhr
f3s6r4StnFfvYCTd0OJ/kgwKyhrEInRwra79nc6zWiGnTIhOBU2W2deJLIkFcaZpQf5rt3S5cgLn
cGSSoWKjsPbn9MtbfmnFhofOaQbZvIcQ+O/4cW3KRNb6VQESYfdsCigkfxePxThecCCfq6WqOPZa
vV+m44TCpCVxbKjdbP8qlXsg/7aZ4CCRV3w1RccukajchsdRTzQcNiYAZLD5KcJRyM01F7unQB8w
zABowAaqiRb8w+ijBzd6vVJ7ThQQfWJoEI6u1TyZpAS6PTDiQro9RyLNJRKejVGhN5uJSaM3YlPu
I5TvjzXmuyQQCHMb/UospSkfUMQsaVbNE6tZdbJlS3HeBqK9vLRh1ZBaD4X7ov7qey48NH6SLL5V
QX9IOMG8RArJO4qjDCLFJPVEQjQcjGU10oPvTwtgphOpUgfxffVSar8mAHGeGL5DWeM1ph6vuFK2
aU20JUZirFiuFLahTzA34bq2MazIEooJ2E10w7Y8g2YGIA8fURxX7Body0HgTuHKF9lD8DHEUYSw
BnBarTDpJtQC6glxBGpTWuhpEs6Bmv7r5fgCo4OBN3WaTMC5wU+LBtiSLWI02NrjoGkxQeibonJl
VCvEfmORTXrXM+eUaDGESgb0OIc7V4YFdpEsGF987B0AHz9N7FCzEKdW7GV9zcoEf1ZqlDABQdOf
PO0FOll6GUmS3qb/ewfm6yEYmZvpoALslHPLSuXnBbwP7l2YshdAz8fELYg3FOuLSFdE6SA0XkOH
RANK65qOez35szFr2+mUi2xbnhwHFblZV6tFOC5GmgCeotbxM8J0nwWi0RdbwHRDngRqZia1sIFO
JSVywx15jxavA6LVnKMChpyoYPjKepCjfeS9b76h79lzWNC5wxx1MSbtToelL7vg8rY+mzZNjHH4
9tQngZ3teMXOCyQ8vA9frDJ6PQ/zDKsQrJvfdjKtFnxWCqolhCp3uDs6j+6FVN1Us96A86+XEiaa
GeEkhqnMNAlJbQUd8i/G44GBRMK0SNR55V6ZP+C8lnuzrQHGVWRy5tDLZ3+Op4In7cB6Pli2ItsW
nxf+gzH8ZK+moFCPq+JpsbsTJkk+/JpcdGiU1E+SrTw0FNeZCBmrVKNhRRO42HWXCy942j+3Pd7l
6V1/X3Jg51GMfNvB6ym7i1gMXVYcoWpMXzj8TTxndVrzZHEe4OkzoJXfwdDBpQ/gzxgiHC32n/T3
pplk4ZhYNyP5V2kcPMR9cTXJr8D4QSt69FL0lKMzJBry8Y2gsPNtwgK4khTyLcvywn0WxywR/qTx
r+HWSO2/B2iACH3DYt4UMT49s5TTxZg7K0Or3cFXVdNvMwkxAH+umf7Vg+I9RqR5lDoVAmkAuTiy
qJ+zyRiCIvvUyilPvnGFDbJSuGkY9GRTgKnP8SZTDvyOyTjdjPq5EghjmiQRfRC32lGIGcBuEZTc
iIdvsz7cbtN0clYcBonsjW6Ti6iw6EuwEtwEt3EzmzwLW0Lr6z2dmEz3cZcaaz4fCc537WLYD1Ed
ZdnPaSeZIbGLMOWtQehLqwYzQG9Fl/3nswhwRnBn7jMbExUXx+zlpe7AaoG62VqA6Zq8vIxg4C9r
sEsertOtuARgWBVWzDdFvpllxzoRCD1CLyoq/3ikLPSxLPDImk8w1jEEm72jju0Iq9thoghMFSgw
hMMo1G2sLEn5hQJIA8749k0QirtpS5rmKniRT5d1Ryl9uarsUIc80yQz2KqDZYC3oENBNL8FS8tZ
rX/ZsruVqOia+SDAl7LZ/VHG1Kq5/8oNietbpeQvMTeuFeIIZxdVPskX/Ha2ZxtjxK9tr9rCmF/k
8lYg2aT9Oje8yhjZt4oLzrwaNmxPZPV4GgRmqR3Lf8cXZok9ibkXTtizZRymjQTM7vyv5GaBbKKH
ZEc3emT7nodRU7E0tSMwSYwtlIYpOHzWFRvv16b1EpJmuVF11CggIEceCkAiuz4hMyEZlsGKGjFo
tg0Awy1+roR3dkuxvY9mtJepD1sY3okrB9JKsEFlo9gqI3o8X5THPb5NFyKNZWf0GYE0RsrivVc8
CuR4giBv+Ga8JU22+r1/02mA9wbs88Z8ZwVaenX0C9SPJOve9ZEcV5ZRJLczb+0UGKaC8vHz2gmK
FgPPWSxIj8P8Tj1TZWC3jY2FOEp9zWwuMxdy1OMbzJOSTxCPjWZOu+Tkq4B8jPFyLQzld6O5Z4ud
MQ4Vqca+gMefGJZFdVAIkKDvhp9BoXHJTFuzavgikszM2776KkwLFO7DyKKkbSwpRobSUJWtMBIk
SvntLa8g6ubgPSTCQtxnowJCMTKvFjpRRdxMkVGIuIlJLdmkxjVwnIrFhQfa5Di+PAGGeuDlAkYC
ddEXExmH+8ONYFcphDy7ysauJGZmjmUYomQeHD0pK6bwCI4bPj1JKIGJQmEVv9BM4CJTzbXeqJb9
UQpnUfTv+L6ibHhu72CWh52ut9QvJDaotu2y8+3VrYIIaUq4C4YJJ6k2jGC5hb8HJqZbEKMlzTD/
Arn80nbskV8d3cJaXCAVaUflpX3UkYunTmnuyip3anobr/MDy72f3K6qhzMWeeVXYVoLSz91eGD0
fda0ecnpphjunb8fylJwQwQw/UqFaVMhPuOmXAPv/SWlMG/TDN6ggjYD+i+K3t6qpfstHsQqGV5P
/QEy8ITexBITxcJ7oXE0Of2w0oqMEuuM9QkMVk3dudoArXb7/+Pd/5khg4Gb5NCQ0NGX5aY7cY24
Brs1umQhm5xNAXojUC4b9IW1RwMyx/euarVyMfIki1pKGIwpxjK5DE9XrC47v37vxsaW/2ewb/r8
8qhWGQ2tIVM7lqH8r+rTOHJTJrrs446oEWd0mmM+Ol/0kSt44qIIASm7q3W7y98zSyHMquZ5Ng1m
d/2cPAGCGZdlclWaPAEGfJmp5JZyOXNWKG8eHMjhKgi3KTZ+/NLd5K+UvNt0+/5ITdjHc93OGZAu
aiDrFt3J4tsGUrLeFi08GjuguXNpUxE6mmAGZBAlnUsO+j8Mv1YF07vT0eVa+9RNr/trr1W4M1aQ
urelRhixkl5+UdNlu4LD0y3W5v/g3yrcG41LXQn+rA5nhxPrxffevsqhFGf4NdHRK95eFDcFFKM3
VX72tGtGgiTABIFgGA8YHV7r3Rd7V2orhDU9UsXMzIH59iXLK4u7I54Djwxhba6QKJMSdz5Yj5C9
TrPyWtNXMRD9+xIrhxFsItLXKivDSHyMuAm3ue2wa4iu/jqkdqCQBaNR5ojGPbrJ/Zt6BvaGOh/E
ORnZBAkIfSYjCVbbL/XiWplQOQhNK3VZzAdDa2nMz11ve6VfBP+QC6FHwm5XazuANUa0NfrKPhTr
laqBinPO9rX+YI3ZgfLI+DQBtXEBsQJNRa0G56Mee/AEPuTqDPhIKVeodz0ss+0EwiIP5zcI09kp
x///Wa9A72HVZy62CGYxcFNpYgxzrbumTL8Tvm+Gclj2q74ze5P1AeL4ieFM7TYe3uCZODKU7m0Z
gTTawsjxPYUwsAmnnRABVZHofj9eHVEz2vaKbxDtva3+3VrQukLQRDdn/ZQKAObuHoCIWLZwPcfd
QLXLAujfKrKqXOjaBMIHdvDUZcXZskTN3AVGs06ioVr/9AJQSYbbh2xotz4WP7s2bytraRTfSfCt
K+DElG6K3ztMykCMuMzzRLQXW8l5eUdCe0q+KVkvgQR+45aO30fXLKrzkaMtkn4A15NVgmInVDOq
0dAg+0s3Jx2HbsAywnPfovR8Puh9KHpLJKv1I44+8DHF4rL36MpSeRmBAMSBbcleCQkoLhR3KnBO
7XSl6NpL3cFwqxwqrxqIlEQrIJs789ou6qA3cdPLM46bXeHEGKSblqjKJ/haDejUX6bk/LplM7dA
CWAaZKHRonBKxXWmyWcgNhnDnywIbFYtl/TM9n3e/6Pg4bQqkxjXIJ6Py6Z+VfnRvk+YtTaGwK9l
xEx207Rtndj9HW6WB4AyC8bgzbusd4Lz8brz1/Q0R12o0Tc5FuL9Td2jTPQWx2+rNiVPUsrRLshK
CWSKDzjbZsr6i+4ankpZ+BcEYVtKwwPeZwTtz3ulnYaV2WVhvdtEZCBWriL/2Luc87wLqic+RUn1
AavSCbYJ1CR0wW9+UMqX1vvyn+ZWtjIGWwPNESpKsahzymPLyj/Q9FuvIVTQ2uglrCXnMZnIB1Nx
m6Xni8OCgFavfYAV/R3S+s453Vn4/K6QwrZVLiKbmsv6BM5sYmSW41zEZJz+Q8SL/kbaOB+0EuPN
5NyjskjXIlUXOSFUylVBVJkrrkE15HiOo13k8eWtqEHzPXNu/haVPyWa95Q123pSU6gsnfzAfGaM
thfOiNzNC3f1TOtJJILmEfYIcQv8c9HcQrF/bhoi/87ByiJFEI8E6ka+oqYMihoZm0aQYkf0m3eH
igCxurURQ7VsCvdRbO/AO/QQhoC8mL3c8G77Bu0Nyn/1RcUZ6EhN0dWNifhEG+Fmb/IphjkAsZGD
HXR4Eu+vdFc3Gs7gVnG/d/+QWCfPhmGwYdOZBvc1lu1EhQUKYrZwxBmNlFHWedd6gdkgZcsbdowT
vdyc0gPPdJA1iBDWR0pdF5Ej1IrYGuQw7NYYyVqtNUzuNtKAejmiDbr4lkrE4E/JBuZV2Cozi/j2
rQtbHp6Gi+JSD3rc4pXvdE6TDYS40KLGPD8oK3LANgDgMVDslj/3rXcInCgBnkP37sqeEtZ4SX5K
GxBYyTn//aM8dGwl2MQJHp2wVS9I3ZmivizdvsUF6aj4VDF8apsicglaANb2OS5C633zmP+L2Zg6
zBsGRWJRTD7GvKzum4EGMTrPtd9K+q7CPzmMWzBf08J9GMGHWge2FF3GuyxBILnUWEOC7u77gLlJ
OzvqAcjdTqcUxO1Esiz55LDVulVCZGUTrwAzWOxqK+6bem9ntWBpu8+xzTrsOjv5GfWSP18luzox
68N4TMZ1CzDw0XDe068E/o6QIrBOL7h0BhYAGX275P8JLw5/CF1d1kjCj6NmLzyS62hvsb1u6ovm
avNtigGM1oWAuXrGG2lkc4mWLarf2/+A8deJNdi74QL4MRvADqWV6GKD90jFswPs0KvPoxE3WdGn
lKeH8i5Lf+9E9Spmj0bufqcThU/ViL3NpsOLDiMqV10fX2ZYV4q/ZVWMmOsN63hXJ9g3FILw+thH
E06rEQ7ca3gbgzX2tddInI+EKI/NXBykCBIkZNMaykG528PlkZ0bJLw082ipc0XMaYZBiKvXrAuY
0Gb0RBe0bcwfoGYLl+OMrtPNmKV7AGgfZUJYw2fWc0mhuoefAX2W+V/W7t9UdHM4i9Z5kh6FzzmJ
eNMnD03CYgoaMgNLMjmvaa6sIIOco6UWMFPFd8RmljVxm4TCeXqaiHBqOHyUnxv0JUiTfCU11urk
jEeMvK8d4TwuPMVoeFHqUVk7ixBHRuQUOZ4ArFvMmQKnY63hId+hVjO3aes3UUzhFzfkrTZYaabM
U6UxxPfjmwqQjcaFJ+vrRi2zKkmaUxm2f0RoJrZbDqSTcKS1Ip2VB1GU/14RvdaxvR5c49wsUyJA
ZBI7GuuF4o1V3p2+INLrZ/fgDmLdjvZTA3wLzhrIubLt4rPqpxIPly2VWuHmgdi00/4mD1N2/jMz
GaD79J4WS9An57umbhysKihvS75bcaaXHDr6JJSDj1Wu6SGN1GuE7n56bDOmdBvYxM2elrJST91W
gPN5wAU9sC2fsWVEW67XJ59rL4l1d9uarUbjjbrRfUhXdxLCWXeAhtA0sTzG4uxKJg6LpvnyTXiy
j7CvDQu5FkWYfXno8n/rgW6mvXG/E59pzSBklGE0SuvALn0SfYzOysuBHhLijvx6j8ElPGFvpG0k
EQgZWdKaL3gn19xEF549tbN9rg/gISrAzd0QteM6jrbof4KkD03rzl9Kdd5pi+5G5SAY89SuVKqL
2uvu1oRmIAjL3N63G1pYlRny33QatPsi4kaABxyPnam0i2uKwDaInHKug6uxUeX53k59avhQChhE
STScrcTtZ4Uea4Wsw6P/IwmpUo6qQue9auLQcrHzEu4O+/s/ljChGJY8x5ddlA++ltrIMVqbmG4W
Tbo9c8TfHZNbB8EfiDelXJ1pnz90BtkHYZnRqe3Z9nuEe5txc4sQ6UhyN9XqSekGqd2KD6oPeQa/
JtFNQXsGIWwQF1443EvfgXErDdshvn/DRJDLFcMCa05ZSZrhWGUHTO87FIZxNiPxq+FpZ4V4x1W/
o8Jw1LL5aGwhpvXn5KVBY4AbEfOl0ZEk54yw9TMukakzMijKSZYPpRRl2xobwFELFlaAc1+2Lfyf
tBA8dxHsIUVZvMqq7Gu2fsvQI4VhojqDUURI8bd1ErfaV5ZXbgSQh7jAzhQbjjiAotpCGlNylkGD
O6euO5dF/WADoo99uUCFhjcPAp0IgaHlzeOWED1uBoei0BG+5z3rOR4GIlhsT6okKXTDKY0igPN0
pBXKqycMyF8rKoHECe62lX2KzudfeNGerTm/h+tHkw6YtvTuuIan/EmNpjYAbJQDPvPMM/8lfVt+
7yKWulq6xou7d08myid9MiRV2AAcuIgycCjXUVBQ3TQcrq23Ey73j9e6+fgwsg5q0wfOjToQPDKm
is8MDn2UKgibRNMUkBEYIH7HgMMfd6CTyLrypnaYJ4IGQUA9z5FKTSYnMMtUmAo4PMe2wafg5Gsj
MfbP+cEfvXyWcqpGioqJP70jgUhd/Yemz+sq8sPsvxynodQpQtiM0HHCu7AdQP0RrpmLaxKsgJLB
+yXFha+VuFJt2XjpjvFEu9AP9yD6VfJfurpHTjSttHMJFqk48xCXdqAzGS31dMvlUzxz/jxYe2Zp
26qIxsK9ffRj/2ggklVzyowi3GznfYUMyb7gixn4LLxJLgc6MnN4AWiuuZXQh9K6wYbqcqzlVOYg
kk50yn/mvFU8FsheYOWr4bvGVxm40WPmzQ5A4qiwtzO+8lqJ2pypEkhUo6P6jqtxNPTjRN+EOV+d
qFiEC4uDMH4YY5B6YJIgBWlyHi5y1POwuWTlaNkefX+qN2VF98URU45P5mCIE4d9jp6zzKsCpWku
uD2xJWDSwGh8o+301lEginng1lLlNeQsTe9/HoUiZiFupiqsYtztzp9iGM/4W3K4q/pbvzcM+3DG
3gJQvGEwXcwmCb03JaaZ3pDfX5mckSpYNNxFvONm2zRNHQDC6RsItTuMWYDs9oOj+IcymF/+qH7K
vdUIkfFPi4qFHA2fAGpAVdibgVUAAzPKriGlNSJlmJ7/uCiIb2zLlT8i3Vei4Q7XlgqX6cMYcV1L
EMJtWgwA0CpogvagyjuC9QQJYt6KDbaogcqEw3q4PXUVxlZajAV4KxgeyD4XYuXAp8XiNuI2ppO6
1/g8dkL84sW5hUnIcz0ikn5zEGgG2R8X+37vDxsQRVx0mv3elS/hHwvbQ5pKgjDqb6BX+EC8dhP9
EuCPva7Mnak25ySzIhrvQwYcgFteg7T0xNr6yRZzVN06nCz7rsQ09Gx08krLH5gv5yYbx3RKwxn2
EiHijxKTtUMoMAi1LWsV9Kmr2EPQZmb3JSiv7FS0vGqAA9S+yF1kIjW+4F8XZUxodceOvJbO5u/v
8fAGIQzbCJcF4EVyBzhUKiFj93K1f+PDmd2nFq56ahknOiei6HagojAUSPcc8kothKIhGjmYwHYe
Pu5nqtaF4l2nFOHtiiQUVwERnldX4niusMSlXvgCsFVmrBO44cRkNi1AFu4E6ze0QZmESS2J66uC
4PHzs6xrEHCKnMNz4NTkhsxD+PogEM7yIBaDNe48oxEdRHUcEDwWyV0ScMvRGoVR2lbDTG+xJeXE
r9dxvLEk3tJTMU6qjIKU6MyE2BPHBp1PoZSwlRBEVXBXy70/GyiteoxeI7C9A9beNlq9iGTDpSif
efJ0xeLQGCS1wzpWSGGpJocrOBb5qhxq1dp4faCJRnnYhXWdkwJywxfwHJPmO/iS5PZEDXVSMI2t
wB1RNBoZYs/lhVMEuXw5LjHqILCkN337VnaRgcG7Q43y2FtEA1Bw3DM85JS/B5hF7S7aCthsJxIG
HBO71D+g4k7WzPckNKhLEUqq327Bfy4y8dPO148ElEYz+xmd5k4X6WxGJ1QJOJ8iqAiTX2IJ13IV
0FIFQdqllK9dZLbQJEbeRFxxqXq+Iwo9j6pxjj7zVEQAJQ5WSxyrsFFP0xtTaLf1cJDeKcgR3B5J
w+fdL1eF+/xMjPRf+0FSev6+7G4WEnQcm0PXTjN4hewPJIp4v8zIHHblzAds1TGJ+KndcYPOKJVQ
TAx+YyEZAPVlhy/9a28HLmsEHyBbJ2spLMz1kpsnjzuelyhIyaVs8dJIiCupjAZbLXnslED+NqnJ
dXVED+DfvgsudAf8DpgVIpbgE+aRN87U+h7I31s2Q0G6VHE0LRw88RPyc5NT9qyPmAtrsLN7ZpaN
wiFUlLbu7VTO6v9EJR9rEvtX8f0WFESdK0BuFosY3E3IW9z3ZTUS0AMFz3P0cXGWtepV1mQhnnY1
XkHOM9ukn6txwSuimZkZprQerhmiJnZV9cxo31KjIBKogie/4wpJuKgFJTOzfjYs8c2pHXntZfsq
xeSVBh1HQmKAPuL0d2k5Ffw9Q9SE7C6kAdBqlNg9ngsvXYkvma+QWNnAgXitgqXDp2x+og9if3zX
aUZebgsqlLucb71GVVppeIAZssLC8b/E5dymDGgXbms1sagLOkuckvv5dTqzJZslzCnhAi5XumLK
/pc3hPO0As346tqiY2xid0Sw2CRjXo998pgcM/7u39ZOj0lDMnwNmrxQfaCaAfVszJnKyd+56FDx
TdkD6oTnj79oXiYa07AL7nKlrRFqNMVjCuKDtH/VuJkWmlaKU0bUitv5ysVp9OE91py/J5fAmFK0
NSIUvcaLlCMdEFV0HidyepgWAbjDrjjqphrxPa2syESnGpF7gNDbcL9zpWWubxZ4TZgh48K0KatK
MUMGe6oPkQZTA1eFlofi4o3SihvpuqAYp616f2loL6KzFYXzQnzyNHkgGzs/TUd7O+iYWZtvuiMr
EnStXiaLk+e7dt9VSbvm1MfSvbqfWvMMNO3ik4qPWg0w8yyNn1dP7nn3A9WEG6CNTuITNOEmba8C
2j/VRGyW7tO+pyzigYwh78w6BfGpEX+mVx8HWKmZw3Eil8CmRDrK/HagRBRTAIQui4bkwbTGYzod
I/tTx/BfozyJ5DOSUNzOA7iMz5HJ8VZ8Ily8e9mV2FfmCdmW5HOmHiTolkl2syVrTCQqQEfaUHd3
dZn9EU3MtdvQ8sMtNl5rT8jwpEXi1HNKU8Ii3fJDJomMovdMstb8NSZCXBmRdqN5LIcUnbkuWsyU
kOULJErAP/nSd6SZtryBv7fYz4XTOH5FN5FkbyJ4bjVqtQHTkCC21HkFkLrmg3wp9jvE/wRy99wv
RFjqnruygEEm1MC7ZggUSUimrR9bqELtBrxWSBG6syb8kwjWwDY/7AOn02XnwhW51tKp3mrhDiEx
1bjP/ca86mRqe5F1n8E0H7+O0jCTPTwCRxsr9yL78gfy8g1TRuQhbMR9/VWTAc9q1oZoH3aCsfbX
hhYEyI6bPey6cb+Ch935a8YVJXAGQyVQ9o88sZkETcpC0W0Lq4TSc9AUIycvY1aeZ9tAWjSclbPs
21UDP1ZyNCu8lKfffBcEWRT7WTMcPf2vj4vFKYOoE1oBjfH3dX4Jeizp3oqn07jhHwdp/UAsNpYK
XpUS/kbm3G/D7TvukZCP3n5jY3XuKwN6HRJJTFZvgUNlfUMisd3IUT9j2sl5n8bG82GailGI36XK
xHOqv67zu+/P7eIfsE4+7Gf32BTGH6aJqp5cyYHzF8hSxgcIdLp93JaXvGtgGhs0Kv5ekSzu9GPQ
hj9KovyuScuQ9yt0azaa/vyaSRTiJ27Rv9rV3YCwn9vKz5qtB6oG4IyegeOzLRoh+CZZs6GSlf69
WHPcLT8Af3DTcywTYGHMn9RBoqzEO0MhidHT7IZM46WSYzQez0El4eILX4gBsg9lCillMGvof6a6
TZ4uB7wzOPvSX8lIF+0B+0xbapQvOkVA1aEAkeJu6BJBahf1Gmctf6bOD186HbyeAVjt+LlMa8Ou
XemTQjtpZtyf76wuAM/+wxHSc79YwQzwyL6Oersi9TKrS94vol/lan5lV0HlTEscC4FHUh9jDW3c
m7WwBZyX8MLFo0p59bhf+6Tuov93Wp0y8lcdU7bjyJ7Xcw4YqtwvTCMx7m/BQ63EJ+/HBrPH0X5Z
+eH3RJHVx5DDzhjSOQcLY/lLom2pXzcQbx1bTdBzXoI6+/V6DPo+xdjO4sb2Zj2j6U+1AxzunnBP
DyzlzKDnJwPTewCdFESbaSd5mkkVhbjXYx8o81YrMp75WFMsW+gKpW9azqW5ywvacqMnKuuf1eOv
KKClNvwABGl9Dgsumea4Z1JfLEAFt4mO+2RxLMF989L28pxQzMRZPe3q2mAeTr4qdeVHnmN3ePTF
Nc3qdhAqVepzy0QmA/wi0vMopsmyznuKl7lXne493F2Xnl2NasiA3B2fyg3OPwxbF2qU/+5mnSsm
aQzFnf9Aaa06T24Oz67Lb/ctM4yRB1RdEN0eILWZMXnB1s8g5r9jShyWQK7rCNFD8RgKBg9L5k2J
0jsqtwtLWT9EwCP4tkKLL4GygDgQaewvmg4vR7qNyaf7tea3KSggNtZZPOEu4AMLQ9UabgFLHPmq
1EQwFN31RdXW4YAM52Q5A/odWVoBuokb1vaidCjNQmfuwsQeXktgqX4k/rpq+bE2igdxXNwBPVig
MMuDltSJgM/9Dm8ENdWKgc4KrVUbF+OjrfvncXUC+eAVC66YQ/19DdFIKegHjjHnaOVpVxu8dIFK
btSOhKwERfO82TCnv0oC1qHXvC/9sBIB7vIpYvXC9ax62kZ3BKtlypVn62uQfprfQyw7jxRnYFQP
vb++OADuDvZyyiSTFlC7mJwMyAcjkaWJu262j6oLvF70s0Ep78axerXYHtQnnEPcCMXDwfREz11a
LZ74b7ehQEGEkuqYq2D4KQ3RgpAyrLNZY4tfpnfkpdm806JDmElLpR9bZJVYwsjCq9qHlLMQ2ywr
wuhZacEOx+cgwOmrjJJ90TuPIzboGVCLTcgEGP3/DzZK9rTMVO7mpf+oy7A8rDGapTwp2y8/lvI3
0mrxPsz38+GGKmXuDlO5qj96SR7gdD27l72OBsOul9tIT1R62+eMOd21RuwiQreq751DE84joG/K
mYedEy1DfuxYwxs8zUaPUtLKdz6xh6C/S8IrSOJ2eTrPDmdRIigzQo4CTXhXahZOSfSQxVWDOX8E
+zxD1UQn9iZHHI4vjlXanjTDq5L92n5poqPlp0lUEPqdXut7WzUxOpzJlEYFf5KIF2uM98m72HhH
JxUv3p3T3qpOcrqPnZIL8DxUwJsAqrsEzyk1rTjxTAtzbe0Uj8bwgwJDBnWxHZ/LIb6/457aSKjC
L0VFyrWciKoOXEaPGfO5X2WcmLcQkj7PhWnrf911Rs3gMJjNuFZGTGyIF5CjNUeaJG/SwIft2Rv0
Sq8MR7VE+6Q5oa0RsWoUpRy7j4BBhcTNJGZZPfCa+uLzB5xOEEXRpJYosZVCyn4RioFhT3pTCT88
JkkqPeioFpe4FtbCr4gHapV9hLjdFZPY2rb0oXY2FuRYdDCM/NOgB7lRog3PH3UmOXQnBjBC1a3P
0T9IeXTK5shXzDlyFC/idhIor0ZHfg5c5n484gU4ffssaWLNnWiDms658vTZ+IjhkRodIj6q+cPZ
G5uhXokQPYhLwT2K91RXp1jBp+Av2sEqRcvaSQNKsrfGpM95FAjOY5xmt0L1cQ0KPKy6qdRnYMwP
knpYur8ceKlxBmZKNZcHTMWig3NKU1oLNfvpPyi9jY7ELc6ZcUsS7FAbuhceJpF6sfD5iXfH4r2E
BIAaXCG9ySn2sTp9cT1Ha6o6qI3rkF1JoK44Zv2qwOM5eHqd/lZ5tmMwmR40zfPioEcLm5/BX83L
Dz+iiQgFM/Ser6K0OWY4vreE0kDxxATmxGrggDK3s6DZnV+7x6bjkNcjAEc5i+wd7T52S51gSxOs
u55JnoMVKHBjXcrwvY+rGro5nshR4QRDD2q4fYQ7vN7P7hX98FHlMuGGkVebFDzl5OlGII1DLCY4
Fh3NTDlVYoLLs873DjFc9TtTGgaUlRMI+AGLhzY1ai5Bdyg+VI2WiqKcKZJtZGOylYawBJdYG8s3
3DVpdUtvZhKVgVpsf1jeEUm/nhtFO9xSA0wZD01colMQ7BgGoUve6bZQcuoiiK/C2dnbE0KLfp4J
5mRtl1ZfJXLwO51jIHT3Qo9utaVQwqoTMVyVs0aYSKSe4NMx35LrTY2S6jk5+HBS6YoUSVhgZHVv
5QUdCHBPFY+ZOTkt0UPIx5mZmy5COIxVehHGaKoAk5nlmRqfYCxw47JgrsUEdYcrUwZI48B/dlIB
pW417gIueaFDdQI48F6+5xTxG4GWfAbVgZSCwnargSIeNTtqvTfAPNNlkDaecS4W90RFl54kbRaf
9w8OvmPBiGet7fd70hGofkQw5n2BTkSzhBF1/ijdGf2Xu2G63ophgddFcxkcR1I4x8T8qzY5RCF6
Xjh2Fn4t4ghoGARk43QSQaqI9nFpdTs8VL3Tw3ujKqk629hsH+Rizq8Xj1yNZUkISWcaSHU/8tA/
NY3hyG42v1Xprz9sa9tmu1VpKAL3bCQsS7i/n9zqu9FgM9w812rIDsDvT1jLdqwTApglAyZdiKbN
E/c8fynCh0Hsvb7o9/8EWIfCWV0eO0jLl390DUoPVejLSJrLQD3RKzzW7H4orM1pEsmsYzSU6Bdg
vgF0pLBeoEMg8y21kIVepUIt2EKstlrsJk4tbwSYcmu32FdiSQmQpuedYNjqePZpnJwH5QSTmflL
p+iY0A55lSqK3B3Y3CshKOEuvM8x6hj+HEw9h7yPZ3rOuZR/au8QoRC7Eav3kBcxSxY6xbyexQ0M
+458FJJFXrOcZ7en1BM1OUPrkxQxOELErez7vI0+tdwD+bMQAx7aSwDVS6d2nQn7Sn4JnRIPel8+
s6dZdyXHXtYxWJXIWe1A9V0RG0KBGo9xrOQADPlukG+vhvUy0CfcYQG+A1HlDZzjBtYcINnDAM+S
Wnzqlnryjq22JgajwN6LwizMsROYV9iuXwp+dNLcWiJSnjIvKSB38uBDi6j0QBXaOn6GVzAyyAmz
bDaQCfF+En0aTCoaU+ocOB0R9/qADSqCAFi5CYfLICSJflEQ5gR6KCdmXLiKWF27hJ8M4I5HOTOC
vX0RKsRiOiWcZdJBD2q9WZ86Rs0V1uoa1GyKN2aKTBs7D2uP2FNbgi06c5Ly9dpDxz8LxWu5KzNK
8/k9CWOjmTfas54O+14I5GmqKZuLnNTHy/dCXOITk3HhPv04qi7KpJheHQW6aGXpWmpdCB/10IYN
JP4ivPv87/dhUxqz35CB1ZCndbMngK9TsC756Gml0nR6VBFNWzPpmYv6jekVjZQ8DLKT6sBlqcgV
Yjo2f3OBwUpyr/BXxEZPIUxplfUeEA7zPQe0zU2OjHtLy5NVeMUdrwHKRz0e24oaJCU/c5YIRuwy
SPvSaFSGY836GAwYgYso5eHAl2qyxpkWGFHdBwr94zSJtQTQSFFJwnJs74PUtEa2VtbfDxjq7py+
jm4iCe0ni5Tl+HtAMxmgmQvj38DRwLqklTVuUH7b/f14ZQ9GPkhLyTbqsa5Dx6bwLvR99dlPujWJ
obGSfJarBg3UbRf30E3Ap9Mrqs5YWgpwaAyu7aaMIbcswokJRrxJew/cSjhd2ugA6Q5MVMFMHeRG
+8Bh6NuXBZexpGoYPVnlGGWX/z6FPdwMQjSg/Y+k/v5vfGIVrdbWghXn0Y79Lg/hVyw4ftz1dp0R
BU0vgutsykdh96N8N0FRCDShCgVUkre3S6lpcjyUFs1A5PJoi+R7Pas4pxTbeXX3RtMBCLf+626f
1xbhcT9PXAmR7e6RiX/DgFvQkhnG6uwdVEt1WQrIMPXh4mbP6L9Wy9PNgyACzcXtMKY6JwwY8vsx
AmNkhxYVM/uukXtAqEm6UeYeVk9Di6KbctLvD8gPUogj0SRkfREGiSzeGNa9AC69B5UgHNSJ8Smk
/whjkMMGrhbGmkUdEHEYeny8JjHLLgPiziMbrhod5Fni37iGhaK01HpFTHOjlgethMJWXA/+MYeq
plrU+cRiS2mW0BJhEElR8OnB3rcrqPEViSEKKu5+Fg54+fKltrkK1dHeEv4s18sHKssqZBJ+EdQv
XQu9J3V4ouikyAhGuuQwFJbK73Wfe+WcWXkJQgc4SJnlAJrzb1tuv8x6+Xygz0IU2tn/+wl3lqXe
B4Hrkc8WrbnQl50oHOFI5i9gE/RpYezxVdUj/CgXIIyYm5BwM6BXiD08zPOFiENtxPNqzBV+8nGu
r8P5WYuyV0D1NRu7E8hmh96cfBipBZSD9l/fWoxQXGq3A79lU05dwwdVShi3tYfeWBWxd3WxM2Xt
Vl2S8qEIvRlDKeQZQsfvc0rohpWcvKCGjK+YOJbIyZl0EK851CtL+XMmxAf+rm+RmzWvQs59lEp/
N7mNrN2v6/5fzVoF9ItICzBmIQofmIl1FkWViSHKhOWd7+GewkPp1xT7i8+zehgaR1wFyKyxaCju
roCzYHWiefULhBjzH/08CpgnGpnXO8xRCHxQe/Htr8Wppm8cUxSAGprnYNhSWAC5CoZLnYbt8wZW
AxazUBnyDX3eC7XltlmD9Xjm5SX9Q0q2L4KoGNYsOGCcU/h8nKn9VUnBfCXbOa4C5rVfqdvbRuFv
/aexYSuwK3CRHJqfKQGX0GWQzZCM1bbHLuTGaLDRNjBLNh31V1vLB8uuUghQS57aMHLkmI4kCF27
aebSggI7mSbyE8Quu+S2d3YNp8e3KTKy9MVWtd0XRTYzX2afOFXKVk99MP94wGUhJG00sZWiFF2K
kE6fm2amlVzOdn5IyTayQYUm4f0T/v1VDTcFRAucYZt3SVgFsiE50119yzPZ/5dMBy8J+ighHvXz
/8/CnNiRcjYLC1uw+G4svuLKDKCUbwwKPgqESxVmZmekURfJqJGqa7mLqpUufuS4w7GJ1hFFwssL
bB4Zpfw8fBMyYMz2pKZ8W0rIipDLx28kIkvK5ALtusDX8rAHhgX2TQw3M2I4p6rk5FJvFUlHd7pz
MLpAYiXtyXP4nZWRi0JozL5xsfPpauz0iAuwbXL3TrNUOPT24YUjjnIsEIGDTNdlRBMo3z/V2zBk
N4PO8hGSXVGOgAVoJk8jS7N0CSnePhKQ75mY3CdNITZ7IZcx4XJyORMROtQF9v2ZVOXF7tk6Bo9O
kepf024LbduaHGfWqhIpx1N8ydoZk0tDVJxLHY4QQpIUwKlrM3DowH3CTPHkIW//fh6+u6ZoP9RZ
QybnB6u9wnLPNZLC0nN039WV0xHw+UtfS41RcqWjbyzwU9/lxqYBJz/ZYZC/TVxrTIxidf3cMcH0
rM02JIBoEf0EEDfiF0OTsWDDr8e8kQ0al5MVn1kx8kECYnYhj3VWgLJSAEFfLb1/E8nV5TlDi6rC
JEZevIPP3EMo1lmlw/LmQnAfXdr87mCfxT1DK9xWKWjUyVtoKbtoZOyiYoX3n0cz97ExGscY6rE6
KEWB0vovDgb88aOyb9FU9EkVOok8sULyBB0eMUQdLn2sOF8tEajZe7BjtuOV0euhvxjDWm66n4YH
uy/UK3FkwvIlfx5MJpCjjFIoxWuTq80HfhaNJQcZ2h6R8679r9JzwiGmgIcAcpqU3O86+YahHLgb
aJHRRKhh6c27q88HUzUdp+FYSo52vWJXW+okIzmthZ3SgaXfIacZM9x2PMS63FHrNYRanFiIqbcl
c9OU55TJPrY/Mh3Mj4WBp5IGsdShZ+LmYPqA6sM/675qbwaJ5lIIk641R2N9OzJvisnuyAIq2yuo
ZwkrtXOzfrCR7lA8Htwp9SRkyq7vd0IHQkqK+Ec4ddZqiDY5Jrppj/JR7wwGrvv9iNpreKy7xQFg
f2Tj6WFN/63aXK0sTFBIACqxejJU4B0WaL3aoy9cpR3t2UbQyH6dOIu59djXIQI8LCiSDaAvTASc
I3Pqu34gheA4ujdGws4YdilQRm5UKnjQ1K3d70DK6ODYOoFC+r18hab7re0BLeI16lJDogDjWyqt
LVRLS3x4YNibIs6AxPYq6aoL9nVfno81cKa3Zi5AoeYO+O00xiHabrqeAXpf/4MVrHrhXm0VQVsx
3Em7d/jvcu0/b94MCAHMOUdIsyFNjjXkMr3w/+Ub8P6IG2WhHx71cLpcUBJaxmkZpKJbAJE2Sf+e
jweVJNHUvncwe/ncYqHinYBEoTU6REQjFPKcr3vFzxnqvX4H/UAutn4PFXdMb/gUJWrpfij2DidC
Adje1UDS+4TZoyKGraPvK22/cqcUTBp3+HJli7DDEvrz4/aGMnYSPpVME0JaFQCXDTJJFC1FbCux
7O+Gzh59vIfJaa9vqe4d/5aQl5CwMoERIIR/eCtyR8YEq0mVbaeRYBRt6pv9kGGExC0fRfeW5W2A
oSdcTwRa9DcxLHwG+VbR4xLd21TBmvauRccRV6QG2uFD7zRJvCvDTzWK6b+HTY3GU3qOi3Nc6Iyl
qHueeanHBvPnhvavsIqROKSzNy72oM5kjfzwEYLriZYubSPzCP4mP3dwAo2nMsH+2vpxtIlNE588
JpZqkA5uLwVcRYR2xSyCWNk3MmnzWjw3wTYY7AFoKoh9jS1x5p76ty0p8S/OX4VWR+x+5HivZxBu
iSuYYpS4o2b51Wr+Bt3HeNZOZRdFCjSDoZHB7ccRdnIARRCj7o5OxT6foARTeEjhT9R2ylI/p0mS
YPVutUZYOQWOfLB7bhVDAXCYR0ogvsrk4ozBdxFrMaKGZa4eaUHxWF45TrZmo8UKE7uGM4WEVhWH
F4FS1eBCW9ajzmbUYaavDf+06O6dr+gDnOAad/ZKWs0t3PEcZFVIOr4WktlxNtHg2KTO77Rtibb0
XWOLKH5l8TpL8B4qkF+t82PnxREFnyID1NoGNLA2JnmsZOytEq0YvYgaQj/8MF4KTL7mbjQq+deP
jo73h82KPHIW/5DpIe8q7FF1m/Zi0Q8IrbDGvlb1jxjv/JetK05yBWzGctflpj93q1XvMyCsHHKG
VepzIei4iAzHqqtz2x6o2uRxbVQV1ip0QccAsvSCU1e1ygIa4DE9dWJhFmBckjZomizo+cN2LHb/
g0RMlOrCKF5xHk5SkYl6iSAwuP2wd6UoeAwNWFP+EFJZRcNrvSLauZCKwzmIeLy+yMkQ/vUP1oG0
VgKrzEFNPPLuVKFkCCyBgKsVlvQtWAWgnzMx/dFYIs2H0kW8yq6P4nw6EtzCtYZVlWTUl9FF9QPj
HbhMJB0+0vgkXhEIPZI1Ea4MWkhQ3zliLRnnJvPxH2XRmxQCCHWULJSsQeg+aAYpoqzepV9Fz1/W
WV2frd4fIERLjnv8mqzB0O7IbdAOEB2XCJr3F646CYSjKYGLKPgWZd9OV8ZpDgdRjULR5quUZplU
+GbmzmR+tRx/QEP5ATRs84Tt/Nbd6r1VE85z8KJ+hsWtnfr+iQ6T+BErsuEgWNDjUP7SNRGV9+3Z
ziAJCGRe9VVXDgSGd5bgMxDdeOAtSWBFcJEsnEv5MECF6ctfzimsY+Tmw5aHoWvOZt7PSeCLu7dP
4YJzM5R0LcXNepqR3UHTviz3+W0ZrGexVrpeLHLiJd2pacUJ7WiCcDdo6/G4kX+y6oMkYm+xUANe
St/uJpJmpIYR0Djv9TOnUkV/PgL+VS3emQHqS+2GEtTaKK8KDYB2VMN2ZPmhXiQqJ0s3ocX9aRSO
WB/X+dwstI2i7W9nEn6GrNE26Z0X+Pm1xPGqRR/Opu51qtOJC0S1COtagIvkxtxvzMU70ryW4BWd
f8b2qLbcL+cmTPbj58zeE5+nvZODFZP+jsPzAdOLeSZetGWwRLPJ+OUis6Gx5t49PorAtIzxsah3
VpLhEZsWZvJdZafsH+FjJKHgzaWd6X8biLf8qpdffYNs4+uO8bCtyKmR66vX1+VK6tsSU1CQ67Az
9rr+G9syW/bZLJ+r04X/sve0Tg8bXsfAYLQhrAanCQLfyuYNi7TKmzse3BsbMWVSt7/9ndunjoM3
5jRASl//vqdOh1lYxMemVFStAYZt0jVwwrFnYQXimicTceUI7QX5bkhgtXDF8xHPqz8gSlLhKHzr
qF39/28ab5LbSnzi/QGEJgDWq5/UUVgMRsyLYPSoKPUwJYYUdZq4erOx4YkRDzd7/V8UNU1T1YBV
LBcgsCe9BuXm+NXXyEJvwC1g8gM9V9VspGMlioeKxnnJqaBP/0yc4B+u28Hn/H0yXGBiPe6L3HYC
40M1h4qYWFbYwWwjTAt3GrWvEbmlhWDbdwqblgZq7F11yAeCuzDmwxInhvOdG9vdTdimFYol880s
fwm5dSTIsK3CiHjL7na2qjQPQT4RuBGda17o48FVI7/yOqh6zqC5ub+c90xr5DessCUMZ+H8+/lR
xGLOoYdD+U61pLMlRjuP4R4m+P1QrdyGA9YHfIpDF4veldmQ97MDs2mQ/m5clgU6/DUNeO/xOKBm
XCoLXu4e5v+8AnmD/T8sJcR5kbq7YVcwl2D3lqpiOIsf03bzY/ibEZd1MXPJ162sSHbJLzwP1rup
wJ/JZr3LpSwyBLIIPZZjbnfz3vdePQb67TkEiYXJLIX1ZBN99tYouDe+6DFu5bxWRb4wqX7f2WvO
Lh9FPQEuJLn5Enb4jrQQCg9QWjBuRSVnQy4o9q0qXP3FtuxrRqs/uGGFYjg/usjPCkIsOFGLUebq
eotecvzQecE1zI+FpwqaiAweo2NIIvSykf2/Dv/bAUNF7Ot5senP/E7MmQeFLJZULuW5JSkpXyiL
EuGIJf3s4qkGo0ytvwN8BkSGkF+vV5AF7CUMe8t+OH/zCL1oG1WDt2SVsbJQgzk21VbCsQZNEvn0
T9qb46c6mK1SjLSBaTAk9LHrNJ92PsCPyUlraNbi65mn0s3tBHgdTh6beb86Kjk7Y/HttIvLyWL0
0UhItoOnPms6KnCZFxhAvtu2f13U77h2ZvxiFwkUVPQURP9eyXb3ev7DkUSBe6WTTLgoJYUJfbhC
XOloZixeu/BE3H/EzIoCItZy9j2uN3NInrnjrI4e+eKqY02edPJfHhsO1OG0/1ET0/7ZoNwKckdI
zvdIgb4IeU3yLTixQ/JybWqTnTQTcvGFm0q8GEp4/LUc/hNtzdf1h+LZtw64yuq++x1KMG1nB+y2
rIFzkb6d0MdBI8VpHXet1kCM8ChMJboPNMSTszLlTcE8prSKyrlj83XhmOOlet+EDsWtyo+N/4+k
vUT1Oefujpwa7aIjuCmJBKwuWCIQz/loNRgjpxZlHrbzy4vVAjunf5z/uA8Oi1eySMwavTefL/JG
BeNTCAl0UaaX6jdQXdYOuiwqB2/c5j3ipiPdGyESbGP75fAKq7eYr6cpOeWmgQx9S9Qpa4SWrK59
rHI4j9faAigZeTajvElceSoDrQ9g3vllUKpvVCpzSVok9y99T3uJSK0DJuXx9aYgDVomHQpPjZMY
W2XAxE6E7JG+3+AVDAIfuCDgsj9iOS7pzfXm0r37Y0KZhvk6DavUa+Z2urPjZHO0iZMBShhdmohK
JCjCbKKVso3jJXsqX3708XFmMyJ7d4PfCxOwPOquvyKmK0mOot3PxmOB6DK0VLR+PUU86b/8GKj4
bQcio7YuezwIbeZQMDhxnTPqsUP3V+RSORVIEfVKoqW8oh2ugnAjZjfC7CZ1ncIvB/z0pjA9PYAJ
o5kkYSNzN/aUxOk8Ay+NvLgyVhsoL46OfpWEM08b+sYxzWUNDuH/qnof7atGLDjS9L53j4kUjwYX
sWKNxMFfTPEWtonZMYJ2/y9PxRkKpirinIVYVBYm4eW6PS5cIVj+UCwyXro5xbrNBGY74PYDi/JU
ylzn7UGSS33VIuQvPO9RdaMu3BCidpBf0Rg5HYRtdp1zpRHZ3nssOpvTs5oTY/CiBYT7bBmkFlvk
kuDrpAFzRp1iqWRbfmSgBhsnLHDE1tizX2Yj8B0/3EU1JfAkNEgFfcd9ToSkpakBym1tMG2p1NWq
5L9Z+yeSf7dw+MdSIees88nwkKvKBSNydHzdHGOYklnjtfalL3l0zWvWzajZ7pKT7yMebSCVElQV
PJcHzEgM1zpFQzqo/jX4jU4o9TvlJP9PfSCYoUOPJKg1cqVl0Lp/m+F29Ymilck+svH6SRR8PFbP
yFWk0OfCIgy9y94NTvPuc7afJwuTJo6BVfHlqxEyd91W2bYonzOyLZCGnygmBtmOKUCTYyDBwWjo
m2sKt6nxvVH26yuAubefq0WUQemltrCIau29XGV8HTiw85ySrFrWt+W6zc5Cki8L3Okv1MVx5Cpo
UmRFvASSeLbUhOGzNa0yqx+chLGZnnADJf/WAZygA0Ix3pCOisNu+jF3JWFl9f9sv8ks2AJGWEMa
QrjMLz7fLOPYyeZ8LS6Bjmk06Kytf4xjF2yxpP3mOb6IccoTpFWpPHOSpK4UotEtKgpvkJOHU+Nn
ITdR78MciABg4L/odqGK/H2hDmEF098RFBk6JQcHbKiXjL9Dk9jfpEXmIPaq1BbPPmW52nhUspW7
XyTH2WyJmn3p2kCwoa6ioFs62n4biE0K8gYWWMf0OihKhSTGIeD/bu6Uy06v9B6QRN8UWkwr4B6+
0c9vIwL1UpER98uwvhy82ISHrSg2J0rH6+Xyo2iAxb9uF46WHCkqFh8bRORZUD3KSCqNkHHGRwAQ
5AoXtVSv1PntIjcIbKqREABoBnuuisw5iWByq5sZHzuq3HTx2NaCXfPUrZ/ZkRdyOLy3AAgycesY
36/RBIcJaClXNu77LL0927tGQOsJUeb9maDc/KO9dH28yo+dYOHcbCZNfFZyJlAsq8sCCAe/RtIZ
+Lok6G3XRShc5rG+yAJ5+qCbhdpQVwTJKvkd+8JFTApHkGEPYP/6SXRJ+/nniAfq0MjTTZfD0IJN
l/d7hUifXs5tKF/9C8sEZUP0yqPMeyXlILTT/mzbJ+Z+Qh07ARjmkEFjV6M8EGZge+SaDPAs2iUC
qAbqi0k5No6MTD/c8MmfO587i6TIYBDYYBJK2j0+ynGKA8jdV2kyY8CUQggwuqTWAYYRnr8MCjoJ
MWA7lvlipdHhqqovblRXXib2pOd5cYYbtTdiNTmgUooutrQdAi4YnQLlb2UYWlhMiAPvJPRz6/nO
lRAecuyGgbbruKa28+LbGhBMcQoczdHs/KsbbTKvAqKFN/gPVsKT1lipDXehca7Wj1pYpj/nL2qk
vemEAiRDcuBeCxOZr3wHjv1gBQ9v76kDJ4nI/JEBOT3dokZQPWqkIV8WfZOyogUGPYcXnVXZRtAI
RWvncbs/acWPLzPRULcmh8pxfB1GSil3gCIB+02w0+XAoxJ0/uEK7RrAT+QmvXlNdQqBElMTuOjB
9LXeCQV2HaenSy1XBZwJ9HX75FbgsyIJVxARPl93mCcFEg+wto+oBygc5SPy3Ck0pBWmCIuIBbpg
74RRX2VFPy2ym0TSpLITlxgDIQU1X07tofm2yuxUzcEKtXZ8AMJzsZfpZp4v4723hrOvKwqS3L/7
dv/zbZowbMfA01P7EIE98Mp2r5jDkafi7mL4ws1u8FmR5kWs23rlEIbAWUtU4xY3+NTdRYltjmQz
sl7Hq9Yu8Odjr7GlUrpMRhbXIpAbF5Y7Abja/Z1y3ffxg1JgZGz7+ztoz3yeoRqORE3zdI42BqGD
a9RUt6s54J8pcufkcK0VqYmX75Dnbc4EdwdZKk/CuFBXjVg7QFonjrcRuYGSWCNB6dESMEQp1Rz+
u4b4Q0p4B/i8PKn79M2njf9bJMgw90RARXl7z1PaLsEQq+qlO22IwPvKTgvzO+MGcFrB0Bkr7pmM
9ZC+LFbh6R8kz3+ExyqUfOBXnxz0GA1OK8/CpvaXEZQy+vvJ/U1QPBysHmSl6rhyX8Xv9iTtH6GA
KB7Fl/1rMnXGz2aJ9sOZ3d2ENnmI1NBXRVyZqoC5FsoFc3fMt84K86sm1rAs9h962J6Kso8bJPrv
u/6ECiqp1rHuKIztRjBYusZwPRUGWq39n/e3qpTsaOljwyKJyzsjSnwE83tzF6X7jl27vIIVHEUl
UGcxoR8PJreWnWE/xRHs7txfexTqa8fi8pu5cVWCYCpVZ2TOMrpwDf12w1/alUvEhxdO9hmFGDth
bQhJSZpchOwDVjIFsaLXU0EkOGu6q12Ycsdvc5pkPOCCnlKCEae8mQSHNU02CCvCohCaz7OLV3oa
uG5S/J8R8cRyyVh5HrELLX9yBtau4aSREtM04thZF2QwkPBg2eLfjdIbSh2oKU6Ibi6JNYY0YJsP
S4F+VPAIkVaUFMS139YbQbdNbMFKMhBK3a0xuooGwfA/CVcA8BzyJuZfkfYIcc+fZNfxtPiLP4jm
f2Tvp//d+xQq3C+9E7eOsu6edpT3sdbiH2n/vH1mFdzOIjhFUCjO0UV1GCDR1Vz5ZQbgLsof/R7X
uF+j5sjLF+hhc8UPHG/Q1l/aixlW6Za/X3uVkJXe/23ZMGGGtvyCb3vMd1/WlN8Ogvt4pRdni6SH
L65NJ6gWjCCD2JH/sb4G2O+7UpnM2uNV6Q6xvVGwc++IYGied4PYDpF6lYuH4W7F9/8bPZ6yJxOs
rhixmGtwI8/WvFByDvLtD+FchyOVjHJeSnQ4UpLVdo0MFisid0Dg2c2kEo+DF75J1oPsr2Cb93fX
p+Zj5fN/PNiNDAPz6JZGCucPcz8EDGjgS50uNCGklkWwBC+CltucLMOe+axtmZtwAynS3RBTfama
BpxecTZpKezGip8YgLwT3fp29xeMZKhQwqommW5GhbcwYaWJTc72k+vCHQm8TureLqp5+LSUGtnL
XhwiRyruc2descw/X6JcGXuJ4M0uXyBKl6dQOBDsJx5LR6pEvRrxytYwwocSD8/CW9s6ag5I5w+4
v/Ot54D3Q27QJJHqTGlI2NVM9ei6vTIq3HlFPcIJlTgIz6maVOp1/uuhXyo5A14Rx6MMG41fdM/w
YL7QfQrepQcaE+HQSJGObpZALgSy8FsEXfgc7RJNIvDEcm/qYg6r46twuTbbUDYTVCtiqq+TjAGh
/Ba1tOUai1Uu36P5N0BQ1YBw/gmJv4sjby2Nk4Gs6wxFTS3ndli2DUOqNo4R8PYvrw1Z34tL6mAJ
zNHZmmOmalx+fJ3dlX9NoXBrgXguCPKuULwS5IrJCVoC8Xx6bAQ8Lu9w00e4voMMSdkAkr+cyOQm
ulsgfOr8KGfJTFhMvfzDKJGFSMBF3zEOcDsa0/QXebdsHtwqGOzGWh5wpzxJ20eUlOi2d46agmn8
ssfJK8EboWzdVLKxyWPA66DWMfCBzgXfz2VR7yFiXkjq/5p2n3ZTXOkDxDYRIqEMoh69UwaWql87
y7kGpTEm+QtlWulyoFODm6wQYDUBT7wXEm8QsOP1TT2YF/gAoiVYdtTXcKS1Zts+FkaXoRi66Llv
270EXNzDx+IE3tscrj38mbmuPFEfXg5TC9m2TNBAsXEK+wgUyLtIkKq8cHaDCKebirAOPIHiVRCr
5Kebi/qF4htBM35t2vCDXsiC3lTDU1TvnxPpx74uC5p/FF/Xg6e8EKPrksl4hmLgFdkJoSdWVfim
wBj1QFJuE7LpBB869TaBmEFtuHhHhy03V34Z10mJVNSN4qRczcWsZKwZdGZpNmxcDvkyt8sTqu8z
S0uBcNj0bytHX9d7IZXjpQKSmSxJKNtnCiJwWwda5P7drw5jsOTU/8AWPxwmfmXYhyCv69ymdVrs
EeEjyqkA7hf375a6aaiPLBAA8w1ejlJZLgviQBihNVTUrcRwFjY+JVi9qsplQJXfgGJi1foouLj6
vLAtx+SEkHajGCkvxDnDt8NNLv2Gtz9/EeO2Vv0NhjYdKTDkFmMB98Vyhp2AMQZykY3AZgumQ3vS
ZFRPKvrNmdDvPN8jdUcJAMe4gAVN8mhkYZgfs5J7i/8LWs4fahi93ytYI8f59xoGwzCUbw5TOSz9
WrprR+j4NK3eBTRse/5QTwm0G41llQClqUlkvTH3RnXrP/2fcwVZEhFxXtTK0ACM5yYW/o5MI293
dJC/tpEnoed8xc6c9OFdyh/CKY6BBzZgXaYKqhykoWrRd5kIyBeml/3XPQlE4FyZI3TVvhGHyyYw
US3lHD5UXe7KSz0nOgTSBiLJB9oZo5hMAknhcgSyem/KmSFNHLRkZAz+rv7FjoFZyi00QuYWKJPC
dN4WqSyN1AbSri/T/6oXyKa6ONFxYJnh3qmEYoliwcsQXcamOrq2KdpIMj1wh7HGacf8tdxpC3qh
3tQdj2EorjWnzv+In0Ol1NPOqbHCB39/DjWaAxC9fBfufNNyoOxLLDpd7quVvhAOMfBBotlbphHw
L7fn/lYv2RAqc2d577RYxvToshkMTSfFqcC7WP+d/1MHh9uCuDN3V/tGqyQ13Y25nIWPpBkTrzC7
30qhoPltg9XWePQzCT5cs1vS8SU1s04lytZgadiMgyeEcRx1OhplLbMDMaqKpmdPLU2eNjAyyuFs
pUjpqxZs14gF8D1mjPPD1wHUXLGB0P7E4PPeURFMxX62f9DQAXbKnLCUHG7CFC9mPJ7e/B+BrSQF
2SB837axgucazrk0k7x/KflcxJnXRHI1u6q5LUu0kJkAQJ8r2u/DUJHZq+McTmf95fJ57n5rPdIS
LVMaQmEtUr9f8HSG4giFBKKIoLZaNyXOFN8nSvB4GUpIwywz4AWNzq9dR5BkwIQJBbjIJukDBj0g
6gUxPrd3DHa03CS3ceZ9jyoznSEzjutIWZJKTHT0kls+zgR28+OX+CmRR+iDNGhC9OD60U7VaNlN
aPkCcexs0ob4TiEP4vmv0bKlnDgyuIWYIgC2E77+hc6m2LgSdWnFnZqL0eTTVboIr8OeLx1oEUVV
8OYPjZgKzf7anQRzikO70bNa4qBenK1umO7iO1lslG+pRhBJhvCCpNSTr8GRyFr9gKqKIFX8TYcb
u92MQbQMECRIYuUy2YAUvvWBiBk1hcSBUF8I5MOH6jJJIoCr2TEud5Up4A2HesUERqd/bXhRhNEy
PCnpWWeOnXtuGWVcgY7zeC+CeLAfERvZNFP0+3h+h1jTXvBnSANNJmFjaXXuKKQsTAmaxRnkBL35
HxQYwDP0kGtrYNk/aN8wDYJGdCSnYZPsxGiRzPhBiHzq6vWRsF7v4dRxIMrOpdNohWXyff94GKcd
q5zpbxZcVDjT0E4Q+xF7McI5x9716ZFSagBQ3FX4plOSVijqxBvtowWnrhiWaDcP5wXR8CpqCK+K
UqLR1estXLFsHByDWI3Wp9mYs1xgdLNpNHyjahkF+Es229RF/yoPZ81nq9GhL3dZCh72Kp6JMj6X
IKakJXqU8GnxAtQ5WM4Lpgek4P235AicMvRFhRZGTg4poMoC4f0mXAK5Nzdocjb6TbErgHRZClvL
FOYnw6bm4cFSefzA9JApy7+PVND/0iQJBxLcoksMrBb63Hdbks3sVuO5PFQeXsNSRKr1QY5Hn+c7
CeTH82OGYaFNSKdW0XUEm7VIi+uDzuzoohJF8YyjYQINsJ7zG8QWd7t3LHJweqrr0++r9MbGfclr
vF0bmfebr7nD2i8uWrnKTDhcqbGa1lMLFdCMrQJ6bDCae0JdkiSt8LIsZPPZf5QS2vallLb5neQv
eTN5fUXDKw/wxf8XxM9V6edmMbEs6PQ/PIFU7I3H42VALhlMXqgN4fpKg0qpOe/+/EM5dRecytnt
Fast5IkhhYUc1H7H8T66Iw65aeR3eUy4dG4LvbaedBJIgKgpVAz+VDiy6nS9vOcAGluKTKJXmvQ7
ctXYfZWAvin6OaDrRghVb4FUPSMkljHXsJDyz4RTrUNgPUiLBAq3sKr78NRFWvsyrzwYO7aaH+om
CsLh1ZM1KjOBBXOm/ILoC4xerd0cofPB9m12ZUX6yw4jevrOeDnVC6/sAl6EFBEi9wt5GKlyizI0
6yE2LUe4JvWlLKDBMVlA/AwWSWJLEGgGgD6SMsARMRyyPKBAyTMUG4uY0obJSeswdpnG4IaLuIWa
ZNBuqdLTUcxubJ/xS+aN/VGjaVmdVpfJsrazmtkdfW4gxC4zLBJIIr8cyrdZ/I30kbo/PojnUm0G
c9jpo9/grVmGFqVdt9t+MYm3SFlZzHHwlnfwVZWEo7qWvJqfw9tfs1cmOyj0YcshkF1IDIJAlzaW
u2x4cAUIrYQ/pdWb5kMxjR9NL+I1h1GXigbSjUmbOXMBomFyMH+URFBP9uGb1b4H6fTnESrbmXBw
5Ex2x9fnvAOchsTdRtTSGRjPp3M6hjTG1VKUIavoVOqzTzeXda9J95YyylPc93gy49nb3/FVesgJ
613mOmvbBP6XX2Cb1S6Hr4q4CMYzqrfNQncBUi1XmWDJU53Dm9d+s+CPLfdIZBBfx1xWZuiP4D8f
hXojqvsN9Si0m9e/GkE3lqjbjm8Wi3BZQ4MmjE1eVOTrRjzIWZ98trKHVX6x1izeLSp11MDyakpS
Oa2MwI7JYRP8mM4pCrImVTS/fMw5RPwG/LciMWDxzKmVC7dDCF+JdVDQDWvNLtvvfthVHCtAtaVq
POx+oecwRTBva8HMkHKQLXagJfkAXT0uhV9lMt7XFDUk2s8Gtz8VnaaD34Zv6RLZUTyIve8EKKCd
7QDHdtMwbeHGTGjBlLHDAsIZL0usil+rGo+ZWBkYknrlblcjckTu10FlIeOE69+G956Cngj2XB0u
nHj0erUCupaWDUzL++ZdWSJXAtvpin9ieK6WqLkdsIvBnuX3hGiYtAO4pFLs4LltUjHPhpkbN6d+
wlYjFlQqwVnqvlqChB00c81niIehv11S2ekF2fd4rCvowEacF899RS5cWHTnj54vdV9Nzwideah3
VkXON3f3n/2tk9FSugepww91D3aOf52m6dTz6G/qRT+fWw3qalCZJjw6/cIKTAujExZ6yKm+F62A
0f9RzzmT0i0X7nG9K08I4CyWft86oepwmNy1+VmCbEB7qZvLSM+CmwZUnNaB9OUIEOJtUNLjmTzN
F3EEAkMmL4BJngX/svmxD7Z+JnYmdpCzCRPsvfSexrWkeMbzXMz4eDblQY3hr9sH36cWnDLxzp0D
VrQz4rrxpN8If5T0dz8kAKBF5VyVBTyLBXNCRHqV6ZsDhM8leOwukrDNH5ES9Y9nJv9kqGrWzkqW
0qKb73rGjPyenukJIQRFodTB8ilc/A6xL4KzDhluDTGWF4i/Is+g7rj+w73g6pIl2GX/3qERXSgb
PY3DLyPFHO7uzuAMKPu2PYDPyT7wVOD4qgqy+YG2hfLczwaZShtcuk/MCUIqCyGOBIqJ9YzyMb7W
RRYJkDsicmHPuhPusQPt9tAnrA7bwFbpI4rvbolyayZNOHldzD1bOcq+qfsyYmmOOXBvkuFwYBWT
bvX4Cvi+otWmcdRmfFI1tqCHqm+gUyv9S/UMrpKdvi02b0us6GVRiN0lT0Dyae+jrppG52KlPmfe
gGv/R7E3uEHFm9KbmKPXkf6QQ65mCyO/AGyWfkN4TF56YChyU05/BdSGouhl33yk88Fx3A91l6R1
aKZ7XbfJkAa5z/E5g2D7SqZDnPXgk1zxJxJ2RQ0jzkkrmDeXSnsCNbWE2YHtsySfjgkHvVhKml3b
5V9TKJP7dxZKzTwN6K+2oRGCYOkOrWVCsPjaay3vEBxSyAUlgAEQRqKvOsHUMfL/JGAiX40MVr9V
Gfn3ZcxZVOSvr51f7cHLIUVuwxVlyopAVxU+/A4YgM/8ssDGxSfLByDkj7wjMbURPmYDJEEqPmww
O0nxMtgx5if0zqbabXguQgOwgWcQ2Bw/ErV2cBlgZfReYvuquwL8woqSlwMhoFPv0xon11doYWrx
OpKcy0A1c5SUPp6GvxU8KZToq7QwX+1QQigXjIbpoX9XNbj0jwLhxOo+rY01Q2XyGgxT54X/38bl
Wz++TBimEOzXlNSF+wNL3n8PqkiFuKunX8BNnGzwGX+VkoCJ2c2pVcYqeV4wmP8Ntg5PfFz+5uVj
CWIvo9zaOxlWCgSWNqk28Eain80kHAPR4T0ia1bjppHhz3+uEG1l0+XG6LULYo7bVbR7DNMg9Mjc
+9YIlhY2h5CyPtTAa4fzs79r5wHsfxaig5r+Q2fLqpWl4KlkfcfJ/GLbiwzK0cD8fSVT76bRL6Me
AuyOkcDJ2hRB0rj9ogW56hrFAwM4QMTTVIHNK/V5MdBG4GbsJSwbRxieQUp4k8xmiTFv+l5YYBD2
03fUXxHITXSjkWGwaR1yPpQ2LUNmMeuE9FKtWAOHKbwyvPfiFfURH4RgGRiiCtDvMJ5E6PDBrKHn
Ik0Ltgj0d/mFD0qYYW0LYrw2sroKww5kLMYMe3xG7RaZjaLALg1cInNMA5dLODlTBU7cTz+oAYgo
gqEbUDEn1WGpQoUSKz5qF/JbvUuzGoVfOJCG9DDsSvMw1iIL6Qy6vgJ6wZnGkq7lHSTad2YDyn4w
hZaEpSajwooFWb8DULpid+3C9ttew8Yy+ATJIuy5YGU6nEXovQERrWcr8kqQqvAIKcO0blbXb0wP
7O/AO9LqDq/qF/eJDvR8tP0/EP5eh9VbeLy1Yk6izs1MfHqZR0TqMTbsZUFYRBQwhnAIo6UDu0tg
FRItleEBDnWCcaXVmpbD9gj75M82yjYU8xsg/Eq6WTwzOtafNQY8s2ImLoz64XbK819/05UQ5ySZ
aZJMhqGraT0Mg3JbDWdGxes9sYx/oU9ySQZ7yJXGqdLXnqRuLAOaqmEabJ6WvUYhuaGEBn8Mufuh
JEa/A4dPiGOnXdxhb+w6OUDOMT3tOrygNCjGyzMKo5W6CBvw5g2pWRlyNEbf+HZgzPBI2jc7OM8d
Wp4q7iBFlsLNZ9EVXvrq4PYWnFtWjjaWSvkkVDpx5Mha/0aypZGUHd3y1QrXMZ5eJkeZlmT1+PDp
b81XXS2S9yNAbIGi1MEwsa+iXYUTJxPcgGx4D1QZ931LTWmMinkYqIMjO3E2cJV4ka+72gPn0ZpB
NvnFUIHz5QrzML0omuWx50H0LemFXjG29dRVCkw0cUlG/6qNMM6UavT/6QdgPUMsggzIsBP345PO
NP7sFSdNWvsEgogXAbzQDox84Xf8tLpSXvZhraEqBnUImEILV0MD17BuUWGngIcn74xfz7w4UIxG
mBdLar7oDYhu+BiRD4s3M5mFNWKyWYm2LWRQ/9YhZLQ8sM6cm++KfILI9kPKxmo6yT3wlQH5rixU
VQ8e6pQXXDKVdgLaLy7750IuqTFOHoYpZu85zZasNR97zKOHIfZgns/pHSN8mLPoVR9cbqFTqzep
xQ+sjG1DRDXwsi7w8n/g7vwRBHrBGcQpO/ddlTkqRQ7i/OTsREk5faZd7GVw6G8kOQqgdlgwxX+n
CqQOHH7G7tXyz9/15Y8Jsq7CXNgxnL/Krbs7eH6pVrSDIBnI/6P0vFMLvPHNp4gUCneTD7FOSQ2D
LNNdjUaalJGpA3G4+Iy5w09QAZDcFgCm4Dld8r2QPjDq66m5fUzT2zUyBkxiW03NUCPU2wW/SMtL
7mRvF06d2FMbT8nGFxxe9YwTRhPMREJqfZ+Dez52rsAYNgJlTG8pLP5bHYlzm/ZPDljh7QEmnVhl
oBh6vHHB89KSVRDUwM2UZlTNSOImHfxkzSAFJMPeyVgLP/eULjcXTO2NiU5D6T2OC8DmqFBOZAH9
rJnQ7ewpTfNi77dqK5IlXUAbA02sdeobBdr4J8snVIyCH6MRZ5wGRf7PcB0zpunvHk0GzpkCKfc6
uiq+LpVFOp25PBM8Gw0JA9e8TUKhDwC6sWWJ3Of1OGCfWciO1XZ9Us4xISzXAWPvaa/LENlrCpcc
8lN7IRY77LES8mbb77/QkkNYLShxuBkj7/4LoTUhw2AvyPUHuosDgwD/14QEfqivAfGB9cJI9aB0
i4ELA/VT6TgWiBwFot1+rstY8GISQ2kMYuhNVOWqn7Jx8+ulABMGO+kgsQCycSM5Xkx6tV77GnFd
ysJ29jq9oYCdrAHZ53kS4F8cef4pJMbJUHibakASD07ho4RMnYlPwDSOCzeGzCFfCJo6GyWvVe9B
4ja57EnPZTLGCfWOcqmKl/C/8aC5Ywa50ggM1NnLQpcQoGu8Thz7FxdrAWy37LFASAtEtxE1P/xb
sMOkipwRQ9pmoBaGvp1w90+XrtLiq1jg09AMNZ+J4ZV1aNvLqePwUynVWte/LYOPba6Wiscpz037
V4jdlR60kOjzu1G+ksxmbhZRV0hhIwvxrXow9exARJFJOHTOhUvbR9ok8Xh1y8NOUTSiFi2ZGx8a
ILLC8OE49etB4G9MJy4lr4egCvO31a/eJ8EcbLE8mO0P9jRu23pwvuKIoEgfMP3fuptlif+De7Z4
77php9Ld0KEj8b0uFDwRSfKZQeycgXQ4leZvaV1Rt2G47fXY97PH0MSRFNbBJRrW6NMw6HVrdlh7
NCB8BUwiJ8YzDozJwlWx41ndbs9tdiQkqy6pRFjdctT6omyy57rGB5VyfYcbUmYExUuZDBeDiQfZ
06HhcdE/E+JRIdXjyhVc0WW0r1jGclqFRQ0rDkKQVPNC0djmD2I69jmiLeEBJgOTq56E+VMtXfXE
6j4YQ2oIw7ht2+HeJOVYtWq7x7sPfMP9veJPojo2rt6gHAPy/MrNKXWArzw3DqmoirQkrlG8QW6a
/pRAUgvUCYY7YRgEY1yC1q3wky6wTq5Tmkf+xNydZm9OV4waiD1/UMOSf82nTRj080W9kVMWs8lR
jwnQMbGBDxEaIw4Mv3h2Hq/gbd1pWLDYzQ5BhT02bNtrZl/o16fjpRyp4B2YEzyqbbArFY6JfQOu
UEki6DkX+PPCszjfSHnU6c0A+8gui8tUNz2y/vDAKKMPggoffzCC3QFq6Au5ZuV1nv4hndM07wxs
cCJp8X/KMdM/osQIJ1aehZCKO/gnIkoQqklXcCj3lQeb0ljKt/LkGh5f0UXD31kj9AOzgyMaTQGR
ldvB6e5Qv6oc2x3rbAaKWlw+qwCY0WXxyxa5vxxMtvfgfaS/U0sWe3PpD45j9cbwGGievlcvll8u
AqDO1z/DLF1Ipr6nCRhr34mScBN6O91J5J2lj4C64ctrq01fI+Wc7E9Jk/DKtfT5+A1f8YsrxUlm
ekR51chCLP5VoFZnfcF02cwlwn/1ghnXdT6eyNl6N9HUg9jeDjfPWzZdpTUhp3Iz1gNHADVHHcH8
ZZwjmdT8H/I7cqDbsZBGHj92w6k9rwLkzzseGkFj2QpYbhkY1nSKrxCOMvkZeNLkqGCfhyJjojFc
po9pInmf40cgIDljYwyAQUpEqW0li6snIMPWILfM3ss8QRcQ+zJI/DyZ/FlHVqzGQ3yXoZ6p8vbq
MC3YRUwJaRJUiI/SwAsM6KAaBuRWtaDDQG+Kdq6K8kYn76yyShNjSz3wMan3LoSPMOBHMJMQVx4A
0FgWFA4hy1c6IsjmZ37nNfP93kwnKxDbL81yPKyQ2PitEDJdYKoOawvnbIwQU1fHZ/IZH6tG/VFt
4EeTPdDCpSpxYpC6wXF/vK+z+S91w9zULsvZOT8yaI2sVO7v9a5Mjo7WtEsiD8BG4i103Fntf7/f
apPgjjEauC0sXWJ+liJT77DY/xwyeBkdleiuFNxHiWK0L42Tozlufko6dX+Paqqbs2d8Tz7Ay8hE
vCPy3dCAoku89KoIycacfZnf+XMopfMg13AQ+XYFwMl3+//QwNmy73fZlC9nl1NCJn3fdbUBGTaI
AQmhQU44Xq4MeYCESR34MyQKoZDCaHc5rTm3da8joA/nD7zOsqO22WbmV/rYajxnzNikbbAfUVEi
gN8X2yVzodTpzIrh0/AJsI06oprXE93pqjqFaeqUqju/x5DVze+e82J2LvuYlMxJkQTBPaqwfmSB
OtiS2LDlsSrf/dJvsxhXs2tgZxOx2HuUPY+VG+AQl5OOBUhCby+lol+MdbU0KRNp4qa9SBuAsd3E
zlnOy9B5fnpBlhcFSxdxtjgGoj7fv0JZU113KVn2+OgT8yF4tFeU++AlqdO34vpdS3qd7IVaxUMU
0Mxb9uMyqxQvp5fnKlZ3MkLakpPNCAUTqpj45w0YlU/TlsRIS8x/AJMdli6BF8TFR3sgH8LU2SH6
oU/fvcOh6shPicYi2pJE42dgy7zqqZz88IMjSscXT7wGkEgnU3VymEqcJMu2hnNdHLnbebE67DMI
nPjEXRePMeTRHZnVBvoaMhOt0yJHphH4WEZsXIP6poj6M5J4v1D/4DckYd6NfSV921UAPALO6ntf
zW2l402vytV7VXncgQBm8ndpVziy5yW5zvXUL80BjXX7SsqWLLY1motMdRJw/mwY2HwOpGH6hMty
I3w5ikR8MJEwRttkuz9dPeJG2Mg3YkYy7P8/LWzvCf+133fuUG4kF4Q/XOpq6e3w+bYmH9syQP3R
VGDHoi03WXkfmfU6/VapwjRLpzGtQ3kpTIk3tDO4WyWkQFdJvZJvG2utqZGmUiX/RwVanMm8Fb/E
2SL5w6391NrxpBJOZx9EFTK/yeV9eHQVjliKH3oQts0+/gsmmuEIu0O8uE2Fd+nxKQMBqULhNHZV
UEAAevbGOFiOmRPwbVW4R4fi7xRBSEHmdfgis715AZgWtUaMn5Pzwg0/breDdOl+yPG5kaoiKk3C
Yei9HHir+TfLk9GZBEWtXdLB40LJvZYETSgnswGzkn9b+Im9qMpewqKNuv/h/9lqLsu55jAgmbqQ
YLZXmXF6+D8pZjT0St69kmw2iKU+Uy2QYsOoujtAJ8hfjiyG67TuoGT6ZFXljDEtgUDlJ9mhLkDl
e53VEawYNVQt4ExqPf0cd25HHpO68S17ZbtKy9g3urgbw3H5oHaxeGLtCLV8gVwAmHcVCBs8cOqw
4cg/ZhTZMqOIxlHGYvdWPS0QPqHU4FyibZXmMlQljKJB9+zWjNLDEpxKqXYI2JWNM08Lh8qeBltB
Iq0vCiYJTKm9e8knN3DowdYoCazgpVGgmcIx0xtb8lKcsW75YHgHOiu9gHUBhvvtI/GVx8dtJbu2
2Av/udCs5AuOo4vSbIT3gA2fWu2wJ1V19oF+cishb4qy9ICvEiRfVEQVr9FJCoJ+dcNyXUFxmShp
s7oPctxn0htL7F9533wXfyI+RO/3UhzM8wiYv/Xlxisy9xF50J50OmrImP3wmR3dvSvFAaP50Cdx
4MKleVtyTNmL2sXrPKGBAtkmc05R/OvUvUVKb7XEsk0Mbr0aEOEKD9th14kihYzG2/4ppbjivA3s
jS2cioLGQ6G6Kk2ley9F1gLqFyx/mXx3/FN+/Spkrcjsrx3iat/38OBp3r7+ATgDfEAQ52rCDE5S
k2WeSJrBS4s4RTtkRn9rXQNi3SGwYMF/L8V8XIvg3+7IstlJROomk6//X6nLHQY133fA9xNLx9eS
kx32ZkNLtyWP6XfD1B1JeBp9pv4UKwC9/g/Ki9npR+/zrHkiJcRYAr0ErVrne75v/ItOfMq67IF3
Cx2kG5HUktPSJtdPavOa1/DiiwORqtT6tXlBgcTdHIWwz+7seKbFH/pr7QPWGPI+KUuvTttDkqVw
Q3Rjwux9O4QEQFogdJQySPP1Qg8Cd9cH9fiMGRF6aDtTsyYB3/XV5E0cSZaTetIP0IsGO5a/VPZC
TW3ncUijTLA0cZcBaerecz+CjFwvzILpMWlfDIeeuMVReMZG6WngP5iy6TuXKwprt01SkXhudfbA
5T3ykG65AAPglVZwTaNhAJTFnMkRQqn5TLcE7MQTkxxun7eZWuHiHFJvRTD4V1+JZ5xb/r91Oe2O
fq9kiHPWv9YK5weq4Orq1+mkoJGaLC+Rp2lpi2cce70MNrPHU8TkR/e5awuF5EbWcCwa69J5nGDK
Z0+20pUWt9kp7tFTHf2wC1OML4DwfoDLUdHEKHvFYjNHYRess+Qo1P4BpXcizuCFZoRiZ7uY26wd
4QtpY1vBzPLVPQqFp6og9aOJX1mgnQfxq81tDrnINHIgwoOUkaz88NgiyHE6M1OGQz0ArlAv68yk
B9m3p6zl7jnqniE59ryPPkb3qh5fYWSTUlv1f3NXtVG8NUNojxJBkY61HGH0JDmz/xgJJ+x4DENJ
v9AibUtk3uISzPP0O02fUl6XfWiPBTq2YAX8HEWBtU5uEEp9BFL5/qanSTVFD+gZeH6VOZCDGb0p
xKDUMf+9RW8epwSF3CJDHIf98nyDDp1+Xlfos3WDFZ548VdQuqJ1JIAKoy5PWoCnUBIW7NEommXi
Jjd1kZY7yp7FrqL5DYcR0L7UtEW4N9ZuxbLXsuMBaut6zSXWUe7A0OCkA2mtCGMCJUokPF8OgM7N
Q2fEM3EOPE+5Y7yD6Z5/wjrzZAW0iRhywHyJUB9tMCKwGRXO0rTpROmb1bfs0xBoI6gHqTU9nU7s
sBCtaPLJhDSj1etlvbsHbjzYB/LioSdEWt/0wj9lGChj8872MgfDsa9npupFQP1NH5DjYbwwKEKj
PXihU+v3j8pvz21w/c8y5JHZL3ym3RraMpnPqxxMlYDDXKa3DT801Qd+XeESfVW/AmFqazhs/zMn
6zd0Z8rLf8yRCANaz+uBzVHf+PhC08L4Wfzn8/QPy6wt6BlQ6efHk//BSRjdfnEO/uoys+f2hmkI
wQhRS58GcYLcXkgoHwgewBdE8or9beUtVYucW8a5hUtAh8Vlvh9O4PJjG3mSnfj099RUaZTyZ3W8
U0qJ/bTxf9Bfhc/6B/sUiLaykQsBhdHbM37sjG47fEzKLphpbXz27IprLBOlB7/ZbMw0EI5n8BEY
fHF53JzmecCYfJ59YhxB1T+mYh+N42xC7PV/ObFP9gZX8kTtYG30xx2MfyFACsvPJolHSF7iHHx2
MP0N2Kp0XFDti/76do6KJxqzU2zJfKLtLYJMP1NkSGU9T61Y+rLygLVHafVigaqiH/U1bFwfeyx9
l0qtVPquPAtLzCKhotyeeyS+t7OcNQJvTffxhpTuw7xo8h2rEYru3sl1roNVKTY81WODrViLc5vo
cUjyBiYyqHzODGXIuG5D90hpJg7RJBF99a1nDHzd4TLQAIKYuSc0JUqx6an00AaR7XwBGyhRKOeN
wpzRABDzayZwcrmC0QoEqBbMJIcAZSYZWUuznUICZRlTlncu2t82WscukDY9hqywRDWm2VU9g6Br
YrmS8sLmUXk3TfY3Ma1GC7fI/MvDKLqlw/lbBGe66XVV+t0/SGWOcE6tV0UMHglYWb1eqKZ5hxsh
MV3tDrgUjsfJj/z313a0ISA1dIvAoVAfmCFx20gL9iT2bTnHsr7ljwZXQcNr2VI+ynXyur+rkWiK
Bg3auS4QKAt9a+GnsEUXXcBMEv8Ys2RRnBcgXoVr/AIgZEdVD0SxfauV15W1pldYtxIKv8oydK6s
pXMmrqo1McuA/6ZGTvyzBKNgd4vSB3dSD5S4rU5yY9jgxVwMw7W8JYLXsAYkvzNgtS8xUhp1LZk/
3mpV3G7XrEatR7lf0+3TNsmHUeaQVar+n3Mdf6D3V6lEgCtKUqVy5FfEPPsBXRBpPb+IuaWjtoY3
KkjLsHLingoX1WliZPYS6vv+D0FXdh48MJwHFBTS0ddt3rUPHPgqiUSWSqPUt9qO+mJO6RB8Zp3i
8U0MLtnwYBR128HR55JVHOfjXfdIhuMIbcdu7jnhPZHoItFIsHCBq52up6juRqyXpqZtM4twfc+o
qamQ02fsM6szZjTjuyaLpCKVqLM3fcPCnEdr2fUgWSlwMCh52pMzsqOCS5picI4HOlOuYFBLmuxS
VLpqmQ8gZwr+uSKv64EtHqdvWzxWE+/pmAesKJcT6rJiGLbq5bg4X4YyVeXFRvKNoqr/GLUSgUXz
gp7HViPXdqflf7Kh0APs5Bq9yydjAexfjwrsKDLttvgkejzqND0QBrdE3+xnoF1vM5nrMXaU3u4X
J7lIWyHOFGbbQNuE9ayfnfl4kMsX/p6WbBXWt7GxFUMaXipr9u9xRAjE7xn5rUb85ExIydyuJWx5
PjPttfDGfeNVrynfWnvQ8ScDHyLCV/qGwjikRHu8SmfLupJvF/BEL4861zwphpdd5QUpPTT+AUTG
0hKrawkrAgXOOCSj0zenyYS4F+BlFlC5WZniZos7uHCj6wQ1A6j04+Osl8RAhl/j7VDnuqvjBjpq
w3G2fYIv0ueF4bdKRLntyMH9FUgqXMQdLlGZUZUeU675+aOU+0917aQRiqusARBb3pnfGjhKuO0R
vcdkfzGY7YCD4WYYomTUzkJuogPBYAsO92hvOBJ/jWa7nHyBEvwucqZcryvqJyK+vjXErjfDoCZh
EWudL2vNe+2Cr+13x0syLVl59JuA1PB5aEB1zxQP2Q5MkSh1d8qq2RXMtr+fljpfWmTXx1TAtaCo
aLqEBCh5OcV6Uo+L1axEzGXORmF3hu9g29+AzdyUFOjHhahk+gxC5B0+d+zz+5eMaIf0v0/utDHD
N6Y669mPPiVodRmwklTndTouTe2i0qAfLu3Yo4lAr9LYipdzSU8I0c5PwSgI2uFRDHloAk5ngJLh
1C5786oreJRp0UpOq5vnHL2qgmAqMavvbQfFNoQNiqRge5BN0ked/MvLPHrLldfCh8ATbTpIHupm
3wp1ms9sP+Sg9cR9Fb6giGU15ToOHXwL0uwKzzW+TPcZ2XevUTeQuD3jgbhPxwgyvzE/aWljAOnS
+T2U+XNkSmjwSMcRTSK0ysUTu1lf8wHvaq0e5ixoIdO0VAMhDkDhaiqkUNnt0vSZ/Hoex0MpXhOk
8aiuHtHhPGaAS2hxzM5BVLs2RF7UwFIXDkF2Rf1m1sBYD6SLBrG+hPL8JAJ6OcoQ9bth2zAr+89t
YXGHfmMyIoNVPucUcSbXY43DL7whWx2Q5GQ+txqX64GEEX5WJO0kdAU5vHMIdu8blgfnEZCo3skK
dhizLwBBNM1GuiqDZ5q8YPAPIlpltqaSzWQeHNMkIwb6BF/I4z+8k4IYaR++BAcIJa7rhCd0ICqi
tuRCh5yCSzVyo/m87IfF0OFejgXyy0N4q2gLbMEE93WMRT+tIRdrHCdF+Jw6XrfH4IGJf80PuzOO
YPZaRnrTo/M8iTIuYVu/p90yaKczwDdE1jlGy6VmXgvVbDzz9EUy1syC389a3dI/zq6XB8hLZfij
gcGCbuNAlCCih4o/3w+hNVSVQbCo6L/mP26omrDFZzazxWbgofr/7oABa6H8K4wEQZNl7+iMuYhA
J3J9oyoYePOLG6b2so+TBDP+ZbziRfLYd7XEVGv4zEjdjz1Eg/ekP3380TFCseYa7gnvt/VgmsZN
1V0aH83oYxgXwzEmpclnBZDiLaLTY7jb+p4IOgCe4SQdHXHpOJg0vEgOO2zkbNfr++EGuTjK7Sme
QrrAWBLzHu9Re6tCJHyx70Z2hGrCqcWdvoNybCa9Y+VvmXXNMoQkf63r/1k70QZnj6lH33x6h19r
8eSGQoS7ZAZdkW/lv61HMmFkcsf/yOtZgc2bFSEFy+613yjZacv6/yvKcyr+7VXatHQLJ3O6HSkW
waBtOnPf2845nicGrrJJiboFARyRAPCPowo5hzl7h9B0tKAX6pm4/gz1V+MSYyWFNshGtZitYCQD
/S0QP6EZOlyCooR2Pfs5ejnT8e5aWlSWy4+cfnyuRwaDl7d3wt960as3LwnittpeKGVps62hYPwO
Po/GJEGY/P5yycZBp5IE4dDUCuQLAfI3T1G/SgPI5z24BQ5t19xfbEjEWmCzRasbC6ABrPzCFC4+
/0MvVu98S5S9DsetAAsb8OaFvtSlFSE+b00JNyqS2QGHE3lUCd//t3DxtvHD84kgb2KdEB4qvaAA
5JnjRIGEkZl8tmGgNDwqwJH1PgOf/1aC0CbLE+E6vzmoIhBVynNXNSQoow9fyrfHPpGxHtdenQep
xDhKMYnjF2O70A0opNmo/NXprBbDsfsRD7Zx9ciQQNFobPwsTPz4zu+ZVgmz93xzwVvruTg1DNWS
Eq53xRZMJc4YTx8XeWukN238M2oijKHuEJWNijQU5Ux0tgV3drxxic3cuLgiSavxp/tFD6Gg4Y4U
QKEoDGd4OR7/nirwMWSdOoBkiSIoyaCd4llDKVOSJshka63EMczT5H7d5Hv95o2yB2F0y3VWg8Mv
SAQ5O0ZTLljqW3eJ3PKCr98fsvFulJL0MFgHCA2twUJHstFFSgvIjnWIEuXznBL58xOK7o/rSSHS
mkFFsMZ0PCIy2cjqHSkJcLr83IDsNo+it5BYIX4IEEAqUl6t7B1Pc0wigLRiEsm5yup0EeN+pPT8
N0cOltVOP4PkBFyXcjZOruDzp/ycKX3PEAgLJEwPhx0ukPe0f5SmvQCvv6QLwuzIRvBsIGdEL18p
SD5WJ/yAqyCHWveJidKnIZHvfQq0oHX4Jy8hJNl0H7+PPc9H7WLRs3GR/jQTpL3y4toHjUjXKCja
HcISU+7fT/4p7hrcz1h3evzAPapOmN5G9tLgkMV8vvWVXCQ5iFO5WpzcRzPyk7c/ntHQvQHYsNVF
NcjBT6LxiTaGymLodzhjxnt59bXwHTfT1B46iBwwj87dnWC6jAdfmdRGRx/KPu/pQHli7KnQlpcS
z/iPND4kfDa2frt+tXU2UHyymHwNM424t5KNOik/FAWC+e3t87ZQ9mo6b0pYWtJ0+KJaYujHGefo
TI4qJRFVU23t0P1mtHx/e9J/OVzf1YmOTro9/xNwOgQ+dGH/vbH+I1yw82HllDQxnVC6b8ZQT/hb
kuaG7sNrZ/O13bH5bzRg6lRAh8Xk/mF3fvBEUFykSlZqoHsSeREQnUvQOYEQ4fUCcILXwOxwORLL
OnCaSMd+1Ekjjd+pzr2cAz53lCSawc3RrpD3ou31WFT+IFX9xx+7U9eYImroaTvocAGuUQms/jhf
pDilh7jU5DMcjmzJwD0W/6mA+g2CCmxAh6feAWfjpQNxXFIVnk+B9yWF9MaRmepFeIPqB0piLRY3
JZKv86j3kwiJmHIANdBZejfzMnBoIhU33BG0lrxzJShctPCBnoG81gEHCAXFkzQMVfWuDHt82YL7
o4A24qjSxh6Dgkr3nZVf/PhP18qWLCRZIlvTBGx0b0ZV3nTosB66vXZVJ097dTEoLGPZX1JW8BPR
FiB0x1XvqSc1JoGIVaqaPA6pvwN8LfY1bn61Ieekv7uIuFYUAFicsr7u3kdg5SP7eUJAUJlZqoD7
fiHda4KGq4A0Th0aB23jeL82iE/ULYTivxEkrXx9koKTrpZcSnvF/fgpbEUB/UDEi8qVC0dLb5Yj
JNLD6+A9y5ZHaSWEO+ItzpIp4PQjvh1W3zxhkWa8IQq1rdwU3DP3NZfO4PevNQmDflkX1ATM/NrJ
XTubcBCH/FR03gUg0wVIUtUf72nQXjUG1HOc5l/sB04ccJZ0VphOQhty/Ntst2x8rElS/KGbwVBq
s4gWNJlye9+mQBPiDH94xDmkzddq7RXdr3wUhSmWqNtdQLxKePh/GWzh/+VeMSjkka6YvQ2KT5ID
s5Cd+DDVuXc3Srct3FiYmx+hAboVs1HZGbtX708fdSUH3ZO9jTVJVoLxQEpUqLOdEhYbxrWlVBFD
/+5rpu/maAmFhBvxRmcw8VpuecZCWhCvx0G6TINnoKtLAsRZIZ6i5MXaNCBMd/5Ktr2p9gQeff1j
41NEj1UvEC828e4tZq79T4OdRRGkTbg8W9hd2Ixb56zp61Q0tdZ0QP5fWNJ7PyH/uHl1MJvozvY7
fYCBjGSpRYDLAaWcudS5wTilQA1DH4HmK3IP8HaPardWPk/Rl0JaGofXxYhtpzQvdLP0eokTe3iV
xKZYRste4PfNc9mdIBU0ZOzGoEu1tD7D9ctBlOMzuIpVRKv5STZysHCdjcShElpdy9dM0asP+/10
wtFSQpqEC+WdlgfEp6/my5A96BtAKgH+VC0WPcjGrUe21tuxW103f8dgNy/qtKgHnRS6DcKzBUQh
Gop0opZEGf7fik14xXQVSfUdZJnAQYRzZAT+7mFbicBdKAy8JFFFtDeKxoFHWFr6EeECtJNubDtd
cRb2GMYfyGv7z4anU9DdWkSzhDvojs8R1TNWoI0SiDf0nBnDWezbBhEfcefd6aaskVVdwWb/k9o3
ZMTyhRlVByErzrmoRfmL/mXgE2fwddQq1Xwe1Xoq1USP7Nn3D955wmUKiavKt1P643ohkN25m/8e
LztM+LoDe5k7GGsAQkqsK70Ibg45DUSsCwTOtzYc+qkd4jtOohUsiNb9pBrxVOYMPjLZhTBCQYCb
vHGlGj3ijXdh5XkOV8HrmE294LlbqHS8M+CmnUgcgwUHbkixP0ySEBquNSfGYYNop7N7gb7MwAxw
YWuHfnc6Co2EqY2l1cs9YTU9t0Lal4/AaHOd4cW2lsqjDY0eop3wC2eQi+cDYYv90bXTKBRyZibV
M4f2TXpaqOCY57Lof2IYKK9yAlcySqoXeMDoSF5SFWGyG0Il3oLo+62UhkCBquTC/nUS4mgHJION
c2gtHe3OyQK7cHMOkeR7yClM4vlsFLftQi9VszE+X7it37szaYT+GgIusQ5MD/4fm3IqXHuxPHUJ
nXWCi5KYLfmKMXWLxdKsXqf34o3TaSsc5LD4Xh5OzBITOMGBi1Xl10286gBDs0OR1gUKX+hUBsCF
2cgAGw2Dm5UgtHTybyEEwrnTgytL/9RVLDAdieKLTWBCnjAns5FI2Cu5JlK8mQWVXtyJKvPhDIBp
lv5bk/sFW97QbCkKgyYjNlrkIjGmemPJLrVKofuzGQ9jqvdeALa7aSVho8FgKBzphEwFTABbdht2
LY+JykRRauFDYXvu0xbuSkOFzwiKelYyC4fQdBQ94U2zxOoX+dYXAvV9E5YqT71vYYRr8BAoRiRV
5LJJaEyZY5Az/HK/151gqjA7m5gghaRNvNXG6WYBvvMIV+T3bfFrAmVMc3dMA4tO4/B1P8NSJwEc
R030OOTYTXlBNrQgfS2t6XExlmUeEhIiylw3/+MTgCkc3/6ftldmbOY2aJ6E4bUCNl1hpS5DJcpu
uuR+8lKjSCzGx+czefMqt2KSYe5GpwljZDLcgv6qBUvDxALMjsiF7A9do2V+zhY1J20y7xAU2avL
SMMcAuaNZtPmVXKriXTRxZ0AtEH/YhNmW1UbwQUBIpDOiSlNNd5vLvETu30JByTjNc/H7MquFzW0
nHrD6o4xFrAmy4EHX5o5N98LOi0aCZqjuQMz33msM1xg0hT3u+AdSIHFift3kz6j0E6erhE/ivw7
U2kla/x3i+RlX1nLCo3MGjLy73GHazexua9DCkAUVwEi9w44jLPlgcO79NJkTkQMs8PbkR6SWlsy
xWVnM5eYhVxa/OhWLx9G5a2rLpdh9nkuCFtrmADS8ousesPE9nW3xCMXxy7UONz7FjYdXWDPSbqY
PX4Lo1y0D6O8z39sh94ywwwBwKfdnLkaBxBNiKmC1Nw1j3cc2Wkrj+RIo1SlsZIi5+8z1ANk9Rvw
+t5r1xCZ+B6hKWlFznsyUIwB38vmjf/A7+4dngU8c4d0wRI0aiJbgP4zi26F2BlsQl46X12Mh+Wk
qOB/NEqj74Bql/Hl9J2uyhRpACOvwGCLbXNSIB5Gl2oHC07tvSaIVm+yGD5T8cRN7F/19o26gEXu
LbLVzTHh/lFSJYRLgnWZuDEh1q8CDhokItgatRDX5iGluoxNesRFv/6GO+kDolCrk5f3S5sKmkto
/MxstK9Lj9XplSUPQg8saaqJ0G4kcb+lukcMBUt8tlMKASK1kMmnjEALnwJSbB0ZXd5ye+dnon3E
kfmZe9LzT4YaEv2v0wFdb+hJevjK0lLJab10vMV9DfxHHIhHZQ+mi70Aam/I4KBi7SrDoVwixM2D
oZmfwzSR5U7tvVVdoX4kMC2T97du/jE0W5sPstqAij7MfJqfjICxRk/PcsGvOcsBJ1vaFWY8roeL
g6eVrAT+FP9XHsg9dR/AqzIvpr4pqf2IxN6OHy+3CW7VSL7Zr/oi5Jn0iLZ0lQCZ3JuSz82uNCEO
RVnalpQBJeFKZBTaUxo8cc5DjqG+93JrvIM49EcWHceoilTXnGBri+OeL2fNyUwrqWd/XYmyNxmK
PfZoxBWAaOrx8c0pYKf9Ju1Qa5HTe4igKyFVEp0pRTdaymhrEsLN43UybxluFsl1IjaEz2xjELJq
bQ2gZaZ61+o6Lj53CXkBZX4dT2CbARYlc43agfrsKU5n+IXdA1CpcZNSuGuupxpL6IaLn9gpGAcl
ejVnVohT7C3guTnEe8iW5J+vj5FekeTC+aEMyLfSv3gEmXvdwJEfMab4tbByzSohGZVhAvDqRJg1
nhg7uXD9rWM4JZnn3rnhtpN0R/oJyA5T1jb8nJrRvm44IvRJN9PSgoSLzOV7M4Zo2aOf12mxIzui
Nz4Vx0EE4Z9hY33YQ6gCuPgq4QaGQzJEdopnXccLYnSFboK74eITj3o/Lxg9g/79crNL8Pg9G20d
WjdZmRvtryilsHKa2WYwpXFCs5bJA5Q+ZY2u57v6C1f8miL5A6yzaaGaGqM9WIa2Kifqh4SSm6HW
L9m11yBELNei/E5KKGUJAmTzJTRKH435llkyATz6tQxjNnqEUGXiGhL29j8BwXEDO+9JGQuL4qus
dmZ8Qd8moklw6QBMp1hdRdEh/uLMxmEmfm87mexF88RXsh/TZkDq8DrMxKLZQwNZ91Z4kGtogjZs
wMPt8Xl3gDfTxxXkYE9cCKRpSFDZaWdlZSfpDk7Yz/YICS4t1HCmM6euID9JnM+MqZafzS+SQd7e
FFETKG6aYTvzf9LN1bftjcwdlcA0L0yCLMR156R3Xldh/bKV1m7X/wcE5XmS7naEglKWrkj2wp+d
Bw55/5gTRqWEzuQuw4DXwsJIEYxlW1bReW61IuZEuqynbXIkqofA+0RmE313WqC28m0MXylzi8LF
a0ZOJliP03kb3mfvazU5J5r7zNHLtkj7m9GFe65k2Ny8tmZnOx1zYtaehwjoyAEfTN7jbwEtmLFy
L/1wRuAsIDncl1O9R43cVRAzggLismjyNOZde4U11rxoBlxUrxWaEZ7RIkOK8Fr3wWM108/ToKAu
l5QkjjLKRuymau6JufQeHMKbOfTseaDJ0tRvjfd3hzdHHrC5UeBuDtINO2azj09plAbKNOBuJdUY
hK+9ncp7n8lrzt4VJKZxJ04X15PnA2vmGhbsgrjcao8RmQRXd7cRMp/0wEVUr17G+RQlXl2+IIin
gw3HfQK01RU/7LpGWfQSh/5WdTBxPqXl2PKl6I3FZAQ3ywxblJhRKwXuxECbOV6fDR6bwSxFayoC
4e6aY34Wq7H94a3rIzMzUmghr1zKpruNLJZr81iEnOwQW+Msn+PzTjsDVZmjxx3/XpQTq0yGvSxf
O0wrzYS92JsI0vtv43+c9xT4U0SpQzRMjSRo6qkPvA56GepOv/ZLsyXnwbDXTqkc9uLXot25VcAQ
m5o4T2Y5O2EDWnyeQA1FEDyDWvKmlMOaCb3OP2kd9Qi+BQTpihFaDAniQTlXIQyn0IVGoAJCOySK
6aFNzXgkP8uCOG4dfs2rel7kvDy4niHPSnB/CO5HrAmMntKQtTjPT0GSjp6LQCh7Hwo1icJyk3zW
SXpvu0dgtr7yy/cvAd+E9fizTjaSJ7qoT4Iu2SZMOcVvxGIh/UHnOV0nVTv8p6quEfnB9qLWuHWo
jm9jXj0LamUE+BNyUypFxhse7FkhlvHH9jEDyKkfkGcyWfeEl+5K2s9SXSTocRlLmmvivQgndpy4
Nx2OjmRyXV5u30hLngI54fNAeQZH0ZtJay+3mBjAR9DpzNrorkieNBaqtwIqg4v+hi5zV4MNr6pE
SQC2GbGNFIen+StRsuwcF8rzBOCNSn7DUVf7BVeRVVsQJj97yzdlRta584WcwPiZrXX/eq5Fjup2
3q3bwaTTHZCZasmQluB0T6pxu1Bj5ghwrPWw5xMhnSbEwZfnEnlAHhUiO78Twh9Z69NHQAAXoJ94
YY4XZgqaOyHqv8WK/a9joOp43Pp9i1K45B0JCPxbwAYKX9cZYFELDUHAjjE1LwjiwMRMluVqZKLb
Fhgek5yeZsXuQGI9SB+fl+25i3ZQAOyqWNHml/bvzXvnqnASQbpSAEu3nC1hyFM7/zDXPWEL4lm0
nqM49/sqeSbvmfwUADTSXtDxS6PX0rlnD14cnVE4tFYkZHtp3MtxU9brwPmUAs5Ja1/4nqsLChIX
Ztu6zySuvNstMUPCNKZ1gREs6t9uRT0aHHJhoNOKfC49h1rm3zWZTnnZUt9RHkNKNjuS/kKqjBD/
byyYW/SmvLh/O4qw2/XEyFS5bQ/uiM28kiOia1/XWQyigOzduWdTPrGEcVF51xXLZURoXU1ZfR0s
YWPNkXf4S8u8EOHaCq1/drFpIbh46e4NrukEHNyYPvEWcjokwq0fQUsiFoixadv/uG08d+oya0Xv
ogU5t526gQwPq/S91f9CMIM3o5u5+GF44s0hJKCGIZYftslx7Qa+avf/lWvejdVpVvgEw0XPo/jC
P2QSwOlyf1Yiqasn/znFiq0Z1S4U6H0W/EvUnxKbyv+yrBNTXq8WYk3zGpLDkjkaZisCfmeJ662K
e+23C2xUxDnJ2GGtW6Xb9PW2KsWHsRHYFzZuY4SLh37DuYYdgB2AOkP9eFX4rhjdrtPc0f6WV09P
8s46GRb1ULAEW2Qboa+umW3uROPnCUeg5bekDqDGjLYc5WyywfH3NRDL8jnD+AzwoFmlufI3hMpL
Ernk/NdoXjpWl4Anu6BxYLGmugwnug8iQ21NEMCwygH1w2ystobVFXImLt2kIBzbl9SOiEgEbe5f
6ctGAgt6q43vSfLt5drzinkOfu7peqjobC8ttoDajeWUOKMyorxO30INWkhVUyXebwpL3W6bio6S
t+j6Rulo2Y4IjDQf/TWuJf645pw4IL42+EvWn0F5ya4O4X4NeGAF3Z/Uc9u5M783UoM9Czd2sRGd
alHbWxoR16S5PsBU77qQX9gC4k8fp7BuJeVyvFbsCLUm/kONsEuSscb139orVnBtE0rs58+WmqQ8
FMpFZWi00x2+jt9abHCTmM6Pl3hnOFytrapJCfJz12Om4LWKTFXyGgZXLAtYj7He7/le1h9oGpAf
rLSzGpCTAbt8nrOUkIUZ5UQNPvZI1ZnMuQ4oLR2hIpoD8xjfEkRUzXpOAfj8EjcMGXj3NAQonh3z
z92zCYzBjOUEvkaEinVT4cyEJoxVfJvqZwL6yEaKv+cPcs1O6kuZqHtrp7L7lv3HLIenCjOIHpxc
3ekOBVGjKNfKuWeqLOYu3FOtXm1CxU8EUxUzw0iIJV0xaaOvgyRUq0UE8ANem8pImXoneadfqTsu
CVSIsJGVzxUf5NVAAT/uGOOvqMfiaOagkQ/c9MA7rj+26OQMXOlYRyAPahRzC+4VjWEwqtEsDaAZ
9D5+UGPAnK+ZdgJX3Oq+xAPDUELU5kE4Ixb3D2XXuJF80JA6pbXXPjcHOg4Rm7inCQxhh8WHjHn/
CfDDmDiHYLG1LdjDptJvon8CNspVRP4tyOHHgy660Wa5R/mroekitHhOgXgA0rYY3RaIVWJgxuyr
v3nAbVJBIkouOTkCxN+EMyywydDAuHVyBOAGSKcP3djZxET1zLQZZeTVANL36Bs3eN3Owp0k//lK
JBpTw3nmwOptJxE0jMK6nMrWZ1pvM7QiBnPUIsYZ+958dUuvYeHxOfH1FDhUdIOktnMKCQ+VW17i
g7cABwTHC3QipRDJmd4mi9S926WsoNl2pJVR1eGmoJzvMMD9ZNA+NriuuznUjvjXrqwblqZkBd0J
wzD0GJEzoiDURB51ezbU4bY79EAec5tlLT7cjtHdwFPgNbQ2DGi76kGKd5C0OQQL8sFwf9HOqCk+
OxBCcD+iXQa80/lpXPbkZOnzBK82crH/TVV8osTaJ0b2hWNhqpF2m2WXcRdBFV3tiXB9fCNmKB4e
ovStieB9lBrPm4BQJBqTLgYdzpBuerSh+WlRG83cc/XYCmwjfGk8LquSIXD4trj6ImqijmjTaBui
Aq8L6XcAba1j5lCEC5yvBoDcX8mjr2JzgESWsSJfn3PZ174qpY/8ymugv8BihUnub0Kqc4QBRnoF
YLTkP6NY0gvM5OjYbW1v3rtlMbF/Mr6rUxlKgacnmbMO96qIkf4Piv0R/iWiGN58RIEw38y3BveO
ovBxGA0uruVi4suMeg9dxVzZLYESke8LDJwNxDwT+2+oNfGxt9PO98khYqonI/VUoO5IDppGZTzV
qOkCM/yF580kAARLKTKbwFXPs046NPHZlztURZsSOBQiromXxNT/kMP807U8Nk0rwCDy/4jx7so5
q4cpN4SROXHCnTrE9/uMNvJXvRajTM9M4nlZWBR388LxmHhFhe+CmkyBiXfN3hOFvyFFPoZ451Er
V+zGttek9yALmmYrVtM+o2LhngayqTPH4/rbMuPTEb3Lxf0Z+cnfFilTmnF/+PY6BWseihJ457ch
1H2MnGWXhMzm99uCI0z8WZILlxfxYAISMfJh0XvQirsBSm7F4lyCyKVCPzPsGR1GfDoyIVKOrYX9
9LmVWuFSHIibU0HojC4jFK/wrAF0GN9B2/FUl8vjQQv6bYQ4xVIKNZd4MkYyv2ufZFgwlhGLAUEV
yWXAm9iEXeNZM5g2ihau908pySM1AHvFyvHcXce6TZflOQyUSsX+CTPEa7aWoSti+xJJ19wo1Q3v
oWXRAKLoAX/mXfKS5Ef7MbqMDbt6AN5SCPQV7d6qi6EG8tF+qDUaHW0BV+gb2V4fqGj6ISWb8GcY
OiWHI9Hngip+oxcO3NhVqFrhL2/K3HY88dLDvLzf1xyxz2X+PckJokVjcQNRtGn9V1teyuHWRJUa
vVceupMfVKwg0vLxRo4V5Mr1VtmWfCNfSuML7NUsvxN7I4CewW9CaAWPP5RSgWTwa6q51+GPWM88
ZOme173aGDBOYTZGfhjR4v7s8cUtqwS0ukigQYUlzaJrgvdgVRDFvITDo/we0fC5IAEC1HChvody
QKRHDZt+8kYR9BV7JLMARZbPZn2A/Eb3HI7dHkXTJ3StbtrcNYGFFNOEMHmKSb3Ev7XRxjRxw+u/
hFVUQKe4Q8ai0uC1g5zpvmAoFrQGnk+mAODGEoK5BynQkmhBkb5U8gta0+2J8mrYWwJ/LJkqYwvR
RA1LuP3NkAQXTYXXrgT0amOnazHkQu0MhoJ8e7hBrVFyDjNLQY5q0Hya3zWKUyuTp17l7FsS5qPy
HCcl5c0MgbDnurwPkmJYgCYVJHMEsOMQQ6IVeV/VpJsycQLuXReCTtlAk6QwzkMy0o4qX8upTDtV
WnZkWcnTNjC/zzt9DheNEV+yom8/pK2Pt+/XHPOndK9DLr5yYD3s2+y2kbxGKeZy+5TiBpPl+GiF
gwwkgYnVb16xnqWYLA4/r6AaW6YpihD981KvcdvllXXEvJHOtU9eaJjRXhv9T1ZxIfzJc9RBv7NU
H7Zm3XyV/Q8sZ4wiMSgC8LLLgyn2KfIIkRiwQzFoLVZnMYlfUr7dRVtvb1bidWaNk9IfU7HTjNnN
JTm2oSyo2zMGIKLTdTY7UeyYgRpQBivwffwUj9xP0A6WfESp9+kFfJ1o3M3zFsmCchDLHuQ8VyYM
l5rgw4CoRPK2PG/WGlD/JrVFZyseQNJkJLphwHx0SQSkdVvP5Vz3+AbntzLUFnCPc7Tv4WuEelOA
qFec/PDRf9ASjDsXqnGroYQNv4SqF/08Yk+b5lBsjOixJ66r4EGlP7yj1zNc5QIPacpnEGcX7Hvf
8QYu8XPXXXUWUcXI3Ke5fPC2pOxeQRHJFd3dV7sG2BQbqx/Ums4WKzL+8/rUAQ/xUNA6j28q4h4E
YVtf7udennm96VMnC/g6MGFwjzVo39rAJIKP6p3Do4If6eb2+z0eqwFxF0GdAllZnKe73Qoa0g/l
QC4KlWyHM5t+cJ8iBUIkxZ6AwvKiOLBCGfBPcJjA4qsQAbFbTTqApdyKuTA9fnxeJdWmyTZneNIk
qlmHFMSZCUSZFim2GXJXwO9uAvcl+a15jwoYOKFyupe/OA4Dogt6fbhKBvcfBKj36TPU+9zRyUwA
xjr7FuPq63tnYRdx7PT4oPzTlxuyb/+6Q/3RfE03nOfIbdVRdSijFuoa7w9cNCqVvH/IEkrJNeoL
Un+vQ13DW7dF1QFQdVYDhWV3pC1d5YsxoNnFrg5F6AgZrbKJZUmQa6RQSTbW3hOweh7Gc/AiLOU3
dC92znvYmcCtLfbsdKzfvQcqfU4ghSdI/FDzcZfBbkYpu2dWOUXNfPtlx1a3bjJZ3tjNaMaWWDFc
tA6lUjdDbbwP1hMiZPq24bRhnaMHWUsbR1KJk/nYnPafU/yioQ0D6cKDSa4xz962rSASV2PlWz1d
YclyLc4DBMreHeSwL1r1hdNFcRMZLizULKVJkwzxCXZLSZB0TJOT/YyUNx7s9YL+/9f9QmLbw4OC
gg3xXdxRjnCKbiSoW+1YSZ5Ri4fvFvgPZSUE8RMdjzpIRhPeI0DtzldlvhSqbYv5ALTYiF/GST3G
PjuNk7oaSsiXhoKW3ZMl8C+UBCltConpVe3w5IQg5+yxcL3AI54/rB7IgM9KpNzrtBYD9s+MK3N9
eRLDVCjbMw0oCM0Geqy4Y0h7jsuRcYyiyzpISoMrEw3khAMu9MgHTUlrGGv3Mq5djMnXY075TLsf
MGFDe9nUvsUmu3Hq8Otij6w/HOQe2dz9H5yg7klhO+0KLC5SIyMkii459z2Cu/fs38vRhGMVoptv
E/WxssP9Y3rzXXMZ3KuA+jlk9q6RAgBNkqCpUtDcuLGR8dPDidJVbOVhrqbEPj5Q+zUfiHx0ZWO3
nRhiB2+VEGoRu4ZQy/fttqyCmkza/SPSqofcjhOiLQvKfbYn6vPklGLlOQ3T1e/zGaiF3dKkrhsc
bsGVQVFYZKfWLyFAX+7ghG+7CsKctxTimVePzTxz+5Nq+59X+sAVPto7jMALfZEJ8/pVP/Vai33g
OP9S6GtCSKbURWJwmChPXypadcObE6CkZhJIBYRK6cv+g/IE5J5jXr9oPGgK91itRyYPSw17tFKi
85mvzo+c6EV6P2ReroZgO/DjkjFcAbvNOlj6cUeHMSncKpaDWi35r21qk0O9TV741rSEyvoKu4/O
iknwwurVD/jkGGxkqqJirUJmCgIz3oPCU4FmHVgwDBaGNOdofyYewV6u899+xwRFiwEUUiIZa+S8
suOVX5oayIzMyOzn3PYON+0E57aAWmEIA/A3DYy+U1UWjRjRum88PxfP9SWjwHZjXuPEO/nB7hta
0FgF3sTPMzuOaTpdZGvD/Bud+87j9QwNWXxx4jg3mQVKfrlaibIjJXe3xNqdG8H7bdg6T11qeNhN
dEJVAQjHHB60SI9pNNqetFnDvH6Itl5CscCqf1Xqh54qp9sWxZFcMRwgrekwF9iNCBaa7vzlD7Im
PltU8VZcUbcJMt63EezOumq3PDsSIyD/plqjME7klxol7VZkUHkNTvF3rIjdMG/zGjjbGrLdU6Xw
zOkc4ca6ht80Jj0D2upB1EM1zGTX5FPpvXwABNKpi4zdYDERMwuhfsyzRdDWLPpyMWnWfIdRE4c+
wAKFtNSVy1qyjLZ1/3ONT03/a0UYChiF/feKXCPZFXSPkrpu954BJm0N81vjvVQGGxJhtF2wLNKw
Cjy2N5gp9QyVYklGrp8zPjWRvmFl/wLlQSGT2Kf4Is/37xjABxYHhThKnWY+u5kwmh5um2nwHab6
5aaxtQiUSKbeISy2rxQL/iysglv/PWasUBs5bJeJabUe1BgEK3KCVJL5GFte7FS5YDcvLoObJ8Gc
zEDxf4DW5FnHcNcpqqajec9qf562f382TiS3k40u83V6lQa5topevvTDMH7H/QkCeLhWigILcDov
HrobOCmSO3XTocl/m13horqQ4qM4+/yv+gAGTtxfLm4Sw79/VqZ3bmZK9NkiCPI+u9wAyzIxoE4X
ybRjf/PTtoZxh3ruWYyEpU86gPgmfElu8x4JUu+Hmg/iIvReWwDjDDJMErm1TQZC+vKHA40oI3U6
FXgOgNzMFcmTasJmsXn1vmnymg9rx7NGi7JFFM/Gjpmg97IIFPSjQjRF6pMtKASl35bbzNXMiEDr
yRU2+0Ptg9z9PS6XJi0dZ4a4urWVgUmh92XmA0sYKhMMfLiKLpqPbYa3Vqg/NSe4qOXQbLbNsThH
H9ExUEsZg8j5V2uXe9UosrTM2lZeisPXspQkqNkAxIGY9DAiZ+Kr4eLASEOh8luKDZuYQgGX/vHz
+7Xa4h7ZIz1qqJRSMbdPCHbu0H3mbaITzr7w4HKtUDieCCZjGeTf0DwJCMlmKRGzZ0B5p0cQWy1b
4Cg7pBK7d83b1Y72jxcWqjVqxcrPJbmlkBjAzYef1D6/SlIZnZlXu8CvUrwWHRpIREepoxMYx/IE
JyhfqJdvbqMJ+LoywtYxvQt7bnK9VlNd/pa17iQhs8Earn+B0hT9Vz/O1iis6iAWQV2ynEma5S3T
9zvbg7GZW3WKKAtuCVF2el/yyYTj5EeIr0NDC30RW/Igc7bRyVE3udwsgOZ6x9hvBsGyFZP2yrRs
lNgSA1hiPBMZHAP6HjYDAfpKwH1gxOCkQQsU/VejpfRlVPQiC9dE7oDyWxAoukn40eOQQC54aQy9
Rs4vjrHsDaIYqWUiNk5vMot+68Tfl1euM789t99OBoCQElUVKSyN3krukElOO3/xCPLIj9sgncDI
Je7XVDSmm9xAu88h37zMAh2Z2mf/VOaEO/v1P4ZV/Q6T5SNmYGJYgBqYY5BJxkYb+azdno7k9Toh
qWS+WX0vgome9WQXOAWTfjtBW7yRm4+3iJjJgjWQNbnor0RL9+2ibW76sBQWZ+uxN5jHnBNB9Q+Z
P1UN3ejfzz+JA8qzLFJLoFGvAyzFrIXKdqyAzdBkxp1OWBr+CizCrg6c+rpnt4qHRObVTm5Wmssk
3TvUBz4XyJFTA/+0S6cpbTKV7K/30PS1dF0Hm+if3/K9wd07yYIw+9Zpfhp3UJKM/svk37L5SNH8
FmMWlXyUSKM9WmIdSdw+s6uSWX/wpk0AvxhGrNcH5K9mRCOHemPPZVFxAmVckCfPENGb+1yMkjdy
zxeZHCVHp2M32Ig5D0CzpsAhKFmF93w8vPF4QKkX2lrDMqnjDeUuL9lwnftqY1m6B4Nb42eAWyUj
OWmBoh5Nb9OjLRzJI/4e4ZU8AjgdjoK6VKWau5IyqSaaEe0OaUjGBJ5QvFvxcCDUZ2OY9noOqjhK
QKq7KJRy2Szp7u1cTnE2rnuk5UT/Zw3cnj4QHu6v5yj30Zv39ECFqqr+LVibu99BTNagFwmBTWN/
ugvGkQ5FvA4N3yeVFnhgBCMxQxDA3Te4XcKAM2Gv8sB80P/6HNfChr0VVgIZvVnvbB6LtiUln+jQ
DbY9NvtWB/dv+ZO4hXhFVYSWsVX+BUtVSOXT2tb/8J5WCN4H6rRLjC4lTcjivarer8JGozaigFtA
0U1xD9HAYzAIdtxMChwEzczQrKAMnM80jyVaqCzQYqj3vc7bO7Prc2cOlhZ+WCQwbusghR57qtFS
NB2YIAeOeyjrChLh16mQmMmgztlas+Qc2cmyngXNpDGQV6etjNaeDZU3DIrvRca3OPIc5dQXK3W2
TdSPm6emIHzM2y/Btnh9EI8hj+ghbYUz2ttF95YCEKTnxAH79H3tr5ZjMz5G+mqbyM/+cwCXGYv/
cjxWTAfpTDqTR+hAxA3txjREM+ogSBixNRpky3n1lId6v4EK2IGLHcabkJsF9TH10duhCyO2Uyzh
Gj3F/Wyi+/LFAHZN+pU0NlEgJYhbD4ecmwb3HVhzfjLDpW7L0PDFPQ/whoOtaiDhD6vrEvHvZKor
U7u1yoFfYet/StN/QMu/60UIkdwBRcTcvquOb1u1j4kyDqyBKwSMJumlOJR0vmFmYmJ0016wiydy
8nihdsuF62sa+8lWv+t2U14nZMYepIOVwphLJDrq959ZMW52j7+EhdQE5FuiYrQ9iyLuxVLFa3u9
kDVdGEPWIeAIe+dW8GzZscTSxs1t5zvJ/9z+0nfBru40QwfrYP79z7DUtzWWsqWTP9OA3nwLbEJ0
dWNUZCBxQsAg3VlpQZva53rsq4PIsp8wTW/hdfX9s4skf5tBeB2gJIs6keUYZfoq+YhTYnpluRnj
QV95+AkarI9nOqaB4cI/DoG40uXx4N7SV8jOl/bNy7jcWpjg7qG+JsIQHIfdULg+A+/ujzW4xVQ+
WA/fzOiTshFBL+xqIhHutdwqvHFDT5O0E0pGRsKBGFIib61z5/Se+HskHjmHQFuzVAAGlJ01u/MZ
t4kzVWfVNHb7Kwn+Z8s+yh9WVjqxO+IDa8UsPBU+yAmfmYPjiCxaYrPp5lyKmwvoXUnEo8+o9QQK
CtquTFWtYTZo6FsNmsd6IYnI09g2IiMvYuYqAVfLjz7iHbEZgb3KLNOMNE6/O4coWNIcrOLRM4eK
BpS6YlpWnAYBxP8M2wSFdGxj4hy7wvTquGOUwoz5/j/8XngWI0ru5Aj5n5A7NRQCNnhdANsG6S/m
2VJHpwpWcSuvGtdho55vllwYwEN42MtTlMEEvl16oMq4TVQzi2aOuMLGMHGTfgNazPoHAsztb4Z7
4/94mJ+FqbWDaknONQKKMnhO+PJkYcz+6Z6iX9vHY7/Ut+BWwZ7sncTITUH/HXVeuYzrqkISP9EX
wYf3JwBy7JZpAuJIjlUFtl4D0b3X+8/4DYKeW0tgwFCfK8M7ov0yCXOUfrPSftLf7XD2yhDS4MCH
MaPBqXF+zvgUIIfKQXkno3HEAVB42YBomkiSSa8qwFGNlPID5XnoTrNyQG8I8F6buywSbNGda8Cm
fNF/Woeb+aD1vxht6IZ7dRQtt3wH8B8fD+xqYK3D8GOiniFChIT6/8aYyk9ZRk2eevAr5lfKs8ed
iV896ieHy0NsRRduKtOjFWbh3uZd8jnHZ3QrCaWWiUEeDvfX4zbTFStt0ovuCOwEhMaPbo9xgKSM
Mc6wDkHlyJ+YrIqgJQDHcai8dgI44Avm/8v0jZXByl56LceCPh/CbA258fHvuFK+BFTSWMN97YQm
OHq7koiGFLfwaNuA+6AaxsUPnkHaPeO7IH+PmwoPd3jUN+kuWXeK5ABhiIZPtE3wErZBQuKf3VyP
fLRzxNSiNo47tdxVL7+V9KTGoDUa7C+42k0vIxXj87i9JDbgo4W1wLZti9HeoygM+Ug4WxnmIWgo
YtueCvynQ2IWBFigMHX9qRVuhKnvWHGMKWHMrKmUisRNbDpJXYgDpIQzZCJXbKlqgyg9Whrzwugd
9wcfUIKRSQqb+l4hoCPgpra28tdXcPxKgWkuzVKMUwRYmZMkEKtmYzbZmg4cfpPzf5cgSOxgeLdt
b1c88NXSmvDT2VVZ7G4ezPhC9lFgatHYBl+0BZsKkg3bYytmK7f0SYX07CuIolp6yLCzMRIhg/oj
033NQc/jnEldXy/ipFOLL5aEuG+/YkK/m3BJ5Kpf8sTsyDhn8YiAVqgLIFV6sQ35sZ5GYbB+pd8y
NTM74T/Tr4MJAbjFUtU8ceeGZbbVVWnGPsJ0m5nfpGFFQAUDMr0kuEA8AAptKr3/T1UaaIRyzBNl
ZxiOiEMv3/J6KzsJETnfvbc+dKlf8nah8jKF+opNgz4HbKStEKuwdCGCmoe/XqwFpQfe/SXmSQZj
fCqRtDwaqXKz0dPBkQ8e4x/NILC3+UufvBa8YzibjcJnOTNhzOuFg6zZf/6xEe4VqGagV8tkt3KB
vKiIEesYEx4uUaLMlmCF0l3jeHyNzC4vzw7ecuF21FJNa86Rdet2HkEcYdibHd6NdALSi/mc6fhy
gyGetooXn64d20Bbq6umZe49nNS6RubW7hdqWQxjbphmXKGQJSuZLHJZkZkHU2jtrwj4ogQkDTSN
6LIsh4F5pzwdECSW2OdueA825iPaPl4D7xdSCV+664tr4yxM3TOXIVI3+ejGcVOvFSLQcG59Kb3U
xny/2eSOF9jxvdqHbjttyh65FIJgJeIbBfbVpYDRsXvdjs4KzgmLRRCq9RdOU1bj3mU0ca+3VCzP
6ibs8ds4EIksikQUBHZuAY2WqEnC1gN+4dHlQ/v8IWfWkzQKqrfVYh3yzuNTtCvl+rWmzrkpZMKW
zq+oGRJnukLdHENudi6llxAyAMCDv8KyTMyl+R1dQDBelD6wDN8Xq2nDwcZ3mcb1O80erhC3x9Ex
2/5Y21qqe4g27MDcvH3ftemzMYuvSck1dglrSCuogdc6WYtdosQ9cxaALWhfysr07nqoksOUVoL/
aCFL9WztCx5C0vtuATk+jhpwRTM/dC27RRglftR6GV2uCJ21by8i30UFgQq0LwjTREgPWlUiFDwi
JOFKVhGbFHfRHyOlqbnpED6HVUgWLuIcA0ms5uKJTkajA5wDM7+ul/8MJUr6m2GAoCyCeMssUjXx
rCP5ARhXFkkbD/lQrFzO3sQF/oi7xstwIUz0g8DeKd/cQI9T0LrZ33fiiuf8HujjbzbPZCwDavBE
EDftiGdjLN9NSrc9IR/7aa9G4CywWYAU8WfHUm1ppAjl/Nj39VPZc+kZdWh7gZan1UxVYB/nOTqJ
ZqKgRKKmj/qV6Xhga2BgekCPqS8bjjBKk/hajmhZPNlB4GCtfN+FFlZEZdnH4ebGX4bul/ApsuVh
Qm6/DflOvMFHN6XOkNviKb0h7ow71dozqAjo45DN2gTCU+L8LdT21VoxyFxfaQe2TEOGb0/C52lh
1F7AWYAhzly3yUfFvSrsdL5A9iXsHOYMpkTROXYwbt9FJJtgqok71fkP8S4ug1ooHesonu3GoxuV
BKMCPq5FDyhT6R3Hup82o8aeS5E1gbtM+fJS8BLWgxcgf7pXqo0sC7rxORVBAmd5Yix/sHUFwr0j
BlthKJLT1LleIKVGWxIfSLKqE7FcTkILt9NwH2FANfy1+lEXaf4WRix80ptH/TVh65IV31wIh+zu
TBtJ64MVEqHdbmaK48l6ROKTNeIUSZs/H1jr+9eFuGeO1VroMwYDg3S3NDpCJmQHL77a4ehuTN/h
qOiBYRdANvuBMI3K6ZdIESyXBZMTqdhYvw9QzpUkzqMk94so4eEhJyHyzkgPNmVfHR/vG+dK40Ig
A8Kti4Bj9Yi9aTEDJZ2PiI4hEGwTamLbIB+b/6z4ltDL4q4XtQ0bBY35fjYHTdIc3JfKB9mTwQBH
uZKxwYfWLQKxiAp97VtvI73SNHsZDTZRtuSf5AnvJx1h/uY0swz/3nWSuIksAqwe2rUi4GetyspL
J8WO0pA8H9zmmqIJXRa7Tye0ZOiE3XdF8T2witZXjbTRow6VkpOfHM4sIveLhpzkKVsZLYkZu+pv
lGVLVMOMOLfjM98hRbOOgJVb3dKUDWvYPaXB4bLYBHY6B5A8ia8rK/HToeXS35Z534RfDyH9/P4I
yqmtcwWwYI+yZFdiADRQs+BUi5BaSlhFZMp2FqGHLheFGmMZzrm+TMsbt/ohiddQppctmm95qhqB
JPcCY1xJkiaLZv15gf9FOQ60KtoPnOkHFwve5l43pWOpG8anBjYxQZb5ue05fF4PAnGdMlhrHN6n
YFPcZeIQXcpEdCaBxmQQt3LECYnsGA64QoWHBxrG/IMk2LXL1TVqbLON3agtyGhvTYCXWEXxp0lt
KCQIducYf3N49CVDZoF4UJ6DipZHdDdj9IcoiY8tvw6wlxDVSu+JQMT9bttY1s48NcM5e1116VkX
TKU5c57gHT7DKso4rz1IoIQGW8nkgFnCcwAWQA/biJ02u2sj6WuTV6YNMHDl69/xQrQSgDT24QCH
PTb2Fql/4PW5UOoQxTfVmo2lfWWC7onvxKzMfjCBqIJivwG+uHC+n5um+FTLHCUqteI6HrdfCwzk
NfZmIV0s0zus8nlZWg7Kt0rGd7fVIQH2ANXAV273a0cC7kosvnw5vvIjIPQmIT5BiX95as5xGubt
nmlYKfCK4RguA63KimbVBpbR5rPxag3tUULb7OvPoRPHMr8diWeazFIkhwxWXM9sYYoD2W1MNosU
aaPS4OervQXRZ2PqKBgNXgtWJ3Q/b93EIKUFEPJ77vMMFB4utzlv9knFsjPqWlS2M0np47Exem+D
5HWSYlJ1K0QXOljIQSEDpRvGOfE79v8vK3Ud4vPdL+CVUgPTxp/eQz12W+VAH6Y44hz1wmZuvDYN
j1B9aKVh/QDjwll0VaQb+mbv767fD6K8u4lbyNcwsy07qYiu4Y0kU7rDwSvMYrVIEExMbX2t0UJM
MKL5Rnoi2YpbED0ktHx7QGeVDVk7s9RrvgO7qflqdR8eOd9G1YhGo8Xwmcg+7jT56Drq9BimFpbV
mx3na2uaTYD36cWKJrtO0kZwgeYOnAzwZJNBWyTfcbDJFHoRiWxenjQNWNKUl3pxi3r6kecQJEx2
IVXB7sPeMulwcE+UzTxmHEEHkeEoEx8OdLb53sAqByF2vfGLK3i0nlkoRBHnXQjgQuiSjGMT3Wy2
8e+iSas1Iby4cFd+xhdUqr4JGJT2d6r71eTlaV3zp5Eon+UVMgH4yHjsnlaPN/Bt+vTofF8xYWSg
r5GPLfI9SUM91OUArMcoAQ2Vs+gD20BlJF+0/V7cU6p6gpibZY1iYS5M2sBoTDE++M/hNVqwbS2z
5iuN288r1G8yK1etMzHoBC0Lr/ebqocQrTlXLEt7HPwk5spXM1d9Krs6feQGaaXA/f6TsI+s9pFF
Ncph91V/HAfAGBn5OJ72B48ybQHAvcj/fRGV/Z69ZTrPIicKdcrXkA/JAAATsvwuki7bk+EKzjUW
cMpuXMjFNOoNj16OcTVqQoEgJI5FssrZPsGgutNWJjofaa3h427sUU56/6atRLELG/PTD5dR3pmx
YjUXvdIspNkw7eoG3JKPnCDmPSKfDV1liXvbCefRS0aSRvfEp4ydOLInLybeDYEiAzZfB235S1J8
SNjsbWT/ecjXJnktHo9AayvELvD4MPWO7QzPw7omFza6UdUC0ocbKAyGYTm0h3f+euLWt+lr9v6C
E+4R77Igx2f4SBEz1H25IIWphrWOVXYEx2E11/a8R8C4xKOCH1wn17a1te25mDyOliDHODhQMgtr
wRrF5HpENn1H9LI9QTNC5knIizMM63kXaN7Ckyry4BRh1keiZusNrZ71g3FJik5QFdCNtL60Wo1T
5SJP3WEvqcFJHO5fmbXc+6gCDGg0Bd3tqba7EhgplbMXwZRYwYGIx1zaP+lqvsVtH3Ne8lv3pfJ9
3ieUZreZvk1VppSbzADPCKvEL/Xz7Cb3HzkY9DLwGFA7eGOs28VfGZIIyJNhnqefiDSlSoUIJgPA
K8+Oq1nfohvXTOFMcMoOq1wAm1Y9EVD64UjQTSfeU9s+EHlT9dihKuSQGMqKUtprBVsTHL3rdCsr
92fP+defASHAb2DqZ4ZKIMTlx4lRCKHdMkYFO+v0LY8cXKIDl/9Puc3Z2P1nV8xLdRjdm/uegaL8
sBpaN3H68lBqoxqRjWHPr0lCmuCUr57U/dsKm+lQDHF6hskg4LvPt9G8kDTWTvDU3GTYh5c9gukR
gM6H9ZCXC764/SXvjt1HPlFcPm/IXowJEk1lzM+AZPOh3Fl88U4/nMD7tAg3mKeiFkPdmGImPG8e
ePToRm7oGf5O0BpR1UPZuH/Qg4xIaaxRMPBuXxwtXCkRcVD5t925Gx9+nw4zU5XpMryMbC59tREu
guVIf+diwUcsMYbvL8b0SItHmXTP0t+zqOu5WUax1O0VGsHeok2Y6vjluSq+7jtqStXnMTCrhPVb
FiEoBrzVpru5SNpBZYOeFI4IB8RL8RhfdXJ2lAa/cQXcUOVHuIN+fL2FjFP9rJprITl9cuikiZs+
Gjp62s/jcTKqpKbzHnrNKphq80buIoyMIguAvCtMbEZm4Y8o0U5l71gC6OPgxU2i1GSEFrYmIGAt
YtCH3rV1KBe+zkiEPC+6S+DVcMz/dCLlMoYa22yiAfuXq4FCFKrLZBmCuA2D85Pjy6d0uQ5zliwI
1WxdRB++a8vk5yM5IstQqa4al4kB54xt+tAiEZx0n7551j0jt1stM/U/E0MB/wHTFdem2Xb67aT2
9c0zZ8z0gUDj1PB6sMVi1O1nuZHKqKXEm2GD/vsKkbcE03apR4W0ih/X7dfFzOn7ayC3x0ZSBxol
vPTM1fmG6U/D3IfVwRuNjULYuDodLbV/X/W/232eJJlypS+05d7uzWC7yyaTcKA5P4eYyUiAOf5L
m8ZRNF4NRaYJwfW1Jd2WMiknj8RO6/K+L80QFl/6elGfviX/2QYmFEnYbe1mxn3Fp3YL+1Wi8M0A
DnzhqFQ+rsmEaOPBlSQ7K56DQgHh80UGmQsgVGkeFnHCk3OojphKuDLzqhh5rj6XVVXRPC56fh63
rtaPIc7qkuOFJyL2P6ox1VtqUD4ewpzFWX5h/yzR96z5CsTgMCUNARH7WCzhrhVSmDU0q4UN+8L9
swSXGYak7RbM3eAOmTr26c3f1zFNPY+q6zy0H3rs17ntWBsxakuiNU6WHAdhpincDbOHPmagf6zl
nnAk5rTj87ftJt+TPwpFXyKP0dLyknDAO6pnfC1LiFWA0epv9Ou3w9r0INJpiMdStJj9wqWFxdVQ
gpx4S4VZM+NrxFMDCmhCHhhJGj/Cy1iTkYyRubP+f5umyxFYLu8IMNhMa8L41XFGZkYEn/Pszmla
6fgQKVfytv3Yz12QTgFYNz+cL/It6wetaq1Ndnji3WV6x9+C0Jpe1fI20nq0H1Za/kIDF5Ddo0T4
6SGFKxyIqjzXs7rL9EuD5I3f79yu2qkad6zue+crOmoRoMmFYdYWs9Aap1UWar4JN4ifaphB2mmQ
gTceECMmLX8ZDLqUoLzjJJ21g0dUwD1uANNeIfYP0GtxOCOXJ+RopNuiFtisQc9h1wjD6NcCynPK
+3u/fM6trW6A/cQ78NZkGcjcV1D0lFxNCWP8Ymll09hMzn4m/eiGVd+GgcWC03bSfoyhq2q3pbdl
yCmxegx04j39hs6vA8oSkaKqgRFECfscby3tWlLrdsQBBHGC8AIbTrlemIbg9IiQyNQDRsGH5OQo
tU4Q5dqz9psw/rXeyxSIw982z1BotdlCwVaE8gLOJSx1EYvcw2cUWpq0uwY4VboiRNU04dlgnZJ0
B4WwDDypkZgk4U09KTyQHhZHS9Xc1FnVTn6iNfnu7Hu4Ft8UUhYrPq6vM1cbNLke+gL1tlkJckWa
pyYX4vdDBo2njITbEHpoLn0q7I8r4yuaQ9ICk2GuKbu2Y4ZHEb1yIqtjNPqq6H4fst9MhiROS+2S
SezaAm/vjOMiFOmb3D5M2y2roJUdV4GZQmudDQz4ZMAztevFXnPMFmKs+sJV3uP6zMWsFRxUvPIn
1OVNnb+XoCMysO+fbZab9hD1eLsMsL8HY0e16OPAxxILjStOlAsTbU3mSjLbWvJ+jDp+adGAI8Nq
S+LeOSt+qDsq1PibIFk4x+mhi+vzKnUMPxP3RHxAwqtwHeJeX0FlTfzWO+JlXqRrRCkNXx5KL1Oe
k31n3mgFLKRDsUiqkAIthtemqvGUl3jqMigxk25WX59KNgwV4A6H8KbG+rb5O2WLiaWTHIj3GvEA
A14nkYMZRr4pdejdPZyiObHvFccoU7Fh6Ku19Zsaal0jjaJo5TK7yDcplJ3usI9T04/5hMVoiPhH
oQixKuG9HgPNWQYd6J/TkHwB54uuZNQKCtOCGJn3gfnzFV4uYGryto62djFbJlXqefeLznTBrMqA
l5d9m6niNVRUmMmwGJpgyn9I3PmoRGIIHaHnKNQMXjtdCwbnZAwyp8CTADP+fChMS7Tw90fDzeRL
hbv6DTxvReIZ17potw19/hkQGDbJFaNZWpoasBpkFGg3UbLts7goR/ynldHNvQKCD7VZPLSb3bQS
AeAT4CaE/83OxHEDU/oF7X94KzyjCPRl8NCMUuPvkBbe944PqPKXeLMGC9b9SgiTNLKp4loJHOUX
jglwMF9srKopHP+2m80Rifaat3PO1dpBBy6vGVyK1jU16iM/x4LSQKjnzjkS8QY7xg5ICbA/9EZg
Mh+0OiKyn0+A4UAbNZkDvpqx/Qe5cpvpWlb+gOAo2ITP2BLz3qncJnARBL3nl90DY/ckgA4C8z4y
0AoTpP+Unpa7fqymTn2s7Uh9Y4GHhEU+YbqjMVV0W8aIbTHbtzmmhtx/1ONtFF+gimrQJNDz38ST
CzkK/B5KdHa4Pp6p9ufLT7pZiRwjUffPYHEwh207ksJ0pjapeCJ5qa51t4mGwxE320Gd3X7ZBfRE
1Trek8D6vdKB9H2hewQbS62qQbQ2/pGUjXN3wvbKLg+UDdfLeGb+SlniYYNGbWJBabMbm3jj47od
w+om2m8J5qw6LETIFyt0VKtFXh3FYuNi9X2PLuo94pUyckOev0BJe0h4mMD+aizydReG4Mbd7Zdq
JN3KtWaxHNTg4Fwi/BK2DCsUwr0Ifh+sx9TxOUIAVzhIyXpgSmA4JObv+YRb0RP4g4OSaXfL3+9s
50ia4kte7RJBMB1D7bqmNEqjAHcZEvBJJC93xRTBwCVnQjSfZXvvZ+Z6djbGNNszyp/qElPGjZqX
3/fP2YeL9ZBBjhzQxJAnjbL2bdHeMRmGO96ILtEh5pOMq6HpK5Ut+wzgVfszAS4XDL4JqPdjndui
mrAc00q+rmyyBPcEzT2sQeYmQV7TerVGX2yv6aDbixET3vV5Eqv1Ml2OGI+24Bz6RdRFl4MNyuls
PHlJozpj92gzL8SM6Qrbcg6NQGjuhkKxFqJ/xU58SQJWYLeormSIvAcb5hC/iCTlhwq+8zymm/wg
hk0h3TM7lYxp6nce8svrfeoj6ZiI5MEAxV2fU/0a00CVr7VIbxUlphRrVJ9A2XCFzoz/rG9LvhoM
qqeFOWdiQSBe1GVZij4CohOJsCQMpU8vM6ao+Izq1Uk3AVXP7GpR93GRaFZRu06HHW74476OrHcE
k9Mi13udc2rE00q/HVKep9t3x6bn7IyUB7pw4FsS5UyliA7Udw0JQVJG0FVxNKkEhSqbpBE2lDjw
LeawN1YDlTkS3JT2AVpH9jiwcgAg9PZs4PcV+uYjq2FLTn6s4nuetlifIVtEBSV+aRnPnjCbVs5O
oYb2l1wsdGGvByLg+OdsG1omzxzbZnFh1965IMgzgIkkbVHThVeU1Onb6kNEWck1hE7u8wKGK84n
KwpApHFAgNS9f3XGc/XJul3eVohEgLpGNcUi0hiZJSKjsOQgbzO8HGIhcI8xN6pws58wCLCWgLKc
JZnEhUv6yeHBq3OYyT1F9pei/typeZLX1TPt2Y0kGvkUQzMJ83bz8zrpuoh/beVe9m+ehGqpBuMU
B0THE2uoYkcfl3i2LKHBV9fCVmUDGgMZPoqb7U5l8PT7xD4OV6097CvVCMiYXDa/N4sGkAa3Ml3V
pAZYPleoC7u29LphNx/kl8c4gU+/8Ojv9vItNcWB7yHYpThYcU5WgVxX7ulpdeIDflWcHSITUeI4
dWMz89hcCTl4Vp6MT4FomB4SvWZPGguud3oUM0vL0SWKZmF0oKZyJCRMbkVsbckJsLFB/wnXP6g9
FiwQBajLGqYH7gmdVTfPHAsXqeri5pP4RAR6JsvGwCiidatF/hs6Bi9D/4pLVy2MB/1S8qamRG4y
9feFxwAEThIc7AOvzTwjHT//jdIu3QM+fjyAUU3jcql1JadVM3Y7tvE4/6HRyVv/wwFGjlSmpunZ
3VgA7TNBvPnGV/50PuH2+NBF7oBVccr/pkRt89c8AwvWYyQVyUJPxhnbbv/OY1OnsgCkKTQj/ikt
c/J64jBMXaPYwXROY+FVuqP2OaekPZF2OT4jjbeNbNybXZAeMvJMZp7DGRpCOq0UBnGglAyMhNTf
jRumNm5nJGGZZf9F5K12e3Po7ns0+VyrVk337sQQj9scZqd6KeD61NOUSF0ME88pQ6s2c+fszqOf
zaivdaqvXmvatwte6wyRNsM7YZ4gFz4rweFOjG4qpfDpq9O087PEfLIxFvonJnc0pgxUAp/qefPf
gsxvPGY9AqYr5He0/vox9O5+JfvLEKPxgh0Khxql0ZvAQb1uMcJnOeCYKsJJw/1TNgQZl3zsQ9l3
B36r0266rZJC8ODnVo3ESKIEEEgrH+52WNl9QYbGa10qVk8qQAh3tNAEBskybtNKI7XCEubstl73
73Wv/2fqNAtXfZi1wwv8GTFTvquLYJKfNqdiiEmfeakkMJkaPnnuUNp7ZKTnq0L9H1c05xHZUX27
fk3K+CR1pKJRQjKE9L+h3GOqq4X2qBrFoYOoaBUzh7/aovxWB6tfJYBW7TyunX5RX60UvAXMUFGx
2BgAbmkXaNWOdEiBw/q/rNFXbGiv6usa3o2KXA1qEQeCKaRpT/0XHKCDbNQhMnhS+UMmh1argsVJ
V7aXmq2ThP9Smwtey1pcWovmF19dk9jcp5y4XZe/PYN1KJBbWeKcU3qCGaF/E7zceFtqo9G79v7Q
fPyWB8tuxEsoN+Tm18ulOIxb6O98NEPQrid1PAoIPgvbiUr95/zDx7CdAam704g/zvfbm3NKA+Vr
GdVj/xCyQ+eI0JNYsCeFwAo9MlM11rcrqgJfVWYOFOHs1+fFwIL4jMQ34EiC+GDnasgmWSlwsmHS
u5Du9Llgcc2LFAXryM6LaZbgxaIIBe1d8d8ScpP5OATkxuiA7j+ogWUL0S9V32kRtQAWr5Y9JtJv
q93yMqcgsxKpM3kdREnrHAPXCVuav2GHORvgqYCC3MZ8fbsrj6nRCZ+hLkUn1zAKZUs28y7jc6/6
4O496XlU7/I3khSuKNYnU+z2u68iV3V540tIq3Aj3pzHPz9bIYFJ91rG8cuh018LEYg5k6BY1FwC
rPsognWXhqHP9NYdz6/8iokvi4Vba4KiSRO+pMJr82rSIjaCbTwo1yaBmPdjGOqJ5QnqH5BwY7hI
J5h3ihnXiCibFl+4VU4SqisdaKjYlDIv7feRzppPuRIhAy/sKESC6MzNl7lAGdEMu6iFceAJ3U7b
kzKWeZkHP6Wa4F2MRO3LezXIM/UlJ8xvxGsLNo6u7ke4Aw8fjRmSmI4jkJYX4Wx9yWE39QPyXA6w
r8uWQN9Y0Y41tsmgTyGT+sGn+s5ugbQ1iefjsSQJMC9kwlMmeHJvNnM1K2RuxCHWDzE3d7Rn8jbj
sNi1HxJZM9K/us9Xx2asXMVzEd49OHKN+rORoBXS+PbrsfZXcAUvuZN01ZdUGn+dsX4ae5nEW3uj
Rk1PQf72/Y9tcVG4tVmkGLkWVxsWrmuV0TISqjDWRHnI7DCpxgfcuXU1hLJEDs+F+SkrYFdnyVeT
OL9BMCHdHp5K/EQ2WFvDCJ3PVkNW3MtUI2ZWF6/6rrlBrztTfit6HlukM3ECcurTyaJxFE1O1xNB
KFDHhcHDJmwIu2CJgl7cxlY2eczJAkccZQThyogEMK65NxV8YC0wczCO1CEn+Zn5eALnowNEYd9t
OWZs32WB81VuZrFqUJ+F6+R9+zcgwgQzYSynTCkcg9lMETNgZhwpcutm9fRMJqPX/br14ICwRMfP
4GJ1Iuj+43UCOlXSSSGyfExu7Hqt1mgx2qHbdGGoyr9oKerKDM2xi2VzbJR90uOo7+Ao3mzEl5wm
F53eKSafoBnkWP/cAxxjNAyiE808e17YBx01Tsn06Vs62Q8NeackZ5y4KMsk6Mi1ikt8QPcddEa3
kS+Hubr8UP27UaWI0W7S7Ni4k7w6Xo5ZBhvyA69r1DordQnUkrgLvOpRKXTXQJaO0DcuBRXoYvMC
vJsiVAraLBgq0GEULty+PoDkGVC/O6frcxN509IpXy9Ko8z2nQpQMCo9MAmRSmNh4ZOBL06ze9JB
fOxBuLTLKaiQ4UDmqtNzaePfQrk5yp0SQYdnnKq5KhFUE3Fw1qDY5sW4S8jDVfDOGSfpk4ViPa6x
cyy5p82WQz/Vp6yNX1yfZXXsuNWSXTHR0E0PqNbu/FC1VEqeDmd/DtN6nJRPN6qcGr3o2QcSK1zW
LFN04w4dcwk5CzYg43RFdBC5Y6pjRBTkQ+1lYE04bwHogfYeHXI4Tz2lbjbqyouSU0MKsmGllnYZ
2bDIRTMq+mdcILLWQkHVHEkIH4BpdeiuxNZIaVPPe8gSg6QDmfmZ6JC58HWOE5YXAOMyLrSNNxpH
iQcvkGPzu5o9YWtXp3VvObwrP+T1q++xvHL3SaRByqSdJRvH7GB5kgfNPHR0QePZGJCqevxAEChy
H9hLTZyCAH8MM/stGpSfpeinZxUGipEVoHV1syJCj8oPQ3/P9NOKwSSoyVUeWS1ksotZ7tTEaRt7
tnREDh0zeeAwLZRM1JlFkAL6EIDndEMHXeI50CswCtJl4GJb+xqnry5V2+rBu4zYrHJUW4b/oI95
XyFUyUxXcTjUIwaOnYJ0NHMI1GDdj1NgFG+kDZArHirJEszl1k5OerXD5lsUqIQtQ4ZhDmTmJyJ+
4bMKDlw+M/+LiN2CA+kV+x8VDTJanfaFXPjKeeSUmFKbAm/2FTMPD0Pclw2ZA831ueD+bhi1Odld
xrDRiKUsMfK17RfyB+4BGOfejwyQPUaIrTTGKSRp7EpEdCiMx6rVE7sos9tF3NoPZy0PfE4QD+sl
dh/EchRv0wXUe0kcA9hBsAdajfJkvenOyyetxotaNGqoKKENGPPAnRKEAxR54QLizmP9iRJZkGlr
1fEd9gC3zWyMHa5lz5JcNZMf6NqTcNi/WaGm3HCuBfc/ylZt51Wakol5CEr4i03j1BSkYkVFalw3
9NcqKsKg1BG9NmyLlfuDaRYPVsQlhouZ/06wiqDcd3eh1EcXImkygPVT1sWS2fFTMIAaYj2TIKdk
YQoIxe026Kjap+xAZkjoCojAOOm6s8fOIrotfRgNt/3KJUaLQi4PXNAvCobDvpsP+XRaBpDl+0lq
mmkNZwT8HCWpPjsEWTt7OlMGdN+3rUTxgbRf0I27+fJUY0oBEd2QMleiZR/RykPQ26dZl8G6ggVc
NvEL22XObNNI41Htn2jT0nZjCXun/YVAhG2xcWxIFtdH/R1TJh8/dDq64+2JQNXADRZqNSVo9AHp
YVEsVMy7bCWqbpCdEJE3RJ42bSA30/W3gAbGPi37OeZREufrCoHzeNATvsi0jJKZujjAc8CIBbUX
l0Y02I2Vb4EY3a9v15z1sDX0/yHKPmqp9/YuWP+YjjP+TxUJr/buhrujult3mUNw1U95R2TnGR7I
Z/h2LvVStpiwhtV+TbPAJEB+hm1dj/WzHJQg+GNwvByc/c8yfd1lXxYgTR7nnHzc07XCA9pOj2Vg
9z40ZVSdo44btTEqlTyBOUiquy5dpLhjzcckTjK7QJjieh0NnfsQ2R55ejeTlkHgSn1JNL+gbf8S
LeM1Xjf64jcQMTGxHpTmsMYUEdQphtQ4VG/6duejYS4/jimGkZx8ZWVt2uXEIFq5RqqzxGID9E3Z
hXSMjAA2QN5WiC9aS/p6xaizNYFUhwfkXLMrsO73p/cCdNuoz7xaeIP9OEnVrdvhZeiMKtYJUy1r
56PQTXGWtxoO69/7JAS22Sb4QZpf7NVaWwVYyo5QocIjarMH6/WUu9Nv/qah78LVf/EqDea8DcrW
J+1OXksdCIrSfn5GHccMcPSF9O4t7FBgWIM2dqYlTP5ifWMAkLbBzPCOMTdBKS6N+iFeTpOEyj05
ZBRPwBsNKjKQWdnt/YNvgKLTgAWWKquabwd3i99pVepR2fjp+27LPi612C0QbnzceTWGyHAb5tJD
Sxqyo1WWVpbtf9/WmU24XZqNwT19Do6/nVOs/I90w1wscyhIiM7qlch5+VZVODGcM6Oe6Ck6Fb+C
8OqVE+bd9Tkte6BPzjiv5pfTOrAg/AH6CwoHahTZ6z6SYFzvQSRs3DP36399KRlNBwT/o9jAm9/C
BcPbeltXtV6JfURdfgNOS8gm35geuajAJoi+RvUFYKdB8GbAawC+hY9JImYcGzptQbv+v1+UAjA6
2n/rP1DPEqhM5h7wpJWAEfXENDTyo0fTr21t7tq2hfxTlyb7bJ/ZTlK6OPQum7wz92wWaxvqZFPQ
1a8XnoYVEE4+DdNB07lyqkpaOta62mb6iKt3Vlg6dd9A4CSs82VFLAB44fsbDZDVw/IiudPKhMKq
1K0QvbXwP0dUk7Uw4iujG8M9hQa3yhDkBweKxnGSGXRWaeqFuAYoqp4e2Kcyai5qJPCkqJzQN1aQ
KZoKDMKS55kfc7id6sFmAgRfWB/Wbmd1BsEy/kzJ510ow3AqQIb1ad4P9SVql2VdwLotcHcOPUvF
iGNRoomO3zrL6ZHJjOSL7w0+IpXft8liffU5KAvpc1x/tDqDQctAkj/d+jxipIpwxpBm+MRdSovX
KL5HWFyYtzYcueWCugJshLKcA3QA2Kcbmp2EjAIvjR329s1bk9aVqbSMNxXdYSUUdUh74HJ9WeAw
J9Ol3h2nT2nutKSGaLRvZpQ1FtIwJf4HxTTHM+i0DAAoLv6UZ+mX9OOI0OoPdRGZxFM/muGA9aTH
JS7o+TgW46xzARCiw7i0/JSU5O/LSpj7xWzpRAIOgDAJsNNU+Q5q/c8VtipPRTBxZORjQoiibCoU
jNmdP9Hh31sfJMN1jyxMyQE8vRMdoK5xF2HBwyLJksgIpaKc/InMaYJvSD/2ikb3NS9Xp3+l6tJm
foQ3MhepFKH8JOYs48Aa81ID+76S1gE7mQQy6NyP0LrUwpPnOZodh27i9nzWKTpu7wAJe8JDNK8Q
FBnF/pPg2spW4u1WAArY/jl+XhizX00itJdRKHZiADubpAiwBHmDfmw34tjr7vdp+i4v/wm6Yk54
Cm4Z7gK9fL8LrW0SJ3iaRFVcINwaxM1CoNaztlCuoF1Inc5A4STWR8oMqG+s4Lq8tsAdgeNGD7VE
ipg0W52jMlGeSYF0OdHc7gfQ+8L2dJFyNVfNNYMHJO9RSSACEJKdxz/qox2DEq3FzsPkdLfH7e2b
9n8z99RJiEJEan1xHzCZy7vnh5xVqg3n0n0Uv/IXmgiyQn4ba9j4MS25y+G2I58I74VZhm+BjQX4
YfgoJJhEKfkiv0q9BafYtylVcxazbGRJMJbhtovTBeaAvVLZ+IvgdSu0vW3ElVw9i7uzNgHDLiIr
4emK/q+sR4H6WwVgC/JdYhJsnW6VBTdqfTL1EZLXQK7OD1p2weZHyB1TlGNh4zT7gWrdLWelh7zo
rq3FHlKN4+CqqtIYX50VJIYde5X6Pk/diby+fyDe5BuBA9syZQPJqzTIt5sXS0vsxhZbnPyRamEH
5if1TPo4c8RHfhQh/3G4K2PePEbfYLvLITJtqu/nXZTwpcrNYBqx3qJ8zhhO4kyHsM9cXU8vLT/T
+wZyK3ZsQ2zSyRuAi2RuvhFXvVAlxtt4YEx0/TdfUjtZmS88q+m2NVTw3CaTHA4cio6QwKMV87oB
cW8YuWoBSDi7+L3OHZRo2N2CmeFgHdkl3KeJ8FyvgUECeQ5WGM5YyCJabU05f3LvgP6wMsM+nYAZ
BjzoOa+TGjGnX5Zr2822CQq4k6p+w1nH7KULiEV2xF1Ni6gzguaXsftlZBnfxcU74Fb8+EnJ1HsU
sXS8LmFxWCoEP6+p/JzlaXisWEwlbGn5ytUyYpots8YbbI56YBQBUOT+iaLgZjY0YrWsWKdOm2Fq
zw9QxHAiEz+WMaZMZUOJHxUgzA7yXt1ES8cq/hKF31Xbvc2CsnHgwkmfI2U/YpoRYRunhhfdk+Hh
oNkD1S+B6slsBCxSMKiU0AqGjcWHjAZg+InSVP5F0Fbock4J4wEGk0BOZqkXAFgFeA4mOUqL2aHT
q/hea/hkcVrTnzg/+FURaNfkWVtmhi9h28beoaDnzANvNpQXvy/CC4JKmFdMz+t+TaDNgCg9SxCJ
s500eormcImUD+eEsNA1CJCjfB474zy6DYDr3yJIkldMd3qcD2RonvG4kL1yMUMQVW9S8g7UtOpR
0JyYOnOyV4r9iUG5WPMWKM5JasK9KAnufV1Vk9P1m1o58NdvwLpmL5Pok2aKspw2aedRINicOv/K
CHF8W8H3xHWeq/xqZagtbSocfq6NKB8DQblktoRpZatxeyEMnVlVtXi0wjFFAJyJdlyW9CfhKBNh
5nkO1zZDeSeHFOm/SBnQV9TeadO13wUFcYatsiW4gKLwYRtxa12NJTODYgiOvBTUci/Y0RbBosYx
nIG/35Oing13xxApYD99StAsYubO1dckLbQRfmCQYVJuiODyi25YiaMCP8/QUt42nzOLUrTi5xa1
voAWYq3gXIxMy5h88QEK7fdktKhOBocFbrJYnbfi5pOKMQfoDP3YiByXUc6fOodWwVii3tWfB6iD
wolqhU4EBbvrCfpoKwTkcpthDKKbxW+T8A6D7Q8synVSAvuhjwUszIr+XtW1IIhiUp+H/YVsbyoI
uZkt0s16Db/Kih7ho3EPiX8s2RWHPuuV2kzeq5kBsmijlCMTwoPvQG3suEI/Z2LGt/upzEKWwbXo
l5xoPlfzqMTZrpCJHVWI1mI842Al/4SShAIqNb3EG/FoxEDbc6uLo5rDP3LVzp+AyGg5p7USxH8h
sMbOSlpucV9p37UlKsU9xGYFVB8VxewOEqXTqTdrl4++dH+/pKjThnGBSECjzuEAOlzk3Ux1dhT5
Qj4F0yuwbVjBP6Phps+WNBWuvfDHdu71KGJJpOJGygxvaso94YJTfMjq0qpkfUknUydc0GNcx99M
Yvr0/nPVR6HAwX3EGnL4i59dyp+8W6zaqjYeaKAhxlX3jzCPV3+AY1lW1shWJYelFRhxpXpfHkoG
dTk5XV8irX3DXVPmw9OfqLpfeLiQkx6fB5Y8/tkbPYCNoW8zBF+DBbaAhksT5ksspE+TtbC/euzJ
h8jIlXxXsqTdya//oGRGZ7kQ0HzQnKD8cFGDYteQ6nIjdcHoulrkSAZ7Jubb5cUuTO2wM0xe4Y6F
5EdwtGZUvGJ3e5gIV3qM65AlMFrx2Yvx8nkJh5fEaXUizulyLYkohuTZWIQ8rONebmq3YUmasCuH
ekEs1q8RAopd+btk1H6Jv+VK3s3Wz19pOwvG7euS5vjBmJJ5SpTX6HDs/pnSPx/TSKOI9WtE+WcQ
w9A/fbS91OZ/kw7N7XNMrSttfZMiqdoCDEykvENS/Me/3SeDjYRVFjyX3cL35LgcBSkLN1F+J58w
tmeIPopob1T/aABTixR+GLMWcJo4/Ag3spqwWLXLRUkJljqQVOoWQHhSpHPrqIk9ezFjZJAotdSz
ffNbfYDsiRPeZqNJLsdHBen8Eqz5H9QTuNePQvs7HdpsjZZlAZdHvgjCAZR0WVn2IwlsFpO6buPy
6OBTjjg/IVaXvMsX+tPiy0Pw9PBK26ESwk8bWp//asDshMwjnTjAqn8yKAbsMkEgLZHhur3GKO2N
SA6zrZG5PA9pLvCCqcpYn9PpZuompX+iLR1OpNdjz/RKKw+3xMclce3tFZxn8sUFmupFDl7hFHhD
yO2WWylUWuGPUagvLcqgVWrQIIEyJFRmht9nsigmdsYrTj8X2r2d/KjrvVJuahPhBKFU7EjQR0iA
9f9n5qcREdnZm8ObcOWYb/iF6uZv35itfhEnzUg4/eCuLEeMVwI0AJWnKDdZTOH3wWdCgiqis/Ga
EPymlEjrAuflDG5+URmHqeokdOiHt9vThbnoiUFzNxSICzXGN7svGRBYfBTz4xPZvTtqB0JPAFGc
1wchGlAlVszizbs8lf823pDQwP72OjMW1S17+YdC4unGMlGRER24SmOtMVAOy4qwDRd748yKhUMe
2XeDcwznEVGQtm2v9NQ1pmzcNG/O+bg3zgqkvHxMF3Wuwv/26bUcuErmIjm6bbV7v2CmxMXzzEQm
P0sLLN1LboYFS1Yx/E9E3uNCq6/ZpA19UYtyjKuE+7GvrJAhTuZnM6nkHc6ewagL9y4LjO1RNdaV
t7D9jP4rpS8gjV7GDdErX1WIBDe/guVvmGhITftwlLdK/aR58JRnaeVbBu1D8cdXZG9Gq1daoY2n
Fj/6YktIhvAy5GArjFWIIoQzyHm+qvl4ApFULftHpbtUu3jGz0NdI+aJ7U/zqbNufQ8BDVZKPR7T
S/wd9Td0Cmfhy8emN1zuQHZweHNQHZnrFNlrVb4YlLPk0Vw86Qg7lb5D1rG2m96B2aIp/e+qsgfL
twrLMdvA4Dfz5qA6ZgSsKOWFC1bErv0jZco7Rmpf82I8O3ro2pI7fRTsm0wlgscMeAE28PAOlwGr
BlrfesLDiOa+zgSOjUr4Pxu82Pie/m6a8MlRKzZmyLw56TsoelzV+O3rpwsmPLTOUjyiVbumRaWP
/lGh5Ge3JUibZiJpao3CwIer0WMwr3J9QL076h7Gu2BJ1x/9CFARtbW/ROL3jlij6PW9zs3cdhGg
ef22P8D9smQoNK+W3F8rlHG0uORCqKtuol7gSzAxvqcOZOUtcHO9c7TGflIRNTRaKrwuWMkMVThp
ySFXwsJEonMZELuVmQ5xiU4LEW0if7AuZy1OlJnVDE7NEu67/R/J3O8YcSHjZ/+jJ9SKLJg7g5uC
sVaSdh18DDtQCzDo7tkWrCf5phE4vu70w2ebxIvXVmcUYjVRG+TqwQ+QT9j7+P6LLgwG1hHK+zz6
XIM5LWPTlCKwpskiM+jd7SW0aqRJ8j7YGDgSI2xnQUEogLMBex78wW1G9EJfG+6m0DcifPbynRn8
OW3DbzkRjonqoqXr5J/MIx4ff9MT07nXkIU+mdPYYUWcyyvvL7mqUGCGHBYXo6+IaFgad9i1KvNA
rvy4cG3FCOO5nr667uxFgXm9KSCQk5LTIUuDUROdjI+7M8PYxxwqcCNBnFTr7JONQvVntEmsRTgs
8USpNCvZPJhotPZfmb8hh7e1+tO8NKV8eaQzjkZGCjOfpGAqveTQ4I3hqgZkRNHIGm4/zbmX4FnJ
XQfLfUlI1RfNrHhKRD1eZEgLtGPHKEfr/R/ZxiEp5FDfE10Rmj4uFqOzKjv8yovjiYAGI0eIbRzG
UijzVfAgI0DNx3824V3y753ZgQmk+e7FU/2n7zhcoxYSe412PinX0hFhi83MQRwrlq5SXXPdERts
+Lxw77rKEMaPJDxQAJJdjNrc9Jp9jM1/H5iXHdghrKsanzJ4N6SBEQStX+lEM/rDmyYHYHmCBhFn
E9oPR9VPMIga0TJPj4w0wAHCYImTLMZ1Xv1HnMIJfSMOQRWCbUNX4cKAp8bdI7D05/FVX50Q0n//
FbF4f8qXypUoxyQtsnRRTTnC3f6sQYguacAfpjtn9UXE5Mcbn6WFgdapocGa8Lp9VOVjodaS/qKU
lVeqpiKxcsI4PNqhaj5WYElJH8I7KwixoLyH0ns2m5TWFE2iU8OfAEsoigguna8rVNODlDilNdsE
YnZZ1oJjf/hg68l4V/PCNDwS0SORaoJwt7p59eYJ9mY2Xc2KbHFYNYvSmA0tG20n7B395NWqUe/Y
JBvLaQfNM2RtjAPP2O8nTXJ/MvsbQD7vaW6ZbDJlYrDGvUwtqpoypZ59HD2/KS89Z7JgGs2YhVdA
quHKIv/XFftfGe1mzeEU6lbVix2h0A0IVB425hSR2q+xtuUbhoTicOBc+kfx0WiIxv7eIXbuIGQ4
HHTm2vLKFRVi233r/CgqaI55e7dnKlgHwz0AWQbdNU2hbfpZAocQ4ZmC5YVjWmaRAtqjQOB55czI
miOnTSrRhbMdfXAQxo8bmeXPI2E5f62g7VR/j1E43L7ihQZYzD+yok8qjvJHxV/XV5YDD0qTXG0n
+s7mYEJYjkCuHgUlPp4I7YSnDZ8dzQ9PlcjAsnuULCcu8Y70CP1E/pT1XBNzeAowlMql57oTSPDI
Q6O2JonE1VMUHwa4RPojZnXRZGVlj8Gyh+4/NONg8WYBTS7buEDhg2X29Pt/c+UGmlVUk/bg0k92
Jp5JrATP8V6pP0xZzzqWnH2Tg1KvzN069H9PsHB1L8IiEf+ivEdwCCERZZ4O7o0rAyh2X9nlgecd
uUzMINS/6Pq5ukzzDZ9jznAxjh43MqhhhRia0CF5ry7sbS0jDwA2RTL0n32HmVSB/WHR89+ql5Do
Uz6ZyH3qF6YLp8SKU+ocu8TdkwVRDeUH2lF7W1Yb64j4+cZvYQ8ef76ABoHnM3qUQF/Jkw33jvJe
tZJiW4t713qm3XphiVFGcQ7WLsX8A0cE6KMjlGV1Uk3QPe1HkFKwQx4LMXB+NNS2XoKLWw4Z2Hpp
CMBaO0iKjP2QX7cUdPJrOHUiReTszth7Gf7esPUlNfLQpQYEXfvh/Wt+7xCUmEXT9N1ThF4L8BuJ
nlDRBQLaD4hw36N3heMYt5eADFrP8/gbE8mPAuFLudbEwu3OJSn7fBOaYzdwXVf3JJ81cKR3wJ8e
Av5Ypgu524CUZrSX+U6l2ANCc6qHeopZgNualCdFsDI5x/Ynbyc0i4WPXbeqFxdIf+ktaC3CEr87
16XG5ESTt73zdxpwITcysMsJxxxD72ajCRCqmkOKd/vKCI1ySHlkKZxnllwmcTfSHiJDLmBbRnVa
XUEzkWcHb9WKgsir3s2K5nmC/alkxkAltQPM9PJVg3Udd+aX6lmCGp4GtgONFNG1HPMwf0LBbfEU
JjxOnlndQQyG1aQVOjHwAUU+05ckmcINWq7EN7Oy1DXJKz535F5J52/C/qolOZaenGvuw2fkblMC
ZbxyS40IjCJWrtg8PkUAmX4XO0rLt+vORXC5cjTMDPmbDHEt4UcuQTH27PJe22NJqPQ7nnmgZ3do
DpslASKtEl4P9IENf+GJ7aAfNhBAdh+YzmTnzK+keEUP6//lVUwJ7wj38kuWNzFgM496aDnKSkLk
x6TlCBCbd0SFL4R09HkSnfny9V/Eh//pQvT6JK7+rjBKQtiknvmnFxPNpFHKzb61wjoK7zB0P4XE
Ty4HHorXdllZ55f+muG/uAYYGJiBx363g1i1NA4wPDnat0HeXTGfas9jrh2CzjNksnQOcTFeJdFq
1A2eJ4D6LDFMrQDGMyQer6McqHPbTOk9A8FWsQCoC7KEKY0475BWr0LCOLponaM6cwaFMMvtr296
aroUBiHXjK+gbY0XEZ3/nZtdt4iuwtaPuZL3m8FRJfVci6vT3piH+6pVvLXZGhliHzt4l12B0jya
2A731AV1az0NEr72QimJELwwR+68xi0fL2synkS+z6yugYj3NBI2WKGRl7PNjjpouvJfKMRXHXi2
3zQbzbostL/sjxsk66OhoGnQ46PKytAO0eiG+acGHU8bMSO1ILARk9+yd4YYW8mJFVkB8HynsWh3
XApAUBo4sPKS/TXA5Qk6RuphH3RIAfzZusgzXlIPj59Rsl4a0+u3t4l4UAZxe9VCDWIZsOy8WBgD
w9ftjTGh/L5uhm2fDgnoC0+bgTa5C0WfgZDJ98xIQfrjwWfBifaB93UI/KHwRBvI+FxxZSqnvKJu
qDnSkQhQWagCJQhAstTSyjTKO3GUOovM8/QwHrLFDNv76/Mhi9VrZoPucNpDRMsGuO2hj1ELlzz3
3AvZCudirqgKLQ1DDui+d9LPFom8/iBNq5UJBk8kFZEpj4XXPAdb5EPDJKFcsFnYKBA+cY3IUjD2
YM3FzNOccSXCbjl/75Pvr7XBNxL7K74EkWol+sAhktWy84byvFsWtrwmjrajEL9V9SOYNCTmHEFF
dha5ldxSTWd4iBenYoe8Cakwoe5ZIifytoLA0S29gmlt3VPfGKkfQIC2RAIB3Pi0qZttqbhpsbm4
nCaBBOiStq/UpeQXiC6tZQ53eXWJ/kqTS4TCkIIvekYzgQyTfmxwAORCf5Tv+OWl1bG0w2eEoIS0
qBonPHSH8NrS0va/yp6QIW0UH6MDakizytiAQ0TXy+MLpUs0ZnVaXPmnjFesRy1ldOEp9Z5QnvUF
JkMTDszNu3kGG36u2Ln13w/8LqPc0NxSchulaTc816RiFdNKTCsRBuq75YlI+tIAD6eaDVS73Ufv
DaQlTNYbYNpCmYQIV4ViRqwnNbrlKp4d/29VsCTnOU8rHnlign+5S7eCm6nLTn49P0CYyfWAlxkL
KoC5kuzGOM3a7xPf1OiMO9rZJELm6RFTUbBoA/EuArukahdU1VesM54oyvPleFJqDka47TB9rNzh
UqfcMZ6jmRZ0jAPwKbZQOZwAuJFxhM//2fl1HC2MY450/WCI1JMTLlGgSNblC7fPby+QwLYmofWr
3v2BUOcgTiu1qlVxqQwawaLOGWivttXzVQ927fKXA4LtFyuOPRoStM3o1XOUJMA16v5Sawlsr22f
0hVIH4qs8At248OmO3IyXN9EjjCnqVJKKfNf3q6/EbuxgO49NOmm/D55zEUws0Az8hXJ28q22+SL
rc+G3W+FK1wPgRYF6bE6Y2gX+zSfzQC3922RnwFtIEq5z/glgMOc1L4suie2cZp37MVoXyfD9nao
fpTtO8xTZtzHntIwiaMfeEw+h0IX6+8TE1yDJWf45L5ll03krcQce5psnZICn5Idfup4l5RuYqH+
i1T1oIK21oQ/MczCK2kOax+FVR5BarkXPu6tiRvoLMjtqU+1gBrTJq7AygeM4z1VGl5GXFTHbigM
LdvJGDIotjhHugb6peCKJN8wfsRToqpN6Q/IjhqeiGopyyY/nCEodW3GtqAzmReZbBrYVxmBOnPY
BhltAF8hopSrOS9umpgW1vErlRnXiEzdlRfkXy/vtWxpSayg2GVS2+Vcoqpz5JEXhUHtM6FKAwim
mAuilzFDtlRfUfutiu+UyR/oGV1V/ebAzUyChh3RAvPK/ilTr8mGkeC9my4QGFpH+cbjs2z82wbU
+5iXH+tBcOsnNPGKrno7XU+kPas5xcJPg4Om76OqVo9n1DCzHE3OdsgbY4kKmPal7HbOT97Jxj6t
ca7l9o/pJAUOh4ToCz4W0IGF3pN8QXU1vEuSY5KntKfv2FPG14GDlaAvP2O1N5WQQ7167M7Gir82
DxrqmF6Or7NBgi5fb95dUgw3QpC1ttrQHyAFqzc+zKsdqBez4RB/uQ+MPOHv0cfgnCMltziwnwUH
HDM5d4OcItNY0LwFOnxjj6+xKtjF2QMO4QR23ehSniKkUHht2FJH1UjAuNi35iW6/mAd2Z/SoWnp
t095l6z60R35ZFMzPFU3+xh+1tazc+QMFuBrinvOY7Mzq609xFAQShJUYza79FvsDO+MooGOyKaT
VUv/u5nA4xlJhGNx6iWX+sleUIVQwFnILzI8ro4PnNGCNyz+Sj5HzpqNcD0iaI8rZ9GuvK34XIYZ
s4K2utRzG6LOouv/kCLXH4vlgSnq2et1BvceAh9CXllVy4nXEePZlJ55kzduq9E3noc7UCEaRu/W
oQjaSLr4XVmQtxiHAL3vnhszBn1js5cgy4QNzIGS7qupt44txusXfse4m1hIBr4li9OtS/Lf9cxN
XweZzoqqxyJopyZpg6UJ7Pc8s//Q9Y9FhSAR8WB+zidhsqsZfKl+OVxLjix7qzUroeMPUGRqbOkf
vzqu9qWyYrHA6++DJ8P+otM2P42nOmxVDIpND6PA5vQm5vs5THiq3toId2j5YXBMDmbstcH9FuW9
h6DVJ0xaLoxQGvEgKKEZVQgsp3ZqGPuH7bWafHzAiDUp2bhHhu5Nslf+IrorfLvg5CdsJMzzoVy/
8fiiE4vvKuy4VJFEsGhzkGi/VRFFJXo24tJUEgKofacyT5NAwcPDG0rnxba+9MUZuyT52NZUvM6m
nC+sxynzVVOj45hmN7KLUvTBaifnJDbfnUPgQR2sOtekmEMJUO5J2tv6kWDCiUdrvSDG1JFBR/K+
pJ3Gr7jvNCCivfDH+mnaRHYHz4cIUGFitEZnFMtpC/Sjk17j2odh0R2MksbuDuqwim+UCBIr8BdE
NYQAjWoHmvTsqJaK/0P+vOBFdRf39rCFbrdVgDn6k1Y3LgzUbYwYHmUC7/y2yyAbwq1iWAUi60vI
f4cvplG4gZvDllv3MAkbVTiEIRSa17Ltzcapc6HIEmeWBLRMO9dnbsZpMAQjCIepnBoLk7Jx5qzU
vh0Zn3lLlVyQXbuZhHV5cIGfjerZs2+eRIt36rka09Mzea8STFuHHkI2uzZxrpnFDNblLdpSPIeh
0tHRVuzneetJufWwR4bSQJlxDhwN9Mt8Rb1kg7C70sZNSOL9oNBkh4s2XtbtuFdJpfofty7BpJ55
Oio3A4qjZB+2XBplzOZl6RCJlxIN85Y3sxS3qeAnP5LvHCmvtk1MQ34mOc7yprzjr3FXnZouPd6C
UJEBMrwQzVy8GTf60O/GlKIoxlj2scxeoCUa7bAMhyW022WHqSCD+lJOV7tG1n/EjdpcOBwiMf6M
aj5D7peXJfo2UF6WcslWhqf65Z7I7ZsgA1C7PVCqnPDOagCeh554ncndcrFo4Ch7+j2W40wGeMx7
TWeT8FB9DdtJtMiOCOV//1dIlU5m3BVSDbicifn0CLvPKMrJWmEkAX/XO1x47RSane3bKnXINWXh
p+Ox6Izv/PeInYkFrqKOlD+pJ0yCI9qY8wtCvkmSYItrTFWgW+KBELIc8a61ju32KS7V7SPC8yky
6fWy5lVmx9tbMpkC0TVg1RjjX5sFeXRwjZYIUt4NAg3u3bHrs2FnvBgIWJVjKiMuzToCJyZRQ786
sJXlhkJnr7ckDBTh+3on5j44/5nat8avsPIHlTXAaV3vGPiTHDYon2KD8CfAV8+FGP7vm+54CipQ
0hRx+ovgXuwwRZ903T3poU+oChzqcV3Sg3O8XNZl+llJ9l/5wKdkMLP/kTcEQcHWEiyBeWG8rW1e
ScCtTPNGFNfecg4EfwV5YgNBF5VEr9jtn50v99Aypmw3uhW4XECjspRC+WPWo9lEOxVF2Tp1f1Jn
IRQn1ZwrUPUdP/G215rRmBVcbo2eymxLfTElmcWFaoGMmrIDtDcO+m7ygYxfQ9dBvebn6Pj3BE0D
96Vqb8N8qrIncnCJJQYx2IZbFIGjnuN92V1gMP3VlQS2fVu8135SqFSgpLj2nz7UQCPZUX5GMf35
D/MZ1uP83V71a9IRmF9kdDhcGqzci+fSsLZg4wOD9HdeSvLX06pNLINr5CftRO72FBUN3cMV8pA4
6YD+m56nGVssYHR7Ctq0P5vgoGg9PCm0AJgUKa5CD7i299qzEB9FKvga6EI0M4BDeSoikB/c70L7
bqqUhmxHV3O2ffCvPuK3546Z3vox57R4HxYG3GdQ/kY9VX2z/qZZ/qDD0MCClFDW/qtLlhIgBrlV
ndg/qHLxaeelpRsp0J9AwXBYySG/777R8pd2i0NZIan3+v8oW6O/k7VynX/pzDzlOqkVVRk455Mz
xlE/fe8C0EBTutD5O+8DRyA6PiWTkiW38r0hRAe1ZQPeB3WAZl2dBirpV4rIMbvHmKG7yIYzWE3Q
3Kmm8AZBeNyw2k3V+lIl//qLjte387hstGMa9xIpUrx6/7mDj5V6GU6fdWgFHQX5SZ9zIq9z8kOI
tgT+MWzhUJciseYcaVTpAKVpSYIuUFkaxT4jJ0S2i+Hm/mdTeIGwVHHRRpM3Y1cBmQF3p9ve/jNi
P3WQnDrhPoJ0XAoDliUI62Auv5wv9WXL945U4BpLQldcXMeXvzcE/j+roR7yf4ZH3hZOgLE1elpN
qcTvEWX1U7o1ubxa+r22u7AyJdjIHM0kY3gKdsjOUB1hs0GqgquGvY3VFnG3ikfEQ3CHFsUwIbOh
VVhs764YSUdeZiy+RMfBcSOk7GVtFGGtmtOV/25tM20LTdnqrgrUZSi+zxKVjCs6DXsObsXvBoCY
wKAsycQ/fwHLkxYCkGa/I3kAU6RPEsvLVwSrSfeaLhkeVckIEda4t9nAAYB9Ztjobe2VQoSJ5cdL
AzRHqj29nLXkZqzM5cwHdA/8cd5104cYMA3wUnBNba2RGcS5BNog0L9KPZ/n02Siwg7S8ZtnDOA+
UPlh7/R14OiO7YCx4m/0ZKWPjAN/rJ8GUqs2/0Jc7aB//ss5pkhLLSO5CwfjyhDnVVzKhs5bZLQQ
ykU2KofQg8tTyzCgLkknEI0uvA0d5lPCzVY4V2sYv/YjzLCrrADSKC0UV0yjfcdCSWq+t6uSnB74
/N0Nh0w2A7XDlKJkHbkpRPOkC3gnQWPa4P5T0n/yznMD1EDg5Jgcde6q+uSxf1sRQ2Bf+oYT5wtx
DJPaJkCS2nmjAVzQg/VjGLLVaWxS+DhOy1T3u8vV+wkvg8Hlotd/SyXR+J5mAlOHoXxJFqe0p9kt
22kuy4DofPSS6xkvhe1FA7VAiJOjN/61BU16MIBWxvwbWlLnXwrRxUQDzIgMTF209DNuL5KapeeA
Dtaunlr/3ze31wKnb0kEIkM4J40EJh7mrBSO8+x+B4ymrvK/fbxIBiKLzY9aHgJIP6RuHhrY1axB
Bq2I1tRO5BXEJ3C6AKg2jZpdzIFsTgWwB9+1rd9wFTWOWej4mnsVW54G7a8GDr48H+uny+WDHXYx
DK4GWDUSx9iZj+16F0FJ/TVxgkrTuGoNvFm0tc83E7vweWSGfut6fKCOqUujTS1yWC7I+iV7mo7i
t+/8ey7dkiR4XQEbp1VgJXrk0NSNKcVxJs8PVa63pjVt7Vx+yDCE2gj04WgKZrLmFVOhg+9lla59
M8QHTFgso4Dx72Vi+GICk1WUlz4m7mJX7mCWfgjuacdTbGsHrhQSX3S0Fyi/gBspAlQDPi31qB1j
v3Si+qkBdHQ+2LSKtOnoJMZViA79AkwqqAe6t0mnsN+PlWxhtqp4oOesYHgevbVm6drt1MbcEdqT
xppOiQFEHb0JA3d3mrO96xbQgCEbFX2pE2FZty1cbFbuun/ARFA4hr6S4ckIaCFR9t7Gq5BZUBJ8
Sx5m1evNp9DE2rDhj4/gKLSsTV1/efYffy2RqUxlc8QIwYo1OTdWRXBVo27CMr98Rh73A3bMXfce
jS8BQSerrqrnsjWxyucsqJvGRq5zj7E/WSTQICk6yuOMDQDuJzNEHEgIWiLtoambWTI1St7OLoyI
+4UGD5oiCiEIpL8nVXpxqISXUdqmco2mr9vQIMx96yDDkSeeN2mrJRJ+saC87vYsQZdLP438feum
Fg314MD/VioReWuTDUFWcJxczw5YPL1XmZY9M47MY8qb9+wstWvmuanqPGJxZ1jPjyiuwc3sRqgm
cCh9+YT+AkgLI6DIFGvo8PH2N7VbeINEan05HatJLU8QzsEaxYcx8WXGxunqNp3pT3OkVRsF2xJA
dO5LZBWzRLPzvk+uriaiX4gnmfQqq2k4jXoinM9BaaBmnXQ/HFgGCNOFqz6WIa1zgy2cm6IzB/Sh
LmyXOCFZYYz3KKKs+9jus0k7IG+3WhQZXXaXx7JVr+87yMQ0jrC/erGYwUTYFLHrx5gf6VRtX7E8
MgQBlmdzH57xO5Uc4g2lNaLzJ415VeKFT7OOqoFyAJDsIq6LLSEWxKNQORPMzWipWbTOQqWX+UbW
5CuncMzo6/aSBZwld9yE/lyvNQEt/GtrKThH0Dfp2f938Cdj550l5ThQTwgUGYkb3O3kQaY/yXNX
OFl7VNjM4KP+CbFmPWsihC2lT2kSey1ivrsAsjy1U1XvA9aM4XmqmYVeWQIRGk9odv7WJZdbM2fI
nQPUyBmhZoiweuL6lgp3s1G43/xsH30bdHSZQNCigQ+17hq7RMwRIr7C0z3jpBAWsHHAy0wxhHk5
+yspyrSe6o5j70MZv43hVrr5U8vZKCaPFo7T+zGoPD6n2r5UT4J2m/9rOPAxmcxDUPwOV0ysIkvr
i4djQZqrS6CfJlzCtpaZ65Ny2qNCzkFSFO2Zt3hQFLW0BiPaOgC2SzOaNP/TULaqnDgeeUbgo1Cv
/56rT04Dbssgqg3nX+AlZ5EzpAVnIn9Hb5pNA7IE0yF5NGqrtcPOzVhlVBA78Ohxnf+qpIXzWakL
U4dVtYsxVVi3HmOSQzDgYqOZBopbcR2kgoMf55cmi5hjTPpOFKU5E3CPWWWkoJmxEnJmJ4C+nH1A
IJKlxdVlpzAVfuHxsWagbZFk2DjqOf/IIWuGxq/MJZkwsmT2Zis9JfHoQQJNLZCrnHD/3+xsWio3
s68wcCgC9XQDt/EOQZx0evGf3a93OTf82ERZ8eu2jXfDwpk1U/42+7I5oQL42wBbrkcgFeWj9HqY
Nb8Rps4GDh1gWRVDkqqMd6K+thRf3xvxAIC00hJdRRtlv5nTqvu9u1Yb8565C2gvfDgMTaqmuFFC
fzYBaSTv0BWbk9WqbcWenFNNhcBVGwm8oh+aQMdTPpzrT8+FievSwcUE7hj+Hla9XwofWEKywpkB
BNc8Mq4L4XlwMPmebiWFXUicnk4uWNhsFURYRS73u1nN8IMOg1BPIVSgXx7bwEef5GKvfQsAjsvZ
6tsKEacNQxQ9kEmdJq/2ew1UARsJ1RmLnk8ocqBEKjzmh516o9hDHXR4KWLkGTXmKMi0NXAsUiOp
4pu4dtGjyBcCOnEBMRIZUdV0eydD91SDIjUkqStJjXzUxsX+aywbH7vDm+vrITPFDCDqCnarI0GP
H32xb/o2WcMAJoP6QS3JZy9OMHI4NICCTgI4VEU5SjE3RnqYSzXlbD88QVGjhO+T5Qcv58G7mHP4
Oc0TVSZBsqvHY7NE6nHEHonN6+DdmCVDslOALLUWWVBmNqYaPk5YwiCPbv4tCJS1gppCd0DkPwoP
yEVxdXTAXsgE8LmKANtH6lTbCcbANMT9Qzl7Zv+OKqgFaPVNN3ZVHLxJRh61d74rnT9Rl4ZMPSJW
XruBta/n9D3QIUYAiUJX+iF5t7DwKGfHDgVp97Dq7y1PhpuXLP7bpfaJblqVGp2P/LdRhawDrVAE
BlihRL1eqpu8LcRVIT3V+JgN1tRkl0hGL8g29J3nBSvK39yHpHphsRRryoViPRLLdEMKNM2FyYaU
McF3rNmNUCOStqjoF7La8St3ko6gj67sC3rZvbS/9xnnnnHewcpgodWubww3+4AGIHOFuIhr2YS0
qGbvlGJU0JcZJ5zR+6X2LX2CCuhaehCklQEpMbS+sAkVoL8QY06n7XGKyoJeX7VKTkX+YYnAHJA6
PEjmOIvtu7JDgVHo7SodX+RY3UOZ0uYpUjm82MS6uI+BiFyGA57w8RHItxzArknUkMLkLNpetYwN
7rChhFpYoTO43SaDns1S+9SrMmEnvz1wiNmBRfT/cb3vjJFqxd5QTjbTaD4k1ewRTvHtdI4SRFqr
QRiCBiY7Y/mWULE+HtbCIaUVIvpo2NHebdloCdq/00yjOZSrtnG8hbbj9eOr9lQomihpelBgEGK4
QOGHn1Nn98UkX4LtXQihAHF8ms+gUR8c2nd3TW2g72f+gT1f3qPTOVhJXYTV0+SmXB9CsRoCCdmn
dvdAmNhOW89GyUMyLAbT3zZXpgrslzkj/NGODDZISD2XRMz1oAEiXywxHichXJqtP72b5p7jAofJ
4ZPs2LJG67CvTAkMXqToQPnNf9VuEM/M9vJudzs5MOpMMP38msKpA0FFPD31/gAByCAh3U3zbMdm
rrc5EXBVhgYbucQ2OYT5376nw9/NAjPAe7qFNUkiNo/W0DGtAA+HCBx6DUjy+VXk5AHhASmjy+t0
NA2mfTIcKDfChTn4pRfcOC2yokKP6cvZGDhG0ypUKTNW38vd+BvldcqDRXmyXlmwCa7ENK7ecBt5
POAyRY6tdV6oVnZfAmdG93r2a1pFCEKUsA4vaRKE+1OT8KEea/jM08XbZTNE2KLOYCoUdBBss43H
nFHyhHv938INhzix4e/mgnq5uqAhZ7EcizxOZ5/4D8YLQYNHr/BbZc+CO3eJUCF1jwvNMwIj5stm
ZY259p7sUSv20I6XFVKO7mBP1GiEKMxAm+ijvlKSaPDwCYmnTgcbw24urx7qojxuAfa+7AlP23YM
4BztfJlU5Fh+xTbPpbl7CcIX3zRKPODdkA+c478CmQ7T0o0Pfc64BmX0cP3CwhULV9ofkyCXuI0P
avIS9+EM6b+fU5a/7FHy5bhje/1535KD2R2AGariQykK2pcCbv9QXjvQ4jZAZkvTcL8k9FOPpkNg
2rIKST/sf6SBX5DEEX8GzuWjFUiTQwPvyHOpNjCwnnlQZLnt0/ePyDQSHIlIGgTEOjOWIcWZnDXM
lC7UMB8mQz3izN3nQnDvAYhbOcI7VNMvslbGPzbQa9UNPJUhm4881Mqedc/SBWYex8uZ3vkSPwuh
Sitm3BufIlWhPaaux2TlY5VzuPourZ5m/cO7ZVkpSni5kUgRwiN9TqPmMPldMRbaIY27Frx6oqxX
aSngebJuopkv8e3cM2al7bhav1FA+JP096f6bPfBuNrYDOQIz5ogf+9WR2jPMt7BKEGUOk9TlvKA
4C7mmsODwrQVs57fXsbl92Dlox+Q65mPT4K+7aQyUv7bI5wIcJPnhsNm5Lfc/KeDH8MaPK5MlP9g
LJUgcQpgJiIY3Gb/iYnJrVo0Bhft/zPZ8ZyI/2mvvuKPvmcx2wB+S327+UgKal6nCf3JUFuIzurB
Sf5m7b7LbVsmErMB/hm9HX0U8cn5jSUYFcKtt/jCdUCw9jV66sJ4atXjoedED45WrDlefTos2tVo
KCLcvN4PQYxjXVn+MdUMinjVGOegZvOYjLNve9ncV4F9D8ZQB5s+A6HwYNwsASb6+UGJOezoqN3L
WUDr44XTPxmGGMUxB7XnJ768pRGRpKYl/vmqlekabWxdcXhGPenCjXZQ3LpQN05kgIjXJTIFvE9x
Ulml21VM8EikL7ZGW0Fc0+V4GuesudJ7TQId5qZTpHPzYmNjEqbiGgRtPYsnzKR1N2tgUg6yn0j6
DZ+G08z9JWnp5iSsym0YNfFEB5qz6oI1v2EaUN0N0g63j3qvEiEybziw8NU7CVFET0IDm7Pzxo2V
EmRp/SoXdKAOCjUWVHAMhKa3S2X6cSgyG62XTsxStBnCIL7CVtgdFEBooB+/kDisez61rm7U+TdM
avZu/LLZPSOUILz9Am907z5VGdX+AAAGkXyxoPV+5GyN3x7mH/Ii2K8NatRsezmapekDl/a4E1Rv
kbDp9g+a8+kZzahrXs/8pqBaNBF8oIlvaApWjFlesek/9+kOlwKZEe6BQZtUi3RNGIzauLyV7sp6
zPOvzgkE+20FsdTq5m7/U277RYZRKcU6SqyTClx9CSyeYP9sxbI3lG4i8ag42NeuqB6x5HaI9eKH
VSkxGP9tCaMi7z0aShOr0KCRWXy6iisuQ14yGr4f9lAWseTuqaTpmZXp7xGKKt9hb2hpqfNEovVc
ahJpEVrpGIb8i9agN2PSy+BkxGQ8IswpHZ43/66MNjNKlc+yR7sC08AstsAj0cA9ioYiWRfjLxUY
uUJchaEJHYxK53/7lsM6R6ntjZHeB7kWSwXRXfocNJjbvq2pfN5vxKh7k9Qnh6E/uGYHhqODIHy4
kzo7r+Jm/aG2YeRTQ0CS+1fFwyqOTEFW9QWr+coPp3e1bQTI9bg3qv2rmTgiWdXzMot4X1TNEwrF
j4JQHmyxvaugaVdsbWHgRigussm9NyWTytRjn1Hh6JEoYXkPHjbo8EFnrdKVZH3bXEW5AhErZPSq
WIdPc3D42YAXXpcn8zal8r9ZBbrEqpdGcIIBnsDwGsDOIV5PTGf3OgCz1faP1YXgfZrxCPl92dwb
9CrvwngiYRBDW8l65y/S0dQPwqS97VNmhS4CqjTcRZQimBcIsMS6RGOBf9IrCYLfY2c4w5N8hJ6B
W/6YmbtRi7cCiU4JmPd0cU5GbKtItgB1vCHcPEuldAyQ2uVMU4dASroXDmYmBYLrpQgEBE3rCt1j
W9/G9pmvOG0/Dxglgid+y0NDusKe6Fl6tiXYF24/aCZtSvEfZDdfIYjkhouTtXLlH5VXsaKliap6
PGjEAFgZ/RxcixQMP0rIRZxjapDvB+LwMUWpPVI26681PgA6DM8CN1gYJqS6dY0OtVAIq6mM26eb
NiR+rCQrqvzG1UNj80sVVyWGiMPwp2N2lVu/SOdYnwSWwf3T50DUC8zPSzJVy6HfALRgzALpvJfK
XfVIQROTpWh5wbyJiwG0ZCBCgiNE7PIvfZan/asHuFuzMxrVJJ8lJaJ8AS3CS+625WcJWXE8bMAl
5B6cQf3SkgGH48Z572WgidS3QuLGF4+A4lGsLviM3PR+nldCztKo8DoOppLGGBtcjOOXU+ZPjOWT
2AeZviw/ZgteAmKS4aA4YImsJ0SAeIA9s6mZB7yt7cGElfFRQTwojMFgBx19YaJ+jQndfVo79lAj
rcBR4WaEe+PjTAduGct3swVULYx+JdhyaJMdZIG9HuJjf+YFZY1skeATMDN6mG3wWcbIeRTDakuq
/9LxLnT33x5Y4xyb4uA92FSGZY+hUAVZ6pfossP8EqMZfhbLlJUu/Bp3IGBzGY3WPhCW0xl8WUHE
JYpL4k2b01+ywQq9VL3RuCnxnsvOduU+hlfs9tRjHUXW57RNHNVA0PZ+Cu1QbC2zGKCKwiLy31w9
KQGJprSstOypWm9Fiwms9QEOCfFC/GTXMHXOcwjJXaCsLBnwduxMbjIv2bOnwgk+sggez2fbjLcD
0VpG2zFNF+5kXzquQa/3kVWekQ/MpCIjjDAG4+6mNpR2dw2M04YR96nhykac2T7hUnW23xq8alvO
fDpwkbah/rl713ytkMwYB3DYbEEFqbZ2fhqRk5mHUR3SXBZMHDzJ439CQeXLkyEXIgxH6M+9fiw0
yyz+b2scAQKE/MCCxvUyMFwgT/WH5k2RWn/I/Ok+m8x9zGMv/xFS0RffSs438PTl01B5CW2k+CQh
WsvaEBg1iAzdkzPbZGoqKYVMg4ukJBapcr7M78I+485Z9TrAKIjwaEicvv2LPtuUxActKWcDtiUr
28spKZ07Blhtn3urf/iIgVcYOknseZEUJPUYe6YWUyPexb8vFDRDZeJIuKQu8LbQrNaYD7nZbqNT
wL3+aWxbICxhL1/CfTxh37Gbc2QCURNTmwO5QsKFCd13rmIQX5aJ3xUv3J2EmOD6h91nXiWsr26q
geVqfpXJh1aqV4siqCwP7tTcuH0ocJXpqGgfHVsBH+Hli/WH/VZWtHTiqf5LIGMwADOT0JvqC6su
5RcPsqzYEO3fx+yd6ktQ47ESkH6j9I6pB4UNCljevdxPmo9tYO5/dobzAu8Dm9Z95qcT+0d049Cv
yR7/9h0+LysJOuCDExoh1JNWM9QMvpkbkbWyKFDd7CAn0L91CDyiomCcUkwsqZM/byCLrH1TmAdB
zwKZfe3Ng91D7zoeJlNQ6Gzue/8DnyIwKqYIIh/8bIHF9gVcGgsjzXIaazOKfC8sfNT/t0zPRg0J
opmkOI7Em+HvR65HauFaLkWbW3z29HbOIT29KjEH7+mMYdHIk8w9QRCZ4xB08xy9BuCKjcD2wpVP
a425Wn6eUBJfSv3KUsLhOgOSDavsQ6Wxxpn+i0KUG+Un8u8WVPvBb9MuDBwFh6E2vfzj8pOZd3/Y
3K400OQclt2J/pzOFFHZUMVi4wwaivgHOnje4tD53bT/W9S7Klw7kniMGlefP1xM8b0/iKxbeSWs
NKRdMNO5SbTXUuMkU+Cu2AHDYRT5/p5fik1ueTLDpEBk7LtgorG4tcUKneIh9ALiVXzZvaYG8Si1
uiF9Gnp/9MIFaoUbeZCWq130lMGSt7H8e/g8ILp/SkyYzw1oXfLQ1bUov9dzRoaYcGKpNxL2NDfj
E0C1GWDsN+NsfSw8I/Dp0G3lVlT3v9g5WJCpoi5F9/kA9D/ye6jvAi0s0GOnan+AxHIRAmubdAle
8xbxO0XJ1uBYZyvGfzpqkzP5oUfY1YaKP522HDqchq1WUt4BgDwhYwwfQ4NCGQTAQdrGkDSQKXiY
4zfADHSfzhZstFgRedHNG+8Lp7oJ2/D5mNjWKDUVOY3mgqnhyF8auikkq+WikbzUWi8ct1ts6sHv
a4GUJ6BQ7Y06Ziqdvx+vE2mndjnyPBo03DT16JRlOBi248smgnqL6aeUgdL18rMQkSem2rm1RZU2
7DF2++0Wmdbi4y0Y88oep7Nq91jHGooYmrTk8mgF10xLw37CvbHjLBfSoUnPf0108pMhWYTDtGYG
2ORWwEmf1Y1VwPQ3vQJsT0IFA0PsN5QBBtDq85cy/b+nn0AZ2Ci/lk9/wv1uBccTOpfpVvTVXYEt
fUijb0d/62MwvzNfhvoW5FX4RIN3whFAJLyVOUoxwRca66/W2yub9ceajcg9RyPw7uYWfgjKKUiT
6U7L/X2Z1iIAgivL8tizerHBDq+VIJvhYyil9z6PhME/xmq4MnxL23rs6YJcmUcaV33lLXpY/tHv
6IRKL5gMQ/5Sc2xxS2To4k8L/ldrXuNzTmoSrOI6LEbzELeiufet//FeybW5zshCbbc9xzFFuA4I
bRakIRFzzX96ARcoMwmOYJVQfuWu5WTVKbWiOcsEPcVulJ6DnDxd7TRzuvXWTbIbaYsFDwuxRyfs
6Tm1MGADChlA5+wZl+eJTKXhY7fzW0Qi5AeoVa8TjBAghu73sJWx1BiF1zLmbSTwrPTE+hZuxTRZ
pVVeqRcy85+3tbktopT+zxgwH7Ealp31ZYj76Xgkj4YaqcUoHP+yC0vJqC3jgJttjkQdFV6DLMJ+
5WWUavAnrAQwL+EtMybHGxi0LrC6DqWZXNmaQbg/pWTvi4kRF33OUuQYGTwTEc4wDC6WGp1/bCTM
4zLCcZNHSA/5E2rDy34dgGIXq7ZnLwjqJDQ8Y+LEeT7J0P7hSvVFTrxnbNlukcRsLPwcJagl9bzh
/B9PP0j3fu32xJPj1zkPISUO4xmhwKi+SpIboFphWnT2vSi2SLuOUTkvpBk5OQclCgEqGN4Man0f
sW3VCF3eIIbOPY4MCToSwZAfp5r9nhzgCtPKv/rLo6E8X5rBCaY3DqejUxtyG0N4FzQvofcS1Vbc
wE1Jvv0zMoaplQN5/a0ma35i3WDfK7kijhHzV5VAAmSmwnzjh3uqedVgy11CRLSO1auZU7tdYu1X
8XvhRNWLL1D5fnDs2sJYmllfmAfFjT1agYiWszSZnU3UNIJAsOlfV2rU8+gZ2LrnBXiz5hmdBLoI
DHpQxSHxK/oQ5+Wyo+cMD1A+Nszpb5hkXBcnD37Q4+VP3N0k7ROy0M/mPJ6JHPDfuaxCND06M2/1
ZKp5sj2SaHwoiCck/9T+5MO3MRZSuu20oJiphPKHoMwrapgQpxPgSWM5fOktknJdBlBnae4of24o
UWv7cEsr/Zy1Es2InmS+INvsfP+YPQvQdn1zVceKEBmJGRCZpVuplziaxOFpaa1KPsvsT0lOPg6B
AYcFbkqM+NGKIfPyuBLsakDxvJK+bxjBtLdJSzzv+TAbL59xSxhy5vj+CeM7lrzZcZpUUftXUJCm
kVtHh5qxFNI+0/uGgkPp+uCG/yhr0+LwLJRCX0tSq3q4mIVqtVQ4SW6p579kPXUdSrZDGa5YVekj
qSsoeA5buZsy27QlBDPuocj5UCuDxF+M1daOB/8nXxDjWbJe2ZiflEZ2/+2MFYzPPx6XE+JB5E7G
1in/49nuvA50ZjTLeNEzoOL0ewdJtEpGQnGLiEVOKpjO9tA3nl0VFGIiQpaONV7yOw+tOochAIGA
QMyyurSoJTLZK1kavo2PHkQz10uuNT9fl7I6HRDeF1wX8y4MtpLosa3CjmRkllm3v1H7DEt0PdRj
UxRCfqqkI5kEmP1fG6usUg3s+T7TqzuwEBjNp8qLdMOZeO/aei8km9FAJ4BRPCg7j0SrpoHL9P3E
6gtRitnc+Waopk8zgigPKHfZ7BY/JbQTKZiUpp+4U9c6+OoYzEH1CmT4N6LhoN4aiTVWbI/MzsYw
iK5WAeodWWh/0XvvNIbA2MdoysvT92bu2fpSS6oOwr8lX1Bm4qEh05k0DDsFL9hv+XeTk1GWLIDQ
666teek8fhfr75gihJYuYgD6NphKAYZMH4Z4X+hah+eq1uvJoYWw9mGVd+FkpHYHLDViQuEvqg0Q
PQoHvwiEnVtNvSva7dgIpmycmWY6SjmVvYjbdFy1LXJBE16Fw3tXJsnCB+yy2eBj4uZe57J7jLaH
5zj7/EmAUJ7PoHCyTVbfaRyECm4pgaROCMcZsRgQx7nRQTZhHG6iaErH+4Tj9+RZ17dB2Tnx+GTZ
gEckh4/zabhnZVWwCOsldtEeRlWju4jSShsmD5gbo2QWep+1ES/GVZ/npMYqQBKn+7a1H/dBHh0r
oggjPYAz9MmXBmfbr0E92tYonljQWhq1gfY2zyhIVKsZPs7dUMHvRAkceF+H2+pJhXH5wBBgN4j4
8JUj2XsENmk8M4zbpmowXHeQrT3cBU/qOX0DpaiLG1xh8s3R/6wroXoAgnKK2NbUuGCEuu9a4f8i
rslaLmOpHJUW74bFQNaGuojFs1sQKuCw3MSuD25Uq7KTQ5j9XogGN5CBa6wXJckxx/CWGL+9Wc+X
Z+RC+kuex4K674DXf8syH4vnXQD9QnjhkJrWTNmP7sTw4BY3zgEWzVnk+NPvpQ1FAGHSt8nBrCe4
rO4AQ09n7R0MXR7rVdN9NhA3CryYfLjg6QrxZ3yu+ojZJSNSOjGyGrTMWFESwVcTTo3WCJohXkwC
wYm05tRD6qsP9xUK60b7C0HkCUYPFO1RF9Rio93pyFesyGYgCzF+2PH+0DJd2oZuPmZDUXYc4qgy
lRbjXqESxOgdLDim6a8Hwd2TPsA5tNbge2kArS59D+xYMecmNdGqgE7Aqyi2S/PqgpkyOTPSMt4w
SukSdK9v17rOuftj6zPZwblIAomNprNXFuKaJZASoADJo6thBojesi8qRV5DbjAwZKzQEYIu9jXF
pKARCjz/346p9nfonlDXkgnRFfHX3TcRsWYwldSLOIwJN7fTP/p+gRgwRu7QFVa6pbuekH1YaN/T
Ho6zI1yChb7MmJPuWibFuBFvHBbyKQKCkqN+48jbjHA6vxmcq8INx1XoQJn8AyaoLK6A1xceguPZ
D7QCQPAMr1HgORkVepbONmOqjjUcrcwzoSXRcmMR1aobUTS3nERDDd+XAN4Se6c0nmvDVYF5Pfgf
F0fSLBP52IGvsc0qf8P/9PTtecD1QqfrweELrCwuL/ZFRESr5bB+OMWYvrLb374vH1EnJHZmnyXQ
GVJrLwrnI4Y/9IEAw3zl61kebCXslhdjKeoGoh8V3ik+rSy8RDBL1XtTxVsHgpvnA7V+7zQetVer
G0p1D4nkbP8T8xALiG3aknOINvRj/rp2yVsV1OWIzRTFkQlEp0rcZCl1EZjlV6qPl+C7ymKQ5jFG
dRx/4VRxNvLNQw11L8fHLMPnLmFHf9bFEEA394PLVzJavncm4/EqQvy8GsP3PQOfo05jIO1hCphA
eApus/dhcBFIf4W67ptJskh4CEigRdL95bHIPsP+INp4sQmqAWYPYpsastMfSEPkexLQOxvZzH+z
L2+Hupe6sEqQ9oU6V+Pl9oG4COpFvAy3s8zgf/mh9IU/mxBMhxWZeiX8CvCQXEXLTwWk2NQ9gYoj
H3DfdKi3ik63iau0ha3iQINI0o/g08LAWsXTugxJNVd5Rxfl1UEBdUYZYhw4f4bOdm+Ohga3gRwI
bc0MpHrP9Io+vZ/kjiP0QwjVQjH7CqhRW116RPuY1GqnbdOy0lmP5gYVpv669Z7z2Mi83pdCfWHy
JlAATgRqVYGtIT+8ct1C9XeMTd/BTuOkbjvWMR4nxZCpVwF9kIVBsDQyeaCzmxqbxcprdXwagslS
J6kROuAie+use22jc12YhD7IcMv4ziWJ8pMfoGtcS2z6Gu1C1/R+ZqidfB4tHHbi+58PkFr3gZMK
ZlOqFcqC65E0q3NRqCH5re1fpTz4inPsvptrpTjHvFpOZc9GdK3LtsSPDp+gU+BWJDzqmgGU8t4L
jmFAosGXYI6i651WXiF/qVdJIJ06noWI/eJ7b2uT/BCV03FdNa43KBER9tyV0V+5ClMAklYaOOO9
zy7EXSpdnHzPDiDZs6sG39eYoPWDecMxxdb7lVcaff6EjoYOTd0hvqbxosKblCfirXZg4QwnPBzy
HxAXCmU/BCTmROjYwQw67F1QibKlANL5hY/li4r0GFdnOTBlGUSiS3z/ey6EzRysTzgN6jMJuEIQ
U0QUzmkk4nb0PL39rlP6w3+I4RhGpXaK+I3f+pDWBm90x37UZJ7hAWoSyoetIW4W5VgrR+dzWWRh
6cQ4shTrrm1DmDTA5LiRmCjlMEgurq3GjOJU2xycCDI3RHcGJs6JQS+Vn1rvGGh52VSd9yPN/FqF
0eRrz1pnfSQHYwIP+6sI2uLOsKU+8SLm7TpU79KgFivvh6skJAaVNjQ/gdRgLIrdindjj+Mk3jwh
eDT0voP5frwRi/zzm2M/XxTsDB4ssdT+3VPLUqXLsqHGmFKOCcFCkJOzvWda2D0kDxrbTCGw6i6m
p65VLlWFOx8gKKwnDccTUHJI70tiB942seup87NX8gO5AeVGLlKTXpGe3BwMziau4WvF77Wp5MsG
zD+wVCCBfTlsFGAOwSl3tL+pRjbYvtt7HXxffy28Kh8xk3f3sIZ3ELBT9DI/gFZFlCmBuU0C+HBs
VAsqY/gJd0V5cQzO5X7J7YuHYnZSHUfzTZHbST9Sa8/ntO8tMxy12zDutdUu8LrhalTEM/1Au1sC
LJc0URygWcNKljCJSqdV84syBSumI6PHtDbtRAOEBd4br1bzZ858uZ4FgmsziSlh4WIAAxTvvRAe
WiMoEgawqSgeoOpb9CJw8KzboPsqRaVnbn9Uvj/LQrGBCNZjXXg2rLX1LmRTq4gqeUQzWIc5tXAN
NrdYYVrNlLRBG7BpoYJpYE+A7UnyWEus0/rwxFs+tcIHDSX7ZtAHiaGMoX5oVqKSbBy96B7AaYmQ
k7upFw4t7NHoZKhLjCizsR7bWsBUrNwXfCdfx6vK1tyLKrflbcDnnnbjmjyX86UixQWC6Jo8fUrL
8GsMB1LidseMUnI2tbNc7qIwGDYm5Fh2RYVlCdXycNhhEZqMmDmjyNVhxS9Si0N88wcrkTmLMz9G
3kidp+ioEWgcP3p99JERqDL9o6jiP9N+HCq0/Xa/fAgwvVcgGcQvQwFZd8ZrUbDdLdi2AVwwF1DT
xjeTGytAFxOSldy2amDgLVPXHMamSPls7n9xKGAUaflOTB8/Wgu5+ojbW53K5xF5ntTOy17pAIBA
eF/1hcI4H16/Fz5DKgROfxM4456Zg99eGjpijwB8QLQCvQJg3tPGRt0IAcn0OfFb/z0wESHNP58s
lZfnadrAtyhd5X/WOt0j6bWsP49//igsGoC9zV02tWh6G+wq1zNOTrj2Y0jz6qUAU+g0hjkWJ4Eo
cW1wShzycemCPemdEEI9hJ9ETRLRRUcwdkgOkfKq4NEq2HOlomy5wlalkNj0Fvo+xkVgSEU/e6PC
yiLLrVbbUnB7ZtBkj3aojIL6cJm2+sjuZfizzLUzlVY7+IpA5lQm4wa8EEEbBVtyo9iu/Xvv6eJz
JczwXJePxvy1GriV/QbN96va79NaXCFoAaalxB+OdzC6JgIdx2snzadtsN9uax9SJcwENON5spAk
48q3K2gHw04VvCmf8m4kRz1Q2YVp04QIDWwpWHlVRjTR4BcaIvaIRCJj/kgD0C+YnXjBzsH1f1IC
cN2CtYuJAWSCY/4JnJRQZLrjDRdjN4KuMS7P12N4F1xTm+u5OFqTDVGzMltbetqReekSqY4kffwL
qkRqbmeZvemMF2IZsXrWu4EQo7+09JbqoRlqW7PmweKaIBf1HQICQ4SnAHuv8CzrE7LSouRGkq9C
a+apEDDsCG5KTvnZFNfWpt2jLRcoAuOurJ/Tak/SsVHFRZoEOBduc3jwgN7/J4lxYSv7p8ukCyKu
Zrefo9xw1f4Pu0PnTKqZwmBC6Jy31xG+HN5y5hX9CRsk9bdawEW2Hqzj4JbyVLh7A4opZ+66qfx6
VkdDLi18mwKWSTFNKMmsUPqtADzk8e7BBQslChmnGjkfFLQP1LREsC/Ae2q1XRGF7DO1PlKpM62P
Dta5TgQDJF7m+T4IDMt1I/odsD6SzJ25k5HPravFsStLl9yEiK2I2Dbx0w/vyjJwRg7Nu3YtbuF/
R7V2QEAwOPjxRXR4aYiYO8FWXIWGvOSrhXo7aKSQnqZ5soqcIdUgQcaHsyOv+JY9ekH9cgzqzqOL
oWHVTY7JSkh7MHQ5rA+AyPSrRirz9UzUAvrafXEHgqRl6Mc+gX40/zrXr/cq/sfNiteP7ENaR9H3
0WeCHalP+a4ZsKl5Uv+6pos9Q0ZYQJ5NMbbhYxcar+RW9VnBH8WxXK3EOgq8Y/T0aOMPbvev6lMW
98zYR4hPLsXLV+5Mjh1sLEFfi+MQt1pEqKqh1ni7Voua0mMpKYKRpxIYVh1eUnTr1GNnppkNVLar
qhdXrwkiW3wTAW0m0YAMDNL+4BqK43P+Rpz8lc8tsEUy7aRIbnOcbyq/JQZoKeBesUN9IB6sTNSM
iFT7EqKbRB1dmV9sgPLdFTA5A/DUOaSfxF7LZJTNS1jmwYd9bROGfX/0dYTyGPP0bfvFfJfswVu1
QMyi9hW/vdqsuM3QnoBV4WjmpQsfaLQ3SJG0qVpsQC76bmDoV2HNdYXhqVg/AdQ/86AD1ajkqGM0
cKYtZn1qcbos+kGfra7Tjxq4V/yQ5584tE0SOKC6U3TZXP5SCo75OA3DQS9u3rhTgsxLkeLtg+1Q
piXoSseFRKift3/whvB1vQtlpuEbAsMklx+KLGkgHHIKjL/SUyXLrCZ6uLZlgVj8co9Upld3lUda
qGjEbEJZV+spridCj5u61KfJiZ2fMHCMR7ZjTgl+koprDgOeLiz/6fTNgupk2JkHfyhOEQJMhcE3
5rpMbXXf/XTfdP2sFff7wbH+zjPVFg53w+syJRwwSeALr4UrRfEFkXHSjXiSpLoCNwDKF7BD0gj/
6FmeQLEBQrU3UOhCqy85ybhMwP8QxFl8JRxr7BbF6Q3a6Ff6xG3RBpjEN3LjeucQp2BmF7N8kMTD
SYLxmwKMf8aD8/96qGiWf2jXUEA/s5MjsDOz0u2bggSiw7YARrTQmpcjRFyLZ+jUOKJVL3KoHqfA
CeGF6sXS0zz6NHtaWwTPSGOa58UBzFrRK4avPh+4DLH/k5EDcUKdPEwzFCP+BOzHJ4wRhCCBnI5A
kFsHfyqFtsY7qET9xURlikLHkJWl7dAC1h5ij8HJ+2YcddwufvZ23RnAYyNd1LxTucprmJqiAaLr
ifRLOW15UC/r7wHFm61rG+wSV0as3ES7cx/BS+oIz/raKt1Ccbn3OlJFvKkLp+SGMGtyCSvbNb2w
QICiw1CkS3ggXdp4fBkCtOqud/Lg2KUvxyahg3BzwGmQVfVeyP2Ac+lAIeSo6IkPa+A/HdUWY/DA
LsKnMhe6vmAv1fOfjmhfh27w0gY+GfjDJ0LwLxXGSJdaDYpHlJsbXu/t3Ou+NYR/BgTOljuKLyjN
0I+95TAJi6+udRrfjbr0dycsAcARtO+89xUu8HViObSaYzGfCICDKTiANdwRRVCMVqU9lc76etE2
WYxWkJRbq+WrVP2dYKQHrSQsElMBKJpTahdgHhcn4angqKog7iz2c0RmtZvsGKL1Z9My5Af/j9V9
ntGetODWhLKrMzX7CvBYKnd69FIqhV1+3d8tEQL/hUBZog7YvRxMyYsQ3JfZjPszhG/PMrX94qv8
oZp7IFG/IAOVWtcXtI1ZDAm3+/bEtqLOO5C/kIl+bYoyIi9zx8kX72EM6hmyr4pgaoTtfpTpdFD9
08e7mO1bry25mZ3/4Z4BikdmC9nSFJbvivzS6H5Vcz1KrgBgdsScfcKlKjSdcaiZCdkk3LoBunfj
9Ax1HwLqqrRkXrxPO2jwUwedkbfywCqx7ZVksrE882g0cUm6JNX8yG1eogZoZrG508+icGfXDUpo
QV4w0ERMCPO0xV2Go7W5N8PtBbrOZLYJNxbu6RWVbM7uvS1FKvdtRaAIoUGq/+EE9Ywj9VEtuwaE
gQzRrhTbKc+fu+szfxChW+2GsoDbZutmKP9KxfjdkdNaomV7zBSRuojwxBXpri8n1Cgux9mVsf8J
5jQuWubxExsJi6hd+oeL+ikv4HpGIB084odVRL++iI/J1sfqw08RCgCt6BH4uRyASPWHjiXm4JJI
FyFZD0ASshew3EFtZqDaMh/2aP3kxlbELyYgjX8QNtfVqGSQiNhB+7Dwi17S+ASvQanLxlwh3qOM
FA8kI3IlYciiRARIhaPwn3VfDzhQlcKrmNVtlqq7DaNJEFxnBVQhce++Kwyz9uM3upf14s8t3HY8
Ar40+hL+9rMUNLTqAvA9qu88Gk1dRY0G8QWwTFsWJtlJaSgqYoUuNsxJnttMcIncjSbH0QHG3PPv
fRa/yfkubUzxhBUu3jECcI7I6Hvcm6GTaCYoK//n609rSWPXdEzHhoGRlYh7y1TGQXZ7TY6/EYJ5
srMQh/kPRjP97uhDneSVDMEiE04Y2TSNeVuumnTZPCNP4n1Fk7s0enqiKmfs2go/KhwQQn49WlWo
DMSebdbtl8BkehL7XC5vuc9eL5nrRMLVf79+8TAAagYi/c+eynclK3zsmbwj4pLx6GcTMYPgggtr
QGxvSn+Pfrgu7u0/yYM23Ul8lDqaxXBOwI8b7GqAvLp+ySwnfsYIdcweQXaKJ3z55jieemS/0+ZN
4wWJ+6UAkFPYchNxsNsVqUpqEHCCQ6c58QTWLykCaZ66iSjB0l6UUtm6PF0BdSO+hf66/gwTITwF
dIMtWqv++irRxSndSzKB3QgHibYqRV1wlCmEtRiA7z90jdCmRgGZopRtsEqKxWw6IiawW18gC0C/
aJlYRADtyPMzJgxxxv2x08eaxQdZ8NenIffeBINlAQlJn5SV5LDLNHAOM/3h5VfovrXGkxcD5YAi
2n5oPSAVYS00MFMs4Q08RCCON2ZH4AcRWTInPZdoEHOfD1ELOgBuceDH3Ke5IseE6z26KKzeF2LR
omlW+XtZhlYnoyUWB7cD1y7IWl1+fcgGUGdz7UAPQgbxB8JK3DCRaNCfKLcCvtgfa8/OZs46bvRR
ZknyQBSsFYVHzi4iD5rGvPwx54wtXDrA2FvTfLDPpBMSeOg44QOZruhmQarYfkQzR7fk2ITYZEz9
IOmwZYKPr4W+3kFCju5Qsd7S2vzPTXxtLW6RUWAQwzvzZZQqAoz3kqvSCVougmyqWhebI38bR+5b
48FFxCNFxQsuPUQ2KwXbRcLPepUoPZLwhRVbpq9y1KChOmHtG9xXJdtF4VwX3NsLl04HYjF8l61W
8dIDoY3XxnpRqDnlD+BqzB/aejsI+iuzxv3rI5ryE5jRzuMZYD7yx4e795efXcCcyJQs4GnOloEz
esEQL7Cg5+uvbvDmVWZctrZl+YwSIVpqibcJC7iqNC00zDRAhv5QSlOkdBHnP8dwUVjhhqI4OylI
oGWn1zZ5oYslPNK+KW1CIkne3Ikm3anxJFSRyeD9R535ryuPQ8YUgEB9ErfBBh674G+WujO831yr
wZZ0MrhWNxfT24JSST0jElcLj06sASbqHJbN7VPkiJPFOy4cRd9EtNaUQBXdJUFVXPqrSnqNMLY7
WnWsJmHCeUIDhroVKfu//J69Vgpx07cCsbENBFaZpVxfu8ZibiE/svAIM9Iwx1K4ph7kuYk/LlYX
hieqMFbWXHrJQDZlOASfRo7uqn13DxUvqysHkQNRFwnrPlrY45IIDaQjhYQc1ch+2k+IgK8FI3B3
PQjOvngPlezFB8qEJ9INawffFhOwVJeQRB93n02U+T6JwccnWfYpkdnihWaZ+1rXYeSxOpAy1x5z
6JaUB9E1gt9JhRdYhlEPLQ7AX1fQF0HHfnc4wov1R1gzxd4dJJYFRHpeIzZZQwfQjrkrE7eYSyNA
hKC6h2qCcd6pHLIMkZRVawXSFTltmAheIOGWRNFtIJ9kGd/bn9ewNPMlmK6MPiWPqN7n7UXMpL4f
EvMaGoD52BGjhc0RJJDW3od9XpFOKcI25TuWAG8Aex6OcW24UKc9gMu6REWYrBkuIuqtfsXKTMXs
yMiCQnlG/JjAbv0+kTibk84MmV1TUuCE6r5z1VRhopgCNQhgvH8MQ7wzh3/zz/RHvMUmh+wi9Jpv
zFu6NQZCABe8isYCH7zKCaB6ZaZHijnDpTrNpugBuX5V67JuStlFgO6OClTq2Y2UhUo67WwVnSQo
4R759ZGdIr2LLug9ye30vHkuuXvyq+PN7XLRP9/qVuyS1ZR6P28tvg7eCzHuuOGv8tN9/tULZLaj
xp6hLM6VHu2FVKVkixtQgd8LNqnHlCbTju27tnvzpe5KfjZWplwzJAVulSgLbqwApSe74kjAFaK2
zETvD389z5NxN6YIz5xb2Uh7cfl0g69pnCz0NQEXocZn0aDaCRvcFf7ionZz65IRTPspyaDvP6K3
zSp7G4QonoRYsxLctj3ChjBjgC8hjukdAXuvwO1GO15BNjaV4po3vqOc7olLYDjuMzmPkPjJj6eb
fcRtmNvb4HN2UMHYy/ecQN/Y4h1b7sOaUZNPAyWPnORsWJC0p6vEjxwTZ2UPHPwwnJ0kBeBUGPOs
/OU9qCMDu5kf3O98B1T6CnJa/mu+P4BhjwusdIyGLeADyP6ShpIHo/R/GPxS0kfc8z5z6zT5qS2Q
2+3xrEDWvQEWOVbRc61EZhEWpwJbq0VInSanLkZGA+MmeAaEye++xAT7qunjWdj3LrPiW/IU9KgM
duIQvkd2qMS/Kj3WzQePS0KIh/XmK2UNr6DHVXKKDgZ8nASZMNnUzAJRA8SnZ0YbePIgHRPORRCi
h92FuhiJE+uUWf2i4Q+JGpvsiWRT1hAiLX6zG4FgbIuBYR352gkej0FTES8ft+HQPfo90D2lvQSS
UyQRZ1Qd/AhPBg0Dsfavbj8PArxhBxGEZBNzha07Lc3/EqV9j787ZFXPrOaAzHkKVOiOqvaz5XzT
IqxNwMkCdwMqeqIFcLk9Hb7fyEzwAtDQyTCTFqHM5qdMs50zETRFJmbNVg2Vwyz4dWubALI5SME8
H2tI8HVXYR5wbMsNHQwL8aFamBopvZYP4JfTPhUAOINRnOeX1FTL54P3ManHvKw8AWDTVaior9US
vmWwm2PcZAx7hro7rxjDuXfq71I26cxzegvgSS9fhqZuxMagXksmwn8wJQQKu7fswJyY6Sh3fuhG
mAfyxI7xDOJzDIGuME8VlwLsuHv90DrCiXyyU8kmDcVSMivDTug4fqp5PX/BHkpnmBjgFXD/TThG
r+Fv1F6VEATIBPCHie5eNdOjzP60XH3t6/4Mi4u+leM45kAkE0cPkDUMzgStf/X1W8N3U7eoWmP5
HZJX4n3QpZ1Y1rOVuzlH2B4tsOUaK+RuKZh6vCbFRdRF1DBPiDX5cBQNH1SxEf5hf7I0P+cXGmzn
tr9/MDXuwEgpkgVaiJZJjv9eFwaXwPVvDKlZQE83zEZ8TRJJZe5kdmPlZtUm3GAZTH/zrtsEmNSp
TymVHIH0pQwh/zHZUVUddpeMnrvMXJEeMx/bgRNtSVieA84gxcsglCdfV8ou70cX9vTiqcHuxvut
bLr0ZEcWJzMkO9e677GZR/qlRGTQEucrKa7xcroMVYVS0mL0qAUrocahXlLiMhF3oqi8xBAlsiCz
YfAcQpQ8pLBakVzdlwkpfRC0Dh49+26qtWsTQQ/760CTuCoI9QubdBDj4gKQjn64yo0/qJOwkkTj
Q9grbXsNGwXsewURYWD6oLO4ugwXfUs5uahqk1CrnYhAnW90zxV+ym1aiZCyPvK0ODND9IvNWBa3
RsoC4Kx+F0e6WT2xOVuNtQtfO+shd0ZGVzHWZROLMU0P1HXwd+AuuFj+PXIbr4iCZJNCj7WB0opo
UoaZd/5ae+8wlw96UKLKhftEq+AimmEFRfVD8qTzFboCMT+K4JI40SyM7riFkwShBu2+dQlfLMUQ
szzcZrOEVXL7YAH3MUoQoxVxSF68VEAuCCFubFzdiEjz7yCZlPi9hEAu8lNU59L7rOUUy7im39Q4
Y5Ka3rSMTyGX1RDH1XJVe50VKP604BZv83T+vxQ2H37NKMO91ssWjPepj10k2oNFta2AcZLkr5eM
5+23X1D65Q8yHUlpKUIcZ9UHIlEE2wG5EYnhOr5uG7HyvJ6FV3+arZ2CcTTE/LgNW0TrcDqdkENV
i9kYJDf84Qr4NkT2thdm+WKip/of47IIr7y2Y3hJbXEwAJq2aCiLQRM2z9ygJaZrT/cIanpbVQqb
5usxeOgVSkIqvYjN0gkNePbgjBof/Ve0x/EfMlcWowv3lRwWLNwnLLNYca6QHD5V/Faea8FxkaiV
d/RLIf/iHklhGB4p6CcE5wpSA0BDjK/0xazSSrQL/vY9+B+CWpnhedAe2bu/DwHwYrR0XcTA40fu
QFQk28KTd2TWF+9BBUQ9echK8pTj/7tdrc4YjDquXiPruBudtSxM0ISy3w7uH6UwtuTHPJFlmoWz
9X/zemMo3oiNS8l/GemAB+UPpDFekpp7ddtxI6uruPge4KpOi8kZJv8SfLcpTWck5l+SH58z9mIU
rPYOs1Kad0U7BYM7PhfgxYdxtoZEcSETqKdpI5+YpWjcBctG2LeovZGdG3y/QW2tW2PkeEmTKely
eneM+4Q8XXXBwJFrAfgRdOfYBMbRwy2JRrWVtttctkq1hcojNVENVCV//I3PpR3yX5fpMfksuQ1f
rLcyE2AJ//0MJBdR53JIZ8lEgck1j1DMA70quGuiVl0ALwCj3wx2D1+k/cScAX9inL3/X7HXlgBK
0RQc0oqK8d4RrAgu/L6E9R78JN7hol+g6oaT+A5kqhm+Wc/7yAj7Lt2Og9afDGNU1LyekGxbhKZk
oaeXhTxgv4huuC5H4x2QaF9MZZevbQn/5ZPhHLP0Vp2rOY8d+nnzP8ROY374NQMjZnSFpFOX16Ra
tgESHEVZHD+rPnKcFrw41Pah6hJEj1N+vP4D2zfh5IBho9+UlQTYaeQB93Z4PJqZsAB9ihuFsmj9
8EJ/RasNOYwyiaewFbUoqKLCcLa6Iwj7GqicNWfYG6chEojcHYg38W497dOyRS9T/yutDSnTenul
tDQ05s67PIcMK+RMCNwCyETKufAVvFSk7aQXD94sCrxoGo/8OFC15b5h1tS8cm6Tyffjx7rdn+nd
WYFHd1Bd5WTvI+mgINroR8JN9l1AEI3dNKwuIIt1HF7mVdZrNhH7BbCOUl1Eh82Z9CTgA6SoIfF6
Q+y3P0g13Dj/qq+CbKpJkFodNqogyqI9w/iJij+1Ba96aVBVm+kIyFIAJoITHFHexlO0roH5mFqc
nhk1kkPwpvYrWOF1SXsqsaAPQJfJ42KtTbJXuP8z+gdOJwUDKCn3TIzd5zhr9E3ExBkyibFSQuWF
vM8oI8tOZie22fr+cnvFOXduW3447x9K8gOPOxyjdkoNfhGutdV+UWk18BWN8G436ygNJUrG6rZc
GKRzcErpDZKJjTlD0ebGKs8Gqu6Yj8l1gjbbx+Q8pSFAi7XpYjKxLyeAmyREqSHGO3svrVl7HTh+
2++xYlPTHmP3zem4N6E0kjceJlR0pUiTi1SfgOAq/J0lg14XzdofLbX22YzfRjFyCyz7ET90rG6U
AQJ8V/Eal1QKtEHh1vfu2pNiHy9+q71b256OCRMD0FDI3a+ElCTL/X6bNuGB1jQSkvnXNKLrGkwE
zszIizYNdCw9XGATy3DN4uVQ+TvNxAvXnpYyv4ouzzDO63E45Wogb5fJh3kyEiHvWsGZKhsIwqod
tfJPkNxRh/g01eYhJfZIq0Yf9fDvdMZlWoVe1m4BAFlYIFFacMfNC7qX/U3zBIDBcwM+xIb48GjK
tzfrqGgyo3pyHHHEL6pttm5qHbzlEQAJKb6aOnYUTBmeX/FiSlUZt2Ad8HLxKebFwwRWQdZgY5c8
gDNjMO11Oq4OonWXATSRAXVzo3qTpbFFNcr38ZNp/XOKyqGFUdZ/LRYALDtXwSvF92Vbkmt1QyLK
CEzck3JX0pGOzY8uShBXh4cwtrOR21EQSCBZna9iLzCF2OIzoY5u5h0aljtZ1GCGDiis0FKFKEqa
yf2V8KH3QcNbsYEfTlFRix21BSfSuZHsXeZorQneVrprtqmKMSQPaovbsJ0zQsHKHAV+Uodh7tum
jOtaUkGHnZ/xWEfe9NdNt5f6u8P0KpX0cxaHBb++Ed3l3MvhjP2uXmtOd3syHrT1BWoG4sqf8kv6
/KV419rQEEnC3w+7fW36yhRLAIYcDZvqs/lUohW5CFjUZjeat12XkKGvrCiW4Q/QhP3Gfl16rJvD
iXRHIX+ZwmZK2klBjZ7PdFq3z9N3kUjjnzFNbpCMzhk+If1TaTKuLBGB4Z33s8m39Lz4kBSZ88EB
urTkUN02H7DVTbAPtEA59LwDC3N6o31aPug3SKKWaeyEXl1es5Hh4ttjyl/D+BKGaFvruJV9pPlL
LAo5zP1V7MgbYbjbvsKZlnDkej+CGEYPTijWbYw6XZGFeu/Duq4ekHWBrdRPeUJczRYBlkh//T4N
94CZYYQugKrIvMgk/Bc0dP0EZs48rT4DsaAVszOTorED3QxNISueIFEzn5BaHPhzekl4be1Zcr6o
dcQn+I3tel8mixjx379mta7crPt0Br8ivT0xOWc3vV9nfGkFz1DRIHp68eeaqp3ijlMn92YxY9Sj
Sxd3MqNzBI+gok34FkB1iT4kUKq5o0OId8fyO0TrqFEYXbX6mICkdLN6Ab9HfXhQOzi7+dmLmY6u
cNUc47fhJLqpj9pT1n+hgo/wmoMcO3+QUq61Myq+hLp7WtQkGJIW7t0ukMheby0JY4Nvu4VSofYc
qDvxiX3vz8UhalEJUmR8ovBAVYGW4q1FzE1QNKCNBv3lcU43KGsIQWuUf2/tRelP/VHEDas8Tuun
YmwC3WG32aKVc1hCkrXI7OGmkrVEcg3KmuB6r4LBgZnFCtWsG/IKQZ47mc057XV7t0VLxoXQR4/+
n80yrFwN7tIgdHyzDicOFBsaXVgtP1bOmLVZea8Sdb0M0nUGHyRzB588OO7aHPDdlP1/e5RNgGvn
r1AAUH6pnWrzWGrCD4d1cllyqRyDcmSYpXppKSxWFzW76lQlkB6oXI6wahTLJufHfcllnaU3NnJG
Goxrc0/HHS4pxaJPgVLs8hSaEHshvJTQlh1HwDTQcs9jQxnkA07kPd1Vt2PeT0do+3AssWkg/gDJ
SE8tdVgM0pguIUqDvVSdLd8PyzW0lKKOZ6LIiUJ4Dwm97NiWfkmhnqiWvsEGh5UyCJ/E2pgW3NmN
xlunFrxQJihzgI7SvPkDIGUAWuqEQ78qUGT4VASni1WDUZuwSC8wkMHzDFRoJlDbZyBgqKPvtwnh
CAuWc/ySl4Pv8yhTXk6lKg/7WEYQCNUzfKS6d3PjhyAqS1aojBFEFLW4SZEffYFnvQPXK1VbbnDG
jR1cfv/ikN74E6h32mXmo0WbsX6S6Yl3YOPU7spj80VYhCLlm+0b5KniiQjtmJ29JNcAd232PZNE
cFr02NYva91za2ZUkP2SFuSyCIror5fhSYXg/n4Ob/UXD9hNWXcfwvl5CLx9QlsLmE70qU/rN5iH
QGaa/dknw0AF1xAQOxwZISVMTVUuTF5zAMoQarbnWQWV8KTlYW6NXxvcrdoqLUE21e7D4JZB3VsM
p1+d0UcQiQ21TLBbYfyZsqUbzvGxkpgcSgIPwxvxffZCDXVAT9h6iJvvwzBXiFk9rE3GHDR4AVgp
3XntjBoCmSgxLCfntdNYN8qFO5g0E0lCABy0k1H0rRFYnymsheDsCOXT3RlQzRmtVqlifJiugTaW
KQHqX4BpbpFXN8tHAriCrd8G6yQIOSXTdt4PpiNxQ9KM8+K2OtmrID40Z2LtGHzhjoCjo6U+GDXk
9fm5HD2OcGA7z7a9KbEvIEGMHTZZhfi20zWLgtXOGL1fdFNyveemC1K+sYoDI4QtUS8UWLB9vbqN
wBTp2TOSyj9VI6yOvENbfopTzDXMafRGj7k/TWVbHsljc4LtMDwtynwtaUcxw15aw0Ylvo553iUO
omneJ32EM4c8TSsYTKK/ZF2OT4jn0zrqd5UdynzJyXY9ss9h/HFOdnAi3PxoYKYp1Dqel1yMyfYB
x8BQNvhJJDql4BvpnmtpZynniWnOIjymDOsVoH/YZPIHznsUo2fIyutAQ8LQ6StuTpGao0XLb7aL
FDVPOtP1lX4+n9aIhcKWX+yAzKchg3KsoBmqn+dGQxFr73+aWK4ybAtnLluF+if6PbbtDOLrench
YWqGZ55G5UJikmLnoppxI7cKSwUpdseVYvWIx4gyi4tn2D9G7F5X/2GWSTg+FLy7NXPWqkf9R2Gn
c0i2SiF1mfx+S42nnPKtSFI5AD6TvBO5xN2IoFhvMAPHE1VHP/6O96v+ELGz56iThn4WgP0b5qC2
V1J+jGeHv72oA+wc2Ci28DMud9l4R0N9Exwkx04p5Gpja5RdGo8HYfOjZTqgrkA7r8WG3hAh7ndk
rodizXRHeFSJFPy2UU6/emKocu4bjv7lZxgE/2gcfbjQzDElQO5Su16mgX/cgWwnNBnuQXNDF2il
6Vnbcq88RLLBCDjOVWjajcXoGnSPQai1pCIk88qjaacjgYE4vigcnr00bqs1JuMW9T1pMihZkMAI
J8Cj0HTZ7ut1HOqrnv91D4H2Ppq7XMuDyqjCYQilzOgPaOPZYXZzK2bUBBmEmIiJAD7uMDPzOdlG
MfgchXc2qzT/J3tF9P06CfIxmRhPRGlSJJ8PYCif2RXRc1x7eBqcZnF1+j16h4ZrSbJvJyaH2FyH
Ln45f+E0YDDpS7SF04wfc2qHGJNfXHKPMYEpTP3kWBhQoZx+FFTyrHETa7jBkEvjyC4CMP2QXfPu
uqerNcP7jgyyCPiHwNuQlI+pzH7z98fRi0snUB/dAHqnF1wpnt01S5L5v6vQxNz0hihcoPMciJyw
ODt4BzPH3DLhfV3RpTl1SmnUJn44fKMb0Xdeow0gak0s37O4U3ozgbFyUVqulfgIB79AJZnqfsS2
Y+Z/qmK5iXT8mnJ5Mz5b6SGQQbqNAtZiKEs7UXRWMEKS7KmP8gsRtRns8X4k1747olazwwqOkxiB
WzO2ee2gyKnWySWkqvErnpNeWRDvA3c+cl1vVtF5cvrGtRkID5pHuaqECfSEcZ/QcfDoM6hga5v6
uXHbkiXp6Pg9vJHGedwx8dayIFkg1PNGiyzoeRhj5FxuyUPnH2PtBCxXVxvGXe0SesLSgQAmxjBr
c+9nUTRJO65RUsNjcrA6tyDuEcCZzteLm2hPfaSmG3AXRyzUyWtN0FmlAQoDcRKjNaDL1h9jaO4J
GlWCr3JLmCKfVDMfB4JoMgaNbmkh0+/JVFf3Y/xw/pZW6x90abT0eNvkjZuA4wEciFuNzHfD06ww
IQwoMfVAQNlQD3jsqEdW0dssQiorOWEl6Cc+ttQO4NI0gzX+aVRpNlVUY6QSOGVx6WxbEdFsTAyW
1OkXYEikD60dkPnNLMcXPs8yNuoxsWNgBA76SAfezcDGoB6qhcKB8wikfec2Poj4bTFtEeEEkfQC
Q5BGJFf+Y4msqQSeTJm8Wg2uC7xphxOxuqlMlUdK1XhDog1Eb0tu2DoA+gNqNidiH6RCX495wK8i
IxjYCDVoqR6+1nag17sY1wp3JjehLHdSeKEofwtfqwDmBkIs2o8tnJiRCav2a+WR98pigag7B3o8
nZlRuuqmJsrWUTBvmqOhBS6dtx01TGzSPRIja5mZWgCBRP8lyZWkr3wZp5HIaXMsD8XuioCJWTDU
kmy9IsWLRr/ByZt5W8DFcFawlXN030bTkKweitce3Kc7l7dNBsW5QFjfzL2vgEt2qTsAzfkOr0sk
h9YM49UD1pb0zq5p115alu23weFUPm3WYer3T9OWdKzbuUJjzP0E3lZTjkpzxsyquhl176YQb9H0
419SC1zsBnqpju8jvF0zBS8bEH3PRe70kFXOM23biJ2mRXZvCEyXXRJHQ/b/TkIMmyHYXNFRTM15
zxvT0oDwtRuAQ47ojMpdR2KLveqZX5g7UI8Jq8IbZt0PQhLdn+fuDTX2OuLOEsl0BZsT8RzV7Wev
kfXmv5+ykMY7P1lsTM+UiitqV2030O4ymfygXMVV85w/DUAGL0q5WWFZUWywrp8mn2cTj1K4p8u7
SftZLgCBnHyyEdm1KqV9p5uVXqCmuTVBA98F3AMF2O7EuoMtiH8cDrGOlzPJIEzGOV4u7Lnk53ph
Z3KrzpnoveUtUUImCN684/qm5vtT0tkWzU2JzKxkxE52oks9GN2EN0JqyuubtLlDh1R2FiHI9NPb
X4bLY9StBPM5AR7+Cc+XMQjv4bhzM3m3p1hiID8BA96bpK6tUcJDq21sxiYokOu/PCWmHjQdlCZS
fkvX9XEcZe4jEnydMye3o58kVdbXdukvB9giEQAfm1WERVO3d3GcDzPlD9SfVgWe4BStsHJv2tPk
DCoz9p9LR3GP71l2imFzJePNPwhI+wz6bbyD4766aZcM3GPbgKIGqTGd/yX06IVYdzcGQmF809ve
JFYomZm3LsdjioinCcRVkMGz7OHks9JWNO/6rD91FATTIv0sOlkcd/EReSsStYKsv4SxSFvfiFKt
CmuJmokthr5ckXMK8rUECY/dHvBd/MHP1kF04TeJD5qO4OB4fBQWmroLvagJUhU1m7qazREojvhP
tzwVLADgjYkEQU5/CMnzc1Sk/7XuI728TxY0sjGdCYT97SZAJtPNp+ypHmNC9QWspyGPysLiV9Wj
veFqrVgFRgpZ5ZxXfRvD/1hUlGo6WZGZVo67XXD2o5fjOIfuo8swR32O23PsX66SVzaCgaeB7DWI
tbPIkI9qJaOxEtMClXi2YTWYAhS3QgDBMOkL6RJ502da6FyYiHf2f5P7jjNaqPGgv80szQ8unc9q
KfeLPnjNqYrbtHpv2gqlWbdMMBCY7vKPTArKZWonpVp5vC3FyGDqHwtvpaGVjLmpIpTFEgsaj0Cb
3q0siLd10Xik9jD0OrEMo3HIGIxoCsJXeftXrUWWMmY3yMW3SHRF1+nMGG06JAookjb6/AacliFF
89PD0fe9n8IwRhPrir0L1oOI2wHEh7N9iwVttIo25UOm5olNx5VfqCxOEEc4nvqwuJvSnUjptXyO
g5lxjCT17VtxMZI6Yd2847ntQJekXdWC+/zab7OaNZtmBeKle8XhgZT8aqP/4FWf8Vx2/9+2W+jd
Qn3usWdK7Z5OH0URowHMK91clSF96hE5Uv7IT8Ti9fHlErOMwD1gTqBGIwR0n0q6TTjSTRy03beM
kTOLi3y1dmYWzyHktEgPfORYAp/ixibXMD9wo7bmg/JR+P2zvJYOTZGIeSXTlLPS1CsV4qpf+BuN
qxEL/lO7A8CYH3K9+IJtQNybJE7lDHRRi/PcEojJWXX7v9cVAjRzo90qbi3BAIjUyb4dcJjr9JbN
29P5xJzozNyTlRuVJ3+9KsOoosvNFDnfMC9ovR0cnImbcuwW5qfo9Nnb3bj1C/fRoG2XKUegMzjz
dU1vEHIky692b3KSNIm7YBAn15T76ZbI5TzK2L6wA1bz5lGUKwARMLDbtuHN/1EMYhQolsQiXHaC
om/SDHngCwfvHfklVfMwaMLJL2QKhQVuoG0QlHFukoCsU0T+HSRHoseA80ZrYEOgNNE5hRilHZWj
OZ+BKMx32dL6BAwZo4BN/t+H9TFTZAy7YCAamdqtCLa80g31d01bY+0wQxoTIRhtiuPfRbLXHtdT
qUln8t6cKKjqIukzLxzQdPCQv5FenWgIqPZkStMTuCG8h4jxVG1yyR4lwiZM9540j3+GUtx+OSbW
qyjPDztQsB/XPDqJOoGE8kWqWLx05gYbRsd+vkJUbskUBQR7CMFjyX3wkZmF/W3ciJ2U7YTxuSMi
v8Isv5m+dCdOuzxnD1LRYoJesHdobYofJEs1fiH3SGtano1vxy7mo4hQ2VARJmrUHisvBJR3yIns
15sDlyKcZ4U2dSv4OimwG1pT9qjsS/tbFqi36OzLyMvIIqd2GbAMRaGIgO72tUHGF7mNu7MH7Vfw
u8/kG9bdd+At8zgtq4upv4NvfXzoZK9rCbi/ls6rU4vXsEdFW6Scz2JLguj83oEawUl52gytgH1s
OkXIFus3runQBAH7PIgOCBk61Gwl47Gy/jmtR/6rUbtj4G2sZSIdBsgzvribMZJ4meSd9h0wHpyL
QvPjBoZKUOAo5po3imtLybVUl36Ao/GdvCtEeLMvrMjzekKmL82qar2sfPywEPntYeF5CN2kI/RW
/Ha/eIHzfSzD19jOQ+vsn90m8vy/8g7b3Suu1VL2ziFJmmFIkl1tgHcuoKkN9gWPNz7B/N3FQAai
75d6j9NpMCyHGIqWqnduD0bB7wpBi2AXK/9SXCsZ2r5brJ9kNhj0wH4Tjfaxr5STom8Izh+D6Scz
GEmJMaBMHb6ikajxYz9IV7UcH0jCJn6J/39+NrCJv3251fsojIMxXn0Mc7rlx2MV9g3OtUV809vM
oC4Mb3N8ETxcgty98H2t1S6PJSpyRCu9/eKQ1P0VB5BF46aZkkog3BtvRBb6ioVftj0lG+zPFiLS
0QR8ZVqAREHEXPwbATpt9wgkGlseKgqk11wHa+RqjDFvQFJt8oio7z4rZi/RYzbpsi1NXpvBHWHM
R+NIa6J7PUlxjBGTxamBU8DU8oXcV69ahOhzw60i9sKI+BvZt19T6fk4YXGwCv3ZylltYMzXu22s
ofsnu700O/kbL0LYenx53cwINzIAT7vz1vuoGutgt8qtU4uDHilj03nHqALLpcszikmIUYGAZj2L
DEUv0L6OTs9Exiuc9iaQE9A8l6pthCWKXJyPqikXJAnpATYr7gnCgKMYoqAsoBVdUt0WkYvP6zW+
04f4tkFG/K4zhe411EiQjLX4RwDq6BjZs6C00uAa7zTTFueqZjdgvcnuSumh2UrU0XqQnFjLSd1H
Bv9db7Aj6s7HBULNb86SixCt4tn2PUdCgzhteximGIwggOoOhWgr4gboK3OaWBKb0iqtQTEVH7wf
i3zK7kYmBQTGVOcm7SgLTUZzsmy1hh/qnIwV/LGV1Jrwbw748Ho/thl2+d+zM2OCLeabU1+N9rMr
FWt/6wGB/kQ87jrlCIF8JkQxnyMmLAf9mLX+xhsab9Cgw/f5inUNW0P+QbJuS5HFyquRwXX2TYJY
q0mRAvdfdThY11xmDj6p1+hxQIhvIc4FSEI4Spq1eL8rB+JvzjHrAH8VUokGi9vZ79YOusmnU4Jf
hjapINfjq47M2ekHG3PaeYJUtiRIVb9eVgAzcnQLMXmk9ingdtnes2bylxQZ9kbe/hqWN2TVyUEo
q3zEZE8hpPi5MQ85igAbT7LNYgQkpgrv+PZL9ZLbGG+IPi45swkiGOhbbHH15c9sMdIZ3XWOUyJ+
miyAP3YcG2TEzmgtES6NBaXntOFCmv6TXqbniwkNsKaaZw50bYsiV+Vi9h3FyapLQGMl8tLaE93u
kjyF9hGsw1l8PNpNB/3JUNZXv8ZouiSFjOn10Am8YzX5tHAFD25hVHExb9+u5gGF++IrkhV09t/F
orTKsspe+imlg/BasPTrO/tVCSWfL7pplGzHOnR46Ee/WIUWVOA++28+SV/Au+g6GmedlVwjrUrD
JxjkAeYmhJAnW4w9iY4Bp3x9wmtuDKmdAuXrdkqvDNfN1XtG+O6h6intTLb5Hg23DlH2ANqxmhN2
MuPAsKNEDQCHnNjdd6YC620CoTByH/B8538smEqCfu5+obFGJG90os//IqIq0UOfRKysciVCGlpo
SpIRb5CC0qu095ps1ttErwjoCWqg/4NaizSl78EuH77QmEFO6PciZ6dPmUNrgtnF78FD1Em76d9g
cefIrddWdZYQMr1p2lI0yMXSqEJ+74d7y6+WHsGMnaJZtT1Q6nrd3SuwUHu0/PlPTClcgaVjNhsx
KiJL26azZezdsgIiwcRq4sAj+oJmkrymrqwdmUxVYyqrY+bLt1zbzhcON5EPpmQ10B9R3R9LIvGQ
rDkX0j9yfmhqIT98ywIZ6fxWYJ/bEjqQaSS0a2cv2IeKlsmWBC9YAJs+7MxqIBvNLE8moEjcc8PW
jNI6P2oQhpZXQtkEww2FOavGFPZNwB0N44N8jFScT5o2G9JbaJrmEfK1whX6NrUjco3dN1pRa6Be
S1kNC9c+BqTITbet5zOOJNY2kAELPnDS4b7/q+QSJQ3SidV+5beWEElAIAMQtFLvhoOJ/2sombOf
qcFox2fEzQWaZEsCD07xq8R5+OvjM92aduc974njuYA/CLt5toctzWKmhjs+xKQsNUU17e1oP6B7
oLsDWvmXL6OWTlMCL873W81WIiufu6h9VbhZnyN3YF53F5mJqDJdfChRYBufUsfzMjUCHt66CkVs
REspOUhMGs9Fik+YwGVcCa7XU1HfHddQbDK4pRMBR0FVMmoFk/LBVAflKC8Ufe67/IPLooYR1fp1
feMuFmOfb6PCeC44oLScUoHpowx0GeFOLmzcjkuSXLfjt0P60JUWfY1/cQ1OmRaATYldOBzYJcsI
2Kc/OVgX0jswlC1oupjSjST+A5AJ/0U+ZaWD28GaJjeuXhW62du2gk5Kqu+MZox2WCTNOCacLhyV
OgU2fgFz9GvGW47soR0Efqk3VTtOaS/fsoI4mKdujw1BHjsIw6mvvPXfWyfEzngVOJcNKszoevpD
/8QgspsHP2YZCHg4eirVpdhaQVCDG8G1NOJX6XblYun3MxxEfXjElVEnMKep1lIAL8mrDD5M/bIF
iQRYCo0O4UHbOnh2NrqENm8JwVwMgtNBge30uzwK4GTSKNxkFjFR3DPxAICdK93INq11TVsPGxCS
LJesDqOywCvdbZ4a4YcPLhioeRA22/sSX6w7OyaEDJK+L9brTHISG1k9QQAzTULFe6+JoDYj4Z8I
1o8KaqPif7rMAumn9Ao/Ydd8zo6KFvEWfJM8GW3lEe/AVokWERuP57zDHa4wp790hSyV2cK7fGYB
gU+VS4HDTFVTYoObgYDzz0gzBW5dKUMg0XMLSfH4WYSdAvve6sC+vcnWn41ruB+lxL1St8b3ROjI
9OCpEkWdm+3E/RfdsiE2Rv7QF1OGo0B6TVNVZEj7wOqaT5jehyLc+9WPDhdxUdihIOF7WRwUAvB6
3GL3tuXBcn5mH/Cff6BBFbJl2677KkxB6MvEBi7XoA0pAN4wGWASixLeIFaaFvOcXlRNMiN/nPY4
yWPqgfgncezTHUXBIHr8NzBfRh2XTkJ2Vl3+nSB8oaK+M40JR1jdo06DdwIHMbo0OCtOM+6DWsZw
URH1Ygv+LOMEeTFouZxhMgRd+HhtkUv+90g+xM7gh0Vt0Qp24HWfnKAb317nQxAgzgS3iC7g0JT2
DV/nuCrUbih3Rd+q1pzuQ1Vz+0rl+a+qwLLY4+lkrsTyafmTw+KmtIbYtfD6C40s1iA/brYZA5zi
GjfQ7qN0kJfIAjjKhOmhai8zcZaLi03Fn1mbkdQV5313xIc+B3AmJpX1yOFIn9wVaS/cd3hwfsHe
0JmLtkoGXCvvK7QXErfAHqBuIUP4/atESza7OjR7Tpk9R4baZZFC+s4JRvqzd2JVnpDOhVTWD5l0
6g0k+sQpZ8HR9wbauL6Qnn8nMwLETq9OUCb+txoLGdA9H4FJoDhQM9OFQYprxdlm2nHfjhTinLLC
QI9U7Kn0G+VXXCG/EhB/ut79zCOo/3Wa+0X3N3q6mHEXwgr15WQZL7bgN3DogSMp7ozXRnz3Hytn
GOqIFO0Z9NjT36cnQyl30SnkdkNX8zThdxOANUwtwTDFgJCwdyi7wAwPJ5zs0G/LDJcqB/DUcTUB
8GyccrKPse7nNjblfhMhONyiNK7b+QO/bVQxQerMsLpatxXR/s5GItx4NdEf6dZetb3w4q2TWCg2
HI4eqbiFIfRVifPH1oC3k0T2bbEbKOB3rp4lecRwAwoTjHrGGNCUTKaW2HvR2XPk4QrcZjO1lK0t
dOgmZw0ey7CeH8QXALQ8eA36TjQI2iLrLlQHgEZBn0g17p4yJAWT66qVMFk55SSvjjcRNZLBUE84
cwWpV8LqoWQDpJH3D8r0dImibGNmJ5z7D+Z+iaXZ4R2+BGsS12SDt8VNZ3ZnMm0gCjR2n6vbcyXT
1ia3nZCq16tp8HsxOXcEA2jOwNif05GCjBIJ6pflLwBFThbttp5RVg+jSPkUQ8xua1lXuDMEVTpn
wVjP1Zn6FGAVS2e+zVlBLihVfqhJfelQd0N8VFJDuz0G3/dD6l7M8jAgcpSvq7mC3jO2/mwY6g2s
jRYnaxJ/qwho5024+i/tDFVm1DVfQuPPYKLNpZr/FkhVjovWby/SbT345aDSN0yPo5uUfRfBTEjH
JfIif1xdrrMB94azKdxPi+YQ5Lypfs1LazWgAQcDX1qaFaRPuEe/tgNZ6wkFe4MhDuMPNk7/1pVE
kMmvppv4dulK5SQPWNanQOQTt7kexHFZ6bluSpNQ34JeXu16OtRczRo7djvFDjvqlqkuC+ThXCAo
fw/pAZCSRKEKOHWyqI/j8VIT+UDxeTx0zZTG6LuF4+1jtE0TSLOA3onf9+/gWaWTFDayVXvMXZtw
3TPUaxy3FRcWgJyP7LWe3rNql2fushinfDTYAFJl825+bksb4DkjcxVU5jRoy6tphBY0/zDDx9Zk
sKGQYjPVrmVRdQ2MfCNOxCl6bh+LwTmL8pwac2MbtZ/7KWEXfu/FXHnmgI1dPlAWZivlcDzN+TRD
+xBCbUbxAHGye2HUdSkaUr1Gp7TAYQqHEs63l11i3s3oHaFMBs8YRnzwEFnKpANJKyzDyBIDZEYd
/ha6TYrQIq4wUq9/5jM1fM99VR9WIxDpdTokqPA72Bm8OEmQD2UT4Z8qTzbqwM8kgY5RyFqCZjVh
Rda4KqXou863zig6+rf45ldU2o/Y/hz7n0xwrEe1xGwQZL5OKX+kDTEdUhIlj5cdVnlf5Tr3xrew
V9X+5KfFFyT1luuA1nwtiQGVgZUxHrpj0MM4PMJ+C46EoiIZReLmDmReJjrcYsAIpFFXt0Fol/2o
dERXW4UP7Ys/Qd0WvEi/IE0/m8hIi7+Pi/4Q7CanFvCXXm2TyirhK2zKk6T8XJPJbaOzEPazb/CA
5QzOP3cdTG8gAMoeWegGybznCOSD5yr/mTOUug1R5Zphs1z+zZuOtB+mnfCb130BjZ6Tel7bWT1a
GUlJQVSBYRcan1NZRnZXBgc+DhmuneM7KS2tMt8aEWMNpt/Fx97DLfTTl7+J1kvkG/32uI6KxKoX
TPnssLr884z5S8hgQumJnrj/ZWDjnwIBWsH2n+vx+PcAonjFdGCKosCBJyw/nAXh0P/pFAFMJddy
NIE+thXq2v7p+Q9k5GV7U1Iatd5zWDL/McH2WKhK7K3JQmWGPhF7YMX85miXqJ71T9CvFjcWTscE
DHFefB9addKG7waCNZMTWu5S2Bw73h7kLKTgS5129DOs3DFQb1sD7BTc7g2FmH/mEUy81TDkrMGL
mOic4P1pj2d8UwIJ21y/458weUeh29isk3dUaYc8Zwa+i0HPc3TPIacUwX1KNWHr2bSgQ5q+kjlw
kBedt4Mp+ssKfD07jCZlxeUwfSilQWrtXoSK/ystplCD7NAhIZjBKsZyUITzx8bM0Bp0900JdIVb
1eP7k+pwwyXWwAizYgI3gl6Kmj+AIEcWpKU6Kaw7Asrg84vFEE5D4zLDwUcGSjueJlzU9fQyKc91
nnvXgcb67C22Qh9KIXe9YGJcJU6cDBNSrELA2qmaimuanM9TzK5IeNHYS8UkqStCSxKOi/STDUtL
p7Xyhlg3m1THJ9dK8lL+72Wy8Cu2Rz52cf3hP3Oq6j1wlM+f4SqbVMfGUxoTs89Lc3U+EMvXeXD2
vE0CbXwYM5GiVAas8eEtU6c3CZGlVePOi5xsHr9mDWlJIHklXdCHFzK80XOFR+Tyx9A+Bhel57wD
Ac6BvrIFF0FB2J2R6yJUTDHaz7UqR6zmyw9tWYdYHkNtHK3gO8kCzOvQC38aSnGtsyfQuqx1wfDX
bV7cMfyGP0ePrpvTO781VgwVCmiVFq7XdF7t+WLIxBDpnr3d8qW93VimA7LesoEixNX3zyOjxkt5
5xoBfxd/3OmQWRq0CUqyOxOiaksHfJi/MWDDutiLD/9v+rTsFN7V8sxo+KrsXaFdW3gw4iepQzy4
TvBEPs/McwBxCUqNt3Xvg1ubM8gsgM3Ydt1CUII4Et+FL4HKF4YIH8rZP4wfl84xTn7pKz8lzRZX
4XIwp/YkynFBAy1Z3ahMwLylXZZ5jEI+0qMmE+Wzq33/0dy9p/6bbUBOlImz3aDAXYhmx9TML7ef
faJpevAzKNkVLe34j7AT/elQ1QaD0+xvnjeFVsQkr08vH97WyN6KTMPZtcp64OpMm9TpOPiP/YXt
Ac0cwnL1TDCTgHA9AMVpJGy/+EmfKqN2Pxpidsp/W/EO30lj4QYou69Gx0Hkr3x44AMEd+VCqJ1O
q11cEM5AvdAQu1S9E+7Bsn251tjjRqrQFieIb298UKagdSYJmIiAJoqboFTmCHycZYaazDbfsnjn
GDHZo1nDh2vH7CNyqj1t3Pxk89m2OL73S+KajSSCm98WekKukJzMJr2OiaagbfcUhcSxjAuWFAAg
n4v7P7ZI/AukDs+Uy2/HQL2E/x3JCrMX3jciekYHuS1lc01xbFqF1pxEUudQI4b9KEiDnkRAhzSr
awFM+fVY+L4VAq3rwdVoB4TAGjil3aOvtgT2bRZIE6xHhUJ7TLobLuwOjeFqlyw896/bCLn1nOYT
fyfDBk743j+DZ/b8BJ2REgyyhCA2WBFgKO2RKBtLlo/Jm4yVupS+FqDVKX5mio65f3Sw4piNn8DS
uhJA1nuTFXU5iUoKZwguFhaNL5HqoKeuNKW5YfFYazly8pqLQ7L4VfAg4Se3bfuh087MFuFkRJ/+
qbzUxcSTKToptv77jl1aVqJJalOE1lE2D201asOlNN6CF6q1W9QV6nU1z5tNW+mkeSgDywm5C41+
hHtms/PIPGWXkbv0tSZDmLdWRY7J4K2PxbVjwLZ1yxbOZ83EWTNdnSEW7xxmT+f5QH5EOj+BJfPM
RAihe5Bo1n5ikb2+uJW+2LkboH1DQyFWs3l5P8Bz/1YOsy3FhctAMDQcnUv3NFTFk3Em4u1AOVAy
9cDAuVlawvx/lmt6OuSEvTGc2EuDUPvMzBvOjvi+jKeFczv4TRGHl97y9/3rRJR3sX/llxleh5vC
HQuNWOqJ55vxLBB9qJ861OoM+9sAta/zqtCYl1fs0+0iuZGpB2ZTgPomF4M4Gg01yTuFWjqAheTu
b7fmXgg/E9C25IR8b1XkI0UxVqXw+N1sNni447J/h7Q6dJ80zOJxsiNjZgewI4iDPAHxUqzw3+8l
ka2j1YHxuIuMmMpC+ptU6ZKuujjpILaKwsmdkit68mFQ9n/vC14BXWp3Z2UX3vQEURs4qCUlFpfx
is6/5nWC3QN290MAi1SOu9T05ET6/29PyPu2pKzBu5QaaLiqHWSjVtfXl+ScAoNUBPT/VWlqD6Os
QeYenCvzgIl9snfWx9JS8Pw2fTvxzJQvmssq5RXfNGScBAwPzk23RPBrpBdXf1wyY2P4Rzm7bSF4
J3wZz+AOmr1jS1cDxPMsmmf8P/YvpyQ62xGUYSOGhSA874vXHJ/+QaTammzyScU7fsfidZ6Hjh8H
9ukdEzN7jyPLpzZMwfZgkMWh0c/WrawqpBVRgyLWr1fieDXXNJ22wONHZQ4v7u0ssW/ZXActwA8t
yZYffyojoXGrXjkCBicWPsmcMIoa7Jo89AaUtTuPMpUxvfvoyHq8xZDZ5xBoSZGK0CsoM8jFJgJv
Gbnmmv79xrve79rrxVPnr9POKfYKWxAPUqHCdYdOAEZFCQTwuH+HT/yQqM4uXJ1zDalCuEAXl/M0
kRiMX5ShwPdLQImwVewJs8q0eE07SJaUPEaadYMfWz5g558aw4N/Lx9dpu8JnHhKrhZD8tyY4uki
V3NzZaSV1QqsQb32nJwhQTDoseuUHzYzR7ehO4LPoYk/2Hwx7RztbK+dlmS2dH6gVfCv96mSbyLs
zPcnAaZlVn0fLF+q6x6aYY3oLTke6MylHm7aBamsELLf5+iYj7DnEcJRTil6T4doozNFPO91Ibxm
YJC1idMMF5CdZhsuk8CWZND00PEiNBMe6d97ZkqYvNuUzZAoMo6dSaaGQ3I8RGg7Wtb39WgzUa13
NQg+i7iicH1ta6oGwc/6D6IXtFcC+WwVRsvKOleVqs6T7lnfqXGY+0JXQ6IjAs5Habk3lJPPxmb4
MEEfFsSCZkWJvQMIeq62TOeFhnQsU5pEk2odAmADz26W3aIEl5XVZpMpd15+CZNSlla7oFQVz+U6
UKCA/ElBHvcRk59QP6eLJCwfl6V9XStYr2+A554nUWkCgLy/ANGm3La6D/AWYgEyaskhHGamkCO8
vkWHI1XnIfvxp2zku6RGf527gx325uFkZRqMN1YXXBX30LJ5mJKhH+YVyK3g2TRPAUK3XK9h/X95
x66I0P9/TadPa2ut/syRa42eIArRZVZQyF5nls+B3LBiHQkQou4g9LVBtsUYP+tHstGeL97w6tUs
yV28DrRVOQb4RGYXeJ1x84v09vwbjQmjbaPY5/HKWZSUCBL73aqSWxyO75ssGO0GZbNY7blJY7Dt
HbnkdBjF6wpb2ytvxHUVDcpNKm1juzYwJqFQZd0JGShr4mhw1IfuI8kwcqMrhsNLGHnButljRTXo
BgTLqgAbqWuw3fKXe5KAvNorkMzp1t2z8m7wRGJLx+kleEPq/+Y5QMXb1FNgFuVma3EIDba6yN/J
AYkvEEY1hg46r4LOadB/nNKydnSCLJLy9tOzhwjl7w3AmcNFbG5AwnX7ELP+6Ba4imjSTl1vFvxF
A2xpVSOpDwpmanOBvRTkrFAv7mvy/U/u2rLnrLB0hwW3XgZLfzlEAm/R1GoNIqoIDs2Vaeu5VomV
cQmcoFhgwd5B51p7ChLsZTY9QQZVBWh+q+zM3rH4YgwEtNrOJGwFyYLJ/Y7P3Jr+qlvrPwhRbEjM
qo9sPowOohwX+XjK9J2GcqdR/vKfi/lbvYxPWqaTmhY+lawXph1WnJbGXlEk1HugLPuJac4xsca8
Z+6ez77UXl24eRm6TLPCN1po1cUJA8BQwN3ICL0uC4cOdaJnUnFJxCi/lUbkTVnhWrTo1jAbXSA0
snR1MptsuvDHSMv3AUfCGd+d4SvEKRsbxdi8B1KPIpoXGHWrm1MAZQLFGmDuNivJ0QCsoD/eHOod
no5QcV0F5jIppHiBP0QdiLIUTYW1R2jPcsR8DJW1Wk6EUemlR++EiepJ286SAQikCJ4iAQUD9DPH
Jg20xUqrnJFBPQLZ+RT1m4Hx5xP0PsDzxJLI/bi8j/be8NOHm4cvjyWDBu4iWP21Jg1+7hAikdP7
oaAQl4Quqyl08NUci0OeADJKptDGtdYG70JAFRt3aJCU404O7brnoMB+tbJ4QAgvo4wWLNT3YcKS
t7T2ZLTSXCvbzoF6YXcoCjam5VhGnb1ejA/SRapmuehleIPCFoXP5RiSSFxVFYKTbLv2F07YiuDO
v8532x2GalxipHtuQlFSe6tbbn/ow47+wFtdpd/0OZXH3imdiZltjM0p5n6KcKuwFSupRQZV70lO
09//B9rqrfSmGF84XMMBRNydcZejttlWYihddiqHp63aWZlqwLWtqZcQknTj7gwlIqX8sU7oFU3N
C53pqXADbyxG+fajcCsBTiMp989ZelqSc7KQAu5Yv7FYFthYdo8qR2UOhp7Vk8831Opd0VVlbUJp
sIpRObA54NQpyNxREvcYKnG1AYno6DE5/QoW3jH0+4ki0Ct2iPBcc/G1SkoYH/2iyQZ047sZNeCu
Rvrg4NcZ0E6HtfeYNPqqUcwD1SrZcoG2FqujpUSAP0xoxrIZoS384tTR7EMi7jyboRGajcivIwWT
rB5ces6DPISuKMDnPsdZvDvddSVjX3ih9yhOsOobXc+kNfj5l8j6A5rZZogzGTZBZGpXW3zrf1m0
w7g+KJwpx6ytNU0s8L5cNsq/gPA3S1PhHay+AflaxuA40nMF3CS+uZm0uYmdSH1QfEs8FZlgLI/y
GPBBc46S+ArLJktY0FQ8BXzz/OjnjCCEwqtUqgibfGyNLIYTsbytAKrML+Z/8pC9vaFuyquYdTwC
9/rshXanIW/8eX9EEt3m1Q2eLrRaFgAMpKVOWj5r21mZJDAZMeJ3uPoEUog7LxJGCDrNi2TFc0UB
0drMh+1tPgqFZ+lc5nU+3ISb7CsFFGotI2k6pRawChPWLVRCFGhBTEuVbLFjD+nU37TktaUibKs4
3CYLInYrsG32a8/NfbXLSU4jlkPo0QUvac9r4WZMFgEsyh1n7ZdDXbJOxOTXXmuPVQ5nPfTSs8it
c+H7fqg3K7rX3Jf0v/nyFWHg285001QxbroIsQ5fgu16a6VhqpYOoxJxY4wsk9OZIZOYPwUDnrFW
QHIXBVQdXpZnG8fnyYwUXqSKXRu0gmFQskKoK2gpZR9468rrhh80A4z8RJq+WSE7Jmt+2/JxJOQp
jR3Mnfesj4O6G2aVyisVNHNSjo0hNhqIZO5ACUwogKwzHM26fO5a2IPx07lOW3XKVnthausste2g
ZQtlc1QeYvl8DkGfblgm0XnXqJR/NhQB+MOI9hD9WHFgw1lTgLXh5cwfB5qWU8a6YdP3r1VNV4xr
D0g4mRlhPjLCbR5iEgYJZcnjfDTl+1Le7T9ZkUjksT+MNKo0LmWKa8XXgIEc9Rx7uozPKwsXloJC
NTwJZcU+zsArQew2Gv9J/r/vTO820Ytlp4JRhiaeXc1j6bDai29T6jeDS7d3Q13XbElMUD0BIE0x
JklBQ+mpNJ7/VgqRDnUxHKxyWNtgs/TMd97a7bp6FCJk9972LpOB49zb5fjERYNrwnJ8SrLp9iUM
eakWV7oYbJKQfMGC79vw3a2zZMe6T8irnUZSr1sy+UjVmbvo2tvfEo3vh/yny3WzTSR2aQfhWDSz
U8RK12qp5NJwEWRmS1EP0Pg58lM2RbD1bKJadfvkmA+UBIGG2x+vNLyStJAnNtTjr7y9kV1X5D8M
x0mExK6D2y+8WYq4GmigE+mNMGzGMBzgPQuMgsdBibO7sDFesZBcpHfZ0sHP1V4ZDYZ2GWVgMUfx
9wg5/aqCO2SY3b5tGLPd1CuH6ZFsu0rZ69kvzZNo+N856KhsxkNBu95d4R3HLPbFnUS2vohCZoZx
gm2EIOmEaQVeiswHngjnhxlqxGDBnCHtW2jVG7hyLKOyTs7Sv3ArkIbNZhamhDYVkZZ3EUOpN20m
Ed5ErK13k3zxctD7QdAftWMGghXwfM1e920Cn8g4+DiILKKSFIBswaP7FwQ5fvDePv/i2q6rgxWZ
HQ/2Szh9MFpk5uEroswb2WFgLs1jmwh+7Mci6oxAzpv2ErLt9u4SfEsdX79tVi1BKAHp2QLWgwFr
Q2c6+8RJu0OyQ3naregUVKrcGDE4B5F4WNJ5tQslW9U2KH1oa06cr0JyRITOyPx5ZnYvMymK9ROV
IfpsTQV5KiGjKKS/7TEIGdRu8C64qm83tOfcTRoPp1dbj8GnDl2axW8kZObtrWBPHbmPb9OR+8fC
57Do4KDBLlfRv0Y4uWllssdHAbdJjJt5+WIfQ1K5Xlwd7q4XB9fqP221KA1i7Hm0qkvFkwlUY45g
faHrXLAr2EYck3j0RHwaASJrHfMD+v1EZIyFGrhbwOgBvgOPXAkGj4OzxxpDTnrdIAe2zrLingZV
FQ5OZ9sV79JSNZrHUvwCOXhX40CGZNYysdCc2uXkkPEYZelMG0w80atcFGo0MOXEEuZwSSi2NDrH
klQPVD1o2pfamOhdpOFGfqe9tR+/L5bGXy2yCs0xfJH1etyLgm1IT7Kfah3uw3uUxk1fs7XqrIaj
TIXDi4E4w6TG2XhEEYueHwWv+52BJRrWBb3Je/nAioBE9Zeeaz2R9scZHChEDXCwsdaDWqB4nn4e
Pqo1KjsSWB7XVaqvHvZOgNeIzn64IvWC16SjPs7rb1wKZvdTYUspcgcnJi55trnwSJbZhGTrNg22
GMDr2TyHmWQq65YPwNp8gVnKLNyxvx4lXo2RNfMvWjm5+4uJAATIDLVeO8IRJ2bKdQCPz9wAUNqO
MjaD1Eu7FDrD79zaQA33ccYSET7TwboHT5ox1jw1GQXtZhdu8gZW1MceEgL+Q4ACywZgG8qGdH6S
qb0bJwQ5sYj9HDVyfApxMsZQ7AvofcKhY0F97CCdoofIZaTlm+DmMfmzCr6ppc03Rh32CrVTJ19J
zuGY6UCDN4RtK6DX4v0wLcbIk52E3zHgis1+P4U4Ex2Td73FKz4P30F5Jg7buFNUcujAHMXVEMxf
3KH2qODTC0H8pudo1btEP5O2UtoQ+SZPFB0pcOOJ7U+WCsUXQBFrHQVUpqfk0r+WdSpmz4a19Tw9
PM/wW4dQDcIiv0U3nkZfCvWo3dQYaLzj4ZRpyeGzZ4dzeS/SLc3pWEfwOdHSEe9+NgYTRIBX5e8j
4HThGb9YtxYOHjbsWSMnfPYSfqc00O7tE79HNbPQQsZc2P9Pn8HpkxKoeEnruOJrkJbV7Vzq8WI9
eoG3t0bBbUbuPVo/3o1D+Ydn/NlaOmxeLxDivsfdLf4OhmIk6XG65U+NDthG9GrmIqI1edT+9NKj
Z7UABXX1BSYoFib1qUnY6+xpRvkvQXCmsFYaAXaLzbdBfRzFZV2nB2+pQPzXipN0iR7G1II5FPzm
F23FiLS1w6r9qQN3N5EfQFb9Ggnco9Z/IPE6ImETtquwJSN6mR736xsX2cJqfCCVBdXF98LPplZG
I1GOlHozebvB8QS34GA00HxZD/OQKdXdoToHe2T21VGAZuQpnDKCwv1wUoIc7fYPHLN0AeAQDPoX
73G6lEvzFcwqb83g/sdH1l7dLpBrCW5QVuW7OUDqXLFTWXsP7O//l+bt8RexQA/X4gMRcarU0LTf
boapjDUFItY+3qdMVO263/UozlOp3uAB89x7bzuojvDHISf9JoWT6rprgAP1TR0A+3gy82kenf47
O2onRCoSOVYJXWZ1Pu0u09eOULzjuLHw2oME15qy/x7j3Yq2aI7/Dtht/OIK5bdyL5Ho+ZF1CAyd
Ah3K/9QdH+kQVOBJxmIpmub3OY/3QUMq5t6luov7ofseWygH6viTGyGgnceB0rVu2G7SDePi5VbK
8EF6NZqLHaILL/amev0xOJhBcipUNQ3QwW9EBjV5CXXUMPE65aO6nvDkDNDrc9QvMjPOsEJ49dEA
GlmP6I8bm7wo7Zxyu9TLidihamFdLBxnu4RVVDNvpdp6gEcIne5CC83Pc23KamfzLq94SkcYVbWU
/z+maHTSpKyUgZuv6XeMO3OjfZu2frple1cHG1DWDMAVSyL/kSTN8A63xsviuxL4xmyfD2u1Kwko
iA4NpYnHrvaffUuSgB3EZ0GVyoNpZOAuDeJx8kRk5++ne3KXZ3i6VLB0T//a3FjcCMqOoFk+DWE5
f70O4AvKCnyNe/o7PGW64BZ5LJgo4MBN1kfOSkzDMSE54ZqxFYB4FUAZuQQEyAQpGAvWxG6zmz7Q
CI1Yqc6Nim5US0jUSHl3XQZzL/Qn5UBSNWckwrnPNfziiF02BUWGMXxmlHbaxsyqAFlwWOhpgARL
8AUtWjicVHdeg9ngnu8UyckGGuv5IxUdUABVjwfyNdSwesZQ7lknf9IS9pJz3LIcvbjrHOrXG7pD
S2q8VpNoXxIPyKtzkfExT/MwhHjBOETCarfk94wy1+HXOvvYsfYWs4Zh46mZnq4aH+c0Z9YGgWec
qqCuostD9D886BMD5khsVFmxc5Cge50D3ut/7Nj22dP/TZ1eJbF5b+u6gXJvu7lFC/um6gY6AIE8
xK1HlXaOmpagmwaM99TH63AiHl8Sb6ZCJ47TLjHqFkVcxNZVJ/VsbathRAG3nOKYHWbAFNl4BaBy
femxbzQ1ubwO4TwUDgzpUUDnwDNAwtmOlOFArR+ylpxwQ/03+l/Kii8KWVc5v3RtwH3z3e5YYUuH
nk5kadNR8s5ZSzlIfyykvRDx6OtHyR4UKGSDPLM7nGuw9PB4tc8+Df+koDw0+MCzI07B7uMH+VmL
bbrpuHmxFq4Li51bn9H9sbBXFS9G4zmDDUKhO/jHgD8JdGLyHqchy1+o3WGT/82UkfR9cbvUTlnf
MEK+gtKuK5UdKQMddcr/qFFeabfMJigk5Alnv0aQouPOADAM1XeDOvu1XNb6rYHplljs+Kmv9GXK
SA+rhiRcRpSLcDPanym7ywuYBTX8cXr0Y38+gy0ybLGBlFCtfk2sKDULnXy3+7Ho8UIMOt+gfq/J
2LgisNKA2glCteSkKElMan+VAk7hUYC9afmsW+w+8yUXlH5hmsVawZKcYwvGb/iPDtEPnNgwDmxP
8S9R3YFk+fw27qZI1zdytnParW+JhyA8N1O4BnrWmKciTYoIXERStKGCvJgqcGLNz/TPsaNmidhb
fTE/+Fge/laYUMyw9KAfzTMv/s/Rd+WTcdUaCE7ZqAMQGBkC1g5b9os6YZnql68lYdoD5mkdLcOi
taWybpxQ4AQOa/QdnIvtktJCiBoVGbqVnUD6mYdN3wAKyE1pbpmM5O9QQn5Ako8kkuXEltGvtZvt
a5N7NvtuOCvrxh3EPZ0F3Yr6jo30zfv4rZg38w/Ocva7A83vRnFp8OPo9RfNYRfoFhw9pcjH4j0U
vr9VEEEO/jYSYo7W5KvULTxtsdClvgcCwyq/6v0EPQcLUrekxpS+h1DbK0rKE+mGDxSsVQnPfhiN
7M9YxNGw0VkgKdbDSChugb9P1jfM5ztd9iXiZfJk2OFGV6Pg80DPww212jBzTpyNnsI8kdv/nHl+
mVsN8LDw4X+18tKoAC0HYohUcnNn1U54im1mGlPsKTXqXR19oIdolASaLo48gS0UlzORxzWitaz0
ibY/PF0c/XJmtGrwTvvUZi/lXhSfxzJ75iQTgSVxwqNyWfLZfxmuoH6fZZob8RxgB7xRm0vH3C4c
VHzQNLg7JFhenpR7KT6956ZPdXX1FYA+4niSc1mP+EhL9+r06jyyLE8RKz4wE7ymXlJOMSB/VOPB
1rHW3A3svI5PGlxNHoFTVZAO7GfDwr5smks0OQ4XriIFglrmdSTzS6CiNstcwcg2A1QQEs1M3qnk
HV4nAiC/Lz41PyaMJiy6bOkb9xC6DziRRc3OPH2jZSppW4Uen1v/aKTaoKEKzCVT0xzON6SP8g48
0zIv5x7FASRGIBUhP8QeIFDrF658hFKu7LxZpdq1DhEW/78GFixR1aMGXxDjfaNW9o4pQd/x8Etz
USzlNsL+jF0QrJY7KegvWjqU2Rer/nUKki1QdF7BQ9PS1b/2I5iU4yt7bIo3MG90ZDCSP/WO6wUO
fMvW8Uqt52uLar+ZtOPxyXOTOABeRNlkkE0Q+HhhMeDdif02+QezMbtDMNl2sxnCZXvMezPjz/S/
AEkueJQZzMCbdngMAc3vygzF8f6C7kFPyHmtZzW4VdVUS+qBiHMyvbj81kWzM0IoI89qc8X0vUhz
Orsc4Qv0ITxF1NvezNfMVnHVzpm5Dv9D9cSBAwGONZ70HFGCQtLoTruCwuUKLhkaroIdJLaLs18p
DYovFz4p8mkOmh1Uz5m57sVJIv9EVMfuOQMxmIPaubB8XtQXZQGNiFPWc4sMfjdKPGTOC5mnmpcn
mDIb1jFuxN7mqOEZF4zcmLA8EuqcxPR1ILjytJF44xrB+5QsyAqtmqKNm/TaCesU1/kWRqrP+vlI
kuz/zTNTtyYvbHvtZuS0qWY5iYd9DwvPZPwwbcn10muQzS/YCMu0Ryf60DYzP7U+i9ltprL9i4U6
pdMyl3YQws+GpggOcHFlJGC+i+08ct65C19xV1SrZHDvJgaHk6aTlMtuKV/qs/9TeQJY0SBJJaeM
5TxWCNOWLK4J/9RTJVgV4O1jltlL3tnL9UJc9vYKzK++hPRWkGLK/HaRBf57WrVlVu7CBUMJD8lk
x7/iEVtWArIkHHlcisEzvqMe8WWQKui6BZoVYqJwbKIg3TGKliupktZs1SjsO8ee3tqk7ddssLxy
1+I3DVj+ygrZphkF3h5lgYJOQ/wnijylm7xMr6fp1ALOkQDxIQOsCv6/0l1VLWIN7ClEIe2UVluv
CgbMIiLizg/o7hAX4wQnz6h4xa8As3LCov09NqgZCtXIW3oN/7ksooPENwFUOHsFvJsd6lIFbhfU
Q0aAD4iSr1n+N+FW6uHvXYAPRAbcz0PG4xEoPqxe3k3MOXVfx7iZzd7i63Af1yDuefca8IhD0hDx
aLsQ0GXK+2qzRJNk0DE1JIWG16TBExQRsG3Yq0LQTWpKXiKacwwOIwD+Z+MxyFnYXg1jiwvV+N6h
G1Ms6YJnx9CWqTQi23i1KlLDWf28kf1rETajTH1RhzFXTjxXaOeC2MTRWNtEIeX+uFrp6CC2pWBO
tdIEQOT+/9jSfr22zLucMe75pAtma0/iTW796AOdv5sSzoua6iGvLTtK7AF9UJBzqPtEXSf3Dg9i
Wrajmn2Iz0hXhadxSKcp73pZcZ76riRiYYni+llGjjyuyAkCf5rpEYPw6hNaHLOH9on2oWHLHylc
PgwgoTkvVgmGKC1PWxrh6Z2Nc5AU0I9HAbS2Glb7Ar316XNRSBBZ90rQVEqzbGOT9A5w806YpKc1
gVxGAakRTfLvbinR3dfIaBlI814HQjHl/9QMtCrf2qNHC8fX7tiFBJSnoEzekXVchMly60sjGXRH
fTvZ2ezdEGpPRz9XWrJMyg9biHPGkPSH87hH75csksDka9t9gkk2Rik3WWtdiCp0Ou5hCBOZwqU3
jZSdYOFmFg4ZxEHemZbst1MYPoeyq5CfoseNK0N16GU8jdeIlfdmivGPLEk1OKrHqF3QnvCGwh/t
oadJ+OJ+ja+SkuzoF+60PVHizSi4zJp3J5GnIkJmRDKzXXX04Q3iFu3diErBbWQMDPW5U+hknn46
3QvYZBuS2XQ0eEKULcrLlA2bb5POjyX5cvOfdZMnIoRpTekuTZPmqlM+7KayRcJOc2mLgqrd9Gie
ZiOSa/SN2HMkM85JsgzB6lLYrfFBdVqQScYf3pcVR3nbPTTNJGlOcegMwvj4aWP7BJSi+mk/BTBg
GdqbjEgIgAa3gP7JEdReFNXrKoRzr3W+sSQvGaToxZFChBhT3Q/ZL+XldOOyMVP/+g5ZL1if0shw
ZouEEN3Y3oWHZu2q9j9h2Hrq6+hjeCaAeuSTT6R3lPgmq0LZG8kYIyRC/3f1fucT1Ot3YtbrOayi
RUXbd1MXTAQyCojcKTCVRABVsjTfWJkUiUNtqhR9tWGe8cylOCaH5uGh9Kzdnqy/IBYPv5/UZDfO
IB5/H28U0wfdlJ1I314aTLQ15qchcf92q/YrIPZ5uJv3A/b7vt+rdjntA2jR3daEcgc/7GTlR654
jT8JSo7wyqBOfWuxtKsvO1n/nZcxxEnoGMfGrql7iPkifdfe9xRZfDa+wSSkMrwNqM0JZXF6RWNw
+vzBeLpSgJ+HSjowK0/1xZnpwk9xWtuiFJZOyBal0cTTpcERBcDu8xHgykB3aZq2vJKXWpxaGDYB
P057lq9HAH95dAarEb9W4FrcMQ1NapYO7UYOVEQb21qcMdxYobZcEsd4FRpFqX3pD2QBf4o86A+P
0lBXwMt5LBgTEq7WoJEi1meqYM6y7GW8DntN78uoNLvB1XF5PbPoL1WFrsbTS+8210udYg9rGdku
MFjYiy8fulMgFIsOUs2PxmXDzcIrdenFMWuYs5tN9SDXlM2smsHGIgksqHtp1yfNDhbLSAm4Fstz
SuSKiAagUCRQzeoFqsuHNJKqRaMPaiI/0BT3KplsWBYHhfTgQLJEuRiTfEMxx6zc+vzLPz0SM5FE
bKF6ypkO5Olbfbl5CvvxyOnIbfZL7nd4xZtr5WoJwYw/d+QLUMl0/1Xmk2tvrix0L3h/xMnRD3et
QKR7ybiPjodzu2rwy1jlMw32Ng0YCwn2PfjLyZStbeuPQPu9pSdt+1MtbeJ2wLW6gegr9Y7HO5xI
0RP1P/TzTf4PtPrLq0wpIjCOAii5ylrVS6nyLwfDiKvdUB3Ot/mjWPFiIlcElFfuVacfeXPWDqlU
ooTXaeVCpoigXAwK/QlMGT/aYiKqSYNGginrJBYYPVtaFvoCJuydq11UpLNNuxiPgIkyLX03q0Ib
uIhzr78lNfR5cseugaJfC8UApNi4Tm7Gfs5u7w+fPQxligaZL7MlM8YVNsk9jjM8P8Xdf9jZ2eJe
JBBk54MspzlThUuIIeq/Py3mMHtJsVCfC+gxfIoHeGc+jKFhZUJ69XMIwtld8QW93QAkq1/0g6UB
oSnhQJoM/z6zRSim6gGpEjuNMS4PV/+VcPj1Y7pcZeZ1O62HHVBoWQOehlI9JtAP2RrUm2xTZj+b
tT9GiIb4dpxwAO8P86F9YP1LquM7E5auqAR2dYW25jeffJ2UZCYf8oVT0P80VIYDIayl5ND3llw7
cnwb79jzwA7MU+6390Ebb1Kg1Y+P049VUqfZESdIPBDWmkCMQb0SbVcEBMaX6gNGJ7Jfzri8fEGa
A1+SeIgDx6luF3VcaIqTM4/1s9IcJ5kNRkcDzylBDrFNE0W4s8xkXfdGfGwKBdHo8qDu3oWc+f+9
nqcDtC1lkxo0l4XhUfy9ePGFghW4Mmdxry+ZphqkCe/Fli/ZIP/UXa15SIzpAFs6FtSoQCdcHXCM
SUvyEdwPLBjugXrcVsqg7nQH8niP8Ka6h9403ing2WWpHnaCrlVhEtiS8b/jDsJ2iJ2D2Bsn4Smf
fzl97mll7yQW/5L0vZDfAq4U69b4V4sXJiDZS1IXzgtzhnrlLclsbiPJ4b/Fp7WccyVfAqx1CGh7
BJf90gnKB4dD1zBFVwwafqQhgpD3sVUrmXKkDOEiOXTuWPBjDvaMS67H7IKDpT+r2zOqh8uMCog0
e+xrCGhBIifEWUi7MmXMax/tq4w3u2kCn4iUYjNtQU0M9oI31IU2bkaZQoknJLpFCbtnkiXyFO7c
+W9gTj1MjFv86VTS/n/FGU4sZ00hEMdui0Hkat0RjIc75wHVYzn/LGQMokFh6V1tV4yIIYdmpTrz
WyqwcBwtHXDzobuNx+saOmeMOf6vWcW4ZxweRqRoBJ7GsrZS0t5qZRhHXk226nJG4cm2EyOCWTci
rTnLst4DXskD/x49wa2x82cUq/hj8UjXMIlUYXMPx+EPj4VSwFgi8JeqsabpmqxHHqhXbo95tj03
7VeVQFcnY0rauXEnj2K8KtI8AQqOu8nmEL/RHb4kF4JeWzGrvjFENjE4IrgA+7fntcAcuRj6D/m8
RVuOL7Q2H3EgmEjf8IFKUW50lzc9B3OA/A5vTFpeNZjXduDqrz0dURaV/0R8fx7LZ61E+SpFXrEa
CW2nWsPll70QyXI/v3r6EzLf65kprceL0CWgAGjvp4Zwagfh+7gfNVIdhkxHkrh03cwZRjpJrQcg
o7VML9cpiB6T/tFSnmEp4/TrHVBtPVhOY0aMGQArxTVo/fq1cUDG7jz71wfm4bWFqBgunr9V5gVz
oR1y3CAytvw9vy0zi5RPS+xQQTqqcwtUNbkm3h3Z9zH+kV80yLrRnzajJC1AG/qY2cl+Bm7x/2Rw
rAw9YgyKtOlHqflbER39Pgg8gg7RbFwbtY1PAW5BrUgrKO9uCrULo2CsptwWMtq4pPcnxq6mvouf
ZlkyhGgwi6z9WekK3INh53lvFB1UXZ/71pO+eKf463ShP9/ciYD80yo4y4Z+JM4SFLYxro5ebt+K
qo39sOJrHu2CevLKGZMxeDi27PYBKe+i4L3/2RFdCv7uNTVjh/r5fnsCHhB7zWLvun7F9cNN/zUL
nz6KfF/3q7gI6sqRMTRYkUDABgWkCG0dW8tW1lhPzHCd2DTDzMXPCjo87k+kt09JfucWJqSwsbS7
6j0uqBDrJqAvmbtPHrUbMeVc1a9cjZjrFAVomK0YX3H0TLEeL//zQPhLRYjiFcGbzFKhCWWSIZWJ
tn0zHhvhCz/VjgcT8lW1OCaV5heJOytk7LipSOIB0UOE2aC+eZ016I/l3tZSFfbecCDsFTaXuVgt
nVFxzKsW8zxT/OEdPwIYysHb2b8R6ivI7PRX4e7wRPHgnlv8ixVqm+HlVyml65lfJRpQ2BTn57Qk
Ai52A/HAltKIoFOcCYbNoaNYAt8nP3NGZy6i6Gi9rHhtx31UtNC04YzytYZfD/T30i3NxcALrWZh
9znG8YNuJufKDw24Qsj4ozp6q9e7eohWNZwABo6gXF0tTd+3KTYsqLz7oqvV0eJHBCltNC4wMr1U
07DgsTRg9r3zf39qAmYHfhsUv4yhmeEckgCQOqsuH8hiwptUN8Z0rK/V8v33KqKYxYBB5bpGSMLJ
0o0jpbGdVMxDBz0pNJArFK9ChjumOfKP0JYcU8nxra3Zx7JMbwFrFhKP5JaAFd7TgNFWsjhx/XAY
9Lt5h+WOJ/wcVk3RvdO9XAHW2MVhPWmq7qTAsUiRR8e1P24DnIlRqGDxcyjNfVczzx3ZIvKcvbvf
K8kIvAjnpN1VSIiJ/7B44qrmGAyIJlx4psvrMRz81w6lAFumjtfC5HocABWeJgpPSfF0VjixsbET
xRMAAo7bZ3CLW8QLJcpDrQpYH09E9oufg6puaErL1pFpMvPB1XHKe9v6zgUP8a+bbw5IC7oTqqSp
ma5XQkxW9LzBF1jt6IlIOXnpe2bZXeNruMIDoTPxkD6+ZKswNs7L4VQFQIQE7Za2ckR5/XoM6x38
Dy9GW5qTb+gKB63i0f70EZKwKcMaia0BLtghwpJI8QHPqgtWj+TglNxOkOcDjPjt6iVED/jUbRbi
2bWzcynSIjX3tKaw7KlilspCKvJ2KaJLcwFRiZo8OcC0VJMoF8zeBZhEwNjbFugtxf5e8srtR9ZO
RoedfT5ZxfuyXD+HQcS07TTtL+2M9WSNiEjolMWQayj7VED39vER7WjAqcmT2FGqR5zSxQ+18rti
T/JifZHtLvfeGSLmBQyQNsDBjtHCJP3C+OL74Y/jZW19YnDfBhwhk2R9DcswNDjAdIF0Q7Ynm6jd
9iqbVOSmu24HcN0zFKbHzKlI+M5qxFp/HNoA8cFXOB3QYESd416e6WNUWGlTdCN/O31OzFvwDwWa
r724yQVLpFuv6EmY7mYV06qFRQAjH5aK/gILAJ28kBoqWRqXsNu1zxR8CPReKDhq7M9BX0mgRR3J
s3iDHNKJ8a1MtpLTXXsdsQsn59HarI+3AYOr+HFAUn121r0C/MGUBeQDXhSIJ1tNHUrnJI362QXz
Az899IN5Yw6tyvL5Y168OjkZsVRsb9R85VMTvz3jASw21ijOcrwg2jD4YN643zMTjV0VY/b3nfT5
NG7FpqLrJl+ybzd+Hb7CqIKzo3waqKKyyE8Adi4SM1FqiNcbzN1yJ/sAE8FCJqb1pGZbQ1EN/d+b
RQ2BM2SClF9WaXsSNKpf4lYodlAN6bcYBPJ6FTQIIOqFekJZRYJgFymexBLBLrbnUyMpCpulaN7X
eQhTL3cGJAiJPFVa7pQKGyDe7/dsHKyVGbbJqtAGuVQT++2pUuIsqFW3rXlbpSdMan5ObtBtJjSO
4ZIbDrcM/shBGTCQvZk7YkjfKyQUUtbOLCmC8ysvNCXmiyP/n+QM5F8hnamzbpO5Ucb/ZoQyEoi2
52dddd3yU3TRAtHEdyUJr0WViDiMOnRWbj1eQkMNroKlwjmuz3Y2DhAoWiY1gi276nQRqEJwmpi1
9T6A7kWJ92VBMlhpHmqfuPaMAqXFZwPkVb9scEnQQ3GrI1fNbmqpyYxsarNfeNoNB3vamkbbnx1q
ZuUDdxGv2dqRMn040qKsIBJ/xITk93gZIXo4toCwWoGtoyZBtv6t73TKmaHaNF7g2Z1WbK12rsZX
J1VH+CFLf5OFmxi4GZzOvzYz0k46ZSXf0NTMnV2q54QVM2N2eB4StNiPQYP/pQQrBXPMYtP1TwOy
AH0S92YrXQdfStsCRC0TQkBDvObkGqZjgi+X6TwFT45yqPUgSejga1gXHIoMAQpK05GgA6Eu4LDp
Q+xll/Z0VcBpNpYuLPDHfV4wGbRvkF2RohezoGbaRCy72ncGyINBkrmNAIj9nFuuYORzgRzYNvjC
ZyBUsrRsgNr3ZbRdJ/C91nB/n0iC+wJY30Ne64LhoaaY0xudBuxd04zysc3divc/Ya+lIEU/MyNP
iQpXIdXMXk4HQTwXHTR/Za6o5Voe/+C0t5AYrpByz2HEFaQDyS2qsSDqvYRiyizjralm2+uM0Yuw
O45ilqm10H/WodC9R+53+TRA1Bn7mL1ETGb0QEqFqYF0pQ89MrpndmED/rBDvQ5ZqZAUjTrqw1uB
BIYcfG4lJVVPxLSOzTMUASZuz0emmA73/RRO2xvcEjkyzGJ5F6E4oeDx2pCPm/NsQKqyNbrB5Tkd
B+s88/L1X5cAbleKwq3g1hHxyCc/03RlbKKWjnadVAHFZzALDKJRObetSq4YamkCTyYYNVoC33f8
Ef0FZsH3wvTgA6/4x3ZV2RGxM1N22mfWTbMcTPrvgUC2P2gUMV4usqneEjY/uhvfR5oGFXwWYtmZ
DtSdWVfYBZWbqrxKLQMLc0b1kTEc56U1GN6A52YO6Nl33Xpx+OKkmn303xjWm/A7X2su8TQ4OvbU
WGJUPNcLYNDbvyBYktWF19bqkIZ+WXZpyGdUQrub6IyQGxuTxBHTFzlLTOycyNsxwJYBRSSO2SV3
RegnPdBtl06ZaRIcOYedMpXHIfaEf8aOsfv0Oe5j+pNqnV2yKfqO4Vv5SWUmc6W/xQarr/27jOQ0
GLNI8ZLez0jp6V5MqtWRI8yC08rKTHtnfIvlzt92ULXeFdQdMcQWcZv+fHc9LCsuPwzTkHOgMapY
L0OLeOB0vJhtzz4D35bloVE4sPkqvIdHHMoWlkcTvXQ0zqI9Hu4GDZ1rPd41UnnGjYKtHs0ZsPiN
sPvAOYPWg1dEMZwmJpvyxr0f94J0QQomgM+QHBrYD0OMCUzXRHAP2LdbaeUzLlpvfdhtMUpCgsSk
MkK/NZkwIMaOVeX5DD2LCqbBWNzGiYybVsRvdzkcA9aefuNk46hhwqXZlYmOAeLTD0gZRkn6EZjs
m0QEy+efnwJvXYhFywfEMVVOFotOIoylmBlRm7iA13nFVERmzfggSKnznlO/U20wx1bGjjnSGpxu
I0aQJKkxfqVZ7l6okNjKXRIv4USO3Km13EhM7VFeKh5YJBd+Phauq4+ZsJeq9Llv/vwz7xmuAoJP
EiInLJAQ92kaXwzZ9mF6U/ocQ/wYz/cjXIrL33KxF/b9NgSfLeXUI08j9JHMdFMu8yqBg895RYTl
ye4kzr9LrO75KPcASe3pnJkyrEP+OSMoEO0koUtwq4gRDh74MwpA3c/Nrqy5mQMEgaNGdLLL07oZ
R4VT3NXcX1DCsRJwKIu3yeVF6lKGoYozdm00Byaovq1D6T5ALr+JtrsyF79x/vW2SgdZneDzpDaB
L2B0M2XGAD9jnn94iLyzGhRC4dgxZM3HU1KPYlBsfdJH5/LQihiAVrcX81iy37OMmOLhIBIGNRJM
24DyPNT2PtRQXjvDrUUpMZMe5n8sRVMkjUUYKQS+Y6U3y58WMiGH4Ylz7TECWi1Ea21YH91TP3BI
EzFlgtC5GcygBLRpae9+5DTDRFVM6HJ0ZCj0a9ZDMhS3CWLBiyREIPscSI4ZeVbDLh+Wiy46/Jkf
0WH5qYffsQg2Ovff72C3O4SHXoQhPh+I9Qb8ue8H/erWOfYevt/aaXcw9a98YcfHCEw3KClwpTs+
cDpH1G9Gwpu17yKMBkp8SGKb3c0V7JfEqt15vNIjgH+K0ZlSDAmLO2ZuU5jPEo46RCc5GtghxfTG
W/mH5i17iIWUyJv93cjxi5vDKgD9eKIEtZYd5xzHxCUAUNkok8e9Yjl1BXwFEkLYRkm2LB7UqluY
sLee0wFETDmILOCFsrh2zwqOeLH8KzWmikiuvB6HkcOZRhgS9u5CNV4EHAhYpCb409dusk1HSBmd
dJV5pAMSrfnBzmVDjGLHFE/Z3x1h+1WCsAxJoDFeII4upD3m4z0NoXPj3JigjiC4FPm90+K0kmYU
2znWsR66TBXeWxDLzV3/Cq1qPGKyZUfcueoWzgp1Ejp4O1Ng1aR7f09G1cxFOjR7iY24H+vQL33D
us+mNfml1koU5sk5f2tgHSFtPL54K3VA9h2JHEJ+H8Vbxkt8XGEGSV8g//ArC017CPF8C+ZlIRcT
rGc/bVzPcOq4c5Ew+UFpkbyBaKIxErybCT8sCR3a4k6Gujlkr9nvzX22lcj9EE1kvHYklNC9db5P
ycqE24iT1AuoWxLqzC6zfx63YAqlcUP57IW047dldSq2QTH31R58ruhJreIRAF7YGsedz9O/7vrp
dLdGIEfQ175zIPXyC4d7KqRyE7JSxc8dFdvT6YmdTQrEWofopYMNuB/yAVCZ3W3V28ON0qEOgwFw
+0JhCwxuLOdKFhJZV0Rx3X+7wnbb7KtISM6qvXX5RPwxxPyBOYJNCzsyXH+oM/rhAD8T88xvFpva
kS40sCp072fO7bEbEN2NUkf/o/G0hydBY/kgeRW9A6yuhOMoVnoUSF56Yz5iQm9tcnxfus6ypIyH
gq/2ZcLW17WJeC4+VcPBWZmNDga4p22aQm8p6m/zV2y48YZ624OzxGKXzgONHoPDkneJwQc0yhlw
0zuoSSw8i9QLFqXPeb+ojidA3JKYh1EEuQD6lbCdFNTVFnhjGZKcf3Ki2PnqGP+gFmmB1NfJjf23
bQKGPmJY69RGw2OMk3s4n/qqR/BgcQ8CmuIzA5bkdKxL9sTe8UZxNtHmRMyUJmKDo5lC4qdFu8/m
bRkA3fLi0jS+/1y7pmKebIEVrRz7vn8yiZr/ZFBhcrz8F+JKFJGmUD8DX//Uet+Q3tElHVK34Spr
FHDcz+RRAxzEhB3ZIcSlyGZqYvSz2HuY39NYhjgNYU+fU1HrBriNDFDX/1Xn5mKbYXKA7QP47A9s
FqvL7tpaLgBm/Hmr65IaTFksuiHY5A6fpoc2H1/wZTLocjIgc17171n3RFzqkjJ+b/pqcyh9flgU
0EBtGmrsJbqS6vN0lfIUH9y/WzTDmT/+7iZFn01f7WFP9hh9ketkOv6RXHR842HjFTqy6EJiuD54
ogEL2rG4D9pZz/gaENytx2jrNH3OpiYuLeiGVIGvc5Ye37hyDPIPrFTMRv7sciT37Vih+GuR1DpK
mLleBtSsGF4RZVYygE7xKXQrzc0hshfaDX44Znjhd69UyddTOm56pmXKUmnn8uG47GmAKQMIlwCT
nEwRyzNWIpZrgaE3gN2j7vw61AK/8VggCI5yH0eQQG0979zgkBurflD3t18HMgzR48sJjwpC6ebM
VckKK3St1tdKeHyROyzOpGbp4eOgx1ebraLRx/P0oelDKrTrfDmT5ehxxv+iBM4n1aCFHqZGMUAq
vDpMThVZlUyZ3N+Dma/Vec8OF8DOmyIhG+whK0F/O7de/4QorF+FYXR9QX2PCFRxdqzHKnHnqxQj
it0KfR7cMSCUBYnavGQ8mBrHuPLj0s2r3LTrCK5/6WsTT3RawooN4fBkpHJ463O9sLK7T1qAUuQk
3Kmgw8Zlrq3H/jtBy42Z3DJ0Xv6YxHwpRjVRTXdqtua4ykY+x8BJLqh/6A6lsOeUA+Wfl2HGauoI
9DU8++Gnsk0SKL4uqR7FkDt72AakOUMngb5CB24Ps3K5Ww97019qhl68SZd8NqCEdX17QqRI4EY2
fR+z+DdnTDiSbzezGiLi/nOlwzuwcosFUV6XcFNIBmHkLUQcF85vp0RuZEAnrFNyCRbYYrzh4iXX
3dHFkExZZoyNiBtPZPQFphYSX2tyyhH1DgWbqIBYo7PjHkNUJU8T6YbT909O0EtMuGu1JHAzsmWr
KeZ35hNlF3H0EZDfnANHnXdmBgWAmQOHElmDQLSWd7McZHNOkLeRKaP+uZO7Kd4VfH3LXIa6RdUf
y0aLKSg91BaJbjkr8JJMjQAC8Uk1XRnaWlhhLqwmu2wZbVdYY+pSD3AWnxeOcz+KtYcGGKSINkc4
A+8JDO6KydXgxqTkpsudmvUYlQRjPzSNh66FTlsAgZIs6fLAn2xfDTaEDjpUo2fr3TQK5r2wT9fg
50IQStGw2RWjnY1b7nYN1YuGAP06XJa9Hoo3T6KOFzxE74lgrOEstodeOHaFBz4zKw0VFhFzFUE9
iACsuZWPpaHCBhir1JJAv23zJVcUAjOGBjO1erLOExyMarBoYWB+EXIzAM2Q9bZZYj4zwo8I1UNs
2c54mXmRTZ+JVVKovW+IexKmTtsYMZgvUJEr/8++5jnNaMUJ6vR2EORfWNAg3wQc829mjHDW6mLs
mT7FIZOQyvyH+m0h7ltccSkFmW1HRXjfBNRcB/K5qwy4gk3rFzM4b32pQ/M8PQgTxl9nRSFoX5y3
5Ew9RpfmxRjYrqBV+BRVLJfyYMIXrHLCczUIDnbLl+IlusS9cfzTj5XjbGNl5P1KN3zUQm6em6z1
PNd8RN11Jsn0ehDTMO73yAkp5txtGGSZKPfoERTJhwDI0G9TsPyox+iuAqAaRDDdEFDCxX5lEkx8
ygduSNetiaocRyjTcYWK8aoIAPkrme6dqLs/mxTpAPuZLVmQ6bEhZtbSu9EttJA8ntHGSBOuvJXD
MkWLEq9ZbppFZMuXPG91501P5ddUBuJ4K67zSUPZoc5ZQ6BbnwdAbj3FTAiOgbaMFkKiQef2xCvS
rEbnsc6sRriDXIIaGN2d+qe3XhIQBB6OU9oQaf+zeCNBL56imTqAaRWrrfrIYIGtc9p6eEHmTKMQ
YB8UKVLKcVK7LyzDrSWp9WIuQFH43KKDqrCN1qz5PiLmMExoXzMHetldCBJsDy6pndkWEls4RJIZ
AjzXBz8yf8F5nwJrvyQ0mLw7OIH5BGDxC05J9/9SXTQS7p18qgUW7HruHVJ5RyR/hZ+SHaHIW7oN
cqBzJiPcDVuODOBpd3pcoXBh7+O3x8DsXRHNG+IlGjmp5XuiiRm89rpz3yo3Pat9zl8VPNpCF6yP
DkEeQFXYV76RFB1KBIcTR6+3LIhADlqe4yP0WehbmXjBRkyEiNf5vvrhwGwPkflXC0W30ZiolUgV
eUUFguV1+gujEtJiRhAhAyyWLR8Cv70tWJ3g5ZiudTW6WDHrhzVtMi/ycpRK27pg5z1TqgzqFDhD
EGgIweO9xyf2+s/mC57YS+mhKqC+/aYy2v4tsqoE6qLs70Ajd7zXAhr4iavKzcbAnAivVRJi/j2N
RJRdl7x9nXgqvJb6XeSmmB67ZvvF8YhogD7/um+RhMy+wtIqi5Rsfmkq0WaIWs9G0IOxvch06BEW
eSpMbNanrW6bW54x0iOhb4z/kGr4kSMsmnz08XhSeVVgqTAbibExrA3KwvjH1jrXkr1ifqSA+3La
oIp7f8v8Twqa6A3ZhaDrQW3YL7e8oqL7Z+odhXwvKx6a/Jlf/uPRpe3yH2mVfL4hd+0Pz2rnJD2O
5PPIJrwojCi4wkNJOPzer8GLPZg7sxvABt5lJ4f0Jva+fJchHyc01Kdy5BwuqgNKuBnjlBy5Q5sa
i+rh9JexlF1sCSg5ecXTgJ3DaFMhwb23PZQ3tQB4hf+qTmH9utcxLb2OdKDd8qxDmqI2vxAH9vlg
7wGhcJghsl9qUF4+G3h4+BARxyNQNVZcW9E9P0KqhP9V6fg/jVtDhSqDZGHR0qGA6e9AonuE9udd
80Zz5IJsXwoIYbMZzkz2b4Cl8Rl+mkFFYDyxrj/gSIYng7XwgAML4/HniqX62h5rCrG/4sNBwiuJ
hHiADVf5QYbEG60bmDy6p0CxGsia8cOxtJ0deAYv2qOBfdgxpnQbhVRkDY5CsqIBuvC5DRUqZka4
Ijtvdd+ZBvDtwgPzrf/bdKEqQj8UE0XMApmdfWWhULok4PtQiz3m2J48zyqlTYn/C15azCaUZMAK
Fc1KtxO1VaXVz2/eqxvBP9Wp6Ybq2Lb1VXMZ+/8NCScCQGM3TlBl+oTiTn0HhqLcJsAaNon1whIN
SOphXCp2HCv3FDbsRvr5b+Ws7M2w70AZz0kF76o1JenJigMvPvKH6ApoDW7aRJCvBBt69XdfZHE3
CG+a3AXCKwAQqvqW0Nx2r8XPh7jparkvA0sOHDPQ8xgbO2XFHECjlDPXkKih5h6rQsgZvv3xqFJM
9M1A68wjzjRwc3jxBNeGcH3wu6mZlopqJ4+ogxUxUwtcjxzjuHSsWt2xNSukQUHAzkfliaxUcTFb
CIxwCtht4/2jwUZuzFuJ9e+50OANZjkds7Fpcpxjf06mXZTIij3w7DcHqbztHLcvp5tAhwKP2tn6
trj6nuzxmehCDMjF3GOYT/nOne6xZVRrOMvoxk/9BOe/JNKg2/hmoxlYdGYd2OFyh5y7Kl7TVhIb
lmF5P+IhBAE+Y2FK7lkN/IJeZPk5BpETnhmXV6US1/VXAp6iulKbt2QuxvBSWR77ENPniFvn5pJJ
p0EHw3f4bUJTrV1ChKaZgbEXT37amTX8a9URLACYLl1c2nXPs2904/qq+Z2LnXpxBxvdTDWiOTSn
cGzkCm9ukQjAPckTk6Mb5N3m8UFcdQ9emPcIPgI3oWz5SSN+4tY+1Hg408uf+uChPgveWvxhBQNK
MdpBzZEdvSB/nOmPM2FbiLU8AupdrKaooW5FQySkk0rN0s4K3/pZfk6Xsoqbd4Ufzk5N0T7YKAfX
yVW/xDGqjupPTRaTytSjG8Vwuoj9dPDoDE1yXYDoRaaNWppddQhuEHpeL7xmyntiWzguJl1AmoR3
h3we5RZ/TmzNdk/N2aocz4jEsUIi4s8yNRQNk0JJzosOmOA4z0E98GC3YVGGDqjShaKvmfYllG/7
X9nAFE4Ff7+sc30x6otDVH8Yly+k16SbpiVbAALI/O+CQuaMSh+x6/R14cnoIR9LdXgzbZ/ptUwn
ghWFK9ZFmr6WnyVfbPW4ifX3rpUqKpIbO9Uwd6aqD5MvMyUC0AEKu/cyG1Dfr/LrJq4l2cjaA0/T
50uXgM18pskjjmSQeqEJbJEWCtNmB/0w24KyyiW7MoZqiVGIXRTIsmqI9v5ATd3P51d7ExXfbhGl
5QbYcM9EbuXkrrF5ya5k2lmpompNC4cPs4fBoWrDnaON+N4CcWNOYX4Z6IPAJ3MIsH2tFBf+AhAY
9a7zAzZMrKjd4v7UKjTk6wTZ8hMGYPNlI4JrZ695iMX9VbmURClUGGEQL3rmApBmUcPpxCcdUn9M
iWVB/maawCZpiTpSjEiQllaBbmhUtMWabvDFnffIoialeQvzCOUuFgJSohIbJ4Fth6dS4ql3b+QT
Mhbzu6q4n7k1qDKilqb+Gnj8+eqeZgTnCeU13sIoWs9Pk9hTSny69FrCeBmihB/OM8+McGqdicaf
ywtQGwkXSpqdij/4GJLGcPRZZTAaLbdYuZTe/ayKYxO3yr/ZMXKtvCdVZY1b+6+V00RjdKflhgs4
etnrJj4qOfLs/qI3ENwomAGF+H7A0dWXqODJae10Ph0RAfyKf5MXNnvia1sI13GLrXMfoutMnvB+
IoTMIAQlP0A/GlOdm/btH+pAmutOSnI2++pV1lyC3wNSUZnTUKSElANY6wlHeOBiwuL0BnbS1Aul
zv7ItUSO33lJcHR7lX5qlYf5ZrWsW2WkXYfYTfP9mCIQH+NfFGBbDeqyp/Te6TvhjLSu0gUxOoFv
H34w9lDoPbdX0Ygz8xm5j0FS1K6KhKVhxx+S6E0iPkWrKkXrPHKWPU9799Rzx/1HmvIuAwD9J07A
qEHkigsnDoFyeFg0q9PvSDCvvbom48MlnWiipOd6P4JbqwfEmTZKAMZvm72QJmUwudITQR0Dd07O
stmxhvpAAX9XEa53ubaYDeUwgdHg2Lmn6hZ2dtrfJyOBR7lofPDloUddefsweyaP6kiB02D95Z/U
IL2oL+4uXSAE1PL6pp5mHISgeGRBb+cT2UNe0LaC9R14PGyZOJqbl0wibCs87uN5cUJAiZR90dcp
v/3BahJ5DxzKuOF+zw8XcFECzMYVl6C05zDc3tVMp9nlU6fbF6HyVWwZ9iLkc9GMnkoncXeWlVw5
wam4nLSB4d2uN93D+ef4/o1nKcu40R2idx1xW9QwxxF2mvkXTPs+mjkWo4ReAxO+Vron9NrdPgG6
VrCHyvoGWDJWUnd6zI2Au59d8HpKn3QZlKD5KAMT7yN4Cs7HSLTJ1RoeJCFOhpJkdj7zqYneRURs
w4G+aDtIDpGIBKqETMfEJNTDTr+bFfdbVsZOD0Z7bumicsn3lqHhkTYqWvYvkHl5DzSg3yu8m43/
PIYT/dAkTZP2zjzGVus5iT7CSFr2EIEttCLdMSo9/P+z3SKy0LP5hiFZMqJ8XjmRlZMN0jAkNXIR
slvulSzWdCvCjdy8n5STJhHj4ApNpeRpfz2CRSePRHwps3FcUF6/ExzNguWyfKXjQrvLSMjURMpL
L1dFUxSVBuKO2eidOr4OlstRv2HzWqHEedREsA7WyMIHgOekRhas+OTUZ7GkntXbpP9hyKqcdfsT
MyMjopUD5mcwcm0klaj9SkUwfIu0LliryKtsYaksEyfT+GvduFTGl8zAyBS/Jsh7JB2+Rm3K1aQ8
lr6lM13WS1+gQZubwAmvPj7CsUtsu8ULfhh27iyOM6og5RHfHiH0Ai4+gqPh9mO9Lg9jADX1FY86
yqtTMb+7CgmDBsdfFDN4tRMO9+16rlPvyVWIK8fxWH2RQAZ6pTRi5391PYuJ5YK2PojqZ2SfeYyl
51L5IbPCj7UEHQlQ7FgKFcg8478hqK6xiLMHY9Ae/YCEDNBST9Cxq3K8KJREgXfR36xH2NXpjdkZ
f6dlPos3FgXN7EDz7XyN4vp1MsK091hPc06VHKb57ijokz1PARAy5320UUdpXPobLqhLnpZroeYM
7wcRMOfdLXfTyH/s45bWs14PDQtSRgZcp8Sv8aR/XFXwFO73VKGH/jU+8l4JXAAoFVkY1Ge2yGnK
h9qRA8XC5rqoiK6vYKuY5EZ23ptr6PBlBCv5UT5IlPaqIq9lyjX0xgyspMHFRXm+PZs2an5vv27u
aVBDT8B/l3a2jWzt5A7/VsLasBQKc0d+hXk9QfbZXtk8t2FIyQEkriqQcvgCCKXYTvowuXhHxN2T
T0p7ImZbH86ReF1KLTarSYM6MN6e1BF/Kz5KP2lFCBQSyagGHKfR1heoyrqOcq5gE4HQFbm7ZqwI
E/ABuw//kSHRrYynsK8eDpL3W8vBc+7d+9SnC+89bqYmIZxPYlYhlKzMLPUbcTG835joJ073vN03
G/X+MCmTqIL3eCCbDUw27QB9v4ZMLIVd6SrSq4zmN7rGB4WqIl0gcxBJ0My+6kFO8R2j42+NKJJL
wghAX66olJKd+jNkoHbsQDPV7pvY0WYYqfy6sDwB8/M2ayib8jMyuR/r8pxZCEvaYdHCa4RIlwL1
/SxhZOh28kk9AUclpa29lTQHzdamarg6JHltI91FnNxXYjmAh2i09ZeiAzeP1O9Cqa9m6Geop5ky
ftZriHudvodP2qey1ORe9VgZVkUNniBbIvgOUZWMAH42Zlm7/uqT3vDTeXD8VJ2xig7IIQ5Xj/yW
ie4AToSjWNbLna+bFn5rn/St5spdDBZTMHbnbGDoYJVpLcA9GRBjYDBgzlLDOYeR/P4HwGucqXYN
MNco9g7uq9qeUmgoFdYdG4AhJFUBuz4CWYVH+XTO581Orl/oT0zhLF/F4EiTTIPRJgejJH8f4t5E
UDTTWJjXKlsjYldIhhc6tETV1A0FcSkzQMzV3U7vfTuCIXljbB0iZzqILdBpuN3AhBXxtuBidsys
O7UVEzFZ6h96lDwWIw90n0ayHeuT0Mcq7Ie4b+6qpSe2jsM8dIHOE3FWdsEU9BadeyLLoN3P+n3X
HeGPBxGsTFYnHy/UGKb+lutK82emyOiDkbkxKYsmaG04Qr9fvv/jcx/5Qq8CCQJlSkkteRV2hqjj
Ovmuj9iR2B7TMOjFDDlKfsMCpIUxqOjOWIZ9x+I0TSxcIiqzVBz+i3KCjMViJsj8ECNk4FH8rtKp
HS+cLCzNdBLExnLnuk2VDzhPgySJbhvmq65lJDgR5DzC4nIwilCzpQQgXF+oNuboUXklHcy4cN7N
QXbJ+QVi7GIyEtb44ATVNB0YJmk+5K1T1WOw8bc4auyKUJo5TOyGrsQHEgszxFNWtia4sVYK9tXl
fGL5SXNLpzgv2Cns1ZRyxwtgtv1VjswnBFqsdAbCNtdsr46Dc8rgdyyCWiuRP6yCP+g+vOXUdwM5
2sQqFa9+xHbBPgFOKOCF1gaqsY+cGf1pykZJA12ilsjNL8UsLXDvqzadx1Px+Sl7thbU8JISRudS
qHAevZvw+gQNjC1tqcp1C2ibUEqw3KBJaZx0/kZoU4hiapnHQtlLWTL+t0cw1lnBDPKKmqFdBB3H
RaaJUsOut25ODzUtwSJKyfiXbtsZaUWHrPcMbOet0yHvb2aE/0nMrVM/yFYyX+zEA8zP6o+U6oM8
8VmDfUBefMunmO2wWaafg4OtDq8DN9WRCpgrEOZ8jcccMrRIlRChsJMeZx0sdfHLf+2bI/FlzmQd
UIuGd9pUGgTutWt0aUfmYjQ69p8p7PIyurOytbF0UAqVBUeErPzOYpwCPPZNm6+dx2ijiK/YeEHv
TPk9IZ7l9kG+U47UCTCpkZNzTOSW/h2pVkE2+8S/K2p/ijc2nRUIbyzEf54BIlLZQ7Fmz3wEIfgW
ljIS5pfXCrPH6LcwZjfjysdEUXFuFbpm5hXmsh/Sd+Rsp5XmPAB3T69uaBjng1+8uy1LSjhbfqc2
Qo+ahpKtILD2WFld85S/CnTeK6am5vgsOVrLNs/S1ZN/5CroK5cA8I+2rbzODYMOCbYrnSbQhVit
U3Ga2fuPSMxILPhshPKU4/Iga1mbNINDvCyJMArsl5Ewv4lsgfb05xyt0tQE8XYvpyrFnOF5BCC6
SZloVjqb6A1Vy6Z52kT8HWcxBQBaGMA+f3UxgW3G0lgkYZ3vic6hepdt3KHTbZ1tPuNSj9OcT/wP
rspCGmmOr4OAeg7VE7QJbGT9SJCIP2TRwAo0+ZByUw7NgJri7RB+q7jSfg/wcNDGQ0qg4yjQm6LE
T49e1xkkQNqK36ixgKc9trNd/U3rK1MDOxoLqr/QjkqAU0ncD7u8JxsB+slUeM50Fn11sAGSFHeQ
Paoc/EeSnHhjHJdl7Fiuydxj+dTTxNUJ/SFHfL4XjvKVlcMM8wxXXZPsIP5PFJbTgRxhwYEcj7k8
Pz5x3NZRVCGkAu78bKuvw18b7aJlP0KAX/3Y+lcqIMg3dBJ5Aw8jHsIqRxGXLVMW6Fd5i2+Jq83T
KnY45tViG7OSLcYSEkQqd5LElxzinPUCQiS9vMcR3XoURDJq4UA7abxe344TaS8lf/FVpvcDvVp8
jXl26s0rRBOedEEgP05w4EOmbxIj6EnD8W0dPrC2PnW1Q7zENeDm2rpeuXQSPmhyM9JUtok2aRIt
RcWPPaOeK90MfjchN8/CV57VF13q68+zCZSBKQ1OJ7o79IUdfzlj5+qmZD+O4tD5iyVyIML5o9qK
C8Vp0/UjJZPJhNZrVnWbKTO9FW2lAewwoBFuNWw1pJMN89rsgo17mmKvs5znjhWPF25yw9PthXdy
+vIFbXhc6jUKGqwmZib84thEVO+wrpnyWtrogSJii/jhzW3s35AU87yYP28b0TYs5Y1XLsNNEgH6
xbbtTZvB/uXT4rdbhrtUeJogkfNts9mUbj/Q//Va66lvr3awON3Pqy9YfXbEJedNRVoRf68dZdrg
KF1XvLqeHjTkn4m0cG6/xrIMRyhi1HcJ8oiG908MExQsGfka3rNYUpdxPcnQCDCKb7NhKqr+eVHk
UB/bZLW2QJId0/4TTEa9Nlvr+igBkZQ+V/2GroC1DGtlvyTpZxOA2y6uaFPAvrIvZBI8Xm/mNqgG
iExGWFaeM5zqZ/446Mbl3BxKcSSeBvPNu+WWzJIBixtNhFLSTKUPa/9KoLXsUQ7Nm0FinR08AzvU
GzQHCc2hgnsgSj3KxrCQ+QuuM6s343/gLjR+mz551EYatmqucQpSPgxXVWkI/HaQMHvTBi+mIUbi
NaDWqLlOiddZqe3EFzWDTVWAdtOsher9qB88dkMEWI9lv/vPMBztBVEOpVXcjFuYLK/mLoGjcm+9
XFiPDLbA+wAakBwLtQvG3KqC9lz9z3WygZUJ4+bEG1YdqNQFPA3vwmrw+rRbSoWsdRjLWrY+UBq/
/+XZYaDZVdy7pm+ml1urdovNX4GJK2oQB2pXEIIx0jjjY+GAPuEP1IKHQuUbu7RLqQGz+XfVdiPM
Bkf4/TisH+4xEwK+R9FjBmYtBxkBUBmiKAb0J1cmOijp55tMeedA6iqB22C7WGzKgwb0Dq7VUn2g
zBlpGjDhZ+m31fJf2hBtgAhZi1n8yj8OW7QtGFkKvnUMPQ8T8OTbDkF9GVQ/sLJfZpa/TnOccE2N
LjFq1rjJRd7skQBiVE2cbNhgleiQr3w3szwfNa2bjGi363vIm+99XCdvvBMxQYyxjP9hHOaxlwTm
ZxjrmMgtVTfkPbxl+sK5AVQWZUpWgwpTe7WhTlJ7NCEpOgeQC6o9O/AED4iOT99dhc2xY0NcHN0R
D7ps3K3Db52XpfcnsgpSC2SvfQdxa9AR9Nxgiu4J5MG5p23Hw6WR3lvUJ/Zxwy32zo5ObBKfRjOg
ICynvutCWCwV00s6DYWcSDELUQoXHcdmlQFlxSTKRifZe525eJ8u0OQLU2D7Wz2qNCMhXWFrFLxo
Yrr/nVKa0aSnGHtFAInZsxGtzyv3G6bj6R41BGEIa34k6YKtp/EtM3L2Haro57KuonMjrZ24WPlo
eyyy51BFVlqchaxGr+Tl6IvIv3WiKpYn2th4PvqgQysNWaejkaMxXDHTdzsexMU/GZFL8sCDmPR0
CRnilYd4eFJneBnD4ohCaYuaa0wRT+F5j2zAAavfPJZnQTDSRKSEG9Hb7Jm7MPv+DdFlq3Yy/Hoc
si+WvxEv9jo+gjzkuB8ifd/YJdgFhQTDA6gpATImwmZvV6pY+KbG04Z9aeepquNd1XWBgUP3nbmB
mY3rV6yBL3IqooUIpWDcnpHs8YKo7tgkjprVaYmpLYRjTkUap2quTRvcsohJHasjCQZj7j9u2WR8
yI2jHaTl8UMLs6boJmRw9F3NF6PsoxOQ0QYleHuUFs88yg3QV+NBccnwE2tUe4njZ/ThZKk7Dq1k
XUOvwgkO47q0Hy2rAz5/+U+hiA0Dw2sl3NtM6mADcbEwf/dQ7RKdStSY1fxZwEGTtrGR9TsRev5M
MYz89ppfZQuoyC+JxvooMh6BBn2frJMGS57xa7XbzFFnqupjHSDg//4OAPr9u431KrBNGyLc1nCo
DkCQQ9qnaol4Gan/eIUB8yMLAcq25J7ZusUhFmO6T1eLY/a/Wtrl6aGsuA87hXbkroQEhddaQwuM
dXaQxTbll8j5nr2Q06/Fzw6gS7AtoP4gw8QFyQ8oyujOtSBtL+6IuI+O3brt91Xn+L8qhqV/GnJh
JFARw192vEDKAsJwG+fh5kVtWtCYMRN6cNglZ9UVYGw/0hSd16I88MjKML4x03vCrpMJ5P63Db25
Wi99MXn2msCtnsi/Qg7hIETKcTRxd1SAh+eQo17gt2TnnaDZAgmKcPhIIH7Wh+ekc57LlMcZL9hX
JLHqeuTTHu6z3Oif1rwpX9zqMThc2CyRR7tYs8+Y/JIcmObKGQnGDBzn+LUl9GQToxbRzq5AVPl2
65s8sR8aaczTWtz2PmoWLDooDB7KwTNQMnhR/eEDgeEEW7cYl5NcEvBwCO6i1Ssw6q69LwoaZJKr
1GbpNfZNCr73+rKxrfugzmJoNmZagg1PB60nr/TxI80CsRMuMvaLDtRa/DPztphVi1HvYTAjpOFL
dTrZbCMyVvUUrQEoq+FD7qn7mU6R1L7nEoyPYhz+h+43mrGRr4c7rvvvtGRLOyov/pkE/yCZlVSV
lwM7SqpiWbw0x1b4sCipPHag98ddEck4uV8BE2iVoW8wDLbs89ZmStJnlFO8of2TEdhE3tZ3t/+6
1WC52ecnm2jzjZO41TDxFGFwRSKEIUMA8EApEGsXA5bRa871M5nWttM7SZi4sBg93ZPpQyD/kZBw
3EDlkMTy+pTPGHAQeJKJDEgb33Z3Lp00nRg4T8pearbQOseob3bUC8AyUOCeYHPGD0KA5NsRdZV+
6JBOKuDYx8v+/zgpZlijh6uVQfb4Km3qXn8xhsn4Un8zXaBatI4L0l1p52l9zJoUu/jd8zdUbDHi
h740n/18twyoMYpasL1AV5mIeQ+VIJ+97BbBLMkWQ8ooKXU1/55Fgo5nTLdAeWt6Vp7uOEsZQsIQ
xNsSayvM7SdUjpY99C31c8sWJ6POG363vQdi49Te0CO301X+/roxTiq5So6NaMeX/wf8T3q+VJRD
IWBPhd+bI33bqzJhWlN/2vWunRanuQ1IcN4u8yGjAnUIO5H3454COJ2cIPxn1WxhymiiseWpua4v
3JNEIXFJuqrfESBh3O88JPr4O8I2fOXCvodcnRcNFJObuHSOaQiFFx3Q1IsmJOLdGTbfPpl7HIdh
lZZd1pQLsuJkGLSsXPkIw3n6/gxTZy1MGRgFiWgKuTwuGCBGx1tuMUkfM100EAG51nv2iVuSuX4z
ED4xhtqWP2AJi0KwpkW0zrt2fQMcpLyiXrOpFSfCflv7Sb1oWh5UoDLdU0Yeex8Ib3Tt3A+UqM1D
NQLPiX84vME3mpInqEEFaSXqfHBi4bSShv4hL0n7geuNIO7qv9tujO3/xClUwenR98FeQdwOsX12
ml/WKUMCz/fwcsBffBKSxHTugUPUcqHTjGHjiWHgr4ShDNudOUYil4zoVfVKSrQia/kijOPwmBJo
rYA1M9ZwQnQveAK7cuUx6hAPwfn0KdTIj4eRZal+QI4zRGZhBDfsqcUNNNYgU0OkyrGPH9zS7uZL
rL7kiUnVzxxkrF3pKgZyeQ+VlPDjSyroxK2gBK/NoiJPgERbAbuPDA1NPCv1PFDiClwKCvP/YHAV
y6GX25aQPFFJ+dXLXDA0CTfrA2rEVxqNamlDWljzrF1r2C1dl6xdxH+xtAQnrBz349pQors+vC0/
v/mAHT0Pa5h7kfJpQ5MVgi0pGzRP2WJ94g2nDnapVHp1VJreWB5K7V7MQ99ov8ElSdYcbEc9yPrL
vN82dpMGct26ilNyA0zjIjs+fSrOdZmQAERogxpG9DOfn3TZGIB/85a5SWUiE4zE1gjZeuFPPCfq
tl9RvTX3MhxpPgDmpJxl3yLbpypqcc6ONV8SDRk2AYxi26uVxQe8vXAlxHo7rUdNcm9KAuL82dFV
NtwrBH/y5AynLpZO07nt1LjogXimUmgVxbqkyl+oqdyEbqpZnqun9xfV5QTQWVl2sYbK3YZL8K6Y
BAFMViXd5ovzBq0xI17Ziprg74kFyde3fgH2v4pXG3IDN0IRddf9+krDZJgp1WYUqEbOGex1Yss2
jAfFr+n2kz9ublXyel7gju0CxIFMfWZh6SjcGzjsKnLCEnzdeGW3TzZiObb7g/2t1ctchc3WiNKF
BYXwGhpMaJECyG0xnummJdFrX3HEI0CDypCxVGvOxdzjYn4iaFNLacekS7Vjvz6ziffVo/sZqNj3
QbAP5mQnTrSa+aHVmMAgrKGJq6HKvD70SJbWYkD5inGqsoxxCPaSJEWZVppZs/rvpl2pfE7oZbxo
vMCdw6Qt1NpaV0cDu9TOPr1hsm/10AwoeNy5KsyiBuYeLQDgqiFgZK63RdH6BVJdh5bq0oUT5xCy
Oo9j43iI/KC40xOqJd0LvLqt1iqMJ/EfyumoZQRy70ecRwXO6oTJHdtP3UZ7l2jzqNe2uLZB8lIr
JJtfclzrFj7+/xU1gYJ1RihkoehO4qe1ZTif6sRrM7RwvrS1sqb04D+EjmqXq/FQDYKyipFyJEBQ
fN0Zl7srqEt7eZQWPhrixNLzzaASmnu3+Ugt3qQKr5G4oYZ9qEWkCH5nxO5Xi5By69HE/F+t86mm
dGh0VBsxJ9wQGPjPW4KYs5KAFSkpTFzLRgSQ9/BaXXQQKrzCnyuSkntFhkjt6huQpxP9EuC+j6Ex
Q4RbYOQJvVfJZFxjwc34I/dB665NA8uLJmENf7mJ+SLU8C7fVdAiazD2QbttycWGQPDgvk1zpLXj
axhFLQEJMjGEoY+KSUY18CwyPD/h74DN9MpWIxcjFkcgUmdL76EdAMoUK7T/C6qbiRoX7jNJwsci
TcUWYXkfVb7Nso+kJR0LhUqq5TEolKNXYDlJqH3LVFcJrVLZlu52iGndUaeoYOAmWaRE+h/pYNjv
YjkhX5dmHs1G4A7GczI/dJ4E9xiiquJn4YmW/2NRmqcAqunFBA+VAKJqRSa5QD1rMQXbpLkiYWtC
qJvPbbBohnZqGa1rckBp3UtGTcBecuCxXyaIV4nWEnuQiQQAPr7c9mIyt0QP5khx9/C5Kg5MEo1T
+hj3RDELGHhCLtfqbxOcsSR8/lHcVuFWiPhtNuq+QuEH5ckgi7aW6dkAUuQlzB2JnnDvdd8j9c/E
BFchQYDRrf5HKfuJc1ZgFsL8kz/WUCloei+MYcIREVHsWDypVIMlAFBuYqMwq5hYdIene7P3r5CA
TcouabgkZOKio4dEnf8X2pBUsNG6dzdtloeQTQzfDJ8mPHBdHrpQ3a5Zj8y+rZapkK9e5O8Mz26d
VOYVHkQ30vSVZqrpAyto26xolkRoQ2tWjHNC6bjjp+vXEc8Y/qW4mqb9TDwK29B2MS5t4B9sd73X
06d5sa1YIJfsfi/eTQ+txpY2nPf+ujiRETA/yGAKFyxaGOX2HnriJcy93Uwpvx7m7atCmyWg0kHn
vWtm9TyrrxixCKB4qLALT3qD2k4HVUzkS2K6nZ5Cc2LsuLqYNzdbAe3bRu3f9OlH04TMj+gI9/5W
KZ0TEHcBtTT1i2oPQuypCUM5WGoMkW5oXgEhogxgVhczzWOFg98aDBBp4ViXWpvC3loHS9UDtSER
aoyuGOQDl2x5Nqg1cRtaBuiMWGnHG5OSFY3/oP7EE+zBu24MQR4W8LpEmk2sd0RfJ8b0B4YrZfWc
nsFFPOrSLYnjn0Mlrr//yAwI4XorqduUa2QuKhWA6Ginzi1jA9fghhx20b/0VuTFUkpQamLDrOqw
EdqFLefd1nyxrlNr6X3NhgIGdaeUy/Ubp0huJxt646GNSnVQUUa7w93tk/L9D/H+TffE9jIFw9yq
HiMJ6QJfbNuOcwUC6K8HD35z6QDBtTvHsD7UEMCVAFv2CMhDj6/zhMdlNYxOV1CUDFWps/TeoT2o
n3KTuAJqdAqgz6voVrBipgNnJ2kOYd60hW6SV25ax/Af7GBS4D+RWIuUZFKqq53LBfirhAghsiSj
GqA0hgljKlLa2xDgd4ad8t3H5wMVuwWeUx77kbwe6wfkXPTYIUiJ0KgdEnWH6xDgkkMJ8rDkQpe5
q3FGdvYTkewziykiVDL1TJ1cNj/t6TTdh9LyLuVJAQhXFLRcgsuNZdLlFBm9zIBleYdHC2wgxGY+
kpVz2VB/rwAXeeO/lLZ0+cF3ZIuuKgHJUd+v8cJNCN5n9qgHKNxPAjKANDnlbrQcFGc02cT1HXxI
u6a1HchMCZwWBy/H8vFJuoMghX8kJPEsgeYm7a50k9vEf3Hv8X4osuEB2WTU3xT3h2vfmPD7K45I
7TsEQ68XRE1JRzd5JEgmZoqU/Mh+iFhclFOBn1mB3Z+C5bWd+iJvYiHOBgZhU1fzCIrwAcWTpYxw
BTKXRDyMZv0f91NIhLSs7PNtj+oU37lfemp8cvMzoLkmbkHqZkUQrgiCYEOGb3D+XWCM+PUluSSd
H4lc966UAxbg4pETAuH0BDohXEYRTPnTS7gxJO4TzsTIkB/nZ1Sk2KFJ2qDnwZAyflzWuMHXMbPE
5LoNVmHQuTKOh7Ka2MVcTImigSNFItzWTNK9XkT1YVm5eYtgh2ync0GtxbuyZqwDAPqiD9MxkYQr
/U5j8gUu++qVCqXfd7B9nCXrqJPsVyT4bEhKcG4WbYqAvrShl5779sEMffT6zDxjB46zTsmJEy/F
GO772diQRL1t0gMF+mfo26RdbFHpGeWnhBnpgU7A3Fno0Mv/lvHNYbtmvZgulwgEsnUGiUX9CGze
jlMADBVYfv7Yw/TpcXHTLxS3AuiF9oDUourS316hlcpl421A9fsK+Dzor9IGg1GfdLw0D+H21w+a
wO4gvGO914tQgCq5esywhhgVOUIXBUlGGxuoZumdqoeC6hJpEYFi+aLOZDJh3we//OTMxq8d1zQ6
eb9hM7c202d2a9HMl9AUtalObMoiPK/ApvwuSNWhEpN1KHArTk6YrkArE7wuyhdzT4l3XjVpfouy
bYX8IezGYICp4m/nfTWISyGCp6uShd6NLs2S8lVd1I/sIoVt8XeD6G3FaIZhbockHX0o2E24yjrt
Dxj/uCeqCv1BJGL38eZVMoH+eYkIrcmMPud1VygDq8qQitHi2Ix9eC7fK5JhnaFprlMea4EuXJAT
gpVuqu3fcR2mV4d2lHoF9OTapv705tKTKDvdaxqmRRCMjp0qWUfFcccLa8K4HGjV5cbIsbkcVfer
RX49kCwrFFUvQfQMls3IJxwFFrU6Hh4CV9WHnWHxK0bnCxNkK/WuI3TKV741uPxb1ZKp/yyOtnFM
b4Tc+rgm1XNiVcyTTvOOykVlRU9i/g3ei4quuP7ck02MdXbHz2Tx5g/wzoKBphaepo8IXXG6a22C
vmPAvo3HpgX4sjN6NSSXUshmlpIo93EpSjk2rKQJW7bbiwCEStgcIISxZQm8cGP0KiIcycApRhRN
mWVeIm6n6xAWC6iWfilEKHLUTZWNe+kWIYB6Zm27dM0nFvc3CtuHH5oI1FItoSnyMyOslGWNHHIB
A0RkQq2zC3ILnSl+HuqOmd8WFlQ/71/k5mXoTO7Rp3e3VctEbFQVrGtc4X1K0QAcjjWpo5tHG1Y6
tT3qyWi9cdfkaerDOIzgBEePb4ZBHCQy8T/eTgUqEiUxNy+Sd+/qzWgNQ3ylHMuobMCeDMree6gA
eA1nMrY4r2Vig3dUf4+rXVZsnBjJOx96Wk7GP2DH6teYXvf8ZIyrV2pJNSzPNjTUxR9clGiiFcfG
LZPeaC2B4thZsQLmjFkRehiOjJ2cP+PsGIk9y7chuuFIqdPwyjMgzPmAGDGmvguz/IJI8HeQB78x
jaYsfNk7DZ0zD6vRaCgO5HicWC802xo+Wy425TM9QaUl/2rNJ4REmdqpoghjY+4yLLjiUN4tEfCj
qzTzWXFacspxrb8Z5V/Fk/0Cw4WhLNhSnwq22fENqgn0imb6TI/2xuQSgw7+skeNJPNSWP7SNvl+
LrZd9w8mPeOoLeG5PPeJ955Wjvj27DGyTjc3laJ3zeCDURC6WEpgyxg0LEC0ibQrL697mUa0Ky4d
bS+OjEAOt0DPtkc1p80M8+nytqKY1rS3Po9JePsECcuagje+7QnmgLNIZwC9Lx+J326GpP4KzzlA
Ks6FmnRWNNHELkDqvkdYiMxGb4TCE7RDBDLTfBGSyGTXCIVLrZj7vdwCESV0aJt5ZhcxgBNRvVEw
I/1aBIAewEjpjxx7iclKL2kBDOcoDye7x8jESXAy8dVe8k1/d9dSstFwkjd0rdaZCUYdsU/uT7PH
5C7mjeBi0MUbThVas98sdDhWJPYutDUC+BYpG9rYfjezZ8vXnqZZL8ZSl0yDgkbFukb0NZwzT5Yw
3KVwtfvAZK+ZH0pPtkKjbwrx16AV5/oAugKZFu7yc6wbQIKNM4fu8cISaygbLtPok1EtcLizVASq
TR9xNXZLNd58jTwGjphYou2IIXHdZuNoVAxfbalZqKutGPKW9kQAhnebhVivH/3xYSEx+6lQtz9U
Kj1Yxzdt/i445GUw4PpsQXxR9GhOQSYZLh1irIB/ie2dVS6dkT70R9HPgsfh5Ic+Dl7Dh5pseYbG
yMv3M8UGLm39/5DR7FLye7MX9TNHJzmyZYxkgEOc+ZRVknmk+WJnsOdiNwNITpLx37tu41l5MqYC
fY4vFE2ltZb36XWqdSRGNJMz4QIaTitaVyMUh7N+82EaZG40XJMO4s2Pthta2WEl50DEc1QFgZuu
2/v6EDO4Gpv7puyFWIy/pmsxUzz5w7PezAmpCSfimgTxE9bFcLqqkFFJARgc0T6+zNWN3H7cZr+f
V2hdGV8gNfWKFkjKplWig8dC29t9LnbIC2kMkLE0I3xUucy//n4f1yQe77So+ZbfzGnFhP0JG+a8
rKzQt82b/F/vNlvWtel/7F5M/N3VZH7QJum4IKxOx4Z+9XWXQXMlWIo2XU0thgOz5I3xOusCxHk3
6Kg2vEPJowacxroemxtx9HnM2RwE4MzcRzsNaqDtVUQJqfz0NgfPHYnFfv3JYWXCC7Pw7l0uYMkK
/ioGvGux9H+7UIOeQWdkMekr2vCLXjtQJPcHD5IB0HnELbd94YJ0aWlNGocSBlqO2PpfRq+0KQUN
uJqQ+XpdXaqOGkuyhagli6TbVbWKEQMMYMV59hxiDyj2rTMnasIgVFjJNyCxxevIst+CeuDchA11
Spgj9gGXhdl2iHGlGePHmNacrqljMh/bZ3lgrNU13WuXNCyckwWxj0p8p/MJmy2ygLPwb9qTID2x
iLAcybOtNV8rg/UjpRRv60EK1RXsJpTaGiQS5xwhZuOkqEPqQV15bPYCI+0GaIxV3Eqv5NFI+Pn6
/qcjT76s1fYw94A/iBnQrzz9eVhYioRdaMoYVhLNYQM17v8dDmH/HJKf/GSmXgoZNJb8kWprJhna
iR9MidBRTeem9MWN42QksFLIs2X/gRjK5FiBVygn+p1qtkXmwiAGSnAObxcn50nmyGcn6h4DD+I7
tIVwxlRbVL3L1M27rB5s9FyiFP4fJotKz2JhRvQDgTKoaX6LxcUsp10XTG/jwtRHJOIyvxvdTqX3
lJUg8QuUGBHDhwxq+MaCuUJFu8XjuMHlXzlMjehWpXHebvuqpsWwpacts+yo86zRxcdjJQ0b/t08
2FN7JnKbhAiPcti4tpCMfCFR31XtDGqIrPOWPY9qnoENN9FIg03p/Eq+YZkr4kkEUtYojf4d+hnz
1eN0/2Ph5jpBU+nxhCeWQcftbc70jz+4MUq6+yJuO8aPqZPvdgbAKPbkEXsNLxk7F+O/QXtOVXCJ
AjUcuUt7TJLDJNEDsovLQ/u8v/+F2rldT7F1lLGirJDDgLqQQTrGlUdf4uMMhER3UnZeG2WNO7t+
cf4L6IZQunyXH48HMSp39GkoylN/hjCmhYHeeYy/LbllGnW8I15FdFUwAQ1f0Qq5Lp8+Afj03Yt/
8d87+xhTpyoR8qV3lkAPFNiCWo6E0bhD7bUN3C9zSp0Yo/2hV/MC0GSbCuEY3sc7FVu9f1CF1p6b
M5ckH0dqZZr4uiNn+q1CJ0ai+VypVryP8RIOXcFlmOjJpxjWeNxEyq/ZUHS7svgEf0LC12AXnCKK
X2JukmVQVFEnkroqAUagMnTnMU4XDtzN2f3X1R2kMXpt9jjUKJWkcrrVyo1kEvjJxfBl68V84NM8
MAR1lA7aoC9njMHj/xgyEXKNsGuQfJrVPQMcRtbv7sHazm4JHQHT3waqSquGHNsAO5yrqRUJ4ODG
XD1/fY1AxN6z5FqxuFK48VkxttD/ntPIYcBGH8T0g33BERnR7n5NfbdLgBBT0DwtWoBCU9uxWF6z
vYGVEuXae+K7vZbBVj+UyLcvm7shPPkg/VarQUCmYGdD8vb+VRV7/VndKhLqYJEATOK9fvF6X840
C128Ia2xfhnvJWh4Pw+96e2X23aFfGL9vNkhDdiEH4LD55FgL683J5Q7rNZY23CmWdV3uFE2edek
8n+hjAozatulc9sE5ajtyzKkB1vAjEYCfJy5d8CM3+raUvdielAxbgmcLHP2IPKIwr1Qf5HqL/O8
tG9InVd5PVeJSfhVfo3qJXK9R/j470+iDc4WVE9cElRFYYG0P6ad9LmhPNhiflhoKSAMBEi4HxpI
kvcg8MMjEOatVPWYB9Mn2JJmpOXi2xLcjeS31Tp+UMgjlVKTTcnTByLgENTH6I8yhFqKPJPM1apV
nCJD6J8eaKZ0FmmCKzg/TBbx6rHh0CJJ0fT5tPF6fRo3TfehH+94hkazYdxzm+DdZ9OrW3d8ay5Q
5dq9g6xd4a41wHNJ8xFn3Uf65WBkAupvWsh62cdydsyMI3rmjpnM04JnL+ZHL6bl0+ehNF+sJo2g
tBg+kyawIvQcjKfNUutLT9yrl0jJSa72GWi1l+oLqPERJ4MV0diUTYrmppn7B/gDpgEHtCZBDcEG
rsXtRvsGZwjoRGxjEY53lvmEbIOh3zCWqwKhrvsIKPAoDblh5NSyVRJqhyCDv32EzFHMMqU93Tv5
r1LWVewCIErfi3FEdqNuBwaiyPPdEevSlDwwqdejYFLnJMvoE15IH4vx0N5WBZ1vM2jh12ztHzhb
ttshc98NSgM+oeaD0JI79fBqI4PQE5auY3VBc9S/E7GxDX5B/lOjEX3cLzwjv4uZGs6j+CLpvaB6
Vn7IhaqoXpCnHs6C+hXPUrc/kTjwWrf0/khBWnUhD4isgh3p7uhKIlz/LlAXIV8MKWvm7Rx2mLvs
4eC9NpFBMyhEDCkciTCSO9qnRWufqwydwAZ+73ajreq/Ay61Lfp+bLa+Kc2C76EDLWaXoHYyJZEy
spyq0sbCkUG8b0VR8XFqWRFXZ6SghP7M4x17wnJR0Vpyg1rLG5hNnpaV0pMzUfNXzjNGSd083A0a
A18WwtD0T8ptPvDqKtmdg8g+1VPFCHlD5Of4P+TsLyDIX/V2ZRN/VfgsIuS3ALq+9AhuWykorhrr
GC/itHZGKLIlXlKu93d/BgtekkmFJr0bb07EZflx8jG+xc2n3paT5BF3VAup9BhwM1WW1s+ghlHk
TRTCGy4Rwh/Qlz+s2N/9dgb9ItOgRuOsCNzo1fsOZxEuuTdWop04G79b3kceBtVeW7vu3R53Bwjb
SpE7KdZPW8+XPcMdlDvlsZFPeetAUKWMm2q8fVPaEhAXMwoyUZKWZZeoMmmRpLjm+Lgk87IOSXYN
TvPZAl+IGCSCPm6nLdi3r/Z7OkVBjDW0RAzwF9mNeFAYr6fqNaQYA+D7xmH72SttpLbErCIXvKCJ
T+x2kk2X4f+kkG+jhTjr1+J/h9DbLwU8ikuSVALYxp2uIE5C5cd7FpTndo1yaE5xCyOSYqau9AUL
RPhVXk8Pjtna3Jp/KOE5DzeGI+diC4A4DKY5ddkwTJSV6jd0B9UhrVtz8xkPFQjlRGVcU3tFJijz
9TgqhZiMnaG9prNzoUilWkuqAch8qHycqrolvbPPyr9viSPJG5JYnWnxc7vJkZClOIcwUqi5Ho/I
CASiO0slU927tWe1idJJ+4x5s1+sLSTuXkqX4JF5Zs3bS8zOKmiKUMeNosk+mjxPgfhpFrqGvo3c
H6mHFPURE5OOs54SWSirgWgbNYmBEui96/r6vzSy6LdfrSBAPSAv6dPm5RSXeReIc5BOP2bOap0+
vJG1WvB7m9jFXl5gHp30a16iJSOEuIS55gcfSbHLN2awiOdefmeItqou6eycThi/XJCTTcTHXnAE
gQz6ETuf/E0E3tk5O30awZYm8+x9LDJH8oQJsVlMMWe1P9PMKfIMawLlweJKphJor5cM6BvkYVMP
T+R15gC9LhzdOfQWfDaw2pvhzV2/VAekUgyKx/0QvmSI8WrMtgHp5S0NYUR3sB69a9yr2hFJyTpk
sUEkv8GMMrtLMXHAucS10DBJlUeE6grZhv8gJLhrWx7a84dOd2k6tNWoieSjZMWDUIVflIkMJXSF
OhmU6LgKIuH9AsBwD52afdPtCLzo2rBcCJzM5Pmiw1E+uCgSjKQEMCFOtV7IDF4E/pDC0I7zfJxc
6G/9mMjqF0w1jbUpqxOWiFTW0uKWYC0YrRrk8r87oX6f27lFwW4O6sm4nN3u/qn9j8yIplEOZQUr
6UGrK23MmgnS0jJMf8k4PDJY0HKd+xEUkFbgDmEN85tBXYzxxFwYoRH6II+vb4aS8aXHNL6RHmtm
gmEMSbxnv7Zy8/wDv8BlT/rjiEsEZbEUwme9vVxcI47SlNd1L4LnzUBQkCGpXxHwrNRm1CZQZsoZ
XN4rrM2zadq8c2mdiTM+25O0GlGDwgjsztUoZHYCrPDJKQIjUDFcfaTvDWRgHxC5e7UBbgGRPeqs
J+cen/v6vjbIFLCXonVDkDRShN8kJjQPwVp+3yKt8LuZgZb16pRBcE40W6ds6e9h13/A6/VE6Fyi
eWYYObz9FtwqcyjiC4p5se41FvsbKhBvbKlMo29RyvHiAiuVKMjqTDisU+KRQ1ySWstrwDZ1v1bS
u9dgypgdEWwF+pmcFaMrVgrSBHdHA3pS3cONjo1UkIPcVN9idC4i2yjMTjCQx66q2LjRQ/rlxmTU
7+BclK5P5HqfcS+h+YzGbmE+iSf7mUXg0Hf6kUrl8PjuSNQ9uSkFLsqETAymWloiCDDj0PNZ2hso
wt4cORESifdQXyPl3dvVcan5E5gDgnbTf6/uTw3xTc3n3IkLao/UsQyZ814CP89BQkR37gtjRfDm
cxGRFXDBPmtob6KiUGH9+RJzf+L+sWTrS669i2PyKg1EjrxHK8+j4tlMg9A6oZx8mQ+52yVVEDKm
N+qPS9en3/G/poBDkrQ61gM7sNXp+YfIgIqE6ynAWsn3uX0UfrsGBKiuD1krkobDzs8RaR0kCYnv
PheX09NzpvJJL5159gSza/lnqjH9FOTGlVnZTPxF34EH8cLxV+jc+CfE7huKdwZlDE4DALst/Fj2
esA5pWEaGhlRZ1AZz1q65P78LK0DW3M2owxHG9aOjpemyXOHXcS6pwuVgcAOMgoeZpJOA2SayBzN
Fcu2OJ+xrJ5baRo+F8o9l2Xc4KdFoj7IRrdoM93h3iRLp+UsyZbv/5NL0MV1SDsEg4GekwLDMB4g
N6wmFNrzLzetYh9wgDJ6yAUpSPOspvH/xOof1534fOYIoiiSqlOqcNJ1FRxq70xDmjjg53HDDj28
i6ZGESswYM2664oU958loUf4wHDMbsudU8a8zD4NaYb9ZQrKSBpklo8pVkipxNTY1HFtmBoySf5G
ok2+mkr47aQ/L/D8wBh1WKDdhaAlvLqDpnFl+/zrsCBWBjtXVDGap6M5gD9l6QaGGONN7Jggw320
nuAzPkIncLQhvMGHtyOuieSXTzPu6j/QefJzFdaUQHRlrB3rnO7ZYfd4BCF4ZGVH6W85OF1ZrY1e
uZHr9dgYI7afQ3AC2BC3lVYSfCnz6dOJOLQjcYuRIILiPyeUTNJFX7+ca1xRkLCi1mgASlIVTMM0
oww9ACvs5twX2bmDYO15TmmUXQSi0MD9BmgLui5+Aw7XH8R66hjzN+9EVhufV3e7d4Akhyp+eI4L
HtVrOSkkonjowpkc4nC3F+HTjWGJL1DbtrMOC26n6OaKt4zBuMyb15UNM3jIYM3OjOFZZz9lMqpp
aiYVYTxQCGPHvnyAAbwbBMsORcLTdhkgUGl1/UbjnnCY+mTRiDTy2UCGaKKgMHcR3sH+CVAObeDg
7xhYu1plxBP+zUmugfHQPAICjG1GhZO8R6vfP411kByfwAn7Yx7er4TxyMHUJnOKK5mXI7pzVNFu
kUJKlqbOkkZygM2c8FaFsEZ3W+Z4fLHxVZdMBAkvMYktw91zVOa1XR/vS7ITQPPrRfUQjg+Kk3SU
1zCLcuJXkNPxxC4wIZrehP4agxfQJjg9vqe9Cews9himQaZWGXsEohbadjq6mTkPB407kGF7QvX/
yqWlYkoWV6Rww4hLSac8ZR2JNnKIxyqbQOjZkDrBkZc92il9WASLmmkPnofb6FsDbJBsHSyXV48A
9IKc6Rp/serpIydtYB5kR9eYq52qGgTzOFC4CNfaZIJVr037k+61iGvJpFbIf/rVum90agYY1yqX
B1P5UVp7SORMq5CBfJnxnOF/LNnQWoViEENVp0vjCWLg3ZQKqibdaL4AUY4RE5LWekn8qj5EF5K0
nk/V7RnqtaB7fovwNsfs2YNDSnSoHO/mYUzh7Ybi8wNu+ttl9P/p3hOlk9qYl0E7rMz/kdAujgXa
Fc5kMbr7FovWh4NaDkxXIiai1sL740uVeuZA6Jnvc+/UkUvKy07qCocXtGvuUv4tXEPcVUd/kfR5
1T5SSf6uemF3COTC+XzgvOBnFLwulHhKQhs4TiBGZul2XgcDCq5QCOK3KwIKSaP92RvkLY4WIa28
sfA3PA8ML2s1sSEkNpuxnDyLRh8qpeU6WTwAitbS6S3VXJfyljnnivelF8FkMqEsBMGPSlhkXtd6
uC4tKm83WqOe6nofZdeSjPr85azrJKSONGa/JOKwLn15P6MUyvX73ZN3x6+uF7BhbsfZDZK9Q+iK
ln38MphDKpHRx0OC8kBkNuY0ae4PN8o7uO4EET2+NGde7BcVvJWdiEY+eLhhvI88xOX3QYWlDMi4
SnoWEo+LjVyexyUCyPfcn5tueWev11XTR3eYBMR5fnJMUhkmyzOvu1+BpjYJgc8oJmS5KLk0i3a7
ud062gAtVCXkPdVg8NSJll/lLWFjLIFjR61u6KTG96E5OaGH7Tgn5zdt8/sAur1e76CQBlknazW9
ozeMpVeTqy4B4XFamivrgR+F8dtBuvupA54UI3raXV1ECAOGmjcZjTW5LJpM7eyjouW8BOC+gNJC
h52K3xaVvGgRpwvotC9u6KThc+1+R0Cgg2UzZtRBNZ3+yd8qgVxjAW3hCiAsG57ODUrlySrQMtc7
xIm5dodwXLWWVtkSO/mc8UDsIODuavWF6ZruTnp+3kvuhXzfJHNy4W/0atOfVhgcnQqWB7p/ChHQ
VvkEcW7E52BdQKhrxHb9klvTW9nHjVxZRN6xUeuSEPzNAlCIVELzn80F0yv6CPpy9o0U/lXUW5xR
+d0FpDflMY0MjeawnfqHZpeYtGzLtbJPEpHrlQoRHCrdoci4gchIsX8ojHTbT2DssfmeRVraeMsi
I6D51nN5UeHCp6FPvPaHN4QsI2slQn+OC30oqEBipFRYOZwwIZk7FYMHHrCAQmlAJfCJpcyDtaYh
KhxL2gEUJFoYijI+RfevZZGd+0TpaO+KssKpX6i2siVYOmZXdYCbZoB6RSC9HFVSp4I34bh+pN6Q
J1/4/MyQ09pANeb7srxIiw1HeJnrSHBIKkiqk5RAsUHwpQ3pT12uxy9r2NWrLGv9ACCdkh3Mtxb0
HOHzSg5Fp6gDH7nV3kCjgEMmq0uZE2CcrLzU/e5N+iJW/ltr83ck4ubQ0WHBaaEq73Oj4z8FMvAb
M+/7VdbEk+U1dO7M1c4tgjduwEEzMqSN3Y2GDbYlZeTi0RTHqgh53p1vzg5wi+9JHhYgue3Iu11K
EdAUQe/o+BHr4OMO07nAYmX9CNoza0dhCtFtK78T33mHZSd2uP5qEztHZGRgqzVV/mlUeW4Q951i
hWY/CunIXxMU6Fr5E75SkoSRYImf0MnrE9vwjLiqRU0gnPOjCDbku/FJweuYJ6tUM+qzDCPO40av
T3BuJ7y/dqytHgirRTVeSGZiFCD5odYapWmGCzNDaVk1PeoW3QwCTJkyBjkFoyzGrwXidL/nYY7c
4NE0ZaBkB6BRIzxEgnQ6DJAhIAGMSf3A4miiIiXBOqrcPwVF/ooegmVNd76fEiN1u0JF00oiFyRx
ffA7Ln+YGpfWMgkvRndaC+aBpOJC186oxiPtycj91NkzOem4mxgBN36DstO91SHckdpwazQi31mH
evqx/ievCylPLMdXIYzLKHL0g8jhOdoj8Ph8rMAJH/J9giZ4VZW5LvLGWwEMFyrz3Cd2I6NtrLJS
BfrJ1SzOKomuz8ZRVfzaffgXgQ/jyEYU9D8X9rqFnxWPQCe8SfubAZ0tJ8vvEwNggYYuY11aLikz
KRYIV200uWgpVksBq69KXuUlZhDcsyPmX67Rs32TeQjPxmWEjXbwO0R9aqxiwY6bY2f2YNgptr5D
VfGNeMk5uFF0kJ5/s7S9LlSi6qYj4lgk4Ey4d1li6/l5Ta1hS7r8t3K5Sh7M0L/dwTjOOno2BX1w
BlhSxJaMn+Zunki4PrWe9Y8l6rhfoBDfGwY7cdUkdKCKOr8+kbpuCOzacPSbFKZ+Zt2h5HhCcT9N
50y3V4GfnoerO5f1QABxnpVkaTQFTNKO1q+PBwUlxySdP5YojwMOZWKz6mJTd2zvWbngrMjpHWKB
8x3nrXXcgjan5UZSpIUzS/X7jTtrM5zkdo6UdpxdJjT02jNTZxMC7ZvNpWjQikK0xEPbdAYwEeqC
lFLoI6FPKP3onk/7VuUehDOfPZjmwxDwcG0UncsnpOWkGjxiBQGg4APi9ufEEipt1Oqal7fo78B0
grm/E32QcNDVCI/VhGIEZt/LSXkffmD8HP/qelYw0heDfUV02qZGCbCw/UaMf70uO5nl3uCwF/4A
UQS7lZFTOu0f0+bzC5ZgztStjzK8gQcuyWK8i/G3D0+O08P5eXwTlilLS86cVvUKuLTK3FxuVyqS
R0c3mIcv+nk6L/T6AecscBSFhaQ/HiuJbLDmXSvtGd0wB7Kjgbsos3aTD/JfFjAeEtuqUDagOeGn
Er9YAq2QLLOnuNayZCLdwAu6sU1XH7fE3rnKYzUP2CzEvRxeb9Jd9Xws4ST1zlXTg+T86XpMQfMp
L3r2qMEwGmBfITsfacUhachOAP7tQEZiTr20Bht9EvZzhh4RluAVTFaOauCKTHrX7DCtPHYkTahd
W7nHWi15qbNgHBtheUqrABv4JyrBMuxXx+odJuE3mGmhLb0xAF4Hz3HuSiz79ibosQf+l9dpwvZy
ydWEUPGMh5DgBQQL+jS4KBbc6+cbLVN3H3L/2aaZx/qx3uWxJmzDFPbD8DLZF4G+M6KbP+3l/wKf
OgvcbbUxMs0dc+FHGIcPpsbHNxDIlSmeuq4cfykCCP0fB7kD19oND3zYCnITL0j/P0pQr/PxJssZ
4vIjnSa6E/spSXvXwV5EUMtUpOGuhLM1VEjqEUmTmhNAkllW+/aLJWzUdCGG8AbCK58PP4BV1FgR
XSqcuQhV8751s6ebPNhFKlyG94w28A28Zq2TBm/NwEQhjNLB5WzTnzHAVKJBYf4D6PzItdrkprzc
Nt7QcnE39DCIHsX93w69qTKonEe78SvpB4tzb4vt4u7hvSgUfaBP3tsGzK0SWgvj1DNSpLPw5TK4
PN5PryzToZ/ZE9jA0KWNtErOp/MfZcW53grzSmvgHRSb5sR+oQGD/3UghZXYKEmcG9u3d7C/KOGE
9qAO62pXL1cyl3ekijoll0oWydA173uQWL1cYYJLebrJe3qCFRzNRFIizKE9sf3xENpiV0Bg7YHH
Gn4E37yrUv8E6St3ioBF0jZ62ClY8t/vTVB4k/SGrFpEQJApj+Ds+2VVobhQLetRg4o7nhQRnJuA
K2FoB2yQwkLxAt5PeylThZUuPHZ9Lz7S7MLOjumfrqEaLD7bZgRRsa2gVAIqcOaavKBOOlTmufHP
El+ugtUpdQjAdcmhwb2JY02rWGiBouMt88SjomnKV0sdKCxOhRShxobQn6ZPff01BFt5HDLtLAHk
J/9Ac/Pr0eW4j3OI2/UuJuA7FIu6zk27NPyWdID1qZc787dR6cmLjOovMNvz7FFTYDXM7Gj7leqs
SdFU7Rop5nn++DbRWjQFkplpT4pYoYYPZoGXdiKO3T1rOynadThvUapmauGHVRS2UcDjRj4G6brL
3N0BZdX92Mic9SxA2sssRNClovRjEuBLpujVImHDeL6CJdPaFoV7uCscwFEZin8d3EEbfEVgjvxk
FCKFRtXXBPx/DErgGYn2fvboy+Ema+8tRA5MROzkHTJJ1Tuc/Z+3O3KB3Mmk0N0+OSERbB5U9weL
Y1ieT4pbwYei4QvPaB8PJcnNN01G3ciJNltbT07Xm6gkb/WYeS45ofJkjIO1g0P9MyrrXxOs2Ulr
hJmk8q7TRy6XQVGco9QaOzXXjQLkX+yPhxJqNaXj29V0tC80SR5ZgjPVQPxZJzFCogofb5BSJLTg
wkPHHPE7Hdx1GCVjz8UU2vh724eKC4SYNujpjFMGSZTf9V43mzoVb748vbj0TGD4sJ4XY4ux7HIB
MpzE03JSLIwSBIfEX4DkPL/1XMxNG9ZGi7y7GVoYTVbemmpwT3CQiutbA0NNSZoJpWthGH+nB8m/
/PNMUkNcoN/1kfMRYJeJG0pd6sAn/wFRnm2+ViGQHMY8MIrsl8f3uAOUXwtNG6m5JKHb7RnwslvG
wjwjpj4E1wCQBwV8zvMtMpExhelWmxXdZxMIbJmc5QqyBRTuyz+ah0R7sO7wSqJXmsw6dxjUJz8K
RDMyjFk8gy2SuwrNRvnXm9fYO2Ur67FbrwxHrmStHuWY9TcJdDGELEEGF2wXN4R5tGDBmnjdlej+
dTC9Y51usaCZlsZsx9XcizvK1I7DAfWaFqohqTOlnVoMqeTtEt6Y6rdGmeJVKyJAk9BfOaWz0bu+
qIeCeThT98TCO0aFBt6BC4lv78BSmutti90fQKGSSu79htA7+ZYWrIemRT1dZNPIMZj8ZYSMjBeu
QIHuIhIub/WU6wMtM1bG4QInp45wkV3NjW9z5JPSoabkUzlQ2Pvm82jEVM512PDeTRB9gm31USf6
6qDmgxCrT3fufMxugB80zxzYkQLGhXSUkzDUMve3ke+qr8d8lQ701sIUQ20IehJPn9nnJEx5NEfq
e/aifBRbMXKV6/v1/r4/lKFLxd3ii0p3hxYjeHiGhFNRbfHvwDB7YQwseYIGxugEGOXS98ki73dl
Su8PQGpm8rayWeTXeCUpnQICCioV/9pcKc8QtRuMQR/LF5enh+yoBnxK11onmZ+z0VcIq+H6KImC
fr/iyCUSd2PTyPvgekFk5bmIAxZQO3a1+MCGWDjQYudDYM2E0kTo7nwuooY+rSNPoajm6XHsrz3b
RLxda0nzKZ5S0RbhSGds79drAgEcun5i5T/O3wsy19UgZqKNX8K8NshiFhzZsxKSWeA7CAumw1wI
Jr4VSzKM/ugDk2rHvewWwfEhK5uK//jyXsCvyc2kjWfZsvLhRIXiw/qSNiZUHR5C3nKtD+yKDNXi
ctIJFIZiWDWKS0ssf0bq3nJpG4zikYL/1Cr261yoUhUevjfvhvKdHkb3P2PtVf7zbnF/y7W776QN
OX2PMI65dHaYsp776Bud0RXaNHc6LueWbFeFG7ovVv4sfqr4MVUNrRLM7o/n1INEY6hoje2bd+lf
lOHKmEeZGpNVfEF1cBql0XmzeIbsH1sH5eRArJsBHcdspkAQKyeLJ2pe+0LpvgUER7jkRj5SqHOc
Ro3Tov88iUm/i4aChytIKHvaB6nqBZwlb2D12hPNy7nyZ21X62g6zwsXUHkSbsZbBlOajQKYd2s2
bKtoTwcFS7Nl2ES0vzNuZBWfbKkLXdJRBSpevnNPiLZB09Aye8oWoKxldK5bUnQ2+ac3VqiChpU8
s4fPuPZQm9OqblguCaLFeY2uzMPeJrS3YVfXJV08CGjibVnq9KpEyB/gLxWMKXqoB5yI6z80GtXL
msu2DAjL2Vcitc8pCfkMZluJPM3DBgMBKuQ8/SpAot7Fzd7GQSFIVuHXMPueN+yWcRwI+G0LSVqr
yzbGh2MJcaf4LXdlOAVVWZKXTvHhUQDHLSy70ucXqDfIV8bao72nJrgk0qExFhjrJNt8tQS0I4f3
OZTEC/nZN/hkPISmqP9YAsmjn6274W7jVIMWm3a+aJxrcAEcLfRSTpjetaF9BfzYFaXg0FrGLQ47
8gc3q1BNM5/hgMSKTXMQOZKazb1pSlUGzjDrAc/hRnawnVmtonbt/JkW3GDYKer3OnXip9UzpgjT
i2gmmTwtAa5Do2FCVjg7W4zOLE/yEOHAE/O746CWjppJaTJBAvBUL++F+ORHRtboorNsteSVUaEP
eiZricIqCsrCAae+gwHmGLcnup2TClXrU74YFyrHDv95Ec6Y5ZNWzrTt/CwmZ+snXFrwkrBwGbTT
l5Jy7zisLR/kTNkNV/EuNtkzz6FJ7y3tB64sZ1e/FfKe4sV5cDZUJtvhW9xeMvEPbBhUqxzi+Has
sj/xeBDUNrrfnhYZ8Y11jAy36XTC89nztXdCDVXHUYACi7W/hbMrVOjruh2pC/LPqquTVhKqJvML
uu2Dms+2hTitCWjAOYOFT8GkoRAKw/WhxlrKjBEcHNA6bgZ5AZaabU+dzVxdOP7Zd1b+ienAiG+o
nSX5byv4xxsi7kXx+FKgefEU/5n64O/taXUC+c+OWKGY5CopHzlkYeZ4o2BBDD/OLoZmG0IM9bvc
PvLz0/UcHogid9x6oA1RiPSA0dQtMaTUzwQ1Shp6ZXUZbpm10iHdaPekOhRrO+MK896aTqTLRkVQ
UrdWV9tiBaXuTLzE+0O5o2dy4fBsPaOAZD1R8lct6YtKPL4trAJ+wZ3QdLhT4AcYlvtq3aKzK4pD
JzEkQqSJKZwF6UpR5l6Ct8gWhYWWDe6hkEtHfKpgjVkHkLu3udDAsSbAGNyj9PuaNNx+1YsYWI2/
yAJ4tXk76V5beW6FZYvIT/PNXkFUzDcKZ0V8fGc5kZFj0Ux7gg20rutaiCCME/QEuLOqGVPC7jMI
3Iq8jIlM3qWVDHYO10nDM4PJ0Mt80LVnCXR4uN3h0iGzuiji05/d/NtEt6gB8OYrvPwdQfzFhqGT
9OvpAll55vA+O6yZhZEdl7g6D2eYCeEa7zzKek3yC/WewhS40sAUtv1HC0DsrhyTft5Qb7+UPR3M
ohCS9sqvrULwabrYbfluhsK+kYYuzomZIdBlNdnt4UaBnlHipLeFf2NvpvQOS2k1eXROGofPGNWi
t+Lo4rae32KyqpSDtH+QXbPyTKfJMpWRTRbsz+VRh+LqzPu5zWXL1GcT3QpniaryZF0zRkBO1WwP
iYUQGbxQqWiIYg136/WGmNT6A+oabWOj6turjntDIEVvwpXFtlakqPNkIG9jaFlW+pcgeNyNCn9j
eMs4IVXuMqDrSMcKaLSRmb6+E/nMoj+ZAvHxc5I+j/7zDLcuwkE+L8SxnS575LvNnNmnLndAbg21
TGCDhthj7ZHQhDENqQ+OhKXmFOlQnWFpCaWM++F4unr2gnjv/OHG3TkFhm7aZTojehy7QIGfUoCG
wid4nzJVDrFnVxfwk2r7RhGGT+CdniEr2zjr4RF0xB8/Qkw+YPpbul3JNZM42APVp88Z+ogu6qy/
MqaEnDKuPsFnAjEjGnL5A8+JmDjbiz0Z4/bw1TWW04vSw+Qe1R/T5CFNH0XcauJXGRe0i02yvYS8
zbMWX2exhLuijPty2EH5QwJ/ENbxT7qoQUb2MsqXmYhUtqpdIMiES2Gi7Ia41x8YgwDQQpLIVryr
/lhEBKgOxecaIFn58q4ix5VNzUOlZyArEMgSCZIAhIFmTHCXiHcGN4uo4rdXU2kJiMzPA86Yjr9H
oQLXJ9UHJOIV+kRHAesZe+FWetCT2cx62Y9Pt+DZM8BB0WCTEIrBuFpe0USr8hN5+N36v2FLy5kI
K7A2RBBHcSyNF1rWE0p8DFWGhCMzCdOx0x2GvE4JHBrD34pdv1EXH8BChLYFGBHERlWfm7b3WgKX
VyPr1vhObHv1AH716WcisGdPbjHl90mPRsH9b2CoeOFJUPIzhXlcp2X5v0x4PTDX+izwLmErBWzE
SWcYHRF9W88tP80/6cskKoUq2Vsp9nEMjEf07HurX5fzYw2V4LPvqZk2ZI+4cNp2bNK03v/QXywd
SOI/ylE2M/gRWdCgb3M1W4fsdgBaa6/M1d0KaeMkPyKsXhrhv6Ypt0rcARUQ6GRhrhtXnU4F3Y3k
vlZ1khKnAofLTpzn3uT5cUdiyCgKFbHfhbMOUIOF7M6nOC3Y2OSRRVVrqzgKdYyXASla0FgncA/V
lSI+j8vT1+2TljC/Dwk9615MhGXPB1Lj9ZGLhFZ86IR4gmYnsVzakmGH9r6JLin4LHSJ6rX1vzdH
vaNlcFaFLD6Se9Y9GmYOXXvkFPpERXS04w5FtktxKNiegmebTQ5gxmluYYeHINputzKAVEuVN9Tk
mEczrfSSg7AwvK4xw4TkINp+1nVgZ1oVHktYuhjXXGy8iRnNBN+JyXOALPNqQExbxKXasMkI4j5S
dy9OV9iaHWnNyf7Lkj19ezQXXVInyH7+zI3Z2YnOHyN6yxXx82HYgP54bqh+nreZUDzbUMDm1VsE
sVqHNAES6YS0ute+Wqg3om/3PSCtKNlAClF56nYrmGPyct+Wrrh9KuFuzY00aitkkXSjjI6m67nB
OKz/+SOKZytWUeZqA5lHbzGDzKQN8BoR6C6sr4qk/IjEwCsXiI2Xu8RrEHP+mRABMpXggUO7OvCf
+K3e13muArsCbkNew+HljloYOhAVcOrffjP8Dp/eOC6NufpgnT76bOas8bzkXzt3gPOjn7ln3dam
JR6KQxrX0rzWVncWXy39tSEZPsBTMs0Ot1aVVgbHpFeRFU/UOdd9I/1WEKtp4+//qwmZPEQuKn3X
n8q8T6D9mILIsk/tfKACJrPbJ2q4xlTal+n9pVMaRLgqGHzP5eL+tE7oj8z7Vf3j0jyJT8xzZ0ZL
KgQ8BH7NxSSubkHLRgJwi0IPK1piUP1gITR/4VBYVv9pI6npnX4HNqGGzFxCGD2wKRmutSIhjSyi
pkTNz6/ctaoTqPFvqeP28kCpfXY9rOSEK4DpRBt+mdD0PBh+YBAPIwlla2qK0EZt60HxH/c/V7Zg
RuFbaikHG4hEXaXo0KMoQi16rUP1cTbpb4JPBNH66Y3fVRlEruiwd5X0uunoDoY8v0AuB8JIRKUW
ItrOONaReP4mCisottbfAOKX6ejVKD7bVDdVaDzbomGz936Laar1Zuj15c1CkeV1c8ZZUQ7fdl0k
emLyLtp4Itr7c9yPSRhZ62B/YgHIDt/iiuuJdSgYtcKd2JkAcqT14/MKdlQ8CcnNY4FkDNMyxvAo
7klzMEqldzxiU1uX89UXEiKl7POAhvuwHnjULiXVRKJCdJgBawDxeg6i17hd6uV10+BEwc3qT1W5
ptLgJtBbytckBa/zvigEPnqM9hZ0Xl+px3ZG0XBUmGFn2XK4CcYzlzCzyiVUimcRwbJsN5INXZrK
hhg0OROXL0cZNTXqO2nJA+cPs+BZKYAzCtJckGys8ksxnUiXZp+NM665vH3fWnPuG/HuIEdu6j7o
V3AQ6SiNP48yID5YhXIO9jxJgkP0wN8fO2c1Zx4Y1LTwmVND7vJzBbFwuPy4nyN8gg1k0T/G0wjJ
uZZA9Ph0iEXihTBjl9iDocacjM6UkaJNCvhYuyOoDAbYI8bkKMsWzf74sDz2OSn/gkgg+lRYWKwc
YWcByxuN46dhtOri3ZYPAn5DlKJN6lTvujLcd1SlLPtVk/IZWkiwFySlWtC8jwB1wDvr43H9pyhk
zs701drDG0J9bW3I6XWuV6ZuW24Il8fFBsFtNbiJsN32yQC203XHWcSf8xcealgXCEupp+wqsaM8
xv5sPoKy9DZakInKDE8rAKjQaeudZ8dJBM0UWoo/o+RRPzvRctC5wpCVn38jAs6MHUEI1Uj4zrcq
Abe56owAlkyRuCTenmJe2HOk+UsQrb3BrFjEiCvwU9/3TQ8IIEVLAiDVA/VPoDfabarISYo7qRUk
LZwtlJogqz7nL52dxw17+Del/4Wk7eDekUPGh7CnqztJohDXclAuZcpifjrxd5auoll0hC8XYfMR
QDuu6EnE3qE4Rx3nva6q/5ilBhEAT5DjpYut3k5kXQmPcksvm4B6O23Y9/Sge0SN6b/A1AtbXN41
ylu3a0Ki/mLjUt3Y2Y6vOzPaNgN9qcxRFW1XQGD+qIPCqhu2NkkKBLpXq/XssnFCWXcHBGj0FE7V
oqH/6/EZoR2rgFFv0Rfw2w9iAcqmXgJ2Y3Sz21usHN5dyKTN0mNOyAlsqnh1SmNnj0kyn0FWRB8J
O6JwWWT1EJJcyeUZtqtpiv414XQvzhafu6cFak5L+qkWb5CxwAMcpZfSSxW7f8iSrHfYzCgI0ENr
sr2oZZUnKUdXiWxVEoNxoVtE2bgGfmqB8NldUr0L8sKv357UpNozHmjIXHJ0hz93SI9VwYq0vLJo
68YFt4aUuhahAseKRtdl1xIXjkS6VE2F3I5hC/GqZWBml+o7eSG7RJuNYgELPKVtJ/ARO+mK60QH
NwHB2r0ngsTDHW4d2mKcnkgS39k5BU7zatL+pvfq2XZkSkaJi1Q7AofQb9znBmMR3nu8Xq1UrLOj
DLQ0NJZGNPDYGaoTs+KkM3uBhlOg1Fld1tYTfDXscsSVVc/pLTfeYB8sdj2slsuRqHNby/0/ZkxH
FNV8HQnpLcw7vP1gW0jgF+ONgxVPqVl/FIpMM+EbpMcdsUvvnQaJU9VHvW+k51FN4R8TRwJx7/Uj
TnLk6Pr4XODOQ1SDH6xilkAFJxk+mAPHKroXq+pmdg0k+gTr0sO/+TaG63XPcm89RehNF/dy9cTo
AJEjxFoNk91Kqpsj0l00slPEhQcLKYxDzfLk1NNJ36EIS3ky+dna500zVgTzrCJ+Fwll3w/SIJ6T
KAZhRaeiwg23ekB2xjUj2h2ApD0viFFQT3XsJusb8IeYUDLziFRUv8t4yLRFSHR0o5IxA0oyO7H+
UZkCXJW5PERW/ZyNHsCQl7wgk7ruh1SfFfGL3ap0yuqErg8rDDehChgtzDe+XhDFZI5tw9nLHgky
L7KVikZge8Oaot866F7gixK5BVlZzaAFGKWe5DRCLvFF495lXGrD8EGJDSYAhu+KdNsewcXaL8tD
8p0F3UBcxGQ3JEPhFDmLUMgNQuG+C+oukozWImaeC8aLNx/Qwog0UoEK53pQi/EH24le1JepNiPt
Csr5rC1gHL+oBHtZcRf1sWVhk5Aa2NHqRtGiXjt4O9YbAjdr/keZcDYcI9YfxtQtzwJJj0GlzLOM
LbBzuVHtbSoid7Kr/lhGLtrN5A+CBROf0n4JnqbCxpJYR4Lt+NPm2ahNlfav4cKf5PwMtdCuNCNx
2eylhGxWjTBIlurmuegUNln2ZanTXil4CXGS6OTMJhloATX1ZSj/cnW/Hr/7rijq/Rz95kkPv7rY
9ITU8Cgt1fJizAPfGzf3GdQmw/Uk/ZuGCH+EvWqg5x5Mi/VkaCd6qOcIQLsuuUTyBeIHggHTx/cj
iGpLfVB11lzq0s28DENI2Vwx/tLgVLoH0Oi30oPqv3Lba0aZrRjnYfRQvXM4IOXS2CSe2ewL97ov
nJxQ4BrO6ufAkEWVVpiR8Ac6q5oL/imncO7+jMnzXBEMeH2odRAnEg7HYyzMk1abqC1RNAhAYGQu
1+6LTOsyLdUGUncda9cMLb3EFaXmnHDuRbN0P1Wa+fTKqk31Si5RWWFs6Ow5F+WVFYmV+Z11jtyH
0U5aJjbepBckd+zem2rwhaZ+wwYVaQvl3VUcsvuS9AMYv4ECNodUSRX1K10Bxo5WR2YNg+GIXZN7
g8rrM0Njd2ZeuuLhi0/xG+Kxb0cKZnzpQ3Dpd1o2W9TFu3l/15l2g06ooP6jkGsrNjnKCXOQ+wvA
KkBXLvT6tjb5DIMb8qFB/0k47MXKzIfLfF8VCVyhaQPMSFokZgPiaZafSIfs8roqh4/p6FWDOW4J
4w8w6dQJ4sNIOxRDVNY6X0fnYqV9HHsN1ki37ol9+FxJgzQXh7lmnILRo32RgVn2xuGmMz0bsGWf
lwNYDUYzKBg/EI11aw12CVg7ZVivXQqNkWnVLtO0B2lR2dNwP8QAnrQGaL6xa/syl7WooIlvLOVD
dwGcTf9i1+Tcnko9r2ZPJgJJ8zW9ekL/Mg5w95B/gK7zbWYD1uK3fI7bfO35ob+HVJZigeEr0vWW
DfpfIhoao8bDNTu4yRPVffb0AUG+/kC33hq4hKyBkoAv42tYwZ6twIFDpyW5AMcJpjEV1MNTlFiF
H9b5Lnr75Up1D6IQPboRyONuX9W7AQQyLYqaiy08iyDk7SnH1aOxkCPw6KdqgAGqGMJSJfLffWxe
QnS6aoWc9j860PIh83pN96N+t0MlTs4D4fO7nlE0SnWG4IwjfLRw1SoavTY/R00uer0lRJMwtnOo
9Edhtb9sALDveHQkxiyuBxuy6/7NPHoNa8NdCekdqyTOjdzwZ9CAtkpixoXFP2TMODlgOWEhLrbv
FsHLAxjTRjwFiA4q7T8EnT3PsQP7UdgPTvo6CeUYjHlTJM+6iAdKINYhpvnTRAvUusIvRH/WCZdr
xG2iHZgZG6LkO+DPjfJDtEbCE88OivEO6DBb48vLJKT3ImIF/NBuSLW49Iim/BBoeGVarTHDPwPZ
1aqXdISpW6cE/p8RPM15wT5VFM6PM2kWY6qxWTRNGzxls0SEuCiapphWFVGEr02yQ/wujJN29Shf
Q8WxgWXatQJbdwufUNJb3zgREu0hOQ5LlCcHeJgOQ3MZy+TFRVGRyr8Uv+YAxIPvuWirdsaSrs5+
+LSu5nquiV//igd2nS/k90UbZSbbGWOVx8tiOEgwmE1y/0KZYpi4c4iFb6Q9lbuU3j6B9usOaPpQ
IHgaxDD+nnUjWooo8Sog2paqOd7SufKb6iEhyrYeHtF3eZQ+hNHJC2xKFXcpAz5ts8thwOEudyHP
i9QHYmq2U6LvUH3lcTB3X7PMpFYwjBXyG2CiCdHL9b5G19t+GU9sOergiBNbpXAxkulckP8xRwlf
fwySBb0xHT7gmolqyOQ3FQRV2oqXgkXD4JLvRvXgJRJVDXQ/8jAF5KOURtogF136rgAX7bMSol6l
b0w3inj1YIm0v06v2Pg+Iiop6ozAzCCNI64i1XirUY5vho238nBeCv7l3WXhvgX9W/nHfdSL4aA5
7puUSZcTGlc/u6ZPj10vfqClId+Vgpjpqnuq4CYUaQTy/6bs+cnG848EFbIs51JzjzQBGK7ZJRRL
HPuSY78R9JzvucHAXNGZfkOcC301U4q6GgzOIvcWofIrxxoCXBDxPuJ4JHiPMKyDPwl7BjqiROYo
tyAqvs5KZtyJlgiwIBjBOnV5nvGYr9Rk/yd9rtXjU4EjfZIhdZa9w/5Sdasrwv7FqNG6bTGtRUuU
CTPt34Gvfrfl69DLuBKmZoK8OWXCEov35FqTduCT9a+/zBLl+fKZW+VMD4hvTHFhtVuVLvpKjpvx
0JO/zmlUuXiAbcyYOKMOdbDJSb0V4RzM1FLjViYI/SIu29RXWrv4Wf7zCfXxQ3UahbwT0CETTmzT
raJJYz3hJJ50kgUgLJRNdRPbKGaQ4BYAb+WssiWr0PLVPk0jKNBRPw2IEwcTnCVg/BiLtQSIqb8K
EDUwznEkdYzgtmf6JihoM0DMLU1NggcNLOESdEorvj2wrM03RFCBt/X7mFpxWbOPGVoVhkeuyCtD
P5Ml8J8xIm5hUh6uFhdBlBf+nQQQVuuhmVnmRoqICwmu+I1dmUQpxSb4mO/Ey87dagte7IvKOhd+
NLWMzP86D2slAayxGslWhf/tSBj8vskSOEYnnlEMNQOMEb1IldDCAdW2V9yyNSiWnVDBsur7Fy74
PDzUWH/z3zp0TwgiQdypc27O7BsI41k9knbJ9ibdJyuxCl7jzo1Xx4QEPi1bLkTxTR2hdQ6at1Ik
DlLljTMA7xAWA9T6o8QO/SjHz/50h29OTHlQxA5zoTgXuPHXyQiltsN/bZzbiPvmYB/GYiX0AHlu
DVeSOk+sGgocztR74wqXIXlsevzC8xC1OEhxKcdjunpRtTBw0vK8SKeVx/bzNlA2jgJDDME51HVS
isiAQlyb9FqI2Rx/bEhn5OjMW10x2ivanuV81vt6wQig6qZvKHSpjQfwoAFMK4a9nyjxrEqBv21F
LV/HuGJ3DSUZG43KnxXmxBLQ/+OkgHJ+xRCqXsvu9AGkh9G0cTeCJSmyu72+84PyP32XCiVjZj7L
pkIM1eC4deB8f1bgafKZ3oMGe3FzF3SOlp0eXxaArM6+92HYS9DIZgwgg4yOHhK+wfa4a3idUQwi
cb/1OtGI0ful7O0s8szmYHQojk4OoVe5m3qjpneBxy2m8NRZhZ+pCsyPnXDcFGT82q6nQmC7ySD/
hoBFTN2SK4UB+jTxZ9SLvGR/owK4qk0FCmvu9be4Qjjc9v2btLz5liREOSysVscMs3ZthFoacvAu
3pfzTbh8XS3aaunYM6JK0iUe76b1vmnrOOAvMdSIBB+Hg+iarH6P2+VENlZXC9OFAckNoeydJD5z
2J4c7+ZjhNdFANLrUxu4HggKtk0RPgp5tStg+T0erOnG2u5Z+edDis7P5EavuN/TbI/aRXU+nSeX
89+N2sojZCB55IobVkmS1KJDjm9y4i44ROVO6tDeVSvQk3JMF/ZVd6tm/f/XMA8jh/KaLduW9cEo
HsKDiF9gwg+f8kRu+5wn6pyTRxIOJgaMjptsnB1WID/VFKYgtQe36qhUhIzYXUk7dWBRcOnfLU8c
RneF2vrQn+QVETL5Q47eybaBBtG+F/uxzCRDaekih+76kAx6fRpaLLKZwUvBHat2/GMeeuMOFUCo
P8hQguVC7ROMNBmehLK5DrbU0vUWYMob7n72Lz5qUDRqfSqDNpTQ8wLB+UYLB0lpU77/ggxJBSOD
w00pUridQobTs9Qc3ytjksDBGrNrICVIq2HGC2rwvLuVbLvnZWerBS6SCytZp3hlLS7dDfBs6Wb4
Gt/DAiFriYhimrOUbDl6hHa/kdAPkDPFfvSKa7WWnT3mtTqbTyoVgRi9QXbaR12XhEljpjB9avnE
ksJnJKga+D/AS+3CMbIilpZ0lZRTSgoZOhwBIC+G77p4BLeEl8lNy+rZs/NJHMkmW53NZvQs/dxW
feSPhN0E0TPV5c+PNOaCdXEz0aU8dyzvdo7/UcW/hWb/F43WnOJssVF/qspup9MDAtdhAlFs0o60
sVquIsos8WK8GUPAMojT+dI+88QOUDwJqA3RZIfqihdGs/kb5o+lA5ZfcnSkluckTDBVYJor0GOr
dR4I1D4u0ppS0qkfdubeftK77pSb6di20JPBHfH/ChwMg067QOLNCTePX0ADGakA/deK1pZ5S2F+
x73zzmHvFC8E5xDFN6siUp7pV4D7nIGhZtHuRmoBa6Zn0+WUjVSVA43xns/7Z+93ieEXT4d4gVe3
XDo+EZFPjKQIIc7GcptzklGzqQeBQW/IRJFOJa+9FkNaKeBPmtEz5xsx6NYZHWqUlOEM8LwqfZWb
PmFFreI9goqQ4CSGmGq2kEP32z5hiq2KT3xWhHNO7G3tiKuksFDveH3IbjGfHXP6sWV3Pl3gwVll
TTQmSgAEAFiR8N37wy7StXQycJevovWjVstE4JEyA5n3G1CHNcDPEJd4uJz7pYiieWjf4D1fYljj
x33qEnlj+/ZgCZXr5VSP3Yz/nIbVHpAYUhqoBMPavKIb3iPWhbG5g1jHkVMFd2YDoy4VCDpMSF+E
aq7SYQmQqROP2PCt2TROELTUgcpbPbAd8/O6EcfnzP+P8ARHHG/cV3z776T+xqg6uCylLmyUqKww
83M6QHvaOiqqbUy02p74pE5xBUf+/DhN+07q8hjivBC1+56PdNb4Qj9O3J8XQmHVTF/noSVc0O5u
feLQrWEHt144HWmY0oIwzWFfL/j4+VgreMHqsreVgd15xM7JwRZkNBPdMzouokjmoCwEfwJYb1iD
+AyQvSxF6RNzowGKp/3f3F47ReK0MZtuNdo8RVFO/OtcInEeG6d/H3DWNEgIfP1fpwV1bnIWyXlO
2dypKCrRGyql4iG4eWoP9hPwlMZUfJ1lqV8Yd5Flk+3YgjQXJ8CTibOsUfeBjneOyPyGC0A5sngB
N2FncJotFkyUVrMCB24JBusLYojeADkYvc9mio6MqHuij03xUAnS6vXfY5yTNr0FOe6dW1drpvAT
kPDdQoPLLugFYGcxrnT97IUTlFcCyIuWYxbnmLBo3HJ7JUrd16HUwX0jwGSbEU956LxrVu+NX78B
XczxVLKOaJcSW5YP0IE/fXzInb5A541An+RNEWa4jWKtRr3LHgePFdMbR9eNf5r3lYfDbFDdnMsY
apiaeO+XxXmXQbL+vVHU45q8+ZL+o7mwpLgGmqZFFGEkBD+ey5JfRAb7Dlmwh3hONr09OoUH8oJ7
i0KZzzdY6fYGBv1nfm7XdVsh2nOsDV4+EeGZX/TI2HIY+ykYQvgRdOn9i0rC2Xpf9gMknAlHLDMV
kanLKgJ13z9IHx+G+6qv9Rya26M+uDwPU6vph93Uqrx6yMaV0FgWrN/yyfLqW0vXD7t/x+bTKwP9
2leU6tbbb54onWY7QNefJItyPCwRjailwroBqlx65Tf2RYq17D2kqSBXbjqUfVn4oDkxu1TiCb55
QN4aKtikLtFSbvGA8nzvE4rGhV6aTuugMlssWooCgcmC2Dh/wNFN77et3a2clsF8lknk70tDwuVq
jAPRK361lWIAk3iQnirAEKE/5Nhn4Pkr36NzWAijT6d72CZhmarlQ3wpHFRmJFfEGQcVSsOJWBpn
LOPozE2pXhKqkUj33Euz8MWlwV9/vBpOeWGqbMgxC5ZGgNPl+HY5R6345jDp4w00KJ/I/VG2mOVY
+zx4hTXuhJRdBzt1dK3NxcSGGHw38GDFcHEpbAcQb/x2tLWdHUOLzdcyHHgu5ych+pMnSUTgX6IK
rnJkWXlcpCJlMM+gn1wkt4qZ1rYhSfb/fs527xcS7TPaiAZbKqJ5otxqs2DCA4msMbqmqp32Gebv
e9zBfOUJc9nxSBxQtg0yjMz8L1mP12o5Sjdz0xc/HZ+eRLy8WPNejxU35jhvQJ/DiePOkI3Sn+Cf
1S3RMKKUocRsdAwLNJ4sfD0fJ7x4jZLPSfGjryOrY0i8/7K8FYbxULOnERPzT7B4RRXpabbw/aJH
F5A7es2WGeVKvgon5GZ9w35jgsHvMPxIX3BkfyywqWziuJb6FPnsVCOcrE05lFvRkNGro3JIGuf9
9EoqtKl/9AX8gKO0ZdIaeVe46cjOXTIhXp7GgSSjG4fxhyrGR42QIECqc4qjvAJtdGjogDJJOM4O
24zlqmEeUhezyTbUP9TyAQ6+HRiKrz/KmguNu1A7AdFrkDU1yfZbi9RcA3/JyuE1gQCv0I83Tt/5
H3KayALMNlYiDVQ4ruv57VWMtLVwIxyaNbuiyBURcLL2YpE6oN6QdB9oO9PSUtKaTEHdLsIl8STu
qqtGrIVKpRj9d8RYQLXzql1J16LGSC0AWjQl2Dgz0EqAakA3pIW85dPe4p5+II5ZCgCc/ZTD9XkM
iFO4q9TOS60fB4dUGfeOaQ/u9F3vAmkTU19DXHhxx/arKBSLmO/ZZdrVG6bgDekRuTxCOnR2iIPh
J5pS1IxJjGWSvs6LaOf6cXCBotGF9UABRpFvBOMEngA+8ukt+ArvLEt4za8hLO/gG5PDleWplDLn
Ui2wSYexwbYBRdLitvqXYEWSciNXtzhcZC3nhAtHzHKMhbix9N59rnaHObzAVRBX0jcLbul99NM9
f5yNVWVc9wC4SLnDR6Sp1mUVfiY1nNluLPFOGD9mP7YqgbCB865wyKLR06Vqasw9AiYvJSqrT1r2
hnS0xEcNyxeLZWDVY7G4WekOxaMj/KVOpbPmKxQkpOk9MBjLDucmpBS4YmUI90unxz5+1Ye5X1g+
qjUIQiLYeghJ4q+eiQoVIcjFyllnOwcPaT7YDdp38R1uXopKd+PVMcq3Mb5en0OZZRQENeIb3gZy
X0Ku3S8NsVdPYn3YJ1zqJYe2f+5Fp6prQJ6u1+ROAed4SrHM9/uoZqmT70RLxhnQX0lF8mHDQhkP
a0TMbxUsu35XjU1xDou+TUGBQPlhKMSPy1U5GOGF5DWvQYk1p+z3SXWXDtmC8yhoJhA9UwwkMXWr
gJ4tB78INVWj4HKHngZ3yi0JPG/FR5pLHA/TGZEeUEMZtRf1BuLrncVeg6lzHttMrkC7zNbF2dRW
bNc0mUAF/EWZUp2b+rxu3jLp4rAm2LA1z4na+csR7Fm0wpm2myXoif/g7ivur2tprHBI1rs7eHWF
lLd/BZbabDm217X+7Tmd2pqcuRaoRLmQ2lxYV1h+5/KwJS2kMi63l6FglCnd1yryRy6F/cCl/rU2
dmaXMcu1n+JsZrJfeXEO0ZsQbXklCHvUarXRjW3PWM4q4oQmT/kAG3O3zRWhh/eMBc2jqDBRnAmv
uzgkachJmbQ0zdRFo8+GS0StqC0sGaHceRXGPOy9aoQ5aoMPy9+kmNP3ylSrP6BaX1yIrig5g/NW
Yj9mFUzopZSwVwH/+K4Iwe1UDSLdH36hPX0Fkx/dvzC6oqmnB1ZJXAY/0HhAKMzjNZgRF+CLnxCA
So/xjCMXxTsXGLNbJ5Cum974nnYQ7V0wKtvbKVdpGLt8FMH/KurQtRiwCpl3kZZYhR3JWppB2s7R
Tch1mOXuJizqPn/wJ/bp+bAJ8i4niIWLr/HaLrBBd8fMk29l2719nBQMuvqt7TAbZvOk9E+OLwk3
ivoXW5gUt8EBJR4svjpKweEy+4qX8dvo33H8dx8/yZXtGFrlgsc9yWjkNuy/hy0t1XN956s8Fv5p
W2p/atLe5cHxVp06qJbOx75uqEjCXygU1/mFWKx03ySEh70zsuzYar8qQHeTNAlNAVcrW7jwSyZ/
27C+R6BIYIOX37e+SlbT2Em67RNEgTrSlFy48Qtjf3k2UgHQKghF8FqePflkW6sir2AuW0LLkZPk
mDKENgIare3vI2Y7ZvUulfzLUgrRPv8xGZmgPon1W3QNUhLK02q8zN4R4SUQmygUR/v8fDC7uKOY
plPVHQ6Uj83YSToVLUGvtveJ8VlVTnbxrr/2p5tzCuU/rE7PyI9FSuUK4ChcBZgbpPhXCaALUNtm
njeCB0wkRBu/3OdyrCkSHzQ1xTqAEVM4P41/bb4d/wcLycKABseuc5pM6PQ/SPY75egiBW1NUDdA
4aeixeln7RoN2xIEo6QGm9zt20xePerWk6KMmV+H7lxqrz0A0EuFjR+JYkwxmAjhgEcStoH/Y7jG
OUSUlxFgvh8ZsWNzj9eeQtpyCq//cWQbyzRGvU2ZRRB5QOpd86t3Yz7JxFPQpFV5gKy0Z+6xyXVZ
+uN1mMA4JGR9frlBY1ffWR2b39KdNw9J93vxt6m0t413pVTPvvjQAMHusGoCGEzWOtChDx2N1JN1
BkQnx7XC3N9uS1w9BTF2ABCAsaj72qcFGAPrgifq+/mXztef68c3+RTBjiabQaQ2bsfK/fhSNYZC
Pvs04QO5VK/QFKaVmY0olTHaqwlUnALNNm6VLtV1Uvcq3LGsmzu9TcOX+DbWwGm5VgtjIcMEHUtG
WcnGsM5vLSWEoIJq8Yiw8T9IuRJ9n3XID2thTWYoUSKeD5zLhKza4jx+9xPW5F2CuXZJHRGcGR+z
fRHZzW2c/kSxWANLZSDBUZ7WsWmtbwTvzkQrX/FOVbcPqOLTLpPSkAktkRbx4C/hvqxcPCTTRSCJ
/IqX0j86gS81RIzpYTbzDTi38VM8iq21ZAzCvBgNA0xqkcnbBJXnhXcsIIq0+f9/x9S4phc9BtFc
RYGaywyXsakWMsXZoHBFbKFFtPJXsROh6VhGYexdhUMOZtXj8OnpWD/W0Qz/uUBDm+8AmCZzwwTK
d1z0maZE+Dkna316C24LPRLggDwI++45ECpyWfUfzu++QZnjvLqsRfgitLKv+k56/BHeBSoiqlcp
k9AnMmjAOdkkzwTbhs1K62mEhBwPOJKN11/dMhf4MdtxlRpiY+BUjlidFfpDw5/Zk3EamVDrlFqI
LlEUslFpzhx85pUYxzYtNl4NvltLLAWOh8tCllSqYHwxQjN27jSUQJZruCQvYmABLUb3PbhTKUNr
wf9N0OQ4bXBaolBZU6RNYSK70v+DCA+lb/Zo5QikGEc1sKd8eYIlfKZ0fZiYVXpcO4limmwOPEuo
IIm3/E/vK9gDHDs7dN+3mg8iewvmyOoeC4yJF1vZXcvgvjFIdKm1gHy4guCf4BvSqQ9dbwDNbETB
gjypL8qRbrDViQM9oO53rqg3RIK7UgZrHUFv4fac+nippOuu2clMNpjKYZsYNNyV+z+o6W9wnPwS
niUqdoaF7n7eFBz2aM2E8E0XVHsazFYZNMGal8ftHl5B6mXVDxy0jVENuIc61fczvGvAQW14OTZE
0PRhy5I47pL0CJf/lqwD1Up/zBQ4TfZ6V5XQ/tX7uOGNkVYq45ne36p9v4x/+4J/slnZb8iV903A
dlgu6LlI0tHZjdMctWKUubf3NM9NKDNSrOmE6nbA0fFxCrN5FTGQS+w2NYzbG41syouTw9SOX1Qy
EE7A3KizJnZlCgZZHcqm0UoNqOUBeUyGjhN1nMJzjHnZOYiYhfvh6eWTahmBhOo2mgNMAxeEDSHY
1sOuWdf85EVz0yvt6/DqeBg3D1LAAhZs7PtLCr+kxcBg77J+qn6dvm/jGy+weh7ldH7OUJglGIJN
E8hy1AFJMqNcOVakHvEi6zG7fqMWXPf4dz90+rgHKcYB+nogm8jtq2aDYqupUZCYFh2b8uJ2TfDV
FDbfb9iLV5nEywjPgjQpreh+Ic0km7ya9EIyYdzQdv7gXHdnrYuJZ4QeWG2C16V3eGhf7Dw/S+MC
lrz3t5MhoiRLDkxfhvltmO5UixGhqpikfIJ/6PlCt8Ho4navKk/B51lIUvO3HaxpLSDsb2dHTlgT
t2a0Q4lwqBRa54JKn7sL7a8TxSInxV7uRwTrOEsXurGMOceEsKnRzZ8nwPeRnGCaErzibmPRztoJ
iukGhG2z78ALCS3z1hQCsJ42RAvHa4Bph5L7h7NJmlbpsYnvr+9hqM2973jFTaM/HPEalf/6kQuz
pI7x2g4ubvTah0mbhzWN9ozHSKlP5/Crmy84xP/52Vrj14IpkaBsSvAUU+2XRs3i4E4+Lf41U5Hi
ZsIWcktc+//UD67Ew46KK/90K1Z3DtdNa9Vd1Qqx5riWnN050K42lKG/XMUizgOxxhOPrhS0zedS
j+rfBJJxRi8XcD+zp8tWo9ihEEQefz/VZccuif89sEAk3pGF0CTOpok7fHUJ3DuFQorODJGMWS+j
RssX05f+W6zMVKmqZM5CrrwgYsJOjrT4tzgNpuPOC1Avar3lNSOJnfsn3qElaKn785JTMl26hWr0
K0Npb3Gt+GlzrfH7lEMf5ggW57H9/7ULJaETwouzYmrhliMJrdLks1Fp3LUoAvPCxJmR2ITcHhS2
MdI9chpnK+CDWf5Ok68Wq7jDZVqxg4XKkAXy2DEsIWayNkjj5jvzTXxyi2DgIvzYJbAhHuINrwy7
lgbWFJiFFuFUXrITcR0K/0UwHdQyo2x3aBROB2Q6op0R2YRipq5AlCEGzQxIhF/XnV01nJKwCFt9
7bC9WHgoQGrxHRcEbk4WyfBc3JeG8aJcoDJthMs7Q8QTL59+LNJGbtIE7mZHXvkhdI7Pcizp+RC8
J/4EDsLifQZwIZTX6RWrGXVhOQ02DFniNBJZZOsHkTF3mC+hrG/koDdmW44qs6nrjKHAFi9q0OAg
MU/5EXC57YRhbyZh7m3DAHlp5ZFxu1GJBOLZuBW17n9DCfzE/SjxCA6YzGbgnEUqg8XejLlTviay
f32Qv5USoftogi1bFdXc9bloQYXoBgaa6KJmxX8qWERWJXUD3q4kvboiKqWj+nPQ2ErZOn7j+pTq
EpF4hHzFCGHJ5S+rFAgiciNcxb57zgdMtTJjTCsM2ModgtM67Ct/1st1lnRvH8KkYDhi5RTGpW0Y
RonSl/xFxPev0dMOf+CaZT3r6gIg5qAR2ph7PAW51fhMfwmPK2ewCv87rCY/dynQis101m57yPo+
hWOIutj+ELOCpJqK5kWZomVrnnE6rNB80C67TbBBbyxGWuOtllzvPrQLTZ1BZUQKjj3rKSkMIt8u
yvAsJkSGImsJUhRit7Qq2Q1oncP2r0Ev210nzUcB/SgrcVo8O46TmU3LfHKssxSO5Dj6Spxdn1xH
MbsaiFL0H4EMx1JU+NWehaHeKoC2f5dO+8gNjJyZZXmytAvb8ZrFCc+V7f7oVh2NMPp+AiPWQ20O
5ePClzqbrb3ulC3zmPjKAeBTgGAXYU+zFYLlzds4mD8HqfDmGewnwnEqQL6t01iihcuRPB3fQjn7
cv6ZGh5SXpfN+dip7ZCoQYq9SDcwMheZ8e+KkGQDXOs+Rqg/FfG4AIpjJKJD+6MtP927Fx6rk+lF
xh2PrkbgqeVsGrFHON/IBKyT7mafqlpzgFRCVSuX7y3dfBArHNZI+fNhQnfE46VpcMfhStmkvkx6
z7VJvOj4koqZ92Ud7O6uYXIjcIZtMk1cHxor8w+Q0ZVHMyO09hP15DGQr4th1nSygPtjvKx1j9Pk
9yR1gIwXSWaQj9osZ7MMCPc9zpCpacIX9WzjPG8hL7huUe0QEdOlA+1JrZ1TZdWM0hXfWOFKNK88
e35dquNeGrDl51MhjGjzsRxhUPvzjoDUyzFhGYD2pR1lXir8Fn7qt7oazW1hBwoi8Er78w4rGJ84
kC1oQ8LgGh0yXfZ8nC7CK++YO9EpYB4o6I6avcJnukb82oz2Np+x87cAjDBXTdLu5dGoSqCfFO6g
TZrsUw2vSisiujhNpPEUGaCiv7GbZ3QNMG+XFgN3tGu0J2/nsVonfTierJgp9bbsZbQ3gDLEipZ5
jgUuligPuFiqU6N7VlSkMoD25c7/A+wgTGTQ4jsGXlX1R4tNS8L1Jgk9KEXQqE5xk5NGlS4jR54h
xkfFSf9zWTbwxPMSKijqcWAhmdS/GdWK91lPY/u99TE6DFyJF9JF5eA3bxl63jDPy4QQYj5Jhcie
R3Cn2PJQi+OCdGs1teVaxm5zUWXnlXgP9ETWyfTvprb0Ry7Yd1xfyZR7lJI19hgm1892NhUzvht3
Mt+6jq1KiHWahWl+IKd8u5FgAs6FtMWdApxKiNskZo6vxCPbApAbKsm/vHlW0WnhYSMi5H2wt0+L
vj3R7zPJ6kF3AYpilUYO82jHvzZWemkyD/xMYH5g/wwbRNhGFMhBWNFEB/w2/bTakx/ze3J9imOQ
YywBbzmoFLet4u+bxUqibnqtlWxsNp30N7NO1n0nKnJyO+/m769WQt4EiCrHDn1YjzOHsb1m6VsE
yMfoJe8FZ80xVLAydoO/727GpA5qveSsYnVB2ofl8U5qBHUQ8c+AtgvMcOBzuOtgwqwC0ziRsNRo
rFd1++8N6aWnCqe5EAKf3SUf6jDLBDXTcOhkHKxBAlXaplkS3mgk3OMsRKtM/yHbIdvjKj5/Biq2
ZjYcy/rh/lYfA41AeoN19Ukf3z77mSwdtj0vMoFHbidhAc6o4ToOLEhG1RPOl9MMHqxZTTX/HAOG
Q19IXuDgqBvk7GfOKcjV26RUFABhs1zb9K6ktPRbXwibgFxDQEcYd5kRwFO23/XUgl93Bidebfq0
ZjOVkF2cQSVlW5bRQk4NU9yZCXGrPyfg+iUOmTrA2iWRcPJ8pTQCzTBVz92GMItvofM79nxbsPUS
tAIv0s8SFQbjPkqH6GizlLKoqlC1GsWJy6zUL45P9J3McRHnHCKlrSL4A+rLeVlim+wmX8VImVbE
KxWsLcWooDwTmjJTuH2NS68mIE2gLeK5ovKbZmMFt2LqKb5i4tU+CY4RXDPdZnZsasU0KN9CvwL1
OUhktZZsTKaqyEu//4WSutlmaquTyCs4yDv+regHKVZLUk4WvP8fOscHNHy73AxnWSepRq7/rAUB
9QuGxCkjRxnf41DSrWcESZZqAXlzzBAmrJULJ6IXo10EtU2LBOxKlraor0wRxksV2xgDhAslBCG5
6vmwd1Uy00KiXZwGNPWxp90fbrOHU5ynNiqqTjMyVBq+yYP5fW8uQvl0pkMacKmvNetOtBJJ1Gj8
a6MRCDvq+WBMMPwNKQnLqng8t8zegDtudJvc9FawqmZ3F2Br3yb1F7R0f+eSavyyFWHI+DDzV0qF
wm0x5d69AQjfBMHaf6CjdSbiJROyCZ597/PxvPwAYUvf4eW9EnaQaVhZUq+qDnsextyIdPwyfvoV
dkkpY5SUuq5VRYQnsWkLT4xlo5oHcr1ty4qKH46Vl2BHvUPWw67qDKUbgxmnz3tAra91CsIWT/SU
jjAePLBHDy9xWowku8XiMcni7s6Dw3asNn7D1jHjBbU0wnfRG0J3nGgBovtXzygwcWm1Xwn/XF7c
AZsGGbF4CPpnUE7mwpyk4r6kyV7049YQt8TrNBasKdT1HzJ9uEpUv16WBdOG/DMpEYtfaIRZ5Lp4
GZYrmYjSGShsc9x4j+dlqgrZWbO77wvjRVD11lxjjjD7xr9qLgXoinYacz5aTYF9DaIeZs+JYpAr
cMAYoVVmbQEomzRiQO3+KSwYg/fdm1kGUBcNYfhFadz379EhhG0Vyk44m6vbQbHaIt1q1p7nAf/j
POt6iPjgHBDe8DcdyVFG+Gz4Y3R0X/ix2pkh5kmmAt6XqWXgK42i8GBc6cIl8J1FwFON7WiWC4Ne
PQY7s/Ud8eCezkhOo3prKry0RydJCcvsaXnnGHG/iIEuxIcs30CylALrnj+110mWFAJAvfPZC7ou
LFJQJx9nFQcbEaEhvXL/bx4YskoVb3M7I4yG3v+sDp+61ADO51sZOA/SWZNTAtrNI/3fkP3FyCy3
lPaYsCVhq5G6K8QJytjDhQ3nsLk3X2aa9PxjkSkypNsi5XYB1Ayq2qfQxnrtt4M2sd6X3gpLLmSF
h7iyrMiF76L7sbjQ1wRQjpbnUW5VgQBBt2GbWd1xhCL1lnA2c5MWFtGdq0/xLtNivqys7izBuM4Z
f7wZm0kXg9/h3xfEfH7cmuCM1NMWkQFbzUpCtoeC5KOCsCtbBzYnbI1EwoBPRvmYqV+JUbCm8jtO
uVBfQ1Ir4U13tU+XTbU3hmwdWv3NB9D8cCwmgiolv7yS2cEFHINqRf4jfeCwEUWTsS1JUP4S4Nte
9Vuukf3KDWtwA4iggl8EEGVeWp+REiFVFaE336nw6tQjIbBlYhY8IiftHW/DpLDfdeE0bDp6IvNK
/xM71afMqGgrGY5itVpyPvYfinOurfTMGvJGk/hbg2d+89euKZ+FpLrf5IxIXcEMIISnDVf1/ydw
i+O6qY6JYlwH9110iDbL4f/4lzmBGCGDiFFuFXhWTPSvO/kPdd8F/lPaIkdc8PGk29z6CBcrvOp+
sfvnSa26/hASwr8ZeJH1MpZHJPMrlBcJDyHLFsRfHJL+C/SCT7TG/+FRtR95QPHKfwMo3ArKCxoc
PyvEfWIRsTHlSd+f581EID+vKTWwbF6Z8PnCwRvEFrgaiyWylvIm9dtIh5DYOdXriCjq9cYryyI0
l7Euo+cbYj9dQlTYAGgdZ3i0OUzkiDwnnS3pA8jMaYB2/rCOqc82DPfRXI3QG+WfA8nMH2iFbNzj
T/peo+titlfgKrHO8Vah+agaA9D7qjiXfK48p2hVy7d5QelyYo4LEg2pn3YeB9Nnrr8vyVzfkH+c
kyOE3PqCn3KJ7vL2BbdKlcVvsOfqzZjeFED0DgO+z0O+YSSt61zwWNHVfXQMpmUcTZ02k4MB0hZI
1x6KXTsV1IzCmh+/PA68R7i15VuBVqTQej6ED4uNvhEvZVIiSTd7t4cjo6OtcQgM1tpWLx8EprQZ
WC+zQ6E+4NxgVArgYYXcwprNWtru9As4qiKQbD0qllirV/yXFmNDmda9/I++L7N59THmr91LAu0Y
6eSeG96wwkHVdFseeneW2aZNPmP1C1RrqxWNHyv5B9iIRoAK5WbRJynKzuFalO0/5tXJIIc0SfYi
txZkPULbsL+WAmjtV6XfgaAfI2A+oAdAFsg6GTu4+FhY1qn9j1IqV1MOUmgpP/Lqyfx7EPA0EDa7
C0EOldqq9xFh0Ir9odfoNZQVV62pLg695IWNRLvRYJLELUe9NoOqrhZWEs6bPapft8lBK0rq1Vms
sZfUQO8viMof4UNuUK0iutG2once/b98Xd1J7uif78/gZaRvvRmbxIiDbbuke+aKmUR+xINCNeh8
QiDS5K3xKVlFSfeBGLu9erEll7FzB1QqLYpB2q9Rshcg+C3LehZnC993wtum6Fwg86DDBE27thcA
ITMV2EwKo+hznOptsz/9S0pVDvz8qC5Qd/Ff5ugOQhrXOJfKhz3gy61JNbdDnN9owV/kOTl9pMqv
XDWRDI067HRFDglMm34CpjQD0E7VpYlBtine7DuOMK0OTxpT6gIBK3Eu0cIytvlPIsQL82Gp5d/N
4hDY8noq0a8PqLOB72R9lf4vnvewjT5+vLYCtPjur6pyr++SspYMMQ2GN2EefacAhg9hy7Lrv6dX
ZSDWaxcR/WoBQNefexNpy8ih+A4wAqYOEuWRQxujhgasAuI4IhiuaiaSMPMRUdf0pDAk8pMFEoCX
MWBUpmisZCpke09a5nEkc8DR+jLFAxRsGEHzu/Lf+b6D4ax5odtMsHAiyUTro9RPhTXBTaM8bwjw
GgKHmLvJQURpQhU1E/Iu3Retkif3q1/Jy8NyZAe0VaKYtqb+QvqTxonziEDWHBaRItRWawQiX5SC
7f7yzci2YKIALYHJ+KGdZgfAj49GhUBANXSt7ImFTGmG9iBuNLRWQUONDZC62Rx6e64dxDE9IERH
0HEnhzbhsXv6fFwPf1/iGXEJwjishwJ1Gf27A0J6dP/kx2gy3zko7fDVpKRSENtdESJjfG/raxBx
zHccQj68j4u/xCX+axFVWUuAgPMyxcZlLy6pk5H+38LrsRhWKPVxvzuUmB/ZEMyZJlXtsVh52aIK
tr4LPk8yqmrLpJ0n2BLvx/93+RGvD6xkkOkKJrAfBtE+ipvFSsJn5zUfedCt0/kZOK4Qple3hfIE
FGBET9kNBptm2Ng8dyIHF8bte76tjkyH6VFTXL66nicHGJkfdui+viWrvbpfpQ8KWZmxX2LxfCBm
pACb7Kc9igMksauXEQmaHgjGHCc9I86mNLsPlE98FU+3oxki5gM9JOBLF6hg/kV4Zc41OjW986uZ
1y1fT9rWZSgy1VdzClVoG9nXwfJ/GufVLCoTk/GMguUuS3QeyS+G2aYO6S9iIAC/kF4y7mBwzmxG
vl3iOz+9VdCa2K7y6U2M3yNasmySQegi4D8UngyREE6MYkFqFH0pLZZrqZFqshsSTUwvUMKkOJV7
c3jHdFAJO0x9WY83rCFxLP4XRUtnHRLr+MP3i/YyUxMdDUCZd1zkJlyA4CzZ7rHh8Lo86kF9KbD8
G6iME6NL0OpiEDehT4OcFGoOquwAOTlGrFKj+tVSuyUh/cdd7PB9ExVaKR1AfceSWrh23zdAcDZw
WgX0RYUeoi8w84ldppI4h26TXDXcHcHEWnjl6r570wG93PkRLO3F7FucgAWEX9ecKEYgwWfIq+MY
tcZM+k4XdYsN5j3XXxtcGIuAbr+vBgMIJ4dF1NawEXr5uXOKU9jMS8MNu/dhB1YwrR2Pl/x87WdQ
jWVYSbXExaTEGjWMV2E+/BTIBpwRhZ/ww2J6KlV9LXJMEI82QLPECQTpO+bO0lXDJ2AZoRIpcdew
LBJAtvLGGnb84nlJ/SDi3Rh8u0yZ/Ro7jQWcVJi/q0QamhCDJd0WpENG6ElVFok8pzOkP2nnedv+
gbnjOWxca29RaBPGLqy90WyrkDmdXnp8k24mXC+fAi4JoKwloj5bMCXVCEocruDcEMLctHbEsQls
Pvg42ceMJZVKvw1+EJHVsaZ5t/ydtyaJS3GAWvW2ByVvFki4U51vnwrDvPxLQT2aPdlM5TIKyhB0
oP70SbIVGwoanRxxMpiSh1EKYo/jG7Dkt6F/rfqgGYwKykZ4J4TLz78D/zsqReMWBPD37joL3QU8
jeFiKxMpJNMZ3VzBfNylmGvfi6YaaG7auvOT52cgo1Mc/HaedfVtqjwg1DSLGW+Dci5S1rSAxopA
fG+7QQ4I8Wcx2JCcWU1pTMBMfQKIVO1Vo6rTzpXjp4u2UrCPStOpXzkhnx5+jSFRVBH4CyqKcKXC
n//cwU0CKdXogZ5KdePHBMTpq2MZqeDt9++bObd7Wx/UbnYz07mv+LIaepB4U3iMueXuLBzlQDWg
/I/VnPWrZRIQ3dbfFGJVi8pumxED2UdfS8t7oAgGh6iJrR9XIavvopxlCYnFYy5GMxa0lbaFlo9X
XKRPk+fFdy398lMG0/8QoviNkGJ0dWWsygDwQbQwfUdSxCJVWmiFJkFkZFqo+elwc5XDBYuAKDp1
WyJKN2fHtG8irxDvT9rFWqLsGFKhV9GEwaiP8JQZBEuc9R9Pq+f98svwoEo0qGvGomCRXZduF/zr
/291qBUrSDbqbduoA3QF4Hqiq7pwKQSp34ECw6KNn71wpAG2ucVzRBgCtirkbwBO6bXoalWZjy1J
3jczy87kuY7yMuklDZ2JbiA+v8EHLRqWgRYPem8ChmhSuRrJXVpki/DR/p3JjmGpUChA54NLu15B
QpY3f3I4xYLf619XGU7VCCvK3UD+R8p0pywuHcl2X6uidDmaSoKsDd2n54ayT11V3eYg+FJZqiuO
JNsX4WoeGSm7HgGvCnzPUi8V3hn2H5QziEnS8alxEjuCyxOnBpHPvLNGZAKgNpnbbR8e911ajnPP
ELEWoHk9cPdyxTqjPAOa6IvuLs6cRM/hb749XP/ucWy5eocQAurQV2kHss5VGtAw9tFFtnMjy/W2
L3BS0eA4qHMb1x9Gpp0e7S1KCo12YvPPvTBLpKRGENWDLb27aYxfBvAFfNUh63ZELSKAg5j07FM2
A+NJ7wh+mbWyGcBAkUz62KlYOqYWI8MfhWRxGNLy6uOdkORwmOdffzXFe9Xf38v3jEN6QVwFPohi
aOUJdwTNa3Mw2rp5bXTSNjDwGnknvMW4JvRZ56gjd1z8Tpeg14MgZL47/eTrzSt/H94kn33hZVYd
2Kljp5BKAL4venLoW7NcI3GdGaKMSq5kGnLFGCv6JF4mT09Rq73h8JJNiwe00mvV5ivhq7Jixzl9
kqxHFJzYsCK9pRrPdzOJ/woJZety27j2Kj6yZGE3+ajXMrE4QtQeIvBiSG+daQ9f7xuiuu87UASe
ngQfxYmsxsV7Wm44uEWDJWQleTi8DEYOzHPL7UBPoi+Txhs52RT2KKfWxNxqRL6hWVL3DwU9SA4i
nrwhszaVrh7WM0oX7DuLVlWVx8U61EkGpWdCn0mef6xKnWT8YWCMaGGhlOW4bbp/9A1gyJEhQwPo
s6guwlrmZk4WY4UOQvQ9zQpnwKk+jDHrXgj2VNEbLxJwiVxHUpW+depbCr+cYQYQfIKOhKqIsxcr
mMOWGsZR5alIM5IGk/+8eWgtEhLcFNh1jAzlMK6yQZYrpcGKBa+6xa9acSQ9P+T0B8SHKx+0BpHp
QKzNtOzXc1UllSi7pfUPuUGpjKYVPzMzAEnJceo26IuzZjXwSHERzyEZx1jKltLZHp4ykY7hISZc
SKmBe7qVE1I/omMDKa44Uae5ZTmem0R8u0trEtBQ0ic+MVpe9Oml9mYIi1u/Lg+atSjX7QERIvls
2LufCuStzFY+8jOIX2MzfTR8gG0cOlMFhy/ZCRaQ0g+ESMEijcWrn0ozhyc28OQxikyGzN3kF/HG
aNDmeOsGL8pTm1SO4oBPOlH2h8pEHEQrAJo25xlnYOjSAmCLLdf3CsBH/Be7V6QmUpfHXDfZUdeG
FUqjBLAY27YUlPEpw5rg0kFRUjItrMDvpTVsphH9qgiGIMY5nTMpIcay48zQUXz72JdL93JymTyn
3x/qzSqWX2vDt0NBZewttMZRMMvqq2NWzP+xQrcyry5gyyIwpYQ8LmZhb/wwIzDHw70PiWDSw7P2
4Qsr332fAJwU8cB3DCxJVmH29yzGOq3K/MDQFkrCLS2sYBFf7PwMaAMPNdNYQpvaoj7qRzmExWRp
TwrtR/4wu9OUAQWk9vHb6BAeXsBn89jJGdEJpV68o9ifabFSra0JyAsL90fFFkY29PWF86hs9NOv
mfGDgP9P23I+Vajgyq2ocRkrbZIvfi8j/V44kxyIt8ln75JfIS4fiLF0DsKoF9K0fjLMTxXMrrJj
O/y7hdDw5MQyhyWfSJ3vQfDrKEJWgKF0XS2BX5OBPnSXvDjGXS4wJVRn4o4DjpHwemaf+89eH7+r
NPPw/m6DLX0ob4h7/QZLrEszcOrrK+M6v2RW9AdJpKCX0xDujZ7RMtGNREqWEKrio/kuOvTfS3cC
rAA0atzULRe6oMTY3TTect+RiIviqpuTSDMrrT1jrDporvprOq/3N9dyT1vo5YidSwQ7BYlNmY6y
9/1vgPvHagnDrPDh2+MURNkY8xhqwm1WlYZ3++5VS9Y6jzlVZJxZbYeGzWj1EFgVwuNCY3egJV90
zgU4ty37Y4l9Da0cZRz8ZBU3dfTr/O4dm0B89QcbSrioinnpEuHaOSI9EqTY/14JYmBH5hiqGh5k
DoGci0vi9Kz9W6Y9DsfpJscTaVQMMy87rUyoppM6s/4EZDPRpLfMXW+5yaMCKHrZK/nfufs1HAx/
Pv5EG2xRLTlhNvcFhOXPWKl6uLiI8NtHNce9mB3khbZm8nxiN71P1Fe4E4+KZjjK/eixRa5hqT/r
7DUhvGtxmTYl8V7d3Fi6QqZvhrPqU4w3wNSD1yI44PTFX3mqZkTnAaVfQhuDcBBTWor+N1JODG3H
HUz9XCA9Wk50dFl4jP3/hJC4PFYilsvVb+s7CxrlpF0L0BF8cENOGELAEllfiGRazIpHDF1QnYEt
X+qU5fMend6WyPG2axLa3cCjZMnKhJehPk/EgDS8RqgNguwfkqDMOad2ZzM3ov4yOm/GA5EXqqjI
aghSN4HtCJe2SW27JaY8SGuo9Kr9/xxR1lO4w4dP6QnkxNy+/pIYLNgNwSCKFJfUzF9on5aOSn4V
y0xqPqKdkPJGOXVkqYyE8KJ65cN+e+ha3hssHbymkPKODivBGCigbQrm3RJlacCsFjKzlKlRek9Y
gO/pbFevdoQ0CdTzjmt9WpNe7TJSC6ymgJpWfBflwrhrWTbHC7dye9Zgj71tDx8x28VXvM5WIP+R
ZunGNyE6mFMieo4kJNnhM6uy+XYhhlyXA9UExKLgwMvGGvGH41qbHaCWmav2V85xi9gUQAGdC8n7
rXvr+Y5SZp93QiHkplSN+DKGQnH7GvE8W45D4aIbCvLLpgbgbaBwYeCZKo30AxhuzAaEwA+rU8pz
01rVYf8Px5Trw8rRORdRY7K4pyoEvDZzohkqD/UCzd4tkmkTPuQX3QQnuMSTZO2RahW3M7YfuWhO
SHQThTKaGjMngYEGwiFxCJopVy1aiQ5jwf4XxSceeoPatshcMLtVxL0wkchS/q81j9wyKFy8odSs
qovoWvwaVt9tKQUOk26OYfNv40yM9lRwwKeIEcnCMJsuOsllZzkFTKRywzbpwSyBgPurdHlH/tpw
vxqSFgJUxkOkPLOwHN9Oy2ax6FaNpxDDZB1TVu0wqcanIgHEeH+3j6w8n7FfYoXYcqsVH5z9e/Rv
q8IRqjJe8nh2m/kBUlbqOD8UnK/9lJuuVe9gi7dHccxqi66SZKlsZvBhtA/t0boeMFnRScf+xXwf
UNRlSossROn5n6Ie7nuFc752I6DWS2/mOO66gOy4JwgXlZVCG7xQo7IsvxM4BMqPxrNsjYf//ckJ
+k338OceWZ4xhic1Ey8ZyI/o857VSELG3FZFxc5GKDO5EMeU+iJexqf+wK3wXLDpkkaOaFIjKQY7
fkt8ZhkguBDty7oQ8kqfobRSNA9Q9krVUgf0+odX1w7iKSwQtHl0FkrYKJrrGzQyG58VFaBugeDd
V0o36tG8+ChMt45fB8IH8q/Qp45ILTug6xRfnoSvB0F7rj/hFkPjBJSPK65Q1gllSKIbX/fwbw4A
zWx/qsYAr+Ytfj76nEzb+YaFq5Zrasr8mvMLi13W7q4d6ewC3FtvIFiFCaPPq2Q9hEOLkjyOz38f
AZ4S+6yX8yDfGRe2yQEo/XboGz8XiImUvCQNe9S6QqCAhv+/SKGQRAoAWvfyP28RDt63D3QvKaIm
OKvgRSRNmPOzDtzf1I0tSh/fG8MGKX7fwsgWgrH+VGLYCLq1LSz9bEDleRGWpY/iP0gK3FbbCvm9
2qkxSMuU1hY04Hzgd4nxdB1f4h7FM9pK+PdGsDfFHl/xhT0tCe/ZfphDVpWvneXz+OiSsrxmWLYs
GDYz9Zw9URBuCaw63oc++jeQmgMEh8EvimiFS/3q4e8Eukn3Ik2Iwd+RPCjw54nelwxevLi18zBm
ojcJ92VoXnuTIJOohuGYkRYm8n8txbZ4pAgkpaUzfaQGUUamqQrmHaXDq7E0fwZ4mH7dLpSXx5Dh
mP9okQczJzaJdh1RGGkfoztEFp7AFdZpVNVriEc/lpZCkUe2ljRCWx7aEhD/+mq6r6yR3fZF88fG
JjPGK+0I0yIeLc20xLKgy4LL6L5FzcBuW+x1hVS4JW7p/U4GaOBMcQLvE8zAgvLwNe+PArqBClb7
B5fLEB+nKFRfgT65eIRJLIZTXgpqnIgHU2pLhnXjfs6GETxdzPy3fv+GfPsPQDAfFjHRC5fHkVOZ
MWim4unvJSkREgdBdzE8V9k6II2fLcC7xrTcsvZ9v+rWxSWTgm4HhReAYywIioD2awyOw6goOjx8
vbHIy1TAO+Dv7Cs7H49o/xDpr9lFbH37zu4MVLL2HRLr70COwDZ/UTX/vXYlQmhYqx10iTcOumn9
1AaNL4WYLhO5QU7zKHtkDsHTlS5qikCOI2cCaIWhKXHNyYTU+cuBfksFW4glN/3xc22qccaKP+Vo
DHftfTS7tDzS7ivFtz7QyQyajf3BhIK/+PPBD9Lum7BzmFKyorwWZKYHY5kFj/tyoyJuzC93bWwT
mJLzGfTYEN3ktQr8GmCOSzuYwzHOSlhv3ekFZX2d6ZAvmUpKg6s1CM6rpo9IhTvYJn2D2TiJH9Og
9d47ks+Jc5AnxZCiRm5WCcrV5XwCqr+nGVabo/p+dLKsJrhvXNowaNupnm/oF73mPJz/YeKjTqbN
SKNvaAyUDtWB5mjKd2pylh6XCq0Zho+ZKlHZSDFR56piYlLrocNwxVa1NaAD/pj4hFCH/yPAEm2U
+5UTx1xym8O2ca+4k/Qr69zwoV8ljuMEePqtsycg3nhgDw8Dds4EbgNWnKtp3Xh9Bdog757jal7l
2F6Aq/KF81e1VU1qHUC2FCqtJPXtlYLKBzeXD3BmuLcg5/to5fqOo6n6bI8PDti1WZVSCHBdLEZn
4HTrvmSkkYKTIpHHUahXK+7PTdbSbByg+0IDC9heYCknBY8SDnYOIo96J/zG5EqOe3HDMMoH3Ne2
9thwDmkeYdhQYJothOprGwhGabwIO6Kx59mxsGrMJXldBHdSRwx1/NamYgsJRLd+gfK26fZQPyrg
Ti8zhoNAv35MAvhe8Gu7k+3MOzU4wlx4JIra3jzLO3LVs7fMiiX25y6s3PQN+JabK2iKQ7nW23Xl
ElmP48a1dGFOEspB8S3eO5ikv9xVY5zVnI4mv5XVwrirzhhwUG2FcU8meYNqottrQvCiK1TX7Lxl
L7b8LRp321X5UR2s5+uHvxbAzQOfiO4gWdTjK4BiNUnHbtaA+uSlVwLnkEVSMs8iQugSBJCJ7cUq
/lKyI2WujNJCUj++qcTyai/KT3Ut6fyKDqaKy4ACT7W84SyVLvKGHy9bdYXKz8tHAYxsHhMwe4hR
vi55gc/kB8qxwU5Ry20K5brpm/wLhs6OrdchPx24Esxsaf3DWZEcwQ4q+bZsz8zSYj0YKJKvYf5g
tkiQvn5SIuSYzTwFKrhkezljdfcATK8z2hh+iz4mSUzNFXOlZ8U18rROdVDZR5ArgQZBDj+qy4lZ
xcVR9ihkPFDwEoEFf1Mu7I4HDTO+u9Ce+BfgDcGSgAzkTOqMfEiA51W3cPs7iv9s0IeSleWJcb9m
qv/MQ8Ej3YsqYH1G6MYErhlm0mxtAsWW78JFh8+WINxlqeqrb8FJ3kabimeeOXU89Qp2DLEKfQWJ
d9SaciREimU5cIAq8AXpoPplb95yur0dQYzPD6DgCsikuytF7/+QZTRVA/3i3W9ruLjKq3Ek5TiG
i6zXkdQ8qYUOngGZS2tkLWiH+xEy5hMO2gLqk5ZIHNz1z3KvzwfRWfFMzvmsGtDVQSJI27yRT9ha
ZQ+1g0+YRj6SNkMc3s7hNYNsuI2yMa467qRITE+qL51VvVXFP0XZJ7X9jS2Ts/6BA7tDtspA2CqV
i4tGkoq7vW/Kw63cBKxlYfwpCG/i/sJ7SAQFZ0RtWT4TmNuU6FttreIDm1EOvTYv55e+CpsIghBp
PF5VkuLM1KhMnV1b5gOnEfS8N7s8Cm/X1FMoeQW3SknSDcwnrNZyRAIRSymhedY7VEawkwHEIkFd
Y+bXkchFDRRPhbO4kyNlBsEk9J87DFuxfZUtxZ+P+fkd7st4kNHIsNnomyFkcfboiWRvRR+GPNu4
BD+dkYi2uVz/8/XuuB5wVLh82R+dTT1pUmhtBqM7sXW/jXQh7ojqdv5KIh+eCw04wm2uxpe/FSzG
+3tbbRJT3HuQ/fiIFAOfbFI+SsHjW37+6khDU/GHKj5QdIql5w+w85eJH1JtlE/vmtOEINX9/c1p
qYYpZpyGsYbEZgzh9ojmqAeCw3/0em6v8YrKZUzwSO5UGaseQ13mxInKEOIqJzm7It7zJtdr7sDI
todiqiehqjNkgQ6E2mH2w6mkO6p4CfFSyADbVo3OwhqLWvsccahR7f6OzT8D25b1180c0t+fxSQ5
49Xk/Ha7sn54GOde5QWfa458Z2L+JYEbRl4lkCxDVefm98SmPJsQFlxrF2Nf3klAI6P9CbYA6b/o
BYBe7nAzaR+V4z1V51RYll1MruRHyXjja7IDxCqGpgZdC9ZgOeB4He4OxkcCSqEuVoUTV85xH2Bs
AawGojkxpPGOvIO1RN7o4+cxF2Z6cq227u2GTFj/EwqTzDn3JQH1WxIaCEQBmjZXxHT5IiiQZTEL
wI59YZlfr5G0b9dI2Mu3BK9WjdyXspAVj5sVhuu9c3qc+ZUmdAPaAcGN5amJJ7v0BmWBrjn6U8j1
9fSQBqiA9LzQhxswtkLUmOvcx4fjRDIXZ/zweTpV5QcsqgbKjT93pRUN/p/Dnsz/1WbZWfqSzU6U
BT+Ds0YU0KMLAlxl7TblCf8YZxoqMjfEegAV1JzK8WVEAVpzO9dLTe5m0nhkpw8Pl8MS9oVw9aGW
2E+dHZFN6GUE++G1ayRxZWuGyPTvh1iqjEf931VARoJwXIVio0YnJHhE8ogb18PdncJVb0WYdNl3
10tteBqm/wg2zNNg7EKWNw7H/3ZK4/D5O4zrjdzinBiDiTLQ3DFIVZkvGHC7/PVHlWPm0hAmzcSq
VowbTuIriiSAZs9RTXVS2Jou8+2gexe4/68WW4N2QI4XU5k8yvqKyFL9Tkc1e0GxWoOma0kuvl7P
i8BZjP+u+n3GPRAKUa2MrFrEVKrX++XyWIT6aJrx3swDqc4K2APE9/nCUDicOCejhJLg+63y8WfI
FdHHDjSJD+mds9ShjLqyCxjw3huwD7gUB24PxZUrM8mcqWuMzdP8/TV7rF5S9RyAVGZW4Fw1pu96
Y5XKJ73vNtTKNIurZVKCHgIiGAVhiJ01sU3ayN12kUVVU9I8vkOzXmuwQtBWN3htzSvZCwpGxiT1
HzKpV0+ZKXLJms7gJx0VGfH50NZwBUi1804k9eNVvHOCyOzrTk6axqlsCaq0vQPnM27KWqd5MX3K
E/IuCmrIZXFSiUHZ78Xo1YlzNT6R6PEhsHUFYf8exsdmxXD3y514hNHpvu0TM50aWazDOd4bL2BV
18BGJp4pCoqQMsFlS7C0dWeWiJZL7MPFRegKu/FA7CQou4rh3eTQ94oXfjaQT3q9d4p6ah91JxR1
efHoAZT38BhIEaISMA3EC1F9tdPio6o4eIGtiB10Fb08Mjw5J4iYgkEppBI6avwMud84arshm6de
hSomfroFFFsjI6bs0IQUpbIjb2qJIO4uKRrARinlnbAih6TfTVvE/ahvFHjt8+ZiznuGiZT/LtWq
bNPAZI5PD+ZeCo808bIk8PCToabuZzem13OPLUbKZibyX76zzdufh6PR+X6cs4uFKGhDpCR8IWAD
6hnMtDUTdDgTI7mClQtvD0xE6zFB61IX3MFLb1O5UTLTeFdvlOtT6RYD3IaFVizrkUhwRC7qT1KD
unQbSIEtSkYYqwUtUD1aF/js9mO84pp0Uoq2iHfjf5rNHBnxkQB0vpkaZys3IjZJ/VyjzzAkxapF
hqIyDRb2G8KDGbLiTuKTLb2c4UDIgiX1lSisPXJrwiwu+j7SOoVPy7VkrmWzZ9Rn8xxe2+iYVj8k
KpgvfZLRszFmEHJdgKI6uJL5UPOvqKIe0zZreQy5haTcdSxHIRcEr3DRAW0P9EfjjBLQBdXkze83
NgR53WI1+w9P5e4PA+5kaa+/WmR4lhIDpT0iZXzWK6SOxkUvNO9/ZQYBVS75JtokT8prnxuBqe+D
ZnlmQiggtrvPpm2Y+sB7c0+FbpROoRs95S43buNu8JpgWXqaW3lEeAXjtMyv9UslJuCCP1bixstu
OsTrnxbZ4IoH8bocE60WhMsVnclT98gunOSuquMIpGlkdqqi2S0dnH8h2uThHPzti7eEw/xnndj3
9+eH/b8+UGcHPjU7bqqPv8Yqgs9rp0Nh2sv+e6SZDMXPGvl961RYowId7Ud1qrNaji9aCXTgOSub
uvWhf7sL7wnJXXe6y1wnS25mM8SrFdke11AKQ7T5lWNOrlarBeaVZ/68de/G3ipswyeYP/owXn/E
/4zzNbZVrgbqgk2jcLcoUJtpeDY820TjxaNAcaaR0xxrg3ES/qiIZaHi0LzPSJN33IGWIrWyESkb
sdhAgO94Uys+jkJNkVNFB+fUabUE8LEyWfR+LOx2UAR8rGZDji4Q9HqrVWc0N64aIaH5BNVj9Fiz
2Ukx73vXVRXfwj8GCDQ9r8tyEpHP0Uiom0PM1XYrL1Cd3Jn5114nj0b0EvjWFn3lwMdirTYnp0K0
8ucwOpz5NvFikD/rYofrCRplgNz8Fpyhaqv/WaE7eT4cN3QRFQ3raeXDPawAIPxHyPFdn9IFqCNl
8Ba0tu+UZs8zmP7P4rW06IQCBpjrIQNRhP4Pii39ClYkLCdtGT99A01J2AQDhrG421LJDMkIJPoO
x4yRDYA4k7KSvZeg8sqUp0A7DCvjqE2bWKZHcCqcXnBevs1EuePzaZ/GstDoA+7aIt1IoLqaS45o
T+n7koJMqINJB4oXalHJ19Fwx4LvENpixnC1Fsf7QLnzuMYzWakJHAd1H1IM55TUbbirHhCQF1h9
/3edLC02EqMDzeJAGQz7RztAEnqoM0jpyn6LfKyPXqvJAQON6yryub1+vpiAwNWdApmLIg48XiBN
gT22WfMU828ZdS1VG6jSPMqXZZQWwYeyo+kUB0OnQQYH63MKpKBQ84/vxywbMdvoZCS36nWWMJD9
bM+ZmgwAy5NWfRneSZlwvP+69xgccPK8x9HEP25U0W4kPr7c6sxqnFCenNi5U3s8+7rB1wbvK+jW
4QVpjyGAHaN36dWuY4sWMGdtyBByeYzV0FtMSEYUT0MX6Xu9/oR5rL5WGzgmN1TnFwf0Qz7NkO8D
Vo7os9FHqVq45eF4X+rwAWwYibDBokbu1t3c1e73TG0kb6bUEryDElMzZLkqnyV/Ke0OW/5R4Xop
Qyqd9oSj8qX0r5Mvo4X17x4x2B2Tv5w83KDn+90G7qr0VWBiS58+oolOiVabPEhaX7m4caMCMb8b
lRFvIJ3uyO2YCFYjYd3bhL8Hl1J0PJwUAw/degnUdOb20d72wZB+1nm7ra57FaTaumJXsf9HQUhP
5zvozyUOAOPy2iDVgSIoj3qGeRCJypf3UzgxyrRpoOSRt+QR7IwoyIoyB+/HAWPZMd8N9K2jEtO5
e3x2C52/3e/UVJz0GmyhxmIVHsyYN9b6/dsvS/gdW1U6n+lulwQ/9Cle1Cnvv+nccWssAzom8l17
Yiuo1HTOyjT3voSjp4piXV2j6g0d7OzeOhl43CDEbS7YCBZRda7xb1Dod1Z2i2fjjEtSXeIthMi7
RK0AvHWnxFcwu+tNyEmo2GAJFb7rcEtKjM+EhJp9BMjnj24/9bNpaTPo5gGkeCarIXZ4OSfV+YrV
Zrlxp+8gkPYWLA5q5Jf8SLptJV/rIJp36Kp1d9CHldgkkogCgTFsxqt7xOoUoeK3HzHeO+LuR+/A
RaA0f6z+MFVdVrz7t8j8KZZTHC4135g2Bas+SJHgjZ/VAKl8zIS9ECh+oMWxSDQqNYmw2hlRGOnP
AJUFxSA8zBhOXb1hBnEyeLQGajbn7IrhYkr6WlXdGVNycsgrdhKmHOKlavnFlV1NMRpA5lrHBMP6
P4q67hFfEXHC9ffp0HkKstyGw3UZeGmK3D0RF+yVVkSA9DKuzwEX4Vd0x3MKBsl5uNpcYSZ7zwgT
j3a5/YBoFBV4rGQ+6xwT/QXMtNzz9e9JYrjs3p0uR+iBMuxxH6I/u9jHgfNeFfHJzkFuiQ7YG+l1
l4k9RSXd8NaweR0/f3ZQ26SyvWhkcfkBXNDREsjZON7AdcMYjlUpcA+ichapyXSV83ss7E3n8CYD
MIOT34zaFhMmXfKQPj1UpozCF/n82VmGAMNZWO2O3oaTYWQOrQTGgJxywC46TlkjnfxVI6hYMR4t
nkG1AvKS3fqItX8PNtqOLgtgT1od8V3rDdV94c4HvwoFn7h/Ud2rnvdrRE0GNeWaamSSEMW2PJNs
Mp0VfM/bb80Xi0GSmIi6YPo/ykcqfLCX4nPiNON8Cvc/ZGTIeI1qi0eoPWqtKjLCiyiMK0J5t4WK
Sk3yYoRUk5LiyhLqAx/HuAYnNp1CfFjTmMH7S8q5iF2yrWn+dvJ/aE4dU+h/1AHomhRp22tiGe3S
JmSRjWCwJSwSCK1DTaySwycaFBCSOpRMbQ/cGC/EzhWhIqawWjmRoESpsu66ypdakRFr+VxPmGFz
DSr1RFoZohLn7Gk/2dDQrhislM5RLqZ9KfJCwfNQuDkJ9xwVAS82B3yMhTSU+lY3L1if6xyP79Tv
ExGSkvTzjHZHkCYSWMJ72qS2LyelWmXWN5i4EaNLQiLrZs0EHMQLKJS0VakT3EKy43hyDxgvj/FZ
+NWxnZCxP4Hb2HH9jWI9wci196m+E6jKQ2ImnMYjyzNQjyuBYt0PMD8yJM/zVDis3n4XhmaShenB
pDc1Wk/VP9horYOWcWBLBS8uGYy4f536CHbbYc62nHYWM6hKnTBV8rqB4AJw67C8d7Bgwy+6H2/D
9gniFG4XZrWWo/TjGNsp1/WhBN16MedSZvAferQerGbS7DV6w9MJ0wbN2Q/pNH3kS6FQwc2GAQqR
4SszPcAKzqBrnFZthdcbrjXaCdBztDcUrFQVZvNGPkAu1toGVqH7peuPhyAJ9ciMtbxiWH1yh54k
zyEyRynZPFkMqMvCP01c0MVHuX2lTNmAuOZg4SsEu/3Fpov8lyWR5g/WIz8a3PzGkvCrDVWacYF7
v5FEq955M6sICS3ZPcD79/vZeshEeUdHoJL4Opdt25WHpF78Q5x+gA1XUnNoPhsiVXdNQKREOIaT
XaN5k0o3nGeY+PC93tGkUT+wepr3JOmfYuDaCoIf3sSvlaiADM1jl8zdZ54b9dyYGizyriUBBrH5
E256TVl5nB//W7JjCQKzb09XK1vLGtlA5TN5zdg5nakC4QxMg08AwZ6MIbunvGqgu9An0lowd/up
nK+sUtQ7R9ziN3QHOVFxvEV4jdJOUiuo7CKzJ11MHAtsJmQ2Rl8PcqlVBum5GOi/W1S/AWdNrwGd
dvC9CyeYEuvGZy2T8+MN/tXx+JshPViHiSQAlnjHLrULxHtFeSH8HrTxv4ANlC2sC7pz3tHsC8+g
lX6PJNp38gUQ6YJgBbiLM/lF3NlG1qsHMLcORy2udlg7bpFY4oxWDrpSWRgBtNnAIJUyh3jTO+PL
W7c6UxdZZkM6q8kiihM/qgryN9737cN2tS5zxhz0uWapoX1d4mXpREqO9D2suZtx6NsBAQoiehUQ
jhkoIQjvMxqznJHQmaLSasxrR0jI+uEnfh9RyPKzM6cwgSZW8d030tu4kyOvdj1XdxXPoAcxqiYZ
V2Yq5drjn4O+cfisHEWcWfgn/I9FUWrLjNJ/SsCvtAYuLyKLsGzeIMYqguU2bRBFbMaQZUuVqikX
DXXVuG2SA65Y65kaxn6ZdA0tWDhB7QckinHzkvsHCnoTlPnNIdRBV8qw1MYHM+WFDtk2cQQW8PkH
j45Sqd4Q62E1/q9l2HUvPhb1rFrMzqrtwu8MiGlcooZCGkq4kMsK8Z1ykRrRdH4rxD2SK63Gj+ZD
fIzacgYc8l31sOIqZ/ZX/ODhVXJjDmAyUH25mRdjYMjR928rAMaYW0SNcIvmgv5btnErFgFrWmXA
0egEjz0KrCooBE0yqeGjQdfhkHasWDOW2fJUucw0jQaZJwlc0A0EizMWBx/DLg+W8hmf4pQu7xXQ
eaibqvc0VfOlMGDVQrdpIzroAHjA/OYRPVQHpEng4L3Mbo7S4nyILyfIaXB9nJk9NvQw5l2GmztA
Gg+sgD4eOn3k6NvyAv4SFsqaThZ59P4u2NveUtodiiY4ZM0nC9EatS63wGLXA3wPUfU5e35kkdcX
QCqbUZwaY0hEFoEhZhgAUhwAFpl/3hVTUYZSoO0hfOWhQHh3fKOstZLLq4LqTAWStx/IsmD1nG2s
xXNkZFvpcqrbt31JjEcEBGcmnctm3Rz1XWPQ8Rt/n41N/rHa+0hXH3dZFQLP9kYkMNBKBKjxPcSJ
1/FAf5AMsvFUuEEYdvhBdNFHCFH9fKixRYhD7FuvT2ESYjf/2fHfmBB59UFtl9qGHny7r2gm+hep
KPcFyYW7SD/qYSiQUpb2XsnbRsdP7OAUwQRA6ffV3BtaF/cQpUMnNeXMXi6TXcN9rQXDjW1ZtAeh
JYGBtnup5eWoSzZp9XHHhkhwnysOsCAVKfFUu/W2Fhx1/fblw3NgY/Tsh2M6r0uBX3DKgggFSvYJ
8q3cqWVLoE3y6EaNPePtWQBZasc1yy+FBS3IeKP7333u1zgzo0t8WVYsqVUEPxMGijKM9X0gJCbA
/btVJxQ8E0/OgGNOpprirC4LgyCI+ztK5IaArJRwCVn7YSUYxetXG0Uyn6rQMDSi3sfLruj8vo71
fzScfE9tPGd6+fVTSWvS7zkZesWjQojZpvCOxYDCH9zTkARgux2qwsWth+k48UozQD9YJ6MU0sCh
f115nY9QVrXh74BlNv6Zgmr2bxGW4rOXHt4h6+fkjSSSwtZWfGwLH5j+RCQYbCca3jke0gUsKYdD
tpEmri0Df85sIsPyIQoh/IxMKaJ9lrM07YvFHD3NjJlbHmpFgL8+BJUA+UaRdSze0XAasdeLRbxb
ZHFEcmDS8ZrRMKxATpKvP/hnvdbVws/WhMIcfQvKSOeGFyW2r+IB+LNYtuyLpl8Bnw2sHdMmNSfv
J1QGq+5K4uxoJ43tRxJ8u+0X6zyWJQKQ+OIp/9RATTRg3u4eU7Rr3vMnSUs7q2lsYI+Kg4POVhx7
1JFzFs02zOsIqUYj0ET93Qlzwq6g/hdfstUuILSb/to94xrDIWxiG5u0zvoTjmCOJcdmS2R+/P/z
YneM45NALxBF/g+HUTZKybmwRvVjc3MPsxj70KcQHTqKQboFIPFSnTo2W5d5afkWA5d1K3Uu9jOP
zMNWHDM9Bjrr+PHUvG94AvCp5BRMgRFZ3KrzpPB3sYl/aupGuULPBSkYOeU0+ZL1RBAGmJxteu/G
K0QYaxP9v0Avja8UN6po73/SBZI6Yw9B+2MlWg0VNs9UBLBbQfwt6s3e6qKwboVjfr0Egp/xPWyj
qUUeca6qGKsndOH1kgXBE0WrwVkiNDmtzinVK6f8+7SQN1/DKcHXGM811AoBtmD6VzrVytveAetZ
67lIILqN/AtKNDhCXgKDoKyFD9Y2cbYSVx4JdluhPS+cFzqci+6du5VD05Y49kHx3+rESwznhRYo
frg0RYZXTxHSrF19RCGgnPWZSDgW0WYnoqB9pmKTY03Fci76xKXNdW4SJ9ayCt4PEEO5RF8SmBv4
g9YzUy3ZXbQEtt6V5uJq/hLzvKsg37dlByEg+zoF5JGKcwmbIRPWfyZtd73Mhl/TrJdNiRjYO2e+
BNTxOr3pNo3pKRzWWVht4b1E4nauQttxlpaDXwCAyVgpOrj+GLkF/lYlwFWrE8gCCr71VogyNx6y
Yya4+OpBM2wNes18dfvNv+FPu0Hp4PwUySe7HFbIMmBYlzjwhf2y363b4DF+BhovWtupawXxIMtC
fh11+IuNiBG4e34nTMbZMTYij6qgQc3lRleCb54qqCaYhGOmVKPxYEOvLO+9Qcv8m0jBe8Fs9DCR
A4h4xvppmGSSglwCcZTBdXPFos2vEd7Fi+AjhwDbsRIyuKrk752bbgGhSruolp3awF6uLyvvP7W2
7synmlQfdzojHNlq+83F5CFiI44vk2TzhZ7kqCZ/p3PUf+ZoSg3JRgaCtAFL4BmwqtXTpC4qF7GW
h3NUvJPLnBoA2ndZ0tkciZ8Eun5pjfLF4t3kdIKQA+972L0348dKbOWqPvFuvQQRe7Xd9AZGLuyN
IBB3mNMYtMfP3c65bLS2Fi/xpoXBVWwUhzajZHnBjRDB/wVh5iN/W+xLOjlrqMFJoRXbGUTq10D8
FsWzxtN9MSv2aAQRxohVvGlGV4Weh0EhstJq2ll6HBeE8dFYPxm2sj4fUSRW2/hNSnPtyiFYyQGT
sGtJyOQk5jsOeYkSZf8O9eUHqySQLAWqMOo11JmlszLGvKdpOHk7fBcnwWMki/bsqX7g9A6nDtEM
SU0EYVrtDBAohnkbvyJ3GcVZD0DlFo7MSjVOrh+Iu3WqEFZ3CvqRDcUremud3+2hdzlij/Bog1Oa
yq5c8F9/B6wMU+BsuVz7K6d9fVDWs6aX4USA7pfvNhFfvv4afyY4w3u+o9XG8S7Iax71FN0KoVU6
aY4JnVK7yW41wv5EhckugC8xHj3POQ5qQKS5zsYIdfE7wiEN18rboJIsOa3EVc8IcIo5kN7DsBkO
p0NYqLbB+GMIm6RpZRgh9/9Rf87PXG1RW3TmpHGJzsJt4WQBe5C0BhkdPUxchuMsVgy8vbUPDwGf
RRhxiu++lIBqFyeKagSUq4dyXm/qBh22JHsksul8LdPDj7EI5FIURq0xWVMU618ViX2lQGN6XBCG
LSKJQPP6iLBgjQQSFCbXswtYxyUeq5OxwnbXBDO8PMCPEN05dJ9jcbsazn6gO/NWtW88w/DK6qtH
lvGZEVBfvyrByUVNPiaiqkhPQ3FpcxzlT+UG12aNHeyk1oaxRYZ1KqSkLBr7fkyzIGl57jtXindl
dl3+Snd3J6sC6ZIXK10z6nlfuAZXfYY+nwWuEzgKvesJiD712Zq6cRUqMhOma5NB6SClxDgaOGc3
rQl4bAEkC3/ciIcPCw6SHeMM4KoAmbiT2aHjbqTw4uYIeH95FBFCZ09IFyH/EFFtJJhQB0pZeOR2
ywNLGffZPRmfC4g9Uql1YyVc3YnDgxd+rtv8pKEb9e0CKaLCPwMUKt+AWxiho5MgVtMZwQwa9fVV
72gNBhif9cDbTKv8lTQXq19IuRn4rUqsyJNbO1/08EXeAk9gMWPHqJ7hsj54kSShyAKYbkNYdqRN
cO3MY6k10KMRwXLF+oT7XGdAjsQ39Y8ExXDB28Rlp2RfHrfAe1g1v5SvaNdB9jYBbEgeE6TVVJmA
n07TIdoU/pDJ6HinroHMPr++nISODUQdnBMOUNc+wB4M8nKmb7BkxT2qKTDPFjYr3bqU4UWCfqFV
iTjeXJAK2vblrthTW52UMdVJz5WR1kAuVD9zAUTlolwBNi7e1nWnlTLEh+cRcSUJQ21O7Jr6Tw6q
chXglmoP+l4Wrgvd3+he5z27cNb2vpQWroQPN1U2pK5O9K3TKodE9UhsYKTM7d9qFCSMrwuLYY2N
jJrxA4eyp+q7Fe3boDaQkwywW2ri0uhrF4L8+1v06gWIECSMepM/61B6wH6tLjK/wUJQMCJ46DCe
wGkwfwk6UXfjD+hVtty8wVh3qpaBVZWaCaWa/8D2m6mGn8FQM0L59CdHFoLIVuswbBz1MNbEwVuq
gmfIqNYe7WJdbCUBBNuYlJr0A79WsGZpoueewJPaLv/k7+iDtQA9JSkzhRGCnkzBtv0EbuIu1fl9
TlH+z0L+taqwCpM1FCOGr3pnxr46qeUk2i5a+N6KSXZv9xg2EYA970aHHSQF8aUfKuwIjEFikYfQ
0iTISY/ImvbFvBs4odCJTp1BXW6RVRGCd5H1byuHfJFaWIl/y9yvGtPW4xfcE9b2X6tvtkMQ6A0/
PPjBiSVxPAEdph7AO8cquq8YXwFNENlWGJJPt+rRTgiGxXo6vRnpo1xwT82KvU7VHD8TOD16AXuA
yrAAf+S71t7layTgT2zajEI/mHR0YiY8sstYnVOYKjPiaycQSclHZUGdYetRs0TeMsNXlH9ZHqcJ
+Ycn99DIeWHWvYVMLFSnQlukNS0OSwQy2Y8WcepJfXIHJo3xVJWqW1kOSMjq+OADZi44ked3CV7E
4/nEZ7v4AlZd4G/YujDmfWHps0kuIHuze/aTGruvPWwD4m+Sy40Neto+RB9KqugEFy+Mr6MSAPqa
mk2GfYP792dYNM1Ae4J+gQWQQ06xfCMEfP/739ePJ/21ls955gAASGNjFIUH5eP4S6vHxSEgMtsF
E8VuLzlRaBSXX0HfQptM4IGWecryXZT24fDg3Y53V17ULxboQV4S/vf0tz2dvX+UsE8QIcV8/dXC
Kp+pn1f+fvi6aX2y/ttpE/WdFy/8qiBNhlF0+zlTcv9GrEej2AmG6ORhW63MBpDXb8+CFMVL2+wx
wLxzYQZgQTW5LsPzbGGja3xsNnWIzx2wQPwMJpVOto08XhDlc8nyH8E4S1qdCGxXUqzzXAZ79f4N
/lj4R5v59WFnrw09QxFPsNZkKTB7nyFDivCeUzgSCRfNa6Y/snGm4vvNTUvgBw0WjdkeLn6gZarq
HSTG34ezisppM6YWBKfPP+FRIx8CqZPPf7BDYhw7qflhAtBn6ujCQK0UrWSXshxclt9BKhOK7iw9
IADU/+q51u7TAry4DoFr32nFVTkdJv52VQaTf4F6tyoslW9WbQdgYB1Jw+kG35AV2OE5uBOAd6cB
dOQHRzKMiESWwZRDE9UKzQ63oNg6sfFw+8Jg/WT5lwHQV3dSmvxoZnF6Xiy0vUgtyXUVY7sZ66SA
/GPR3+nW9h9X/vpxw84P+J2vJ2yvogFTrjPXDGScJnp/gX3L+jCLjmybdlEvBmyewoQ+91tRjLQJ
BeMAK8nMjj/rawC+NI4jLxYVxOWLK8mWggnXbUH+9HGsBCinq8fV3d28y829Uydl14X1FPmHSKDD
O54qYet6gZhy7vy8F1VU2a+jMC3bc7KOnSv+DS2Bu0aDurAay64w8YxdUhxoAZ7rp4W50L1HK6Zc
vGu/olF6Cs/ZYWqLdqNuDzoxXdEuuT+B9pHT00UkQ56RPW9lf6qhqOTyiSKf/WBt6pDlfFCq7mc5
u1uwOxJrKL8SuUxsy0uIU5JzdPEqJN6Ojl53KEUK0EEzTVKGK2e9eJjO2MQDshF8H0CWqNh1q3FC
DGsZAW11aALXgf4vObxkKkT/lTPCpTcqfC4KFybGAEyeWrCsux2vcfYw/Ab1uerMRKSld12h3EOG
1ON33k9JpdKCrtNXJpxx4gBaMMYRYKmyVvzSf9sEq3klaBRePt95gdboBWYRun7iC2tY6cZ+c34E
VInfUFxH5KbWd1GeWRr7PyEFiDBhyPDdzCLqWB7dauCACcUDlrtOmOPXJ+VdgUw5I/hqiCoIZUod
BFomqwom7ztGRYlSdf725rZZUpCPBor5dGFA76Rb3Ixy+VUQ8tSQ3+a+CGNYQ8luE+FcMrVaqkox
0jbYhBat/R9+saPy1985xgY75z9YduWL2+7KuCZ5a8INljcY3SIZxIvMAyyHLGrIDhyBOw5dae7q
VtjUHhUm5Mo4CcqpDuetYZxjg4mB/Rv7BUJanoFaf8e1wWgxgi0S3YnX/NB355RYbhc/ygYIwljz
fszsJHUtZzFtjDJpZB9EPR6rKwh9XgdtF1Yu/SeKURx3iZL6QxFR2uxEUoK22CFp9RmZbSCyqXEZ
b+FysS1bRextIvrrNAPR7by/QeGbHzapTk/5wlP0E4jOLlti3k5vmijRJoncRv34P+uMtSfJxe5J
g5D0+y9yGCeK+zLsnFGetsMCDN1Y7pClLghWYlPEntUBYTua8fYfpBJEVzSBhfKtfGx0kilytrMR
fCyxysTCeDc76PtR90kas8cCpVCsHrfVHbDWck2LFjjOu4toEKgD9nXvT+DwU99Y9tAfQ/t/DCe4
w+iRBf/31yW86e0faY21o8M/bZEtiYGiSPKamK7YUcRUpBUBH1hUCncxB+QbcyjVrDmXnHEvrwvD
wiF0fgElFiG08DmEesgYywP0NCGqE4jsi4+iPNkWMGvBLeiJwzyKmDyqnYHr+oBtoO7m4MUsHAz/
8Xd+H/Jn4SqIsuRUw2Uy1AGNcGA327a02bPHGGy0zbkGN7lq/ty6qztXsoQYGp9o/3M+w67EY88t
VfTBflFp4daC2xYINikSQl6kLY5g087lZx2mzcAnVPhxV5IOxaULg/bpT1FeSQKWwQeT+J094ua/
4+tRLg+e3GUdm3mo+TVXy+NZ7GZXeJJsiq5Am4TGWu7kVICDNAbJcp1cvcN3+3v0bvey5MhpmT3F
8uQKSiEcphCtf/x9gg==
`protect end_protected
