`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
X+PLjbpLQyVHK2THcfsqD9EK2Ow7djF7nNafejHHEPW5yBtzLrkh49egp3l50BesnqPZwnRXzTBg
FyWMG1gUxBwZyMLrpTMrt3IptUjxYElsXRQW+sj+fUyAMvFTfAnKQTaI6WSgq8/gRqVBrZoMzyPl
J+if5U+r/9y7nO8PxJMJ0P1PNbdzGSGeOjSK9FLMkmT1fHA4mGDfS+hrlqTfeDTm4ljiKauHK5NF
vmhTFQdAnaOV+AodA2eUpEcG+efBqxC7TjBSvl+xE47O9IcTw0Vb4YCfI2m3oBGR8bx8Vrupu7Ma
SNT67LWWVC3NkuDfe3wi4XnmNPUOqZ+iMxx1yw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="TUMdnRRcuVJXljaV+T34akgKMKi2HlEHDmzdQk7ypVQ="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37568)
`protect data_block
JIpfj8yjg1YQIA0mEUhaTQSxCNegxIl6O7KOooI2DIhnL/mti5wXJjYvrbmzoElVqxa6MQOBV/7I
pyfPddzE5hqAdQ2HFQJSv20QmaVDn9cVeJuhBuk9X4JIP3GeF9RQiQ1rd36SJCUJSQ4deevyNNZw
tlPxtM0cb5WDyh0UTtxKxd1+9F20OvFV5/MlQ0+UpG5ddwFL9RqJsbhFn4cNNTDoIdU2Ti6woTg7
KunZmEYyto/6QI16gjuJGcwryyvXmUo46HigZHXwjOhvsINwhlwgAt6A4l6dFfYdlInzeWbsjwN9
d0Kp3WgTy8Auqc9uoztd+EfcFjf6mEbdr3HA59W8gOxAiuBX4b/aT6GqeE76weu56Fxgh4Wj6Bgp
7rXOpDE/y84lZxixMCNQE1JDEuKqFyxcihMe+ENzz6HPwIQu7yb1bC6NzDi0Q4OLd8QhVbJOblFZ
rR9Ci/vKJcGwtCJ2EoYN78HjwDuGrEqLcuYZSiIvP9QjpXvHpoo0zr5yiL4ROWJtFvw1RzNPVGTs
/U456pIZQ8fD8bvw/ZuHS4Kp3FIU7Y97eOEwrzjhcejHjQ7sskLWNzgAmuaI6v9OGauqWyYBeMo8
7Q0V8qevdM/4Vx9sv3nyw1M26ogoyjZE/o9xJAQlH2fhzll9ZaI4jfrF99FA68fnGr3escenjT/m
p9WB0W62nRxVLMMzcUZZUJCKlRHANhn9s5CyA4nFIzX1rwJvoywIy/YPCfXc3Y7rfGa8wrt3I5hv
OAE6l7RhfL4xscNFtQAEQBt910ricusRqbAGz/hvdh8ZCBIuBAby8LF5QsVv/yOYgrNKAgGEqc72
IM0/d2dQisUe1uHiUbJKkM/CUQVGifql9qan6LsK14pbLuablN/+AipKdSuLpA+32UZ8xhk/xAl8
7HjIC/1gk+ZrNOphYniTuXHZr/xiAWLrpc9bZpffb7vgQFVcSjb1N/dO9Xgp4t8z8jiQn0OmmLBT
JJog6VMsKAERceV0IUgRT9ZWB0LMTAZiEsPaLkOGBNj4QxqWtzYW4JKyqMONQjoqraaLezZkNy/j
pceLyCF7YJCNwKSa8+l3oyqAL9Q43pNELYFprpFf+rUT6CrFc+fMoaksbWrIJPo28Ql542tijcLk
X6wFEyIhg7+9hesK/7+dijZl10uuxJOe/ibTdE/2LQenrBFKhtXefhJb7EoHjlH/Q37ZM3ZdZp2o
m+Tnultps4MGjkakqIAM/0d5M8MND/mVMHJirpElSO0GqlLZ7jG/+98rrxSK1Yw6C9H2Yc+QfBjA
ZSRtup+WktY1MfvQpeZTYP2XejPTlIutR1i4s05n7Fe2sB8UDw99AiuGyzUCaH7+WI1xKPWZgptK
8xBKUqVMlGmixiFUb2KWrWOUk7gc8PnTmOIERu4vWGdTfFa8jRYtlgErrmTrsqbSP+in60F1Bwcx
ryz2hmQ1EVFYCQms+17q+6pPH8ZMXgK9ZoGhe6FK3/BmWZ4LGodfXNlszwMk0HotfpjjdczO1ZTs
XyA5MG7bPVC2vPN4wB/CvCxK8g++lPX2Ti7b/hoE72f5JfOHoNrQiy5P8dV9Pwb5/ShY+BbzhmWj
wleq7/H+H9nguj44dI/h/+XEpkrVN10MbRe5nwE7+ZMFw1L3PGPJsM4o5QRQVgXrNIVSiZxcKVmC
KxWRKH9T7PSnG4zSP8O94WmTbimWkyBTRcrpcIWsJD9n4e5G/JnJhu9T+UXWhHimNrm1bHidFh6G
aGLcr+gCIo1hupcX7f/ciIEM3t37n1QOr9fYdmPS8NU2hsn6Nok7YXeGXWDBHfLPITYyVZvDU4f8
jTVppg5HC62l7mCIpTA3kQ1l6BtNCWGk6b1a24YAm1Y8PnnMb4UUMKaW5KJZh8a0k38roKJX/qgV
7akODfSqvRQfzfY4Ope9aY/POP9LYUifHU69hskvgEewVi3GOw0UdWOhMZxd9nXYA78RXUtuE+o6
14LgE4ipoADynvCvXgyrk6m1BuoWd9+BiCfO8aEAdIvIrHhtoPeJTluXeh+9aBgv/z0LIeY9FhKA
s+7AKMN6z6F/LC/c9urcneSkeEm1/K9rrEs5RMcb4/+ewwPrDEi3Q6cwttUAy81T6I4TQoGg4xBe
WGg1Hj9yqPabSey8dgfTOsqYmdAmak6+Ivoyh/gRQ9n6aQn15aNWVa17Hkx8qx2/jDkTQgKsStSZ
E68dHZ8Z2c8lhVzFsaEz0dqRNZAqdGsWBIJOmoYR/d5rPZNVLPRyiiCmlIUWOKK5YJK2sHWGRFfw
2YitenI03DCFA2atjF5VTIRb4rObGxkAX+lFle5P2/3Ojca0qSfFGc+DQb2/SsKAK9bi4MhZJFec
NGCcsR0srxCk8Oo4Y//yerD3sXmdaekEZctP2+r9efHpN7KSpOCvMbUCpz+h3eyFQ9u2nMuJulPY
cMa/5cKiM87aQV1M1r0JRWIsJn3tF9LrhwQe3xfJlmmcmOPzUmi/ggw8azb+JG82KIdaNxlti3bT
Ca8OFUshjARjZfUAJLTbhLa3uWJKVPyEkAhL3ZFR6yAXm9YEuNNNL1cajV8d1JnHUXxWpp0rkNh+
BiqmAfiQaBFQ8zzalHK2j8qj1XMz1xa/P5G4++CapBfw86qPWwIsj8vv+vSC76m6IZjfe3k1vWO/
LC8HXoCH5MqWv1EAZk/mrNSxAYoYzdWopFaG/rEdCvGppgN778MUAirnMFBf14F7RYkq0fo6o7wE
yswqCHugfjdEkujVb1xZdHwImnzXh7hteJM0OADuOgEgaMfBwPXe4MyXGDywo3lcJSEqgI3+FH++
8wjCt9JgXd28W8RearPng5nbvgexiSOoks6wLV4T5G5NE52bKIDkd6wZ++JaN7TCW5S2RTD22VyM
ZQ31hMKxT//N4dQdlyMjYtjPmHMhT5jUMoyQlPCUiYRjp4aGGO+1+1GqZxWtt/Bx6wkoZzOacVF7
jB91dx7hn4SlLJRteAsMDjE8jPY3u5X8py1H0+P1YKrGUd3RWPkZ5vtnDpViWqxVSIkWH8qVrg8z
DzfjSjUdPh8BPtwdSCuZVyLN41MNjJgKSntpg4rllNdfAzPgCzMSfSz5IHtzsi5qttYsIhVPTPXu
ldQeIrDqdqmdwBQ4V/DD5Y7EGnWUx4J2HmQ4dLCpMsdl1cHq+ONEwCFmQsMVnEtinPy48DjHgWNM
vZjD+P7vK7+5TK0mznzUZMyU2fpavISU/hkyvyle8MvueZzfXas9bDX9yRlLWiIM/lP7UOfP5hxw
GVpesOWOt79XRSsV4WMSrFLOcZ/rw9FdPEjvxAwLr44Hrz2x4ji0rwY1M/1crWZAgQGZR2I+gMzV
KHIujfFzcsX6MfZyUM56vfJ4kCUFitl90TdlDumNQ56xqo3ZDo36NexyxQIKt4PMknCUG+tm8q/D
563PCoNzheAS90or1F43sp+KWGdZpBbyo6E/hYIBteR7OhjVBaOmkSn8BCXiuAI8J1w5Jo/zamnI
6SdxhzNnkOjftZ3caye7NvfEDg0MBiYGebAwV2rWvjGXLwpjNwWFgRceKh/r/Q7dLkl37u9HP9nV
UKJy4e9aMgSs2tJ6OekfxkJP8CJh1iA2t5GgZ3BVjYIATFg5qJ6flHgA/Ebk5U97Yk9wCBKvqVR3
DcfG41B2TYb9ErviDMpwlTTvznIcldBeYiLnKA7XBo314iGucW7e+G8iDn95986F/jdpRD9z5AVO
WF5GkHqyCPTsJ+Tz21GC8a1/58wDJ7OFGyDlCDEDwF6ZwbqixGqCY8Nm6Qc2i8Cw5xvnt4TheU0x
sRRDePl2cdRqze6umYG1O6/4sAiy5RhzblI4jBAC3N0jkxfcInydkoUTCoVmPNMU0JS2hrV+17QF
PfuyJP5g40Wqn28sHnFcL0mRIJib+kn+KFT6nIzsm3tciGhr9HmR7jGeXMUScbG7MGMnyGJh7KVc
/NfPb7EYyHp8X6OhxWFrLTVfvCLfKVxHDkbmaNeILj4hXh/LPmxmtzbctC9rVpmoSmELqsS9GZBm
14J8W5Aj5475xTkvow5m79ltlkXGJJF8kNtm0bp/ROsw6mWR4DK9AatlLy/EYhnuG665TkWMzZ+A
J2e57hGjJvrLk4t96swIZroLJkYwiXAfS6V3QQXZRG8/f5aGgrX9OX6A0BBwJwODyroLLLDCbd0M
0RuXYTwSvxSdMbta6ntIDr9FbiKWUGAE/i5kdFepi75AdlaRj/7/JUprgyexhGGQSKGp6cYa2wBd
EdAfmyQH6LX5PDNq5jG5TRLvaOYwUiNyj6c9knesM+cdcvnb0YiiOLjNBE9h9YNcA1yaVHeV+N8c
0oCUISTX/gOcRtPMaor+uQ8uQ+JSL6u7foE1mzlRrG273Dl4A2IrtYEBfjTBWQdMsZrj1KE1kim/
GsID/Uy34XpaV0wptJIFisPFI96ubNyYuCYdSmT3kQa1LlJ6okrW5ejVnfzi/ZFGYWALo1BLpOLT
EgpYrtg5z68Tkx6APwpf8xSbmq5exJlzuec1n8V3ATw/lgViQBYPJ9HAVs7k9XNJbgNK+n19dVn+
h1RR5x2syKBievNioPDirJaMw9cfyrW/rJkIstlvICWLsPUKT1wl2Py4Ftn0GjnTXUW6ctjpfnUr
QEreTp/Fv82kJF/Ccvkc1tqyKuLFY0Oxf+2mKa2F8wp9wYayu7NS9GIzKfTS1/hhWLs6GHICqnyv
dvLu9/qh402jY1Mi9neDqkDyWOl4rzLL3nDTdiWH1qTIGKcgHSlAFMhVhrQlCBpBHwBep4vMXZlo
PFFeJi/9a8yElLFkzPdLdMkSXMyoRI2RhH+kcnxFGzQoORC3YMFempLbwnEd5EEWFtCa8MIkneOe
tGW2vo1ESL/tJHwE4DP6vP4evVmGf/OTaGmzwkZOz7tCT/lpm/YoPWy9Q1NxXgSZbJhNer7SQsSM
Bt+egS4BWZj+uDLIjqqZ76Cu8yuocy83ph4Z6rrkjsQ0ikZsJ6g4q49Ldoiu2KSSy4JAfBBhy45W
B+ceajd666t/cb0Y8mm3ma7/ekLadISGgGfINctzfp8K7sNVxwST08ECIOWC6dKjnv4IA9IVNGvd
cVfsEu+PgsJAfK0gqmXR+3ACukUPVzKH6pQS+qfhGZgIC5iw40k2uUvhxvUsH0ZwwaYwiOlCmhYu
muVUuPLwiqVrq5pUOu3zpoN0LQIeW9IoewvAv0CQB7+Ee2MD7CN2irL1NyuJaTZ8IrTguVwuyjUG
d+yL+qH4o+AjaHVNL54mhP1faVBHnEUnhNioCOL4juzum7IDWcD+m/28ecfeDTSRObGm6aKwSYoE
j3maZNcd+Vqj9Ek+pqLFgS8jeCLJz5Z5COSAd3JdJg8pMur9yS4ieVLw5IYIGXwcDIs++YcpKn/a
NeUZzVjTshDL1AYtqxWUKs5lE3SI+Rmqxg7bfDXcgi/jQH93eTkJycBxsb+wnySe9091xK84ZrN6
CKAgm370/KqjSgd1BAYgsN3KsieDnCGbDxabhRJ0U0d6APd6FyoRoGweSr143XpT0BQgZY6/lhu8
UVzaqmgEfzyaoksmFdItidsE+CpObDFRKVUJGA9nrqG6P0COBUmYp8b5efSEjdKoI/M7k9ye3tgg
NuoGHFW01ZFPTupY/6qJQkS1tYZ73/a/b5nLE3PRw9kuJAjrpj0p6h5p28kFwO26luhkF+nRsiVK
bpFhd0yPMbqSdx2soOPaeyw6ngjaeuNZuZ2qxYtVJS50L4kAlgAt1zTPELEO8jEhyzAubBZ6CXXh
fMQQNqBUcFMMkOjfnghSCBXbowkKm42tSjdEKDBHJkzotv+btCVh/ynQZQtoXCayHWLwPUuFSeMx
ZJgwdZSjtMv2EIAc5QVNOSW1bzYzp49EWMpBPmdGUCWvLu0v3xDQDAjMmiI1HiZiV1nr0QicIkyf
PTdC0fDQjudWcPkoDJrWP5m01tUjqcFsC6UsVvN7BXs96WQBHGZMeJ+ORnAE3P0/tfkxUCKQHoVe
nrJyI8jG2VX5sBFtiqzgtG9laSBVhYA5IBTaH6tZ3CyxLP7SGmlb8brlp08XEs4MVtk6A/OUgPqM
KWYVuUstN9AGABcx0faTg6yMz6vf16TRZFd26gyte+6MrH9iXeVyOzHd/qF15YdpVgQpCOTsYLNe
w9P881frUJHc70ck7PQN9NRVOYE7e8gUzyWzivJVb5XAx34U7Ahx3+BsUIHlUfZxQzuvudRHdK+K
8CdOfNgtuvIfm3ndKvGthJ5LICMfHrA19mWz3fJ0r/QwDNLl075sB2qlUp+3DDy2ZEwT7pDw5zQY
H6Vmr4Ml6rNcuYfXW8Bv+nKnOnbLJXlaYvzkuv91G1UcpiqLIaHoTIjizmZpURQ7Uy+TcnPl5++9
YTdaBTDfEoXsbu2jI9MiRW/6WYhibSc/TkaJPH9EN5m86rcxcMDC6QKjy0Y7wQGWOTkhVwE7TLw5
ateK3ySGgB6eD3aQDEYHgjGd5ypKXo8LwDo89kMUw4Tz0gYe+ZQV267bRdu6WAHpoyJO0TfcF+ty
7xO+jiaG66ml93cYikZnu7PNGQG84ejxGnutNFX2V1fbTo5efyaxHOTtYfHnExCZ+/vx8zoIYSie
FxIw06ggDXHyBuORmiPUgSHJIp32GbFIV8hYMD0me9JKxeiP1WXG2IJTWhmhYvxDLdpFEh64+0r1
+xY+aJIsnXeMmcbjAneUtrUl20TmzbNVwkbyCeVIlTxQt3xAPSxsFu5A9sCg8T+L4TK0igUebmyQ
j04Nzvn9eAv7I+hq70Jd7hXQOKdEPilyIYeaEKD95E5Y5ZGTn7h479S1f4sucU5vwh1jz58lcFKW
bc+/Mt8VTkN+Wa4ujvB5O8O4ETeha3YUpSM7u5Yub3xF0lXuYS3ywpT5l5wCZvjA2FQoMfGyv44P
JzpXgnRjA9ntz5C6cNqW6z/yABIBQfPfFyzD/6VzKvBiATQP47UEmuYIP5QFaMuiBHDC+rip7aWC
SX8p+lH1vjUFyksazSRt8S8+Wf8Zs37dzAr63kGDu/br/WCUIquE/mZvmdi3mITWLZ40p6IlSMVr
rzA4NumBeF6p/5QK6Vi0FZZFUiJ+mEUffs1IHLSVyPTP7Y4rjoF89IbVr2lQpKYwWbEO3zOIaFm/
047CEdYxT5orfcQ5Y9eeK62fp5KdJDuA9iCC+hivnzYg1//4+thOb+Z0Yf7qa5NVqoLRYfLe8fSx
mW9PRqOdh5XunlX6I/qwY/BRL7DrTMPEW3i+eE/Fdyviqelm/JsoZHqZwaqNn6EVs33IkETQTEGy
IQwhSHdbEmXOmZja7RLI8F9x9e4n207WHgaL29MioOhEJu64sYxBWC3zSYjn0w6rej0kttXJ82DP
uThMjXO0JbrO/UIQGzYacXl1lffHYU+rXoZ/G87Ffbfosh+wr0MHPc/snR/vxTRC6skk8U5Vqwgx
QBISe0fk50LbHfDNqJkuQuwjmoAig/+2EggEn6BMP9NV+eDcS5ZDL6MhpummpKKKKmQeiG9x6WjA
Vc81SgWX8aZ1+REZ3Sern9iuBgVJ16oimlD5NoK8NBHMzdoYET9sya0Q4G6CCDq2kufHRC3sLZlP
xF4QLJImy0djm5BGOaMkZBSi81kQFzvZOk5spDbGpmoQaMNOCxNA7YRJ2/mJBgR8NEplf8Xw04Dr
V0CVIrr+EPA7gok+NPYOn5UVNWpRz7YkCbBycMrt0zClY+1t7mDLc8DKMm0hzbEiYD1xVSf6O0rK
zt1Kewf3DSxNrjShpl/VyRxGFxXG+ZCreaLqWX9EiUk1V6gi5IPNcELAd0SrM/SUJGm2ODwrsU2R
ymSWNkTBi8MzxvM4SWRe2pqMS8/sv97W05ldJd8QQK5VrW+6rpXc6EPb9HvOCJjxcakDYBWzVIH4
ZKocZQQX8e8qaG9ggwtskgpgvAHmo+SbpEdMLD0VksmZzVbPk1darzU0n7jTD5tGEcxyVrMBNZb5
v/vIDR2HcP32pwpv1fe+AneGPGLzGZ2QYx1aEWqGxRsrjU4UE6cOM47YOJOW+puS3cyLkfpQTMG+
LwPQAuZJ1eBRyRHIoGBR1kPtEKjDC0T9o9bUAOz2tCThidm75ae482Q9nj8pGjiU7SQ2AWD9YXsc
xLjBNHKZxiHazcevP9qePUyXlT6hBwyEuhSMx95VqGypzfXbZhivaH8UlEk4Z4sjOtPunaxESUMb
63gRoFvB7EwmiAoCG3XOyGOWilPSfseUIiXd2LD8MaKLrJk5xjRYHzmvg+Ggw1HyA13ZzIDgYZ2R
Y504+c/MYQOZafI7A4DsDg4+u3G3sj5dRXVPvLfe+wYVU44q2GcNzb78oe+Q0Oj8kbo6bXbnJvHA
pQKXkdeMmyNd7sHtPjCupNxbNNBoUyHPQgvchHVO3ZIsczIgTA6Bt8wHljBr4U9cH9ftKD9+5I5d
Of9mA1+k5dFUOSxlmMk/pFJXbnFM5YKJIzJXjnAaAzmg6Gt4IchU7K038L9KMdiTVrEDmykesKRv
cfKdorBdia4JfOWq6zifgAb50BMkd6UcDTHwRAlvHepcfVTktG7yEupRfFAX0+ybXZAtVk1Vm5rH
RDeDNCMjucb7lUEnNTBaR6tNsHf+UPOC+CzRQLLnb1g57VjJZh7ora0OOH48Qs2rv4xkMAnNaLMx
h2MVCDRfCB/FCDxkhCcJpDUtLFbLJmKpjlquFjVr42+iVkezx49uDERl3fi44JU3fl8/4PptpDWz
LfPJeFHjcjspxKotLR/MWOMJ+D2rzPbUmLiydb+BnmoR+GJKGmWovgVxXMUKX0o2U/Zk0mlnV8XE
celLmH7wdEGh+T5Jyw7aalHXaX+YRZaskFjzt7rBdefi1wtpvNc6IsNBtbSPzEu/KCudS2qwXEWI
w9NmB/f4jRbmaB2cfQWwJxcqgL8pc4Vd9hU56xQuvzSi5VbGDJGPiZ30faxIEOr40U98s4FXRrhZ
HnxsTPIqxhhrWo2eQJmmP59Caj9wDiNJLCRzhR8k9b3FK9+1jDFidej1xQOG6JOOj/C2QtZ3o8Gn
dAf3/rMkymNWMbhAnQ2wkHW0/SC2ByZV4qMSDQVW6x3X+bS6q5s6gu8WEoflHOOQogWtWZ1UzbRG
OoPvn7jOIVd6jlVj0HXyk5bCvjJbyHB0CsKDr55ozAR0yCumUqHjtIOxbSamQVgDYFveRgWVmORp
1lnM5ivQ/ujZKIowcu6aXP1QFMSHvdQioIDCMCN7LlnzeqxQL81/166Tu6pAQgZWEBKtaRjpa8DP
QTEPI4X0t3yZ5UP9YWUEFvmGzNkF4J3Yn6qz7yDLP2mnroRu/dF9YNy8CCBaVsjPE7VsmzDPNr0+
CqIlz8Zt1v9Ofh79mVpG7xshWaqWR+rkznVm5gS5WVnNVeG6hO7DkWKDrLn+Vooard5orLoNKJ+T
fZ/zjMjQN55wyJi4FPVT0ad6kB2ILKL3BlArF3+RzVCEqf6jaEJQQlGqm/BUTgfGXtVeixhgOh3r
k3r/lRaW2WNfMkKXmP97ZNAPc25JHo8CuDtYy4G0hu3uMAcnp1m+GVArhh7ah5Kyf8RIuhauBQBK
jQo5rwnmHf9XlJm6LFpkHcbUFy31RxTlzQc3XXq221PIJGgG4V4QxcGbymyFsRrciXgeWd5iVyf5
1x9nygHr+AmyezenNqxP2T4tnzQKJ5p364SiM12ULoZEZKkxpYc7yFIazTcis9vv2MaaCABBukVA
nlIpXBtwx4HSc4tEu8C+FELQl7hZGWOyZ6VShOtvKjJtPmEWjUir6kyvLG6FpFjtXQAbA5uuNY2+
EpNLmTso+0RvXeS6i5ETBuKDZiir1/7ifZ0L1sX8rxut7sGpR6PkEF66s8X/WDOvUpdCKsN8OaQK
v68fqtRLGecEpZmcMtKRVuesQvpjEaZQVYeLEH/XeziIgUzbrHuobxfc8RWtiSFJ5pDte1zfNgVL
tcLQsxAPqz4s1GaLZjhagDH5oofVLXbXK4f/2PcC0X/qVddmSZiiu2puQ8BosJo1QKLJqnV8KjwL
7o9N1gwU94Mxvyvwsyhv7qPbFczmvCUhYQMwyIiXUTYx5pj4cxA08dm0he0ukRoRHrW+tx5mKN74
0C4yHMeChrNkVdsi313qdGgfVm8esuEmHzgL1oUq2ZEWYo/e13FU8DsFugMggSL3F/SM6+mmWTVQ
4OEJ6ZObXPzYDOx1MZz0hXcRwGPPx8jF14GkW9CqSuXNF4y1sSea46ODKeV5URU9h958aWaV/gYf
xTvbLkkjdeYYPree/DVgeA4sXUfeNRT87URuMvOu/pnunTBencKT/d8HaAHyoGK4tEauAnlcAcix
7xhm9is2n+6ll748LZ1e6D+koEx0iEjdZNmSyVK/I2Mfqqy9qfC2ZB5uEworAEsvzTYWogOsltI8
OZYdE8fmd3tpeHKuURHwQsu7lgguWfCIsvCxi2dFNzqZyejl/XAZu50kkgYyAGkb2zkQT+wf3dsF
lkRLMRR/IC72MYytIJ7TilMFkmXHivxE5qJuNVM2rcaIaAImcaJzJUzhKzL4yai/oQc1JaTnjSf7
qFxVw5YUSxLzqwVhS7MUrKQDLjgbF8Q+BhyuO5jNhgy3uIYqgBNXmSuogke7EhwjJzGRE+0suYyZ
kZtIY4v+p/jVZmE/4DFYKy3oT4VvD6vVoeAm5axshE9LvtcHQcZ+ujL9s5HiniUZpHUsiZagqBfw
0U0Cmztu2m3wABxM9nlO98/p0n4qI1VuZrJbUr+TatsMQy3yz8jx5/2s9P2f+DCAh0CMGszLdkX0
5bWBR44vuTKyqIhl6EsAiBsnSBzE2Y9nEySFRMmYRImpVFz5zIyLoc0Ph8xP98o+eDNw/EIdbslh
AmDDMf9XqOcCk8EEBzIL8U0n7Qxqo/IxgwdU7T3McNIdJfyUUxth345GNMByBmJ0dKWxilwuLLxu
hrfsEknjic9gUSGaJw6AzWzs8ceeURKfsd2Pm/RVk0sl8WrjgqUKAHqjnAIWhZSVN4b1WAbirN2l
BFIosHWniBqHaldMsWSUrbf9EVfyu5QqZL64goe61ByKRdSECEuZzhyHwKs2q+cTX47mHyt3nDue
t3HlHuRkSEK97SLLZsumzF/A0kfjlntUwsOivAIPF+IdlU4VFqRy7gUEK1EifjMjUY2JUZBfBgCl
a4rDiubNzobqJmEhltjf8HfDcw2ZgLz5FdiWmklBcw11J0/gzxUZIuYc5TAlYjqggXHYiW5Bd6T6
0rXMRA4KkCV39xKmQLjjPbG1Yakuupc/IKU5MK4B18fKg0tBwVYxsToIM7fwBV++AjRZqDeYVEzH
l443xkCZOVOFLiZq7lI4DGKRaFoZsdzS+HNF2sAXrgaIbowHbPMKJOEnMyY6xVePZGDYSYWK8vOx
q+0wiRrxVWSxR8S8SWWvwRMQM2o+n9qMmWgbHagLmPevi0i94WLa1Ay666ZFNX38QRzt33SHdZ5u
KogiT6WmDKGPTnzxfFzHwnl2QQgy7xh85/JRZ1KcNTjIxJtAN0Nz1HJURO+Xb/xy8CzY64zoDlgN
fh2bB/BK2i1TPjMUsD6Ya7CFp5QVnRDruNpbapebSjt8dshgWLV8j/7Wfw7oAh0td78z/db6AFhp
e2GaTXAuxw4WEBYMaLTAQlR9FbilFwnuXsm4J0bUSXBaeFPohkNvFkljIZsy5cMqbf8wzkG/iPhH
z3cOOimsCS8aT6SAPsgWw+RF+bMu58l1p2ekRxVzr/yrq/tCDryf0jbpswFERLvoq59bdnRxj1YX
ta1f4wKpsBVCD1cEWh3DEUfKobClLPA3CIr1DCupJ+Muz+vxqt5f5j1uHbOwjSFPp8CQQlI4N4m1
OpxgrTRPtfPNlbnnFIWh5s4m8s3kdbptDUuWJ+BBeMOZWDccF1c8RXmGYqCUomVdq8MPl4uCQgDI
XBovi+5hYpyUbBzcY2rUyfR90EyvL8DcyotWSRK22hvUEZ5FpLDQHQchYs6Zo1LK6rL+s3bBxjtn
mDuN1dbu0lwbtTiUT9dVFWWv6hUqsKczdeEmEJdYUJSCYQF4jF6fsPDEnrb6md/f4UlMAcU5g50c
CW8oKm8QEpxGZKOfpTgbrE2mrPZm5X4/GeoOfAGuPg3ZAeRLcaxtZHjyPXBZYkGMai2nu8QkCxwp
yb6mfNvmGOBWHlTldlR0Yv2LaYFbN1I6WhVteqWcab4xBZEK8n54KqGnEO+r0kJGJaZ5JLqXsCBL
ZzNIRy4PkQC6fyGra3Q4/FGNZ9hdzuOefvz6i0puq9eFshQMciH6Li3AaTTiHX+G50QhxYm4zoUQ
yjyaLbU6S3JOsc6hygYGGKquHxn7Vy96PF0199LTAGYvFEeH/n6DnIe6NjaW7znlB4HuRrEtQ2HB
6ykUEXFAmZQWWndpKjMnZTZPpeIS3r3FmHL+m/J7x7060E8agn9Gn1qYLqz7PaaAW6EC91V/68s9
3k8i9238kPmh45o4xB7ZgyqqMkIWJY5fUqdDZ6BJn0Z1JkGctmK3Ml3RpVkfjyAL4FruIv7Holja
5LwgxxOIfmBX8Nh8NymickZdlziV3IUVndJPThN24ymjyBMVzEJ0LnVsKm5iP+QyNpjEDloqGwM+
2N1q025+eOytIZZBEmva+mwaGcOoUYsHUoAownseeYVK5MX92BJAFNgiG1riK4X2jiC4apGdkPyO
HSeGvKKyVxyO0amYAkDF/KOLLH9d/K4yOHicGHkEhh1QQxdfDEOmH0c0dh2ucW17gDA53byleM8Y
g3v/43Q6ivVEpb3TVQY2U2ZbMflK69QRYOcjR78sZoGtzYCJZ/z/BjyKVUUdeOzlEJmXP7Ikn0B4
Cwga7uGK/Li9hRCrCQ9lxNZmDnoKCd4zxkejbh1iVLDEIWqKpywtlH/rB3VlhvIMunV/gbfC4OeT
NYd2WkEry5/SXkyG2PBhO4Ft2Ei+S212vnzxbUG1VuO76T5cucPfHzOe/SldDwwxaIjljisjlAvf
PNPytED7aljKf3+CnD5+8859165g97gTWoTY+V27gfPiCcCaMXl3h2BINV8Bv0BzO/sj9e0drTbP
oOnVEDQ6U7oJxMMSwy6BfD8dLJaxRxZVmnJbYqs87lwIudUEeacF1byrHf6XpvudDN4sdT3Q8Jz6
D3ycygYov515IL1pgO/sm3vZBp68sq5RZdzsKXQf7c1EVrTEKPL5/6eoH1IkF3/h96/P2XKDOQwE
jgji7YE1likWfjXjjO/T8sLrV0QSSH4Rm0ABe1m7ZxMfgxmofd9Zh+yQz/jFJGJQY8ggl4MhAhIV
ISHYdKfY59euALbh2/2jGyZi/IskbqIbs8F5bp852luNCgpXWYj6CngeGSroVEmCX/V7DJSmt1BK
azdj2myYfv9k6qoa/FgxTNtTjZSMNPAyNIQQB3RwR/59xi3QSx8OkHKQa97jCpKzWeehMEQo0sr3
PWcqbOjH+RwtDDhNk1dL5gt5xnxM6a+AhsJfmLSr3yWeV8IfEjHXDsEFq/zCD25JhYwVh9cUkmHc
kpCCR/RuBKODUeieFL23W8BK+lKvlLIiKSV2HC7E7m7v7UxFGrmQ1acQMeYl+8i3I0AzwKrsW1PT
/k8KrA3sUiJ59zlrr8339qeGw6LYkNgdAL7CuzlCVoYAEzq17hsAsdShM0VjDuJ/lAHje3YgHBKR
rLC8eXJ+cBCpuGSGw19G79+Wrq6/LPJaQkFyNCqZkiL3d8rTcPsz95pQIwexdILPRNPSAw7Myj0/
LS5YjKwVy+q+kWLxs92Ilg33SicnwIDSs/c0hiLHgQ66cMAZWzs5h5qi1P7xm1eTXDJxEPNiz2Au
k0VPG0NzHIB/pBDnpZitpf8kusnGp3TxUU2QmhJHj6Evjthd/DNxgZp/pu2pe3jReFrQguUjYrkE
ZF5PODwoc7HUJXp8RPYucRrCHvQlYs60iwMvwjTOw1JEfRLoREgIy7oBAw9ePjX0H7vD03nQIFRK
x/cxRFfNJr3apsa9NW4nknTqWGe7rUyYlxF7crpgoaWD2iLaJjSb3Bgd3DnrW7lIC6K0Y878l5s/
Vq3lpjU2hGkhTu5QjpFAovIR+RCyPZOroSDPIm2XCQiLlvWQF2174wglMzJiS48Pt4tBJqwK5yJ6
WLSA5q4ZL5HW6hdFlKQkp0sqJWxjmgtD12PD4aRGaPGjK0ObdXhIMmDbVYJHe/Z/Xd0K0U1qvn2e
YK2cEVQcZYFAmBNl9TeKhHey/5Qh+5iUjQoTki+VNN3KrJ0wldpsUwXBWKUiQlxVMvW7Gut8W7xi
OTmccmlyVgu7wWG9RUCoLuN/gwLoaEp2XoUyQza0YL7B/hjMPAp6+wo5WbffwI1bvBbHSJ1PqbIV
OduMTghkqmgWrrz8q7ZycFQgjQ1bnunvaTNtvSTBOi0rkftDmT9LopywP1cUx+DKHkZr8F95Onbt
/e67w9rVj3/I/j8BNxAPhZPNiRWm4B3NkbBndDewV1VHn2WIS9WvsFPLtkj6qEyjSzkZyc+Ri4dz
2QMCZN0+/SbEWMxBgt/lRcJ5wytTi9VfZjoZSspOIiIMWCwba9FCJUaMmrFjfL92CeWGBOaLfoae
1ZHl00rkxhmnTHq/C4myZCTZ1vKOLGjw4IM1aDAeX043fXmx/480DsP3wmKlQdbVN+t9EBWAiiU7
mVgjT1CqwUz6cUlJcx0pcjXLWOffFTHHgLoxdbDBFQHiyNFOuCMMKSqTj3GWGKNnBpsz0KCQnrr/
nXK2+6nhWvv4smOxjPOrU13uJZVHSBdCvidS6OXhKm9mAFAgvcRW0P2X1WruBlrG6WuWx8CCsJ71
XrQCCd0dIjPl2NlDxI2nOXFcDImj9IedwT58/CDRbmiJNQcPjnE57W3CEeQL5FfZu49jf315yQ84
kST03q8YOVY2YPt2lvu/D0i3BsIG4MHQySPTh+Q7nRaBwptYyh+abIEyVyKx1mli8Ie2h1wMDWF3
/OETboPZXABPnUZMfOVDIibMhuL/20fzF1EPLlM5QF/8GMAtq6YVTbXPJNkcpJ4xZulaJAbLejev
23k9uH9ZThneyqn0wUXJV6On/i5+QaICCvIL7Y9iiHrxGCiPnPYXt71DXCAbCQqWKZv399Xc0FuS
U6HI3lGbbLGUadb9QtK47leQDTOQ34S2iSjyzQeQlQHGEWq2dgTb5NY+rrDTWAavjjkJ+RWEfJed
47utAReuy6i2KMQ8K3HHspgyHC8/Fz7SGcFN0xSoyP92F1eqQWjoaYt9uD6RiZ1NBGfoiKzqv0Wq
gwt4n+Ms/m8a5PFB3OBcjuYHseJKvoi2XSoaU9dqaM/9VRJt6UkEs9Z54xLVBHfjSmqhxKu6WETZ
QZcrdpbrGxc1hba8mAMdZISybqhQv120z15VYI0HK2Bm4xPJXJ0EHzXnMULgetSiZCMJmYLXE/KN
3f1NV9Jz0T37kQWJN224MCT7Mr4daQod5yhKJ+EzPdLuzgklyTnXfGqgiVMSf2F7ePjKGG+iQBfS
efZxfDetc76H50K8y6R8IjxeAlhjUsODAGkzyIgstE0g37KmDkVM+XTnCh2mwUa5nz3OF+rWRUs2
umYeDJUGeo93WdWraR3d/tP9QpcAxUeCC2eaOB5gkiLqIQqaUCJWjeWr2CRo5PXrIOefGnjj/eS9
Nuc21PZfKiiejifLXtEfU7KRBOQ+7Ely6jnLX/LRQGZFJrjnCUxGyxwWTol8Hf6rNEn8IFn3Dapn
2XfgelBMH/gxXHyiVCHPLuVZcarjJm7ZEYoGm6GTgtgBEpEnNITGA251F47y7vHjAsraLbHI8CxG
16gWKAQar8JtIEKS9LXjLU6LNGntk8WAqv9nfuiT58C/zcM5+XwqppzqttayUqN7jk1spHgcgwSv
jBOP/WAH2nr+fLFRA5wNp7ZCYmsUqOAEYlU52SXO1fGE2QVhTEEWbnHonLX1ViaVjolTwevYMC4Z
lQ4rjNj51usD5L45tD+cPzRpKhiSvZ3m4nQE7E2yxddI2zHRoSQjHT7y7mqdJIgdG4DqltHSeYln
DGvn353+JEqE/umBM1gmXTWi5i15IqKjRDoGI7G13sm6BYFxv+QcTflI+U1enmwNq0+5tHQt7efB
vmGDh1V1bHw6LW+eorVL8Gi3xfP9cvJYCVed1ZIX53eWQzu8k1OjyBgR8W+sicRi/ErWP7S59unz
LTGKdifAqk3gNNaDvbL19iT5974teP0ys1XVMvUZkWbLRViz9qagoowBC3FMa8CdvTLYcXbG7+3o
UdC3zI+UZ2CpuQrhZP+WXZxve/koK1mAOR/iB7InYVt5IumVlyTd+zGdprBc0Yjwr91ciDw5fWtF
GsictI4/acttoBxqLVgLQHywB6fpyA6NAB+A25+cmDWVflllcKIWgLsLVxk/LpDVu4zpSlL7BPh4
k98rdbI09EOxs8qgSubUszXcotR2jmW3RdlxiQsw8A7R4Subg4hDdyvBlkfVLF7vC6vRjmRCyW3W
myX2IPdg9IYl6fKZixk2tZlyx4jobsjP8dbGEkCDMIyAtDWw+mAF81Vf6f2UeSobpLdGhtwad2Cw
jgDyY1jm5huQXtskKZZnVt/s61qKFKIv9l5Nnur/rslhgQylEoj+mILqBM4PIl3Bv/6VJSGIOzm4
nj1P3NCVX6QwnRk7nkpSwPZDZeuoFYM6H4IHR2dQlBikv9DMMhV4Tv9G7bmqOEoa3EQFBNPjodqD
7k9Ue2/iskymaSZf8gyYhR/9z2D3+1yAHUv9yHpweN0VoBDjzwXvNLMOHK5kZmpqPj6HingWj0EV
qpXFFv+mgU0czDE6vcRrjTyeN9Xsv8vx2kgOY1Pi+e8Yi+a6Krc6oCQHphkaS7baQSwTZYNK4aw2
gy6AY1dVN3a3GTXrIz/VPwvKsWr22FZprv6cIXzkVnIcPAUaaboU3FCgn3s7lkDCuY47bMPNVU3Z
DahZgZz0BriWEQymazFxiabhieA1OFTNbpZ5En00CR6DxD86oA/WmrcXrxWPwg64hDD09mwNN1Er
XMmqE3Q8WzA8fvJjUfYiTy2mmZjOq1E3z1eNk+A6+SAq32nXjZN/cVn9v0ySo1D1DTlOzHN2DfOD
0tusGoQfL6ZM09v4V9FHzspeZ7825w/yNeGRnOP2OU/JqF30dHUIogzrgDz1HbKD7BuH6chRL7Lu
S9QhGgehD83RSXxtDWH5RcwiRXJkicHqfvzD6YrWoY4gzPWjH9rQIacbFj8K50W77dYbBcYSRwol
nqQdn0Q5Jn8IlcIxfZ5q1W+AmFSX5jv0CkSUwL8ytI+QGoX92B0AMpbQRm5RPkIIxwLVW+2/6x9K
kwGpUaGkJAGb3ortY6L7Np/6F2adH/nSZcDVfD2IJZXjz+ZUCnu1GClRO8WLfbPt27PoaBPCT+rF
/X0NJUbpbxiBgQetzoZyzxmrwO4z/8EBmglRYvgS40KiPJgauWi5AKmesKjLMa0QbsKCksWi2QX4
xHkHUeLGucBu4kvAITjCSb5dbi7S1wa+93J8Bf9BjefhYs+xUfk7zbDA4BBa0Hl0til2N9M8Evnk
BEgg60wTf6zsKEGEqr/hAYAguSjb7Xok/jNp2nKpL2phGlfCFuCJF5E3IkHEyVrjsvgvK6K7k6VO
Al/Y2l0xpQv021qI6G6g+wWYO4zeTXP6WieJyGFfu60myixoow/24q6w1uNzwh70YsiMXYvjNA0p
vdEPhg+ZV3CSvIP2KwyJ1SYHqrlnifgQkw9xNPAJpX50qlBQ3+I8dwYX7dVfcagtxnr94G2b/8ku
t6OSK/Aa5sSmh6TO4Opy5QLpyP0HBJxzTLgMrDTuHTlqI6V3wzgwfRFsYn4IVZTLGUA4zNYm6JFb
pZTRUJsoe8vv+4juwUdv4+rO5h9X5Q52a97PG26VGOJfe5yqlCwCzqbYj+/TSIjLayvA63k8twx6
IANEg0El0hftxEhHF6XnViLI0a64gydZjW23U0NbY4/ovKTKQiZeloEZp7A+d7L7nwi3bPmcEOm3
OUnn2QNyaoDGJazNvan9HPnxpocRixm7xuStXPHodJiZZ4N8QBpfbLoVa0qU6Cu9lISYDunoqs/a
Nwxi1/L2Gzeoq9DiUYxJiQQKbqkgkTnuPtXvC7VLfmptTm9TlVHCz2RCE9uZHbK9bkVa+ih8yI1c
IM0JY7Jrs0RcgFGrwmjBTGnkldkkLTJuKml44BLB3Az+jxox0ZhRY+sMr1L7Dv9jVT4/ttMQ/p1D
x2J3/4I4ztQ/B9snNpOhlDPRJmbXzvCYEHXbPDEm0Y5opDwmAbPINYUtE7whQ1XGVKgkdjQHnGqI
GRs/uS17v5oKp2JWF4Jd3aXMUFERuXhTNN8RHmKf3BOfzffDcM/BOBL89dZ74zG86vRzd+z0eNYk
SHB7hXYVfTXgW0fm6IMdc5onjfOUlprAsXk6M/S5ylAuG/kMWBpvjP6m0qm9SlVtCpZM1o/ccWcd
ny5yLAv+7JMkzjyAsp7ujo2tJ/j+kxgf1WopqDZoTirkpwuMynpa46Ka+Liiv3z5maNpE0VusGJ+
vi6RCLL4h1g4gt4SMxFGDotHM/m4gCM0j5WbdGk8U0TmxPobAtvi1j6gUFLmYQ4EdmbVPTcVGskF
b0KeIJYdyaV3CdzcqT1RiN3LuPsV5nieXNCVJwM7NC8rku5Zphb4TR+xvzG+lmZQv4TQ+EXZIXii
Av5yGnQFifRR8Isd0YxEGYrEdVaKLJwEG7eL9NaCRHFvhhEBP6vpSoaGD/IdNxYLgKviL9UXOUk4
wzawcEHuLs6Hu7uuDBhD05HrVs4jruevFhzBaKxWT+/0ptw4mx4fqif/tXhZWJ/OPC6XzoF0+h8f
4D7BZKbw27/H/g00Hn2ptRMNfmrfRpnSshuyX1DO+oECRzGDMA2gzDgPePEo/9T/Pv24U4+yPcn2
PJ8KNolxepDtSuBhG107QlvoGYyL4nhlwdF4Dkk2Wjb4KP1WcxLOb5dxcRIopVsRbgHlK+qLQpEr
QC2/f2kLN226nBpN+XOTFigyRld/1QnbM3M3qr+P5zF+OfYDAC7t54MVVy5lpYAZGpMslxRyezj9
QlLnrr4RBSP5gozlEl4BEcGp3xAsH0vJWbDpBB+C9+3NAhfezuBR7+p0uEeBDgJwgq3Hqy/TtmI0
88ZuB1+Zj/7NtVvWYZF71MiMiiSZVBl+Bx57g494zHhSuEJxvcuRglcgAuEOD5MUeBaQvFcAMmm2
9B+aXxn8Ivl6qDI6SCSDUO2hXRVoZ1EJD1ihdVxScrnfC0YDuhtl/nWydY3mvsd30t3cXXd+2x4J
qwOuH3K6i1F61tGMUtLsFxsx96p+Hg0ZNb8K6CPZxTVpUGLjCy9a/kezvHYmMukGuqQOvmh7Xy70
KdSNLNnjEklqfurpp+iIsP8bb198q5pIy3hxqq4Ten6+C9xCd6W1qq72CF6P74SfUljSNc8Fv/kl
lIrvliizjnXaI6aqz7d6A6w9fTl7szFmx0fp4d3DRRIr5945qdm5UT9wBoPHzx0G8W7mYfr039tj
VZsV6idr+XTLTwo1WoJHDbZMYDLWV1W9xc1zlcvJ+6wITDVNmG7j83zicCg5QYxk3llZEVx+6LIt
Ff/qx7+4HHKQVruaaNrLVTlzNkX4UQpu+F/vWsKiuBGKSmsuKgBAZGeRtrR19/NeT5S3ktXxgqQJ
mJNeizRZHFo2bXjupRSapojT9k24ozdjfYfy9XghFlgvTqtsYrx/6o0/7nV1RyvW3AGoRDFTZduk
+RasMZyjp1GDDR34+NDNzqUojySg8JTLUfirfJrEAXYqbJRSC5+ypMJHnmPGnDg0a8oOkEg3cRSl
XFs2vpRBlXWoDbStHz48PX4U7vjWDobSfwqeZuF1+sCw5UqdDTpZNjI86Kga2LdCIIPo/P4UUlZZ
mAlTMgsm7g2O7pZ2xwM1ccPtOsNyR9BwTvnf4VQ55ve8oVmVJxp6Bl5sCo3o2MQgZMSJSgy/0nyG
hkIgiPxITsJh4pnL+OsghL0vtoTJC8tAdq58k48o7WYSyPRS0YGsfTd2ats2lXarudP/DErqWLs1
8Gm09r/lGTn97zb5tfU2ic5O2ZR9sR1+1M49xhB4w3V1WSiiCAIi5rVqec2lf/SjwgrHUTtDL6P3
PDT+Ann+epONG254epqFxBMUenGnD85e7/leI/cyFFs9TLSRqTdjyrSb0bKa0uKWtmObBhtUFZ6u
nj8m2f7/Br2oljhVJDThYP+sATwQ92ZQCakrtOBTcG1KmDip89x19v2u3EvfUwNAgz3VAOTfxCOi
u3VHORXaBjNliXW4XfZCKxUUVHmEJrb6Zr0GQNbixSnjxiRvqqIoQYDt2a9T/TyVKL3DFEp2wr7i
TJcQG3cMHXZkKCC2hfZINLsKW/7P6V8WMcfSQZ5M3aY11L09eXBNVNu30s1P1YpCv7xEXeZptIdX
4YjjwUqm9MHPA4DWaM+eLtzUjJV3BDbREgNrvZAGFUDR4jpX7E+IXOIDmSbZZIuDLFkSRhWVzGzF
U8BXSKZGMWN/7TZyY2nvdeTELpvn1u/yjt9kUFcVCPcwZruIHAYJfwyREVg2xxxPcL4o5WM6h5Tp
KZQEIr7VcbSi2hCiwKlEXaUJOvih/SyyYnnJQjuIuMkVlQy6dXnitdVRAZ7hj//1MUsHZ5AMpSGw
avX0ylkynI4p9Mbd8tPPfMwB+zgJlfcpmHF+ltnGk9ZIJ5DQ8aPaLkpsOBLn+cqlbqfDp4paZIAH
yhmhpfONzIqO/PFATU5IvKJV7Obi6kH3NL3hNPdKNiOjhgH8aNAXKjF9oaARiZaRGgZNWvPHvMJ6
7Dt0/Y4YWEnkAO905S6MQPfSu7/6yUM4YsindIW/xdp97nCmsoWmiR2AXMYbXgWnjzoMosBwhLVW
p2bevXv9UHOvjFbsrePEJMFf33QSk+X9evhZywn0gN4wkZENYWTiZ/93FNtj6cyAmlsJxyqIaXaE
vKSwFHuroZnS4B4udKQgqt8Z+JDpYcXGk0cmgAx9vDdZjmNE1fcEhQjxGTJM5wBmLWFEWKv1lMZk
LL/9Om/0wSHbQoMnuwJ1flyA2EVkviOX+etmZ29XvzsM5CAv29aqFRYEFOF3mo+JP7nAAxn8dLog
ROnX6LTFiCwEcywXMvqw8uWLeJ2Dy2jI2MR5DqXlOBx94Ua0Jy64By5HyWbq0gp5N/Hy1h2UjCBg
QJrloVeM/OjzndPMskAZoIYmS+SHQuRDL9aoCwUBe1aFq1yRtuSh3cnH437AbAsb8Tts6R+bjgAs
KrOfkIBkE6O/Vdei5abGCoGZJ4oHtQuTTt7rQVIQsXuPvVb9ocdG2VVQX5F9zE9C/zjOS3InngmB
hpatw67cCkdWmJ5pKxa1e1iXlAnb7tv3VztzdzNTht6xGkgYWNX2bhU96wk1d6nrlF47ZMU5FoAY
KvIlYNvJAyM/NWpvM6qViycoC1AmYU7M8lP9GHTTgJjzqxJCkw0ypK4aDTH9+Sh22qxuKWSuwYbe
HcCB0nMpcW0yUJoEECi7h8z45lKMj8BAWA08DIq3DUCZ/A3+q6ql7QQpioOIMlgAzixsteFH0/f8
4ukZA26JRmqNhcWOqfQ/jXH46B1GkofqOVB3dKz8IS/0g76js6lsPThiLfW4XwOrqU1BF0KhhmMR
mLKomyuCZPbJexMmVBLDCoFVJSHzw/ZGgWiGIngGmZZscy3oq+OQA4XXjS+V6SMWP7T3wR8o83in
D9gU7AZl7J33Ib06kyb+i7EE5r4R8+RONX/VTbeMK2+qTlEPa6dBxZ99poER22Y19BRlAK4iR8Cb
jwVwyRHsN+LqhCHdBZB4Ir0kv78Sof4e7zm+pxTAUZlRJV63GLUJmTxWaHH4mQ+EFomv5xS5sNbB
VKsFoGei4beJnnEHSCOL+S2xJsyNijBxb+7VUzwjS7vs8xjhovI4i+IBov35+wpuoEOnxn7mD2Vu
6qNmh/8mMRXtfz44Jn3C9bny9NI3Fsq/P+MOQa1TVQV7SP41FsOzKIG01OiKfsC1oChyLvVKWSrA
ht3oQRPrezxRuy92CVxNcqeGZSTrJXQFzyTiV6nQkGmUqtvk3+Ae+Gw2odThY8XH7Q8SUrv5z+H5
+ob2dtb367pr2ARjGJIcZq5JDsYWZ35McZDi3cRFm9wWUuyouodIUxNQJKkFKfqh1GAw/1XTN+zc
jn3skpGFbx+eCe+mySk3IhidghN3grREI4MM/i8qGkNvcI1WUloc1+HCZKmEChpuf+5gnDwJ4bbe
BO/iVpihUA29mDS9J7KOGd3y6YcPCYGLBjNzubzVxiPR4d4yUjhatbvr9V3FsjGPq8aK+gKpcsr4
A3ySA6mv5W24QMd8boD/Ah8Z4/w8MdBlPCsS0+6kMYfuW5VELRYbrcDgaw3rklu2c8KtBi/f9FQw
VorElccgL3IKmDXMm6v05yBIL8lQMxnKFYJlp4c6a1ylnjoUfWzuh/niaqFSW2P9wvk4X9QneVTr
uzdhYjtS/AsnTPfLrxIgGEd8B+YBZT1CpLrMf/s6xrVO4TNaP2Hl568nENkDH/n8vKTvFmC/6OOH
Kf59rh5ioXpBYU3dJrlTMgMK+1CwrrIDMQJ4gbSxVqVogQHNk3bytuMMP4VqaIjteH6l9mJY1pAI
A6r0zkjKpsC412x02LySTGmE+T2XjcTP9sNknTa9D601i5WkqlfggDJj+u4/egkubCGEViwIueC3
TJXebsRtntUWwK4wdcNqPRgKcVrIxAfoGOdBifkNXdNxZVgwwelqnIwj33dinSeP/W/uncQr+7oj
0k5prfdR3p78hJ65XPDVO87Rgi4vEmEpdUvuuvpYbDbEEuon4KSAKAe6/ALPaO/TcBd617ZAgrUp
aopiWd76ppoG5Gs5fjKK2BrJ+vMconj1Zph2fG73GIwjv/ClP2KyUwHr4jKPRwnQ5fTUAl3umEBd
wSXsdAIqsbyvYZt/BTZuZ37evFJ9mCnk5IiRjZkNSSd2yEom8/Xcb+iwxlgTiLHkc8NyaQQYUJ7Q
Dv6nCNxQs/6Rho3vcShwafjwS5FmdkHOdw1pQwKARugH5wiBDOChAtdXDMRMO9zD5Je0vmp9quSc
v3UjZOUqcILeLZ6S2bIV94e0BMrcvMA3n9DiUYiRyopc8B7Z1bjS4vwUv9WOEMUhUhnFm2kAuMJZ
UGTRndK+iNrcFzfETKgbxKH3C581EM3M+hdC8hrKbu2Mds7FLsg7f6VuGaHPoslRPvavbMycgi3q
JT/smzAZkoHUU/abqCODhVmbDoMfg7olyQhNd7gJPgelajflzz8IFvKWBjvelKM2zQcOY0YiBdgv
72zHBVgXEO1zkPjs5JvuiTxNLaXDEfoHKmJ03ax7EQ5W0xsklAFgp/s8SzbsbvmDlb0CnT7XBwOV
YoTf8lzaONrzkbTy/LApGWF5Mm23zKMhg4WEupozMqXtQ33o6kaaGdFlOGQu7rouRBbddcO8PMYF
HHKbhKKASSG2ce5nQe8DuoEojsWLoY1HfkxKIS9baGLTCHygfaXMwa2V1AeWTSy/CBd5x6IAKTzf
aWmJh/j3ZrKtFCyret7ksFbyaqAKs65XOeIk14xYeY9nbSMfnvKh4HshWInuxG6rVFvrMuM8YQGf
/VIQtA6rYe7OkJxlwkb22hHrwIIjint6V8N7cUvmBH29HTePbmn0rQHoIKyNTw7Bbuwh/sRqMjjm
iW11191L+EjiU6oVWOszzaYQj0dkM0KIH+habjN/Ie8HSzQ2roojhouOtpl8PkUkANbr5ZqKoM3i
vApKH8DwxgfkjnpyElWBouVROVNHpx8GIef4Ee20Ls1E60W4aWNGYDy41dbWQO95DH3CtvWQ1kTK
0F2kzjW47sJ95MtZifz2JC/AtsN3i5JCSGAdEMhHUWZXTPpzA2dEcLy2o8A9xF4ombwKAqrWj2Fu
SAqAdDMbvjqxE4GSQV3uvMK1i01h4/olYZdWrFfKZG1S/9Suj0mV5/g2xyKOZBC47uw0TTshuqd+
4IThDomVS/2fU5CdRQu2jlrdsBxTPHNuyAJd9LSXQCm1u8c8naoSU5eEjMt9BwvoupTanXeMJRQD
IqDdZg88miqgvxAtZGdht/Ofm7CFF6Ih+q686THHiCBYEqouw+obChb/cDazWVR01NRmqTF1FH5B
tYKwdwnlkNQydT+oWOKHBfRMRG706H7UNEV2OacGEdBuLwfU/YY4NCBeZCO4QSGeA/sWD20yu6YZ
T2rN5/Mij/IxNS2dULqouuI3IEdn6rRPSB/4rsMOE7GpF3v6qCXmOD6dVYuHb9i2KU7YFNINdm+B
gzH7CNVXq2W0flZRnq5BFpZNIsnU+dWkx7LgDu7IB5nB7lb2+1bjxhq21pWHfBTyDIN2upmbWRz1
6tvyuEPb1rv5UifCnpuK8kX+DiukYsiMXBfBoACsIhV/5S8z7/OqnquLRGNg86sSA7smshRD/BsC
6LaAdXZFny8OJYRXRmGpndmsxNoSqBcvxE8GQT/bKHOQJwNLQRZwGRr8dMhxEO2YLvIm9IAJSQkL
HGe96No5tRsyLLsTLSp7e7xohmv+Ka8g85bbaAMLRrHJHIC6nPgS7oY8lin3kLkuAWjDLZQvihJQ
FJDE7+L+dgrgNxzdyG+J++haPOgAZ2cc1AoFxf7Ln1AEVxD92k++4S4iQRkFiX4Fc3qd6CFdG1kF
kPKJuxv1j5NxfJ0ttDlDM9A3aLWNuTD3xjzpCNarYytBYMDtr/gMh2l2FbQ6fgwrguC45zpMPPg9
tsJKEg+6FO63OwA4yveWKDGPJUwdB4VBgdSYUoRbXmZZYY7vcnASQs+uk7oAu1H7GOh2eEv4LGev
JVWOUZuI7QEIhsOlTNxtAP3+GTcvboiROaYONzhwS5fz+M7BeCN3KzcCWi8lBI03hC1f0EKnRpNs
KWT8N9ZqgtjO4wpZumGXzE/GqJapFDCcSQnPiJ2ENKoKb/HePnlwPFZIZLAWAOOUfHe/FiMR1JPr
5+blRY5zidz1NbKxHnM7Ick8MbqLkDQ2Hn0AS2T+HXlxDgivfbwAW4/UCrTYl1fEu1k8hk3QfgQ6
41roYl1NyBIxw6JnkycDjwybw9rLVm6qNcO1UxH9m960jAt95Omr32/Zs2XEDfum2n/YmI3ne1g/
1ROEoS8ucJbkjpnlmI5lCjQxTu3vp6J2j/ysRwJOm+hzAcstK6myV7JTzivcxl+hEc9VC3DK/A4x
tc3aIZZg1uB//z1wLDYzotcBfEBAfoFyyMEuBHYDI0mxPPfz7l7pQCVnmUDQ564bw1Bc7Neut6Ax
cFST/m1a8hHzYomHTGmn/hmW5uFexCYAEPjW4aju6Xp91ZFHRcUbrZY7AOMDKIGbmnJnVtWNnUO/
3Qzj0bsUfQdfx+ieggkoVcEKAJLSpCz9vNaErdjQZrvBuNkEKowjC68p8S4e1OmwHnsjsh+6g3v+
rlo0GmTSw64kEu12vk6KKMrAFE2FWr4YJOGfO8M+UTCvtpp+GlN+s4MPtYw0ERqrFvIMMT+MN4ut
anJL8X52dW8CO/SSpY5aTewoP/WIEnV39UvmXfKgvmunvoNfeMgfaN7KFXuW0P55r7aEGY6mKllp
+XpsT4dftyWZEvCSSb6tODeLtxMBq4oA2Zjx99r5panuMuPKqX9GzIukhEnd/iOBbOhV4PYDzpM+
gwwBSePCwlxAWyAvmYpAeR+mTcwt32MkXKR85wsG/r++EEI7MfAM8zLnlttrq0BkmrAoa+ttM4M9
WToIA9vTlE8byhhlbTeHQQPg/+Rryeic/+ggNGkak8FQsvfL4s3sEkmdAcJnxNbAOmlNFFVgtV4q
UsqLimXjhvWJI7zJ2mCXs3YnyVGRYxzXLAcGfZ/PnPL1H13uioOU+F6aT6dPLiBHjGuhpJfVEMgE
Klsrj16HSo6HIRSL2DTP6hpzWgq4N0fnCipZdIWe262ndRbgWpQ5xy45D7EFPlh1FsVgj7uuWmRe
YqK6//306g5JR0/6HmfcRly3GiBgopdeewFKhIYRPd5AZjVNCIJ7KoYgNfPTudAqMlejZIUHQOOz
16TJqLhUQojzqb0STs0BBZHTR5c7exWhFBZRV+nr1Z8u5Bjwr4OxEzD955Ok3Mi/n1BSBpJRPsmt
XXDVRUMMOYYQAYypNiZ0q3LHMpy5GGwOeSTmGkyl7tJpGy3RuYk13EBfuZm+MYU1uRe+2wY06owV
FTqG+DPrT4HT9ibPwRsOeSGv8yDqfPYEK3dVbIasGf4AsPva6t6vQnPGF7Ob/xYAeGz5QmGsEC3q
d3v1n+0xIPWzxyR71f6Dy2j5HeIQ/sRjqd/G1KrXq2omuAObBTUt4Yc4KbAEajpR9KTEajlbIE4q
9V/aONsEV1Go8+X5kvVK0dYhhod2ytNcOgq0V/Wo+sfvf9CUr95xrIx5lGGMymTO2+83n3Mldnzt
rMlWgGpp1l7bLAWCHRYWCzxNoSyNhETSZyFE2xs1jPx+DHMI+KAUd8JNYSphomzPDlLK5+FSvCyR
2vU7x55PP+QNNG8UmwcVkkdkqpL5irTuYx3I4LN3f96rFLJCRuR6IwByKDRhWxUNWuFlNhaTHBAC
9A2h5BaHX7Mo6gfrkRcCLIrgOwF1N9VZVb+km4v7pzKYslgFOV7HV6w5+Q2MwbNxic5JnUXdEmcr
BPivjH7DYhJNJb/ZGiX9X9UOqr85KlQote1o0xplvSTlvA0ykwLDAxBAX9NUFFyBl14wLjlqomhh
qhyImCfQvbbmpyJ6/JnjPh4V4mbp6owHUJteEvZJm+kB8kth31sYgzLg85WZKqlu2tk5T/vsZLPy
RRXNe89U0efHlzDHSLBDsQPrBgR/8Z2rWyAnZ7Xl4Rcx2MdDhgNL975Vt/L0j7WLc6HgVxM+i0Hg
nKjMDAYdaGYdvGBCqvYuDuisUhpb92VO/SpUC8Ne1R1tU29YXxxRgT7lxan7vQcuN1LUo5zS81Yb
e3+AwVQwWR3Ylj4LwUP4j7t3mpd+0Qbx19P1oPjPdOOG81SNyH4XsxbInSybTZ2tHuu4ctvMI4oO
cUhTznOnxhiCpgfUdaqpgs28kewZU2DICHHASLbEzSy+LFGxquEbNVXbdgdmTGOnAJ2fHSaWWFWQ
0zb8ZswwANmlTXzpTrh9iVteEhiRZ44tmXADVht+3KzFffneEKkIFvJ42M+4826vCYxTS3El5vo8
O9nRG+jLlivT0+OXf1YxPgbUfsErS9+B0WlBxlerCfAk5CgxNjG0L5isFuPty5zHqr/bYmSFOSAh
EDjKabLoESadj/Wh4tWg4/58QGVUU3fziZSwNY9wO3hMNJukNjHcq6CKRNXeSFetx93H8A6PP/9E
MY+8iecLtiikkNU4SqRnHhWMPudflDJ7kJLuIq+B+FbN3l+tSiSccZRsfmpR2s3wUIRFLDpxEU9z
yW5FnEKNqXWRPr1w0AV/Vcg+fyBRA7jOMNkNVv4slQzFVbTGSuU4Ytb/N2dy70iradESzs5tkRAc
Tsydd2ASZ4MIXY/HXqZODgcEgG9oVq1dF8cymV34oihdc27W9RD1ZyM7vo5wXlRZjW39knEX1ZqU
ZV8cLC1i5a6SVlLU4DJidCmA4Lme4+MRHu4uaeqIqqUIbbyqfu5OPHa8sFFyrY9o2RCfJSZWr0cB
uEEeM8Y7lHit6CFi8jZJtoEE4/m01lFsPHdng7dhln5/J9/fxlb+FicRoZXJBtjDrxBq/3Jic7AQ
OAvHvKXX8XtpkKCsODqB5zuwVeStDQ4yKUvWsRIXbXkGsMFvi/RfFCrkdm3CJA05QopK9QQBQjGm
NpX74b+Qvmy5p5Aq5mO29Q98Vdo48/xvSsQOKrMxayi1zziAAgmeQQmu9LbYxzlpvzA6uZaNapyH
osp3W4xFAKi2tfsNQFqrvY+8HRRGpTx2lhSJ5+ikgD/Y224hh1pnpRQOS1gkDuhjGq2r9SZbBnzs
GGGvB+oJJPZCUpLd4T4Zc8tos+LCnJtdCvWWskE/Cn+KEOHBXDAOeEtnKIWY1odztRLt/Kg/KdA4
6SY2JvkFTdZz7htb8eV/bAJL/va7ZBEn11KA0oOQXikIlf7slKy/o/EzA1DUf5jXBLJqrQFG1zLD
Iyai85b5u1ldLJZDANxx+z+dgQ4SJzxnV92Zo8OE7ZA2tg/FDVZUAmrg6SojEK5Te2LNy/1E0/P/
/OWmI0qypfp1uR3I3Rj+9lt1zVPG3DLVplh8n0iJSFoUBv/Dh3TRU+sWVOI6mH3NEsOsEoINQW3H
55msR0j3yESsw4v9K1KMEjizhDNibqQcURpC/+yhyKD9rCTDL9aQjJlGyia7VD+A8lqxcY1kNSIh
xEmrmKwz7tCx4nZi/+MHg9AxUGX8Lz4DyRA6qIlrhiFyLHSLtAko40TxLIIfovErfXA7Je7cgZAr
N+Ua3QxLMQAyIxYii7qckEM+NoXY92VMYyXrbkeX2pvkcVyqnz+ZfpDVszc9KlB40X3udUMohFvO
+4cGhsGTyd8hqgoyQrMhVxnPQX0mjFn9aBtcy60a1NyO3mDSjEsrwU/wOSGUQZaLJFgKnjuvFsUE
tNEdzRIBbPgVQ/bhP7jALlHHTuXRPGrCA+5spAotWA6XAJylYlFf7Uti1xsmMl+KxUxjf0mZyqIA
V7XPhDHzf2+5O8MyFc96w7sCm+AM3WgwtGi+/7t9ZvFg7HkUmTO97lWHLuC4uUNTBooThTZe93Sc
QiL2Rw4NUbM3Kh1ceqrcVgLuOyF/oKaF0reVeWAA3XJUwTp5vzznEQEbyTQsM9dLBT6HQbb5+Rgn
/DKmNC9uE4szvLHn/MCXoeab3ki0A3jHJkdLrBu6TGaf8ZlFdjMoEWhQE72ehwIjuXgU+ndeY142
6tXLhswBNQhqf7pWvRkbTIg7Lz2+/TptZJO7KI2jB/L8yIyf4lnONwnsfN7/Ijm7VDwDBHi1Y2P2
85BF5PkZ+CMSmfwre5v3bvHwu39pqoM+ahSh7n39s5qSsqACw9NAIwOH+rHr+6LajB/HCqJQwC2V
53ufEfz3m8A0yVQGpWWHOUc9OLDxCjK7GWYVuAUEnXEMd+iHAo9uBrv1r/LDExIAqxCJXE3DnufF
MOz6pcWcs+o9V2W4nhr9NChNHE02UejzFXRZ2kBX/v1/6rKJOlirBGkFT2+Ma5kMp4LXaJMBiKBU
cbWXTjoTYvIjWD30kO53kN8kIG6Se74MYw0yaIu6eurd8JCkWmPfXS54tDcnytTSWzTJgXDCa+qH
3D/XAKSTBNgBmHFCFyxvybqtmuEVmvSG7iflpKb9GrWNgPcz0obqBF/Lli949s1pSyBA21XCg9eh
+PgVSiL+s8+bsewiCkrUJcTuF/IaYlk9WBTVkTIQNAe8mjvc8wQlNuJTqRU4Kbe++p+sLSCPfK5g
it3bfdUUZG1987Lj2FDeR/VPJpA17mMtUDWOwLVUUFrFeT5n9V8d53AQUTtulSeToczgNvHLcekx
NcHGzfXzyZ8jT7Zrg3RW1A2Vbx3yJR4MI+pRIm1GOoB6AXY++dBTi/ZeEtbc77nqQFXB0tNhR3hS
QhrCnNn8XDMbLAhoD3BYEs5fIcr0D0XzRerXlb8TNX7HHEbzVE8KE8AMVL8ue634zozjFuFXkggP
lWHB/KT3Q0tNoYfuTMc71vBJulUYJ4M9r1PdWqBRWTSHN9ygOknQ3Y4zMEPFQc/+ge2oPg6TGhps
sWGXon+ZH7Dk6AVjUp2XIU3IyF/S2GB5oxbWDE3x92IHorCxmcEdbwWtLZHfnTAo6fXVd38Eg1/D
752RnCj+AnZiSlz4JpPQgHfUe+YRFZDljWgmXp6Rj9lnDmXr1FkuvYkwl6FsaXi3Dppa9OuApAR6
LGZbVQCdi1mps6o9t49EhD0A7C1k5o3Al7ygdTlxOru8LMFKMIJDvkVcFOL5fzI9TvYS/I2i2PRY
aminPheX7vxTfCHOMoP+ZCbRAIyvt3+d3O8DVcHfaf0FVDYvrxiuRIyhTyTvr492AMr9R71u7Qk2
k9akB7PlUCCb5hNVfk6BKjcp6rx6B9rPJZVmAxWb4AKADb/9CZTCC9vsSk4re5Z1tE5fP3ftGfeb
ia9FxPAFKgjajyzXufJiVQ36dHa0D5uhFr8+lFZRvkpyv8xhYcDPxJd8akOwrWcj1wn9HhabFnPw
1u8afodvjAY3Inx71eyHPS7JOvqzHECh5RkGm4RoOdocdwT1M50cVqDodmrivkHCSRSJCirbay81
Ux7M8SKeK7pVV4Q43n0uYxSusMUIj1hW9vIQA/U+rA/OmsIBMVK7jWUgDyV2XUdh5daKCHXrTtYx
rAxw/1Kt2x9DeWtvdbghCz+5X499IRoFWPlyAu13k54EpAW3OYcaKhRfb9TE93nsoOOPv2zPdbnd
AAcGGg/AFVlV0SSbaWX+cdF7BGV2tm1zUaGkxsgqF3yimCjCxg2DBqgbkViC5JHRIJjWsFt7mat8
PBtnCOMBNjeOzysz2+af8uksPagoFqMJYTgjBlz7vtXVlywzHsvL31wn/eur0Zq45D2JL41a4gAr
HYZioBiXSYK2bajmvs4ztoxrKiCUJOYI0Dtk5Pr0ASmC5eu7sJL4KiNKaKqFNtkRGRMP3Bqec7Kw
xJaKSAvzQ0G+UOyKXwJNPwsYKx5xNY3F/bR7MAF/ZQjI2reEVlPMzA3elXX2AcsylEJFKVA2OcDV
JdtkP/q2t3YzIXidtbtAS4f22YpTQWdyyPSYHWODXTatTkjWAKoZrQtmR5nTg7pd7oIBTQ1JY/Re
fbfrdlNT/erR3nVqQdHdbSIVD93pX6/9m+j0Q+xcLcJIYV4f4974ckXhOJntR+hHClMh08tcF8vE
0RiPoLYTq3V4Y278uPIDjpdwu7Dq4BNbdR3MXaCjFBYsjrdmb3BSC/ZxDcafFicZS0dUWnnkLCPY
RVzluumpPQmZUaqHUmI74BpUhFCHtjrhfOInkSCwF9ycqG6dzMG+zVJp7syII8tYU7nQdSn9lXJ5
9NYQBOnuJHjDFMVhCHxuU2456Ut6bEsll3NR6jbrViDnAZCBvULawFY8L6uu4Wjlex5tG1JssvOx
QxwXShA/KbsE2kudHTEt+Tl0uXuveMQRPLNCcdMjVhMc+Zd91x4lRDoHPP50wg7Go2hWEiGhCKu2
vdaEIgRY853OcoQCAtgo6XvRsbAesUVKj9sDiksxvQvGh+IXGBpi1fiw35XgXJd9rLwCxlpAoDSp
VxmS95kYlOn7Wp6HnsU4pxq3yM7orGZpQDfVgyFljJBTW7xVkM01BWDWp+WA8+oC0kgS+qp723Io
go0C4IuQvi3mqKvJZVcGnTTYEiGa2mpa6W+tP4L6ly85d7z4fsVERLBBbX0DAwRNVwqhNoGDzMCl
SL63OtLaMrnRR0NJqm/9IM7QaQO02P2PemzA37k98tkdn7csR0pInqQPQ0MoeI3r1n4ABfUzKv03
ZN0XeGDMKJG+pul1cFpLezlpvlmzvqDahNUnAyEiI2AIdpghVHnwV6H7YFerXnsuASLV5TfITyOH
C8KLmrK081yprCLpqN9sDC7p3XLxyP0nLlf6uj9AmEmoMBdzAMqbCRhjMVojCRMX/SrYwstthBNY
qDh7a5KUxXkIZY/E8YJOI6HDxMs8a73a63K8srImHKKDGl1VYzVay3CHlrkt2iwChcLdS4BUKiQq
zf8cv49B1XrPx/DQQg90LXmKovQgl5E9QXOErfDtYlix97HrzBaHfUSDU18vdBSmgs+mvnrkH+EF
SSec1g3ocUzBw3yW1NhJerr7g9rIdnxAKz9/448LTIBDznTtgN4MmOKBkZMM6g1BNjc2jFIqq6lZ
zk5LbrXN44m4DhhOAFYBJof6u1ulMWSGAgu6zsy+TrrLUBGoDyrpg1LCmzYLp8p2k17dMvgpSgnK
PA/yx34VeLLCTAo2gcoKsys0ZrUP1Sie0OIAEUiB1Eq7z2ijXWf0bO19bvmtOouGX+fuli+F4BlJ
RdIwJ7cL7judol93eqOWTXWzdYenze7XvrbBH93/95Honucmq2gTu/Q+abrlKis8BnZgh+fVTCO2
lqOd1xMKhVptJIUHkXbNWaniGTVAeSefAn2J9dzhOpUCWOQFqhwttMabMu+UTVzW9n91l+bj2abY
2ExDJVSvPLcJ6gaqG1ArSNeIvaakBbJQB37YDroIV5aflxw5rYjq4JEPuh1IwGIwguQW1jBkcVhk
hJzjdMVtyCmddhIcaUrHw1tmmdpLw0eLSM09L0gfCNY7S/p6wjntCEl6QjScXvrpyKqlGyLIBQv8
dJaxJUQO8W5yzV6X8VLG/kjTy65avwv9b0W1vSkobKsNsk0vjYXIDh4eadDelKXw+CCresQWoJGE
YtxUpqqMULcAjc/X+7XTRpV7kfr0/Mclnp0NdObfcE+71E43DTJZDdF8CH5xU2JGsIcOYzLuxwAz
d4FYAXo+aaIKzj/H6f87H6+q1dG89wPem9x2Ucww/jtBgCre70GScvKkobHWrYaLh70wWXOBnqEl
u4L/K1O85OOUiV/4SyFNLzw6rsDw3mER/20ltz2DWWgLhBcxJX6ovhwGinp/KAwd0L6OzVa0qDmW
gu0sJVlwup3tlUHEcV8p4Vged2k0UfVpCPbNREV+LE78iIo/kUk7Sq5lS+xwZRdWTi2H5N+ib1db
xXRknu2a7XnWXkfii01V5n1QVyVeqJATi1elVSgojDJmCj5Nki/NoM/aMdFgp0GxEMZrKSah95ol
vY/7Bclw+7ZUoYh0vRhF3bZXjfLY5QEfBVOM8Z6OCXX8bFdmiKmZhxE4b6QM1stFhehOXsRnwipV
dfGjfdHk66opb+uebDFWuJXgaj6Xa3/zTC/t8u9TvpbnM42P3TPRB1djcwjUEXzzvUIL51Cu+ZEX
Rt5aFnBa60dhhOYm68ROCE4L7KTBZgxsI5gcvdjtxwPdYHZlHfig6kfd3qgL3cNT3Zt38uZ9Y1pg
fjJpaYNDYa3W2AisCMWgEpvKswHBcI8Hh+xzolIaLOIi/tv4d2PoG9xqC4LBralU9oHJX1gDxePZ
dhIKV/Rc/hv7eZagrJEvMEuymYvmzAmlNH5QxvtgzfOnXqJgXhqXHvHwbLecmIDq5msvgJmF/WkG
eoHHnrJIqcZeyFafW8STlS/TEDbOxftnjkgzobUr69Ir3WJ7WjzaqY0D3LE1JxjSjCZFFSrw6Moc
wPObOg2JKbLHKCtpq4obtUs2uRW4akxPBnRWY1zvD4p2UX//OjgUGh+9vmRGuBm68+vL2u5uEDui
BTBlyXFQOe5I66CZFhSL3XMgSZPTHE3fhgeXri0+T3PEJ72+Iu7uMuc8HmV+2vfJ4s+HacVGP5Si
0DLM+ds++VhgQyqXd/uncvjohcMGfk6TJeuAA+mOJVjAiVAg96u5J8sW8D/USTlJj6jIDDYDgYdZ
hRvMbTUL8FnggC75Cx3nmvXH6UPBnVG5ln07zrgepRPZI3zXfvBLQOh5SD8ZJt3JLV45MMUVLJdh
wHCQfqm6cArKpbaLOEQFrGTy7HUswRFutErXfBJNyQoLZ52lpLawXndiq61os+dYhn59YR4WqixJ
JALwhP92nK0V6PjynykLnwfeaKsUk8rUGWGQnfOtDADJIe+awRzHCj42EeQ5QP+oZybUOUppUxWX
g6APQTbhMmZcsosVKxaJyFeuC9grFlmWBKpwLJHgNS7ZlAZxYUcYrry31mJO9x5gkl45fDXYIGNo
srzOGV/qdh+aKwHYHGYUi/hkB4raTrLdd5P9MYRyJ8DINahb6mofLAn9eB4d9P3TrZK4c7NmG3p7
KyhrY0u7XgRWOok6cZXUeyx14tZtIkEDbOu+z3DG7ADu11LWN++pCR65/BFN/gRkgKhmimS4le18
TC06dSdgPESxB0znOopRpF0rpjXJlfI4rA8SOCrH9VV6UziSCkX4W176FBD3OYk5HuMRkk5grteU
9wZyGOwGViN9tttQWQjtMcAO1foH7JUDDMoU4JSeaTm8dbHpAherYth80rwFoBybzFLFPZ9KTB3Y
sZ7LnNxER66VyHk/IpUTvQK7GVF0MDeE8YhTk3LAWAWuWwk2jfiJcEqNkNuBzFsB368oBREru3Lg
5BZsZPRCEiKb/sjKEvNguPIVtx7TGJ43NvHBNQEdLv/MWalnSDKA0Yau4gb8isUHznk+qmd12ulm
fZMlWqnhMe46044+N7qBaCkbg3lYsJEBfrP06zJi81tDjHTUy82KMkgCtl2XR9girX56WNyJ1zi/
r5vTuD2611G1dVwkezuNKB8LdLogD/iZ/On18ToSFQal9jYEaWvtb9x+s73WMi0b1hNy/yG1nSct
vu2UUkH/WGj4dRW7W7HZVz/I4UTxOZ099bPukEpggGRLe++wJ1TJJM8B8p+PVnfprkorOuvNBWAC
lZ2qx1J8+7jXe+txAZNW++KbjsEbC8WH7Ikya51RzwSPhOE3fYHfNMYp9JCTQDup8iu8DZYUOinD
uVJUaLFTvF3EjQ0JcUYOraONjXUIlTDYJ62GPANbXBxJ+HIMUcFBzxELyvwSgcOqr1besbvPcPHY
65dCO7tehR07Zm91cIdbiYYNI1pgnZ1u680zQf2g/7tcBdAQ4rCK6zGKqqHzLg/yzwC+N3qw9/tO
YuXCBuASk9wit5Od0HI0WQ1HovQNB+MJ8QUeknWYLQtpoijxG6K6BOKF/mJwKiCdEIIR0biHLWC7
KtK7ARy1bNAY2e6qgFe0LY7bqra1mX1nfpYtlpM1nssFbdJYZyhU4P/I8c1MbLL0mBo10NZ3MCJb
VLC/cbE2E2IaPzfQK9M4yxgH9JE4BNkdCOmy3bOStbkQ9XLu3REK++IgrxJ4BeC3Tu/cdAcZLVrg
zlfVXuKDxIkjaUq4eJ78ZpShElBeLw7O3S2j+z465GtR9cOAZxcZ89pjJIY2vdw5JyL4in3350yC
aMXUAY2wp6Dr148RN+DUYk1L1pcKSusIWul2v7u5w5ogJMw3Qov7AMoJuNpuRTJYT72QsTxntT55
lJXNj62sM88o4TtEnq6IuKrSCZvxs+JhlI55Ph3GjFzPX4i9Hi75oml/4cQZOBPl3Df0RcGfBJHF
GETS64geNvh48czGImmgJYA8RLqIr9u9Up0HXXY4K0LZ4t9VW2/4+/C5QHvGlhJ2ow9AFwmHkZ6E
OLFp2MnmdDo2SGK3O80U3iXoczWBoSx3Omtyo6POKWjP3Otrr2ucFSfyFuhG70R9XYyGi9fQhXPG
X9b/BBQb2c3UVk1VM9IP/FHVmeRQTC70k9CPwjm9f1u4/jd5WIwrGdlFbkEKTCKKisFH492+0NLl
2gvEpEe05Hj99F/VeeQwgzM5RPlqaXUOPDpEu3gpgxtQMTfZR0ITm1oBvnYKEn6ApI2AT9pHupdu
U6O3PLRQIowCfG6FuS156JAB7k3p1QGjhhNYdIBG68MYtwTkgWEKH4QySD2EVnQt0YLqHEvDhwoF
i/Lv3wvzwYovj1c3BQ/h1ZOibr0Ww5wDbUx6SfQuNc6+aEKM1cvN8vEUj7/J0iT8R7JOshUkgsdz
L6jD4pZOz6M9IVbdJ+916Sa9/bTb9szvqAwcVUyefVUtDDfilha/2C8qTFQNiIAQNylmOpMTfH1Z
EwVIo2vk3Kg3xUA5l7qNli6NgxWOJ9gcX6dBT05lUhyXKsCZ/3iDr3qyqPuN6CbuLrOrq/1adoi/
Isw0YzRpJIemofu1yRJL/nSSz+ZDWMDAnAUX03zfRoVeLGKnUWOfnb3FHKM7IIOhJs9EwtwFD3Zy
VaCtDbPWzHY5slIG6C9px3Wn1sgDTBCaTyec+Sj+J5qEEOCjnlSWVHUN2VvqFez25GdGDyxbHWw/
rNodDrn4Xpb8tANugFxqpzbZz98tcDbOg3ulAjjEPilG2EXLtWDHIIPQGs9xnnneKzxbtcFtsxH1
vpvN0VSHZMa5hKhNUz3bvtW8XROnsxY2JYbCO0YA4H55/Q6Bx0W2IKjvb5dKuzmC3TpCSTNek6Vy
sWqMNWrNLPUkDe7VR86tZcns6WQlVFATLZSWDhU02ODSDPDW7judapqagNQ1Yktkl1GgX7FQgh3X
vAYK5+pI3wYr7OU6Aj/trQlSPBUcmIeXuuaR0skAPOE3HnSsId+VxqOQir6eXkZUAD7zYTODyl29
N4Jlyo03A81i2W4Ak1RidtRQVVorMdCOzTR8OZ5YzC83YNzt4GjxR4z+V0cxDZAX258U4HoIL+Mc
sJZuz3v5xLbX9BbgV+/9dz53GDbugyCmHO6rsqUJrrMCSEPbruU9F8ftgdgCWfer6Hd2beACepPP
0E5r6KdXQvyl1yUWVtvDIDpwuqBk4vG6cfHVp1eLoywriK7zsLr7wEgz+coIipgyquliQszAHcW0
o/I9CkJgKzLPR8apbXGWgCca5vJkSFoSvatkdIBDjBQupDvq0P70YFHQXi+I4CUnlce1AO3yB+/w
wm+Y3/2KlYyTGWGpLLibqcBTFSDwrWMogFWAOGT4cY3rWVNhV3w0bRzCbAlWwQusyR4dt76fMv2z
YrcgK3osV9Jz3FR/jk5isGnwq9Q00vLBdVo4djfeCGHwHdR/PpkF1SpkuPWM9y3v3Cqen4BdAIVO
42oPjNFdxpnnS/VkoPlYKWrl3SDPWAjqtEKZcpqKmNabo9KdD54VxlxFG+CjHe/qIOlX+H2beyXN
UNsV3bWAzhC9VhJG8/ihtCz7jixRzmWF4iVXEx87/kv+vJMuV/BORrjpKj+njMJff/2JOvlwUzQe
iKddyGRIUA/ocMqnkWG8TQdwFq1rQuv3EIJUxSG6/SLIeXCxrzVFSmLIL5hfrMMbzMEyG2fn4PWt
or5FpvRLQFOvZ4YCeL7QtaR4Ob52wcI0mZnjI67t0PB9chVOyZPgGV67cYDI7L4X//KI5EesRs6p
ybOAhOJ9Ot5TjqH1+4b1hOYlQMRN+S3l4lrGpotVcVu9GwG3gce6SRTDV+bKu9o8kZ51eJVcS3VY
ioS9pBfqZCvJKFlgLGqi1GPb9vXvrJDRxFipgb9qCZO6tpr5WpgScOpuxLUEoyjD60yJvkW/eNpI
3yjw4t04RdrZFdAukSpWnd+xSuqEKGGXSEILvwPM9ruvev3H6JDuNYjcc67sQ6rq6ngSVI/Int4y
Fd40bcoaxbTeffOR+Ryn9Acx5pUoVCaGf524SeyuzI8OXt2VeNLHfcwLQwOwBd8eGOQtmMKZ77Fc
lDueTpJORFCC85ODwrusjfGJA6fEsnS361GgPyJDmDAjLluRY/z1voml0BYSiCL5MR3Gvxd1QV5E
HMGiThoQFM2hwgvIQ7a/y8EHzk7paOCiVO3NRD039mhBB3ZAbx9ny4B09ahLQiLWoEito8CvsGOT
CkU9DAv1MgpvVVFiKsTd2W5pvOCggzgOK7xKhqdg0G6NKOLRT536k2m+NBJ0/VRn8vVxNJ6XOZXB
MqM+RJ6h+GDR0+JZO8PA/FOMjqBGYBDdUHLvpULzlVfj8JCA6/vF4dWDnBoGIIuJ0WlBvahWWv20
nR6X6nLeSzMr/JD4DIWOvYjZIofyl4ypTP8SgFGtTghlKc0QOLrnxJGghgyUFS7xdh6KjRP/JEWZ
MaJv+wJV3jN5oCEqoE5MEMWcE9yRufsBiOWPgqZrmsbQbJeM+t4JLnn6W5t7n+mqOcZfCqaeKQOm
q1LzQqq2fMAaL9G1Cb7uFeSqTOBNLE1zidJ254RSi1lKpepys56POkeYpuVg/2fZ21AzlMpgMSCO
i6uTvYXVft3oS8Wms9UeLuHfiVnYgH8+CYTBsFN73k0l6SOtBXiJBOznILzN+2d11S/ufMrbS2Ky
DI8MrNSrLQhXhpcxuFRQIOTQ5Sss2lPkerRdNP0tYuiWLTzWMt1VFuE/h1JHJ/aAdmwQSAH03z0v
QTesSZ1HaeMHAhWewqj/ADgd1kLrqZo46RhQJoA+vXfaPr37w/N8U/K4nSk5U13Q8Fmt1zqoeyt4
1jitG5KwnOI2eg7okzHTzFCLlcD0zmGVvKa4u6jRNK8iLJ2gwmmFbXAkD5chw8g5qxP4sObg/enY
khFcw+e3DiLu3v1AtboHTGlAqmhpB30Pn0KeK1HisYNEFrJb13OnS7fKbmy0qfL/NoUqdHd7g8OO
/Bd7QY+sF02d+WysKieSG9OrjaCM0R3kk/xT6QOcKTPLy8bSdO+BGRYQPK62fYjkgImQUcKlSOzq
yY5qXebePa2sbILG+CSmM2uc/G7o+yWGiiyeLQVZXO+XaYDxBwBvVdy2S6TD2JXtCrV61D/eIiCq
xHo6E4MzrT1m9W1zuWM9XAU88tw+9ID6gNVMcTpDB1aw7XTxB8ITDn58nwf4uJ1xNLmMTth6+RhP
LwRNmSpGRCW4RvYq5MQ105foTWXcwaLMjhIjmYlxP2flzvpiz4pmJSWItMSwdkj+BCEP+Y0TNDy7
5dl6+jBbSrlArGHLo925G6pW5ywawCsb/r/5kVqJ3ycwI3+st+b16AoKLKuxThl50llfUr5/7FFb
NXXPpZHuy5i/WWJuVIv1MskKE15grqNGquanmwIp/HtYrGAzwCCtCCgxIuKz/VMmkRJB3MWMp74I
0nwGI344Ys4OFCzACypzGMyyJzYHgHO8Wqb5f1lXXfxc2r4+q0fJCrDAZXJGB9awUGAY5UBr52dl
fHOEQZGcoDeRzpsZwsQcKVpqE4iRAldXgTTlRxCrreW80G7G+sJ/QgpsB2uI/PibY8ikZ/Vct2C/
2jeGtfD6cVhpQYN2zlZOwgUCFVDbUCkIPie9Xnxj18Mge338ml6DXiCcOgssFR/PXFETfmyHf3jY
mkhSRofMhQ3D+c0fPdEmxtTrsNlAIOEuYjsBa/n/c8w/1fxjfu+we3d22oS6KzJOTgSjW+wSoQql
nW8kgKBNnmPJD9jaxdHGfVl/k3C+lZSbyTU76HyUDNXIJwK5ch1axI5ZJwpu8chex+qdKKTs9y02
TBHdNCx9g9xJmnPi6OrFyosqFxvuBc4g8/qeIxi8ZpC+UavopUbSkZPjvJ08gs0I5rNQ5TMDmV74
4dNmvCMu3eyKFg8RxKe9GjTvCSdJq8KoC2G+ySU1f6klZgXaS8V/UpvanDxV9GjWdQpZ3B7H3r/Y
n7ODxVuVt4S6compfcJN9JEdo/16XS4eFBIV4vPEvAkaQX7Ms+FTzQ0Z9GBhdASmd3v5krMFVCnQ
tNjHuVPwE/mwGS2xzXnHHklXzB2UDffqK1cd2iNcFhviI1ybVOq7YLizP/RQQtnFDXQxsac4Kqcp
8A90QCfUutkQsmMjFVaZ0AynJa9mvWntqG4eFeu+WIHBcUr3nzll74cKmh4pHu2HxEBw+6Lrzy50
ehh+PiDfGIv+WcXS45p1BK1/FBQPLbx9dSQ2TCwjGxtCBU+fJyz9SAuGAZAv2n6X8vzlVpOK/cNL
QLY62WWi8ILnCeeq/McZd8y+hPtIT4WjJE8hQhSUHyJYTcxj72Fi0uWC9MA9k/WpjwwTFWUpreqx
E1bHwY/M8P7gFbHf6mZBQw1Xogl+XB67BHwkeB4hT3bmcbx3tNOqC2Mwfhvej+vjLm6cowaWtzXz
BuQgx6DSu6A/kpJap3lCoo2go7/ZQednyVgGVBVSd82UoTH4lCvHsWimvv4qwi5JSn+tyYeFPdnV
JkhsqP8PnbxI3L5Cu0/guhuQXNhJ9oi7r5LOsQcVNJyN/5RZU1jhRAwCf3W/1r35bI4A1ePcxgBH
cQk4lWCcuq1aWla8aI8hTvFcZ0x2wPVdN5B8XM4PBhM6W+cJLPCOvQr+ixs6lPGheP5m+WEUEXvb
mlVa3EDJccsQuahgmUivQ5nztHUYtUg88fdjJm06EfFD3VRbnh/sKwthU66o9/jBWxq657Gl9off
opzd/cTpXupU2mMjOZN9/B1UEA+Sc/QBAdwcqlI02/OUxHSkc7JPZBEgC6IiL5SqK19VpbRgVVo9
2im556t6O9j49v/ZcuabBIEke6iC+txVhs8w/PdNvBd3idHW73Txk6wpKwq/RPWeHQwmq+Gqgry7
j5TAoAveeZKmXW6/vhKOoWJjvq3XRA388Tzh5fZZOn+BtxCfQI1aQZu7jNuxBs0hfv1JLL2fPAD1
lbfXr8dDdzLRalMj0ba3oq6HmNimLnpOorzIUhteAg8kEtyaNxZU0UQYYCStDo/BxYP7xKubOmP2
uwtnGFPeXIQDVrCpeV2Wu2yud9JAQ8oItfwnp8alZoEsdq3kjM25wBUTcnwDe1+jfju0/Cl2pjYp
QTTlwad8w/pA4tulJsqpR5Fpy0mWizIfsWtJsrNb3MtyEvkqKCUrxK+AnqtMTlZJO4z7p3fRAKn5
NNfZXRMaSD1NT7QR2vadcQY/AOtRgfM7YGiiTKAQaxBltBKlSpB7CZBbRd/baTRKGdvhiJKd5xcW
YAh33kCSYpAyzrvV6KjwFidjOYhT251lk3z52n8JvDosARd5jk77LFDT0tCall/9+N1bJIOh2uen
owJqxqCqoAqPgoUa95M/RTIMVgdIOJyzlVPAToAfW2P6We1Yd2PO2wS0dEGgmzwM4BZLds0/yQta
R9aULIB/d+433I2iArWBLs9K0XWaDEUBt7XOHzgAOECIIvf5XFPRk3jokppcznHSAg8iDYI7TTKm
7rbzn7ApvsHZygwyoEudxXqWbZ6oib0vJlHV1J3DQNmhFF0sTN0nLT1KH0g20hdYlw8RJCQntD+9
0OUNiyslou7qcsOZTJ0maIMnYCS9/E0xMWVpl8Swtu3HBjh0rYjzp15G0C7uaivkM1mED64SvSzt
NFJg8qkvcU/dy+78hRVc4QNp6ENPjap2eHWd06BTnMrNbj4MaN0QBclsHof6KI5dwoYAL3+FrhZy
korX9SDDBajmwqDaA9TvcS/6CwH1TyK+ZMmTslIYpwhnMcu7MJyq4yn+xXFvx5FQgMELAMpdbiXo
Lo4vJBIPCyxpIdpbY9DCTPWUslhJjCSeT2GQu5UHDoMW/WinwMcQs/DtuilA1w+XGm2+dILcOgmy
z9WTFdPZl6omC9HUiMdX7Ro/IIthDo06c/l1XUiyLmydToOspGkUWN84mrlvURfb+8FZNLqsVp97
Z0CgtY4YtmasfSyLxGEJRJgZGWTXvVn+K6uLUzRFKwrw+4K/N9hEI++sZY1qFRmhkHT8VPvLdpla
gEzNCdawSoUqL1Viyr4USmhavIyUEkFo3CctzMI0Khtlvqxi1M8RXtbKeF4YvLuK+Qn2cDUgGQgh
IeCf65yILQCM8H0VnexQC/bkZledixqsu/TC8IkBoLzVr3Ae4EGWYJQMcXaXO2aEOUN3tZR12Ogo
dawt8iwg5wzitcQWic3eogM/aAH2lEUGRUMLXAhWGAP6CkrVDJ1NIYpUwSdq1RqcQbQumKEFImex
t21RuxCOO4023CNQR5BdqoIgMAFq521mfp2YQ6hYki+hKa+QaEYVn1FSjIWba8ix3Lx0nU+EDtuL
Li0vMbOI7w2CnhY/HsBvw1KV0iBDurMJiJZXz62t6zWDVXr7w2HDJF00A9ltdJR4jf1c4GeDO0NX
hRqTToSHkXYq9hvwOPz4fJHEI7vQKVhhShwESjE7VO0jl/zAfhl5yz+cINGsIiOY/3mt2kSc1mZL
4CwNgM6grlmaph9/9E1t6mQGL+glRxt+X0CWmJcycV11H09rbRGk6N5Hg093iNr63W3RrAfHVRSW
7RnTsdc960zOARaJaM2sufeET+yvq6C+InMxGaP2WcCpdVA7vKgaaZc22tg0PGuZp3TSgnrX2GBi
40VZLBV5SpA6NkL5766SiWWzWhxpe0bYLKeL/JgDIm3AQlmzQQGeMDH/tHHVUZH/O5YiFBd5sUm7
J0C01AwWmmSejCxWrbawaUNBD/kBwNkxPGCNmobt0VSuzkmKFleDEWuwb0cT9g9QMylC+3BtgYY4
ZuIZjEK2nLw7I9XTm5qQbtie7Xv+k1Kxn91q0vauRxvj9UoClB6y9Jrkqdj7w+C3cpm3tbrBJ0X4
R5kCQxNURibPCr/O3SBFYHgejxfKid/v6m+7KlSq3MWHnB+J0FoIFjKUhqqodcBtlRTM5IEF3p1m
gE03WR8Gl1tWicB0wT8jhVZ8ZSiHvb5rzrXx5OJTRFIpTelBOH0b7qLiGGrRW7PVFvASZuh+AjhL
j/axTVPuspLvj4FPTEVMBO1KUCdsYUhmJqqEVQBVPuOW+FcXD4IFkMSNDEyGYnEPdwXGtkH3Hur0
vpns8pMpet6xe462bEpODJlxKwb/dhtTOb6rEskseabHQCt5qnYheppWMca8sjI/WZCHXTEyldzu
KyNgeLuR0zduq77ovBYp7p6vZTOHwmeBfzfRLndCXv2HAYU3KjVaok9JyWaBw52iT2Z87GJHFwEP
mUYRtpoBY5IBJSBbNEdHoCguno2n1dTgI/pmUHgU8O3iP5ZL/DQJet3j8kPDuTpOGF34kzABirxO
oU1lPiXc/sH2cz4yUfxQecIDrL8pmTdCl1hi0ce1TTs/TPGc36UW9H1T8PD1Y9oXQdWUtD/FXpQ0
Q6hQ8kmhz0pJ5QgrMnfw30dLrgt6rgoDgutPlrJjrPedlZpqxGwna6EV+z3FHtpfwQujrHoRrCnc
8hbeMXv8m9NiqoJNqREPPUwe+4YrXCaGfJWpbdieuYj+X4KuFqE0/uwrXzyn0AUMNYOR7QGvmC5Z
KBMDL5/XzzeyJtbIgoh8okZf5+rpRAihgDCntoqT/8fAbHz6XqVl2I6tuTwgjRzF9Tvt8j7sR+xV
1y+tQFcHTpE//B0Ng3kMA3+G6uFwuwAwLDefzB9/47PiJCNW51ZNHwvf/AQ1GZlo0QO4CHrNTOub
xW6Qq7rdtLuXO0pkof7ALR75NTicpT1fQajtPMeRQreRcc2Ovqn6oyd9fbwvwu9yKvK82pjHPT2N
8k2x9zQCs+Ma7sqGz3mMxmYmbe4yZZLGmojz+SGE62Z8LB6YBpgg2mZcoudG6fFFIOWZLAr5tm35
ZKt0rNQL3L/ug4wXtjS52myUz6cnrMs+2P5kseTudw+V07e4UBsvnb5jFOBvGZy6mA/JB8y40fEF
bmJjRAltoVaTkVQ9nzlMZudLELTWPNieRZR38mtlw7bARssBc76uuWV5XBHO1eZS0GkbBC5iB9mV
l6CcyBrjuaAGxAmtnT7hLQstNILdSI27QdWC28eIe+j+CCF1t1hwBOZInj5Z1xzSwPa8gWmPEl2W
Nctkqe7ioZJYn7ucwF6Ha4Vwzvl3SFeNJBeA9h2ws0McLJau2HqGT+QjjjwYBk15RwYfe4Lqfcl7
HkwXKTttm7I/dFhmJc1LUnfliR6mtawdNjmyCsY5soPUhfes5ojLZ1L8VYwnArjbiTqwg0KIMvya
B/JXf7BePvCcxyfg1YKgOFI3yHheJa+U4UhR8a5JCy93IlROcKTu8p74VaGRMgZa8s6NF+jVwktK
rLJofBLefNmUKXP1kKe/LiAOjnS3UEvYzfAZZ9Nf856UXWJImUZvHQzStgXOXjnJuCoLiEP33wSc
2A1huDmukosli8U91CAJfoRjipusgcE4zMa9j6jy0KTUn0e7Yt+DzwAb4RiZCygZlyPz2TxgBcGr
5Q7imKopPUzmgDj+QRLbhv5cMN/kDO895hUm08xiUYwIUyrB085fRC6PHpIp9GYXbZ7Tr9fULTf9
WJFgCtzKcksR9zz+0DJcrkGJn1X2ZmU1XPDRbi9GmS79Iwoy88+Lo4HAE18f5dnWQIEnvb8+5jTo
5NGQVMmaoPOYOMtOeCCOJXL3Wb1baAggdxlKo/4napK0EjBQqOeyHVA7YCVVJ7jTYbw4IPxOTk8V
QMszSTchVD9Q5sXlu7nD85A1XqKBkDQFYkVmoxMqCRMm4T7BMRAXCUOQRrb/u6AGfQek6ci8hNcR
8dEvjxPnwM9Lu0NPykFbjOSLpZNtMCgiAtuej3Q/Qy5U8hwxTc8StDTpWPL5YopDWYct3L9TiRj8
WVLrNRJEiCq5BCXFu+F6H5TECJYAaNv2mJgZPpmfSaZG7z1EvJCKjQvss8ud/YZwKhKRIZgC5hxf
bmE3eKpB0LX8iZeXn5geH0sTIJpTo5rZFxOTGRkOm+JWA9T08fehC/r3ikFBvMlEA2yxJTWmZzsq
OQx3+bbHol1rYgIoGN7EBhBAhmGO4M7uAGkkvBztrw2dZdu5+dgJvxGGOCfxlmihlsMhTKbnykt9
UQttfBTH2IjD45Ta+x4UL30x159eD9qKPgSAAWubBSX4XO2Dr93FLbliLZdaYPBlUOzVkoPPTlGK
nu4kZFuP14If7it/RIs1e+0fRLps8oimKfQ7XXv+nhuW/gY+AQ6m7KxSOxiZ+3h2sGyfeSYRlIvF
rQg3pOj/xwzTwWocndhcGQlXMo0oV6c6thS/wAeaoL0KS3u2OFY3XHT5BpkiHKit4joJeEu8mBPC
cgqfpbGIoUW5sHSJEUqnne+Xoc7ecPzpLjkxU6+4TPjZdVI4AYQdDmQJm60y53doz9Hs/rR0qEbz
Qe7U06AuL/w+fdskQNGo6bE3J+7PlQ+oCwsS+DHAs8fSccctKr70s1wiwlywxGrTJF+YyIBZs2zS
LIh1Rb7M7hZ6u0rmI2MH7L5ULaLABm8RcSmtxLMTGzd4qS89//DRShzI7HEF3urFzPh3hDtIY/BX
YEZwSuN+kcHp2WzAFomlK1c4SiyUrcVld8ekl70fguI1t+sPwzGg7V0UvK6XxWPrGwXhVZ/t1eXK
wwf8xeGBedcDjZXtS1meMT/kDEi4Oyuejq7NT+a0XSnZ1WX2bLJxsYmGmChF3IQsZdNRVXd8XC5q
52ry7AobhhSWUQxWikDoTTPSpdszVSRV13Bagq3WCRkd38uloAJowOg676pIooJ/RF5vl0BlMPlX
3+x+2lspcwAZxu0nv9tXMKlVIn14XjVDjmwdj0g1r1o+gygBgrCwy/0DUoAT3+gGNK3Rp9X15BCp
wqwz0i+ImuQ2Ju3fPH6JJ8d3PCzrtUwwfe1BiH+2A/fGU3ZE71YgdhMb3JeVP70rD1xonGQtcGs4
orZfIe6XZ0JKr/F1ys9kiPkrtgwrXWiJGUCB5fR3HabJP4oXZY1AG/oEBG77g0WDNSZj9GWwuPBf
Aa1T847s/beXmNU+vt2Agznoxpi3QHd7fTuZMLxBq2M6QgiEqGm1AvMlH0RLkCnGzYNpbhFjNc55
eqzbMxb+3hXhD6Q4dOvCSrNXG56vrgPS64B2thFa+RHIFVG35ui/wTAWzegx+OdxNgTxCHCMIKI6
XDLC7sRe7jh4Iw4rVS+Ep1WO4CcPveN/QnGcl5P/8NdJM8/tAxD6JnLb7o1X1JB4QY+p4co+2Ho/
jozcm7Hjl0m09xCDW9TIAmHoH3WVx87yHz/89J8wfPoh4grSBD/XS25q3KnSHSYQdPcFCRNLVHjn
P0/pXzRu7h75VvDje/ay0Ci5jWxcxE+j5Fsf7G9rPFwZhrhhNVxuXupxNznpnLokF56Re/3r6aKj
9HJDMnGre+n8439j6uE8Mj9qoGln4hIeOtlvt1n46S9sm2vhbFzC/zqSbIOBJ/q0EvMd5Elp8hH0
oD4IdRFdCnqy5UVAC5+0b85LAr3aeHdHCOp7BIRtIU0u1/eRaA2x+OxVOUde+zbRA9w8ObPtReAH
QSyKHLN4Nja+saslNd5pj9tcx2c1Bmkzy7biSqTh6GaW6kxBk4ki0EqBMVophDZO1h4hsxcnJqFE
8e99YcKSsqzK6UZw6/N8d2pmXKz0OCedi9EqVCDe4yqvaIyon0pRG46Gv3JwEwhgN2dSzXCNC9tI
CQo85EZL8pL0bYYf1jvyQysEm/tGL8sQbf1DF0hMUtGhYJXeFll8sMaxNOMmDwCyFXFpIpIfxCYZ
efxRZlXPAZm9cE22eG7v0rp4GelFM2YsjRfn747bw5XovaJZ1rSxAatpkHlKTxvJhq/1Jx4tkX3W
oaVsu3IEpwULKd8jtoNGHtEQWL66VJC4ZYfsjvN2ArUVI9yPw54tNEM6CsbAKKiG9KZXeiYRQMmc
RawIB44PxVKw1nmRth8c5XqM8OpfYv+zt3bHqYg3NodUGkqCp6Dv8dKRNTQYIuxtl8N43ne9Xvmp
OS27zYQAh33ZSJIQlAD6Z1qc59uh6KPs/RjJ9kb0pL4kMDW+/s0wMqJhHUQW208dkxl7nGXI3TAe
kb9V2OFrWvWsvZRDynkRYM+PzEEYj3jtNyfoZVXwieD9FJan7w977DIHOOncfZB3X1nSDBJ6qmoZ
YEXwv0OwIKEsJCi39VZgVGVhTdUg1PbQVgOAa2zs7SdrWCOfJLj1K1Skp0DIiC1uouUYUymp4k6H
wAHnfLbTUAPI7Sqhf1+TUSNhN7hUpkUUFT74WLxpKrrenK+OzOUhHv8pdVMEOOIqE52wZI2nbdq+
9NRMs7H/nT27rd3A1WLuL4Xe7pUmwxfya6CpUcTWI3gVYnV4KrtJERxtVS/PmDkWnKDNpFwj5FDv
yRLNw3bpmt0YZjZ8iPZ6ebHgFLhj0GxCtwR7+OI++rgDQFId0SiV9d5eJf8h9AkA4chPmpqfO/ss
BQreU2DhXL8Nr/1IW8msNOd7FGyFj+GahjAT2c3orIIo4Vr3Y4uULVnaDVH7A8Z0/Aix6VFHAG8s
hFm5l8f6NIGanFFtK4Kw/7dXzMgKlutLJG1YSFcHmta73IYL6DDTsCh9n9SeOF2/XAHJsaHg/3Su
AGFv8mmAcE+yxZwGwjGSfUvjE5EV1ucGPcpWEfQzK8zJxtXqfjJ1eiKAmGPI4ID2dgoe0wiBLVTH
BhW3AI4rJ0XKxWkiso8dEn/8FgmZUfs+YJ8Jg2uTyKd99qT8FEwLByMYv80tWd91gS931cdBAISF
UZa19qogTSlaQy0bBiNrEmMLUDZGnEV2tnNpl3M/aa9qj45YECfZ/Lgs2k8hYc/wTSapOz5F0XlQ
OPPv/Ryyrxpcat0oYdTW8+Y178uN2oKS3TORsZt7UJd8NNp2d5G8keNKlI3jonvzbcYwzlZPPvvv
K5qW+PlxON/VwenD3AsZjfD1QA0k+OhrVMUK8BX3BJ6j7PemgtFU1wWkFffhOL1E51c8Hfr47cUS
FUXy8i7P3gDbGXBXSpINP7jFnPeesXJj9JyU2W3ed5DNbm8FLCt4cafTcopv7B6VrvgJEfww/lKH
KET0zNcR1GBBR4yclMN3qdJWaIIK7zEwjctVdcHeM37hqlK+aia29bc5ySEF+kE1IGFMdHRliB/B
U3h4OB/aeEV45cck6JblILZ6n7fb/R+3ZArhMW591hzi7YTM6Dm0NGCjSa9JeN4oH6tPGQRPA2CS
uFeDAvbYYFB9kwB5KJf00SamgHgDNCfxxYPAa1GOXKAIc5bysRJeluPAPDls71dfHyUNNlUC9K5A
OC+rXsmhYUobhTmBDgbQw0D5wbCJF/KUUIXhpmkYsqjCMVRp91eyuIPwoBAlhCqclQUrnVxuNlbQ
rYA+gW0sgBJE5tvgkDXJBfocDfmSbOB68MQj8AXH4a3Id0JW7GT5vaGuVm5lsHqpnLAjEnis0C4u
991sQFvqKygkU+3toHiNJ25130iisPcPzzv/Hfkl0iPomvQuV3rj7FRJ11RT2xhjoyjR2eVz8uK9
+i61jxga0HiePgpEGsAv2Qmkw98/BylMM0VvcUwTbIhb754DB87r3I/s/QVNmlcHD/ECOuiQM6ti
5Q3aczln3XLcVA6QbfvIetTKeT36UU+YiCEQTD1A1U1NXPofOXemCPROrgbWfQEdocBoVv0UBbbS
71Y4jbyYQcqoHA7z5YOtHUTiJqR0I+q+c7J8WHUs9M4boZu5ILautyS49pFXKtltnahTuk0s6F6Z
0mSQQEpn3m1bvFTY47t+9/N+M4K7J6b8JFLYg3w583+GSLPGXR5NhAbzdxaL9lQAs3QzRFDK4PaL
f8hTPXsu4v6EzwwXdfH2qee5jMnAQaAjf/ZjZpNWlXSGF/dUoMgspTt3w9UA3jHMyG6tNdV6x3cF
oensaNHPeD+511ieYbyKpMb2Z3JWvDz7MnEQ0+avJ7zqyvImmVHb9+YRLK9GvdtwSsxvImM1JUvd
9mk6YyOSMKp3PsMOehvwthfkTv3MclC4aQtjAajYo4mz5RG6JL5INeoKyTPeFINIEKo5R2aHVTG2
2OGThdMxUK1vY5OcSMSBW3SOCNWHsVlpyrrW7o3D6a5Cut7qN0XH5bFtjw45fKv6H+fqSnoAbsJd
I4BSh2k1fkCYrWZNncZOtqMgl097rMWSjOxtgDBNhcBJLGJ6Dv3g4WkyE9NuNI1j+UU4dzb+pN/F
91AWaevPasB/gm0lRXSX8tmBUaEkYxyMn8xfgT0damqx1g8SFgxeX6fsAMbL/2Wkc4srUPzciy9N
FcIQ2AeQ0BLcsYYP6dvUXz7djh/PK0HmQ9uTkpDgIbfzJ3okZipZQaC1QQJBuIs/Mzp7vPtrLJC9
hFD7J9ovpwDFH8WoD1BGuzHKRAC4UHUBG70WeR4/v+fRUGYhw0jDNvZ1r9AZZsu2XsmYKk3Tov56
FWmkfxOIgcZmh1uptkTc6/KfChOjVyj7VY3UcxxgJrt6bn/XSZbG4pdInj8xOhS/21+hLokrrYge
Y3nTYYEgh6vsdI9qe4Dh++0pY9NhLyKXnynErslLrQAG2KNcdEzSPerbxN0PObpZMmDcf2oEf549
2Y8LK8mzOxl0EBCw0hloq40uOVfKk70n43+gLmo76mSGgIhteEH3PV9Gz3UJVUNFbJ+3sOqs/SJm
+XdAIl5xPvAnI1jEFRj++4G5utkTNwowk2V+zUct79htyJF51mDFbBQKiFKT3y0ce29hzGKtSd8m
BZZ/AR3Q3nRk9T63y95moTLPtV+FUw+Y40byEoQs7/Uye/3GCNptjPdDcAaNGSQ9SSHG6R5Jx1g4
Jmv9TrB8z6LwoenCkfD6uXe7OwjX3tMXmGBvozvSUrtfN6Xa6brd4jIKyq6piqn8eYgOb3ur91Nz
vl4IjHA9sUvMFxh3OkhkrwjoRDE/cmuVFCiuZ7RRCXWxD0Xz36UVNqp8qz++LWFG8fqsCJaDqHME
a9DaafrOHGHBz4V/9Bd6XpYwq3d7IFm6m7byAQrWCDX5MrZCzJ/i/GvnmmkC00lQqj7acUbkftXe
IJ70X75opGVOGH3JGGUADX78HSbDK/+mYwuibt9ZxLjGWLWOzZY6V6V0CTLNYXhYYJCo9GK+Rbkn
5hm9aNn7psX043MZDJiGDOiTOPBu2RFmCey5Vz/Jb3Y4TbesuUwt8rUwRfuc3a6Z6eFfKYm+bmzO
CAwpDmGNuIgtdYSMIcqeD+QhMX1mUf2W0rTUzx/VF57iVF5t4PkYSLjxIKYOLi7JbhfF0QsKKzf/
1X4ejQwvplpe5NFZaTtTPmDpzMGl8CGAKM+dD/GjuQy8qF4G4H7nB/sMOE0b6eYpddYU1+ULH1+K
g7hOiRqI6Rgbu3r2Bq//1nlmIxbVHAOONgMXEOW2Gs8L1WtnWPraLf/V1LYNWpFBnFYXESIO8221
1nE/jhzboPBWg7dBux2a4YCy7gWLHk80/F5JD50lCTiJl9b0McJ5LKFNW285qV6dfiSFtGo91Ti8
8CxE8z2qpr6NfGKjRxNqGvT3QZeaiawa4wALnH3Scd9TvgHmn7PbdB/XVOvwK55xWmFOeAvUyln9
ygJcrxtuYmiE0LiDIkc/NipklpCiTrsgUfUOJoPsmPToXYAqoybzvsPlhXYWNbR/SlQcJUI6X6Nq
vFMCvnUIsICdYWtGR+4PN8Try0NviztAlL7MqEEozRMjmdnZIwnry2Qs/lBTJt99zYNaYFR5t633
/WguSt6XCqd0TKHAD/sTYVZZp3C/BkdzfR/ZaB9BoXduQFLTGTTm4oZHazIB57Tw1Zeb5EyXrOFJ
p9MEa8XKSinRYgTdDYw6m/5C74XRcW4Hsk2iBeWoLGAxe0HiRi4NjPIHrrX/d4FaGKw9Sl4vQNVJ
04zIBTpn8w1Y7n5TonVgMHoxo7AJxscDm5QM8z1RXIlDIIXtINCCmBgPEFRnDa8AjSDeXGh/kQz2
FSzS0tY=
`protect end_protected
