`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
YjdD3b0So+PqyFMLeJMo9BoV6i+F15b7G9biRH9+5XzVhriSW7A7texyG/D3LLKCvW4RDcQsy+PA
nkuryoGQcKVYC4VWADwQfW2C2DcmjfJpkMV5sx0Yt2Y+Y+v3O6EKUqWB+wtqBF14fYu1jg6hCqRh
KbW5HreGTCCHGK8BXoOqLBZ5Bs/eIid/6ZV5okHccUsvY7xR0SycX7RZVjfhtAWWMh7Mrjp5frb2
3CNdYDVE4VhzCMwNuAHcyzQqjL+0ciJIFQNTaKCE5655XUT/npvCO7TGzxJ9rjlfmOP8izqi6S0Y
mLwh+ENfpyDoZrvjEH0JQVrCf2djiK7wKAT+iw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="qsNo2rPc4d3lzkjErY5+pF4Y74zJJtCScFXWw0RJy5M="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25168)
`protect data_block
9J/F0NQrs3p5nCM8T708CQGsbwni4Oeq+EfpSOSjFIdMHQeWC5Gtc9XlOxvqrGHRqe4W2bGQQgM5
3gAMAMTVovCM6ojxYzqBxntkOi86xLj+YScF78ERPn4Pb62fQvwqNyZoJWkgUqK0oYoQeXlXw4iA
o7fZQdOryYAh4R4+FBAoYDhZmuJcsT0EeIwyPesulKDuIMDMOAF5ZXdQqVLloGfKbujyObmRTI7p
135XuN2ueyCtj3/Ta1kaeISn5zDgiGf4Spip3PCcWBDWT/8SfdHNubzw6eAUcYBFO7hWgFJuZ79x
adk5UShPlzhRoaMRY4HpDXDzIB+a0qmLP54ZAlWWmIxN4A6AOZSw6/HjnZ7yb60e+d8CC1q39E31
g6lY0fFDdSGFA/K7bJ/gXBtGE3pihIsiyVphyuhpi9wp2HzkCmZvOv3ZvHpTnqTn+mLMr7RbQE7U
t4c7o1JXIv+B+GwwUVA4HSa/zh24tYrETY+r83JWOCs9aWyaDeIdx6VJv6+C8P7s/hwiD7v3+KYP
RUCiwbMq+0xrgWtppraWkZ8ARyqzagnyfAqs10lWUb+xJ3YnGcFj6iOpSgjVKiGmWWu4jQzXXnh2
UPZ5lXB3t7pOZR5ADyTl/rngr5aAW+vaVLtvxZLYGZCP4uAPnEtAJw9jQbHW35dsoH/HyKPB8wbv
Ocv7VdUQZQCbOqOMXetHo46F5d27VHRbNol8HQHHzpYbsoGpPRZPSVSlwziPDSuLUhZcgEMiXnbE
jGz2e7PlFOksLQaoyFjw1MnNrin2g07aWuxPj7Y6arkOKcQs2oasDBtwvb01SjbaJlzP3X2ra/f+
dj6JX1FGCVDikpeC7jRmAQQLeSNEAhxYmEOL2ML1c93n3ljh8CLN5kHfdWLgGSVG5WfEhTJPULYH
mH1jXjm7UqkbNp6cPyL+vRMrO3A2f9jKYYwJ3Dauqzp8F144qxZGkIqVBRsQ1QgkVsV1xc/H5d5h
NRNnpvhp6ZjvyuGIgZO0UIu9w3XzRQlkN7ElO2U2YO4orE+A+Xq9umk7jgfI3qRCybDFZTVb1+UT
LrJOb2vytLqF/fYKm5MJJvlVQ89QNbZTQ0tvO8jjzmOHhTAAJnzG8aOBIbaSZl5gyF22muOzLpzX
kYVr5jjAVJvmAUCsXw0m7s9dTt7xaAUlIolX7yNgCyr2w21mEREZth5SkdPOmxMx/DvMbya/eOP2
LZ5+1zrxo/lWMZ+Y//1A8JUHOT8t87qYUeauuXxpmIraCJ0qmjSe4a68djIRUR+0jY54+0Ay46r7
K3iSMGZNbCdKSmr5TyPF12jbrjJBVA4tJHhEayH48picdh7qsFIX1eetqlcQSJEBCIerDgJRS3JO
xJIedgW0LuLHzI+Iqe6jvKhgixxTfQ9RigAHZt3AdESsE/oojd3iTEPb5Gv537v0HsQiWROLgbvr
XpJXJo4ywuoUbLw7CnDUpCpba/CtX58wUhkMTBTxJmumgpWsq6wcfrnr+h4F40ebsF+Ob6vw42EY
iKZwCLX3Bei+70+qrJMRJ5ipu2N5/aX1twzaTgQ/VfdOPyplkErkkV4fMv/baIjBlReOoR3wUKPj
ak1OZgM3EF8Lu37ALSJ/Aw8ebQ8urRK3kd1g+/48nuExFidHWQj/dvE4w9yLY9nF2PdoscMPyRUI
ihdFjcZtEnKZKGatq6B1TT02WHiA8sON92HbkkHmmp8NnoppROPdc6ofc7UtvQbI9AYgessoOm/d
ihyqwxWYO6EPWYVDxYamCrv6H7ZPR256Knb+CG0pBkXO8terDpoTV0fj5yjCTvln3zOHbYuFKIqC
JeTt+TmSZ0sDr7uWmbh1OtWHT792zjLe+MiTyLo51rZ8GRGyC0eZPnLYfU7o5P6Xdh1cbZuA29Su
juDwB3lTVgfZ9LE8b6d2LVUS/geGi0vp5Fg0ONmXWv9fYIQHNWCbBMCo3RPf2mnsJOj0S7eFIoIy
cJVeX9qA9ZrP/yF2DSq5JgkxWVrzIVuMsLNK11DQD5qzxt5Au70sNF6jeZHM40c1dcL+f9U2iZQt
xeTiLZYjvAA7/EtHAvaA7OxFYj+btok/1pstwp6C3uz1dW2FIZ6VqnXMXP+AUxJFOSzpnyH9e29r
s+yQHIMRVguCxr10mgq0Cnv1zGxygKLem6PK2/bQ2fArvDWfkDPsII26g+9dTmOdgU0qsQXHJYPp
vRG5/1SD5LFZ88Wj9mRmUhbvphPAGd4JTfS+bgEYm9M2kJl7g5QEHN2KBs6YMZ7jJAN05oG+BG46
/Ah/w9UXRd9Z2hidPoKrXLC67rQ34je2esjQwfxG84En2htZgXTRyTAZN+v/LhBDBS/Iyud5iy8W
TRBeWag75vqN1J1wNjH+mCVNbTV75ko3pimdzCcIVZuTi+uWvTs6w0geex/lLVKvgef/irS72vlq
51bjkh1my+CWBsHPq2rrn84jdOiP7n6yDzBhehQTKLTXVzJqN3itQe10FkFi3mjcUdbYETQmaayb
sJP0B3vVK5AN/E/r2Rspu/5MRBEIZj05a73XGDlOi2X4yuB556zynjabIZKXUdxV2mMgIz6H4naE
muCC3OL8nXzu81qBqRyQNHGujcOCZolCaIdqZxuj3WHnX4nfNFD0otV1HOo+/eOoMSPvtRY3B/IA
nNcvI6bc9mYuoVcA51LJ5O52hh6Uo6tljGhVr+mzNfo57nbm3liaTHp+KLj4DxgR3rm0UIOsIpvv
PMkJ0irU616xeueuxVPtA3Fp/RimWbi2x91aE7mroC59iSEQmS0QF+wUHfCeInPOZb5aNbFLm507
aNkJAkHbPGg2dCnyrW3z+K/cJAg3HLo7Rrs0SgWPfL9ytRTTVvCNGGHsNTdVjGYEI4EZ86IilZ+g
sgQTDO0wmsl4QEXFHYNnLx/aeYKljXYfggVgC09qfcttXjTVAzdBCCgaE31tBRlV4FlE9aamhBoc
7d/5+wUzR9czPrt0RwSn/7mIIiFRr6oHpj5iOGyXcwQmlOVxEucyv63OD3eJ7Jo8SewRnngok5ye
PzTrjijX69oHCxSXONtDuFR6guKJJxDaEv0T7c2o3Jvdhh/q63p2X6ISRb7kSpYS7ipzG64ycZtz
GEo78kgkWkiF2d3Xsy8gi48nr0kVh/YfaRFC01WvjIjZtaJAKnqd+L1ssEmyEco/XLEgMVFQugn1
9TSW1GEMiHdcyChRo4TdGp/WyaK7x+3kcBWSsfQKYUOZD9ilBx6nzAPwk/4rbDAM1k5q/3fkvaF5
AW7VaUBWiXkmwdGDa3w6p0RPnZ80P7rqadrFjiZEL8N+CSs0e8k1f7zFNSRSGdKuvSKUY8m+290u
XFMwOrZhlm9ZHdCWmD2+o6eHJ+MJQx9jasONkFkrItE4vW++cZbMatqzXomBzcdpNjq+64W+Zd7M
sHXfTtxIOO3znbACwj7tSFzVzuvs997nPtKk/zeRye4mb14rDY0UGt9tjxSOBLcw9zmSiRpGCxC3
9qdd0qwdhLaJyGbzle+r7ATDY0E5WKTfkyqZ+RJW290KwuY2CcqVqADp9klOOh02/09kOMHdtvlG
P8xQdycHZ1t0GJw1EdnWoqcZvgzqaAD53PHxebd6IO82CBOEaY9dMv3JarOxcICRxR0XB3k7icsP
HDStHc1HQsdJUzigJN4kLvBu0t1KcHREhUAv6LkAT2rBks8IVuGDbGuT4GcqxpcSrlyR10HvjuuQ
iLzp0VUjHw9Ifire2RSmE7/Cxb19E+36MMsWvR5yWsxhQEfXGvoN/JB7CAX8+0OWSpkDk1Tavni/
54s235ovByaIKWQVkqQGUKx1GkUy7N3kG9Uz1hTFL5f5ySUv33pcUVykU3i4CB5kKUOAxcubd4h7
Z7wNos83XbvtkYtIsnzVkW1oCVRNg8a611YVIQZpPIVWcRYq6e1dcc/cHUvbpx8K54lbzOFUcCAQ
osdCh6ohg7JeND8QwlpeLhAWMEx8XXeoq3CEdg4bRwWbt0tZic0H6uypzSoPxb0IAbazLAhq3PCe
SGWHQBGVGnMkOwki0etEfGnxXLGgD6AxLRgabcOMHcPGwfVNeqzn4J7YPs9+5eXAh1CPRnFiAuiB
7tHB5aut8gVhaG406so1CbtV+b3k2CopmlkwbeG2xfT37IOisJGjv+kf068VCQX2XXpnR0Q/32DQ
MzgULE/zu+6mWBgfISg6DRHRc1WIovpQ1DSLc0pS2yFKk824Anaa1Nn70l220DIkc9fwW/4sCy48
pxNT78dnjr7ciQVnbyl3MUE6GE6sswiMdtBypw7q8Co+TDfpSFm9f1ZwON5IuKb39PSJ79RgHpwp
IaV2xRKDlYA076Vy/q4UVuKzK61mqKDKF9Q2ghu5u8He6R18SbQrbv8Ldr1GaoeTv6bw66z9eGi6
uJ+cu1cpQtJmKFKF+qKMSaiBUhA+B77Sa6MeAcs0CdWFHbwzKHB8SBo7QsLFN17hjlmuJ+Jys/DJ
vJ78wtJp8XJG0NvwxWKsifMYq8USoc8FLsLpZWVHWNQ0ZHL9HIRcM8Z6DHcxCF8QumT0vKubOKhU
9lm8DsKkWzCjqy1WEQia1/hPrlyl3aiO60Mv1cc9xAtmchhth9iaEEeX1ZiYriT4tFsIJ5JD8QWY
1GyBAc1lgHZY9BjhXQUIMgHh1EILHwe+AT9rQc6gpDUU4yCzccFZTSJ6mUk9sTJI4WLpSavgRoO3
q8W8zYdP8xCKY37iE0L+svfuR7RYcxzxrLbfhtwunS6IAJ3Ne9cA3qrc18BstWlZm90dLAGw5YJK
1I2sdRXat9AmHV0WQnUsX3Md1LKmFoLZ+hqhNMeFNsLyswjN4ab+aDPfyXRgZf95FJ7+0ASdJk7K
HLWAAY4818ONdaDOtQYvUxBumv0g8j6kRFYL9eokbgea7ceKAAbawoKDpg+Wr/3++qVyyWU5C+20
y7QcQNEZ1pRB4Uz+fFO70RPbwIV8feihdy7SwvvL9hsaJ1L8FicYvuRgREH9TD3CjZs2iOEfW3/N
VT28784rAL1wm0cd+Gn4i93nQBglcEqXQi6n9xwW6R7w4EyIiDsa+3V7/wXCggPqb9c1IGGb+wTp
WLc1GmhRKOiyDU/heXkDjhO2HO4n8tXv+/ci8o7dMzLuIBpB1AdhQsRWuXcRVi9hSKWHG+AUxV4V
C5m8PLYUZ3dwrPpCGVjc+Hd2piMFDjhgM7qNDe/AMCcLYicQNZc55M1CAKoFm+8u+xJIwd+5TpVe
gjIzY+8251tS1zst+4fLaheOWqfY+Ri48fuNe1ohCVmdrdsB6Vu6qIlboIpXpoCseepJSQWjHo3s
8pvQsgtBcoOoY8DTGcx+lwgBNatZe8fIxoB5MeWM6wyx802ukQOZwijUwO32MRYrUHVRblLjMRqw
/vKqbfrk814GKd4p+11niYPT+FJQeoRbL53CRzJXADDon6YINjNwaGobP1b2BSZIFVRK6tXLVkZO
rtxp31gjYO6hDLHKKEec7wL9UxGRD72yYUoBuJNwLa4JYa7p/uqZX88bxcc8rC6jO60TRFUWjx+u
g1W+L4f+9uMu7pNKBcsEPH2CmuQf79aySdQvMYMvVQd77I3xxEgKDvl009VXGBQvZvAcYxSI66Xp
lpwDyrQwlkdRMjoykxTRhGSfpjqZr/M33UidgNgv9ZEsZhJMwwFuGa0AkzJ393ZswJGwqP+ekJZn
BvEB/RfvhZhRmZW9md/3DgoJxAlxlB4b4Mzjw7bFfnzVWVPfLvGnRM/5Qdp38MIzHZ7f5NYQsjoL
kLk7o9qYrd0+KCiZPmCfE+elzJT5bdGiOKpEwtEGcMXi/7vGspKgZR5fS/rW/8acwIDCZWsoN2IE
cHRwEezG8mEXCBd4Bs7M/Z3WKuIgZkzKPVIOjSV8Uf4IdV96r/xffjjdcTLkF+GDBQ68SxIxW2iP
6NIShCi54x464eKEGzhFaMBTIOl+YIFChRxyLC4sw56i0DsHadBcKz9ne4erGsPN080dd5r30jG5
9QOcpElvMi4HigIoDjeRMU/wmWnPrKapr24y4n/6YKfKHOIByNBRqkiQbMVPNv5rPXTCcDVye2Xh
Yrf7tgP/GGb64TVAxI7u8eypTI4Rg9D13QW42KGOHz8QolQJxziqhYQiQ4nJlxPF/dIFZiDzsHGu
PilpysTSuKAedaj86avTV978LZMFvn0L6O0QQlXJjczkFea+5sDy+1uueSfWSEFzftB+y8Of5cHY
V/4MNRwbiAV23fKDYaM0Zx8Lzuy1+5nNSo+LyosDRFpUyuPGNsodjSLzKLNM6h11JK2jZNIAStyk
ON1VuYohyEJHmes2BxplJ5tKutybtcXqGAqHJDBmLLHt7T5IhSl7U7X/WaoqkNqbXcgx4YWh8znK
t4qq/3CwElCNUPs0vXVVlExlOAAGNv1C3lAh+dDgR72jsxDNhXDth1GYAL9zz1Io4C+iN+DrLtO6
VpUOFAncQUz9bv6QBWpz52pNC85D0QS4YWvdDUQwZBcSJdgrYX99E+USAudqWeamqOXyIjuYxVGd
WuEJuPpHAd5UimMQOGDsysANsJl0qiMT+h4R1vMA6rGUW/6Fa2iI/C0ir3NGLJWr7FarU1lMbeCP
KftR6ickBOz+rPtth3jsDMb2zlqcD3hDqr4tNz/Nb8rrGZoCXqWRxJprLmnetC+uPwXzL7Vw5zYM
klUxNXE1Uu9ad57VhntCEg3FXVqTWr/S2WsUGdp/h0ZSlFTS1Qe451lUJ8SskCTPm7Rc8TXJ2tKw
VaIx+1hUoo+ByOpCs6eOeZEeG6XYTUQIdd9cQBZlWWIrnpUkeenISB3LfNqKs8Gx4flR6rHpNAMP
mN1aTfPkW82cT5liaogQtm1/xC0hdUmRyNrbzjxVSVAquEzD+MMLbA0gGHcmCBUY3A3NRapxy8/n
Bt5qqCu15UXAKosMSkVsXKKxqZvxdQqsSkEPRjJZTEKCZQuAJmE79Px4WDQS/yJS3EpqZbT6vbxy
ilPt0q5LsYi1wDiImrOTOTmQln0Dov3JYaYbhVqournjHCK/XUFVUg1mpJm0s9rUWRK4bGw6YxAO
/1vOrxEHExT+5PSumOVayRvHc0yYe6EtuIPt5/NmNNZk6aqImCwtWr9GidsRswM7+ZM0Eqh1qUxo
mLo6OtZ1zSM+PlxC7ltJjJoIH93W4xjT0STgyMb24SiKS7lDD8UnlDB8A0XZcVdEPCkiQ8uNtio1
SOrp/NOrhlDHCr0HuYGjozNSzMto2ErLe7KiYP3HtfeAbCMFHss+Ac4NNjj4U7GBmDWiwW5CDS82
eUObi3yqEIjBMIUkt/A/eSK/Q28mdjqCvRB/Q119pfUPACD+lWlxRaFXCJJr7Zwtc2DKcJgAL6Wc
B7DlicTASs9L67oD9hnPw5GJuMpbBUojDgGnMh0GGGGwF81Bnq2gpf2j8OcqJN1MsTfwq81Pev7H
GOPsBjAEeo1zeAa5LrXMAHYsrizpvEVmoWc4TQVOy3IWhVCym97AM9bAik2aKn5i3GobWcIl3UHc
sQ9XcFTNO2CZKjmOhSbD5E4lEnPLbqG1ajXnE/LEdMY35vsVcU/zpi6CBz7tmf8UxtcbTPfnLhG7
PEomJSsChMqsscuLIE88fNGVlEH9uLUoZBN2qWuYChOnrugm/MZ0QZ6Nz9joqYZmT68a6xhG+K4O
fJvt5TA+5L+HAedtbQblIG2yoeLX3u7D2OGUtth34LTgkZyiUyKj2B3mzJCTmFBnReutWCYmUDUS
DK0/wzQRj2pVEE3itQMWL1POfAwaz/kN4t8FdlIG3zfnZM/xkzlDOxLVSfgaYZNSWIM9f8fAlwvn
skkqFoBeRrRbPVQoPsjNQl37yQk5moRgefrmAVyRxrJPuJkHkyVv6ee0svWgF5Vqo8AdTuRxTcyR
QKJgYUXxsYz2fvXCySzukumsFHGqInQAt/nl8mq07/ZQUse+YB63FcUNpC4z942Z92TTK8/1DAzM
4ycLyjCjk45OemUD1PDxEhYu7H9iZMS8fryOTxcsUlhk1n83nmZyWS7fVsGFO79Dl92GZqY9hRy2
LaiePbO7Q+15vvrQB+MobnZ+xfXGccFTzsiMPrJWSSNHYrBPTW2OXZq93g+PSo+7YOQhNet+KhjQ
vqbdb17zyNzuAZMV4MINaMm7vumFUpjKaBf4L94PdvLbfsIlGhjo4TyPhU3ZhfLVosw4C/h4xn0s
Ly2E07zJri5kP5m/gtO1qwFFBaxRS9uuxCiXJKgo83sRUaiiK7YbQkfY8OJEL08SPUEtNs3sJw5i
RD2TXd+YSIV+ll73pmWkz4x9Z+8YumDgA+8eHCw+q0HnfGIW90ttfeK6HtZg25vNSkTzAmwuFt2C
2b1F1vvFFUykvkg9nC4Vo0o4ELOTnVE3ts0TZ00BsIxqZoGVWPfD+xKgVyshv2Zn7l83XNZK3znw
HyMdjb+m+5tEIrPYmDcM7vLEa3tEeXm4YG9iJNL1qva+ZKV/x89qVjm6Mv2CeFsPtV9u24r683dT
e7mtlFXo8ai4rQuHv4rKtVLsxj2yewVLdOHjhjY4OAYY4vxqeV5q2lP6r6zPb61g3VKHqbyV0Etz
JsadmECM+yPQ7DGzlQlJqwDCMw5sCtse98kB7SncfVHbVkyXrxXPoQ0mI9i4U6fNHL/0h1f8k2Ty
mArYEEeArVDoDjscOSmHFRhMvqMLn1ZoqoF2j+m3iYg0/E20/0LihuUf7Sar146W8WS0DmKl98vY
6SUHcyRfWOW9Solny/np7vrq70fb4o1DAGajQaqA5tZXjXydLEnhFa+2emePdWb2XRj3+aj7yRPO
LN+heq6Rbc3rEifQ5Q0Bds1g5ZC6OiXR78XxvkN/8wCsgaDTqASm8SeJErhRU+sQ0lgzQ+9gno5T
V9g6vRj3mbRwKPewPXrfEWd9dpw/9e6gspodzl9xK6GCgRIWRV49W+2zvLg0CyUfC8szy06XxGZo
81IzsND0MB1HcF5HzmgxfgxkRhZSH5EYhtWCfWvTKWcTPJPJQ8pvecV+kn/lOhHYuB+XihaE41S0
w4gcJf//hhOEEsAXqci/ZRixU/6BCpvnC+/JONlUxmsAIAY4heMtStPe8eX0eNaT+ZpNvDHh0nfv
+rV4+4QYM2fmapoH6tQR3aKRMyvQ2XmXLmC18SHPUWek025IzGVGf0mtwh8Ubu7evNKAhRf3r+Db
WM7mceE5DbatOUXwQ6BMlPB5wSgzW0Aj4QZ1SC68b7gCtgKVN2+UXh9nhUmzjnM6CLk6SqmkXtst
pjbBRtaHdmaE3or1xliA3DJyJpFj0FeiNgTM4WgBLtcnVLywftaWGnfUw5g8hFHgNIz489fP1NUj
7fzhaQ5FdywyxUoAzjCk9VBjJWwWkaGSbRYXqaY+pMKnj8P7VYGJPznaXBDs8fxWz3BrcGbIKdHb
QQN5GFt9uPJW8dcUCzEgNXXl8/CxkLvuNUsFXK8FHwQup5biano5vBmC/Nx7WaENZOUhNWcwujTx
Egyh9RUfKJ0EzQNZMdvgJafcqoL2lJYwDjqT+m+s8pzDeJssus5Pq4wjIATnU8AQmjXWRE/e6m5U
x9SZpoTHwwhdHxKulFWvnIdQ7v0PLoyE4rQL4jyRlk90/MHzDTdBvAAqJ7IEdYNxHK6CCvVqPHnr
ULIjQ6pMdljD8oYp6YBdkIxPuxJXUOFBs9XWhOpKWeKZCsqEqgDoG2TOZdFOTwLcd7Lj2te33XqY
fMArEmA4dtOapZnU0FOygLbtJre2MP9suvJMQNoHcSOwx2o3zqZRqdWUWvfONdEglT5/ocxp0rjo
p3wnf308IR5/iLjhG4oHrPCqPtDFx1aYfBI+himv+tESvR9BIb1VNVTrCB7Q7Nnd3itFZQYitwA4
p4PN9CGhv8e6+jP+TjkAVl6uMSnHne+aRTjDxlj4YYghMnuAjQK6wVAaJyKpZJ6S/s2P+Rd37x9+
4hg5s+ZFVdEy4BJElAnTQqvnLErvPSB1Zu2tifmQYYemT2KjjS2XWKB3aeOhaI7tAgOZZ8rYUyU2
Bs2NC06e/E3I5VlwoU5hWh0j3qT47EyuBETEesuYlaf1IKozLcLQYgV+ri1Vyqu3wrwebtyrnt/Q
b6lXRRPsxwdHoEFxHdEyh4h2DMhnLEnmEmMWbilavDyA6rC8l/ppoBnwTGtbh32UIR2aCMh/rEe5
ZnYud/LFeIc3IcjCSrX4jJMrPTMoDrUWXFHQf6zFuF59Dd/tTxkimkWUijnzQAN73qOQBvVEjSpo
RKNhaatwt9DaseWJ+oH1iYm0u0onyNGZ+HZmaeUDClH9rKPs7HZN+XtWDFr9E8taI0bhXcyw1ruc
CDJ0tLODxqga6epYBRxdfl7OKS7LT8hDQcqmwWpK2el9y5I5YLRFJ8hr4gBtYJXNSOOG9srSzt5f
H4OwGIZdF9wzjFQPYtxUoq+0llOoF/+HBaiSq9D87Pf1gIcJBW9QjW8inXa26AJRyHfGNMcBVjkK
vpCgJ6wfja81PVQzXRXVCJxYI0rPxL6IosfTTU8IZZn+9olf+wgibZGdR1Gp86VbmCZk5muBAIMt
3iei52L3sEMIK2SXT3Plt+6ZLrb4x9grGcHfbBITRhjjMm6ne7yQk0rhJJHgrWnTek8x7By8bQ9U
rzSqH+p+5gWvGGDzmt29D/zTXMgO2ZYCaQ/NNZhXE2mXB7RBYuEWqonAUKloBYT6G5Tp6+Z3PKkg
kh4Y7Uj4vTcO8i+4wiWSh1sCC8O+7/uDidsEsLd9U9PgqaXAYOUtQd6EYi8MsTrFUFBoT/Cd92dH
OoX+ZuDtpFifquHTM1HfCXA+RxZQyj0fSNF4bCPj79lsW6mbq5bY9IGLVoymAgAzRe+mbnlIIXEK
4GKSaKMRYOGbnTE9LeamKTivxWkb4I3GQuSZUayJf5V0bYbXKBD0sKLjIHn2aDgEB733i+kVdTz/
uOhc6Guvfz7vrwOmLYAp+X0btvoVsa67CM6Nh4WwgZ6yT1c/QwP6Q9+pg/XTZ4Ykvhf9goYrN4Vc
xssjONHDsNCP/mbk44imTmS5kva303YnTHmOcywy36qKEn7V54Kf/xT9Bhy20zHPUiLs8zbWbTon
FXtLLXMTUISXkNg380ktLPaHDq90vQEb8AtHPdSb+DmWgExFLXd2tPuwKSfJRtlEUrIzwI/wH4Hp
bU0fwG4xHAZpn9yj18jVeOA+s+Pz99yLU6bOEtqKaaBpaziYT/6GpBwBpShh+i/g5cR4CephB06/
ZJiLusHHb16QkuTNw8uvh7NAX1mKOsZo0blUIREBdG0JfN0X29PXMLtHLuafXYUTRWufzwO2U9BD
ig96u5MddMk5P4RUIa67GPWwSqoUvXaAzeETl3Kso9upV+OezdigSGi7e5RQ6+a8Wb448niYNwPP
p2aZUI3+YdajPfW71ndxVZT51uX0PexXTSK9LhDHkWhRHb7HHDxmmpcAhvMJA41yqV3tYRE1vq/3
90tGpkQYOPvBog+KTB7tCftZeZy2hcxuiVK4a+IaCZue4fCQi2HAdL+hdAqjeiDFTl8rLPVKmACh
ogns7QAC7AiuXSI4ZSEsyz8mUPt65XQTiqGaFpgCDhWPwUc8DT32ocv9/qhVb8O6JL0DyGLzrFjq
cQk3hAgJrKFprELrSX7IPP+Nly6wH1/Pnaq/G25m0zkyoQ2u1GFHiuDQgROhKlqPBp/ZeJVR8/OL
mTixMQyw1Nw+IcE2Ai9i2pNgKwq0v1HhGQuKadbmgxaQGKz/ToFgFImgWKGtuRI0gqWMJ74A7XNf
1rLNY6QvA4UWr8ODBuiCrsVrXSFAsVWlWzJVL1ngAHGcIr+fiq8ZfB1ukHIEmGqdJMT0t0ge6XMg
SrNGqgdTdnuCgIAR30F7K1P+5SD2TehlpD0y9ahFD+Q0PaffIXPrQGShrlgE6AG0AcFhhB9xdkLX
yX8LiylOeKyYcoMoIyvuRaO8qT5AYGwSqsIlZwEEMv4+Nza3DoUQF1zyjDwKUvog/1/AMa8WOvD2
mxUB3j7eREOgRoZXnc/yAle7wUrnjPC5rt5XlMFB9NygaH8vuzc65zvu+JThETpIETprAoSjNVsk
YmecgCQGBKVnONOWutyx8/lw4jdu5mzkzD+D0lsoaKq974lO1LyijM1NnQ9jaR95tlDOp9NLPVJG
VfoUYYaeHjPOWUPtZAUmoNDbSbBJgQXtZttPjyM0EmK380QVeY6XyBhuYhZanRBbDP+qvTMp5YP8
LrNkX/X5w9g1tlctVWmX3HPrk2gddR0PpgoP0r25zxXgNl+sgjt7YNJNwIaMIdJWAF+0HtkNduvm
jO2fcouSsZMhfp+haH7028pnFyQQBJc1dtEtAAPYTKi+vjGNee5Rfviq57snLvnJ1ueqHV9vOuSs
6DnjoEHaGtjTm46QNxuE4pmZjhaI/LT4lgYGlN3wLKe6v+3dl15D5IqHcnaOANHq5UKHyWYY1Fsd
jQ8ko+UrM4PxNvygrVqXfL0+2oDmzPkkJqSZqDPI/n+xTvHsRQ4kjM5eRvR7HsiqxW7f55vOhqvR
WkKPIK/4sqxO/TGKcXfB6ayDFJBWzlHNBSg51pmbA5heI3ReY9+fHUieb8S/Jlz2BHSiFypz3iO4
NDicmn+i0u4AEw1mQevMY3LoJ37HrQjMP9csmK8Z41P75jc8b+qu175iG+yuB/9Qd+UH30iRnAxP
dYSYI1FhsjG5xM4fpQC/mmL4J8uUbL+yu4IWOu7MXRj1Iw7MDgkYTdFWS9LL4spbwmOQ0X7EfImS
qLSv7kENKlG/B7P4ptZMsL1MfBMyHqmd6Pg6quPpLwa92sHP9xXHSq3Y+JKXd2832hisbu/DEOKD
RqrSHUViEwRgbn7vEKY/l2ZK2ueRfHaT/gNWXTai9J644T/VAGVBzyaFEcIehR1BmQzxORMZCFGx
W5/n+CvDsO/CO2rAjB5D5fFN2m8M+pCE/ZNe+7xjxA4/7G6zn2h0qwYAOdTekfb1mDcZuwA59O7i
ogCvO1TFGg+Shp9xdI0tI/6c9yFf7a8fRc8mgEMNBxv22hSESRI+ZxU4yHrI0ZPc0WK3ap+dqXMg
NohYNj7IW3G+CNqhzp01XAaaVmePMiracR1LyCrPANHg4VwNYtJIyLDlnZZesfj6mX7eF3DN3reV
rudx+DpKhsvAVnFmvNmL5yKojFH6bYvJelV5/ykmvRLG4dDJScYR4GKmx13ZDHRG3ZuAqKEbwnY2
Ru6dtYu95Z/+fUm4F27xCMz1C2ZcEGaiWRWGds9U/dF+/dO9q6YYjGTQMCoHnsnBlhkxRjhjIxn/
p+IKJKirwEHAIvFeyojpjp1BJY/kuR6lKXhF94LwJrEXw/hh7RJtz/CrmGu0nnQHMLYsiC0lFp0w
S04utc4Z7nyZSqolvizMxUQhnZUw/m18nWeWK5crafLfX4jB6zQdCBJjI4qvLxUYRbJeDfGsWVDf
r/+NwJyv5UR2Ua8z9nvFQJvimTuw+XVotJcVPmQugwT0tuAY96C72t7Zq3Y7wLdY/BxOXPRfVvpk
bRL9kegthmcwPdTFMb0yifc+9cZPcfML6+gRbRBKI4csICVXt3gurRJrV8ZWo3jslVBY6sIm1j26
ynU6eKQEZ2tFt8l2Z86020fbuipgXBqYQDTv0Ci0Upe5HXv5VTuaVZMZPib6djgeHfe39OEDEt4F
GHZ989T4RwfgBza0I+Zpr8fsRUHRJr4QXiFBj1eG88Ea3QT17HabecP0m13sWM2Gus8moD0Ue0pU
Rb4wvcuvumnISLdjJj13Rr6TFizFY8ObpuNt8wYAVWxII+Ajz3crHxOMt61Zidq4gRHUIP0J2Ckr
38WzKtxfJR+rXQO+hf4faxb77yrKXb2bPqLWeZVCk3CNqhQYbGTsq331mIftVy/L9CY1ocRzop7n
1nnM3rXDTCQTXx30XRyhjC2S/RcufAgPQUzH0yEtEae4sSFf89zJf4AFpPwy/AsfY1Kw3E+nZdLc
uKfShdJUi+sxV39FdeGOyGiHUlBKpZtdUO6mDFPqS23gVPcRtiozadNRgoUOGtMbAPdmdjzPUHOp
uXMoLD/GeaV+yoCBlOg/M4jID4ZDJFlEJeZd+W/sy0raIcGhoHqsz3zLcpqgFhWJKqqMRYHP2rt8
+z58cwiEoSRbYLpGAsWi6bnQTfPJlrfKquJA4XtY5Rqer+aK9JbKPFfLqOsnkNRMyQLVz2Zct+sS
E5XqO3a3Y1ezHclgPaviK3TqUXnyAH6L5tM6AyxPZcAAQQW4fTu1l8Uo+MdGh6EZRYVEcKtxW7mZ
119vzww+1dqc4WgHSY8HqkiwTj2rP123553L22lp3l4HiSyUEi1szoxGGL020idEoPyFa6C3dk8m
gbjuO+kSNgbKAuvFHGyTF93Sh1QAlKZ5rbHhwTD4FN1O6C8fKW+B/URVZK3bCXOX1Xenc/3T3XF6
SXUGYDDyJtz8/C+szNSsUlebhgeu946+Y50IU5sy+2zrL4Uik7mwJ9T+qjl9Kywv1owGabenVw6V
WWrNbMkt6pRyoXT4wr8ATItSrl3nrwBdj9Wp60B4HAFD32eFV+MEvQwlCizhW2R7aDkmdVjlNPSw
n9PlQzW5TF8yC+O1Vue55A8zk6KsvDdxLloJTnuqYNTHTSnaPcwPedMSTW/E8jccd97C77x0en02
NHWOTGYtmG02spo3NOSQkPuqjomXJuZqWh2YoXylK0ro3+PRlQ7SLXGShzg3fm+b6FA7sKl7LLBW
GVaI5QzTol4pEhFAbZBq2HEtHrRfDxkhKCpdOMLbIJC9Wr7Sptuy5dq/NVwOZnrsA7Ap5dlXdK4b
xCB3GkFZRwtm8JOveQLDk7jXLtHQoVftr0wAyypdmePRRrlsXg/FJoZDr34PtG4r9d1E+L/3/v3f
jQB/+gUpeGthPHOZ7i5eIQpQ60BaNHzJQsBEckSU5oue14InKKF4qS922YRDON7C9MK7AUKLJ3gf
PGz2GwjMl2kMWxkmyuV/sYbVxA4rucJB4JV6tuTkeR99lwhy+Ior29LZ42ix6aQvqKifabI82TPe
Z5O0HS3ENadk+kBzmrVzlG2xWC3jMQWSK9kuHVS48NcZSV/PU2dlcwdnm99FS1bnLZv1P1pqq/Wv
VCjwjIwfsEzksNPXLSmvbTGrPu5KIGSyt8NLQqzvABN/3z6QsCc4awBggQxdYxk5JXpgj7H+XrZW
YVFNVguKluV6zmtOycTz2+9WPyu4RfVK4EFfJlQFu4ikQAYbpwqSMTICNcJOmDwf5R7ymZSNb/NN
uDKQstqVefihU0ZcSN3+tV4t7tcxI64f49SYDbPMOnhWh0w4RHfeD+bYBcy4u2sSdlBQoiePwzb9
g2hTqA5AHE/lxgvlTj132ie/fMlruALztODYiS47SFsv/XsAGAxmo5vm7qhNOtFPzdCECd/URoM8
p0LV+zMzB7gAnmq1WvTQficDTC7JCYtP6daFHT5LuRihu8nfsnKMuBMliWEvxcOO4smk7agKSN/n
m6eiD3ixtEohmNhK+T/rIbCozSlXlGdetophbIP0ATmjmBYe5DtMn4Zg5Uq+bzo7mUioEhoLR1h9
OAGri3ceEPYqenxdvZbEICapzWEZHL8/dabR439JkSJWnHUkC4hI6EW7qyIEDFuJV8frMSU6D3sf
ssoXx/nVvI4b3v8F5fhMMFCE/Ly2NueI4E3fz9FhxAnxlZjEwkSHrrzuFqSlrKHXjPLR6L1bImcu
Tw3EC5jEeKMopdumZig2q3f3HwzNPuYozLnYRkcTKa5htPswxtk7DIV/pzaKPwqZ3LgqOejEAm5Z
r5VI14+1+cW0VpCIob08ebctyJ/2ukbcAy4HwV58PQg39Ivbr5/DahlBW78b4OJ/H/K9T0RqlrvO
KzsDZiYeN3dFUBCPg1hapaXBhv1rYZv6p+iJ+idMpobylwGcgM/b/Mj86J8pGfn1Dh2PjtSsV1Jr
eBSrusQK02n1Py3lrCMlq3hXaZSx9S2cowpFKcq9RgyaUw4aGT+1Z2uASp0JHsUDQ+QMeCpyFsb9
5PrIj5npgefkPxoJ+WWbNCDnhHLIHD57qWc70disNATT3cd/Qm5uXjsdZAE7MkHRRG5w0fUZ9Miv
Q1CeMHel6FJO2CqDOnn/2E2haGOorgwOVLznsfANxI3ooMV4/sTMJ74ZtvKdj/iGlqQfDY+UiqAe
JEfKYZ7PsWvuOJ/T13KQ6K6hE4Y2PGhRqFzgBJ/45NXGUn6nfbMMQiFsu4e3I7AcbeG5QU8ieCLb
Gjt4mIvt145vTLjdCUP6U/EXmP3x1DUyFne89Gld2aN9JNYv9/xVgsyGGDKqhR/WwhSqaloZeCcY
hWD1hV18AFJpcOVn/5ei2GWCK3tDL2j2xq/BuFUSbL85ew/X6iPEP0uB3cXsTtA0jUXBjj/d+tz0
i6ZWl+9hUW5cuT64TkbupAGQTORkhAPyYmYlF4mvhyU0xuUrAQWMeHmNqujWU1CKguU5hcK/c5a9
zybpGdg5fqUjQ7d+8x3JuPo6LESk2vr3cIGaboEGzDekaywiaXa2x9160+FOu+1Wk+DonQPWakml
zXrEWiH4fnXP/mMQaWr66uK9buIoFG2WL0KOM5ninI1+QzumWODMKqBuY45obXM1IGDnpJkX1aUB
oHzzPJCrWEAf1YkBnuhoGguVELG5M6x3rhAthyxODx9AtazLTrpYuP8fPtq+HsTUrtpHwMhXeJo4
HGzWPDGWbfGqJcSo3y0Fl7q2MWeCRk/IcLoXa+BXYcxGOJY98kTH3Atxx9ImSSrUL9EJ32KnIyeZ
cqUeONk4GlHJFcoPPBoWMUXR+T9+m6Yc8xzVx2mjn9m7WgtDaS2etSpe3pQXdTayJJpvzPQF/KxM
jbObcU1C+BR1oB5qoWjwlKqPb+30WzhvdWL5R7I/VMQTuXW7Z1QVqQaiFdam1+UFU/kzr4PuddO/
PKoeqJ9C7XnrlUq5ATccRieoQmH08f+enfqATK8JGjAAIcrUIe6Fo75cByssRSekGHwObqLENqHy
Aa1yrLllVg6PWNaBF3tz9MSrKJDToezj1/3wglJrIksFZun9+JO7TyYreTK9ga8aNsOdPk5JTMXH
bhgiGZok8RBAOKc3o1mxOPxrjkVmSXD1nY70OiJSBlXqMWwxZNxTEw5EUpWjkc3urozYv1VpPGgj
sKAlWKUIsIYC7zMJ8+0ccH6WbRmGooXHl7StKT2Xymc9UrmtpQ6Q97ZxOahcP1udSTR44nsfEsH5
8JAq6LPCklDQ0GM8fupAknA+kKbWwv6YNim96SUq+rjMs2dMSkK0FkUNYZlVLV75UtGUOszlkTtz
Jg9iNyw/IJdrpAlACNc4VqnI1BveF2LsGiooh0BBcF0yW7mWIB7GL4ywJKk3xdC471HTAq9GGxL9
Am3MOl1rhbWV8F0q4Ygi/UA7xWAkazT1jo5NjyuPsPmMJKuSbJIcsc9hWbDyCNc4Hl+nnycSdZIK
s5LZMTcoY11kgS1lXypB9cqfxV9UAMOKPLc1efKbK3yE0jXTlbosrhOEJC0Tl8q9NPgviB76NoyY
HMAYFPIDNkN5xnjSwa+IY8d3L2MUR7bn8uR2+657p3T2awlHRFzIOHVIFcvpK/0FM1Z+bNs+wjUX
/Gf3GYFMebOGW9ar8oBd2Vmo48/V15vNBNXDaDOTObi1XQgC3j0iWT/mAkWuvwdDqjN1l1RDfhnq
yJPzaKwMblksvTpkJKwXfiEnCgSf1tRVukNGPuhA7qru2UH1BefJsKpeiHeVD8rNnOdWeHMSt34Y
gXy63N1Y418B8ZoLJCrq5lsRXtw+v6YtbPOHS6v2zTHYPeTezFJY5ljJ3S30U7Vg1cntwcYKjeRO
s8ENUay9NpNNktlT8P/G31t9XBVGooLrF7IurW2DGAT4g00FBtGidECQ+eVS3SfNLaxGPD6EEgpe
EVw/cVj0kKpcNx9lG5QSeVz6bImb7MzjSIfuUwnfwpo16pMuCGwMT1fcTFPPP135Aoy/PMepgC6v
r6jYTtau0PWXQiCst/lf3OBEjhifnVRF+xk9X565LInCUbeLzWfmHp0wRi3sHfWZMucCdNCQrhNl
TRKNuPRk/9oyG/QSUiN2tekt6nl21+BQbd8LrSerHO/12mUZlcZNDBSIN2d5nmbsCLm+EAitSzLD
3hE7Kqx65457x/j9/sglSWbMxeU3fNpJ0sutp27KDjGmO6JDIfNbrVUMFStmfQSuPb6Kt3QVoYLt
BNhSc23Wu7wJQNvhmd1BXAJ2bpttRQ8wR29IL2z/uDtloHEUkdLD/nBRTbcsUKX3E5FKbW5iRmmd
KG5b1X3s115R9aHyDStdSV/vNCeQ/CxwuwbbDnOAZtNgC6zw4+bjdW98Z6buXJ/d5NpBY3anYbEU
6/CSBcG/dorfC9T4vzl8tV+eKstcVY3RqH5mgvt96LRLr5ZK9o5xQ6MAiRD4gHFTFNIDzZR+jNlO
Zo/kGrh6us6osMmo2TMijSA7z/hX2R/sETPDwZ0w6Ms9hz9B34OWmDIj8aZ5WowmclJWUaLcvF3g
D8AWhAFvHhChBOQiIkFfREPhqtT+kWbasSRMUjKBag7uDjVOYAZ+BAXho3DbDu/y3LE3PmlX6xRO
VaIiR5a6yLuXuv/queQ7FGjwjnv5ngC4SSZo1y8/9lD37Ozed5D6kyNfFtTTOkPi6K0wTQWagman
aLpnl1xlWbXdhNyYfvlk/jj8C9nDpjP7CiEua1gPnGe9ek/SwtJH+04qgpSwNzFYHKVQxEh5H5zr
xuGztzZw024dOl0uKJZUPSdF3AMn5LZmURfq3u8uJ5ynUr8NCW9QGj9L7Ucnf0DWSz53NvAzc4Dn
OLfGBrwhcpJq6ucBtm3BFszrfeiDzwymDz8EyNqgFME7+qgDishtvUcPOtV9H3hIFPP4Z5evEsI5
0qyX47La8gEDHztp+jmWsly5kiA+dNgriQPQTHDxXpKFcLAti+v3aUZEstkaLh7qLXCmdLg/YVDN
lKWtLjB2l+1XFVEA4y/RM7p47ICl4BpZZYiPoZgzfVBIX/icDPzxMIUqHciVnbwRqZWkCAdZvfFP
YXB8DhFV91EJxhsDFUyaQ7R0zYFGiZ95616zebMCw2Z7o1SYSw+vJ6CpHY7e01avOWioCkiyyB+g
oMdfvhPrngcD+AfAw6cceI91ncgtiJfcRofKLQBTgrjCKOgmGs8PEV23Oh+1nl3Y03ys/vlhRGKY
E9cXyXHMJt9vrfiyP6H2g0JOyADtsbMQoTekF9KLpmskheOLSLA723GzvHk1fio+dvYHEPrndbFI
R36xRyeaGM9Gjn80VxAeBvgGOTIFYRSJbQS+gASofCeqpxCO3WZDHH0NUZKA8taca0gAZxVLRsX0
RytQ8Jy3C+Ft8rycsOA0HxKaMcEUnqHaiU1ZtxllWK6Fc9y9AmPyrrYHjA2NTOMG1acEDVJd/dbf
cjl9sQBaiS+DykKQpPeEcxtuvcdQlXVcRAQmhf/rwe7gyKsVBDdtOPsDRPA5GnqevWx4O8ug6Ypr
rfDYGy32kSazmWIedVvgwtR/C/N1lu5BWi2x71g3lHTrOWYLqN1wUMfSpP8Tue0W8o7ckg4TDCYC
zhbuMxh2ZCcw7kAnFeLIetSul96j/O4ziQmmfA2NIQkIrgbAvFfX1PVSw78yymvNQI61RrLY4sO+
KvF4WFh6mkCKpKBIXVrmm+MnUbObP/qHHsdnB5+QtgL3mMC6jBTOsKOv946bg+oPNCABhZV3BcxG
ZE7TL58etwj0X9pY92Qeu61T6enQzjGlzgp4ikrr0VNcfzkUjenzO/6+1IeXhAXedistuFIbkBl3
DL68V+60+z4O9YjbIXxDNfE8XJAgexMi3yjvVSUxmRYuatOIeSLJhihyNNH4W/i9cvluzNvgmpvT
/55g3zZDkJG+XiGVwIO7Q0Dc9DrGUvzYag+B1wkfG/GAUdAmZplBexWA/qLFsFNQmOBZtVVfBIfl
P9v8IWWpVZU+I6xtNGC23Kv41l/CYGUkxV+GRbM/Oi2cODywGYKIpB0jvkX8jlPnFwUyNh0Vhuci
jJqfWrFioBjHQoDn2dt9y4gbRQHzaLmV33lbr/0gXSHNluTADRkXgGg7n6va7QBwKlEjkfq5T2bB
z9Q6LciHOcNnP1rNJ4kXQvEXWq2zuyScQMGaCocG78b25HeF+8NMWzTG7ALO8zW3JD5RVOuXAmxR
BcvQU0obTo99KEXEFaMu2YKQX88dA7OWtnp6sGVTVstA3qSaGCcGbbKTzt8naUt9r/y3QuCD9YMq
fcZOW1pK2Luc/6mKncUOZz2+IIFVdsk/QrvMo3HFmJhuO8OUPC8UiMWanjwNemhS1mG6BlEcTU2a
dMm61Y0wfET2CDD1p3MbgsWANT+sNmQeE5/l5blerSAi/nLkIQkZPsRqFg081zYu6NXPyOjk8huy
ZF0/Vtvj/HX4okV82NyVezobCjPWptLCQ70JueNW0LyXfXoNnY2I49+6KMx77/dnhkhqxygGq/F/
PlJXkO/m2F6VhUXdrAH2K5Qr5t+moG6eKeL/FYVr4s3P+2bttQX7HFaWYfrb4qWvxVVFGLxlLXOv
5wuvxSWsstuygYI6EKIoMkio5+Edkn2LWtJi9D5Brh94xK59mulJO/Hx7ZB5q5Hg8ooI60qVXIFS
s31U5UsFkvO1/bXxYK3gt6SwKNdlzsvq98+TLWUeYsGHp0tiVULNek7vGEv60VScjJxUNANgJWrY
Qhk8vgkIkR3Lbui7JpkAoYUWymSL5Tq57BepIaEJewjcJWLL5xBVzrIl/JiYz48uf8vHh1qkl9xK
1YUYlpCU5Rqy0pswgEwogzCht5t8f9aIqt1irHtvroz7y3rqQQvU/sJYNSBekF8QTKUn8XJKZr0G
4KscnMhKlnsqjqzM1Awa7Jzb0idx30bJTYTLa9+O43qDQvyl0ddp833ZYb1V8YiuT2IBHCqzVq3C
RuFTOO55Aw4IVurkj9Qpl+bKAfu+botnG6GQlvWqxt+Y6iL9+lrbJ3bnYsixePiJxPntEFlF41qd
+R4f4LTESvC+89WKv1K+PNYMfe635HgBWd3T/fe9S4nEbo6V3/fI5soSmDckRvRdbmjPBqthsmQY
JLjzaeG3o7c2tFvuYpqAErmAaIVHav0fuLRGQWzZyxPVzQk3OlWggPpXjBm9u61RLM2h3CxadT/2
28g8MnzhoGyX8PJxf/e8fxbOGEJW3gYhYDxEEwdTnzSvF0HTDgXGXOAXCiSgHcRCiMThKEtfPcKQ
JHKLDwz+4De3Nf8oP3FimelDBW5oMSCXgXF/wAhJKA+ufW8XhNthC+yK5nQ01DAHyNLQwu+Ur+sl
bfRIaf+FnlHEgxdifGRo7X5B/MDfj04ga9dcmJvPvvMiRpbTHO52vmB/y2eNhxtFGmlOFu3FTvQt
fCDNcZcimxQRWS6pRIMYu8l5ptPUl16Oeec0QPPsbqMtqeqCqHtSjII7pYPYiae2BGmY9NBCQOx8
0+gRz8fi2ozb/zY1tdaw8w45Uk9NnOUxfUMJ9U8Gue8v51d99JUzw4zSpLoPgDoVO5OFcZXTUWJk
8NLnaK0oTf3m2TbiD6Pj+Lb14rHQp9EJC9D0aOFSE92+c+yFqHrMijyjGC+HVO2lVWZxj50xFisx
ZD4LzsHGslbdtYy/4bkGhrcXQvJ1D/bmbXadMcLZJiM8RTunmt0Gpgik4sSaIEPZ3nhVKFaE9DgG
WR7FMiITt61AL71u5uGxPes4Sfph282iEZEUjmWVdV0spttfj8qb50hKD8lGk56p+suwCZW74Ass
GSwhHDx5FxxWiFH7RW5+bjMo4EUZjOHo/eQVfXjqgSRWJ3BP5dtHhz7zq2ii4QKg+aG5GrSbQZ1k
htR4ia9sp6cso5lAJrxbxonGphII+CryoGZMr6twqrt+Llp+PdW1qtY2szu4d5fZZpkb4EwDiHPK
uTnj4ZOx0ZgC3M4hu1L5hJ4uoAAFo9XEJRCA/zvOMcpRtohFoCg0EvXgWeI+6K62m1QkY3IVk6on
iJXoui6ccGgXcUyJSCNXmX1Q9YYbJp38+8h17XSiHS80AkBrB7M871ASCIDMIH0/uQmVgWu2itI3
y6TvJQQxaHOiJmnywYG2PwWM9/a8Ep3Hr4xiFb/6qP/FtquLWj5IK20sy5HJ9MokKJvY2Ef1MIyf
3oq04IPW5eE23N8xscEZC4r40NSZldE4J6udohCIOLnlPRWX98heRE51R3Y7xKq+nJMlIdxmhCeb
QKB/feEWkAYCkhA+qRr6gRpM+E8CmlM865NmKWzmMicf6OJ0pDB7iO3U4ky601x6pHccGhITLf+P
oBOZDkYhO10NrJt67TAB8NTTIAInVUfiEeBd/UNxUoof+HUioM72nLYPT7r3QOfbNEZCLw6WeORv
PxXdpVxJ5etOFZ4LE3MjZMdWatY0IecDt9pWdrBj7eFBSGWB0PmsRYyLDYR8h+Co90OivASkKOuu
hyDOV/3hKT2C7wNlKsX2V96YoGGSinhwJflgxzye5sVVXjVUegUTQEQdmKK7zG3iItywvC1eap8d
BMwI3OdbCW8CO2M7vDVrgcPJZACh+bHcynyu4fotA4JvjcRYHiYkpsF5biyx5aqUbf4++I5H57++
gRaV1EIjo/WYokFjo85r7v4Js8hxGM4lTHKj6kV5vHs6Em3LDVgL3TNfs2S12DBD0f6ELtGh+T//
9++vmFGR1hLgtVPc77j/ZXFdJ2GQ3qoBR2qORpMfy6Rp2NfgchG3eJSZmUDfzK9O4wYdNpD4gfVE
c9nJ0YzGmhyUjkKIQBieQLu3VhF4/ocVQcChe4VHE/yrZ7Mdhr1bREbRfd2I+7NAVrZ/kZ2nGMLb
HJ0xbDtfrwnRCncskDMvOEWMrUjEL9PZGcTKFuqVPcriwd+0AeH9gHRnuvqVY2/LkilpSCEor1+1
x+kYoVWWRnDdmGwlDCmoFp2tMym8ScClFj456bIIPD/I8j5XK55ADLyYwCTpgnjMKjKECKfNKWG1
wnoz0l0a2DJUkDzbvFl/hz6oaN0FEnleJeIK9VVO730MSyw/y11OTVAprlD6vYvPJ1+l7u5HJd1i
CdCd1L8g84CKzrBO7rZ0AW5RolIXR/L3raJvHnVGjfzeF0AHP+Dn3lkDZvEzsk7Djv3gPvptjcTf
VLZSTKcvkBNb24Bnj7nRgOW1+yUdj2uhQ69IHKuO4tTHB6C1q0Deeb1Syq0cv3LJrkmPyhadR0im
Wim6Qidl5GY/yMmvQQrgq3e45kPloepvCLSrBJ+toSYhUo4bKX468mnKMyEJM/wHNW8+eII1yf2I
cw86Y1Cik8YsmfH9WALIlRtZjCGU5krQl6L3I/9QBP+PJZpw/OLXOEcY4C+3AbrlyUpIW99j0I6n
6PngPFuWbLZYzXs16aLXRadejsHWkINCgKjjWmKH/3vZg884kAUAL3jhc0q1bmjdASWT19FZFY+G
JLVekpFJj1HIAMcNVOLUN6OITHy9u7KXhPFkw2yoYmJBOS1ghyhw4CS6KvajIoMSKoTgyYQCL+Vx
HS/HZBMr8ajJKLRkZK9LtB1KlfTEjCy3O5wlTeOGAEHzOY3WDrwAdF+udjWF9EwhocY+zpsS/ut5
DJ0FoELgz/Qsxb7X0z0rQfB1HPEwCJle2nm8I+aIpUSHO3MTqswm8Debb5dAo7eJyOT5WmZFfNzF
wk6+dXEMRK869wuZkcegzhAdA8857dAbrplOmo1YuQFlrRslxolbUj4uTWLhFcNfsWxXnOfJBSOs
EDI1mLtyk9kcYLBSeXvt5EuV9i6xM/LbGMbCF+YJlPBHcWel8OcAdb5T5njWLnqglfb8tkUvn0vp
Ucao77DhenUOfDbTDY9yc5Hjw2/vmPABMgoSc2fIB7ZgN0CXSfVyFFUArZlhsBsj2G9mpvT4wKMY
d75YDAA8mjU1JWq0TXM1GqVwpo3bVl6Ki0DEESA3Ppk8xN3S7OS1R/R6G2eXVvCES91Yv6IBR9MT
uFvHEXcMyW6sb6PKu/oyMBxJDOeoJYp6gDYpLU1sDi7mHW8wrpr0Bi5AAQEZw8lk7j1n2mLViPLW
JPzHP0uwKo4V8AaamHQoCtQL01E0Wd/IvY+El2gk3+eFln7c7+fsWO5/AzINpdg2Fc1HaSw4UMU8
9Mp5bFZsftqtEO2q+2ZU4uOBwU+uFyP9Kwd9ryp9200XMyADaM7k42alFLgcZEw6obuz19x2BjWO
64lUhJpyPDNL8E4WgB/3/XtfPUqNi/Sp1IeMkhtRcRuNSwqwV0PlbJhOiiRmYtwDWVJYdt7k/6cf
dtMDJfMI+NNLX8Z+p4nUUIjBQiLOEPGA9w663pZwJ1dN/76N6PZkhq7MpNBWBCdvjXoCD6hJZh8c
4+pWvPI6e2h4le039I+1WEZVIKiXNaYG+UllPEGa7tQNY1bDC7dtwhQ2j4LUPoD3pA1PK5PKjmUq
6WdjHu8PeoGaXD66e+E2hVeqV+TV4xUchbQh94E0JilPxa6JtfmG7dRAnOqOF5uZQ4hhvt1ndH1V
Pjx+WZdaXkh9WueOOUerhvCx/C473logljzdJVyC6jc5YNDSy2afH+M+/VheeeeNUd+aAmWX/pWo
///4rmIiVCoViRgwFnAl6WM7hrbKRMnqxkVDxZN6Nx2hyJy3anKhy8LgZUXY7TEL1El/9cpx2Rsc
vIaOjRajN/5lWJnC7mMG9UcgS8IBEhCDw6RftCrzcFejLbqxg97XoedNNtjv1Maf1x48bMeeysTu
0LxWw2DEVAbquZ7wIqsyFh5/X9afcMbeHwg/DDhSvHzxkVpeSATIFHNPdXe80X/f10ZAuB54ceyj
yu07/GzHJO7WIhigVjl9ZnM5fHXZIlOmmtke8g6NwLBAD8v0JFou1obqHSlajXvRk2H1MECXf/8K
6TS6w7rdCQJHB2XJKzUv3BRrQtYr3qpOSMu5yHaIrs1CnR01pAF4OiFhPqvm75+sSsPUW2vQWiW1
DAB9VbSpdXuOHoGa2Cdvnt1J/5NtGCJ1H/P+8Q3iuo2NHoPVFazy4KpWapLd/zLn5drE+Icr1PuS
n9D0qwcM95iu3XDWXHy3PuQA3Tza182QclTR8XiO/5LXcPvzjj48ySm+i2dI9MeSIkShQfjjbs/s
ANs3W+3UmzqENsZckuU+S/PFVlKDnQkpvE3gGAUWLLe6AbmoQ34OPCVBbZwUfjvgDG+VOQgOuMow
ggkfrLY6zwZX7NUS5n0FZSlsz/+eTzJlgmoZPcRe/30YW74+cv9CD2zNXJbRZYcMbc9NDj1O++QV
87YzvvHrQBuEkITdpAhR0JbfJ4/Wun/Az2CoAX0Fx/CWVmE8O9fjL1Tn656OeJgK/Jd7p3hRK7ng
BKhKSc74P78+vzVrhS7BW9O4RpaJzackyMCWAM5kpxR0EmnP8L3R+1Cei2cWTaD0u1Rvzdt6CN16
V8ismC0MLFeX2qA0lfVLtKrmyOEYH5cEtdNCqHKU2DZ6VhjFxe07T3mseaXDeLbWOMTLv3Z7SDzV
IhTKWZKSMz1nFjb+YMrCkR5sEVCXyL9C3Gj5VpVLjHwfHDprb/9tZRn7jIzwd8JBcOthlG+3VW2R
rtZ6B5ijE2le2ZDtx5RqZ402LdtsV/8+DSuAD4ZFEZVnpdb0CG916aRKJK7QTr2U//y8cyLzXa2r
nPUsef/nbzK8ZMhJG6dTGH+hkIy4dLNqtH9HaoP7hjMASdIxHM2NSn4sxExWeG4CuRk03Kz+LR4+
NXGQ7j+q4xMPXcYw8TxibtcCKO4SRwHSfIk9qcH57h+ObN9gtxhiptvCSzHcU5Ty0pHMO8ehiB7X
f0BUzvBRw9gYS4MCy7gXYDrcIy3De98a+fyXgJSKIGqqH5Pe05ycQgdkWz0v1fUlCpcmZ5ZL0CY2
znFWdD6/pcMrbNEUKddXWvgZ0PNqxygKzDL3Eb2Rf3FfHEeXf1YoDNGLu+tge1Qzv5qM+m5MJltM
RQ9iHJpTKt8Pdv3nn/wUoe4PT3plyg9AurOKVIPZ2tkudIY/FAnS4VGil6nZAu/zeKgBMugwyTp+
Dtu0RomVVmLaRmSjfTwAVEK0uPFJ8gKgarPN6UtHazbu99yRQhYHO1UF3BMVtPrx6yHTwTnME3aJ
gFReYXnld23Ntw0Gc+U/h3AjrmBFcJ7dEljQWFYx0C4VcqVAbbpvlD2Ha4lbbWCxaS7IkUtgXLqy
9MepJrXhU9VsghDK3pms0p/vyzqQy0vokipLNHTtqQZM8L7hC7KyBnGNRjZEGLNl18KoJfRbDwuD
GhKDcrCi+EJxkmQ2lENyj87JpP35L24ifjSCFjM4FrFgIkOCXqT/bXJPb2FTRnVvdL5si9Zoof0p
ER8gYDXKbaeyaXeji8mz6bNezjmPA4RhadI6NB+wEyBufw/XmpSSHRnsLLMm0Mck3GfeyruannK8
2pGDF61wyRhWyJqeYsuzNdRcykwzCbFGll3eSuMX/doqbXNoYHc95qVjWeF4DVGJ/NQpvzRbgVL1
hkfKEYe3oIb+rkLzJjm19bAtyUdUfGfHzfT8OqqKPJygrejI3kCpu1ea7srKIl7x1DYktWhosb1W
VfOmqPyXD7FqOjk6uDXXefQS4HpBIreTRZQNEvCrYjVdSM55L8vvdCnVZfS4t8iTIa33gi6kapyQ
R9W0k57GAUE1HceKkJap0rkfYphh3JEwbGjmwPPSjqJl4ihk77p9J1dBv58shq807mJOPNZ2Oh9T
njZlBTf9irKXSXqYzqtuxb3iS8OF9wK+9ceXv3p6SiyVOFjfm03u2fLCyFQtDWmUinlq7VrRiZzB
sETQo2PP3L6X1P5Za4LiyD1rI3FlstOnC3PAvsb1vE2g1WRsYwdd082VZyv8bxiHhEdLf90xyY9k
YlzVFqamFJCHnymhA06hlN4bdIGP8PVyCMMCsidbdG4aE3tZJAsjcUfnW5V3N1XCn04gGKfyGKjz
+PJpaEtcbftyCBpQqEAgD2SDmt23kFVAeOiTY01TijOrGT4MMY1e5d6n74449b8V1hgnqpzWJ8fp
CwhDRKUEf7M1Hp2/hwWMTFN8xSqOnzR9pHWfkuqtlGqtw24iU73uHziYAvgcNRLacFu6p/Vkrxod
NUmbQIpahcncUN4ueS+nSVzgDkc8zTU5z1mEXgr2G9Cxj3Fz2drIqAP+c8DBUZOJRDkQELwYayMq
XeRLHuMwqTU1aOL95YWPVBai27SjRHn4lPiwiFPmpr/c23HhSjbw8kaLuTFY4HB5iYR7gtU1QVLi
Xzemc67fIM5FuuoBKHFmT6plJCIW6C2hg5WJ5tPdW2yXh3Jaw0ke6vLdZ7XttrteCEDoJiI+VeO4
2W0D4kE0uXMz7gvTsOnYGvFkQeqNfbbrAXLgPxjHk8mLjaT7HXTDWLqNQN7xxLkivqtOpAa2MqnN
MEHqnSPFFdPTJTkL1M2UFQM912x0yWEcrweZ0JBvQjk2Yl3fmIVheiji0ydvxDuDZ8N7GAu71STa
Mm3WhAxR+4ZrVdy96mQ+j6iMakxKf36ZOi9lrRRCGx5Jnze1nhCgEGueSg2KjMn9i/3YCXCmQJqw
7+/+jDMNv0hm2/pQ6q8X4t03bcrGBSZMbTnun0Xb+P7cauaZwp3JiWD78FPqCRn36afMZmHc0tNP
2e1w7m0yLT7tuS38VZ3lEVWom7C0/RY0RcPx+/4pyMODa/fop7bjq52NBot6L/DNA3vnWK+gJiKN
T5Q0LO4QkM/lN4TalpdaZ8L9fIT1qwjRG1ze1eHYQ/ovcoGNI2+kOXoXWuetQOvYCNKxRDYQq08g
Ef5OwZa+W7poHOem9AexpbklBmbOtSc+bcLKMPh+EUrSRGwAEPl48+r/QC8fJoCY8NqBdAR9D14V
1uNtwrj47KWGlwqWfmRBTCCK6HdyMvrLz6yhmyRvzMjYkP4PzN/8nvYY+qzTe3nKJ7IBlZzqjZ4Q
a2unE7I0zTrig7rA4t6BQsOAEUwT/ma7TzmSOfDEGK/1ggmUaz1Xco6y5lYOFAXXBCWkxYMWIbNK
2qkqLxOwirZ53ZdJUkg2/8fz93weIv07BBrnOc+LXJYkZPlpz6qzYq3+K2tfq0Qft3fIc2+2Mlaq
6mAINYKIR94ZD9McbhsgC1HpybCS731q8baduDPVgMZx+mgWN0MVHuIboTh9A29lsXdyqZWUHpNr
8be/GaDyKZU/EtaiKyZ7iCU54+7YJKjxYxadYAg/e2v3ZfHZzqB/f68CZeB/OgaeEFfpQf6YHt/c
QK/k3+v8HjH5DuGs59VOgdv4HZr1SxYYpN9Y1SgIcFqEVWwHz4TOqiChz7vO8BFBKyi0Celtov/o
fJl3GEPcHaPB+Y2vCsB2azCQWIrMXkd9uA0rypnBqpnHqSd+7BQXm5e8O2tujOJpHo8sGhstujsc
6NlHYWBvW0Hej+27xDMLni7EPotz+X0BPN7Ewc42fLYOH69kLtyTLVqSGKQdBZ0CJBIGZyQY+vLx
YaCUXC1p4YagqmEJQF4rNbiSpwC+RwYcHq8LhUw29ysIEaBL/YuOJGY10sw7jQryBNBfY5r9nOF2
674ZqVR6ufumhvwLhEdfpgbRtK4YNeUSS+a6Wr2HO10t4rIKcjsg/g7wkkIIJuVhlONsDNX0LAPs
LDKmYIWov7jD/TMQwnJel64TVLfW5V7qYYkgEyFw71eYgQyDSwX7QdwlJLIZx9duxd/ofWpludLS
E4eea8Mue61Q48Pmw00bEYH79YBMgTs17ioYzVyCqJKAtMYoBeeWezgRrVFF6TOPr0WkVlhaDzKX
Yjo8DR6cHO/ZL9avA2MoBgjN3K1hfA6mrIAsv9x8q7a/tLPNpMxBtVcjJpyM9gDPZJv1RCIX6Vzr
O+WhQv5dclpaPzt/jZpa5XiRzx0+qnN5PzSaaP1itviWn58oQdNQhDMHY4io2H4VE9VgSYw6zhbd
8vk0M+iZ+hTPQMK1GKHLmvhBGEu/GXqRjkKQx7wIoGeZNNue/9VZ68v9w9AMurdtRPibAnDQhuZU
q1EpEkQsKFCCc3AnFiAVgGq5dfN4QZRhq/5poIFXGB+8b//oDtO8G4ooBQjoCHjiXZEpBgFFLlhg
uGk5C+MXuk5/lvlqmRkk8V6ydaTWA2kBwq8Zh7IGxLq5oFBkKjzEz/5RzYcL3RTRk2BELjizX8Eg
n7Be+tTvJuGx0ES5kbxTnKLjYwICwUa7IV4qNF5XEWP00UVblBDuOyKoSFkfEL4p+Eg0jivDbYSZ
sV2KwsunaUaqCtiYtVNPGI7GV3gia2ln9ZEGDzzLZUKc0bXhQAoZIsWPI+PpXTXidBnGBu51JjzR
VMOYEQqeHfVD9gCnXfrDT/5/IohWmm1uFRqGUyxxWd1XC709hT7ML+9mmwofodVul4v/z/X4XKcr
ahM/MpKFhJWgqtSye5uPHqk2WTbjmNxCWPKq/G5h+8wYxsVn+R88CIyPyTz5oH0FEJUh4yxwlNTx
9vKb3KksBjtJJdDs7HFhvNKFPoTByYxLnaNE4bRL3/XgJLBeK99XosKxAPq9cJ3kZS6FRXANX7kR
nwPHls4zXw63Qy5asRguW6vhqB9vtMZyGouS4maIdT7PKJzjOm1yQB255IYcGIzvaDrjFIWf5LB6
u5Ql3dR0YV3GCRKk0BBe87Qlr8LJKj1biHH4sDJNLlzk+79jNzrQsBnOTxWSmvTPkre7+gr+AS/E
CCA2bybOrUkhl456KR4btFfcg3zyEhgSDNx+guTHYr8S6WiC7spcSWnXWz3ckDi13Mz++jQ3ESJn
kLNlGucKwsj5mHb9KJLLYKUdREcS0GqPZT3qsToJB24No11tRZYbKTyL5suwLulQbuefTsSVbxQi
C+s1vfVeYxwZvnOyKzWxUzYFqpZrcUISSEx8eieQIUjkr76/QfXKLUKBMBjLt/Oo8AS61MrzWVkR
Y2H+FHx9Z/zkxKxUpjjSLjNXPeT9ORT5gYnfhB/hWl42VgUN7IqLiEzCGYYMjwl/kePkUVIdOTtB
rHCQzN0X5eaFxZPZN+B0MefR0n2KLBbE4pMB2MRspQ1KRKSYfpq8gkjpcQac7L2aa2j7AOi4Qnvx
2frn9PhnJsMw9D9OOne8LzBBX6VOU6Fg/AfrVd5HYfNNs/sgPZ+9SwnAPkXS4Zo/vVgluLalFZ7y
xabYHTWWSG/3QC2BY0eMvodRaciqZpflTf68DHsrKwlRHDsdLOJaeSTDC4yKASFFL1964QqFRtTC
EZY+oJ7N1H2wxwvKd1V75lfY2b9XH2HnrohwqeJkEngz93a7oq+s2Pb3pl0a9pByLb6+J8HG2ri7
k0Vg9oKyYv3EROhyC5jTyQsK5moF3d1Up0+H/45KeSXhQkAYuPqbCXF+9nznaSC8e0RMlpTZXT1k
4dQc2rdyGO0cxtLUuJ0hXhk5up2Dsrz0ZdvodgqR8ujHm7r/TwZOezHJMNkmAC+soDZrK8L4nqBw
NUdOJUxMt7WRvAc5vf7FH9o6zVBC+wUn0W5bl0LyFRJtTNsPdruNquVkXXdldi+NW+lpwb95mu02
1UMXD+3ntjnjJOh8+SBSifWJGyDDT3DjucbI/3Dz/9cYFAn4Pk+q9ShXvK+AtQOrJRxKsu04aNU8
kD0t4xSdhBEnm1lKA25oCdQ3y23RcpEhs4mtQU3rRoIB6srweuJ2lOjx/Y8a48hFS1WU3rekVYhP
joskzDsB6RHWWvVYIRFTdGxlszYFvTosWbeSON4TCvQu/YY8611iqaRTI16dhhVqJEgbPVZU5485
UfpggUpxgFClcrmQ6KFMAAXTq3Qk0t541YE6WEQug0JotdFrwQIiRc1Zyg53n2MEcL5O2yv0u8eG
DvSyeDoXnFzxjfzM6+vrPbBUVTIU1drUjlrxXU/u9lS+YzYGYeY8dEcpbPrSbmUMAfiQRhb0qQ14
IDqF5ytmWLV0IUVX9o3oGKpFk0aEWMpUA7vmhEcVd2PUjfEMjmr8VbcQprBtw1qKu1Vdck6jbksF
0akFR6lxsv8qGqhtxgT9IVN+2ysTrZSKBdzrLTmng7tW27MuyrvSIKJYhqS1IFiVtlii98L+7eER
wtCvD4OjgGLl1WEJWYytEhweH4GwqRxT3KMRSVG8nKy/gFyAAWAF/WwqBz6ULFyiFqZrABrgCL2P
DqghKa1bkKV6UvDCM1y+j3azohfyCtAFKPL8jSoOqbnqxX8DXTIvxgMhhyOJg5+GJFxg+9CQcdOc
eI2E3n3sjVS9MTlJ5tFoMqXULuZw+1rr2x2Pk9ZOJj5E7v1pp+upHztHTbjGvY1APSHhq8LhiI6+
qNuBPwEdwoGvDy+YQCJjWdsBYZfZwMUn46ycibTvWUzFNhsVlnCQVGV9yPNWQ/oYiRnmjC9w4xgM
4zNqXZ9O/2I8Ww+uxkCOzd9xldQY6tYrxq9cKvnARE4+ZM57FNWZzkJ+/c0WZ9A7D7kCTy0WFjGn
5myPnnYzMawL0PI29R5uqJ6lXSBIgiJ2+drH89WA5eABcQJn7310toU6jfDlHRTfu8/Pf1ee8cTG
08Kc/wokEm6NkDTI3l67jqXG0av3tfRJgeNOmv+xOD4okKr+uJ3jZMLOjPQWehoxfCIdiky7PaJ9
2LZPudr0V8mRZhZJXWzSWQf+pyC4K0I5lUAijGnPzVVTtZmc5lugtGECD8hUy0LmP0uRV7eueq/i
otPS5eHn68Z5VRcO1QZ/nflqOswYmnUnUpceHGJTRvLccfDxG/q4cCmujUxSgTcQandeedkpbvar
W6xd9/1Aks1dlg2+ePyD8ufKgpKHel5hqEEM/oLuzJGw/ANtBpSOakYd6OKiib85zkhOuuIRpUEL
ELpSGqOEENSk/6t0YpmwScCTLpwvWSjxtp0FUFNXSmI2neR7Q24Np89PnGsTMZMXwlSHpqGyKjBW
7X9qSO9zMvpwoH6htILx2frOEFUUOX+h3VrjA7XmY6fXuNGrGxfPHC3XbdjburLsCIDb3DgIWj6V
CywBfqudWrfwCc8FgDzYWXKgrnZ5npy43j/OBDLd4DOYPkp9XDDkNQmuAbEdcIr+kE0iL/Z2UGXL
BpflYDTHO1mmSZ5n1uI50nwrF47D7ebSlN4lcS569xjCQZjZFG6GiUYpbjTebgdeq5lHcEjut100
fHK3X8wv8WzLXfhvBKSpzVbeHZ7MiHMoebcwFfk0wu/aMu+qTaRXIBzeQquhUCCyphEDssMaoxLg
9i8Z7YQ06e+ZVOPilvrgrWX5TGNrOIndbtX8xZc9uNIozemHchLSaIdCkCWn69rrCIY1WMMdUjXN
ywGLSPNRMOF8FeAszKUjh3g/dxl87wXF0LdDUCYctcFexkyjAPKhyLzcTaich0kGDyk0QzleMyA4
1BFHExPdlO12C+TR0QBJeYy/lSI61zcpnpUrLtVs0rdO2y3rydm1i3u9UoPpKjlh7zxWifcVrZVM
vSA49aHvUOwDeI55p5pdFdgU5zt8ZPDg4O/AUlzvMjfx5v3PljA3zH0Yd+h7M4JXrDDIjafJZwHu
iN2zitTOQq3uYZrn3QD1lo3s6ARme20DHPooJMLqktoLdBr32xasXvz3eKwjXRE0qq315ixxkUzY
RlHdThbDSNcUOxyIR9SJFGPwf7zjNGPYisHNI9guMeVZBIPlxYsBVNyHu+BcmwEvSMHD0kNknN1e
V0u9mnAX7BEGkmDLb6K48TnxLYmHAj4M/lvQETnx2bMST6JgAWYzq8vNEh2xAeKojwWv9nsVBoiQ
a9NbDwqTCHSAZQHMOASW3un0Bxf72y/Al4+shCMB72XpFv+8RXRvoGAoX8Ho73if2Q9IM1dgR+Eq
ycjz1Ae1dcWjAfCThVU9BLLNyr3KQH+HIaTgrJoEkhwd948ljNm/Zd/tvDdaP7wXw2VTVz+WNMeY
XMurVtR1eexxOjhKbXfYtxHOJ1gE6ItDDgwwGPhYGytIKb36o3hcAy7r5GXvZGMAaaoMr6CfIwmG
Kw3TOw7EA3RwgImxQ4ez6nbh5DZjRrngKfn46xG0J4kcR87gMHvbHruu+aAv/SMJBFL/HTB3qUUi
GnqDrVh2gI8Hy+lxewBZiljlRJ6X8fEVtQts7EX8WLZ7rIOimUWgJRDgZTL15MWBVbefXnQJwpxc
PEdNIFqtGYTFKtHIy27OUcDOwl+rEN1z9XjP5y08/zaj6HpJkQwFDeKx8C9k0wbPkn5DrTSgx8ow
EMu91jDk8zLL4+fPLqGB3m4DcEtsqdyuh2pqtYlN/LNQqi/n42Ki07zPirBQ2kL3GfwA6sLo/MPL
E4SKIGVFB7bBENIo3XIQlx5YFxB6YDIe2PoqEjcIl0wN+QP3NZCZqKyiZMml3IyZ2wYGzkhqPA0H
seGGQ/39XhWfm8I7IU8EkUe7vcXoOFxr5K0PKCosEu3vBMiO6ZdPibTnKtM4mZ0VXMosUGaY/F7Y
h4imQPoY3gPnDAOy/WjA7SA35f1TGcuy5HpW/lYA+iL7nRET3DFLGkXL5NhoIvz1IEgbei4r464e
TbaqSgocZvJm4WvezvXkAHwAY6MTe6LKVMPK8oQ9Dw==
`protect end_protected
