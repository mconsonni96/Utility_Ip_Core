`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
GvCnbjwVuvdkV2sE0AIbuOR0KZMLn88RQ9f/KvOWBTnzX/Rb0gov+rRg1ZCsT/NlsldccjqzE2x2
52pjD2HKB3NXk9iDNeb/KG1QJU+N4WYX3YGMmmdibNjtuXgGhf07g0BZ/VWcZ+uvaN6k93RCsuMx
09M9Yi161HS4BAtwp5Ce73cA78gCNqAnXOvrIhMdLxunUpuxMIIXTwNE6QgigowqIS63tfMKYMnL
L+po4xDjkyZ1F2CU/cOVA/vTdo3BWBuCeaLd6NIWKX/M2xE1CFaZdaYAFSLcLf1DyEf4ZIWFr4eF
+lCA2ndUvZlWDk7gbSapEozkkHhV1sHX+mWy7Q==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="kGf3oTuPl/cFtWrnhONlsbubmR+BNxvGUDVNOuDND7o="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12496)
`protect data_block
9MJSTHTK4RnEXpnl3nP7DBH4hZ17f1XYB4Sf9x5bsaoxBAlmaZP+gUp3LTE7qtB+NgDgNKpbITzQ
UWHykh4/PA3LlwLkqOTQ8ze21OXpdEIjMpxAFm2A76QWsOZCMWvtF7NJAXZhy2vRy+vUqlJPfh3B
UWAD9pfc5eQ74kBFEnpf6LpW6w7edrUwoWb9j8/X448yo8c+glS4GF/ceqrT1Bj619eiUln1MgsP
ATzS8xn2zNjgEAD72yav0tv05tRA5vVFWz+z2wye1uybMHhHG9lgh8iYfCdF4Jzm5SfnvTIqs76c
5DaDE0o6zmAy+MZmXosIb9Czi/oGNUg9SL/czuuRLIeaELqxMMRtFWP01cqVPcMTyuXUI+UKjwQP
Ob44UzhRK+YLbpUYx+yNQRfJ5PZXSBtIanu4zRQmwC5fnyk3FJXhB3GcSnhdFLArKYk5VWR52RaB
z0AmQkMFEf4RavMuPs19Fi1xqYdDQeRemD0lgTor83YLvMbftrJpGvUDdToQDcF0F7lZKTYHl183
8RZ/kCcnFyle3mcP7HQ+UkX2G7oPY/eyYZg31QP9S/jqtzZ8yyJEAwN376sWE+v4mP7QsvPVDulp
+PVyECFl0UHG66+D5cSJeT3vKhQliJumVNZMp1nJEf41fY9auixJG8HekUhPgzKUJ0Z1mgekXD/B
HpzPyT5ux5sot3ZPkmey4+LG34kMoqxrREt0Iicz50OWwS3+zaLDVFfrapz6CeboLXCl1J7TPZlt
7Fv1xi9l+sNAEdt4Y8aQrNK7C4DEd/t0sr+4oE9k4pN4d8v+3CTeM0RHcF27RKKVXKdga8WeezAg
SJR57Wxplti4HEP28DAlOTLqhUOtatS54o7C6Hp27zgPfoQbZQ8vlB7T4I6PvM797ACagIw/hRHS
HOO+VSqWPJycT23BBMn8ZHpNxIiovD54Gqke4Dbfcrtd3pRZ5/DnQW4XUs+X0IYn6yPIMFRx6kAu
I7YUqQvLLVS5+R351wvzEnM2sJc+7FBCubccTcRxziCKdlxYXp8PcYVXP2+Eg1IuGHiqIpzVTSAR
0GOPveDZbecgPzoNGAa5ujBOtXXo0kBQrGqZ3dzWuBzuGQv8tvwJK4VoDxOeBwqk9VRvX2xC/dmt
4554sop1pAcrE0w3TOAp2yatVqmicn29bjrAOvZM3rygKOiusKlpaLqSrvnuWqaLN1wI4IU5/LaI
gxg3tJIOXop1+EMwSPxPIigQw1tJ2cwLlxwg1ByOmhWqFx9qW8Qu0m1/U1l4JmT1mQ/aTYGj24JP
K2fLn9LFy0XjkmDFRzf3eHjQrf9DpFrxLetSghWpbNc2VYVOydC3PAN+suFHY0WSIy4bIOFTzW3N
ujfDtf7mBSJ4FqzHWbTEtjfaU2+vqtEAlbgBq/1FCz/gVRDrd6bVX5KyKZXkI2FXNVJBkIgGMPha
iEpeuA2Mst00G1T1qnfIj1EL1C2AFq1CHwE22Xhml90GR1NfuRFtxNuAY6FLaWO0P7hH9m+UF4iY
T7p099MVjAQ5vNEMcG3t1Kmn/QGH09WG4PfsCiD0m+S3hkzyHlVhnyN9EyjK6TkQjXMzVJIjOPcZ
SV2qZ3MW52kwPAYSvF5teYniH0OkKuVSUz/5/zAijy5uP5pr2we6wQURJRdMiJnIG6NUBHCVVB5w
Y+23UKJ9Z1qS2aHulZseWXqIs/UwzBs22ojJfh13DH8Hq5bfywmdKaSr7FhszJZ9PeEQ92b+jnbJ
yp5cWFuwPUIL5WcLrI7vm5+exGiInDOKNXaX39RN8hllDNBZyWAWuYmP/jKFnB2e3HcjAkNB/VHm
Cmt+2I73R9OoLsdgHTGNQIvBne07swJpWH3KSy7hWpLS7O7pmhOadYNBCVzUSm/XGs4gYFajTbw/
S47K4vsSKwCzOxw+FpJTcKy/p+9xDyWBrTxS1EJ9nJZZdnpnWKqAWhJAop/xRGw1YZneJ4c927U/
RZn665fJggcnSzWf+S3l9StfV98j9VU234m3xd6IvzcyjWFtc/4/YvETqiXGJlD3+x5qLc1sXHo2
PuchEEBvUznYYcIhCk7tKxNQcNxdnkRRHD4ImzYEAOLoUzoPGaivZKnPVJ4L7OhSVXy1ePZ3XBfP
Fqxb8CfBS/0LIYblyuTJNRNL3xPWHowN7Joi/NimShDs/mdul6602yuc9P0wK39vusdE1bM2fhcF
TiFWSP3abEVDlFE7WlqLk3y1yCSMKisxv2syJqRNiH8A9zK1E7u67vEDlbUjJJHahEALbNby0nFD
79K7YIOo4vzHqgRICfHdFyWqQvKW9Woo0Em5bYIOAc2klHsdkVYoP+QO1N79EGA10ADXPFG5DatP
a7MAHSHBjy3nKv3GxpWQFpszagaDxgDcfJLSp1yHq+3Jq7zY1N2W/aPqzycaJ0rQ3hiPmd2xa1LO
aFJK5m8Nu+2DCSSDz1nrYmy3fpvx7mUyjSQAY8STmBc0bWUdbnMHoOKVgmHAKU3YMG8C0spS+Lzd
Y4NaWv7OI/tDLPVA2CaB/UrUU0sVj2GJfUrXaXFV/eBQRJSHeENdKK8T28qPfNBifce5alESj7mk
CXnu3vAjc1NPDSKogX9Am5765kyTSvViHanV8z1BrOgxRopg9tHknbr6T3TqzHExPLLGXtSVJ1Jc
3csN21mCuRYXB3aBP5BLm+PNTT2Pz9J8pXxA5zECNLCd8lVrXEHA9DxpNZktIWtNqSgOeBKf0tHB
MvaDmQbxhcZWFtKHDO7ESwhkPqPwGNXYO7hcErPbeF/Vvxi8G/1CkSo8tLBCIWCmbhGo6Nx41O7e
ULf1vIsnxAoR0vPuuvLZ4B9/MEmF++IsCgGprDXGl96CceMyCnJmrRgPm91Be+o9oJBql9FaxYFp
0f+Inzk/vUCASNb/OTcELEEU1SlhjUX2NtE0eje46oi6z45Au+v4R/jNRwGVn5JucPrM1QIfX53x
rB1heV2OmkAHxtNJN2IT2/w0X52MInoQx3RI8QkGzCXFA35RdbvS6hiOoABA0NkicAPc3D/i1lEn
pyUKmSfe9FuoZoW+59wC4WVfa0NefdwPtqDPsXmpXV6591RDtHQD7RZvyQgD4rbKHoz6iSSil5xY
lxwr34LDS13L9RdsL4/FthRVMmUelqE8UQl6WsocdlS1tEbUf1ZvfljvfXD0Qgwo8TBDMmlSeAK+
/4AAoUAtr6DOKmzMquHbe8R3abYahsA8dhzQeO2Ga9nH/4MeqWBNIg8kERuGd7/itemq34q+PHBQ
JQKALWyVK+Vvxv+/OvacM3zMT/WprirJiElQmo4LlnVeks3mbTEgXQ83nCYhCk5+OX3TCHvIhkqr
d7mDi/tKB13YwxK7pC1WpQGqRP3nlo26PHFD61HjpZ/7SGHf1MVBJTWbOiadHqUthkng437nQoYZ
nPLv6nrnOAvvz3hqAK90eddFhzazD6D9284pkC+Zi25SFlSFVALcCBGRLCWM6hQJ2bhCIKqaOExj
TmqKcgflpC9O+FRbZ47c1Wn018tDEfJpLyBBO6XvUG3Y2Z9ysYu/XAQ+baXSAU/NGWyEkIVUuXz3
FVwU1ocq97AiLTR1tVj7rOGQwc2EIQk6QaSc0xgBQQd9qreax3EdmIzogemgeCQY5BQtUw1CuVjG
bRVralWEVlgfD7QX0nZJB6D1Tq/8B5MuvEDCRBMZZ0c4HLF2qNRiN0kfLk7kS++VMwq3lRQhkBhZ
cp2Lwj5gA3Egm2IkPtTgzYFk3czb6o53lDOjLv7NxTBSZia3+nsT7LSrEdB5Yrt7vA94LqsmgNNr
AiJjbqzblBWg30Xj/eaiJHlswV8f1HtPGhr02uIWIZmE198ghpwCa4A6PdZoN5ux5+/C+oKl03mO
LeqFM52ROmMToMdVjHjtBt46HbwwC67S+qNJx0pBclD5Yo3d6wNmcG3ZvTgIqW9V40cI9Ee/sSBg
T/uozPBuVEXmTnCuFnp/MtXg50tJBt0B+NDboI3AZd331ze8OvgthSgyQoj7wbDQNr8uljJqzmS0
2z+bAyGWU+dP0Ce7syANRW0MgGIr8kbq1aaEyINPi/sDVGDgdAHTBzYrsGniEZFslYzJ4DlmJd30
szH2P0/H+tShP1ZIyCYUfinrpmNwOJ0EUzVLB75DBduzBnQPFmtroJVX90GzD2h/lpNVvEdC3oi9
MCtl/T1CNwy5OG9LbWsbQfxpjTwGe4ure+FJjU9B3/NmUp/6/7vHpy8YuBP/dD8gDgYYVqmTaFXY
sv5Ohn/AtUiWG55QjjN90muk9FWjekHTXKDdkUo4uoJ9OPRCHnqiKy6efH0UR4xC5JYfBq/jVa8G
2rCZiZO+0ynyr2P9qzYEU6tEW8enZfTf+fDDZUr1bAEWJD3XHWa317yHcT9DGcQKD7gN3V+fXmHP
h76SVMqzqJARDR3dHBUbFp+zG1mspDf+wpTaFesQsB1lMkisMnG5EceVx8WQjc6cIJ2o40+oo8HJ
5qmgjaGdEIPgVb31hhSwxxaRVVweplhqSas6FjU4WfcslBOcI9mVhNE5D6t7bUECBZn+yb0BDGbV
4D9EOPA07f4m0TTY6xKabG9IbhoMpZcViwN86pIUJ0FeKSQaKjqm3nSN8yeym2MpY++/dFsDetvt
7C39QJGRdB2IY5n8aYzrfUZPJL2GBmMNaxASTw95G1EW6xAPQN8LikTew2AxuGmJAJ6ShHkEqbv+
6HrOqo6xikgh9MaBPo3kg8yPiWzOOxoiEYsi90r+kieSBL6y0R93iNxDeJUh8nRAWYNOvOWcXFm/
2tGrp+cBx9w1oAtchKCFTO4SDC95CXCw3VQ1Y2tCLlIU2joKuT5WX+Avfjl2vxQBcBIGyT1yUpVU
81r7Q/AN2byGiynW12/gCMec8vAZyBRGZNsO4tLA2WQO4dr/7cyuiBWtX5SSbgaJ+Rl8VLbkRgsQ
mDkUUJr/zlqRAgwHrXLGk0fDSjbgMRcNK129nVHXWi7ZxFp6O4skxA3U0A1YW0mHzdgGs/sOVzAS
mxcHlC4EcWIvWyyQoFFQnQ1WFPT5kcIz+5ADQWLWpZOud+6beuNzkHaeUt+VNKiOnrNvvkK7O13d
QsQjJ6GF6Lm2IaextXjSUhZPmHRTEIwj94RH0tnqx54qOJKl7Bwx5xaW5tDjbZnyXqQooCzfXt6g
haQbpw2mhMr/WMIAnJ4dK3K0QZRy/kgicZRAeJkN4bnUs3UZc7IPxFkePLGLOTFMZZr8aFzSRVVM
rGdIPsIXgcpwLwc5/TAsYRMz8QBEid47ixp8Qmi+N30SemhXe3rSDDFuQLAo9KVZTy7GGuqdlnyu
bX+odfJrnIxelSMDoLY1Y0NBF8s/DasohoZufJcv/wW2wyHWqAG75IGmub2WeFE57LMMVdRkpSg+
jaC/qSzmxue1lotS9fMh8QzCFNuoY+9DmJXZnxQsdrSHyGbK+7tR/vmvTE85ZRyXL9IcgTldjAp+
JhIK3u2eEJxtJocZEEOqg6JnlFxwazqbAKD/DV4M1ZzPvsVQbIPubsmW5dgqzDWT1rNNTMeOF5dC
/Hbu2MtymNAdFiE09IfmIZZ8w637AIYAtvISJ7qDC1Cj254ffaxpQXkRY1CTO1Oqby2IO7Nd3ylp
zJp3cVgbD7mCejDxvp1bEa2WXjpiCoeJbReAi77YzDrWxgM1GTaVqxKUN4s3Ckhs/sQ3aX1W35jM
RaUBO6QrAcylB4JkD3Ea3H30doKja047rT9/SYwE1l0H+OjnRdv7OkKBlOMBDMW2c4BkLaQ8EW1K
qGIsusMUhxQ5bnTMO8K3ixmlQuMq9v+zJPDa6xHjyCdW5fQtBZ8dDj80NnIEclJG6YFTIqOzZZPM
U2sVrgZVO5pvq7IkvwrVLG3kqgVDx2XSKccJ4D4KIWysFISOi07eHzR4AONMJsWEKSm7uesXPFfA
M0V5Ay/XEo6XYvEHAop143/5JVJv2aw+K/YhJJBflyE9xxtbpKwAWEUnx7P/7NnJwZetmnlnPqWK
nc0vTkYbdyd6AgE6Sw9FYWtZikezSIr2Dju+PXkQlasKYFq8msNAK3ZXJFDxOYFL63xZX5Fyzrkw
jvlMoATU9m4Ktnieth5sqZhpxOPxFQr8Nxgr5mAetNO48Wk1ikQPzf7hfRTUWM/Vh5Xr/xghXsRN
IV78Bq1fx9Svuuq1wuh6CVdUwdQ6y+742pWUYZ+VQomzt+k31bUjgO2eI40+3wpuY9MuKPditu/j
LcLoPPeJopwMXj53UpkLIpMojRxgmXvmPKyIwRAKNDF1TIBdgvCcQJb1vnHA7L4lymk290BycAdB
qXoTS7Qjii5O/O1R+NI2ae5cHGfIOniRwgHv1EvEvcikFS9Xt65evK3A+mFbiylDUb9/X3BZaehS
XbSo4FI1EyOYsZggEHTVZLwNX5CkyGBzG3gq/CkQlRSFQvSKkqMjOhxOt8OVSF8LGvC5hIK18k62
XDBXA5fWJKhjiznmFg7wLK9kb0dFujzjn4Hx3pzepPCqzwMtre/2mU6Y5oBdI177Jgb7p/fH8+a7
I1BsfVF7ssQI4IUzbaA4du7lr+W7Yx7CRX0lEez3yuWyvECUcH86CgFi8dKKOaflU0zVNVkxktn3
McspeyAKfk+gtEY3ay9S+0exPLxiaDxp3DmxU3gjK5CCOt9bnukRYaiFyHc6QGIqFlcbr/bwGk21
c+2mbtiRn8Ble1Cf82/zUclDlLPor5TMoIuKG0kG2WqrYXSFkjA9jyNQjTzZ+a6RlMRa+u6D0H0R
XQnrhIOm7o+TiRagTeDWiojdyDbWCaeRsc7WQEgEdIW1tzGBMOZmxhLhUnZfe17xoQKVg755m2OY
VLepqk8QQQeT8Flse57tCO01Qg/PhEo6O3X8bmVQ47c/1OvmJJg9PZfpyHFZ3AMRTuRu8FhpH9+S
ufclGkcH3F/PWQXa0fyfgsuIIWhaw3/s+FwheixSEVTZFm0K53ckr1ToeDDQuzfbZbiMXjd45f8F
qSxCbQDa+WzbzOGdEyLlII5VkeO3QjyQC8+5GuW4eg8x5YoBUj2Bbgg6KDnXS/yvP2WAamu85kDu
NfeAHNqvUvNiuETYcuXmlHnG+MpYKsr3fTx+P8sSOoELkNWawmSmlEjLd861nc8uW8tvVc2J6mFp
d9QNj+/p1mS44dQyPSFRkq0JrQXX9TFBdwX6EP0Rq5nvnUZFJiQLbFR2v5dZ6y37ItZ8adHIsqBB
a7tu0KjAfP/YqDr0mSOBAB8np3c5QrJ2ojskq6Kg4oVYfcWhROLzMHQ19klf24EJY0vdaAW5NaN2
CJtvst+YLoLamfl9PBMzYqDpROXUONnTWjDdITSY2zehmVVdYjS1YuO+7FyL7DwUlyxdFBtqWANK
mWcdn0++YFJhvamYCzhl3nViJVdOXVN4JqMUq1WY7bEXLgdJTO2nhmdBMHegOGibzKTYypYChS1x
id09GUOST4OTiOwMipzlcJVZGCxWxZWion2WExDHWB9RS/OK0c0DhiIPV1boONvRRf4NIx2Cjog5
5nt0WXkOzB57dEViWD5cjjKm/MqHk7jGfgwRVJ3siqYuvrNnsbn7aUuT799DsD0si6tzPLDetsac
rXi6JCoMX9rfUBMJaxiaTRADKG7KWGVwIO/W7TqBw4XlM0MOzyKej1lnWshpPCedsH+BSbKaCqNS
SZ4qOGn4kpmql9HvcN6W6OatxQWR+cDpQQy9EDpHHrmDLRLQtG53g68AZ0y4+taqTpWzGs+ghs04
FUcMp4Lh+fFqLS5qJ1lyoYEUWYehtzHHEePlODJlJ6xfFn6q/q5tF7zi5tjd/gcwc9M6yY1hC+Ko
ZBnzloKDfv48Ne5BUwQ7YgIIuTVYixCiEiRt9q8S4JFqdyQxHkI5Vs5LY3Q6bkvLbGjDk73tj/MC
FjEknCYr/XejE5NyrfXiQ/58j48HGdqvnWQ3QX/y3B8fvAQE3lXZZEdAj+iSHRF4pwlPNxoo16CH
G+aQUfq6juo45c9iNm9weolTcmzxMsflS4SOg5aTzZqbZSxqONRAx4XnXFTv+snVftGO9Nxk57OH
N2MIlfOTXdJnBlY5pXZwW92jYVagFBxnoHRdRZLfs51UkQZZVVzH4l+gO69uo0GJTHYRTlbvKsVQ
mI6FO6UcFCmtbzLwwWFerYP7ctO+Uc/EHa3bNhaffzv0ObK/EGSGwIPFxeEjnMoRItT0GON6zgFD
IM6Ek9p5ue7HyuR6kviPCCKaHAr0MiX2/ufOBPCqGFZDl/KsqCvxpY9wfn0p7EoBPetHmNwcDonh
lEH/CBq4urhGXCCFq8DylCU7lN8n0OQSSm1Pp6wJPFFxAN9EHLz72CmxlUfx6PgaENHZ0/dDhGgK
O0NY0ejPqETymx+xf3IdpNRsRVTXCvtiZNV5gRJfxJhgRf0GgqDlrKARGtRfo+Ey0oO6+SuWF1Ch
BWErxYeyYz3YTByIvOCNSVmOiobfi9l7pM/ur6+tmVeeq2oB7cr9vcIOcTvw9yYSiCGlvGrFNhS+
gOrGTcodZ1bZz6RKuXvbLJGct7EfmND0FGqNwNlzRfQNKt/s0uzlndVSsI19syHOBvwlH5LmptZV
Yg92V6P+tAMr7SkDdWfK7QWaK8/n5mmB9Io13CnXHZgxVrNlh5czWgj+bmYUEYB7wX7AiYcHBpBY
TvhmUa13gYBU0GbACKsX9LuCkoLHW4tbkx/FU3udeXxZePSiL9FCfBdWPhenoUVXYzl4kLMicpi2
oKB04zeez5yPUWf/H14FAGQQb80p49IgJwUBFvidqVFJTf4uSKL4/9zKhwKiq+ubAjavMthEw7T0
6EdZ54qx1ZxQ/+cSNNITZ+5TAx6Kziz0QJokOXfkSq8iF9wWhxs/FMpghW/hWkPbGMR94tjuVEEr
8mNBTys2RLfdHhCp4JVll/5TvDRRpQAgGyzL9Z+puvorjHS6ZelTVunirh/TEpk363wvP2yshYYv
chODHAkJ2/kEfO3NXdnk/dO3HYbn1Uug/W24W+z5xu4ZOkxsBIVpKuj51WKph2YmE7suP6YaifPc
xKXfGWaI62uV3erb+k/i72rnKzDnUYG8LsoU2XiRZE9xNVnKH6m/uW9wHo2Xyczj3vWDsQ9GHMYC
LT1+6fgOPBP4ki9REhop0470R/UXCTuRviGxPJzis6OVtI7Y4M9gvy5lM3bOfSnbBV7x3ZZ/bwq5
FbR4/5hsUXJEEBqRd16a/Ve3TZgRQi0zodzG0Y6ZIdOTSvu0fYNHshYqZqFNsN8qVeav7P0fB7UO
/28INcdnlYQG1dnxa3Om4Itn+xBiwIuXjyu+m9gdd2GCQXKIzSPuupJsLZA1AxqqYK7Au3adtI3E
AyCoMH0uDiEEQN6pMr3gOSkTZkD+ib5UQ4wdnQQGfINsi/5Tk0uVZ3dG5GVipNgjNk7a1nMzbrFm
JWAqAEDjfbL0L3CsEeoW361/eGG9w0YYopRK5rsYe+u3pyZOgE2gUH1y/TOBeUyFM5HXRt45+aI3
eMcsy6IssiCUFrzt3agIghR9Rhktln6guJ8rAdp+BAzbHxOb1HxsaAxM/5b3kacSs2kNZpj3oA2f
dE/5HmzL1IhrR72QQu2CWS3vPSbHyClEivpYmzmF52aJUBLH1Iyi0hCHEM7FlGjZK2CZJY8LDZt4
I2wd6GNVZZtaLmXvb0wgnpvVYhOCC/q3luNtVW7lz8jGv7owOfpn1D84QRBaJFFoQINj2wyIo4Bg
PGsZ7hlvoVgr6Qh7P/XnGEqFTNj3NgE7/aJjYT0VWp8+aVCs/lOTPtdtLORuBKhJGkPHg0BRnURu
W8oRusl7E3Qa102aIoEYr4F1bywGOHSmfkvBn9uxEXDNcoPLeoc/izmPT7MugXRjYMIayJCAnS8v
rNnxvbr53KFRUe3iylQlSI/d2a9V9rsEWqJbrjA45t2LeCL0RbFrrlX2koZE7IPmBP00PVD0WVdw
fcNF3k9mHYMkz7VjSvQg+oTRQZMvxdusSrQrbXVIxhVeueN0h9tBcwvQ/pI/6F9KQceurX8mwyiq
hHdcElvj1kzavZUFm8BcbCDK/ZzlWptXEFGB2P6WCwSpCFU2fcfE2DfEMmj3Qjt4JaWpjCR5+pX7
JyS/W7JIKqQV8ddVEY+ktfm8hR9qI2LqsM8qIbfvloV9gKMHRHh8lDuIfO4UNz/szz/A631N7WxJ
WETWEurOOWSPOkhjHwVtX2lXlNbvcxaJHT2jOxiIRqb6fvlr+0BuwwFOb3RyWtj+nZa3FKwnPhda
mEhgtpUpEPqmU1A53B+PUtAi6Pb5n3aPdAw7ItSXspoY68w7syd2Lp9rnB58RgD70TA3deFd4uqR
592Zf8KDUIjpmME5Qvzx3TeTSMdL8TV0ZDwkt+6iOG8c9fDilnOJgjtZjjf/+UZCQo4lSovC4oRS
Da/mKF6VmKE8JoXumCwPW8qfiwUMzscuTibJijjmvd0FUrtQQXQTXUphl1ol2fJzVYSCrt3TeW2A
7uimeFUvC7Ef3dd77G33C8RaH3BovB09MYLBTTQnOLosJ5loRxmzx7WqOP4gtFhCAidb8zbrnZRn
t8Y0wQRc/3Y0JvC+o1ahrjIV5U0xHhJ7pE0JSn5J7X6On/5lxXFjAMzQAVr9luRCOjGc4EJFIiW3
y0F8quKhuXoeZl2SR3s+eZYewNxU9mKkDhLbo4x1QBSpOfRtjZZHzf8hLmXrEKAUmGH17ibJgqxG
toARfKUPS76zCKHThdz81s3qBdYjgBBD0OXp8kRLtpn+c3wYYrkzG6QYO0znh7JxoRXRhoBG1giE
JPbAv4jTfmYZsorLuU5bADV4OiKk6Fj/+nIThlWi+zh85K0MFU7yUAGSXI8AiOLkYZ6vnzsSvqQ/
1lovqjDpZjt8nDIqBjiB7klrQh/uAxbUEetAcm/7uw+2mer9Pd01ukW3BhX0uAsYg/kyiEsPp0iE
9N6bCEXueqZUjwsqCLLZT+N6yTPB4vfVnzvbbQNn9vXtP61CdoGI536jOvfVlEcJ4reYwC8cd0g9
nxyvM4kVurROsZf6XVMKLZDMoj6nJK96L286Vet92tz4twOKNTtfUypv66QmodJQxnudeDK236wX
B/8J2luUakPsJRTkVBq93+yxhG1fd45mRtHHFViIAAhvGEdW4Ldye3SuBzwzQ3lSaN0k/5q3JmF9
Z1jb8l7dZ+yVKb+q4Gkz3gyHb52gbzC25kWgVjHH5pnOH0N//BRPFLxHbMK76tdv6TbzUhQo+O5A
ysHEzU3mBmtLi2maPmdx+qsTQJzdJOQRHGJnAxsUWBCRve0sdLdT4jf/UplzjlDC4Kpxzak4X4Ky
o+WFMVeBHeaeNEJ7KTQyOg8C58KqnZOXgzPZTax2q5o8gv0oB0VaE9B1g1AUtuojmx9kudpx4tta
RI5zHl1mhi0ysXiLMv4f4rGY/shSy0L0bgI3RlUr91ui9g8mtP9bmipPza5R5VYhmH18qj12JqX1
dAWs36HTTNWITg64ZCkG1ZbB2lSc5B+AbgXmURqtzWrlYbPA9c06zOlbM19mt3j8Sk8TwJ/AYbSg
os949hPgZUThbx84/r4bZAqhGieTBXc49jv2q1hOQcKqCQm4y9DxQbiu+m8cB4JqlKgjZjpjMjC4
gfO+4AjnO1StyFpSR6b2bWffIPNJWmXkbL/QOENrhG76NS1PqAsi9w264phoZ1nqCRGmRPDUJZl7
DPD8HbRcwoQCW6iVX96oMHMlSJMa5hFFn9iAp55mZw4WCu2hpar1EawU3QCbsugn2NJO/e8yW7LN
53/1oOotnfRsVQCk9KjCgjZiykumRvICSpX7K7r6RHwmYobeazofc0CiMfW+ucLruAttOi8gsmP2
sdg0KD0wKjLHvrBnvOZwOaTtltC+vuSu5Aznj+9IeDfw5aWoMlwyhhomHp1zGDWF+rjQ8PqwKbJH
05B3a1NDL7S0vipG1Mtmqf/8pRCTmtJIh2jZ4BXbiN1lSwYt3m1bSUpsraO9TTpuggXDugUJslQn
x4DzEBD9tqSMVTlUY1V4bVLHhFTpJIbRzxaLr4Y/73FYh6w3rIxyNW0OxXN1UkDcBM7y1kHZK94F
ckqb6s1D+5/hgoVB3okPwKovQgp0mgAiB3U6aJ+0BM5O4jk65/quIOljuvcn1dPRWdPwMTPB90vw
hDLpTMfL06cYWxjbgoenwwVqmtIMJGkuHZ/amIy5ACq3zxy9AviEdnnQ3eA1VBSSyAS6iYm+P/XQ
lCXgpwpxPmMXfIxxYFfYMRxvXCmakFcwg9Y01KNZD4m/vQKbPLnJG5LdFeWPdADydsQ1J9/ueAzZ
MC6Kcyq4tagu/9fdx0V8fOaSe3GNmG+pHNUhPK8eCyK+Sg2HFmqMHQ99n18h/wJd8OgYkd9bNHdf
Pe7fWvAx/RLzxIsvQT9vJmEgkmG4wPLVMDkFvqAtxNBxP76Vw/a+1PDHUo3x3VGmhOd6R/35LWoW
O5EDxtlY6wSxsoNFPTAniMUNtV/sve4kpuItGetJ3RzZfF2RRDCZX0CGLkw8/GK5gstG5p2b70rT
5yILUG6Fid75p2rU6AvH4pYnf4a6OQaSDIGx5BQSs2ySBltv//o90lBeTUW6zSVsOPrDSAt18YoD
RKOIYgY1fnmHvuFwcVUyEIOOiseh7K+BoZh0M7DS1W9nw4EDiLhTcAUPOlulwInpaQyZzZrZ+44R
3v6xu7DincWjZ3Es7CA3pkgZpHqhoEM2TOCFLZS/AUbJK6e5YUL+tKOGzB+DotLYtH/dENOGwhKJ
vVnA9XXgIQkSaW7N7GRWzk1F66cXqXivDFoHY+dXDSFl09wLfIzY0YSZ5+b7yCWhSqOBt3+FuVcR
4uJTbWtI8L0yox6V+Qos9+wXvx/5Zl5BxNIlrnFpZ5liWqznlNJsq5Sw3jCNUlOXKvriZwQuOfTY
ptR8nViV6cqvIAiwTxxmJlYpWvX1plZ7bABvAbQvjcFqopSTB3YGWRORNQI6It+uueJPRmPNK4n+
HQl+Se/2KJPBiY0g//w9M0Sh+ece9hgPr0jV42vTPqb8tkIeWhlBoeDdavbKwuqzPbjqaFTs8Mxg
iEc23wZW3YBgrCTOhkbP3CR2vflKNReSWeYGfUNCpOxKYRHwJLYUdJhZEsS1BK2Ppd2Qoxbl4t6e
sk5dqHdmcO9Ie0FbTDOdQOIlAMz8uwRPuCBNPlwZ+0xx1eUCsbAD8ClYAggonD3s8knEeGXKCyUR
kGYnATqpPTAONFs8kPiQAO7OGiJ7wVf5lLd81zDfx/xOgX6wgq3u1SDhJ9UR2kjUYRmBSJqDCAIe
59gjHR3s0kV/3HIkf14smxn0OZvIlxvET/Klg/j0v/ViytFiyOXxOMJLw4+Yf3unaW8z7IMTdSGL
AImvU5H1+a1TPYl0JTbQB6FoOaben8YUXrMjSJ7QDa2ytRpoO8q4295gomn5eFloBS0SEOIVVh8I
sltiQYdo/FPLoUWXR8etdzhiYgoUDQNEjXaGP7UbmqOAEpK/SwVP3Ehi8VlYEKKS1O4ZXIdtR1FH
QwWrUV1+zto3YXm/qOohIxGY5qiUz5+ToEYFNicZUMG528hd2+YuZZG0hMrPVMan/76AQ6UlOg0e
MlLH6FAPwO2PkWWPAABPYahl5AKG6wka1QOY3w2r9XElOiTwKpkdOo2rdOMRYYvtrEIuJjM8uNtM
/gJ1tQxRU3pqyw4laKeCN5zOk3n/PKHHAYaA/+ukBwLzzb+QJ9srb28eenQANTSMtTbZVFqaCrdt
uDFSz7a4+jqeiFbAgb0g0vAi6d6xWlbJJ8IeQ6Y3fljy3Wl6jbCINhxczVjHUFaSkOxA/0DgsTLn
BjgR2s7lpeLg+dPeRmW2NjFbmDkedJ7L/MCH0VLgVZV//gbjVXI0w1PRGWoCTOMU7wf3MlxEgeGR
6kx1QNVESJBGeJ2KN9JB8zcqF6KaKR0oSlnNwKteBr5dCJjgFs3UgZ98TijOb3D4lt31yylen0gW
3rYgbX9w9QyHxCqQdhU0jRwZnf7lE89B1YfBvfcpIFMpvG5dum8n0L92+3CsLUsnmg/6NOqKtuC5
D9jBQwaTpsCr4jbdYbM5LDppnwr2bcTeXBfkvoMA+5PKp8MvncQQ4mUp5aQVl82MUtdlVEGhO6vB
enTQoU6jUYO3bP9YwtnUZUJZwStbigy2kfrUIkyhU5AUklcp1AeKsxCd5/t/4w3zp43p+2sabUZ6
9mv6M5wsKVrmqv4Y/r2qNuHdYZX8AWiT6ls6mGzcBxc6yVYVEr5yg8Dz5cBO7in0yjlsMrIxMsfy
ipTlqHfItPhwlACvrACP39g3EP8ufFE3KeIfID8u0zfutgVZmalCr+bTP5vgZoHaJRV0EOGjt6eL
AjzPelDpw3Anvx78LMyQORP1V5gtme9Zv7NH1At8/T7kPo8PGqYD74TZjX0P1AYdDxvxVtjbb+tE
8htMJRVVQvGN7SO2wrew5lGkFNqFtCfAbxXo8z7o7gVKGzt0Hp+GLt4kRHTYvrDvqXAj8Kf5Rue7
6WCsi4iiPra2JJvPG96iI592ixcjKvnL8H/lxnKaC0+83OmcIDIoIE3jnqE1QDAKXRNe4S5m16C1
SzGO49iOMTQhAprKV/isB1+C8ShSr1a6r9Kmu6bO+Fb8i2MkCvPgH27O8lpgaFZrEudgITW92VgF
axoaU3REHw+CZ9RCSuB37M5B/g7bGeFofiTWOMv0GTeadVBh9V86MLcKIfzhUiPaB8rCC3C0aIFC
pbp/uZ8JqqkN7AVyQ1pKceqZPPDd7l8r0NTsBCnssaT1v2sSYilFFJZQx7k+0caYQ6Os0whRk3rw
yhj64llsZ4sYqK3Rd8b2x7xVyRdFQkv2lKfB1lC1MTZKhLcun74RZRmci22KKR8vS2EXUzIrWJOk
zjuUEgzYzAOSBDme4xB4/hCKXy9T1s+et8/boAMOA51oNVljQvNfJbQNO50XbDKjWcnHrLPtwjvq
lZ1f+LM1DjigSofro8a5Cmdf66w5XpmK4NVczXcQowiujS6YJByMq+/lsPVZ+YF+QjJDhJbma2aa
IpVJIMmjfrY582k+Y0+3ez6OG5fdHuyem2SQ+LTUHFoVdZb40rkpxfJNDPV6cWL7rYpsV22Q3Yjo
RadHBuVE6AiLRn7GAy3ifvkiOby5BkRULidHkcZVvz1IQG8pNRGBvfx4m7z49EzYrDAlmU0NDQ9C
flmrH/mqh3D1O1/PUN//jRz64XsHJqqnhgJN70v+mdJoQrvjN9MFjQAKo+FhvhRN3rzR0ptjmdpB
MigVlpaTr6uCYJ1ExF1zOjCjFpK1U6X6awUkGL4dqOUF8J8dRaxErgClSbpa7FBGgQ6ya2Uz2/oQ
XMOE2k5Cq6/Gk5ltBU45uRxqz6Ep7k2+fiM1HRGsBvQYZD0rIpFapf5k6ngqppTx5XnVs2sD/QHM
lD58Rk5HRi8n4+i3XJl+yXKPNp2xzP9jkEQH3FJ5zvFuxTSyEGUzSY/GJgaar3sX3A7BNFD6MCZS
KYG/sJdYBm4ktYISRP/axEZNqCs8XGZ/mwx1GSROgPGEb59MphD9wl9VT4dqVmexOLHBe+6NyOVM
+KUEOYvEdbw6pnhGmSuJ7xwhDiDzNPkSBRnaFUnSkfUprNpKxHlCavOM0szBJsjiNnYQWZFqcbtw
56uEN4Ynqu8UuFyg4HWgRha1H9QwZCHfYII2l0sY2FfGtlq/76tjum7eEZVls7tUUkU0t8LJWQlJ
86rcxLKXVMSY6/2qa+IoDukNkTlsCq8hNJI4EB2T0zSuYiH4zoT7Pj3Qy5UlE1ns7VhwDPxlGaFm
y8AylvhabRvRynpXKMIFBccRLc3ZRw2Tu5vI7072jbjxIK21KWKG0VN0e9IbrF9hiS/VSpl1Nfqu
LKcmFpGOGHoY+htve25LzogwGB92EKHZxkUuiY8VthKYWH49FbHRnAZHyd8iot/fKShdI9yrrCsn
51srC3BhqM86o8aDT/jVL2MAp6D+b4XcGK1AePTan+sIDnlzhJUd3wnHQ3QBZtrAHPyXbFP9yWDj
eplAxNMJqbHaUIp+tmQpq7hUCFZ9FSo2ZVEItjJVewIyXNG/nGBDY4HLTBkIqcwOlslcAmCVr6y6
wEhYV9H6c9ox3WCeesdJJj9a/GWQrdDlCM+qYs0BRhw+jdKLJVeZH0tbvDdX6pnbN5aAl6qENUzE
MgTSBRYhnVMtPeiCfYRjv0IoEHBnC0t6N/e3M2wp2E8u8OW2moI6tcoTnTtvOyiEcJFmslnENced
2zD/Crqh4oEHu1caKlWZ4gUThMJDRyDuQwvwzvgIuYUAEQNGmHDIUJzG7tbHK1/Jy5Up1UcIlI1U
BukI/W96SoBiyFE6xYbope9cFGqOH/F2rtXKomePi0XoALYqS5I8RNfILQOatJ6gUYQFQ4JHUFb5
wwiHVmCD425JtidVIDACm0KcAvXwbnOdfxgHpmwf854juYmhtx96kZgC2ZMl3yJHlhyHcEouN+uo
rYdUbgHk/TVj4QzYX2wUK4+r1SAPzzln1AMM1zTB8tMq2uSy8XDygpOiuYhHxWrRc2B9br9e3Gxb
Vbq6eYj5jfEIgZECxNqBo3fpTOlWvbjBUBdn3sGhPYdZPb/lwERbJ9qnk5FVsZtPIuIxCpK3dri+
8bsjJE3u8wsHYg0caQ==
`protect end_protected
