`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect begin_commonblock
`protect control error_handling = "delegated"
`protect control runtime_visibility = "delegated"
`protect control child_visibility = "delegated"
`protect control decryption = (activity==simulation)? "false" : "true"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
ZR8V0zJd8TtLm5a/lTyEa9whXHmd4l2tlUsSrfsrchXIjHHzFnqZwz7pB78BdALmC0rf655u2QDp
2ZQSU6YLcdpI2jY8C7ruSSQC0alMqLUG12wCzJreuUc8ai0UQhopjIT8yg48IX0OmqN9jJHgCtdk
Rd0GZELOXeVryNtX7sqnUeDhPt/ifO41AdlIwvCDPpohtl5yke4iF4H94ACWS54G1+gJXNYPWXjX
dOxlxxalY13ikQTO9OkoqT8wZVNnvpBcZ8Y5WFin+E5G1XEUnH8YFu0NjRQbZeiMQseVulWChrsd
dBF3whkp95k3XFsKRVpY3OW2Ct9ZB1JAVCGvFg==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect control xilinx_enable_netlist_export = "true"
`protect control xilinx_enable_bitstream = "true"
`protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`protect end_toolblock="jpzFg5pT42C0yu7J91ACfR30CfKR5ChPl4CzKwgHL9Y="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19936)
`protect data_block
uFFpdGbgT2ge2LOhP7+fMjeWfLePV+Xj8lbNBVg97KqjbOuVCNG0GS4FmgBbdvc03vXl2soHLwuv
0REZVgF/ChGOJ6nMT9IeISgqiW1O1qidgp/0NCDEkSJTufgXlIw6L92+rOiRHpgodqv0l6YDLWMJ
Lm7L8M87UopLJlmqCcMcXRFzgjr/LroQiDT6HrQ1MNiSrkJicSrVRTaRUsdXQmrcp8XPRyi1JB//
Dyic3lv1OrevLShQDbQxAvdVlVa50tHbvFWOwR1iQOFpQAOHK8JI135eA1b/lokolcGG97Z9+h9I
M3c5fJIJHSZLZD30MRzYW4S374laz3IdURBypMv5fhdFqxwLvsXsHP/VM5UUYpk1/U+uyH+SFjrw
/7xlG+eUSaL6y8PP1R02NwANJ3zaEf8K98V32HAlv5BOhIDl3lbaXoc4TawCSKdciw1/FqSMPQX6
8d1N5IMndBl5ue686TIKVTfXedh8tXbnRpKF1lfcp9Oo/ArsiV5Biwa1NFQK2GScUOr3/CJFdLaf
aItL2U3HKaIZMNdj5m6iQfWDBYE+Q8PVgA28DCHtGh9EtjR01EqkKu1lJLNwSqZFQZKVPZA9GBcQ
t/4yi4jAdBucjd5L7B71zotmqAtRpzPuYMngD6Qb0LwIPQ61rrLk8lxXKrLEY+mMjFo4K4J7ho+R
w1UalepjB+GwpaohATV0OqhiZoeqhLa8mP3FNLPy4oAMtrJRSLu7xrCt5Pn6wMhrPRgkpHeK6FVd
b071wWsVkw+/GM/D5w7zZLW2ivAOAk5RKL8ok6UdX5rtPAr+NytAXZ/oC/LkB8gz7e0P2u7N81RW
BwQY51JZmhGeh8l2g/ybk3nHISBB8oDtB5l/ERKrPhCx5rKV6NuNDpx/KjsyQy8iEcKWjH6oFv9x
QaLNdhwffEzQG+u1aKhpNqGDFkNskdTrAfq7WNtpVcNYowNDO5J9kplENx/BjoBWJzm93Fj1i6HJ
NaDONhIT3bKjITx50/MQWVaOetBuBFqvS7rDSmCyTQ9acPAQ03qXlnI8HLkUnT2we+KEHMvWcdTH
lxMu+kDnn+cV+M6kwUONyemO1ZMcXofQWFwV4HQU/SHUxL+iPF4xAtLlcgcUOFYuCtqIhh88Pa7v
VGTiPauRGT5cgwK4v2gJCCXIgc5eUPg9nNDy1uxrUKw2M4mrBbPImY4V6NMelfRL3vOoCtjHKUvo
Hz5JPx6wiAXPHSCzNE78OhJQi/HJ1tMBb2tpB+0fWQy9HJ7IIa+3VMA++czZottl6bKLYQXLCZsO
LHeKJBsa3af2dkaUbc0QeQvFxnUE9nrBlEQ3BTEkaOP+QB5782Cn09i020BKzks7t93bWWgaUL6g
a/G6x6EpkLZc/q5NIQF9HEO4B/vui7TmJq5u4+OoZ0UOw72+u9PcE1M9I2bGddT5g5+hA7lOK74R
FuRx+Gb/NhBVBg1Q3/CuwwGtjFGwAoWvoqmq3iSiVS/rVmkQJV0MYCUhhkVaXAkqLJWeVVAijFOZ
WZCrefEtOACasKVKrlEMCg8THOBD7sj1QTkQ7BcyLOL3hyCYCVec4Uj/TuaNZF2m1kdbjD7FJpN9
FqzlkqiDoza6FlDS6NNgHty+w4G+dRTf3DK8Yr4FxS4QuR+JzjDoKugYetR+xzi7FoDKh0uO+8+u
wiSHUfb/LJcgk5UX02Enxw4fvz0I+4rQzAuvhnzJn35PnhRf/md4dmfu+IzyYKSJf57Z03DNlE0D
WGC9Yi9IB+8Gh0VNuYgdzmG/n74HswGAmfok+2IDltMWXUkUyVHfzDDwFDipEzlxiCHCCNvO2hBI
iB/p1sfOG7oxTNoszam/oHIYLWcIjpu6hNP1jkEgfdSmf9dzZX49SddkFlyzHstSC9RAkxGJ1c8W
kcXetBKVljCVw4zNn+I7DEHizVzhE7VIr80F3IiaV05IQEJU1u8HWbpXkG8EkaBk8aX2m29vUqMS
xYsQcnIQ8PXnejB77/8xOGa7fPqj+qHih69yCCar+jMfiGkSZ0jQnhvBoDnX9X9F/sHXJNb1NKA6
+rAbjojBx1D4bPathQhSfyCZktxSuA3fDPozeBxYiwrLIpCM+whUXcfv5FrJydEJiA4O2FRGG1lT
tphMf70tZRL5FxXw5uKSznvrWBAanl/+QeES3vKzuOYnQ4NLLoBbTlvErnhdHIaBK3xunANrZnu2
EvSdcONkcjXnYHKwaE/vwUTqax/8qwV5RPRot/Il6jPYQfG8DFPf4k84sBa4xVSr+et5c2dcZ60f
XP7q6RiWZf6u8Rz5LPi4EQonWnOku4g7ebgWj5hy1KymfSo5aeSS32KJMN70RlttNHw3PEsLHE3e
pHHaWU00rYrXAWvtghiU1OHUH1NaQgvpSj5VCxAYJYjDtrqJwTRJGGaUkvQQgzcbfqKw2JXVabdO
y5Bbz56VWD49Y0yRPa53MiHtGzloW6O2pwgOBcw4dEnGFyQXvM/aeNHTvLNmEcY4d+NZ9KG9oJx+
m+WBbgUeVvB6gnFku5LtFNyxf5Cac9ZenU/QmAOjbheMv483nfZExLaSQsdYMArtq1OS8XvaGUNK
aqurAjSf0Mg2CriZHTYczgs6arBxv13JTBn7ze1Uq/dSqcWbKVfkj+H+ekuxbosHvj3qajMRcUSK
opOoyrCX+nCC84S2zpwhp769sz52NjgnV1xCb6/STu9XkGPTxFgnhFcy7g1XgokOcMlI/AyH+7wt
nBNdHkbmT/pf3fw+T5WAXlp3O1bklLRevBiAOz5TuqUsZN+WbSZGSbwCjOPHrSbrAzu3oMAx6y+6
O7w3OrYwmidaWWYLjRwUEi7nhzCZweAVLPw/t+hBxj1i6OnEx6fptt4t8FOJ4gffSMel3zPi4vDh
I4bMs8ZFoyGQgYJsz+AOyAu/vhZ/rBQ9gp/JEcny4JOTg0tC16+sRcA0TlFC+c6AlpecO8MtuG9Z
8vNkl4estATaDpK1tqqxgQ+3Fx+fUz94YbOwMrBlriabc5LsmXqd3P4huywojc6vakppvsl3kiyG
YhKnqNmVhkQC4qF8gx18POPgdT20JvkQ/Tm+pGlC/l3XOmY/PPx0Dtg6wSetMQ5Bkyz1TY0Q31T8
krwgxIYsPJtTfqhfZeIf6/MU7lGh92Xt0W45nWdUsuAp65jMxszA8GoKIH3RtUsFQt3HxNQ5WJGM
uzbexeI2j+tuhKSes5E6UAt9ZEIBowg+hNbl/KSY/bEQcI7Lqpb+09C+jeFELRimD0nA65XaP2h4
I04thkqASHI3V5SaqApQR88OWaSzMClQOFCfYZKVs+WHsOBzzeoWqDQ/JI99zMRlVEU0Up6H2y0p
pwADvXFYAJAUpJAJClmYK5LN978/90l6RILkmskb4hljZze44zWDLWtDve7dzyXf+Q1TIFZM396I
wkzVi1Ch+ht60cORDPb9dX9upgmPew/kNauCVfM0RLkEryBIhjrDCN74GYWhK0+VYFGb9J4KN9oA
NJbWz1OKP5Rilb4FHofCaZV7/UNez0fD6F8rsxkce+fFy1Lo5eQLeLjAesBd8TuOcO9zqZK1wiFy
Y7bZk4QZL5ooWHACVLaPxz6iRP69chGHn6LsEwnqXyiBffF9ZcBJls5BiBZbkkAaVQH6ZPE+CUr3
3TS58Y0Vc33To3PbijKgiq/xsZ3AM71mfimDNfoG5D+VSwIgM2ExUeY8xLGbWL8psW/PoKk7V5Zr
JXGjUV8C70qM8ubBWcD3VPkL3hi63efKmtV0nVvoMxswhXQSgGRCt3xA4+XhvYEJ+1XfFmKNpfHy
bE0XooGvmVPXSplFsATbmHR617++MNIa45/iZ+SyGbf8LFuVAqG5HMJCl9tgIo0qgtFIOb1SbN8c
6ow0Nf5BRsXxBLbbLHh6jKdF2le4cRVuwfCVb5cGMCv35RBrOs4pAx6DM+ZRlXO4REOhL9lQ/IX9
nxn/CXHMqcoTMMOX+5e/WDrEGrom47J4qtzE/9LGpettaX8nhcyagGwEzy/zQ+wM0HPKvSpd5tfv
c4RFdKQirTYQVnMkmBNYYskHXWyDwkJyhxMcBD9YMQzySmrxm1fuTj6aGUwE4ERu3oq0BzGs8pVl
Ol7uqg61Abg3fFYXWAvPOYF2OyJPzZrOrohTuUhKVNOCtLsIKyKffCQmkNaOE4B1efxL48z+CnSs
27uvv5J5e/z9tKX5MLL8mRIotTlXTEE9j4y1tXHATX08LEXyIar8+8RFD+5QFWaBJPr6iVV0OvC5
EugrOjfnvOMQxUsw8Ky+GAVkpRWOQMMhSW5VnF1K04zKR4XQdl10DTZ5hmj+mnTPYaiWqhoXHv+p
KnwKhq823I0x3xBK562DHTsdka/OAEHRV728wQ4DvFJj/dVtRTHXy2lt9a+3S4aerDDkzIF5L2QS
MG2ytYDumXTL0nEO/RWVMwUIpzq238CSjUqaAnnIV/0JntSHDSNqbnvJ/5yU+fjrb5eMKJ++sEj3
yOxwj1USm7hjYGrPEnPZMtgeWtwo0bLM3cR2CufaNEVmUofBJOsEN0Ubvq9tw89+tBI86okttpfm
6EPKW9zAEnIe2WAgaJ+qKfeM4POVdPco3gdHDCaGU2ptKFeXmtSJ21REECUoAWZ9R3EqBmfyVOrf
l8+vu+Ai5LIcPn72KjMkNTswPrx6P8x6oxe51NyCHy4+gW7kXYZrNhBKSKHc0YaFI9HWJhMi0a99
qemnHcFM3Bbwy5iDF5uCY4BXRnN7ktcWDvqlISelGTA+cvN/r92MUMOBhgwg234mzmofpuwV7Kqz
jdHrALJUNuPonPXewBf4hs+F2wkAY56/YBfx+o3g0u96CbxUSHZ0qsyCfL+5epP80OoyyVHz88W9
1aFKA4G5yv/ixFF1vfn8nmTkwYqC2oz6t9vxe5VmqJo7WDtfysY1c5MK4oIR/gh5WZKbNRleHqoh
pMZdkrgoEwztHWyAN8asX+Nzg6ly061FOaXMFpGMLf9j6gXI7kYCebk5DRXxekiHhIJ5XA1DZgcj
nkOcuTTO2bYomFExlPhydcmJP6VXEEHgTUMP/s3LP+39Y8uW4/bRI2lwT6J4s2PcO41z1NbaxmUP
FvLgAyqbbO3JMFnvWGC3Ky1t2hwAH01ViJzFHZSAJQyKy+XVdP8tX6Wr43dupmDLMGlDcz2PjJ2d
n3Lselb2zxNUJvF27/L64dXMmGAcrJZJvDfTcrZSSrF4PDqR8ScmbV8z3gmC0Te7B7fWqaBGEOjF
c9B+6+bQlTEhtQSUYLBh6gkBtJjCMfdSwEYDQ3zwmyZbki/x4CIUm4Y0JZsAkAQAPrcQQVsZeCWo
dKIlc2nVyygig/fktqBQsIO8eMMHegSxOwJu+E9sH0UbF1hP7/mI2REz7ZjQeg0OQAXHrOZ2t0Tb
wHn+MVK9bKyogrGZP1J6PFEfrfHFab+KcJlXbKr7+ieNrQYaJvZFHlHlGIwjV3rZ9lUSQea+irmv
1IewAQOKka95sL9yxf1R7wUsA0gVbYOcgPIUrJpNO3eOF84Z2Yzfi7BmFveD5VGq6VbTMT1DvlRe
vzG/+JMdu0yPU2JmiLyVb6+pvppV1ec71u7dppiEQ1kA1lcwbLgtweD/83QHsTobf9C19jutAd8s
yDCePG7Wqm3jxzePEh68PMsYrdHcazxYN4KvK7+BNkfUpp95GrICk49ei21e5/0/ePDphLsxM0Ap
DPFIJVjGKYF9cEoTZqlVEKxXMsWvzZJ24+Pw6w2jMPWquX/bUAh637UQRuxzxkHq3gQIf8fPuqic
9vhLpMmH84E/5nwcd5cbAmR09e6lctZbtSSAXcT4/EJIe02BTsyDPVdQqeAS9tExCek65ezA9v1g
0DYooOHZpdKsDnx3VKyZs81R8ejk0md2UH1AXgEwQmQSWl4XXR/xQ6fslp85QKrh1odzphjpoP60
bs3z2TU6tlZUJQRE17NuxJ4mesgdvHougVutuLp+SoM8DBXg1eCvhEOjHd8LoajJ2jYGe3vCd34e
eXL3O9zJFipyHICwKaH7wviJL6buMJPU3/Lwo9xKoiPQS4W3eeHAislaaY5cpnTcPEuhcDzfcI5D
aJNvSxfalAGEXd6lAna8JbsdviqzfIA3Xw2UxFso7JHg6exLL88/VqXRGhxT/WgQ7CKZx5BZmGAQ
V7Wn/2vHoKzbe7HEvPGE9lFSvpg+HT/bO3I2ssHO0e9RyTIuER25+hemd4w2qn8Bdx3+ED0XE35F
thuGqQ4JtDL85Qg9lXNnUKpIpbCnEJ90+jHQbmE8wUlI/o+9WwJVIaA6HDJ2Nwa282ibSXvW4H9Q
i51ojJsWX5nx8DYQWx/I3H7HUOzHHVtjRKqEv+nfz15ib/LATb5DDNt5ntFKamJxA/EbGRoW5yZQ
0SYrUnj/j4XR+9wuieMwT/iZN1R8f5imS9vhe4yVxqpBVMeHKBFfr37MePI3EiayrlHx8/49P55u
95MGJvATXJpXP0z+q/DQNI2qkeN70+Ey7m8b7nzxKjmthQMulYfUc9KBBkAlW3ypqW451VDIA6By
gZNpQRC1dI9jeRKFyKp2lxEWnC5M/ZgQQWBZdghXLtHivIYM1f2+XnXexSWVKcsjyrPJ2RyAJ6TW
kHtzHtRil3o0mtnXsOs6xldc2sHP1JQrw9XwXXIKoZ7o3acadUscXDN7iWqFuChY+CKgqBY0GlC1
tLyc0wUCLG9iwAZfOsQ8wV3p/Vv4jD4aFO592n+ZvrvFEbCjOyp2OoMUdgiDqyaDj/rCbMdQ3Nal
58LvKre1FO+hORP+jI72DQoMyXb7a+2KUe67fE0LKaEuAinhWVMzw0GetM9GOUAP3NuJYPQs6mFb
G4fyyLbmI8CZ/kknxZOa3Q9f3+eO4B9q9R0UDwAz2PCNOyD+6BlouGUA2r/gtMs6yLnle1grFZj/
+Md1bkrjHFFBFe1sdt80QTn98s/0SdM4PzXdqksYJksgpc8f555xpGsVGNMpI7kOBkOX2WKr4n+W
VLoCudXizZxeNO9VzNNWyz+xHXZqzkDpK6ybhkPlehMz87za4qz/rTk8maxMJtpmgW80+2h2nRsk
M+SXfTr+dk544TRESYU8RTl2EQMfHZf6k/I0dMqL3ykUCm2eTCeg7WqWuzwh9+pkfUQJik4MNxZu
90nC1ynvUdqFIt9f+rvPC/nIedt6V5Dpcgh4elPM7ErGA6LVgIgPGbEAYBa2Xdn8azYxxPn8A75W
WsRCIY4vmZ6KdnpRzDN6HFBI6YTUkVkjpF8fyNou7JR8WqKR9SMRUpvBnCS+hYHVexseJjXgeDNT
dTQTfwljwhLaCuBNbepa0jZbTewMfUDTiafWLZDm3DRCiI5JYU9Gl2pdf6Q3gr3izbK6sa43+qqm
6XXJNlnnLGCLeUpLNpicQYDS/CrsiNx2/MW+62+2TIy6n6I0bg050RjBdaaS2A05KwUIs1cg7qC1
+pLRdvxW5E35EP/9w2At4xo60wOM1gfcoy9NqlVGoXHKsflYsGrnterTjiJP78fHnhZ5Sncn+rtF
QH75747P9qVPf9sGmA/cMB6tomcaS2OfB7ok98QMSfjnQQwjBbXIrJ/F8zYZsbJv8KzbN6EwV7IF
mpMmSY7BwtKwnHbV6jeeYbUggoKLASpRZiVVjkE2ijkm4UAsArkSf0o5k/CbEfIdBP2e5EuEYlMj
iPNZhavqOlzJDIL3IlSl8foQxKMUOb+ze0UbgWN5hlw24y1CrTyQmBoMiXhHPsEuMIRvYIn/WhzY
d9bXEQ+ptMWW7XU6uCv+REceukNkLdtS2XAWbslWLSNIXQ/JIJ6iQHV0gT3eVeCKSm1vWJ0VdjyD
heS/dCr3dTGo4KNgVQ2Rbwb1OJZa+i0YWCizqovH4d+Ilk8saO4vTStj8phfP/s3tC2DchR5FUT8
L3l45weEM7PauKuigDflODeKGjQyY4he7yTMM+5wkrxrrHok9xnttOXDeTdLjAvAqcToHc3ywXes
1fXmXSy1nUKITdFCpv1WzWZoD3vzVjNnjMrf3KnmiiF8cIriLxEdjGkQoIIMWjBUQCHPQvCLUva2
b4tjWe7BDGIx6NtTbN9ps3anjasNDikUyYxC8YUt25oQCzjEtXe3tPGywXrFGALRpLDxLut75ak0
xsBP2k7t/4iPhp2YR2B5Fh+GbQofqKLB+kxle5roWdAsrxglTmKLMon7mgGL4dtL7tir+mdMyfIt
GrhqEOiN0JB9CvQGV8opLIp3tR2od/24UBtCD2LeDW2eNRDpYA5gUHsxcQzPn3FL5gtz8Z0LUzsL
X9OMxgNLmZ9XlG04aFF1l8uGLwZ0uGdOVZ7ilxyqnUMM7MtrFgoHw8ne+jRmHHzaQCr5mN2wM0u9
UPOIlbi48gSKtCgFOsepBq3ryxhx4uLJmBaENFQdcBY9ap8sFZ9B+rHOEefT1eFjjJW8T9YfV525
pSypIB1de0GGtxuy1wLvRkdnutB5b/mw0FhCZB21cSeWG8/mJ4z+6NTNW3ipMWln3/ZLEUf5DJfz
h0CqXcnR6QW6xBIbi2D5whdrl6suJhJjF/7vYEC9r+kbNZIK2CMtTquMJXnbN2TrDqeryBxSBoRj
hnTQnBv10VIfduTYb/n2XJ3eNg0fwLy+5XtFGcCDh5k8e+4teb/34Yz0wK4UomAGP7dDc9OiD8HN
Y88POK0l3n+Gz06ntcawuSmmOx1S0nnjSUm6jyxQHMeywk5Ytd58Os7o7W/RkVxgEFd9k+sjkLjX
XWta8ugFaXpnUtjxSEkBlg8sXG4y1ckEErtZPLHRqcgBr/ay8InOvyggtBW1vPh8JpWBOMfKVCMe
hZ19/60Szn7oOqRwQoLiseEfuInmUsGPS33I3lHztyh0oZX8sif7LYBQIcwYI9hdZ6HIM3956Rlm
i9QNaDc/hJHb1L7DkbPzIn+pM+LWB4MgQ9urdJu84sXHjkvAR/VHEL/Ky/PsINPTsvwYLZT3dxvu
ZwMl2VovHwwgA5nPwacpMWddU4OAR28hUqJmuwbY4FsKALTcjlvnQa4QkefMENvIPLYL4Qps4n3F
9YnrbJ/BHAadFOP5uELox1OmMp2M5/5mIHZXydiCOVajnb24yv/TMrPOccozoh1/YKEWQ+GE01x4
Z9oHHcCGb+zwEGSCEkatxV1NGN956wYjX0iYAiSkOYwOlbSGQys2Gvrp4/kDJX4pG0NOeCdYtLVN
91TbbP1WUBMbsmo1IicbAtxOOiJANmkXZN/6hm+lBDuzz57Zq6nF5ATihrFUuMw8n7PM2HTo0pUk
5PhF6iSiizjO982eJgoqODdoU4p93riWdj2WjtpQuxkfVKTx3c53a+Uy/skGZBIi/aOuJHtdT5J2
4/GCxTabCiBfPo58DOdryTM8ky43NzRal9qP406ZPe1k+gu3iWitzwz3yNljjObTptj6Of58d47R
pWj75A56A+MSTOErgmV6xxv6wyG6k42BadEVK6/Sam1j95L14S5O1NsbNG/UFmnslXb0hgwr5AVe
izPgyz0BIfdnzGUvUh3GgLBGdsJuglT8KVu0q/2r8cBqj9KpAAmI/sHz8hM9rsG+ks8PiltrnSVN
2EP/wKzx7iRJnvFTqboDlT3bAy4J7w9z33o8iLKHwAYAJdig1RSIcp9D14eZ2arzHCWTraoWoDrv
bADwDQOHKlcxJB7JKbIiBhNjM3gPFK0UKxZxtusEw7SS1Pdf5vHh5B1DEWQFiB5mNH5C29FVqIVu
A8sN9Qk9oMjgYB8GHjoAW8p6ZQWLpxr80IRolAlKZzVl28QqFVr3qOr2pvhKnzbIKU9HX4aU3YHH
ZMomG+ly6lVAoCl9IeKSd1N+uLBOdD6yJRcQjM6weciDwyf1aSnILa8zKKCcTNONE57iOji10EB/
1jWZCIup33adgXf4fgNSuX0xllEcTRolcBwqUzFmBnZJK75SkDi+19LV0/1K0+SsiAp4WZ/MnHHt
MEKvtDeoEe5YptHpcIKvilKOY+T3htq71e9QLPUny8BGm6uPpCOkLFhXtdn+0rV4dRmxT01f8ynh
vkpbN33KhBOSR3KOxh1zfgJnpNuGp8UKXqUeIccL+8ERKPg8f9AI096EgvVp4DxXqeS7J0Uj+DaZ
EAUQwws8wCZmkyYFzVfWx2GUQOXTmJVMjhOatmHEvM1WpVIweidcqKwhEUFpUsc1+KYHqOPByswd
KLu6Onnl9od1adTb6Cdd+ls1XwXOD8cXZw6Mnv384tGd+QMrRiXzBnfegGe4fogJGZUvIefhDWoZ
Ldv4+NxrK8TEBSuW7H96KQTmX8oA2ffwX1OCmuj12Tlwce7kBJzo6TieuLM8r41qzpG3p4wttEXf
VT3sZuNLs2FbcX81t34o0uNXtFtv910g4ryqSAdPLJzkgSKsuCFzbP72fX1gfb7ncZxwVoFWt7AE
FG8Vxd7iO7N3Wh1VdMqSMtHhC+m45KGccVRVQRqdeW1t5Rlyf4gE+1JnvkMpIZNjPW+iNMBEUEjd
xvpxss4b7gFb6u+rVWU6yGcW4sODv7hjD4CTK5O2MCTIRSUtuxGBC2zumZ5Lx+up/Vm1u0iMDdrI
TL88KQoYoakKRmZb0sQFcwkkmFOxrfOEY29aCMtHftY1YCBjJF7B/z17d2FB9xuwJtrD0aonDZ7a
QLlJ9NzS8VijD6Q4SmgfQNbnE1vFITh7+qkfy1KxsjBWN4+zRdSdgb0VwsveJwGj+EiC2pMwn2n1
Vo8bm8MxgG8yhLZWK3N8tDEiq5Q5XyRvOnuO0Z/HKHco96jR4QbmmsKv8ADHj6zGEUm+yGoGYS7O
grP6poLpwD58WAkvIWbCSONwlIniEkEB/DK+a9SLe03Y6XAkCgbOyWuMb2+iGbmR/H8SIzNG/C8c
ZOoo1WY9yK9WGu0RxmvjVRfqV7Xxv+hgen/e0fttJKkfIUf79C9am2VVyj37gdWOX5GTxA5oIpGC
ncmnTOI/a1X993/giItzCxddTyzbFSlXDoyEIs7fevYPuhay5IjXah7SnFB0Vx86ky0bptNZrfCQ
v9bk3OHdoo1du2DaGZxVRp6rM44LQd5TNXk/nTOo6vKB6lGRceAqLOf9NCfbqFxXKZUlP+ziInca
gnOtdSKE5OqfXabqlh/tN7kYaanyob5HVERlqzBazLMTi6GqEyq/w3t0Dsa5yl7eljaqKtergS+Y
V+6c/LdJtcm7iFQ89/WQ4jbuUmYIMh7/pjg+0QTnirsIdYOc7edwjXkUfoNjJWaxFEFwcq9q5RRy
KB8cU8aL4jqjoZgvml4B06xbcpCO6luLfStT13FL/MmWsBnYZcSxMYVMWaLAD6DwVl5lwt4WNRUC
cFi6YWuIF4o1i08clHWtpe6YT76kkzOCFPv784l8M9S+RS1P601bwyoXGImh90u8KHQjcb+rsTDT
hE5ZYlYKy9dksdjiZre1GjRqs0/AUjtJkhnst2zyfQ4TnbcFwooUbx02UEkn9G1KfliXYpJNec20
eJdJ4ky7gMfs1ynG9k+cMHMHrsC5YKV5LuQ9UFZzUaWKhCDMObKbnkl7bf7wfovrV7L8Py77/WCP
VgbG2wgyRintxgauxZ7cLbYVosSGDsQOEu9QiWxdWC7ylZMFoTnFWyfXyVTw8o1dlnBwqxC0pWKV
/Vry+vHz0q5MAD8i2pgOAhV9b2CT+foSV/wR0YtZs/od97sE47VqEECaz2p4vY3xZCzv+KMOY2Vi
ozTFHfYJdUiNUuhVGnyKmG66q1XCnOy2icFhoTwhHw358ELOT5fFPeItjejRT9uIgM/Jhu/FDCJ6
aNlj5X7s3FJM/L4RoTIV2mCzyW5X02ggc3ANXI2yIM/ePYNkxYCThrkuX4hk1vllRXN17YDEhANZ
eg4jTRanY6bpnnXqEz+ao4AcJoDAk2eUeFSXVmfuAlzwPD8B31go+ER+hckmB+gH12QES/UjnN8P
HaV+jE0cWoppqGkdm67cgDFIsAqJvglHy38MMwoL1MtS0GGM2mJCmB27XD72d2REWFtdZ70DPAEr
Wb/HXXtRfqr2B0S3Zhs5XtwIwi7Rd+9Xnom93b95U0iqXb/fY0MVn3XxNGr1y5m/nB7X5fzZlz3J
m+yy0rxnX8S7XLAHVh/B0rAd4Zo+mX7DmtW2X6X+DSAEheJurVhZIZ3wKp2b0cIjwHL09M4chXoB
JFYBezn9j5JwHmOejFtL0ZmYNaUjAdF6qptmfEWoVqYKLRj6ZJdifJwxTLg4DmC4HpqwhDFLWOzc
wRcPedIyiCKharIFGNO1QfYzPkTyWVOUYuJC8T2PV7WQfEkMKPIN78AiuCGS0Pb5L9TbeG6MBqVR
gtb1QtbCR7oHsD77lq7GrHE1Rl42PZQ8jthsJ79BlfXzoj2ZqYDhy/5Cqw+LKNHSVIRxsJqq9PoK
ufD1jZvBjU3l/Stm6BnwpieAm9kC74DYIVAj2bRe7IClJr6OON9uHKlKGFfFRoa7Z2zv4nvWdxyL
VIujx0L/LpRuH0G1XKj1HIC8LYyKfb6EwrCKZ+jbm7hH6DHPgWm36lloow86cOZCRTCE2zbW42MH
kCkCxnBZ8pDRkDeQC9O/y6ni6iTGwf9b5dAg6XAxC+g6g9qx7ZCeSlj0122LNiF/tuAxmWEnMx0F
8vu4BZrMSGH01SdFWPMlEyz4bVdwJBSYldg0dp29Vns6ekwwYHwu+2cb+EUmmafodO3j1yRTotcn
fpuuLIq5MvnZEA0NSrPXgwvy0bDIL1dZAGRK0zXPYZFtIML8mSgrSm5HXpyTjDYl61SGXsoxGnNV
qXwP8Qa93XJnNfX9Z9kiwYbXJX9zINQIRGlNVhnknsf+CCWZo5I0+MoghFflpswiuSsRVpOAHynV
Kc2bQZqFZyizEeB2XpK/FCC8p2eJldytzipWGxAjb9hJyQyAJbDV8AaF1i7e+z63v8QpXIVe+YT3
p05EDp76CsynMR/Q9Udi6tnRs0yr4pl1GnjH7W0SWNHqhDWqjQB7HqMGL2kmL1igR/CIXmeCNge/
hbXfaUMdwg0UzCkS111VdVeKtpfgJtRm08JJRXiQIDGBwxA7HlMldnfpZUklNU69POXaVzp0U0s8
hh6NjAboSvG+iwnbqIJsog8n2Wsnb25TAwij2+sqzwLDTKJLpb45JmbPTsbi6wxn8x3ehqEjLSGy
c4uq0fqqd1wnFukfdSILoBoPAwaPBSXOpI8MxCv30Nv01/KnRyIY62erKjSUDZ8C+0iCQtQFXZOp
2IZBm4iJTGA++7MjyAP2aIP+PqgSXKLDXTCmEq8feDKD+ijzeWLh8zob8Zm2NYzCRqkI/reSCLWP
G9J3Z0wxwZ37swq5uFC3MJfKpcnBAalO+i0zOoZGjbV34KGhM5FrXImU5W8VXee5RXPVDhc0Ko3I
33MO7dwvca8wEUNZxCv25i5K4uozV7jgoHCrCZHecjSA1WQ3bvu/0IvkufiCOX4KUTJyx3RQaY7C
lLjefUtEFofHUKHg073OjPvko+5gTzfJTWoMF79zTc3tHhcfMdiLPtb+gW/psTNhZ2LoAc/WWnrE
/kH57ZvRHhJ+wtJPMPXagniI4Grrbkduqh3y56R8h+gtiXgTxM0SrCjE/Jrqd3ZW0M7PelixH9MB
EBg1Vxz+fac7zuKS4jDKuyODcS7y4Tsh6/Scbuq0BviSmPx5POjEhNwiKSxiGiVaQqqFDO04Vxc0
1jpHoXhdCKXd+ccmCkCQk8dcmlaOkV1nXW1+yFsbDyGngrVAX5kGgkawkcz3JTjaoTKfwAeO3BTu
ZUUGygbMP7gSFY8h9paLldXUx4uQQVSRlR9HVAAsWv94wfaoECA5PsF65yi7gEkMxeqESKezoSJU
l03Hgj/b0OqH6mv7vB0c8DaFmEvD7LCRCWPoDSe98irqZ3ma9ubQ/DLcoJAcODlQyfsCY1+g8pC3
kFu7+Hf2+gAsHP26u/5rC5ESavKxBLF4gkuBaV/xZ4n/p4LdwnVkndp8xpxp54M2Dlhsp7tykBdB
EXoCOdtgii09zq9y/cF1VrnFIBObZijI/qenHdReZkdLjbjgPoXqAjdvVEW9HOozCLxyusBwCXO5
SjPb6ne44cGzVSJBCjzRt2BdcSvotrPrkPCAgOMexKPfphSHQrhkk1ZUxUvn7kAvXbF8qwxwGo7X
jsKgf0tCgSKb5dhtBVOuWm0ErZW+2+P0dS4eQbBeRX8C0V6yCcF9OZSpQhYHpvLegNzRxbezWGzf
ZSz8DbDlDOGGRi6U9EiDHnXWAo/9hkAdtOpvpogibdhi7nxhcAnqk8sD4PjJ/gnZz3PDdyBtt2WE
89Ytn46dnuLNo0LpzAE2nqoNiJXOXQ8Dv27/iN492jP4IGhCO0eVup9xAa+V7CH3tkGFrFhTXnDu
J+W492Mi9ACGMJhwKOgQQ2xIjYAs1Y6xfpbjz3tLP4tcWeiVmdxbGzM4SNjoghihQFzav9eM5Ck0
I1yWeYGS05ntKnt4m9DmvhgWWX904wMd1uDsb2BqV+pXFgGIVYARmgsyL1h3jB4Zuy+Eq7bZPuTQ
TO5tCefuf+MfaQlxQ9ES+KI0Pnf9zAegMhMabb1TCReBU8UmxiLRX8ij6WyFPCuNWYaQPl1DDLVo
cC5+TmG/uAJmqNTJYNBTvEI0OimM0Qxy87p4a11IgwDF5jU8BAc8jzxxTz2OrizczPPygBA1uPs0
2x3v9aA/BLuVngrRVN/X4DUHeZA8OBj6VPTnoNsLEkJtrmp0g6eiZVeScpkwOx4g7M6UzXMIeOp8
asTGN790VVNaTg8Jv1RM3qJHAY2ZlqgYvEKyvNmwlZQSEFG7VLK23TZC8kDCaRtfHLkpvsLAVtMA
6sGXty1NWYDxL6CUhYOVgGF9skXmzpzESUZS4yO24z4bFdpQ8lcTGc2G5tmMuJWRVVJEGhXTKv0g
SRFWW8W9fLsiAEcWg+G83qrD3UnRTBvjcx7eC9lQh4+VhIu/vpdk964J5ih3Rdekxk3jxgoxhb+c
MHmujGuHyAi+rer5Pue9hZ983CMLZx0cZWqAc3PxBkdjP6t/YYoc5BmcAjcFgtwtneykE5TTU1dM
zIC5sUXmsbdVxog7WjG14EDwbJMrVXiabLxZymtEstcbuk35yN7G/S6vxnm0Rqk50uYigIyGRXcJ
lrtkCJOelw7RV+eG2RaXRPe3QlLkWIGE/JwzmxX4pcCkXYuxQUFPBe+ka0UwepEsdXcRVu7jtEiW
fCDD8V3TbGXcsSZ5Znet5Ax8u9oH6A0kFA/twNnLxl5/IDVJz6ZrLfR9p1j29tAKgsVWkAsHwr3g
nqg+tnE7KGMEhB4HOfnU7Ecdg2dXRPnBdSvalLdXiBOYtz/D/H6VIheeT/Smir/DRQWhsjmEwy7w
Wvr6ZJ8yZDxOJzgcj3nuXxE8b+BQ6IChOEyxFByMQ2bekoh7vOZnLO3fz53Y+zIyiR2qQsdW5BmP
egMBhVB+xfQwvMEU3wk4RBLnl/mYL2HqxahnVtmP2mP+C7AXRKMEB0WjMxDDK5GikDBWbK3Rpqe3
QarWlsB6JWqx76SuP8CmUHgiVFVehyTdWjRQvyDDgJWqIxdKYpH4yeGGH70xMeZKXRI0ergW/yF5
daXZozxm70SW9jdHOy+DfBbSeNrf+e7qFqpCFAanoQPadWLEIOzCMaWDsH9gr0zhOY4ER+XuLCV9
XGMCHZOeQVlgW3/ubsN0CKwhEe4LI8HXtvldNSBhIJqvb95DhxYowIqn6Tb/ZtkG7cdC5cYZwsPu
kWgRA701l7pTin9lNlvxQqZFysa8A+GeDZ7f6evm5qGnBaCoERGz8nu5Dh/Eimr78pUTNfJ+iQpj
ibU0t09N+LXJaXm9pGqzrIPXVcmhyERY5I1VvWP9SJbioNIPwdGoRU0HHIZ2vXdm8Xhc5kQUOwu3
Pryy3xTMzjw746PHdh4DW08ZnjGr0Z7o1TXn+se1H8a56tmK7mgibN7YFpMlAR/ENGYSR+MTQqFH
Djhk7q3/vvHJ0ehpEKm7y5+rbKg6GPL/yhrpsToYU01jfkEqmHjHEMfPsGOAJH+JKuXKsAGR8+r8
mTyB1ENen4wpEDt/7x6y24E2NVVXwkOf9/o9Xeg8s8JQBc9nWlRm8LGLX7oU+v7QCqAYCHR/ksIs
EGbmwei6xj0XRVc9Vlz+NAn8/iSAQtj7oPh97NUu5e8G2nlTKXyjJtGoWttmgYol3HCPV8V2o6pl
VGB+8sCivtS3Zkmjq2s6agGJZV+Dk3w2fALl5TeA73ftvazkCSZW39as9J/4M1lPHfRQlSrNnLP1
B3oNngd3MnQjaSBl0xHwe5Drl3jz91XNqKlI/W4tYwexnfyKLZY93sNcsMEHwOvYnqd1l2Ccf4Pg
CaYY/Ep55Fj/Ry1YyqeLi9MxSvHgWY1Kl9kyCOFIX8k82HsW5G82l9KRy24FnOSrvsru3LkL3NbF
Qv5I8uz3xOlPTFIA55gSmIO/PdgRt60vK/TQAN7ZPpKtjwQe5Ed1f7P1yKxSB/3vpSzuz/l6djao
3pS0YrVBMGAjwi3tZXB6TZ0Lebbgltnz4R2faLVDgxdRn9ttWfJo/rSFAGWzUjOluIX0GcB2oxrx
QIs0QSS9ZdmoyXaXLVI0mHcVFMIldLc7+3rJeTMY5FbfkWwkpzGWVwZ7hDNGKTsN5SwCWm1kNbJd
bc2ssnN8EAX/TFH/f9fzYHhnNinN9L0I9gzjdlAFXBQJerUx+koTTUlCSSO39qYY+n1tbHa1ieFS
3S38m1vFN3McztWSAPzrL8vZhS5pYQKoNWG0oOLV+Mhr9Cn8d62YUnSubR/0CxVDIraqFBOTCbuj
TEGFId2iWo7EMpUgnRvUlRXJgki7nYqrRx/KrJtF5o+ynAyKLmL8btbkeNw6UvaAIJul3UILcpr4
zkFBBYEcAb1N1hnLsB4ZsxnSt0sci/gKcvPfIzwR2EE16Dn1q9cwbnskOS6TJrGEt59f14OfHWpK
z04xdwtBFgqEEYEvK7dkqWHGkye0QpCLuzHc2tH0i22wjsraleysqOcbd9kUNOZV99fjx8OC4zLE
DrMZxlJp+3jUkwcnPtkRNqjhR//6z//juNPgHfL9B5eKxD0pfn3JHSgDCayaM3cdF8gVq6Byihl6
l4kvT7+kaBK+V/D088Q9+3IcR/z8WyxfdEO2xTcr9Pn81XXiTHidEhGZy61CTToIiGXig+rnbk3R
I661Qe0gD2Evz4UJ96lPdCw9/CmyeVPAlhCweJJ0BGByNe58iJg7S4bRjhPbsB+KsVvk+krooMcz
El2H6Iypc7Gk3tetrLloruoSGlOBy6tDAVA8Aehi/qq6AilpU8+LdoSYIOqhRzdlVlFcOGI3eOrL
PWZuXwA5y2GQCPV0fydaMl/AQdbCFj7qx9XY4xfVagV/E93DU4YZco3LfjPkuxX6s3101QhoRWIf
C8SfuC4z59CKnTBfg3m2k3CV7J50elSkQ5S9IhE/zJAl8dJP2qIc+vfLoTJecD+TJdWKAUypFfEb
ji41zGjuAEiVa9guRhPioY1jnOafOXPWjKtvIsMQaGbSCEr5P9r93sNgbESA7OdHgQInsKj++fpL
8OE29MmT/mLRiZbhAqBc26mBuBtWsoxXXJ6H2JFtFzQe/BuQ7VTV8uxZYa9cUXWZiOTHX8brVmX9
qD1qNv67FF/BbswQ0lW5y1yAMtfhuF7I+9FfCYEMWUI0a+kWJP3VPzLz+ltZ1dkE92L6oFUcoI/B
FEd/o35fUi7COAusvJpb60Ys3cC1addvjT11N0WuVGf5yLUXGDKnzaLP1oT29NW4zydtGN5gff8a
sti5aJyR103EiEwFZ98I/IAC/iaWfAJ+xLh2bBxBOWOEw7aLggTI+0b9puv27x5GDBVZbmj2MfZc
i0q6Ouigqiss2FPhbnucbdaivIMb7dBWgaXVEl++aOegPl3N4k0+9V1AIPEAWR6WXVoAGx88PGIt
HQwQgQQl2QntieAcy/XQEchD449rhvmAuh3OFmYR9BXrRW++PHoNjpC8Ds74o5elHdyz6iUB8jkB
jS0bgWyuJ7a+mKzVtmjV5hgFY/W1t1rYQQ8YSVFTETCUdR7WV81amtAQW7/g2ocQBHyAX1QJ0cfy
wfJRXStigB8OEPgP+dQT/EBkN6yRhxLUWmYzFJvyPNgJZu9eNmPtjb3Jn8/c2hStkrSRV0wuoveX
0zCJqojNktSOOVv167v2rgrcjx1q19lqABVR10RID1koi7NMiaL3b6mbW7Un7Eusx3ojTz1EBuqK
vMJlsnDA50NtZsaV1+ytGQFH4J7x7tya/+62FezNqImqg+h/w64iKXfe4Yr7Wspk1oJHLxxBfr0n
O9y5IzkZXnGkAurYI+eRAqW7T9pb6JKTG76phTa291t0lZbLHr+NC84e2AfGwv0JI8qyA8jLuMN4
imjlNrOE04pYHe3gZfLL+BNdcACxCFav/PE98z95t94mKhm7BCw38O3TRMC8jJusGDR5eDfBJqNT
q6XD4glPAxj5XaKd0Uiv1nafJagjOWujEV1LcDk9gpHlFhIljVaEPqwFNUA1KL2I2GBiFrzn45MN
yfliQ/xQyrLF6dsjEFApHEBRBUwZQb0P2Fn3C1mO3RPSgJn1Usc7EIg4j+iAHxmSG2YsrHlsYqDo
bUvgg8fudHxR3ZXVH8bK2pol40GOcr8zxCLMet7ca3QtpvVctt1pkolCP8zrwovjxsmlozX3qPXH
b0l04N2Uk663MBZoT2HOadK2KEkjQczJ+GBRbYz2jdbL6ocZbk9hjODps9kJj4ud3CnIDOrnw3Je
aerjJdqBt/UK4LQbY0bO8rqRQOuV1TeU7tgAwYXSlwK63iOUo5Q6zQL68ajNJeg6jcCGrjnG6X1A
19cE3Qy9d/0rvFJ/bmo7WOsE5sTPa5y73qZRYYdLoT8r453A8TDWT4hUR2cHPoxZC/Yg4Sr8fqXg
SVElQNeh3SN2YeA7GH4+QZ6SIDZuhrz+ZFQj+rtnsu6u7KMSlem3BJAhgDoSPUw7dQ9IvMl4+hA6
ZprV26VjHRJgWCQOoDK68DFncfz2ELzyHKG7/Lo+F4WOS24el2T74IqqYWO8S4nsn0VE9pI28zzd
8OLNX1iO8hYVMKrcJWLCZdH1KqRlSn4t1ADW2cbfQKbSSVwGhhiza/2b7Z2mDxpeOKD6UPc4YnLW
xBx5sEy9fyjws9VgVx6iI1elnl6XDsSsDbmsk3gvhYq1CzYW7qp5fTOyWG7xOp4Fck070AFW38o8
YUuuJXE6WnPHG9/qgqSRCYT6uiP5VNf76qTqUJhXodxcu/NM2LN0pOr/7zZyTaVMP5/TCQAYkJhK
VKbXAT9uXut+0wk5rvBs2T0FC8MCwpRhJEL6i8qIsYQWdAfid5oUrgOFVAENTljDWCZZKapGmjFR
2JQrXDHRlnEg4f8vOXhPH47qARMbn5dOazN3bW9YCsqqW9eLhA9atJ+mM6ZKPFpLcqN1Wc7nOpvN
RnkfkB67E7xVOWN5mSPF2BA9ZPDY75DPoZwBk2F+55DOL5xB06bYyFFz5QUqy/1OhPsx5tc2d/6C
ooyZI/LXdBXz6G1u40ZwHrBEX6OEbwU6WUpZH0JqSN4+yFb8RmBSrkDd0zNY6AW5ZDWhO01BF3h5
Tk4oDdd7nWCpsou+KX3wvZHLP55DbZ7EX0psnTWccBMR2ZnG4fWlRxNXkzTGVA/ljCakGqX3zN83
WqLybkgKdp+lMeQtGkAV6UF0W7qgM3o/FXlIG7kvrcHH+HdMBfviUkVibY0ilikwlWfWITniQksW
2JzWVoqTXwqOJT88cwHLDGw5WYHA6R3FXvY7ONnXA8o+n1PjlS3//Ilom1NiqnEnzrLhizXAdXL4
fAGQgU1sLQ+QMAh/Vvq8CfXOiSr96tPVa3ma37zTb0j5RiqIJIsDxwG+e+Wz2llEyRdCObTYr20X
UqalnFCC4JjBGnSmOSYR/imoZ6hSOe1atL+AZQWOppiLXARXLtnNKrD/xh4zDcJ63A0Cxe1yTRa6
Jsbi2CsHiXGuM2dDYM4gESmweCge6app98tfXFhpFPakCv1wWGef9/VGloKcwDdIkC2RlbsrP0Ns
Gmybjm27E2VnNHKemrvoSrZJj0CxJ8z74GZK5XbEEGVqcAHsRRPGowhxSr6HT9xfeotieLvmB/Px
hAVlea3+WAiZK9tOK/l5L/KwCE26La4QRK7QmFty4vO/fp5qLASHFfMPj/8tCJ2bWsszcnD4QgvL
d3S7IUdR6rOFxcWIuIirF/OfQsndOK0n/jkW3oLqIQ/c3UYRPjSMrcAhHaUUQz1xJP8tReoy9Nwj
Sr3zD/nOATTKTbukrnhPCMZQAq9iN+c4TrjsvSmW8t6zOd3WaIDEJ0K/NHDc97LrLL9LOzz1CoYP
RDlB9Z4EQLWEnln3Gz/3MZxxkliXtD8THlJ/Br6AbfQxyStesZDUC7fE0eHaj4kCz/V39bebk3LD
5yAToVOnshDuSex6gLb/pBVTIeyZvrVn8GNNwOmhjndAAQa81bIEwcQnkVnDPc0Zb/0nwGdrZ/YW
p/awwaNbEdyydgVH2aQNaNen4jzoAMPYljniOJbVysfyEEXyUzD+IDWnNh9tvLbRetCFYtraDfn6
3oc/K2Mp0ZAriDpjXYNfndYyk0uNcIys+1jXwYPvAMCeusgypsr61Cg5TYh7CDPHDMP/2WX9nxDA
arVUZfuFW0CEjn4x5+3KmsrbDtcaXWWtu279b3HGrMjacDDieTTW0VWs7hXmut/Vi9XqYJrPpc7y
pILe64nJFW0uo8KxAGaarPoAaj3veSQ+cusBzZgjI8flIMr0Rjd5+/QIlvdLUN/pE90/GOxBshHK
hfj8Xdz1rbEIm5hxUGbxJd+MoupYti3L87tnyqCQ0/jFLMES32Tq9jBgJXsQhx72vycnTiwnrLIR
GNMGo059ftIeMiAcLynJVQJSAb0jCf/WnaS5b72Mn3x63XfT/ArpDGtUAEJ7UTclxpBnhpKDdL5i
uIBpNYelu5ndSDbX+QTkGkhkJ2EJTAQRFB/8Tq1VzxwfN2cSVabYYRExa3m91IPHNuefMyal/Y64
Xbg0caU14yzyoIAfSOwATybwFYgG6z8y5EaRZVxZUmaV8ogLj9OCMkHkHD9asohvWiG/L+Qf+YUK
st+P+mVHj4xF1adRPZ6cwThCkfJfyt96KteY4M4jY998bYTod48k7XPbMQf23WUHuM/FGsBwEJfD
ANFiVK6paMUXHxCZ81nAsCTQLIy8szIZ1tpGh51SP/1SBYAOJtfUXhWzpS1Gg6rHruWnSXaAbASf
p93S3NyNwupG3uc+BUb/nKrImxrhFVYwzhMLTy81jmaBcW9Dn74NJ6Rgvt2s57WoWZU+8e3lEb9k
9P9VEbBE5eekcI4kzQ1Gb/aCwut6DYjGKXGgaxHHt9Jv+6NPWfPclcFF6xeLkMO7APWjjbizTtZZ
03+YUPytYI6bJBp41Exb6/bvIeQcTNWC1nXO3hwOgBDuWt+oDGBXs842ZTkAxx8NZeLNdCHUoV7t
fViyivde2lTXoiTzasCGw489u55EbEBdw9s0Giw3f3P0eMKIQlvhoXBEDisQYpp8pndE4ieo0h9N
6uKShzY/7nTV6VDEMxFL+qElQHNeGJN5xPoL3kOzeoLzc6/03uiWSZf0Ox9/GJXUoh1/zdYx/Bvc
etbdumDYzXwVqL+Rn3dreGPDP6Vt0n8yrnaAF/Fio+dv40Wk10mtWKjTiTtYYl9bo9SzVjZgS7K/
lEcqObTGMsLaZcD/G1JPrFvcnM7ylURfF4MZJflnygxaiXGtz+cA6DEegknkjKsBdquSqTtP8srY
sv1Rtt9OHfbLaAEcNmcjcgOXoidg53/lVQMSq2H954Ox6b2y8o4KfD6wF7shJwW6BPnf3WxsTem0
HEkwTeqwM+Du2Zv56BBeKoCNFE9FKW20hgSbHQLM0A2xgn3yGJm7y6AWTOmM5wzPIVE4flnxMBND
yL8nqb5RR8x4/HzG13kJ2PzTUZbOTcmeYPnulbhsDuYWtN6qfapJlz9gnaQMR930NrbtYq7TQ4ao
BT+n9Bx9clm4CX6pZcpU7J7l4l8RNRqXo54atENqq+zGPoGzC+hI/UwVMRHxa9/9A7vnfq3wU+yq
OTlrn4HXdwrq2vyeUpA+oktkPmUqH7GMEruKd8YTWoYSBiEo6qKnaeEW1dHLM7pVw5wn6zsL22BE
usbRCh7Yry/w3hls7MNi7ZLu0V4NCElTBZEa1D5IdcG65ncTyGLMibIIBTNcxM5v1wR6rppSVwDM
xLcNVlZSSsb5MVUDAvQ6sSWzTSOTR8Bl8hDTqtl1z//7aGFu+05JrJ9QfC7KHJQGze/fyBljQiye
CWDfOXDUKk3CCjb+jayCe4VfWAnrzaoYeOig9wM7fkhqMq6FxQ8H/mjU7hMP2tLUTRMveb0d2VOa
kF65l/OV9cp2xGy3JVs4oCvPILItAzbziFRReiX5fKEVHqaXb3PynRoPowZbt56zorXsiVtHrMNh
pSGzKQ32hC9ApMUY2cg/EGRUGpyLBmnVUtLHLHuuIWgQXhCKa/2Qjpt0Y7qNUsYlXVahcOrZL/0m
eS8zwqgIeycPGVPe8s5z/amMrGGYaYZMMGz/JnFat5KuMwjkrFLsjbSPcNWZdHxCNrR75ADHzUyp
dwY8KfbslB+9MrWz1ERYdptjWHo/3e4rvWTqiR73/GFSgY6Ot2jS+G/kxKF2PGSnyfeuO1CDjH/H
gUG5xr8D7aEscOcGfoAeFu6Fi/dLPeLIML1nkOnf4gKc4cOclzhNhhb0Jc/i6G4qrEONoR/0nCSb
9z8ajyNBZznab6vUAVTwRAkDSQpsqyTb8+aK+C/V9Ks1poYIULxRPADvx0d3QMmiEIQWgpUdsMrP
5Ug1EbWwIkHcYdpadwZQqxc7TPRj6WPTeVWWoKQw/XKSSsPjuyKcpexhm4/DWPh6u4iuZfwR/0Qc
ul8RRoQX7eRwKukagkeL2/hnQ7oqDh74GzbG7fUbUdrF4SQeuDP2C9lBPEQFZkHCmha2OOTNPfs6
wx8D+wkI80wTysaAvnGCz7RdlobydpBbzzA0RNA3X6M/1Ny6WaHzgdxv8WNlkdijyooKqZf4yCKZ
xq5ujhAYTcXVtW0VsV3XqpP+7oySyTs7YW9aFXDWZFGQWid5g1Lb3znXmqvFXWakkKE4R86nIZoT
1tPso/O0KxINkZzj7VuTe3TUaDESEoG52Y/ABY7h3/dfv/FC1xXndVsp/loIdOQ77ltpOH0iGk65
Vw9bxD81WWkWZClq9FCW4JgzPuMR8lizwAIAXo1ZuFh+6/XFX3IavXD9dk13g0pFIDMvHCArmbdU
Nl2vtBEeO2ArKCn8FDZ0k0pZqkesgiMcoa2uu+xYgp5E+tLr1SlbScnLdh2aoRcM7VKDvxIlXt7P
VPWPc3BHmdcPI1FcTF+ssK9FBSbnJFGz2AzyAIgU3Nz5WX2pAPryhBiMSKM0xinev48IWXtDkpKn
sTOo/ev8oby//EqWhkU1wuqy85q7/eBit1r81e/FvI7rpD6hogjgJcdm3+Rp86NZLa+l8HCGA4u3
YOVUNgw0nGEhuamDxgaEZOcFd2yRqqvtR4n67G1eros+xZ53dm6cNLgPJjF9WM/R9evZHy3IrV0x
FWfpPn9gejOx/pItTwz0XXg1D2v27xoV7ssIhQ70EBdPpJ36mexIIulKyQs2Nj68dYbVNw6Sifkg
VEd3870IpWSDbw+1Cf9rSUUScSyUlWvYfXYSeggQ/00j0ikn6nf8Z6XDqSAYhCR9qcpE7A5wGWs+
ruZ2M8x49okUSyVIX3OhU03mXG+juXJCdLPAhYkqEBFFM/+9Jw81UgFulfacqTeseyuuFPjNhhpM
kmPRDLvxL1I8RJqrMXxvrnAzgdV7/XHXT6NtkscHoVBFXLHRWZvmNABngmglkjfxZQY67r/BJEF5
sLHybg4p4Oa3LXEGj4LqgKYQZRKEgKGHwQxaEB/h4nb0qdktdms3ezBhxrsrKIl/dvFMk/rlypFq
xaVAThEVP9Lkf7D47a8FJ4mcRsFlQNTOIoI/4bF0cSzNrEEML3seODXkdapbWunAmlNPocE6FVnY
wY89TNYmkiKt5YSyxS7AYbjNRfE2OOq9ZvikxIFPHXCo95a4qZT65rzwJtkTjLh1xaVndBZg1ldY
KRX11oGhkIVBzW/5TJPD2MY0YlCmHKhjWmy2oh8S+VEivmCezcQVH5l8g6ucjieBAVigRHcDWekN
YXB+1s3vNCARmF8gKQ1p1JO9bJ3lKom+1lZihX28xXlTcszUCno9huqbkTbRhHp83R0tAavQqH9C
u1E3YsTqZbTXVAv0nWqyLnHn+DcFiCvA1s/tccHqk7wXkJPDk67QC69WjDy68cpjX5Zsr34PGsLS
qaiNboTze5ZU/SgTO5N2cSwVsl11ZSl0Ic7nuio1R0T6gqF67N91ELi7asi4FyjQL1oGRe/rF5c5
Xo1bE30U8DPIQBhfopPzu0Sr5JQMbxLOyiU7AJqBAwXsXBgSpJ/veUJktFGg+7fHKbO+hbalvICB
ZTrff6d5hRETNBA+/bOFeA7m44y3TWXuAs5+WQQcE5+WzAPtKM90UsC6MxCFXic+bGbNcMcJ48LW
hMuCPfjskoKtyhWr01Z3z0NSNxmCa9zfweMquMPkAsxEbtpVDoynT4sIWWTJPHYbbpUQmSaFXXLy
U2Bl/LUmp3yi2mQnqeUUvlFf+m5MVKzep0G2kMr/jOB6BQqmRSYMiAYWwHkdSv0CXNTl8qz/q0Cz
ztLWtGVcdu70Rc8ADbRhEMhSY39z9vmeFAQ5ZgpMCthk6LUXdhb0D40KjQV4nr3M7lnPBdx/1iUH
utJ8fRrbBrdh35JIWhQsZoQQ/zQGdDLs3XQVmPor4t1bgk4TgfT5i2cYlQnK3spf964/D6V6wwpp
zGbyM/AHq2CMeB91brLybgSszkoHQODytZzEft4F27JNySXsFOvodP70lKCxFw8FX6ZE5X38zkWW
7dt9/lgUKkvfX3UZgf8oslq5wVrY0lmOroWeywYB3J9QBZU4SKpFLNOGBMhU216t+Z1Lglv5AvI6
6BIHIB9K+gAnqEs73g1U5zyHcqz3txyZxo5n6YdHbewztI+5lq3cJJlntM/wRgQyN17jkj8fI/mp
f08Sss5F9l5rvnLSaHiboBHzTQp0Gtrz/Chg2zSzdBl4U5o0kFpL/mCBP/QaUCrigbykwjCi5mIg
AQmmSvhhoal7IXN1/yIkV+Bn3o8E10X3XcKbGPyU2Vb1pUm8O6xZc2ROifddhzTY19mTavq2RFGC
W2hvSEIQBV3TK2Ntc30LJ64lhgWUj0ez4ALCv0L+FvxjCS3rVfPqtPM8WKngiW7nOzaPOQY9mxyj
YSYcGSv5137IpXJUq8mQudMYiLmFKU8ibWg6vFaKhECfdlMosnv08te43pOdLbj69pkhspX7n5Qc
3cZpidwK6SeL6y1jubcUVS4dkAnXCffngo8GsP4N9jh5CJoAjqaIlnrtbJWNesYfskS0L+iqTeL4
7f4Lz52Q7UG3udKjQlEa5w4B6qu2+A5bSkpZWcMoZ09h7fFiuPlTYsBTudVWt0EQe4bDoSu8jbRC
R39YgCOuI6qcCaibadZwEaitcwxoLJHyhVmGlYuyh0AjJ9wc/mra/uMMtLkwomN0/TgXNcuMppX8
8MxD30JcOTHzR7dpfskC8VSqdJtvqQ2KkV2mZAMMEBE+kc7q89sevFq0y08icw7xwJJEMlL4RI8j
m7JJ6UqxehJPLuR1jY7yvy1DVg1zD5ILZYuk+E5X4ZLf0+EblhckdibsKgvOnmhuV0cKImaFs6Jz
NaTzyB+Euh5zsV/qIvfEaqDWkLNmU8E7KnJrf6fkWLVUtHgyVRrf4GX/2OcDuCQWrllC7Y8rWhAF
wdQagqoM9xE/MchZYMLqzTujA56MT33hiBdxw/cRydJ2FBtDi4fIZLQzO+Il+gE24vumi/73uSCo
D+nRbTMj7mdIjiFt84BEBH72l7jtVq9BrvpnVcEVso3FBjtuZzbaxEYNFgrgjld90W8xiwcrAjm3
OWNPGmi7LKK1bl6jrPuzGjaqY8XBkZUvzhrwt3PCO7XzZHBvO2Tc9YeVhk49CcyF1uzeGzhs/lnA
DL2cm3mfg0G7geOPDurgpYq+e8ozBVF4cB02ncyUJM+3ZqeO0I7EIXni+j3LYOAKhAE/YPMib77/
V4Hna2aqq1W4TcfP3FbNSFZcj13FnR6xSDBNaYcFcRAk5wCA3aZntX00+mm6lI5983auTI7EBVID
hOWhU6D88QxSIF7y0Qvj5AdgHDaEGn1kfedazhenbIznXm9b8+KfVPhVpgxl8M5qmHTok+sUVNdP
Gj5Y0vY0Idgyeg0rmQfrPJBCrSVE7/Nc4KPHEAX72VeRiSZT8tX5y4tB4UsI6JsI+lmgCFTeWJWB
X7K0i58i7KzOtamKB+9fz9RjjWvMxDVzSOxNUmrXYE1fxLVlk4R3ydB7yQ5t4WxmvudDln4rWSkz
QIauodEyaDlm/fEnyEYiVZA0bmhcXcSQ9HnihBTWbGeaZCjAbAx4zLAGcQ==
`protect end_protected
